// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ZM2eY/ukCymbWJWYCt0Zd0fkWNLixECqdDOJu8zas38QdP3haAf/i8xg3+ChPnLk0wyEUDvP9Q/U
DCZ4PRP9IXyY2AQueS0LPUTigxHc+kpRrUbjusarc+c6CgnXujUqFROUK64FttlX2ru8IdCWmDlS
ShSbsYJEOrXRZCCZ/6LBmfjBK/xx74GytTM1fFbv51FYMPVIYtUbHtpsNfnJIJf7q8/+AUuXQyJ1
9SANxC8SrEvjOsvwi7kdCTpNSkfY3EqB0y4cKHI9Cus6VVejgN8GWB9Tc8vWcPI2sJjVCmZWhSPr
GIOmypgeu+yuUA4P7FivV/znzyuQAFXTfggHLg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5600)
XheZRDsWAuxzkHJnQGhEuJ6y4s+MnXtX6XUvqJhrRfdN+ekpmNuxlHcl9fp5rF9ndiuCTDIfxko0
FTbpXfBeMCa91QOn1gTgaxdt6RZoLbLVGwhVymVAqAv7NvkKT6W9up06zRj83sQdQeSDo7V2PtPd
dFV4qbmrSn5mw4PfdVZFoGJAU+5TLyFUlDQ4uaybF/CE9birp3ZDx/ZHhxLtfQudVfjV/o6BAQu2
dh/dMuFZRDIYxSbc3q/kco+1GqDToiCnOaSYIfEMUnncqkwEW2bFvHFUt2SKXK97FAhOxc2CUd/9
8doSB4q8BicCVnq+Gxotzs2ITY9NXm6ZVX8e9OXVeInkUQ+xvw9Xb1Z4eU6OdaCG+4ZQYaZOzQ+E
f2wf03bWQEuZqzIemmjdafIQJhts7yXOHJhZqAk6QImywPm9KdcuWt2mpB+NBmDkNzIT5Ke5G15I
gRGgULBp3m4jCVbEMhxiJH83YCHg/Vk2Nm0z5Lm38mYqTXww5Bi4KgIQQOqSsh0Up8pD/WDRy0EF
KIAV67lXuRuI8y8QqpUrrVicgdfq7UMa4EIyKjTBXr2uQ+Bcwm8eyAvY+dRZgWCDFGbrH71uQnnc
f3dNP1eQWoUypktOG86aQmDbANvHhx/xD67HKfUakL9Cj7Ikq46RNAdy9eSDubxeiHmJBFeBQvZp
Fyd6/6/ms0PU2rd9iT03Qi0N3SK8hFCkJV97/QPL/1xumAV5ICES7pWK5sxy7fs+HE3Yytxyix/d
z5sTLwJOYWAPYZvOnCHuvWutOpgdxkmlQhfkEKA7BJxdKJa+T2JHV6VevNujZDu9XhckEg2rgi4Q
BjIc4uZDxm3+E3zZ0RTIk6Mnv04Miu9m1NHprUSWpvbQkRdxOuMGZe7pHCyncgMV21VzCksaBuJh
55WwcjVop6hvl4aoCQ+NzqPiWNpTD3VUaQ25Jw1gRKfMkKR2oU2WcXMsrI8H5A9H2RRAc3UJiVgt
JW33pem6DmkV/T1PTnJ9mI8Gr0i6nKdUjftodLgzhsM2Q0uu6+sho5rgkJabnsOZhNghC2Mngdke
SeHLuIw64uHpezcnJN6cZ50c/4mBuQdyWxHosB+LgHv8sAdCNnmpSJqcAzfcVIEz+5iV6KM31xzg
HD26Cxnc5UHddtOfU3znWb91e26zQHcqkvN7ZFUFWh/edurYART4nWnmXxj+ODd0jwKiIiqN6KV1
75yjgX7wLWJCthyF1wR3ajPi+SeFcTiNVZVcc5f6GlGb7QByZSReInlfH/6JnTHQShhlHyY7qoT2
3QX2UoyeiYKjNcNK8Va9hWfuwz7u83vOl///iMv2Owa2VFFH8091n234sojuoASPdUs5tjsZvxD3
LMi6105Id/tsUT60hCiEqjht4KRtgPSX4QVTM6q4Zn835AV8t6lrRgeLRlLGxrHdpX76+QsOxrzI
SLsiktEmdDO0DMXKa02foPnzKJ0TOm/jPVgKv/MBztl077fy8kBmAwQiVNheBI/1ZTpPqe1lDtZt
BQk/Nol+dAZB7/AEQ1IO/ByFCBy2MAo6WZgBOHeBEKI+lZMtZjBoIArDlECBZQ7zgQaSWKmFBB1H
5pUJymXA/+iyd+vF41ASF+8kloyz9exnaTHWwNDWVdBtVSywbkf8ftQAZd4Vo6A1qDM45xcnPG2d
nqK3uUdBXapDmDdWgv/rroJhqa/PbXpVmIijpKg8dpmN4vpRhbBCqIWTV43mbqoqYIDt4KSdA2+D
s4sBUZSw64Kd0wtHcU8NPDZq6J8zf8zl8yw/unBjvTRf3wCu6rVMRzjJItxRQJyuQSkO3c2Skp+R
Cw4a/bgAykHsuFegw8SDle3WpTtv0tmZJcs9Dx45ipocz73BkS/6FJj2Oa3VOEvCWq2na//ol7Ya
+VsvvaAa4373rZgV1HmHyNDDM7+0NCyrEHtK8rxj+sjZr+cn2Ehn5Cw9MnkKouN07QEaAZwPFHje
NcBdpv0QB4YK/CPHnUe+gaOc2Ip2+XiiD9+djTz9gxahyiIiSHt2nrc3qN07qIQKIW9CP6QYERZt
tBdfKXytmJ9b4lqcWGyV5+LlOsHczwJw0oPF9lUBv3nwHIlhzyb4zQOK+8vtTF1zg8jGLI/1sqR6
gSwQ73hKUwsTbwgvczgxqdpnrM7mCNvNjr24sbWGXyUHkjEM/46Wag7Cq9XB8gBmqdgS4fmLCBRN
ad39QIKqEqH1EUKDDgJAv5q6l+eVseXhHr+5sHd4U7NV5RnEPxrHsnySuO+3LE0xOO69rkQvolNH
+v8p2HTFedU0J205dDvRjtT106nXWMoSRk6I0UL3xz/YdG7Qczf9vDOCdmoUEobWfnspQsFh4HuT
R4Hxc8D/9v+YJoNwllc4DtmAmwQ6XJQ6dcIZ9OXjq2YMz8vx921sKvNz1jH6UT6QZEFburJzhln3
QxwpsuE8GX3+uER7KNvzDNHgLFmzDsWfNTCi86dPUESaH4ohawOKvHxbTyE4zoZ02jYyLqw/FGgh
dGCxQJS1A3U73VeuCG7xDWn47083PGGIf9mZl8LWfXTHSJiDsiY+fGYCAMBzQly/+8RBUIW58XZl
XjuDzaJ6zvDotuNMIMXvaFEQdRmRRJXWjc/CGLp2NtRhn8m9iyULc+Ii6Um0MGDPQgcQTFrgJz+m
mQ2qlBiNYVj9B3ogXLvwAupO26MS7NX6ufXBzY9m3Ro/SEtbei5xQWHRc8t0x+lWD+eEi3FDeJQz
6RTqyuADLPUBSKzMcAriYe9bLR0z69j77dk98dX4di5fKAWOFjKFof4fWniOu30Jjp3y2KgIV/GO
y0ZJhzSiTQw+fM8QrmuoqP5yN6nLtKwb8vXYSxBSrVXJ+M0U6vXc2TfJUvVJv5+Z3n9oPOT0cS8a
juF5/M1dZp9h2737hQ7SuqH18W18QB9AMxWWzpnbpC97r5GpwHIR85VDhd1MHtqs4YPTFNWbYW9N
YBB01vwuFK9NkGBzwnO2D0TrT2P7mG2PBxFXADZnhn3+lirdiFGkygjk030aYgolFUPgZc2uwjfM
74r9dTkXIdws0fiTTz7X9dyto1O0kOr44t/pA6Hq/ew9dji553D320LkID7jbxZ6zCHIuDyKlnNc
Khh9q1CW7v4WGwrAEtGoCzTOljR9QIFybKTZRMtk1BXv6e7gX8XPYSUq2RaEZla6v4GCTMxvOqq6
odGB58iD7+a0hAaTmt9wnqrhhQOUtcmTudnbHfLw/UMKnvZmuHMv4t6GS9b+CzzeJqO17kT7VWMO
ABRUIuJGRtN/N31+5ZM5p8BV5NhwbwUzJlmmAYFxuFX9e9u/1InvTxOtMDfnmsxk4rypvm7Z6KSf
o/o5MayhoDyn32EaZZmzVqWl+jM2yrgysDrTZjgXx4RwbHLnSf2MyVCsJje6i0eFBUsNpNtij+Tn
l32UXxpPAZr9JVoNxW/SuARAo1Yxu/ccqJ0SRHQppaLftQBV4For4hnVBmHcP7HMbjruYhaLMD8c
LnIgYGE+goozf8XYZz6ZJSpCReIbLL/+lsQsgkygLRWqBDCZYg9LYDr4DQI++T3fNPrBS6PZ4wmd
tx8tX2QyjBNVGgwCSCKOtB4axrrRt4q3fZky85E9mOTrJHcdIDpjPRE5PCcaL8GzNfrxrYM+6dkK
CMmDp3WlzhP8H28TcSfKzdnzH5vbHZ1SD+Fz0O5iAphgTgqG3ML7rpLw0eAxkgjNhxSZizyFGO52
4/qeCICyl2a+lhBo91nicFXB39eesmAJLkiYPwNETAevt6fu1e/Ip5sRtX3vqyETbRI0vtsmFXyn
+lSIjWdZOodRKfh19FiusK+FDHWybS8+sKyBb3A0ivYzy9d/0I743xxbZMaLiQ1TMfuP8FpzgmCY
Uh91beD0lg9lRGNupnfx80gybB9TqakXf+7+40b5jSnFBbDud5GUNxbfrSa7hlXAwh+3JfgU9B23
NO1SIWBE6cysXmECfLEIZfM1V2MIV0yX1wRqEBvxWxPkuv3F3rjxwW57iTyVObg2ptMUz4/nuNLb
EgACC1g82mgLdjbkkIjeYOD6tO8Z/u1juUc0X0Zh+wzew/TADY0cvgSdxwWT98ZIGmB/T28GG8li
EV4UKE+WZ4M6ExZopmvxH9sfYrCLa04Wkw8UOINFKcwexrpPyHnAVkm7JJoxkx/0eTZgBWq4aY9D
ntDKbk2v4IZxUmAHJWXFkig1TBklQ4tRNbHPokr4U/51yl4sUF3rJ6adfAXhdemLlOVxKnCYNEOj
ftchSET5DwAiBdBWVCm0qB0z/xZdRs0xDLf55143XjibsAL4CscYiUzcBbIelWUtxFqLeVKbUE4N
E8BFLGDTU/e+U+wSEZ26exRu/4TrnLzop1nrufo3d6hdOWMI3MjjK2vyUpujZLQAujX6CGtDgxK7
zDctIqAdyinQrqNouC/iPJLnSU9AMad/SlU3uAqd/Ngfqts/QGxoCyZG+GqVTtvg4Es9kTlUbYWc
2c0diJUonYH/HPRXHDmzSrHtT4i0meZT7VqLbGY+n0E+WstZFRMzNx3WW5+AA/oA90t8vrz8i5Y1
2meROycAp7g9cyramQ0XHOa5wG/co9HZ8UV1y1HHrdnhUMIaRkRtyfLyWtWP2hAR9pKRxoW5GlLj
PijvGv0RXWaSgf0ZiycCgndOLYGWB7xJQSleezXsPVU+m8ulOajei6ngUzp7zq7D2D0/cwU6k7df
4028HWc8cKB8N930updLs4IUG1J4wzcbzDhtEBhyFHuc49CaAtD8ul8g2pUr7tk84DyixXYlVsY/
XFwigQCr7/vI1qpcwxht4G2PCQ69g/A7sz8ax9+JiFGIMJjkYHt0JY7h46J/Syw0goQEQ6dIsk/k
MHn5srptiAPzQI4tjKznqqkRaz50P9ElOtWiNu9e+nQEbzQDaOdFYNrZycU1FSU5HSJClVejoPYp
4FZ63PRqgTBGGmwB7X5FtRFvgX75EClOZQECXc5Wh5wtordfV7V22SAZ/qNFEkaOJH914aceDC31
QXCKW/GQ/5+a5HwvEHr1H5k7j7WiTcqapUDMQn1Lrytcj+UQ3ADHSw7C+oNcpOyefif6UaFqSzpp
SeqyuUtEd6lEApkX5hVEpePkfjS1JBQJMyamZPsGTRrrk4j2Bs81oKQfEdF75e2+ehFsdNwbemFW
L0U3XT+ATXwwW7QrKM9p6f5ebMufWpz1q8bJal4MYDtyig7yJNyCXTWtHjw525Em41Q2KgAnSBJA
GI44RmC1+XG5c2I+QVOuAP+eDW5xCqvXiVUdVN5kvqyMO9oJtH/ai6OhWQKzGZiSOkOUTF67nsSI
Vf9uD44z6K3zlxlq6NaJWhZz5ZdI31hT5to1mDoVtTpQt5NiCK1HdKIrAFRsdmmKnYE7fQXDl/xM
hX5RTIER6p+tFvDb4o1gu3/lBgjcDAypDbXGaV/fjdw0RteoLc5dcT3GQMsmfEq9Z9yM696T7NM4
KyMDnNZAPx85WWOgVjy4BN1wGh0ouBBOBG+4DONtxTC6T/j2Op2eQEHa07v5lF6eGjUP9OYs04n1
QxYftHfPju2doabboZ1KE8sSwIclzlmtWn5k+2ZKc/TxSXeRRfjyRCD/4t+z5MBRCqJ6Elwf+Q6D
rFkJbRQuj1vH+o6qpv7t03Gz2C9bsVCM6lIhN8VvfNDc551QNzSkX1u8rp6Qbn5mULv3iBKeflbp
2DNVoNsOsCOO9L+g4EVARIqE0AEG1u0YniBeJa9mvW+bBiv7jDZg0FaW5E4gbIAfKDCC6oHSB3Wl
Erq6xMS2EsnfWMqiakBDFxCaGRbcJJlvraGnVpLhpf4gt42Egyc1mjto7FYOScyQVprzjVwsyib1
Sud+EAhFgExuxTFlKMRHpzs9L5dMYvkNygQNsF+DydOSI6mD4yRytsRaJoE8RBHI0PBst7YiYyCa
KgxouML6uHPziz2dxBezgjAI3OzQr7LyV7f8Ecu4A4C0yAOks1BIhYqb/ObaIxAtQ28gpNvTz22R
zrbh05SNSzJ/eACUhuAtX+Jtes70TL0PXcY4IDHfzf+61948TWfvxSiBfi9W3WD76lK3hPOIpE5x
5hxvsd+93JoHvv35zjNd7XGH1c5k33zcQy82mui/vWuqGP+Pd8QMdWWhcLMMEeX3Hnw9UCmLtaQD
e6SkniBlO7inzsoRncHOfGGYQLX6KvanjeZ+/M4TTQVho5Mpz7L+8YvVQAyy8yDelECycmgET/31
P1RpeuaQTlsbakE4t3SPX9lNTzW+KwLTAVcne+olK2WR+WjBMD1mpssOQBppNbArMtAx8UUax0iP
Dz9a7Kh/qyCihmrZstAclJAVZrLfyNdaoKpSNXcp4yr6uvJK0PKZBWuHb13w8vLlBwpK7BOgegxE
xb8w4c6opFvkzrLyX+HlXdHehR8Rx7nc8NDdX6BtIZyzImMW+sXaHqXvnQnMtrt37+pqSedcgscv
8UIhE/fTc63wsv/acaxy7+VnscWp4hivJUcVoaU9/UIsEi4E4ecUZIdV058IIlfYSPdjzV6g8fbd
PPCcJxBu6pznRHCx32WE3MS3+zZen1uSzacQdXJ/R/GT+r3qMbcnXKpRLKMvxFwT4cGJSvYXrvTb
Oun8xJRKc9UZD8b4O4Db+4rk4Cdj9k5LH3IB1Df7zrwJ65TZvryexYTQ/PaBh7q23pXjNJT5hONY
CetFH+1gPtHU3sLZi25X4SUOySjDD0AHHRq7UcG+RIk8R8Tl5QxuQy5pVHaLUciWTZaR0cchAPxt
bupMCwyTtwmCvEW7WxXPs7Cok20vpI+eWuRw/ramiU3y6nqreu68nEQ5MOyya/LAf93VGr7h2CCQ
kk+45THYAxhSJtIJrISjGHHBwWTBSaOLLyu3calUdu/n7L/JJbFpxgKAD13tNdVX6sZXGIs7saYV
M9VfoMNy2H1BD/aoGu1NxYWpCzxJMvRX0CBtIB9RdMQ4dv9g2jQTWiW7PD6mLSMCLNZC5pBtQT0S
EnO4cvxs9Fc2LuSQKq+t8e08cooZlAWrRBFCFh4wZ8tDk0aRSd0WMG6ZlwTePu12S/bOTj4NAGSi
I591k1OJPi4er5Z4F5erjc5U1ByrUDzvn8pyYC1/Uf0lf78z4ChIiHDHTW5c0rUSunmR5B9D6BN7
LjPNKlb1CYws9FqnCQA/bYdm6d53KU3JgYUrTS1leajP73+d/nWiD/4t8boKjkl24y52Ax8U7z33
jWD+Zcu5Ce1cKKu9elj8h8rTnmL6Xy+wwBit9Ay7rQDgHfMvc/7bxY3vRObTu3GdpGhx2MoSU0uD
xKEYnFC1RrUVnYNVlfh3xPFmefS/RcqMn1DSB0HDXcTRle7ECd0fyLdNcMSotPUsCZN8CrFSjMjy
+B9Q/jeDsW8ocAINNebQmmxKajS6WsmeN5SBGSfY/C7wkOom05lI2cbsrttI2UgNHLCwTsE4AQrz
gprV3QbouWxKATVoD3Q=
`pragma protect end_protected
