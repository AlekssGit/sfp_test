`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
UrHea9Q54HQDFxI/ZsqKPtxbZ6lfBXb/lBF4/4O8y1qXYkHdyQnoaUBFl6IuElxV
KsuKTBotDzidZul0D7F1idBkKN65Jsv8D0zEd5N+kUc1sYZSt2pE6vKqBCtinCF5
sZwjUNEjHA4/ykpcuCVbc0N+79pSsZVdeXZLgGixOzI=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10752), data_block
mPFXnUvmwcL2vDppFTS0jPm2deggSGqgZ9xMvJqvNIi7sKYq2Fep+Kzkc34YB5K7
WxMt3rpCSanXkFwgmyZwLcz0dY5mUyW7MUhD7gFzFYbb9mrLbkq0euT/ClCWl6no
hi40qPWn18NJ0dln0Ta74VCfFgWLvFD8p8gT6ELwHpln7glYjTNwddfeoBu6psxY
VP2hjbPGKQMcZpNHEBflS3/W3YSBejE2H0pR11rusJSN6OMXXPJvYS7aS1+TDL5D
nIbevygOd6nKsURjjdxgqkLsRXTd1YI3OsR/yiLzohYFYY5FALSv+xZeKWGRX4l/
tWEwTyPYs0v6FLAvpp340aUFN9k38k/aZ+5opUewJ9jeXr9qemDM6rxfbBXX1J3i
4GcQANY8R04iW+/wwQVPYfDNh8AwBRVrtx5P1id/dgI2Ds5xXTojoRKolRO2HQ3y
mm6cjDduoik6Bn5/d/VHix/U3jylUpHnlLGlenRl/wVFa4lT0JPO7sreZpswcwQV
85V9YokS4B+Cv0xRpZf70UW0oUDCs2TN0Mz4D2IfBtq7+aaFU+09iH8C3ax3XlZg
9u3C6HkLgOEwb9AAvmFPf6y1lgYy4ylDrtNyR2aqlNML/wZ5WPF7vUVtFyDZoFC9
MLYji+lfoITgudY1lai57P11spDuHyKFc0cN+RmdOa8fGJ86rwolXa8rSjiEMyzi
Av5yCXkvNZ+NqXPnWVV72lXQRmxs1cPEGw11tZTaBfha1lZJL33eI9mfqDyYT52D
jbnp7gYDT/7OrxDDweyLRX2nxlwbEBqimzIK8r89lY9e4mf+t++JIy8iTy7Bat9z
aBJwkSB32HnETIerDg0hf4BB2eBtDQWWpzxUQMxiOMoFu5z1uhsITe3YXf2Bnvjc
eKHVvvJygGzc2ZRME1BdUO5qn0AHoM59ma0bcKtsUme9/sqzEJJt6dYf+OVxjd64
gQivqgAkrTT5eXZcaai0G4C98pr7Q41MFn6BL4UpT8ohetPcGM492zuzHh5aKB/4
iqgxDjHO4EQSiHA0eKEO1lUpYlGj4vOn6M0YOHkWejOH2lyIpHIySo2+1Pv7+KJM
hrXRKQgS1eHhjf0yyhf8eNwn96bdRGKrq5xZGZIWHTI1eTpFHv0pAC1wMLRK2KSk
mlcIUwSZzMMH3d/MWkpp1dJjEo91UXKi3Cd+rpO/voKBpWIAPQYw5GmX3FGn5rSf
UOf6ATD/I0DlbIzowdECLkckjYQP5MQUrTZSTzuRZL6DnBad7Q8L6TeezI5/at0u
H/wh1AiBBb9KmLSXq4SzCg5IM7JL5Lw+d2HczdBPaNbRRagn3iLZDCpoYWJWPrbS
RjSfgYxqsegtLJ5uXFAkcK2rwW/2Kl8xKBJcs2RN1t49VYJ+QD/LXGiB2PfsC8d/
6jD47WCiRvhHmPuJXvF0F+ifE2q9D2OZgBzDMDWD+BLoM4LjWWWJbhnEl8KtQyuH
P3obxb3/HTdJLjG5yYi4GyBNM3p3aFqW1mMFk3y7aT/TObYDjd+ja+FZUMeoACvQ
o/sMCd9i7mGM4ZCK4SDOwrv0TVLUyRIemnxTtyHAE89KT6FOF6L6jr7nxVLYPiAM
e5KHd6CwDY79aTtWlAF7Z39lICI5Qq98fx1eDiM/Dslcjx/U7/zG3XJfKdOZX/Zs
TdbFSf08bSqYxZm+9ccStYggTCY3hTH9Oy3KQcLTSwATeIfcELSVtxq002T+rFwp
loiBJDYluvxjYzQOvQg2EpF46+gOEl7+/FCiCd+J1zq3OZbcr1Ep2mk682/OHKC/
rT2KSdMbUtG+8t7x6F3VtpYyKTI30zvfqltkXaHJA6qPcDa/TvVNlIPnV2ubLkZ0
8MWMNVnCo/GqXGL0rJZrUrcnpRZifLfIqCY5DJfBxRIwgv0ngkBLKI2OEK4vjkdc
z6T/0ykG/zdK/hkFp2VxkoqnhAh82qJkrEzaHd4plCTgT9pzDx3IC3zjI3wd4zkS
yyhkofDHcVIiZlWtyR/zKBxy5BBvcgchRcs4H1Qx8pM/8ZToEt3rzO/hcyHvmldu
GbnHCDAX38PuBiLUFgGQydLggQoHTwhg10KyK9h7kWNV8M7pZfAN1SJBXVsv1M3x
q6et1xYC12/Qg+XdZiNfZRAamD9KZzNv0L4rVppD2gvTgA8Xl6GW+TogTuqHm2MR
35yLi5tjKyw/CuW2EGTCbXxU/hVHGM7jr19lMCzXiuiOycoCZU0RkRi3axR6Plg9
p03q9P1WV6Bqvj3in59f9wm9gsH94eJdAr2Fq9MDJQSORg1suVQD1RawvXE/3gUG
QisoXBkIBHRm8FufWzBg49Y7owW5sb4qM2v3vxrRz25qpjIhfH+44fgl/hqgFPFT
ZIosFa8mBx/39vyn41UVjQUG9SFwKB1yu0coNIMlf+pqkUl55rPcFgA6aU1VVuiI
mNbykFUIeB62k7HfQPIk6Ij2l182aqOpC7AsokiHbOPsTzxk5gkS8YnP4Y9k/jon
6b2MMJL4RXxsAvsDNNXotbTJp6V0w67DoJge+hwYWhF2kfTr/vsPDjRt7ER+I5su
6AGfkgNaXYRAWQa8DH+XcbRdp8sBoPkWUxJ6WVD15yXanc1QBl+fFZJtzAq9TLuv
lhUPyoH2W30ZuTY2lK9qbsc8kkyswNz5IPyH3L4ZVwu99IRh2oYEto8cYqWVPbQc
rwwixn+InXem1Q53D4HylSJuji7ByHqSrtuGYavRjt4iTr7E3vwnnufHQW0e40w1
Kq490W6TkfdLoGaSGI8d/hRjsS1gOAyDvEUoRJV7Q+UHWJc00QWdKcyTTCbhOTJQ
3ahVnAtYmlOKMH/VsbD2pW7EN8Z+NLwsmw2byy8jTIm+IdAfhyMTEyVXEBP/iUnl
on8LTobKmSwLzBatceoKXJe9KQMlFyXKjC5ZiV7l0Gzj5VMEWqhT3VlMqiJb7W29
4dFoA5VfNN5mqx+xFZeRU6Q2imLxgP6mvHMyg+NUbQgFW+LaIx/7d3U8mDvcRPHC
3npiS9qkBZz4kfbPRSynvWeT4k0Iv/gzlhtK/pZKtdtd4gp2819JwqPB4TXOTWSz
JuY2e94+I1kzMaXhPJlm4/eKPXY1aXLfKGSQ054CrhEEDWiZYXTOFGD0Q+w/ZpO4
0vkNyawkW+V0G1tdlbmg7phmIpjwV3pojgivaJvHowZTmqo/3n5Z1iIOHBuoW8KM
BlHY9lMTtYLOHqDay7wB4W2uhT82zLg0ghnopOi00ewqGEelzJQ+ErkvQepLYHX4
NeO1iqiye91sHDqijTJGAQ1KxfCLWWGqSZLFlJL0rCScn/QGks3Jypnjy+rOtG5I
WvSVqynJghOX9vWAlBrG/Osyx08JtEqq4vfvzlyi4T2pbgrnR+BT/Kag6FeLyBWU
bMDal8R8y+xAsTCLE9v8iTHL8lDlWLEkrjDrmVdbwkyuMyLcSjjDGwV1njvPDEm4
Gy2+fdgYdyGWQXkCNgAKQ3UgHFFxIQi5Tt5hHhKOrhCCyde7D7iAMXXcNUAU4F/e
RVUgu/bI5EXZqHJuBFVeCq2Bcn9HI5PtKtFMB8UFz9TV5dtyKVkM//E7d0E/sOAY
A9cncgaldI6/YP6zdaIuGmFxAwbcY2duewgbtUAUUI7+xFxy/yz//1v+sNpYIM6s
SUDH+n3uy3zOR1taVNo4DujymS/9RhlKbt5ZhegJDOa+0QOUv8K470Sz1WNhogyE
BSYdGeWQozsxS984Xx++ZtqV6u5QKUO7KnOW9LzZmLA0q6iGYllOaDxWSqNqSgKT
bNj3Xoll8SObGEcC8E/s+/eRB/Ul2lfXhThSLhItxq2X1YLYtIIgE8JUFCR4PC3+
efc1cqORUBu3SJtg90E0gp2lAOKHhylQkDnvvpGWjOSUZBYz6wICXsuOT3qU1PJX
tYxjtT7PTx0nm6X6tEGsF7G/vW/0SbkLXF1TLMOQlydLF1oIF8Hn0yfYLWPhjDe0
uqVDP8xny4pqY17Ir7o45OtpmBYU75vycAbcMqWS+k82SMugsfXzsKt5Vb9P2trc
OkfeifQhnzzkYN0xrseczIDpT6lpbISJXQwigJvVFk4DwOaM6r3yWFBg4GJLQCs2
sxwwaXpBvkPdOPDh+V5y8/VqXxb9tGSHG4RGH+tqhFObruDSIWMsTJ3lbMLHEjNa
1Q+CHUoXyQBz4SxI6O1ABnaY2BC9M25q84o5jOWnSO9orPEzUs4z5UY2Wr5+kQHN
Sr7wBA3C5xx1UG9CjhwK6fuug1suoBdE3cD0wDX8rroCrG7cjv9xeZFVG3xKL+q6
EHX2dX77QDKzovkJRZcVttd6zVQcsDiqkpBSCDMeICajS3jbrAxmENVw8RlpcuqR
07aCmRVL+KhgdQFmMz9Bi5iwkIwX2/3gP0cMyzqWjRhCBicInk8o+GfEVjdM9Dt2
YDzfusJqIQD4dn4AF7ajsxahRl6mEOJMwTJYEcszZ1X7xdt7nMZVCpNKSp2AJUc7
Rbx4OjmRIEOF08JMTNKrds8e9ZyuEziO3GVSA4jwjK7WrJcakoXDCBDVxAHSOWkG
7DuamwPNNCvRo4/Wveu1K8RRGBtpr+nh0+HUgAZOPJW4z4jdDCaL7hjzfHBfqrku
ho0EgTLIiN+/dTrXnBI1i5iDuo+0++8Ifv/o+9eQj52+eKBw0Q2f5y5USMFNg17X
teMh9TF2OYJclAzSQ9lHWHGdDXoScvdW6kw74lznzfdqenZvVvph3oxD978I5cPC
HGbF7o+bQpRSC4Xjjx27m+WgrNzDkFYe5i/G0/Z7trMLoC4HnJKX1uZAqHuclXMb
0MjnaMMIH8JDGWi8gAFCpjhUeRRMrCfDScyJgKpBgDM+7Ie2eB+R0LMedYW9LrXP
FfFddfOfPZKEHfrvILh9zJyJoJEW12oU2lJPXBoowMxFBFsUIY9LFFiMkI9yQAtQ
bHQ2gazbPCoNxsnK8WOiova5dMLM9jre7thn7OCmCqfSi3MNxamFDU9JtKg78Xth
xjRMgywPa+JnDBY/OVDoMbfVxOeZI11vsW8aSwKQqHNy/1zjz6vQnohV1NAs5jiB
rxz4364mw98lNS9tdn0bMxeyRBpAx5Kaz4tlwh4A+B5QVO3FxCRzEejLwnkIa3xX
bsB2PSvJGIKzv/o3U2hePb7GDqmq7FuaM0wxzXUF8rsFyKSdWSSGXKV8P9ScDz9H
uRoCF5LQkNY3YMJ+L8TJ98R86ik2IgQ1PThGcA+eTv8IcmXmuiQK0KzuzFN+6Z0Q
5/vZacLUTE1x20cRHA33LCQ5GWb+k13rqitYPRTpO2edV1tkPN5hUE9fGtATb68u
ezTcL29lQnfsQXNmdptr57I5pOAGZKJHOP84uLB8joRCEnJRjK9fha+vWngTYx1n
J4eaCl5lk2o4I67Djj2qIqmS8H1ZB/39JKgXQTfKSvWrKnlADRMQJ1bgXobHDmH3
G6ZBWkWRvpRU5O7cCVVqUYcCCxegq3Z/DDj9PaUcYIA8di6c3b49cZ13p07SEbWw
0x6axVYmiKerum4IhoC4yA+E7uXxXclBTQazBTjIOTFhxyr3HYfBQfD+29G1fmLY
HEBAtyNJZcXrkb4s9lEbjGIGHix1yLtItk6LaAMng444pdY8hio9dd9cYsy1vK+D
z+wEJvnRGFsXgH2a6473XklddQuAJ5OZ7zFScf0ZzCKq9WgPKqL0+Pjv/IEsQE60
/kJUq6sIeNPBZ+5c8OXTOmD/0xQcuVnb4/fC0CLkelwMd/COq8z/5mTFQuAdjauo
xp/bp9/LoCuf+5mCPQnx3etN6dAqRh2653fFYzo+yd16NhJsm8eceuR5LEsrSyo3
AuDZP5GYQs/7lTB0i8HZdUZxXKU4cHcevnGGIeDPvD0+CArqx55D0heivzMP69rz
9/4K6yUumZroH9PddAaTXMLt0MmJNsVdnYKwaJ/MAX1QHuO0K3bTIlGRVv8LA8bg
WmqDQzSUr04ZPtZ3sBNwG5ZLAEQ5oJ+KnOPGkYh8lMUgrY2prhWmwlavh+28r/zk
CVy+DAhgrmj1LAYd56w14GaUci4L/y0dcHUYfvJPlAopUXQLmfE0Mhcn0o5oQ/UF
7wZe3ymaAUrDh4bFMCBiaP0w9a3kEgeJ88BCvhLT/LvuDA8vlLhWnzjegQFCfsig
xoedXcwz5AQqPAXRIzLsEap6C93cI/aEUC65XTofeTZHlzp4eD0NP4e38XOpaVJI
Rc1BkX0p6PPFE874h8NfjWmkOqhOFThI9UxFGn+zYO+LN/UNbtsUYemOT4juN/RX
U7P8/kHK9wx4Nd756f+7H7X8aIxUKtjOEVW7GQRZMJPubJLnmCDeTX8i2vVTMHlY
eTxHY/Ul9/lbBlwwZbNfXn/IMQCZwqEEyD9IQA5dnUoQtA3ns7kUJikbVKDK9xR6
vfQESdV8xICT9zq7m0ey7xJ3jdNh3D6hnhdQ7r08ESYOdT04xObstwwGWdLEHVea
0ZlOOm/MuSjh4Rg0RjkeQMSMUrPAAEtykk9IXAQ//+CxToHbehRHUraEirkakvHk
x3MnP89JdCt0XBtzCWg7uMZ+eFlyicuy++tOUa1PXfh1/0daSARcVjcNvxCfgY9j
E5ZkhfwuUJsCsPnejChxEEtC3csVquVCO5z9j2xoGwi1JbRPPNsFB8sDqQaDSbEp
naMOSYuOcL8+KHkkibTPsN0LrZs6x0cYrl82y+GUhgnap8d7+AQUDfiW18Pv6B/m
MNSVgkhf4QLv0LvMI7KFW9QpxXWUYnjwOVrYoahdVF72vFIM+FR7EwPcM4mUDulE
COA1dQgQCcWmcadfdkAUvHmYRwJHX/h0o1NRYVGV3sNQCsVTooxNhsISo6sm85Jb
p0hDHBDBc8L2w5DDDwhkNaTNoP3q8wKs67lz9fJmpQOxfOrdkW4nTtDQI/es2rDS
EEIfVMZTyqVF+rE5eiTFI1F0j7prJ6doHUjOa4Gs3gPuDy4MiXkTsRJXF+kc38xA
K6FQwBqmcaZAUZxAsONbK7Wqv3alKFVx2muH1GM4I93KnfiIjC2XA3WzN4qWK+kC
NWr4qtQrtF41/94YDvT9Q4zdhhqmJIhPYeq6f/VbCniYfW9OISWCmosxPoW4Seo6
+9/emkJMg7hVAe1Cu07vnR6HwWhMeDLpFc98bU0sGknUTDYrZu6tBZPETbWJ1AwO
1BBT8KNfeYIYq4nOZBiRDsRt2cn4euWkqCG6TQd0+QLo22uJDifJ59icJVZn2ofx
xa4BV506x+htbOqLRIPA0YOiHKReqY+nxi4REb0260FVWRIwk3L5MUSGMJRMCrNt
EbbWsg5rX1HpaElkyre7d8mJO1OgzMCyCc5LHGiUarfYstVNxUTG8Em+Meb3Al94
j45dtpYu8T4rnqw3Gh3/XjuA226ttDpnJLEzarUfvm2BTjP+nsYxH29EGK5iMF4+
bJnOiBLW2XcU+FGMpUj9ipx5/4Qi2SLNsWriwMkrKtgbQAF7J2slYa9Lzl1S1KqY
+04Vu7t0reDKb+CFx6cGoLeIoA5XLJwO3tZATbyrtCI/NdB0n29DQfM3yWrOcnzl
rF4ZGWYQId9NHlSCAoHWmrwptGKZyxO12zsTOfwcjKHkpYQcvjC4maaZAnn93Fys
8h8NhcN1KheQJfQC8uQUFzTaCN7vAYJj4HydoXted8sDRZppeeVzd0l8728An5y8
fvEeOWz+hqCgMrrgif6vL2o2WEzllLI4RCOTC5lNm1HR4KyeKVMM/XzPLgyL0Yi4
Lh+pFcGlUDu0gWkMG4NQiX5QLHdod9Mg14i2I/LHCQB6rDjgzd7yu+LjtKVGRZaq
N1kXAP0MMSwyud4K7y46Q8Q0jas+KcDDj7Eb+inZjOrrMwVvpyyRGIDSKi/tLGE1
IyyNqmfydMvcXuKiTUuV2RV02R/mXiNXo0W+GSETYBxtbiAImjTS4OlI56rhSjys
hbDKKm+KRagE8cIW8HMNizJ/yjc2ToMDj9HWlB84i8+RgjzMq8YDcHRsplbysaCN
NIbEBhQYr4uZ9aL3v6BHe1WAgLgg5nP85fIeAe3rlZuL/KVidpKQv45a/Cyhp8Wd
xRGZ2yq9LrsgHACcfqOLk9dxWEYyX42mcSZLkkrN5ilZ94SQdmoMU8uMy5L9zxN2
Vseef6dD37qjvEXGxiZhi5kisDLC2vWXyukeYJxnaWD34H3U6s3BXwokGyzPrQ6N
TA6TGUxtdssap7Zfb8Ghkp3xE+bpRyNd2S6w4SAvhkYOO4Bn7i+06qD6GXmajVgd
ujxcNf1UR0khhgdi3Pb4tlo7oMVtifm5GccotBX4Bedc6Rih08BbTb4xWN7RkjKN
GuZLkv7z/hQcvoqVQtOwGzl4xQVKZ2+XnJ+HtF1wXU9j2DPR2aXegrnenqvLfBdf
Td+1WArUCyUONbAcEdmHJj1ximx41tWeVNuc9rT/cZNhjnyZoNIWin4AcX82u5xu
4H/JJ8tPDgs/bLY9RYLsSekR1i6HNTl7v7ox+TNirtRqhWyn8Mox6Y+6EIQ0lpKt
8hfEm2A20GM5VTI6eRfwQ/P6iETBuZDpwRJ/wo3yzrAUBDQZl6YiqzRa6jDzH5Od
XZPKy6bkIWpeyeo3k7UtPIUeHOpWvZqzHKeYSaOFLT7qvEK0EFD/THfenpKXMnG/
8YaXtbZiVeCeo9NpI/9p/avDr+6AbEv3a7i3dMEMoHdGsCQymYOQ1tcua8+VrtyV
MvLn+TcTbEe3AmLB4fUeJZEeD9aIRlwCB6HmNhP8k/fykCQog7aMcFnpq2bk/lNO
8G4ZAnWCy07I2YaC8YxnLn9hVfH9C6beEnVgCCESx45hz77rY+X57ziMwS+FMULP
WzTu8qR+o/lsCnLiBVBT8y5sku8vNmLjzPL4po1irYyss/g8QeUqvZ7VQFhdQtlo
4rDbw3lsswA7p2i1sD2wzNLBx2I+TdwpM6gb1maO6CU6Hy7Xotw2mUzHg98sgeEW
x2iqSzSkXXcFFqJWTdbQAeJP2RcDr8W0QxF8M2Wc0T+hds+D80uuj6jIHl1/yLkH
rMx3k+G9Q1bFvzHNLLeHa50zzZw8jjHr8LUCI46C2a1XOwLFNTMjmxIhpPIOA4Up
4Vu7dKRQQx1dbreCvK/GoV+F/EC7W6p/g6wGlE0j0Vmmj5Sb8e1VggS5wA8ByzSw
Q/7vRQuKBF32YkkEbLg0+d+4oCtqw+CbYUuZw6j6Mqha5Kdq/DkahnMlUz+GPB8E
qmyWJy5yEWIrYjgM81a7hEnqHShsrPpbd1lk1kv4esuwrOAaKme6UYo45tEkjEqP
+A/07CZKIfqmHPwepg6JbrT2ilKY1ULiyZNW+GzAZty9Ig3nMWbhktTAuCevlL2S
maPf+HspTwm8nRj9j2a3M7kWqZqwTyJy4TTWrAyqHUQ5asEVh84EK0bgOEltNDyw
bKLOwObKQ95bsNElZCCfouTBmPtm5qCuurWHjYjy+fZQ9Xe6ehLnzPWs0eCypEGl
vupY2vhZDFZ8r/dkJVKnV7A23jGYvJi1+2SiFSRe8bHk5oaJTr/y+BvJElGKEGVi
Z+GPBquaGqIqROSZZHQih1gfn2mUDoe+X+YkuEDCJwakZLny4Wdk7GEZecYVyNak
7dLJJr9FpZcAReqebOP+ULIr3Sy4DRSeC/ngjQnUueJL8gQmXpaygZfPsP/x9kzJ
Mholv2Fq32NUOc1tQyG+hryZjS4n1QDsqREjJoaHLrDGgLvOeZb5jixXAYa0ZABH
SOE4oVp7rzDwkz+ZVIdNDR1eD+l221F2lGVriE9JrTLr8KDCobKzlxk40oGPHT6m
5nObELxWoFSyCmghVAdTKYEKyGEVxTogr3ncJe2Ef27sfPnhP0EFdwu1GqYNCsxy
35xgsYv+cjKgeCbirr9UpMXGt6gMB54ZqTZbAaqzM2G5BuQVNY5TE42RhpjeIS63
ICXYiUDSQ1oGIqQq2r5IJEDHuEXKmHypdMF+Dmm4cfRhjCciXcsKJU8heRaXytRP
vhUStcV1yL7k8J7KjSeZS1u+3pUKo/7W3AjAtP7Wy7UFDhxDx5xIx2wm5i41HC15
Di7cTza9FwCRSWbmBTOFuGiBu8e9CBlsVtmlc4yWZ6H6bVf9mlUOb3xNt4Cs9n1o
KEakg1FzLdC7/5E11sVfMmM0SfIR6mK+5PJ98L/b+5H+KGKvHHbYodUENJe5zXp1
kDkkkeDjajAF247jdJLnIWV2oDLJl9KWShazts7+1Pv2ysgub5uiQ6m66HIAZCDC
q8YrNVlnk1xLRI74oT0h6/q7fU1/MjgOd6XpKklhJeAo+MuCG2T4igRqyDqXKFzW
wlX/4rHT5fIrwvjMyAh12SDfusfjvty2cu9l2AUbX+XbvhOdyqT3G07HpWMz55gr
SnPlRR7JIbSJkWRXtB899j+gcRM3tXUSivnhObHIRcAvw6lCWFeIxTpQXBtbZpQh
6lthUgXCrJVlaSmWA8ihpEA2c5bRV8RGdpCStHXHlHK6Yd+5VYhzC+D6p1P+bX7b
KfzmuzqW+qS/5lCtSeGshN37AaIrdTkWXGPwUX62nnRLDy6Iq9G1q5Xm+Q9RyAP7
zuPRjUZtNgrkVDr3wOqLbi3/oDZsuRRuWJPJl1hzjjfUf3hq/kKGVBXBqVqrGQ+D
061t9Wl3Cj2vO/M57BbiktcDYdJZMKExljqVV4NU6A7mqi7HXl+ctz2pAbJKsBUz
acUQE/xxwHEk9l+uKh418sk66/X9cmw7M482K9iHe63Aefrta2C1Dc432nzZpwCX
lUlM7ik2KYa9GjtDx0MnHG7mXbf/2HheTXzO0ZZLfD7MD5KRBohdhdbZs7OIlnlI
i50sx73AxBRIu0MYs2a5nSSO3jUnBXZfI1AgbGsX5qwbGOhrrywU9SA6HA0ehYyy
+mfsAerrCYpkiB/NT3kSx49PVfEmL9M8VrEslbLtVsQHo09MxVm8dmeF4kPQbIdT
+UKms+rUAgLLyIrzd14jy2U+oINE49+37Ha1hmLKRwjPfn9ro0ar8DqKyND2Fqgc
jB+Vnka+N1Ryy85BfBqSKeCHnAb5x1RvAkOqA5n6S68FJ9bqxprYgx8rt8Z82FLO
nZUyANs1fhVu2l8YZfFQTcse66XAnKsN7eylmclVT7hbb9VxuY+982sTYnFR+Go4
NE5qiU2beMoPxfqnxp5661MOVwjMnXevHUE6WUTwEIyMIs+SkhSdBFDNpCvE/7Be
VuO+6v1euCi9XfdmY5ae3mrKLmCCXLVhLXmhkQDDQSlyq+TYYYzyKSPn9D67Z43e
g8f06pomARe1kPPmE9s3EJwaezUNwHF3dLWMfUkeZOX4fM79tDuRxOMaVP8fo5QD
hKT8+NNaqpKN6giwd9ZLUT55Q3uHnVwF8jk+UAAo1Hkwe5Q9slggfQKfWckLOEIW
qbHDTzgIpjiyxOUh9slw+Z3q8UQ97r0jae0sT669DyvBPxNumNxW0oRjmyzGKmuB
lG1W2gM756hSODCHn03T4iLUyQ4tzqb7fESl+/UdeqNoWtni6QWeP56gjagkZU9E
2nHUdf8AiQzS5HfUv4I4yZbBTqu/2FgAdPsrxQB+dB1v1XgGsRAtS6aikjV1ET3T
fGAElFHF5KBAe+Fx/V1QmVU53KoZzX/+C/M63tX1Y+THeitYX+tUoxMGxBkGa3T8
LqpueAaLP4tYh/CcIrpa+vluVPhxWP3V5fS1ZvySF9CbXQWHW5ZcfJNkK+NrOzBV
fKji3aa9SpamPrBkTqd5ts4/VDtrdfqha+MTXv+w2XQsrUDbM+tnNjkSDFzHP2Uu
L/0MM+tSTBJ7okKsotrpD2YZd8U60c5ri76vkus+dwy+SEqVxm+eOHVJ0H9uiEwH
olcuCeMkejm9DYkaV0VgMHYa3odImt8cimpNFxtJAQ3+m/j57kTHAEP23SXcMROK
T+QTgTxtkew6w0lNEXpaFJm2OnCTH2FTSBEhJj2q3pGFjclXDK6REmwpyNVJSa6w
mM0MOmx7ahF0DgP8+rU5nC55rMxv4XQXVBpivMRyQcshKnQ8TwJgsilWlUfTxAMu
F+gbKUZJeo0MieY6yOO7mEQljgXCe0q8BhsLf8gKDDfAeaxvN4Xz/ZWzYP0qRjWv
MU17HdZAhFEMoRwttmPhtVoXUhT3wvdIz20NOhfDScYt4J40QgcZypfmpb9ilEyN
KKklr8Fi1X8uSYjxfhBhLqbuiVEKAtAuCu0hBeQSToyD1n8INQHRhN2WegzSkB/N
lfUGDBotIfz9B40uIEy9tUr6JW1hKjU449rcUyiTNcUCPvzvby/TtvQ3hyx8LRWO
O14Qz6xBdG8ckk7zUFWbTNVIMHyHVWIeGGIXVkfTClMBuvnwgm3E3WwjC2KPO50S
T5UXDcKGWOqck9qxi0++SBEYpAZz7XV0KsOcvWjT7IrvcTFRNmSy3OKLLZeNhSy2
13a1OcQo0Ch8njaX+ZsZaOorJUML6UnIRVHkdhNLgMq8Mhc7nH/TweHMGqMDiSHn
evHBGBPgzb1QUbjWO2YNMYjT1T11zX603bmF6m0S5YQyLHdIttdVBlquiiQs0MVz
n7LwZZJ/BYW0M156AeuPb3b7putjOqVyI3RA/PfEltppwbZDygqCu0FZMF5Ar4vn
dDKQzFSpp32TVjY2+kDUEwsRivMv1f0fxOOovMcbgOXZzQUbxp3nMAQo0lXJ3lmt
5wqSTsxP5373W6gZC3na6DPkG23RDvyy6y2a/HfgXlLdC8DKIwBq5AIB6sp7PcKR
WEeXN2JrP3sGbOOBzldwGAChDh2Om8/HzRx7FY0pi4XaMGlEtuyEGnXHOSxsc/FZ
jLPSZmaJ+YZNpheaDXQ8QyLwgeRzXlht+xn48cizMjAdQmwScADc8NZQycB7zOz1
sxryWiHkS15wx17Q8xfE/tCfzJBC5gxemyuc3AQnuPRMzba7EVxdv8MqyCNrg+SP
K/6t8X0nXxFh5W+UrITrkp9lEtsikzv/ZF2ZKF31+2QypCJ0mQtrRd5v7shU1XAc
wo5nLdz0VFwwKiRHl48eUiOTX8LDpQx4fgPKdBa9OvXfCR/3nCTBn4nppCfrqcCq
xV/GeEbm893ram6k+LNmvGVSPe9Ox/bakSJiRPzsG0GYLmcXoMQFxoilyGWSUJQ5
9ZNKXstrW0Fo2UYaPsF5Z/B3X6HNDj/7nyiJwirk30hLc54c6F48vUqEVLbxNUuA
9sA4atn1ZCrJsPo08KkVdYxN0QI79O7Vwbn4HauxT17sxDtkMyFJoKWZENNcPClv
cLx3CUR5K6ejAFc+aARCncgye/pVLtOqjEgyazj07tB7y/3hH7akWlo43CFo6EzH
FOfJHUZ+FIOMkGydmXoMHV4oKLfCc83l53UPUP7vkId/VB7ebsDtVAznuIOMakZh
BssIREaP0Q9oB5fzdfuFFslR5kp6wGwGG2/HpSCN+VtN1jtlW/m6g5/wM0X9Mfpw
MMXfLOg3bBOXP1g6qtQzf97nTssNSGehOG2RWTFgkYPaxItkF+ynPvie4qP6jLQP
9CxcbpxSTK1y1DG9SoNDuwFMr606wKXIl5dFc2DkbyZKzOjSWB7An7kb8BmR7X/i
/a5uUILFPSwuk3GzZ7r6aqvGtvqV5VK7sJuLN/h+1kRROHa6SQulYq+qC2GJma7C
xVUZQqyX649Aj6Qs8M0BBu2nWnbz7IdxMX3rfu+9UzvR3eClYYHR11gA+R6PAsjL
rKq1CC4nDyBGxaG1WjyIennzamEef/HAt5tgm1slksZhBMhT577f3HdufEiJeLyd
HMzJXxiE5AY0WMo8Ad+D+KD0/rJkwPlJc8srbVPXGpEdhhNbAXFrBIOOlsMXO6G2
CJVWqsk7bPSSELRyXc7S86VffOTMQmk1SilcCcO90B/1kq/DFpkB5lQtck63nRkM
LBKX1kujxyo6LPK1ogu97LtsoOWA57qzDa4GZQZeYPnMqylP7TDfT1mXolOjc5x6
SE6lc89xirgzsbSvnxJipGYKWcRtf1US33T012nd9N3pcMkSdBZKzPSVdZUuTOJM
Zxf84ltHN4tItSf+nH9OE9+hNZBVP2gFr8PT+b3uMewrRZU7T6UTDuH1gxfa+24q
/eUFTOBlzmUOxu1w6oHDlz9GzS1IbWdN7HAJjWzwHBHuXho2pYLeHxgYJzutvaNo
f/2yvW4NyieIqrNa8ljbTkps+wXUijsBqYFa7qUwQyWfXWqOrYkm/ej+Kq4QqqpN
BX87kDbLe/XvYb8ofG3DDQqXqw3llnbRJZfQNr4YzZqPrS1RSITx7nv2eA56fsDz
xLrVSfocZyKiTUC5oYtKv9ouzusWmYkQOTR+SLRVy1cozqTLzt7ohCdXLo/7cWN0
`pragma protect end_protected
