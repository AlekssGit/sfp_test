`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
Sa/Ib1QnmZ1+dFoMCzReiJ7ltprGcX1WzU6EetNr6Cd9ufBM9SWBcks/CG9hiQKV
qbfxzY3k0Tqb0QWy54FCQqkMAcLmgDQAXq8AXMMtZxlimKN900xYPJZrcT/uXUAG
jxGeO2/K2REAmU9WXaln0jLnBkjZP0SH36JvUMgmD48=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2022880), data_block
knWWIsu8ILdDdKFbUAmV8ak2C/1qJlbFKCkeh5cuM6dsF08yy57B0lM6iN86Vhtj
VLSPFnIw/yidUc+TxOXdPxB4pGsE896ujeI8lPAiLZFrTRL/kU8CgoCzr6aJbeYX
lk6WIHogVrJ07U9OSYdIN6m2HaiWwKjpB6PZtLZt837vtQ/Sw86vkKqRYxRzop+W
P/ykUC2T3+XedL/sHbAPZ3IPUCNh4LQzXH0ZKAQ3+vn5ARI5xG2Y/LzgmuGuAElq
YhNyOfUWI0i/xaATQBTdDbOnlhJbMtT7ByS30bx7ox3EDtrR7GgMqpmwx8BW8ecG
xhgYd74hJfJStrU2OM4XN0x6IjbTh+y9FFYgz6rK1zaR9Ep8p3UKzsBAkOMATYHt
pg5e0SQxX+CnjKIww62Eg2gzkCR0RHvXuZlB368n1CXi+eNUcf7WzhpjRvZgZBBT
aLzBh+zXdyfRKPacPSaMoGe4OzHFdb0MzmmflUP4GLq0aj+90eQeXFASmDW0OlIy
90JeKOm6x0oOd07VHkJeUNXcKFLew9bYrhz/tGhOPc1vpBMHi0UNg3H6hcIsQoz1
3LtR8OUX29oTUI9RUvDyVWrGORG5j+41UYLOajT8yrdc/QUtszjB/0f5FObgl/xW
KTDh8gxAOk7yMVq+1/wQoXj81qdekW4/ftsMrbX35Gexk46xPZX4xejaYR53QyZY
SCJECO6/vzDDFx82W9UeEcLyl626hYb060QWziPUv5H3b7cZ0XwEjRUU9E6aIcFT
Pb6bmb0MO/f3u8/Es28p4uwtX+dwxRU6p7fNyrT9GdnwNc3IQTnlXuKeR7zvCvs4
+bOVFdBhbaPosO816v64NFexeFklCUeFyNQ+NFti0kCEyKkUD0+h/3YIiSUcKi5u
uXkytohuj9eevsdhw8Kn3E8WOKRJwBds9vU4ToiGHsIb29aLDGfTNLDireaX1TV7
JF6MlDGExE8NXCWYbDmTNbjnUna/TgkyIl2DGlbnhfomI749DUXH1/CTUBEPB9Ze
xXlgzEn+eO15Br7C6CSURChAzteX0jMFTq9BOKWSgzkQc56o1o10UwRyLbXWJw94
jT4UgSZ0gOwNkx3ngdc2fRbABnPZc73Rtkt5dtLlbutWNk5GRLrHC2y1LmfdlYb0
o5HYdTTOwoCan3AQoSGkn2/rZb67/hpKU+4jiIX8Ui+EVvMklrb49ZkWhuybEQ7U
t20fQvQaPnDMqj7X8n+72BQUtKhgbhLCS3PB1WO3eEWER3481T/idNHXwo33ACqd
+oRJwNA2AGok+UnHimtcsUZfGtL0mNtK6CCce2DwPqWuh3SDUt78r1igReai8rZb
/joeygJmjUjkRYBygBZpDDRRXKs7l2+OY3RWdVM0GliWA0wKs8KYJM64v54xIMXP
u9mWulFmhg+QAKnX0bb+LjNZyDffyekadxBEfFAJzGhmTq+hYBV6RraGV9LMubrW
a1uYFg7lstnD482oqtHpIwjST2ADGPwOVNBu6KLRXSNsaveIoyEKnZ6NBEJzRsP6
zxK6MipwvuP2prNnYj4XOOZ7s50ylOFQDkyqbImiOmpejIvrnZQ8hvKCmffb+AEZ
7s1UVf6v/YjM/E/zYA4igFv7Z3ZimRxG/zwbodawGXEid4hCGXF0wcXGSnzF+QbI
uytgb8ya7ZLELdmLzz14NgG/+f6BorZ1NDyV4+gnLJhSpdr0RDz7Xw+wtIJn9zo2
RNG9lUi4ccx78cH7+xZxjPhxitpZse6cMA6GRFyW6F+Ok8iZAjX2PAqlcQR/z5nK
t5sjo//7E9fbM1ykg5JdC48X8WVggTGTsGT2rjQ2aoD4gCJiFE3YUSfEP5vphg9B
cjAzFVpmOKkQCryzEXV3RxawWHxLnMR+jGzbwDVo0ZqEqu6YzZo/jYJM+LjDzvdE
o/hKIR5G9RzbB1kK1bkpbp2WqjlM6F6vA7ieeBENszZdMJj4z4TVP1Ep/bV4yY29
4k3cmXhds9xuOoI2JQF8KEd2ZuJ0919aYI6FuzHTpFDhp3BF9MqwgHtnccBl3EHp
/uGeu6rsp8QRdjBwHW3EfkiqBBMNsJrh+Yify52CBeifQrqZFx8oDfxePbrvQzMp
pM+AsJtL7T8ZCnPGPShD6pHxJxm5ZWBoZNpxtn3kX9AypLoywLl/k5Pxd6NuWv1j
3tdFriCaSJnO60NYp0OkMSVg3SfezmQF8+lM3htDvkwEpDABsMaQLOG3nGHWXFFx
ZKzaFLJytMOPqeFQ2njeUBy9PCIkfVwBlnJKVhr6QV+ScsRRRZb0DsIokzgvERLR
AA3q2d6+cGEDLyPQvxK2iwPpRXmwl0z1+2smxyxDKz2Dpx+oIeVU0+s0le1ppZvg
fsvuzwfM8Jk8/CU9bD1rc3f3ZoPhN1QHTMMNHQOGL4SBf2UDdhgbxRhE9Z3olhF7
V5z55ipRItSEt1yGEGB2fQZx6c9EDlkQOex4MAM1m9EL6N3AVlBPgRkOX7rFCFFw
Be0QuRidJYN7zETBYtEUtcZZ8YCcAj6AbTJ9TUMZLWfc7XjojlKMxI8fyRAIZAhV
nS8sDTdXB7DqairiT+zFtXKaBFqAs4PdKTtZNQG4BDoRXsO35H6q6/HJNKGNQAx8
pKi/x+r7ugPhsW07gt0I0YBot+nElYD13Cb2iIIuRLfjO5EGRgGc8U77mMNrYSEu
f4EUghdD9cUEFF22jKegTaNJGe3OQPUf3nA96yaBGGMiQKfSDlR4lIq1InS8IKxo
NHDsLvTntgwqBCkyTulVGPFEF5qTgmEtVRyvteUioIskwWjpbAHxT+RljNZtWAqH
Omn0KPhkg+kD983SGelGxaIX/vaJl7qy5SjMSV7MBi3/XnsfZTdsOGVCEOTyJxVg
FDasETGmHGtmw5pq7OrdVtZJtrgPqbrDeR+9wbWCKEUMwLj5wWHO/HA995PqAix8
Znb8wfLz+r00wFmllsbNKSGe2pdOEUJHf0amMpdwy00qI8v37YD9hywEFOfsNcco
0p4bWcqLebKzdNNGdsa8Fd2bw450i0Kuu7ug6KAjdPfbezZj2Ud6JRZ9PPPlCCLl
cyzkt14o2gb8n3SWxN8i91IU3rogQhcVxODIVi7STeyGBhAmqfmRqJyw8zdgupk7
bkyRCBd3AHsVjtPWf/wi1seyAUyd9g4n2bOuxQLdP7jIyrfI64hA6ejfkLBLcEIO
ehJouB+sVgj1YDHM3y3m8x2gM6umeN1ydjaBrCG/udD1n5dLTrmHJH7DE/Foobji
shvGKx+lcYma2wIv+LiqWeDyAoE9uPK+bv6ujDz63wtO4I5pth7idXKgkrszLYH/
UHZsDdP2QAiPztDwlQAcpwRCkWAKC3heUGGuTrQKA9l1igmcseh609t6ulaNquMl
/dIBc2tgC+Mq5mNjHn6asZMs68T465kqzbdRcA1SoA2+lzApGPhwF1nKeWK7lI+f
0JCRo0K5gZM3TH+mAiFKiw6iE9bpMiWdh/vk4azaI/dv3FsZFjQBVlzuuTbp7z2a
2F7NpUqG+n+9kB5yvNEQ2YXxyGSdnRQS1MzALBhRSAuHNN1fEM7rgf29VI4ZhAzR
H1J+9EdUgXVXrVxo6dCO7LnR8rjbJg6HyPfRPPiOBk7bcehf38Lx3deQ5b2ISeRA
R5YfIV2timuQYHwEC1Xf5rXdr8Hiw/Id+zr4GD4YpZdQrTsdeUecXmCe5flMJeI/
2N1ABmQQGrvIb83VQX8PfKMW3dqQ6WQfTMjGGFMDCy5X3Zxio27IbPWW+oWcRV+g
1N2wvl7nNzu1qDYUS/V/TP91mXP7Fc9xn99TIyG15Qzy6mn+V2F0hy2CNzJErW6a
d7CiduK9rsIbugt0OGhAEQLvb9dnAjff5iFFfgzhthg6P+bjbck0H+WXCxgEjXET
jdB2FLn7Ln/YyNiUHJLZUDWcyZ3KRrd0Z+W5L4D5eRr4+qWWUhAjz6ite7BEOtW8
OWYx9B7bC13006icncBEdM6DDAogu2c6WRsh6VaOkdTg0Xcs7OHtFgWHc/Bqgo3e
h8pR0k7G/oDNjJtDhWRn9DRm/9QZWKZVBKaRo2Lv5O4/Jateon9cidkzRN9A+QBy
s2mannx/XF6JlQF0WLeLhzv9pPZfeS/IVCNR89ERn8b5BA0EYoYwh696VvEp8Oop
ihyLEZuxdW0WSjhx/XSnmUBthVI3mgiTa0h01tENZ0E4E+Hpt4TnI1arH96ii0GP
BtN7lxpC4q28WE9hACTTd/1HiUwhyxo5iMg4XaaaM2y5FTahIULnvdOZ/K9NNm/v
xZL/BdKmx4D5fnqrOQqrBpOIfg50nP0MVVjcYxDmETMI8FJhwMp9gtj9k6OVw6et
TYhwjogmTsxadildGF4mj1zBAWRFduiUbnWu3k2D19hyw9z121kJLN4yUKgj5Fwh
jcbARbQDOCw0iJ2YJ49DTGrzY1L/gtIhctnyuLX8tcWoUnUIMGWnwy5HbYul5EuD
6CyARiyibTLoPh/kr70ioG6pSY+xakbUL0u3wWOigaqfgbl5RKbOcIC83sY9yZ8v
0WfFjllQxC9bqheDll9larhSYkvPQCNlY3gtH+wusmRhAfX4UMmpESudq2EUEx0L
gmmYQ11gjK8jwHypGgfTJISqmJLI80+4GlbmV5E6B+FHsBHzWTCqanfVGVvqLhqh
sVyZTuDuVtMeUFLsNnS/FiRgoIxeAoAE1Pp2GC+P8yuDFqp2/cy6J7jZCTmBKSDa
PSKWRvwStM6DSE/IYY0+nAmlFdQs9p6cKK0eY0LQetkgv0OX60dmxyl+4jNHHRT0
E2T9qAAbsYaRwlwS9OL0rdFdwcsy6r/L2qxVJl4V9c9E+1CeZlUlPY+570eexhye
9RSXw/yzBprFEhIIPPCJMjIa38+hXdW1+dMGD8Ij38Mh3MpIkQWnGFLH6LiBL72f
yuqEqQ3TpEuTyPsqnrc1wX/CYcw0BESCMrusfuUJim44tZ8AtyU0rVEvU8A9oGls
2jeBCyEC9GtOQ+XDcKlXdsij7T/86ZTgz8iF4L1b5dg4wsfi1zfT4NXQy3CaF5Z7
j4fwfL8ujWm/8c6JMv61m7qK3Yy1GAxI8Kly4MUcQHCBKrJ9aR0JKcy/NCgTJ9lw
RHOZVeq7gUTwhK/5rEQAFzMmcyktHTJZs9e45E/UJ3YSCnEKkhOWiR0FS5lMgEBi
Uw3MisqmCuhyBDOH4vZggKBEgN7dkKI98j9d79OLmKSHynQ2yIQr8gnHT6vQpPG8
6QyVckglBtElyEnJBf8Qa0uZ/zuhK10YnKs+QhQYEn6kmsqAN2Bc4Bo2aOzI+sxV
pFlG3rpRggOY0IC/j2+cVlHnwISKdNZsxke49PjGrJzhqNgTGfagNWOHkey7cua1
L6HpR1VwFMnFBrYJerGXTRX/UZoBs/10QB6cdovqcs0gsIsqfE8W3S3GvQ674UYx
rOZHEiWhCrhNp+Quw4ATIOEiRjUO642IrLclwNecE9sjmg1PViNCQdu3DHEvjofG
CrWTWAk9r3xn1T705dgPE9PaPnq1UeEEMGgSIACsg6G+utvGSSTVPWhHI/T3YxpU
I75Wy/xHg6xC720dJ0oOgpYM/hj0NfAVyGl/pSTxjyEefTZv01S0Nu6u8/3ck/QH
Bn7fVxckS/xVrH2chooBelf8RcZW1SIpHNf4FQE3mvUY5mItQAhnQbxTvvmXlagF
DYEXi1c7VOrDC8oFoBycnPJlfjTFjWjf7Qi5vwk+byROcKcx60yiP7q1HN4VcyVf
BrEv7gtNyT6+1pk5aH1lJ4iLLUc2Pi+p/gxJvmEiPWw6/RPaYQ5FTqVcDkupAKKe
qEU6p8uHehriIRVpvAib/V57RPgm/Nx3mAPNJ3aw96Z2azyeJzj734+gdZEe04rO
xkT3Sw/uwyz5GAve+la9RX+D1Wk2gnbbP4jd5U25713N6Hx8bmSEp/XA6OzdWh32
ErD9855cwJaYvAc1O0ZxIzYNswb3E6otosnvdo+Z7Tav0fzfi95qPzhOeIXziVK6
5tCJ1+IlZNwd4zt+Cn1zyxqV141K3AUTO8pKQ3SZX8b16l/dhN93QPq0V6ND4Luz
V2xKljqcOa62EIDc4MQAfZlKUMiygECY78JK65tsaLMNvS8Qh+NwzPvMaY0egV/Z
BvDhy8WTdH+68yIjacS92To8RVEVucfxU7n9hN1nq/tBGskmRk8jx05SRGs3qF5G
+cYhaBd2spcSmeKLpeAf/SPtI14GC22ZiyCt3E8Usjhjj4oy2w9DH0z184+QRiQN
lvBWOHeuoU5K2dR1Bbo4HoDPT2B9YQ8H/OOYnWoN9H8Zzuz1+UltlNa7ZVHAVt9T
QGWrY2Zaei9BAUU3O/BBdzHeAoR7ljwUAqo1LgB8Ig9pTeI+nOgB0iySRUYJwp4Q
gkhi8IkQctcyRGeoovwtOW1sMLwzpk92JoPskXVREHKRfb73S3tvQ4AHtXNdA2Pp
tMIj6ZehZoSmGDbxcwrKLcf0h0KXofIvg8Yl/12LY4e7HLhcpo99rTN/kRSvk0S1
Tsvp/rtOa6WpM7Cd7lRSky3HbLqhrZq7Hl8v6lH+Rn8ZoIr1BH8ltI806yUmTvG4
uDmzkmcIuRs3DjkXcEEBFR0GoXjtXQiOAJksm2b+F9sxB5h5vqEzZg7Ic8hn/X44
vd7BSLYTIoFedgw62eXWt8+oFUjngtZLMLs9XQbpsQfwEUhVmC5P1HqCpWPeAvxp
7h9daH1wIu1czzwMEPB/OVTkYywvl+bLoQyb0jiVXScWxzpM+Jvbabwa3W6V+tzx
0UDP8PtE4F4IEmY/pTIWnz4d3c07ePMy29MNPXdp5UxJLglK67vGzNfIeLkPzQ96
Mq2xfcLu3bIJp6TgeOBu3n6VtqhpmuYotLMqK4wQCdtctF8yTS6lHeZnorm0CQ1N
HEUykQwOvV6J1M+WGYcfI0UaBgj3UnnW8yFYsT4p7EqqGxtcUobFapqBEtRzdeDN
LB96tKuyxU7qKFOlGSsHflhztqLL9/OMnSq50FvVrToA5STsBKV1jgzUfHGDv3nT
CBuVw2TWv7rdBilwumzGhaOm7eSKs2knH/TtlRLicaQFdKDW194EPzvMwOXV6Ngt
POrrZ2Ti1idhxk4j4UA203bRDVz+0hmPRtZcZKIlN/fiOd8rDWfK5NKk0Rx2PFnI
ysdDwkaNz5xN3FWvaoICJ6Hx7R6KnDyFD96UeZgTYIjbkPVESYw1gjAfSXtk3UzW
x/49R9mLEVLR7fBpznlSRFLe9pQg/0sKCQVULG65+Jy5GIxz7y4ptLykwo0h+wZ6
xqpUzdgAZP0zcy+TS9tLNGP4JxuB3zt4W/6fWTsXt+u30ka3xM6eo08snCFF67Br
eEp8r3lPArXYLpc1dv1GM4lIgSpD6gTNeHzFJYR28N32Bs0hv61uxKo3kHvmdTXy
xONbdFxMTXIYnnhxc5iRnS6TTc8jwgwUGhyTT5xiHQRACvMNBafp0ZKUEs6givCG
k8CTXY3GdTPvdLAL5ywH21ZCY+/EbD7lzav2rAVuvaOZUV6IyGjn4KrFd+rbmJcw
y4f1aU8BDOBRneNYhrFjNMXIRiuADdbR4cfL7DmSgd7sJQVweCv8IiT4HZvTyXyu
mcJ0KZn33125OSYEJZO02v8ahYNZpNhLByP000fgZrVp8mIm5SZpAh0G2TtVr16F
mXjSQVvfqHjLQuyFXksXPAhIZFEc+keuzS92t9PnAhTWHNraqqHAI9GQXPNxoB45
JRV8MeZnMneCaozaQ6jVvoVuesD1qfhXS+vVPXt8iyrQlfwmK8itb3qz0jnBY3L5
OwAocfqH1Uv0025DTmdTMOavZEWecCVLeTSzgHlIj9XRFM+PtaLBrFDhnfMFYSnT
dgoPHamLmXtFyi/lGsu7lBtFaBWO021ZC4QWU342bVqxeHBDFOfJRXNnslAAU1g1
uLXx2xFrtfzRxyWa2ACzZIBpuHVoFuRFfl8P+GmIa87MUrNgW94zo5pRmwFj1EDx
GCLfVS/Pxb49e3RR9/BEi3YVBPMdg3M6hiFr17grqgH81biXJHb1VlBumDxXGoTl
QMaibREHdEnM77kIZOPEsbrvXvO3/sH5Mk803HkzuRkzMSmV2zTlTNg22KVFGEbj
HzaH9gvW1dwxO+NBTFNn0W69TeJJehAY/xXFbyd487f9G06pFkMC5wT5BAfVg/tT
FqO3H+b9b2gP+F8SFh1VIBIuKDsLethtXj4P3/0OBUdAR4QTaeeSvsY4Mb0TfQKA
elSPA0PIC9OI5tGnGh+fj+vaR6YcADA60axOOyDlcnoE117JjpPDEqcsG7jmzrBO
36tOBQ+/RnxXSp68bfvdgrOQe2p/U9WFcMzWKABoxS5eEzBfIOHGpwndeNo/TCA7
42nosVhT9ZdkYKlGU2wqEKgwzF5x14DlPXj+wTaVFxnRnE5h7qGX7zs56UMqMhsg
NefPMBs4X6uNDfyEypqWXJ/3+qUjeDwZMjukrW1j5FwsX/r2XACIUw/9IjRIh2Yt
O5TkVtmiOXCrZvWl2sBA4ydy1nHgtOqxQnu/mr71sdFY6pZiUYSTwH1VJicWHvpN
i34TuQ+qqS2AAsQJroPZtn3OFpzDKuJOu6TNeaFtqTlF6m1l6qRiX2IzVo8D8sy3
zBj6luAhz1Rbhtv7lEVo3kRSvllG+DAuMMWfZW1byHnICQOmeMe/xLFwr+ddMDyD
bxAKtC4ovOh4PNGsx5J/0ZLGIWIt10M2GYUTqGIWvrIOkvvREKMd+Vv3+mBicjpA
YUO3nIScsGTx9JS4nHLhw6cGhHw1KeMIX1wOk0w+e6m3+zpz8iBk5wkolNJ4wxyW
u515eOZ/58u63eCBQFUxpTa0Bv9eyEt+iRPmDPdCyb/Z3/n0rj/PAF18IQcwV6lw
bmKNiI892OJxt25xZr822eK8yU7+L8OpnlCWD32eSUOzHlvpdBk4rn6klClCzXqm
g6/ZRZIvdwYIe8gvJO+OyiQr0AN+ilZ/yu0XhHjQHjrMm/TBT4D+GgjRk8DdQiOx
u+16qZleJwku+LrRm/WB+AV3De15+Fjlg2/PBlwWJfgTA67TCdMiT4N9gi5cTaFD
m8qQPsofU810ecQHCxOgw9SfPy5xEz97dyVnSAv9xIe6lrmEJJHCg64kxIIsyz9Q
j40zRMfQyyDNCoQDQPM5JknodClm+uh0IjVV8jr6mohLijQRVm+apzZ5FyH6IZVa
+CgPkjlutEaltNUGS51Qx0sZK0BjXIAKpaI8oZdrghggf/tiWQDqXhLayJ6cBdvW
uVlro+y3gNK+7tkIPsG5JRsxioDx3mksOOPeqnELo5TUtq5Dyg4uguBgtWdNVMm4
Uprk/gcb2C99qYiNTa2XCR4UeZ44v9s0ad0pK9wslNzQX/9gyttGDApn03Jrlco6
48NKhtkEVXeSYhnLnBYVpGu+bGlnVOTvN4HDBWGr2CSL93tu5mTZlQdRwlzlT1JC
gQGM/S86SHy9XOZItgud1e00iOiIRXxnP+Dtg+nROeRR6qlAzXa0NzafQ14pSnAw
dy3fwPrSLChKDy4EBdQuaMXiN/m3e/hl4pVaWQJP8CtcZeMQqiNL2k6tW1E06aRz
m5oSQh5f5wBT3koOo2E0cy9UztsjJC83Lb3s+3m0beNRLzTjRt6oycjSxp3Rw9vK
WNMvWmdUwAk44NdwqbyDa2HzSyWWSh2O9lHuZtbh3oo/IpI4UF0jemF/0RFT4iGf
c1yDVbVMByCwSkFjx65qf4Kz6S9ZNMoEPfIeF3nV4KL++JowhBeanAYtoZBRy4sh
u2vqfPWb4j1x1Y1JjzUQnqkETFKWWENUazoT1wZC2lEFfGlLGQKrSvYX/65dNe5d
pPgafvUrZOrFCBCJtRCi8+1ivhj0KwscPV62jf/1LuG4YAiC1nwWYMBlAurpTgGA
2BXKRBR9X3MXxVy7rehdbm9pe6UagSA93IKP8FR4ODNpeNTCS6kCo0Y2hftsG52s
G4/lwCkea2o9+Yo3PjTsk9gg/zL2keY3XtzJmYEokBAuf4tCxmNQTxBoZ5+AH3IB
jQUh8WVuzoI1dfDIQ2eo3xwmOWinCO9Zjp58YJ4o/yx793eilqA5eu1ZDdmtUrkm
gnQEdQD2buDmFwnrw+F/jP+67y+hqFo/Th758KpBP7BmusySMLcGsdUNMpGsB1Y6
WFVOnYKuk/U4F28ieGGub0rizp7AHFXRe7Q4LJWDneHgEKlJ4RJNQffkO+HA7CEp
W35CjPSzTiI79XXAEP/a8xmON313RAr30IqnKnc5osxZaqJTjjFqFYkx71V+8Hjt
U95uaa7XyCMFn+hy1k7zwXgPAplAKfOEDByfIYXsj+psnbKFTWvAp4KZ+Bk2zWUh
EctHqkjkzw+vS4q1fcVkCPZKmqONf3pwg6peUSyZZD76CToZdHeFcUrEB6QKhqhy
GLbWFP+pWIF//Erh/40URF2yNmnPuDClNB6DQKvbY9eR4phXTohUqfDuP0MS/KK8
BuUz3BLMhbq8SA104OTgznbxkLXMsHIaB6ERIASJUFXw/Fk2sAYRBky5Tdw8kYIG
XWVr6NwfqPn3ltlF/IKg9MGTsKvwolzjRUg4V0V24QrEG3QiRru1RSVropDvJB6U
OTubaOB320tEocyOFXnbYo65Aezf0CnPnNOVZCMPiq45oqiLF91DScJx5a9uccy6
cp1gZSYjYCu8zYlXGmzGPsQP5UWiJR7zhLsp5vwqk9zICcAOofNKa216/0yoG/2h
LSqwK7jvmN13yI6PAQTmrOLPA4ynlRp7FDeGGTC703JW//Mw1IYWVWClZXjeBLzI
i/5k80xIwTg/7um4f92v8SxbCZTxe+QActMWoBVdPQ9HOboo8CuwlsDZ29E07R/o
TG1LtFObpJSLoXjw1rwh8jZu/rr4VjZYF3yuka/92DpUc+0dqpIq5Q37ps7Kytgg
Dz4ZYX8sftDWo1Z3hl1wcsxmlQlbyGZKsRnIFi8Kg48Kv40AmWc7BQ6shtF46tqa
CCrcsvCQNRtouiELlZNuCgHiT3RjpI2YUkeTAofa8OtSqG1GgQDnzBUd6fQ0BxgZ
P/bZdhxxDwQR8eIXRAF/cRXJFenTUkdYd0r/8Pq4FXjY3YYzbpHE0d2XiZT6GA6S
EiypH1pMSAuAtqsw6LtReeFOfWy3mA/TBK8pS4CFY1evqPnds09xCckcHmxzdQPN
Y8brz97w48h5CeWreqA88Q0IYPBEgvLA7M0dI3SY6Wu0th1dBq9ICvs6fNxAALu9
D1muYfckRWxh9XiHPr5iqVCVFHPwLmUNnVOYhgIPZ+mJWRht++U1+zKiyYV0ai/a
WDlRyAE52Be3VaUOVjFv+7Ls53c/JXYls6K5sYQKcP7j8xLhrRHPUMyGC1p7az6T
Clv3u1N7BLT3EuPhO5yNDlqqVL6xciSLk/MR3iOZyyw75TfK1waW8cq4SVGXXHal
0+AezASQyfneUb4YbKHsERLIwKUySAr5svnBZY/EYcFyCOPsKS2zPbpSm+jOLRIC
oAaRs4CFcYFTHbNmBSzY1My9wNl5mHGZJI8Mab2UjP5vKZc9DoU6/K+yzFLEJcdi
/dNtve4LMMoXfSxZTqwk5u9mo27a9e7Lnj7QPdFKf5rLxFNjqbea1eO+ivCV4RUK
NEnVfZ5C55GGAuFDgI34bNYSfZwt01azyIAeDy/g2/SQYfqJNg3cLrYmQhBWa6C0
EOb3AGEReevg9dvSEiASeul6dSHuZUpH2oXPGTGk9w0uiW1o28DTGEa2Ydcz3xRI
jfXWRXqSSBDWPc1hpmYnR1G8VUhoTzlQ3FhMHjbyd4Q2JxpoxlFx5tRujDLlHef3
MF3Xh69VM/S8hFXOywr64kUv5xyznbDdTM6RJnADqsT9dhlFLg6iDxvQm7DPE5rE
sY0iAlsqPB3mG5gl5Vnn66/Nx9NFuqS9dwHAeDC5tCahsL7QYCvcQv6lp69sWzaw
nSbMDFN/3SJ2nQ/s175O9CzYP14t0ovN3oT+k52opRHV1rgPmhaReLucUzF2IfhU
5KYDuC6AXwCQlJWSwYYB8ZwzddmRtNxL+tdw1GHVKJhs1aBICCko2FF29ftuvyDz
EnxiGylfvasO6SkrYdz2YBcoorMjXZhtmcW8RqH98tzEyzNkkZ97/eRLUJxsUqXp
YHxW/Hl1LZWUUFhGLWtzFQpjCJi3kQ9ysKPpcapqrtwh+5rmnOkjnWlSHjH9guhp
0K4H4JgqoQeNga/2CbPt9TLSO01E/BXjxOIRivrv+gu4cKjNK3wNTxEegmzdUkUD
y6DhZlGDwtFi32WVV/52P1jzxj9VEp8anRCRGsJOEykoYXdAC7zUo51m8tPXuLpC
2CCc9I+Wd60OLPwJ8pVyuCpiT1tTa7j7Y813b5+QHzkQ5nUgYIsBNWUrlMov8T5t
s81IOV4v7kJwKrYWd5lYrSoe5hM2qqe8C8ylf5PiQgP8rqSneP/m/Sy5zbIlj/3M
HiyDZYTSny2FXA7yge9uMPoHNCGvADca4SxadSFS3Cc3akeQEFtkAh7ylZ+w/wpS
p9SSxYQgPDbw+Ki9oujJUaWNmg3Ke5NQAUjhYhiJdbOb8aFlVlAqW6fJbWZi3+k3
e2UC14Gb0FDMbUrUf/PK0wkBbC+csRbLShg8efB6WDSD2pMMvLn5WbUnqPhmH/v5
JeK5HlV77pLbyb0TawwarbemiF6EAnZ3MDcE1nU445AzUtin7iIhRTWy68+YpoVk
/3VDRQiRp1P6Upom804xVL/iPx7ADHkNi2Gqejh4B1+kt20iEGB4bdu00wSCRWuq
0xv97sLF5rJqh1Gp4WMTnj1getxATCtmyC13th1KcAe5ojYjv8FXECL+yDQjxXx3
hrgrQU3+tOTVTwyKm2LvTSBG9K4BFQ1Ej+3KpAqcPj0NWJx/Sn8wK6p45fgT03DY
1wmZtx8IDaQmrHnzdqoGwGsXzvV37ku0hqUetLy0e+IWnKnMoQ090xeMX1t3r2/O
S1xybCs3Iof62NprwluUkaZYNoU4mNwM7BahCZszYzvtJs53qViwS5PiMTcbB+LG
tfaWTw2F9kjscrCAXlWPEkrKcrLxb7TO7q2p/ylKGN4URDiu9LHmwMCu8KQaVK67
bH/Hh5cjifrEEZWZSgTD7IlCEb0wtT4ndMGCTBQCYihvHlJsI2ulC3EB2hYs6ans
hnTI9I8HGGiuKUe0Ly0oTsKY0uNlT8M2lxrb6DrnC8vfpsNIDlHCU6qnMIq/xEi7
RfF4wPr/WtUsUSDvjpaVAS/sWroj3oRjDg7nKyuxS2h7305/w78D+mT5oj90RMER
/tzIQpmrFmR/s6M83qsLnGaYJM907CS9nLJ/1qoi0VGXVQwGBE/oRSUsUQfBCgo8
1Mof5l5nJ218vx8B3bUyASR6F9pUdWYpT3jDyG9Vn9EvnRBl9nYmepcEeAcVOIdi
lNulmHqmkXeatuuuQ9XV+/fz3beuGAjO7KMoNnCTfMBXDl8HF2hMOWo6HV0We+nG
GD/XI1K/pBTTgpuNyzCr3KY8kote/9JAxyBvVrLYXDRAcFSlZ4gBbVXtkkimKbuK
DZT3VeYOxOpoNU4fBwut/wLBN/MAShIJsjwU2UjHn9TGYS4IUNmv3//DgxXIfmwc
SxvwFJU8gKxVQs9WUKaq4QK20oNjjpsQnlhXnvrAlFoxDfLobMp595PKFow1fyBx
SmU3wDWG1LKPQyEWmFNLU5cYypWqtIgLBPykfBIKeYjoxbFd5GoMc9MiHXbsnfzo
QqoTDKIM4mSxVWWnQakOH2oiSAmEfnY8qjXxB1VaJVVNwe76c2x306HFbgjHGMdp
HVnbtkvgmklvolV6qUPgOwfa0oT3vzLFaGPLCOq6cWra45bO07bGAxH1tZaYdAPL
QZBCLsgZNlJW/JmXcAEvFIbjjaUTwj9tbnC8vAvnKcrK/6+SHZ2+qdkYo8/Ek7dX
wc+PjspZAqqwHtscNUnDufeo7KsqDFm7yG2F+FyBxsbGjABZE4gp/dloLQVB+6jr
ERbnGn0/lNsJjMVEoKs65EfSkgxQQF89iujPck7LCuIl7HCOWS5j3KBRCyCsMB7r
TnJWKYclrs3GQdu5/a00k9iw6uvrx07krz6NSsBJbsz2i2S06gZgZsc7Qd58TZH8
SC1kTfvllmAndgvxSAVdy0r/ZEQYd0WQho4YpXUSFAOxQlgp9glugtn3YvwG7w+E
i2TMARMVP537SMZLUKFvZTsebQ7tOlupstKs/AEsbHpjq66kQJticW/iODuQMthu
R/8sUg0aBWqFhpFb9cXkZXX8dL+XG2LcQSeh69FKfQQLwdoXnVHeGmfbSYIhkdJ7
K7k+UfdRtH9dGgPgxfuTbCNQGu2WF7ASRNOD1pGqpu+Z9t5fHCo4g7UadkKKActt
NdXcNBtKr6GJrfUAXBZsf9iYug6gDwLjKLGmANz4MfL8yabm+pUgj9g1gLmtELOu
XH6UygWRH8d6Ub6dnn0ZPNWTHEdhVMJlG1Ac0jjkn2s4GJQJso8bl7QRK/XJbaQE
yznzj75VahsjNz+v8anQ5UgMFmL3ifrpNv4G88BS4RRr969N/FoXpoQkVY81jgmI
mx+s8Z8c3Su0/QN5UXJol8l2EH0LLwB/jLLZQzjrkk1nX9vKZ9bOsWz/U1+hQ4Po
ExJsyTDE+MQIqRrk6toHNbtVq3bAlVsoz4NhiEpbe/eK6VKwkftjO/l6d9qQ6YnU
fqFtxzsd3GELsWHHj33m3/TlSmNVCcEo+HmHZNrepXsIjK3KB6a3WJFa4hYB6Yp0
HN1p2yhzYHO+OrS0TgDg4EpsfJyCILoXWBtGfembh/Mt92FLbY85Ocu/Al8KTRm+
DqfFDwEFh/N30pt77TmdnG4oyIWJ/waOF2HxB6GMQNVQOms93O+ko1teRBZYDel3
GGXb2ssTJ9Of6gYaWItk+Z5Fxz0wDV5LhaF6lsVk7OawEwO54VoLxTDY5l896F6y
vFUPBEef7t6NJEaO0hPJxBBfrjRwWrEuWeP6jG0lSpeS/sldMTwmiVMxTeQI9+uB
wyw9kFcS2ymhDcDO9T3DEk7eGnezvBkJQ4jhhHDboVHh/Rdl0cHXgke+9hK0BlEV
5SsdFr1Gdy33y0cZsBRfiitSHGndlM47GYoMK11svWYCyqkypE3/DYIQSj/4Q6U+
79M1ofi72Bg/607QADD+ZvXBrY1OwpTMnP0sc3OSDQ67BqVGtlDmYh7alzlkrG2y
z7uEz181VUSXNLeC3gZsFSFiVOqfuefMcj9/WAv1gu6S9JNSXQeH4JmL6hKFo4N9
bETOr+ye96RKf/4oj2GWpN0mbBN/bNlQ+aLhEEy5AB93mUfE8C3ugQBFdhhP6W4R
tY7E5P6/YrCWxzbaoA6bJKh+k1vc3lhAtGjKUCpAngv4kHlYLgutjlH3bOW8oWcw
WqFU3QZdedizHbrjVUqC5LF+4bhL/LApG7moNnpJ9yN7o1hcybb3VYj6P/wPtxyq
E0ah3aqXE+bJcKavGac7t0dDpHwRaRAlCRIMdhpK6CfZqlObO16hLEtF/c7zbday
LX5OnXg4gg/fwobBojT6ryFdi3ip2f3UJDPRXL4qPJvGLuFAUgu2qb11v+xwzD6s
V6fgErC2vEXY9JWuKfeORRG7E2WQM4ypX2+16HH2MN9IcONcLA1XDGqnaHGcS+1l
ICu2tRKj3xK7CrNvwArMfgdM3vIMQY0Lox1ef/bjq/k7LmX3AR+CeJFJcqR/K4k1
9SBV3rlu2sxvq4YmQ7XdWdi7U7l9Dv8aZlVYrcd1ld/hBAQ4muh3Q154DTV5DcRJ
H4UGtmZN4d5yiBAJcHZnMnawxYaS7FLudvxDW+YRExYFWHx/VO8gPWD4dkOSFyU1
WOorR6fGpDl6Y9LRLrjKvtaftLAQevlJaVpvoblY9XgZGEfknh5Ba8vqwu3TDztd
0Ujffa8AChFPAM42uB647t0Beg9KgID5QpzJaR9uqi6FhZyqiQ9eRCyexlhhPSNN
uK1FoetjAWC0MMvf5eUssEmPkf/vQmXxV1xNmU7SDO8v39yz4VqwAznZvH1Dnmi+
Ei/30R+Znc04PdEM9DfcVV/Ro/p1tMwDmgZoaq1PsHS5IKJF4yteN0qdou1RrzLJ
5vmHfHNMlsjS3M59otgWnhVyDALb7RWC2CBj+6gMXO7SgRGY4L3edtshET85F1Be
T+RAV6iBxtPUIke5eowhrvHM8QNaIfk3UnGEcoLHlJ/DIKlbO3gYviigZU49yMgG
w1bzNyF8SclKjnT6X6uSGWCNevSB4PO1mVO9qOVxKP9vBwyxiugwt8rH4ylQJYnu
jipOWo89CwutdIE861jOlkxO1S/EfghdjyvSBrfkhpa52OmRaWqa+K88aZZkPsF7
y8zyO1Ul+db2zyb9mJe3hWYKpnkX1esWoH2R0ZFD7+UH1nIlM0GPZ2zVvIme0mtF
efi+MKfwMsCs2532xtG2WL6bbwbIkJwj/j0x4KeNgfempx682hxBxHomeKxutPWk
L2SsSwUV9qPFKEHsCv9mtZY9KBavLrgOsiIB/GPcNFoHZZReT7rInbaige95wiUU
3MjMqF16avFDZGqiqGnT+a+1V0kDWK79+0j4A5H0fYeqTRv/tz1M9Tscj29/cmEK
OqP885FtWwOzP6tuQMLYInF/qxkk+Q7xk9qKiqz5ObtdOatGWQmiNXw7EVeuQxI+
sxtdI/m45KucaJrWEPJFV3vbHJawychvY0roPiI40OZBVBLgmqdLFE3RZS5TwDtF
kHqaH44/xJO6TpiMsb6nk1jdYRPq6t4SGTCGq2d8mSlf2CfnV+U6vCJ9y/ZsB+qm
S2zaRVuTsZfxTIKwh3+Uzck5gyW3ABf6470TpNNFC63g+PUrKOfJmrA8r5dnLRr0
2xvczExiJiCP8O/Tzma4VyFbRbdo1+GHHjPjNz6GAc9KUao4Dwm39q6I4P/+clEI
QKcHIQlF7lTfaZS7/YPwEgyojZjjE9lekmc4YAqY42gzZj0D3SgkQsrhirzZtgJA
YWAqJpk7Y1xm7Wv44bsvwJQrJrpgzE3aMHejplAbVXuy/7lHH4vKwvJH22df/r5Q
bnPYcFqB/uFe8HulDlz698iXKV7wFnBkJ6+RN40q4r2sz55acCQtREZXy38lPLiU
W19T3jSQimDvoMR0zdLtjicbjGlcvdYf6LUpd/9rBRh2x+QYLOL8CXFZJlDuwgmJ
j5QKEuLkcgcFbqQkgIUCLWhB8VJVoqm7QNY+ErZ6yeUtvrBJuo9X/2OKvbB8O1xq
g4OhlBw0nMhIzMMpQOe8EyTHEzOWchPARaZllWC/8RfBzaBQPDjxEoUaBF42eVri
PNV/or/7c8CaNFI4FPD0eF5I7gBdBd/V+7wJz9udY8wYfqUIHX2jupUQdXP+gstC
X/RtX7de/1AjZ4xbKcfXchEETXodAmkfSiZUVpU6zXv6TlWEadH/8ksEKjGdXgMf
i7DALtk2zvHE9XZ9/kIxpuBUY5lxvDNPBFy3G0iWll862Y87iij7mJEH7ywbwZDd
dPiF/L1I56L4o9tf3RhqtStGYC+qUYOR+JBIhzagsESzC+AlbvIKAyoMe2yjh9l9
2FtWr3J8AQyy7nvinKpU/qZ9Q2jmh/Pwd1TiVdjeVZ7Ogb3Y+MhaiBGoGayGSc4K
0LxNUOek55q74hd5VLmz9MUBFxfVIqDz4mW/P7YAtUVnWjYM1MDpXdREEHtlneZR
DxFkXhDROkaJpMOVFSch4yDd9FVG9bCGIXc3k0o8aJ2loQgYs3fIHdO5iruDnNXT
+wSclHwZmOlcYNXQ8k27o346JxT5cw3+SGthmAK8su4iQD/rHsrU5Y0uZnyQh2s5
4GU5TsEjRsgugpuMW0oNpb+3x/YRcsaitvJ3amvSRLq1yy3G6SO5kiJaBtmc69Bg
pvT2l4l/9ZTlVZBSnrvv6CUKd30u3HJNKbj3iOeeCWQDAdCEIhcW5hYaT5hPVmHX
cUAtIN4wgd1YrRJkj2ser5LfYuchMJ9USNPF4RtH0PZZUV/hgDxyl1ZWz/lk4EfH
Tnb6GCn+j9uBmZ9nDxR1UsOdEqKl1u0Vp2Lw4vZeo0QWXgb/ba2GxoEwzzTfDtKv
v0pzx8xncEA9n/gRne5k1GjXz8klg/D/kCv95MzmORLp4jUeSWNZdize444rzC32
m+1RiQxa7b8VIS04F66JjdF4s6z+11+pj4VC5KgNC3SE6Qk7J9yGAGAhUbmKU2Ap
RnE3X4pcQOMebPZ/pL5ZFAHO85VKr/yqK14lLa+9p8yR9rPJttDnqhiu2VbrImHu
yoxl1JVYQ7HAcckEx0SOKmCFQ0ivJAeG2MlfByu+/sGSL4bt9iRC6vMr4KFW7ksj
HhLGIG+6BbNZRpx4YyTlqq/OTc8UClAAFXIc79Wyc+bINpkBmAR68bj/i3Unkn0R
qR/j7ekRVK9TV3YEqMUm9hFuDPlZ2CRFeu5w/pMnRUXHM3SsC18K1RpddisxzpHc
wxnX6Sf5i7Q8YfZvHpjKQTPoz8z/RxhOAPvWP/SDOnfDYUGc8xe7RDj1ux6aN/sY
vSnFb09Ly3MPA4PFL0E9Y+aRjotaFlVSybLvfTgIpgxGyDquwgOGkRiXmj5jeCY1
RMkI6Mh2FW1T7yeP10BSA+cUWV9DAbjPWDpylSDaOD1Xe3dONuHcy/VOybBpYCGH
810sAaBPmCX9VuloyIoLSmjgfQONRh3XHLN6qExtd/ihehklNWFMhVRAM4WzRJeq
jMtE2I4rPRHIeRLvP3nbVGc+m1Hu09/TeiR68DCHShFeoCg074DwJSd2Vtpkk7ds
y+nVyRTpI93KqoC09mf5XVeMqHpxVdB8ayT/lLZB2GtahU0k07tfRfmAKyAaTkDS
06L3eMeuNrZ3KsONnTXhO1Jb8MiBdP9LJZHIANmSf1vVYGEAWsFjMJDP0V5vjK8Q
6Sur43RFXb8+BdthuYd1CCVCF+yT1aJ20LQtvO53qbzP2n8kiuQpOe5bag5079Wz
SkGQx+eaUEX3OCs2hk6gM8e9cgypMzlSe8l4Wc0GULNSEaVHXR8uwJiFFrXpw11v
aOiFtciBRtZuXnauKbN9Qp4pRP87hEV5ljP4asIU3uWj6rnApJKSYIWdEzVRnjsv
B8AypfP2S50LnrtlMMmYWy+ZC1D0mUfm8IdU65+DnEyQfsKhE/+/cJAV0XpugBS5
UKr7UZXdeU+hEA3YxXCANCbSk8mCYso9MnGQoX7BQpUjZvMhMnBJJHvITm4R6fHn
oq/BX+eQf5Gijavn0VDJNuQrravAX+4tDlMG0zndsqs8t8uMlLPkMPTvhChFaPUZ
pUmvQcRKJxdT1wY1az4XJFloRbBKPW0VTJToVgKvqeE0LkfHhY1CKsJmZYv4KXWl
DuM+nMr5uCeEUKURdN7NFJzU1bMklE9/dIHtT9H6EAGHnIlUkujzFSrqFEsSMh4K
/5ua+hZOO7rRVMcwwobCegu/QlqiQdErUqM7mZJ6gOqdVGLc6pbDt2pDcRd8X1gG
uFOE19SbZ6ydY1aZqB9gFUYaQpdPQSiivQryoxEkVlZv+B0QrAJ5/JmbVSphs+cT
NkLby0Z0PecBah55gPUePbBKwArvjH4j1xjeGrFWxPa/cx/S+0hgNkFGyEi+PlZT
mxV7XbkkQTR0kBKmjKLoCqEX6LGE265DX1I7WkbaGW2+dj8sp0Q+OowWvTQ4ZsgL
4yYWgYgUOtC28xmfoYWGNMtWWHln3RDtSDNqMP3GbeUi0E4Q2Wqv+dcF1Hh7g7A6
zpPRj+DE12BzPvi/IFJmDUKjtkzMEiDX+3H8BFBNYzCEpiMWBR5Vt24urOT3edmm
mHTutBUaByQsKGmzX9+uMOGCVdMxoqZUaATobmY7nNAL3Q7n1UD4cPFcj8+pKuQA
ouaNGu18QJ46fA1p/kjrnaifx/04uReYVRiCNYhwUoBZ78aMkVuOACo8WZIBTuTy
kwkmf1K/gXeCU3r+LN+elfaHD4uJX3oYSUHfuqZqlKs3prDaH45GNHZGpGBj7lIg
h5Z9MXLun5ae8bk0hMldpLaEZTzJ5F0gcPZYBQBKx3B30hYaNPPeVtkJRIVo79gg
5j3OGeO4YYG1QlIIL4kEb/9coqF6zzjpCFNWesQG0RbAzelOGbHka5CRzRUIUos5
+HOliJoLbjoWJWlUHoDm+YnNyurJY06Je0oBFg6em7HTTFgoPpyUJM9RTh+cu7sj
xl2G0p594/pqxXPb3kpjtqQkRwLYL9qvqOPkvjWNEWkqdUJ2V3xusVtw41vJyEYp
1ejOm14w1e2LbRjIlWVmPlBBV6W9TX4mfYodYu8jJWALW20Z7blUDH9g1euyXSwo
LwffpSY/v0gM0SGapfS1F8gy0Zy5c1TGiikobvBvxwcYlykMYIejtc9NbSHyYcCL
pyu7rBMDR5bdLbCibqGbRQGV9XSFMZh2nXZr2kLPp3W1iIY1gH8at2YqfznEPJaK
cvoJ+xdibHWdh2AXPqbzAvjQ6BC5T0tSmy8M1SHGPnEgDr6gJinAzxMzkNAgJZWh
28EqQ7G2fi5k9Knj9qGm8itCsoCknYrY7tkl+SnSrdpwcIc40cyRNZe7d1YS6bHT
CYl8hnBM56eTrxzs0ccyEG9pBRCA8XCoYA9vAP0cfI+GtNivMHeIl4vcacrZEVMz
9oW00B+lI5reL3NoQmZznOddOGzH64IuO7bsYdwCN75o6LqSWOguRbRrs0Q5KHN4
2bB3eJ8KT648o2OvRO2UHswLBXkaWRD5ptJCFf6ChvktBmNIzoeuxKI6fvEbRCmQ
Z3QEyOUhhBPKLkUJU6TWvNRNHrYaGgo2YRl951124CcN+n5aycidGIbM7m2ltCvE
0B++ODHAldjwzhDtJ4YT7OX82DkTphIhCVjHTyUSu7idOROa6BNOSKiyYXmXXZ5o
I7y0XnszxM+clswwoml3bQs2n07bJqyxzoNyR9m3bNwUhKs+YDt0PwL9q7Qkfv44
HSbfIGD25DbwRJDGtelHEDIZGBhDB+Lp78aZ+1k/dod6dA2+6Va58CgT83DocMnI
6KIArbxD3V/49JXK7rfityVYRAYAogQDb7WwgJwRAvek1UC5mZZc7TlU7gfT2M3f
K3BZ6pRgzsgHWB2IO1dRqy+YRkYjj/hNCIXM0KDsk5Izt9B2ao7UykYbQsDzhgI7
hGrPjNR0v2LMGZRu9u6xSqlZhePEUBHg6gxqTpOsZ3n5bZ867HTVy1eZgs9XcsYR
XERHq/hG5RS7n2e3cC31micKUIPLofuReB2w/tTR/fkOHUL4cEaFKsTOsqDZG7vw
Y6k8x8UTt6dRoQ4KlHDiTaP200MrfMbZ+3Dgf4EuT0oj2hOxXwmWtLEyoTDhE98c
tuFbA9oR7hOEyVPWa4orX30mT6I8dAoAqKTKx9UR4UAbiLFpA2Bz4ljzGCRVnGLS
Xznb5Pje9li/u1jK005oaKleKKjoS8OrVwCeYFXzRHJs8OK01MweJJIAzVy/HQHY
7T5Y/XYN4RjLuTZKXGbQHxn9IUyV3mOW+SUl2j2ONvvqP+qXRGuABqSG8ttTW2qE
ok/v/ypYlcWHSJi7PMSBve3W2ZeQ9YfprTauGWz2Q4iNCBkHNAncbGROJjwZCiZS
swKvAUvjzdrUeuZNrxlYVI48+ub+uytmxXIvZPYs6Sux9tfadL2a2hAN0Xy+QE79
L0d2sq65F5j56xvVvTgDY4CVrpghb7CI77dAb3kSImicU0W/mfPV/Qth0vmJhgu4
BblQ0zdpnwDVvGFQj7VHu706HpOf8iYi4d8+TXyZq97d+b6LiRG5fr8dkuXqpMfE
XkEwFBWNr7TMmlv6pKtUR2D+HUERdfNCiKRq1+CSz2m8XFp7x3YmOZo40y/LEM9E
H1ktafoDxyIUbcAdptzm8X/9l5lD2Qyhi2k+mK0kZIdPd7xiASf6h2I5CrAfTxhs
KmoHcTdbHUJ4T65X2xVo6N6ZXJpZ0uXxpH6X7BOnxHQlMfpTzW51gzj/0DuWXcXh
C7Td0WThq3UgV488zkldeWGFoKHgVgqo43Zz7btvr7bAcOGHWAzZCwCafGmYgCLV
BFGusuzvuqCnuswLZ55Gfrau55cPPsmf2Be/MLK/1l9vJemhfQornW5Avxo+bCJN
K9VdR+BVSkTQO6VjC/nMV9OsESttUt4t4jgWxq0gTzyd4mdCTLfx7XQrGqejEdal
6WScpBW2CQIBEQqm5h3osj85egVM/ny8EvJQV70gmzMypuLtsCh3xjMHnF8Sg6IY
yc5kUZ33O43LhL4lH7k6SebNqZyzNAvNOa1X+EdoV3wUc9Q4CNTla3Aor6LmOiZx
ojc4FEiYqCKP86b55J/8BIXFbgSjThiQW3VxNmSgdcDcyYUOllx/m0wD0EBztycS
hYU2DNgM2VL/ELtoJSJgc+C5cYh7jnWouVy7J0EX1fjUVcpFPcmOFQRUXdZMwD6i
NR9xA63bQdDBvKe6jNjQLggNTQSF984b3ZQtYbNoE7JdiK1jJBnn3LoqbZ8svl+l
10cnu1vA9a/Uqwz6WRWz0/7AELeiI2HhrESNP5g4Mix6GIz9BR3+AXhC3TUoOJiK
DzT+OTXj0nDuXxuLK9wWXUdF131SotmfQ5SLJwhlfhuApm1f2smotrlAR+C/WUWG
07RkwOY4dVfx/Hs7/cIIafZ6F7jgBi9RqGSXY7wyhJWj/r8Xk5G0+uuCst9yltLH
dBydZijHCTPl1eE3IQSIxD/fCSuNn0JPbzoeMxK9slwH3sPxA9UvGwFFSQcXj/4B
bY8XaVq3oYY/pMQbKS/Ta+pxymPJOEFbs+IoyYgA98bw6x89OZtlMnNqd7F6RE3T
SAgex++kJSacKiQdVKs1OIZo69sS35BcZA4RYzVO8N7FyVQQiicBgGVLbRtJ/i89
yc15mGI7RARuV4Al+r6j1FgO1BkG1DQoYCwrQ4xghSJkofbcpFqkecMoimRQDDmj
jySHHKXdqD/TLpcgO7RoAFqOcgCcJU7UbAmjjYwJ7jkl4om5hwjzUGQyLImHjScG
BYQQrK8P6BwZSIeT19tIvIhJezfO6tgjnxxRCJGd8fSX+IzE9XtjHukE14vakP3u
1PMJJql5JaVeb7sPEFIYAiaTbjbz7DeqNiPwPkXvjL2JvJTgX1Ljp4TDSZAV5Rix
5C4TbWPeaM7iIO01onWIpMZ+uV47OMD9Uzxcg3h4wPdLUJmD/SGUPnk5RBot5xlQ
W/Q3tJITvFgWqay0Pmya5zlZWnNi1cRDLZFADZV55p1utni03XZHtZ6AohOPEdSE
SG8lQ5M0G/z/wAFeQfXIOWZ2yBW9HFwl0nXiafRr9dsVTe2Xyjr4UZyNJQFCdpH3
fd79Y22dpDTM9xyRdbN9PTKYYcGb3N+euyjqOWph5+CB4iDc7KKnz2mPtdy3/W1j
SLxq0TP87TYIC1Zzi+LqMyCkRytBNHPaRZz1Ir3TdlUmIbGddeOZonSG9Em3n8gN
ATJ3aVhdmgaxQn+6Y8IJi4evaWG3LhWgJ0g5R/ws+equCq55O9lFmZmyHiHsL9Cl
jNTJ0s07z1RT95sC1iOs2Y4YB+KmG8PdXQuw0UT9wNNKNd6E5/0FXXNsZc6DWKHK
9TScvpMufMsTcAN9/eud9NO+9lBbdr/j1Ez/QQ4QjprFUrr3TFU94aNkYURJxZQc
jqEw6gu8tzMHG6yxxAIQKAcmPRPeKv1dOEi/pGWYZXkvx6p9/MNYnXfM+uv1qXvt
Wvh3KZYc2/dhhJ/bMBZAkmKCnULQvH4PpFJ8SM5Sjq+X3bCa/pchDS/ym6rT0vYA
mlqhZjX+iBflLi15ixbsZKX5LTDwdHj8HWrjT+jA+lHsNOF1fMkJiPpkGL7vukUl
aus8MNoMrMCsq0yaP6RCAq7jHwARRdkIIxxAF1UwGusPYoAcmC0flGtP2IrN4Oc3
2eaPejsjq30TUpBKfIaqMq1jtuJFrVUEA+S/y8p2Gc4bIC3p2XIL+jMDT+vMv3mJ
mv1PqKxf3LZsEd6yPEpKKiSDLf9oY726I+iC2Vn2mwxjewCv38Pu18haeIUYdAKS
goEBWBreHRelJEhM4bx25jooawC8OlDcEDU4PNMVvU9Mw8xnUZszmae79KaFLMmO
ZiWX58YZS6csZ39Jp8KRrLJZG346rjcxpNK4Oe7OfsO+UH1JlMM4LQs2T/mBy/Xe
xjCXbvxMh+KTpED1nzVSg8oP8ltWTdMbbExyCf9qGqY1Y5+0uV4gmF9/KjXmlW3B
rexaEkyUhp2C9easvHK/xss3QoPQY8O0g+aze9ovGkt/9nwc9cvw5zMO+tZOooHg
RQWuzYsV7vlVUemxK86dIjlePdtN+kea10u2KD7kQ7Q84rEOP7VkUOvNLiIkE7/v
muB7g39xQtWJZxKjUzM2zmwMieF2qlU6mZnkr+JXQb7ac3fApoGpHT2953sPvSDr
Y+k3IVxnI2wjKllXMLfH/2T9GgYSoiCltpY1i6HI4yFy5AUkmTIZPdL0Fg7OsDNv
OiXQP5GMeyliTCY7e3kkN8Ato/h2eSiiBZaWO0n6v2BBPpc+gFy4VkS4jiViOZTp
v/VQaeepb1wpNc/y9d2++NnGNG/A1ho7BCSMF3HZjRlvwMFZWwzRstNnVSqChP9g
sCcoK9PWYmM84wornoGdBIUBZniqyWYKOXz3I2+7cZrmM2Y1Ik4ox0DNoYlULCzM
YuN6pHTVxuOul4VJTererMEB3M1qqFBKfavtQA2Mu0CeAhK2Kd9k9J2UmmqGoAOt
V5UhnJma3vs8mZq0orect5WOBxqVNaf3TC/vfb0sRNrT31hDYhZmdXuwIScMIRpN
3aTkHTeEiFtTQXRBO8XZFz+lcwhVEk0YQnpUgqoHScvTCQB2SbgmkFG4FqPwBWtP
X29GsnI8iRBiIRaYpDfCzbncokVQc8W2JUPFz6LXSoGLyqAE4YDhNubTyEJKwvkv
LdKeF/nmyWNiRcqcD5CVlgGcHwPZzHhZAk9CybgM0PzJbfn8Z+L8RhYKyxU+OjEe
obdX5IFLlpy2VZLnm+71tBCBXG4qWG8fAYxa+eX4OlJEiwdxs24LncVX751YVGs7
Q/yWioj4pYBAYRWv/Q/IgSR6q1Knv4gLo30DzwcXzw+M1PJ3RVrOjUzVlKxCOehp
VnAQT5VPFgkBOEzGoaQnN7+4ABv42WnnKZ5qFjcy7GS/DREGwf42sIei8dE7GQnw
22n3NjuAHYIQyPQO8zxMyyF+TeeigUdYMQ1VD0n7T1ERmLARCw2ne7WFIUh6/Vji
MtG6eQWi7HRXMkhnHqGO6Lss4KUXgwK2wS7HF6QE3LmaR1bzyWhIVZtt3qvFrzOj
qG6NgJ0mme18lalFmqJ8UYVc+PLx07ND0YXWZ1dCNwGMHRtpeLv4dN3MXSR1HDLn
EkvTWZizBJB6+NqgQrh0G5obbnpOMrGxes6WbAXlbTnB+3KoJOLMUNPVfXytPoMS
ArAhRRT5k00TIfpsRKqFGul0yEFSRhq//e871tsYIrIAvbL+Z17bVEM7j0Bq5c9R
yqNq1AT7fAVJCkK+wqGqD02x8GVwScvsMbvRHhkytdoskKR5iCg/+N/jaFlYLq7A
zm8a53id1gFltqLWptoIABj49RzBp6+GmnBJSqHZ9RAvAWkJzGrABmn/mOfxFR/q
0QoBZ/UblCisuEcZhGOPcCC5P04r/ATgzDulyqDB6C6jqcHceRONvUJjVtKXRuIJ
mSB2BySv+GeYtqSH9uG+jaG4+tRFdKB9EdGF1RCvI0YgVGFkugui8EkRZmyrTh/A
YU2yjuJPlc6u8xodNjojVkMtnqwFP4eQOIsz2n9eCmBPBEgGJmRvDPXjDEA+BWU4
eFTPR3QpYXQ9SRb4tfR5QkZiT5p738wrCgl5/qRsYNsEeTBzKMdO0UiBazF04bHu
HvpSO7zPJgNwujwXP/ViG0BdV9wWdot44QtoEFF/Ioxjd6Zmk45AtLYyccnlf4k+
1qjZTzSWRUKDaJAE+Y1QtFg6+y8WFOpgonm9l59VsiLaQ2YZO3nUDP5vAeDECxqq
r6PunM29nfo7gD4BXCvUrPI3gGUWpg8KoM3mtqT/s5KS+/LLcZvBEfeX5e7ps42h
5bYgM66mBcci4J9zJlUJQ3Ik3tKAd16GmhZvKmoViSUR7erYG9UqI5J0odLOM+2U
v9ZnPNKL/TMhGv2bRUQwBg2XJCvgVUgPupjoAtYOCQcBHieYFtAA6GHwSR2hpwp1
R0H/FbYBnEz/pcoN58WMo/zhRbrq94L1MKhHpRR15/2wLYWsGYym+B7K/WUrfTyv
I8I4CDv8O1WgBBEBo+Uw9TjcQneFOWY0hkIU0MDZd8vuPq/SAHkRFIywAATtWfvC
6XoOjsyR3khAleyP5UxoDldVLUwDTqDgqfph+Clf/Ys7EvOdFkFZdUd4UWETNWtz
RZ2hZbSq8p6prNIeE3SBZeIoUoKb6TGE6gEOO0eCp8PVsydwAR3zLrkyYRCIHBSg
56KCMx2amemI2xdFvvvKQTjDykq7+5Fm/+ArI0/2alqqXzrhPJDBHrIT+5BXzHhN
9PGdxp+120OFP7SI8joJjkor1TBqEhBVuaWAx6KaTJ2xRisx+5HgE0ETBJtINRQ8
MSjqzOPh+2iiW0zIGaJgmDc/rNIh/u820lcRwGmytZhzyz/EpC2jToS99OGYscZh
oDXrk5sNiXGFoCUQ0vp8h4Cwa5whzOUd6HfiOVB2ZuKGZ/ATDQWF/jKTEDekT11b
+ShfQBJA+M6rXz+7GYwZyK3g7MPOTxrVjbICEOmJnQMrTwZSvf34XjQGyNrWDYwi
W9EIIziMHVqaFlfbFRxCtIUWcBlrLO3VhRjWQVYbmcFQPJPmGCHlz8X8QbfyHAtF
KvKu8KJu4gYZZfncr2zHeYQklltFAAxBU89CT5IkJQLidVea1Hp2Dgk5qjo2JU0B
EIryWwTpcKjBtSebQlAfnMLxVvoDkOVyDQGJ1/4JGe/YJW/kC+2yq45WBqJo589x
p0qbTBiu78xPNtlCr2/iqTaQCXwwod47WgaKF/eV2eB8aOB1DthiBCHXI/uHkIcL
5u9vD9Zjy7V5L/H49247aUzdXQ/liridcFe0/tfiCJXkvm+iswj2aaCMXxsqQnDc
+O5ZhOxb6GdR1zFayxo+1ZAzxNW5AgXDqg+Fe+NoqcoS3sxjMPZTlUw0D/Y61zm/
iPQfweplE7YfoE3esDhMFnrkkcZSOW8Sxm+8Up1iqtVvKYL7fJCsy1drblhtORM2
Q32jFuFgPAsXaH2QNySjF9h9KsMfdRy9ggQanb5WFQ9PdBm5w3E0dByiuI1a3cdj
k7EtiePUZ13diUoPPAQz36QAwOwLwfUnLpRM5yiiWaQM/5zsAlDmUv+Ye4B7KHRR
bnBTthCTE+WU704fIv6EcWSpIzXNpNgf+FPmTYwEUEj+W/EagJpgb8hobonGT4g7
aigjFgQFv72cajv7vLJGGYl2M/0cDRhDIOhiKkC8KjC6MZksQrt1SgCHDJN0fWhi
zdAW8ZTwcFGCUsx5rluaZqpwqLu8HkJ6wY6aAXDjQEiH+lrlsbAtdY9nf6hO9lBz
4Ppiq3pOPvv+ViKG9O5bMOmSKszXOX+oPow8WdcPB33ZvTVW+VROvZgPgVBI1+AK
L0R4assq3QKXuiPqbq8Jwmaa0J+QZNxhciqPXL51cNXUPniFaeCFn5FQkpzwQSwA
YejiitaQ6aPH64KirlUrleNpNebQKSt5zc5EV38sMqkhZMr8GDC9MuS5/Qu8auYB
FjXoo2XuzOPPMNb+3OdRe7lNVEr/ri+E/fQxxbQtNl/Pqfzgxqde2imTTJYf2vKp
YDg1L546Dcc0afWT588Aq8vSiohzTfLsfk8r5VpUsjwafAAc8yQ2QAZLWWALMnn7
JYiq7ZzPQYv7P2NMY21/Y18hqAZkKxBUvbKHnnJRUBBYO0p5YqDEukdaVL8BUWiO
s7B8l6oYJYVawcguhWuH1g9OZhC0iMWjp+D75ge90O+GbV7wZKczNtVGPGmxWp7k
W4/7PgLSt2E5obtRWDAOxuPA49a/hwnAkC4Vxm0vZ15fe1GYZg2n86L2c/x1nsCO
PcjYf03R8iX3xH2G3zLDdp+0ZdsBiRR/4F08SAxyfW5SbcWRoLlQDORzpnv0DkBG
sKLrivpuf64x+8tLPOZ3VSXt7DV/vLwCJmj8G45mAuFcTvP2/lYoIheYU/FvCDLE
mLcYCR3oQB8E0f16j6LgGuacSFZS0WBR40cl3o1V53k3i6+K+cxu5JkOAzaalN75
fY7Jy8SPz3PYKIzpByMbOtV04fbTAXpxHUNZ5ONABirN45rM9HqRE+AhPZeJdRie
qld7gdxo+gs3WwajERMOGb8XVawGc55YqUfgbiJnMBawSicGh8jfgGwWb97bG1kJ
SmYw12BjTMzf6vkU1nTvpYKBQZPz0GfYky8gOMmOSvW3GtVwaLUJWpOIiybH1APS
Fv7XuTGLRuZDcngk+pn1TNHhW46RgBafnlgVN/kIBEun2kAGplP2dbeWYVT+ffBM
0C6nUaIG1N5+DMtTCYflxbTQ3sXKoV0d89jOEG+xjolD9mnmeXHqNi5ELtqoTdOD
6113tZw44Y1tFCpXVVK8lsyc8efggER8P2nHRQt9g1xfL6/qKDjtwhg/ihjbUWR9
pyZCVzJhoQnJU1yFtAuAgMlfKu8zV/QzGU4GdlF5roFd7xI6vCMt10U0djj3FRbh
fvL+WnbekQfHIZJke68DPRjqTWeZ8Qhx3ZlugwE3Ylbp53MrlUqroB5kA6iSt7Lx
Pyv3QzBFw26Y5TFHT39h0Pug8AiDFxL2pL/rkT7lzywkQ/0IzcM5r4uNtzPC5gcZ
5Ik3bqkcXsZ37biIv1ln/p7SikQ4NEsImX5+vE3vJKTlgeqEKWkMHn2fBHHxNbTd
01pBNqznv9iSzftefZRojellt2/EcC81fXJnN5PRuH8hCjlSExOlCqwvitq87DlJ
VeT9KYFtZRbwBt/U3WyHRcRzTgPPz6+1rkbvJPCZlw5ALTgoDoVydNiU7S5weePQ
8H7oVyyi8x+ib8lPimcU2mf79B7lvtxU0jFPAfE+35hN6R5mrs9+3krt8ckt64a3
NXinji06kE1dCIAD5hyZMFhzcUkWdHcvgnYaVzWiGUgu2I5s2cf2MTuFpyBzOony
FDeXxt4MiAGSXnip+ZpwEFIAnTsJ8tYSLQfM4SyhX06Uk53niVUDRm/WB4cZH3aB
E2etAk9LpUdqmayJbEBINit2L2j1OhQ2raJ5Cx/dTqfNBgLfiwdJFoJh96oJ2sux
e4iWndCimM/R5xRXmWsuym8LMdDKzw7h6A0E8FxnYJCdrv9ybQ+8ERruXs8VwYZ8
Ud0jeEEAaCeZVVMH0hsxePFEMm5/NankDFABYXMpFquMqv2rWrqOfD6RDiDuBIre
QDX0HGbZXU82nGKaauvXs5739ypo2QQn6vqJ0xtxCxAKwVKD2CkMrHkjG486sRMN
EgS5ElzOFJ36I3boHWgurvWy7OdGivp/4Sbx6Jg2qdO0DdOVJYGI91EAqPF0dC9k
b3pOqXnh9meENTnW7+1MJ4xo2Zel2K8VsM8JXVPlF4iU9yCpqNzXmXJB2/yP4ZJ3
TO19SdDbEBt+OFwnoWMNTNZM8P5YhWwigA5ELxg+POvd+WTredpfS/kapYXN3gp6
w4lTRQd2mhGSK3mNT471E08hJ7Y9Z1tMwiECYxziRWIVZQI/NYjMxkHydR/51b40
uX5jEOwRaxlkxjbggCJiVs3q4e8IURmeFQo/uekoOkv5SR0I7WdSttwHhw/s6x4S
Z4QJDJ5I0VOh3rGL07h0GEmjUcFbGB/JacEY2dam9Sq8237ZqujAYTdTyUMXSMfM
hfaI5IF6vFHR9V5kR2LemcA/wk15jAo1hcnuP2A9BJbB6zCdgrw+DMQ9uRqFUPP3
uqrkkE12IzmU1IiPIO19gOdaFlHb1L/E2MFq42b+ta2RJNeViwDZtdBYeWUuBdi0
qgeinzxxMkqO/Et9IW4+SRzHiXE5ao+ywIganBO9EinMc6qdUbTLK3amqJjX7DS0
Y/xS76H9ceTcaFIRVw8IGPOfZypEFZUJBNbj+LriwpP7J2kPV2iWbYwa7BV5Pq21
NThWhX2FtqTygXUmB5Y00pe5bl7m5jobPo5j03Yj/xlApLc6TWY2NksUsfgtdofu
iGjQLM+nZQjWjft/pYeIRmH4ofszroh6mJMwwoxzK2WyaUpA8uPgQLCNcTqF9Qxt
DCQ0R/Dx1IaoOGphasbl07TXXicWI5jVzOI/u0jInYXRCe7UvFLl3O4juYxtWjG1
rIVrACZuL2zN4FahcAuWXbu3aN02LzA4bZnIeDo7Fj/JXfkCxciU3HFcfAt/Q3yY
2AaZJnx0gDJxQMOQFWCKxL1wM/Bn4E+3s3hedcgKDZJva7RRXznIcQm/EYGJ2GT+
4PAU1FHO0uody0p8SZ6GNq0YrptpFeoFPEYxNChfdw92QSQP+bdaQ8m3q0ABkDm/
7CvU1nWodvzUcmlx6pOLIHEmcqjeOHkWU/gF5h1/gZhYfjZrEOeQy4+1WTxNkCWQ
tWl8gZtwTm7imEAEnLAeAHeD706caKOIxai2KozoujYgR81niUCCgx11I3pc09HZ
PvsFee3SSDSt7RyPfZHUx12ceBXfmQBjosFD/dElAGGOb1Fw6F/oX33hD8chzgSX
aVZlycISO+eSEF0I3K+AeFS+Gtk7mkGPGrCktAUsNSTvDfgI9fu2aEZz4/e2ooqZ
TqKIpQtSSjn7I/m8+LyzC+vfjJKb2S91y+wCNp/ujWBn6GaKtl2VZlWpZWoU+WTd
naAt8Wie6eMHzGfv/RwH4jxEQ5d2Eo41CijPZxbQpWxIE/tVX/wd0vUbqYpADdik
N9KK0JyHdrTACTlKI/ifCrQtUGL4+ocu/SUuj9g9j5V5oJe1r8kBoeRVcAbZ7oTM
wJGVP5FS/Iw++jBXvxMtF9f0dOwI15LZgEWM0UlTynuSKeVYqrZKBMDpeS5U/7hk
6Qo7ToN7t7wBr84CnNXf9W1PW1KIC7RkvhAjG7MTW9RoPZmb6vdbYN5DTMIS3i/g
LOLs4TzLHYELUPpYsT6N4tDGce/zv6sgQAHkDxfEkOXYjhyvVUuFx8DOjR+3iI7r
+ZEgeDRDBqVUZiRl3Xi4GnibQI14yHS+jBXViJYVirDpEs4cOG44ElIS8q30QBhq
vQrp2vIRu7DFgsie85rPd7s3nW5UbF11rYtaO0w5JPnpVeKxwIEwCXXYLzdG3ie5
Un7K+IypSLaZfJz06wQAZQE18nEC05V9tEbAs+MGlOX8e/gKsiZ5F0xGXVBYJHXl
qlWIjLW2rf5Xe0NOXMW2nSUFuAhZtNp1qXul778JB8gmkbGYmRfb0Q47f2uvvbeV
DWroDRJJh9fjNeDFa+YguLhdWnPVdbuTEeI7n7Ak+lscB/VlaVQBQ1bKckzcXRV4
Q9IACwDkDuX/bi64UXuxBSx5oYHjqKoqE8JI94CpyHRkXGfDZg80YnRdaRilATGM
50E6+enp8oAv5DSjgpvDgvmKMt8CUW6O59DZfpEIWjgNfsLqyzliznZK+gpFiTgD
mSei8DDK/ItcqlzuqyoYZQ/7aSuFe/xJXO2NFHpY8VJAxFQHwNGMT6HZIGIcAnEl
DQ3nY6kKWv6LZcsVUa5MvbJ7cyAG9uvkVX+pB/ONzxYjJw+bF/mIoSCtOI7Rg3Hv
RR281YcDiAOAB3R9oGH7j/CzBeFH3KHw4Tv8DZYY5O0V8QKovWME1U5FNcTdu6NK
JXXpwlI2/KQrgS5OMsivYRk5ZoEdZQZu1Ztdjx1TcfO8OTlECwM1gbdFd41jhfG2
jkevA+N6FgyCWxv44FfR54Vt7JXOHqJKjCjXov0XDpZqa4QWCB0kyLghds++DjTj
T6xcFm3IqF+aE1/hDlIUvWkItnILjY24yDCIXCEBOihYkIkKjQzNXMaYPYzs7d7d
bPUImoqv01rzB68PLnTlqioe0/Fr6lpyGzVTeGIeIwzTLzRkBgwHI7xSoMQBe004
71harf80XWipcANY+19CqdlQxIupTNUgzaUWt2DnT6qNmWQMSkKn7fRAV9ktZI9+
PUHnmMMXVIEujxBl73ImdK5fxDbGybYvLgy1zMyLXysGZwZRnRb7bsqWm6mNzeI6
dtBtt1EohL7vpAReV7wiCveRYGC8BsOm6QBitQ1qOLu6SRoSb4HzaYbC7gMJtU5P
bJJWRpaT0bhkvSRTcWVA5UgllYKfenYNdd32+lCbihjICzFEaAaHIcoLEmRSQ8bA
hru+fQM753wmh7qzU7XRTfJyoMe6bXJm37l2o7No2cEP81Lok7REYQ1MeSKjV7sI
v+g7zFc97w0f7giwPAM/5ZAJlJtE0Npc+/rm5Ta79Ngbq0ZwaZYzhE1p8y2op/Mc
dR+mkyr75Ga80B/7vngzwaB5mFgcmxj9+CaXGVM4axCb/pkSEeb+PIzmzi7JAanO
Sk3m3hp6c4jwQ8qZV3hJLXPw+LbTO4ttT74DHutptTwtu2E/TgEil8RUiMVPP7N9
6bwx3zTG6gOSLoc6Tf0E+7FDumy+TdN+6J8UAUU5LlTFmceoGlzZqXB//tc0rmbK
tCHkym7hzDeVbLSstUYBRz5tVtcNeBd7/9J97vfaEn5s76Mkrpx9tv3Cj63vBEnm
kGQIyAlaYmQbevtD9mbZU3MeTEutMwxD/3hYf0OYsI5TBQ0RDqiC/TIsU1oJOZf6
ZvLLSW7eX8v77uT3GJZfYcnou63ek44B9uoYS04RoddIC9iu+GdlH1b3P/HWoO8C
fnQhwESB7c2sg90DpqIAKHGbjU+kkuIOWELWtxpebxTgXe6Zko1IBYA98cueS7CU
eGsIoTmkJzZOxEIOYv+B7quf3JGVi9FC+uaznq/HI2rgt8HUKUETv3RcoY3KeDVL
e+AnttjvRVLtKNwY2olEQtC8QqheEtbImNYFxqfz+rxsiwu3ekUydjOjy6BhVtFS
Ldfnlu9D9NSa/AS4d0M3EA4iCgGQA4rKrId7sqZNmQgmRFORc30CJEVRuW6ZoTQG
YhVR42BTgNyAse9peXb69yjR2/7t90/NpwiAeHXXlGk8iSAlC98O8NBzgrUjeAyJ
pKtEnoCaC27+Ib9iv5vPy1jw9eSBGsreQNXsLSYVQOIiAfbIcOR4ufRQ16FeAEJX
g1XOnMvp78h++DlQMVdrimwHNrHbKvrKw34s2Oihwh+61a0uRjiD8RrJkBO6l31U
NlADWcGp3phCIjixRE4gMfh2Acz9NE/ufsxJFuvC/TMWqr4ML86aM1/i1g/KfS9y
+gP408jGhxP4vvZKTxSENuS6rXlqCpfdIgpLLgmiuSxqWBLOB2kBBaol1SQ9xHHn
lr37ORtyB6Fvnt40lrRQxIxRa/Ahu9/JWIKGPyG8qsfz5fvG7QVXwTFIn0N/MJXR
/L5azQCEHdviY087LDovXM4bf5J32qh5pPsGJXfZ7gqD0wZ6o29nOKLda62qunjr
ZNqZGtRVbiq5czRw0ZNqeVyf5nqD8ffvt8HAOpRtmFsmGDFv1nhnXI2ZytFSz3Fe
N9D/rMlbUxFSI3xjVENFtPZGL0VXpOXb+ZBd6xpBDC7aA2FnX+L4zxVJgrhM9wPm
A/+ACL6nZjEGi+GEAyFKPwS6KkuVb1krYv9bT4lPFG2xXrslR/wN428dpUQU9Yd+
1WE7jNvgAXUTtN/ljdGU7d6K/8/YzzRgBJhrsvvC5HPvZw/9wT2JMJ72kLXBn9W5
BZt2of4ZP3xwqK9upE7O5Y7Bo0TnB0Sc0i7ZJ6AcMa3WsXCLBLa/ZhMD8BtjB9i5
MAA61mJhNCk2nX3cUxDstHkOylF/TAKPYwOcpt69S8bsdPr4euKOPUN43qkLAfr6
WgCIM+eCCZBHa+vcOkxPf17CbAC8cw4Z/9V+TxKzO8eVO33nEwC+tuPeNXqgUmAT
53UWQhsPvT+dLzWzf7+YyApRviRuHGSK671yGbXSi7E3tA9xf0KITMMRbpu6n8yN
Plt+7x7wEd6xK7ebWRr7ak9uYondJDWFe0scSZdkLFP+WJDy9eF93KRM+Jyr/b+W
Ev9/sdT7b7G4mbLpKERMScKgrFsl4lQpDS+qotg04QovASjPU7tB6QnngQBFJzcl
RpCx/f8kgEMO5dPE1e1Tq2AOxxs8Rf4kvlgF8jqqU/HNJz8Bmz88j8Gwn9pOtGnI
0nSir/iOzSZT0QHXJVX0qn1aosBv/KM+LjsMr+db0H2UKe+w3js9dBlV9oY225Fe
eqTblZLRdVWg9kMGwcMEbSnTvqScze08PdBnoRQ9k4CiOAis/jPx1uKbPoDfbkB3
GH5/CQG4ev4uTbSGLPmwGBn7QCwuSFDSsr7Mtiud9a2Ulf++dUnJCW57GtkCGJAr
xdfdiO6R1gxKXjxovKanDpdeM/txfWN7xtkIMotrt3xJqNGNFP5+EwsR93CeZSPv
EKAe+mwQjXc0mE2Ow8Zay2sJZ/CiiRKxtmkTSo++/mupXLAbzdbh/nzC9FJdsYiu
P7amvq69gRJ73P8WfJ2i5SCCuXLHfkGEU0X3EqWqeMc4qV0Yhr89pSX1KXatSyat
YwnfixQKkAlG63M8kHVG7hPI6KjFN1IxmIia1DVW9mQzQluFHK1axy65PuUXyy3R
GA+8QtSazAKLtWUkPcB/azvLyK0X0Sv5MRKyNGVX2EXpYY61HY7/+yBhp/M4yepF
1DgHZKBfvYMsfG2hQTdvkI8JN/3tMSRYbk9UyOBZQTMnuuGy+J8iEXNJi7KlULwm
VBTAHZXQQNQXzS63EEQtzyYbUbSSEt+BA7xftJoM1RYn0Ydlp2e4aHeix4B3K1DJ
MBz5Y2mszMqfFWdHEGsT7ITduyGsy6hDlDCSIp4dIr3SSDVjtMQlUWCv4BraKyTC
J2ZCwWREPwUFOn5/AW/IWBLuqcOInyNjNfksHuUlX+MwvpISAHI+88EmMCAzgDjc
O9rTDQxPe0aaHIKhJ/rQEcCQNMMoMBTEdWY1OFrTW8q2KMOOXrdX5ozPGwJmolQu
B3WFuK58+O4nAMh/V+LjhjL903Xz+LAdZfgt1J22eXiYkRswmoELQNmAKfbzeBXQ
iAss9dL2AHhSEmlZ9zpqwoSDcQCoGvnVKOOKErrs9tOAums1tDamrcRG6hvq/mjy
SvNWIt4T4kRfCRyfFE488J4wgdk0NZojkr8XN2E7DefwqWWOiuKyKbvFxWle8rnQ
2XJ3JnV69l31T6JhHtf/81mNmpRNGOI+DKxq3k+7G+ISRQPTb2Y5WV8LCf88N1xk
Eipu0dIoE8NY1fWV1mvWpQOBjzf84Yka+s45DmgwuMTpY5TcH8NWRtpI3hhD/yzW
FMrg4ngk2as0kVMNBnzmIY5KwNxUuw5qiJIi8HQkF08gk6Z9Ag4rAoQ4G6Q85eKV
Ra6fFGlpRMxRe7b6eQnXAhrQbEC+OoljWe9PquvfnvdBqW+mDouKTGkwoBE7/yc5
Gm/trmGeQhPtpNjnvBSLe/XOWofXjPBdm6hLyugC+p+5Yv0C+oWQQeu6z5wUKAiL
L+FWvfWnFCQ9kvJ6cKt+W5zGxurZYu+sj1cmxFs6W2tDtE6E40zCxjhluUIqurPI
xvJ6uTAMVd5FPpW9MNcIZA02K+PlIkS29Cr1xOwZmpYA5FZnrfCoEy8cyyuayPjA
+ej8cIDsgXxWR4cHC2ALA1z55ciTuP7zT9yzhRsrE+sja7xDpRIkls3FXh7DDU8c
jm50MHzhBSZp6Siy0Hn71IJ/vJy2TOJHY1YV8B8cFkmukVvIOcDACFuifMxIaN73
+IFDXzVeNZcp/NgzB+zm90oB1hq7V8jxj6r8nT2okGnQ826LDL4+v8hcaRQTSRlh
yqvMaA7yJhccrBqGTu4Is3cgDov3abIum+CTnwC4jzGeUZg2gxbkt2tkv7u5hXNQ
8sD82OUjai9wVhD7f8rNieNC3ASFZ1dxpCWeOFqbKoPg5JXLrQ6utiFOnIZImJgu
sFltuuozKTRoKElstRKdysVw4D8nnnGp2LQcSrS8sMAvMBakVC/FKTjeIHHLEQgd
1QPE2cssdUMCt0tTISFjujTqvE8QvQJJ747jrYtkLqd0yYD4pyhrCrY/Ty4PmP7d
M4iHuTW0IL+k8EgAPRva+s26md2s5ywxTvqByOxgWDteEw1hqYigfebp7cLbgZ2d
TiFev47qjJuY5KcxVsyrKbUerYp3P/sqdU5/Cab6tPKmtemjBJLyVc2zS5Lq8+nl
TLZN6M4EbS4vVDMsUDcmSBKRgylWTx50jNyAmsbCj1WG4fP4uVwC/cb3o9stv9xL
Z1L4gUcQQaorqUap15akmxUalhEAnhxS9UyrgsvyXxzRtRfolK8f0e7QDOnaqOKP
6bw0emcOJWfDjH9Exd3RZCIZXAWUllyBPZQtX5S89Mr/HCHClF8KPfoYX9AxmrGW
vkUY1axNKlKZiW0MtRU316+/qagBOJeXVrGdi3DdLdLDWgAo/LM6jUnOKMQqvWYA
zrlkXcSU+CZ+v7wf/IIS4u+Ouk1mZcFqqIlfWqOqRYoG+1yHom6ZmAswaNNJxj7y
sbb91ea/vGaSZExEJ5bZ+MkWN6s0xVPPevgeGp5MCNhGJy7qvKX02wmilu4PjV+D
CWW5L1N4s00G46MgqeLLp+2rStO9tsdczPNCMw3y/EfyQGNfa1oWd5n7vrTtukGf
S+LMSCbv0Bf67cnhRLiK+wJNz5CqQyAsFxZLkshtgUDCqAjOUjc9VplWgOOJvOQB
ddTbgpJ2ua2pzlLkJ2kM1A3Pp5d27kOtJmLBY6YC+nSmQU4aHPdR551ewYpjZLJR
OoY+pQamUwcgi0HVdJPbdUzBQHphyuUpYCFlT5GnJUEEMJZWbWX3mKPHunRC8wqH
Uem6c/fr15xfhsgsGlIimnMpQawIZvldYD5gONnRlSsRTwnEVgSJIYcdTwS+KLjU
z59C72+hgWmBOb79g8DaU0YiSnrNVbGC0OF/MQ3R3KdWiCYMgjy6PewbotFn0OLi
Hm2R/HXt3ffHtxYZ+DYrjVidARg/e/BpSGTnIeem6MsjQteMZaSRG3gGml20XzSe
EU5cfLTlT8DrLO7srWgjAjHqBTKSDZK16uCp+Zg8A4NhU4SQ9IlcOJAAoy7pliLQ
dvMKe/z1RKeh6H2sljYAbW3v7sVtVZAADK4S+NxK5QwdFlmFuok2L0nKwZ3i6GZl
1xIi9XtE1wC/qqM0fmGLtTrVwW81As61+dKoWGxPaDhdze+iV+iUxldN1+Pjuv0C
kxsLr0589Bj534cy/JVHPJizIC/C4d1U9Sx4eYzTNcglznh3oQVHeZ2K1FhYu7Xr
NLvaWW4S/cF80jzM2xBHlb2k5WQCfmGmvs2UKcLBzeoI29g6ogfTnpK781X+NkLZ
Swp9HTOVSu+ZlSBwUVV6pFMYstgCdb8AMfnas+GG7HB1KeOin5sTUaZqjNPvQNqa
WSy46VW2QfJ+VjNq9RYHmLUlE2Ui0mfn/nX8ukH0BtGDnaTXiJ1jofux5t0IIIT6
VrGEJ1akjAZSoHU8PhBkhSLmHuWz+vTmzZ/pYd1DLNqOBHfRnHdyL5n+tUOFwB+S
3sYhqmmVc+vm9WlmPjz9HqvrTeuPLH7Il/eQ28LrxLjs5IGkiJZDdeJ2DkIT9l7P
ZenIHGdA0G6r88qL9etq8JEBY5VgGCGW65WF8iPUa73bbHKeUVLwoUUoQSPtskhu
i+D50aOan/R9/0sDaCUHtW7Ebscl3xMgot0XiiOHHhjl4T4Dy8F6y2iSVTPpKso1
ysKtG2ke6vgLlV7dTmisIyRyTO8b2+YtHfYM/nkMmcj0SmFbWEg0EO7OTHG8f+Ot
dmh94iq+CElGNQK34OAbh8pHA6iIk0qlph+jZx33q3a0YfgEPjxo3AUe+V7m69XZ
WEPMCMfNGf5qsxfDewaO8MrlaVLDO2lFSuh3MszUwg48NsaSSfbMs4jSLfNgkYRR
mEch1hieeQgavnGjv6o5fSh5nCA7z9MGj9F8ILLnJI7F8VS/DJNLiFvatI3V13Sg
kt6Io5p/KBWKQwB1LxJa+Z/WjxJV8gWoKmhnq+yaq8Fw5NwEB0gMVIJ1k+NSNoza
2OHPb7bkOWLtBgxnLL7vDkrq975YJWOb4jSat5e5hP0JLSgy5Dp2lMHBa3s8+fp9
omOg6T8/q+kVKZtmCsQgVpg58wk9ddEuaX8ygxN7EIhiRC7T/WPZhRuhPr2+yIMY
S6F1fTqxbZsE48g4NmsOqcIlkwd3F073Nva+zI206F3kit8oMw92g2bIWWvxImt7
5+P+PZEseU6ncGFjRLnh0/auDE1rr+L4J6bBIZmEyX3LYvrCzuHMhS+Hd5UJNm4C
WYTVIFintncWQ8skqxqW3Hx1DxP4QJLvM/eFYotqVAcd9TChvXawTesQ/UGr6j63
WurVYgVi0D2FFD4zHl9gQAIpOSa+bS3ZH/Fe1WRJOJ7Jg6d1bWAJK2Pw2crwI9Hm
c9qUSphYjurAspAMEEoScyxRIIqFMii1bNfMpQLMSnb0CmMbvruuBnS5QTfHkRK+
m3PNuS2yXLP0JWzpM73AFinkgXBueg91mTvagfNbZAV1KRJhnraDJ/1fQVS4HOlv
/3JJtyjjcN3th5gA1f9/3NIIl0RN/tLOz23NXN2Tqbdd+ZIgaPIs0OOTaWPbw5mR
IUNRtyJA8DNd7XCER3JQGnHpFtAPPWo75Mdcvc8O9bnBW6M2FBRsV9JQ0qezOnii
JTVYaDAC9LGvpEW9EBb19AB2qUpprtdZPioSSqBLZ2lzCEYV7iq94N5u6zaMEIm6
4gnMToJE2LBhAmHyk5/s2NDQwEh7dZ88VjZzO/taXYK+BTrSQvGqYF4jHc8nf5X1
Isz5POgYV9fk1XbEmwOSSb4dv+IzDXQbVHthsATc+P6Y4p069A0C5KuUbDOh4e9D
D0CvJD8T8t+jkEoUR4BxCFxH4vV+RJQrDvtHCxZDsd8/15t3/d1SzXAXwqbvHsO6
UomOg7TVkM+FhCPtdHc3duzjBJIYZ2h2d8T7VnwwcJTw//hVaZjAYFSOaYH+ghGr
9tpQyzFikmEC2gkKzQl+uW812P5k2dYmjP3sjUPSotYQB23P7zb8XU5nXqUYNtAv
B21CtD6NuaAhYNY3211daAr5Kp2FqjRUEdkot7W4nrZ+VveGz4jyrLQayTXh2Gux
D3cPuzdHdGR72WT0nwE9ntuCHRJAcTTnjSIyCfy5vWjYVIgNOsmzafHNLkadFiMV
Uyo/g/M7yHeS13mPqMDQna2RtCICiMJrVk2sorVpE1LjZ4d8KARBNp1U3df0tEpS
+6RWzSh5IxX4h7wXQ3YHiXi3EYN/B6Zt2tZSNJtNi0b4DamvvIQTnp2whkSLKQWt
W2Fj2JJjb0EVpOOLwVGMsf3qJ1wjAyas667IpgBFPJCPRNMdgciKzb77Lb3Rqle0
gl6Osg97wQgMY804TLxcS1nWkqoMiQcWuDMVNXhTMmQXI4Km5wm1mEtyo5MoatgC
pUirSb7g9pQu5coueVcdJgyWMLn8mAkhfY5bPt58CCxk52MfHEPp6AYVf8G2MW+B
/zSlQpXAxdHi1tzCVI3y5lNMkvcH3aEgZhpTQBltlNJnjcWZxNTbt2nqBpibXCL2
i9AhIIGn+G7unNb6O9WMyphLgZJxhe60yIcLpMawZTyk3aEs2gZobCwCwnHf14tE
P/bqOC/BGs9536p7T/nVoW/XddcGrQnGo2c4TbU9Hi8laal6C8fD79YjjOL4Oejt
tI/XYS5bHh+gTzhwsjyL2sZI0fo0L42div6vJbFJD8ajUb/mbvMe2WT5iAZWPHvV
IWZfjYHO3Uf8JcagDT8Pryhu7oKVaYyOqsQ9awr9YfclUhaIwkx4M3RgpVkgYnrI
2OLDBk1zCVrB6Zucw6Q1EPkVIrbJUyhrQBjG9YLd2OFFh3/0yl9THVy5Z8leyfjN
9EuTRpreqL8BZ6KFNOxcLq+YfNRO4WW1iaB5l+K5tK0sxXgYaTv1bBBSr22u/svj
n4Aeo5gauw+ofWONtN9aSo2NbPtQU+nZGFO32DFo/ehPo9F7xpNCd/q90siWfnKy
6jdQpS8QkKnYDu56RwANEYIUrkVgBs3YdiS4ek2AtehEUUJFLZlSYGKOHiYAHT24
+DCUtKmgGEkOTwINbp7f8Zja+uFLM1Ee6YG+VoA8dDvOSW9n+Io7Fx0xtIUnw5Rj
QDVeew99e5h3KzvooHqYACofiS9dzOWRgMdPkUcuPH+Ovn8gTuG7L+7sMgAqpzbV
q6i0v+wtHiBmzIosjsWx0on63GI0XSsnY8RnoZHTR0UWGgGUPIwD+rPe5bRuIwWL
WgqIIBFs+9fffPp0aIR7mEZjVvvOvKY5Eyc/jv1jD/MAPCCLpfd7jG9JLHJQ340G
1XjKgcF1R2vZII4g7WLo9kdNynLuqRFoslPOEo/36gs5xIZ/dKNNwrRpZfJ+MwEZ
j5bx7qg3phAlK/L1/22ML4q7zNiJmETEvP9lvCgbTXZgEh30dhRNz2yueblomO2U
JfX7ZMBOa7fbMVsTcaptmwj/4OVq2htRKCnC796qfue7E315sg+IltsMQtOHwRQO
XbnsdMT7X7uMV34/D1ijH5w3mfg1eGEL/N23hF9RyZSkt6W8E56mnrXU698kquMq
u/S4Bo03tMCPXynB/Okplqe0veFjHbLbBYweCqaZTc1FN8TVJWuZHx3TKtK5vO0D
RTE8V+r5NfhbBkCDgQ7h10NKE8v6ImjGUSsywBmjnTOminKorwOr5NXFm8foPSh2
5FhjX+FHl1YtOHUI37eaCRH5U9bYUs448lkvlP8PdAkDMReb9s1A08su8s9hyafv
qaxTor8H7HQbQW84tpWQT47Tc+wsqi0P+7pVQ52lhSVzOHyrRi035x+pAZ/9VPEQ
cbDuLEqdWRUbOE1ZOXUlpmOCeL5LsWynIvlxF66lxzh0vPHWP9SViBmOO5JQ60Dt
Q8fUmJyqwff+rvqC5qA+ZoXVIo1/qjPtb7nZ7nHB+Tu5L1HRA+s7RaLSMygqxR1f
rIzUNLE0Xk8P0a8UIaym8Z1TmEhO60EJ0a+n3JZOUCpsIv2qfy2QJEwh1GDePYf1
o9SFFLseDIMyXAgjzGVJzi360sgMSsil//dcy34ejnkRKYzw2UXI27bSHL3/8bn5
HrXlGeJjCD4x7PUdxkCw0ncXpZpPGrx06EVR8e3qZSfL+bciV/8mnBnRmHoodr+A
mQoD8hw+j26vpcqq8R7/ceVHf0BqKuTFjxrK4u3W/T++dvHKqiLMVVIUL2bRjN+d
4HOYAz2sZCQixebwX5+/ZyWRFdbcRFCGlWCHr+Dfuc07pT0tYtKdwfrE7PZAmE5B
EbaikmsV3PsIhAggiWgjF42pEz1G2Brvs6ZRWFG93G2D+1d/A+bMUul0h3eir4c4
2jUy/Sz9q1vo/kctdYoeYKKLBj7vKA0nZ8vBiSVIGWLS5Pu44nMaxBLVm8Wt9wZL
hbbe87gt0ki2wlpICWvzQ3B6Qs+NVTxBl2qk0Clb/emATwrM4lE+oI8WjiY0dI67
fx/TW2MtYu1G6bFnZfH9W61aiqgyne2w3n9LFXOgwdDLr9sZSxw6jNo+nhLEZ7cQ
SZ+2VTorsgAACvHfB6cYXpfJo81IoooTleoqkISWEJ28rI8Ta+/x2/PCesaMwlmE
VFYK9MxdWiT/TDFUap7nHVaMR8/j4XF9qAPLq6Cp+0KGmXEGVRZTjuDrxsD9ePQH
qfYkEEC3QOqucobGZXZkX+Xp/jd3i+fBRucpsSPjwmISoulsYZdd9h5N/EGHc6Lq
m22muSDRJolic4YZnSZcMkuX+xWs1DCkL+MQeR9chb2SjlwS8SY4KQJTyU4k09DA
FixrzkMJeAvhUeuEx2oDCqYkU5MFRn5T5qgrGSWHkwIEi2EEnmFclgUNbTyoKMtX
GQ8Db4/boyzefbg89M5E/VLpv5BqYFETcFSfJJoub43/s8f8268c58JqJkac3hbz
77soefd4XDvSGeBc1HhXOP2S24J3lrHtPwRpABjjI76498LD5lBnJfHConww8XI1
ds2O72kVq0S5HinC0Rp+hxwPcNdRxlmAoM2ZG1urcBZ6wkPK+S3tmbuP6seScS5F
5qItezDcKE3TBkk6SAVO4NC40FEQzW7EbrtTQmaYGx+okkD++XIUkazAybOsPfrG
GgU3AxOkGTo0XamhyFfcMom2co/OBbWOFMm78Cx+S6VDVWKJEE9S9If2OM8kxvnr
DMVi6anJbl03zCJQvV+xbrEgLh338p625eJDuMoStshcrADpgY7j+/L6EASuNkR+
xFz6xLOuwRfU2OGR2rVQPJi+sfhODG7m0GhS4JfevI/UVV/e5yrdEaNzDn80eRZ+
QdgAKkUnLsJgRqIgePJQK3ESlca8UxlcA4Hv1QYDTJe0AnFRZy2I0HMeUiPsh4OJ
L5hN88BGSzdAsssWWIP27D3fr4KDqARpNl5nTaiQG0tTRw39nkX1Iv0BInryAKsK
3sEIOQ5aWe2tAN+JFlDwo8BYI6sZttiplrHXgI3CXQp0vOqU46V+lHyV2R32YlJo
UE252ZSTwgwZKZ7oRauR2ja+0v8S1VfcprXJwKaNEuZncWA0ZBkGxvCV3RNnuBtz
StbVTXDOVaDB/Nbz4Xtu+bNeOY0y79SV7NdK0sdvOib3JTmg3DUKw7bEt6Bga2ot
ctuaDrfOMWVC4+mFH/wvHqDt2n/5/HgdALxEvnNpAVQ75zKNnGNHUb4o2eKVTfi7
bJWkZeU7yC2vfvnG6xjgSqpqEaObYSSC50eMgcn8hBjhrxj4YPTiwqsKDAR4hYqw
7w+2uzVwUn5DGO2wykwAIuNEGHYEor7aSJ7tPIIAIamPK2PFQFcaB0YREtgv1JAE
gQznn3LH7oDrWzIkiJNebnU58UW4hnHGlFTN0aA/DWsICbrjNIyUSWEs83IuhyYw
X+FJ64XO/cN86ewsfjiXLuRPEkAe+kTKbEkAGU5bwxrCnOtVQuHMa5Jseem0wFmY
guyKZdtP2wOXPU+zOr7L2AhpMKu8OTZi+/hbz1tNiPpRWs6r0U36rLJvD7zosI5j
uNog0KkJpH6MZd8vnBh0zYIljRQ1MX2KBVQJ8qRED927QAZLOhaPPqGfxe7d2k9j
1IoiG0SHWjS+gB10PmLqRgDqJlfoskgxQ6Mbvx4NPd9aDWNSud3tWPMqCii7OHpG
Bch8hjSnn8wSHLpoZXCIfBrl4qJ1OZxLPgDGjYiZzcVTmdUngwUnOLFXo/6VAB6o
JgzvKAWM9dozRgKLisdDKYS2Xl5wzSWEEB97Hzne/P1TEXfMe19LM9rvrd/4cQij
+BmXtGyYZX1f9IOfnKlYXAT7r/3HdwX8nCjiXKoq/fD1nuUMdNbhkOpGfJ/CeK44
lSPMhhiTwQBQyp6DV/UleszLK5hW+FIPS8se5Mz/oNLs+5ozU5wgn+BrliTod3YW
A1PSHjDLM66ZWqCdolDNCwmIQSRgWO1yfglrYl8IPmEJiQecZcn1rZ5PdOzWqiyA
0yVL/5d+XjW0YQ5FI63ie9rN+3whfdr7PNydi2Io3V4OpMykBKkKPFt80VjVU0Fc
m00tf+V9HYT+SxCrmHazdphTy9CbLsRwqEdEMlFN99tNVAdma1Av37xb5i4ss4tA
C/QSd+ge0SExXZjI2ODgNtuChpm9TJGr24ayV+u1c72rSo9CAhCWjKeQ4JqhNW7/
IAL1D/NBtwvQ6BKHtUGSTWT7SXLrqzYEd583uPkSPDCYwj0fa2+G6q8SM6oSu9O6
zHIPv1POXixbGp3gCVYMwzaBhxoZQyDEt64Fh8KIQFGV173b3N/w1dzdmYtJH+k/
BsTDPI07HPtsoHjKP9SAUjcBNIe+bXgIO1w6aWzGXLJoSPICvgB0ILIsW3zfTGC8
rSC+08pXbh6p9yOwMcT1IyPAml44p68GJ7hyyJiu619cSgjP7XGOpvVnDA/F742s
WgN17Q13u81vXb3kc0imt9XLdKLuieodBw6nA/qVCMmGeI7G7vmT/04rn6myIm0F
Xg4uZx9Iqne9WRlEYWr6ppTKag2qI6875uaHTR1IZw9+RjFja4mdowJwBxOMfdiY
daoj6VKCQzRd55D2/XmTrW2sEp3IpHdZJalrGY8aoevBJ3BfMcCj6TNFkmkIPZJM
j/ymTOTk8l6fhbHgkKgMkl7gDd+rc5VpFnhzfWOx641yvlVsaNSdyjFyt9R1g266
+fS3h6l9xRv3Ap7Wf24//ZB8aiowGM+It+WdnNh2FVvfNDhnDK0fkWbNdPq6JGJ9
BL2LSA55GXF2U4yxR4o+x5RPNeXLsooTy3RmCWrjW1TyrWa7DJKGFkkvGP9TZn2t
AngyJGMO082z3PiUK/qJDA40HnHvV+o3ebFCXELiZEVxn83yU3y8xBodMyK4aumd
PNEb3GZn2RPaOCrj2K1sdlTdGcZq5GyzosPMK8HnZ7PaRJVqimjjzKkQU8PmnLLo
KsZJm/P9xq5OR5/MZl4lemaqZfNjOiePttlseVxc847Yum8aikzaTUeONOszukzj
/EcovKTJ4dkDWVsQ3cC4rPJHF7y9NaQOuXlqzGVIbjIVHoQedocuIJjaKi+t7sMk
0nthvLJWqn4Tc94Kt5lSLG+XRosb4ShM3wymzk8Hv8xIynI26BansLOZoUjHdYNj
T+/+b6HsXEpO+3XPq7xpsU+poDVjqOBrTU8PYiaWYRDpWQCw7fZIrCOEVZYo79u1
KqbUHXSuRxC3OeYRrT0RPAwNPvlyjbD/3ofuWb1o5hDn/cBZQsxxrt8gGvmaK9Ph
wC4oSiuYIgHPPLjSc5PT5+DeKysgAwYWpLLksQ8Tj1R2lL+nUt8xLxsP0g254GPL
20K3vLEWl8m8K3FAAwGmsOilevfUoUuQ25QW5r8Jkra+oSSop2X73KVKa2gmY0c+
D9i9T+mNmW48wUkSXiSK7bNoYaRlva3N0zbTSps3k1GpHEQBsiYtlNqfV2ljzNwX
eP5HoY5csU7kAnUv3n5V7VmGAupF3io6B0b7RH3rbUv9gGGmuvyJPTr3roTATJkA
IjMoKrWpusqeWG/57dMywgHMtbzUIRNIF9b4xZRis5Ukg4eRauMEilULjDDqzD6z
bqQYN3kpbITE4/jB9RPPTbRzSH8P609i5nAl2lcasDSdDxhnDkmDO8zD6y3DP/bq
uUpAxsJQCBqHdQ9xrwjaJdfdOUySkUUN7nRhiHIuvkAPDcZWdjy1zOo8nEzqOkrn
yUwu8xxo6WrxRZUf1EIA9ftCqMuSuYMzGz7T/FRrqgfT/o5y8+5oTQD9iOrFjCfi
R02wCKqmCzfqbVZPzhHeUM7ZUJt6Bior6vvkQLUOvdm/AUR5cD6HllNtlN16mh7p
rZFnG1mkEn01oQIGFO6oiJiKOlNhL1s+EHg4Tigf/eew5GKTbSCM9pa612zRMcmP
/UYOW6ZYCdSss5NaKzQkpmJYIV2WmNW23dAtyA/ArQGoUfCspqBAjqP9w+rl//ux
NtjMmuQwYK8sJ5n9RQ+uPMSyTYthS2aBeC8lj9dmGcX1+O0xPIEKbV/LBj9gRBPp
kO19YcSWLPRUYuxhw6Uyy3WOkfucggGs9K8NCrrISg8ucNvhe4Jg6/DODHlOynFG
uKgjzqaj07xsJBh9fBcPYccHq9yJMJ64sM/Llngnmmb4dFxGhSmAMI9txjKWpA+T
5c8hKbUtV45rOBb1ZIHcpR6n/CLVdLsztkPyCw0g0/Ddp44/38GK0/6DOEeU+EoH
nDX00XaGI6MtnXCDpVzti/pPN84za9ttIMdGRXalyTykbfN0RkeKHmfXPxJKAMDj
K5KjiXBliYYFnMPyks/er/YkgJzPEednekKTeLJ1V1XoVp69dUsSHXbn2BZFUtP0
BRZrmalh6ZnzqtdLTQdwmWsQK8Apw4EdNMxvivj0QhwqBaU7wuP2Q40OSSknPcMh
KIRczWlVdz2MlBjqaHKlMDqSYNijGn5VxP8jxlvToKX8pqMbiR+oqhcODrVOp4gN
gm8zBvQKYU1lAHaAkEcC729po1cYnX9od8TDDkhs1/NL440l0aV/7OjCJvt4UW+O
D5DO+1esofvNQ4MJt/EAxzE/lQWoKNH3YoubKS4hQl4ZB0vwBPrHV2+eNeiPQ4/S
1rJGTRBlAOOrfCm03fR3y2iFuZWzj+IXvekPPT4G7rgU9qc2+LxDY/Uz6sgmZzfF
gxjfLThdmp9weSZmKrsp5Zko1Dq+uUyPyW02EUKOljiQeL22+HtKN4ZjVwFzAf/V
c4LE4xiLsMevhf77xFAgGv0F1IluBY4J3xGNRMP39dOxd7QAItE2Oc3AUrg5ufGg
d47h346L0nrtl2tKms7HunUAiegfEleta8BlLkF6Ns+8Rk9J8If/muN8QLFxzUCR
s6mNmW01LGG/ZO16y3ltNuJJ/uF9SaCMpcCw05b20EzCax4biXpmVh6HO8ld3ORU
uhk0BrYk5KZ4/qoFcEBeUpap8IqGcL0+LwfbeATWbHAP+7AANtQtO7ClbGDy9dvc
qjIFsLXz3LuVYLPLCCUwkipNE+33+EsnHDJ+RyLZVv9kLrDlmpjbssr8PREe1Yp3
GhiH3/IiLGwBDavBsVYuneImvEwZqagf6T2RPOcGCQ97dPg+I+oSpGLICWajarIU
APfj6NX+3Z31DMbWLqqXIiY+Dme/dIIXIcp8+qmEfYhd3m8BDkyPfVIHORXkkc7x
hSKPL2IVVGjKUH3B8M34S36q9HWwAlfjNX8lpfdUhgjJd1FhvBtP7UuEzRgdnnvG
l2eZjDrXLyv1dvJ7IOQUA56HpJklTATruIhFp5QAOEat+1r25nBqndlHe2XShfSh
34/sQfO9UozSX96Q3yU+cRvm4T/DMqrsa08U4izbYszvqJG9yPwhOWUC4vys9Ax/
MZh3leihlf09khM00Iw52Y7MawpAwUUry2kRcEs9Q7epiVaNweT+I+LNoAUTClGU
oIBAIwcdNqFgbtJTnN1Q3t0nhKwR1khl24nn7d1ULptEe1AfLGkuLxhOAGP3oyzm
sNWdYHrCCdrBbe/aaWcZ5LWgerxAA9uI6QmGG7k7d+mQ+lJ7DN7RpBZmEA8++e9J
JwdoaW+vWWe0WEm4gPDVHh8eiAxjTYLIVx8mEroaAHKZFbx9x6cR2OvTwyJgzj1F
zKlnF7h7k/rWzby+4H/bpQXV2i+GmibsJJG3HOmNJj5GAzg655bHN3lt0AeSqtTj
ek1qqEPmYu89k0l4OHEGfJFCFpuNdu+lcjdoVXX9M0Aaw5cXxkqDvZ60Ol1bkCcZ
+V7KZX6CtpiSjD8BmwvCx9pmQ8jNIk97UFqKQPlPPRle5XjnkZ/XrfLmKIhDg2Hz
n9BKFkPDDDPdSnSCEbrFqIh/Wcf/cLu7V6nS3VrjbLZEjQDuAHmF9WtCEkLNHorO
0OQDIhB1L3d2V6OITIns+PanjmRpWyugMWkcYDblFFRaGyAgGsQKBEy/W10MEXRc
gF0ANJ0b/erCXtVXl7DNnUb1hl0mDXCG42hlpxgw2g5w2VWvATFqBFdesq6GcI6g
2bxak3Ow+CsvclJz44LlcYnSOc3xLI1hqoJdhc7rzirHLQTBVIAWolgotfRyVba8
R5Po46y7AoD8nsSIrZtCGViO6lEDiFlyEAk0l48ykSv60IMoODLS+AYU3P92+RRa
xGb6imoXdbHIXpmFF43jp9ltJK1eM2/8YBRY9OMGIEWhbdqOffvOFTtZfJ2buogJ
oC1mqQ4TSjr6PTJAEI3vS95X5mw8f0czM71/poXEqxzMo7bE/IjE/OoncPoeji8g
DQLzk1shiP1mjFzEphKw3UPe6Oy5H2wsO2p3YUNlC81hH2j04bFAV71itIKUqCoD
U77cTqI6bTqCaqgtNSBnlF7bvm0PZ0mhv4OKatla3fDyEJJKoy1/0rqWpbtdVXVE
WgdTJCJgTtNQL302Ew40REqJVjAYLNS+MB+QFrX+rfSiWIxhWsf78iD7KgTAjZoQ
+YypoqJqPvI6sMm0llwyClkJr1oCtsWPGsiPt9wwdFd0gnB4AcvfwB2L3vsq9G53
qMpYpsPa01If60o8C+KC9mq2CFWzNz7adjneU2xSqL8swSQ3fofXHH3QXnz2l40m
7PxpZ/wkyifjowapEi8ir+m9lo49lozeWnt4dpQGb/19WsUi8sdAnJsGCzxMRZ4N
hbOuLdwcbwCCUhASsJhQzoKRa86fQK2Im6hg9YnyllW2Wrs36G2OKJjLHBCJ7KRa
cye9NMCsaseBIZOcJ8RnRMkC4proAn5stzhOY+XG55GpwFY0F77OnyeGR6Q2OI5n
v+0N88QKlPNSeu3sEZlgc9xvoGtfRqJZ39nI3YSnCD07jFp/6gZfw3/BZmtIPCNY
6wJxLmFMnV+ajElcw6XOuyg/G2r1pgxTjICkG2tkk2VwRr5elNTAxfhf/Qw13gRs
yfLbL+G7AvWO67e4ZP4MekKWDHyZb2p1cbKorCsQjx46CeuN1NuQmbSDOIFMeuq+
XAFpYJAV2CE6+6WsIRGWgVLdj52WhFhmj2mVZbT9dvk1gTdlNDqxj+ubOZH6sFrn
4fQ/+8ZOqoOSr9PSbd0DuFDCq1ueb6YU/eJyVD5ryNjKLW1YAsS/uSffko9z6bxE
Jq24hKhnCpsY+ZIvaIscekaaLPgykapwyb8Hxtrqe5On05Xw4h6qoSMUxKg5H/3N
lwjMyY1CZp/v7soB4dyyCxqch5wT6FBIjqTf7F9eD88LSSLB+UV1QiM+eT6IVyDA
yJwe/S3t9QsgafepueVTQmRHZtb4TCQOpOYz8kxZkrVkxRLVupGku5woGDYiHT70
Ovuz6ExVlgrvWaUzuEsmlkH0ApZZorSx3jo6oKPWoJzPOnKn5LYR/ViMJeN4PcTG
65/+DLbe/Fj/gJ+I3FEzBbloI40dF7e5Gauw6IFOANuP5t5giZTmEJhYH+4mpWPr
Dk1eKlQ+djZnj+bdKKRLDXbOQlczNUV+t/i9453jNlwGbKf672tUL7egVJR2XTdw
M0/k1cl7jL+kleh8YrBei3aEoHxvz7G1Di2tGtyM2qRhM+GbFvP9knpNkBbIIk0P
xOJVCN2RML3PhoEDJdhC51ODI/XXzbIhIQ+6Yet9vluJmQuX8svWwyr+FMEm3G8S
TtCKxUjvExDKXOo+F5XNoddqDCHWSU/3bPCTN+19WOiJXd8kFIx8WPXrMmvZ3RH6
mFkKKJ0ECatwHowXA3Nse9At3e5l9Z6uD2Ey+DQgRfH+dKOScVuPyVdrOZaQECPK
M4VCs9VkeWjJkDDGmaqsIrXmg4z4UBmrNTFg55s9jp/ey/TokpOEw9Ax/1khzhjA
ho3jflwph1qODJYUwhvu8y5WHNO5YVfanpMeP6JyLW1WBX9Fa3NwzJmK1voT5TuY
ueDZIt1RuWwOfF1UkF53J09l67uJBvt26xI9tpS7XACLCAbdCXHY8JXiWck1keGs
6wrr/dCTGwBtsXDRrTDL18Wb7FBeNLqLJyonkXUU9xP+xakxjTvCr9Vm/pNWFCWU
Zr87AXOtPFeeT6TxaPeuii3FSS0L95Ij0IW1bfrFfqHQJ6TqoI0Ls+VLHu62NMmH
C1rYL+sSEfJjixJkltDHqdQCdA8SZ4mseGWIZd+tbfPBUtsKnQS19mvcFNum2Ppp
w3vo6gktl99izdQTyWY/35IcX6fFuVQaBHMlhSLQXWEmOB+OzChwneesB6CvipEu
jo5VmW+q9aJmCzzMmCd8ZjKiSd23CQH5RM0mEhg3cgtj7N7lxJePWJAGgZ7j20hC
2ZOLKQpE96z6/jhAZxNohMnHhcCTML5ZFsANWb7tn5JGsIzVirEWaLppdWBsmsLa
NDoSrVEixwReSIdaCGmGernBk7ED2DrRkO/ht6rVhRAAWrXjME2JITdUQXQ2I0sW
ahcZcL9/+UjtnuqpStBkNy6yQWufd/yMMrbyZGC3DbEXmszuFqVB6e6Mjhk90Pox
U3VekhS73aR5aa/wiaS4TtM66DmgA55jXN3t48BYQ/m1SloFURmrln65Pu13508H
5I0rRf+2l+XiPgMl+LoRIqQVCjaA5kQxFN+DIoUfmj1kCcZJlPz9/WS+cvv7m0Kp
4HAXy7kmjrCzvwLzTDenJQqLNttZpX/MMMIjej8wKdV5gStUZEeIhH85igw7tuQf
KCrBmWjbG9vDR8emKVCLLYVOhdd2Vb/z8rLp9VM048LaOhqMobTLqsuImBdsr9KN
ae1qe5rtwHXxCPn5OpA00tY/JEFGjfaJDs5ypBcJ4W49tBRlAITmRy9/2EZQxGmr
kGG1tZXeGCDae6NrxrRBkzDZcPBXUIen3sonadlG6aSJhaQRV1XmZcCrC+l+BAKW
maxCgdSqsVNEv18tzs+/tOt3gwhn+WFGsgmjTm7Wj5yCUqQixBjHHq4I7FfgC04f
gcZBiWxSXEoZdlM1FDwOtzLe2D7cUj9ye/fi88+qqXzvuXrZymGyMWQ/1qffntYs
ipPieUEQeap1jVkQ6+C/HE6veQCb5VFsG2DOZK9RQGX/h+/pCl+dp5m7YbiROOmA
0rGQz+mc7EcUPeOQewVOTZC1ulsOGi4RvfGT7JZLGkYtvhRx5WFySycuCpPbtafj
QdUChCH6nUPAl1DcfP4rlVANpOElIcWt0U6mEiCMTyFD/+H5AYaJ0g+K+Irp7Vfh
aUi2uqM1etC/PH7xyDwtqSABxz6XjJ4B8xbx3Q54k1PMqVL46RD17iFc83bZawAU
WyWkNejnquCumibS50dxP7LUun8cibzGg2fGpXKgf84E7iayJKD7ynzrgRSU4IwA
FBWO3WKA1OEre9/Quc98kEdWgPVU8DJTuIdf8HyioqHRGWKBOD7Ufk+HXmxgAkH/
CCrsjxjIamcdyIE9q3SfoTmixrESpFWy3fafASpKLQmMKKp5jTFZl+dBhrcBkZGB
pojAvsyJakBc1kkib3S2auZRKhPGKMURhkMJdmQiaFO1bmo5+WUcL8EtYbNwIU/4
JxFPmHuMOQDe4QKj8saNS3jkcQDU2HBUEQmal4S0VxekpWsDFmlzyrExxDZ8/bi/
W4GsPPfOK3HIHpAenFrfkzLw/EWbqxIjX5zPFiQFrfwUv1FF4r8hPDI6CoRSO4U5
yaYg2JebkH6zLAhBwMNqvE7/lOsetTjCSHeuN/bG34uOVZqRSRe1MISnVQoJP6ps
fG1kqJ3Zcm7iAtLifL6QsdLKDMZPnRvDuxdMrDjrQb3LQgArfYaGZ6CNRs31t+TM
a9wtr91jy3Vz5z6Ps2EjZUn9++kATdA4UIY6rSqyQuhw5VwoDip8vPHBzl4jqmBf
wXlzsKf/l5i5KCxSYeqMLbBK74VggWP2QsdybZg869kKTaGq6nk8I7wKSa9Fh3yk
RS/EuzT7yKwtx0HF78JE9l9VDHMrJipQGEszwq5HwV3pjboSzUngB6UgCmXjLzAK
aMJTbEvM7k/cimH2Lrc6ktpP0E+LClJWzu/nhA6ixgqyUma/e30OFJZrvjfGDcCC
EJuuLNFnmY+F0Zv73arDVIcRsi2nBvrZ7FnDC2kbWE3U8UZL2xCL15b54w/u+oq1
LKTlqByE2hg5Ywz1b3IPir3ZPpFWnbtIaUGPTx95NvqrY19wUqiI6v53ZpVkDYWE
zbddbwNH9WNy7XMlj5Bw81X9cUSzwQxwl7LFsgcEJg9ld1CWDEqw30my5EWkBunh
2fWgC4Lt8E/0IFGe8v/V15uCoLHAL+x2pVAMvRMxJ93bAHAItb4wHS4vpSvjvzsy
XBvEAcMdclTirBru5bPrRU4qFL4v3vB0hZkI1EgcCafkeNVGa9kGq4N1YVaePZiO
BgCAyqgHbTCdgv6jNYB/m5X4Ar3/t88MSyeq0ZYQi7YGVvjlyZV0ZSUuamMEQx+d
kQtErBrrNWE8lUbQMUAGzdMNC17ITJW5a65Om2VQtuy5EZ8rUA7JuhWPwaWNNKRY
7X24yuIzyV+bXIMQK3Cu/9Ipl5QgYowxhHil8yS1dWBbbdq2fHNe8KntisRi3dSD
Y9ISOMVYuuijVbogJb31bd0IMQmZNo4zQ+wOeLajTIGf1i666giXISBgT8d6QNEk
hC85l3ren+sfGpBi02Qizo70spvbI4kYzor/N5XL9pbUjYtv1brOmAOsK4bTWtpE
+4/aE6AN7XwY53v0BXxHeUVf8cnUmEaeQpl84lvTcfD5pdwHGSEhKviVW+394Sfc
tAXfZXraniL9TyRT0pCr5LrpARAHG17Q/TYPbxu3AxQ/RPTmqwlUong50C+q5DVj
WSPRR1inpZXY+66M2eBEjUSNEz2BhcbL0Op3trBafiWeqJ4ybXHjYpsrXgi8zNjw
Uw0qLoQhfhA2TGusGXdSpKbcNoISvIL528nhgHJbxA8wherm9mYJvvkTf0OwL5iG
vB1QWp5X3YAFCbT00XJP/qBf839Dv3hCN8n7w186hmcrfvJzwL+DxeQTo25B4lQm
Fcaq2XSnCkPsE79csd31MhDCu9EWYxtnE48cfFUrPnocMFEehk1Y8oEzSl0I7LuM
m9dbaBIUuRqtYFTeXiJpxVsvm+Az38KTUau3uW0gdiPTgAukJz2GgrLW7Vpm/o/u
/LXaGO3igd6tR83YS3aIjbI5xEpwenXd/FTBWY3QFUu2CL8kR16BT0hw7vwy/sQq
gyeY4YyiREqqUw3oDzCsgbaBdt8GHAA0TOJET1/QPDFUFDHpkuD1zx3FAZ89CWp9
mDyYYfY7nZI2aTC5bEcW3dv15shtc4JDQAyyo/uuYN/bO3hNTlPKg10NKprLSghU
kEyVDr9dTzuwQIOSyibcwh76YctNnuK2wo9SaUyZBK4Su7LPnnjgs4aZO//LqpDV
HGED2JnHNGtAfFc6RMbhF43wYaXoMPSefLK9+XSD+2E62nF4+wxDUBkyJGIcxoj/
8qlzvANKt73ZRZNOJrYClf5DClSTr38Ilx3CZCnrmH9X+UUeXzcX13eDy3r5ndOp
NdsH61kcONdflCrPhAnI3EpnrzzMQ7MeeamcrESXTE7p8w5AwhsrZ0LDfY/VdeS1
pX1qG0QXd234XRCsNzHbBrtPd5PlQ4OH4QYNv66GT/qRpx8ZOpRXC+3MHmI8yFDP
HuCq3eT5TR5ga+y8NDE6To9zqp1WySuYUDh89lVJOFpk6SUlLWOdvmQu7uM3oKp1
+kR1xYRxPfh71He3FhIT79QV6kX5gCtiY0PivFJ2fTKB0KjANFNZxDcrdxmdzKin
FbtUlsxpjZJSuHX8JWAZ+iq5YtNbLib4zCZUuxTUaymRD7te8m1VBSEmKgR6SNwQ
9IBJ6M8GH2MqgiHSbfgCWFq+fK4aNfUbmI6Fil9bnQLjgeXJ57cSfigRy0uLcHev
kBuElqgOZhKxPnzwE33KcuIjhU576+lN72AP2vI/rkLBRQXhlHc3wlVSTMhOWdGv
Fn1+114pyQngr4uSMn6YJoqzUQZz6DgS99DdziMs2v7TkccHMRBNGMehyOkhm9hR
RCzGVQiFAd3ZSLX/vcGpvHmdj6rO5V994lb/SMswDO6xFTfaRFfd0KSd1G0D47jz
SZQJOELzA/Q8eueLYBzmLedbhloJX0+iw7w+BVZIhvNbj+TJLKYSztYyD1HX7Bs3
7M53lIXQa50ypYkQ9XH3a9zbFiOaqH/e4I1GBAvt/lituMptCWpBfYe2HM2ka8JK
v2s+hmW6V/h9OQKS0OWI+1/4TjnsDQTPhd1YjEMfQ5A8i8yk42HB1y1tDtM5x2iJ
FIJOCOqItVfitaACZlV2/QLKg8KYHXpNVTkxBfjYDidGYAXYVyxDKvF5Px+e5H3+
zluYi3aJxJzhUYF6+paBu1i36/APBEje/53A2/smVoDB5K9t1GoC+4/Bb1RJT1nN
/EunADfk4QvGqSN+lqMjpZXg+M9XPi4AMNAb8r75JtfSqRuQ4g9AeRd374dq5kQo
BsEZVe70NLCMFOMm5tfjPu/SfTgXaFalZcusJ8uN8cKed7PwqF13k+H9MnRWrN/2
XMP/yUO1ATfAc56lqBbdTiAUtsMGTJfs7X+IJDUifXOPSh2oX3p409G5YTHL49vI
efZFS+HU/SeTMNzS+s+qzFmroSRgqSXruzuOYDhmr6Rb17mdtOFy7ZtXv3MBcJCB
xf29opfO+IwKCvBf+A06pNrJKVtnl8Uawg9fgStAYhjJnzpfL0RjGe9pK5Eya10F
QtWLcB9HIWGZvHzSgFCawUEm+dZcHQks1Dfabww3y9trpM/hyshFrYSaXNgHjIU5
KOrVIJ1o+BlxgrZ+BwbstKZlFRUYMsC3pHcl5gAv+VP437wrcDYqPKMty1TZtDVZ
IOEh1OqdDxZZiuTUOEKRRa9ndLyizRlq0yD4yEMcx8GrxHW1txtfPr+lZcQRJh0d
KyKgKKpGpiUfTLKqXr4kH00IaEVTJb/bGmDXJ9KXX2u2vJrvYvEmMAf2f2hY5tbc
KFP+80aTbXFc3eGGkuortfoOAkbd3b9c2ySKBlptPqZiomgde5cjs5U7k77mUPBA
sZB6NvvjY2r6oFgU2aYqU8oFO+p4R4vRUXoKGIg2V3Mb13oMIelC4jNFebDT1zWr
rm9u3xIbh2VH6Bogw5CnWSogRPqLqt13cKJv+BTEtPzpU69SX/uqLl7C8ZewRIQM
0Kzs7E5r2xb7li9flXAxDsNfZXSFf3BbjqBiVkR18MNwrVHc8uY8kk2f6WRVp7J2
6zJTLdBbyWtXVMp6Mdn6R+NOkUWHfmUKgJKTabl/S9qOANVcSA6SOHgLhjGYfyU7
5JrTw9e7ocfGWdZ6xYEl8B+xTcJDXgeZGxOQPdF2rEa1tnQr1xDx+4yI4IfvX5Fm
jQ1weAOh26meRtYkgRGNIQCu7tj6P9CKA0/yHXsAPr4sdcAqQvBuRtlJ7E8GAqqh
2cj1q8pG2O/xsHLRoLxTj04dDDgQJ6UQ/WPtkZWjXC8sMjAjhY12UavadAWx+Ujs
tuCvxveOG0kKbK9cMk/bRi5murGukKVo8iP+u8LDBtDotK7oOAF9K1eXT+5Jx7WG
Ps5PdNrfLskHUFaRFUEuDJdowC29DJIlvhvoHoYOOPmRYJ8RfSQ8Mv7mqxkPjiqO
6/z5Ep/xs4KKsqVEv9VtBgDyQ05jE8cmtgl5vVg/elLduNBc6kQImw63cszt1a0k
itE/c06IAXBQghO1oKoga7vF1nxxe3hqqnXU4Mykgd+JA3KBWNtNQ4XWfkCvTzRp
aD6DLAYNFMxNofM7EYsF7vOMf5jmpZw61lGCFY1PaNId8zInfjqTKecCZrscyt3T
xqrGrLZvu/H502v4OEr0Ro78GSRMKoxomY8xMLSgRXoZo+ZTz4iwxPA3N7WeSrCQ
CZ628vqfgSaVGHYTKZ3VYqlPRYTr9iQnfOHRDoXX35kC96hiYsRU7fgTKIpZmQs6
4HUwCSSjx34Lkxcxg74/yWNXEbGlEXHNQ+6xRCRBa02+savWMuZORredDjQniMtL
xDq+Bxg0sx9w+3zjO3trXD94y4IhgziYFocXdPCdtUYgrWafiYG0SQy2GZ18XIyA
yym1P1HMTS2Mx4HEW1xfvDKuY7PwYrSaMR1ndV1xNiEmvu40PodU7iZQ3hm8fyDI
vWKEuLenHomCr694naf9KT8yFK5JAdQIamB4RufAPZ5najKvZYei8atuKUbRywVo
aeNxBCkWbICc7w+jcaSPkgZbpJQYcrNN2rAeUnyicOgCzmILMFRR9xjlVlthj2gk
mt4V5wddh4WOwq1fzM4fyhlhnW2tLBVDTf3gCNihYlRXj4eYPCz/8Ctpll3GAePz
JQjJF/ANNhCU+EdqUXnHCdXCeAQWxlF5rahWkJ7+/RCAt71CEE8HPcvuk/eYgRHp
bKOddSP2OjVkq6kb8yYgi7GdsTssRWdcVuJxRw+4kQGeL/iHw/Wc9KEj/oa+KIbG
rb85bULdZJ71CphEC3yIcrBZk8Hh+5jxMgYvSB3ZaSN7l+hei7XygfOnPW1osa7O
egB1QRFu1dRDCm1XJ30brARE89sny07Ew1Z0zGGO3GLgChb7Jo2NDtMqksrJ+W/F
zJLrvoMYSfNN710dBtlDSufaI5Xl8ItIFtSkxTETa9OerJZY+gvcw7VvCE7meWUW
GQyszT6hFMybwZxinhMqkx7F4Bm6c25I8VzyUr4YJOcWt/4yxVA0XoPV2iTZ9pvT
FlBw74CcL2OSzhjpFzA3wBj7WJTy6VlESO+8Iu92OjDhNbGmD8SA6GLqZwUNtUkI
9uMhD1O741KdGN7+TCEtzdhJC09sVzNnX9wBONsGQ+wl3r550FV+fTrLfMF1xqJ3
uHspY+EQ9RiA2QphurI1uqR/K1f2km8lXd13m7mG4EzgGFOHFWhLG9w9hsAtx5a4
9EcPA3IUnx9pC5crT8di9dhooA+2i5zK/OC4VyLqzKGOI7fIL4KnwSPCjSIJVDQl
fRtbBsx/md90nguNzNBfWFTNzR0WpNpcWOBMM/gQ7RmQYIUYExu0wl6QAx8GHrof
iXVhnFvovHHxg94YtDakfwpZE/YvJJ6eT1QLt7ENvVv/p+5la7mUkcl3OwUQI8Yq
sqHcVL7s35uiVR/Y1yR50FfJUNk5zrp8sv/DcZbE+joX3r/HgpYLjIf/bD/k7ZZp
qkFE2iyBue/v904f2IPqP+j+tY+uoUdMcJGgK/C/WLSsV0bjoj9p+6HauHWDvi3k
jNWi9xN6F2NiTTNzEHEmzf4eHdO/TOL8c6222fk31KCBgJNxd56VcAFfWYLog0eP
mdijPU8kWg+tTYtcAEoHr1YbEmOsTkFiNPvBg2mTv4URG8HKpK+zyNYKbfMipkGO
S7pHrc1fjmiYZzZOCOJ31A0Yh7EYL4A2flrlIXyMlsRepbQGxCNmX/YKxTDf4Ehf
UiBJapURdlAZY9XOSHw0u8Qm9LcQLjsYdOhMSyKOsMr7ItK/gm0GSHJYgsDJDsJ4
bvIlJnBw1nwx6nigEY3ewhJovbGCIgP7tnq2H8enAOIpn+1GJhPOJqNjwQY1TAHO
2fTXC8OyVOU4NDK8jy75OCzEtvOj3qMnT3TW8+VrZSXgxyEQDuh3xgwzcW3CKt6w
RAcvOrKNceiYjMdRIDeofj+4+64YfWaEhlCr243RkTEETlLT8z3lOqbKsONDBE2+
WDZB2h7d+xWN7UDCjXLpb2aWkxyxaPPd4o+b7bnBM+6aMnV6dt3OAbzNdjPdvOsp
iHdCuTJhMH7/iEyigsmd/NC4FG7Nzlsric3xznBQj9Vt1T9Zc2Ce6Hp+fgbfR4vW
PkHYWtxHToslPNf4lak5Q1ZIAGOLCg7xanmwW25kr5LI9qF0WgLrU5bYrNlDrs5S
9aKenYZ7RLt3/4GA9w1stOPvMAi8LhW47CJR+4Cjk1m3gqoN+CKYSbwIaKs7iLBu
pBTEL339RQFJ0w7IE4UE5/8gNPNmKyYvgPP8nP5DxZnE1z0rfsI6GNI4uDZ6MHfb
0nlvVk3l9YE+ZLv2gQuwtXMIoX13q7Mt8b3kwSJiAccsf9CoMrrZcELfj71BIjUP
PCqryRBm3RhZRqL25z/8IJknQNlKfA2jJcWYUqQTohxicKoDCfWZYIYvDBKUVAas
4Ps6iAxpLqCTzPSUqZqiDvZtr/S9a3jP7cfCEfo/nEuW8gvDKbDKkghSVm2QYLb7
lpr/dReWcOpUq5cgJQyIgpiemC+CK4sFL3bIrnGlE+c87Y5RfrEpmrvgrVvgTzyp
J0zDY/9UDE06+XTz+rZ5s1xAamHby/6H7xJbyW3rB2XFnFz46dSLcHQlAIzcSjyQ
kI7Vtrg523KsHY7hasf3A8XCdaiZ00dgUiBj3v0D6+a7CU1vERHIXSB3rYYcaoHE
jGa6guzlbhNQhEcnxrWcMjSNWm+Ilm9Ue8vt6w9cgVCr/K12mr12LfdEu2DgbQVZ
Y7ip3mGVQpIIvJ8FmvXCQogcU2JdIR/9uXpam8HkzU4UKURphU8xipxrzo4i8yOl
jIfSLm33Y8YW469GfVOt4q87EDLMuwuvUkJo7+04T8akfsCn66MM/dEsxFPUMudf
bvtjgiQEy/fkvAb76/ry53kMADlr+nmK19DlA7VLJAEi97oS7s25hvYJg5qlGMQ2
D3/ANFP/9lMkb9dDGAhJSw0RF7a20IZokAKTNYkhH7n2R2tchrtXlYF/4TWKCqmi
AO9QvbKM62iFRJUuqhv6XbE9zhdOefziP1OS3zisllmGVmoINh7FOhWCfjJtjwLC
QkBkaHj68szOpequvX71Sai+gaifM/n5kRP+PMNFlAUix33b52JEsMRYsiGrJKsR
QVCxkHCy+ZaSwrM6OQdKeKf62+srGq0YnxLrWtwko29N7VM/A8NLtSwO+dGTIskE
uAIYi4QKRjNsCLoeIvALSaGBWUkwXLCdp17azXFCwaMnuCEmWWfNLOnMBNP+qcyd
zDtEOq+YaBYELUisS79/DKx83chZj5ACzZwWMaa296/1vxueuHfdeWi+Oc8UB08/
XwT8m5wBx8Tn2l/Mc9m2UPr3KW+ObpAMqsVr7BMYAY3IqcSe9OmeJ2Oj3voHzlhn
5cWiG2Gik7ap8MiMZOFP3Nfh/YDCu6HpfeAZxTZJ2PSdUPK/izAiDFqqg2MG3etJ
nH3AeOWzBA9kvjz6+7Dwe4e+ZKVJUM8XOD80SRQMqDw3wv2ZTsLR61BdZH+un1Bh
OldlhrHYb+4AGS6LwhMiRXKMYGSbM9nZ/NfYfA2BswJZcWf2+Di2+YoqzjiGmcgA
WVbpCAomPLCRFYL8vatY1K6ymh0iYicp2FZFBpuKqL+TglSbm2N1yRvumzPmVE2B
y14c9U8ykmdsmow14FtSoy5sU5BLjaCBCxvr3GqW5zkjONbHfNeExdAIENiIyHrK
yQaJYAG+cJQEvTTxcxUP/p6bCZ6ZAGjsbbIqTI3jyMUU66LicjiGDIaFlHi2k5sr
DNCqV7ldRAtPk1o9flXaTHjdAX66WfBqX/EvCNExFRmjIK3Lchq8yZrrnfeFkzgd
oamm+0idWqCKIMquyrb2wf9fPGGGogmJgym5tNLwFIZAfsORmEBDeqHG/2W4AXx8
cd3c6Kc74DhLbjifZB8SspufNYUfuam0r+f7Ezy96vBuGHqX/X+eyY22P9J248Y4
XAe4mN+eHns8/UunNMSQgiQq/oqMiDDOaTefEwqZ72hmstdRKWyDiBp4MQGAmw9r
DFkllAcbhyXvGyVtl9/S0caeXe8f1V8zpLzdyY5pBcZ9edD00uR13WRVLpZ0/0E8
hY2DT6vzfOXGrl+VuKfgLXn6+kdLZqbxy08LFdWWHktquY8/y4X+gatA5C3dKl0j
yoGJlW3tNxYuPi2bYtSqIXjLdbVbuMptDklCkf2n3x7kLxKEdDVGiN2yYWEbtp6F
sNszXNxWl3YLvfPFqkffkXgSok8wF/kQgHrJb2+y8K1T+cvbVQ4rchCkMNEiA/wP
/wxnnJx06li16enK3jyn6GUQWe2endtnbL0jidd0o0bOyYwWwy7YFc1Lg8jvYtUU
oPGaPOmkoSv4+chRmWerwHawcUWA3RLedep9TnIF+7NlUFLFY9TQzE/3MDNH5E0m
amny/OT8Azo0X1TmWdRWcAXEPOY2QYed3N1BpcEDbNN3yHIDJ0DdCeqOEvLbe/0M
X5Nmzmwi9SIGCBYsIP4/9SqkevDEzhnJYIVhGeZnLsUbf9YeXXD8edgwgIv2oqOC
Md24Fsbd39yP6dRXL3dLbY/FhI293AF3SOZMwQPCyJVhWuz1E7mNu0FEXYajPqYK
wEuHi/I/E36UNbKyKLL/EsaHfpuMUAWx+VbGwRYypqUcrVIw3/zxRoeGQ0uTW3JB
Al2dz4UeXoHzwX7SpsHwGCuIy0s0TaoE/TbL+VVNqAvaMrN7pDttfud/OBphlzee
FAxzIIQXyBAFhzFOmeSaMakTjGEVyIziTT4X0c5139QFK7aVAQrpa33HGnjagW2W
eCgfkVCGDbOmJAvHR+DmiQXC1Imrq2wD9THa25Z+XguOHgu+vTBp+RT1OZUR8BX5
D4lk8W7aiwkg+o4N38ihGzDUDL6So6N9oF4LwvC+9Twuqy9gUAbFOO7jf6+xOrha
XVnZgSvM7m3DlDNliwKUQhYoJk4eTxP5lG0tIif6qqhqk3ko4HaKtc827QS9ybyS
tG6MnOCNNFxk7xzSSA0TK12OXkJ5oVSirHjpfFe4AiXSXAsDAqPplxEbflMM2FPC
PQk/7iiBwG0rjuw+BriCEnzIsuxiLxjq3Ia7Zo8xzvqAF3Jr23fX3Di5AGSBVWAj
dlpy28aeErd3IFiBG64owQW54T3toiD3ZbseWELerhKvcnyd1AGFYYbhb9qYHShi
pYHH6r3Ri3qP08bVx6Y28/IyhxZFjP2xGTpMI4tiMYCd4c2HM4b7Vzh8sJytHrCm
mXYL2aueY9TPFw/QrcdwxerBqRrpx5vPh6dKdeojg/FzfWuIOS3p+MHPm/Dvmsj3
FIuMDvNR/dAfgAXoiBY+tGOCdu+vDmikf4xscNb9erCrdHK3FFy6YPO16cbbzGzs
TCI3rew5XKxeFktTv78XrZj/HdKHHERZzRj8cidEedMiI0LbiEf2jkOyxi6fmL7h
iTHeCSKX6kyAVeRyJpk+s9aZKCM0O9GEFR1O9u2PvIYjGdOE6TVSjBL+BoUNkovn
RqpODPxTdB9PXzndPKPYEKhSJAWUXiq/ys1iWyGi1Qrc6ultfiy7REWwFOPGaGZq
E4yEIDbHXppVZlR4YEJOtNfKHYKHFz1je2VSCxUSUi3tNzmxVChGTxZB/roHFGYD
rGfTEXNPHcfnuhVdmms2qilqCLlTSJs8osUca0KQCn8DpkPEfY7b9QVC6UJmmaXE
inBrqY9jxXxDpR308Pk9AuP2kwfsWLEm262KTTr/2F0p/QATnUG0ggRciUs/w8nI
zMHaj6YNd71dLC391vLc4gc2CjNIJGHfMv7eFOJfny/Sf7Ms3bI2JEsaeBThzOzY
DRNTmb5wlNeQAsNwvNvCx93FGeDtt9m9ZpaZOODU/XudzJ7AOq3u01KzFPoU/Ytt
f7+FjmZgib+xK+EUmEC9owiz61occEF9dG7K/bugogplXxgTCZG4DH75JaqEzKGs
YLTsun3PFJWxCquiZYCBmaZ7BYm/oL8ZGEpTUNaLH/CpQ7uS7tiB5XgtMnn3pXdY
KmuVgd+NLYqQXulfTB5878FDbbCaWPxLXuehjPXyLxtkiQSpLbMNIUilRyQcBSnz
lnBn1PH0psKr3nHYKOnWneZUYQT52TOMW3Opn18fHB8fhPkmTb0ImxwVPthWQDFg
XZZ42Su+SZV1imMZPSVuUbCf5FzLd7K0U1JBHa0d4MplrqtLSQ/hD6GuVRPoJYAI
nnDkaaW0gk3GbacNaQogNupCXx6rSzOweB1S3nfKsbHfMaAAc5H+Rlhzo5D3zsgk
cXTheI5ko084jGs/8bYClfADpao8oP+oYslaPPu1/cP4Dy+SVg9GS+bGv0gcvOxb
+sZYmkVC0+/Tk0SHIYVSlBb3920HFvN1sGiV0ZdZPAOIJxexXe1CMWb1YN2nz3Yf
mrlqGD3bVZmg3ZUy65V8v+iWSiDf+hQyI75AfebqCipeQqcR9AAzdviwmMEQEE6/
/lVBHiot11MCKL0sQ9ZXx09C9OnadZZDPALbOfigLjlt7m539VtJwU3IaRqiTNcx
/OM4Y20v5FfUXrhFnR1eWAlL4ZS6vedSVBfg6o0/BZKmZ16VWqlrrCvlcXoqfLro
/+RqYJOPkh2PIc20AxMwMNTOUhpmL5ZHKQGqfk+Yn9ccpCek07NqcfsdwZBLITQp
Q61erpqjEprzF8MUiA6wZyBVJX95orzj9kFbDjwq/4BcRyMNU+13yRnAxSpr2uXR
jF10sgOA++GOT4UlEQ6eb0FyzGJ1icaQJm1ViKffttriGCyk+ebWhIwPNk1kKYcb
9kuEywpuozwogpMpRYIqHiWtgMcymmyv/1jDwPhj68oG6Lgt6BAXIf9RYXynInER
COHXjalCevNEuT1clv+XTS4I9SArKZXKmaLUdfaL5NufpNFWtOIGvlWTF1f4S0YU
4I1FKMJXFqh9wVTaNw+5VnvYKEs4ucDNQUQlOdFMPJTQfkiPjq4hmmI8o//pepCD
RLmiUB44jaETpD41M4sDWnZyTd8fiM2Yj8gbsjy4VkUUXjEbwUsijHZe4ZC2W/1f
xAWOEkdlV9olTHCEV6xD1HyPVN/uiZPG/zBNJJbtpYnRdzcHxysJ+9bxbAOlil7/
GZjUPfALt0MF41xexL3m+xN8fO/yyTnDdk5YsPeXbJ24hls7tOt7VBFtpay4G3c1
SCP/2W5FiH/zMx9T57bveq/j7Hl0MXuDZW9aYKZb5o2MxPxnBJ4K1GtjXYwabwGZ
jQD4DrgOS/2aa7C9hwEtEXGVQMc7rvB5z1KBPqgobU/9t+Q5ryenFgwEsyEuzvWu
veKioouv3ABD5FRj07FkMtJzwxvY1+J+eflvL0yTv63AxgA9Mz04MFaF/GabLHV9
cdci8/7k1GmI6399cDoF4GVDnHobnq4IAaLDtOoFZ/Im89TbqUy0zKU2JBlFeWbO
AbJzs0io0mLRdvDK/lX8JDvno2AjBFAw8CtUUtpFgkbXGHE/poPtg2cmLJTfKkRD
5aeb7xep9QDthrtc74wVPSJbhQFLA7AeDKLfD4ysCK3Z3z3xKio3UIERLkPEMC+k
UZrh1B2xb6egBObjc8Z9+mr+PnWGZFB1R2xaZ2cUJ4fdcx60Y1PBJsq+GStg0OLA
yEGj5ALeIt3R0/bDZEQ8feMH4w0QH/9Sg8VGSyRlYFYerzoZvvjEtTFXvjowZLla
RjNp/TPpudFbA/V9gI3Ns0VE5SNqY6IX+GsIXARYUOhD2uz4sFjKy3yDZZyTQXvk
Egg8HT7W6PAVt11hdA0jH7+FQVJXGuBsJUgTypbaxvTxDPQncZ55BPiPGS/3uezR
+rYcIoYjtG4o2ipSdN4UlNP99nMABflE+QatPGOxAi4YyJkshPfV4v42wtdPKsth
w2H42F7WCOSaB29FwVTHTkUp/jDsCnfr8ELYlXTgtxhEA17RlALAvWfRSQjj473X
tyTjpmomFP7PEN5Be2npBRGRnoBNcLQe7FTYAnjnLbfHPMQ9t21lQxvP/+O2VYf1
4wb9r+QyO+FaKQ1fllVmojMegrwN3jDJ80yuAOpA66DvlQQOg6cUlfS2ewfuzR5d
zF6872aMR/5VS3cKYbJWzdAqzLDedz1bAWqsBzJdufmF/xS00fybuQnhgRvtyFm0
Uo9sEKxw0lBc89NMFXLnmtzwS2Smj47d7FDf0VKCHdHT8SqiDhlFqNJO1ohr2+vr
SHzLJpwmvsQaiwk84O/adnM6RTgu6enizeEWHPFKA/ChpdkJOqO1r/GWNDj1LNvf
Wxn7X9+OydknB/DUfkiP/7QrNHIz+ljHu/tuNepo0Tz7xkW0SpGo7lx55DX8Dw8L
p8LZKx5BsXEVMerAaoTxcG4OLD7M0gLyOSTKjkqAQ1x3Z0ejhhTmzvcGyE47J+I0
AFg6Ce147xONDpggHHE09gOPAP8HwJ++33uZjtvJAtyuJoMAMXgDGNlN9mTYarlb
T88rA2RvLNNB2tRn+vQxq9aoj0ZPB6NbOypcsmwkzzTbzd7EmY88S8apkcOOb4os
IoCMJsI37nvcFid5qeP914ram0o5FlXgJl/1p0KTkEsl0891AlADtHBLexForq49
FV3fEJ7k9f+sZA0ie6136qtKv6JQ2fLObU+z3EEMZVPLq7fGKK+SLI1hkeqf48k2
iK6Eqw9EWxtV2ZxL784xAZ1OWsvkkEYrjfTTT6Dk8WMvnGlYvTPA1sW4QAWuEaAf
Z61oeareehl4he1eIpWCeKm5eppAXya3Tir/hXKpE/AgI0oVnqt3dJTQR2mjRU8i
TjTGAzl0ZAaTrVbKBWLL4Hs7zZJod+VI+ch9/ZR9C05aCwGZpDGuZWfeIkLFm5uw
QWJ2ZLNb6xSeDY9I/k7kcbQI+YDBvk/R76WRuO2I2lbvBVzZjGXBKh4Fs287fc4n
Dlc5MaBmR6pcHo3SkO4l/93teZaxjQvjuTICY8yn0utOJQmEqmQjxlfYT7NqkdT9
DvyXRV4Qodz6sWIrGhMR2CAndRWpjboEwaUUc4FruZ+suOlqdENgETpMYdhW8uRj
mhU6ij6+OGOHjd5ruAmbfZBEI245TCD7NOnc7lY8L4/xIzo8uTpK2utxjm3wg29T
jPeJ0eVWwNwfEdc2SeRHw7S/zCoOqLBGmdajVMRVScaknvLIErCQksfmnUL5CuHY
o4K/+ADm2nZ/qpLYtijMboxRAR9udQQNw7nsaXpMBz3qDw5d4jPhDftN4pCYR0pI
DRLhSzHdaE5WrjDWE81CpLYE7w+Wq3uKuJa5GpmVpIr6nq7H0G8wLnabt45h+mUo
vR053hy0tJ5UHlWGKy7qnrEGfmzlq68rkMavz6kpxo23PYZ5fY8c3Wa97OIUPwO4
B8o53XL9C7K5QNIcIS8n6DVuAiGnopUCoX21ZTGab3noGB5bZPaPFZLlStsCgJCs
dqKrTAYWofdaBvxmQrMB/w4cFgSrDGSgPqVEIvL6edNIsH0x+GFumBoz3JMY4Jdl
NXKn8IpAehkxcuDMfRRVaXHada62/GghcPX+F7UHVnXW47WyLztiD71CUBSMInkk
Sa1HVoKePKgt11NvMkwSYuvDDns8gpHbDTviieibmDkCEl/GVKKUIllo8y4qhiql
TcmuX8rflz5jre6K6u32Qf90RL8KE4vLG+axV0Z1asu+rcbj1kKZLTG292X3wq/X
SqNuqUIIQDEdyhHNXT9x+idpdb4HVvRs8DZwfRx7Gh1W4lhuai5oI0anlOBGzOSi
6XuXFzF0E6+b8ApTZU25EUbWLtPa0JlVJOBqIshhfRB3Y1yMHWCwbyJ5GjDs3YGl
X6J9UEgbxNuAaORcETsvhDCRmJUPMt5dcHmhJIkq6FStosWnEjROgRNu8lbw07fR
7mgV3OS2bi6DHQnfwr10jqaRlSU26m9riH/BIQPH/FercOiSaPq5wHSGMzn0G2an
zeT2qotiVE7G+i9x98aZqt3MS6pPs0Oy7Qe37fVE74FO1sQK6ZQV66ue/Xbpwsi7
8O/DkWAeKY0c0Sm3xoWEngB9Pn8PDQQllKOqMT+8srmulFWionZ5VoR4LBIEtMX0
2W1q3aYsCwohZKtVCrph6mXj5IThws/pIzsMbeML8brqOpV+ifn2HBPYtHOpqU/4
3kR5kmVh/WZIIuxg9ATavo6WdjqqGwYCdkd2nRWGOBMUvhSXTt6dJbJ8z9tUH/j4
s6jE9JMYMMBJPSqA+lHKRkYli5ohrG+aT0KxweGTRZrAltb+05NZG+axzbHHkQmu
F1TVsB/JvqPo9xpvT276DicGz8HapBsd0dOpKY6euEF2gEiMUqEjnsDma/v0SIrD
VId+R7rNZq7x/fa45w6b2TFAXa5klYm+8RgAWUlCNPJEPqpUaNVxmR01zb0JpVbI
lBOENcUoJ/ENWKtH7Nb61ES0GNTNjYS8s+1/FmKFkF6r+B/MIp54Mw3tXKaazP2L
wb3t/xwDVFxHGrrpezbnGPwOdfq9/pEGiMWjzFZCQcwOPkXt54NstREngTXF1mxf
bpkBPOZGxvihYekTAOos/3wtq6c9zKOqlwcLZ1aVoPco5rRCuGF7iQS5r4cVQFdE
AImdqrb96MelaDi0H+UXu1xCboEhzp8z52w1wsT8N4O5d5L1PNt7exf7CY/AT7Zn
0w1IOOWmKSWaIXkpVHMMhWfZjeMwPXr/jo6Lv9GFzeIuBWtJIeWqUCBdNB/OlmdP
UKZzvOjAm0xfcopkl6ZXofg1eQFLZn/hfRXy8p0kvAk2fz+2O8m23jp+qf7na+b2
2Md9HBinFe2D9RkF3T1Q5DhSBL4qAA/pToDyDb1ejvMllwlXHMNRzH3bltz6+Ran
HMZs2YIHEKINRcHsQxPXj5Of/Mx3XFSpSWGzHOSjzrmTs+aiVLJHPq+W9lDNAXAC
S4f+P63tArbV6awzRZRkq6laQ89kFaiyQtXR7lCnaVUbgGft1f4zo81R4bEVGGHl
LAJJF4d7Dpw+FEMYtB/5Eb1WiqIh4E35LtInB8CuZkUZEJvpJKZjxEg/SZIb9Bz9
hpwHY/6URRI0QE+Py+1jiEVyx1cICj8H3Qho8rZwV0k7VWKjpSEvjAuY8Xj4xzhG
ObbKtqrZweCLlaTS+D29mGYVC1Mi/QDAfwPmJ4Y/K8b4XcSoq2/7f0meL7MnYUWi
CEYmQdJHylf0YanQiUFtQt9I1Sivf27PiV52r3UEpLG8cUuJX+QuiMHnMnrMBQUB
SSm/3WOeF4a8FvlGNz/FhziHlIMaQMiJerSxIHRf3bbXVBNNRAWpx1YhdH7o/iPW
3UOdo1XlNJVBVcPjzPIPp+LQ/7rRBN3sFR4pPIBSDq5CmS0vFq4ToGFumDOHbwBO
Of4wcTt8DRRFTN8/5+VLrrG68bsDUmjx4NevN/++7UyBASyHyzapFSpgLm7a6TX9
FrVOm0C407Jo+tOrli/NVK5DwLFx6RLTPMunp0gw0oSzG3gSrdfi3dIwDzQhdsmC
PFouRz/xFxtgEXkG58eRDbFrF/6GDrVGdryAsfv4LELfrHzDzsT8dgOwlqS8FVGu
gGOdmZnmYnn+I1OuYIUgR1RzBS36lxHVrlTqosa2Mk8UmEW26x0D+F39v17G7GME
V7qtgfQ1zp0A4m0zVuTlom4DhmY8xYk7wxPKCOicPP5AAwPoJMooASJD/3T43VdM
3V2NxUoTLzbYfsXYbYe+8OSzQt9koYgQWWDSj9ZDQAzTJprDuEFcSsa5WDaKXaAw
bDDGIV82Qa2ReBAIe7GnWyLBeGgVM/MDFfKfoDAABF7lYzMFYifJOeeXg/Dorl8V
ejyvFupfHgDXbzQ6a4Q+YYOegS5FcJLQZvX9DqncENFXTyoQouf+cM0P3UUzeWcd
t0YhrB2cn/pQpzyyOU5ffBOq0HAFLMBsg2lum40wsUtf84oMdFqGQrHKivmZtqbE
AglyitNdkNhr+WzUwuzdx7KcN5qbXlarkIQBCgm5MSTIvf5pdnvSMFBL/OoOt1R/
ARMXXtH7GQ4omRcoZl4ZPRA+JP6ADqJ+AreK/aLFhpi12Q26lWzwocjR90wR1qTT
QyoUMPQdaa3mDaN+Yx+J9L4jyWfflD92J49djAaAU2FbqYpwLWSL9PNFuGaxqBQ5
BpcmnoV3grtgYGxqQb6gD3+CRVfkeA0IenrKOzfWxk3JVy6lGcn8W6n2RRIMXptt
fPwO+JhDDqSgd9qXenc3MRSvv9NCrtHVqaOiZgU8es4E0p6ujkQd9ww8miZRecch
zR9RX7E9sAac40a5zRQFdqIKqnKlX1khwdhxgoDN3uGvx2cayxmq8+baUt70omkD
PI/Pd+KIKT70MJDfmtjoApzuA6F/NckwUy2HObi7WbldUvp0d1nGqEfukCoDAX/t
YFWeli0TIQ+KrW3Mhf/2AR2RAwsATxp3tWBDSeuBBsGMGe2a0GA/VlaFjhhI5OnV
YJQ4PgL7cy4ROsZSHiFsaStSPo71Wq5giAjpG30HguGaWoyaP8lMjTHyp5Vqe29z
dVMg7MPeRVNOgscRT7aPfIgSmVRY+6GvUW2AyYcp1qQvFqKF/TWYUoOYZOYGkTzg
2mp6DOPYdRYN8rz5TV4nD+6HxkhEZVeo9YKwd9PIOP2233fDKUOIKQE0ydKF9TSv
xqN0cCbc2lzAG3t6Ewx4aJQirDdnaSHpl7Ponds0jX1r39nFpi/p4gcLtJE65uSd
IsvFGeNUcp1t6VPxIBF2C2GnI3T4tzoJCmjTcvbjMkUS7fkNDaFc5cU0/fQzWicL
NJCfReNml/XTIA/bUTIFF46WMc02dGTTr2PA0laynvWRo5B0+vGDlgOoX/wVPNcF
jhrbU/ZfJ+oRSL8FGVzkI/uOeKxc7Vk+YUo4vLBhql48MFHBASU0n2mWnfWBREcp
b2QmfXMN5Q8fYxx578FHc3hT9cN8gwl1przfY3EjaWMv5an7zT0aPMapU8eDwR0e
3HJfzzrRB8hbXxHyNadL41LtTxvS3tgackCAiJpLsh0KW8DoR+qnRWFyy9gjvAWK
BunvPlP4qo/7ufhZWcHtpp2tsEYA/KbPNLJduJ562ywNTOWiKVG//EMwszeESNqJ
qaqqKJP8eqc0sSFHt0QmNENYS5zX6g7cdLCToPEHJQXwf2PiZ08pA0GMlUh64qmD
cQkXJ3OzzQAI4n2lOFruCwPRba3o3R2Z/2eq2CtA37dzndvn/myIs1cdzVsnGmou
9D2hyLVEKVRYuAHmrF1LSjXHkYy0z8EK9WGAAcK10npVpAW8SUy+5PEvXlKi9ISz
Q4X65WcTkVlCJtYBRYi7nXnl9uHvxGL2p56dB2Yepe2WT1EVZCHKieTSRetQYqid
CnAptMGh+K1G1yIQP3xJmRsOZZJdjvWwfY1wYZwZN/Y8+p+RH0atSX3+Qp+CMCEC
s1DCFcZq4L/XUpW3+blw1LQn1B555d6V0O8PR/4QkxVuxMYeP9NTgpE5bT6tzuXj
YoTap5Wk6wypTpOB7wvHi3BKiPzld+NbT04PHiBUZLqXzZ0k1RmUgdl4INQZaH71
z5JESbvE7WOMapRzLg+z4ToIdvbUFFrXw5kJm7kQNBQbDuz9Te2GAyszT783MwGW
BdIa/mt4M3pCiDo//PDvx0TE+kJPxjfbYNeWP3tZlpTcxcarByczFP6zm7L+zYhE
GB4hiq8OmpP7bDs8dYPbOdrsTxbO88ZX1rOhG2YLOuW5cyxykrMyNBmdqxgQD4iW
8P+9L5tGU4oUeQDzGhevDJwXz4et7J+iWHchzHNW4BJ9rJHQgeqqMI2u+Sa4R72h
x171nAxyyEtmzy4vcVcOlcx1nOOpl5eHyku3okz4Y9mdKEBsfXnDtqqPExr5DDGs
Pt+3Igr4kAjgwqVE58N967gijAFcacazXDDcviwITiMxyjx1FWgUSSYb7JVcinje
sNGab+lFY3Q7a3iFBO1+TbqZwPpFwZeXNfKxi8RVyWKppn1OeIyff8+PXUAN/ZIa
97XmQh8J5muqSUFxUERrJEoaO5VYixGQMkk2aSfc4OHjZ4r8w2v8OCzTEwfs3U1z
RCJ9B7UjLjyVqEnCBfPmugchjmI1xx2nJlGT5CdmjmFdc+oF7NsEafjgLmxB7HHF
N6Wo9eWNhHsPmw18AdHC2EtcMgXYKWDXwi+oNErtVW2zupNU7Ae3GjqOHa3ZSXop
3OM0eBBqDCOXjtOMHph27AwCAMPgXLCuDk23tI/+dTRf9YYH6gbHLT0KIIbntiLO
1JaEQkOFq8RfEGqzzBgeHvJVIDz1jAWWfB18/Lb08KtiGZceVESl4rNuLEk8i6A5
WPpyU3WS1Qj8PvGpA9Wmv/doHDkRQ5hA2lC02DUvdM1t7yxDJnZC2pjuwmCzpYAm
MwBMHqOtMkRU8e4n+1Alr2ZWXzPh+4kGgS08UCEcS9CjaK3saoqDzOqLM2V+2v11
2QpO6Sv8I5zlZs8FvwkeAudLtCWFScVcRi/3VjKUumiF/DmxHnpaQzzCmbSEkFRq
s0Mq4c602ZQjvnA7GqoxTT1tq2UUPPnKUb0nCMg5BtEDghIrLW01W6Hu3Sa1SMeJ
m7rv2sFLTTakeM3uE0+rZ4cN+m8wpxq4TBZnr9oWQq9zb6d9BjLyHV+lrxNHBlvQ
batWkPZRXtIl78TWgVwH0B8CC3E1KMLzKONhhAL5MEYHCGUkndOWVWFk9lGFZWzH
o8kQpb8VzjOtou3hRnjnOr6QZIBZbPGBhham2Iqbk+aqudHrkjMCMozO7pZy+Lc1
g1TxmE8qg6WVC3GpvcOUrT1SjJH5QgruVwxYsD61zkP3IgzBbTCTTUJqfKy5kZ9w
9Hi+VW2c6wyjCAmGUiUJrs1Wh71WHOmQGtwDczOjGokMLWZJ+9FjzNokg3o4T8Ho
Emb/w5Y1SGaS9TEs3fSjb+IcHz8mRS9ozbb2vnBlGm/m9JBzJkmEbkwKFruRV/qB
4ayi0UhRt11nF9NEzWKoopXat1+2V5Ympj+T8eMqmy72WM4ijNTEX+x2E/KGks3B
six0ZkqK/ONy/hxWmI5loRyETMd4eozN/aQgpnV8MA4jVOIIE7o6nfOSowbmg3i9
h2XC60sPARvkpoL3Fb2xaYQkonA3PKyIoJPS2lXl+mAoqo0qslTQLQhAqYHyuvd7
p/+CqGDfT+GTvRTrgvRmxuLUoCX0vfRCHZEMkzpYStHLevPG+JO1+aUmJ5irkzAx
e5Cj0YDhlE0Yn6C+2WPntBUB2weZUy/rV8HNPnTuMrcDe/JpCJLbxcPhwe3fKzTa
g93nHHkLPOesofIIMERZixbjk4SYe7H7CAeHq9Tzv2HfI2Wx0bk4sHjqL8AT+SFd
cHJc2PEaSv5gZ1SGNZdXwT4hsWT0vQZHkF664eBTtu6m9Pl5QdeWLFZf0wqrFVwY
w3N8irFDurHfFQYmRZgiUgPcsesgo+RfScM4AtUe4iTIOzFqwcupooDUDG775Whl
HItnoyXZL+GOkR3W7y43hlvn5W4GsYG8O2mtIWeDiKGOTAysYo397Q8khLuXjeVX
bMZLVvzzY2H/7aZeod7FvGQheNq1NsOGZ/ipvRS8PaaV+y3jMFUj8XYLNijtuSov
JI+0jbcYSJGIyltYiv6303q6Kegv9csmfHMOFLbG/EPwzYNCMjomdIXv1qI4fu4Y
7SjL9fZNm4piBJ/l4Qa1mh38G5gLyGAczquWbhOzOd6o02+woaKTYEoOGRwyYwqA
SnO6mm+DMk4gRdFWYZYKYsPIatI9j4unFKOi4ZBvQLvYOcB+8yM1AOX4X2BD/Qyp
ThEz1AbBcXeVFv9LRWMA8EnFInuuedBUY4P3gbvIlc5BTA0eyE6AAavpAKiwgUU4
DtUhT5gFWD1l0TJbzLjpHxMlv0+xIoPrkNOE7yhid+r4FN6o89f9jG9/HTFHIT+C
Ll3rmfKrVDnT2MSvIBTx38xSoyCGrjrRNQ3UFRqEO0j/FsDeKU46H7NajbrQmDyH
9H2VEiaBlUNAfnX6sA01y8IbnAMDw93gNE1LqQpod5LSlLRTF4W2n7WI6lafD4vV
PCHDjb6BE3oeUlRc909PC9NUIWG1DSoV0j+mUuaEjtCUKvwGkRytK6jRMIKr0XLa
zXEtaclqeaBYo4hsfoDomX+AmpqgU8IDo0XHXmtE0q9jNymtUdKY5Dha1Ms+PoqQ
5bt98irdSQtefMCyHy8qqexRNIHrMcwjwLw4pQXoCVvx9oQratiMPiaWNNSp8FC9
F5m8n/vAEvjsy7i9TDISt0l4CKx5+0NIQt/H6GWk4odsZUt6oNQGAk8ys8wMngBc
ORqG5raAlO8JGmJg7ajW9fDaYTjFEQkqj1Lay+EPeNJ3XTqftTMJdiGIZl2W1tD3
bkk88R55cD62j5xxDmYh8QdPq3bxk2m//upKur6sY/Rnos+9RpnIwW3WSZ5OmdW8
x6rhWs8/C9po0Z4+t6k1Xbxomifl8v6BVc19KqLV4/s/DIX/tUYYgue1gDdAKgIU
Xzi9uTQqQsyoPLWHMWGANwGjT1HsmctQIbg+3zCapl2DlFXKsKZyUMhmajDvKGYJ
/tMj3SEpgI2Io/yY5BnNvMybwHnGdfh6BfC6D7+JG52Q68/6+ibSQ1lF8+pPcKWX
ssfM+07LUvp9BG8LMw/uhfYGHxTdVCggsW2A6v4CgEV5dSqgvzNtOgm9lHxAt3WS
iNzkrHdzeGaMTQJHipSFX4Y7uoFU7oCevVcDnDDClb5izQG9ZHKGCsBho3Nm9C3Q
8/bcPMaopbPmHN27CgB3lrWz8ZHDBDPv9MrC551G9/m5YuJorlV0hH9KUpl4zqXq
6UYlDEOykwGD0oaFHgWMvo4Hw/B/+fQoZtotdIgCv1YRy2l2HWuN2lkBfyq2BcY4
5GPGHRygW9n0crOhoWi8IVJRD1YRX28GUBX5uxkLFxckh7TFxlQliOSRGxfyJMF5
U4fml2o/JPGv+OsmjdU2SgSZo35ExOXFGx1i3AFHgXB/yfyyeQGvZSTjQnisSq2Z
ID/KtMBYzx/SCG6y1zwWgnHyjVKgk1jIGzxsMWzDvqc/TXhbm5+M8AP5clTAp0QK
GdcN43q8f0lvNz9W0EhluD+vKv+W/tdsXkAAzFZHz4sWhPbf54fzQB4dsia9gWMT
mUj/w7PGQjobEYOPxcV/z4fI5EdI0fv1CZk/p+YZ3j0GLaVYOOvqS4pmy3sbFrqX
B9Qh6QPRVLZf2WGcSM0FJq0dwpkyqcoqXc9UYAzyfyOlZHSsMSIDuRBDW/iKALwy
1oOe+wexkTJ//xVnkPHWl7eHcbiFTQ5CmKvIc0GC4wYMISiFMEmWJVtgOrCgYj7S
vyUQtmN3Mi5+JRQMr1/9O7EMl0pJtBundf8kZ6WUTviNcvShggFpjQr4bT/rdXYB
uoQ4UkBnmpFWhZ8VtcGg7pOuBo8YUd6sAdo3NElUvlENuHsnKSSHfHHQfomKYnDb
tLb65G7DXZ5rQ4/LouAt6pN9xToWjeZjnAMM/z2jUS69yNa9qY6uBvgnR9Hg7P+F
8OEL6q4fyKTFyFe5Kd81zyF5a+/TPSChQpeHrLMuZqCHn5Ng0J7lVoCsr6fI2DTV
DMAYHytpYtyjFNw4UvwICO/HhtOekmhGW/PHY34QU9Nb7pOuNhlr42kzoVCNUPpz
Kvuas+qMm4HTUJCUOB4HDDFV3MNS/14qnDlGjwkLUp39jlXEpdpGCPCV5YUMynzM
E8oy0l8LHh56T8ydDhF2NgolQHQ+rnqMyvUdn6we8GAiJrNrMT6iecdRm7x5rE/1
zZlqkha2QfWpplrAClslaV37XmH2nyiyCiGXEPBEKqEp2h22t4Ku8g/ZkQuKPypF
d9+pMs0ny90u9JMeQXSNDNQj8JpV7yu4zIEhw52nXeZ6dQFeuORrwbzIq83xWxZz
oyhSJPn9sVyIwAYRO+K6I27lMId0MoUulbegE2YizGjOzJQoyqDmGPgY4eyRr++o
an0AKlgjA3UK4P/J83G3+HsETQrSto5dOXj2TT9dpZI6VR0ipH/4KkhWDojJmCq6
zIvc8GUNd2RpyNYtn/6bEhQitnRHSCXPzihNW+TSNFcSNT1+ptpIVegTnBiCK4iB
1NN0s4RKKd2Yney5r2cc5/nunn9Uqlah18reVpz5EmK2O4md6UU5Y/YxYLtzL07i
/QzfpZ10VA6B+253WxpIeCpefvGPrjA2Ax8h0UF8IT9nBZiBig8xtoM+uta/kLJL
87JQsbLQD5W/AMqydw/ZV2X+ITUlTPr+GbD/bfz8FKT7Drz1iogTUZeUejtw7X20
FUNpWUAoQRuIdqAm/rOApdIoN/8cFuO8nCGVbEvCLrH2qyIOAVmwkcxFoeW3ylNk
8vUPnhpPJrsfDJX76hUnno5UjYkyDfE6k6io2OEaFeWF7+civz8MXsQ4eJZth86O
ZMec6/jD2+LENERFJ1aqc0wRZIGpha6wDeF3tDU8ehKiEGfxD96wPoMjDbwRi2W4
gkCbg2AC+dMwsu5Dpiwhw3+YcV3gcEWHMl43W7T+HFENKo/Mk6eNKKO//0lXQ6lA
Vj8KKkzZKhiKI6FvpMTEk3l2Bn1n5u8kjd0cQy9Cqvgn0b+2YpiuQxFzU2MAcQ8s
/1z7YbvrRNByHiHjsQcEDP7OeSPW/6htj1ldCR0WrYvr9/Naj3AUzZqM+7e4VT1I
FJAb3rJPuNNqsywvbOA8Se5I8/GpzNsKcE8TX4Z0ALR+4r0B/wCbe8TwcCa66GKO
oOuSyf2MJ36VpXYtiWvvEVSllb39Viba1HuWW/AzIuqxqEOdkiYzY8l6SHy4B2og
2TKKXUu/GhhkdN7rOd5Og2lzzcZzVumCZmDuwDmKgKd3cZufzUthRsOAY/eGeS5g
9FgL7DEDTNCrOl3+ZarwftqoH6i/lb+BOl4JqnPQjs3iCn1wpNkRqVxMDe/gIRCH
yF3PSRcBDKBnRMTnQRoalTBRcNNCYNO54ZH6cTkM4mzVl4eTNPxs1/zcd1kicY/P
Nrvb+QeEDqbHleYJZUYyenP2CJjL2UgC//m+CH+X8HnXAdn8p/4UarTNqwndNwWZ
K+CUhNQTvCoirOMwOuC/UAulqLC+Ca/WRzpWtBujVT8Qr3pvFlOOABTIB0bmbf6m
KQThmWcQzMU76vZkY+8Tt70dAPucEOQG22p1/24LHv2+Bj66LTpzByRuXr+TK75R
KUsXv8C8Xq3s7/k+zD0ppVGWIOyHXwLXAPPTT2JnxnDuF0rHuOCmvrcIP1a06QZG
ojbR9FZSWShk367uLW3nB98+pSDr/dS4/A7d+mK37UcwgyQHm7BqfIjTqCoUD0F1
3Aq1z7PRHuUblZ8qgbfYRlMvmDhj5xryBcBssUJHmkW5DjEHuUFsKr+RYjaR4HwY
WJb2GT2XyBJVfXIiF+b4hVDU87HSQqjqzOpVc+RAnaGrOeIGKARfnE4c0J3Wf1St
kUVgKgFH0Koch5BlnwxdZa0Br0y6H9We6XD6plhmFokZSoyvf5I/tYazfSZIER3t
Z1D/b4gyRBn1jNMo4h6I6xvAeyisUnwVLKATLJGCrGhTcOT8lY1k1z10ub/NqDuO
vlVlEtLpo1D9b+TP0TMRUgM9miFdyKKYjKcdwc4PS3s5JyQ8l4a7ggBqvOOxFOb2
rV0l8dc2AoLjt0aKPOBHIjz72SU9j9YVufqgZa9RSgReLhDtdvHeIzhEqSZUr1kn
t0uFDpu1u3PxocZM99O/DEJMCqvUGzP/oYXHLHjlNmCIa6Q0hkInIDNbc4vDwjt3
dd7A7A/ftmpBgB5kTsWMo4YoIgYy3qPxF5/GTyq/QnLhAtMsfXpN+OHoPRby/sDZ
Rk4PS7jFa7sxJwPnspvoTfGM4CrC53NTXxw/rMIZW3yUj+kCLhm8XnXH1EUMMeAP
XSKufQDcUkzt4Gyh6yJOXq3J0J+1heSmThCjbealX6wuVO0fyrMq6PQoQFugAWH1
nMf4oRABFwuFzyKX2kyWGnlF53aOfQ/UR/T2SD08CD6Qhg680OydLqPOKSAPIAS4
8YKNlLet+pUxufmGwtx/+m5Rtta5m2tPra2rdtPe7J50hgFP9Shqjvf/943O3Kni
+K/C9fC7YRIoRn3KbL9IBzEHFDmVmNswow6fme3Basj+xn/9dua5stgcmsZ5GuLm
hCfceYwPw+P+0l33y43dEtbQ4L/E0e4noaMWJgaAa0RZsmHwcRcYL1XpS9ZP+jUZ
MKHf8wVGvxdM2FMWI+Hfn47b8B3AF6UmFqpE59jluzoC6muSyUBY5K5f0BsAnASi
PoxTooBPKVMJh2c1+jMhaCLxFOlVmc/fuBMNdi2pbEnYVuzarof1L6EjPlYS2cHt
UploJ/ITlhAU7knzKeabt1s3K/DW0AT4cutNRf8O5YiHG/BOkKdTesW9+39suJlt
4JdWQK3tqoYZe6A66n2rIz/QB6GN9XGpNzY5Xfdo7ihQ+3Wk3YOAarZXYfoe1UAQ
CCUu//fSjbJEb4bQIhN1cNWdcF7WECZTS4nNLqHKiyT8LNDC11zcX5aWnbM0jSyi
djTV+INhdiYYE7QrEdaAuTTgwJm0Oi1yYHQNONgby+hTnolliGDy3IMgUo7GIrQa
wRKQHXopxPjf5R5BiqplwxWPUyQbe0pSnwS8j9uvaDVrQB1LjWhWxPF/kdu0W/E9
YJHi2V7JeYtpUvLUS6yAiZ5766lRFeFN6EAE+7najyoSYj25P16L/OZXHGgfPw5H
S4hDdF33u1x7v3FkbogAnNBmfik+/yPbO0CFF6zv/kIfwSM5YW5bIdlae4AgbTgr
DXmVZjG+eGNRFoohpZUkely7ugsF2g2WA1agZt1Ud+ZDHi6FT3iVruY73b77a6va
bzyPWi4k64OojsOug0x0EPNlCSvmBAU6gNngvo0GTVvgFQjVHagfVDooJruCcgE/
2e1OlsTys/d/THprhA/mGITvG0KtYg3eionDfHA6J2WXhdZP3SmmMsP+yDFMnQns
ljAnAJkDbfIC68yGL6EdFbonb1CcKEqIWt+priv41C4AuEYWL+PDOdbw7bOUseTV
jfdZ9FpVUXHG0Csfv+XB2L6aVM9aJUit9FOZHAoVy8N0MCrXE2mjYWEJd6AD5nQE
mYxfkwx5aKx/80/WSwEW++8hL/EE/OkFE7DSYS1ST0xkutF52oWhfjynJhXDBzaq
O6OpQgESrbZ3qkGhpGMmgF8YYxq9hgcD6ue3MAZFWVWE1kk3BKKsUj2VwZr5EuSO
n1lIGW2Te1Dj2As/WOTkzZW+dgYvAF692vI7BjsN/6n1iRX2DpFxnERxce6EBX1d
wPQ5UN8I5I7pLFXBzi4IffRTXlBrgjhKuEr8lihW8AU7pQjW/wziOLxnqsrrIPoR
sRUrHfKkthEYoughh0kb6K2YIaKjatg+oi/Ipx/pETiaPyHm6NlmgIHZ+jmCJiwi
aLTngvoYbSckY0tuafORTSqqplddrhhGi33uUx+J+NNoJYRM6BKSpT+ruqijlAX1
xr5IFhEopxdLVqtV6pq4IZWWg2pa6/cVyWi8l+9AFSk8FBhcIGQ+yeK86u16IIGH
DOutz3Z2HGCeQmQOi1G5N7pXa9QR4so3STbw/7ffkRf6VdaW2TFOSEtLUbN7Fi/n
X6PXOKmVpDghKB6OLoTd9826auaikD4YWjmgPM2TRBlt+fNMWix/gDvxrYMMZVGR
4pBvq+zf6ChQPVcNW0CV6puNfwreOX6O0iHjZZd53YRKDsLJ1D1uQLSxDZBOuEL5
jVhH+PLQIs9XTsC9L6LCU61nUj3fvx2/HDkDAvDJK+JWifI0eks4ZXu8j8/0Wl7J
7xvJI5LCt8H8Hj9VnJKrjkcobvBbJKdfXwALIeZ3JlqANinL3hnX7RtdwjuQouRM
hETzvOhAx3mLg8WDEfGFXkAJw49b9f6zoo0sh1uEe+xeUu09+o8ltcA89BEDzBhi
98WndtgoxWSW6HZgcXANJ5t3wiABpAobzmMF8SG4gh+G4x0s74yAeseFR7QJIZR7
o5dEN74/MKmRSTYxpy9/YQwvlyiDcHq+Z4rl68/S2z6P83palwp1OZxVrEi4YRwO
rN/xd+FNDbYV7pK4Qt97iXWNaDsr7Eomj7eYkYoDUKAeknvHdnHIdpvg6SmmV+Wf
C1EsKRNRXAL1iFWCooopG+BsAdh3mLYrl07274v8usWIhBNGKS0WXdlWg+A9p9uD
85cz34g0v2pb7Of3vkHObxBMpQysEy6MQlcMNpsVxe+QGUMA/JHRevcwr3A5hPjI
PRxby5eUHLKe7LF/PD1Ok+DWmD29eKtTX4iMrno/BEOrLeSgNG+TsJkd2Nd98wNQ
MUxj2CsQGZJDgXAWR1NF6lStiatq5rSYBFx+q8T94t2mJPZEZJEUkJo57QO5h+Yl
+TYM73k6SVgZ26kAt5Q70bHSP8Do510aHZGhQ0HtF105d1BRCVXHim88e8MOjyWX
uO4z65+rJobDJs8gXPBn2K/vois9Z0kRsz4yp748AD26NAESHbhON5JN21c/Hpdg
46S6iplHCuZCIPza7fcdOqNOgBqNXctqALssnhJIqS2gtBp2GF8koe8WQGqN2fue
UMYXXWRrwTrlupycK2SR3pqcV5JcITJ737aE9LlF82pAzyJBOXQsq226FMRzea1o
v+V+Q8dfBMfQwBV6j4mbO8uhNtLpGqtZtD2VztizWk201s84S2ruHmbHEA9WiWzt
AjGm8gENI4k0cZ8kse+k7ie0AceYIcnJXzvw11haRFeGFq8YUlkvWS/EIWEDNxSM
2M56iYg0CSN3V64HiP9NavCYUL4iOBLlFspjK1UOCqj1a/0fq3PXJMLVDo3kdPJa
b0w7lLUUO6HpBX94HPDQK9X0GNmcNgH2FjosUs/1JVJXgpPOeDbY52TRkmjB3RzL
H4d6KmgA7Un+ZpaPr02IvKjku+DO+x+loSu10DPy5jlOY1Xgx2CWpVsA/geMIvup
uFFZawuDQFR127IfIosfQ9SEVeao2TyPFiLvRnaF2IM4vtt2qi55qi/9BMAtdwK2
u3d9xtMo9lr7zivu8P5/KJThxljUrDWSGQl8k/GwS0lz7Oo2BNtv5n1UexD3fDkD
2yUROz+JwLVrUfz4uK/vXEleMxsBWxeLH8EjV0D/p/0DSBUgxOcAdZetyRvYaWNC
J8koFmnM5Wj6EFqr1pNAOBHvRnJKuOGWZIUPHCF/jPsaMEabMijXCPq/ND3SQinV
kCpHcNDM3XEs4OWsMjYxH6rLy37yV55ZBDbcOvYu9jEfbo9fZRk45Ie6zr5qqy2+
yo5KZAp4vGn87RCN7LdjgDWuNe9l0G3hVkc/CDvEq0CeBLaqNOlqSfwRwq+2rNHa
23bIXjX+ilV4Ii494O7NEjzymMlSpa8AQH992seMveNeNsE8ZZa8yHUwlsTxVa7d
3lrw88aAcNM7Jy7ztfczi6NATHhhuMke9C2fLPuhxG8L4eMwXtVZVwDBx9TJbgY3
QDapoV++Me47uriqPBSrqe/yxFx0FcNE9FfClJVtxHiICsv9Dp1ovpLO3rjh2dT6
L+5rKzQ42Gd+h3QZ7Qatv45k9w45YuKIvGp1mns0MVdejh8/acY8Y2h7E7nQPYf9
pzKtIrfwECLBjxNlRz2i5MYJjoNMwE1l2WqTuj5bMyQPNEIiIAVGibFaVfmJSV0E
32pN5Facg4bkdxcGtSsC8iYFS6c7GDsk9nl2psDZ67BwrQdzo1/5/2vfBWJSNHq5
WxuiVC4Wop9G2A9OIlVH/UCCv+4ZoRsuvfuaXPGXc4KPVm3EZJAhiyw0LOjk4oXP
yPMadt8z4mufOYt/N1QmuJXVEVG1y7vItxF0yr9+UADjXwtph9N9dcvgl/O2uu73
AN566wDuder6GGf3XGjF1G66npKdNIX8aLQAGbdiqXQQr/0SdNwwMaH8xXrQVYYS
rjk2cFYzBvdgukuEkgxgY/xkskip0kOGHEhqYfrB1cF5Hq6lQLD2/B5omGvdbbHy
Lwfv1hTTvvJY7fcSVQQDW4atKYMBpd/On7wslLcpg5mTtQdMQzeF/AJ5i4sReEy3
5trpaImpZcz5aANi2pajQ4p6HG9KrpZHujpBQbK4wBUB7RUWd+HvYoJKoletArW8
D3tQWMMNmMgmcon9U7LuQTwl6LB6j0Wq638K6GemVFsQa5761NSAO0vWlD2Ismel
mX0w3EPBd+ktNisg2ozFJgGOWcYKxsQUsx7+7d5mEaPEGHbJPcUUGvhIU2YDZy9h
hgUN/Hx0CKYGQN7uGTDg68zcjHE2pIVdHX49i4pKv/NoJ1EzI7+n2udEdTrYaftK
jf86OOLoQJPmDG0KTVaW/cXs97vleQGK+wjrelahBoemSfoycL59YvsvW/6RVzQ/
mKW7sgY4TuOXaM4IEGddkvctjG0J83iJOizF4CTHLEBuAle0LL5RljeH8IIdwiC2
SqjM32KtvPdT00Yp8vbw2WeFatAh4Ppf0WDXX/1wjAgRvsBMgfWDATZ8wtdtflKw
2RDs9SG7JDfyEZD9rcZzcJe3tq4Qxj7ipPUoM8uucdVftYaKdY4ikp3p8CTTHnzb
Y/vK5OPsNt8QrJjI6/+LIHWWCquAW7F6S8SB7fX4w0CYSshcpbWKMlPJSoXoxunf
UDHSUjuQpP4MfQvorPYsLAR8CY89e05iXoPGKJxfzPcTQFcJ5TGU8IgP/YUGxJVW
rSvR9xL8iztDWCLurDb1wfgklKmZohUJEeJGf5dr/rcIJ0jPsZbY07Yx1tM0dfau
lfPgDTOGB/2MBEDbAz/66ZerUvzxzeMZQgv4yhuzqZiuDGNdVFjAfkydUYpf4xgl
kZwamakp30Dvbh9fXWQvKys6HMdCvwkhnUz3csdiySanEuP055oJRzRHzsfQFvuT
Y5874P/Cx8rN4yIy7t2xQeDF3JM/04A07C9jjfyXezjPhQgHYi4pGF7atZLRhRZq
0npJl7YsqtpcSv4iFrvLSTnjdF9dcWc0yamw9Gaa30xYLLwrpr7x99U6t5W3QClY
Nrp1BbeYNJ7RlxB4Ozj4FbAJd4yxsVw2GEU9bRMpg1nygIloke7+J8ahYW5zSTxw
Ys2z6n/TCcg6Ag49F4p6gX6UTzpfO9doGMlRFUJVycOlFIpqN7uK/LDLY4o0Mftp
z6C19o2CnX7jH7WcrDfXaRvCQzo9itmBT+RXQWVgXWh64BhhtkKVnShDoYL/RJlF
OgzIfRHCOxDLSNxLZgqAsxhBwdw2iPD9wVwisKN16SsMyV8/zBGuFGoR7/uGnsRz
lvnyMaWLimR7DQU47Mb7r/INnc249wXlj3G7V/1QhZcb3swEf1Lt2D9qznlPZxPi
OaJJxxG2keuYvNX4T6cE3UcxVZZrCtSbZ6O5tMEAuVJmtavpa2ijEp6OoHfO9Ci2
jW2tV8nlLPGypg5z901JI/DisMoDcFLPBJUkkS027SzB5o4G7e/Z1GMRSKjRrzL/
vmrTpUEAgpNS4Ww5+U1709j4AnKd9DMHuY635sBsKufErs0Tvtgv1lreZuAcexyh
VF9zKaaNzP9HzkQsVHaQGf0dfJUwsUItXc9AW7M7DuatmtJlt1KyFn6MvOQeSNyp
EDHizhic05d33pxw9nE7AMvWPy32jap6+xByiD6lNehgyKKmB3/1kbGnH4ANsll8
l5No/tlaXkT/efJLrd0D0dlIJY40OiGlETkdQVToU8G+rdCbvZMasR0FtFIvAIxJ
+/tCxccY+F29ZAZa8CpgF6VrzH/Ngsm8g8Msvm+FJoj8ra1QMP/jEY8kshHLznHv
+98sTDSSit7oiqNaDviRusTOd85nB9RZJ5U32HquikIef2UDpizx8h5QpuFgNiFL
iKwjvQ4wrTS0kbETUqe2c6HzgsoaozmJMmC/eGSnda25d9hx0bYhKopa7GwWX+qV
IVG1QOJHdjBYiy8AmNYWhfjDgTk7ixF8xZW7bxLZldUlOk4q8TsHrxlIDZ4EzB+b
TcipHJoFpsxQNEUpyKU5ikjfb+tdYGsEedkpER0ewZHQze8p2Vujt2zdhK5m/YMz
8+FtF6hpKKfgAzogQutVVCfltMqErq0COICQBoJpfpvCtzsMz0hmhf22zLEjPzbr
TP3xeDwojFBco2ncYHuP9kFjX5t01jFTM+ICrXO6qfN44oT0TB6s/+osEmh83kGj
SkLJjoR8EnJ2nWomeUAZwQXRw0YtILMysZSZ5NguiYn35cWqEOVKRqMahNgiixiW
Wcdoy8KXWDq0NJYhfnVE5Xu3PRUvTs4ALO0PulJd2haQOP7pTP60OhgqXlYirdS8
DhH1dkd4S5YeUuvC1wY4poKsaphnD/4ZAFsX+/yB35luhy7IpadrP45bX1dVYJ24
icwnE/mIDGQxJ3dmtbcSyCej8Sr9g38TMHH3L0TRW4WCP8aypV5csZPvJ/7ac98a
uZlFacMlhiYiZd011MQInQKkBuqYnzcrxvXn0+U0Y7DBWxHv5q3KZMBLM3PMG5fz
zVsRLTVYeZ19kLrA4ANqC4z5gle7luTOJdRbisvXn9MWyvhQNegQlEJ5+1cEEvPH
GGVfOGZ+FpLUftp/J0jS1qxC25lZO5sPtAh/161jej+CW2Tm3ZH5gypPmNaz3aVw
YcV38iEnYX+AIRBigcYyCvU1e6exn02tEBaeFwyuLnxmVQXhiDFNE2BAcUJ202xG
vh5HTsaJ+W4pdUgV819B6mmHNIY15YMDBbaw3Rg0R5MyLeIE15r8xh1HU4ToXcCL
5Y3R0wN1HGzUIlLFPyHc3TQAqVkyEmpzfG6Vah6TX97/47AjAryMkJhiThWZTzik
9S/O7sChZOOYcpFoAdYNkREYVHN5dZcZoqXGwC2j8llehKODlQfHByhsYBT0P4rI
cTFI1RvVMlhUhJijEAg9bXC5obpDeN178H9UJYEIn4OiZ35vH51YDWKv3nVwMLcv
mjm54b7BW7fOkMQU3HuqfqI+kXlAB0uf29I7l/OYwvQhgk37BGuZfp502Fw5WIze
KzYqWENFzGl4xmBSegkFdak5kx6aVs+1dKQEHGTzYOlNWBslSPkwpd1oS+pH9JFL
UmRpgLUUz2OM97kP85sUx9p7BQwOw0nwp4zqVSAtdolBJUdiG9WzFQQdxAYMUOkQ
2KNXU9iWoT18jtmiH8KOaqfFP75mSWH8vIDcPBALfGUId5pFJ3lO71YHjWskxP5C
nIniUGDSwyw88X62R52HwkG6NIK+SR5/nqT/nSKkHyqtgVYEWE4XSogDwhk8+nX8
CoP5Q4Sm8bACQA6gbK1fCEmVq03pCh5naLX0kJIcNIhNZFZ6338KsDdUz9wUfkYW
xSC98bxFchFCBTLMukbJOMdl94IfhdAeSp73bkCyyGiJTeR2weuxPI2qakmoTTl6
NL8Jk+Ds1PXZdwi5/eYwDd8RJNdSEXFotajO9RlPrz2TESiuwC4Yy7jgHyFQExUE
bn3vBMEKptkjISw35a9JeDyA9kSmr34tS/0ODlGy5tAy0Xj+oJyGonU6/kc/HrYE
2++jrU/rcxfX9oxvAi+XAhMZ0Vm58w9W5xP2VfZ7zpGe/odQZC56a+eDyboAw3on
Lwp4ml6bnnK+5vY3MA8sS74r7HxMRFDAAGTbzDflY7G6NEegmYxdi9JP15mdlWfx
P9FDk3soIfFMlbO9Z7+bAnJVEXv75bIucGawQ8i1tgyu89JXKYcGU5Kdr5yi8g0F
0Rv92xB5Mb0U0wV0r4TmYEAA/rzow9MZ0+EXK6Z1lrmpyUxTTQYE8ZX9K7lAbscz
UBSI+1vJ8iZg2b+LFAAG6WluBbQergx6oUN4ik+2y1atqQ6TDRYAxu/wb9TApUCn
YCvJDvbC7eK+IqX8FUJS80oJO1ZpzNTW1vfA7bvHtfazYBKPv+u9B9EfbrYIG6c6
V8GtcgUwU9dsRshldRlKiYIXoWflKqNeWFxdY/mr7b3yj/2kvw0hqItF7U7Wu2Ql
pxV91pN7QrFKRhM1shCICZ5LMXwoSKJnDnFDO6jVUlBNxAf4I/i5CfcCrYVQJ6vq
d2YwufLYi08PNwO0H8/fvzDix4kL4EO2uvwiZ1TRpKjTDm0p4lTCl4GMiBuWWZZc
vVIEv7VWlhUXlhmsNRBcGYHg7jcd9pabA1SyiYBw3fuxmy525U/E9WQ9sBEul936
Oaxk+he42NrHSnyHr67b0+DeL6ou1Lbho9wSIk0TLr3LO2Np0Kp7ou4sLi0OTi70
3cNHsqq0I1QS7SH3czMALvnYNjGgaLr21xH0Z3kOkwFz/+tWYlzonzbv+SftGbxO
yRTXm6r3Whpcdhi/uixqjqdJmr0c8R7wDmDYPwsq375D6hG09kMttXW3qImqkErf
OSGg/LZRUyoVh4EJ/2tKDNvoF+tuk+7WXGxQSqtXG9459ozUt46MTRWKkUYpaNtb
AsTSEHISKh/V6uv8fRUo0n147N3f1Bdv6PxPqJAUJMURVFuWnv5emUXuKiVAubtl
NUOA3O51gtfFteSO2E9pAcG6iJYLLO0s84vj4SOay3FGSEWdY0JUD2Mj9kD+INuq
Y1fElt/+Juf7Ng//TKkgL7AiboJUDJHMAS9kzVe+n6xr/xQXFLJfFOUBb+/hqmA8
5O9IGXHAfli6ZOaY6JJj1dq7scNd/E+puSh7N+NHjXcW7dKQ7jx/XZO3/LllIOei
t06lbCfNHVJOsraP/pjbTwcaBSSUliUsnDA9AncaaK/7jWEFeNTd1fxYbXC6ZbRI
rDurtgAUo99JlE1ADU2dBvJPU7kjvYckIFYPiHhBxmYnCeCF1kUT0jadJsw9/hzI
dd+Fqst4Sytec+gqhO0zvWbZzOT+lxXCuxEnpfHEBnaqsJ3FudtXWQqZ9q9N0Gc+
Rv4W/PGY3INK0HytKJm/E4pjwDE2W54Iae4rC77puhMootUSK+vatRQPow6jCtZu
vChcMpuAxQVmveTzlKARSDmVh08irgZy+25GgnkUNRd4Z52OCPL/PBlvvzkkVxK3
eWXTGjNxGHfg8sLQFNqE8+ntlQzAA3Xo8KiEv+rLqsgQ3ifxfwjjBk34ftfkfnvN
5fDzV5/ur++gYJStbpyHbRJL3Pf70x/Zlp8LBtPpvrgFoeUX5fjzpyVYVCIzHSUn
kE4Se0G+LrVdrLzbDl7V6qlCdcmdYg4/kDwEJXZqTa90PKJs7Lcir6YJ7+1hAyIJ
WAvODjO1lDsJ25JnsuakyvB6B2OPWI7UHRWDjGduPEja3zxi4WByB5zIkeisoWIh
uEHXnTpD9c4WIEy5iz8iTkTFkFZQdx3pTnDa9ezg0g4VsZmnIcXJwrvQw3X2Q5gR
Xs6cNhqKGAHg1UYxCpKUEEcTNhGpeT2Qe3EikHNcLxx8TKg7UQLRI38blWGsuPFi
vaet0OLSJmBdI+TE2cldYDJWrRr2sOjn7HXrusy1SK4MTiBHjvDOSOVSYaD/JaSi
A3g/fh+9UeQSK9He6Shzb9GF720Pmbg0gdOTaJ1J7q0DEI9uZ4ijzwzlkbVae5Cy
Gr2cH5CWNk6giTJX+HBhS7rOOsiysHISvU1Z3uMKd0qNYwUsDeyolUSMkO5jcmD2
TnKTAdEPt7nvPmbkhHR4In5mvVv2osBQa+RzkyNe0ndCCPw5Cl3Q9oztzUw9tcvT
9IZYly/UlHF0ReLR9q6LoisRnyx/xOlgEaLwUuEWHTX4wqQRLzNudpUhL2n8Ajqx
t1HZtDMR44hLaPkNWSSUSgjiUEo66PalXW20/IW57Sw+4qUIG6AXVgkv+cgEZK+n
cjNJTwc3NDucB5VBj+FMIEb800qb3IF7WdB+bnuyWYRYhl2/W5umC59XjVjBg2pV
YDmlsOpiw3ZGJkSrjapgQuzgR4kW7SuztRheMxxCQRgBmFSG9hKsRHs/k0ap3ndx
xFvqdfEKZe9EJMZI1Gprrg7ITNVgSZjw74A77t+fDhneYbh7uM8VL3BPItzi4erd
qR4TGBqA8cOnCps/o8+QozAp9Reatw5tsDV48pCWlkW+RR0MfnB9xG+edDk4zkX/
1DEOOP7ZxxqnFiqJHTvzuqkkqoZAEq74on16ia6gr/wQNSNjvAKpw64Xm999uzP/
vOpZsLi+ziEb85ZH3eLrHIpzsxOU6CGECmHtEzMlVCDZ+542rPnroGFrwoEq5RFb
BZx+RkrWDM/fVfOnRX5Vy0tlEeYVjhXLrNrmsK4Y0ygXsJv9aVvWmmtELjttsM24
dtB2xhjI0CobXMGAgWdxyT96rBRWagsnB3AZ9oQ6Z6OtNQHJZFwUl7iSzbeAJYGg
8DTQloMefvyf8ST4eY/DsJTsjt0uFUA5sxGU048ATEHh+VFsvYPCGVmxJqRSorwm
KnscQ07/zypicEYl1ymUvt3AvR0P7Cg/oXrehBZJS4oTGBKGaKSMOJubjv0RNGbx
7AYiFD7Js+eVrCCshgpOgwONfH9X4rDkkT3xrzddWVHkfBIzcLq2CXJDaMJ8u25w
nsPfnXK7I0lXlwrf3Zano+nX9541/ivyZP6ajBisMdq/UWESEk5mVxUtdOcSAUx4
TbAQFYfkCP1CYxgleRho/hE8Ym+rTSEmRGQMmONU1IU4IEQzsK0kRKT6PG+ofe8C
D5EckBVTyGhRpPLr8IOdqqPekAUqvfrzMTQdMQvKQQt+nscWwwMjMxcnYGJ6Tdkn
L5TiRDcX7D/5JEbQqA4I1jEM1OHMiNlpeeyVX0mGbB03kgvD4PfmJmlVEZSN0Psb
qigqgHzMOZj0xlR5n4WsLHi5pPt18dGEqU8hHKTYc5Xg2KBYD4livM5Kubn6TTBo
6DlV8uf3FzrygWaawgljPqkkqTqtBVVhWctVMmBhIs4SxADUbJXN/1l1aTkSojXn
sLlG2cxwJIW8I0jzkpb4T2Qs8sq6IFr9LWu0VFfJv/gNoM0IHNG/A35u74jXB8gf
DXA4Lpnyg4AmLiK3bKX2h18J3m76PXMdYo8M7z4KCT913H2LITO88X/D8aRm6owZ
qLEqaLXcwzQghnZ73L9qghctLseqqg/kdxaD4qaySXzkaiWxZ8qPP+dQwFsxSMDc
VrNb4kkV06tgoUOZZLA86r+uVtlCIp+CZd2aeG9X8cs3M76K7ZJC8e7JbN87q+TL
VDCn892uM0Xuc8dQlSCEBZFKwbiPa0edkibCMNb7Rd4HysPlb0WIOcb10pucsL+c
ZDiJvCVpyaMsfLvwTAhDFaS3f41TDS2DeoEqRTVDXDOPvwcKcf/wXeOHzD2P7Yk8
2bwpgsOSVVHJz4I4vPnV6w/08Sg5wUNdKVLD++R1J4kewutTW0JThuEkJu0k0rbv
SbnieGiJZevlfuFsJeUzrZT3vrXeCIpHklCwSH+PTKVG/kFf75rYw6aKJzE9aRFb
XEOd2K1GHPJZis1hMiQOtAT+qdZoGant21XE7HUL+vC7jt9rbJKrGtDJpKfE55ly
qIYBIveeSwmYl6j2OiaLPJq6rdFKrwMDC0wQ+1Jg1E0FvMWVDMCGramfVKuBsurW
KwnwqBFimKMdWdyNl0NGXxZHzQUxyxQIAMp+NBz1ZeVnY0LiB0VdGLNmmVmj+jQi
Qk12FQwIZoDgHUPI6+zEuKC+78018hJjIk1Yi+kC0TL6ZQhOb/X1wMeMgEJiqR4g
5hmS35l2KlY50kA3iZuQI5pLgFCsoyZtViZ6JvvqHw6EORk8nyn8OU/28o08THOg
q+PtYyTgZKMokNP2oLFmdG7N2GQ01mWHzUuvQzcyhFWdaFmqjMU9eVdtfUNgXS8X
hVgQMMsB3pQA82kSSd1rUHUZ92CrhxRMhdP202jZdaYgVGhqnaX3rEKHvDeqOuKB
ddxnrhZMekjAHeU5D0uUqXnAuH/FWzNtaQY1rH/EQ1kixOwb82FhPmea0ia/RmJo
Sr1S/OZic+Ad0+abH96r9c0lCxWug9zUPUaowqVudCHPL9mLp3tdwYmjpKMbWBXj
90oZH9+vCPqlLY9k7ySWP36xTiaGppGIv+X8O0/ObTyHB1c1xmoSiGSDc6L8eRGU
sQU+gDLn/T/jU6eSAsTsx50CD/Tf6sOy7lBjpk7+PTQiL8DTDdCgSRRFkMZXz96F
3CQeHPQsPdh9BK16/S9p2lIKNJqopx/n2TYd9sQT1CEfQybJKzFpQnq/uekr5piD
V1Ga6KxOLOef+ZSe8o438WUsSfNCOPhfwk3JuelLNnl0DTQEEvS+NwuEhsahgxQY
4fRqBLC3pSnuUtFHXWQEAa99VByFNd3ZzXusVR2xRLSHTbJZeH9VAvnCNy9HC2A3
HERN05r36MKnhD+eV+h5s+99+Iyl7ukXyzqAxARghN+NzPDWgQX8UPlMYDpm7j5J
ZzQ82C9eZhr2OuerA1HGYlZYIbcy2eZ4vFOzTbUVZsUCiQUUTkWIP4iOYazjwNHT
jarGjsDkk2imzUeNixfzILXxJtfslb/8/tYWNkF4t8VtpuyYlUt5/E0fISYZYTRn
Jc9sa3WdhXPDNd7zHO/HG34KtyvH871MoqIybJC0vj3PJFvvp3xJRa8F/xCjFwL8
PC+CMPMrjDroJW/dKZiasLXBT5988CMrTdK6EZ1Ik4vRNL6TMSdVz4SxOhXnEJ+6
WatQsJ1LhnCFabnwrP27zbj3TfhKCDNph7AfEYnYzgbW0fZsfIBMKPITXTTPl52/
pC+LiIqQWl52dU3tQaxVe+wS3hXB7MpC1jhn+vymlEV1fi89YwJMJGirK2Fyhsxq
yGSxw9i9w3eujHf36mPIrKitDojm0LBa3B5v4nfrTT1mCuGxQ09u3xIHP2cIDoUj
IjSGox24Zq5/MiCisRu+hmsBprFA3TzdfkJv2WoGKULkzvl3cCMktAL+011CdTgp
YvG+3NPTpxN1G55liMR8L9aeY9abD1ec+fzjUpyWh9xMVPWcSd/+bUMc3odngpJA
AbYhR2Xpft0Mz9PVHx5moyrEqP6DbddSlnY/zATsPlUHhhyEDBPpF5iEnYTIPmNO
DhZ+95U0j5T41NOISJWy2k8dtIvEuPTcC0rdkhK7z+pyUj1cLiLsh0BX75xdSA7I
ooJ5Oim363dmC6WnjX3cbL2ENpMrUXcVLiud3Bj299qiK3/SVi9cotD9+E0VYB6/
LCpjGmKFWLNSiqURS774CnkWOm63Sznb4smaEHJ1e/tUl3IsCAxwiOcUli+Srzj8
DTLBB49Ud8CSNq1+dzFt1K7iKtCN/A0M8d6wE5+vbaDLkmNaz0VE9NVKr2sww7LC
9hU6IIsVhU/axv/VfAqKlKMaA6qZvBIZUfNGK54FqkXt00wGB8/ULqgXP29JwAMZ
WPTV2sKptULByrhn0DlqlM3fMe06yOIi0GdLOFr5cBfZh7c7nP4s2Zn8iPfsEy3P
yOcr7kjGlqigI+l9EB1kCBYxQermBOYy5P+9WbN0+wmEOleZDP9byKe4jsfpDtbH
t8IfkCvleoGRLR+Qlc4qdX/NlZ+tf4MsE9Tyx722YhVqVcgURKX5rL++zNmMDGeq
lSWoeNEiz9GUMe8/W3AHC/LhvF6eLh1BW9IiYZIkxiU64iCuaxrSsIOtPMojQrzU
PpiV0dtgmkOvOBipG7qXFa6YnMMQF++BkGlotN0FeefbRZm4NVZiUcCeVJNH33TT
BsRiD9IMaYTgA/BEP9lHkQRVg3Mp+9n0I66mpaQWiK4trlqYAx/10+qC/HoKgGWz
ENove4Pq6HPhFAaQLfMVp0XK4imnfq+aXpP2Qemybv1aWIADmHcVkpQ0lQAeVfm4
ho7SnkBaSnnpbMQVPyCMsIT9k1uJQR4vevqcpe9CW6FoSqMN6L8H9wqm1NGD5ygB
LMmS2DMcyAb3PMigswAkT4LvgH/nSVBOQj1C1+BIin4i+O8itNvJ9eGZpT4E/4RQ
j6kI8n/eqqAy3W8q2h+JUUfBJbtBCibX7zfzfDYncpZs1/Jp/VR/eUijN8BNUD2a
QJqDtnYiMCXgTe0xqFeYsjnPewKUCEWC3u7Ic7srUlKrB91pH+NURSjb3c7fumDM
nV6MkSS6F421yw674o1MTQmvkYbClwc3zrXKDvCvup+Vc94PIe/RDU04IadQ8pBm
+MiynCM3bshRmxJIADAS5JDYAvQCu3+27ifURnXjKHHJlgPBLtgeqgOMRGawbMZq
HS3ZoYGHdwoqg1qcVRVH7TYTKC2nR3OCzlM70cCxM0ZZSxHxhGJvpsBaEUmWUKwL
FvujZGa4BzNJ0YBclfv4WSxk5WjeiavhvkYrkXx0qpjr+z3M9mnAciuilguwN+Xi
nQ58Bv/aWUtafE8+XAG35zljXlB2y5vO9pvvn/l3+odzdmtSR5FJ9ZHhs3f8ahz4
nfx4y76zgl5E87qtns9Gsz3l9f3xF/8S3KZESQl/w+ZBlKfKhAOICQ7uTOOIT9Lz
Hu7PfsvBUdseL6gCpgUXEgeIDAu3ndQKBhHyQhtMwkWY1SDKzmg72kVwvPMz+SNZ
g6dmn5x17a0mafvhFe48DdF4vAeqH9UrNyMRbjEG9Q7EohOGb78HFjKklfeBNbUC
O0vQn7bjKT0Bmfgqw7iLD5+dUjicAL7Hn9d5kdDcz695YY+OY8XftdjMbuGo6s6D
in7Jce/4NK6A24FseP37oA9YmTKoXltY4MujzisgGt0SvYGjGnah8qa/mNsV6e5E
YFt0lQQLIS/VujWi7h3fTROsfAiT38zGZrupes5ExK6P/Uet0p315xi2naVpP3G3
AhTGJjc/ulAx0DuroCJ0slap9Gdjt7mHGXcdUq3LRcj3nvv/0+Fpv+6TW6loYvyf
oLA76SkXXWfYGBk5wlYTyIDHz8XiIp8SAMdDI5BsHvaL1oMGXkeDy6RdPzGUE5Uw
f+kWZ29M34zshGMA3gUDeAhKEYOVGljE0I8f7u8ERwtNc4JzXdrpDvz5OlhrUp17
QhqEYcf9A9HRXRRqtzAARflIFaR96YS+Q0pLKPz7TB/mJ3R9wpRikNwXqLynJAJQ
e1rQRpZwdxFs4S5tVKhyqn/A3MkUEbO3r3evmhKO7a/Hpoavh0m7iOWvSprKtXE4
ME8828iPEK4A0F/RxJs2qJrEJv+8qHzU2hRSKTW+3iGR8+B3qfoc1mpBK7CuxzFc
s+YHeJMExRzFfxIyzlg8Z0yv3mZPdA+6nvdpXKYzdENGdjS2mv3shWDFlo+I10E7
T9UNvwYn/l0WKsM82x3VMtB5YCXrGKEwd8tVpk7eBlm54ngdH667KMz5tn2IoqpR
WvHoS0Se/U4fkIngkCxwp1RyBSSZAlSRbVyaaxwaeOebRFw9aGH/im560v7MlSzN
HMg/63bA5OH7P0bjrbGDPi1l4aFg6N7dU6s8s7DVWbEmwCzARokoB8+Wd3d5zakP
LVZJsfQ1NeKEv5kEIEO0JUQTetLNeYjNRni/YJiO5YHHZ9VuHpnDWUHeUnzbkXQg
qYzVKiS0Opvqmq5vfma4rm8ZOIO1GMBQJgm5n290j20e++WYnlQGSCiuccxd2eez
+Rq+vYMXQV4f9k71qtQNodd46YUeII6SO/s8DLyv1TipJLRE+lSAi9a85YRGkhtk
FONmeD6M82Kq60lRnBXlYN/tOxutnNqnJRJbv8h5NjYPEH3G8vD6VSbfYLzs4J7n
W31/eZEPOAMNify+Pcqa1YsOBx8Joxkky13EVJFyDojuiFgPYaNK5/94HyvBesDo
S/UFzjTiv6sR/rE1sGRZ99bmJd/rYJRWPR931KdbrDsMax11FjV/K0oEwqqC1ABx
JV50Luc7yH+nw8ugso3g7uSWJU8WmCoecOWIFMinYF7zNtfFx+z+FGSsUViEPYFn
VG2vnXaNubeXL431CeCRQR3GzrF5lglVqDpYXF2cZfsiMdUx9H3uCvHkLZxntPmZ
6U3dNXl1HU52nXQZjOh9A3pDMgQmgfyUEUngUKIteBNbEpCqXfRLlbqmkKilOc7n
KQwEkMr2by411JcDblxhklo8q2JAObKcsFHtdqNWIAwETAj0i8vpWoLkXl429PeX
y7Fmoz0rjoVWfv5NLuiWm1GlZsnzWQmeyzbQBTpRqffTr+zEE+dRRVW/lKWPeH8r
1QNQ27yYa4HgChkwt0z1aNuYbMJlwtSA7LgmPyIqiwj4vd87sGxFTD1fbpmxCyQX
bZ6/Y3x1qglf7BZdAvs5yt2WSEIVNN+oqztwBfm2PRnOQv7TlObOBXUNHMuxvWLw
CXgCdYK3u0nfoAKEUtjnCJ31l78DB63qJxfv5KPcEk6rrpsimyK/WVM8fq1NBYzT
WXc3QpGCn7iMZ6xynvCbVTvXU1T3j5Q+uHRL9PcCuX1DMutknx5tVwmErxkUg5Ka
oUCeNSTh/MhQyV4OdBRJBvY+c+e7ipNzlx/qZLvHX+v1Ng5PGCInne+skqxkBfSq
lv/MpuV6Y7vt1Ia9l7P/CK4CmEyHHAL4706Imlu02Au82OhZo0VDTL3TztM8APds
6zz8eOeWIB89/tkQi3nRWRc7MPT78DmemU0kQlJkONJzs8GVBN+YjPUC92Hf5CJH
cGvXUEakrOkhdS2kuOciI/X5Z+SS3KKrA77aFcI5/c2xdUPx9/7/v1iAvyjeaKMY
G9FaZu3RFommW0+kBSRxWWaHc5ZVjYbGmrLIoRG1SI/9EohX9kh5mD+GSN9Hkne/
AQbXZ2nzFACaONDK4OYX6lHfS5bNUjvuBpGHYO6CFGQknWQke4Ay8Gb4dRLKwgit
9LsCaXqvhW0fhM2jJ1nGriHzwH54kUvN3sWL5/lds1A8QRyNqundFfIYkaY7swZI
qSCb3A33DinkWZOjbbpqwvGEt9xMJtp3BTg1f2LSuwIxDFss4dhczf4eAwlrE6gA
AVbYm7UkBUhdaL6WQ4W4OHdEYEM7qFloANC+lKI486Mom0vqcxNcq/vJYIyhznnd
3MKmp0fTv6pu0gWOy+O+naq8KePI20do5A7R/lPYHdSWAIFjRGMrRkcYIm6a+Czk
x1MHipdOaLFh+ZPbM6Op2qopN3YeWBxEL3BiSNhedanuM0QzC9G1RqSyXFM0veJv
YZFU9cv0IwNEiBlj7xu9Y2cUad++PWlGzfnC4AmWuNmr6f0Q4xodVij0AZC0t39h
d9HMCWWRb2JEhvBc9hz+YUquS999iBK+sBIlavE7888GIxLhIRGcjSoG9gmIhj49
fXVyMjwbGiyBd4ig5ZCG5Cs03wAAXy22J7rH2WE5s2Fax0t7ZFCLhZlftYKfXdl0
ZFwUg8Pi5wPC/XBuM3Qumv+f6PTXLIxSokGjpkD9VxyAACkPHqRvYOMyRCpavxcb
6snsO1ADJ+dID7Siy68uYuNkhg13GCDaMbtW2PizHjYN+Cz9PNrgiQafN8qVYAIk
7UPBsdkfIcP0o+PY6ePE2uSwFkcRD2Ow6zOmqAQogtCijqhH6B7vipzEKco6rugY
e/xrF7uiLb/TbWIJ8QgNHV63A/FwE2hJVn8kE9oFZcxanCkKLmsqAppqzpgyoxFN
LXor5BUHw0h7BmGyLyIKGyD6QvENGih6q2fJ8wpyEe+a+HvxhyN2Mus+2eLRDr1r
2SGRwiNanEP+TLfD9Z5wq4n9fpzTiA/TC9jJSWgnmkPBXHVoXXxqfiftzKJZ8cjp
qp9HfKOmoMEolku3b8D2hVGmZcOFUFmIZVPAqbdBy4MHDlGCv3BOi4KMJTXhqlTl
A+1L5CHp4T8ogtvqs76JqivgjAlCsFqJXgzveaJ8xR4oj4YOEJwHLyKpWgZbNbtm
7MC5QjOqYrWrQZ8/QW+iu5mY2XXH5U6KhayhvQaN76sSVq6DcuBV6ZKkSYOOe6zz
UJrZKfCwiKZSKVHQiV4TYP34i6gvlJ7y0aid0wSdEzJIZwITUrlcO24UGFfc93Wb
WNlOI1gG4DuWy/ZImjV7QmYdQPTYri95ySH9txnKHGIjlwS3QEp3Os2c9nIAFzP9
VL7Wmo86HrLXaf8uaYg/VocweNhytMFh0dHdFub/3emBHFRdHmBNxX9lAHsYt6Ig
CHNwdEO94BKn+mJFwrXrV9GRrF3wcTNCw+PofWSIbBwLeRIuWJQYoPMo9rISPXJ8
a49Exb+IspXypashRY0NZWQwLe2ChR2UOZp9IJUpzcN/OLrM4dY5ui1250H4uaN5
RaKAVjlD+0t1Brb50OiO+iNgXrSizdh1y87VuGXkN+BJjsekUpA4N3ty4v6YvcSZ
cyXW5ampeDxD0hqNs0GMoLFbOqHVEDayrgzl8TAz+EhF58ndWKJnwPMY9DbvNLcs
Dyyp/jOvEgdcvjLR6iK3lrhfp5FyfVt2kQK2iK5sjtjwELoYMdWRT+SkI7PmT4Jz
N3NOpQD7/UkUYz9Dl7zqDCsrkklt0uwjJmNKGXNCpZeLFNVwgXQdwcEzw/AGRLFY
WHFRMr+YB5FXxnKSYf2hF4HtmQcqtQgiwv3Ew+2bSf2ItA4N3tXsM8wByYWsj5ht
oJBFPY87QktFqeX+24jTc4UeKydD9QV1dnW/bwWHkjnUU12vkaUsfLpaJhHOTtYh
xSEUVk1ct/IdgSRiaUX9mxvUq6vSmjAllZgG3dtZNFskhZDoO8y0t3XRkMKXSM3r
e1JDrs3WyCymntqyIDjwORkVEuJuApIKbYt4LzJGV2YFnISCLvaok25cQM6oM7Md
C0mhMZY5TXK+erDiQUZgX7ZUTsYKY+qwhHJaUCJycKRtMglW2dy3mE5TYgDr/xdd
9C73CwBy1WYxDJJrqoQxyfq5zlp28SDrBnHj/g38QDfW282yaSCiIAa7ZbGGWoTz
lO6X8l3ixG/UXIPaM6kEZlXQqgmvPBQ8N5dSAOCClKbmTr0Ny+4wuw+OWL2jrjkk
ldBzW0O5SGHaiBEhLY5kgdK0bXK3mzVovwxDmcORMuw/D540GDpCSxETnPHOTelX
uGx+Kx1Wa5yDkn8F3cwdbAZ+ddiJbXwsXlqEnON6VpLZzMxpz0x5NOlL9RMpoK2s
2/UtnIMl9Ex8ImLDU33xSxxuznOrzRsHGst5Yzkw3DTsP/95ax06EcNmq7HS1bu5
BOQ1LK7zlh2yTfzeVTAimqA4DFcuj7uTw0wtuibZfiwUdqL/aNyfnPaHDab/Ckho
SjgBeEYOA1ZW+bdNW5R+UiaFGzo9Y4eYE3HDTDKEUgXtKAX457eA9d7DnJfLDG5Q
WXlIk1Vpl9qigNdtKuVJHc3u6qwRCJCor6AACrj5HT0DSr7zcEIswW7d659V094b
VMdDU05ivt+QXg0Owg91aLhxPZ3f2VdLiTcum2vypOeItYZz0CMbkm5t4LevWgcF
E6MgqLdsr2XHW1/Uo28wHyaa2jmPLB5dwhMblyoITZgOtvS6ZwqxMlFSrbv1OD9P
bfEBHHURzgYPKuZVt96bo1OukW+4wlsqmWpvR/xjTS/jr1EHGc7jbtnHxXe0N6qX
o7/Z5NW5R7ejEH6lEbT46LaD2AxGUWVdKIxHy7D9wSdU8Gw90ECm8er9I/Hjgpxv
t1BKDfu3IkH9JyhJBhz+FO/MZYAuMDO+c+zisM41Yiu1fnXr61gm1XMSwEM/Vfnn
zfz0xAYMgPOVdR8bEokjIdZ8eL4krBJ4fKgVEaAyuKaye8eoRBF8Q70hUETs9NQn
NYgC6nkGl0lAZfDzhWEcbpM8ab5c+el5JFN5rpAfyCHLvKqbABgy6XC/nfja6s1d
8uIS5CFwqUg0gihwMpQ3T96YGpkM+Ivo3ews+03kjzmWcbbsv+GDdHtX3AVu3aVj
YSUeKZ9rJP2pwku+DMZbngw3lBPO9lCMrPBGvvPlC30V48v2TsTtucKU5H6LU0tD
EEHFU00jZE860WsOO/Sbmd4mJTkZ2UvZRgV5KQGzlmyxM7X5TKv++9d39S4UJAX1
/0WX5LccSL0fjiSs5r5wGH5xXHrOEnPlJ8wM45NQT3ajfurjWWYbKnOS0pfKVax0
b6qBeB5nJIwcWpepXV2x45Pkh9hCnj8vlhcG06h7VUT5mO6d1sKV+jAN/wWhA9By
4W2fKE+4sHLq0/bzqY+JMH/46/dXKeCi1HzvlfnDXz7aHjrmBgmzdldU71yDVkGP
hmn+PkAZdVwShO4b2DRrMfzMkXYqDA/9Vq5fx79vmP5Bx+KfZF1KGGqBvLAeOsNl
TCqUDoCP1+AJEYynYC5B/xyqHDqibrXsmRzceqOiTT/rTUf3hCXadQrMjnlqJKIM
BJ8KhceRMdO5Zi6onHBv2cMgh1HQugrM6/onQV5Sz9zYsl6XE5sMq/J6IyglwAKw
Rqnz5HXLbt8N8RqetrTiNNHFYdRBIP61GJAK4C5J5hwxP/v1NOxpWavbTvKo/R2E
iBsBins27SdQafH0h4eFMwnSBq/sZ+Vd3SRYLok2rUl9p5P9LFedvEP+KpRk6g0O
/hi7lvhY2K8ZKrr/eM+ZyGnJgKeeRWDIirxNUehFZOSXsncUagpKWUXP3+mnaqcG
W5wCoGJn0B1rQhD7Qu4PM4Q7J6GrwiZcC+cEvqt+bg982s+oyWO2E3dj9zN4CBZh
/V8dbIQ9JZC0XJuHv5rMsRjkup90phkCF0OB/qwJ5a7gRTGBDbpyn9IfdiOHlVXw
RUVdedE9JkuDzlIKXFGm7cBVoQFMMS2jI+JVP4VFvOAzqXZzb9nt1vNu5yDMLHBM
Fi4zCTj9XTvdMRMranyBphKqlDfrKTd++42M+FsT4OHzqiv5PrbV+E0PyrbBbkZA
z3/B/c1DfDEJt3bDUaxF51xy0O4StsXqBMiw9yl9lxnIPccsOKEmuxBJa1j5A+i9
Qi7/snrVA4DF7VLAdPoJR5fc+QYhPuolP3IooGEYhANKbHOSxs9NdkuQtcWHjv/G
WspROyW0B5iw+RAGuPnvt4oAOfuESh/kZaBTEkn9VBuTCFmmyHX3MeLXXHhdhmO8
12I86xn+WcprkCmjYW7CC/AfL3JqFCt7qdTCbjLd+6zoyqavc8tlkyxYCUfjs07h
XdJRSOOuHghhi9X/HGQ5ibLY60bq6b9eBC4Et6dZPx04TwyL/L+Z4633BSMjAGgz
fIKYkT6DBoR7StXNyM6cN/W4lFXs9YsRlDRw/ScaL8WQgjZl40k2Hktf3JJtT40X
hYp7qh8vyi/x0hZZATi8zEodJVm8t35UkDDTkFm9kOT3KN5Ba68x8XpC2t/uwKHC
LPQFARO8EkKk0uqhnpPCXEHJD7Yt6bwkiSL/y6uUUEUoeItnS/89EiXb5fhBvdWk
IyM4UgD5trk3Q16HAADbHOkSDjVH0caBRaPfKT0IV0n+K2QbrjNPT09UUD9shS9Z
b502BRVj/St609wwWcM88Q4CGvJuu/ww8r7DZrq/lWupgpYLiip+KraLib56w941
RePQzhhaolliY6v4MX8Cqf/tJjXJZxSEnxlXbjOJutIoOxAh6fXsaSIKb6DN9e5b
XHOQFb/pBxdX53pU07iYQq2TQlc+aJNh/oQcbnUFWlQu2+UK61iktk1NhNH0/D7H
+zAeTGRuXJ7VR1NChpN2EZYS5bHQBpqHQR7N7IbSXIOAkUOjxSPymWfarkBoLU0H
uJqXNXxSBLJYMiB3AHf5AM781aXk5JRInimTHN++Nw/LlMNQWPcQ32LMjGNTQA/Z
DfbFUFZSQyYu2MutscfNch1KPe3YG0TN6Y58jgAZf9YeWVHJ7gepsSYjFXWgn0ds
h9oBPwzcIFlg6cO2VTRICbien5yFjC1KRbNrS3lq5F6Qw1nqJ3ImPz2d4hOtaYwt
pjxfXfeaN8N4Kcnuy3aF1QVKUKDRtnZAbTb6AGxUKewpZrnMlJqopE8koKzRy/q9
clQYUlakmtjo1ilNR/ZYtDkRqcbAz+l4Vopy/8CYPViQvmXfQdAU43qyd/Zs37+d
degSQVS/8lghd2dfj8fU+3DO0XMrgYNaAvS21+j2zriJ7uQa/5Frtgfp4QafhG5e
LBf39DzRS2VRyAVSaKukz9uXbfeBSQgioo/AUINPpRjMy1QjuxyIq/7Z729ZQhHS
YwGLR1LPHyY7tKVIcRx701hwoQu/JCZbGmRLP0xw7MEB9It2S8tU9jjN9udzYaKK
4YUm54kaIlv2gNMGI7ELXdRI5gwjqeXziEitPjcpPEb9d6a3d+OE4lwNbFVxZvFO
ho9T9XokGRyBrHnaLPW7sMXkJw0kq2UKJ/2FY17ocoOVdKRmEmTCVTI77zZCDGum
CYCJREoReulP1BxR4G+hSGzEqii73xQrFSRd3Gfz9DD9SQiUDL1c3TRXQ4aJSgUL
xDlBwTm0E1/iLznsb05nTesWH3m8LGn7K14P9DImgjRCM0DDR4oJa1FLQq9FeYl/
PxBFJCzRb85838QBrpQM+q1B+Gc31Yioi09JxAnmEei7C6dsJ6SQayVGvR1uDete
TB1E8h4fgZm9SUTGP7SU6xqHO/cD4JkRJvIU8Dcdxm7RQzIhZnxhrq3nUX1HSDNo
/ovADy4SJY/MRSsvwU16sN4Fhcb6NOy0JwwUZEA5lewqwdVk9NvT1CgP3sF7A2L3
LXkcJYwWBKoRvh2Fx2ab1VAkoShA3TzrZzvIjTKY1rMB0e7ttqGeYcTMMvoNXbCC
Xrn6vsz2wARoxqS8NLhJ96BiXAADmsQA/4nPfmsakkyfoQauOv4IRPxq4pNTM1yP
OvRmfze8iLlm7MKYwOLJkm1AZwgdapE1vc7nJ/+92cSfOwLOCaAud1NMKgADWNEC
5Nba+Dq9xRsebdTakC7lh3JO65rWlubwaUM5XwHu3hoJ4NLbhSqOSYPKqDQ7+Qxk
C3RkawK8RerwW+0m369nX3hz0dk49mPs07oyae3o0PcEw7dowCP9MtQGoOjTcuL5
ZjJEI1P4VERrG6Wre+t41hx6JD+2lXZ1cvVaFbSpAuUiiAtguRRHzZ0GuoU9xVhm
PJ5m6IUrxQfA+giTf6bVDJuWYZSO61F0vzPtCQoEjkpUUgBvM4KEpv6t2tBbRLrC
aZm0rdB+hO00AcFVg5/BvFBtG+wPTVzA6ch9M02eQnbXDQg/zSyM8NfZh+hYcntT
MCc0upcNreLddS9dQDEvKBQrhVTKGqUVEiwWSZcbR7fpErQqSqiNRMEiMQKxKNbv
YZqeUUIsaTPPIcn7OUKlrKfV2Y18UsfCNIPcQr0d2Zuz8leGTKBgmTOS+3mAoxHV
c8HJgUEV81m+xDAhDLaQ3jlWLJ/vLD5kXQHDoKHFmotDrgR1qPa9ysxi17stPHlx
+KKv2/djnekxmsHAwODJ1SNHLaMgyDa+gDDTPK6qJ43e9rdHPl8ygOy7C0ayI4rk
NY90ox0DL7fAEdiaRmoxytVvlbYTT2ki6PN9FKQ5qg2tbJwlbdyUhrJU1dqdWAgR
ir6tpZ2sf8j4EK4gEmykxZ6I1XGIvQzmH64lymL+Sazr8C0435Ka99HC90ecqgK7
tj8VbBzMN/2g7M2VntLr/yfQ0++dAcLj4dWN+mChKK6ZBV6bhJj0KPKP+YsdQs3J
8+21pTliSXZwqmRUU+5DR1RmfAhbHy82EOvVL2kY9U3Z+jINmRDe6qcP9Et5iKAE
tgtlinceFOR0TrrbzWjUrQgH4jMvamX8CUjbdPLOFZ03FtwUrNXIyI5bTSOi7Eny
XNdLbFlqnpUJ65lvcSpFpauAwpCK7/irkk3FWHIrpJrd56pj4GwwW8pkxiD2t66z
+LByRiNQ0vxuk4PQDBmfF8/21RcpomokwM1RPxPM9spuyq2CVcn4S3qD6+32TkOA
9MiW5kCM2MMr8NdDhaxKTdaagP9H4X9dZ7PuvgCG/FwyyKbzTroUDHZA5nvs8tHX
59KI6dorFMq5QEv85iQS3bk6n+3B3YL+RzVECBloQONelnhdIY2FC1hQI1rMnfIu
h+bKykr+NSWXgyGbBi+o3ZL6xIQeM/tJCa7/0+cqJxXYZ3hFooxyg8J1yLPSkQsl
gbsdQ1RyuFMHCVURSQ4GnJsBoDsdQ/oSYeIyrTnzI+z8TIqNZCw5WrvppmSRSqUi
rBZ2xf0PD6UnIlSkkToVYV84R9ofwTnIA5TTkAgZ3NDv8CL3DiMqH+qacmGydtNc
KTvNbYl3E3O+sZ9qK68fwc4QgFqlE6Hsw9oux142qKWLYYeAgkPQcof20+joNlcn
lZRJsZeh8en7I2TyRE8tz4lNb0DoOmNNwwSrVCsy9Mq8a9mDGmLX5kr8srvmS6AV
f5hqg7A1+REzal45i16ijSw5pX4CU0ieE/RxvwkdTUN30lDqMu1DcnT+k8EGS7gt
q1ef2FaQmpsnyJoXa8cezrYfPTUf6//+vTcKL4CBHxQwtDNekNksA0H77V7qrjXu
hytGpS7ZGiQPfeIUg4gyt9+7EuODjCPaBts5Lb12r19AmVGchS2d4dzfTMB6nP0Y
B61Z6Z0d+F2AYT0Zf81SzFRy5yw/7q3jRx0RcIXMVGfl3t6KZJE6sAcTx40HSOZ7
QLYhNMfxZfqfWhRsReoaVrQk0fSWtMWkkYCF31FoEoEfLVEW+/1nzL9q8QQOqDPt
rlbcx8i7eg512JfHijmtCaiFwtXxkkekzvFtvW7kFQ6s2uPVSPM+KcQWPF4iD/dT
Jnrkbxc3BeJrtnjOv6Y3cFyByApdiwbD7BX2SDTXJzaOg5P8mdvVn+b8NovDNfvA
T8Fp+LcT+McLfLYgz+Elew9SZHK9t9j2RVwSdRU0Npj3QCmSie+R53SyE3xTbHWT
gLZLEbTZb3RMiJDTfcUUxh8tzrqe28Zpuv54RJc/4gBlxnIPsUFW4MNOeNrI+d2K
oBM1hgxFkVogYUkxl63j7x4KCHzRBNCoZZQ8Ir9lRZ3yf0BmgjUerW2mN+7s+vCd
HNiXiUabnXupRTWztONEY/ig55pSwZja9OvDks33fiaV6rIzXvelJdIQfCTb0aAx
C1c4wCDJ75cNPMhrvVPzxqUQWhjUW69fVQx30gVF9rnFspEGmEMLbRVvQwS5IQNs
jtYzIp9ZTdyT2BoX8HColUmTMPgwluZfxq2YMufXo69FcUmaSUUSdT9/qBfLLqF0
gY1j75ljLrtr6wtpyQ4RZb3VilEu1T5pQNkX47F6UjVyUXiaSrYIVAgYI1h9L1vm
ELG/hjdzQLY9LbO/by2EzVaZV2m0PivdBYVtiIuCvAZOBJhVQZjc2+dU3xuV6F1T
CYfXJtHiC5VrPV5sJ07whSdsxipf3LVKI9+Arg4RQ0dr3OjHI+bYNZK6JlFGYs5r
t8g1qrZBpXMmw7BLRx+Zoqb7NZ+sHLp7lpUMWjqpUTJQBdv6FdW35P2VaQnL5VUL
CcUZMEhM5db9Te85O4OzabHu/QF7BeEyKkxqU8l6D7zGATUdQWAuQTr7FEToPJlb
+FnmrMmhmuddbWt6For8eEI5+uNX5dJRFw/YX2FUMegj5HZlZb+Cbp8m4ir4ahvG
3cfQ50eVUrRMY+w+hy3mqxeayEzp1QYOpXUDNkZKhxv93JRpfEnSjlphX+x92oRR
CHzulyaIeOGa2llps2ZYNDVpOGn4M7JB6dpZTJMpg7kxZytM4DAKMwR0RFW+opP7
OXjJS7nOdRCV8yRTliM4puWOL+c7N7Jf/uIaIHfrTDfvdSuJq80l3cBXrXzPpDrn
vQfMttNE3o1pj/I2O1jsdY++MlScKaPlXmY7uPYAjGlyNjpOo8ioS84ihJZ+QRuO
xDEcLk4mInsf4Ko+2h4KeKbsh3aGyNToEwq8uVOO1jDi3rP02vjJMLEnHsH8RLWe
+BavD7kAP8hPZy6G9adfq4pmKO5zBdv1khFrzOWFU5dyEb9+sMvR2oq3ysU7l2z/
61g/pur7/cS3JlVxMHB3kUum85YaFGox//EPBOOY5Q9ytBRxQFf6xNncQ7WTdpp8
D+4igRPH7BtCIhMsK9uSKj+FnG04WV3UkTFElByVHGx8+w5Mv6YFlqDgo8FSFWkC
OUeki+5DwFVZ2h80YLwLaGu73+Os7li6OtnKqm7L1DVrdSayDpXsPKhrxfjRPZoU
9CZ2oB7Nhn8jjZ6f/9hHfqMA2k9osr6g/Sisep37fJ9NZIfiEMHvYaRLs93DB+8W
6JbaVXuozAgWdpSx5o6I019bjnAlNd+xBO17Ie0gPC5PpsikW7EpaZsMwRjxM9or
Tu7l8TFcPXY21yR8dS7aZjlFTSGbXsxPm/qnYVVbNVGGpj8P7tpg5mR3W23PgetV
BCwqNfnBPRJmpmr5ypjyj3TgcuQ1hcHM2HdaAcusNgMZAvcy47J1Fqjqg2OkBX2Z
FzqxyvZ8grGrF8Dss4hNsMPmpU7Iki+KmmhiYfrNoui1zIBNcsyuIRcFuPE1Tjuq
/ORXM4JcWc1piCMUuqaaclmhxdPmElgGglMu1VZcQ7U+UWbMm5JvqActPqGCD0yb
Mbr1+QY1+Jw0ptWPeE7Ct+2gYAfEypyYp6fDPvn0PrMavNmRBlUUfEN7KO3STkbZ
lWsZ+4YugcOGBCvw6dmbSMD4qhKojuaMvec1HjStR62Id3iOM6e1ludWnnZ8wz0D
eKiR91KjG1ls82WGIGQxkIC/7ElqUjXfhocUpDnZ4z84IZKTqc5d6Xjm/1a/wxqR
HRVEomiuZkAIkuLN3I4jS+NvbxVV3paU3h9q7pFNsgoKvAhy0qhMbbDp0NKYESZ9
EHS1Om8xep6ZjC27OautL/L7VhquBOoy6Pelg+AoyUieqvO4ueqTau567deXsllj
T8eUv5Sva15SMa95+vskuP86afHyb02D9yD9phEKov0GCsedDpYe+GvVKW5lLCUW
gvbw/qD/oI9/hqNqhy9q6W7wLFXkAAcv8ysAGuC7PdvuLqsIAD06pdemN6lLrnD/
uFx9KAUmAMXMFWGuEK5r1DR0sKOcL8V3wo8Cs8EgNwX10r20/2g7pbLq06VxeBiD
cuC/PIPC72FLA+JaIrFH9lBIvI1o3g2J36PYRbkZo6hJdanyUKTEWpDOSIiOKr3L
LH0kwQccbEY1ETFKk4HT8QCnjeI1jusLpaId0N+Tc2rgZ9UueSuKuVF7t6K91/sm
1lWHxQk6r4cvmNag2HtaQfNihiy8lxStwDnIVLodFSCmEFlAKijqDFSXl0nHIrRp
yqYrHEj5psisBXHt2eniXKuBq2CeNo7cggtQGSvuGyb4gvzmuiWPclKITAJErhsR
YlMQ4RFbOsOIjQ8v/tRvy00dHyQzHQF8yQAA1P4i7/N+toAQBhB1Rqu6hDJi/bX9
FgtuWQkQEIOV9BaVO2rOBs1mFvgnIeTL6J45Tss7tZNPjo5doiypw9IKy7beYGic
tC+vSn06OSNZ8j7/krkpTM6jkdsQwRh4GnxhM6vwZcn8oCKwr4G26KFb6b4lD4dN
cj4XEnok7aGarsqioS8Cr9omLhxt6jgUOSQWX83ZeDH3e91e+6byOEcVc3VzTGwX
doE1p/ruSStfUN48z0Cmof9LKZHRZMmp/mDcZhfKJ34Xw1nrriyI5JDnLg/9vTT/
DVSXh0BAUm4q4GgmTo5VjpGwDlmkexh8xz1pwryu2RH3EapFegDKdRIzNzwsV794
owpWldckSZ5hFJL7Zwo2TmRczryD+nqkxcvOCheI1iSHP0LPXdaB4vPWFXd/stl9
wYze684TyR5F7nOpR1FcTx/q3efIcvCkX6kgswdexl/++WxGt4gtJoJJNGpCOCH9
Rn529BnOpSH0Mgp/LeS1KZFRUWri1/fPP5kJgUSaWSPXQvAZOdFyQCvK+Nxfv9BD
jL3/DZ1lv37C3ruPwA0OKmsRydauBfNjzFcKufacwmAvRsxnC1IAXc4ZTS43byFf
xfROqActHG8yG3yhiuS9HFNcfWBrA63fcORmWmOQHIVsOpvkOHR8/rppSXPz6oVS
oowsmCOca1u1kDdJD7ZjEWE9KySi3qApGB/qe4HBwXl5nYaUIwZXWoKwsm2YF3LV
aAh2WPfnxCBv3umcQZioPSsDLZNaNW62CCGxtYtDP8H0tZXqoAmLmP1Zo3TFBN/k
48Kj+zHMCFICPnpHmGdxE1TMnkkjhR+Qm9qXljfGL4mdaSvv0oJG9gSbLdSzlE6h
wfR40eV7+Va2I1taI1yEAXCNL++N+jN0svQ7V+JswsQ5a2aQQ499Mz8frB5A+Y+p
LVuwcCn0ZRCacfwFfvbaOTlSCN1O7bhIX+GJ2TOgBxzbM9MlWhRqSoOxJBfvqFPa
ABD86jy46LcoiuQ0UTPMrEbrXUMPLXKkaju97UnMZFwiglNI/wU8kCQVUkmoEoC/
JW9WnKF3CMG8J3eYd/esO4L3K1JaFgvTOgp3gQliucfJV2njWygeYAFgIcIEI4Zh
EX154a6wduv/DqvzmDQsccy1BieLTHpDM69cGU/lrdNDhKzJenpNwD74BuKzH6E4
D6B6SMHvRrYhyOWRpVjLNEgXQO2eKlBCsSB/6qQhx85UBx0mTcrIwRVr1CzvUmc6
lI/UjWVkKMqSwBIQmX7/bmmDlbZEAeOEARWFgctcxHOdPqLwAWaZ2F34XBXnkljb
0bPf7WfMuLvv8O6GvNRrjHNBPLPcQcQkpMbGhf1C1VbxURU1y9ycCeg2Au7ua9qq
WbfRH7SHllbgjKcDldu95Xumkm5oGBBq5gX+sIO+twtBL4Pf6FGH5vzOBoPUuUaC
X3QX1MikIGZFCRoJcs2STavUBX7yikAvpKoySJj/P1KTxOf+fgvfu5Bek3EM/iZb
GYuOW9HwJl4QcC3jjqOMnEkR/+4JGvS9paIlBPpXbxZ0+gtnLFzZJEmLBpFh2y/f
7GU4eVGMsC8Z9HWLsTiTGU/shTyFo7AI5ZMPQ96JToEqu9fwSPgK3XtAzFf+K1mb
ISH7OS7sWc8caDG69qMCPINTJuLnIwXVFsNDYEf2gHhbOCRO7f7a6cWbNacHZx5D
vvxEcNTWyCZbY3s0z787wMa7nonmKtLBJ44vKtPiGvdXK5eYQCTzXsmCSRWdkhLS
XYYeHeMnjNXUluQSlv8ghD3JwaU+JbgrYcXrHixFPdBQA5Pb0MYJcksoG5XadOBb
tq1fTvtbHXivIT9Z8304qUKKyARbskyCT4EA6InRcHIJeVil8xpugM8mr+Jnnw/h
6v5CiWbc9ZDiHwzz9/VRsjIE+P/rMUcr/i8nL1vEiQGjV3RApL+E2eyLa875mrFj
1NgrMVU8KnnsjONNXLHc6gHrjmG7FYLqm0py80HkNo8vZpNLtWm7hHSf4bUfJ6Qg
hJOaZ+91BwX1P0mH75KGLiuM9yg9S3HfdEdgGpAGH/fmCAkH6jKUD8ZGLzzuqtsL
+8lVIdbQcAz2Fyfr+62B0R/TX/yWzGqfUGtZ4wLLMWizRc8+wGsKPUFBmN5+E5RF
IL0+/wv+aA/jPntBNbsLEB0Omh+ppewvcOo8otpLXheGWfODqeEZdSqbGy6T1PI0
bcJNcWG6RIYJtqP26BIxx/izkZjWrKzZuLpRu+KlsPDtwkzlUHUtF5Rp67eTH0LG
7W5YZhEfXjoC+wqpe2lbo75YRJfV95Sg+OaKtceTixgzes2Poq3PU65Bphgu7Thu
ImvNVNRUcnxI2sB/LNQqPbjEyUy3dz5EXi2wgkedtpBsgwGDTzS7FM4TekMOyUNQ
941oSqqpVWG2Ws+YgmUMiLdYETa71b1QuzySddPD2qARljTR/C6IbONwizxzPLhq
E7qSUdb3gJdV1yC7bytJSnNGCVkmTiQ/yy/B/vifNmGm+0b4dJRHqFM4TVDzi1rB
3nu88GY74JJ1ibAvbJLQzZ9keuGHuTLsoh+dE5EwHfYvq48OZklpLWoAzBuVqvbX
ZWIPM69LkHx5ekzRafX5eJIjfqYmGlQApaxAHCYdj9RsfQHHg6wZE/7tMuGRk1Lt
JHvdxj8wvZTzktttcGqUIY5W7NIvnY/suZZLl2t8ZL28S1pomvFCmark2/h9dq9d
YTIREoeE1qjsQom9XAIDDGsvLq9SrgojaxiOikFfY56VTgjlsUzFkG54NEPtp85F
gPlhClmyRdKdLSR0l0vfF3h52CtW45L7whxCgmfN2Khv5VdaS9NyQmbAJe6KFLF5
2dOMaH7nm1XZKatr0nnuxmS6GytlVOBiTdQyjyFy3j+gB+WYq7YTYhDHW3CHzPJi
cLRAv9i8f07z7aglyDUs/HyeqXnIeHbh/qgENv+mPHZDu3NyLL3Dtyj0fWMu3kM1
TnMHCj5TmbEYMYbCFOZpBAb70frovHc9C5APbXQR6mVjG0ExpXSCb1i8NZjzYROi
vxmKY6qSv/wUd1NbYmQZuWQc5M46Wcpyb46g0J96nPXeA29aq1OzO4ETxCCIXAsS
MFj89QvVMGojSWQGrZl6D+oEtkvP5Qb6epzv/h8JN1b2Q3miJsznA7Cdb4r0EZIW
VYI7CqpmBY3FkogbV3CIHF4wLfGVk8Q5UOmEdU/qDNKhB9aGP4xCKTtZzAJtc15b
g1+SBkeSdVr0iybNluN+rJNxNl9CBEg8irA+eCr6vJaURw5t5fd3TjQUc/AREX09
kq4VhLGTF4+DHH6sumHRZfysXuA8jIpeJYTT4JAdjs/uLzarZwwgjn5yljAUg02C
MAZVcAARilvHK1hBcFklUt/CydBSh8mlTkAHGaFukzeNap2h7o0hNdDFGHNvgszL
A4OhWL2Lb11RLcPYBXMWtHdzhYxzxlAnjLTTapmM/Dckn/2W/gzddwCecf+4cr/b
yTpVb99ca8pV8FtwL3UdJmqb8JH64tgB1Q3+qJ6IriDdZFaLeZeuywPwxWyj+jLI
bKTXrDScWamVOy4uyAftxHDHaBFhB/v3m7HxpxK1Z6FfXphHldHLlCsDU3gUue+S
q+BKG7ENcXz/CMkENYIZbvX7bQWSfg44oo+8QD2yDFX8VxpHLmkUvGD0uDv29EoF
L/bee5nATUisV80cwnn6BIIsGTur5mVMIrLiOWNJJ0KbhyuZHaOXYt3u2v/1nX3o
qCM1i7AWhQ0Eogc7TCKfEMcKgQVetnhdB2KYGaF2FAyNnS/XaK2w7oVhgvIxSutg
zhKEUjzhb2fIqtAqWSYuiANIO8pxAiFKKLVgYN9zTn7MiNwN6/2qu99ADbbY0QDA
xTD8GuUzYmSzg+An67VhRGnKLseiuam3kmvjZyzHy2nEEWFRFNE3YA6MRcgcSKeu
qJtbL1RT721QtbCwlW0bkOGgwEJr7QD0YjNVnLLW52C6WxK3NpweMXOodakAwM9k
IRYSZoUipJkVzejuQpNT4wCMcGt8O6/G9r5LZuQOs+p4griG69BSaSeYrHXkRKtD
n1q+F84Fbqw8skLD10tEdtRTOP+NUbIaOLzUblioPvbHnzmmgUy/4MklVyIdD6SI
8Nd3oKeoEPqNIxxILKFcYrlZgsaOVZ1pojon6eDBaliXFoqJOoE5OESFjAvX3Ru6
rFe57YwihURGYmYgYNqw0VGePofBtEiDD5DVweeG/B1EMn4gCt+QqvEDalzN9Z0j
1n0XV+Tu5v7Ebde83NsUjSbrFhnnyjE6BdYgvo5pV2X3KTfHcouvByrcdPjArVkp
/Wr1HvnNDZE9+0K5it0zZWeWnA0DK0Owv8vmZPvxaxJ/QGqonhbzGrWzATMEN0qi
ixw3dTzseEzt110GMwXYgg0z80qSLoJ+Q3XTEZrpmsQdpI4YolKiWZr6dL/K2KcC
JbYNgu+FTDBG/d5dd3N6X/DQbVus7KP8YjsInynfnrp2nQVn9tybZYiSxfCRKIXy
FCwV0XDJ3jX29xmLqKGD15rz9SjI7qatix3hc3NAxM+Lpgnoiz/655OXXOWPDtnc
S1d9K6BfFnpF3tXdaiBSv37r+riZk8y5hbNPwGzwVjPNR1nXNi4ygqh43lVhyQHw
dQ5q+5lVB9mb//VsDYBQdARGzJx6VoDitgb+NXxv9ta0K5fc1dLaQwDaUpxbVekM
BAvej34XwTXKGOvGihu/ja6DnPXISMJ0YH7mHAhj96nAvfgk3YVYCJ0zrjva6N3f
plFWhztFsOSkrpTOqFy25/JRyoBpVsGv8ns0ki/MOUTIIfFJk87GswbcZ9p1vOQm
lRqDo5jORH0ZM1JYBzzCtXYpsZR0K+lphokFmEUZQQSKr/2MyO17jHGxztGSDsKN
ELoV6JduWSgWxRlyTvsf0hj/s3lyLKZiPzZavQ/O2Jl0L8zO64iQI55s0MP2ndWj
a141wJpjR+lx20+6le1mRSo9EDS0X2RHugHExKgQ9N90j5EMk05tE8ZGuLPD1oHc
I3WiqxzcJ7UZGnJmpZleHZqiSKRfw6lUm+0Hl2qEB82e296LXPOKoxPDymnNZ7bf
f1D0thM7ZDFhRG4CNvi7I4NEY+XRRWQVX1WE1StEoa7NvgOgSIIiQVfOP5GalkXR
yFXUBzaoLgq/POKZ0Tpa0ThmlbHZNHFHQmKOuZhrpixn46it6ECzcJH+jH40a3x0
ZRuTIWBOCxvpZnlLt/5mE25AFleK+MQSpSFycH2GjLRtLVnbKKN0vp0NqbRwoTEp
TFjTRlC0LxlEJAFFVuoteJ7qC0n9qgnZyQTm8x3ymUaYHi8Id26Pcm1EFVXfDFUt
SyqdIT7Omb1pgR//EkRd75CVINjhBMiOxBBWJrsKcvGapTWaYgDIGzXbKyqokppX
ceKuvjWjpX/TUjwr+HYaYAcSQn0jHBoRLu3s0O6fFr0vQqEDS8HnWA6/PrUOvHJW
mNeWX57Ga6SfnJ5OgWmDjKSVZNjCxrWQusPN+LETtUGjZjTKBkQplbdVt4eP870J
sMa44AvYL8uISRvORePb6p45qiY9NIpttCUy1/LrCvxleUh8KpW5E04USFJvBXP3
jR8S8K2WUwy/Px8w34APQwsdh88Ub6Vwnn4ot6NUW2RwkigaQ8W2PNKqnXP6QvX5
B07wFjLA0v4uueHCM2J1UxP7uH+ShteRVCbSYna+uIX5RhtSAB2zqyPCqc3+WH1r
k84zUhZIz9x0Pil7jz89u/0b/8v9StjC6wHcmvaJlD6MKKYIVrfqVGwzxWFpMH9n
a9Ul3BQKka+Gxt4W1CUpJ0SjqAwj8SAxyksgkXi1qyP9rchL1ie1PqoVI0IcMmH/
8UhNA5og2QM7SiEzetGKeuuGuHnVmCAHJbAYCHIcHlyIjoC19DqMCQ+gDz8FoHRP
l9DM2y9JAEkbxiH+FNCfAXIZa0BmqbuNy5ivQ1mspk21GVcEwtWaASov5rOx7JAD
J1JZ/A3pKX/j3CzpV4rXf0CdXrtUlE5Mju7O1/cbzOOM/uzVBw/LvfH3sImj5/y5
ImdRb+qkRuEiaCm/OqYmrlIVLrYKJ6/lNzy7fdzg+iH6BpJN9JzouqLTiKs0QxFv
8CtFChYWkeHSpMS2KhrRXCNlglTvcx2B9DRbEBmXP83owNV5Gz9zufhB2tomnOdl
ylli69DdSYn6W/zp9ST0urDmaO6CYeyEBF4QFceERzf101HvB6in8g3Aze+BH8WW
dNUJQXlOZeTe1n70fCPosYU0vhWErtsdHeVVfj0YrvcIWROD1OGxbpzJye6ziptS
kR/aGTs1OJSd/GgxZyL3SpoL6B5Yov2QTOqx/ds9Wz/DOVdG1unIR1eqqYn7yUH5
pkqg32ib+YCDRf1DS4O+BH7zCNvUz/MzUktjApQPUAy1ShMTaPE6ePcnMTzsaGtP
Gs8A/hf/AcnpqWrPDdDLPVicluDO8pHGruQ9xNTIJhx0t96E/H4dX6A/Ttw0yLxM
ts6JMv2GkVNARhhs90wmohoEVayc2LykzvHdm4lL7FrmUW5RdL3pcMM0j5sXuBKt
aIsDLEGSLpWvIMJQgNGmiD6Itav/fZAFsePidyy3buIwWNLpVROo925beVK7awN/
/wT5rkk1qfLD/gQS0V+wN+ZeEE3225ViXR9k0kuNgV20SNwAvphQ/YEoj8h0k7ZS
JTA4IFJMBcbJVOWqItqnd59YaCmPaNqq5ZA5dQ7dvcEtYtSg44pCnIJzAPoJkh2N
G0kpf2uf2NBwEbH+ah9AY9h/9vqgRNU4d73q0menNPM0xNnz/DZOVe6pYBkWzesh
K4K6Rs7QoGBtsBZMo+QdBASwa/odzkQC3KX0UcuYxXTp3pmWzqEdn4cXVM5b1xVJ
EPuS+mlH5R5xh94r9f9fnLitiFuA3sTPsiO1I5bM4eqdQZbp8qlRfqELjbSHnct+
1XWJvIKC+pOeDaVHrLXBFOlz6kT99ZRFxOD9+EEwQrzVaGpm7ZIj0FKNkaztOuls
wfJfzf5CqDAiJYPK76ZHp24q1jqOIOzG3sqPVL0rxaNkrmR6+nQs29F+s5SyLQBp
LCWo0z57VdDwmMBlIaAvf2WLhV2RwuypEx6HjY+d600jTs48xM88gi0pcysAJjXR
xu0LFbxSEiTcy7mCOBbHnKHuoUoAIKG2qG6s4D73euWsSOsQpD8qnT/yxmfCUPzp
AtmbBKHz4zhJGf2ELD8Vgz4sqbjtv0akSKkFLpoOJtWQnls4H6+8aTNywSDmroxw
/b0Y1tX7RY0DxDh305N5ZDIyqO9wV55kCSwkdMzYMto6zORAZx8EP8A8rkGMYsXm
nMlsEdvuOq7mGUZztlF2cfZcGWKmn3P5hlKicLpc48WL1zafO4SC53cHA1Te+5nX
X7qUNQ3il/TTF7K3C7fagWG0q+uknZsMUWHA5iy4mOzWfu0qAhnCEm0RgzaUthJY
bmFbg5H8RTUNkVlEf5J8dxa3QxYcaMFMJYqesOf9Sn1rTiKmpnu+FdRIJmAbMzZs
CgxoF5tIJo0AA+caJKAFLGgyS/QhszYS2PH30UtjN53W3/BUvy1D7BCBmVtkwaiy
nBXp6nCpP/tzj7mE3UpYGs+7jKrJdNy3y/tjIXeZef0xd/FhuWRJlmK5LK79dHkh
L9mVuDy0QhKfgB8kr5IqU6DPRype7DXsXok0ycgAPYdzt/zB1hldIAf6oOj08WcU
josIyixLIuey1z5T9elqe1lYlzW8amMEUWUlWVBPCvFjPhFtBoq/sYBSDAWd+DVL
qk6WwhVJ+vkbDH1dmOxGDYsNU8nA0T70JdJ+kG6P2qjI/pfzrf9ZtbvCUdrQXV/v
0Gfs65VZpATSZe53pOsy46Elq8rf1Wi3ts2Y9R7rgjMicy7hid4Ti+/QnA3sg+VA
GOMkI1BD3uHI2gWy4yZI4OZmeDcfq4pAssVae4RcRn0rv84wM9TZCnpaJxwid67O
+GdnHQtIFFm3NOsSA0QF/GbmexDX1oLpIqWRS256w19Jc6IjZD2dJ6Lq3htfB/mc
i+4EFSXOb2PoLZoDVxABfnB33VQJlDSNZUmctZk1KL9XTDr1wxsk6FpWEpcKEAUr
BwnOxp9zeRkNP9vdoFqm+GSNwne4AZSM1XdYD6hyadrI2d208eYhghc6gbBUDh04
sZrAGWWpG7fX1zKYwJwVO5QyHOZ0E053Gpp9m/4zpac1rl8aDinOmRlCVn9hAgZ2
aTZm88l8dBpz8Qnp690bP8/E1MZdUX4mxE16BlSPL5383z0Sq+LwB9LjGj+8jEqL
QnYqS/AQYBwYThe3YFkMoPGLWsXYFq/M7++wr0kcwW2hR/+Gc8mZc+NMvXUlkE3J
5HenBPrSejZFcWVyQ3JvVQPXeqNEqiHGdIySC4d29mekB0QORQQhkTKSLxzwLp4n
Qi1lTKa+lPmv94haOMvVGXnoEyMYp4Ak8gJO56F2qzehJoPUgq/kHt35IAuNxttn
hjdgnqFFQFH8NjNLT9+1fEwAics8U6lxfvW2+1jLbhn4ZiOxz/TJWmSMC6KTR32Z
4BOCCx0QJBfLJ1zbcP6t9b5sI9KbXRTyRqSgwYKyp8f6j1nn9Zq4e0dt927HAwZn
bSH5k/MBXeEkMtTqVpw1VkLJ/LU2/MDj86Clsp9C9CkHNoTFDVvdSxxZk9MXn9Zs
x96ILht+oDdPk4KJqpSLPu70u31MYWPQevUE/9OUTLo0n8DjL4p0xU/GtNx4qZui
QJavXyBeQEVy7pOdmIRIE+3VU8mdRr+EP7E6xcYWs3y8DAtv82ooIzpOCI9SrtHv
Jlg1YgGnRsN0agxka+fbo1XDxifHZXc/r4l+yjPhhnouxIvlmFSxwzie9CJ7WTM2
Y8wk3hkz25AaOziACdIS2rPrCAbXNi/eQoFEDYr7L9n6kXmS4guU7RBs0XoXqaO8
5geoungK5/LrEaTWUj0KbR910DjAb7dB9UXSGrqsbgOTZ0C4LIBAP0x1Ij7EX2HT
9e95IfRqUsmGcQAnVP3qWBS0yyz+XLimQoFyGUX1UoW1lHOEvBvDO5uPzUT6+qQA
aU+dKiLlp8YvKXXBX416guIrHP37Aio/g/nZ2FqaUmU8lATfaN7Mpy8MwRdqGEs8
roXU3lRS4MKtjD14zyikreSrNLpOT6UGggqZi3D1uvmhBetsGXTG9zUDUp4T7HWT
MCF2QpOOXlxw39VxrDCvYbDg25SWv7eiDusg9ivZDlL1U+ngnwSnOvJbNg/lGHfD
YeYjKaVGCHEiC7xg96zVWMdfM+5b08jbN43WRvBOBqv723PnwZ/oWooIrgDDQCnq
1eI6UPlRctyrddbxUDtET9NwHEJRQgCQEW7HzsFJ5DeF9lx16J7KAA+tETFIgpXo
pW5sSXpqoAzD01ruS40fesDbIPGOEDZgEc1bghB2LnHSvzoFRWGBm7lph00G7yl6
kWVvE1ibeBuQFrp7YMPjr1yiatipYfs0yb7D3hLBFKgfGa588uix3uOanK8n6ec7
aXtwcmCT0o28N+nbO0mmKxjY/XcZCb8yS1f9I5Ayg42giAyLFdmkatkLDRUIvxST
PdtrlLhmEhVFgBBXd9XHcMSkJ3rD5dsAoAgSOSstU9bhiIXap3hh5ltqGbqMfvhU
C61KRZEW3MsP6Ajw42fF3kZdclH8PKiGAPvZWUTxOowWdAiW6NCtVoMjUb01Wt2x
dernRxlXhM67HrOTHn/H9jshGjxQlaQz5KYljaQgzTxSE9OahKLpXKbdSOpMA/1H
C1xImnutgsggKRJNaiy3BZX3baExbkIt24MtdvYL8cOa/HwxVyj9LxGH51yYluWY
rCET05IGvW2Ir4DEgnqq29IKHF3UrGRuZHf27KgpkmVYbsV5JrltfMZEUkp4cCLC
g2nB7XlyIIWRHENjv+NUoQ9BkhqU8HNHr52Z1ZNE+fiEomPFFHGf9JaR3x+V+Sbr
auDOk21VVuBRTweCWoO9zEfUfGAz44zwOeg76qEk6iATMg6cbLerfamE5Au4YcqH
KwPiXcsy+LBXiYEeOqo1pK4LBUXbIJPCu+r+ysIcpJwPNlTly/3E64p8F3buQ1Ur
3d/X56mwSuasdVJ7RxeSTqhujH6ZVVhj5GxtQKviKmt+OUUHsfRHj1jkZNl31gbz
he6uEttjFs/2eKDuwh6n9vmRlio1kQLloCUXFH4gS/+aEH9ZqpifCq8tVsOkN9pl
Lj9w+q9n+G0O4j2ndJJ1PQKxi8/bVc2WHNsnCYPI92J1XLXnjK0Zu6Jvb8+kEKo3
rSt8NBiJQ+4w/TOAcMmzlzxEykl7u7SFR4pnleRNDKbzgRfBqeFDjZN/wQnrud4t
08YaTP4oQj0xQymVSW19ZOhVJfJYlRhz6Lddbvd6/5Yj3f4PUifWohKBbWR58qUz
7K9J1BbGoCUxXYsRlkMUSz2+wgh90FbBX8OxPIb/DlGPw1Gdxs72iH1zh2a+ZOEt
keiKLCCqvblOdg/Axc/yXtR2ATrhb8KKL7Q4Ug27TeqFXGauTVV5E3jIlyF6ssFU
a/P2LyZ00NwNPfTo7xd47RjDgzOWUoJ0GbooGcg2XfoZB7NcCWsuiI06zvJmyVBP
yOvvFpBh5jnkSnjsd0b+Gglnkn5GYttQp3LyOdZ3AjrwnpnnbStHvqwOB71sOYec
4NEbkvnbrWY9JkmpRn7ohyVaLMrz1Uv0BIQjZS6ResqZ65LK3gZ0XA0B28E/iX6A
Ulbc9hKm1TgCOYQ8GXhuxjacEdL8N+bWjibWL8B8NJNelbid8uFQqTfEOvpBipsu
6Ti5RmN6gxIGTDmJGfQNyzoIYnD5MEXWhT2B5217o7oemvo98U0eU0Bve3tu+GD4
0GUXXgRMRFEG9RiN8U1EAWKTA3nEym3X86NNOduLM3tLSBrccnEpkGvkJycPql10
XRRDcyY8FPskHy7WgsGMhNiXTWIi451jETqNtRI5G/cxfT7Y7aKxPdLoN5Oymycg
UpSshAXSAuYzpq8I3SFZcXh0cWkewckR/020p+TZdXxg6CAE5Mvo8+CYrDFW3vD7
YvS3GIKkY7evUSxmD5+Xm6BrD6SQHFe2M5+hPiTtbNWFY1SBL4968wEnN6/+BueG
eeffQQuL/gnBzSucMssuzkJyJH38hDHyhynAATvHN2npdGKuauaWeF2/w967NB6P
2byoC/PRRBoRTmtVmr+KRjaGmVyrRMxR9Nors/YK/eIYyjt7XXk+weBDr5ERLcrH
Twghl6qpTV6Zhaqcm7dV59Q5UB7yQgXmvqzc9x1rW6XlNMLz1GL5L1CG+o6mhCPv
3ocQ+Z/O7NwHEnck7TERtWQNLqYtzlTMDw5dzjzJwkR77eULVLrVV84WLEjzC7ii
tDsmn2Tms2JuoP2vuFV6kjCsnxQAQz0wjbSwi4Ns7QaX5nUnbTBumkAgwxlbF7Lw
+RM0J6AFgR1+ODOVElisX59AokTVWCCJWJsAFzyfjUcDkSRt9a5DUKwSqflLxfe4
GG1aj6H3mBFNOkF3rGjVcbz/V8WpCgs1rAWI95gRi5zi0rohBfHgo9jwWsDeGhBP
yOs5zKhu1UwV6mY4LocOT/ibM06HSnhyPnT8tETfYJMF4SZspO2m2fGbrsfVElhp
HRCIbkOdU6lKtkxmaQU0swqvZQ6lRkiNxKOlQ5bmaNwq4dVMxbJ09Mqh6HJUUbAX
z5PgAEyMYPno/7uyDmSDLCY1y+uOn5oK4QkYGhrzbAkFK18moMKjAQVIUfsppMaf
0dsM8gGcZcHRBdSh0rCQB9lnzKAtdQ9x6STUqNR+sRvAPRqVLsPLJICsmrFu8q/Z
RkIZLhdpjqHWNu1SE8rQy69jwcfnXk8RrIvdLhV/Myxd3Dizdgc7/pjic7HlSfPq
/0JGSepDMfwT+oAk24oahCRFNtCuLyzVOFaEOKsQa7D13yFqG4TOeuVcQI6RP+FI
yU77Zg8eQCAiQ2g+0+b7LgHt5Rh8/qlrY1RiqCZB5r5qLYNdlYT2U+MeftVButpL
0XTN76NrseQ+zXKDalpxYmhiVCbemGbZ9vibO2NAH2I/AA5pEGDZ8afng/Kr+SWX
S3GL2JdZj8d4FnYtCti41ZELNvXO/4tdseev30C56hI7sxBoGAuhR9VspUpMqLJc
f4av2IF0j7Cr1EzEhwfwbSo+M2nWdt6oN1t7M70QVX7JEd9voobc5TUNWT9PqqOC
gyNoDX2EU4ow4yMX3VYQA/c+ip1N/CwOBjD1aM4ArBUqxWCYLeDbMnrAIM5PzdOa
cRbYqfI/JulI5MceSV8CVwp5rjnfqd/TvQ8Db199gvIt6uT6CnJgcS6aAjdwA2Cl
rm8Ck+zNdOFDdhmxwlPNAYZBj23RrOGdv73/uJldVjvNARr3ZhPEEeWkUUtCLiDa
RELj3PbN0jCtSc2fu7GI8sIQ4bZJ5oPjkVBifzxj/d1WtDBc+x3jRJLY0erkN7NG
n4ugTO+ZbWcSY+p9/V6ZYwBZkjXKyv7CDkI3xRfb1upHXko2bSQmlQwIAxvha8EQ
ypV2eXPZj+NbQqFxEn/DNlhVmur+Q5kQijXuxd6jy+8GeajHLjQbGBHSyg9Zsb+t
7oH0Rgpyr8KDIFPUe/jiYaW7fgT8/KNhVwrViJTOEIGi8jS0S7T/vHJyy2XWJTP+
/Xf3bJydTd0uSN2/HIJvdX9XQBCDkOgtuHhGpDyBm1hiBfQbsWzc231K28mkLEyY
Q0QhS1CmqhgFVQkytMlVIACWF08CmXJ04d0AobjBw/wjP1tRjXVPf28fLTKvr3cd
aa03HfLYaAmkXhmp9pXGM1SLRIi4QRfMo9uEtuTrUAftEPW1sVN8xGd/hsEM/EzJ
/C068oGvNKabPw6btuj6rQAalQxSgpd+EMdnITeGpp2t0zflwJTPvSxZ6Gzp4712
WZMHQsii7UFotH1xyOiCMiLg+T+dBHpZEjS99h0fMRtpTsYVjP01g0uapwEiV0fa
aVHGaiNe7IXX90gkjDxcjPrg+84EB4FNYGgX/O+NGMdgWBEuR2RzD8UZlFfCGo0d
742FBN8QKuddkefKZTBD1TRrnfDWONdfkIp+9Yuj/1dI238p/WwoKoi0Wlxk5V2W
EgOBTmnXiVF9eyT9/Vxz/GQZw57qw0LrcL0pGnbxjQytVQQed8XrJZRcGTiATg9P
G99TdrzhTo+nhqMlDUn5QXK5T5dEthrrh4Hq9VsX1Jl/g43Od30BYldtY+GzPAKq
5u+NLZSAZSsANH5hJtwd/awpfBCAZtoEXoTr0wn7m2qLVb8XHzzjwLcrCQoRb9tl
U3FmUGy0q11865IiUgDzncmsrQ/hW8qq+SHQtyZM6L/GOlQ+hC64VAGO6/cfg4Zd
VjoOvcjYJzqAZY2vuXs7w68TbtfwTlqhs1NfvrJRHhafmXq7eYhPVimzEW4GxImq
HzDaeyS557i3z5lbWIasBluDCAdkTpAjGB6jaQna17D6OaT2kT/WpqSC6pI0/lUO
s4GWdFwtmWPDrDS9b4ukORV5K4OnnqtvqBdxxRfeEmTaob5Jm89TRn9gA2zn1YNq
+2CHbPvH3gXyiXwuYCQZzs0mxT4F3z/fgUOQApwtYa9IuCz+HT7emLKh+PfJBfXv
8AO+1PxCqRAhar/KabHpuulgCM+nNknQ18o1NopU4i3YFvd/J20lVEOBjbpACtch
kSRizILRC2yiQj91V+aD+1dYPv0qcSKAQ96vLLmR3XHHD/k5HNYFW/ukEQhHyUwb
fgWgcBAPwX3Ebp5I8COOCWOH5nnQQNB3YfcdKBSP8BCN5gkj5lxtAAAH4AdAHsvj
8FoKcX839fl5+35bkWeDlBBvKkVD/5Qm2lUHzOUj5PkN9sIdQ/swKOy/7zHnVw2i
ZbONGZ+LxINlkD5r3+IHZuCM01iVot0UZgXxW0Mpt/7xMTJQFU6TwFIya8wNJnVi
q27IcJA2o5rs2C1ESyPLzOXozFaUES7lwuAbKf++qbGCGAlYT3k0KXsRRCIwkS89
XtumsHoKRkeoJ4jaoyWYsoA8x8To74NcGivXou+4YHEmGpjwdbB34t8BOdEwJ1Xp
2O3Es2dq8Khcmh/K+5tEGBslHz4AMh9LgJfHAuKABnd6HMDAxm48YhnTQFdYMWWP
a8K0lsgRKaRSiOxxl4mybJQVRucv7ziCtmhD+mdXKZgFxjf7LKC0lnRFr7CwiP0D
M9AUIR7gZB16L70ipBrJhw3KGi2PpdgPEZPgr5UIzpegtcLGAjg705poe3VMEdkl
9VWPbEsIs5f2kQpP9ekIRqeOxcvR07zo9CL7zdVqeg2qPT4hE9MFc6yCSa33bmvM
l63YpSp+/D76/LUoL0+qfTIflC+VdAj9J5O/7+SmYGOu6fy6kDr6vY8/akSnOani
rV58aMHd9ylQlHt1DoCDXmmaErKpbIkAwn+qeRzrNdIDzCldnDCZYfK2v57wuslN
ROmF1ixC8/KZmObSC3PPBB2JAc96T8Pa9j7Krc35Ut8DFdNrLdaXwHeSszXNyRvA
g1q5+eQJRSghVbyf3kES/Qvbb911/XPBsqEed708koWw+mIAge+gYgSef6V2xNdn
vUI7lUBSzMsbIrGp4TleRYcbAwHYWHFvVxOl5lnsbyFos1KoGeOoVhlsAj32J4LU
ar+NzIHhl3ztJANOThOl4zL1aKgzzK3KcV7PJ2IeE2H/uRbld0fO7vbZxNdzgbtM
tacwqJLDbvmxCGvLTy17f7YmNs1WKu3FOABbrSJLvwiQsJmxG0vwj55ep6CXsv5f
39fDiPYF/vkHLvN7ddWKd7dLeYMiOCyKzBPnVVCLXPSrlfX2nDaGkrjqnUkQYTln
AdyXaynV+Sp9lz/m9W0zhDS2XMmSp71/G5oDq2L/tqnsmpvmAaDtP+mOgsLC8tRJ
5h1liySyWaJ4kUAoZVFDZmED2eAUamAFhSU+KjisQXDyldfO+eh+MF0JJPLwWgnk
HH2V1hw7fp1DwmPV8NuVj+fY2UofSw+BqjcT9nh9Bl5OUibfy56Le0J9xQsl7t3+
lIqjG8ydkMRXkFJKlymUfRfAtG8b4iKx736dE2fKEbJ8FqOVdSsosHRXdHPLXlbp
hjzUgysucfj+np3zw0x04QB5jpRr7rRzUC+1qKF/loCcesKgB7rXEHdC01Ur9S9X
0BDoDmDwdyM2IOBYRuL3qdZfuSUPc/MfxCP5JSpQbMe4zTefAVstDeN5NfjhuZXR
SBpBaeNwqL5nI/sp28gDSZTn+qW1/0yCFsjiN25xKVPHSLUoCdiq5bm4jTs5PacT
DLJRLazNoCYnPvbi9Y9Wt44nuw/x8OLh4SZX1r2FYIjaz4bEh/SEkgVNVCLE8BzX
AIPaPhoo6xQF9aCqcvDidAl5g3cJxyUhDIp164WXl1Wz+qHoKfGRA8WPjVndXHnT
cpe9BCZMp1a4IH56pnxAzx/yfvqLtl/lIFj/O0PMR0J0q3xf7TadY1r/v0qYdk0i
dFaeD2TEvZGb+mmixa69Tg7roGjQDAQELfIoX8g/bfIgqHuC/joo0M0NSrIT1PLA
ds/Sa6ca6SezJSn9bL4D2ACnoTEoPAeoYnSQO8IdzARDiCBVfdOdiez+srCATIuw
Oqe/AxJVfA2VWbDDp4WJFMDb3tYsAxtwcCvX3M2Ux1U9lDz+35FErBvbcV4PSktO
DHEBNifGBTbVSYTEPu/M4YJObrAF3ZaimLr2GezwfruNbNoI3yFV5MktKn9wEaqv
0AH4Kgb8qSOF4W/6xHZHLgCQ9Z+vjjh+x5ZUCDU+uUbCBlGHiJIip/yFf6po4Wc2
hTlg5zO6h4ENtInJf9zi9Ve5cthb0Zl1EL3ucUlqG3w7rUKWHmghmxJsY9ysm6TL
uZy5sL7Y1ME2SLMoJkOL5ey0DaQ/HJv3bIvTELYzJR88mQwS+s+wrCiIKS/Qrdz/
SsLTxrScObkaPXBqwxQlTPhnFj2JUrPQncovt8jZDseJxVvsOcsmaorMuM+B33PC
uXbmbJ+GRVodBNLgG5uAlJyK2PRBGjM0Pt4MT+Gghd4zUEvamPaDT59H5OG7NPQR
bqP1X64Y47iImovYsmFUB0LI6Pi74+ThCUlnzGPOdOeu8TNMevHnd0cjoQ0srQEu
IQwfF2EY4CdidIQGbB+Ptv9R+dU0A+fe/H1+B5Hzx1awvdUCwHUxLZTcUpj/GMuo
S9/SS+G3fhVeUls8yFZRUgNVdwq5cQA818ZdaWUnXIUgVfle+OCDc7OcyW6c1hZ1
g7VhyZocuDToNpLGWa5GACqsqpi5/yrIheW9HrnP69ljV4XV1AJR4wWVBKtRVwVZ
Ac63FQH2DXKzVVUcadODDE65efaO5MYT6tQ0ogSKP3ZVIMoDZ1HN+JvKXxfNXswq
gAeHwlpZ9ccZ4G87kqY3ALmL2M0WRbAKp/4XnFeVS8vsJ++H1bmbBZ7lgHRWRncV
a9aX8E+lsasGQzuvv47mRxZZd0gZ0v6bLeSiwxhajZcy89UGQx3RZqoDESEffTqs
2/pmYyrWAX/ijh9FzPcltR2mGmtVFOh7ek8UV9lGE5XnxSZ8GunuOSiwwQ6vIHgS
/YFK6KyguMeav5lCLzjeSyIgvFaBSPgEixfN5J5N3RAjJyGL5j864wZ6q/gLBF/R
3oJAXfCyzxlosfoDgbLuVN8BVDynqwUEH0KW9nYvk+BWewCotoIfmi9MwmJts2Xq
YL8YqCtFIwc9/iyCfQFCaakcsrM4SZQRa6Zje/xTtPf3kqc/F8Bp94dcQT39wUNB
tPBOsy9ytRUfp+ktfyV6E33Uxk1ohagxR4hzdueZZgbi61cyBAZCJcOPax33Csrn
jC7aQiBwE6v9AXO3vxk8LicWeh1PPqWAVIn+ao31oyTPIYFLcOE0sfyy881nkWLL
L/EnOc0H3DDTa5IWFdc+Y/ugp4udzLpYfG9TjYymm4qujHkXvlGpw6mO37HR8uMN
jVmX1b/Zc79m+AQJJwdDzCBh9RYu1A73b9sbycCWPyzpZ6xrPNNNkf2uFnapT9IH
gx2iJyT4jbiN31udf6H6o9US69qOYxt1u3N+Fg4lRxSVrvZvNs8Gk2OLUjm17JP4
LyZCdglI8ZYdYHC5UsKorCXn91xJQJHR3MlhQrsQSsEhzfdsaXOSlknc8kseSuZ6
tBpH68O+fxhLm3EQ57/1KhA+L56NEerZZPz/CqqvdS4Am219FHZGsgJQc5ylLtU5
OCQhA3LRBLkIzytxhv3UL7+f/gyyi95VBCKxLo60/+CHdU8G5oT6rzrNe3nisx0e
xCNUJwp1SfbNlOoGoLbUf+/BupQ3EhymB/9M9E3dGYzFKZE7wPJyNTpOJvWwy4rF
myNWhZOw9EZNlzkAqkGVO8OEOgq6ZbIds8ihSMoPeORY/fKECrnayvVw9vv1f8zv
5imBBeCwiHNB8vdjX1sbZPGgdo2Yk//J9mjVQM2VTVsGZ4wts3EJjUbE86bm0Q4Z
4ZIfKBHIbEU6s3BBZm7hIrVVFR6J5oMV3LUubOhe9B8GupDage9XjW8rKJPDQzUm
GdP3qpkvj3C3CStG0JhM9fF0KOrw5jQpYS+CTrFVgZeTgQqKNjUhlYx6KI0Kfli3
bk4Ssf4VoPhKSvcmqqpEZr0Oi+atd/v666jQgomNMVFn5/Esm2DRBkCJIejDaJCN
PoujsFSUsLmfrhchIw4PZ0/F+kptn8csraJ9fRAWoH4LQMF33D0oGVlKz55apJi4
o23xigfRfo1gLuDIUlfJ8g82ILT5uTyetJ8eXsWtujQVfmtZcTVQ83U0YWyE9pB7
v6ZYtiznv6WxKo+GM8e5RFmnffsgyQqFX8DfD7U4eoUNdBd4XHL35KRQgi4mYEtF
axagysRLMUJh4dFwRgmQqcadQj/bAJ8AW+3SjUKdhjjKqulKM4pIeY4BAxaPAQxA
MmXihTSG0wzDJGFVqaDCB9BiXd0Mlc+jnHZOeJXDQchCVON2IO8oNZ83ahDKGNdT
m4ik/Ml45hE6kEb7AcQcI4pZvzn+XX2aGK655CmPVDessf+fkSIDLBMGn6MDWLD9
fU8p9g5UQk5WzhR6vtsLRJS9NpXmvEWkUI1ZiA5KGdlzr63PNG/OBLowx8lc2EAF
Lh9KcYPJNOVdYblZgwAF9N69GOrfYseGmbGw7+EuVXBulntn+o+SfxNdDmWWN04X
LgelM625sJSop2/s6+EtabTLrlENU02E3K0PSUIDTmxKlExdNqtV/kByx0H23QVE
g75CjWLeEzzwr+ek6bR4ni9vB47Jw22s3jOy05HJC6aqgqU7dvHA8MKVnMZnkFq+
geppYhSk7jCWRUsDGW14YIZOy7StzjmcfyPe3XckCJfrZDfJj5TgGMvNuISCUM1c
1xAYs1NRC5bAwOSIDO1pgOvMBVBDVAowwk1O6nH+gOcZRbmiJiyI4BtDjmpLc0nT
K45R87QOYEQQgaOusdGwn1QVRH4mlh9M8LlRdtqZovtBjnpmQBRsTzmEVQucc4/w
wTSJcV5BCXs7BmPtLuJZcQ0x+bt62JV4TmUE9PaRu3QhX5MCsVXkmbuayrXUBN4E
on7abFEaFTS55kgAPJv/k9fnInXfuJLaiXHoTxPO5WlLfU2vRAouA3YBY8xQRHaX
MX047aiZjOIYdaOkHBE2Sd7FbDiVvlYAxMQD/KfMGbvDlycWCEEEptLJcpATphbu
O/aUiVreBKLznpIPRw1zwXC4sPgdzB+BiCDkF4Gzj/CmT4Xu8+Ldv9Tzvu62EDR6
iRIEg/BBYFNZe+E5YMum/74OXPYAOiIGTeWXAxXxcUd0O+kDQYd/0w+MBO+TViTz
Ocj/O3sdKZ5jN7qXb3+8bCh29sTP3B8bvG2S5If8zYI++QQ1aBBezXrRhhC3pbgo
Gz/yi4R9GWnhh8nHQ452cXzBfVIjiy4u41hxPqf1xcLUWdN5QWk1wlFBSC7RhRK6
sN9BWpS/Hf6PN8SlHdPIbssW/AyS8PHoauDlkVE0Kwqw5eItOb59dFZ8IUpZYsMl
+9zQkz/dFR3pGUHtu83M0Ug7UpcSo4LPgl2MlrVMCo8WdIqONSkNAOpySoVBoWtr
pKz+MS+fz1DTh06eMNYPSJRb6K3iPtPjJ37PLFofP5dClYZCO49Qvtz35EOsGCP3
CXwt6MCscIbgpEex8578Zx/ls8eoJOnpfK8Ld6LA+Mv/O8q9dWYqg3jU7MR24F/k
25Q2tHhctBMiqM1ZgO7q3T3v/IDlW/zNqEPNfl26/alpv5kW4WxAz3WRG0OB27lj
OdTKKMSsFcJKPjtApHCNv+xqEsz0CyVDz9Jr4kBNADBLeJcZr7NcE4/RXHYywfSb
Hm+G1leRAYyqASQlTAuGEDjvuu3u3zgxIkm6c9utYxndpxrI/kvJt+iZ1/fpDar7
EjGMZFynnSZSSRIlUYdImJGlEZEhgLTThCZjDv7VUB0xP4MiFI0cKaZq6zjfy2Wa
/HRbObPPKN2w7Jb4UkucuYARhAXFnXYY3RqfZoAcCqtSNcXD07b8d4ucT2VbIx3i
ueyUWWK8VdKvWI2wI+OvnH8lHOpSC9BbJEDwwWYDeAKhYEEPSjf7bDRPr/MNA0qk
F29Qb8dPZTGlL1+lQoST+hhoiRMFV9B5ZdUa4gOTNrm6Oh5RrX0fuSs6Ac9lPVvc
13hYyYPCOe7XkHMuuwnFh0VhqSrFntihw7onFNixMSEdWbpC6SNCVZc1mScKX2qL
nlDsD6cKF0Job2COmgwZZ6DXKH38TMqe39Lv2OAWaiEuPwqLjmnVK7QQYFJ5V0tO
J074Ql8gjM0VORwVmOWKJ2oLbGLUpiwKnuIfYO+H0caKG1gX4ILm2EFM4OfkvTap
gQwFs6tGtqrd0RH9/eb2Kw2lxnWfaTBu2hCflliLPDy82blL+81sFR5CXb6rmeRw
zJxiPlOwzuAvdlP7ANfkp1eI67loUJqjXsjZZR/lWSp2PlChJ0CkLnF2iLQLWRJz
2rz1DTSRIxBO4EIazm/Bc/IFImj5k1UlguaY6SVs0XFHrqqvaNiyUY1TXoc6N3ST
wLit625iGA3nIneAxNm9sVPkXEdgTzi7kFbqN/dCVuEDNDqXYXDe+PkYb9Ao/Quq
PAgsRnzRj2ZVN8yukeQ1K6dQB4OnxEfycYS6N/TMZCrQZ21TKRjUQ6D7PTfxURcE
AZ4qryh8ZyqVHV/WSnaIH1KXmnN2lqIFuMYR6bcHpm5Sfa9c6PpfPYRq1IJMGOzP
c0IzHmebNufVR44i6DBAwQSiw0CLER87l7asPm4/l68DdtNuk9xq672dZWyGCcU4
K6Fr1su1QGHJ9FaysSjXRvzOev8lVrpdd8x3K2XOW9E8H6P8eUyAt21Eo84ZJnq5
4UTIx+5F9/rP2kbT33llvDFNVX9a2LzDWv2qdWLwhPth7H8XmGoiCrpWXwHXvzUw
LPWdmfs5k26XCmFEzgnBsyUEZEWdV1iPqw4L0qqeKsOeO7TGWOmx0ImUR8qiHArW
piV0QCXtIkPoYrQ38jz/UHLNiOVwNrLpwXbMVaySmHo6n23rcgY0U+j6/esX0Iga
ZGgmh0NNKmhDYcjpgL+djxk6xTUofcih427f0DX3F7EBab6onMb+QkJ2Fdlgy9EA
P+BOr1+lKE9WHqhbG4aG8yq+4eYZJHIPz0nao9D7qzS665lUUn6uce+3hsZXldZW
nGVo8/I5bYU4h11wzjg45JrXJQoR+Fx/Sj/a45VKXVdTmoNSPvBTfxn2zZiCtzOF
7NotQY4hd57FC8OHTLLyXJo8xxT16vtaAJVW7bIOvbHOUUTYV5vgpEIXrHHs8Jbf
ufTrviK6b8bbdXehpCRogo2A4z3AidcLTI7omGkq4PyA9cdQGwHnCnciYdgEV1oB
akuzhcOZm8RjdvXcPOsla0vNRt2ihOerBBoflNDA/FoV55mQqgkePd8lC9YFRDTA
Zs15Z+a81Aq6hWVn/ltcquUVWJTD20imMu0hrgxoEvJqhijIIKIaHRhogRtwYedJ
7wEC5c95X6QztznpUzgnfXDUOO6lyPmOFxaab+zQE8I+odbbIvzedhomPdhbDZsw
lBdkU2xc6jCQt+GYt0nK4f0CNNEFI5uvlCcCmZSuB98NwQeWO2f64NrBD+y2qteh
D2+uZ4IPv/skT5LhThmuiwTdsnt5Dp4QrVo8TqYZvdp1cRUIIkai9Un/n2spC28p
9aK/KgY5xCdP9ewITAzN0nLq624d4lJV9DtG9qBFGpT1hltDzPrCR0Dg817du8cT
V1tMADnk0p7mNNoKOBgUJySuTIjyM+XqrTpgpqHqHFnzf9p1D7jB46hyRwSSSdh2
jAGVu0sSU6INlgPvMGXt4zzQIuHlS+2Oclhw9zbTNfN3HUGw4IyOGzFzZnVr3boF
8xRtvlPpmcisfFbmKWMUW04NFUs1hmIj5kf07q+SBYcB0s+g+xLZOtk84OW+NyR4
bSC1lZbuW6WXnxAE8UVOLRDC7UpwgNyQAAVmU9uOHzcDCoyCMF1rYeR7CU2Eq9BB
JG4aYhotmj9YoPSlt1lZmG7U1WweyRwtiOA7Z0O7RIPxXp7RfKfTHysrTbddcV2g
zsSH9+eSeny4C/3aR9Vycxj0PRDjGUbB2OJ6nrpe4c4Po/Dvem25EFZbGz8WQol9
3AUsb55BXM+MYYNHEVYX+easflELzLWf6qYUT0xEpCva2/VrejEauDZPXRoqSHH+
Iu0By8AzFNDoN30zq+V7oidVNWuMoKnBRezMF6L02ExGOg+rVpEew91214kmDURB
UR7NJVH8C1GyZdArV1g0ZPRDodKqDq8bGJeQ9Xx2v6GDupk0GxsWgQLsQBAR97IF
LkzhqWntIMUeXC5/4k1vxZNkq/+OyMusYsOBBCmEiREfd6MtmYDonTIFaPQvewxb
wEUjsSkehf1Q0djP1TJBE3GfQIIxBI1Y5y7DaH1e2TlDGf91JI4ca8h41jGMF+zM
RAWU6TW0Tol2ny6RlUz4V6n1+qrGOunRYclDj+p/kMxZaw0j0dBW7U3v1eRLBWwf
1MC8MEjBpYKH7sFtBTp6z2O8KPJmKxUbXHRikYyJ2t3XPzM6FCxC5ScFVmRvpoym
29aXc9Ue9Y68mAdSoNCySZHyOF8Ut0C+jjSeJlRk6rrw+qDYnitPQPu4V4I/7QoY
SNE0OBGMNayamtNiRXZmiBU6L9JlPZmavR6Jbw1MzngvHqYA3WR4ddCdqBwMNGsC
Qggv+1m/kTRHqWBMEP6/4NptdGy7YoqfJNVgHKe4F2k84dkB6xPFe1Dp8q5cqwXR
99CLZerOL9Fw7mExasv1AuvdjbzRFwSaVoU22R/kDXRq4ITlNbhxuTbQ1WzXoDRh
6CCAF0spC7XqiGQF4exprDsnk3lI5ecw/BaC3N4BjbNdlYH4FMgENCwCcTCzLCM7
89lPA09yaek+nyh4LigBvv4m0Ik/lXuiv+fn+Z3DdWYwVetLg/QuckfPLRhlqgVj
I6B3W0vk2QUzATJiKmgmBp8gm2y+KQNeB/lq9y2snpodVGgP6e15skXucj6limhF
qQVSnH4rHh/empA2I7NPQSOLv6bmmih2/k7QdFjWpcM6pk+fdskSlhxButSFgsS6
a1z4cHrbQzwE3INmWNV0If3CzY1FstsCuaGnz4WM3WgROT3QhS73L8MRMsa2qxsm
x1Fz46c/8Gw6FdFKs7O3cVl9nWtlmgorXcUSL55nKnEagS5iLCw2oa7BoLNTFUW4
SdiUBfL0VVO8lIEP5G5igK1vc33av06BVT/q+/fsOY6nA5XcoOrSs7nQTAc/ctI5
slNtLk8YABGLZwnCxBuryK5dtKwLeh4yuwSBlg2QkWmoP+ZyluUUSO/889VdPEA4
wm7uH3CC7strRpN3L8dNwu5p6AWyNgp/jHZEm2XYpcJKTOWjynAFWae8GRve8Cke
AF+HWi0Wl6QyPns45Ev2xH57QZz5DLk9jq1CKCzqAhSWM2Ymo5S3lHtlWTVXSze5
IOercwn9Nnn0TBUTxerZoRItgmRnpfVA5wSDnb9vZUOl+oToWVQiIS5W9YeqEmTp
q6MxVTP3743X43EiNu41i43GysFyEve/DHRWcqqNEW+Efet1CxYzAUSlEkoe4Hm4
rwhC8RIK3aoMdUQSkT3H99PL0jdJLI1TQ/t9VHJV0tRUCJWl5XGJaSf8I5Ndpfgi
nS6UBD8IgBVhGpADYWizlQOmc5XquW3olsXcYugjSbBowFNG3qTNKOmvTknL65lE
pBpOeR2rY00YkE5xSUiX6mrB02oVImG+PCMeMxkaOvsDGE6JYdZM8gnyS7jPwTxt
huqOY6LXVHXHSf2L+zD4X4gErHd7tEtZJWC1UxXk6GCRJ8ZS2bHAqM8hb3fVuaDX
ajc+1UDXTxng/RoIQNUCGxkKwcA/tWGrC3N34xiKT8lIwB0ecOBmEARPEvHUtWn/
mzKwP9UBIe3/zh9uzn4lx0qZDIgIE/KD/iJyI3Wnr+cLKgby+MpGen/uo9bIj3IL
Jb9P/RRGJEr/piUrfNBuVBAp0eDzJUvxTXY5C7lyQCAlLxHA8gUpk2nmdfCuLU+e
ogL3DRcsuyuZU8D+vNT/Y94tj7VXXTMOJwrSJ/7X0VRHc4wcKi/rtrzrq1WYXgou
hsdoMQbJ270F3F/GOasmWFjf+59m2zAhgRAFA8xXvgM7y7M7hM+hflhTdj+0n88i
DBo7FDt0q82TXaLxhPNLPsioX/N43YITewVUCS5SwcpArgN29oMGb2pIsSdNA3l3
7p03On7j9fa5avTG7UQG5DFwXIOhLv7jhz96lDNiUMhQs/gXZMVBvhkjSFQISsQ1
FZB1gNdFIGJVUjIOLdElVyKaIRH535PF1XdZ35KNgAb4uDgVjoUhPlhpvcZKBY7i
ffgZjxrl5Hsi4nP9hvhxxzd3cfIAMLu3vmyGxvBaRe6i/Wthd7TWgLu2mTPF/Jpq
0+6OsUjv7OVc9uzTze4K3a7Frhs3ujuSOLGhmzsLN5d4Vk6KwUYLsC4H4CXdu+Mv
hoBem1jnQ+E/InlG1bkppqRSqvJMPv8mzpDfwuQKJVu+lBCvLhitmeid1yf7KQ2F
h9eftptLru/d9JYjrkUDFcOAEWvi9g4lmifCFN4TmTIYtWYHz4eyBaRjbfBMU25X
mK1hxqqPl6pDeho4dsMDnvAgcPsl+cXOmrGF6pyiSg6y/fqy+Szer6RJDARKL/u/
WEtlStJA1gue0mf2OOkxjn7l4iKq2nkTFusnT2BFu+FoniAYpN0f0l3sq4JabZyP
qYIWif0YQWGo/6r4hr5wUsfoUJy45O/8tfCLhd9/R3ieLaYxKdTV2QcpMOH9HGgv
0ifXIuHIj92tlHxD+LkHlV4APbyPDnKjs8ylWSUB5ONQIUxQYHpth3PTDAQqiTo+
qos05of86MQCJIZHQWdcDYeqMmqm9DI2OTTU+qdgLtC9KB9+pTpftmvzyVG9Lhco
T/yBIdT5465oYGQYULQiNWEKU56XLceZyMC70gonAlekihgsHTskQcgmerhTnD2i
XK3g+VFkTyf8TexNm/S/9D1nciYjVP59t231jVUJ3ENRcuwXgTQ3KIx3KAXXOxmF
KgRz8GuRKhK9eAMAcBVd0oKZ1alvTP6bdIMS3R0JO6Nr4S6KVvtcwbHYKmC4VeRw
Ouy92lOp3teeXkjaOMZ5JpzaJXJyKBvVLB3Hp86gVgo9m01VTL+CCci7dozmY0HY
uLUe4fkeDV3PZvR8ZIubAq0M147sv+SmkKK881rNyVLM61gMhhNquo+AYI5QNZza
lAo+UkUt3tClpCWouqGyB1ri0gf3+bliNGiuBhEh+T90p8q0u7Yl+yHhxPVxz6sf
oM/RE+QnWY6co/kClzWjRqM+ynP9vGJIpBBtBVeFkL0cHYWSxnGXI4Ls6QmHNH4t
hMb4bphrz5yHhAw8usToKzEz0coX9+TaTkSIp61kDM9ZqQTWLX2Iwww+eq1x2b8J
+YNzJKj+8MDsy684bv+nGq/b/GrGQ1OoW/SxJ0Zn/vzyBmIB1APfLITOt3hH/T05
mKqdewz/tKIp7+luEHr4ntJvDpOK/nzEFRhKvSEH8Usru9sTlRdmNSoM/Fs8rRDC
HAbJuVO0uGgTstifEOTS851+vI+1XDJ6mLBCoE9LUQzdV4MeskhWivXUYoSl9HDU
+so0PT0nbwltGzpU/ICAJbRqmZEV8NfbraaFz1Wr5sfKgDdOQH1Eva6FKqbzMrXp
EWhoRD+xBh/cyWzsg+LjGq0FsmrYwTxNZwIQmmSthcXZGAXMlhm0PWQCa0EVbCFx
OjCQfapK9pg44J1mDYghLOzBq09lND7MtnXRoK83w5qrEx9ek8NH2B0vyhZm9nUy
2Tx6Rul3WKhNzTff91RDgHzfUZlkvJBj+mz8/A1ZYXFCI/I+GMozZHm3FvLZUZSu
23wrQnQxRbYZs4Z2/EHgsYN+QoWGYRFc4kDFvzCul3ikaeDocaDnoLikTp5MYYWy
vyvm8lKviNVwCirY3QATApuRBYQA1VNhieN9j6l3z1uk2ALeRZr0iFKdkBpgYKWI
rFvOrkclAjPo30uXfXaN4WCheJf++oiGWbf3QcZmeowvXPhDrSlYp1HIctGSxASm
HzMUsghCxwheBmKI7bV5vsm7MQaKds+a9rJKVof+CluLzUpxLMBEn6pa+G+7x2ui
BrILzreeLnE/Mu75VOJMlpYbVoMgMLO/qw9bbU9vNX6DbeeTX+Q5XclGIDj2KzmZ
FqzOEEPLT1Uy1wO8Tf5nJrn4yicinN8W/F5gGqoKKrzR3w2SFl9jvcraYOoX4mdQ
ViBd8jxH8J3BJl5r7AIhDOpWdoG48jomx+/lTQI/KZikn+W8mMrtBtiP+VBcJiXq
YhUxPaOyxNXNfLGAisitjKc+BIN0+mhJTu3e+5lmpzennK57M7eSYRw3CilcWfzo
DvXMMfi5gduDyCaIl5g7zQvZqTZRTDmiEl+qualDNEl0s3HrUI4iRixnpM7RpqeH
cvx71G0VmXERnDv8xK3INVDVzJTzeing11aQ2fYnNFsRqr9Rb49CbZlIHVxCSXWL
wm6vDM+3Rhmr6HdKKfR4y5IU646tQZhRmZR328Tzi4RouYUR+QvWjBwVxOiH2zO3
4q+flxuVjF81D6vJOq3r+IkhNWnbbEIzhS4rslvDccdCK9/eI/2ymw7bjVJxUiVg
R8Ij6PXS7RZdwfxBhaA6tYgZjw9OUAO21H4ycQOww0PUHThR9uNC5NvI4smyDeX3
hmSDN81lJlRo0BxUmvcBmu7es00YZJySp5CBhnn/z5UJei+O/raG60i8cCJy7wuI
Gq44McdC0yQ40T1n4ohgeVX4piJQu5uobm4FyH3+2C56nJCFyvJCFgIDfyFf0zFM
ESHzUxMvVPOt9W6ggKOfh7BCne2CvW99f84C6Pt718pM+LfV2nGcfFarJo9m7I1N
K2rJ9Xn+S9VjthBLTydeX5Q8i/pmHlss961FXEZyLcFqSK0gL68omzsnbarivhpU
hNZ519fTiFn1BeBaC1UilbiaKZDgMXVSL3sfpR3065G6wTWfl6VIeufuMWZWokBk
lZB1qNsSJo1dYM9uHR1d5p3jbpoGW9vjhx5Iqj7qaD2W059hXg13bQigJjdW7Nal
4a4gxzFup+HN5flY7i0lt5g5Std7uPvHq7rP5MGT6Xip2hYfNqCHHzN+9mFjOBZ2
0Y72r0ez2fskMqrls1CYjT8TYL1fzpPANKv7sTEiNYIQgqGkU98m/2+tZGUyWnhw
ftJqCd2Es2gHBsXKY4TdrS1An2zjbQXCNZGmD5jxSOREP771ZhoE+T/u9Ipw/CV6
njnXvS2vBo6NaJcdB/refTQ5TwJYzsPKSTD46xZoBj1iek/SwCrmmREeu68EaiQm
Y1kCO/EWRG+UoqmlydaqaEZybO3LnguuTV2FT/K3l3wfa5nRuHgCdM75Y5YpK7Yx
g+Abisd3xvEbIdDK245S+DE5g2d47zseqTTACaeS+ve8XA3iL66Pw3rGGXvjtsrT
GWhXLQEmZtqD8ZqBqSR69BaTL0h7WzzdvTHEVYTOITHMZRGR2Nrqqk8bN3HJf5Xr
BHv0i2UUjGLN+4osElJwR63DM3NvB2U00tQSfIv1tuViRpY2G7uVMeU1Q5nv+7zM
DNjRNGrQI260EU+vPrE7d+lTsBoV0LD7CGeeqFIRud5d7N2mPDjxUa0wJGFlFDl+
996RKH3cCGMB58mTlI5Z5YQLLZ++CrXfTUdRNBm49impazQ5ohf+goFtdSQdZsAR
RqKYvP+b0UsOdP4NInncvW04X3f5iQ2GcuvgaHty53SqPsUFivlXUlTwEsXuUqyF
kp8/oGBDCVCSnCCQ7KAdPfbu101pVLtcM8niXM4XIcBxxQOTUJyk6KYK9vDRSoTl
9t8uQzBxejzOtCdxKML5YGM+1OSjkXPW6gNWxVlUBSC44tuhsHpP2SQsKxb/9atl
ydXh/YsFoU7pi8uoLhaXCI5YDigRY9SLdAs0DK7PiR0zEgaZGXd07EXLgf0yTwIq
NDlUY2O56MeETN6cTf1r4D6P/mTvhrvYYnsO6xzaPLZIep6CmL0c5H5jAQ/14nAo
2qwJsY1yauFs1rYDERfnZ+LTxUnr3xui5uR5khZrhMURJeI+px+aqC75K1wsAnni
DbwZxg80fJkrDmOKvKwnZPUHbyu1Qa5AWMo0ifeT+BTii6UOG6mh14SZnxeKNeh0
PEsgs2aUlVyWsi2EGuMBEXkk7iB+nVlkS8ML0QQkoZ9NRgUuyOyZkiG9T8M99LXZ
RB8qFGW39L9aeXdZtRUY6OTL0qMwGAyOh5i7rJe7vzxw8wenEtiQJwdEQRgJZHlO
DqUxF5bL0FmoGxL4gDAUVem+QPIMJf/Wp5BT+VMS9BUceiUH0QUNyrLs+PUl+vTC
UZUuSPMBgnPMfjnA9Djef3JvCVU3ysCg15mOee23RxS68RK4aBjqwfzmBhRPsQ+W
BHZCL0x+o3e6Kxl27V26J0tKe9iq+WdOA2Gzj0XqF9eKbyrTRvMtRzemKtlgxv0g
0lvW6SDNgaJlGm8tsefuFPraJBw01M6rpzYrDFN+N85IJ73/PANd2HNkYpzXpkHK
CwxDClbdsv8YNnUFwfT5mbcu0HLb55Nu3ndqp01afC74SVAkn8RtEq9iby6jKBE+
AZBWT2q7oRdGAai0N0pNDP4/Qy7nxuLknyXzeY28d0E4sXCgGS20CVbpnXZxDs3z
Q89MFFkiPHe5flbFJezqVX9SXUbG36Sq4FY8jtERUWsjtxv6Iuu+AwvUob1fEW+P
lpkRY3i99iNvFeRLqLRB5ks2uvCBQUGxydQZZJuOYWQ+RvSd0g4Q0TrmBlmMiTjM
vFGFtPCz/McVaslYBKIQgnQQSoVGqT/x4nWWrN57zF017EMoDnJRuk0u7QaRurkE
T+phLravkHeQxUDg+5MAXgWD948duEpkQneP3hVHhjDElGRh8dgVdB6s0F8ifLBm
hDjD/O3Jz+cbycHPPofraftHElv7iYgC9HVGyEp73sCj3v2skdKKRX4h6QbkAMen
0wrXtgZfmhMvJze7G8Td53JKKSJZAvihJcaT2qjrRH960cng6wKipMNlws2RYovq
yy+jF1BN6e7dP4nh4IXjwATyudSTVBv2xtT+vlz6gQu4yZXU7ItOPq0qnb34i9NJ
it5IMuavoH1Pp+2HJPpGu4rkPoKVZ3SDP2uGOcNIIalFTZ8FhD+cH1VQjB05m2/T
pQHjHyzi0gXBT/LYipz/WW9ZUaxlLwmbpAG3uzKEvZnlJ6c3qXz2xA1pZI4QoKzE
w5IOmMXKMv5OtCryqMulmw1xTOd+U2ZlgAtAd48bvKbPTXwgBjjmaDJ1wxu2Vkgv
JN+oBojLNHluK4lkuLSqaUGTCt+29IwUqMZnH+tHDTynoQGeU5yx03XCIlzEykNS
5zWhy/rehCqRbxymWNapQVAmczYoJr3sKGBXCurhrUroYJ/HfK9nT7YibJDpxavN
qG1vP4J+YwJY5GbOJLZsxGdBloBIMJmjPHMuih1cjfnTR6cauYB71233iwn/oxkv
YMk8/AuIUD5KQYuKCgmH3uPoxavUniNRd2bgI0YQxqSf2YnBVFoTgipvi5m38zll
S+puruLfrYhHzPETt/MSkoxcTBoBW1Ze1cfeAh6/wMKYspuUU+U81GdVBITGS1BW
iylkHsP5RUWYSmE+YIwEl8gatNc9XhAt+qWFH+TKidp45L0By4vsasi3e+jtzLVE
41SwGGBENEpeX0Ga+fmyrOrDB6Rm8PZhIFGwHpV9OSh2W2e+b0PTSu+piDEDlLr+
NGJwNEVsmGFrd1UO5Er/KEH7zojPapMUUnQyKHFGUSh8AKnVUUHezZKl4Y+lH9y0
fS/vvmUXrn6qz28L3KdLuP0EH7Y0oG5ZwOkEUYe/rS8VzaiieWTaheGpUtLrrmQD
dXUnxHKZ20CU/VWTwuSkibPyk4Lmh6n+EykuuRguNRWAb/VUAf6/OYlw5mflDhDI
0sDPyq6hZnYs3olgHKUtuqKIs/2fxmFsT51ZMYn9jMHnHF5pe0S3AasDDDpNIBzI
1urV/9XUc+NKJ2dF+e+xQuaF1yDG46NfzMRuMXK80Rc7VpVafJRtamLoBsd3SKeN
kb2pLuu8ruc6JZEbAUzJKpB5NmCs5QFSgHTShJTow5Eori4QwdGFfad/EgOfVLXy
+wLPML6/s/vEL71hMoufupEedJFBTZbamM4AZ9auvDbNgUWneP7u4kizkfSJOXw1
l4yU6nT3k7HUCjSSmgNJ6XCTH8qQwgoi98kmW3fwAJmg1jHx9Iqj5p4YGaBrMpot
n1TDdoZr8xHvmUA70W6WyJF7KCQ2r+1H482BQn61t5O+xkMdWSemOsRXMXRW7xzt
c/y8OtrpXG8OkjK05SEcOosQxd9QdmT4Vqy9+Q91vxNecO6NK1BjiuscWskeYkV9
V0s7lGH/38z88NXKHjDBQZqh6U1j8ZdPy9lAASF1NsbE3G+S0xQWwVtspObEcB1z
OubU+Wm+w3ssVek/zgOrhIBCuxuisHv/QxJNLbmDE15pI9JVTuf1rh1QnbnZGthM
LJ0uOfw13CA+siMoIFPVcc/52bdiEmJ7AYI0/p+nSv+N2kYcemYefMz+cbjQEwN4
Jc7LxraJ6Ge3E5nvqmnaiy6XUG+ryT6PHMYTQ/PH08xRsm9wFGISjsH/i6vVudSn
4Mh7BULXFEaJogY2G3tlrmf3Dy3PWiVVWY2Y7q2FeV37fzk5HcXcBNx/l7As9lxe
ojyQOE3cuVl1qTHOehe5Fu4d2/XXsU0bIR2C72Xdc/Nv//6Mm+/n1teVGhCJo6Tv
kTvX0+duEt2cUfFpsPvnToV76uXT5A/j3mszKng0E75hJLwyrhiYgtEqbspnGht6
IPs4iBqApZelgM5vXpIVrKQKfwE0RGj9plergj56Jh4Z7FgH5m5GvPRdNxximtP+
rYe9xFEobexyjUzsCYj8IgJvPlZ4bBd0lC5Z8IDrBbcuLrkEICLX5JR9yVnUPgfu
v8+/RYTRV2pCOKlPQzLCQ5usJyPOU0FUM6scVZHlcCZPq1dpsqsmhD+WxqvMWx5Y
aGQCUzdwL3zrt59+BeFapXOvXAWx79OHirH/oIBBVKt4aJpcsvTHZjF93jkKoQ91
FLjMhsrWF2owtNRCpsiAiIunH/LBhIsAl8CFE5wdkfQ2Yt+dr2cp16XEfJXJnedC
9fmkncCicOyloj1hPO1HrzU7rYcAUzYr+Srvp0AjEJbOHuMBQIOBRTP49cC8Xxa1
ZVtIi2FtwB+yR4FqJyV386TiSwsyd7PxID8vvrLsgFy8TonbXLaTcf4rl/N/1DMy
+UKk38zlh0PprZlfHPbHiX+BOEtcr/duz52Kg/DLMM5cTSt52+Vpp1NhcR1pCaJd
ynbNSYtr7BhE+CxQFJz16aATlB2SOcXOzQpHRaigOzFK1wd09shhYL4L99PvCECQ
+TdNclk2AwY1V2h83uKCGMG7qvw8O6HTAVlm3B0PjHcSLp8USLN7CxDUgw9U57mr
VlyvtR4iM6npMiO6KOo0PTsWXZdDkRDXMcsJ5JdkbjIBP+MPZwNUIJDURmDqUhBa
C04TYHbQrafeyuz85sXFhb2m+BJ/mB7l53T17+bG0/wcGKS6Fi0Eho/+NH4Sx37u
69bEY7jbae3HsKrfXprksnE0LxIOxJttM+KpRuO0OJl8EfmDrgLlWSg8A2jc357t
cKQ4KNv9jeujQmZRNvXp+IEUkDho+xDVAdpys44e9xv8NCltIAHpQLiGEIK5dhFd
7Q36bpGnorhDsKz4s0sikJr6FiN+Fwa1sbhECgehz5TwxOJz8suhla2QXqg+Q4g2
ulldezvRjSqtpOlMj2otHK0Uu/qELHQj4CVIZ6Twlgt0Ys0uRpl3M5yAkCjoyDo7
ce5/u1VkLTUzR+NVvjxdo5M64Ll2UyQlFaX2bTYl92NQOMzQtYSlPk8p2U8nEKNX
xdt4WkIr1xmUkssvuHYKKJh+3mDq90UlDGqd8YXBsuapsrB8nb1H3Uge26OLrSrq
KUv5umtWHm9DGMPyjEKFYmsNwj5S8jNazTqbjjaXnoJVpFyLQE8LTTB/ax8iDlsV
nusQvRZXBAnKvzUK7ZqlPD1mF25MlYQyQlNvLMBVW/ZXVg24D2HKeF6ia/xefxTX
jWdC01iNnMdRe9Wwc2BzKGlitTXzIO2+ntWQZEiH/y3V3WxDRbdStzzixvbgWmC9
esHFN3pQYYRKORjsuaLtlvYzRF7i5SpyTyI00By/WQQszbHuZVTCssRQ6OkVPmRL
mnb+mcISDrmIBw13b+Is2zOPJwK9YEBCqQXBhagcp9MorWnn/MnySHoLyOX6U/Nm
uuhgrCgcvy9Cb+7cybRrkz+tKqBgEBU95IOY9o1V1ckemhLVwkNb+ajLQuKex5Qx
JDJtJiR5ie8ayLAYcCsidNHAAMXV/4JVZU26692tr80ELL05l40gvVfOgtqmuPSq
skmkf13Ies8zUPy2pwlrw0/bdwDBcZSx0atMNH/2zlLtVVMav4wDDWOjl7OijPtE
Ko/9DHmUt6TLObU3q53gGmXeiY1mXW9XAolSqyHge5OtjCi+P3eGZQGRUbDoh5Dm
4qIr2BGwr3A+jlWK3i+zB4lDJ6JzMDNaHiUuqJqKMUi9RcbmmF7lFPX4I18pzOmX
HIm2s3vmzJYzlRchKo8l5WzApmG+GtXfZ38xckXZxH2F2LR3Sn0yXagYBYdGJXQK
ZX0bnh2iKkQGvUiwMZ/uAjsgNXYspLthZ7RxVQzxD+w3mXDOcdF6OsuopPCTNjol
dBn9EJdrxI44q4L1Nl1daR2uW/ICUbv+NfPNdUBrY9tJs1+vCQtIl0YNGO1i16gP
OKiblPcFoOf7b1MaCPj6ZHvALa89y4kt7zPmwVF345/t4Sg1dHRdTwtHMf1fMwPe
XXw3/pr2LwsyiukqPjS/ZeSuqyRylktEpY6pNdFSSbAXfDkR3m8+2h05GCeBTcw0
w/U2zsLn3lqcT8Q/q1MaTSLxeOmGyRtgxnuOeVjRkfvuBhwounZabpfLRo2k2RO0
Ehk6Jed4qXOik6aumQSSzVaElYsU9qDqhdKmlNFzqBQ0ydeMQbs/PZK8f/jg3O4X
W2PhW8ih7izgVk0NJW1Ekr7Zr94hA0MlfieFJGJ7I7TcTQXE99kYFgxGG3P80H3F
yAQr1ewMRzHLv4L8sSLE99Zd/1hg+Pj9zOe+nLKugFF7Y9Hxyv6lk1+ALoLJtxCD
kUvLircBbrXl1THWpR70ZDOFs4ajnYdLrVIPJ2KuD3m+NIuH9/hOWewWBrzvbs9L
z9Kw8+YMaJitXFkZF5mhssiUareyi9qd493pjwFN2eTuZ02KNKF2i7lxyum8VMWk
6OgcHTgO+tErIrAwLfswLQgM0VHu1VC0EB2U9znMZ/xxz3wU5QzyhOacPIuy/O5j
NucGU/ZGu17KrhuY+UrWpSRo2Kga7biQ1jq+QEnKGC8Iu3lMIWlfCmTIuFYZaMOB
wBJLkUBiOJnuJNCk0G4fN0AVwZTwUcOG4lVDXoJ8AG6eZE32RImoW9lY3b0NIibQ
bzDTf6SBtfj1wpPPrtC6pXLTJkFBYXPmrn0zqA72EvhtOBV/4ba14EDliIQEMFbp
UKhFr8hk/BnVc6PLSE9n3UOvb9Fdoem7/MTk7il5LdLOup43MvLOsZu7i8NeB+q7
iw8P3qRaz7nCSEi92ZBhsEGgkabTWbXC/863eFKQMNshhNwxH8Hu1IL1lF42k0ML
MrXwYKNG3VhuDXd7/I/EajLzbsZzdk0e1lPDWXCu/nQTmg21wJH02x3/chCul97M
IJvSRPQMyiDGjq7vqqmIjMIPfBVi0510t8zlxU65IhviM1CkGxshrC8k0ZURU2on
c7Sl1/zT/ofcmsgLAg2UrYc8ozI3VnH/LxOWZurmSZFTZns9J6uLBRCITm4vJf+0
9T57UKBxhaPhSCHw5fsOr2Ki2aR913g/H4IhKjZd/RB6olY68tVhMmNpf0DOAOFO
aiWMW3j65zm5f6D33r6OxCre7SWGvjb3Vp5i79CWQhBWt7WeGO78eIsCl+oQyJO+
RVhcuvQuco6wZpllR2A0KjAQ1AbMofhgtdG9l/Rkalsc3SBouTCzLWagkl0r2Ush
CLS7LGux/kLMqQ3TlD4GtNmkCMms3Hph4t3hm8TwzQjIEqBCEe28DoZzfNeekFBr
/gKok5hYwAZiqCoFB5734USGJXXNV6jWc+cWa0XMMb9mmerWz5Bso6i7E/NVpfjz
KrMCSrD2HcGi58qv1OBAHFS4Ok3PMrcnT5SSrXgfl/ZMdra2WAQtMiy5o/xkYpRz
XG7sqiAtZSLbiD3+1VT+nmbNrF7EsL2JMOV0U9M6xXOuqScEkQjvTOLRuhEi6DB1
htPNwQEkZh+gGmyQXfuYLRR7TpIjB7Wa/MhG2i9+MnAIHlj7JZOVRzFtwOfoecH4
4CFrIwqi3I1HASi7ZpbCJ5TDvuX++HMhMSuLDt3cuoPC3Y7LA805XK7iDj7VyRkc
yiQuD2uomVrEf/uOgRC79LVEqUfl1W4ynfRg1YFBzmY7u4MMJILOvITPpg1OSTEN
tpxrCeeZDfZqcp5kb2nx0VZ3rsjQHXPdJRTt6Qkm95c4t+OS5cflbgQfFv6aZpxq
XjNeUB0qXwm9Wa49sORv/HAhvf+g/nPUhB0eCosw0SVf7vaDwv36TmQhgaCr5/GO
7wpPw0V/iFnpMaVdYOC2i3pRX/z7MZ8SRPUdghjQzNpNAW2wzZubt/vIGydE+4UG
BJ5+L/UHDHgj1lwYrbhyrDnHQgLRlqXInvA8Bc/x8yb5PNXBq82HwzrR7SYBFwJv
3uu03pP5BNV5ngPo0Fqm3bgsrh0CuU3vY5RyWfasRzRyUDeXzkcxH8GUpGke8k2c
svvdYZuKKRLKZKuG5YfijUn3xIU6lHeJitAltkjwvxBaIz3sF2EAlyQ8A66O2YTP
30MZsG4M6eKiqq9D0RWKdatgKzrzLxQO0jTSoFdBPc1xV5Tw0TveOehwrrmtEO1S
Py5f7Z3S/PBgBLhfjU4MiqpK1bK62rPLClmEzGfc2D/lzTJwqyRKfayXmFPyoFO5
ba0e+efCqUHzpkcsCmS+oAxYPazqychEHaEOgDcqoeKFBexRSz40YIDDpJp6yZd9
jERVJBotk9COybUyDE/+jq9Humiv4YO5mmLtvyMnAhVbKxZo+26L348iMMGFQ3Cp
grfmfMkO+7CbFYsu1Ou5OAwyxhJyuRdizlN+dOINnX26xC+bPIwir7ck6fH9HCCB
ajVjt8xv4u145eFhXPwQY7sr3gNR465K6H/9tsJrr/U1pIvKbWDsAM0zWT6GJYqO
ETS4jd1Bl5RAH1Jw9m61WpZ0Ic+6odgFExVJtgEbYZLHoWmXY9yYtIBLpn56SWXo
vZbnURt257msEJxnkxAVoCYLZAxK1nckCgenEi+Rh2OYVUBiSjB6WDGaA04Ovjwu
mPt2FvEMkmiHDwpI3JYfWmnID+0hmgcYX7JDE82AkRY9XHB9+te/XfIw+kFBY8VC
9FtqOYo8ECvtDVZVQh03g8CgHsjWZCpufRNlc/Pyt8xnMH3wOeQqxVMN0tUTD9L+
2hP12+JJbwYnQU/2nTOxdLUd9aa10gfri04oL5nTQG8xO2S5/Q9baA7S+ZgP6QHZ
/QlpVDWnTVGQevJd30NXaKp5iD5co1/gfaUOXMW+ETFNyrBXvL5C4Rqc/V0IlgBs
qOrOx5VyPtHF6b10nMgo+Nwv2cHgPhyEUnyv+Nb+PCIkc0QtpH1F8+bXezNb9VWk
fCEoEGxgGS3CGL4QuFXdXIDEYFRTnYdyVFxnnMjIdDbwzTU72oKcgiZZ37L8FoUN
u3v7e6ybB7lmGAGldbtRee8U14O5dQRNWifHQLoraW8kjNjMYZpjiJgAb3twhOol
1ywqo+j1jSg0ecHBF9Thu0Xu7nTevYUeqbz2EhGaxT9jRSfwfqPQZ1vqp0+G0dwP
1WrIhlPnGidxCVHa250BQKyZ8JOSZ/+4mbs8H2MSSUYoSQpkrhIzI346W0U73R3v
d1yPk3YDXoUXCzz6gnt91vo1chbQXyJc81dAUrGvubdNmom7Ut/f/TuEPowuAGIP
ChjUG4MPYV6MjMVwbP+FhPi0m4VsUyMbh5nYh7CUB7c+TLA9n/MClqfy4gKceP2m
MuO6OIDp4oO+3p5n0xUyXod/9uA/1s0sNR4EqVYRpgEgWeXkaY5VEkk38n1bLoOb
i/v/fA60RazSuf2ifISnjmYlj2OFE6JR7PR5iANLStmKdV+I0OMC7SiBvN1pMGb5
Mn4nHh7UG3y2kM5rAraqfNZ73BAUG1r/FXkeY+UFS+AkIykSR5IZaTbs02Qc0z9T
rCTKpgdL1HdcWHK8DxyJiNlSyqbVnWKDjYVdr67FPPyLmNXTwLNBeCKv9/O9zDJ5
NEH4LrkFcHLv2pDIv8UCew1RezNSmeG0cNwGx1hrrGumcbCU4sZRqwxHuzOPKWs9
BMHtDEs9To4mJiL3PgZdpMMpIVCj//OYIPZqsdkwa0G4TSRVvK3l8tTw02/l9xG0
9kY17yL+pBowE36PAbWv+Y1Vl6S0MXFCmSV19+Mhjs/zj5BJNcn3XHkG/NOsqStN
d1M3wC5PajdQLLIuu4rOo5XJzg4iMo8F6GqyqXbxqfCBf1ChHaaSQEvBbMR2IU8m
dFn9AgKwe3JKOMlHHXu4DO9Y4DhV+YGobobgxORvHXVIDqe0+iJ4wrHgTnWjMHMT
QbQAhkV7fq4rKI5aEYnQtTh4yTqP5NYaCenpCe7cqvqvDEsn6AoPmY+geIMaA6P+
EsWCtlwrNj/EQwJDeLNbSrnO1EuEz7qanLdJnP9eCQbeYIcL+o7ctBERU46z7u+J
7nbBYkCNkIZpKshioT4N7rX4vUqKBcQKfDxZOCGMg507aSgs4sZZOpcNyzXrA/uv
dFwgGz/dVyydIWxMg+N3XTdslUaeZ5kOyhHhRPlDy28oTo1vP+sRvccHh1yosIUz
UXUqagWMghtxX/heW5F8NZJqkx6p6rM7af+neROEpx05FA2VdaaaHBLAK75UflVI
vwrb7Os48EMHcI9kWfNhG8Jy4Ro0NvA6aqTLZRmeksKPrmqj8DDiLSXCbn/dHI7F
70DlTIX5kMSAMZUg1IEmFKaV0/N0ROB/HdBPrgoip3CtAM97hUEE+STnJPP9hdUe
Z/rl4OyY/Ia4RyXSVH89RatqRKfbk938/otxLuhsz9jlUag1oshkwfc0+WsJPpsm
oL/mLv1tyn7Xt1lho3QttplWOFTkbtQLSmfEzOt/Whr1bYD98iAFXaBA+Iyw/FRr
1xIZwcDhPM3GLFUgjxJE1S6im9Fe/19ya//H31h6wd5iPmrf3cRYlpuy8sUgV7QG
XNkWPz8cNcs1GQ9KT5KBUqbS4jsh7ddvrWFfZyKBbz9bUYdFv916nsEs95hhlGTh
7iLiTYSMWMBFcLGmsoSuZmvVmGDSnKG/Po1dwAKlmnwNG09uye7odDvO5bhiVNRg
pbchzMC3YQpDvjwrYLzThVD9mwnz6CvSYewsLYbyEqZr4/iXyiG42+FVyJWFoU7K
YXkFejLohyJ2vNbUR44jEPFlecK/3FyxtasGFNoECAGDC4Jk2UDRxCHu5AA23veX
uYOqMog9yILOgCPnP1WSR/5qjYLDahzNF4gjo+YajVCYBUFt/ek8dMhmmmHSVPFh
M0cwWE8zdzjyNrSBQaeWghTFTV2wh/obmHIbk/DlAhBa6ttZwih/JVs6ZAHjfet/
COpf9jyGXw1lFscuJ5fQs4qxXMmFVVSiqZAXcH/fHo4euIJUJvEuh/I/6w8PgBu5
FWI6Sf5eHRE+uYRjPbUa8taYYM/tEXOkQFkSIlJ/21cx6Ib1ON+ZCnEOokB+ZUfZ
+0vZo/e7lTu6R6x57sBSmqYQ3mFRtbrwuGaLiBUA77IQI0OK9frR9LiTM7/tY/SC
y3aN/isgv+e83dxgxIlPne9kbJn1e4iBoFbdS0CEwtWt8daomtexHcm1qppui66t
jY6gd9cWrm1QGBZvkAFLJtoL2Gn8an5sPpkpR0sd5AY9G31dkkZdO53MpvlF+V2l
uVml8VoxnzBHXVsjAKmyIAyXOdaige89z+loj5CyOFbzNOH6G6pbxME/spfEv8OW
bjBF7mCH/PoUhQ9lguP8oqY7hQYqBPDwUyC2opzzaF4bwlDUQlsnburkOwsGlPxD
UwVob8GnnOo9l9rV1x2BjCt1QfJJQ4+2f0fU8i6lsnZyMGobFeodV2Xdv3+jcMV7
a62/LGs+HHWm4vGiVJX/xGB+4RHsLYsw4cejNsga3WnFTK4tc6vjh/rhRYVYEcta
44Fx4U+B54E0JzGvE0/G4Zu4DpZCV2gWIUlKfngWocacBtTH3gK9TcDhj6vV1IWT
5S+k3KCtuOrzi89uGSQBk0MKGLrRM7N6rz6mm0hbcQUUkY+8ZxljpaoJMVi9JMDz
dy5BIj1LzUDgVDR+N77N18NAKcNtAKjtfmjEuLGxnwvPnOY1vb2IoH1PaFHD+VUr
eEoIo+SFQ/hnlMWQ+n0UaivdBJTf/TKZcWCvHbsm4uB5mS2cb8Kn3jBMFHj+DK9l
gtVVM5a22rSCWvWb2QOOhVYltNanoXp71LJDLciY9RbjOn7dxWU7LIXtjbOgz4m0
0n1ZpTH0yomU5fiBx/yJvM79XFTzCl3WNTuMyNzgSn5DadIPvtlt2p0YsMlzOGzd
VMuv0Cm4WJyT2b33qtv2HR8T/rTLzKVYhnBjVlWQJs7NBuKEtE43yppNrV9NMApj
ybossmPGBhOTIjhceS/8WqTQmrL+QeGCOOroLZdB83n0g51ZEciJ9gunNBpus0nE
PxcUsCFsHh7FUg56vSQEAZQKdQm6F7qUJz7Vs9eLBNWYHKdcZ0kZhghmKxeUzAtc
2PPiJrZducZJDiP3cVNvx33CF5fpAMLjvKokjtjxNTjkkFE0RWOfR+4SQVoIr0AS
cgwwoLTvZnIb1B3a1V1C5BokGx7NU3wPRCtQMC9iXsKdEGartYqrHu5MrUcTllXf
c4HiQOJs+lIzu/WIuMdPVtqPiN8UYZVobwSByUJxJ3yXsvhl9AdyRVID/Gseji/J
0KYIsHrg96o6rqvT+bwCgsVlz4wLureyisWMfQGYBKyDmz/oZuMj0I7hO6EoiQU6
KjqWFI28vDYxcHo/XH1zUp7M/HJaPYucwY1Fy6GBoEqmA95BOMFDmEQcqph+/0eF
FhUvEIy9XsBE5rKYGFYN1KzzyrsA090k7RCxwC5+bcGaqS4b84KrK0Bhx+/x/ciq
bSxcEtrWVmsLoIVAgimh52pH7VQ1b+ZVAoTW8mv5OlaHDoDnC79TUSAzR0J8iC2r
dTvv6mBdqCrigbFGmCiNG0eJ6SEUNAJwrnOvh2+oUgWkMFDfu/KRn6m6eGmFOSpz
+1opKFvxzLES/WiMKC1sK0GDrWnSZtD/Ujmp53pIBEklfbF128vkf5AKIE1pC1n4
xIDxtA8vUcWEzGFCZ3IYWWYXmjS8Evu7VfF9d2EJ+RHPhcdgMouBS57rvKhtPflC
9vKMK4aNx4iWTnGaeCqPIwjTYciDnmEy/Z07OFg8Xj2LUfiYX+dDVmVBKq9q8RoQ
yPE3QG/9RfC3QV2eM2jx0VDu6EQ7erNfSXl2ggbVf1Cfaxxxma+2M0G6clzjh21M
S3VlTTJCOo4xCiuhEMsrEno+dJ0Wyfk8O2uwLKs5jn24yMfabvScekjbv0nX22EL
nz3qvphLnQU3WUERv35Tszgv5w3fswnk8tcbgDbMAg7xy6qQEx7k2vTUvDQWfC9I
s0BUBLv7D62d0FoHzjeeCKriLR4UCm8tZlk74p3irIl6mssF90YmoltUIrEZWJ/p
qd4BvkEYq5umEjbYNJEffy502Vk9IljuSUN5THG00fMGqGzhxmv3qlxM9JTS8fWT
LGhvPj8mJAQCKDByvYowJzA3ZoXb81fvdddYI7FJm55OtLNIv7miOfHbtkLVXktZ
IXpYqlnEp/nfAJyUh3FNkMDiv8kSkQekvrXUJpZk/WccbUKcWLkAMqlsYkBfN+7p
UEQEp+/VCb9coyf1YpsKRoDpSQ4QpCFWpBp9dctRzjW5fzjHBNgFeXGhlfaiXpKI
hGTmDuG0PBg+xSa6A9TieXjEkHaavj8C83rzF42sD43/lMBinrvGEQP4NbH/EGvO
q1kIWmNcOx29fIHDxRXzOxXFlQL4FUA9ENpv35AKnJQlqhnLG1Mr/PX/ULk7Qxb5
Nsdrmy6hTnLQNjFRE5wc3QNfcNFkxnGwCD2l3DGuWfnIKU/f9TQiWf5DWH52Z3KH
CDfoEM7tViIxRZTgDsUaCnsfsEcHdqa9f/M/h3yp43NQFK2wupgtJUZU9I7UmlGP
IJMbhrlZnBjiCQ3beQEHwIuDCeqROwcsRCgVWgwoDfgZB1AGWHKAeqZ5MfbtvyP9
NcOPz7W4R0+NX16EhZy9MLyI3uEQkGXtnYUfq1Xoiw2xdOl4pLwu+RrXY01ZQ4ml
udVhS/mT+F1PCYOvPmm3YVT4pPh9R1/0/BgrwCjrgI1Gc0yUWJJ2qp2YmbKfaZhm
cXco654DDUFXTA+LZvXCSk2825Cza7E1l6j5yIoNJBRgng7mC2hXGQpBk3bK5BtQ
+PTToAG61lmK14An1d4BnTPwkl7SaECU7FyKMOm0BZY1B3Y6SklnPb3hwPJ7WXwd
hv3t3EiMGNthys3lZQe/lDQHJjxiI7WpoBnsFfxBfFRCkK6E90mS9ua9zREsAVRQ
GlRqdJoXiJSXAmYfHXBweZ7jnidbgTUY9evttnQmIaVI35tbVRfCsHJJFHPL2sjb
OgluGzHG0l4i2ePidPw9qz2HMTs31r9QC8GNypXtx9drvRbWomWWXnn4K6wQHO80
F2Gh27y3lB8ad765hZBDnokzYatMKwZSJ7l4CTwuSZTi4HT/useQ+ITf/hoGHXzl
U/ol3oCrkTUvXHFVeirwTjPIAM/LD55KD6g4KL7nlHg+32mjabNFCFw0pNTgHJEb
vm06JPQb+OXhbZw8h1xrI4rLd9StsN44IyXbu7gxaoNcKfXI2pGhSQEr2FrFAvQB
nyrM9mC0MVtjt0Qh6lXOl7UDbGsgknV7LlQ68qqrb49/WHvxIbpwM/k/4jatKt2U
2HrkXVYiUlCMLSoRYu1wmkoPWlxMrK4RFKDH2PD75vsrujsaN4wvymcpfsweybnK
+SxZ4KvvuJ4Zu4nxc75fDVEmxzQ631EbmOu0nG65zg0cNYIa8K5WpRn4ys8zFi5t
okB1fW5kMgOfHXJpdOZJALdCLNB8pgeMoQp02yh5ONa+wpQfiyTNsUqNKWXYxhz0
E0pYJJXGF1IvbkbQkor2/5NbLcvlVkbNTXhStfvBWE7qB/jjJZik1PrE/+zZz6BD
fxA0gabIKDdoAL2ypC1J4kz8tTywS8Vs6FPYvr0TYHVvyxSFtVSxgbLysoWPGGjH
8DrYuGW41pG2XlwQZjj7C1Oe1873DoQbPgGafAWVeNyNcvnenOAIWinhx0pv3FYV
vn0HTCGhHnEOTwOVhnpm0dRlPN3ktu/qn/xxWFc1CGX6hV7enwGnrCjim0nfGavQ
PywKatAo/bBU0+ldwCdLrdad72mc4jcP1VBd7ji2Y3qP/A+50CXU+9Oz6CwVjhk4
jqKaP9IxMRr4v9KcCU3sLOcyNZhEcE2UqQArQMasNJnFZv0b/p8lp2JC5mdwxlcy
/lyt9OuMAZ06i44hYRaAJ2ebwRX/rpKgux18x6OGsUVWqq+99Re61NgzXaN5T2jr
kHui0yybaJAlAk4S3Fgz7gKxUP5jOTqhLkLnhNpch/qVyr2SA+913v+P3Fdtz4Lk
Aw85VNGblvGEyO5ksYiRrr4K0An77cMt+JmZDrccgH3TMYROaRte8un6q8nlAcmw
Vv6+F0hLHVcx59gHxRM+pnnm1FK1FiK5vgx6jjLxCn8NIh6lmXSxUgLgNxg64CFh
8T287dLgdfgnrG/pCdeEsUFE4YYodfzbxL+Yvo/x7UzXSPyhuaMCpSb0WWoNGkDw
lHsMSl2ovsNESgvxAZP3CRd6KNoS2EEfb+778uswkSnjrARYraAkZkXjYSIGkqds
VN8KVnOZQr60cRtzuNuQ0/AIAvGhHDa04tzTeNWk+N6I9RgIshBQWwKbntvMy7m1
8HWclTKUYekF5BW4JDCjruXXSZmwuiZfIv8OLCoEMVVrfHk1yeUS3n4T3J5Jmes6
2Tfq6whkg/3IyeP4L8chKnBHcrbjZ57xAG9PoolPor97uSRDP4ITykJNTKAoPf2t
184S2kF/GydIfyiISDJ3io5SeaDBmGj2dBw2pzT1NTQDTWtnlgZocQ6IDpfruxUb
h1BDToBpWJX4UJbXLZiqedcyXI5JXqq+2dP4I7deXMJM1WlD5sDlQLHuYNgIFeHm
iMLBVHh7OROZvyWdG2V4jqEHbhF5ZpZAc06CTwCyT5yKRi9bjedsZ9dd2HFgzUfE
zblHDammrXXQBXm5F0CbjjNm6hsQ6FqNDHOOeSUFWkveBqqAKaUyn9oeFOlFORUX
x/lSYsxCVungo3/UiFay7B3R7vE00gxr6vNcNp+QJhWzcJbJ5UuiH1Z9jb6Yjd9S
BaMCLndUpKqwLQwv3Pp+93Zsb4D0gK+XdGRq50zEbbQlKee3vbaN0ORZXk3xELZm
o6L5LnBxHSVC9vg5fBRJx+0Xc3O6M2zO8qxsBVKwQw21KOqJk6oWl7F5Q2UrUkhy
64UMcAmgnAr45GPABbTjtivxZbxKv7QezXXXCa8pE6tmQgS4cvG7sQL13uCUWLBy
jZ2p8L3aMkIblCz+WEgadzvZu0WdgyuSEOJwGK6uKxKP1Qy+zPY8x2pKOPvuhe+w
jpNfwHI5Xj781ClowQTimWrpL3KkZ6wxuw+HA9KxxRG795rLnfwKlP42w+BH4Iel
Oq92g2Y0KhrKWI4Krdyhn2kIFeMshAT7BoBklG1CD+9qtY31q1AydBcUUQnohM/c
pZpLf/SquMLZi7P+0H+0jILSyDDNWEE4GpnkNIq8NjMC921QLCI74WLpxLldZS5F
xlHKwtuHXFwdi5L6/zN4gKRiuPtYRDUWLfST3y1/8t3M9Z2TAKVJWsi8Ox9G6I9Z
Np/gfxIwenXqEWhID3mNLLO3f7FR0aizAceK3FBVkvrAlqNWB/QWqE2GX6r/1jMk
+3iV9TbXpdawW4p5c6vbEV8edQd50y2dfbHwJkGaFwW7hNBtXJQKQbA3OrIgJ4Mw
I3DMLuzfeUtQZaYeKNHGVa/i/u0VetjhEuTu+6YRSMZEA/0i0o6XTGNDzj5u4r43
mJbIr4ZzIv+x4XqFvkAmmEVuqDHk6hNA72ygag6cxg48tq3VRRvUmOLHihHrXGci
fLY2u27Y1Hxu0OhFx4txCFpl7lqhOA7CanXhOK4UBOQadkU8Dxq+OmZ3UvbWgf/E
mRwN/tWU2BtQ+NSrVIu4/fZhFxCedV5kt/ZgCHzvEf+JKRMA/wJviBKCpFS0v/Rb
axuPYZlCHLD+WTdzA5VgStqtCZtJjG2oSgENf2GVnE3FZeI64zwYsfQ9pjqhPj53
kPdt15+dtE6cZVh0wqwMaRDw1Y1wvt8r0brpnS78iq2aPdPNU0+MBSF3XEHiI1qm
RdLEBNQjQVak55+CtMr6h0DnHQ5eSI4YasdEvJkk2q5EjzanLbfFz6VdiJGBDuwl
v40Hi9lStQQrCB+zjNm6h8rt1U/SC5s385i8tbzjfzew3e35HDO4rmuC3FNvhTno
kzkFkmAuhhhNx+GDr7aQtF/+PLQO6jAh7BB35/pF62A3PTUzNeLYcxH5HUOCSdMz
3n8z+9dWrShEvM7Rb7ePTwSaAMlpQtDaHckmuXzhHfg+2J3+h9PBzYzbQ6l/z8u7
PYOXOb01R74fXe6CmFZ3iZhC5qvYmFW9RolRWvcqOcE7i0LkS5ggqMcRZKXcN2N5
lvtCMh2kMiC2lo81IJCNTUpCnCGGX1X+FiqRT+Zdt8yJ4e0wt2+7HFN/hl8Mgtdq
lNuNMfNSgQbf4XKI3PsNliQXm6WN7cUzDyQYeTBG7xOQLVcQWQ2Y+qZdOilfxdbK
M/cLCLs6/SYZf/Q4/az5mX96pNxwKBByD/WsMPszqa7rjo3PQCIyLy7g9hgxC84+
5UXhFGNkNKDNKLKBxZ5NnqAXhb3fbTluvNlBJuWyeNMh8E+b3DT7rnNlI4tqn52m
Y0se1hDlFCkGcj7GNccMqdT11OlsFYsrPlEC/LH8RSAFlKQJKqm9BfO7gu4ggIJp
7em873sZnbMxTil+xbIItwTkc3JYHA8N573PT5BS23hbu+FMugDt66GbKcu8efOU
YWy8h9FIc4GmyiOv2Lb7UrnNuWIzr88LNalAeUliNLUsorv3U4NbuzGSIM4KQCaU
sBS4+5HCzCDouyMC/1KpImJaBs6srsiUGats9xniL3pYuiSDPxwc5Jg25OWnI8nh
0dT5zNJ4dVzanskTwNwdlvoblsrYp+KP2JwBRrJd1q3OuaOZjJTJFZ1vsfXFMhj6
EsQN8nbcIFZ5NVjl8vfPhpZ+xLyOdwHCxTxqLktvm52yohLzDpqKeyJtrj6gVk41
xLB0NdefRv1ro84NgWqdj9pmQWAXbarVRaIbroxeqsTQPwY7d9f3ih6mpBZgs4sy
v3bUw0Mn0/cjKTmK8QfD3R50+fc7w8/eXRURoTFPvtaTUy7Z0KKGRL2SiqghspLC
Y3tP8FBEQlmSAGLyF57Xh4/sYrVBBL/9Lup4SnExd00n8dkZqXOhhXbQvV/JVWBZ
eBO+4Lidiv9I/jCmxCTnhTzSo5hQhjhicWl4TcfJ9pnH88WFvLVBjKSA7Ti4B/pW
HKOe6b0W/K/H35bH+cc2AegoFR7qc5C8FfmbCYTTDzgqMUQC5miRiDzvjMJGFphd
jnGYrfRnU6xP5HLrQEKoG0b+suzNRBsJTHmsPkYo/V37b4QueiSf2BZeqxaq/Yg7
04Ig2zj//6CQCi5/yrIl3gdr2cTpTjbK4LhMArT7yJrkus28LdYKLCEyg0abxgBd
jy2tBBSI7bTNr1yUFiBT9KRg2DEyw682L+NYe8Sc4JlqrKSjAqo/3XBxxdZ6lKBQ
SAFIjklYnuGr4BLKpb9C3lFHxiJ8us2Q/p4Zgt6TRSR5DvcLRmwwbQqXORDvTrdd
Ehez8lGphxqTs8j2UV68nXBPCC+4vam0eohl3DnnKlYmtsI9MvYaQVvVxtGTSuK6
oKvxhsp5zzhzyI8Hz/IsyhjgDt9MkdiArRSzwGUlsDU6pAzfttpT4gBFWOA80Bym
HWCTRa7t9mLYFA2RGt3a2MeS/PuMxgnuasVzzCgIHFj0PHCts/K8a1chu58mnhBB
oPEGv4Zxe6ZE/uF876W4dxCyr0C9YZ8SKA3R8QVa+vFevLnkyxLQiosdxhU6T9Ww
fHjDnpvQa301K2aIGv50H5el9SEa3U0tzn1qK+Qbc3RDisFf11sdfJHD8zgZrHST
CPHjGv+MjTaFgbjW8+DEkoPppVPWl9FYH8jFCTonWeC3eFF89dwmGhPBy0LWAHn3
bDQ+k2/RfxlCCO6A0IU3mEtNyFKOHNamjuat+hBp4ymnc26x37bcUUCjbg0Fi3o0
bJ8tog9x+DO5uiAC08A2kcMeJd1lrWcOmyYie7thRCbRfY5uf+Hgu6+CKlnNbqvG
HbOZzdZQOw1r1G4OyMaRfkO4aLOsuNswEqEvihTRA59D07Elh/qQWwVUYN9utNIH
vNdtN7q1fOHYHxM5rzSziB4oSopJZ5qluFLQ9IhXdtPYis5ZclBvodUa0WTr8v4M
Mr9jX0qiEKCRtjWUkTMgis5W1aRvS4mxOQJVZgzfHi5hHoNz0jpbuBwY/QhVw/Js
kPdGJfjGaUNbCTDaaX1Um5aGEHLmcs4YbkcRBqJlqC1IaSTR8uDq7XAr9rrSfpHa
Q80sNlc8nxPGe8nxDq4g+DyJiIJWrmhETjIR9VBL/owz38+3yNMhRuMnHhzh+bSY
J3PvZ0hyaS6sFplBM5nP6XJkQ730jorT5/x+ZsAnNSRMJXOoei5eSDzmCjoyoC3H
VgLwIpo08v62qeweLaBWu/c5M0Tt3f5V0BM1iIe/gO1R1nxVAd9vha1njIRkZo0/
KvMK5CxorFQiWDC+as5Fnv5oA5jqQ9S0GJu/cSXx5uYeD3Z0rhzH06hWL3ecGKLF
JigG3UxcM298tTdAQmjR9CnZ6IngQ7fZDwHYdUSosM8TVy03i+wRnK6yLPeNlwpv
A4TojLmoM5VpNLxZzxACAcJ5w9t0z6NEDJdla/A2dw7Xbd08YY1myf9gpTGvDLHK
AeFsg0myp6gAOzDbVMjIZvYFQUTMNMwLsRMuDYgLBTY3nMQfwzs9Ec+8A4sF3Q30
3yspiPLAcGBmi8khWUTKs2BzEQbdgkESpbGYAdRr0M1vBSecC5kCd7Cr5WSsVsrZ
h3xL94v1b3yzDBC7TbRPhb2+P+qO1YmjmYm65xgLWe+NQUnW2Q6c0rYGR2WA6fkr
c61fjVCApn0EMEpTD6ZmElystVZZJYwWpVXSdXM6+WKM0mN96gyCPBBJVeawjc8x
9bvEP+p3jgEJN+y2gvfEhpc8SFRvtll0YaMIQouY2gCUfjF2og3WEXfzC0kalej4
jkPiE82MzkH5Vln0hB0PyA5ZTuvqfXpQJyh4QkbaYItca2tuiSa6Z4nOAQpHGYry
VIv1qLCWw18R8iMkpoQxrn9SEvKOoPn4Gs78RNKrX9kgGZxRD3cbAdETDjP9t2ok
hhar8qbm5z9l5HST0LmEX6buM0dtyYExQAXC0cV1ZucUuULJ8k4OihXyf+UdrkLe
vUEAEwNe57fq4MCPrGPzyXZba86KbBOKWkkdVbpbTfrg508UkPc6i/R1gGLmlonZ
RQaa5sfmxY8RTPXEsOIb3IR0FJsUkr6+tBhUod+J1sGK8U+BwL0DU25P+Tb4DY5F
x/q+eA55i6MkLPmxnG1uXjHzH1plQOm7j8FOfB9yJ9AyF54P6bQ5zWPMYdCCOa1H
/ZxgcCN8mqGbvgfnH/xyazOkClPaxzGIJ70FaIv1unYxk1vYv55SJRjunIxPQUXq
wfoT0O9Dw46kvxmUWmb4pVEL6fvT8InKFI0XJMHPuV5PTPz65QkVp4jmbBQUX0wu
NNIhLoPDgueqNCaRpojaUhy6BVvhY6OskQgAxUKyLK6xLCJQy/WvTKkyhTBDeCyr
phHifNdqIHqAutt6f39P3jUNKj9yx0wzbhFVW1zMvcUVa3J54nlarRgeJWYQb5cW
Yn9NuBt/zFIMTcnIwMvdwzud8a2K0XtWo+R+eygIBaXL24+eFTWqM7axoUdBWq+W
+XRsb9/T9YkJ0i5RhnfLf958k64HRXo1I8t/A5if7S7dBi2fvOkA2cIJjOntwxjL
imT8lu/JD+4MrJSs1+JjTXA34YPEQ41vtXil5B3hO8fR6Sje6D9ZQMWXTX/yItKW
ePe/zn7MwqkE5HObdpNe8/y46DpxA32KU3RCm/yG/fAnndOSvWvzuLcH5kcnYYLj
ipV7IS14Y9gjbA+nIzQW1wgVFABnh9sAUuV9eF19VaYnJ4+CUqmDXPmek+cBxfo4
qpk19/RJ62mTvRt1Ld15LRdKHzZO8kKNC22FOeMGKwovVprXYKI9OnSv84hqGahk
ldmNoXMRc1AgXcOP5QYicIatUoUwYa3qVSrd5RF/2c7uQJlcRP2s0JE++kNX9pmW
T6gc2yy08TdaIlO1B5k+jVTZJwNdbpAFoM/pj4GDW0iAfcgQrSf7ZRkH1Y2ed+4r
w2PgIMFSHG56Mh7uDUEQVeXz/yelbpHEPdkPRSDKbU7TJOsnw9Wmc/nTHbk8WJyk
0H8KstpEu1NkyJj+0w52yG2E7VvMQuQ7N6m9OCnndHUX82cP7iUwUCQRrHcRhgze
/E22GbQZn6m+38vK/8S9/F5OJ92nBJtdAsHXJ5ylYxeFEQnCTW+/71sY+N6tl97w
4OlS5wnoAS3K2Aumg9OYnAy07s5dfrUy7KktvsubszHRfxzHkpb6eGYFoMgxen09
lp30TX4pez2XVRIR/fStEnb77WqJrfFexWmS5JYDK/RofTL3mKvbO/5/CtJko4JO
FMv2h+MO8Lk1Opfeen/bur6AtGQNO0LQZb8J6RLVqDvJyr9wORsq5Cnzq/Hsguh7
+d16FFYlg/99snddQiStlK556DlHomoHqqCoLotQ2XMzDOmOD6B89NYDufQre8V+
47wKHOsEmExTarlCNNwk7/+gxPkXaDMb89sEycam/+RHBRTyDBwKGy5tvQ8cKMr6
k+poTOcQ8fXPx3pcLYtPd36Nxigy9n/TIorhmDtQWL/ulX9tkcdTX0PfzL/yUVNx
tyB+/yy07jeaVNrmuGQnv4oz4upOzaBmKhwk0yHQaDihA4aJXCoWwBxF3LtdjwJZ
SNTKn/05VKDzT2hMWe9TQ/aROVsN6kx6YBepVc1/P9mVK/5nrST8oVxNqPjG3b13
b+wO+RudO7c3JXrmpgDdnW127RyZFFZ+PseZ6jff1gp8R6bxaIhkI5Ehvsb4SCAB
qsQov1jTkWFpoIPvvthzLz8cxWxInAuH3dBwzHoPY6+sdB4y4OP/EKMqJzrCNwgK
FLg7AVtsFILdLHplu/SBRgPmqQ+uGKdUpQ6oUsmuJ53uf8spEeHD3JtMT+KKWWVC
YzaKRe6zRUxuOCJfRem9aGjinGMyIwHRHzD7n+bgPxwpT+Ends3JHjEO4XNzrrIv
hWtjLUOEu4gDWNC+DO9WB91bhsmlJZLjyNSC5HQ5XzUrZ4wNEs4rs0vCOCicUyNx
rbQbmUEl9ORB8qBxblo2Q0mGUejlODEK5hHI8FsaN1sPXSzGVPKMLZn8T/QgQGy1
Uv3CofZAF9vrGU7C+j7cZR9t48TM01BrmO3IsJI3d22qPO/BxycrKyFo5QMBo/i7
dYBtS9yAMxkQcGg2UeOJBZGfvFxtvqztMk+7S75RyU4iSJOWmAkPUK7VTpj/XxCU
MlaEvH9gl48m9ssTRDyrDTZFDcL6/J9GzSzYxS5JOzg1YIxVyQXZRWkhbl71Yn1E
dAGmrYGY6U+hmPgJbFN/g238Y/ONS2rNQyPrZ8Qo4YvsiWY5IBhFg4nxt7SMzG68
bea32bMX1YxH0N7W6REQ2GP62AqkpNdZry0YiZXw9RnZKRqbmBJkUcBResqQhNT3
kp6qnTCloHvrfNEIkZ5qXaBac3UM1fUsuIQnWUVE/VnSAURIB7fy87t5HoIrGttV
/p+BiNlgPPFyFu61vBRXWDAdvvd0uyoIREl1rBfqcbNWFndGLUQ3RT2C5EAYMb9G
hWwJznA4lnpbXL2Ca9nTL+L2PWMZmy1j6P59K7DZLcnOWJbXqxtuylyVvTFlx0tM
5OzHVxRwxTlldonG3WshBogEoxZkvkjNlhVv3FvcOhqLwnT4w9uFtupvG2j+51lZ
wUFcrEU7/T8DD1xXZnQvHOTPh104+/dqbK/3c4ko2oRDOQ3m0UPavlnaG+vGEDdO
ZGP5SfGVDaudu4ZzAhMLAETcUKTveD+D6kb4wnyxXARmqLNCbIcr0pM8WGVhYdcZ
DKYPTPyzkOF4xI++unzG6czxU0IbjdlWRO7E5lU5Dr840F7ZSFgtaz7XvlmBzAAX
4dfx1gLAQKulXBWN3hXcBRTGwqR4/yj1bmDFnMBDUu2qQiP6ODLQGDmjO445JR5P
G5xnxJpmZYJMUSo20lEkMd1Az5PUpAD168GaDwqRnnH0hZHAVSrOJPQGe5RdBhEZ
MStIC0O7MkzqjP41gC1NgRD5sjTu3igIlQ0pWgLbX9cLUueEBhFU/3X2FRoKrDue
aU/ViDk2/5+FWS/0sVx0W8bZFSywUL2g6xdT/fIoVrW/njMkIZ3TMWa34SjUoA5P
6qfMlXvqzjh+Cc91Ch7A2qPNVMZhEM8uhAQ4g+qInNJZWl87kuOgd+1BQLAhbV5j
nNClxNpj/Qj+gnN3jDZhdfpW9UljMWRaLaLDT2GttaQudGIzC1DjqqYLrwZUIK6A
Wq+SI7CLZRglnZoalCIOd2HAPUUZsyYpv8Lt3nJkafu5TVTDCcxyjuwBM1XpmNII
55S5sI65I/YJI9fqzN9BZHMboaHnFSmY+91TFuQU3xGTf89DnU4bkVy85qAOSaL5
iOBmBvTJQP7FqHPzva0/AAP0tDQfzyQnuYoItf2KgZU2oJsRGYiNTxXOhx5Yr7Sj
YQn7wtEsQVObLIDPHhTdlILeON9zrwTi3owfuod4k7rfhqIBd1Ci5o9oYCbifgW2
6sW5ttEfFZfFy5E5Ig6WKoI5rSnoLitaCm4qhJn3rDnaYQMcf6azzMQSVwOhbsHD
hdi3bsE3O9BAv3Rh2xXBRYzAZXpA1VVdFsZkHuYJgKVcWgewiEmx7VWSYGnx9LMk
Q4IMiKfJGgzyiVsgv3kneqCp4aDE92IFCLG7rznPqv0jjXBamaVlm2994WGMz4kx
GZhhP6OSTUuyCBTVlDqmuADp0SGqIPDqnlU7EfdxwwMOZq4ilLRF0+KshU15ssV9
tGLDnZ0tqYx8hmjmTelRG+HuGzOR4sRwK1eVzBYanOE8KeQYGqzltMF6U0lo2jOw
4ksCCcMYDp6hm4arI/nWbJVIjin5k7vkUshd2CoVb97A4qlQUTtmF8+CB+jneY4F
O1jszFNTfra9lfz+tBMywyY3uqi4mvYwYmKQyAB1GW5clBA2i2H9r3GGJKwnnaNt
ZxG+Ekr43Kcc8bvUq4l8fWVzUukGQXECJguXRSGNB1C9+VbztdaInrKOf+nD4hpV
EBhOiR9AX9e02Pc7MFdkWddNQdxPM4+Ub+S3ncxy9+DDbIyLxkAGLzYCkhn3770J
zcX/v91SKDLM7H+fcoaKbogLnvtFWEinBxJWMZ1DrsbqZfuc71NqPaCDSBjvkdri
wmgoucKR1kI6sv2frkCmBQgTRLAjtc1IGw0KldJRueLRWrEhhIBHY2FgwkeXlJ/u
Js0h5iRLDriQvYv50CdV8aUuF840WzYExjXVHt2fw4QqMNmswwZYSDUGs29fyhxl
bRjmbFOm9Q56Uj77LtxQkMVoxB+qw7UO7s3PiXNxiqK2t9hcbVGRSqZT6kvH3VV9
whTAhy8P8X3ddRtRMkeYQXJWvNj6Qb1y/c+QvJDsBZ2d2jNL6DOfXDjFLuPoKX3p
/nzjenZpIjyh8ttt4CxaILDFDNedweTKUet37Vt0cnjiL+K5OEexS3omuDRPuU8O
wQo25x3fUKf5lJQyGE4UOnFp0PcalkS9sBwZcPtttWZf3Dpf9Dixiq3SpMnsvmfY
ssSavjSzde4PI1PW9NtphY/PND/41H62+s8qayL66Lt2cv6HtKTjftForwWFZYlT
K2zwrZKhOA/6Up+QFp9rur+sfReGfuZvqFvWqg6swCSvZnu1h68/LCeNQfrO2I/x
IhY7K0BaaObVv48RAx6poCzoCN2hrJPfJpMlj+JONkdClLfC1Bf4qG7hfVXWLf/6
XqI26PHUgQdW0rGCihknWalCeIfWYLge2jfPb9tldpDwVmviEzDVmbgz668Uknu8
mUdvmDibeoNK7ovnTjITNmBoR2eddNM2/kRWfHZexB5YTBvH5Q6//+9NfX/S63h3
hPOHCUlcpTb926Y8sp+pw97vm3wwtPn9CPzqA5CHBw7jZ8/1vnu/g3oMa2O1J/JX
tozna7DHlP/+9WjKvbNHW18wNWz+05eaISTw3Ov8DGkodRsk9Y+XBo+6dRjxxAZ/
lHp1u4FcCdvL1hWh1sgWwQoT0ys6WdpG1WdaatIfuI4xmGngR3jXqRTl2onpzD2L
Qrxo5F8vvROMPlX4iRIWInmwVR7xuxc8qFTjTvb3OJGPWhJeRXhalpxWS4/zefcm
OwaKnl7nuiJoYV6PpIeQbbIDqB6NWXxrkSxofPSazvWq9wRKWxMhoAfgpHQphI4x
RMnNNxU+ezeCFcmQQMSK1E0x4sUe8IAXSanUkGeYe7cvm9ZoxVShXErg8jbc0FdB
7BlV3kCdQBJpzxteCuRxC/xa1cxrkLfYlCcta7N/GfLu/tBObco0FWnlfbP3No+Y
GFJku7j7YG8y2ueKCw+FbBfi31MdeECwPdIkMbNlydqhmHVOyqqZF8l00nb7+7cG
24CFV5vs+Zh+UNfCVG3+OQfWtqz/BM1cLzOYIq3xN352y+xjBGeyThjW0c5MWId/
rYBPwtIU+zsLVT+aCPorTFcBGQjo/sITVrVjcAHpVjSIiKURb3ct/pK2q+mruH6d
vxtQcVXXB2oaCYHzG9dYhM4j2yTymJQLJf94nbkSFFt2sIxzYijdrdqkh432wgAu
vr0xLTLn6uWGxP1yNhPHLfuYBrkfp/QWUnIzX3AwcZf88zRVTtYskPClIawo2SyA
FJxw4z1mCCaZ5SrrqvqkU1cSejc4QjrkR8XCBKscRKWsnGqCo+Rn9tbb+AHyFci/
Uv/AACRpb9ldNi6Lsjtl7ZK16x7/LTzCScdBEY9fGjjvJhfGVMX21lgakdXn6O0F
hAVjCWYWx29VnAnMnXc/kYcXBWWEvdyAWT+npg4zZ6zdNdfHvS3gKvQ7CyzM6CHO
4RkiCEAa9XzNpWNDtqq4lnakm2pQORKLe9hiYt4F6O5wZD3ugbwuDA+6iGQXJzt/
5lI58MWJN6+U3wXSLdajQgKgSiKtalOVmr20/fbGukt/G96e748/rFdIIe4dTq/N
7WeREPnL+zin8XfO9N81AyZcfBd6pKOoyl2Dd+ZxFgYdUvz+z/sKwTuzlXnxGlts
fjvw/V1PN/EgzFbFtpIl7u5YnhLwD3Q9jxCEeLeWxXydxa9a+qZjNBOREA3CcxJ/
QPWFCULrZSN9f3LAK33wVeGtXfph4MM9ArnSm4bYOGXk/dcj5UPRthN1cd5G5VG7
ybM0HZNJyO8fZKTADO7p9pYYBUlliWw71CAhm2iwHflkVPhBSVYjdU5S4/RhqWaV
NKy28FgIH3BWpHE6OIfkoNUw5vk6auIHQjffQHX68FFzOcHcwg6YHlrm/90a78e2
BOcTVP2GbemlzwZio59rmu9XG7+CsCx3uhVUbJ8fpHh8EXgxyL9eLp0jjkw+RUL1
cbRTfVmHXuPrI3Ni8jb+DSGFFmnEFqfbY95Vgi8RBbtPfXytz42o55A2gcrEeRVO
P8SwsIwE/zOKvclPqqJUKwHLaVZH0gqRXc0QE1bMWG5s/JaGINfqS9g863k4QBKl
h96irsvR/EiByWJ3nqFSbuR91WUQgXSBBJYwG8ANCT9DyJ4XAyV2mIZsjAU+LNaq
WROPAdASWckt8+Zr0/jqgRJdJwql3xPrY8to/AoBPIvVDdycPNn+LC1nT2ZjfYTf
QhoG+UV6qqkm8LJnFuT4RwAfITq6OGFW6z634Xi5tvlTRstFRj+ji9lNf23PF8sZ
mPMAHA00TQCQtKwwRrvf8kEDI3xT74Y4DobW0Pp4qup89XR+KW+1MukQ/S6zuRM6
ag2/Oer+/y8DydFf+GKVD1Zsct9/MPDThm3rVUAoLMo6+qe+FTJ3DnKtYbNfERZD
htrCsMzy1McwLAFERJeWwijn+ZppX0Oxu8MdQnt+DE5bELl88Au3zBCbiHE/FMjS
Z8bns3vf57D5wsuMc+y8UwtE8cmkr268xciGjEUOpFIqa4iLXBTuaqaO8n+AT0Dc
1UFkWu1J9vJFc0LOCUkHTqj98LslBERuLLZcxc4pKJ+Pz0WaZRvYwj89btEhuiZl
qiyPj4HX/xlPAnD4FG/qaijqF9JhS3H34ePIqS+8L7zsQanSs6VM+B4lZsiVhcUZ
jZcXC2IOUIM1BtMdB4W/9iD49qpegcKtdlDCAgQW0dmHa+kRGmMlToZWV4Lbk9IC
2UfEVsSzk9NZStvFlqjxpVeaIs3J7eXf+t6vzdsL43Kx2EE5pS8QZ4nSDGdHJ+4b
clkIp3Sb2TLJqy6Ms72vpRiN1/dkj4uzpA01GVETPFvll8oQRZzWSewWTPclFAu1
6mro2V3NtMpm7OsIuu7xFJn2Oe3il2ixVY0uQcKHUZv8TwXUGn8WcwH4Z02wY0xL
ZbyYfpGAVG+oEGKVPAAO+M7q1mNNCLfRRW6aY7s5QDwWQTkcbm4LrT4jViS1B/Gj
hEKDJnEBHV++GbyaSdUjeV2CAwXiXxNdoOCcUskeqTne5Q4rdi5zQMk005crDscC
vT3lAvUYZYsRA6npYGOoweSAhdaPi2ozlwu9QyP743FsbqbMAakzYt4QeaOoHLVN
Faiq6z7uFKDDRdXgp9hZ+NUCAXcsw6e2hHTBXnB5eS8q5P0m5InxmD0aMb/B1vCq
EkVbUNp39/aFfBsinD8yvJW1ThWoLHP9JSOB7u98eGc7rBhLzT57mDNqaInh4UcZ
Fm4tbdQ8UqA9f5dmpZ70h4yjUFTVxYoc7SQzq11dCam1IYwZgKM0tdOavM7VsF22
Md9/PhPr0j7Hj8xov910+HqxO5mdaaHzNJ//KG8Mo2eK8jkpgQIVzGXuF2RjO5p0
GyPiSe8uFAMmEiRpcajbJD3SFHQsY+0isXcl3xN0CNLxWFfIoFqKV2rPqvRWd2nr
Q4RgObujyqmyZop9B/tCcYVaH32EgsIHmocQj8AQsaw2T75/viC0HKELAcKj84xV
Br85qlvMRNdyoRE8lDiwr89O6BFtNLDZ4xHiDlnM2ti9FImDkg4Ppmot72tfG/FY
yzqLZEegyFbAolhwggoIkjQVJcsTUwD9YxpcMMyB3eThncxzKjoUK1pT+35NGQi0
cc1AXcIYcD8CBWp8lnhHj9N+XQVvMGoZkgpo9qigubQF1BnBoGz4OTGRC1LW0aHp
oW9zwtbxNUzMHmW/tet3bkxVGo6v6NhcLr+s0EBjIKqvYsGRsKhUu1jQWuHdGvaY
3qhWaTgvOKzW63I/fnXr6EA3VzhQQapgtLJQQK2BnP+AdOkeQUSg0D0LxR1ONXhQ
0D2prsMpzRoaPdD05cobdjiYYInkg0Sce5kgZCJ/M0aj4eXpsf1Uzdj6HiSXTCbr
MrnAXtS8AvcTU3VwWX7oZ/WjZep+r8lVpBXpeuPP5rsuw8PiD9qs8+5b+zZK8cjg
X4ITfp+rRCW1kU6egO5/YK4XzokMfruuby+Cqeucx6obmTT76sK4ZkQRCgimNtQ7
r5RWMMu2kLDnGX78AFyUciAWiJu+Xqi+9NiIVIS3niohAt1X87k/pD3GxBH90UTK
gM0YT5b6VN+CLwQyrBmypdh8ymWhBqF6WY94zdlmKWIZfSly+Bv/Fjm368cctSEi
bGzFACJkTjnbsb9zw2abOYai3SGL5jzKVd7cVHTrR0a0ZCAj6AUvKR/XGw0rtbvS
M1Z2b1b+n84tcOHHqYw5IboEtZjY6sb3D0n0g3U4Kqoak0UTv0lNa1Ksd7MnkrmR
7toJ3BzQwt2TijlHK1u4iiNMZ1BOPK9dukqjkI7STXFCkMIPsAY+KMVLMM7JBFDl
OOh1Veq/cqUam2TrlWSW2vCZ1ABjpHBHJTLrQiPu3FLwr+ohaC8TEFFecKnN5P32
QfiAx98c/g8e9HEsUWL5S9IanAeT0+x7ADkm6sn4NeXyaE7CmALYlOHAzH1x7at0
ScFb66Ow6BNlJ95irkkZAL2Adx+TfpnQGPXQsEF64mM/nh/0ErhwkbyW6KwvIsIB
sbktsalTkMYeVgpYiuLCDsdum7TTxs1NtJQojFFrtZiSFFRMiLzW3OkRBiWRiM7k
6ASXl/lPkzKiUiIFecRHH10GyyKgjiThqhBnX/+5jiXko6NIe/D+4O/sSrjHKSgx
sNn06U02uOguNrjBWxRBX16SUAWGMlpmOLLtIhU2E1/NwPwMaWW1EiiCu0jNRqMB
cdV2s81q0snA+EHtyi0zEf4xFgr3bEhFnkuIR8DHt0rHw6JFd2qEC6+lBlUFukw3
mx+E8tCp5/f89v5mFPnVVEpHujCAbpiuObstszNz4UBWR4mAagTImQyLyS+HOwRa
ZH9rDpbQ9TXHSEVT1O9STuF4DSywti8mT5Ca4zfiqhpTM0RtEJ8PyHbZpLPaozQl
/1TLiTAgtJsM5x6YhDCpo/ed4jTc5UGku0N/5Br7JTliAN7sQ7UinsbhTs6GD8Mr
DAkcGo6GzFuDRHmfUDTetF5HrbUAtH14KFGqsopYfvk6HUHjnTglHSeuIm1/Z3fw
rMrt00jEIZFLMRlVPKq+AOsPaccsoH3ajQjYw5VikxwI0cy5Ajiihlg8ppf++8fQ
M6m6vl5s6kMfEJ3owKoIYcL5ebda6hfvPQDTpQ9iE2ctuJUeq9nX+cP+O6GcwfWI
GJDNYvB06P3IOtaLgJmVVnjslG90e1h98A5WH1SpmAJed0ipvWtDvI/W5OGdgBrV
/ecZLqW2N+rWMa8IDB/aJGELGGcgQikolhh8q0pf4B6Zna+U5E4B2vmvLMuaypHI
p4u16DO/LHFQO3GZ8Gk+iIZCUxNo6f9ZvX0dPdn6bOeY1JYX0hArKddD9Y+I6rbH
RI9VL/dAmb8Brn60tC27L3BoYB6sLYthDQZ2BAoJIgpDwjezxo4P+3b0CcNPjwLy
GxRGZV+/iCvLZ+uI8a2Es7yTmTb8vZmFnzE1+ld6la85/ARjzIAhkw9mHTeasNhi
LNZDT59nofmoapDFOsv3ZoSN6wERhbPeQY80TAsRPz5JPB2wAMtyNpEy4BxwE4Pt
yadhB6zUdJr3GoU4dmQfECTBeMWuGCiAwxv6cbNCr69kRe7fKmmL5fKp+11eIX7i
89N5q2Xc1LRihi76OasSXbhw6jjfAq6hbZArI2NE5UHoamExMT6tqRNKjNEJ/Rv/
IQi9DYXUmarLVd6PLYUu3yHS1UL0FkG6ZGyFMrBBwkm7OnhBiLDa+RI7B/lz8asI
NdrkVBNlCCUMZLJKvPKdMjHHDgk3/eH73sX/7xlEJw+uGrTJu1I766Pk/e6XMnhi
0NPogYWqoEmcmPg1YA9qpvDNN3M6dl8gFew4RIM2k7Glt76l+0qO3xmhzpWwV3Nk
XiAnBJQl0ZTuGcbj2LMZ6PWBDKDqfPXZoK5fIYAdss6P0NHqpFaOpbQS5/I5E49I
sVUrxWhGth4Sao4DNT1/pZWff+KJIVFHcX7DiGLnX6gUftoXzbNE+iK2+Phy474t
nkqvqB9gc6X4E526+CWPeGIGyH2vTFscH7tHB86Xq6jZmNY1FQjBL2LtP48C6QFr
NCOsUsAv+JQLQgX1N3f0X3jp2XnGhq8FbyPsxvTs0OGAcUiOlPlj6afGdMHd6bmK
UvbVZlxjUc/FmO+NMLkPpwCTtO9xkmsrGFmi5ARBGsljvvqwExCVPz0eD98YQQQk
gh1MLtlGebcyfCbW/a4L0yYt8U0bkk0/reRtD+h3RmMBliE8zN0Ug8zi0rHYiK7U
8TuY7rS6SNkCjLiQGoSNB82Etd/tYIQriV8dBjxYJGIGWL27FJ5lq0Prk2iMhIxn
V/UD4EPAt1gmO6h0XCFrpKDNbIbfHqmiCfzrFBi4qOnQW9kPTdEVz5hOw6Yq6/ej
rFIorH8+FPDMj92mPP+57Lg2DjxoAYwzKcnKmKws0JKoII7G71yndDd01o/fO8Ro
+eYdAD3Mwt0iAHFptPtfmAPWeOT3DzBacntFrk5C2cu6ZSexp+N7vNWTSRvPDkVm
EGZG5ikjaNwYKdhZVaqm6sFkM23ei1bOc0iMGCf5MUEmdUN76DZJXv0+A6qAdJ/0
7qpWSpvC7CyD/CE6y7P/ypd/P0AGR3uRsOYdJO5avNqFojR+JTq9QCMBDGAn3B6R
FOdlZ5v03bRuBO7d9S+HKBCq3laT1zUc7+Kn9TeV16e2HtkjgWgqCDQYu3EAk+hq
zeSRKWYref67Ggpx9TAsV7T1Iebr9hOvyWfWqUJkyhdbcSFSwOsP60udGAzz0LnM
mML4O9/SimwuZ6MCKtrdWojBmf9beplWquKQWLWj5QaZwzJwR1t3eJ9hv0idrhxR
UvxCNrk0YTQ/RXRLojC9sJQzqcDZxYYpcgcEuq9pQ8SGZeDFbOz+iJXzA9DlNZU2
hNZoK5t3B6TJY8wrxtzMPSQ3kDzoIki4hUu/HYTi5u3eMEEHj42qRn3BVX5QBn1A
4gQTcclUp4QUF44Eob+UJz7oQdA2rc4DpDOl+CF0rsF4O0G3p/3w1rfYBI4h2pbZ
zrdyMuAkR4LX+279XaPiPjjHjnPrKj3auOGpkzGHYpuauVcuomjZMyaTaDX6Ujwd
O5eQn9jB+CaYlnq93RZWvVtS5HkePFBQiR4yFpHEnh/ieMIsyUIKUFIhs2YazRL+
8liXrFVyBy3R20llLFDNc066WPZGtS7tpS3PUOSQ12fBHJkBsmCAYOtgT6KGvXYI
mTgpUVevzIr3Pfp6uEJXa9KHotRQYEkZhQvJ/M1LAf5ESIm+Bj5La4wwRbdPaPGY
7RcpU+8TJ+uCTMLXZUnrGFAX+prKf16a84vaFDjJE+XPESPpjsBUVmgwgq6Win6G
aQ0FE6p/j1kBULejj6wsaWx6A8S8zyUQvZD4HDf+0ohjGNc0hFNxmc5m8etRg537
LSQLVvoZK+AyaXjtrsCRGnfBdT/PPcEeW62VYrsvIaQ3Ejr/CCMc2u3l5xQIfV7R
UwGUzy9PGDylht2vjCcBCZC1tplXI/ShAJy3k4aY6znJeYPSsUsnXfjgjQxEdkz9
zj/rz8GSrWPjRKMNsd1/UpGa+AcitBXFYbJu44KQqfk8eIevZ7Jg5qcpsXn7tiVP
M2fceAzPXWF8IWVDFXV930j0EMeP8Vn9/I+WwD3jD4sEmVldJRn5Q4oMamB7RRI1
vgdDsXn1U1BUckY4eLKuqTPaPrCYW4YJYs/0y00A48U0/vV4CjUwwu8vTSgXQmAS
4IqbRNkd8SpiteubYDygNQNMGNn+O/00BSjwLhNvLciG9FzvNVIYOKy9kRokhK4N
hG2sR+EIZMSfpIs5cix0xaKyK7bxQAH9thhkKv/u1yATXUhtqQjlK5kO5bUaDFlU
M1PA8O2GKPq7t1V5Bjg9pj7BwHgXA1FShiWKpdckCaabLyizqeLRXRLoEP0PuiSt
aN0Asza8Vd8hanZp8rNcQNsKeoJ3CmMnZGVyuywpODouZkvHSk+FYmWc6P2hv5zL
MtU3ukux+Qqc6M+0nB84UIGzCnrgs4OHREMY7/4cBPn8EJ1/lT76PmjpysuUu88b
WbMJ0gdu88xXUGo/j4XKUy1LjtLxuRAnZjujC4PPE85nxdl8LOBphLUPXwQjfPbE
N/JZdrqaikrPjaiHOckS0LO77XmCAtQA4rpuZ8rq+JWURI378HKMWabubUwGFkoQ
1SLygZcBKkNWgQjXPlIxgw3djNNtVXdDNTMXLzIL3PFOZBIFZvJWv7xz2vkUlLnT
milPshzM1pWQ4+f1sn8uJs7npBDs0tJmWkjj/QcgC8v7uW1AXxiI7pn+NQNUA8lw
YIwFFgKM+rY58xcz1zR9EZ3iU2gI5SdFIGzh+N7HRPScTpPfc9v8oL6FcEKjR/AT
zlGZz24474V6sUF6ZH5CdGtzaqX8S6LH2rOX5rt5sxfs4nS1xb9R+h4hQIyIgFb/
MgSFkKvNLkQI916PkgvsW36OhlCvc+RHDm6ZqAPVCh5OfgfKno9wFGzmVbHbKo9e
eaKkTVWbyzHhROk5lOXhr7SgCiHQjXZFXtnBn6awMR58/wuLAR1DEtxJJ0TWrND/
sy+RyHMizxjoQmAB93RQwca3Wclw+lYV+EaOAS9JHZd7d2uGLC6nXHzWzU1S8rMP
Zg1IEM22i5lwcQ1yykC6g1IJJOiO/w6wkpuAqcjd4FKIHbJc+ng563cM+bfD0nhL
502n0HKtvRx5PpRgTKZ+PsEn/pcaMMuDhvVxW1NHylbA1AWj4ySznvpUDW8Xn601
faxXwQeStK0xMNLS+aRKNHMTJuGRx7bR+oynvPee/rjpjv2FN8aefe5fPli+89eZ
ha3d19gNyYvYiWErsKc0rM1zxhd8TyE1udXZq1XbnB0UjIiY01Nye0vMQdEOU5+p
xwOMUFGA2jve2UM3Ou1eYGkR9YSs9TQZVEyQwslX2AkNAQ7VvJJHBUlvcjCl7UOT
w2D0OkxPbn7YkSHn6DV2FObQkFuwxWrREHOWJ+wRYkx7uT17m85FIc/UhdFRESLG
+yXdP36WcXfEbiJ+p9QwvrBCgmrwvBEdroGY1GNTlUkJux34iXLWLVBycFVQULsC
yHGo2U3yqHkZeGWt/vo73fyG8X/4Blg2WhbchlPrsmK67W4Jz70Z+t/Gi/dL+pgI
VsQzz6vg0e2ExDnQOpmH27e5iilXYF9jZzGj5uHPyp4furYx471WDFzsbWSL/PFo
v+gfnBIJjAWe/WKNeB902va9BrQHl/Tnokz5Q3E2X9jFqsRUJUTk8Ul6wZ+SWIzq
sj9ncmdUk+9Xshym/MycEN47Oyv+mqxkm7BrXIP9IoI7HnSD9ZvOapwplEFmLhz+
mOO6IuNd6ycrLzGK1RVbwW+9aRc5DSTj05JQoO1BO1VsdZFiYAXwVPzD2TrRAeHV
M6YJM9Ou6ulxVuvDHZYa/dV2waJdHr8lod5uaYQcNTi/RKH1OsQ949DJiOjacPpT
7DMZ56kV3ixo+6NaAQ+Gr/RHj9t+d3EqYWdgDGiKkZlHam6pOdV5dWXuJcrlXWom
dPBfDY6lTLv1hhhK6KRJuec3TMqQ2uq5Fk2zuYLgwgOETnC/hpYIidi/CzXRsyQm
RAZeLie5PtTaJNa8YHoiyvInk1fBKwQcix5SHXbCubi6HCG1pge8/o9gT16J+M/b
m3BRIH5lTMNfmvGYh4xsxKyGk1meP+6RN/wS/1TxgD59ZpOrTXDUGZj/vCx1o39S
FdI45A3VLMfvosC4IdwqLmookq8OZB2gdx9FJ/k7o+U88IQG5Fa7FO40ZA30JYzi
mH84A6Vb8IQR5vsuT3Q8KvnIbPQYblpIIkhHhBmVRyk5im0qht9yyAD2rnmDFDe+
KDc23K+rJUjx1LNHD4H7aBMcIG+/ndliicOuDAXfQmMj5/b8tUvJGHK1zajva7Y0
hPdpk2L5OLYmehAbym/tZsmkPE1hmhcfKl5ny7Tg01Q2VLMf48F8EdnTnL96/+zL
/ao09iyvN+kDsFmYLl0zcYq9ktJBwq3MB8jokHu7po4oS5Pzgg7bgzOyv/fgBJqw
4jCQYq5VhiadWyyV0rqV18ErR+ZLpzV7ap5dghNg7lu3tq1CuEn+uVyWdeSjLrPu
v9jWvCQGKyy7+Mae5cewOZA0ifG1UlYt79TQe1lyNXojb/SBCF6q/UyGsf3qOoyz
SP3CvqdxbWa0XDSEVuMHqvO7C0G8AEbxRYZH3da4QMPzSmNw+OIdSHIf2eqbfyoo
1TDLAHy8gqM8RhsnUIJh42QyfOiAXyixOXhkdKYhaEJiCyDpLPEzKo1yB6pD9MhP
hxj2JhtQQmCICIYLGN7E+7ymBCWbNWC09WxvzcpWF+a4sSDEkhwC+/bFGswyPtg8
H5Y9VsmxYGLwtKjmlPVMmlzEyw9p0ouJHwC65Yr+nosb4fEIIl/A2W46iVjRaRBu
Ga08u7sDRQcwdleG1LVkE/rsXmxZ3I9KvzuvSCEqMEiGI2GdmrEi2tUHhy8QQdBP
wCzdChYCmimCOosaqF6xCKgqJdbnCQPvYryOTRhP9nCQ3LBvDvwkn5+kZ9kZJt1X
gMJZgBYejtzW4Oww+9hsQSLeBP7EFbYirG3Mr/2iQ+uWAKXzqUXRPJy2edaUMaAN
3cso8ZL/6E4eQ03khqbRhG9559gTG+uckzrs4nTIT+3vDvdAfXfmahb+HK9ukUwl
Yt0+2qmp08WjlClonImcwRcPpUduunXUlu5kyrNLZeSZEL1jc6Og5NDBkoVjF9Bp
27Y2IB4X9N4z9cHkJwGo8XPiff292OZqgTSoBtIQ7XT2M4tvAViGGOPZnkoBP4IE
arxtPELMbKY/DIk2B8OtEHS/7ybiMsdVej75ticc6QPliyHPM39HoY5i7FWLxNIs
5nF7YFx1AzrX9TDxCGPUdUjrBH3sKLblCjy8IawNJqFM+f7oJrCRSol4aUejisEb
UN8+mpR8FrVw/162AhZ2m/J2YhN+kJytv5zIrJJunflT8OP1qxeHFaE7amdW2rJd
35mLW6azqJgwAbsSzfMsQunmp+T9XKf8z9Dw0Jgn/5oBBHSaWdCK3VQSYIKWRKRJ
Hu0kLpjLFmex/AfiMXJKy5yWMtnc/Icytb1rg5/oAUgSKfw+AlRPjaP//41qbaI3
sowwE6VCMawZJwXmfp+RfayqRPWGosnYN48rdc2xBfEO/oo+j8ShfPICuPC16ecl
Bn/RB8B+2WyW89+lbFFeGIYwwX9NBRBXZSUPvKqsDkoT8vOE0nqskRTZ+/JPF6fH
1B+0m4pgGh3RQEST0l4IgP13eiI1AlJsYnEdnEr2nJfsSChfy4iCsDEtNtZ5KIwb
z7bnzD1t1IEJK/Nz73vT5vjh20VC5pGyBX9xG8YAkWfZc58HnIKf5NKJ/xOOsJ8L
SXpq9+H3FAqhedrTLD7/k2stDMCZA1X7iWGG9JVT10DruoborfVVI6hAjVL6BGRL
2E8UcdRR6pvkmfPiJV5j8t8CUtkq5xw6tdUSqfogD4b6fHcNTHHhBdT+SgnkP7MR
J5adfVK5t7hmlo26hmT50eeWRQPH7OKh8zBdFAA5JAvHaFm/rgz6GTohTgX3wFHg
WnpIcD7LssgPmJHaZG88ezIVeAfoj2LB4ms0R4oSwTwBP//AvU8nOEuasbBvgNoo
PbhqXjxcT8iMtJeHkAj3IWbJc4FV2EL2I33rl7Ki8ieTaP6Tq5z1mne4ie/T4Y68
UxCzMl1ZyZRiHaFQZzrT858CZ2S68on/yDvHcEHSY8mYCt+ae8UkQUDEWPoKm8Y5
wfWmho3f/h9gZcCDxk2wGA339x7UBWeLAC0+iWAP1M+j02HwQw7aUv+dui3UctVU
pq7Qv0I1/3jG9bbpfbRxlZmxhKr551VXjWdipUzC07qCQfbrctyeiRStl9bBEu7I
2bOILxrskmCshGNKqpFQkR2fdtgUKNI60ImgOfhpFy3jq5tHgGDaZ+mfEwW6i2Qj
gO2XViHEwCuMG1K7G25MGHBcHZqVqXIdWd5RNDl6GFeD7KpvXi8NhVt9VRLzNFcm
uFy40m6q7yxaHL9Woa4r/ZNHT04N5SnvM3nDqWoNC2HxWbOC0JCNvoyfnBvNNgcD
XvkJ+pj5hkUqm+km1e1pVVOITmPt4q7wuGJoseWG/Wic5bXPk366khTLvDZzXPCa
RKEoA9VQzxPuDSgLBK8Z9im4P00b+CS1KrHn38WrvOD5K1Hf7N42ifOXMjF+BssS
8c1QbpCgEcJzuSun0aFmV+lGdu7tLmhoKTFUQThOOfwgm1gTHdIyfdob7ANyFcnr
xJvoOVmmeYzcjihMnzkJdaGs3rnUU1yK/D5US8RfKKkHJX4x7ElHYYaOPymplbY6
Ymbzn7yk1o6fNTUFusPPIFsgKN9F+tJh9wpzLdyMVeM1T6UcvYl3dGMyZ0TQh3E6
oR+w3RNNoifnsh5o5vJuUXyFvUalaG6fz0VTAnEicsYGM3cLPLM86l+P1OfIBFmi
zV2cgNeUf1LBOBOEaMCZ+GOAtwUtUP8xIpzg0RTWA36XAglo+emNuVNFpNQnwdiI
7tFSn5PMDgMSKltsZILrKQ45wJQHyeKYSZd77xvkjtXKvOz3MX0+9N+O+BL7KENf
98R3Hbh2uDW4NeaV6G/1N8sPPvKiiM9PcLHOUZZmYrUtyvg+X502VnFUzxuVgqQO
7Z7uWYSWQYBM0DNvmIJ6TPFjKszDT+s1w8RMzRQjj9FeonuyHL2shrxxHC1W90Mf
tn5ZEYLoVu2RW8o4UmdEZE5vp8BXlcNjzt3FYWZHCqM3gWq3wZQzHUiT9L/C8n1s
7Ntqj/RtIObJLzOE5t6Ax0EpFNfo/HhrfaxOt77HMgDdvmSXwwoHKl6xNriAASNc
2zTe12IwkdDTDckeQIt+iRQeHbOd0/5Zy3ZkwCli/un8SpycBByFrwFcwlG0vQf0
oR7WyhGjVbIhKgzIV9/luTazE7ZJE9XI1iUXRrwHUF68PKqCXE6tg/q/c/++YMdt
BOHbpM1HLs2khJGeGNXRIS0oXoiH5kKoCUIGHLCXBdQdP3Lm1k5PI3zuYFnZ3FEF
IP03otJvlMvERuAVhjw6b686nFeot2foCrlFusnBCOtLvVM77JL9hrTdEqSN38bU
9ZUgN/gzp4Zqy8a9B2k58C9uxkHpg/w8yfAc8fFbGQY8A9SAxq353olJ9LpThPSV
SLS336yyT/uhVEKE6/YxkRAodczTUPviP5XmrwNsJVUJABbLIRW9VQCLepC1LyOM
3MC2w36ZLAqVriU5xgKaqJJcIrK5tZyW+0d24v4+a0G6C8BQUYoN0kHKm8CsGTLY
7gBEQkX/sdU5ftZxjWHbwFdpsL7icrhzG2Vl9enXXdWqyD9hbmXi1WI0ErdyDASG
8KJDLNbEMjsqFpVfHSWy1pOcGJKKXAFfirwtMhuyec6oW6lTTLv1/ywYFM8E+Z6Y
ABO+yHu/Ms4RGzZnd2gCQSrA9xFT+6sK/5H1vbZlz5Lr/s0LQsfzauc6I0v+iNrS
/BzKeW3VRdbN5G+k/9vyyl1cGPuoUXXrX4Jmqb2lyJQi/dyBNoSgL6iBtY2w+pxE
9uciKQCE6parVxXEu97W1erfG1Hw5y279y6ydQ9SHE/aCc+a4tEVm3ozhKKF3hK4
TgCUgDUzrDb+IAExU12BW0phvzgaUTxOZanZ+eYWov+CnhomnOBflzqHrR8wuBYZ
ple/Eao2svjSx2Zh0/lqQ6t+WZE6F6UejXPUxrRPE0aIx6YGkbANRsGiOetwyNUw
eSkyQ159a0FKYKu5xLGiraZJk/zRQlaQeRVgdak0PIt2ePLropHSKDyyvx5y8Zt1
x7xmehbEaD0XmlE34F3RdctoQBKLZBq4pngxeDTDBVXvk9YC4OI/7x+Wz8D9Uhqr
LPsUOXOmzgQKGu7Ql1F9zPr6Xha+LE55rvKar+g8IOKLpwHSTzOz59FkZGzE2R/f
d9MNbWqXg+NJXQElpnqT1vZHsjnfKzKxd3KnotUUN3SqW84hW4NA8ktZvFW9skDT
lZVP+jSUt7OimixkkTM3xXpJWrV6p8Q05CRSh0ePVpju/6RgWBGHa38vtMO8EG80
sIL0JsECddvwCF83H9pCY+Chf3Uio5vR9hv5JywATByhChi7izsCS/D08EwR+6iy
pLIXC0PVI7OA4I8PAWbTgJZiYphkV2GcenH7jk7HMB0dtLHRfnGHdAzRvMtYUsDf
wv0bBEGJCSS0yPJxGjT3xofvKT/Ga5xDL1MJbPlX8oXDe3UVRHHWHu0A6qsTuP6T
GWLhRS/E8qtWBgBY6+Vr4nzFpMZsqq3lrErnO2uU/oCQ1SFCHRFJIgYGegYmOPic
PYEY9Uamw7pMY7dPekVXflzVt7tc5W6oVaBnsjJ/HhVj5TrYaZKe+k5yA29buLx1
/JvNPoU3CjA+YHKMLfZQSWpu5eHkzK2dO88TPlos6JJ2nHjeJyvlAOzTNPyqv2pm
qXG9Drl2c5LRmgTl14u8VySe0q2S7Mc8/mOpZdBqZyFxykijlI2HSIHujkL9HApV
ebFUsJiVEWje8D2Qq55Hsx6guuYSzb8nFcZmncRUBhkqX17xRilpc6r5fqi8m6R0
Uwv0CHnSCndUn9wWp1lSO3mV1zQHfRo5P8DCNMzyBu2IeK31MQ/4KO+yOeHFccvt
DD8+s7fDZNXemAT8wU+M8pR+T45+tA8TZo/c88zozIf/kCou/rbTiM8smXb2O4As
+IMf5/IHGkUAXfEsrWUI7nAKKXoI6YDa7izVTXd8R2kOTL4jO3DmheZtr8eq+6rE
jpKTD1/JMOD1bLWFc0GhGjMalwP8HRfJspOcnCoVw6XrDmjGZGHvAYBe5qUl+cpH
diHhK7vXZokL04kernvThPQ4P4hq0fRG4QQn8bnYQnaM9ELl4AhpmflAxQhHssYK
k31ZeNq+LAjmIvfWfSA0e1yBK3l7LEXhHP2vJ15zxNZuBey4576lo/mme+rl3K3P
L6yJ+vHbBHq3CIIjvIvFxQI6WLnuOpc1O18UPjMZa6jyLTYz3KqOeYbc8xfTeKIq
x78goQliKYTsMkogHraszY1okwpkBXxgb78WIWvFvlqaTR0DDihx6cAiI4dUcDmP
adHCUuoKqeaM5JBIAKijaadvt81isg1Yuxy2jif8cMrsjqcYAxS3zI68EZIuX8HZ
14Pk13m32xHbu5+x7pDCb9V/iyFKc38Rg2edib9a6c20un8yFStdyhzpUCuFjTbe
IHJ6LZoUloNDgy7Ygp8t43/EEmdOelsaHmqkXSG6uDRTYc0fyHgAQl27JrJ4Vt37
KfOIOEMQ1JyI2obEcgEtq/F6FaCOHhg7MU4BreQA3cBmxropPpX+xujiklChqU19
xiJ47bDDg75/+/sLCfgrRjxSdHfMMm914SbdA91C1+9+M4NGbt2FQE1en0Aed2i2
aMAOv66NRKNlFxwrCjLbjLloTdY4IFxAG9Oxec5E475uE3MF0e3H5yhZC8c2UbUR
LlR+gvqnMCjahhJIevybZBK8azC6llSEscbSExvuBb/SF6+AMTafrw69cXpiBczJ
656Yzbj/cHxYRPj5V+mauqCHe3vIK4kfOHi97Vwl57JB+/ny65S3dWnowyqDToA9
ADUz4ARmx5a+Yjsg0okmnXz+BBvcLj16JqtQBrLHKnC0R0WcUziBjJa1KWjGdkqi
o2ve4vcEmdePb5JarWTm5k1KtfQorDbaOB/utn3KXTQwyEo5kVnCvMP1SfWJMddL
2ccgl01TNj4YStN8malkfgqnuYJ5wQWJ5V+tdxB5jCtGVByP8JW3ltqk720jMTmE
vI1K+x0dcTbluaASwcb758MwdrDEccx9ijkKfo3z7oiC1xxEHm2373NOBiZHonlk
P7OQOl/V9b9gGbwemc8d+y/F/Ez5qhQwqul9Ngi/cTQJ76xXdpG6xxMP/sHn+JDG
ySMF9tASEhYtABdB1RmfSlUuylxjVw6uLgmSU4HuUXhjhMMV0ayqyxGYYKa0YafS
Q+VfzPQpqVyrnZaDIA50mobtq2/GVlzbk61oFcU/0v7DxIaTXZzNq0sH9py8kKAQ
dR7Y/F4kgNXHUEAJcypKGw6eXfczOOnsWxJIXOFzTA7UEWxIhFy6NEt4BW5HM9xW
LK/VwPJo+Qfq4TZXA4gqMKiF/MC2alNJWGDgePdRuBZ86s3PlhuCe5g2cHWkGn8j
px1Tqn8Kp3pfkfZ8cFuvQ/EE+0MzKb6CAWvLd6cudc2qOQJqgjDBXDhN4+rSdw5y
um11wnExhLqERb8MUU7NeAoKqGOuqtN8n6yA07oDmI09WMwptWZjRGg7Tu4MRu3x
c07MoG6DHy7PGZYv+WjgPOggURlfIw6FGxrlHwxfpbHRuqCLhLUT9/Y6ABcrodSt
arpj6K8NAG4ETE9UZPgW4Qor06xz+KMu1zFgDFtTE1AEpUYBBfaeApxjVJXJJRHm
EbjTbJNZUX8588SPoVvNhE8Wuw3dBKElDes5m/KVJMrlTbkV9Gv+9VAKao/Ch1Ql
O/+spbp+cGbTq9gurrZo9oS5S2hqL5KDF46oxcHURJn7OljWx96uISkbyzPOIp9T
G2EWIGHlwSJMoEp8kyx6LEKlJpCDHWYfjJniflIb+1iEG2SX0hqY5EWb5tTnH2an
ZDorvL5FSiFGE0/P6bk4RgRBTQ9+0mIeHhioTX4MJpyGcKesnIzaPVKXP5sxQM8A
BzXRdbzgUoDf4Bh7JrEpSKNtuVahhJsQyGSKZ/lnfm1fwEGsVGWeDxD2RCXjY3aZ
cUCLlCdSmWtLTIDIjz/fgqTNF+tsPMSCyS1dL0yVwBIcmymHhGHl92HTgvqM67WY
Aq2jZoG6jfhwpJC6/eyk/71fBWS11U5COL+VSXbakZvluqEtAUNXml9UMqhLHWtj
3HPN6wlRkrZDghwgxFzXLRn3btp2q8mKA6rjIHqi2KGffsup4nSst7i4fj9CRE1+
YTfP/XB4iVZGUdP0QaBGKf4zCrz8h0HWpeM8wLsgKzxx/dKbMbFG2WKONpC9Q+MF
oOnI9q1pE7X0hIgLmOehm8XvpjKirNgQ+lSm73aptQk1JgWV5WLd1pIrpKGq/1OT
GmcxBiEJI6sM5SNeCsmGGfhtEnXCXOebBMY1xfMaS6EZvUNlcDqP0oa3sGMlnsGJ
TEgwikkddMzd6IkW7DVd46j1+6P7Lwqp8H39mq/JkTSazl8/lqr02XcEmgz57vCZ
CvP4nOWEyHnrg6FXs/KmBaG/I6BFdo1I818H+aU8J7Xl2t1LyyeJiT/UbXMEH6Kl
6OOkqJN9ehYOKJE7OmW7BWdsL4b3WgLppJQeHU9mbhjU5ovMpHyi2XJHJHeAdw01
c9IrCPnir33cK1c3mDpBTrpFCpKV1T4IMTmhbXOlJiNctJSRJfzj+5BPg5dQJNni
QIsuhx1+YFmyPDn2xUqMfpEOiuSMSqxN2Lg/52j+XgNAl2ffd7JbD+7cKHrD/cG2
hwzLIx+Fv0q+JBtLkWF9ucBwjXVDKHGiWklqQld4yHvPHcgTqZR1fqk3FOmYQF4G
3wIARyig0W5oQvc+QbWUyuYeHxMB+gmhDwXvTISeyyfjTOheFWlT3e0RnN7BmC9D
YMqXRhSBQLsoEfZcBSWzOsUtmvpelM80tXgCiETKvKczU+EDkqsuPbWf4ELZQ21F
vZnahBGGZP5cvQOS0GdE7CjuU0CTR7f12mi0bT4cc82vhIczCRsUSRJRYVOOVtRB
eXzMv4K9pX38IXoVrcRr6AUPVslEzb3CYAkAdtODwyb9UgKuBd1av9Fc1CUc0WI6
zJpVvUiDI0kJQrkCBsVW6oHq2ZPPprfh0eyDyjtSqFOurOw1eSRmwZrkltw4G9jx
brvo8+B6CHiN6/lKm++VbEsesH7vBf4imb1rzlE7iYTyi8XIO6axPaF10H+p4Gc4
inpqZy+ESWwT0/9nL1hc3Eqqamg6urF595g9oyGp2tJdQlGjOaLbHTwtGg9bkYZY
Ujyhd4ciWoO/1T9gRYOCaIvMH7Df9pnLwSzHbyrAOQTMh6Ynni4PzZE1eIxbG1zd
6M2c/s7QQowU3XDb1ZqE0AkcAjeM7Tp+CXTdgZc5gzrWhlvwd6FSIgPUgyh0pbvB
BUGW2i+A9E9p0sVPKjN76cDWVHTT0pNBv4b4koXSe4GJKLYf3lkd3NOr9Znp5jlt
CPXYKHYKQ0KeG8p4e9z+6IoufPzB27G7zFsKJZm0EyqUwR04JN023xEiwGLB7JzE
vgzPnWfIhQHTXIhv7rXbfgzivn1/40+ngyOzSHM89ZxtcwCp4+oyObLnYpX3XDhJ
1mBImi1g1kn0JcjU7iL91FB9KyBpqyTJeFWudL8dlPaSNCNgD2FRUUzJjFf08nV3
Kvw7W75bJFeW/Ty4eilmH6OQ5nUq3MLucqaEPcjeWh+rsfZpl3PIPDyFLPYC7Fo6
N3GfQnSOi4FSuLh022EiDVFqtpo9OUQryBcRjleMxYAyjuOnIjynaUj0daM39tD0
C/MMVdiGQUKwrrrCaF+DmAcG3KfQHaa1o9MD8DrtOTMuGtktib2XdMOpbW+p8VKB
0DeTorRLk7QFyKDwSgJdqmjvbhAz5N8Szv5NYUp9TYqcM4sPMt3ZkbqdkQe9af/E
O/twLYlA9IVqt5lwkPXA9drVLzoRrJ4fWUJ8RNTM7bLUg1avcygGipqUXf8Y0BQF
lbjzqWBJZsxRO12aoS9zV5Ak/pHUF20x6uFT6I80Tr+tnLR9uTE/hB2h03e1qGJS
rHuIR/rvHo8trsUUozixOi+2GBQaVxghHcSQYYPhQYKhpeAK9kP+4vUSmpKwsRRM
m2ioS0FBvJC8pympgg2583KBf9JMKnNKOdwV6XZwHdivTf6cfRHo0JWBAQr8TDTQ
zhcBAcHbUavJQlR/IYXnJ/YGwqqZ3V+ggfNxRHFQ7+kbuHEVXcsm5KRMNj9WSV91
KP3eOY/DYfpW8be22b55jIpVgTAETI2rZF4+aOoUVxJupbvXSfaifSM/PDjTrnUX
VOi3JTjRuUQ6yPZu5rXdUwneMWmNQWvq2EURimgO2yhjd5VnKOxlcpneCT2m75dq
pMZMRp2rE1S8rpLSTffAyXJHqJbMmZ1zOjQZWEvRHPG30jTGdQoowrL/Tlk2Q1ft
tqrcgzuw9zgBhqqS+Dq2FCXrvW4AvTcYOH2v3shATP9xIpnee6Cvdxk32AgUapdL
1qJux1MajXrKCf06ajbNro3ujTMX0khPWLE77FMj+T1oFzQO+o+xR2RMVFfmll2Z
qVcPLUSUo8fibBjaaGHmxtCGSQNECfS3d5zOFQB4LkVNv36+35fTcvjmauDfJbTA
qNK8LjeNlK94m+DqARBcZwYDUou+t+XQJyT5Yk6GGuEH+y5OMLIQHUleINv44CWU
rii/tqddZ9nyYJGMq5K1gorU7oGMywrDPlU5t3E4cqFyhJsSkwoVHKVpNcZm+sZO
eyN3NRwOKtyYt6U/XDjmJGL7YcPni/qK2HRKymR+Nae5bkTYxBhXHdFZSRzkTTk/
w41blCkuqZZrkmNKUnH/bYMbmMoO2dV0cSQHBHR/2gFZP6/6hS3XzPhLtWt/NTXq
woYmlnYuZneQOiiZVI6uPjShkHl7Vp3FL7IU2XygkfChcrLsJxIt6p8fffyF3+1y
z4NYvHFFLjxC0FgCcqkTFAZvWl8nNvLd2S0EXbFwsA8KIaa2x6sgl8oGn4+4ASry
8iJlsl9T9NhKs5PwALcaFtF8CAbXDtM0szdlLBMQjdeRYdUXoddtBA28D1GkV/2m
7BjprroFMxao+PoxvMbb769y/uurcbxIzabY6wUo35HBRxzqJrFqfsgy3VdY6h7R
680THmMupN+dhXvkFIPpcUmRzE79Yt1ZL7ANJ0Tb1gnc9nJLcTU42Htnq0ds7L9C
o+FU1sU6G7lkWxuUbgwulu3b+UiEvL6fXdbwz6jaV1oqz9gZ12pzCNC6iN/JG0lL
LuwEUOcm7ug3FNTnkI8d9LS0mmlOMO57jEq89J6DAzRFxb7Wn14vpwBKXZuYQId3
6AfU4rOTyzTU3Hs4ID+CGubN1KLFmE8GBQwnBIGCPINeZL6102tjnmrxSoQmtY6v
Z4E8HMM/AIOBZycHvYLD2yhVCHBI6mwS5W3WuySho89TaKGmAFeNivtlIWiuQ3LE
7q8mW5x8sqg9blOMkbEoKLkedXd3OUqffwBiwpw+bXS6UjMg/dZW87/vBNHtV6VB
DBpbrhCP9xaWFcRcpFoLC2Na5WI6GIWGL2tYKPMzxuTCvIU6tdtmnUBEIvm9M7Yt
fv/mjSmI843CNHW5VAOGCAZXM0KJU1Ect/k9kIKFrbTgA7Qu8vCuhfzomRZmDoFh
1JLQX6NHLeFbuqob4ZxrPdXfFHyIyOAFyyWU06bBv2GMZ8dtf4OmzzokKyHsdDkr
nGQe7VwsfN+t8sQ0maS030Lz201TP954QNTiD0wHLQC5g0x++MzeLw4QEOQOoVWb
kbKaQGBnlOVr8JboDy6LrpoVXBYkwx/OQrElJoSB9LjehSnqwQ6TPp5//IyDdD3w
oMiq9I6g+6Mlk0MwoJG7vFoWqy/qvvwOUIOxoi84a+9t4YFwKTlzEokinNtJTAtB
tIRlnQ5tFXJBFBJsH09NSMVgQUB+HDyfg2NfbTGFXHJXhZIN14YwaBJbet5t+mPU
TzEYcnvek6+J6mO5Kewe1KU4UbZI2ALgMm048/7ntmsdq7KVmSl7plc9fdQHpGvA
DXgmjBI9Q4/sKVsp1RlOmNCKhd9TQ43EsSYQS0usJyYrkSWltrWv0blLQJZG8ZXi
4A5P4RbW0LH1ctTwPj4BcOb5p7rTOw9bJDcnmdnQ50VRkRSpZEBg12s9W6bwsdMg
7sCzSzl3vliYDaz6wB7eL7A8aYaMm2nqHDJtrWWRRzlJNPntLVFaBZVP61O3gizo
Rnpjco30w3GJawTeHuYvWk3mEi0OXRYYyugiRA2G3m4jF9hRLdEtRlLTgPwWYfJg
AtDGAI7UZO5lttxyJJVpfR9Hoh4uPUNJoFpD4xe6/jerZuOKaTBDNLOUll4uJVfn
kSsMn+OY+Wz+GdRQgfWSqwi1rtZvtHqjvuXZHFD5YbJcnEP+kflMe3LnFob/Vvop
QdkV3hycQPcKsYATYr1teaPF/bA2kY48Nr8sfaXk6f3JViaZdDNhwayjS7M9ZaNu
8yU7A4KzWjVXSUUB9JOiXI9vh1DXra8LGHljwt9W+iZttNoqAp8EurpKO0NxpKsw
Ovp9n7TWBfYD2YG8R6eAOwe8pEbgZ0jNNLL8DtJZoeC5utWhVo54fcBTtRazvnog
FJMznrTpNEPO432O57MHta9qwHZt8NxXBETjqL9KKFlqBehHVVMUg29/rx5yOEQb
AdaoTFefD8/2rFifGI/ikuUuZoRRMMDcwhfyH/qtmrgDkB1vb142W+5lsareGCUE
6uSki6NToZYS2Hf8CRAF6woMjUDgIJ7XqTu5eaddPM0kkhSj6BpC14SHUIWLPLYZ
eReFafTplHFS8UO/aOMunwWSzMcz/3nPEaPqbf2JJ5cCN54B157GZQPRar/ecY6a
57YbRBEIRkTQPmNyNs2QESV9e8ya7Nx57/kHgH+TyeSblDEEB+t57DDwwoM2q7Ur
r/1Xkr+bwrkUWbTfKpxO16fDNcC8CLSzvdSyW9hAel7lTrhHLUyLkaZ8wAsMJcQd
httx5MP/Mv7EIrBCFbi4zOgBjDlQAfvY+UOK8wIpOTbEK2RzGg8wx++Sh+OPbENR
gzklqHzM+gyp+TmRZkafp45eFiOZHBw6xnIBt5gj3PGR7vTmnqqq+flPpBM5buMh
FcVl5Maup/Myy9G+4o3L5PKhx71vf5/jG/z/USytRPz9nIKHUA7OLMoN3XTcG/XY
bO2KOCrFKmpk/gdiAkotRgXLy02g4/l4b+gZmTzxEfiCErnMD2ew8Iv0UuSlNC5L
xI44Fl9XN1mD/M1Efxn7PLg1snMdHOm1wKPinxlXRctFtCPfVDjGffSZ0pLWalNr
fAKQvOzBLJDom2AgxLrgXSeMgb6VpXfNlIOkUbg66rIj9j9iCp4Jkqf9B/pBbVRr
gcfmVKAoXEzPnLYmb/AdX7/He+whDF92c3/8C/j57pVGYPTJIgPZwVw263g45OBP
+IO6OXBFHlZF3q0AVp/n+IaTmc3804m+zloj8epqYkw795JoJ3RUmAchI3g3S+IB
YTo+b741JGbJc/CajGTcIIM7v+UQdsnY6vPS/tvLqSTZcaqZf3CZVCYu/I4Om+c2
WNaha4PV55tUtkqEV8SEuLQltHDSONo4xx5fnZfXMxVbzVsPah+Y3gUn3g8+YehS
J2W5hTFqNao0+JUmrTIMG45a5aIshiEw3w78Ji4f9tdLpXhLK9DRU+L7BjKFZNHh
ck2VoUF0diU60A8iuqRGTYJHMxcC6+Ukif+9fch8NqVnuVQ+BaHDf3JIiYytlbNY
/KRvUKfuJ2NZ03dq6Mh6uODlbpYDZCEpQnSuTN8Ou9ymawBmJaMfjmM1bKylZTXt
lNYh3KjIE0n1kFdYiUHP5D0DJGDxFj525CxWo7NGuahZAG18Uo5d0IFJuf7jCN0a
1KGCwEl+iMKMejVuZ35q/NtLwQtxDeNOC0lWrsvAQCAEzPJgdHcHO+3CtobybkWi
RSanF4i5DEFQNask6YPU7TJHw5SGrHINdaax8knCBEUXJPTFlbgg+wZQeEN0ansn
yaMgeEC+Jd2ca68Av98iqEuFAYFGT40HLQogYRc8HYqyqk7i5rT5Y3DATcIup/DY
sIL7SvIkfDStpnUL7x/JNH1tNZQpaunSe4pylIAwa/yFO2ObU/GbGn7W4tALhq1Q
up4N/+iJpRlUpdUKGM87wmUAvw8AacPmU3PYV8/3iM4PnSoWqNkDiJJQHw6zTKhk
GAsky6I4Q2gsn6mfVoxsBHUkj5Jg27zCYWKs/6ZqgCJ7964XZJBywikJzPnnoANo
9DA0+aNo5Yrr4s6xMOq/KAJ4Wr5zrd+5OvkRqjDG1dtlJ3pAdlGiGp4+flugPTyB
NBRwXUFGPodlrfueYof8C04ntSGMs3Bh35Go0lNZUomrYURtQuVvFhSzyHnsrZPl
+19Ghtqu3QhlFtpF4fdwDUVaHTT8NtsNsG+M05ongJSDnwl3nnZ3FxdeE8vYZtuv
zMb8TmEiyAENURs4NhkoL+SlsNLAHMZ+buHERS4Z3biJhCG/9lAgTe81BeKQQTFg
NZU9MofDxwxf37Wuwmb9uOelOwQYqIAdV4O5dkmSk28clK08JEYZueqyOCpduyoS
UqGIcUknKCKpEfRLXYCP/W4bosWinG5oaxhxXfcjMpUnshYhD/9csybdAEeFQrqb
LzFmCYhRJnhoLYEx9N/T86SNhuAg+hrPULybRdwbYOD+sbdGAJ/66gUcIp+jx+8/
PEyqYjfAwZQ9xSelSCFAHjcX9zmKb/879RmoyjY/lvelV298PuaKVn29jpLIZduO
yqJatBc0K5EoRg+S621Snjpl3XJ/O+qihv0BGjOl1QEbXKmO9IhVnpEHMYy7sOvU
V+Bqcdy8iDjUhfPooS5KMG8AffgesxpP60bXZNGira7bnV8Z/KFumcWYjEzvlaNN
8R6s1ilrOpFUz0rnG9eJQDwFyyNoYajJHGqF2YkdL2uYzLwv2KdoOPf4T/f0Si51
fkW4NTVBnSEAa2qidkJeNMDJwBCWoZhyWgbNHx9o0o2SZHHk/ecpCfW9JlU229gp
Swcnqsl5v15zUHGscSG8QbgEmHkOzSW7qBEusX+x75U37etUsmxmpk4K/UnWKBg5
i3LCFerLUQM2HBpfxA0BKR3wpRh6wSzS50X1s6SMAjXwqIt2kwQ/prdeCoOgK/I0
eWZibbvtNFciml+50q9qw0Ly8Bfu/BMdilcO3IUHyY8RWbNPIJ7MIk73KOd3VJpb
c9TY1fJ2Ak2E20CffcHRZSqFR0/JHfpL/DE/ELMITH3cVOU5DnYklVha3B/xPEf8
FGTC9m2NLGhi+KUy8B1/UEZh19ha/tDd4tRH2ZTDxDoBOaUYvnNrSrhbPeencqev
f6yM/34B3heYMcWuf6lYI9oSSsOBvfuyizvyhDmjNexlB3X1yxpLGW/9AzwiX9ip
FaaWAy4dimBtEPLBqNR4cc4dC2WM8AMU0Rtt5YUO1zQ6D4/GzCiAVn0daeixrCJE
9wnr/uyytXN72b8bthxRac5U4IjJWsC8TkTANZn81nd3i2lncIXLRjl3oqw0HbPy
FVPk/qGyfxvyUo7zzYortYo37u6SHvIu/zhF+UBSLH0+nx/09z8CM85xwB1LAZlP
q46YQ8Yoh2KMBaKNa7OEDT5u7fvkynv5P0MzGJy0ciQd8ASKgpOViT8r0daMP+CZ
cGnGKyXBXJwzB6pMJCKodpXDFGTpaCy0OAJOzJ9PlAFk38hyYNY7RQkGEcuqE/IR
Sx+PxKXQZKq64pfW7tWBW77WOkUi2DtFiT+LAUr0wbJpXEjmH0cY5ClniAM6jjd5
YlLJqttDieKQxHfX3PP+qxZmAk7drI3CTz/V7nwcAuZo5iLEkIOPQwnjht7SAnvu
7sJ4EJtTlNlANp1JZOQsURZ/avQiONcv9ww4364okfcbQ9uYYyBvMnOGcvuX+9n3
D5Y6nLIq15D/GMaz2l/PMlxICkcr/mo1GV33XXLo0qay8gjvVMpclHxEgJTAz8/u
Wq2gG77FabVcnwP/g/6DQ5IuVJoY+l+xRKJTB0Y/njzwzU8SayA/7coZTC27T4wd
+aNm86OSHw+IdRx0/azUPkx3MlHr4RSJzV1qsp+r5a6Vm35/PCO/4JY6vdIHVw/K
7VUAf2RG2XTaTSU0YEkLVlg/9A/trcu+jqByhkvVvYWiV9TT+W1Dnyyaay0hJorh
oi0UMXaPD3579E5M3rMUFfm0nAp2PaLjXQoaKPzpCUaDlTCKYgiDBUNQAxm0HZzj
bKUJYfph690CqrDoUj3bhorDPfhBWPRGM5nNsjkjNNs+L+P6Khwj5j8MlmaGitu1
Whp8w1elFzulYOAEr8f+Na4TWn3vqde/zNvCQhwjnxBgtlifexb2A5i/YhWfnQ1q
dDFLPM2akkzh7X8ZDD5xslp4qR/GPT3VL6obyFQjlXLyWxkwPPqNx1jlAi9j/t8C
uaXWO7KO+Y/XIX9BhPASVWOf9tlwe7nsCRqGIyyo7OZUgJMW644R29eo40qARJ74
SptywiAPbMzQNyoYuaIdmYq4s5ANhPtR//sbcEd3/X05x0lojxXnuUYga+xw4uX4
1WIra4z5Qr85lKdBkf7ILbMdwIEtYRnqKZDHuiLsi9sJay1iRFoszoRSpRLPBGYA
Xene652JDM07niCGZL02Vcw6bwdPzXrvf62vnbGxTVJBgOCT6VYBGtBUYG63CAsw
H+ZVX3MjrGdHPVO12MsCY0p9vir/Eoxq3/nL7Rw5rbQgvirEYzdf366Lvn/uX13y
ubBDIAKQ8+ZI1GTNO90sVP6LIeFFFDXCl2F6q20JXu7IBRsAkFZzIEAdOQL5kfuG
8/WQ2M+Gxg2bvx4WW6hda6PrSeZUmAB0ebPQn0/JK40MQwLlSLHSAVmtKDKo1sGO
RK0nsedA9cCtFL1TSucyos1gbzhiDDGTXBemE3Ub/lxEw8lEyzMlxzgYe5eYVh70
7A5dR0u+9iZPmgBplbuiMpjBmJcJDS3uIVYNxzh7BXU7PAallStdWdFKznQfpFPn
0DIiSE+Frivw6gAyb15nDYfk0x8ah1idiObxcqlu3PjXecOKGYagezHWey9WF2Cm
z89SwLACsbZos5ui6ILoUXlK3rr5Fvr0qUNeI5sGKn35LhfpHxmTpqvXaHepxZye
lJnL7CBEXNmeZrMvwKCFIy5AjCnJhDBt7D50FKUGTRCAqdt0O5l4X/5D7HbMcNed
pYHs0bOqtr/VlL5Oc/wpldZ7FpW/AU4xKHZSAynh9cTSMcNe/LUI0XBKdqvXuqlj
c+giGYdAn561AGVlHS0lNG3bC6+YkiTwBZVWPYvdMaRFba072dHyuiN+r8kQ/Nhj
lxtEmAYTtmjeCLpI2aQCejyB/gWp+Bwwhe58RmBmuZFfj9gOTnpB+63HkmMdHWpk
7AUINfGdp1vMuSI03/1owuUiApXIznvSi+puOQI6jfppti/UEGGw8Qc0ItO6OL3E
LZi3NQB5YphJDPUXVIxixofuW2Yt7GGY8LQcIQIGOXRV3n14V0tWaJzNGKcScZ7M
JdA8RbN4a3C7i9nZuTTftVxn6HikKakDwvc8E7mSGEkLq6X6Tc0PfyDH7eBKnMtt
oUNPqhrgd2TEtSWKFKgyWfauBbOrOMaaZjsivWsfG3O7HW63KPISv+AhC/3FsPsJ
FbJeegiVAX7v2nZitjF0RcXCSHYWrNcgTyRFlGYq4WODfAHXmppNlv5qsOL0v0Mg
BkoBGcaFpQgHKNLhxQvDhH5Quu6Ib9G14IpC5wuTGjMEFLxKmqZFHS7ro2GbbuFm
uGhMOuzKuGx5Ul7lRSv5VRirBzc9WMjX3p5/Y4hrzVN5MQSDLzvfXOC7GVwPeoyf
suzciiEszfCeWkklpCLPAB8Zx+o9dyqeH1I/SIy6C+dx9r+17JQGn3xXA8k33QeR
/OyYs7zs5+a1dI83sDRd1Bxf/uGHtPUn/V2X45EndLiEZKj3Rvr6Iq5LDCMaGuxD
CNdu6i4baKwcdxMTKn06uy+rO0tzy4C3GEBvLczRu/BkyokqNO0AOVXJ6k+vhhp8
heyk33iCz9ACpMXVyFo6B4V5sY9xVoYjB9uT2zCn3L5UtNc4fJQBJAWMN6WBRy/+
pTZqvw+60ZUZK7Vulr8Lx1rLt81y4YARRhUHwDZrOge1sG0XU006qDs2vUS7QLah
lvWoyvJV3WnNPjdHBns8seAFgnvbWjnTVxXcMrXtjwFFxpd2PpJTjPiBAqWRsdtX
Trp6vDoMh91dBbNFVX0v3prIEHGn52eC/OfWRfMnnLUR5A2hKrmLFl7dz6k+Hybh
oTPVCRwEMTCJxv3v6Gnxo4WKI9r17p1eDau44Cnk3sTE/r0PZDZ8y9bSmUiCbxZv
+en19ps/HfjYJwGpitWu1MuZMLPS+m56MAtJS0vQt9vEGdotRBfdyoR5UvMwr2Jg
Me71OPylWVtpTBRE2s4JI8W8u2lhzAAFvFiCHWY/Lm03VVjJMN5D/dV++C5WTWgv
mqCTsApC3ceq/d9IYmnFvpZSjQVEMmNRG1XNnj/iUaPVBbF8316Svd51fN1ImMma
aY/zM5Y9x8anJyLQb6K92yXZr0sWI7twEhcmCf1h0PV5xe1HN3nHC4+iok/0eju+
Nnv1ePEMAnssFNFaw7/WVlCOmP4MKsUYxb9V6qnYgeV4BOywDnNJ4IcC8vvBy4kF
31FCzdWHZra+jcn9rDhjyVJbRUHyV359VP/vzbcXDCo5ohwVlumb42jct/5G5hN0
0eUCpluCvEN0Zp+AZqc1g/glC6wXLZA8BkyRgiKX7pvq1NWAmSXB4zlGndlflxt7
JsBCZTqzGveyXowWeWcLwfZjn1dqrcc4ebKb0erQz+hA3YYbPalkN7PzNDBlEMQS
417ArSx6oucX3y4IQrtwMLegrTWLxz5Dk29nTd9x2Y4yVIH+Af08LdSPBSkmpEtG
064u91UtRRGLIyHipmf/4ufpCXq4XooNIelnW6ojb1cN/wX5hg2/mkbpwCSADPw7
iuFIO0LAV4SXHHaUgXnude0CicFQUIYrGrHnC0jUK5g0UYZUKJHXcmfJtvtMuxfk
E4V7BFaSVdMn+NOrk8FXDVIgS/+5kWm96cLdsMI4qA+pqSDHVUJXaCaiqvioxeDU
fwRiJ71QVxs5lyxfIWcq+VOEaxYrynhnlaS0bJUorETZhD5IpAtLGl0/wPN5D06o
KVJ8Z84TRfsLdqQFrsjmHivnLZnu5p/AjfH+ocoEWyZxwwyUIWnfCLDcbfaXUCyh
hZILpWCj45nf8XafgiNyvwUe81/0E9SdHjFSnU4X2E1qaDRn2cRVO0cn7POG15l4
/7/eAtX8BzOchcfl95CQmSQD+o+qdrNp+akbdB70uGh1GecSzK0oathIbdtfqB80
jDcmRUlmy3zrkS2c8Jg8bSZAx2qEPdzvq85XD90y7ZuYD+xeEYm2txq0acQwSU4e
MitmZhyYI7HeOqOOUo2KjfhSO2FJEJIEbnlMs+pK7dD6yzYGkNECuFVeon1mrXZ1
L4pNap/0aOuqNpngdD5N6BoTyFgNgghqlkAX4/QPax9sQVEPjlZd3a1m6oLis5vy
9bT95yukEI/U4EvLs4F3QUr76NhBST9GFQ4cPhD+WTcGd1qMnSKH3IxYlZu597uw
tfLZLyY9L1NzkGYStcKuNA/f2adkC8EnI7qsA0AwbfZnqBpYW5x2e/FOITAHFTvT
3UROOZaFL0q+eOsQCrtRSIZnO630hPosXpkkzJenrNvbN9SldyUpJY9lyJBsAlkv
OiOrF/9WCwzc/K5TjXmPIfxr9PJXYiMsxJEQ5tX5coAqCjR3HeY0TK1c9uCAjR71
QfQY5cOy3p48qE2xBeEkULi9vaIwhiXjDK+nn7tZvyZrouWr2PWrOAEL4l2OQpOS
17k4WblunHpuqW/2pb9RHQlhgg/uQtm6DNvLm7LO1lA+4uuO/DwfKxtg1NsDTsln
nLmqYaShutj0J7LZ/iLwECW0asYqiXRQ01t44g8NF1dvABNcbKxhr4h8WqqAbvDk
ld36Eolnr3SzqvQR3itlh5ly+lTFjvvT1rEA1JKr3sG+LNvgtoahQlEE5OY9zsXl
ekT0m9Yye1K3TZGoyL6mkg3XeDTN/B//RiskdMJq5hALvQ8+h8K4DdYEHOuSVttN
OkdKpJVhUbhyMRAJx8paJG/rJ40QltdR89nkHfrNqzQM4hqXIKNiPVsCZjEHXQJ9
MFZAElXhjPUx/lvHpjYGLyJTqc6hsUnNpQwz14602zOtQBp4w9B7+6zeGpyZcHvl
VK2Eqz1PMWfmVd9FsGPvEDvE24+fuzyCFYilts5xtLSSMxCryQrswxS3ccb0Krl6
GYuIqJ0BbUY0qP0ymUEvtou3GA3qOFTuFVmrd1wqeFvOpa0OG6rBEtiH/0PhGapK
+q41064g4cd7WVw3HEMAFbmtgnERHHPJ2bqGxUtZ4coDd/h3fCz/GTV7FLKGWTPB
g4AXveo5gtddKWLceK8OPIAK9zF80kk3ESe7YIeqDDHWjCkZ4oyVRhQVA7FWhIb9
rg3Cm4u5APDyYAIw6ElfQh5rccqsgqrsvQPIJq0Ot1TJ0Zd2k91l6JuDZs5xjtsk
427kynWC+v84rAcwR/iq9fmsKO2146+Afm/Zm4r3HaVCgyINb6qZMrAdScUuv0RB
8aDSiDG71DqLDPXF6X9i/hXLnFcLLvZplJ2MCSGWrPuiovYV6MTrF5KVbkj12iFV
RYAYbIsl69v9aRlSdq+xXApRfFMb+AyNSkOftvvsx5r8l9E5TU5/8R+I2e4ngtGp
f2W91bqhyAsXAfHzF9R5zWvPfaHIpOgKnFdpR2btikxuRbIlvkID9dZpbVEg8F4W
oPynR8dchk6UViGL5gcCQRMTdW6qi+a7870QnDE604aQM97MCaGw7YSymmEY3O68
+fpPlockG+fVDM3xTEPV3OWSoZhNAWEfdfTpLiPCK5l/KTLlNGUmTFp5l1EnN3oW
lL5JeaaFQmYVnykRDE+PxtmiMZUvr2ZmtO3JCOCFsTZ4mBdB27w4WEBkyxPOw/ca
003l6p8LPPIc6XD7fbKaNUNZJNhtFz8AvH4mx3Wv8+1CrxMbZx4Tyy+ONnXt6I/F
qpld3EStxv2R6zBnkY5s0iKj4keUAhAQ4AbuMxk5TealrUaMMaLNLLlFFndOc2Oc
GwhgNn9/xItOlhMMOTG3CPWrvGp6sIheSEKuvfLLnGm7e3uo0Dtieu5yTnhtuw6F
ZrYV8p2J/rYu/PyGTtrgpK0QpJOq+sOKKri1sdP7/uehI8txdW8m9+j4bQpZRKK9
bFc5qFoXccCgPdNYqTzA55t+HzkyIKY5USrUBYSku+88hPQLsuKK2o87sHvxExNA
CGlb4b7yKgBcvah1JWovAz5bWDpSXQv1ZDZ31b8TvmnK0wqAtx6hsams6+WrL8AP
uIBMtpm7ZiJChO6BuPpvtBtFAwySQJ0S4yRXVU3mCgCQObfRL/nA0l251RJw+HD+
gE+PKBpFwp3AG9I6hPJLLjTlMHGLSLXPtRUHGhqRuva3N9dD1pz77I0yJ3LKgI/M
MzXcmvAx28vSZTAuXGQmVGbV1VPRTuFEnWyxhdsJOcY2+vRA1bpRJwrCMuUH+3gS
2PUJgTTBFQiVqFtaVwGD+SJq8l8hquyl+cTJImKnBJC3f55Atp9IcfKJyKTfpfvX
B3M7nXdkSfIi/QFgtOrEKHhs6jsGjCrpPyMOC+0qM/VcEkiwM7Tfe5dyd+iWA/bC
77BF5e/hJQu6ymKYoLo3f3HUZkf7ozctQdaKuddiXdGGI3U77aUN5AozoK4ZuBNn
NkJoTk8KKvoU05QV/6RpGRggXrPOF7gi/pI1IOJxBEWjDjVT6XOAT+wSfZu6ZVRB
9cYHhxeeFboxsNT25m2Oh4S7vfBMB7TWX6rG10N93AM1A/jSOeiqMmghrlIs8/pG
3/4VRi35tX9t+Jka+FWAUIP47M5cREkadIJ6naWngRzjDt0nAtxsr4ecMaR4fGEq
yH3tw4CnWfp4P8GG+Rmfw0dIAZPrY5UxHJL2i459D418LWRC/1TJJCtUK5AQjzFs
hEe5zJu1mXXROPNId8cpNTlp5uxHBO9uSwz6KUlfRAHDt/04/4ydsuqVwnx9MVGl
413+KKH/C7Dr+fzpuowuN6Ja+lM1GI9BugMTshqYBj0xrZQ4MXMiNVZwrOgi0I1w
pEAdk0r8OjzyLJhg/zDlA2V55KVa4pcbR0+vK1hIrjtUrGDMFiMckkr4NwpOD1s7
gDhXQumWi8OwReh7lXOMK1WTepukR39gucXNoKB1xZ9v2uUruYTSZtiFYKc73nQr
qhsmACwl2IjZxTE8I10kRgz8E43+vD5KE0/iFH5Rjtvc75HzGiZUvd/nT2rl1EfV
+x3bza8+4Z2+T3eItuw5ppAg1darbtXwVwdWcIbn3HM6mL6f9DuJyOWGaoShHCCa
KOhApRDTtBfjq8jkGrBQI18LOVd/pkPTm6JsKhTiotS+/iCEssi+4h8X5BkSBQL+
WbwgkXAsvkZcKQjlEmQcM6z9tuxVFEtdo7ifN/jp0wF92hpoVF8EML27T/GXVjdJ
UgHEd9r0+XJBzJo14kiso/VGejgFiK1mwemfuKvbyx3aTnyjCjOYGp+/P83TiXQW
NLIX5ydiw5g6si7+nSg7VbPlRFbZ3uxVyi9eR5VK0OauFd3ZU5PMIRBYF41ul4DV
qigEklRQ6cvonyfldpw9FJ31wcbPXsVA5XzhbIFQxqhDxK+DQKIc0I6Ty9ERmf4W
S4P7zDOuSy+42z7rVmKkIOKVeq/WOmrbEFRR05j6tG60r6RXlz077EMsBaxIQkpd
7EH1Mptdg8LJlDM3aSt7zPY9HJ7EXRtu6aCKxsq1XEZ8XdIby/mzypAioD7YO5K2
TZKnMBz4nztHKGlS3XJt15/ASXh4GECqrdfEx7WRyLaWAc6yNTn9QLUTQ9CPnANh
BDlWqC5z2bFLK0PKPCk0uZAuLcXXyYBOXCU9Du1F/ctkKsuw0hdATiCSriIxBTOe
QmsPi77Z2xpgp3aRUadbN9O/FYikc6bnBBcK3r2dT5m3JTAbo/0pxidt6pUMUowy
Qbd1t/nk/E9+rily238OQEL5t4zGAnqpCDvSHoQG4xMSEPlau3ZHUZXZR21K5ItW
6oSiQjpkyRT24zes8ecRojxcP5lY0QnebKvudiLMQcrYdLH2vEXNQ2Gs6b5DPqVW
z4m/6kDWnASdbShkd2BtGQZHC+eKPKfTkbcbNeDA3AMfhcNQhRoVjwd5FVOzzs6d
ZJqPzfeQmnfBZotBhIC6d5s2sJJYvF0fh5E6iFycGC9P3+IwpNx47NP3ujm1IfsJ
6nJpR/Ynz0cmYXTBHUkE8xRBzolWsLmafhjV48YUPN6CAka9U+o2TUyrR4uaVAeG
CXEf7C/c3412AEdI15AkQoV8wkAYLSYx5qf9xbdqQKGpU58SDdO2CISxp8Iqg72B
YhS+g7l68puidsUtGCXTVT2nZV1CeNhJxCF5U7H/KwOeyeCpwUf73dLDshr2Kaka
/Tn6WU4us4/4B3lbZANOUcEelMuA3LsTRv9mHFF4G6vHrbFgGUzYjCzO3yXLGQGE
tvrb/Aer+BtUuPi2y11TrEetgn3bNyVl474vXa7h+JW3nSg2NiUiyECkYA2TLoTV
6arN5rL7FeB8IWp91mXeZfwy01qcoORhXnNyB2tQILrFpnaY1EA/qcBKiRghNWkk
BuRYsmU8fsFecpNAC1A/y6v5QzDvjffkl2+cxgC6VKpUHFOUMGOi8rTE9S3PjkrK
baf6xkboywdLsDHQtpxpm3+QEHBUehLhL5DKWVNGooUc3MQqrHQEOkTEQ00BlooI
zUIShCyUfGjS2RgBPmxmHuZIYOeiGbfOpfVb3p2jkMVibC0IphqRQqCbGblmkKxb
K/PZlkfDCjXmhUwrX0JquZx8LfmsNF0QfN5DIEDkKNEBY7aSnNhtJgG+vQblNqgk
6x4Y9PMDTIflllftwO1JtNY6VW9QERapY/6MxFqtEi5QzpHBdiCUwzNBEtm59322
iRwIeFDE/fhkE3RIWGV2TxuFXj0BVej+tTyCTiKfzKXvWrBaInVCd2EUTA1INnEQ
wy4Cp5kiQeJ/XBeW0GxKyyJau2D50vDBXFbAWb7yUl1ybpsG0Jh8M2geExCUksOD
JW5FiPmAiqmib53CQ52XrLnTQCXfrpfxRMVt3JRmQ7c5UNRvhsQzkmAC6ns6jNmX
/Ua1qLYr8TTWMOB1yNwsRCxgyccNcaUCRPDKGcfFFJFaUSD1PzyCTVtYfJZhtMF2
Ya2ppz9jIlLXQ7MmtFPm9FlSIsbVHJrozTpxQv5VDNNbTRjJMwE5Y6y0uNMZiRX+
vl0tafpGfm8LyjywB/FPL3qMMKcKgCgqqrWOqv9NIxWLZ2xISSIb22Gu95tYOIi6
BowGFXm5BhpMD0VDAH5adlyOkUQYWJ5T/VYRe+5I6skB8uORG7TWBU7SlsStlsH/
o6FFxyNpk3V4tFmAGUk9euZ2tlq6l08ZYF5d0Iv8QckU27F5XKtXu1GqRRfBGTtH
p6t/fe1ZiBqzHUQolcdxgBFVcl3DUMgnP/huMyO2zFlUxcKYv/LYl+b6RlLHaiDE
ecijqShoSkBv5Lgdjc2VbDH/OAvOh0dNqql3fon8lqXAHxB2KzMc6glWjGNH3jJ7
W+c5CJTGIiHagU6NNL1e+docEggGWnSWaugMbCFzz2CF5hcwHveFpK5hKLxyi23H
PN1k5hYo63mosZXWXpvrADtBPghLuBezNKiiCqmsCQbzZbhIWc82PXN/j/DWQHZD
OE75eArNk3R2iefBy4Mzu4/Q9iXZ5JIEZklh50TeDJgeLI8yTaK0oGlI6iuMBCzx
KAAJvScqFzyiaz+gXW3kbGi5gvlObj7ywpy4X/hJQ8ILcE61cXe98af3M9fc/H/M
dKT8O1BdfzeGcW61TCTBQ0ZHO+hzChwkK61Y/WoYtAONOBNUnRElH/Ush4HXShcv
Q8AdiRBjYCLxLNWJ2O1eVDlMB4IvCu6wWNwnxV4g+wQDw4ehDIW47Dgm86KRLg/W
L09A8MbpQP+T1HncK3KgsbACC/S2PEfO16DgK4as4nUAUMQkAvu6PlXJkhwwinTE
P6c912R/QKZtbyPOtN4pZbD3a961VEtBp5MGWUadr8nbhW7W8qd95aW9hnsG8jZx
ycjcGz2Q6He+sO3uzfLHinfKusduZz/qtF7TVJ/5+nwl7LBSJvln4CnglEpRJsOt
EVbnc3tvvaUfhz14zFT++FfmcNMqWcPU1pp3Rsrtx6PDPRn5SVPiKx7BwelhnV+z
F2rUp7zy+8eqTqmFfF2FIh305TD+YRKnPhVQXpe5Jg8cZozHQF+oXoB74vnBsxq/
kv5YIkveg3+oHyl9/cM6MmyEttIOiVTHXO+7//dBfC4Jy8ICP28FGlX63UNUd+Xg
Yjdm2iyRj+ksUnplie82g84Ii/JhGNsBZtgx5RjCh3P53hVdHlUvI2srf6BLavZ4
OeandFKaJ+rU3CGkIdxStLqxlR5pPfEWC7jj9b8rRuc/gIlqB2F42XNquvIXb4DD
cv/Km6gXd9FbERCQMFBNqAtYjugO2kgPWG04jqBP7G16sLl66SPaQv8tlL1SwapI
C7a5dO6gns9hIZEvgPSaq5Lpe1mCa8USpQE8QDmomdjwGYXEGy2CK0bbMYZQPIBX
VS/uRYBa/Nc+Zm7iMkAjLz4fVLr26MgssMuTcoTv/zxGTSw3+DIjOtYmWeAjPaEP
dp/8dQEkJwCWmESpcNMw2dL5lElwzGEeBXvS+T9gxPMr7rXkEd3nCTJYitsS2tOY
9WIE031lo45HTRyRVNzKh9H2WxsDYSyS+jELdwNoOYberg66s1qHM78SxumQGCxZ
bMLgshFk663dbemUoRgUUvi3/VHW9KjCxMy/kw3Iq7SaggiDMMwfuF5xKOMzORQ4
0kqrrBP2PAwlYgJB0xBQT4hmfR2bMY/EoDvw2ZvcRB1k5RHcNjvOfE0G3F/8/ISC
BMQZPskNX8uCHBuVCqa6yUcvuFAryoIj2GeJokgjuQ4iSKSe79tOuEttQ7Km3tTe
guNpQrln3H3QDMxaMgmsIibGyhywFSV8SNzJ+pFj1euYQy0feE9Z2SkU64YgxV50
EfyLZWIm9td4qieQQs3GzL9PlskYzCaC1FTlYWbcuSNOBcAVW9wI6kkWEKSZVRci
bsDprHSryTFVPHWIcsUiIxUgieIdBnHJAF7ndbcnFK2jwk1qJrx19BJn4ip8R5Ha
NqVpLoGcGha3+Uk3sPOUXc1FlsAvy3L/9jZz76SnFmOWf7CNtrEG98fnzb4Urck7
ygJcUpcgKcSOgOm8NMJEk0/RKFAGuqU9fjAzvu0qsjOuur2GuhHrpBLtaoJ1dbzT
F7UKQ7NDGK3GxKhd4D77on7LT0stzRTiIWWvS+5lM1+syR67uzzCmVWtn8Ivm17n
LF/5qqxM18NV86UrFXM8qpMtvWiA/ee1iF2aSzfDNZdoSwbQcSnljYUD1955+1ha
P/x9wE+hvmelQnoNVsDVLuUivjrrBT7glxkM8wrDdm0KyR4zHq5gl618LrOrmre7
ne2vEeqPAvsnqk68vyTywFer8rGiolJC1FrjUibDmoDk0ErN4Z8jBt6/spDPpXBF
Nhr/lKsPc7D5CGIuLGJ7eOu61Qw3YIpnX/a4J/eQB+aNHyALTHi/PE4O30DppTx5
UbWt9JPQoGau8lSh4x3PonVmLIlLEEEbILLkuE0mWPSInFR+A+Ug1vQPtlhzgOTs
nCVbMULHbHBFIjjliwwkCGvcG5LthL1CvNhLaS6jdmNsnYw1RPLw0petsvQu/8do
UKfCH9WjW6JGKxkf2geYuj8snLcocWkoi5pmLUX29nGz3D0nlTjdTdJE9P5dYewx
l6eBb2VEakQdYBJEkmtkqh4Jim3R5sKkSuA3lkmAqjb+q9vAkATHkPqbS2tB+rTV
KkueJG3n9Uoy1Os5pZaQoNW+++hPDOH+2zhW2Sd1oZV11JfibpGwm3AO7Bdc7inz
VEv8cMUcE7JrBi0xZ0Qr8fKyPHjuKf8NCyOqmAEkpnB7dyAu9frc5T37yfPMixw+
/DiYcoG+4MoIbYOpGHPxGuJ4/uzWH1KzDzGS6qwYMEfzCT3vehpHY0yFqB6uCu6R
4Xa6vQP17bGGWDVpa4HAy156n1ZDSlvVpQ0iVVahWANaT43X1qngusamFUeH/rpz
bbAr9bN81EfuPmYfrZamnnluzokSSv/syDeXwjFvGp3lf27a1Um1Dr9wvITBD06n
gq8FOLeW+jw2dEJPpzVGV2QUL6QqoiD47vHcjXTjbqz2KVHFO/LEBgc/SZ8XOa9G
ZhsfPxx393PFwoWPmlOKPDf2dyRtDvT4kczQD28Za2Gn6xeJxsx6AcOC5CM2CJQc
RlPXjg+0I4NG7C6KUyZLv8Gn/uCFTdcdejHQrvtZacj7l1+YWT+G7jRoQRYQLrz/
VPIxXQeQIhZxYWIWdOga3Ky3PzOuqsCD6KsQtX/EWn8/8XZ542XTI13qNRTDq9iS
GGj9ZOfC6LwT9vUlM6JIYGvZonIK9H2Zj6hxRtwhsEOnJorUrXShzdHjLtIVFckx
iAiaNhyUoFGIqUtQH3P14y5nBdzwz4DA7TdC4sg2mkqc2GRtbSqdkVkPn1H3Fuox
fdwVKJJrbLbpfhCge0f2mD53Cdjq1/TZzJ8l9a6VeXzcOus3/SgGzmH3hG3TddPm
EnFXlv1xclSz5pdQKhtwesz6utL5iStaqpYsPCenLX0l7A7jc58jRPMxCLSDRkXc
WFb+w3VlLR97/xhup2Pfyy0+E+ZmdSI6GzluIGhbhx5SArFnUaWqH607S+4sM1JW
tAdX4pGH0kM7RCUPESmrgzovs4O2QlwLMH0+P6NVGSRHPcmyliPa1eW6HpsZiWXp
jQ5npv98ONtiOVy05N0YnM1mZgVncGV9hvHRYohbblfF3GhTZQ7aA0CfmPH6f0SB
powyXD4kYxvh8Uvmw8vPnq45PTsuTaCmOl1Rlcsy5OW+lSPy9KiTnxSo4whlHtwr
pY7/Ho7s5gbKlLzRLTx86alVcquDxSstPoFsCipjcb0MPJ/OT5dWXNMpPFdoJ6Xj
TlAr06Vpryc3DNf0npppCup6VEdKju0owJBf5dgI+vsvg63dItkRuZ48wvPef9Qq
ABR9a3uwP5+GXQwXED09KRzfjCb5rg/Tew24ve3O59QBu8dZ8Rk2FhyNmaHcjs85
NCmf1FotABhNhmZxsOba9WvzdkFZXwfiJNB3HbWZZATumGwD3tAuP3o9JV0cLtVX
aoj2AqUgtVONb3i0eeU3ajmF7d3uvA4iOFXbj9hq91EJ5fAzZ6CEkA81YF6EzGLC
ZkgH9zMahxhm1/EYgSrVvL+bxs2T+UrmXNcfglrWIt1HFKxqDvSd2HiGrBIESwKL
wnxBUh5+ACoQEgLHDOkKjDkU/znYKcMYcnn0T9kyaitqOrMFUB96BZDGMzZ+GhaC
fOTE2Rt+3X/ma5NdB1FAJxUhZF1jYQ+2+tD1utZWm3yYZbhhQnCWAnBmw1XZ2XyV
CAzP+TDcUyckIv+Y7PO5o67npmZ/4N8U86eRB53Jpqou64neBP1/g4xc4RNDoW13
QKvfmIsnbgveQEylwF8swg9Lv69wBtpxJj5/wfnjveaoUy3BZ41BrFyqRCX1iVQc
Dimdps6VkjQFLuzL5E22Oq1VNW2FhRFKrhJMmYkpTJ1qExfTZlAN9ql1qrR6qNDt
rh9ZpklgGYTBgjb3XTeTvNb0j2+Kd8rObevd+bojcrEboHWwQTxySAVvxe7udFIY
QNEsr513NOgzcRnAghJiXcPRtjYx+2H2iMy3B29/YeYBLKojRxB8EW8WkbeGgKph
pb1UV80T4Msempgt2pm0ZOM+HGlFu8r5QJW4O3kwrixfQJJKWtse16ssfQNpih1Z
MtbXwcl4IW+kB+ONuqdgtoqpMysyfazV9yxgG3z01v8OtXhbXjOJD/NBSSBnpE7a
J7avUnYdL6UXcDuhZIQXkScnxuZrCUO7Qh+vLpQa5iHmBARB6wDiTHQO/dQALTo+
Kj5D5dHmea8nc/6cB00JohNPz3/P9iInlHuC/AfTPP2n06oOvDf/syF68Ord4uzL
+/aUgkW1ieBmUQzA8gT2GBMqPkEvgU9npszTCzV9fX0KofiLxIX0KsAQ76wIVAYR
VEVEJJrP5ZHzD3OoL6VYDma6of8aeXOwJDdkXv6ojDfV5P4diUuhOhfDhxkc75IW
qM9KNajtLEk+rCUhg8WT9w8HLKCDMtVAdYjBD9clShv9cIlyPinjpqj43K3yPvs4
j/2kTCJm91gnVL2DZ2Fuc6KX+ABvW83ZiaKnEam0Wdc5Rbzpq2Zmx/QNM1FijlvG
K556Nx3JVuqnKNimZxhhbSutKPaIbbQXK04ZswfFHEwONicV1FfR9vQWxN7FVXY0
BZCy71q7CgRKJGVacj42Tb9pGwJz/NEdSjJRNJ84AwropfDzNSXwKC/dqRP8snbG
s6bZyce+qlSVxPkVLk3xoLBUaSqS12C5aASjoSNpI5NSOMJWMhGgPr71yvScVwYv
oyvMjWIeJy8MI/6um9AZIEFv8gxg/9eOWzwFL1GyXms+DX4ZS5aGw7PaijGPVU2c
1xndIDs9YCBXB1rSuBzTlhA0n/loCoXXcvxO6qUS2tv4GXriTmhugeDkcXXiRY1S
PXU8PG2lzKrtkLHkGrLB31CXKBEi2V89GjdPnidclaJDHgDhyA1aroVzpRIcDHdU
h7R4hSe0rY/Y77vhFt3tpOMIn9mcSNmz5IH2bL94xVVSZNFg89VlVjFs2J8ZtTWW
uPBx03TcmVzHjGHqf+WKeGxTa7gxpjWZchkeHRjVXdfAQY66QZgw+5EkPcCPWa5V
QBh398hh5s2N+aUkt08EOTr+I71XoWH0fi1rmES/n5lmMnMjrlzyYJeTDliAcfoa
z/+Z1XrPcDuUMl8Wl4Zt3gN/MBq/YNlPhzDoyPUqkRg12YuAkljcI+/ai2ockxgg
6ob9A+89wjpO681O+Xd9hjRcC2QUJhECrIlJJDa/CcxmtZqE0cNJqEVJXIDa97St
iftzg1oFYV/dYRVyMXPCsRk/pvwTxf0QgGnrFNh+gG78bIz1713rkT32EarVvPvF
df+hsFzLDxiNC5EpOI55ZqJ0BpPklqm3aUihYZav2Etkv+NiPNcA0vlhZQTYflxh
u6GmULEAonOREKaw8n6XxzI7VRq/0aY5VoDs0CElQpWx0D/sjmrzv/EyFQPNUeqP
wh6RNxFQzgi+bmVD1LjKPSpnl03xqbovgh75g/4i9rBU4Tza8BpPuQKTyyMLiC6o
Me8Bdwcr1ZGMkEn5w7o+lPFDwwLnWIA+2kkwqXXmr7tEI0EkQd628V3cpoXZ1kJD
u/iaAAOTbNOcTvyuQf1cBCAsgQSxQ5xM+h8iFztgcX4VcifnGtHkz7kaPs+giIbA
WfEbY37e6k5xRdo6MhT8gfRTP5ka1TB32TuexmTkEQtM+6MvyjA4QIuXHmvOcfFo
5ODnYZz4kGsVulELFHKqDSzCg+p5pkrLvPuhYkmIfLENQmrkZM5XEblqVkA4FcsU
7HwxDDy4HzDkbfwLO8n7flV/iu2Qeco4kvF7zH7E7vHnxUnakv9cNSDYLlTJTCE/
p9VIKLwZ8sXb6cRmPOwwGmOlpJbrx3XsKEb+N0eavea1UdYt3PzyySiEKidedfMu
46nCnHoyBMyOb4nJjJ3dyEPeNEUvQ45hvwlLRdTR1MaX9Yn8d1A4zVVQG0IIldQJ
dZyae0tk9S59soKUp4TTSLXRW6ZZvFDvPSunFT1o2C88UoO2Xk1tYGPGP6/7uoHD
Q8Gk8FKQI9bxuBHVvefZC/zJHRHRY/NF1TXfrTgRbAl5S4lvKgLDbKK5wBAnBn6Q
v4f7bmce9+4pbnXT0cF/MtFORPJMbVLs4QlQ68wMIMw4LwsZsgGYA6QsS5fJ+Nac
//+FoDjNIecB7g8x3OlbOIh9++UydEDrT2oRKn4i838R9XXNy+G0GEbMASx9gXFP
V0Oz+DKvTLFpQP9eaj6EKzlfHqKYkAj2CQmOnSsrJphIB7vR3+7+6QRI/IOOHef7
ODR1gN0xr4DxE/WkinTRZZeqL0VmwGpnym72fhHYxDhLx//uUCEbh7s/AtDfhgeE
gF2kH1WG8/S2S/NZNYomV/LS8FUQl8Zlv6GhbztZQt9FSnF3qGcE1wWHwRdTRWq7
a135fiE7uvaVTs6wQVmizoPhIPYZagRxyzWvQzYZ2GxxqDgKnSJgJdxnbhYURuEX
LT4oXJ1gIDB7hV0ZcG8om6Rn8F9c53IHDaK1ufHo+rLr7b59KeW9MjI8gyWnH6wY
Gu9NzBOstsRmS6hkB/PtdPH0Vny5RO8LLfF2asBvnycGPsc5vEnCw/kl8AwHiJSL
Zw9eexAklEDXGZX9AoujJhgk/svo/2T3ABuUiUshuLS5yeM7wlkwbu7p5wyBrZjv
puN6TtZ3pSJn5SNv2Od/I59EAmjWy/IMA+dK8z2druqLUpygtETaA4FOp5TrSfET
H76wfDokVnO+L6wM4o7ar95Gca+kn5MARTTLQ5iyeBtRnSSW2qx9UtMg7Ziy3O7u
t2gnVwoiDOvOzPHB/G74DlHIwzPPU0UBX1t+anr3Tx9IqK+JmLdJsuW11UxqgI2v
tzdH+ydZtjVWHZ4FNfGr/tHco7vNVkBX1gSbrV9gjwK09g30Ij4gv5RT5+6GH853
1QrVMfU/+Byibl7FtvUGPn9gRKerMn4a8qFLTnKOXQmmzRKOcwMzxf6AT7Cl6Sf4
7LYvLSpYNwA0dlBnIP4H1QfaY8B/sUsQLZhohqnI+xWkZQUzneGD0jZPYMFL6zWT
VCbNVZEWAcTFvZ0khJmCvLtOCUgFOqq7yIZ3qCCxEe4VhJDnDxqEojSikQw/iIqL
noy1PSxLRoqNzF/dxsPiPkXu1c1+v09kUjnQl+bMf2szV7UDQeTdjHz4S4Tgl7zY
cYxjWb9vmhskG8zT078DiSvO8lFVneCRs+/l1rtzslwSQtxVFUM6qCvtQUu1Rg0x
cyiwl48FoSDi4dvJYDUlmVofdoDJUNBaAKmb9tmd4ADnzkET79dufCDUhGaksxHx
BiyCIkDVCPrpVA9NYKAs7CMWKFHwg5YOaadLmtYuyqYEosIZAno6KapEUuEYAezP
0vS9yYJBnbS5qnwGWNG8kun4BSdota3AyKpJNwefWGl2pwcvnm6qilYAUvk6+/vt
EpCaYMMHtWIJE5V1Pq7bi2U8ZS+P56p1yLtf5Z9JHpAvND07S+53/59gjwfMV5fB
yY2AEBp2eeFEsC3Ku75PxCVFxXScVFsMjt+DbiCZInsytuzYwdEpGSUvuSwevJs2
P+MzLXQhm0USvchTMOMQY+BcvIaB2udhW/RVyZy2N/zJwRlX04Phw5vwrAwudT7j
PxtajcEmmgwdMFEHtdj4LbtbB1HtPu0fTOk5gFx+PJ6XNAJ+zEcxtchJdhqgJx8M
k3MQMQ+1KMndgcAgyib+eio6PzLayO1izNZZTJmoaishoM/VIHUJ4vCqioRH59lv
rHdidrMiTO4GUBbpp+mMuRLlzmjp9AzmKtg2Ped5uv162pMQtZvZiVTEr7YhHunq
2WyIK/KCrYEwUq6QkpyDBchG6d1qIHawTKa19aNeQTTGBrUqXwZRvYDGGH7N9yrL
cSeJMOTtPP1KeBL0F9782b9GmEmJAQZBiQMPMMIJlIxVLSiR7r5HyQph9d9RtnZ9
5EH4Gikv/Eg9toL6Suaq3trxyRw0aOvevyLVfCVECqMrEavZHVRa7/ZH0+dO2vMb
0pe3PwC0XyMHy8DKLKYmD5VocT5VEmv9Tt9eFavglTn49/aYOsK6IEAZZajdHg8J
/gX9NrkncGPi/bU5BZYIyfvni8zVddVblz5yiPJf4fpQ5tXO3lTDx84JlKdpaEbm
C4Txkm0D9CZy27EycFvPw1ePg1jdqlYmC5FcabpA0hzYuW11bk2q2T4cZ7OB3gLK
3I3qJ0OjUT3N6xURRmWj/c2zaeKISXgovzXn5VM9oDX2LL8sRBLeekmdvVFNAaWy
yMm3PtIZLmMOZm5+mWiVez4fJODDDrC99YRldUvtqwSqxMmxvx4mvCpqdn2ESoR1
EOS2vMJIk7dzmH64+QzL/O2NeGwwvlJk4zM27pCLuDn7NeOVS6jnFLIA+6CuqRcV
XxhEGbhb4s5aLWrTHu+ipKZFzTNNMv83B9g55M9EWFv42UK4tiggxtrQkCE3MgQi
uG1HlYzpBkCL4Wnc0ZiFIqdNr758gBhE3wRMN+nyrbNyilpVkIRiYtKsFLA9BAXO
rg5wp27K5IpwWl46UeJO8jX6NCmXlsbPGTltBCe0FTAsdDZwZBrTjzcv42oRuAAi
6Jfjucjc5BBQXvR+Wzwt8EB/FkyqIaqBWhhkbC0LE7TYhA0R/badF4FV4n0o/uIa
TX8huFAtrYZGzeWto5pKewrbOUDesbs1fCyaUtw7YRTO3eRMalYpBXNykc8DAdqF
bJGwETj36bVN30lTQeLpkXQaCg+K+JrVy7tB3phSOcQfIAUFgdYgLDn3Dz+lR0tH
SzsEIlZCjAf4+LU2yIj5IDLQ2JiQLygqEktXCSDrOMtIE6KWhAgUuTUycBKYG4Yh
Xz+uL+EiYjoTWtd1d+HF7ZpcW3qtQV5qeFNszljy8PAhmRlLQmGG6zkcj2GeeRXC
gtnwDYdGQ9J+59jR7DRMFRF6ObaGgmzyRVep9I9rTInQ0tld0u5WL7p4U4ay42pE
UVqVQdL/+N2ucZS8NrF1W9YMoKMc3pzIdg2/m/Xg6RFnbWkl+ocVmG8L48V7tgDk
a9EmLihI6LTS9ymFitkFRyHoUGxjZ8FR0JcOWNiAi8+GYKgaWyRLUH5bwgO8lCpw
zN3q5Ehi2OjcxcDaDobQyZBrkIoVjP7iJE+zuVx/NCDRj2uHxHVdGubzIv6lLNmT
oDY2dhZ5S3bDmrTVZokyeNprjihbdDgrqb142qmPZnKH8zdgS3ajsJSs5kdeqvWi
dH8TBaNF19fiCDkoWrCadLUtg6PHTqlOGOo14x3DZ95A0uq+fWi8jbvfl3WFmsvz
lPnwYnoWVLm96rLXr+Mfqee6LzM3H32GpdxYZK7+x/uwA5uVLfetDdOzWbdwsekU
CNNaZx9+3ygAvie3WonpRcjAgpSiyKMgnT/rxTFoY6hifQhqyNJrsRQJH20oYvP3
0G0ghUPh5RxI9Pwn5U9ovpvqPKQm5lonqWAx3nSjnroHjC/eUezd5t60ZsRIbSq3
eKLUPQa2dqAPLgROi4kt9Vvb9amd/jQrvTpNmpvxMg5mF+fU9h+jf2ZFrRYyS8ar
1naIinRJoR+bHznixBCLykdTG/4QMz5xdDeEhfFVb+wAzk1guue8q3fsAE3Vw1pr
4eRpZSqCUttHlN0A2tclyF9AKSLJQAfxUarPPLyvdrub+nXyNWiZ2KTeDVuKud/I
rPgHM9tj064uukwk0pFR5T6ChLl8k/U1tIiFUeX7TF8GDsWVHX/1A4e/E/Cwtoo1
BiQ6f9pPZKyCGPgKSJCzZ+N+B9v//jt3JuanljB12zJdxSlAIK7pVyhnzkdEGDa5
cDJxRYVk+5s7IRUb9JJcLzxb5VrKjqEnwKAu4KsPWg9j/gFR3hmJS9xpJ6ezkhtz
JLac7OevKggfScCE/BdRZD71CZZres6umRQQF9WOy7vespBPEBzS5/AQNsqWvFgi
jbPOKemx2Po2i6iWQ6Y67yIMvbaePIvaeoJvZ0aRO+tWd3dxOiRtyqYpZdG8+hi9
Nf2QybSACGYXFpgduKxKasfsG/ln2ja4s/iC/otF/WQ0lyMplmy293v+3j178lC5
C8vyWgiTwDANjKsP1FrTF0FIKUYezmdlLZcK8VxOw0BsNyDLtswI8FY/t0QgLm44
0FlHVVN4USPo4vxYA75/aEzZ3MucQZNfy9bK1y5uc+mWJqEnqW/C7vjVPCmwg3zf
2esfYp35R+PKptN1HVsUHwGys+YIlmeR/I2P0mZxeRk2nLO7WuztrOlZehzgyAlQ
aVJAiEr0IyIT5eOp9H6O+mEmrLRNHEb0em6BS6F9shEfa+aNwF4LF5IfrReYD7wm
keRXqOSVq0gKmwNI2Oe1wuuY7P5ucPHQwNYw56Ptmd/ZyUn21/LS0NWwCyvWcO46
OFVJ2v0bOz9cZXcM6iFZ2I1hkrahJvOACSvaOEHSa+l+D55JCv4kInWY5awtIA8P
6oWTY525y/EjT0uyMN7llXqrhyVqBiNRYScfObYNFW3ANCa04x7o1UOAK1uva5YK
ucmEFwQFyUubT1RGh4ojJfX9k8da44I7/ZMVKhcksQ7P5WA6znIMGyopF1slvF7+
vf6rGSJqQWMnPHCvXYN1xkmle9FQqdI+iVH1YEpkTjNEk6vDv8HOZHL6xkzyhPqC
0cjpkZ7s7y96eiwzJSUfZtykWXdFoL7ZOFfLkUKxBpsBGe0QM2JQ9ORUb78/Hi3T
ZS8cMrvgts7BhjAzt3iaKjny8/+tFNBO4x1O0bImg2eQ+SJ1mMrjmSB5qUVobmXy
+TY4E4KIDh/DS7NsjF8GtjguDp42e+UMJMyChdPJXsdHnb4ZxWEkdWPLDFyBkKWJ
WOydV7ifUN6mW2YvzlivHiPw1DZ9adCJntoTdiBcsRyJGI3NKYMmpqLmtkVNrctu
8t2agb7LT/LczmyeLPMRKtaDok+byNXHV0ah1F8i7QUkpl3P+0X+7KkUE7lQIxoC
92dbaMC41efkHzFDp+TEhPLdztzdPtMUqqW/rKa7xC1DukxP7Af6zV7REU+sQwYP
6Lf/lpmkHFrcA8SJdLTWNW/Wq46t0CR5pqmMTDJ8ZmSTc4FTD4fJgVFhM0VxgpAf
aAowxVI3ik37Lh17i5rPJCb3NkMIdpK47YRDajY9GuBaS0Rgds9bjs2FRud5CVhu
5bgCLbNoRpsSlkfuW5v2KZrLk9zQyyG06ds+VXIzUyoouxfQr0ZmGfdcweqlqg+/
y8jj2JPIjnosXN9iqu7rRgY8jbljoHBfVwLMdzFxAVYv9gAOn78eb/YhMpZBnBA1
y/utb00L6ZML4a2rRKLGkGNzCdLmRWB86/CiIxBuqO6UJQJVTXuyt7u3KA4wirtK
4sa7MGWg+LnhvqF5sihlz3qpUyiHygvD7zIseklylJGeVVH+DLHuW8pqHO9YKZo4
2L4czkyx1j27TkZQbDHDFwKnIg7c239lnVSJpVIMF5Y+TmqqUxwJdi6Yoe4f09tF
8xpfSul9S3s8ccy9jZfbvqkYwdAJ8I5ryhDxrxU8tL7YhBEDRlK6TNJJ9T2tUf1J
IKdrbpP/PF6GwZ9o8Xo0Lpdbby3eF0HrnHZpUGFShYDR1RX/Qwks39FFo/kNcdwF
FF4m9C8xI4UFJhsp5YDcTHtr5CA5R0LIWPL08dWyCEMJaFz9fhV3836CPqDprk1r
ELy0hirAVvErTToDSVhGj23zCX7NJShYsdVY00fI/G9lzoUKWobdJ3gkNmL2hmL9
2iLKzHYIpTRjhU4q1C9QXpx3cw51q1aYdE8q4Cc01N9RLXVxCA6m+Rgg3N4MZ/pK
j1+gUV7Lo0BT4FRU/5dZKr4XUsQ1O9Pjgd/VpiS0UPYmr0NUeYLLvdQ8HGMoOIsf
NL5U4G3ioSFZa5EBWu6Uf+SD3Fmpu6MRlwKrjW2H5TggGKwvMmsbSqLm0YEQ9MHr
sMJfajoyFgeGh2ckncYUl1pHYJdjaFDoWTXOv6G0N98cXT4R3MhM3SWtd4ak23UN
tapRv5rBkOuCDNquO4lMUTfToBIcVNi1ssc1QGFGnOHQe+tlCxSjmuh3zpQd/lgU
tyZV5E/085Aq7XlpoAmh7GJ6rSI3mxnmKQEW+4M66VzG/l2DMJfNxVDN4DVMqh/k
ILrw1LJP1ios1yVl6kxzAej68ff4BFekFmepWaQvG4EOGZO5aqe69tMzA85anGp+
m+SyjFdcFCRopmWjtYQ/yZbKkVUpTlgqe80YLDZMTFqs28cADGwIafcYfD3x6c1Y
CU5/w/Z47z96IURMDU95z3SXzdfIeIeRR35CaoKW6PMbysx8otLDznamM5UpvwTD
kExnKLDjcpk+n2B8oHSCqpXYO5DUlm+TkWukp+tt3/eydVWqnkdS/BSDv6d88hAv
i69uiLUsX29H9B5pANodB331nnrt3GvTuxSfF/McmbbsrApUfqM6+4JyzTwwqcyX
JcjnAUg0Skf4XuXN7/U1jQD3og+jOpxk5R8o7g4SEONWbrkyx2JTDXIGWfLicg6J
b/YuSIpiWuQvYvHrrdPL3qwJ5kixTQYbM2m3fXhzO5O4890WUw2oENE0930xBOND
cqFthTN8pj9hn1epgn9K2HnPWcjwHt+hRIsl2U3fjdii59q/X604OTLiSaS5j8TR
QeDX8cZH4uYGrYagKlQEiTzQqoWAj6Z1VsgNmmtEWTL3H+2G8pyhXSJC5Xrw9SRC
m7YRwsWrrPL5wUZ1ZctLmKpdZUkqP3oZT/cBxhIVZO2L03Wh1w9CP553Ns3bpVSg
wJW4QdUnV5XfmVDBFcf94PzkksBQRZPOhz0vLRI+mmPs5uHsotTIl00F+S7vHnow
pYl5ffSLQ4BNPTfLuewu07kK9n/695suMDqQx7WullNKYduBAT8W6YXT8N0FFBL9
/ATVgLayB+LxXf6nNsIelI5jN7w5/XunHrTd1G8QVLQpcJgAbGhdOy8fRN/TCmCJ
GA9eZlGEisMHwb6YJrGUGyL3BJWyFZ1T++9VE16HR1QCrAiwghkdJijmZIqYU7M7
XlnUoYB9ahew34uZZX+ADSPiRfFtYcC2T/RvvUGjcuIvsq2qDwjdA84L+Q+iYt6m
zxJ4dOwnt6qDYV7n4tp3Cdn3SXhG9jEVz9FvFp/iTlyMC/m9HOFAIHqPX1eLYahj
O/fvLoCFhiHP/c20iK+jez0T3E3PhLXkZ5h7UsJZbyxFwDdt0ODqzbcx9iIhFHex
9r3Jg5RlrtZ3TkRIvL+JP9Z5xu1x4tqFNO9SVCtERbLEoHM8mMTqjroIGqQ5PE8H
ouFdtDNt028P0ghBT1jldpL8Ay/hKLvfOPeRFsu2n8iGIvOb7tSjubjhYO9LUJGS
Sz8lIAC+ejuX5NynTD/q3ryhL1YfYrGR+5ZHVNuK+U3cOsZlPRB77dvca+tJgSNB
p0L3zeUKNxAQGQmdLCQMZzDKGU0lESuOZtag+zquiVQsthCYcKSf4rtCG1c57TKs
k1pgwjpruJURxq75me+G+HLUJhxl2tWjj5qzeCONr5q7YzcNrJ2bgtxgO0MOxEW/
9BnCgpxHV7h9Vh5GhxVigYNWplm5Ec8ThkbbtaxYDu+REh2u0nMrx1PXqlgZrqgc
Ctv8Yjr5rpd6tUF14JKvflAGGrecj9ZUseUlh3c9pPHoxuNCrIpJzfSIPianblTY
EGwDizHv3rleFEQPeZXQVz7H53NMul5szH+auq+RtWgN13FZ0hgDOaC8bVvQGkbD
pkF+d4A2P/PcwnJncITkNss62ip9dnAT9itHJu7CVEHXAHPgGqElFhoSwPn4aQOj
NyIwHfzow2QC1nSCzygk1seiXLsN3sczcOtEC25GtTIhe/tNsIFNOJtBf9fbLMJp
xadqiosIhSAcMyM4UOF4xv+CQPcMRJXC2k6T9qNRq4zwNeQVINoIyX9KRHajru+D
+uy/0cs74PCSqTdQSTJOv/gaMBtLzCRK0lAOM+6kAt7o+LA7rvjMhNWVflnKAfdf
3504ySju1g5b62wvyGjcPY9ZhSKJvWdx0x+DuQ6hdAXetmDxZbR5R/VwmjJe3tAE
C+lC6IvEV7ds4hG/HmhZ4brK/gx/cDCe0lfbpfGh+yBL0PMsYral0YGy3WQMb9H1
BGfSCkG3rdmzihu9Eg82KnIYrqj83kszDv1XNr4gfbLmhM/vzQklFKnJx08nYGKp
RQMF73XBhw26h4bQWXd0DefI1wuR+SKL3lrnJcKRLZa/jRwZSkiJqQ+QWf+zE2pe
OJOPk8bUj7m5MjTrdrlAlsGQyokJgrLkVuLi1XAI+rnpn55lBGTY1sdX6OAiPhZa
26NwlGvh7HPdakOzEYqEg6tyKcA/E6JrW5QXPB+HU+j6VfKXMqV+NE/AH4PWuz2J
A6VFZH7nP+3qim0qgouu37DQwri7nUZE7gd4jsGaC/JWAUkSNvOkK+pDrIqQHegk
M9sAJTaMIY9DYpa3E5hQoUV0QR7qY52AFqYNzWIvjPxaTmNaJ/WNdnUwbpTbsT4G
/eMafmA6SFx8hIlGrVo+69+e8bkmsrEvjbTCmx4/jXyJQg2a3baaR6xko/leLroa
3oCGSbtLqfO+Iq8s5dmCvYkjEH1EaxnIDHjzsO+hqT15ioq3xhGIy0DuBuxQbJ3Z
fjrlZ+NArnkJ9aFWJCzr03Oj3Jf4U/5+giFg/Q79o6kyNRs3WucodpTtUd0UUZ3l
z5OtKvuPxfiFVP2VvmGzNPkJ1khZ8u959NhkUQc+V7KMM4TMVoNa0icwyIuMJq7O
1Yb0d42lWbrzniozEcSGdFmqwtmgLu0luRhS6rWPSdseNHrUGDrq8T1ia/NWD9xg
2EKr0PO2GRagdHholy28pq8rFmhYj7msNaKt/UKed90wo0ak8AA69lmC4VhIKRLV
V3Kh9XbQqljee3kG3MQrUA+vqICkT+UrBrdj3RBrV/juVlFGEVRDUcK5Aj8TI0W2
A8mdv5u2yAbGo/S4SSbkwDDmTMQPrgNDqO1qcxOBX5sUqd3W0xkWcJFwIkz+ZEeU
EGndCX3j9WIzbV8Zfa5kvQvm7nCVwP18MXrqXATwyIPPvDw5FHoquIXGZvvdKDz+
OLFdwonJnYMYQzo4W2s1mBy6WFOrMDW5ibkU1inE7jwHX4IFk0KSbUAg2w/ma3w0
pYd29hcLpJTxCIYN86oE4W0zH4wCHDWCrAZ7/o1OLfWwi+W5X1wgDUFenRuLNrtj
vbMgY4Znh26p+MQBWxjBa0ygHlfLZNkiAC5Rl1gUxbwo6oCjgOYrMlKtQE9zl1Hb
gZn0alre2BnSESXgtXMTvqpwGYgPzb+ZHF5fVzWu2GHyrGSAoR4AF79VfpO1osI1
BMZIK26c1kuwzWuF1o/1BPFI/jvVc9HszTq1V3KP+WUSdICe/ZmZTKdUIXy2LrN1
52xNSGBsx6A8N36dpnFKRZt0FTu9AWry2tQWKG/9csP0OjMW0qBe73PIMqDECHh4
nHdfwq0JP7pkVTMJGk86KjZP9UfeozM3rnWbhkIh5fSz2YMm3Z9v4h2jSJdTJwOJ
5W8j711kyLb6ECwLMJzhm8KSL3RXccz13QRv+SqWsqfP31jiM8PJ78wdw3N9p/ve
Ziyg6TcB9WygieQEfJQnm0tqUn+d7jLxfPbBStPMOAj/du2oPsQinHJitT37OX72
PtxVFdB1agNaxH3z3m/W0+RoqNvmD+cIZEjF7PeW5rBy7fCieoicAxWACvM31k/x
9bJQ/0/h5IW4XQpWAXPR4zBhkrkMoH5WSUX8e93yumkHrBy7lac9iJhO/o16wZad
QEfemRm+YIgvMHD9Q/lxP3FcmafGwui1kAYp1xQapMFh9mKKoL/Xeahd65/d+8Tm
smzMgRJvQPr3M+PDJnKXuNTctcQvODQYbOLqj1VWj4eDAeeQnJRh+GOmRdzvXsl9
VOzXItj/4XhqOn3WC+Gv/BwdBNdxMQPIFy5ItU4cizspSnFkj5ZVGT+lBWdemxw+
rCvG+Fj5IoWSQlwZOjY7TtVZeSEobu49Pkfy90/5BUpFdRh8KI95GK+faPRFzw8A
pDO95Dh0KE7FBEBTudfOoOkQVXWID8EAkHdG73ahj0hUr4gEjCm+Kv4xTFUQl5Uk
syzsdMejef/2tS1UEac1VBjLyMu3xF5huWClCyO9zXoVbQqI9MOG0GMGaB3P97yD
m69UimDTT0FZA7Ijkm6YoOK2XCG731WuvVNbhaIdwqK3iZ52gy4ozVmITxU752y7
CxSgjpQNsnjJTh1ZkdYM1sDQ9Lrf4USi+epv2Ry1op7c+18TAVm5PYqfZwGZn8Gw
7Xtk48YVuQwQD8Sx5CCjMfzpaq4qpUuxQP1P3guarc9miyAhr7GWx+H09uF9tQ82
cJD1sj5f1cmpxZjjyBUCh6GweAxD60gpkWZAd2D1O1szqWax2UOgz4GdD53EP5/c
+IMD2cZLsSDYQfIKYteeV8RD9B20brQB16LZHoLrSIvkjEOT9GdUJeGVAhOich3x
dg2xuXO5MCNUnr0h+1s6VM9Z+8IcXcP19qiE1fc8zUIKD94hYPqCtILYQhoWGI1H
Aa1rcnZFRQQp8bK91IV55XD/JD1zwnea40RvjGvnlSmPKzEn4gFTytu8/sKsZlkj
eamKMzkZ6vlGsqHBVWctCjrlE18TdMorEis3xn09Elg2NsLc1pdat/qOcfi6aJBC
OWAWPkehqv/0M8jZHgFKAsYNefjHCzahArBUbIxqjzGLP0gc4352OnYZcpwKE7eI
BIk3beB8NR3zXaL8adhRVA5KbxXrMW1OqUSmSLY6pSVDglth3V0yd/FY0DMW/nnR
BoeVhCzVjrNhLV1Vt0f4s2VhBgCfPX2mOlNf1XDCYeYrnQhzQkvkcCRq8vXOQfTf
nXFU2EWopDrXFmhwPiPWniNVvR8GogxZmFtrRKn4GuJ44xR00YEja4ldUFqYZUVm
UxbVN/psw/nPWVQPZueyNA8LI08Mu9l/qeIrRBBl+75cs3jfxgh2jutyROuqO++O
edyeQjIO96lvP0uC+X0YDok8pdCCB69lHwzod5zOJzLsaDnUubNfzBuxsOa2SEDN
S4SHXvKrh3RRSPE5z59yUfcKo/32cm78bNSltBfNALK8X616nsWB/gyb0Q9KR7Cb
kbjAm+ZQI8gLKFJyLW5EnZ4skNjSITB25GDCHhWU783/y55pGq8LJcAnIKbJPhsK
1VCSKpfBK2c0/Q49Tyehb2x2RA8XFYJheOcqQMJmxz9A4EDOghQZCx3Tsa/QRyIF
QnlzxH9N38jF8WSwecvzbBTdiVxDCFXRzhaS04pI8z/dVf+CnPXRJChvzUJtHjwF
yzqV0wiRiMv7TgLdB0WILDNUcxm5Fbe6v47PvKn/b3cycHyr+VWbTbM7+Klvt5/2
xkAAorlty1IBr+9XQ7XIzTg6k4CbUPhdaDTo0QJJPQMxQeVcC8qDcxBiGJnBtcIL
z+bjBzea/2Ekbp1RdF0AIEd9wO64PenWUVnoDUwJzDHmkkHXM36nD68f93imjZzi
VxeYTy75AmPYW8/LGwy3L+K0oikogYz8a8njMBaYCiXiBexaJLuV97gGy36Sh+zv
jCYFUj7hw1F0JV+k0J72HUQJe0LgzIdPR9fZ09GWpFZMYDV96Xbh2Bxt/DUgcmJ1
AgJgd7sdLak4tDqfmi6EA7w/dV7l8ekVTxKLtwAAocdPXr42dD7IFDaEX06M8z+S
dwlnBrOL5OPIYoEtmNwZbCBSv8rmVWOcu0LJTbZIPAAtB6ww43yF3MKzVW7BNKSK
f6yYvS7Hm+53+rvZzQDe463Qr/OjwiCzuHytJGRWxv9yKpFHgv7upnpkUmuJ8KY1
R1lTiUXXFseOHT06F/A31vtBVh9AJUOnjjVK4rrealJbvNWLhYVsJCDz/9Zk3MBU
ZOjbitBt6RaYOl63Uv56w1SYiiZYq7SzkG3UeIUsLW0Rtz6FzhasBAGISmuBMvHT
PZMni0AZYP/j7rKhIAwst9pwa3x+o7ybAEJ5QK7apvjd9KC9Nmm/rsV6+BsZiWAI
ZWlxrQ1lZZC8mvv7nMGLVPgbDONIMm/j+kK9Mg263uPMpgclXYiRjHvwZFPco3se
KdDDGsr9M+ekoJyGVOm/TK82tCzbM0XrzDn4jcIGB1B9SbY9QN4vhVc5E0Wfkxaq
9SEvNgrYdBGTtJS0MgD9Vt3ON5b9p1D5Q6GVfWdapGx+rRNOj57i9jD+RBF0IMOo
gxHWYBcxifNbZib543q5JvR/jdPaFIDMGnCIjy2px96gihDmsKye88RuOmssLKpd
v3Pwr7qu3Nc6GDKQl/Js7ekZw1HLvp68N6BgkD4y/8FXMqqwVIotfFHEHy8oNDlv
8Zeu59efmWvUXrhNm/ZSTC7j3A47RnQWx8Npewl8e+HwhPJJjr903TfuYXFh0Xo0
y4Lh8QJfEdFMgvRdWCjyVQte5gbc/G5eMXh05EDh48D/91jrCqGYSygadLI/Dt33
3QI37RMlPSCOGeKzWbPIwSKMw2jL9C12VxYK/1cIuugyAVptWVKxr9zRXe0kjhX4
Rgre5rA4aNckeR49tWwx5qEfdNMx3oe+t2AstupDVGc/IiIWSc/D/CHesZL2fgX6
TGOpasKYyFfeEyWufAArWhnZ5dFGyxuLG3WR/D1JWoozt5QI97B5hjrTRRtIn+9q
cUecA0wALDXTE62webU8+5EPTwTc34IjXIaAF/v166WqqvDYfHUjsWQ6pCcSPnAz
x5wAG77CoqjqFFcK0U69XpgEz+chdp5qBCDa2FgJIfT0QHr0fABVselYc41NrIrY
AVC4x0al1e4CTIi97KLN2QMSEpPfDz1XSOowEPOFrRrh4jp+No2wa/9y1RrW8h1p
EhGfWkGA34RU2P3Um667GmNIGiky6rGx5UzoYd2Q5Yqgb47gPheN2yH0dBynzl0G
OKfCH2ogUGFNN0JLyYwtZEfbcfghllOQuTgLHlbMr7Jh/Mb5Kmw0IG3SAzUxNdmN
x2exHajA7NtWiZXIRf1YWr5flzspwthDkYXhVCPqWH2BwypzbW2pih17uVBUEb/6
qVcJxEfCJu4nfXWTStj8XH3uGeAZPrCu6pxN3xyrru6mJumQs7fc29hO6JJeYh++
rst/W0YtmV+AYs4jizV/xTKGlk5JFf4QqiSA7JvFKuCvlKd68z+VJrLYd6nLvISr
NyP3WaFE6wzTeKt/PlkiPNdhwLYCG6UGXU4jTRhW+eLH2q4xwJwSbkTEfBBZkmul
9Rv7Ulj1NRgpZGYFfgDqMbXttkmgOuiETTsM7as/atanEsOM0yoC//COo2zKQ73k
iibYmDRUhnlWKAmWmkExzwBKjrq+Cw12okoEFG3/ciPWGHF8scNeXoMeOaSAisWM
ZllF0ct9hhMdbpcLForiqRafa42dA51I9BZWp6FRfpbdtdbcUPmDbqFq9/o3X8B4
EnCFsu0a4Lpei46sPqqAa0NC/ZCwx3ekfovnAGPV5H85sm6KdwwJ8LFEZrGh4sf9
jrWjaL7eyaSYwH7eC2U6e5lb74vx2bWByyWsICBnwyTjTyrktWgchvkzynzbazXr
NqFSLBCT1UKrAlBz8SzLwZpEmdOYW74DDOR1TFYCnXMhR1kpyIDppKssymuirgVQ
owODYB0Hz98icjGGNAMOFpoAoxmK7wzXKPMXdIg4/6O+K1BRvNNCUpsMvBEZwARV
hWBx4b5DINK7f5Lcx6ll82Ael0Thuu4+FJWhwm+K+YXukXRbJs+E7WUU3Q2kTtL8
RDcP/Sen0YptdfwoVgSwqLQ//HqbLdZ5ZDaCTAgl9jcGwPQuxzqQQmqhENZlH3mf
hH4T7/wwBeWH6zYv5+G6ESdppjFfABSwKjfHH4eAVjCPzc49IFTLErsAm05LAFEA
7OIxifUZmBMb4xea8EuaTn6aF3HwYSxasT6e0HXXuVffSbhTNrgWBlovi6znRo2n
YanN4YozBOZEeT/ouKmvpyKX6fsHYZERvKWSAal/xDTEtaSQyZHkWWgPw/lUaY1S
PY1kKV2bYEnBsdFlzYJ5QVDzken0XUa12BWekNHMS4Z6M9Dv1lRH5sHKBd3Z5/I/
fobgKBrCK9uN7gaG8C2DbpdcVMJVLusuX5rGw1rWqxTw79gn/A0yCT4fJx5VQhhn
bBmLf6kLWwE9xjgaFpLkfrl65N2kBmeA8hpsmrAYLo1S+kElwUYp6YMru+OZjrpy
s4sP6d8tXiQizaa6Rk0msf9TEIA9yi1MM1sZhaCnM+g28AaF138drFbdJznXJ28+
/Kf8yZQ+VDCUwfS9m6Vfe0wWAzqFrRguarau3ytKyODkdhPU0jKNIR2oJdKbVVhE
Fx+JctLdTdQkpTZQCHyTf/rPDeqU1LEVMM6wYevIvgt73SM6Fu4yPVpDPgQ9AHh+
AGsN00U1r2AfZ9cMBOM6Re2xAH3SoyqK47FPVTAmcDOWiZ4DqaGXBomGBhUN2nXQ
VJgOMO4vLPgEga1l99kjpjdLzfibbRXnr2EuQ97e96u+yDfpgdVDi2r1Gpa530um
agFazupeWjZNqJmTtExuYNFEiaqzRxWGI8VSyHoFGDdIteqWJCNJnro2T3+AW/zp
6Z36itVDaOGAE8Ay7/u6CfH0X3++domO03zYsxnO/gNgv2xJm7ARUF6SmdmPQ7GQ
ddSuwLn/47TG25kirErIqgJTKxl24OgpHd7XJ+M2TbcNX3YY43cmm+b8uW7m+Dlo
OIr2LyDbl1avZ2+j4VxMq1TNK20ShyHChktV8T5xH3fVxrGhMX1zI9R38+rjdc72
Q4zQnFBQ/9phrc/DIgL2Lwgbe3t+68rNlc6lbcXUr0tcZf8j0959HuM8mqMki8UW
QR7G0FnkmwRCk1Ubm2C8PNx2sM+lTiXtIRrXDb7Tg4LUzwrYIxTku8DSNyoGJerN
WD0wiBFOQeTM0inCawJHDRZ21niIuyGIHfsBBWh6mk1FOdbVPhToCp1bIvIeUf3y
/uHOyBZGTS39YQjYu0QdYdj+RSn5HmcLuPpLuNxGDAn/uc7cbI/REnWqR+0mrJmP
kl6k8cfpyx5H8E0dtCH4I3a5cH2xMWvmf4lSF5Rj57uiEYNpqQqBU6EufItwYZf8
mwk/3bKVD83o8rdtM6G7gf+hz37tlzPdtU2Y+K6pHjIw/UZHmnJbzz/gl3Sg8SeN
Y57E/VjZJ3iBwvL/y7xM5D4IK8nD5XQr/C8Vm/NP+Ioy9qnBRDw66ZvI7R/WY+v+
IWKkdkCYjm8xs8HW3/NY3ROIG7s74Q3WdupYAXX96HrsIIr9YFzcGpq+BxCe+uTZ
1SeBq00ENSrfnlN7NJJVTxz8CFImJuhnU02uvfAYf8ddvsnQF+4jOm7JBHfN24Qx
BRUx3ge8/Qa9YDarlVhnSupUtGXDzBT0zZUndJdFKe3M9cur9XOzrkH393fq/LHS
rs6R0AOVFscGkOUagd4ReJC7SCje5dalUzE0QwTr79NgruLb7yS6K5BHqaAE6gpB
buVD9KDPhSW1GGo/jIUg+io3nKsU5oQUcT1Tyd0OffnNtPzVrdqMT4h075EzuHsn
ZfA4ID49IpNXQ4REKIks5PlD5RYrHT6Uy7Q1T5rgJRBg2Dp3XJoFxxpi70hHUfYU
2FaNWnDfWG6oq2oD2ETxjScbdQTgAHHceCSS5srz+R7e11jAcqdrNgJXs+a6wQq7
oqp4NfIcRBlHOxUElfEWkGJct9T52GdkUHMfGNLUOtoMR1vz9Wfa2T3g1yDHWI1U
/skfCdaFsWTUMFCiEyRtoq6dQRQAZp3Ad0DN2LehRlSqDt2omLSq488ckyrXS1o4
c9ZM6Q+1rcI7CKPaMj8ftwqnfinQv/Ly3i36g1C8FGbX1IgvopaJggShMLnzZZs1
VuDucnkZRqJBvStHnaJbtHWyIiKiLAkvuMH2erRDNshz5agzvQ1dTkchoNd3rUBK
nLJxyneKlDaIJwmLEYcNseYUOv/e6GNpnvnPAW3m+DkgfLNiMggWg0HSG2nyUQxb
yrayyVLbD/1jHKvvPS2MaCHySYOVttOawCBmMm+bmq9hrx0Pr38KstASQESrpaUg
g2U9TwnEamw+l3lccgJWEvFxy7Qrr1VRXRI7ITzf79h219BRlLsKwPPj+RpHonu8
aH5b/sv2KboKelXO7lQU+ceZNykkdFVKtbWxeXsP1jgjierlSxBHrTUjB0nvPg8J
gHrkGGrzHRhrtecUxRvbFpvOILC+zrIakOFOw1+mtZVe48mHp6Ga4p9lhcxJsa6b
SB3V9ihFjzKUkPMo3AAY2XjkC83+l3yF1pgkF3R54BX5It9RqEZubo5lHvVR6wQy
+uQuyRQK4A73ndoAqPUswcDS914B+ViZsjrgDqZNmr6+01gPQ9WrKisiXMq01RBk
7xznzEjKI2J1RL8ApPahWaOjCQODhbAw8BZ27LWYZl0xnCw+1WmnjVe4+8NGm4+N
f5rZiowQoMRtSb06MAOO36X2IB9EPNXKl/YGp0x5+z2Xfr+l0NgGUW2ioK0Vxsmd
MdWzlKLnCRe/k1INJb8SmixLY7DiukzOFpWWh2lgnkkNNMuiUNvQPzQTa2r2Wgm4
PxjIxJvWaoiqkO3rIDmgXK9A5kDOPPT/2iu5y04D7y7OlMhMO9UdfN/u8nim7s9F
s5IMvID44lbyDYGm5qVWckMtSDpA3svLMTN+6KhXZdGL0DwxzwJdaALuHdXl4U6y
r7Iyh1PPtQYdI7cmvLqzjpbFyhSFlszUcTaGRSRxP39NnW4sjHviICfnKR4lgYcY
B8/4+ZnhI7eFgx61BhAamJ/iC7UVWof/bgzyKEeTg6Lp4Morw2PtBEg45KrsPdVS
4jtPpGdMNxbyjbwe/18HP48i19ULRQ4J2Bf8p0QP6YE50+YQVtoKNKbHYw5O5zoO
9fXUAgiHua5uoiuq2C2ebroIbLxZPhNvIfN9S7ayjd0+duQqerXKkSzXUSQYRKRh
VsDmLXOoMkArDSypMkiK3vXnecbX2P/FxOx5dQEFr3LZaR4ogLlU3gn/lsrHopbu
wplYJ2z08edAbhvxkoyfCJKXtQoXfwm6lsi9uHPWoB9NQM8Jt8NITx5c9yCYMpAI
K/CDvhK41yBaPFKPKlC+EFMH7eYoZmyfMUb3dgeFwspDoT3HoG3cuTFpYSCxz81o
flf8vWOfpNFMAIHF1wk6dJC2HecrK43VU1KGF1gjL8KRj2t7BDbdJhgckAda40Ov
mh6TLxMMXZh44knyK3yCSdn4C1y7i9f9Lj9YJT72cfM3xSNv5clF6CuydnLdAAoh
ag6HzDtazkJaqdDqdZd3+7gDMTrqurCQHxOHtgfwVuNrCkHzvRf3QNoGezp6dI19
IfLQuTifqjPHiv57bOSXKybNDyDNabn+mXsAlIUTuyjIfTZyr4gZU2ndr0OWSlVm
RKs0c/+tKTBpAybvr2d8EMkAq0f+NHRbYdRO6yeRz+OuzbIXLf4nmr1AeuGxQx4K
7b7DK48sZebBbFU2XvEmFxGa4aeCgmJA95LHsolscV8dbu50bzMH76Zmn3CYZQHy
VfKM3crS2iBuZveJrnY3tydmqiTJ9qmuvSGJDkOgLu9Rpuk1D2Rz8PmgMb6vPGJV
1pwE6+KK6p5MYxKi0zXBxTIuhED+ysNPiJK4WaHS6QGW/c+GcR6c19GJJnMEsXId
WeleVQbmuM1pJ4wAbUjYYrNAdV2VGlOUZdOY+eTdNyu+ZTUzlPbSno0Su19C32nC
rKVPwd5eCbzVvbGpOEpfkrRIxbpP5BdrIavZ7cKfteQlLL+rFE7N8hxz5wxUd+hh
hcIxTcUm04aSSQGPuuUoKqH7gXi0F/lAJVlJzrz4nSNbxS8GdMLg5xB9+Jf1cyc5
dWpC9V3E8/PWsh4rDJ2w3IvS0Wx53hJHujhaEgYysUwrfP4e/Pyqz09izg0+fYUa
So+Uh60mYhjxCVDSL9g+7e/XESvP9Rv6odQSpoGExZ39nBklZpANxxASnuYtFP1H
lVSTD8Cwoso4wgMe0V39fQK33CeIrVR3p0UnDM91uOZOmDWhytSSlR4Fru9+2n2I
LBKNTQwneSnZ/xhphGeNoL9yajE3NaelsZEIRmV81TIJjBGtDm2Sv41kE6TcybPJ
gS9Lv0+OiWgRMaMYmloR5MGCeZyGIEuBLpao2SkH1l8ELPywnOIKOIyovqhGzlAt
60cjfsPJHuxHs91/PF0JoOSrU+I4SvbWhlibhYCiveU4lqocpE1PxwzKk4RhchiG
ftlXUOfADhbqopYttV48JqCQTW4ed1n+nZQUO12mI9Gt2Cm/UAdTPR936TdaR8oU
LYA2VPERcK/wVLc8Q3Gjw05Z/RPbIWMTCOlnNAW2Y2BpfLKPBT9AHUILmBWXIha9
rPddJHgZ+Q8YRwA0OFI97Q1sDjbOFLc760a/sCSkOczNDgLBOVhvIPwyhgALrKaL
5IhuAjB0HOw7G0jo9nD5h6ndV9OyKbiQ4H1vHb00nL7MdrZurCpEWUtWIMheqPDs
6cdMqffekMwh9Od6Kg4NWQXsFwVe3jiMk2AnGMXfr5ffaoFQAbfwjFAGhhGaPAEV
89+JCJcSg7o/gcmLnb3KpwDLkF5aYv85KTXBAEC2hJsQhb0eCjQ85PjRu90JdANR
jD3eiLsj4bMvoHJFtnML5IxkjAvJgwXPxy2Q/3eJ8gfaL/03UeMm74BySOUD7u6b
K8vOMyS2KaY1bXSSMGD58wHkFJbQTNWSRwoSkMroiROcVq/blP+7Yqt0Lv8l2Tni
xSldZcKbt32VMCllzqdC23goAGITIz5SnKZq9LK1OYCvAbkMXYEJ4mJj7v5w6A/x
OuOFSmToxIVgSh09c4iiHqPb8GV8H75cnS7yBsYeMGodBovV2X/drjeKnZNM5dR6
kWED0hNQqR4tL5tt+NhWKps004llexRRylrvMBL9LEawgB7hsrLNOrlqBYV9u4m2
IQmso8W5uDsmpkFm0CoweLNEHjHovNqG/IMpHMuRpZdvqkT1QkHl4PQRge+eRDsJ
/nXbhldIU6XKqFjiJ2GgTRvzZgjpOQ5EOm1zQmo8BJTCivkf06ohXeZ8x/Un5m8I
MtIWwa4Q9yBSb9VOto1wHYuQSpJMEiVm8e1YKMyzDrwXLtNxYfjpc/FFh2fnKBHO
9PB8e/q1JNrjxFom4b/N6y07Lk0mhLxirEUFLEHlge5BnsOPooCzw0/ESVZzkJr6
GILX+jjq+78MJZZesCrH8+OME96LJ58qhihLffCUevGi41VJBjGBPil0fRHfYmmX
UueUc/Fksw8QRgHgObdZ1X4wbj+cnkYpB01ZS8m1ARsaRhbCvlvBQ3DFC4QHg/40
yQ9y0WabrSODD4sSlM4VYie7yY21KHze8ZVgVtJWK5M2KurwKEndhGuG8z0dQr4L
peVhdWHMW81MpeskH3fJbR2EpxaXE3qEqJCOpUo2UzuDoMBdl2ngJbFjt57I3PNe
ML5KbOft4aK//U5UtB0Yqg8jnFYSh0HOSmtroDuHVDdMxHhgpnx9IklOG8gzcQP5
FEClXSAlujU40jRsgytAFASd/mHBOUgQbUX6kEEWhI2kJJlFXHsRHh/PF3vPiA2D
AjH/0Vdk51SRGoMWqYdKLKqAj422yT0MucJxzYA2J/hc0P5HKpzBjzg7cO0jtp1F
vHuL0W9YdPicJQXdKqjfaLh72DIyeFnVJu0w6Suu3gh9y3/4Jvj2lqIKaAeMkDnj
8MWqYUk5k5m8ulOVTWKJBTlepzR6MsOB0V/rl8o3CLTRisAX7MTWn/zXt+kPImIC
Md6V6K3OhkPuoccNTBM12clq9WJ7f4PqL6HTbNDybov9JiQ/rS5n+t40jUErKqGz
ExbkpC3jkKZF6YzsXW40TL7msRlga4ufsGkBtahVJWexoB5dzYiAAQC++/Gs7mNp
DLagiUfCCFn3//X+Lo322hOMX0KJyrKb5uFgx/XDrFCvFlHOOd3LZJQS6EoI7BVB
j1tDlonoOW4rq/2UEUYPl4py2UL//LhFxkdo9fkOO07wMy3SgKhI0ST+bBJ4YMe4
vSUQ7m32RPlnjBbMdTETdZP9zcV9kS7WQoAe5QUIiKnkampl1fIKZghmwTlqR5gd
grIXE1sOhSc1jYP3qB3v3KZDmX2kEMmeFn6QBfkK0xX5lfBDRZ3MH17iSX2SXM8H
0DBzW8g4UzBU3qK5gWYfFgKClaOILN4Joi8QhIc8zXphpoSfVf/J2p+Eze5rXa4N
x2Fh6onFyMkxLkCgErnxF8vYvGYhNAHC44BmP65E96808KF8ACrZr/AT5PYwxq8k
sZixMqo8vbMyT9Gb2QvfNIuzKwDtaNCbc7FTsZgaeJKDt6djv7Vac7H/aX/xHrcD
0nc7WaRq9O7VU5xU8sM3ObnxF61df5EQX2So1INhZIyRhOADMSMzeqGHolHXMOBG
zMODf8xnTrBMA4GAIDWqOrR7X4hbLC4WySOeQhK/mGR2isGyhLn3LGCl0NUG3yQO
LPyIJYBjkpGbWKussDp2o3NwVRw52M2KVP0RgnWS5FQrGAL5r3aFGgF2uyyMVYXA
Q17OlAebE2W1sf8HY70wR2p3+ZbGhviNmPN6t6gWHPaweDQuDIPsN+tcR1FZYI+X
iSL4Fmzqr7B04+fhY91yI6r/ZX0HllnU9t2EjrRTdMdeANpxEzroGRQv8z37QMHG
UJNweJQnb3A4TFlf9ICpSKdnqR68F9cgYN2bRMBmfwaMkNQ5sOPoT9h0rhUrxyd3
AG/BJefyhcr3NBjoBVc5BXBWPoZ+OdsgsZ5NdlYoPvUlgVy679xtJjRJm3uYNpEl
JqtOFYWSQOqFGp6o7UrugM9JYd2r0IdtQk36JbmooCO4hlSz/+4pbPdYsNJmMdvJ
P4sK4oskTH2h68VFm4liRtZvGxL/b0bkAlJqhbWj1Cn++gnOhCSrCZzYj5YLPxYZ
o6PwmdALs8ocHaH0ys92o9ewOPFZ55VNuQBuOz8Tmdvvcf/t+9VGsra0/s49OwMu
4xrp3Oi4oVMgMQ458MZqNMukrKoBkHlniMwbBQ1sxb360uGZWqxM92GcOJNluVlF
ShWW6q1pWK2C64M0EkuznnH6QW2aYQoLNGMwk5GHQ84ImmZo4pdpzE7XOsNhx3Dn
4QC/tT7GgxusEZF1rZbXFiubXqkcH/lin4XsLEccxf15eTl185BnYpBXl/4gqUFS
ZAQUPbg36adGD25U1wNgVUzdCKfL36jNOTuZsjrhf9HjscWH51C0LMxCWth9gpKj
HEF2fFRUEGVlRiZdjndSQwmS2IYcvBUdDbR5Ct2Sd99/gBOHdMdflvjCzSmMSJBH
L/UhodfJrbXD1yjVn7zd2gPR18O4OO9U2rjwy9/0QQr2891y4cP2We8/nVVLNv4n
CUbzoUk7mgtZqTN7aQJ71uY9AZqU5MH7piYolZobXkRIGBdYCLHb1PMKMDJtFrKx
jVsXWGGNpoG/cXbgNsVI8IC0WJcg5D8K6cDjDqAIQSFuErkc6hFVvw4IyYJuAymU
c6GGvCYyFvW7h8wBXMhWn2aJjMe3RRgsxKKOVBjIPhVe6XQ7750d/uzb7HcKkRSH
FzXKn5ov1ygje4hCEraX2qBpNr51wJ4bDzvEErvJa4RwVGfToaVrzMzklpiJP4A8
b6hDG/PwuMYvoguobUrfoe1GTfbmWn5hyT6cvySKudnvyGrHNSAcVPCQdY158u6m
CYTD0rcmGgUR8BbYbFCnJQtW8PKGfWKb1DorvcyADYcZuFSb5Loube/gQO/fIgV5
2Y5jERYS7fM4+kKwTfo77Hd0VK8FBCN2IwHLygAWqcjfhq9A9haDGsPNqWK88bfF
KeZasP9AmLnIvU+/XDUQZS4kVvAj6LOJ6PxA38DYRN20n6I22uancetGC1SoJVfe
G2T2/5XciLZHHi1iqE9eliif/rBglLx5po7XKGJDwB2XtHuEcKBZ/+zxw1L7dqQL
YRTxDDoXfXHkKvTgrgz9Gon9ZxU6UwpGQphPv3xZ9Fip8400+yfLkgD0Q48gaKYl
7Nmd8BMDxMFxxnZqx29PvvwItFz8ejQCq41fZW6+AywIf1BdAA8aq3dDPMLEn8s/
HJE6RxkDnZaftndSU4EAYDQU5DeXkFBSBLNzFpuKorgKGx8wN2R36019oZQAWeGm
Nmg1b71cL6WUMyRVC3CxOw/DQURWqNz6rOl8Y+NuJgUxEKMRAT2zY4HDPh2y2o/F
C4BoVdm39zTyiCaQEntOIPMcUjqtMmVqtV2ekB/Z4pjNB40B4aYLJmq3iKGwAQqr
8Ojxclcygilu8jTteTy6prxjW95a6ToFBU77j+2HXpcJIB560FisDwffnjP5MXmt
6zpj5zNRRnkjqlvptpW3Hk4BdMxZkTJNxS7/1sPZh+QW8Uk9Wb9FcAevqVnJwYYr
bvDQ/R1wSyB20lEi/b/9nVyL4MKvyNJ2nDfi/29Dxq2EHc95QSZrEsper3C/Qc/1
z0v9JLO0h2my3QM931EHhFJVEAlDzTP0HfaL4YRFzNnYBCSutAolOXpG8/WjmM/P
YHFpkMRZtcYfQWsI68JGylOX9Rljyf++ibmmSJVzh97h9WohFi9jupBKaRL0c+Ly
hQ12inxu8K691irFDRHNfiJDGG3Y+vDp9WX601KphmVji6kJHACJsqbWT0JFKLQU
77XLzGPEnn36PQOYrrhzNuc/iwAqEv+3laEtgosmUUurS2KeDenYoumKH4YCvkfo
SX14tUqCmZTd1QW6/hJxLV/DLnTaiK5Wa0hXjpqx3xuziDlW+p91sd5XkpCgZLEC
Cs5oBRbvh08LLzQDSeagyNO3rMkICOCBnDOFYCgXHQAksXw3R4XVqSbq9g8WJ8Ml
aF+Wb2gFTtsXnx52arPZF52GTjM6PvU96rqanOZmECu932vLN5PNLmQcCTmqFRiA
3ZT0aJ23PAr1f61nB8TAz9PevAlQmuYBbSuCQ2VfO0V4v22nabOEW+rbz7UU8t2s
kvHRH4VXU7li2/ARVGP8BkTEZgTIRmpDiPOIYk+wkswycuf5h/igOsOkjo1JQu4B
baiqrq63eDo3J4CdOsatSx8d5ae3hzHMYP+tNL4I887mzTAyald6QZY/+uvvhIMj
/MeqmFf9xhPgRzXA7TNLaRVviGeZwI4XHAACDNqxRQFhfc0nAZ9Y/JipVOJzecVc
qyTESZQ2/t1eBL9Mx3MYkqYGgONiineSTE5CI1FXKLffmD5w5mcQWR3IBkdqkWZB
a6oOhet3VJx2cmPUAfnRqQzi91gDuhfZu+ropDgfMKhnnndHd6s72PS5Si/MYKdb
6VVOmqZoaLsDJ0NFBdpW/WGx2Lr4v9QFXNrC0gxzW3kdPPER88K/q+iexr+suSot
CK7E1S7PkvV4RzftM3OjUKdvUVjwU5epXXDnbf+2+mjg1DP5iZBAorT3P1kZLYHd
A36Ul0GSg7RXR3SKQBBqtrcmU0Ir5vRiOgBuAhsivRBxhJjJfHLof3LPrb7Q4hSi
mtEJVS/mCRrKlRWpnX0aSprpdX2Ub1KqATUmsaVcxqOjgVc4qHzyjFrPzQDwVPsr
TW+fvEBoz2m4lvMBJA9QQztlqIVjlaA2FRRQwoJMIEXvzyHG3ih9eAi6R2iO7ZsJ
DOVamAo62pIN9QmrTbJpZROo2ZoRslJgpN/n5yBXXxy/wMTWW1Z5DvUJ80uUgBI3
zKX12J/oGR3m9fBIerz7u/j1PMZIn2xhWm/pz/cK+mHEW6bgneCiU2TrxgGcnn1X
BACLjLKZ+asYmiB3XlLBRQnndz28cBtr2asM4rmFE8NswL6bgeoXFx0HAOIk3BPB
9D2rukerHC0KPZhsbroF40hYZ0nM+VgvasIqyOsLZivvFGcc1N5pJc+2RnEw60Rl
8+mCq8R1N9Dy+vhF27Sz8DkyKf5KeoYIpqixIGyYSTL51YrulFDQAyinGlhtqTXx
dM022t8qbMuQ6roQxMcT6zTLooVxO9oSSDSmSJKvDksBUyPoxZj2kqvHv/9vpcuU
jFSMzdmDjg3CAi+1dumAvesQtKD8HcCjoSVBtuSy0fHK0o2UiuaxLfqcg6U4+4zY
SzAda3k31Ms0dPERoD7Km4Blu7ZhOxgICw1+++5sCzrlUDkq5XxAoeFeEwurEsx3
2oyWblsYSphVTaovBOXQFFWW2hn4a1MN3RJsfMfjnRLR1LJDK6KZHHeXR0+Rm/Sb
OmkcJnq+5OS63vGIU6w2xyyifw3FfKSRMj1cbOys9YIMz9G8cQ2o+z+gNO3mzNKH
GVfGnv6vYF/6Mhzm30ecOk7lHwCaRjfWstf4xQmfv9eQAShhH62TOVqoJetqZXMO
NQEd3UPOdDM482HhWwHR/yt+LECmzOK+ouRvWdoW8VmMLeL9STDUW2e2ywwkpPMD
qgZ9qzK3ETaqWR75DryPceE+XBmQLN7tbycFYq68GawJTBpzNHC6+IFLlD0dIB68
eAXHWu7358uDtEuxOUx3lCQM0jzNGkFHTO+rtzWaYqIA7uvbLCBUd8vNJ40jkVZX
ZE9Ikjr6/rfmB8HHoIZzdjl/FaGaUwz1gwGhq+r1HNNFwnEyOOlgmwjpy3W1aESK
sx+MRL5zTJDsyK6zpq2imBTbMuMUm5PSuUJLiJhA0MjUJ+xrJay2IpYRD/w1tznZ
R/XVFN0YS69IWnOilcqWYCLrc1Id7IZsiMHhNdlEUiK09xRsIIIfDFHgilnfsE5q
dG+0TxrH+9Xe2SbD28i/wdWN3CX2fal5jVAUwHX4TGTzoS1ueTCQsCyy51p+gOHC
cLTl5bTkfP4Zb8YCxdJj2prGXGhwgN7FBERdqLmr8veFowsRkjb1NKVnsy2fbkAg
qfqlBEsSQF2P1vmV+c1N47TtqIOTnle7Hv33ruKBHn1ArlZstqtAHRSYMDkC8+tT
V/OIMkRx+w2ukhlJ6WiZ+a3PG4rmTWXmv9ozTp1ZQKUe8UQSih/PZ6SMmfHeui+p
XUxslheW5a6fSSN9mo8AfUig66qOxUhLSXdSNcBTa+1Udpd6Wo/qdW0d+irnCVsI
gp/TQBrS4oIRyZcBQXPv5FhiKq8K9QOLS2UB8FHwvDF77ZojlFhlFVZEsNuBDz4o
Yq4/zBgjmpKKxWS6B2JHSFXfakM23g4pXiAOIBQxSOWe66baXDvixEnvj9a+CW0d
/Ih4wJMhEmpouxbdAOve6Filstr2i0fVtSKElouNgGWYj5wHbdG4brl5TQVFWuMW
hoMdhp0EeFdVbTmuGySBKEKlq1zrVHAkhRqL6DD3ylfbnzmD7/IyV4/DO/cIIDJ2
7zW1jOoSnAneqju0ay8PbkpbiiXUlHPdI9wmpVF8dCTA+0AEKgZLIFY8g2NWcSp+
CWN0jkgjUEmlTvDTxfgpIJxBJ1JcGYoKjSIkVUTWCZb3TWOVR2MvQqNekQn2EfXn
3n96HpGisCxU4G6xU5eQDW0P4wcGsd7qqpd/1Y/J+tHuNwdSgiTLAq5+hUr/BhI5
OPhPbVCbuUtoOB59rDx3INcgmXlAqnzmAgeo1zyi7bZzxV8mTAUzc8cwC3gYMydV
8v8Vo6vLvRBY67iODrY0+xxpVxXjD6yOv+/Y3ATsVmq6PZ9xgiAPC0E0QyvjVF3O
V2thvjpQrpiFrkvIZaulgJY4TKW7POLPqGagWCj8i0kGwSWOC+f0pRldwjR9X6cT
9+Wv2/20dQkKZ7LubFVhyWsYvkQdIRLgeio0pgpijgaSIvoZgpZ4AR2Tx/IIfe7N
sag2lZ+khTEvC2RvtHSoI0Kp1Dd03IQQhzpQeFPItxcQqYwJfOeXw8P9XcRVFTCd
ebn4ZRALrZNFFIEc+67ze6cizACCwsUndmiaUZ3coRcDhmfjpKaqqH3fa6UTdByG
5TifV+1ohZoGQj+vdyvS1hQLY2iN6Bn9VzfgAtb40LZtQ5abzKD0OOr+m1tg3lpD
NlRgUDYNHSrgzJqTBDiqXyE/yecXJi+mK9ly3wzLUb1S6ok5ywzLcA0GIR8/JPnz
xhLedOD8kMtQOV8EvlYqOuUVrEEGGxB7fYPqje9fSwxSdYPwuuaI+aJy1mZTW4sO
B8wD0YvbeFhNzStHqMC/oBO7PPFOxT8t5NU8xKMzdsLkCj41I+ahXXcFZtJspDJz
lUPalyDCCBkaSXzGBdbEiWyqJE8fq1sqmSrpyJYChHCNkVPRxhkB8KundkvvsfXJ
Cr924QepCHTenPnfJHJdlUhEoBRCi68uLyRaGXHNZs9Y6mpQHU2GPefeW3S/6sU1
NApAvcdDhPQ+bhv+VgRQfW3sBt7TzvCj7jnTkNZzUsUPT4fuaq791gUIWbg0L6CQ
VPgeCpWdW0mVla1Mup5BFaF90XgxcYnxY3mNluK5sEgyxKy/0PdkQoVdHoz0lLUp
VDR2QLY+v4REKNpUkb30oJAriLIJdl4oiSUWtJgijV0YxZGg8I/eRsPIIOTZrs2G
Z0No71QQIGPXM5cCM7YEAoeHFIy+bd5Rx2shxstje2d7StttkZvSkoIG3cc5qx/c
mD/EXNoRGLAMmmThG/OWLrUd1Qszi4mHSnABDYBUF2ZIeSDGpwCM3oAjUFDY/aB7
OOYACiSETIavW+W414JAchHKQdPPRChd4s1TtrmSGnCgOjUQIum+AlfJhflM+pWr
jn6YSNeWn7xTY9di9pH6hko8rMSN+rvIZwMa6wdUY6neTS+aLpghMAbrsct3YF0B
c2AswjILiWDW/javJTzIVeinB/ICwU1LEbc/K++vccUkE7bBQdwDUHC+Q7jkjzyK
V+a3ERoTDklo5kOS/fWmpAmd2eqikm3m5WV7fzt/tXzYEutk+VA+oP9Ee9hknZL3
q8M61MkvsuWiIlY5l4W0amN1A4nCuIgxQftT0e+fpAe0TMNzXRBSRZvc+maKhvHB
3xFt/El6ny332lep2YNJnjbJ6M/zqiICyqXg2+D66Q5yKGWYRR/pe5DIdgRk1Z9f
A3srNlRNdVf70UTx2gCXIRmgyLgd+7P2MrewwnAMeL5rxkAMBobrpsUMolchWa0R
Jh44jwr7xt925gRl8iwLTQp3fXjSDB0J8EwfuBtBpVd2yxsvB/EWK2+x+gQs4tcA
zwVXUVXLWjzUCkSOnMU/pm0HDkj1KVFOl0VjE85FxfYrOcSrwkbTAUclvPoLzqMq
R9jTuYTC3f/hJwx7Jpr2C4G/PCFGgwQmjuem/CXdAcYMHHCtnW4y8zySaSybiaKp
MlgTQ68doWygRgDBVFgH0NILdhpTzuSrQLVs7Y9x5R91GkoO1KhHGfjZwh2Smv8b
hveNzVXuu78PDa9Ul7Ib7Sc7M5hIsYc0Waemp4LpU6jGb+O6IjFkJVQANzo/J8VX
YAoTmb1xXkPz4ydhL25V7vfA5SnpdGq2YiEGzqk5F4LFjADp+uWphphl4QN7eVcd
lTDDyJGKq7CDRkmEH5JG+98qWVO0PHnxq+ISXYraWIqWT1tp3Ztkx+TbrnpZMNaJ
eE1fTmrXQqIPg9U/E5Xw5IFdNYjkAywSDEawfKXXuGo7Owq4JACgyR7UZenfz8Mk
MPXN4ClVvETvwnAyho6t9u6zLpSaPdVaUUS2gd3k0TGYTVeqyWeKR7EQU7t0IV7T
UZHvSqAdKp9GqHoh7hVVqz41Xf7EytO4hNdGdzVX5NOSG1fYzbRwh1Zwh52ja9ln
zz7UAX2HmgzdtsgvDjRGBEX3yWgjRAmqz5S27dROnC7DOViLr2puWVotxswC2h6s
jboCx8HEgOPYG3AAiFUyH+UDbMUxeMo/oObD0FvITq4j4VaKJu7EYDR5mgkVjcAq
+rIgtSV28pa2Hlg8n7JX3MM3CwQBdGp56kgbeJM7uEslEyfWhdLxT82r3EGV1Xy+
V+JQlXqq+5L7tddtz4rPDNId8dTAP8UROHJ5Z1+EJF/ZXrr/W17k+ZHrYbC5DqU5
BLsWoqWA2ySCD875uh9E5DpzfGnhvVVW4kvcxHocRmMv35GiaRJUfEsfr/7TACAJ
JjL5VeUoIrt6mdwSMun4mVlCBg5+ETZ2vH2UTPFjO1SiXljNc9ROwfAh6aJ+G0cR
8Tdp9jNykjGl9vdO7nlYZ1jgVY4KRFU7qy9eOMYeOK77ENxrkS1jlzj2h1XZeZ75
QesLz5ckOtLfxL5LfaTBFEqz2PoLK8a+UdAmcVBISrBmsqwHOD7E9JC98KOhnUhg
UI6c7vvrqVsZ/a0RtRQ4D0istO6l6h6JmgoTlaWhLYQkwMjxsNWcT8qG1UVHUs37
i0XX7r8kqnTOWHaAnB+VB3y0OJqXOerqBjbpxFTaHQfcZhTj+zozD4r1QJMNnDJW
ISRt/VyXQH8SAjAgnnAy1HZYLWndkwcJO77MULetBRuJd8WshfupgNmBy6sukKLL
vfzljvINAR4jSnmZyJT7p+S8k5s0/NS2Vp4IeqKLSxR8FVmHX4m0n9KM14z4+9hs
RHGi6yXdBPIYl7iBDl2KY8CJ4V9SY+yyX7GSnhChKr6vqXTLpQGbYY9I+28q2bAE
rQQDGBCkEMzgLqoJvPXd21vHuwHREtM2ZhQavJj8MJEyu7vhqsSKJ8h68PohHH20
Lghr9SzsR8Vh/hxyEwE/UPKwUJViD0rsRmMT1bi7erPBjq4nuwJvQcHjP4DO7uJQ
gAi+cvKvmjQ39I12uYicXY/L+9y7hvHbc4v0pLGvwnUn1tGzBOSxLULnfCTeDIw/
/K1+kXVW9pxGRKcY4VLH6BPlaCzYW3d1Oo/Qkmxocw1r5LZXU/Ppnq7TdHYckyO2
IirTrIEwCZD3LMFXITOJMNNKzbgy1mFHiWn+oE3DTk8jtoPW4XuBQ7IAQeHGrOST
JmfzBoc4kRNvj/SjoF6O2jvHOf3ZUblGHq7zoABC3EpGySjKIdm1PK4fp2iP6H53
9AwUO84G2NRX2NnCvyMOROp7juKhpH15XFv+9HaQQzGlC/VKJfv2BBlZ7EqYDDKn
sCuseqk4NEcdnk5chQ5xzKU99oRGmXaCY59r4H4wfFUccXTHYyt7xZxlsNz7PbvX
1QiotEvl2uP+uIcZ8By2mqLvDtPWGnx/GOHVXTapfdiXO1b5jOVxn6nGvpajXsbw
xWeTeNXoglsT+7tfR0lV6fzSDfZ0i+HjCsB05sNYVwNe3EL2SDUgivTuRv44KjBL
WhdFvwPdGVQeJQu788ay83shEOn2pel+y0RzsHLkZwh7h8rdGenSQY6Twlzx6xjF
yKtz4OP1agDji0KRBHWFQE79Zfzv5Y3HiKaoRZq6puAnKZj9varOZfsiouHYfLDj
8MtKZAGprfvqcxDolADI+mBaKFJ7s8lp7dqAeUoejjObViHRBWGDjrZEeSjHN/vq
RF/poP6iKRY9m4IiNo21onoUoZphhQeGc98ok5dc0yoOpad20uy8UY3RpQUHuRrS
5zCF+1K2TdfXvSyoE8ArF37PIcayc70Elw9OL3YyIb+fJSLg8DSl2M7/LgOfNB1q
B/t8Q/8Ycg0R+jw7EPuZcxtUFr42S8spotrZ3Xa/fCY042NkRlFmTlidVeD97lVE
9QASV34/ALRrOV4ukl5C573HivJxKN9g9dvV8yT2XqqDZp6Pv0rxBBwBmlDmIsUD
vH5+5jYEg7jxz/mbRrL+2/P04JM82ZJ5pxecfGzZeVLH2Ugb+46TGIna1Lfh6Y8U
0lOkHvoo3VV3WgbjykEwQOf4dMKWUCwIQUjx92IEiltp4WBJrXhQ9HJZuJvcv3U6
zUt61vj6JFvaYdj8s/SPB+F1ZCU5M3TCu2zxYj7f7TxfJ+MKOEvlUdGt9FpeygkZ
YocgydEmL4v2kaoHdpmFgdseGrTe20b5VdzVNHx3tq1+fG9hxEyAqdouXx+Th6so
By1Wya3igPzd9OtVdxWvX9lC7JkwaqDjDY3B0B+Zb1pyxujEtUOsIqVGki3H/S1J
Kuwcxotmx5ign1W/jYP/4PxK791INTDYrqpMAjWCCCo/ZDZWbW21Oo0qvsC4tTa+
jbyPa6RA1ip10s0wp8LSSmxt8mKL6XVZvWBVNrLJPKdVtElEd0WEBHj4Wvw29Qa1
ejboOPgl5+9jUxgX4MMFjgU+mVy+sTdy/lRGRyXkWHX/chU7b/IwdH2xhb2FPdD0
HKuHWgiw7Cttw6VMrnoXY6jRIcU2K5gXxEWvlww1uDkVEMr5Ee2AsxoC8Z6VFiUd
XSV+NlJisBEdmIS7bt6Yg8Lic69iyA2beO1LlRNLpdurmBgX8W5aveeT5gAYFb9V
n6H5M4YMcDWLIbz0cStUSnKAhL4rHMKY6bLXrgi2eVtZpdkVMDX/nH6SPD3xLetY
du6wKIs2JNd0JZUP63wya8thrFn6h4YD1h0nJP8u6ZtKav+B4949AO84tM+Zczvn
X9Plzdz2wQI69QBjbO6NyH/XHFhapiJzY1mP+33fv0PflxqnrlcCSLmTBn9FpGwu
99jX5gVnPYPwYamZ2vQWWlaZYiBcrHDeuLOQC2i5k8hDDdUdxLXH7G5kzGdqlRvC
MSR91bdK0drDG4T2LVSEqgOxL3rinRIyw3xherqQN93wpF8t39fm1B23vUzz1agS
5lG1EYSO9N5EKHhOxr3TumgRuZTkPZk5rZ1VMqWI5Vl3sh6FJdTxInPobSFqzjM2
K8okvMp7OmHDS/VqtY6d/5ybGqD4zECTkSJInV0ARCmZV1BDU0vcCw50a9a/Tr9M
XFVHHfxzI70bo9+0Tay9qMyp1n69yEgw8whecpWy6o6rHt48KPEYBT8JYLSJ5Llc
93yuYrNIAykxlMDiWA23VpQle39V7e67iIxf8oOfXwSAofk8z2rr9ne2euafwHTY
nWTR0t0o5e71eJvHDombar9sPHFmD/aGqR+Gur4LRhg8mQEsngzl3ZWVcbh7YIYp
sbEJ50gvFYlIvHu4gbtfUohLS35jmbUnwuOew6ygodi3xNXFk+2Ua2cr5ohJ/3+4
12hEHSiK6rBfXAW2FQcmiBGvStLrcq9bNOiIDAdWMAjyWGxLf246H0xroX7PN1jp
pAYiHaTg6dg2kc1Slix1Ki+Muc9MGGeHoJD10BtWab1QV1EScx8mOY69inwBpLi5
dSOOxqHDuHX39BfB98hvNW5dQWNHFIAp9RnjMibcPdF2ubujfN+6DjB8nRZ2QEMs
imWxKpJ5b0K8hfILCrPYP9lB5zSxGtFnCV/4TS074qwZAddSPaR6DCzMOXpCHJXp
Nv9e3GvXJ3XFk7a9SCw6gnNtpvEIcS5QQB8LtPOuWcmGiDvTrS48KsLrsdt8Wtcw
i8C4VcuqanBnAtaYtcLHZWlUSa4wyx0luvYD6coH1n833niWuwZ7TqbuTI4GtnGn
jrKuQHMqYIWiOq6v+qF0zrurBg3wbe909qEEGbowpGleffARIE3cnqLvQ5iPeVXY
VPXqweQc7XAKzwTOXxZ+iNAywl5cAYnB6xWDin+jte0czvd553s88szqR0F/euD1
8dxyimxdJQmAtkZz+WUeENUpiJvjpWZy0bIc75YEZiX0cCpbLbKgybjdR811v4Af
S0eMuoYMpScAMkWuY89Fw1a5Z76/r9l8xFmiAgeQOZpDXOQ8XKXIIztNUMLXFAOi
27quTj4CsUlTNZZeMcIctRidf84MfJGh3L3OqqqmtQVfj1vasW0dnfwtGoj7skvI
iP3s9NlG485b7JRpt3+8jkRZ+gVRUlUa4zKpJlSv6VCf0eVKfa8QGxhvI95W5Y5e
/xwRvGTMRhmmFfzdxHZ3D+rgl34DrytZcjTSQN/EZnbY/CEXZPhoa3dmmRBBY7zE
RAgrZ5bwXEG0icKpPc0N3kOgf/qD0gYgtqVDLoXYbI5xcKwicF9M06FroS89r30Y
wi03vLSM9AEK4PwN0Ihv+s6cdfDIdji76a4NHY3fBNUKWMcZ3+1p3iIyEnuaevI3
ZCygk8n4QUyIcn+DzGmL9qHfMIiDWC5JDdDIsxNGkOjv9pbxRKw6OGuSE2jXo39c
BCSnk4x20h1rF5VogNsG5l3z6FAMUKXF0aa9qKEzCALICJIIZBhrGfahpztvydHy
tqP9qBeqMjTqD01+p4Ymw4oL3QBC13oX88m/vq6ltz4udPiZV1/rbhl5VHGA5Fhs
hn1GvaMRGT5haI6IIqujNiujHkohggpX+jthIrtUy/jSA/ACRzP1kMLTMZo6gZN/
/DWElXiG6kb0GE2tZ0bBYHG8pK/UoHXkwobMyT0Tn2JuTWCdstPuUwn9ebSjh2tI
7qB7/YveR7VWvc/bYuOvoJtZKbmNGu7TlfOF5gmlQwJdA9wkSMnwDNAjDBCn0Shp
1PS++3ccRu/Bvvi2Ieo468Xekp9vxLi+i5aNabjMRskFUidDYysGW1aAGIfMw/0G
rg6fFX3E6fCxu0JLyos1YpR2HQbNYwC6jzDABh4qIVjB2A7FzvLDLAMRKwIU3Pjw
H0HW/AeusC3pk6KVGx71dDOqIH338qqw/KkWrLHdK/Z2/eHMcRCTus+c05hfSSO6
a6Dgm2i1g4t9SlZMb4eXwgJ32lmVBd21H8LZO/UM+QuOJz11b9M3daFmlMaeZ+0p
sSjuVUJNBi7PUSEswKxdVO2qGjKGv02wDQ9jU9l0+vTd/s/R8MBLdnQTFy3AHPxm
anTUJPjSNrJ24d45+p+sQCvTv//o7dQjarphQ1zFVxnie5XcAbHyp5lMfLyWegCl
5VQ4LCYTi6ga8+rzuwItLEXW2vyS6orSPZvnjdKZRUl4ATAskk2Me6FhEybYixq+
R9QS8LJMckS3v7hIw6Qspkc488cJrYT+6O4MbJk/tkjnxX0zTSqAePAhidEaww24
4bsPUkj8bpuFnFWt1qGTrmp9FHwacODom8c5aK1U3u5K2aCN3GVyuP718dmVi8FX
TO+ZbmHqvIhF92cb6aHv38LarFvhKtDyvFBP5C7inLdAGYAeafftQaoneA8h3hyi
NaKAYkpkARJdD4jBNam+2vWUZy7U4sXbLib74obGiE3y8ANEgIwHvB5271uYXHoq
Bro9Q++U1q2O5SMb/BPhCdRGvVHflw7+00s09wZUPJCQDSyZiMpqZPcsaGpcYue3
MD1XIjixOwBcdIUyrfwctJ8N6kOU3o9o6vngxACZUJZ/vVdhcEynyjgCmt41Thd6
hVmuM2Xu4Ef3AAAfJNtIkWDCZ98/eDOOSS+TXzo93NlkSe1iVACghjXPNcz0zxcd
/DSKr7yGWlALRP6/mReFAY4PwXHhll8/zCmFWkzEEalEFUjCn+bOhQJpLccpmi0P
yc/YeES/dj2Cqy060sgyXdfYn6IGIDj9Wo3TqEJEaoVFnrEo3n/JmoI9x1/DmltT
mmD1YiqO/xIGA4hUEyCC4PUPCfOKLbDXs169jJ8Q7Nt7uw57O0iuag4TCTuoOCAx
GuLZnu8ZMk6kh599RlxkrPHEYnPEtKIjDqYmCgC4KeBlZI09XJAWXKLmC6ZXKaEl
pfuxjU1Mj47Zw+6Uv1OgyEYVkFgrhLuxs6ypAZRmXwPFTDf3D72C0dOhKVBHf4gv
NoFfQ268j37HkunpBHI7W9kAY3yb7wUfxSgv40ONdcXnCCdPLrTC+Xn1ZmNb52Le
vBJ575WchE7/t5LdwVv43e/QuiAjrMyNpuAOYbTttUEHlHqqBMnqaCz6LWUDUeox
/PZJmj3yWv7YrXV338qpAWTMN3sYnmCiHRgg717bAt0BGnC74m5Wc4TNV969K9X/
dBEeLeb9IRRP5U5bY71fScPDXPexL0wG4WXlkfdnks5hCNwTPBhpoM2hPzakI8vU
Mr9voBKrdqzy4ABuKYDOU/uqyn9JI19+npGc6ZhE7V6iZJKE/9haL/XYdW16A/FY
o9II94CQ1/OINJQ4s67nLE8ooVoYgOIZHG5EsUzVFtoRVaOy2JcWocMXPB9Cz2Tn
Y4V1r5Uk4TsTNDQzpS5Ge5Xe+kSK7zSJFbsMVabQfpIiJ+Zw8sdER1RvvyQP9iup
l5BIODlFpBIX2xFbBu2DIvA/YfE8aQA1dKDc2bZpoGhave3TOL6YBnyCET0P6Vz+
HqZiOld8An907oG7U2jC0JYx11Z59KJY+QQuMpTiQH/AouEwTNdAf4EbwBTA9nC2
E8WynECK019z5XXXweT4Phv8HutVfwg4TPtFOv9QivDYynbskYYfXXhj+reJPDqo
0W9yYoJMIqF/pJu3N+vaiJ4b7Bc3OLaQvomeANXG0MxaLLhu8GN7D0nPTiMA5u4K
jfvKbUqfXn2/l3j9TLMCRBTAAlLeN5/s9/Cc9ALsa3/MvSDVjeyxrVgTAuwBGEfd
DLPuBxUnEjRm4SONzMKVXB34/hLKiJRCWVVz7gMvNjWK5YyDbA0htX4bwDi/Jh0C
EyCc4/hcf4FvobWJ5uYn1QqFe0TOQzRlNdi6Jy/PkEyVspDAI4XarWDbpckJyV+2
oHKeggcj/Ad7pRNBdbHdNs6sf55JrOrOUI246cYzgk5cOz+x9LygSiOLihw0iDaa
/uJAqkvWZJDunNvsK38luBzVClJqQfo8Nii/0Gvi6aL9Bizgeat4Z4TwnxKJpFB5
3YEAV7UXYJg/Fxb0AVsH9vj+NAPMuJw20Y2skAtV8koz/41TFxz1qOsvJ3nyZ60V
uRi7s/U4rmIIeMWvdeF2p0HZDhwgebqhku3AZqYFC+JbKZdxpXRcTUKjsQUYNoAv
jQeVC27wfZZLr3O/iRGHQCGLLqTSGilQfFvwgRwGzJ61TQ45GSaTN3jL8XmfyVOk
L172XOa7Bw5n8RcBZ0n/P92rpsMxHmiVkHwLSpKmaKfjZTCilo4+LJTnWJBW5Dln
Jq2w0x6RuxVuFISPrZ+1QsRSVyN1oZ0nP6rjr2gGHURB431uBwi5SxCCX0lkjISf
RKEEZSrx2PevQ4mLGalnOCyyhV+S0BdWWPMbfKbiHxGkOUw+TnRSFII280X4+qI3
4nbZ7pVkD4nCP72K3zU5pav5JWbcvqzf1zQpOXGGSXrPU9KDYG/VCIcbN1e3PJGH
/noN3nD65aGj9YPLD7zzWHQ1dXdBikDrhyrH/lBpdXfYfSd83z8r+50QpBZt1d2N
YclMfaS0azZyFZ8erCH2y+OBTsukb+9P3k7k2IB4umV4YOdmRSo73SKSdP1LgtRd
zsavXa3WOMkij6YJqnWmA94HTNjEKApRvZ45mT6ToNMrXX0RUHTaAhgXSIJwEpVl
x5CLc0A9TPZJG5eWPeqZj8dS6fgx0lWgc6iUE7WrDAUopKvd6EcBUVe/5Lx9KH1h
M1xaskWvGqaTefYdi2palF2wB0rAb8xu/jxKCU8rrliUwf1URYKGBBJfGuZV6zQy
16bVyH5jyaFTZ4nEuu/N94z0CMmvFUFs2OQQMSuf6/T4UAq7KI5B7IwsgMJokNVi
SBh5uUqILRp0nhYlI7TlEcPk2mhzPCURBjhaKPRopx3LzPhjpwYHH48n0n58mKAC
oThmmQnoStA4xXGsi8SGXFUbTgdRyiTZD1aE8cBukHXi6PGEug7asZyUUtxrYikY
PXz4HLQQFlzDL+9FuR1oFR5D2ES8v1Lf6RT8chDa0/6+BqXeu1XJJ3LXLhOv9Y+L
xSdPA0OLs835iyezQghIGk6OI6XRfXTjl/8aEzQxINun0Qu/ROrZIbumrHc9ZJ5m
T2WZngaqM9Ep4ZfxqPlKPcLjzP68xrNSM79sR/V0XlWzsJlBhi1BiHVk3PSMT6Z9
x0Jq4j3BOn38OLWctiqtPstT2L9J7lTMbFt04AhJgyLL9NtZRm5x7EleN7dCIsJP
HgZuq7pq011hkvDy1RJIHRty9EC2VoB2uks44C+oniHTg5yxj7A0TQQISqiTGSW0
nzsoqF74DdVapyKjArn8AwDWxt/PMzEU+PZnkacFFNA5WnjAh0By9jVp8smkUFpi
xmh2s0l0NNxb6o4WOlaT16ZGFnM38lMsSf0JAEcQzbDNXSz9cimry4SFrJ4D7uuj
ajwsQH4irHoLr9kk77Bs9XNn6e7iSFpLrmXANIbkClNJDogVT9CRN+Wc5BtZ3cMX
WYiQdkrTsn5yHodVFOlztrH4iooz83+c63ak4qPYrjfqX+zWNWUi6NMBlXTUTWWU
Ve2r8xmNyntk/+Rlw55WTzen0Ph5O5Mbj2bywwhsb2KzZbtY4XLgORKWYzT08jx/
0QfCqt0xHMHmFEG3ZmqFFFBKwlJCjHXKbUzqROagcTkZHnRyPZTcJa7XDl9WDicu
v/LLI9TFj2laB+q96wnCvruZoJWfQ4+BGR0ZReAbDhrwSToxIitFpD1iq7XWihNK
wclJtjEaXlrjP19kfGKrcR2V86AY+xuULLjCn1LcKgIXZbMpruJ16xHOXwbZkNhh
1nzs+3USZBzwShesXDy5uk+eXb5bJ8mcnACtRd6595POj4LknLLp5t99LyqB9V+4
2hgH3Zx3utaRHab0a2uQyZ3JLHwL4FPUrlcNrRT55G7Qjpb0Bkr053B3j4Stw+6o
RaFpNN6ZdjYi7koIAWwVjvb2DRAxB4+k04jJ2j1g4f+appezAddtOKjIE+o04mF3
b+NRweh92X3Lu8ppPhllknsY4QWrRaS/k/yIlhe4c/c0Qw9QpqJgRBGoB0TukuRZ
gi7MV4Jug87wHC03u1uWJLUvpkkj+nfDpuIVhlSNwfiDommw8LiMtd4mHuDsUhfR
qG+IyK1Wqt3ZLcXkvK7MzGplqLHm0qKq+vYsCCOGPegvkNnD7qPZuv71rtNko0pD
vS3EOw1bJj+Mj/zTH/0N9blortol/PzkzP2Ps0ejdtil5Ax91du1xwdIkmrGIt0+
dfEYpVo7nxewNc7qaru4o4TsiV0pkLU8G09hMtzDYh4nIB+YIAdHVyHALNTPwV7T
dJS6bIWcn04w0naL1j2eo1O3zdosK5R9y8XEsrPbr77dL0SxJudEaQCR6rSEDFl4
qXJUTlBmerFcSDHI67bNnuKdjiRaeqDhScU4aj72i0/t/3Vf4sQ1MmZLE4BoiN00
5NbX4K9RqMD4rOn9hKAC/gSZ6YZ+7vxvr6x1RJoJQB48TSd8P17FasRIpOTueSQA
dkvU0bOBcZMkKDZFUfOs10V+fWboQrHco1xQNbqwTlG4EohcONjOmJmN6ZanPtMj
S2gmmrQPo+RlE7G914cCptGkvmge4ntUmh9dMIv56YR/fVbE0t4TsQaJLlmkfbpX
9/2GvCLSuRLlFp4VAkgPlLyKgxfw/ENGOEYpVi8u9DhkmHRFL+2uPvObn9ulmwhc
TmzAYqMdUNWTRwCDnyvhQX6T/3yYGwJY+nEUS8jm/zXL/8TQ+Gu+MQiy54pypelk
AhneK142I3kBXgMizeeNDrzxjxrchtiWtQ9PD++MaTDX3gcOJHdCpAht33fUnvwj
wIbd99NZvkh9jo7gdJBX+4vTWJQhVffijFWrph4VflwMDkfH9d1PUE9SdDNUB9cO
4yYGmfBEJKGWMKniEXX2vOKoImy4qVYzAKn+4SKF2VXoT3AIXJFoVFHKN0vAgkvQ
kofJh3t+PhnIG4TLwyax00C5yIjWiKsoAhULsnh9Cx0PHnhn9pbFZSTCtTs1FzX8
zSKNcXf3B58A1VVQpIznyw+C8BQqGrA0sQEqBvLqfVRxZ6TqrZ75biri9MFZw2b+
jkcsC3i/vHNVVNfBstZwc/8B7hvytiojYq/T4MQ2cnojRgH2JJJbYK6IFFLbfTV0
rRDbnPcAyLbdCzc3BedzEOy6ickfkEwLguR/Ld2aXDoO+0ht3xH/eFupGzhJWED7
QE/suOU6XI4qWlklRf3KgfwTY3xtLcWojkJZHf0whSSyXzxITpiS/MOClUEOOUh/
v0MeczhY7+jWAsM4OeBfzFWGs0zrMI0KVbWw2ObMiRmn1hbiuYG9llSVXeSqMrhB
I1FEwdcqcymJGmEX/QaT4emCoCxo6MTyqebApks73l8VsKgP0BEHmSYCUEhSVXYD
J1wHYPz8OZRngN87EaytY8O3vmcI7GZCkYORcXdHhKwISDYTDW/Bg0FtqYkSKGa9
pE//kZl4iFDUEvl6NbxhRx+pkdMhowavz9Nr9rXDxJEVYCgl5HgsUXyRJFIWXSbZ
2YKRPD3xIMDFr+OfMqlBR7/ODh+epk/x6v1g/RUksqWjXzk5v352/EFvyTbeqGE6
u6Ak4tRH04arm0q4pV54KQa/yIhHLzDadZbhQwdIjLxX9QAD+5nSjXRjsROVX02X
378LfdROuWIzp6ntHd3+UHm5jExm63CgY6VB6b9numvTIR5L8WqZgZcD05Cz3MW5
GJ90YBiFIlS+GNY/xWjQugTvxW11VYhzmQ637NFc8IxxrVpZ27WK4XlIGM9h/YGU
QNTgsVJlbOIYYGgGBa73XEbBKKxt7XTgfuLNk3wqM+BY8ac6APtPC7waaRKV+16l
8hXzknrluBpobfe3ZGyDzrJplXkz1ejoCNKmWz1Lz6Zqldb7/kpu9z3o6LjIQFQp
kbjxS1HOEslSYHArdJPxYcpSVz+12jrbg1ksgMaRWHRgFcZ66ebabI7/5mBZxQ+a
A2nZlBppTRpE7qn6Uk3TIB5UBo7VVVfHKzbhvuzWYVnGKm7Y+XvTHJriHiz+tL32
j5DdIidPsdFs7rxpWm/YhfSO8TobMZrOin8ZSbOEWtQ1Io2bUVhiUtNHFrIkSWuT
ESrgNhwB0h2AtyCtr6ckyFhv7Nxgo3mAFYcPBMCQt+HLxBFumxX8VWVDvNoWu6ru
kcrFMXk7asI1vEtzFFEgtmdkWuZEl2ZNn+Vwm3VpmN3e2bA2m9HLNsRYrqD5QStP
mlM4v8aC1MsP7GlASt1FIBg2bNOcgBVhAVmgLqnlIM49b0256Q3azNtZ5kiwSoV8
/OrH28q2Szf5FoFocyPEEGaCMnbUPPnouDBFWvEWthYRY3cpzLBB3f7+D/X05E7x
Ap78ZkIiIRFGQbiM9nSp/O6R+NjCn6BxwKjwEnBw2P1dJ9DfiCAmujdHbUC2Oaux
9s3/79msXn4mtJ1uG1As4frbb9t90zSHG7Hg+cXghzDkVKHbcDZPuetQTyPGOtDr
sFDTvNw2dzxG2+KPoHfoP1gPbvByRaq2TemZp+5upXTYCWX1YOtQ1kOW4AEjwHXC
fE9aXqB2WDRc1rzvhVnX3bCcIBAxjRt6kAxrwn3SYkF5pPJccLOXYm4HyGLPriR/
yVb+CLBxRRe3dWGX+UIb0lJv02TmKpO9U2SwiHdGXexL6N4ExhUh/qTI/HPyhAy4
aYaGEC37oIP8ntvKHEcxSV67ze7tIdDh/3zCUdXMak6nxHB2R8LaP7tiVDnwkXKt
CTVgiEdc4xpSW3k7fxpc19upIv9h479M2cOcNJJXCFYWj/PfhIlBXwc1Wpdz34Kk
cH583EDLWte4T87FYQ0EQXAPL+PA9UjPg0tnpWwFXAMcLhqrLYn3wLm1cgaL5NXS
IgzD4cHmFkxfmKjRzPqI6bEf1Qqu+KWwRtW4pJ8IOza1yMsQb3qadWHhDslktFPO
Z68t5xbfYz4uiguJQN8yhRlWXFZ2HxLeibcwTNT9WUk0AxXhI1GCh0+OqYIiQDda
nprOIqNJCphSJVlobB6ffsjEOzSV9ZczsiZdmx2jMETr9J3yl39CiWivvUqOcxw3
7F0711AlVV+bTdcNkYlIMb1VF1yZZ/dDyEVjx5khIBrbumaD2on4iscEJgtlKZPW
cujFKat5hUqCPir9W3fS5aI+p00jEPujhT1P6+1yYNBMDeiF+uKxTMv9G4PDENkD
kIz2KPYhL/OqHEyfoGXlkTuEHuOSQmTS0NT7a38kWndkPTu5rERQcD+9cOZHhCeX
BxmoZJZSaa3o35SFH4VkQoqLNdDzZTT1PxXbisFZlUxxJ6Aq+A01P4h+TT1NbX0Q
oUXCrco3dsFbSVFOffAx1J4lmgNw2mv2pq2KD42s5u3NdrujWxw+sAYSfAPRhYFj
kZln812KhhNKwQ/Bsp4ypJUe/MwjrH/9B+L0Kpn3IVh5hSPb+/7uxWefIhkCzten
eZIROg2TiRd1J7bOx6pBtX1tDXvlfUBehuH957W5BW9Lkw0chZOa6unM2yxqE8Ap
tZOPK+wzhAWb3odPMzLJblUKfCjfpW3C2VYrXNW9u7LE0XGIcYvFlonkDDOBFPJY
iKAYUzbkDAxBzZ5x54/kiGZHQcd3iON44OhhVsgsDlcNxLcKojuQh6MXXiHJQAzZ
2+gjp0fk6Rnk5PhrryluSGKoyMB2CV7N1zPlWxOGWMVve37EFag6An4oQstnLbqf
tiBWkmnpClRZNqypkAdXfRilKrfR5miCUmygOo6kXNdCk4rlFay8VV5xfaMkoEp6
4B4LjNlvN8RvsOAd3KRtpVCfkOwuClBw9eOOD6xW7bpZTzCwOfqrZolCPp0rHzq8
izkk2iPZgfqo67W7sM8/vKXlfmkspW+sj7iczDkKusHuhD3cp8KZ82A6/ssemdhy
dnYSEjiKGvw/WKySFFIrK4u8IkGlDVbwY6rHfosA+VkXDO8PPHxHqqZik7AZ5kxh
xjVj1iWzWpjynHKHs2GvG7/b/gljkXj6lEQclShuSwGK+JQzsKzH5DvtYJJYYUHl
I13pTjj4f8JlKbZ1JpimTKczLLv3X/+VoHzvCs7COImZTJwflloJOp9xKzF0bZdb
Mq7pu48yYamPvicSf71eXnz/Q83m8EztKZfkFE6lPw0rWqa+9zRxCc25zPk/Q2iQ
s2It/A8Ihc/HWbTGZLpoknrC+lywGxj+7Knjtc4LrCs/tAXQNJQcfBqrKkROKsAD
PXzvRfkBDVspV6d3+0NYt/PIiYVQB9OoTUh4RL2x0RM6iOmhKZrIfjXcb83+cv3N
QsNsnd5js94L9yG+M8OB2wdDYIcIHOhQGV6FAzIVdxmNPHeaihDDus/7gW1k9WEe
M1G/15zUPeKFoEq+BGhxnYpcGTj6M0tIzEGPWRBJIoCu/2uy+UVcLbFblZV+ZLfD
oN3GOVDsQvj3hyr1AY9zjmIOgCBrRV3i7nBy6x5rYuC5Z1oJ3A3jhwsAaNrCpiaw
9kvFXukk3gfpoVVrD3eZajhJFuuX0u8liqSrBubuMBRJYUrnmFeWH5ENla60SwRU
EVNMjJtCojqtwjv5MK43Vpr/HTfLud68GTlfkCNMubTlplr0ogWO761QcIxeg8cK
NxSWF6w/vwV8rL9xhvWRcivFu8cX9iNoXHN5T1e7k0dTS1Rk3vOAS4Hma3gkgRkx
FZ25V8A0SZcgzKRlL+Dz2Z0Y+k3FJNBJdDRWZW6VCfNrHA6LZPdKrGyqQMhDTE41
Cc9BWl8H+xNriSsU5mkCs2xQmzdrx55iozVjWVhC4kU3xMscliNQBcDi16N4JJDF
eur0Mc5iy9iW7jzgvT66ACmwDhgZrfvr1AVfwyW80YLmGQMqVJjarP4CBorYLeig
H6epmhhLapUQWwn9sNgWhbGby6M72H4d9FR5l2ODP6LihpolTgC7HenHDj102M0C
z+mOg3z0zM+n+RQ4qFwIX1TuFDRTMBDpGkYdt8ico/+tJu4PmahTMN5swum/1IHm
6cj4pKwyalsyOYf/ISHlD9dkZfCgDWzPv7f+epMs++DtC6030FCPwf2jn3Mm8MS5
v0FUxCZfFBPD1frLsCcSi/wcXPPRhZju7SQ1f4W1LsoovPgPTdX9pRo1jqX3mzZX
kr0LcqbT4L5UvEuj56gUKk5hPiYgNc+3iC1EpXn20IDjQhAn2t1HFJKvOVQ+jBN+
lY6gPW6YYrtlcjnwjet9VcZMeeE50lTGu2ElthoeNEHiUoNXHQHdxV5DMDtG8L0Q
PAkwlrzm1c0PGWbhVuGHcMZXdxbwAknqyEQWdyiVyHYQaJGx2k5yRGg/Nfh8FA+G
5r4iFBLBIntv5Ke7RZZWteeJzEUMczjsXCSYcomYLnRrdPdbS8UInH0y9hPpi8cv
VyvxQQVQod9A+Ewy2BmqWf7kAVV1uQP49sx5WcPayW1+9CFKEP5ao46VnVwNUKPw
9rVlpACZQdf/you1envOxgD2K70uvtollGwEkHgyC2xhR7sk6oQPFbLWChjXyI9t
lWYxiJv4BTF6+809TDLsRKIvidmmHIpBuPDngwXqZNxe95XvJ5klhG7vXrymXghd
0gMz+U4u65Ixzcl3+JFqdVoA+hgm/79K+DDCAnw3GGn1kcTHKd+YgXDTGI3xYGaH
wdesAlgSWANMXbwxG57ik2Dy0RyUthspmyAzVIwUAqWRijc4cRaGRiy4oO5Tee6F
FxNcv9iroX/aLCx71IUBMUTtuhQiYjOe9gtVf7IFs463Ls2eJ33d5OloccIKXqLb
aWPyf7PB8bMq2ePH6Y7vePydIi56O0elhJu9TnrvtyFt/0k6m3oaEgKjp8ZK+BBP
Omr5zmVhObPeTpDSTAv3DIb0sZN6gsG8kk3s1VgUzDOATLX2qVvhX75fByzXr/4M
UWib9nPdq+5naUtE1mMcQGepG5Y/uS5xCSFh2FYtHCqQ7vOScLAucLCdYeQOX1Ny
V9ItZgp94UhHjL+QcQ7w3KuEkYYvo2P9WUD84TMso6u7A0WgkhpN+ZS96bOLST4L
O3wwgRe02z9+pDgzpjjTDjbgfBpBk8DUT9AAqdweEaO+Dqwpac8Wwf1hM9V2lfjg
pzkZFzbPItDThS2KJ0PfsYJrakq42yOztyPOk+r/WoatXSuFObPUBpk9ZKUu0hjw
xnrB4KHYYxCfv5N0fcUm6jMvAsYdr+3seh1nYnKsrsIHUONh/CPJMW7Mj87jPmip
MUBLGW11WGKZ/NLCxKNUwTg+N7UowRZw+2/TZAkC5lE6taMKl+kMTOXhUOKKMtDy
fo6Vq36EL6hqAdt+jlf22iEM6J69V8RGs+EwfDI1GoPAnc1WPZ4fv85AWhqQxYdZ
5ZQ9uzYJtjx8smBRv9UFyEcfztI6LSHecEMXzTwi0xE771ziqZ1vxdkpCZ8kMVkP
lBIVCNhhsFY7EgNAMqS82mHDFDEank3SokTzut0RzrsOcnE9OkA6Zaqi4Kr+KyBc
0hvmBGV9z7AsUIr1YcPVrLHKLeAHueG/So+0gazt8LYAf1q4+fDYaawHsDO7w01q
+2nWYRETAAyqsXTqNyYO2is4+0MribBT1t2yWjNxvaTf18yalOyKHSIfBL+Hgvbb
Q3exk380CVgHpNkBRqTRQtyL/CqQY8S9RvH3MCSzFRVAnTg+nUp25rQbh8W5yMco
YQ08LAfllFWHfg7PAAJRAXdm6pwSFqPzpa/YVPU7da5M+rAnoLi21/O1Gr3u53C/
5btZMIiQyfkwTiyWWmM2zuXnDY9lds0tQ/rVzdmgFeyXgV7cFAQtdouDnnz0o/tq
iE79IofIgCH4yRi1LyO6uo8MeWI00xG9wqoH5XUS6t4Dzw0FdUkx3XArqNSym7MV
5MJjrzK5961UJk4Foi56t55jdi6ScsaPSRd7rTVn9T6vvDdEXK22rdQLMBr6M4jl
F4l+RnVHNCdYw9pvn0+bWzgRxmXcw4ozpNKxDDYOv+5pMVLkDw8yZ9k9VM2v3FV/
+L2jWFc+R+2k+FipdE0Yep1wkrWCGx3II2b70aiYcaQT5sc5IytffRYblZSU6sf1
EQj8RXn7r5V2KAc8jKwD7XylcXLbN5/MULGHCTKHrYyhE5VuoZPJj0w7qgNZ6vHb
2awVAEApK4vlc8GgnjCJgDpJtdbPiDUi/UGaaqyTgkO0gY2UZ6K92BSK40bNhplw
90JccvN9BhKqTCZ74+M2jEjxqmTrQzOs5yxFb672VzQUdMqEVV2znrvqW/J3ZUB2
Ye22s7g/nrqO6cWaARal6JdDP6L0GrPXMjyiCvKbiNoZWbelidvEeyha/Yo5Jniv
giTQ2e0LaK4Kni3pAgBtqiek9a0ZE+8B+mNikT6UbciE1BjD4ajqOew5vLN//IgD
Vvww5VT4NWIZY2nlJ+biNt6IvTOGzIcjkbYrZzE2ojolKWHuYCElWASZZpk2J5qe
1zYR1mtDTPoHU/lUJYpFOPL063iZYKMe99r77o28HHy1ddR1OOVDDT5WtnDBw0sr
TTd/qR4kOuQ5Ccr2LQ8l3+TsiB+tZeYp9psBSVVNPMMVnPpjFfCxxtwQ2JGOsysH
ma+cArpvVHuWps5BeVyTGZVETYjgmAp05RDZ92uaOppVtfOHF46GZ0wBQFahExw3
/M8Jp6oARfd3bYEiul8nC3T7pNn8ZFBN57uBXsxYdDNLBImJP7W9/JgMyE8HEUkJ
5Zr4H6v1ch+km0/5roiwxKfzaIlYI3/P7cHqYPu75pM6b0rUY70/Ss1BVaSqIqf9
Zu9bVorq/ySgZ5mtGN95d7EKlcfYi1ksW0ZD3o1Q9saMK6Gn7LMhYdZnr34yU5xc
U6nQ8Gw0eTXmknywXwmYWznlhes+Pl598TSZir8J5/+YdW+2/GzZJ8Kj7miRKkWE
W+C7pjcvaomgqv4VntIddcMqxSDIhKC8lUU4kSlhryYjgkpxpRZMOnXeUlP/X9FP
DDzlH+F5X2Y8KNLVuytrF6Ga36rH+P+NpNsT1PNPjglOUIveAtbyGmOEOYKuIKY7
zfmVGUPFukl6QNpnWlocHrWvcUsHjoXGR4wn6iB0M+F55DVCMKlvDxvd9WhtlP1Z
MFxMwcepu+bDo7a+0dF0YvqyRI4VzORQvnZGFkvwHfSog6cs5swhJiNT5SDgkbv5
Gywo7yZhx9ybsvluaCEUNql/hBKZg8IAretu0eQjzr62xK5J7FCRiHTk9rFki3fb
2Iwo2F2BJQeu+fVAtyBoETmdAm/vVFdC3LIeY7xeKIs7XUAtr9b4PlPc6L9Kc6mY
xMsU8dY0lU+sIG4LZc6t5sjslb72gWJPI/qlC4uFjBl+yVnmMIZQF6HDLxFYrhc7
7K7ZU8NsVAqFCmtxn7tA9v6+V8eK7m9S42Y0ILbUM7xGRkcFJ+Um7t5WPPSqaWQY
uM6WwVRwTZxr352OuEa3YWrb+6mM10U97GtOae9PXSMsaRJLQPXQ9my2OGuGURcC
N1DEGajks/5PiQ6FXrT6/6YZXw7lbnFUYeY43kRBMTn3nvTJ5+WbatI9obj67cUr
eAzXzTYsxzImdh+PcHTxyJQgQna6JFrtYq7U5/pul3zFIUYNA0Gm9foQKzpuoKNy
tbcViouS/Zj/rmRHprPaRs7Yc0h3vdJf8pNTTOYOKp0e6UkfXYPHKMgH36yoEAiJ
SF1mMwAn6VoXDMOTZaoLoX2uPb5KOO/IuDFeMKDoeR6eUL5YUCpXwUdLdsE8zt1r
R31QOFV+fEYCrA/PErf1sAr4VxproCG6wYBdtvgjAmObTdpr7CI7WrXbOt1pdDr5
rpSc3aqSeVWd3CFVhBKmhoSrGpJq2cyK9K/5j5/f5R+d/Nb0VopzmMLWroMag30W
rA3dEV9t7Pot5L7ju4uzlZvNvJ9kgUizeoFDlT0K8+Bioa1PjeE6+kXlNlH8YFNy
rYhGb49S50xmri+Wult1Z0N+ZpoA3hzjAlH/g1sBy/72jt+aatDBaDJKZGGDgZMT
xsjGZdCgQoHnWPBFKk1O8yauvWQXjGgERuMyOBstDRIb08RSpDSSs4KDogFcEFek
tQMvFW5uFJ5isEwqiZWF5oMXNDcp6lomzEpYDDIZowN2yVlFVsmd7w5vctmc6bf3
l1KvXkWPcn7xN+HLqx34byxc+wLTHQ4cjzA11PRQCSEKofrn+FdMNC1z+HAPgUl1
xJzW5WW5OQCa/r3i1/XqE5+1sZT6xBZZSyht0weh5zF2ovoPukjt9o8MWd0V4EdR
N3ARyXQh7W/+2JmbULU/SfKDzsrIQCA23Sz0PRvKTqa9k0tMneZ52DnTCqY3RAZd
vbDCQ7utkHFSmTJBDqwi/Dzuq1bRTQVe4PZDaSjEUlexDx7HosXTVIaH5QYAP7wk
RphScacLMv0y/6fvUHuRxVuNdkFSwmXqzvX063hpg42pNOT4MtdXCGjuTGksiR9d
zKCiClBZKUbNTigw25sq/n39Dm2O54PsjSoPW/mnkke3biinDG+og/wgDvWkO9de
DDEVaVGI43jiEB9iRDZI5mL2Eb82ik6jcsTMgVV8polNihMfqvpGdTH8u9XgsLQh
FM08AMncUxIGkDYpOPn1qQxj4h9NW0B+qqJ1SEJHKDEGk+LpBiIitfNpcrxz6uxJ
+K/WjWyxcUw0wN55Z6hCmYFI29VNSZw7coVEwEGREyKVPfYM66tI3C/r0s7J9Ax6
dlS7BgrAMF1uNqlExv5lU3FemndGlSErlEtghjtfkf3ZClpQMi/LEZ0R8D4RSD4b
Cs6LpLptJcEsmSOJs3vGoeRY1L4NsHilC4/7N8VHSf5jUqheWuzKRSqVjmfkbsWR
izv4y4Uv/e04OdQtf2s0b6bZYVo5Cz6gTMZOq5oQUEk3aQNUoEwQr4jQ/vwaZ/6p
HZRBOsIlTOMs5g/HiOOWWFxYlR68Brg8v0Zr4JQypXGSsG8/PDBWrlbE80DbmnQB
ClngwaumLddj6xxtoH1Wc/LyDSMDPJPdA85wuopm5GnJH7rLxuLF5wwWZfwu71T6
7AfO4DONBlEO1mmuYYbdGA4QUTh3bx7rn+aTKICWCkMHM6Rt4ECB+2AqB+LCBkOf
aib4AQYL3hKAvpArolNIK2ak+FJG9YnuQCrX1BcUJw4iSbpq4c+t7IhWxnBfqtnx
F5ym3x3Pf7qoFpS0VpRYui/0ZquozzKavDIYPiD6v8IvbT/oFNayvFQzxgFwWcj1
rQC9dKfjMeBtYia9DH/qTfyw9DAAVYchlLYQ9pank53SYLFoTRK+1KrCKa9gyATS
za0E5/rsfKB2BeH5Ryqxc4AdExP34sRTTXzUoGJIL5UxNPxt4Gr4solz4esCFm+/
nFbnpDoREQP8isiob69Fz8Rr+SGZuse4qh4Lp+sADxMpoxJnAk/O6ECD+xTlOx1W
FxbFwdcmt3OVZXYA49liefkhmUw3guAdK4+jQu60IRkhXex65yqUKUSUJdeNOrqh
yFrOKOCn7L0zgLk9WswvcU6lMTnnrHM93aaTpV2qhJpNyEK3KM7UQl7np4wYpgI7
3LpnsiJjua1o6TyupH31UuunZoU+NVEsoILa9M9oLOsKUiuiUlaK6HeLsmQlN27Z
SZCLY1qhntK+hD8MBsYUfMuuviZmMNba319pIFG5z+idTcwg5UdZvah4r1VpH3UR
5zNl2WRuppvRZA9tzMyfRj/QUa8QWQH+cFIARpf4AGhjh6iqR6aO0lXawmTRCP9d
/jiBZ5Roj8KK2lh/8ZausohfMOLUedvJL8Q65HtWQjOybZmTZan7N5bTNLP22xki
aA9vHFrtGvVJ6c6poMwPVsjZdOd+NoH9Ge/lAYaKpr9kqRrqFu7jhR+mSxQSEasl
ng+4acPa0VJWt0KqQjvrtqDFeFCNMe49mZNA9FMU9UBCCiQ76OcuF2fPKCRAcyFq
0Dz2cHUqShbYfTPejdaeOR0sDEmxvFLMXC+OM4I2VIDZDUYO4+rW94HiW+8guc3z
Fc8H2U3QDDY1PQBd0gwvoH2OJklAuSy6hl6K8kWy+j0uLIA5WrPJWoLCFO7af7ah
juvs01WeROzNEvH+V963c9g+gs4J7Ktq+/fXjmMiAfeo3le2iOhnfcHI3JkKEXsl
jTRpLKtsY6ySUerhv/T/H6q2t1BF63UsnmULALUQJXsMWv3qX0NsF1lF596pPFiQ
wlUnRe3HMcteWBnq02Qg1zO38YM/0gCQQu1O0ajt6naMfMNgP3GoiPOX6iihzIQn
fuiaR9TMqSfcebrOA01Xunb47owKaQOi1UuDTs7NPr77VyCWCPVQOt8FUCyDYYob
0Hf9ZzzbwstHz/eSYmqXrdIj1NFkUZUo/sg/UO1rnCAGZfD2CFJvbWPqUH91ZxGD
/dZ3zhn3ciGT3kJ1ExUJMnH7ClBXTxB+z1t46ZH2VaDYTDxrILjK5a0qvdOE5VAM
1KzM/HD/TQrQ6cPA3XS9qLXfwCqTcBsWBGUqEuv8K9dVaJMC8TSBa5QkRkZYoL4Z
lanYXQXpSdahw85OOgl+dJiWDVZRa4epI0IHqcSJFciwBGzq6zjp2tF68kYe60fT
4rh/tespjS9U+GQkWqALdWaI/9xRUqTmR3HeSoh4edBUWGRSZQ09+VBiXgnKjmBW
8RCQApsRB7Jvz2/wy9ZmIOGBzeg71sGQ9wz0e8Yxkjio8pS9uQdC/FtuVHFBOKCc
NSrYb032EmGaJ+2Bx8LVtO2xJ6ubE1IvuWD2X61eLyogP5Bh5+b2vULKyU3jQ95o
sUkFkvELcPkvv+tfuYrcPE3280y8djRMohsTEhUaP2XUJC5yU9Vd5ByLaMpSeJZ9
VTDF6y+M2LaDL4ov32tafF7gpgtajnj7IlCUnsjCLxu06/tXeGbx6KXbKKDju5Tf
SPwvE+m3uagyXOjWmKSayUBY0oExNQybecDFd6wovncSUMkZIEmgYwrdItmgqTLu
JjP3Ka/vpNiX1JJJv5EmqrNiH7UlfrgOsyOUcsjtA/DLpt3K1QaVC0ssB825n4fJ
2bYXOTJrX9o6nkulbOTMg6+eSHVSc1NCRLLa1RxYXihmQWaUOybJBhHQvnsdNfhz
V0ZTnSvvWOWKlu4G9zQFQUc5Yn9tjMlFmGw3DAZCXh/s2z+8aG5QDjs6RfJswTM+
mhmdWr9QizkUwiDgZfyUa4ZhnOPeilr8eaAry8fZCbTItgeiJnu6D3HL1N9kXpcd
vTVUcBVU9j7NkB4UbYyjPze3B/zzTv4R7XhR9bUMcH0g1CFrW6pEgE4+ybGLiy1e
beBSQuZXlVwCSW4+8qlKZuy/AEeJ7bVxbel0MVu8uNPeIWk3RgZJtmOx7KDMRrbu
QO5Zerc3XB+Moln1yuw6BRyUg2RbSK3dsgEHU+Hz/0V5V7MTIqTPp1xktngfaSfd
p4auxygp2vcn29PcPB4ioxoQY2c34KrCttkU7xBwzbTzai71bHKjvD1/tlR6koGg
cHyM63j48y5iBG3htbLMdQ06/0Ynv8SkVm4tq6bbc0qQmc7NTicFT41pwkQ6NdFu
pbmDK7lCgO5/NLJjrnHUaZeVJhMyWGjfVMkMM37qBeJZ9yk2y+AydZxTZOkvvPWf
fFpYQAcOpwIyNmZ7jZua6tekutS4Y9Pq1wN0AT+wHC1CzHqTC2hYln979wlt74Lr
4TZeNxdzTYuePpeJ6R5614Zfaj2sQw+28p4MHDzu5c/lU4WtgtGlejy0tn0frAw2
a5/25PUCJxfEVqt3eakXFeiLfGU5oJGwymu26iFXCcsl4RW3vbL3RjAujNojYOUQ
O77uNcf/f7upZFjiOQBg5ZAHCEGBpM2o1GVYj708PdsoA3TsWM9eIsJ+0T/JDSo0
A0ga5gXzPy9UvorJVe8JAoe1Mq8z9bvRqta2gja8RoKgRUYD9Mc8U6Lo9rYyvOr5
p+cVL2eztXJAnmnf+b2wsn95rJUlxULH2MBV3kBVfkMpKAl6HMR8YbKhXaoPOFPz
ebmu/PdENAdOUrx6KO/xK1mXF8ZH4AlzUksEFL56VdqiOR/yadaDMMz5YKFSnKr7
sOjYRt2Yjf4OJL3WRRaXuuvINgzg1mFGVdLfexniAfyDYrH1gRuOjcYlkLOAsQd6
prjcDA2NrS5eU2rbSrwILH0pNX5V4sEXSR5rWsP/HO2h01mr6WlkCsn7igz9Xvb+
ZKhdWEOgN5jYEh1JU14MYiRyYfzrYVn0QJhFFjfMbU/RL83TOWYylmc47zIs1Tk1
1ZxyE//mVoy5QyFJQBeC9Vx8/NHEHisEZzwEKgx6Aozm3Rat2EpOqvZGp7M8V5Nn
WdSnJ7n0bpxuSdt1W5qAcIP0sGrWbkqrbecAXKTIf1x8faa/3Ajt5bhlbe5P3gAp
s6UieuvZAJSdfjudpU516Kk6Eg1TOkLp9c7KFMr/lZ7ccL6mj+BJQPUutLy/iDta
xYYnLAXnqoWuloCdPq9XijsvJrCjy0jPOGu4/DGD6C+dkFO5Wsfhq4DxLwi/xyVy
LflEHJVKjJbC2y8joRYlzLaGAY0duLO5csBPlm/XzdTfwhztZpZxFpkFKU/yhI59
FDBqZHIN5DDUByVku7eBQN/XhYVyk0wVnaOZCjt9dcR65Ud8qxBLbTlWMtIzzy1m
UEp7LkNMGkTVjoQmhDFnGIRObgDK8tE1rEMbodhTBK9FQZC929WiuQZemCP6xEus
XBNxEFmhzJ8qYyxfUoOAofVTN/DckafVuUEiDe0R4hmUIfquaNSy99KdX2D0K4Vj
Mz+8YXT+ibb3Gf6evepqUDHRbnW5IwV6+xBwvYaf3XKEJKuJplvOtNVPHNBAAy2C
Av8VmxsaVfzqvrNChRBllxIshQbjTxoGbjCJ32/EkjQYetE0zW7eiR6GAY9p+29n
epKS4Yo7sHd3sT9Zj5ZHx9Uzuu65oDevpcQHhiHloXsVlCOR2pFH3M4UaO39D6zr
wkBaj+BZdpIrFoY9DuzPLGb/WsVouXcw7w+4XMdvIMOAoe6cdVEtY89GkzOYeKiI
21MxMFxFUcJhJrx371leiR4PY2pN0DrupCYJ5aN0PZvNENj7OPpbDTcIBl4eNLAE
RBqwkNcSymBSxjNzg8aooPU5be9MvCZlVQXmuJzFDn4IhlIjgNHLXk+SAA6M5DLa
bofcFExmqES59i4N1tqtGDFGtqJAo09xilHhXkGJ3+0K6Cgb9+nql33+Bnb4ptAo
7sEcXXSpd9Cw19ccLcecPpO1ErpktuHXihTGuNhomHfi/LM9KCcPVuZlx+obZIwx
HUzFzYDG89B86seZ1oRI0Xi1Y48snyAQKr/JYjg+oVN0KQBAYgzPKPDrEikRz72N
ubeRlRryuZ8Hm3k2KQokz1hqjmNUbR2HZagcZfXM+xCAvzCDQ8xYGHTDZiGuesK5
W5HbhpdUTUjRVddpK1QU6CMZEi6VXbelPUCbug+qMKIfeRDvCQIYA7vtoLNaRERx
hdHZc75kwuIfKp5NqBwRFM0UcwgqsX6fGSmIPvHMcN2kIv5J0DymeAE6FbmPS5Rt
/DPCpVl7Y8mIJZ5K58UZwHno1CiBV4JWg2cRkOopVJPBLbFemsu1WVAoyiQhQiHH
Lo4eQxrFWYRX7Dmf7uTOScKsNJZoIkCD8nTjjRyjy0PVBcCPCIPopeTRemdiU5PB
8pV9mVMUGPgvOVOQn/BTn4/GSY8wtPCTlxtqnAFzfjvljm3elqqbUcHvuUPQMFvr
JSbPC5jaNyCOFmHWcEHfYrVojnKbTvqI1H1gvAR5y8WcigE65KZWyJHvdXv2+CFg
3G25J/K5hY2d1GxFKDG2lBA7uejzxqlOYhEvzhZlqQ/PvbEBsSbV4pmDnt9Va2b3
sNukT1+R6YHXvGMh9hyGCQ/7HmnFyJM7dSfLy3ijlmOgF/Mm87YKH6Xk6XfH+2wd
faXzzCaiF7wtHjxu02KAW22SuhqKApm7C3xS3MCNLCTZbJZt7S5/dS59oZuBZ0k/
BH8zSOZhmUVijCjO16r8L4xxnJpixaApdTMfEH+M0LmRDzHm7MeaGJhwGmuTrZjQ
soa40XFlkizRv06fN8DRa6e+z6Sgky3rSOVeSjvQZ/t+fUciglcvxqvGlrqKgnze
kuuWVQ0eTGkH5/ECFgMxAEVCYF+7UOuNrFF9B/2UkTRwXUH16Zn/nyf0+Ocqd/Mw
WbpQsXe7KVBIL8bvpXcpN4m3SiQ519HmYvaYIbyxhm2i01Z/hImWIdI8PfCPYMX4
rxivKl/avOYDn3AjS/ZhVYQZIid4xoCDziVM1fBWj2FMF6oH9mH7Mt/jn3GB/EHS
bhH6DiB5L++4gdtdypkPmTx1LGhu9kg8XV/21944PqrysBlMFipjlTNNBbKCHYMm
dTbYTZnBFAv5mGkwYdYk5LG+DhaSHT+g0+aRcDH4FxNHCptOFfIgFHZz7F0+BYMH
N5PDuO4/2r6o3tYhF6FXfyo3RRnibkiXQInwHSTO7Bh59BOssXDQZvsMybHcJPmw
3NqnXwNGivtyM7+HEbtUEsk9fBa18zWjpEwerQXQQebFVd0ydgDJYL6Ckp+7ztDy
zJZWFje8CKi4qCwVgiO3IwosafYpwyEy/7zbzBkpse6wSd7BSZocoITHft/MeSIu
geoCeHoZ5A+AH3Ve4vD0cBJU2B2yMw/1S7xzD8zFiZ2p6M+Kb1p0SJoT8G/8phRY
9wWDL7HSNWDbv1/MS8yvlCTvyX5t6alNDiigpvlc/vYoKtwATQis/Si5Wh+lM537
nM2ZoldVeWtDEtpzTAH7A4GdrUdZcjd8keZOTn0xFrPi5UpFa4unQmG+B7ppGR/H
YP4ex7OZxeLaOgfwQqNj9z/k+q+HmZITXeiPmkqObjCSp8JTOHvz7ehpyZrzSb3Y
DWhHiktb/ZtBj3/on/EdnpHbgYgIkrQKMn7tp84Z0YVWvPksv/Y8icSFVpMDrTKa
JZageHQ4xLjcZEILnaI3ZpdFPoGpzJ50g/NVm+dw1Gm0llBLP0PHR/mueE4t9rR3
l3fIgn6FIPuB7dCZH7DVHD3PKbjephdFjTEgcDWzsJSHyuRoC+qv/cTMNLc+iAuM
194rT0jU0A2Ro2pPX2f3M8MExKWmIT7olx7ckWa24tE9FguqXVmTgekC3hIk+FBU
ibforNqxHXMs4KqkwJ0lTFwG8xAcnW8wX7c7zxtWn/TVigaPsbNi801Is4VkAQsH
zc23gsQxC9U7I/+0yodH7mz7X/6toHMGQvlYlSCwBO2NoSLZPqimgWK3pfB22daZ
tWMuSJY9hfOCiDhOCT1AWxq95hwaOY0RRilk1wmBNJR4a1o+ovNXUXHeucHgEB4B
u9K6cPA9PyUR30mZObnrWjI3t1N0YglJPVYLqGevy4M2t22g4VrW45K0Y7/7VjIu
dQ9XTy/iHby7hnor9Iaw8GZbcU+9cIWPeMylfEeZlNyHpAZH7lcbWooC7Glh9UJi
EO5aHvnxJ4U7lYlsuplPx0erEUMft3iiFiIKA9nHQviKNqLbDGipSdb7tTxtW1mY
ZcEz5NcaIrPaUi6XGLhL8/X/421FwenTZBM56Zx4G1NP84uskmo9ez617Ba2b61C
heTRnIgMNjCU/0kqyUlS3mdm+CWTxL/PS3Dpp9G9QO8UdxeHwt7owc/0LDn53QRu
VwaWkD5GMgHnLy+jqbtL7AdRXHNxUpjlcQvj0K8EcyqxjHQ9LMsmy/jVDnVn/CRM
pUbE+r2ggiMIZipFAWVzVJSTGt0VUlyJ22gqABHn9Ymn722Gq5XHyFJPUAmAVcDX
9pY3ml/dzG+4PAjz2ErdPv3t8aNYuWIp9aVFbUZtvrt/+lL71fqhdweOGls2pfAq
H09ojVExU9geYl3kgzuFI15j+b3E1aILrDqqD72dyqxB/jp/AXp3vrGEE/fl1Q/y
8bybbaJbhmm8077xrIgz+F3unD1f+pG74UjDARGhiyk9+t3qRQ3lb1ZcR4l17BxS
rgpkpwC/px9jVU7midTTDQiR2GVBRMqluEl+dYbcGBifT9Zyp6IJa236zGz0wzv5
N+53btjVW4vyb6oTWLVGL/nYxwpaxN//0W/R2F/IniLntw1N4wbHagi5uzmDegwI
xMjm1dgBXLpdy9pOmgCbkAtpD5ycv5S3WartD/HIcHDcmynMrYq8u3mMa7va+blK
seHJ5dV3wKHr0g3zWLa3dE+g16Iu3OxP39DQ+rippTBxqNyjh/1K7nAsOaYJUaHl
aExPieyV7Qmpi6gXzsanG/lTlw3aeUdPb2bCQxgEmzOMcTIaRldiyaDKm/XlkIEU
/A47ziMU3BQgGntpwcaaR9E4ud9kZwLTb1T8E5MBcoeavhpYZEqsQAwRFLgBj1gs
IXI4paNprzUNLFdQWUi03AU/D/e46kR/iPpCZ5ebVK9KbI6GdrQ9YfUEeHF1YUCM
c+/m7oZgPEbS4t+cbVU80xwI3/Sc+gr9k7patRBw5KQHmtnm8Rr7v6VzqEk0AjnO
efWF35VR2q4d0eDh7IlMwmrAzp2Ni024Sur7H4O0vEhJGU+BH8xTs5Nkm1cFP3bI
23YvQfhccV8JQwFOsk3iYR7mVD1diZdpicKa5WwKX9ForyO1fQGNxoJSxUf/ocMj
u3oMhjb7lpJ+mIdmY4tvFxgIoDqQlLrxYPiFYNEPJNXqEqkq10MZ9OGgqPssoY+U
0cXnoFPaVCtyhKeMIFZbOzSUsDXYYZSCJc+tT51BEmbGd56BUlBj1dPoQrdV7o7n
eaOT0521OrJneRl8eJTGQVM1kOsJI16SgJBlMO4GL1h3MWGjnYhw4zd/jPYpk+dk
/2kmRNTmhukTy9+A+1L5Vqn5I5ZCARRniTC6rm/Sof4Bgg5i2/zDVdfCc5prbAXD
BpUDkJ8vaIAO9BFxegUcxzjIylksVA+JGJcutGuH1H0vuPmMmHBy+S0+V6VC4wka
MBRBEGAspqQmah3C1MAQxEnTNra+LX0dSNFOQLbmF6KIzQdukUq2AhX7MS+x3efU
77+XbhTboLhFLA5ChlcFNVUt33zACe6PkSbIybi7He42KVcWpiv40P6qqNndpCKW
VGNB5FRFvWvmF6yGy6zVGf0kD6D2SKS35jiGGI8wtnT7qfnE+gyoJQhsjgOmCCwl
OVxDRBIE3cddQM3GQbrYxQLO2NrHyXjHDoZTaXWftAiS22N8UqYKR8NAuVmmn7bU
/rrDGg8dv9OWfiEQh44B5vWdF91lAcon9vV0AQa+MStJdxHQFTEH75r6sxXPnWge
hozu2g5JEyyFQkZcgoIC6T+ZFaSRfz7GTE8B0dE0Pv3WgdgCWpJHMvTQSf5/DIa5
BEM9aFgARZnrw3VXYYGUbEvKupcQ/5SnkIqz0fbv+TWJrbzKumkcotDtJhKWxhMg
s7Of/NWlcfHxKjr3HiG+V+UCuO1VUtJV0nPFIMdEfm1Ns3isuKtFh4XjBDhCfy3N
W0iqr37mAK8t3c1dNfoB/4/qh6g75Ld0fqD9QN/bS+E/wr6XFHjaFjIdmH+vPDFw
qctaLdrkxfZJI9DE9U7hdX4TiaNM3pwN8UO3dW3WyDXqbgNwBJU0i590u3AGGmgE
mm+DExUvnHFsUrvftuQ6tCqF1y2Kcwl/CQO4J43if99S0QAQOgKTDWkWjNST8Hwn
kWf/SzYAP7kbu4i/cgAmnuhYiX0TFeedcESMs+LUPuvGApvqZK8n3vDSwfmZQ5sc
RqHl4nanHsvqoM4fMJcnP0YoLgM8F4PhlOwHG3CRTwob5Y77r2rEPjQzD+p1Oom1
9RSS+FNHwM1XkFZtjKbwqN/10Rw818OoEPBn8FCITp/cxefgMfjR9hVPEGNmU2Wo
J1BKODckSXfCy53nkhVaz9ugxcYErF5UCM1jwUgo7x4bE0rnOuKym35P1MY1qtgo
LHpRtagyvxiaabeeILJFtyGxj6OaRt24lWBUtv1n9dqV4Y99kVX2YAAlHWaYzdPW
DXNi3svJjlUHhqwk8h8HtNqF1CbxHuGDTBfXTU+KIIzC2P/Z4MuMo7pYbGwNm8vp
KCrUttC+Bby7oySt/EEQdYFKGYH+sGRqkOpCZev5Tn6UgAtJ6B7EyCraTbz0xv6H
3E17NsizUHvtMNWFmPCqD4lgRiAk7FMe7tOaiFpem8YeMfHOuHXQkW4Tr/PFQPJK
I6sLLN2Kx87MaOpWZDhzg+KL8iy+6g36el3HoopjTXxTywhKKtVnkEiqwMISKvaT
pg3lpDM+lrIjPTuWiOh1UuEq2Zj3MqmFkUnY9S2jauauXx7YLn7c9rRiVqmAA+HI
gnxv7UQ5cKPOOcUYubkECfxhtWJyPKolMav7CzSWM7SIKLyJdU1qUtMfmyb1Nj2C
n/wgQspVDEfJCX3R+06aLr0GMUEgOb/ybD3Ihz6bXtBqO61OYiuc6VoqiOZVpmRQ
4girZqLXJav8md+XTrI2ye9pozVa509ILGKzdZiguM0ITQmk7sZtVrXYRsn804WD
H7wPJtEvk/vtXfvsYTrjX+jxfu/to4sV+5HeU9gOZR6s9lHNzg+8oeIAf/rvpghx
OK2ekFtr9Ey5zS4fORs1jC0+xn48OQe2mErPlvIazkPhO4En9pYfFYFLPSGLzCLy
AvNIedLZyKNmaKx81ws6RSZ1sGm6vGeilxkuVkwVcNo8zfu/tIYKGAnyk2jaSCAQ
PxivPff8QiXWzS0GzZUITUMtVlx+23/+bvBV42rcz6hh+N9OTjSgqk9X2s/ysEAt
G1c5HRXDKsgYELI3g9N1veyPVDfoz7nQuOvkuDDurz/l+1EmRtikJtvxbW1YYYdc
Ux/y3dI9PhPoXzlfhTojKdoO8Kr6V9MCrf7ZSxw05yQFAaZFl7CnfKfPYtzL6Duy
rafL4ZlSopuGRolSWvH49FPqKxZe5rDTYykqZ9suaaWxV+GEFZksv3QJHzRD2pU6
ktKgevEmSaXbj4njvVEaiir+gQnYdFT1GU7Pzx9kwdo8O2vbW2j90QWLqqhIarwP
+Kg0Ofa0i1zyZwKQ5iDKXMzv2qu7y0W6vNv3Ad1zuuTwKsL0M806A49RQNQdiSBH
sqJdJT5qGstS7tN5UjGPgPcnBPk8aAFb97qmbX6lvQgZ4e2xBA+604UckbnU7JRh
5n2p4m7HvNB0riWFbxxtrddWHDXt29UCReR1jQ6UJ1Q/AQjddRvBfKBdz36JsrnL
fwuFXXXE9KSAR96UFbotn3CWlvqz/5ZZ9KkLElQcmYCrHlpme+nFX/5iKgD1jtbX
kMKKkqw8jin2uqaAWu34LnS69UpG3JIe1KPzJgF1Nr+5NjyvFZ2q8AdjG7SvwhPr
XLWhoB84F2sxKflIgaiiI4/o0oZIExB1ahqUML4LddLA/7ghedNrwdFxtr21T+cM
/B+35Ah0dorypvakiEQKuvw+ZJwxN2Eo2ZOHePqrP/8K+wyp/aUIp71a3Bfu3om3
nb0TGeXHERhpQmqqL5LwE65MRwhsAHxK/nL3g4aLozusRCQoYWhXmzowugbhevZc
BYD7mEblSAdHCRsSr+abCRkTtsusPAm/OSJ7LESTtEycwpcgJN5qrMPi9i27kSqv
yQ7Njqe23oO/9KsPee1Gcx+xdEPLsSobw/Ct7GJkvGNJX2HFG+9aPUxjF6V7galc
7JCd0u+QpBeJJRW1fX0IJwNNaRjkr8P0FtmReVM38YzIn8nH0LwhwqcHFnBwd3WN
ZIVfwrU9F77XUW6OvbSgSA6cgz/z8fOuD+CMVhbhwn8kCg1+T9sTdbic6J83/F9F
+ZNjtIVQxG5tsnay1XmMAi1dKjmDdd3J6Mw8mfKIgdhs8Q30k65avWzLT0w5ZG/s
kr9WRCTKUpYgAmAG4vHLkPWt9/jiOU5C4JmTlKWSvrRLpjK+hqLFvIPpLX8GYqqb
bo5gvL0bCa0aBq86sKWFL2PhDsfpdykG94MbleVCOgpUUApeZPTgRlw8bmKJIyH5
slD0oy032mkH0+dcQgkG9TytKPkHnz/LoCU/6kFi9kGOkJbzZDaaayQNbgi9bfoD
SI2S5dDFZvvKJYG3npflo3F/tFuZZ1CBB/g0DZUVxhZ6pKeNZUagu0PrBcCZHCJ/
HMQwUp1gfP+SnPR8FcjGYqdJjF7Jy6aOYQM6sH5EdAVGUnteiOk5u6/QpKPpcJRY
jHxio9SNy5YcQgVCVoDASpFdZpwyF/XB9E+7TRZDVACMtDyZe15rxTufPuw5sAbC
FPiEtydUU2/mD8wJ7o8ddrFz0kEYmj6bwKPJleeXpntuhMduQxeEhX9Jpin1FuzG
qLrzdpHKhgPKsJuHeDtA7MPWMYulCypXo46lN4IPcClQgCOoUQWkZwvM7hFepIma
HagJ7U8Fxk7AAKL/h0e6tY6HPRJD7vHXY3z7eFL3DLnpV9Xx8sP4QHjAozioNH0B
aozwJLN4mncnPKwJlcPTjODqkNpLlXwIHl4I0VIs4qMNgHqeAZJdIkHn7JtqAxSg
WQueRwuSXiXFej+Y2Ss88V479EI/PPG0QZnoMxvvkVgbUxY4nGZwRrG+LmGM7Nf+
GfVFw4mJTW5bfUO8XKjVGqx6CO1qFAy15qdDbTy6rs6kIKTRLZajXQ7xqIm3Pd4H
grIKuf4oxfbSBl3oixY6LV3WiL+d1gMiAv+Xh0YRpuSHe/K7+Q3Xk2pQyFGXYRTV
3kefGC3DiRPqcyesS5tOEeC1+ReQK3F0G9+kgkLd41WVmbfWM60tJegC7yBsDK74
tkwhGM+6LElxr+87XLOn3uB3eSXJOv5CDSLaGDdeKIClWuK47OJc6cQioEYOhtWk
nh7LQOgjVfS43q68bUKuuFah/1JQ6Hpk3SA12l3KfKKGjHfTIFd83g0Th326C06l
Ntma7uYMXZLLgFA9r9BRR6vZv0Ne/Amccsh6u43k9p3XAzZaiik9A3UP1J2zkN3u
adu0sCFLciuObStUpMPxvg/67oTcQPKAru65UTxdIQ3qaYw1yzJL4NeFHJOKi6vq
KBZ3LV61UHtE+zR+GI1T3FeR757NbUfUcky7x0i+mDcc/9XnOkFQfm95mwr6x/L/
Lcy/yApRA6vefFhRR5e8TSJqXi00OP5hkgAF1FbKASPeidxqPACZFcUZ69VD/XOP
NaQr/7yFCjGQvJCicu/jLrxOn0rOTAwJX3r2Nl5eF97pdNH8Bc+RieMV4SCLfwns
mZMYAKOQr+F5Th7+qZM+yBIoM9BxG+QUf3ZTHUeabMsknh9hOIGQviefwSGrQfrm
KefukEM4U47JQPYjd2gGcyXkzYKrOyU2TaZjLAW1nIPJYKTgqFiXSzdtGEmXpTsX
Uc8oRE1WMEMyGseV46Fxy9D5Nh8n8cYwyEl3miBucgrkmr5Tw3wO+hJ3r6+m7KJq
rhE40oTNCaf38jQUuxH4mMdXxjOLxuqg5sfUgokgWI/K9POfaZy6EabqAvXfNc0a
QPw6e2W0X4QYqh1E2ZSKTBjdYv8YJ2BWOXOjmS0cd1A/onCzPvwWZ1LGqxWFlVLl
dvsx4+pzgjS1XXAZ78xGF9TV6tj0iXIx6Q6eJxXWr++zriGCsqRxE0tfWLYButl9
A5DPQNj5vBw1ESAfdQxctn7q6jv2Ez0PgUeA9PrS/x0lbzDDErZ07zBkdI0sSQKq
5lh7pHgoIXY7Ucnf6zEJMHzbRk8OGd3nW9tkZaUchyOvrE5WEJsbGZeFhDHz/g/z
rvkE6YtL1ORt7//469fxAfzxpOtJ5u8XBvCPff9dvcBcXsWkdedvky9vw1yAYpKd
gYE6oE+NFr+kHu804+qo2IzcP7aOB+WlOgMAznItEAaRgJlpxoBW/thUV+IpDTz4
A6189dJk1ATgSUwFCOHYt+QJdkxJ/hXM16uU9fQ1Nsl/rlA8Vq+my/6XSHNXFUFW
dT3Heys/vFN15CXb9zGSrV41BX4eZcUa6tJFDMFbkK31p6smRtkRHQscb8aQRUo5
QexDicaFQ/On4t+195ivQ+QtLZZPg4TLNnoe4HPqYVE3b1D4eOkcoKXtrqk4Szp8
c2m932dfeTXIUjW/5xJjhBo3clW5vQEHUlwAxaUYUXXlB5+7TL0wqjxHMEltoBzk
bwxSeMrw04BVjkYLMV1moUOQBN93POnnVtCymOyeLct8jFOa+IdLKX7SnihPgB/7
QNid8YGicJc1Zp3EtWjxtApKGvlLELT38OBUg7FvcaBrQo3v1nkuPXkTeNvk3ojO
7zTwI4HLFY312pwHAVjIOB2FzglWEW2uKaHqsI8dE+4JjRncPdorTa3kRN7fyfRC
jh/Zer3CR/0Zl++/wW39QmNGIo46uxy5xyDMosxLTOThYfoiH+6xVa/y6Dlv+Q7M
bmQoQfw3Kfh/7QxlRZufoEb3D47jbXeftYws24HRyW6oIlFTgGMUA+aU5L/OKwKM
CGHUFT8sCSxTN+571KJ55Ug0aBHKvA7jUAbhu2pROiz5tdUFvw5w9GQrfWws1fja
aHAPExbxQJR0MN2nDgYr27wwzVqiiVa9srBgqWkiqyBTL/CyCsEBIorCd+MmmLIa
OEBQPsRpsvWfdoo5JsKLluxEkN+EGf2McqPpA3cDv6Uzfh57oQqzW0dO0c/L53r8
Y+dTjUcCwFvO+33qqBYz8cGXOq9M+5ZT54i8bFKt2PdNUW1txKG47yLgr3hpTTw1
b4amVqgbUqus6BDTLJYCjxiTDU7TMbj5b2sKvmEgDtOz7dvMQD0Lzp5w7Q2Z6KiV
YOTXvkpwH+Gy4n/50ijMKaMXn+CBcCz8IvDLAwIUJHUqB+QGCQR9fgEKY9JlkMRo
bJqEYOVyGCCUgyDP0NlGPf1A9RniXTIcnCrk9vxGPuZUtN315EdX9dPsafy5QVEz
EDeRLG6HimgfgvdVVxmlSRaJxc9qtqvNI93E/SVEGQJeJmQT0Hb030Lmq0z35fkz
wnLUOr/2eGiPvhHIPC2OrYol1R40zO6rF0XWg0+fyZCGsctPj3K+59nZdeRDG52n
RlvEEMKr8mQDOwQsvAaxy5I7jSJpuF+TLEccVs67JL3MwXkUCcYChuZ8tYs0xmjL
llHa3nLJ4LxoOxl3nX7RL3cZLGBWaBESm6AeQytYHGz2f7ebx93KWPt3mG5Sx6mX
PNJ52UlpdwxU5WLmmGTm7uN/GMMuG+/upgl4hCXwsufCLpjLrUMaejfM0Zdreh6D
zsk9MdxW2J7Nj0ur6JBugRId64LsXVvaDR+E4EQIUHWbfDue+J0CtWxNIPATcAwe
ssj5JwjFw15nr9hSvGcAl4INni85byJT/h7vcVWwcF8j45EU4jxGEkpnmd1ICHat
rQs0c47HrdDCRUSRvVFgXZ3OZC6FCEvf3f+uxbtKhiJ+VUwU3yZJ744sa6+2PAMZ
1bWvPlihCS52pYqxdZWZG+ms0pMyOW2Mir6x5V7fPZxrE/fUbpQwOLR0bH8Pht/E
5R4QdsydTPxJhkBWpTONd+6+DqwO3Vm66dJCaoj+c6hoe6AZ+ZR469UwLLcIpKZM
gJnH+axvCFu+RKJ7sBlqHBO7EHtEGu9kw8LM3zKRFWIrUKt6tRq+J+qxc4CU1czs
LSn5yjx5SqDT9tx1D4E4waSQnSI6pyPH2BjAta6NgW6FGplhL6Pw/sB7DwHKYlYQ
rZS4JCu1EnvgdiByKnIK+hnzEhxHzwISnEusPA1pjXBn6D9PR3L3t9IgXtD0RwsH
eUlICJ0anzPp1AOjBzzf/wSf0Op7JBjhZc83uRR0KWmN7rh1DIAOWxjyD1XNkHxP
r6RIeoxeJV9+1n+DBNtrLpqC9MJ8foc1HNTH2xQ5z/C/HqOUvaBxsEDf7TwHIuqi
gPGl4m/9xPsakYA7BDukjbuf6cZiL+/ylMfcWPo4qrevFoeE2jV4enPPpPcGrB9K
yiygegITqD6K1aLYy6Imjj3u4A2EZDya59xKto5a5Xexbm8+27154FDpiW8QvFRP
wd2fl/8gqMUSlNsR0I3x5SC8AJjWIP9vQnRktPXTnIlj3UhR0CqYXDOI7OKjmQDq
VB5Ha4ItC1N/glfrfx+8vxsC3SynnctlWwsYsbFYDz4kLOzBzjN7z6HGb3ic0v9u
NOxFNwfFkrqXsRASmy9t8bJgtlgbOF9BQnKaWwJ1TdBF/o8kIFHIclUwzPU9IVcw
YYxiwKeGipgiVGAsXEZ4mX9kt3p+Ax+Jd2dOp0Xayk7E6b95nEJwabq3C9AAFzLw
ycsJdCmK2z/Jhn45MaR2VP+l9a6W+4Z+pisVuDToCiBAgFK0cAEeEaOLHZVwdAKV
GSXBPf039PxQHOOsqoX8SPQwzmhgepwQKMlXY1DiivmfTXz1T7QAIk3ClSmO0VU4
xMaLALbdEpl16GFK0DGt1U8Nrg3ZOOtrtKWJ0inKuwb5q+cPaJ0JCfOSEqiWhoFz
j42YL1ZgpzMF6OJPH/VQF5dZexc0yImOnfazFVXsZ8pJVSR/UhcoRQ7/lCTvA1cP
ZMT7RPnJvXjQLqgsRQuH4gyLXVHDl766Dui13PkdlwAyfQQjX+B3xUAqCxm5O5TB
zRod/4pURFV185Ta8Cp8dP1uUp55IRmALrbPd9lCtRDAAtcA2F0iwZk1KhVA6zq1
7z7P3hn1C8riJA9/PpXpO/9mbVzC7hmkuurWg1GJ0vvs38y1RXTcWvOBe6RRTlK/
I//fqMK0fxKu1+o7IkuzWbxH5DmCHbRwBZHXGePJsk2Pya1KEqQa5xSeKoRNBCGb
BZ6hJpmSHwKyTqrdmx6rP49TuyZ0RDx5VWlFG//jWahX0qUUeonuvTBRMxHfUsNQ
9rqZ8V+0KRkcdwCU1xKO74JJdabX+tGM2A3PzLI8iXoXNYK2wWMKZ5M/66Lyh4bj
JCy1LBLV+kNdsH+iMKNT8Nd18clLZ12lVttm0C4GuA/X4nzDbmDnzQXo6tu81OaP
qvT9a29fOXkvYzscSx4PHLvR+7sxs4tpSR6tyW0hRhubsfStYOplu6XGYPtApkVQ
8/IHLzc7ZsGkKY7eWRq/VZMu4h+DNc6aihtpYGQJ1nl/DFa1gd+jNpE6G/DWz+qf
pcp0ryUmGO5MgfeDZGEnWu5ba5dnU/HmALbgEI6T5SvfouBeaQtPOF5nofwuCgZA
V/i4odtirqQKJbHcqaCvuTd5ySV3JjmMpjCjCHVIGxOenChDc6ebaAUmpwI4elgW
MGwRct9ufmtOz29OzFJcfyjeNomEnZJOEJc92ZXf0vBp0m5XeL9vE2xoqfrD7RTq
5aMSc4PZyfnHJhJUq4d9sWXWi8llQL4jUbS9q+w2Tp2P+WtGHZwEkfMxBwvlO5bx
S7RzQ0ZcIcA4ACF3u52ftLZrfw9RJ/oUzkucSwNXJ2Cl9zSKUp9Ejg/J2tMxJq4P
jINNpo4I1/CoSaXCOrgASsAgAK2GZilnCsmjm2M885ePWBY6sc++UHnC8IMQurJx
wLo3ccDZsyICIUOIql+0KeN4rdtvxcwatDRPhCV4BUJX9YY3NjllgQxm7WA5KEet
J36vFLgL1ySvlBSuPqgnjVLwWssnjZxcaEGlelNr8y12p/U8JSch4iB9h8ty7G3Y
SsQ0/VZiumWYtdQ23MfrW1RFl9MkhaJ0viiV1VSLahzmV18Yg6PeICKzncS03jmy
xVJQ/Gm8pWAK8Bo7mD2onYpDu+8+Eel3bKJY1QgeqOEjxVy10GdOnl7qcvEOV4eg
5QntGD4J4QCF+y6WtGdwnNEVRd8yVOYWl9EX6uG4IfHsFpmPTChK1rxbnRJ1YCTb
gcCwvAVV/p+NUIlYUOIvOPp1SxashNEz3AYu+3VjXcUIULv9ujkhZkvqw3yTOuoT
E2hg+Efu6i2szS2XnUmtrrUZJJoaPpqVFdmjrpylKpTdFm+M5P8oqNMDuwM21zso
Zouy4Fw65Cc0SzFdh0+gBMyeE8jQbj/TkxUp5a2HEBfHbCH8CR8MUD+ZcusMERTU
aV4c1IE3H6nixqK8gvSCrauNOS+SJJeBwDmcvv7B/q5+LFZ58NyRtwIXjxSdOmRF
nc+WIRDUGkPD2kJeThDqX+mu0GWbTzaYmK63lSDxTCcxK1cJ333r8rnhUZ/Ur4NW
tceHdHd/440K900+wg5EHuRbwtNfPGPSs+HhSDssK2KEirqAkzTw21SLKLlqNCnU
rU9T9YylNr+YAI3X/+2DOQQoxNgoUPZ1E88UFDv41SrjDLm3aI9TQhYtA4u/7Qd4
+fpfOXWXDGg7l0n1cXUQKs6AaYAwj0mdw2IIZHSb5uxUe8KhVF2XoN8jtuC9A4fS
UCB5bhTBpGOql8uwPxIqqXQMyBi4Ho84NNL6gqG8aySqEDmcn1+mWona6X/KiL64
7vNsYkuVOstWeFemX/CqLkJoufr5A/Rg69kXSNL0flVAlClAX7IPZUOsGXHPTM4r
p4kP7p1C9urE+3J8EMg3UmOjP3fv6b0q7Z6owajUI1OKNKprR6PT/5D++FWsRlTM
inUcWQThluEA2gGOeJnEojSsvqZZpmq2vBWIl/qn+iF4bC7xF75GmonYvYUIyD8n
z8zigT50mFx/a5O6ZcHl/5T1cQe9AZRz3w3Q8cQpGSQ6caVIgRY4X5jQlK6OT7Sz
Pm36XCaPHaeSxPvsO3fFwk7X6Gwb3rqIIYqBKM8+61pxFdN2wPgVBLB+UUDhQ5q5
U6t4KfjaOKMSZIsufVFHOp2FVtMZiFCgZPvvQu+c01aXL4O2N4cA8ZEz62GIaZEW
9YJBrI25xCegkTf1gMVQkocduvvEdjOudam3GMjoTNM+2m8mDdgQnMCh3lEOZeYv
nRJyQndKYs8vG1zfHE+iNf04N1ivVkyHfYLMr5iY6So5RjJvy0skk+izWmxOXTVc
6AHiU2WfRnPz0a2f82OkNpGFXfQw4knUA6wvsC1vu2L28vRloms7IwvwScXLPWOW
XLbuWzx69pD2m5Lg/rLYDigHzEDcuX9f5VCqwEReAf3niYJHCuj5NjpREDvuE5p9
/2Lvw0ov1d0I5p+biCEApcW4Mm8gP+6CedidUFzJK7DjWiiG1ULJFq1otIzJuot9
b7SyuXKNuD5HwqFPdGS9rSIGnZUKBXy6RnkJT4OBvxLDjgufXvQCZzLiEBNWE7/T
3/QL3Rd/iBxODHySR4ntWzYwfp6tXJcDImhYES9rEzfD//zBbdMO97mo95j3gQKW
e0MfBztr1XkNpz6lrQ/zo/LhNOXMpTUyFuDRDCDXPrfvupWzNCY/DvAJka13A6sM
AXmIu5yPWP2ENLWXmFQWU9Q0Q91LS8kkZlkZKxtEms/BguPvShTjlbNshO9bcH62
c3J6t2MHJ0rUDhLdUFZL45gYRvrFlBGDcj0yiX3aXbrFnYfXP+IO+q0jD/iIynZ3
32nH9cc1cpeBRjeKnGdRUdWgdaaN8tBQuZ5CcaUqeSdOE2pg+y36RVUUYeItToJo
YMJXObjV0jGcr6ZzsvLOVXFELv/myiR2mNbQ3H6mdl0JfgcW8jCxCyztLtlBGo3u
sQABcDEBc/kk8dVaVga99vJJDdwcPI/jaSv8sv0JavuGEbKFTEPRDxO+FZ4zXmud
Lk50/dyKF+uNMJ9XqsTP6EkyWPZVA2nFjT/gdH5dTVadmMoyLCGmF/dS6C+K+hsj
lHx9FZLLUY7p0tp2DCChOG1oZHMirv9GUQo0VVDfHH+nbk0NHrwMQLdPqCa92GMT
85QEdzxgNUpk1+M0AX4UrBbjOiswxiysp/zOKoeTiQ4cyqfFtzDqqbpLyerk+ZGb
R06MTc48bW+r4VjTCb21nGp+paFYQOYZ/ds/gmRdpuua6NhQ31FcJh2VFF2mnqns
54/wVJDFn8y/PnHCAnppjUND9BNsBPJjhM/U1V8vMdFJvGPydGTLUZ9mLrOAzXJc
ZZ2GoQXd1cDZ8QF2MRaxYFsiIgNAOKB7oejSziocTth+SWPRXgEfuNk+pzKaGDb1
hCNDzt8b1C/ZycrCJFP/gxAj2O0OiTdqAClVF7AVAZkptGaC24f/b3Q7JJiNuwaU
TDAi80Zbp3vM/0Dg3VWYs/mDcoE1xHYrSjMwSxkdZMqnvsle4HUfukdEV6DJm97e
5idNMFaYSaldUeQslDEGRtRkjlFYOYr8BwYvxuQrLsBTwe1OA93oUdvy3bQuWVqY
zkEqspGGCrOaJtwUnXPa+AV2BISG5t7w3hvAEalDfIFLimzKqBb4EKVnfGueVt1s
7j2MHj4mFdqBJ0+hlw0vLksKUZzJqf4tX2Z0Fj3GKLoEGmqgJlBDoxkmteWOqkBn
FY0AU/JDG3H+JqcPaVJoU3zGB+7xKNPbMOT9JsHUdevcGbbTXIPgR+RWMUq5viBr
YgxISUuJdUE2fNFySsynmdOJbP+HT4WAlPx3+h7JAtG+zMKfb9cF14PuClW/lnae
FwtJcot/s0RZaYKoK6Jt1Zx5jii48JUwHZAKb55EWu0tGALf4a/2lq+ljz7ONZ5h
gc428kKW1VW4KKucNH0p/DJb51ZMrEIq9mpkr23W8zYqDuy59y4n0RVzEWyDb8M6
rYDAiWtVmeLuCTg/Olpj3CyjL1YM6QqcNz66Xs+TITLw1kfzByfVW9uJiTugB6Xm
cpZSfyz/zTJxJg7nxQqgZhgmJcpdclTPBMIF0BoeYMgIcF5BKyHiEPWHX12n7toM
Zr+YjN7gWKxZHYO25q+ph5xe8wPh/kEHIlF5A7znPEfoAXKSd2XOJwfaKZ4p9/B+
dXt2f22DpDks+FzPoTt6tfMSzdAh0XpqcwHNEglOaMZ/FFHWuKbcrhf3QwhBBEe6
3set06bLFOSV1vmay6BWRzsvO6Y8z8zumdpneB86QJC0I2ZPMjjLq3CBu/zmLLCw
tc30Ax1eiUhYTH+Yxno2QwNNvRJzYoKOUTe8/stYwLJKFbDxnnjbJiaJmgEDQiiK
+9NqW5bXNUJJSAqzo3PvKFPCX51/xjO3BQfYMmS9Tu5xEJa4WM+zN3gcVLbsDCUZ
oISW3yRiBYA6LKU1MByV8mx3fB27tgfj/shdLKgH4FvozjRJGXJypvAEw3qkhcWl
UbVD7r3tayIic1WLc43//EjlTqtjiWofJ25tbpalM8owzitcCOfUZIpf6aOunVhK
cktW2q0IWdNMb8jN7kxTV2g5OHE18Op6b0gtJ2St6EIP0z3STFGaCCC6C32SANdY
Gk6gNY256Hw5O4kwsY7dgOhUFRu1fXU7vC1jwrBJjo8VXcyFMaQY1zZ0saGyUJny
33Bv+Ytac+M5wzpNPQ+aostlVW6K2XVtpWbyyHn+WWi2wqYLdwwfA5T9vXLAw72u
nt8YFfmr7PAaGVbzZoyoHDXEx5Oe/US6osfQq7Gdm/JUvMH/NoILzE9GesR2kI1f
8ZQ+iWGMtwCv9j7fDmnSWvJY6KzeuswfVD8CKJG8NXJ3BNdd8GmehnRLjRs4zRi9
f8NuIUmCTcvSUKBWGcptZNdtymOUn5wVz8lZu7b4uR3l67WvFu5q/ctl9tJXOaSU
r2BbULynTUHsF4sG4eIyA7lZIu8JdvfXqeVDzb4LqK3E5AmKmfJ6wM18Jioft5ww
eTHVrpK7KJ6eCV1vqf+Ucc34w9I0wQb56CxLNgaQtIhQQ/AxQqLGE2i414mNqzY+
SfLRl1JTz+4ky/r1INPdBcyKy6vokXzh2n9i3lnY/HgSq/+GK0mbL/G/th3GQJ6G
MvY0cZjHYx4y29dB1knMsB3msY7kjyVDN6G545DMWL/lkluoYv8qtzXv3vjNYmzo
pa5JKdMcn17DmTQsvgLIevlqnr/quQox5iT2Ff9vzf6BHw/gJIwj9Yt4jT9u4z2S
NCKYfwLnNURMXbJtKG/qvNsfCwIeFSihVZZsPANoV8effSFB68RIyx/od5sB9+0a
RufFwJUq9udg00REJ9AX7uV99n+eBMxJCTSbc4Qf9NnWrJbCY/NG7+BycwIz35b9
EGIwPzu0oO76AjpfbPQQIghXScmrYmdVvNJpdlTzpd4WN9giHm0bAEWnZnhN5E8O
hrpVuryQZ/SxPXQbNhzpA/BDmW9vRHxuLl5ey+HIJyqUrOLqMwsxZG0jT6wO2RNH
vwX0qu/af9cgx0kYGRLAMa9ayg0wVBV+T7CG88JF8fzHaHNThL9VMawGcoHr1iwe
DBv9S0WUo4GqnEnBC7g7b1KXonucxPsSnzHRXo3xn7CYvVg8TqU+Em/6urLXzE9W
7MeGDqTGNdYDInmT0izSRo7FsKcjMgeTSirCVVLk0PTcJZEqv9nu/lxNhRYF+0EU
Uv+ExvFVPnQ+Uppmfnfh14OPWySiPBkokl9C1mGAqLh66wRboWKTW4qlG0UZNC9s
AoKUAVCaZpY+t0Jlv1FKgY3/5g6WijPVXlY64fNfRD/J0dURuMTsDnAUTmNVtgiL
Oj27f+6KadcvSDZD8hilnnmT9xBeTymi4FQaJQVKT+FHbC6pWT28PGI1vKxMAZGT
gFW8UCFayOyNV2dX4wWXTZgNrFT5EqYnRoifIemdQY70fdjfqKY/i+jAoaOLEQs3
OvpHmqaWUssH6o88nvSKGVFlYWO1pRxMMOpQ8SYBam2jiu9IP8KzRX4aRZreGx+9
8HWguXdo5U1k3jLp9eMXclmpCrK522Cs/RVqDtI/9gOPyyBn/C//U3JoZVJNHkYq
SVY75P9pnY02nKWSBWu4EP/AwmS+HEC+Sb5BKSwVIA6Zpv1AmisjqFiEnKvSAdkG
3pBMya0ib6uf/4IiIH8otIlzi1Oo6qq6EB/nank/8cKSnaCTH8R+ZM3hom6rrswm
Bc+3ovosokh958I40Ul4DzK+mgBGwd81kOF5y165LTothJTbOiUMatTe48cpPgEt
bKCJJoXygOI3oeYj6HBNPw7w1vbs85PLyKn2PEk+Xj4G29X1Qr4rHGZ+mMDNeRqn
vv4H4m8rvsCj7Cjt/Ax4UtpguN5H1N8KUcXjtEXSmCM9FXEZVHWVHW9MvAxacRes
7Hl16zHFnQq64BEWz3TJdKGX8dS4xIceZdEOI+OVrMyhIwHcteMYtx0FhUdElFUF
oZ9TJXG8uUiA9TpWOKgKmS6IP2+7q0EXP8azZCJhwiqJBRUVwNK2i9dSkyN4wY0H
erbfuEAtWmDz0HuSGAeyYJmxE3GnIqCkcZdnxjb3l8eM9oOSB5KQKzqOuT4AH/nW
6M5S18+WKkaPc5ftuXhdrvZVILX3N9jjsW0/o5cf45Po9FbdgxODUY/k+b0R9FJh
W+EAGqZjfUOu6R5puuqlZ65SZ54yAEFUcQmIMkl+6vD4WX9hlILLnlW95Tg1m/KO
p5FJWDAVR/KeN3OVQjuLtb6bj6ZY85DDb5MhJt6sPT8D+FUcKwJiAJPLur4BP40L
Rfytm0EtxXfO4HzDeYPBEHD/Uj6jUmhynRQ+wlroUHq+khAMZJhwPkJ1gzwuJC2Y
3GLRq5GHmP6XP+BVb4LEzE8HTX+b069yC82CAKYco51wr893KcdFf3ycJTOLk4hU
6692MwKucNF3s1lg3CqV/7YlcoKLTPeFdAzGZdi8Fh5SMcMbozNXFnhYV6Sp4yer
/QpVyRmKoBImlbbSjNGM7FGF4Q99HVMS62wToHY3/5vmo6EdMLtaWLN+pnzaaXyn
d3Hzl+n/fOBA1wSSvEBOaSE8Q/eyg8eHQMMB9/+JM3r66eWTctoPj+jSAhkiP77A
5fMlzFt31RQybzVpWe4U3E0ZF9YgrCYtACh34QN4Fjcl4bhtMI0p2T8jhDNxK9iO
oTS46i2zfNg9uND8lH+FzMES984EntmmVwVaZ9HJupeB082LHmI82HaBlaA7kHUB
RP4oCJTp+msbQor92lzGUSReVGUqY5UTms2jqvLarMF2FqeIgiORe/XP2b+bxCvi
jtgymjWZN4XfP2JNtb1MCqV8jInthdU8tu9pjroAoBDhzwo1NWb0dTcHUcksnihD
PccWwDL//AuCJEotj3cZTurEEOHT1DS8NlrwkV3i/9gIvJdykrSnJD0RolblaB3J
OGg6/LyuX2CEALAREJJSRhhlPBlrsKX2Gf8narpSnJA0J2MRkK0f9HMEwFWNyzWy
g7imnB6X8bKRynfjwIp7i1xpDusdQcCgecFGeB7aK/ZRPuoa2Fs0p8zxu64ZnK1L
5vLIKWXPWPSP/80e/AAJuhjCMXpTan32ZXKCxs/mI6BVx2kan+PBNnm2koheVzrm
qjfV9kMQD9hBH7skbQIyi/OTlOgRE6+z0cUD1W1gzNuUvjGtY1PPpNAL6YQe6IvA
DBtzgsTcFI53M6fEb4QGpF89UR0MBOOxVZSPBPO2vnfFjX39/D6HrrZYo8cdHidz
4j55bNDfwe7oxq4peBiNJYP84iIm/k36qn61eh3lt8g6plj4ygneES5T+4GNuiju
8iy/kW/M/vqUtuoswxCDkz++Na6rLGD4PeHC+651wtk+5IwbjUoolNCM3i/waTzJ
Gyiti0eBb823PC4MPINOoZYkifjyyxyZB0Xu8OX3esFNP8euLEWabsXB8zXTYnUV
vwabVW0J3szPUKALGGSdAsIREJ+9M+El0YqIb0pkrxQkEBKLVpf3kvEUoUat7KQq
2Gng10kRC7UpaiQipOpmjrlOJ8oHMpHY8yiNuFwBivSoiYDwk1dvNw5geFU+vSoI
HyI/OxoPbUwZdQZDZSgK2B7BaQjLxyevYtbk7qvTNQCfQ02A1E5MBrrAdDiM6xsQ
kuyS2hgRLAJTl/yHYOAaiAgJ39A9/poWk0QYR1FyMiuIYqd0GMagMpodOsJmo4Dm
BnNIuLa2HWabU4ZUbKr4R7No5BlHwJyOJyAhV1KiN2MWimNsEgOVp8IE/x/v+z3q
csSwTJspwibx+632W+HJA7ghTco93jpjP0aXNOYE3jhVcyZSnvrtuFqrHHMxcgjm
OrqA5PziWkUshvA4YkwiVHRlnvfEKfNqIl4mGc5hC8qRbTgdhrAU1ADIgNa27Dux
22RhdLiOI+LI0GawvxjtdS00+Qj2WTY26+hazQypnk9bLyr/YqGeHRE6u2FR/HcD
HUiP7YBRfIHXJIyBrDpw7go7csp0qSA9+WEmTr2bvklwx4P8mNUG4Qxi4eYTXkqu
4BLm7BO8zNI57IE8fiK7dHaTw/LMNKkTSjoP4qV0cFNyXu+LY3shT7j521jgnC02
pHJzliEBd7fGqug31FW8PJ272WvW1BquDYHp9t+8ejYN8pwbEyuuZqs+PT0racG6
eRZmYhWS3dEGbcsi4Dt6F8ahT3dfCDkBjJPNz00GMYxrHKS9lxf4RUhPVD2+dE7z
qgQCS0T4WgXTb8B+27CDyMEdgUdmAse7jrJkWO3EPUNHgfhYazxyW8LQL86VBD2C
9qVQeSSgchUQZRl6xGadc0fo7izMmwv4BXsHXTREwht95qxZZNriLZZ5E+SFZUcX
UScGO7z4WIQdAMvD93BSs48l1c09UAZDNNx3MxtPCTlMkqIVaB8CIRufQT12mP/N
wI2jBzUf52j3NdvXGmw16ktI5Bzy63fYse2+flQzp4CnSrhZozX2XjEEYc0Wwbjp
8GMU9ek2z0G0MCJUcmYLUiRQeLVGWmNmJ6Zu/AEPlCCCZWmXe+o4iqlWrPGAYHDP
rZ99iH19aDa3hOQpfSob7UwUq+5IViVGOFA0gn8rP/LrDMbrSNSKXI2CDri4Q55Z
CHNgN/ERDQaEjGWT4nJB43Cbq0AVbkJCkPozbNT1xkHVb16x23bRVi4l32309sjA
X2PLRB4EUWVmQopm8gfqPR4QvpC8dz2qQoL3Jr/kr1mR4woN5wIv869a6VQzRBIT
gNrkkgAhYnvLDCaHAA8wgeY+yj9J5k5Ijh5MzS7G0YXcZb+wMJ0QZ/HH4nPRSsdO
e/6Sm/vGFDcp4gRLW47NbiMG9Aog6h8vY48VO0XQ++3Rvu+EKw7i5yoy83mmOW8T
ueIckrHgI10LX9kdFa2Xp2x29nQqrg/pDto1Vk54m9a+MVxmIpLicKv/Doln//kW
VTyTK2SvOT9xs+DaX6e0N++/6nO2MXL3hX9VOTQ1ulBImJZwSL9EkRNFAqedrRr7
bdAAKxrZhUrGb1T/AHsFZnlnwl866JKSOBpd2UOuu9hKR6bxOdJkgmq8cgKWhYNs
VijQQBSN/xUnN00M2COHHyhdNSYWnZYX8aAtLRxP/J9MEkYGPcYIZIs4mP4hw8fb
JKYjgyvbqK0pWXRmRIhmIaYWMxAun68JGr1ApG4WSLTr/x+DUm5efdSSW7VcbZnI
07QdjotEsZmm4AXn/CygbqyDrAVgvfw5uKCyXfQIBaqqy16JGBjOb9f2/XltCiMn
u8oU1nKi/CHcPrv/jxy0wzE1LKHInHqAWJM3rH/I3qSEUWfiOjBTmnOGaBjBxzL+
dTR9eBi9mSa2UmnOe8HmnevLoeqFBB5DpskJPJs/psGpWl3Q/qiqhl4ExbryBZ0S
SpowifUmDVkCA2wbaV4lEDH+Rk0RQ1PkoXIRcjxvMCR3Lz1H0vm/fmWo6QEWXLrh
PYAPZNO/7HBl3EwSpx4J1B2R80F8oBeYSk1X7gEsL3hquhG28VKaaxtEUKq6FQDr
/I1qswHXcNc5qVeiIsVWhdR6nq4LegrhV1ZZwyBTq/oDC2hgeQuBLsyWDLj4rzav
2I7ooRc9tykk338uI22M+DSbyrKwYpKbn355eHp+pg5EmnedmTlJizH2lA2Ul05D
/wK6sYKeQdrvwE3pNgegSVJF5h+/clecQKUanLQfwTd7o5Wixylb1MZUfSjbXY58
85TYf2kOdccCYkdvHKpGYkVkU31lNz2dhmez6GXnaVu4b7aGQ1DeJTGMAuXiEs95
7hIdKl5GNnjJp3mkBsIjh/lQYNAzPcOhxgROuqGYxanMHwYcBH2bsM2gP6Lewzzr
5saj4yoZV2sKfPp/huAkTUIchA6jsFUT9PmUFyV6ZIGcnvZ695cei6e7qrZY1/B5
tOFh+cPp/Pm/Q6rvenv1nUjEB9kGURXye2esBDnaGLH4FqvrnqD2G1o4/3+JsZ66
3Vg0/VO+g0mthwX6f+5PiHV7Hf5mjicuk7SSPHM6adr5qRVj9G7CgYdRC46ZGACB
q6QBTEKnDr4Gb73audGk2gcXSTqDXhSnbloTXHIfPHR5NDW9AdXKrscJv8MoNpUa
FseIWlXsy8jZdhqQTFqJwUvG3/uZtP3EZrZ4p+kzseTCSuRzJf8ans3m451038LK
Vyf9u6JpOWA3Z+A3VjniBfFSrIaE8xovFfHcgMw0QvgOoXEnl7pgRgQZ7MfW2mp/
0QsFagsW/GWMgaSPRjC08G+Fu4XVmDLN/foW5xyKPQBUNOgpLGWdyONGtKN999zW
fG8DtQSPxi4k4i7D3bD9AJTFEIeNRkUQHDjxhDxSkpfBDZ9M+TrVb0nGNkGM1Q93
9xr+DbQRflz/zWEVY3JJNcCSncunwlp1gmkBpIyeIn9ncV2u+aTM9/AlGa+7W5gB
mgTPGGZGDXFth1LbwEmF5onDEJ3u2DVk/MgUAqWsObuZfAFQPfncOG99eTN0CYcp
GZuvPrnNHoUHWzVoUDRkGdGyOpjA3ioKf+PCecjFZ0j5zUTtDMOwCm4KuSOb7DmU
9BY8DovAtwNg7hwCA6d9DqPoRcIK4+FdGFicOMiBvHi3l5/vvaj6aypZN+cBh5wC
8FItVYwJ0T9+UDHRPZCiAAile+TNiGMiVGwVQ6ctwfuZIlpq4s/sLki1lShC+yRQ
9s2MGeDGqLURYG25PWasRz3wU5Je6pdOwMcgbJWRT66UTEJDhmsB471BGTbpmg7E
F6eg5KzkHWPGY+dy3C4mPyT3Ds6CUMv9nGaymfS7u/t1C5SBrmGuDw8QFMWvjrbN
k8MZUSSCw4K3INVyCctw0ygpo5A+mS5L9e0ourUhD1HRGwaLToIMDUQu2sUkW/1b
Xnu34UUFyKCO8oom9cdQNpOFfGUXnjoSVTPjbTyHvQBAhDNOyJUqtlvPeMgpRW24
NFmqx+MqVN+eglDSlvD5XPuhg7YFsGUGS9JQ4NaJTrGHrC7+mJlZck3mTjwMgfH3
b17ZVKtOgVt9QYcVO+XP28WdoHbaAXc0BLicYSHcAmIW7SZXhXAV8obbDq08g8kG
OKsqYnzJhL3Eorphb7xhDubhR1g77HC0Uv9OQ6SYbwAKzKZZRE/rS15wtvA/0RCo
DjV1u7DZscaaNe6jBCH+iB5vrsmUj0m4iy9e6fBb0Prq86WQHQNs/QgsBhf3aMG4
lWrNG2nJxxYtCyr9PtS4fWpO6WVWDA4vQu12Ho/mxlixDRf0NmV8YNFPEGfUqbA5
BSol7nvhOW/IhpQ4gNyuwYKZJgyM10rnZnkaUzjR5HNA6tcK8WhSJ3lwIIKKaF0q
evBSafg9lz5YbhkuiAt9TtewyvuW9/llPOV8uy6t3GL0fYfhduMelvcmW5oVh0y/
Y8SFD2rF7RDZsX1abkbCnoou1mF2S0ODjwqkndniE+q/Ym2RGpWB2lbSZcx0vlWo
3YVAZEfoT4b2yNRvx0lrtSrm2J4cQyL6h05NL9XrTtR4M/3HCC82iqalTS5TBMIB
inYKAAGxdHf5jNryjs+dOtyS8Ufe2hEoT2akJHHT4BzHVK9cZZf7nrYm6AcIHcuP
FK+WqGhO5tSu9HWzIvNeiMg8TuR0u+JqooglbffuHGAICzGFGQtFawhZlIdV4lDb
0Sj+C+y9kNe53rJHYACnlvBWzqDMszO4w9uQGZCX4BTdBdpOyUAAy47qudVweek8
HF8UaoQ9P+QOB/UycoWzzmzV+xmSJXFP1rQHB1ljgsym77JiUr6R0cQyc+WViIMO
t1RxwEnuJsciF/2DbBHftavf0sqI5OwOgpQfWdgF/PJytuiLhOf+QK9urxCD/vxp
b99A1TQSn95fl0a6S3MnSc01dw3Dcy0nu/7sbE2ZDUmaGU5m9YfX0q+lTRo/jh8n
zpWoJz0UaDNOEhRdLCT3UCeQFaduVnrSaEhLzfgQ9lOhK/ioiJ380mJfl8v/5x+K
qK7CD1t4SICmK4LpHzI+cykTIGCo4jy991Hfw78U5D6T0QFU62OWKNEydJ6S3SS2
kWWzhN4bA/4EYFh9pXHFQLJ1rExwYPofNPWWK4ul5FrkOplipFdGgMLnrPeHlWEE
jv/dy8prm05sv3YQP4KBsRs+g9eK0jg5Xf9XGYcYhc7DbRBfABRHP43M4zi76urS
y3rhRX3yc2VQ3nuLNtaMLlD/4IidIFrZ0U4w0j0bJOASM9jZWu9lbyT0apGFAJt4
PRgco1M8Xx5YPQUBKMw3ct43fUlVv9ESBWttNVvD+PyS0AfP7BMhfydfCBEisg5w
j0dBc0RZ9WF0j7ppzyA0YLCUaD4DAJppB1SfUAPadzc1F0Hza+IfyDi7TRnb5bzM
0JTddFR+oDYKIctP3OXShgvwQ52EKVTmI5Oi692MACCOc+z5Wd4tguBNmy3z1Km4
b433ZrlrrNfwZrP2yVnf5SrL/GaDJQXTMhSGPibp+Hwvpdfx44DfGE1m6FbHL4ov
R/cPl8xN+I4nhUfF67e0ws20migAICg09VX7lmd3L4Sem6FLv/7lP/kD4C8dGOAE
jDKklPhOADKoYsYWi/Ei5j1zeJJhRMzX6b+zhX/UF+lrhaRZAnyYa5kVb/3d+jWh
A4Fg8wfmYfAmmnYNSgGjPvTz0McTi1Iyu9tlX9L8/COAyiOzFyXsO9VS/bd7GiIA
VXqym2an10bRacefkKL/ZGvkGXOJCNlUwPuuouGWh8mSK+wpjwa/f4DGUTEbnuAL
zD1jKSaTVqvBy5AE3JpFpc1D0SVcXQutX/FF6M1vDfvj5XuwabD6LIO0ty5SZ31k
9t8zTO7dk+qAjh20g4RZdreVup+kHJtlGDaLGR+8Uc/bnOH5zmPw8RUbyc5cKF0C
htFVka/3Taoh3rqVJvs3hACF0r/eGTQmfF/d4AFxbPQB9FOlN9cx84QobrjPqKMJ
vQNvQe7lMK1T6DuwzCWKfjnv4ufAJd4OTJzN7BeYyP4JQVa6k1wv7ZkjcwKwQVok
8N6AQz8U275YxTsUJOqrCPG8Sw5uQrG4GauA/yJbZsy3ZqOwG4lAZZg/6erXWb4B
8Pr7J5Ugf3hIPg8+7p/nzpRpi/Tp612pheZVumCzxf42E2nCcEUd281kKQErtNO6
j3iP35YRzQfDTU7o5Av4ruGoGw4CwvOkQ8Uq33NF+rj9b36eLBtSlE0P6EQBgqWP
ggAchpy99ABdNeo3a2wT3VaN6X9UVfOHnrxL5rQfpjfBI+xU/n4/yfWhqZ5PCzyT
hJcWU+biaHDwShl+h4sY8bJ8IvOn/Zh4T0snNaMiLZNIE7xV5KiCKgtqST8E44Js
3Cq6w6p8zZI5gPUsAKCnzeZHC53W7ZP+9PhqSbg8TL69eYw1rClojUo+TJrylKNG
S9e3OKlousxJoSSritBFMMGfYR/hcc1vo3fj6/N6Zy4hp5K27aV4gk9S82TqL8jY
DSWLGVz7YFe7paBpFGLhOUvqQmEcXKPNbVkPTWLmDbb8h/il4xT7iKh9tQmKIEF9
GpNLYgGX+4HzjE/FFf9faQp2gRFKXV0EWQLm4oWnf6Z8fuHOpkT4ifQE0jpIt7T4
nDxtqxVw5oKdyEZxhiaaVmfyXty18oXAt6VtSdUDTABhrTPQWl7EAbDC2ynqu6Mc
Az4213ERosP+Mjlcp6P93yeW8fAZZUoEhChW6WgIFTApKCVHuDCRdJpkZKJxYQ9c
/4xj/o9LmTQFStT1uRc012Xi7zMGnrxR5L6t6wxuZlgUgULtkiS8BFxVBjd3p7LE
YkiMxUfYhBKul8rsjrH+uLkg/t9hoV9xqA2Xm4DrFmxGbtLlFGS+OJFTgyW0RsBC
Awr30cZdMm/Ru+8m2LCqBj/MuGN1KoiaAFZTGg84PXKYAP6FwJdjeEjB6+QTPJKg
j5wJ5GOF1de08OxwkYTj0swSHWLwb7PPBBkxyxw0zH1Z1e/Muw9TiaUbi1pTKoBS
D1TYj1dETisY9qeuzIjZkrEGbS+4/p7L+WImlUgTsSdD2okv7zacMz5x79MGdyoz
MLRlrmxlPrD1WpYPurGe2bJXYeP+SI2TvyeVE1dz2iIB2zw8O4CWDkIg3dCdI40I
wjJVtAL0p1AC+eGmUJGhBjAY/QOGxMvHSlyQH+GIJUVhP+a4GkYTwYLDPA8enHdH
BnYaOOiOAYF7s1Uff0QzYh9GVTS6AUTFPMy8menYo6CVXLMAskZ/ML0baho1W0kx
gNBPQudiwUwrfZwvagOjtcym4XMY/kCPvAB6qe5nUF7HN4gjuL8Edptdv2ctlcVH
DGQ3nMe6/UYi0DorAiB1eDrygioUuTiEpP8B+NPjue1cEKKUnWfbhTyPbr+Kk6cx
kA5lyj/P0pqauoGPVOgOj1NinnmD9EsRGChv44js1utUkhTMiLsp5uC1CFUd8raW
xlJusrxvEV23cIaQ7/Te0VxNTkxhcppfiVRJ0G/mtt8Fp0IR6PNdD9gxCxdwhAj7
mXfNwqfj9KTCset2WPquDtvpEHhut6XfmCQv48sHWg2Dp9E/hW7ARLHFjlhYvIqd
sXh1u98OWT85nq89SRAY6KQuHhbgt5SLhYTtuYCv3C0vMMUqSQhRALsCcpg4noGX
QFt+IVYCju9hiCdo8qGHEZtgMWac4EqrgKVUUUcaYQFtTMxdHrR2tXZu60PwaRbM
A4QNR9tS3yKizpX7aiNUf1s7GEy2ldzg7PcXoTnO2umt9BG6suI4yn7e+OZ3Q+vv
vqBqqP76Wc5Wb8A4jFPtEfpGvHG24+em8N6Rk69vL/eKttcCT10v1De+ABCLw3xJ
FwJmtZZvhGCv5CcRe3femGQpp+F/vyEzsnUd165SD6heGMMHi1nlI1lRfLvlevJ5
0YAGhnU01+7xoiRz92orkXzodZyF7BEVQnKYMWur6/pzRGoh/WDIL7Mq3efK8Bt+
+bD53KqoZbunHVJSsOvUsTDVKFNzvJlhGDyb3o6C8kQlHiVhZ0urn3ijIMxhJHdM
rcDUT5zVXofVXgcd3stz0L7v4p3EOSh+GVtO24CKL8Je/j/bvRbaICC3XKN1AezN
FfgopCAetVEhVKtcwEojbd7eL8YZpB0iCC7EU/lbHSLhbacuwvhJwmIsqK9IWnfs
m8K69eDSRgmUCtGzvW4LnorVuI8yJLNiCSkLgtz1l8XgzE/iaEVhUdfwsKwcy12l
eUObFO37hgZ/t602L70rTpVGmJfiLFjAK6izqswOvLHTnyfJNr2zfOBWqqes0Z6I
j073xO8AcLL3PaGxLXaMGl51ErFu198isaRg+h8CVxPOVegcVXZBF0n0LwXkVb0q
aCH+3NOx/CE6nZNZOx/cgwEFciqQ/i6U1QmPHiekKaGGWetaEJYrGu7Ajqi91ZgQ
9mZ9KW/Iq5EhLe5oM8LTHObJGcnFQyUZuOb2uYPm+WiJhra9pgW1dz4jgUNDvPgo
cVeqf5uJF9oNA2/JFzOubWZFJJpO2LLrThiQpS2SOhMEf+tbRlDmd+BRt2lGrmR/
/mGS3ujmgmL1to9ICTcacMtxMqPyBEKFvuoNB6cEUAHDMYHdqDFQf//2jMNUQ1ME
q+cgUv8932BpNYykGygUGyljpEby2lHpSj+Gf4wAA9JrqMmuPXcfxJKyhGI+WZNh
4HjdkQVyiTzEci/qKbdp5LoF8N2uPNggH9oH+nhhD6obtVBH5KJhXjVJMUeHMcLn
n+PMZ79PVk8YpA2y/MMo7loZK6EVj6FgSbt8ZV9APv0wYnMw2Y46UZ8rF1ilIH41
1Zy6F7M/FMbFsLnuYUFcb8DamTVDsgxBDjMphXy76iZHp0Znwxp0nFR9pkzey7b5
K0xi3scph4tArXQkIPij9a8QXaPfUa8yYB9PuB3+7AHhUGS1+7/8E0AXkGMN9Zc9
CrVPAjett1tCwPIA5oKuJrHFvITDc0zeXIHNChR8rRrxHs5462l6GYMtcSWtBKny
MjV0Kt/r1NvKN1n0Rj120rH8vapnKjJi1j+MfF/fT/S18l7iBeW476uBa7gAijx2
FBtFm61jQ3huRtnEpeODCwTTZBtwYy4i40PsI3tiqQEsxRIRMY4P0Fm4hur+1XW2
tiZmIn0nrE4Pm41Xq3ABxfLQIOO0FNKH+gKCjCtJIzf4fC0S/xqgUbSko/jRcIGW
ADlRqsgXP2DpVSWBzXe6csBv/VRBkpK9/W+DBERuPofBEh2eNeO/5cjOaMu4HonE
TW260LMe0cOvOci8T1b5VZMlpL4v0cGr/uRjnFTq8ewugVp6QlHGQc6KB4LfDw8U
zgUzJSWK2s78RHsbiD5pveKtyQPRjckzx5qEUsRLg2D4ETUiaOOZ7bJ9Gnt4YsW1
PCAFeExuh5IDcuzzWfxKGbk8eL7Do334eQGvbf0vCKa7J3q8/+SfecfIJ5CvFxS1
mIhkVzLohbOn1bduWmAqGks44EdgoJzKfLE25M6iwTDhEGAS96uW/wabGYx5hLb3
wI1oMzHuJ4m8A1/VsI4AGbKkykrwOK1woDxrpI4VJyo6FQdxfgUJkSJjemsaL2cw
+h0huYYOr1ZfWVQO0KoQgrY67rSoOnqt/ni8nJrUTzXUH3gSK48Wm9/UHks1Glk3
BlV5aKTp4DxgRu+6fbEW/61iCrEtXwbfjZ6d8BCg0l6RHh+xqezgIg2tcHhg9Z2n
Pvz6uXD8+JtN7ECqhCR3983h5LMDNV15vKaT4hIfsf6Vn4CTXoNWWXIYI03mLd3N
DV0ch5KTjOy9cEHY+wOxuRLSlk9UY8XgY9tGf8SsEFKV8i65X9JihRq4+nwHtZEH
sZ0c11bAWfWrtTqqddjcKTOzKcM+jSPKKjYPci43yj5WWGOTfmXDFjbTditZtres
KdMsk+N55j+9ne74Zz8HkTYEevbwAoB9FaKZA4s14wIy6814lcPP/7NMH9Z+Q2aq
kbErCRT0f0srqu3niTTN2/JtLheTCxEQAcXsLxM9HbIMmi6ExshMPkpLrYfGR4dq
gUfoIqNjeXTRPOhfAsxz7OCF8ppHkulo8Fdzh1ODxOZ8o3pufezdMffHxGIs0gOm
HfYTMSnYFj9+ORn7pd+IaqiL/CHxYGsP/0XxT07EcVI/6aahGmBra/sgmQVgn8tM
SyWpC+uLrMmxlKOhCZDT2M0ovHMIwtBL8z9R1tCO5fL/GxumEyRCYl+tuo5DQjdd
a/SB1GSYA2Fe6xc4WS9DWLbM/uXm2htYDehj6XVJKXemFHAaU8wYkUL7CVbMpf0M
GWuEBFF8uL3KacaSinz7pfr6lbkBK0dVY3sMB38oAecHTCxIAnY4WH2THnJrGyRB
O/q6JfVi7fxsitW3Vl1xIeG4UPtL79xLV0qgPVU40lI7svUoE/lz+lBmWWMRDEZr
IbKcTSzJTaadCTckynozsTzGGi/uKfoWpz+Qxj/VBx2xp/Z1XJ6TFooevCWDGr2R
jrEgvbSYF7Eu+OhgfYfJEBeMN0PPXsMyutgtcNxutoGAR4rNBcYdO+5mNaAZh/c8
4E83LGIPSkRJ2XNOjg0CRmunS7jPtqIcVRn1MQw3kg2WL1lTU1e1rQ2LD9kWsTuE
Xi4NffSLVr3n4xNTgLb9FMLGzP9hTmUKTKBI8qOFG0JlmFybwSdUp+VLoOyl3cL5
D8DOm9HBVJbf7oCW7TiPL7Gzrv4rVBXxhdxanTeeQj4KWk55IBqTVjL9EdbiwK98
sGx83tE5JDrboHIQaYYfX/OGhiNnuBaCzRSYD59eQQXHdwttg/FuUV0LN+/3Pc1R
zU6SlPoVdbew4fm2gXk53ls+kodlaixkAl2HxF0WFLxG1fFJwY/HYrsgPdyqOYbJ
fOl9nuWmhnLEXGtrBLaKaeJLGzuBmqqUWLkhPJHX2MPcSdymDZhIR2uYQ8QixUFi
x3ijsyPxO4ztOoSc2YJ3gTYn6hbl72tRysS7qC/XZfxrF0W/4YcXYZdBIn1smFwd
E+geeoPaFp5yN09CU556hn0R2ffmbVRFaPgkiWiF4ooB9RdBu2QvE+f3wUzeJoCG
OvjOMpWgOWIcsb1i/VNBbkDO/4HJnCSGCi1PIwSOMFNnBD5hiHT29IFxiskgFr5y
XW1/u4q5SyvOE1wQmdLebt6OudqnQdEJjQMPESthzov6DuE/pnm/sy4c2iJMBRA2
RMDPU7jJD5k0LppGPHzqKJj5alVSYUGC4/7zQM1ZCyCU4Cv+BfEmrDRavkANJ+qQ
nLFRoPshEI4HFFc2p6geCuu7CXfJgUzJspN0OTjt7OCXCfV94rLdxpoqsywUMppm
uakr4tzbCVpnx/rwJRWFVbQajMxxBvJ+h2canyTe20pHhIYa3EtILWT/ha6FbDl+
BRiNlsYP/tPyMl6NeCTcDzVTo4KzEGqK+oMV0VIXTeWRwSHj6FctT5wstqNO4u+I
j8C06mCyh567uRaSbOrDFBuGp6sLsN5K5Djc5oBsMlMLpsydA9I+gIPuX7I9YZqe
Bt84o7yN+di1R8OIlXeY6aV3P8XPtxEQWmsZPxDGoS2AEWTbY096DfNzO+D+x5QI
p3tAMRZzCA12S3HSLyvmUratseAK/f3AtlmVnrQNMhbQorEMt4mQwBBtkvKIQc6a
/7jExpwcj1Vk3aS+j2AuFnw8MdG1oR3QZmqn0aNThM/phFcAeBv97gWWHvmbJzUg
sboen8HHGcDo/ksZApi6quRuaq4iScw9oaA2Tc/hCgSL9ym/V8XZ3t/q+WWEAiAZ
r5GpB2SSwDOlGs83FAy2VmP0R6t/LqNeG66Hrt4O9AGCfJFRPspCPFwLVHUfztfo
CeCxDMreh8XbbADfIIR4AFKIo/41G0DDbPMS2YTEwEswiA4F1fvl9HRWMLw7NNyT
3l7XqN14/c0PqyiJyjLhJiR835rKJGxNa/G/K3JcSN0iut8GCa7gq6H5Xp/gRdhm
glEIW62uw9Vm+NEpMaqcoassoWuNxqJwRQMvZELe4QQtCgWdVtzlNGLvow/wwMPv
glNLYBcM/apf45RYMBbR1pYGma0KQVVjSyILzYCkcMdGq35EcoIBkjZLj8ZBuN9C
y/XLKKXrBReNbg1SOuam0Okqi66bQ8gMls3r8CjyQ4/AV50it3C0AqfJ0kIU1KD4
sP6UvvX4c2EaC5tOo5EojDibCMQ0d2rrdS6kLOoIEF/E2F7myKTSWoxQTbvLA0KK
KNAmb/btf5oykSjYJd9S33Gf05SPuHJYIyoSkN8+3QVVjDSxdyX92CdSTotKR6ff
55j/1OfPpjl/a1fWzl7EmgHS8DIvgmeQPOUHDQqnaCJGWTVf0oTswxYoQ867AjiE
ll2DFWaj1ufoeyutIluaG82o4GDeCNT/BrOg/OsyjJpCm5r9TFwn60aOpJ4pu9cz
Q/FlMMZv3Mtz+V3dPD3f8bjih1F+ehc2tDirVdVs3bOBANdMM/lxWOu0Vxltj4Mf
EPBJIOsU0b2OXtmcxTB3fyCCRTpqfPznmMggXWpjJsKH/NG24PhknRpifs5puEQf
KxkYSex65+dTdzCtYpUulDBqeOMcX1vUhtKnXxNvLafbLB4qo4j0ldBZxkFIeOBB
mAxGqHLk5rJdL+0ASQ/ZVpn74kVYzVNasuXW64yuALzSzYg0JL+c9JOkCkwLprr3
RK8/E6YvDKm0Ab1aXxgMnbtuLEqelq5N/2vi40YNQnHmKduDcLFmxtJ/bUrj4p/B
UlR0ZiLmt7Ptq1ECIk0wvaaBfHbPrg4Tbr4oWfsXrLiSWyRw81q3vDd6YG2lWP/F
OYJJECpGl7O/jhxewjCHEF5mbx44L4DvQMk7tScZj4yfI1PEhdK1YBpobszv3zLX
UG9frfw9PdPbJrSa3lSpz9X34d3qLSVzvALFXHZ7l2IWsMLR0OV+SScQpcOKpDza
ZDeh+YnE45Fg4fCCIVkNGjtisOJSu3vIKYkOlnNiTS0Bu+MVWzk4JPSsCLWKmdLr
JAL3ERbYfx3uVN6J34OtNNfHSkHeS8Su0+DhR5dTR/8t2wwWqQUxMgcwNLCK8sEq
PkD8n+WoM9yzMSVIGywgKncgpQzwLfb19a4UjKIA/MOR/0L/HFGBKlQ7AvbG+INC
FlesjIBL2CUg673J9NdEKSbn4kR0jari4MgdRyZi3KKrMh22mzN2VrYroq2Rv43K
PdD//gFt23p4E5bRw/KK8SVqC0drSPidMFUHMOJBm3mMlULjOno34TWKW2tYzdqu
6rgBkmPHBegE7KUv9TrTUtCZeOXZKTpTPRiI80EVhVrJf4BYocc+IheKgqYP5LOB
C9rNlxa708V8er4bEQlQJwAcf+sPWNOrSqYCntw4OV+8IWrJ/FE03J5jsr+4E/YI
SQlkoOuRoxhi4ImfB3roUeEXJOYT2LpUUKxS9HBFmHLXfRyFOAm8gOX9/valtV11
g4lmJdqTVrT1OQbpSdQXKlxYci/1cb5SmwHWM+aGJWaJEAGo+JW7747qfaKF7bA/
ehYbgox3d7xkSX5inlXVYm9b1LfeZ+3MCiBjziOMS25Ok2Of/PIQMywZI1dt6ER7
d2+s9dDrcNicJHEbNnfFVxv2Wozr0/GxSZKpfafkFcO5klIMHkDn8rxbpi3u50bh
JtLvhF2uWVYmAcUzsqVedQGKE1g7UC9ykMlPD73BbJDZCQOJm3WzxSUoknLIc7Yi
rJPgfsp26TAD2N4sNjVQHSpNKqfQL3Hwg3qBgfRavaWuUsdTu+SIG4eKyUhMKzYC
1bC5emFdPafn0jbJIU/ja0xQAe/3SzCzg7Vc18RmjAAJEK2mImf4Vz5P5Nf2TETN
3ZPgLeIdLMoNe5nndaKVgvjURAfDcZZNbnXHmHerrBStpUPQWfTLn+ADkBW3MgSX
CaQ7PDoZEh4G5Ewmwr8TfPhenDy45TzsfvWJl0eqayJBGMz29pE1JHx8uumF5K8L
HfUZBKGccsOKZFPl9FgDUWb1D2KT0hYId42OhvIrEZ024gAN2Fi7ZPwBFkY64Ker
zb1dIRxDpBSrqxuy8CCMuqHfXcLnHhTdzcumufcxjtgKcgx0+hWFh/aJPWzUxxuA
6DoVKB1D2oJPJa7NEGt8496LiiGQ2fTGdYvDFVYymT+UIJ7r4xwmxp9k7PlnVbYt
F6cIdQNvZOAKRNuLQsaL/QNOqpJCMcK5W6WiigCtTfW8OmQTvq11Rxd1vdQqxIUv
88cv3f+theAwig475l0cfvOMbb7fUcRn1oQ6e/qseBpaoT8dSJFLZEXwKhntHwD2
Xxn8vvnKtEpMuEkvdtiyImynDIpqvoLXILx78+CONBFnHoVABl0xz7he9sGdD1v6
2P+tAGAAmnYzE0tmFoKQRe8CYRopOjy+JBcu5ZOXKgkEuEftEPW+I7tCiE3HE+x5
bRGFNJjWme6vojQkvG+DvJdfOnm+GKLkCWOcwg+W0FWjzyzfTIVnArOX+EEzhq08
GNQSXegkHCPahxN+aY0P3dGxQoaqDz+Db/4PC2aHjHS/iGd1YeZW/9+w0+jne/sh
4M0sYE8iO9zlUkGu3Pp+6Ype4fHwZ2m92TPjOntDSCTuC31sQeenJeaiVnV7XSdy
hRoHO8/Kg3gXp6R7Ss5OYIg75R03HtonARyLVvvsj0dksNH/mkkrwZwp0TSfj3mv
xJQqCoaYP8YLr/hypnvN2i5b1J+hfiaFXYPMP0SIQMA6U2cL+/Tv0Ulh+PKj5peA
QCv4tTrHEkk5xdkOE+f1xwcQLYyoaFm9QYx7XOVIPvl8J4x0YfNDIuOPAoKn08d7
zsz2tJOs3X9hQBKWQ+mB3FAPF1qX7e5hfYwEzP1+IHyRcPiizE8h/ZGGQ+5L08Ba
V55f8U3JC6kCMwVxWIg0RYj2cKnxCM+FWfiDyssWEoF1xygPIuQHb0sBoQ6Zj/H6
XzYQcl9s/J8srdNryt5kcSPxQdKVniHDqSHXCy4iLG7ChCobOqRUzUB1H3vHTxX8
zv+lNzG8JMowcuTDMvsoIV8Xo0We/Re75UwO0mMd1mKnlqbIaBTOnmTGL3Mlo0Al
ZxxIT7+Yk44pJ7luqpWbtUw89CAOZ1XISSZf3JXkZDRJN8c4IDzJKU81S6H4lRjZ
VsIEZBO4EwmFIettTi/7pNoXEFzrCqvu7mPwb6Uu+Sv3d42qywVLzXLz3iQCCuiN
LLStZZAnQK1RL2ybw1aLOVZ5qUJ48CtbAEG7z1NutI0FejQHdv0XSJqNY6jesuHm
viyLL7b7JJlBC3Zj9BqcaxEcdbLVdLsapNIFOmqljNLXrkaIjoEOSqwh+v4hOJ1g
ucvlUa+RbXq1qHGHLVw3jFVRenLpmjfiE/f3q3m26bLWtu7CRkrg5lSwD1XU5fSJ
XH8ypHDaVzIbeZd90LelumuHTe/aklpDmSVMmUM/DurRCiYHEUYJouYFIr51D1wM
vjdNlHf5neZVUSdPRb5Azng+cdlOTGRYLr7C7fBZxAgOHj88m86m6U/ekP07jn6p
g6W5ckXn42WMdh2tAbz17cdDYBAZh1V/kutmGhQreGPp8kwzk65/s3XpWVTbGmm4
d5DS50oR5znYkXKv8EboVjjUISvzwVDMajXsId9EEkfXvNgY2+w06SxQlqKySTD+
tXrSlfD91ShupG0WJ+whBtB3mApVvF1flMDbBMhqJtyaJ6R1xlK85hwDlDhaBNJS
TGmnGx7cvbeisgcjGg54OTSSp2DksChyeD2/+pPT4eQ8cK6V/iroe/KF/t9F8eM5
AcmSV5XkGLTXGHfavZlGWpx9QRZ3K7lO1HuyCsIN5FAfql6ogspMl4h60ZzwNRrt
SdvlX/M7xYPReheZ4Ngr3BiyOAQK5FqrPmHObvLuujXpO5R96MikZXjblLP1/1el
a3lE3yItY85ALWLeQs4blV0AsXu2uAN897+bouOR/5E4dGMYhB9n0iyJbg/uP9Yj
1PQG83wM7ptvax/KqPIbcz9adSIeevMgRzN/XmtB9DtwwxkvArzhBNwYT/6xftMv
pTESUAPcw1J7AZISOrSUieHyblf0R3uWmDfd6hVAnzKw9WgdMLuXM/ZueaX23Mc3
82sICRiTdUnUXj3Wd03wGmrEBCRCOMmxt8a6tRJhJORxPsorLkg2oeewTfffljH7
so5Ak7GCXsHYjd43JCuACNafSE+/ov2V7p8QuOzsGEU+gmGaIaKPDc8MvhzMnl9M
viZDjiFt1Qi3/V+WX+Bq3cYAa+5Iu+x3hnbalySsgf9DrX3QQo38qP+5n9A5gaUY
NATc0wzxG6o+e8jmdsLoG0QEpWZFeFW4x+4ab3sZyty2CagmPZnoclPGfYqUoGzM
9XubAw1o8yKnyCew+/Oc04H4EHc5zOYCP9jzfPgVslm3cZL0+122xA3DwqmzL+yM
H2eAPDYTF/xYmHMGkqfSpSZhNTt5Oc4vgMOxRvEGeZVsCG0r34pdNUmdrOHtlz2s
F6e6j5ncdQEnW0lkmUDgz9q0iS6kFucpT4tqgMxNTe455/OM+vyTfrGhUz0cpaBx
ni6R7qgrBfw6GWkWeEsphA0XNs0wBJa9NnnJDKNtkxaRC4patx/RhlPduyXQcu8a
C8yLEMLvTSx8D7BdV6aBp4dJd3CRvglHjUveQ7Du1Zosb741ts+TnQ7AQoEHb5Lm
/rPBiJVQ8VvLbWzpcIejpGjG8FtnnphqVElLmOdYt/VuxT7SqTpbu1URdV3u05XD
prO3aP8HbUqN268p6CZ5FpTBbL/22yFDE25kjg2J+skZO+PoGyjYTpZl98YG8v5p
BAaaFEwA27yxcKO6cCuSs5ZzzRi8qE1S4RCUxT4OWnMwRyq4hLmz2mbfn/nYm072
Ib4Rq3P4rHZ8rF9DXp1WCvxyl0OKYFlmZMRuDowqwYCuTavwzOlvPUNnb0hl7hJH
o0UGelrkdxDVyC40ljsRK2hLtp8cN0LpByBr9qh1jlc8CZVADrDVUl8PNBP+jidN
cLzkcG9OEmri9eqouaWj0S2GsazlSi4bHdomCz5RKTgOqwPqDhwO8rqvgkthl8RN
BdD8O4IbCX5ZFyBTd7ornbQD+ZjjW/v6UVZ9rmNuZiPw+gJSOF4zajK5T56a2O8T
VJxyhwM+q5qyTLh8l3ib+vAEczeH4obA85W12lZMVMTAQnNHM64D2x4u/54+tBnK
PygrLOoHeL0iz2x2xAR8D2zf0z4AiPfOZfFtl5hEc+eC5UmABVUy47skmXug1iNK
vIbsCnTpcn7syXk1gxmfdakt65mG5RwmWOSa4hIGcS75M0KG0Zyl5BA76V4cgifs
idNimOCykjccTkg8yHrV7IG4nIV8qqziNw72XKaHYRVWXm5JWOe0MudLUALK/zUt
V2vbWX3iwwc88fBd2ZY/Kl0MGGY4Q27vbuZdfLvO7kvjWctthLGhNNBP4erKD+/f
3apDLDII+jCy1DdbFMfDBXrD+6o4prIUXHzDl32G11gIrcCoLhc8YTQPYvXFauXC
6Z8qAWxXxEzRizSIw69Z+D6/cLFa0hjLPA+1DzkWi2EwFlOB8r0TOqdbl5INvpjH
aY2A8IcPZkDaeouhP0j4yHPcXo6xFxHR+S43EFlKbR4h0wmUjuXN4evgbl98sEuB
ymMMbNxW3l9QbENG+GGIN7XCzZxS+Wl6XR5yOK2VvYsYmwuhDDRqpxmu9xlvE1qz
oCxJ3eAM9gICYcREvc+jKg9WVZ8yiP9SlrjHe4jTYt6QqednQddoG0dCF1C2Bx7c
Q8vRMb9ahYS/s92gJZPws8DBk5YHJ2lQEZlYK8Nsy1OljpummEzXcD7MRX4PLd2a
9jjuTzjuPdPkOYPRorBFQ+kKcfOh8CGmPEPpCXGyWjHvib09b6u79Zg9TbkSeAqH
S/EapDuRpUWfHKZjAb87vQLrkZqennyOinE/3m3TWhexScgIE5aRHJT/NxtHd729
MulwqvoMd7BiQfhRf4s94Ug/e3QLfeyYti8CEEOGcvttT7zGtq9/gB5gLHVDMdPq
Zl9Tzy1WOuIymTWbjOh5Ch5OP+3wwuJ8JktVfOBomEzc5Px0nSFk63LzPBNWrvHh
fUZhYvOonTOBgbQWFbJV/dWcIUGdvMR319eEjI3fKUC5gjl25tNtMYk0qPmqeiSQ
lRiscIpfAGltMWakNY1O6F27UmKm6IiQbTSTT958GWrjYZOwHzguwq9DkAExzy8V
qePh1Smaq4MIC99vV6SaA7gcvykyysSQQ5Q8cAKfZA5McYlyIR7NSyX5wLRnQfKR
gk5WmsAO1XHdjzzS5IOv2WqVUmDjGSBVZGKKAM3Wr5+XKE+9kuvHG/7Dotb8hhm8
n13uKckSHWaBPAh+BBA4O3Ssanr1+/4JeG+OXpRpTwBHs9SeDq9qdl8xzqkhxo5r
ZdHQ0oT+PbI0dipqfduuCOTYOw+nogwoVJq4n+sKVOMd4r3Ok7IiLgZ7RL994eJk
DTM48+UAiFmisaJ4lb4MZhta3CZ7QAs79mPf8i9RiG1SBiypQtXx6ONPD6qZvxnH
XwDj2tzc5nF3rLG2Xb3Z0xBTvjKudtYybDPQGNGy/Mm7WROR0gZkqaCMTW+HWWKu
fOtEhORvD3wMZYn/c7cLgk1MpgIBw+yNR/Wp5puhug+dmxpOWuXIzFprTHPksFjp
kc3U0/c1W84lvHXGY2SJSWlytrJUPnuLVXRNc2VL55WihyyhBHVq9CA+GHRqpG5F
+8puEsUl8SPKLDW6VCU87zDEGPc0wcOc1IRWian0Ucp/YYiUz159JnoSmlyU1iQy
FPc0JCjY42bLzGW61OxNdNbkPF/1IQev86SA0LlXX70xGjam3KvbvZT5M4YP+RqG
25uDOdTIOssCCBzSwgR+yLh7DQEIZjr9TGLbSoBt6PQyJ4M8S1uppYV3pMR67eHf
0fVwuepJo980ZUgwTCgKEeh2c9oTY/KMNc0K/B1tMYwNocIe+zuTU9M1KLW4Dvpv
FnOIu2DiEdCIRrAgURC2R4uuehUJhZK2iVHEhuR9eTWApSDpJd9s5434ptVDEDM7
wMnlnD9ggRl4OtVprD/mZvd2Ga/+ly1+7Qxsak8GU7ji/JIVNUX1wJlI15bhM3fy
jmx9tjnmYkBMnhVl+5J2u4ia1jVY6sQET5WT4XtqgjCuGJKl290L/MFPBaeg4139
wU1Y3qjoG8Bx5oJToE087N6TCVaXy0du9tNnOB220GEPCxAdH/JMw1YpjIZH38zn
xV/rSlOV4VmSmK/XsnbxmxqFYIVd4Nk/uhV5BmTDk/hCsYMMgIbWBQsp2vwi//hb
y3GlqypcfRmkMuq+Nvmcy4kMW0mUd6i9d4rcVqkA2B6mwUVcUrLVjkHSWs8k9HCR
nyXya787il2AjPC2QTVFB3umA6UKXwhgeoZncAnWVd+cAv/2kvn3UXPkYkEAFi59
+cW3B2hOyACcHb76dnBkpfik/r4wLcz5/mtB5Cp3I7pxFQA9AvvhCyG0kiRuIWUZ
Cz7A3XdtC75ez0iqe1BWGbk8Fz6iJc4LKHUvmveu0nlDR/1/d4uTFjlyFSMdfpw7
ag5SqxqNVk3eOTCHNiRoiAprYnCYMuLF5G1Kyj5fIG4Y+i5lTPbjJ2wmHXqIX9K0
T33UCzNAgkHi/o+YiVjGq7E0NnWhXUQyZyM6ANtBvE2nD6s9oXJ9AELNVXnF1F/k
rPEGB6uNPy1jH9jFyQC1MDUNsR+yUYNMrxWnizes1FnzFXyxCQNdTyd2FkBgzpR8
6DCzn4hcFhv+64QSRlrai9GVA/CcWs/QjYsNnr/YSU60zl99nWyPmQ+vlCVvE4pZ
1i6hetW3Px4LQVmz4ZHJL7yun6XJc5+Tmz+bZdtGF/GTKxLrJLCRyQOLBRewrDhZ
sDUH17nKM0I04PV2OkOnqz4kj0/Fk8GLA4diZOZK2/ub4RSh25cctUYJ3p/eYqxJ
Q7xEoyExbw9eOPGSqGyCHPtj/hRljSpBERn9Yj8iw3KTYMqlAqzid9RHaVlLlqZc
FH9/QIECg0mQKzJovrdkiECwaLZYwZ9zVUwcQvWVIFXtftfhsK/dxkx5E0Xg727s
C1YIw4cf+OKdrcvqlJ7AODrTlvjOHB0kHsau19+9acaR6A7gz30LQCYD8rxQlvlQ
/30MlFEkDpsPrD/xE3OxIz5NNJBfOFfoLKq79+mwE4fLAWZJcUR/Zw2AYnC0GhbW
BnLfQ3WsPeg0qyzgxG4WXSxU+SU7DlANmcTOtB3mF7pk0YwYbc+fqXOY7hz9wflh
bi+oaDwdlzG/Io5XIh5o4yy849ce6rg+CYzybM+riX327YyRnapWUSzm6wNfznuf
cYfKbruK3JRvTGhkMHNPjTTqPsqd4rVpblU6T86dzCInc3jOnavcTfvpcHkYe68Y
UQTBq9Y+1qj63zPcd+xStRM/USBC7VhKFs4WinLHNC7gL94LXtOMkxSoAchGoSiS
FZwuQcLs4TIsjDhHK6xPnGnDWb4xit1RJQlmTXJIsbID/iupjVRJLNFUOryMuDUw
IRlRmrUibSfNeU2QEA/hBjm5CeqOJrAcsfwJRFHvcNNB6LQjmQRrVestVkZwberY
cayLjiubQphmOKHi2YEj6jbV17W7At2b7g7gXJIjrdEAmYmeOAMIjvTCF/84G0ts
4VYkwLEfs+BwMfJLMYRa5VMsMtRMBjRKwBvGit09HGBx25qq9XK9JU6xkS5sHnVs
yAaIdRamVQCjuvexuGFnWfui1pnm0lh5AMf0pY3lOANSlSP2dzo9at/Oz0nTD2WG
U1g2f1nbRWBAgSt+LwRIdsmC2Qko5CzfNl3LF84/sh6sjOSVgorpDw6/3zsMBEOx
DnIDaQOiJyUOIEsZB/tVtXNg6JYMUMnIV75qdnIug8PyyO0ei38sKaxQvBBu8AiO
EcxtPvCEKaCZqaLtkctVU0YXr0c97wH/quxN5YiyEsWaiSmNhXbpMk3I9CEO6vd1
8Ds39mCjA91GA5Ce01bzuOp+6+z/XmRg5r6eqnAlD1XgfjHoNf1RipzSSPu+uGKx
wix9ZQQ35y6jgxWzb/fnm24y57KRDXO/RpW7h0EJ/xwFdaIfKFgZQ/kqH9USMoRt
27BtV52nia8Db33C3LWU+tG7MlYspYxd3hdeKh5fZ1xxEUy0AwFxu4Jh1FnPMPNk
zZ7u4tgjTrVRP+VUC6X6bmtL2I8PZA4qa6u8MGA9WcvFmj0tcco2NbMJGYYTV3rT
raIiEn+0qkeIC3QNyEPqLi6FRSnZcZEX8sifBl1aiBK/kkjHEVBlG43wEKH3voIg
1b1UiOLmw+hqfLCjNi+QRpXLntt2V7276cNZkagcm/3U3JYCGCYPWQ9Y0GkKjxT8
Iv2zHGQDehek0NUrfFlOHd/u/tMmQrAvJl/N2KsGLqCINkWxQDtxvCFVf6Ohwk5z
UTDNOT/6Zq9ja8VqFa3yty9msCKHm64kVFFNFhr1q5+rCT+HyKvmj6XZPiZejUme
Hb1rfU+aLXfFVlNRIPErMmdqpme72BNjtGXotEGCS5c5GV6uaYR9p7RETQejxW42
zf8wOP1ZKpKd6hb78dQzUsUaqm+WTmqv0OK7Q7QyQct8JuCHEqyR1Jcw2pK9KTld
Kxf7wqzRSa8SbXonihq8YLopj3IJtqy16eecz2DWstX1UqO/37QSD1BBtb3X5vS2
OUuCARxw9md9DsVNqvw6ym9f+o93H3unlMyrRIHIQL5cm5H0Fpe1LnxS9d3N2XT4
0dfd9u5Cz3XYVs3npoXjsGGgz7toDRMz1s4hblYRXGLJITi/jTgRtKtEp8gu+6iP
pO9j9qUATN8bHUrqlaLmrPnQAvK7YoV3kB3i+COPqCQ5oNrIRjN80Lofowott6c2
MYaGscwFtc5zGA1W39x3k//1ohZagGAD3lYN396NertaIojrQCRIDJRtXnZ+Ucgb
DCPUYiHO6AyH3HvRH9HSKV8kM9L8bBFbVa45xLqTGPdasR+QDD6UvJEHBXoUxIhJ
MPt6cfHUAJMWJxBAMe5bYo7oNEsK+tSbuMFoSQkM9jugffSelb+trzEVR0BlTys7
y6TncpEJqPHhD099zzIaSmcbGubjGO3OS0YFOIVWKvWH7nTH3GRwJ6FSpVPk7OXD
6QLxvGQMK3XWFsIty/4pu2LSH3rohK567oxveRI14WD0SePCL1bNXgjKh7MaCsa7
qodfea0GNcnKvpOQrOJvEMKOzNO6Vz5AnowXxv7hnD7njkBmj6QGjP5yhvvKNACC
nyayCkF38bf6+mF+obdCbIxHnfBwIuYhnhFWnpV4DBhps3fsy+/PvLpz6sK2Uv5q
MfGIspVGovnsmgiFRvvxvT3A5mYiKxwbRlIJI2vLk4HYP3NSCl7/ai0BmiGeJNpq
wzgMuLIb0N66vfpc7D1F1VhAC8vd/A1F8H+PHfDL7YJDal61KCgCwI1sBq7HxKot
VAeOeTNsY9a3b2vxakZf3mV2rufIOZsYM/d35r/YqEvRhRvw5k8I14obyS2c2WVN
ap01AjoQDaETxlqB8/gb/aCcDJrKi60iorPxI7wnND59/L/h+NkRx/+UYJ8u/AY4
4UjsX5bqAtoxZIIj2EZtnmv5RffrOlOWEA+Fu+8FeILQ9slRv6TE9zE/X8+ogdxR
6HILN159ujsfRcMMWJnlEWZeEydU78aS6FokHJW46+XbHpZAO1ijc1B3O5vrI2CE
NYuYG/cOVejqbKC42gaO4u3AnGMtI21RvUSGDccGGp61c7/wyMRUc6LdIsAisggv
N0q5F+GjROk3LgiHpGS2pso11Is44bK/DsK6/mXVy4ZqDxiUCNlDGzamvFaqgJf9
0li/GgHEg3+ijkJKFcKRpWM6Io88UphJHE/mKO8B3UI1/+mzakZolJxqOUMZi49s
6E1ml8dtqj1NEid98tfE+vuzPpJ/x+GOVyVeSawcUzxf19BoymE5RLKV1g0w2E7b
4+bDuAaxPePKapOhi/YOhXwxBGGbvsO2rJzyazjKOOxMbKKACupg90xffA65Yb06
lCcxeUHgxLWyLTuOZGH1aGzH2qB9aBpbxS8pfWpPTuPpeD6n2UYb5XZtVep3HJhb
wLCGtXXFQrtQx+md4manqw/I2D0/PLHFmxx9qD7W2ELvTwsGF5GUbElL7W2B+f1E
1znly5iVVayoPEGmGDSFjCSK+XLPFc2bzGZ+qD7IRKAkVcBfO8SS5ozpiyt6MLw9
yKFgfO0272b/FYtyt5YDkK5YZyN+jJSsPz8vGrBJZmvDkvRFzifJ4yjCdyMUr1bH
gcvXgkdOq2DNMk69SrwqakBmtj/b5Vpn31rgQqvcS2cSjd3EUUNdJdVaPPQb5E5W
q99glJ2+ASPIXobZbB4+MciWkcTSODpyEcuVTAO2XDfl/bYmipLOIkEUpK1falmB
PbSxeRtwoBKm7QuSt7Ca+W46dMfPCij40bq/guDt40YyFD+M5TUVtntPDgEg2K83
kQGvHe9uMV7apDNyHVevAMIANdVR2Wa030rf0ABzqF7rB7PDMCy9Qgkm8pHrizCP
SGffP95jfIBYDXIgViBkdBeelHkjM3uzovNWnx/zcTOYwiZdUMfYL0flBx3/mtFS
KqI6o6A/SwuTvmV7cIpVlenxoara17xQ1lnpaAngyxatoYAj8uRSJleD/cuPdByG
GlGQKweGiQYhaHZx+D7aZnuBpOfMn6KQAdFa/PU2tnLZdPC50cYi3h1EDQrV1yrU
GpxnljoOMGyFykdL1nC9cHXcyisGUXGAmQgwQTKg6R2cyWdU0y075YfAER2vkpgM
14Nq1AApVOmzKYBrzEeeEoAEwM6qY3uQhvEsSvohgXO98iuzJLNY2nskqHbIVMYw
UapMT7GB+IM7dkqRQfynKc7U6Mt2AdthB+hQb2d/wZSIt9ksrF935ZyxZU4y/10o
qQqBeucGWx3cMPtpwZC3bRyjhh8m0llK7bpDy38BD28af/KdK0P/9oAetUcc6PoJ
BduCOXtizWeyUYVn5truMtrCXD2bz/rpBs91RJm4Nfymc63U1w0GcQZXmZJwD2qc
Qnora7Og6t5JICORMpa6DK94hjHOBhcUuWAFOOg0Ox3SZKalP6cl532wIVPGfjLb
5VAHqYHB8jYoOaGpiDKsFbZdXDRa5pQtaRxOArduWcn/PPAsfd8zt4AaJyiR65CX
ScIVv+xYGoEdj/xvIszr1xBuCIW8qJArGAu4Lt+k0yQe7efMv7PY9imVJvMsXGBz
YAHZ4FfbCmWUJGsizMhpcW/jW4NzSOcx4QIfuklS/8ROjKvLhwtunZIbYWLHcHN2
InX6SoKCOAm0tPpTb5FjUb+v1E1sDgZgyNGhIjkxOSqJihPag3C3REJzb2UAcj8x
cOmB/k0ftImfy7Ik704twMGzw+tpGc3GAgM5Ed6F9Wwjx7i0w1l6v+ZfDw5LkP4P
4e+Ut8ch5QD752ybpYb6us1kDoCdpxnAofkH3frCSeLNGayxQkQfqQdaHaQtxWhY
3Riq9TP0U3rnn8uNNYTRBLg1Cz5icJuFlvqOFte6oZSM4VenZb+vJ0C9TjscpwlR
HtTGbPy0T+KlKQ7S/P/qrobh+RvQ+65zj/oNbsRXXwEq9O49WdjBx+V9vwXQqXBh
OVdGFqSr+RXp+EvbW44H/Wf7LYYMskqzLa6TSSdd/umzgkZ6FH8b6CfvZzXyLPnI
YxJp6sw/+CjcdgQF3f9yf8bDUW5q93eoAhoNuzSfvLkcG/JHVM5mxGKHsyHlmF2r
Zgk15n3157l4PaFN5EarMzi4/SOGlCL2RBp/rrkNckgG/9HC/NDRaMUwWISl8q7c
hXu+EDUMSZ0F1HKvIa5zQGrMoO/b+JkJ6Ej6aMk1uhjLzKgluhoMfnA/fg5qYtN9
//s5C73KE33tSzaRYHheQWDjYZ8ykuySJN8TCQgumOf7WfDuVkrEFbFbTVR1v6Aw
s4HHUU1+rP6PSOuOM3Nu/I2eKAldGMg19YeI0ZLbXHecNeCcvOFVNA0DsvkcJafp
TkbSbwksNpoLVVAmdc0yUz+9V5vl9Q4ZcjoyUZ+/R1i0L7QOm+ZAtm0m3tgt3gHA
bL1BE+W4numnK9y8zTJI9PA4EoN+q0moc0Vrw5dQ0xM1lpXsdBdc513z+g9zFqbd
ISWO6tjpuAAQUskYYAXAQeMwUNWg/0ylz63bZ77+hJiOMR4ssu5eZnomqS5cgi+B
D/zksWlDTzP7BnykDaaEl6B++dtbiTt9cSCaXMtjdKaKcHRaEHz9YKMPd0l2p7gj
yf8OQOTTs6VDJ4Zi7YbwlmXQzmiJ8tRgLdlQMc11qSOo0IUXeSfRBLzeMOx0k+Vm
5v1n1uQASbHecbvVC2g8OAM1CIk3Gc/wJ4m9bnvJMi7rzTrOLQHFbJGZXcgoZksz
fvY1LyOqCUj00vc/ngeFULya6VeY4jiGlOK3JiefipE5ep9J62jMr1ZBq7mM8bG3
eP9VWg6GPtL775Fhhgq9NorHlYk1PKp3Z1XKAWnKAlBzjel7f0IKVd6H0M6s2HhU
ZM6aKfFFC9kD0o6YfdxpR+PUURS6LXRC8WA6U2U2VqE7Gb3Vq+2w7zHOi7wtqEt2
8FmnK6cfw9GW2m7tP1iv1j5yToq1nhIImIcT8OPaSbQbJ9xqoer6yz9mkYv08Dz4
WHQ65PxmdRG92NITv/vSlxeucH3UEs5hl9IUm1pd3SwXoCq7WWyCym1V9sJ9SuUm
n/YSmtft21L11+kILhyLLIMXMqE1VAb0gfwxUXAtydLNMNDRVWVHkvvbIFQa4npl
6ZTQDr2RyJ+Hx1WaeKRROn2M12PPdJBpM0RMTfstvMmP3pcGXDdRx2BUC20k8+dl
q7CTLzBvqVbdyhlYS9qIveVMW9Aq1oPl5145rUeVY7N6PUO/ZKx9fk/nIpFOfZQb
nH2gKRV2tagFTYQgQNN5a69iSODP/2X1iFEV4WH0qaGD2XrdYCNtfAz3nInJPWm/
hIiIx5hXMbHV4ymmvx9z+qgQt2VK1O5X8wzSWw8fA6BTS5oXn7iZDNzOLwwzFq7z
pJs8Mafra+JODAhsuB0lBuanh5HCZBQKoVaSOCCreZpo3DvqXK0fvYwqnPtmyPRB
T6QaU7k/C+TDbeFxUh4vYdP80tPI5A1acShBfKJ0d8YdjQ0X5h2c02RPbvfzLngi
4pI/yrE+xNbAG/v10bGH0FuoCozRnOB6hKi0SNyHjVjJB16n2ymFXj6dZnOtG46t
9dzBjpFWx16efwXTDuGTQEan+p8uEak66GkZW5SKIe1P+1PJ/Cw5x99Nx/HKPqV5
6Baz4GPLgwJ/SBAFuA4Je7/ENspz+8nBQ6uDN4Yd/GzcAElhNKPKoLzlqR743zuR
rsLiMBqOvu2hB19dMbxHhDglKZ9/2q/4BjkYncVsVkqjRvkd5fdB8djjP+T6UZ4m
2Yq1ehj2KL6MQBrGFuLoVfW6tQa5A5IWcD/JGOzN1oUa1hs1gEziBWyNC9cGpF6G
hTJWUg7gqR+MASnce8Ck2NwMAr+b1cYgvmYWB8mC41K+iR2DOfQAuOy7fkEGXCao
30Gh6Ys8g8pBAdFGy93sQQMKnSpqfMjSa7/zImRDkFAKcCnKpNgCeYUbxI/26zRh
qaNdO6g9WXaEtkC6T3L3EijsFhhHx4v6jasze8UP86WIcw+XsmaGH/u0KkJY8jSc
jRP1vDvfwKxaGr7wGnaCiyLd6IHKkXltQPdjoVaR8RZ1pTjgGJvpDDRNfayAfmHV
s4fLw1O/EvthGYMjRf9gKvioi9oDiE4kxYYQWO0eUUigjI1YPB8PjSobA5Bodzsp
8vu4244dwtkZk5Z89Vc9t0ElGO4dyRiSWnG77ggAWEpFrixfuBZM3FLyFVDKV4qa
zWy/iBk5pPr+0i0ypKRb8Ka56UoKw+Xv6m0xDXkeXd9t9fCtNwSrD5S71bS5iSK1
BPRWWwRjxTfxJHA08acGxRHglT7NKsT6aoXKrvd/wIlRgebnFSVeqxNfAUJx26Zb
vK9rgx7hLy6W3/r7vknHIC7hUxxJMruH3x0d/RXTHtgnnxv4hq2TAgWJybWfrhmb
HicsGtbXgMVYU1IB646ml2h/pSBx6hqms0PBxU2/n6MYdV0h7TB/2t+3wJODA/sS
so7RtO1rGNx795U1OeQgHg6yB6hx0PHp0dL1EvtFsxSAiChv8MnOW71q2wgFsUDs
NKpNd12IEWy0k/9av+OXLnAgadTUZ7BqtxnqK0vP/B1kid1IVVlONkkixY1bqDTT
MfXFTpZGpyBC4icfQh9mzORpfO3zUzCDlRYgbcM1x42hEmj3mkYtVKFIEBMFcCq0
HtL4bUay6w+hFyb7k/DLtsAIsLL2co+d2kF6BxjJFeouYPKM4tpklkjZoFewL3x1
r6L3adAFwXpOJSMRO8pginohlpftqn+mNNE8izGvQKXr/w1aMZZJcnrTdPAftsd5
ihmayw/Awac420wz6+60R106gwtfyqrR2uGs7P18txv3KwIq6E/A0t6WUi45P5Z1
ywem5YKuPkNiLYNakJgwewDWTjIJLrBsZpqVz+hmS13hNxIdl5xxKl5cj8hZsq84
m4RCyKufxSLADpF8JfH1vHHDoLBQfaGgvDvzLxugnq6xpRZJZmHl8JDvg/uFDSKV
QLNEhSs1iZK43GPdtixG/2DAw4NEZjXUYxkute92ZHVZHFm+/tNL2/UnPoDW2a8x
UZ8OOTjFpiKRIU/E3TH/+WMfr0PRdcrBLUDQgxRTyqXIc1BMO5W3t7pU9XSb41o2
5Kr3JWypCM0LB3TKoih/88B5rh5e0spWjgp9e9sOcHQf3IURxqin2XJKMBQAaUjU
/cr2hlSxfvy//oueO9nJjGj9k3w4rS9BqSFYLW/HVBiYVZziM1omiPMHg6MPWCBH
WSm2/2op9lKHUjpq5ku9SWBExZkQeE8vvZa/FV/ngSpMIScfhoZiJjbSSpNpVGcD
lVuM41UK7y+5TOg0JzoiTLb+HxRC5v0IZ8nKwQcEkRHruGyR8UrTfTOM8SyG6x42
ogVrBmvuIu4euOD5FfgVLxiwEciiLMFmVsWBSCM8y0ZS1gXKLTxs6euYqdw2kWm9
hphONqtiW4OHpb6AWw4hRcgfFiRVT1zwyDuWaZnYan3AljpOzChcOTQd8MkAgPCu
WLGfQzeLAcRBwgug1DG+3BB9Ldhj2jOZ0FHcTFpwWMxQS5ZilxrBkBPQOotKRF64
pUVUppzhly6dUmRC2zDRqAFMPE6CymOwUYXqIjhVJBXCA63NDN9sU0FsvcBYQfXm
Hxv+JlUBDImLm51A6NPP9G1Yn3wUlwdO8MzdSpOJaX0z90VAFghhoPCUYl6aP+4Y
wbM/gJDJ2sJxGUOxvyBaIVb6w/fkDaXBlbhTVFq4sTgQtOApufQnvmDLhj8/AcGC
rR4vXOFdoKx+qlm+VWMR3LrFLVkaIM8BGp3XwcnlQt/xeMmhxGP1N3ClfKYAzs+f
HfQ18CXID13unzpiJtNOWS5SNFSZNpeLvjxOLivTwhgvsM5m3M5lbRUnpOjpy5wv
B52sMmCRyklC7DbQy+avwpC9xPZH+MNeORXDDUo04H3ezTgj8nMDY2bY7X0l1vG/
FnlGC+mm9swF3gSRwFUuskKk46bs61cA0OPUQTs+3UoFpeKRgevjtQIj6krLAxoC
VfCdw9kMyxeybLmd+aKpD7LJHVX4F6g1iV3/ZaAPt2XaM9hlh1Xgt3C54AIFit5k
WODvankB+NyhFbRB9WuBV1jCOALeiuHjRgngepu7D9m/zJ430uIfJx7UogYVsXrm
kJJd9KCDRckmnZHelon6CyD+dBBkrgFtR6kCUUPhG/eU1FNR2EY6FEi0EJO+krwm
/yHQBKZMTgiN2CO+81aIyCMCyYfT9z26F8QA/L/6DGQCE/5Kvq7YchPxvbmIZLjf
ZGD1KbeIATaKN4B7Dnnf+dEwvlvtM95ozaQx1ZQK1qq3TV9IV9Vg+v1Rc/Nbfgdn
6sTY2FPlF+nqruWDmml6B2TomcpG7x9C1qmuRIS9bAOM5KC8CjZy87MwawAvvqye
jouj4s+D6Wgy4H02WlFaNGlBGaz56VkDXLmst83fNIa0sJoRRW0XGqSvNeTBSJ3X
ibvpipoT5IfaCkvpqFq1GNMR/3rtPD+46kpwCngmGE3M3ilFoqwljAFKVzhqCMMP
lR/d7ewuTi/RIfBja4nBE7lEzij27QMmo/+IwvuQ/3YXqbfxsTajDGaiCiZCy5Qi
RBjdi8FbLL8sIf03NrC8e2e4jOY6DVI3iJVVvBO7fBtKf/QD5BhLw+B8M2HAWGIn
lOOlfug6SsBEK9HflbOYfINHb6d4PvbhH680+cqYI3RhUGaSHxA7AIruaZa4Firl
Va/YBuhM+0681+MVuHVHwXpppHAQxMocZFyteaeyVil00Hn3ueeJLmmJocLMJWsU
mT/iXqHfy4ztoHfVCK/8wLHOgnOfExEa83COsSJ7OVRuZ3xQgGfuqp+a19d58L7c
K0+weC80RkWt1MLewlUfnDk0JWs/OT5g/2/0WUPbsqxg7SIjARZQbbm6yQr7oCzF
G5Gt/fDDgsdBftu7NWG/v9Osek695ifLvpWNRWqgVwKrgHu/q1MOFRpIvnYzMxVv
IoWHufP8MJeaV7Bc5aOH5m34jVy+7ye+cEZk31AevpHmUtB9RFbGKQa7tV429rrN
tw+ZhJeIE/hzFHdDAVe+9OLwIAxOMNYSxGVZB6Jd//m8epeSsufPDen8fV5KuaZl
ICSl9eX7r27GJRFbm/duybUg/hHZJhn9SB4gt34GVKj2skpvtAOba2k1DSMIYzSJ
8Rc6rtNPFolNkCRWn5GqiOhrD97aNKGeA1EbSgeJOFDhCFUUzT3X3qjyOX9yuOYF
QzTPnOfY64hv01+2YHZwEqnGGjcoQZmuHxTjAxeuWMTOZR68Sm6mBN9h+tzcRgfm
sLJmSSpAv9hgAnC9w2uzib4+ZT7HciUethx9MnZFio9woWbqRmfowrZj6uTalf+C
ncPTy5BcBwY1tiJXizvtWxUVesqTNCNkmmfHns5CYD5t/8d5E01GHBAn32RRUFss
PDn9kG6Hg0T06pxPpL64VL8J2RHHxyIjlfxEbz9GXr3RPcBhdF6MY0rwNBqB6sMO
bwwlvp194bSq+8nvWiAwYmLFz7Xjx1wjbScKHKMbJVqBXndE7yB/wcHLTASwfhBn
GCRqgXX+E8kOECdBjOXGeeD2ri5Sffayp2CUQgLD/TfNQCB6g6dtvcID0A2EgRor
d5h/fuFta1zbND+SlwmOu+oPJqD6TTB9/ffyVSnRPjvBMajLkwOPY+LQK0w+kpRX
lpicYX53eYlDcN0JVIIyALVcmPhUytcdxAC2pt4Yx1RipTT+7aquCw8d0ByKMQtx
rkIgUIiLKdts5qIxOYOv60dFeRlWWIkls8DW+XHdaKSXfD9KpOU5OxrTs5KDoqI0
sFya1/5y6L2ooXuZS+DqRfv1N2cXVnAC9f+pOsqTEXY9jY/9mYH0TrntM8vd9Ea+
bMEZV07s+EHqFx2CzCqD4TiXJDd5fb8Ur0nuqqkeNOXlFihqcirWU/cLURPjibL1
SnGmNMmx9MZgkYRIbc7fgm508vKEwyhT8gEnIKJ1T9wsj/i18CrUCpzc6VIe6f9y
zWXre4Se00MLNq3eDYCkoCZRnzJQ053TO3Ail2gVXMvAGKNr88lVujhWJ+XmxZZw
ylskfxsUa/q6Emd9U/b1Wjj2kNzJvy6U7E96kD8MK18VGjjTYEyPc84sVAHwmyfL
7WF/a/KeHiWAIlTJdiqFvnh+zonM+RLgwJ2lHYzba0XLzigLPv4t0lmz/AAuuRY8
QnXfC+7pqB5ApuZqqm70uX/LNcFdfOenvYcHcNeXVVAkCn4NKs5qARH8CSGWHDU5
wCKtCYBm0ZKH/0p35Gts045E+t8aAh53DPmBM50B6N4+IolvfnWOqf6Sz0xmxgw9
4LzKNjDDjoDqtykDr2EqoSuXGb8ZsICTizXevUTZiXznbKm/vqFIc+ttr2Lpp5qx
So8F95WA420SLJweJMLhoQ2JOVSZ7l8eRAi+FNvruONYG0HUffcMWz+qmClIU2LN
TBqV8wkRea+tFPX/nqAyVkm8AkzDM3RHEAjZ3uymvSII17G8WV0e6KNzrdglHBfY
kYPx5yAct2y8P0dVBDoQzefMqraKjVY8lp2pQ520sewC8KaalBgnx7r42vcNJmLJ
qtP3SfYBSFszfQLp2ki1TD2xFt2Kap7/tVulvg9vqjJqi03dMxkfIrH9oxySGM+3
6GAdAgp+swqxyCcWrr3i0UcYGVdvSaaQf0BM2hTuie0ehOhesD5EQqsknCxwV8MS
aMz5UJNa3yChnihWyobqV8V73SnlOH5YlIZXNy6MPudX8SPTMi4mbiKpEBNMal3k
zK3ncgSbf/tWL4KXjgRf2a5j/lsmS98GFXgVE9J3tiRDBbt0IpIL4qM+uN/GnV73
Z3N7BC2IhNi+T32IToRHUPXt/z3ACpE6oci1DVzOyLH0graTAwqG0fEkPz1VEJX5
LNlJTJwiOkzXHzIxAAQtRBvu9NwV6VIEPP6LfVljTqGjA7SdE/J4sPtITeL0oNmq
+ypln93Fx6Q4BpYtHddjKYsXDTew07Z1/jP4MMF5mdcVBCqgVUpRm1LqWLGbrCj6
FvHbdTK9okm9515/qIDzE1h4tf5KMgFfUZA6CSmQE5jO3krTpZEHDSx0kkwY48oh
jXzjj1oIhsmbajIY5BstMUYbmtKAQTpiD72YdCupiDKkAGM4ecPfrw62HY8LIMOT
s1oiBXExnj/DJGTPCKJfeNlQsD/guh1ZmZB189T6Bq/+fgWIeWK5End4xt3Lc2MR
vJ1JtGUzeiRWV1YtzxK2Ff96ZSEAqY1brTFXlcWk4KdUEdzF3iE+VYcqp3IIkukf
iqfDzB57C6PZeYncdy4JLQQXAS5nqS7W3Xfll+fEfDVANic/DDjGwtJwl7tnTTgp
YETbUtG1UpYsR1sSLi1RRn/N07ftHZJMchx3wqsYK0FrOTrYMBikt1K3Os62HGf6
VS9wfOCb7sxYBn9pveo3GGkuXDghVcwr5lo1kJeESiU/J5TMHrvKQchI/tRbpeJh
w2uCl7wTb0qt73QoHaVSmeIoMQwxUGmMmq2JMJ+urQn74JKunQq/GIdi5a+zKT60
N2jWByAobuDdfgWLbmFQHMzWWdT7xST9WLffjLbZcMuCEH8fVLE5GDdI5Iz8b0hy
lv2o13Od4Geu8NMs+71xgVDnTCoCnhhDnwK4ifLRvCNKn2p3azIjUaDEVwfyc+av
vtMukZrZ7SxhGBwgZxvmH3a3YiHMumHWtBGHn2be/9B7h+uIbf78xL2Qqzdfl6iI
wVeg0dulHixmbrmkFAF52GVblEApX2elgKtE6ocovDOrQXafIu+aJ+JevJSlttKQ
DdKG0SpDB+ycc3GP9CbE1RhzNmTpINxZWx6XAovFKn5jiS0TXMoCiv/90CQIiLn4
Nzm4itimXBZ9wtgjkndiIpm7dh3xqNcsqEBqScYVxg35eX3ERJWa76rUl2Q8C2Z2
cqXoAfuQMDY9XXfstPK1Gm89ajJkBYo2WaLdrDz4sfre3al+OfSYq/aOqi+p6yjC
29a1S+cjzCHJkYGHKIfnzK9hI2QXTLOtpmiwAmuPwhOdfXc0j0EmhRNF4kwTzGiR
TLVRQ7UsrOBMX1EHRa+Q13OTxeHEc3UwVNffatxL8d8PzNgPztZXPAACZasPjMVU
DgVkv91DRk536P+DUAEuWzEr7MZndRs5VNH/e1GDUZQ2vwWHoa6Tj5uNT1HfKEUb
d9G0P8SEp4uDerKJIoFzDT6sEPt/nAzwh4qRznffVzy7JXJdSoydKI+J2VHvyplL
qlkPRoVDxo6M0hMY9Nm9APv6wOF2Ad8b/jxGkttw+Cc3/KZuXUgFnPyoPuTKHonn
snBX11OUVG1aMk3BPCEm1Kp/gN3mkDrd/xfhTNNvKai5gf6BgGBMj9wnDS4g8n6m
jmRo590RtaDmVQs1/HaGDvWgpfjv85U44VGqLUPQNfhVp+BxsgYIlHaEmU5Q2ABi
wu5LvFaHJVZGXZjQikUjwIOdat2b6Kx4Kqb8PtWKYjxcg05/VgfUXFKb6WSTj+tg
kpMAg+QnCX0fevtDvCddVdSiot+MPq/NnBjExlBHgv0MYcjEwgYDo5dWIDB2d69e
GtnvH/MreQKf/1+nq+BUKU34k/FwWah2vjaQM9HDylYEme5LWYwOgQnU37P4BGIA
WmOohtrkql9TJRDP3NkAoOPMekwQg3jDSx5a9jvLucm4q/VE2LQrdOTAZwKIC3kv
S5EBml07I3zOxzPDbHRry6cEXqKY7FiQMjnkqSKCtiP54/pZ8WEPBB9S+ZQ8Hs11
AzKJKqoqmqV9KsvCnD6dAkZdYH/8pV0EEV0D0wted32Ui5TguSPOGc8vrX557i2J
8FcQcwiuLoO6vyPYjw3m3NeOsBAsoN1PAUDQkO9umce302SKHki9eglCwEOttQQH
USqrf2bNmzjJZkpvp79qd/pykdqZOCCVCpnYthrNQnzrt0sZNnlQOpowfgxhtw4d
lZGscJ8E36e9DlE8wu8/90XkIkOp1ROvBd9r4Y8v4714vZF5LunjRZ4MUaS+rXRI
Qp17qwxVyAKKOu6jtA3XO3Wjbhvu/wGW8VMIOUtQ8sUUscll07K2oxAsFadW69HG
Y903d/vZ4AxVtnsEPGMz5eLVsrBd4+Zxkw69RcL23LCdWYlwzvVelOSaX00gEWIb
OSA9/60GJR6lf6ZUwfL4LQrUBIb8yfWBIO1cGrpmcq4y2m+g1UrT8k5LgMRxRVJ1
jZIuQ3rnRbNj3MV+r0HxRctTB62YS5ozNjMSzGjuXI6lH18k/mDyfPUTRjmmwjwR
HF4MZQyaGsJouscA0+KHnyw4fMBaId8caCBCKQu6JDWLsvlRSgIq/UfFLl1nCQV0
piCZF6d8Ce59nsHBrDs25ObI6jXKtPkPJ3fwcc8VcbnnzuCsHlAY6ppJTyovhmiA
Qm6IwPdJ3pS0ZMhQBOVuYfR0UZ0/0hfOrzGlTOKeyylfDeXSjuMi0U3gE/24hoMF
0Ua19iq8VmX/JbuXTYFp0vLe6JH36BdTTYvNFBbMymryKM1j0hIyAa+ciuSb689t
2O5zyqv1qNtA0TX3vqIBKOMs8TxKwW6GfpNO9Ds/g3+hH4p320RQFO22R6iQfqVr
Xq0lJuzJU+OxutL/uJ9w2zsB6OUKt5jLpjZwm1k3X82pGb04WyhYERKWV2UMJo0J
bG/+AdzMcXKt7PJb/vcAQIldj6g0Y55OQncZUrYk+YDPis0Lm7iyV/HKBY7Lngzw
vthJ6O9iD3r/Bot/DVXmWuZHhjXb00fuYMNkXAHdk/lbhvNPsxy/MH+Z6Ge+P7S7
7XQBZCcq5N0VzkZ6sEzOuzF/t6cwaH7vIuJ+aMrqQWpoWCf/FqYkncne+GM5vSbE
yKncOV9FExDNIx7OHnTdCe+bfuwEEtk9uzGO4bqEq246uVQL1wtZplcO1fRp3ZKt
KxL/3RnN/rf5aHsB59ZR1YXE7a0+4KC5by9Ja2AoSE0v9yfDCtGiQooV3gVC7zH8
J2LcLr4c8vWPt9L1aAJLkILEZlxb/rk1rQQFNYZn5NDlbEfrz5KbzmD1jkzoIZar
az7OGmgHDwM0GPaoXOo0D3t7wTWTsjg5SLxLGEgFEmYQxNoNp4xSoynKdb5oLXgI
RBJJNplaFWMZVtGFLucD8l5VhPQIEe7EH5RmfBkLN2ekm2u74nGKuYK3jQU8Sthn
xY+ow3MSoX2TaWWEbJQYOc6l+n0R3YUVcPUyfwxQbAvMgCyeeLN7NZfNmmjRsUyv
vIZqf3r9NN/doo+8OfjA/+nOxTOSeMZ7/SXklXxSax//ApKG0zC/sSIVQEb/lvWC
C/Hwurwm8i4zD858GjL8Kzz+15DhiW7AHx1hqOkWovaH0KSfGqIRtXpG42brvEpC
3U49ABxBSch8TJrH8fZokgJb1/0IFtJgidmJByJpD9bwRomP7dFT7B7GEKufpLsO
PlraNbVwiCH/Ju/GUTsmjksd82TPJvpCjslovmf+8TMhWKWHVr6DZ/q7c4QKKsD7
kEd/vP+7HMRLwB9mgghAJwaOdemmeO9B2ipsoJdgKNPlqJODd2QIpc+dM61tVXDI
l3Ew68svw1QKbwucl3qjczPApRdF8nVzF8pIxkAB4vOA03NMkgpwnedODrSyBR6s
fUzR/ohJVG+M8MgY/0aBu45eJKQdX1/n6c+nrN/wU6Hotlk06Y9N8k5Y+vOghNAY
swWsWQIXDQ1iDEhyGv4OoHdOG8175TPUFCCiVlBYItVlAU7yhj0PYBfWYSkebm78
bt+XQplH399BzhpsNqoQ0JHwPW8/+aV3dCqGhxZ1S/DA7uLo+TjhQwwAME4R2sp5
aqnAIxH1PjbJKCRlYXhYIyfzn15Cv0irWEXHOUdudC8RK+bb5uOY9uHbIWncWjtg
99QdDEI7XbQ+0aXLLdUKvgHtpBad7VSk5pRW7+0Fq5VMKMg6sflcAwcygY7HzxPA
uNnRfYxNS/ZjIJ2QuriqtS8KPHnNzhEbxuGXnAILjfHvz7Ujow2HRtplbH+nRM1j
PDAo+pQZKVhScyXAB480siVlkQumm+MQNNndhCDsPBZh44hfpBFqESjfdWuJNo5a
yRAR67HtXoBaJ7dcAHp/7vYCVMCY5QJC76irRsiouFAquj46XkNKqJJy0MNrTTgH
9BmqcAW0xNnjYoqgdDMpjFJYpj+XnLuOa2ZAD5O8sTvB+P6/9C1UMw6ozNVS3sNd
bNXa4gFFaNrjBDjhvjXDhl91GQdvx48GnWETXpFmhAvqVqvu2UpIMdoHj/NNoGSJ
WFyhVMjvHDNsSXqLBv8UdnAPqekpMLlSW1FNtautsTZhcUv6z8yUOI20wSja8Q9v
RZidfmqW5VhIoRxctDNHAJY+cwIariFkV086q5r1WLaBGmlD0HkJaC0Vw1nlaAmS
zx6d9oKL6r8s9j1/w4ghex1mj15Y82LeOvpjoWJUjfNvbH40tbO/LHA6tXKpMR/r
2lbphDnX1JMDK2ZLhBB3hM7HCWPr76s9hnDHj5Ar0ALqhlKVCZCOWzuA8P+4eUPV
PQgkB0O+K8xjPAGpLRKrGR3d1DBwr2ePmn+UiuV4YMVd5LZ3Cy5fFASclvTluGCa
rlOgAFhiHkEgFCoC3VcMNB2RZyYpfGEew/xbJfKlityZhYN6hnffyXS/KWyFXT5n
9EYhvnCBdyB7XoU3Hmt+3356/FevMm7CjIPSoxoois/KRBjr6YJKK26J0z55sLXu
wTRSvPISj6Nn6PgjdXrpCCrWAep+qQ9UjVjASapNGe6+RkyA5oOcx7fty6ub+gm2
qZq264wMRbvUmGlTf9zwIcj6ydy4K+kE56TqH7jr5lR+LvJjDq+63Nw3/jMUx1pB
jRRfuJDSFXebZTq0ykxxP/mpRliksvlxRffZXMuy3NHCGiVTbzXPItOkucniY7Iq
n2G7Ayiemb5vv4E+v8brPJMwiJ/iKVsi7WUBfpIeZ5RmV6buvbZI2u9bYUthTA/h
WqM9KnOVg/AOwaKgM1uYUeYQQdMIkQJ8whbWEQwQgbKcY4ulrUQ6o98qP5c7kXNg
H7f++sINrhdJHmJDnbkZjjWGYfulplTqmtD5y4WhBdgRtxl98FZZaDRrMxcaf2e6
m/z6M7bwJJ5kRfjUGILH7eyAm4/NLxIcD6r7M2FhvCE++xoLXAdggSFt5RGlkYBD
irodWKG0RSzcj7IQt0zzdh6NC/G6RuNpy7Sv2jp1x+Ytc1pSlLntnowZntpPKAS0
oJcttVpP4ByjwD6YjuiCOrR9hH3CU2IPojKMkyC4P/LNNxkoF8DLvJaFQkY1vyS5
vkayRxo/XQGcTB6qGK96vuguY6/lVQroMLvluK1zqvf4N+eZ7KuSCX7iNbHghMSP
7jbKyLrijXvatwCttdcsOMwPJpr1WpWTAruUSLqe4+uAWMDXeh0hEgYhEwa4s/o4
StkgFbrMggLyzK2vGPMZ37JonALIZRmWlm+KAfVhqf5N/Rp4wffRZxIbg8D4uBCz
APddaa9rjU5nROyVkAxJd6FaEstk4PB5FnjQbnzvvGKrIV2sslZk7U/wzH3nbXgT
hZ1ZyYlkdzpIRjJF8NTY/gPFPoD+NORxAhMorSpWFZ8H4gaDkeSVxpNmCD7Gqboj
11yXBvUUP+tVTNsN3nkCu3X3Ikife5+/18RjGT7hWdt9D37XgHV+u3CGgSA+P3NL
4088DULhQfZj19pj4FKiKmTnjv1KonUOrt1IHZM7OmiX3/D1F/AnXD8Nu2ksfJIW
W2Z7iau61we3q9yZAZEmS3N//xlcII+6ZfHFruQ+4nFW1etniG0sRkC4Fn48m0t7
2vIKFWQjF2I9Lgg5Z5R6QtRVzp3YnWoV3kaOfE82k+NdLUHQX7B9QDY0BOf+aHRn
KK6m3NLPZHwG74yBBDLS8eAkbrUkWi+XDnkbzkJe1fqnCGV1xiDoWl9VA+gRVjFo
DReiH255HQBAqYmcV/RugRkTb6ftFoRJATuLr+EUFY7nX5LY5o1eiKefBdjvskD/
lJURdTJEu0nWvYkcb7iBdnBFiA+1HW9ZtLLi85YAWSZH0JYdkRBUvHNxYK5NhfuC
7YbQ2UbkRiAIv6+yWVk64qqtVnt3fPhr9I6N4BnxeehZnhJkAxVabB3kWYuneH9H
K23V3zM+g8gtfoc2SrBAmtcJDED/Xc6EmDrdW5UNJYooCwJjWPlktTq0MWDHlYke
flCSD0QzIxbYpAwwI6JKr+mSK8s9UMIrfX2nMUG1igkUT8MX4ZK3Fk/ouekxO92N
6W24kaWlyLSUNQRjvnD4qEUakV+cvmaRlAzHFUbC27H4VJV0pEHOOYJpHVtQy700
K4aV7/BYW/lD/vPgH9J3NMPAJ9eRMmSwFOtaydmJgZ3gzslQL2iD1SphvvsLdnJ7
f5lIlSXYhsKbPzFp34d5HyYmcVmXe14edc6PLrtM47bVgalMMIsCrOBvYlShtw5p
IAdLneahBTd4tZ/UnRlYYs81nUOOA9aksqm0iBnhaaEfzfbGSxNazp6QE+fGPJiU
fiDYoqGVu8BW1bC6mmEP2AIIjM7fcP73Q9/SHUY6dMpc90LDw/+qjyAW/tjupLzQ
kKARQknVzmYtJyeJh4ONLururhJN7TcJUDKFFFlAiPC632rJH3YmPw97ndDgcic9
vYSNK5cDE0+c7HRxbRJBvoc3P6ORnr5Cmoz5SZAx2sNwFtqhVqqpG3iCE1BMkxc9
42fuH04mKF9/gLa8FdA7aLFRmn7bKlSg5Tj8YC0hO9hPC+nxGx+oPslq/06M6ElX
AqEG60YAqnsNvSaQwZH7i2gSgnZ2rKFzoXpYnTK9Nd23Fbm3KFQS0akPgFkpUC42
RveJ4Ibl054TibmkV5yKp1rXwEHFIKg6cJqKlpbfeerRo7L0QPev+gkYD5/TnxQ9
NHgfS43z7MUAaJom7aq/c64L+aDqIW259tUga2Zm/rT21xleDYaIFMVoi8BF+mo5
8JrYfXCjwj8qBoZmfx5YNSpu2rb7S6no+GMQiwqpgB19etb7pvzZ8HLV7KLw6lk0
DDtDL2R1v/oQJI2n+tom5+otoU1IuExzbOxesnZ17Rr+Tyg4MDpnIo4XOrbUhJcP
Cnt90OFtQNfdWi+yVndEvU7mLwoIqL795lfW+OXaHkygLWERcC95S2PgTAam6maQ
WJuxkD6cdkhVTzLvDXnVzZwXGYOJstT9usQuUzM4LRT5BbTaj4tq7dZwFHMSL3ck
j55lDK0PaLj/pXLg0Te531vbUq7AYZOo+uxcaU36yCFnf1sOz5OM7UcOprHfRDZH
HekjMeB69/MPdOllCrQmtF3GZs+9pbjwKpoH0rBENrSVGmzSCSRjv6ceDZcWwBb3
Y0qDFlwuCGPNsNBvHnkqDxRp9Rju4Aev2ZhTmPjWgaE5rkvNOeFeSQSPPzH4ktN6
IEMU5h2lpcTUV3GL3RRGi+gmR0WHMd2KGONak/EE/jG+SULBp0eHwMO0LVYawVPg
u+aWzIHUd5H4cAul7M4gmej7zGyrXkXwxqoEfYNmZiPqZJNpncibp12+va6nTLb0
Bdl5gKAMtHIBrKyBeTVQLGv0Pr44ZhE8Ko19M4y7h6cv4V16RFnrZn1CGpMEhiCO
hMgjtKpNtCv7ySrMgBjh/je68G2v+RtEKNv7UwYsJOVdD3mtFr/PVp3SFZiGV9F7
R2V8KqarYa3DkTQQtepzgzOxwauyV6dbkS2oFmG7VIsNKe071GewquGj1KTJ2/LL
8BMj3ofp41S4kvrcfLa3FcVUSxNGazX6BaRy3wMXXvLEXuaXZ0tF68mRRoEfS92e
1ow1EahBZWmgucRcdV7o0OqLmNjYr1lIIgRLikuvVv1doXLzP/sMR2OqmTJdhlCJ
dI4Fvw0LVsfItJqhGyQm9zWVDwrYeaWt8P5U1e5O1gxqfAv7ctDXPXw6fT+iVipA
NZ1pc5qH2FjH7cknJBSCxj9QKgVIDiLZH/jcLtnGZCIMpt5rB8+qye9KqCoFyvKK
IsjhobjsE+yD5s1Kj/hYKbiPsCA4tagEKTcK11adS1r2KgnRASustAPY5uvGwzWT
Kvs2IQ6EocALS7MShOK0l4/OdQ0tYZ/qQsnj+3PR0Uc+sTeSo1VojAo/iM6Joua/
VwoUrS3NEAV8v0UR/zdE8wt5PlC1xm1iZmOoAXJYv91Gz1DmRQ6AGgpIFz7lvRko
1E3jMGRt3WB3+sYbL/Byd8QJUAQpNtOg/f0QJuzOdj65I1CVHv7BMqMwiiv6Gxyx
fu2fpWuzZqFRTx2f6CO8/NkvnC6H87NtOJks8IEUC83Ud81gSejtMzr1SXEqSNTt
WJAaS6FlRlnYoqavH2U1lpg4MPDqLNZuZ8VrJXnDw5+VfoaZvRwrBq7L+vyNXEUY
Tiz7I24BgLLG9N5ww1qqn7AI5BTT2BOqeIgJH2s5ynuWMucPSHLU18hNQDDucwJ8
wR8dvCUeYxGHgBch8FW/xm2hCCDogFxb6wx4POoz/EJA66xqT+v72QK8Uo4eKoVa
P3OPRVvcHq5MHZx/j19RC+l4NmXX0GPErVKm4f7MYf+gFj7IUCtKflkNncOEm33v
2YnpRYlZssQQrDS07CWrhPbp3OFUHansK/WUAqjCmwVTYH6yKEeAgQIVA2psXx3T
5il8lRYyUibmg+zHsK9Rml/Y20QdN9T72saLyUOF968KoJ7hNXGCh8dZOLWPq1IN
mNwq03+hQHCnYP9/I55mzzXWrgfyNQM9Sv5BtKYx7G0FPinO2uXK+XLkQ7O1WsDZ
sxH9OgCTPnhnGeb0Y6sqTecZKfYyBIZ+tlNmEKZwHi4prFD9clo2LVfAfb50Aksj
tBIlznQ3stXIvJXMa8P7lVFsmBcwRwDvlAdhJC7Buuy1rG4a3APyGCsmlfr+Dr0m
s+TVMD5vyMQKR4ubuTXeb9xf9PXFF+a755rur2hc8vqdh1HCtilRMQPpe77moTDQ
OBN7nXbb+3vIPG9XfvWtvXgwDlLKeoxd175Fo4vFRqK5D5LoII2yibVb8op0t1A1
PN1t0rkf++V0FJMe8Ud565VvRwA3XSIw2LfDB7tYIiQs9fDqWH30hOC6rshckprR
4xTiIMFM+fIMhTEa3pg/4Ydn27tk6Z9dAN1ZZaK0dlVk5teR0u8rbzsORoPguZl5
xmfwIQeVl9u86s9hT8/BrTwFzc46PRm0LRvwa5JgIGtsRkY6imxMRrHFgYuhf4ep
uXzvPJkuLkOmveza5szObTmtN/FiZ5zmT0JnLatZ9s/nLbOOwdSLwvsNJc2Dutw3
7JnZ1t1xxNZKv43ZCNXxA2pQ7NM3zLddsAFpFt7fTBAPCAwh1thY4z+3LJlmZGJh
f/JqJrhZ2KMx1edqWHcMcnjAtVXmOs0pnYIgHWXIfCADhSxzs9ePQOuZ7khQB8Oi
jNssRcFn9xuRiqKGbKZfpbcQ55ol0ziS4MhUsn3VE70qaN7+u6YOGa0EG+U8Hkbe
/BneWJjJeLLzOWSDv6Lo7kD295ZqtxmMNnI47snIruUPcVfLOY/j7HimEncKmLhn
ORlyK8EUVLL2+qtdku5nkcrif0Aa2nLX9N2fkBq3TvdaRx5qpeoBgAf44tvEBdGi
05I8sqFRCdpE43QGgBiBjoqnQ2330rdkbZ040dLFHhUPiuFkY51icd/smsBV5RR2
oseoB2AGUxyVeovQhZ+mf5ifF1EZ9WmCjnsM6Zc1xCXibxXWxO+83e7KiSVkALtd
t+S7UcUzWpyDDj20LRiwgMzguz903D2yVKYcph5Vc3f6O3bmL2e2KMEa5RnAfPIv
bae849RYVueEWzMSjb1TaqIvjkZdT1h0q8wKNTHoeJYleDen/0FW4DfN66v2yu2n
SfGXz1a9F0mhq2war3z7nhWq+Co1Ccof9m+ktEkPr46fCL5xbRsZ4hXRdKkwfetf
3mMnGCWa0Mztxi4CdPRwM/96XkGi+easoYDdUr3AtMIY0zkU0fJKMih2tzopPOgF
OPRB/Y7Yc/88s2lM1eRrp3uxu1CGIcqykZHhwOknSjgNmHRFI3va0jJBMsZXR75A
KL0U9eKQ3KfjOPDpZkklpyDWftwW7Jd9Cdxcu2KoOrHpZdzDVIgQRZ323KH5fruo
svNDqWeNwL9Kctvc8bMBvB7S1ki8t+u1nU6dsyaHqgAvkoZcy/16Psz6UwavhnYw
C/o8d/IiikmreCV8+rQ+e33VxWqSfXnkqu/S0qOy/DmZ0cis5N1J7ITvCxCxS0bU
qf+9xMLKsGk6EXYNUjEU2OOJy2XM++MUi3pJHl9EF7pwAPBOUKSY+WBL5o6diOXk
883pd0OcGekORLHfMo/BhQ/YneMK2X4HwtZR833OgkeOj2y9aWdJDH0sYoXdq5th
HuXLKZkLPbr6pnbDsl2FIEL5FoEjF2JbqguTDTM19USB2NIXvHRKRQEbxF1ecege
ewyeiiAchEspKhH1b4S8ZeKy5WsJUXBwlrN3aG1dGccCNxTpP51FetCkb2h5Rdr0
TcBmfUe3vkjgCrXiT1s4H186ee0DC1JDQmZcPSYeYggfN8eTaUBJGDoOY0K962vq
UZvvpTK8Ykq0DfdpOe2r0gNdJTYer/INhINUu4Ov7CjyounvbIblR6LffS3hPhR8
HGY138/nayD8+TLzjQgu/Vn5126BiPunEndsts9VycgpUWlsAV4L+sdhjOgoLhZL
J3umr75S08sLpRbzork/JXKIUSfo5yKgUFtcES2/laxFbZZ8cD/Qj2G2m2XIxf0E
keLML7F2Ej4WxRbf5aCaRQiYevgeRgZRt2bUkROiZoyXAs+Ar/5mH2nsFrirXM2d
jh7xwJwRq4h7wto5sPm40SrQnZY3X+/5wOR2KGl7oIk0EzMy5OMfMTPi8Y3+foja
8iYgkFst+cdMf8EG6tmuReX9Oc7tOYtpp2QfZG9ZgsKaYa8YWQv5cF4PszUj/ooh
Qd7OdohQbrpfbHPBU8M/+D4Zu4VH7d65kEVAU7Fl2GPTjKhURe6BS50w336v+tWl
FmMQipk0fCyAxRwEHDjG8m/vl0Fz6l6y1VrLQ8dx7LNy+gH8TVvaqxNCx0gvuLVb
ctkiaEVWao/t7ZGMqidQO3BY4YC6IIIEzZqoW3QXGXsdbJ2zrRaDV8hW7J5hFLlm
OP2C1p0qxNXJhUGxSOYqML/4CvAa43sGQLkwoH5z461QVyk3j2Utl/N/CyfRbbmf
4Ev++1/TK190L99vDblyfMNc/tBxfyiK8dxUVjZ310xU4xVcD2fHvaPa4rGXCV1p
sUSNweuPftodDqcTZIFBkpc5F8SBgI7J4URKC3NvH7FMJJXi8kcpRvmHIhGZ3H3i
q0I0fGs7vnxxLsY/jiqidhM5Jg1hHgM7Jb1Bc1krINwB5NPFxWmtagoLflSk+YUN
cKmlQx3tLdI+hq6DCJyPIIdL59fmQQ2X0ygUGYcO2H6+pVbcxp48WsD6SpMiQSyT
dUxH3Zz/ypTW9C/yh+oawp/BVVrV3SO2lAv7ccZSi6oaztVMuMQZXwSDUiX5qnBD
ij67FqAt8PmAnDAs3qoAiDmLNevnnBl1J1WKJC/uYHj3mezd2Q0OvJYiMzVwKG5i
63HTh/FH/Y9R3wfJloseql90d27Bsr7YSXWpPJ39WkHczn99uCDvC9sQd9dARzoj
CGMhFPacqgcLUkrKnBped//qQG49hXaCTJHzlaoGf2L+ODos6IRAHus161ZaiXUs
Dm0ZfjTtWYEZxjayr3B/CKWiHyngeP7ebVkgEcZVVZUSqlOFCALRzZ6PuLoYc2cU
dNygLWdl1EW6/pNoWAmJzrYFYMIIpdK1fv4Sfn3xCBWDbOW64zMg1q4FL86oIGCA
uPwmzfNhydGq6M4akINZ30rgs3IocRSH4axGP8dJEf26icUITtoEZX49WBE5mLxb
OxvQbWUhjhYSTgULnsLwAte/2mmFGhzMc1J5oXxP/SNDA7aKKA4KmR7cGUMmyxfF
H9MzxsIudOQ/wFpLP6YNq6CNGvFM2vmeLlYh4PrllOoWsmeVj8OyeBqua5G4ErVo
8ezOSb4AVTi7Svz/J0nf/C6OmCgZHpM3q7Fu2cpVJs4IYinAzSymqLvWUn4QzW3/
iIoC0Zo6bvyLeCA5QxS6MmMRFUWY6dAhEisV1mrYoK7CH6WYKweEdsPU/R4EyYUc
kxBb8ZOccFi8xN89bZcBgpJSYoWbDnwrgVUn0gFW0c0ACIpgHSPmsroCj+UYQu2B
ng+chpDEFKzHR6IkrpGpokR+iQL0Wh/BTveSJ5tOimkTQQAnO4sNNGzIDgLp0VJ9
OmBKTnnEe/SNzEGfXXsO6/BKNEAAJdjiK1+ALwlCTvkQz2I3OnFTZQ64E8l1FHZr
kmofCgD5Hj6U/tvEnUpCOMpr6QnkdugSfJyzkW4gszExPcOxWPMxivawZRk+HCmy
QkOEtVEwXQC2KaIRjQok24JYAoqr4T+4NnCyWvaA2anaU33WTmKXoCdaeqxOGMzr
e10kMgelC6PJUNefhDnj/FY7lwX6RebL62PiYNDPrci7nwAlMW+7pL/E6aJe1Odr
spES5z5Dc528K5Q9R1pX1UaWtZq5bMdhe4sMYr+jhSdn7sQNROyOA3irFpHW9Pgg
/E9dBb7kT5KjMUsrgnoWktEwqUnoq9X8fgXXIgzTFRmCMXmHBr2ROoGPvFOmS0O2
sftXsDCAD0a7q7GBvt7eOMJ5P3Q0KsrGE/AGoDpJpyFFQjQ7CH5BaskkDbRQfDvq
06jCsGba1D9acbCimVBTN6BzlksI7F/+eFMDpYMZCuPW3xlItH9BDa6lm8hqGRBl
UuiqlM5ilte25/PWueAFLTQTnY4Cg6Fv6zTNYA4HKR0jzF9jLsrsNietw4tRpKki
9qhXz/nuweA+IeHasCcnL7w11esKscZ5POkgWYcXko0ttMEt57mgu7ELY8ZZKXAh
sy2bWyWpOI1+/n9sH2DNQS8sjbPX6eZNzD73umo6cqpaj9M6w8CFUaa6AGpQMejA
IGBi1FdzhsPwLYBKnfzuFpy6bP8NNHH5jjtdRpjDa7j0hNaSAzD0OJ2kIM9f9sKL
L4aDoZQJRBuJ9TppPqoPE2GdrfOFNFiwdSKBDYag/Dm7hGQLkyMnF+AxBL1PLabm
XV31eH1fVoKSBCF6/i2EZUwyqQolE9ZL2+KMK3zp4T0QxrSyu/+2rL25oT4KbPgm
trdxl4PSqLrrZ86kTh6viXbBtCYZUFfxXsDJgUnPUVdgR3J/E+ZLKAMa94lxgtLA
HxUzotaRBANpQldHgMiD2SuDieoSi2Bi9AU4VZ2PCJCnP6pFRNZZrj941ElH++9w
D8KB8VR2S32tDpMAfWpFkMigTGc+OjmMyuaKifq1p2Pl+BUnr7QIB4ky+x4Gw8L/
MT9uNfqiyObBknBFQ6e4L0Zl+dKQ1rpw1dWfQ/lMSCRK7Fk8KcX2Lt3SM9MCaYHl
4uMtA1GDKK4H+vKkumvoU5vxiF45c+MN5ZI1tXec1zKd9Bzm532U5lk2tNaClvZo
ynCE/sVFkKxTN9c5nPSAwQE+D94Dt+8F7GJzNRCx42qbTtcQkxFS/8Hi652mqIcg
y0W7S4uE/k30B4ejRaQu75N7vR+9liPqcBsB950S7sRbdi74XoH7qq5oq3N3MiCj
+GJ3gc0CMwiLSekF030rp3b2CCHIb99CQCDOtGCuFFqzGAUovgek7G7Gsy0GwH9f
3voQz1wPNgDt6gKI+v3NVBo27ukwyx4iSlQOj5zmPObFv7aio1wlQsrjr3g6Q32Y
DhhG7Qfid7xWGMPIfd0OaE3hso778zXFE6rh6FHH3mwbcDhuxyNtpujjfuxEnxgt
9F2doJdnIcmwRqu9o/7oj0gMhHA8QgvllsasyZbZIIy7PkeUCrKydT8uh7tqXtqu
oiPVvii4xirpqLZPi54WIgYA1Gm7WORXy2A8URGeVnr6YkblKMDa16e7O0wVTSDU
lSscnEFMzkwVU8gCZPYDeWuL7uNSJhMvF3M8Fw0y8+0X1LKb/0Pl/17yxnNGnJ2J
EmXaMD0aeCcqmVUyQ6dz6gW9mYk6M7qG0YmjNcdhzV7UPHJPdZHvMlT+IIhVcub/
rUnyBL9L1M4wx0UfVbUO/ADtwNNRFDG8HQ/2gyMKSEiAJtMwZaubtPNgSTclsrwa
gT9JuTbxN+rgY9PQKS1Pf+RVnRDMwl03MlUqfCVXLZAgredxQNMjqvdJp0WbSo65
frYGs4uLkDAWoB865gETzPnNnrKjzO/5U26i04HSyUsgW/59OknzC3JmOZDVM6Sj
t2KgO4YFrZCVWRCxbz9COQ5te9uR+rVhRGnM4LOU/PKSpXMcqwEh5RH6fIS9DYXF
nrzYpVmF+WRIR1614X4hP7JhUr54TQrRGIw5j9Qasb4WsIyPuJF2t+Q+6M2twfJ3
30LszTLhjhZXhZpV6/kzotwSOfXckoJh8TdD4sxGXghhVuOJbWjpWl9Fcbxsa2qd
zlhbaTcVlLLNx1vE9dAkZO3idKrdBFOPdp+gEXZYftc86eFQLOrTIC/uljDCMt3W
Xgh8oAPqCmEGOnMHTKrLIzwxAd/fNN9m7nVJlJzFWlHArOzVnKIUP8/Xyhj6dvHR
bN8ChzL5VJ3GrM2Zm/GAwhfqyzBGT2pUZGIAshCmo0XIfo0K5uSt7K8If/4A5XpP
wrpdHv3wLKlyhlq50CsQDYPZyKQzXQkTWMj18beUN/IgYsUBxfSo6pH0CM34lG7a
EzsyqWrPgQDupu+chW0JKienW5WZeUZW778IeTET0/TAqL/D+9KDxOjGX4+8DWUv
pKm7pYMYHSOt68FzSI7dK3zEgQv0Xh1kzsFsaz4Hyu5AQiBd8okuguVHkY6e824o
pmMzUi4/xIpC1n097/+yZnFxgZ/CL3qknxlkVdv3mh8UGXrUFMWPg9tEK0nqhdNB
R51y9qMhqZUdWqdwqIYURnJEce+Mc+Gl6Y6b+7b7bYqkzjC1aT219QrxEaoz5dEl
+f2rT7m9qgyDIb7ULn3swAIVpi81AJYziaQU9VM7IkBb2H5YvE2v47Wbu43onRD9
oK3bA1CJOmvUyATr2lx+sbX3+rOaeY/cBGGjSSSGH0djkdFrxxcZ+59S3H5XTlt1
520KCrC9r9G8dKq1VY7XUz+bIciD6BO51Q9e2pL4Pd4MjzQAvvgVKXG2onOC3eep
VQkEniESoJD/ckJF+P/di/ydGzjSa5nh1g74Ux/M5BIOr0SMawqTrPAq/c9f+p9g
MMHbOCk59GsXyHkb+e1B0aPKY7ZW9dvQhbLhqFksNp38csdhezvPECv4kJZTXTxE
LoFYlxMBKGLPxks+npSI/vY3fBTqLishRvTBZmFl6kShk8SdLUFAbluii4Pc7LBi
Ofh7SmcZNW1rxEhmWzwD1z1j6j2CjkzvfrqsL2HZTOHm1n2D0XEYou5StGEnrxpJ
Bl/pKV+vSGs0N6O3E9KWiMA/gOwLZHSjE98pVkyD4QWtDPvbYSnDhCFAGvUPW30H
+THaJMIObJY6hHxkNkMh3Kxl89pBTM4V951/Czm19O8xhrJBvriUGdhPhGSspy5n
rv4VivnYqrHK3eU4DGnH4w/3qI+s9vB5XubrRsS2t/VsKZDbcEuAHaopiXW8JxAm
nHFuYnng9U/KT4n+99v9pxrzLY28lmg3l4i/HvsxppO2EHCaPkSa+hIi8J1uCrxc
UsTDKSViBNztQeYvHiderJ0lXPRkpx1UZ1AP6P3NNmuP9mq6g54JSJ3yR7ARphYh
QRcnJbV+EGot5+GBv9HcKrzFQLaCrwv/k1oFzYK1uDsdbnWYSwZFb1uLmGNQGv/Y
XO7WbO/9FP8/+nC+8uBDs1Vj1q2hhBisLJvsElEnIwAaSml9varbRZZnE/z6pOxt
p+FiuS188/FFBobgWjoleRPoRfgwldUvIVw2bnK3ZLF8vEhvEpnYtQk4Gh17ME39
+FqI1MZKvEDDk/J69ezMlXuS6L7FRc1K+QrXoMnOIfeG9DJNsKl5OnVPZX2ZbFkY
Ef9Dpfd22PF0A5J8afnpy/hZ3M622AoH9siZU+hfqdukebylkzyqfnu8wHwEWJBC
jTTWu64Kqn+TPIWSvcufP9q/8OafvdWHEoqPTQxpnTlY0UrKYQx6et/DVaqB6lVk
p1Pq+ehozjQsEucg8g8plIQckil1tzIvj3bRzHjB8Ibux6BqrEfTIU5hmo50ZVNx
dIFj7oV43j7H3gF2nrazxU5tKK/akVgrSq1MPFmBF2eRZhQbHwLuLQUqwuCmfzhb
F3SCRPldvoLFBJaRKgfUYfYo4fBOtRfpf/QWlqZw5Kgx1UeEmY91jBbWCdShN+C/
xmSu7ES9kkvGBFT5jm1zlW7QiODbOMxguLy45KyljVPF20X3AUrblk/flfYvOArg
fVhDuB8R2a7Hop0t9YkRXWev/gwKinO/xS0k9Cz89dsyFZ6uwizAlrBf8g92npsI
2x/MuVoTvqKv4ttN8hSyvVZOQsWGAfE+52KovQ2v3+GYJIJn0E7Lz2N74Qyet9uj
fejYvbuDU/da7Cjj85+yl/0JYF7KYLd76SYLqYcnpiZRiGSwFYECdwRVQy5WMC9z
1Q3qV9Qkl3oQyxWFACUgq5+IJD4rnswne2Ct5I9k/zG/k4nEUEVm/n95oxmaoiyp
MiYa2nfolc2RjBfGaA0xaxXXYvQsv98W5azMszLBkIvmqA03gFeB4ZrdvcdBy1cZ
yLpdCAzhz5GIMRSMIVTO1H969m3Z615BMZYK2Jxg+6AIBVRFuSK39ityxFyIPrJm
L3+RNHZzitAPAPGNTMhE1JXKWNj0PFUJBk7Wtixcy5zmuafcgeQF6VTivIyoNj20
ctU43nWlHEZI9B7VlpraGpW1yOzbgI/UiiB7nqKzwbDqtS9BW2ZJKIGuM3W1pWkt
C5hF6JEX97XfJiNdYMz+3lqC7xQHgo4uiaWc91eP+sAZRhK1Xnph6K3/okmLOdEZ
XtU2WM8O1Mi6Y4ka1um38zOiiCp4SYeFXkvnu7QQIgeVz8xOQYiQX9Q4p6khs+tS
9TnJbLkVpF6FLn7rMyq+GEU7hCE2BKRSQddUOS11nziEleXHQPs0cJK2m9pR5RrA
M+H4Z9frzd9lZ873ozjtVx1AqybXxxF3lZwqDOAE8ZgP0uBuTEQwlMbKlKrEEMQw
bSCw07gevD7yZEdUjPxY1OzzK8FozP4EXM6hT2XAVO9pEd5NKrrJiqOBDfdHNTY6
cHEiaoht+iKpKCPsFmdzWsUrj6Ak4uGO2d74SGY4ZBk7o92P3Q4NOJkTTj4qqWzD
CM3PhG76fEDHSI7MTAjdRztKrBC8i0ffnW8kR7QfQncVE/IGBvBDK+yEz7v3gD4L
ZsxEZvrCYsQZS9fGwm7gfncPXDMQfAyc+B/qo8CS9Fh0NNsb4+wU42hPmh83PtVi
jW1J4+Zy6PXfp53yV520aCorxGeU8qMpecmZmJ1Idq6mgxM8cNUhe8EXsgyDbFps
VWFH5eq1y7MHtwldBA+ATpX4O7zXrOS8Jml55neXvmM6MbGAaR1gLvqzOcds9YNh
d13CNfkjxO4HiC45WUijlacrV0VBHc7wV5N9u60zLCxMx/nR0ZaQbWJwklDpxHkE
0lLpmV5y9VyxSgISiL8RRFr3JkOVGIGW+63O9L47eQd6bs4GziKTwixWc1qLY7ls
LdeWictg7Twv2+68i0NIkSLgAyCQ7r8XTOK+jyN51SE3JWN+Z01UpoVFQkKiSi7j
Yoojo5h4U+YM9+dMgwd+aRzGqpMi5ayfBzAoGddNV/MYpjcukLLvdRX006hakOS/
LoXq9U3IghYiS0OP72HAKS8BaKiY/++60nR4bDy3TgPHp1jjlgEw5XDbhuW/DIqT
eQMJkET0qpyfLqL2i4SvrS1S/6Xg8r8CWSvEgP0aJpmkbRlcwmsjWCMOcQp2C3E3
qwyr67i8oqfCuKbMWM4qFyHXTWRAF0B8IxjT8u1GG3O6C4v45xGt9flt1MBx/Sa3
wmKpXHDlF1gqn/LaoQH8fyeQ0PA5+6sOdoJa3poF5B0f+095Qkj/X0p8i5L8cSSX
mQoSYpwGw7geH2TMzMKlyvA6XQeZ0M7mHy+J6pzb/A35NDV8Snd1I6flvqQzZWe2
Jv9dTl4aDDjj9MvV3vnc9EiRWT2MnUFoeHtZCjAZi84Q2t3HYGoP4Qbv8kX0RbA8
doij93eSS/XDTxm8TDabuTzv6dGVOowZrmfNjoqMQfWbspC3DXH4rOZ8l2fLiDGP
lNRTgOSrssTef8vgB/DvbUjKZj+xx8eG2YGiwz1ZOsf9CozC6m+roZYc3Mc4D7EO
ygDhbMR/FjamScr4Q8TM6xrKOIhSNx+DV8exz0TWwfTRddZyUNqZypw5fG+YTG4z
ZBaNNCL2UXdVbeRr7ry3gL+elLFt/8nyGUQeDsL4EbXxF/a600U0XiwJx4jaS+XS
kIqLuPykow1T8yZc8hg+EStQ7wOKBrxC8KpouDzmQP/LPRJOC4PcXjsh5wUeAz/M
Hx4ZM9X6mbcKu0w8NvQ7z8G9w74NRBiwZWpTqm+sgaPxAwPFC75CETiRI2gNNnK/
CK3Nxfeo8U8vq1yXkifqogLUowDDe4CJYpv1dK0X0TgKvZaDUKMrHpo5T/OGxYgW
SDoYKh17nfYePRQXVFnrC5zsHSL4mz9nD2InTqM2MrS2PpvDr/ediuwU7F+zu9La
1eNK75hVFGs8HJFYFhCW1wDRCgQTgGDq979XdWEvK7Ytm3XUqQTVPMXfqSdX3kG1
YbRaOFNLVcfrmE7Eo8Z2hyjEds/DFXm0hPgN9N4c4962Fd+ziVXqRe4JWYqpf1wb
DB/SPT3UqHmpUxJgn3H9mGvp/HeSNSVUF6vHUXgYg2Pj0nnZUdbyHw75Uo49QXgH
XqlG17sB2xtzbfZH7+g+0he46Ya/NOGno5d7GrAXi+F0N42rmqzJSE2K9Ll8sHnL
o+mZdmhRZ6JNMRObCRMRC1FYG33sTgiug8BF0mNKKxKd9I/1ywyuJTVzcF9gGK8P
v50wexrxzYZo7FqgI9XxKmsDuH5zqdk8JrdlQC7DFW14+SThrldLZQJ2Kw809YZq
InKw469hntP+MNu0eBOIO+7lu8pBHTA1PG7IXGJB7cCy19TjZZbaS7epjrpKYzmA
qQGXZHrSDhaZ8WSyls2QEZnTbpOENEOBN3/tz6SXoHeqHZJFxT/6HcF+FheRXrYX
UFJ5IzRiu2GjuUyEv9JR0fJX9PNs/rV7QTjNzK/x3vOkjp/ijVzBrCr6lYuLmQR1
M/CQraDt5Vy+A6dai9n8bYX2RI6Rnnzt88tOV+/zSDJtZEtyXA4TCmSU6hGuQuY7
LjDJUVXaMVyiYk7STCj+rIQQZueeShlkUYBFfQ2kQvp6Lfk6IR0qHgJVdeb7yjMU
7dVgihY1reFF71NTyOgYIRyXHpqGfk7F/0CGYcFLsu7yHUfdQ8XlfDDtn4pFaLWM
gtB6PkocmVmFVP/iITZz3RDJUKgO2tGokwR8wH1/xu4jul22OBmEY7GkS7wC6A+h
1KHuc8/6+kRRnqfZqfODVADYtVKjY3a3SYJtHCP2bk/qaUsJ23qPmzqHwD6i1u5v
ey5OgDZ8BN8rLzjTbEOl4ONhPNtCzgQHeouSvHmiZRlzJh1SL2ifPaQYRd3OvzCN
lfBOTpZySTr24Gw7QcnElY8VVIilyr1A1dTwQ4DdGw/4Du+N3k1iFK7Cg8oWzyC/
8sT7ofPxqU5Fg2RhCdZQV3zFS6VM89kD1ZignEJmKRWl+tAWetGA1mUSXmfXkEpU
AGGw3y56pZIdgQcQPSnknX4eUVtS/t+0Y5zl7o2lumlaGmbhzaWX72NTAj9rTzCm
48eu4sNcuH9f12ib2LbIponCvCfiT/B/3yG+XDDTlqwizKghKoQNrArr3K1IigA4
6PdGNS/j7Js1x/SkgK10yxIfXdbAIvEaI6q22k8Yh7FNT2jSkz85KN7+bUmwU11h
tm6lL7+z+4UsTbiVkHBuXMwqe+ER9S0gHOfCVfR372ukk6N69+BQ8r9+jX8fylj0
tLjAtrcXS/RdyuUCItXwfOLNxmRKGqPY3jjYOKLnFKJ78LUqLX36By52kQq7hNXX
TgOtH2XxP2saY5Zm7/rZLuzH5MYSIny4jm53oyYXEIAc3F3rjsq28Gomb5vBmtq9
r8lMVnZYyAU49zZ5qYdQ0CV3jafDDM6gOEKpxQZv1r88U0qsm50VT4oo52azsDc7
FI+TPUZtnqYeUDXKp98z/8MQIB2RVPcDDfnI1MBuGtWTOgSoWh8lGGSKhpgFlnwG
8qv5+nZ6Y02UDUKiONFPAAoTbKyj9ZuPOsLEypTVgpuOCUFwdz+RL8L3qT0vJ//E
fgJGzUiqd97ZydZYI7l9RnMByX2nloM03rW4SotTWNBBCGfp1M8cz9mfIisBRTHs
2gQ1Z5n+vUFuxdTgH6GuAapOrG458Ko9dH/kmDfl1E7NI46gSGaYnXPsegXGQN5M
bUBTdiXz/MRDq4e/TXM0K653oFOX3A1bmJ66iosISk1Plf820JFT11q9qK5L4jTD
XUgBZsp5AYndFW1kCYoCWvv1O0Ry/XkqOjWj+Dfj6hjObHWwUe7F73/D4D0vHnd4
etUkxDZahA9qx2DIcq1+qNShue616vJ5ZC2RvN3ju1Qb1+rosPUJG5inAoU9Ucgr
MRCovm6cvsDI7QHeNmdNokQs/8lhNMPfz/FMdeZsXGu9vQJ3P4XtyM+PRuOgAQ66
YQbciO/COKVMX665XoC2qvkvNxVGCpoMmj4Q61KCqn2vSp4fKmu8W1LmODfbZ566
LashdjlE04UUiOjZiJf6sWE1w9ONFon0Xxg2HR4Ks35F4voIWuYUU8f0M61LF7Ot
qYaVcRmc2oiuBHNAekeQipR7uN7jTGona4CNRF3PodOQ0x05gs9LTIUJeUXt3f4C
c4jtc2ljXD0hJqX3P0KfcPlJK8W+DPBUcFKb/uCPqBnEne35TZ1u82WsURbks6ze
EWzoaicqLYR3mm+EevVlayO1CFAxvElT1Utig8waG+dCjxlii6DoglZJD3FfPq2O
AlR+x9QpgH+bSesdaPj3XFZ91t6Y9qAKkVKQQO60kAZpaV5/E9WCUR8q95flpTv6
1dy6tojibWq6JMpRRL6YtS7YUNq4kfMR4ce7fszud5lPykfjU2HCOy2bCm6ANsMI
FTI+NLPgby9HWvmAQwM/MAdehNfvy8Pi9xBTyXEQFkFbaS3F2P8wTh6pz3CvMK7O
NjK/gCbP0LTvam4uCSNypaBK0mFORwUq6YmVM5u7ILcKFEyaINYIfg7ISMLqf9Nu
oXxS2ZEdNepM1noNrST6sRSrGSMkXvTtXz1sq51LQy+JZvGlGmZBEKCCGUPyWtxi
14uy8UpDeUYNwgkq+yRX7nEXP5IEF5cJm3mAfUPnHRfyqGq/yMQHfU7PnH3AvR2J
6bIjduF3aM/mgu6AXocvO+DLHJGRP3IoCtIOXYuY2ASigKDeRMRzcmgLCMxg4Hny
duV9BPoyVwHYPWaKMeZwZJ/4w+7WugdPSMfvd/6qWZ9L5Wza9h+SFxXinjK/i/MS
xxV8JeXG45Q+8trMyrHcVQmzkN157BZ4eXc7IHLA4RykSuIGZH1in1fBbofZoTt4
JELsCIs5zYHVxExqwUuYyha8smsLZamdkFn8+MlZJYbhLPZ2YYqk3Syv6De+NnXq
ptOb5nof55KZIHcTC0KurJepWJ0HFmUICYEsWetnBHyV054Wp8sq0d286xLDBKn5
KZRn1q+oq+H47cWZQJNsyAWvZjZEXmOpsoCtDELwMSW+mkfshzaC8n0It0jV+eWj
JGr2AF3JMnI06VtFousYxgCJC8SJmj0R74M3fSa9OUbuMEGiMFSSzpvTW5Y5mwcG
ee2IraZgDbWaxPvd7Daqm2OHr3t4BH5FPPWsWbFs9Drsh7YwcfKHMeubbQHZnZ3K
SEqpdjDnOx1CUS11rwa3MUNbCTgZGpjLH9YySyWldXDbNhpaRHDdbZpNnVkAg8wB
btKESOxqzaOstcAIliBAxQYLNtfZn3kq2d+kSmaJHS1vpvZM7NKgnlBaSxwYuhTl
oZlrjrycK38/dxfOTfWiO7q9ENgclfTT9RbtivXkp225y0Ou6BWryG27HUx7STRC
SiedYBNJ7xhucA279+ANW/p1AVWZ0IoZ84ZNoWxOCmiw1bRuVMXaCLdqDuFOTubD
nbjwcen+WhdAfOtCXunDSRcEN++w2xG1Dajvyj9la8zW/6TJdfxjpHVxhWKoYfbu
oRdvbOrkZAb6mqvxJBIm2BGZy8ixBF6to1Awj28AenZzWEuhq88EAVncSiNDlkMd
qqVC79396Ow+sDjqvEYuZdor9IKun9q8oSlk3HdwYLnYiuLr5W9LqfFqnLaDmOGp
ej6kNt6UbvCxdNFh5AxTtLFix3bxzpB+YKz7kmcMmJxGN18ROmVTDfw3BLP/BKVf
Z8Z+itVuof7JhA62iPUDmAyQLflAzMprdz24W4TBoP4lSgf+GxFuTf2H5COIlMPb
2aZjw2LoMVZDu7IBgnvqodmplftFN5I3fbpJtH/lDyEURo5ynzFYajGl5Ifh1FQf
Kfkm1nZZDurEOd1hdT7xsYBx7NS6XATN3oo9lPe513jCgMLxv3jVsmCn7yI0iB3F
m0jjjhklUoU3ZJggh456QUT3mZWAUpJ2D1GZs/ara7bPcaypMx/7BYL7k9F97Jp7
Ex2YN4iBQA08r/jxtDXFQuelUZ1IQfcEKznhJui9ERvo9gXeVgR4vOZaQo/uTngi
GdfPKu3SkqBYjN96wR6LaMFars6fVv/8f/lTwP8JX+MpvxRd7sFW47sN5WCADHcT
jFjZYEkav330dCWSllE/SHpF8/fsBZhhSb34zDQo39gQz45OipGU6EhHdkXz4SRJ
cnrl48n35KAA/vpN+zzbBIuwuLQEOkxLogGHYSbJ+b3DJuMhBAdnqEZGpNRoMUtg
4NMeSh2iS1vPEbdxwAHl+cpMHpmmpfIfUCTtIGuF9d/WJA+x57DrMc82pnpsDdAo
ry/VeAfjdiM/uK1PXU3U7tYT0HZ1priI1ZGGhdCVcpOuLo7z/f5GhdbYUAd9I56z
DrU8W7u2WSn9fOYYYrv7NeOGci9Zm3C9Av4Bvb2ddtup8HhTC4O7PUSWoMIV1eYh
+L3Y+T0ff7mY3bPYWX/lpTJNs9Jjyk+diRj1NjmWJdsJfW9xUe+aZyzwxHrAaiK+
dH5VaEziWvwSNl7atofVi0wLQlQTt/xOXIlyU2Cys+RA+tgoLf7JuGb2pnA+DvKc
Sj2I8ONNOT3wlnf2n37Lqc65ANGtFbiC28WvgbPVuct/XR4oJFbWlbKl5Xu4PJdU
0PIZ2Kui0W4SXBFNP0RR7eioOxbX14n/AATpdyoEL1Au9mTcCjk5gCvUSwTuwuIC
Ur8POK9I6tWBD2rHSeNFU6b62Fa6TLUcGSnZ7DYjceGUAuufE/bgzUpgHOX2gCY8
bibvZzIWo7Lm8LLF1pMIigMDxI0fMydAKjtGpFyTL8UzHaAvlYveHxK0Gg9n/FBh
FU7638Cs1nkyiCdRNgDfUYrvPHWZde2/RPmlTqMNeHbIxXYwmgpdztsyXRoBDwXQ
xVx9gbCJ0OAnZ/oTUK6eCU+3dbrZKUufFHMu9AX71AK5soXuZ831nbyLNFTOheQm
QIwrMLYSFut6p5cDbT+ywfGBUPEzitO3pXidV1CyMuoCwO2zUDFTCjKB/jtyE4wq
1M4A3yq2Ly/XIYVhzKAqlfDkf2W1tCxjFmmU7N+swhRpK+n2c5TqQVhM/WsKOtlq
xZD5g4KtW+zUZxcMGBoYyEr2ByYclh8t1GRkf9uSOAaerICM7ZXUTPNlzNrYulnq
me8T1YRVomdrYHJjlkWcd8e+D8xkkMkKmrkkp1UmuRJtNjLEGDlD4FVMOXWe2LDm
blRHjDK65o96yYVLdr9SNvcUhYQW0FeQdeqL7/a0Ur3y4tDq3DXp82N8ctjK5zeX
bzxrIlKSc+Sg/mJ7gGP1CUihzeTwKx0OqXhTC1bpFPY6IlZp6fX3lm1SlDmHuWp6
xmoDCPLGsHLe20BG3YgBITxSueeSyOvbonme4fn+kb6iOPZeoIer1hkZvYtLAMnY
juhP4Z+amS6xeqG06CWgxIT3emA/k4aOqskwdCugeJ7nYgqnIsOuHLyR2pKhslfY
U4U4xD569KY+AQeZdP4cEJ8V8d81wbsbR9NLMn3KubNp1BSPQ/Yd4wwJv7Tk4GtG
QiDJ5wUR4vvZHjJbVlYbzEjHO4+35flmDZCClkLkjxWoH4kbM8aWdelG6Q/JH3lJ
6ZplnGdB/1YnEQjZpK0ochqohFOd3jR4KT6QClYTSmm4TwIW/eGJcjC+3cp88Z9I
d8Lsxoyh2P3iUG8CsH6ZeePby98qIerpXrj8sktG/IsCtKJ43CJTbgP2DcDtcjtP
AAGOvZfNeOSP6JpkqXZPTY+lpFck9FtnU2LOpzkEs6FGLRpQAyfCXE5XX8UJOGMx
xvStGWvUofSos8lOElPOjAy0tW5SgT3e6YAz3SUANwxqTVLRY7YTwlzW19+dlUDh
4dO+CANetCWFuk5cFFpVwbvrbrU8BHt5iIVFCtfaik08SMPs6XH+F1qZs3/SxD82
iKgLkqileaS6dox1VmfDc2gjIrD3MQcBK29ZZbokaRY5QZwtWz9X4ZQTt8C3RsHg
c5Vl8dpOD5nfdKgp9otJOlR6/KQmfzcTSfcFW9ZWUvjZ9yN/bKXQ0fRoEu80Ekyu
QkiVQaz9fXbvrZup2uZUVif+ZQckMPFPrm4Fc3f+UM/bTmtJnkYYi1kI4W9B5m6H
MjeoswoxLZDDSDm0wpmV1F07SFAjMCnUswuBTc5b74zDUPd6GMTo4Q7wKBIt049C
omX6Sk07jatg00WrprG6BlYFhe+y9kmYMSGEWFxi4rPjhIWHdGRp+aWdrBS6TZku
9Z5Xt21mBqzKv/ZqNI8Je0j1VYFPtIYaNUmUbeRsmzAEg5jlX1JqCftFeT3nCt5T
0VbgI821Qk2QtHY+YE6xlJ76q/U6Q2jqTpMwZ2gKhLj/u0Vg3/ZwM0qx/PGdJJw9
f5hOBTIXrFbLd/SVaN8J0m6dVVBdbiOZxQrTCpD+b0dCH8ZAeBqGIg/INpRs6qQe
XZ/SF20OsIiu1KF7442F9bNTcsVfi/B65xc0K9Ih0MGRcHprdhkXT6URvD2G09v/
MDnRp82ARscnqiT1r5+RjV6x1UMI1vSWkMCnCYqZH0Q3l0ocpMcH9y4Q7TZ9AzV/
WbtE6f77+GV+gMGmkQDsAuugXMDorAze1gp1K/g035iTCNmmj9eKqby5D5Zlr3JD
rQ2gvtI+Y6GC8BWzQxOy0pRTR2qxDN4s+7xPzj7kL2Cr1QPUgext66I83qL2hUuT
TZUzU4Q9Z1XFt5Eq2nClrE8sroDDvlhEIjJL4zW/CrIslo6UJ9G7xHl6d42YY0KF
Cg4KRypBj4p51HypK07UzWpB17U8Nm9ETWmJ2DHvoj8ZamU55v5aVk0A2CHzh4Lc
YG1wzmabkgopY7Dm4Cw9moS8BVKe78NwX/CJAnVK8vzx+tOzkSbPfmToqdYMiSdZ
RBnG1m83dPj9tJmj9c704vJ+pcfmGRHtK90kNWExb2LjPoa8zdqUBvRIwRK8Jfl3
jJMjwvL+qZbiI03QenNwvnkUJRz0W++gagQOJPqlaWiJ5Q/4Phr2mDMQ8yJ2FRAR
b9x0eugsGaD6tE2tZqbb2kphQMTepk3D1RQr3q7+P1WrWzbH6k9sPtXCWMJSL3xF
Tw1Fl3CWSlUAzjJGxMEh2tFUOsTe7MSW7Kdqevm8bT+B29PQ2iyOmR3MBYO4JfUS
nDHHGLcIjcPiK+t/HLRUZQkJYfu1PRCuy4g/lTSsP5lesmjLNnwVfnokKPYxFFc0
kx0a9PHeunAS+XwATu1F5aycQtbf6G4pDErvApAlfB2Oes/Y/Zl/5dwKuSNxk7/B
sr+XsYk2qCAvv+EpgUsQ8or3qqzXIdnhmobSBrENiVd7bjkvATxYu20fagC+6TnH
Xe9Elnjvj0jQjxvMbm1/NmoyaJHUp250l4PzbLVNvmZNhKMKDMAKsTMqRnx9ryS/
OoVR9X7lwsZepXm5Ofpv+rdomIJajc+DrTCdodvP7Ex1iEbdqxscT5cBBnAFDl/V
4OxEBXNTyd7x7ZvaRoDNOVEhylvjWi057/PvAZWiIrUpGa9BVH7PMBOWol9FvFpm
JwCMcdmTUckOU0eWMpSvr221zIzY2gULQ/OrJIRToBVlDGmASbDXxzJxNTS/wwqX
wq87vMniMf1ubKRQMKq5eeSjweGNXrcP9ujpIK08pyQSSe7XPn3gqQGzWGhCmhOb
jMbj74n+IgQnBdXyfMLHld/ye9cidntwN1UiGIT9Cq2qYvOUL/xwiMhRWMwYaCvp
ZIXwA+v3zwhMw89Moe+Q29oLcVsyFs1NMCUHroqOFP+cITfN5di4/iqzR72wjQPf
y6enVUsgbY1XNNPmOeyknGtcx53PBTTKwSR6ReMnCgqp3EyKtsMyZU6iT4ONSwOg
WbFjZ5LgLgXGW9jTn11m1a1e4xgBXBREhP0dDzoK3H1n9WLL43dhCKOEA85HIky6
Zu6GEYOXJ/k4bbkXzaD5ThOKdbU8yJnMh4jdrxymWPqbFLZA6PNYHcFF8ADLt1Qo
iiXe3C9DTe1UYkffdXJwccAfI4no+ZUxIIi8OJWD4Ng1Gc/XU5y5n+ECL1BweTD2
iG7U5KBI+te4zUzfJ8KSsbdoTd6I+/dkGfXZJasPMAGSN+eKteteeNNGTvNdc/vZ
iXYfdplU/g7c9eZHlq2AmoWHCiUncmDT15JKAZz26jZOdAzfoabxQ4ba7lT/SFZ3
MNN9Hh9Zn+Ot7vrsHkZIh1xwan6eWZijqGnSa+kZY5w2w3Fi3va4He+FBexRyKWz
9C885FLfVZp7d681Svyn17CKZl3XtCEWKPodnsuKN7iHKt9suKOn8RMQRPuga9zr
pUAjHRqE+caHg9nc1GdNlxCl7tj2ruoKlJBVp7tdC+xmNm74NmJqe9ehTdwjO5q7
p80m8XtnquhNWb5qgvb0JYfFQMZJoP4dVXZwggataN/bxp0t7UODx7xivGBFQ4WI
1BvxaRVkrC6rhA2VB8xkTEhUumZGxoZNxnR9EMj4Syc/Rg/VE0fSj6cZRbzjeYId
vUCLvlYjsWVaY/6BOzv2wUob2/+5EI2tJHE6BTqhDV/Q1S3Rgk4T2vNw8/tbQ93d
aNBvuJnyNR3bWqxD5t+sOLONN9zifZVxM6jeLXRBGK02KXo57pN0VPDOro15Cg7V
7tYN9JcZEXtBpe2LNx1RjkpNbFCHXLl0QU4nrSl1Aa9uW9QcN37gXOjxwTR2xdQb
zzzKeRTCa9O1diGA0ZfBMUAaw9koraLV2+r48SpZ+SO+DGi0+0pAtT5XXSeQ+6pl
Lon/i5flFqWJ/tTi76aDBzt/ee9mA2tvgj2CcV3USVrV7jJCHyajatbFBIygDCyr
i8qwHeFjFjcBysAUhKzyeaqYHLtO5XPJq9gRVK9MMM7vNXO1dQVyxBEBmtsgNZHk
aSQCWVj1I2lMUf6zKv9UB4QhrXYB0YdsvIUbkr1/MlNR7S6tXcIinAjhFAxuPbNy
lu4n1WpDRREYyy6nRA5HjUsSzDw6tl9PNLQSv2IN/JQnABmKZyvijLw0biuSzxHI
yMGN+C11LbIoKJALmDSO8zz/Q/4sTZ/ZZgTSASNJBIQdxXGrhp+fx9YRPRC60liP
y0nMasNX7tGvFrKRgIyjzySmCIwux3UvMD0J2C+7mOdmLBZqw3vBM9I1d3UVOEt9
0D6k240kEbNmCLTkR9QjLOxUOq63dGTMUTxfbEOKlDmIaqiIh+/JFgNW2EnWtjDl
vGnCjkJ6ByK6hynh7cCDIUycmdrkkl7Pq4h6uwm+lauju8BpU4R3+BLtIdP4xJ7Y
qMq/91UQoogK8VYK0rFEssPtDmaV1R+dwsvyjZd8/fVQYrMV93bqBbPvSbA+v678
q2p3qNAFvi1Di2hfcsnqstEL5IJo9uh4Y7CQtXYdxyx3NNeZ3uHctgorzUqCXPrX
+oF3lbJQWJEu+Pr9pvjBLcU0c6RlTaAlcFeoQpFDnY3TJFdiN4UbR/zQcZX9NyqQ
2WlMFJy2rfGLNwmzCdUCFZKVrPD9Tmbpjj0jSXXkfIxTOl91EyamXgGHweuUhFKu
HSjhX/LMglP91xBaWy+0oKh9/N14l/S7qIMSjj1SPT/74lTyiq4Eo2k7FyIEEuhD
QL6kJ55UGjR5OUJRvXHROC4QyFzwW7M+DWsTZ8plr84mt/6lE24mklDE3Jwd9U6P
qEMcN+sg5Dsm5w4iopU4lnTsY+w/w9G6+ug8rtc+a2aow8j9G0OEWMfIfFt0BEdm
jeIiTZ3cjqaMUp0IvgGEtKsxvN/f2kMT29HZ1q7yd7i8MKBhzma/2ZAROSopqojG
jVuDLsFTB9JSfqEzuO2sjNp+/0ALHTaMEj+N6e9qi0Okd15sNl2IKCcGhU2mfsGx
AizNgCXIL6C1bP6uy2jTm9BoyV/QkOgqGt+NKMIFzud4FPb3a4PuGHuAOuqe7/rf
vdj86+32NZaue8JhObJ6IY3+xyFnEkzQQlkd2eC4tZ31Fk3i52/aKiW6izu+AYfw
o3F+tl659h8iAuRTlA2p/uXQr59cdy9RfZRhGHKG0/X7IAoGE4sSNhcScCCIbQez
RLQGwE8NlB3i9mdAvSbHhSebfP0XtLX1fOWS6DFMwBINBocbPUx8tLOjErG6leEo
cpPSRucKZnLwKmv70fM4sNKT+EZgh5eaYj+nY7R8K6fVK6BHaa4kkd7aocH0Bnao
0aQMVkaTmfKJs8snzQAasDfkL5U2u6NQMBDDbDRtjfViqmtyDzEAvEsGBrD0UFWx
sWO8lPL9Wz+67WuNNRQpIZWH+w3pOQX5nhNoN5H2NwaQ5BEth11vC7Fv8xMdKDIh
Or6q0Ot8rM7rPWVnyz6i+tLnB9LsJTjRpYK20wnYR1c7OhP0lnO+mmlzvGfnoWkx
BMs+BZlRZxQ+xAADODMw85kFD3zqXaWXy38zePpGePxAFsFdNF36rGHGM4u2Dhci
ekgwd5xN21P89fvUT3B7hJ7nXHRaVTZBCua93PWcQkMDheAT1lYVnqXip1MYSq3T
ANnIPjstR8Xit9EEzpaXdTOF+ljZ3GapFbYRgRbmx4dZCk4wElhJAlZkoiIP3GIz
d/Ax3SNr5S1kn6gIceu5AFc7Y28+P+EUJtWoHeqYd0IXLMdLb3ZNEWatC0LOGqxh
3OfFxTQZFbaHvr+bb6GgUhmExMiQsD8TFyK4WlVkPOCmg3v283zXImlMnrMZPzDt
u1vuwT5u3N/g+8d7NvsFnRjYQwiRtOYalZZuJTxjJ1Tn8aPZXqgwSFtEN1OhNsJb
X8orPzfxgAgQlDyVokzlCiTmwKOxiZgOmr7QSQye8fTidvkYJ7ZP1UQifCY3Tm3o
4CKbZ5HvvPsRBuYAqUVo1VPQ9WW/Qc11S0Y4AnFrCwL6x8VAKTw8u5nn1vvjL0Zq
LFdwVKyULtDtCwfwrMk+3AsHUPO1LZwycF7csRD08etcrHUmcSewgQ5FYwralv63
ljcytN4TM0rFJLwm71XsYybLQtysG3rQX+Fm5xjq7rOgJ5Vu6BDLfTQVhkrpDUkR
UMauNM1YjdGL2fhoxKX/gV2ecNi2onRwBBOQMuAIdnV9IZYgZ+AvUCYMQ5WvqpPt
fnAzFioA62nr3Y87Euw96jRrxbHlzKGSCOpfKsoa9VTc4/Qobw1W1+8DqmtiD8mc
4138aLQ46+aqt7C0ZeNNPaIYIx6PkykBRoAE26W5HdrRAvIfKD8L1AuETAe6NLi5
XEbo4BKjm6NYIuURTJRMx0nrjwmiRtpHr0yTustz1GFJpu1/GxpwKvmodfWwIRaL
ZNYdexTk5Ix4kn4fmAtfuOSz+n1FuqYcz2NdB1mvRCQ8gPYW7yo6cEAMZKDMRlZ0
oLco3AkE6x+dzOYGXSlixsK2A3ss5oIAKP4aS0EzfB5Bb2geRmvf6bhtm6pg4rcT
6babH9YhGn2QLX9QxXtKNsrVVJ9EW2XpCVK/DLifjY58Do51m6bqOzpYGLsvbDS5
4WQxpPQN97KwqR9/QFA99bwMiTzBXmTJddOQAC5JXWIXZazJEofD+CMQqbI7X3Rq
Yw1LWyVBr+1gRC4E3qduEIWvkRRgnkAJoOH0HFkz7FKqiFzBg55wPfmYYD3Se7Eq
RBMD9+qtYFpcxbXbMuLqNLz593Za29lOPFqV0jMesnMf86CW6s7PsARyO7eNpPrj
NR5fDlLXGv0SD+/VJBfYi6NecSxUc5+VphihT8ETnkN0aRWbf4n7Ntq/UXZhHCbq
6JDjIyB7+m6YajYoaHRWVxFF+KRGylnCY4YUUdnXWPmnzSDnSJqDP/W+cwf3QYm2
S6ex6wsRQNCtJZfMtHEl3fZYEy70vRE6M2qYS/oPwlxLamHwvxi1xfdQNj1W4sHJ
b9P+dS8YL1qB8HwhDMlUGnrA1efhFa/gN87bHmX08wC1MAyeacKZ5VSe4GVZCAre
5p5YBPS6mBlDo3dX6Bhl8YmRRc1LMKFKrv3I++yz9QHFSw0BmG6eB5FrapgymsCO
1zT4tU6gMO3C9kkmDHTa6bvCAov879hf8Phgd8enLQ7KKG5XbBBjHhYcntRSUJkL
WPG7IKJftrBZs5+q8rtCz+l1mrs5LGN/G/w5Fytz5W2D8mHGvWeDoBKNPvK3o6W4
KlYj3gRZa2cT9dRFM8WZ438kOLuOhdfpEBgONxKiybeeMpNFwEKMShcbmc+U9ILi
lMUuRdsY5YuFUje2RpuF9RA64RC1jAOWQB/XqUotameytPPex+5j5imlYOED78Cd
yPqkPpYQI3ITCQgaGvb+GEurWQCGH/LtxUeOI1qR9Pn8CsyHQWBsrFuW5DmodMpg
P0FH7bUhsrRZ9sfVYKq0NNfyYeDNw4tvxMD0caKAKDF4p0ODC5AvvdmyB3t2XtQc
dsKXlOL+I0YwBhN9urDCFLZMg8TgXh6+LNGjlvlbcifxS0jvW1TBbdwmtuKywzQf
lXGEEoKLQdfdMTuC4vByuouP786cImOdpMqRld7dCbfp/70sZOf6+oMvkVnXCWxQ
yMxztUIb1R3rs3/lncP5i6Mo3S9adw5o8QN5vu57e+UGJlEWDF2YyfVG0eE6H3Re
uCnPIiGfmwicb6mMeysFD7yhXamxEKRSlNPVY1tne3kOB9FIoC0j+9gD6qiMlw+b
BrjvEchgdAK6I6HkZGKzCc4X9umuJ9kOM/KOSOWRdJQOgpFcwuDvvQILRp86X6WO
vTIOFKKXlg6dIjwugZ88zTu6bJ34DDP91hEsrT6pDsaWGOmoj6H43EgmVXMlNEwX
RCKEwjLyxxCZAbuFCOxrbR8kDHw4CKZQwk7qJstqN2yD+ppobRwBOXxu6tG4GhDa
TaePSCvvsoTT3nWqcX7Vq0ZQjC8u9H9l/i+dQXV0FxZ1cXg9MgurZzlsmpq496Sg
zPDI0Rmfgj55CTnKhsRnsuEKA++IGbxniqg6YVCFQdW3+tsL5/QC6FvjKA2NKo6r
rV5wp2hZsqRTaCVh60y+7HE1Sm+fBvWl8efhtyLmllmLOyfepqf47DuY7nizEFC3
b7JYrjJ1YbmsZF9lafrWEpc59cbKJwXOwtGUIbsimwzmfGb1hsLaXvogPxuTG5lb
tz7VBdFeLE5PIpy1wnKSh5Gj3ndB73HUDY244VBWtrHpzxoecebdVEQeSJlpFDnO
iOGCfhcsc/WKa/bASFS9AYv+8/b8YDgw6Do3Q+hk2315muaP1sEBc3bmnuvWx+Ch
PY5Xs9OATUWHCfrA0Y7kvj/xZJqWjj/MMDcEMewdTV4vzHsPj8yHCEYuKXRvymvV
BWj8rQh3hdAmxn9fjVguAp+I6vviEiAj8GSFcwDPZFiNwIVYRuD1CRLy1rgQoerC
q7+PmFVBDjj5POwcKA4LFcRkMVGhf+yryeYgXSjLJCYj3IDw6fi4xlnWhB6PYbB0
58hOhK+4D//qLXDFgYqZo2YeiK9eT1fzvf1jNT3Krn4zyvabSRW6p9+ANc6PLh8U
iYkTZS+xLCk7EE6KcV72mv3kKDtN8qLC4tDqe4IGtj2ffGCTPe1R/iZobSn6ysW5
shtCDf3NwfJFnLwJLxwRPjINHCP8Kx1LU+TGOXDhm/HegQq/akTBobJU/T5C0W9Y
BfnYxx2+xkJB0OV09SK3jxRCq2fFu5gs9EOBNyE/WKetlXCS/Qy1P9OJ/EwlXEqf
ssJWJsoCjBfoFvjrvcz1RMksRLogm5aMPuQlC0FFNTwCTTwv0Xp9I5MKvA4tWmW/
BAL3xNH6uw3gvlDp0drJGWSfqEU7tmwJhxdIUXA3XVa84xh5ib0+ToUWJudLn/ac
W4gaMr7l1XqnKmOLTPJSlmjD4+QxpodK8itdgznahH7zbiWiPfRFk4ERHSViN9cW
ddHtUGuZHZR5cF9mm+75gSdZVprN3aTcBZinKxnhG2sn2xgt/0C1KDk/JVIS+Ca8
5Yeaso2HzUs6pLsVQc5R3RsoIP67sa0iaUfDQESEY5tCxFlNs1zxzwo0OMS/AlzA
BU0P58IOSXVgXL0HkylYsCskDFD9soyOZB+5UILv7gLmkqgDJEE6s0QL3PxUpVKZ
8Jy3DjH1svk0gFx1Ckra9vhhAOOSUtIF3rUYvEvzkofRZVZLQTFh2teKYF0utK3M
h3mu4p67gCWCO0y+90GHPUdtrBjK4EuNwzteo+NKhxiMLm46QtSlF9K8tKZNaE6+
csEvm0JEFfz0V8hFuRxd9ZR7Vgivp0nnPNHQNJ/1LUoW7FAvsZxjvJ74Z8RVEmDt
WPH2c/QeN1T6HSDngqDZp6BFikZhI+zN1G+f2CwrYqlFVvU6trRhVh4JvrmWi34r
o7oasntkpVznYgzVyMel66jYpyG8XO6G66iWT3UE+HkXw0mE4MletGN88der0ABt
7COjP/Om+nQSHmyXqAqsZXQFSJN6vU7R9kW28JCIq5RctEnCaIcIK4EYuYrqBiLE
Vo8gBmbeUf653DxvHJOxWTG7QNZcQrmw5RtPAbVC6myVkZ/g/2DErEQtH7D4i+wh
rwzWMp6DHdV7HCbnd7HlFu0VIicIGqOOUlM4NeobDivDNWGTB1wGW9/4YiEXLeZ6
1oG2HZyHX121JQ9AxrF2WgG1MLVtu9fl0rV9MqlCSTnpANfGT6Gw7/z531fDVX3F
awX4Vrlc8XdaIM5qlM6xLBZDPyKdt4XkiPYdBgIw64ExBwRWBG2cmHQ14/RNezsX
MGZUDiZk0wmTPm5qSsTImyUzODJB7Vtz7Lqi21q/T4a6KJzo6UHFG8+HGR6T31rf
PpypC5h+dcq51BCFpQQOPzUqaI++ETWApJjdcuiijcHkbU9O2cFWJWmXLFJI9aOe
NwnqsvielMCue0N0KRxIGEVzSrghXxa/iaf47fZpAaO06p3du3h0bhVk6yDP7KjS
8qXohJYqtMePSmlHXIqXdVNEs2+Hq/Ziv6/k2HN6X2uJhwSJM8T1WHoHZocKkeUh
/LLxOVZOacs+p7vfbutvXzKnLDASBWWjl3R1Q7Tau2uZ836HGZ+8TtekQGMXNkoW
euLUApWBocPKe1RfjEd9FdvAfmhde57v/B7RUXn8eswKrst7O7OjGPIYVaVKf3SB
1DDplUNVMRuO+Jo0Q+Qq14VXT1Axn8G94srIHpXzVhmFpEcmXzJHetkWS01Ey9Z3
FpVItOXSHORuvVT7BaYkfCtjLjAeLxsOqM+3YA60H25euC9aX1g3Gb+R3HuqWjBv
LRJ0iyhfICBjv6yzj0wE3h55el1dGKHwmBM75vz0Pss4WaMNXIWt2k2lX7Vex/dj
Ya2f/ujuy+EYEjseVa8kz9hoaC6/z3mO358Yqxvke49YKAvhKfYDCJbEzHHHm6B9
n/dlK6QoBCkzU34+iVd62CpS7NUawKHnxPSRBDmq7B2+PGHnZgUTDJEELwBaLsHK
T0oXJieGxc9a3y31qcaaDhMjvNplm9sv3gWlw44Xyk6Cs3wo+N1kMYZ5FI6kY8Dm
nMAI8Z5XebsxyOccoRavuk+I8SdlGHTCmcDSJ/JBS7ogh2nqJIFjPox/Yx06MPNQ
DZ0l3Oqoo0crcW2X9ph7OYNGeT6/xf2NMTy2WMHEUw+FCRuUEAbxlsD7N4LRfr0E
rC2usF2/nzzziWY1HNBEai44J3PFipmaV+Hexoh3oKGvh5i6AjGwCnLAsPMtsgbt
3VuBoKSK2kTga0n30j2pfLJyuy/BCwC5lR7dm3akdCFVCqwr31VfpSluN+Qsiw5I
g+z+pcpzbCM0GoWOt8JFWQvmYqlUJFUAY9rcFTPWIQ+qcp8Fz1g1BQa1pbO5UvGA
nXrwlpDa1Vtzxe9huzffvkp3KfAN2hl9MzLRvl0b4Y5D8If+rOuC/sDRt11Chstt
VUQycWgW1hX/0rz/vQ730ApcyunZGAR5JBVFMtc4SjC75jN56NALLQGEtkuDGn9A
mippOZzWgFg+sAnXdPWvKpto09NFWpUlKO6pqhYb2gIWOpKfxxSsH9aAndT7D22Z
BnEt2RmwQlsIqhATEb6JiCymFbdI6EsK7TaCczu1ps1sOcZyPKS8RnFSZru5+q6l
eo0effYSG8AY/vkSS09uQs+jUMEcAuf4STil/3VBNSStV7464mcwDESno6BFvQ4/
vqgCzFiKpVjqzVgVKGcl5qqY+xPub/Oyw5qNDVNnDcLFfxVhvLStU5+r0PoaPOTm
g12VLI2Iyt40aX4Quok9WdP2DqP6O5HdyeGFZXoRgxy7q38w08ryA2WoK7eLzIFT
rVugfYvmSkmxdF3dInO4X/Rd9pB4aKWq0IBYgSPjziEuwKBq1zNz29y4flyV7AU/
aci0Sa/Of391JreLJ5ebRLPUlJu7h2cIierJuxLVZphyTQZgqLEwrILeci0z/pZ+
76lsTQPVSzh6+HxW4v/z9icvm/UXrV80v5f5C02VB6PomuiEXA6QPjonK/HbAEJQ
qZBiZPgmFnHG21piNM5nJb22YuIvjXGMBN0Mxq/QjXg4CqyTdj9yEwzwA6MkbqKJ
gg9fdkQnLHVzbkMRwU0qfBSNHKWLqHZHti44DWBvI2YJSlQb3YeJ9u3ReCFd60YO
lZSdi/k+krmthcosiNQ5YyiPCI+LV+2HmLigdxtlvoc6y9anRwh7b1YRkZIXlR93
j6FgvotYHDTJWftxF9mvhfwi5AaiGVx9p2FLpVCV0izbQwYFktZ4oRJe1+wFvWB+
iRqtGSa4AhsRrz8lLSzV/9P0NmLa2K/7fwzoxGS1VvVkybklgtsiDLAOk+wBUK0J
d8tRmMPrdjqPWSViZXU+o77ZI6pSsxEr7LzVh/shH4L2RtLvWVWO1ddcDpaNsP6w
nKZjhfLJ1HQU9jslglDUPe9+qbVaxn9JDzLqbGVI7CFRFcikcj0WbsuGlw8WvwFl
NtXCwigwpRZdtJbM2KLVUeHumIaBrhKxNJZXAH/3hpWlHME8OcZ3+K7AOFxTihik
n2wjk8Mkl9Y4WJ61GPRxOIOvWE0sPPqbONFtnHWgOZa6Vs84BQ6dT95ZUzfOiZDt
h3M6PthbAUQSEig1wR3uAREldUqhv90qD+XF6YoQt6ylDsqbqkdFysm1kIieWZJv
yCcNXQrdlbxwqyGcMc4Dmk7kNlwc6tW79AOzoo3L9SfzUjU8230OHXUV37WNf7dF
5j2h2xJ5r0SSQAfp11wJgrkg9AHJ3HoWB5Ghm1KRktyYqH6KxTyuNnQhU3GIttYY
izA1OSDmmDeEbjwpLta42K134u6fl1OX/kWebzhoGScl4H0Fs/UCEuo2eQSN+chO
10Y6uf8H76C88XZVCAlck5vbtd+T0Az90GKS3gEqSP7kYtWowMBEx1mumnNQwgI9
td+rAO1WWYKyaiz+tuqzVaUl8fYGNrODtC20pQeZ8CvOo+K5JH5rHx4Dg14Rp/P5
Y5wrjPn1K4mWaGcRaRInWrOknv77BnzwaCs37FqCiehFbQQHr1GfePQsl2pB7O8J
Yh5ae3CmHuuo5FV1UnelyV4zh/AAcYaU0CUIcldliRHp70YNpR9sxrcYKEhlu5S/
9vpsJ+TpzRk+B96KtRaQNT71kuV2iSMkhfUZMfrKDSP3k0Yl5Gb0LvB9CEZovhbR
17ml/kuBhtqDV2BRh7gO8KiixhPKJjB8fy/8maOD3nZjKXBjkMO+awiKTFNqbQWv
8j/z4l/BwF89NiWEuFJR53Bc1IKU/L4piMHEkHbDSO9hCve8V1c29kFhH4rhC2Tg
ykTNNADku/MseRdvq5f5tN9FUaciZXOaRyb0tFa1+KbCHJuoJV4TLzdAHw/aj4UL
56VEiA9K6Yw1Ujd5xjTcbeNvSBeyjfTr6/gQNMBXjebH+ztP8gQcY5Z56lSSadqr
9oB2kWvZZI3WIFKCqreNm8p1i8FvZVJMUMGfAToQKXoDIfoUFOhBfA3loolVY5sC
WJ3vql0rsPpaPHuKtguW+pTmq5cRtIk8juzB4XN7XXk8UgKRUZRX/9sJc+Cmmgo3
SusJysKbCJw4dVGwCeLJhtNLhLgAAfvawJ9GIvsWbZVu4NJER3j34GcKI/iAvoTd
VkvGNMDMaWCCf3Mk8d1NdY+XqNumAtm4+IhQNjX8+JDc5t5ZjG+MyFHigwmFN2/z
/nHlz7S5BV/kK2cWwsBHguuDmPYBCYBrJSdER1lLCUDilgp8J4uje71BctFYDafK
bopZu3/P8byBycDqAnr4FVkxx4CM4l9/4NAiVENlV63bPJU5jyIOZeAPwDlckT24
19VVHsDdf8XWoM399x7I8y5YcvHw2w2qzfyRxxANLT3HEQicLa+JqzEmm1QTPpvI
1ARIYqASkMQ/FTIhWqaIUYhODqw2L0dest+njtpsgD8/FZNAhJrKmJsHpdRln2lr
+un8bukOcN+Dou/Af0Kv7qbIgCDOSyeYSAOymKQ4JRpTPztrUHIrPTDCTSEHen4l
OtEWZL+r5lDQQdXwmk1sdjH/6sFP9evliqO2bVDA8fkAUVFApZ0wl519Xj1EX7dP
uc9KRfUAPBg8lIfZ8VstpSXZhS9YweOpm0Mx+PhwLiWTSMf7AGezh1LGSdyP7D16
qzEAF0sB1U1js0u640axIj0QymLxemRJVevY8/6ciediB75uSPCH+KDUqYonYSN8
VK0X1zxkRAUM+E7p0WrJKsw3XVjOjX8EL9T3Eo7e78RX9tAuVynd808DmjAT5UKu
vxSHDnpsElw9s8KOzlbzozNznXGjsaN48pFCNHm2orLcI52jhB4HMvTfXaV5z6xo
X+n3rTkRV5t+kWC+IB4PwcMl8a7S3CZZQ8qIIc54mSk4gq9Efi99WJT9CQHxXQd9
6K8ddHn6SyO+Mg0SXy5Ntc1EWlQvkuGrcZf/KFxtxFQsCYATsTvz9rVr9IikMU+L
1Z7QwvG2QnGKCCPvaPnFE7NzvpIMBaeoaM6nEMn8LQZTiUFcu0RWy6Zfw70R/SVK
FPYBFxgASfy5qyaZiBLkvvhlaRSJB5ziHA1KgwhvytJBDP72R130Ep9iwqhOT5/l
zNojlEaLq6dxjFh56ef+bqBTT24dzsFFHpFb1hmbiUk83nV2NvxWq04kLxqT3GxR
l0VJcb6nP+sE7AryRnAY4DlhH9vROkejmscVk3DLbncc5u8O0/5NUQ/sr1VOaaQR
jxjLc1JclqbCDU7CMz01XgxSHBqIiuXW0VZd+Q+Nh8nTKzkWbwGCaet6XF/tU/6r
CpP8O5xC1+r96jtr/MFHGtJEipeCkROQ9eq9tctCJUuDrSP08P1x/UQSXQVaIKbH
HE+4AHVOQXZvPgbJCYHKiYygjQ51KuFLgI5DJDnMSKe5C1T2OSXkr8hIQWWtxMyB
Xh3/XrzO20fTMhGUBkjYbqq4FTIejjtps3fQs/4s1WKcTPNagfclBQCnX5gWAjhm
RwiRYxw+YFDAodeYvMv4WwkPAFfGJ/De9Bz5+zOnW8Lhz1wFJJak452fy8whcNxX
L24E0t27V9eTgJyJPVh/OYQcXyu+QD/74et+bB2Ko2ykHVVxz2jHruyqWMgGPMrg
T2+fWBgMk6bvzQIFwb3ONAQG+FPfGpEXKJmAAt+S7qwJShGun5dmSAPKZ6Cv4h0E
33PMx2ReD7jnWmz94Z14enCB/dVRmxPZfxRYfoZVK2AIbeupYU3HBD0F8eLwwbF0
aGOoq2iNu4TTn+HYGxb1KcuopZt2YFCWX15qblDqusKMlCZtFosnfw4DR67t4gNx
nOIC70g4fLMKh2ZS0956C0KhBXPoJtGnRXxvH9pWHyeaib6z1nHvqiUp0yrzg8Gv
upfLbcmH4AplAkHz5sPr2XD/yuhk7WcOVihHPzqf7ysbb/rUyPwXozerex1SL70e
vU4NhN2udyJnEZ9oeUGRPrKwwJVkxtep4BmHPPgTy304FXD842pEWPM60gBae2ms
8eTKFYhhUvguD/L0Y92z24M6PiJIOIjO/QmiW1FB9iR6LrhfSx2mOUTyeyUla9pJ
Bn+Byebztx+M5BIN7Dc2fpsPIeY9xpZCU8wF1ba/yNCrCIcWa9shZE8DSbyEhWp5
Ai06mALM2vyD4mW2g/sbUTC/+aPUpSkhfJi3xbLxqQZ2bpUwYpxGaIHlnv581aGP
HAK1GQIq12B1bYKll2tfTi6ZLSdufW9n8x86DsTFdY4ObN3m8azdKheSh40Z/cYl
xc5rEfmZAJdqbgEgqxMFSljefh+QKH2+Z9huWt7iMcD+Ul3OToWyYfGAWQFTyqhZ
MwnG+KRHsq9LwRNpLhhT6z1SbuqNGRnNZU/uLWbwsFhfmfmXhi/ciT3ujbL9DlSl
5snZdvyjD7N5gZnpz7sXmTMEJ4rtISJ0uofFaGN/f02sv8rCFmfuKmo4QPpEjwWv
bMqzwYe5rLiJFDYjeAfsqZcCkn58JvbUwI/t2rKWLEWn2ZI999GbeHYZfs5h5RhA
vSef/I5x3lyKT1M1MF3zDGbjvGc9FTHZXVLsYnFLqv7S1ZZ4nIRMwgYA09fJTNln
bVDxh7xOcc8+wpQrYZFUENZLm9ZxhMuh406ILqIlIQkiwdsBkQ9ST3jKs+WXqoqc
Ulk0YXyzIwU8UF/54TLqrQrVh62R26eUNBu6CRY9HqnAyTHmZxZA4mDa6pKRN20M
ff6F7mfyckd5ZsHP/UnyFUMgOQSVShdEeXtzSPZKgB1tLkErnILjHdOhNUwBfOjF
uzEmRSZz/9YeYETHM0BZafyp5GT3G9SL9ZLZqUSzwnoaQbUnw4WJBD1w17wyPnsG
rFr/iyRq6oQ+pg8saJfYox5Z/2c1l8+9FSMivSn1gvgP6GvAa7UmiEVxNYp8Pdl/
EPLaxZCUVw7HVsAkxMvRy17KpQHdmqGxFFOZwm9RtasBaPTC9znf6xXyEcqpNyC7
atGOklxESzVITjiqtMY0Nl0q+//WeA1kBwkw58w4kVmMk4wvTdVS3WX7OikhsO4a
B2uEtnCoBEzQ0r89rdHJBcn/mk/WMyRYrz2IUKrvbCFt3qAAt4uE/dHFugFMajkb
4YkqMKFtr+zHoZdp7ZZsKL2fp/nFKfztl4FP+QYqCWdJFqbupqbUXdjbtDMFeK22
KKHL2W32oCYe3F3NEuIjl1/sRPIDiKdGLxgoZDd8di6R2ArCNJmDPtlgqP/4P1Is
1oDoQSVVDratzgV90xv+yRiMU1rEyhqWzDpQdM6OXou7SSe/4Nw8dsgzKHjb4wTd
vxv7jz9p8qjiR2iTkSzPg/PBc3w3fm27tjES/sJ0aM6m5qSqjp3ME1QiADPVABVl
Y8aNSpZIpISroGQ9n+Nsy4Fa27tQmmg9QtOa0xhyzeMyl4TFfphScs9c/wm0a+ky
Nfx/Nbs/Czjw2sTxPbrZJsdQfD3FORQDwjmz1UbBU9eBZSnSeE/yH9bZ3KmIq+A9
uw3Uy6tonj30UtT8yifIRmxrSFVeaPrcrI2jpmicvKV3F1u0Mxbq7VVHnMhKdRiC
BElKecaZxZmi6xI1eFJs/tdTEPL1qVs0gsbj2teNzke9rJ03uuOVXLpyzeeE/oUp
gRYaMV3FxJohqOEkqN4x/Rgc32Cy4adn0LS8a2l+HM7HBHCCVnR8GjR4P63/l+nh
1jdZXxEwnsiG/5pyhB4SKYRmqfNY7WYlzx9bhwEM3KqoqVjwG6hrtsym9yBJNYIN
/c92pwTCLe24FTLluroD8Moxr0JLzdHmVN9lsiGjQgKKwSw6yC2gILvzNCwIIcuV
2uP/VpDSa1gzhdgngfg1g3ZeCubRH5JOebFFlwrXEJzYIK7LgeNrvWoS1Q6/4B+7
VFIJUtpn28pqPQZwyw2gYCC6J4Hnb+2iJ4/J8geQmbfo4Tvewml7sjrVv3s5Xf1c
p9azVmb0sjxVrZbgY+qKXuoZuTURmzSYbAetnbt9boiOSO5uPGuT8C8O4DUK1oPv
fc1UkcsLoUhdekrr3UuEHjqX0+aIUA/S8PuZgEZqCQMxxEl7uiVyYsvafSqzA/6A
3zsR7J+N4t5AwklNcj8MBrBjjindrQPs86ZzEXAzeTrcidyF/S2g4LzLjhzQeMdb
mXSicygnY2ZhTw7nanLuJdwjVq1Lx8eY5frw7+Q8HHXw0tFuI1Kg9zTd1b8LbWI0
QCrl1mmHI5Npgse1pWZbw9Yvosblu4dNMqnLZ/UCF61oF7Vya1KMS0LR9u8/khti
Nj/4hGHWQWCjarov/14fWtCdu0zVugdohxer0dOaCf9FZdZGcDK5UGMt5LoAtBtj
L5cPgCY2hXr9sU3phnNyvQO8Rn28dSBsMMhiLSSgttJL7gxok3ojxYDT8CJHU8pv
ZzuoTukiQfh+onlaGI7CnggGFUfvvQeoOfomlgvrGYEFpOq0bIC5aeNtMYfR6FXb
OMSjEKo4fDIL67HVIYsQN/DpWhO6A+xeY+cii0SJP6HG0le02U9+HZoZm1Li28X0
sybmE5WnEuzRA0RQsApEf3E9xGNXgyXSYuRKjGjtFDonMb3nNEtngQu0r02JoGwE
F70eSIBSNlKy8c4oWe5vHe+NRVf803RRpjEvFg0jJeDo/ma5tdLqXmxAx4uAyPQu
jMLAtLrCBvBjIJflysg5McORWIpgdqFg8971LtD31FhSgHyMWQRMBXcfyiLd8CiU
WJgv25jaj3aGVBSlGw0FUSjRf9JZSu7CnVKT0cKpHeQ4XMzr0oQGDL9dc7Wlfy+B
aGpuGtgMT9UUXCMEHr2q5HUTUMkjXdJwGijGHQ/gHPWgLjpK0IFQ4RN5Do8puKNW
/NhNPEckyUr+H273CBWC6/VOUMwuvUkOGian+PqJcCvdoYcAd6hjKT1BdYz6nL0R
Qrp82HWBH8Y31JpcSyFCyUYEOca1piTy7uP58iSVSCr8RHdGdfNeWfoJYfwnXoAz
nrl2W5DSp1YKw8Et3YVO1GVE4WAN37IB3+a3Icxm3Kg3jIsFQiix2+F7OCkaCg6r
/ShPC4WdUBOkjwt/QrE9OKC6IP/rV81/M2Ef8GyfXMz7DzMr31wpUaB2+og2l7PV
l530SKuMPSXzoOngB94Jb+Vdh/OBXwLFh9yBpcfviVGjvugwU0u9sU4lAY3qW/0c
xFRNqZ6rUIdkCbciaCAo2PSssLvLiC4qC0LFBPPxdIVFIzhPR2zCmY2GkFjhTvyp
5OUV5j0VahQnFc3YD6++QVIQuJyiQmqGHG2OVo+86oaWhxtus1rOFpnnbgz/HQH1
XZJzC55WdcMzRKaK5R7crYv9Mc5wRNphZP0g7giGjPm7IALg/wMl7UOdWuDCTOcK
vYHpvD4rGVapxrRZtRZLgaxHVxxrfLjf91i7uAjesYMSgpvvnletcKAJM86yW1JM
3JYp+upQbRe9PxErgbxmjhQNwdcOROC3ZWPKJN1CjsMj1XB+sdeUGzy4Gpb+ZKeB
oYW80DLE4RN0sTWnKFaLUxIFSSzjmvuQjTHnpbZk/lnfiMp5ySU8MDkHA5591w+z
VrSbKRnffjhoHWiHZdlZ11m+86h4WsENF0N1O8G2uhGGm1+g919gNLS6ipT9fD5w
l7aygEA++YwimKAUw9LAtW4DPXWRqJOemrL8fXpvGLB+CXT+937NNUOsZarBV3bM
Fm6w/nP56zoMQ20z737oiMZ5aehjKPISEVyS74XwcKqWG0xaXfKSktXnU8Gti9sa
mTwRBVexnqZSerKV+C5N8DipoPh5i5G3g1ia3xM1OOEmSiZWwtMWzVvv7eFD4LSf
E96oj3+R3YtFnEmQ8yHSOanIQqz8XuutDVlCRS1/e0JdczHCG3LP3KFK8e/g7fkW
a8seuifV7b+J7dE7kKsi7IsKlIs4hIWzdQHSiBSeA45gxE5R8wXCzy0NEv1CYAKk
4Egg4nXXxySYc+PYH2p3VdZP8jvlJlrGr/jNCdosuEF6k9YWcXLvD+zKVyS/cgGp
vk12EsncnRJauXCC0zfriztqI8OqgFqozePG/NS8U3wt21nUZ8AcL8lQ6Jchzqlr
rb/cMAqLInWJH+RTScebMuJZ2W+qKyN+9PnaxawNJzLR2VRA2aV8DYHTcP5fRs8i
279u6iAije3WYjVAjlIaursovPsueTHHegsa5aybqNXAzxDDO+/ZsqEKx+xNwBaA
vbl45yTq1GRfsyg1FdaijwBVAMg3BYhAiDcLWePg+2PsiDGgtzLSpaOUKytN36PX
kXGkRKkR/8VyT5fR8a5JVb4ZOAvj4aohLdsyCwM6O1HtojDVDFTo2g/xn8u7RMVj
D3MqSIS6Tl2xe3BmQhQbIBjdcrgd+aW9TzWa/gDchssG4BCbWZ2P3xFABqgE9+SH
4CznGojTFcnao/0+953Iyufb4av1far7HLRPm7otSSBiTaHjKP7FoBUobF5dsUZH
XR1Suf4Bsd3k+hn4n78D8ttb80mAHXJjj7OL0p0CPsrS8nElVFhJhDsMEWZfSP9I
3hah2By4o4D8HjzZcG2y718zc8TgjVBehq/o9eY0SNVZmea00KCS8n8pRQ5PMDw1
VTeGDvfAEbMLZDk2GqPzdPi3ogwrwpahTLUQvy1X2uHKIh2waLn/vcgl/+dXCv1+
fjXePA7EPQThlrpg3FDySeWmQXBQvQONQwytzuR8nOC1tZfjW6HZIMOZYAA5E8sf
ZgAmUEKBmzcMOVmS7lUWP8gbrllovzY44/qUQ39NdKSa4pnkCgoh6CeWi1bVq5b4
fJ4ZUg0hFJnobkZu3GKb37GjmUJKaEfWoZpcyUnmb3eHMyn0BcwYLl+xNk0tBZBx
2+nZajomK5z+qxD7cW0xPqmo4eMbwTHxLtZHCvo1rff3c7pqf60U6tAhpEW4WF3q
Sxe85LnR0Peeo6ARhH7uBcx7uKKobb9R6s6sqEqL7Gqlr1QCYyDxy5SoRsdUsiJI
6iqx8B/gmxXaUx82lVyY/sd+D45ocBPXsnOBr5C97xTuyJyYdp7vg5xqZ20TYAPA
uuPQktGwMSJlK/1c+5BvqVCmy3Tq/fP+xn4f0kPbPkmny5TyDF+rPBQjBXnkSIaX
bRxF8hiPsOUPcETGhEJgklaxP0+vwsc18NKS1xgirvClwgAeyYxhXY4mAGw3ogsH
TPmJVvaNgVRY/iCeoSMDQnxPv6nbx5nn6tvjT8j4cVHCVDVtL/RtC0dl5J83GLog
JHGOMixX2v+qO54tuKYWOBfFV4PJGBqPgnpcQrEtkWY7NozWuR9E/BPk/MzP8f48
u1GqGKnn6rgc4Rd+KiLcza2SXz+rphsyuMLrO2zHEQKMhhVjh7xjwqKj/tcFxwj0
qDomYVuCzXnHG6z5y0pbB8qcXjaMVjb2PMBe4o+3tjJwF4CWsxU/y/V+azdSlcMz
s6bLp0eBoCDkq8RaNdjLFGa8eDrXOR5U+EtlkeGiVA9UzjJk43UQsSFH340SulWF
pWWD+WG0n/2gTa+mRBkimMRKCVSJA7C1k789QMZJUQrH60Az585xQooyCmbhgW5T
NmP7nOK4jJZ0JcF9NnUyNy27NsMI8ZxC9yBVHGsP3xNes7IqZLTpTixfvGen3ns7
vVJ0u6qeI7avd3/DkqgLzs9KZ/SV+wxgf77RExbctatjchLvnagDYfEH9a4uHk/e
swNBgzEPpS62sHLaRzNIPuVXxIPSupzANRXnOmMjjktCEjmcweXS2SgZhit09gIn
EM58LVEg1DD8ftlwhEOYQtwagBUhSsFDLw5ytD0yhQNMiSGOgWoEKa5BoEbxN7HQ
mLHmfizPrhGMwJIiD9FkEsMx+btnEztOHMekoNeE6L/WgCndi37UFPj91MftFnBE
pCnnJnKKc86R0jnyCS0rRbKgbYjO9vSu5hoIYX+j9AvY4tvMzFK3NS61RSd3ELcH
dvYS6YyyACoe+bl/RAfh5IayxDFiRafs0KpTe6phPltMPdxBhZPD0u0Oj4hbCaJh
W70C/+8Fibt7BdGVj3gsNOh8NIkrRjSLoY/lMvs5FfS/7mEWQum85PzZxop1LcYF
vV13fx4q8ukCyU00TmIMigTri4wIkgYQVPBSEntjjHzQY2k6uTcBIbQaS0Q6q9o7
OeKZ4Mhzm+3/EqzxoeoOPlKfK2uCsyUg/oTpAz46pJnxRkPQ5q5Gi7ifGU+msztS
4JRZgAsGFx40cK9lhRMs7VNHGagtmgytKckfAZm95KMZvRb0mbIy6IFETrpMeLnU
x+GYgNi5l9sFQKvdX5+JDTbLhFGI6b8cQEkd5KnKPlpX5fwqm1kXaAOdPpegX69v
kWBycko+WP5/RwshoiyuGH+oJ5RSvqN7ZceNJyiDdpJD0vLO6l5JdpfPoW5nLBRb
gXu4Xa1lZr/tiPuy7GiF12SuUXfqdGDOt/gX1HExkJV1fkbHwwXPIQqHxRzActur
k3Q5SUezvQkP2HcWAoIEYiVmHei7wemh2HLZamzNv2XQLYQmfHNazWl60xUCCdfb
bAmozZLSOqXZ0o6ZhuwbJtCtK2LI25a3NwmFC46y2jdgI3JAU2teUpnUB0N1nGPJ
vKdzaWmw2dlZ7sPLZ2/KP7RAdwFMX78Ja/DAF5WmYjE5EqHHDtuK24i/fY1MP88l
Llj/T+xVvmAHpY4AQWcJb5wq3x80m2VQPVfVe/N7YoASphn8JABkmxWbVx+/hI2I
IB+KDMCjmys0JuGW+jCnk6nn/aqaCF8aTfZHuNgmacl7ez4IWsV0fWJZiDoEJB37
GTy+NYfiM7sT30BNZaEuDvL9VJNr+65XsGugRX1evsYNZR9ps1bZUxaP5stMGbtb
8urlNz65x47AX93suMgNPUfG5IrFz71+jvpetLWCMswduJPaXldT1PR+sJjBTyxs
6uhZoxtGQW+EDh4DsDvvMTpG5AiZ9780u2NRP7qhqMRFxZDeoPUnZk3/d8D9d/Sg
i+wKk2IbWaVqWdTyFqzSZNbDqp5V9vd6JrtWtj9ltgsHlYTMFB2oriQLXF1dpbXG
Hbef3Cc/Is5vAl5cfQ5MP360B43h7j3isgC1jATZgTUI7KU6r728xKj5afr/Wk7f
+r0MD9ZbvsJ/LPgfSYKUYmGy2jvPJryxKo/Z4kAsNucfOBUsZR405Ut5cwnYLows
aRTOQPi47ipuU6W9vFswF/+LronrRa0HbtRCpMBZkbRe49xR2+1gyLEpXU7zdNql
tOOGsthqdtnq/1mKL+TiPWdgkWT9UpCCpGT06TyFsObXc3jGPKAUNavT9L5xz1rv
J4nqQVkAVqdiaVfGUK69QezvHD1yZpLIOrhfp06FZxSM6q0mg516DnV6UtREtsIB
XkjhO8dzUIZ9iVRwiLtqJk05IxuzOh+n5YXMjDqGJlYtGbaMIoCMlly3eKuY26dr
h0A4LX/NNF+lrwtb/uRYCawalZYZCXARp8y8UgcT7jRi0StXzat1tjdnSKx3GsmZ
RmjcxnT1u290c8MH5REzLx11qkmMlDrPRv5Bg9sIMRLlextIed6Yq1/VncQSACpy
rP4tgx8cjHdS0KAx4JUiE881ZOtvQ8RVpTh1b8k+FGESKNwaAUdOe46jtAYW+74g
Ls37vR8HaJOGFMXY8JslDDlEzX9GDgP25sMUmpjp/mCImJFUIYJ3u4n/wtDzlmpk
JRO1pVG7oeiAyGZFUFr7K9xqwkiB5mOrniPc2xHMygO45Lfnz1uGqX+8xmM/QxXV
o+o5kpAMqJXcpngxfbWs5zH2oAQdxTw1jMz882e8masQXi7UiFdAku1seJqhZiU3
Jb9Eei/X3KyNEEc1Uef4dXg/wLBhRhvG4J/DN+xNaR7MDkrEpfUt2L4igsD8w9Cr
/IBMg5sP+ZGaSDUSH1sMRjH36RwG3IcxvQSfn7uBeX5lcKW046qET74+ckk0XfCD
OJlKcFdQ+tX+nQdcWdsnV/mOq+gXI5vxVbxk8Ys1B0yWCjhTv8odlNjkYkLrKqn8
g5peR+p570USFjvjhD9VE0GFI75l079Zs1TW/v37NtI1oHep3Sn5RJbYI1ExW+WU
Ett2Pq4gS4PtIL3xjIo5vHetzHEY1tMbYJv/SwaRk9E6if4xWDL98ngjxK7O8oIH
EMvEkJsmm+e8MZp3W75+8TqVdNmxSG4lyxas+FceTaLLItFox6QWSroGeC1jA3l6
1ZiaV2kyWCjHgykLnO3M7eankYIu3qazBjNPxSZfN9Hu1lbTqQpxmhGgHgtz2Ib0
Osu+u806zWHTshku1K1ouh7iU3TRuuQ8gxbQdF84WxtgqWxvjZK4mzOO20Rt3CxW
jI6lwuYf/NeC6Pm0L3t0ap1h/Lcmw4R3kgKCe+AcNf4bEcQ3WNFizVRO0RNikRr5
vlg9GsyRTaX146B9zjwysy7hLkcmH8wyR5JpzsMU3mbzpzcTAuuWbWnIq0R547iM
uy4NVgTAmktiUKcFNn1AFhTtXR/823RbzDQBPRVnCeD+/Pg7wvE+uUZ9QtObxSXB
dSUDFhR7UG+SaLB1UJpAIc+8d+gFsE+v453NoKjaZSnX/3qfsmHkPdWe7Y7Pscda
JqhJBxE3AyvS/8LSgII0prYt8rcRqQXtKoOA5YukiGNwM66SS8xugsJZe7PUqspt
gE8slFXqyqiKJbxkUpkRw8W9N/JO803MZ1sJIeoCsOrzxdSdZJdelcSy2ao4H+b/
pNKp+Zvs2jO2glLErl2yZFq7iprDIZ3yWGbXUNSSRUaUAZIP7kXRlZ1ZzQ7ZIKXp
5eVH9CkqLmQmkn5bXvz4dEfAhU8icR9RlGN+206+bxJ7rORakHauG+REy+PFUwgd
HM+SXSGZSqsdMVWikp66DDE6h9FuLOD6rZ4ArpwDF1lF6SI6905jbvlywJ5FNkUs
qOGc2O8YoBOCd/93Qt7rR+2AC0kT5rsVr7EBVP9GgTB7iGeGmLIvECmJktwS53FK
LXZb4S0GNoLKwPXbojvkfHCEDMUcAjS7wZ986W+GEkokuZYLAbzRj3VYQT+rdRbN
s+HSJ6ozseM+xPIlS1nWXQlJ7TuxUesT0CeMGgQuCCH1dx0SYG3IJhGMoyMWZpxc
/Mjz3Nlf63bBi6H7jk7ssa0JaHLXDNmQc8tESttsq9w3z6ygsvZ2gAF+rRExzAgf
X1RXe4Gt6fmq22sQIeemKVxLNja9DouzNksNXAPxLXOLXwMNWVHNNVvwybx9l3rH
hQImdPOd9yZ6cRMtIjpPIhPAabUQ0QQi2QBgQQIdiULqXezCPtSFcGI7crm1CvPo
DqYKmj1yIdcHVGTBl3gC98+1tcg9dWGFqJsCrSbLhhDsTWKgNRgGjCXUNTVq6ao1
7Grl5mGdagAJJ2vJhM9BzYC3GQpA7Fy3B7EiDghh9QmhH8vXocrePH6MwJNodw1f
FkIUcydlO1/+KRFa41sCjT4PXYKTfGHa3Mg3S+5I7T6du+3quXOf2gI2U/2vsx4Y
p8Fa1tgYRiSZo/tkQ8FrcoLjQhuzPYQn2R0q4koJ+dCaRfKt4yCiKmw75x8eeLKb
mKw8dWsPiq14agRONqrwZJt2ON1wOKNecSOwGXEkDXyA377rhDu1782xfTCbBIob
JTGflCrrpL1wfM2fw2u8FXpq071Sa3I/LTvFqmG+ruWtL+9lBZgwVpf/Sqq8TqqI
jNjPsHaHBzH0nJIUvBxjNH0OelsA+oTqbJ1Cef7hDic033GZjHUXlzkqryWigbqb
3nL5xLlptsWu+9jMy5UyQfDiutt/LWofJ/sTZUXAsS9FgNohIeSeycsQ3ocw0JMe
4odeoE+101bPb/NFqthrHs6t41Rn3MooGUvhyUx0qYcMt0j4CXqSM5Ry18Z3s45w
RbnGiHjhWA9T71l78ojE3W5vDrcmGfGXPQkppFvgxsghlu+9pKmEgY3d9v/mq9q7
rNI9z++t7+k+KHPqpWJHDkxz3m0A9TF99WWesMTdbdlR4C0En5q+CIAin/vFyM83
+eSFlzVXs+onr+aDnmM6CpnmynpWehHKlvzqSyZfs75QdXA2vkVeARsgG/sef3EG
dLzoNLewfqLOdBZQ4WSCbKkndIe1RJ1zoEO1d7W9eMecFwXEcrq0mE2J4q5+nmNg
TD20W2rCvFogmlZljg0J5wm+BsAm0oYP8p8WOAr96bEcaBcT7yh7emMOLs8GxptI
e+byZ3ns4hHpcDNBmjOPHJtTZJAzGNcYyKJSZeHAcREsOpJv4HPPO0xSnw7VK1b/
xM7laZRGy73Rg6zlpbw5l837ZeaQgPho0JY0ktPm+ppvEtyTEsPrYDWjVq/UX45h
7EgAaNxJFfm37/clX2QQwR739J7SVMWCGgNRc8kFFEELA9UXx9eVwZoRZ60S8oTM
Y95E6VCQWvN0q0Tlaj4aIa/o7LGWdpGItPTr5IFEpVCdJX5h0FEHzIEB4ijFdhZb
UVlWqXfKPE5eTDQzzhH2WMfqXx50mXRG8T2CokrxT2JXqJIESeM6WLqsvsaXZ/K/
fSQZl8l/WbG6G19YdOOMSSppPJ3gqrmbGtjGDuTZaK1z1YrkazzctSNQFWnrEg+A
aW3QM/ymEKDfYuKiuhCAxj/C810wok6/3L+BXkXtThtPXVKus5U6FQCeEK5bctF0
sQvTyTFiorsabQDJqQJkHtllcl0HQGVhbeqoBs3OKeN2uoQmort756sYvKFy5dkC
hqZXdDbxpoWFzohrTKcSqstCG9bzRtTHWuYi3x2OSVfLi+QKdZh8HLWgnFy2qAvC
//nrg6YtgHtxPVqYJM+OGh+XaBarfbw7BFCk9SinokjYiEfTHTSx2hEH1fy8Hdhd
xbQX/ebMJK6woswqZkGugvBxuW7+2thIjA+otDBcaV7MLD5D917FboHYRVfP3VS3
aZphoyHMvuvv52PdN78KRYF2Ogk9pMTQNn87TrbfPl1ixvkwDeSOXLux4pWh/6ke
3bhICSaip2jrAbfzGtjS/0bxxuoaerAa1uL0xbeRclaNPZ+b/TEydjSemRLotGtU
KoMRSQn2bVSMAOysdxaA5TerR9TuX4X512AadS6KOmHZXfpo8jLltck7CufyC4ce
8xnyPZpCagMoaQvPHrp5Ot6Iv4VyzLV0F6qF+uNx286rBOu07Ui8k/31uz1C1T49
luhJUbNHwYL5qK3kBVQRwinpOHCZTJ7XgXMUI9MCVvlKf2lh7X6jBDuaz5r3el3h
vNwFUgMPhDSxfIDUV3Z1qSRmVor9j7tameLeG32WW5ofLy4JKdckzOAN/xt+heXF
oK4dLKHWcT/z1PANdqGEeNeOjYmvKF4/3iG7+yizoo+ZfCgomsD0e0qzRB/ggi5X
9PbpdfSEWD5iO1v/iuLE4od5wjkRbrfU5lz76h6A5qTRooZOuxVcCveLSnlftbHX
x7qZVNXgRjxJxVCYp1kb60Jm+r7m1upELoE+oDv3PiYTe63ALGzyeGBS8M86P7eI
xpGMHiEoTUhoXHP90LQgQZvPL7DRYKK9w9mLk2oFV1PBCcMMewNExlybKPzf7Uel
LBWCFluqqvM+8TvSvHSd+w09nMxgmP/mycu1xHLCL+6JzH8IazV1+8p+wvgkZPIH
A6CxvXruZ/hps7IiGfJ/ZALSQmaxStIE3jlz1uBMbjaLPEZaOMacYU3BN6kvzEbB
BBiiqEKHLVXdZC5nhSreudck4Ypktei7WnE74YRg7V1q0ypVW/biN+Ci4HS5yjPK
wegbbk4Ko7ZQujJedmJtaPwnkUYY5urnRqz55BGxAOikqSBh9IlFhTcbFsBiXuE0
vxfjcq9CaVxMGaW13x3Qnf9F7LmQmbRMqjb+9oOozDjLG0FG8jP6jZ6gm/7tngxD
kC/UtIvcqg4VABy0U5OSX1lTNUznDufRtwH6cdJi8gvu5g0xVm+AnWu5TwMt8MNa
RcEURg9QRavxO1KTqbq1juHUClzhwIPJxwbOrYsSoyUlC+v8qVJAO+A9K3fL4E54
42xpMeMWO6uwpqMMpsZGBUcw/z1LNKfoTpSUCJMIXVbKwhqsrYacfyn7TQZMWwHi
d/pUxct1rOXjLmENYgOCxyZz+EIGiiqdW57+9QRMI5WE6EUXQ5lF9uc6LfcCpRUG
tx8VnjxdPrLaUsws/XUjseivfOikzWyiqWKor5x8FSR3Z/cnvozsbdz0rZO/O114
exkrPU1JzIeniClw+DG8Xbo5g+mC8UBy3FJ68pQg4z8sfl9KkMKKkVoYgEXe3Sit
+hG3UD/3lRxwGHyv5Rvl4jXT3L15sm/TFeRDIzxGcYygqqE6TEnEnQv5b07/AN5v
knD6bd6wl0f5Eea6EoqRQmT34c4Tez35trDGdDLB5CLf3q7rt2W101xeAe3679RT
tfUAPN9Be78n8RXvjinTtjo+tnraa3kygjqU4erfr4D/nTpJqeTGcIX7oEc0wq/g
yTfs9YasmoJ3yNj0ZYZJmkzN6bqyOz/Wp8/S7SUNvGETvPTEn+MozkbVauPcj1by
o13zjLuTr73v4wFxZVBLIDv1jK31Tj41N/7dlQ+Rd8viDQZifd5Ys9ZSy7xG47kp
VPLR76UCNMYvW3biyOhkK1882yX7jYvi3pWVRNiVXGPlUQsQ9tNl8IuTo4HYlGel
e/6M+BXTE01ocm9JVkpzGBsTwcikh9ccmIqVVEJcF1pW3zZdi6CwB+0jysCyjMZU
Y4NeB+BvrqVPiRiHUVpUAH0GYx9HIoD2FBStEbslFHJH8k4w9xhX/pjlmOUrCGnV
LuO5UPxlpE6bi9jmGTulVL7riOXv3/IyRggVpc4zoVlWbIW/uEJfc7rG0VUzRRO/
fItpIiDhZd+ZCdhN5rzJyI7xSkqjUlgCOhg9lE50Hb+rJOcLmn9sPyJGRE+Jz2Sj
3lhm3rrH4jJumStShv7yHDQcCZi1ADy4o4xCeN3vM0AgdiKZLF9FZxQhwvTOb4zt
vcMSxlp3kXgbgkgcV/memyDzPvoduEB6I4utwCNK/qHBTsYn2DWxJAsEpJ15x3+C
dcX170Y8ereiDkFMpNED7VSRamvLSABSv1+c1L8QMxhIvJ1SwxbcW8acvP68u7zO
QZZ8ijhM20MH+Tb2c6bes30PvRZMKpIA++WXO1gJTvMhHTqTvPWoHTxwLXmPxa8B
nhoNMuT4qJ2lowieJGLA1C9RwAca2ESDVpcKZR6ANegoePKj47UmYdfjBDlTDtHp
CjZM1pvlXX1IV2Cm5VSjACBPRxiaVxEfG5ATmHFMoBgNQeipteNJW7ZWRVruQnqF
JTay1U0ZDQ76lFdw347hww0pssByHFRwhvwxXy4ZFmWN9i8LbBdklWU4orKItDyA
rmDfezGIPis7K4ppQhV7ZY8sZuuC0/b99fxM1ttpU4dCr05v71smS3gN//Ke/dvV
OPl44XtyKcMovQqdA3h+PARr/8bSpywzGI8DQtpkwSRzue1hpExZFBSH5Mxsh9Tk
ExAHDewv4ChY4WOpxSRZUssryqvbafbBbAkAaYrdi/sjTouhraxXGiJ9ClGnVayn
+NWns2919gNPx8ez89i+rJDHH5keZka12KYshNNI5Py+GEA2iPjluKmAzEnpnQCF
yrwTM54VKkZToXMs+5guuKCQD6kHEEZxSJO+onuszRaoEJ0TQruxhU88T7f9ojA5
yDrTFUqQxhezEmqA8pezLsaSuon8R+Vq/Fe2POVk5b5UyDRiP6EH0yAkSp2MxEez
16sVXvpLJNf4KkZlliV1VW1OPZryGTlxTKXNUxJsvoD87eFMwstdJqvVzYQJx3zP
HC6lgXdggE9BL8rUelp79wl+MJuhNzgJA+zhk4e2W2nSqRpVYDl12lxuKDs3081j
Olq40oCYBfs6j617f50jCbzevwTuxwhpAYMpL28H59onOU1wr1LuCcbqgUUeVyPK
rPj3E/XluMJl1dhYezY02krueTgjmsv/0Js5JFsqTtd2mYDXqhSn2V6TbdFXnXwM
M1eYOpWwPDEF5850MlhgaqgX1RUnaOY4K5JfOlQSmHaumCsBsNl6LiRrP2JrDsWC
JmgO20MswjgMlEMge8BPjTIQGbXoiBvxJ2Bm1AcJURFMlRRah+AWjomMKqNH/5Ql
hQOMOAnmbGQ2OGcxgtyXGCCog9AKKwY7JcQLJ9TWx99wUCfgkQIs89QSGs/jWKm7
VTrkJa/1ej0DsBZ00yjasQgielttET+TR7mI544wotW5RI7qYy9/rOhfojbMUKwF
8s+mRWbnmc7q7zw6c2hTSn2JOuiLXky+3Agvj6/STJtvJxbASZ59VsSYtyXD+dLf
rGLd+RXHpRLdPlIbE9BoeTFxDIWScAZsfEeeuJfN52/k/xSG4vuma6oAkCHqOazq
h2XadaJqvMn2TIz99NX0FYgsjArNWFcIE+GjowkhNQgm4W5tODqQEcJUmb04pdYQ
Y51NDu99ZX9RXc6OzTUOtbUH+1G634F1/UD4mK9W5pMPAF1Kvq9z/J6fIiRByef6
SKrV5SVz3lSBXid7nA4oJoNXYOzNjtbbdG7zuu0AlNvhO8ZHXGJhFg9P8GbRF8OZ
UH9P0tiAKtxHycqdOks0Xoi7RsltBScW+fO1m/FikOby6taBjJHDe5oUMcJViQsQ
lzJZgmwIbX7xp5v6UoGOgpQbunBF4mjpv/GJKS7dqRUzzS/fkN9nL+vZmbV7J7hY
UkyJgG8ADDBbBp5TluRl+fCe1GRgK2FdH3TkctNL1kGlg1W4BM7mzez7ThZCXc+I
pRijeVQx+Eo74OTu0UMtPwZFmQRzCH9Rb8IEC+bSip9/KcxKPX9h9JczAOv8vKg3
+U/W3rytteRkuMSvC6HBduYx8HQzpwwJYPYV8X4U1h5RtvW7WN+QO56V8thOHUri
NSRSe45ySMLvCi/xtQso/bk5i+1AUasF9Sf6qmjPPM/TX3PYRva8NfImcg9nm8Op
MzvEY7wtOXg46tkQS1ZGpp5Rfev2PQZm4UAbhg4EEMUaWu+9B74RAIcnl/BH0FUQ
k0AakJi0RQqv8gNLHtgzrBo15dh6i2J0lRRBnlbQ64PJXf3fSK0r491dHMcSG/1c
a9bwtwOPF+esy0Xpwni9f7F1LEWK5pUimrGu1AW0jwibkrhcfDeonpz9YWK0BZt4
06Mv/MUXqP0CEBARWwLdwj1f/xcKCw69PlOIuH7EnVfzjXCtvBPOR4LGQEI5ekYZ
PpBl0Wwdmv5xuZow92NnKOwlMufIIDYWKMu3xLsdCs1joqQ3C/r+vqkxgbVitPtA
pUtJyEawJf+UZwONiAAlZ6r5X4g6TcoLdgToXaO+lOFu6lecH1WcXB3GgOVuyDAb
I9VEFdnr9TZgRPc0Woj5FH9r2ikAsQtDBnE+tepC9hnmhhag9awKXUnMZY7eKBMd
j8lKU5InFwb42K745bCVRRPmt51e+VINMwMz+0iuaSN/airQLHhNYz1Z+VS808uQ
PW81Ro+q9UCJzg/2DFAesgXMWmj7PmEPh8rLZ0aIvy21Cg17Rp73IOjJBTGB8ufj
i903a7FKPVbhwIEzdkZ3TUCkUVMNhekffxN+UE3Nv3KD1fpzrxXDzGOXl8grcDQt
RIzI9eBEBZ90/u5cCAGF9m1WN9bkrH7HeyYwCLwN6ivEE2JyEDku1EB+BVtqWy7D
iK+vZPH4sFDPwZ+42Sgxl2G8dE0hHeITv8Mx/1WCGsLSdOO/s1Z8FcJVzjgiN1zn
UKr2f+MlT7Jjy2evwJEwTCeNnRlG6iZzLivISALWPKXwOVRpZBFfu3oaOS3rsP/T
ObEr6W9r3LdG5WGIEpp8HYlLCOLirccVImxMUHlj4JvetHfZwUXC0c/8DGWba0bE
KVq0TD7cFQGNvK9K13W3JgsA282QR6aRa7HlHsaVJl339E6iVkSKI1EfPBnye/WH
QR5a2BoEkXIKrjS2XPxMewITn42MoaOeOka4m3dWPlKkJ5UFZR5tNiSoGq64Xsxd
OGZSi74LCECGjADzJVKzhxA9M3ZMKl5FXPxOgzaS0PSPbm4p7cuxAtMCnLR2OrZd
vPeUpkhWJEzx3fRZsv0p3+KOge48Lnh1XWNqoh8YNTiGb86Qgefs38cN3FF0iMVr
H5jZmGYa5jHs9tia/KhIUIPpjXs2uG21vNyv335fRz4AA4OUSrTj8zCsKyKvmjyi
zLV+5nJtfLNiO64BOzyB2EYZ6CZV07kLvbMA0ywTIwqL63qDcEnI30+oqbTGbfU7
Md9Rxo56kOHbLfD0372YqZaJoz9T+wE6ChtTTDZoyKuqE2AtPL5UUF05befFfyfv
kn8ylcAl6rq8DMBGEfc2+6ThJlWQ9FI3+WIzNxXk7p/xm3DDYL4kc74Pg+QLS3Fu
+2rb9p5Bi5Xt5Z+KfXVv5hNJDB6+o5MtqpNZuHHf5NnDSNqrExasY4Zn3snPpX/a
lkk+6Ihu93YMAbJmb0iJiDSLmqr1qeJ8jZ3XVd6VnS2H0yESZ3Y7vWTu3tsieIlz
rGW+Qvb5CvIf9KdQF00Qb1d/4C80K1LqwG/9Jox98Qb5k4iDSClKl80cObESUUyT
ZsezVz2HeJzJyoPWMK8D7V5daDfMul0qYEC2+6y9Zk+e3tw/CA2iH6VU2EUsBE3m
xSQ6uhpa6N1I8A4oO92UsAd5YkINpKpAZ1bF3FTtB7Fept0c+rM+6gkmeOQ6DPzB
rd21nUtx77jNT+Exwt3MqAeSlu8AAy8ud60HuK3Jchr1QkrLZFqiVZFNlkB+6txB
rk2+9jVJfSFSrDmbe0YZbGCNsK1+YnpdWtGcWg9DysFomT36KFaMWvLtt7eJySRg
etJUKw8nfmJGm+oh/WS9uNBeOtl+HnhJCO1NoJhyYiUxnJbJf2klVDE6Ii5GZPVD
NY2GtV8u/KefU19JYt9qJqHT8eTzkv+2RSBXrakKtkQGAZG6F5u/pXF7JryGiu7h
nCMmRQHPDd5ztgd0iNm3w+9iwuDxVAwT0GdrwrRwjnNo5euDo9SNMnQoajo4rORE
hzATnJFZ5eDvIBSA3ZJOhN0OGI0lzTd7Faw5L8SrjEM/91sZW/llouU4K2iFALCv
WcaUZ5qLikacIAGG4zNDVgevH7rlcaGfwIwdQ6wHKg28JnqfRiew/WC/rlE8oWjM
MYKC7e7v/UQo71Lh0lSOpblUUniBd+B4IYjrAxQsFbmiqOjJyJnh0ZRzPDrNDH4w
uCm7Znn62sOZcAUm8pOgKBvyhRH3J/BSBHhoGYb95hOjcKu6kgUczEUvCrdYSsz/
OkYoQ3/KSZE2XfLy9Sg8w0tnODwAkKQzzBI2se0rGey4Lfw8OZ8sWg3+LLRuTzlM
zFIHnZpqltGPMNdJ0qa4IOI45cILDFPy8JRU/O4MFY8gtTgl7+UvgPfE6wRTqBff
k1FqbI2FgcU8XY9t2zEzprXIsoCXcRbkFVbDRYSpykFgQYgPLKQzB3qKavEo++Lw
NpT2ATdzS5VRtuzvvJOQTvcOpLdDkrCHDzVCQuDIqLUSsaVdqcFEVHGMZwSMLCs+
xZ6L6eh008pLqbfskhkYVwhercS5M19zHaa/4I0B847sIZuuy3J11Sw2ulRNz4jY
YuyJRXxWyhHpcHxFEBaUYJsVkWeHdwyj0118OAemwDvlA2mDK3TObiot9jzj9gRq
QAZxoWWR0OL4ORSxYYEzHK6/lzjc3tfXXZOYcQutsFAp7X2FrmH/fpGrcIXVe9p1
GD63kWnoe/NeGqm6Usp/mQOfNNhkxeYKNr8JgqDtT2KACHt9kpXLebcwdd1KuRin
LBPnflna0rdMJpXFa1G/XYN1B+pfSCxaxE4S0BfE3ZFW6rmAW49XQ8dfc0T3TV5C
7HW7aPP0ed5oD4g8rHvSiA9mv6UutnsvdkYrNmBF8QoTG5LfFOe+Bu8Qr0v99i8H
xncnCNaixHp00ivCTr1h70TDPd+XSQ+rb4jvbmBH87d2L7YpxqVHEFwQk51yO+69
Q5ECvI/RfM6cdGhWjYYgp8GGqzhL/lnQfFXoCA0IXj5X4XTThpxHVFSDsUq/J5JX
PXS/Iw2EXap1DtpEAkCZ97ZPDrooOADAwUIoTH2RAPFmfjbvdUxANGk0+FjYvrcv
PpNsq6RziEBXL6q4sB0E4sdpzhDTn4EvGIB9n3Q5s3cNPgvXlLo3oi1okXt/LO69
YMXr7pkoz/FqqXUNuSal0S1pkeNabXfxHqCfkh14SQEC/4abVSDC5KCR0Zi8EFko
feU3YLkBQLeFTOWgY7nJdxqQC7ICgWWDB1eaOPRVwAmjeonRhaUccjHKg4X1jAlB
sS1VesdVooz1+pKujUnBivwZugskCQ1ElqQJy0Pt+OA85Z60ekBosRRj/ofSSiA9
6AYy+Zt3z0DgBlOy/R+DeXeoXuSjs5zol7uBURcAUV1phgXXQq5i4fitoIILBOfR
1e5yGT8Bp8XCnBy1IBVXerZiGwQLatzHQXVHmrFcdkSlPootrOZ755Uk7YG4YtHG
fRuFOdq5KtY+8S1bd/TAyegOdaDH8v+cRd60c9RWo+1SdJ5OQl+22bWkGMUMllCA
Vrmk48AE397F72LaW/0LO1hUvprvP338iBcjG+AGNxNb/oiH8zY9PSwMkYi59UVh
jOnBTNzCls2BIEXA4a5qpS4Tt9MCfVuzukrvVhqGpbjk6eqKgvrs3A4pdE3cOmPm
WwpEWa7oZGsY0cXWspXkUOrDUp19MyPaegZDCvWPZKa0U94DJ9A3DGCb+PrwBiIU
04BDEE4PzUm5HEDyslr/ia80rEcae5NHH5BnIhqlO+6Ixt49UOOXLNcgfmJNSU9l
jEwRDkXLc7MpET2qkAt4PeaPDeqtktaNT+/5GiT1iYzvqEpK4I4WnONlfiGitTXL
1P8zYKd0G3whhlTooBr93xwblkfxihglLLsEqVCs2pJF3fYlfVdg245TtIVxT8Dl
fmFy7+9ScnFGui62o4c6ps4cL6AvHPlY5JHUELnrgc+1fG+VaM8557BOdHtBwciH
/mQ9/8spOM04I0/lYzCCxFPMcM9IvXe6QYyMsfX5iTY2bLNnoOI15YYkgFV54g4G
UOCQG2/v7YTBI/38elYFKx8l752MyC7LW1d6tkhQgGkdmsiL5P25yucCTx1z+V1J
E8O68DMQr7E9FvQb9ANMRvUAqxpNIJYPAkQhpN8T9k0Zvk5pczgvNgWQ4DyRiC1Y
sFGJCfMRG/ep3Ez5nCvLmSuaGuAaT9VE4Os4vER1zrHGN7Lx8c4nwKQOzsakrgn/
bfWb1K2owt2M75PRpiC36PSCIEMRN9ZNOi+59+3rluGGDWpG9AGCNueqVTBzmb2x
BDCcQiIVTPKTSSlYSNmZRGSlxKM+WZDA3muAhcBr/cbYadsqIJw3/wtrgOQ+/bWB
zc4jFoPus4Xo9Gay8t9yN2pztiCzRahN3JC7a74KbGkpnN7+QSYSTEwBOgNi2XQO
P2XWO6GNJ6DnvnXx2LQB1aH87hfWqKIdm5z9huFsZoDugZVsn7i+kJExC1Sdb/Ra
Y9pCv0CcEyok1yeP17It+c+RDPe74yONU165nQYO3k4xm4ttIM6LmQYIs1rYwpCL
MzcOvTJO2hs/+BCeE6JCdzlhK9nFgUNk1Nq8w/W5AVQYh3KzFlA1WOxm01zwQQD3
RoiFbdQHi66nPnqxIKLk8dAOwLZT40fNJZQvf2KI1J7sWq7MIVzVFM/1ci1nu5qy
s653Jx4yYSyJS6rLYtUJ8JoLNiDm9KJNCx612SKYXRTuW5MHcDnkxVJeH83IFy0f
XRI+FFQXDHo0La1WCu5LBop7oylL8X68n2e8Co0j0CEM98RV/rjpQEGoIQb9M4cD
6tm0FcuSWThKWp4/51IwpWNNeP97wuwcRlGOk9Ct5vNuPIglsgHpOBeou/hEgz7x
Tdqu/Uxe9/fh534/Q+1wKTej3nSFyrDpFk8a3fIDZKugPZTQQ+wBhv2M9Ro6TRDG
UMv76fKzKRr9GUACZltMGWSG8iTjXyFIonr5FuR4lyOBwaNpgleeNbSbGA64RkHI
0k74qQU8V8OS5v7mHL/NNbwqi5yltrqHn0SonU1asB36tZAeM+3atXlP1au5cLC6
OmzF8ke19QJqOyRlXmpof65znbmBAF/WeSQBLUv8STE9Er52B/g0fcerhtrryHk1
xY7Iox8Mjaekhw3c+4LYGZp4fmCRP60nawslnaxb4Z6lnBmeffuiioEIzGUlnrkt
fT/LEvkSOfuDbJmEGIbVC+/H7UAKYGi+2D0U2ohZJ2ddwr7IABkuaYveguP6AK32
NgZhhyzO6El+vWVtgBjOWEq8gkxn7+2X04iIt88Ecv/rDxk7DLmWslz4O4AYlTTx
9nzP4QA78Ky+4Fet1lqux85Vh/LK0JIEZtrYdvW47Po82ScLWkNusj4TvMd7i0UW
DXkH/h3hJdKb8zxtMyUHoTVwtgfOgYkVST1EHz3x4ApctYRokbmbwLUGDbvS3tS6
Uupy+ZjK9Na8tNqhAPPXwoyu5rTjiKSGPvUVKN12O5oxvfnWY+A/TRhTpSdwSR3L
HcQEggAJ3+ZPgKP6TM9HlSoulbqjdf2uy6AQGqw74QEC/A73bIHhI3wW6Ya405k0
PTgl/19JlvinO7ltIr/esSROedhmmsnrV2ENy6i9HKjysV4ZXrnu8xdtxbm0o2XK
INGbCWPL7GqY8UezhD6knK4kVOwJQ7GGJrRnEv7uTIl/KfUqhHkmsDvu1abV5jCQ
5wpodgiHcYtm4aS3LMg3kiU6W8Vdww8ABSKYHHy3+Lwntdqb48CktOe4Rd2i71/I
+9NEtBWlGVRWXAVHwR6MeYmEg124ROhumbR+ZuEU+h66ZElQqkrtQWA6qzhJiwO2
8Ab/8zGApPVBjDIr5946r+mhx3rc0N0FDa7NjnlTVR+AqHo1wNSuVP7s7rk6GgWa
oNoAacO1osw0y4fRhCq6rTJ9OTSxdqON1TjP95mrP+VJXO9/Uh1zJCE3wUSKdsiW
v7wcEdVItqv7cmLksG8azxG60ONpxXcTOqVpg+txmSHfs0o5rK2Tz5blP0zSgwj/
LD9fA6Fwqsou2IF+0DiJw/7gKvDXeyJ1j8oOTHt5LphD4q5YQOvWfhDbZkBe8Itl
gm2D7gEfscFmodMCnmm58D4bB/j8zDcOL5KvDtja0+r5esprYERVBRIu5V7pKTg3
cYc4l+lfHc6uyEJuQhpWXOS7X9aEQMcpymfj3g2cVbc9BYaYUc7DdIlNfOePshg+
no+y+Oh9slAqfi2eNK7DGeryD2s24rBNOIvqTHQaVPb4s0rDkIST3s7A87pKzuW6
FeGAy5I8uQrzCVud+TCRy77kP56YBGHkdSK2QLWOgT4LzKcwnQygJmMPh4a95Wep
t78o03QF+on4nRitX50OfmueljI2wYJAGWGoiooWe+7DYF2FXdUr8U/xonslYUSE
fm3tOc1xInYKigCeKE9jFBcxw6ynpg5C4/uPRuCwHu/25QXz3fS5RuXV/KW7n5Jw
IvoXnqbIo6m8bU8tc/r0yJbO0exJdf1jrskhTl8T5qZUFjuePBH+4nwFDYy/BGgn
6X+Lu/hNy956p/mFqi4JloQWaoPlYwyJhOD1cDwlwI10naK1IQvaeHgCJR81RA/l
Ej2xmEelzxxtSFzpMnhXDAKQJU5c+fgw2hK32/WBX6VcsUNk80TS8+fsFJ5Omez0
n9/Eg3tnFcgS/GA5E0OBfLh1WtyycNbGAl9R0cG/V9ciM5vlTkO1o+WWSmdtwUgV
nUu/nuBZms5zwqGjwYDS9C6IsSglVzBb5CKNiXzdtvuOPN1oIiDcjGPJBTf9s79U
mcrVfPjOpL+hj82FGjhGxVI1iuADgwSio16H1yd4jZXA6kaGLicMwH3uDmbUJGO4
JM6JoyOmX6pwlTIRnAzgWEOlabMEMCOREvvoYaDC//7MD87seNvg5Lyq4NaRiYRJ
PFwRfClaeKKzDSwjgH4YVB+im/X/NaD25p+LtaFz+n3OEfhDxu226eK61CZAeHr7
JGIqnkPK1bbm+SYKr+rKLHS0sCpxke8yeJdBQfeH/bF6iTNF4OYt1KYXG8RJZC3K
uKOlYH52Rl7lXv2VOmvv3ETRfFrCnDb16cE8uM6NHDwyOjJbstddvEPBA61iEcdo
0DpOQLlyb4N+kVLCzPMYv5kmVTXO8D/xk5hgOC2dCWhLZqhMW8YkHThrZqKOM+L7
beJhvPxWitw33BqgqQk9DkvzWC+pxDNmS1dD34IM8U7meykvoQNFlvQ2OJCly2Qe
TTB2aMhygmHqNjUgecPTbxtgJ+0Gxl96u4vwOFr6c2cllEc2LGQJ0W44kD8Ld1dO
azMe3GoThepPr3H+wBYz59QbS8juC3UQbqosTustKOg4cQi/2DgXGiOZsjkxEUR2
lLNX/aUxU9pvU85OcGC4jCpwUBQMx7sNB3sigdOlCam3s9XqMb4UArYfzBt6owzP
jkO+nAwzKvIVz2irHvC7JQD83ufR+p0XIZw5xajmr6bKx2X7gFu5+q62dsGWFFWo
d92WEpbakHa3EQMfFytwrF4hWddsELsYUP6oweB0QBUtwuZuXIhaICVMItLbqVza
gvaZlmaiZisAbLtfn5Ah4dWuCkEIqB4tfKrnBjWxf1hovgAmlfDiW8L2q8spsArA
sS+20zE/jPU8OdSTuxtH82lQFfDlcbCSehzWzfyAsPMeDA66+DqeF+P+g2RqXnDA
5SihKwPiXHUwYYcsn0Xaauqy27ThiUh95kAVzMTbr4UImekHhdshJb3hwEGX5t31
JsVLppqF+wTkbeqOdXcjCnDdKMgIJ9/IOFJAYG1SMmse/5wJ5KIEpqCNrFq6fq+A
lubYU6HLtcQZoYbmGImCJjX0NWTspBmscWZAWIfKlBWVd+yoG1zShIBlKUn5jS8y
10JrxE8ypCM11XwSxPLQvVeDtzTEK173ZmsMOuUqpIi785ichXZI55gsD7HF4evf
cq5spvW0kwyTNwZXD9lo4izFVBFDtEbhvNqtjXZ6YSb7G+RXFB4VYxtbWaIoThnC
GOT6Jhx9Mi9oLkYieBinTW7pmAad+hYYd5xX6pFhCpDvCSW8YUsDhMkiNX85HsDv
sF7YxpVg8Dd9gCj2EKyZJwIrVym42MB1j+eA7d2CaTHK8TaTWi3ytA/aVhfHCIWz
Do9YvWznqg4D3KaMQz7Z8Mom/ETXLT3ZqVutWmHCXmyGG6vc7haWlpG5ULuaqQd1
MGFXZiku9pSHjgSmoIvX39fjUDQYBbIiNIVgDRbT05BphMLU23boLpiGLQplQvza
k+tqgvko2D+YnInw/pwJewcoUrehQg02FbsBtYfZYC3O9PzyD3K4YBcf7oRdJ50o
GUc120Te2p9RaIFtqNVPoMMo0OFMrmx5GW4Dmewss12F/bQaUZ3aFtv7at8ZgCAW
sghk/QgJEy6hDb4fEMrW00VwKe68CYwxkC4xswjFpu8TjM8kHPv9vacCslXtwWgK
W3bl2WhJo62xGJEptopvzNbx/GzoT3owA10FLjYenzlOFiyNqG0lUUCsVLaASCmB
pEPXyuF0e/R2Eci7yrXr6oSqISQ9Lh4CB8BCNvepLtpHHdL3idarSprBViCoC6PZ
yuUSTYbrK5y0vsR5KINJ5+s5Vrc4HF3Pt+fftKmZj7LtliKM6DO7FpqvoZE/RQBI
NFbL8p2YRtHHyUaEfWkq3e8aOJx4DQ97k3W3RoFg9yqmMjjQO+wiGNN0WZHb6jR9
Tk4CfCHEYjI/h8iFqPluqr8i8fAWHIJ6h9b9unxnw1732vI1/Se7ZOkfgUFxPiCQ
Cu8zQhocPILCDY2VZh0FSMKBbZND2+D/odyhlz2cXzzBrOg1BIoESP874x8PCvNd
RckiXV1qN51+g73/E4uYJ2QKKQOcuydXm+aTQn0jhrjxXCAg6TWTFAB0ZeuPWh+c
Y4OPMIqMjcty3rt2nbB+alZeGjdIogJiXKrxb9H2u4qK6SuqjLA4wKVUh+BGmXfI
x0vzNu0vYoG5NBDeqZSIE8Ck2Z/KA+aMTIgGWmKaIBTD87Dmja6FCffYLbz1VZQ7
x92BqnWikfgUwVOyOREfmNMn0gWiTMfu2VX+r1OwG7RYP3Q5s4u68nKnyfwjkMIj
KhLpOSOU+ZjwKw3dpIFjjtUsr5MYrhUOXt6igoNknoTSIPNgkckDyzthHrXxJpZL
7L+a2rXMRw3hf5M4Kj0DGXpM+nOFo/+wmzEV8QCn1iE6ZCSf4ezS+V633l0d8IDQ
TNZlm8HBwfx84eUf/WkoGZa4hlg5yiRc56JD7mj6dryIrVU0xbRKBaIbF4s7flpV
FrDvDPbf9WOpWFJULnafI5TxUhIe82riTTLIactBdYJecPnP5Fxe7lTsKjKhDtx9
IIH8dkFfhHdw0MpV1tKSllyWzu6P9SqKM6udYNu6Tf4rf+GPKdH0XjOvhWxnnVLC
Y4SKZa167zvFwtNSBRCkHw1CnBbDvOLfRlPSK8MNymnGCG9SSvx0rOCD8QzoqAd/
opKmshmvuZGrknMHNVrvxXVtRBOXi8teyyDVlf1eNQ8NOE3o/E37l8JyetdK2Po/
4n/yB69lxLBB1aJGlPUBSFFT7esXcKusgbr3npHiw1UaphvA6wkTrR3UF5PHrLaS
d9pgJmOQ69PiCMO18JCAzYbuPuXqaxXEgs8lkw1/OI11sUyv3OvkDve3mFj1Nnqd
Ry340D16nvgLyNMPSrdYpaWGVibBb8wFNoMhrIeW2bxsHA+aGYEEyh+68J0HwpMB
Uvyvvjq0/nIhPnMbisZdUhQfqGg2da8s3RC4CA3n+Bo+BHziZstb+bcERWonaZUh
T04Cxb1Ibr0+VNzBK/S8YytKUj+seXpQmwAH7YwLYInim7T/BPRygmji5tsqMVVo
rvbs7eSgyqDQAnG/TT1TzFAQVPx1J28m+JbX2rNPRPflmjsvFGmxNZvb2Svp98Pe
xlKTpep8FwGzNd+eQJUWUIQ0bYrGMxjAIWtIcamhKnsB9GhsDDzq0z4KBSGVxkb4
AjHfecnL5BQtuS0USTvAbHx7zUXtoLEouIZDklJmZNMnPm0Foy9CQj6NVu0sidNP
Daw5L9nJb41Rv9otYyeAU57jvGHJYzMeXZLFbxAvGZxNAww7NSv4iUyFbUcJptFD
dr+j09C3GzIAeq7AuQ9plaiQsYjLnLqeFr4Ltgff0sXsrlQuvJwp+b17U9C8cIvz
4UG6rJSVKPHmNJAHo9+ryKwVs277KGtz99xnr48IzQeATfR6RD/nz6vm3OwfAwSr
LIkyInOncVSAaefGx7Ocdvo7OXSYyXp8E5g3bCKMbiXgU6tse23p5BdUzehvdfPP
5bTGAZZmmMY8NQag0MpDlsAD1LDzQpwNl9S3Ujkom2gW8a/1IdpP1MKcdYSnV/Xo
Brss/5CJumUqkPAvWGBzB21CvZcXXd1lWWOF7gKPe47fZjRJirWRiD3Z6/jwCwbU
3dqST/ZXILr3BtOkmqvuMB+iOj3UyJwS5+E0eAkksiknw91Dcc82WKiJ4pN2rwKf
0+xwGEic6GBbmyoHpkl6m7FKteV6l0hDaDqDtMkTcQXraPAYsZRwEmR3cThQrWXL
KqTlr+0gmdhx/gv/FwSAbVyfJWOr2+WfSdWIi/yMrm+mJPpx0kvrBVGPXpmpk8mk
NXAObbReyfbYth+YeVwzAFVMZc1D51MLE0CTR66pvf0rL+jzZ3Z56kcmCPJzGPYq
aahLmBqM+AQ0HQem/tn87X2mzqu7GFVvOUnu6EscftdYgQFD60N49eg6+dpANk54
hYJ3tNocGxc1yul+hsXvUohM/ns4dJgkxcO6Mrc1p30PMvo6oqloLJrrOz6ldEgd
z1JGUOe23YI6vdMAm3IDuknHvpm8fjuB3Lfs2o/DRcyPeCqVZraXkSkI/CbyCkq0
/cmqzC3eoKCR+VFjZ6F4F94Y8DXRnFKNAIAF3IYCMiOoE3bjODzTz6s5jt5HHhB4
0TV8DUFqIQ0q71wmH4ZQMJHsB1hXhvJ5kFCcOA1p/vG1cS6xATl9y0l7vtFyjfx7
HypKPA1UquHyZlL7ZWv7i8QgHYSZneOXnplkblk1ji6mVFJ9NL3DHAk0oMJp5fWR
6OBF955bfNgKqSA3ayabSG8ygZhzapty2VSmc8dxLerfRKtXBS9H/mHRtwHgRsGo
5xa/1gC/h6/LzRFiC6LLXGoRzAwN+Htx8itrfS/8eOZm5USyA5Fk6nJa68RtjNRZ
fDIvl2iQXPKofEWGBqyeoqhTF/bBdJ7xqTAn0/+ZAIqny9CHxT46BMIiCXgY/v9u
jfwoLPKZJpNKzYuyvqcYGh9ASw99SN9o0XQMh/tzIkRDxFsaGlr17cD7vXTGDJ5v
W28bad+ZtEw2t/p0TmY0iDiyE4PsFM5rHd3qgIYEO3CYXaEpFx6tTs/w2XufGKQ1
OofuLGSbpuNCN3WWhQMGSHTxgTMypIH4CpOCQCYGjjgI5paEjdHTZYHcoAEF6LAl
0cY2hyWhKeR3/AEx7fWIt6xwT5A2dTv4tSptOij6mmGfIck6XMC72uxXzDRGwO1G
a91eK11lT7QNkzvSnnGJvviEMthz9TaIccTWP64Fp0ukPFY8c2XM0mW973AnPvaS
LAbKxm7sJIIV1WnO5dWuRpts38vn1sxjdYWQ+6EWk/DJgzzHXtSMeMUgTd0iC0YY
H9K38yY8f0kadgiIIy1J0ZnjJDHoiJ0aQmSVj+GfBk5hBHlIi9H/SCvSSRvxzq9N
hyvkC2YglKFtDP/o5vc+REkepLq1Z33/FVJFngF6r6jlG5dC8MjZvvu0AoSpH4HD
OS4wi//53+vuzArCWrgKiwPfGFCl9WMFWyPGb8Hvj+M/mQ/zq0QXTtABcaGoPCm0
mIXzMTHg2bOFYFFJLxNQmbdFVgpngKwT+6H0NxkTQpt7GwYBMu2baahq1oHEVi8S
zq7rQNorObqiFaRw0dIpD9Q5LcTJTVaXya2O0xt0S0c4b1a26qNz2FSm0hTPLHqu
yOjIeU8BXlTnoHkZK4lGA/UanV0CprzoqPUciysh8vbLWZV1WnGnTe4bpQ1WHUev
0WBqwHBPOjgjpgB0l4EMK3UOYl7I9wSu9Nr2rN0+ej7qLxB1TfV4vwybfAjbE1H0
l6TWGmMOe11BZnwnR7TlISNiKuKmF9SLkJZwbVZNfK6pShOtPHY5qF090S5jtdyN
bPCv7siw+GO1Q6VDopV9qwv7GEtcrr77cC0xbWTqwuUlqjCcr2e3pUa5n18XfBVV
4JEDxDU4jOzwuOVs+yzEQPPF/SeAsrJCQC5NX4FhLYuGt4aDUj69ZS9ZaPl9g9BD
zC9HLhWZiOVK8ZMnY+ygdBrsLpmSZgEpLcB7at6jtOQt4kirP024gx+D+qRisGLu
e8oEW+B4jEqlf9JazwDox1yXhaQVtMKFionBYepP5UxOZROzyS+KbVnXdXHrd4hp
5YCdrYmu9UzW9h4fzJ516h8HIPCIzwi7Lj7M5lgXXQnBWkwY6u+uiu0tXht01dNE
EmB+93VNXO4yipXSKi23YB9O0P36dK0deTSWSlhptfDHzksMH5rAjfPZBMLfrW8g
T4mfalVcG804mXuTKhnQdYEJej6pJbRgiFgFtqU0/besut7vuuWriQQNf6tiLHE5
a1Se2+pZLYGKKJ2BWMDyBQPrcRVFi+04dixAzQnxXpVrZ+YtjpcA09CqoPHimAxs
aw19M8ye7ClBbAvSSevxrDv7G8JLkJEQhkJrV66Zh/v+VGrewbM2KTNrcpyDnSRh
NO33IjTifdXgPdXSEa1AQFR3CkEaK/K+W3dt0ZILse1uur2KeJ87Cstjb9VxEn85
MtUC3eNy+6GGvWgveymhMP27rY3cYAYnK8ZZH46IJBXgNim04AnXjy1lkLWyvtU2
dZwSmQCUPcHO57AV0Xn0/BNnseT/BYDJaYasRmEcCkUVbPOfELr5Kks5kd5K5p8a
YdXVHiIMbIdPOjkOQRAfrvBqQlwEXh2xkbQIdBLYvUN3QjAcPRo7G5qgi6K4lxtA
ykr3lVyzZFt5ZYzSWPz97tnNB7ZDFlirV65alFmq7qEYgAuoKyQzXuEQTXu9qVKc
X91brh9dWWfKkPK6Fczzxrh1xdQHoHxnoKmFtbOdLcqQYIccJTCTYIhhaM/jsiDO
yfrXxD6QjlWq6fDzkjFqHYkNLyV0FAKyykIsKCBFtHRj4fo19Cr8OnPyZFcsyV43
6SLY4PXrZS92K4zwLJXpGKJTBCGk94HwLleESKXMihvn8vji2D5luek8STh5DBhK
be5eBDonWQtvQO2AjSu21KV9bgifl02oVlThkNmG7RYu96RC3CFPoHGUC/XynBCZ
L08rWXejlUe34Q0nbtsQrFyqdwfPZI/ACfXAvd0LdFxFAjrF+wRimx4L1bJPL6vi
wZHMxcGNH8/jvMEyZzvAiBlzrJe7iJD5awD9np7LinXSh7qhE29iHsnEuFjlZmJx
UzlhIXzLhIlmJg6ZgPPhMbH2AnxDzzWQCByTWujjCjhnrS0JqHPhxJyRuyICepwQ
iustcuS1K3FCXll/y5eVtxmWw6jdHntcL2UDDRIEgFaWl0xm26GTv35u+vBODpUs
QBIlw+IpL0+5eaI3jHyJYMagYSx1LGPMumEAa5pQgp/6zahTfqllIzEgykKA7i9Z
XVMB5utjl1yChYSQizWAP1ep0yfsfFwJDai9qQe/kvZQDj7w9FJZ0+FHoZODseYv
btjYuP+pV1bGjq8Ios4jrU5mKSfeVVGAwnslnQNbusbTOoJqbB3ofNavMFIZVnMs
skZtnO1d2LiTecygBe+hUCeea7sjMfC9SWwAv/mdXHahUjlVh/7wKeA+aJJAz7wS
qyhZNaSNeEKafZT4rpjzU9JWrFc56NsG5EJJFAoyECUQ7FfnGNusdZF3pnwaoQUw
JJaQ59W2Wk5Yd3AR5G5Z2H68uVlrFpe4dHItIsQy72oKvPzsbBZfTidbtZXw4JiC
1AtGTbgnQSlVtMmeGcI9rDI6sIbCpTBWUWWBIvC/EllPpGgLGu7A1fqcGBlxrOxv
JxqscedKg6v/8a3esZxfsqrsjOEok2hL/sJt8pbxfNzTTpU8q4jMmUljvATQtefe
LNcSButUAWxBSBTBVXWOPki3XtkYqxg6btskp2L5FJ42NmD9cnRYkKtrROFL6cHJ
PWjZhPOB2w3tB/vH4Hp5atxpxY79CP84q8dKmwf+MQtCFKGXnI9sGlfoUKFaM7Vz
T2E1KEhZKmojnt2cgplMHncmUwbnjBKGPXMP3rdz27fS6TXAAaQkf6Mcsc2mVZ4d
T53eMOjUrGWWFwFuL/FvDYS19KtJZFDkjLcW3locMvAPh4WKr5mQxZYdYXVPzmwb
ir39DksjGdw7EmZRkR9Ms0GetRIh3h+cbK74cyvUf7RBoxnoDLooIZEQ3ovMuS8V
JVBr+tYndspyiex9rnUVL7vyNOB+jr3snQq4qXXJBWmWX/+vZpU50++j1zJKTct0
4/AlA+PqJCdUIppRGvyZwMCNSsoIa+H3GDShXMcKKFQpJaLvsMzgLx4NTgn6qfin
WBcWa4uf3oIsE/JvgCqlZSho+YJy8PbiKh8buRCz1YAvKZ6TxEMzd2w6lRYCcUYr
Br5XC5q4vjKQQVAaYcODkw+RRztjFwRJUf6GeQOPyJRG6e2YJ7EJmATmi/7RfMn/
a1wZunV00Ihbm9UbHGJIncwdkn36q4gH/4Q+ne64+ErQQspB07LAzPYEB365DUAf
5olNWsPPB9o/tsOrlGfxqy2+KCGE2IeQbqy1aFZxKts+MAX+2iXycxcYSrXR7iH0
WCimQvopRN5nG30sYnyYZDuZKPwggkQ01js9ouy/X6zwl+QwC4Qf+FC58c0x26RI
QykopGBmjY/qYLm2Y+op7ItfR5Z94xxLFTRAqUBNYY4PQfR89DZXeLK5b57hdSZ1
BmfO+0eRJHb0+52d1xW0Bmdz7knJ83wFopn4tqmLhbjrdwy+hnqGwsqP8o+8X/vX
SLgJk51nZAMHZi1dAsQ8gugkdvXy2rK1yR3yhInEIDSrnV6Fc/H988BMsv02p81Z
ySDaxgPkst0COZSBkGycQJcqL1BSBIeKSmOJcFkLWnwAuaebTr3u4HE5P7MKjWRM
bPO21crp2BePEicIjaXYehvv+J9dUz7NfnOqy3J6waQ6fGkcKThPQK33cfvbInWi
TCG8kUa0QOio9nvcgVRmO0Liti+pPWb+5d8X0kMDBfhi4W3eBg/JGTb/SIQpNngT
/q+D3ej32rdlQ6Fx1+RjIif2VScb8LXzMDESNx8vzPwVLX9Ilugj834bA67ZqHyf
dYkU3o34lblmCdBBd62jBXycRwfSyndSzAeiI2Hr27nRjZzoCxG0p35g6eeeiFMR
0Lep38Ae3qHuA5Th3UgMZHror2N1ktzPSS50L3icH+0fPfb23eI1xfzBl+fIuXFU
H7h5DE63zHMfIaNsOniHQC98kUNKHkjKJIjePeUZ0E0atoTtrN5T2am+UMDnLZae
kaIfK+l8tv2Zu72W3KhpEgrXEOATM46sonHrpoEG2npozlEMqsYgJinUSP8oJexu
HWFh9Cdi3YxpERP2EEcZisVBqcyOZiZAiKB7jvDH7t4VC2s+b5J/WP/sf6neq3f0
udBBhN2zKxBRYwtp3yi+qPTSqbd/qpfDOZawM48fvoOb7Tk8bITkaoTzB+UPG25+
kRwXj2RcG6eI0U2UkyEyOxV4swUATV2erIArVF9QrKXzbfdE9KZO1NzmKtu7ZZtT
xhDx2W9n+OOYR95K4qZ500sOI+pKUGOj4BtGIFlauxYRS5zPNMZoikpiAM5g0ppt
UZZPLFzrgvUlYjwTOhQUHAZhFd1v+w/pk1T+yQUc4au7eH/PdcDxMOA5EMI8y5eH
8peXKpuIwod9Nvp3+I2TMp1sHheRtVs2SoBznHVi8ou16CBV95oIaIA7vxEboJza
1G+DJnNmB+/EE3MknYbf9Y4iFHzPJZVqW99J5t7lbW0DIXx16/ML1R/TMoubvE8Q
WkJAiu7f5iX9VptiRTxDKTRDCoeE1u3nf6W5Vr6C6ArAxPUyqItKNXYfY/p19LMG
Z8A0iC6tw1hzp/FIjjAADTdZQdXR+fhAM5Ek2lQFbBe+q+MXSIMywknkUiK1M+22
ej5rzHOTKfQYhdcQOEkwCmabWBYtV68unhWTbhJ7CeJS5RdGkLBlu9PDvv09G5wq
VBpDfnr89pr5rrJfZn0aSvd7xP7VD3LF5zyywkJs2S+BWMVGb2RgCvNPn/9w4exn
0uKSC4aMY9dKlbEEIVjmjgyq8Ep7Bs6iK+zJxvQFfRtFUFCvTlPuF/Ibl8+bz2Yo
93IVXTGYJcpe6S3T2KkEiYtPB5z/IEhhvFzj8UDHPZOGu1ri97M/FBaR4r1ldYZO
rLpJPT/8/mUQM5n1UBLJYR5BYfXsUL+6OVJg8jlvwp1mc/8BGFr+m+Jzc8gK7CVT
YMfHDFIM+dS91Z4SsvAKJqPOaSMyuma5pYG37LCwIMjWQ78q7Yt1DWR5vamMwTym
OFDYuwZct8BQVE4ZjjANC/m3cLesLj3QhcRT6YUvZmnnyk+5nfAvTL71lrL0OQjZ
BAeRywW+w6b8hR1x8243CSzsbK21ms/XZnP9ChgTBpoMjZEclJeiJcXncwba0E1H
wftg9zp5sndjHBoldzCDnHta/IuYOdHCV2asuSv+2TbDfV3t6NVpna0J6vMRhitH
fBh92+ysOwHmdHT5Rphyb05xK0zPHISXYoEkiZWmodqlcOAbzQzk9HWYOyrpkrVN
ZcBXheeeaps3I3bO2u/wV7C/5v9HFBxCfONzyHTFjbiPCQaDfBpzQROr5kTY3w1W
w0fsT3YIJeg+bRqEsM/zwUfiOYFlt6l7lCVE+Q3cr1Z3E+cUWlCHKrVw4Y9BxDcG
pQzo6DilnIC7wrGg99JzYVIk65DzxigVs9+BzK5NmWRGWFPBAR+1SxSRFWs6OYoD
Wj0+XPbCRPSYTn1H51eZou4xTHX/0OojzgzBcOgMQ1RMHEIg/k/U5oZ8vdKz4Khi
JqyyLflDFY1FKg8JmDhg6b9sSmggURVy8PY1F62BlYk/A+Rm71PBnRsoXMpD1Sl+
Bsq8tgUdI6R9oQ1gMZII2R67Aj5KDhryiVXYr5QXpQves8iLmSy73bTSfmHLUwnJ
/DohLBkANjSYl8ZaWLApkd6TTDjiTM5GleV9cY7k065w/+2rl9uzqx8X5hXm5ziE
BN4qX9rylTAkA2MQdFLBZNyO+qnCGFXXURDIKAKj7IoyHpW8t5VQ2vrQxkgbABEj
Pz3DZCk44GxefaDG49SAnX9GYXokMNY2lApNNU+0DWSrp7/bOAmRbkZ6ClasSGuX
5yK3+DFYzfAA0r7gYL0L3KKBh74ybaZmsvcsxS6c4JTy/fMFbCh0mt9YWwzRXDpG
85isHzIWHyyac5w0SS/8WmzXzsGlLamUd8fDEEatoVa4NQ5+6H3odtveyvcs4LJR
0Wk0ASAsXvGTrznsVn6LZpSlBa7NE1089P0sVkgJw+lhhlrJsiOnpC72b4zyszOn
1vmBNCojkLjIVrrbHDOQ8Z/mIT91PsOy0/ZaRojOPioLNkqh3XA4DUgoNGpJyKC2
14qOfpPsaLysLB0ggjlrClvf30Oag0zqPp8Yb+oTaSPOXgDk4OQAspxfnl5wr9eb
iS4dcEGS01vCXycoczfDWgkNd24YlOOosbzwGf96ZYMiAHcfcWwU2btGcwD2D07P
LtVp2ZDKlgbnc+I/mC9i57LIcCAhfqiu+LhxQQ/BrczFnaxu+EdGScGuZHjh8KuO
6/w4FSA0abANpgl287AvXaOOnRysams+0Pemmh7TzMvoqGkQycOqV4kab2csKOJM
F7+xsV+3UZ1oVKgIFmWhSJqRfWpoIgBfzjTho2v5m8pgyzqJpyUsMo7D3eTdn7aR
xGtDY+4jFQs2iPw6acnz2wWduORDMenFGAhdEiaihEqHq1XCiZ/y5dzS8wC0pq3D
QwH/0YwGcpsEE4vY+omFjo26W+uzbKY4h5RKVJ/LpOKl+V7+fpLYzkC3qjQn7UY5
j/58EwdrYwW820FK2Yx9nleHkhuEocJpVp2YRmDQ2DzC6HFMZFcsbkAo/+VRA10Y
S+r5bxd0xuq/C6R0H40Vswk5cz2RoIy3ozzxDJSxPEtJTR6Wta5OnrDn6BE2Sqis
UWPPRW1vnUdz2Gf2zQk8HmCE//Ufm7/m/KrYUGB439h+ODIcS7hnDxvlfSGSmLpz
Mpzzq4qq/DsU33PoFl/8ld2bGgiMe0rA+yNWI1Z/FnAc72XGVGjjQzbxqMOVPmi5
pjM6qsIXsdTniL43LT/6r3qaBZjrAizfdVGCPMacdbwn31BiCM09wCFXxaNT0V0m
x3PYs6K3liPvroNSKOek8THhMyIzWWKMm1/k1Rim7FF2OEYkgQxzAzu1yHEYVkGX
r028gGJ5n7qbcmpO9kLiACQOXvS7IIfU612j7tP352XqU+ufoVaE6VrjMBQT3u2B
mGxd5sUavPnqmuKD8vwE6e+l2jPNQND0OoK8Guys1xkrGEEFHxJE9d9SWIW3ozYH
GNMx5vKwIzdqGPtxexNCAKKQUT3zOHWLmLW1T6bThzQmgNHXk4k9OJ3xc5IQkd0Y
dzktQXlj/aU2hADDGOvvl/EkU52J9Pj9i+ObciIoEKIP+Q3+cb1sbocn67tjLJYf
KRxapjWY7YT/+TMqPqaiehJEqIiMtl+yT6Si3MLj0Bfr1iVxtYJyO5bj3bV50rrs
Mx+9Kr3tH9S4M/7Bk/mt8MnRiD4jo9PuAOhkfPT9uc7Y3wWV+s1gVjld+3mMz75T
z6CuP2YFrnoXyRTZvEg54VdkYaRGisgRcVfH0xlZROSWz6P6pyYCMUtHwkn1tMrV
U1NGBz5g/CDDQgTobOVGk51g1FOv+Ta0EG+xuQvxMys3FMsz8T+7NlWWmuSq9/xt
5YV+OlmbJD4hgZHzAUId+gUrXtH+6lzzZpaqrg6WLnN0t19VdyuvHH4VIOZzTVPf
mIlmu6QPMW8bNcVMGCjT9jvtnekzPpa9qQwzUZhCCZ0QgkMAp00uDxP6eRbjcMAr
tIXWBYp61M0DoPcxWKoUS3hTuOYi3991TdXIz6g7I0ub1GhAE67ESwYeFO0Sl2hy
xOHvE0OWv0fuQXY3j4FNf3CgjLlmiEOkp7cy5MPZiGqvDW+2efrPm7tGF3NBvqJq
GgYra8YmXnp1P6TbBWkAYlEbT4pddTzc+CBE+yZq1NNWyzAWgEc/d6XJvENrcgOx
JY15huD273RfuQaNKEHJwk9eV29k4W9gS6TCj27Prz5NufrvqlP+qmrUQOOpG5rZ
Po/SGVYXXxW/2s2jruvBgxqADsETdmpIITutPxWCRpbFS+/2XhdKzEXkBsF9dH+O
J0YnXzDP0XeJRO97INYOeloeODg418zQ1uJ35+gc7gmQA/zO/wHEeAXaaN03LDPR
U5AGdXcILPm1D68K1Uau+zatJVVpE+YCG7b4YAMmbgBfztsTysT7J8N/xiQ1HdxT
ZWzvWXnV3vmkIuCd0VKNZNrV8y3ygJKy+9NQnEROBuB2NlJcjB3os/VulFGIbMeD
NVHci2W/d5T9xgNc2Agmq8xYW6PuurS4ROpfTCWtS1kKdT97nm7SB91Fg3UYibL5
kE46xKjA0ZMHCP1b1631NS9lIlPi2kRC3mu44dDvqaLSDJJz0Gcmf+CxnZu2ytjK
0/iJeRCpH9ZEAR2bx5lJbdGXFclNhuEeFGbgErkdruseAxnGI36E3nNDMhlPEU9A
wa3gDBJVnuYFOeKrpLii9EXHdLsLSlHtjrxugGjLW+3W9zmVd8x3Eec69mK0yuxC
n2xdLNO8GCVdNQlM1cnWP8AupojMQlBtu1Avy/IgX+CsNoh8f8gB5K53bujteFEi
W1gPbrNTarstKaIJgAeB9kwbit+OoMrmzDWFL0D5lF2W+L3sCQsdeeXps2bOi+lv
kR2wMcqTnLObwqdbdySCal7+ZkdU7iLOcs34ljkhbaM1//pkT2SPRf/RssCaiMMC
UCjY+gIbpz00rBlkConks3Z8yG6BIGcTL3ei8V2Qpu8Tmk70rQRbwoSvm8cREdJU
ykDBu7LtsMQ8lhtu+gg87rqAiWO5yFgUw8a3pVXEK+c1wvumGYZvKYN1d6U2dZ+y
NZlvTh0ZXfvHHg6K1SW8YuJ02hisq8qdAl/rD2INz2BCVsZeSXyPKN5wU8d8/UTp
fi6Ufdg9cafCN7WcAlcPJNMSnpp2xk52DNGHoBt9Y3bJXKRnmy8Mo8uOtQZ5/HIJ
MNzF6KzilriuOXNps6CyKadzSPYX5JQiS+DW0HwxXMmZTj57SOb2quDOMiNKIl5U
TddkPaUA8gEcWA8Ch7gjS3tT8v8VFdCLLHb0NsrVjol4o75PHZXC2m8EzwOcXO/F
2ulx5RyfukLCom1qvlNzTzGOinGaB6UQhZWfV28GlLsZ1gsYUPhXbx0beRGDvqLQ
InhxVy/RsMtfYC1daFkTPxWl3fcdLLkG+rkmDkbluKnJWbbqj5Uxnlq48JDzBETY
DaJBWAmlb2HNxVDKLQeuBYn3lvjnxMMBADg3PVmJPYGnpz7yYyMCZODYYuLS4ByU
CFicITHIvnzaQF88Fn4Q3+KmwlgNMABe3wZAnee1yKDni4kKPM/twk7Acss1cFss
q4HOzDYSHodRoBkbWm1c4CAMxlnAASwjf7y1qs3GarjpL9Ut0qJlXK5yiP69B6Yx
1ZKyIL/F0Nxi1d6+Sl8iaQ+3SmZYKl8/uUueB+JFs3AFpRKDzPIOXsdCf1A1m7Gv
tIM5Rl/144BpfBoowT/3Q1Ytp4HtdVEE0FwhjW6p/03fP5VcE0x15fo0PKZnz6WP
BwxKgsh/AfjnZyq6AoB/Sp+sUoX2lTqoIciTDdmktnFDGU/c6TmqAXaMGVPRlSUO
XokGReYFp+8IIdn74k7CtFFn7OaU6f3xGaIsgyKV4BqddV3yZoF6Tcb6rdG/XmJ/
FiKVFiUAWKJrKHYs4DGrDu7jLVnXSjHSU9izMTElh9/BIRph9wUjN+PnQs1qcPAT
gSKQ0CXE2c9N5LxLNNQ9VgD5b/9iY2GY6x+ZIh8GyY1IpmLoBYyANnOs3MxAwuPX
vnAsneTt+UfergaMQkIl8hvv472FBzfx1CuY13sD9qg1cnRiV6EPlWN4/oNf7Ma6
ON7cfUw2OaOde491HfRDOOT+4iQDkmUKNRk/NRM8S8tnKMsMJUrdGHuN3iBqX8M6
JnsST4XRKoi2HQgK77f4sCyeqtvQu5IeII9uJuhlk6qg1kUhiR8XKKToem/IVVTd
O5jLiozNrvft1OU/5eqdRV7s6vBiICQsf/5b38Gv7qwBj2oxKfwUKvmZLpPMgKPW
YI/ZaWJdvqv8abSbcZkjg/KHxlcItuIy/6Au6AbtUkEHwOZ3UOnILRq92gQU+lij
3xjG506YXWO2rQgdV2zIidSkx3l2uTEU4ZD9UHrpukuRutHbI1E2jdbNgqnj2yBG
Ap2suNi0Aeiy2nMxkQx6+1h3Tz+YftVrJCDWI2paH+gzA333aq+HYX1Gc7PRnu7j
zcAt6sNsoaFSivFoGcDNLes+tQi3OwDjApf3tnxw3oCaKFL8xTnHC8m4Qp7KZGXi
7sqc4+VrTIyoxMtWgnPj673Z1vDEju/ixhLN9VzFILQrraCyXliC0TLPmFkHP9nY
M7r+xv2Z43cAS7tlwCfdiwAKli7SQz6fgw2pyDTtJ1ZAEZMZ4B2uw8EaotQGNL3h
we/+dKE+YeahNxmy8+/RCmYgITK46rG+NkCtoUrFR8YZR1DfI6LU79xWuTEtiQXm
m+pI8juyHeZOBvNN/23DpvJhvK4SlDfWQWcYrr7Dm+WOGwu9DyXhMe4sO0vGjr+P
rzaGHimMlBzB3mmLZ1hg4qpFbW3aSKsaPX3WFeW4T/bNs6QXdyHZByvohxi4Z4l2
zZgU3QP7UceREJGtDlayXJDE5xTIsBUA+5VubWepx+ZB/UO2H2rSfJmFt6A/+bA8
rufd2SinfFaEHN+0o+mUCaoLwAfSb6Ju/jVI+ZW6/lxRgiqB0wqG9zDm34NJU0gG
CdMoiMJm9oaenmMuCTHgaazXeCfcI/ywlNAbAPtdhe577rY0yVFzWzvhRpGY+Zsj
dtUa9M2NnGmR7B1I/3bcp9PHa9J8Zu78MbqB8tBnnTUjHSC9qMknIPKVxZ/y5VcE
1pTWrIsV5uhjb+E6aUIHk472r77D4Y9Wz+fQz7S0eYp0E/fULVSxVewDcou66XaC
ThWR6PxzPbzCt9VwlvNfvZiNPD2865f2tZZWs+gU/SyQHLAQbCBzghBMKZwg4ATA
gTuuxQBcBnO+HtKmqlYcsP94rAtES+nB6AsAcYd8ly046fB/aqtPin9dybkol5GB
7X+Xz6k3q5vflSLQgaJbnxoJ6N0OxfYMzj8YeOPL7OELucYvZITuSjzfJwNICQxQ
TmdiSakoVJNXseScfCCJV7twjlOTeT59AYwkW3LXOo4NF9JrlA4+Gr/nkAiDp0aT
P+g57xy5KxkYy7GWRbTGChWjCCmvb8/OefnWojxpHq3s84uB2t1HEbBsMnYyuQ7f
9I2o0/cbo6D6DkSnyxGR+r2bDta/QB/NW+q4qZ1vVvz6naNbBfekgnzk0rfFmB2M
P7rG1YwhT6kNeG1zXR+XPv/46gYpXgOYqbJdi+qwYjmE44lClXPr70MevKfprzQm
glzkgDu/bqgMRuMo6MDUwFsRJfBZh81VYU3HkQhmLM94NbmyKdsy41PIxeEMoeI5
FUGRnvHSFdxbk9MDnRM+wtthcBWwQVP+2RnFr7JP2IUOnhZegjJ9sCg8LyZuxMst
rqcPFRJp62sGToNZ1MTzZx1TWxmaH+3lo2PLhuRrW0BlHJTPQ99cdPwgomPqM4q8
SJjUE5+PUNeXhcZOyfIDUdI3GRUTjfZY6dqKGPzcZIoofZ2NqVsaCdPNJgdN8u6i
JW4w2lMr212eLxHWselz0YECouokGOnUtlol4HJU1OXba/RFCGbbgEmUdw1tnRJs
6Elv6Mbi/01elNxMJbmjgUHpxVuVO/MXBO6MA7q6VfEvMQUZGkNbB9ZYc+AY/lCn
k4Zc/lr2CtLO+0d1DVtOE6h8GXzH/eRb5Oa4nBEIK0CGwQ1d5exVrno1GsxWXmZ8
gK1K6kLMLGr3f9/8IXqpZDpPuuWwJi+K7Ug8bik5l/QPtCbEjD4NBXjSjbEposns
xERis5TpBuT5ZoJNnXULBXdTe4P3MUCJ3QjBVQTh1YcEmj0c+YQ3O3goB2P4yz7i
EIveri500LvttSfdxaf7nd3gMfuhjicYnCHRs2K9onL4oaGH2R9ESW6IED1JaVqx
6zZInxDoJ+YBaAV7r9OiWRVgYoEJ7R98NJIv5PWmo5gxLgvFmUXx8E9/V65UeNpJ
83dpfK1ktHRyZO0No3jWpaR3a9awo2mtC51EBC376RCb/0kYE4i8kyoVYiY0nEeH
JkNBy4QJOgrzZUzlSFDaMcUDIz+fq7J8BGnJj9kKvZmkhtSFHz/nk729PqR5msKu
ZNnWUp64rCDlFvEepFX89W2oBJ/aqfhzZwwcDoWDOrgOw5ri1E8gxXNMbAWvE+5H
TMVgEVrfzbG3STBmj6mrHFaxqwhQHGiLVcmAQK3eDB4J7FxrS0JaR5xgs2C863e0
TcSEt0unWcjhlAfE+QunnQL/1QpmYef+cs6KVxl4wwGx6Bd8+rClvX7hhcngIrDm
8Uwx2zzB1sco8ftuT5TJPF1eV3mUPRguMH5YVknT8d64Dzt/Q44v7J5HVLUC640o
Sm5EaG7Tfp4mHXh88wQroGmqjCW9WViCFtzqKMcCuRqBpzcSbFEmYZqsylFlaVV1
6y2OrPv2qKzJDHJ2KK8uYF1KGPW2GW2hOc+v6qAenrmjbLDXjNeFwgXme5Z4vQut
36d9us0HDnJ1eg4IR5FEsh2PN6jy/88tuLOkfoj8Dbf1MeP3HMVNbmZxrE2uXAzL
HAE9WjVPDVfVkL5FPHwV3tneWJxQCD2stRklK1f1ckpTFxaExbd3JaiTn0ugHno2
1NVioCzvTEOrLDy8UE9e9T0HlgTDpp+dzlNRpgFqFZdTMfE9I+A73SPQTXmEZUwa
sYbjEV8zmO+kDNWMJACW+/n0tF4Jonat5G9OHfT7amdgWCXdVbbYqVH6G3g7DY+o
axoly0aw40ss15YmWfZvijTsVVk7WBQlmJFn3LTCSz6QwaPaEnMmRWV+f8RAXCQW
vOxcoY++s3fKHSxZb/0OqhT5q8/fqwZxs2FHv8J04WdHfcIUG8QTkpBngEH9CmUg
+k3Sjg6Nr6OjggBmybChu0GbQ456qc+GMdSqBBq6HPBvdtXe0wFZ4eS3IqigzHDK
2XF3s2U0YldU+07wDA78esJb5SpG1HZvQx1SIBO0hFaWFcg7/AojT+5TVq90hYlr
OFkcvgV2OgJxF+ueWz8PFdEf+0ANtUngMWmDxgkb3wezg8RG32DP6jra+RBHvgXa
V52m/YTSATD6wrhg6C3Gq4Em9aFW2n0cCazhy2cORtIeg5Fn3REMYH64tsznsoOu
NYVxrZ4WjaTH+T6x+rsbavo8tE+CIPy5fSe/vE1dxRMHaj0OwIPKeFwAOyGMAAGD
y+oHO8DQSF8YuutzCye05AZhqr2lBYAWSH9LHnlCi+olTglXrI3MOanSRGz25odV
5Yy7zWwBNd4nut5KRFl3koxcw2HUg6evFcAnqiFkY5k2AjbidLrL5y4FQxsU0eZR
RP8S6AFcZvCfiQ0kzV8udvGpE1nH2IF9C7YcnO3DjKuKcJwn1/LuapqClRBtMVGt
E0S5Tb600rcP79tLn46dYJlMfqiFqNH3DKPyEoi9oDNOT29NUa5NEoMGzRGX/VfL
c+oOEaJmbFssGNCdy9xmUBvIoFN6amH7xTduXQ+vKctSPj+ZHYgufc1q51l7nyaT
PI2KEN15sotdO1pQ9c0RB2IUMdem+oiyciboQb5NUL3N6I+8gyP0aNyNZKa2kf8V
MbmjVZcg9AyQSjI6gOfGKaebKEwM0lW44afvs1GI6nTfUMABfrlJzmviP1Xnt6ua
F30frl4EuKt2U5epoDZnakgh3u3uLIlQ+Lg+bOKlnXPMvC3oZPUfl8NhMfAXVKfe
9S4WgUGj39j8581/t1YTxjIqinb42ATja+KfC9TzvvQ51AtNb/g6huKl+/dc1cnn
BNe+Yis20faNLkYl7ETMqSaHV4Bphg7g4AsYC1eyBtZnN1KfT05yHuE/znEEvKJX
IAdUyK0cJqdqnzi4lD/vpRD8kv0Ky66KGWCdvIBLhPUK2koXlrN0Znu7RE3LycJM
UgrCbHATVexPfU5T93ZiOGKy0zMUA0vS9M6n7MI+5a1KufF6oZ1y9EnvnK8O0hIs
o7LQ192KxS4UfNOlC3h3W4Yy9QmO6b3xnjKHFumV7W50npb/AnWJ61mej7L7v9Vj
ujD1fkYg/LiF7DwiK3ARLFNPX77IRxFtP+sdI2n6CIpvtQqVvgjLtMsxqjSIJaXl
4xHbk2bvuZWFRH8fddj88aJ/i2DacGdrgf/2FjRBEzZg1ZMtEN2JBBCuuG8I1IxN
lNOC+qiKAEkqPuAjqYGpesOTFZ49uLLi9mY1YqO9eCWHjK1mNlMz+ORR2eK/mxVt
wAv92IZHiMZ3Bia3GxcLuOHTrwx+m5TrGPnU9wwYVyBEOc2ObuSXkAh6IztVT3+3
uJfFdwg4AI+UiGKp4fIWWbWNkTadh+8gNdry6T97CntDvefB/Hd+j+X4BHbUKyMh
AYezxQyZgojrd8oLxG2a7AILNCcifnNKzJt9OZ9WZi2UnICzS35TPKFWMxLUsXL9
IV+afrsMyE2DxR43fWZeBNxFRXpvVsC+CslSi1F7UmefocbGhm6VKUEn4Rt0cUdh
aZcKxmmltUR/iGxULutUikJgjvZFFEy1CCH/dTzqyadwzxJaEPTnkWyz8wghl/Dc
griqlRUJiJ1pWPrxslQMVyAy7udtoJWIWOnpcJyYCJUlt9daE+tnGs5GeBndOUcv
N/o642IyNieNxpKpFhb+MswIXcuHbIuD1z86Yip/ZAFxm6c6dR6dGujTtJ7TmLIn
sZ/qpyC7ztlroNTiTN51CkbmSjr3v97jJp5oqsiLYImVducZB5TAdC8hQI+Ko4/C
UgdtguEZZ3FEtvoa8t/oLpnX0t2/wcVlGPevxE5R/0Z3cMx1nfpG+fynLjVEVg8G
CxD33Yq54VqlTYoAivgUHTQo8EPnwdtukwgLbteRNgqWaegTj1TwurdBxV0G7UoG
vd0q/dWrHglFJN6pLMpjGvfaR05MnNd5gy0PB/6zIYvyYItd9G3haMPv/CsDiYwV
xv/HNazBuz2MBPXVDKJmNw+JkudK3KzErS/mSPOMXhvagiZHlh3oa22cjclQ4oSg
cM6FNtGvwRYvjMEum1lTq0pUA0uMPzn/jekOfGhQrldDjMPqnH4v8YYI6sOzp8yH
WaFX9n+yL5axCMjMlrtfpi4ezMUiSOKU/t9WDBFbtWwG3e3TCYh+6OM2FkiAAbH+
PsANFWU5UB3+0dbQnWpPtZCqyNRXJQlzjdMm0RJZkKA8AVG2dpL5vlxAABNY1C85
BsyikZvfBkTKbljYjH6ku2r4/KAt7J0gaJvr/0HjXitSiAHbOWtyOpP7LMW33ezT
cA3er5B0BGMaK3U0F3ySKMl+3VOUcV4OW8Xq8PSrsHiq+OZR9Ltsjk/y+gggA69g
m2fq7jL9p67zlbJs0auBbH/3Y3kyHrvDcwhdADCLx/kwiik/nYECFIU22oNcqp3Z
Q8HooH9pqA3cu0YA0pL5oJNYp4ubL748zHFK2JYQj2cwuxlZmI+DSCUda4YFyFNC
ZuYnuRguzK4/eDFU8/aotuV0hFRNfWQdhmSRAqhBHC/LoSZFZghHYnRZylmcbtb9
PGp410KlKqIHM2LbXiiycJxt0kiHNux6KAY98TVMLrUmkeR6ijOHIRgd04wBPPP6
+k1DDCjKZac5+T4p2nmdRPzX0dD8mwINeQPw9qbm3XoXF482efKQ1IyOXsm0G9i7
WLzDzT7pUj1GUovGcWYNcQyQbjC7jkoVuTIxf7HOjdYdUKOU55XeEFNATKp64XTY
BDc6Y74OI5o3r64o42nIqaMMhNTa3Ga1PAz6cdd7TEsh32nqyEZ0/+ID/Cpd0vhH
pzWvQDDF564YcadgQU4LQqrGj6Z0gcBOt3770lHMtkc491n/QsZcRjh/XCk4NKQs
DnC+gM0gMAwKRuAuFSfPDU6VQr2irxeD813Oxrrm1PiKkFR/bLpxNk8LLSnXjHiD
xWgyE5bVw4FKrQPpIY7QQ8MwASe/qdDgo7P5asxTSPrro0nyOernky8fZCHFuOVI
kAKChZjGi49bqYe2ggwdu0OUJZfVif5Um+nmm2YjHigRU4ycb5pO53iEWkV09ug6
wZ3kVXE6XuK6K71FN47KEs67ra7071NNr94httEJdJGicndaFtlbht5x2QbLRGy/
dDgeDwFcHppU4Fq/0iv+vQtdWyv29sEhHMqK3WSeA+oaS6woXGEN3/bcGKCXmJUi
1/zVx5sMDOd3pNTpWCH2bdmjAINSqlgsuWMPA2JaJcvFaV75EzD6J/tJFeQlUkf9
NuHRlwBI/+LfOVQUsJ8fh3yRnd3BUN07UDy+WtKaQWaOLpVzk435pVX/Mps4k3NN
BPFFLaBAehyd8LaN5sgaxTLR9ZiVA80xKVx7oXFsO6gNqgnr5bH6nHw8XsI9UQSx
0wmo8ywMJzRcDI5dAtAcQ+ktGEKVKUCNTsTD4otl/JeKvyNppzt5oX6fkZxCp1lM
LsLtP4Hd499HLa8UGUm4Qz1FyH0AzobkiAExWn9FCGIAk+UlBJGg6iEPySNduVYg
b1QHFwV9pW8xIw40RZnXu7vrm6Ir+7Du7WYIbeiOHMoTQLm7JY04bEZWMijHb7zi
qquxbihyVzw+3Y0jy3c8pKzi3Jrmjx/N51QV9dSoudbid7aGSQncDfvAof7L+FSa
r3VylLGEG0tKx9mx4Gi0nNC4kNUNnE/rBdQmIdiKszapwVtwmE0vcz6u/35jz72+
LJAML4tEZsMxHKbyEnlKbnIdh3WWFWgxEyW4XPTNQ07ZyuIIdP6f6IhFxe5PD/Jt
4JWz4gR/LcRJMJpbavmcJiA/j5UwsG+YuqKiGpuXYR55tkM6RVkNAhR/8Ap16cja
Flt7rN3dYh6r2OgLujobo2W0lUtVVlai4U+rC3ViAOfEEwJ6i26hyXrvF0CJD3sB
mm7A19bawWR6moaATnxViZSxbmZQywC+FVMw2d1DCFbrduttsuiX1oqYaKHeW2vs
LvWvaO5NDfPB72YoTKvXdIDvbPKVKdnMtTQUUOymUshlIiPL8LCKQhNvljRUD2iE
m3A5SCcbl0YFhGe6peNb/8Hegr1aKciOrg1V7xqgDI6LdHxAEM4DctfNfyRxEF5s
6wf7oQjQo3I4jxM2rKs5DrUuz0GlijsqmCyD6mttRK20XWxMl9vf6olxwWWAHZxg
kSPM2UiIXX1rj+hqZ8hOxqmew1mPOaAAkSlIUN6poQ7YBfrnxKsztuII6I0ZhSqD
uFqldso4rPDEcHN4Xp6/El4m7wwdHlTMq/FpOiTMpfg7whsldVtn+efoz9ayp6Na
QRI7CqJ9tfE3MwyCj6Ia7dVomsN6z0t4ka5qtTIvRSXb/fleVB+X+2j/DOImYebb
Y7GjfHpJSz9HJCcZS4IlYi+K0PE75dfdNMyB7ba18/ndehRMyz7uVbkV6mVOuVyR
AP1HwNYSejqCVhr81q221X7SljO80+RV0SEUBGrUUDfU2qOGvlf7ORETGXAGQ6oe
EbofsQDTImgdTPghaLnhobjdrJhnEnecVobTCBkWjYMqNcIlIk5KqL0qFoe73m3t
m/iSkwUhy1gWXZMv7o4Az8a2ZIHegFyRPkRa2FiIaoF8DtnmoWDBl3EThkeExgrA
q1g8IApcETNDTJ/1T3gs+grSMC470tfwGeG0gKQPtjwOTo1/ZQLIpx1qMAelXAt2
034lDffxE6qi/206/NbVfu0jSYXsTyjQQU4Wp1TI2ZJ5ouECi6TNzPxth8L05iO1
bAKAjANsE8PnrEbQnu1uUeE9A+IIsc6kfHE+VflEvHrDRrlpVROxNm31Y3HoRHSg
q7sVGTKSZ467y7k0rw5RbaFZdvauBMbz27iIeCruabvrSszRXuZC0Rh2jGXMVtaH
20CRQXxwGwf46js4y4kD1LnIU/3WrTCDx56V98poDuHRC3ziDK+h2wNZL26CKD3+
e6L1n9P+q0Xs55VOVLLzLCWsuKdEAS+jn+P3LhUsZr+IW9schxyjtKGpORo/E9DT
88mh6eI9bRBkGbDeaD+bZtp4KHiGMYQN7F3pZPsWB2gCw7vhAP6KtVxDft0x4tAH
a41xZeE8vnTVvMu1K+nPF4io+xXO/ouMMI6bVMX1F94KUUxU5YIEDC+d90TOy32D
nvUNG9EirrCBJwWG5hpEYuKhE7mmXupz2fZdgitbdq3R3RcPmji3IyJ3J58q9T2F
3XWrLt4o6bR1Nd4uTGhj2WgiujjgrCTY3PUqkjonqV/zBI9aX45B7FYXECN2mybV
4imLdyyJ4KtWkgOIb43/17z8X++KBkV9Ha4z1y8nkBAFyJfzhCLBVrzpsLXynPxF
CcAudoUz/9GuQ2x8tN2hJd+bgcDmY6aIbrQoflMddSuilSY/j1MKYyyH6NNx/8WH
hV8ucV35DYd7AyC4Tr68qUEXMi32ecNWOmpHgxk87jNxrD0lqjCbqlOvzHbwN/uJ
7rKlrcRmh7n9VvfS5QWPJ4NeTXgSh44b5Ttv0VtXPOh8NxwEvqYa7Y/qUZutwjys
Tszpd1DEXQ3C159jBV51YFHxk6962Pw6zHq2jZCkO6OeuYy0xkE9Ovm7OrA/nfkT
7OBV9z1vlUf7g+6DdMbNuWJu2289z8lEc7TNqqhwFx1DhuNXfMXCO3/KfsFj5pez
t3ocuByo0GWrUwUMezgOE35nowp9lr4tabhwbLgDPM66Jq43ZDIvE5Bby1CAObqe
Y2b6yizl+MReIaorpygnw4drDBmsvte92v/49aN9dj9NPYljHh+Fk0hfHVsMGEJv
VVX1ons6c4hQlpRDb697R/c/a8rT6QKKLbzqd8zpVZcHUdINTkoqKPbhBRIAOotS
z6bsFNddyWoNzo/kvVDEJckaX0HuJ3mc5SVNZBQPHTAv2EjvJ14Fww/pxnFJhhh7
24LhF02KFTvLEvwhPmxvjq5nXNSZEOWLzdY/NhK274+sl9gsQDiLaYHL3M1RAYnj
X8KaTC/Oob3+6paXZDp3Z2bCpZN316mj8FjYI2HhxDDwERLqTnOsarNP5rBnFm79
CwMvsy0Bv62IqseQ2KJ+CpRk2XpKmIeaEBGK2FQrhflzNJUuNnzIeZf7EnUSBimv
KPEVQAXxAEbN0qTq29YItldEm5leWrRF8/zpR4h+HaEq4xBWx1JgHeeeFX74XE/i
YmJEjjLQtBZuy++yxq/2YY+LUrHXUdIZOLwzTJiGfs3hNxRaGKjaT3xuBhN2bgyU
BIFInpa4aTLjMrQ+9rTyZKamaVSmVfdTY2c5XSW96VZ02pSG0Ff6qEkRhOv7RilT
hgsGMkwLvIzr4CUkZrMOkfXvPkJ2r0/AYN78DLiLgLY4PGDFJBXoh5WTeat5tEDA
hD+q3mh+NDYFXAKgx79JF34XmSHY9h+obYANW8jMbccGu6S4GhGYLnNk2Ry+Ane1
GCojpSVydtaYd7HdBwtm2Fuy2TGSHh4JAG0gf4qEYrsPHMfRgOtCPks1pnNBgu0o
wNN9l3hXOgSIL19EttTGPlykl8Y9qXjrcsSKYFkxOFKgDzyPCQiTA9dth8T9iSOu
i5AfCFrW7m1gsfHoFlm0Z0M2PWTR4VZjz9KWvt332qxmfsjpiARr/1Aq93L961dO
/kQPpv3cyDBVhzCMnWLFE5WJv8BWwWjB3lAnzSj73qfMwosgVj9jVuoZEZItMMrb
XGwqDqfE7FkaHV3iGfxFyMOzASeKaAGxivBhPtmg/vLApkdDReAoAU7F/gdrqvGB
UbfYx0CdRULE8GyVjDy7H5AGGyW1iwV+2dh6DijQGon6+vRDhwj+hRPVSZlt4Q2s
M+WkqNhctKEhNfpbjoEeGgPMiT4UUqTnfgvFOFzUVz83ACrs5UtLL1w2vnhLVU0K
IBE7Q+SGdvTTvwio/I4cNfkP2beaKKzSssOGlcUfHKFSjk1NyCMi0mCt8Ha4/5E8
3XQ01HqFRJuk75kE4uNSpe5qTTKcBgOvn/lInXFNoGk8Y9EvOm3xz+f0WaDbediV
s4LqRVjYqucWi8Y7cktINb2nPchVE0KYYHsneE9ti3IJDONmcs8ATQYO9zrIV68z
sC84Lj25B+KZy56HfojKrQrTFBNYwhCL5ZdZYjGryVsmMSTHHtK0HV4Yo0BCbMbS
/6pZvTK1bBC2i1ubZegSFLR+DBiWQhbVwTAPc4khWMamdXRkdO1K+hEVogKsITLU
v8GTP5QMYZ+OSyp52QG6Lm7rWdfOZ3x8LiBQ9xjuxcL8fCOZRpEM5n0/c5eR9lia
24CfgMC5vom//bzF1slByzNigp0AOywwV3h6aYn9TGvvrTvIf5+4Dpkx4QuM9cf0
I/Km+p9Fjc6VaL7BIw0HULAoiLX7xWKl4R0QIFWSiigxJBzcZeBgG/yucbz85lKD
ZYVy2k5hLWD5U2faoyr7sU/ikWOZGpWdlMx6Bjs23FO+WvgKwndid233xXfGhQ7N
p+8XRoqouYq2IFBPtoanvOHc69FOpXG6tBv5bfiTbatTSJR09+VQq3vXuidJk5wV
CwtuURJG9HPyR83IxkaBUVZyrHlmwf3HRGZRbTqvPO4FO4APJ/y0vwzJSqJRqoMd
ZHk06GFY5LLc466pUGOPYKKFjh/Zm2mLhkx0H+Pq9JsvWdjEkgumxwdXKg2QSPCb
DpcHlssbxhsgUVzBwaBQALHJQAsn2rhZeI40fOthKW2SOZJBoFssBCC+7+fUxBFW
48sBokdWYmJK73N9SzCxcb4HizjGiM64JyrDP7gm3asFBjj+Y+KAztvUrtXgkOya
DQONP6fEB/gcWeZKZLgzHpKiHRNe2MI4PjP9PyauBj2K8pkchPvBaZdeWsIGVKdp
UqroZkJ42zmVfrSOkXn2c6LDi1tMIAfNcl8QrInE0reba1WQWfCXjrcmvFA60FuU
L7b5DWhmJTSGlUNxcL6tsWfvJw+qJmcCjH557fN+luG75IqhUVnhbNY9qWzcLnZY
ZAKJ9geogJjF0RLRx3KxOhZaXvbOZ0MYXkzSTVgwhlSfRVPClemffZAjXiTrMeKf
ghFmV4Qvdv0CObeWm9wHdiu8I3mt15fh4p8uHyvzd1tL3THr+uN/4fvVuKCqaU2D
B14GcGYOZFXiq9S8POd0Y4ST36TfUkoHjT/TmHTxv7u4Pa70Xs6D0XIo967QAtg7
R6tQNnkxRpc2kusKT/C5B0iK0OiabSKSEZZlJ7dE83LGfAtN5s+1HodpVeY1W2S2
alb3pzjVc5MGZ6QnVSnapNuCJzyhNGbH4K7HgPjPYt4vQnwhUp76OwcAKU8sk7xy
2DAvOlyh2KXXFD2Ag++gYrR3gRHFehs48T7oknJVhqrIz3TtDj4+La0Dm48Gmkk5
a8NsFln4dGL41+vn3yRf6rj1HJafVFhWvI/71dn/W45OPf6SB7ak1gNG0RJXak4+
8rhgwotqY2ZteQENn+rusTcFizsK+pqWwsybgrlfOwZwgqL9f8HFVdiQaDeXqXBe
Ay4q2ac0IwzS21gPsOW+DeNUS9HhuNGbUnZU5HVzvbHzQ/sCIn7GeGs8aY7TjIg/
0uubXyU2TjpPbMczWAmR5YsBY/h/n+AAOYoG//RviZ4KlWm+PWUWKX4+OY37uETw
JDU1SSwAD4Fj1zVtW4MBpjABiC4R1zt3sM7RdI2BYBw/zkA+azZVcF+hWU/iPhTk
JsQz8gc0GMLkdDrFCjmIYeRqMgiStbou36lORkQHLYaYpLdkhXKR6qDq/7UeR/nO
xlkK0E+5WoYp8MWD8JE11z0PG1w+fwWs1PXCAb5Bb8RK4VNwRUO1kNaFRZElipZy
ATka2lmd0mKfaF8O4Pe5zzSok5GDQRyTySy63TniOfR+tLHUJtsc49hDfCuWl0Sd
V+KsKrvNQ+RZ6754w/3+tFPX+XN4YOx5a+Su3jYuhUkuDfbqtVXatWeWPkanEvl4
TqVRS7mWe8zCsKknknjDoskDad0yOUJVn2/svffcuO4YjNzwZ5UdU/Usl0DpSU+6
uR7yGu3QkCbNTncswNTh1xNBYqytBpXUCCi1pMTVJPV5gMZ65e3xVxWgIgVntaqK
9QKbezYeon1p2zn/vNuV8VpYMwIyJvn8VSfdVgl1qdhLaBC7hywOJDFnTsDtuLpx
EeGVOo9EsRF5Q+c+gyGCZgROC5N5bCMNjTMZubK+VSG+ivf4srl49PY1b0e+Pmke
n/2vC3m/vqw9n07XXGtEVsIeYQzpoyMuy5vwij0+Tr5TyNqlJg5n0tJby625nM3m
ya3Ah+CzFJBLY5N7/aso9IJpr0KhnlFkLiQcijDCCfxddjSjTU0xKZqXXHn7s5W0
+kSucFmKOjhZpeVnMM+2XH5dGrTyHgzHxPvEb8Xfv6V30KcLJ+WMR+nl+h4GEAoO
vPpxdPgS9sOIS8vS2iao8cYhWbWO7ELm4o5pD4eqBHZswKHMp/lq1AeU3euKw+J8
6UWoQNHiSoyBvLAqfajHaWG0PgmCBny35uAkZD9XRn48RgoqBg6SrHRz+ueoYnbY
cVAGRUQLbolGQSMJrkIw+rODXlfPrHZchZuOGLPejwhT4DQ6HsfzdRmfaH/oSupS
twPh2354ffizI5YjVI9xNE9+ID4upSW5Ld0JHgUV+Rm45WeaZ+zc4ga6AxpA4CGp
Jlq+HCeDoFkJoFQ3TU6E02YtWFSs7qYr97xRO2CAX3PJOY+QHtIImsRfTEIWAnfT
QAVm5xsx2vD0DSOfOJ1kaqc8OI95gvEeXXkshngy2whdSPcoxJY/a1Ewnr8+bXrr
Y2sfoQ7pwggQuZAS7S4nviaJm0dF2sNXfMXbciP/ro7FUr1t3O8yF4tNX4SkaNPK
DDEHz5JL6kUA6xZqcPX0dJ0kUOtBe7n9VS26IzjOaT837w3wh8cfybHBhr74Gf2N
TMwsnmfbqOvnPprAlQIEbbovl8V2EIGVezynfL19gUoxbgC0v1+kWov8EbWYTwZX
XK89SNRtiHWVTwaskRCF1lcSCDeDhNq2WBDO4E0yBKZpQXVo9pNSgMrCIaR5tBK2
oQ8KenCNqgd174UhuWLB03+nu0k/XRZ4LYHIFAigI8Mz9rzBkPMHuoTXhPdVbpG3
OHKKwzmZ8OSInx3Daj5FgKtMsQLOlcl+9VdVItZc8QWyjTs5P7U1Dh4RlFmE9Dl4
4hD3z0lRkXRyGI5LCHbp2WLkpARoNB9sM2urlkewtkqas0FL4aae0XhpJe09TbPd
bm+HMSicqkPx+3UCNeUsjLZvJYtxLybcAjo/ZPL5+haj3UYkPX7l2mjtzTMcp332
IKupiB3pT15HsIw0Jtq4/sPeO3/5v/hqh4JVhvcVm68Pbfv+8TgoEypmkxE78mWJ
BB01ZSgv09SFCaJOW6j2xcFNOh3Abak2Cpy4r4OedUbWPIL/RAOeGwQ022G+9mxb
kz32WnEzRzPmaZKHRPtFCaQUEbfteX8Xu3B+uJB97Hy7u7n601Lug8FY+BLm9xG9
40N8MhJuCV+o0TxZOrSigJFEB4GGxVFVygTt93q7m1PVnslH8uX0fol0KzaAKLWc
RAyhkGruWknzy63LNZTadJgCIWt9+dV1pdCyJGR6eQLYqwJi9rSyDtaCi8qCtgco
4UxNnQT4LHe/GhqETcV/lV9Gsb5rErik735flsaJauPjlNTthgfzUOz2KLit95Gp
7DdsrdbEX9gKFF6q0WvTPnEEaMeIktulZdoFQ4A7nIfVJ0Ipv8xmChumR42sYEaI
u2gZfEk2WHSWg55TYz17ecvIsNtQYTatpdsM2r/u/UxC1cf0LwSO00yHY4zis5ns
n99pl8Zpn7Lfp9bQ6jIBcuY2whYzHjIXM0NBnXGrmCRFvyhl/0ESbYHsS9ZhjG/P
fOzCrZdY8H4rKDTW+4KvKFDM9QTXYSvDnx+upfZqqQLirnjHjAyGBs3P56xABAkE
+ZTiiLKSFolEqS2KvP82iDCBD63H7wKKEZoPGLuNjIOUsAPn7f6zCMnhCDwO/J5z
vMwvzablq+mSbVtT/ZTQQVdcfzHS95/jSFdD0XXj454TVI3RpInsZbd8sfyLVgdi
JZTS098W/FNyfCzImG13o4p7xjF+iv9NxAFA1B+ukQ4OBPMBbaaH2MOkfpSGUHn5
4oGxIyorp8RhTTwoJC5K7F6Lm0hldL5W6hUuVLEDsWMf39oqtDoG9JXyAgq13dEx
P0/ngs+T/jLHXv8b2sqOUtb5T8nJgwn1n0OKP1ZSO5QrOKfg5QU+B4SWKQAaMRPz
NSJ+MhBS8LPTO46nsyquBV032fVcMOxYcNpx3iJ05wd1Jh8QHET+baetnudt2ufl
qtH/diPQGawy2oz+CfkDkhW9cnWXmmh3o71m+0owENR4RunvIVAASscQ77F0jEiw
e9nvJAN0OsTFwz7wzukrSEgpLkzaKgdiEA9tt85ng/Jn9mrrell0pR5eKIsJJ3rV
YN/lsqDQbkWlbGR5yn0m1b2UEGi5WcuArfkwfOp0EHfoCYzZ/QZ4cug+iSgt+/fB
qz3FZgrxMrpJP1azq8NxM70OAbStzbCnPjpOSp4ugPK8SmhshpRQXMLuxS1Uec1d
bbUSy3RbhQhFLsXb48v6++GXP33EUMA+X7u3zyqlwgDjqonuc4edoaXDJyLpkVse
avomPQnHys0JfpzRNKQHB8tiuHJMsCMw691/cRWOVT4YVFFnq75eKbdP/Muv1if5
1SbTxdKiswpwQ8ONjHNI8QbsoehvFvxbi61RcRF+Xm2JP0bOiCkBWt5lU5xby/qh
n64mO5/vLhoGy7+b5Jqoo/hVDP8EvOHtW4AMyCY1LOPeS8aJIHqjPtDKtPXVcuai
gLEZoJG7p6fXSSyZ9r7iGcCvWBPfCxhLLoKqTH7eFOxsCKWZaDDukzXTJ+fW5wFN
zGl1GRgA5KKsBbIqwm8vPH3oR6CsJ5+jMOrKP7szNfTLhv2cZV9hPzJmDW+SHF6j
zbG7LMLx80pHvMYuaTe8WnEzLQd4U4DOURfdxex/iQ8GOx2Agl+itFzJO8dXzdZ2
F7m5iEtqsCDkw2/vPTU+n1kIt8VC8EzGhrTc6DRO/eQXNpRGbXVk2Nugx6gMbgIL
bwfUpiCO83Bhf5y5GyLk4HURqp6aX3DebtE+hrVarxCXqJw8fYl+gQlTMti+dqgp
gXPHD8tMKWxnFbFwFzfVgd6eRLS2quz9FLLPUkXbnla7Hakn/FlzpVOrlyzo16+m
aGHQ+X+SojG2B8M8BVGIklQMhScTHE0ZAkLYJLRIU4UJ86+65QEl57SR4+Q8qISh
QfdHBu65ILeuX2ioBwWRGEC6RHp+BHVNG3h52c0xu1wRQnng9lWu4YNp90VzGQHI
fUVLKJT8XTKdz3e7vcYqWnCB5MI0SPv6mS4qLaPKuDT3oblLEqIJRScq9h1yQxfE
SxNO4BflChDNrqEo6JNFD3YABNj9gzostoPsxsLIYTik0TVRP6LzN7X6HplOrIVx
YMqa0jsR+LvBqtsJAHL57mTqvy32MqR6WJZk2A2b4wluKj9pt3bkg31sdcng30RX
QC6PumIFVAdGn9bIYIXHLdBzsFlJd2ZDweLJb2W1wq32cfPjkBoX6cYrziwjF51n
MlkWqQdI9JuPn4EdYOWtoyrsJDMoNpmwIZHjykFyJV2dL+WwsrEy9wpVEYub3mrm
vvM7VWkFYJLvj+wubKfhxpP7rPUnQZKY276N9C1cB+J0y7zt74PqKaGy9REpPI/F
4RwLhiNC1W2PaMcbN5IXPneyVJELVimL2/x49xhJcX0mc5XqMaVcIqaWQ5ZII1s7
hHjCC/HrCOvWExSsvzexqI6kFyUkI93m4jhvZwEKLIgjOZAB94Uokr9yvWwuyCLp
i4r/VHqLqCl3Xz6SKnlejKsVnkL5MThRG0hXFtS7y1da1lhwjkJpmeuJxQvkPd0X
L58IGtVHqQcGsFRnXt7qHMDEHczZPB32vv70OuQUU90xVzAr52//g561FkzmrLyL
c+4MmdsJAcX3xxE54Vd810gCRuAo1m4dBTmdqs0thhHyCtFjanV42LTsAwCou1oQ
Ab1Fd/lnqTambwQT0Jb5EZEB9bq6iytRJ1zKDTGDKGJIARxrP5JNlbt2l4dvd05R
aE99A/VbPbljouHQY5qTcpWfET+Pw5OCAlB2fLQkhb/BMHTeI8lSBmHEmOPOId37
pmLOxjQI/rveC4M1yXpjxs3EiCLJ4LLjxHnx2piYi4aKi0TNmFe65b1y8kf/1ALC
FIuR/AMAnJifBEgPYVOF/P7DhkAMRpiUohgnYcmDRFtXHXbqj/qkMlRF2DJWAhmX
GBHPBzIIjU07ySVXTv5bCzrxdVX9BD6T58d0jjSbWZwytTdv4I2kxfbtBbeDowek
gt5Tyg/nc9v07NbQH4HvnxS0efnQD4PPjPH3i7mrGvNYkShQ+MuiCy6jn1gxAhS5
hRCNo4z1Qavwampe3YS8XGElCVaH50E6NoT1hi/vn45S2TM0U5EJ++Co4iSqOwzZ
vBjoBR5t/4A73iR/fKvU4AR8QMcv+ZeKXpin/EBYFmSNH17IKXoEgMqHsle+suxw
aqtf3z9WHwN8wbnGjLKpTZwxsk+QV9qKLzzxn94COQCgzJysQO6Z1YQQAamzW7no
VXlX39b6rtDIwqGngUx//Mw9oLyfr/Ke0FUHxF5FO7fsp5P2ORFicHkZQSjKKxGP
Ji9qaFBQGXtbOd2OEbGmIEZJjQC2EEbPY6F0jit3+9x+Nyvgpk53kMQi0HOLgLm1
rsBcvAOWBdTbwRP5HP6JbfeZ7GSPiM9KthzL6CRHCzBmzF/dgvJQID1BdYyAg+Ez
U3E9ylJfRQHVPJpiELo5aUnHir+ITL5+577OHuw4XCnZg+FXXKYqqrQ2Ic7z03Ud
XTdrnSWFjLBus4YgvXAs1CPMmVdw+eMeMQlt5yBud3w5heP03traxeNC3J8xNy50
N6cm2M0n+708mgNvD7IHAx+wZtZtFubwLx9IM3VGDWKRd6jEbCFEoy/JFH7atx0g
XaGrkR0T4egcL3voGcCcp8ywPzEpn3tqkUC++54nONx//yj9smSZjZsACjBJiKo/
Suu6PNT8AbyNPLKdf9GP8IWcHybDWBXAUk/lbflfzwa19mvI4f5JCef95/22WBym
ySLDN3cEuhTqADN976SClmnWuTy2Bf2PKKZ6AOaURLkZ+a5Mf4nvRu/zxHmJZn0V
aQG6E0vWCk3MP1DFPKAbLGlYxweDY4k/G/pEEiPj+pVSEZ9ViQbaHa8/+4JZEEoU
cwV303C3itTKYRxsszbvzDBE9rcYBD1gFOAkFQstfBvWViBC+GIblp5M4E2jTLNX
4ys0mm/jXvAr3tQYdcsu7vwuaxL/xjkzqEwuxeRVf8Rvlk2Qf1kJoSnRqPy7U+wo
q53MxS/fx2jxmFNg0yvFJCsBBEKb9SN8nunjlvM/pa7Uy47Az/pd4WK/WXJXPsen
sQLMepmwRLd/mE7xMWgaS4Un93P3Cy4qEfvf2VmGqo2mEzAXF0+FHYKRHp5HUxG6
AVzrFRJuPC6Bsp6VaJa7LAu7ahxHXlGnEy31xyJvOYZNwsIEFvxKqlxVIhF7e0n1
hRaxXiCkl3Bz6Ntq9koGLWlICgK3CffREMhPojECtPYQBOBWPPNbAAuWXMxW6eOp
6bcxKvB2R2Ko0BtxgZllcd6ZBmUZE3W6tvPvssjhois8F381kZ9IEHLZfNdKKTru
JHp+lnpSGUz09LXmJfzWoEK1yvbcFzJfBqRNNTyhgw7a+Utyel1zheHU2o8fPI4n
hemsnH9VmvUoiXii0uUKcfbe37SBrmoPHUkUmj7dlXsc6rodvTs8iWNrs5x2vFZk
tAVougvPm0e3KyVpzzXOHhCTuXnFvhdGTHQjos+9gEBmz4CHmc383pHSxOLRlK+x
DfOaqWWM+2pGlOL69bPgUw1pYXgqRln9kEoshnmkS3EvnW0JwnEncFwDcnQrzWlv
NY1Ca/B6tN5FtEV7fcZloynOYMP3LogLhyBCRW/wqdZ3ItjQbeqrGbTsB1Y81QrG
pv7V5uK4CmTsOZX6CqfDtnkzG/+RkmNIN1zM21WzsDs0f/YVrB+j9SutzGLtIKKt
RJ0J9TjNBiVyRl+hh28KVKtwOyrojgxUKyUuXEH+AWmt67vTVZYb/AQPIau4/6qP
7+gXPYgWyBWmYSIV8Iu55PCBIhC+IRoxHQhIvMEpx30qd7NCGw5G5ITbCpwHcrQz
DMdgY4PxcrQO4pmx8/bEfAg5Cxa29cknTPgP8/wlebTgSvKUQx3qGcMqN/D/Tchd
TRpIUD/qWcLltdC3js6XzzN37ZjZGXP0m72KmzPUlgwffATod/ujjjzQBxgEUWxL
IkuLPnYFUstMB9/Q65+1UO3CNibWNHP3Qm6qbD4syyPaJfbXRBY7AU6LyFcu9ErD
5CFMVvKMOOfGpY4cCuE4bWA+q+wgAYk7amzaYL45yoJdaPn9AXTuqhBU4qc9fhux
RGHhQ+EOLzKsgIQvL+nlbzuyurSymGNXUWGTjrgyWuYXgQXlOYf0CtUoyOg8cIIO
kB1duOo+RFpOKRE051m/HGuw4LMGQ0GBntotGph8SNLn3Lt0g1YA5tYqc+eYco3M
ymNgfHL9VuI7cMXfaQDJwZJQTRv0epWe8v+48V8D5sWjeGPTX2AYcTaBXtUBG5E+
NgUtGIxut45qQZdO5fIfBZ3KrB4cf3GS9XGwHgsYuF5smF1Z53M8eIEEgcm/sqXl
KMvqwrsgcmb2R9CW082ZVbK12uAnNLvUqKbOFaUZRRAfHLJ6qKGQMdTFx2XTaZ72
iPCJn2ObJvLT2WEotiMrJ2UMdQrgkVbW2jz3DRsRudb//8g60nppCS5N+IWv97uH
Q5/Qcb1lKWl3KkSAUc8tQCh71+FNrfx4wiIVAr0k2kMl29U5qsAOeY63fm1srVC1
aLRZOlgF1xeDx9LqJZ/0Dpe8YLObRBiqM5+8c3HCVhIpX0tWKlQExrY0kQa8Cly8
BaLazlw6XgSEibdLTPZZaepyyhI8ZMU2dqbJ50dXQhANo1lB2S/JeBAAb7+FDUJQ
0cSVjJmgr4t73hT/GlbU8iPYnTgUM4Ph8ThhFDfesg4BMi5CS2ik+U8kSgaIE8q1
AAKjsQ5GXrBvDv0de9MMuTbbgDE5UDP7JFOQnYaPSFio5LJaQfTPBxHOkVXMvTzT
0tj4CyYOo0Ib6jKmVwkeaExxgGz40M7Sbe2QeIRwam0Y7NhvkCVHIX9czWa3fGyz
Tal+NqnXmcaDEfaMkAurO7cYw+PR8wB5ctlLsRzqkmT3kNmUOeDQL5icaAYBVHmQ
lSEGyaZCiKNMXbWdmAVsse9j4VkP9xqQjF6BN1x6kwsD06wTm8pCfW7bNPjGyE/O
qxBsb9vou6UJKRy5UO811v0Le+VQyoV1ZBzlvfKuxEdQuuQkHyJ2yw058phmhbRO
H6bQU9WPNE/t9x7PHng56j0zvIi6vYMvktJa1sNGbLN63U1xJq6c5Cy5BtGJq2Vo
jppW60Pg55A1b9dTcF3bdabyqWY6J0WHNkHd7DmkNwbkO31dWrpgu4oWVsWNw5wf
HTGsPtDKoT77DAQXKUV4GmZPV1dxydMFnQqn/ZFImqQFQzy1TKI1Pl46MXoRKSoQ
3eNYdXSGY0y35DZRl7EVX4M8PhqAAs2W0Kel7ypJf9EgZInsi6NQKbnf3WuBvDH2
O9Vf/tb5o9jO41xm2z+eqKHqYUJN1wnBUKGdetU5A7HSWr/+8u0YQIMijh+BrmC6
dLbirdrr5sopwz3VCu/9Z3VrXEBGt6WdVAnmS+tSP1lkzQjiJv+uIxo5Qw/k/sPc
pTn8GTjBzzx9vCxrBXj6euSx80Ojh6V/I97GZExGxSCgBFRYJpP0LLgnlASkh3Rr
Ca4rJhmDcOUgoV5Vahz0wIdReGyy6HHF3EG2DHnCBOI0AGnptt/g/tfsbf58qZOj
4KPmXU6+KcSGKnqdvQM7AfiwFWeQRqkgjWDFZFqaopLL99jLbGgluemG0ukLJDk7
U7WJCaz690jMalt9kUhF4MDu+iWJEZiOo76U0zV9/bYk5OF9QbN5PkEPfJEeidOj
4i4ZNKVUtSDuDU4uZVGakwutino2pdhGS181szVe2FpouRcpq9HJE7KYt+X18JYQ
s6dUEoXLTxIvAENf5VuA5sFv68WzPYnN/4iO/lDiAde2Z6f51I+nLvR2c/WcvfeT
jrsfdP3a5R5Umxc49slWQwbzDIbT5qY8LjjJ2pXh9v7UDr7200QYN21l+nqeUg7l
ntpu3EI3d3bYRPBrKqdMG5QpVe/7AkqziWIk3j8pQlXkMU1GhZkKJlBIq8Ir1zf8
42SbfWzuC36a+lprg5x72gsEfq6Q/oJzbPnUgwUSTAt1lAKWjckG43OfY5VTR40O
IXGq4YMSPSs0e2/dyLIL+X//QRKm75sd5YBywXR2iNaNsOKf3AXr4gRMk7gTbB8G
rQ/2T24joxwwLpNUT9EBUWFvLygMLL/uvICcIOVQoMWk+DdJqeVILnv7xFEr6YEN
rm9iuSMBHAwT7813BnBUTLRGJRxhxj+nVcMVDNFa6lB81JURjGzi69z2Z9gHrBV6
agN6kHk3+9IXLuMv07LmulInip9pMnpS2hEAJPEP/gt6TFhBhMzMdXOJWDyEMvvw
KVt+Osf3LBQaRv3p3dg/PIThbdC3hlFL0FQ8bdv7CRsvChGp8NSPAKS7bbVhmZqx
Op7ngWnmD8J3fH5B0h16deTvudHNTGTVjnCC+YZr4xsbjf/IQR6cNSCqm5lsb/JN
oebMyEUpcmbZ745vPahiv4AwyBoN2WlVHDAKaLc44nE4fwC4wFvyGsbrwWpInshd
vraNLHFOH8ohizDfMPfrQmvsLgraW2wDDO411gb40FyWXXabtoxq/3ume7Yg80Ke
UvUB9XmhgLkpKIBDDIjiH2b4eNLTjywdFfCssCN/TTsiFWE6kH5xMkeMgTLC9w1W
/ay10VCwCbcX5Yp9LVJutADWzlfoeB7yIS/e6zyLiI4taaAAdkx4UCM2z/emRjD9
jy6gkSQhwTQLvaWex5MyqKNIOJJCm+QM2NJnM6BQH/OmoTBhG9s7x8SDHnsLjJKQ
Rl69JNGMr6Fs8K0u5X+to5N5uRsQlPgYh6FK3wZpL2cr1lGGXSEIRsE1yczwY5CT
1WPC0+ilClGt7zdyw4xP7oVwFby2iZyolGo5pI2ZVKVHxoctd0BhZs2lYK/oH1/E
m2S6UGbLphMIVHl05w2dQEfAlgHs3wwOocs4rb94aeoSynO1YyuZq59z5wNwPTRv
DwK76avQTDOc4tsaCAN9E/4NYyqwBZaB7k9xrQ2wWBj/zLDVRDAcRXPRqUvMzRQ9
HYa2+NZNkv+MoMryfVD0B7JNgcNHpAS8sAKU5B1uZ5daM88n/ZspQn3265k2Rc46
Uw1iX43i3Qvs6LN0Wh0IfA7qMfwFywOYP6mCUcCAsZxvmyUjo8YU9bHfcviOcUaj
mDWFnEaOUXLWrt58lkWEaMyyHm16peVCr/Asqr5aczyg6hT2IE3US34KaI3hPcP/
vC4B6LQV3xuK/iNYfzEDBGV2Bh0v9XNSoWUu9sV7cilMcGHvyCklejkjNU4F6tqE
HrMn5dVhFTzd772TwIitWUVMxcABBKFcFsD+8q+nF1+ZYNS0ftG6dSaAlevwcCRc
3tKbZcSpf25nFJLBZq2PREVOZQ+E5nHO3A5dDg8w4BkerrqVzUWg7LQ5PBU3eOyH
yra7w2HurS3i6XxtlBMiOla8brT/43SOHiOdX9eDEJ3cBigUSsAbMcPm3mYl56UT
YqCQLKTPPWX5IpulMbjaRwU9jE6sUb0qvbTRd9NAabnzqopVvI83Eb4XoJEb2D9s
J63FwA4UtXXYh3FCl1ZY+QkU63cN2acoK1tNe4uB+dKop0VRnAZvuJfOR4MmNUQw
0t+7T1ROm02J2xuIWjbqzfYX1EkgLJNqgNnWxg0JHb3TWbK/3Y9/pEY2hGzbMeMk
WW5QK5kaX6GrD9BJUCdw75oUnwFSOyKepUgE2qT7DGpX8CJdijvwe+ATpjfe8eJD
7HZe7QSoI+1cZm3skrhiIoEZ/PkH635pF3b4at/bpjLtw9v+W/QYAKU9FJEbFl8d
ApreRqM0dTs+wUiDNhcUmPYnBul9O5xUkS4/syzwwgRfnv8CFrNvrGoDqAE9Wm8z
YImuGcD5IOGWyz87aT/RI3b22aUTbAatGaOTNQqyqdbDdBZNzRTVOAMBTyc4Y69j
ybjL5OSe48uLyavM7uzjqODmwx+cha4+Xhr+EUFag9zTb8nJvLdXDSyxC7XbEA3r
rWd781U16w/Uj7Upx7qULyPZS2RIgkb+1C0cQYxsnBXxoMMfAq8JVTlRYxaKoBgt
O1zOIVlA9gSXOTAf2OezP5EfsQ3QdozkvlMqMIxEK0m5FPy+dzVKpudTvPh5/I+g
1mUK0oG3vM7wDxcRid8BJi68e0UbOHHZu1R65pPLGOXnTKytR3icPlc+0jzGZBtR
jL82NCUYTY03PqG3A0MpbPOawpOfpTFAuzU2N7S6vkee1LCVnEG+0tfkakqiZLCY
6J4bpoCQWm5VkEY+uY3P7nvQlmmBletmsyYksUVt5JH8Z2oCUoSjwQCEPzUY4RY+
tZpdJqxOaMgpgabQb4Zza5Wp7RKZMHej+Jz/NIhUpDOWJN91hEF3d2i0oV6LHtJx
sbnjfeOiMXtYepiOaH/wFKCSZ3tav7NfIpK2XqHZ7pcT24HpZ7VgSFwVlE6QJFNE
lu9pwiFN2pjA6kaU2aQ6NV0YZWQ7X/U4hqw/Ag6PtTQDg+ml3g5Khx0m+RLL+r0k
eaRD9WizG+MEUeyXeppp6IGzSwVINNcpZMAnvykb7cUhnXoZ5UopTKeRftVy7CG0
MbeSN/ZJtAZTYkD9RBA4bY/KyGRiJr+qtx8w4Qvbk4/030J3OPE+fcIwkHREmZML
XEwj58HLRN9A+CMwJp0jUiysxZ2TkqmbjakI5adeXXwiagxiX8ovCYBPW0yjCL0r
KZ1KGvpz4ud4sekKLkSmnVKT8CFDvh2ww/N0KPuT8heFMJin9isT9G/hUh0orrgQ
17tVCY95Z7bGLcOM4yiS7R6yKKTnZ1l9Baf2SoHr/yNWBc5HOy0zqHhAoQEExqWU
kqJE0GecHBb44NQVLek4Gq5BQh3idYXtIPHgs6mcz3faEIXQo2yMuFHT1GNEnVdr
yzkhR9f/qxXJgmDh5TsSRK4wMrVQldt+t3P/vcriBCQ2fCc0s4ST8cIK15+5Mgtk
tMENKf1DfmsDxyt/AYywA4Nx+52nPFyHGeEdMHMxFJB3pHp56OC0qmcr4KjK1zo9
D+iOB/JUuQn0PtpNSRQjP3ABN9sp32uWhJ24N4T2x1lBatEiUVJSa6Ecm13Nh8ae
X4DTSkWICMzK/VLsMdZMksfQ/JKfLGEtzmWFeFlmV8i3cuIbLtA4ZfdrlK4wTsaf
l9Go4UpPte5MeZ5VgX+Wo/EWeJhIxLk73a0wX9KjhzVC+8PjzvKuJH0j6uzzpIOe
+EFrQ8IY+455g7XukqCCsEjx/Z7NzsBSsQulWentRMl239r74BCwASyNb5f5C2IQ
fPnPx2iE2PsNT5hcjqb+OvdL+LskVcooM3zjX3dQ9WksxvprmPcdTdNrfHZ459Dn
O7w8eoA3sqEaU++g8cRX1FF5aPWuMYYmtEFl3a+Fhf1HArERBYl5rbenNlMvOG/S
n3z6w8I7rb8g3CULxi6QsNRMqJybcoIIiDL2y4l+BYT5e2VwBQcxzKrCwKM72w8P
XbqmlpjcBOa0M+HYwdVJR7o0pqQZp0XJe4CGjihSpFhDXMRWclfq+KKxx+9Af/kC
iDgluix8B79o9WBz7CKSPEz4hlOWes7jn4lF9AH4I96D7RxVqoMaap1gsNw40Bd5
Y8DiiDjOcYr6N1r1yoTmshCKW/uVdY9vIiaOczl3WwwH9Dx2HA2vqV4ILjC4kR9y
8S4dNYvVbfcrC8xivUkM64um71VxqYDNZ2Tst7XS3KLVbd+OiE6SQb6Q5iRhd6/F
dwD8joPhytwF+alx4Bttdc2MgLNOj5wWpolyngou71R35I8tGno6VYI+jyP7ea91
OaEaUnqNFYahLt4V+lhIl5dLPkqbnnGkX9I2w2x4VJbX22K0UXHg3M1clSEK3clK
44zE0sA+iCXmAWmLIWJ/+wsMrXnN7verzvsJm7WRoJuLjm0SmJMkUjm0xn8SlMBk
9eszTcfRFWklq+6L6CjLxPvcNlc+t6OYjfOsXtm5zuokGMBgV3mKLUd8ISWtk3Je
+P/bOvx997T18JRc64R0vQed9nsretvs2LfrezG4F/mOA+6rRRxQKgMOZ5SYC2VP
0CHhptJENm8pX+90UDNiHQb3YAVNg985L5nASgheWthnfEOhf9H2FWM6mUpIil/l
tX9Dm9T/lmylowGijCyyRAapd4SDku/3SzMPaUNvRA/a2opx3E1OhwSPgw+V0KeM
Ud3Uktg6QjWSqM/+g2p90a1qiqaUcOWmAGQ2DAiZqG1DLAVHJLxkIO/eqZTcjqcl
buBDxQFcxKxPWSq4ZLYZTGkWXJhwDrQHNJZNFAFhonvJNWI+wfq4DAmSJtOhITaO
gGbJvfhr80wrKFpjG9DyzoQAOir8WkQIIN4WDUk4X8q6rk3WLcjk2mLY4vH0zYGx
xfvNrkJlwTZKEubS0Tl5bjAviM+Yiccme5lDJdyfDW6KfG/xzlLQzymZc3/MM3n+
bajyyAO1b/9eT+gnWNjkBbBcVtSE8Pk/A1Q3lr7z9u0s/xsYE0IYP5HXKR47f9XA
skW7jPGIgRTa0+3vzORZhHl47bsSp+bLkvyD6tW16BZzemgqovHTBoUjGREYkq4n
RQtKDuAioiPMxW9FZ2oOONjusIKdm4s3FfV5L0UeU0d6UmnKJ3oRwpiJ9B61aJ0U
RcUkYGZjsoRkenXscsFAFh36rF3jGTftB2VB05N2IWvwCHPmibKPROD6qesHntPk
qiO6BkXeaznoKvPDJSHHHgoU6/d2PkPX4Fska28Ypw4QhGvyEHz4QqNOb4Bp+Y7J
ik+AePKZHoSOr0kb2x+pmagp8HKSNg5Be60qFTkLpcwU/qTyGr2Msuu/43zRMSUo
YMaBvn1CBdc/eqvM50DA2Y08OaEPtl3t3HNEzhQ5fm1FuXz0tsbp2N2roaTULuY9
Im81stxb/AtSRza5Vfwr+t8ELTXsHHlJu1yqTUR7mnh1kAdSNiKq1sqqOJxfD+/I
jBYO8yMHiG2TT1q1jkA6FJPhBymdg+I0hPXIlIGLpcqngtMQn90qPIQyZOig0SfM
wqRxOjTQR7vTCankXFaLEF13QiFJndyKf3r4O5GRhnKbWdHJHGKnvQ7i+lO7Nz25
Am3/Z0iygft2slDXqZ31AphjT3kyrRQdTLR4u1nyosz03p8RP985skOMp9JHvaSx
TDq04Xn+TxuHr+5UD8t20DMkJ32TZO3hpYKG+7oaa/s8pl8ATVsgxWuSBXiLGRHU
YVDgUqF496IzpuvadwSDftyx7/vanFyrmg0TUkn5/yYjZ/dzLZ01ksEasmweI4Qx
NrWR7NjPO52h8xdwc3FSKhObWBtho6uKh/PTejK5mDOhq6vZYu8G2MbqKMo9C7M6
M5+K/pGSVx4egBvSA0uI9e9eklGLXZx6QgnCZHMpANxfMeTZZFDEGi3OebjM9b30
CpTR9IkmeRAj1wOxW+tjdRdGXfJmLfvxzyvuRFvwum7rLgi4xdS/FCjY0+tGey6I
F/IKepv1bjw0s2worIIybdm1Bs/YKhfmwDmhZ3MCv0lpRJMKuEI+N9lPfGABis16
yVpINPSoSjFAyftcEmvJIVGHrot23mgI1H3weTln7D2OAJwgtYlswes6jyYbXQAy
1d2/G9QAosCMih7TKok6ge4v9cBIxnmNjvjJMcthZQlyPW3OfiNpuO0f0MH3wo0b
8yUhst8NJeVxSmKy6KHWi2mV0L568sTuiqjGPLeIXllAfBsVt7FyVY+lhHIzuHbF
uVRgcXp1Jm6kg5ZYMMblLFnMVfVZRNzFjlOdIrl3Th4C0uUdFMY1AlLAqsS6GcKv
ozOfQn22VHPb4JTOwX3lFOEOtQSjA8jWC3kmyx/VkE5qn0vf2V2M/9CizSWmS+Rp
fTIIDH+YFwF3Bl33oPxHP/3l4Tznh98S8j1LugLKk2hTariF4xt+DdPjOVo8snkC
DkqNPRIz+WRJHWUG93fv1wkOqx933n5NL188/zu1GxLoYUQIAoOE6ugreFLZBMdC
ipxdF6pm9RIwQNZnMs1szX1B4Z6UbkSIW1+RsH/2nN85/up8fUo2eiljoEpLQIVs
3UX5YjIAyd75y8DOpNpietfv42uzxwAuQ+DY3Y+lJSblVqI6aFos/vwxlVqyVCss
CEZ5ADbFM5aITqqwrZQ5FyJ0OR5l4wENq6bGpJwsZhgPUCwBlVsJVvLxBArfmi3q
6qBm8dhge6f53z4KSU4jxlt22idUUddnDQHKJ/i9ZUfB951nJuU42bb8QcEhbBOm
itxjZWSAtsMTcTMDRR8jhMbdmv5G74zXqiMWAXeJBhV0PaAhGUumtMH3ZY7wJ6It
cCqu6IQ3bk4753RUzzP0HZxic7eoEgTndK68HMNiD5mE4dmdLciq2F/TtBE9EXbd
kZ/ougF3IoEDwZpkF5JTXM2ynAsqyAZmo28X7RdcuSwfEVMyLLNInj2pdY3yi/9z
vbt8PTrrpePei+fveUCb2u+mGE0ZBoZko2XpBQLHIZV78VUjTYj3urHmp2+8WeBA
Y7szxrbjyRotBXr54Ut02i2GJn7s+6+LKtHlKYsXZErxog1WMrzxR2T3r9K60w6x
+UermKXTGk/t8+LTMBA774y6A8kCy7hwZ3bvkwyGmWjnIaW9Yv6SVEYapkD8X24h
T6UsWouEFW1ISal74gsCHF7ZPBBWe8nDIUY+EotXj1zX1laTLr131MVwswO9GLYv
f32Nxjp9Tq7AthJOKZBBA7HJbmzkZ3HmDkkmSF76bUopdvLCZGlrq4x55XVNwIQ0
Nm2hBiQdIKNRACVz4cedV4wfw/rC6wTnUPg9OrXPoRDA1Sz6cpagsmwR4ofxVFPk
IRaojB2H8gZoevp90VplIE0CZ10mt82rLuXnZtZu1DeleCK5QzPhkyVkfpKa2cmp
CE8FReH/LjbfrbKwyqRg7RQUAILC5FnLN71IeJzX9oUPu5Wn+UfvMy3DdYljLKLe
Id2/DX5RckrxUkfcV/lXEGduLDImwBYtlRZEqfqDhZ0fK0NLV/DT5uBOyQUPxl1X
yjjlNV8kmtkUzctRmJ7I116I7+XkzNSIM3C059nem29tnRSq5ID3euxsIAs9FUxT
sQXsiosfqmaLIfLNRN33jbqm4gOGBGa3KMHPjYeQmDhEYqa0v9p6AwXRBftZcCwI
LpC5g5tYWtJt5/hWhgqZCLW7jmFL77ijyoY3LV9HvDKgd1/uC6sI8nGQ9qirivsz
FBLuaJFTGNxgBPf1xqwKpw+c0Y+oisS9Gzw9xmnUyAWr9cPbCJUz86ly9fnqgJiM
MNWUQJ5MZz6Tzr61D9OuJzO6yy/tg/Tu/23TRpsQH4iJgvTkOswH+rfLZzWW93pa
/TNvieyL5ZAkUsXqcRpI3cTU+kUN0Q4Tpl0UNS2aySfGOnAxDFtuVcsQH0WHRf90
HY6u5upThenwfSLv1NTa7j23xHcSbKr7POnNCExsa4EytYUCfrOhtpv8OKGSI/94
gw9EHlSmrKu+F6UarjUGs7EWm2lg03E4kNqskIOsCFGwegn6oBs8u/7msoTJU2OU
TjJjlsxYU3KxTSznJSwqKz6xhQ7Dls2Q0bYAo8RLNaqcROPRl3yT08uRePIXORBg
xyqVtEcEKVEfOoEkzLpyVx6q7/nYhlQF57PlYl1lvh7dBKATDDUAJ+fqFnROfk6t
s5//piUMRLZQXgCUFSyhUolKT7immsgAYcTpVW80/Q93l9IAM2eSjXiZ/khOKMI3
DZAcqh6Y8XbkZ1qAJxTcTx3WU3faO9i+zLNmYprhFmVyCWaH0s87p/EEO5aTawlN
m/6sD4Fw5OOilVnuI9Eb8GopPiK0OpUO5L6pR0nrWmvbv6JGhcu5qnKwnNtJf+83
fnB6vLWKlqLGdjDF9JBHsNiMSIvc1FIP3evOFyHlVC0leXNgzmNWN28CjTH0xNfm
cAVvQPlFA8D8ZHBFU4NDiw5Uafu58DNMaKVyWND/ZEhg0Nt91RQE9fpOVuf4Z7GN
HSDrZad8BfGHndRZZ7fnSy/Zp3Cgw8h1MirDwjBSkQocXeDjxL0ARm3vRHcvXUss
nZPQojJox4jKQu3VDZo/SnHjTqgjoOtrmU2stpM+uqo/nIUbqaOOlG7ltRDk7LVh
NfKlm4RKnK7v8AqMCDuuuOsPuxLrbcERTPDtR8x2twcwwbUXqu7M7Gcnx5fJmMrz
v8RKVEhodGZLNASNp+s5Vap19/e5Gqp7tfaKZ9yUHa9kCIsDFV9wzgEvm7kE/QTo
g8yDsN+BhSd1HX25X+6layfr0fj3p8y68iaSxGbkuvWUHjqNvTG4wqpll2HliEnb
mddx9XfxZxc3WewqySIjpbSzbcDWqn8dLW3SWJLdpPupvcBoOfS0ePQ3RolItlvq
veZB8zMxjs4NdUpZ5KiLF3zadi5pq8ShKIE/W3ij2k1XRDG4g9XF9jwYjfL/PcSX
C9bBAWSFXKOesF+gG2MOTUPlXA15q+tO9/0ufsMMSLI1VdonOnxbhc7X8+Ul8GI/
jUM0s9kzss5Q5NAzgdAJRu2YSpiukMxy6ALP5fWWbb93G+60B0ql8rop0pT4DnO7
KyDVyJkn+FUr5edLmGVqGFgkkBLi7tNPmwqgm+cAGoVCc/1HajZiZJlZBzvro1Vk
u75UAXHdIYUyV7sZdpH/rk2iOPor2w5eFfasTIcaWqPJxq5OwKWeNnN8905glq9R
Xl+co+vFVTS3ZPzqKKomcmJhyFOB0PBICQiKwnPH5L57BWch8kDQsUo9Qe5/kKQp
f2SxpQaTMJ38PKo3RTOfdimtgjYzvoP/voE+Dto1BPf83iS6+eg01pQImQBIugdZ
IO2omxVHUkw8n3fAcv9XXK3NblGJ+YamWn72bm1fvDLyPfLUuZFUjolZghDjSmHk
XRz4YjoNaUODsCsTMPs2aNzN0PPCVgAYp3bbugxN1sBu4NvJwtWeEWgh7yAJr9kI
ol98gGNj95BzjiNKhW1f/I7GLTki5jrhFSem4Hn/NG6NhXwAtYc+fhPnIqHIjwl9
cw8U1e8A9FZxxzJ1CDcfCtK9t7p8jRo6ByjJMeVUMTmO8eEiBtgwZVrttIIX1DXK
sG1yIutCSfzwFHutsgqieYY5ghXHU3nmIZ6Vt7RoXR7m2QscbxKv03mZ3QdTJc6y
le6cCcTBNOGYTmbqTr10gC1pVWgvMUU/+QsVX1thiz2KcfGWb6g5SmNurDzIrR+m
eRlz08zlT65oEayw/T33scOB1SSbm/4LPwfNx6rL2HxwigrqjMAnispNT6HYrYJw
4E5A29Sf2WJQjl2iBR+N5bLfPOeo3NTHz5XdMFF85wcMB63T/VhJbIsmGHy40ZkC
Gy94eYRLG7SNF5MftQ0Xkdcw0+GHm0jUcOe/SHjVWV4k4s4SYJicbVel0PwbArwW
TTtnLKoxyIkMnQhEUK5FhdPHjnZj3gnHSTaFQzNJpyPqKk9VqDsYMj0fMde18gmm
c0GQtuN3JcC+v73SX25x+xsTN4YuON+PZBw2ysgVi96OkMvPOO9mbVE14FeNvmAM
X3Uj3hPb5OPsKCWooum5zNBSkhZ97kfT6kIjkGkoEqDEFIjaOikX5N/INiI9RrZV
X/xcWz9pX8VSGyXnvld+Vpba/TBKKasDrkuqU8mZxNbvD5kJ/If2d/FOrKzZrPd0
C8Bc97y7cCsiyIhsSSREriEIeic7khbwemkDwIUFRdqzokzz0et8w5TNxPFVDQnC
qh0nNxY7j2CdE4CxhMOEnYMSjjxpgiEALb09bFzzjuZs49bBz+gtqE9kEgY87Krp
8mt6J+Zyex92CGnceCgLKSBBOAmbZeJEKtSsYWe4Ef4Mrja1uAnrBhdRYPDKCvmt
HPpkROFbNprgHE8B8AkREuJ0spsGELB+w9C3xWbpzLAX7uIwtohT/jD8E+3VsvTg
m40JwFKuLlrmCxnNUnMQlQVSqkz1L9g+Q4Y2SuMcl0BYsEdyacFgK4FBMejwyupD
oh5CR7MZQl1CP6EOJHvf20MFsbMDq36K/drKG+6OKpJVIF13G1HavTrAmj/khqwn
+tVt4hkOj6EadSVLldy3R+mXShFFVqLPNPuMTfh5II/Fq0d23arcj2EF+MrT7XqG
loTwqOVVR8YVNLkPbWRXvmYk5CsXhocKwePxVQbKwCF0+2kOqqNNeyIqH1U75v6T
oaCjkPgpyGVhjVlyPdYhJjdo2iyrovMg7kjw6ACM9WcCmZrsYU7gJTeKUVXbfKkt
Uj/Gij/eamoRjwv2FLa7BZz/eBKa/aJ5PKi7O2JhSp99Iq695mEK2A8Cl0Gj3jVm
NchExtRiNVnZNcJuxswCADE+sguHdBWlNAZrkVsHK/7/TWHcnJMeNHH/QcO4tgIY
hdQPsV+kdTn6NRtNytyR1OcDBskM8igJLYBtiW849cmIG9LckFMh1sGqAu7sL3hT
QtKFVwsn3VvZjn0ZYDCfvTQOEKOvzKfUqLY8RNNj9S/+cZ2ak9DMaREcXnorGjg1
kKj4NJFBC4BGlChzbPYlG97qxYD5lZllXmYMm2TOmdr5Ait+zgiJyNBBMb3N42Tp
SJmOzaFJyf1EtnQD6w91L78YfkmHuYQOEibdckZoGenSbr6FSIZnLGiUAcp29Jts
704YRa8TqvvNpLpHx6Rmw8S1ZyXW48z/MG+E6jSPSv7doe5S3VWlgvooo/BkTq8U
7yfpJfrGGwp4OCkurqI8gsXAIASCC6z6dCZSBbvqHbGBb3P0LsuMhTE4KxSBAW0j
Nsdn5hkezpY03SAD682rCjKT9ypx278+eIRNambf+KMEC0fPhjv7zyJNKPLHTS5p
ZqC/6YNULuYlqyOeh+H32oGJfRnxune9g8JmdGxWBq60V7A9BO8P4C1E4k98iNtO
vuodo1vVsyw8bp+05TslVLpURDP4r4Eyh7fOHS3WQ2+cZRnA1ENek1oonz5T7zW9
K1XoM2yWpRN/MC4qvYfBNpAay+0yZCTvJwc/ba2dlXJrGcM1Kfv2eati4ItRtx57
e6KhB9ZsCXDhKsdFq+zBwMQNe+2AB9ECMf2dbf3O1y52DUdWoaRs31gE7lp9KsEG
SO0mAsjxeVH3buvBTprt4jKx9m564JcZPVwSl/m7ulhQewpAE0M1HkLZaQkIupc6
gINCHAEN09yj3bAQaT1ocpza/48mwpt8ZICmzxJr4eA5kyeSEuQVlejIyEJiPhzn
Ockxn4VdwIVGMv6wPghvocTuVRl4s8/+HQVeicSPMQzrIpG7bddDst9LVUldj3yd
0PgjyV6iofDjVJ2CP+GXEX+ztanhVo0Zid/RJXBgQSyfJg6cCADaNilwGIR9LPzf
fpbgsvRDephtG2dBM57a2oXw2TWmKpvHF01nG8vImBjUaDhKI/k5sGeocabxYaNw
r3JWXD5Z8z51T/TLu99LPljaGCGAVqAXMFE8Vxclj/8Ve/1lw/kBokCu4KhnZ+RE
sGSv0LgSyNge6FpWXTODtRSJwzfyoBjEIwNQtKfn1UwwQ3mbVLvxzoO9vXsOecfR
eviMRBMeogOVrkvAG5DEDi/qHau2DzFqO5Fp9UHuShBcdW3nWNyEjKdpEtYOUspH
cJFpNa/QwGYmqoqJoROjux0BaqxqWWgit1BdxxKH/ZKUQp/Wp2lGczCwuqf0W87d
AKvHUkez1bXbTRk2777WKJ+Yr43SS4b2siYMfDx7TUpAOCaYSIa2E+tAhikm6ssD
Ee3+7nG2D81JN1ROO0CkI919yO+2SPE7MQOV/oMyHTdJ7IBuaF43pIX1ZiiCBkYK
fldF6BbrvX3BPBnkJXCz5owMrlNZDf8s/QtFzjiUigEiGXVHMiGv6fNKvAxt5SA+
CE7KzY/hiyjXu/FbqTG00rRAI/jJqMYuB8Fb9jLLAcQ/1LciiN7JOxqkM4cDlcZ8
Aw/9DXKnGq1IQthUK5aFYe0qZUOj1YgIhHdcEOYNsrsHiEf9ctXbM8NalAX07+s8
SL+dddgx5gOGxxlxRKSvxih/to0FM/qXDVlgypsGBCkXyGiPiOZ80I/0VG1HjPRb
V/bxrfGaqy3/rohJYjsXjmobsG+kiYgeDtyCzkvaiJW5luxNzePem68yMBX0W5Qh
t37mhn0YPL7i8op+jVNjHsMmfBdTDWeeFCRATnpKE3C7OG2iY5SFzDkjoJR0ms1h
SilVM9+2U6FFapPOETVOtZCW5nxuxO8BySRc4vT0okxPr5rMtfa+cusCW/WhAvCn
T6jLEODi2mJkBoVGkoDXPBRY3TzpdzF8J97vhUm810I07QKGo989/6QbFHFxHzpq
MZBRlgvg/QFeZPVjD2xP2H18O72ICnNRiIhvk7kHGPBkVDqVF2O32ZG7cAvSw9ZK
OAyIXyS7bAtyfB2GAF/X1VnirZJTUWaR1BWVy+gtSgiSBzMI7yLRfRNjaWF88/mp
OOLgRQnK0oFzB83+A9D8boscfgBs338e3wfJsCAvqoJyox5G7HGjvHpEJFFV6VqG
cz4aBs4dtIVxVuTufQBwAQz6huIy+WIIiIPlzkrqnsr9HS1+DGbNraxPqc9ajzJE
WWO1EkB3YaRSPTwRajhWuVLTEohJ8K0DYogPCyA1QUt5HH5uJimc+do+WjEZykf4
34HKgKkbalDuXn6qJ0q8CzsU2RnDZgzKMPH16jAo/sX4b7Wr5egRyqTkO0o8oZN0
5utZSXyhHNvh8fLsikf6P/A/4ouHqxTDVb3iKqKXvLO3vHWktw7BxuXLoHvfBH+M
KuDfFq19MF3Dhdv0j7TNBZig3Y31pdNC5H/wUMzZ+vQx943FRicJlF6S/haxrjCU
pLsM+YDQNPCwxzOXQFIUZYScEKJfBe4E7H8nh1anhyt80LPMT3qO02PNDwG4kkrF
R1kZhNPTpNPWZK4gbhfBzd1w4LVin2jAMt45+tzVNntSzIT6l4VwMnP6ZCuQvxJg
fAqZghkjTWO26MLOVliV0r78KmiKzbFmt5r2A8wKLkdnQ8LuHKY1ztkh4k8VNBa0
5bStBFAyOY+g4G7LzfBhqYLpCiOSLgkWw02WV8ukOX6jh4gSmOPPW9PHVoV4KuGJ
6MdPep+WxB8GJVwn151fNlkjN9IPrdmtKKrnRfCDfZKFnDUOH9M5R+qacbxfsOZA
MEACNXVyDyPqqML+o41KoUePKeuAUAwjXAdUkuFertntwU1HqRErxofGZ/TJZdGc
9yWyeP0D8i2mSq4hfZRBnarduhy+AWLNP1SnCgGbz6pt9jxQc6cgNFcEaxIwo6FV
EpgQfoS0KEMRYx+4VecQdCfXXIvkMQeIiqn/izT/eknm3cQJQHWpowiw0sLF1a4v
YWdzSQPUKMOQPBMoKBKNXDzaI8KOGcTZb3Cth3EEnaloeBZCIeNKBOz5mIX237h2
ZcYx03IZZ4aCDvurOza/rNEgmel8/j7CmAlyT4wKDJ7EPYoTL7trhrsclj6oEQQ8
XHhJdzsSJo8pewfyNb3mdkPgdQgQ16QPDL7NDQUX9+2a95uGCLAPml7rhHWHsPqB
0JVVgUdV2LCR10mZRZ35vxpcVHRJNjAStmp0WGBVVhIoeOzcK5sgpZwgnuozdJY4
Zm5R7PmtP1snPmJxqzZoyVRPEZ97F27euiP/9Owed9aRaD/j2HaSTJumnpaNzMlb
+ahvtEg929HPv82p1Ue3cF8JJ4JIPFFIjRO2v7MdG81pBXtgxbMWJ5nUe7Lf5TT9
mHsEgfpV79YUnPoiEXyAzemCLYSwZSMUbYgXXC6+ZSGqQz7YwfJf6wSxSccrQhXr
D4f+RxNlUFTie5X9SZldOcemnM6uHy7THz8r5oGrBwdoBhQ5NqNHH3WeUthm6hxw
bpc6MOP7rCY/TUXnd/XDJtn5HNpQoBxhxMjMfT71DPNl2spYia53aBEBSHTC574s
jTWE7DGltvEujA5heH65yGmLcsgP9AoHZrxqyQDMjLmIiRC51G5Li+wEFq4FvmYU
ud2zPSpM6egfhi02aLsENXMnks/SqzFkdFsmcXEO0xNGbY7CtJHRj3itKLnHHX+w
yCdUkvQFsFMMlWdAdiY98QDoBpAhVz1HDFq3hrrFGLqzfETtmKXbIX5ypngnbSQY
l3gLPnOPFEFAREojUWScUeSZhzzlQnCskiOxNi0m59BxS65Ixfk5FGSyPJV67dIL
8QWpi0a0xJaIftLykNSdth4tr91X/hu5fESmjmyLTG+4tj+xCc1KsnFypCzKVbz4
GL9Qlx4YLTWxRZp6+Nou6KZv2kcM25cgNXIWzRkcksSi+ZFjgL1RMunmuMdEq2Ug
nF4LvE2qAhytm6VbJWVNCB07Tn+eqjwKKHQAVaoKJCvxh1ctKT4oT/INgSXy1Uak
2QvNXXs2n9qozJWF5mucap4yOf5IOhwoCXgrNByX9ZD33VAzx+YZupbTmVP955Wl
niU//laFlhDOkj915GcPxoRlud8aHS+lBPk/wO9RfG1t58RRxNKkPZr3nNQIesvY
uGDrh3vavqmq6/+IB9GN3/QEz54ZP5ZT3g8X/EpikrFqhhdPKqat61tV7U3CjEWt
Nb2J8pa77YyGBI6/inLMdgDfuVSColQcVExgAt7XkDIBiiyI4NN2SsMi5prup99B
62NBTUCu6E99aHTzoPQsl6o3H4k8pi1MJ0imi5vEDR7D2N01x6jjGGnPIr+m/o/E
uEM9jufnmGp8S7MOyVEsri7InFpEpyWNQblaoeCmXydwNJNauHFUJoj2n7vlmJcA
dJRj5kJ+Et+KfZgZTHKNGcvKVwQW/CwEy/KM2vyBDOF5WTziY89jnKAqbdJT8+nf
v6gZrJmfJ9yt/HU7CNTx3E5oCq9sT+qCZ706tV9dJo9ekMfPvVJX8He9DGpdABsW
pGuKCSY5CK+p4DWjAVTicVQlwC052p2JRAKeL/KegkDUXeF2P7++Vil5mz116wOF
B/ZSC78Ijt93L8ubfVDBEBa1EvIhpw6Tf9HerPaIDNlm0yTBLQ/4N2hx5AHbi2IO
oU8tyH/Nm/LyI+ZK17ESZ+a846bfYXxGJZjjzHsLBZY0/fACsg+mgL2TuaVaYBc4
4EsbaofCly84bZWlI/VOr99xneRPAV8B9UuUJICF+dx8mlDFZn1ykCIOYRDo4eQY
vFJs5hAH28QQejRxCIqFoRuAgsJDtuzbqx/bFI0tDYdweAdlC9+jgF9dEUZN6wt2
3WGas/6cpRGggb7QmYB5xkAs2kmF13yNIQ1uzYpC8K9FC/JFLOYHNaqDV6mbmnZk
XXXljhbfHiILqQFhWK23mjfMxnfFM+fcJuCZrs311Mlo28uKmcI3B37MrQ0cjSdz
H55Z9vzIqWJXAAPTHeKW39kBUSDK6uMzsLWPrPnktUIJMx/0z0q9DtXiSTHiIbEd
/YkZ1n15MSPumqLPY1PMsHTcrOT6eTeHdVIy1mKKPzgVEBD4JZQVglIbTcy+Rub4
sWZ8PadevctQXVckE+mcqavdAzzbeK5WTSQrzSv2h3tMfRNRKb3KVAiJaU4CTa23
H50QGyBmKuGLSbyWyUTV3TmBuCJZc9E/G927xf8VKbAmMhtM+QjuhKBAoYNMB8eV
1n+dwY1C9aj0Uba58UKuepUcGtcen30a4dr1MHS7d2Bvu3V+OW3+jFPzGuDUAnry
/M8rgECGd1GA2Pz9Nm5giQa8HZeTJEJyp2TN/PALTuM1g29h6pAgx3sInY9Yo/tL
fUhcmiOOYXaRIidtYT8FYvrt/UtbQou9c/5a53PCwalsyRLGLjVK/YBkCbzl/6Dv
3KiaEtsL0aISthmDJFUCoPNn8S1WNfXh6G/zrW3CS4YYUiPsZTPW8cwv1DHgViGG
6nayJFFjLe9pmOlYyoI7VB3Ofic7hJswbRhUQS0hqNP9f9FPxPFZDrZFbL7szDnT
ZK2Tz2c2X7DFF0DkcVyi1nY+UihlmQ1XdqWS9DRE+t9MmZmPLKbvOo5wEfGgC5l4
BlVTu01HosrZru9kvjN82hWPJ0OSglMJUJlHA/DeHR1bocdYwhYsNy/db6dC7MPa
/1b1l+S8Nz11JTF5PbM89TOcfEpIa9E2JDO7CIe11JUAuH7QorZ2YKZH9kvvo4PD
l1XpUYflsrRqeBxjx8v/K9uOZtgACS+yoG1htz15sYzuohtivJgI5U4RC3V5An1O
lsxOuCNJa8X3DejnpauOfmHl0d093+XhvlNmIzxGyWJc+2w5CPM6TMDkspOwZ/Nv
tnm/92uz82iXJGJpvnwLQ9ktmp2LH4VN3fGpOB/uqYSIqvYQV3s6GtBInEXDgE06
W0FlNV1kV/mVZmVoWVFzuYoldIwBk5u1r7kxVy50OET1+db0MqUPANRPS0udWHSH
HtcsKOphnw4DzfMdnsRdGjPg5/N3574rkdPRBgLTbMnFATgjXbc+kmuUPxOQKoZ6
dKWSR1corA1pe/OOoG8v8hgPA1GH3vpona0Okvwf3r1RCK3DuxLor7cyJih987JR
LW8M8MaM27NR4iYb8XRtzdo4d0RzVc89JL103vGK51w5/QD+CFsmMuSKX6Q1Xr6J
oO0OSFh9QzgHozF6/D/+/5C3MXPPmPupkhEIBUGILiwDbe9CrzmVccrK+cVkTsZ9
3imXvVX/q5ukdArHeOx+YOExu9sEw6pIFNaze4TDojLXS39WN2yNHl2WluhKcXlj
Jed1Oej5LpjB6rvzM01GbedY3xcpIr1Y9SCUdnAhMRhimu4K+NQBmpCSrTGwDlgB
CZT57Oj7xc7YDcRpjwCWRjLb84uFT1amuQKnVB+Z89CDuEYnIfSjm1iiF8HgZenn
JYfP3PonlpmmLP5TX5zPEoKGi63VPoNPAUkfkNNavJkDX3IkazYin6XFRpA6FF1b
Wnm9Vo/IiSz11OzDZSNASMx29Kwvn655r7fhrUYHeF8I4j3CQjRZEGtBryAylewI
SjCHXuGj4eoJpYiCPPfX8iWTVbDcahpGuOwtIAgcl5YXcUTnQ1/Pz+G2ANFYKnZ/
SHIxLy5HaiGnvUQHEWQi7LS6JmAGpx37riwG34Pl9BpyRJ0DBhWdnPdoKSBY31nY
o96eGiE8jC+esE0Ko42B58lI3/C467spYcPd8jW7wrdENEO0Lh911gSPi1Ece2gY
YVFY2rjlWsv6hjdM3uBmYl1B4+BqER8kCDmD5M1SF62Csh8Px+WfQuPyCacxXJBD
J7Xy7Rr8SInIfoF3wQi/gIcaMQda9O+Zzb1BxMn/ByKcifarLd4DWuuB636KBbUA
KywLZuYBh2/DIg8N99Dj4anqtyC5BK/0WxlnCmJmdZtd1X/QybsCVg7AQZJD08KL
f7OnTAsCo2G9jVQz5dhRtGUbTncgmgX2kDoH5JdYqK0PzIcnaegoAjF1hju3Sqwo
tfHLgv8sTVGIA93HnntG3W5wllrgfqNcuxxPcSc4vK43iTfasWFJmbKByTu35rfp
SQGvpCXygOH54iHLJ/pAuLqKGc5rtTnhhEoULabFhGEQ2cDyZ+9qjq8jDRTYx/kd
+/EEek+ea/yuEY4FFT6hTnjyT/HJ46S7JAhoT2ZBox310udmrQUtn5+WnSipy0MM
9a94rCO+DkDD/YdEmt1zAhJogGkOf2PkCdMD8GS1BYahqCRGy04Tm29aK2rvusqV
h+JA9XZHi41qiucQ/MKxKNFd7IuVJv1l5p+xmiWRyW8D9sraOMBlXlr9v9Z+6BUz
KdpaJQ6MrCjp0DYkjV3MpN0x55H/709Q/fWCBY31gUvWjw2pwVY+NkPsMNtMy1TX
C5dmSJF7W/bszQJAszBlncvnYCQzDvsEixIt9d1OYKKPrLchFLvdNHNnJkWyiEeI
alE4rsu9Gj9JdqYm/p1/fgX7kv39Y0DjbWf8AEkFg+EYI0qRDzqgwT4S8kcT75Ns
mVXUzBeq9Gu+O3LpA3/jXM6kBzPnVBrut3xIfHj4vVH/E/ppqtvXYSKSOXmZc4VS
8qz2mvJh9k0F0BIO4KFT69zWbISHbOi09KIo+p8iSYkpU9tO/HVeTD4UvGb0qVis
KUU1JHdaZeKNKmXIR8y9GgPWeDwQPf7NbRhS2yuvJwSPUqz2yqEbaZ2VvJXc+03I
Jp5yltu3LT32gNlkjt2z0goS3IJ1M5pqORtkm1MjK52sX2/lvrnS/kgdKEvHdMks
iPdIRdFTAuJulyOp1aJXAlM0ODlOR4sVnxZn69y95qDm5cs20d8vo+VFbtdKgvLw
PkE2oyTb0uH2dt91c19oesBQwxwYhddswyQhhWGMX1mWn5B1YZP2ujoKFNM+i6vj
8vTsiiINw1etAY93d/nwYuR0guzQJn166ZfSmP1fuCdU9Z4yuPwxyHi0+OKtyJME
/ofYnH/bLb1/db6+IZta+eDZfqvdgYSNQ+B281VSllUIPR4lYQKfkyD61A2Wdbeh
yBSvXvt0miC6+rfIMrf2BesA1dLU3JN6sdOTavapgJY2+IHs04/nLWUC8p3xsGVd
KgNFdiFXYJNb33WAvGUDxCq6R848hiIRBMoxOit1lOxCUFVhfRG+eydiSnBAUbny
vpIsR1oZKXg/ygkox1KmaCxRr6h1QM06klIYH5vQHOVfzNAStFl6Bhqjz3r62Q10
BrF3nTDTcbvl3HfwYa0+FtzvxwTAkG0n/pL+eZP5G+An3EreKKJBgPKBPXSzvZCd
VNwEIT4CF6V40qowYWzw6tWTH+I8UBaiRDzXQrVzb5WEiudg3n+rz5HhEic3SLoI
Y6GWA7iD4cKYUT519T1FanltpqQc9v/5Y0Nn+zuUJL3Q9EfRMMSbzz2jM445Zy4g
k8yXf8IwZXCW1OQJV8fhAGNMFPp7D1s7cjAIyLe49PpudM0AjmUyK+cZ1+ANgyp7
9DpUd2zHWGHIprUcEJrMGZ3NaN4NZkQPC+F8sbQDC43rNEVvX748dYTLQyiTr85m
AFHKk/j+/gf8sD7/I3kWD5E4CwI58kMb0/XhOINibAbAr79XW5Uhs7vM9TYchYaO
duccgK1I2OkhwHjssKo9So3BaYLxyfWmugNBKIOabpgrvKzWlu+oyBeNSHDlwnwK
qsvoVbvpm/lEW2tOxh2te+PXGL8jSwhofwRYwpMu3B1mOpYRwtScdK4obK6ter+U
58ts+gNOriedrTVCoLHfGh0YRpByoq5t1vKpJaLzCYm98PEh5+xeqlf29FUbbnLC
S7U74IbEsTFlcDmaxWZ5B3ouClPKT2GRtv6WyHsDSQzOENCOz3omagH/hRdzvLBJ
x8bAvIVIAZkRp7bu9tv6vmDwS76dz9oC0oqYN5AA5YdBucXCOK9EdAjH7iIamFLf
wRkv+PpK6kpItYuGCpDOOzKVimUZnWOISR+73KXFBTllAC+Re7eLFRFM3NDm1cYL
gcld0XisWC0Y9cBt3sfoLx0yQJGcWGhq+qkmVpRMEBBHn0TIajw55glhfXVIFivC
1ivgLIVzTBem/CwIk8eS35Qtyt0vNeWl4MIt0feGUMg1jX7kxx+NwLBbXbnx9sY8
J/zDmdmipeg85OsqBpfrMicuI/6Ekqxg7mIKw7GxAMPyXNHaVbGsXItlgekMmyVL
GlJ3zAISfcJaqqJMHq4/fP72qJZ1LlhNTAtPLz8zVuPNcD9/rPysZxCEgjNFLQkL
fhEMhZi43AuIe+EpzJoNb+6gS+RTpo3/An4XTpNJeGCTprJF9vUqztsK9zG1g0Wn
FN4nbtnUgk1UH5x0tEWUckiUx20FsMLXsUsmaeNpWAj76IBPk0qpYh381l0l3T7W
3brnvJVa7DWpErVfYBeBa5ZksMqCo1CAk8hSsRFE/KutU587cunIUJERRqFDVx10
XoVA/AHNnomV9VUUid/duqjc+GDSKYpHgCDc4ThI2ou6ZrWto6f9ELjcB06ImtJ/
IeEybgJFIJc+9rfFQBpTpNNlrmijVkNq5sOC20YeWkboFL/V4wpHxkp//L+oHYls
lxULcAOhhMW8ofRJKvNUG1eDx1f3jk0ceaaJevr+TN/ubrBAcMMum9rD51RKXZxy
EZiCCulo6CgoSjVTnwucU/xh7B57cq50WUgPBCC+i/buIdB/PGQVYdXcJcVLJg32
gg7IvarskQVS0oFAqHSOxJdhyzkJ1Tw+nNI8diyOuXrJU2sHM1vzE9NdYoPNqrHJ
Z3XDvenB+I3L8eOvfBFWdrK4gxJ5Vm3nt755kjaIW2ENoFPbu2pAmBUmezUEAYFQ
5c9GzNT1DafdgSvf0LD5I6V0sMROtVUjRk9K/c0LH/42OdV8MEAb4zCZgLcyI7UB
Dt6RY2mBzD9ZC+uXV6IPzPRHdgP0sCN3MVonXTLmTkgKJh4S4bNWEz5dp52TEjNr
tTpH+87Y3IrfcM++FkNOrfbAB3HiguA0+Ypf9SURUZenqDZliCaaLMsrG8FmyvUN
9wbv2KK1d9V68OYxrlL0n144iyyeaD23XJYYIEEqTLeBkN4sGS7deTV6lJ1Vphwk
dFcM/Q4/DxKNb88Z1AGxNiKLqsZi0n5mDJMC8jmzvhRsJriX2n5/UGnChWF0kqS7
sGtcLvqAUAePruyJE1kQKW3l6fgjspHd/CTFsJgXUtnOVNFPGsbYlGokeAalv4Jg
VJsXy27CvnvUkq5apyCj5AxTDjjcBaDBxHzn5jeSGtHUFQuPFsM/Z2PFE3DByaHw
HXEYIJxBu9Sd2KhVGq+AV0hUWISmCpmXQQVSvm9qXBlJiL1RejRC+fhw3aOiAYjl
K8Z7tCo6yNk0yXhmU/e7aEo5nR2l8waqi8/sfUxBunCQ+mM+ShRiXwmNRGEJlZIb
VegWuzP/qHOCIM63HHCekOvZ0psgGnma+U51g5RDLnoC/6HVAo3AV+GfTMOsZkYA
qnRkR4uR7r6mj0TnQhTuyCdtbdbEtpNFxjoxYHFnr2Jkc+CnYhYSZrGvd2W9onL9
54kYF2P3oa9+YvbytKTqGcsdrFYyvPGppQ57ZuzbrGzTrLv+hgcGOO4dvjzuys97
EUPpr6NmVb8EeqIbE7UsGMdG5ZmVP8QmAyaCgXLRuc0Oy+6wn6wRJFLdkmgscj8a
cRQOGAzFeHRRaUwUHstNDPVkK5CZsYmK9NMiWQaInUTi5w06J/7Iqfshggq8jmgO
okItJCoqggpOtkrnD4SXmsUtFB6rwSMmY/W7A20h1OU79KpqEilHIkQyxELjCXwQ
QGhpVpvnJF6NT0NHtfauzzdwckkoVQwfc11PeneS9R7KVdR/c/EXSKxwqWa5cIMy
Cy8SNoDnAphGkPMPe6uAQ2+jCcvYngpWcT3EK0oTeljESEOoH3QWFDyvcyF7XSFp
ht+ayqJDHsd4TAQo597xgXULLeJHpFmyjDotak/3J2mWj/1hObApMAHWrTO0AQKZ
RIbFkIiFhHlYSrjNygafmq4Vjj4TTkKh1JzEcsam9npbenwdNceor2XMz7+6H4ka
foESU6FjWuKT+9gVreOL+L9Ie0IkW8tYSXSzFkC4clAs83dzb4pvAysS/yNwFL9n
biz+bF2LgJIpOgOh2vox8BnlFRTW+33tyanH3qUbrSUdN3gmkeFG4cRtDkNA3KD4
TZ3mDnJ1lOunLqUa5t0+/20Wk0Q4bOZJmGo6H0QG8d+w/+QgHRI9oiY4KGiER+X7
VROqplWjWfMYnXeGkk9tC6zKIkXrWy2DMVHrH3KLZKpN9jzXnLkpgxxaqr3SVQJM
hho/CRRUJee1dXThmkycatIM2ipaAVXjR05NGDTCO65b1/hc6t66JXzqZPQG+At+
DG5BHf6HJRIdu6PDzdtv/dvcKnRlr1fdI2xv2T3DqsxDaBGIw4rUAehYuiJhoBOn
Y/TV/Gt6PRnAu5TSjwmgayE0JdStd9S5BwvCqCfUFWWinAldPmUQ7uXkV8mfygYp
ieJP1iPNGehaIQrDVsnx435pH69SXTbr/f7SOFrDKWLkEhVaTynLIkh/zJBvy0np
BYRISUNk1Ep+2krO8590lpcOdV67GjDlTl+O7rM2cyd05DQAIJinsR7RwUQwX3Fa
KhOBRb4P1kDycNpwnLunyFfMEakiw59PhXdKFh753lEWc81RLPX/m9iMK8cSZEkp
e2ioFfhzzF299ZxQspXBLiQelGgXJZjJ+9BMjhJ3hvYXq9LFB+bD/57yX/qByrUL
EQk1jUNIAYZNQeVlWu2bEY7TUzYCuFJeE+3qKdNxb50il+ZssmVZr58LZ7ickNSp
A0xEzpfjNHwgPzI89/I/GtBVRaEtfffDwXcx1NxewG3PCfuIKYWufhBXZ3USmkHe
xlBW0+Yd82hTL7knS0NG3ls/4Wyy95quR/lE3XCH7yRa/hwBmWSpuvMW/xkscwCd
sC7wXAgIsVdyrFE6QbXeYh4wg56+otbAzMrMSItAOSaoKeInLxZu/BwVQnSyGgPZ
7qwrj4HcVpKbuRMBJO9qdNyQiTChCT4B4a2C6lH8VEml3yiTJDCJlgKm6D+5/BtG
ODVfSsnmlmdMShPVBMuNhH5rjQOhwfT+Cnil2vQg6pO3sv69rwm6ay8uNrRkewbw
vhxX7rG8NffZA5fAiSfC9PyYxTEw0zs4lp1M0yUCHU2vLwu0kxADO2OZdcGzTJln
w23UapUBqSEQ4U2JeUdGGlOutdHLTDh0lvhv495M5OrIBW8uCXNzNirjT2+XHBJ8
oB6BoZX2Y6+j708BOX3dSR5H0GGeQYnwsIB+sW0QfrdUEqobPQqNv9EkTZB7oB7a
eIKThf7QA20p/nl5gqKMV8UNJALpxYFJEq3la3VoQFgGI4V04lQ6YBIXVGawjKqV
tzJg9DvtPAOyLtBRpzw80O1MFrbrvkNs0ZNNt+dGrJeBPKiEq9Ab3Q0Sm8ZrYgqR
K8IvOG5X0drzr5qjqxZ7T2/PCFx1RUIONUiEqFy5370NvsBGIak6G8/AvAwnEyXl
Dr1nfbwJRfyxbSILWytwpuXgL1lzKAbXO4nnXKkzrzRSwA2IYosYnyb0QsNRUW6r
r84RFpiDxknvoCRyFOC65EN/d2S9iaMgyh8nsO5jNHsKTFs1WPLaW/MjCnFLt8AG
MnubUWiKqT9oPD9nxcNqTHF/ekHXI6wEfXQulZoFof+EkhKJVjZqy701ev6bxrbb
PjIjUgsgUS0smlLuejORLneLo7xInluanYcwMP+71onwDk5MSmfXHq5OozYGT181
QlhoVInnD1cdrCXyxUuuaeMcG1tYUr7dyY2MsYNGd9vt0IijGDAWAUAWd8VvASGS
WqLQTGRUjC998TrcTODwKlQGQVwAEwXYBZehbMabucfb/MOmcMBJFpKNBQYzPPdD
h2+me34/PN01K1gsXBvzQCN6uY1h1ShaB+TeOJ1gazJiQoaGZ2gpGFFdytHEiSj6
VQmhrWRc6wPZhLUiFukyxW9Nagtv2yqFCUourRoGdX3Lf1THraJnnAcKMArQOx6e
HTbOwEbrJmPxLu9EQpKjFKGh9fGfI/O27tvL9amP8108tZYJ7u7pSAo/jhUCNHUQ
4gh1/0pT2KtuekR1lGAdRum8tC3tOUYgM76RLY6J4h1hlBK2I2Gy172EWipTwMvC
d5GLLrfWTYCFDHkRp3t1/cMoILPM6QJi1PKYQVbNl6j9hlsaQs/SRRruBAhw/YHx
Dn1Pfe1ExopMddn7OzAR34VgD+ZI9ABaAYdsMS+7vLaqDsXS5Y2uhm94yzc9PU2Q
nPjvpKj/mPmoHAO/JBB43gjCYuwQ7D7qX7N2O1xtwT+TvfwS4KcqAEda4gDOQiAH
2KegkhdnGgkp3WETXIEMeMyGI/YqOaeely0+LFhGFEdQQs6uhlqJpmopIT5vUFOn
4H/k+U+lwvD18FV6ZajdE4oBcfhXe64i6rijWQJzMeac1rCR7MqHn9BNRw4IgSg0
nbhJl794R4BQwAPbPcLUWEMHP9sD8mF4tM1jVAg0dv1JwjEee9+f8QeGbY9+7Dqq
x+53laF56qDK88xIKguCBHsLk8sVTuhrOYR5p6HUdFIq6C32fjeAwjB8bwPQU0Pz
FVcXvZ0ascFkRsknzrIGl4nPYuJRV8fuk57G2NQaOEuXHq5TUkAS2LpwV81ENCmi
MGF6fQM3pTn+exrAFaNFQpq3hOPxwJ6qZnnIfA52TsCxLyKI7UDThADYQJft+sW9
rRqjFm5YV35IO/7N3equegeid2gF453/9lIwmz/G+4gd8XwNt3NO8SAXH3V8rLzM
hL0HuFWcyXo0UbwMGSDzr06BfdWxqLvqbq3eWctydnEUWmQ1U87qBDaelyTZe0HF
r0blCn/u9ELsZysk9cQ37HqgZUY8iuFv+RdRN8Zgn1RWBUR+ot+L9Lf+zyyK2wmY
oeVwlxFH5l4S+XpgAMC+rh8Vn/L+m7mVtXkzGpOUF5X/UjWkjQzbgjBqTTKjMEqE
hnO+moBF8J2oYrkgOaEsCyLjVeQDdB1BVua2o0kBCKrH9AZTwk4OtBs1Hbta5F9B
ITjRDdDVxi1IUBLYsutg+QbqWHqn3U/hizuFPR2UuFUz9lAasn08Mj3goyRkF/S1
X6oOkDNiAGWJ27QoVBQFNUJm23EHJ83peUU/94d8IfpK/pxmfWJzVdRWujGDYj+e
ZEs41u9WWy1xdAA/4Q1eKO27Z4mni+M5NW5di1t77I5qfrncnT6emTdurJOmyWhl
0Sc/TUUXm9OaZP4WaiJ8xjumc1g5UMcnN8mrnDQcnpr9smW6hCXbWAN4+9KjTLPq
ivcL3YiEN9je+TrmwaFXlRbAYvq58Lz5Z/2jT+pERXf9myIPnaLNP5gp0/bYLYXj
nqxxK10lw+nAkYcAa1TPLqdHCt+MbDrvQAYGD5nZMttMsdZP2q58Nd/hNS9vm3AU
C0c4KPSibVkBYkSB2o0wm64Pt3YGf2kmU2X4p7uELSX4JDVFHdWdeXJXZYfuzlmF
y5TRsSxz1bAg+HdOVqkeLHPM0gQ2jZTPt0XzXvUUquc8Qo26TsO40ybfgRF9+7m6
3gwkpYucCtUn8U61RQVyYZzmhFtah2+5d5/G4JGpiWRJNdRg67DSF9pBhPPCALds
y91QExV3zZzNKjcNL31ht//hAHkeF+x3Oi3jtlqQdhJN9DF2FHiIXIPxfX43scLE
uuoO9JC9ENtXLSAHu6uSI/OYZiKFuOpTH0r8LRufzYj82i9vD0VhekiKW9npvHFM
lIXt12QpKCAfYr7eAl4XugOz4StiIHsYIEzpoXjvMarUTbgScmHm/IJwWc36MOYN
yx1rpqWqZxSZutwsT9TEs3tjUaA34STVQ/fXZZTzFLL6EKQy/9BX2tbvuhjJdvX5
48x8Bs80VpY7WYBeVPEoEKvKt/cWV/ncT+xLZdW5wYzzQGfPWpukkfVnCuHJdaVQ
a3CZ0WJ3YlJCZCbQJ/QGsrxB+j9TPqOMbQpKYx2d9bl6rYMFMYh7CmVVgaToahCB
KuQJ9DL3ES2ZjgoGsOfmvcqT2YhyVZ7xpAWvvfKKPST50btev+Gnak8SeVTe2+zj
TtqROufRw0zHLXMD5BH+F320d/uxrcXv+2E9nVSnYkEQv1Uxwh5Bx0e2PP4nkxF0
QkkCHjnPhI5eN9Twki/p3fEk+1rXvemuzS/ysdh/kZKX3gwJvu6CYU5MdEXEONv7
yGsB8B7lKYajk1TAWXMPTaDoCYjBJXFjSWCS4UMTXv+WqFRykLmpTCLKHJX+Ly4/
LQsog14uzSxnhWaOoa5d0cH63vQ7bjMXk4YQm+S3I9tpvOQrmAUM/zLCBMfkUm2D
ZRwps5SyXMNHqLzWnJVtZrr7VCLN89/CMccoAb8xnWZm+u08iL5yaHppZPSNtWi/
U9rDTcAkIbgJZPowlCRuLO4M7Ag5eV3nl7pxoJEqeZsqg5SAr1Ug1M9yZr+0I0wF
0KJHgHFVz/Q1BwDhBDawQkWK0f1OyeG6Th3uFlQyH9xSciTGgDwGDgKPJdPdfSXW
hT4NDe7w50IVHG87vFTjUsch5w73//oLfLMPd6+Lx7np0lmdVJTo/sOt6Y/0hVmE
HamiBfY/S7JPiaPeMZvUwYwlE26xaUYS5Cj8PG9kZT2pEWJBaClsuhEIZeB6VJWn
PYBIEPe3eCTNQR6xs3ASNselxPakafLpzJQDw5R5zmZz/v31oI7DP2W5MH3GYoeb
yfmXDccT5TamXq/6Gy5j2Z0nUFOdlWKMdH4Guhfyb1PEizu9BnXMkod5WACWeIHZ
10SImWqguXFtNpgTqPE7TwqrQx3SUesfFUHuGzOPfWQuHTdWlGaWLETCOrg94kbq
S2aZMlaF+c56M1e4qRetLYsthstRRL1iXzRpY9aiT2jzGFl6ORWfDnXdoOYPWXIM
WBVGQR/YvGKXLdsAIY6Y9fAKxT32vxVNtrpCdwZZmOoyEVzgzHtQRbPAO1HfSkR+
BA6BgInz4Msm6OiEaeO0ztcJHnD3xYZzmeXIFIjd0yGt5ioHonmJFlotT86JjoLt
hzPdvAVj5ql2pPKZ/enirdPJ4FMakkHbz02S49Fc2tfkPkUF0+lHWRTHQww1YD1w
yH9TI8YDMMS6RJUzx+RrM4pPlrGaDrLeYxPVR357/Vt4VcTuLt3lRms5kOh3WcvG
ThVf/dqENod1iUOXWMTSLfL6PkkR5sllukvr456NkA/BU91y2y4f7t5WADRVPuGj
cwRpS5gjp7cfmchteG5JNXqKFdCAmg6OsHJ0W3Rojlq/vfInDCFHSZ1kjHqAc18S
TcIv2RKkbjlmxqdsbx80zuvBgW9OUEuhCXEIg+vZOPlMcnZBn+oiFZzagtWTfPbg
bJCMe9E5qXT1h+IER/7DO6O9cvqAJ4GrN7o4QguGKQncqGVSzVY0oUEpp+6P7447
7qxD43Km8U+Ho5qllByS52E0uHJIj14XKTykZUGfTvOmTiLzuZOiHB7oHh7vceuW
5FK4m9mHM1dYSy4d7PcrzjfP5SMj5iSyEffDXTKfLaBXORGfShB9JsbIoVdAGRXc
Ry4OpgLsBnIPMaJqZFLkXdCMfuao/W4U6aztG5TstY1GXxDYnjRMG6CYgnS72bY1
XHuzhIdsD8pPT0xqcM14hP+Wy4KIv9ZSVTnU/xkkesSTYsLlznuEcVMYprsn47bw
r/vahI9BPeCZvt8h8sqacT0BvH26dAkaL6UOhHB7Kzr2PmZbGOQsY1wXNDmTAw1n
6/JJunohb4WmXYkR0+DAFhTZlVLmXzYjtp/aZphA5djhQC94iIlaF3M2S7Mkmi2r
x1viwpuAOinJqXDddJGB0r2162XtnGu6c4oZluI5cHGJvcWtawbb6Lxvu0uWHINu
rejAa7CHQcTe6xFAp9z1Zqw8xPeNXmy9ukzbbWnEFwAcO/R61zWjDnVNuxUTI25j
v2QwfdrGXcLv8TxS07y82Z3w3LwvdgnZtnRCQOHVUz9rw+jTepdpVu6fBnUs8QD+
YglVuj+CD8CXe+mA8FKyGqSGxD8sjhBmAvWjWbsAIOJmZ5f1bKGxidg8fHSoe0zH
XKPxZCJmm8BuxBlxF+NBBdv1mc0DTk4TZsGyvO3v8w34GhS7rqJrN/f4GGtVDyhz
6zR3uNX/2spRqTOIoOZOB2WFDqQjIX6ZFiTX9VUCmYgePPiO0HV07pBIVUAPA/YO
q8xFz6vIjSolC6rq/AW6UejCJ1FyozP0U4dMTlZIech97KfMLNx5GBnMi/RduL2J
cU5NWyysDnVzH3nQRRa0kW3OX9Maclh48rFl9pRYdYB4vEShqdqdi6FAR1/XBngA
4ngQ6Kgv/27AE6F/pCMUSLxwwTl4QuiFWRAWns47qRYlL82aLsKL2JLKRyNBV15L
RHAcxJxVRGboUHoipuRggbtqIHJlVPSAaovYwKoYt7WHYtPB7Xug9WXbDRPoLevp
nhMPdRy+JwSy3OYFnIO07AV6+EpX+Vlx6psS6rgLHme+X+lWYr7P1GFHmPn8gM1b
Bj3JatYx2xtGADyhF3HaWsyDBVdYbg7Mi5O24t2ZW3nsm0mAvpO0OgnGSjC2Zunk
SVvT/uWmcyh/QHWDjhnsWkGTwYU/wbiAK/g5tGn34Si9Fw4o2lcQEiQmt/Q0pYsh
haiumvVWPQ+tEeoBbqUv5AOJPJ/Ho+rmBzOjoSxoxNnoNkepcSbJyXQdBBGLKrCC
e24ngEtQRMPemKFkZCOhaMP0+GJMScGjzYJPwEELx7KhvO8Oa7aEf04YqaEbrpxJ
1JHTMCHtTI3SDczwZGFM77JVgnbSMQjSpomfq97/8e+jeEZ17uK9RpFv0pZQRxyt
Vunna5TAOKwdVikLl4216zUistCCIk1qBHzFBhwz17iI27mShRgzN6vQoFhnmDVH
ku7gexn5pHuLOFMLglmrGH2kWxny4zoEypmJxDaxwwpm1Vyw11ktdlff02KFE4sE
2zh4H6TNx5wSRfr0TvFyuNtFfKSjv7UTzylhLN9KtwD8v3SMfK1/MuvAy5/hSNxn
hczuYCEvCuKkuZu3SwtOaknPtG5wjwNUew9sjkFWTAhv8LYzNX3G6Ti3Aie3ddqH
eNqA+IqDDVtQeo6dirQQy0xZE6hQtWviwoubXsZ/2EE8yoku6xWe/j/b8pjldbsE
jCUXzzstulWTCa7kWmXH9SfsuazZOozSacaVw3TI52P5y6TGI8vfkRTIErYxUPAj
GUoZ+NTTvJWpa8u1xCYs9KryCtczX216cLJK0gM6CKmRZZt9uYfp/XgPr5Lkggqd
Oew8IUs9EaZPo7+XjJysE/Fqp2mqoqFRrp+wKdAZ7vpgFUzBDvsyzlH1VVojmfJC
GA+CujZQBV0Gh1Io4Ez3ZB4GQ3g4WROQIDDfUKbue5+G0e4boMeAm1c3p+9sYwLO
eD4ICup/jfC4MLijO7hzanqJRvH0zPgMW1UtchpkQBFh8xvl5KoXFqiMDLcCfw1r
JHsj9Bg64UyLiInbj3UoP4oJfEyqpD23e5cJY/mGM3XQ+pcUAXOTRIC6IDec57jh
lxn/e8aBtPmAf8rtF8jWGKr0Dxoj22pJ43v34xjFnmNYsvY6ICFUPX6vzwFazbtT
epatGRyhokr2u1AFpsuKKIEFRTnhcvcZy4a9GSWMXpcmjeU1rPMse9kLlxKweEm8
pN5mnyG2xwqg0R9BXlLz+yfyFICBeTkr9ewB8af1euO9qhDzphe9xX44NrgFUv5q
uuETwOoVdelYMV2dn0uNzzfTqLslz7Qs5vei0am0QEr8pHgHXqTkarvY3yAnAf+y
FxZ2TSGGtjLVuJAjHcdCv/4GR6Zem5tQeP+tViizYg4hZtfqMgayLb+wz0r8YWoY
5rj5WGB/86ZzRf4RtpzP/e3wevtB3o1eEHxLUZwMbxcElz71uCkHhs2ccd5udmKD
oz584VTrg7lbHpUCfYDCqMPlvZXrU7qxVJ0CWz1Coh1xGg+iBzwNBPGwD+Zni6Rk
fjijh6PH53ABCQPxB4dxQhCS905mpmpTnooqzc7nD6oYvCc0OQmdX3tje4Sk0tLW
jzbYPqyJw+6vCIo7nyG2+HrZW9Zmax4P2bCIeJSiXsdxYYpuFBjeftuEBtCoJ7MO
sx1OxfFjuiKLjL/rlzfHwcQYQ+4BYN6H6Yj5C3OJXWBPmIXOjKacfnE+rENAIfz5
6f4v8jdvBKtLa7XcH7R3OPxzKupYvvc/4TLwvVwKX159m4ealxbrmKad2/x0RwrX
3rTXtEcCjE+OdmEw+JPiMStFsWG7OCl2LWzYRWbOh8fki+9CUIKFL1SK5ai0K+pR
NmfnpkZvR97pJvNizNUc7SYc2Dmuvaea716yCTEcOyVKix2tATCVsxJOIXwv6l1Y
dB+ARt7dB2Q9HOsO2MB0ScTvwB+2bwlgPQIdpgRfdkwfcDWshZ3NoTW7aud9TB5m
tgbaK57XVHGKq21V/L4jRuwkNYXoZ/SGRgawWamZupS4Q5J9VrYaOA8Q+IEVLZPw
xuJ+EsaqYkcEpGn+ACn6qkLg32W/FlvF+FlyOx3gUM5R6OlBkzRnRTRl1DMJEjN7
FJPE+1QdlSqJnYvzZwYH1Nd6JIFNfrZXe3z2dT0OCJKtBYWSjqoGWDtSN5V1I6aa
HF7lawHw8wXPtLqLYIid2Wx93Hvvo9HmDr+4H/nLutqKy0IRZRkVX4qW4BM4jvwM
Ws1xu4PMwrp5iE8UpfwhsliOcUGd/DyGu5W6RvYshm64OPm6KYtmYcKdf9pB9daD
3WpdiBfdrhMuCmQvTUBh6Rukh0gfrLTZfuB8KpRmPuCbHZ2VKlikpqktuz/rvcTc
LEVH5CunsiZh5UbIgJCOUzJcqZ9Y53d8kWzMMsc/YQXJc6G/uI5urlzAyd1tZ37w
m0v+WI2CFRClqkkViQ6N/KiSIwfYr2QHpw9B8hnWWjBsUJ6uHZB3SflKy2Plu3Oc
I6Rd3GuPM58Rqiul/iSuR5GXoPejCdesf3S79b9rMwcqN+KgxjtMFhpACPEpNxCT
fVwAkP5UJ9WKPKtF0qItp4NZIL+Ha3kwsc/BvKI540MwOFw3+ejdxWWrFJx0Uxhc
//w5mL1zhvPoLLbIDu4RpC3DsVheDugPrUnN4A6btKMqXYSHZ9ZOGRrWB/8JUU/b
Jze7MKv5C0gY8/87Oq3AMcYvvNNV3pBuMD38LMprPPppBljdp5fg87esm743EltD
dNsKNl1Y/LMYb8m15tNOWdomaVoPW2fSQGFd8T/Lc2RcK8KUHNB0XWNl42mmdDjm
Pl93nvUdOKje9dMWY5aiTF6s7AM/76520IusQqwXO1GFYU8kAqUC1NN6Gd0VqLHT
Q9oG34yZSV3MFKLoUG9FuPXsE6nBCYewQSP3GQZJDzjOIOjLO+s3hyfkvvbFs3/F
z4Jaju6jXPHfZat0R7xI7X0hrxbS0O3bFrIX4tiIXAPdbTt12wT1wXRr5F2/MJki
QvQ8uIKQhVseSsbiUHXfkrme9G9zdyjA6t0Y0O8WCMcvNTqQ5VuX4U4PsOfGNr8d
ogZMwI8vcL9N0t6huVYJ7sCTgsgy4qIM995Ve9Mo7Mtj07v74TTRihfJyn1Av1QX
S8Q/5NZIxTw0YoqXCuwoYOYUJVY7otdsgxtWmSGATI2mnOYzwV7oxOURbJYs9yN+
gq1QJeza6G5Zm2ZkWqAfTNmTzmYtRsZIi5J9UDCwj0W3yuDwV1wH1RSaATo4xcxO
UwTusu5q41RWzFAZOefw62egTJv6kj8cpewWi+5CMP71K3psOHVn8EepaooP1S/Z
ke3A1G5MLSQzy8w/r5udyUNU7cLvD74REVEIssE+iWxUTqWAbxbcg4DDfG2ItB3h
oeN8lkh5WH7oB7ysUBT646tmZa4hZOqmOKEIPwmeyYUdg9pU4574f2xEmPyouIoJ
00/OvK/PAsPfyLKtohifEsIqlLwrMRZvsc44Ijy1IZJPtWTCpd+JCDf5MZfnBUGl
MQt7N8FKuDK5V13qtFKb0NaVzYkC2kV38wn90TtqSWa5lqB80m4psveOlmnThgJ6
yx43jF4rgCTEePmjibLKbf0vujtIPGEd66Epr9neqNRqiJumUfHXxyGcRQxQzfhz
y5q3FswJvYx/a7snaqJa0jSjswCr7knURbS2DH2D6oa0uXXbmIyRifINDMka0CD8
EefF9CanoHmAwSvAANBA5mp5PuUiG6f0gf0VTkbxHv6p9cKWQtskrjStNt/amhs9
5exmS4pVpdkN+dVrlHxSovo4RI8HNtcnPMIewEhcXFjeEZYx73SqzBESFALbpg0Y
xR9yenJ5YWsU634Lx9gVeGuBVlymfoad10/nBgRmV9AMZ/YcKefWWUli+ixWy22A
LsLpKV2GE5BlHNX6qO0E973rT3JGNk5sAc60gojelFsyRLXqiL4jBH8Cd7yTHP4o
er1FXnRM0McmMTBNbwTe8xfyuz936hMW2Ko7jsSh7izFyn9KPBzXTWHkH8PSQlUA
7CVaZ+wimsmAbv6IeNMJebpGbVMSscyGlB/9qoWugYbc8w5Z7ezgs93VXdz2/o/z
vUB0wrC/Eh6rr0Amhg5pqqElTGjjrpdaH1Ire5JqR2RvVwoXrOYLbjhaJgJY6DzQ
uJrOmyMS+ZQWRnaWAWtsi75wWiq11P460x9y9E36cFrkahai8BdwCjdnr5maJcFJ
6HI3je06JSgjWx8udPhtgPNwAAURgXAvCqIWdkb+TNxaf/cpewBBhDOTVnXRTaqp
EWqS2KQMTJmvN7ijVQsv8UXBZFZsz2laIgxQeB7dx1VtUxDoozBou/WvXeApFmGb
/C84jwNVC8N0hw0Z7CBlVdaX+TYSFnQJJZh/a+I71nHbq+oq3JgXs6WmLtbAfDSo
7+nbigg8zLu3IIFUe7KxXJZsRAkQzcGWSTkJYexuP0FiOFUF3jBH4XgyG2UY9FFN
Ij3729gofyEjjXrkjdY890vC2iWBPV0Y+5RWjJ12BuaFNaHc5KpXNwv8fItI4IrP
yA3xeTLCvYDNabxSqOkle/IyK4QqQgRpBfSCcQD+v1QeupjGL09F1czv+PqNzCdx
bRL/eCyXFl+KZXp9Nj9bXyVcvUn6Dus+BwZk43t3AGQd5E139PNbH8oYPqwMqChL
J5xH9JOBtJRrFQeEYrE3lESrljzec55i4Z7TWO8Ts6YygxDp7xCbCsvVV/y15Bi8
toB3ZNxjXdXQwZTm7Qz4Czp7HoTxl/1P2eovKk6RjiXGbc/W85n5sL8ZdIUtlIZi
A+rDDPio//YYpMhkA6fT7xxhHTzgVhusOQVmVz6MAgqFWHPiTLXl+EiHATE3wnJK
gQayFqSjffu9sir0+hTjljEI542ImtwjSzUE9cJPuF/37Y4FzctsJQ4gVKRXJHvU
9SNeMKyVtAo62ar3VcxYK1zNalNV8GGmSG/M0FRWdeLiNhkkHCRY+tHagiK/om99
yw3QG9QpmrOufDMD3eS2ylSPpiJUIrP3j8e6RQv7gxwJCkHPS68rANWt4L/lHc5b
TOZ983VXtqS4ch28OZ+DVgNhJPXVRvxOH18tXY6i1OTKT+N8FmTqXWu70ipttj7H
9Y77ZED9utmoSAH6LOCqdh85G/pzWV4sAmmsj/WMnPMFhgooOGjNDss5fXKbgs74
EiPSVKmRgTmgci+DV/1h8PUVnFddnJc4ZVkteexw7nSj7tereJHUDM2lVxMJ3Szg
4FsaAYvD7j9fBmtrzV18/nqAy+ymVSC416fmgK+tra/wJKjCYaIGPylM7VEjBJ2j
UvoLQyoqjb/Q+6Z5YBhK7EqnOLMGg6MvZFhw6FcMEioccdvld7CN90xByTWlt6oB
kp21RjVjGZMsuommnZeJM0GkgydE3aShUxzP/S73WDmLZE1D83JFJbLtsp+8npF4
cQUJOV2JV0ZrsXI4MHIlUovp41CJkmcuWgU2XVlABXd0qHxgSOlUmzBPTDEM1Uuo
V/ozypDbw/kwAEfSEw68W6UaGrCOrcuhHPZKr6YQ6i4PQ3PgonC6szz3KigaIPGY
WuCZU4/5gMkJHaMQO1s0JybBUnpPD0eAczTz+j8BbKzP+nxu6PEPIBO9cGLuqH6W
GGSmtKXOT18AUnNyhIam7I1pn2X5ilN25l5tE7jTjbJE0DTcKXomz8jI1b7yKM6E
x2N/zSLNd1SKoTCsCsETnJQ3TWwiS8wUWN8Gjr7YWCPcDho7kd4FW+IV7DrvgRqn
9BtFvLn4FX6FdMvgmtsWvSVYalZrwnwX8wEmQUrjIbMyrfewl0nZBJcLtBWlTyKa
nn/TMC+6MzqsSH/3vmNXbXUgdWbFzlnAEnfVhWaXRF7aYH3BiiIv3zm0rVGmwjW/
M8U8679KhWUuUS0BO5GB5dF/yl66etR1FVFoc1WchfV+YcuOoiFwtlNKh6fjbEVD
IE5IIQq3l4qBCso+4UR5OIpxdXLrN3RRh1ecETz4tmn7NBl/P4IkZi2W22bNUj7t
aauVhvxiqflavEGPRmUCwWJxaPOvk45Bu7EKGR05Pek8C/vEApuwJh6dFYbSqzxU
gfMtFVIPBZRZ3FhRENPXadL7P5Xr5IQ/5kfqH8rGeuZncpynPfFKCcC5O0RigejZ
FhjoeZhEvPJfPhGB/ffvwNYTzhc2gF+yNh26dfkOslFvK1HzqVRuDGjdf01oU/CV
ojc9Nuss+u3L1YjTdYin0jnYpN4jYYdu5DNYkZno1odg6pO9dWHiBVdTaMWhv2q0
Y1gm1W+lhhkW4uTtUP37qhSRyl4IbD6ibY6L0qXnexzKDjX8+r6qwL09CvHZTDEZ
ZhlZWt+pfK/djFyp/XA9AwTQnjpAgwWulLBAYaK5hQkAIGliOGm2IRoqXVyfvQIM
8J1vY1KfWM2ig7jIcg6mBXt28b/BDNcPd10KMxQteqmOCplKE6ImyF30LBchWtd8
sZbRPyT5YV3aTkY9JBA8nysmFEhES0FwXx5KhX6Mq9k9oghdszoCHaHKZBNPcq8v
yZfoNNdlNIqysiULmReZOD8+0fVVshbsKF4SqSdJvxpCuDnOMGETRseixqua9NUG
x+5ao43kKA8uQMfokvtsTIVeES4oz8se0b2nCQsdViRhl3iCHbHVBFkfh+X0Fxl7
BGrJRXvPZEIQmnGsmcfVcKpZqmYZs9Cz1NecRkUE6+3oGx3d8+h+sghNbsMkN8CF
2e/CdsHxzSU9ofPh94sUtUNEbBeQ8pwsz29xuOMEZdfXFh5sBKU9hTG4gPOvaQnV
/UmNgIYP+xXrMa1rp+a2vw8/sb8QSDLfQFFv8PavJvEDDfCic9sdfxbVHvgl8I4N
gkBIou1QdIGu72e3X8iSIczEFe6mfQ9ECjspWfJu4GmHwGDATgNmHZXLLOWPjj3u
z6Gz+LlhAxIKmUnx8qcBoy7fW2xCJ/POHSRrU1cvTjCTsY9I4TqT/m/Rd11ajdMA
W4foevUh1k9idkmuFhVKbyKvyhJFtu5sPpKtZjXcz10jFM8xv1+DQEJ4OZKuYTlm
8nYY3Mrt4u2ujIgx6ShHaq10Rmn1jGlsZHieY9595jEGUVNXF4Chxs4PUW6gu8qm
Sw/IlL8tufnwKLgBuFnY5T5cT+jLVXlUFnJt79EmRoYGK2ccuiQYsSLgaVVy+ki2
f7eQ9j9k7zt4ReMAVeb3Mo7tV6PHsPjqypyATPI4/r/TvDSvwJsqwFC0qcsHjPU3
Jwgs3JgowpdtqIEjvmaPhyFu3MhgKS1keO+XttJ/Z5FJUVED4O/h43O7YjFXvDLT
PSMFE+iCGdySRlgWi8pXnTZv83EwH9NGuTibQ8WkXWAthcscW8YYQSSKt1GsSQBz
R31gCDuTrFV3LnpJgxBFD6Lj44KuKY5J1gUyKP+mKBICk0hDKkeMAP5PW+gf0owB
Kv8E8DxfJQbRw50tb4PLBh7XQiQGbidZmS+mSV0uT2yIflDcIK5GLMChmhe3sjTF
cxI486AKhOfaYv6aVRlffWdo+Fuk84CSBbng9svT28C3sLtUmZk2yJhTUkTrbrCK
r39OOYMaes63wDIeBTEpbmbXClLmq+98DnZw7lWdx0L48Ea3oxzLfZmyQXs8f5rT
gsqv5BH9a4Gl9UtvkBrqmhZX0RCCSycs1iBOmdM05owMH23dBkUlCC+doaxNlSQr
B9o6a+Q0Jgoe9YsPnWQHIIM8HzbeQ0h59wVOBAkPR/oQZVI/fyOhWPLHy1FVoYQN
9dBgZ+q3GP+94yWoXNLR+mfy4TD2NCA1eV2HdGdv7IznCs1d6bp6miuaFN11OtgL
82HlSOVJHut5LIXHty5MzcDxCExwCq9BouFUzeSXck8RR/MoiNWtdRybR1Ui8dDE
EKkTK8zW7GFeqAiMutBcm2ZurKM4vW9pVXDvDRMovPpPy1SxQRcNfPuWjbyZsnAf
ZpFWM0umRJQk9sOXyCBvQCWdM5EB7aZo7AQ4pJPC7RxR99jKQAvq3M7P9UpTRoDd
k8PTZjvWHOvohhlyVjMGjazRN/XjbxfqWnhNYTVecjh16twagh7+BEE/OdgQ+KZf
h6d5F0RpaC0C9HW2225PJENqHcAGtKu6Gpu7525h//0FXDiAQhX8eK9iohGNCcj7
WKxgdezVAugxOSkXRls5VY14EWy8gz1/OTinpH4AILks5xj2G2Q0tK2FzGw8BhLl
davPHsEG81+AwrU818SB1nowa4vBlDusYMFq1E6ULpBSHwmahT+bf/ad2M1ZDcnI
M+VgyUDpJ84e3a+LM8GhUip3Wr6/ys8Msx5xS+cVwWIWkt/W6kzrVrxQW1u+ttzT
JVzHSIhjBjFcypfnIHe/gVjzvXlKwm2G5fFsNVpiaTKSuvhTdSAEg1ikrQpj9kJx
HdibIpR7RrNz5Y9bjY6s+ZJjDABq0sZttXhOyYn5Ntky6y/zFN09PcT+0/K8gxUe
2ry9Vf4zSEd1s8FND75kMaB2M+IBWk2UNPIEmXzAqRML3r2tOc0ZtegbPuBCw0dp
nM48F0Z9eKw1YKxWM5JhdZREA07K712k8k5Ptlj0Tkow0QLJn24yWCEJbxwhBL4R
xxs7JGM2o5aaEm7sa2aKHZuXe+5L0PKlnYag1gTDDjIfrTXj4nk6jzGWO8HTr8ND
+jg6SLVV4Gy2K5Agt2sByrDXOt/q4jk1cPtijMXoRDoBNGauKJQBYRhz+cOgE0ND
+hzMTjeUSpIz5kbU9dyRJQ8VFV8vO8NvaegrPvk4B19nl4q9klveahNzSImWq2mx
Kw2BSQzRq0NBoXmY/88U/FjXrOwByyyfqz/81kXrLfqjT3ht0QcAZil2RlRrzbtd
gp1/cei+TtmLkwXBpA8Zsp3ixCo+FhE0CdTlL6p3vh28d3dxIkQPfm5LoSXGJ8Yj
+0zjfWH1RM31pI7jIEcZFJNYiLguC4bx+eMLyE05MNuyThAuR21nmk/la3RvN0aE
EHR6DIPKenKoacIUZFy965bcZTq08nq67iI6uAUZxRMnitL57dB1CVEUZ554WQ2B
4St+evtKb8+CNF5nw9VNZQUrnMhPjcpW9jK9IVXrGOg/ylSBM5z9bTHTFMzXJgZG
GKReEkw9Pe/zNLJG35vTv7I4FW21t7BCVMmVlDOCHE/yeai/lsDmWR8Umd7TffPp
q/lyrNDMXEgvihekK20Aq6QxFM8+32elaR8P8wNlAYFf/05i8rdeDmmx5GhQvTml
xf0UXp6ynrpjir2XyIKIJMhsb/iXH4c3G9/dsPcUHdfVN6lr0PuVwxIfXd+TpyTI
9+f496tN5X8DprqhsPNT3YhCKQSg2gZSE4L6P3Nw6Msh0aCFI7PI1h5Ybl5qm1hf
+4kq5x360bBYm+j/yky4L/x8MKw7acpOCNILMzuGEUWpcEtpp+wfJbmE/EmKMVxw
zagc1jNUBpOWDdBNbin/Ky1Xc1w5asAXHSiIvozupwX4FptyR20QzNkCRW+0WonM
V9ji0xd5BeZRwYGAJlsqBR06fKWogwvGAjNxK0sBA8+Zote8D88BhEndG1DfpAti
DwdEZG5B+yGbiwX+224reVITmkC7EK5TMkVUTAlGPpeEiSJv6KNaIqadylNpgraF
5YsGmF32sh8VtpKxjDoUSrEx2FgZDVcyB8OfsmPfLhqpv7Cwqw70wqTVH/ROtpNy
wkcVoE3HBJoZHbyWJGKF4yYM0SZtdQ/IKLosA50a8RJbEJUwZ1FXhd4p3wCmU/v9
Argi9UPtq7g89pSdysouq01Hwhe1NICkEPJ9yeV7rrfC22chYw5q3colozfmoxm7
l6CR6W6b4ki2OJcXWQLM7hLeWoS7J3rm9zJHYoWjb/mQLQ0fksXa8MYywB8TBLhk
Dn+kx0MqpB8sQzMgl/pabTGB8SQDx02TC5D/76yVqwuBSJPlxy9cI/U2BQscqkg2
1x/IEQJRKn52kGOuXCTo8mDbUm5UE9v49g6I9ZEWoDb4fBIvC9gPt06fGcUpXUY3
KUtSof4N0dWD76nGyEFw9MVGOMb50X74UcxpwKIdLlNJFDGx58WDpNZLRMOBTBc5
uqnu8Vfoc1besmmxlk0tIAUggD1IFX4hMzf7JK4U+MC1dXJ64hNN2/1DWjM4EvQw
BnnC7oZXbJ3MQFAKYnx5lso2fx1ccvv4wXIGBu4yPQ+FGcEbnmg55nFr1JDrQPJ2
7qqPaK835fgq109gVVUFtx4cK+HbFeK2pk3hpbil16COBsXfzXBFuKUkkAet4mFD
Hi/PWRMFaLTU/FpRUq/6IvQueTLoaJQ91k7eDLS5dFRaq1LvnbvYvmDh8h7W1r2K
uM8OJ7/WbPK2Q5migSz+7aUNWiBbF3Pqi7V2eSn0gTAQYiN3B07zVdge3TPmzmr8
im1KDCJra1mcfBisf2Q+cLnEz+Pv5pjQ4LHZHEVyCEOlzRDLmP/Riu2Qs5Odeh9L
awFDheje95lQhHQbg8RO/4IQyIHoKuNNR/7j5R5Sdc40K8vcPioYEXaL18l+1wPT
NJwL5dIIhszz6moU2lK7pP2z/In+ZxYoZRDlf1P0ATQSrNG1e1M1+/PAnQrmM1+w
tDZkMgfIHUIZjBRP0ptRxfx3/KH4L7NT6AgQWzunXuSMEqhDfzTiAOMJM/NxQrDG
gIwGjiWgiTmDPFa689e1C4HO91HcVhlg+PhYNjbdFpm4kCmneKyIoSEXkuDEPYEb
KYKtuF6y4dbyZs1lwzAPy3C1jnHjn3h+lHpTX0re4+w5pRDGJG5fwyCEFV30FUug
2p/L54nCGbvNSHBCvGiKxfBcxDfFIOTwUMcqBbdiY7Olb8odcCP77p03HzF8BtvU
psObkT54N+dW48HRaBgEb/ZHc5gh3ayFO8/A6ho4E5eFTDmtAFYgGbHxbv04fB12
Z1AbKdXhsXBZaat/1NP/TTSMMknljJXGq/zR3+lGmi1pzBKK7wjlosOk64rZA8jc
PFl1odNLO25YUZGqKQS3eE5zfd8AGOuGSa3tfCpdtm4BsoqeIAoMOvm8EyssPxXA
FCyhH3jwvkABzeztp1eoZe+pENWv/6sMB4tQMz2/zqNOHeuMZcaeVTqYCpmCMAs9
pzhUlxPoubw+pqB2XqDieW/j+HB2Bo5zmt4sXAwV7x99HS8aM8KM2/MO775vJckB
CN2dLDEepXPAk5kJArGUrQLiyfqrf9FHTK0qSOBw9kYTgavYCCaNMobO2s2Yg0km
m5ToX4dGWX5tdKfmJbE0S9dz1X6tbflKPSaTecQ0BXuRzN1rWy9E+WykWLDlF1dw
dDCW8Mig2eHmb7rZL5sQqGTH1+M4nIZzVe1JJAwNvG3Qyoc3zdWOrKIdlV0xYmeh
UXrH4qG1xvjG6xHpmtvM1QQkkhOn5iHENSpYnJ6xjQogdiIXZYWuxZtUbNm2KMmB
luonk234js2QnK5kNOroNXpqJzarjYPcesTinYPPcCOwH/pcf6FnzWwvEyk7uoIL
gcwtzpJ/gwKiPg1+mfo07hd0berN23U1hMmR7W0UlkwXPrFuL2M8b7HQ0DXdhrU5
zT/DwrtFJQq27ah47rckOMNyT7oV/Z7VMEA6syvP54+8reWge/Z3jeNbXVFjQ7E4
n65bytoD/9Ry2IijMVLZU5NJ41oUyDMP2cNggReFYwDh3p/o4iTbA9ZltCpTYhGo
vAgqz772hvSKX+Xr/shVrIJpJM0sjRbCMWhiPZx01TUzCupaSJmpmAVAGgeAoQuI
/y8udwXLh4kLcAYSPP9xwSs/GQouyr8xkSaEb82awcznkWr87TRuEdtKE5JONPy5
Y+eHu34utb0hHRerc6mcsGoqEUicXSvRTvAxrkH0ovft5TZmVX9tu5DsAHpyAIqW
wHNLIPX5owETyLkhKPntNbHQHrXYXCAa+J7NcFytjXoICAhEPfIMa36Kf43WdMmP
meeFv5TT40jXdOxhAtbUISvfQLwofDREWPED/avuD1/WVQQqCmTLyDLudLgh4xr2
uoG2f70XegNuy4fXmEGYFhVqkQ3n4rdEQQawaQSK9mak23Li5u+rY0+YD//9wCuw
IpCRefRjxXIKi2QDh0h+fA+xor7lsB+rjNGMMZKoc5fxXXWrQtq2a9L+elZLEJLc
moolb+gx2VeAEUrKZfXmV6tXSBodiBIfkilEMBvn7PPwnCoHkyvhHp7fjXAWeSEJ
e4Gl+20qIxMI0EOoqZXZmqBhARBQatVL85vkXml4IZSNkmQU2Q4qpU3Ed5YJaC+s
sNVrKoZHToL73sz/KE/1RYkvp/KzcefmaUYLKlYRfI3aj2X8EZ9Cn9O9edvQGmcO
JQsuOBDGk0eK0ztPNaJhLMz3srErQSXL4CGaiEN+ugQ+gQrUWFdJDVIxDoIAT4ls
d57xU5BD5UvrUPoA/EMF1bEOT9enrNgFvsSbcHCsq852nWjvfaWzcqUL4s4SnGii
aZtkyfe6+MBSPGhKgiy7KYhtswsHvU1e30ddKbPIcpDiTFkGptYuVmxHCeluPbJk
6DyG+j87s8aU7dcGH1wMj4L4wOM76vk3C7BNg4AE4NdvTvlG2RPqeGwUoW7FBuZJ
qEnygxQCBNlf15pCuIZQ9B2GBeWaczlT4x5wSljJyI7o43PqdumrEUwN0oqurJNL
sBkM8znU1CXa6f/bS1ycpQo8DlEicNnJoOD2O1YeGS/x9NcMUUnGrLYziVpTIWDR
3Ex9ymzAMDiK2AZs3T9j3vI/c/YQBZfOatRzyiIgiFPZgQid7x2rsN30UtBxh0GM
uBhhc5YfvTs/EJIUa2ADqpiMmXH+Ay1sJcxmeY/kRdgvxbnS3zQVHXE8Vzyp5xVS
jYf1Stt3Z/gBoMQ6bjWdGnw9NAbscjjlxSG5Do5PEs/bxNIS/tYT96DoxmQ9/4RH
2F3FCpX3zTY006OOaT0s5aoTFO006PuGS62NCfuBJ3ePP//y+za8t13L7G86bhhD
SVqiA/JFrtAn8WEZSYrmIJkcOv8qessaacK6voQ+sBCPGG2lYruUWz3hCDhSufrH
+UNNf+/Ksr4i31mbZ0RcnnWrHMO9RJsXkCop2Cpf+k+nNrXPP90aYmqHELnedO+7
xT3pdD53NRpBOb3wMe9yimEJy5vdFshxpIDlUJHsr6oHLED//C5V9O11Imfp8Nj3
GtqYG7iYk3pbqJ1cu28T0rPqMRgK4Ns6pUCdZ42sA5H3BnpNziTlg1xZkJICn9H2
oN87J8TEZoL+/lXKI/9kykkZMzpw0Xxg+Ov421YtSehbMOX6DLvsNX/G39ErfVTQ
g71isC1dz/qlTsA2s/eS8rTmPaIRYu04OP7U3UtH9ycYXNqI++/kf9aCNekliBec
4fq14i4BVLYbHRbJqg2+JTIEZhKR1GgptUWDJ6tC5F/NWR2COmvT7rMIbVy7/6br
f9RGWCQrQg7aFpjiiM9p39ObeoSvQ8AFLX/cIqF9VmLnCiA6FsrQAefZwZdeJLM3
ThD1d/wqLQyu3vlObWO0iOI0ko4N9l3q9VCiY+sTY6bEbBegQvMighDKMbJaj3bC
JGVUDfeM+OwaXQB3kd5gRFZKP4E0sPw1Hc5k1WJ3VXG0Mtux7LxfCRe4IJlmDqPI
A9V1MONmbyGK1Jp3qqU22pB3YKpjrJicnJzqlmSFaNJvQjiZBqAuMxspwrW8G/+m
Pde1VcSy9u96ntouDdEgT8MKbD13AvwrGYTgE9OKPEZEuOfDr5omG9d+RLfOQT26
3ihVbDiEmsQP7mBCYkf16eel3DMhvbG+vcFHc4jUgFRINw3FnTpusrB3UNcRyzVq
d/IW+WtfbNuHy8B30/uHdEiG7VtAwEXb1qzYLC3//w8+5L+cqnJM1n2LPyLBEiH6
vsTGmm90qq7n8AMhwnR4lo6bTdSy68WMPU41JGJX6J2REcb9X5OQkTJFzu94BzAt
2cWu/pu6H2jl4qXomUTSrNOHHNHptxHbWn/DHuw7wJyOfsJBbVerl3G6C297VabU
Z11+RvRHy4xzFBIzFS+CumoEXqTDQ/hajaAE8/qWU/y7mzJQXnoFpiPtup+9MTdg
Qahfhd06cWdmuDezZHmUtEiSIYFPglWubJs1pk+4tAoU0VQPTpsnDmHMSFVaQCeU
K1haY1DRINciX4UDWFkz1WtQgKPWzw3SbFBpydmoMsSc1JYZ/LP0YJl5+/95EdUg
z4J+yQYeXk+jR89FUc4r6TptdsKmjdJOsyGVVhGsMJbAWIRqCQzNeZD9eR8iPB6U
v/Sz0vZ7sPnXwxbeNmXmUEDEftHdAwYu7z3SJbZMIxGgHFp7YDYGO1dwdUisLVWt
3VQ/+UjE2lzxvd4hROHTaSTALFRTZjtCr6WdhPQLRGqMP2qcZIxm6PJXNB968crV
1VUNRmjetDGVb1Z61sSUlJVz7K2ydxbNRegR9zB+THNMMMLhed6ot/78imdJ5cpL
JVhMVIrBQmdzFjCKNt6WEfmCkEeRCB9q9W8IHkt7+jFSYSZaLbhVRommIPOKeZXm
qVEDLfzoG80Ow+qPiKdBfN1LrhFLoyDgTjiWbxxcqiMGIaBZfdTAi+G8q+KQZx0r
BdSykfKe7Me0kYguqZnJrkEDjQkGWF5fsUbIIisXMe2Rs3uoTJGon8NtbqIw93D9
7ByB/G5js72IW3Jmu0z4DVsGn06/5vSNpWi4FeGsz4w/ClxhWf6L+t6+o96GoIGC
5Jf27FoZsHFJF/c5TpEx4C6OehReF0WmtGjZ/RiKQQ3CvOtjXf18IWhzHthVfYIP
n/fgUiM41a+ZEli+ViTLohCQV21i8o2T70KIPXPo1bUYvhbIRrrUvSmL6XABPz7j
gZ1ipF6RdmVPVLbA57DYGNE/FqeVe9W2B47xZzDpCIqZ+hE65892ltA6kpC3WORI
G64NmMzFfF8v3KFvSiKxmnFp+iVTp3ekwSvZhMgaKXz3vBxoEP6zu/SAI73vkdQu
ZyvQso35nIqbO03D74zgm3C0NrBvYqBmgT4K/8/y62//eBJANYdvgFTDyGKO3URA
mPKdoWFupWnWTdwQgnHKMP2oksPd5fsIoyIr8WODFDQBVTKTWjbA/I/kTMhPJEwH
CegSB61/iTgsuuCLr1Wl2rlM0cwZypB7XpFB9NpQ2LSlh+lhBYk78UwtgukmCLfb
Zw7KVTWmfZiUiR37lJINERsaISE7w1WQYwebpEorFkKFtHg2Qp27/mj68EfUvT0E
V6o0a8yZ/V+3bB/WDpKzXYSHwbIpTV3/jfYuiShHKwEx1/Dp+rdUfORhArc3TSI9
zEvK/86hSGtENT1mGcCSvb1XHsjf36EivDRg80hwXMFxibiaHPtF5I825XUkTqI5
zBoHaJK1BwSw5Jx/c5+Hdv6fJ6+tDCBICXK8ltwtHQOBYVonCTw2FxhNjEzLhevM
DwxagjvpmsKbsRJOWuHj9ru7F8irRBlXTiO7xuwxGhdi4gHlVKEfRWBilHUxcj7G
ycBUZdqLAf4nAalA6ncsYaaUs/1GUtbnY2kOWjLYU2XYdDi3DuL6jxzPKHoj+Jzf
hR0KWQdEogxI51NpdK570eIjytAkMYly2yx/N7Y49cEQ1UsHWglYr8JC9DqP7eNc
i751Tp6l1Ff/t0tBboYYrZIXCxtRQcq0Lh7p6XcY2p6poKr5AZ2Z9CnzQ8at5W9J
wABS+Pvgm7oVW6jJ4i1vi0tScA5pFAzwNt0zIyXNoGPYooH0aNiuBbWbp5tLCj74
d4nq+tN2jsGXRENq169zTBdbBxGE7uEOH637C7FOxhre8ihzN9MSLIVLwpTkFleA
whQzeGMoAG3UZ9uDHFuHsTBS2eQ9xuXs0nVvKGTOe+KXLhPakoyTUvb8i/xW2Aba
4EBOGlrzf1o82TV+GHUZriI2ko0WuqOrcuw5PUi98SZOHNrhJspGyzwek9+eg5qi
SQcqg0uyYH0QD90wunZcQaYG6z2B71J0EogcH5fZnK7YdivSZXagHEAct5dNWnxg
v8dJq01Izxk/3fH7p/YOXDsmAn+1V1qv0hZuwfz/5qnSOBx38ZzbEv12p/oZrdfN
DWlXH+FK6Ft/aUdH07NMeVXffUgWClW9+1ofasoQHH2XPcLcgdrB9OWi9BBdc6Nd
o7UORlHD985USLwRvExNE49TBsGFENnTMXDpDeuzHJhr+ZgwXZa/YovRb9bOYlFa
XAROuKbSxMLdrCTb07NUyjv+zHHFQsA7C0lxgcw1HiIs0v74vaOzTc+7d/a7pwfY
Id5JQBBBIdnLqAbbdd7n65dBJy2jdDHcWkXOxAo+PQb2uUSlqHZ2QQsEnkgKoMB/
X5IQsNELENxUe02zTnUK7Vsk55Gkj5wfW/nXN7JiB8m57fyIAaWYxcMZfR58Cw1r
OKEwkO5t2m4vAguD2NdOgMBjpYQt6/OnHU6YZkKcRWIdMinvTRklJLsng8dxDEb3
K695dlv3Sw6PkD/Bz7R2/oP7uuzt8IfO2GNtpplC5a8nCO7rVLQzbNZccvf3Wcu+
MxJxnsp7c69uXlM6PqWIpleR27bnyi8KvZenXDolaupeA3nSnBqmsj/5eRoKGvzN
1rt2nh2tcJBZ2znGjUWT9pbMB1+bMgkV4Uv+1L7/nsop7jBP/LDctstxux+8mTci
CuxNcJjA+3XkB86bh1Fo0GjirHh53R6lEMCMfmE+AZyl9qMCDZRl5JiFuHElfMeZ
YhE6VPPjV6VaTR4gtFCg42Sw/vpVwCcPQX/Z7blCQXcPwApFBXdZpQyMpT5eqlwa
LOG4hZU0UzQ3cn34K2Imm2On0clq65rnIq72l1ACXKMeX8LNXIv7o3YrzVD04xEb
B64nsgXrAQ771ZBvctQt0rEukvnqKYs8WBdrgOkGtccj7oSCrodCSnQjIlByTbFN
mJlUkqO+bI+b1ogunal/w7XIt5aicNHU4eDqAthj7xtTGD6/o+L2ed4yHOK5hgfm
p2mvi0bYrZC51Iw7sbgGzc0iK7ws16ShvNklyHJnELG3PVIrmqModso8f9lwnSa+
IfqbvYPh4t4qmoP+708MWcb+J2/4yTU0cfFd1Z2D4AQcohwSzKCfLUBKvRFRt9VY
QBmaP/0NF35WdrHs2a/MOlilF+e0PVs60sRxZxOc+gnkU9t9MZFTm0CkwD2No9Zu
il49rqRd/josFMHVwOmljLb73lBQYIFCXhnaR/amaCNZzCiTcRYxbhdtOPWGptgp
xk5jeZrAo2X8zx28BEQz3qCxILiVJebr5ZfWOU88I0/fADDeRpnYw3gGGdwAbsY1
Rdp2FP0mIODBc7vfDjDu8W3ZoadPeqJDpkJU8+ojQgjf8yoAlVo/bkQZLNiwk0nk
4YvVO8ikWzPh2/r3lM2bMPbbTpG+vgAUDrxo0RDmlu8U4AEltU7jjTEXmuqZfIes
2Eoqq+7h4L9lCCp5kRApX34kZcZGp+FpWexrtYY0Ul0u1Ei9Z7UpmlGniUlY4LVi
iU7l7FokDz/3jon/iCBTpAscWQ3UtdCxZeLoI/khk5YuvAzAl1z/wOZ+r6gZTGoq
v2TfBr9UrIRpqNWWvWY9mGmOJWHWeB9WDAtqgaDvpdvyMGa5GQkWVhZejRu6kvzj
RTRuilt9uhj3t3oW+Ssvj8z6Tu4+EfpeVn/qS2r8JcISLzJFudxWTSnsqb8ESb12
8jXLpR4qOqhW2TyoYjZwo7dE5eRxoJcZkbVWwv83WDJjkU2qP8BQ3pWcV2YjEIdX
zqKf05I1qP1Z8fpd6jXKyQ5MVAUqqyc+UoZR9dlnaRvkSJV/rmnivkHog1F7q+O2
DjOiFl0b8tGOPXoxb7rIyizrnido+lTPz0f5MG4aiyGbKpt32YcJpdaI0oNROMxF
0MCs/SkRwUzaA8vsN9do8Pp1DZCGkr+ZlBqsDvDrpGl0lCss9lBUuFQHzNXDG4tb
G5xCwqFAfzg3yEfE/Ig4wf4BIt7VlCJrxd9qRzwnqJQxcLC+nMVU/rfGMYju22sd
9Z4kllz7tDDAZZcxz2/E6xZhUJsZmJUvFyBPw8wqxjyh6uQ8WZRXYEFsVl7SiF8k
tijseKegStwRVs5F/7y6x9GMeIjXRi2I4UWjZiCQHyMFw8tYY4kDmkSHr7GVkrUI
p9865Pni6om8zmjt3BLtu8cdmyWiKmewdFFD17F4tGYmi4xiBgMcstWisOOsFVgz
LdzHcTA+g/m4XW72dI5CMm4j/A7AtC9QxMsWb2G041PxjdVVODzkDLUyzKAyO6eE
daKrdrCBoT1WvjkmxyCjnN6CFzT6hDMmZzDO9q/6c9Gkrm5l/rM/CfxwdLleRc9G
fH8odeGflI4qpRFumeECm4VsLUCfm2aLkXY4RstDKIXke7ttniAu/gwAW71sF06T
+xpMbiFdhQZeXMY8BvHZO1wFj1Bu3aNGFdWqxMXa64EQEiSAwdFyOWQLrLlafVo8
ABQpfg0Aar3W5cj0Cxy2O875L+d5rqUFsiQxxotIKN+er9dT7XNfXke2VAVHRdgi
5NxeIVdXgXpGerE6NmLVqHLUqje50XQWz1qU/ks6t+Ivr6Qv4061g60X1DIPUeU1
rkGxy3GsPxkGpbPV/sBa08UceZQ+IO69lpXoohIGtn5KB0ey00tkaRNlsLak6OOo
k/mkRmAVNBV/UQncuiVpU7Et/fjzpzv/RTa2y/IDfbXjGXZ6RH9gL+Zz2Tk0PRVc
0ViJ2jPn8mI67TORLfs0b/uIhIR/+cGDMIpNPB8zuODoWJ3mlv0qw0qSgl/IbZvR
clCWOO3XkW6t+Kv8PAQkMcFIGGY1v6tiLJ8GTyM3NRtnEFma58hrlivXZmrkL54b
glIuvOkae1GjBMFhYJHa7PifacIZuuQVye0t+NTaUewrpRqE1N2P25S57GPV5DzS
q3DYnlXtHF1vJ69vVsmoCQc7YBjAj6/ilk5Ng4w0pOcwPwk80jEhNuvCN3jYYYiJ
tEcv/cg/QliFnpfC4zBSCKagvoZpsRl3GSynca7tjlk0WuM6rcUYV/W9iVEOI9pk
FJh4P49ziUnWpAssd1B8byJXiel0ieYmaTh8BVWeFVUtdPx5vICA73mPXGddcBjO
9N+Xa8uIvyXyLTK+3eLYGlAhlNmzs9kSkWgB4g0x5lN1o9rdiu5ag5DhQT9w8i8X
0seq8MyuBcc0CZx/ZbkSX2+UughZCqxCN+cxanfoiQY64Z8A3oE6YarPfXY8eQT6
awzRMkrM8DOpkbt/I0ngs0DQTYBLBm0doXAR5h6VXq0wkkQvOL4IiJHob95Ac758
mQTZnrvpdg6b3EIUDSso6RRk+041YTmE+P/GJMYUk2AJSGbRrK447GBr4Is4lU0b
2UdQh5TredNWVH0K6akXZI7tZtj1RR0yMUrbiYIb5coEMkbA/P4wk9EdpAuock+E
t3D7YghnVll/1fh8rdQWsgb8z4+njWmrC7WcSS9XFHKszRRiKkfXJeoLHjU+p4dU
0G1qXxJ7eMUeg6C8o0fFNoGFSja1ldGDdVUlODEzX6ms8A9KM9ruMvVT8kNWMvYL
llQANow6X7JY6mJ9E5Tnt0TVWGEO3zIzAPOOTtMBsSQxPibEbCl08ZJd1Czllun9
dEBKFmj9AecijaVBrUJH4hUG42IwbFqqBbOBVS5PGmkA0TvSuCwpigqs6xC4BH9Q
03JzEUw8W8vqpX9/8Y9UR7typqjZ0uj6zh5k2dvjy3FKd9rDdbCmiB8QtIEef/9H
Dl3oW9E88TLoZRuhg0n2XGS4whji+gREw7se0KdyGrmq1YlHZhsdw2a9hqCoDfNc
aerKOolG4ZSD1dXDPwCpJl748eRuNzS15UMHRJyiwyUdFIb+K3mEiUVf/jh7ENVE
TphWXZVbCLCoXxK2dNqMjfEtB34Bi/YRYH+oF5EC2kK5WgxIXtS6fWGV7/sPoV8j
6PrswDxeb4K3sIUGUaebkynZ6MBHjJGc339ixQ7WCGhi6+PkjBTHAUg+ocbpHuB0
2p0bP/WGZRTkcLwvdwX3zU2AbjxqqvGVHJ8D72wuPXXg1nHBkoYQzYQ8z8qCzHF4
9ySlvwIfBFvbsXuzVcwkiSztnKPMiN/dpQOFBNbiw9fnu4ASWGJ9TLBC8SfDXI0o
KKOXKMagK+wvE9HP7OQ7vHL4TJzGdAlpfRx5kUjyY2Aq+PjqZ86zSVKv3/vU02XO
+Z0y/ObkWGBlBG+e2lumPpcBsMA7C9eIIs58ZlJsHTh6Jl71lAV85c5vfa4Xl+Sb
Th4vBW1Yi7F2iWCS6F4b7Bh2q3Odpuwk/MYOGbad+EctGu6a+pL/2fEKSIUuU3UA
jUpylTFf6QziPIpoKACxV8kLcvT3ndsW3Tqj3KiYIDMR1HOZc1HF0v6bNQ+uvIsC
UtcHsVdbWjk9fmBdCTZMft08CG2lI6YfayrFEMt1GpAd2c+gmebWbJKS5x4rA3DF
f2sHeoK0xy/efxCGe1hCfUGUE+BFzcRW/rE6ftSZfDtiO1GFd4GfdyELSsXt5+kI
7KfeLk7mqw30iak425nG7hS0wGMU5ZrR3OpUjNXax/kI0GCfKimaxaOnd9pQXhlV
5DipmIKLHzepD7ESQc7/4ivxuKsogys1B9y/nJ1oPT9LQ+fsjwN7ovubWqi/OWNz
DlpB0bHXWUMFI+GrA8uzjVSBQIcbtX7jMtwnW1WMk/DEj940KiqJGIopl2ld8IWV
mueYByaIr7eWgcfIj8QyjYJePYB2Yat8ANxRmIqdllhyQu7nhQqT/omBYD0ga6bw
/sRuPo7b/SyIDZI8HIaY1pG2TOSxvSK3/Jb3SBwKC7SFZT3k31Cs4UwwHnX24gV9
nj7boWsRR8b9QHDNpnK2Nkig8z54KJPP5P6yRvGCfe+o9HEV3pt5L3WX/Pee7SCT
Lk6VakZsJnG1QQ8gwOlrA9KiPS5oJxG1L7/lWwHT3e0lMJolsgJDDoIUWC8BFXyj
HAU3iSDWiCDXOi0tGS0K+97MUuyF8luT6cd0UxY567E/FqqKZKUHwSDnhdfUjH7F
NUDmRMzMpKuaM4+CMJtwFTWasdyYpitfhzicrJb7yOS0tUH9vcW/TR2gBLztDc1x
JsyGX5ev+hdYdx3WhlPe2waOhe8JMMeZgJAQL50Ezr6bkQDm/xWGQdd0n47Dsiin
+gKfH+JCubJ+kUKglQdZz/DhSk/8YUqk63OKXi4gfvZcswp7HQftGi/515wQgEPa
Tebk3aWVyanOq6/yhYjpVZQbR+BEkB9x/Y3fV/BEPS5JTmm7FSinNnoYUhe29Igp
CPgDDNH+HV9AYkACH8U81RB8Lp3rmsXjw58DpsaBn0Kq34bxDa1aG35su9dEOq35
inRme/y5wHk3CKNWMhdJPUkbTLlPzo+/CPcEMX9bRVWq9MI9HE5UbL07NBeqQdF5
7Dd5kS49wL3jLNSysLucY9VF3j7iqslpJhJr2y5GjellLO8cJIEchUPd0nRWVkPx
Mtf/zYLo1vOkPI/f+vslVZLlvu4hOlkb9DhPChHgygWT3tr2jZSJ/ttbODDSvTYO
g0cJx+CK88TWXW1iXM5j7znGtdXXS598ieZkEEPobV4vJZypKa64sNVCBSOx8kfT
QAdEk69I9nmeUlG44A8Gz9D9NOKkicxcwgL/uyHJGBg9604G4Kua/ooKijPbhvwa
M9QgnzRiKsvo16I2KSyR54wzqyrFeR/KOMH1DChCFSq11oyZi9bTW4CmdKhg7J5w
/TDqOdRN1mRgEb8aO979bKu6tZXRgAVyLDLGTuQcGpNHn5xnRM6AGyBRuDfgsFV7
ZsCTSRY9xdqAtmsYlwQxPV77xHwe9gF7MtkUVBunR9xI0P6U5MxjwuLSB8vXj6ry
rvgRV48crl7U95Lq54rJz8GSfyaX28hcCN94ObCJd8iXJXeMxSk9S/F1HmagugrM
IkuuG8J/T6HpRsJ1P9WEnyBs3GfXxxQyj6VtkbYnZyAb8OSqArVdUsu7doVLOb4i
OCMQAq0LkcaNPs0wau6SfrDzDhay2tYQEEhGWOpwK6z1sofUoplCJBop64WgFHPT
PafxderDqUTxfeIoqwTIxGTlJJT7F8e7cQnbWGfbJsaPfqexB3VmY3PdUPQloFn6
1/6U/FjatW2/5LtvXDS4/hAH30YVu2myOqGuTRGc5CavBSw1Kgti9kgX+s0IBPIk
tXLQ/Vtgfu1+qzSLFfpzmYZNVvoEtuHI9yY+lFEfuV7WoZD6tBxXNNt+qw4Et/wI
Ik2RsXsvPdRYFe973Wrk7vhzEJ8tFsgJk6l2yiuHb9V7VW8ZYxJ/htu5t1tqmMb/
xblppzfn9iYx7q+IZASQCDR81xice9/1WhYnDRr0nZlDNKFYhR29DdOQ8jr9AVS8
UXsiqpoIksJnOuq80/yr+fKxklOmMT8Dr/XaIz2ubV0hRWdeWp6CW4QDqKd4safy
uwSzM9EYYVYKw7h3L6nvJiXjea0C22O3rRUfzPi7JyixgIvaMez57+jN/isw0VN9
Qpk3QViMUVir8dFwEr9Oyr7WswbgzLFNki/K2ltxFM7vyhvHToHRBqBoM7bQxGs7
Gqgx1HOQ9oYryZzfkjtOAwpsX0RnXqgva6jCBMQVDfh2QQ9b+BjIpC2iUmY6AHh7
rGR1mw+jd4sjhaRQjIg5Nr4Ru2KlZla/23ExebkQATcN5/YG/ZTKCKd4SeUDxJSu
hNyPhIAjfGcMybeF5JTL0vX+WBWpuuw+cq23i29AqWuQaYEKYxX8mfxRqHyjPhiq
ThwW5VmWDXfHWJXA2C0PbhKjdm26tIoaE5XfAqSZ6Whh0wRpGRuxJjmAooMm1C0m
vD06YAhXT4A8dftBOyvSeV2qPhDxBbPQCsjRa9ZyljEPlYSGxCAHEZg0m/qizFK9
jeTRnr4Me9AfJbeo4U9NXJBuHV3/6Wqt9bNPIm5HAKh3PDPKPr7V4wtmjNh9RXUV
nHaIlB39F7sXONKofUOzNNGXAUBjQj7DFSjR8IlICtGAmm63y66PQDzNeWVPYaBc
iQIwz9IPoW9CjzNsuNLrCZig028MRYAT7Ihp3iinsxeFFmgDku77rAfXx2HxTiS/
qDg/yBkobFPvmHs9L5QFjCKEEavFLV59H9XteAtiV2vq24KKIMpM4HxSsCGMOC4n
YaK7jI+Wj9EfJPWa7KepWk4siQjpSxZfKbe0AH4Yf34Z1kaHR53l2Ho/xHgVo/aA
QLhIiW6LAvXCR9KfAeYuP9YUkS/j4VdSUYKTAQ5w6pcip1LvufRbs+kEg1NFc8jX
6k+QZqHePKGFG0J3eUzbddyEtvbQLUe+UCR2mpZwj1AczFmodhzTUoLcm8ATKoP/
QwyeTYPPC8KWe4uqSYrcNsQLb+PLVmoAhWWbtgNn8mUYIoRnb4jC3TNFw1mzIn1N
abV7v2xi7G3RhXZIS8AZs365iEfvPXfub+gbhqiglAIzc/UfeThRJF9b6LA8dM92
aga8YpQlml31haxR1UJ3ApUN/1UACpqn7PkIxcfMzVFpjWvqUCjebskLgG16BjbT
+IvSLtNGFHte+8Q5utG8o+E5RnExuA4DYYJDY1SanequSObu+5wvrJWYv2k9AsMI
OX1TuPzmnDQ0/21L4XWuPHwg0FAql9x4sNtkv0evuoerZDr1int/i6aQdLVGwanU
HNqZm5tpEElgSjrwrqif5vat+KRPoFhElLLLNj0KX4puTFAPZnbx6K/wm9ETWAi0
3oYmsiXgG+0Sfxdf04BCS9BseFX8T8J+6x9Ff3oUgghj3T7ZDpU1AtNbeYbuHZTv
gZ4MlfABiNL+xPzVsN1qBjjSV787W1PMDe7WWxw8wS0/s2GsqkPPDnvvhee42aMx
dwySowMoYGEUOVVV3RLMfFGXIUj//lOJFL5IxK5QGjvDVl3A7IyqjBJWlxq1nN6l
KL0AKU7ID784407ez7bx9IF0eXkz2yCkQt7Bio0BTToddjA2/Ba+0JHMntfqxQAW
WaORIKlNGehzP1qAkFwNtgPtp/WBYQOkwqYDrK7qrc9Dl/A9QolBRaLpru5wi/zs
bVwES0zyRgDn8ML/vJ2wSN/r4Pc+ddtDkntQEYDTrw8Rtsd3TJ6JyShcozNIYqsm
gsS2vmjjJaSCtVAPspBbrdjdL9AEGQGs05zyYy1mzxkg8Ecx7jwFW1X0EhFaBa2l
yX+D8Bc9E+RGrGnsM2q/wNZlQfqDBUnl2qY3p7QL+fKuFMV4yqUCDBj82lewtcCX
dZlmYKMsgMuSIqs7omOuWv1zTAqgNBs15I0RABgQlYR5/qSsQg0ick7LwUtxg1hj
+Sq+j1OTcIO5iSW8WlNB6Emn10dsRZs5gfMvOh3lq3IgLBl1YDdHtQZsw8xuxn8K
PMnHFDDHT8aF/uhkkLsO3gTckCeCIUyniEAXz/7/O5r/aQvs9eGANqcgCnUl/0Iy
TLcw6i+kdVmc2+j/ZnP9o8o8Fpxs9CVU2o8MdKfsykv90MlosStr5LXeJyJWG4ZL
8aICj1mIC2FtHo1W/r4IBtuR23i8uRl9A08RQsnnwqJrTKVfxN8xBrZy5wl1v40o
068zj2F06IxmDeX6IKeYMT0dV6e2QOdq1dCd43fK1aRwCf5HeOpHT4DIjKtHAkQM
kacit+dgj2ir6Xh8nrRQlWA7DpYxl4oWBS8IrL2p0YxTNK+G7a30zb1TD4BWEFXT
7QHARA5P3lY4XxpjxO+j7+tXjaXgeXqdIB5+52CSORqyTBtdTB9Jb+haQrwzZPb6
7PRww8GcQ+d+VLmQruHQCvqWPkyia1CRlZVYzPtU2j024Whz+IEO9OLDSvCcCBZa
hnexulCtlNwje/ao4DH94RI+pbph+/aCyvzAh8pwvJQM/5pR4ez/DAWbJ2G6USxl
apEhYGHHwnrlULSb/wgW8nFgxIbqJyLBCMP5acsvcmnou9iDqKLtKI5qfhdV1bNT
Ghy6sSnETJTIrAm6ZjuAj74rZcVzcn0/Q8gG3c/QpkMLQgrn1Iej0I4Tfg7UNJOi
kF/OO/5QTsMVBzie/c9jC/OkwT6XInd6tL1E2KUdzdL1DjChkmLN64jPZKXI3qOb
D6wELJvMK7o8t6GDJkSMSWFdkaKu+Ap6zX2FoI5B2CXC+hnzcRGsCGb9LA3w6s75
wbawB30in9uj8qfz+stNQayd9Dbo6shIyfxDHPYfZ8gH3qv3P42hs+xTn2rvR72M
TKNRPAKs5PHvY9GGIoUneSEdysgbp1eeWiEpuAa0NNtReaIe7GOEPZG1soh3qSrB
uEFGGw50f2pzSF8qKcqmVVs42uLIFtVj6dp/A8udR6XxHWCseBZB0oWKwtJ3Z13v
IpZptRnQaI6HFMvd4MIUpG16D3WX/V3W5rwUqdmFGZfsJ/HfNdDkrKUK5M9BvO9r
cLe9M8l/PCk5uST99NwSy2Bi1TCV+xlvSKlyg6hjTUIydcSFcqu4D1WzjgDsU4w6
KqoOVVRZkiVuNvt1jQDRl8QVIH/9U63enndjYxM3K8WM1RkVSLcIg5Dw/qhjdfsd
Q0b6VfPHlJ8PsNd00VQH82Ozjk5nRFiXxoictK343smfSPrNjpBr4MmCJ++R6Oze
BtOf21CbPPZvsOx4riebqji5BXBjE5ZpATsBgeMLvfEv4nOkf3Pm+JWHNSEG/iqO
Q0P1eCngSPLDPERf0ExvZKvayhv7Hzt8Ae+rwTWPBE8osyivszEBLKmIrmRCLIEO
CWvPjEfhx1cI7T0aERywmq/UYFhmLrc5MZlSfhy/kmRz8WFypjIJQayoJGUPJ+v9
GbAhxwx22qGduciHjO6z/AVxJhdi1SZMewId7tjH+CDHOwIpNhwl2DtYe95eeCph
7uD11cwWZRPQ6hiUUb2bMN5Zc+xXZxGMusZGOOBB5eDxCHNWzhVmkOZicSMIl4dy
edXTytbJhefUdOuR+3xb60W7YR+sulyqBjs49VrA6/5IurHckCfUnXoRzI8gIDHO
xz5eR90pAqnWwMaqd59NPKIcl+CllmHf/eZ0Crw83c7wnRJVa3rwMwpK/Tshti7y
O6Ccz0Fhw3q+YiKIhg/dHe+UBjD+Od7Ga8w7c3kZssUn0K8DDezgEWSVq7qRaaXd
6KQ1PXrMGqbURxj5WxdFKGD7Zp9vQwDSRMknL8vJLCULa6Cj1aRKyqDowhb2dCaB
QbqBcL9vnYBhuAlCWHWMuXBZj63sYrRNnLYLxI5eFglqmPEIGy74Rw/O+pbWUWcM
LkoKrxDmwrjnfTR3wE2FMVRxpVmH6leFQwkTmp/ctGWJjsjd+qKrBTbCeqHKmaU7
DipE5DvN45L1H8sKSpyxQld4QURDnQ5XkkBOHG7y/bQhf7024j9B8VOj7Mx3DwKa
qmLfsl9ime+hu9YnW5M8cnwf+GLaE5X/4qUi22I2B5STxGz8CaIMyjR89hOhOIOm
El3S0i0MyxgGdr5A37fONaw4tMOR1KrKwYe1fIXgpWJUZX0s4BFXSwh2ClQeYxxj
N/6n+QHySUxNGEpdA6RnNDHQriClx1H7CjOLD3ipu1knay4RBYxOBGiEWZgiIpI9
QoPknkC/WTLwkOo8NYvEvQb2TKDmCmvw8TxpTzSyQuBwkqsdd4+okunBcsqVQIGa
imQO+P8KkCxcpb8kJ795r53Nbp1ZwGJKwwSmxVANOz+yIGkv4m9no9/QBsIb1nju
VHgM3x0vxnoZhaN0dS1qxeqWfYF84lGQhfOSs8JYyWge25CMPjgXcq0J1SuibEdO
K2ZqkuRk1Kq4vbdC9QyL4DhqgvmxMEkWD7MnFzAeSX897Q2V03FeURY5Ji4ZUcya
UBaU61vKC8WrgZxHGKuljEbXp86aSR/vWXdDErn4UA74qbN+SnRzIO/LlUYDb0VA
bsKWi3+SmKwHC0+FcLr2yKTA4nmTYOepUmH06ohEbD7+iDkAfjVKG/WuT9YKmdfw
7i/6QUOERvE/L4CBoyyaCCSaJBBhju4t4wVbmp8BGyPcDouwDDcXCwI5rqwsN+13
ZNgsESr6MWe96Q8PYCcW+XzPHugUHkwLbD71DIwEMFsP0Tqjy9SmFcPpfIDzXNgC
J35NYAzsHVcw26ejQPqT6wuNzfbD1cJ18MHQeclvq2f3ispYa1Agn3ERY880ncT9
mVz3E/L6nSLz0rmG6bC/2Cg5TdCo4SrUF12JLOmmclWB73ki+ZcrqZkSqVCOpnjB
YShuVBtkWZaRqaGBGZqXG6n1YNKquLPohAAJdrnm4LCoy2Q8sJxpmqvqafq75Un4
05oQSAsclup3+dMavC3bcT8Lq4ivWWJU/cpm9ADFvYnQPm8vK+TTyAG2Jf/S9MGo
ZgtlDueaJ3LRnYw9AFb0KoyVjeVkYnvt7nxHA0O8b13rftR63F8nYAdXVMu9T7aw
qFaaf4S0DEubEuC2ckvN2HPNC6p2veNizQYR48AfcUC4FWq8hCEGYYlSg8d7Iqsy
3Vwh2DHGHGYUXZ+2MErQahXLtMVzT/cMMniq50QmO+Qdh9gZkeLevr4hqxBzEqW5
DnZLlSSPj9sm1auYQ+CA71A6faLPeuV4ry1OHKdfkJWXMiXzRVlLMWJys1bYdGdj
dgQ78vQ7OOfWEeXxsMApFrsodIvouPcRnEUmGdps5qmmBDmh6r6utJDUOB1TxwEy
BPDg4e+I7KycEN0J3MgxVL5ug7YCg5qUfnY5KFTPnFbvTW7UYmxPcZi+aMHjqUhi
6nq4PBCCFd9CLKOrxu88hjv3oRi9dncXURr6AWOKJtlDbOuwdoaDQOrTQduPvtov
Wb/h1MjdAnoibmf5MV/niNe1jyjbhEJUd1Jn5sEkROJhs+TWBdCP1SJuYr1G2XM/
CbtqMhM+Jc6r9cdwcMvX6B/A6ElU0SUuewxmXCg9foQ3ROksgTgIPdY1PZ9CW2Zj
T63zUP/CJh9LkJVv0m1DxxKECnQhRhbAhOJ7VI/mpY0YbapjBnSpxt6TQtaZvSlG
vdUKjUvZVF2yAGxYSPVXSFThzFHQGfc8Hqqbz+T45KXmESVyQnTcUMBJmv5j/50i
EqVYogGy71r/j/dGo4ujXaCZJ6jXeh5gLFLXJ1bzivgfeyUgCFErGnLRPL7/oi8A
P41WjqA+MHn66oRO1+zDQk7Apmzj5LwEcnVOENlzHpwZbcF+ivl0Idc4h5xkF8vT
EY29wUlHxi3cyF4/kH6Gjb3YIAbORJTM8UbyIZtgv4b7L8rCqyHiFBODO8i2a4MP
+7WRrk+GZoyI8k9MF5FXl+pltp+Snp/DsEsp3oeotcHSKR8AUAYQrLHkNC+/8/zI
RaBGsPQY5eR53O4ytuOMWFN87mOqZZ8oy8PMbKVPG4knWFghZzh4o9u6zNy5lWPz
CRfBoo/Z6LXofLFSM++fKdefT4mm/uPON2ljahFjHnbAK3F5KSjXbpEOxnngO1Sv
DdjryF8zSUDLxrT/n4QQhh8ASOr0sqFKcG1vWhRdBAKx0mDZRq8RftfGPG0Tv9Fa
bPuCjdNnWeTMtkwBz/yFY+k2IDWR+TVBtvS5+D0KQf8VwTDa5uGeoOPw/3qVW0YC
MUPKA0OJZdzFkJoTSNL4Qm3qCpZgEA6fHefBwNRS3v396Tv1GPygBkghFVybEAHv
7ZNr2EDRAMJVWJRe0oOmChIVnNUHFpDTBbJQqXu3XnL3JRTuRy4UniPUzF9HA9uf
aV9iGu4PzwtW5z05VLjX9mAfXEiDEZArmkn10U/zYMvSet8fw/aCCvI6W6HdZ1qT
9F+b98at/Crat5J9TKhfKpNK9wDHfwRxu8DMhFkBLeRUT8Y2LA+pQbJuGZv7mj4Q
+M4VEn9lfY8Sr0eQwjRRfG0Fx69ctKY2V9lI388sYYkz+5zab32CJUe1loP7aDAi
mnSVOsqkME/REMGX3/raRwTV0PbB+1oLi0i2Yv8PUeedfj0B4gmc130Swp0DfMqM
GeiCPdtce1abaDPxJXAJM84lcBEwlqxGNMyHTEd54KsbgBFTZe1y1R8POGwCl2ek
/J7zHmSLSapS/NxOAHIVlmWQf9Tb4pSjqUHU+FrCb6DMgq+rC9iRzciEob2MZBNk
J8xpE9ekfqzjbFqy6Yp1KZaUW0a2TRNHKLjpVRrarU8BBNz/pVMUzBhG51JdtUbs
9muNxKyXUAgN3n8A9Jn12me/M51cC4R1wnjx4zCpsACt6T19+PViKCrVFh37msxd
XWsgvnj9pATuMICl5kQO8r3AC8+QOev1XVNHlSV6BB2t38OTQl4WN8OCMK/rpGlq
ia+MqNCoR5j58YW/LJ4w8IScFL5B+w3O7wxaT2UWsp0ImJjDqw2xrNSDYmhx5IK2
QT6jRViTEjPWPqvVs7/vt8BGwK2fLyafoHcU3102YhtoYXSkb1uVUhKHPBhgSOyD
KsALSLNxw9YZ0PEOJjsx+xsEaLTKaEIDCItm6OoeWejb5y0U4BYLY0m3cGsycgWw
I5wlNGx3YD3y0OHjVtqfB5dc/euy4Yxrdifp75dc3m5J5t/qmDle3E6RBjdsaGY8
dP/JtBTImPkU4J/RItrMwoLNbZ83y+IQtMVYYepFJSgYBeC1aUmiKRg322iVKfGw
BA63s9pvxbB1xzTgwncm+jnhhZuiQxCKmGqkN6AuZ4eGIgFjnr7QgOvv4Z8PvwBX
SXVJB1X935B0FIfOW9NBhbNdzXYjoZIhFlTsIMWkLuck9SAS2BNsUAnyqVhj27Lp
iInDY1N+S4crwcxvt5oaUf5zVv0QZdMnrL8U4Ihk/BPm7t0OcaYKqxItylS2iZUd
sqOqiNQc/d/8qrveEEH0YG0oTJCcqcCz/y/ESM8LlMXWQC/LVAkKrQKLTS/EZSgC
DHDAuNzdxtNPze5/imy8L/mrHyI5yRZSIcbuGC/Wftv56+cdW42kz7Dg+nJ5sZVW
pgQZqBAaKEF4c7SW9eVBItPk+ed2eJLvxTzsZMUw4+mEQUxnpOPeNYtMan/04t9O
2OTcnCG1sB0P8xDFGfYZtoKIYKzJWLlnpxMqk2vFX/cgvwElYs6GesQJFNqq1AbF
IcvPQ44OKftwZewsdfRLQfJONoA87NpyYKR9D1HxgVv/zn7KJ1m1fxOY3enuu88M
ZglerU+NO/XHp/j56CMq6ZpqpcYFrw+Qx1qpQzFGlA2gVmWCFoMkvoWvzPn1yMiq
oDdFEl1IqjSL5fWYxkWcNZun4PkTgDjtQGpaxxsB3RMqTlQka+61oJpz1F5qTfEn
DzkkMGZaHaTRlszx4PFkOmD8ZV8r/ZeEugadCWQGDQomUu0RswzHmSgb7goxeadr
Ug41eNzj2HkCUE2qKRMDWewxafqZAFXZ2xE2C5UIJPPy1erR+ajB43ZNW3A4fIlO
/Mv9wMc4jHCBcAgBDRpIXJV55kxDRpnQdhGZvw+JjGXupOCSdEq6NoKw+FN9rATm
ck2lWk6+o4e2DyJVFD8kiIx47I/IfBZ8VduGgQADSMKOvCexBY1K8khbuUzxUDpn
ETAWg1O08kZo/PJxC5X0fGMN084AZSEv5KTsVF4kFNtiYuVX0yYACHiu7pjOaBcf
tYuhZ1bHAbGVK5RA7CnMVinovmF5oG/8TFrjV42zAkANQ9OdNiHkTgCQmzo9UWo4
Pi0Z3kdYo32vIrRcP1RIQvtLp4py0ODyTs9CSfaJMjQOznDg+84Wnktt8f3QAARU
coXhb84vIW7i8RAWuT/knscMMBqMK8YBX0ylRqffSIU2p7RClh20E+CIgJuDX+X7
f24M66TzcBNql32vEB/hJZbdgn2DFf6ammSKCD6/ha9kCHO61Z2gKa7CAqgnQKoJ
E++q/IgYn0g3VKswSG01uM5BAKXaoWapaUbqqmVjSRNYBhgV64jOizigsP50cRCm
f5StgjFk8geHH5D4mGLHdHWP0kxL9QiEwuD+M2sJObgC2R2Zt6DYr02u9OYAqqJ5
Nfkq/B3IpSnCxuYZxnVaCkL5c19q+426jvZKg39EwrjvjRlH4cB4V2Wfw+5lFaHD
1/Eb+lBXsrv2mUQV0JHiiyL8Ik0sVyK6e0C2QATXbUCI19G0eaYVg6C8kOXifaYQ
lJkgAXweobMA1m6z0C5Np5bDe8/Dy5MSsNMOJbVngXWVFXLzEygOnF8skO5BMFNU
kIhpjRHZgLnzel4yTMCzSTWYAIvUUTqF25WbW4y06OthhDXDHdncK37JE76zZdXW
10/kBG6na3B6rpuxp1pzyOnmROSh0VjFRaxLnxO5ntMO+B7AQ6+4qa4j4pEjyesY
XucxJW/a6qYk4j0MxnZ06ZwWxoXA5rvJS747wn0fKPJ4tW/A2npiXu2N01z+OibL
u4Rdy/bUTCcqDtR8k8vkTraL0zm1/rZblYKDvjnU+8vDVI1E4l9lAvd5v/gheJYi
5+xHNxY0JPLPDXWRFGh99Tf0VK4jRv8QJkSn4avIBpIwTlsd3Qlxr/85rcN+pkcd
s/Sk0zl47a+6gbcUUi+E/nHPOOn9TALKYxZIwJP5sxadjrybjtz3/9vsagw58NCw
762FSeJNryUU/kQGFxravfXHxyUWVO5Ex/iWb8+pBmt3eBgXqOacrP8sj3g8ZK0C
rUxGWRDFsx0eXFCghkb/AWlcj+zVoVfgim/B5spRRsEK57HBlryVlcN85BQp/6Np
OKNseK0dOPGaIHTjsk+ML+WO3QiDn6XKrdPSSe+KL755i08ZH6NSjgPEypsmZiXo
iAZRyXvw4DHySYgurEEP2IZLzE4gPEnDvZE4UVAu3wUxohSiREl1TDqpeZz3Jyzr
fetAy0sdM4/2Xk2/5Ly3T8HeU1g4806aTvP2HXax/HNO2oQ+gmAxR4WgShI8Qw1i
jceZsgUbB8zoFx383QWyxNalZ7mqOrVWHrAFHhcKv++sWhL+ZxIeJXSOu4q23atV
MA3oFK2V0nnR2Qm1DAjPFbOmX0tYSYwVUugbsx5lhgsDV3tF9qaf+4fOGA3ZyKUj
D97BcjQ7VElLgaf2qqI+clfCKP01wCpwzC9nQC7ybpNnbWckCEulsjzNmdXegr9f
E9EQsZxTFgFXoDkZ4o7zwms4c+nccZwlANDagZ7Q27KtKgjNwu3QKUnWS9DmYOti
jXGWi8bbTeWByd2bme7kVubwoadUAn8zS6QOqogF5svKLmpiuMc37Q4aNnfJKsLM
bW8kKfKyMDnwH9GvFKEmTqefcoAa/KwhGYf+j3s3njmzJIWhiMKPgzrKBcQ4IVB5
lKUqL3lEJu+NgJAf/i/ycjceDnIURHlI5aP8JHdSn/MhOBER2S/vwJEUxM+Tp4l0
cM7ad4wn8GfxiR5xMk0wPjEqIb6wx2oFbvygF2MLFwZuxxn1wV+jn5ymhWabS3xL
pi9lWu89sIF9osEUnBhyRumw4mL0OqTjFJWu1jeZEdBKGf4u+e0+rVlBrr6cKXKF
f9of4VFALeCI0Hyk53zqbiyms50hibcuko1aDKxp1j0zlENU0mjIpvpK32BUjMQA
J/ejBDeIxxUFPTGTTsjjGicaxp9SlgJtJwz6nFevl0IXQUikrgTTB7ZoQP1YJ7tR
cu3kKIYLxlpUhY7VTBHCKeB1oWTxf/cq+RvWh4F2Df2P4CqJTWhhFJ/Bh96j3ZTP
fmUFGSKlCNy7WmNhfWRfAFaBMkSG70FC2w490Q2mliMTH5fGgL25NxywOlFRlKUE
AoW9cMSEqW7e/0js3VyC30iyt/ZT9UcDXwrcUqn1ubnAQvcUq9NcsPl9iMXU+vcs
rem0UrTqlfRcaNtqQj/l+r9Y8kFPoMaexYJ6WanjO7MbR1cauPacNO6+a2kiVouP
8XDdop7L+91aMoIlCh2YF0EFhx6U46tFFZOpLaQQ73OUQ1x+x68JP4b6yUaMdyUW
ZOu6O/ZGLs6+hvGR0gbEdKdV+gQX3XtANh44FGU2e2l/9VctEucM86MjyaCrXXj1
OFXPy4J3lpJCwCHRjVf92KDIJvu/OzvzGBsUNNqxlB9Z5S1TBeXNUK6koYd52JMt
vV2sLl81GanJSSWlRHZftBU63q/59gzURC7jTsk6kwRT+Qe1ESvYSQE1DdnYMdur
dEB7x0ltZfnd7JP4dvs1iVtau2gcZUlDNv3KMG6ljJue4SwHLf4uzpI5hjEMVZoc
iRIwWXO+qAOvt59tUlg2Q0q3McUQ/R7UNLCsY8l8X3N2cqrrAcRWZDJpQ7VqsyhU
3wQidQp/iJcL/n1t4AUa0gO9slUnlkfyTImDGDz4B4OXIzw7Th+Ghtdzn1I26Gkx
bG3/S64o4S0PHRFaiy3d2J+CUkt0/Xxv9h+VkvGYBwEySZ+QuM5XM+z5QaoE5xbc
pCb7YlShIeSnSJSFHfIC2PqRSfJcA2vblcR1hB/jXdNdRut8/4tIaQzCjwzwXQNc
y0NE6OdBC66NmGP2bM8oOw7kp8faIxDOH+vwZJjsExXoXRaKx1iLsqvE3ptyc8gu
XYj2cuxF3O/dvwwU+OM0l+IOL0hojVxMBYYtFHBs4AS5gy+LGyJJueAYUQMI9n8X
khkQClCyQi+brmu/MNgH9oqnMUYWVP6CsriiagcS/K/glMqbWVVYfh2n4sWdhTdE
Mt3otKo4tKIMV8ztbpqiFbtOBzTuZE8CMady6kFXloPdABvbrvCedg3YYdAna5WR
fon6jxr6VGaJgqXtSij6cYZExDMORmESBwicjjjVMunFYO9OP5ge21BAjkftkAkX
Yd71TtoqPizZeZ8OgAEDn3GF74rYfM6kMVlym2Zu0UrfQFQoBdky5IpoFelJ7zAC
0K0Mi7VkhMQG7PLlAJbjtiyssnbAGaeBPPJbHB7C1vJ/5A1TEqL3X6m9BBf0xXGx
nf1F41IBBbJvYCJ/S77KpUfTq9bKTTtTErrHHeBXRWnmj3/f2Lm+sNc65QDukA+9
iLJnzsizDoqld/kSUGW65NfQ3HpapOOoDRUtXZ4NiiRNVQkIGgVsfU8LhcU185Tk
NUafsS9ovVB4jabJKK/U654UcXnDbVYX1dp6pKUMwhVYxGZgj9FcO1y7hnm1Y3o5
RoqaC6Msajf6MUgCD+LrVdHMg8rwn7s7vUWweyElDwDembNpSntm1p/+BXkYWh1R
Upmh1APTYvRne1fWg657mvAO00VrrDs4zZJjQWC3lx8cVbb3Ynkk9BTlJ9FiCKOn
YaRFz6OeQ0eJ/sJ2TM73dw4UFp2W3u4B8dQWSMa+2nuongGpRX3lf+7YoJE0qY52
Wxm4ShIvKRx71RR+Efv1EEMtitVz0N0dOdslIYDxllUbCB4CqQxRR3DRUXJ7otmK
caSJkpjk1KislAcMhqGzlVveWAFQDrPX8DC/07pEaUv5vLFcg1gL1SBXf568x2St
sA2keL8edQ18R7OSugLUUtYRt9ZSIDjmg4zxz8r31mzn3gM+fsZAwxrtGA7CMOzE
ssjIFMXS3wKDNI3kT+l7UcmBcYhgDoMkV3eMjo8+m9Z7YyFJ9CUNMutioEEb+k2R
0c+XVH4TXDGJpPkfT+1yiLTEwexv7kAkYqGqtTG4n2H/0hP0Bz0dFzrvX3VpRQ6l
fH4AMNNxg8RZ0rQANaNMw1rowoZjzJNK7so/GKMRplBTpqXrCw+N9FZT+oPblkN2
SmtI4XvlPKkFKcBm4wI5PNgv25vvrqA1tlKyoawUrtZtF7aliwjqMa5I4/D7zMop
uG9sub9b91W4elgxMQdjmHeACMRxvN8x2R4eXYDsz0cVS1ERyUvhcZ8hJvWijg0M
AXSmtuxPFEt9yKT83ViNnfLHWJKzL3La4Kc/sK6jxzKJKxeH9kLDk9xS366paTYS
IOjZz7R8L0jEp9xoKtoG8xMMS/jKm4zi6QlAsL+rbW3eUJuzOK18mT4/+3ZzzVm+
Jf5DCELdLpawyh84pyLMZiXQm0Pwt9SaftCCylHhSum5RzUnJU36cO4JmYO6jebD
ZgS3sfNGsFl3r7XME2p6q52x1x+aWwXWyvmkMw08vGuS3TTVnktdapyEalTa9qFP
v2ukMj163vjoUX4nbHW9DLwtBHYdWzC135i0iLihLDHZNud9M90y/lU9dIWU8jK2
g5mVcPxUcoHAm5jYAm8VY9xv1i+WpcChLrVT4LZBOcsszSjDKtxjY8xStPgprSPy
6QE0hyFNC0wJLBLMaSqn+ouonFx+4/FuWDR1gsSR1B6yHfOo+Cm/eK7NBwXMO+Jf
n4RjwLkgip7T0ohfI1jkiGGCTogAGk5uX/tzX1mYoBcf6bBeJey+KteCwJd8fS7u
gs18RvyLon5JTs0j80BL6y7GmhOojvuwzaXGVr/Y7duO6pg0YuRqrdE9pkARzN/V
MNWtsE6CSZnVsHph43FsEeGCszy+6fAobeerqozpo5qORo4I5j334c+HQXaRBIU6
RaCsdy59oU0ezumpimd3RtdIL0i3AHzG8/qqyDFly16ohrR6fb2qyT0TAXUZsKAU
jISAd04DBWg7j8UtYrJThNz9h4e5Wc1/eQPLDr/F/HtciJbTqAPV6LdpxAclEB/F
e6A3f17uejYneh9OrXLRh3h5XLC6d8bG5WpIWt7TxhdfFT/Lh4KkkwkWcQtiTX8N
Nz7Tz1LQOms3/Ngc/3wDL72cVNGxYPD29vIP5iSc8FcwcqLEI5RbdaCo50a5tCPl
g2783iBkUWoEU128UKt804Ca+W8iojZKZvqhvdE6X21L5BDxShrpXCPwwvkVUrFf
QlznN/3hgkALIsLum05jlQKV9WdlNULlcmTeKci5PoAaJnTq5YZBLXg3DPoGdrxc
1RShRdrDrtXX/vF+ti3/i0XI38o/lP8J0N/0UufX6RcJWE5JZt/YWz3wtIr3Kn3f
DfZxRLaANQvvnQMhMKsYruQ5GBI/FSpSLQG1oFLTA0X1qy+ZbcPLFlUjHw5wD+kl
hMl5NQGzIfmHEmZQ0+UI3VJmg5HVc79fkFIQ7TU/QamjaFIkL/soHpoQiSSsH+F8
Kt23BJf2WOK9uG7PTakqVXnkMWzKl0/OnaJ//FWWHbIYTw/jxeRconuiTmrH3813
F4g5hBrrxHVY+ODajjj/5TLQk88qkIimUkqv2q+Zj8NR8paEBE9uQ0tlBUQ3k4Oi
RP+GXL2SBg9wE5JyTfh7FiLgq9M9hyjDhuX8r5b7zPvqJedmF/xA58Sp7ADcM8Di
UuXxJzaOn1VEzEtMIKNPeRuLMlUp77PNMUx1WX842vO5Bs9quX0QAy9PcZbmZBdu
kgEcCYoMAqIF+YJf58kJMzn6Gqb/+3b6VxLDCaDp7kzxNuL8Df6y1yzvDzHYPLos
HpOyyUNLN0t/sYpEwGj131CRRPZF5lZIvOg4XWw+EL6ajIz1hS1ln5CGQCIdzwzF
4wtlRgiBSb4QfsCiBlUs427dQ32/bOuSejOEN+zzO/D0ConpGeyvCONAYjNJkwGU
gvYoNvGoEEIJq7FZgdezo0QPmKUUA4vhcuOBk5C//tWv1dViYl59GaMJDLIvICGY
SNifFk09YoiHW7L62vsgLarTZoBQZ7l8XmeCRFuoYgfOzm9AiWH4iDIBQkCWurof
pZhPInclsQthiPIGUfsqZ+aAOk7wDDgMd39GLjtWBxDhE6pRwfzSprB+zDOMdk45
zlG65xIfUuTODfOnkXhqDB/lOAN4AkQ2B/GwJ4lQDc1Re3ImArieDHP9/W30JWUV
wySCo8wNzajy9WJh+J8lhI+IKZqpPwiw6ROgvey78gJmCgWZJpOXXZRUEOGaX30Q
GcKuVqFlMArDPdPUs8SiwMlyM82Ex+a/k8dExFGY4Zbvr74LRKNNPhjpRU+SG60y
I56FmU0cxjSHEtjH2ODE2b8NsLwOJVB6SEEtuFvW/SqJpPeFvvcZ0Xwv4hOlQ33m
5uPnIioSpPRovPbp2jSrW/Mb5HciCnEQt9dK7KsRhwiG8BuRqivYgjDzcf5t7vZw
qCQX4Onx/yI2x07k+xqe2IugvXs6r8z4cJKkc5uiUfUOlu5BN+xG/SnyBDYnBQO/
bCReGHTb0/1fbhqCXjRdXdNzwcT+yKqd8moov73XpRkRMfWHl48pXmFhJcW2w4Om
5WmfPE/s9G7LCVsHF82qitrUxegMS0sYlee5/uNvnPUoRhLbg10QJ7eemoS8/gm+
1VjkPZzMKl1KCxtudZjn31ZfZgTtPPSHQ77vGNHoessJi9WuoZ4sTDthbu7Fd4Wl
/Lq/JsaSWIl3vm5KA/6/FYeUZs8FffBFGDNJGv2iJwR9rM0BcQm5j9CFIs6Dc4vz
r9aFsPuzPkcQ0U1EQrVAAj2FeaGwhcgCbvMMMrIFGJM3Mu5l+kY/nuQobFkZadzP
SFCZXgDZsXgYnBoLgCH7ZYZ5b2J+0LyJbEzXlebxSpN4VT7vAmlOOtGpfSPTmnR+
pQj97dA4odCW0A9yEb9faXkFNENEK2LYATStnj8UBB2Bf+VKR9y/ORu1+N6cgmYq
/+tgX8FwyopDR8ahI5LdKcFGOimYk5WG9aFitdUYsIkwFFyWWugMo0bvkfJJkS0F
BecvNZbWXKuvssuUJZwchOhMl8B4cxwgDjIG5omeQBtb8YaklX28V+7K76rySjRd
ruhd5/E99CPtYKndxcFyEYejuNetLqXYGn46Z5vtRgNytZDBzGOsEz9WEI7o9O7O
UkbhUbVt8bFS6ODjbk8LDWQ4LhtsXfis+JWZS4Se6HBWrTdod938f1zci0d1u9wJ
usy1jkUrtfrG1wxdEgIQCy6TxoOCUsxWKF+yKTcGXXz5WwOdccWxhs0opp8wIBQf
LH2DgkMJdS1838vS0OwbGqWF7KH/vZtpRfc1TUC8X7uXpnGiGV0CIkn1Xg58vHBw
8iMclhfAL432lJkaQ3DSL2xIzQlKfmMO2gLk3D7uKbO/7VUs4wd/2/t+GKvRD7UL
mxc2nQ45gD8eqWE3yYM/gq6PWDiKbh5kdrToxRsiRGqi5rp2lw0pMti3wUkVNG93
w5ZtOKksvQpdjRsP2jF+BgTHcfh5RqUXUXa31GG5RxlWrqH3/S086CCNNAmlzl+W
Q1SaMUPQtVTfe96En4cjzXi4dsu64dreiWwTzjB/L7adoPX3Ap/VhwJUih99l9B4
hcFiSkOK0EZ/4yQmtkc1F0rdlySrnfGTwUnDjHprYsZinkB6bE3zR88e+t0rdMg1
MV9qdGbC2SPHnRuEvIl2UnDiE/BNJfBCZrfKYmmQLU86U8+ZmzQW2hFh/0vkkPq1
M/GkR05U5YAlyfxQsf1bO33xjJbvibdVjraIuVhFUU6/Iy9vqKrwuuL8kPfypvTy
WdhIMipfu5Xc9KTc+8oKmlBOxqpyRv2CX8bAVd4I/ywpw/RXTYTDhW4SsrMOvze4
jRtsxiJPVSR/9Mh13OfI2EhKBy8Q67zRnroyQ4vLQz3qA3CqKtWrGnjLkWWuTFAn
NNT6qOiO1jvcsiPfc7cD4m+U5oFRNqfPqZpiKGv86ZvBGDVSeKU02QB+mUZGaBTI
494k5RbNib3UNNYJtMDyO47Qzlwu+N67saE4z1px0lb37iBVCzzsPo1raPwPFRee
2yI8c4yD9zbIEoVpsOp3QpXixqrlpUaxxJoqDjewy50ClReOinFgyPLQ1qgk5cr+
VIYGzZ0fNxLxbj+Jmedf8pRBdcltqHFkgQAfSPwfyHzQy7idbV1+l9CcpWG2pZB6
njFSTwZ9WsK+TtcuwbU8cUQi8pYEMu1vrtHx98WZ+wGjOCa7mIXXYOQsuOKTYuOb
emKQJ5/C2hDr9B+Xs6F3Mpwb6lesGLxcB1sf7YrJfF0eFosSoHTUMymCeNGScraC
UaRorxijTWZAY0xkJk/X684MpIrcSxyubMpKA0ZibXdHToGJBvGwk9HOjJ2WDDGx
iUH3xVQ/A8QLpJIkAh4bfdMMZq2GDcVBgAAmP0nubEo7dyWafyGJypTZ/oOMcLsD
dgeDTojePV5v2WBBRF1IrAY63p5GffOkDQA1FdGr/fbGyEt/w+u1WUlqJtQt/Mka
j/cRDCTz/TVK5q3H2f4Vhko5vVCtcQBEnC6AntAWakhHBLbR03OIopYe2gDg/vXD
6ba/yUGijE5F8CLkPaDTzECq9FzyxhCulEIsVmz0lbHIbp4frvv/WtMd4QTGfMeB
/5u3aDLXy9eYtJtZb5zn2S2qaWlr1AIFG0gZGCQTFMmzlLZEk4Lu+rMdSYx3nM/i
1NzJ//7MioW/d0iCA6oLmRuBwdDx3s3Cc9KlRElgXywWfDBFBs7RHuPmawH1dHk9
r8p6paD46rYiwdoTqXKVAoj1xMA4NCgywkxUIDeEWl0nGxgx1I5k1Dwp2fK82ujF
U1ViLRRximWo5/y2pohW0vE7KyXmTLEA4xZgkaEiAAXE5zg6u2Dz6XbC2zh6181n
9NtIULRmeCexZrOpw+QnW+t/QGqRQc0KcmzuDaAlLC8soFkB9hloSUV1U98idu4u
FICLbauSevbZmx7sZR+ey5sTDtOf+PO52wtWfPNto97YrA80ywn6uSujajGvdHh+
0F+hFIhj0SEmgEHImMPng+tyQSkAcq61wy4Vf9qDsenmvCn/b8kB0mHWbj1SyxtM
XfsjeWVVALy6mOJLepkp3Gs1LVrhg93jAJMjc3RBa7nucsD126xnLU11xLAerB4D
eu+kyVZHtxEy0IH88vCKlJgoqt5Z0vT8eGQtxvgJpPGMOsQZV22eGCM5Gf2YWmx9
9gjYn0VzMogb3a1gDZmFpNzBzOuoWLo2BJrf96JkzN7bbV09m+dgOsBDOuNlvo8l
J3OK+z+RhPGM1LMzylKAbxDDrmrNWhw9OCJr5JHviaDzBk5qZ1oWSJMONJmp4/vL
DFUuJS5SSBKH6nQc+nv+DCtKZjsufmRAtfV0WgpNZKJE07eR7vIr8QgXv0X9rwAy
fCuj+MQV79vDtJQ3tMVtlKHuefLGL0/ryzkkJrthBmYwvHbo3TRVsnduEsbf06Vi
z8akzVOBAEtO+p3N9UxgkOOOVNeCMML6SOo2w81kuzB4uOHlCyBfo9iigBoDLxd4
OtdZovAI1nwNfg0ZBbG5wxqa0RX2rFA6/Ii3GFWwdaTvR+mu2N1ypum20zMldqfe
3f43MJPwlWB63e0uT01871sFBsxKC6La4V9vPfFUoPzIetBTYfcIgpm0oa7enHA8
xj1OTAjj/WVdQqad83S9vbxiIJgfgMT48oNq+mKZfYrI6CGlhAv6Yt+lzThLedT8
DAUwqwZ3PlsIXXSnWQWd/bCId66c6FUgYzsVZASkPiZMMX6GOH23E08lQch3FkDs
zZsddD8AXXf2ChEB9+tsOH2FxWom37KvsTfav2IP7O7cFkskXX1Sb4Ky2EnYPvFM
ut2cnpJJsI4nmdrvaEn7/W9pXN7MCyAkI3aoCEt7b4anydZuA7l9Cqw5yNsX6O2I
iRhYVLniXG4akfSGcjzL+Ge5DS15zsmaaiTzh+rQVcM5vDC6WHmMW5fxWHJZPi0t
B0GOdgO3bKq19BQDWTfIzF7tAeL/VlNMnTyI7HjP06z9Gd0o7i9bY9/USrTaiywf
qNvD+XhMHYnfjiEGOvF9/JBa7kMqHlVU/bfbTCRY8jjtdy3X15wV+f4Bquv3j7EE
s+TJKCl6RRew+rHYl6enRK3V6qAIVdNM0JpC72avmj6uDI1P9bR8vLqeL65Te8o6
Jwpb9J+QCLnL7UAk3l5PN8q7AWAbu3zanbE0eXRN3SxFRSIzbQPVK+KUyjCwNC1Z
V2Qke30TtvZVWLCMUIWadu5tHIwCF25plKy4uzbKerfA7Qvnn+o0xWViTnZx67JN
uEC7U+DGYYt4kW5lusDmMtfeFimz9Wjm5Bzsz5GwAJrbUROlLXEtVlWZ1YjPnlkw
p687S8kq8VnOTk7nvGpWVV5uw6R4eM8S41cdcTZFGE4gZUKxJyFeMWDBodMsA3NK
dMdeaVHu+KPNh44IRb7iEk3nj4m4Yi/ccxVMrrqcu07mtuMnzsVVmDVaDm+3mxav
dFP4134DwueHzgjBgf4ZT5j4NlnagDea1KWOxntTxCQZErPg+zEN9X/i2SFz7Yr4
0+oo6XsXKgzvZaOXtBw/BujLOGX+j0QqGYqec88/pjQwYn5RRrsdHeyDPxHS0bkV
ITimoyw2SDE+uoMKHgNQEXAjMtRvOrlUuJfLL1rNBnNl7gD+9C76zcVLdEMQhkfu
1OD+JnP3PmF6J5bNWo+/qCykxICVjuMTH4st7O73lP4wYUKO+nnQ/fQ1J168yxS2
ZriwRWaMWK53xByHtJ6qqW2I5ZCqg3nzXCi2Rf6D/2Izu6ButFfsV0INhgRGAnML
cR2d1pAU8MnnFmVmgzxhrjt6F/VT5vTcnywHYgG4fq4lBZ1jEWxAKmkXL7pwMoCr
wYLNucgs3ixLL6bOKUN/XUyAcCfT54/zpkWaiqHA9BUjeLCDFNwKW63VDpJmA/QN
nXx123s35SP2yj83kEMlwPZe9TfpoMe3ux5q2sAkjswNolyOaG/1Bs7HSjgwsc0u
fydxqL5BmXypT43Gn/dYcW3hTqZJfnxP5C02aGqwiOqn5D7wVhE0qgD77tT1jA/s
7XZ2LgbECQOzJKHeZP1qwDRnu8z5Qfixp5UniXtHniP84jmxXOD0MwfnkwKuEiet
79Pb1K8O0nuVp6epYBymfdDN07acNiaDr9vD0Cm53DBUC0dwyjkMsjSZh8M9cGe8
/iSv8W/1nNObTo8xBzSC4wLL5xU+cpmAGRH1dDUCw/cdxWTymBg1+E50JyqFXll1
qZ27uLLRHT2toLaBuO/ie5s9cVDOWxjK1gnnmKqzgbg/OjSQeVX52VpwkIsAcUMJ
vaENyBp2QibrTWCd1iJl6yyLBeffVC1XGjUN6J0wuIEpzL6lAb0oN8gRxzOJ0uTp
J564W/8QcAW3usThKdANF/9fD8PjZUlm6eDiEjlth8qgRd25GPaniofz5q+DVS73
ATL9oOrmEOS70m7g6PssdF2hA4edCJoE0mpfwQI7hs0pyCbiNaKOsJvbdybINV8Q
suIy80JPBNhlx0aBgitZfDVAicr4cP8sGt8gakifh+os2gNOHf9d1xrYJKneIFSc
xStADousfJ7ZPBWp67SqMrG6VVy0an6RSuh9kU8E7Y7ktb9cXukXEwmbhynCIeHQ
tUNQkEZAAnk47/8uwXETcZUKSbBhcqC6+fYFag+p66dqShfz81fjLfRrhY4DhTNe
i8y6vIfssCT96aAqRE48wAMW/Z7QPTeGiHqvDhxN22k97551Qiz+HuXZL2g8FJsv
0Aw33Np4T4HdYg0wYQla6vOvI7qANv8meo9vk0CpPaPz9atjtArBAS2qb/XN9vIn
3qowklXzUFOQagXm8arUAK5qiGHm9li/cTXAuvmtwxkWOJf7ENZ8bDLSUt2eOPWW
QZ0vb9hrGQ5KnFRfpvgK9ejl1k1XEuPP8pWN1lY209MNYBDnWdyOyjAhdV/gsh6K
8S8KPAHnpXNzQaiy9qjG8tNDtvhwiO57MFX5us2IyZzZFSorNG0km6oSAjXRTEwD
2kMoYHW9pM7JSQp5HDFuZtkrjD3cW3MxrB0q5dCYAGFVOk/NncBuYCnS4/L6UuE6
FBSE4ZAqMIhiPZwQgAZltw5ILbhRZruOm9fvEAbggDW8g0GMFJJq1D9MEyXQrhXl
BqFoJBkDQrhi/vkpt9DN8GTSwWtuvETgNIfZvrWWe+goBUyp+butgCXkUn4usYvy
umez54+oBHdfBdgsLBoaxY+EveFISXgdT3gURyguJ8ANwzP5scX6FeLfdhCCxLku
GN9QgzPgDmntc1j+8CCT3qW01bftyLVroEyVOvl9u4jr4PHRorFW/jsuzp/tZ5J5
TBio89B/0KZjRTVwNTRGwLH3YoV4OC0G+/VuZDAp5MVqqxoG/VqzgUGNfiyx4hM7
okShIifpISXrwNwL6OG0XRKOoUomSoOdkfJ5p8hXYIPaDdEAsxgYJ2n/1ABTkQ+G
a+MyaADcCcus2/TEc069Kw6M6KkIPp4hozBIe4OtYEPr+G9PnJsK7C0NQu50QOJC
O8pmAOok2cIJgVBz7NTC0pdQRiBRc7OMc90vlAKEYaugi5tXS5lsdcC33MHIlLqC
bAwdxyb88SnKTMCBA2FWHognrVlLhXqoFPXkdGwmPlz/l7UHD+MypwTXH8Z+nHdz
jzjqiOUjrFTh7My+Fbj1/whK8QNIkprWu4KqpC8OtHhi7R14RAXf52Y9g0sV0AeK
8PzI3qknMdIGu+qn8pZat+Zrcj3xg5NqgryD7H0pXeKsYTlyu+9LaKYQH0nNl1xp
KnOozYUoiI9HFEJZx/ZSirTRH/lBFgjkplPz5WhyfrQg3I2Rsc6YXocokfFsGJtp
ZpPGoxvVqS84c9fa3IoVMlYDGM1TyvQd2bxscbKD/l4v8K0aEi+kAq5swy5absSF
cOKLHalvdPFK9gPqOQBOC9ebdv8eVF01l/maKZpzez2u1WkaKnWzVwQ/Z5hl0LAr
wWJpLFR+8bGxN1ld2Oy29D5QVfqrnAgp39dA31MtbYY/VHU5Zov/Ks6E6DuBmAal
UIqhnYA/8iue1b/PR9IbR78as0zZ0wvxm+2TKZrndtKqwEumdBdJd6hXvIZLjdlA
inXI5b++CRRrJfPReynYuQYd84m0u+x59c4vo96NjTGEQUWHpkF9ZnWOkq0wcKZa
41nVZgRBcY9CjMPNCHeBkMqKymHKLi+U5k4AIdnRnS1RoVtl+4M5JJx9TBcl4Trm
y8mWHUOABj9z+NPxHLxCzdGjItirMqPsT08m8cUl1CT/q8R+pZAV1bKYuPn+Dxf6
UWaHmbtl7nhkQznrL7xqVrgaOZ29Ejz3NOWZamOu9KJudhTX/Er/gi/nRVTyWeB3
g6NgPhOZLK3KyM+cv5TU7RE1DRj8eSvQyiyAJjQtLRd5WBrpKnBW+F1dl87n66jM
+O/YvX4k1O5fbawpccsC5vkWwFbZR3fSkuShWN75HuFwnAbV/RiJ+mUI7jPOgE6X
K6BlTfnkdxYQoX2lXsBTg/pACeVKNzWsPO+ifMECO5CGmyMll6qkZMIdSw92EKGE
2us5opjRcPcc7fee9uWVxEeM0WMna57u5IhqJG1caA4PhpvCGV/7ALPSMojy9lBz
RL9jyxw4KowbaRmrxlZS6Bg9OEvEim08uEtvGqiTw0vi543TYUPSxsyd1feNB4MD
k14t67aHCYpV/4niBDTeEzTPPg9YDZyACCRXPrgMlXyI6MCg40j92VHrIwgpRzKy
Q/mvvcogewMUUjkBbo1pWghsPlJwMFtWtN0BGDe7H3nP5Ua8B53koQnI0sGe6mjb
l1UoglGVfECxpTNbPrZDn0tl/lIM7SGtK8lqqUC/DPqDXEBUPRqqguxH4/YHD27e
z2NpUFhBPHULKSm5rzoi/iVF9Xh7b6MD0+dxHPSavvZ8tzYd+9Uo7x1MuHwzScPH
8yknauPURB8+wvQ1nz+MUCobEyOc4XfLdA4fAYPI91l4s2TZySOyxXyPJoNAinqN
TumuDbg/CZ2dWoTFHw85wTC6cQThu21FxSNSwyEsP+hIT16LK88E+vU1pMvbJ29F
1RXacbF2qpzv/W5+xDGRLOAXCUI/fFCfaZD3abE+vic75+iHgWVe0/Cs9dFi2P4r
bw8jdSUGHaPqyBLlAJ7nz6L+PjYzPGlTZj5wrR8MfUOU7JCg+J08OOcEJ1aFqsz/
rzKXrubtOIg+t3Fo79mW48M3evXQAGcMhGpurddagvz8CJYCd1mUmZGrLWQulW1i
T6U6koLBBUjx6AsodVpV5lAehNs0OIAKqMYJIvuFuxKWBwEiC6KI/d9ocjFJjPSI
V+tgvqUfZ9QVz4hUjDyYaOA0vUbUnCvt91N3Rrl6naFznU0O8bpWOtDHyxhCAfct
VSfTylihjAdt+zJFeOwBtWigRUY5BhUMn2LVVkxwWX1jehBw5mt0H6+ShD0ZrO6Y
9fE1NQqtrpxa/H4E3DtHrP24TJ7vMnOGi4hNMVIua5uQJvztN+FAaJCz9wMxYupl
yOca7/xorAe0F3kycxYzBxHoDHLITPSmwT9JN5FflgE+mUnz0dMhtRJ0dEgd6I7R
Ho1RqYBAJHHQS8UAHFUMPBUh0M24VlrE40GLXIwGPj/BVQsb+uBCAfoRxXXqAH5K
+soPz+NS2FETIVz5bbzIlHoRnLwvJfR+jpzkr29CxEdM5EIaFzbFgh5wPXO919/5
if153VREYF+6SmBkJOEbOcaSfCg3AsA+AnC0hQLhWBQ0q9Dmi0DCNMQ59fMqZnJ8
S763iAAQqzmYKGa7Xh8pevGlKkaN4PxDEP60fyqWDp5+QXd4riwBcY1I3DIsUQ/6
Du958duCNX2KeTQBoqC2oaw84+QhTo6PI7G//UXs0LdQUnM4iId1XZzR7feV7J/2
7KgKbiJa1YRkuPyP8wxgRutrUPqp80vxnApmuwA0INJt0fbbetBs0R2j+MTDyEK4
/gkSpy1WFY/qWUfoBsq/7Zyh17EUp5GIOLvVvQ+JtLM7yyoUw6a/WlzECLAXfvKn
UvWAHdXvqTufvvexveylUVOoSd2ZQDqFco40Or48Mok238sJb/vx+tk5M7Pw8JuK
flc1qNuj12W4pfDQan0O97TAoLyvM4cckhTjiZKED32wmJdBAsFFjH5iYqlJ6EIm
gC1ArqIKfidwEnPPf6ljRsaLNyFMCwEFiUg7otSY2qtnvp9WeLPzLU5RiM6XiHUu
OFpWoS42bRuSVRUcPIgpBJ09uF3wzmLYHXSrNuJxEQHVcE1MnoA7So6SVsPHATab
cZ7rgWpQHomoWBpclGdEaQpJOa85uQC0Lg2/sgRs++qOt8cppNXJjRDKzkImX/gP
zBZckXicm9HM23ApWdqZyO2nPu97hPBX/NyoFsQrO4G5FWZvvz4IXV69czTGyK9M
JJ9yvBXUzUQC+eT53r6GtnKpVuqu7kGvOhRyTxGCVemImXUil04F9Jkt1zm1k2Js
g5cuEyNTNGLukwfMkaNor9JmYgcVKpqgJRBQd6QIS+NUHhBPVwBAmgasG8kzCmWA
G5JP6/zi+CWjqsNvqFgWBOhZaEV+mFCK3XWx0iz0ozYpmJBZh/eN2MbN435QpfZd
8taxQqVqYdPx/W5SCAhaQ/Kn80GLGpPfkyfeqotaVbpRTd2KsyFRCBG8oGWf+8cA
traejy/kFTmhXCHKdi4G7oUEBts6wXH2thtCVIsIlDrRmbPIwTFIu3Xpa88nsxBr
cP0YV/Yn/Anp4EkT+0wKsfp3Cfd2S6x0C+7JYv9B/tEK+LefFY4FjQNGr3gNxgUP
nW3lH84NBOU0PEOsz4XMdn65Z1BFeJ3jfwRBXnztBK+csIGI0Zlwe1cOmL3pUdz9
/8mIsH8LLwkO+4yLUvmmRamUYmwWawPYeFhIu5io8ersyY+SNNcwNoc7ooOx+yto
PKJUkQeo20441PUsvtR86Cio3yQ2AfyWnC8F7U4FMCm9e0rzP3zmWLGj9NxOf1gz
yzYI0PKZUn1HQi26Z8/CMZOT6CcArW68SXC8lzjJGF3wnqUuwilXHrXRRt7j806v
5/LRO1v/PamK1HFeVIg0ZQuKYokOVHtA9gef9SjGMaEjFbpQjs23BudxL/U2wlfV
5o0YIjG4w+SI5cgQB/+xDlV8d2N8i/ohE/ChZnR3Yq46hNNJcgRTbuJaWaqEBX2+
gh6ROTmnQA1iSqt0XfKo7GvgzD6m610/pdR2TiyIIdoNmAzn3sSKsJCSW+hKCXpT
FCRPPdRTqloJAmVx0Z0Of0TOJiku3GGEugx8lyz3ESYEOUWuAXSEjWH+oWYJQSma
Dvh7DJ5mnFy+vavaP7MBIVZnr9BVBdGJamwQkv+Ue/FildQ2f7ONbfoML8yYpAl/
2yKQIfQXLCAbQ+QdAQHJQVy3lcgkYwki+dp/dot97ljWudW8/2K84YA7TyAEAtoD
+cpV+3bsUPRfXMZqEfnNylQZGSmdz0Avv8OlnqWqGFXU+ha8IfLeQ7tMbFb67AjA
0Na85hFuttQRwgWIAHZhxnfPXiT0xshU7EhkmaUNUkC1GuNVUv/tfcr8w9ak/BgQ
o5qkGGtjXDC2uqPjvNpeu+P8qZFvXiarINQnpFQfDERtRNZOHBUwpo/Tj2HZiMZG
+8+PQ82ZX3zzjRu8EIOhlw2Szrqo25mHJ6DfTmpPC/Z/TbE07D7hMmVgfRXuNPCv
lnxMitMlQVjaWHQCB2mIB+xiHs0dUbmJFOTyydGmHQa/KfTb1ERqS4BIRGDm5K9W
3/jOTfghFdu3LYdSgC9BuGFnv/jlN3YwFY3PBFtH1wVLpKoyBj8KPVrTDJ3frB25
Jpkfy9/t67oWef1Zes+80ves7lY7Hc+Czs9HEuCMggMQ1uC+Olz9YbVqTz8N9Ons
hcI9+kK8St1dcfx2pD2LWYw6pSUvkZA2HOh7hIWvS+pqBUaQL2BibpDvnQCi+qlB
Ms6vh49l+M8HO93ApmnKPungcSvOaZ+wL2K0CxD4KewbdNkbtMiw70FJ/2Vcasdx
gkLF3+Yqe0DtzrVVIxKrHiGWM/OZ9Ws7DFmL2qaRb/tWwUr4L0tbCglyWDV7F4Sb
b43HgOuZt+ERHjkYZWluNXrjHR6pcsQ2F9HvBQXq6FmHSG0A1t5HrBKQMNEJaRif
0rCRyl2r3XEWfYV9TmoK3UPvKaLxbXram9MXq+trKQU2X2NnjPHiFqlPh5yZDCMr
tgZUt1B+yaoI50gjMHEEl9ABm4MJwUK+6GBtE+KE4YV+BvkCbUHTDxSULg2LfXyS
b/ydPjSLec8doAeJcMhxhfBZXGDIw8qt6S3WNmShpK8Aw8Lfbwn5ZpGPjXDkZEtr
fa7Q5IDf3PPCaq/viGAOVC3ccQfUfCH4Zdrq7cZs3bDv/SThgsWRedOnxalwDFHS
0IHlkzf1mg7OLwujtz6iHfzuduFjZ4VQqfIzHQzWE84l2YAzJ7d4Asge3qentOvZ
5knDgYz5sQl5GlikQxn5XkHt74AUjRjVQ4rJRF4z5VdbtP5NtUXAZ1sphcU4/dk5
oI7ZISxQ8NnvIhPVUrRuINw9wspMcC8vHuXtmqrovyZx0nNWzXs6CHunoZikV5qC
+oO5116YAL/QhLTXsb+8LKDGrQV8Y0ivomNEp8MSfvWuYUxsG50SQfsn5e7K55Yf
x2ztWhLYCmAqdg1vVS5c2JRFKI1Egr8qFNMSroHu+CRqJeXLkwHuYdMQlf1H/NjT
iK0zdwyl0Sz7pcWSc98wk5Xit7+86cB5EqlU5Yi++MZ+NqtdH57NkVgctdbPR1wG
I3LhYVGpuEkycVHw4vSBqf98OfgcKz4Wz07M6ZJBo7HlfMfETih9Voiw/Wl3j8lq
GI9ovBSqivwDirqMjgd9EGWcpDRHAfg3UNwm/iLVAFEQjn9lkyLhp7nKTHKaWyIZ
Ji5ITrPDvJX5bMFAQeLZbW5vPMwDZhuasg7yZ86UcmHzxPrkjwlVukUGAA+hcxgU
xgJrNN9FZDvNi+eWulPesnGKTQlu4QOXvzDkL2UWI8krYpP1UD/YqXI4wueyGUvA
jmFf+6x0tCGBZbbvBftzfDuuHKdcqq/hv2Dz3+42vRfwL7bRHIwc57Hh/ZGMFkfK
pUaI26j0htz3Rc9xzX1x90P0WbsoCJghW+D5DMgKbVyrubKgYcYcglGGIavPb4JQ
da1mBp7vt+eonGSsgDVqSclcEBhmWR9xYBeXdrfLSK0tDR3Iwqf1xjq9bzvCV9jx
H3mWbLH7mlgjc6qCPpAIEPb/icU5DUA+Lme4Ewg9F0HkvaygObazhkhr64OfP0bp
Ol9yXR++ZPgTrWR+IuN0LJssC8gU9oKWLcQAt+jqFRVw/VSe058sX0S+cFhp0R5L
yLy9FNleGal+ulFo71/BU6e3VT3RZ1v3mzN1xEUTi8IaP2LEcJGBDIibOkgiSLJx
MuAgdcn0lRy/4GEN8QBFXrX5yg4yARriNJF53i69swEINGFjmZn79C09LkIwBPGN
5bzz+hOjc3bs1pV0cGkJUMLG2M69ZVLt4n30eMjBsowvdbO0Z+QmL8+6fWTgxJgC
7CGzzeGUepNl6sBC2AsNnz+kAF4/nt94DORX2soQSQbMik+dzmm3c/I3/HGjgd/3
d/KPiY5ZCmAORzGzaDEq4DTzlKQXH26EzA8yY2/HTK5l7z1nwVnOwyz0jMpEwq0e
jpErOxOLMFfsxgSGhmPcFzV1cA5HpX0BADaLVjvGIWCJFQssr8+RUjB4FSQ+Ofi9
U8P9HyX/oeWuBetn7RLrqUDBj4n3jS8uHqd0ZA84QSyNaktyUZSEfLHQdg2d6rfK
raE3W9JOfUANu+tEHTpzJYs9z++1lp/ACdYUSyOpSUtcAUVni990NwQdwMJJ8N6i
EFLfdUouS3wRjXzdw1ODXeOGr3PEaWPqGrmrD0sLMv8OPIlgnNUhWx2k5QuRySz2
+Tl9ltf7ZojJvMdfwberRSWNyQOhw3gIJdY62BPNa2OBOVsGCnbjJwY8YTmcaiUO
t2E+g6dDP3X3dYpA8b57ogw2yr9F9Dr3dKZoWaIn27ajwZmC0XgWvOvTWVSF8zwa
E43gXiFwwP5+4IuLsp+U2OMRgO5/xqH9OarVVwVIHp7fkJGuJgPE9hGDTk+61joA
RVf7uoirIlAsJ4VFJPxj44/O9vSkQSs9p98Zm5DTJhVv3vRv2d6agc9m8NLjFyfh
fvmqaYvMkbQaH+khl7lYXAbQHwGSX7Vov+823ebxXCjWR5eF2h2TVVd5JVSMZus2
IV34Hp+HsSzaQD18FsHawjuECnf7ZKfTFtlKo/hNQ96bZ1rrcZjIbPQ2duJpmcAm
V4sBjIDjMRhyiRgM+cJKEOT8lnsK89C/41/okFLy0uY0ItrUIRiqGOWn1YIVoP0e
hqpfEtZC15Cb7WMtxnAie9Z7kbeIgtJ3VgiasQnU13nta3vVOI9vJNxmkMpJZgeb
BqhtBWqN7ZrW/Bz3ZojJ/w/jeq/T1tlWXeTYyKcjD1gnZ5D6L2jOYBiK0iGTta8L
Sal16wHE0trizWwDv833qBBojY5lL3tM7qcwPO2mOSTkDNd85DxRs+rDVGOncEUk
lFIWucJSWqYuoBmod17fwgm+2UBQ4QYxlg86+ulv8SLDGn5S2n1iZ34g7P1vFycL
gU3egDydDJDIQm8ENDvgNDU1r/sX2L3W+X05nGRyd3bVecdDNi3H3S9bk95FVuGP
MkMJ3AC/qACLNmdx8A3Y4AD9utqCsfd7MvrRP01ox0GO8/3HNUOnVZ7qEO0f8nZV
JtAKoS4BvkyiMx9OPzJuQRcMZkzyotTXiX5SxzJScaYTjume8Mm2d/LkvRDMFqfM
q1g89uCoi+pjaJ5hA2tXNEiYtnmE3TV/v7bx3EYkiGIrZnlFtVg90HYTnv6RU4lN
G+kpSLvk5As+eaXqfK/CpzGDKj+YW8Sijp+/Bb6faUs8kenX5yBD7CCZQ6O7VRxx
FYensXR1/XW7uOhOhtCWG4XQgm8fdec//rlu3yY0x4atTgwjDrzXm40vtbCmxenw
7JLr7o1WTnJZWDhjtKEflXX8gDJfbPb0k8XIpIbeUGI8S1EqMz7mqL596eLi8PjB
1wYk70A6BACXYuc4ZifVDGBvLR4lGEq4EFlnaoxtcTtQwgGRyx4saTumgDLAdEot
EQ0UN0nxwATPaIr7GpCS/xETRdtLcnpHr3mbY+hlAPe/VjM/FpzI0jsu1KoBlI4R
4gA1OTkc/9TmqmjL1vF79WDxz+qfGPx0OHxZvDcdY9TtnDNSWKHt11zqL5o+2t0/
p+Ni/xwxJg3JROQhPfdcyeg2P3hh4QhjnoHfiRVMrmL3pqq+b4claa1UYDtRr5ag
KReAeMxyJdaxCJFPAThHsn9yaPOdcBT6ek/4rDqCXqXjC7FVhXBS0bYJDzNFEnlo
O8ajoljBzk3H7g5p9c0PWXJ7YK5PD2ctf6oK5jSU7RYGYEPRodYejbMrEEQMaiWW
JATYoxPhPutsGpVsvslalYDGl+ioO6v824V5pzjwoxAg8VkKPUaSOXNVD9+jQ6BO
VzZheTfVaxz2uTddKIfUGDjr4uPyAm0WKtLCbXKywIuI/xmssfesNHZ+M236xxeE
1NzD9XrFJjCWZ1EnLdNDvT0YNHEDt0dWV13cDRp4ebvt6xqGRGsr4AitT2fPhndz
f2ktvcV9oLUAfCc4pfnmdMy1PSvT8LZ7oBspHxUmVHpLz8Mrsh6ZFB5WAVIlSSpS
GwAcGLR8j07DVV3kJuIITBkVCHIEXAZx4ZNN18AnoTJ9T1w7+40E1MDEQ2AS8Qgp
SyeOrZzDL01hYWuWHi1eTcIRvw8HpOkDyeK9MQuYVy+NGRXGotsJ+pPd0SeeRL0Y
HJe2nLieMndUWUm5B97sRlsoAXfd5OAU9HtPGYbPLH9DP7aKl/xJX5Bz1A7wPeVT
B122bThZkO1Vn0w6Oz1wEO09+P6sy6tO4wfoz34T41oLW1dxo55Xe1j50KkxktUN
NxKCee1jeLA5/hVIxLEMT4iEMdQpSE/SXQCgjA6zMv/Ngu2FbA5tRJFuFnN6WsYS
6dJXx/M+rreQ/x0YcBh4VaiC3VAsY1s5TY7aBMQUH5wvP1wLc5j2pBIiViBBLU4w
v7/IL0r2WW9660L1L3i7qXNUYTReildaCZR5Cc8OzshI8s8yfM/pZYebaiYIFLor
SSX79vYDdjdL+NCdI81aGY0ujTDK80Wb+kfcRblzZnIuclixuIureJr4rWkeYugh
lnjSvTuft2GkcZh+N9q46ofrZueAxJMAQjhW9kh/GAF551Kxo/M0YyDiqVnzJ+nA
PYmQLelA1LfVex/dNmbWcAwyARk8mjbGhP6U6hYkEZgZQ1zdvCAblYIQH1wiPTL9
AzfHXxCzoqWjPFVOC+d0l6ALiayh6lbagKbsoUWepJSNdljmYF0aHCDQA3oXcE17
9ai3ijyE98T+GDK7pyNwH4aUOBJkcpBXvLoV+N/II1E2E0gbRzDZ5u3cEHuNUF6V
1pR/IIY7WRdR+t0bmOAhgOpXyZfIkYCsQcHVYrnJ/9tY2+w5uwzvnVywsm71e4o1
nKfnZw6XjpznuuA9KeuY2ZWn55mhiGoi8RomZ2eMw/SAJVutgjy3O0wEHyOaChQX
GATJhBBrKjil7yqylRgWQPogTEor2F1yfRQZcArA0FG1jK9VrOTyW4fY67w0NmVM
S5uEeemJAJRqkgtDW6Zte29U7v4vHMXr9MEMZo5czYhNiUY/W8Ctc8EdsMRpgmvB
frKjkAzJv+BYYn1oyz6HxRTzKGJIgaKJ3y0DAtlPcCvzCcP+lksK1fDE7BguZjM8
XsOKFZzJtO8FN1KAE5a0Vha4hl3zIXFZ1e3n5EPV9gMNBh6Wlt2ldH5QzHBHiEcl
2k9XDFjZOCjgjN0f6P2jKIFdymTqlXo/m+Oy+urxB3AK3jMt/mao0aol+vSzq+lg
H8Vxbr0kl1LqpBCW/x7sfDU+7rEezf+o+DkVNf5e008XU8qais3TDgiNRuPotwx8
Oe7hPW2UAzXIeW6FDDKx/ksNEBxqx1Pr+FPXLKQp5l1dnWrs5GPCdtl0BWleJx+Q
TfciS8DFpvg7OVi99ONtBrLl8SpkuGPd5Bk6EXKwR83gIbHA9ZHAHHmRRBkDQjjt
E5kQV6oS3mlFisvLnwjIERVdHLk6fSAF4BwqUBqKxSWDLOq5lYQuQU0uL4OYTrNn
60BQ4SoFfKg43z/qBmNRoBXT1HltLvqqNrscfRGY24HziBotkxmUU0Swrz5ivdfs
cc/Ien0RtsrsCm22r5SPnk21hNll+qWueWl2ecEDQ1+o2YNMPvDzgG3mVG5i+iM4
iCjpmR2zar8pcwqHgeyvsFXEsdbFdGNCllxiDYHUN4xyZTR884GZXdj2lJEUkDac
zrcvARQsZ+wg0nX//1LgAdIjpqBHbpMFoiTCW/YSBEm/jDQX3+2WEvU142XAKu8K
fN4UFVlOGfwXjZupWxxmfdWrUwKZtJjsAyvVV8730/bcmeSlsuYzIGNODfQd365b
H4DZ4UUduRursTlpyVPuhRaMktyWX8xQg4UyV2juDFdi7K7xm084W4ZyU+AvyASS
Oy0ZXnOGdhIrF8S9jhQlyUPIgEyD8sryyZsQL2m7HfLCL56ISCs6JULyzSWeZPQY
uUpnwmLfejCUYRJs5uEAnutYqYIYT/uogv8UWNmxGWssgGUxPzdRA3gzBI8luNJ7
GVqRVQrqpAAVHS34dDAnmQa7+351QemHpeG7s/sxk4u2BLouG8LbtrGXB29jOkET
UMkcw5AbhJ8t0m1G+UetngQb7Rs0tTc0zYgLl8CaUDlNYfXe18jVqW1QH3r5x7Rh
FjOPNtTsJWpW5WcJdd578T1M5venIPJaChNlDldHJiKOha8pVTCtTJVr758z5zAN
vDzEpP7UCqinA9GFYDXVP2XkQ+sDkDDTooIY8TP4xY5rMwKT5a6nSLiXFVz3hU7q
VDzK25DMm0igzQIRP+aoKnc8DKq7BRZwxilnwdERzowQY2VpRA5UO1Ji9+MAmKJK
LFjMagSMRjR4fK1cZQFJvLUp3Eyvpf7hpW+KGCRYl6XK7fdWPg3QAZcVBk6gQxuy
Cnx/A6EthHuE1I32E8C59qwp5AS1ciLCZNquhr523J7a+K458UX22D7bYQQHQGeF
KyYMw5RiJuDbApqWItNCUcEyLrQQVurufOHnDik53/mzWURPdnXD5jJLMEdNYIsY
KhADV4lqxXalwoNN2FJwxkgzRA95SZKVix+Q4FqjFX4H6Dne+ynHL6mU5m4O6BzD
oqxOPtCjI95dwOOZQq0rxUuUMtH43HDdjYhoAB2VVIXpp6bsTn2Idm2zngauM2u0
Y+xn1mcOO+2kVV4+gpsyNq7jOzHUjD3ehoMhRIlJpKvy0ZrzaVPuyyeL8KJaM9Em
A1gwTffUmQNY90wT0rifQsB2mfAdt/kJ5VTZH7ivPBXy3BOk29Ba6oWRCzLf/xSu
cESd6/VJXdDTOMdouWxtOsUzDW6FnoyB8+YNrgx576KMF2+AVJGZdEqIXZCZ8h9J
tX6h1dyvshPtEYGfPi+PYGXSAM50GWJFJlWRbyQhGCQq54YOla1qVIyMdwn83iJ4
2DOWR/4TO6rc5x0tb5rBH8zt3XHANopocwUDTg+OX77MJGMUhxOqb4tMWtf9UoLX
4g4n4DjBIjjZbMMz8+hYmtdpSzDxI0p3zhXQncnGODwHjFuPetc6d052ciezdFwU
wafL3EuHnyCdppIzo4OQ+Y7AGrPa4YatacMgJz3hu15y0VaHIjhOzph63W7fobMf
FzFqgWt3biiLgNbWLTrDi0wtHLqbmjsXxxY0VtNvRVRI/ldhTiM+c3x7IQAPv1Hm
vkrSMhsbtmv6ecZYMtW0zTTmQjMDJGPXwoB2uSJd4gSD0J1CQHkw2KlIIsjnqsty
VtmB0FB+hF9t2HwZrVDc8jwDiANCucJav9mCXwv92067qEFqfsalR94Zkl+YBbdn
MExLGwUpod1S51PjN1IizM2DjgOfORgTidPtoX8yWvGXdHurwEEkRlpEuD8mwVPL
WbP5pk60TTXr2Tpfontm/jxOH+r7wbhorOeiGEWWFgtJ28NGfNx64At9zu3sL1ug
FJs/CXuwpidspiSasq7NOGG+fImFBTmad4vTn5CHZC6xrQ+OrjcwuS5Y5Gp0JcYp
iICuQ7tl6nMaEy0lKsgXJ4DXOOWZcWGMNgI8mDJNUVxmnnAFixjcBwD4mCf4J5e0
gdmzJhG1sSnJvtRZe11EGapGTSm0vTgckv7r67EkecG5+y+1NgdmqqsUhI1un5Pe
noaa3GFyZw5RhtSfe1gkMND7tKvANZWsSwIMMQ/fZpSH/iicIsBa8LTKEtikRegq
AY23w32B5lGsR43ZWydxkFlLFlYlcdoBGEFohR9pBEF/PwWhf4y/IsYwgwEM/KJN
dim1Ou2HjNbq91evDX4bDNL9vrnRpEkbL80J2NCBScmkBJbgTMu+ich7mKxpDFEP
eiGyuCy1BjplcDFfOG8uT2i45s8Op1SXOP4g54BKxzRpV/yfZX7f9eOPAG/Kb3Ix
ANjhVdVyssd9q7O7IxxXADZgESwS5ky32ULDkOquvhBO6bM8yHzmnqsYojUp82ry
9yGavOi4l0LmoH33h+DYGd98kkYw2xaISRi30etFJRvowTnoCFblABP0wMDf3ZUL
h+trKhzDRGF4yf347RyiV/Nzx3uMKglR1wDV9QWDy8Ou8NsOql+oZ88znr/J+ZZF
MkbV/uoGBqiU23yt1yDzoqsTFKSxsbVOghkDef73qLnaSS3bha5a2cNGYvwj8Zw+
U+Qz1HWbCPC1nQfyv/ZBtgaX99AEDQhQCnV4rCHjQwBboDK6n9EU9kMgw7VFqZtS
wiwNdKVu9NQVa/CRBLhg589i7pUB5mw0xJ2iHiJDm/5v5nV8uqNWWx2eeH36xWUR
Ghgse1YFPiNvL4qQcf44/yMNAnNE7+LZlFBEXXh4LMK0BncYuQiruvdbzVZrcFat
3oh45vWItKhP5VZUQe3WuVOy2xwN59r7WxdDjAhblnTPgsye4LjTRiktfFm3KQTU
t3jOGKNAGn0QFeNLvDLUOU6A4MFtIemX1kK/vTJhrPQoeZcBSy09xl148u9xwiZL
kv2xXmn/J+1Gw0t6bxr+bQ67hs8CsZ2QZ6VkX6PC+neHyyiyn+NilVYcKNkJ1OER
5bsija4JY29BjV+W9RoTNp3RJ8EDqPYR1fbz9WLJRT/ce1QlHnTvbQTqR0ECZmZa
S2CXFGvlZSDwomZ7lMM2XpJGspjttWOXvy3x4gomyG+UCZGddCF3Ko5V2BIPj7no
mFpbQhRZrFLe3HLMG1BsjKIKN67ZJnQIs1XP5Y+R8Dik0cYLsekgW6Oy8hgHP3vT
59a3eMIwwe/fEa6ldBnwEuBL9fCstOstymgRxw2WRDoXqoCRcHAozgcZwm0sZPsY
va0yDjmmBteNvAeMDE+TdDnU8dnMG1S9RxsuZJdVhIQiiaHVa9ujqH2NLbZghHfk
lfM5Ks7saL7kK0OzuL8UeH2nMx2cFgUNyyMC/AfwIGk7MuJUMw2GJo5z2V6xvJQI
OVpvSS/n9DdmxG5Kfzp+7oa9Lk1oOjnHzzn9XY74vdFwBGvsRBW1nnuRdbDhAKLm
Jp1hgt+KF7B9AKyeHlkEDPOokE4MSmWJlMdn4w2h1c5xtXI14H/ZS76uVNiwWQmv
3pEKFtZUPqfn0kk6yo7IYkFBlv4Y0IOOVMEYbuHxWadBlSfbws1eMhUU7eRywLAD
7Q/cqhl+DoWM56fJeyWCeOCOt6hlv5iGYBI2P65DCKLA/jclwsuUgCFg6FRvIDZl
6eaMM/1ecoaQJAfKATyPYLXRKZYTHMJ4WV6XfHNnzTOpCFbS8WWJcXkF7lSnU2t3
yReCB5PF4fOGCPHhrwHhiOBYJ0IbZrWZ8TDTHEdTFECXzAbsGIbdO0LujJrpaAUF
wehFZ8kfoCl5Ya35aVcgagB7BZPLnMRLPRTzjJG/2+OQin9ScZCfYarr5r29fUFC
Mr7wfRcaZzqFL0uoN9PRLHKWPnjfsE4V5edOTkTvxouGAy25IxnAzQS7QAFpffDz
pi3fl0pVZ0RPCoV34ENquXms2edlFyunzb3wHlqcvKxNh7NfEe0Nl+kmemiDgZeA
0XTZv6qQ2kaQjb1YJ98a0Ai65+La7W6ly36klOa0SsTkTfilfC0PDEEURAXfvJpm
dwOMpdO/2ToJ3/aCWPSVN/XY3Db0sd+st2LMI87/MmeeZR4DHHllkVhQK/dSaNgH
9/HOSW+jyjW7OeGoVFrJ0yhSitHwCU/tE9ZQ67YdfgRMUzwnI95bX6IbnP65l+3q
LPhZKOPoPphts8p/EauHh8vYzl/OyefWQ00MfB0c03OvQol4JXNgmeNQg5fTrxYa
GXp9dnHKYM+IkY8zXMyCtaHrUOTt9my4Rv8l5l0g86hQA6bp7cc9V4mbeFrMCg7U
5YVHf8tMjgA2uAwyXm+MEQo/6H+sXh+oNUx50pFO/KzwBMg2Ivc6W/7K/AFt1Vbv
zsw7Bh3arWOKIJfJw2BYG5tEBU27g60z/k66XEOfqWitBFP/iT4izOKmCrlcPXSa
BdsR7Yei1YTsbK5y4KTdClV3u8RREFuZIOudx9qN2BTNn9s17wy7w1Eqr1+OiXJq
8fIyOwWvLWJDKjt+dL3mEzsfKjnIGe/dGocmKcCsY5hczrh4GTdjZGlMGRzpgaWs
vPj8n6/f+b2IM7VZDjtdqe8+WSOF1gLmFle69vd50jcvKko1dNQXwPXw7EGHA1fa
2qZbLsPREskdF1NoD3qssk8fTQezjSEthgbTl+WurXkwL4FjqRRAJ19jlTlJxde8
vI5N+H8B4OTz9CvU7Z1NyqAVThhPKZH7FMicFxZYEsTbaphZQvQKPvGy/US/FouZ
l3iU+F6RkXRTQmt0r4RBzpzqgissWZTZEAIwIICVsBy2//dmPfXv2ovgTAPOL/yQ
lMqkboxH7Bsd4o2UGPBYBUb+gzgVcFKYwxbX+CiQYUwNwykKVy+1sV3FqWVk6Whz
peV/lFrKTod3jYDnXuYSqykxpMYgRJW5Qffy/7s6aABrg1E00i9c30cGsUhDiAaA
vvt8Kv2xKzDHjuTfYbRuCjdKzrpx59kwm7uxoxu3qKUWpIPzeUAOQBPxgjnqLTn2
FGZvI4wVo82Z4/qpbIJ8PmJf09QA2HNr2ORoSUxJrvjRr0FrUDvO+Y/Xkfu8NDjF
2WUoL5uTQviduH0qw8u4AKM/nt3jsquap1xjU55WQndo16NHRdJc2SVBYHPHoDbS
iTWgWsh9m7Y9K112PeNM3pOvDyB3sPO5gHYr/bqvw28q/RmDDqPaVG1Rx2mDQjSi
9Hr56hYaX9JNdHIyWPOzbQbJi+nq0dE2q6uQ1xguxVHucPvHHkg+3FxEbdHG1uiV
+uCHrOSmS7PIXFDnZRP9nkl9CB5auyZ1q/A9BdrxE8LYdX5uTu9FTggE2vIgQXn0
lW5pvR1xO5bWFjoj9gLIfg/ZIQG1F1c73E/iHzePoTJ9Icbbs2zPiibkADFolLVz
DGjLxSRtLMANQluupjT4bf8jkANQhXmJmhMmuRN46M5VjiGbosog82WCjp3K3nVW
qS20L87KoGX6qJReHUd4XfFFpbGLdGg7buif8b5jSeTJOdSp8xb2JAgIoMewWQi4
nXFIq3ldwo+lFRO6hx3RKjbsO2J/4eN4qcFlEnRUzNydcMXFLVMQZHa487qoNgHz
KhDSIuy8JHOFgneXn4S8YSTXsaAKsx6pEH84g37LkJbnHw/tHUzi5crSOEoyBaXH
jdpYKbqyownkx7vJn3pH0Z4oyfhfIi2Gx2nVH+ThIpGcYQ3/HAz+0FgLocBGvIXN
gXiz/UjEXItLDI9onwL7CYrPAtipwhJW7RR62sx3pXHkimhdP5i8XzuCs310M0Dz
uxx3sdUoEeRNoASsKHTk7KR7nlExMDYKXo2vk+OC8Cou5yj0A5HPiPVZw53Bxw5b
fx9wkIBe+28AeuVmtcGmKfEYrgKtJg2cNUaJiY7swAvqqEOpTecwRcc9rJ8jaehG
zxdOG90shldQVwwthApaIqG8cDUhjXHshT7ZyTD3d7M7nDyThYNQziJx9sFpB7l2
uLYv7CVJ+w88KwAUrCtd1jVScwy5GJwuKpVcKij71eP23lcoEku4Lu2BhYc5WHUR
y/snv7YytDLNke+Z6T5FusBZTOpZwVzPWEgE9q39NhCDBBoBaQwUjMQ1FH+r7DgZ
MSgMfily9iXUN5Uc/g2c5olRHz6uH1P9n7Ty8ARfP2CH1luVOA2rwhnIWbMc3LpK
saTyipWNj4qBHwY+kjPmW3A7gvtrUjGRF+d5zZfM1eF0H2AA2sOCYK07sFQfbKt2
4ejk39IBS33ozq6fPoLksGOeJRbKWbLE0Bw9MdKkcu9NCqea8v+BsGm5WokBDfa6
2iH37OpnEOU3gMFXE1AEXDmXt90NuI07UQCiz5uk97chnEHl33EZ8I11e0YeAAPP
3CyWq3YD95jH78OFKjvmcsYatyx32vQF2ZzJ2+5X/RopvXHOC6YkesnZgwESpO1S
O3yiCTfc4PSQ3MY9+kfl18zaXQAIQSuHBXNHP4b5xMJoS0/G1YrxWcBn2IjTe1wn
BOg/DnFKg6GoVQvH+sswbRwVWDRPNvMWkCAwXMFzJB+xdpXPCFw3i0zET3uirFDS
d/D795Qp/lmXNLp6cZcwXineoOZNpvR44wAYqPM89WdWVlUuJZDE6U3iJ96muCAs
3WcIc4pYekGsJfocSn+u0NRoKvPwe7R6FPjPMDhcXSC1kOrkuNu4mbLucmLcVKSS
DkxuRUvEki4xGfBZ+uThofYRUH8Jue+LPxnqVDqZWjMfJmJxDkgD+WPwVeVsWGCP
SJsSQ9K3XzIaCKJw/2yeryorsmXN+23vG3YpWXFFEjhGal+nss6TbCtvBkZXLXKm
qgZWcljvRNVYx7VIiELVD8qN8g713surmOwuUU0Clk32ZmGwvMcKXITtzAiv++RJ
TBEQwfTVOyUlinhYh6dmpDb7nU3wf2eU9OsB3NF6+poHuX+64xPMkX0j5pOo/1Zr
oTm0GqZB5nfLSHaZeAmQneNTCX6K7gnRFfgK7ijtoFoBB9nWoFWYQRnun2ewOLEK
G6pia08nwXsr3LhZUY2lv+zo1yBVclUQXyQbBBZmY2HFvulqZ6GmR2hrYEyhtH5y
zairBqzQ2zpnRwgjK9+rh2BHgluEcGjEXkRQwWK7Ffkjd+cVLf44a5wWyEaBJ2hO
RVqjTSNPiCzLwpVXsKWELSOUb4Hpytou3MV+xj8elRfh/AQ31ex15HM7Aotle18G
ZtODMPgpaoHjdb3HABepVQDOlKNc6g3XX0pd0mgnZEOFo0HqmNFbUJUXZaM3U3sN
BHCqNpa4zl2TNbRI28tN390ubsU/0zCjG61ANSqrSZXQpWkA7075ss2Ovl0uWzKq
kSxgWFPOzbZoQi5y3+mFyT23GdD+6Fkmo+LJ1+MgatEiKWXqpWmU/UV2mW90vOKn
BCzLIHn8lJ8v1aABrCp8rqDYX9NFEL9UWSeH+Wz9s09O/Iqp8821lRDwRXY+2ACl
Kd+1OIgZk21cKsGt2RxpHJWsbfOTMPULkd73t7goOd15ukTi3T5oav+p0D5AETZR
95Amwo1mgKQ2FgPt08cInyqAjc3umR+4ZxCBapiPZiYdWc4BdJcq+2zHrd0HrIOu
bXpT/pgqXItfmhznfw82q01ZlcWESajG4BsSKsMCbE8ctJtijMRqu8IdKj/sA4/E
LJDrAzpjrN81J+MSYXSszWmM+YNUwU8JwJHXwH4jNQv2t50eWusp94eHtd1Q7tKA
2AI73Uqqct+XjRKa31hbQafff1L06uclsQwQAt5zKYlqDsMRFKfRTnuDRfUWTavU
qtqoU2XejxJAbkgVQzE+ThdgNyzndhcCDD62MMBE+MA+Q+IWz2HM+Tuc42fREBlK
lO1RK2NZydauxx/Eqx8u15Tv2ekbDrGNOoiRzQVWs0HGOuG4SzF4pWCA235afLu9
DoEDr1f5zGCbn8DYYhvSSdMiUH3aZUOCyLAZ+zvXugE1Ypj94k60ysTa4PyO8tO1
o4RpujbfMqfjAzOUAQjEB42vcX7+OPnD9StwIu+lG0PqLmYQ4r4frJOQ6Kzp93MM
IR9uvept/CZOEuJ+sdvnklAD+SEgEGLKJL9G4aHDNhZDK+ZVaAd5RpR/YgJttjeK
qI8at6qTcWo+JGERWi0MqccKvcdgLPoYG0ylyuo+YLS5fft1FzZ40Mk+K9lCy6dH
HLo+0YLFh3Iyd8W8OAmt7fSXSZ3zsbryn2TDPOOCgy8njQdXcxmuPJBWZn7O4Y/H
5+jYOgXe4dBqdtUYwJdgKm6i7vkij+1+av7PiYpfscEQ792cMM+9/kIpKKGfwavv
POyXq/BF74tSZ2ph7vkfRQ1Xqex2ogMKRYoH7aRPHX63pBYz8EAZtXCPp1Zknehc
O39+V174p+lZUOTyk5s+ucUHqLE6DJUFEV6S64xiGcqH9Yk22LLDuS6mAGLkOT0U
8bc1mX762kCClCE2WAMtfN1tgFCQGbUPLQdg/WzjbCSDQxyLlXNOJND2kjNOGV6V
ASeNUSfjbsLRlmXkT39XehONBBxUl7EjvRVAcdulz/LzU2A2A2r05uwMD13Lerrn
EceTnUGTPB3LWWHtPTrcsDWHs9lci8b7e1bkWGFif4ZHH0HgvyaUQLDbUNf/cNk2
7KRB6Lthl/K/a3B988XWj3D6nssDCFoNUmNWnMhsTLAoCMRtRasX+TdaUAMhHmMn
nHJKl3x/B5e5Lg6VEgOaQbx/Z1rP56Hf0Qs4YX0umZ+lNA5M5Ym4qe6LaEbYRCsB
Dd5fxz8vU8De2gDQzPAl1VZ1lj7Q47I0Oh/1IbccI8oR8BMRrkOsYK/uvAL10Gik
6TZq0theSKUiLMj5Va1OHElWCqTnDkuG4wPmpmGa05GXT7U67jeCojMQ4132wOCy
STr8FOlVjXXj3j/unbKGhYhtNtoiv6fQgALwiNqFvtTsD9qLwmxogD6jR5AJ+dMW
DgWblqMsGSy+JUbGtCyjE+71ekDwE5396GSce3Z6vdMoNsa7N44mUamz4x2+Wm/7
UlPzQNtdpUlEt0chsHb49PG309BPjIXqX7EN0dwGPk4kqb/IZk4+fUcekBTtuVvg
KaM9b72RTKYr3X5rci5068kqoAlhhJ5mTX7v7MCbeCtcnvZug713i1iSaLYm3uf3
PAwS2NhyGHGMbJLbI6KQUqMGNg+ETEAupSyYw5xTW4mjPThNII47wxIGd2sO7akz
CTwbd9UyNNx8YioWIOY/U0FSiEpjt+KwmEZUwkugnPZi7UdFJFJ8xS74NL2HKVjr
vyAuX0YUsJ+mqznNyIkmTb6hiek4BPNxVm5Hs04oExJUx7bwH3aUXxjVEcD3gsB+
vgmVWfBd0s5x2C5oyZM5MBQw/JEFO+XmTLaFC0HjC3KDD4gvD1C7HX5mK3i4G3aX
2pvrU9tQRCWgmlSBjrn3E1vTXCpGyQzPq3diRs/mY05vtniP86AAh2MJDfP4oBey
1IoI5A+Xh+vi9wCn7/JVxMUUV4vrOLEf/3OPZ0tcPIjmZz4NBej0mwvDFq7hoxpg
r5OzvvRIW+2owMKvDFKMYg48gQ6Xx2KexB0rzcFgVlGNeyJVK1RIkgLUb4EhfM3b
aUqdWGr0kfkGA0RR56+7I/owlOLeew+zyijCA95PUkURCJ7YinZmri+nKxstDUHQ
sg4k/RJjrwYOicgHruX75AkLiXH18bOxjrhQbMV/L/z/Gbsh3VeFuVyxB95Dp9bs
9E2VEHAp2rZiLEGPxr+hIuJ9CM1GmMGOho+/JEvhXCTXpqezCqTR44HKBqg0X6ol
VmtdILcaED0ef+DmY7C+3HQB6xmyo1X4Yb7ggyjhBKSbSD6JhUJhZor2HhuVDbs0
tmAStldcClTBz9sxvdKTXgeFiGeEJVZAw5K32nqJqsihph0+9cRyKBqC7cX994dR
i4B28rxzxypjKg3UsVokzIOftQheKXG478pbUZdUZx22n/feLk1s7vek0Up9SsnH
TjxdKmdJI4wKPbuu2Nwqkyh0ZtJNVgqUQ/yEuQLTeiAzjoHxNpGNQuoCc6czHDlT
zDgyhM91MdwitHifmpLy2B+LVCxe9RSrB/T/nKqho7OXgmxhNiz8BlXTVHxvG0yT
IE4UoVB+bNsBBva+0Z+h5TDvlfxWDIihcpiV8SMM26p0+TZ6kTvRdf3bqKjR6sq/
TQ5eff5waV33bAL9jd5vd0tnXpZeu6aog5xjDdxwL4/w7itu7L+0u5q1mjH7VwL5
VQK59d/FrnkTzZMiJaI2Vk8+yAqjkwmFUqHPB+ztDoX1b5S+ocMfT1BLYQ1SQAf1
4icSP8mEguBTrwCZUxFeGiCaHsSIKqhXcmAMtTTsa9FxQuu+B2ziX+DjlzHgLTPC
rHtQMQ9xi9n76JfTfscQuxcFtW3R+BRQUmvKekB1/dskIuMKm73VtDTMs55CTw8N
/TNTHDROPaCWOde63SVok8YkJFKPfuSeKQEl2gmpwmSaVO4ej/sKIEdbhn4VTWvh
h1Vw5B+zyu/SM1IyjLOLT/gQVmSyfm0zikfkiIHvGgdUvwKTuP6VSnUBYMN0+CNZ
8pGKxEYtbJk+ZOAqvUn79Kx0/A1Hf0i7mqvICyJYZ3IE/C51N25bWuHF1N5U+nFx
7e26R3NDQ4tUtPeF5DehozvcLgzdejXiFMJEvra4yvvdj8O1bKszOtQuUdeM3gUa
v1vyDKZQ6wtHDLyeBVGfjTN7O6zTk3PP20DpNHJTLc7WDDmqigSB9a5XsWMwWSh4
7PlP59Kb8VxauPoc3tm/yA9T3UtWgGpnsj7ni/BSdl/pCogtjfiZunE3tAHkBO2N
ajP89GjScxs1r7lqACvJrr1wlWq0whS3NNNeNvZXkEHFKoY0zRw2V9XN4EGP91HZ
Rozg6BcXvhTaVYsLEgbQuMbP1cGrWZ5Punuqa1Y66XMritLCBGdE0qrLL26Q+i1a
VeUL9EFUmVZv+tIeMEt3l1dzu3tLRyhrCVmf5FJmeCHuAOOmi/b7P2Y0yvURpHtM
3diiathUFBxGRxNRCmKX9nTyyTJ4xbuFz023IZ/67h4syQXiuRvO30gryJpWrjm5
hnZN4Bg3deOWKdcImJWvCjRFIZlbrFm6mwBUQS/UrekgYeZrHTuMabFwsWu5osQ+
XEiei9xkYM80HIPyRJ1kkpAKjlQ5/HjFWxSeflfvdimdzO+g1votH47c9BuuJh9I
DS2YDb2BOXfrYvTUQx94Poa+4TYqjRlddza+OTkRUAh2FWl+tuJaH6IvPy7L6Uit
d8GZtn3AjrEwkhnhc+dAkAuXC5cZCcrLuFDho55aeVoRDZsHUvgYyr3DnwJ82G5n
wySu2OpUSBXEZKw1AQoCAxbwfbXCUR9R6SJ+uoRz//buY3QhhUcrCSWwaJwtAneM
pCUZMnidpPQN4Vr/uIZYsurmRGbeCu/2h/7a3qZpgsToHC9pU4u52kzVescrBVj7
b5rFpVvfy5DbzjpjUiZE28gaFAd0eMPp8YMghwyFywjPqgXe8Y96NQZuBd1cVl1a
7FB4bdWOr2JcxH4JSU3RCAplSQB0WEwFpepoStOMZvfuJ8S36LAeauJAhe5T7PWj
fUsI1TEcNNiIEqPpnR/B71d2qtX4e0ygzL4AlKMazwVw2OTbb0owL8KS9g20o7Cd
ddSDdof9R9WLQDm9zsWH56yYUygmgX/bd0u8vA9BiKtpSaIJBrM4qMahS+GRVRkC
5SD8kbaAcmqHM8rpuzbEsxL9QLzTc72czXGWDCudslVHEe2KdwZT3Z//bxQHYoej
oc5E7CXp0KXldtkP0K5pTajOHyDvbjCVZwhojZATrxFdDVip9AbLunRtDwE5WNBX
HXiaPTVYVDUWdPwJ4mie87gZItvyS4549AN639kSScQlatdVJ6tUjRpdcaRaXyTg
MuqDG2Q/77gGUni2wvp3UK++UwGDkAsJ5LXYAwTbm+82atmk9+4g/Sva+rKdrVaS
wYteg1+22q4+Klsb6Z3llQoWSSjaN0Am0Pfxu+WQ4aYe7v9qZaPDJ+Hi0HtaOSDv
JfDj6JL1rSdQQI2lqAo3tICOj4Ij1mCEAkOrUeckRejuAOHLB0CBMVQ4sAO5FWF/
DAg0+ABwbHBAIXnGB/v9N2o7Z1eOII1z3H3A3GOCXJ1HZ/jpcYyb4wGyicFtlqsH
IVTd004RuGcxe68UIhgbizkIRVY7P+DzNbOY1yeTwP9FdYDI+XsJo0yjDm9Ip5Xs
iI9UI4jGCxKRXUOIvYAoDIPSZI8I2m85xu0kFuRpnJpUROZGPdbDlfTgQ56oy307
ox/9IqA1ZWwU3542/DUT+aSUFeBt2yl4zIIrT8pwJ0HcTWNqJ55yoxUHhn222Xl9
kSNliX/xNs4VLCJPA6CRjI9hLUF7k3UKvLrLem/wX68z5W1ned8S4qR9RgpAF6p1
xHValUWNtFiZFTsFNVUq8KkamIWW/CIb6VGpsMp+CpQjnASN4/rQo9y1oh+1UQSp
i1GzkS3yNpADSL8dCKjR3Hxd9bBsmU117MzMAWPtHx4+Ara/bl/9PghJ4vq9AGYq
OdixWQSUYsCJ3bYw0iR0zjyHxIF9S0yh8+eeH4gDk9YO5GNTp5nuqMeLMutN5dRJ
AYqnCGe71T+w9ovtTwDF6BpoVc9JgBLfIujXfbYJoQglb4CNKadnFJtSlRwOafnt
vfcFTpDpLIAFIlzXiwCLSR3ItsgthHkthNwOl0Kgkg65BVKGVbbitm2/ncsbusio
YwK2hpTZPqctOqdu5rDZhMnuJ6td+Rr07509PxqXz8WQ2aF0kH+AICpiZALkyv4r
NMjmHqFqF4MmFVpavd8CFOjmtVoKg24Qhe6UOGuh90xcZ7qFio4NqkkcTCUgr4+3
usCa99Qf7oRV2Wm83o6BZa/5ixuTddKh3yRSUZo7wjbfCwwzfbi2sf2MDHwyeJL1
cueRf+EKWQO/9ymYF/1y1HSyAFfPum8i4KlQzg/nNF4lbGMihK1WuqgbKKmlNtbK
bwAGLs5e22biB5UWbwfIsiSL+TLOgHjJ4uATvs1axcvfi8mZskd/yT2ikDmfAzBn
L0eK0tB4zqtG0CNZO2BaP3qoR7s0U2ttwZNzbVfYIpmJFFYtB9oo8ZgPY/re9VxY
8/Xya954jrFXzMITTkaSnOp/q4vK/QoP1XrXHMuSaKSN6TADaqmgyBAxni4HeDs+
dC25GDH+yQwZ0ikD2zz1b1ADm569ime71KgOnyrvG6NN7npR0rjoKWoyC5ESzIMI
hVvfAnBrnT3h2XDBEuCKItB9BlYnKnX+7Ip6U2Zh9YGOeBOjTOZeLB6O4vgl/Qdy
R6lbeVeOXPuATQ85DZezwbkCdMicXD0IknIhn/eEqcJeespfs49fmNLa1EMHG75d
CfN5MyEtt5dl5wlBR74SlnTRbDXnzpQyTw9tFgksrJFQXuNFfISvLkGdMm26PS/f
2CWqQ55DBDJMML35gFqjGWSu+Cz5zieKxn+8MssyhKchTExxxlwg8h1wtGTSeYwP
cCBoy5R6+N3ACOmdvI/BfNNxTj0J9bhw/fR1eR/ZHsxY7IlWgEIw8QDrvfxrea8e
IfSWNPfIq5qfpBLDmlct/hUU4N318BXqacKwhRBC5lptpv9ENO4haMSlGrUiDnw9
yNHqD7HIrXcR8tuGW1w5BDwQ82TmIMVMVqK7i6yxIF9I+mPEjTQX6iay7eMZ+B5k
dDUTHd9xH6xhwWbLEUquzl0G3wp8/D0I0PYOlAVqinmSaitjmHarlACGhOyweny8
JKcUowAreFrJFo4DWbgu+tRvpLurkNjxETTExvYiKS6LE7ciK6j4RG0g92PuA7Qn
tdN+gQlmx7H8Emeh8cla85xgxKbNGbnQ+P0MCLPw+q79698A3GQyxTGX7+eVvnZQ
RszGwwzbvqYI8F27IVryNvH+hYkbVRTIzm24ONapfNqnpl76Y9Kb8iqfjXA/KUPD
Q4QqnmyAE3f8HJBXfeJaGDEbOkeScSRB38Zd9/12NOdBBPYH/NcsxiNIC5mqIafp
cAGkwdZbxAD9V0I/n2VM7IrruQKziAc8YSJbVZoigOQcmlpq98sbNJU7ElNgnZiI
AVsN0Et/nDTS/7UmTu2fm/JjJBQTmS/12WUaept5/jl5tXjQ94EgFehDfkond/oS
ymOb3OuKXgsXoY9OI80AEZIJ7MKbIsfr5exYoLFmFcfpIhOyPlfiZJNpbKZgtw3D
GsCqecuaEZRV09W5Ee/ExRQjUvB6SF6s2pAbri/hKBegWkZMV6EfTEpNxtPQkOTK
PDK05RWJzNK6AhAE59waPgPLVLHtoaWxXs/MdPuZep1yjQHheUFHMhpIl2ThMevF
MyNcS5Az4bJDXErJ5f/lo7oiLakLapu8CfmmlqL2BJZKBq3SQGQFA5PTjEU1nApA
83+KAy4BXSMC7J6SK/Ds16/PIIHjfsmuV/cUbAhKIHK9ppeJNzNN8SMEoBLqxI3j
gXRtcQaMOALPcqTZjx+HffmqIMRWy3P3n5xNjcsX/DbhFOjjgiZwdc0yEDVIHvMU
h6Az6OVCXq3h3/rCYbG5SooN3STLqLbMoZ8uGzX7eAbeOhMerv/cVYr5AxIKnCYj
v7I8w4MnP8tVUt78McC01da2MldZtwqp6XCvPXeZe4e6Y0LanOUfeHTcQX5jQNLV
/X+4SS99oqQDmeeYaou7MkIyR0AC6dLKBIYEVByOKqSlCunDXxsZewUB4u1pApx1
ZaHHHveI5AqFNdkIMYlEWh0AZ7n6kkFMnOOx26hyh+wu6th3yZWEM5nRVPAt0ZOO
KxxYIDIDmUChteJUwjwmEnj0MkAlWqnUvcTrgotHRDS998X1o2iHxZ01SjWAaZlg
K/9eKDCTozhSYoehkR4agO2g5y1ps1QBwJv7DUQk8dzNdePf4PMHt9VA/AtX59JH
yDHgfgusUXSs+5hctSvuOpDlHw+o9SEthmXxGyUAXQPPHALSuXzl7vgEnrqZskH3
CAc5voy4RFu5/aROSgD9Q85TIrsPmBbaot4av6GL2o5THmvjrAXJoxh+b8ENv+eK
Y5DbQQTLOkiQkgES+IzuNFdgrUZJLRTGo3zsnYc3gIrC5yhCoEcFNeN4n/qocGR1
J+2+KdaOuLeTJhNFSgc4bFq8+vPA86Xr4gLHuhCgOb0GmmCdsnshhlKRkzs4yhxO
MbhOHiVHqJVmPY2MjsCExQuOvWPpKx7vrnJi7lNaGVf6OScr3DNbDkXKVMRcLxhO
8qJW9IgA+xQJ7Z4XraqFyB7VTCcaDPIB6aCUq6CuMnJIxPFrnMzuT9IHHl1nxs/1
bmfvhBKyK9pAb6+4PO8HMLO54TfSNTJQQTZ/aUUVACdG/RKQMtAe+48gM3PkIHYJ
YnbT3ufxaHLz/eSeqnZX8WkovudiU7j9az9CbSJTsW22VrD8fds0P7qhjRliXZh0
d1n65evtCC4ewqRv45Y/eml4tCoZaIW4zG17UFMALHWVjS+AXqQm/Djse/nHPsXG
F5kBgtx/2sG550B9UASerK9Rte/oHfdvV75yY8M3piU1SMlDq6OE9hUHIg3BB/Su
sueIivPvz8dgBqcKs1KxTsfnx3hXy0q93fJQv/15njjmx1zLn0j4CiysuS8MlTj+
X27zYyrdwvRTlYSShBa35Bz7Rvvjnvx+dgatlptPLvIfvST5vbEgw4xOlg5B8I1H
8y2R6w9zFLxbK+oT0j4UjEc37+0ksDMBY0Nm+whORlcGP6qYhyXZEgJC0KtWwJI+
G2Vx0Y42SWnOod6pFFzErZIq+gMmpuZjE0aAVql5ncN5weK7R2HO75nK4ZTGMTxB
OedqhJ/NEQZaRB4znJWRl+mw2RuJWX0Q3KhB5Cq60pWj8AFs8m0cF0sAkdFiU7H5
0auhnpw6TYmTDFJ52UTf/6DoAttheIV/tCa96rXmtYX3IlaXSlA7WJUGEcQVSYH5
R+Yp5JiHT3TtZS1psGsmhn5Gv3LzsPOevZVBIfxAWYXHCS3O2AaYzt2ocm9kmngy
VxG5t83/xJSgRIy3tCU6L24XEH/dwLk2/UEIwO2VhQuXN79Hld1QSjPBhhqrE4w2
j4Oj2SwPZ9t+XP4E0RNF5KMkrA64muYcQU4Aw8BvEuQmZR8dOxKaj4+wT3hRa3hc
+pDZF5GkTpkjCnyfJR6EpmAwMPNM15L393h5lHg0cYSLtEIrlylrYzZld3uDX3bm
cfozjv4Nk43l4UEISi6xichQs9HTUE1hoDDIVW8ERDYfXxHcnkJd9di7fvcqVmsw
avr0NK9qYL3vQY0DwB2jefbOFyEtdAElC0asmC2lYXx8cQAHsSjde7To1BF1RuGW
Suitzi0sz/+PN1bcCQJegH5Lwy6ap29TWk8Plg53FtRrTPLquCJLzksadmBhTU7g
gbHK8kFsokghNHN//y2Yw0rYkXZbhu/s0mWUG19v/Jig4SOV1YdqCJScW8sWDVw8
AhogKY8+ApoyqYTUa4bxw9qm0K90e9JkRzVZ5QlH2ywtTMO+eTazlosu31zpV1uD
Tw9LzShgnwqUD/FfDJxq2zILm/R2B34gatESrBmCQgIrFoPhElb0gMJ0k+LE+zaj
7ZBNVis/yU9/arsdBA9f7qREbgoD8AXQCOGP9ZowDRKR0IJQz57/T3g9LCUtyqi2
TSp+GDCtWXs6dbOznvUIC7VDYgngMp/xFumoi6w7lzZ5acBJ1Fey/SeJqBqXVmzW
LvEuv0whwjdow+vAYO3hkvtV40pRVHk2OiatW695SvbgzrP2bJvbJJ0vCUqEYvNZ
z7AASJwKslQsJ41oCvJsK8AUBPAJW+8TfnRkFIUQz4RtGj9aWjsbyMiibo8XcFut
8ivQu3/fxGSIugdfeg3/7w7N9bYGCX0jCcd4tm/7lHQSQW4dQ35EdWHsVamYVffi
3dZ2Du5eL0eJf7exi9QJTlg46hPJHVh18ALNz8tArU/4VM0i6p91VI421VhAjd/0
KNaEHgl8wKlvFYuiUg+qFG3r5Ntb1FoogPSzrEqLE8u3fX/DUyf4pStvLRlgHHWf
QMIAmmKQerpU+OUsIPLdHKWtFeTsE0vqxs9EhWsdRln5LDytReI4/GknAH7r3gpp
stTnwt4foAcuhurQtZ+jhok7UkLyBHHV7Ys3Wd2sk/vBW9m6z/4WqRFfRZ61k4gX
mS6u0BnWjj4ijYXruVjQj0S9Zk3hXxr9Gytg+CTOhPVbYZ5UmX0XTmZltYLA7B/t
F61q5n/9EVzxjxqUSxhcZkxFj3nU4VLCLJOqK31jh9s7xzPFa9iiMLGc2T7KwK4l
ZO2xVPLF56Zi5ldWEhQAsIybXXquAnBpT9V7tTncjcFQltS7hNEw1XMzEdwkL7/k
ylY3FgqCPtFOBFl6uk0C8gACtfuFi8Cdjp16mHbrFTAWEDSOT/si+M0Agt1ehjSZ
cbW0aWPyCnTNHkGlNyTkTzsdD4+hFE/mwwrIGMOChDrZ6LEuavurxfibnWtpqhfz
BUv5Gu2t6GRRE++Uzbbi44wIl4xUKPKhNHhiIrK3oGOqa1da9RH7aUtJo4kd457g
dTzJ+o8EdbJAR1rxc5QNqHUkoSJil2fN+TMt0JYQBOP3QUK/MGc+LVI1dly01ZVr
WcBXOobY4OCauGF+9FOv/YrxXs/7VhhNoHIZ4S2qeWSya7OeDoKEcL4ge8LxO8Nb
CNfR0FnAIgiQqmL8rvsi81ueCXu9ya+tXvm2uo1wxvzQaSkAgFPkWnbaqDtzvesq
AlCPQEhUWBMX7NLW4Sf2xdurKOrKEBCOfVbNl2HcBKxTVRs9iyiuf/OaxIu5KWv5
kebfYIcE1dX67BTsb18sN56gpwzig3D6jLvxckklhN4rjuzmtWa+preDjoCViNo6
UNPxAk1zN20ZwEAiyyKMasJKuHb2/MtoaEdYBjfa5p/hj/BAPaf5fUZECJHMgAah
QvJJ36i827wA/rdaINFyN+C9HEUriFRW7ylAltV0O8+jBWjGUhfOXLh6+eUHFMFm
6SpmAibvvedvubtpyI8XTFby+EWcOg4INoy+TSxbkAA6mIShjKSOxBaBAQvW+Gdi
MU4StRcgdBMyjL7Kj36FvNacjU9qrzXr1y9Ua7T4eI0LjzRWrYWrZL56MMkrHro5
qb6G9fSMm9V8al1LPJpFpgOPrHeq6CCTsJ2W8G1zZ62frlJ8sdh6rAeAuEVKUCrJ
fHN3XIyP7dit9oPDOlibS2xwyuYB63VfTHPKcwncN2TxFKTIu0LQiqd2EMOPQ9FU
DpJ+Zbdmptpwev2c9QsEDJg2Vak3uWzt6C0Lu3kf83tcsImnsmnprWfvrkfhGtqH
7/28qsMbAt7I7y1JCcrN4HQdL2IyI4nNAG3hW31snjLGKMq1KukmAL0yT+p2ZzYh
nAo0Zvuy4B0Fk+pt/1LhsgWY4BTlqGyJohoRdz0F6ceje9gLIPF3EVSagYCToQrg
aiNeTvPYpiRJLLFvw8KRnZTNXycgDuxcxSNuJRmOaDgnsefy3N+RkAViFyNQnuCY
aoQSeg/pLHJR1im3Nr+wFTU/L2ocEDdH4YKB5WQ5AtRXWpiK89+gRbPPI70J8R4G
fRFoVFtOBt0W7JxpXFYaCfmWU9CWnx+B/IUm6e22jO7thJeLFuKiaZ+lCmj2//h/
WpjLGipmyUj6Emh1cD0ngmdW/pv2WbikscTeEAbKvMbiN7D9+Fj9Ve9JEwc7/sr+
XjtbwQpAjvgUzoQMlzDsbiklQ8xw9BDjQahOHxQtM2ybbCJzuexohVnNhJn4p+77
0sSXuKsD0n+13lvK6nU0pinZeOdGTvSZC1udFaYkzDWsrw68SAff5lCIKntKpskA
qCBSrGLZaiDaCoUMpnNoO/fbTwTNkRu3AOwo6Z25BhI8NfST6iviB6J4qVvQKku6
y+GDCQi2XuhJGOnC8WwTGfxx1Amd01y1GIRQytIV1KscE3GiuA5hc6/qOsdgOVYB
v6e3PyDjBB1ButaKqTp33L9gRnfLam9fdrCNLepo2UuAcavnODjzAo4nOfjeEVzk
ZGCmdBdn0qCigUR/oHxAluaDPZ9RrvxwX8AWXOtFhW0O847l+fNi5Y+v9C+Bf30B
ll7nA/jqaIlBKvH5zirY/iWvUOKZefvmC2if6HHmWHOb1QFQWJieLU+4dRZmg0lg
LxSlj++76PfqqlXQaMbmBxkFwMErI83oX2pq+r5VswMxKSLIpbg88L+ZLHjavrez
tf/mbfW347r2cL6SF2KewWhSsOc/bbdsn+bGTUZSY+I1XQ0fsCKI6x/TtiT4wUr5
/2mf2P2eGh+XOoMVDDrn7Kb0fwPaZlJdsujq6hABgKl8ATgpFykI5RL3Au6w+FcK
JD4XNY57CxqiQw25ieZWDs+anBNhq8vv82JQSRpxd2lM18vAk6Beaf1I1FA8de2r
8xj5FfL1WgdWHKZOXdpgBsYsaxUSuzgfSdzZsvufnoPdGI5Cttm/japgOqWasFpw
5XhjdsuDD56g7Ag9l+OSUyfYkhRbJ4UeS1XYqN7lN9Lf8qYL0N3M9IY69vyJQel/
BR5wekQHUyAOJvHvqd/d0UCMhMCIpFokDf44+H27kp79QAyCZfZGHocTCOWgEvCE
qnUvQSAidiQ2qCKDILXzZN3Y5SNMncaAOVq2+io8OtXZRHlgq8llySaFOC5SZPfm
/aFxI6eJw+ZfJxKIa4cTBQk/0L8hSAY+Jjq4gFlyXTUCxW7LImkGSzJrpKctQZ8W
GutlftvEpLvNIpHPjiQSjhNJ6fo7mWLEDUUe4V1AEiNmjxAIobf2T+TomITdolHO
RtgomOunKomKtBebFGatySKUSLFjSSJ//Rod+26075rkMd2xGmjrGLN01lnRd8gP
CPi2sHEL/P3cei1Sx4L8Z4kgXysvLbRZhhC1cX8nD1Zv/7Z9SQK5VfTG+2srTWwj
ZXlqQ0V/8TTHlX28w0RoTdde4D5dkHeSn8D5gZwaZK1V5pJY/2svz44RxCD02WKf
RhKyjgTEaml3lBVMQdBrsKyG6If6sHGeWqn7El4173iXQpLRuhPI12jGIlNOLyZx
3cPolnbVxMwX5Sa5gpEWHeU2/DZF6CfLL7JAVKDGHbhGxPVoLTQIsEvsnlhLU1k+
/eiaG9QzYOoty4/EarBfZr2RqMzQV7q4R9I97lsuwyMUSeOFLt6ckknbbb4p59Fp
9inX/zhww2x75jc5yFAGItjHOPpmdm2r1GD0M3wSwXhbGRKAMck1bsdTkkdrZ/gv
n0q/h7QRaWSaCA7Q/FhEY6j38f6M90o8WoXCCWb44t5I5+jbIRfvT/u2YH+yp+FB
/tGmbxeghDABr7kTOBg1kqk9uQBt1nt9bo1fxh/ed86SU0Qk7/Ev1khXxldXoiRb
QGtRX24DEr6d8PyVevGgoTWJHjx8K0ixVrZISQIKvQQbjiYOpv7hYuyqB2kA3RNS
QmLlEUv+NOb9d72FeO4V0R6Ih5S7RkMJ+9CM2qBfHhc9Qn4f+xvcAjjk9ZB3JQtW
ogvzf4zLUdczPwyF2M8n7QsSJ4s3A/Aj0zMflMClwy6zVIj7e+cvt+pDMyCo8Fmz
8PMcZ/MceBdT7fpvb4tT+La943D7LA9ne5d5cl9OwfAdbn364GNIqSRutCmehba/
yZMKTaDf4Og7F69DgDKmntbL28kj8pa2fbpCyxSnihOu0C0NU+VvNcqbxWQt8gXB
uj+/rAsIUjHr61SZuyuKITVdCEnvwRjHA+1kEvGYfzFn8dBd65o26FOQOrUYsiIL
YCqhH2+PSzQGJxQ3hW/iU997m8baG2kdYmYl26rfSGgmQTr/p64zpdukKAaeA2yS
7jSr56GUDhGP8Hoc31cgAUCmLtODkEgRvB/U6818a9Hcn0Mron0J1JXYcg+KbsHC
x+zN6aX1lPKSTjZhsucq1Y3y+m/9/9FFl2Ht/eYg1KcNagNmNVQERAay2o6SZeUI
P2vyF4RPZmewk4B/RhTa19uQIZjNllQi5FCR1KZ8WwQxMpiDTXtvQ+8y3e4aSPMp
OLWDa7eLfxJ4D0AKe6XD4vvTCBHEd++Txg1/Z6AKM4EX1TTUdC9yT2MZuLgzdTlM
5Aju2T/lbjJg6btwGDSpsZifg7o2/wUpOaqrGH9MsvdZvMPTa0EisVMWHJWf21HP
kZcyDdH42J+usGYZzs4DQWQIjF0eblwNR8bWNykDL7FIS06SetMT2rsWuVR4jJJL
r0vLt6W9LfigMnXbEPU031d6WSnD8Z0A791bD5XSR+woVVS7qmDDZFGtFg5BbbFm
8JEC9VkvDDyGlQWMAAVjb7Rzp/wJpMMIrhev2HgtnNYVCDftao22fPjUe5IddX6z
NIM5NGmSOwnAaDvSH2uGnGkR3mJG1xgdKl2dkZoeAyHyLJSWeucWTd47G0A0I+FQ
kdbFbRERRutAlp+JZfTQjHvMl9AKVjKhyx534itUt5i2ukEH6Z6s/8EtJDCo+1p9
Nlen1BtZosfpjbG0UHphowg1969I9fDy0WNNzaaqJbqBGoVs0PbOO9PL12UetRmm
ABkypMKNZUpB3gC3YpsCHWFQGvpeTaU3AM+7bWvQ3s7BqNDzbdYfoS8eVlU2RBnj
Skdzzm2IgYkBiNO6fCF4dt+uri+xEm5YG1A5j1TFihC3FtO5v3kYWaxyJ1CvBMd6
u4TqbKdYoDXdB2MJ/WPVN1U/6vKDdKifzSRomswdUHTcqizQmcVDkhKHSoDOWhjE
tP0ibx0gQzFFoody1ADFx6SYUjHQGLKC9fSAhYVEGPDo1tdPD5JX5acHo+mIR+TW
j5kJfXgjsUKK/QNUUIFLiLdPJRg15GF/0C6AH+tjOr8aZSZRROx1mr5PckRQbsgF
DLIFaglwB3cA6LCzWn9ma8Nt0hoaFVtxRAPvoxPRppIt/ewE03oxUfvFEcj/5i6D
ED3JnubFr2lRq9cp8trBOu/3EPFjeVabznQL/6giZpK3q+Fpewar8rt3GXlTvg8B
AvwheixlVSjS6hJPd4f3OTMCAR8qtYb2oZtu9niWfbSV82aqDytvoi7KaGhIavBX
Zl6X8lCmFxEMfoa+Z7dnZz4oJNvYhEt3IR9/zt6Jtz6uamxNOkXD4P3QsoF2ZxHa
zPCRF/xikjFDXR2S1/wYI5QpqMtDgaRqAyiHuPJbqcTFFuaSrnvp4aOVph+s1xeq
2AoHYoZuNCAgYscj991ryvZWfVsC2s6M4CtIVuDeBA3eIDU+/7KRBlYRDq7iMCkr
a+fBnuGqsvRP46G4qth1HHA5Xk5i7z9C4UyKBbCFf0YATPW7FiLNng5Tb80/jzNQ
IWkIsoIgCZzt0gGSyL0+S7AI2n6mP2GGoRRMga660z3tWyI+hA3GARt2VlMYKQvY
geuNUfEjod8mG2Md7nyUyJHVGhczdqOiSSSrsBdwdMgliTQQ3PsjGoDyQpCb2c9b
aN2x4pvvhYe1PPciJ6KcrMAoQ7aSRLr9pGtFZMq74v793W0kLMlovSJDFr4twox8
gQypwlNJ8XBrFHr2LVHTYOujfPOtBOgP7drQsF0J3xGEtQLao2aKjqBaMp5ht7EU
2rd7gkJezK7wdWdBzGHPiGZ3Da7aN2bbfm3XRWdZNGkcP3RglSDCuuG+TbiJAD+Y
/zi8gOgAr7hQn3ORHed9BW0syyIKSVV2a+EOreBd+Yri7UW/eeN+SPadUoZ1rl2M
vQ2LATfCgBUP8aTZSkYN4nhO2dzNr58wFmpDeebBWq46hcc2S3OisykhUncowfyH
csP+wGxAR+PjGDHJWmO+7BRK3AJqykkJ25gmIB07VjoU/iXI601t7dqe3DeTBes9
OjyiTaM0pWdWK+lqL2aLXs7scYTyv/8cTBR6+2pZDA9qHw8lCcglkqu/Zj2ZAeao
kU+KRjtjXTnCWjd8OV+NLSlGxXYgW1BMmEHxylxSpOCJkE6/MYaxf+f/MB/XXJJJ
QIWCrbXHplh2hA7uX6oVOoIEj175zM02CZLURc9sA4qEKXhRG0BoFv7sRDgB9JCE
JScqMQzi8ldKIYnWbjGrXUIXHbfF/YZFUp0whztBR1PQDHtWVbULp1z9HIabFfAM
5IneVRdEu3pFswiJYdaKKlkBAXnxgtqifprmANMQFZ1X5CEII/omWZneiS6h0GLz
EAENItm/Tm6OGlzzpjz5+E8e2ibVVcshHptCc9MXvg2QzXJvTSufsA2EFTAoqC7j
ltStI3TzJJSHOd5yyHDdALyT2LSh+i+i5mXptyb2j/uA5XN9P3QZFTGAsodl0YmI
rSefuZYGr91zl6idyx1zPwMp49lizE0BNcS83Cs9Uxxn8bVDWox7KeJGsY1lL+dQ
R7b2OJD4xmQdXpGRh8PZn2Yd3T5EoacX+pe0pbuERlU1NGO2WY55iViXQSFgrDg6
Pt1E+4A32LUF0cslpPz5wSHvSnD6YliMM6c1fS8xSwhpCFpVvMC4t0W97V9atW9j
qQqOb3CileNIj7JCEih/Tf/zZQvUdEycDSGXJvfPineTURv9MoshcU55ykyPShHT
2QbC+VwR6520kZGA+W6NzKOOIYnInCQSrDuP4Tmo4sbkzvAQclbxMzHVBnhCMsez
QO2Kf58B/WicLeWNDD3gij93w05IlRyEen//SfQ65xE1nlNlkSO7Z/D0Gn4Sfhuk
dmSqPzo62C1wNaVrU/fsbz7NRoqqQJf1JdU8J0OYMr5Qb4XcWAtQPbG7tJQdXbVn
yh+PeHXzS6ZF3busjTe9j8i/KJDbzahsA0TjUgU7IFZigVoBaMwflWw4mU0OQHjV
IpxQYEdzMeZYDyy8HLZFUV2sCxPLazcnAAJrAzIh7LEQvmV2l9GsUvctHTppFC3S
XhRAL8eld9e+93PgYATECCJaSGB+ODXq8A0upV2lsyP0g+fw2ghnyJbLozgUJMes
oNfsbf6R8NwxoKfZ+DnaJz2Vbx2EPxHxSXdGFbY0WNPS0AZ8sI1yWcBSgJgnKEH5
d7TZF93YUbUriywSyLkVmyTz/W7YLbIYJcA3UBspCHQ71wM3XOjpPh0+05c+BS5f
hJHypoS1HqajtpXHW6Rf7QkrRnZvgyn/+Agh9VEvo5Fg7D+OkDChAuKbIfZAxgWI
9X/puxn0Fil7GhGKX2aLvcAmM6stUl8sQZM7Fifv7xM2kJYm3yJ9XaT/NDV7qCAF
jsKZPDkp6HzeI6GKd1V3TT1MhJc9GjMN0D3ZhZmVE4xmm1LABrmh9302H7iWPfVD
/Wm0Hp7uHgwjZ1DpC+YmlZVppbdg6/nhIJEVJSFPuUWu6/EqDbOsJxUcgfhLDpoA
hdQ0tZIF0A4UhmWkU9zVVpQdKkg2bSzq6F+518lpH9nOu+hYmBOfs4Q/VgXuRNcM
E0g50yhfdOxxyIXdB8/FGiwbdWBhpFxL0zaUMwa4S9rts0cfzhWiIgKsaFGpLD4/
8EBOzJMVH7FFf6bzQQbcGXWvv4ZUfzhjormV8sfuI5jVt6PVyCR0w1X/3sJgbGBt
7INy1jlZ/Ofs6AtS7RA7tMAepsvmNUXN8pUWe2rAFNgq6vRtDGGBhCCGl/75TgD0
urecFATs9X36y7Ii0faHpClSLoMoJ4zB4a6y/vB/zoNPHVIbW0QtYjvPa+E+nd8q
hlJ/xVRvK1nngRNZNX82CU2MRuugbecXUJLP5fC2TkXcomVcf7wVYumfiL6ZBJAV
lGWBJfpb0g4Q3BF9UnMITwv0Pzw9ghGkn7alOmaCkI9onHy/qX8OoanedVbWK+JG
izjY8jassSsQsUJTeUbuhv/IUgxQP0Brj+Up78oMz6JO1dyOyKMg2Gz6RVeCX9wK
HvWZoy/3ZqYzShbU+2rJOpQXICBgExp8DSjBSCRk0zjffGnt0RZ06Ep87iR4Epc1
oG/CNZKF2v5g/rxcvjTk4NLdsgIQ+V5nS7NnZ+rKLDQiHG2khUfYLjhr5ftF2bUu
cGPAGBScYq9R2bc3HJtpxwmCQ6Gka6adDsOy/+J6EfXUfYKO2JB5J6yuSYAagSew
DNq26Yx0ofkbt4mn9dRPzNcURPUUxfMS6GXkYR5khpH5y/tgYtN17ExUlEWu1N/I
1jXeYyQpNxFl7pXsM248vsQGIjMh6AI28cLiIqJA+sNZLBnpWAK8iWb6nOmLtzzu
mI06OmKD6JR43j8UinW2hA0kyzXlGYMldRKOeM4glM7cdTPAdF1aISC9Ggu00RD4
58i1gtt7CV33eD/6b5+85xprokFZ1+rF8BPZD9E1gaQTZ/a+RU6fgIr2VRLniPsH
19zK9GbA8kx429qMpXMczIEEcT0SvhY+EpxFnZan5C07cU+7Z+gawpBW9gNLCVU1
57QV0i/phlf0DGlUb2dxP1bMt92hcMCeYHE9pBDwePL5LU5Mxz0+aNxXkYJnVkf1
rsziYXLTanoSr8OnU1kn+z0U8qIpAE8KhZMFBC7kHacwUxvXjPFYc2mRW2J+KL4S
Sx71HgoQGhxJL8fT04Bg414HZSDlw2Ojy0W0+TRTZzS7QY4XHqjUlwnxcYokUHqG
+3fiJWgDgIhATkf3E507KNhTrPGgHGIJyGnu9DR4oIvvYE7GhgU6zwpmSZjLktLd
b0pFayMwVelkXGw/xNycAAI/M2uQAIOYGtoG+BQ9N3yFfwMemKjTOWCg9zcdLOPy
bMayj/mrldJc8ojsTi6BK5dnhT7MJkyRAdWubuX55DINgWfJkYhKYECDRNfiDQ1k
vDn+uuLXAVDF5V6KKVEaNcznbiZaktUFvCoxAD0iDr4Lo7V/h9XM8LXkH8aYURUR
RS4uYEhTxWuhU2zUfvrNhKQdshpJ4skAPQUWFdaM+jjMHOelLwLiDyqOTQelw0ro
e+1/ppRYFh1qlW4A9dCqLuGfisOVkBfPxoOGg/5ReiSRag2xOxy+5GxYt2s3ZCTe
IwDaPg2LLJJs2wCsTDvsXyiQSAdH6XAcErUiMpc9pZg5pDlSCCSRWOMky570/U/5
H1BP+pv2NYy6SHNrKqzIwPL+8Rg/Vd7gea7xAsYrDO0pCeAwKYivnzXAWR+ON1Tg
MbyPAB1VXuVw92SjnIb1mEZDzmYtkjPwriyifWMv1QzurSpkET5SVJPYHuFPd9AH
ohXtDepc7INlTzOdsjZFrfUfxIozK9EJhryLIjNXzyQIJQ5/niMjfA2dwRkOckhC
+dkfb76zXjq6SNGokdCn2TuS6snJfAur4FWc/jaV4yxh2KDvZWsy6SL1ahDTeHuf
PXXr82eVOA02C/+EZeN7zgy52MbN0EvnIDl5X9SNDxa0CiYCYI/H5q/ZPmDps4Ca
/jgBw3a2ozoPjQvd9mWuRZynPwMiGSU7/VIPNKtDOptPzE65SdbQzTtEDKV8+F6T
TwWHTrYKqTsZCOVyCaQfoplhNGU8yZFSmi8XkM8ecQJJxwZOTorqxXlQVdl3MAQS
UesWeRf1lq1rWxat6/Ymr7gjB5yfzT6RBYLI/zksft9HVsIecK8ONOsyy57mkf5Z
4prj8uJ/yf+evS+kCxd6jMsX7dpY+T8+bkXfcy+uXCyUYecFIlmB4uVEAMCvpA2x
zWOsq7Dwk03s37ARWd6+G/WlykvKNsl+QV8JvcLmKqQhgeNnTTO7e9WMVzjfyj7W
jsUz8hYvCAQtJnNvyagD653pXeh+JSbeluSxIP0vLrfFCrx9mU3x1hnpxT3HahSp
aufMc7zSNtZAcfgvRtesQ54LihhWmpM/a5zoD2ke40pVgjiSLh/ZXcJR6CtU1Yoh
PfptYWrQ3Ft6gXLQmMRQon5skHEQlgawfNQ5XHojj+JZ8N7RBY+lde6FY59bYeW2
nXuACHzos/ifbpkGhaV8h9hb0nMDSThgobHuUid7DVKE9vA6qeVoe+kVlzeAB8us
5aBucnRoSVmeVYvEyb4IS6xN/PTJ4WQqh/29vH7Vu0P2/C/8eojDu8UWVPxWIhuy
ubCncn8A1wYiQ+Yt7xpVesMA8eDaroYLX1+BAyuqVZ4fJ4MkW/6l4U5hidHCxR51
QVXmhR9zPsBv8KQQHP1xBBsowE5WfFXXPmDctBTcc9LCFeFhFK3+KE22iViPbhS3
vnFTGfo/x3WUj2ueokIokZMvLoWZ3iIfE76uNJJ4FeytpIV8P40Z1mhQGlye4Tzn
ZItC3r3AeHflnra0MFkZiRIv3hObXaTZumFlOI6/xcUUq1NwZVZX0MoibPl6pY7C
h3CTm+Q7HwI6FiJcPhou6kC6xRhPJrKVxCX65bgIlboQZ+qtdhB62q9xzxFZt4nH
xOwoFDljiYXJQX7emJ69xIYXhBbXZACqRomLymgAXDIrv8hBUl0uN81WhaO32OXw
7vbswBdkUwUHWs25CJwmjMudyt314nTg+gncOSStt0WbE/QEz6Kx1KbzWQvmlw4K
kZOMEJaVt7X/RtlQ6k8H7LNchkLl/FIQfBmW49egOSPTp+gqpNQVeEmTO2y+WILg
rMY/LGJ92yY8gCDI2Z7YTq+iLTiNSi6+NngerFLrHH8WxFpDnOG9ES3tIqJt3T2g
RPeeIYPdj0jCxMe/4ikcubhFDEcd9BH7EJeHprfl8/8kRl6yJNKSuOAnZgYFqNX9
f5ciTSI7DKI2TXEDkPzrMOuG3xhxSVy0zYHd1FTfP/wgITMniqTXWKwojE8pjSmh
3VVEq7zUdQVjuS26DYWWMzvzHaJU9BJuTAcSYFB91+uGMERUW/Rm0UDjATuu9a9b
W+H3m1lpB0NRnuEoWn+sXY4/Iz2AIjWqRaY6Usqqmy3yUbjwLekvjkmStfjCoOLI
wR24MUAHPTI36z8wJQgzBEyOTza2fWefsiKcSlhZVcrvu7SF7RY5zDqvmE+9lX1t
vx1JYvYdwaKjfptfhmBQnCz0cV/2uROtnlzfZbmsmuYx97FlLvdpHB6CTxDDNHEw
V0/RazB1E/ct1GQG30vk0SAN8628DAbdhSgsBKDnFvlBeo+bCkd2NHGkkvYbRx4z
Fg9EsglRdLfXNJsV+Dln0Q1QXiBLp798HZaiksySm2aLFlmvIbmx2zhoGbF3ChaL
HKc++9zfjWD1deGXkwsk9tPPazg+iPJKhkYFvj+fJazYTlixO+78Apu5hw0L3HIW
XL+OZZw4cdom0MNkiHexscael2Phl5pjTB7Zb4mSbP2SKRP5vRGvm0RSn7NgSwZt
Pilwlk/Fd2QDWrAN9u1QoE4QnG8pPaLdljU/gOTJDcXn9cs/bY5ITM3SlWzWMcDg
qxS88w2L1WQYpJANujVJ/10OoLKoVk9XG75nJminz69x378DVH8oWgnA9/GVkmg7
gXTwiCkrBIlZdIu1br6xOliNljOzcYE1TpNrudGSbexvdYYXjNa5kSSvvGgpXCWO
Y/G56HJG39ea3bokYub2jzekIxceTMMW2qUzlxVe+BuTwTA5DVA1hK0QiISzUHMp
f96czx7dXZP9ETJTU7pCUBsIuCV2J79pS8GE+b+dna/PD7PtjiCnQ0SpSPACs5EC
5dOXH4orJEjxDSjRkTQ0BQDpfvlqKoyhOGJU2wz8KLteoCR/VJZBjPUIGHfI7bOD
TqolO6ctQy/TTklognEPhprvm2u9TEHc9x1PMpLrGfaMs1LxqcN5Ztq6a/POsyfX
PFtWtKidd3r8MbNTKmmbM4zPBBeeLb8qZ2E7SYI1W8OmciN9wbZT0AB2jLSln0gF
DYL46xlhvFK59EAvtP4G6v2z5wQ5N/tijdkL0aUSdq0QFsP4DrmYqkd5rMeqgEaS
7kv2Y1NG4XI03KKp/7n00J3I3wP9UqikPn9CGUN47LUdNqXf+8ycuNLCv/JHbBc+
UfsQpkgFXzx9hoZKQUdb47/ylTnW8YrXBZ2xKX2RSiD+LD90S40eIj7FJySKYnFh
wKkLMrCgMCwA8tLMAfP5xB4OB4EZ63bOR4xo2fP/DN5ujg8jiIpHv0OLgUoI/lrj
6oyYb5CHxYYqpr4gzCVxd4pAOCKK5gSad+kSfTNbO4b6URbJ7OO2pYCRj+BvME3S
0SXAiSRlk9+Ab+vydphg2gJVv8WoHocC3/xNu1MMkQEMg6vQAi1MKI0Tdfd7EzFb
Nvb3aID8+bFVYoUGDxFN1RR2Uf56WXigmKBK/iGN6UrIIPgepuOZaHfy8UL6Uc3X
fl98l0vZ7wPbBF905lqo+gYEWPCF0ePTHlOXoD6y7VBhEvi8ZfFhhSEnRDaFys5H
EY6T2hUBRldrqyr3Za8svkgP77JtrHOvVBt759otxMiT7e4R1Uy0ToiDNlfuF8m2
ITXX2YvMN73xW9tVBqnMef8Wm8kxkF30sqsWM18HfHNeK07S/UyqYrRvOPUXm0ty
I9yWkFFwSgwRdTf8vqw0jrmBz8oA8QY6iJTwyqQ0IOIyM/Q03zHXjW41vfxyCJ0d
feIRGdZdtHRXxC4jPpOhg2cQfjHysfMjih1vcvGsu+w0tzENeoU1Sv0SaLqXbewz
wfWx/lVetK2j8v9POFcGou19p3LDb7V+4uL6N8YYa+jOZFZrKZ7mIk76QPPsBIWw
OB9D9F9ch9cq0YB8FKuxSgaOuQFblIu8Qa7xs96j3auzLehCHpWBkUyXCiitBRQV
12hecXW0jM6UaJueYBwORUlwJRbgQXL/nPXGDi1ivWzDjBRc8X24tzU6F6vFZqwm
FDNvV79fbpFo65Lx+kGLF03n9UZy4rBcnRu8Ks2HaCy58m4WvDTo6mMqY/ebloIv
fvEFR+bOitxeQFVN6mReJN3gZVVIz3Z6kfN0O7ihAJy6aEL0IEtDiBzyO3UJ9g5c
pgujpXH3wck+gWFsO+C4IIpzuIBaBq3iA3kHJZxuX6wwB92oFXZIqgzCO0u/JNaF
/004WtVMu/v8WC9ihuCOror2BuDzbzCMWaJhKQ1kpisdb9coe/9EFZ+EgE1x9ccV
7ItKs3Im6wOqF9chtYD6OxBp33yujLI6MsgpvscZqIV6430KHizjY+wQ1IdKThrZ
5lqhH++XhElfm20C5cNDXj8SEZhxquRJP2Rvwq70gbwZjAIWq/41538rUm1rL4tg
l2zKo0uhT4qxRoVBKSrB6jyHE4MdKjiJm1J75zMqDtnLKtiNPAiqbevDuZx5cA7g
qiOjI/etv7kBkurj3NHXVsoRI4fS9Q+pMtmqHYH6dbutFAzfZRAm1VX+lwsWTSbC
F555sAvPKJNTlRf7i+3WUtA91uuXR+6cF8Tt/JKFHwZthddGiT1I3f345FcQAijh
SAxElWZAdHy8kWZdxj2l8/oPQKW/qb4Eb3nsvOQJ7/YSI7fCcO/1bxIIjQWF6Xan
vCAywJ5m9k2hyn/p1bSVZPj+voio0vXECIVndqyWAWroPaFRdN+yADaQI+e4jIUD
ASk1j7ZaQul4wp2sCnjItExybqOLEsjGpEXgPkM3i5xBoLG8g9xMnCy7Mbt9/tE+
a2lVKvitAZngJffd1Kd4IKnLzJqYrQUdywikp7XgWVUM3yeN9LM1pYRm3LPhDBCH
1fiKxHSqkdVLXuN6GVWZnornli1S1oQiiKslnenLW6uGhzNwESA//jkT+q3gu4sS
Sux0wZ3xoz56ORNGiTnM2NP/3M7r7Z034JDhUJ3ryWvccomLcLLU3j3GQf4N/28Q
ynHCkJ0odw+BQUe5s2kjrto2tlCUedk+XZjnSUdGpXi2W9Czuxfe61stJmH0HZz3
vbb8AirByZndLSsBjY/GvFbXK9ZAcKVMy7v+llXLK/9rgfpy/RdM8TOzXMPdcSaq
dk3bDRwfx9yyBOgD025a6zn8DYSWazF69Jo5stNriHCVuv+yYeCePlPhaS1rx+Jv
UTvAG1+c7kdRLRGPBLd7aclxIdm0mY/gigZxsyOW4OMA1niJAKqFrF/ee4n4g0r2
sIhiYPpvnwd89uHqdHzRk4jGAjXKSpyffqnYhUto1QlKl4Cnrdlk6BdBxTQyEuKI
vy/PcyAhKC7mnr4Cr5R8Ns9Qm8EEbsTY0RUYR9q8UvI0aWjMIHpkaYGKxOrBjmmk
kt+WUr9MykFsSPZLAdJ7NyDcYM8Qtc8GGM9nQ0szu1Yju4aAWf4zE9ylqAdFsm8+
fcVP8hGCRSpei+4tcBqZiu6JCd5UhTVxoC+XquNc2pS74SB5eiZqtVaT90SeNdfu
p48k0JY0BQS+9PuX7x9hZ8vU1pGrUZ3NbbXM96GQ+7oqWnok+tYsU9nfj7syObis
rwFj8P/FrgI8SvlGtooYhzv4csEtDRalUDjjhUvh1nVkYogyExsOfHA3g+HabWxO
exOfndBP2791wlnF2fksisxRFGF2Kx4v8L/dUj1t5KW8YNqwVJBpknBNwKZ+x4x+
U7PwDTmHsAPrv3isHRrnDIQjvKoQbPlSEbQDlnbFYpLglEKXPRl6tSxgoOa21hKq
7M7biFVLFyMFu35kQIUEZWu7P8ViKl/lL8Tyc4MIg0cDba4pdAt8mmwKMSY9nDrr
RD5pA1O52c+hk+mlce4VUFUQv7pS0P9jiC+hKxx2D+EhqvGYCJ7V+bPgAOpM1QR4
+zz3AB5np5nma/egYoWJYF7/twmOGIDQE7upOGtbh/OkFC85cV1GBAOZsc3ovqex
ArIxD0GOi//P3sfvnOL8CdapXLY5ZYLExSW8jKRCsjVOSX3+En34Zsk3pKcZBS+K
EN3tVb08cFY6s/DVo0f65qX7f0gRK3FQrgZzK0fpZjO/sNGuxBxspBDra91RlmMZ
eZeFAhqBuSJH5+S27N09+8BNhZpx5DXDDfxhH2j/S5BZDskq9VpbJaWacZ1spxhy
yl412d7pFIpFORmi2/D5AYMD7LShZ05OAdFVJtT7IxCllwdy60fUyv6ZXYOIRLzo
b3m5oE3KshFiWMiwurVXQyp3TbEUuDjsHtDkooP+SmlHlHQv7QMDqrnoJBf2cWQm
xoKlg1YHwOPX6v2qbv4pnkU4bH7PFcN63fxWibdHe1K3IBEVVk5/HWfdw5AkV7x8
jt19VEAN4dGkSS4EJGJ/tcRpz9Jt2rCA4ebzNBEgbYb9dOYii2oVhwwmB26qR5Ee
t1ODQbL5kxqn4ndIfdAlFiPqUXldBipxdkfWa0ubUrBxppJ2cM6N8lFVQVlW5314
mQZK4Idr0EGsPHfaORPt6WwNUgKGmNjGXqMPnIv3kQgiKm+YsNzBpYoU82RP4bWB
RgwQX1JJm5xvDWhkb+BlDtiTE3VBUTh3NOBRr/sPEsKuImMayD/reHTo9afDQBYi
qWKq1tbcCIimZNknofZopTpDyO+uOXJvoS1br0jKPNtROUx1NNJedNT6g2JCklvP
vc5sXpmNOeZ7hx3ZKpgNAo6tOBb59nMnZRiQoJnJughlOPsSQKQOKOpttU0QNySQ
pQIg0/hvxJHsuzbuPlMJ3mksUx32EoXoa98nqur8+k+I++VNq/DE2zG1ZC1zsgU9
eie0kERyM/wYrhxEKC7LmDDUQXS66KGW8+jGA/6f5HvvxsY7vWGMwSixokB3zY7G
lVSUyQJ2EDFhHHKLPWCIbmxzDCYVnCRsFzJHv+7tQjggdtz+9jTPHWJBKrrWxdOA
cAH/a8HtRf3dXRABwC9FFizWJ6dz9UE3vHgrjwId46par2QR4EetqGbeCNgoUKha
kyRhxA9+Vk7PazNIFt4HoWU0G7FO/3r3N7xZTuG7kI88GGc9Y4kgUt2NF4m1we/y
siWgsRS6nnGQ4VgmNIyzuU7yKkw3UNkTng9jIz32pZAmMSQdqLbNE3hyG2NT+8pp
lXb1bdHUQ9cEgA0WuRMhpLWIs4FKWi+Sol1kyWK2kSiexgXGPfUDioqEwn09/Apz
8H58W5DgxZEhsX8odHSAnDPDgGt/x7vNipBkMCifqpCBt0JlVd3hKC/oca4laKk7
M9oRaQH468i75QRRHrzNGoHE+AOW2J8Zurop8m6hdTZiIyyNQbOEYTWusfPrlG7T
rClQ7LjMtMh+iGhWNVDhWSQupugn6GwvdGSzZxCUs5n5k48W4+pPhT0NgpnEYivn
3I5XWHw6mfEKg5EucRlKOt2VAFpF5CmaRuu/SKl7tJYkbcJor5/zRUJlPk7YL0cC
6U5I1hRNGueYfgs5+kyL2QZ/V+ie4fivDarT+YH9nCibpddr4kawNFujr6xOzzN/
+ZrqeTDtR0glQaovRBAx1gCucTXf+CEmaUU4TEHCwlRHNp4ZjOkQ9SbcCT9q4fWq
OtNFA6/6TpDC0dIZHuhulrj9+Ew5ymqkvneweb3gYeGAC4dYxSAU4YwZJxXQrQBe
//7MSZqiW5X0kFl7eVHcB+7grI1Hg7b8DB3lmCqyFfxvRw0l0AgBXoE99O4p5Btp
hnyW664N/rAfMub9v3XpDeB2oKi+yQNxR04Fl+ZfkmyeiXGIqUR1E433fo2XhGu8
y8iLbRCfour7CaSyjgtS0Vwm+MSg3Aq5tQUlTTezJGlaskHVNOQ//IrRyUjLoKaY
I3VlR7vef/+GRkMvsC14zxn+Y79aKwhy4Q8PFt9kQE9MM2ZwSWtpbN/KHhTKU8ot
3r319wSpkHhBYGzludDyB3BEtsKcFI4a4bzwsSJnNqk1I0CLUTdwNXmCo/tQD2CL
2+FosEVgnxTvP7kKbPW7/Kj7S7mhmukCw/6nU8qPQDOZSTjEm+De8U76+aea5ZV3
4uXPGYzAp4ZSmLrePM52TScMboYSzY2GtNI2lxU5mYPnGpkiKYSB1rdaE8s7HgeY
oDfMaEzfARZGH/wN/Qs61i5M8YhmpfimqGKCEWn4AfURIhdhbrFQ6oihf7ClIsl0
WYlNp6wRkJ8SxEBg5ya8EMLDLEmrbApIZbXc62VzYQTReOVwiuyOleTwM/yA56vE
6cNeXzrb/vljzPISNhF6VrQ+wAU3nPyMZxuAHEAYOrqKBA2bUBv5jxGkhlFRWLo1
6wFrOvMj6SxRMU4usDsj0DW54LnmroZ/0NMlOfMFIFRJdIoNYndq2lIqc96px7DX
DHpFVchAS1XKcoChBCQinzF+OIhI5DW0cIFfppI5uGlKumE1jjC73WDM+9UniYgj
Q/F9uISRL24k/3dHzQDb4Y47pY1qzHNAb8VDVwCd2rx/S4oaU2IXh99lf8CAMU6Z
F5ZxQP7QrkExtXi027sFdeHPzzA1dvesIWxKpwJ+LDAOdAoe3dsm6aXHhMPRhecF
GctiX5REvhkKqCDtukNjAq6iTx5sPTaMDhJWioQ9Ex62yLzjfxjUNKt/uqWfD6l8
IDv+crIAUReMei3pwW0/fp9AGCFLmp+5ZTnR2W2SDqKR+XzhFvxKlYnvS+cSzikr
XVOwUVDVJwmb/GnW7IxatOTDSxquwsXiN/SA84VQcQjr8VBe187/trOjWmq5Bfy9
QeR5ofpEqT55YqrhHAq4Bf84aqH5E3cREu1AM1vl88yZgjU+HbbBFe/AoMVqnjnt
VSLjZVL3UfU+bfC+FfROLlf9FByQ45DhtYmYmcxhArqNfTfU7ehwJW0UZFfDxRf/
6q1SkvaCVg/C0JcZQ+M0ETI9JArOSnP58AdrfhU+mptUKWE44edfZs95FY0AkEOO
gk6OIgryonuD594K1njXSUnV9HQBk4l/2FJqwthgoQnXLJPr6cLfL9ng1UJ551gS
sLI0D67QLgXFU1HHWqVujjIWg/iXTvYEbYsqEdRG9Bd/ewuR/NYfOwmKE9NpXH+t
/S9dlywHMEypTzbKgR4rN2Rk7BsBhAmpQparnsrYZ3hspCzLpWdsWIG2zCKozrsK
NBosfk1D/ys/EvFeszHCSOe2OKeJKR1l4Jp/5MnbNXyRsqUS+YYAx8kQBk2x/iQE
qSZVnvv+bfLRZvGRKFVBMR7CBZDblFyJXJa3KwC4qcim1FUzaK6qpSYI2Rdmy3Ix
KhVs7iyoPvHcybq5xLMh1GhYA36B4P/hVxaXc0QrIB9TamRM0n0QvR6p/MtyXRot
6JbANjSwZ2NJ8QNHnSkSAxGKGv07yGJ/M3b4APrOXU2/uTLg5fVtIkO+AK+FT0WF
BBtKQ63OQMVT9JY1/V/gJY3meulbYsEtT7hg+K3/HtkAaoMaOLak1GXWAGTdGe8p
DkD70zZzH3jh79Mpv/edPgRY79zb43DXmB2TyudFeAn5cLttK30BGAvENdZxOKxQ
+eVnbyaLQRfcq6wK5JGAAtffBEYl+5+C7+A66o5lbceoWS7ePH2wSRXgkXDgZfWq
plsYtt2itDx6kdIgf5B7MHUhi+1mb+ux/AOVsHfBir2HOv9VjbE4l8Y3EEONJZwX
udaO71OA1ydY/mAwqMj6+IoV/ysn38sgIhvXBix2oo/goQLGDesd7XIqrnGb3YqI
AhbMgyWYQLZn0jwkQ7zDzFedJVNSUi142N+6tsC/A3QUdZMxP54XnSnfKJQb2ZVA
lO161RWa2T+L0/3iWgOUY1n5jfBsiLqKyIaKh9Ab4jhtjyYQKH/J8AkZVuC3sV0V
avNoTgrHAeLvCpWOylGUicSGQxqlw8RJvonzzf5ovGcCyaADAw2IGt6JIbFcwUgl
DNrPAkDiXPnI6vvngDUB/Qb6gMTwdiAQMzW0xvLC65ey1DrAz9ugG3R5ybUfVInX
0FVtJqNeHjkuP1Um3NmHVZsNpcNV3X+5wYGYWQc25rpqU+fXym12usMjcb8j9YdQ
el487N3pC0g5IhS3OS7exTFQ0RdzVLLIayuFq7MPlHT4U6t/WhRauMqejLsXuwQS
sEgy/iX0Ltb1Ny9eGld3/wDKIJaiNi20MGvwcOH+Ncpy4CWBry5phDKg2hhRyuxg
4oDB7aMO5Ol70McZ1unwKYz2DscBjxh3om0C3iChxk+wtUOiqsXoVCZb5haihBis
OyBH9KRdai0NEiPg1GdHDYYmLxPcbUwuzDjn9MuOPxi/Z+KgYeVC2XxXrRF42l46
6UOthWW/K52cJ6S9iO+dgnRzJQzoDQKBOyAlIyn9Y0dCgO4Ks7SbwwOAJFSLBgTc
OqMBW1iakZhclKjkkUI8FfwBi4nVvjodrrvCUr46W4mp3EHnHLzlfGN7yyr9N0+k
MygeMboi8lqN+iABo96WHXIORx3RyzFTwBBzlHaGVwVLF80V98XfxRDUxZdZyGZc
oWSi8A72B/Ecl5a8DHfdgU6kmb0GkZLBV5886Evoqec5R5Lvp8x6FCjN+eIN06fP
WwUP7dSbj3S4ghLM0+NJzf9ZsCPYvJpQmTVeNbgPp5aH/9yU4Tau+6GwI/gHroFy
qS2jW7v6WlMQwrlACZfJWsiQw1WQ/we2FqNv5AGGbRY2MlpiIfxQNefegVrs83Fd
xD73/YPdDEJYa0BuijJgVj9xQJPXDu8RYDmxFd3mU4UYRn3jFmObAy8AKbsPsOWQ
1uncfrCgwhhFLu+QOCS52deFOQDybirM5uuuXqNJ2Oc8mavdWSD06spFuLEvTmjk
UEwlx8h4aOmFNxAXjezDU2Ivgebgy4aidbNljO3zTQTYeIpWL92gD/dojQqabzPt
gnnE4FIuuFdorKWExi7xAVq9jw47ES4/BOufryzCkF/inGJNOG09AAMbaam28E7u
0ktXBUfTpVEvHfJru2VbI/4m/Z1Pfl4fWScc+6kdqRtd1rjwO3WAHNkATBltXeCm
6IkYw+oivMhN3VHvcdsX76ufIusb/rzp1i65pTJ5svOilFYZcSZOR4sVPnltlbP2
pDsNGNtkleqZ9C0IwyiiIIo+B9duQ2x3WMuqiDMvML/9//FAvAHXtSV/ffoLAeyE
+d0DXfY5FMxvHoBCoqsqQzMOyUxjgnMPpm4c3r2G2IvyBy8LEN8xviw/jdxb84jJ
7uU5SZQXLOwNLwiiesBZSGpejlON/Wn88pGjNhXUTEnVg/9OQBOijFPXNQl2e3u+
ptkHmUw20teNvNVHrzm7IWkfFuTGO3S/xxzfpbLB55oXrxd9hkEVEi9H59P0XLVm
xVDpyyzkU/8wpzDtNbRjM44eovqrGjcKzNHdvxsfMDHDMau1nRoH+uAIEt2c14c0
sfCdCT4bkTTuWzZS2kvoMlZhpf45poWvFDKDS29N4NFF9rNTyej3j9lQevvpOC+n
B9Zc7FnKQiCju6dRDeBZMVBV7hFFUPaxU4FO9oqVcHLno7EHmpMCAflOxkJ0Eqsz
CiNNGX6SBH74wShHFt3jzBQNoytH6/XJa09EqxxJL75WMs1fBtLuExhsllok/kj5
DDNCSOgYO1r4DM5LgGmGazvh4f2HXtjayatQ5qsDReeoDLV3s9zu1Oc/AoFepr7A
vHzMhN+nGnpI/NbjwosCUZC1++WlcWtOG5f8PBW7+e3X3w5Z6sU91nszAR9ZsMIK
cmgwy8djhcPOSFYgm9t9FnjewUwv+uDUHWQqt4gLQOUUwKRjC8xz0se/lZxgdjnx
AVuS4fKZU9dFiCpI1VPWjBPA0s/u5pUlRnj3qN9vdAxJpTysLfkV6ESEcmy/PRA4
k1Yi+9gHrVdnjgGBtCGMpYvuY/RP/D6awB/yvuxVvnU+4sHUWM5BcrkDr/GZhsFi
Wq7axgvMjAm+4U6bGirV5idK+mA43NqUYbaonVXIqTXWoUn6MJ9DtWMxi5+rt58S
xOlqtYc5+yZ2lJhB+2QZNprsKgFUFLKPJaHIsVEZkYgnvi2CxiQwxdKb7aaC+m/G
s1+bg26xP5CBCFrwKBMiUTjfDh33K+j6vyL2cqMkMMTTO5fL0I7EXgjxmsrRtCJe
jSwHDzht5n1m1h3BEzfefItPdQukZln2XSz0iXXPR3oCpMMCNZ5XKr6mID2V03dm
awiKCOQ5QcnAD/93qFzoi+rKk1lvV6Qx4+vds7ubl+kJkSPVUtEbXoVkrlFSSNrk
BWj/h3bulTxAIjtP0w9LrjfCw3YqrsfPszm7Aw+SHKVNGRsk1imMqpN9UJZOQgqn
tVAlVQ1d7K35zHltksI1T0o24rFc/eeAz9U8X6VbZjR2wmFyDZstOVy7f3lzXWyB
cwxoC19o0yhiVjLVwI+DhDOz1C2SfbZWsEr7UvARCSFChZaBmlfUhmygGzur2XaH
fNJQPItkkyQjnACK14zI9bT5PZFc1QI/p8Kc7ZkO9SvkvkiugRFdjsnonEz4Z4J5
B8vVyoH6iOTcLps0EzwCUmstP+k0SocuprQL0WQABU1kj1co4+mMI77JOmfPaHvo
K2n4U0eXjwoSUSLxjIJJ5LzLqL/YYEnz7T6eSb9EJkMAoxYl2bxY/a91ngg+Ninm
toELF+fLwJRb3e5EF+NhEPY6mfvJsgXxUcsSTDZOflKzC+RR7a4LZM6WO2F0PFOv
6mt6dVA/b9fJ7jS/kdpGZwEwZnOK+NB2AM25lZN4hsDy2UP0igcOoy489YOMx5F6
gcISN8rIMM+MB8aFJ6dTPI9Dclh1ARGWuX0aBFkIz66+CnhCR95aL9q3ukTb0xam
8cMDyoPx+CqUUwxiRLy0KkjjdI3WmYmcM52oz+qE9f3UIP5m6RaBAWTM7Mt63cYD
eE6C/glQzj8NhtSw8UurvHC3Bngnw3vscl2OpNz47Bf/NgclJmtx8opE45HE+rI4
XuztG55S7lrNeaD2RGToxXsxHFkonb62GnNtOqVhYrdlIAFwbgyoJL8PrsnUY09z
6mzvE1/E38phett34HnV+1Kw8lNqN1G8NZzQtGbh/a70HLkSFpGjIZUivb64utVN
qSqpeyRg/SnHWzdTEv85LxEm+xadfBiW9Z9cTRroEGRkvnCzv7/q9hW5VT+LOcbr
3mdUZZO5jEqZzGFPuRpuYFqwtzE477HJDytuWRrmtvuRpjrRahW2eD2ZO7FQ2nfz
VNfC8m7fwvI4tqQIH+pFAE3SYKH55ENzGKSvPls1lFXmSgR6cnW9rzjaVx2HUCAG
Ex5/xkHb8D6PHQ36ZJInHgRHIftg1Z83sJrgihCFifphoBKbEdfQvhIMLr8VEJRq
H7JIKL6tEYre1Ba6c9g3uSiFjCcAzVpww0TVyXA8FZKjkbVY1PjuX1RhdEtm4aVW
EAhBHFISLZnTTWQpT47IOtSfps+r3g3i10IlWJk1yAZ51pj9+MdgmvcOTdw+Xmee
tx+UuC20CzVx5N8L77esRw6fOzdYvqes+2RmRHhPJJLbBNKBfXFr10oQHyHP8X5U
aLShh8739EjUFBG8D9oZmimDSg3nGZziVGBLeQIgCvoEZzl5G8+fOXZ6TUdXQB16
bdFQw2Yjxe/wNOd7+8eTLed4HOjAL69jukwm125O3HINMC12ImmIC0egU1fAKqWl
6om93ewOtFLdUE/KLQXVyyfs0xUuAJlj3SVNFLP4q6XrazlB8r27UrIxOJeQoe6I
GX6PvgAyxPe/ekF2uSOdO2fvtrAr2EukR8qEWY9VxhsUS1d99DU5Xsdh07a3c4hH
GN9ZN3mKkKSZ03YgTGuSaOOf9qAbU75yfIich0sN7gxV91MzV2ZhBT+mtdZSETnU
0iNEyt+rcQno2nxeVMyXZKPwJBIKvGX4H8weuAaKyo2+9xQjKs3mGhcKYyTHdPUS
Z/m+bLQEIThitc2eSV5wSixuNNDHQbAzxo4LCEkZNU2FdU+vlCt5W9II84H8zXlg
ApHkjb+nUFHt3Q44+0z3lwlJQKa1j2qWXeN2vjV1nu0X6acDxw48NJkdpygsfuOy
F/4xuV949yHc0QGPpAN0/vMFVLwzrh3DAOIypTMfRu2rBcVtOwR6WhVyvcpbS3uc
wCjfe1KPZAc+biCdisKzVuJ85AyNwbafOPwjt9K0mcOctslh6bb1zPaJgBBXMJVH
NmGb/3Xf1lqSzzm8tG1Fh82gFq8SY/+fON6fmE6v2tf8oVhpGVBMM8PA8Yv4bVm7
FcU5xeNt18TIb6j5YKWh0vxgs6tx9eXFLFVW8INmAQdd/avWS2bojiC1zhnpYe2d
nh9ij5rmh8eU0/nBwiSaC9NYLoKAWQot7+AWnr27yv/WhbaSr11/9xX1qZb5S+Cu
+53vU/mUhPPxgwnPJ32RyPWw91ClUmbNpWmWO17JA/qFbfdzh9tGuvQC4ajr4g6g
QfYDRT+dicoJoZhpD0x3YJiLuPtpf1xrCgSIJY5Q3LCaW2FVKuQM+23I91c+a/Ka
35cxHqMJEj+5VoPZ2CrNwi21ayRRN2oPoDAU8gWcZZbekNmsr0nNopwImdeEi7Yk
KacXCJ1OIP0+zq4gBDg+R+XKZQwdvSqE2hhWLL9L4kumh201Jw9vv4GrpxEZEOp0
w7x4S0kWuBBValmCtzTCkvUak0WlaxEitHqrQ/8NTZUkHcbiSjUiSTkEI83glzkX
9l/jltkbGV2EE1gsRVbeWALKC300/47EWUn64ru/jTYX8vpDcvZV82/gwRn+xNCg
yGM1XONvrJcOE1yL1B/Sp1Dpl4eIRW6OAtoSgxE4hwXR6wxsTEfNmBHsnl+MwQv+
go1j9M4dH8eaHQvT5qZRNjG9d0UJ3rlwj3MyZUWKsv4ft5bC9vFSjtvL8sBfP5FA
HiBYioGzE3pGsXymw/n+nwPe7YEMa5mbbpHcS/E34lavPQBHiLlrqJguDEfJW8L3
mQCcOR2XkkmdJqN+qcHgylz7oixHCK67bo4poF5vGiOw84Ou5xE60EfBk9isqGl8
ECsbwR9wGn8X5L51LwD8l/ez5YOshHdmLPJuHTemHF2fKk+/KokuO04IA825Qolc
pCNVEHiAenxvMvXmf/Wivgw6bE4uKSGU+KFe52DzYWx3cpDZdR3qaNO7IifdDo3a
ok75LbzIlFeDc2aaHip1lsachMQhA5hQQFQb6psBUe8IYKBBf2gozgOjTTmuNCxF
pVfov1ZoN3vshTMewA7U/GByli3KkVtRqkFaDUHk3RLg5GN1DX9U7k4u6N25oldF
iUeoWRp43rTcWs9EgjnVQDUpo4+H+z5e1bNI02JoJ7mCxrymkY4d5Q/ykjWuWo48
VwsWxecFoXDMcqtw6MZE/bNLLkUjdrbtSdJ3R7HB9QAaaNJKTUjHlYWaW3wXkXXK
RLaO5uu+FxcedG2M7RK0OoJbMVGBov1+DdV6snZmJIMUwdmN6Bxbt7SnK/Jnr2oE
KudvTS8FRaQyi3VY9LEcpi7BTvgTex4fFqE4odXkWwTTElZvkUQ5nFBbgS9VpcVA
iMc8JCID2P75kUM6Tajo3IabLBUcfKrtHBOyMm6cTqarwKtTZmM7JtsMbhboCtWi
IYikx+IHC/jXZoFI78L/4SjQwegKJzZyC+xysvbSwbJR6zS0NbjZhdNNtDRay4wc
OdpkEEPMb9/I3+Z7Y5+VjFlT9WiTRhjmDYVPmWsGsVy8WeJilq+m6LFC6hEtAW49
ICYGpU+JJBlQeso6TJxRyx7LhWxw+VxUBnypgfK6DJimKYR5Twmei84kJlF/dn85
kbPP0P0TljJZ5yuDsRKA9te47i2eptVzHSFqFZkuyhw1yA7HKjq632HlT6zIfM2s
3xV16I9f0fuHt0+xrNe7w6QkfNFG0IVLJM77V5SmtkuJffraEH2XgniWgTfuTPDV
9CG9yx4SsVQ1bFKCQBHyI+Pc2e0VpdT8IY6mOKLXcZnwx3I8aGbE3Ixh+7o5wx2s
UBtH+jsj04QyyBoT8OrZb36iuBmYD3upqlhZw8hnpYfBkAWmUSV/SMRqVGRSP98o
yBfEKScATt7E1U+bSn2W9OoMd29nGGa/MlCIUBwcFxZP7tgrbD+7A/TAci39tXNI
e1tdfdHCfyBRzAf31cjEQ+ckKXnXl/ggLp/ba7m++0up2bBPuWP5eW6VAmnQH1tg
qiBX9qBlqaAvwkhANbAAe0woylqWBBQZ0YzQnr19jld6DPbC9tRm3xGlP0TxZd7G
FKrL0DiaIYgUDiNEZ4C6rf8htFQtpmSsYtqhXROnEljRxJXsL/zvo/YSliv4qT+I
7b4qr9ODj2uoY1rOzjp+HOR6gwBySwo3r3HrNwaWoFKaB5u9eOqO08BDt9rCLmc1
dJwVY/nsOTOB4ra6cWNlp7/oUurnbMQcvnjsHb4tey88VZmUF17kCuNfh4nnekKU
en6dn1UlXbly8jVJIvxyxeotKtqpE3DfTR33wjx3E6i4173f9K1Ljt/BkZJsztBz
zKwtacUp4+n94lZ6mUZauz5d2NSWvqHqldd4zTVLCk6qcpK+U3ezixceSb7BJno3
CftSaqEfqgpaTgmZDbmrv9aAvwAGITYjhF/EBC1yqUpNXbqcN6muD4JvmbVrwFLk
tVBDV4Uj6VMpJoUmPne8EC3dTu0w4Joep6le4gER8I0YwMpA1dDvc5v0T7MZjl1i
vvuHX7xaOCEDKlYvS14XIJNIta8DZtSh+ptzc/MmP7dL3ysr6WWir83aJUbOOynm
vfXDimnqDF3qesruf/97JKFEo7OqJS04QCmWTBdNlKFCalNLo8dDHuJybyl6O9QT
3uqyLn/M4fXFY56ct8EckqKY3+zJkelMJ/+XtQrFfG+VZ4l/A2LFJaoi+f1jZgwt
QPH8T3CG0HOHdjw4Te+J/XtwpPYXybLa4e54i1c7kFFZNGLRpYezF5SyCTzXiHvn
P1/THKPSYSrXsav2SNEwxFNBM074UQpYLdGn5bQpmgnTyvmiv327Nd3uWJYhbOrg
HRQJrO+qZ8oB3uEZDymcp8vV0oo3ZZFOQu/mrFJnTUZqdvTedN+vZzkZMAtmVaor
JY5i68c/C/T7tKXO7z4FTEggrPO4kQcdGRXc7T6wkwo1PZHMBP1omQVzTk16kpi4
CvJjnlWj3Umf3L1SW+jW8MW9coixv2uaPXFPa1FGOE0vw8s8LCFMD0uMZsdcjAO+
mojRJ8RlDvViYkQpUIKsZMHjIl1oUCGYx3zza8NFZDb1bBULS5shiGiIMj3Khrr7
UJ66DNaqz7qgkj0+iZ8OFvuLv54ErMlATHWO3lRp4lj5a050Aj7a2Mlp4caaAd/T
ZZDsrTpt8RpzRINewwxeXlnWtKsgXMWLcCmE0nEIjmLcBK0MEoNrSOiupkeGqQzB
TLnYp7FZJrNA4zDlnQq1ImKzjv3Ny7YQ4TB987GQNEjFmJCWYazTntnvmev9ZwHo
+8+uEgKTrKCVHyw5I42rvhuruYht9zsKdbUx4bzzL4glj1s1+d2gXEnawIt/dDp3
+pigthmn7vAV3vfVCIijdpQQoEejaH34dZj4v6tSB0zDVHltUjr6RCmse7glUL3v
qSvhEmVOovb+VHEJXE1WENaUecbhWsy3+hRao0F9VJ3Ef/5+2xZ2BQMXpzleydj4
L+NlRy4q3gkwKO6gotCJGwUzLDWXvezn3SLIqp5+mU7Pwo4RQe63iarE/LYLbBMo
84YHQcMkXc4pcQmWu7ePR4MfUhWDkO0yp7IxmhCGy35K5b9Ia4EqqjYWHgQuiND4
AR3cckWYluR/pnHsaGjthSrfXA6lM+FSgrr23pA4TzABOwBRsf5mT5zE38FplyGg
gR8NKs/yULdfkcM5Wfpc94oqzUArbG10A1w5Dc4gjewwJB3kj2J//yCaK16O0/pu
YhSShsM2kr6MmyB06FW5fS9wmT/UHU3AsFzRgg1sdw06ijyRoowhSVN0dUttce+H
2sXt+1wisnHA+zaO7NWH3COenqjUAeSFoeSkjsgM3+WT+JH3kkBoNCRiAnOwItOU
1vA3+WZ0uNZfEdWwsZ/a7U+FdBd+PgHRB3uOe8FiTtQZzaIxm9B+0+u+dflRMIxU
vNo4kYngDIqs+sNMAh8j9zqeCPOR1UxP8hk5pPP07N+miNh+URIiigvot6enHO8q
ad3HBTND0Pi6yHv4x0Xv6LRzF+wr4RYzYZpJx0tsop5uIiK09Mwib//KtwDAQtvm
ogx5Prb3ohwKyxLN7UICb6zsXDDoNJyB0SP4Bs/cWP7db9QbgWTgZgi+pWdRTJu3
PdwGgs4KwBh3SQVi9hA+qgmHaTukDBbBsvrm7Xs0pptQbIdh7nlKCSZYPGm+gSwq
fouYtyQwRUqm8pUoyrfXLmkQPs4dWx6tdjLpDlA8oJidNfyxrwuJ+XpRJyq5G2lg
vHWFzNWbfz+Y2/mtCoEiJW3PjZcpzC+AHEhyHoMOlh5PQ5fpRXdDyTAQIrYDy/DP
j9QQdzbF2lAQOyfCE/4OVpsAuPM8LSbrbwLoBlMGnqffcFXF9L3ryd3kTwLZkgBo
CpbDzf4Z8rFTx4bHfSpVD6LqXRwMCmt4Ud+nHMUha+KEYFgxfKVSruKEzRG9yYOG
swwpP6mM9qLnrz5q9wjSSEfnF1uspE4A1KbmmoxU4ob1NdJMTAkYXX6pz4qSSRZi
/YHX//DxvDufaQfcvlmCnPDWCuVe4HjpHDELnTL3gcsCH8hgcNT+0aSltabxQJcv
RByGqqr9nNjUjjqAY+y/KqepjKXgL/KZDoRpcmJAqXEBuvBsAQ5ijS3NLv8VAR4K
4XiFMl7hUKAYuuWcmyRyl0UEn6tmw5fTVvE9BcOHrsbiuwsd9yOqeyYSTaqtOKwu
arNmaVq417XlsP1XpcRXdN+O4zrWmoB47MD/g++FRJ/gN5If1Aegc28akjPUGVBb
YKcYiOPyaAA18tXPEt+9Dac3mLZWOe/cUt+kNlbBgmUU3mFuO9mL4/hyNEBhWY+Z
exeYcOW1j+Ewx3NDunxO6nPJ/Iz9PgFmyyjZDUL3HtIXGwSvkNFRNorDcniWZjUH
yfgk5C2xdGXxSOs/SoKMJAwlGzpxTxU176fUfqVqzG33kmhSYgOl/EleyDFBb508
Ts8aS65IAi0svXq4+N6tixayRxX0ZVZ/oKF5ox46+lfz9PIPZS5FRzIJidoZh1Gv
2fpYXNLwcUsfi4obb6dfOZ73jc64Inwxes8QBgYQqMIhBOeZ0RGsp0Fe3H3DzWcP
tO2ishUx+XMoE0FbGmAmGtU5s2L075a2bwwAHqoB52+kRvpoxzckY8M072ncFIhR
SChFnQIwKPWSxNjRaLzsv3BCb4+PlUfOfA8vM48/5u8aItfbIL0ghqvhyZYM49t2
02YYSp5ovDUgapjSJC/ac5pNDV8qkOCZE+Ud0wMuK6fyKSqh0mvf8zAf8eUwqpao
V6dq5PU8geMKOnqsjzIdfzRIXVIhUHoM7++d1K2E4yV20txjSYSbXYXrXBiUOCRr
ZtI5lkv6bp4yPXtDVdOAtT+RE+wmYjaH9sguhYLF6OxwJcDNOy7VrJwS1jckbyUD
pLTiaDVrypth/kPLMQTE8Tr0CTd/lTeHEqHbznIsNCniYc8rWrAuiGbmtOPQXplB
7IaYdp/z3uBbKj37Liv4h4QhGBufn+sA9WjO0Vb8EPQmjcfMhhWkb+6g9Jr+Oxe1
n7OGLcjyuMHl55doVD/n2CgWAQ26+P3FizYkL7xxLdJXE8FjDR3CiBRaKw5tcjws
3alqOAoQRclGGiGH/ohjHXwvkSnFNYHdVDjZBzs2Ob8lXxvwPduTwS7FCpv6W15b
RpmbDmmtr1vvOiR1lCFWfxkt2XZd+CRXFUM13yoWaNOuVK8dFOybp8rx/BYiaDe+
8pQuiZwedqujr+tgEcfE8SabwgweeFuVgceSt35vwDrtQldqkwHJQtw6jMzBbKaa
9JtT7t6iPvVIUvyfEKI/hEsJ1r9SaTM66LY6ADRq4mfD0OKuyItOfPp4W2DGN4Lw
wUWkCpKV8vR1I4bMIr7OdZNRwXixPpSFi82/bN8sNdADd9xRhWkSwkz66ptGKCY6
ocmSdoEM6r3NSSCwfoIPXhfVG9ApWZ9LeYIL2tZokCVS7XXrvYfA2DsQIe2ABHVk
CH8vfouaTkdlpdx8np8qpFLpliH4b73r4R2qRU+wS6y2TNeh27/SZ6JptL8D4k2X
WnjFgeGdrPysHXIYAq+gjpgafs7qwKkekhtaWjCOYGQwJkLou8V1EVbDxG7UQek/
mJPJSRVrscmRVaFX0kjL8GvVCQI8DJadbxOepF0lx56ajnAFWYRovINWZlMfzbqJ
Erk3cwMh3dFh1dSjglou2+XOL/XDlhXVEjF5WvBV1jHBxzVeu5yA8YMWFsc6JONZ
TgqRH/mhFegCxH2EQypAUxhAa9kvaGjuUPUf49g6uupra6aSKjsD5JA9rBde1saG
WM4iy1Xka0/1Z3I2O6xXllcgn8HSeca/9l7LrS4ekrFju/luELNPlE5q0rUqwfU9
EweOW/M/TA1RW8RHw4ZmjzIp22krAMIRWuqhyVips4iDEIq+mFlvMqiCDbWIi6Ui
7dnBCmN722SG9pDPkBtU1fUwIBjKdCjTDbpA8r0w+qfnS2k4bdNIoyng4n9v+SxB
btALluQwx9fVbYZe+nCU565tg8JBKucGpCf9KY+aXPfOlrKTPqhjzmUQPfuS60ui
Mcw44FpmoCDwbAw0Nky6Cgiv/oovD1ozkG16WiBAEi0lOugwJXxl9vfK2Hpz800v
i31vV4Mi+1JzfqfRjYjp/UTkRneRzlqXCqM5Lv+YaHtqIT/4BKH+t02doclqDF+V
6uajHoZv+YVkFvdNE1Do6pSX/oDGSiv2/PzZD/eIlfRZ1VUwD20Lkp5cTNSl3CJP
Y311o6XaUZ/9Ni1ODFULiPj6hchArkXqHTfhPe2A8VyO4fBA2D9ny9myRnfhqr4k
vTnwGbIQaSlasSFcUeIox/J6VjYqxPaVizaW1W5GhFvf7pjsVVN7Ac+PQCaq0Zoi
ba0EZX0o4pTpGJiQvcum90f9ElPOpSG4GePJImdxVdlltJiYJUIsrVr0+JZxmt5b
MoB/Nb5egqGkBi4CIrdkKWwa9Kzpzp0W2uy4MfVdZIoY1L3Cgkq6wzpQUi2Odnai
LLiNwycAZRL8jkqQ2oJaAbLUqplTikiGl4tegdVjLJEw4i4eT6M9B8sxmNOo6Wwx
+MxppLbWGT+HstvBTg/+F86Nx07C/L4Qk/ZtG5bJ3TY6lHTDQZWdahS8GwyLMaPK
ntpXEvaj3YXipF7X9WB3xdO1p8vMQtUGCdUGRixoBXJut1iiH0BYuey8UE4k8RJo
L1uW842pe0wX7lCh9iLo/4P8ZYE7l0hiYdwdRJhNkOH2Ki7oBLV5sGDq3Si/Lzls
sdpUcf6dKXzfe6I6cA0+V1QhgKjfjfdrrVgKMVvz9hxJd3LCMmVpzmmunKK0/+gb
dUy+jPeUsWuEmVNYS/Cxpbd+Kz8VsKJkAx3ti5iEv2/V6VK1fbDOAvMJ29ca1j8B
mC7T7LUapxYTsllTHu5CBeRF6uQcs21B69TWjPEXXuMSffKp8KNKr92QY6wzm1hL
3pU3kVfInX3K554yiUIvcxz0AZIou1C6OFZCM7rgPzEb3zyXYbYHZnRz425MGLHL
cvwlV3+YY+GTAujyYjRremFQnERTfAwOwdsEId13jw9c7ifu5FkotOB7W+87CaNR
j6Vf74WnasSc7KXBBuk+fAse1J8DJTGmoRBPTiZuoa4eeKXr1O9MeE8FEQdguMbp
XCW14GAyAZYUpf6CDgMwVN563Iyy5jIBde5cP06iHwbMBQ2WtnllMPBoBWceXDqS
qKzKybqQvE+6M7OVqdyP4Xh0wj8qeT4pDbt32dS5egjArGRHbhWFRVIh6f+KI8pO
MLTSY83YC1ZhrISlM+6awt0/ui140v1sFEFPDdNeyUYe+HoAl674Ltd6kcxcNQQq
1ewoUiRdHLglQ3O0RkvMwDW3LFuWemFq0ENaza07L0phRnjQjj/UFzGjL9VCb0jM
B9lr8LLJCg4XOlEEgplqWSiIDbvohUmWWdscVpNQsqA/TeSx2cQwavLebXUoElIN
awZw44mtxdNWP0Nym5Ygp7XYCqniHKPAtRBlAYAVpx+710RLzp59EXDd2VHbQZRo
NHu4tA59fBSM8J9ZhM2wA3Ymbr3HIVdv2iACoGp49PD/XfCFF91L/1pw4MojybnO
IpRcZwC92O8h1XHyT+fYxpSGeF5BFCjlxPO1UpweVCQcMbmMJZbLRkEqmnL3zSst
FYygxdLbhK3p4Jlv4JhGOVHao4ASSygy9EE2688SmcDxd/N+PlavQgwLaJ3n0XJB
RcHifmwGWDD0QGESbfEhvPljO3OpilFnrAGbcMlxpBLzgiUE0gNb/5d5hYvCFV2t
AiSWdVyGCyv9pQVFHmMBtc7HciauAQCE8WLLePQmFG0toenHY0+qise4PxMVvvtu
fnzXHyPeFAgJPKCrcHwJEvFDqgOl1EvHs+AJzhIfp0lvE1vTXKpkmiJcM8fVkgjB
dJWsX+m/+Ij5bM/h6ZaNwZBZUiuHxEvpINaIL4m2VX4LXrH6SPELfkhV5q6h/Rzv
wpOGMTWs06zV/BquRvKrBp8GJYv4ZbxwGX8/xW6caIgQ6BEllO/D/iAc3YswHTtZ
pmDIhza8wgIqaCdYWuroSR00LgP3CafJagLPYUH0MLA5NOXzGAHI4z6M9J7+mvHY
DKEssrvgFJ6t1CXTaumh5daE4b5Q1WeH4AR2CsEfpINyLESvizGvZjVli1tubBXh
1d7HCTseto4sOYA48mhjRzYOnCoA4zbKQGr/bEFYQCi7csGpGvlIeE1p8jrwfnoH
xUWLeZVgU8iHE9NoSpKz5sFzjv+ruYRnq85vP7yJt4Sdj4wpF3oe3MZ3NFcAYht/
idNv3vJDBtEOMRQZIPTkJPZZSZlLQVjsiyywq1aZ/IB0ePNiMEc1kFl+zS6es6Ir
s1UYWj4BTt3xhUbnuwxe0nWsK2YQbp+PsE+LA6bj2VT8boBRMjnE/cN6YvcJcM3d
hKAXPrZBVADwjuJvX/QPG1njG3k5qrsY+Sfk0xb5K9O4ZqOFfqwPZVtE/i8xYPBR
VNMYQa3oUp0rEn9lZxCShOezou/NQWn6P4w2JL4B4LbYgy5oZaPAxnrnKuWzKXUK
Xm6YO0QuckPwSdlbuHgj0An1HnanLJXtvaNk85BumCAnfnpcshD+vKkBz8nht+eQ
Jbb1q5OjTU0tHAgrOfWX6/hifff7DvCr40RXT50ew+v9M/yXN8I+3uzNLCvbzjdk
Q7llWVr60md5iXjNh6jHOrUOIMd/zHLbOhrWef8wZ5FzHQsSdQqepQnU9r/fQtny
8KnPd06DyYgOmm8rc6ji/ICwqjHA7lZ4wQgXIIw/C7iPlvGgAJD4xXwqzux+HbN1
G6f98D0IT2+SusSjFpE0yAs/r7uFD2ltVlLWZLLs5SSjv8SOK7JCqxRl9wOus92M
8QyBFcGfk1xv2syGqRKBfFSWZQRsjwJl6+vu34AkEzLOAyso9oRqdbnFJlB1eC7v
O4/R0hAp4popj0w4gFfWfdcSTaourX0pA8RaqsMv/EPy86tZCammipEQAHUuWgSc
EGfcokyg0XwrjS/ZrlZObFEtcWc4WFm1aVD1h/GullkbtYb324c9Bl8i+OYSkOkK
2HgYnphzKQsd4EFELAxGwZjvATZi6p98owM4WlyIxa1XDJvVRH7OiSntVOxiUMWl
0Z3m+aRawCT+YZaUe92mjpfp45mUIfdQAdsQAJhrk465gw17bBhOBYVuAp0ETrtY
azMgS3g1t25vKUDM95ghqRYOAViuTlL7B33b/nl5Y5n8EK2EfmhTNI8L85W4BXB8
FYOyuoUH/OdKr4gPK6IA8N8WpyN17P0+5Guqiz1W+Z4pjfG+eFdmz0wwV/jszcWm
mLWfnvAivkWjA6I1qg3ylRTqVShezv+TqlOpkXDEEoSXUQ+Y/pWegxV0jVcVsKIK
UhX2JKhfxPsk5bNNHS4EMQyrP2MN0nppKOpLhPDM1ygMY30mpCMxqYLyHs7KmbNM
KLAM1T2LnPR2sEfsWtflBiRzm4VgUCwpnRza7g/BK3GGwiwjsV+xzy01PTELl3Cw
UzZ47cZQBVXQkdSZJjmti0M2AcXofKaW/rhjRBQN8XASJ9HCWC5tGO8bG8gLj41e
wRkUshQn7utPwu+rHhaB8e1MIyxZR900qJFBJ8WgXw3Pw6EglBHxrzeuuH3+ILaZ
LNz3bTnVty+9IHzrF/ZYb+u6fH2B/Deex9NBr58JcHTg0dbp6cOxpvNgZuJ8ORai
w9UKN8Aj2mz3e+QH5fafpULX3rXFFWJhk73buTEruHrexYJYhaoFrDVaupiCc134
s+vylFeTD8Cce7rQUXuI3rgKx9podmUiLiQ5aXFrdKGYq1ByQvKtOf8HtcxiEayQ
9EVq/5xcL4uwxny+Zw5YrlQOasnU7FVa31Yb8R8v4zpZFHMVHfcztTmQPKRDfTpN
1svrd653S6K94Y7kbmab3YXRFQ6sWBUIUbcuQfBtVHfF2aUARYyTPMscnaCVBBSC
VZKA8CNWAvjh7K4MrqauQxOk9EbSe/mr109gdoDqYs/YpphocCLKzyReN2s5Ek5o
CUGOh61JHM/9xWlqprN437qdAv660LnDZXR2UXtKqoNnJKdKT8pAUqIKbBadHU6W
pI0c8FpEYIKfPGdSKhIh7x8CM8jVTb1I8iy7EA6NHxXFO60g+NUVLovb+UoazHmK
cTCPTzkq52N/pozieZ7+WaKhSZrZBdtiGJhckqKx4Po9veuS65WEHnHPweV75x1Z
JdWp+OkZn0YU4tAWYRFfomwoy4eF1rn0YbJLK7jJlchcv2WS7NNtS3KDc9YKjrOa
3AUqcbVpS+OjYf4hneCJYvZBF9aPuXB9a8As0+hK7tzSMBzwBu8pC2lA3RlGjtiC
c9u2u5xKLXgEFwbhl2TMaiIvzQjWUSz6RN4+tVOqR98Uh8LJqbLSLQI4FEsmCDSK
DCuL+6JaUa6yQRjAX6RxM8jKpBMoCnMryFKUIj4pdwR5mAyCdjEKpPDqEaQc0FYK
/Pwo4IWWixkz8zQST0GL7YaQJBrsts7Qw4oGw6rCIl29B7mdjStu52yf9ibF553m
uTjEJnMZqLWdylH3/s7NBICWiCi3nAApZwZWC8PXwdIb4KgtkQPN/zGRAVwAKk7D
PLgpWYSAcbvvuHvGH7n9GRiyw/UskOeHnjVdN5c+771T0a+Hm3H8zw0jD7tBunSO
Tq0JVJHf+eVFOgZNrn50E0jD7M4HnGB5zES+iJtFmgVSo+7zsDFVDfs2xLBUTel7
oWbS+XpJN+kza0KpYZtIyyGZKC/M8ZFht3Q9bCcdJ8CoxlTdRfEzcwmi/ucD+kRl
iq+p7Rbov+vfQwxHTFG297SB+jgXBd+oy/jf7Kj9Y27abHS62R66IKFNiXtJL6Cb
llWZ9pEmqFfZv26mOuv3GUtwXcnMD0yVXsv/9cbrxoj/sZmalHkEjp2Yr2UlfYqW
W/2QToFiquLbITr94HNT2M0p5mSi0zlt9XrLpguN+z2laacKcwyraHvxXDFhYOnF
lYv4wr52FbJCiY2te72VuvvnEjHYUi2L1QH/VV5Ren0hq6QJLYI/CBHott1HDWNu
7eMGjH8C3SOseSzroduyJ2FZhPhFboipCuiKU8nnbZ59gs7anix3nN14E4FDkf64
FM6Dju+4b20mo9Wby2tcXXlmnh/Jq6sCdsPDPvTcs1qd4I8asyVTJOWmiUl8t2H8
lWLD3IYX7x2vXt3OnqdmHzoJifC2d3OmwloQnE6dQZRKIHfHLx3SdSaVxZYdSHu6
WZMNaKPpkZKDqT34I3/CFfPL56z3B45uZaPr7076hjyqqu9PGkqz3WwVc71/4QVD
6pAalVvdr5WrPTKQQHMv590WT3t7CSsBRT52f309vPDddazF2X3CQURup5J2ycuF
swaf4ALSA9v+CbzpJl4oTy6+TlbKxCLDzdjzCqvuTPTGYDOQ1L8IDkOGRq5/EW+g
lopoWVpDn2I9N8B3Gl+K1kdJtZ3H8grUnsJJeq4nbtsT7kW/nmUt90CkVrdOg90x
1AiM4hb7TQN0h4yd0YlP8uMVpviekAJ8jyQ1TWm4jxhMbdvDMBbq3FNcEfDVf5L3
HtfyV0p50Q5dNH1T2zuV83bMBZ9SlOYhZDJvr0XuEiBailjUzYZd7IzpC81Kc/W/
MqguSEtEyRGSJhvK9iJLmqytAxbkENp1oEw96LsF+iMsFhlBrbt5yEeQE5etDieA
FZ1rF8c5vTJ+BVfDfXnwwGzWJJVpZN72IrpuQGeOCXxzXlB/geUREp1Yv1eO4/bz
epz77J0BTvkE2SdEq/b2tV71ThzhxXxHoBwz2ga62tECWR203jkeoa+KOPmB7AIj
WIksKWHu1d3EpkWanGTFrIGftvut5tCDo5uL3bTIiBVB/LwkZHVPruV839aCvt/j
t/cw1LSrAzuGK09Y50UpXOd6u6fOndD2op+pboEUPk787+VBsQIhPRUE4K0GcINl
ayWS6y21D+Oz5/9m/Iq8MlfoygZ0gC0iQv61xGC0Bmzp6WlmnT/8CgH7LqKmNhHm
J+g11BfCxeIC72vJp7Gbs9Fvpg8wRSX96HHWSdahjI8IPQ806/G4bfmVtU1TUdTN
OCB4qzP+PThXoRfIKEh3hC9HgX19hIeaUqBDm/w97v30BWYXxNYnCUVxUOedyGC8
T3Q5x1xA7u1qIp/Mxppi/13Ul9dUUvQ/ZFsanMhEHt7NSqjAMRkkhagpyBp0q7Xq
ZUx9yAn/AHYuSKJretn7HWUqTJnpR0P7R3/UH/E21evO3yxmLbTlTdqugAJ64pne
AGu7/eSFA5wkCE1nQIcRuPHXH0wM6qyWdwBDZzrKSqxu8CxqyQ5Ympqtdpb4p9xU
YFqHuV3EuzHIpOc+bV8z6dTOx3PJLw+vZm7TBAljo1/xQqlgtzg4GD9+BYs+XeuR
vrWXXLGIYG9Ar7DpduSjUn/Hb0fI4N6xE9WXXEg7wFcbSYh0NR2DBcLgRBNokIuP
OkOgO2xT8o8DkUyDzdAQfiNiSBaLceoojx5gsstmkmy7K8SiH0CKksqbWsZUYxb7
zkocX4k1dimqNOKM0S+VpyRJycJ2JZ+J+y/Fu6r48f3m3V4dEoZ7Lkn91WvdyBDu
ks36sG3robmdTRkwx8iibA7pZ9c5KumC5hHxNUTu2+vhKERGt24Y+j7Crn7WqztL
qS1YvyPkeI3agIllKc2DRiJTh6PCXbkvHgpTXBEuhbL4+yb5Wxbg+KUiy8yNr69c
7WLY+7PUzREBA2Itn8ugCz1e3MmniAqQ37Cgm/dKwz4FWznAD6+y9cObDNCeDpvk
wgiBcHob2qXvu7qB5UxEf0J5A9SxDyoBtO7x0PnHtbMwvypFZ7kcrc66cDr9Uj9f
GFWhBVaS5jnlBRDyM8MGNwZV+bqzYxnTyhVoFkjk2XI6f5HTX8act/V3SaSlHM2x
AxPw5pkKC0+hHIxvfEJ4daboilp2H+O3nW3fd7SOL9BfftWopRP6JAifstcYaBAq
kCnIHbdSWTWmJfl1YgqqewHFm4EFhkcHFsoK+/hvWRooGIqd60R1WqVx6q+RkQBj
kdqLjrVlznhxeeOiNG2mcF8Hqgcg5cR3Kq+O49p+NHTpl3mPV1+YwibmqsiGTLYm
CQiANVU+wVilOOubtVv+Y1Ro79bZfphYWVsFvOcIk0OauCmuYaTWzTTUoWyCQmsd
1EXjYYm6ARX8F1P6eiCHObBy70gBqoeTMg1ZvaWQbkFkSskhjJsc621BfwiLSb2o
gWWtVl+vrERFUKE3U3NPPTBXE96UnuDdN3Cks/g5sk3nZfmJnyKPgkBYcCnMGPVo
M1ZZnIWbstTO6f4TihqaO6ikNrdohVCspWxwLzXBFswRorsVr4YEaxRtSeKrSLGj
gamxcMsYFOr0LPqHmIQBVuN6YdEd6C178V2A0n5K8nmk0X5HMxQtb8ezTuRs6ZoW
FzlH14WY5QLvamapG3MWk7HaD92Q7NPDgF2J1igGnu4nDt5SRSyl4O3xeZb01vDQ
fpdukfmbL7PERM5zSSi5lc3yF84QmFkJTt7XNYPj9qRYMyuUjtPuBUdVQJiYjmmb
H1L+9AYfm7ps+CDVCBqwSqGn7oaOXGgfcKQ4YFVF8pto2yT+zGTZtN9TZxPuQ7T0
l5DMwaGjrsv+p6ScCSV6ej2UUIxdfq5eApAmQ93SixiP1Voqz+Vygwp8N8j8fzDh
HPHLwJnOh55J99R4T03OBHalYrgqBVXOwynLfL/TUFR+HIB/FOr3b1aptVbe0p5K
ENlculw4WCF0dDu2SeMo5YxbHhNg2KDBiFdwfeAHdkWWG2jtRXRCG5kZfqrkmLzx
xcIkIDIt0CcvfKPsGvBA0FZKHmFWR5EEACIo3/WMrLSr3itMVcdkkkSY4Xz9xN/U
KFl1bz+Qqh88/ARcyLpwSVD2JM6y6kMrLjFivRvMHFbdLwYLZWjWTOJneZ5OY+jX
wamub5880uAHbSk+rXdUNPIFKBtUb7g91XvbC0ThfAaPn9iShur3R/ZXZ7IKDYjV
h3b8s7dVLRKS5oPXDBQ50ko2z/rmaD0qKvuuOwhcfQwmPtBtCz2t8BNBiUL4WoG+
AyGO9ig1Q+NYcy9obibsxNMZRtifl+5KdY/sYTS1UPnXDEA9nhAjefkmdY2u+zld
B/7wNs8Z6UbsAycNC2iLlQfz8nWF+tThzf2WRWRh5ds929LeF2iFg01A7+Fm8CvT
koW46x/OZ2LwfvGVQfFP1VVo3bwwGNNjQUBOSVYVqcdhJp8hvdPq05g2s8r6/boj
Vn0i3fdKOymq5OWUSl/1I4DublgI+CoqW7kvMG8SMvn3mg5z18nYqGJx88LHYFj6
rtkjdUHsS07a2g4wFN72U/nYDC5mAnSEfaYq+BH+UPC9nK/03NrjFWAGjnT08ckE
ZderG85kHbKw1kGc/ddut3tVWtD55wOhI8IMhu/vNw79DSpD21h+asXFR0p0QQXP
dLqvNTrFwbzPjXFgZASkaOxULGLOpIVMUWpYBsmxmwBiuu6QYqjm4xCGdx0cWkX0
+vPmUASpoSMnkcRe4s/FrDxCfEJldPfqg1BheceHwYF+BVEwxCgGC0VXqgKRwGXO
wk7DY44Jrb3zW/wEhS7wam6IJ7ly5vWWb4wyJrk3Znn9dIuerAFrmeMqQN7a54RL
94Rzu4xxJUumvw1VFpvyjtkSYTVzEPdwWaL9CbGUVC6qxUUtg3yIL1YxtAqTfs4Y
xbsZfr4Uc1h9SXC+3gqht8tpJs0lUzdJpcIxrPiLNf/HMzJeXpQfe/rT0Y5QxA1o
XO1CVB1hX6NrdtilcSlHZiMv1LrURzKvoqm5BWLeds2GDTFKhYyKYJD+KTs589mK
vLRgd4/iox4gMGxNijXAT3Ug2AO4UjUHQrmGT7cAnEQzvLDk5cFSiC+iUdbEV2y4
YVxnM+GKjSa0BN33KgCuTcWK9UkYDnEKuhKGn21rfE9aIqOcAKVavy1Tda8RTruF
NuWuPhM4jn1OCBlF1MuHVVhc5B/QrC/FGwZW8PdwwjNGj9XSiIGRNjh5QW6RTfze
WcHOCg/3lGNpRb5DqEPONtthCtdP3NoU61NoySpCuNphfsjVytAXzwF4t518do62
cHwsclmeSkBEdwcWzz1N3d3e3HcoAP4Kn1rSJtFUi466eevcUL3Be2LW/68Vt7Kg
P/TvlRruC5PhcTbN4aF5TFGCx1NdKUTk3XgEEKDj+KfdT98IxmJBVHcxrKyl/ofu
LFrPlyfJihv8iYV9GpIzljGysPfTEeWoFnWH9Y0R/U2JMTA9vIFxwNi8KLQAblX7
6Y+8c4gU6eOWTE+Lb8Du1uvmYfs0GIxtpwBVa+sfb3DaX5+beuWZKjEEo+1IYexs
CfXe+qPULX1YIuEvMIn5t0wDRU5/d5As8ACMmzPh9caQNh7i2agUYMejoj/FT1Yv
ZQSRVg97RrPxJUKwkvBGWDPOTExavtQjlSOD8qte1U5NMAj0+YuS3mI578jJPZQ6
Rmeb48gKSvyQ0a9VIqgvr193I7i72p9V1WaVVfBVFdtfB5w9f/LPI7dJHi8vP7LN
hXLrYMXqAJ81SmHH8H6eiitzhqaCLm7xhkyxU4ipOyYLtQHZH1o3g1/IL7umt3II
Z7jfWNIZyOJjDezLtpX0pTFLI814NlVFtRwdX1DJ7vYXJJ2UtivQ//tg5iC/QeB8
Mfxt6Fqkyq5y3l0HaO1dYihqWBzF2JGkpC59UqG6pnQHEh8Q0CNFU1Obx7RZZni8
xjyzoAZPo/jt5o9mq0+U9lySwjUtXaCVl2FgsH2guKChjqTUKWDIa+jxUOA3FXL2
2N9E3EM2ZC3P55zUNm1d5Jz3xmL1LekMeebsSTRcYKS4LgIvmCfZnGw4CnXrEK9z
9Am+0+W0paPVfIQzo3g9o93hwnyQNIJ1DsKSrxSNjFemxsFycRWluWwSAjdxTe9l
I0oeodvdGzPTxxeAR61nO2vS1bTdoNnF8JDO6DBDZsLNFFFe67fb7lnhtOpTwJaY
+SC2on8VTJoe74MqxKQh6vXrc924VC5T8p1Zw62rLsDhRB50jGjkBuDM0bAbSLHN
dRXbqpVsr/PhYUE2tE7C5jIXUnyl4aIA2MSxuCC4myys3v24OrgE0GNtN7srgD2f
qW3Bl/ytSUSviGBGrDOv5EXoBxRIVRwK4eRtH8nDjXyOoY3fi4z3P4N1aimN4HQ1
RV2Rcm73Y8E+X0+vES3JWLSSIshsLjF106ODgEDUiY8mFAEkRT4L56iOHTHBv0oR
d/LQ0cURidM1PO4IXWYF+931FpnM1DdWtz8N7f4Kz3gqK8+Hp+ubtFMlKH4VQvaY
mVrH+8WKmbe+owxj+DSwCOFfUxhH+0ihYXaBwmrDlu2jJvhkGiB8MPcfzuz4hCeN
cYLuZQoTu0Z3C2m9BG6iiUE3Sq1qoCy1Hv0yPcr60tL7BVKH1AH0sqvh1G+kQRHD
POwit0jgF4gwZdxRa37KhITaCe4N6dD5GwpAfPs9t9WFXQuM0fa7PMYMSUTM5GdJ
anTzgv+5lT+EIsLtq2BHUDq698VrpL70CfM+LjQZBMaWv+KElB+MXlRgvXG4q4jK
FcKUshYFymu1xPYgudECeuR9nOyCGokwdtsxS9BJGwz/MpuH+hdM4wTQkg95DTyw
9I+58n/yMYynKYgxfj9BSOBMo03h+4IHssK0WlLDSm/qhR99owb/F/eAFtvhzi57
LDlDTkAZxm/GCRH1SjWpFxlSznQ8mK6611zCG72+O/RQc5YYTcVn0VmkFdM69FEy
5rSVwESoYhhao9Sn+C92WWv+rkV+Bf1uDiqQc49DlyuT8FYfErJE9dWKdCN978or
Nm97oeGIi5CyVXMeBsvN5tONrAAeKyv4eSAK8sYB4Ie+YLAf52PUa6Etvxwa/gAT
/GJOa/15gISEHmt008+W9viS/CMZRVCy9KuR0+7/HMm/GwoEjAM97aJFbcwkWPmA
RR1N4lwks7RkIPgSrUGEbZmmuEfBetYwahG+RdOSRYQW9LX6S/hHm8Cx7glPNy3w
N29705lu7v7dCItopqvQrBRX6abiqCkFrS/sMl0bvRPpTddsaOyjs8dMKAsMDOWq
vQjmIaa1Ky4JOnJVpRxu1hwA8JK5/jrJlq8Rkcb2ViWnpHqW4C8iJAu/3sXop6EX
gE8wbUdQAXonNli5Fhm3AXCCDJVgNKDv3rhH33MLuB/bRdXUMZAR+XV/m/Y3QBiV
JL6aPmnu7N7phIQemEqnW9bFOfAEFVSFTzgXepPG1Se90AhKYwuMkbPIbK4WAxUW
dHGHWEUJNJSsmPML7swDPhhqd6PO2kq1ULQvBh/VRgmKp2JDoGRGM2endvdDEfwm
rCTTiTw1zpRms0QlVjXHfcdhDEj7mkA0KIVcsSBAUR4FkgmEoxMFUDVEId+e4zeb
l2pbEwKa2QNf37f4jpn+3bvAD/hQrhjcmq7Ff0aG/9YUvRMRn+MCF33S80xzOjZ6
BOa/8WgMfIGWr1PJ7eFGSJjxi3ml7a5lCe+FTyVf15yFdgkqkHRIARO+8QTPEkqG
AdlTeJFlx5uRiYlefCkNt/T22KtEYSqBTXxbIRnzqb83rySDrCVxb1VywQIvwkK2
mr38p+xaBiQKXQo5NpJ2awPdADapsXo7nJXDOE9xYq5P1ntscFGAUP/n5jx+Y6c4
UmT4IuvmMFyO9qONQLU2Z6drdA/yTyUQEUVvSSuGCX3KSazSMfQYj8De5tUmwAPf
axSTDFE23B6GXOLlg9UIVQ63cUhSy9LtyaS9Jt+atk366WN3PSR+bFRslUABvbpy
omADa8u6Af94SnRvC22Fih94+wGiByMplYzZYr0F9zyHog+8dwYgfc/tHnmlnr4W
HncVdhXcyF5oYDAhed4mkVTu7nt3xbEEBW6RRxe9AoWVyD+JzwFgqxMSUqiD4Asl
w5fevVTKwr8T983WqoAIzrwIL+P1iNxPovZLrQVYC9SyDJLs2mOn/tV3rWyJVAtd
C6ISpDBuXOTVmUbPLtZipvuZCxZrmc3yZ3bXKG/2RIqNsQDTZWdk9MbGyGLpf8tA
FfpJPIfdxRhNun/SWMw5j9+wW0gsekUAeFcDi7McPxO2t6sbw7H6Y5+WDB07T3uA
3D0t8z4yLA2gbXFyon52Ykhu7gw7ZJKs2I7xkJD+AwNK24iY6XnGw4hZMWttnATS
y5TP3ZcOeYY5wRKhfDwxgAjvYmrQQwAWI2jtvpnZeHzurtljc24jH9A3Vbky01rx
yjBK9ItkUrEcSIO7AIctvrXWOLUI+7v7n3uzOdAbsXHc4uEeZ6YHGvOOdi3OWGsk
lYY8s/y8hJ2cblO8x+sPt7xlvbPJVgS/itYhWukFpp/KpOkw4D4CvzXQmBpo4dDG
ZRYeGg1Z12BD4Pzfmi/CtCFCs2WiC/yZ7Ei7n9HY+aCF5cgGRCGzeK/rijEpbdhM
DLQ3ZFF0bWBfk2Oip1vF+pB7Oeu2v21afZ880keUMdSP8GlJM6iGxGvWwphuHFHI
gLub7DrKUgM69783KXGYy8gmTollUfs8aGg0k5qIeM03ihp2YmcCwn/GfFWhF9uR
/8XR8OOGuvy1B4vhl4UidEjetgghwNZCwWKkqYfB0rZ9nZTgGAR7VkslBsD+BNwF
E9qvjo63OPb6Lw/5fjVZt8+LbkW/IG5N775qCsGYGHaQPCitW9Jx7fybQd2sBycy
fyqEapOPGAsSPHH1v4op5+3PMvzOTUmxvwAkN+01keM7TZnW2WOmwfUjhRBJOtPa
xesoVp1CiVXCX6Kz0Tajh44vyX0MZT5jr8vxSbzs8COYOmf/KTsfEjoOjBEv14P4
QH83SmikXyh9A+aNQYKHbtsiKJB5hNKSCxe0mLv0clRMATh8RWWtLasWy9j7V2St
34Ed4KXmGY/jnXIbSTfZNI8cSn3DCWmR47Mdm9o6NVpRJ9eFMv5/epWNUf/3Fcww
dcuBcq717VbMlI+d4ekn7bO6dJfl4skMhDRs5j4VtKlNEKEvAp4YLNzLnPucPpGQ
X44JJUUNK7e6L2pvJXxh6LaTTS6UIPMlOZ8l3BfPfr8L4GAwk/oR9PThRT4C5J4Q
i1N3iXjgva7KRlXAzSViLIMzS5ZZQtjmx5pN2WHsBjQ4iqOunshA4y7AEGKpG3mH
Px8NcTIg4NqCbUELSSRLvHY0Udy6DDvU+HpPDBKmw0wMdcHB5/SLFWjFPjbX1I6a
SyiAZTa4teUsqtXSsbnKe748MOJ/4p367oEvzlEJYJQU7C60jZvQFwIBwCZPLXQY
npd01cgM3gCiRUwiGQY8qHUWtaM4weFbEs0eBHOmqpgS27q7lOoykvxMU4YyhC38
kPbEgOdTR3NZtNDqdUFeKmI1idQBHIgYUu6BvzcPXx21QtjtRooJzodWnWuclIvb
ZiiR9fbAx347HrMxhv7Oo9qbbNZXUQXVJi+4artEqBhtwdMiv3pcXkyYGjzZ9bq1
AR1RAiZ+b1x+vNC2I3g12qCBwbnze1mPx6FXSn5PZFdmuVkARPq+JNwMnGEKaU9U
tDHEktKjrj+t8GFpf29PnP+Vhy6At9ldJDeEWy082PTH0gJL77YgTtlJxbQ1tBPa
2Z1ZfgcnJwLrcR9eMVeA+Kjj8FVc5aKW5bH68SlgIdiAPBgzE8k0/ZADM8k4wL5M
4kCoSJ/fF/A/QTpl7qAvaC3HatA6GQfG4lBCgA0QzVUvfXK/r9GIc6dV0Ma8Vcic
VssgqwsRyGjwHSY2b/HDBPr9Sjas8q2pH/pMkigsDp5P3hVWEVNshlvUyeqHRpdq
3aR5HZ9zZdrBa/I9GHpHojkZqKHZmNeZQ3XroO6kRg2A8DrU/Yjvbu0SDx89oPuI
7nfELFVp5kcyTbLc6c4ywPEHxz5gFhxl6UipXj+MfxSYn4ofs4hgRBpzviPCIqjo
A6H0irLzH+tljPkMIU2t8WInfWvlgjX2/MUmThJopuymwT9sj70Wjx6T96dhz6V6
bDkyBjtUnoq0GjDuHiuipLBT1ZYLkc/SJYXnPFMQ/xNHI3dIqqNr8ag3ynZlK+bY
2O78LJzvrDPOiLL8mN612Yg1bq6Dyp9FlvJCCj1BOlqG7AoiUkBOlTJG+iLHzQIQ
hueRHhRgxggtiNj+zArFYCE4I89A6yMCWhC8Bv6kiLyhmALmGD46ZVu10V1JqWKj
+/RmZMMB8wa9Hrs1XiaPl72ahzof76q2nNRz+csvtHMJJB7S9/RhiNcD0GzDPldd
WN50wg4jiKXQy5e77rlXqixJS1zuYRurGuCqs+XiDr/n5hck1Cs04xXNaODAsE4e
sHNxwAsx7xhuh60x2QidEoWAY7LEEFC3T9xYUHFgCS5jYcOVIgZnp2DLWwyZo90G
s8gBq7K7YV29d8CHFmaTMEkl9gJidywqUg2TGGpt33CkGpbI+NJ5oldEPXmXJp0G
O1BoZgR8fUVCLn/nvd2+3qeqsanARvCtkax4aFNhiGzSq/EPQECETjM5JXV2LKgu
wpw6NCW3qr2v6FUi4+X+hhN49vWX3a1YFfaneKrXevavNOfNIa6Dk5FW2hiHQqvk
jZjiOAUFXOPV6mH87K22tyKlbXXtE+8dwLTjNhZoIC1YwZs/FuXYt/I/JCKdG3CB
P1ouFBr9Bfu+Ww2rw9NqDTOQZp+o0jXocjDcHbvzfdcPnRDClFe61hQgtMvN5HbZ
pcoB7rfc/xaoWJHK7NqlEnWcCJk9Y5kF6zyFGcmnFq7iMp61Vfm3jxRPXo3xOzv8
TM2Z/xoqHhBuIQL5cXKv7qre3AUKSLw5WCJLrNij8hoLL06Am0J/tZEYM/5aTuS1
fWNTiyu6GO3MmTjvjVPnWoMeJQukzqfMI3p9NM9m7PT2nPQyrRUgjMUYq5Of7xvQ
47YmS0RioLcG/ME/hYjNoRFuaCk1MVuK0R7phHBmx8cHoBthWBlWZDaV6O2Nq/iA
yAhBZwdF+i+YljONHygkGC7JAsitoLobfDTc9ANESKc1taTLibz4osChYiv80+Zt
lLCr7JJlLEQ/GrN/sAzbHTrYuSnrZQScJOG3o9hnY2o0cUkISvrKiMG+H9Mgo6Rd
KOZeSj1+Obv2S2S6sj1MUELI0Naw+A7gP7pcFrRUKPs59HZF/2TpMTwEgQATSjHW
50Sd+bCrM4u/5fQ6ur6sVPEWtcfM4A4j37pxayPWP87lGq/aZgBBmUCSyN5k6YEt
B+W1G/Ia3otRc1AMHsefpmMuWa6q1OzZ0mRXRKJXTixGFwGCifwuQGEwTydvgze0
wP/7jVV3ARTk8p9yKyxZdXMybJNNNSMDkPxKjKqovfKAhF0NSUz2nJ5WMvX2qib+
ckMGBVXvasEURVJrBoUToA/I62cGiSymmQGFk6HAV/ZA7snf0JVAZ9XF2I+kd87I
3XQ9qb8iCucHaR3cau4G7B2mUnoJPR1/tQsL8Pq8BZ7sFOPQzalYSedHEwKfpUvj
7rxA8ITMJmoaBDY7Uez7Zt5gHsNu5DcYLwXSBMHikIXAbQYiLn/0bGw0KhE5J9up
XnPvYYjU5NTA7H5oMDLDauD+kyEeQ9kfeQAXyJBNORjmbc537pljCSc21+nG5SL+
1ogNDQ7YdDXXw3gmwo5Flxpf0pFx7KiKFyPp9+5evUSSib/dW45vw88wzIgPqy7W
M348Io4t3kiFLsgpQVV0n2nxjzYnk7RnEYqi1S7gJpGe4+59XgqG3Sg6D0o5ZwrY
FQeDtre9fWyq8DrBy5w2ZlD9b+lKGk8Thix0i7ueX0ONJGvfyGVbIO6YZ1qU9vjW
eqEYegfaOWd/sb5dyX/q2Q62c+SHBPK3YoahtRJ02ExHjJkTsG7IDo0JSxjyULtp
9tCsrFOgiq4q4R4Zc1GcIyUwsB2o6tMXMpmUJvTH2ELKx6XFFinhlf1ET4Zrf+Xk
ySK5/Sg1ZN7fwb42usG6aVG4YW7IN60KYhyVTPGCvB9PaRdtwqHEuLD2UPfdLLza
H1o73YJnjOLz2cgjEfGF3zVhQmIL4VTLffouTADebF60tvkDMwa+t+u+fV74fZKd
PtVbP9UB1XU89Dw6xes0Tj6ZqDxAxnGjWmeo5Hh7SQi1laiKWFz7S9BOtH+Wf4Wu
HgzFiEs/qTHYIJ1z4byNRE7uT9z/t7oLgIh+goF8d4j4DBqfRTxVYjep+cH0rkwp
cFJxUR84wb+43ha9EAfqBEEp27E6NZIrmEXBVpHeTmZAyJ07pf5cmoJJXQWs6fjg
VILpzxDrGCmGCcGf/B2MaXB8+QHZSQS9MOyx00rHWT+hVsjm06IuWeOF3Y7IWpBL
waLc3nhe9ick1p43dydCVcju8Hel1VerOiHcf4Z3LcvKo3m9YnGOwthOEBDbX/y5
Z7QYK+SPN+otc92Vxa/uVBCxBeqsfXVqYlWO5UO+27exVzhJpywNu9AjaA3bm7xW
uG39FKI9/X92z+IC0xN3OVyh5IuIzLYFQvFRFxtJaH0KumABkJR3LlUyfsKYn3gc
jgJwH+0bvNvH3TuQ2geFO0aeICMgnWPVjDBFsfVILBL6H8sZDAYB/HQPUWuMjl1S
XfVVvvCIzs+0cDYijEciu26OqQoG8h0W3u0GeNvkfGXrj6WkRj8yeArOcOzWGFon
C5aQ/BjrQQgo6Y/gxRSTLTUVmcMwo84BP9crkBpMANMNoFR5TWo1DtIcJFB2GTQs
4PgODf8jJ1NDRugj9lMF9LKs+SY+cK/IR4uDgZtTpNCRNwVb5rO3b+dw28ZH05KE
NpRpa8tzvx5OGrx8qeRj3avGuGjAaKazwVayERjuAMdH3dqFiFI/Fiyw1Fjb0u3+
S62b5GreKVX1yvBqsFCSalPmKeKZVQ+f+r5s6E10RTSeZB5qnvm83VY56NENpoQ2
gkjiCYiLj8SvxNDuC4brJ+m1B7VQZPcUSSKM9cgGaDhQDVagYzGZqF3TVLJS0Ktb
y1Aiz70NLuoHJXPq494yaR9rUlqZZxuYGQhx8JYg3TDye+BUAnlb2t91Sg5EcF+W
M0hfPGg8Pl40+uhijVZ6h+K58lhix58NmjOa27WUULy9DLg5LJPoUtf8UkmY5/eT
d6tKRqCpfuJ5LgjY7y3SvOK22JIO9kBDr//MBgkcX5uoCLtrnOHXjn22QLaQ+vMu
PJKGQkKOcoQp5i+lYMOFLETyta/Kq3QKPthPqvX6cdSVuJQFvK9EUzUQ3QG73lUc
xcq/P6wHHpv6RhA0FebKT1WEsonKXscHELmeqZCgCxKc0Rdk8iCgENxNm8Isd7rF
O+IP8qYEzl9vBg0MUaIziMuMWVyVvXRqvLAay6gthJXuLMDKxrlagh3dI1cNviAZ
MtNwCRAssXRLbeoEMZODFCaV/F489xu7CEqIcqsHvf58p3dW35MN4I4tT5bQwITU
wdYnZeMAYZyqWQXhCBruszSOr4yJMQoUnw1/8rURvqsKY2TIxrD7+Rtjj91lTqmU
buxOSgcFDG7K/Z6AMjzNbdDUbNeZ3YkqosB292IRTFqAEbQNfY9PO5fugg66DD+6
tQ6AGBC4hKzUL8aiS9Tbf6LFkhV9yvHx9ML9LakvpSQ1V/QGZocowRyOiQQVXMs3
sV/FeDK/o9WCWgVU12zk+iHNL1PI9jU9hv+A5nCBhk2vZCLs67kuMtAeysRyfpsJ
AqFcfCizDrU2Tk+gevLLIGFZ7LFqIeZgfcsPIrsIRSRMMAdQDGjkfCXi+8rzT5lG
3RfeuUCBx6wWuQJe4o+PssDIToW5PDiZsBWP5cq6AQFQ4mZoG6rJSa9i4nDK5zwM
r07p7tuV25IEih57WWqvolqSe2JrPKYC190s3dhwTPaIULJqnTZRyY2GqTvfCQZK
XjXcsC3rM2aoyQcF/uxk9VtZ3l8IxCZYJjkfrLdnutslOJG38eGsFLm8yN+DNKun
KwkqWDawErcYIDkdcjEY3vaXe1yOvb3oKb1Rir+GIXMECsJMYtHG3yKr2aN6SmSV
bD8Bu+/1NPYlbmp8AeMkGO05hChl/lzMrl0qLr5AAIcmbKpkI5+Ock2Uv1HgHr2P
6tqcnQ7CFUgnfvA8D/hgipE1PDYvXIR7ezVozOKmAbyeu56MHcT5qt3VGblq8Etj
m2t8SyfRWY3n9WcMPvpL/1kRju/8o1P1YrO+R/qX6zgVQ3Czsm3JRmD+MFNVAkAr
0xUVxABXYJaE4IsCur3i6y3yqq71FQT9LTyDIF6jbtIhSFaRwJ4PbxVd0cMHJ1LC
MwjgydXjPpjR8Z+22H+f+/P8quIfwZhb8N2Fpo8vyrsznLDKq62bguuW/G30kKKh
6zhg0apZFUNYs+I/abo9EKseMRv52j9ahy/i4hAqTclJHMNnttDPBZaldbG1vyuO
o5BufOenWAt0qchSRYa88aokYFOpdsGK6ppnTZe/qzd6ZdbUcO4Fm9lfG3blCOHM
AgucA+p0CZ+BogRq+Ieb8AZPSncd2Igs1SQd9uw57n7512tqMYKg7fNIKdxPVoez
el3WmI0XzU0TMV9NHxXyiZRtEraS+zBxhXWCbCqkwRaOucywESNypi9Tn3dlVO3/
yOgnefjL+QCf0qXcxICoRWU/6N1978NqfjYTZ3uwyDguEoaiEh/9vEMCjXGsaV3l
HJXkWRMisV3vPM9B2U7Cgy2fpNvMGReZVu9JBiucvILtGRVjrTL5xpiiNX2S1UAv
6BX0x0l2HBvL9IBvWThh4rODlTbEQudFUMPoJIS90dxf8LJC34sV+P0vNdWPEAvy
OEq3fXe0wbUTTBNCH6XR1ewoCKNKqrmDPsu7/S9qH5vjvVdbFpBkH6Brq2k4FGp5
oEdURSPJ6GmwEb4flzr6Zqzy/wYIdZ7kJtLjdD8W4Kc83McmDu9opOcsEZVtTUdQ
cK3fwmDIIDwAxe9rv73AIlHYht31j4dFPBTE0z3w0FFJjOakmRKFvc16N2yKUl5B
UF6cKmsYwWjhSI5ifk2+gfE/bXadwlaUDCrbpa7pIq0Hfj3144Edo7U9O8IPwrkb
EJ7S60jgxYodfFeA3wQRFdX26RKPRHUlvzi2bpAkUnJviG0bLrAthkx94aMvo4H2
jT+H26vOQFpwNKJigTbFHftDUjp7mRoQTMQlqamB2RSdb8ip4JSOS/qKBy9gXvma
4H9285zJseTWkkkiMl1SFqTBoOK7fdMn+Yja8ATg25UA/K3lq/Rwc5/gGf44bqSs
MQpkUDi2Lol3p+LrLvIyTuIXre3ga5U/Hja4dF51xtznoNePUbA1lqKEx9yI0tVm
CsUqMV6fIwjUrvpZ1MZCop3l4eqX45/YUSPL1mzj2ShT6o5T7YgYNcuH+fpPYdG9
MSMzz25cLUOtUHkdcD44zl7xwL9WnMYIJYyFpc6Ve90/YtTBKqvwU2fuhXKkzkCD
fO2/lurwlRG1q3cBBvgIXv7AsVRHDdceE4S6jxzlw7dZzPyAiFMeNdnxVgTgyUj+
I/0Jk21p9bHZjakER0ilJtg0N2lsoMae8V64dLFHJoETFoDQho95rfTQCu9Ofsml
cwNRCF3cJuSnu+crtN3l0n2dtKfRkd8eFt4PVPj10TwsQgXFzS02A3tLqEahVYUk
wBMBerHgXjM6jxfBlcQa5KEjCfTrQz0TEh0tMjIaXBNlEGmA1sPrxHNP6xUYGuhL
0Nm0WmUgvcfA5NYkV0gVT7/w6sawFLMoJZJJoDtt6RT5VW7ST7hZEPkTwOf1FefC
9zBsUZlppC+m/QVRBkYolBdhdeBWEhO3brPqNVy5te0fmWN7ftavYQv/A5z2Oppo
6CHoFZLLJontfhoA9JRJl6bKTx+VsQr/69PvOdeQe/JqSt3pmVUKqvwaxQIw0BuP
5Mu+d6PA6PlFjmS1c3AohFPg5mUmI3pWBdRVPeZZa6tjJycxhFG+4PhR8linn6dC
H1dwa1dSQrSDkoyzKUdev2DyIVuNQzlpyHc1qDVKshrI3woLxM3QvYQJcXWqrFvV
EtnQJBYbMMQbGI2RDFf3hMGEh2t0+tpl264PRe76+hftjwHFm++eJj+ic0KdarYE
Nt9sRvO12lSrEli5CKBLUmTAoHrVY9dTdQwYmTZOZU0B3FLgRYU2J7JDXI5K1L/U
bgCDmR8epARE6Izs6EbfuM1wHIPjJ5UDW8V2m0D1ncPWOmiagvTy3Ea4HkLsfPkM
VVQxqq3Zuy3lXHsUrsGBNqAh/CuI89XlN9fNhhu6KE70ifK2wA/2+TzrOHGNx7j4
7yK7VwoKvuUb+lX4E0+p56TY89vJhUoXhcxIa1mSAoPQXkE5JnQva6QQfx39YzsM
79xTAAThyZZrfycjlWoVQhP4RQehCWuIAKXTlA5j8HIeNZdAyzMYV2hwTjewG9fy
DHgU9p6rV/o2pXmbeENnfmESDwqQjgoB+8lGA6PlRj2goLdhv9aTUZXZF1dwIzMd
Ia2OHWcJugyLYWo7KFA/R2JQAc5tVuN76tloB6zzaSeDUyHlTA8bFp9lGaP260Me
d3CqiSjCC72CsoCKb2E0jlc/5bIPQGvBpfsY3q7p1R7n7NJZdg6Rr2EtoFLoXgNl
sa+GalC+5Qx6AiUgIrxUPf2B0g/XMhjbgUhzQRVcEPcFUQn8UVKa338PtKlSNSis
pN9/kUwJ5rOTGzR8h80ObDFFmH7nBnSDsHQ1qqb+c2zDM8BPaJoYqay0fZ3u3f6d
XvG/PRreBIY0EphpxRAL6vQpYskDkE35zyj0LDT2tac7f5wSAsUIWiToDkyMa30y
cLE/dDD55zYCpia5LsdI6dGtgPodWKvIJ6u183uUwk+XE/haC2w7BVmoKSTzfJ0L
vdw97KhaCzAA0JDVLHw1zDbIQ1FB9Z+2fvbvgl8sdK7K5jp7KAOQpmUqyrkxXcGC
EwpfQfogE1BPCLTgcgWugWkiwFUkH/vvdx3QsUuiuFlhpjPlXgGw5SRRM5jy4e0X
UJhK+789E/lyQlyKxOS2pazOtfu/ErCm+KnsdJMonVCdCs4vA4XP/D2M35P3FNo4
281a9pDX8Ayf/YCLk2KzLOqZICL9k0vuVfrGIIg4Yc+62v4y7fDw+nCizF+/ny1w
GNlV3+0eM9eplKqvyqBJMif2zhj8mz6X/1ZvBLQMM3LW9rKLACygc04csCRNGnVT
mbsTldTNuyuVepSyHqW999oSpCuVzjuIV/ISfoOj52k4Vb8ytgpHHdiKdGdYEclW
rPK1lUaq4WoBH/H77JUub0ua1eTSyUCrTBgSRUXhRqEcVQomjutciPRgsh2TQmC1
2mR+Qy9G5aILYT9qyuyBRRustQ7UbBFfRxqwvW3QEs+cMw437Fw5cIKggGvnfCTA
qwZNSwb8NLL3gycgYFof7/LqhgZQT8i9tjT/ECVa/C2qE4oPL6vE0lrPS7+38pGt
V+A4qKjlochcPudd7+mmQz/UC6I5ZjE0m2/RzyxXmCj4bM+F9HU/BcpEUwxi9EAT
4XPHjTw0DD2GSQZTeybkQ/XUgJowo2OkxpIri3GlfnaWAic9M5HEccTCYg9REioS
nQKA/CvTKvNC4hvz2xJDjPRKaVRYzNoDeWNiRsVPDcKlG+rpYREz42tqmaDto3L7
Gxa7wCkk6hh57pa+VOLGMNqEO1w+tghJRtJ3oyQMEciAUllLCYRfZotHk3auq8t5
4WHZ1U6pW6LxWqPb9Xb03WUYPGgLqZ9P5YOJq+BBnIYVgnck5khGCwf6itEzJ7AF
xNWxSyROX8+vWse+2L4utjMx85PxQosGiZkX9oeUnud0xaph3nQ+L0mrUQxhTHyt
0R9JPOFYpRtBRikfhrA586JnY4ksWx4K6xOOAWQIPK3wKhQ+jPQT+IThq/RMkn8K
VZtmN2ao/puEU3n0aiP8JM9KNHV1WCvkleRuYi2IJTcKksRzutieoVUSl1tPtmik
gE4Zol6iH8gbMFolZuRv4RmoJNC7cCHuXwqv7Lbj/aIQ/tw7nKR6bVkFKpg7UMDI
t7E6xgCwM1EF4ZTF1V/jgXZcrwsEGLrQITnQCZ3XP6aSesRcQ7V2PcDT6Ayc78yx
A4FOWNGGb4Q9PQ8hVRjo/7Ixhs5HmgNVI2cRfXK8XeNjBRMVkkoawVsV+o64/lNP
6MQRsunuEOq74lD9TaMBA2kv6yXii4a882UvRWbsm9W2yHHwMifvdu8EhZwjodHS
rdYDhG7PeCQ/hnIuofPJg6/4yaOlbeN1DZEb6MS7M+eKAjz51f9UavzhnM4zpIk9
6zAY5PKxCbe9b1ilCCbeWpeRMu4OZ7njhFbDG2l3SQi9mxD9cWT9ZD3m88Rllw01
99O1mMSEqogPL1cw/54NmQRkBhLBdEtF+tzvggGCWTkXTU/ZHz9WZQthuqyCMCIV
8HgGDw5wFCIEDXN7PdLMJZWDCLA4dWrTAYlsNdUTcNb6ex2GIGUPrOISU5XC4T2B
JBXzqTz1rrt3A7Ctsk+ZvkYVDTMXTufhq6eC2FIcIp7hab05pIXhCYdv0GiXkPHC
ubaSjNMIB5huO9uvFTd7EQSE+QngA9rn6D07dV1TZfV3p0lplFysnuAV57y1iJZV
+E5wVROIlk1DTmC8BWDZNgdr48uBoCiBj7Xb+1LiVV/OyUrO9V+RyJAGHtnMc8m2
qkqDq2EgUj5H5U5Q37AFDoiM9bXY5zZHt8OzjiaRpYc1LQLDbyVCTiefv5+LH30Z
495zjOstILmpREp4ONjmEOlgb14fZu1xKnlpFqwbeyHauNQbQSf/lZ/SnWELAq8j
d71RldTfsTReceWtxX5QebwVrofFEshhnsX0cbpmKBCmtTJLyoXX0AuVMbtZWmIT
g2/sP4ND1vunn2gnrSSwwpDCGOJUgWeDpYW6nnK3vWQFJd16c6bPaJiMX0z8zyth
psLImekFZpxTp++kSnOB640s2rP3mGuAD8kce98RHrqNLYeQewllzRq1XmzVAm0t
G+HJRRYfDIbMl7+6CiP7p7nyGW8e9uWkoZ89YE+9H0t86d2n3NUykv6FGQXW3K2K
hIPLdSI21WkiYu3VC3B2Nk8lYsHIyt89IdnbHJPS5PXjG/YSd7s8hzryFRby9EYF
GGER+SN8fVZoUDWQaIUJ0Sigh3PrupqgLRQVhdHAq1XZnAjSxUmDsvy3xrQdzG9D
4isojjCrGZYstOUWRAa/CVI1xqFdbAqgMgVvJw8dYpbi2BT4MqwwgUhZqTsxYVeR
/EEMLXevjx18LAJ9Rgn8fsS+PQMM+NglCYb3VlsVuSy5RS1gJ9+vFHBUob7jQl8q
9KKSmWamfLO4UiKgMWbPPrEX1+NMiK83VVU6oa/Tya30eq2as25wwir/nvtR7V9I
wdJA5ryCA8Xk6KEvmI78M29hdK3BVuwO0Qa4RpZwjGbtNqKZ+kUjDEv2/BIHm2B5
R1JIyg9XAHdX3gGoVewj4ZetcxARLTlah2DYYje8cSmoMydlW6emCioHpXLeLmaj
ApwU716iABZwsLy4Edx6n2jC0iY9TLDzZ9x3dUnK+1/3JsOj4bxdzwTt7du4vm/J
fLdPtBURh9QLY+Zrjl6cOheJCABpfCANW429rvLvtqUzTDw7O6P1Al/v1vCUQcI1
spNOmM7rjLQxlMyx1MtmCm+J0NgxmOKNp2+p7mrb0IMLZmpbhmKD31sXDxa11vmO
P+ZqyyhAEUFq05cvRWK8TptfmhxruFXnN1AXwTq/hbsuoDr0LszZIAnQPpUorfsS
15qAj5y17wnC8O1sPg3p7Fex7K997XCxgIqg/s8rNtoZNPyP5lVfpzO48mDCrw95
bVoGDsXNMDAGDYjWqWg19Cyqs1dH3pm8aQQxJFgUNVWsV35WYi54HHMYbNueM2kE
+aUVW77peuFAHR4Ky+CzbkOjH8KpYDghZ7kwOF+uI8KGc0IyseQsHm6s6aD0li+S
GK4GMNgzH6ZvKF+OEVrpX5uD/iQ8m3YqfZ1VV7oRKBsPi2laXPUL4YoSNQBMVJ/E
qcciOHdkeAFscVKjZCuNitmqYxgegbjFwbS+s5C2vuLAwh7B7iyl6J796ncUBsgu
GE5hEMw/GrNmQBSPj9Ank8NhHmDc2LleY0YtY4XQ5wPLl2RvpY8IPB81D08/Z2Ea
HoInNEGNtN9Q1pR7uSWkeHgdP9Ji61KCS+W0Pc3yOmpaNGqKsTKabQc/B3LenqCO
RQwJfWRXRHCRa12ao2WZlHMgld4sfx4x7OTYR4GjU1QPws7oGkgxwfEt3FqSjDVU
CTWfwwfvvAQ+Ku60Z2TADSyFHd2kXfCNwTOyHzOEEPH/g1XeNZDYS3zBq9OoU87h
HrFXNUytpWEhLIgHzozskx0IUhtSljiO95ZsdSZgScWe+Mbh2I5y+x1mVYVhRx2m
O5jrPzq316XInja/B5TVqJp2JcG+uMAtnpUlYmXPstKxllbkAbiTfYrbFGnR9fsv
9UKZjNruBrtijYF7DITIDejxO/RyyFsA426+Fzye/M/GnUV8jpPz0S63oxxIPp2s
1tZIlrU/O6DEkeTCbxb1EbGqf33qhSZNB0UCPZpFZ68yUg9Tn2/AVmun2RTKdfOO
f3KufhNr3cOew8u/I7QiNADo7ZhkSjDBJ/vJU2p7rhpC0+IUsWVU+g2mtW0yqSJq
wwGsPx0CaHHu6LJl+T7wNDL5mwaLhuV4JTjrhb3w5n1n0b9fJUrfK3D8yNgVNq/5
Dosjzqg5EytrmURAfI0ggX7btGxfuiERBh1jMm/rRuh+PzzW5k2vqaiNHoUflXv8
nkGSN00E3mtjGez91VDzdMvhGq4SaGCNY3vW0Hs+wO9wJmBBNJ7nNWnp37PrQL+L
1Mv8OB5X4Uqgc/PEp0YMZS3CNtnO6BkdEYuMDj1eUeNHt/gLjIDfQomn9/CI9Eem
CEQfbpouBUucPucUA7yIs9aRtsiOsAI9RtfJ4/UrzpbA08y2tRETq9ds31GILT7H
dc3SylO6Bp+KlX4ATBqlk7BsVIp9ZCwDzOHLGp+4mO6W1g13Zsgv3ZANrfsCRSUT
zDjzXw2x0sVJMn63gCzO9Wjtp6XShY5L/1QjXBcaBqwS5hSG5ml6W0yFQSiCUXr/
oc1QUvq2Huf+U7iKEv6hM1HFbyoTJuRsEAjCi9MqIhOZQjPQGJ1rINeDeCUQtLtQ
/Tx5GPxh35z40xWWOBs7NZef8xYycLdZktNS+JhbEUyRuF7Cd+fRPRQ6V2kmLvO/
IcV8MgIuvEg1/PJ/KhYCVs+4DY+PCawjASU7KBpk8SDPk7X6yW1F4xPpmQOr1aeZ
VNDc0/1TZHkG860l+xujrMouHFeZtNY6nEo3o4DlQNSTqOBN2XwN0mf+etHUnT2l
XTiS9KPZsVauVytPppYZASZqau8jHrtUvESleCdkP9T8tdb2UvfrXFc6J9SSgBF/
Yv+lmundOoiySosc4o25hlB5rYe4oMCsV7kYXHlJgNG5HRfic1xUul8e1B63gN3p
KrSYPMsLPpU0U/Ukcy6tZkrIgCvOOWlT1Iyd292MN8PGUfZodri1DId8krAHYcLY
NL0GdujaMRGCTcGWC4ImXuoMnA9H/jj/FQfhGv+1uUACiv3Q0wxGL9Omf+6tEHa+
ymlOSJuut8BndPreK/O3jf7nn+YhiHmsbEmkBR76kp/xOtAauSq7bVhneUE2Hqvs
VxL43CUX3OfFacFrp8LBZRNn0ie21iA9hMxcQemNcTa61UkKcbAIrr3QlClChFF/
fzIfz2DxU6w1JQp1iD6p09sfMlMCDlr85ZPWzB47UBPWnucAhXigswUAyGj7l047
q91AUhRqPYmLrozqP3Ed1kGIlmJjPn0D3FliQU41HAn5Pbro2yP86dxpL3+Y8XMT
dnQ1i2Vju0xz7M63MbK/w7MzzBTPwpCGhTwOhpTM/clcF8tzSw2Ulz3VAKyeDFLk
rQGYzeiv5pyaL9jTJpWRLxEwRhmtpcK3u7qN3oMLWmU+JuDIRf64HDtYiAvV+oQw
hbe8zwo1KKTljsjNRpWY2+9VOckJ+m/MKrXgFV27rWbbPYauJ6MW1vGElfH9m5q+
B3cWmQW3nHQNkYZUKjiwe+Ez1FFqG4x5S+IfAlQUDpFWO3BjuginCbMs8ysTtwxZ
zmRhkuD8OUqy6jMAJHHKY0e4TT4pJ7pQrvidLDYlhfnoX+EQ+JQh6hBR8g4LUVyX
58cBXaoBccd5VmQNB6nDmZfp0gWRrIlnr3hAUyKo4H53CV8OErweu6b/wHjM2kHN
+SOIfV/RY+aDHOZODgRpLRk0o4B32TTTrrvNKopkf+g0F/EbcJ7VqiWh0lutJO7R
bX0WZy0LYERV611Wa9DUdV7nXBZsnG9SwsBAyDPiJ/MnYABs0UxLJkR4NrfbCmY9
zZsXw5pKRRLmBQTmx7YaGGawillCewcfJ0xUX6OnCYHMxNGJqABGWR+dl39CO3po
d1OQi49d5F8oFFqqHmZT/NuMxjnfG+nLWuxgZOwik0hZ3k8fhq/kbxYguksUuWut
IjLrXuBwREXhWqB+dSNbVev5jVAzC2TpOUYVC3nEWwDOJ+jppXwoIl0SPsdZaBiL
nLQAO5MKxTyXF11KtDEdP9cfX5snlCyBeWRkEgD8wVUJx/p4/IK7jaHs8jm/IGza
p27QyMop0m/2D7LbMw1hyPwYqK1A2REYqLSyOmOvGWifR9uzRKZieqzbKOmO2CT0
rwoyBeWnUUIVC7GkWvjKsy/8LmcwooxevM3IvAlxs5sMxMPMjb38xkm//pEtqh4p
8MC18P4xgcc6uMQampoPIZ5j8bMU2WYvUAvGj5C9DXYkhi7zdb32MjozOLiI0zcZ
LgR6yJJW/q68kQEfJCnA8ahrbYcdx/Kz3Qa1DlMN1vwX23FCEb/Tyb14FP9hYAq2
YoHcRXyvqXi2WVJSKIkpp3cjwRgI0w1e9VRJ8APUqRFWyyI24vsc40itFoiEpnEO
O2HZ3SQSHD5sux4P+rm2P9zRe/9ObiBDXRQ3GdL+uzC/uoRY/Xyz5Ned9wrYVY+b
xL0Ld5Q9Yj9g9ZQXSMB43IPsh2LHpiCGli2npENCtkutGi0SVpob3tQCCzMcn3Jt
PYOwOTaRn2v0/SE9mUAw88uB/ogfVYjR6+/ouFWXjKQ5YmygaJnaFz7l5wIXB3QL
wJ/OAnW+k/lqUVXClV7AXVneTRmZhJEVgPcBOC02JST5d0fHKjOfCsG95/uaNdLZ
supy0axO8/W2n9F/TG/bzwW4i/PSg17tRSASlrPFfnh0nOt2+enaIqyCuDtlFYTq
ThAL2LmnfpVQXaKbQ0V6+aamiokfe8TcCzyss6tHGX2gK180zwZERScCSi0eIM0q
itdVTUXbSfeJfNIDRe0OsWC76a3P+b1WyWxLFLthiqmafOFt4x9K7lp865ypjozo
7B174LrhLunz+K/XxN4Jf2T00YsR05rwoOKQ/rw8ADPurIB48xK3Xtrmn66iBF8y
E0J9AXJBcRC7BVCeojafCI6KgPBwTqo+06TP54vI6HlXu1l3zTc6VeoyXfVYBex/
xte5nxcEbIwIwMtCdZvwEhlX8x3WEcSSDjB7LzB2u8GDbUkeqGtVgFCkJnCh6lKV
qKiF24ccTMctStbZpkMw6czUEbKJIS7K9py8dnwQ6N87xYPGjiONSgpeLyPFByQ4
Il4cZnmPA4boaneMHnMWFebpuUB7hE+RGRb3vWjifnpQua3JnoSBrAMBLSeHIb7I
z9Q/BZ4u8Xj9TOKhri5ygGB6/DyP6A/Lajdy31f690Xo0MeWioRvCEWyJ+l6pzB0
lgH/uUJpInogp9kGYM+IoD3WUCXQGYWM8D7hs/68aW8UqiIcDgDV5LzbreekL961
qi+4P4ozw9hWWceLEoYjcjm2LPNZkrjz/qVf5LrHciEWgKw3R4RzwaH0bPafa66L
o+IkS29Ik9/STlKdul9dkiHJgMcoGZS0SO3xitfEkLDfRCf6JVioqwl0pPU3SVZd
45P4YGE/jUvodlLQLNYM+MRFrX2qMWOrWw7whRgPu499VX3oQanZlPcqcf/EbyUo
TrWp3wzHMbiF8132WjIRuFeFi3+tGfnLmAoALlGoTPA9fRdplZ5bBdzX6N7od27Z
/acXXiHUCpNGUwPBegEeE+Pr7MUhfMQVlj5y+SKQZOOio223VShf3a74oRt7btOy
BbHJ7Y7SqlfXIRNUWgwbGWHHqikigPHqjRFUnfRE/So+SeJBcqYz7CkOKo0txfNT
zogVIvZAlfUcOPmBK1dvJDi/M1bwngL85Odr/Wyc+S+8ENNhevUDsSBG7wH0nFpf
d3qfLJcNHeOFqkw2By66wjZtiNFbSjp2s3bSLIYBW4XaA4buIMaqPB2NBrZa/Ksv
3Z4xyETce7g+sGp1706knj/57Z+YWkh5khwN+KHz18cfLhjuDvkVThvyhpWcNyRD
QR8sdPW33oXqxU0Qy7L1avBMZm2FHvuNOmQTk0PF3xK8f5xx2BaVv3jXRa2PDFXm
mUOy+aQvCVL3p/N+UIUeimq6Llt3SQl0V6yLpLm6EdB0P4vqxybPdZDHvbkHI6yp
PFyECAvMqv4Nshstm98N35WRKFczwyCr7qTEIRx+ZYoX3Ie+pbgCpd5hChY7Z7Vp
XnAZ6Deyi0DEoImYnhshZ2hnrWmKGMYtUimNIYoA7oWjHGmwF5IU+9B1qf8Xr8UT
YCCmZ8ZVT8+hOnnXbzmA8LOCUPTg6+Q7a4JKuEOzWKTWFJCUukm+2Kzxik8SSbdZ
1Z1BKjWjI4JeTz8lA14FKVbsdxe17dJ5EN9b4cSo0/gPEA2hmLtBiAGszrcLEKAE
tWXWRhY6SKWfE3k2RQQz1YXhspi1SmMEJPm6a9OE/T4ecide+ZtBW4/WkVRrKLgF
6wdB0KqwJUz6MfIiDFVIh3TLD8s2YjtvFKAvoLpNm9BbbVEd08XIDm8Ze7p/fzcW
ZGPDgcpobbjBN9EOGJv3HayoS0nfzblo1jWxp9XGo3g5VFNAoxrC/0Bdx7aJrg+V
URxVP/QGAVrVIXtX1fPyy5dFs/CFki89JfoDynAKXPniz79xHakqZd7C2spMq1Q5
cVTp93dXoZeRe4GjiVSyTDjUPr/Dlmup1oxsxRDznk6fgT+h81W02Nxh7dBeQD6T
LHO486hh5PZOx6JCHwi0MJS0/P1eE0FAGpFR62IWi/RltiPxezqWxg4K8rHA1b0x
Ym9cTmat4T/sEyVYQd9N4xvB+T64UfcBwMyZDqu4SymXEMCfo/Q5NpWCcpdOLclD
cZMd/3gk01cTs/GyXaO4KMLpcrWXUiL2Qy4ewRE1nxTfP+JzHGzhSGu8r1HnR/PH
BrD8wma480xEyKFoJBJXmcHaio/ZcJRU6ktHMKcxYcZQhVYJcN4Vsdl5u+wjeW+8
9m30exA2paFW6QnW8/wQ4nXSkc2evnM7wXjtIdhlLKd9GQox74uWJ3jaR1zD+aM7
PJUaiqckEvuSl5IrXcH3JN7qeVM4PV/qWrwvM28LDeROwlobHfDX5PLrmzaWIREr
K/0onrSRo5+vn53p/5HHYX1EX0m/y8nlMqH1wH73mnVmoMrT8TYhSNEeBGkoq929
VlZv/kLQWNO1lU2Q6m/5zzqAuIPZT3Kw6OXlMsPDVhGQnIFxT1rql/5AEFiVOGtb
s+Vyi9fe3OVw9UccWTWCLeFYbrRmpBop+CrfTNZSfjc0Vb5luZxf7MmuV70d4x9r
xrUlW+VuJ+GWd0yLerHEoSD6ObdH1z4wFxbPRDl9Nt2r4nst/PGGvqx4O0xYTRsd
MQppHttWhFPBCPn69vywgpwCQa+7Y9acNapvuizRP5qEnephQGV2sC4f5Jplm9lB
j/Gjp74bMUiS8wUUmWAQFmZHDYsTbX1ANfaBPLKTzyX4as+qzUHn2h3KnAHsWwoM
oVDYMBnRwC8mqGDBzL0z5BwwZUEnxPiIyRyHV1mb0sWdlfLFJH+ppz5K46cySHtN
JcJ14AOzfDqHeNnzK/sPhVA4+jwOMEIoBTlo03rF973dtgo91WTrDbaWW2HX7cwt
S/euZxLRSn0L42I7wOeJECFShVa2WzeY+5Y8HNFMaL9188MRKhmFu82pTcohS2KE
0LUgOBtK3fyU9ZU/V8tSQd35e1vPmFvGdbYclP3c0n7XOHvegKZWtFVwNfFTEkQe
EZXHKfGSlRnE6HCtb1h9Caxn6a/DRO0EbcjAF3AYuzUD72FunGJryFNE9c61JFoD
BoJX6jkiDhvJktlwsmMaxv8cDHB3ZRnNTHNIWaM37MDCHPObTRHtuP0vDY+yMg0C
HogMdXKPmSudf7Car5/GUS7pptk3FOVYlgy3eBemeGkW0vU9//GunzZ3NA5u750K
dQc5pdPymvuurkLOfiV3GJZ30h730vLidi6lkD4xHWDNrXlNMILs3ev4ltP1CG0p
U19+DM/F9SarDzskOgDXvJ9v5yQODG//nK2bx9XUu4X2pff1b7sw687SWAM6LVeV
enSqjxFLjZsZ5DVFXVctU3SZH82kCf5nX55WYB/6ja1RkoV0R7euBIwa6QRYpYX4
kEcVsQx7rNX14HMDhlC4bB0r+3fhMjLyf6+wyB9dKg34n2SiommJN6EUueKg4cWl
nbA1rPbLz3VHY6AyhmalAKfpGbcnk7cqU917DJiN8GYGffCg8jU7JPp5GhqETzgY
iHPdv9PeZQbr8GT30JsJQNQ+Ns5lvf+DqGkECpDOp1ObAca4gsNCeeoTlo8qTHzz
54oMIOZN6RGbP5xfL6uWH16TeqlV244TUC6Sxn1sWqEKO/WTzW8H1J4wVCKl099K
cbAW2yr0GSRcL5u/nt7L1Lv01wuaiG7JqnGZziCENpzsXi+nvWKdXvDnDdiW8CxU
q902IlHBqUM+F0MxAqPZL7FBY7puMp83dZtBNk/A/7H+vbsspLOf2kmlQAaTOCm1
FLtTjP1J1Ykg0yhP6xoaMyZljMsf9g7YciDOY4As/lMa55xnScg1Es9gL9igUO16
TjuhcH9uVv9yoPFtMgFKx021DM/1NF6cOu5TOqJ8UZUBudYr/i9i7ijOlSEm6fOh
qOVA5xXJpQ1B2+Xile11wDlKDxOAgY/EM5X2LBRcUNSXfHA85F9/obBLvwxDVxuN
dQUDhlgOeoyY8FXxqaUswH9eLUICfAURmFjpj9h6vUM/JuXhIedUfTkwD71svYoE
7WQ2o+xH/y8Qv7ZwELnJdFcwK7fU7v3RM7MaomxDE5eyNyDVtddGu72ZFANWns/5
WvtnfnYjRjCL+r5yIgYGagVZ/mvB5GtXok/CKq6JsnJZ6EaJKvQaKXEzUU2F1/bW
9unPBB7RSgFD/WC3uhMhPBw994Hww9yhhEI0HUzGPSeq0vvgtosMYv6rotuQX7B+
VLNFGP+NCYOTnSDUKLWM9Ce8GS5OQqhattPxtigtDqXYwSULQqUxW/Yb+fpRoHyu
LL6agJmnOOD6+j0KyzyiUMqElCKUGp02ltuBEM2agdYJ6yt1kKu/QZvAxQPWPzzx
SNT05Mi+QUHnblGY0dL6g18W0aUPS50zxb7riiHKHkR1qxHDMhoBB5SyCkMN75c5
jhAHNXrGvBl12cwHWqU173rvpFWxMDfKzXR55xhvLIgLkLx0KtUm7GuNeUcdsrRY
lkxh+NRKsBz5unhPmQOKYaWLVf8GiHKIV4pPfwGZ55lH9w0vgM2F6ynV3GvgrYHY
TChw0WDPzqQNjmQGjQgnbCu15bvFM7I1+6O2K5prb8MH9QMpHmCnKe80+a4/kChE
2HLNdjvjmdUdDKeOhstZWns8yOsdMxJI5W2fXGsXD15z3LDK37ozywLEF5vuHeOP
I9bkL97EcOrjl4YoVmby4ajUuqxTMjyteel9YRS53RrFpww5DLm5S6QrFXXaY6/H
mxEH7dvJAnCUA11DQmslfCYoyRcOA6LmrcVjv4jUVPA6P24Zi7S/AEyRT56mgDQ+
EmdNByeXnp3oPYociGXDPWOIHRMPnnSZR6Ns3rNOc22bg6v6OaRL8MQC4N/IGvFu
cxrJ7XxMT7ahSbnVmINCqIF4HSU2wdAgJZfKT77PjzU5ZHRGvIDZFoh51o/A1Z9Z
+/RH6l2v93KKPgEIUK5+C95F0yC726g/34GpZQj6zhuvbHeB5tclfUnnN2pS/REq
F67lJGaA02tzHSAy0oxdXYMz7wzF3zLGe5ed+k2CWzTQkyao13/sPI27X8qfj6rO
Io9S3fM66mMw4XsPuho5W8F8L1KFAF3DojrRkk/VHHi5tskKnQTsrlKgDp63ZCWZ
E7w7TGBztKSPQz9P2Q7UbS8+Z/6174MunkziLjVh6ime3VoTvorai7Y1h+ghPisU
/8Q3wLt3Y97+2A81RQ377AVfDQx/23zz1hOdR7LGrnuFtd+wWs6j14ot6pKUcQYN
m8LH30b7xeqNxXzrC8J48+bqwvg61SBOIbzUzLpzBmHWrbSqzqx125++fUKTqMgG
r2KTxYkH0s/Fm/TSjaXP2V3P6vcMr5lfWH+AAth/7Gy+QD84wXUhBRHIEtTOzMZ0
92VQU/wzRHIzftTOCu0aJ0LlkJgD81bicAW8IHor4lsobumXu4ww0lg0iuzOKC78
xIVkLlq2JQoLghU3kNIQTyh8CohHRbtoqP38yKXWOMyNi90HxtVEI8a18mg+PH8u
StOPYjO5tdQhEHZtDqKMOlduj2Q8Cz/Ta5DEk4SifARxxqpo8pijQo1AiNt/KKc4
SAN89hgA4sBETaUTQ1BCo+FCJ4QGx0znaEdl6jGmdfvDOvyHGX4ZgyEB1sk9rY7H
RKqZliNWBbuoZQvL6gJU2/MisC+e67eyAM8hF8ap6wCRbWjVy3iKG2OUb0nKnlon
mWHBw8Y3VRPPU8w4vRFDkCAu41rBt5DvUO0MJMshg45MyNG3dJH+m7y9/bGVqHmZ
d7H4kuNZr9y+bAwuXyhLMRvRhqbEReFx89CZmh5/vvz2PXn51PQUAKLWwlHEh6DH
ZVPi5KNP1g0xOV74QX0G4iRglr61X74UtOYBE6OJU3PY2tBFDnkw0lJcDr4CGh9o
4jCNsup6vJvpW3VCwUhICgCvJZLfVMM1rVH/QIlBRFtoAR2HaEK4xvz4TR21VdS/
ZPioHXliw346VUEoh59teuVvuLGKy74U05uglEv2NCCUd5cKGGo0w6utldONBLt/
HFvxnrw0gEUFTZ4WTa5LbwBpWD9fSTvdHX7YZLiDZEdAx0QTWafK6G+UXZ6VnYiy
qo8qfdszHLSrq9r4Sb0P25xkGWVOC9rJLcIoPxJ3JgxYKqYq123ZHcmyLacQgnuw
ZR5FAS/0yMxmgwERfF1gPp/iKehYG3Zl/Ycamyg2B1jtVpVGasG6c9/JLzb60h4l
rFw9/2TPk11xdHBnYvk9x6dvl9klu881rWFkmhamx7nAc6khUYdxCAng+5nBX1+K
Q837paEY2nkCJx7KYLz5PpwV6hkUU5CbJwdrPuOG/R5kWQzUAIoJPXUFs/J3RNTF
FBdQnvhjrL23UNcAzl/i1+ovIJH958xxs24Z82bBSEOp7Gf8ssp+WV0GrAVkf7IO
azTChOq3mAkIojvEcjW2bJTxi4G9Pnc2pJJEIBxkhKlVeWKczQsE9k73+GO2wQ4D
Sdd/ursukNCgvpTKkJgrGibQU4rMQC5vUTcJg8Ya8l7WdYSeZ1yrGrS2pJrkWvjx
Oh8beaqGwsBaRMZtIC4Vs1k4BEEqdjb5a/rOleSsgPUZeQVq9n9N/VQwkUJxYfwK
azBfUEUgCY/UfuX2mUb5j3/Y+2d3UblL+6/0YZb2QGrAICNz9TLISx1G5zbM+yaB
iOwpsDmHpIMZZkaq/Je5Bws3aD6vsJ8NSQ3Yum6XUwlTcHzCzPQSYiMkVIQTRMHg
59LYGfyx9D7Np3MnA3U8KGuliWvaUTxY9vxGk/q6boOCRbHA/EX7vxZHvxM+HlDT
O2w3sy0zVOvXzwdtrVF+pNARzrixF8SWo96Irzs0wQYr0xQXVZGsS9GTKQzS/dCB
rw1gV1RT/1xlII6oVLtR2IO0HLQ0csob9pj5a8KykjOLTaXK3Bj0Y8nTpW6wGOuz
kMq1BLKcN77xb/uH0UHYNl9BfkInLMQFdJ44frhd878LUDY/eUQRUdZpEnWKp2+G
FCOc0uo+HZyCkh5u+q7hv7f+mu/jjfsQjNagD2d6/p8zJVUUuxviFvkPMlPsL6Rh
lkWc6g7T+KxSDb3OYSQMAnHvwGl26ub5uJIeTRsOhwMVwfp8krgr3r+pCpQeOTlW
W8OLYxU2XhpFtHTq8R1HeSk9TcEO4Tlp13TRXRTJqJUIj3a2Cwa1Iiaa5LU+cK40
xBUxHCdjv1HMtv+Z0bfqv1qWg0MOli1vfHhaZcCDAAoMPqyiv7RUTUVVBsgHm2Fq
jDesRFICKQVYVimATnxBrv8EB6+M+LhviWlQX1QWv7WxDqE7f0OUFFWzgHijggZb
2L/6wWM0Q9KmYrfRoVihsVqeqB9KB/LmBcpUcoQkbJJHrp4HRdl2kWynvvJUY0rR
/Purb+t6aFhKFK4ZRYB4KbMj0/VffyOtu2GtLNFB5EaMqHIqig41aeBiIibVMbC+
dIBH+9znXSqdgkbltgZ99Z9A797RbFwgJB7ctMHNi0BlW1STNvbeUBVfMIlcleYM
k9NTQb6rxQgbB84q9t5oqG/1aqE8FtTxMjRZGK0DaUhJsGONi5h+qqxBwJc9r1mF
ek9/AhCqNEdw82jNri+aAsIkgIJq+aNJ/D5o1oWIkznzwLfuRDNsvQRUkAM3hoZO
WPSG1D1SiA2KOHIpO3HIjWqNT0asK2dPkVhPg6x9eds7v2L8LjBXbNZaSGABkQac
D13LVuXEYRNJzOB6UBxbY/NW19eKpNZ11uclwR7zG1MtfWSV3ITgDMsEBto8Cen4
M+UhjotwQ50KyNyjsOF8JPme4VWZU4M1g8jFOHlrINq3zGcTGZKe0qPhTGac2HsY
2cq3kmCkXR6X7G69Eqjg+3QkMJ6ycao01v5f7vYUUSvMitX6s+GtYnLSzm9OVSRa
4LX3HhP6yhO3KOZPUCxPB+Xm55V9oTGI+ftBrLZLA4iRW/JFEHngMzDXftqoXgKz
VYvNakTWoDc6reyEH06IIlCVWYkwHPdKq++3rtnkqBFjzCN6WtmMT298ybLOJ832
A4gUtVBmMufrAST4tqmkVpQaceNO/DMmgfecuAh2fXUwkclx4CGcLRM4zzA8r8Sn
+HIxJi38C5Etys2b4RcPSY4K2JEEqc41UiCggE1JrI4/dVpHpQVcNJk8hH0ihQc7
h3xxRPCnER9RlA1UsFh9bnryn00GTQ5HoZw+67U2DQL+B0yWsziUh0NbkkaLw/Wz
bIqup+GVeTDw4/3CuNfM4XUD0qvURegxseJw4KPEi0eiAGDKatTWeXD20T1Q/8fZ
4+d5aV61JbIi7daH1fRbpj6msZTgKe//rynFTrJbJoYmZt7TqfQ2cR7v9e2YfFX5
TS42QChW060/aXlhPH5uxgspFKwyX9KyTWMaWaxR9X32+PWtwmbMn49djhvADIWh
z7p7olDpZJAFev9TLvkXMC+o6h4vEYDv8G1u/96V3mhyJjtgNzZTshIHy3rj/zs4
+R8G2atL5z2gzfqoIoiuW9f8IJ5fZaG3hK8UwjMVB2Qu+iNfl0ipIesxIqBx2sgj
NWD6EBrgd40orcD4Uw4zFiIZIsa11r3jg8QftiYeff+/bmr4JHxodR+ATHgIgqQe
mTo7Epu/wdcUvaFeyG+Ms1Rc/krYpRjaC1sZDD/QH8ZgBJpOjBWparluvmIkUkjB
HCg2KiD9TasJL1aXZLLxzv220TYeZuru5cKU9PceHafku6D+b9O4It4mIYjlGjPS
LmO/9ufcf8nhq5UEQTZ6yYuSF0oJDZdTOHICxDQ9m+Bd7rw8dlcvZKgdIMRjPY/Z
ZhEYQViAbnal85EpMpZH8uYy48hFuQ6+qill/6lmV4axS1ntc2qCyWQsnyk1DRB7
CO/mUuo1/vZ5XssC9NdfgcKU+s8i02ewheY3PL6we6e75gvLV2JLhjAJYGoAM/HS
ka1BbzR/nsR41wds0J40wEIQiP70sK/ltt6nitxLvXAKNU+ThpWZ+8XnXyrBfA60
I+W/ayF5HWtnbZUdei/Bw7HP9qHv6mjRek586DWeUNEgiDQO0//RxPMkyfVK1Xi9
3zzCkTKQAIAxMNaZTTsBMFLffT9b2KOwQq4Bd0pJueE7F99m05Xzfjb+JU7hUPOH
VC1J+rVKujHi/U8I8RUDVmxNZtWBI+G6n9/yTAfFtFkrxCC4BzOr3j3HKjIjD+Ty
fyP671xUB89bpoWrwml7llEiqVhos9UelDz4LxxmaURrTe8nJS+2KhSsCXYHWkU2
IRoMvVnQSCNghRHKw/nXoUvjsdgc1u2ciKeyrqUhmtGBZUgWAEbwpYq1dtvYAtHv
I7Fz6DVs2hChRlj9N4dh3sw/nThWKwxMjra13knPplLvt8QQRWZcACYiUwLcmvPb
dYoBCtxBoIYcGUm3PpbA6URBsFs1UwiYck6O0weL101InB490qNC2v9TTF5aZt+h
gonTlGFcLjxAjhh8htiZzI9fqntyM3+86VTASiFR7TyNXqa5kvrhyFT4r8GoDvPc
VrGi40tZlMRx22DO1YsKyi4Ysu9zJu4vapPOYEv36vY9kkkAoEHDqLmamZzC+7J0
OX3+zpBJUgxJZbvVwqJSJT9BA/sRt1vXGUvbxouuxyISdnzYaL8q9beyCXVnf4Sr
OY6Ruo9ByYdQKrwiuoZ4EL0AAdWZ/I3Qw32IUwOVtZvzdSM+bpGXAClzBxpnZHVR
KupLHE9t/Dmb9RQsGU7ldTtrAtXWkUUARXCWL1HNjKMMkh+VWEKXxKMWsrsJyEUC
FTy1FkQHP5HNnCAabBK1mkhm7XSzRs1bUOaLMP14m7VHoDbVj6fnrQZ4aJcjVhV2
BxmhblmlXUJzJx5W1BBEmFSOwBZKXopsjNyExBHhEjIM6EVJQDyYlC/sX/Vv0c3f
/2viSjsoWc7FzmVIP31EcnFXl3w0y0xAi5UXY87eljkXdcUpVq8id082dW0Abj5P
3dZk6KRILy76Nm6tds1mkmoWcsyleTZJbSUYx7KSUnPixInKBEVRXQ+pRhT0Qx5r
MiCr6a62NFU8l+Qx3JwYIhLkeILhurzCbN1PRjo6oQvQFDdqeBddkLAqyHmvuIlT
NyRchFpTM/MiJRtl1La/mntaS9SjEtpzI5I79A/AQUacbzqqM0rtyDFgnxBk4VEx
3YII2TUq0J4/UPjXyRfabKGn7xMMeeYowB12w/TJskhB1wvcqRqkeoF+CJVDZVMl
n33gbScN3L8Mt+/B28EhEnNrNDhmiRsygyr6fpQRopvS4HqqzOfRwCstyQjwDTuv
0HAXdo0Ly4fGosQGIftVnieHFJFbe+AIB7XNbmqMqPqLxK2jOnhpwK/CyYKll3+t
H1z59Q2uRrpkfR1qmsrb983iXtSxbI21MUAE8mQTVixvw8Yxz5yvzJzv6LvoJ6n8
x2zMWwKyBm4ZMnZOMQzl2o3ELdtRu9r4zFk4/AGc8YhDrcVJyicP4lxlR6z0fBhR
PMCz3UR6A54FCUr4nBpnqAqoFnyu5XdSwlGzqYOVykpZLeEJwo9uBjokKGxN/0PT
TZgG2sDnroXKvh53a3cCIBvZI65LlucBVMRgTTXssR2eZLeqzVIVyqJ3DydZPjke
VnJhfV2VkO4NMJbfYfGaKznuYbAjt/mZX7Z/BTW46/e+PhZ0YkbBFqx77e0VE/dx
5M+txoafL17qWP1rkgc48kbdziV65cDmC9/KvkCZqlU5MNMK1g0/QUXZOHzYkoQ7
66Jog8dJvIbrapoZWmrdAYS7DOKFboAwU+0arame11iyQnef1cODdLibkFi+Uiym
94VyeZaTAmsu4akt4+paP6odqChF+Es7VMpRJ4Q1N7ZWTC4hgjOVZ7FJMzk4hrwR
F9NV5CpkJf7FUaTvDiv+wOAEqHF0rtB0DA+krPhBALDqfThZAZQtCtgCc23XK8WT
fRKxJaZdWBn0XU2JB965re9PoNWzaRlFkxdnUTjeO+uYPvA3QqKfQjm3mqnqFyVB
QGu3wAtKDRf2kQilLg2jdKvk6OOu+jrEmk9um932FI7JrC4U8ky5JaWQgma5q0MY
ghLoPh+/4QBE91kGs0O5ZOFdWdundMI3KvY/lGzzi3coy9u/XxlXjEm7+qgGrUK+
cFZowBeKWq1joHJLIPsBfq8dhsLsZSZHsONMEdYSxnc9+W76f8b/Dz/4PcRaX23m
0DvI3gjZyMJPwGWbIlxo0BCI6yMwT1IU/TfZBDNILBW/AQC4y/imglAyVUeHjBFz
E1xjAZO54z4EiM54eoq6k5hEjh3dP5CuZaMbgt6/cRCvjWdSrDJpIdtzxjM7gwrH
5t/YF93zs0Elz5nR8aqlKVy8T56zTrtfxElySCvwtuu6Lu2ZaMM1Qqrw80g5fC9B
KUsdOvh3kkEgIe/WdULmBMcM0bi2y3NHBM/8HX+J0mcnzXO6c0hDqwUAuvpucRA3
uWWPCSS/w+dB6faCAz8aSdMs4doNnhKfyIKqx/Qa+/SH/ZhRr0KssT41uSstwvsd
o3Zus09K4xVSZVsJK49optrZcLDz/EO4uwtBlCiLbzXIkfkn138g9Sb0F0rQ89E0
Exk/UUntE8g0NqirAyVdsWj3o2eTCwA9BmYHAMbzg+GIkeLfEqHv4ko0aFwbyRGP
KclLeahelY+XvMxYargbzW3cCXT5sOfBmeaSJQq3Zl1wdgMDFtEeRnjngxfSK/KT
6JZ7vxFf6USdyL3JDR+19+a7t47Fg8IACJeVF5mAcYWlDtKzQictbhOCTuhtI7oN
cE2E5lQw6Z+PNKj5qpPvoGIJISksJSpR2jI0WEILfat9/ooAb05YUO3wo29M3vrp
juOc2fuqD9LOihMsy7FIAgX2hW/NrYIM8mGEI9Nj9SXM8YtIkGVrJfdteV6FG9Rb
RC2wLgg4uP0Sxs/IsE6u/qDGOh74TXYmv528OQECkQ8+RiPIK0/dlWmffcl5Ja3b
o66gGjaXlLVyYQyQdyUsC8Y5vQ/tqriM+eEWitVfrMljjYWo5+aqZA46nxTrKy4A
aS1VCwk4XiwGXeqGVeSQx8f0mReOaBh6tPhS95y7r1aiGLwD1KYrOWmdM8GCkgTo
jhfsS3eam2IbNd6BS/ni10wYING2hL/jb2LXzH9TkddR80vDG7Iw2iUGcL3gFX3j
AgtWN5+39uidUt1CmwFTk401/YrgtZj8CaV6rGTq33aU3dsp2SLnLNi917m/ol2s
MLBIdPjE9qz6C8UPug05BBCgC7phrQ3O1vn6Fj1I6bEZFZ/2fPsOzidMBra2277T
4yhhxnJfwZrJpfhu+JZwuER24byRpBnjh1rgafhG/ahW8QdAMTS9HOphoCi899j4
J1Qe9EMXcWdOkoyoMiG4ww2eTvO2x0YBKed6/5vthLmKlu0pvbd1b22O0hSO7OJ+
iYvlxRiRzsFaNxNC8AdXD2w6alltt/UsQbyZm7BgBo2T5qENAWCoYSzioBJaK2Ac
0Pzof497oOAq4373BW+jkiULCXhCsMngZDTDk8dNkGhyeBHnxnwuOngbCTcZrqhp
c91gf539mkbTJ4vL17IqpAACTBQ1iVoloWe/4D2PrHeyuLz3RBMwzPYmg3NWu8R7
B9BgZSb9MXx34wD0/giqe4OTEZxRGU4VG3vGaZObJKeCiuvccCUNSwv0/WPkPHbw
MUTd/GZtDoAGfsQDV+wukEl1hDy05sWT/lhZ4vFl4ZjrTKkVat5EIASeiyEKoyms
czGqJbCPJBpMWWcENbRMplzi0NaH6KJnyKOxEn3s1+ImI5/fib+aCLtZaEdRe/HJ
fudJIG2FwFddj97KdIdozb3VwCKPXVxu/uar1JthcYboWVXCpjkVS1uC+a4HZ0T1
7Drf7vrLfbpF6Hd3Uesv6rlFmw/ZOKg9xevXty2/lRrGCFiaZ4JRz2hfEYhZOpYP
kuvxA4eMoTXNrue6KbWUo79MC/tul68vXu2LuvDXgqKdOANVO3KJ1Mt0M9IGlV4e
XRJ0xrtNw6zCiTeUVAJy2VAAZHeDW0LY/flqReDsWdfsw+S40JqsoCbW/w9Tf/hB
GxVvlOh/ur7K1MG3MlPfsNQK/lig/9u1riFHW6y+CDa/gMwCLmR/NHxAmMqPy5WI
Fk6GGOOnk5jprdoIbu83GgKuiwh4TGyZWnAc47Zt1+QFDMx354XWJ9sCPK9dQoJ0
KMMcfwrYkOhZs3tBCo0ifFvbPsExPdj/3SLoWLh5AwzLYw1/AE75h5k0lPMYlBau
SCJ6lXkFnCaCIO00aQKaH08BHhiCKaZM6lXTKhHI1KjnW7JlH0gwmz5MYWMJUhYp
8Juzg3jCjX73QHkDIbLxiOQbmpoE8+/xNaWx4uHVMNzs5AA37JMza0fBekAtTyRT
xd4sG2Zol82C1qyit6/W4JbmgA8wT2VEWXrBwOxUB0dSr3lzgrHssQIuhjhKGh9z
YeKJUg9bXfaswYKbW0E0MF4fh2Gar+yzmwlVVoMQcL7hftXOPK7f+O1l59Ipjwek
BTHZ1E2cayFjRJj5o6XgOltnYOg7R3fe8196zyzbA+dt/GsghiP72DYJrUhClj9J
+kBw/PSWjNlLnmjNJ46HNR4OYHfWNqJIdP4PTo73u1n92YLK+DCTaWxClLVjji1F
aAZNcx5kSdcYAS3B/r52Fwl/sgGGfghDPV2pSb26lx32hyI8i7rGL/vlWTZGas5D
Df8uMYvAPdp2TfhmVisGw5A/he/uBtgGrimVL1r8XkdFemRUJM3Ev48wLmkwU+eU
Gt8pjjaTcvnNn4KmpEsh1YqREPHzuqCSWVmCR4ndL8+p8Ux5oeyzwgTktuJzcWp+
HXl/6FJW5fxYwdK8ecnE2vjMN/413iS8UIQhFvtT4hLuOjYfTq6K6l06y5VndjZ7
yk+uJfo3ObiMxcwIWbGn5uqyyfSJBWwhWx4w5Uxng0XLj1Cex6pjQ4wUH3RdsS8z
KQOthizTql9RwiwEA+0FYkwyC0ndzDUbTD4IfBvNba2zt+ijpLO0Ex5+Da58yQWv
bG/+rjz6Ad8jA7jPitybGZR7iFMo+RMnCmaRD1lys1Kh07xX1TagTDcP+ZlMw3Mp
LGgJl1INbuJE4of5qVWOLmQH0dZyTcmguijugEs4jNuS17Shb2y+qLBJUBRX1pZE
mVMyiVp1epPw3KjjSP370t0w63f1pkcBc3ngDmW9VLIWWcdanzwnQwDmnD4iQTWQ
bj8yqxL6Xj9U7pbSirI5GBgqrhQzj3DzoYVAv+yeDpGlz3LprzBqQ1mLq/FjQYwb
MO5p1A7RXPsCFMRCMfBtc3WIpQaPyEzxGTYVBmt4H1pO5/ETe6l4LKpk78Gc6t7W
N5ddFhVfa9DzVjiMCIqVmKyYjPPSrVFJFfHf6yPe9qwzQeUG2uoj6/pxahvKtW77
L35dMT/Uu8acgNXR+94cwKoLfIRCFWr7mvDerLQZzTM1gvUoeJBZMF6Tdcyv5mbi
kbAzOunnspBCpDmme+LgDmYWCrht/L6vuowxlpVbQWlv/YGiNUDdJs2Iq+fIo9nK
qOx+YnT67p6pK58K3FJa11hoOPxwZdq4SAe5fbOTr0gnP/DKEeqvzplbFgcbWex1
FFHfmKjkyT5U8fBTX5cNh6uyzMtAHM9dzWhp2CItDpL+dNygzS4ACwA+cZ3MDxW+
2Mwog2MIKlKbjOqa1gnKthPzxKKPRaGb1WPhEPGUSfYmdunfJ6xGoZ7WrHLGWg3u
zDBG2xfmOPlCYmHuFCVyZQL859/gz8Bt7tIBgcLsYx9FJJHrPPJR0cCZrzfnZLuz
Ke0lRJ8sfGPzlG7gRbCLLc7haUVR6DLG+FnoEoYTrrP82O0lHgayrp6aCpGi4tJG
rWjICWCfVhP62nNBTFpFMBFv5lWavdj3sX+eRSjcZ1m+/bH1kaQnTYBGRU5ZlVu9
fewg65pM/j4ZcikFrqgstpe8T+4GDeMziHVTa5eXIUwYllsCoQsynB5BktgXtBqW
rTojSZqnlwDEZRXwVJCHwKpk3xcnLYRdrE+rXrZMUxvGM/ZglQyP11ZX8+yToVTF
QMVj+ebDTMDoFHieU+Q8lkl/dGwRRWmqAaNt2VYyIRpYa6UbVs1Eibvvszj3/NUN
jDmA9D8wUuNZNP+lRG/gGBLOD2bNhHegSfdaYHUNf+yYHCbz4+UV9YoX+LHVFvJ5
cCo9PSaxAQQv91MTKfsR6cisO/6uul4nyRmsdD6ASxXZ5ZW2XkU7NCoxXUWEJ8yt
hInvnLxYs8UNJXVmnG2OXbMx85ZiCeP9ffYho2KULteFoj+TmUnUJ78ytx8MSofg
jnwbo4J8k2kdbIurCGeIHWDFiC4Z4niomAKe7fSHy9CoF2zJzUNm2RBfHPF8UXDx
lmoQGag+3DlXmyo8KMMfHDc6pnQZxQm2FaknKWCfUM1JusVLIiGPkEqPdPxBJ4RY
oEwK98KnKjqPzcEGEZWUfFQb/3RirjlV7NJwOhmnSMxbSVGTYSbnlHXz+lbkhndi
qO49tlGKky+G6HVLO1pRHU/rRaox5Aivqp589GglEdEx+xATufsVKYEY2QOGHVpg
rR+K8lsCOfpZryd0hZ2rq47IF9iuTf4Y22DoBXdxdRUuiVJOUazXdUfDMr2QZxgb
pmgGLy7dTcfCzBtADA3gTEPKViUea3wfKNH23SyYoFfAXY0fxjfoikvpJRwFejb7
hrd/FrHlp++K2LnGzIFoPQxFhyaQHj8/KgHCz0sYdmTDOQ6fhXZbIH7LGXWkQfCl
I+fFzr1YPHQg9eZ3BumDrApXzM9SEXJqvmVSPkdG0791g49BTXxDc02Uvv+kCZRg
JSxt6WJsbrCLw3OHHd/z8uYsyQkPBLoAYQcbovxbLbZU5Hp54KyxZnNN6PpcDp0Q
8k6mnBtergjVYqaMXyw/vNP/21pn4xHyNlGFAt9wVjlvrpbc0YToFFHxJcb2t5Ef
DyhcGAAN9BPrwQEqkNwrL04oBvINKjNO5bw+IK5Z6WSzZM2dVIcqRTkySMVG33z2
alWSIMHULuxLIRLdIpqOEb62PkvK7bA9fICxQcri9LvtzJj4VipcthwTPjrXFfFg
n6Ad6FPRgJc/9r4jOGhFapa6YgeOQx2Gr2f4rx19z1NVY2Z7fKHPNWEPRV+SlUa7
xsngK/WtYEQ061BgEP5A37dc703ODSVTez01YNMRlVQCWoJXKHMrn7aNJ4xtswIo
w8O0XP06T2xRoDqoIqm9+YVZuu9+IWXyQxbxj01iyA/Uog/YTPK9YOu/ljtNMqSR
1vWtBJwFFMpnDccLmBuxnR7I2238gM7uHtb/ho4O8V4ji48Xl6UPhJLI/rQp/gKW
qK8RBhwWsXlHnwWojAdfiYvT2WO/MbK5ZPLEXA0iGD8J/ZJTA7b5YXzpcaamk/Wk
uR2DM2UD9i303cUyevnm+xvrS02913sjOsJkfNN2bQUCHiZDFLge8COzp636G+9s
mI06VVUw010FQ8rjBPm44ndTMUl1RTyr1WfG7vuEhGSQCeCUEyyMThZOCdikfpbP
E4h7Y/L6qv/oCpG5ofTIHHm4y/SRYCKQT9HzKvPnDCq13ho/AlLZjH3LedzA8L1I
XNHmItoWaGJn22YCdDUsmvKHj12N21O0S1ktnHa1m3k9HMpLI7l6Xceai6+b1Zo5
eFg63weZM6xLFFU7VhsHL6g1n9IYeGpm+xuw6lPQjM8OMEIa2wVweuj0xWwU6RSh
OQeZ/ejffRxS+3M+CaHV/KIgs0HPyApBi+UxnmBcuxdZCrXjI50IOi/UIzjC/NXm
ZWDZuUk2kNRCNR/XEH2fIvi6DgvlGPNcckxxHYPxxT9QmoLgpD1OEHimal018JEb
ogrYwGZzxUxU78Lphd/QodFOZhiL+ckg5smLRrXFwr6n7f+xxjTdxY+GKJPHYXDm
W9TgRyaGInuGAK8fUQ/XBYJYBYf5lyuczVJtT2Hb9O4GxO10Fiy7RDvIJYfZX7w0
RVLLfN8WYNMVulePB74TfsoeYZQGzePQvTzsi3ZKucX4ak6P0lf+iJTjqXyHS8gB
ysXCjxQwE6LPj6yL6wwTiR+UzeFXN+h7SWYSg22Qgv8yWDXX5SQGAkD7+LqLq3vL
c6gflFb4dDunPv/PrrIiohoUZCqUgPCa5Efd8GlpdreE2S7nPlJHNynlUeYOH705
x1fAOKFq+V+XRruqWUVdx/GZ71N7ol0Q1N4WCCZC1Wv95ieEQ7T8cFOydTzuIiZw
6Kdm8/Rt8VzzOB/SfBmKHRknCRYbkywtawnwSB15JAWO1EiZZRsM6eH2BczkRrkW
W9MGVqPTmszfRYHi6Wp8LJCKOlMZ3pWNnQqIJqafJBgHS/tNohxiDGFjOMGi5Aq6
rQgpFB8idd20Kb+H3HZHFkdR/hEvGlhm+abGV3FuWOjjkghy+XtRtBoDg30CkdUF
jXiJZHgjOmPmJI+irEZjiV3MlUinxhAPdogy9IdIdEXqyOh5YvHJMdM4/oJ7NY0p
ePzii9ROhyY/GxTz6U6cTycpkQY0c32vp1YNPra3QoJNrEkp24WivTPcJSsZhVUJ
Oyk9OVuNJfqAJZB+lPr9z4HNcHyW+tz8T/xmI1zLIedKv4PEwLo2SyUHu9+IwZOM
1d6NwtvD5ppX377nsVWMdBRz7Kpdy5c2+SwAYMdCwYiW9Oz61EF5bcbAr9KwNOT2
9GUXJfOQrf09laWyCrlT5ttCyx9qv2kBD4SERL2ZnrTRaFgA7DBrmlxmJ8+31Gw4
FxWxxAyKO3O2jSPEMHwpW6kJJUDDAAsDBXWDALJAtxi2b1D0Xtfsn0Wm9pjJgFh+
jAzXkN7xtVUSakkqj+sXndSrg2U1S5HfhI2xR93KVGOZ6DLEfyH6jXWPH6yVkp+d
0KpMyuoxMdvEsHrAQEAfVl15Qb2iFfo+asqywPVmlA30026d5pqRmkoD9xipEKdJ
PB4kYeZkidFhJhu0yF6RylntbDp/gw1SlbTPIxj6r0JgysYauHPXpKLqyH9c6Hv4
RvLs6/WoA4O6NMECsOyFWaZtOB8Ek9M/sSLT7UGF9FUsjNuFlIDcf/IyqHb1xGt/
b8rYgyRsPbnfv6aZhNvGJRpg2l3knsWDkMIj6mpx9aU7R8VNp3B3DsyN3FkgQ2fc
wyrmEumKNJ5hhU/Iumrp0un2YUDun25tOdgQylwuiM+w53PVEl/i1mwEv6PKNCvo
8/EnO2NnPeCV1APsG7ZuUkjqAjeuYqbsewXVIg0NjlqjPRvzQNWoiSTY9sHvRXcq
XP3LCBPZIjEHepE84vFJYeq37OYuYVrew2GHtudiWz8RMiC9U27ZkfiIsamrd2B1
MwreHVgOQnAW2HXECI/usDLuy0PoViQj8/F/klkUM2MPcNx2xAmjapjfGj/BToKj
oJt9Rso7unPfd+XaQWds7h0wBfufuoOTK/zuYycaxigQuSGOWRedzcpF1+O9IS8W
qntTFx1fCxFHYDhcYy5WvShcc54yW9e4T33Lg1zn4dXwdOX7eDU/ZdjckjzXZqPI
v16YxxdwombTWzB2eMkSLPqaA30Q2YkyD+Vm3CEqjJEtw1x7zD03TxRNlOw9DCFB
qn9/5ad9U1lIdKkOsyiHJytnjozGIQrbSkdZnjCTrbEvgNJRpYS7VGhFlnMiNmV8
L58aeJ7N7vN1ZDnKhwwb2ztRNV4SNq7oFZjFfUHfIerdZ6Uc9cFuT4gDKLJqY9l3
GogpCFfsldb68WwczMhFCCvhP64QJR9AmykWoHbUR5Z8WuYIIGI7vQFWdtwHsQTJ
OUTA5H8UvaxGkBi5xwRW5tcErULXUzVFUDydXy5CleHLqFUFyTay6Day27yUxrqt
Lrl5TVTliT2qG1BL+N/SiCh7mm83wrnUoUrnfJpAfls7oVHKqAcJbQUZVpILjz8P
Kf22oX0NLPoyKxtrQ7QxwtiEEwiNBA0gkNsotJLmSdYeTXr6W87iUHa78dqk9om0
/rD6XZwd8WQZ5pU8mWDWvhDF6Aw4f/ienhbt1xgcKay5TeQz+FCFpFZdkeCbr541
RCc8TQ2SHQ9uUZ/6s+MTfbLL0AWKNxT/Ke8w9AZsbKB8VTEUeyDeUfcTBwLGx8E9
T6rHc5UIHOQXlXLK+lgOGWnnhI3iZOxUzLDJ4rFmgSnfl9FOm/zQdBbqOfYYcyl+
xvP34XaMK8MVS4ZQM86NHVARE19aMCT7fonpix1uOjdU2cxDqRhu7hciFHxEoWwo
nKB+Q+B6v5z8I+KPagI8mge8mn/gCpAviDUSnBBWJ3phhzg9t6vgBz7olFKz/HMD
bcr0+I7JL5IYFG5azbcVRsO1S30Hnx2nq6pBvX/LyNjnUaosNx5CZdGFv2Awkr7t
XBAqrYd9K2t/xYDebCbNa3etbFn1Y15e0YUc2TNey6MwR/jK31HXCoFUBbs4MkB/
N+Q3n2ob3RDuDwzipOcSxLM6nsIZljWmxX5efokXx37Pf0K8/3cJJhh7P5b0ZvNT
/7O5yeV0LQBzo8db3EAvrOgE0fspAGvGJLkwe0CCwq1MiJWfNKCc6FRy3b2lLCyX
7HXF2VFtn+XU80ZNDCRUO6ghwwh/32hesBTE7bFzxc6vI2N7i+SNyYQaO/Dn7422
OtvM0akn+38X8SvOayMPMADto+2PxssgVWFOR3xRf35XvKqNBRw2Xqjrt7SN/WKo
/07tADjYsAMPZ85IbZ5M62RBtWT2mXTviK0zB5mE+v3OEAVrQRlumikXTrxi8yot
KjR3Sd6ieMYtI2maG/eVoJ6fP6HbBwmU1NAtShwPPx/V6TDCg0CT4qGIDzqJBzQF
3ayAJ+t7yWsmFakE8vvtsaC6j4KqW4g6N6/YQjjnmPu79MKDeJPpr6WON4JUyoTw
eYMBbyh8AbxefhY5OWH6D5V/s0ustVjGnU6HXQacupJdid7qlzRy1ziriJQKsRTY
fGNqOEVlmReQRUsPO44LrmLnhD94uW1EHKOirS34Dy+29ILFMu3M65eSVbwyQPSZ
YkwIS66xlqUvqpDGR1jJkpD4XQIyEaJ9NLkZGPbddxozBS1vVmomRWmbAqfV8FBa
Fd2kPZTv86X78WKOlWBippxXSMTVu7Pe1WQU5jfT01JBenSqug+EnO03ctxRmd1p
lPlmFTLmn3ZzdgcpNOIOnq05j0AnUA49QRAn7iqeHH1vBvqEzz5kyPzCJ+5RLAIM
GuPq5YJgFQByBQpbUM4ZPk00q8LDTvrTW5FDritjxJ+p/YWBjwtvEsYa5gZFLYzz
pIcL2QUxGlrpSvut/KlmjNMP/ShbKwaClcS2HLrgx34b0AssHq0ELcOw7t+XFREt
ZOZlf3vd64NFmYSnDqA3eww40VFfmyxpnu+hH8iyopzgttosrJ+y6bJilUzof16h
0ucfeg1QXZwMgx1oslZRgE4uJ96UaU18L7JT66wQjl5pyFkfQ/0WkN3I43AoDZAV
yT6Bw5aaH0Cjtlql1Zr4nXuUODw2aWIpAYjiPQ25aGIvCMdXAxCCGlZIO74NlZKH
oCxN55lHwnRUnV67r4M+dSz+pc2SJQ01hLINCSaEhV6KWkcHJsqzG3mmicBQ0VZi
wVG1nzlGIxJsRLgd0Mh/mLZ5waoFc4yVjWP17u9j8TAVWDzYs9xCNLgPmWOHJAQp
B5bJd3zfnVhKWKtYpcl2htPTHkb9H4tRiYUYYhNSyzi0Ox7bZ4BEHSnGXKdTleco
76oxXOeMpngBoWEjXCQ+QfUEuG8rRHmeDf86yodt4FqD7rtyEnodcyQ1b803gx2N
xIP4RTm9hvqh3B20PNXK5fAyhXTDeE9L2BPj72efoDrBwUEAJvayJTgwSk99gyqG
YnPacX57ZJIhK6EXo60lnkvLCBs7SJeDpUhsqNV/OWHNmPsJQmLktMTd9qFqen4g
PH6kAT32578IQk3V1a6OSOQYZrE4nI5d/TjCdeKEXLXpqz3sjl6xSKbepjyGnLVm
GkDjgOgQ6F3iy6p8IAijZ3SsUO6km2Uj7AUjlXj5e8KB9WAZchSJblSy8HtzlpS6
BNxQH/VGp081p2yTPqOOP9fqtES1Cn8rRjHztot1kt4ryVSK+F6LvPg2/dqyw5lM
fnbZJ1C22T3kcKybjl8O8Sf1zi+SJ8bKuHpqHaYgfX+3+4t+VPgf8K6TkKbR0G4J
eGzV97mFNIdrARGyhPs3D+QmWOxNBqthKiO70YB3FEQJnKWyLDB9dKYlfTaGbwNW
zCsqO3f7S7S88RcgAWkYCUP0sTeR9I4mAjNJXkpJD4ADH2mJqlbHsIMR94/ZzwjL
OwcDW/iUaIG9dMtwLa42nml4Wn4Nc4nrNNLFEOdl/4CgqK6VpPUwjamN5HWkL9X8
f8QdBtylwfTPRS2L6QIVx2TXAdPHq2li62Z4ow/INsOF3Tl45kpdvHnZLqJKZykW
q8SyrWZYd00p9IghI0ROie5oQ2TDSVd5Bjlap45aAB+Kcu4PMNZr8ZlN6yiORP2f
s28OZNWdeQErJxyHFYeL5ikSYL4rBt8um1b0m6mscEPBQpRHxskhpO7gDXL2COP3
jbSTZq1nAbpH36aahd95Mnvi7wQK3iYMLVlHkQuktsRfleW+zCKbRx7+T2iWGwvt
r8ilKtl0BsBIeP2pZXgAkVhLqGcmTZATJmaqMOwDznntZ4mp57IEQBS7ROqK07wE
n+mDu1GF6tIWaP8SoMmu0bw4x1MfRacUV+TncQ66M6+uCagycrhux2JV59O3SSys
4/+KHKlA1IAR3QXk38e+2GZUlYO2wSsgvMeCjivBLUBD/luVp6p7Yf8yC9gdXHVI
fRvndH+OZj+YbI1u1QVFO3iSm4/RlZH5nCQcDaomfxwzQv1ppIXmgDyagpSXWp3r
0q0TiQDFmK2GmYBfbq/BRjb3Npuey6YS++E2bo5scWO/RrZESs1zjpxP0uEToNxg
L6gXvqnYdxH8fL4MjCPRqEvbX3UPfzk+MFaEB8SD+gM+mZTane5KKG80r1AotyZH
BD3WBS5936QxhFryHeYnWfB9fVpPBOqT0osRj2F/NUqSrBocCkiOrhuAXpXm9ksF
QkK/5Yxt0w8PnjUry/+GgPBDL1F47JalkZ8doVkiusWNcvgrEpk5eJapkP6j5hgK
1DBBm077rw0ZiaVhZodIvdSKT/6Dae0RlsiC+WNqrbZDQDxhz2LtoXUg4EE7P+07
zPmGRXXyLvCxFM4yK8Zwli3/b8FGb0WRI8Ex4dw2FIAnPpGTSYDJWM4AtZ0DkWHp
WjYCvw4vf287HdAKz82SQJ50nNfabNFr6gkNJxZg+05hkS2HN/uoZgAx8MhR98yp
YwMlIzwxJzzdBwZl6cm3ivxLVPFCOUc7w7xLO04SLltwq2BloVZxJnxGcmdK5FDw
GZBFU31nGAovmC16V+BVyHSMNMzasbO1KvLa693rVTlQHWKzT7KUf12FxXLR7WCn
TcRgvceNoNvFRrPIOIZskSNhY7M+1tZ2Tl+j/KF+07vTQonyxrRT+dG1sRYQoNyt
Hge2o2QrBxoEJgWhp43qx/xxX+e6c/j4+xksiBifxSXiCVw78E4rmLEK8S7ErKTW
0+7cTVcYIocslb8iHPsgI044wIrmycS8fovHevnsvObXiHNNdej2mpi8AnWAjQpy
Jx+1PQhN8hCL+KT/3Z2n57RzRi5b8Mugk6NkvCosEwI5nQrXsN/a3hlqsm8Yi0oK
vro6x3ZBLQqbWUnOiQ/3HoMGZ3WQ4P1QO9hu1F+bqLv3vRdBVIEq4B1Mqz4YuEmu
Ymi5iHu0uB2NwVlaHLgYU2uWgfD/VDTFN86WjvpADUnHF5zblwSsKYKsqnLawjHE
mgO4owhboQFm4aVTLBlm2odqUrb8Hna+CrVAIJQpM1V2bo05+VaP88+GuNq3gHl8
jmzfpxlweFOwmH2Z/innW1rg9GuKPRSYTwnvJYvjolTzKVmcY60sdBRIJ3D9zUB4
mR5XvXzpABdyS9dF60gXEuVd9GlQv4Ci1XMzkXJFRpxCdIS/5B79C/uiRczQ+Udl
Fd9q5SllYYWj0OgTxl2Xz+c3zOZxe8CVnidX3Dc+wdQoM/zKWy4jkf377nj9qyIB
oMi3dQJAJueOFPvSGSpkL+lJcj3dRkB+WXxVkI2d5Gh2W9HyptzEdL/olaoZVq9N
qd9GmibzMYYje585T/EphzfbkQiNDKFLHQW/R8NmOlnSU63g06tLoWSTKwfJa11S
4/bb8jpDcl5izEoLqsAqLD08VROrTdcotbMfr4k4rb+PgrUBqNqnzPBGBNqi5kDQ
Xl2t5N3e48CtfD4XgQVMFfXnApxMe0YEmOTHQrFBxi5Yjc64nccV5/0jAjQq/krw
902eMglIKIAu31UyV/jhS2Hj6ODZlYPepyDWVgC8DZxAOn9TovkkFKQFjQtbtMLm
5q2Eqhn0xKBzMjbn9tKIe2fFstvdmMCQ+aXiJxI7kPbCaGpVihf7u/1jUQ2oosBk
LzBWQUOSycm6Eyz5xebvdNdFfX53Bzs12P/RoXij/4rxFBDzWMrcK45BS8Ab6/cR
KoSXF6AEk+x3BlblmBEYwqUbhKhbArs/eGNFAHJ47i11pd2mjSeJV6QBc808uZHE
leFynAkJP9oCmgYuEm9zQZo+sK3rDuRFv6irMIe9ADr+n8RNVsQs/uM/StBJidUA
VlQMvv7jF4bemnR7UFWO6UO/MDUHpaI1AXhBzoWbkhACqrGMUWDV1NoJqbSyZRlt
bA6WZs1QaTUtuEKkQ+E4ufcS4ZRf7iEXneuvUM8dBYprV37jfNfN4w11nPS8G7+N
CeOSr57m2bj65dU5c0JgZMNzdSaiZ67BC/4o6Gm+8HNpNjQemWrY0QqjHqPkZMGM
m9NCjWftnXjy6fScVuod+VLNBFmfBdmXxq/tbZ/TtR62xBuyEjleAcK1UZO9hxHc
oCJnPtUlve2uqIY4mTfRH3uztWxg13UfsIAbj3ScUtLzfE0Fn3phYovDib/jnfUL
BFITwAoL28dy26atSFuGj75Ydi6ujIiAn/vf172Xptpijku2Mx/yXNZ5WZRXGVDE
pim5pafScsAFE4iclCXTQnVrpY6RFae+QcYVHyNo5s2s9wlM0L9OWDf3G5sbQW3F
3EcWbz7Q8eWHyi8vOLw8xEOg9zR/gfchs5EcQztLiS4FnvRrxDrwUzX9gfrST1gL
yWi+BcBgxXmGUmHIh/iF7EA8B41AsfATjQjGp9sXI4AjkBn2G7rJstXieLlw5Vsk
YmoBWc8Ooi9T/Xz8/3QfqpV2jNRVS+rvnUDl2FyGjTNgNJP+RMs2xDfN8rNKbntD
/JPKvt412xYUZDMoRisfU7Lba0qMERxEWoMjic1nGh7fyxgZg83RHeReSzx/IMdz
CmNHUs30X/lfz1N6PEozo8SW8FXW13f2UCVcgeMFfWFttwSQZZIY50w0pb50WdwD
6RULrGMeCDVxUjRuuGvmicfc1aB7NnTqsbUInsZnZ1jRHaNL10aZgqtR8QRyD+AT
WFwY0NdfdnPzbu5AB2H2SLr3wpvpxOrcrX862GOdKAp3QVRbJQA0o6HrsQakQgCD
JqCWd/ljYpRCq7Sc2ig9TN8XjPGKvRQyZeIaGFOtP53Ur8dt6O/J/qAxcfPiMyc4
NCxZLgHQXuqEgXhGcXxXxs/a15Ds5FyuWW4zOYRpuZ/C6vhwDdZkpCyE0CQESB1T
xhqJhpHsX/pki5XP8x1er8dKMwysi2AH+BQRS/KGwe0OkDcu4mst4SqE3ISj8Xxx
wFj9J1ymfr05L2z4mqtfXSB1drAd2FgS7rLWrvPaeH55I+JPap6YmtFa+a7RzqYb
iWrQaToedBl/qr1IAlPMqKo6PaoiLNysKBntC5FOfA33DEolfM/4V10GsJvWe2z0
dqfzDRI/VmKXT4jzVOZimozTqjCiSImK0TwiPk27IXMucXAzJS/t2u+1yfbyUBwu
UxBidnRIedMUo0OHZ50i+PTCrDpfWxFCnISGyFu+zQrqGgdGTNgH87rQgSiK5Ds8
qYcRnkEfZZy8C2pfi+2xgVf4GIJ9TIgHSApMI49VwhZAPVYBasZ4DgRK/Z1mycCQ
J/tkFejVwGiP/zqpvojXbKdNyR1rbD0AVLUpZP8/lIZYmBr8ZLBQxQzirXl7+9GP
KSUNLpNizAA/BthavODJ55DHdt1COXOkvQoMThLyj5/Q3RFTQMkAAr1X+j2DjzFS
dfuiT7qXUJsAi0FUr4+2l7uwOTB5Xz49je6sJokprP55YJrlwguD+5npAbP5ozK5
dIooyO8x/FElXQTRKQQf9RGc5WxeC4sQnK53s5ugRGORBpfo6uhAp24EnHnFiVse
bmEL+dva24yxqa1qNY0Jm13LEHQ9k/x3R919c0Us6roNkOITzkU/KMl1AOcHS8oM
0F5PxvpLOtEeXBYXx2NEGjm6oMi0WY0BF39vmMFkHNRWWIxAlfNXMy5us2NHQc2F
6XUvv/9d4EvPm3oEKbigkd0VWM0qOpeTCvmTan56Bs09wikXlqKItTbcz+8O6l5J
Fy+PwRjNlQzlWGQE+0aKljLiHxRZd7JNtZU6Am5+h2Ayb4Kf6Rl4G4qMgyb/hRip
xcJ7zT8cNrB4AptsUYVoOUXdHtYieNU4xIQ9UpTaln2/fa4uVI8OHpMEBdDl4uu9
H37J3yNHjB24QgD0K0hRmvGujyD1Fky7v6s4K5hq73F5DkTHMQnaNmUVKe0gL+iq
WySGOUP8dAua4Nbe4TEbocJOA6U39ckw7UL9aZjJIb43etfk3OBS+Pq05hT5t5da
Ljjzy0f5elOzNHRkH1LmJchnTGFOEDVbiH86yr0nnB/FlAZS37yiS/QcxlGaOWUR
1NM5e6Nw/ctv5ARo7xHOw/Icjn5QFDnZ2FQrcjyNJ+ryYJsCNu6ABnmHK2sRFrIY
zH603A7ZiAi2WoNUCOicdjpULi4wURYqCWYvh5SgULdTHhUAR7TAKQeM/6CmTjTR
R5yGZxq98aDc6A5/Gokp/2pmlCrSiNSGSGQai151v53cQfTMe8+mCcCNNq+av9/w
F13rnNG7WzVH6pckIPAcKsiATBXzqczfzavSuA1BFpt5zYBZ/QJR8r273cst9dgF
WckIouUc+Dr7nh1vOShLdJ+SysK+SoEtGvL2Tkn/WejhuC6TFp1rvg6gGl6cfOHw
k4NeYNdEBmuQ+5GL1q2Wr5jGoAyMvwAcl7CZFNqjcnwaex8NneHUyOs3lsNdmIi8
OOjEqATnDqN73aXeOFv1VchPPpOt2idQduCh77UvQvYAyP3n91gNAJRq7aJnyaEO
zDLp3BMjZz5H2O1VFyoru8/0v188Gk7Ox5978dIStLwEubBambCPeawmkasoomll
lgtmdumMRlR4ipIzql6BEJ3+SC/aqheB1m0xkOhsdkzQ2CTd4avog8VJblnNW7wv
0pihUpPvRtNWqzwceECt69TcdFptSxr1g2eUdN7dqYJt5L8MWMW2zhMO5PZrpXvG
SE7qY/0Ex7Ixic/gbKMl7xdwb5xiOUHZorBAJjtlWYIpBO37UFO4N0Sw/aumFR51
AuD9sjdLv9SgqN5yjHQb9xxzZokw5vBe2/YarSl4PLYc1t+psKdFI12P+Cqs0adt
dtfGveUkW0f04+kyin7l5HQHbYace84Zm6f9j7GiJ+Pt04Lh2gTrE4SeFpBdRrFo
fdES2frtkHyKURytj0vTUCzFiyHSp0sJ+6eege5/jiXwK5DqTxmMks7HTBDeUYRT
fyuDViyMgpQPe9jLrtwgMZuoxba77OT4LwWoiHkapoElhL5oNFwKz66gQY5wWx7G
3QPmrkqHpXp2BprZYnrIZxkPFEasvjUHJWA9uhaelcL2FPrpHFuKNQJhc6HmB3s5
etlL8swdvdtiAzHlP0fppXUHJKqSCN3On8GvjQp1tMlSwcomRvgkjBBqb2q5Ti86
5NEgIH9aJVhfBoYXRagIdzAAn+6Ijw75FC9mXEdSVSU91VnaYLDavALVoYcRaTRS
Xz/i+pN3CIYVR8ZQlSMEEMQZTZs8SAKrFD0PIT6jS7h2KIvf6lQsAHj7VQlOj4l6
+ffrOsQ7vvXPee9nFrHnyqsiHz6DXX8xejS25qgi8Gh1Znbo1NgUYx3Cn1F/03Ux
RgcEbLRUkDUMdFhcO+aDEjeUwjWTJH9c2rxrAlWzOdfelYui52XxNhhf1UORyQjT
DdlrnYJcA+YByAzsEeI85BM8hwZEWATZUXz2YqZC7Dp0FggiOOkHyqDzHJGM6YQP
ybayLxlRHCqPXqCio67fWRlA7vK1M2Af2axJqnREsGFuDeoX9sCQYWHn959E2NyR
YSqyIOJmc6sYNGC46aNlWjRmk8s1pbPZglYtVs/8FMa2f6wQxkpk2yMFRvfEAoIx
Fssp12sCsGzfNJR03y2eEJwfq2IxGIUxSGRc2l0kWoOgIVhuA6sh+c1Wy/fIFD8r
65JR1i+byG9e4dMcX5Plp/uhAtPfintuNO+YJ8GAUyeH/E9sqweYfPmuNrHNRvJU
3b4oy9j7GVO8U0el5k6UNGWvoQ2wNFLsByoJlRQbiatab7tXyEf2/pAjMWkY+jJG
N7eWMTV/1WoP3qQoJ2j31thszgv8eYDI7fv0vjJ1evxUSMFlkyfoRpfwUDgjjQyA
I5xsHfljiZeB0DtKwY7zdV2jAfFgFMZaDX8mFzVKFSXzrhgz3mjzZ8AbY3Oes2ST
fBiV7tadDC+edpbACQwb1FlVotR3Ufvuit6BIhQsD95GYi/RFmI0kRSBd6YfHnue
AAwiU4r5C9LyEekSlzXkifa+7sFA4dtpn467Gq4ybEoBBc3bu6SgrExSc24Y57OK
NtCjVV8XGrkbSNpY5dDs7TXcUAmSG+uYNZMflrWVgQL/Y0FgbK8+DfRuGF1jUcTn
210mFnY3DpZUlNnEckll/litTMZ/RqYF0AmMweoFUP7/mnp0+M2yB0w67ikJCc27
8vua+sj0c/SNWlCMisKpJqWzQ7Whc2Rhlxn0qdw2p8oukmiStBeTQQTaeVYBCNia
0nEPqOR/hpPi97+f4UjTa47swIjuBdGZZGKt671X5JKh+KX500PSws9sTduy3QPu
B188jlR0SLIXTM+lCvGKkvwoj/C5c/P+lkvZFYiQC/hDbQyJ82CqlM95kFcmF3FM
GSD0CQd8bsyzF8TytVcmEyoQ6FUEsgifClVTbut2XP1d9G3gSVf7HcRpUxjF2ugt
42/DL5hXtcLqaDKjIMuaPv0QimHC6uV7i/PBliX8wbXr/U+aTGOX7Dg1Tbmkfmtn
ZMw4Y1cERLqjltJPrAxuqETz7bj0hvMbs/c1GcFce9djY3j4OUICvIN28qLaWZcJ
up/oWModjP93rOk8FW1At1S16JogN+hSy5EHbb5oDx5dpsAM4/84pMdA6ocxITlt
nSMRnV9MNv8a3m6jwo1PHmXMiFnI38Jtq1ZAmagQ6iupjw5J2uN3GSnYwqPspAQ9
pYJU+EBY1xPnqiUrSsmsuasJXWGK4O8b8kiHEgozNm0ES/2H6LWnkY3JA8rMbNbM
AMEGSn5s2UF3x4S47Axhmk+V73/mTT3LLTp9obzYCEHvoEi8xuBmXkDD9fLUfY+N
srRZYrjPCwYtdQpjr396Ez7wq5wM4M9hxmubTImWJnE9+3E3VpmtMxu4WH5OFvNk
vB3FpIzy4GihHXUwIT95daQv+4pZpCo9Mk9UQbS9mV4rcdtzBRslOah7Lmh67qL6
+MNjRff+AqWOL8HB5A5eRgompFB9Uxq6cPRPvOS2QYWYxh7liB4VnGH1mSOIQbRg
MIOoJBAHIT8vIVPZCaYOWgo4Ts7Iz4s0yUhtfuRtoBIice+e6Z0o3AxVtwRWfXlH
zQ/r0s/2KC0KQ2P5Amv6Fy7mjU/PkVg/Sb1b5fmm9Gg6rolSNNgEt+DKrJqsWq1E
JXNl2YTQTBZBi6HYf7LIsVfRyqFDGrfJuneUtkwFu0PyOI5I8K97rbwa/YNbl8vH
UzEgJZ1LIfZlGU4bFOBuIBdYJHEQ9q95VBzNIMMKux9ZDdZnSXBfEeNQohtmV3op
OVz1xgHcT2xPaeekbLviQ5KBtM+mXEk9AvJiWIKkCXfkZ43NBJaGbS8mBxAFRclS
QPotDp7VbzugpaQmrzD8AKq9aDpIbr1+LpQunG03L1cd/SCrrFG+kmxvndAhEhzJ
wJSQoUBdP/6z4pHkEQs0fNXolW1lIpewlr0Xd/1tc0J84qLdELGL+m2S5i8f0w87
x5roc1advozQpcx8IeW7cLKmxBxQQJKPKtk/IkwDfMjLtUNm6FpzvRVph+sluwxd
DbjpeTnaEVrX1KsRQNFe5MOnVjNB8ZeWCvk2KN5w5Q1AwPEgbKh7gF3QEkXgJRvt
vBiLGtjUkHEvuGtXJM9HHT3haJ1Ae6+Dwer9E5KhjZPJl4S2VtdKPwuQuJC3xvzs
h5eEsuCLLD4JU4+cLGs2ehQSYogPeaufVL9Zzd0KUmXfaBGKKkimsXRkDnseBJhe
wywX4sKL7wybIwL5KTibVYmcHzBMrbxX/63+tyGoiACcQdX+i7UBDaeHiGlnaXqb
k1HnXpSHZSGVcTvFfi1fd2iR7750ZUk7+fF1ADMs6NF/nnNzQiwBE9VbM3kG/NsC
YGn7l6K5vXe2fXIpTi6H2kl3R7g4FO92qkU6QuQJcu0q1HngcNtoo2Vltmi484xA
do51QyD4Z5g9B+Y3tiaDjSHLrUKOCLK2SatRQmXwyyaKDOTmIonJ/gPP2UsXx+Lc
wOGlm2EHPTg14DHEvCxF/pTq1jLJ1830aqunNM+ze9K2tZw/X70J5LQNMPn80rt1
m39Hc16duTqJ7Qf77FK2zrRC0U+I48OOOqyjYk+miDF9chS+qmY42cNJ+jAjzJdJ
KgJwG2J80ak7eaXp6fCke9/E1ot6RL+w+cs2mgObAU08vR9ICSgxPuFMMqufIU5I
jNRx5z+0NppZ12j0j7W1ABTtUjHQsBpTciKGbFcrRmESKd8/gJuCuBJS7DKLmLJM
yA4DdLPVbGYlEzM2E1mcWOh43QMJSJvW9+HexRo7WE8zMKEQO4uwY4oPx8W8u+Sj
HzEGdfUfvODuMD0O7RdyvChf5dh7ij2WLpjiJnL3wgzXE8msOFo0wJXB9ygShV6+
Obq3oN4gLSafGL4F6xsw+9Wibzb6k5T78F8WjICzM9NgH+g7kHJjTadlaiGjByei
Cc87ocBosvMBRbZ06rnCeiyfIXMxCVznez6AfdTnZTtEkYLKXTGRhmVOD09wqr+N
I88/7hu+JdsTF2n82I8Aad5Pl6scvT04KRTA13r1MwqA2UcQ9dTgxJiTcXef71WK
gFLDyO3Kv5GZoELdBLc6lsnJriZPdBFPtJYCpVUwPj6iEeTjWB5Id0CJ39YXMaSB
YO/6kwnfZE+PzcLCHNKnvChURgeO/6GnsKyPoqTkzooriuByPp7gf2PyjkKSb1XK
VNnCCAyrYHRQYW6ElCuFvhL0i3hXfYYZyuGohGHR/nuSBl7KnmKYyozpM4xwZ9HW
QLamt+XW/y+oPwyO8jvL7pe190j2ClyW/7fdke9DP+fYQOABPEkycxskFiW+TP99
+TzbKdKs/lJTMZvTm0eBDbY3xBQVZTbP3t3LlgFjJ5hW3HoGhgnYP2XgcW8nhjX8
izBkYjVtsFeE3FqcSynx+JzTLgtmaV3xvV6LCl5LJwQuYSX5Eui2XuVZig1/qxmT
ofOzrSu3MmKLqXDmtlKu1AG881HEAEOC1nKr7VvhE+K9kPm5fO2BNFCltY09xNoW
pJ8BkCsQmDEO2YQRP8Xla16S5c3DE6gCKcmw+c2IMZKWMEmDoSX8J7sgNsXcZHoA
g7+zU7aAl1eCAr+Bznjnli2pFdpivLbLjmMtZherbPOqerVTCQsixH84RGfAAq8O
Q/wFCp2mQtbGJ9JkWOlatB4V47SQbYi8qN7MicsZs8Btec/edS8RLCkYRCVdvhxk
csXE1Q3886yTrc4U662i7GczXKpd4RIBlZ/zURmFb8UxeoXeiYgkAyGnzIj2VoL2
7WGK4eu7sVAWx+zk9qMywhA3dLnvx+ungxzi74scCW+DevIyo+ZETzrfz0QNuNFm
RoKyhCSGNEFogq2nKibIiwxdKEAVA1CMdhe2nB92D2oKwwGmuwpMmG1cHLiWZ9uh
/AdQFkaNrD4ThitmZMRBhoz3MxFfExOCXDsSni6ZPrqqZ3tDupMV6XiQN7/a0JUW
q10bLoYB9GObRctAk5bc+nN3Lq7MEl9w0U2Dfp0dxPqvgWeVCRzmyO/p9ArHLekO
dWKuIgMj7wF0MCmGM6y3a9HINkvXmveEbSSggyXONJPjVTp9arqxArRvYKl4P/kJ
xIVP5FQ++9m+Ga05zE7XgOtqGwJxvpqf58vjdGoqD+ksDbHJ5FACFSUXqxEUcdc6
plzDyzKB4RiyP1R+j7Xf9Jpvpe3l2MNEfjOGBFMwCtUAmo0RQtZ8MTEHLzEf+jqs
0lEzcT3AjBQONeFFsaLP9Wz3tsBW4RoT25yyIBY1XFen5V3c+vO3QsnC4sdGMnjM
76kDgAW3CRw01Rk+VdeXWB+U2ahkhVs/9b2pULqv+ZhqURxm1iiIScCffLHJWX5g
nYBOeLyWiKHTR21hTtJ2NA6yO13hTRpbwnShgo9x42vxy0uD+iIaPElNm3NshYTv
X/xcZjiJpTxtYSkX9QIYsxN/qJjM0BQTXD2AXfIFB808rbjQmoHuXogEfkTgEAYr
aM42mscoFGX+uleA2El0M1qVHafpg43A3QEx9Zmg6JbytGio5ZxnZUZE1fsvpsaF
j/jX0GWBtMCtjkkh/2/2QOBDGFz9suk8Evw/BSpPpy0YOhpIiuqky68vJiYItcyK
gha5akiv+WQ2wePEpnSxThXIL0Qs1Kj3U/4EV4bR48qUS8vRIEmcsS49PeVK1+up
2yH45lkSkU41KcKoYrJWaWiQDCbAqFSlgl8GxLeDATa3Aql2cGr104ci4I4dNk/w
BDCz5zSKeqbKdoaJ9GC9qvZHkjavNXnOEmJA/019CH9Jj5I+vl5nH66B7hg/8M9e
ey+6ZBLF3Sdzq8x2tdQRbtvWAeBt1EQSn9ovSDo2Dy0K9xEFZoKJmEDqzi02WyGW
+SB3E3uAviOCudzD258EcoiZHFVAxb3VQZ7w4Bp80umzrREiNTM+kvvGGEGVbPlV
S9qBeFPJp0/YRX9YRTDgY3ZaHrPLQEaiD7GYQySDiy6DU2z9tfVJXEJW+d1hvupC
8mhCAgSENNHfWjA64vNNP+ksk9/wW2385YfEr5NQKTpT7qzfHZTb3n0W4MGfcI2Q
3E+vBHXhBHByd1Hh1K2V/YyMa37hVXQ9hQcR+vp2W0xwYpuBbAkF9tFKuTPAJ2VG
lLSw9dQMM667Z19EDJIPV/SXYfdiHnpbV98QlhytiAfov86Ij8/ShKgKjlbtfa+/
udRAiPP6P031qfliQPG249hR92e1fVyrKMuf8uyw384F92uPRl0ozS/vySwmaWxB
AephdItFYss/Jw9nluHUIS7rbvkMZuqlnptTXFHy2iTxeKjAbgnp+4JQf6KBLzf2
T+gt2V7YTQ8fk6VuiSfrBLvOAt9d5YBOpanPTikW7Ui8nKP1dX3YuXqmhcXh5ETW
Hhn7iQdpBWbRx6xRKJIJsUJJa9kEfFNtc9nNBiEhACjPypJH+mB/D/qZ0SYOm0Va
i/wNUMMACF2zb88J/mHwY8pALc/+ZD6LOFqOkNbqTSBZ5waNLLw/2sKHA9k4IKt0
HOnePuQb+YAZsxFCb3/vaLwiiunQeNhqDnlGRhSZfObAm+gYwcCYQ4swGSuQkWLB
TXtZm2WwsPrD3u9Rm91M52w8aX4RQX42cXtHoVMXfQ9y5TujF0VdO14FPUBKyOO8
XOqmhhQkrM4RRlS+FZHJBAabhdNWsmUBs31a3vcG22U8QZDpThDUl+gGqTDrBIw8
gK59YZ8LGdmmp3doxZPnpYe1/7gz0qYEAr6TxgiHnZBngtoG3jScASU8kumJQwAH
HMTPJpQ6nnnuDctNaLYdIhHDb/4l9tTazQNElShHew1bSKd/X7bSCU354MMM9tKF
TaNKdmivizG2U1n1693EqirakvGwUSU82t9Wo93QpJP58zmnZ3k2pNUkM5tvdY0+
ZUDtwZt8R56aLYpEcds+G4BXw6TK/gHugAYjkQruKnZjn6REsHTZwu+5LglcSLOe
7hCVGJmh87jBAJ7ZzaSI76GuFdc1hyvvxHRx2M8hodkWovHFcrdjcWJCCVI9X0MI
ljYzK6RqYwTaLNXyoapwLItRUmTAsZJMDQpk+5ifPNOzr6nibnayhCsdcaaqINd3
+CcKk7bXLvrb4gVggOHCWVEOEaMDmvs6ScToIa2zMCGLtnb8oc/2HUl1YfjFDuud
gn+Wtug0K4S5nsepGrwo7EnzKywb8XlotAyrJ1JfjD1FKZe3zZ1xmQ50KjT9YWr2
PckAuFnoI3OeRILy+JQPFl9qbuhKiZKZPrJie0R/nX4j67Bx05sh10QjLPK3n+BT
bpXmbAuonwPjMpHGIagUS9RBW+RUfsppxTwzcqhppam+F3R/okWHO9wA1Ygefzam
5gu+cHP5f7Zxi2DLd37yJ4ZA4UB1QfBVs0SnWlAH8Al8ExVM9UYvuAbo7f+fUVdr
2ovm0hW3DFaa9dliiyZGG6E3QwN4m0USAZLO3WCc4eXvAnKB10FW1Ly9NSE6Fs9T
K3fdoKE+kZ5Z5FTm5hCwb6LybaUlQjqz/4ItE6SIqs3XrXQDFgATwwR/N96maVuv
8eY3n11lBXWUfzYtHFlhW8gNEnp7qe9/sO1fBZio7A/kvI+gAqIf9AoZ7eH+/ZVF
OsTo/Z4GZ2MYJD4c9aYexK79aERKfotSF1q1BHTBdOZyPH6FBv3uT3VvZ2rIt+SW
gmkktbcGbz0Xed8E4MivwQ1bmLEpx+JDK0f7laNZH0+E2mkvAgnE4A1Uc4VMzybg
9Bocb7W8DVAxTkOVgd11GL4gK8Sb1V/OMdTg16JqWzGh4k+CfyQ+54MGdkDqMXG2
y6CbZgvi85P0WkFUVohWSrgBVTlkDK4te1uLlDvHBBcCU9V7eEayfvtY6mq45tS7
956cWHyEiPL/wfIWxImCxSDSAM4x9l4vb6OKXnzaCMwaSB4PxaQmpgQnW9E5TfmO
AKDD08D+BD9an6/AMCBJH9N2d1ktgJ4Oi2R9HazGRamB0DjSJnL4ZNLk2+pP3mTj
hPinwX92dCPjB7k1wT7NjlnjZZ7d4g8AakB87G7Wov0OdQcCXJRZgydApW3oO/Hx
nbNTd5VxglEOucsthMAis0fVwjdzUDFRmLXYMt1uE2CDavt7ldothGULwt3fgwbh
bn+5mLPg8xocsoOhF8fTt29cug6VN+77x93euXzN/ICwQ9ElDUEZ88T62pLOVSWc
yzw+53bnXOzY6GQYtiloixE1NjSYVnOIfBLIRQ3Ao0NLyHhnRlhtForIjS0OKIZn
F8MrZm084q16aXVCcKOMRuZz0tg3hkz7FZMyL79YnYe2eIMOAlaPW2os/7nV7o8t
iXKbOueNCepQG7i1jdgxu0lsVg1w1oq7GGHh9UBnCKItnJ4q7/CfDJ6iw3PseNve
ygx0Xa6RMbSbnNJaOvNdoEFLl+3f2Y5znkWEJpMVhz79pPTQEsDvWgGH5FwYBMB3
wcHpzpTySOuz0z9lQ/QTJewZIu4ydz+gl2qq8k/+MCRV2jGyVZ5Y+kl062lU0+4H
SJHRF/Q+0jGbQ0Plw2XCuQG6BT8h9eZ+ZBgbMS6vu1l8Ys6Q3TTRp7N73A/zb6Pd
XrIIx4n63jaRJ+4M6lJa3IPoR5NbMR8HSomSuZUo+alNVnLtlL+W9DP2olQbkG4L
08Jl7KRH57xn5LMbhckx9kSepGO90VaeWY798Q8qcX9SZ77FjEze1FviRuNN5K9t
RjCB78nFscBnJQYdWxD+76YMIvqxIeI/Vcz4fqGnm+imhuJt2bgaIghaALr6lVM9
Z9OPPQpsdB9osldNyiZNIPMYEZqtlACYHsiTatvU3go8Q59LMWmbpcOOPhCPBXRD
Hkj99v+QeH6/lbM9wEFWR89ATGaacz7ltmuxN9OGJWZV2ld2BmLReTzQ/FfOF5tY
86nLobqrUSq5pnPV0da5/ENetiBAGZb0J7WUAPbhiiZ7vzZ+kY/F8V9bLwp0JmZ+
Mqm/Hu/gN9EzULU1en1PmW+IEgycZtIINypzeYjBlX+rA9uC4+9qxzkM5xhaeFl0
ioeq5b2595VjICkLOe4tHXowqXUPYfj14THTQT9mXcY7YJU60eLZKQqeZNhOfg8s
w0gtn+zSyxQpEbO+RFdFK15hwbN4rELuMi827JhQTP70nilU7/cPlXghmaz7eRIz
2+3qZq/a2ML4v4ZNuFCsjn2XxySwuQjupPEzbDR5/OYSTXOkxrZri8xkrtiar35k
1K++EdUAnEwcMaxT3mW/FplQEMCA4H6mcwlNlsmqC0clX1RQmrZixMmNns5lGbBM
MaYIV9eT7Un5CyzzNNJbkuei9lBmL2rSyshtlld5P1RAPUeQSjTrEi9mjqnqiPrP
0TxBaBz3SPcUr4LHrBH9tAkG2JSLYffoMqtosbIxyvxTXfg1DDdS51fp8QBG9Mh4
OHGXyr/REZ709V1SGDooiZNJGwyy3WjjwHy7m/3iAHrZohHGzOuuhhXCTDEDk73C
bKQm9VO2NlzxIzj3HTeJmIbz+WeUES52WsezdNE+M8hVa3ZZcpt661NrEafHE30y
R1ubnI2krec4kM10OMmKJYec3ucGNT4gwGcNz5uazQ8snaBgOeAg9ghVdbZm+B4d
xg+upDBL5O0OopYGrCKKn5/EpORbH45JqqT0HvqDdLY0CqTMwqTbeCVo1aYGajY8
ohkyaOC/kzviZqPorY9N0KfUHyzUETRaizeZZGsoBWJgVoevKV9HkkrGFukXxeo6
TJweUJcHJEv7APF/za1JjtR+RvTFG0cCqzsNOBWZn1CpVJRj6huHBjXxNBaXlMJs
7P0BPIy9AT0okH244is1RFgpcpTCAcM8+G11NFckhL0HCBCfthao1V1ugyDEWb/h
1k6WkmkPXYlLKivYenExaTprOgDxtu8CTVYzM0J5fsCCCrPFibNnrHV0Ft3LVWoI
4d8FfwFTaX92KgXMwVGaiJU9apqeyUyFb5qyiAQ4ljlzKl6JLcahGi47S4EwP0ET
CajqWjTn9SDq42zscjRbbrd7SMgaM6YpnIUQ4c4efgwrhRvjjL41zCpJ0CkBJLoz
Zdhbp8upEl2tqF2saES4TXWZ62ov2+2GqwVVwhi7kXVx5Ti8yUJ1UoxT7wXhyA2g
lEqbHVy4SYSVpXbLLgDgb05OPP+YdPrUTLWrevyQFoyZVPQKbuPKlnp884z7ycT9
dCNaR3L3cmOQbG75CVru7Tt2iSIX90hbohusnCVZCm2r4khZLLqq5AeChL4lzASH
uxhYCXU57rbijYvsje7QmoNnP6cndkdeXu5hF127VKneYagFVWI29WTz69VwVIg+
SEemhrJYTVvaQAPw+w++f2t5Q3UzbQ44WTp1KN0+8o4QdQ8CaJ3v/4EvMpu2xNtV
gEHfxFLG09KJ60vice26pDaa7wSHvAiOOixbxj4EU8fTFEUz1bkN7RO7Mnbu6HIx
JxFCt/aUj2SzFabzwd53s9QCtMcAnZmyReQ6GvIJdDP98pM2BhvUyBBQ2Zye3FpO
kjTSNJpZoqnU87iuwR9QDxMxpnzuzcyjZ6gAt1aItMB7++OtxvnAm1xQwYtzp8U9
na84iKRRYKj4oenfVbiVG1EadRDI4ScRk7dO/h6vT3p4AmCyVvsvAmR/T7x0bmPH
48WCBa/LcxvC5uUiqAaWHNOCVrNdrE+PD/44+s22LP9TqFCquOxPoW6bVPUZnlkK
3OcwhhRgvGkbV4pKWpI5c/+ouk8/f7Dz4oSF9EnoEyFNwNZ3MqyOBLX4hMBFPa4C
IYNTySa/ew6pzpo1jN7/I9Mhw+9b/6E/C0dECT/YOsFffUSJZzX0q08oFlCRB7bZ
YbxLbOyocftmrTyiQy/69tYNYC18XlSzjSROnJA7xTFYCYsAJGRVSlzX9F/SlaU4
arSEQYOI9J76XM2ESVasRMmWUtqqSA3cUVFOUo/yt6AxgS93/f1O91276GsOzqfJ
qtCxQtHRdo5IVeCFqZVvs90sa6nN94JkXZyI83vPmZzLPJqhvB/F3IqG8DTPTFMU
QS9HtKK4+UobGg9X8i64Qmh4eeUzqC71YmTYM6ED3JibaA7xSPXSesUSM5I1qPpV
Ufr6PpG2CI03snwVTsU5MCVd8+53x4dP8WTFEUN3UQcLvIA4+CO7BEkqjHfftEgB
0CZTjj7PqAdhbqGvCT0po4yTaYbSYDRZppHphHdrCCE9CZ5GDZ1eeUF2krCjmTz2
UL1YTu2U6rkUKZWMtGKcV55IKYeSVwSEBxM4V6vIyzt4fJ8v+mr3vKoZKpoCzCER
500LT/cseNkkr4PGK7ZfrLhwqYKX5ZgkAYCASC+JYcgRu7TnboL6d2cntCRIAcVa
CJ9HMa7JkrDQUOI7JEoZkaqaTJIcTacLZybegId2b8RhgmeE1w467kf+mN9QsZ6d
ZwEppzRX3DkR9jt3b7IAEDrcAaGKzP51s5I4rHYhMuorxrWOlfpQgqpgv+IlQvfe
3CFvXA2YdYfPAbKQn8yy1ENjCljpPDFZdw/90Tz1YYHQPe8FTUeOEb2TK5a5gJwP
e7jUcZdcv8HCRxOnwif9gwJXQzdZGFfHX0tlJgFayxZsY0bYUJlYNOLokX+zUkZr
ibXG4JSUOOcLnxafDJlDt5243mrrBmHHZiFg+865bu/uEL0fKwFm7kta5FYm5Dqd
K4LqND4K59m8JREjJUJS9ZjBUmR9ha4zYgajI5DRe0BPauBP7cIYcoSYyuI2/TkB
vkwHjFfOLbfH6bFV4dZpyPTyPGAlYVgjSkNl7PYwvsa39yU+EoEmyefh3x5eG/Xr
2Tsgw3alw21FUfbtvESULXcRPklTmWwqeQInLyVZw9qVI8r4w51bLXCuqi6eMcIo
LA53tGJu9OoB40teFc2uj+dB4abpI4bJuvq8VkIWq7Gh00ZyJPySGfqIpTUTL7TN
EIDylOm91iVGCBssd36T2G3ZWmzgvijYKI53BU06QJu53N5fv8zAx1TR6SCoRhNQ
doSPfU7DXIzYWyQwkYl51dVsm9Yur6n+swnh/cS815Inkj4urqXeCedV0eiEXFtK
ZBhDD5zsHCyg8MR3htiwyTgEU0XEVPdMm8TJYnxfu5ethZTWgeabc8Ko/uMY8zmz
7maJMhSaZr7R7Qitbucc/W/340M3E1qCCuuv1Us/ef+Ai9rlrSPpvOq++wflikz/
gHDkk6QxZxyrPd1L7xfMqlHCwVPe4aI6t/kvjmVse7Q92H+e6HGd85ENZXX6tpV/
kbjRgBG4Iv2ntM+Z1EWUR3q9AduPb/Z6zO8POMdgLyBoiqt0h5z8CEJYveuiAaw/
nOX0h7a+d7hOF2AKlvBA+5QGINb8WFbZ8Mz0OLuj+aIOCqjD0XJa7M4tW7E7nI6g
00ZwUhRR1isY9KgNCRFQTc/qsJxO1g3cNG+45Izh43VVhGMapJbDhyBfC/jIpaOW
7L4cIQPjHRN5wnc7EEUDPq3IqUuWO5XBozBhSe4h3+BK6WuI1CfdMJE++FXO/vba
zo5P51nwWJHhVYRxY9E8ptDnX7Rs0p4qdp3UACQPHEg9f9f0ddUNorOTc43qprsM
sEtQgjnfmM493znRjOQYtVuFqvkzVnF3v5Xe4yRkGgMkUKUoy57RtXdrj8Ajusol
/YAnzRgTXFVjzgiQ4xhA2bFjbaJOSJEDwLlZHx3jBx4mLPrpz5j/DGoSILsyeH2p
GSCy/obhiufcqNo8CfrrvVBAYHzrNCpS3Ac5nb5pKA/cZEcuOkBur3vaTEsCXmWz
OVxwGCn4hYYkpk4/VB6kFlTrGunfVd6yRC73Nj2omBaKNcrfDUW6cRec7NUIUvcZ
2K8HcCen6m+eyhl38PwolIr092jrQGm3rgawPlrKK8oXxOobIFxuNyKNEviDZCZf
P1x/OEq6+68s3MwWy7VDcDWPwzclZ0B23Ogduw2dMzbUtNbRgNMsoL5gBxHhwv1o
IqiWTF2mqfEy0GDohu+43dPrdBmrnCaxXTN0S4SiU+kbnyGeSeY36mOzhWtLxwrI
CFIhedUfWFqqOtjYYOhq9WoiY+Waa2YkiqCnyST+nwHwKZLqcZtEGHWGQDP8a9vX
SR/z5coGy5MR7CGiwYsP99HQ7tV57QFKc1Uvha5qilCL2Bwhs2nf3VAlmii8ZsWq
Up9nYv55uJ44C++eDQpa5DIXAO72JY53EYNMfgVHBtnjuG5567bBhBEmARhr3+B1
cIqqdoO8P2nXj9AOPkY8/CW/YnFyX9p8UU6B4JJhhKmKgBk0PPgmi6aeTYPnVKTK
xIH3povz6HYmUF/Mditb8qBOK091IVE0kTsYw7AUo6YS4HjvII23AayF9mJppV3n
k2ieiqya34hNPkuxoda4UqXeNMIqxOi/Q2BWrHK1BrSkxzGpBFMXkV+aK+nDHXBc
TD/eCosfJNwQidGdsXiSE3CzOkBRAWKgMkQVVe/Is7pljWmHUZnps850lIlxnNNK
E0S91IyKPiWJcVWhqmgBGa5CJXW7gKEAiIfEWRBsl1a5cm/Aw2fNeWBELuxf9ki/
4ttci9NekpkXhVW0MLbokN49S07Bz71WaUK9iA7jnXrPtu0jKBiZramG8o6vAzsA
d3Xgc5ROWx5X+7Vi+5by/w686IgqoGsY5jqYDLZ+vNETE4UgAK4gH0igXBpn/cZi
GuZOVbv9KNKxkVkPC3Qx+9al2abBvSDQDdqhUUDqnEwxNfX/jX6Hm16XjHT+mBNl
PPrSMhbxW+NFnHtz81Wt3M4RbrIL4sJPNgF+rS/OhamKw/B8m1JYGAeR+VRnCIJl
CdHDcznt1pI7b0gBjBqCj+kx3cCYUdcCLMtJ3BHCskPpHJPUDRqKMeLnCQj5RULi
9OjHR1p/PZjv3DPBItxzBh7dAKfc5zG/X1EEVCN+fXuZoFNp+3hCR5N89L9MSip1
j02/slylIYRpOfVclxeMdtjzIScuZoOSxpOdD9CiHxGylapXTbIMq1Oci0JDmCmh
gswAyeg/EveTrQdctYmL78xKdyzlXsoHdgXzaeBbvqiv7ySHGLBwWPHBS/cGuz+V
7OzauOl1nrdtI9bP4dByK96vmIgVqTIkPRl2VfWd2sLBZwbKlt6iEPhuUB7YNYvT
NaIahmjfDFh9X+8nlUzofvZ8fIrReDJGJRuActWhdZRafoULU/lULkE5muixJ1mN
1usHNZwHi+tZLW6xePTky7GRAhFajIbSznMUtZZYaiMQFnCnaJH9lTmDAvuFoG75
yxDPNU4l7iW5qOvKMNaun+vVxkxeSm7pm7jB6r2e5n7JY14sMw04Ja2fz+/O8ErH
TvzRM+FycsPWKqxIrAbm3W35jGPlgiZoiyuAjbSLfOZRTEYMC2JsDBkKyhKRxAty
h74aD1MoBVFgVSlW1JPMZoWTvx7urGrWg4XCxWJSzpMr/yHqSbrfzGGOfmP+FZHc
lpI0KYcvv9pUnNCoxJzKwCDQdG/thBGvy5aXsucLZEDNWJCDsPOHnPvbsr+5hU8F
cKfUoEoWiWGu5xFFyA63SPlRUMWKSGf5aGu7/rRXX5jZEG/5KSG41xuEjmulADwR
aeHbKuEmq8YwBETsDVlQCMwkR6oPht1NzG2rjWRrNHYjQruyRFJA1TVOfQTBWk+I
Q+SQfxrGRBlME/GZpEuA0mAEvs1YkQj5dUnTilPN24tYJ6I01i90Nsukl7RJsOeR
BMA8hasGw36Fp7CLZQYQ9RgCOeuRtDY2MZc34iobtXrxKg9f3i3KO1Kf2RJbJXLH
DuXhuGYIWUL7uRCLn2cWotc9JgI1hfxJHFpxVFSKAGE5nfstNbF5ff/OyG2I+33n
f9faXXrgeefPanZXOApqMOgW/lE3qg3hJBdjkRNoJ7emA/j3eErXBEjDS6JTHRMW
VzxK7iLPDlELGMtFp3SaxV11Cf18j/Z9Tcrfu58Rs4jyQO4lny7/6QGMS47wfyfU
xjDdkymzUfxwRND757LyKhxknTW+a/BiqV8rGg4ehjejJVU2DeEu+rca/D8r/yKe
izcajn+qt2bsHfHgIbiqt/ogpdgl5gXe6FCYQJ1iTDkD7aQtptyPC+lC5CEcfWvI
k27+bwV5ZJa5u2RpkzbhKwQw6/q2NTkgvqMIBjPnJ5iz0XNG8Hrw4l6sRNf0JGaa
4YwYF15w77MMaBKkAvY7gnBEYjiie3aqqDAxp3nyoyFAtk3S1uF3FCHFIUJZ/4Ec
MMvJPy6mRH0WGY6JSsDF3JBBzYwVXkOb/wChikGT3CUMXAUoY1V/+xDmbfizyb75
YI8DBpACAPRedb13SufcRppiSgfBTQQezwyopFy1deECnhiIM4fwALutRLDNx1wq
Q4wx9xnJjyMqbPGc/fA/LMm1Ua9maErRHXbIdKHzoQ3cjTqfcUBm2mQ/R5T4JNmj
YkwD1BGuOceuCA4DX0hXrge52XFqaesTuziKtDVDt0pQrhyRFxWma5K6OCHsnNRA
CIybutMRxV1wDCVTpG7YKDC2QKojUu/uvSUwsh4RyYnxoOkBPUDuoLvB+qMgBCeh
P+PqJJSQ4KKZ01s3KXq6WpTNYqI1dgR3awfE7qGDkH3tGiU3H0krAlu639HOXwFc
NvvuThU/hZTxyOP7ETV9z2BYvUfJqGqmGcfpeFThrVoikX3R2xYl40veI/0A9wVE
qu3PR9D6UxVpzeJD3mXhzVfP9Lzl78nqaoJblvw0qHpIXeGUj/xpvb4l0aDQiVfN
SuYtp3MrzWQnqP6O67QKGeijbmoJ11DcJUmDhtAMFSuZ5fARpWqe+/fGnOAq2kaO
lsSrW76t7JPV79uATAp587koGv6j63p4l22etym/h4/hdCHlfiz386eLkW6dUbGS
hf40MxAJEfnXHzGVv7l6WISjmegn15gD+S1EHWV0tjSLTUrOXgSLtOPf2/KVtuvo
Nb01xLzuXJAnttFtnOcupyhJ1HKknz8sUgdo6UNXeTEN9MZUOFEnETNG6NBYU7N+
vaqk49cLhs1gH00N7S2J9eW2PjBcW/SYjECbkikk8Ldem8YY40kKEgCcIH9dYE5K
rE5+wXxp62D4D4cogl6mdapH8rLK4MUTFtUe6xMmo3s2yzHUj6RLCq6uoXAhnNcv
ABVHErHmPdvnYj3ml/AdXXW8vr4KdtiBQHXiPNy/ilc/KICljhzqZXCeH707GkV0
71mqfQp4Z0W2A4RexMKQ4mvusfLmYHVieRS/v3yeIqbcwB5yK+35/ouOq+Nwle64
Bb4LTOJJHNsmhMv0dp51A/qq0ol1pGCUEfegPFQIh+eDivhzbxYj1gOjLSNWuY18
pAGBQshOMeY/lrg92zMIdr8brJoAj6c5CatNiU4QWXBunyxMebKwVd90zqFNPruG
tezK4tEZ4MogVMCpayXkwSXXrd/vkwZxoQHDBDdlRDo1VnrSEccMNCJJRQ4PXk6D
/vHduSo0la0YEfGViuc8OzBCN6wT4tfxjTWWraP1tTY+22/BI09tRMDy6btJRAi9
eq2Eul89Q9cRIIL8/sX8xOdqTF70YmcGwUAPFqLP8WaytCERqzgbKWqxVRNmc74v
cQ5ut5wq0oe+pZMxFLbZZuLFK+r9sFMFdzuDIexJnKFLVhUqgmXThMfpfr+tnw/C
ZGnVGwYc6VxekwWNv1eFTfdysEp4VK0jkzsD1K+sZCaQ/NrgDr3ws+QvRmAnWkhK
j8yAB/vDwu0doFuFFaAkIAqrhWxD2nA006bW6VSOonC0pnvEwLkqxCU8xCk06eYh
J5YgJb/WnMMopZW0BNSN2zl3DNQQoAWs3zw7eUzYgia78twsvo1RIAeXOo7/buxB
yyxDPtsmzYaxAtVOXiVokclDCHzSYt9ox6ZIFtJxWex4pLXo7X0Pm4AxsRGZl/st
U0Sij6oGo02Q61aPtb3GxQDkLzJ5kfXYKrlHawIBRazLYvwa9jKeyWkNBidLR8Na
7qKCAYwHYhAisK3/XGCUgpKG7EeOUPAkolt6r1Sd4T8kdac0foj5hwsEeVfx36kn
iKRr8Ea5zW3uZFJGKEG/WKksR/b3OM7Eue++nKa6vl2kGePA+/Vp60QFP8AuOLGR
eK2o1efOHvIADT+f873B820qoLSFsfCzVHEp1uSzLyxRyIOT+2oEUPgNdZ+QQEev
Rc0y7WTaLEdVuvfO2U73KFtU8QP67Hr9PFxYsOSwhJ1JTzpGYoEUcSEFFnCNcCtJ
q1WO98nHiTyCXExE3P55FvH+mInYnjE8PzDvMvKw1NMMEegx96q40t3wGgnA+4gc
DnVn5NvnhLg+/jIUEyPJlZUMo8NknRI73eqSa3n0u6sMRJdLi7Avv+WifV01sfVX
jwPgJR+eKDEZ4LblfEanN/XlMgLglpStNeuX086Ca88Jh7cfn5Ln6dC1W2O4XU7+
nK5YVx6DXTbCL9E3QfwOyiAnw2IY+sRpPsKIav7OzukXzB32XyacDYTjOXU2VcQy
cuWlZeWXgwj7o4r/tDFb+YFDhJ2W2CHbD3wlWq8hZ2Hs0SczW42bBkOgBEcAdx1M
1WbjCLKi6y/PTvBcFPc96WDRfDTsZbMQQpFGA1Y/cZcJ9TFPVLiwUm9sb4btX2Fu
hv+nm12mysQzxhp7yctIwCxM2GrUdgdeTREOs7qIQoBQiCP/nITHPmO/x5+AnHES
s/hjLUH9XItBUSihygLVO5pMR90E8aC3orkrKrs7rq2S8I1W1kNZNpGwVwV+EObm
pMUKw5ZWqiai4KPFprfcCQ0YZss3nPJqfc+iaJCa7pjG6VxK9onGhhX8r5JEAiMT
y3msM1tn9o3jzqAC5aPsezIXRy6qI98ObMb2L8vzJCBCTGQd52sTFyvYjyZz5Z97
e8IYQz32WsV4g2bdHiQDOFbzr38hABP+Fu+jnjw5yvcaOnUUIWn64h/I5bTQrZQU
NnNupfwEq6+OtxwsdB1IR0LoN1CFtMimj0cCfmZ5bnPNDGWM0Wg4O9/wxYFeIRGV
UAjjSeG0/fN6MEWocpdKKIx3btpipynDW/V5Nl1Ls0KRmUHQ/FOJP6GnlO3Zh3NH
WT6fX7VHhHDLLHoZORxzqEo9fvc8y9nXG1rfKKUuAP9kx2Wv/G5+zrKG4bsanWQU
G4ZUy0NtaGJ2ZbDf6fZ53lXOSq0rCbX5kPD/yOABF3T3oM9ef93h/QzZg6zYO067
6CuOfK0jSi7TCtHJyP/Yrba7oG4GT3a+DIqyoJfYDjvy4/AA0eULkJDFX613KgRH
kVWIGkQBcLfMdZz95PeC8nJdt8oMSwwxIa5cmEzk1OfYy5mDKFm1bTTqEfxQdQX2
RI1He7WW/Ck30nGPKh9I5ELPqxhJGcumqUuCY108EOjk7Q2LuM0GkUXi78lynmHp
q3cSoTFyebAVOwPiIPGdTz1UUlfydWthrOnJQhWOLmi8djjeOz/v4lFNw0NuXqK7
e83RnrBZ0R6DeKdWzsd2sq7qNqPoVimOMwyRUAWj1fNzt/iHJ9pSF1OtxXeuBEFo
ZRzFarHWDBVYmVJzUOqaJbon2FmJSX2tubcFvOx6Veog4aX+Go4dYq0mauu5A+Hg
6RPF+JJ+4lR+E63ctAiXo3VaDN9fFVrGkzXV/fiO0QAlZ2C9oEn1am9p7AYVt9CN
gUgf7SYfX3KfTLhWG/agFhNT/3/Cj7bsMb454R2nDFb5oVePkcwfBDyieON6uPcV
hmchRqLhrVcjND4Wfhgbql+Y2HnaNiAG2F5kqvCNHGFbdkRqB9B6inbzPQ4jdgFv
746v90kXB3w3lF7zwRBYMOun/m/kiuvkFeU2LxyPma28dlCmu4CzcUvyVM9/U8Hb
Z3pCzYRSkSOJedwMnTxj01va68BlMJXsx8LdjP6Rq3NAbwUfy9jLZPk/EyuxSkWB
CS6dAXGyLHpAhYnllgr6puDySEqKh5oGxIAzkQYiNsuf4rAcYMdk4XWhwBzDEsUQ
n2sVeMvhVCT4TqBJsXzOvKUM48YUQPWCVlr6L+enj7OJ7q1ZV+0LC1tCWAG4OBtH
2BgnJKgHzHAaX+kzXz9h4ZvA3yCl49fKVcEJb8z0YsfzqOiPdBUSYTw3cjFH2+Pa
/5ewagE0UBkSXHCjmUDQg5EF7LJFzy+k6gF1f3iAYq91LsZDvKcyGTY3pEj5v+hu
KZBvGR94rxQq0ARh4foE+yDGOXScbKEDYZFYEIipdJBpBphdSL0yJqGQ7PDY9un6
FU55Wx4aVmjRqAPt6c3gxjZwe5v8qQdkKVoBRW+yTYfdcpIHAJ75m6bA07rV4hRL
39J1Giql2edFfJe0wZxq8VWA8+yWEWlTSW0A901F3gqHAlQi0zEtyQ9zBY+lsE7a
3IPFmsgd5JNo/DNmZ2NIkHaZHfZJ/159z5GGDonQFZ1GFgGlBQ4jBVEb0oCHEKKX
sPFg6XeBk25852lxkRfeJCIqlvwulWh0uqyfZWZuYAloUSYQiz2VaheQSWf2i0hn
M3wKSiNDPzAZqLvgORjF6Sop3zrkTZ9CnUvGLk8wWdPUL6u7MzFHxzU8NGWuAPkK
eY1CiuXc+NZXOyoEAZWi9Yv+ErB69wu7168MZVtZMCT8mb/CqmbF68rErnWSyKN8
0NMEp32yIo7XcnEiTavkGCc2oM8l7TwhZbtUHsIUhCLLmiFmaXa0jApeEfvQuOLU
o7FiqkImkf+GQ9rU1GdSbhCeooSHBNbqzuGTSv5cuveiPNSPQVSIz/rhg1McoYA0
f/TtaMMCsAbsiof39RTk3/SuBobqq/Dj2KtHltAIDhiebfJMgeW9gWlapNRuP1gN
F9WOB2db5XacTRp7nx9WpmLS8z/185CLXzsShLZZp7BFbf3dUwH7X+6Chf7vi5Wr
D2ytOnssUNd3qTdFebfbnEP7wYulvx1auBucqiFuACc9CJYa4++Ypa46CK6i+S8Q
LBWtZAkm2VUqFBNELyVK5kYTfNQkFO37M40RJUpcg72aXZZpgpyeS1ikFEz1/cuz
LDEi09ecsU2vilMhKBXyQSGA3ySXHX9DWmX72mOUG12p+Ilte5xRTLJ92ldFisPF
8sT6ywFMOgmnpS4HVfMCDfn6x1EPf+jf27fvXi6Ma7vhyBTkZ738yi50NxY8i4YO
Dfhlui+jYSeEyNyRHREys/AKSfnborOWmzaZNkOGCVoI2KgceD6EiO96pIaf4Pn5
CbTrnWQCs1U4PDq2h6IYqUS9gljZK2VMZ+/RtFe6m2sIy6nGd0JTWtZ0i9CxzPlo
6ejkdEMBEqaN/CuNu7GS13UAng0yBkHixSlnE09RjAP2/8t3TQgK0PcjNw4/GdTq
vjAb9bTk7ajUdx0JnHxPMv7NO2zCZ8p++gN2WJG8d9pX/YQkEBX2QQfD6BBgdvYC
jUpljrdWnoJZ8EeS5nIXnDrv0YqHX64GmPIiQ0Psn3Mv368iu0S/9+rBlOsrDgrs
x4YeKbKUggFy5KsCu/9ZRY1G/bRoTOPs49G0jYLXGpaE0hu/fP+GBggK9gy5HVD9
uW46ZhyET0ScLSvqPrWXxaz3v/vTHUvbRpxlLGZ6jAYRZ0KdUNZt15Q9ad1eIJ8h
4DYWMP7uEapWHGRTlg5UlefoCuoeLThxC/JFh2GBUgzpLsAngc11VXPwutYX7nrI
sRgKZ7OwnG+Io+NKW55p5QmL3XRbpmH8D/ZZN2/nUewcd7hVLoeKLikOk88ePmbE
ZjirQNb04Kn07P7S8bRL6OhgbiUU8XZRQH+/MHXqVJ9KwXNR1sqS1tCjUVudX6Vg
HxZ0e8DQMSr50PaVL6cjfcTOFnh0vOafL2Jgv2xbzMJs1Z3j8A/gmYP+FSKqRgVm
N4+xgYykcVJMZbAYDRi5T5GH+WxZsWnzazbyXqUB130BL3f/ALpZk2Lw4S2xS3R6
0AxlVaxGsmQYmvz2VYqlr7R9j0FvhQaeuzC5mRsDCSYkPEa+uzWYk/RmD3IxVL1O
ap8VH99gjY53w+7/7IU2/cZ+nBSNYN//NRcbhaQFX2iOqusDeyk+GV8lx/K+uD+r
CW0rPjdgTyFqbn0nsx8Uya2ud9AucEhvPS8zdAg5xazl8lkv/qfU1CYMV16Efyo+
7lD9KIIyQku0nYKrEJul2+LQB9Sdo8i7hWs6sMBdkmvt0sGE3YSc5sx9vzDeoUeC
XnshQ/n5bX+Wqff9CBNSjj9FbA7+NH3pIH0GpoV/hjG5Tg8ePsoZ77T8amintTR4
TIoymeSZdOHIY5HyN3eZlGLFhdaU3dRC5n86OmtUZ9KAIPUkGoa2Ki1yP31O6zBn
L2SdmXWosuhhU/yx0vMG9GmgDsjIsW6otJm5+2Mx8S1YmK1Y4loiLBtdB0ZBNvzq
aPx14UwTokZCtAFLTEe5J+wk0EYORV38Chywm4zpzbThJOIVDaEEnM5asNbr2O24
WbBPcg2QVJqQOgBHACMqSJRwv+vGl7AW5N+/Ipy7aMWTZoNg99YQqTIqlAnqZqRa
8g5WBb4FBQ0umBEXdDt7WjEx4pAjAqBvdtWANm6uVO+ID+i5K7s1Bit9Hq7kX45d
rR1WJN5v5MJkmu+SUsth441sWMaYvDg/W+8tN3mCd149dSxwXuwPp7YAslWern4+
7fM8bvSmElcMQcp5uzwWtE/dXSLAytZNdMKkoRNYT/F006E1h8OpheA4x83K94ho
khJhe0G4t7wE2vY5N1uEWiEVJgXvQOsKUOBWxeFfhvnD/HxUsswYpFbqb19ATd/8
E6H5LqMEtsZenK9aqDmvZMKyoi9nzccdeP9r6r6meEH7ky5CuWaWaN7J9/nzwESa
AJ4BwcoEEcHRieQH8XO0l6s33RUnqCwx1vCTUrsqQEY94HGU4oZYgobKMGNEx9AL
IGCNP2nUMqA5LCMac5rJJP0/tw4/sgRYtIS2yUercNgUPNR1DY5tbhh69C1Z5ohq
ZZYYfwumTsbWVaWv1T27EVnYgOM6Eh1hngRKfmWZ5UIlQfpIxpWnaoKunfGeRJJx
F5bAAVrZVi+YsTUjbsWYDgdsXMS/4LhpAbZXOSWZmNX9uMa0+A6LAUtGex1ZvIBv
zh+xMYYF3FmZRJ7m6KmH8VF3bcApUmLsHdJoc3Z1QOjsOu8jb+V0gmOjO54ce1nZ
/jLNUzwxULcIpeHX1twKZE/EsHr0QzzncqsG/XqT/s9gWqh7OJwM7s5UkPULp6J0
4qZg17CUBggJtyx7ZZBV/Fc4cTYcyznU1I3x7Hi1y9Y8TiMHI8RbvZ3SneBlqY2v
RtXCi/QIPvVfViLvkpr9FazxKlTGobbsh8WXxYb1y9Xp59T8Lkm4WgrbtCocqFvQ
Y0tWj+XyuZN4gNhNUOEfqcdJR8kE4sn4lyXHEtyJHUYytpW/tEcN+GAbbPE02UaJ
qKpG5GEG7m3RBKEaqFV4tGgEUzXaaJsTvZ1h2RZHmP8FRBYp2AbT3eID1Lwbuwzk
rJ96tnv2lcuujAeGVoPeSU+z6veq74om146S0NpJANDgkigHtPXbdtOgMHCSrQZC
xiA0Rj1AMPG56oIDnQ2Pik8E56bBkqU0udXCSf8z5iPSh3pqRAVn9rTgK67ecdwy
+eXjOznT6wqzxZPkwR4MaV8ehEEVo1ruZjZaxzDmj707LfyqUn1ZgOjS8+eJeSWC
qkRzFkcEs2xdtClDEXCXIyhvX5caaSfXPnjYxXEJpmA9W+W71/qpq5PVhwt1PTfg
W2EsrTK8YlJIUjPTINaTUsIs213Th5a76LS4hGNuO95xhpbc1fBSu1Y/HrkawevI
oDKKV6vHu5X28SW2HMLizTyC7szJo/M3j7PhkbvDqNp5CbU4bjp+Wo3F89JIFRwn
h4VT6U8qwTMh30XXfi6GgNd/nUitZTMkFrGeeiKShTxwN0Kh0UsmLkm/sLVNQalQ
yVLfxew5zLo9FLE8Q9R+jHaRFRjmHZ8vg3MkjWD3pkLmvxJL7jbYdSERGh1KenlP
ztOEEfk94UpKW3wzwV6IuaRKOs55/9W1O6cfFGVu8P/ryCPMr8iUUNyZgNR0Nv1Z
RELUVvcaA5gXEA/N3qdde9PH01tY5jzxeA3ML1T4GT7XP53nkhP2gcf1JBhWYNFN
aQrkeXJjI8qYBerRqb4X2aiv/zDSkGZh7aupD0ULRat+bFTCzqgdFEQ8j+15eXbA
38DS5j2b4oP0V3P0L36q0ELIFQNSo8o7PuYqc3us1N102pd3YJiGWbfnt+uRy//c
dDH+EY6BrG2ibq1ypVeV03V8hP3/PEEtZ8GCqszAJhrY/lH3D8nWvgn+zCJId8YO
tU1Txh1gzdGNCcQAe42yPsZ/ss9vOdML7w4xroESjmMoeooNORUFVpkhDhZDVrP8
jiBWDc8AVtc47l6uqD3UrX2oCOPKvxXmaF2CxVP81ow9VfUGVrN6VGGaQpqm2OxX
wPRVYf61VzKCaRi4dzIiaTSeDvqsZ3q39OE28T7wa8lMTxEYeEr8qxkTwKm7wLz6
o9aRr5XcOXLcUDrNSei4Dh+DgkhM8lkLTzSWNuyhdnyOkZ9CBHalixVMRprFMynU
jelJAAMLtUmOUGMYQpEHQrQ/6z6ES7mHdB5/PJQPXLYAeuIJZZOAvSuI7+KlPkw7
vHL2XlQuzugAKJgHZKbQxuBNmdNxkrHuh+E97IGoitkh8Hzy+MaEqz3uwW4SS6zH
JPGPjjCQUCZMOCQRx4hnL2iT2n6ejyicQqCgCDcUacEYTTskJhtlyziJDanipidk
CTmdSdDwBWkoqVumsK0HbXG2hoS7IfUonzT1mrKgJ9H80S3ti+4mvmfPAvmzA0ok
vaQibrd1AFrcK89+CRYOUut7HH6dyg5PugZwF72xh7f9fthW4srkB7jrjDviJGbp
EsmIVZBYDoMF2hhXfLjimjUGlcZxVppo36709a1OOmD6OVGT0HLMcNaUoe1JRKWc
bZxtfuYMERZU+YpuVa+mfG/6hk46yQRQmKa7RnFE/4OLVHXMhmmizP9mD0xk5Vhs
PXoQL7KXcAyRpPaBC6hx+kPr4KqityEUDy+tcc+QF+gtM8iXj7KPBUa8wNammEbj
gEtNvnl3NYS2HS6lgZhb6TksYyOv2HQsRYMqkqSveF+MH0JApSlmPYAs/mUz4gpm
ny4ioHqO89NTLCICukAHlEfhLBBgPj5FgDyrpCxwnXgr7qzTReg8vxe94Mq9Qg/q
krFJ5kUB69t/FP2ImRS3dj1+fTnwnXr7N3Jv3VsiGcS2Xh0nLmPD92Wa28HlyvmK
D4AgzRoe0kAGsQ/TQw6NGF9bGoNau2lSiIsuryeP8uKUa4i5L2x3co3acu+Rv3fM
ffQUIUf1HB7tOxPF4Cr0Q0q4sscew/aLdcrX7fdcahu1ziGPDPhmgMtvpKdH3oLA
H9wRGlEefURPUiemYH8nkWKLIDmT7RQA1JE4v9cX5FA9oLYnnyOJ1rOnF9qRnG2q
eRf6J4swHxxlXk2hDwVhwNHg2v3gu0zz9wDJFQ1JF7p6z2eKzmpvzscEyjsYbH8+
nSAZsZNzMgIzKbRS5cccEvHur17dcTew0ocF7mQNH1DL+/PYGc/uNeca7zus+Kvp
3gUbdjQTUGVkVEHYcCUOSVDL9DON3hLTAzBKH2o+F7jfCbjdsXHuBPB0sGP3W+Ab
sRmCSUunl7DKXygsFXgASkiCaV67SrLjDgv/c1fBaaAPv2KJAdkETiKgltpHBAW9
rHXkQ+9Li0soVliYgcrwgiBJQpuwQH3Wh+18dOy3WldsHpxbMxsuwUoibIXsLEyn
WdfU1TpIlOl2UoCEecHLFr5tRgcOl0/ETgtVOiReBWvYf9ohVrNhAfEhXgYSa7NI
nfqEBeSNVewv+cQO0+b6WH1nzUGOpMB1XYvAxEIDWgqqHdftOPA7fgvdCZNFvvgE
r0DtYYgS+WRywU9YvLYoyOJXwuo2tAISOGdUdXyCHY/tbyPbsQfTKm1FTnTyJFMr
ybGieIwKo6OHYLgCfzL9sp5r6zWGyVE9wz3r6xUAYdnUIDGX/sMF1B/TS/Th2K4Y
1SgQtQjJJtX8Z3kjA0/4Tl0JaASs1RNDiwvqSOEpc4VHKiaF66BhILzkWaE2s4tl
6Rhe1oRO9sbR+b8Z2vk5GTimas/peNLzo6YXy/Rw4cEdHarei8wlYu1k51oSg0CM
DmNJ+gg9olf99gCgS8zPBLb68IX7K8154zSqqCM9XeI3yx/M8kSM+WjLaRUDPSpz
YNmg8TdPg2NRwu6l2rzTQEO23P70mzoWxDr5DVDN25FQfEH7gJD4TaOT7Auzpves
umsiZnY6RLIJwTvTLE7V8Z/c8+SyoWkKk5u0lhhW8J/tdsZwlLKvdQc9b1L6//H3
04sW2VFjF5N+GgdGNKhQZynqFhIPzUVVXqHBaZHYv5OmQ4eucopJsCdbPZvJhw5f
/twZH5JKFWk+jxwdKvEkucNAL0DBuWhVNm6hBFeU4kVIj+Ib3dGx5QxBHx5iWW5U
p/Qlvru1GBjDneH0vQhb9edwXSWoFHdppuweBxVer3pxwG+EbNKchUeSK5TMHxL6
Xgch7wImz4bCqn4N+gLI7t0xNgY9u8Tp6qAL2ZkLe1a3j62VJAAZRKP9sSa3knjN
RoEVS9Eis0ZleyDiOWSzWF2hqTKwUe6v5tgEvWGwBLMyzCp2GYItBRnpZzzC6rxs
7GoeMn4l6b983pNuCNylYlXIt1kyqhXmJRjqJDBpJ8KlbhxlBfjYFyMmmAK1Fmhl
/e1AOI7FNzfLJGn5U70TswXlKimrXJq1hckHRXRgqxWpaU7hO+DpakiOA0uD03F5
MRiJn2GtW6WAHu0HW+3OApaq8/em3w72DCIDU89JZjz1vuWSHpOu0ubWFcUnDw+o
lWCnGwn5+MC9EVwJkeCULST6MSeXqswMqHokEV/RkD3xjKpH3z1rGax69SpgcJvU
0ORYljfN7S0J0CiYRqUDgC7iWqKBFdBy0HrEzVBWc4vIIPJROZiProvJ2SkRU2uH
8JJ4JWQGdZ0xyWKpATusR1mWnsrOt+AMEju6Hne4sbaFVRRPxfnyUl5H0scmBgkY
d7qVoxs7QcqhIZSHG5vEcvMKu7WcXqXmErtOyOSDyeUtxY3cz9shPpp9fv0KtpTh
bwqt6ef18qz9aqxDt/SJxq8yraXtL5NKM9/fyeMmtHnZ4wKYIs0V1hWkOGk9fjoR
aHf/LaFldf9ki6q4X0AoRHsOqVay62y+TtktDu/0Ndyp5Pt8X8kjz0SC+JrtFp5a
sxWRILkNG2bBUyTStqZkbEfYR+LIyKN5w0Tdtva+sjaPwGYSpQ3n38VF9OHzxQO+
y/BVm2wjV1LKtdAhLwSYycqdNFd6Fs4SYdYdg2KfTAPhcwlQUmjelPIVvq8z9brz
JEiYGXiMmOUw4jCMKfO486eZkPvhcPEAHvHDkTYzOebXUSBNjBXugdZClRFHrhv4
arFMCCXYOytmeV8b5Ej0LFkRfSavq/WqdmPPmKxYF+8zu03s2kAtioYinMfqjekO
VmTkYptzHEoLtsu+M4qqfmip/mvZEEPHTGmxaQc3/ScmUnzis1r8W3+l29fs6Gsy
a9FrLmE7t0uCyss1BUYB1TgSSsidKgjDXzzMXsWUXysPvcmdFP4aBghWuKl3by36
nQ0B6wlGEpxml35tr+FSja4wl75lTCakXjZeBKfldAWpcGDDTGSok5V3u2x0Hg1u
o+tScxZvZ7JFWCgC2UfptRJSLWzqgNPBLBPhThoKStKMp89MWh6hiKv50Ip+3E8W
L15aaY/liyLK9wndWurScsWyJ93St+eJX1vo9rRvUzRzQtPrc6qcVHEtKsBsXyyh
MSz/2fi6p87BwbbTs7SnxjcSpTxEiP7b9eWMj8m2pgpqoU3pYicm5r59SCIySylJ
0HJkY9QWMU/tVI85qAmbI4M69XTL/AsrtfkCtDXxEWsL8phc4+R0lP8fMn0O7Es+
0z0Ze8naNQehMvUw9hWqD5sBCipuocMAEwi/4fvfYWkpLgCqJ1ReGIJvaEk7ueoU
JXo991v7f/r9KlqVgjmHEcNe6B6NOpQ5Xmyp+zDLk0Rb1PNj1JoJqjEyZXpbcS7+
es+ZO+qKrd19wDHwiWCOUihwwB7c06x7lliqySKh5ImN5H2PpW6oI5wWKzE6vYhz
w8Jn1X0RmUakfYnIvgYD346N9tcmzRIOwZzoI3NTLLluw3xQ3qIKS+M4zVUEmDVO
SMk6Kx8vw5vFX/aGtOAfCBt+vcgTpI9D90z7Cbf3FxCzFWVEYbCaInFCCcjrtzhj
urAyjJOgeikOFFxjQALzwfTg0c5c+gOJHB3fw+CjRsFEwkN4E2esvjUxS0slGeRS
KHjZM87xfnyprkWBV1dGo1O935CWGEaldQgZmU1ZIV1PRwb3nUlhXarGAzleEj5O
nZJ4OLoM+dgtWK2zJo7+zSLDEJxAweuDgTgzMeYVxenjmsOVQcwbHwORtYEg2S3+
CniNH+mGGNZdr7KlMHKCVTHz54Mno/EtrHySq4cOyCiLYrJQ6nHwmJg1UFBhzt9p
PanGQY9cVQ597MuTu4PDPZWHDYVZt0k9wtXxf7bwgc7xzQdHfQr7Y0pUpPnZRcrs
Ne3ukFwCKmGfa3ZHm7Qmf8eWA+dMxHWtDfaFzBm6mfGQaxa7MP13pBCDwK+tGViS
NLl1IIFWWxW+APjy3N5n0UCHNYO5t5aFV0Zz6mk4W8Ra67EAR1gcmmsT1iPaW7R5
0yic0OixPgmsVQQ+HyxQCYGXfDoazHJeiWfzrFi5eKVteZ0EBESX/cKVvmsuhvIz
pTTvX22g3Ey/a/eTqTUIkj6vTJmN9qjtVrQumAkwX87GnmjeUJWc5ANDAUkcdCh9
20zvbKCY6hXB3hgwLuUiXynLnLhrxpQNFFzv84fVmrbg3uTizxUIrW8rddY/WQKc
qa5VFydq7hDd1jgX6j15Kakb8q0oZkhUrEp+6g/MrIguJ1XgIjDbfIsEyOLlhmrh
OSO/LhBftM79ZU5quwGerK0qF7ofYCilgLZ1hkY7YewnqV8Yd1oXIzZ09uh77/1T
0kC3NcokKzoCt6CgDEGdXKKxDaTRee+H0o6AZhZ+mtvW1EGh7lOxl+g5P0sfJzSU
6sZ2yuDTgD9/XGTZ9kv/yftbGYB6fLHp8voRMDx0+Nyt1oU9WT8WGnFV4PJgGQF8
M+ds5h0Rzr7dvCNrky7ALqzM7vCTkYxyUXcsl91u7RLk8J5662MkfCQ2+rm3J9n0
dpf8PgAMYgieGd51uH8BBL7v+ivAhY9RSJYGa9FqJa1uy51TqF2mzabXpAEjcxEm
sG6rfdhB4B461YSRw40LzYa7worpkJEMa1wwbWrCGuz62y0sqQdHz9peM6K7yA/A
LMj/Qg0REpWWv3ZfmzbjaKpizvzyvJYVFWAIoNU1idamvFLy3cqpRPadbXlH7STR
6nhVUABcdVNBbkWfaK/B3rcnO1JOWLGM5jgHkEOEDbIZPhsgaTMAgBgfqCltHn5T
cUYYhNcqQKeLx1FCwfGogGC0ufscbUBzA9eB57ul9PefVonQqWiU/xPUeQJ+K9W8
SVmWVL2BRyJXOTqDl1eK+YpOHDQfL/66sXT36p3N+mCPxzQj5PhJwJMDZRdtqDF5
tf0pLlrMRwkX0yOAts5ndNMdxoj+NOmWecZPZvHBkRNMtE9hv6JGhVVKRH+ZjHCV
BaPa6/kVme4BDf7FkqjX4BLQNh3PZQAZLfFCubgdrfeQZ4KzUdAG/QlXjpNT7dxs
WZ2SGFv3pYQCAVjjYEWf+fqurpD2jLVZYetr7d43rHwWwvKiThzr5v1GBDIHQpfA
FzCwvwYz0TvSshBla4rhR02thPLE/t2MzmvCOkV6JMy6LqSH1okindOQurWIOMN7
GFBvHQQZW5phiFPeadSD3iFkv1hnFX7YFY9NXRrxDaUVEHHlfpzhFBAMIaSFBT3j
VuTQ06Zzy+LNa5bBrO77zzX5EtLvYFeHyZLkgrddXSPBsfQPuqEktzQZiKGwVi6y
vLhPM3Hw65XDjVVfqkGvgg6TDLy19ZmSMIQO9RdgmsNmGAfW7cWPNXQC83EaDMx+
k63BIPUrRte+9vZCHRGhYj39NLV62AwFZH9Pmr7Ce7rWUZEzRfirquexRFrswoyq
PaiUq71PK66q0RHsYIfx9Crkl0xJeUExLTq2IBewdsLD2l5Pq3JlgU20xSEc5WHN
h8ena4AB/0QmD8oxoRjd3pCfqya2ANSS4YRZ4/VohU/pmd34//jUGdEh7VyabR0W
6f5gHEHictAoDg9ms9gjwlxebDFnWZhhHsIM8aEvA+UrHORsKS1c1Tp5YV6WBanB
io9k0ZKpE+jBo6dV8ciGho9Es1m5fxTi5ASfmZLkYrtwoJ4me/yBgkHDszuDch1A
nQIEWU/wVgpyNZ8kwMRm6YsSPVv0iHsK5Aj3hY6MiKHIzjNyHb8X3vwiOjm4XaHY
X/iOAncWsWPG0CcX8bRclps25ifSEvy9hckmvif41VpEaOuiWw//y5VdTe6U4oFJ
3hbHBVLYYzxYi4I6iNWV+STkx1OuRm8hpIiFp/W9yR+JsiCzQkAreQ8jXQj2DdaX
XDqKEf9E5guoLBBy7xevhmvawZ6orda51+ZlQkBfiTlCWzAixUVkIFsh0qRMlkR+
WzhZ/GbRvY8bANBjHK0Pht5WMpFAlOxJKpc+P7NIGBKcvzkjJ8Usn/0dWbLhx+MV
5VPhHUfnkFjmWXeqS98tCi91zKY+DWzofNqMea5rnHCVAsnFsLHKLG8wSzOMiYPY
X13uWsRLGo6QvXseuXLWS9kvHhv931Wce3MJdm1Xa3WeM1HysCZDBmqD0pCcn33h
Fym42/4n3LRJLUVnZ6dqwBme+CXPiULVZjf9MANHss25Im0kBljQsfYGnr669aqP
PAkdha1dc+qpUAdPEadCyb5IgQgVkLZnm5p/lumePIJ/8RIOshN/QzrMyg4UCKYL
tbkTnRYe7pmfMESEnIDbRZg1kEqlCoGqOWSUepyG1N5RC1ssUhmJ1GZgAf/7GbGC
PjnuR/yZARdmTRu1AOuMa/JgjUOBVAtpNBjg0hJ1hQGhaDeSVjmFuYP7Q84vkNOl
xGaqR/hRHBBsikRsdVbiiDMTU0KP0WMw4tmNAEZH8AAYaIkMQ71Xwi69QdV2LlEf
uXdsd8AGc+2YFvSclX2nXd7P+6E+oSvz+hLLK1b0pgGzbdBj8xYRdFWuWu1iSDzv
uhAgIpscgZI/lBCbbS9w3D2+enlSazvXAqypQLfVBIfFF1EHe1+eqz3a3j4SWN3Y
z8ugPGDdi7eR/bIqVYfOHK0tf9io8kQvQFiXIS+x1sRCV5Sh4qcoxSVLOUaeD070
qj+xGxGebZsUOBGNPAugujc62CeKYtwODaBUc6/+2WQdSa3fmYeYO3MxPMEVEjx3
73xY2YpUaNOTeP82OSySWboSYFWasYuiN1J/nyBfOcCXyeLKg4q1Uzm1CaCdpQvd
SFdcS4E1rxc7A0giOEV2Toof34O9TO8Vul1LvjdRvzbE1Iq0fBUulloO/ztFbHMC
R1+O+qUfoCk2gz4pB6Oz1UADQYD7fGT8CX6l69kliKqkqn2i/HizcHm6ZJl0B4h2
d0Qi7Wicvz0WwrPWgQqtM7njaC/gxD6YyWC+ZGHWo3TLJJlq1JhaN/WSu90zNZGw
Dgl3IMmmOVE02O8VOvtPqJK78flMYJJ4hD8oT30L3vjuTcLF7yVKMjgMOHq977Ds
gkiAgC+WHxvko+qMmQzlnrNhRUTRa4t42kImZCLWQPslUH1mQ6EQ5RrtguHCJ58s
en9BfWQXQAXs7X4lZ65dwtVkBTnvxWLnXYCaNbyd/Gt3SOlxPBcC6evntudg28Vv
W1U8RH2dawxzC5HCtSwCj/F9rt9zXv1sceMWAdO5e7apkmvJ9ViFLkmyoEwd+92U
T64zsCUed9i2TNFACwn0Aei1NID8L19Nqg9/Yt4SfMjgoj2Q63i9D8EvQUyV4qyv
UHGwMRyuUakyrqBnvtNRsTIzzfegbbbZk+ijiDszcaCI3DM/ngKc1PE5tdXJuZ6J
J9vsRA9VSGan+UsScHCDPewKPIM+D651bfJqb6ml9WxHRMTBfuBKBavhgTWX+tNg
N8W+L5AZhAF8iBiiUXpYVtn8fLEyAnpIs8jMaTtnKHqmNHC/DKXhf2rnt/zYxxxv
UigW/GB3H0j80erLT4uVvSNYo8wbAFsG3Auf1eEeDtGH3Z9oKoFwB65TtPKFjWp5
Ysh4LdkJvIoDFmyc7PojkuvCWQjnavPGw5JWhDo+c/qN3TZUHuZcDTb0Yp/wJxTT
ERUgNmizCO9NsuLprQFaN6E95pG5esomZXMXLv11VBrzM30GISrtkF5WsPRwZwPu
JQkbVjHCC/sdTGLM3leer42di1HvqCdyzpFP4zsOp2EKUAVzooUXQkOPoC/kxRAy
JqPVxTjyW4+52iVQE2TmQzptS12aUu8iGndFU8rry7vWXL6OBq5wJZK+0xTW2oeM
ObqRvUG27f7t8v0b7pW2SFBsZwltLOFutlZNRlC9WONJGcbB51FVFtH1ynwJ7Mwe
AY7wwgx4XOQuaScUSX7gLjAcYoQCSt2tHRI4TujvwGk8XO/4KGQiREtey1MlMiWq
OYzwO1+h1IqDFOzA+fASUy831aSXGVpl5OB+V7RvojmPl4liV5kS8dzabOIA53S0
vkZDxuWZjl0PsCc+8lDckc6P/KVqNI7oaQqxWRTUFh2bgyqae/17eBzDfdBLEUNW
oVy5XXlHgqoq6a8NMCTlwY9DCsnlWch4w+FOns21T/pgKmwlA8YXig5J7l5Q+4w/
//aMBjT0et/WyIm4cfui2KJlT4azQYKihiPnfHHBgq9a5PZDcTSyyfFWVYcoct+g
t0ERIR/pxt+KoNvw6IM1MX3/WbsiDOHX6sT8JM4rU775HLNWXTN5iKDXv14VUGqA
PqxWBZsgLrAGK55e2LcTvqwxqYT5oRe07ZOisA7WIxIjQ6gaqTiq0+Z00Ac0YKeM
oHdS1VoArNnvXeMUHyMU9wKXPt8gLq5dEB8kyiP9Ld/u7we+2mXyPubfM9opgJ/i
BnMthh2EUTubSBcne0WOhQjF/zcP1mcVzw+9Hfogf0PEvuqSe9TfFPyHCmFaaxTU
5E4oAJpSIVjwFHqWksZmzkEadgitudOL3zBOC+I7qCVKAaNMWtNK6zA4+IzuhvAb
5VILWtcBczAjq0HsMi4xSKJ8Tab66GA81ke9TOgQoRefbFr8XKp7xw3UxSOyedVY
nh4AwZnxj4NX/MdgZ28aLrEOqW3Ya53emNFNoXWBMRxYhZnHPEBiCQ9LlXULyL01
GEFdPlhxpAUNoMzR5Kh2dP5YCrWYTm6ljhopgUQs4RZ1NjlEccieCJ+prrvRnR/1
0zHbJ5K20MiU7vK/BEcwnP/hwmKG2clqWpFPOP0BWSqwE5GOqp2+XT2pQteCz70+
IUmUIGaxzP+X4YefNhvzbIN5/ijvtldD4dhuanf8lte8kIii0WoDcCssaUCN9Tnl
AaeOBspao5DfcTXWR94wT32xgGfGoazkQjwbG3yBDzeBWytLRYkiacKvk59pV80g
jA5FL7EJzg2WD4pMHppuriyYcSF4uogDnQ7Tz7UDjOf+N1OzlSmZuE177CA0UpU1
MeOxIf9BPa0r+gPIV+XWOaRPggW/70FO9n18+FNLTP4JYBQXhsV7c4AMXffu25fM
93NcSXiQXnKRkuzkDs6c0XWtSNFFJQ6DL/4rcUxkB8IQnS+kh6V51UItbmu/sc9g
oPE4oLC+lApGRoRmOh9ICPanNOwbysNtU9IU55f3ETc1PBsOSqAc76pxgz7qrzR2
5JMafyloanCNAcB/mq5I5sx9vu2hYXEErC9Kh06illMJI1Kt1ni/6GQD9nJ/iav6
GLe+Dp52e0lPI63SmbigDHZmXL6x41APAbQONFQeuBehyMEjyGlt4xX308wXvO3X
dY+jfQ1Th0PdYhWYngFMAdabsGOm81+GLoqK9laJz8rVlXfDw1+LxcN/szHtpmRe
NfbPYX1vgkqZMjSjSz7LefL/ZsbOjH+LtOTkbC3zrVfJ5oGsI9kPkX2JpPQJ3ahY
FNVOOFW/8GGksa6FHNZVpLLuRkh0J3W2xxNg6XkMIATVBic1puKYO2IWCDOMqZo1
3sLjmjOhqF95kNqJXp/7UHWnWbh4w8VqzqJJ9zTVccpv1b41A7tA8Sytk1gbqdw9
x2Yfu4N5HPh91XE+uAVeCIJ09BzDqdv2TvqnXH8m+xmEjhyQce8+o8eur3GwP3dv
qZSmtCSw+7TlfYMNml1D3WWzCHfUK14qp21kUdc83SAS+i2E3ORnQqiLUqggjO4K
CALOixHypnkmW23vPfb8FSzCwyG4RXQfMdB3CpjUGqXLD+cCO1u0eSqI9irVdddI
Q4UBSyVqLPX1aeVG5shpxYPt9pkUH+G3+gzuEH+QlrDDPL8UTtQs6UJVJsJBwoON
24muv4rvk59i8Rmh1DLtlECQFXxE4X9hnImLshzuuRtLyWX3zQb1EGk25oPZSdHx
pNZx4s4YIUVx5Fb66ZKpfVtmrYrKHHFmQn4tIetNnZbB8CCofSlbqf+GbuguH86q
aQezAYOf/suLH59x5U0btcxF3XzFUs+svolTZkpxDflQR4QvcyOKrPZ8Erw3IhQf
ctF0q0O5g4DMsNSXVjk8xeiFx1eFAE3PWJNueFxQyU0/kHLczHj/DYmz7Bf9FL4S
ZDJ7FGUVE3+tSKMGYZMQ0maNWx877/p3dguxspUSNIkNJ8ekXYoADGUIESXxCzJw
YLvCNLnuwy/7eOVT4906Dv5y6IhELxvHCKxu7OZYFCRTOKrvSe3AAWpjl8OHfawR
dzTqI6L2P4kbrNLILB8AoxoWMar3nMYLVUKF21xLZMWHk+Zx9+8KCtb2PM6AOif5
mtyGEgGrv195+LxkXNorRwc31i05fp0/6/BEI6dqQVVsz7s/XnJfiL0aJKAcYhK9
VkblKcX7yWRw/wKydnhxCd/5VCUTiOUhyDOimdA5G4W8gWsKV/JAkv7GLqWUftDY
QCVuZcn8hsAPz8fGFl1gapRVtX98/YqclYuq52hkPmAQXk42Jr8jps0SFc1tBvX/
R9IpruvTI0RE4r0KPoevwlPCo8Q619hQWk6t1nU4FNHpDmGaHtA/wtkvCCAuVs0C
UY+WEgUFQcsGwdnuBSs5mQ/39RWT3rYB/zpKqWMrwrzeYMmVARb2QORXUwc1Ykei
vDdjrNoR4TaU3J4K16EP7qKUzvG7bGPJcoMmvrZaugDxDgUd4SL2skq/VVPiZHrY
I4FeWJrylmY7LnNKYs+NU3oi8wc8Ghg6fNTDS7+4I/rZrowaeSevw0Bq3PsZcYXo
GcOuw7okszwaIFYYZ4Hzt6kBuh78oqEGE1cfhTAP4/9TdFH3mpecjc2AIABFlrQJ
F0ndhgk6LBWn/VzSG5cCehv526yh+2gd4bnZQcXrISsyiA9850OrG+NF4RKeVyPW
7T6K/yPCDRl/8Jb+076XMk648H+YrVdmTqd2kFQTGVOxvXG3L8dRXmVtpEIKBY1i
eibg8GVGLJ8793olwn9yvOIUFx85uW9xM5oDoq77xAkM+UT5ZVkF82KtEGAJBlCS
lNLxni3zCjdkfU5ROLuaHJXT7NiguxYQz+hPfh8e9w2H+XHHvn31M3fD54FMDmEi
4ZiVmrO9rXqlDF0PQvfx2e1dplI+KmaZ9ElEZZaC0emzLt+N3RSbO+eDHA4Ddw7K
9I4Bh7y0gJYRtYdwYZvKNtK/mgMwdGlRwjrmTvKuh3fzNT5eccQS8HQeidD7Wr2s
BSKn/zuBa8APGCvw1JwuUDjCPRmVmnJ30yO9RKefSUSnVNPr+6ob92t1WK3W06dh
joeSynNwQ2Gw5c1cuHb5TDnoGfx/CtTrFzm8xBPllKzi+DzvAfInnbQBSdrQNReP
4ZnRTRV5q7LyNzd2zFX9nC1px46cu2WCMYzjLliPRAda24kMm+VokrpFSpRlxuOb
05/hWIt79Yw6kC8lYdG42ornlO7a1qQ9KzDe18LmLXxbywlVaPUuSe8eWT4FkOlD
inholV0nIEDKfmZj4aVuFyCttouWgrrrhCga7JLNVldS3lm+FrgpBdFPvX+LDA8j
f1fvzSp2ESobVlxCoKfpCUbYRsuvnVJBSNVps9+SPABZU6Ea/j9ZOgxfwPlzmaL0
rcQhhwi4WuQY54iZaAVkYRT4AsYMgyOFeiPfxLAd0cAIlytJbzbg0s+ob+Zkn6Sz
eiNfYVMMc0+7WZ53H/HPiE5t4PVHu4/P5tlfaXfBXcq3BhbHY9iJZOvK3+CG5w5S
5+1/L9kMcA2NpCNRjYj1Wxep6qfDbVxZhW/AjQtTYldK4ObNNsg6DTcH02Mo1vgZ
6m16WwbLWCF15KMNXAhglTYAl4TqUVwXaTRNetqCH+hoqpH8EJHvPwSlOxQSGvbd
18EGUFJ4cYCWU9KhDAnNHqolq1LB3PMov4Q4Z9/Ueg4eZDl0wo0WsGKFoOeeF7XE
eoEZaEC32VMtkRHMpM9PYjFKcTp244787hplpNQlw/QHSSdWJClnyLsQEPF/YDHO
BKNx33qTzD1iQCuWT8Dv/L6K21EoohorSyf0DiKdDacQl5tle7ROVxZ5L17CWCkK
9yG2jfy6QN1A8T8QeQbw3ZMsDkejIXLEywo5/inGpDlPK/CF9FsLOo7ySp6Fw9RO
V/ytqeFcaAfr4zbCkcXLaZDfEafFs6DC+oGqRHgi0jhxdyfDPsky4HoBCmORnbRX
kj476iFD0NHJxZavyakFMlX28t92NvBzd1ttaX5mrfCHqGrbg8ZZg7fJ0LuNyUTM
1N51JQq/oLxmNkEm8xqlC49qfIseOPX5XRCJzgYo+/4eorjRVej7KWHOZjw45v9Y
eCnnLxtraVCEM6eV85zvskpzVWmCN3p0Mq4NLPVtn8Vim6+9BXLLfdn5dogjN+hH
jazoUon6jZmw3IZ7cMVPTAfkVBlcbY692FK6BQdURinuPPuEa/407oXfOtjBQlln
yqNypgFx6UocPzxv4+V5VghCkN3r7dEg7AtKkLrt5TuNMvz6nlXaSuMhHJt/duhI
mNiT7ap+LMmM/KWcTgo+DK17b0Qn5x0SlgoJwgQaSCymcrBPkqD1BFX8BL2Ylofg
Gr83I9WgaANx+CqJklzGGnumaD8PfLQnMQC1jvE6cbmLRAk4vsv9rf5O4UqQYf8q
PvYExKCcX2AcZTLl6QJsjOms8tmXD+vAiW6qn2MzqvBh+s9yai5ynMm9/uehb4pa
qe+6FZqiEkK3HhiKHBEqplYThD/QcS0YQ9mG0OJjSplMlxC9Px8pNdDxu7jLWSLA
22cycHftrZQ9oo+JHEJ9xKwirPTbOhwNrAoipgQL5fd5aCVFSqeE3ZeBYUaAmSg6
NVP6uT9JSenzI0jjnYW+ZeJNiRyRIzoIl4F4QbWWW5678ZewFemYCak9xczGXHmL
w2v4zMMb6+ti1yu9uW3HBSc9Z5JsEm9ZLE/xoVWANjy5x2awQwd3/DdBDMmXpUkj
gyZaA2jNvgz3vOsHuc/mBKdoNJxMKb8n1Sl/K9rf5/bcjIXiLvE8zOkei1Uq0K/r
jJgboCZpMg9hU7kxeRK3+wEPEHv8e94XxRV+lxmV3ia4kZhsRK0ZPokJYi+DgdBi
bbFIRYoJLu+or+1fVV3ovcFwlHJvKBFLV06heSovS9z/sGNrELq1hGUwEqKn/MaB
ijvNPJOtCUUZaVmEaQANDw2AAujYzsIuW9xdzk5SIoM4q5AvocGe+MjPVp59ZhWA
xIWrk8uGVAaQB06VhMqIzZ+ciocZXLHr4tOKW9gwZ9zRdhPjWupnmlYa0SKxoRgj
kUn0UJhb7P5z/8rhoZ1uVVJBdVPdZEr8/jLXnVnqzIQ/noCi3HpgftykcTqHh6J7
0Lijzd61eH/W1YTeQ1afG+u2MlDGybGVIIwsMkg9oOmQMgYof1HBTmoVNzrnE++V
YOHHedq9zM0o0AcQDPHow+ySZ+AklPNV4NECwOqHJpFdrb1QHuKrR3yYDMcEmVcj
5gBmVkfIMEhbomM6jxEMe0t5MhJ0Ntv3bjna7fpfjqzAt69AQXK2RMhNdpqlgn2c
8xPMJJHjRwbZLtgFN2oxAtjgQuKSSf/r1+H1lS4Pm2pKL5uVmaQX2FB0TtT6wO3M
xSCMc8X4OkWYWQ42lQUks4OvFunwIppuisT2SW7wGx41BZNFR8/h+Or7zteP8tLs
4zKLke4E49pF8XvDeCZvMsPMeB7O+9iAeiw2crMmckDdI1oZtQVEdZUwo1/9futW
osrbBcftypqSrvSpUB5ByWTBI/mmSdATqC62fk+nTRgoEKaN0XoswW8TMA1/Y+p/
w0Ff9SthTeX4EeC49mdnqtmfqDDRAJG58rotIhNA34tbLMtKaZRxhQeRC3IS5GUm
wIEUFo4V5msl33PA4SU71H+QXS4Q3eqST5DlGwQmIRHqrnLZp5rSlKZ3Ke4GKdGL
28pD37NWlV25EYEKJ6GsJxgL2fBhK6xMWPoOvIIEKCLCAvHBhcZM5Mb9sJZNfxSV
4W6hSAjGXa/mBV3dU1GcWLEpHndgNXnpAX/Q2AjCBmUQUXqUz/mUG02/kGmzE9xm
ojM8TWrjC71PWULuHu7rt8DP7kvFf0I2Jz8Fb5zKyp+hAAe0jM8uVFBv03aEEpYh
7TqgLz1i+q8P7h9ie9uCsPSvXEWLL7KRrlij5m6ROP+5ydN3OpdHnkYlngg0Z6Cy
Acgo3ulpsKAqkcN6VRU0jvXd/cvneIqmKza48JIdct5Zp92hkhqF1Zfc8q4dt0ZA
YTcISQyybZiigK8m4GoCVQlcdaz0SLgLfuK23e9V2mZCZmaUVcqh2BdX+ilmW0C3
kN8HK+inwvMLewf1EyBahw7IPezLwH4eOhcFxsQ197s/9l9Xe77rY+CiHC5wU7Nt
k1724XRYyb+GQp3qkitIBiwjjwprGo09Tae0HyLm34gxdULAPXsCmfix42LsGxaX
jZiOSrA0cU/24sxdi7H4OBpH29l1u0TGwWKyXIKr8nh0/eJj9eGDNnR1WN761rDS
Rm057Hix/AoOZDIP85XqRKZBRtF/Tf6VAWutfdFhmUClDWNu46Sgg3mUBH9An6qT
ucBotRT6seF+fSNRbku4Xd4xTqwAHzm0SJ9MuSGrdvu1DhYi7v9iVmbjtySUv+bi
GkU3j8IxdgtbMnshpvqZgQNbcAGAyNFWedzdBnoNISDEj51fHODx47izNalsteYB
4J/ilvdgemzQvAAO00GTZ165grqP9ZD+gjPy058mL+i4amDWCqvMZJNJRszPj9oX
6vSiXf0Fr1psU9MOfzNbliEFxVxqkgLNYHwi/wGssnFY9TVTqp5AI0o3c4U/jR5R
vUxvjpdhUbAXUSMkjWJ2Lz9utUi2OYOlSfCwbWtSF8ryHI12x+UZX/OZ3uW5b55U
N0Kt7C/X9iG9PGFHsjlBUWh7Qxcmy5IhcvqzbT1jVE7AiDAtUWfVkyeZuSX4UKGh
507/I2svrutt6eAK3BV45mkgScbUPKQlSnz8yneVG2JRPkcQld2qw86j+fmIqmoC
oHgu4FBOudn/pC0GIInhZc4yNZtUOGhpLPw0ZwGEdTfrY2HwtZPsR2qNWSZKGtkh
iHY48sHnlBNJMZNP7D5eLlh861IW+rw5CdiRUPSjavKy8UGU3HUzCZ7+ovjNdL6P
IaFtvmosg2hIxsSVk624FX024sbf/+RHwLkXxBamExK4pkn7GW5oF1OcAGEsVouV
la8DaYO/VydI1wLFQS24nA8CiOPx8QVTB5naPcQwWdhfn5TeBNwOFCR16zxVYvEd
XQbeaPvLAYs42Z9vxbVp5P5Zc3Okygvpk4+SV+sqPgzdmGqAl0IyHU2GYGHhPoxT
/RE9t+D1EsuIWSFgJazAfgoruSVbL3oIWM1PDMipBg16RIn/pT354PVsPzLyFDst
aElTvYAzwbTXesTSSL8wbPFFUvV25pIUEh17WhSbj2e+6+D61CLh0ej9zj03iyiV
QApEL/dq/tlH072hoFicdY7UG+dRbTkTrwKOK8xkxzk1AyJ7Dja5XIYxvtXCeCND
GArnbI58aqO6ZiYtiROduyGcrE/JyG25GIE05niZh/swH2bCfQ5mlrFYNTCFYOTw
hQr5EHVMOvXHkwihYymgBACPxaEjy4RPBk64xbRcfJmu+6p1PhvrbzsoieRpnp5O
kFiBY0wQPuBXvUJiG5GubNO/MdDsUUGOW0ZNO5byE0EHkhFFmCEUnCUmkvhghjNN
b2GYxmtjL8NRk4RUqldfgBIwzJvcIDNah8FZkWwT4acIYH5qVZ/0toC/EjoIoVRx
Rjz+RYizoWEtG54KY63ey/1r4YULtTwfLL32aDdGu9h2KtEtHmGaRsFvRaO2KDy7
ViKw2Hn4pN5m2rE2Qbuy8ZQoE0c/omsTXHK7xgEgO16UpFdXT5N9SN0eepDWIQei
mSINSiPwVq4pm3Kh+QA+7nwEcnHD6kIuHPHsFnKhloPHNkvJxZltGpf1YsKmLdvk
gy+UGcibtgAgxcx/q0oX0nsnBAlXsYUeUgI6C+Bkj+HbfJhnBTI3wQB0g3TyxUQg
kkBvhR2g47ckB6RF+rILYxWRiUMlbQFUem+Ej3+IP6gm/n+QR5brVZwIJ9Y0S7FZ
AJgKajMhKHTKW8PqUVjxTL8Byyez2Ie/osc79BoCHXZNytoZXwkCPugwgtBMhHRw
obf0KCEVYqlICusS5zPP8RL7i1aO0GgQqS7HtpNQxBtlqIlc9mVWMFa5wuUVMo1Z
e69kOX01u890JAdP1cjGMT/2EXGnzS2JMy03dM9ZxjztT9wgA72N4jp8SvljEGtC
lC/BsuVf2Fsi7eTIzbmxsh+a9ovqxTsIhgkwzwEEJpECvK4EEXUnkQU2Oi8Nb1c1
eTagDJFbIvGns1qQAMRpfk7OBExiXQf41EsZ4qris2AChmrxzVxbvs5NQLwBG1Xs
7WSLbg2LsSUBXjpmaLgQKW8xkHX4Ffq4yQ/t4kh+3ZPCYtenEBFo34VK95mOOjyl
sFRuObMo5qXYudwEjotmW7GkHPsKhEXPvCfQIfS4+Zs+mB3sUsGFzUysYzeWE37E
Uddw5Wezaw1Et9dBwXOwYjGICALtJxJbMZulwgA3y0CuxmYi4XEoc6ehRwwAJQm+
zRGovS7pTwloEOSEWykTlwzS4KZRcwPJliZUZhGovmBAnyt7CyT7/UFSVs2uRSBq
1lYdiO4Bh6uIpV4ZgbGxeEcx01o+6ssDJbSSH3Rh1jRAPlFP2qy8bXFawFGbv4uI
/JdlYa/yNOTAZv6oDBW0A7Z9adcC/N27yTPjl5v8MpEDn9oWnrOMcJtfzqYrGW0f
8+WftDV/fgquGqkbMvDqb5m/M3yCZHBUVdykgkvmtFppohNwgesInJHHkqsZEcE+
vfXMcKYFXdp/LWeJrHn8uIxFYHEMYaqKJkeW4o+qT6EJpHxeaTPK9lUxfkUOqOPm
xyVeDPsvrs43tDmNgulNj4uGAjpL0PdkxHBWMvPFyB6E/dm7fk77La0QNJkY4K5M
IA9EtoRvGs1H1833Yo1EcrbQROpAFWvXb/7s/CpMoHMu4mwPbc+lKtsrCwwgb5NE
owvbtLEeocZwa/NN2u3A2A6QZ4qnTE6+VEp7e6yRUs5yvKXErXONjuU7GlofYs81
njYDFByRjw60gffiH6S1jCmPddfCdGzVH5HnWo3rkRzraE+G8JnwAeel2c602m75
LB4k6pjtrXvHOvCkiwTQSipf5ls864iJB5JXXbt9UxbSisj/vPoSkr21seDZOwss
AS/Px1qS4U7aYx4nC/i2SZhir4erE2bGDY+H2KsofKtRsO9gcstgUCqxNcaQBsk4
gxhNHgnS1U8uXGTUD0WzJeoQhmgKMhmRC55bWvrm2IKpXORxCRbTurNjEsZFpMD9
eQ7X28+WX3gh64pCKTWXa+9CJ/1fsNYlKQE49D8T4pSEX6kkH04m8UQtgqlP0lVE
B6ijVqdSkkOZ16W4HVW0rWSVhE7a5j3VUxR+o7e7KhuPxhsmna8oM2VlndEtKXWs
jYIgDhJMTLEIBg1OHFHmyoQonmCIzRc2RdsgpPdxYWq3RLJyd2M0Nb+h/k1inCBy
fKlzF8qo1O3M3R1tuszzHj2hAYjShotI2579iSFpTO0gZX22vqxx5SGw3b4xUQyQ
eIuaiCSc5xGUnaoFDRDVIQ1EblijIUSmXDb3Z+6iH+gdeGH0UPZlXiwfBsw4YLt2
nCGkr6iC7m96rBPV2lHVpWVqg6eQs5fx8O/c9ufz8Y/UJYHw1PwBRlc0HGkEwctd
xnropTW7AcyrBge86/3yYZLYiWaMpXWsKlCNykYr9oUhIczxyue3u/VIXIzHOfge
bqByHzKUnkKRwgCEYpzQGuIYgcdVPmkqK412vn/IMrIRCZ9x5DQXqGjW2tlPWKT8
JUiUFd2qn15giY9KNNbKUJtl6sfQDftb7NN2q0oGayM5CyVdUo1ZwmPoIIEKQXa0
zmqKyEboCTnf6bu6iOFxOiGTRofjJgDmL69Gb6wbnJ1bqidO2nqEgr5oQm0N6OUP
kaPnme2kKorpar6JXXQU4JxB8Xi0DjtT+Ce18KPt5EU8hXsumxbEQSI/GxBlQXNf
jzYkuxkEIjqBRtZl33nO4EtMll0perjPQicWn9QzLkWPp6keXsRJLno1sJcCFEtn
ekrXeV0l9h2hgNCq7/lj0QDTet1wrZff/Dc7ELNr1GwDSuGBoPM/hORQrjZnZ7ru
LgNwjNyzE2QCQwbIibnrNSGrTI6ik2LqW4R/g33vG67xDPPKA2dOW/7f4rQSOeD6
kpkA2Pedzo/Tg9+zl+x8nJxAKGQKQUFrJmcNYWbRjNS77PD9L44HZIf28KHbNioW
QSff+ceqhshzCKiFC4FYWHoLPs2Oqj2Zalz+VN8DAWnvoMf4I8gXhX6Uy3riOiI+
hl+tPp95J3sXHW5SPeVYmAard2nGUaAqf82NGPtzllryqmZMpGA8op7nnsvJW6W2
GvqzDTEICbhNCt7FVmXvgsPC6UENl+AWGvLjM58EeF37yS1eyrt6xklXT+WwVP6A
SD+A1RmO3Fx7tWZbRM6riCkaMdGFRy7/bDJW3sk/VyGeWdorUjDdT2Yk2REgAwqa
zMyZZ10ybUQUPQQpGtEIok1lV2pNgiXFSqxdBvvGZ+vQ5Gn+z2xMGpAoB+3kibDw
6XFsRz/2fdreWQxQiLrLBUWd4FByayFuVsmRMSuTEYtuIMljDaFovBLMYhzLn7kq
sPphUd4TMkcIg+ouQo8NK+kCh0ire1Q8lduT1JYMDxHVAf6DXokvAe9zAiR1U+RR
oy+FffoIGr4I2omIebY+9A6w0/8Tmh6FDGAI/duuI7yA6YAgvoaPWH6So7MJ2taW
789AFRQTk3/VInjRuftSZMYlcGjO0rYe6cgr36pP1U4FrJBNBQFGJ38y1kU21f3q
cI2iuPJeA9nbnrwg9yt3qbFQIwqJ7AixDHpCSGjCpIXd0p0ZXSVkGkD68F9b2UNC
RvwHt6Gfaz2MNoBt0zWVT2cz8qkUo996PhBDFj74NaLI5G7KgGA0AU2hbgSKy84O
bDZlgHIXDvlariEcOrENSppKUknn3VUYMRuHzx6ERc2DcxzkzKLYonmrE+p+4wam
n3lsMJe+tYybWbOmaUaidv0MeQEMimQBx+Jgd4hEk5RbRbv2EXkotxPZd6XgDG0g
1e9rd9ZFcptcBCHtgfAvkFhj+5NWWcI1B6XCT8DfvGi9X5Fwiwzo8fqA/NQuF6lq
82UlHiLU/fTQm1IAdtsqRGg7kv06IGzpq/oyaVVbLOJWZ7sKk9Rzm9ghGz3fy6bo
UIU/K7hjbG0xXfIE8+e/XQwpS+tK6kVXflj9Frcm28ckVdsNh7QOPI3WXOP/v/a6
9zMeCHbYoJgBDNKo2nQwVqJKkrxtxj4h3/zxTAjCUFXHE82aGvN40ntyYwgcUesx
N6Ys6Xv0GdwZxZDz+i9ydBar0uEetEb5KCyDGSuHQ/P03SzW8jxk1wiv71biSOzw
hBKWPkRlFEfbCXjKFdFh7Rzvs+wDIPYpnfNyezGAihaN7Hpz4oIBDEO5JI6tTF07
XDj6VtFmZOIHYg5nBbmR12+8qjWr8g/xrwcf7PGhEQllBvkQS4Xd8KaJEQmusMxM
fbxfvX8OGlA6Ku4TVoaAzzo30bHhIfGEomD+9bAbMSKUUkktsvlfm+eOhbPxn9a3
YQctKEbOdev8SltPokjthaC0prneuzxOPLfOQnHmE7QTsbT4YzEPQZ5DRgYCZPSw
B+JEKulasUN5p9Gw5hCXvMN+rgYuUENhb78Ra/W7Sb4HmLzoN69vxzDYe9r6m/g/
Q8z2LZQzh4ScGAMm6lz3h5f11V0lNWKR8Lzp/Zs2J6YdiUMYh4tBfD5YW5YqnzNQ
bID5XDbQfUy9Jpjl/FI7Y3bbFheY1xPA+icJk4hkzyFIgN8+t1YyrOmoAdNbxlbf
I5dSMSvbVLZZoFF2tmWfb08dHEqmxafPZq8LQ34lXKQmKlWrgO+IPkHg7Tt/cbn2
6K3orOWSOIxx2FWYgXhhYDMv6MtzzhHcS3uLRkknmNVtfE1hJfz1uOlHUdVngJKF
p4V3gekqowYV6MDeZMvQ+XcYedI4nadolD/8wr3wZx/S9jVh4uLTggarx+4qh/NB
aLVFAeSM5u6/wNA2Oy7drzE40GJGXyYWm/Sk9NhTQ6R/TDhLqaueAe4IIaXj9fba
sVYw1AT4TwOaj1lP3U2bkHIHDtS/kC4WosLFjYDb/WQGrhBAw0kpJT77ZDTcB02l
uJNEbGZ+ySsykcdM8WvMbcr3r7A69fJGoxUsVPVLtPRAljl/PD/YhVi00ZzsgXZA
IiUUEhNRwWLiWgWA7/oZhEkFhPpscnwaBe+ZnTg7j4sTCEdrf0oNxdL2EmaPuFMm
Lb0uakxmKWLDUiIs7YqJSzOyCso8OXKrrppooKW++Futggv8kbWDWHOcFZBlZ6M2
tn4dgB54gOUBOmUqIohsyu93HgMZvLZxwR/0V440QFLzGsRIT62MbRy7O768Jf98
SGA0qcpSU/WQAkhXTS+L8RM7ynYuYcAmgvKPFiEUhZDhtpVWN2gxEjeu0qMj9Smj
N/YIBF4fmSYGFE2vG3lGze2G32CnrusK1CLVR187BVapSGYQRELRwj7D+8w2J+Iq
FttjYw+lDpmrlIPiSUtM0/6pAhfE5qsTVzFqcwUXYnEylxU2EzfOgTLHP2CWmgqZ
uE9qTLbFkGQx+vWKPRQE1uJ8wAZduyc6TQnZtnp8A6z1u82U17eFqrphRggIxx2n
AWwGRIhKeTi3OtJzjDbH+xYs7ZxGz7h1PoX0xSU2GpeaHl9l542MsWrizsKPAh6E
jTD7GDdsEayW//tisW7lRlS0TFBRgWyjxA+bLAmifS8feyVjIHKTwrha7lOZBsSp
YI1xBqy0egMAPDzD7xNpPW5XJB9zSucYVydVYiknkRZSg9XFlNzNU9z/sAwg6uKW
5fOV02GKUX7OR7c7WbT7CuWg6UE2t72sjITUNjSJ1mT/ualE2Wlo6oDltY4n/nbe
hPFbDC67ZXPO6t9a9e6WGEzs2NZyv8jyP1B2ER2HVB4KDEJ/khs3Koyl7kIuvhHO
r9Xtcqxz5lR9hUMeUdhzprJU+rBQuHFGPKLIniS2iepcWy22uR+ZN6nzf/DbmLEk
owEabjoYrBEyt29oaiM/KDS4q7GX2veJccG+gTq2reoGXOtSOZj9E6x/BEn0jNj1
p6jpQlE/dmd6S+vwc0/mJDcfr+PKiexHmxdGaCWGvXq1T9kWXnmOBIIwfHwnkDaq
HrSstjZm91CIx+CM04MbO6YzO/eEMqYJPMqQLC1o4t6XvN08xtItRFXD3mA0tA0E
CQAqhrVeSW6PtOHiuKmGlco0r96H/gGaCK4fAQWUF2lk2vuw40oa3ehVx8LYWir6
zkmINs8kQiSwqcC9m8DFfbv2VPR8Li2yoAvt1tFgDZ0nKLVutV5MNmYHAH1y7tSV
FkRA+mnp2KW9mV/n7ka3uOp3wYjbqugd5XSlvW7a0HCVqUXdzjLUDMdvcANcasoL
gp4eFpbw2QlrXb7VYygZ9B0/TOb9nUkJLwGLth/NzbMdb9uEny/27W91cmCjbENT
MS8jfd5hJxJzjT1ZaOSdZF/OQ1v9W0dN7yXigcsuu2oazHTU/Htm91Y/HiyRNGG/
Gx+V6TqnKXFI7EGp701G/QQdnPR3vRFIrv9+W2nceSUw6rybeVpqE5KdnmO4Tj7a
jXt9K5BgjBa9krm7hnpBQIbwf2MxFJ8290gDof5YDvDUbjf0MuSmA5MHbYuor+Om
dfh+BFEIJDyZyY6hOWViFcp6E71yaMLQoE53XD852F1h4AyPJqeDMom4k3C5bnOz
vLz2Z5z8vD8W6BDKS7rQ3TAO11V/ZeygYgkhkemnvmnnx8aKJQojEjidm0a1z48c
6NfUEl6DmPl9K0/RpbszDYEQnSaAb4qzYX7lzbCRv6ZhEW1Wmh/TehhpCByqcnYx
f2kWFECX1lQJyPu9R2oIE4VmEJJ1Ei9jTHFsYUXxe2KAWs+7jJYsFOn+3fdTO7JG
qY7dMk372yRaVxoyguPCwRzDw7gATneNvUx1R1j1k4whjECUoe+ce0na5qRNlt1Z
Pzk0s2ZYqsqWRD14fwENT5sBErhMr8ND+v8qsM/AYNY0fIaL6ntDmcf6wHaWZaGI
aMQ5kbxqjfckI8ix5OX0Mx7d4dFWH/4OW56DEgArbDYPGJJ2h319/cWnTQWAIgvY
zeRXwIdOBCEtykTK/b6j5woO1eyfAK2O2GW9CFReJ09knIrQOx3GNWWf9bK/YCvO
SkI9V+zqBmytLM1nZPS4Q4uDDt2qUSmc/nTOJ+vS/Reqmc9qbcgHD5CwvFdFpXU0
6hG7DvYQygNEa8cC1hKqU4gglvefSYVbptKG/GhjYYKBBSw4EubPGc4n+k4WX0qK
D55y733VkhbNCCwCYwA2BpDmCdmZ2Jnmd8Ye+wbuzLMDsSUbfSJzj2UwXgBvdBGr
FsJcyvJB/YaoY9MR9H6xSxAoQ1mR4+3giNgjptvCsCm/6vQJ6/Uk5WYr0Qz6+YRV
MEtZPgVgNDsUsGlzqFi0sKbC41H+wvadtRkLf52Xy+5yOLye3gDxc6Tz96dBJy+D
vIpOd557yPoWtwosC23a99r22lVTNJPfdHjo9nvvwkEUZJYZwkvIFsKOvxnNxnm1
0368P99vfG4vzeaz2cUXfF1XX5fyKHLeeawGk0AjHpKISW/L7S5bef8HOs4yelI3
sOC+CXw5k48KCuw2N41sZ+feVH4szdZ63QgCaVuGZIhescaMP2aP61LqNhuK8Ru7
8E3O+uXK6t7U7L04MQp5ld5KUQHNrUt0MXLYnezrYYxDxJCwv+c10kMEIVKuqTfn
GnxPAkGZLypDxXRGAOO04mfORMMo97zQ/Klf8Zfn3HH3WjxdHw0KQ+BE8RLqBAYV
l0EM04Bt4tdfLEL9PVZiqAt8HrLF6egZdMinpi/g7Tc8DAJgmZi1T/yCe58fSset
mi44jWqNYRBzk0duzlX1JronnvHjfgpaWKW0qEH7SnlEvwRf90aCsBEhnTSV+S5c
nz/iIPPk1NZeJys+dScPFm2/dJhy7u4aafhNvcw9y2tNARdlUzDmTV2eLOFqXPO6
Q4wwdyh9TmIPVc1sfDuzn6Q9tYiPlO1q43qbB7TIKXjB5iFEJkZl6G8fS1Yh8bjV
xosdKKkmIbHguaaa5+KrmL6bN54gMync/u1mccgHa/WSJL9bOLU6wiIACPjU/fph
bT5RnIHURAOF5b1jPtcYBX15B1n363kvZj3OgCh4WcOcItXOs6i2k3wodGOdCG2c
mt72YBtFvhZvvXPIi514qhTFx/tNJkcesDGBgqH4BS0RrGTRF+2XhZbPorcfDbdM
M31f3VbZP9kyfn1avbdxvB4rfS1nEfd5onWz+zYJf72YFCpK4WuOXwfUTsrrDEIP
GJfEYnmW89smLqykMUczOr0DEoMKuxhQPw7a8lAVJTp+Q3mCTIkiCCkqhf8SdG/X
/NxmBq6NpWqyub2ZtPFPe/kKqoMFVWr+5PhTlTG6lNep1ruv3sfm8KcUA1wIzCHj
DBHosKemPGEQtIjlTZC6FOWaIVQJxovnW2vTrI3mq1pOD/vKsUbeHGf8BUxlNisF
mHxfhUUGgxKoU/XKuEuzT2ThoSTyFFimHE7Ea3jBe4EKadbtziby/z3xwSOe5VKK
45zEAx2R4hn7BvNLL+hZFLglRgjXL1XIqZdHThTLDHuybc8h6QM9NsJwFtYa9+MW
kqAV8hzNGNYakYbqCJ0zzlj6Kfg7I4r6hMjNQPsKGpa5kA/3PuKTYhz/ykM2pt+K
yX5Wfv1KDh1L3Ia4huFZpgsxb+AkBYaesc4NWvXR9jRTPquCd/XY0jshHc7Dh753
swJQ56y4GqFL+DqFcrcUmM1f7vbP/EWoJx4y79v/MVE0EN0hXFMVgl2gErNMzFA0
GT9y8OgJ3bhPZcWfKxYzcYS8mgOYFWX+U8uXYVFa1qh5VNz7y8IYsturFYM2Jnac
ce0xQ+G4UNnRf1C+kJw89zc0fzvy2W/KheghUCvZsGwP+ys0aNfZ/6LhHqZxFFGP
NjL0Y1TYBAmI6kI11eQQma8ghyWFiqHUyb4A3sO9kOWWtSAAd0TvbS26YSiyGyut
hNrN//EkmVs/2EUMsorXwtymWnEd9Z3bgbDt5bU6xYusv7b6jawoDUjG0n8r2vVy
XW+0ndsHCugN0p36f1oyg/RwT+XRtcjKnfB0bk9cAOQ+kPr1dIW3SdCUm9a4miUE
BujBDXv091DhNHQnJXqGwhbMISqMRX7B0FQDkdzGdcGz9dxLCW4wmcBkDRxDEeJl
SWMs8Je+4N8WRGADP0RPNBMO4HyIKmfShGibJ+/eA0nX8RgTuXSn1iSgBvProy3v
e49hHKFGjJkYCHMC0hrOwvemb8kL0HXwmOL66VMp//MJa3FgzG33n64GoZOEQvAf
OE4UIZ2BAJHIEFw34Zm4LZ+9SkZr4UK4meOmLdKPv5/9Hqbb0BFOoOOxDU973VaJ
gB7XLJXA1r5bSfWsKEOXEwBi71En8NNXUi5dMozTH2vjpcSgVmjspFfVASLiFAqC
vJ8XTlFldB3F9bZow6+MSDfcWr+McQohLgwOu8u7HC0nqIxbj4GCr/6h6covfscC
fag7mIwg1iUvE9zNaK73EgunuHjjnYiy+TdLOgv9QPf0bcAtics41HWpsecUbNOX
TL2rxiybqRVKKNW5kuP2g0lrAvz5WbAzC17MrqayO4HtDPOeNmt/ecWzULWahUcV
iYo2PcIvle+ucQTgSid3nQlK83SrGtlzWz5l4GjGYyRLy1zs9HygxYk1Lg8V6QUp
olQM/rAaD+iVJZxKsWpBLvYeesEH6FV4M1gC10n6lJt6ykqqYAp22AhXzYgqaQNP
IFqH5aCx2Kv9TcdZD/TE2HQkSmcDZHea2t5L+Z3XLbbqIM0E0FgmVBeRFJ7/XhJg
1tQdIgwDLxUHLj5JiV/m3xUjayJVDxJsDrlr7wohvm/I2VU0a4xZCZDTg1igXDsK
vsdMCTajknGpmeXkr/ulCT8mEBdHjy3tNrpKCEZ8zN4rSKzYZixxYVVy5pD99eJE
Lb2mWt98hBzBAzEmIjOmoAoHjIha6qG9TYIvwQLH//B7hkcUldc88FC9G5jV5De4
/AiVd9VSCQONSKdHmpUQ4+Ey8Ii4FUdeEdnXgfhLeq17udxdpoDpmnypNhkxj8mj
EUQ1dlcWUT/pBRwS8l22pC2rmxbKSvA8ePHRG3GfKL7gL4Hd3b1UHyHoj3D90yPM
6+yG6AmPaQZ8y7VcZk/n+Y2RD/L85P03Qdgl3Wd2A4YICeJLwsI0ayWCKg/q4vlu
diN7jS+vjtsr21d5yMcGrJx0a7kJUqe7yVKIzODCzXaqo7St7ejaCJlhmfvwuYh1
LHbuGH41aZ7kkfRB4QWz3KI/F3Xes9muqw+enqa9VYGITziCNnjAHdQixzzfqpbv
5dPTEe1xCkRDlfa9TXEV+ck2wzbvM9EXxBvFASlPmNghXV/2OYS4hVDFVTgTeo0m
dOPWBthIN4pVm4Jv+VmIvxFbUcingdoSRVlGKPYUjV6O9PUaTMRGO8VMpd9HkWTa
A3S8xo+3OMMlU8nkOW7RuaAfzXy8+095lXka0po/SPpC67SuUjJL5WXRdORPc+7Q
6jkjUAAOrmdwr19tB7elsVmw8aAXWaluiIgPnLhTyLDF211gWWIcjUOptgUNzRyt
2ZHqHxV4OyukxTP408kd59XK+bRkFEY3oJxgOEkSHmmfmzp85fJfee0tZCCo1H23
CPW3qkRwSbGjN1B4dZHnvKjxXNMjIucciXSi2A1hlhNNWDJoRJsOy5jZa6yRcM9V
krlXluRa1rB7FUY5Afu4s8GMK44AMGpEyKDQPiahZ6W0sNh7tfLtDXd9eAfgbGOK
E8J53bxL6YKwY+dlRumI7uYDd6K1QCD/lfBGcHnT0i7q/G9PouJc5rYuUnT9hgfv
7yNwst8dRgtXWrbIPosuiGMpZgyvTmMGfnhMccuqG3Mpamyw5oczCOKjM7Fn9qGq
CxKSm4zEf8+RodTuo+upoikDNVHajOIGhCNqsRPU+UqZL97M1zJYbkMQngwSRVpp
cGjyohufL772xE5JoDXAb9GHFa5GDdZz673amgc6vtmVO62pCYJhSGxx3Ge3ySO0
zpyoMzblKkjbQzVfWdKlFA9iVFuPA/CFU48Hbf+WmvA2Ip/Q0/LP58Gsb6lfi+4I
MjQPQ5h8mWLYm4GrnG89vW7/0eShnpWLbDkf7mS8aZCIcranCu3TEq6DS10yyTgF
eLthyb+s2O1jJWY+a4f9Ya0kmzCYzIcE/IEjkuWjBR+WY5hmXhH6gieOBEU5/brb
1/3jqE4UKItA0bWbbRygWtqUdlRlHUPWXtbxLtGWQyoKMJollKCeQ2ZYzmB4f6id
ue2sZTPCOJZPWoMyi1KjxOh/2e0MrqbV59rXD1GjFCzdTZSuSS4sUaEA+edRyY5m
xU3qOvQPK64mIH6k3XXq2Cn/d85CRy05hFg2FaNPO+tArkp87/12+McZpNhctUDh
WQrKlVoMntCGh3jo/WDh+OmjsJam+DsH4YQD25K/90EhhWVIpqnJfOkdheRB/kTV
s+0jBiWXucSb5V0eehkcVWps9cb6KOeS/nU6ylt5h9w8ueNrE+b9tdOfEqJoxrWZ
IyohSSEqhzJ7vy/5n/tc9joEoSYu06mIBiGZiKCyj4vDroqZgcVXzwqjTwDQbv7+
RjVYGiWCKxHhl3QQZ4orYm7EItwje/l6YL5mPe1pgcCve0C/hUKk2Vd9SCax0mFy
TnTxdaTRsXbbjk2MSY1WuiRgTMeTE3H8pEU0O4fLjsy4SbaQ6RSJJh/AlV2a5X7m
eCjI39dwin7NXZWnNlXPwOfPuQaX2Ijh3TH8HJze2i0et/SxQ5L0ifZ+qXvvvdDT
BqJB9k1QsWdMIYNx1b5f7GxBzxLDTT4+g9NtwdDjIds0eY1qwHZ9aaLME63zAEW/
7RpLx+sbOjlRqkfWamWukFFyKC3XKrL9564RulNoevrXWsO3F5WZCezhfbrzgzP1
+/whbpScn1NqsWQc3absj5akDX7XJKzV3sZvqToSFP1MXJa0sLdesCl+PeyMvnNm
7eOyphpQCkHBxPiESAvavk/q020jz/KDU2gf7xf2lvJE97Ut04cq1btPiGHo0TjH
MLK7FKhpgrQeHQzlkDHtKboVDXsdR+HwgIPJtbC3kwpD/UtoHXtcuyITt4wwezVZ
iIOAyw9YPyTCto+GNbuII/1hWaR/PH6KrhuodeI3HnCOMM0KxXkVgUOdks3GV25M
lzjdRy9OBcbULzeEtcOPFKmJryxGkVKokSaQ8TV5JpEOZVgu3WJp1fd/h06bvzci
zglvuLGR4kZpZypqP6aIUvVrloHskhniF79w8osPHQHTM06FUL2EckRxA215NbUq
rYl3cJojKRtAZhCQ4wjbaj5bhiOi/kjbQgmS1kMBgs6OElvB9o+Dk2jGcS4Z+Fwa
UiAe3x0yi93lOyZX0urAsq8YhmWC66X3jSq4p1jNj8e/uARFNiu9zffFR5Dw1SLc
1N3ntUzBOsUQJFRIq5moJydRwwxE/FN85/Vm7MvlETK6Jfx4i6m+4bmMSFdG3ZKU
R1vakSXzjUJ2UbnG2g9gMt3utOCTWQCFQQe96MfDydity6r7aj6rrnIj5icf7+lI
nnD/TLWmc+wZehRVNEIAjNXwKWb8QQ1Tmo0RIztaVznr0lFCZR+Q0jdZdIc9ll/B
n/+NbI7M/vx/NQCXP0kdJ0idr6ePrAVM6uTZ1dC0/rAwMSP136iEh67cFHr0B7g3
oTbSgzTfG+ALCj1VPg0QrwO1RhAOLSSHtA33aH/CdrBXYAuwVuOSd5US7KVRcyqE
PF3lhXIvXZu++atHhDVAjgpTVmYir9uqjjxGQ0rNG9DNPUrroj03N9D5nvAmNH/g
CiTH+rv4f2pEYQIrfDbsk8BPkZIysqleh7ExfRVCqNTCmYDjl0iy51ROvoEWjS1+
LLZtxuSuXjbyQ1i9LyNtL18/FzApCF9SLxFZ3dD1DPwdb75yXGlSB5cRnQp2vKEf
+8PFejBXq2AFj5GoZv+ide48sas69+pDdEarWg2YToB3YPwSq4u+UmGaPG7QjhaW
MWIXcFH0t+aCW560eYVoUdayr7gJNjrDCgFbFW0cJKxtQjJgZC09fJ6JyYMbCFCv
7ggsEPgHMezsLoi1bReNui5PplQk0NFg5hN4nTqNIj3Tyf3t2/1MFdHapDIMlwx/
GFbYPszGHoh/Sc8oZj5JRCDd5APPVoZ+X/S3z6zls4Y6RX7Y9CAG7RX6zWF4GQa1
jIsdl3MkdYrhHP4CB3+OkvtHnJQNF+yZu9xXPrEGVCqMfeoz9G6KdFDRo6PRBcyl
cf1eqtCdKscG3wlTRymULVmhInWg7oLZm2gMNGmfBwWWsyp+M65Zum4q89tvAsS1
d7NRhNYPSdkjfwP92qyM7YDnjmNsR4Tgstnu7sKnim/rU+HsxM4CpiXEBUrdB25a
6G39+QHiAVGtuMvH0/oGPjJPCm8jZlrg7WeaAMmMDTxw9FKOano84s6BsVAfWiSc
84TKA23Ne/n/fGDzWRoV77TEfSkU73oVRKAoZJAX/tF0VuoobSZZnPKmupqeL/ZD
oPxSR1DdDqHLGZhOFOjV4SZQn9WouMZ1hf/wbCw6wBj0VQSbmEf9QbrGC0EKOv/Q
QdQVCXORp3Vva9OBQkw8K6OwZ+NJbTVO22own8Ub5o/z1/svBljfgCl/WgprV2Ne
PI3eek9l9Bd+teW7n6Q+xL+cG59Ay3+ARWb9R2+xK2ofIzdvzNUZDq6mVhs1WDWC
pPBj60TawhRf0a0BcosHHmT+HtSHC03GLsxVaNseWxcXRGO25xwo6AJzztHAp31g
wBg1SBbwC5J7POkEwe6pqjevszUwpWGJ6eNKOqLbf6xbCzZ9rtMyCjSuYrpWvmFc
giUgkGq9iWkv1w33LTyvkqmcPnf+r5lnz2XxlLNpGNoMGl4d+YfmeILvw50NnDrm
uUNwtoAu2EJE/GPFTsBi8Gh/jHgeoXZstiXcaPVvfks2Qe5dZ1xTuZgwGNwfKRFl
/WYPfE31qFJ3nlDwwIDWCtwkPZDd5cX+lR4LivLqgGkcLcu2dyRiRNGTuePYQeZy
eyZusxVUcQtBRPEHvzzNOuArtH+Tq+2QvJVJMLIG9oFUyhWolHfJpEcp6PxPygDH
J1y8YTO6fpuuu8BUq/ih/0khvctK3FNO8/FDTbCzipLJNfrV+h1yYH27txPGEX93
iTFSJYMfFI0rKAilht6LcXKKvmy2qCZMml6IWPLCgr8TfJ1MCvvoUt0oeWrfL8Gv
887aR2BfcrYzBwFh3PAm7oz9Ys1oXmplPgph5AQImiN215FknimAKp4ykXJbi0Dc
6TX8BvLh/Um4iNll0EpepO9TYzAONwHjmkmSrKaWWna+dcD+ChhWQJs+r7v4N4zG
DlmcQ2qdWLLBXboUTsY2qDQMWwd4XRriHNytX5dOaXoeJM1IHHyH1Ni/LkIcGhVV
2gqpAy7xvePVSCucKlQfDI+XjkjrKXKEKaU/+9XKwKvG1uWOOld3TqCpJmuKiZBZ
1G1oHeYtlTQHkDNkp316DvlBloZZG9HgK5eOYuCig7wDyA/SOS8LDHbFZob0dpY2
c6T4HwRDxAx5GlsMI/XtVmd6ieBh3Gac4zvRw0UITDmio3mBSBqcHpakJ9XRL2dw
M28p+RQKFmEWqUh/q1db7Qwtb5XVVMbDrwx7lO/epeOIwqg5AGzlv8FZCK9tam70
Eg+0QQCuEwFHNlZg4FvUydlLctk9SchUHwhmTcEqipYMAx0XAszfNDE1XnaKVXIv
mr/h/OS3j44s6cj5IFDK1dGifCUpH8baw90rKhoqmZ4smvXmnd3XRKSlUa0dh/Sq
bhfR9+j7fEDHSBT/XBYyDSekSD6wC7wR+yYSti16faNtFfyaSXfLF4IvAVcsrHKW
Lfk52rG1JPYywM/PRp4HG/kvYLBnV6+aRtnDpzh63Ee/Q93W3Q+a8We47pIbpVpA
Dtc6bqkS+sZ+4vcKyhrclU4Yzg49FvqELR5qRchDOlqkYoHfnP/Axr/6KpAoTREz
1Pl0zB3R1RWcYuHtZLJMJUJaP1SVG7hoMXa8avoljH8cvxrrCyybZFrMFACoxlnN
v4iHWvcReMFRYZqH+8FNC+ENLxpyWOkoOSDozmYQRmiKRQwTowC990ql9WxGz8O+
kPQPkmaCS9K3t3tVKeTNLYEpktsr2lbpz+vxllJAlcgg+4dfy1vde1Mv/BJr9/Hc
QZgA/zOkuLvkn+b1wHZODHMewYHE6+fw1C9E10YOnLyovKzXAFSn8jllN2LGczEJ
R6LCitGy1PVCSKUY06NsUN3vHkeSmJSaTsCF6GigjvERNiZ47pXN0NZmkc7ADnPn
sJvuI3UF/o27rG86g/sGPSWEevpgggk4eS4VB3vKbYvvh0Gi1R6tPtPXaP8DYeoz
Y593pplLz8e+WQS8A57pshLnK+uldLkYBEAc288N3AA04kNTkLB1QgEEv6Cz4kgQ
lX8y67as6mRNgHb36EiZ7XfV+gjDgEzchQPfUplTY/N5n187vXwlmF6EzjWe57lR
sEbXk0D8vPQKWjZG8BNv8wO3ltAs44lFQZLLGYf0xFhIVgxLi4pDCnutZqpXOi6c
Cm8fbSI5nr6wxxk6bdBBXcBUa2T0MDHRJizRV2i16chYJUg4pFn+NjCLNQUHdMiV
pDtj6uAqueH/23PgC6xEQRQ/rCmo5xoQyERn49BgBzDCW2VavBOBHRya9OuzfxWQ
T4PUaDzRoe49OhMEqGcDz5l3JrL6m2IjO924McecG7l1NpgvgjdxAg9MbzKDb4FY
NsZdVKNgNM6e49B3puxVxg1RgT0/A2d8WIiOUR7t6eS6285Pt4Att83WS4XhuePj
J8j4xKwhCUhc1Ms9YQQH40b46TdhM4fJz5O4Bl0GfiN/nujWOMOmOOEamdX1vfoo
f3z24Mhqayj2LGFYFGGv4iZ7Zs6rJ+g+HgxhHUMnnRo1AyUeNTQ1cwufVPhLoHWj
SoSNmLxDyYFIWrLOsvhN0PVIqrZH7OwF6BnMtXTBsD+IoEzlCBTPb0EG1Ivjah2A
X/tj4RfpQtHhC8l1GW0UHLAj+lATD+ZxmbY2ygdZH1CqXW2FTaKSc0jui8Ypms4L
ssFRaWPfzARomU26rif7a8cblPiBjUOQaOToc6L6Pf5tWOpB/GSOFgT8LZqwTvV7
rCDWESxVUFWUWMl7nVcjiGEkcBRN7bxr8y4i/eZ2qe62pX0msixIubX8gWBYAPco
StpneUdpmVjDP40C+aWlvp312PJ6jWjexLr8jsn3Znnl+feK6+zUSNZ2D1pmraHw
/VOX+BPCAKl6/XoJ3dzg8+S/6QCcpFKqez2wC4TtzYOPDNO4R3Sbgtco/4Y5iTEW
sDol4vf6DegomFJX3u+E59AjznlQ8H6g9H//WDh4JPgTd8ZS5bn77VTpW/yO9dYq
NnEO6jQEK0IwGVrTqGxIGScbVsJevzD1VdtuEt44uVt+0wuv22Ug8EQsZrWEtmJz
E101MYWbPBv6woz05qtXHiEWJYc2MbR2/drEm2U87iApZr+PlntpEXsawT6dBobt
CcaXSfYJb+Xp4fqUZrgbpuMQsEG+AkbBvqjoeL96jmhnR5nE2eaj1lYi8JomwbHB
g6s9UblQzlfPHMyGV11UYhKMZlmeRtEEyFMnJjnXtS2JrOjcI6TaTDWRw9KSI7Ol
Nr4tNBsLusOOOKSeX9lzD8iUXScGFS3zVmf93CWNYmPBWaGfq6q76iVJxvh4sGw2
+EtJ82hXn3T9wKUBqzgASPfhdFk6V6/if9oEnbQ6cM30GBg+NUt1elzgulKcwCo2
46GgeB/GrueXjFJSW4xpes6xnIRsCAUjQjqpDj8xUPUlf5ktEg1EfWibuw/JTHNF
KEdFB4mQ9yNvqDRH1ejKHU9LJ9tsdqzrJUvDyDxmt9P+xaUQPKi9MOFMuTO+Nghv
F0Fb5EUgq8ZQAaoNBzrnbQzcF6K+ZhmnPCjGMYXInNfDqWtvnvaCGsS7xOtuGjFk
E9mNxF3/be4YNuecVQ5DejzY39XwyPBP7h8KP5n4H5mln8Jq8GqMGzA4RTcbgY3l
15nfQKciCEBTkTc273+Wm7HBeWy9XvWq3N6nK27PzPVT7HSMrpNrvHnRd2Yikbsz
3KcaPBbuXkTewNgJOq6TNPHancdptyJrjrQ49DN2dokU3p14pVlZUXSH16UzJdYZ
LbjFfDTQKGAJJ1Ya1QymoYccXDLOa6dRvDjYf+6XuXtrKIn1TUwWyotTLgutLVEM
ybK547nAFFP+rPkLxVMt5/Zs51+ydvqjATHGA5RUGkDQMhz67wh9J17Y6a5GJ5UC
8qXTtov/yXZV7/p7VjIrF7nktQu7OWGfOIP4yGlijP5P7/NVrji708592BTMhYlX
9VsblUGJ7650uqAifxAMW+gpUhTL2iMvY8ZMIwZDLyg9Kl35UbNRLtpi8sygblX0
82KrV5jy4DejuQwHyFYpF8BYK79JSU3HHU1CYTCLyXcLxpV0YKBZeXgz0HXtz2SB
Omw6vWBYdKEqr6hqEiP7UrQaL+OkN5s/S1zgQ7NkBjLEmy/28Vnek8vkMwnX6sdi
n84xZHQmKOhz9E9t7GDIKGQJMjybr3QKuAj8ZXr5cFiigUkTJrYlKD1JQ77f7pD2
KnETTotm1yMZigLL/93tS375tHkjcUNLFz3cOmuYa4+vkJvz3mGjnjT+mG2fNBnV
mdZkvsNEMsKoPtb46aNSeiWvxEvIp9nHAb4AuoakGNZYjGP92L/XUPwEgY35bdG0
SG/KtiCNTmKoCohfJgNhTFXJQXRi0OGfs4MOH0GdEx6M6ojRP6zzU8ln39z2L4l5
MLIK/IPCXBuLjw5m89bJBA487g/Jgu/+6feFHtOC8ADr/6FUp8/oaBNkFSdONn03
2tnnl0FdHrfFwt7CmM0mbcRoU5FyNG+xpOQyt9ty5s53Xp1R/HtE3EgRAA3R9U/j
EES8NNdFnjMdUkHh4z04gcVz/LPMok7fzoRuqGcJj+vfBHZ8fwemGS0nhV2ZJfgP
q991Tl8BJ2ikxxGv7oDKcHqqBkqLAxg89fcfEpoJMhhz3Rnhia6fU2QGl0s3mK7K
MWdOJ+DtQwvccRfHuBIUIKuN/hSCaTwIR4qOCd5fTw8RzMSFaS8cXHq4yRXQJGGb
iBULLo3M573eH60RBbRCDKu395d3Txig4kYO8RRC7tjJBOpkSlEh1iqlsVVei1Vf
LFhXSpdeKAKnADeoqaDD0qb9qt+qFRYHUL6w+k8VGrutQf/eRnTNvcmdtsGkXlxz
lvsJv3CSKiZZEYNGqDvInAZaffzaIjQESFsu/HUVJmhDK4FJuaMlZ/ORFRFpCjhZ
kfvF2TSdNSXa7MbL25XftYTcxGcear67qozJUVJdWE7A77C0ir2zO6mtgEKkNZ1K
Yj7BQj8seHCzC0j5jWsT+2wVYeKnpFRbjQp3weSv8KDQTpPdfjC5boDrEdJCl/8z
XL9CyestgRcWzpDnPnmONKfY/BWMxzkXmexvM74Q4cFBkNMWUW3zgdU5D92rAyKM
XmJBIHu2yFjEkstkxgYCUf5+Ymwg+2KBGNtWaQ/KAfmiQE11ilp/w+MHuxN3YuWd
sC910pR8wnQcgrfbuinMP5hTcK7cSY8QTD4bUIKO1/oi4KOZaqMui+3ah+lc0IOF
vZXpSQ5TtyUMiJRn8j2Fz1JwObRtdKwQDxBRbmUr30+i01hUTXdSOVFjezJTLOTz
mnrfF4lT1oabFR8oNfypzB67Me1P4Dq1cxrUufJ5slgbbDX8iF6iXiHh3w81jAbK
YV1V6NMBf2cjv5+6v4E5vZVXMTRQwGAXzJWx7SQUYa8Hajt6imZ6SA3N3JuOk7ko
qjv3o0dE30elI/e992kLk0Fx2H/rOCmhGJOsHoDA4achLxNwTP4RHY6KFnzsLlOc
AnluUd/DJEww7FUAs3t4Iax2lqeDWqMkzaPUXr7Xuht2e9XItByIXAKi8DmgI8iF
QGY2D95nSos4tGCAXKxkW0NJBK7YI2a9nuH4k03r9Bhr1jnN+4H2gWFhCtonm8hM
fIuud3s/fzol/yfbFoy8YbODxsvH4ZCVjR1rahis0DqKl25H4hqIEzpj4Mom1Y+z
QbFLM3AfS842exK+TLuvXgjPIKQTsburw2hfagdP5C2b3p6xRo3N2MaTE4j6GivQ
lv/WOZ6BgKymaG7VT1idKX7eS5m0oCGbh36ivclvZwg3Ub4Slcm03g1tXknNCHqA
5o3vLuJ9i50vdA3S0iIyRomwSWXngAO4QvDB6kVER59B7OFinVgCFL8G9qWK/pFT
WBtenwgnhOhqWJHkH6/F4dk0oZzmwl8BQfNGZO2YmZ1wFd8YkJKPg0P6UjuSivga
lCp83/D9cNPb6DtsPre7uyJrbn1FXqVmvee15U4GPgmx3I1s+KFohb5x7pq+/31Q
Mwr4fOJE0SPTZMrMQn+Bijt4NAHi0VTS04scMkyNl8uyp5W5pOzhVCDKcuwgSDvE
rQy8P97f3TLeiKYPS3x8D9IPgzYFqmd+QzGIxTccjEh4V9hhplYT3Bt0eywFQeLx
wjyhXdxQBVjPeTTx+d22FfoDUvhDeQ/PtjEY9ArgkJGluJfz1GFbhrB31DdVDklh
oK7cRcBIYe/oKiDC4V283vJSnbTHQm0HjevusCazT7M75TwtKme81J42PA8qoogD
54zPmV6KWX6l8H9QGe2wejAYXEnpw5qFQxZk3FDnpaP6P5PCb9FCKBDoVOCi9HWJ
fglQaNhAxQU4JhfVOCbZugAfWfkPQUUn9mbIO1h/gnnEVK8Qvv3+FD9/uvKGlhR5
n4uA0u9JqaBhGPKLoUOogDLJCdxz5lNIJlbegP/G6qFQXsQ8q+VITgDnair+3b4L
Fe3594w/MTKpdtOH4aaM0h0LWSNTLCLCuFYsd8ce9ucMrj36f8YJgkGIshfuzJrW
HG+DrqlhTHgm3wIYJcbnH5p2dsLqZEbofoh4T783Wj76XWP11NHzbnAjzFPHUYXV
HPNTjM6MkPonDDiqJK1Om9tkuaVjbcfQKHp7f9cE7Czm3thaI1MUujHb5e+n3UGc
75Rx50WEK56OcarWDknY04c98AeWA8Q2qIT1CnUzCd1JG8LGYwUzciy8XlMURewp
rBhhdUQRh5dVjbLj0OmU37psn1oTfIaCtdj/G3TaWWE5irFDJBp4uQn19oIXwC0W
d0qPdGcuj1evbSFnBpS4W2H2jyGF2ZIcOE2tOQ2u34H+uYGNF41zXqFsgnGWFUk3
BJixKPujBQbiBc56G2rppnxJJJD6h06k5KhGAqlrmtP78mWQ/1jb146iDRhU3Lsh
tZOPHiFCZ3O++1OI9KHo/WPVp/2lpNWYTu3Drq6Yx/lsgGczjU4Apxq/krWx9RUw
sk+AkQqZwBQIx8RmRhKMzWFQ5jwoDxTz6mlBR0NvGdUeguY3zQJPM64pgpbNFufo
ES4ChjY+3R7rK7TiwtjGWhEUpuidSRtOUnpjKh505iDLYyqsv8Tg9g+bRZZvEVDY
ZSb/wtSccwzECCtSrkrtu0tMecUcQA1ADVoQlX44s13cykG4mipT3gVL2eA5Gu/i
vP+Vd6YgUD2r713bQgSHPz10t7W+QwgxmCRwA6qveRXzO2TY1iCPJ87/8Y7ssnsq
2bMj/4wFAiPXFLEQG6VEznB4XQe+vQZxWS33CWZsrw2FWJj9zeZL4ONE5UYciXro
okWvKiWNS4N76Anw0WAAJEqPfxBDaYkHWJv+25daWi6zzjIg9E2BpGum+5PcQMGp
SE4P8liKFqap12i7EQX2TnkckBhU2Zyzo/pVYtsvn20VElCTQxSMptHORXe3B28r
sLrPD80vpXz19b0Mz22TeOZzC480aimtdUFjLxoNOjJr482A8g+4MCfoUzx6C018
gmAaEqY2FZ4xSEHTruHWXKwfIz/n1Z4ZmX/I1DVo33GWlaezSYsAw+c5wCkqLVbT
ZlswjE79htAkw1fxUn/9zuvvK/q8wIxnHccDsYyP8Tu7ZVwZVvN3Dn7WcQvChi3/
gTt3J8jVzmSGgSdUxDK0OqqmUu9DQ0NWdXpUOPuQS+8cusjMxfxnxX4gB9cdh77J
4IvyEhjz5mZHmBn4wfzXrTCad1FDWgMWJzux7agoPJNGgd2uExg4Q7pR1VVh06g/
iTwN7MQwdy78H4Xl3+0LfUxY2P4JRKPWTCvQhuSJoXKXiaKtdyvrDqimVplhTdnc
ooxr2kl7M+Mj51tPl2GPeywJJ16giujUiyamgsm3EX1NNPrKneNPuaBKtPPqTakj
1TPokCZfaT5+opl6thd2Wb3+MmlzXs/GCGLvDKXK9eUT/rvAXh01OutYMP4xahCe
7WxZid0h4Fzv0zCCtXpKKNuXfCWTiC+VfL34G6x7yXZleQ11W3HYmxYEvCUDbVZJ
BxCUBnRQ8sGDzY8X1oMchBgBsbRWqpiTkTSDGcXJ2TDlx/7UJSpdgCvZC+Xjm1Nw
yCkJQuK8JqUhWyDNnyaBW6Gj3YcH5RsD6oygREvY4tQL7EK9+Nd2uOVYcP6OWEVs
sIuks4TaCgf2dfRo9vWw8gU2aAZ7o7URDYo8vAfkZmtfAw9w6QFbl4YMPJcSXz8c
tnqAbxkaht5o22BEsymtV7C1FnbGCRgOkldWzgyVwhKjqhSsldwlcr8j63oOzPA7
p4jia5bknsPMVxj7EbTgf3+6Xl7lwv0uxqSLrkCXN++c25VU6Ic6rAS82KY4cmCN
QAR1iuDCo87rJbSQF4HNf5+0UhfI9RYZ+Rx7pQZiPmmu8/9L1XjX2sLbw90pKSAt
Z8Ze9VO9xIJJuH2pfk7KTJahG0rx3V0RjV+eNxTJ/brduHVDXc2NowCqEhq+0+mz
nDI1QQCkhYYd1s+XRFS0qg08mg316A/XMgAoMBlykRDvR/1vgCMHXw8Ch2kyIVZb
Lh01011GzdQfp6NCtx5vqhzjH2sHJ9GXRmZkjkhA3vXfbMU4CBKln425EVTqmCZE
CiV3McT62Li8MAuKwEywdXwXH/e9FtIEKdTuMdK6Gf+ZN6G6SxPkykxJ+jUUh7+Y
U/m9gcmZb0qVp4MbqJroouT1BwZfehqN0zk1gzn7bD2A4pHhmgCtf+lPnzLu/QKu
wyYdYEEW1YZ1eA8Bb7+pa466yOYO7FfDu1fTuv5oybN3NRAg3KkhNFZjyiVEtDeZ
cCMKDI1PdJiOAg2it5zKR22Lky3zPY5+8YQFNItHT79NqoB3fRB/IaGgvVtvWViw
PTlmHp+/3fJs9r5iH0NsVQdZcxBjHAgBCZoGGSu+Zgq1yPIKHielNvgnrZbosAKY
HWaPpGxkwLSUyOIljBDHzrhxFg49gH6woklfxY0Lb2X0x/8rQB1PB08qP0OgpMka
jxfAOYxlD2CtRMlveITtdi/PxUZeQEEK3PDYyO/b4YVjOMtgzzx1kgBr4dXkFi0s
iKyyF2mJVsFFbPzqj1XfkgbCAscDCEN7QvM/e3PRRZ1UVRI5G9Gdal0dGkfxyHmx
WGszz0DjXwMNlxmnZ8qYfd7t0jAgzYeCDR/UHe+1N2eB1EcDW5NLRIRWq30nTevs
5whk5xzI4ZpIqv7yP1UoU7BL8mx/21aT+elzgaCxei6I7h+jJi6P0tjs5d2aGhSF
OBAQvy9N9bo0xEdErWVbMfWFwVnmssBf5TF0Q9GXg1OP5c64bqRrAU1rlxrgLszp
EsPWdmx0ZAG4Mn6hPswgK6lTP0QticdyrhcAat+FMhG9p65Pj0UuTmu4mJYrZ5cM
wxv5klu5lg0Zrmag6jHp/Kc7hs8APO73OsaiiwzCdWQGiP/T66zFlcE/Z+nM70KG
SbB2io9sXHd7pAj0CnmIfJmTilYuyp1x4i+x1yYeCSui3yGS4zi3c6a+VUu3sIPe
rGcCtnnDLWRZRnkpH/c2fLLJt4MO8qiSpsI3buD7bss6xwOdwOSQIkgHp8SPIJLh
cOOt4bTV7XjJIQPVWdPz0BVBs7rtCGVysdMjfb0AtExg6iLCo2jpKSR1VAQEe4l0
OBLKNkiLbh3ZV3seTUo7ulk4LFgSUqqvn0WhCpcYpZYqOLHrN6HhUq6pE8dSB4u8
5e8S800S4jA8N/rkaSajb8dvXF787PFwwSVtpmPHnm1NufSHLNufzBa34fTZWcq9
glaVSetHjfkPoIT/7qY6AafMpdvCwP0gX7FANvfuSBWArp0KbzOtApLXEv48CVNz
8LA1GDsG1hWSUPjYi/O9GqjJ2MtSJHWr52FTosTK6CgGxieEFSpc9tsT0g88XM2r
uY6nIIBS54Ad3FaXSfFhp9I7XCOnEfNgHeNyY8CxhsZzX81hEQcYqSEcf6bPMq9P
XUJqM421WRBX4DIwl7X4UmsMCPZm2O5VCAJOQL1iJCnqZHH+3agPBJNE1auCBJDj
6zzTLrrmR45f3pmgsRfyY/v2aL0E730dPIGkkI55BbCvxtJCceewXqZpUIvhR84G
f7fLChnZPaI4Y++iyqhQDLsbdAjauaUBDDtXUI8YoTfO8ilQsg52Lu/ZGa7Glq8k
6PRAGfSUQPC6fLYakNqKHyEBrh4uElCGpQx/mKWEl5YIibF6lUElPH16L7g+UGBJ
Cwbi799HbWfGp2+v4mOALddA4JF4KwJV0Tg3qu1/C4lgn3glUT+cH2LW67Vaqotc
fK0VGzm3mg+ReKeP2WOVg7YG9l8AgfNTwhAPF8yrAadzuinECDKtMcYjT7HAsxcO
fowDCTApXeaTK4zM2szJ6v1KtUOIQpWSHveFWcZ80+ZI2modypgka7jybX1kFPEp
McMSmrw9GKe6KQnLUhIKwOtuYcPIn9mkAUoD72jmmtiGpCGttfY1FyMchVL4Xs0j
dqIiQ7s2XdR7EViqvFTMab2h67jx6S1ixnar7Dek3giAkxMTll4lZx4qNNuqG9DX
oX5QVNi17A+HhVY8NbdoGxQp/vYIj9la0uOj2siTEceU7qbqzQV8iEZntrojAkTz
YsDEEzsyNpInqZgodeQusZqT90bSO5T3GYbyssa6KgzdTf6oc4Dl5u7EuV/Et0xL
9NrUWxDqb8WB92Hj1JuzXwEcINedVlLvPitaGLEcWo/RNyndFvutCmsGjW4QPQ3p
sgX1S9G+qryRXPm/Juuu/jAKupQmdwqb8kDNGNe6QVQMQE60Rf8dD8b6rsL8uhZ2
c/xePEBv2jDOX25eFlLYQH9g06PSdawfRtx5E9cYWYdUXhjWw3aChoXfggNM3UTS
nazGolMcK/rS/E5QUaYZ45kITEyVRmrUBD5z43u/KYsGtvoHHygrXJXilPrk9pnp
TQ4+9tH07DSVEBCKWFqB4CUUNJQSEEC+JQzu2jf8elfw7zyneLYER5B+vCD8T5tR
pzZhzz1xchC54NGbi6XLEBlQH12vkrLdy9A5g4beCG7qGyRtdyJODiN36DGDU88J
xMwTTu3nPvsBbOMD71CTvw7uEkrqcn6hiXkSs0t8xJUwfyT624gbdeYoOLjyx4Op
LnPCjgvY8cn8ahPhDQSh4ycXvcuWJYoHThGwxzzSK5Ro4Jr5vvxV8hh5Bwp2XqZu
5Zat3gojfFjNQw7jQR2FuMqgALaezULBf3gSqd47ghXY+IbRwysgX2JztJ2wiIhP
VYSksnHTlJCkS8crPKUOsEboP9tVQYJ2aJnIn7f+F30wnVN9VTbbg+eCICg0UFx/
TxZPsEN7erb3r3m1CAQ4yVuiSmFgeZVKDQecKkHwS4TJR4ZTr/HuHJisHvLDfTcL
mLHUzCjAfgxqqXyZX+r2hS6V9W5Sn5Sc0ex46gA69mKSRt1acwLopgNQPTzd8ePo
CRCvffAWZU1gSlKAw+sMqKY+BclaJkLHLkIs6ULUK/b6ROGUIxWIWvpGRE1vcoXR
mGw7JANYMaDxUrUH7wNR3wqL/BGr4L0T/HdbGoojr2sjaTCcGlE80b1c2ZENRkAv
hsNKBjvs9Uqa6ngSu4wO7/+WQGErDAl8/kFJefBs0iPCSgMuaWczFkimV0+Ani2o
0zoK79MBv2X1QgJMDGGXERU9L7lgy98AW1QvxSeDj03J0SUqwDvnhkLkVJqDcK7I
z/qndEpsJEpKoWlX3UERWgw/eeg3sLz+GkhLoXHb3CkcM873nWyJMfnttVTXYl2r
H3af6c3LeJqlloydYVB2l69YcJ8zWgsedhbAtRzn4rHHsZapKQT1+/oHvrFiXLPP
D7mSDiyHHE7z/kHrRSCMWXbQ3jQ6wPwtVPUlzLFyliqGeDpqWCHhmzoVybQUJdjo
xc3+qIJO5KDQwB4OUxD+5OZoWFpnIGxY2dYCShXFdAhzhUeeRNSJUVHPd2uwpb/g
No4Yfei5/WEotSuXh9v5fWy67b3YfYHgaKehP50Wd0+yaCoUw85RDicxepWRariJ
sTAi+qZKhe4ZrCqG/S+XyMc5/QVd57n5TDgwCDqpNa+iR+k81Sm9+lO1BOraPaFH
vzcdqe1I9uNk1nWunRrgwjPY/idbAVoqp0J90Ol9HmT/oygNSiGsKGVZyAiZWXBP
b1HHl6B1f2GUC0A654U+SpGNoh+/qokT1AfIboyD0+5rsAJmjf0i9AR0UQ7XbL6Z
Bwvaz4b1doGHE4FHW7dUPOeh8h+buUJth303ZfWLBFcO01/1Rup/0R4qYaPgXRUQ
7iN7D8G8tFCjkgRRR0+ZHKOb/D+Tlkjp9vWqoFBqLJrUHuSMFPjYiJGnEAU1/1NF
fmnX36c7y4hzJiA9LEa5E7tn8LNNsFgIc8l4zExRwOYmGvnOr5AJhcHMZTr4Vc8p
xT8pmosEz+80DM/ZlTmnSlKgUvaroYhiSXfvzQ4IDD480RPRhLOXMEGKLr399qNB
qeJ0qWVebc/jfRuoka7fIY/Q0HbSLEoRJBscliAAm5GtiWW6zWWtjbO20/VnHQf8
l8bWtsUfz0AwVcnAGzVQYVHofDoVJf2XUGp3etGdUxq/Yb30w/AB/8xmWzOdTlKq
NuarG1z3HNpwrhf749qb+lMhb96R+tx2KvFO+H+rMOIF6nF22EPV8d/0l7GmzCwz
rcqe7GdYPrpVps4jPw54J3xN790hhP6MK3S78WOABV4bOamhoolKV+PKB/uAjZe9
2awnn8lmIWTBU/JGJsqIGMg1ZJYdZc7xJzumWMWz5rQ06jp89DQXXvwhXHP+8OWv
+4+eWnxgSGqMb/22bcAw8NkC/XDqxC5ar4UzLxeCfIr/B/ODzHkMCSB6m54bHP+T
jLzJmwPkZys7JYKlExjDUt1vgEaZVwpwv1bv6WiyekqmET3FOy9eGX1ruziVf8lL
YeA5/3E7SkHVe2zPI3pGRW5K47CRPgaUIcmRi6czNAVDLV7M9A1r0cyznsb+1Mrr
UtqjS5II1N8LXz3r9MD37KCciA5SesEE+tAxAf0WoNmBP4gN10O180k/3fR0a9XA
bZ4UtawKtExZhsFn27+rpjTUwutqsllntIHvyhxzIJCsFxoQaH+QBbgh8H57dGua
5KmsVWLfbsP3vZfEo7bTV0jFjGje2iiDiWNd6zWdn/bEHodMXfUXiY8OlCWYZwhC
R0X3yOyopiX2ZP4UAc9lri+N+Uiv8Mb2YDiitAc9sqiapWnfpIhQifueHZt0I+VI
uRBkJWLCwsRxVafZeg8iVAVJuSQa8Kbh4TDqC9X5HOP8R/6A8hkXPw+zlyBK9IqH
A2N7yuht2FdoM6zKrW7cLDIOBAMFYGj445ni3jAZxnHzirFJnM4GhYzwXaywA0qM
k7lDuMB2lDwJoOA/w4CLZfi391w87hsUy6jY7eqTWlFSqbfgpB6xJfye3ze8eBhw
UVIB3VZ6dZ8goDNnpgmTdHtBXqGlRaL+AnpAYOXsrHRPyIKRTgkLdE9aPLMAgQAM
8rHvRhumKGk9Bp+jS2RggxLFoKifNrUikVMhST+md+Vq+wPvYeKTP0/zB1211e1H
fqe9CRhZhfHdGH1YFS25FwUdbGZNl2c4yzfnF3He8qS6CQnbwEZ0naEEaumzq2C2
pIvChlwCf30T8kKwTEfnFfz7QNMgCK+o4gkJvC8/toHvhn8ePHGzRYbGZlXvxF9u
c4Vo5M3fD+FrdF9oR7Nj8sv5X44c+SiMLwiKx3hio5HLpTBdzFrxA/PT4zMOlqvS
cIZ4OQ8NwqVT2Km/gCQcF9mPXDzW/e1koMqMe9/+0vZXh6RP4uEMI8rMuAnotCPl
o/e71uJl3AfutfjsoL80jRLVeUIlIEIkVPFhOZpBMJ6HVOBzM7qonfZ2N6UlRiPE
KjI4nGHXCztVlgMHHB5q1nue2b2Pmiw+ab659uxCnEgUkvkn+kmFFFVxWKlhUwkW
FhKtNpg6CaGMbMjfB2Yo+8jKcJc1E3+NwCC3QItmGFM4SzLspkpyQrponfGfsl6C
X9D6IKUpJ1Cg+ZkyAdVofiEVQovjqHE5L6DjYVD35lLlpDrAYZbQGE759xdm/0BD
g56aT8fLFLE93CtGH/w39cx+X17bKheT6WvdHVnEyvWKpodJ1eGcvcarWB1ZPJDG
nYIhPpATFK7H2ajsYw+nuy6ExiouhKK6aMiWdQbeu40z7l69azCJ6sLIngNnlXFy
z0mnFd5mJYEetIt7BJHWNk97XuQoCUeao/O0HtPxXrQNrmwnWekWzzV5hwh6y81y
dSXMCgXdJ5xEfacoMMUjJi492KmZmxcJjycOXX2nNFzVQffg5M7kqEWXst3jQ1f8
zNbYPM6wVhcxWEpOgbA04N216JRxuarSH4NgdAwDU9LHjitMXKx/kBrOyGDpa3qU
0lvVURkBppCZqtOgq6i7C0YllS6sZLgt1AccPHAv11GWy3bQaUahBQgxec0m1SsJ
osh36+fTofV1tdeYSvxDFbacDWwzJduioRyb3/4tGuTVSNF77CEdFFw8N5+1KvEl
9hj7b7CJz324wrZtl1PTvQXOUF0mrmXZryWrUo7tzLxHMvL9Wv+LenxD2vEe5V2C
8Fncjwh+nyAXzqSxjJ6U+hWhuPA/593iVsbIpEYgxfPVlFTp4QzuWxw0ZehHCLSN
eEWCUSP9+PMm6L9betU86Uemj22muXTAZhGVgSHoAUXzAJbUQzDHYwGIkBkRfSaU
D/gkSqxCNrzVWoaOv474koXtSmJf9XyhPA6HDVQivj9lUTMLjRNUor1WvkN/O6p2
TncpygWPFFdPAQSTpYHqwjubkVqFuR39yLpvuUIDAuvUTYZL+/UEuwZ+ljAQ/j5u
yIXJNhqnqYsK+EJHz3LLngI9eO+JSZWkBybCvK/YeDps8zXLdlHndENiVSght7W/
UiQF0yP323/GccC6dpcliSU8ImkRPR6l3m0noVP7o1Ligeifb3/zjWZH6TGEcjEm
DU8tGik+Ky6Ig1cvbWrbrck0GyTfwOH/TwNWFDEx8tcnBKXGxkjIyj8nYPAC22kG
dfAoFXwsIgx6M3CgLaX9cxcRxPvEEyCXj84VJrBzfCS1KD7aGkrloLGZsg0Iw5bI
DmvORdKCP3S7UcsrMG4/VqQSpldep9rivktY9wK9HI6vfimFWot/idlqXfWCKxpQ
e5cLfNYHXNWQ6Ca+nCpt6O0TzIMWURZ4SzYzO05xZ7GrGQWW0SASMT6b1of649Dn
+RfJUMW5CekTuMFyWM6wMjnAHQbXgaWsA/l/DD2TlMbSBTiodUMuJ6iLrZh+XmPI
AjixleIX5/jqhuprsnatczHjKT18pxWZsbqQQDUkqQUTdrRrFawKSK+6cSTyfRjh
PEXWzAC0w4YWvnu6V7nLPH9cdU/Ud5ithu8q5+ERMODZhsoKhK1KXLw1VRhU2xGr
WVBPQAmevTHk7OcwEz5rfDCQmbwsdud/4RREVAvpcNFRrwHun3po8wbp1mehzd1K
K/nyDfk0U0e8fQzQiH7f13qI/Pq4bjt52Ve7XGvcgRfq8ppX5QSuRCJvnfoXyd1E
WRFiH+ODSORegQVqv0kXQtdPQr6njLKF9JhIeTPfPTzI6GtCiLGhntBrA2GIw+nU
eDXA31ojlMsosYqWY5qj0wqMgnOHTono4bvxH8wIn2o/BKAnR29b266yJyR6yT22
C6/1zPhe6vCBeXr9237jHS8gfcrr9K25Jft8VjzzsnK2EZBrk0WuayZCC3RFVEVK
ZMMXOozUobTpHHkx/2O+iZUoPSwoSNKKYpZ+3t2ueAx3KGgQRY4nrx6PRwBsr9kr
AsuJPUXljLURNRl1G4T+hb5Xzjs/styjOkKpNBV5FsO2mXunwoIAutQgOXVZ7ZBb
0FsbZye34KEYzr1u9FniZPJFdzjW6nJWe7hw+Ar/G4R4lFVTrHubAOKGZgRLZ9az
nIDCL9yUy70sPG7nYEv6LCgq46CgXrV6DmX3GiSPhmhPs/JAbEiMsDyUwbUX9dg4
xCMpWJVecUmATSEJnPKz2xPR5TuV++qJVp19zF+srcXX9RdXaVRqY7r6WxQF08rV
N7IYkz78dWURmbekZG6FXg0TCclh6/btEGZe/UNTAref0p2FaUPI+rOL/IOIJCsn
wvtiAI8sPkvoz6zi01rLCoNiw2GRCtwFjsS2BU78y7zlukz2YKVCnRFIl3RUbOuE
veJxVMfuUT2az55XQiWamsFR2IPag3KAglg0XzGft8b5HqQR7Qy2wxOmPxEs55Ey
71nJnFBehO5iZsBJJYhPCPvfxgaoP7eXcJmT/GqsOjtRNUzlbrYdA0GkZknyDZRH
6lYMt1xQ9Bf0wceWnF8hjMrWgHNtqQXvS8fojxAWuXD8qE1kme/kpseAfx7Nvzdr
I7HHPHQ8Qz9fmG4ssmsLubL3qrXtClbWlG3ukJQ2lmkjMWqMbbOtEpshAodDED2W
ZXTMfQhy8DNbm+8eDbSVSgfwCYxSh0kiylIgEy+wurxeXsw/URHam49KFStHtJlJ
yH34U6QrkePrYgmO1fgWGvSCFVH9x2LmWEo30JDL9yXzX6i7AQgisOxoqFcnvdEd
mNYNkLnMJhzTVta6D2JT4FAiLU+OKErv6/MJGAIdavCcht0ScH7ginNOHCVHYQ2K
YqCMBeFyZPymLxw5eR4lSsQRLq4wMROVdlyApY7iTTpJqTJ+mcspGMJeV6fLTRcJ
q5s8DCGIQ/yW7ftnfMQLlctVFEEgygPCA5XpTkcbvEfkujToqKg2ikWSypFQ45ZX
rfWYoHSNTt9J8tfzLbfDNACAZkoZVeK7fB6rLfB/t7SMbDajIi17V5Fg8ccTEEJC
Rx8xF9PncvjPKJbyvrF6YVbj8SSnj4hUCWNYIW87+tOHi6vJ8+kKnOt5aXmPDOwL
W8UNYcNKUe532QQt0RmWvwk27uGgmi4mqmfsWtTDLlr4Vn8OooYDj9t9Jpt4MmL8
BEB3sSKZ+2JdhvXxRfshEUhsnQsVE0aFxwYkp40pCzBEmBsXUOwvdQx/0V3tFCE4
xrfiT+P8tC/QKjokWmrwzUf7asHDX8P1gKBbjtHJFZuFcJVOOk9wRXOk44ou8xuf
1v0YtbEsUmV01rLSFiIfL529yfQYPDz2vV/2XyL4edKQn3LXeeyWgweSUQAceWP7
fjtziOJhmkQPOlO7OqJI6SaLECDM1wUiKdYH0fqCyz/vjpC1u54zemYxWW+QdS4D
+Cr0sE0pEtCnNcWjuOl3l5Btgi/38+AHbCzwid8ILM9d3WavFbwoymthUGfeIlTK
ZcBQMTS3lRuGBT0CeLXLHOeNo/doYYv99LsCFnZpwy5vw70vzMSiNWwPB8/Jfv9t
796v04hn5mEi2udT07+7ABOb1Pcq7WivW24E/+6kQ+0SA2pGt/BRBySSjFJsIeiw
0QYfcmf0RYelv2zrokMJh1Ox3DLvWDKyxt+wQVb/wnjxeZiJqFIcPbfuvna7xGe9
hKr6Bq071KVH06isPSLILjbdqcYKfiNJm6yPrWpDLwzyhWD0194dMgNgjWk5q9Hy
UdIx5AoAZQfCTBqtoiYovo5C4fFUYq07dfF8BXeExdZ3zRcoAJVLheEQ8PafModS
aTuxM39wmMVP8KTMQxIF0s/o1clmhFB4AnOCXHro4nB42RVJmUqM5I2JC1A8txge
Ws1TihUmpnS0IZlNDD+FpazSzmEM5YLeYM1dJtbXXghMwqmyyJaBtQlWFmxqWcSO
uf7j+fw76ldcbHLp+Dw9M7ccnquLIpgGyLVUvJb8YU64UzZCn994xp+hc9J+S4zV
PMwDeTbrE8K+Fbh6Wx+R8PRRoa9GkhjVB3stPmaehibWpMAA2jMRpVAYbpZAV0vg
1sUQjlD6GkXNGEVVkht1Ao3yTxSy0p3qF3RcdZQJd/hCTj/OFy/S/U5org462NUY
uE8f38d9KRLsEVTci42OZ1+4hlFYrcEW6hbrbELjozq/eubJO1hCStGovKE0lzGF
TKxkpq5H9R8OlU1BI3CApWKHO9MZQJ3by2xifg/jUedQpoA8H+tYCnIkLVYkUHAi
jqi7HDdmIpBPPpJN0kxvQ9WI158rE2ZCymqir37yBo1tDBsQEvbSakhUEPwAJSro
w5iqgWYAq0PrHSqSq24xq+TiMloNf/WL1TOhrH2FLw49yCwHSy3U4SMblJfvjt9b
G3C9KX8rK/9q5WSW+Nk7hldueF9DoB0aZOsN3JJsYP1tTxjAzrW+MDgE56LDWosQ
egHebTpEEzs4grEyzlLL1Lr1yHQaYc7YxHDqXm3Th4FavCTiz4ApoKiyi87BKS8W
eT2JGcOAomGAcVKKWweJNhvEAb0bQC3H+OfR2Uc/dLv8PbqOVhENiTo65j44skLN
qU23cfgvhjJ8jZYnnC8Iao5YSCYpbDsb+KQUU2CuiD/w983ccFKAg8rwUWTkbIS+
cq03YShk5/pbwrAlqOCzLgPX/zEeIeueqnRT93JB/o6tPn6vWMV+kIFYvXLaVVqJ
wi5cz2nqCeETE/pwuUc9sfE7Pp3jAOWeYkbsDpGKCSeipKQAD5B/KmtVqw25ldkZ
eoD2rYK3XQWg4tMKCVYPOQ7rWO2ovZ05jkW8zEw+1AAPAHZOd71XekVaIcHGyOrS
gKAfV+iH3fJB6y+cM30DyDg/g2+w7OnxEtuMZTKbif7UfPjchldbC0fnyuMRKzBw
M2iFaHn1ai8F++4SdtTAhRmZCEI2exWwVluXwPXvQeRX+wvb87DRjhU8haI5f+WG
gkFGktTu0jaX4K5fl+iGhvne9hnpLWdqIrogVDRZvhxyDZo0Epi4+vDZgE6YKyVC
6BDedt4vI7WBTJQtkSvLJtG/gKyKKPT+Nazy/WklXNx+knCkbUTtlQmpsZTf2kXO
7qknGtg8Gz4YbidxpYKFm7/IpYw4nOsP8OH0N+UmgeWFFr4jZo/ANADjrlIv3Z+Y
zoql4sgm35s0KbR8q8pUVNfPEOrW0RKWcS27CDfnjZbxOCZY4eNsYgwb8TJZ5oES
1daGxLJFIBc0UTOdfdAWxVUd8BsMCoGHZAvNFxZ+kpTXPe0s3B2yctGGI01202ti
/getkWEba1IZpk26Ru9S8Qr85XLvroT8ptQgZgdTUtkN+xaWrPNBHU6c7hrn9iSM
yWZekChuP40fN4adZiWtc9Nbwh70nrbAuTucEIsa/5STZtXPluhRZq3ZKqZt4IdI
65LAZ1+v8eplfl9Ezg+fcenWoGvMKv9S9gV89A5UouKpwF0+0PLgJk2e9iu/OuAh
clTn/JYYR4AeCmuwMMEtSIBJ48SWW4mlE6tq8iPU37o7DVoIK7AhGyHyN0PKfYSU
idtFpOjaWIyuNdwlYx5/L3emyK5O9fGQvaqd+t2ehxyD4TkrfINorY8y2fqj5y25
au246otPntH9MrDdzmMGqLydC5HKSptucVU3Kz7BfW8EAIZh6/zKCQ9ihqvFxaJP
z2NaVKG8S6fLRQdY46tShyKMOHkWaU1xnjY0fp+tn3jNgGHA8oSVwpadGFkEcEsY
GogUAzy8S+/PbdnvcY6K7zkKviIgsKbH5i7pif9xykCwX9PVt3J1wyqevkxufWqg
E7mwTurxdwZqTbTTXTxSr0KBLJ6GuDnQjGPNXo/Nt0t2L69rBE2Y+CxRuhTZjURK
hNTIYmuJuD+dWl62cEimJkFyZ/4eH32PISZqJuK5gj4WksRGOMQY4VkJpgl49R78
slp1tavW+zATdWv4kqTC6P6mPoePGVtalddy9/yTd1ADDDVp8MWECNkA1Njh/kQ1
KsthPM6zXF0PIwC/2wY9cubuvlO9KXr5BjyHrvq21Vtd5qbFzJiSgweZX5b0PQcJ
589H+isj6LWGojOCdQnjgyPfQr2lPGH7Rf+t/PR1tvvIo1V3In7onh+/rDhA+riY
RIf6LmnDuc0rpY1TXdW33KlnpiF5knuutSDYMEeaFuS28E+QnAtAEAe9pmYGNPfH
eJOAlnjBuV+suCCpPiGIpbHz2kVdqKPMkzPS+qm+q86RA3unUBv9Bcs7Alsq2fn5
2zlS9wUU2By1XcbheJAiUOec/xo5DXdBrX/Id+a6dD+7aAyyJ8qccc2mzvznbzPa
2s19YpFVhX08XU3bZezqp6fqRqAAUNapT5pv6h6LqVdlhybJj2LEbjy9IjHY4YXw
wnxsBKaCTG7VABIFcStyW8erOi4kBtntaXrLO52naVU0GkeJpiramTBdwNZ6Y152
eSecXJcDMWHq4NrQDktTErkJfVYjH6ENPyHZn+dkwQTAkl9AoqA1QEnyp7wJBK56
hjIVFklG27igKjOpSUrvxthfRDJf7jLnXCIWazBtTeCcLlKRkezj2zbKmoybQ/IL
E12aRH67eYkPFtmQlLrz2gL+rhuEW4acPKV5htNt7kELQV4YGq73VraNuBbwZNuL
NXX5wmLrjDOORAt+WbW/l8/5OuPp4LXRuhMV9Bk30LdbfZACbp9mRLYgljpOr106
VbzGICRQc0zhALO2lUOicifr4dcO1I5zON2uHa9RYOXiGPbNuUsDELShUXtzK1ur
h+SjGBSmP4zMtpkFWgXfNE7s1vBmu/p3YLT68LHfkJCK8Q7yvDG4wKJKn2OVg+Ab
Xi16fkYkYyoy9Pc6748Y1GPCLqN+UfdzBU/GE9tpli7Ro0RolcrpgJAIsgi39hQA
MtJs8cOwfmP5yYDBoMisQCkqgVXecekiVnuDDCY7/dLHct7N3APx7uZ0nEG8uFbl
9IhXGT8thwtvC1ZCI19IVxHFbVL/akHxYcou5tuDyBfJ3nHOhGA3pBTeQ5kjlgf0
/gJrq/l3zhCJUAaBOqf8Mw2RopK5IhvW7TNstEcUHxdWLMiH/n3oHz6iQ1kZOvxS
jKSm/bsYWWBkdnlCZdg5+PWHeOzangfzdvHEBCIpdElIi+HG4trABhoS4AADLmZY
zW6iyeaT4z+X7jzhFYHMwK0oXwe1nsdgfsPYveZlBaHRD0XNFGULwggBS1N2UOzG
3Ue6WFEil8HSpJRVjkBnVNL+eGQ9eqgvwifAp8rP0yU9vhJITd7FxpAcjqWutG49
+KGrjeOrUVTqjwneVp4rUWwUTFDDwJYTklX+Xxid1ZLDMNr6XQbtdRW9qhjABP/J
qXZPigCViuS41dSg6Hy6IhCCK2176MMrMbT2Sm1pIKKS0+2UX1jNzw76KCq9MO7Z
HkGH32qKdre76w/ktD5ats/8CmLNm9fqsKhZ0Sj6kBYc8iTEg4G0+w5gwH/tnjat
WbUnuyv5Z7ZcxO9H8lIJ711pqQJIOP+b+79Penag8gcXxsBf2rPtDWdfs0Cc38XH
ssDtTgzOQ43pCrFRT2nZ+JqYi79CNhx/VdiAZNpM4g7KciYORmmJr6J73m+KarcW
My8NZnxFdCnkH0pH0FotoFVX2jpsisTwBF3iywBgxcm08KJSBrCFn3lOgsFB6Nwb
MKPiLiEwKXu/zwQAsaFf0a+cVzCgD+cddfsgFkSBergX/bXb9t5V2+3A6h5YitB4
cPimNowTFDfFwWllZDoyQcS1Gx5u87Fc6gpJ7KPtVonJF25cAzvMCWerXYMh1Q+V
qLcuZQDXjh2Sf5BFlVIGWKjfPttK930U1nqDToyDXYUr+/fEL8cBEjhkxak8rVtE
fZldI3/NK89rxjQdRl5TfsOprCoIqY3oTpxnrFlMqUvy1k5DfLhJNq61tylFG0OK
gmyjxxRr9Gw0P3Xf7K0pHJQ72eGXCLH/atjXxEaDZoF5Qrml68Z34Io5w+e033vf
c65NF7fXjZsEOaaO4Zs40GMZbgCFqVJJwXKEjDRDO6VVL8OPP4Du/7lgmrZwh18+
jiFwLuuNzUMm5yfDhUs25uM18s0ZinDjIOLxT30sWQyN6CitpgwgPrBvhHNXxQKM
txa0Eq7eBc4cUO0JzimtInNy4Rl3QsM26WUR51perphm9AgTsYJbXzKZl3xA18l9
Kb4JVFX0U7xM2QjQo6OI1wRHIkqXRFshAlqresU4D9AsBcWOsIb0ZwRh9oL/lDSH
4/Rpfx/ChdT2TtAyzwnciJtXqLOeuk3/65Y3Q4DhdOMFYNYd9BMi6dg0M96w6Ikp
2Iw3QH9GZ/LEKez8/md0Fo8A68+DPzy4DnJA1hEnN9HCZ6y1+DKrA4H9hXfKIqsW
ZprCm+BEZ2omMKWxZ0RgbqDDhsGvItttBLaMMTrkDzOIqiUFn+z3xlz+mGoPTphm
hlWmDX575CzvRrSYaNhABG0qwkYX+EWk8D5DjY5cKEFTvIr80nZD8OZLE9XMZR3N
o5PRpJ4sbhWLcA2MKBpRKdG1D7efGs8KeTndjjmPZa71dUDSdis/S2Lh/72mW+Hg
Jp8+BCM+XL1cp0DRKKJ3Jj1k96v4ALjLmb16eb/Q85FbujkVjF77sHMQrodVdrV2
p1l0/7JTKs2S1EjAUMCmguUbwh1jJbn5tgPBnQMoKuR6NN7q1hP6GlFrNYtY8Dyz
3AqzAf+oJGf4pDHSa3sk69cPDGg8IaNkul1DBKPjiy7b+Bt/Iyg7tBl5GHfGWpQT
Jje7J9dSRvPbkc9Kd3shw1rBRVhR6XuckitlCHU2HfvysE5oXFYGuzWO0avcnsxd
oejvC55Vo7Jgjo6cDAYqapVsO6AufWowW+ILkCyt2qB743Gez5IXphOGrI/sXNin
izGJwTLi1Qa7OeY2RoVmUda6HrfFkoWqwWGONMOMHRRLj5V7GdbJ80NUlLHiDoI+
4TqbtgHZTamrXK0NEXauKw2VDsAxYQ1a6rmUEaTdvNRowjDSteMvwKyTkF3iRNFF
4klnuMIaKFFNnpdzA66GzTNZsY5a6oMBSpMpl2LJfTFigUeOXjUZvBPX3VYVr9ZS
CsY88g+6CsDrhppU8ltEo1V/rAPJoTlyusl4I+1IJj9IOxKCeCGU65kxgUv6N1Yc
oYYW7R/nhGnkjCjhAWbSh6cWelKQMUfHyS++63YgonK+tvwTlKDMvj2Wf2JECjBc
Awk9fA0auxmqQhBzCsPODlaNP6hjoJsiABRbZFusuT34qpWm6/HiHR4fbv9il3wM
iOZkNrPSHIzRLud3x45q5Y2shEHeU9nkX/dPgp6RogKXoSFjSgmu+zINBfSHX1FL
9vyimcgCHTf2BCz8+wQPiHSBYCGCY5gxlrtLvYuOiCWR/ygdggZmp3nRbb2Fiifz
ndANwQuV55qZ9h+pNvTfIgFqvILYQzIhhCwuXyODoIv6Uck08Pol8kFqCttGxBw3
4sSrBkVkB/kq1o6lT1ZGO1H7FwWnUjjZORymWsvPTSlKFyy7rFQ09jCAzEzIu8ge
guC69CZ4g6GZmmQey4JOtnbggr6lIKWuFQLue6LFfXZgiMM9cGa/5CB9YuonATqM
MApxSsSMpjT8H/76QFBk5AssUO3omudQPP6UhSsRiZfpJzy4bRq0lJ2Jc+0BRLXc
FEo9On1enyGL9xfPkKajgqAu5W3eFbcRq+ntYIfe2a3QgfgwOINqk1eMQHUtATlw
OoM2lvkyuYELxYrgYneBPqekMW05BLAEksgTiE06qBvb2oVCN+WUPjnsI8FoG7r/
1fftVkvPp5MFexaHNMcGZtmXEjwnHRWqX1b2BDVLmxrB9pyaiWEL4X/foehxOqN7
A3TtX/nNRLHzDUqaeDQc18BQGMU5ahmx89CKRf1WUiiWruMq4mMSK2WYYeWPIaHk
S80+4jqKp+ypttSn6PWhE9Bk3m3PU9GPgWNWth9OjxfbtswcPRisHAHILA/4zF0i
ji4+gN+syz3CcPM4p+XFeEnEutph5PORiVDBaMBl31Qnd7h14m4d5IayowhmhEkP
eGqHUN7VhmTUGzYNdyFVJH/+KpYAaWdS2a/fPECF98tBNqMgQz32Na0Xwjb9LpG3
FK7LRZImt3odVb/aSbCylo4j7f363ESt8RqQ1GN0lr2D8/Pe1HFcLEPR53OLsGBQ
7zbBtSPin4JkbOt7K8qI9c1uaCfJqZ0UzqXQrjZSrNoblB6MNnZ+WN+2FwTHXh1D
Gw+vvYbbMJb/F8LpPgDUJh3rjVhOVlReOLyjSClz3kCykWgMDsRtyyyADUvPciTd
8Ndlo8VxGskVzYpRzGJgRFfZrIsUlsloVE4P4MLf3nqWJOes7agq+QB5uZbLyxgd
+ltDok2tqF01JaxmH86UQ+jeknKCXcyh7J1OG1YVi76Yct9Z+V7a+j21yX0gRrc/
oEZErBxrb0/YeuTGUahHaDFhFuUUjtg/Fj7IZFC3nR8ugeuLbQ7u7wkDfOK+B7oM
9cPz44isG3xbPL51uajJRM++q4lwgwrRFp1jTa5KP9wigHSCk/iIhzEMys3HZ9to
e0wuf543pxN/3SNnllDdeND5HhnZybGClT6hJD+sN/XDTA13vtIneCynGBHiC3+h
zpcBsv14JsNyLd124jgNIS6JPmcLYf18MY5g3ozNzqlMzBhluAqLdBa5L4eU64jh
ZeqGdLTEm1zt6DJI8blE261wGcEe9Wz2/5j+jd+qEW6wxqk/vM3+i0RT3FX89vjl
IEy9tI4Syjj4kmHWIn3A6ONq8O01usbTwVDFg11LjEl0htVLFtkK6EROOsphkIeB
sDWTZKNU16QUd/RvB/MyvW9P83a1jm6XmNlGoXA0J15g5LMLDltB9ImR1IyWnEbz
/ckBYffn5FJAn107b7dzE2WsBFgQ6ARCs9nliUae5+T+McFWEuYLg/zHCCLUslWI
Y7Oly+Cj0h0XVpOhf6+i5pLSkDyT6ME4SpNRBkwXDYYBxodhC99T4MsNK4GoKkW5
XfQso511GfzQdtxDN6U+doNVtsGErtP4a1hC8hKTHVJCZ8SpAS/71oYvnSJUB4Jq
vQaMfJx5JP5tCF+Zkea5SOMg7bJHkJC02UcUKrxkzCFAmS4WnJytSGq8zY5TDSKR
fZ8X7bkkjqZrnq175NwyUgn7BVFKbWI+G/qpvJJxQoh28FzMg96Ci2mm3nT1ildk
h8Jk3qlXhRwzDBhu51/IxdqGQDTayxx2hWL5bbP1v2sq34QPB4PifaCAajQfGT5g
HgP7zDvRjEy2UOOM/5jDxwthm1OHUPciyKZHuQHSp+FBzpvE5XV3yckmUyEmaGD9
SBhKjqJi7qb15LvRQjjinT8u/XuCmTfqt15PAQq3i2MKaq1+0MhKdo5p8fURwozG
KZJ6J0nTBRj4n5uMtGw9P/WEVhKM8JdWi+1PHncFFG1DBHmBWLE328Ga8BfNx0aw
/IEK+TwnyXWBYKUkpydr5hBaHKJAzIVH1/bWWshQM82fyQxlAYkuy5cddqVLoMBc
9mU/o8s3xRkXYumdrLICVihMDOmZnrJ1CMwd7LGikAVKf32a46AUfl/naVmtRc4Q
9kXFo8Pz1M+OFAZIQJIEWUfycHHX2cjK341cbGEuuDs7oUV48ClMBfU6zkAabpbU
VwWl2k9m/bRAeElMF/hSWHTL0i6JSppCqLc8H4jhhB2B6YzjZmyM6xLMUlkYGKCy
teFwA+NpsujC1OzGuAHt0UOTIHQJ079GJue6cqQCTZAaX3bhFrjtP/Ek0EEE7LCd
U1lLdv/KyiwDfczHm7EtSAawgB69tAucWd+JEjkz3+4AkRq2rYYSvyLRl3e6M+GV
9Fd1bwFiCUrLbY31zq3rDOvmV5I7Laq0UTkcL21iu5+Lfw5U1pUqOd68rfSEJLOV
6nRxncIgViEH46qvMq0pYYXcvObVSyP1tcUgpabMXiQLyKfz9wW8aRjKVRUS3RO7
QhJBYMvty0vtqQwuMegWJi5TPBVkpfF3RZ1wyqSBZZ7uIFu5GkO59j5pJdpwDzC5
sqp28qQtpfjrd7jQf4Cn13DHrzyC/SsFbJk5tZFhWjGwTLRARzW9hH1NLR+sdphn
Sh5ASZ2ZkcK1j3j9br+IaqTluEyc4+ybJo8KimsY3gcyjf9neCKLJV5suPWzyQxN
Abo0R7Xoi3HpNMgjPKJceocDKUteUiadrTAsq+5Gm4vXU5wm2ebJ58Vldfp7i4KK
p9lEVedyVQmOUBT+Njx53OgRAXq4Qi6z+guupHOe0f/D40jm2eRMfMnwpyTCgn6x
dvtnG08qhuYfdrJQGfXLxDNatdamV1SnMhfcNPvLq1GZJzK3o74BNAUibK0UN0dR
C1tD6bCsIFTpr6lri5HWYhZ0Adi41g9z4cOq5PpB/NQuVMr1J5Gd4fH5u4cvZBjD
nrcnzFFTEa11ElBW49jfGPrlSDyli6H1r8vjaxrzwG2tmgfDksB1XMMcUgXdPGum
K1KFxoHM2MHdM1q9j9sz9OlBMtXdJVkpkqXUMddD1MiRThayC9y85UlfDDUvg+fm
mnkMQC2nqXxvsFWc1hFgJ/8HZo4yBGQ0JLglotaIxJe8Huh1o9V3RGjlxTqEOhJL
ZKrrFO9wAn66XVTmWcqpDtMsGp8YcrKOQTwveXBwevja6FWUacRjX0dEuPtr+tJA
/sTrpgSxeAsNotVzMLoNvR71VxBwa25fUMBKRXIZL2lqcvIZuKZuHG8cms29fb3I
v9dW1iB3vasppppY0cL8ufBCqXYyyMN7T4oTb122czz7N51TLzFo79U/e/j14sJv
7CmKxrxiwuDEbHn3pkwInwnY0CDoJIwFXt1F82Zx4Qq7Cicjwn0ZZ7mdXtaGuko0
s6aoVGMLXLLEJkL33JjCgjzcpQJJ4dhds0N/+8QfoUu76CVQRJeSvayW2CeRlYmZ
Iyu0TC6PGAz6GTD6wYMYBAETeTwXpMDPzR6qhTXGNXQp99dClWj4DQzo+N4AwCTR
fw7UtHjkCzQCZbtXnSz//ctaPUo8uZyfO0LrVWitnx9P/1ddeiqigqLbCZhTCMwN
f1kZ+o0s9qS5xeE5p4qboNuL/XaQVNjpi1lXhBw3N0ibpEQ92/aoo6+EvLlGIx/q
hfIAWfK58Ubk2WnEwJSTI9PfIR5/qyOjx0LYMUUji52eQiL/ldKFb+ceudhHtbdg
J/RUkGiLvGwUL0yBOvj9RinnhtZAYGtx1bhnigVk0C4mjtNwDsNkrIRnXcjZ+j2Q
Bg4EcnXvOYNMkAU059P9F3FZ6r7k9z5k82lLKdS9K8WooYhCYvs+HCzq1YZokwc3
ZfSammWH96fUSVnxB7TuJBiuM9lrfF8YrYGvJnEe/7IlkJ7MZ4r9JwDQhAKXz/V0
ziZBd2ngTMHZODlq65rQc62kzM+bYYe0JsXTLFgDFha27MJCqTX5sBWWYqM1H6Y1
RxlwzDkIK4V0Ppcl6SzlIMPl9r522G6blc3Mna30600RKcrS/X5k4xsJsBkEiiqR
oPUzvRrHD2BpUhiCNzq7/EKLNAbELwj2X08du+IngIKeyJUBvuMC7ClADjN3BcR5
gJlzRylT9EE2u7DznCtv5ddRJN7Ub2tkdgLSNtF12Gxuv5eNfQJkUQ7U+67ZoBCV
b3kDi0NDHTkupNsHlJwrszK/kwD4ojpIZ6QFSbRka9N4X/hb5HRqrnOsA0FwQvGa
C2f2TugKTcrX2r/PEly5NQStmXvN4pwHEkUQP7t3nvIgEkRxG/KAkavRWUj7NniV
zrnTTN783FuR2rKF2nKCmNNMz4YU7Bo57rB/JIcxMc3wCrbZs5CIh9A56wWTLln2
2yfBeAe7SQbTqszBGksc7E3dbgd76HF6YT1+fpeQR3zeaarBukeiNE3wH6TOBQbZ
HVtJY3uLMkLu2+eIRJDNHe+lj9S5xynjy2VhqZUx7NyEGUxdbutn4tnxsAuq0EdN
bmNNyZbYGWZRMKAlRlqtwO/9hpJ3EzKrfzCI3OvYUPHroGXOpGRSRmBgS+pB7tYE
fOxm6SsHw1qRacyIx2J6S9DS9PGK1NTfGSNqM+66kUf+hmhPWq6J02jdrYyWoiUt
k4wm8apDZgtPLdBAffPVg9E599bKe56PKsnxsrLZfoTercVI7KKANz32K1aU//2F
UOgc/zjJCzLIiqXvP2m/rNk+Ux7fNDfG3c662NcPhydmduPu39I4LwwdClDd6kl4
0tu6EisFUKDW2OxaHQhjr3XOhFSA+hJRXhm1UEoN3A4EDysWGpVNMkOCRh6vzIn+
pazmQQ8GdaKVwpEaBtOyto1PMZZ2YpMiV3VoCjdygsLR6nBGIlHNclRfJQv4e0Cf
77W/1krnccg8Giv7+Op40xbPIHuv7Ai7e01X0c3yEx3vEKi1N487tJhCwnzf8373
wlNWvHMIHxyUGbH1PF6sKPZKo+zP4lI+lOLmOvuE5MpZT/ZXVNOd17PkgnrUcaDq
stW/xVKY0gdtXeuk+ZaC6A+vKQbUfGXp+5QROFuplxUx7L0mFTtXsRX5HryaOw/D
yZg0YLRvd7YdMkyxA7Eqn8z1icKaemNLSRYCvbP+t0SfKhc42QBq17rWrvrNTGEV
pjCPVKdmKhDzNUevqYIZrWjaaQCg0cWWNg2HQlOcwSglInKAoUz/gi8EGPlTPwI1
sr0oeSfbygPalM7HyKlI/RSsUuy+wLYPuEP82f5lobZWaIIQlv4X2C42QNaWNJAq
yrqCkFFavqJeQvWl74/e49gjwDpWo9kx3ZWYEdxFymL98c+n9MPipbqHu2Kr5s2N
sqvy+oei3tx9BWURjsRWfxBcA7snAVytDQjjAvEXW+LBp5YyG4bZyj5FCFMLNXms
aO5nCmvFxMrnT3et2PX0LbIk+F7MM2hgBeOQb/ryfirEY101VgA6UoFH8BR6k1iU
ERoigXTY9PqzgNtBwTZfluuTy6Ssjc5CQO39AiF0pfMCUJSlmry7dfIDh/qfW+QC
u75NR9oFuzYlAOG8XpOyMVbVfXpnSTaruZTyFVVdPI5qvq0SGs9ANQMNPXE5Hnox
CorpRHsbImiqWzOz4CSdOipdaF0aU90lXJqcwuJKKL4KD7a+GBEG2slquvhdeDWF
jw9rWXzzjbNvN+5wNhtaAUpPf7c0DCvMUTG1/EjwG5T0LJV7fBqQ37BLHMc6LPmv
oWgJGd7we1PEqGIzTAB1Yxln6sI0f0IeLQoYcbERYXiykRB43KgxxHmrrvSQrWp1
eaSrJjdjfenYorsKlreyEXxfKQDItskTFu+oX1OCQeukx2W2E6zWe9p8rbohOHhq
WyPEcT8sP3xTUUoJMJSyKXivkYOXrpEMwrEDRBWGGn+FP8tepjjrgdFLn450bldE
5PaCKBEUa8/CH612TXiLgkJWY4NGcb6bXdXZg2db40hwOv6OD6b7lUsW/pprINZi
AMxDeRopfErih+UtZfwl8usAaFrfQfPlWzZiQGdQKN90LZjz58Kt8/7g+rxLJ2HH
xSSOLP4XauIbU8Tee/ItWVJR5O/M9syd9Ci/dHCLx/TRJXI71HqI5281gpV/uRvp
utJQtqy1vw3RUmKhm2Z72rxd6rTHpUbZgjT4s3sXJMNtQqUEk6gbXARYh5tFG5Pa
odT1DGzt7HCbzChZMU5EgjrzSHF2KRzKzaxPVEFSCdKn84tMaYyPcQdjnBN7l0pZ
ZYC9Xi023A+DVBMqwepXQPkJYDUHNzg5CTymMOXeFdqj3KryqEtdvJuWLA+8mpNN
e7ocMg4DdXBIi4mBIbrzQNMXsazThlDC9F6TqhVzKstuWd9cmbQYajHiWnE4oMO7
vsd0aspaL8OnmozVGaVkJ2pGMZVGd/DdYV8VpFAJfQ/d+S6Cre4dSVqkQuxbScY7
6ZFV6V6DzTYgKqZgO2YV4pb3lSHNis9kzuQZ5F/bpS2VC5aJrcsXd3hQFrCYeyPn
P5RyRCaOAYI4uGb+8BrfMU/YZjTzYhvbD+4BT/AROjBeNQyj1jt2N5stQQQqqYeI
6zXpAqHnRqRTceVTDcSuFFhsiXNDMDfCzngslmdqqDptFGK8HF84praBagdPmsWf
d1IV+5orR9KfN69Z5xrFz4sJvM7eMJZQeqXXydBBI9K8A7W5QKoNU/Aqrld9YSS+
0FMyPst8dq2ywNRWFONPdh8sUWUG2sLWvA/PS2S+E/cvLpfrI4vC0rthgMwL1AEl
kQOEXKUNdSoBKIV6PLeRNOESn1dY9ZetQls/brqwCw2qoRxyhHH3XrhBMxJgoVnd
dY8HvpAoFCiEzL1ZbJZ02ZHTYe/qNC7EK2wXpuv17rXeojRZCWU1c7LAEYCtTBLb
kJpNMLkCdDVoTiheHlBLT5PgdqHvQpGTOghVXIjzTToNcjfCaV+6NDLCw1yUgXAm
BhCKGiQVY6h/JtJBxNWoHfOF6TZXArBWzlKDlqO4z9UuIeuIOvQxKK2zgJyAmNJ+
y0xg8+clW5F1yg0FqqcmrMqqBRQ10gICjHCzyIFmUSq29HvgWrx0fz75cThxLcKa
L4YEomDyGNYL1L4PAM9BdbakbQQWu8oO2n47aSCS/AMeeffZ6im0bremyEpevwm8
apY6b+ncUDBtZ7nEBXXb2uI9wWyH6d6tB8FXc1jNEBANClRKZtBxdpXtK7sQRLqj
9n3heF3uhiVURZQ5lCJx+G0I4BqZoUPisbNaxQRFxJrRnwyWt3fmIz6wpftuZZ93
UVCjuSdG5wWK/h37F1t+mfwwpfab9EkZR4MnzKcc4PuQf5k17O5WgKi7g5VIEAyV
BXNhq73eIkm+tQiXy7PF7C+id9n/0yo+wes8z+qwOZMkee8EVoTCvULm5DRMdqYK
hFUYwnL3G7ZW8Uu0UOv4RcptHM68akXHFoNkQEpJ9mC0qh8FhPoioXoKNJRPBxbK
IR+JKJjgp+5HHNILQyLkMOm32gOE04aXr+lcvyd3+hmbnjt1kNwhQ6D4X17OCaUl
LdI1XCavwsta/LeiQzsUwCC1DMayK/AdQ6w6QiST+nJP8UaPk0eWSnD+kedaAwHT
jIeJ2XpmTOiKrPgoECzaWwL9uTD4160Uv+GdMkSjv0ubOZiY28xSaC4KY4sfYu/6
f1JgsNdkXzM5mTfYBvaqeC5BUE/9FRYKjNu9ohVPkZBLGd1PBy1ktclirTJUthsL
MZiEkBQoY1H/cO+BLjRXal0BIQyzWAGPDKNy2ALScsgfvQ2HqGg+xjYpPIdY45az
b/BgenN4CIV5yt89vo4pwyF0dF0UJ5PmaN8AdhkyCgMgtTH4SQ9XaG13OAte/suV
zQGNeUmdUzVWcxdDQP669R4wNZedL326NOP4h9SInMPmC0LTYafGepjEBE9mZcR2
QsreRqkiRkmIspGkAQqvoJ19MxEtJxMYVpDT5A9VVtS5yvArLwyPn9LgpiILvPax
fmYCmoWDXoWJcuyOrv2nuqhdOY7iXRNf3e7YYq3/kt9Z6buh1uHkdhBP+YUCxkBF
qlQg6N93K72KpKZgquZNn6z0Ex/YI8EC/mg9IbM07z3P+O/2iMiWPFcbeaJM5Y67
55ZqwBW6Kom5fl/MADzQEXKLgnrV8W7OVgfktNFGolf8WXqVfiq862UiXj9YyJQ/
h686NGBwb6+QsxUYiTD26TZOBRNwM+vxwr8j5wxhbeM2ePqmPtQEm4cYr1MdfC2c
utXwYklW/8Ss02inF6loMzjORQu0gyjzPuJ2RCtaY/fQdwoL+sJxswCUL9SzonMi
WgLpm4CE/ZVfHEog+ZRmN5153dcGKn6CSJ1PvZErPeksmZyDB3Cd5OoNK7Uzodgu
4LVEG9wIrgk6X2bs4gAtPgj/+ZYGjXRWdavdrKJlLt6x1Z5GxLIT/tizCFWQFpwp
yDSfcx2Wh8MDmkcC6eVB8wqLwXEaEbRgw+gjkSEMpG3I6AqJnKJkU8KI6/RpzxFz
Gd65/ujcLbA/bvnpNauMBvs+6sSz9xi7zvm7zdbURovzZtqUkdNgeE3/GvwUIfVF
uH3UAQI65zti+SMFma8ogswIuMfcEBV8w/xf2dQ6yEJfJ0123dNeo420e5JeKMNY
4Zb2GPWk1dUvw/xNBV6bxJWTrXJjnaHA40Rx83leMDkoWJ473SzI+Cso8hEHHJK8
6qoNFrN/5Dex6cIp5Um3tbg62GOpY1qbfRMz6HsLRi3RyChDeEXjUl7Yy09vjpnJ
LLI7VT1FXcA5EBLp68ITg0ZEyB/KybRSkETBbU+ZetX3cQyCgiqIz1DzEoOz/NOw
LqtQhskrVuo7IEkxrQq5sBr+z8KmA6/x9QmUbQkaDfbblvDILVC9GxLOGkPAo1jZ
hlet4cFcQWzzioOGnN+Jkj8fO2xK2knPN53s+cPUGA0SbVrr+6JmuJGtF9dwaqRg
p7fVE4v5gjCpyvidnZFjFEUmG45Ld4sIjWCShedT/L/DW/qNZSH9xeTLUE4FTuI6
8oV7Sry3sPAx14DUOfujUqK81yxTcvyoLcU8XpCwwbE6qozkAsmb+Y6a0PrvaloQ
a5opaZw7JSxWMDOjSDcV4PxJOR1N8b5W3AMXYvTur+px3Ol5Vj59IrAUJY3hR4Ay
GwvtCebosEaA1+9CMKFRQE9cO3rWCPJIq/vxTY20897AhjeuubnwTchCky8O3vuT
8ZH3jNyeyC1uI/hw/NZu7iEpd2VtPtC8wrbWP/JPjrDugAQQVYIhCPt4fD5Wd0VW
cS8DH70iB5IdBPpzW/n+3xcnYgH0DI++a+JjRRQkxD9U0FwSiJOjn+OHtrjyM3xR
+W32rffULULOdt1G3ll4WFoY+odq4/0LKk0xKpk66o5W4F1J+TKnSTmKg6tHytJz
nQriI/s1iiR4XtpWZQnyGoiicd7Jw0sDVkyJUtCK6/SvF0dVpIJ8ciWiHzSHqVf5
/v/W6RaoXNb5kSJNcBk5GwrmAkdxavy7Y6pE8K7Sk/8K3VR513Uq6vFD8tzP+UF9
Kiq1xrwc50mQKih+AOKBr0JPfBRJ1YDV7tOjBFr9bd2F2jqLHwjvjlnvFJM+FOy2
qTD0d7s4LUkKqJA+SwStfbvtDjPcvC2PD/m8xjgNNfwiHjvEEyjQlD6Zj1M2FltY
+6SWS4GyJ5JKpQkYeOGROpUhoyhM0fJ3PcR1TsHy7j/Z3zR4ae+jU7WYPoHmJRb+
/JmOGpawAv6O79QRmqT+9kT1EAIZt6sXCJLmQlUZU0n3xTilJQHQx0N+J7Wc3AUQ
TT69fhKzz0a2Z5bMu8a4YQTd1tI8fcL5ap1VQsuwZVN96A3NvuOlutrgLJrxMJnp
imA3UV09NqNa63cs/je0yg3MG+RBQula7J/5CQQUozPFfSaSK6dju2d7i9KVoQcc
/COQ8B+ObC5Kc84dR/fjsoRABzEtE8i7VU0eiEHOGSriHMeOzT9abxIFkA0Uglb9
AJhsr/QVJqCabKtdS03GyU+CelPuZeo6xN/svYolQWl/ZkiJebid76OIy57K0FN+
shD9Qp0kGB2qQmvyE56WMQyZi+5Oq1hP26++5SD2MYu7qR+dK4qAn3z0i8nB2qwX
A3WJmydmIYYueybOGVn8s+s1zBGyiSwsi05JcjAycnz9kgJAXs5yE2CT8QLqVdQ1
uq/BmUJ8SMWSmw/UQHYA+0Ph+o4cdccml1tFqOHPm/sQB5lM1EngBUAhKbWPg1MX
K8qTp9GeBZpNONmDqwVcqHkLyTu4Dc46/sJN4YdOL+RZUDLtM9Mv3PFZWrmHrdQy
A/Kf3h2L5xkz4ORNrDCwjOg5axOw4nPM1xoxwGGGrYae/rl3DfGxwZ6EToGD6k/M
Gs3h1fJhuzugZkKE48bU76rgytKaV1JYBU/CTRYuxZVV3xu0IMkms20yZ7UMFNhA
slSeWmIF0qL5Arqi/Rv+wpzH04eyxiWs5Psegz06ilOLrL64YLtEd8H98f4W5Fb/
Qa6Gazp0EQIQx4Z+BhHMO3QzIMrq7OP558UzVLDNQZTqR/ZYg3onZSor9a07htkv
eNBjt87nwjdEn6bPptpOLqpCelWArON0OVN/mUh5bYfmzyXhLjTKxFPc9ivHizB0
CKYoGohrG4liVEo+XdIs1KfgdPjKlF/3cfvypzObEWo8nRTiHZBaylLegaqDNxB4
CBcfFXy4xY+Mx9m/wLm8UmXcJqKgW3xrAomWEhhCsg43Szyb4ToVQNSE/uYnbzg0
hT1XVHSPKfmLWnf1JWA0r24lvmMGacwlwYP+O2m0qAU4weIcFZ2m6A9gzHnTeMMm
MEcFz5CwbZEpmkRdMtGXB+1/U1A1iORd/x+PRNUlICRhb1m2cRvEycitvYSAF/hd
ZZI4+OGBHDEwGDA03N9HjZHgc1T5hTK/j3RsVCVgCTki/J8mqweKmRhiUZ/J1iXf
msrAR/DnHcClH/A9vfx/TzZ2FdDzV1rCOSUwUlxmneOnNN9ukhYeO6khiPEjjDsf
TSEM1ealG4x8JYJslXfCFqxL3AKYuROurzl2xJiXkFPoCBTKXehSvaosaqQtM7M+
I3tJhwIgFxHgQgS/C9IORrzq6UsPCKwIKJrKyZwXlxx5kJP6qLC6u6/CdqVJOjUa
oYnd6h9OAt3+oi0tPadwN9G5WXgUAX7dslkLNhdTB9yHIxIbC2zqE8WTlsoPESlR
yLbERfWwatPxPz0brfiUaed0KMAn41i1jBQjbOb5CJG3BrBH+fXnjK/S+RWEMJT5
XvCFrSQ0160C4+medrrqkCySY5Q56x6i+Vu7kqMfS0tZHAWTT8Vwphp+h56sR/Z3
Ai9P34mI+op7dBrlyoc2Rrw3w1r7aWWLKkko4r47fV4tfu8WpCdjPXsOc/ZviOPG
+6Yi/dJhk7BpbgYgi8EXPFxQloeolYsDF2cVRdp1ukniUkuI/GslWgBZ7KWp2qWA
cei55RrpvhCEvXwcfw5xy6e+UZyzrc3XVxhaKRCFL4iqxnx6/tyuLXMnaiV2ioAo
TWxs70/oLymzqnJWY04qURZklHo0smgdNmP67J1lIp/TXwf4Y3mvv0vCsweDjaic
4OQEuitDpgoUaF1kMLiHmMhYaqNnJazagQ5jfNoz7sSk714B7oqkAKsKyOYeNM+s
amf9Omy+sgGQcgrM+KlsprNwo+dFdb1BQa/Tq5uwp7KoeOh/HRl8tk0qXvphU7Vo
ULUcrQMtgpvzUVfBidmqXP5vqMoTe4Hs4LxtXpvY8Y3nWGewGiIcFeid5s/Zf1fT
OQs/6+NcWCk3jD6N8gFAN6R2We40DCr7S2x/yJtSBb0xERdEStBn2a8+cit2O+6X
3OQu5fJSG6x43fARTItqC7Ry07ibA9C7NgfTtxTs0h6waDf+SnEMYe8/y8eclBJg
YVgqEqDIKSPdwC/5f8e3taFULFBqitg0EUuWiOEfCgyOW9ufeZDNFijryuxrC/G3
dr+afSP+akD6CmV3eywup5Octy/VRKrSBjLnaPeh6aXZKdPjtSDQmAbd5vE97jT4
qoSfYI60G0BuCM05i3qtiqSmVEInnA0IsvaOT2FY5lL5OcwZWW8LiNI1R5LIDll+
lx/NDsxyZW5G1AnCrmRSG/4X/X5fgHimWwXarBB6CAIXgJdtcnc12JzaFXsD0Vet
vXCRZCc/TcJkexzcmLsjCB57bwFRXy5KhodgA9AMTUCRipJ1ti+dMgTKieNa2ujw
M706JZbdCTlmMWQcKRIWJ9r8vwPrIdwpyrYIVUem6XrR5c3O6Z15uYEPAqZdAxeU
4ziiobNJxHtkqp2rFZyW9mJS3KJp3ixx5j3hHFwXAs5L+zRrKGE9se/l4Gc2qRyX
LrJpTiUL67yWYjSKLuZ3aYdTv2RXGRVShrSMrkJPdaQjl434za1aDuQmKT4oHu2m
5G3A5VkXxR3kqxd69t+FIQt41BrElNZN3ZW3qOgdLLcwEZDIW6wwxFKfdLG/EhXd
xORLVp52hoIonec/pOz6REEvIxuWppGbROfCtJPrGFITEpsKpkYQxF0ltvZloAOP
fVH/mSO2Ppbhz5S5c5YKFMNEy/LTUlYV2FOXCALAZrqoPIJIzzZ1CiytRdHiSPqf
8wd7XyADM8zBNPW3QVxfL2jj5qsPbrv+Ch0ePOTyvvGFVz1mBg09KVj+1uI05Cpe
Z0pwZhURMtlfv6+ilowh8bt5JJkIp0LElmFVXU9cv8aHUZwk9+gzGn3TnWdkLrXJ
iTq54Dn/tcQuvQ/TKAwYZ4iuDK13yd8NFTsMUxMaSTbBS0582X8OWKtcMpcYXwVS
IxDODtuxcbV2ze5z3KuUh/OkWa3nTIKDHp6HCwmj+/7KjYoNaUtLzg74QMPF9tuK
wsvjmYgRJnlr7ov+frZ/LmOgdh6Hj8J2sbBvJUbecxbOz3GP/1raKrgThEzlNNGx
BnsVOahhQXncxwvqLpIYk6RuMDgrEmDYnPBGSnBVblcmvDqmyo165tzPtbnFlVBT
vXcpM2eDgmmt5W86aphrB+G2X1aTZqteh9CdiYiH5YHjpWVxKjXcoawvs8Vt93wO
Ug+9CxvY2DHH1q2fKqF+T2698NyjcY1FZgU0BWz+9Y3WeyV4aAo2HDkt8skJeB0r
YXZAs204zyXloy+bvBOkV8GoC0ZemTdvjgemzWbB5ktnsfyGndFk00HUKNzYLlMW
35rOz2lUtR7Dfc0cRPQYmNUroVOZc5zGYNkDJHN3F/j1AH+c1OtY7rbsI5CGzaGm
5eyUPAWm2jM1dPcsJbdBBSbnU/tzjwOChocfbHN5XrtBt6hH+SWh5zCieJsDJ/9+
zVMPY8TII4nOdrB4Bb6aIu1yiluvlX6mf27migQyl4cBnlFbnQxeIum0XOcddUQc
KbugcCpFGtZ2yrVy9jB2WBOfXLDWXuIkXuvxZEB9iDSsLSx0PKGS1zPezsFZJ0Zz
f3vTdmlqojWNf6hPmlfVyfnHH+Jxss8jDawG6zHraYCI8gVe2G+nYLqQpj7rrMky
CSYWWGNr35EKQ9pKsPyLZjHRBibhvhADzOs+HEfVxAeqqBX6mVUrq6fN38rN1N2w
rU6Zefbsv+ImzxR36TzFVWRydq34sv85hBzKVKIstYr624z73ARcpNnQA/eiHQgk
JwTgZq8JfjfMsRjYq3ZCegsnb++Zlf/vqB2j+CO61Y/0AOhVA/zXk9PpexVMplIY
sBju3a3uOfHdzlRG9/OrIImBRUUYZuk9sCsDRbxDVA9+IsrJKL0RvUi5594MiPtH
zb6NryjBCnJq9hq5vs05RHf+jn8bwNRpLLXINlMhTMF0rCsRPktelBagM1LasGgT
VmE/p506E04kEVKgjBkMIfyvn/xsr15LsyZj/bIRvAFVMVtuyKpMsTzcPz+k1NTa
8wMKqONlUJOLWWpCl3huOSEJDXfSTrnWIPUzgjqqpcjj+I3pm6FJMHthSrvF1pMd
njV3+n5HU1DRQ8Mon801AHP7d+NGLqn1uw+SLpbYhrmIXUF0E5uxSumqIGJoz4By
KzRYrYbZBUYV02/dK5qQjW0NjdnTV2Kc0mPu2JFGRwuFEFrZsjelXSNPMTKxhB91
vTVmN3WWLcXHi726TOJZm81bia/3z8tSMen3mnUTJSLvpgea29mCC0fNEWY2R3ml
M8EolPoCMjpnR1LPkuYyNN37Y2iRwRHXH9XnNVNGpskgZ5boR6YWBIg/ejaronZN
evXFJoM1c4A0np+iT1REDd1CyhpaZdavylJsGm6eKOnTv+b0tSks6tDb9mjjFHhZ
jQHUudyVQIxnRzAMfcKlU+k2KQLm2zC72vMg/1SPG2SljOUKkWLZVJLixPGQKyl1
X1jNFDuCdfnr9MOI83S/VRvU34ryHtP6RuAUwlaZxMobVzyjvicDGBzA+tsO4v3w
zG0vyBJDoCzUaxsOJFqSaW4LmQulYpttA2j7zq8t7+g4oMG2VcFgSolSXPOrsK/U
K9fm/3AgjsU64IJ5IryLHUAsCnNr2jLuNV++HGxrm38VeY1LqZqzwwdVn88N9Qbk
on/0WqpKvqR2uJEqC9AC4BDXBtXEMTlMQn7/Qgskc/HYXF+kGd56hTtuxq+uIBXn
qg5iMsqrtYerw/8iJDLzZgDGA3noPmoEzbK3u554gbXMEftykuRmUw2WxsrEvBx+
Rlo0UKGT+RBs9l6fYSgJCmGV+nUhgxArWNxEUYLniI8+n9U4H0YU/ehkeREUGDdf
/38T+ZWc/FI9ciFDgBfH/SKAjUMLJd7Cod3agBi561uBgfBUjH3Yi6RrxN5dP5e1
RcYyrJonfi/pC7KpuYcLT8jtDVjAy//4gVKotLsEThuisVeklphylyadHQIdc+to
xvQzOTkxalJQXGQsc4DF+KxKTer5n8GvN6ERtAJ1eIl3KBQuOIRlTw69lRuF38Ep
nRgkxGCkijgkCmzBL+50ZarKaV2Yx2yeHNBDAGoPLDGQfay3VvWRNWE6N4kngCyM
ISmNqvKG/mzNZti+h2ZZHaY+zT4zxDbC86CBeId/kkqLnWa5HjCsKa+IHj7YTM0B
Esr6UVdKf0EoCSIfQRue+dx5ysfs8kaPWny3i0jxOicnafQpVmatZUKVsoqhC3Lb
dbDMe6Twar1tRkLW3R6O2/RqCOHuleNEpE8cXqZeUbg1QTr4tW/H/VuHbUjKi3hS
uDMztm88H3zYL81XNu9sNLm6yQYN3sniDAy1fuXb0gu1gBZo7ikfi8c5M3/HviMq
tIInxANE8XEbv3tEeGlah7B8l4bQbTJmQk00+ylLk6QyrOanO+hKiR2BQ+N+H5Mh
/IEze8TPl1/r6adyljDwy80QFq3N1vDl8YmpCwN74ZquW5gtS6/kuQFvVJZYFd6X
9T9Ta+VPURX4r11yFUWoA5CSLVSn073K2nl1fVJc+JLTOxTm63DZ+jcBhPJFbM5U
WD3HPHOc/l7vhqsMDeMb20TCbFaqal8gueksFjR905rzzGy3Z6zrlsAJtNfTiBYj
96TSHoXk7AGlXFHKHktCtXBlOKlkMYzXTJHxXHszj5bCfHmbvydTxh5GsSRUmM6S
o6n5EpmQ5Ulglel3AAzmY+oYKvK4DdGYO6IVsa21L51neM44x6+G+r3lw71GW3ws
LzwCilCPfDPbCHailEbnOS4ewwAKZWsqBhp5Fvowb+5beskhFpZlV2i8NuKlK5Lp
CCG+5fbGZKDyHACB9R0JZsYRrfoxRc8f+ClaaG7dt9snGydvyi+rdCAdAOltRM79
AHS2LSV6RkjVXGrN/qoJHFoB4Qw4VBXHpZ0GUgPxLqzjx7WOeM2Fl8lHGeAG+yym
YBuxKnKqd/BVIZS44jpL5/oNQzRQH1e7iG9S3kaSaNWl1cfEnKDtlTLciIpfmW35
lVbgT5iuYeU4NOCGudSjNZhZthQbg5MPPNq2GlAHYAQ/PxpD22ufif6l+qUQaBL1
KjM1T4bZj63nDXdaldf7rOTdJUfagT+b1OSeTyl4GUnvKQiWbmd3wC7/9MJgrXjJ
6OnrwCj+0JJxOtK+Pj00Y2HSJHJPGHMBq+/B8ZNf7k6P+zHTruLj0FfMBDErj/pt
DcIEsnx44um6BNNCebIlgMeDBV6KstLB4WaQj6JkhptnOpuAlRXhMlKhlEtkr+S5
cqrqT/UXo66ZgG48kZvcVufj7CpOReNt3oCQDZSbODaGx/B77leuJtvXikOuTq46
kRnek9Yp3n7BxksmTp2My882uck3rKqBSPEskY9xIREU0njV/6OOuQD5iGhRPE/V
92VanPJ4/hhkUPWsBMmEQum5FRQJC+Nyd1pc66Ud7LXO8lNzuM5Lpat+RawANrCi
O3YzJU1Kt0AoLkHkLyfRsvqL1AVOzehAycV19tSy9movYVYwuH+wrnlwK+HmJ615
pWY7ASs3DjZBwCURthNb52iaCNJXlC/Phe5d3GyV2dTdz/HU0yCtzzU/CXO6PKiU
MpcD3jrEXG6HF18jbRNHruatfHbvWHG081lgQFzsKUrKeAHqwCjM0FTY3c/EdnLB
8XdGA8kDonma2uSQ1ydnoydDL3d53pOs51S1hdVd+6bWgSO933LC1znKX1YBAQYa
AUCx4OYNn/LST7qvP4O6T4UTNc8PcApeeKyRFKKcINe/CuDe/dWJO78yJbfimx68
PivBmF6K32KA8788XLHim+NQKVWhOgNnL2xUnZVI7ndfWAOxOEnSJQZXKyOKWlnk
M5mYeQ9GiOx8uNxASTZQqiomdTqicCl3xGPH1ctr/eF0QMYQvvBoNZd4yVFOy5yn
peL3uH0u2HkQr+ogu+73PgOWvsmTPOm9Vki43hCCGHtrAp0viNEwVgguqf8w0Y0/
T71pUzaL+nQ010E0Bvfw39qlJZnD0OQLWQdLa2KLIVXOURybxxXFvgjex65eaeMs
kKMEZDFNIzFzuWMThJZQTL6EOfV8YfSrNewuhFu810O/lMcoIdREXzj8a+wc8z7/
SEPOyLx43ZDa+2/DRUX54ZhlxSUDdx8c5/6h9LJC9q1ZtSTF/BvsV1RlpYaWE4Ir
sujBgOcjqI9k3JWwl2y/9zxUYcEah2IZPgSlfM4CDTCCh/4Uz4RovIjvM5JqR3zt
ynbhUR/jBOYCeKVoQN3U+C4Skbnl8H9jTI6nf/VfMwctH7qT9PILva0/ReKAyPhc
TSbcxkAFO6M+m1tK7+BOLt/HFk+XzGn/Q0WK5BdtvICJy4+OoFE2aCVOqiAinl0S
yvYmczb+igaD7zBkk2Mz7xQZoTMEE4cHdV8CmsnV+WKTocYpeH22xn0uDUcJyTU6
uEfF7563dxolwF6DFpU80z3vFprKMAYElDWncW2ye4PG/oSk49rnecoY58jzwCF5
EndcHTK39H2c/fssmDeHb8U0/JRZNZ33/8uaZ6E9XyJC2Snde+uaISjShYTvIeXH
D1adSMYsDluqqrL+f+J4C8YydpDF9Q7LBQ+ohhOZQKrvNzsY8qa8jgGLVdR59Odn
r0Lbd+wqDUBc3CfFrPGPxEQ5hQrpWmSVFQ2ZyTDjRABaeT4bxjlT8jIok/3/YcKP
s6aVbKuTCjpKMJLJeitUUKIyAYdv4+3GJoiBqhn+twwVNmsn4u/Cnpb2ul8R8BNE
TFTe0FkzsLwxTzczAZd3kSn3hXeADHdcHdN3p4j5Qwi30Ik0cGm7DfVdm6a0f07/
GAZrpNb0hg9d7E1lMP+4k2GNP+7cSmdLAeSCrtUYd8zDY+8WTr+8RjNB5KnCAO42
qKnHDG2iHy7dRoNfURbdsXkHndoFSmUDh1zyqEWlfW5SFbi3qpNukRykuHxZjeiF
ii7rCQumjKLva1PYlGaL3k68dxlnXXScvqKEUq6j8revl5sFTle+kRtiWVQeAayN
bIToz2IYqoJD11hzwqXjNPu4xBA+HUHnDj6jfgX+T0exZKb30NcAOebD7GkwWNUh
GSQT7IyPKQQ6dPBuDZPqYM4UFWGU3yGonxku1uKiU1CP+It5/kaFVDPSzQacUB/Q
ko3l5tWN4U6WLp9S/NEWA6AzQocVDCWrpIgNUmQ4b2iaMkcnOC0Y0rBhNu+09hFw
8NpNYEbEomn47RwBFm1Nc+9TaxzhnnDoL0R97D2+e8qFEon7g4mtNyZrS3kaa2dP
7jLGdZroP10dqcoTliInnBJbC2nBlb6CYq93nzUTzJmhWE7gl5SHD6TWiJE5xogs
DREUVXZeYJ5ciwx2kayzcR0Qb2tAxT3WdLEp5WMacHZ/y7GWtnOR2Batq/37mHz6
q11vtWVIhKQpOBVgLtb0VTbAbf21UxTxrTyHONaPIQhmEPifWekQwitVse/gtWtP
5PWkd2bWuYqc7sgKnEzkPLohSchtc+nhPTf/yYZ1ZKNJbuXC3y+lItY0wP6cRGMw
44eOsILaUSfKjWQPhdDUUcWiUSAoR0khRwYIzNiXJ0ScVfK0YyuYFmxk18lDyoyo
BoLY3bWqa8/jvNi0CVb8pKqhJNF+vuKdSp9IfYfblyWeVDJFQKpkqvAS7LJoeQ5k
MVCdIyPtOhin8LbBQnN+RdSUMKxJvIoiUzUFC+ALcgQsT3J1hu7fgPiPkTv20ZLB
NMyaWzpf/lwUxdz5m5HNyoMHEf1pco7sxm087kDhn7ckPrcbk7SiD2m6tPkLpvDw
p8TPP3WKsU/1fLMUtk9BH1PiTLrsGJhhH+LiRasXYr1CwIQHkf+1mDv04MKzBZDT
VV3G7g2JueHCMtIif/GiDu05LZusjrP1IHZv4x910Ab2kumCaNGUt3Do4JJIQnT1
w3raEMvSDyR651R/Y2ywbj5pt46Jjva5xHxkpPv4S8y4/dI9qS3etx0LDAZCDad4
Rqyx/DJ3J08mKfsiirSiVW2RvLWU61xGmoCNEdojTdu6jlthI2WslvzZt3bT0vyi
PUULSiF9Phyo29gMXUwx/+jCvjxYwTawTCTmT9QQlPqJBgR/WN/dXRUz7YF6uCQ9
gq2N8LSzpK17kQ8kLaAt/a74n5pkz+ynwYyLTleqAsS+yDb659Xd6sd5rqdG72NL
men/EZovdDWYPTIBuedoS/Z1rwBa+i3PfIpmTOync+T8lF92O5rAXybQacDi4yYK
MiEEALRFF47KjqoTBdimkzymNSACxZMl2j9PcBN+Tpq70/wMAmwIKL21QxIP5nSb
HgdXiYr64t0IoMD/I9K8qZFJ4aDD6gc7DVvuvKAw2JzEN6UdFVcYBMzAv+8pRDNd
JdpVoqEqW6R7i7efKuJWYECUAqXwn45rlaJNXcFkyc2kUWHuGJGUvw720VID2Av2
RQ34bZfs5uBO+7r4bL9nK7sJ/55Ksu+04SkgWf31P0X7B2aRtvQSzRq9DYIMR1nC
7wo/iceJaW3fFkhcF8ZaMxZsG1wb8Kp4FAQGK+nq2c/59/Jqj6nbtsO+/XVTeMov
qggqYVH+mO2MYIjHv4OR3vSa5qk/i4+fl+LkSIMSS2suPMUZVDwsBMe5Vzb+5poy
j+DIZV4aiI6nHtxpx6EfCW6reFadYvoBUavDmyduFxjVGECV0IGbkP3PaZpQfT5t
GmsJxNTTkplA8C6fj/rUizZ3mxGGvaV//23uKszAoPdteOjKR/4GQyGeHytnQAPq
QqF7XrndYYc/C58H+/hD0R0+XzwQ6WkdCiLZM0WUUszbkYGHG9mHwLzbLzPLcc+H
Ihb1l+3yMrzm+6nI+NIgQiyE6FLxquvCQWxD2R036tSyPLXjdPSBCjhs80Mq9tIM
Zejoh/W1MjNaU8i9wBf7utDn86eMFQ+Hy1/g7fOb6x5lB3RGmiONAcay++PEPPnN
xS7yC6CM08YTTSjSUfUFqww/YKjFIidSG1VRkGLbB8KyiQEKAIZQH1l5sk1iLqvy
eXP+EIm6vPQvP+SRMkKHFDfe5sD2MTkKEiNJ+kwaI5DIUtigDiqAYrxavpw5dG/U
NKf1nBiiRwqha6MzKsZyURxnD8swr6D3Np5HIMyOq6N/1XTQbRV2KZNSNRpv/QQI
1QT2tZmVBWIhaB7JBwnMGdvwK1gt6HvpiwnAGFfRLSxY/+ANpLBahBiCIFyDiPe9
UAlNBkNywYuHxsVP6AUSQYu/wUP6OyIpRDQB2iCQ1BUaA8YG4Cs78GOEWVGlPj9z
gHCj6zi2NOsJQNJZra3mVPTEMwjTPB5Qv7lG8Ss7YkTxqbQ92qylveqI1dLdSwv/
TgkqRGzTv+HIFxOWe8STk0K8xH5KVrtQyIr5ONjALdxmHRSqmREc3sICmOlfAQOZ
cms+FHwPuL/yUf57iJgAKIUy3rfliFHbevso68tMtGXmV0SJDnRmCAu+oxROXYBY
OJN/xIoYUL5gmBKqTHHbHK+TKwczSBuvpl9at5xOqlrQofORKjzgZr+6dGcUm8Pj
G7fOgiaP6RbO0UVgSVylz7YIUvJ/WkgGAJ25oa38RIr+cT22AlOUkU69XIJQS/RA
c/QzW5snFObiO0elolGeF35xfLjuxP96+obYreA/gAqyHtaeyteWE7PCz3bpYQ37
tQPZSyx5ogwIwDCBs2mRloK0HlCbPdKOzCJ2Vyi/NgtqQFsFJLkPVdADBAyXIsU+
sIElyuB7dIfwNZsyUFKRJ4PsbWhVtqWQavvZFUkd0jUECihUsLUmZHRVwh0bEzn9
6ZOBMTAu7ESS+mYxJN5ALR9ji6LTyz3KOaiX65H53tJgLjfREB/arSsVek6rqgWH
Dy5LKQDrr7Wtn9AWIWFWHxy/VwEaF2HcC2WSh9zigXsZq29n3BtfbQoN9TDzgxy0
9+w2NuNzPilN7LUAF8zljRthpztIlbLJvt4RKif+NEldNzBbPgLX1VGjXylwEXVu
7osel7T8/N+Cxzuc2Mw5q91oGtDOMq0qd4rDRnQ3qpE1qlQpn81SARRxmRZGfPqi
8RsmGFDrVUBEh2D+k8xhbNfqaLlULtPqlrVbKYc+kejo9B8NEVmRwarrvhIw4o8P
ro5RY+wTXXaHpZkmm4QaPH3mIxwYXy1yc1E8PeBMTMj2mOFnlUw41oD/+xGtzbdo
orEUjnfGMyeS3QsugpWtMoyOaTFihgaWI0MBjUzpI/kCCYODgaUXY2RoaLLgTwNb
T1hC37Co6zgZbWdrNjuk2u1HO1v2i5ZBr5y6VyPbfoaSnZ1qz7IYgrGMxzSMs62/
3djD9DNfhyFERAFTS5c7e0bh88zIjM5fMuq+xO3j+BWod7mlpWqJleFW/IBBAV2l
x7V7ip7qcy+g4GPvULK5eGBfLsyaXnfGuhH3VDYxmxPSZ50InrT91YfP+OsO3+3i
3eRW90cgRrSH0o4ZxKr+Y5a7RJR4yWIIHc6WMwgpsQhq47Lsg+iuTOxI+4ZxdrvM
0PptbxfnSwM77l0gDS4IoQQ149bHa+H17uyGC2hMKjMXnZXyURe2Vi0j7pcA8ONt
FCjROgRP323j3zpMJab2JIwz5+XtxhUvy9gOzK8tzvZQ9wiehTcpDGk3ZtKuNbva
Lns/bisQDVx4cqcnmmlNdfID9dKd/ti4PQpNGBcbSaWf7vWxeS1qwjqkY+/cqegH
lH459/q2Kb+4utJLKONgTSIZCwS+3/dD5SN52zWjV6GclrzHLCNU6EKcT3lE/NNW
81j8Uu1JCupzUI297pSDNvt4I+OTns1oVmBuZ+/u7BPbPrgSffBg0Q4RD9ZX0kop
7tzoyIGB+PwhQ2h5mHH+zec/W3sDe8SMhl5p8oP04Ze6SZxdCfiCdIxIsGRln4dA
2c0B0s0arXUGDMpHMvG7qP6WmI2chvPdrkYdPiHpbNqAbqI1NR2wBQ1W1QoUANeM
PcBnR1zpWy1Alm3PSlbfJEWaPpLADco2lar6zRftgkZKqnkPNnC71M6maxPZzS6c
WFXQQIkR671m5gLtmZwrk2zI4cRxMfrfvBTT6zPYOVkHTrMX58EVbvXKnCx5uusw
uiJO6jziHF7JhUw54jxxS5CbWgBRtSnWToC2vDa4jAzvyvCgjSO/xCq5vqh/GS3B
TzpAhUjf0pY06r1TGAOGWsKmKjVy28E59b32N9M9wcjGjNcR60+N4WPxtqAG0qpc
OyP2ooIcyQX7zhKHUvy+MnJkE/e+zSBXQvtd2pX3cMSqyAQYiIEyEAhxLSfDX/wV
Hha+e1szS8yspYS5SF2DZWgVPa1eFOF0+T5LUOV8h9DbXyYf0iSAbu8eGYwJ1MCi
MxB6zQh1iwtfgjX2/P/OhaBfza+QsAeLTYq+VXlTT8TjjaMnnsySrrCtfiE176iZ
rdRi82frQuYowNJlCs4kArNcRKprqv3KEfLVBkHq5julAmH9P+MFEHpzShVMtQ6e
o1S7ngQDR02ZMXM778Vet0UDHUdykMOMas6VdvPxY4etCxX6MeRFvj5e1IJfGTD/
Ymh/y+RTriefeFlFNgDACISHghwXcMXnGGqw4A0Wp2cNqTujB+EFyWcK9u8rk8Mb
Gf8lTvw+sNiHYCTlbwcO9T3Ay2OZeuF73XXE74LWJP+Hv7dNu9R5rCI3eJOhpcqu
dQBO4T/BSh8XCRd8ksHdnCkDM740CA3UK2aCffcv7/sb1i/2JDR5d9ZFncTpFy1B
26yidyQCD12ze6VY+Av3ThyjuoNG9RUEufxxsCuQSfNIW365a1I/OE8+1b7hKffy
AY4kO5lKrP8mtD6LCdgYfPSIdNm1ZM9gNwpZPgEPokdk9uU0tCUfmtJMgQJIcTRS
tJg4rt5SijSEgG0gKqrUOXLn3d2Xf17HojvO/4xs1q9WvupPYQs4xXEQDt1AhEU0
Td1+C01R78ksu/eeDkZSZruQSU2pA5F4UX0IXm4Q55vTDPGyZRNTQl4wKVL00ZCo
3Dm9n82eEzFObkNUvSxb66zS3IfTuyY+7IXAosKTT+n3Pz/UE6qEF9BMeIfaU0Op
fHQI2f6QBkq0IhN1givP+lHrTmG6WTtbLhYSVcRCUBg1wiV3CPJjwxqE047Trj+P
2nFAdaMXlToBNLMTSwHDbEuDninb7TrrxWXplerd7gVe6NflIEgzjcJTMLJhR1Dh
BLuGGMm25/63ERJ1FgQutfWE6ZkJPu8hkn/howsKAjzKAzYsE9+nkNBBXnlqwLjC
yFNBjdT5mpj675ffjsSzMyegThgbf7D+1ha+YiDKk3IiEqvP5wIH1Rgc7oGaqsbW
XnQ4+EqHguvTSowy1Kna5zPUfWRvQRi7wGcqSdqpC0NWN29PIjRHeKwpC+JMj1MS
/d63HX+Yr6JHUTyseI912qncBFo7FhPL3DjWZMrYw6YPjKvDLbNeVwXJotCteUfY
zxBgTxrG/hnw581WcaFQbVPqCVsiIQK3TlEaj7G2oAs6ESwDx4/nbEpQiuViH8wC
t4PHdJJkZv16MebPzGpiqDCROrWyb+pQTJjEr8yrbfzb12bWW5RMbx4TRXt5mZM/
hm6gc9C0dtOTJGT9wEwu22Kcb11eGHWh8uch/vd5cYu5TEOOZLhx+NvBjALgPFvA
Q4d8k2wHef0wDB9fpytlCNzZJ1igaHybpmnGcOEpF7GjxOPIf9X0PsTz6bejcvqo
hohShTmpjfxAzZiJLrpaWnKUvZv1LcrJfE2lM5dZZsFenzxNdDljhqfD6J5tntYd
fi48cysooJwLvgtHywIFUW6n13NRqk0Nage8WnqMfk97l066ggLZS5kfqg8WOWdR
20lVEIRbR1SuzSDdibqgy32y3ptL4JlkJ8CC7pd/UfBf3ZCMcnxn1iweQlGLeRgz
Yc1ns+gSke/eqWUXLRPkzoarvfxDRrIhMUc4aNqirTTPufpJNJnAsaY8NOjZGic1
VQvl7d+bIjI0a29BKDqb608wUQyE499Lhbd8f6vrGL8Woct6nkLurrt3lsayPYzu
5Uvo394pitYjCEQTSG5kGd3geGi/REqxRk6NbMU/bmlePTYS3wTqah57x/OaXDLt
7NJhuFu6OzCAKHIAQ0rJqHwvRWXvpasZgqJKrbn9ME1wqZFHGbNoRYNNx7RuS3K3
4Xa3dPIUdsPKnprPNXKe/VA6+PqnQWn+KuQr2EjlM4jO1zAnNgO3jIvXMk0wyUcZ
LZ8SdstaNbvEf4n/Q7Ai80pxZlSbZ1+RrjgtxeuFZxkRHeGdTYgGQ08TQwg1zYl+
R/aRzLZ1kCLS7euUmpQ/5Bvem1otlV04n4yN1OzIrezkqZvvF/9itEbYmE2Yd04z
H43ZZ+3doTwBMJKQWHDHAE0Syb0YNMG2GZfcnT65j72a8WCIeEzpKkBwyMiN6mCN
dPDdqDYL4SULhe56BQOAuTPL9N4rcdE1e0IoyrTU4a5zo/FMRgEZd4OHuuAfL1gO
LO4cVdxa/65IIP2pWMw3xWnVmpn3+XRkFwrIpSa10LyityBZz5Y7klgIkx8y46nM
rm+c6mpWjhWQb0niYgu+aQ0y8klCVvjhSpjbgmIrtm1fA2q4AMwdb9ZSO8rTmvq9
PjGfYeB6clKoidQ1wfTxkASxZ7m6r8WmSTmawssyYcCEPGMGvdKSwgVgViWOr/9N
n0s1HRxwLX5gJdiJei75raHSCMQuiusv7qsRMvtdMbt6ivl3jEDfYMc04YeP6b6n
WW8uz4zvmGSOhb2Asn8it4nLBBjGjKNruZogYNXSpsC9D64jjwOc2V4+rHZR8vTT
HhqV8KGoiPemQ/OEr5JSAZWxbvfaKNf82WF4iXnQzaZ9u594TY0O9UA5LBS36JVj
HZN33iUYgRl5/iiEl/Ve7WZHy3gSXatbCS2SwjSvHNpODlBIvkxBjXDyT59L6efc
FKZUaQXTxhCyjsIUuUEthiS+CfcyWJnC0W8vdFqUeVNIijq2WPytzl4ZRAjEU5QT
javJQ7fcngsb2U5qmj9iB1sjOBepaoYx3AOSUIsEXNn+B0PhoCoujOjWx/C8z0fq
CUd0Kf8C/28h5BPM543Cc6I7yMqsPRXsWVRvGaBMaGUC4fLmmEEecf4cPD0dnTO+
BbGHI5CUoIfGU6hs3NO1zem4FHy5bQPhhQb6dD7Qn9yYT54EgLDTV5A9CS8K7jiR
UvMPE3XM6kPqaRQeqi9CFoX9RS6f79QzrXBcMxw64k4sV8W7SUvPqOc8mIxhQXNs
KvS72bg16ZemiRZCNXQAVVQH8nuoQ3EvTGVFTb8Ec86zJLcI3kf1Jecbl4jntjYs
cDTRzdtsYf4maDFQC6w/xmbEsBQBBTTnT1npKGhkwZbrka9YTjtXZ/jvDTZNYxO0
iT2qma1KEGgDlJ/07TV1GzN3uFiNKyoY8Mc7zynEhuamsqH1XCoZ/gy5f/zgK1GY
q99m2fKZ5HyTKsPtO8aXpB7IwU8f4gnVpVJ8AOqNyISNJqZ4CMcGFp8s+WgBHRPj
9kdG0NS7cHLbyYFABd70XOYgYF4MoEAvt43nnnLlgmOg8lUFiV3EmEChonnRPupZ
XMurKd7dVKashncx8Eo6lr4IFIWvShh5VrSSVaEJvU4zNgiZ7SbaK6v+w6Rnlswj
lZ3MllyvmGNBOACXRPP2kSNm/pOZsKfA6Xu2vZKXzXJyMbNtlg6QU9MEmBAqJ6UT
HrTpFNHOIkx5orZ6RId8jrdl/oBJ2sGkMnZ5tCLeyDgrtphqSm+4u1VobzzrKoBV
rUuOQ9zSMCsinXY+TY90jJkgcFyucfnJeVBFFBFjaCaBGwDujNQPU+Ht7ONhBWp4
GwAozU0FwuKahB/4VoJxjuUTG2r1xNOiPHhzaULMkI/2Q1J+aju/oqXJCuvJMp6K
BWJKcdt6nOlAfDjfqFRIHHJEZqX7UjjrF1+mgk3vRRdPuQ9dLengR4jWuj3Ar+nj
MduTwD8zVJVxdumOKR64MRvRPCSnhImcpowjsau+eo7iIAmYjdtPUHr3tBfi5ZQP
NHruPcBXR1qOQHKV4U4FqiqjqU61BRk3+OwtPrH3u5uySAoxSiTlMNkXNKEVNuPt
m6GW7RUmP/A20/WhLZoEgtz42Qal0gyn8EXzrLzg1oDAIAMSoG9TZuOD6Hh6GGUy
9kAbFsNf/AEaJx+pgudBupGisOZzp2x64GPYpyPswio8oVreH4ymURd/AXE4/F5y
E3bxOx8AnPk88elBPkQpAstGhieBF/ytL/aTkLOiwiprnsqJaPPMHfMGd48d0n+L
M/vmv9VwkRfMF9SP+NBzYVA63zeST9DqDSj8ijWzO96392pUCmvk9PEWYYpeRu6B
XsJm1iVPgcoVNvf3b0tGp1AwH6g0jwx7B90DkHszeoOHONjI9D4qQc7MBfzzc0KF
J7a5i5mmmuesqU/OaFJZelTglPfYvSK9u+Y3GmN5B/jh3JjPvkHfsUBjee9FhYJ+
V775ZZUVMsMPClAQYDYfTDoHi9aDJcRcBOayu8OaQb6TWCjIAJwn/Hi0rAN/1qJM
rLq0PWixTgWK9H/viNuzs8RvEwGqAQvLhFBTTYlVqEPRMi3JoD13UBxaXP98Zrdz
+MOBSAri7yWAEWjrqH2qmE/9VMfIQGRyzdDDuR4xJhKM0hy/W1LnaP639egIosS1
k2pem10pnA5e3ZrnqX2L2lSYjhqGSz/0LoiVCyGqrz6pnsOPKKGS69hGnoQ6Pi8l
etGOp4bm064INHPpeKHafWp98BK8D7Csb2mQeBj0PVddZL1VfhL/fDaszbB9qBA6
YOadHZnEGA/ldinOfH0FVQq2hDwsRa/oFa9rRuqVseSuIn2QEeqbe2vmY5DFowIX
tUZ9Vph6FK451qCZzwG0qrTY4+EMz3JgRJjM1sqFwwInUOwsxk4AzA52H98WMiuk
4hhPMuXByZLIPoKYx9Xqq3iBoJMWrSBog+B3wSXnJMVPLs9uoujptRI63i3TxUjD
QOSsc1JYhDucRZsKWWMSBjWwHVup3oji9UO1l5JGSsUbDcQGPTuoo1sE23f1etxn
1Q7XFp7ntMKfkC0w3wxFG5HVjm+tp1UDi662gj5xg0kOPRtRNblVYYdwvkQ2rRfp
6ZA+B/dOZ+4EgAOEgR+l0cp7CgPRpM+qtFbYBepVk9pgnrzxET/xlaoTU+S2dus1
sNCkP48IthNh5hd8nh2mpH21KrP2aGoFA+/GvayGdVkAkEl6u/JBtLxt4m0LbY28
zId74bfWyJDyr2Ct2aLYOibmqmQhPcScRKRJaZ2JDT5NjKyFCUvAfjCg9HpxnUcp
PT9cxhEGAC/Pvly/KTHAY/ZEJVBwQq5m3qEh9xPZqMmaHKLs2h6z4UgADr1yHm6Y
LZP0yAAocbHmS+p/U4AJZ1QxLqxMTMhcSFdLg4/VIrGC6UVd+uNxvHShr1/c4zQU
HtNs+kY6DNla5+4YFFl3vWKO7vHr5FP2B+bMcP+3A3+9A4xUQqvdfiZaKEhNrRQj
svAmmBSKn9R1F9dQWP1PEkEJ72trTB7oIZidA+CXR1Aopj9vvgeFjAJpPM9+geYg
gIZtIxLCQzdyeqPGr7IImwuoMvXSN2NkWAnkycnIPQe7pAerGj57iZUjhK1IePOl
ct3qaQVqaMqLXB/fzUjoFsWHC1kXxVT0CNNxR18qR0ooW351W4HStYMJeoTI8Idj
lutps6KL1Bh9D2ke9Y/Sy5TmHBCXolJfa0nOIqn15C/I2fxLSkbzhCxIHPkwWKba
hNNTGpTUFSNlkihydZUJ39Yw8SAIquL2jCH6Hk9zX1vU8GudJoov13CKeQ7JDuME
JKVn+Vs/bR64av5h4K7rMGKvh7v9nJNnfFIetXDVSj4Zk1FGHcTIT7ZfND+EV33V
7q+jZbwIExjkqJIog3C/NXGphrJp2c1zInrYRrpSRIaf0+lbv84bqb2XYorr/ScN
XD/jwzoeLvv4hpDFHcyILwmoVv8DaSPi1Cw5O3a5EiSCOEdReZRNAG3fFr62js/A
7k/E5ofVvQOZ1AW1iLRmIZNngvYkSLtcvVki8FHu0kWTAdhtFSD82KYp8592/4zP
4nA1NyGKfSp4GdDpS3GMIwaYd5HDxsEapoScgTKCN136N7PCR98eBqXu3np84SMB
BhVhYsyFNBYuCsOrYJrGq8oJ778anzU3zLsJaiIHARW4OSPnvoyWTU0ylZlDm7PW
r2CyQd0Qbdj/77CuetLOYpYswx4koQPOVmFhtfPqYPcHZ/Dz7qe2/0bEDvAeEJFf
5g5bvd8CHh5m+FAiHwnVXXvc7c+28ro7YNhXR9tP0speBihvfzgEeCRfABJKyWTK
GnH/8+h4dogyej6UYk9Vsmf40nhGC0diOrmVSbJATnWtVb1zebO71zAriJf76Dng
6sexedFdOVQ0d1UXFTUp4aeKoCy7ccjqiWAnzgr1CTFrzZ6kYLFqVzvTZH/ZfhBx
WNV2VU1qHKc2K9i6dZdNGPqhxqiS/phvlYWdnWZKAkWqJgIspGRNGDfXGAFuUyRL
ffwoa0q5w/T519OHYZTcfFzwgZrdeLZYGUiJC34VG+ij8wkbZdMT3y137h1H7qyp
uQO4nkOaWU5Zv51VvDox7G71zieY6fdq6V+VxJ0mbdnGgsBxGSpqcqjjpQ2j25tk
GqCJ9swHRbuTHMeH7G7xVZKSP9xFc7FC7DGFixHIaMvzN1ABPRhVrnNM7rnqp1AV
ZQZxbLIIpWny3P+k3d1stfJ5tQbYIRqqT4CfW26FiwFtbJo1lJwzZpQV7xZSNxES
L2ZadhZCISiv2/6joI6AZdZWD4xq5KZQvBkI7i1Kg3+/QRxVcrormFV9sNwslvB2
m0b8ZVgK1xwaTl1h0SQgdt0xtuwH7t+B13mSE1BBHz4vF2keCvcfk9M2Rh4eMgi2
Y8LyrT6fDJ2Rkf3H2Up87LaQlXBvIMWDffDXA3Pf1IDV6+rcAzLFqR6PmDPWkw1Z
3I5zQz1LyUiThgWAYHHsnaZ3NSiTLme1G2luB+vN01FVLyDpQVLS/WLIHRE8AYEo
oRHeXSs6hJ7Q+UeU+J3nodjVa9cRfJ+p6LR5+G/k3DOImO7zem3w2OoxQ9ScFcq2
Fm7HEqiZki27E7v4Sr2BYdVYohMC2DC5dj45eoPmn4FCy21hWfRk+RpFkOgOgFrq
IrJrC3thf+B87gMeaucdJ47MXKu2puUDSpDPDcqs4EyexDnRKHvVhf7LBzdwnSfO
aJT2ZF2+AyYrXgk54jsgSu2wcV6+TvTHZquowB/wbR5HdyLwR4Dds2pwjpzUvOFz
nQSxaB5gVFdzkfWkS5hjSVNLEtkJxUN1qYOR40j8DOP9hxvXQmhF6A26WSOjoLs6
VZGAtJVcgFMKEbnwSjQqpzseWvK6pbM39JVvh59twmwHqdedv/0u7fhvfW1IARhQ
OeIcTobi3lv3jo1AO+X8/rE6OGduBlnDaHDW0mer1wqBPNP7iJZXDv1X2JJbIbZg
MqqkQVOQEUme1V85aB8zt5Bc8qciCF+4AbITps5150ZpieBRLHd75Rh5QnHmyEXi
9cc6avBFvg2QDUaV1axJ63eqJbeq42601AlaztwnFIWk9XD3NJ7h5zZ15cDTTF+p
FKG2glSUvxgYN8nnBeyZ0Z6scoScoPN5j0EOVi9dU71UywaV8nVDfyZ4j642qgRN
At3e6V28CKgyUZ8lwi4jkiwhWr6inoykNtnDCHU/XsHxnyufXK0kIVthsckCV2AL
YzzV01pH1Dm7bOnxXpMp/SvikfNL+mkhRVgFn4kzowAmQ2nSu/ppylJqnx8xYjUm
0RLm8f+6NS+V5I231UwZZU1VucXRQCWHg3V+HBZ0pL/RRQm3Uzog9VbzvmwDGI8s
VBLH4VTePB3NZA2PyZFh1csqrIU8wgJ6facdMyXI2e3WKUwlknqOQ+zF0iNsdD3m
TtKmaSPgT3mv3pckgcdkaQZ8qiQi7d3C1/1wUpD2Rd/Z5edcduX6oKARhBmFxRz1
xDbE0xv6i+ydOAKPZuENrNVryAbxj3Sqk8EA7cjCA7OhQC6lx2Y/9P8b4JIKO3z+
JjxE9WReaxUecgU383EDbG5v+faacNeRRxxz3Ngnh1dkWLUXheTZ4uljT03sptkK
HV/uhYGSczNeGc5jOfgYwzEfC/QgXrKRsvqT6DLqYpevg+TkhtGgj9Yykd2PUEad
o3C6Rw1SicIakAzdx9uP1O3mOEJ90fJSto8P6dwy5g3iZfQFn2vyqvzhJQODxjZ9
fu5H3UGiWMHDzFXh47cHdmnb61l2CXbxs8bD2Zzjic2WTZx992/76vC1Ko0n2HLz
WXFu4wqSHPEZ4s/bnYjuMVCgdpV4e0rjFssPDKXi9r93VN1GmG7UZ8bmmezJMyEb
hFEz+Ik2fBy/1MCogUKDu9s14eRvVVwpx4/G4raJQq5K8ruXJSWo9JFsT7eYdPht
xnTKZpfFl6j21kVOiG9z2YrMyOyrHeHosgqOnDdhUW8jHlqagTXmyGUC7DxeKEtI
qUgGu/XjIAXASWw444Fve8zi+wdYSJApjnt6EIJB9y/8JkGDAFQonu28ZqyNSTW2
1ZMcW9qUftQRfu5PglUZU5g4C+BaGOjw23P+pe+Y36+u3ejdwcD0Bvuc9ZH2v/69
OC7G5Gaj+i784VphsBf8j/bmYMO5lwZXFgfAUlR77ghOu44Ep0zDwVTcq9H+MZxs
Lm5SllO4ChRVQY66JdkkwEibrxae0iBqbS6u/FDmj6mPZ3BMUgYJwXPHEzZL0WiC
X14JVEXSu9vfYpvPSAaO+TYlj3aNu0OfpWhyyesPO5Mi3UBzTwzWyRA7BeQPzg1Z
C6OEzhWRzliBAreWsc/RXalponu6lmwBoE38kua+2iPj0HwfENnstS9dSLl6Jkqh
rBv3wDeaQx6IchIkQs/FN4SBjGzWu/dQX6Ufwy/0aSHBbBamBvDJ6ErSiMEm8vh3
Bmd0ksP9XOuoJpjqD9GhWx8DTrl+q06iENkpbjBfKwAcKirE7FmTyhKPFv35/m5I
BqedKhkMNbVTX/GLZ79JGXtybMyQdnOVl+dxUZBDz3ZYZ+/3ipFuduRgonYhffq7
mIl9jD9C6UkmiZkoHyg4fqgodWwoTS5NBYlYG6SCL8vKp6NHOCFJgD+CTSEOoz1d
GjFEoG0QcPOYaK8yodGiGvIEf9qRmGtwHNw/QKk8VhPrwzer3G5oUb57VaqRrBmN
swooGK2na/WSQPTvEx4T8NoDs6DDSvlX4JIZgthcdWhGKJ6WdEPuoT1yMOz47rby
+9WfcGyioEnG8GIN/WeypIFQttKjmJpyQ8LF6m8aklxpf4AzJr+lAYg+YgyNi9Kc
LHzWzMlKm1eA5VzExu4yjg9MGHOU2p1C6f3IuJtmcl7k75LykC0qqgYrr77l5XKb
ikNfQo3XtxDVqkjjNPhLI92fhZNQNhcjzhSBU5w7Vs4rlDuxC5+KoaS19lREB1k7
SMkZYHW0fLXXFlydCHUKfMiogD3oicnZ2a3il4+aRV71rRI0JMNUOBJci1PU5qt9
kql4re2caS0dFkV+EP/d8sCy9aWJ21ZwCBYnxXlMNKr9M1JEOBwsD0Leca39C89p
P5h3hHGeF9KA0+EX46a0Kea72aBRbx5zKIYD0kKmst/PJZzOwmZIl9cLXw5C4SaG
BqEs/QYEAlmqxThr/NJrIqTM8AG7zoMgwzc38rx7fSLAfA/v74ulWxTW4COWCiB8
DbEzqR85eCZsT260ilwf3v6wNxDhBas63KDdUr4Wa7KGsE22S6vhbpZzUetPb1r0
1PlfswWjvIM+EP5TDaUH0LkrHdBoVsi3KN0EBMxvznGxTGsuWIppQ6mS9Fl5NSup
4Y8DFBRQ9cTIGI9+IIusJIkR7S9dY0ER1zDYVn19mwA6eZ1gcB9kaV2ZTLbWHdEV
WRaHXo1jJJxZRR46ilWui6drCOCWQY5GLl37zGaLoS7UmpEHc3MlD9J4ug7XzxAB
BLF0JzNmmp+bvhwknhPqf8H81r2sjcwwEWYMtoEa6bdH9YJt1tXfLlHmA7QSZ0qa
LTSbpsIkibIDjaFyY0rWdjiAscbCnY6dHcjGYET6g1JSsFUgtw+A9LIi7GGCKEqg
XS6ZJ6clAN4+XZV0cdttDOAfAqH41Rdm6TaxXegwgVC5RDaO1FguurmjAGBb03mj
AGZuHOmDyV8L813S/kVI6/okVgrGwn8LGJ1bCSWvGGO/3IPB1NTL8z51wq0IZBdA
CtMxNs3ZY8roWmh6B4itDos7m0vTVfMcQDlPeMxx58H1N8nN2ZmxOSTVWHfX6BdM
VN7EMf4W8lPaP+p7nfW9ddum/ixak9FasPcAKJGq63VVmn5JmQLC3RszN5tgphoz
CWm/FDb3nSgdSv6zip2pLq7c3aXASJa1m2Xa4ACuAQE+hfvm0T3n2iUjrs+uhycf
URcwo55of02v11nngcRhIO3SPDVgqNCw4Po8pWGq2vt900UY78+Makk8fMAs/WEC
h6rM0QJY+BNAzrJpYLN+Y0HeBEwS/mimvqrHQvjib9a11f+YlmMJdpEcFhgmEOKX
n2xZCA+ip+ZYCjxMOx6QIoP7qN9iDQ4TjYarq7tEUL7GPjAJPJtIF3YHHomyO5CV
jtrElR+WS2WhNSeI3YMd3R381LRm2mVlJO+f70hi+HdJ4+KztfHPnXRuAAmXJPNa
sKtL51vGPXA2RgU02OBXZrlJJG1QgNQz5EszV+nfNTW3dqwQpgEqOjgz73T52C4U
rHVIRWyD94JVTjQolZhpK4xbXlFkCNzT7RvWDNy/QrRaSeaLsjVShjHvfQpylNV+
V6FWEYd6kaecBelXNZo89iHb3dkTKSMwLlmgM6DYS1okNmtD2bJ8Mb2czPpUUUUT
KL6R7He6xd2qJ0qov9FRLvgdvKaogRJWS1LolGxex58Snh9JWEl+4ESlIbhG4pub
qzTG3kQOPtBRrAmW18yxv/KmNA6TJjCN1x1qJKZR60m0Lo6iHLahYpUv296bMB3z
+THqfNJYLHXny7sFY4pgfJghIIoNQGSvkRHZ/KCZ3VBxW5pwsY4a+GAzvY1Al/E8
M7ypmNMczIMu4eLbAHtbnrVRUZ7cffxT+hhzLegddiKvk27oC7aSTiuI/DKu3V6g
ubl3qgRXpKpmFEUyIiGvfGnH0jU8AtaXMTl0plNlrPRlRqfxKZc+uf/y+I/pxu3r
pA1zi1qJ8DqiOO08L23lTVFQQPU7svqGURkJL+ziy8M16IwZRghygIoJJppXSzaO
f7StSkel0xroF7igrshJtvh6Jr2OEgsLXcJNXsiqkiDXmIHxbN4f9savavFED3fB
kHp2dZ7D4Or6MV7JwiqfTSrvuTnqC2Q/ffZiU/6UUYQngfFVxvdJD6CVu7NIagh5
JRJlR91oUuKOS0movcFMcN1T1LILRpNbrjR9sTlVwEQsav1n6MHy2odFHYfxSRqr
D1p9iKKMbp4/WYuPx7ZGA2gyIC0xkywd27QgbFBXZrpDpRLX+BLcQE8+BzZNp43x
LGm84ZRy4/RrHXr7VoscIlt0YxYZPf8lr3fsV4B8i70ITm4WB6IJjVbetooWbIju
WC9wOKIIINOtZk9P71ne8FJcvy30R4qdaOb/pRTdfP3/W4zYZnw/LdKT+H2PFSJy
SEn2f+4XjedEetnDaxY1bnHJvlsWLq2kIbn7hJskcqYMQnSZsANQh15juGO9eVSB
1ftnKY8sp5WIUOeJA1zxY3z4zozDI+hz2R/RHZ7az+LGrAmKXxTIuyeFdazYvBRW
hLn+VxY0hjcyHsp0P4yBrdykkLskKIxZnEYtek7c9M9A8JnanAs1SIbVX1oTvpvR
5tZ0GLTOchhdvU+IebYw3AbbsrxegmNFe0doeq+omhn/EoX6BufaHsyIheF5NJU+
HaAvtQXgxn2o63m7FO9wcbfAuIv0AbEtFJYTD9/dwIxgoJds8GxJYPUXSZ0rt+cs
uERSUOJXRWbiOe5T4ChjdZvzaikyrL3oBB71W4oVwwAca3O3bYchrH5vPc99XwRN
xucyQPtGy4J0PW4+8LJaXEqGfaTX3zo49l6MM+LRMZfmTVdpQlOOKIp6j+/7ay3Z
m55KbssjgE6TQvgrwvwkpdm3tiAAAKUHVi5KRV195/d96xtc/C0UqtZE8rRaPy8R
lhZ5x+N0e2np96i3mUpv4yKwFJNEJSs//RgspW2RVXiefrQV1apXLr+OYFUsA5Wm
EP9GhfpV/nSy1BIKIpO0zj4W4ug2qFsC5BKVyh0x+IuPLI3n4Bs3Z/uFa7YQGL46
4OiPhG9dzJNR1cP2XHTioBTS2QbzU59RNnYtxJS7QPLaXCWKHoH9H5wC5uzyo56Y
IFLQnJFWSv4ZCy90rYRfaYa/ODWDcVCBTCZgXZZRG8ljq+cr9ezEl1zgXrkXWl9m
vSyb5518O2JzlGQ+2C7N+AeWucHDZUbyjujgielB5RHzT5gU1Gyle2l5GzoqoT/x
Xbapf6APPE/2PVZIRTnlsSG7HY4GMg2W2yX1/a07gYZEjnRRguvrfZ+OvpSzQcg9
P7uLkKwCc75NBZlXg+I1e0Kcas2e4nR8AuvykeTlcbQBzv1YENB//4Rn6a/pu40/
u8PCS0DczVPd7hXnIeYbBLtyZEDAhcWpCyZmjdWS0hxCABvmj3PJfHjpmp0GP7hk
L5CJG/vMLcM3oR3hR9ZsFeRJrNxT0s+7FtrnPTfuW8lypb/3bbdml9btl6inHNai
I7r/4gXVCXbHq8htLTIIyXk64iP+9XbpKSH9IzfWfrQZSXp976I2DZ6VWajsHJQO
TCfQCgiB/ux1LesSVm15e3tq6aty2Qrd+s3CfdCcUXYUyDN8u/Jto8IMlOzNgH19
OON3FL2raNKkJmeGivjozRe0BZSvtEAJifwV2tZPNFHk2/j2nfRMXK41WHfOnMOk
uuOdzJOJwsrlI6EF/PvyupmBOetNEy77xl93k7tF7fUm1LqxPiaF4YMHcn7MvKK+
UEdRzQDUOVOjCyimbV+x67ibEetoxZU6LZjvbsUlowhPhT8l2MYrtU0sU83+sZh5
U3rc+bZnaR6Mx+BsQ3/r6//G8Yob47ZUj99NNLYAErGzd3qkg/Nk16kn8xEb9VgI
cp/x8327+LjyjXtLCXWk4TuILp3d2/radduCNAy/Q4DFbWpDDTatBT8p4pfQ4Fzk
w3a6xciJQ0ezeVExzdeNBbQqOWytnlcfAnr6FzrmkpYMNvvnLSIGOSCZiIAgNIS7
Tx79J31H4TO4D6K2omq9O5FL9I0iqcM6i9GU5J4H/zbNE2o15MdySm1My1Ygiy6j
nYgdhxcCPB6KHaRhbRIMXN5NSKZqF2rk5LEikCRkQux7+1yzM+Pvk7g5c3V+QRlP
oOKWWKeHEBivOhfaxQbB2F7ytuqqBKlt/UepkaAcbT231epFdM+4mriwRBWT3GxQ
u84DLJYI5mYTO+dtMiGAL46jID5Ji7r4X3o12I5Jap7/fDj8Rwayn2Fjrvynm893
WsjKwvixNM35gES1c+sg+FjqR6B2YCzxGvBpWXW6EwhzaM/o4bMmBjfO9b6XBgQS
ZZnVLbNl/vtMdA+X7lETQQKYMmjbPOfWP0IhqIbKbnLJZGyxNeLjptGQr9AHcgEv
P1LLcscnpdzO923ztjMyBb1pxcL3VA5P4To7RHRSsSHIzGhMo3HSKyD5ca1fpw7H
3yuwRDBLVvPJjkXknr6PZw2ZTpn/cL7Z2MRG3hLtMms8yMKGjopFZacvN135CPoT
h4EBXToyCHN+2SV+tuYMD6XiCR6jn2k851L5cpTSY+FPNN29HmH9sYTtMYRklF5r
FC8KFBXsIBZ31684rfFKiiEQfUXdHkI3XX3wmtE9HOquHLeK8RfltmQOBuOx/o71
SfuKHoiBfpW1AoBKl4oVTQmRFrmdFIeRuQId9iKwNMb5cFUVY/NtaaQHGNUcUxO3
fS3NXWmzS6HENbD/6YLhhdisasCBsikKM/RSelMRZ1NQABzraWm28gUVrTdgZ7fp
ebveORoawlX6LdUjwKYqEBYAw6vsIyz+4qlnreo4GM80GGIc19YlIuP4DRy/lagM
VpSwHEb43Ty4DYbc3lpxLBwbvTsX0HC46Q8ETlb4qU2oy12zkqf1ucbw8t7tQht7
8yk7xXFwp7UXw2IC/AMnjXV/7PDniQChbYsDcsAjQBM67CZ7q0le3ShGZo27u62B
eCNGrRAPeOcWzW4kg4V1Vbajn/haM5qM6Yj3Irwe3BghJoWzKv/zTK5+ZVWtmudJ
L03vB3PJmsyYhSnJvxzFGGHCvSXDR2dQwwuonF5fJKyx6hJvbCwoj1FuMIfNqTHh
Ila/TVsgnPt0TPKaFofYkRfNHp8WTzkFpVtNAMzEWUlC8vspX5iNao1wHn0oVrLc
1oKs6XpZ9uylUhiZH7ojROTwuLtGUHM+1xkkGB4WiG0IqKq0oqQ41WlXJTwmGA6D
//GS6O3B9DsgTpSf3946mOee7EQigCnYC7zF2j/CZCo74/Clwo4AxS+ByIwJI8Zl
4Qr0L/i4Sus6ylGEYC8m/qTHRdgzNU5Te7d9Rmm0nSQf5c/W8Re/LsGXyYgP8d7h
jRhA9tJgT7cwB2RI4VVCilJy3P4y5c604PpPGIchVPq0EPE1rqlUHYfMlDrKRAMs
BRFmj95t6O+ARanbx0/8SgfPb/PIwowmJOtXG0zLURE2kgYuWdpQzILO8+uya3tl
xA43Irsyg1/afOMwUgqbzN8sGeaqemwzZHZ3r/dMt7CXBSiUo7JsD8hUCraYtJ+j
aHbZpG8vrzzMz8fSFJjUqU4e+vjIAJfo/SDXoNC4zcSvZ2WRGZss/jmLZNOLzUHE
BCC8L1o4pxr+p8nkj5T7TdnKWbjO6Wg+W9elu2x3r7NhX2U1YLAMD/EeVMmO2VrV
ONXzzcckS+8ewMlYlWiOKQetO7Sk/spiqBcELzOThI0Vx9F3pHbZ7v1iCojOjd2S
hLivIgVc7KlzxgEnihFFnJqrW2mC6vICTLCWpk649SUsjQPc5SR5enaYfvOp25ga
EQuo2ziM2TuytNlMpGymA+3o2qNs1yfRQRSsmJCaIqWCmcvJVe1lTzhnttPu3R+5
w1JL2fqcs56Gz5OKFhpu+F/ccPGD3qBIcEzfOjCFqdmsYvv2FbgBzWy4UKewcYcK
xUAM2iZs7eV9hcqgiyVPBFl/ayreiua4vYCVVdu+D3H11rW3odbdk3is7IFpINZG
M6sCQS2+LlTRBzwvuFN2vNeis+rJF0L0oRxnRDLteDvuIvP6jMpRkA47vv7wEjWu
FvkjZ6VR4QM7QH8S7E985KrZ5fTxTTeE68IpN+0LwCivOLM+Iaajp8wgYdNJnQ3d
t3hwxr87/3pd5F8R1Lrs4KM4+10IAjuX9MR0CeGrizIxVRWXd9mnBTVlBBB3qkef
Kr+HAG/j2BLPtEy2xJbnkzGqCoYkw40DKsOpfXcBk9OfVHg5GVTkjcWM/+aSBDuI
0JRBED5K/XJ03hvAiYgw6IgZUqjAWJbp2wjOJdtEPgzj3LiEgNyGsYVF3HwQW9qZ
4xm3rvOGU0ZB+TnFV3cCLNNsa5GDFKDXYxk0jpYliufpcwEykkI5PGPjo3A90mLZ
BmtnU7T1wunY4lwRVDZ5TkBkqRWX1v0JmHF+cO8ZPm5RsZyBv4Asdk99zcAZglGq
sFPmpyP6oFF/LcgQsndhMlBcXHF/sx0IW3VBcDya1ouhHsdii9y1BwrHOFItk9jz
nC9CevRa8hy3Apgo9W/wdR3AvThdJQRLN0UBwkX9eIpqJmZ6/OlMlol95v+5/CqR
stpsrN+CDvfbAmeOq0AhZ1ZSabh84+mZxx6kDrJSRGci6J4CdugcUV799TqUGbHi
+n19ioMzV7vwdQ/dgBgeSttfv32RXQm8rpoK2m5kWaNKn6Tg8bOHDBylzUC9DUvO
D/a80Kj3V31BOCW3tXFhjUdRuGuLu9t4X0/LprD39dp2JRIKxuN3lAWiHHWQ29BO
F+H2rq1Dat4C0XZ99bmlgDVpDAeMXxsC5wbcwoqO6VABUqgW4zKvMGyWUMSDvl94
qPnvGSX2cmh+538jJdz9IJN+q8HmUq5bPQ5AROh7vA7RorzsJCMT+1ZuusAYdQBm
QazWL9KAUAlYX2kr4n4CVzFQogy/z5Ci15SC+l0ZST7qx39uZdM8obOEvB+SfNhm
dvFfxCxbPCEibb04Qu+Ep/PXtqWIKZu8R7ihLacwinnbvcF9HJQ08NyHkICC2FU/
knnzOorOAga3AD/NlBY4fCy6zdK5l9xNm3OwMny2SxgegsnGB/B4zFA8xhV/yIXq
O/NELvJtY8oe12mk+i9NpSZvSZDTsyqsY0e7J+ADOo3325SSDdF22j2CTLuFKwoL
RJjdpHqdlPCByecjUF1qhXMai7ior2joZrJEThnlJ5mzjE+Ri+WQaiLMd75m7/OK
QEQsL67lmB0k4dFLOkPVwyFEu5g0sOPiI5DT//j/PZWUB9W2Hlcz86dtAxfUZIm4
0/z6w/eYRuH9qF6htuSSxP30h6Yf5JrqGVD1q9F/71EYHk4d+Fozg46mI+8l/Qp3
lFHYai6PAunqfrITgvdKEVjsLRTPqZsMiF+PCTvMu4HxiKm5qdNat7auZZjo519B
t3n7uIJrBlz1es29jLg5eJ8xF35yD35M5kede5udpSnw2T7t/0OmX4uoxKsGZcq4
TfOSU2M9BoxuQFlK6ggK2SRvYwFNihMAqEv+NZphyrkilsdhwqUyfJ+DlSkR0oBo
VzpH/2nNNCzh2XmcuEJsj/udh0SusHG0fbMmfkUAN1z/ewnMAyit/+WtBlQAvAgg
phTgvJr3GYFRwFAWy9JUl+gAzJi9L0NPPWGOqYjnieuS87kEmUhwNkvq1FZbO5oS
weJ0Hk9uXoQaccpSTZFKxTtio12hONI9E9qbR8nQcSFrp6VTImVVOxi513YUOArE
dvDrGwD52l6JLWBFyFPrAAoBmlHmJo2v/03hJir1vi3OVQ2f6EhVGYdnn808Ki75
amOZ9k1FBZ3866sax62PyA0aCWZcOcE4sFawBa2qPJzNbam2jg423W1Cge71C2as
C04Ug4v5yW64BO03xaHCtYqWlMjsiiA/84Xm0aIVjVtlRQNQCOv30Ychs8KrORi2
qUYY1anhmlDnLDGLHjY1CdYu5b8w2/3/xevcr8djc2ZoOrFzM3xpnc+RjwZd/voA
Pkx+5pEQ2ipXLfebRGkofH+XgY0TDwUReWYa+2mKSha84snb5O7ljm5NqZc62Das
nLlgQ/Ww1PSWiA3Q+Iub68eXe3XaBcxY4UJudwWjKismy0gg9+6L8DG61LzwQjh7
vXdakXgNxNLRRjMjOv7EQEOjnVyF0DLHEsmMeBajWuDHUfb6zgDLy2exBhatO3do
db5t0ppuMTR9kBRmlpUYZZ39TGPL8Ng8+WFE55e5K6DzDWZaVhKm5Z4WN0xvxVbg
Dr/yV0Yd0E4gS4QE3eCr20mbDyC1BCQ8fBHQXBwEqTvSnyAcAlPZBKWoy6/MkVR+
PwAy1yBIgohWu+9b1SHNc+yVkNfOmeP/j+SkEd6lDzv8UY+TSj1lq4GWOFKKg9VC
CDNiO1kmyob6TXr22Cr8RhcuB2D8D3HHjp3Uky+ZCjPtJ+CuFpDEs+WxpQnw3Muz
mH2eraiQmTH+Je2XW95U0QTbwrT9CUlFwnetVv15nPRMfOaBO82U7L1bdyViaANm
6pl+Iozxe9MjI88z7wE8e3S+GcSkYYPg3741G7cpbCwDf9eFSoxx+KEpCHrbo7Yq
r7nbjWav2GpTN7hPmPToFnMoYMz87lT4OUpV+TC6nTTVNrsiddIOKA6T9cAbQkJP
tCcN4zrjUiScNeT4dJwLjOkKHzFwsx3UtUdaV7kt5lhaSA8LwSUEweg15VK2l9Hx
nNd/DwpV7UmUJ1NNNbp0EoC1Lk6ZJXdbjqdvWbTTBHqdHu7r8EfumqyuefLoJl+1
CQ+e/Z9OwcsuSF8lZ765ln1lKjz5oeuGeMKSlmuOFG2b/VEN0+0WJkHQEcL/xfDd
UgU6XA5daBAk4vcAocm8ogpo/vCYCFYLu5rmB4CJyMRQmkFAxAmiCdcs20S4RixS
Do/5V5GUuGapGu5rLfPkL4B8+aDnZdifPaMN2FTWtD1pW913nz2cl+ovaIYspR92
tnlTtpmG++ESrPFetDXsk1xxki+mqODHZZdAyYSJOtAlyKNoDnZNLugimZereyJp
i4wdtIquOZZQHvfNueLCN3Te5wPPZkxuMVhPH5FfueDN/5JOIUK7xpRD+TYivfOT
Pd8+Kgy872MyNjZEY7mnNWBPZjPN8e9sj0yIhmLFu8KxyWyUI/6vi7xheOh7Q2LZ
3oWDfZCy6C+OjZgfzOcesTR/0DBsxyHUXT64OM05Rh9hBvdvrt+Z+URP8MTnkcwf
lnRChfTF54OR36bZxpKhgzDA0tiUXMEbCaCy9VtKW3c2LyJkwZ0mFNI+ADaR4nci
Qsofv7rzXm1vlKne3S55Xp1JHxxFkactpRl4gT56J9iEu2Vvm8SAWD+nXO3Ijt34
2yrbUryEmuAuf6g+WbiAWjMz1OC+kRmjIyJZjIXeDY8vxeAwI/4GgE1o7P8hz0be
XqZ5Z318DEbLb9vRRNuzTEOHZB1vwOOt6YNLew1BDjoz71uZd03cQ4bW6mNiUyKj
h41EM2Ix4nRBpziZRu5kyzohpGng+3sCM6UH5+VfFFe6OUVocqLfysUhKFq9HiKa
VKJbk8ibEyY4vvetM3I4C7B7g24hoQdORuokyUlYTBlGSZNe9Uatb2nMeSt2CTbG
n4yth3r4RLxUSn7oW8pPS4Hl4fcJ9pSxszvyDbj8zVHuiGYK373G+4JhOKqiuaPc
L9t5megX+C+3wiILGg0wQbs4sfSQmwn0FUhaknt601SH8Rxmv6c7C8GxrF7zGQwq
pOn3rJNdmnUjGzW05rukzkzzfMtE4L/ThSHXKxPatthBmQht+URwvtI5FxrY5rQr
HEpALEG6NthQo5bAxBT8bRi63ADJRkZNfBYyGwv8FFTPCkr+l06eXz6xJDQskuIW
zPuj+K9lcjBfZG2jnaoK7PVP3VIX92PE9ct6dVFdRvVKPLJls79AOheJN6CEbxYP
WKmRfcX7lcgII+nGA16zuZV8GXNZmbMQ4MmNyOIQp7hZk9axwkriR2t1/7VUEqoH
/ufuFFkC77iuEZF4RqOePu6Z16zYY5ebpmCck0ZQDKEYeVLcz8JDDGISQBHraZ92
LdgGMM53kdF5aTZsoaF7b2PV2goqZuAHPrV5U0B9uzMTaPpaEYI0F+3gFcNx9con
KAWJcs902UYsWx5ZZ1IKJ+0fCFGOyYTWnXhUrWx5+Ba0lsc25XXfLZh2KgZr0i7F
2Vb4M9bjoj81Dxt7+0TbYix/Mmx7J8qASx3W/GhBXeJ3/wu6uAs4sYOcItCG3HxG
n4Q9M6Nqtqdyf0d0Nb4DyVN46JQVX4aL5WqWnEg9Xe1LJiMOa39RGVeQDur6ck8P
5K5qaKsGpzwSN5Te3gp7tf8Fzk4Gwq7i86CdQlj1AQxVBkmj8eJwCSFMH5SpTbcF
tW3QlgkpyXQDk7nTZvzXlNpR4VnX6egVWiN5adLZf+KM7LNGRdsuRui0emo/t8wH
nSDfbwKM+BNjZkSq0Hd8vZFS5pBA5pPYlTja0+V4OrtMDjYByhM8D2q77jYKTGN3
1Erhrr/uduwlVNuhvFvqWG9QH7IQIexApLIti4efLwcQIM15wuRuSEYW8aQw5kOu
AefWXe0XajniIoaWh3i5luCjihE7EG1/nO9pAXh0DaXZX91zPkHEHO3YbMguNvSi
c2ntZCoZ0GE6ZUNHAg6DajROt6pGfYGFmNLumS2oS1Bw/fBFunmVQSQCYJ5tsf85
eGLeK/UHUn/Oe2LC05Fe4DheW0YdS67mtdo3uxiML3OB80155h7uiTefGhOvkk5X
sxsL9cw9Ryo0tO/h6ys29frqKsNGofmJQocFsqjdbl3HBIQPHzuoCmYAgoBDabW/
fdq3U/s8i4MczkyJJR9rhEvJiaL22HbptYhgvhFC+qWRlTi2/n4zToaVLE8rTFq5
W6aguMrF13PNG+2pCinAgLhpbN1ofDqx7+IUDi1imns4d4biOidfsGqaC4rGZF+a
m/0CoH4AOpFBsImsvmFjBgPrLuAIQW6EE1bgo1C3PV23Qdyd9iDJ5nVewlXrkPhP
hbg8jydiUd5xFIQfyMTJMWO2hHxOY01nNMGKufXL0ViVvi8BQR77pckJho+X67pS
jZcDH4n4xFgAhhBArgXb+3AV9c9O7GkEwYVoMY8F8uvUuwc7GPIikZul2ytmMnZl
z+K+szVMR4awpliD3K2z581LBSNoGhhSJ0LzWEueolIQWpdtuvkXMrPiCl6Awlms
vC783ADCOqGU4DXRmo6KRjEGNHZ31qPNOLgFr03EKQWtKnqUbEhtivJWdPAl2YgX
tjmjMTJaP5qjuYoDogNuDJjdFaps0SLy5l+oMJEk/eTq0HClRI24lcg76uxcunON
NMC2BypWXDU6XgsOII7CPV90ZqUvcKPUOuZGOKyuTOvZryjjRZKbatUZdK1/drOm
L19l9EK3jRvZwhWELCTNSgmynrFWIVzIzvXqrvefK47xpjN2JyLb3EA75V2r9Yt8
lyICiFRjLSGJzddPNlnA1S13Ipbhp6a4M/u/V75abWIb5R/xbijto17XG0jbHta+
iaDj8oZApUgr+Y73S0WjHw7OsvZezyk4pw9kxiciysqVHdL+uCFUufeEgelZQy8O
So01aJJRYX5xipY/XuE/4w11ksFk+2bNG38CWBsGLbrXijXIgL+SHqN/r8pfra1K
baHRqnQjv7rVHSYleb+GsgP5TiGP7mEQJHsnEDy1DQ/ht5z4dk6iatYZQCkW/il1
zNP7c7oEJ2EkCFRUD1XHW6cjTWEoH4BEmrHLI6SYTmG4q/z5r2xMknTmMioMCDko
zV+fRRtLrM/rgXKsF6lNckJowtQjWmYLNUTvV6ugWHKUNvQXDGTjP/el3M81uY+P
8wl3IL54awiHo766n7Wl9bo8IOpgYtIb1AkSauRwXw6lMyNyqBtGo9N8uaBKn8ms
h5bYUqbJzUjHRf8ELen6EdlVpEuytLkTl7o+JUFeQyZ3xuL++95mlYJAJb6FA/I7
4ezmAapYhjhMa6KitwOJ4Dooo0TWjigaGGRz+YdTUsqanPKb9g86laW3oLS4VNRk
RCnLCbJqQJl/0hEAcAH+YF6PobYLjlgo6ruS6L/W8MUeY8r4IunehZAja/HFkNmD
hxJALHA+B6fJP2LRNgnmwIPPgbRCBGadoZazlTDxmapY7yLXBN1V7VZFxSvrvkVu
lJSiuneyNKQqSgfXZ3P56gjQhwDkBfYqOcQICw7sZUTiHMtMQMZ5lEKvvLBE09YR
2aOKZSEVbxK1IrH7Eiz+EOOdOAPF9ZLBPpulAPTjQyCkI1gQvdNwyz5HxsilTkID
zFk939/wMTQkgOzzEgSbjpRuHyaF3pVF8TqxfUsCB5+VDHLpxgm1rwTjKSyxGb+g
Bno9OYx0NuShmIgWplquMcLVBQcYMbl1GgBn6B2Wc7q7QGZXx5/quxOTfddFxNJI
O3YvZq9UNTFmy6yuDumbacDE6vhSXZDKdtgfQKX5g7CiBbveNbUzxysRD2zfTBWn
DtBlvanHzl5ZClaU7J57WZ0GtjXqE58qqZgN6zvDRys1Jy7H9EH+cMSdRigGRBxO
TD0bpkwtMzjhiMICwOTfcOoTPHJvfzQl/iEmmJBAchavLTdjZ6gqJlA/QVc67pPa
lAYE+0g1erTyL05JMHgPhFmeEDa+Su96hLauHTA3aW1Vpx6TSkc9jWmiBWV3bTbu
c5BnVgrEXUDeT/bcE3fMzumlqP+LDmNvCdfJ7GuugHT9oJ7WKiF9rw9g4wxDxoBO
uS/M+3z/5PqoFGiQHY830V7KewEZUVC6zmX8WEy1xjwXA4hFtDYlDiHhBiFhHf0x
f/MFoSz9ljQNigpDlvG1SxzTh64Nww9RSPKy+scDI9J/+DrDVYj3d8AKks/k/HEM
aoyf7g2pRMc+JCult8FCg9k1EpdgWtvi3cSIfVsu1gd//0UouH/YB2y/9w8xGBVA
BDp3iNApeCtl53s6E4DvzZ5TTpde6RKuuyXyPmIfbkHDo+BObvzK3dDZu/Cjs60q
S4Y0GjzabKSTd3V8xE6Je9Sku4GgDKyoAu2ODIWJrB5m5xE9ikByMJtqxeWbi9yB
JXUjeuUJU4VwJYxgr3OCNmIPs8OLkE59FP5sYvEPGhOF+YhVhAZ9IiqXWfBKWB7F
nOUdYBpsuUiYlmD0wSRjW1qi8k83f+AeoeWG8lbdlq87IVIuF8Oy1ucZgkAiPWvq
x2eFPnfInSn7UNPxcz9TSty/ZLQsEyapyED2rS1eMKVueNH5D86l5lPbdZ40unym
jMsBpFjPqH3sL+Y/OmF64Dwg6iUayYIr2C0/pyVRirSp16zOoD5Ee0xFsi34r1T4
tOwRS+6zQS3CaKdEqfMXzy8d1pDOnsaSMWIkY1jIywugFmtOD8lv0fQyRVKR5aYP
+UqEzU/hyAHW71qGKSBP+2VMPtbrysdiPjgFhDAsOMjIfqC4Fp5GO/yJ2BNnvWUH
IKYzbUnX8/C9FmIlCGgnOqrBFSoF8W66WZHXad1A8yL7czqKoR8ganRnddFg5TW0
Bmm0AtgJR6e4bBcqJON5Qgeh7as0gGpCRedK1DU8/edlxhCFp4k6QhTuZBtqUXtB
WO5B9JTPBaKlDf6jhYvVM0JPl7a528I74QTnLXwOsfhGouzqSzL695KH2gpJRFxu
fSrNgW9or++e3VrMg2qIuco97WtaDCejSCiAvPX5wsjwnApwAfE3flzHMc/+ZJI3
oFYh7Qgcns4AN+wz7S7iOly0SStW+E5I8xsB4/XNfGWRi3WnD7caQ5/Wge1VnODt
dDm3wpeH1VHtqUeonxw/Oyj0zCnyoEcRrFoXt3Znq1HiGIsdFcU8bse5DbNPreG0
KgZAZyKNC1snFcCbHnE8rlyaaPPlWayFcF6BtswGgxDLU+Q9MNlc0Yf6HdCOx2NM
AN3p71SvJdvPWRl2OhwA8ycnLUP/6LYjxQXUKklXnS5KHBtJVrWaySQ7MFulMlH2
68mb97HSUnym3EB+UD/ReFgxcP5xOy7A1Z4qF0KUFTI4ZpquqdVcFx321jgZ+ZZ4
0LlwtS1mmfj1qSmcMR8ta7+PUMCrNZNa9KlwGKiLuu6LLoTRRX/AZ/4bJV8jecLn
RPTSz3TAxRAnfoPP7TUDN7GA3DKqLwlxEAntdPUKK2UAcojSeGsjJtxuorK+OVTa
RUcU/RxUKFgCEgqXEzsn/xGyPL8zoa2Aw/i2K3NRgaeob7H/vl22hq8ga6Tkpre4
HBUPYK9duESxCLYv72M3cE6tlAPZovnJ95eAGCfC27yPI921DKzEekzHPmvHh/ZA
Z886wUFufNGR6jaC2ZhcyRymAxct4J7bTRVa1C1G2fHSo5LMR84EpatDxjxeDb0Q
tz6wdQ7AfcOf+4RKx3OCWLH5547xIkBkHolpPSGbcDMEWERo0IU5tU0Ld0TXU3u/
Jm2GezoLKPzs94xZ8llbp+Jb9lX29iKTXQzieUf2rymJ81mTsoL89m5ZiHXtYET5
u/cQSBL7JpXmyFGqkJy1SiwYdZL2ft+qU95GLnwbCINTxddGF2r/asl7dtcDsndL
SI9lz3loUB8gPCPM+89HMJcjtYN2a/vDy+xQGHxjychmi7lPvkP4PresexJGNJrB
grETyEl50lxA1/8nLG1EuAlnOBzBGarK+W/KguZd6dJeTxfIZ7et/0zAVsdzaIsY
xvc252zB10Krs0X/A1ikoEmwu8hfaVc+sckKquWbYAG4QgFhLq7vszPJNaNkt42K
tJYuoeMERVSo2+wTps73oyKkiE+4escL0Qq48C2gtnZPI8q9i58rHfk00H0QuK1C
xwsw+qnxIa5URFoEj7+rlSmwImCk2Wk+X3/U739tgHJ8DWgk7zuTa7R1rrko+1s2
DPP5rdu8Xv4bT4C8xzzlJR9gg2E7qFi3LLhJ+ymrnWMLVhTgkbn76PFXR3xAJKg5
G6NaPoKMY6q862m/SPUVbFc624RSuFIoQThWRzVbLJlWS34RdqgpbiMGOjfg7ec3
6wcvO2VRjwiWKvfJKF80n7wK7BXfsOn/E66U25ONSdqrrw275YuMTQ2b5+uzTNQs
IvnQWrJP3iVWQOhq636Ae1eM8EmBjm7gjtgr0iUqyMpI9uYUTwQFOOYQ69PzJjei
+8e/Aa0AnLRvCkJaTmsNrQEDVr4cIJeL2WLIx6duR83+SQLYFm0YxM43HZxkxu38
+LHCaMuyUZH/fqmTKgrFQpH4BrpzyAxHi27jMwYTes9VmUEQGjkXxS1MJYs/NQah
N8wFwPwJWSOcvrTWlbFTW3Wu4QeoUQWveZMcuX3IMKZHMFjyIJTkuQvaWRz0+w0B
CvSxu3up4UwcbWS5HmXuh28joNyfc28Z2juRapslB6/8x/qJypr1nXwr5W6DSQ0m
rg+BvxE+2H2O14KgSeb+yE34nIjrjaTQyQ3vliUgTgD7ThJEFb+GNQMBqkv8+jO+
Oik8heZR3w20HvqauKeYEXTGJI+RkGqxgY1f+NfPNjm1XWVkTnwadf17KWE0XyFj
v3TFaVnFGgeEn96PSU4bkAgrXva91DmwLS1op89RYzQd7j6r6QGyQu+hc0RQcQHy
1wh/w28dYSkF1sullkm3NpxvNEpOMUDw16nrFtJe52uqvk6z0jxyE71fI1BXb0Bl
H1AYJG1/ukVbpEmJ2e3XamBRNGN98XkfSqNJ+bP9VmeaVTdKzUZkXcQnzv8VSamd
CU6adAOPACGvOplY6T5fMVJbpSnaeqe+NEKVutWgGFAxQga1lUMUbpRjhfCNgS4/
Q+2LHqAVLDgWroLMD/bQDxtlpRxpNnVgSQ50RcwB9UMsbQzmprheoquv+3iu4Jiq
TdelupeRnLBd6yDUQK3kdd+E6efuX1CFZMiTQmwOIwM09uvA09NUVMU2oqwfXKBv
/aBur5UFluZRX5Hgxakv0T0jfxKtlb87PJKrs4Pe9FjFtL9iHAKeqsNfxNAr0NbA
jReO31FyTXS9Et0VJJKdvD3CYvj0TlTvownBWmR1VqCMINQG2RVlu0B5+5JTkCNt
MWAQcnLr3xZzTQL+ws3WSO5OxUUcTBwLGy4ZMxE9d/9DAlyQ+oYloFU45lYwAnD4
hmQ4QVm789fyofR8TnrrDEWDdPxB6K6Ida5E7vmjInscxPETvSYS5T45w+DYovPX
8R9IrLjOTUUjw9EVwDV33vk1TZACvmKD2jaK6G6fFl2H1OJRTdn1y0yLQKYtBLsD
9zWX1IZHzi1GgRuTdF1DIpZjepuMy0oXmiedxibMTgv3fYlkn3qAdzQI0Lcn4GOc
4yJYI3CCvSl7df9rFTSfH/EgF3XeTPvtpHANLOrW2HojKv+y1GWxi7bGE/n4acTZ
EbmaIZ0xttTK6pJ/Ms1PrE5pAXlaAO52OGv68wJacdTWSsWdHGm8QmF5XH+FBD9L
m3NPtENzFlMqAnwjsUhrHsMYlqavI/rtwfBXrYVhMK/uCsF+JzLrVcWekZ0mefvH
2+3bfkokZdFlSFVH0MaHQuFSKaWoJgTVkEL/rMthtdqtMjYGDXDhw7954Id7JOOw
ClTKEOM6dSXZ5+zZ67GCw2W40Kf1/Df9ZrAGdBbiqyL8MUKTCBtKKuvTdTEGjngF
ItFO0f0TbZrFoWZWkw51gY8ludN4eZf5CjtyOkoM8lOUQhwSaEnq7ysPLzWNF5EC
FfMRCqKTCHLxN+aAEadUkIeQWoWMe0deEhB5vRKShsB2r0b0AZjCTBLeEoqinTpj
oGh3iwvnr1GXfeOUwJPUxK9CqKfzpEm25O5eUyoFtMuOy/BkGzXNv42l8RQ4SV6S
n5QxrMxnmOzkfwPGGYLRfsUVEcl/JYU1BTpgaxwVM4bOoZXp1IQRdYKittJoVowz
y+3F+HE6XdD8qTnQ+KgOkSZ7Hs6MadQBbtm8K+fzF2qGGEd1jB2tCFDNzeSdgnks
OW2PmUI2mZ1OnJvHlXZK99MjApwANMPu/Y/L4Vw3dQpTMV3abjVZ862WiXsy0zpq
WvuqbWGNXT/zsO2DE+/W7mFAZvFnDf9gYFK9GgTlUOzum07M8Z6vhweHhICa9txO
8xlwhMG8324QxrxcPBHLijE49HxdviBMGRfjvF77azIYJ3w5OktXkf5xn9y7so6y
QVbQQROxSgVhzA3zwk8UfTmutGU/iYEutb8Hkp9y7ihaviXo5CSjsv36CVUZTxYv
4ODrB+fb7Sej59+NU163bxB9OMmYUuhQ9316LpbeBKsDk77rdkOMdEMax8WU9Xnk
fvx3xyfjAq5n7u5zhn92bGWIrB/ByKMRVOP+JErSl3v58kKkcqNm9z7dbPDa6JLL
YwBKtp4bKyBdnwdpmkgaN206T3D7geXHGczIYG9EXS0bXbON9CE9TvU+78ocvIK4
SHvcqcToyt089fEL8XfGmpFxfErRhaX1gG+p16+/Q0M6H4AkM3Nc7fzcxHY/iqBX
WbAXyll0cus9lftDjgrPa/dUMCNGN1OLMrDy6T1hAbv5AlLqGaO86ACSxUJTneTu
T0RFIVNBZPH53Wijxn1HOj8a9HxOpECWWalqKdnX0vl9aLQfwTSSULDyIt1HkGhq
8mnipI54w8e7BTmtgG2/925gBZvbe6p8nclt3obwxT9QykmLaKR/GlmPYJfxKj1b
1imfouBJH1PfVbrHM186Fz4S0vs9yqbmfc86sEDSSIYSnMoWxck5bbQe9Saw0wiL
K6ZLQKYw8zveOEBAXPjpybowlP9sLcyiCBMAdC5bD0Wc9ILWJkg8yDrtxdQgfDF6
AsfJhwW8vz94vOzHO+GTzGsgGtvm+JHuENpZMrakqIqzNXPKtdTSiJ0uUxB64r0k
v9Iya4hd9XlYSKB3OsK9DkFgAY/By6HxYxse2gWE+1BgoIkgEMyXLKv8IBY2fBga
3E25kj7qrzmHo/IhEhb6c5H25+CxCIyhL1V/TA3tMRX+bm2IC6bD+bwqlKxSvCWb
kB+6SVpP2JGC3e1YCd572woapLHYOze3InpRCCGwDcRHIr+rA8e7l6x5LgisEscO
EsSxlV0Iauyxo3ZdVK/DyabWW0YasssU2h+FvxHyKj/6lUM16bPVJFATU7S8XeGs
aFHq2xMO6QQN38CI25sJPYIb2JLgHgEh9m1CmOZEm1MEYj2uAeyaKOfONdnWKsjQ
YMTB37UAvg+zc6iAc+WLH7itcpJzHModFppvXqq/O572p7lJ5pOvfFIasX+iGlkA
r/E7rrl74raKntEZD18TANbsrohzZrGjjJ8jeiVWJYf2XHqxjnqPetrzhQVRSl20
XNydebudp/OE/cuSzn82U1FCA1Pm6KogOGTUOQfCm1MBDKy7aDVnFAMhk6ZGNKe+
gNZTRXK50T1Mrs3i8E8IAtlLGcVN59uXv8x5fAi3b1VcKcdaOgNIGd8R7U1b6t+h
HZC30QEkHjLknBVY6XpHJeVeTN5OAwyqRBpPOcwaDBy8BBj6Fp7axLG55Cm1V4uU
mPE0VubXJiaTmBCH8pbuPW1GXnBgBmds+DOuSgoVWjNgyC87AOE+xNBzGRuIBS03
vyNnghmFxln7CaZfZap+x+TGl2noaeYGs93/KaRlco/G2QkHK/SRh+q/F1uK9u+I
TTa1LLiGIBrOR3JPW3WvPg89LDK4yf+Thkajgf7G/TaHY/8QP4cqysQVnyqSElBp
gz/vul+BP3mEIkIlRUO09HYuA6FPwoooYeB8O+CrTciEa5JcKP5sDKu3BNK4FT9g
nB1I0DX4YTOB0NtUgROJVoNzlx6/rYv/vcT4a4OrHQkV4xyzGO5t7AFjY2LNF112
GXthrm102w5GoLXKo8dAuLy//ijhWIZ628zQzpndiyNh6H/PRX5rFGh2X/pKtFAP
mMeXDqh9D9oNwpX0W+ULpJjWhahJ7Vt+lFRudLotmBWCrztOQmu+ljQ9RFa8g6oy
ELIhuMrsTXF9HbeE0ORsyX4lc0aTLkfxJeXA0HCCD/2LDVodtI45kABp9i50Wdo9
DZF8/PUSrZg17RRSRa5+INshXhtaZsRo7nUeGMsKmEwkH5u/Rsy57yC5fA/1UN/3
V0MH5mfAZYDq4cOK8xG5M9SFFAVwh8IGQFQpfszTnlKUvm77+xkpDdwdbA3e3P9F
rk7m8OhrOqcbwPF9XUuY0GZnEx7+X1PpwngXNwffhsjYOvHlJvL866rSR8XsICwt
CUi+b8Bjnq9G3ckke8GeqCRfMQQMMiFP8/zTaOEJ1R2IE4O4/fvef0m1sdMH/xar
gBGMrtZs/SElH6aEpT6RF9ZEv+FxoNryJCRgui+NFV7i1MDo7q6a/FdFU1LaYaI/
TwW2HWZPFm+fXesXeOTepAYvyGTWUfwB5GW78dTAxEikurTXGwrMShxongiiAMWN
M+LjIgXTLfwSeO1B8+T93Crd051VKbc/SFw38fXEGjkyA9nOVLGSlHs0ucVGR9Xr
hQimNv3NprWu0X5z6+2EJY2BoYkj5+KxkwWX10C/TrdFw0yzJGj2TnEJpa5Q/3Cd
TTY+SLdsPSB+z6C5iXqIpKNz9V4ojBcWOUPmKTMDJZqAZ3cYPK5ixk5F+Jdfw2a3
TlcEup8B+yEGr5yjsC/xuvqdRI7vioURCATZmqRVk+ZCQKDnQSYU49xYky/wIJzg
fkyzFXQMRHvmwkJIALifomSIEfvAJ+QGDJlTlJm8s9cAYFFTr4jso68bgdFN8k5I
2qSrLS6PhU8sxGHoQab1mPucv2s+pzYMPq1DekE5qWUT2mRywQuj8Zd6qBnKcgEe
tjrzpLCJ5DckprxFgtN8VkO0lS/M7LmhT3P49nVTCnQxuTsssDFETqu7HobW/WmO
Sqtf39rk9SwQ0SCratd2SLyO9+MJTb8B361UU0kB7HkJkqviH1bcr3m5Fvql7m1a
jDxFPOY6c/5bxwv4UNEEfYmL1TJlEp5Z71y7/pik+wYQBs93xAl4dZNdtHneHeaF
98OLL+ip84PEcANS8Z9AKBdvbEzDbvKn9qPa0z/f8f2ZVYgq9i7mX7zhsTVsGlYM
2FrPFkYpIkvov1EGX9uPiPJlXc96qh2zUn9OxygjGxheNvZkiikwtZ0r5OfuvNOi
B6/RmOqfUi6545g8lcBjDfgXExFtubhdjgtI7pLsWwQg2CIdrr//CPnS9YIJO0rs
I5E7PnU2oZbAkGz6li05797nGKz4P3Bzp+R/nFL7H1uiFMpBpwrpmiaxYhhclZhA
WEPdUOU/vceZAqS91C4X6DrxdWwiT+gqSBzNrQd9bpNX8z4uu945SvSvR/LzmHMD
SLd24atxnm/H5TeExv65dr1zc5s7DDIc2IRvH4um2vbpOKQCQFx6Hk34Vtb9y4qb
USfOMgOFmtuRIr4c46LCrvNUSFqRsougiwrbPfAKD63KmwxggWo75447ayZbk0ly
FtATelznZd2QAxd6CjOTrV7cIhAyVCJ0fe2gYC21Okcj7Ngr6+Oj2OCWor8CQcPm
009HTwLJyOc+Dkkblc6l6KULjB5v5UrIiR7j9SbZTDlZ9LWXHt5xeCPS8N3t4ubE
p8gEm8A9F1eDquaAhVolyu7McLC6k6k1a9PlbnfYxtqryb6/o6hZTh33pefB6Fkc
n3KKlZi+NpC+kNReJctD1loaGBA2jTDkgvuv068liMK6VxJ/deHSB/CUB6rtFhs9
+SuPVtpuIxY4BxTold2KbDpo+B7OWRI2bLJMwGWalkxI6aXx5PkEQKu4ZFTLluz0
XwEX2gApflVPAxATxG59F3xVGXglozCTCpEgxyaykBuIRcbp74kBBAti79c5hyZY
fFDdHlIBSl0JHgptjQwTSFdr98uG5R9eIUE63emplt5RD8y8MuUjTjyxnmYhOVgt
abj2FsPBBhuzHZWkc9cx4YL8VybC/6RqNYSgPmd26zbmNXk47UZ+Zhh53RxDYicD
fB/NoaAxK0sACbAyVrjw90g2iNDsSWRn/e5TlaIvGaeiztC8wOuYOf8dte9umM43
xvv1q9/VZ1cRzPjoD5hQxFDG+rZmTU8u+BFAPvR9M6QH1wp5PsLXiOOs72s7XZqL
iI3lp7lfHFGDnTZRexfxutteQKcrATuGTSYM6fBbBvsp0nwv5cAkFN2x4TgUJJAg
IvSZzzHyKXJxRspeA9uWfj+oUIrzTIvuMHE5prE/bRWDvEXD+SXgFnN+ojnblXUQ
znuzjJrRoOx7sD9WOvTm6bswFGIMgcHa5WqhKWlrGGoKDKZHP43pyYQE/uJvbFnB
x8aksp0AW6Vwe7DODcPo+KN6i9pBd4XlytKiWr/yXeLBMJpqKDsGYSNW/iw5SbyQ
I6nhnrEkmHXsMTVo0WDb/UQi6Jt2Fm5zqi1y0cYrJ1hrobAB6ZC8b/8WvVBmxIk4
i/0HCVnNx7rXC2Ehk8TjrH8Lc88dMqDV6MrOf1337ztio/y8+RgRGyBpfuemLSyh
qt4IM6YOQFOXnqFniebXklQeCUnzxDI/yf+hTRGzpMccvIRtR7++lwZNSFWacXnc
l5q3amSTz8cHyWFz9Snp3Ip4gPfVTy/nR+rA+1BZUA/fg8i1z7+8UjY9UjBrWucO
rM9zFX9cSoVsFKjgz5oIAOFoze0FVxQoPsbznr7JtgdTwWW4glaAtJmeDYFtSJ3U
SfpQhg/7+lwfEyK3biRbn6H6EbP4uwoD+xN5D+CZkEWQrCBNHUUfnZIaXjHxpDPj
wmMBnoF3MtVQ7SeMk2sqZZqORnrUxrPKGxFUb6OzTvTs+IYqSUnJVW4Daznet/3C
Pfwc+mnkzBU+UVbMZcEbSbjHgkCqYtXIykKhrDw9srBB2d0OZL7gwT/aqdacPN94
UNefdrPvpDXliy4uNQrwkkTkdLcTTPX0ozKiuIY637bA14jQSlzoonEgAiSGg9zo
a7Rd2PZWQK6sB33QuyLj28HX2Oqp8JpKJlbAdLuVGK3J5/adeqck4iEDefplCyS8
6d4nLHojfSlf+jEotU57RqaYrH72K6tWN5tflyL+4WbzfmH/qAp+JlJihpMSsx7b
qHxNOTDUUS4oLq/Kd+3sWxNwDUJj6YgS0+8nzUX5p9X26fIEPQv5iu5JkjtTw4/m
J3DkGy5c6TcvqamgpL5cT2kirBayFK8xp9DYZTU2+O7TTBVVn7nz9oCVhQXSG/pN
4ziN1vCRhvXJAqP3TetKWK//k3dF/9DgKveYyc1BHmfI8bSoXmj3k9J2kNeevZsm
VcCUjmqgkDro+JzBUABtVlkY6YO0rBQBXgzKUlHcoSpFyaGKlD913jM6QCT9E5Vm
qvpPLETDlVA0J5v2l1Nyc0TEskVpD5NAwfQ5NeAec+EJY36CdJgekSAHp+TSJ8F2
IGg+fldswbE4S+Y3/P2mKcGQe8I/0TUR0ao28RCE41LtFq2k3YtoQq6EDjvNOXKD
Py8dHL/NDdR+HxMPdg4iZX48SqFir8h+p5v8RADXgcfLuC4jdQl5VEWWUD0glONV
shksQz7imw/GCvgiXbTy7rPNZH5L2eNSppwJ2wcq6/nHc+wzdPmCsOOIxMIq5E4C
QAjnM/P93uq2SSRh7qA5uVqQYzAqtv7tdVu2aANBEp111EpE3sAHe16574tHLQ4C
YgXvgMHeS9ykAJ+6S/el3MMdJuJYIImPyHnFjcXEGkdECNraeMraNH6cIxYICDAG
+qk0vQz6wdyzapMv3pPR8C2NBCSFPzlRGB3pugMOPynXWO9MvmCDMZvXr4TXTbNM
TFGSo6KYYPN/MZyHUXP9cPI8gz/s+VPYRLyuHu4/qPkn5WR/3AilMcTUtysxbPO+
Q3HiiYEmzVbmJKbMRsID3XkYuN3qd8O3USy7miiHreag+Yn911Gwl/pASL//S9Sm
rWCbEu8jJg/lOhVnv+d3GFEeOf2o7l+z5JsqC1CrvKAD95Eb1KS3wtDuDzIhIIoj
uiCjQ99cYjoSdv50jOIyQsNOqE1Eby1SaxaICzD8kcOgULy+Al7uPDWG+ZCU9jwa
HX7NjBiavVKul2mAy3GmJvKK3d3IvkwSTXPHvMhnDF1tN83AtDcn874agZHu7zqT
uuLZrU5KXoJqrZrch8x/dPLLGYfBKiln91+o8t9iQBmuWQz/DZuK2X13SB9G45tw
JofXsz6WhG3bnkzyl8WZ+bsiYGeEoeJxpx0+3T+5wZpoxNmnRONjTTOQZbC7/DFf
VmzAdAdMJ+GwtxGYEAbokZcL2Rs6jy1F7cfmZnh4dYUagsuIj/ELAJmzeD1PZZGT
t05VLiBja0wywgJC6c99WeFm5DoYK34VbdTngPbMnkELTasohod/L+cCMeNii+OT
u8JiRlUaqSoZZTYI/1qTpNSjlOOXAcQLgZzH+8c0H/RyNS4eHrTtwVreVx7+oB+Z
wVORgqK6zf1hQa2aITTDQEFMM33ystP9GKp9CxVhrUZcUImj801FDsskpGF34/7z
4UQss4En7BwktlIUIl2srd6O1UYLtoWMpMA56gvIMFS6xXScvJc8jKBfILkfFmlp
knP7EXTHNWzkpTht2HC56yZg7Rnkc/2bNWgL7ilNPD6eAVKBUzYp0NuLVthMgreh
XFLORhKmlYpqW3qBqq1IwGiSe2AnoZB2fQyrpCRd9uWU8Z4IjH7mpXRYJ+ylFo6A
hTqWE5bcMV+teZZ47R68+Ud19jW8bnr+9gRVsKGnRqoGvZdoP9PcGTaE106gguAI
KjB5Cv1ls92CKIdANfRV5DRYT0mBGpWKKAB7jVnFbrxg9tbhEbliHk0cA9wRuHFH
lJrof+pZss+/D93ULHDCyIbXgbNleVomC3LbzwOSImdV7rb7bZVNCxuBvZSQ2Emf
KWU+luTsW4UILZWx/bMRpk8V4prYfHO6oASnj98RWoI/mm+BdLOQupcm+ufwfMDA
sgGUbP48HDxqYNhzY/96uHBtGAHeArDEqyEwf4BxN5D+TO2AJ+QbrN5bc3i/d5mq
EDc0yEWlRVHA5zRaM0/sxHJXS+/8gVP9px5Og3CqqYUoa56Nyvt1fr3rQ9R0Y2fd
RnAwrWpcDULMeFTPkiNNrIvXAMt4Y0DWSk7wCchshqktKTapGymbYagYcdBuNllS
v2rX8ToZXGyuG+FqXyujzfKOh2pxDQYSBHYQAkNT879cc27sGC3mSVnWjsYoADNY
h3nWj8t52kaJlsxVW/HB37PESKuHrG7rFzAzG7PBRuYNBfu/VcBx3/AtVlH8CFzn
/CcCXA1QFiTKgmDdnsagyxoybO3BYv82t8+29oOtB347JvyIVFrfYM4jtBjq01rD
h5xXJpu4+ZXwxi47Ak1TInfqq8bYK1+caK3OS+uJM53pXfRRvHEjW1fMDf3Hdg6T
5ygVHE1FiXVS3tZpgMy/VsAAdNDn5XcLbrlrcZsD+VaFUmJ1JbhOHsRfXLKWi6pp
mmcE0L3KIZtb/MOD+mPfiaj7pqNJAI5xDwDgn2TCkhKpEswY2uHpdlTrkPi0v2z+
9oI5qkaHvBmOHNNREUVqMhQQXBM3TaTvO84Vjf5D/JdGxrPWM/RXFekncSv7YtUo
wT8xH6xRBzQOoxsrfHvBd/v/W9W6JvY1ICPrKSI7PHBBObq97XOqRV2hYlCQNJJ8
BV3aYpIOBFTxGY8B+7XQf30Liy2A1o5KfAmfMGsSjEjtpNvpd6mGD1EKN1IcpNMk
To3tLxhF9jts2RlzMNWVPv6xCPocxEZDqAtI1HwWMyzGJ5iSXXNVjcFTKyxLuOX/
fA7gP1nUt4iPMJJAW1s5HBug0/ngP1WUvgEit69u+jr72hrhigrCTN5EXuAX50Zo
epkRMpVmsBwZLTFSq9bScMuPYUIkDQAb6HtcXbIrrHcLWmUZcU7EQZ9WxOTvZmg5
9DRjkY9JQ1Akv4UOvMLrop6RUOzAB5eT0rZ6Ai9XwG0si/dex/0znhx93H3I0DHX
EAnciTknZRUjesNXzjEuE8KufsEcMU0kgtMaNUHzSmKD8+9z2Oe3HWzED8CBYMlM
jJAuiTv301hSixXsh02BnGqyiQ19XR9K23c6mAC+Q91hXkLcWqHaxYEKMTmn2m/O
ax+UOpWA5cC0vGVGyQgSeqjSwXVuOWTCX5Y+KguwPF/bPbSBGb2ZKS6P7KYzLzrA
0OmFZm7wPA7jyr0LxjLdjqTIzs8M3gJLfeUblaSHnE7emeHfCf1arM+QcXVrZOfQ
1ltvOk4DHpa84fq4g6OTJvjaQ0hbAkSP3dSIsQ3gUHhho4l1HwaomV3zo13/CfYt
XF9yDuvCOMZ0R30uYGJkfmhgjeN7hkqgwvmvvEJyg934gpqUpgPfEocnuF1ZDExJ
KXOb9iCdlCq7CddqfLTBj4XxzCVnTno08qsUfej78+nwKV2D3wXHhJnHfhN01Kvr
ERBIXhM/jWZpSHBBar8wnWbdtay6dJ0cf67gqd/2sKum/B+DcQ/cLI2PkYiVxgpm
Yt/Zf1IYKelLbf6KpbJykFPrKN3HwXjLLZafp92ywhKSqaAlJL+xiOR21YI3PZB3
YqdzOQM9sM2uMxH6TqxHyzpYRH09Z9JD569KuaSEps1SAqWzIaxlL5QXFfDLX6MY
86nh7SZmqZbaxraX4kTzAQw9PojXIddcbqObU0EaI75pb4DCDxP9F4ND5GRx7Ew5
45OgqEjBo2nzZ5Wx76qkftCXxeb62ZQfjo4mR4Q8D/ONm3Xf4FyLqilq51qrXguu
rriJsY+brzlb1GYOXZ1B+6QYCjtcRDNXFlCfyoti5J2KXaDOQohXPCYr3cP2W5HB
8+5qk+L3AbxrLGetoaqdUFM2xG/VtsWifiiEF/Emmwq9YW9vr5g7qUp3z6ESGN+H
sm/NjuErjHa7jQrWzhH0vrwsSCGqiOzsSq2qHuTSbXoUu/Ky1cUzExnPL3Zte8+I
UAGL+Z/QXrM4VRMMkerMNnWvxPRMhG5thiNjYaVjpj9taDbNWctPqnB0erfAFX/P
rYMPnCvgnsw2fAzOguvg2+NXvXS3Z6ZAXHOecjLux0s5q4suH+rnI5eCtn08rBu4
pZ70RNFBQoWwRj90vWEmVRlmN0x4OWA3InnZKG7IXO8PJ+7WqhIBck95kg/B8lpY
vsSTwieLlBStQ04ldrR3dQBS8Xt3axMpLQ+eZDGNeeyy24b5vQStI86O46lmRByJ
KVZRqttQGqM8LyEE/U9aQK9Jpqh5OarnMPE3IopsQ5/z8YBX3H8Jydcy+xhL87dj
9ypsXDgM6+gK8yqJQerfD23PkJ10GBA5/fq7Y9eGBvPpzkaADF92CoW7WO7Z+xj0
75RwZzRtfiMFrWZnUXYFn/yDrNU6CRopcNi9LgM5j+2w+H6wr8gasCqFiS/Mcsqp
8bb5vvUDFI9iHgV0E7YOZQrk63Hnzo/nTrQY+IDq/w5lG22mF9LEi8+3TW47ABUr
GlF3/KJzevHDhHMn8xVdTSnKKUrb6Fpal9o4rIw3/I/q+8Jl5NNWO+4S1eTihbb6
80Jho1QrnpiuouFYXTwGom9DgwDIgh/glPTBWH5xRFipigB86Cal8odIrXY6zKt8
5m+jRG2gkqjjlFLM1Yk7yHa9PIeVVBltZCxDjsaRjLvnFHI3hRK1uMZFRpapiDU+
JdrSVQJ0LWUk4MzR9d4rDlAc2lF+nmo7FIC8V2F9Mmv3bZwkLUlXbwKtmAeTNwb1
kL58Vsv64af39yaWu6D/1qm1wwh1X/pWwlD6rSU2/rS753yR+iD6fu15FMvACWPQ
7CJNzMC8G9Yrt/cikyLe77+wxKnwrT2VIgjAVlW0pQhxd6EcEsA2B+uuRXL7Ue4U
T4hxvIeJd9EGwsF4MVtj2AZBMvGVfejKtbbRRDwYuB0u1isX+Z411yxrFxxB74lp
5s6uZlreDJO5dtLNPmajuLOpeN8hPqpCqA0mAmElKv5vrwTSmU4JzSMyMRjOfmF1
PqLJl3jbOuNU/S8MH/2wsRkhczXzSgVWXrRc5Y/RFMUx6emtpGXttTnfs1kfw7nM
XS6Z+q8t09guF8OutZt06xpP2wefO2blT9LAbezJiYVmk//fNoF+DPP3EGE9Cpmf
qZM4jQz+ugo2C5lcRV6/p03Fw4sdru6ucpi0C3HzBYGSJbzGn76SKVwrydr462o8
scILRfYLRfbgXkMR9nwJZIV+zyZDqvCxbqFI4MQGo/NXxCNw9W1XcbNz5Z3ipXjn
UukQN6qzsk8zI1iROqeFEyhM7n5A4AA5ddk1laOqKwmCUiwM/xqZUkvvEZ6JoiCE
M74Ib9I3wMucDShpLDOYtn31701qwSsaUXXNlJYk4AiCms5fbxPU4aRgMowLwY06
V4e7Ap4MBDNkHJtKiljrpaDhqUCFVdg0y3FaJfcrWFpCfxQ8x8RTDT3fLUwZESKN
TIbNse6w1Ehi1KYlE6dL2VO0VwtPEGTotyshJSahKa/G7gXhQmO2DHKCRSf3z8RI
SOM1suSpUiYmi7sWvqaAr4MGfQLtksKy7mpH4/rVo601XnJDR35Jh0Oo6W449oCW
5neYJ8baezxJ8kH+YAGigR8cwQEMK6IFNUGAjWMiVVUIGS+8KEcyfhb8Txa3BIkh
QGa6Xntx26ThJCMDdzo98Hl3qnV5NeBwYjcVmJVi7iP/WLmclC3ZeTAw0FXwe7YS
yfnA0m9tFu33JaZc6eMroVmZqJXaqqAP9j7d7epKXNo41oAvZGHtlrUn2xYTDbp4
ewbCfgH2oGyshxu+WNBBKmQnb9bVYTQgJNlzDZ0L1lc8DZQ6UEFrIfGvTMlt9EOY
xFnV+CxrZvoindBMhna8IQarEwJZvcqB8IhkoY25854Pohq3fOe/xVGpKHuqNwZP
8rww9+6n03/ORUkZM0MNGGghb2hLq/QEqwDdCNKfXU7IYgRMj/WFUCWquNirk9hu
bxCCXLj0mS48OC6yZgxUdHdA0ZBjNkftkKrHEx08GEZ7EOBThGunpw9JT1wM/LXb
RKR8zBdPtEc/w++7cuP5AF5IDtm3UaKnHupzTuZxlTQ7uJM9hLxQdzOQpgnM8BE9
3b6eUtGm4txEC8thgyVEkzED4vM7GGnPC0SR2E4TNQdLz7TgYdDqyTbvrNCCuj9G
RmO0fxqNxfrWkJsEKCP5G5HH5i2m48Z+i0nJJF91OFDhmcAWb+63QFkc8jttP6/W
8lC+0PvaZErW2bBobAw9zGlYLc1WkF83TifkrFQPzjg0kYvH1/KFeQt6cQEBX4z9
K/P+UT52VyTeUhVmCiUWjtAGN6/BlH1EKRC5kCJJFFg3o58gkGKVw51C63ib7HX1
PeOz5LChkiYwgd7eFTMD6z24pJ9NVMrum8Ld2Rqb4iwnODs0KiaJ3zFovEFVxsV1
gGC5rXYPP2/FOD93ZMCSVhfMDC5+W97CUGqyjGuuiHIKxaA/HbRZWhr2Ka60ZmO/
tlC3fRfBx9Y3biNCbBV8Oau4+oT8GUP1IBSjhuPGntlp6YPKM8vtNZqXgDW1HXns
3DwHCnslmcWQn2O4mZ1q4MbMxkug8qv5W7yYCqAXecmKMz7siVHlR8orpSpGZmK5
BdBmKs1ofUuUBhE6ilu6J83vhnL1PP9WfFJah8vgGPbt3dOZOp5sIFJgljIJt9Xu
MVEi3TDCMbtiB1KwFnvRkuGJQuvR/jOIrBUFGIb+3qCrJ4MZveKnr0YIZiWMgZUn
xibFgx1jxt6jknG0ctp+vYLUlxrcLTdYCrodVxibRGK4bY14hDufTO2TM7swGCRL
cvFFWQyXb4+WHygKej2guS05GuJVjrAdbrLTPaZiA4HwAeKcIp4qRF4c+kGuQdRz
mkeus8X7h05GHk/V7w79Jw9Dv8veAuMUQZS05q8vXGfN4Xh/ZqQ7/n64Uv1eztkd
V/79+v2tNpHVvXe9LUbq0PGsOUiXQr1r+thk3g8iX1rOVemkt+ow/a1i82WRMwsK
G50ymTisT4QjQ1v4/3pOMS81xUgYFO30oURmDIiBfg+XkiW4eAAPUvlqot7glNnp
KFKqJpJDdGiwQxNTjwLkk/nJUi6L2NMV/CtgTLTWDcFNH+UIi3CWYVlOVaO4Fhpo
+y74jnC5Sz5APoWTAgCZUIp7WI1tuGGaNQQvweev3E2Akf0R+60KY53jgP+jvTHc
ByMblpbQ8yoICDMehco0bHy8cy1lCIZNtSM3bE5VthaeJyqPy3PteryGo3ur8S3O
G/mSPCEFhCf8NIXa3ta1XpOVvLNZZvBiploojiOHU9IHN/hC41rfIwRSTEZrUcJE
CpZA0EEtnCyHTULDON+WMK56Gd0ldgC50BiqddpvWTBYDbh4zf7CCiK+WuRTr76U
CdYsrYGoGp6rmdKghez7Ksm67x163VYoQJTfunkNhmo1l9i2KYs4G2/gVVfke+5i
uQgfSeVj2IMmGkRyndW4FSbD/EkOa4lVd8h+G+BhRfr7WR4PCOup9nDlAspcyuz7
8D+yjCZQ8EqRAV2p6gg1eyKkjD1IfuNcFNJkAdcNN55o3qzhz5U8hM/XqzCDduXv
NqC/JMnK7cjb56H/pBh4xiNdjkkJSoBylsb3sSzAdSdPRVn3TPFl6qeBCNurqN8A
3o1dCV+xd3Ve5qkwcmx7YbF8yx4LRCKnfP10JnrcuCJPfue0kNUubLtHH62D5BgB
63gPiQSS0HyQ19O5mTEy9yEELAdcYWjAbzZ6VUt4rc22/Jc5tvXB8bvMUjC3UUBV
wFqxdNRGtg9CwpjvIyWrEYVjaT5yUTOeEwVb5LHytRuKWfaeaJLIRInGlHutLSFW
dVy2gPmL7Tj1peDXzvsuRHV9XeYDdUMwE9YOtbwQy3O5/q7P6c5poinL91NvJegT
eWVNYh1fi0NXMKnw2aZ4nhpw7YyNL8qZFTQcmIPSxpqvXbWQdFG65L9QEUQdnVp0
zJw/uxs7YtMBer5HrTld5LcfNFa+FuhZE0AY3f0WZ6WwZZZlaa1KEZ/Y6HbJv/tL
3GSuk2a0Dnx6pQg+cwnbW0gMzSMnJ5EDK4exU8KElhUf9NOfkqezH5mUJ+x7SNRD
n1ryFZbqJkcQ7osfzLOputwEgZh9sLBp1fBJCUYWlGW1tKtlR7uSNKMLi1/wh7+m
dXOVn9uzv6AhXMgl8QnKxaAIHXpz2I6TwUESaJmUpybGDUXd9WZL65bRJn7qK6vp
Hc+WYuXdVCgui2KhBVDAG5Dk2Vfp9YZv404/rKJMdFxN4ZgPLccGSVuacZO5lzqs
x1Zim0NpssdKlSSyPsNH0PCWJhLJ5yMLfNuTYpka6WmklpvDBbMlnWMCgMB+ON2w
6hm42e77jJr363fQDaXX8B2lI66ZtUQQCaYnjFObSTsX+gcvw4+9TvFI8l+bC2F1
ftCAw3STlmfAUxXuy/RXO2WLd2KKtUvzzFIl+HwDOENF5Y1bQ1BnKcWYmCCU+gsD
1JjxgKAonupctI7Q8L4M8VMtPcrobT39rU95VwGA0oNi0jePTzK0eQsYWL4Rzy2X
GViW+I0txHmCKXi1E30Mqp0nY7Xz+8MwsPStUEl9LK6+M6m+Vrjkpiu8nQ//gEsr
zyffyKvIsslDoi3zdEmLAipzjAdrnBh5JInLVnlQ7Fe7KVxpSv1fts1BDY6KzGUu
wWyoKu79zt/KHap7HvsHBhujspW0/wH9TRp3Ar/xmd1Bwvw8kHiKqz0QbIfH1lO4
7IftSU9jNHeIB1lmwy/qehudjbxk7TLHFOW1leQTI6F7BxGTelrGsriFVhLEHn32
z5G1xkTq/s58EyKOtighoALGfdl9N4ajGE2EqjwzoLNxdkBvHu1ozYf0/7iz8HPZ
t/birBBp8PgeKxqkLErUaBBwInZ4zslVq505owXD7FztdRfz3Lc1RdvVYxk4Pft/
Kx7/JrjjD6wu/bpHpwECm/TQxz4TKrDOtd76gN0GBKh5RPjJpOkmAx27SBiIBLGm
gp4WkiVIC8mZZjbYjCSQka42Dbyl6nwuxs22WNUqXzUfpCTrWjT0Cz+uGJYHKA1q
CZcor06V/MJrWS5jak0LTe0aFjpxYOGDQIEsBVEV2AAAWFNtNvRgqcqxfN/4f90R
DG8fT1rEPF/l7397kGCc/q10eo/LytFz6IkvFUSdFo6Wq4B6ocNFMirjvGW8ZoUU
paINFR1xzZK6cZ6kDCzQ1ld0scHw9N0eVxctD+p804e0zkC+9g2VKDgQcKIRk90B
H8CPBh+GPw6q4ZZ+M++sejnfYa58FeK+4wBfphRXGtEKC7TmXKAjYQ3B8VMFigxj
5eZ4pzXEJ80jkmDndCEPLAkThga3jv/HgckNCc7uLgCaZESyUi/+ohDOLVrENXXS
sTPAuXJwpIOITbP/fha8n+pNTne8pj5SArqI4DRE34pa+3Ff8K6QlVftd9ECXKKA
7C7DCiq3HKrbrcQn3T0jwTepUeW/st30iJJR8WhIM0R+ThoHnv7OSrIu6EORw1hx
xYnMkuCFBUwf/KVkhu8JzmxILuspvYFAq1efvBnV+HhbPFDkSOjLs9ZH8YAGgA2M
b70opZNTpLNl3xWcNLtlLVvepKNgvWUpv1+ayUZrvtgXJ8F0XpsuSDQiwaHq1+n8
halnYu2lD/c1OO7KyKpGdlBKNvPZ4LZDZL2qPZldawPdUohD85o8JeEmn5hkV1CG
jrLg7iI08FbpDzPKp1DxbHUu4IwXetwtl27NAAqkDfjhcsrZ14AsC4FvarWtRGgd
6wOPgnGEg4V+wPU6PnIDy0I5GYtfUO2iSNN8eEeSDUsJEe3VVVZmOiexmq3WmcpI
C+AUbEWV88GSLLspQIUntwbefziVxyj01XmrAiz/CVcK0X+uKsDVWsL90WYwgDQf
x7vGTpnlx5W4qNnuTSB4UrUun/t5FTSDAuvEteKO6pzxzNqTzEqaVGjtH7Lg0zkg
7hC6+Jys6GQ7z45mc+uN0raLtC+TH93Vc8XrbBbrdP5Xqs4XQntLXZxJFMIJnNy9
Iyp6/EscoKAoTfg5zWCyF4num85Xybawdi+Y0tNnFym4JJqlCWGq7JP0t/LYNKYs
P9IVZcqfHENUQAbn845HAaPnixaSExA4/fsegvFMkFdCxwgTlKn3LOTpG0bPZsZi
ABSeEJvMklyxSNyqPUmvxhm/ybKA597NzQ/6T36M30Mw267GqvRdwdsfZ9mrRIBe
nwoKJZ0y7utLDT6bCfBK5z+z57rgedJnrQGOUrSlDpi+bTzw5yJhHEm37BbQ9xzT
4DRNwH7a2I9jwZ6crtF0mv6TBlKP2Lkk1mdRX2V8uz3E7GlCnIq7nJThe1LsX9xm
K3+DPMuCrqSLjx9195s3oJRs+PK5zAkeOJMJXKK5b0uQrPRJxKaNOwPSEMFPBU/v
2jqiMmfvceIxnGBCgCml1mUnrQkJiCmzJbv/m1N9pPgNDutAMP2YvXR6F+IZnOpl
ukhHI1TYlZCcNpBaBEz8ttPTZX8do80MRDpzyGUIISWOcYkSj40euBs7m3zQMsPK
3Z4F+PXZCrE0I/plWJOYAGtOjLMgOcj6Ylngsz7MrkjI17+1Sb3PZfJsJlTPZpWO
gWRaNTEeqHb42nYqjVI0VomY3Q4E1IwuT4Fhp/q5n9YrPpcBoiJvVyNi4MVeQQIw
5wDNdZeRmMIVeYdSUQtTme8owsb4K/Z9hH8XjbPL5RN5HNQ8v2yZ7ue3MAQUORXF
vo5ZjkLGflBM/GshJ50ilaEExm1alHdx3dCLFK2mtkjqtRfbdD2ZovLZO1YqDrO4
nUQ+8ZmAOsq8aZ/cn6PC2VCNT+qRU/2jTBsX1ydoZ7qSvZ+7yYIuTfbX4uR72jbl
Ibu8cXY+UI2cSWutZ8A2Hjd+Jcy6hNoFb1n8LQFImgtA42H9lghXwR7FJOaZk2BQ
TPwITMfpDn0xPz/6+wcK9/8R/ULrvHVMQY8GjRGjGM2IDNKIgJiBZ7nfrFV/A4WF
LVp8GcXGP59I6LCI2spGC3pvqvMXTlpCwjZeaUk9hu7IbIooa2V2hdfrRPTZOpC6
FeuYXD2NMQnG6W206zVvb/dBSU/p3eHjMnuSHXRZHl626AeiskOJHrZ1SH6QYD4d
72HnoqttSZkD9LkSgQlRTa/n5fu1aE079777qW15p98WLNiIf48lTHggc2iWFLJe
WxTxRQcfdTDZ3c3bXeSiY/uv8BJ2A3AEi3Ik/nW8p1mcCb9Vrbyv0FptlV+Vouyy
bUiH4LRWZUtOY4WSFlPZevqDZQ50h/tcw4PPJtLKnooCPamAq4RrxZ7jvzoY4lSp
BRbeid04XC7p3mMwhVKNS1r5TMuq9/Chq/8cIngn3gsttlfZ1qGpeIKwI78hTR3D
E3bC2PGgxNZrVYkt4oGH3UN986rNKBdPJgFCdmXo1mUL8FLJZAo5e2tjnwmXhNxD
vXcdnq3Uk5nnYxyUjDuKd5RVlzDrKJ6ZnZFZWnFAjlatFLYRHMCd/XvUzasbklhb
hlYgFGc/MlsDKYKYXEkVa2eXuOimTwDPOZMBQLk3SsPehrWw6MmaIcjp7zWFJXEV
q7BIOHXbYPkDT0fe+mwg5MQA9puPxU0nbDO2Cp3my5wjlDqNieE5GiTe5EFPXCeZ
W2TzXak8391EJvmZTw4zoE7u/SxA1OLdzqCyBTla6xGm/v2LhQCl08QRFAeevtvg
TxoyasFsjz9pMSyYavX9lzbqgmw4pXU2UGE/x401XMSb6+4Rn/c9AUxfsNEYenRC
Jb2ytjKTYZkY1VucrI8Leu8msQFWGap85YT3LsQtm3ziYYfbxmQpP/qAvaBDNB/q
ZiNNLeIlpvC9X76GwqEC4RfqtI+ANoGiBYVRan3FHLhr2c5eeTIayKe8383hiP4S
gGU+VaYIW/xdvNCjDDRbGUlHALo4CC6pjiTXTAppnTCXEyyNnJ65a0PCL8szBtqA
H8ESSIlIyI3cC0I7P5dV+h9vUGSIo4zLgoFh+GBN12T2c/wJHnZFZG+uaYT4Z57p
+gd8CfxOAGgrpJb3o0vEwMacgjGuGox56uEwbnkYpUh8kASKKrSIpJ8Zcnq4e/Fy
rqW+SsJDW3KU/E59jSYfAz+7e2WI197ofLZ/Tts13SrDZgJ1wj7Ca8blhY6rq21d
xZ3q3fwDnB+AJ91VF2PbepT6qqaW4OkTPmQwDe+E0kLaufccy0DieQURQnjvPWoI
rL3c5Bv30donMq31+vZMuLqTeQs1I7nWwnaEBEWswsqulmmU+a/uG3M5AZOY9/PJ
4+EzwetrGQRjW47N/inkZzp7VgVEEuqBasFy1w4lpJ6CVAyWTM5zQL8gFZfM6tBf
1D/ntZp/xEFQ9o7rvK3Hkronp79GcEaJDNEUSnfst5UtnL6gJH68pPiGAnIShXNY
PYr5y12Bv1tLHgcKFU1buTM+6JZns+hJ5nzuoJelEEkaXuUArYGZzzQ8QA+Vl2ze
uDkYuIJV6ULFnPjrj3jbNfgESBFwdkO8aU1JjkFPJqaqhq//qlsiwyAqTf5X60HJ
8ODa7IdaH2zjHTNINh3aGDrzXW6gr7rL/AcA1MRwt4kSrnjZ7Wn0UBpyOYbUI1WG
QkS6H7vbVjOGj5GQbHG9uTfYsjgldUmtCCTurKDxlZmr1MDJbNjlxsqyDcCuq7tI
Fxi0/+DxNwmzu7V3xmwSn4gKWCGiUuSRACfknDfvC18OOONj0sC9GYD43sSR+yd5
6q5+E0DnwUtzHVlHnpRCNab6OxpmFLjiG6MiUBxqgwVKPyiM1nWNQw2ZWGpB9mSp
6w+rrAczH+NeWCq5VEpRpNgJHdMU7IsyssPvLX1WSJPxrGKbvlHchtCpV6TNkxgU
euRYl8fUalfls2dOpbbwHOvDwwXK4dV+GwGxNGQ7pDeh/y69CC6jJHnpiHQ5t+55
cJd6K1QrBceqTHOrlr3d+f6PAnMeRmyhLHVOSBVb2lybKWr4yPLt8FJLjjnpoKph
VokcZFyalcVHDRTDCF8U97w6s1zSTGDU5ihsJeJCH3gn70hAX0vvWMFiA9yl0IsK
6OfT+/sIR95vBTOLbXD9146ULgKyfNC+zyO7L3TyzSIpfTmLuXWeNFHwSwPrz8Xc
Ef1KxjiG0pwE3bomaQaRPNZSFBEfXwPUa2t2AtcvV/GpsWb3YwKbwYEtViRDQSFp
5oIVcsRP99B/XJglPc5Dtucp6ks2GyBsumhMLxWhPATyjSs2Txo/bfbCIh6UyXWj
MLCLMmb7Q4njbpkQwx4+DC8JY1aNjiiJh68mUarcZAx2m7bwCyM9maopVUqaOMEU
VvGxEa5EM/kpWW/m2skRB+GIDORzOh+egqeUF2Vss547YJKtzBERDpRw+YCrLZO7
2vp9EAxDnqEq4bsiplPj4k9W12Mm8UbLYlzt15jm2EiNgaokO/vBbfrVwLgeHEAH
cT0D2l65V+NPbmpZczOiEzGHE/gQmzog4TZDnihdp/uXMQrksYmPx4qfsDOKOQ8r
zeMTnD9paxxYgtySYoq/S2JZmjQjljRLpFNSZRaXLT74dFObb6jO2R/yGH7P2xxu
ZU/zPGI4FA3/gXfknEZZja9BwW8NDkBghw/AMs5TDzfSRJwSN8g6rz+IYGkxmSt9
b0jcsXUlrBsJ0lX993ueTRJEUHFEJV0ekX7c+qE/SRWF4lwWNxE1az1L5mlVw7sI
Qs5Gv3BKvA2ich5TefHeX3CaiDCAQWdtUA0oxjkIgnAbxpPm8iPZJ+WCzjmu8KVd
clfJP/3AOjQFFgLV5TSK2EwrewGejoyXdRWDsZyFktTXu1U09fnMxunC2vJAb+WJ
ifqEEoItG8uHJM/loTj30RCeU7gwhMzs9VzI2QnlqkAvsbDXnzg2wcMCjPewkDCF
zficI53NOE5LGUyh3KteTpKSY1x7iQWHw5+kppYcHkVm3brk7WcZv6Xdm/x5u8AS
LnK41mk8BRjfoxZjomVNnSzToiAvdSp2Lo3XkmCk6sCollAu12HwT3RaurKdiU0L
auz+hTJWzeO9gL/6hNBtNYTD7JVGObD7+QZVpUjRQcfS/7NuyXVMPzk5ywKTOBV/
EZHV9IXbJJnbhflucU5ps4VH968kZUTaqmVldRI0MaKnK0P6A7uxugf4Ab7fJ89L
EZOmTG30wEHQa8Tg2C0u+D0EO1xXbO84fkVvK9krTJobT8adcXQn12ZgT/pZPNgb
KarvaN0nIMmRchvDw9gzsToQm6p6TH625OBqZ+PwuSok5jMbWW06PS2DF+9R6RYy
IrCywF2Pk8c15G4C9cXcS8Ke4wtYiMsg8fk6oxLLcrBLVSPoloW604MjVRxqflzh
tyJrK+hpHi0nr2x1Oi7rSBVjJ0AXS2eGizjWJSgqYwvKvbtS8OxY8YAqIxWrH5rj
M5bfyI3Fu5PS00a60ePt5UYEhwfmpoaLJRMbISZu6l3yDAdrUhWC0btCYAE9bydL
5QBX4Ep9vaR05I6uoPHOsmaM4FDr/uBtXtV6/0M2/Rvrj75KGevHthfpfhsFcHIn
2SB0/dlx9uxlXE7bX5rdsMpvJrvQtLmyfTkIevBK/KE4NzWWVp4pBgwCXMtwpGm8
4dst9IiCjK61afLurWxyyrpLWcdLLDNyjOIupIJDhB/qJRJ4Q1fZr5emvLObgMVs
gzWXWHru34w7x+KCn7qEKFPYemfX6PKXMC120EPmJ4jOXP21g1vbwmWbuzAQFT/I
rF8cJf294mZFx9glZ3s3Z83/E4GbY4DS5mLsWDVxhRoJT/YowdaZZoh1QUbrQisC
PgWTjkOoiQ5Hb2/THLOzDHnBkmfa2/vZufesZzSEBpmtcUflFeUPfukStp8Sxosy
gNZU0U72Gsb5QT5YHMnOvfKE7uwlOz4NZwn4aJHJ1XVWAuwVO6CydoRNCrtqu2kQ
VvcTBWPIdcoJpkzxXS/GaPQwT/Kyntj2Wgcn12Mt9Ldhjw5418pgry4N0AlY+/xE
OJuKpeCgAuKUIo4FHCIdQXKtpC7TK789DgHbKg3ge1SqpFWcJQ9JfHTENc26uzw1
jWjwTKGh0m0vDGEs0e/odIxAONhLEJgc2o4VrEZp6x0Dsy4msKdGAIgoZGC6LWEH
T0SKawk0ux7zDnGC/E4EXr6hBfDccLeugy6qY+9VME1pqvEaqdZapPRcsgn4YTVB
yQN2E2yauJeqqgFLA7idKBODM1Y/zXtTXZET94CLXasq8hFV30NcCZGlnIF+XfsR
Bcc6UBEq6rY+rc2qYfvAti3Duq7yqj2MVIK7DsGjoh0CgAYG1BOkiWvN1e+hfISV
fqKOstS+Q1z0roSVPyzI5Ysyu/ZL08L5rPvuLZR7EPI5A+QtkxC0YXP4UBFtXItb
Jj9Ti5d4VjoNB2u69u86/ahQLOqZAF2fvQbsicJ3tQNS/vQBIq9RYciR+B8DFSqx
4ObELDKrpHV9K/tX2xLAHzG9y8IXm45UQtnyC15XzYsebvU/+icrOsGQElDTwxcL
vgIWrxVW6xAeHW/SF7sPdXbNd5YMxKFJ8oYLJG8VwIoqZKdozSB9yawEpfx4EnpH
i4UgTlse/a46moDxL0M2rYWPT7xtWGEm/OuUmg2KlnRKw0tOdTXpS7y7uT0IP+8p
TzO07+iwMybzxX03XF+cRqhshhApySn6fAhOqmL7hH9Q2JJ/0BTpvG2W53A/LfGf
pnM9djOwin5GRghL3jLk4MKL9TjFiwiI8+0Hq6XuK4GB6Godv2SkuqgKVGEa5nx8
neyJfU8xZGE2AdJWF4nBVlm7sFUgRlNdgIY0dvuz9YWFMztBMxBq/xoFkEJo33An
WDWp0domoNZScLXuh8Q/v2rg95gfgSJgQx8H5AuS3rLlsgpN9gFMKlOx5ZF2vw3W
nuAj7EfvEbL29FiFyme/8bYvXfCh21caB4RSOhsOmJIbbmGSrTXlQGm9vhgOoyt1
eJQKm9AV9u+IGOqfvdOcc1DkrCUrhSNQopGo+BBH9F75D2zE1in7g1UjNlZm8FoS
bEX0O//u6jht9IIRfb3fTvu+wDNYiuvVn9rLz9SjV0T802kqmWBPDEvRskL/yShc
1wFeeisrp0E0t03dELTE9Zb4WUf1a7fHFlYVxn7aVyXCKVm31EfGdiLXEG0HUL6n
EKdgB6vmZHG/kzZw0csbYmIjpWAqiCJP3rbWMTyhqDDDroZ0OrY9mBw1deBlN6Hf
T6Lo4QnEK37KE48Dp9iOGzngiWD2ZNvl+iGW8SxbkFkWg/Nh44C9Oy5GrwVhRbyU
AT54N65XE5eb8nRq8Y9nQ7KrJ5L4OlAWGZpFKZIaR8c8Tm3Qt3+j2MA3nu1egdSs
9ZFKrdFr0iFsrjW0QRvoDPYVAURCjkrcOtexwexfndEtx8dSmKX48DGTLYYHhYhG
LGrgOUXrIDmsh+WEuSd/00TOJpQDBii7DGQILKiUV3UhV5+6ga0WbK2TwCd2vCW6
HhUR2rg4Uk0l4CWYSiaKMnF+h6lWa+UrCfOFJn1ZqNLD+NsJmCThb7LFMBJ/lJb1
H+6tbJuzPGmyYIONIONstF4/9xGbaf+P/6MkWTxE7jCC7Y2Bxi+X0GQO1byckddr
O42QiPeDdEErtLxroTZ5t/nr6nHJ2D7K29XhAhHiOqcljQUsmQKi/HJtxbCZy6TQ
gpE25WztgUUJ+6VDlZNA/FfYD6Zyd1tBslxmTwRVdUu0dPeKVPnUtjyiXjA9rSMw
oy1CLWXTf3qjniWgcRSygPu/UDHxxH0URlqDD17x/CWQEZjVQ8sEJyUphFFVjsqE
fm0G+0Fp4JrBzZjf2xhnyIucBg/MjZd1D946cgs/prdGGLVAKhDGvES2Klppuvr3
Ms5ebrYx9pkiAbEivStXYVh15I8Y3xU2BuX/vJeXVXWwHczppYd+ngVPpuey9HgD
YBcFjCc3101mF3DeExcvLPZlLf7C4rikcG9KhS/2w1ORNU+iZFlTBpZodTijwHwT
WFD9kLklYI2Yx0wUHiKxXCm4dV7PmjVe4GO9RAWrH2q81brOKTnN5Lj0EgNFD1cS
itNk8tlcAPw2hEkQy3QBhmYHA9KY3Z2LulcaFOitwNj96rvqtM8SYrA3x+VFxeQ4
qfFPWnjQkLRZsnN3RkKsBmIBpagv7qzesJM0v4QNd+9Ew3f4JPa9dJr/BnueP18G
vDi9aiRYETR8ntnTfDdxiyPktA5nNmkZXSiWHYnP6OdSqzuBDK9ukZoSK6lzn42E
PaNI4MHn4bfh6mu9pvIq6HiZdtvZnXt/TQjAaDEBsi4MOCRd/BYoGfFCTyM+y0PE
B2cWglXYPMSLzWF1JoMoOMI1x40SvE6ZwUV61pw+3FudV3wB4wq5kafl37A9/0To
GYkS/BDwpctYKUiY++IA+//qR8urqgDU6sQ3GyRaHwTfT2PaBWgzH3XU5vBIjNRN
mOe2RfiUdSdHw73MiHyypcfCf4YWPlzp8YNPHBCOqLKIWkrh+rL2PcajB1y4E2pF
D9PVtTXQ7n/NnYYs1MG8HVRmjcb98/YvYyTOhLbCXSE+ninRwBBvoeQcSXcWudup
oiBJ38boAeQl92eYY9sHd5k3KPSZbV5bG675nL4gha/vPRC6Ky8FKN5ZtSpeUwTN
Ygm/lRlgxnTyd9pW16t1Nk4/vWnFQPA105x0zZbDuy2eBdqzyF2KQQQYYxg/WAIh
4zJ3YFOxrYQfDgQSryTaj760bfCPEkfn8LD9563rRon2Zu7BKw+pqlEvh50CP3ZJ
Ty5hjdT43tkpEb+8FFkcoYT3MPY+1vSpGKxHowJm9Vu+KIJrHCCM0ITkkVQQT9RB
ZxbuWv/DCo0bBtY/VjlxA/F794YPd4Lv+fO6upUERyTe4/QGJSZio/KxIGwkVQwC
jWbFRUgtFAd+fE2X5PlWIfGPZGXdBzkW8YCzB1rHMvHFHSXLqKRiUVvE002OpEG+
ow5EFw2iNOCwiorpMDAEO4ukb1GrixfS1tQg7qszSH48Kj4co/h+lncAw/dTzJ4W
xlzWYbcoPsLMa3lsfUbOUPZomlVxMU1pEInyc61fzBckYL4747TTMLPeqwRgSsBz
yYfxGnLIZ7Ns/18WT2spNP4SR7ng8YlVp5N+zqs8fClWe90DAO5yLvi5D8+OaD52
BMr46LTatNinB+EkcVJgQLbnePzt55kGq0T23bytNfS7tyCHjRcobDaPFwIKT5Mj
Y58tm9R8UCLJU1SkxTl3/oEON7w+fIC+PqEVFJnFn124WX2YSEdQrMAuZyRcJcMz
ue7G7KSE344sBHiRh4bIShztPf4cUDf/mBx7t2CshIsCfzWr4rxixNmEWiKYs0yf
1O+GwS5xxDOOXSHIcmYi4MdRUuXCfcS1MqYK8g8cimBiVD+WdWwe4VX3VHJEdmJf
sNayGsCdHyqXvTgHGK6q8EzvJ3JsuNSOk8RdCcnt0+3mOZJLe4T0mhPACM0J2zEM
SnloHWD7DJn4yhtJZW2I3UuxpNHcPsqOIASftPhlSGaAWpkMQeFTZDyN/O1MeH7v
y5sBvGH2s0S7TfhnXc8QEZAxuD0Moe+fpb9NQiPPmaJ2Sy5e68dIpcfigfhYAW5M
PiTo1cj92Vj4NKsv3omXj+yQH/7Zvay/WFqa0V3kd6mXkTVi09DC8XuJAJ6yYKE6
EEHbQhpnQgNHLiflsuTp9tdOBXGeLHf8hE96dZUr4jJnh7NL+WQvBV2wmA+FlWWn
e1FGtqnaDs84LN8dW073azYIJ7eFXPnbvKKHIZXJ9llkSZW6Nu7w1s/rKOYuVW85
dbDkWoyvU1J7pxsGXMwwr5IEItkybnZUd++X043aPvzL+FNYLMihABt1NoBywylk
C2/HCJB8Ian+wDEkgY20NJPVzJXzafduHAMQYSZiROyfEoPMPr0g0D1hrTBrQ782
3zIV+6BJbI7jthk9mA0MHQbWUEEOioTovjed97IDrDuo513d5RDOYRltUl88Vm47
WFQO5BfhyITYsMjCcWQMxkHhwU3RBZIisSTYAdtEPcoIouZfLPvPPati/BK8WDuq
pPSVH0+wdurHsRfEaRjgtpeELotCpq4CtIALzuH3B2YDiU+lKzk7hF9G8mYCxPyB
nh+jQAL3V8r7ukpGL/yvX6rFnqcvxwsidgf45jQ+fm88LHeX0uA3p0PoznpxU0u2
nFOMH9ImJu/eOfSImTlcS745l/QoUOJNvzIbs04qL6lqu9kX+rMsSim4OBl/ZhVj
pAhroXRGZYZutDH7PpSvOkx1EF157N3bC+L1uvjrOnTjsWLJlxbVtnW2c4u+XIBu
0WvAqEf1qC2eCHrB4mHOEzi1OEiPZ3mraPtsqxW5/v02N0ka/5rmUw61704EWeO9
C3HwLnSSkGbgA93cLzzS4Jd1SHKIDWehMxtBqBP9UBzbISuEne/T5vLGAxOmNIvZ
KYW6zhvOVr0M0JcNf2OvR+r67qX6vfo1qxdPGK1Z7SkpeHPXn9INmkgodjyVzEYx
R5NRj29068yC/r2qCPRKEjnJb+fIy3wX5wVwfMRal0Tna4JHqO1YtPFm+/yjsu0a
RrsreisUesGA6hQnjLw2MLEop0e1ZDxSVRHezyUbko0Sjiru+skiQIVsttu/F0BE
EZnJXyfKH1rxRoa7RNgmJOoj48wrYPmavT1BgeOkQkG1wlU9XRdesGPZqepDPxz2
KJYVmPIpKHaUdNQdO3usiTsRJ8o+1eQKuuIgndnW8yeHfl0U0HZFEUYp7aiMtd0Y
WnMfaXEmC1VllEyOaW2i2PqbRuus+POW7OM5un5jtoNYa/XiGyg1gXJ89lpRIX/a
TmB37GPYUUYpk08tR2Aj2bmVDSUrTjRBe4dj7BR+2Kxuobr/9sa0lFfORs1KiyZK
DrO8UDeF78fK834x2zrytf3fA+PQXc6wYNfkPzhjeDXfk/q84RScdLLrWAkrDbMF
nudqexvareEcgnQy8RJvMrwOukai7ElB4TGKq18wfm7W1fsc60aL6GIpeaNjMUvt
r5T35um5XNuvdkbUkScwaTWcySKQeBZJr0ReBQDsPK80wSqeqI47ZgjRsIJdOmoq
jo4UzAVIG5ZLGHn+9SSe7jPwabSg1W7ZVD0cr5IfjuHWGKOcFw35aKytnky6Qt2+
eTPkc5Y6QOym/3sH8IXZ725qwE7p2oLScGAol3gPfp7qq1hevR5Y27Z6hxXO6JXX
LKbMurEPXlQdc6oEOI5HDH0t/8EBqAPcOGN5elUwsozbUA+rXpOkY3+uW6gnD47h
LjJO+e9Y1BOX2sTk4xOn8wCjD3nARXlxmjOZkxIz4PiDsKl8lxzywnkTwB4ZYEK6
Ad+/JSi3Nm93t9NhK14txJaO9GdBJy/m7P7lPC8DPAA2JPlXW/rEjEmpeDvS2DSJ
g8eG1ntCihK6eAIQknKVJifJgtf+TD+w46ZFtIr28tDKBQadnimLgfWxVw0MSIKE
CB24+TbHCgc6yYCR4p2trhNulr+8+gyVZo/Py+gJIYTW+GGfwVZXEzHgkYXpMfPX
LkxCfmy5xEeM3+6UWrEtolUsBO1rxHecvgyNwDDjHcrEX2cWrObIXu4N4AMKUydZ
1/Y8ZEyoilsr5m0sHBHZL+PusyrlLxdxyU1/oPLINVIzA/3I7OqAfDvn+WJvjRCn
FXR6+QR6aL04NXZYyrn6FuRkV4FlZfuyoOUhFX8HOnhmSgzXMLx22DI9ctIirqG3
nw4AwIcRu1crWyhlFi3WyHAh2aMdTwYgUMyaiUPzbwwkVHnrUa0Py2gP9Z5JDSL5
rgfsI+PzIjfbqeCB2daiUsX2m7bqhbmnx2avcbySvKvE4OW2i35534dpTWAiJr6a
hzCRvJmvgFalksUR2YSvNHX0lh8HSqWMFRIDHp7dVbOJLSo/XRLuNSWms4m/Lc5Y
4f6H9P+2JQV5Ur5W0Ql1Sz/BfZoRYSDYYdtC2jT/0Z2cKaAESoHiK3xmf7pOilcq
TZqU6g6gKeyPYq3UbRlWsFe+vzUQ/Xe44NuI4X5o8btplGLmBLEBPLD4iND62I2T
smu5C8ibiW5qVQSpXTXBCtMWW9D8iI2q2IHyQgChf63xpoaP4xLqYNf3s8ZeZZBg
WgQfPwzLMjdKApXaoPfSwSsp6BV2eaJbfInqgwLX6GEvjjYspdyPadKzOmuUZJkQ
nilg0Cwx/yQsZRomIB4zMMttb2w85n+vhXVHwI09iJWiY7wD3lUJBLvYby1zJRR7
048rihUprBLjf2JTflD7TikVnuTDxTsMy5X6EyrLT5H5cpwFKxYLnfjpkuE2Nfkf
bzmTJI89wRJdEOExmJcFAK0QOjceUPePl+qwzgt7hA5J+jNxFRFiApTFwTVKREnD
LObd//EtEIHfTO44k7257tynDhLf2rowUtI4flXRxo6A62sTZ8VRqfUzbbMieSbj
5h+Ll1wOrYh+JTwpoWXcvIkrnEkS6dngpQ1Xtm6Ivc07HQGIJY73eHUGM5Jf1jSd
6EvxEfnLtgHPYTbBuZrWxQ0ZTSQwVt70jkKX8l1Q1iMc6jtDogy3foUcVPKEqP6j
kGlpkyDzeUEl5eEutpHu330hTgT4dfFO3r9M8Nnj+MYWCCXDm77C9+swAAjW74RW
VMsPcS/MbxZP62I6609W6LHXx1b5daJj73suHoZ73dKGVwWxRjovuDTdl+NNz2Aj
8D3oyB0LdX8T09eIekOGEe1PsmEcojJVId1YWjuziq19q9Q2yiElXbWyRS1VTNuQ
d/SznlE1ERfqtO7TcPo3uUCXnb/zxHMGJGwrl+wKc3qfmcV96WkZFklGTHVfQ/Ry
3ACFRCAKsYCu14rGeDh88cDSHf9/DZy2AZh8bwGOJI+2RTHDb8sruTbwX2zxyAbj
/QD/x+Z1dzQWvp2UWmo+vD+KnN1ksX+mie/TLxs3bf2oTWkICNF/0Y/9AIqJL14z
Nm4g0ICFoxc3186ixNOZF8zRhu6V3VV9jpG5uTT7vSd8bDfk1Uzf+Vu93IhM80pL
Tepq/QOZ3iCPVeOLWCKd/+eEIy2vfPNsnClUDUEDkdrhNdAxiIbWqqfx7IvFi6Z9
yFYBuGPDE6ebUB77/z8SWGYKparP7NKFJ4WffDXSeQpg4aY0v3wXhh69GrgXKHK6
gFaDdBs7OiieZ2pPKNeMihAK+xPVHFCGlseBOZe9Srf1bygUYoJ94VTBNauyDIE+
HJeftEDK1lQstvClYewFY3cYOyVx6IMbE3P4oco+G01a67zAnfHfto+KI9t6oEZT
AP3RTm5AQI7T/V/PonYpWyQ2kSByYVZHJatYO3mtWsnuONFRM+zb3RnblioYoTp7
nnDvbAcFPfwGWzfIFK8F+AwZQ/sN1X2XWw3vPfA+lXbQvVIr7t2SGBWsVLOngYt/
JuIfYybTjMLyKh4yXbd7HRXcl23hVQBFuZ9WKYFcQZqnxeFK4IYS+BP0R/SRno2F
ckr6udxME9y62jWIDQsDnTy/SKeyQNgVdyJGHFcBXMoAETmRfBBaBDxJnx1Pr1NK
mDOG2B9NSBINT0NfoPndRq/0DzxImOvuXvHGJvYtysdgtqYXHhRrpmgRtlFn0Gtk
/eZ3Vt62k2yvb38evUgCELgelKVeYJmamdAmyNvdSHeE4zLWQtTCyKD63wYzkwvU
XyRYP4ErE+5qHk1fgDiICyEOy4jRYfPrnSGORyYdn9rZ4HlN0/ZFGpPtDqKDnKTg
Jj3av3YOst6ks3wQImIb9NUBzBI5krJv1enZYdFPILOr5H8XM4rs72/VFSwSjA5K
VT5KZI+I/75iCiPJr4q1n/Ox3z6PD9tAe8G/umGAHLkI1UY/BdQNv6BdocG9zd7q
96Yre2lhFhAZvwm0Et0+HQDCgScYlOsa/eGI4LLizvUIfHHxnisHY4ljTredBN1A
KCwwNdswpKKJn7bJaPQj2tKVBmOD/f9u6e3DmM3kxQhHnICpkgPdiirBl+x2V6RQ
d44GSsA5lpUV0/mHmriIsIM9BS/CwYhFh/jHtiMNY5sirZJG0G4UXsHKaH3vMNZn
TEO90u1OptL6EnaaPjAjMKkrhLEWiF4YtMNZEOMOGs0v5ywxrO9ijhmE+sdUWACL
Qry4XCoxny9zozJa2EhquVDHvTROGkN5r7BxsjxQjJLC0T+MsqOl5f88WuTQ+8NC
RYi3o82AjKtv7lSGrsMSn+Xni4+pXjr09aBO61TLI43ZaVXiIBJGeGQ1PArbDhvG
5oDM4PtMwz1aN2RykNCJvOjHFlAg9TlumHxKsFMTcy5uTe36DLIasdRNGf0g6qMi
RyE2R9tLvIodtaDNoVtOPYVxWGbGiWzU19F38Mr80kIaZDr6bLEYJF4oLFJVOgax
QtN6rGoNhoPeeCbw/3XHXbhwu33yeAKZzmlV9kP7nJwq8CFi4/lBgRdzcqSRaTbT
FwyVMrIM9hUJtCt4F30zTEnx6zV8Ji348jtJeyJZVqe12kaihHSSgHFWl4yvLnWa
NVAC/tNWwpCG8DjnD+zNLoBI3V0S3uy0hXqgg2pIcTWKzBUubJaEqczYoxyX+GIl
nFJefRR3OkMam7WyP83wL4E03Sv4ltqPGDLZOzGj3uSL7lkUAeq/zFbkxdjQ7ZiE
cNjSBn4icF7ID1l8BpaKct/elAkgM1FiZJks9Z8tgdjxfe0BpSzkE7g/Ng/NUQZX
sisPUyPEj//jqApgZ1LgJ1ohg03eMvIV8lHDqRC9IF9GZ+Qx8bQ2hnDzxgGTvVra
I6xmiXM0rERNXwRPTi2NijGVbJvK4QcEt6cXGoghgmsIv2c/WN1V8wFXBN8gR/08
jeH8FX02Mui8podLQm6qhswDUVYopJzyi6RLejZhLBxxGjIRYqaawvl1GwX+kqp6
MThg9uM6ibBpdtmvnOgx5e41g34A4bE0vpJuTKlgYNnwoQLUTukmUIJp/zor3Ehk
DwWC1jpXExLBmcRprytT1lcVU00/I1Jw0nU0bnHUgDl0ZH6QpPHHwLW3ss3Y1A+4
uwQjIYknxmUvzNnATIXvcABxpzl4/pgJlNsHxNvHIWRZCRIdqfBJ2iteqIfXbM0q
3HRsM3F5QwbLrRt7uw9lCD2CfuBxh1lRID/fAVn3j89Yg1FNMj6ZLcX2Btlwa94g
KSmP7qQyHD68aidVAyOY9Ug7Fe3xVrjlxnZeTVeXPQlNlnjOWXZJQIriZhf97vxa
Eo5RawyU0MN65y3NKSRUNr45vGNf5LtbDeC+lUVf4yxD8M7+ChIH5bjvjZ4saiTE
op4ztqKVgyjxL6UwEPwattvqTSr5kcVsJdTUmLf5Kro0/rDp9gXrTGhBtAXoOudw
NTPosHFWPi8F13vkORq4If3EFvhIk3lw6mBuxxT3luAVD6edTITBveBqjYLOFf9F
zVloWb9fglkoQi2Cuugh5iNDDfq08irRSyYz6ZeSpv4l+fgdKEqwQ65XzARu1Q1m
G3FVKNMgZYEfoVW3WWKXSTcTOL5fkBcIL1aJojq7QC2TFH0hHG6mkD++dDduGxKp
4bfs3pRMHbaf72W8uqG4vSy70gzCSxYBoIyhK3oKvMLhQ+jVWJI3kfBhVk94DC/u
dRUJ2Tu7ZsJsNmj5h7d1NhZixJACALtsNeYMMwYh/PS+TotMWn7hFMAuYXOG9kRu
JqMxA4hYXNVJhwYwu9nuhSy1Z91eH4X8yNSEZqV3VLQR9bR1xPLxaaYg0NF8PnYW
Mz6S3tj3noTKPX05VEJLD9bSxd28E08Kck1qdFgGwMnoh74VErNNEQa7VyEqVSnU
vH/6BCTe+mrCFE5PqsbF3QmvfO2M3rKXDL7zQLBIpl8uiWbwP4iyDNlDvPC23oN+
zg+F4nih5gzqkkMD0jxcv1HQXHu+P929a2pGIXUxAiECzsVbJgcOJKpYiFcJE8Sb
iUJcC+dTtFDuTcGAvU+y2AV19TYecUKcEAjgmSLVO3UJmL5fpqeHSLkCWr82vSKB
jon27RkmJ03aAtZxyuRarabkd8vZsb2y8Dt89Dl7gyfCe4D/7p0rsztEGw/I/CwP
H/Ii/ZU5VCDz+RpwFF9pO5UUO/KpGipF4/4zYGAgGi0iGtG0/nMhH7RTI1iceLRG
Sh/CH0ysdZHvW/5k2qMxEMEjONAo2DF0FsxHq3IS8rSS11VboffEElHfJMs7xlr3
ZzaAfiHs700YR9S5HhfuLyAsU8Tf9a3B1fyODLtuqFTH/IVdGODa9xXXguFZ3y7a
PKp0hN8EF3x9qlyTfuQBlFdGPP0tsNf+tZwgjBW+5PJaeBug7AvBh1axqKLFqW8n
shP91HA1cZBKkD0rRlNpKPxVHw4JYaM/fthf7wDsP4uPh/6mT0zttObziZKW9y0W
u4PzBN+qWoWQw0eGB1I2NLZWhhzYXV/JQH8UVIRBj5Qss3Wn//v27Ovv9IzRN2dO
IEWXilN/6Q/jrMrMTWwgwOvjjPB5qy7HRSEp2Pj0NYYt4VosPX+BNfLlT9X+xM/Q
8pGgGl/GTKokeG+9uUkBALxQoJRou3xsSdO1I/zLMloIR/BaFofWdXTNuVGLW/kq
BUHslytDtu7nT+ga0Zv5AKBMEm8O9tKAJpUIqwGjkymiQq7JDQ2vpVqe7xMIMSlI
TlKCN+YCA4mKLnXDutYwIxr5f+KcuB9U5CRqB0DrA6ccSZk1ZxHH767xINbHS96q
nARHgLK4kJV3WIxWX1wdTcbYQF16k7kp+EcQvQy8CvzrhsV873+WE8X9FvOdvUTq
3EMzZq7gvim87s0RFVKw/tVb12yICGhTeHTsLTeN4Z4n2hzJcYUCd7sM1dMRO/2o
y1xeqM0qWWwChrhdWvanfBa+R4HwrJHGxdv2sG6+4NtexfVvn/J0msAoLvdR1VfW
d3lPRAgKHeTLUPkK3DhbIWRjQavoTKd1sY2DWTsuUOi034tykIffVUtu75TezuJM
fvyp0DZsJl9hEwcTD2P+fd3Bw2PsTpmIfJGxdsiwwtQAHxSyNjOF/Hu4PwzxSz9W
lNg5RKWi6Bg0qpqcurfU8vFcaWuK1AlIUwMQ9w6zGon5iaSebcB2sZePhsWs9L0o
5O+dvexzn94NZM4/7kuQJFaD1pcXnBI3J20PLw/8LfMgUrKKcg3vwGnBiz79s68T
8uvBlFcELzbBW0Vpp4Mc//sDwSyNOsbMbrefnQdomviF3m1q4Q9CAF2TXZZ5O8jw
SYb0VMTL1SGvcX9sbT25tXEZtJkKrs9gWDrJAqvppHnSx7h4YpV8XMV6Tnd+VaQP
nrjNzUX5qgR9DUG/L5KCIIX70LiiZLmYoVo5XUMxbnHYyobSUUFKCK79S0QaDiIs
pDeQiHW5jD6Fj8N4NPxvBqLZnvRXyXI9kUJJSnL9+L6LgNigy19KK9Fh0Keb1kq/
PCIrnfHoNMKFnyw5sYq/bUZ7qWM55gn83bEaY7d8XFmFgKNUyGujqxG3R3iJJfcf
LMM/Ik8FLKI54lHu6L6SvnZJz4v/1/5T3kQJY0XTwMgyCnnCBcCUV9ulX9qeP2ol
lUd6KkAFFixinziQfwrdwdGyGOXKG+Gl4JE2e5NuXR58uOaiBVxe/ZinE5Pon2D/
MY8MZMhK0klCtGexN7jPA48HyDpFBUoVPCCzhVkcCqZZ8/StpcwVwEsYV/QRF+UW
pROVOiOz+VxcumEhI4Px1InxHfkxsKTLZup9lHOBWl5lMwKBE3i59sQP4beasJo2
s0IsoGTX3rZkwu/hRWl/vwd7LHxX7b0cy/DR9pNinFF6c1QQFgKYMKdhI20jEvYy
TBbx/bxHFUhU9S7dwuJ31BssNzlUBhO9dLEUJcOvKoC6NPKUIFpQvFJlwBlvbT1w
t+7kWsASfz9DDLfQkb0xGdFEFjhdKGLY6BuHWA8W3AEOMT5iP2O5FzOoceQpdWPG
10Ohqaq/Sni3blYygAkxY6NW5DRmkvqfGK9ZQ7+tRzruzoeWS1cKWyTOyPwgB+jg
LIN4U1Erw7pakLTNgMpUDJPWh6jEGhh6jcMXGcQFrarnHE7tk/Q7wmTkjwkmVuOf
IT4TwF5GpxUqh1HtcTVBx6opJROJEX8m5xUUUEuV8ac5H3uMQKkGYsxY5JvPAVCF
YE6hVulEXa//ieyKI1dpJh8au+RYwtnRWe+LPaonLhaK/PI6xPYg+gpihw4a78P2
kdqXIxUaoLY0zdiPJJ9EWMg9iMWSypV6TEjbZZvSheQ/JeRVcK49sj4DvVyW1HlK
OpwdgrLg3Xmjg9Oudd+h7r8uNL/gqG2omsSfJ96+++Kxaib++qMyeonYZ8Od5UT7
ZmHah4b9ZiXW3bB9qutjINBS+RFh/oaR1KuT6tlQy0ZEbE75iVNU22EiMJXGrBbt
9vwbCu6iS9uybz3+QTPZ8W/eCZcmL90rcHR9Xn5n1t1RDM0uY4gnBdbobg6YkF9P
aCiTeNaJnxjBEiGwgeuaaftAyuZ5K1E0ehAzTjCtVR5OIjX7qcRH18+KJN9shabS
HinW3fLvDKuqlIMgslkF620Ymyz0bB8sVEeb7DLDDoCTbhYDwNYWvxBrxePY5GQb
3W2LHvhLo3YGS94Tiefd+EkImORq4jNQRfj5ydOGGYjMx+JIsIiMrB6OyERIq6nF
3OkbMDnHEauEwa4WOq5NupHhphYB6e+9PGdg6o6fpUU1bLhhaXLZ25RtjdeR/IAE
5y10r3TvybmwI1HoutM89DU4dMk6XM/qJpqNL/BTf4Q+nVvMIiovsQ7SeHkFhpbJ
iDL/cp6M8MJgLOPkS1Ox8qaNHRAZ+Dr5XwdbXi6y1HDp1h+hGXY3uFl0OzT3tEmp
qKY1G5Qe35fsNkCCxrZ38QuzFYJIbryFVy4S2oTP2BsI/F7p8Emwr2i35Ta7I6aS
ni+pzOWF7aHATBuJ9WnygL0hBHVte0bAs/tISiWV0goCIyrSdiScwsWII9AHrg5A
qu1dJ85dC/EHehqrdzqGr0f/cOPfQtqsxcmYlYYHFddebi5YvPzimpkfK50O8VR9
3PIyA/HZwP/GnKhGGuhFBRlmtqDd+01B4DGHv7zVO1hDr2OamZatgUYeA+xDALbh
A7mfC8lKYWWIAY5n3gJcQoEp575pgYYDZs/LJA7YGmqRgPYH/Hf0W8qGx3L7wKZz
5XYLW/VpHjOAoJZRvbykZIUrtgQA+jKhsmjEuFtfGuo4KYf7uTbtjHpvhL5pSFYa
+pToYp86B7FDH1paZ4AhF5QCDztu6Gr1VsVMEs7xMkz+cqCvqYr03U3mlZ3nbzOV
X55zTu+1O/eohIEFA+HLxZg2lHg/qz6UNLLzJcqqLRXVEncgOYw/UYDG/M3go2CY
cSlFueUkmpVMQFkyEUNq6wAP2xHr8A+GU6eZKbRNeOqa558SLrReIdQBnuvVerEc
LdprAjKPu15ASI5Th1jNvFVdmOQND70iA6uFuoDK1tBAEmsPM9OwFrsC6dTmvWb5
42hP113Abl3XsCBgeSnZaZQ2zUXlQ4Go+8v7tWm6eHCmYxofO+QVa4egFT7RakQZ
zeJOfySOkX3rxa7CyD6X0HaCa3kKhjMbhfOBEMF6ZrBS+QtVYLjgT2k/8mz0EnW2
w9iI7exsTqZzDUwWXzfmcPFuWHeIvWhTpw5imhhBeEXnnHuGKGLkgSy3cvdp4mwI
8uKm7ZYvSPiN8o5RedxpgE1w2h/swXYbhqn08Da9yzFZSApKpApiRNEoamMDEy/O
x5E1uUGUpEZ2jr0NfqHZPfchbkp/fWdeZ/jEh40lxLJk9qVwbTuCJslQp/UjxGA+
vAbuzs5Yw85xaBfVMjGCK6aG6Ur0JSxcox8qlO0HlACDuFoKIbDCbkpBYzkoQI1J
sG4Zebkjyyvt0TVoH3UJQdouOkyvW8BhIoN8TUcPzDb8eJKWMi9aq+PSmQE4dppr
oTkLKIY/WNXih0LVhrKPdld4SDH4XGN/uhA2bCRV39zL1vb6lnN6EYfJrZB0SPvR
VFiAAFMb8bsAsGjfYNI3ZeM+IHuO3eo3/q2pf5IIFWh3N4bUHKG++l2d8Ssk5LJ/
BskEABZQoa06kfRWvzb9W2Ijs59U4b4thtuxtfsnzq/rYgnrP3+bN/kaZjCxeoiN
DgvEM2iUN46bsNXfnsRq9jsRjg1Xuhe3625ubFM53zwoTIMLwq0MMjm//TBYwIXW
HreBi9V88AZmL3l2apZDVL9/C3PB+idW5pj7xaxyiM9+QYMs+m6FOnEy2+alWBse
rOUewPgahfd22hzy1KhMW8JjpMbhIQvgbF9MyTkSNX0J0Z7x/0vAE91g4YXML13M
zmO+FDK0vaX7cSiCOyICbfhkEv/pUMFQrLdvbmNPa0/nK9dh1KELo2OIXvBXIZOP
cZPgyPnqgHHzNAAh2Seao76lgaSTh4lH2fNling/5QMduxV0ASmq647u/qG2X6Pb
5KiIWxJ4wKBAr8ivQG/i1SDcghNJRp3t2Kpnlf9YNJ7RNPU6UcWbzB1RYTHcVVwZ
PJ5KdmbOj02zgQnbX42vH0b2E4b1F1ZpahmF6Xc4bYzrjyOegko25CnsLeb2XzKV
9lY1mogoHIYeHW+vhtHQci8k5rWjLOUh2bJ5SXv5G6urE9/AXwKViYs4Fpqu9ZTV
sKXn+NJN4JUcoSYbbrDh9AUzK3538U+AU/pOB7punWcgEVoWLlLTYXiqlf9Om9dw
+obqvvy2klACFmcAePTTgiWYJMte1XV2Qc1wQRbF4VTWfNIRDcBHCfSYd+Rdz7vh
zK/PdKoGeTnJm5Z40y+lakFIilWlJpdQRXR9XUptId+RKPbLHFDiLWDhmR6c1rw1
dVW91kw0ya+SJ28BkOZpk6qGVkLY/ARuyQ5rnPtPnf0BD6QTpX/fKnVZwGKpwsxn
K6xeeD+f8bcXXIaux+gDlNUlzEbbFwokr4Drqj+3TCoCjXIEhds5ingEzVsqP/Nn
kEBQS9IF7ALoGPipJzwryN7ZBPlrmwC+Auzq5nJRl+acEQwsZL6swRo7e+f5qQ7B
AzXpFTdK95NEjnu1LRLtfgOI1AmIYvfHONBKsrhRCxP7mwcLtGnL6dnjnYyr1A7+
T97LmlCXsCEl3Y4+JibHIrKMg45MqHSFm/b8czUgV/ltUFwX6gU5a2oYZFW8EkED
v+Gu7z4Mg7cwMngE+zVuArAIBppfpOiOaXrwQpuG700VOTi05z66N6RfeZW0ohlk
DjdV6PONceyUjTRW4OojdtGGvRkhc+sp85ZSjVWTsRTisnE5uNPWkiaNgPG89MUD
sO5S39OqpLJGB3N9G39DTAw71dS9bDtR3cG7QVtSZwpcmeKgStvr2BaeouQi0cu2
lQBrbonQZnTUN70iEH68P+Uwb5lji7eqvlYfMa/IRHk3FDs7ApEITz7o+2/MAxiM
FD4z4STJK592nzEsBR8LgHH8adcvFpR8REuz1WQkbETUMZ/V/wqfIEobTGKRfn9X
fK3lW7nVUP8Lo1+Wyvm8aaSA0zaPFQIUQNyQt7DFNQqQ7KsblO5RLcYMQ7RU+Haa
JSoAI8WgRkseAE+1O7CcE00tMYs/wtQYOT1McDinE10g2B8Nqi+Uhpqvy6msEuph
DeaADLhHfXS6InXcYEUbWhJGzu1SDI+ME7OE4vMm0GKkLiq1uEIhdQ8ONCicb7Az
ibnZi6KQXtTinLmtK0/O4LMbJm4HlaJAVWJMVmHqbIcUaomThxGjVH2HcrRzUr3J
DH9rKrlNuasnXHsX9i63b6xKW4toj+QwmpJiAsZQFs6Po6kM+oJlUDKcpHIeFbWK
pSa9s1Ct6Z4xdfBCA7zfiMKRYinmZzTApt9b+Sh4p9Wd1UKoz3sAuFRGiQk64fLU
Xcp0+l7BA/Pru7iud3Tb/BGSSv2mW3EeERnVn0cvG33hqMLDMXOUTbCFkBpB8HUA
w0lT6fhyzH/T4cPYagtqQj3fgi9FPx5ECJpUdNouQ+eEP7RgjwwSF4Dut6ACn/E1
CIQYKj5wrJ6rkBwTcG/x5z00AcNjQ2FIjOjH/O/bC+THHNI40CFxwuz0Rs69WZUy
Hhblvyk5HNhfp5PCpk4otaX/Kkji7hVwqFj6zB/6GJuKTaD8K6vVWsShNtdxsd+X
oa6P4NrXBDbE/iuYKv2QQG4FAS9oj3gAs1STEr12TyBFk482+IwUgNBsmV3Huu74
Dj9QOpHTwbloUCueHUFns2UR8Z+Kr0ZmxBG5RB+OGh+k9KRvok/hiSsRH6veGt3m
ueh6SSg5/+Pc+UG52TBnMmGOGLbTSejDg17U/TWXbjZ+xCivGrK7+2SrZtsJ0YEh
DONVia5mguN9csiIr4DzUAv3lVZmWYDbmos+JYSAmNBgK5tRPJU/RBHNA96SOmKr
RRNDHebXuhDq7V/cLxi5helhSVnn9fMyhOcC0TvUXPXnrsPfWiQP/egmQuUSbPUs
9GSJqTz+e/6pdw+6xkxDIoGtKBZ+JeDyXZdWsQdbB4hMLfCiW4IWMV2Nf0B4qKtn
uv8HKSey7rfRBPwcbK0Q9OPiPc1AuM2hn0ubshEE3DVv8bDEZFosZetr9j2Wi/BV
RuV/ivPsDU8O0CtqXPOiZs+qJ1nji+59vTLi5WvmdOBiUCXITeFWENpsFgd9KFec
xSNFKXVp7ZXbeyWMqhvyd6anFzEg8DVKwf3qRfJfau/DWxcGpkkRq885ZyhL6VfH
P1r0+xy/lGsOtx8aMvyZoHmhoBoITGiNEQejxFYsSS1N7e7XGgN6cW/FXxFXp8Ky
n2DiAAWB+lDUIdyHkTnzW6RC44V4bm6TZGw6dTT1+72RkbfeRy29RiwBsuLUbZBz
mxJnLvhCmvcStXr0590Q94xDng2t98YwLRtF/C9kJwznc4V3WhGK5+nhHKtbKcN2
fJYPufx7MCfO9YQEVCzQg6cMuI01/uq1klL1O2mP2Qd1i3KxMDRFYkbPgztjxm95
1noyXAklXKslwolKF5ROzCrc0pRRO/Nyn/7LDf53Nb56BcKyFKFgVazytppVNzc4
RBCPnClolPMCdlPNGE8JbrUj73cjuq7cBlyKVyq4t1IuCRZurS8OVqa0jSADpUUY
uxhXEtf6geaWaY2LlDNKSaZr0G5vsBHvZCxvgd+DwuPYOtUpOv6s7SEj/FTohpCx
B04OQ8zrRYCfKbXI0+pDdMxsJOI1QLffKJbnOg7GdILDfeHWQg7cm7AUlTXtBAXc
dHD81DnPKwdU7Iq/sWJx5kz0TO2O7xuh6CJgizFRhZ+4H3jwlNQbYtv4Vvw/ufhz
yHxn4qrIEPwuBR8AkbBPbqh8LkWksotetG9t7hIZnnhGHMfiQXtjRODydDOZEZYJ
X5BqFuSo+iKAJg4wmch2Z+38gckcgCqFVjYG6OUHHbKi47moFq4eK87PMrvIcxbJ
TsPjnvHDV6YLnByLcqb8K59ciEZtThEnoAnNf+ILAk79ERV+45KaPHzD9B3OzbSf
O2gGRth0uW9NIyypq7jo4O+JOU5bHlJN4+AN374KjOMGp4DjGSXtWbT3HDpOR7yM
OE9xeWpmk4UqkyMDNOcvux+zRk7UNqu4o8nBPyw6UWccbbKqHA1CZS7RNEg6hnBS
iYqjCY4HaB2q2xEUGNxSaws4fE6yZjXc6wK91IPpZueoSnvxHdjD6amjV/BVE0z2
tErBYlgCC4QzrWP1cgug6LENcQCfqVC+w/023JkYGZjXI2xp7mNAh0GjzMgpdoOK
DlyNYV2MeRq51DA3wegy73bu74T+1kv5XveMzERuKfrSEuvWIgM6l2QtUwGM6yPX
RkuhDECyK8PL/uX68LZ4PEcZL2yLJsr/OqsR9ntkDt+FkCv0VpS3dBXNIs/BPeO7
0bZXcw/vg3X3I0jx/CD/M9t1mA1w0R4/jMuQ5NNGRMsaCv4pptCElVroH4kATzMe
Eh2ih0xUTaZX0dNzCmZr8Rn1oiM+oRUeO3xgsbcw00FOYFVOb624DuKAaq6xLLlH
hcDdyVmvRaG7vkBT+UlkE/quwwhiSMMjykiLxKukRK3Fk3ub726IP23buc2FPkkT
BL8xA3JfZKa2jZcDRfh8yTAwcSQK9sqeSfqYNNBDfaytWnZATJExYS6qYy3SKYvB
2qiy1vHjbY/8XyoBre7b3Yhjz13WMF+Dl00GVNMKE1yuvru5eSrSLSOewGNXbI+E
raBhRC0dHyl249k2PsKYDC6DnZRVjvE7M7lOFBHOMSEycNe1Rmryo35rdEy6nRkt
ydVz6dzSPD+eGBlYCcFPr8TgYDsHeGoVakVc6VzVbyvdfuq+Mt5djjP8XgcQZKgp
ubQGwzwaO+pvnZGOKomISxMdd9McynI0RHomxeEdhzbqzJqu+vekt0tTFA1mJSIK
pnl8VENYHHk2Icbzp2u1jjBDYC5bPtDtNLS6yq2t5Klq6I7vwc8QuydqJzojciAx
hlMjwkgV+oYgZNHDxDfDJRF491ShgPtcy55jjQUawwpeAC7HUdBthBUVEKWk6t1G
pC9K65XHyOre6DS4+KYzmZWlGOPnBxpSqsMqDoi3ykji+681jdzIqfL3I37rHc5v
o9xDktyLWzUknli5RwgC2sdEg+tE6pgn2XwKgaYgXFQpmcoOyCzb+iUa2LgGHEqb
GI21HUr6zwqluVJp9kudFx0Iw2SybxTrPAAyr1d8ZcIcqRS8eN0wkkRt6LpS8hZk
nidv/IjQu6T8BlOggM3HOTJ6+dUxmlFU2tMm9sJEz5AtNWSoshXcyPfHHlMqbCvm
RKF1m2wLbp821eE78w6lSWh4nvzBSVek92a/wOHi+h6X7ZPXDPovOOSV0oKOK5Ch
ZNozv3iKXoivbN17EbEgds35gKoxv36e2jCt2eANP1AXxxNau1Lgrjrg0LjoeOm/
f6qJwRWI2vVg3Xhn80hXA7ZRGE0nWNOzhmgUFHPiuCZEsvXy1QvzC0Kj4P4Fn8yz
JKcU+utW0nSrYbIZqqXcP9+eDl3PQQ/5GEkRi3Gp7FG7qUV+nYyEJVqooCVMnQ4z
JxSJ9lVf2NvMupKUiiouGeGLMVU+Niyxdp/jGHStfBPdjHHoRGOa7CEgjEf6XHjj
O9PQfmkqihv+KuHvKzqBGJxX1boL2xa55pZNqbFJucWSuSyUKv/Rerlre0AxpbNe
TX9XP7JpAk/TMNUbWYPOpasjhTMiQDLDCQlZtdM8UmYbhKTfV9PdjRzyzggpJp0J
gdkdVxMigmbvF47n0Qj6O31AwVwcE/v9ZrPL27gaZNwDadRfj4Uq9SUKW5VV8YH0
96z84vxMZIbg4INXZGrC9GjDgw9jnD+SqeWo1n2SVdJqOBBHm6Ml1oPcEVWEegWW
O9DmnytEphpW9/EuOsRbvz/ZfhRCyx2V+EVz67ALw/5z31yD+0hlEmoumOHKar+a
d7XPkDJFlxVMUctWJH3qlzP8z+W4skA3wk7bSCsqLxOnH8jCzh1xDMQDC5nHbCBC
EhvUxm9jhphM+1zGW8E9+Vwkdrd6M/t4MAhmU7CDEZrWm3LhhFLs/GqXDh4Qp8UD
NZZ16RYkFyk+fzYCsmteyHwoZRhDSXUgzPovQBi5+qeT6o3Ore1SXiz5ihhT/A8U
W7PpFRrEC3c9vxC17rCeQj716q++rKKTH5My/pnrHV7K0obvlkAHO9kZNs5baVIh
L7mIYer4+dZfbZQ5UOL/gASJkcYi/BbpiifCO4BZxzpzPXVOQqhOn3G7nmqSQBdo
peYWasIv7JQtl7LcP9MzYIwGV2wtpPiHClTK/Tsgu1o1S5q+JcFZJdyYIxcxAtKU
CALbU65XFBE+q1SxN1zht4qXfO0XqO5qUsyAZyIZK2Fazm93EPVjrh2NckX2PncB
dcXQhQs6k2SHZwAf8V++UleKDYDe2xSIhFSMBR2Aa+YZSPWni2KuMOogxj1ON4Rh
UkO31vKEZREMxzHEgVD7R0jkQ8QzcRPgA3F0alA7UFq+pA8zI03dyIvMF/tI/VwW
T5DVFXk26oeDKi8HmZtMkhOusOUzWWpogWTDFZyaLfuJPyvDMhRAkq+oNIZCQ9+L
E9DOdtNEGwalWiNep4zE0p+JxGJMbl+rPTkXowGb1BZpkf3j6ifsCYbWToHCbJj7
f075CDALclZxLswrjShsJdDJkA6h+iRaqFOLUm0k3wGKQLLyFxsJ9OwxeYUIFe+6
XNuuS8Yy7MuanG0Gx7x3A72lUYdos8ZMXFfhPwEPlUnYiZ5zsbKJH1/ZWBoMUEHX
hMH0dC/1lDabMggEz/CmH9OIcwkBoRdxin+yFHhgHR/koGUejjMuo7V17+n6Smsw
y0Oaryqhj3lAxaPxJamWiB3jbK5GC3cSXY4EuvE6HNTgUTwMUhpl7NK6fKNBjN4b
HjXFm5OwH/HvIc+IVDUs9REL9DyPtXNqFupNHcG7cugkwMyK9ScY/S2A5VTPzkNp
9TQI0c5xgBMb7z0T/djwwyshGk/SWFi8oO6EZ7s92HYzFqutGsuvC3qsWCNjX1ai
xpw764ThcTk6QsEJLrz6urVZrKzzZj3VEJfo8Wzdt7QLeLTDkHV5YaC3tguPTks7
LFBC+O8ZJoWhpPyfGJ0/QnPhj066TE9HfRksPQzBW6OQSHxm+NiDwZEThzc9f6QT
ukQgNPX8t1ZlxefiuWwpQj+4fTJvCzM4M+qgVMK3U7dd08h+J5fS6PHXPLwwUNyh
SKlKfrU6Z8V4/uBr7N/Ae280hrD/QDjT4tXRZrswZ651AdA6DhOjty2MdUngjDn+
Zzi9QDYEoFt3Gl8RnG0Z72JVMTVA6q0qKXLgLdtRvMaUoanQTyZk3zAVVxtTbnod
J3hvhDujH8aWR0MVP3i0djueo6aCCkIqGg5MuBqHZFACoDZAyjFi0ziO/ENmWsCE
Zzdc1kTFwjiyjGPU+Wqpxlw/J8j/immMSZsma6QmpmtXCwfJmLFqOnhV3vBrGH0V
XO68qz64XhiJrVPnkxdZL6mAdZgz4wig/vidraHrMer4E5rcH5ndbkPZL/5yOAEG
eL77hMmZTLQ39YS6+MZJqKxPM5u0rOkZCJ207kZmWDcKdAFlfexSYbzpO8zhPrPu
0EAa1K76wzbVuyk5PmbDhkaYKxGxQWdestCS0h8oI7ukfyVTu7mYl43h4EIGtgPO
wd+3ZsxGb00SrDxy/Ddbi/cuUK+JSqvooUiyrpF/uWfxZD+z5JNrxbOtjQRt242h
XuT5E8NK/mXR8QY5fi3/fID15efJVfm2dkqdTM4dGtem/hOAnc8K6DWljYMbzT4f
RUB2gyuyx/DDCFUogMjsfEFkwwcnhjWFCnnNuiA2yKBM3OoOFmjZwpnUBHIYaKnf
L2w42/ziRpBcGoVgv0tgLV7gRrSw9ui5JNnoNhupO9Lu4hCypyxxyaT5lCiFfSZD
4RhM7cF1J3FUatsU3PVNwcacBz1w/hPnsfb9a4d1h6vnvsDILs3+G5qEIPh2BLB7
Q83rN5GQppBH+wGYerz3iSrXvuHr64rfO63ArG9ekO0aOyMUGInVPC0wlomQh4Do
gpxTEdbArKKYPpjp4tkXSCoPATybqCfn7xoEHSlCKbQj6sZCRTyi8ohNZgbPzObs
LTapogpuZZI1WEf1hq3eZ5PfKAVR/5BfzYylc4THOHJIREtstJ0mCtjvUvbtYDsq
/gs2koHYtHK1O9P+HcCu4s6Qggl9VoToBIADV8Fa6e8fPTncvumgRIERtmwx856r
byOJCcWavknWhhKnspLJtCshZgFLHZNxD0Am6jlusmqOpEpXI8id+LyTkTap9uUj
WCiavewvnF4Qgow3p3sd0xH0wemFPRAo9TtoKD/xBzbo/uNtsRhsxDI2H3SkhjKb
TZrL2dPQi2jgWeaN1JN5ETOKbEQHyKQ8U3Zb5E5pa/ceduG78yEsKuErKn9TEJSR
S9KvdTrczzv762H3BhcpCQKEMmRwncyTd7K3jNZun9izEe5mWY2SXCwbEnT7uDM/
H+nljBBkprTRnzSwNBC8AnTPIZS7ZOKYWbcJ/c9hcuja6+bfzI75LLB1H9Z9YML4
G4DUvJn9m7qf04GGSqXjawkVyIpZqF+/qRgaHPyOxAIMH51TVj6pP7VIsPjavnhI
UbYNtiF0y5Bxdgaa8pGRZ51Hs1SHG7u8fBJnBQnI7fXn6SfXwZHdj2XyckOxSVC8
xYpa4O/znAAZroy9CD3HyEM4IUJjPfKg6tqvatLsx5lMtTk7QpBxcXeLTV/VZJkH
Ymd3kPjkWhe0gMovNFsrTO57gNxlxW7qRCEUFQ2atil1iforMXAK1G+mSZBOgNLJ
RxJjHywpKaMhTzuJMaJWg1IRb5Bl/6E6M5k4BqqBPcCngsa7HBWr6KL1JDo1yBo6
zv9B0QAF2cEOMQDl9qs9IV+PHQx7q+d0E0Aj1mUP1MxcD+yTYWg5bvwcoG83HM0p
f0hb1J9pqPFgbzkO2L1Wd6EMCl1TQSe08+Ef+mYBu4A5fBLCPRGTSXG+8C373Czm
PQqmPHPzypXInkHNuSjf/hXP0+FB79gcX0RVVnz8+fHYFDvXLkDpqES9OTMyH3Qk
5ZRhKWw+HfeoIxPJimUH9zVBpC9w/gsuOlKzukTIQqbe8NqQSqjfGm5VupljzcmQ
ykA8XzE+KF8BQjDjkZjig39YxG6HoViYI6Qv1uSRV711t7LD2Osvvgblhx0EooJL
C96ycpsYspK3H7T8cQ+qeHlROTLIK/T/fAXNXLWljIT6oOmOEA0aU3IdkqgPsM6h
BXNJmMEvKl2EJrbFRuuPaouwBbmH4V1rvMI+vkttJokeeNTe7npDQFjrro7dvZmV
6/moglTL3pUdPcMdaHJRFSRP2uwevDWMBxB1HKn6jdGKG4OidJ5bIXc6gX2c3R0n
5Zn6DWNXMxy0cWdzXjctogUD3s2GAQTY/FAhJfB0r0rdUllfEioK/pi0iaqZGsKe
Ej7JuMt2KtPXCW1/dnjXLHDA0/uIO6BwMHODDFX53DR+1e1FFGOEYchz1NXMoUwm
oFK6URjPl9qDQ/MHBxQ36b9nx+RsBNkmf+gXsF4JTtmop/0ZzOVyFKbgmHiL3sbQ
Z7lUhC1/WGySaiuFZyBsOfrpfqocw96QLUoXhWf2v20rlKYQa/bRKVO+9LKUbBHR
//AwiJPss+vxXNKFAMUIH0CihNHxoXZtMOGztXhXdU2nfQ8kdG1xMsn4YXAI+ioz
WXqmYPhmBxrVZz2o4PzdmyJ4Lo+lxiWPQ7XBHKj3+JY1FKbSbw+u5Q62gfYooHy/
28pZ/AHzO44GOPsrviKE3ZLPR12nv4PPLIOLVj+XymzL9cC7+4IBjhQ0V5ZnvohM
rx722QKZdeSKsVTGMrWAVxCoiXdegSM/go9ymT+xqHH5edIn2LBxE3LLSsEidNdo
50kjRY6t6qwFtXLZYTfWC4q+IfqvhLkCfc/gs4bR3sUyJu/elyw9TjfNVYfq6YkE
7e4G/OxTNA90pqfYM/bHCDnkW11i5hpm3TG75k18BBxHBqRjpg7kNEseBuDlNBo2
HB19+0kumMKJR3UvQ1Yt8J4NcsqQzGf6NJFLVeZH/6z/7GFL8lPiovYkQ3MWqQuN
snQKWjt5is8U627FtJ7GyPHTCdXE4mwi6vEZ96bU+8x7qE0o1oqRSQ6Mfao+MiG/
sy+Co+Xmx0G+2UDambNM3FqBhxRHxZ6Bte5pHPe4O3gu5i7I19ikYUtMXj8cRfSA
TiF2dqcyqViucGcX+QrfdwEqaKZ0RxE1eSzSTQn5KHp9OCT9vNVZQ+yupcHyUyvm
ALZ8iq7jqWDueNoaLtQQPnPrAFU/8/VuLA65dWVynwDW0isaZ+rJ7pc0B8F0ofmu
7qwJLuLLBVh0id0T8RmO/tESasfodKGWlQ8gFoaQIrCt916Ih5S2iphvjIRsoR2c
jYbu/r1wJ5+jy9iuTHxyRd/Q3coPvbH1zNTgv/caVvQGlPZjnJ0VcmWH3neydvY5
+zAR236xf/59NnqdxtG3iCiOps1bgZU1WCftRbZFG8hMqeRUIVQiGU/SkDYxfhAk
buqCdZWIXVAYyjzcB38S3x0IUZx2akeKzPbn3zn+VtCeEe7ijTgCXHJhPVmZiWuj
oblcgQq+T3ABvR8hzQSL3wiX/DLgNLbajxeQTvZonnQPCjmLa0MdVfsE8VJa26MP
DWfM6WAG64FmWCSpclhSmk4gwJ//gizDvKe1j3KoznGFcVW+ixgUGTQZ/sVdOfDH
awqf20CP+f2V+WohhKRMxcRpM5v5RPQIF+XIQ6/lIYcBpeSmFq+Nx9SavfI0ufGs
xOqnUTsgThNz9rCcTPKJPe9VSbCe0o18cWM6hZb4pkbKP5BwmJHg2mcqLlWZwaYz
1/1hyy+97nTJcU5IYTf59erHqQpmxA0IyssS2rLZAiV6G+inc6C72P4RS7JPB631
wQsNBCGKjnPtOedudHaTIGodeFprVzFenjAI+/6OAv3TIj78R6XHckhIPeaTFeuR
u6AY9m0YArxliznkAXqw0XCMgwXlHa66kmyaOpHP8Ef8p54BC6a0aDnAQI9A52te
tqeeaEZLn05r473eFqqwPU8wzNWGiN81cU7cNcJuzcXGUfYI704/UOQfCItH/hz+
zuFDQ/HyzM3GACozW0ty972SHkySmWIVJEwUUxKc8z+Z1TCkgA/+12K+iHylS07r
18dyssvZYC9ViE+o/koiMWU7i2JOTyq5WuP/CKCVne6jXWIlndzAMvR5K5aRpfcs
NEnLjWWBH5LYpMHv45GHd+TE4V5vJZvnfKhFXm69GyRg6fgr+0+3hYGEpoBDb3/n
c2bg6g0ek/ZE6x6rZ0rE+9DXRnNspn2ph79hkJNQTaI5u7++/FkAzob6+F1+6zWm
N0mEVu2j1VVGjlLp+s3pKwXewA/SGCBczXKI9ElLc7ViuB5YE4NaImDOBRZ/QaOv
zqMG/zieLN0GfJSVDojN1Dt20jIEVShUlmsCCv3v/eshHfEupxuMgFe8SmIOHTLg
RO6EiriH3jepSru5NfapXDRK8NVdJUVC8AZ2AqIRzwsBfSieJe4YQiNixSnaK48l
MfjfsSdpI1i4pCx4Ww5cUttsWBo/EMCyqQ6VyBc2Jn1SKLCEPDiIcEcv1LEVrBju
xuugDJQdNqhCCBn2XBCC6MOHvmpRjwvvN8wQWBRdREKIvAj+CbnraPmKAoaDY2sy
iMXNEIJc/1pNE76pOsbWC/416gz6MqBq8IznH4ObeEDAbVEQcOT2XRkAeN4sU6EO
EZjzvMw+5jp0/QrBlae6ZtCejw4CjtpstU1oJX4HaJaSQHPFSUMzrB1SQb1vIizY
oYkTUAegPira3qzLTccpj8QthgWfzCh7uo49AvWZxHksSwWB8cp3fsKo0Qldz0Sj
+6pfF1u1gYSYJYlF58F25TROwQ0uIl8DupUchkF7Atl7l6Vor/flhypOQmIvTEeQ
b9CzM0QQGjIeAL6xlguuqpcLgMk4mHoTNzsgy5SbC2Q9W9S3Q5ppzTc/uIL37+eK
195MFWg9+oGaIemocpRxCfLSnHU8Xa+o8ziXo/i+C79+nFkvEy23Zqyu0vg32EJ9
+trch/F2ktoWqJFm2ylxzF+3LAO+fNf2hIG8oJzvAA/vi9wGyUKVKJlJeEcC6Fgx
gjmez/0PVPMxkbE0lXtLRhKi9+GUTyu322Xs3e/MuNWLJHiMtdJLh05wr3EGmnoA
YgaNbqKH3cLe1Wci01bJbqpLoCVTNRetJw2S6D+/dEqahXi4Y2fbsy5w1Xr11R7D
URgw8ErWWiBWpCoXeYo48TQscvViu//eXoTAIGRDnDCEPgOV2iKYxns+TSFgJY+u
Udj9+3p/YlML4iAt/mZVZPSMfVX24gemF9cABTAjYt8EPwaaY+3XTIYLS4OWCKfl
sVqRh89whKQ6ttf+ve/gONbW6xIcVUVAc/PeecTKGbQngOG3Aqk+KMJ17qddYjXz
jJr56cMVh2U0OXGfPqvMlkww6hWoKDGF+ycMvTBScHsVrvrCowWpxTZ2ao8bOCrx
sBx0q37dwKdHaNz4lA3Vn0gknSR3uQBbi4oQ54vbxyJiiIWO1E2pijftbRTIHOsy
ffytfm0DcmKPHGQR9H5Pl2WTWBj849fiqcyH9UbO6WQoSZGUoXvA2XcpcsUbpUb+
AZRc6vJEVe0WqcReMjMfjJhzRv+6yb+PFZL/yDH27DLuHLxdYkT1VXs/aSMuqB0p
Alt8tcKhAWcZSp3hjvmTzeKN3vydVDDKxZWO9gzuP73L24CTK5MMBDnJxkEpDGQW
YqL1M14QRCrUymU41kH68pXcuzgeLQ61IVclL6iwOpSl1Q+Ep7kzCvkcP2EruSXE
cCuYEK9E46icdQMc8+YFCkDAN81PyO1erumpWLRgyREsijIG2urHBkx4b0YHs5II
qbZxmumfUjC2DsR76EnaiErsFqDjo6y1HdzDssvBWrhx3CYSC1zBjbyHkqcR+Yng
hl0wEV/h4tS7KccA2t9riozZtW5jOm3yHL5pfbRoYjgtSxVhSPoCV61hkgg9dR4a
eZs5OnX7X2LOx5FFC3m6rbDoER2Sr5jVwOCY1b4R314XoL6NqCR7G6wtnvMqipaI
KZHPguRfDAOCJMGKjmC91u7k+HS0ZaeY0ybpfj2qDoFtD8s7xEwReCpJ8Jho5f6l
7xl7oYwXFDPl2Q3eRLBCkOLZkn2QzOSboJaVqeaeaKG87U3jeXa+1VZa6sMX+7+L
oNVyya756CdWJa/Cikoqn0EfIJWwbXBAWOntMfuUkycB6jrsTIYL4xjPKETpL1Sc
s8LLvp7+84Et2Ysy12lkeQmQ40Rr1aCNrCLPqTdJYgPQf/XWCre2v8w/pVacpHpb
WKkanpWp8LNq/cbSTbF7W+t3SnAjEDdWw+rZCbi0/XQ0VMSeMLmROcAK+jdT+O3t
D4UgUS3MEmd3tyAtU52NMw2p/s3hHyVUHvMPwyeaGFV20LPqLPDz4x3JCR/wQ+91
T7rik55Xe3+L+cJg5ExYhK5dvke7tog7LDMl0xmhFLm9wVJvBASJr8AQvnE6IpYz
0l/pAVQippt9oq1mh8KOg9w+PV9QsGhr9Ik6ozC5g4WhJCE9HJA4snWOeLIvmq54
k2gZ0F38LXOzOzUB+IQYQ3nQ2cbyhbKhrZ4cCJmzJyEQyWTfk2TGp/4wR+6nULZp
uBHeQgW88VZ1yQYzKP3nvP00ETjx9b9uYl2A3BW+PL9KKRk+D1CVQpCUC8K50DZd
0rSpXzxEHBQf7gxYeb5CckHdgnyYaWebOgl4eGQQFD64rasD5ttJfbntF9oqs9SP
pMVu8qw3c3AHMMw+vNk7ohg58Gs0+og6PNzIi7m5MjTWT2p/ME5e1kh0qbiCJD5E
wU2igZ1WP/TfL3TgAc3S5NGmRsNMwbDPqrWcbJRhtCuW776KL6MOErmv46xt594+
fJFj7AiBuK/QmGj4uD5VPxu+U5K50fsej179tjfLr9OdT8Iabja4wvF5BAyDlo/m
/puZwEBuyuBBPG/sl2T8ocHBQO64agLSG0hMvhTQgB/l1nx0yzQmUfy/K/R9iMMj
X0zNZ0D2nVv0Qvx1DWtCKC22oM4PYNgDatID7XcgW2Jc+jkJiPyC3RjJevxSSrgD
5kkWIQK3s4QIvD7mKcLoi+3ZA1kEFa+5Z8/0GOVroT3VyMeRjvzrpL+8C3aXrSCD
+c4NAG9rJ9q0ZXiifg9G8amQ/UnIR29+FBP2x3PuunI9dJfAP/zb+rJWEa8EcZXC
oOIOLtHysoccho+tkv18vccNQuI2EXZf9NU1PtrWvxqf1lsXNSL94BCv/U1NY+UC
zZYdrni1frhhTpkS8FYDGjPZgBFqQB91MZQDrFR7iw0XALx4D9jB9GUSmUY270M5
b2Bz/COLO1c+wBUEjFz9o7GRZQZY8tLP2e5e4hktMxPR3ucwkUCZygIKRw4DQMY6
8patNpBnxve5VuCrDhzfJZxnVNchvn4Qye9K5i5bCJ4eI85vLsrFk2oM+fALr2yP
kxciyRAGlh59Jw2RBjuKH4gokll/3p3Dij51QhEnET5C9GXR+VhKNJVY+y2iMUMt
Krn8gKhQcZh6g5k+cab13yrsLtLlQGuM7CoXNnf9EsSdPcpfb2YYdrEVdlwT6V/P
SbxMKASxWUzq+RtwMVdldQCDHlZ2KTSyhh9gyXClwwt7EFW13x4XB06p2IdLK2RI
cvbCegY/+6B7J7Dqdalf3HB19YuD3+UNn5ybPDL3FqLnqSMHKuBUyMjS3/U/30mr
NMycTmupXEwqYUTn2c+3oWqQ3jbathq71TKyMb/o4o/EMzveO3u2Aw7+l5WL4J36
Rte15WOHDV/V1Ma9rLtNaJtkypl57ncfAhyOn/LOKoSEHVKT9mSQEgcGHo4ZiivE
Nk3/EL+Z4rkIxzXwf2cupoyMdcmoZ/sJyjsHGDTm0XevqSZI8bIE+Jtqui8R+1Q6
Ub2KDRLVu1AYwCXl9Et/M0bU+cs7tfvqdWsQ1Z89n7+4KoDyGQnXdHF/3vpsdRfb
1H+nrUZ/UrqoMmosY8gD44tTYUindG7XYq20/IX2kTQs1Xx1dO4h+tRd6tV+ZGzK
hGSvmOQ++NcZgb+SMavHXrnO/lwfGL7a70bh11b6IefhnkKl7lNL0DBjJQTQUFVt
iGb/AQtXFwqtY9r0d98xjF9MWq0w1BnB6ZjDxBNUPAF9OQVV02SURiM/Ermu0yMK
BkYQcWyh0YLDe9nQejIu0Jasr/Pj9rZR+A9RCWIfKshZHtSYOhlI4VX4BcFbLiyF
nTJKog/l9RYNnRkloPca/YBo8dwkjinMyPFMW+wsE89grGTxP0MUYdc1bPBm8yYJ
/KG5h4vlLEqFI8WNXLPpvqukDtzq3QamcvuxEgkLcgi0OPOp16Bkmd75biZ+Ij8B
/t9ap+7Nw08kXbE06h3sKzSstV4+u5pcohrBoFJnLkMF5pEbF524J1PuaifMmhYD
Isys3jHz7Ir0kv/nBWGVki+FfM0/ys10pXH2Vx96u/EbNOSoOmfqXab3IXahMhGe
vHhVqpE8CvRc6mz4W6NraRTYtgzdzb5kvHUj9Q2QLdW09dLzcBr8Hx6Jyk+/jC/Z
GP6F3yJh+4gITSq6SeplLKEL2G3rsmN42KnEz7IDpLBRCk8m6bo5Zq3qqpYjU1bg
niZ67um/a5EDZa6y2g0yTI4vLsholKUh9QrsaPLxA/sKuKcJc2bDeW+9QeczBvnd
I1zgbQVzOm2wVBiJQF2fBx1PyKX1bC9auSRGAKsl8qlhEGN/GJ2GVWoBVL4OKuJH
Nyd3KVE7fvsiPTI2IDWm93be4ZVw14NgGkMkZfOJaxTzGsM8L/LDRNUThIOTY+u8
dHVITcedoEr2eSVBoWxkQR9aQDoJ5lQeiPxiwHoRFX/Nx8p5fZ74meA8xcD2QISI
3aTyEUjro4SmjESFw1wUWu/bl5wKa67wsJ4eutnbqNbrt/GVvL+Gzxojh/10I/VH
7Hd2EP4xqTz0RGjSJU5VDu6AnSLViRWnuicMtVkUdAjstFvbWBVF6K16sz6K8SSv
8OVkAF55eSLUUAhA3pqsJU9fZ7M6prGYtvoYDw4zIYW61lRRrAqwpO4ObJSLXanX
Iy1rGcQbeT56TgIdQGWeDlxhMAwB/jodnmidCS/GZL1Xhm4LXlo2rFCj1SU208cs
uQyTHYKEejWEgJ1vgXGltM9PBheUstoxC/nIs7ubH5GEEoQe3kilIMQeISQbfzOC
rVjDcX7+kf0sGq3itvCwr2RLm4rmvdo8uH0uA1PmZOKC2j/4TaxHQQhDZVw83kK0
GZRda//B+kUcH1i4ZrGoUKVv+4d7G97Ae7pM4Gb23f1KtTQvk9y9ykgw1OCv3YKe
E8sm00GWZmzfptitfXDw1B83wgKiqesZSXyrYmuBhKzr0GDALv/du3m4qEX/y/sg
YK0QxgjEhNM+na/4jSFdakmRutOS4V6yqW1ahPdxKI5rPXDIdVraudDAbG7dChyb
RNFY2iyHagoxQT8eXQDGc/3hGgE6J4z1+YchcvfU3E3dY6NpBi2pV2T+gRgto6cR
3i6OhD7vSXxox93lZByyUYplcnjTwM3T8ADiufahWQ5Uz1q/uVSvZcaAnTZScOJd
sds9wwNXcXDCSBOjiDJpn35jAB83/NykZ8073C6XPwCl/i54AmN8G6jZsgYcqGGJ
RgcsDcuYqrzdonOjyHEwsayf+uIctbsbSriwwMg241tL+R9N+dsj8I485WYqeIU/
lW01yaEibBimFv1Pz6JOZeBvBN9WiH1RZZ9ybwBePLqKjr0TK2KP4ioCX6EFE1wm
5oe63Ap91Arij1uZZKlINuc/5LKDaUX/ITXJd0t30FiFvjTMFz2XfqMurgQZoxY/
kCjsS6KTQZVWcxS3T+pX0YL3qqlhcM3kFimJ2hPqsQOgnzOxawSUnw+0kdtgKzwD
PHtAe/4UXjWd49Mp0aQrS+mblnRi4K2RcGIjihOyUDeidQnB3qjbqeyd1ShenkKG
sFUxOQbaam3w6yUePTso/2KFk0+x1ToxMBcWLsyMQlgkj5qdCw9vHkkHJP1w3Xwk
2grCwoan8F2DMfhWoVS1fLYhylmaDe3H9xTS7qo4u08C9vyT3zU2fH1ss0l/mD3Y
PsJ4xOaqZAMWgZSHIAzuNvsi0Xh4L5M9/SnBmSMlC8CzrhPYOCd8/uOx2MAiIsp5
nOY+1TKWw/RWKfVrjhTC9mCmIEFih5QJebmuYVi87oNs4D6cSA6zjf7UhUTSLfjV
9wLbZb8Q9tCTwikMrZza0I3OnHG+1xQkr+FZeUdSbOKYTPZl/BRaKJnfT3HSZpSE
ZoJaECcfo/miak4Aao8WsVL+K9LdbDNUdGoIy0SUu/X7tDKosi3I5ss3F9EIMtuU
ztvq+asJ3dQMtcyWd36TDN0FKGfMGes/VCDa1/zgBfQhY+kHof8V4NVlFpprC5qe
4fMk7JVQTSg1vn0+dNqQtc/HcDDipQ95LjIkdtBFH/FHT2+CJwkztiNKs04EEuWL
NFHTOd97zgsfGgOMhYSmRWETDfS9zJrbCIZeQUVW6YIuXKfA4odYkVgJlQIO1WDo
6PLHF0/XTCndTmjxn3Z5MgGgLZ85gtn8oINY5kOEHGgnWNmBDn8f8bncdC176wZc
p6+sw4COsjUA5nBzZNHtfLIVSK7aaiKeVuivPuw4lwMMdf9HlaPZyiKsdcPM9e7l
lX2j5UWYiT+1E/qanLzsOdGMGeglZvUOb2kChfJDs13XUAAR9HSPEyqKscOspbeJ
wDKv7mrZeQY1gWGQ7pZuQ/7RzFVPh0NRlpxS/h06UEvUgKwP98GrcrboIOmhquOM
XJ6OUCpP4EJ6A8x3DpNVmGOch4zfPiFPoXA9emGFTgyVdPChorcOY5QMx3tAjick
gGO9ED8C6CX2Ctu/TGtlhnlbppebMmVPictzM+3gp3Z/dd6BqkKPcjMKOr5Hqzz5
G7I3f7M+UtV558TcHG0TcujczH3ByTsNBFXxpf/kMYmbEgcrlha7MRaBGHiyDbWb
FJmFlSRJzc3S/I77QZhgEH/MpredLwgJ7Q8hGqiapo2OAZWpfof5xWfigUAlKuBf
o8G1EiOrLUsNOQn4wu0SHE6DsFQXg1AOSaMhaCHjKVYPPQJod+UhMvY5gJpbnOLm
qeAs+SAe4ro3jFNj40QHqH4sZoarA3RJnS2iEvcOGC53R/w+CRzKKIscB2ulZ8x+
hE4VU9QxfsQOCU9izt1eYXF+LpDbi+FjmYVF5A0rEwPzNgIa/lZbWvN3g7Lh1v1N
NqolxvkN9NtRawnzQ5UaB0Cp7lJMWC426dyyOsnOeyJ1/kv9h62hdWxxfqI3Svp+
3rJ35vJepiDoYS8/F2ekCGKUCprHbVqdMhjoeALCIk44MEl1cYpJ0LUm6JTw/RDS
M6gCfKgeMSVPqiVUyCMpEN1fAlKC+qZ6+v20RJvVqhpt/jvRQdHR2lu4vIU5YQ/M
wQ7PzStBWI1qhx87otBco8clCLECTV/lRR9Mvlx51A+zevqqfoS3WNR0Szj+KX4u
B43V/Qbp1a/8QS1wpGKmLTvgUTPu0qK2Nr4YcSfX5QyN3x/IEBqTxSrMQcxoruhP
HeKdYH4munNpr5zgW8DXSKHlxjgdXkRhZ9AnftEcWQwA9ZVy3j2ywPMRF2jl/ywL
MxWuDkKiUnYcu5/34juyXF7XCQpw4SRpX11LfBsLpuHHf2EvNdaG3qC73J6TyKf/
rMI1zqJdcBB6kMGIlsGwtledjQYJfQjnU5dpo4xJQOCj1F1FcE7kQ16IBFrP6su+
umCspCWjOMg6B/2ch2Joyo+M943NKDOw2hAY9f5EYNetvSfe7qv99u2I9dH7eD01
BfKJLLcIn6Wb1ybzK1BdLyXqm/mPRxyW5dsntZX8lID6HbymE0fI0zDQJEF8Qf/d
KRi4Kbqfm+UK+bJ1a9d8zH2bio1fiCafP+MCm90z8OJVWp/NDHQTJE/f3m5vPVfC
PaLYnffFVApIZhflGXxU2Lj2QmCRD7FuRNNxx0feh09PWJuEU2TR8trE0eKGKYdJ
lHXuEHa+Y7Hr39SR8dhpdcZ2VZz2yKURaz9RtWnjIHa/pVfvjPyU7j/Kb/LujZXI
6mCZ4uCGGEkp2+bsegcOR50tLz+Hx2YKuhwSX9ReLr7rm5rRxqWwjfvGkH/w1NAT
g/W0mrAphDGxniLuFrzxA2dr6KE3Hz6Du6Z6h/8gnwFasCAcgrvouRnyz/5hf10J
fBUVlhxWk4T9pJEFFrHdAAGQe/GB9+ULt8AkP/5BUtnYy6PPZVHSj7CAzgg0TVn4
xZuwc6Jq5SPXOsambnpvlaRRWTxvhp2+4v7trN5YcOs9ZTnZKYDGzVUFwgyua/Ye
+KClv9yY/mJqppUxZ0OPJ0vNvR6Y/MgjQ66Pk9pSCJYs5a7vuVFX8QtJhsRcNPNW
00gpfiaboa712kMuHzmZnbG9fKj4taCikBRGt0ZqaZ7P2QMV11QatTuZ4fSV+JyD
trHFPo7TcqkhVrCBsqmfl/juFMJg7z+7wN7fnZtcN+YrkCDgsvrQ+IQszWfgKx9t
bxGB8iCODmdjphhPC0LkNijfDJj5VbEAl3FJmKsM9d58ujbxEJbvLM7YF0xPs9ig
cJ8nmszglklMR/2tx9K2bc8t4FypUw0UwQpqqt6FAK3ApYeD1QuegYLYN3O4VfFq
D4YQ611xjfCX6sHfYHm2ikfg5HG3fk7l8TvAGRDUIBuYvLTXjHUIqTCZXWJBBsiX
T1GsPKMHTgGpytiq2jtUWHKxo3xIxHGSQQ8Tm+QkXkZDTabRO6LPBfkVkq4RyEWB
CnssYt1OYisaMnZhfiYf3YVzv1U4LqtCLwKf4mZa+XwMQoCfFbXLo1UMiJgSn2OU
n41g/jRbhmnPTXqSqmilqV+1KRbcLxTucEdZdF+0HG1pgEIBw20C1stIdrVLxaj1
eNClRzQlFuR8xNALwu7cCGW84FXxwJn8/9elhPt/LLGrknaERkCICbtTc86P4OE6
7KlvBwkb9s9mJ4wQWGjgpk6uFbtHml+EWPalNR/7FwCHZG2YRGxzPpB62qRtc9Yc
vkD1oQdALrU/IXQjT5HYFvL5msgszyv+zpWIVuYrAzbAZVSpTK7r54ZD7eZ/Kn4W
xIOwDhM+uMxZHabbeoZcprTevAxZupWZh4SzO0mpgirps/jt+xOTScBdXp5mCbHP
pl0lFUnu0nAQD44FQtkuhfrsezdZRq5yiNpS4vuCbCqJm9+YoldXTCpTxntzkTXA
m3d9IZ9qs7BihKa4rBZpUAX0DiwwTMLAUurx0IXRWwEP8lDtrRfsHrAPmziUjV0v
pr4KWfM8TVDzxxtcEr+GU9lvTYiT9oOF8Gi66n/Li7nbsSgZF8QNYrKGQRC/B97b
Ajx/RpS8dhCk4/yUYfOCD6Gg7Alm4SAmEUTTOypT5EnpTzKPHisvymU75N766VPR
NojMPg6bmN3AAq5cvqQ8+kpxWwEP29+8024ofTbhXtRAi5WKP73x9ZFgLDJ8myHU
0ekgpJfKZ0360E67I6m+OGf5CLbbuPdWBSWaF9NsLdc9W6Q5m6BVPZ51OEoOgVIP
Ycsz6yuxhYGWD+8a8/8Y8ZZsxft2jYmbX8uc+HxAm/SHT7pI0NSa5lgsg+XEW6b0
Ikb+kDzes0MVmhR2zkKmlNpyvMClXpFOH7Hyz0gmvUXePNmqIq9CcVQ47jCTfd0w
bf9hvLdSNgrsJgdlhKGPq/K7mQ4Y2+WxCH/O1W/UVtyn8lazjFwO2e1UKpYo3GLf
ZRmWX9fA7taVPRnN6g/yNHe1fLnvfmOh81aHbVpfsG763aAF5jJY2NdJT4CcYP1n
onqZdFsYu6UD5uQwAa4mqly4siqMQeupuFklT1Wi2dSXS9bH7Qz+pIxcaHLZzIii
1rxCljtr+0OJfLSWKKgrQ+4Ms8W8lRAW0o/A/L91YI3figjTFemBGBO01gBgzFZ5
WaXt1Qe7CvWwoGna6yA+q20cYPcAKfyo5WmSb2bKRckcp/N8kVISsntgblPdiG14
9wzilaDKzUNyljSgsUVij9IsQ6N1jtBeEFyslgOIRTxVo/i9ZoZhC7+eBl3+XgmO
TV6ULegobIvSYxg5fEOIFCdzydMgblGVgFKVNkAcclmbBOr8b111X+9kgBktQVcE
PoPz/2OzxxNpqsn0oJX39sMFMhwLebZc5jLOOqqZZJ3kMreMx6FcWmXapl1E3Rpx
xvunKQoP/FfoCnO6X8QDr3s3xVE2bu064Rsc4HBX4y3V9GGucAHhIJWLgyeO1xEU
NMHtaJ74rKcaFEsg6QYlLGFZT+P4Q2HRAmNqIfqbyJTqhZW1pVtgnS0yxP9nCjV/
t3N2S9bsvA+rFTPdm9xY6LW+3jgbiyD6REFjWM2PJ+T3Tkew1MoZjpIdHYlgLQNU
/zHJ8kMpD3XCwcRZA3tHk4UHOo5d94bB3rduOTbeHmz1K0nzTuoS9AKRi9TjBCCw
8M4B/TsYj/86qRNzhboYf3VvJnRKeJS6Jx9FfdeOqqLmB51D4hl4lYMmD7CoZ++R
Vgx4BGYih8X5TwRXMWKWLCvkuu3RiNu2rQ8gznwI7YDtP883Tk2tglzI8lMGUorm
LfaIVVupkDdtkeihjL8pATJdcAz6M1eznD+pfTRB6Lt000n0hT5g9Fx/Rgt55OvN
7vGTMt6sDbyG1gf6tiySurtaaKJzoKvIl0822aHizLEuOj4ZaRNZBxZyxWNB7Fyr
NV8DH5jxFZR/ArOTmtckiI2qIBIt/5VCUDQbp952G7iwSA0hrJrp/nqmMule6cN8
SUHiUuYKcu3URTvXawkfpGSX4mEDPnCMQYWlYRboywYzTtWjZ//gXahM6nq5nwqH
5SLpZDjxi3Uza3PUHfLUzl/6hnQzXbjWl4pOLXOoiIOCTg0vlYrPNTtqSU4Jdhxg
rmrbP+GAzgPcXfzazyLvpLSMILqUw37ho8IC2mXcGJ5nWABZp1WDWi3q5w+02fh/
cSYGv5NW8C5A9Boa37nzEuVp4umz+cJ2kYTMEYMmqsA+QEmJEyYQAmuF7YjkOpwd
TdwqnCqeQST4W0+FRBP5GrXHhoQKuyk65PXqgZtTbKOZz+adyTrwUm975allBihG
niJmVn8IkR0ELTTADeIdDzY4VLElZiWZEzBqVuMFzNWwvWgoX78AuiuPcGs6v20h
20LFuJGYl7eAszjQkjEQNhsPunZsbTpVTw3CusxHFRBtsL2jIP47DKJtFY+uPIGv
2YaLEVFUihF9mxwaBBmqvdftKjQx+iNSiJRXjJjaao5CPOLmBhcbAwHTmJDBmMn1
4wWTh6/Cvrc3Etcap2YHkJdJXG492QMOifwFEq7tQZ1YBR6p19YUWDU1TYlGgq3d
EoJEiwWxbKBlNQWtlWv9kGWBoP+pbB5Hu4/01U2gBPcyqU1e4CNWfWlPkKk2LygY
+UrkK4nI00e5UeOOC+ji26qBHGxNNgT/wIBaLHoN969ODZqwgV4A21SUyUbtCABz
Xxp9rhYWJMJq4ZjfUZpdCnVKtiO/VU1mpBEksNyi0czJhZl9F+5BwXyscFW962Cl
Rp8ShV/Y4qYN6nCsb6NK+GJ4w4uSdFuwSdg12+OlEz4MQkHp7uuhLCeWKXqvfbzo
/B6LXe42uYHMhdeifI5M/DjK1dtPzo+5JTfm6elNFE4TbfK7w7l5Vc83KBJrN9j0
mKWtlT0hN4lX9bMy2fldObBNKzykwIbPo5LIKfuu5VnaITeFxLtaD10s5qQ7yYfK
K268+muk51PgY7jfXHIEWOPySmsjkSosV8G1vtXZdSnxuawuLB8uIlaXKJYTYN+k
GP4FCgG4tJneXsM+jja/1riLMYc1vzMSH7HyzwTFcyWUeRbCH4QyADybIWpkgbft
gwG98TPX0isFYFgpQoeWSLxk25rICUIGwGRbkt2hIDquoHQH/s881MUDjgPJ4trL
8zONWl2mVfUhONBykN6WCwvFjr6wHNF4XriIilJ5+R2ZRJ4rnegwtGNsoiHHQBLz
QQKiU2w/H/S+y5HaLllfhUHt+S8ZadzJDlKoSPoijxvw/XJBdrTQ2KcroThNM0lm
h3Z0/NcCwGCHuKgKgoSoRm61Tt/rrSUyXakcB/Qc5D8kvF8xeNwLoGCXrRUz4KzU
GOGnGdF+ZfSIOb+PkMrLAHWcGK0sBHtq9FDBD7wittOvByoQzaAXGglvSbyiu8EN
J/rOmZ85sHHSZD8RyQ9c/7dqH8xmrUXIuB0iCL8QdMSqS49nHfIC2+XzHA14B2gn
pkXIP2iCfru1xH7urPRSKn7KBYbnO8kG/4DyCb9PGx6+qAJcaMH8DqqZb/TOxlIc
Qe5XxV0EQ0/iIu+3BpwN0zXBfSGmiH7v4wdITBV8IxE55wQcgExoRpTp2bZd3bPN
nlYxcgPMK1ec2Vi5HsetS7JvtSj+A/jDQfZLmCmh6RhbSrmHn6hLTxQtyAFiVWBE
HTMsusS5Jy6Ivk/DjknzY1xKxPK4ErXc9V+XrGWSiqY5fSwkLvPlqPfE6+WgsDDY
ZETAhffDyDmgJyylwyatgD6pgcJKei4w8VRdk2VTXeJhOwKQ34rJOQ3A9D9K5X1I
4jkHLNHTu276r+u7ZjFVg/ngS7dOjWk60GSY5mgjejnHr9PhPZorsWuIIYqq9ChL
mBcEmoJgTa+2ttcs7X8X32hUE796SV5A9BH5WzXLuIQqKDh0RH267GsjvHjIYOIX
7oqcF5KMkDEaoU7dal8SZB2mHZpuy0l3bEN3dWkpeP+kUtVldz62/FqeXZrk4i4w
J1Tg95RZQP94LDNReFgAuDtJUs88hz4qyvy4YmgQN6Q4PGzIVTHNsGRkQU+4h5SL
cQsRMxcOEBfSHAzpGTEQi6ApYkQGRFZ/Jc2qB2QScEs/sGSv4qNvMSkNGdEMIaPz
AKYkH4POuWqamStlc4YHNtzGyO7dimtmIRvsgrO6PSeMNy5HYzLOOYNRrFSOV+03
fTup0kQbOd0LbsStsiUL14VkL9vPLGnMNb/aYqFshSfZ8p42NUu5niCZWcQOkmeY
m7yY6kjw0lsjdKIJBpUWR+cpv54MZhoaC96P2hzQ9x5cv3wCxzHEU1m5EE5SbRj9
BLKRQ8ciBtbdu0UpUcSnKZtsSjwV5KRsjUVPIv1Xi6DbHm3f/HW610WH9fSn1Clb
qGjnQ6KAETSw6iOqNM2OAdk2UoHgQey+prj2Vo8awnbt6XTEChZWSGuV1O6QB+5K
DgHqi53MluW4yjtJ348EAbb1omx6O9E9UC385x/2XTaGoPrDiiPJ6DCtRyCAaCYz
kRMFLnfLfDoEEwcTqxW4lCnTKBs4n9BTfbFe6Y/0MwKgfXJSmdO73gF4bLjCHYsV
ajS0A9jRm/cq618BZ0ZlDhcnqNASTlLBb4KTO2WNR+5zRb7wuzTqaFS60XVVoH+D
IkOwh0mEzaOEMkugSbiy2IytLk727xOu8kA+hNQ43xSCw3ASxY/H0Eo1OxZWHJdQ
zR8/HCe2SDFvZI99+UkCdIqtQ9zfInLJe9fgpt0mNIJUx05qkTtlJA4KDS53LaiA
wpf+rjyF4oNpFne2HNTV78frYEOZRz0wnMWVgh4AtS+m4hygTT5QusHFAtMRP1Ay
pCYJm+MU3AXx0F8qR8V6EZnXQBpjZ6KbMoyhKBasIpS7l9m7/KLFGnh5tRrctDfy
6eLZ1LPG0qQbNu9mgVMFSBAs27Xgez5vrL1Ml0+bDmE27KU+nz5aPUSK7GqgYmQy
SksiMMAtHLG7ac8+B3KyXiGM9onOWH6YPgENEBzZVCZxAKDn4aVYwrW+xZW89F12
cKl/CQxN2K7LIMGQp25vJJckr/OVw5pH6IxTvAg/rqXV+4MKZxWS16xjZWdHYtyx
pvZFAX/YhaQUOfQH1TGu50l3jCp5Mi6E7rqyKRvSAHwpDBPbY5+wh6xOFBvaK82H
DDAJz3feWekygAO5dy7FBNSiMNQb6bzz+zJxKD+kJrEBjEjHxILAnV8Rek5+uYf1
JcfS76/p54yqmdzQlEsf38lK6eTcpN+zn4NQHAHDuwLNiviuO54gx7hfVvgxj1pD
k5T7lxhCYK2PR73oJX75nGx9XfKgoPjliizTUrSnDP4LWmhgC5ZeKL7q5IfURK4i
Rs2A3I0OXmu7eVDbKm9lnPMiazDzi4UpOp0OYLuOFR2MiDq57jEDGZDy3Rq654s3
6XSTNByQNBU63VbQXSOet1ywWwgffLDgzyYaEaqsoyvzcF9i9tUtsItHV7SFRG1t
1aJ6icFKh/TWVixf3W5v54avcqfAhAc73RtrWJE15JxBmoM0A+/lPgkGT+3gVmI0
srfGmolGeDmYV2sN+z86nzgbMuf/DLqsEyIEuTTPK/Kodz6nWraXz7czcICUI5XW
GSi1cO+qOGhMDf0yD6bu2UwcA6FaMfljBvuxtvUDqV+Xu5e7YA7KKduCqxkTLUYP
oyWs/HMlAhKw+yWOkwF9zRx0yzrj3fWsvy9Kw8Fqpmu0Cg5Q1XHAfagrvx6Yo18A
6gU5eeE6aQqe8F7pUOP8Mgy5HbD+4J8oJRVBUab1/H5d7HmzB9x9e9pqDzJbZccU
h/q0V6rp+VV0dHsxZzF9EUUbDiBuDEZHWSzyI6OUHQ8s36Hn476LyLS3eqHQXtDz
IKAY1VC3G9sNFP6qvehUOJdf8oMUFDXpouMBhF68QDrbggsvkFeBgEEFBeneMJbH
tc1uMWgbtCgdjhesI754falM7nRqUMCPSc2jbUTJsfjz5Q9dtUNJAo09m5X+Mj9D
M1/mhJGAjT/JyJO5ht92xOka8wZ3iUH8o/z+DFE71OdKrfL50yc7zkCZc6CyJbS2
UFOicD+9OAGyOnoY58rqpqC3r4DFyV/x895PT7u4pjAacg16L3zqoah7FN1gl97L
1awBVqB1oI8k0YYmsQvBu8/G9nhjsO/kj96GLiIL2mPfYN5q4658yvrwWNp6Tx97
MOIrD3KoJ5VnYE9NcIBzHcYI3ASKgWKLLSvlxuiduuB6Cw5BkXIPEUvuG1kM4cDr
JsGTOr2eOWSnsaxUbvkdAuCpZb9+e6BrhwR4kDhasGJIn9PlyOTm+x5D0WfVHNeQ
C7hmFbbd9xRwYx4Rl6pG5W8dSitgY6Lj2creYbVt8vCaoSy0p7QLqoO261M6/RT6
6Z6gNCixdxMtJutPJiUd/YFfe0EzrakPCr66UPZ26lEUc4vYuvmvVleLyuMkBavs
4xg8XjIy8iT9unusUOG+NODf459si/g90RAY3g47PzHUt8BPy5CkeGX376hbIxub
R/9dN67kmZeHu260Gkf5RXGOKMAr4ylLqa3vvuOEmg217bZIP+wqLelDEZ/Yz004
gLGl/5fnsqStOD1Fx2jVWaDhci296MpueUFJ1tHK6U5yjCF+E+7hs72sN2EvkCJ9
bFdqkTEGJ75ut4AXfAF7uQpHEdTXwTp/oH9UQqj/Gv2PX/SZjVD8sPrJ4pSEAw8X
sN+FDYDclkEHfWgaITfh/dVN/EX/8Hmeq737L+68Ey8yfHlUMALk2f+2Y2J30IV+
W4TQN5XWeRegSS3U2bOej/0jpLuve6EWHoGr49p/y0gFH3pRCZ075uuN1qgp2YIg
l53jZOMGMBuidH9e/tzpIGAkAeb6h5DRJD0AlNQKxDjgSMHv7L2lNlnE27D+0nKk
Q1C5nvYm/EAlZqI9Co7EFXSekGv3WA1In1mv4O3fZkSA2mGNqgjgsKfiS1pBayyh
rQx6JTkztKdUo/ZBzrrzgoS6+taN1IH5cH9Npo46AnR/rtVIePs2/DUW0UrzrauO
InCaEbm/cryofZRlyepUfWDir2fw/H8EvYQpdgrU8ds2XdTQxCy5UuJj0B3C/bno
2XQPgVsnz0K1tNz1s1XHA1fBy+IUUSqFl/SjIXjBT5fR0vNGaJjCuCfRU+70eiyj
LEF6eS+6Mcy+CoPdemxpKQTE83Ee5CamIXM/03xyz/KXBrmcpd6l99HSojwvEUb7
CIOY3Ab/6GUUBwe6Mu0H9B9i1FGcFcD5Wj5dqi6uAUfL96wngB3nZTrlwVCaM05V
RaSzxmH7TdgwfGNgG0u7m9+HtRjZJhXS6OvslSTSUrOUKecI8TDPgSjOD8EFJEN6
rE5yygfGKvH7D2fk1hQf7ZMr6ZIqwlt+9YKIfygeVD40OQs2/D3ItUMO42q1NSWv
BnH58AdwM0k8Nd933cJap3qn5MHy/6+FgE2liPxo4iGfgXM7BlqqGur1W9SJ3T0A
qG+a7RpN+eSLkhb9cVjGXRcGO9Imb85KXTwlWW0HZAru47NSw55WIxN+dD64kp2X
YYtV8DIXkK+7ct5AxRnmmud78ggSAIqSMl0BF9kLjHoV28VlmOkiKkANL6JCFNLe
FKhVEUoxjsxm6IzqiOzN6b0fSAynbnh58GecCHShhoj+Hv9N2//ugl+XN0mlpF02
mpf29f6dhTS48M1d+x1NermaUE/yKlSdmmcuSUdxFXU48EyPI8K3poR9dVXGnQ+U
I3XQF5/DQ1fADSVHqGkHaP43BMCOUNC3c2NEkH71Z+WfjNk/yM7sNgV5OHqG4oEw
OdV4sjln++nzw6VXjJUHkhuPJ2B5ugR1B/wIVv583NXZUmf9uWaixk1VAvJQWjR4
WY9m4EeNBANx5uCoWG2yw0dc8cxvAS4cr1cyb7OwF7iLYAIzFC9uaJpD0yej77Bk
kF3moLuE7EzTsQQZtzlL9opBecQPxDwLhMxNFewZrIY5YheqzwVzLY/GywA20Ahh
vhr+fzLUbMh9x1Ubjw0qYTv3L8CUEQE7X4gOQTmhl0K/sRom7qoS8p97gg0w5/Qy
yzk7Gg4DK89mDfYdjAS7Abvj3AL4IhIuCcrKGppwlIsDbhGge5vLX02ekJ+4lgiH
vPITSBf8+HoE5aTAsQECrNIjxBP6XqlAHFDtvCytbQrZO2h1AG86QuqBHJccppKR
RovGjRcPVbVMk5vYZf4WvxkZgKB74lWBI/TKtb2Pb3fp/KxaxhnbmRAz45/HTkDn
3tv0p62IVuMyuZfXL16xjeOsNaenOq/bd/n+tKU15tDMgiJYEO4H2FCNnqTpdOXF
qxamgtj3xE+ZKUBtmNMve9S3tzSvX7SbDn8bLKvlRoC19KEh1Tc5+c0hw6Qcrlxj
ZgtE+PJzDwDWWu61SL+Pymuf7MuyW5Pwy5PLsBxh+itkI/yNzQ34BIHHo65OIWxN
vwHQSVN3aMAnJEQ2xud43q1UUpq+vGfKdNG4qrw3TQXf8tOQhfJ4KpfPVosC+zHu
xREswZAQ3zlsqJDyqIJKTPs9pX+S1ANCC6UkFR0HZuRewsiM3lITug1+TVszWLok
YoFq1/ewUGwYoHqFAemzVx2B4h580hjJ80u3hSl84ddpWvYnycI0DH7jTiTM/NPi
hmugmd032GawHwQJk6wfRs+Bchlh4m6N3EojPjlDVLhRTjqNOjUCuHD0Wb9d9kO4
wMBhufc0v+JHIdR/xFCbpj/RP+14x46jXu32KC+za6AKnBHzdbzPjEjyntbOvVih
fTrHt/0f6wd/0uKkGsRk0a5sBCbKmXPA4n3alhMd/jRklzsfwGNgBfm5A0ct9yCi
wvf4QXz+Kt9jQl92pq7ZL/TkYG4XHWSoTCeTyq9tdHqpzhkb86gM99NTqM3JNX5l
pwHuqtbq3AuXzY4lvTHPMf2H4pT1EIeN1qYFGsoJJ7UnBH9F5ndKMoajKBDxpiH2
i7AeWujTifMoT/7VaEVnrEzQz9q3p1riAh2/U6VT+wQtoQTuAe6a0Jst1mzNuD5Z
3Q6AC6koO9V7vs2rMKPIMPtP/YX9IBqHVMV6ZTnelRMMNStqGwrNqxvNBv5pzZBz
0PlJ9JVT5FkBNISFNvgrFslEqcNDAR+4Y8oj7/zoEi43kmUQil4a9Dz/GF1vsYOD
/6YRLhGiqkPDtTg5QaImW33kFcf/ovhBCh9imTMUYgyIMXdYDDCdgCzsh9aSahS4
X6ePNcwA9sqFYrIJArGYgn4QDs95Pu5bWxDYdqOi4RtOEx50sXgYgBxX87OxW6g6
XJONBSw3s5XMsEDhZZnlFBPTGmMvKznRwr5cCEe7Ku4URIVMeyIbpyGuvC6KWZQL
bH/ZRZiPbndxW9Skqh6rhuOeJmOqAUmXeT8mye5JVE3MjEjXeqctn4asvYAhQoOJ
CrMVLyfTvxSbxjuS8pja/nmfVOMxTWw9yW39BrmpBg8J/yUyt5gPHXKNuC0KFOVe
rvcH75Hft/Tzi4PkEg4fFy5SJ4ytnoE+9jhBdPD6tciDJ9dVOqQcXVHK4Ozv6gom
3xBkbCK79TwCAwMDwnqxAMRS1MivmGiyUgFFN6ekl1pbWuLDikqixaztJojcBm+P
WZHr1l0kQXk5zWR+1QYXAlPpNz2UkC5QxOnslWhnHI/pA+pAZFY9iOQMYHQ1UwCR
bqTLUsjBf0JWbmpTNd8jnMhcZvpKqdtbiVVX0+NHNOI4O6qJg6/pZsiNvAuL+03Q
y4LmZXYCaVC2H7sXXk0GrNhM5SgjqU5qkmlNYNXhzh9/wVB3QQLp4fTIU5cSsqte
ZzV8zKH+Ne0Hk0eWA9bl4Qlm/MUk6htaVnu+YP0ZkmX2QquiHNjw2niH8zjR0OsG
AgLM1H00QyFf+cs2734T7N3Rb9zAVPlfO+GJheIWec/fOalg8pIG9MZRMBmhiRNE
d2R5tqz68o8/GIORVIIHfmQgOEwfwek5tDD32VBstWBxDTZsStrttnw8kUt8JpAY
1KNFazZ+Lr9tgGRN1v1MzCo3wrg1yrOyZ/bDbObZlGSxgb26Ee7c/K57pBDePm96
o6L1PG+r3C8Xl9BgBMaIiErOegonloF0pV4MY6J/0EavYHQAX26GDeo4yATmvlH5
/xhY21JivM5GRL3Rbq/9VdpyiUkJdLfpJWElxjJvYOz0czHW2JSxJ93xgAKppPhe
nuWO7yXnsGR7ijjVVdJrKUFqIZjAt1eBPOYAT+JifhDoXvBNOVhSTEi0YFetQZ1O
gwOQD5h7Len0HaC3fQfdTTaPDzO3lNgaryeIPsr506iO/L/yXUWvX8v+UNo5ITng
9c4RxUv3FnynKv4ow5qh5Q3WpmjVGbbO6Bi7PYSfAdOtJaW9Q9nGr1wmoWI7uOA9
VFqWsf6cBH4JJwjVlSLIaeOy9IGeJww3LN3II+qmlLNevYuU4Rf2PIhOBVGAnnHk
MeQdmV7VcrMpoxIMf9ry+5QGW45/ip/eOdIKp2yoDBCKRqIh+/APOIZzAiAYn7Ej
aq4UvhwLMJG78J8znLdeIg4lJMqEdw0dzrz+o/AudjJfQ9CT9vWNKdiZfSnHdQXp
NKffssRprCvNxy4IeM77g81jMgtcgJQdc3+MYzVLN6CCOLnNNVsAsRlW5JGZFq5N
es8UuGZlONCumK6TKvR99PaoHGtXWzAG1OKxz4NDQbGHQ9BVwoPGQNP4Kv2xfizN
jmxx+hmgnkURBsbcCFlcnecVhBRKJ3iDyCSRp9kU5ZR1bUFLnnZceEHLWwqnnRTt
FEMVK3BSGWaSxQR4OXMQPdnopd6sbdF+AARHG7KDymciXe9Arf1raDig96YP/x2F
qBnN+4whhqGCocVhwri2KZaRypxOzGy5TvG8jUvRonDKrU8u+dIN89XXNX+JlNzK
W6cuin1e2LDPCzeh6KU15CJWn5UVNtg93DfJNsBEAJHrPB30nwCMlehIHIsmt1fU
BbW3Es5B5VUu5kKbZ8qBhLkn8/RnNsr4EMaeiyfxefbqD7iFtroSxbAZWxiMxaBj
GIzetWZ0hX1aq8iPSZIlDrH2E9NKEhscIopffyKRI8KtC1XOu8KZ9jeL5Ok4Q0nL
WI0cCS/1g0CgxZ6GRBcKGKH52/uJIE/NoVr0M/d9QN1zvCuhJZ3zqixare8Cvf3H
KjhRY3yOUcWWGKLjSCIhB1CI2/JFZe9H11YKnm/MPQROTggmX+mLXKtzKRt62Cif
tH1tdnoT8A/7fauwjbYPLq8QgWV/ebbGC0+BNZ/MytroWgWfSltGKYU//nmy/ujX
uwz4FK9o5xq9qfsWPzAz3zb0iSeEjVCOy9K+XBJIFxxZHf1/jsS1Hh3se4hK3il+
qAtos+qe3Uvcrv6jdgmGec+eTCks4mDk5NziVeAcfUlPedKpDZ2FepJym8gD+iEj
W4/5OZXSGZYrGHr5NdVR7SynOopaV13Cz6IFgvLAbcNST1ZMfbkWaOHOLlZYL6US
Jb8XbNn/eu6rNp9GayiF3KlOSg5xaWtlpx0HhHTfZPc0m759fGzUG1C0REroAQ2/
EEzuIO5mK7SL4b+N2nhNNcQVQ+vatPJCOuy4hMQavAeCQ8JygQ9ARDa4skd/SD1q
58mQ3mLO7yNBq5/YVrlKKGtwj0X2u0+oGqQ58s7cEzLmOcNZiHab42WQQL0hb8bN
vTGuZ2BAJBc7CfcuEZ9PoLNkoR/H309F7cx4C54Rki4PqXFE5nSjnx80DzrwGrW0
QNxTJSOgG/qBT03R5m5f4LkKu/OyEmPCr0lk7HSX+ag3CP+QEdaE3PckcBlZs1j6
kJeORbtoPK6wgGbzfq/fEyo7aXvw8Irswn1GBGm6oaKdsG5MgdgyLBidgi/bhMdP
AxVYbSQNHduz7pi1hve4lm910Vth2OXO4j5QkVtCzx0UQqELY3CS6g1vmytGYudP
8/9IM5T1yPrrqawLzFV2fnbJfS49nofWn/rue63xG4FO/Z746V0qQbz+bHWUEqWb
kDAKxwzBGnqHU5kC33JnVXgAmruCD0zfdxsYbBFBkj2IwXfJ+u1zMfM1SoqSTBhf
0Coai9pwITq4xwEozZT6ZPAhtDD/gT3qOUa8zLFAsvRSlx2iRTrKVBujuzJLhQoj
DuwX/go20nHHYcR22FVhhxuuEZhl826wNXda1tq2RAVrBOaAJol63Fy8JC8sCI9/
Z6U7dmVp6zi2eugrBW7QQtf/UbYnUcfZHKdEgzxtkn2eL3qmdpDAaxf/SLbGvu93
WzGFudja7YqAgdbOcAguSH2gezIwT2EAGmWIKs+4rkmX8u+O3ZO4I3QIm5fGP6/1
N2X3Yi9/RTR7eYumYa51UrMOaYh0gA6GbMJdEqOhfHHKHFv1XXK0qd6BsFyaR7xr
jTYMW1Ryc4AlKFCyIrr+ch7RuB9moTmbzDKr5FC6ikbAMPOwBDEZt/kSe+SpMTni
LbDxdPQPVJMEg7pmclB6bSJxQySC1LXPjgWPMjS3c4KEwMbSnqgRgqDLDwd+fTiO
8hTTjtU/7z3YhMH9M375kqFue3GqYWVdEfrKLZIY/Qz/GDNmsEicrYk/HqrOLvwC
u8GSXESRytrzkA5J4JFo4EOdbS+0E7MxFZxOaVjiZH1vEDBhIWRI0UKTRMCFUq5s
H82tGNrbytSu8nzZUhtLsEtPK+YKcid4BSMXGaaqqO2r34642vzO8kQQYlWtwCO/
bC+YPxN9EArDlDDFlRJq24KmZGZtCrT0eNqkfACgMN3E97CygxcslHuTsVvxEuYr
EPnHCIdbQGUx7kD3WUQ2fELTAlYG7umU7BXIYuIXjvZJD/FK3PmbtZbkOsEy9jw5
vTSd28kiY3AsD15rgjDALmQGphwEgBYM0NoK81Yi0BV8cICU+5g+/dVSSfK5KH6U
TfqB9WtPayEKhTWejz+9gn8vukqgLjPHZordu9y3C7eBpLFwFpl10UEhB3C5zGsW
BhMG+ddtsqZxVcYeEA8RetV6AFTtD5sdcYKW3gpLikYlKky8awx9fZf7phDLi3H8
lja8Wma8ioq85/Nmjd9a0/RrkE4ZLizM2GbBVtuGPd7EdsvLc7MEe50/rpUaaFzP
8W4s6Tbz4pxGFd4+0QuAmancNGRd3QXMRE4zQRRKZDUwe1gg7iAKgS4039xWq9GL
fBgVi32LMniTdjqkcF3hiuweSxYKzLDlU24TId3xbP3ilJQtEYWf4jnjbwY9YFqz
KImkzN6eHcDuA1m6qxvwPfNSO2SVGz7vzO1NRqjeJdBtX/y9wcL6sqNeRtZwow0u
jxQ5Hxvj6IYuCnW6yynzwxqogQT4VeCcTwGjJ4EQJq55uAzeZk/piSUrh1ONbSUe
ph4wYo/lT2o6MqKCk62sfQn1Hh4FdgVkHKS81ZGpMZ+NIRvs2+/kPjQVSuMCOocG
yfNh9gVe9AkmU3DImzMwmA0IC3swZE2HZEPU4188cm8OHYn0Y5X2t0V91pgUVv/p
eGVQXt62bFuPcjQkqfKndMU/sv0mLjCUHPApNZ496KRqnnO/6cpklxRdCg7/ZXfu
a+grnck9L575vWlqLXrUuQL/VS6Bi9GeMT0tdBowUQm/fwNi4VcjtPpZzPAJGYsP
gxBu8t+K0K7tN4ZH/UIHEP1txRGljkvqWxzt1UuEbVSCqsw2Nj7ZQlSP5DHrHpQD
+jWDkx+HC+HnKZIZBmhwdG+qs7DtYlX+9ikuuJlPU34oWoTV7zsUMSZNxQi9TCb0
gcqRoOpDLkefJ+8kP2CYpnrGI7g8d0xRFLRNShJShYE7MUnHGFaKG+Mwx+rl4o4E
1mAEtsXrJOi8vrW00zYLYd2wjxowBbCw3iu7OSfw7Fqx8DNobOOeSouF4HGfrhEV
dFVWSj/VKC30Pdk+5xlc6W9nISdPEG3wzs+mmHlRxTztKWTFPx7z9A+pXsKVVg4P
+cP81er+48wkX0vOdspPsY89jlz36lvVa0OV0GdGK/DsuLjqG3RKg4vwrj4tdMm9
pKBpK4BYD9RaPJNDljk9FsVI5yKoyeCo9Et+1IfLt42dHEVmOWdrCexQ6xCySwwI
jAr2cirr8DFikFABMUNCCxDFH5cRnINv/F3y92LO/asyEAKOldmX0DJlvJXZbgdM
cQfJMWgUF2ietWU21PnKsLFRatYRBdgOjuRzOWL+2g3+SSHS8vkL+86Wxi/bfdAV
rsGQmrV7+hziOQXnFBa938o/YTBmr/Jme5wlZ4qpfXNkQI7cUAcQXpoR/3Z9p/8n
eZm4V6UURW1xXQmVnmuu3/1vzU8UxLfKhGrr8Tsnz+5jMnvLm1uVX0pUV0TmHxUB
w8rtuIWW1ikt0d9Sqe5Knkwe6NkaT4kTej6wYgd+JGs/RuvOYS+60b7qR605oCtQ
TKXTND1m3+6dQcP57rDNC5KCIS0U6vJwHxXjTikoF2DK/lCyxt6wAxrMy4VUCMKZ
sko3lANQOn37/ELOe2MEX67DDn69eh+0V6DEakBU0Y9BP+kmbdyFlDelNz753cjj
vSuJk8FduZqkikQ4XX4pDKIu8bXGRt203fX7wJY4ObONUV4uUZuAvf4UTpjWJfJN
hoidjaxvi1dGAjm0uds9ILe7Z7fSwstmfmNB/tMZ7vhrNU6xhLwsv0y8fk0sf0tv
uVQQJQwKNoAaWp5Iymf72dkQDAGmf9ulX91fP3/5r6wyi+STaDfrj1oou6EpJ6f0
X8AV5M09w39xpHD2N423TrINeRZC8fDie3ZNHsBziLXjKi9XPskkP3Hn3h+NLclN
YI9BoLkso0yu5O4x3Q1TLTEOnadrX02xheHZvpWk2QjvzEoabbRPhxdZDBMVqNUr
WcQHyzC/v+ACBSd3FgAOgobzboF87mjSBIBeMonbisrBZ8Tmh29eB7IKXqt8LHbE
Cj5px/prYisJGKaNIBQ8VfqrbhuW8wkzst/ucGeCgvSYnZ+TCAEhcScoR22NqWlN
Z5zJM+UwC9LrETy2BRUlvJlmWaDKyu5+F+cvPmDSuYtStW768u40f8kEh1GKwus8
5C4jnj1ayU0G1JSa/rNb/vF+dyc6hC49o9n7txUKvcXvBAhvUJ6rH6vNTK/qL7Dn
fko1W12OvDuqq561bGpGQqYcJhWqQ2r3rF/H3oMoxVSeGJf9FAOKqBXb74y6uhH/
tuTbjktd749hriS0nyqn89rc0/ekZVo24bZn/GBW1l3GXD/C5GeizszpQwXWAf9n
28fUbmR51nBy/zLYhHc/M3vGIgmNRIPNpwL76raX9d7rqAVSyUiPH2orqr1XbHT9
KOKqliXGzancllHbmarsWNaw5Pbjjl3O5xJMAUbMAuXzHyylfodCGdqDwkQE49bZ
212a26MG9tGSoPlBAQViqOxz+2ncLsOeJN9YzAQYH1q5wi1qcwJYfMXuKrr+QL71
/LzirAllTRwo+xgO53UbFRWDO76YQvN6N93UmVUymmV5yKHhB8dhgCXpR7vMZR20
50KD2yVhkDdAVFtku7VMLzKSgxnXAeouTKYqTKJzggmknTrh8zRf6oc+N/+1vRDN
ZBJoQZliD1lezNvYLeeel36i8cbkHYsMZq/xbKxiexkWjbnXtKCHKlrJoUyEnw/z
atxFRNpyF+TgMP81bfo0LaleXSYaeCMVI6K+ofRKQEhv57XdWvZCZynEpqNIF/95
hKYWwf4fsChoJxOmMWN7cRmsU8hLw3ySb54S3/mrALYPFxbatRRvT171IxK/AURb
9bIh/HdfiD02JgF7OUyxtF38JTOI76Av8h5QGc8t/kQFfjr6eDtLuTEg3pjd3fKS
GTHAPPv2EXozVCmM0LfyQ9tZq/9eUt621C7sYtyeiaU1WbyJA6YCzkEwasicmWQI
SYNBY8fKpJcrpLttxALqRNAmOgSjwjTh5lREkin24Q7m1ioulTcEZerG1W3ZZ0bw
OxviDmnLKtWTUsRTmcK4UH1hgdtQAgIcxscnp1MZvZ1l6tmkyH0DXJ7GT6CgL6H2
kjlmWlEj/lxTLnHJ3AHKzRfdW6pUh4EMN5uRJO4FV7spkLGhw/eOm/VzjkkAZCOU
CcLqDidiOV4FbFs6d42nQyklo5ClXcCdj/GgSCUp6LupjMnGrov6AWRY3v2t4jeC
1h1rJ/LmfxqE/FaFYW8jAf+JiQ5xl5gsChIPtACHOS/EnjpY/lbLQjIF20HUz/kL
yDiqmEi+kdgDFaQmnytsW3KDfpHVMXqw0k7xUjax76G0o3txu2iCZtvd5t82pHX0
NwgYC+UINs7vF/f6GdnQH9OfenbIbOydfONx4OrjszJiytaNqUACtxmSq5XcXUn7
1OA409TvhPiHOKPjifrB27n6ta+65likzluEGp4xp6iuNzro5smWzKJ40ezueYVR
lsATXvvhcirYoNkT+hqDdJsRiFoTuDuR0kdP3tk+RQjA1DwpXz2FH+D9U/vmfvBI
v8MM9srWRd0LGgpvHfWmNG82f0ffbod+x7p8lDyb/YAqX0Nc/SvDp8s/6lNoZ8rX
0IyiT98J816Rc1KPWV6oxAisSghq16Ofs44g0qE5tE0p7b6TvJOX/M7zEbwUdgMb
4inX24cxUgnpoW4pkw2i59hIX/KrYFTEKXh3bJ67UcPyPsqjL9RBYWaPVfhYqD0m
VVozrYxaONCq/pVBW2SRmhDxlBZgoKS8MRFp2Eb7EZhkXqf8s2a0nBSmNwNXOp8f
56T2JLZjHL/62PBPyf/vA6vgtAhjctOG8iUAj3XJizwJnYRAiBatD9bEWuVgEdZp
YGjle/J4al5tPMPjPt2AzbtGSOEzt2X65TH2GTriaPJxBWfs3QCVflMlAwlQdhOZ
MwZW7ZsFiaxcaPxYHsM2LLtIB7nZPr03d3m0qmCXgCQC2wstkAiOko335woivbGt
FdAfCPeV7rl6IbNIy+NLBIWbxYURqoaQ4HvJVlgkcfTLMk14srNhQ+xUHBux+JUl
d8ZM0Zo2kTR/93ZJsY+lawxus2ufP56XXW6OsIFVbSGXKyaXquY92rbMy0FGlFhG
Ij81vLu7SfgvtvSg7mts3Bp7jyvd8cJa+8axXlh6XDJPjTcQl/RjYKOeHzT2Nhvh
eYqvX4RZ/jJXhI97ce0bqyiYrRJJ5RV79M99IBrEsBf976vq3qI7eRJNo1BU1M9f
MDlCs48eU5GzVGAjjCSopDcjHjsgcsr/HBv6lbUpbQ55qoDJHoVE93V9PAuCXjBU
R51swU2DxNYQ7gqhwPMOoE4jaJVeiaTGT1b3Q2ExLENCq4Kn1251GGtlauRP5YLI
ESq4BynXwBm4j0udflVDDLGyj2o8EQxGF94k74RLXByYa0Xzpwkm4u65tDR2YL/y
uhZonMVzWIJlsxU0jC8AgqLRyQ2kviACPYyoV2Q1BEqCeGF2lhi6b84H9Zotw5WK
vOOuEW0+3Gun4UXht0C8ljMtK8UZVeECxF1m9BVZJRQPU/u6Sf28BdZCI9T1A29a
q5WXHSzJk7xawIJylwQAAu0ctEjMT+emXhC0xLxQJcDxhb0D5U90+MloUN6QjMEq
MymR51+/4ROXxPboYS/WT1oVCuANeGLWY5QV2lSSIe+7W8HZtnKTg9ZX8ZDS4u5n
84eCb0HOdgpilfXDDns1lIVJVmwaseJ98uBgAj0+NZrvN52hunYs8H24LlQ2J75E
FeWDu+XS1KyVuJ3KP6n7O5oXDV+U0pj21LAKGS60hPp2dBCPiNQkv5UECFLjpmWQ
p1i0Yaj3FeanUWQBqJ/GIOPb6fyUVVwOsjqEaawTDt4dItXVn5ZmDcBBjuYS/UMZ
HvjcCnWKwiz3z2PQ3i6EB36lAzrXBwy4NndKZ3aReQuL/1cuxUCn2D5YPjQWvwH1
lqs6JpB74jlhEhg+UWKCc7LhuMMeWIIW7HdwjAjeq+A+53hgYpbbtgFf6Y0blEVg
/qKmziLeaURu+/seJOLTRGx0/HiCWqExJPtDb6Wo5JgYD2hfrImWlkyuu4LeZv/n
PuayN4sgGYeFPqJFQQm8Ubd2ITQcYm0qeTuU4q5Tj36i7Cr9+0FSzp7jYMQdVIb5
gzs3pSUq57o75/O5LXUYPQUr/x6/MISUKgvSVnMvjg+qN+GIjeBkpKTWeanKL15H
Ez1kmZq9Yr8gvmZB/BdoLGB3YJvOfQJCMVH/PugHxwMxlZ/O8pRAStYUWBY6Kc3O
F+C3vN+p/jhNICSaYhwOWNQbFOtcnaTIp45F5tdEwMs5UKvwibMVUoYTkzz1jGqt
zkZCjjEn9e45qtvEVIlrLqPiM8LzXGSbww180iWWpnVl1ItSe4gus36Qd06QqMXw
CSTKpVAAlf7jMxOFgVFF+FXmsP0k70KeKvajdILIyoerNPSrxUt9+yfenpYhRfo1
RYVDbKnAwxv3kHkrLSkffVk2NdjIfRyREVkMoUKOWvbJDd9dHiNmqcb4NAGLrNSd
ti1uEmYUylz/vNGBG5dmcEflN1LJgoi87nF8sy58//L7Tps1GS2IUn56wCuc3Q5R
99AM22Oh03Y/fvpsRZIVsRneHCpRMay2Sz8I2v0NS38xAxCZDHlJgpJp2Uln3DKf
fhwfaaYd5ddkdtybUrDKywXHoxqW1MZb7KhYXnDh4feeYYVXamH3gtAsPluAxsIv
Z8sPbG581zW6G5HlZYcvyhvJxEuFhqjY18OSdlC3/RzR6hH1FeT8O3hP43EsWLkS
0EZHragEnoj91QCbLFwYWGQ6Q4bFneWmlwkrak/ChpDutK+K0M+AVJywL222Rh3h
uNolW4TQMXU/EuncXPczl0CS9+N7GjvCSbzuecJDoVKLTV3YVIek+impfgkSUFbK
Qk46zM0dKhNhBWdxU0v/cGkhMpxWRoHZwn8zbCEYfLkZpvrXO74/wlzBnWp0BlmP
Bo0SRrajLdFSAxGjAMq4BnhT9yCXTiJ1rEnnVd98zWaMp/8RLRdWtr6vezA651CV
RxVh6kIqNB5YuhmO+vOCYhcTNnRqGyjqGoQzpkRDya/F7iDw1iaVu79ztb9364Qj
sFVi0Wn3+Lwpv69Np4y2lmC4RpVjhhYTaeot23gEbi1nAkI47bNbLFhYlpjczyaC
Dij/Pe8m+N/umiqL9d8OtAB162tNU3bBM9HD/dU846DL1ewCf0BjFHoaVBSTbGbC
NX161dJuczubgoF/+RKs0PcjX6VJEpGihJDPVaPmyTISheIjJ297H2/T2Ye+SwkW
uYRibH9/64rD4A6XSKHy0AlCaW7NMwOrPLEJYMXx+LRY9yAGhTdTV3IpV0bRKplb
2bXlMctZuYxDuz7dOs2zMmDxYIEHjIFrGjDgFAanWoGf/dPfGGHbW7+ycUYQrrTs
pS6reC6+GSbpUNXu91fO3tq/RG6w9cftDQVpOoUZeLMcyR7r/uLAb7xc4RYUZ0js
R6UyfgRBk1bAU8Cz0Iz1ekTie0UbJ9AklxD3Pfyc6tJMr1UNAN7lXgQpGwbtzYsH
TYHLpXGFEvsQHPzU3TMV78S9PINy8I6vaEacRgmqHaEKJKjAKPTJrcZiAHVRVe5F
3wsEP3XlSK2YCtm2ZDta79qmrYxrnbi/2jH07cEJCTUaY70r00X21UIS0qcUUg75
5Nqj5x/EEApxjZJR6TldHxbkHj19fN64YCT0dDjGbc1+Wg4f7Q6umCkaql4FG/FZ
Z+mskHYZS92UqQWJc2XOu4sC6dYSyp0gH8RnJPVkWj0CaTwfah1MxpH5omucmj6d
MYkVW88RNS2kVAj/19nTXLwEJ/kZsZuieLOTKC3n7pTD9Ol457KM0kSyFaAHfCwx
3yYKohWlswH0JAYHtrxjK5cZvi840bHPbbM7V9CJ/usScKAPn36qQx+JjdMfyq8O
aBw9s201jJybPlgowi8J09dVu/LK4zQchHYCCL+54rJ4TxHkc7Oa3XByhxJ7D2rw
CBsBXokTqwfEGGaLvscsCqEOQviGC+uNN+sFKYftubVATNik2Nvq2ChmwKpgtYjP
QTiSCjFdgmOAzllk2uJ6uNpr9Gt7IaqA9K8USvANfgFSOSulkFOutrMkpivco2rw
2O2yId+M1lZ4KzB1e+4e84kjDfQhYQlNWuxkcLnCX0Qh4irFiQ0rdbhYiP6/Qxxo
Ixnp0C8SXiEhU5VWlKYVLOipzwWdg9Kqg+rZMrGAPlDD7fTiISrO/IQ/IRNatrWF
Qg9nGo4rh06UKk1amRZKePwz/Y2GSLfgIddbrhSpB2ktOa9ngOjrsJd9X+HkvOq5
4OjmDAZQ7trYO8R012wCYZeI4J6yqWwUYL8HC3S2s2SnGJorqlvw+77yyoSl0pM0
+TFtVRws5GjFd686OqvAH9TDQb1koSFn+hLH8dQIw3PXfxF5jByDTow9/WZSOjot
o10ljgaJga4x0FQ3OOh/0gmRnV2gBXu0EqOMP6eSeQ+Y+rWZxgaGByX8ipAn+KaK
eH/KmsXUBTgQ9xmpZmulRyZ0Hp4KZhpdndQi0/YN1BjvxKmkp4tt1MAImzNJUL04
aeQ+jKLgug6aOxVeRy9XnD/7ZM6GFfhUzwrmWLzhRi3euAqrf9FY08j1iiT+lz18
btx7JHZhPvfnv0JQxZM26YuY2hdxlHPRvSFElqO1xYuzcNTXJ+wp74aHg5KCGoQ2
7nVmJLUWzNrduPMPhjmcpr1AYlW8o41z1rX5KwNkuVwMfulk6dMhCEXCjSf0GUGK
bBnED6Qhlyo2/fSxb6pRh2c6IvhK7UWhLh9g5uRwt6MwgS9J8vIeUOCMf4LC0x0F
q3HZU4kuznx1ESJu0Bv/A82T84gU08cSYr7mvEL41wae+M4gND257VHXufOk6AXP
rGGys2OymMeGAylPCUSYfSLqSXGVKje64ovS0rkZStU+Y3VkmqF28pNwCMf8M7O1
bMXrhy88vuPDHkQWbNmLkYX/5XWXMTmOH+wHqY0c3ZKeYgGF4kGY27Pmhs5HJxsn
N5F1FEyRmDBi1KC4tCqfXf5Pl3y8/nIMTVRymqudtvMiCr0S0LIamF8fTYPS14dJ
La5BjLtChOvilfoHgaS8SVxRvnkqV9L8zHtogqqbJR4yPXnstf6wW/KYtwKeED6b
pVofDPfBhwlJFJHC+C3DZvzJ9/+yO6SfNJalqCwh2oX4I+5WU+D1Hsb16xNCSklF
ltmP2DR6w7pZ54TEcBRTgaN6ZZJ74c+Xla4gVipGN3ujQpLnxxwGfH/VHY7S6kmC
UX6GPhibOZpfEKvoatjbA7jMmgfSM+8ih0B/T1p9cuqG2NkE2DxhXgDrqGfblrpV
l8ORQriYyYj9kfpZGziCLh6MvKo825fhRZQacCc/IyvFxI4Pkwei4QH+rUHMnZRK
gj4sitD+ODBox3pKsyW9z4EnlWdCSB/Aj3Qoijqp9/duPeNrfjQG7jSNAqNITwOK
LyxU8sN0O11mLixL6lWWjEMMU+76TNzWDVu9FxLJkYL2P3EYPceX1rFcUwIeGPK+
j8VAMeEsgCqdXmMTT/3D5zwq89L2NosXwxGoqepTm4URKbvpknSEgx41y3PcHmwT
3wFSyT1sP3NH8WAuWpGkkj5bUkZqGtBM1t4fg1uoX/Q5EOc9TXA4DvR2lLYZBzuE
lsuC7M+MMMMCTQNQga7DvUjyzKtbeAMK/6lOg9vKQjVNmA5seeUf5Ybk/Eigztw5
/9RkUsKfZvVJn11fr1gFig/4rbUJ1jqMoqx8Pv1Fw8Tlsw2vi6Y3+84k1MXfHjSR
SsUpNb+1y4PJEC721ttz6qXF4ByTrOsmOYESTcau+dr2M5zSH7CdqJ2Nna/4CCGy
QWjGeKCnpY1RQs5kILFcK+nK1mSuuoXUqwUgb+9oIHaLDdmZpzul2GmtrNANHjvw
0ndYPnORs7k8VM6PSWst9bt5atF4iGAb5UYx52OvArNrFdx9M3s/v5dt6ZgaQN8D
llUoNHB2DywGomR0/oGdf3c9FHX9B9spwlM5nHQloms3pXGAekLWRDqNVrFfwohZ
BtRZDbAueB2Sg7TN5/+Gb2jtrUNQifsUDVaebJ7ZlnqZOIjlUffKLjVHE4NH7lg4
MqTC98Roohr+xvwIDoKW0G7mOfU5MYOnn0ERFgXuXWzxjujD3YGj/Sbktg9S5aU2
ZXl8VLUpfkmY59LrrjN/SS24MOciozITXN6VqsE77QdXALcv6hH30GJkyZMy/TOh
cCg7Qi+wdKA7rPZDHzdc4eMt+hcpEKahNHQz1JsDH6l08tQg4HQrNieJbH5oE6bm
4hGvmnuEUzpMbPm0M3MWl0O3nvVa7RlbAe2y7fpTDc4MDsvOJ2sLFavJSAdf9Tsz
/O2JhAJBhIG4X9YDz9HmUSWLkMPUyKNUdQeBCrEINyWQ28tw8gbAEj8AUv5TFUK6
UgyRZ6PmOuanmRlVdg/G4nX+Y0D9v+RIJnScLPoiVhtD/5Sgq9Fkx5X05OCLR+rv
zyDaJYG2tmpc6+lKyiAgUnM20yMJSLydDOPqFByu/t72kW1QRB0sS01t/fa32/Fx
EligfX2Ktz1UoLZNRuPiMXf0IIP75MHECYQUTD0UlVQwBp8n8SZsdGYliaDTHPU5
41jUV+yDN4CbyIkt6fhV5ZOn8CiFgiBn3WyPdoJaAJHl+Vjlmg0sbNI7PJIG3IWy
EUisHVe8VfN/B3szmZ/xSiBUheK+uqVQKt+m2dDSiJsrJAZ07PZ/YfDSrpu3PNyi
HL6iGp6D9XVn7DkicdmH30xiADfN/k6MGP2h8vVn8nZcr8JyVTm4goL2Jxo31wot
0P9x6al+RpIgfPvgQ0Jq9Bf50825fELNxfU2SivJEL6DTxjLXT2oVRYcloq6Uwq0
McElzvIlyu7CjY3Uw0EyYBbG3WxXt2hTJKq2gYpaWPLjj+fphsV/Y/0Zkuh3bSnE
Mgtz05pb26TwF5L+8GyZDIPr6uGrhs+Pn75bl8Sr2b82j3vYsZ4KqvDcAXsu7QLM
qpro3oLdPdik651gvJ5TszMnGvviuVL/WueeWm0K+8kJKcSZ7R0dAsEgH+uvjd9I
K6/Bfpi7XFt2qjYEkXazkPlVV8JO1R4V5WJ5TG9gdhD/4Oy7u3S9qSOzb6dkNKc7
Co7q1XFGorYY4DLRPcKH0DR6krmpGk3pJ+qXdKUl8lH15DbyHT8epdJXK2LvW99r
rc2tP2ii9CAkx6ORp8K5dmDlnjNzolTu/8aFM+83YwNrzU6Fd+P0I1U/t55iLaJ2
GhYXVMtJL189G5D+6nR6LwXPlPON6S595N7QucMedIbqxZOfyPzST/HZRN18UH32
Spale3+P6c83rJeF72FSKFPRhQGQlCPwImkjE2CgQOkwCFf+Hbtj5Ra/p1TOVwvW
fRO/+hvO//gR5Bhu4Q3vzTZr0sn1GnkgIbmkbQ6lX8/6ZTNmPs14W05Xd+MLna+V
6lGPlKPlCcyjyVXmCsAeOuOo32oPEfGKA2hYa4TTadKlpOiokd/6KNSvXoPOev7L
6WC9jfFly/iX/x9gcoNbpRAeNfozueR34e8gBK55Fox0QSgSX59+18kV/rS/VT3t
uHe2J/KUQjR90jPg8dT5oluMkT6cXMtgo3UO2n6G7+lhTnMARVFl1BTwDtAUCexG
9h5ft731NF8y6/jIt1bHCZUUxDY36dJXe2YAh5gAJdyY7yssEGLMOyks+7aQotYK
TdOZb2+exKuGZX0aH0tETC/mXSv1u49g8Nf9keo38PU7EYZeFaKlFFtr6a28Xk5E
hv3pyEx43aANuQ90TszOI2bQeFBZSlSPsedwRC8GWNxXqhz9+2hVAw8s1Y7PE+Y5
A74TdoqCvljyE4lbagBA75r233tkRaDqymg9OrauK5IkftMNKZnyj+d92DIzkKPC
wT1EhTbGJSuN0asIE+RZ39uSagAPWz3HFkaNBrNUNFd2PMo1jW90zdngwShG8IVb
Qt5KZQGsZ9MXD94JBiW2B0tZQz+n+E0dhxnh/Y8P+1SuhXKsjqiCGyPlZ6ePUWZa
BixbI1sAB6PVXZv7za1BMNO2NIJGUVHPgpNe8Nw7Eu8qqOvKC0NJKIQVZizvYg2p
uEJ5bYq8d50rKCqOXd0kmcXrfxFU73NKlGHXxqRBg1ixVY3NOZ4Z1u3XFWaU+mzb
lrnkyXvtq7DcYk4S2vTevMqQBsQmxbgwDy2fwbLbrTUOFz3hN62O14uP8z7t2usV
AArrvDC17OyfFs6KW6ChTL5oXJsOGrpi4bluNDaaQKmmT9d08u5udmB4QjQ3lgph
tSxSer0mRIFermi5iqUlmQ+GcZWdAl1w5qot/ZX0ZfPy7PAUY8Qw+EtsDfXqiI/F
fYLReKfVoMUlBagiaFjrM6acaI2mgFWLL8GFcM+lYp/qea53hsb1EfZBabVuSQHu
DEcIj1RvQqfaizxwCkW4N0SExIT61tY6mG8DBP5QWRhXv/BHOLP6THpjCfCIRPiQ
JXdiBvmz+t3R8KeboQBeJWzw73cyIIlVqpaoC5ui2eEc29CtHitO8xdi4lL2TCd8
D8lcGZJjkdxbiyjd/pBQqq9BgrOYPEw9IvG7l8+ZdhzxCv/JRIhnWbSgLlK61E+u
lBc5puJB6EOnlZDIOPGUJdz5FxSCRLWig47kSRim6BcUK/Kgs22yn2RNNvQY/rpt
jj8/nXkNNqjSAYnZ/jjUXrqRlvup/jUln7JvoQ8gMTVAd7PnUr3pwZycb7w2qF6q
lsw160r1moB7UmHRZCFkO2l8tHSeQGY0yk9eZmtx6DZuXo9R8rbPZ1or/uVv7Etw
AnuEw9kBYrdLmyU45BE5JCmg0k7G03Nh3P4KZO6Ay7aMAQWfOIWsu0GCBjRClbtL
dMWO2NpkLrFUgRie3wU2bFzRBk6qBuxJJ8pE0lnqH5FDh70Xsqg7DtiI+p2SaDeJ
tRtfB+TPmCMMH4BUTgt8+lOONbdlqZfmDuuW9tqgj0hG3dLExMX0qWI896iAAxRp
s710o8Pa/s3r6PGpTr0vmp5c5tRPlgiLOKgcA2cZopc/BU0V9PchraE48hP1yj9H
hN/XjqQFNi5N7KhZUV2w+kuORMh7BTronLrNlEXU9IDK+Ul04e3Zqy1h+E6b43fC
9UgRMq1KwpkzevUTOdIg4Z7MblrSei5AUMvuCkHltVcKG3ym+NDyUgSCuXIDGMv7
+6XHMMFFkKMYrLLRlNCit7161NGIyfoslMSuF1ooyAVpwWpLOsMPmH8qxl9FZigq
+T00qxrm+CnNLGduCZ7ZWR48rTj/lK6RzE+l7IlLb7yqqS55F4ZcXc4wGQ/Z6Xw5
13pvTSBKXpgif6iTtHEp6kOIBG5dnl0Q9qcN7IioFvMmbH9I333ldsOPn/t6i1rb
u9GF6FEYhOWzzKRkqaqmmlkD2HAn1mR4/jFCMsbAp64YuG7BTNG4Kn09+5qtuspa
umrHowhYgiZu20StqCWhO3i+hNoNuv+w0GlwJ6qJpKidPQrAAY7HdDHJw1KuyY79
zUmSSjzeK4/ybHDC608oEWKx6YclGD4UlUkSig01K+mSovB5SzwNsDtRCYcYBfuN
mrwjPMEfbyfEiPhoPBKQ24Vjml+xp5CDYzHHT9EVLs7aYfm03L2J20VjRpp9POj/
NyE2OpwerwtZXe4Pd58+KYJML7s0X3DwiZVMeAW3dkOHkEapWugRFuGT/p+BXX+H
KmPy25GobpI/BsJ++0Nq+XDNwQFHIxMa5iOYSj/HtM8Lo3Krs9M9YkW1/h2KMqwO
rzrXWPC8pryvHuT0LiTsqcqisr6zZuVvpo+bH43i8O4nd8SNimG4UEVtJ0bPQoZJ
SZMEmMtY5L5yPeT3UcI9RXyvTQsaJBmI0u1ox017Ra/Omml1aZzCCERd6CniwdgU
64AnEN/uRbkpU8M0WeUS3R2YeLeUIyH/eQh2nOUa4OjWpfl2K5us/R+UuQJcPe8J
CApa9QYa/7dyfS2SF0b/gZAtpVc5kOWWh+7MXC3A5GlpaQitsNk1JzPmHhDlCQuI
O9j6x7LHNAofM9TLyILBnYFw1TN3vEkCfIWkLT5ObonTYdWpveSRjhZAWeObb3G5
lP8ozt9qfl3k7qlTUFsWs8NaMEc6nUkR/ILcaDdmMyDRw5HHhSTsA/HNF61oZq3x
sDa8Knjq7xoWj1rS5d1BG0k0y18Ah7YU+WZHRuCDboGcFHz6IbckxypvOFa7YhjS
YYyYYveymtmVJFoi0c/FVfws8508jny6ti2k+Ev82wJn/iO6SMUBxLxjdzXZdoEL
JbiCLyHigaCe21jJgTgNrkWIFrikMQY8pdCzIgFtRbR3tC+jDoLNRAe9L5cIQsFL
3Ymff0ztl6ZCNwkhtBBxoJlcn8JqvE4H2kMkXzjsWoNQ6cRbX1do/O0EHm02MQek
gbywboIVJQMhUYOu0g6xrLNzzANMOhSONS4lmD/twkBmZOW5wcfQpRHkCI9YzuWb
5CqC2tFKSsJ2xzNwRbmT+J1ZqWrC110pI7ovAJFGcb2GWSzoX+OY355r5zv7syrt
bd1t7bSP/ZPXtxBSUMHl9UsMpSG9XHusJVg1ljfK+oPQzz2gE6/I9kz32fJ7qsRz
JC2G4vAri6Br//l+KznFvDkZmf8OnrfjifA3ob82SlLJVRylbLFPlPoeOmDUCwzN
JRf1EwZZ8eRpVp0692fUBeXCA8p6q5JQEz/8LcN7PYG/Azhc43EPAJ+2Kyl4WmWS
mBlYHYBSyzkwHPnUnlOgeYq9mPIY0yZX5gKfjYSidlG5toG9Y2KXGRyGALA82h4j
EyGqOYREzZ1ej2F3BtGAwvzcZ/KsDn9btCCSTcHH0l7zZUBFjKEMKXVK6ivCwCCU
CR4YL9RLP+B3yNdYI8C6g5BMRJWrI3EEQc+aNw6G9r5M/8SolZePjNzkYWPS/fq8
yi+1OsjFLA9eVc/seyqI1FHQfRMo1vMwvE/+ebSKxp8GT77KUJJnJgf32wLHvKyx
WnME+PC1tAgzVo/MFlJ8/0z3N4aOGWinYW5JkHyq2tmdYupFnQfF06KjMwpow4El
vVxl+ZJtQsx3kriO90hYX+kweVDvRVRNDyZ9wN6db63cwkXAwm0VVr1lMyQVOxYs
kTs/jcHONBYg1rq0nfdBHQd4PZFvACeUK5RoGlgrbxbW7TPRyqDRku0YezoBVKLK
/qic+VlaoNt27bQfKSWJ1Qp74SxnbwifdhaZNWuMfBG5VUJuM2j7YDWvHcMhkMn9
kxSwXdYQL1QsKkpGUOmPGdxDx43iCiNjgmn5heGM4qMCb3b5C2H325ZO1kb38+4y
00d+oQZFCb27IMGSgTaZ5BjFd+Zv1RNGtNe+bRz7lkHsOf5I1vHVEUXMC7M1xlmi
UB6sRq/MXSDf6Pul/PhFM4lpWThvuxWRt9RhKEUWnrVvqTS0psXHPJgaHyzAZBMq
IzE/nPa2RV5zLSlh5FeAo/OxmHr3pqL8pQGo3fbuFKdH+HH6LoIzY2tOzRnWX5Bo
4CKIeH7ocHm5TtThtL/JPmMtI56+mqaew6T+M0obHv9Sfr5DS+u+Ge6mNndxfdnX
rTOlYN1p6s1XwvxLF/CNK1chVBv8UxvYIAmrSgvivLFdcxf71YZ+752eQXNBuNQv
FKZbvEl5Zg7pBGJP9GPC4NoU4Na7uUMBTXphuOnLHOMsZUN3xdNqQnLSKxjPFnoi
5FfrZ00Vq6GvZR6UBqzQomuTspDip7MEqQMUycuPFEf3IdOwOuBsMmp+cxAx8F28
SkEmEf+5RjU3aKtwtMXukxuGSMCRoSnQ/w7cRGQpWEqiXDoIc6iHjaMZ0hllDoHU
/hhT2rQ8K0zhYC/jXxxpZixwCX0BToj0m9Kh5fGHLxH/9YtK0WJqR57xtfy3j8Iu
zvLNANDEJg/4+5uzWeLz+zZ7sU9bsUW3SJ/zl+qKzs9WCMm4MM0N8gX9tKJnW4ux
6y3TTJA/N30GUYBTWyjR5Aoh0e3mORLaj9UwpYrClvCv44ye/T2/NKqhu8H2fPLT
2rHuNEcsroWgf2wSczPVRBdM9mCKu6M7uvilHyAV5gVB5jtWTaHn6WyKF8UMlRkM
r4uV8VrviqXjvQgxJ8ZByDQjW41NchY0zMTj0H5P/6KgG0/I7UCcLv2RM4/8JhQ5
fOI5JKIbD9wjMnuriWT1wsgfClUSeqifSbiIs55IjrDithV9JeAjNkD8HW4bP++V
r6ADzFqfOu2aA3akC15DE2SvpdazfRJJYuJB9I8SLnlsAQA/y7Ktp0w33ZnRXl6s
GldQcaW40KBRI3ZdTu6TedhxUTmicU1bi5bxeD5mRbMDy/cMwpMPXtkg0XV9xcrP
0MJUP993zh4yXZGBKZ2+B6AfMx6IR437xZpcQ4WBW/0dGogWdwsFNSX3zIrOqzi1
vuFSVw110omdh3g2Oc1Eq6kI8F09tiBWJmeFUiZNpGAHbfkpB8npEJIzxMWZid0F
qIILTJ4/IpVSjb6w3/4uQifyK02rWS9+gs5BLvMnI2BkNi1LQnNd8UcDqIAJWFG+
jwJg/hCHz8lcryg2P/eeVbsytTVX7h0N8XWHihYTtMHEomqeFeO9AcDKG/n7Ay6g
QKLGPwlq5EDmk3gc2Be6QFAJIK64/POaBkmHgM2r5dnaZCD7No6+5vVekCXaW0BD
zByY5Hzd3ZKmeqwaBjlA4Plh+BH/rr4+a6D56WRu+Kr/m57W6TIriF6XPbXc3bAi
8TonZlo/Bp1abZmZ/bgq3zaOM365S5j6mIBEIzojaJm2e65o9C48TtgrJJcHxgMD
PzDrwmpWdPUXGmXslR6nh9Pzdge1gxzI5Pfes50nfJUZeI8FFJDiqtjb+TcKwRp3
QKtrHSDH3nXwWzyBt0qx+tLRXxNs0aVSIyNslb/Z+coXRhxYyChVajNusqN1Foef
m38mMDOKJfy5Q5mDbTIsM/TIRUWxxdHoKnH09RA3YUgWTpf6tiuWx2Cz/2FzyLnG
Rrks723tI9EKNhIHoqT69A4rRWT8MP6dI0c+xedtcYBDgvV2EuqyrcGfGEA725gm
0IP5bIWfUB/y4xkOo3Z3EmxMWxvkeiw7MTY+SfNXJRRTKHHfawlhO9tTuhG017Hn
hbRTWUe+TqXTcplbd2Dsq47CeU5lpfn77FMCt5NGs5HaF/NIhWdRN6DjRFAf4VGM
tURePbXv2BuJqu6crEeJWzEWJk/MVPQY8FYeWo1mzg25Ts68YEhN5rxPTtK28bxn
3VXcI5qKjl6jjtXEVDFHMF2hXyVD/OQ2vtmSh50rv5MQUmK5Ek/yAvs9YUH9RgKC
pQtlg/c5CFad+ej7IhwrQ+zWffReMoEXZaJdLhyUi9i4Jh7q4BVdXNQRcufy8YFp
bJOCgQyKOZ+AGunvjF9J8m7a33Ga0V94MicgO76BaLe3wPhTZqbMRs5zA3GYT0cQ
UjfW7DKZi+YDEhCeqglaj9pa2vj8Z7X0zQ0/JJWBhw4CwEByIPedSqTqmn6xMJvG
jJWkw7Giua6gmfL7zbqLrYz8ClJtmrU6gJKA9F5yQI8/DYdXIZ+pGkZCzT20j2bt
ifAcc4C1lP9Pu0y+dGMremWc11XWdIcJRRp9ELE0zewMo1/yZ3ObzPz3l6nSPClO
wtjeKPyWWVpr3e4kuPw7Mo2ziKtA/d1it99qVjkaq6RmqCVeLxQIZmKOZlWbGMNv
k5VYTTNGYtI17nMPiMMyLMW89NCdquQgYOHcVGp0CsjUlBD2YKbsk1LhPG3xfpvG
eKl0BO+iR1JTSUcheFNVM4uV940cB7s8CQcmPVhoFciCNKakcWGi5bM3qT69zRVU
An7Jj0d0dpTQmGje0/q5uhnuqqTJA41hHHxwO9zcpcb/FCi6JgNXWsFLIVJe64Ur
6JjOyJkI+kPRjPGXudoznHruFzbxto0UxIi6Fw02r4Sz+qXJhOXBfmHjIPdcQ+iz
TxMkoWaXgj6Z9KBeCtoRW48laEaY55EjTCbyW7r0RLeY82NNawvYPOYziDXEgvEt
dwRyNyOV/Yp5YBDqFyKOqBc2gBgZ3EpZgA2Sc/mGQnfQLcI2vOVD/6JHvLj1KSh/
Hg+YcI9zwGLja8AASSr877GL5HuAGsVvzbpRj9D6zRKttvfAT5RuZm+AwZucOWek
n+KCDNv4BxtIxrKfYxZT5gGu17uBLNJ+YeZUFTEn9Y6+ZgvydNE83DtE2iqTvjF7
obmrY2ZpmEWcCSxXRGGihhAWHIarR95D/6nFi+k5ubQl+YRO7l+w6L2piDLSzFxE
4/xby7qk7647NGnMthpsYRE6RtCv3QYfiLB6W7CZZ4TjUYBL9yg+Zq0sWe3Eod5c
lL6eXpejgfwmzRwRUZR+RIk8PgDTkzbAkZlvfYETuFyzJaFuJyiYgys/7vnwKt2+
OcUZeTJ7e9ruhAM5q147xhPS/9rtQoPYdiwhut5Ursj3Tyqg4YkfvHWG5auFOAVt
O4exSn71t9wA/wUTkrW3QelvF9fK7KrNIdHbnFb3CV6hx0iA1ndswyU7gQ4CqifO
4hlXO/wWLUe/LCDuGTG6rpkhefKmIMgRS3LUZoKcr8bBOVcVmxVTTURiUART2cE6
5AmiDw7QDIv21tERdAL3Jkt27yOrRNYLhsqr8/0nb6z3E3/+EWSaTCHy9BhAPdo8
tPu15Sl71ActUiOiOp3Q/hjtr6anlRToyoGaETZBoS+G+tMtJQd3wD7s1DnXPBS+
jb8VgNjeQpIsZmohrx378w3ulJtVAmlULXTyZD9UsI+oBrWrhtfQUGvxB+lqsC80
By891kKb84gNWrs4makaJ9PZUmQL/9sVTiLVLYfdlBn5JT/jBOr9hAhm1FC2fjjr
AnMk9n3rhOKNdc0fmdHgPG2lslwBPY2MpUiQNgtbJWbi4+q01auMS/5OxwHWfuIf
JqCtN/mxuu16NJem1J0p2I0TknhRc4SMH2x3RUt/ep+I8dd4YyeLJJfKWJySCCiP
2HIBo555dF2+YwU6b22rcEaZiBT5JEZHz1+lPHRNlwe+zjHaSNmJBdRm0CatPT9B
rpeprJskvlpF7GC95waf3Xt/5SzlYdJr27sODMlfrdXjAUG4Co4VbaBYgEY6CeD+
LSv54qXN5cAAX0OGelrAwGNMKd5Jz03qY+h+qzVSH24Aa2BaYx5CI3hOyEqexogR
TwTrj4MLprzBMcj+y68eJK8lO2kRMZiOxCmSEWUfIMQehhnCrbxzfI410y+8fza9
kaXyosu9UwwDS5UFY+8u2okAXJzJ2+N/TLUG2kjVtx+guX4C+mAlClrsIf7m2R6C
GGuZVz4vR7onawrRj5VrnwlL4BIxLzUc2YW6vwfgHRsfqw7yom8XGPuoAv/kGg3x
wPCACbuDDdXoX+B7J8j2SwFe9MnKfpavR0WPUBEPy4ONxlgC8XFBaXJe0fOWwLzl
+48c9t6eZLipixzUUVzveMgTOb/AmNd43yWGR2N14mX41ZxGQkbNbJTqsOldz0BF
Y1bUr1gYqxjbdWxflFAjkRWRmAFJOc8zwYVE+4dqb29muK4S/85TZVG5XYBetQNQ
ASnsHFvUoj2xKPKpdZkAnoc6opHv2aUu9TWD3kcQIufs6VSrCZzSZiY9Q9ECoLWI
+H39ojDLdYYc42AhfZs+dCBAvvlUGVbI9yB6MZx47gqqafqWTsbRNwhdL7zIzdVQ
EphAk0DS5J4iv+PD6q0HvyqOUD88UMQ01FRyipannPscwQPhuQG22bT1N2OxhkSn
0FsumOy7zd+fQxjY+4fxsO/cygnyHVcUTKhATFqgI0CrbNt3kG1ZXdsUUtPLXj3m
9oHstDjFLajDOT70dBNIcYB1ISyowk+KZYocd0xCBDQmt0XSokQKD/v/tJ2DDf4B
7V82jYf/M298+xLk2L8+eafD9W1tFn5Mtq3ZSfxAvLOQHMfGge6B9CHMCrmJRr9r
BB6iqkdIHkiGGK45WVwvVjKOclvGsD6AVLQU5e8PWVHynfQJhzmK8klF4fVUovBu
xfRibn6ZZxUjQqB8dvwkp/qI4wCi0lJF5Ywc806xAwnm2WTdtbmlRvffqHC9INRP
cwkO86KmhXCGyNDnpdiVTvNNxyCAfj9+P7CtQwTmkpMvT8TY8VOn5YUxMmhA9pfS
59FcIsW3J0CKD58hBn+jgbtfl2sTJcyMsRSdWLTBAIptHHAUEKsOqC/W27ZHX63x
tiaIjS9aK6c9CvfIs/GvqtedYIlfpFRJhGHOrGEvb50U6Lur4dhRbGPWzLWTpOZZ
4aD9UuqJrWYlKTy2y2AF7ER6mqvqNRBmw596vAOf5g1EuW2TFOSNfhiuVG0B5V9J
8V9ffwnUdtT5C9ObdJnHfcqqBN8x1kHBpjw76T2//arQYZHRMQpgG2f2Phz4NCNA
0hlk84lJnvbQ3noEcSN8OFm2x7LPdDE0VqHpFX+MRsoNEuUg6sTjl1IVgZ3MmX7O
eoBR163Q1oNpMOUgCfxTZ3P0f9ZdVjOLB4Z0+uILdW+rmeSwwpCNP8lwJ5od7tLs
mWsoZiclDTBKfZOMTTVzLg8T+8fZtexMy9m1lTvujiz8XEOwhXpBpwc0/E58h5Kw
ugOdJ8/JwmQLnwhi9rr+StmXcmPTBUS81iIFsEDeIkMK+vYetEMb1IhVttbSPFUB
lJ3l/TS3vi/OK8qzBtk1IPO7D0Odm2kmoULrNpJ5Af+O06JuMth7AaqV+6R8yJbs
jxDzdoeko10aiaAp9GHfHMvb6EZVix0JGNEwYlLVAKhR3Jq9NVJkezbxXEwMhnQg
kEu0Gjk21HnruU3cvaNjoqdWVFc0Bgz9RXQtkEjjcJhLjCAewcDIl8oX3datObHG
Fe2RG+qcEJh5o7tiXgbaHZp0R91AeE5kN5/Na+uL+paLIlMhPU6afiMa94fjs045
9it8mQzsrj9jaAgX9AorzcXcBgA3PdE2lnG+xNYwpJ39ycYKw7Nl0uJGf0cdIE/G
4ZcdTWIxAJPYjzKRJuDQruF2PtjB6w1c8JdQffUrbPJQLN3EJBEo5iHFReQCg7QN
ApnZWdpu30SxWF1KWk2ndMWoRAdaMlFm4gzsRHnVxcQJ269v3ZdGROrjm8/5S7aA
0LHQVhx22h+ANCa49uLaUYDFyGqourTllnkCejt8ERLGN0dcMWo6UPYVlTKK63ZE
tOn5/NpmK7pO08JYTUVeisuUNCki90MjaLCmtutElXo8sCsvc/cNeMJPHDlT2r/t
pVdfeIFlXczNhGeAtRHoNqxJLAGyCbMKEFxCUJEVovx5PmrYE/WoKGwEbEYhPhoZ
ilqzQLdKUGo+HMnM5jhuy6z+NPWSeyxiS/QgTEfWjP1I+kSl5lVXLkrRt2zO4s4M
yu+PkVUMbGx8tnLPOqbosWJ/vLtPDYlU+wH1HyW/8JXwXRDHgfR93rFL2oe/XWit
5ejDk+/RkkWteL5hjhAzPkp1rONBcCRH+F7BpbVBSPXW0NrhNzct933xTfS/SDfo
OTDxX8i3ALJ8QEATs70BGEbcKGYpLda/VVsxY2E09oKNHmr/Px7h+JV4PvsnMVNu
zMsVVvkkv2OHf4MQKoYEfwpmwff+AwFxRzYF1wAdi+QNbzfHZFszPysWrJv6sdyC
+WX5gG2tMvwnNy0j7PsTHy0dDL0S+3LdCphw3deEptEW7hPti+xbDHoJ3JE3DeX+
prx5hUc+1tYPzdK/A8LUOmv6pRJrk7mIZPd7mUkIj0/URgDBV3/f4mTdayw2rvEB
2rtlJzCqQ9o0Dv/EDNNfuQRHUwUyzxXA0frLYZk0OmNVK3vD0k48qTxXEXuTwAmd
KPrtZfOrU18deVqsWrqXmwvbfkMt5qYuL129V5ebsJEepIdMGNIWABzr9ERd4XAW
cXjbinZC5X10Y5BvDz/s8TDln4PE5d9sgxGjGuKD0gn5B8qRyM6EIGoTbxnFmTFJ
ExLGatVBQJcSrIERnBQTerZqYhuA7zV9lbMd57vCa0KNoDdZvTOZgynob6sW5HAw
bSLUcMB8+sRdLVfFf8XxXcS6C55tA19Nbu4cuUBsV4OD/UFv5FIocTPBOH+1qP1L
50TtzK6lSbr3YrDwsmqegrPC5SpN/z6Z0OS9FaiQIirUgH2qiWjSu4TZEeqiJprI
Unt2H82Eq0El1JxFPA62kRRXFYbvIupT/Xi9J3D1elU6s6bAnyBv/7pSZ7vfEQNE
JcJS0lsaHgRuqLD3FYK6Djufc2bujIUEzBfDiGXQOKcsFY35t0tgIFJp4FcIHanA
PeKlEdSLREGLZgWIY+wBc9GpP+zi/AOJvT0ZGyZwtfcMoKjfTIzCtS+eKP8h6RDJ
5cQIZpsmoTm+bcAetwel/O9k8SdPm99ALE6r62AZ1RRPJYtBkl3S42TIs3PsUVlv
nU9DMlwuc36af9t2ft6EQV0Fv+t1A4BKS2+r8bZF+fyKl89/5CmTqXhioEKTfm9G
v++/NUOmhd+zwv2pyERcSq8eh8g1kaTe3VByTrrx88vsqJAGZswivAIjYp6kz8VO
Z4eKk92PTL7yRhTcbobPtgrWt5ROmoEcPqMXBrv4KHUUbxjYHQXlok/A1/d8hYog
a7tpJxBmnwlmDhtD8dRGetmrdsRcCZa6nBPmil9xZLOhL012Ac7GosBi9Wu1ZsI5
r5/A1csHQQuIknkgwvdq/+hE/34R0smSNXmLToA6UDUvHHGgdth4uwJwPhzK45+E
5TprK0kE7WS6ZtXJqGAhuOGKfYPAwu/9gV5L0vtsFtwN2hb1osZwvlVejobXSxBn
FnDFXTcoI75j28HokuGqK6Vhf1EQn8USHc0b6f4SZTCWtJLhptfnTw2bp2w8pdIg
DQlHJRDnmGkpuRlALzD6Plv3CQmllBzU+OLgYdd6/2tfgWfH3ucndMa0XP73nJoM
oNZC8ml37WktyNSaFlU1QMrNXdppMNCFRJuHA/L1h/N5v08pH7Zw+CS3KuX/kTPv
l++rBKSazzjVXDR/Ig2LwdFkweWmbmqrl8xWrdpuNLDu6dcSE6qb57W3KnaDcbzQ
yopelOLUqAbfHiweHbXa9wJpCpxp1jJ9r3n7mP0COLU8kaGgYHLYQ2rxO2U15/WC
tfP8hgt4qEreHvG3R2aypLU8wfNE5l+wZ+eni8LAuNOzWRhiiw3yst/sxUu0a0G9
WEWuTEMtPMlBJhmjTAs39MnnY1gP0fD8wVKs8hAB+yR+1rVdSX8lF54VbZ/DhMch
NVjhGkDABCLt5AK8nZ6/gPwHGeAR+73+10+XcHYn3wxCA2LvN2WJ5cjo1ep7Szed
v62T5Ip7W645vrpwyeJX46U23oqBrKJFc4IO5henpEJ3+/qV3/JA5Q2gVylh3VCr
RyitiY9rrEbZPXU+JEPikjGOaNXC+hauPs4c1VBRhAqsg24VL7sLurbhgA/jfAPX
HUVFQLoJBskEEynPXGW4Uu7UNM7s0pNhX1mSoQE3DO5qX974MfatxDy2tHnwPpDd
y9hXNgYKStefdkChE19lqB1XL9KLRjzQ/iwmz7hY1azEkTqpjy6O5PEL/xvlEeKp
X/cZ0JTlWc7lmu6jRHSgjm8W7kcC3K1v54+MVh1Q4FQSimM0rnr9Ousspl+zIsF3
2pOa5ZOCVOJti2bNQ6hy1OrLEpsjd6MOFGCdhO7i8k/b3Nj5F+UDbC6+JwrQZVqi
2cJoEM+MkRue5LuFPxnTWNJnwhpEV71DnQXG2QpXY0gLlwMELMBN6imBbna8QxwI
hz79BtSHIwZi3qJpP59QwPbtKDPk2Dr0y6RChZV0eFqFgetViaqOdu5i/xzQvHMo
JNP9M/MvhpX97R/LNYow13smMyLbiL6ImV25n5GkDAZG6rP37WOxF+x/LOgkdr7J
QLcyZ62O+GDu4RIut/tAnknzhi6Fcn3Io+Sre8pujnRzEIn/bkRmlRHPk28FZgoF
CMdTkAKuKimLibOirhc02l94mJimjktpQnid9Qfh4BGwOUnLkWbNf0R6jkRtIxxP
qu0apc56npRpXHr5m4LjW56krVdfxSswQml7Wv66IvtseKhwWP2mCSfmmcP5T8DR
kaxhwKXTsof7rNiI/P+k14XLOBICkFUVwTKbTzeKPMbrlJ/+UL57eKBDUN+a1EEj
tJszF2sz4t2d+3S9si/3MpTKYABsWH98GSiAu9L+fg+Ahos7ktpe2L1qTU0yd3pu
fgWbIMOuL9KdhTYWPx3Omh06RamRqw1uNGWaetf5ss4gAwZcRm/ANfJ8hy4hlICU
4Vuh6aZTLlmGrGQt5rSxAC6QuUxcZTXESe/WyKf4pwjIiF/gfdhlSO3JxlOwUq8y
46ltd/+KkWr2s+yQLCShSp5xyGgMat31HQtBoO0mK4cptvQ3KeNvOi2tzxqatZlZ
nn6VD3nxHJjrJy5IJ5dGEWeqIgpcHo9UbOTJajoIdRSiznF3kpwgw7ACDN+SrGcl
KOg3L3RWKq6aGjmuMOuR5PDUpVPMDp+T3qJ+yCaLbMIVl1AxX3SP0fNHX9OaCT+2
1RvEg/jvHhF3GLeED1ox81KsJfI/kwZSt7qltkeONgQ/1B/NAgeyTJAwt/AwHKNv
Jv8qqCaifZSC5n9dnn86CZEvxEKLLlAZNmnzYXI4eDl8ymgT+fzURK9iFCAjuFW0
9LZlWaiwkNJCrJ14i5L2j39pBZiH/pwOTP96JxSjT57JvOg9H6pA/BWdyVNCEQ2O
CL4NFXHUw9LU32lZh/C+Kr5wsEnY9CYt+zwqL6X6nBQRdKp5UpGfr+QiH4QgEJbl
YUTvRSVCzM3wePvAjUBlMBX3ej47cJ0jf3qfvriraJLTNQvLkvjENPE1iTFglkUC
VSMxFXt3h4rvwjyDo5g076lUC54LpQOLI8zZ7DmEyac36f6/dXYNHvgg3p+aHtus
ZtDPT21gO/3f/nVjmT5tRW4mp0HpJwaks2ThA9auAmJuZSTMzROP/SeT0RkdGwYi
YUnnSDEDp05Akc+eggAB5v/Ve8BCLHS48VAUAXeN+1cP0zi+Qg3Ca4K4MFgCcFyM
3FRgNlxgOsAlx24XX+FHH10tdT60yZckWqveVIvuc9+h3wWgwWIh3tdZl4ICUucx
2F1BWf0f75Ox9w3BXvrsXDW7NaFg3yF5llzj2rpuHOq7KBaUroDh/ZuDMPognH6E
Xug2anqMJPSi0SHckebuOrQcDpGRG2F0VYg+tcdsQKM1oeE60kMEkmAxxjLPI+jT
/e30cfCBnHvSHEsgJDvVemY0Ley4ivff/X3HVnkfEZ9Th/yxsrxSGuVw6m46PMg5
Qn12+w8bl5ONoKZeGSDmvS2hnft6Il186Z3FpSAjBrExS1awlxW7nij9QZoTJfaj
vEpOQL/32MPnat8seT1mqZVAYgMwF3O/anFQYo3/FTYpdqXvQclWzIeXmN09U//O
uEcHhjYSrc14yNp1eQK2FBDItps5SghPgplrRfX+b6QIGQM/jcmFOcfoF3I1Piip
fvGdC3WNNKuKo55xEDyAw2+5G/KOjubu2imVS7n95wilnOPHsnoWEg8VqBME04a+
v7LwZKkt9fnOczqneHpzKHb9KpcgMJRC5ZEhQzX6P4NVqcBi0CVynZO+HAMSYRkd
SdJ1BKvOk794cyIoXh9Am7+weQP7HahDMTJ7ZIAvZy36rCJkddzTAV0AJfxY3m0O
PQUldirgx0KURK0KIKUKkDCUjY8DaELnwORlhZbXa812dPGVsKIXOlY8vEUTCq1X
0JXoZyLuZdx+8GeohrW/HPaAb2ZqRIZDymv6LmCiGV1bz7fgxZXjag2moHPKHtQX
w2euL1CiKY+V2tERL26KI/wPPBpBpSSF+aMQzelKHbO4Sw44u/3I/93UOcvWvwBG
VDJ0ttAXOa0iabhM2WGQSNUDv9S66rVxkfpKN+ers195eV8aQAitsqdqM69jw9CY
qjH39m0eEdccDAFuEumRuPj5SFu94x7QlUuYw1GVGYm1sGZy8REhi98xph+GILFr
/mipO0Q7xQ3IWYuXU3113NafOI5CjbPNaZRIrwPswzBntYV5nlHEncEE56RMgIgQ
9BBiKQi1fkFgHkwYXXStZYSFVSrLSKPjdGKd61yMmMkhS+xN4tHpaNj5AL5/hciA
ArI/xAO6bXIAIbLWXEB33+BNCf5DvTAdbxM/BundcI9CE9K2nEFAL2TLXaMwGwNC
V3Bx/neEZBRKFKYsE+ye9eM7FAb+RpMJX7C8QGFr10krWZZ44Wie3Zc3X/mrROgI
G5+49g9wAs71NFvpZV7OvHqk7jW5cx+rD4w0Kod2oBVKbW3Klxztq/7rTGd9zKZG
8thukyBzUmJYm36OkLicdoGPG06UUxpN8Cu8w2uAfi6eOA+R3nqMtkTBNAxtUEBN
Az4vbSMOojp47vFcS0euBhFgHfirAN8FkHtC1RUS7yDB05tjNUKKIYsfUVzicJZo
ud5ZR8dxKg8yd1QMLPkKz9Vc1hth/LkZS0XNntid0i09/1DB+Wk3Na3q2wbY1qMG
ypcllbbE89Gj6uhclaXnaY2ZBY9vrS9g5LOXlEF+aIFTtGMmUdK0o75E7VbFnEHL
AYDrJv1pqtGPViZYOOZ4MqXPa2faDycZReak2PH9T3d5FthjPUJUMsRScTFt30QG
f8QWFvv7vmd/axi9jmgqnXusQpACCOb5z6AOqedn7WWpUzg83Gn/pWhVBtbRU3Jz
iuv8ZatH3iZ3lhChSFTzvnpTWa4nSxvG7ZBgF57n3uDCjaZVV0bZch4id6CWgg8M
Z4BljVAQZjl33n4fCm7g58qp/Z4PTICtq7GVmJ8x5k9um5xmx9itbfY2loNG+9Im
VQ7HsSSchynAllDELYvW6yH9X/5CYaL5lXtbpuvcbm01M2VvH59JxamQLgpLJSdZ
juM8XRlkG8A+5v7YpBgBYt2OZO3IJld25MtrrrHAcxOP07dI6s1KIaQFyHDfERp8
wKEcaxiNr8S1C4DsS3idY2i6aEU7ke1hYvp4MnDxKE2pO6Bg84a2Ty2T8bXpT8j7
YqAnGr0DuNBXKdKn5noPp8slTPI6gmLoPdMb9GD+ETNGQ8cVLQLaliJlelt3Ozt3
NRA+6LNKj3jpElMHsD0KvrdyFGZk8wy51NPfV2IUJhOUZEi1PSgX4fzF9zfuVf9W
zSVBljKvd5W+SD+4BQSn2Iambgv2VJ3927ZtsNPl7ArU+YEHQFd/aTMb1+fQymjT
iA3Ti7kU+5ygMZM0A3XzVYUNguoqsJS3jE96Ya2IACw+ZVrptYcJcRleYJp/ouEq
e8u1g6PXyZhhaeBsM49hkMFiUHzh//wsI4zv6Kt0ae7tTD34qFjZ4kGzoHOV440m
EvTXJW+FxSKgWLGsVL2E/u4o1tNNWNEhQqf4Fida0fE06tfLoRvx5LfZRvjO8w7l
RvcpE5SsoWRrTTkZ/Xj4GCuI/8QYfkcaiYxjDz22eMsrKkmdaxiggUwH5oMPufl2
xs8j6jLPg4z9uSP4Q8xQL4x7b5N7fZ3+2OzJAuURVCUPJXFC8gmeu7HbdAiURA8X
dwyU/OvCyvMg1I5k5lyOaxAacHzFc2/A+PEJZGx4ovfnay8TUwbgr3ivZnueS38U
sNkikjyM2H+6nDKSJFu8dp/iFQDQ00Omph60OOK0PVQUDbtcF6fWOXReNord1zBa
lzfOEGbctT60XnOI/YLsucHbkoSCEchv7dy/7c93wIc14cfnYwj8f5YLhWPowG9m
hZELvkD/tgvGqGeB3llt6Eq8iFsOIhKN4KCW/Jy+UvNMMS1feaWmJ/EQnMqFBt6t
3z5IxLHLXfz7njF92HpFBECVnnIvtGOzFUdAG227S7cRh0kW0u1FXNBDnHSIad/k
qiR8atHoAK44+POOttyBFHBGUOQwpUTSPz7h1SJ1cvFCc+pBEpzgCOrypRQVK8/L
KcYSMWr/PMW14hqT0fmRN2e7RuUh2pFiffYNlxsrj+ntNkMYH46WPAT/kZKcLOGB
CtFMcJ5JoJpXQnJqRRbkvIyENmwjChsRt45IgS4cY23Y0IF601zEhR0nBUqbOL07
jRfKKVPZXnX1EDygtdDtjgKHr8JLl0bjOm7QvoOHD7iV+8gQ0BQKUYw9uTXEnJ7+
USgaVQcokeBq5Gz7FPk5bysrJXw56j05JYEzpz3F3G9z6dVWkXyux6mvAtrsYQh1
MbmVA4Mb/JY0SP3sO+PMXAyB3BTZThMGg5/530WtQ6jiNQkqNsyvbI9SmA95BJJX
196QsE573Ymw4+IghdVGtQzxgBmnld/UMW45bazhsmICZ5K3xYZVpN4ISqmeGEqC
E/Pta3D/vJvCX7Gg/G1bfneIU9PYYxzqMbYXtR/V6aoTHwGb48zZv0WbpiQlqz8Y
6HTJSTS/nDzw5RI9+Guleg2YMKRsZhpuNBOIdbVJNH9cXPyC9v3ON6lNfNhEHKol
V5hqd126Gzw04Tn000mwnXYwWiUJru2Glu1Yu50FUJMoR98Xs+5hnZrmqOxUFf5m
5UX1yefebgL3iG2M5RSmDMYmWQs5QhaE0DIJzHHqgAUUqnvz43U8SIybliJ5LFS9
o05GSNf39sRIMLIK/clF4RxvX93q6san9J6DvQwqje+NIvmWCrRD+HOZJ1ZcRcrR
d01XB9Ue4NLHfVNUfJqOOFl/uCr46dPPy2jJKMKlWwiT7doqDwTDkImJytKCQmIj
6oyEKW33u4b3LWSm7RsM6DhplEi2NosHrhIpouFPQUv13KRsNyv1sUxs+csHkInY
U10Hzrdnru43b77C+2OSZ7jIGhGKM5CZbaWqW4jO552zVAAOdg9TLn90j5OzCl34
98a6gLnRaB0Zog8KthwGY49t2buy0FkYig3ifrHNiL0wh+Cl/vsTliUDQ1NUm3+P
j10rBoF3g9b+WwGteb0kk8u6U0ZQ54w0R3g8Z7z56PLEmP014qeXzMNklz7LsSFb
/OI7GgKl7voFpeCqiOdwoo8sZM13LZyqQ8wTVnRWGz8jldVIGAxNeG97ReJpwlD7
qmmRAqDND9AxMykt//n1GA+CZflLSyN5421tui/pra8DkM02ALRSHJM5Hehd9IaK
ALB6hyNmE92oEBnmlAqpICF6p3Op1dwOmvIfcy6atKKh3JgD5sjeSYq0inWCXrjF
AMAZtJ/a9XWHnJWiPD/NL/PozNx3iDBEAm6feME4bHYAO0aVvPLXcZoYKWpRHUX/
w+QA15Rw7n/Nv59iaCXpz71yup129GI2h1mX7qYIjNaaFauo+7azPhsn+ulN/F/I
9JHaId98sYljcX6XpJD1x0pl6Ptud3qtzRvFdHsGBsncsdki+SrdpWaa0LGU9Lr2
7EMXIsWt1UC9t37ABwMPisRiAVZ77xrrcYKZFRfJNV3vBFVXdoII3n7IqVLKFOfZ
fotWCnOok3t0Oi1vW+pX4T0EvY++flz2jlYzXt4Mb8g88xH+hrp94XR8JnjGQnBU
JGhT26H/GMkTeVSusldKJ+wU6xO0wvFhWadRJa1n52NfmTUADSEZzdeCpjkqeVkX
y1KKLFEbHxhTJU3GEvC4hs9R6338KULUNS18lPG3kA5J+TMt+auDF9vDernHTZjt
+y8qzRgVzdacx5r6zInBHd45FbZMaJ43A8a+nHJVPv97D9r/4MZTeN4T+vt2carR
YJAJmUjVx3TZMZaoRVVsPjY1WHUsEC5eZQ04gVGAdrKakMxI7nqMjW49VJPVyny8
xXmcJJt/JCIiAHnlhEVdyfx8cGNuNddl5Ux9wKuQb996DkUJUKRcTKxQ4LT9V6Xe
U1UoBAdj6RGuv02VCoMHK6Ebz85uvs/c8DAuW0xMA7c1SIDawHOFODmVJ2eR7X49
Ycd1oNCacHvnBjAOTDxgZNrlPwJLzWob6hSVlj3gqQUNmL+Yu5sE4QhoqrRrcKjZ
2XllCxCluRQHHI2nMQfHd2gHJ7+fnK+LrInZlfvNhHCNN3L79K5JfhAy9Ljyprmn
kl8GtkgpPe6IeezQQcUKI6naU6jp2qFj6yxQVxS973UwFjS77kcGLeUSJbSBWQur
+g8sNbuGK3lbLjwcdS9/xuiooPbV6YF67CUariyX8HjuWC2tWi28UYUxJCm4fHLI
WMh1uBzYxi+STieiWWflxLZtg3mRwju8HbIMubnTQ7Sk9k4yRp3rytNrKpOeacUD
cxb1sjsOlSgsjlq8B3pbkCnG12E5XQ29IJwcskXY/USe3cy4YcSilKwk2gywiCYq
Rj1zqYjQKE68uzKI/Kp+osUsO6unKJOC+e5MNto2Eka+56FbXw6/L/1AUutm4VO2
P+DjichfA3/KB0uNHnfl/DkU80JFZYffkxXlLBHBwsVlHHR5c7hLIVW+M++l3C0G
kKCxHo4kB/wSfyjAMMvWHM2qMdlJwF3+ZhJh0Guf3uWauPxNkcfh7iyO/9peFf8E
6y92SBeHGOcazhIgZn0ExQOMhBWleuDj7GsUdGL69FGur68tMogsicmtkye7meGm
WvGpxeYAzkqyffnEwDqVPmeZlBjrvPsj3epHvja6kbF+tBjMFY+vKsN3xRBPfAPI
vGt/+Bj8btLnVJHrSdRPpjU8qQRsgPp14cya+IVZq/JdCueaD+72VwOQEQN0Z0hR
xQ+QbSZJ4s9d9G4Y6wGuLKlTCgtPpF5mmi7x1zImzFez1sLubSa//+VN6zj8RLKM
E5m0DYuY9RZ5/Tki1YnCBLjZxdChu/lM5QWJ/UZiiTqC90PQ/03AA2F4Ue37EZq8
P7INBzJZvL/tXrTcojhtNFm90QK1KLlIZ+hJsb02uPY/OrYGy4T0/2GGafeypRwn
NYH/7kyw+1kCkvzqUrkqH1upPnMDQGj0B/A/EudZZtTCB5mLRLEpeKKyQMYrFzoG
TURdauwa0HemFdh4Eg6zAAbUrRZbTxl5WNkX4ngb4JkP2t5gVB2nUQIUR4MDnPG2
YBhTJNgF4dFq/3qthKXaswXrBoqnmplRYQnUgFY/0XTAhxMqOE/8OOm0Qunt6EXV
qEBUCM9uikTNzLgJXMchsOa7hThMqjCsHOX6vOyhRgL8VbPht4dCeBfMG29HzPUT
wpMnJbTheomo1YMD8/Ve9RcCUP/6DmQvISSHv+WSGn2XH85eMaGNaG/YElEYI7Fm
K4PvaOAzwiScZkec025vkz/3YqxveVvtebfbhaKxCY22Y99AsHPHtFsa5nhamYgg
Jzl4Ytl9mzJaVZpRn48gLp5RrSp+wY2n+CgCCBUvAS+CBJjk6nvd5EZgaooctYK+
WBrg/RrY56HoQDuWSsbK4weMaA0W2gTfEB87OStBwEhafKl4//OQTQtIDxSR0iIW
OHmBS+nY4m84IwDlpP/oD/wAXMD5tmcrMDD0xxEj5nXnLrqMcxA9bVpiTuujtJga
qxTA4s4sc6afyVTZr0NVn46v0yrUXvvwQClSoMDwHh10x8fHKooFY7jltQ3l2L7F
95FKOCzGR8zmV2bMxnI7ab3Gkrv12poBrD+90bYqYPTUpQEH5RMqWI1ruHkheT++
v10d8JTmffgB35h53iH1LfcJIJSCbK/ubpc0IQk2iXpXUV/aKqU4znPOZnEvvXGo
W06XVOEW9/jL3X4yuWzgRbah0US71CMx3+pLbyLWNq+YdGwMYFNj4qPHpw2fESYL
IM7hBfs7BNVXf+EKvb6QaStVm8oRPmlYZFp01f9vywnIcur4oNA8rgzwaX3Gk8Eq
JU+sm/Haxdv4MlWOAfM2/MZjTFoQkaE+sTX1WnKni4k1bU3UFaY/J/x3lR21V0BT
L7WR8wW4GVj0ZJJuWkO137XUKqYvXNtXhNsDe7Hj6A/CoGTPc+aogoz9P0ZqLXJn
9CU4ApkmmO9OvCJ6grzNxqIH8Aklho7xyb8Sw82uR05iZUaTXak0KugnWAx3TieH
PHonfMtwzCY8q3il2i71BSIMrEX9hIkvZzGcLy1iGyrWRZPnjK7MMnBHeu47HoaE
RpgBrb1IQLC8ZxgckQe2YN/4o8Eg0vn3dkL1hqDhGPuGSOF6RitXWo/JGIEVP9+g
Won2brkDbkmKv7G4V/XAIiRZt23G5jtbwwWP2IlvS6EJ6hvwypq6OMXKY2Frxq5B
z37HKY7W6LwDTy3O2w+n8JxyeBtRY7FXFj0N5yfTlPwPGDLCRpmJ8pAQiJohHbIv
0v5oehRciXs2MlnPZEB9qrK6mk47A8PafYEWqvFJCgmpCxpialVUxhhEVW8u4fVu
aS8VxSg3iC8Er5qtKgq2kUl+HRnnXmLa0vyBk5GKHjjEpBDhM2RFdqcXTgiql/X5
YG9bjhuZKOF1mSiAXiCCf+C0GG7VjPhhkLGvg3bUnSlcJuMqSy8g5+x1lqWTujmu
iE1IBjPtxyCN7gGa2NKUS3DYa7zkvCqKZtlPMNJt6heRPLbqYQdtC+daTY4HPYXm
gwBPGaQwdiFBUJ5T4UIv0v9XS5KoOGKzvCfcOhLcWRl/pkew1z5GVwMaymZULyM0
NvYa6WAimgx1M8nfBna0OoKJXaBHF265Sh0q0arJTZdQU8VtCD8eLQBbC/excC8j
5RUf0XkrV/taCte/j3kzBc7FhOWy7tvqAZZEs0uYIQnHfJ2ArmjJcL+by5OUGuCD
mJpGZ1cL7gxIpiopWFRYswODT0hwCXGZUmSvbTmBLowemWGIA/p83hYpRs3jKGvq
bde1lYYa50lBnZthF00nfDZK1xVqMzNhOUmR9OtfckIZxmX9qYUFI4+gbHfirh1z
bwA5+jOkXdRAhfkEy5iji4+R3Og7xvC++u7C9hP6aSBYPvV1wEvFrS7KkOxNfSGk
foh8M5Af5S9/LSJgWY8/DDrpWDUz09az2f7m84Jj4G+dE62Ek26YJPC6m4jx4UC3
SRJYepqF97a+FHejsgXHlik5vA+HkrfbCwNnDuXHT/3jK3EtkYF4+5dxjk6Bp85b
G18B8kQA6YY9J8In8pX5whJ5DuQ0+I8rcbxjDSvHNDrboURviJkIX+K/t+B9MoVp
HeJg5kLuSIVGXYUeYT2K5BnPH466w8BfXWICXsGbrHTGAWnMNAakMo/eDKAVjTVm
5VAae2klksg8P2kio9Wszyx1U2w7ZelShGibtyGW31Bo0gBPh3RS4OENx8aU2MUm
f/k4acEPaKDm/50IHm9kpFqlXu/jqTZODdZ9KutmyxQDJEQYh4dYIe2+PJpvMuTK
oUojRMM4LMLTwOBdQ+86clkCO3N50zfRaNIUV3lHoF3W/ozqOfJObrdR08K4JPoE
0W0TKYAbSK8nJO+I12zqpdJO+mi4q+eafPPsKuyvTYFTFwHRcxbxZNMet6ks7KCx
BdcoG/6ycdbuWSSu+nqnr4Oupx2sanOduhZ8pj4DPH7GC/cEP4Lxbt/YjGBJlM72
y0/5Xgw6BHyqJbJb/V3FYu8oKF61rgu886Gl/giLyLmqndW86UamlZtFsfZplKe2
GVkQu6eJxnR7e01Pnol9HWRhyniKJ/ZncOQ0N8ACNsx04TkPSuaOuA+2G8g9+qeP
sbrcYKUcQwyPeICMeQpliI3h2sfgoRWvErxeDX/IUxplZioxxgxE7MQCh03U6l6W
BkZ0ZdfKqSpHo9k3IKaHi35eMxX/6Me0wvn6V3d7CT87cBRt4lbBXLVWQBh5uKO+
8QSNBTklid0Nwt4mmXC+jbCmIJhUzu0jSTCs6WDBJf/EDmrsXtuBSbJf25i2agWx
QZzTkzQLWOXXEhOVBgK3AtJ8OUJ5irGfx29w8tm9Rv2EDQDXLP2eiFaEDnC0OVYr
bgojPWGrkWov4mRDZnZq+b4Hk6CEPbtZdaCzfZiOMoWCGxO+r2IRpQbEaSplNZmO
NlOhGk/c7P5wpjgA92Lnufpx4viKDo5nuyZzcw64eidIwX/Dy3BXl6qSNXmWaUvc
xELfTG6DzCMgb2VzCuYnwrk0205DVSBbh9oXLfF8sE30rmZwRZdXHvfY1/3KqaSV
7LaEL1kmpxU7UwfXv5tHozifx9WNX7q/3fyI0Gbs+oUH72+1V5yVRXbEZONyOwp2
O6hKNsm1aaaky6sjEcB+JatfvFNc22DhtcXtsu8kwXWkPjKDbCx4e6LtZG0MqR7A
pocVbHsatNfblIKJeuFR2IiDK46MYHwub1OXA2CwSYVFIL1PlYUi/Z2gXAAe403e
o9SoUqbaq7a5RZCpiDAcbXeN7QUI9/Wq8EesRIeEA1102+X/4CCXPXD4NeIJBtJV
2+nNdqUmUvtsVaz61mJVzvm+nJ2adEJBqijmb3oNXuPOFDRc/bhdLkRPbBJWc4uC
YGsC16ffGqQ5DpkXgpmCQoituSsGW6Bf2sotrjXvX31U+VXJiqHnbhf/zBRP5SVZ
2meDzCBcdHaCqVaDiSr3JJLij1p2i/xGdqW2eyG1J7gsE/AVRkZ3U32+kjuQfagH
r25rTHHvuDvlx2omYOADEa3nEOP2Hb8s0vdui//z0fSNWCXJGR9AGf8JFiRyBG/A
jIKDP0mTus2Q8Ma6tWMk4gwJhhToWDrM8B9GEZh4M/FjYkvPBTKpvn2TcPHG3b9y
PAFSVjqtKamYn9fGL+zG97A3zAvjV6wQh/O6qF/vo/SgT8a/owmTLQrs8q2XWhD9
B/nZWi345ikT/WvlwVBwTJdOcYTLYe7uRpnzW3CH4z0PqDxuB3V9/2AnSxJLl3yW
/Qq4KL7xbiamNMrH9fY7NQiaES1jHVWvk81YKj0dfyRViwII41n98DX7Jm4V+FMl
HQONMtO+ELbcDePUEfaZfFUKzieSQ97IucS53EUuWVMxEPC3RjrkurNeeCx18eDN
qOaENcR8vD+6g03CC7S0I5qJoRCoWg3qX+wgPHPCZiidhlwa6s1APOPfJvDgG+bA
beZBQDhUufxXZKG2gXBdUpySD4elPtI6GdDtHd46ClZSixdeOoglhgHfp+856JRQ
jTgaWnfkNcfSITr6h71ARrPkQ8Oobxif3jBqOvN/7Aoc6CITvIrOFtlmMINuBWwA
8Abul4WHa+6zoOH0S54EopnVdIT0vlZVQl1XdNFBNuXTlYQVZop1040ga0xbbE6Z
FBCT5hV+c4AB2KrSbz31l+mTcTHsZY4xtlMEp4eJkQHGpCZGhVh9YPKCJpmemLcF
8R34zd0lYb4/1ZFGsj7QcPVhEkJpxBUrmBb4LgPeL9xtGX2tkIPy1u8pdTz2fTuR
J07ojfyl6QzoH4qUitrAu+/xJ12LIrCbtcyWjuI3AzZaDzFIhqFcz+jcG8WTFXBx
aeowsVt5lxW05aSuTb50I/q+F+5GBWOkAHsGE2/qcCQOoB7APoGYSiAnbWjw8Jwl
0n4IpsXLZbI/U0uh1sG7xgT8KV9r0z5JHB2mTO8IgZTuoo9vb2A8aQJGf9l0dHBA
FR39nQSWZVb3rTRrf2+sqTn5zM6VYlSIAFcCrOegqxaMciTqwZqanlyp8rRxZ/H9
DbL58q6W+osB6k0s1ezAabWAAGX76SlSdB1yAuljbCaL73mDS+YX52JjZnD3sQag
1ZvlF+zaY0Fd/IQjDYbBvA0bSDLzbATGhPbQJNwdRVinUcTU0bNX5IJfx8vWqU2s
9rggmYc1LbJ53VcBylNJoMaVB5ClNmEDqiNnFVO9Znke9ulQLGFRSWtzCgu4tHXq
53WX2u17iBJQL6b7D0l5fxoL8jP/HGm4vHJ4klrWFbVZDA0+CYuazjR535uEsiEA
MAWr6f6Z1fdYWlxkEv458ZBYQYmamIMc0qFcAAGE9Xo9ouWgp5bAnA+5BC0E8ehL
HfbShjiLBMhUUt1Wa2FosZjz356+CdspN1lJ7UPGhRqfMTAtlxQHiPuJ/V7pUbc1
BrlvXTZM0exkL/01Kh3/9Mu/CwajodRypoUsqviCAh5PUoVrljxBVoK8No9jOeIK
VZP3NVIR88grAi2zhH94C60KoAGwU+7YS8KlgbygktRcuWZ83DPwcmDS4qS/lEXc
nfxvgWRZYGuFwpkIhS5jSJvhi5KV9yTZIrjLYU+bNbySbKJ1OJSLYDGD+QFmXuDX
96mt7elJbEZ4uDXHTv820XPMiU/2o0ZnGn6J9Loy88KirgaqIWGqVDS7R4ows15+
o9rrfd2EA9hrAGth+oF89D1xXE5JzG8xd8/NKC4IqnrFDLV0KTqY74uUwQ3PQ/Zo
C+55gE+rRsqo7HCmNBtWgDn6mwZDdNgp9lbBshFg2/xjZtbJ/IhwmGz5G+sVTMfI
sHSIh95Hknbpn71nlSyGJj+fuGMyQGmvxCHJIPkwYwkMz27WBu6qw71idNKDk8ag
h8izL/d1xOcTVaglIH8AsKksIFLkMHMz5Ghb3BbDDnOxOjFRWsURulEvVZIxvlv2
DfjVBXzWqlMg7yt7h+ZOSjbfwOhhHW6qed0pVJDPm2N18FimNeNwelZtmr9JQ2Z/
U4y16lC7j/R70NBvuHeKB8+5iSs66ynpbZkWO+qzmYcoSXxFpZBJCrsFwKxUQVZX
+n7nx8n63f05fKOaIDSL3Jmcbt4mi15d//M8T09+vcnXvThPJxe/BlFikn4say7j
qbGda+qqET0wr+iIWCqnXs1xiCfakrE0NVR3u8+7GkPZHr8VWRB861OdAwQkGn3U
MTpuHU1gWpl/A3Ar9xc8CK74z8Usws20EUrnAHAYtPJ9QJd3eFCZCA9CJABuwrjP
NrCh8VIjxhItoXOpRyB1v2wvP7zARnqdIG+19nZH+SI//klbTXhrLoD7BPaNzc1X
dIjpU1+blGvfRDc2rXPV0OfCUWksJcKqfO5YLeGpcC+OksBrbWCmQG/zn4x+l/aY
YxZZzfjiNFtXlZnibIIl1TVJqbPx9qiStpAAN6sTjTTgStczLGXAZdKSSfr6oSPt
1QcY1v/vuJsgzXLkc+JHmJaDVr9Ss/Foz6cmnp5OJJh6PfDylFfCm5Ozp3y+qeSU
VH3tFnD14fY/i5bi/n0dBaO9l75LCmXVh91m9I449us2rzp/uh9uTnlKXW4xS4DK
aCq8ReYNSKLbDL/GYC7+0cCdmF3rrLbj6GEb7p3dyi+wUpZlMj2ZvOC5xNfHA1y+
/ayDvI80vKQshiGGY0zPbPKvrDnlX1Av0kZjgePXsYKN/TVMyGh5NTFUxEl3gP+M
Q3ohiS2DqREn9dcG3TtHLhwv2RkLcdGdEJyOFFerOZSZAuOSe3qNju3ZqTj41G65
+Lt2rs+Dwv13LWsqwCB81Dw9uCnrLKLZI3RVgESCJQ4vPKw4ptsBiCgGuKG+XPFu
mTOOkAn7xCh/hQKlV9QGdPNeARcxNRMrRvIDX0thOB74NO/zEwhXX5Us5NUYATiA
mR6u4PrZBdO0G+tIGDjYpcAnuZID9Yn92Aqq9lGUM2jirZsEKN7jkmK+AcGnIEXw
jgARCz80vuG60V2wXtVmQqXDtBuuhOhDVwp8q2ZDYyso25u5ItxS4zMuhOC6IX3T
G5cXAfH/IuTcAtaOEwuotvBWEHXzHyrcIJSKrOTdIOWTz8Tq4RMnMyXMP7AzYcaP
vsBrB+nHYMmGkMf6StByT/64WMK85QohN7xZwLfZz6d1zVfkxeB4BYgKzWg878Yj
T0H2WBAE4vEH7C/YNMQViXjsON7mAqO7UilgUj3Uw+ybJ1q6TfSe4dnD5NTbmcGk
Oy2ymn2Ua3oUsIFHmbFbkAIYxKhBkt17aWUSoPSlUVLS7xxh/tqI/do8PESyViBE
gFVqRo76bcutIdTEKb4AsLFfRSyxQZZQqxAK+8Zgbee9u0U29nCSHQRMhofDoSTw
E19WX/Hy/X9acT125F62hm3GoSRSzfx7/NtB4enRZkv6OowkbiKu8szG9H7JgICx
ga0zKb1MGLvhsJ2NSgnlXnY1wIs32Dhf87PeaS0ds71FXF9lC+aC1sDF68SsnDJf
WBZ+CeupqCySOPtxwsX54umH7ocusnFGAM1PYN/VyynpYrm6HsIQjTH4+gdG2v7r
pWL1JhK16RuZZIiDaKcK5ghv/djzU5mPKlB79nxIZ2nPJf6jdEsH5WEzuAKG4uCY
wbeEYYhAFqs7qgO5t6KZ/fGPaknHBGa2XH6sD0Xgrme7wcdy6fVfQnlvOMiekHbe
ck0/WmAaaLjGwO/e45r7Dbx2nQSCY2ZKpK0bX/WxgLuUgbtz8YEWPWYGDZTHChY7
QkAze0bblMRLeG2uMmgRS9Y1kQtonKq89ghZp+FHP+BNlibrJkGRX2VX8qM3U8ub
P7Y132NS7OMHouLE1tMw6DFN//sIpZW4xfmp2/D2QzoqeqCbsUyvNh1VNG78nAh7
LZ5AHi7A9zDtvyv+icsXlBmUAdmWjkvfgzhmCutIeZwgp4DvP683OGB+uEWlcjUU
L9j7+PsP6wEnZkbl47BgT7iQ9+etDWh5WUGrJHmM5BLEZIEfdWX3GG8Nzgllb5i5
7JcD54XsyxsQ2U95NKK1xB6tVhdeCE/KFsRqRfH83svW5qakopKt3Df1mhKfbsK/
+oguyEBhzZsSznfs9+c1C4aG+my6tmm10p1hjtt/MAH39QteLv+2W+v38rU33QL3
GxvevpPEhzX5jjRWYHuhgqdniOcTTxy5WcQbJ3sXZAnoDBv2eG557NagW/G6wj6I
5gUp+cOBkkbcbVVwnREVTxHnYghbsldjBibK5juI2uX11Dg9QsHPUrJ78Y9WvJ61
wjijaj8zjaSVU91LbJ3OtxmHZZ29kQHg1KLtSTz2622UAsp/eydkf8d2UgWQlGfG
8eivmN6K1WSA7SsqsV0lLurhuGL40AwzreGbgw76IE6hAofVjo7koKGei0m466mX
tCjpo19n+GpyzQ0gYrXT41PENcgOI5ZW8NttEF4XUdD17NTU4tbw05Fg5wQyWJMX
6Vjj1yNsxEZhGvnuyoRrtlv4iyOlazaYP2WNibx+nNTqYHb0xsayAw8VTAE8vpqg
FSgtgOSbJXrADczcmllpkcG3cM8BUlg1LQpBaJ88UScPCRRCltGwtBnfWPmFmbf3
4i9qWMb2H2dPnQ71l8WybH56LlR/B9S36WN44RxPYlvsbTvEDtMO7cuw8Wybnr49
x7AwgE4vNyEj+obFdQToGILkzo0fguV6N1nHdT5rJrn4P6cckWSNiksjkjsBlPf3
elkpiCMU69+UJlOqfbKxsYZRsCYnFvzzWxlwFF15KyHBNpvQziVgdtH3ErPKcZns
uo/0jNESoWFsPuhGgfzsFyc+Z/ZjJyMlUGe9pTzGUO4gX2uUGlIBHIg5qggQyUuM
ai0+y+uKbY9meu9GNlSA83wieqSnuxFVxEP3sxxqV4sSo6Wv7pgdGKoZatB/ktze
VNX1/sJl3dy3WX6hxco2loXyxxKqc5qJUoiKya5EDyuWpY2YJrGm/zOho1woHR7l
inIkG8iVUbV3V2tZ0pHdPyeeAPcDS7yUhKnNBTyWwz6cX5MV2cuasZqbieKHmI1O
QOffA9WY1xz5DbHPRSFopcRCO9tMZDYt4ezkgfE9isjHN/Ub8EVMHgvX353kDylh
VI5XnZrPh7p65Pn3a3K8uiu0gqoJGxVsAkzhzDjMk5XYhSPLUBdNGGy2qEgl2lho
gfSuE9r3tQ30G3Vidrh0ZJwOjTRNaRtY5VP/vlYFA1IlaANQMls57OUmRl3RwTiq
TjwbbZ2+q6kIF1y/UE8oJ02GgDJszhv09u8pFmSCgvRfR3dlQMtCcU6C96Wksk4h
0/J15f/3SPG8tI2JZWc4oLaaXXG9AUfd4cKb/ApjdlQFJ5BSJ9iEPacoaEjf2U1G
+6dtfxWAPlyzFggyBXWXHfBM6KGjVDfgFaoULwxLChmuXHnIdlxuMosNIaU7sjZl
eaBK0kRgqlpWZEqYDzswgXuDqMJf4nfwgt3vkybXx4cyZfK1f4UeumW3uwH9eRAj
d7VGIUbfrEL4nYPAjsOQ4sHNT1RXUNrAaBBWl2X+eFUS6eSZhD8lJA6ewIxSDMF+
Wii8dJsDXkq7qr6S4rF3fDs4KHAmtMkar1kZzEH/Fk0iqhnTQfcNzG8FkULpS+ao
swSyDFni0KGXh+zbAbR+emnS4V0hm8CffR+h415WjaRdbSRt33poqK9VrFsRKALo
vMlbGiuCM0mBGp6P9xnjpffC19nz/5QHsNyXIXQ3plZhKNAeAozrgoz33Lkaga/F
BHxOmidRrPz68YWb56fNthsiGvj9DB41WKlrUO5MfwKZjjXJhh7oyF2pPQGBCz7y
/ra8LbuoXEYP8+bSssy3iB5+cO8feQH+yq/3reWSUnYZxMC7SoeeY6DvNn5WjKxv
scfrwLM7FNhQVY0X7IuHMLU1g1pu8BVHu1o7f/S4BoLAGrwQWfeEiZhECV44Yxp9
0I3ELyJkofiKZaT3iUl7eggcP/9jlrlWq3rQ50nBqoU5PyPk0jKPQaENPr1D6CoB
FKsNuQJ1GPseFTXmz2DqeEgSFWZak0d1mE05sA7am7PeTsrONXCWER/skB2gRVKd
J0NWPmRaW6ptSLR1WnLSpiLk0tg2czVmgclUIBkbczP9ZkKqnccZsuGvwl2rECu0
1H3o3lKE7RGqhK0YqIWOFyMoFC+/kXpwCwXX9bXlQ7JYYnP6i/QOwPwQJNLQGBHJ
hOhBa1FkVCfT9PrPh30RoB8EUybloe+580gKIkhUfM3B7RFYk/FRQ52aQFEqnxCq
abmmhXrxM1qKbiLvD2+CdeR9cSHXDVic2MLTCWQWvT93COH1aXFi2tA8tYcZE0Od
7PsQ6usN4iWycxCu3jd6oznSZai6pW7L3Wx+MLw62guj9Jwdo7QqCDSBE57gTLu7
CX9KwmAqotx2FJA9tQc64Fjg64y6qgGFF5li/UN6bFL5He3WDyois+rc9gbiF+JI
kNjA1k0JOQuGEhBpo36XXzTtjhrP4P+Etcisj0rXFJm5l649ihF/4LrpeENDTe5/
9m8YZxww2WjLPEGjmiCwvQwqxC8lV1nvlAhvYqSG8RhgjnnzKr8QXGpeHO3QhjFu
IZcXGWI/1fx7rowUV5NCONgahNXNWiBugWro3ru5MQ5Qj/i3dV96p4edbO6+e65N
ZpV/1ZxP0SpbV1qT94MqES+8w0DY1t9y8+PzUWy+Jtk95WPWitPLftA1UEDcS5wG
FdBdw2jPgFDEPcdQQTDNlbQduFgir0KfggA6Mz+i6CtUhgJIv4xiVTbOOljcAhue
vtb30b3cj+rFpGkqU35Mxgcm6ukikfFToK79VTOfGNsR/FOQjRVHxqgIi10VS9Hw
/fncQeTTRu8pFNn2/ORbvv91gyxZmE1kjY851v03adTdFJpDtfNyDWNosu3Ro07h
476i1cHvTm/V3h6sfs+V39iIucnZIKq7u/J07ypFa2s+kPeIwBDGDjprb4SgslED
wajkjjOZvdRCsgqVriZaagIooQEdI+d80pcSBtVHVzLJyxS1uxARCJzhrYGLnJd4
yGfGRtA7RgD+fFYqYogcb2MdSt70vo1wyx/3OSmsmfD16GYhf9lyB3qq/Xhyan2p
Voa7e4ap+uSbTzO+ADKzsJ73F+IvEoDNvWrJr5nY6B9vutfqVabkC1XriI9XsfwA
E+7lD5pbNhkJznUTokCGed2mj6rdGiBEd8c11MJ71gGzY3BZ+8yo2UdYFDifY2/9
GXgILBZEM8UzUehbzLmzFbVKlI5K8lybftGCcnKvHHbwcYsYutJhItImVzsge/5G
Mm0M56WutlFVNY/qNx50i42fWowPbUInFKPjs5IZXHsxEbhsTLqwC3zBwhSDISL4
bOliGw349N45nFVFb+lUJQLVXlOmllrtlIu0ifg9Gu//Ry9tzrPMMSQgLZbYjwrC
xnNN9kFMQottkwU6TinSWYuS4RVvomxmysTEG3Pho4FEx4aODI4BhFHga75I/fhu
xHwvhKYSZ1V1giz1NmXBZmvYwj7crRxvRUkVyP2fXy10R9fk2d5Xgnhqspv23Z5s
YxCg2H9AqcT6BG3dwcB42+TK6uMlv8ShWshmj0wNeaYfuCodd2jxgVR6NrST09dV
mqwzFOx5Wu+0fBKY8H6IM0lczj0sHXOzcm5liF8G7ar25i16yxYqxIf31HDTNDAO
owxyPP2U8SjxxnC5SsPH6uoCkQiJAzYGSk92t6EcTuoyxLw0w025CODsBtXtyU0e
kQPI8U22aGhUptPM6YVWLK5nlb6ggFdhkvKMGQkSU5Pej3HMMaonwtJgS2mEmBrc
eNOPVrU7mSzytBXkZsb21PXHhQaw2EaaIa1S5GAoACz26aM+PF1+V5N3s466bLKk
xmrhZpwbyYx5WpUeLOcmLkib93hAJzXrYrtkD7ndqL6qWdEHrCJr3r5KPx9EYgc7
1LYx8fFkYYJPAu+yJ11u/soc1zIH55v/S3xdpkX16LAxjDFHgfKgSFNGVl4Mkom6
7SNSqJ8P3YJEqzF9p6A9OxzrptDNNxwZoeZHhqqkesnXAAjZzxRnVBOHLIWvi6di
Hv7JCZkCEGFlSxdww6j2/m9DfTcRzTSPGdrBYz705rb3pObBkY2fvHqqNmDbPBlQ
af5rzGm8jVfchK25P8TSE7jpoy1ZZkM2fH+vkDg/vtNaD5QWIdEBEY+Pbw6nCAN2
tcgpVYv1FkeNJ29OQcgPNX3u5yXllIVGA7CbNC/tJtWY4TOGtVAPTncmdr00PaZy
/NYzc/NuB2hb33QpxF71wIleAwNArHFYGStkdeqW9tPejAl6hw9Mt4Per+RnHGb0
3WTDVEgeRgxkd+CLn8t5fQZT/6vkFqXwGEFhaTaUTWa5icdqmuwFpvAN3ILs1ZmT
TxN51u0T6Y3knaweGPGJCsbcpnodTbEfWv5exL5GqrUfNbU+OYDYtCMJFQm0wp1i
eBsaZ/jRGoe/l3HkWC2u4uaYaV6xu62zrZAIQCLOeh+wF8V62QX6tv5MwFmUGvqu
j9s9BfKShdQ+hmGy4dZf25P8P085+e6ZZSg54IFhqajp5Xgz5lZzcQVWv0kyIL2a
CYh+8FUtO9m1diQRsOiMhyyH1WaczwiW5yvQ0+TQIXGbpotr/Lbfr+WxTV9hMKC3
QFdbJad3eEHOwfBNFdUKq76FZZjsxTZQjvokrGzlRAu/U9Fg2Ny1d2ls1baaYooN
eLd58F01gROdawk+eImpWWbHNALOZD4exogJvAJoUFXrIl63te31MTzyrQ5gofK/
FgY/G+ZfH+AV5ERVNkcYi1Pw5+7rnUHG8o3QkgQlpPe24IUoz29/lmepPpxDTHLy
0o1gbmU9+Wn3za02ygpQX6mA+9BSNbM3OcP2MzmYE6epbZ12L4YTbK1KOZN/ae5I
ES98BRbm67Ili+y/NyRjh0L9cLOJGoztwPRvGhYERTGQLP3uTHLJX9ZaqXYgWRjk
tWCWixE/WStWUx6nzs+3qzpQxCZeCJrlQDNgfVwHqu3G4rpbVeohb9zFamNXwk2R
GbLt2zg6Qt1pfBDQOI6Jkzrs4NAPHBVowdogUBcTXJ+Irbg6VvAP4WSRu12RrA22
YagvlcwoHWA2TjIYZo1PwkEhLQYXU6ss3sG/HXvsJIZuG+S9e1HCFMgqD0FPzuBz
GuInMmZODRSG/f6uZbDc933jumXBhYCvjwrMCIKUd2kIGTJ9HODZdcVVkOV8MnHC
DFpcvK4LaVFdd4490KosbxIcs3FDWlxgGFT0Z9Xkrt+oi965fI6jg9Gljh37eHTv
3PenK6c5dW41dtiuW2JY6exskmNRBsq7cnC8kvVuDVbjkmaD1Zc9RKgRJY5Vh4Zd
7DWmiWiwoWOw1n1GYCoaYqxpw0PxTt22rtEZo7AnzH8tKh0CmctCYoR/Sk3bKoph
Mk1laXlZg7MB6ItpQiU+9QzMbYTZJp+pJJ/ToUSH2hgT3UBAVd147NhNiLUL8bLA
Gek9++peiFfzy1hk40RUoRN9LyCy0rKT0zM6t1fOAsGHCTBkYJ8bbpHCffC7o8wL
z0e+hJWXhlgwv9+j2kvARNGD2O0BBXq5qxs2YX/KKzUkW7iM8ZXR1MqxRRA7+KfD
mNiH3IMgzcGQZWERuL+BZWSTtXAAZYg7eLf+kxweL6GxPg08FjFVLRBaZ3DRIQRw
RGN8WkK+gbSsHbru84yeZ0vHVjdKcOLp9ewJ/9WdPojFVzdhHyAsg9oa0FKITyKk
jZD+OJ8Jt86ZpOqu2KdYGUot4cIm1K+uSAljsTRta6XX3ZbiV2mdmdYj0deRPm1y
55VGO6DoqQC0ZIQnW6tT4or91yIjry09dgJsytC59VbzhvpBvBAnPyuWUJHmkUol
e0WlIJxG4KQcBBQ2XzFpfYoDBV2vYqsqlmoebMRkq2Yfxp96iYhWf+eeiziKZflJ
wrLs6W1gqWdATUvZwM6K44QanghH4e/igv1TiHdd6L8ih62L5Jtj/lqRhL03efw2
+keToUueLQ927LNDYvov9tMy2VCGKyuCy0/IVM5cRIlXBOE2FeBpzsVtmhgI2dS0
odlO3/XPWXzNfLeRRCWXZLLp0KwJTbPb02yq3xFeFXnAoToM1V87jKRoM6n7VNIl
5eP48ATwTe8Wg5LbgUMzsDWoZPSxVfq6c3rTiYXmK83rHF0TS5wq1SxpfrnGlJHn
qXiq7a1X9cdr9KPdeN33gOmAFFWoGrSI2ffRuKd2tSdDizUyX8ydBLrhjhuiebE+
w/s32SBoCfMB2makBC9EeNvTBy0iXFgeVct6Oo80zFiVPnq/ZP3UgujGqpG6ySh/
kOzWAyKnaMivRIxjTfB+mxXQG7dumTxjpv/ad9i3dOPL92OnS+LA94E0cKHKJNdM
gm2uWeC40dKCtCU56QJaRkUU3BmLmJMwq91QimzCoBD2PunWGDhRs3PVAH9UAg8E
Gg+wUl1zueQ5JwehCnSIdPRW4VYajzxd+RQthAYObobw26pj8fkehj0DM36OcnG7
ExNnZI6g3gLXvh16d/BUubOZUcNRXC2yhymA7Lc04030T5utWfJ3a/rxg9jilYc5
wuirrfkV7ymZRz+nuFesJQP+WW3BvNLjobUEHpambUwfvhZ72MYQq4/nE6PZtyTq
dTK+iZX9wLQWEBtxleewFLk/x9/Q8DVN9ikt/8I5ByPuNpC3dqSRYZ7cFZ4FMhgd
tS81cuC1adbrLpOo5tteOpFCadbrfja5B6zTc71Du0u3Wu6fMLgnJxZuv5I/q2w9
TRbu+c9zRZlgo5IU/SdeQaQddv2oBu7lpNDHrPY/GmwbH3vpx9GpysHIhzLUH9m7
Q7YXIdDwgwc+LePeqjFw8lAWXHxL0jBLFGgGV3Ak2Im4IpBzKXtAvwNAcCpqixoE
GxXk/W8zKDznwfEMusGvzs3YUSSkdwg8AvbnV27fh6nqKpuqr2Pbom7GMWe6X2Vy
RXPpp8ww5bwKCSCxllmXHjeACeXgWoq8X2xrrNuQBl03LacA1Czdw4CxM3BztQim
z0qcvy5gZIFSkDYmnknByhJQ3jn63tpf/xo26P/2Z/CtlGrCIHWPX7JKxKNRu9oR
L3sTcuIjQdvIPOdiV3oWaPMjJqDRFTWe+Lt9M3L6hP5Al6m2SneIZpMvJduKeI+/
Few/JfdcFI2RsaTz4/BGzVrUclnhGE9gtCxjIfQsR0uAMgmSwuQyhouV1KQVwgP/
0JUR8RC68OkmUBrssKrgz8gfhri5MefrLB1B8JhiWutnZnnOqbRjifJMbhnzp3Kd
Y64BGG4KdKA/7zQxI4OB4LQqipHikYgJ0Dw9UhkMoS+9X3rF52H/baGbhf5WDJwV
oo2Vrn4o+3HaA52SuD5RCZprGcdebvXbK/iCDXOFy14CrYPZn4wIuJHGfh61eOon
OTPTsMJNP8OrgS34giZfvqbvQ+ettCG1l6+XRTKoPJsNhi4imVrKrfTPZ6AwVajA
0AxQ5+hcF99uTKAv00oBZX5o466V4jla50yEdhhMtt/clbi/VhU36aYykT2tR2KU
izxIkxgMeck2jJutJ1U2tmy9Y+rxlleHstGNYdB9IGbShWf30kv8fcflgWKfFNg7
iyIQkYKW4gUsPMwXEytcc/oIgLgBN4AqkRXn/HEyzv3HoLMddGq5FX+1RHDZb1yF
w7Cr97IvaAapeRoTKiBXqzmdWq0vDdh6jpmybHGIDbK3jTUTNhZEN/ACRaw2T6WU
qzmZsnSL4IcT7dNwMnib/E9SXVUyxWf/nRDTGBEghJGLBsoz4IuiYoAOzvoE6zCT
VpczEk6I53zQn/IT37hnRzRV/Hn9gh7VpDQK3+DjofJgkMcwYqFsIViYlTsj3EiO
bu3JKJoZtBRX785tpqJg7xQZ4uUtKC7TEuN8KfKlHdUlA9GjhBwI7tBH8k/GtedJ
5zEzuAlAvS/7EP5UaWkr+nNngjL6MApJhnJz0vyWDzfIebBRlsPh1C54mvAAWgL7
inRydwnvNVWaTO9uBeYweE871hHf1hDZsXu6zk447f5YlHN6TcAs41vvrxspLd1W
SpIZd1ZylUXhEOuId+52FR3j5PUrcvzJs1z+81w9RJzmlRjf20ySGYTT/HOUeICl
7FhF9aE7GcnbqQg/htZeceX+vk0QpFE5nBs/SpwuSsiKiGAXbR98LIVkP4kUW6kz
n2/BDyQnSTs5iFH0ax0PRlfSSSS/uKt0kmpTlpFvuJ/crC6Wqs+Jc0n3Lg9aJ9cz
7tVYlsuX5m+bXRAi3Yra09BwkQssqWiETpxwlrNXCqmYyb15sHbzTN4F43+EdHMz
x63zLTOB13Q9icjLKnqaUjTXBtcNQfMQB4o/+ucGnVrDBlg7fZsQpnQs2Jddhbzx
D7rtnk/QYgzCEJPjyL7hn/OKYBdqYxhEzJxUj0gPCIioBlnfyt1EhE9N0aTMXoIN
ZQRsciUDJN75Ti0eRn1rm86yxth4iu/0qdT/Zd0uGpkv2ogJ1k5dk8+k04fuQGsl
bFU12H3NswNYRx/RSUyMKUfadOqdFp08pI0SnB1lZvzBgd1H2x2VW6sNVP+nDXba
gbEgolaAxPfUo6HeFsP+V2/ugqLkFi7aMp/+SC096dTNgz5Lir2wciw54Nu9xbmM
46x7lIXFam8XiMCcQbH4GtZh2O9Jgs33babcjEPVos+vFGbOyHUF2YZxKuboCxbz
j644SawlLvwxvCElSQeLu51AREtYdXpt+gWl7c1LjbFGxHMVLT7qBTP6RgY5q5rS
ahW9zo1X6y4XOHNkGYcdP7dUbTfVVo3UFk8BtVckTATVizjWmDQmn5tj2pdWCsLg
SiltVGxDuQ5A7uqmypjz4vZpwnJD+wUeM0QgVpoYvgVjY+V8FCfTSRWRzkIEqwfa
VJbL15dKPLXaxjEWxZGtIed2y15GmUNAbD8ATDk6pNxheOkcl9VJFSA938EtbnGm
EJEj5ivq5NqPTCbb3G4TvRzd3beIj64yhUTF0PcC/6KLLoSDbaw6/jkjlIo20uDG
+rKfJxQVQ3AEoy23CPo52nvppU6zyAZ17kSSqoMQ6/UYoI0S70gGH4Bwqt+ggbOw
RGKgag4lPhFriFrXcGqJ5hR3G/hI7h0TiGKSr6W2Vw1oX9RDn0pyajCeE1XsI98I
V3miaRv8dd4ulZpahwoclYYpsgSCQufNAZuM/js2KBjpTS1iJ903I60GFweWIX8+
P2TpkqV5LjkOA6A4MO9YkhV2oCfe5fHMd0gTmEnpLYUEHyrIDPZKnJLJyj1YgaUs
xH2HRJo1sj1NaHQ5BY+oHRHFg5I9qI+4dtFZ3hR3O6CIgXhgd075+IE7PG9AX8VO
otIMUOWqAV+FartfYEk3caP1XDcIAWvsdrEXwct5f4JS+o6v2m3/wtPwYvKIYszt
xhf3cI5EZlOwMRsV+Jg07+8E8Yio0iWrSiGM7Qxw68nhXd7sgZsKWEKIWPQe1Bw5
d6425L2q9PUu4Q+hxdpEPc1YZ7xmj4gxgC2bnFuAybMF0WscRe0LBUoSOvB3giew
5m3rIlSSJcaj8X+Q8GCTrKcgmPIvKPtXkEYN9LNWkLym0XuPvDJRhAcSDelf0bNz
c6JAzzXUKEWQXm9ca6XJi33kGIn4QbOaVTNocTPOPkQWop3WCPyCSdD4KVkNtNAb
9i+jEnBy9UhAlIlFcGvARhC1OyYBL8VDW5ZCkv+cPFR2f2UTg3h93X+Y66j5nYV3
xhpu9w/QI4ybWfXkbyf2cuhCTNyrl48JiTWsrseELz5lQNJ2tRTC9ubhaKwTz+Mv
C/yADQPVQJwEegVa90U8eqKHD3z1Y/IpnmT0SdiQ7/C6+x6fbmNCOc4uIqcNtVLE
IeuVNTkuj2movVVnl9kOWpjEzYuq0pRjU1PlsVfO0xoD3Bhi7Lb/bHtxEjabjExk
Hqdnc99QD6v+B0OiAcI8Ke5TgJQyfQZCYkqvRARR5zzABmx90nXF3ZzZmlOF3UC0
gXvqYEpKI7gUy26taVLkqprUlv2eKozW1UKKZ4mGm6Wdim7LU40EtVqSYCm6BBqt
DDyGtoiYExPe1VAnlp3rqOLpsJC0lPd8bliOrDoe55rYkt2HU+J5QxoCFFYZfGQe
9+QRW/aSA8wVMu1GcmSW7rrcxfVw2HhQqXZiJNZTFtNpjeXZj86kQw+1Aq2gglXT
ao05Jng+y+/8RGFJR80Mdn7jGyGLrw4ew9wX00YYg63QB/UyeXnmnZbFob7aDbWj
Fpo220wIiLrN732cCfagZoYQ4f+P3GgoVdoktG3bd8HI5mODoNSIq1a0oTkNk1Aa
IWTVCL9mobnyi49ASXHoaRHH5H5wSMOYspOaHSFhd6C3wqxqwAic4Axl2aEURWos
w5o4TduNR6CU+vyZmALo5eBNdiuGkffpOlBStfv0mxYyEJ6O8yHuW/hGsOrrUVih
ZcPsEKc6KsdBLG60mY9tmAVVnzv5LMSCyg/a4c7VeML3K/J/pVFZ4pfHc1qIJz6C
w0x9hGxwL6DtmPIxCz/UqeCEAoekSWiAtg/KADQedW4xw80Mc62CZ1Uk+PkNXvm/
HonzeONQOHfRccIgccUb2NVsbbLkG6BtJl9Bw8/153KlTLlr8RIubsQFBWw1GuX4
fvgeMcnaXUP0q1oQuCop8ygjA6V9ufS95UDpSI7DFxL9avTSwVi4u2yzZRJAds9V
gUO2ClPkHJau+WASdmQFlQYlCWFjcMHv/+6vqQq3ocMPTltB4cgn0G5LDhyRuL/c
9yqV1q5KDRwkmPVI1X54oeppU8Tl75TtjHeverKByKe0MZiOwV/8vVnA/2De7BYb
7ep67zctT4SyU2OOm5mgQS7GgPiFXZ1IhpvdYlHDGH3nI9FC1+mTv6RibA7pn+bQ
j41sfyqnXA/zdcWtzJC+0kXGuzCJ7GxzQCntFK4OmOuL8bE5CGmPIw0suIq5NzER
piw9/bsv4dTOGSW+Z8NzWs9XLhc3ceyMMnjnCkpp8GDf3A6vr0gyT8ViOZ/v8ZGm
d24f59cKdx8qxd9CvlzmXX+evlT0EppG5AYiPUWjIZHRlEePycP+jVVGbfmAdAhW
dUEU8nq+lQ46VRSn6V9ipRWq79O9LO/D0BPT7pAs7HH2STfz9XkX2U5kyo1RVnhk
bouwjNBFjQ0cMtbB5+3apGH3T+DLmtwHGC4vnsVhs8Od9MCL7jCE88j9wAIzXRTK
kcOEcw/QBgCglVFhS8aizUPz9Xv5VkLeLljVLMTuY2yc3nGD+6y8Uohn5LRoIWW3
yS5copovfHB7jAu2laAgiywwTHP/Y1bN2W4o9A0OgNCJJ3gwM3KaQ7zsqV+VwLQy
UUXmcCfaX6gQMTE8ipsX0uLO8OY03PRPnQXEsrcW8mtwjwDdjk7Ns9tPhmtpEDI8
BUX9ILKKh0mOKikEwFznbmzJmdp27GiIwBd0UG39bOXl9OsicHsz539jMpHkuCr4
UJH+4TjrrIQali/nEs+30Pq8g4L4Eypuy8I9mFiGxd1+EcoEsYDTNs/be8djXqOn
/Dded6l806aabQQ4jCabwadUoVq8/w5oO/AT+l3rMcn1XkvtE+0z5rMfdSjsraoT
3Shv2Xy7mrybI6u++a055BaPBGgk8EmyEE72eCMFXkLbok0RgNq5av+ZZEd6UfKE
xGFtrB1qL8cvj+Q7FQal5fmvOb3y9ijfVzP6rv7SmhbfVq0iyvwMf28xhW3pIDJG
H6OtRspiZ8TEubrr2wVXH2gVSQ321hF0orLXIRDdmnL2p8eQpD+YVpwFQAEh1s29
suDcvVkSZ+Wut/CF7yVpfYshCFxCqM5Ji3CEbJw4C0lCIt05Z2AZG7Wt+u70v3Lm
ApYTR+d1G2TjDwleym7wW9eu1Tu07g0mODvaqz408XVpl4Gv2v7SDE5RkrNkHH3d
SFvqQd7nQHA7X5VPbLVjD8vHwuKw4W2XpQb90lckrVJ/G/RYTv2T7WGnJ/X6kWGg
FywGO/1I8w7ltk2ZybnFeVAASoTJ0zoguP5ms3mVVYLsRrY3JQv6OGqhtlNbmYHI
86yRl91gPMBviex5eDUe4/LODBSSm9m7DpSaBRAiSvcLqsnQicaeLmpFdxPb6yNd
NvFFegDS36PA9n06zipD6ffgXYj9A5LjG4WJuji1TV415Xi6HIrvtJp59oOG44G/
hxD6M1PJmddhnR0NChnfGrjIHmyNjUFJt8pSYsJc103U3GCFpKNV2WGY/GijIcD9
+lMmYEWJQ68MStlqN1Pc6CZvsOaCXP76TPtbKx6AQGA8drcxTBmxbxIGTfo2ay8o
BTCr5nWloWZ9sr7RfWMKMl+J2KMhxv6nALgzKbyZ3tUrj60bUQizShybdoY27ZaQ
uI3bJwiyDn5yGDugk63leZpMvOd9/7Ta/llIxWy8F/7pTri1afe3ODnvB32IdCf7
78GKA8ScmVkeRo5k/u3rfB4ZpkbMNH7Onk44TeTRWaK6G0WOrbW5A1l8xexgZKF1
lNDwSEM7htpcfOPjwX88QxejgpugPE9cORDCvz0tUgtKsknuXqrDcHcxgMNXUG6E
6cjMiQ3uDMdWYh0OlOtVPy2klRTMsHImlIUn1aztC79ujnfoK8otfpauwa2c5nZU
ba/6Kca1RdeBLbGPsb9oNo5XeR2xLEBUAFJbkUkuckeOnm9Aurrw6CHlfqy1tAVs
YG69qs/SdPC8TNydDNH1GVhr8z3pC9SN/iTp4rXboJHo+hyR2bKguafSx2/Vfvi5
c89W9JZ5Ww/kHZCGV2vKVSJc3zEq3yrX5uTEdXrvuOrYem1tI2qOimV5dSh669Ts
ApQ7MBkRj8vceBbe+kHDehVMk8fnnwKXTEpjbvFiSWrrY/u5CW8mqHv1Z/+JLkfy
RHOBT0bvW0LzP8+2t22PcGEYfWdNIVAirbq8e30WWDhYyR2qRzT0QuoJ0vcyF6gg
Mcp+E0L/qPyXR3RPZrHz+5Nuqu8ymh9kC6gZ2WxkBQMlQ6pMZVtKUhGmVwpD+O/W
rFVJJ2PRKarAbqCmrJe5DalONZnK9o6V6xKWlsMf/yvAPCzk6wW+J2NDYNlAGt4q
b8Pgt2/7fca4kQF7F39MghODo0kPCDAlZ7szqS9ZnmVK9Mzds7PeQDhaoAhTeAyI
je0VtSEXMm5DR+4g8KN5jLhLoq/YeB3O2fUHgQi/i3q+uMUb0JJH0xN0MUbEYtZo
eZbfVsb7OfF+ZGpHRrd/mkBoWqbNUpemFDSAypumLC3zmL76mKGJAft1f9JZ0B0e
iXtsNmnnl7SShYMHwsUQcQhSmkb5Q6T/CxZrCOx7ubW5gBtA8Mzgv3a76Ou0LUp7
webRpRC/cvM6m8NY1F5ep6tDrsvF/UPoTSsbmiufGK5fjMOcRMduhg7N1zvGTunK
MJ0SNbGY88ORMYo+6MjlKL5/rUxADDg0fyI6U1sfTzV10TzDPP3D2nC7LW+cBQbf
pyRd81VtQjZf8+5ag/fr/cxqixQDXWQG9IJPZI3rl9y/duCBoUoGYGN27mcofivN
K+OJt+ZTH6DxY4/5gAm/JOO8Awm3kDsMGnhh453vShNrx7YEW1n+mT2KD/b8p524
pbFsDWXB9LL18Tbo0zv9l9Totr1UZt6r2cnnvIw+kf2ARrHrdQBvk7bFgWR/QqGn
J7/ZQGsOVDSXXwokg5v3J+vxcDaZ3oJ/7ySiPgnps9omgnlqVQTrdZHqD/PWF8Li
s968XkoC0RTjPv+nW5nFg0HxkBVxHE/bTY4behEJ+TqF2qtBETebv88DacK7/Dqu
ql5ci/9x9OwQonTOYZb1JAjOy5lKaPJlwjNN1FtxjLNvZ8zB2luwhdYvvRo9+Vqy
o45p9ErvZa+m2HVJBiCqeO2/B1LsmIFfCLVTUeVwwPq9Bhss/Lr6hD1BUGYtgUmp
xhEiwQ9S1lzaxGnYiRgTU12n5EsB4IHlFOEJ3z2LSwndKJcl4xxBVeYCBqN7KPqE
Ldf22oboomtLv/eNm2X475gP2Npiowqr4fBahvKzCgIyLLa3wK2ESLmipNK61+N0
Yp+u446ozc9eG2WwAqZ5f1Y+qt/nqI8MpbZ9ndCQwvmSFrN2gr4Pw7kb+HiErIHi
JgRat9lUAJwpLBlDZ9vG6tGH+G8Vjfp3njq+6liaKCtSFd92bVpgN2K806tG+63Z
pfvrnu3/hzvV722XgTvNmHZen389sHFjj4/OOCOWSdAu6ZqQLSA7gY1zCxIq+dSv
nvRsFjgrS+W+cJAR4FP8HwUlAzMz21VWm9hk+7d/OWwwc+S11Eg4bzfjXnTXnrA9
EzLiRrgIubUhmm1IO2eb5Qem0QP8NyPGsZWq+RxkpYsfP/gf4ogD2lsKX19JFEE0
Hh29loK+dVYnj795uk2aFieALCKPfXIiH0MJrbo1BTBanvdnNK0jW2SQ1PNStVFt
TMAFZFkZDNR2uEwKyKWdK1ptfQafbihpx+ee9idTdod/72seJ8QVvKXvtSldXpke
a6C/WOl8FBtC7BtkQgrDl35740rylyACb5tfFbnzJnAwY4K4UYM428RdmJpnszls
hU53WprrCnCGL/lm95DKyCBKzvsJ0vMxwoOmhwIZ5NUH0WiRuGqnzvOpwaFKmK4u
uAVAsRieKbu0RaXwY/rW3t/Ea1WNFCU1JDgyrFutATb9PzHdqFrA7Lgu9Kz3itCi
ROszik7jnH1qb61+w79woTGEk4zFUWEm36BmS37wKxJsO/kh2efbZs87A0qxvGcH
5CV57m+R3B6SIr/+8iXheRwvf8rlYGh6PwSxQbp8zuMkRD0221hJge+44S+avw9M
cR7QRmTs/W4J17RsldIklyk6mNLxB7xUavzwfeKo8CGPUpDzbQgZ/CjYdCzMIXaL
JtsEk7vz6eV/aA8qArayQH+5az3V8NIIvrKod+d4rXZL/0mnd4bQlGwhNOmlTUlb
j6MRDnexg6n1fzcyuRaAxste9brLRVt6rTHBfQt0urxXjHsTvW+mhnYxQyxWROjj
Y4ojgxMH34Eb+mdfBHY/Y5hrIvLdE1WGovk3lhfLUnu5KJbSqA7PEx/ayyl5BSVi
J6FIM9umAVINrF8Hj2Hq67+lwnrkzjWhufIbC+Htcml8XFeKeIdO5hFZ4X5tdCTp
01aSes6jR6+B8iRN8JOaco5oGkxYGgB4b8NQNVwj/5gyqjZDQuSnqLkQvd2qJrY4
8vSzS+FHDYgmqiTxDrRN1YYYFIZg5KH6wsVKGMty4uFc2tN861yZMUg6s/7aAhwl
i8ArS6+E/HszXMKu70LZg6Fk2MLLXGcqw0jq7xnOJvgoX6eFPT+cDjWRLkDPOE5x
iSd/UlhyUoslD9eAwbyLHvx+9OoDskG3T6XFePXxTBO0eT24qdtv0ZwDlu5alsLg
Hf0LRmSKeRktc8/szm0xnTIs5+96sIzv8xFZL1Cs+Pj1YyyAk9vjZQ3oKt2MAEk0
wA4orhWkobO0Z9KjrVKJP8KCwyYoFqWv58XwUpiXeRU7WavJ/Rc6aj6jBSHUOUat
eT1KpsvhIZkoIiCz3K8pR001NnUT3ZwhBnr17GtPbwoGvsGKjBnNwKN0skhdpNCu
dVOx1iZ6aTjl8ujColtg9hDGDWt4RRpZyQTmSs+wD2vmdhk1HYyQuKd2P5qNRngn
Yn2Vf7t/MUIdIlWjSlIAiWG25wTMNr4OfuRmgO4JXlNur9eWuobmscL0zXNdvmE2
p5d1gpyluumlMiW75dTGr6xZi0M5KrEhpeeH4gSRw7RwokY3ZykDRDH/VhW29/jZ
IRLyaQoX4mzhOLmZsa8OmD/acgmlltSVxZxrteXSG3sgFCsFf/+W0qxPlYHPZe6x
9JHZR5vTvaZTq4MQdW7hDNFblkAZMN/pU10Q1Iibk05dyyCkoFSvnx0H3Z4LEzrV
Z8F/nkosc/7VaK62D21+tGJFv035fiXcLTR+9N9PB44FKvdcGYO3FyGLGjtiZctD
KSGgOtR7dV6Glyb782eoT9YlJ6oieWMd/kp+cBOB2VNb2A/MREPSRCOCfkM+EZdr
SghbNdr8d20r+4PK1EXP162nmy1dlbSPddxReADhdY28RbhnoJonRAFZzUCbA8wr
PfYLxSqZwzJ/55iQnKi/rIfQ2FJ9I74iUI28DtBvHwa2D0YkCOm1kRyHXJiYlFDn
oCFa1JECqt3rg4dGIhFPa9Jspvzb/PHt+KmXFM3NInE0DU202R/IFNP6QMffMZLy
7XD+lMtC9fo+euiFlRbdW8InHFDYQTL3+wE/mhziwWRaq4N+S2kvGUl/w2jhJE24
qUqwA+cREUjdeYJ0/S04s6655RrX6RHiHyORJC/TsDsUY0aLZ08f7XBkEWFy+YJ6
JQXEsGfvQZTCJPaSu25TD8MBM1Yt6DBH5ZO9DvtUIvg3VLSCU96VvaW/x2+fsEi/
xotFTV71fPrb2e9et1TxaZK1ZJr603SgGDklEgJp2uF7ESkG5BUtjW263FMlzToe
aCZsfTVIIROiF9yKKQpwCUe9PPxUbptuC1w748jWyFqh94pyjdSs4P/M9zg8qxUE
TeDi7q/aV1DoipRIiWBt8XC8g5dIjAYfkW/asGU9BV14c8O93ecCoSnozSgxWbkm
1cEZv3T1aEkpqq28iKXyNaBJb2vZQI67ZFO8itFRjWv8iiuOclqTIHWgL+CJsEzF
LpTys6CiBOOaZdR9mVwpKBK/ehYrTLbUMjGoBnzC1s40UrTKOHW6XtNHEqP3CdGI
riblj9BJNKu/0LA4bOc+kvu/KA3D43ujnSVWwB+LlLK7LbdCEVKo7Ksb6o7n9KPZ
FE/K85f8cNZln0KfXhh3WnAYjJsmgd0y9gZgQt929bHAJsjPcnlsrk4rwVWkTJbO
v7Tai0wisYrcYf1YvrHZii6pD3rx/0jOQRKRSYCCapnXT+QgWXEeBRdLcybZD2ar
r6B9nCcRndgQU+wlOFgy7pLHfig/T4dwlDIL3fgRsiJbC9Hm73Vuws0S7dbAvfp0
2V0qjpJATI/7QfiG8a3zJi+k+cbnqFKGVjnmo+Hgda0offYC5R60OJiWlmB3KxM/
WJgWyzLR7xFYKjp3eOQfNk11MDWOwBspPQuiMeIEOvzDuJt+U6BIsQR/D8jt43S7
PKcIZcLj3y8B6V8o5+USf4MsMvs3X1mTs13yJhcaSN66UCImRiC81u4ndVC008mU
9MzbZlWmQbgdXHWT5Y4C9ma8cFn27SCiwVItMGWM/9LcK3YzQXFG0sl+0zHadSa/
xraBTpJMheBNYb5MUOSrcNp+deFrOPgqN9VQDXrdACaat1gR1FBUN/K3sAN1LbuJ
r5hjWba/XnebvmbbZ1qN5aTHzBkapB3BD6X2/XL4AijcTYGBymX4xtN65jnv52Xp
sVwgMvf9fXmNAp/Jl3S0b/NL1ue+zCQIcA37cf3fOYy8Oa4SU3S7EQpUd/G0Zw70
0aZ4OdgUmCc+WJjHrH9trK3G9b8KhhEDYOSw9wqppCx9+t+FzPu8lX5T9+HgqdSw
v+stBSjNkYWL7Fif4BbhLpZPMgAAdXtqNskBfmSjU6gMk2LiDS7E06uR+4PKJeg8
yykm+k+wqEv17ML0ozrbO7bySQl+DyT17AOlaSWSfdVrtw7LNBKn/cV0WXU/uKI/
4YZAWfXR+yyONlUFh1ea85pXpO/+n8s9sXVj5tc1DoQumzX/sQH66PIf9ASFJE4F
eYRhiMtgbjz89NvzYuHmVxU+9YZU4m1sjmqZFBprndKgcmv/Aa+zuT/4FAW2rIeq
GL1BjEa5MK8pT/I5iPU9r9GjgIS0DKd8vnMl684GwdRDEYMkrexNIlLgOLqEijKm
tS4/w8hr2k/ALsZqX7CvXMRoacoGqZw0SgKjRuK3D9PiwMYgcJuEB5B+1cr4J2NM
vSJcIK41yuKLqzArTGVXoq37vZMOgE1Ns98FvZ6hsAA/cfkv25AvaS0JAKe1oS+r
UlVHM3u+kLcocwwzPpS+oU7+7GXWN4rWz55rkLu5M1HrgHsv0I5PoxnW1FF/q7Hf
MuCRU294ASToKjwMtYPgCXa3tBD8ahYADU9RxFxhEBKiw//u/zX8/V65WMnUC+0i
CRDhU6h4LNY59Li88Ry4bcCR7Zo4oFacdsrCyr0iB8DQZaAkqFmAbpLSlz0O+4/c
DsP1kgYeQTsqt4Ckho80TcQRjdriSVUBkof4nbwmL4gajeHztGIUKPnV2+M27X93
UQ8pTVAxYhepl5AFQ5dEZWbIuSgO0MWnEt9CuFmnPWoZ4lZS/KbMC4o2cwI0NEdD
Xzoz0UYu9bZkGv5skJbihUNo4Y7irvVIMpvwmU58OLLBeTtMH2x7KeVtVQJVzSrR
RqysCHrZDYQtF/VqPzTKnoLbihcIcP3+Rh9bknwTPj7TAXn8VF7QeZmXxZ7gfnZm
esQTYSVRH2ArUg4rHmWScGBMS4IjOLQT/uqc4QOVZDIMmV6Nqt9+/lUZo8/fXr9z
yIUc9F99tA/JbpRaOzD6mAUK4wge+OIrVE6kE+KgY5JXXW/QHX996YTUvnBlEUME
71IBxmdDw/OiR6c/HAupl422cIYF70zg5Z3CSOp4/+tcABvc6LxLeNue79hq3oI4
s9dp8yEDoKMfA9Op0i1Kults/4mwuhG3oksb0PU4P9eQOrVzer4L0qX6iwaPKT6U
BLGk3jsdYma/ofiEhDcb7etZVvPQccezpnAI0fhvj4DbS/nRKUZrQwXoydSJsZO8
6+PKBMlnyYE32XU0/QW64uCM4zVasXAeDQ/WwqwOeUsOtJ/rD3gD36tcwWismE82
1wzuitsSTd98J+lEuKGmVCa59JmlV2izeUPSCmi2JnolU17o0PldpdkEB4fi1TRL
l0qBIGaQ0waHyjtIYldxZs3mSFW6NMg1FlHr5fOH2w8bSrgkQAWaya5coZ3kg71E
hfkQe6wsfMw/IPiYytcv8AvwFAqpVv4Yx4S0OKnyi5AdQ4wMzg011fC6Byx4PRLW
NTynGD0yuftOol1U7c8A6e+a36WaJdgLjmgscWH0x3aDYA9EI+w7L1/xdSssR1Op
Ap16dfXYAc2+TJ0QPtrZs1wmWX+EefzNWvUmq/adUhcbumfpKjxBNet3oEXrO6FR
Ixq75eLyJmr249/PF9mgF1OecnFKxTscvHlqKWBZQTSmWW3dj2Gmv00iwKm89mt0
1IyjyZKCguSBAiukFCn85rVQml+Z7nnteNCoo6mCWAzOq2w1QGTctllxTP8si533
5AdyemG+qJBOUUuiyFFTV1uMWNSzrYpcX8BsKh4RW+tCCwnI3jq2M0A3h04mcEc9
6stSc78JgVFntQX02evl6kphsIggDo6gCuWb9t6uxm2kIoOJg6AroaVj+GzanBSE
A2XzRWAdoXyceBAzNTOBL9Z2tvF/THtuS8TJEyFkgPLSkZKL0nzJGDpocsJneLcR
LGxiH7vL0Grwve8QYySxwYjsDj8fxUOIxf+lxLRIn18zUlBNt5QaSOn/VmqLLts1
HKGweeolEnyU7aI58w7qbAik9Ac9ndEQm+JlZVPMnsSh4YP6S1HVVQFRiW0WFvVr
3abT8C4kABP5dZJGgMMQ/pqhWHi9tgwtol633cWrngFd2Gj/aPb/ac/lyDdHjvtS
zJOgNBlr6D9lSMKpcvetyeVzZEck8fAGk3sbPTxQ/XdJfUeNiR/ruQDWY3gdDzvK
P8O6XUeev1watGX1PlDSaDI2SF1hR5R9SdQOEbrXN3AsZoPdCq+Cy8rqE4qxmSh+
Mj0OnCM0ca6D7lGqamJ1TfkGHOdczdKmj9Bv7L1PFR5/kCXB7mc361/4M1lJui9t
G/QFTiPW6CkihW1WgL4wICJ9X4uCP7xpQfWLUH17v6DW0tn3hBwIZldPFwcn+Haz
TCAKAYL3cjYSGgR0zdB2Duy74a9kFkyiNdzitXl6F1GT3PQvoOArJeExBicR9VNO
xwVWltkE9X+BGqfkLTC2ZDSzC6+9G8WduG897y1nQlA4Cfx0FRpfGONBLFRhc1wj
xpy/r2ZLQp20kC2xoJgX98LqTtFP98ujES6/M51qzpBlvCWzKm9cP98rR8hGqns/
WSjzyfg3tI6DYxwFWvd/Ro6hSvy6HwBK3HSKbQEe89HvrUb6k/VZAs34f5JKWhEx
D19EnWpkY7Mj9GKgCYQNb7GuCH7qOovo29zq5E8YKRFgvDH8L9McULkey488HvbS
fhoQu03PLMbAVnnio0LybWKC8i6D4WoHwpYzbj7VUQK/A6fIuitQNPg/eyz5p3eC
DHIBYklzkfyeS46hPs7Tz6bplHLQM6s63z9zGa8c/uPXV9SKgrI1IK6Z/WMMwitn
sB4JUm3qEpRjJRN/Xds2LdoDMvlcQza4pDPj/dNux3DXmEajAPDAcbY6kSr1WY96
4rvmdiYKeuUwAJAYVZ6Ukx6yif+Wh4xRqJ0oIDz0+FXc0Ng2Hl5UJTK2lS+uZ3zQ
ssbAOk64xMenfAr4LRgEfQt8u3R4SbLbgCwIGgl4u6U+xr6FLCSxej4mXw8MAwCJ
p0wSU4MplGXa6lzOrfAnM5ihKEkbqlsaExD7cgm+graHu4QQ7fuNgRGtSQKzddEV
Iqcb2Y/DdvAnA5h3/TWanGSberohMpUTq8wUg+VqH/J6Lf41Sbyhc4VuY4KnO+gL
gqHIxvxeknCIMDL08YszRYR7Kku1lh9AovbfYUTunhBRspi9+J6PdvpU5IM7s3Eu
0ZQWT8GGJ14BMctWNbVtLBoivQy4Rp0bw7l7EievgX8vDf8D6vCvEeT/06GG56NR
0r0nWdLmcvac72EjXkbcgQnM2tDmLgkLndqJV8QnDAya35HYvJuGrYy+6gY+Xx7s
rSIWg5RgDXSy0Swcfpcggqy+u1VV7yfsIaigGSL15GxwyDOL76l0KxFZcd2bCdwj
SX6uie/RPwTn6R+I4UvoCB+QMFVjwyndaSs1ObNkB5+3TEf2ty/QzP+7OaEZjmi4
uYiVGiocPeHjqU04Ngz3GNFJ0pZaj2SurpEgo/ZQRF/SkV3uOX9QWTeOeFJp/AbW
j90GAYod4LR3ci8fRgBQBs9RdB8m/gFReo0gwlYdE1Z0Q001geZ0IEgJy7LWSd97
QV7kCLpOxyklgik/IKxe87ExUUDpEh3Oj33C7JYTOwi5pJt7R3011vq81G0Th0jl
9gIylzVtQ1Pr8R/70E3yA7+OgeJVWRowRCmukMK7/7MXM9lc8Ni3Hh1YK60OFvgm
neXt7Qtj39ayCkyDh7JzYRWSf6K1EMaulPbO63LPVhjIY9oGAiVcpBtPPsHrgRxk
OLkcD18U54ziNPq6iMU8mgsRvOxaG8284ETttx/4QiiQ0uLA83lyEIc/YBYX3Sb7
kIjXQ+vuMsgYpKmslQars79MOFqEGC4parVK4hZuSEHBH5B3fQn2s8NXErDbulB3
Eu3ggcIr7txDb9jmZGe8DUcmDaQNGIpl4zmObdgjuNk2qN0/OtdEnE91O5M2++Ah
yvx/SbgpKswHdQL1ZFhTTHW5hkIYyBwSGzH8ZdlrEVYtkRGzYuY7hZ5Djoady2WN
ggJnX6LLCTCRw01hchp+NRXFwkqQujvFCQgWDX+0CST3f/VIeF9C/jUlzAfFFXub
KA1TIlW4ELwGSAOuSnQupZobDRMs2eU9GldCWd2FWdEcY5OKe3Zp0PB757gt3HeZ
dCHLnF1Oa77XZhHAMJaX+FNyj8/NJ5MU86YteGF4QAbgu5SihUiaQj/oHgGtir8A
CKlFADQ2RL9gltdO0gGA3Cemvd4FH88Ty3rA4useY1i65WkDpnrT/L6Qy5SAmFzR
gx+6SPTqVjg4eFluvX62H/kB4+OGy/Es1NO2gxNMu3RuGA/W3OdhlpJkUp0Gg6+M
YR7v/373cVeGoB1X76Uff/H+dWXdgSTdMOOKGD96Ri4aPqzF0XOEm4EtxP5enuuc
Uf4WwFtqNJPq05rHv9Y/fUc1m+dnzuPaG9y/qGORSAhfu66fWgMk6ldSWRl3jqDS
WV9g7d9jotiAaenBetg1/uqG8WZfSCJoVqQ+RUD1aXC0l4GVuHxZFnJMISa00TkP
ODeDGL4q4C2jNkgprO4o05fldpPjXVKnKecNc34U/Na/XHpDUfSxfDEv3SalYArj
DrPvl/o47o9pbBlk4gg2+Hv9971KA0gX/8a9PWW74h3W0hs4gFDVtclRHix8peRj
h2l74HzyDI9apBM6/EFZxFtltsa43M/tAQWtiPdA6eoj9WXnbLHFM0FiNOXq+1Vc
6aqSKbL8NU7YyOEk7atQmVvI+oe9jAPI7BXGTL9xYFoYv3yJX1g5J7P0UNXfamGI
V3AcGfXdF8U2kdB2Z7o1jZ/d9JtzNuLZJH6jT8bLdKMEWjfnn7Ki4krndBV3ztNp
O+IowYQY9Dc6PJMuvVErhxuw+L1YJ60JmZsW6SiAaiO+Xvabf0c1iehiiJ7HVnPf
B4uEnxKXPKlVUa7x6mcmK94UxXZBbYSzFIQgKEdXPTqiSqFL10t87Vah+8SW0HI6
ZrkISvj1tuLuUo4gP6R2vhNUfjE8mUJw6jolWN/J2XWsCKf8L2fldmkta+jIdQyZ
phG3uxjrzyfCVjLk1FGVpckRo4W2xvvHc373kptgs+W5dtXc0iweRt5ivvSPkzSV
oYFqM3pXk+kuI8TwGpoeOpl3NbAfGgdb5VKgpvEmaLVWOlvb/5lpluoVpM13yvG/
G247Ayg5pV7rej0cpJAGrhorjW+D9AvwOPdOK5dQD/sUZrXLUxtzcfspy9b74LGb
jFxRPXZUlo91yopF/k/LfO1x1QWuMrqQ+m7g2cNHG0ERWcmbsO8KICtFRJIJc7nb
O6d3+ZWqKfNbMo/JvqYWIlaMRQEYCN0k0p+pCgSdJd7GsiVYAHX/ZkqU3go0BJ65
m3WlZq0m9tVxE90ZPLFDih0ialKFztkS3FFygVecKN74kT9lLyASwyzsGk7nIcSv
YANEbyERoN1oV82MdA/KoEKSbjzK6DpVnodec6OTLV/t7KLGCkkS6f0EYV01RGw3
tK9qbl9RU41Xew4AiZBi4j+592y2glpDUnfkAoljUlflBEbBRFLBBtESeIfcyXRY
vqjjoVHuG2ePRGBTUDfWks2LqOo+0M2zn5WZ/fe9mMUL9bHcxDaEB1hJgzEFamqt
cArm5vW3/lNLzhfI7RLKMAZ1a6ipe5bK7WA1Ky4qf17+5ep2u54/t3UpRpsk/QIz
po5ntjK5MttT/4ntAfmHUGzHu67funYDrXlRq1zLRIUG33ti9nRvQafxsdXJodi/
PyDESzrjPm7sTJpKxP7c2crVj3E2q35MsZTIPjNkZiidlXvaMKeS8h2QaqZGubq3
0uRtJe16G4rqc/XnNfpPcjdQQLQQCZt2xanRCcPpQ7ey5E021iGNhOXKljbuu92R
WUGPDW/9pQBvn8IOrnXNzfodWyyzmxdUFONeRcFMIQOuheN4wwQ4Db6VuKnOQ0nu
RhGaF42DbR+t0oppe7VU2tufOTtDzvnKXiZ88PWGiX4/pcd2be5/hgVFWYR7oYKb
PpvNFbT/P3RJ67F4d/losYv7t6e77ETodE3rbCOxWjgFpUHo1vWRxXprrZ3TxDWj
vRe75+kAnHdrRvu6lmjx2cRYPYdfc/A9VvyVKphp6sl24dVpOkQSNpaYYqnHAPsG
ySK98+CLTJU3CRA0dJAQXLZMZarGmC0igpAu2LWKCG6bHwQZXBC+hE+fyl5CtFBM
K7sPw0/M5KpBJtFn22Cp8yfMGEk7iLJUXhCFtkd5bqYTxc7AP4w1zM/8r3vd+mbb
UficIof0p1Z2Xay2tmg4z7rc9aWXklJ0WdOdp+pswMCBR6PgA6I5CIwYFzCVvEvV
Ajx3xT6myDVmdv1Q7PZUrSPjJW0tOC+b45EcFqVd8HCHd2+IlGqQOHOgbRfn11BL
bjsLi0gyvK7wxe8L404kCzwzXnuBprNYXfLdfEEG8enC8tIRFdaHASXR1F8UqHeN
YP9ciH5pdJCHj5j36twBlvaHe7V1oTbYNC2PzhOqZ5JWCSTg1xhnRhKxRDoCuF/A
OsOAIepEVqpsXXPM3QRVJRzq4VEGFyHcg3vrXAKt535YqPh34kA6TiUUbiefms4J
Pb9lDvcg+YRkVuhXUDuw75ypBvSObOZJeaLVBf3waAJa80HRzwUjKXes+G/fO2J4
/XmYJU1JuGOMU7lUmY/0hxWUWkJf57ObAfkCK7m1dfCQkQJDaU/fbHfAvtvVS+1F
c17/7MhXtDHlFoWphRUZeIjp97Z+gzhFityztUq0RL//vgqBHktRX3P1La6eU31o
hd25XodZ/CjO8eemqVOyGdWB07aCgIY6Szv1HMMCsTcXyXzxIHN6mkfrp3NKR5Yx
8ntiOBrCyoSd2t0EXlD/FklSvMyeUFkWDRWb+QjAtMNePzqy7G5Ni8CQ6DM2p8rE
pIzyBdbR2DVXXtH0DB7WWNBkSYKbTieYWZ39tDW83S+7k3QyI9O32WeNtTZ+B7F7
lZ7qzxzahLqo9eqO2RLAZF2ZqdNjSU+HVhT3FINg/5laXJaZN5pxpQfts/QVwZ6M
29OwAyy/hkk99cXOEInYhJK1xvF3BCOrOy0PJJOAVscwpEdNZG18H+bwNQVVePVG
nTgU6POvZazSy7O9n98eEnnf1vwZ9Bf0ya+xWE0F9TtNZiU3pp4ScDXawceCF1Sp
KiOSlOIlgzMc+auhNRt+R093fKom0INtkBMjAoSWMUah4ouYCH+4KcKL8yr+Wn6S
Y1oMX8pJwzxwvmadxOrw2PsyRX3CWvpERaKIVXZ8YSFwDkGZGDqYhWJSHbHTwjc2
/IrtfoX0hA8MG30yR4vPenRd0C52EceXC6qbYWJOTrgXVHaXj+yCjKI7yJdCYDm1
oTanlwg/0QIRBs98EkDP7QIVCFKMieS0MhgBIMrOTB/suL/KpcNrvOErYAw3CQdB
zN7g8Jiir5LtSD/itOZ9axdTqC39fFkg8LT2xX5EMhB1RJBO4oP3vCI4aq2IEaMd
GTK4gFSQpJbfxxhwrWfLTYqVhWZSP++/BieTojmdOYuQH9wyF9Hm8h9p46Vov5V+
4Sfj/3xVjYJOPyrhrqGBMqB3cPYcgX8SIOkXBLLhrlAciSqls7bo95YBfvDm+1Z1
//z12d7e/husZZICZ11WtvwGJasnxWkzIJfnYZQ65+6EJbXbGu4QVhnbuOhrPcs4
sQo8gvgxoUY4/c5Xs2KZ37NNhnvbQ0Q2ZH0sLzNCXQNjHuWrYeDzFMBVWjIBc2Fo
9BHqpOVwPR07xdgazMhDwuFVju/s2gys7ILdVPQG9lcuUM+JZKPPiJ2tCdhLex9D
mWeCkiaExqows7ZCwZsZB6C9AoLLkvsY5i+aAPu9l/fuUaeQhtfuaH7HCBW4vdIO
76QLJoSiEwWWwtyzwdvAFAAbpPa6x724oOJtgroEiek920rHrJ5w28CX80ndR2YC
9qnwxqKUUU1u2hDrg3zNeznmGsjSTgdFVORbo+eD0gOc8v8uI9WoEMa5d17TT8gU
nUSA/ScNqoFzU7RTqMLOVSfFNydLyFx86MoSS1KSA03xRwZ3WkQx3Osgy1eP4dPh
cKaGVVzjMIqedMdZSV8e3Aaw7NaSwJd2E9jP+I40OwAO26KuVIxbhbZyeYu/cRAm
C4dvMFiPw3i8H9ia3yswiQnIWqEr13kh+gXI20lnS/unwNl88UbwAdYVREcRt4Uk
Y2wkDGJhCuP/e7EkUOyX8V7a+xWflKGIKQqUv+KHS+xU6nh55TRo6vrBYbp+dqXh
0sEpdKAugMb8AxtywXxoFvvWLtMZY6EtF5Ltep8KjgC5RkKEe3VRz64m2eHa4cRw
RJU9p9Mahz2U4wAZ04QHz0/hU/ifWu1oB89gR/nnNfPkwp4pbB/zaMsjFV7au03u
SL+L84Wif/j9mr4Hc3mUIWejYXbRhxa3ss90N0wWtFoS94GgRhOFgqmbwm4eupC2
1PzkhfQuric0f8nD1oXhgA/LP0s67ODSZMovZZmGnZbIOGQTYV/u0/N+N6Pf2e+C
RgCGm7NJvPbhlST0jdESEaQFJAJXyb57U1c2rA1BYdWMTVyQX0LlzYNRWLzKq9wL
TLowcoaHDc4Ih4UiOqkmY7KRVTVHbp/OH8IdCU7VTvcPt+2ML+3D2QwD60U1jBWp
LnnKKFZ/pSMT1WlumYwGMcxY+X7rR5SlVBQ0RwrDpQ/NfDHREeQVYKc5zu7DHmtg
DE0P+BzvnZdFTV4h/6w67mrnUHJbUADuCvMmBpYkoinTzEEs/9PT/oEM6+ZQARN2
aalMC6fTPnd5e5KrABDB3cgHy24+88GuoMBNoS/7H4lA+FfZfeT0X38/wgvOWnAg
FDQA9DlI1de2WIZwXqYn3Z4mPbDCMAMyLZ7nAoPXyHwaDVGohGGMPwTKuYOQ2VKy
UxvMnWsjjzEvlTjWWQ5aatRLIPBHXeX+xmXMoyWLF69Y7tz3qbcBnXUG+qEDd8QN
liwydaxVloK7Js/J+KQealPLCcr238rFfK9YC3G4l8JlNm+R96ngVti4Ku4DvRBL
8wvI8WOZc4quNQGBa/PwulIE4FedJMlzjsZL2JSXVcHBU7Mv9ysXCMoRKlFO4OcH
6YPOJYovabYQGbr7pcgWHHIUcQRnLcDyde9x42eOXetCQQ/Bt9KVksHAFlhTW0Z8
7IImP5/S4Lqs+L5fLtw973Bmdiqjiip+LB/AoYNVqiK5hOK2W/pS6MNJbuDPBFmS
M4lotXdIEC2gc9gz/kvYGxm8+OHmzD4mZ/hZq0tQO16L4g/aGFdS5oaL00U4lv2f
1K4TE3tjzVeFiBrI/68BuW03OHSl9L00vmZZdZKuUzuI7O+4s6GD9gEUbkl20ZmX
fgel4bG/Jkv6xqRnypkhDJhjCW+7qATNZxYixNrDTqdD7tb4SuOTYKKJ1/gA8EjA
VFYhjOvR//wSOSrs5TMYXDj6WpjwMN2ISai8+68DDy/qvi7cZRitXHr2aPzUyQhT
MEnRcEjg8nqpcKBbbH4jrloRfO5YbvcFhGc96ezMkCua+ubFQm25a8UAUr6xhp0g
8WDM1bQSREi0MvHc27LPR7l4PpokbGQgICFT4hKAr6B6Pr1VmefZlEz+aUcF+gf4
BXXYv8mCNsdBNbx1yzgGYu+xo1fOYQK0B+XnApUHXEQ7AIXiP9NM6EM5O20U5obR
4q0YePZw5TYAC+qEC9hDVcj33XAjVcs19E8p9PQ4U97+mdOvw3SLsyVqtx4iMtau
GasP/GmyNUqrcWOnEh4zULZxT6yTyLzy1XpMu3qcacKrYA0/x4eK0Iq7beFWGv8a
9pFLNd5MsNdn4bUOyE4SUZOBV4wcsVeB37kdloh2vT4OaNbkSX1YiQoMc9xRJmkZ
WYk22iAedziV3iYW1v0h2D09gONS6lD4iKQ3GZ1n72P6WJC+mwLteeMNPADZIY1I
GNm6pfTnnfYvysbsAY2D49z18iRUC4VisQcFreQK7aUIUJ9BaVb5y2/DfrqmqTJ0
6B2JgeXW07sW1Cd9g8Z4kzFcquss84qTS3D7Vq3sIbZ2+wh1fsYJ3M+TAY37jMCt
U1ayOIDFOfz3/EwS5gXtMpRtU8aaHQqPnAKKJhsWY3HC7wKUVpDCiO1AmZl5iztA
fVwq9gqVcRnGAlYlg7++/8yLw113qx0930ypRYOtlAkCdCKimEWT7PIu6sHts51I
HDYBP/tKeGDxVhDJIgOctzLGzHCkL6TOmT8c6NCa6QJKVPuMpw2PE5vyj2sQal8l
z32ezJchZTXVViWywEhCc95ZKH2iR3EqMxI0ialpVdRCNv4+pelL+1XMGIQ2Ymog
apQMvA0BrfXiEwupzxWZIUPArSOOlzbI+mK3VSKLfAqahmjrCN3Wraga9k71pyQI
fP5hXYoSXP/w0JlTwFqL+OsKyUgMFgb46laj6hnWwbseOmpTv2jv2kBkGK+jcEmo
X10KdjpCPaWtWqRkF5tP5gUhwZ4CK9iNChK4g3PfdxMm2GNexcRZ5nnnRQ0cdBg+
Ks4LrHV5FteZxz6nzkMX1l7hauRdiKWjA0aFOuSLi+9M1SuEzrhJJPbyKVPr4ZPu
wSi6qwH+yuvJbtv133/0rLmRmpTBKHPb2jlsxY+7hY2U45zER9oAZm1/ucwCCw/V
XmOR+cWcTIvn9KYv6ZEY+nsBWntgyRJNsmkhLIGPFqeRMHmReEKgyH+HpYFB2KV7
+8RarxttnXA577fut24BA6Muk9Wu1nCQOUXSXZiOvXIm3/C6mnwCQschWo5D2Jt0
9RPM0+at9rsKks961VH0K0SL3abDdbUsUUQ63Ai3Q7QSYxKk0JZf4f3aIPapTkiQ
weeNKr/VDdzQjSEpHpbn/adx2yFcTDZL3+TQrGRf+3jIFYbEBTv4Oh3xc9CbqQEf
IW6Zgub2RBgTddC7x3bVoVpc+d7KIXU3q4OkqUuHnJ+L4sA8zpRh3NaEkk+KkbHi
SVUQfxGzcVK4Y8mpikKHHkFWpeN61bImG+K7nUn9gc1GJANJ6diLWLuoBYjVUOWa
mzM03X8DCGqB9L+x9HSZ/QQGhVonr6EBeUH3qs3HOCwKt8TTpUtwyf4f3nyscPti
hWzXk07IO7VGgYc6lNG3WkhaGSNenWe3GwN7Tw3V/LF+tdpLKIDBqLL3XlbEndOd
Mmcd+ndGJKFE2E4p17/purJFQRfijEuj7zKZ9NVuE3OXhk41tACPo6OSCkWaqo1n
xBZabb/OXlTiM0gJUNbIto52JVmO91eGgVSh+rA727Mob4/wk3ksZ2ED+tGimrdt
DpRQHS/d5UxIzXEUELMV0PqgvOgpR8G4YemTsvCZdLeleC/Zma2TfPEbYCJm2R4G
F/kefs9qpChFBT1+LDhh0z3rovURpUZug9u1TLdCaazYi5m2gGJwzBggCrL5CNHV
Emsd0hPeoGFyS+kJx2gfGM0RMXG3AqCL9OCKDXELq3XFv7OwCMMf+N4yzdvRY0DW
QHvwReldu3zW0SKZlG65+xwNO9ceD0o9KeUr1RsVRSV50LpCn3Xg5l4VB/Bfe9jW
D5mYCNyRc2qm8t5D1/ZVviHBPjCwpH26McJQ7nOqdZHMQDXkesSh3norMZlx7jpn
WYE6B/3sUDn4+tWzgYQg4LdQIUBBDEnHB0J2HluOb3hRIHwJE2Boq0yBoSqgMmTe
4OHHpNylLwUZI2kgzXHzzipUkoTrmD9pMUgAnkqJWbDXE+RrFmQjk0E1SbLQIhLj
7TtYKwl+hgGoMMwb2fRaOOxEKjnMIcu+l0wkRU49aTmGqEblLdccI9QJT3NDFT94
ZeFHrvczB0XhHdbtlTWDagi9mN6WGpW7tUraJzg3y+WI01SpHNLTdBaHocfBCd41
Ow/9+yV0vbMAcNNhKxHa4/9Nbc1KXykcjrLcYxVvDH07MS3TE0oyrYZaLLy8+o47
PlCWOnBmJlll6L5tDm3l540Y3BTnzaiX8IPkfZEh/YTEg2yYmua8YxFZZs8j+WEq
H12dsCpt5kOjNUcAK0yKCpv0e3brxAMvrSZz7ClpVvnu4Rc2KOCeDvs/GHBVMWza
MjRpGjbD2Z2reeLR+6yU5o3IVn+MP5GOD9baWGe3upzA9tNzNEvjp41Bo/5qmXc6
gRh6Bo8JTENTa7eqREliRWuAI3bw9Bc9U1kbsz6NfPy00G4SRRBgtU0rZdnQQOFh
sbCbcaF4IhYZ3gW57Ls4gBczOilSwmgmNsGwCYND1PMEH5bLoSsrSxhdcCZnyOVO
/TlDEs95cM15yMPYGlQcNVw097MSPkr1IGb/f56d/hHYH3PO56EeBFeQq2kz46z2
AOZR9UyT4T35aBck2WNRrn1oRR2NeobWhvYyNbj1XRDDp8qJ+yZ47B4kw8Z6vco1
n6tU21dybYOzqFT6rygsJVEG4UrF2x72UWUEv6pB4bfS3m/X6yv7uaH0YqK1JrZd
vjX1nhwZbOBvz4CqhOCE7gXdAVYfITB1DNleQ5MZIFmFCoNwZycxKjTfvbTYFzgd
HbMQRpOO1iixIFPVXFTX9ovTYuI8IxXgkc3NqIKWAQyja16CaCaka+50kK0svymt
nZM9DrZRzvutOqddQmy6S1LCDv7yIHsmpS+at0fiUzIoeq1T6bEum/f3accJAIVy
20qE6XeD1aBvyo4MI6lZd64FKxgPI01mL1L0/dx9bB/187cxKW8wg0Gb/YdhztaY
NGVt6Jlsux6c/hVb4/WCB9K6UAOmyEVx2dnsul41XEttgi1J9VQ0XNXM5FWWnHQz
iXBcJEdGf7a38mGUz2rfAZD7xd7Ht+k5onOkSXtuBCxYRp531N5Q8TG6O/D0rGIh
jQE1iGhBv0kKXTIz7eYChc8jvVNq2P7MPtX3TzvB9ZzVzw/Lytk4cwkkxPw7Rdjx
HvQO2LTrPO4dG48W1alwgRuTICyM9NyzFhqGemUAdJMwVE9cua9oV+S81xOElR1E
rlfF/2MoOD7F7tl58gJ4LTyrw4TqRJXbnCPk0yc2/Wi58CqXWdYEcXCEqLXhcxGe
F0UVVYDpOTu4DuyPgfmQk9XsQIA42Jr4ceiYMA2TsjXIWGtm7cot/NYJ3JCodTbA
sf27Z+x3/fF51OUTyNYJg20tVZM6hvGZOWGNTN2PhhP+dvd/v+EvrnwTxeFRJKe3
z+k3YDZFLGY4UvtDt7f/JYJIFmr2Gh2KZk1fcban0ptuits11+U0I2/y57+Xs3L7
5G4vkUFRuCXlYE9f1dGEQXYO81Po82H/W84B3kfZJ2YuJt3noSsqc6h5TjAye/iV
JtzDBilu8iaYBqXf334wucm4iY9XQJLTIyM3Mi6VGTjRLkHvcnB35SqnXF101JN/
jOsn/HudKFUKecteCRc/sOmHWig5yHAQ8bS3wUzR7xG/FhgFc1n7cLeQ81EivXkr
doxZ+oikeWiRVCdMfLlcTsKKIMmM2zttF0K+y0BsScQLgID7nOqHY6NNO+htO4Wq
RSs/f5YzqAaBP/hvoWta1+qOhOTorKNHe69LyoIYRfrx8HHWeIeaRO42I3gx+rVC
EwZPOEaJWrwrJILYYhZ+Rlk3/IIJPpwcnfmRT52wH087HW6/sxTWqfQigqcpdHpR
0DG8QZIiTlV0DSB1Jx1Qx4Z3wNmq2QYqbv7gm+f8zXulZCrl0XTTChhbFpI4oy2O
nmSq9vs9pvSDd2Oz+AUQG43nVMBcnGqn8csEvcExSpu8H3C/ojhJWmgt5yV4m0S4
+gET0zy5Uu2YHCxlQB1THzzVCPTaEOMiMPVGVmUCyhLnvP8Hno4aGXtLwZcsupqm
g7VGHWhLh5NNvSmkkRuydNf2403QpL6CiwqRMNXE5VbThLJ4KtRoxQxIW35Swpv0
AJmI7Q6qZOWzRIZMzLiyCBK36h/vIbyzm778RfSD8d/lcnP8oN5Sst8qpH1x1U36
qTzdu063RC/NASzIRzZLYFCln8icLQY2R7ewKDsjUE/jpAw4B/QhZhPlwZmkDPvW
GxlChKOLc9IXdahUYmxJuKjC0n8L4D4TRO9XQU6CHxdjBbMJA4ySKjxd0rIAnTR8
o7H5FoWJbmP3jfHb1HEnlm9HMBpzpZM/zjlvY7AisL0Uu3Em5bJSKvXiWmtSrY/y
r3uIHJ/6807iDR2HouG+YQhlVg2cjXcqpngIR5pWeg13X97kvRfjGJgnsTp8Jg3j
0NtOGaOa3xStyVGNuQe+h29eiejx0hkKu7Pf/siOhqAu/YiD/jenGuU55QAtetn4
PjYJfgTzUwgvrZdhv+XfcVKlglLMiZzN4OpOL0ql3ggkLa+mh2iFhXeF8ZXhR2zF
1ia9N32n7fC8NpS5EBqwqdgzIYuT4cEWSLxS0zCjZRvDnEf7t4sT5DkdXg7BzNXv
mndjV31VP+q/C+Gj2V35KyeT1P+mN+eOgxgDYeHf4QhRjXurTOkcDbgJuwy3WEuR
9G/nUmPODSvJdviKvmeeglUbJJjaKoInfqf8PZy4v7rDTYjGJMQuwW5/xtlEveoI
wl2Xv8z0OSGMNl6Yon6gP8wlr8G4LpeQ3iG/VwL+Ni4+OM1JVftG+/DoAziXegvA
f4LtoXQDtUBgPAUwVFVcbsBGJBD6P7mBGPNFqYhbbR5g6gS+l7JARSCMUNhUOCQ1
h52mClnahewE7PUKpOowHXSeXRpCGYj1edZoQ9gNT+PypfeCqrZk4UBRPVj+y8Ei
irN6jIDzeYI0q+oZmScSSdOfLHTMzcoQzmdMPm+KwUHZPSQguO5BA8d+ntE+dU4x
ugCDOjbb5sNDdEIopTi1MxoXf7fDVKpOd6h3P+bX61ZT66Bbx19kmh5vuT8awFvo
Wqr3PdS5iou2bSaQBMdYi2EaERrVaBCZ4iJY5MXyfijdjEtCOCXn72IqLomly489
d4TkiSxxLf+HB06UQuHaqr8QZ9jgd1k1j/VcMvqdn17or01xJ43+G8BJECCC7ni0
Z663iH+YX8nOVvTcar36Wit/CCR2wkQnq6wNeUuqcoSK2HyvX4Bi5O3yciDKYFYN
ZHUc5xTHsRUlmhtjAVnBSiGmozokUHYMr0ZAiM9IkHIgPkQzc3MWj+mdKSq1bSgA
Ob6qr342mpc4vS1GBGJXOXFxhAMUsd+oX8iw0B/UjMqXzjPyV1JhA4Lq9Vy3kBIL
l6iu8P+rAr4i0Tzv0x/w2fc3tnPrFnndowLFnmSZcMNfcEO8GWrp9mMCdp+stOiD
z+RqIahU2ZqdkzqMJ1FDNgHlcsAPJRvJn3vEiT4hD6WQWtIiRWhhMFSjGBov1nxH
BKg6M5LzQz+2hKTkEycj2adBHifI9Vg+McGTVUVQal7SixTNMuGE7bax+7Umte1S
pnRL3y4ircjQUfp6YqNCPWhqX5MVPYJOJzPL4DDCv46CWJTmBCJFWK3Z8zUlzGVX
TaFg26Uu4sfDW7bjgLz2XNFOdkemjsbSKHiP82HP86fcu5CvRKFzILCs38gEgZp7
Z2WIxavthd6HrcWc9TfDD4yfU9JIJvNVkPJTtplhJlGhRiiC4UWJ97NOnWMi+O2y
vf/knoXt1tRzZd/xNW2KQaQMD+zcvAcNIwqamWmYZg8eQqx/QA3fuEnjcc1VKlgt
84/3xDdxI9ONLTcGYThsu0CHej3qSK0wxWSTXXvpWPf+xx3fGXKcpDqzRf7T8ul7
2QxoEhlH7F848dfCYbd1WfM5o/GYKl1yN1f8a8MhRH1nVCw46UOuK/8dYhpNQl7f
w1mAFRIxStzTL/Q3YJuT3R4/O4JCH7o7yQWyq/dqTqcTduO6Y8rQqgZ490CNKf15
4oWxMXA3t7NkhlkBtxghypW1NVWf4eGckc72T8kSI0fO5EAECNPjHKMslSa2jlVW
KXLE8LtdHxeKPE3qsFyGCGCyYzzzgAziKK3hvMFE/KBWhVQ1xuuh0jS1dwSs+1CO
rXgHZvkB5lxzmM2jYi9S51vB11csNN4QzFIiODR3KxGE7Jq303rVT2V2gvEZulZL
y0DJ1NWdUozdicOD3PXbgSX7yTwG9sqR+5GcrTu6SihAOYHJp7X/He39QjdOQ+bP
GqAWyx6HdigFLrrT+lCiwBJPweqm94mDIK4JXzTt8hTNsd1UybEEvhTmNDvvsLg2
PykFW2kRb+smcaN6igItko+nhHnab7jDe9gJWkQGJXO6e+eLOghMnRTJYRusnBMF
aV2NOSHQ3oqy/l9y5K62jAlezTLUZAZcEKM57NRD6chJ/fqu0Kq7e/RSY4pKrOqF
g1We2HUdFpCh09bRhFibcWoNIyTWPtFY9Ix2pY61lvSZq2EwH2hsUTZ9Y1bxOuJD
auqRiTqkrD6fPwI8xvvFmcXMIO0FrWOIajGnWhBYYncDIWx60YHByhao74OeH/OP
+dxiYi7wOA1zVHZtwAULSAml+93+XFkpsoL1DYDQqnSyrgLBdzhOu3RQwelCRIu4
UtE2HNiqWD5lmEecZLGZh49lkt4Y8SqPGhLic4LKhPiMoLzEudgemx+S8R03h/1J
ieqwW4I1XiHHs8W4k7/urNdczqXsezW4OkvXirAnu7S0aPcKplzWlP/21diCzw2l
6gvr7Olc4qV++fCIN/iJb7t6vuRRib9VJskCqa1lFzU2TmoVij6d/Q5gg0pkU8tL
IYRdzFjoh3O9IBiP1HKdBnacJVuGWdOI7xe0DglE+rYr8z6TGFXbU0/M58szMZX9
BbNK77kBt7h0lPLmLUxf8UaZZQ39xMM7KxX/mOSz24eil7tx6eb2rGtmrRwNE+QS
nlbflzEfE0wqJcERTePghGb3vNIvyJ8VJMjBG98ud67OmoYKDte0efVNH1h4hwuf
4Tv5Rg6pIc34LdgARL9PsPBx7ayMAbspy2ZnTeO8+eyyavIXC5C09WkJ8Zt9gU1X
sTI4Qq1GcRw0XQCmveYLNxcMGt62IEsKOhuj2mCpeIpFADALZXhKmI7mvgykECiQ
gZpTZF3bYKKkSAX+OJByjLNxn3t/GcEiwnGV9rLsOEUbCmOnUvRNJRlEGceRyI6h
HIZ8aYkVIQHAa5JN52hf0voQ8VBfeupOitVyp+op8IiQRRYZA7oQ7nIUrg1ZVmjd
ARXCRW+wZeOSbAVnkXGqC+NeDMLUhylvhFdVCAZHNicoAJ17UWp8TNVi4DiR9/4D
kv0g/VQhLeLf3GRSNa6zTyFj3j1SOr9lenOmR6bfsTLPJi/+k4u6iDw8FkZypxQz
yKJRyiUm9Hd9DYHTxCmKEUK4MErYOST+wPVQ3wj+k0Jj1tjJZUhvxpjgJ+3+2qtM
oItkF4cbU4z4FBCY730gUj0uWUHmP7wU1SVAJNkpRY/ZiKU6/mnxOmapZv4fhn/f
yYc3wJsQTlfg4Prc3Jm/A4k03fNxB89fQwZa6Z/yeXyQRFsUIs4c2LAn2VE34xKZ
p5D8WEP/t2GN8zavYWVXXBtYoJ8jQ+dFmFKup73lY/wcSVBAYCjbUg2S9kUXQEZ5
z7GgO+/I1qgt5OqQElbJRy0LCzxd0KLPmPDLUWlxS7VmIZCYUqoE1HvQrJx85dyv
wxCnYWfQtkff7a1pRLzsb+NXDLNQizETNGxhars86+GDUfdVZRoZDVFpbEdeq2Xd
HKIQUwX+rxHdXa+ri2zzYhh6M4XLDjGghCojtZKO8WVkzr8BsRUECcaoqgE+EEIt
wjkwC6EH3iXsUcHRX+DEeKjKufqzrxU7IY+b0oVG2gqOCNCjUvfqRV2iHXNSPOO8
wU4rAzKfbCJ0LrvL4k1eev0FtJlc7K7IfZKNFKBiMCXDs2RKSTnMJl+bXdINNOlQ
aB1VWQG86lXQON7nP9iRToqz4Q6HXvDS/1DjSeaKgJWW4zN0QJj0pcgPdkrSuFac
/AFSwGIr4o4r9R5d3RgbTU+gidYED+xXDpGn8P9X0+n8vOBD4lYB9FN50TzN1w4y
fKuFuq2g0GfAd+3XC16LhTirzog9ki0qKoqr0C+Fcz5IjHoIxLW8X71GIGdYBM9E
/wFP14Nel+HjlP3Jh2+ci+kxyCyFSBDhikbZ2RkdYLYfg0CB+qIZfwBz+1OAS5OY
PnGiYWXvP2xt/JEEGdPjnCKE2swo+7jYstBRnnkSeocOS94/aTF2EuonUSBGJzah
EhE+CnAufGXxP5o0Y6cMIq2q7ngqfZlzImSOYmhkUoGA/OGe01oGqnXzSobaXwmF
b0wjkZmiGYNkfqeHVKDez/BUPgTZ3L+5g3EWsXUdsjsuTB9eeRhNeVA1vTenEwVo
dBS5x/vQRnW6vaThwnwhkQ7nMeXl4RI8e6sjq6+3ozowjOM8RRdga/ievFAegnvM
Fgla3Llvlmr7eQ9KhXcojppQdSOikbsNN8sFbvf38sqDIBWP2TbXC6LRnUts34tB
C5zaoH9Tfd2qBZqat5QV4tJRNCQ2EkcwTg1H7IqEG6/FY38Qz2NKdzf60SiOvJYw
/1I4tGRCRK8EWN5n20U8weMeMObC8ZXQxTkliwczu1n/Gp8dZ7kfOBUP1BDuNT7Z
GeeGpLl0LKpf8+x9UoIak0rlT7iRP/d+tTHrX1BZVElLPK000iRstn+nBPQg3cXs
pN3bZfj3qVvAZGlbbkcVQjacrNrfZQMnZXbhme4ujHGfYxtC2HEn9sXhoOfg/aYs
Qw9AD4OhhxHT0WNZgpIOOW3J1u25jTQbtLyq2d9BZYNcoTTDUXqpfeE2wtp29fmI
YXEKAivINiChzaqgzmUYJFynpdgC+m+CZ2Dc1/09H+CxB92ZjPo0BMHjUpDaVs6p
pFwudq+DIQCHZrNkv7m7DihDDAK1k38l8AdQHKeTDucYUG+qM1edoZny0ww2D8jG
479nyASX0T6jgv5D7JTv6+ZYB7T9tg/Xt7ZQvnV4cZvtZ7HSEimiAmbm4df7gAu2
ACcNV9i0XYjd8dS8Kvvx/bdxX99ZpJ2TRavkuAL5ZdPXoAQHfMWk/m5zDsRSmYBA
j4xb19/kmrvxNgpdkd7cpCv36vwgUVcJZWUIkYYz+48LWORoRjSrVOO7DvGJWey5
7SY7PVAq343n+XUwdhcpiq6P82bk8hp/rYbGNeUL3d4Y8lVfRAVrWa1h+Evxbrqn
AILslxccsOMz3z1buQeL79tcizgsuJh6YygMRovMtAt1kv6u4NWdKQKxVK05sTD/
ONkxJVJ8cPAjeYU8i4/CGNjfLA/mNx54Z9GxudjygT30s0xhfQ3Cf7h4IjLlwwtA
DdCLZs7Z0VqQQd/6lQwTL9JkClYyzLlKMCsBorpS94WU5JI48qgBMp0mhdFQ6HFr
EkU3CoDEGi9lZKgUfLGIEPERsQ5TPh6O2FKOrx/+Y6tztpT5dVEycCh3QATACDz1
NzjTttS1EuVq/gEXFhAm9uNbq0wGWyazcWSY5Ge4Q0vQHcUlU5F86l2sE387K7gJ
c4ejcS4T92Ydm47KUL78led4jxao87y8GXq913tlnJ/8z+sFotOTG/Xz1nivV1Il
hkKZePU4u/zg6hy/mk2sJl9Q2t47DajI897PaVqncgAy9RYG3+IOjI+fb8E1DbI+
hfodrfUW8hGCcmTHaLd+nqbTAXuHDb8Qa+sYN4ok4brkxtOlY+RPB+QFOkyzAN6X
1kDTtKm+6/Jti9ouHhumYYuFAb/K34P84coI4saY7R1cH/NvlYdOfZB5WFYWgPBh
LqC0Jevd1N2kRBtRMT32GrDfjCfoOFQTs5OVjd5CUjQEhu4GqfbuXd/VmO8gY/bu
zjZ7deLjXLANQbIx6iqzr/LxMn6Xq31kCTPUOoZGeRcHvLcSW5/yn8js/N8HXYSB
ctQHlTdMtHrXGpz/clcWAg5PqbMM2LhxSc/O5WsMDeT32P/Da29cz91VBIgoEJIl
rQiJBs2pcDb67onfNPa3NOUpkOla8N52fvvJlquGsykg2UF8BOU6Nf38afjjSXNU
FkBKoHxdfjR27GbqnVgkjZb2TiP2Zg+M+oa9dGDtmE5rYqgmJWtvHQU73tsjp62i
LG7lhe4hTaBj4ANH5zuaEdDZ88AS06MDnmzNk3cWsBjnqyIkocc7LbAa6MHrD2tC
x3cbfriLuHufqnpY+O+BBNk9QgbfW0HU6ZkuHBG1khqKS+iDDf5PPrCiOdoOziHb
cYoULtXH6h1N7XBRqBFj0kqQela1s8js9PRSFz6YHKNndfo1IY8gn/uEWchMJs7B
sxuSJRPFaIi0BSpqTBiGeNFowz5AO9fxCMawNz7yp3J/v8iA3zoPm/Hj+UhmhaWo
PVtQNPrCG1AwXER2+wf8W/kJ6MDWPz/1w8V8xBxm6k1e3zF5hpoLn2bAEV8p214Q
BHMlg0ZjukGdYKtVgGYk0xcHMONj9mhr177PpbvPTkQyvrYJJoSIKr/nezvD+oBQ
KoNkXzkcWgfV4fa4V0sqoZBTqvJzM2mcQsJaFCW/KW8F3GMz7rvVRDDtp7spxB9n
bW/3ryGj1XMkcizs/s/hSjFqPYdEmEn4yZ9PHxFHTuexmO6wd05X5kYY6kPsp1VX
0mZJBreiGX77cUAfEByhU/VC68eEBnAZfdHCkFaBJwXIr80ppnm32N205dGm7nj9
p9JkZhnJhiaXEuw+EwzZ+YX2BDMiw31xs1Uqeg3gZyUaVxH92nfrseTTpgUnTKQl
mfdZFwLPSSj4yxfLFZFS2IPK7zJTr7/LubpNm0a634Lcf99TUllQSUtGzgUsO/on
HUSARfpMKIoiKjB9fGpeJJy/0QPqWu2OGzCyVQ5ZNuVfhLrFGjgX5daJiagkLBqP
aPfNqtYZ6073MWs5kX+YhHNghCTYgPYhWhLDiBg1UF7pBwAWYPGmpas7ISGRCo2Y
VcGBbGu07n0qfwiEjgM4VT6O77EDD+uKgcP6xpGkbrk94Ager0q9u60FAHD7wVGo
82BlrHpQNZoeyD9rShwfBu6pk5B58O1N6lpmVJeLIlT5sX5lvBl3JgtbliGvm4E1
Pykx5knviYqkxzrvyIljzkPngQvy4aac/nB276SZCSchkvz+rA1poBDEW9/ksL0A
Qn4ejhaI1v1yGtFWCg/LTZ9Xj2xAjCAwkGyMg+kVuPC9/tthGo28oxv02c3O5oTO
m7WVl5TN9cGL9GIKTQ/j5p2YCT7wl+51JYNXXZu1v27LQeTLIkKLi2I4KPqYkTWq
tEaK436kiRYMO1hPqkSakoizyWGyt3jTIbUgsSP0Tqa6e6TWLiMPtmqDBRxGUXhU
0mUPZ3AKOl581KIAwclrARIovUKRAYjG7OagsYTIzYnyjPqFvv19cJazZsVQkFLL
jtfo26EEXpgob9DNQQJSuZIftDt2KWLcuZEpO+Bh7lKySUQvLKovDzEPq5iHAh9u
kV3NQAvyRyhzkdR61lBTfUXXIH+MnocOm3c+gw2rSqyRspziZRLYhl1tA20LqhVz
7rsWKEjIrMf7Gf2NbffX5+HOSbtPA0VOAxL812+Z9KY9JoRgX3DP4RmDTyrqg7JI
qnCo0QP+t0tU3DmetSdoCm0e/9aSEpM2mJeJX0AnjDCoFYz9XZId/mfyF2+gQjgL
bWJDES2g3xp0q9zeup1sFk00GOVdBptHn7V3sof6HCBI2GQyl3FT/pjUlb/PHGSt
7TKXLBHjHar6UU7DzZpTLA7g4FbGA0hrbfWAoY3QuTulPHhPz8BCOjmp3cyY3Esc
0bwvSSjhWhkhV8xRpskwC/1aBdaNjI4zfFNsFHXtcUUw8lnTUN8qgmW0H/4+6t0j
lAeT/ZsVIKx0M8pdcLqTQzowxQCShAmZljMtd+AW9HP5Hshhw/t6ukqFJ50G0cfp
N3rRgz6dksA6VQLsWFXPm1jnxrhtkzFfFoYZUPjTuxkMxe++dGvcZaOhWJBHRlEK
ayju8qte+Pk4TAO1+Rla2ohTGXFqF532ktp3Lge4f2PG6/rYssuSUGzY7InWFnCn
T07YzqtKxhYBsS3vO1imKXNz3PuFA5TsQoZEqtdxFt2ElDCGjCTmd13APRgVI+aq
U+PPPChcUsqOPp0hMEXVWPn0DE2a28NhEmCEcIIqNWUrnARqSVaTa8jI9S0Rk8Df
DuzMu+azXjyQ5S0dci9hZs4wrwmQK1cnLfc/dZIYX7u/fnajGTo3BArSvDLOBFWD
c+Rmw2aylhidX8Mn+3ZEU8EDEEDvGdOV/5PbcXaGE2Vx3Rs8ecas8MFhBK8C6bmg
u/939TRCG34my7FjYzUNBSEWJGBlOBCajiNNjuyXaBew4wjgGF9BXzQn5gXF8naf
kIILgRRX2aVwycLLakd2tDqK4Oe0RMM3q4kULyv2EJmlsQsyofGq4KPsw0Enxo0h
Basv8yqAtlEZESSstJlPT8CnD3C57ktcGjikWN+RTn2xyOBSkewTGapi5gHRtEL1
8sYnnpjD4ZLOWRVBIWKHEbGrV7sb92QaP1l/w6GJhHcOD8VbQ0qofv33/63tzlmU
nXQ0KoBDZbtDNZsKrwpds9gwZzdsc2aj3rhfe2tX8fvN01iHY4COfQW2snFmOt7v
vjTtfDz6gCLxCFnLYeZpop6KNO+CcOJNQfMKBExhwpc4toqv6ACqKz9ZmFWjLAZt
EPjhhqkMa+HjYO5jp1gMS4NZC3wCqLlaBzvLn9FABP0kPtjNDRI04S82C41PWvbV
zafM1wRvNeg6lwa+pCYIuybjt6Eu4zJVVxhq3JF/uscVPtkcgELA1k+WP1b9mMKD
bf9dslXmEesoVfevHCp6qMsY2kVpYjZUpAAI1yDx0U6df8eRBLzUA6Hak8TyvVk+
ogdph959SDCtXWU+qwVUsxB9eheRMEobqTyXpI30pBWAxSC0EWrsTqEuZaXxYXnl
oZASbC4R7KpT3il1aG/+hUkCv+mKhnU/5KZIkUC9VcqTUzMIv15P7o7P+V2lCJcS
+4Nhp1mhLOhjObcjFxZsGIjZObZ4pvMkzz/Pbq47Yr9T2mMsxSxgjtRaw3UYmRiD
RybrhvJTIFm4xWLBAcSJtC5ye7mF2MbffATjuFiWXDqJ4min5XqB3u5r/Y1iPm5r
0tzY+Ffi8clshrpmy2p46tFBCMBa64AsauGXs0Lr4qr1vARlfnFiHWTrUIOvFyIb
ucON1lpeJvm1G+k3kjXYkTFxzo5lk7S0hPKfiTL7sGNGElMc2Ufpp+76rzA1WAqm
6soqUsG3USLxjfNXA/SCaphjJ2oSEYWrXfpY8N8h4o/OumNl1bft9ylMN0c1PVAX
JTF4GabuG1zV4RtCQuvaClLrzzP3jB6ytiR4MuX6ms+/qWlQj3EKC8ClZ4KpP54I
DWO7TsXDgRt4tBe3qrzqqRTSkxVdrONL2Zwc1CicEVHRRu+t5gl/v2rLMV4QW3x7
uXVrRbH8JIAPGD32pHCvKm94Tz/wcH1BybipMblNhe2+ZtDzh5HRhjw64OlglI6S
ZpCHfRBKqB+4rxynhQqdrKcIEBBfBLjNX17A3Q1DSHnswqaC1Flmxd5bYcgBYxMg
9cRvAEX6e5tLQuuTSH03oUk5Xg3fZetYAqLdHIPTUqPk1Lg+e4pWSDP/gPxKlFdG
4Nm/SG4PQmkeFOiGERCoX1j4QtsmzxNv2NZvXqe+DlmgPOtTg6m9YfKkRs1khbE6
M3ydX/1K2e/gbfLCZg8CE05JhstRoLRCwAnQvtW5D/XF4zQIMQ1EvP8RobSgL8Cq
aH8iPn9J79L6MIZzptbR5zBc2xqBiMvZ43CGheOfPeh4DjBFFBwwmK2OotlIHmWs
EbGUsqvO30s93Z9fCjzSz7j7Zv43MpQ8Zh0cYnGCNg7eS4kE/mKgA7U7hsu0Li+H
yQje1xkbPy9e75JwXhYi4phgvVBIV1Mp2fGjOB+LyVhps04A8Q9us2kEKqT26Aly
ha3IMIAUnQR0G0kD9CiNlGl7FP7HnHQ8lhQ4kJHs1EGDzP64zUVkMpmYTV+SoasP
tNbGouT3m6hmy7VrnMpQZfdhfGRfyUgIA1pLDnGXu8nFq8xliRZ5dfBJ1/EiWxdD
X3MfZ8AQHuA+p39U5DdV5LZUXHMucJGrsyk6V2r+mSja02QxtlufUi9yLvVJX1JU
k9WQ/E7ttDj2OgVTVzXwYrdacljq+7AueSXxFAkdn08o3zES7gEj5OBUGZ29oDfs
/sCCxIozfCFh8/viCets760ZPWv7HPyaANPDH1tyfF/GPBIOjd0DVnaXz41sdKZl
dHlQJYKxqcHEejg8Bn2qtH5PSTgg1TO1H++OdvmOJ9tnQtyjwMz8WjLCcusKzaeW
yCCuhBzhuKVATDLJw0zQjMOEOKMEpqVm+SAb5gRd1Tca55thcKVCIg6U42eFlOeC
nMZqydFAF1NHQuGWzYjEcEmlwniJkFWtafDQN8ZMZutVFkyPgXbnwD/7C08L4Cat
I7aisKWIslDS9bBXIbkioIbfRZVYqRz/NUIt1c5F8J+yHXXeqXy9yxj+ARwSbjSq
PkFJOW1adMZ4Y/SqJz5iPkb0cGWPLw4zxYx8rmGCM4t1oy3Ii9gT/Ravrs0exdZb
wRBiP0qQeyQ3QKIpniih8PES6TBoDeSg9F4YG3Xk2KS/pWJpTHCHvmi0jlyW3XQq
fD+FSRlwIwJn2qYVSyQ8ribv28E8PdDvoDizyBofWa6l6aFoN3TzzzdqDGoHHbUv
DF1VBqMzl50fQ8/4rFtx7Kz50r0EMYDnoozLQaga17wAlTpCTBOsjtaUVh73I16i
y+aB0x+Yf8AFISR4oeOoDkLHld55/6MPzB2mOrZRbSK/WByc4dtz2U2sFpmuVjoG
FyvDQn9rzaFc8ZkyiSkyTYFSYOrSofjWCRogMXxEthdgdo9Jf0HaX8mIZCj4rZoZ
fptI0u8kVmoSaKw0+VbqXcyYGPQL56vrBF39vtySTk7GjBJ+2W4rjxtueFcdA5kx
Mh3pyTnYZ1y3wj9K4Y+3X06uLflUnRmfA5ADeUbZVZX/sN89zR6TkD52VXQcsPVV
DGwyVdiy0dJDpblCwpYig1HWyYZxc4+2brKwCU3x9HwezaDXFB+tWzlnf8nP6/hZ
v6vCfhy5CukPfiAp9VcmJSZTG144O9SM3Zxj5t5nUSl1tCtXjeF8JQKthoq6QFJx
vbcbh1PLP+BU663obdZUn78X2QoqJbxCuM6/tNFoGREu9bzJDWo/aQ73duFsMc5k
0AxgC64BR3BdqBDxN3qmWZ0Go6Y4FkD2oZB7X16pJ3IkOQlqLYWvuww7UcVzYKSh
MHJXVM4o2s/sz8+JLKBcSHBmcSFf81PmVsFwzeE/N5EhnzlCbPNM9BJRJ1tVMXjX
LvUlADZiE0dvJ/tUfA2UMA4U599FuMMhScb0YT5eRNOyPvIVfdcevfuKmQfUpc4b
27latdcY2nyUidi6TIcw3LXcts+T3PY22H1yQwDL5wVYIWUmStFEiHajj8N7rnbr
GLFRYYmKxI6bZS8M8RVGhc4P0heRl92HOWnP42p/pD7XFHsZKuTyVJBh3/lAfCZc
wQFLjMwgXfYEujUFrfNHxleU4n2Fq/8rXs7dPsb9Y1IiWrqZdK9dyz66NN2fLgAL
vGdsNgsYtQZGhvFDMs3qhJqK1/EvOGATGaQGLHp7VUV91EqdctaKmOuc8mXRCwhM
M3hHxOdSZcU6mTMWbiVSHoTB1zY/lth0yOI7F48/kgqiORVIT6iOTjrVb6VISN3F
LurNClCdu0zDBqsWtxjdiPx3wdG+aEcwGdTN6V1nznuxeOMrVxkxIU3GO/t/mD2T
g+sRYlpY+PtohZF6YCnqE6AgFRUEP2x4jFqMAasmXfKUerFLW3vuGvfJJaHnt3se
DerX1jK4QkVaxHQhwTG77NfKgj6uJRm5pPfbNpuTcIURCvYjXhVWPgJTsR7dqhgP
umI7FgYdOEPXIUyNpYXWADfjPWfefu6106BITFjZNyX6+C3zOZ63tkf/08tzQm+P
PbpLOlljCpHeOdN5pr8ZUmkiy23i1StECBjBbA8VTo4WO6c6pBsAZ1QPh2/AcGAY
GXR2tgbNAL3IH6PPIM8kct0iY9uLi35sWnwDwindBXUKY1UOrwdkf32r3rYJmcoh
HmK9NchWgZJF0XHDu3j2ogEMCB97i3lM5ob1bPRvIAz5B/2H0ChuXK5ecT8vbO4S
fBwLQLyY1+/fXykkhM7vQIKRqin7B6lrA6BglpaeJDgMBYFxBXcXv9E3DMf03SoS
aEBSrX4NH62GWt1PokgXMVs0nRhJxGO8ir3cpJG75f9HZrBMZ8MPZLH2+OghSkCH
k4U8l2PBaNvZ3nWGUehPgEvVs0xXzy0yHK/Md1T5X1aeYOQpl+1SUK4bsFV9lwQo
fU6BL7E4PDuZPZqddcuK+X1Y1gwqkugfG/awsImtFyGxNtyq/zcAaIXsV/9AnXrh
3Nke5eBsP+uxXov01FQWdNBUN8CUI6VjSspi8eaCt1Idj6ImCinMrh+EzQRIoAFk
NhmxXY+Wu4kPrpfXqVPFmjWbdWXX2FrIxGeQlDNS6SjB9kt2qvcF1PTtXI6ImJhl
2KwLBXiB7E6NZWIoqJJJn9j1BRriOEZV88si7LiJZT0ClKI+X04HjnyqjJnCPz1s
s3QIoaak1ZMChFW/2Al0GzUuw5oeGktc897L3xiHInsjaPnJ1DoppwBoqjxl9mt2
odC3RGes5wB6kgkZkbmU1lS7VzmMCcQ2u1J1mIk1p0DDXC8OL6RDBIcYji1tunrt
0fHUrPP0Fjuvnazdop3CAJk7In9f63F2XQt+Td/bPLfX0+4flmLMkts8ThNA+I0z
A51nke2T4O3rmyfI47D/tCbYbDPM+6H5L2cxOWWQy3nwkp5clue3VTgl1RZwjCov
l81f2NGj6BVjwAHOsPCgbewiQD89TyXDHC/M949+NZCvBYAJ8mXvxqMpd3z5NuEI
p7TKuFf4E1eZ3paNRP2EvbiE/xI3tp7ty7yhjgEygvkx09gHQHyBm7srPBbrZLMc
TZyhWjoOeDBXa/q6kXcTgQIaPW+ZrDbJ8DhckGEUihKzi1rztw333H3EhT0pUqtp
tneOJEkEAgUMdfGbbj3sQU9vMCH/2gQeG0LfaMAfOorXK78RhD9hsVXFQOtPyP7C
pD402PC70Hg1zmRg9Ae2Xza3/JG9PwX3AGHDu21cgBKMim6zuMZshgznVWNnCe6o
Nc6e4kDHF/qIOqd7H1fd9HU+Ra6bUk17AKy7BJOj9BTNth78Ul8lF/m45z9Zn9gE
cW82R7vWHmDk1pOPZBzl/UVFVQYMlJz/U7f5Z5r52DyMghxiu+jrft2y5gZbdyfG
04lp8snSV5akJnK+ue+R0FKic83MSqqZSsXn5iMlbNRZtagK8OvuMTkIRkcLciy3
Xnb/0ZOm4oFE2os16WXr00k0WUkEzFD4MHK8fbG4EwW3H7+Qgj6+cqHUF2PV5Mi3
GgzCJi6IL14Qcd1HVDLAro70nhDVR2rF42r+QjXBMAMc0uI7tPjl2LUGEADKJ2h7
CQBV5kVUQD6+8L9c+sTjXQ/O7gvM6EWoXPZe0V9VTxEIDg/WnYTcBgFID3sEvTx3
wKzHe/vTcsxWSUXECNDE205JE2oSmb8qfbI5+XLZnkw/iWrJva3oI0bGtw4fFdC6
aAYYp6Y2qpAJBtV5wMMg7wJUEmJcYaiKJKlHsjNLR8SOgV4HCvmpb7ZtePOdg/Au
KaJI5OGdQxDsJM3uonqypLnDJ+Oypk0pb5QhKWz0jKhU4vlg4Wf29lYplTvdyTEE
X00vcRcJSb3eOe9JzCt+qlGxP0bY7iZDhdEBeq2fExoJRkvzHzzCrzl0E0BSiDhx
EEtX7NcCCNRj9L5hqr0fuy/4SWI4puzguva745USzOA9UZO1jC6IlPfVhOdnW4sq
D1n7bx+ho1zif7ML87UeN25YG8zINcMKyTylhQPO9lilMyhbDISGz1rYkcp2SGaG
mtNK6vkHq3IaKFKzaHP3xkN2xrf0RGLWgfPC2Er7A6xXcN8wlZj2cWAN3KLHqMvI
yv5diCHh5Sx3eijXqdUKUl+py6seGyoakCL3nPvVExdvge/CM8hcQDwj1S6d4D4E
8LevAwz/dn2831qdLIr5kqDuEzEiQdVcLywjCbYe/SAbSqkHa4QoQTSDvTGYdDlO
jOlkzCxC9egt6O2pkcfGZqPXuMxQx7YNBaMcPBwHioNpPI5eCAkpele7SBxtQxYn
EgHLPeDR/m54COztKhUbu4Uus9KPsMWNZzZHYyNNl0oXXW33NBtlVrhWV++LJhzG
r7/DA5/V7RlLZyjU29xXQn54YK9d0pwkA06UKp3YiLj3+ytXVtLDHLiF5OkG/4kW
Z5WwqgYxJvlqPkxd5Ok0JwH+Zlry517W2AK3h8lu3jXf5EopBD0ZzF0kCq/QWC4F
ZxtHv6FotQQnIkwRsf4LIOTd1MbCpRlLp1TKwJlxrz4CLWZbK7LtY0bWI9det1T1
j6h6CqdA1GTUaGap+llt0DIriYsbOWewrgWReKxxCoP2//+p5iiLyhdS2em2WlFU
mDCaNUQ5MLm7sZDhw6zV47BR9g/4uPhK2N93Ap1gfp5gYKEYNm16H50xltbLi40E
VoiI7/SyTRWzkGr+TVQ4b+oNgY1pTwsXFBHFFf7Sj007U6eNmZz+F+pTX6CPOJwz
rSKhV3gqfEWrkXfbP8ZVn7osfpgu3rx9GIs3LqG/LXUbdUCAnYdnstxnJC+Km6TH
QJrisZld0wBxEW9I0ln1YT6tpcW3AZ6G1Qp2YAOg61OFX4HdBzgLBgMVCvqa9gAN
nLPz1y/D/Kbx/9Ys/Mmd6OWFjqkUyVrh0n2gjCmsAOGTYF8MbpIwCUHNpIzWou3r
OdTxtvYccGaKYl2Xov/OxcDdXCN1gGqFkQ7i8YIStVqd9QRqK8o+pXPhOYpNBHDm
+rGhY1KMD1T0EthnkJQIanAFffN20Hw5IwY+xAvb+Pud7jOy7euLgrbpEOGkouwC
h3IGsq58RVP6uopEXfkBIuo7UXSI9KLb55sSz1juBVTZsD07gBH3Ee5wcqqbHGuo
6EB2Axjd/7gqlPW6iVI7F9YZdN7uLenQGRULmIFoCTmCc14rgcS23E0424n/7gDs
J3N9ZbzH5jk72y0XJIT/9+S/twIQuuPi8ZfGrih5CVU1S5PolGnlD3PUcNh+1V1s
OeCmTS9JuEw0QMED+lwZ+4MuAb1xeHv34gNYcfv8a9I5LjcdTTMB2Fnvp2r3nc3Z
YeBIFhkOot2A9vefzcB+A1p/zpA00raCZ0rlK/pNW2GBTZBuVyUQtOZIk6evtjkU
HVpKuNSz8IjqAfJLIqnl82CP/2HbT7TasOX7Bz+PG1cw1oz/JaDy/WcL7jMw/u1h
PvaCj4HUbbVr0K9CoVZLpIeiJS6k/mKBcreks3BxbpQmAnvqiqFJ81L5OOzSk6O+
6v1FFLf7vfPwKqkhz/Tg7SfZeCBWqZ/BmI81krHOxkmIck1NW0pjURYEoEyAQXXS
/8ZEjZcMzbY9FQ5pAsm7qbe+fYM0MnWJe8H1ugJMEMUqX99qTOroJpDgTXmGkjyA
xF4+ifyPKBJT55t2Q51Pp8zE/Bxz6V4iIS6NIxWmabxhCNqW3IVMrFEmEroUItDz
8TpF1h8t3IiXA49OVSdETREiazsM2+0kWCLhw+VGfokXam46P1JNXPx+9VvX2Nit
H6JEBpn7RimbRQ8GARuujiS/GvbXZ6c4PU9X/124AD6bwqyHUlPv6RGF5i7eKwKO
+2l+LgCwCYc35XRdij2/9iM0nrj80EuxzOfHDJUeaC9K2DLxCUN58CZVNLqgmWht
XRxSOYs1/eacKEu9fn47kXIkyukXSwklLKqIlLcJSnxeC3jWO88pVulkUVfFrE28
RiJNR2T199pP00f54Ko8DpAgnTTC0TUYU4Ny4wUy0yjk5iMide5mkOKNGgDoCK56
XdVEsCMhGCW4Hx8xYxHHuLja/NPlkOVQi4sxgo8PzVS750a1oxzchkTUow/eMCnj
Cgj+To73tlGiZ+rYgaZjdhCcwqy3dfIbpwqcOJrC267WS2y/oCosbgL221BJ/dau
glVlZFQcn1OpQYAFj9nzJ8pkHmo8k2girYn4MMsVnEP38LJp+wz1x/ujKdEchruY
l1neylv0AMmQqyWRcd+tcSRi1SLIHMcy6say5/KYPIwRBcKOvsl2aadADdxaBm2S
Su4peW2X/82jIeZaOt4xaM80hhJyT9nBkprGIq6w0o5blcGn+5o84nqPYanqR6lJ
Sexklh5YcjiL2xm3NbLaD5yht2YEAFxAWGJMA8Bn13SNAS7+FYRKy703REScJG1z
NKDJiMbNW1S/RuSv7LVB+GYi0RH2rvMxep/nk68W1h2ivGHuMCwdk7x/gB8eqhoZ
5cMItvXYuRxRtxy6q+Sgh3a7Q7bWad93PvbN3dst+bHbEJfHxaFUezi4H6wyhG6b
z/PbGCWx0MaSxC+MxgPlIbUr0s99gHjW+3dI8YrWn4B3HqKQkVly9ypgZyHPGOp9
EOZSQyKdGpWZgeqwAe8aIhTD/qUNNUS5Ce0cLeEyDUATG5DeJq9Q22GLeysyExjg
AZGdetYOWvieTbpdSgM6xMTPFoyThdG4c7o2SSEzM2spZQRvOKqbAueDze2AJizr
3LTta1ngmLPkFWBsp08B3+96r+Lah1zAUNDW3wvkffpRT74oyWs7V+/cBkeJ7HGu
JJ716nifoinsSkN+tUgJtgLdhFTBXx5iHxqJmRlarDVExfqM7CCaV36wBRSnFMA/
H5G8/gvQdGNFbHRyb/M5ZTM933NprY8CQvJqO+8EAvWIby+zMSX7wbbQE7TTnjnq
Nl/YBjHwxip9QcAp0FtHDFIxFhy3zVGPAn+1EbNlaZWTn2GoRXjJp6fTlEzGpWnA
oaUoLi4WMAk2LKh1W2NOnYF/uU2bVyGbQeNu8E6frYxNcLpmnyg8qtbgp4xcEa9W
3nOnDdTs3lvyhhpV4SsdKoT6WdyXqwtcNdf1lqc7a7hHbX7HW73YboGXA5pG2nsn
UVfrQWzpcM8cA1bUaYr/BM0HlZyD/p5nc517xaKqf27jvu88C1nZhJmt10318e+R
70sf1oj5K/TaDSCuVDFZ3iER3FnuZMeA3xOYczkhwH2zno07bVGhNaPoF/YqUhN6
cCdAWPJ564+jp1xz0ltY5Gll47YeyTr8uk7xBxqYZWRIHE8gqhxGqJHusftUpP19
LRKc/six7T/HxUC0Ks0CgQTn+g7of1Y+/2zjXjUTlq7Mx7hpkPgxscqUkjcvolEr
pVE5hDxftaXPN9YlQn1i9EAzxMx1W002HcWX/r5A2/WM/MuCWeQ/JLf4N9fWHWhL
GbbaB2D0RELKrKZGWVfA/nUvfhm7vJhZuZF9OQPpvhGuXBcL7cApyb2NU9WQg8HV
Qj+9oeVnrqR9JIMpk20DKDDnkHDLzEJzWEqR+47959Skyy1wH2wzqX81UyO2TrLL
/onHTlrV1kPQOgFnJyrk55qx/aHYSKR3zlHNA2NGKgXOgJ23msm/kwszu3c8Fmpq
EAWgSDyUUDErHnb+Ol1dGbyEEEgHlxS+A8CV5tzrmoXNZkQnOHS8JPx3KnqkwY42
aCzU9L8p6uteLpxt5NAvrN+odPb934bjKPTXhe09McGMeBYGUjhPUumfVYGEF9d5
No1aXFMK0NwE7PX/avOp78xxr8uvuf4nqWHNrI33VXJSci76E8kTXXt2DslPeHcR
p6vGBFKHUGegDdEODUgaAxkt0uYdE9FzBYgYqCkg84RAuzMkptiiz8OmXeKp8ndP
o+JiKwRGBGyDVy1CHAE0IQJet5rykEdFrV2ZLOJq6UH+bq7zqqF+FyJuPBfzXJSI
FGV9iFIjGoPGFpOi9tAgzcvSjRuNCmYEp4wpiFCaxWzHmqsq3ol+sswD9LP5xV2K
bc2QPRjkyf3zBPYo62rmiTsMsGvLieJy00SEwqTS2y+DGMDc32adaIbdPnncX7YU
aVS5dHHLv3xlPbDMjpgvRDFnrjZgiNuKT8UHxuy9bwMQZNBkYKt51Lzem+2KVW1v
xOTsen1hp5J0r4E6MSMnt8sSavpv95OgxCwe21G/TbtTuFhUlTY9YK3rNpfDUrK1
j0iDvZi3fCREbUh9iDNk6aYVkfCjSOLN6xAzu2Gdj6U7vj3zoMAg20WXGeQZpvYT
viHRDHX2fMHa0nKH+5j9EK9Iz7gZ6bQPs4WgDY9ehICEr7cmu7IxLy5/w5NT14vx
8FKj/+XTnGBlFz0Ze+PWgjt/sn0c+dmuArRoM8DDWz4ZaaYCnW+XtfzsEIIAqz3a
6aMBfubSGOSaroUQ5K7sxbYzMHMXGEdz78+cuye2hq0IKoEq7Y+cmAhJ1uLS0/y1
yUPaMW9mHp6WqO+5bEMTaqZofpOKtcsf3ZHFsHkzANnkYpYUT8fBu6N0oZ36uSJY
OFjFXQQvxFDz+FJFd6m/POtxzfGD0KSR02P2S5fqFIaSgNGHmXk0B2vpRgZHXyEQ
g2EHh1G1fUM6yxlWTMpQNjuCKIhtCZa0w2EDfm5a1odYlxXtXtaATMoftMP8GW7W
dlfe4JPvdqjXY0NIbi/zKzpfM4aTg062NaF9QwgD5pDb+xZZu406aVpa0elmK88B
xRlpDA5hVPng2XL4HMwCr9CdJiEtiWWs0chHrufUJp6dEFTGAcpgvNmVkkjChqhx
P5QUUfv3eVyiKeatzO8m4pIreMAxKnjJXgFiN2a5PYOOMJxzAo8JkY+r9f2Xutka
1bGguI8S2EBsBKu0UhJFdSwKhXmcleKEp6Y76/oRyvwyLoLiIA6C+BUJbhBtYjZA
ytF8KXo/qymiU6TtEa+1hDllTZ9bkNmez5/mZBx1lUZTKU1ShXoFswO7WgYT6ogs
sH6iyWtNJw4ph/SEdvlTyjzD1t5ZiYmNXZE/q56WNRXG4KKfWgVs92wVZFsgSyvc
HUF0tPJ9wrdk3mC8+vHq4e/jriDIsagILdhMx6dbvonDjykBkjSarGH2bFwfbhhZ
Bhhz84m6Y3nPGNFVmztN/JAOC4G3Idx9IZRWcqTH+2BaQCwfRgfpVkuMHx6z5FR9
MvXQ7q16IB9jgnBoOl5jQcoEnUGwoHj49bBw0r5Ujs5uTAUYbleoYE6jBFN9CPzm
vzq93aM4HPjPzGg+D215srl1fgGWsI9zALxLCf2G7RzBdrKWtKZReYEAfeeMUL7V
IiwFCxDtd7bzfPWl0dAbcyjhwXSTN5+Nt5mvuKBobZjdJMfCJ5mqqWArNf/PcrlA
RDD7JAXDCBJ7Spo2WFnOaRfcsFmmkWPWVJ2N+L78bCWPyRSjqG+2z6n7oGJHCJtJ
fDw4Y7FM9njrg1ns4BfNrI6qfWbQx6QdA0ZxXXlvVwIw4kYp3zu5LBVQ0uW8B5x/
0hndrQD5RWa6aVCwbcuLB/AUyCkDNSOIqo0R64JMxmyI/rsUDNtaLVrXivp86pAK
l7Ues5msuaMAPfFcVKokPISLYCq0dntYvu1tCHYJTeNQEXnmzi+9CfNB3RynrMOe
PFcekvRIluWdKzUqOVrGGkGYh8wAWoCtVBqCNJ+Ajs6wbS7hqPmA2GJw/qLvMV1y
K5lps61zIJo3TTLKvNxc3zpYNqOtWXzLMzEdPDi+eZOXvpZP23zHaU2zsHI5zNzj
VV0y1F90xyGK6KZM7/xtgYlYPCIQT8xsaqrUAWhUtpRsBXO7J4o5ADuhxGqYR5NC
U/yGOBNBCayJDe6E7SuEfje4TjtOYog3WL76ckRHVBBu5lzH0c5AWRrE19CPW9DS
cGK3lPf3mMNdeKuVsqsIekxvaY0CHnUMCCq09yoWPkX5FwEQ+JVWAHCRtgyn9jfT
5FMIjXkzgrgr4K1p/vGrpr8UHTxJBjaW4b7WGNFp69Y8d2ZVEItfVFR1zmOWuFch
6P7mfGKYLguFBhGnmblbTI+J1TnBjB5SdWWJTMyRHmlSOJvLx4nLKRjjEWNovyWt
PJVGCrCKJnrN1ele93EAtxkS8KGT0TXgCWXDPyAouLDxi4GK8VGHXvHEM/WdBB/1
7bS2YNHYRHrZZ4g1AEX+x6IZW3MrmHiBtX+wWNPhxSMANvFSVxPOXJbSLHrnxd8P
szwvk54Lg+OoNI0iBZ/6nQUMne5c6oA/b5CZ5VA8DPbGbTYEwwZD4LchmRqR8S/m
A31yU0jYGgaOnsviJcMnQBP+AylN0sukc/7M9jBkSbNNt+TOUuhHxxdFd6PeQLxT
aN7DBGhWkZNetpqW36s1p/Ibr/pTV/RTrDAl4n4UUmWbqkSjh1XZ+vJARIUqhjLB
bNVCXAtXB087uCqBAkavnsB+9VoJzU3Jg/qBdHTuWpeKJpWp42QCUd6xUGJlLthB
lOJDAYeqjG/EtsbcpKFC5aN/9Vs1RIrlA9t/C6C1AJTdsi9MAgB8FQgXbb7su3Ha
AIdQDBMxZiNwLXtO3tZUurINZw0471ZDIcasSZ3hBh0mT1lI112rKVQ7AyHlWaZR
frBz9+Cc0DWxLlChq6+9LIuhm5hZfsVu41+i4T9y4uCUr2CxofU+FcOwcn6bPMa3
jbFD6rumdH88EsZyIolKI+bVteMnFcRhJNuiWq2BuBr2DD4phvGjmem94sAyO1ab
jizp/xMKJw7Gge2hUPnvo4v8zHe7jUsQBkcR52tvuJpE+KHwx3PMU/a81PeQAlrJ
8HFHHWIv/QRZnsS7yPKCIl0lnVEhrpQGe9JuzRe14HJqFYbRmdVP2hG1E652aKh1
jegpqOhPM6lEFNkKItxwhhC3qp76xZyrUTtAmKNEn+JL2eaBQvD7Jbgkyo3yukT5
ZIxcu7BONknrSXUfRxMxZSCVonFAdGJk6CFMnxJi3QkuLAzL9z+zZMKDXHKVzn3N
I5ee6Jupit0xqyCOoyoFvSuqgphNlvj0qwyhIkUNHMJyoMZB5yujw30ufMAHPmm3
qefuYana9kv/RegQhWiJgLBO5YECcIqWpu1fOfnUXVsiq2YMcg113ko8PqDJpW2s
eMzlf05iMPogP2YygQTKl0ZWsJZtOGulcpQikQ1dnjj+caBDD0h6n4/FH4X+HU4M
P/WABT9rW7848ZapUv6IeRPsyBkBUUweVrX3veKvcPqL4pBQBy8fxz7NC+aMiHGk
KuGronfCp+8sNHkqTFrRh/w+naxPqO8blTzPZux1HJA7Pf/qailrjV3XWUn0KD0N
d7TePgCDgm6g49BJAj3rH98tHfkF3Hl22oKhBpryhLHl+xxH5RKM6bqBUcFx7Jy6
TI4l6cp6T8jXr/pc7v8l/IMJvwY7WUxuLTGNde6T65OLp5UAe0N8nsYyPLK5tDGu
rhy9BBcLlgqV01vf2xjI5XDF6xTp64/1E2aoORufct5BPvrT7BvG7cUWJSts7Ntb
WdwGKsX3L2Irf/rz5/2y9/y+0E96S5x0e7ObI1dmBeMob4PfYr3MS5Dt7dfIzqcE
f0YmGIJKBy1Zlya0KloLMS+Y6qZlkgSNie4Q6t9Vmx++QKVWnbJKGtAQh1hwai9O
TO992C32m8k4tYBfMpzBijUg+GHwh8FNUfeuo6WImtOs5ICcfGLzR23wu/wrWylo
mYStXjliZLUa2Q3VCQMy33JSMCFfilJvk+vXld1J9joTvq2gg5lpYdcqmEV4bsLw
YSuX+w4GSmLrL0s6d1bDiuo/HT9v2hgnea5hjIVQB3YAdQv2/f3G0r/3ly1EVeih
UCXZUSEVuGCIeJsVRfEQ2XR3riSLWgRUkw3t2/xzvLlK4rOTVTACux3aoJjMK4RY
SAJQ+9brV/xQJQG9R26IqFIr0UkrmIqfUaCFPkxneoURkqXF/sADtxPTjIsO0uwp
q4m5HhTrailfFQgHFc4JkfEP1t1W6qKOZaiXgEH/HaL3wZTzhpThw57zdxwfLQj5
zFU7zhT0qdY9faYOCTXGOknhH3/pQg72esWytcMUxKQFIxi6GSH8SGV09eWgflbN
LG1wxNZrwaWtAFN4iZuHO1Ikof5P1HWbUPxSbC41fWv/xhtKRB8Tnlldom8eIBtV
ieQyNGdOJLq1cAaLm8GnItpqJk0q6gIo9qW+u4niC843mMvgPMjxpRO0axIorNi9
67Kt4ih6+DTI7qq+JLmG6TDmwMR9YToea8cekTxTFgKpi+a2D0217wpNOCIpKZvM
MQkVY/2403K8x6Zwh515S9RPTFaMXPQgWz/Giiw7Sd05kau1nWIywVObwAcSQRgS
WpTdjoRVXVcLTHIjsovS9jBrSzEzU1anxdAIfqFTHtkSGQVOgyWedy08nPUSBX/g
545mVrDra2+513tVJWF1OXtyMSavDgrSCMOiA4obOUYq7I4g26IMlCmNPFQcuV8H
BFxi/FJ2p/LCePtgVKoDCw8AoNbli+aiMMqK6Y6r/ccuuj2jVba9q7eYrtthF4i/
LGox7H7wOUT3SuQOTox3OutV6rtoC6BUbXgKpt0q3AQUurDCVI0HLcgill7kbXWm
UxmxjEabHqPNmbmUes0aGgItExbA5Cx4PtTO8ckSJLHMUHPzGoc4zZziFCngE6gj
wuV2E8TDyOzV1fTIQBjVCyq6PHcpvbMjs8jrF79LpmJV3UQQvYWPFrvTz22236Id
Df+kFr1mD1Rx7PxvsjeNxiUxxE01eieRVtxURsjq/iylw0QJYAETIKaSPPeoBGkN
KdvHNPx3/Eg9RaYXrn/bRsociEEsOp5hiqAV4IheNOMUqA954JF1hNmjAVMi/HQk
hJ244Fb5Haug3lYOOdUm47OdKpWPPVRWvjAciCxujqeE+an0V53wCDtXjW94sdzg
mAEETYIziDggMNbkDaewNN+U7bZ3vQysJZyVG9FzaQOO+z4VELhicGVyIyFFibdt
4REQa901YNF4MuNyBJTGncmEgLG5NMfGnNlnxbpy7Ho1YTez0on5/q1by58pwTAH
4MQkvueRbkkHoGuXiE8ZSZ4AUpz68YZpxCPMQrK7ms48c40gCpkzkkTfawmCohyR
VtMlAQxL+zmyDzpi4oKhiDtHbgntUOAMpo9j3mUAnM53Jqmui/9bRT0q5ZNCzukS
heCBrJFVxUVlEGODhPVVv85LtLP+p/53haJf5hrcsnrVS3uE3Fcsb8YDROXJjyEv
QsryynNE1CNDFkCcesKJN4dbEg83DLq6NLbRKG6vFz6JkpoU+xOk+pEb5InTnZQx
rbQWjpaDK03X+GNz/supjvq695XU3OCw8CN7jEu2O6ztks9yHeCJlhgTCUeEt3CS
uf3oR3RGKG3IMJ9Y6+CbPxsPRq+HbTGzOJg7wlVDYgkLVMP/j1N2B8wvlRZ+P6cA
NPRic+cVP9vWabJH+BE+Bk84Tx/DzHN+r94K7wu7Vw4dltGqf4uwvO/+tmY1PGuz
v/i5SkIlXPvaID28tXzBtW2gcrtWM5L5BDQJ2CLWF+YyegHMA1GnKm5igmp/GcbE
IWTdYkTXnHTYULHkQVOvjAK2muljw+vMZTc/TiG4Ula0itMurHImHteEbwRUJZTC
NXCWpqrtQqBqKpqhdJeSoalkuFQdgu6SOd3LgBXZ8UJz0JQenlUpuBICmhpJL9RO
z7toV+pNnDSFHzy8QvCqt2iOadnXtcYG3544DNs6e4zVRpriCnpK26F7rv8hQvsE
neolUUVFl1Xchql2G6dDsgwMYDgAkYyUJ0hn5InrwaDIDY0eka6P3s6Xg/FmYffs
MbmEmtew5Cs5XJ/YknxPF7DGe51GWDE1mGnUCRz2Ro2p4i776cPTrxDb8V2oM7C2
BrEQVLgcQ1EqSXUI8w7Xx88frvctdHy2u0b5L3UpEBX0GTbQXeYRC84rJVJbQfiH
OYnNIZw0lO3kusYg8+6pSxyYKKMOIODa48bg3udjHkSP3O/s3V+xQzgqGMtw5PBg
hxedAN5fE40Y6Iwd/IwFXU21Nj0nWSpYevVHaJc+jd851irNp/4zeMU1Q819fPbe
xzko21QTtI42b8IC/iauqhTwJzx+nlgr7LCi4vasaXQxmdMd+TsB28qIeQrms/t4
RQttLgXFcuf+kIKKi+qJzq0HsE/xW4P3Gy96jN8dh/O+OmQbuCuHXxK9M5V3B+zH
uHuXE8S8YjKuwzNAGDniklFf2HM97dW1aQzTa1Eujv3SuVQbW7GTC21baJLob8iF
YCPHtNB5fsVR0tu/+L5v60cYBGRFXlAbbFl8pNNmz+sG7wD+tgeT3pk2dhRr5nD5
2CegqCRSAkJzBRKxsj+u9ELabVFw2JjiF2FDxj8vTambqOQRcOJ1p6VHxz1zQOgJ
1IWPSfXMU4/8sCOcIuoBOCCJps/c6sUZ+UsGJWeixQCGC+2ivaiRPPap9/tNrqLT
32PukJxWmhPSsJEfuURyCNfISLGxdHl81z1CP7KvmbxZrFlzRUHoLsL5+fghYW6M
x44wutNEnNXFlWD9igNw3dlJzZEnlhtSmxg1LhhhCW56dpSz49XwXbSr49TazIbW
3OuobjqQwC81bWPpBCCroVhDuzfAC7Az0CNpp9qjVHfLJRkdcI3dbS1cbZUVu8//
+LPALRiPqZcErohObtGjEkAIMzk7ScVuG6fGNyk6S8okezAU1lsMTSDPPbok2mX/
pOZQXbr2Nmkl+JUffIoQgUbZhJlgxPhNnm5qnVYaHRmKvw/uSp4paoJK5loEB2B/
aXkANMjrWRYtZ+aqjcX7VrtD1am8V0evYK/RIqYWzTK1sSH5gb1Zt4slpJWO5nlv
dnRruoOpTtfRaSGXv02ap76DRrYzjZHKUmLzi1WIxe4NyJGoQnyq2JQIjWpQGr9U
yLtBq8J1Y059sLa/gOwNCLmzFSaIPMfH9Sx1NyooJfJR3XGtaN4raAx6ykWjSnJf
gCl9bn2YLLjmCQwxSfDECAOfQGVYhNrmZGeyLWjfga53uAj0QK5pcFiFFwGVF2/e
T4PlhDrds4dbIWvMq4L6fpxfvtTwADipK2Fycj0Vfb4yu4NkmlZ11vitmYVK2/Mj
ab+wcbqX9KMyHtYC0ODnokWfxRqnDhhkzmNEzZtcxeVkzfM3OvRKg+or0FLq8R72
2Ik4zeVgZrIAMRosStDE/+HjOJ1UcCYb864arCPl/gHksUQi0ViIF2FetUF9f761
VH/cnNGNqV4fCd7oeuo9TDBtNuFblJb1iYxcfwP9nnXx91qE8btd5Jq6r7P67G/f
x5UHprIHTG9/dWmo76r8zr0gR5v+qx133D5fuxQL2rt332IWtMgNfiScblRJ4OeS
wiWt7vWOriq0aDaHGm5Qv2EOlI6+ljE1vdjacVwKAAp1ZLXzWi9AS7EYQ8y4fW3E
2MWJFino/11eg5h21uoDp9rjHA3xTBWiTyGMk1VUsFObDx/QiGRQwXFdiRH60t2q
qoAv4Cscdiu/pbRm08nsiXuV2qzMLiLhxufdU+aay65G/aT+HEQxlF7XM0/DLDoS
TnsZ2OyMEFORN0+BFWHh9zQEPV9/xXB2rD6uIfDpptSFTzAoOoUxUKAFmcyhzVj3
tMijh/iFDbpesuwJaYP14A+2Hw9IU0bebdLtihbCIg87ua7Dw8da06YPs7yUD2tA
UDH8RLgwcGCJM/RpwknbUwnayrhABg12OZyKZMX2nPLpHy75WA5IrqoyhdwDZaZh
kTTWDRr4AIUrDwLhwT6P/Ttt2WasM02xQNk8Z4zkCVclefAkLEfVbCIsksM9hWyt
4Z2dK6CSzwvLmBPltkJNITEeKSZ+GvBKSsPw7DP/NOiuh41nMAStI2iPBacASTV+
AzlvD01w2YY9ohvxmmy4t6azRQJbCyCSE3IJJbyfexqP/H+bl4JdA4UAmJcwILeb
wIg56GTqCvrd+wPmrqIBToB6wJsCGNAm+A1J9Rb7Gg5mNGJ5Qd/Vu9yoT95FNBvz
0tl8ALe6hQeh8q7+Q9A+g1rYefVca6qO7hx2cVqN6wZC8Kxll6ailh6IyvXP3iBu
1WelR7k6c6smqEqMT8BekB8J1Jn228cD49MYaIDfORlMTFmOtTjYo5Nua8eJtSg4
rFq74QOqbezboUABhwU1zzX4kChIwG9CCc8VR1Pw09VgqNBfFtnTuFPQW3A0eyCz
Uh8KBqzD0QDxZyyWYTJHjk8GjC9olGdG9OJOOljXjPRlG4LMdKGqAOP8iz0VJk3a
AoVOLvhWrqqZop9bHKvqk6MUovvsC8tDSKF5ibX1+9FYbDjpL5eCih7kJXyC0/Ii
tBdVm10NjiiIhKku0WHeyhWWEcCs0H1Zp/9C74aReKiMx7B7xj2rheUlC9Pb1Bl7
W/BXk1DPNTdkTmVdrORRe0i216NlL51aBqqakkJtQSzjU6rMIQtNHjM8VFiDrILS
8H6MJosdNzGPFPHrWT2Q9TBKjj1EwQvZ0RLUdWtzt+alBLonhvtYhKa1CExvLkTk
oXMWSAk8El52c/TOh76+W5fArl05qyAoRjeLj4kfyLvRaVBcG2w4Ay06oONU7vAZ
hmzFuK5Ysf4Am1sKe37fala4HrllBmy0c33WqfxYaK8LiaNjPDd6asfjy+gmd5Wu
VFvpyNXwM2+SUq5kwLcgLmh0Jkt29IE/cKssexSGMfXQ936zyMO+VFsrgXcN1FLi
BCrhJSyCNuVuptehpyBr3zFGieZggMCfus0TJebz/iAIvjITNyR6IlT5waT7tF4P
Vkit/Dzf4HMqhuWf6uBSkR3xO3TAjQNrj6POL6G5nFqkSW9A9nXejOEyN0Aoy/v1
tdmhis3HimsDb9aGTfkPpOfl5VkMFkY87TMJAn/JIiTC+dXMbpt7syXh49sL8eIb
ULQ7IkHW/s+lv0Cms4hUs/qWeQR6ktbIfyk2KuGDqqFq/SEwDjbylNKSeNgVbh1M
ZNUu15vEuPStSkUZJQ+nbffEFVpOK8lYbxF1Szh35zL4ScygpXsMZ18xhez6P1Gw
ZRfwRQCK9rSSoCyQOYQk+leJzH5rfSiVkkjwpTS0FcD3YuMJNMtzEwlpcYRcQZvm
lA74zo3lZWijaMQF/IsZGa6ly4ZCrTlFXPTT6M0VpPR1G0Aa+M3ETRxqMUWFU7/m
QzGBN5xQ6NB7h/9+lOVwOYpoGGi1JEeus/28Ga5R6HfrEV3+F6WPOraGpG2RKGUD
cypgXf0pRoOpgByRu7WesZKWyqMtuOU3NwvEeSkm6SS4xIzoD8J+jFKF0Fh1G1jg
ffoO0ReyArx8K0BPQklK/KL8meMomGSQRQSv2QKkvBgQf2EagjA396zbRNUoNXyE
BmrU2ytgv8m1fhzClcKskecZqtqAEZSw5tHn86DMyMXelN53ObvRzXHlc5t+K3Tl
r9TMInisvz7bMy4da/dxnhgHiY2nf0MZFjku4jLWHu6NNlDtChqtrJ5Kpo2VNKSH
EFk59wURgfcCEpPXK8vctPvtXq/1IEeBKVxJngAthzBIqo4lorAiQW2DMgS+De7q
mHLn653CxHF7N0bqDH9kR77Kd+8yt71zk6N7yWPWMBbMxQmD2+cvNbMHa7HLkJWz
s+hPdTTiN7qA1WtIWhXpAjnRwpwNjmvxzfNPX3Jwk92Dcd+3dgcZQvn4f+QjMwEl
tDhyIwDSrCbTlbngxlKuk2fv9yCmo6VgW6k87NOyw8Fv5lvNE8498WEa8060fAwv
lCy8z68nQo5mqfbOl4ImT6fr5nAgqosol7P65Sr80Y66E2Yo/weqATcLNMzUGRtj
t7zxkGZv98uA+kekiHmJRJFN6/EChnE+sFY9ViGFqyLL6NRrKcQ59jFRKclp7+jQ
JZ1i72YQneOezCihNL42q+qep/N+6RM389pAcGdBZds2b1meurd7WoeHvZKKNCz1
I/07fepYrxnCyqBr7Z4WW8uZtwWZn707ny0s3Rg/pKnUptkTyrCdLxfnRmBlavXP
oFbPa48ZNDoU8oBrseE1m9hMVaPR0s0xo7DVdh6z7gQUWymoQlTR1pCqHC+Nn8UM
zfgq7D+iZDryTAij6sKdoOiF08/bw+DilXi6kCGnfITWooP0+LGTL994JypHxlU3
wMeUcV3L06DfHXkW0iJQdaoPn5ZhDURFn6WHg9hujfj9AqwlsM4v0KYfRiWiSvZn
tOO8yKvVcKB4mJ0xSpjA4NDbH+7U8Gkz/D2iA+adA1IAS7qK1CsyCNVRLwpmGjIQ
TnLvaIvpYVnalql7K5AyrfHcWsEIAG33hvexVXHgNaPfVdDxEHzI55BekX/L2Wel
wewDgiaNZUHyQdTIwqOgukKswfuC9a7hZj5VF0D1/qHvFU6Cik3WbOsOZSy0uFSZ
anGWGsnJqxi8J1WyAb32T9rLjkKLAK7/HCYIddV0msv6NBJ+xXo2yye3cjhYAtl3
odIM0ayXohwXj3jZv9Oiqdl8NT09VAOXTm8Mfm+pRCJ6Akl5247OskMteKxccnSK
EdEhYIeogvqiVX1piZ+Y6HPP1ZrUcl67Igzj54PTvhci9mqWF00C7GU0xXCJZ4sw
TJwjXZd1zUeOwlFj4kxyrxHanbsO0/reQPA/QOGjuJnNvgU9JdzQL98otUh1bxaW
rFIrI+GXLTqqkXfPqJgo6UXJZwM3+sd2wxD0VpZ98uqmhCaAxNnxq9VzgqFrLC9z
kBPxw+N6X6BG5norvKiOCcPeUpOZ6k1keShnNCUvHn9254lKmhxxzEzSXlDGtfJx
Kpppls5vKc/Ot6f+klWU/YIreRDmK9cNczRlXuRfY7uLVoLEm0tI+VRcqyRK0pYT
M5LGeynNW4mYUCECvoM4gF2+MDtuAKvyVYwE76IxCH78Z/v1CC2UX6+VKuyoH8IV
d6h3PkMEcXvxVfOWx5LOBxXUk0G1L6Z0gWocEeqf13oZ+Kq6d89RzsxubpflE4pR
Z/uJ2UUEJWuXGwTPge6HEKHvG/eg63ruolEeDEYS9ESiv90GSuxtZdILNbSlGByU
HeXvKYN5SCOuiCjT73mVKZIME86reCl1+DguQFNhPN0dH5wafcfrv/npiA2htT3c
hWGOuOQmHlsvhviIMWFQBl9kJy27A34y9idp029qKMvL9IOCPd0PHPOijsjA6mnW
C7c4yjPmc+RR+OPLnC1aYZfTbwH0Dnlc4H63FmfxMRVdmS6aOao20/5oosWRen5T
1MPBtUdwln79ZZr/8+djmpx7EJOpZmH9I6wWmVjZD1c9O9FadQAevLLFwXwlOme7
zDtyZXv8fyBdFBQHt0Mx4sFZikVf0zudgWU+PpIU9yHub5R4PwrE/UJsatiYVa8W
Kybd9XBYUzjLdSIUHmvsgvRyDk2HQi0deasJGsy1+Km4I9nRMKX4Suupv4cIAr1L
ufQao8Xecqn7LsSG5Z/JofdvU0YeZ2Af4w45rbDKfbOumK65w1T02+P9ppaj/1PV
25DevaYI9biHT30T91Kgde5ZlAXEUfmXOTBfgW7euzCgPB+Z8kl6K3gNGqyo1kl8
SWTCvUPJIZjEAK1daqz7L5+nA2XSM1gJiv7ZrvYXril1h8vT4bp8f9PZpahT9CqP
NPGT0Qp5PwBZaI5GLDTVp/EqqJELTBDV7rQsDB4Jth8UdMywogRe4T80VDXcMY80
L4HMdhn09PNNj4ALXiwfmSF3piuAo9DQ8Z8K523kczK5/QhUGREzHy5VhKqrdK/v
Ppc/7iYoajrbaXwttvYynsDBRxEJr40XbpuhLA9o56VoNGIwa09okuEriWRas3Wf
o+w24YHkfoDQd1JYfUKDOz2UONNpDalzlrOvkN3hNKskJFt1PEWvcNONDzPhC2Gq
Buj8xjeb7tSpj8SljOcdBWla5kQgbW1Uz7USt3PyQjpYHnAlYlyNnCMRJGGzWoMN
gjdzSKKxaaM2i5b7T6MdP+rK/g2Q+lRMKerXfNJeHtP6YlSbtOaxogl9iMJbzuxv
GaUDYiogu1EpR9dnNVlSCewRs/D/yZHKYw2qEmuLhZCKGANKH+7lWIqdirfXdJXF
ExnyKfq3XPfunK9z67r5HetuBuizsX2L3aywLCJ9+mEg1Yn06s7s/mrHYKZYh1s2
NQsrCB9EXPmWZFVSnun5NAycvZHOX2OE3HgvQpUTEwYsckQwEp7FUxi36ssPGB1N
elqZhuWchmzMnp8MTfNfGluqQHoZ+IxsvbUjsnumSFepofDlVaUwjeUibP9+WWVz
0RfDg+UM9WjXgVNURzYt0Iy5wgKkMHx7ila/mRRj8s8bhKrih9JiEv4pOpZ9GUa6
lapovFs2B4F9G/IL68zL4Q0yaBZDazL2uPIM6NP/7I/haqK5d0ja/uN2CPwf2gMu
CFppqLqcC4XUwVtM28cd+4WfNR+QgyGWTZ+5MHUO4PLKXDiqmLzDkgqt69f8Lmpl
Dc5J1P2MU6/tbySMarTQ4EWAiULuuavYSnEmXxVz3Eb5OTnk9FjU9wdsUcHl3jlL
WJ1B0BzlUh83KOjsBav/oqnXOZNadEqgo1rt0bH++2JHXohXawLMYdeYmNCPDqQT
23PmAu5Z57OdxAOfCs7x50x5qF0D8LFHDdL9SV5Q72Zgk4JqW8mibtHMYQpXcwGR
v0Die15pe9WxX2cNU9kmWDN+nFW7XeFFoTFv1PKHAiyOShQkZ5bcaUbR7lbmxs+O
cGxhlyG/VAWrlnVlPjP9hWkGguG8ND2jlwWocq/Q2cBUdwXR/5mz30I/z+FpQ9i6
eHkV9aAASOArGILMUEWqjjyV5pcmX/TcL0N8RTZGpE3YiHLTWkLSjOy9VwAqCXPR
a/QtWS1ZsZNGk6MRcU2L2IYZ0eLJvFKV9n3BjrqVLVqAGrUGoAMHG9QxHLaU9iVT
/wGCvM3sPZpaueZrjYGNaT3S1nlHxxqDU7IORLglCH2eVL9puINYrbzFpGXMgRKY
KCwVXjBjPRrKZyK9CirPFIbZZaVVVes9o2pWDp1VGgcqxvNaSj80ySomTQRbL5Ab
9MVNhog+nWNW7hy+EutALkbdvraogX7cgc/QA3lXdB+SUWFoLUsTYxFXEv/Rcb3M
vNQvGqFSc+qS160BrXtE4N+vJMWpj2BCGpnWGH5X+ESqcWswhdeswhhrdinOOX/w
OzoJyWjTKcPWVpQiidoJIwhxSGW8GXRtsA4SDnNZbQIfdHv7JZ+DvursEyQ3LlFU
o8QmNZQWpG4fQHQ6cx8YbNBivOB33BcLHHFyYWQ428vo3UKvDyLN/Y4X9ZIhDBHX
f3XdAKxVWw6rpu9mbtNKEQcTz/EAr9geCF278hplIXsYaQLPq1peCzdkr73gC/T8
drEF/oDIFwqf3ySCx1M6WwXqAzgqGqSRI95br6KNIdRfTq87ZHRuyKHR41emS4jI
jXT5q5s7sdr5xfyM2oR6fzuq4t1QAfCiavYa6LVNB/M1yRA/1z8k32kA2wrYW3m7
F8k66CExVCMbBDNm18fLOvGDmH9w2vr3EG4Gkc5pajOQFHckbTBefo6JH//mrVUb
uvSfHHqJiIGNx643PHLE/Yfeahs2IWxGTYEcVXECYB2sucVN2PqQTpKDS7eVhbyU
ILL8iF9e3llRQ6OqnkUQ1Q+mfMf2/2ACGWoCqIOQBF9W9hFSyAOF7d/2tXHVKlYo
lBBfHghohsw93CzxdE2oyDrt2yk46aj2ysiPiJvLGQV6GAehbyzLiWNR7QCqdE/D
Ml6mIz1eAUHj8lNOH8VcmoRtNKdltT/fjYoYivbZL9N1xz6LyUkkDnl7bL4VwHLP
7jjaDfDkJNu0ShwE2eP78fJCz/J4BhhmJmqu4mbZRWDK8ktN/g7t9lbP6jGqgmvA
L/3MLdCUKrWnwlh6nmP0zHTlbeNmwGq1dsUYmVHzPCFg3ePmpgTsPvaFSKELiXtv
Y2iwKt/LaRNB+mpa4tPjXFG5FgmQWhNwihBjUNQBFZWXyUzs5pWIGS62qe7WzHUf
3TQ5PohuQYSmUmFeI3yNSlhIfRGARP9zP4R9IFTgKq2DB+NZUG1Soaa9JHxnERRG
34p0v9cvCX6X4l9fcwgrsbemKQospi2yisdMIkKYpvyw0aq6/Qwinyq7hx8ljllL
Dp/qMMtOlpziFYyS7EwDi4x2BFcW5Fojw/aqqlegl2eccXQ4oRK5cFaX/O5xXrSX
C2wBNpORHruCi1utgyizdWJrSb1dBrmkkFiSs1rC4/V0RoZCQwOTxiM6IPTmnvbH
K8Tn8dQyov188TM/OCQCn02OLx7Nz0L19mlZSlBuhLKtQ+L05SptC8UbgHkBDPJf
JpHAyxveac5HcKzLRwJ8dD+B5iTjuLg/dLL8lkanpUwbkT/IJ9DQ9FS7jtICUx+h
Z2Df/HSkvrmoUqFYnOerXcfmRXoK6io+ftB2aeIkLlzahVqagbEqPw/BH21Plkll
3DNe6Lm7zKiKbCJgUFMeiWocfpLwi+0a1878ZTXqUUR+FFxFoK4eEps5vm8BfyGT
rxGVM5zQGq5L9DbauP7oK+HD7xi0mfOwnd+QtW/IZTk94QfvTcJ27Z1Eb+jyDscD
NzteUsDm3at8EExp93V8jmKDCFsonBKJ3WZoIISVn+jQJ18nAKnm5OSui1CU4idp
rjSilF1oSY02NXkBgcxlck7hEL/o1dmugvE4XWaSehxyZmpwekZwY2cpyeg3seaw
xLAUxbN9tZYt5oY039Zo65Ds1w+bH8CkD7T39MfqaVBD5toCOc28PAuwCpyggU0Z
6Xf46Dkw90ib25m7ECsjOyhkogMmOYCDGI7N6BnAncawRHjP8WKxSLBaDNp+UMSL
kDLa428MGQ5dBw6Pm5JYQ31Kri9AHwgOOUKjSG5ftTeaTgU746elgWYlMVyYZDJb
HlEq7eAyF8GNZ0YUAPCu5Sq6EJl0nwKEoahLGW08WsWtJmDV0m06qqOAECmSIrAO
HUiS25IzXDXiR6oy4agEc6KSquakSx2oA+w6dJOfSbs10YND3t1aVN0pYlwGsmUc
PsE8FsPU6rq64DbbQZUXialwiBPR7L7eJ9hYMejGMJ26IXPmoIjTcvAWz5/rFvR6
JdvboSRMJ8uIEGOTog38EqhbdtZ13P5K43D+lTdGMag3VhddsXi5TfVybeYMwJKE
ifXuHM3DWRnzDCCe+76tD7uf+zZfPi9eLydbP9nWehfqey3x+070IgpELLDkl62C
VcGGOU7GVZlE/kSLLXHcpLc5cmQaQp0yWksG78zAKDynyaiDcd5gbT15zm5H/s1r
bZDH1WIyKXjJoD2DviIeCnvvC0PB2kXaS+aWrQ2dAingkxfjvT8ALjosG4ir1C01
VyNQqueM/oMljDCUJlUkmn1EPUFjfV8LiwYwW9PNoxFOnY6ZTiGkBW1kW+c4+9oC
Vx6flIB2FT0VDudIXIkiCusRZK4IEmSLJFZFzZLXO9CxS8QsuQ7nbU3qeGV7U23n
MxCR/6wWDHE0BN/UoeWJZSQCB/O4bE/6dYLhBYmPHK4jf+WUVxbiEdFFK++mMhmy
+cEvoZSG8M6Nq8xWDsdX/2/rIXHp0zvovZGvcx4BsxMkZSizLL2gTVHTMYavhANQ
3m4l+YzkYqNw/yMpnYN/UdWjc++IXdYweXHEfWYU0MhDjklFN1djxzD4ElUCTTHn
eiKYC4dV/f5bOmA8iz4okZg9sGLzQavEXI91AFpww7GjpBuUTaztWuuXzRWsGfOE
AD51M0JOgjZHrr3EdM20OiudvIyFlG7hiKooBB3BzZJGLDamUTlLEKNveOug+36R
0OtQzcnjs4ge6/czY42hIe2iL4vC8oL9XYeKBBghu27TG6vVcmDuCDGSxrANxz95
8Tb8kHg1adPeCIC32kImYrB29Mvf+MSbrK1eD2VBJY6z3ntos62Mfrrx6zgvTJpO
ePsHTX4Jfr7cHLWjzciEgOZ4Ha6Wc1Mey38A/c3v+/SQk6xMG5T4mCpHfsgHGoyj
4pvptEXFsx/3dycoywQKPY8Xxn0TjuyJmOluKqIoTF9sxfdEozYdYereQmuh+qvf
66jaLOZ+yQmFgl2CJTRt8bI9XdTNf9YLvqG2NuozQJBOi0VNILNK0smPhsI2q7om
yMq7j62nEcPiSh/RP/CcGdzfYEMDcEHH9qe7GGHW00SB0VnKv+OEabEhTIGonmsu
bm98Ko4AywkDdjz3ceTLvDwfhgTWYwGvRPNH9CS58RXRkDy8RIWpbWy9n+Bd5wKx
RPoL3gaoaX0g7AuokxQxAcjo30uniT5LhUhvO6y4WjvvxZfMVhGP9/Ly6+hZo8jB
5uWNYN+e5Tk3EzNsJZ9syhRJt5Ynla8jfyFbzb75ZVYk1/ctbIqqihB3gN3G8lqW
adYP+9OxKhvY2fsEqJd7oscrpW94Xf3AkchRKUpsVtvZgywAucXPrhEJObo9tkAM
s1rhsTq+Cg14LT4TMmKnaX89y7FB5O3P7o8PZnHhwWQ6t4Yv22GQBP5zXdOJupMH
+O08MXjBL8VV+BI5AbP53dyRZ6VUmoLvqXLreljuoUuqxiQGZXgzEg/urlr2wab9
A6reQyA67wsTWHTf0Xp4qgwUaC034GKQODMIU4dNVsSHwt69rbm8CkSd0UO5Y2RP
er3Jh8a9DEXvqcgBGAw8qLja8sagfGU90KSbvnS6zCIATZB0SP3uS86RNb75lTtC
3q3MTZBh+MK1Be+fxn3R4f+BUkIJcWZx1F/v1m0MgdMmQjM89Q2EiIvYqvfU/NKg
srqsfz6VmqdZ+37zbc0S8f49tySWLqlfat2Mztl4zOD8zfpEgWB9RzsmoYRcFuAf
AemN6XQHB2rrkmz8XpMdVxbYZI5rO6AITRXY0KidiLhvdM8d6UZEp/ElICCR/Mz/
3s79LOZC8M+mYytFqDd0Q3TfMqIO0/Gr2PiiwrQWOIMjL+HBqXqg0CLhUhwSoU6g
GzwYzHzQouL7iFTHpuT2ssOvRdJSG++eSO5NTiirCtu4TUOxhaXsWHfrR+2DWxCH
q0ImcOIlJ7KrWjfs07H4oelspql2Gfj9uheMKUkVI6lTI5tIvlZ9F16F4VyoiDt1
sKmEilXmtirtPJnvIy7g2F/0XWZMn//OU3KyDN2i2zliLl+eljAL1JzDU+ujOqsD
CjDSQkePCoeW1lliuxGq5pFMqeUb0lou9R8ZubK5IJMxnQb8Oh7Nam/cWf/9Y7TD
MLBpJxFtonVmEPY3qPR2j5gIUD21Xa0q3cEMz56gv8sOUMRNG6krRvmhApzXdkZ5
3y9Kn7c6jcrQP5u4pkz52fbtmnzrG6ojVnSbJTxapUUBbobWp6hJZSeX/MQFMFUw
wzfF+Wf09d2iAqOxy+hvsjNX6mp64nv8WdZv4sIcgG8+7gC8WwyQ/Yt7wTY5BnbY
q2tjs8JEIIcHBW90l/PJWxxLiQKRVrD8vOVW6LJaiBLbSOMXyzN7jQovDlj/5wwp
fVhXpPpfykmj3A9QUinQCocHcQqz/EMH51jEZX4NLrTu+Css7Y9wRmo1T9VYYikS
5czf97JqvnhzYBdStgdt2Jwb4YMZHj1vtEOq5mVqSAkWHhwPd20xdFF7Wx4NqqGi
fR/NqSmPOzdI01cNd0VCy94Y3EM4rCbpEVRwDesbCF4XNql8ekNfeGCWukD9Lvz8
C2296/p2f7o7gyXQRzE2R/85gMUo7qxp8s/s7YOUi/5QRvZfz4yH6pfDk+JOh8+B
ANYe1pJpOIJn5ndPYU145xbkr7xgbo2gzgNiXVbdmrq4NmBAZRipopPn52lXiH2F
ect6+oSMPisFMfqNk+B/OpPtKVP+18jCvbChmuhdjzzM+3xd4id3bsHvZmz06TfK
3ICWB2EMOze1+4Aq2G5ejtVu0g132waXy0KMenifeAzwQwsuANDYHK+yb9FsPYra
L2/U446RG4vFZnhWoLVJA7qrxklvPz/7LeYNMd2E78nnIzNdi8mI5fe50LA9vEb4
bmU6b9ZjI5qXpya4yLFOoLgd9Fefaref7gSGz+3Zdrte7wuurom3dw0RY238Zdmg
B7g0iv15bZI5lqUU1uX4dPTOltMipF2/i8GqZvSLvG6FIXwUCDvGnZgUGaUn5woy
eJMGqYOqaUk2+uZQoeswAto68qeH0Tei/2WDhlakxzY1BIDqhBSlbopL/cSj3A2y
/PL7h9Ij5LlyByQl5rgrKcDJ8xuwrNO7h2joLyRHbOZGaFeI26Xy85yRgnbbM3tw
6YEleEmVwpZI6laPW4pmIxaK/huNgi27IPL43zb855FPf4B+kJeuiGfSLblXAUei
JswMG9T+yum7QW2eyIaFh6WrXBAdA0At2dztglFOQabws9JNbs6QNaJw+3GXpaSD
31jpYX7YlipuOW6w0FDCPr3YJf5y2shY4KZWhEuVhXn9CL1UWwggew5SvyPdmuJX
qTtI7IcNHmYsViSbuX/1dVAxGYVvyvx6gXxpZH5pctlLfaUI+lEPq8m1OkZW4pER
FkjaK1tM1E3lGnF6PE7AKQaLGMg2MRcHvSsRnrODtvb8gNhIa7GSEMOHz3nN5FLe
AKhWs7XCH/Rj3Dj4r30fOQi+ybljSpOQm8Nrko/GwvNQU3GgOnvlXU728ViXSomq
Gx1ebD77NfAS0azyR6D+Xng+ZdrmJsPA6l6G7kTvLP6LJCtRkFzSwFmY41O/V6aF
zrX4MecSDoahUjX+IBIDl/hCp5TWOFxnyQdwvrD1JA5H54V+8XDR+hXE0F8qAjOE
osYYWhDzbppfLVYTNdoArpDdcmepFX5opsa+GbYkbnJahHDVup0S0DQLHsZSPCBM
Os4VrB3SPQrSdscHsJyd7p5a+BwnSnMQ7l96f/dZyh7BrOlcYxySqqgOd+ay86qs
cWZjgeHww74i1P9e+BAMQlQgd9EIvkxge+glBcOi6lcnoT+vXYhUrSowXr2ffA+d
IMtvtaTthh2Xco58icr+7g/77MS6xSz1eGBbjDIeA/0oNkhx1g7WvB7ChP5ps6b1
deiBZ4LRmNRVycUfIKqMOqcLYdl8/lXMVEA4rMFPVxymaMAzObwYrhX5rnRPZBJY
row1Qb5t7Cyv4UqAktTGh8wEmrD3xaWDbTJF/cN6nxT4IZX9aNoKxJ+4zoW9U2cw
iO5yIfn9SeGKtxTDbJcONqaoDQCDNs1HoHcIbInh30yhlX53eOQm1n/xLErsF1N2
L1RxDS5CK8braZGPoarxFCudpdTVLc6FwI/5CrO30CwGlM2iKNcnNvk3cjJbsSYE
h7veycPNzzbyX4c7cUjDNjtQwKMmh5ZI5AdPXYJvDxWCsHeHHCbLttGxnVnKz8c2
TU2IpnohgxumUfGRJEC0TG93NkpYNYpIxkc5d6yLBBihGo67uZeI2siRfHb0cYdr
NjgT/WaPpBBKcZBX/dyNTICYp/U7vYQFmZ7kZLFY2vXumop4AMA3KvQW6fFh4UJY
d8vGbzCVS+eC2XA80ONtUHrx8huA2A6wMt2LMmVLsm4Ypy26ZJBMeOKfj9eswFOH
haZVFd0Fyze7K7yViWBLKiaiihnweB9J5xsfREi3bQ8b9EGqFArJYII9eSsPFB2L
r7lZghNkQ4uJT/ZCodCb5ranI3aBi6D6EE9lOF/QwW4srgWdNMVkUm32Ou+1gcWq
4uSz1o5rg1CnWxbMm05PxLkbMhBlUrvT0jQRsYDtfPM/XN3ZPnUjBucsSpy9wpme
Z1OtQ4AMR0E9LNl7OtbL2NhaEc7U8YJ5kVrlmQWMS3Q/MELasXmKzoY4RlhPlaLw
bcJ304Z9QVjx8+wL4UIAhlyIpdVrN+8q++lsKg6HJkGpti7FHGkLhdB5z5cnug6h
1hOKvSlnwPkXbUedBZYBRI6a5LZlzXLQbo4iIdvMSAuc8z9QA21S63A2+y25NrqE
m11RIcnF62/PnsG0EEkJ7tIMq7vXvAdsWFEmGHeNV2CpEAlwDDgHB5eHcH3EB398
onvuwndQJS0PCmanr4656ZLggTQI4Lxma9ZpNznBchTHyyWp2TBr32xWDZlwWhk0
NymMEio3UtDLd9MaiOfFow8vgiJEgjQeDbx5AFHY9tPL4MCQvWursgVmv1BBZCG/
uxusIyU9/CUnssWV6mtiVQFIKYwCMA35yXLPtNIdSMIvnCysvNcUziKCNYiVkB0X
gadZMHptk/+WWvzYBmEoqoT8Oar4o82wBgDnT2MjMpzwL5Yinen/YR8yXgEGY3Lz
iNR2kOGZK2R87r8XxjKmsswhYGxMZsDUE6Md/QwDRGE3T8RTMZacPDRs66uIUGKw
Y4Fb0s1rTSCErjvc7qv8UjAwe0kUf4tRgROeCsVJ5ZunIq5irVqx4iXIen5I67Kj
4UUef5DEp/RSnXO+mIkNpXxWeIev7nr2rnA/Df5BXzchkBfaq+fBW92crsc8M89f
KrYUCgy5Xjw8cvIwIJ+yRR+5aUuEG6of4s4Q3Vy6DtonwJtBxRfpOKqKHt3idd+B
TH91YvD/ofYdjyi9LN/i8NkgwDi86Fode3GQ5QZr0ioIskqUL0lH05x2SU9044Uv
oxIWQIjAxvi1PC1J2mUTjjCDaiwqXRPmddMUiQiXBk6EAxhEul/Dv62OeT9ckhwS
VGUPrDp+wlMe/HXijZdg42TRt9kESzICU7VR7sE1iQJwc8DA+sS6dRNGtche4F4e
YLY9GA7dGD6oQo6x0ijyCvebNGR1JnOTq8JaeXxh8KMA8BdXivYW/OcE7qtgi/Dy
4S7aEf2glvRdUcGnJ+lQ+dHAJKg2Zjn/7inhrVrfmWYcWn+bjsyybh27bAZVIJI2
rCgIgNknFoHnmOFig7RAbmJmDAyFLv1r5R5iNRdyJz6zv5d5H1RXw7uL+2SKQm6y
+QtAEMGh8wtnxiZ2YKtBkDojuElUr0zcn4S4YxLKFFQ4ncIoA95hdgu/8AboHIHG
dSkSzJ6Ay5NHFz6qHnPiNiRnFre2YZLOpfkFtivxDWIpo/LyzP52b8c8Hv/ziuD0
nxgHDiCh3d+V0UV/1hKxBUDn/mtZEIwtQ0NLrIXvfVrNqWJTt1LKByyQsBVpmZGZ
rhgGYRdeWw0vyTs7PNsSM8/MX1Pfuqb5KBgtv3EnOTkH1/LLvf7EdX8zOCmVDPjk
eEFKddr9KOenbkDSmRWz0LgK+kMrJA8oD3JafJYcxfKdwvkUR1hvDB4Y/x2EfOjY
h/k8j7gJ6qoblr7qWcPgPV+NCKJN8awjrErMqj7aifshPuSuSqE7uVunfjgHt7nm
yFWDQFq8u1+WzCHKX42uXD4Q6GODc0lqYvwVxrncspI6I+k+/DF19RlauNigSvKV
/PUQA3yv2XeGthYY/OaCQvrpx9GFb4OzpBYifLkysfqUxKzHbl4hXsp6b295iSj8
47ahoMCea0ZLljE/tqBI8/Rdf828mqXpGYXzz0zjajZ3R7TzuexyICmbUGTGZG++
Y/vYUPlfgChyYdKfu1ls13DyLYdkGOP4pnclaGNkhRoKC2fbzUAoJdTx6PdvB0hD
YGNHaNHQdPHjNQCQhhfyawBJZO3OjBX0+G/SjliCLQ0FlIFtAXwwTRgFPWbAE3IK
GDLWLBy/phgxGIYNv0qEyARTtOu5zk4H5POd8/WuxKBF8DYXG+JFDwXLZmiWI7dS
znf20X4QE1sbvfEfYoQyDot3a3qwPrAE3NlDlk2Q8Kf4Wxk8NhxZKm6VasA9gBC7
MYd/30IP6HynLAtLlP6EwFMhRSpLidS0vNTOmGas3tCe2WcF8BVTkr8fbzujLIYo
RAbvs1JrB7sZ5OgXSNfpIfPzzHL+l3juPSrEkGUtw7VfKRoCOC2tZOprKMtFyvpz
lThPUmk5U64Xn8rxkDyPhkq5jgo0sYfFaAGOelJ8rbZItkP6fcNgD3HODQYvI79y
uAJ5DMczfs/u+IMfWZp392A04rhaVFfNEZt2Kf8yURKmNADowu8hU8dLHH/c/yZw
lkNSaqXjEVZZf+XMinGXwkRY4ULn4fYbjeT7igW2fGjx/X0ga31KAI83gJVJbVMp
Vvosv3m98YzoY9EnuclQ5p9NU8+yW7v3pIZC5wNzreemLH0E1769pmqlqIBsBDPV
t973up4ndbjFq90VHoEV2kPdHknHh0Jj/CQkJTrl62uKW/zVEVJyIFJwogWzJUC4
itXPafeyrI5JaJ6pTbUFX+EuFGk9t5NQbB7N7TRD4fIUlP6O2UawezaCRDtvsxej
x7gUlLw2TfQAlMcd8akWdRh2YlAHRXIyEwdy7DrONafPWbRtGyY1Ib0Ygi2bW4tK
gawFV3fo651QfkXvs1G33LXe2Oe2aOC6Kua6IFYp3NaJ6521cVWGmLeRZPlDhr/x
bBvTxgVrO4YJjWFN62xs1aYqFPoUgUzccZL0WLvfKEkHimUjxXUBzyHTkKcvBSwL
OgWvSS3zGpQt8iWLDlIyF0zVuvXxDB6zHgak+IvSvwI3CwJd8+GdmahZfKTCRTNo
OHgWHH8dhQuX1Foryb8VXcIsbs3MiYDhSlUtuiw0didaFbRo5tqFWLEOevdloOIs
gIfDvXKrU4kmbloCquRVhn6L0iku7On+qA5zd+jwMSrCG3zRDj2JsYW7kI2g3ds5
qUEPnInx7qkzpISdEF0RxS8zkBZxEljXlOBqq6NE+dyQSbcwG3E2ihtqHqIoIpZQ
wiHxvFi2WubdRG+K9va+vgXcUmqZkrZQkvTrVNGYrmsIar8PqTCHons1c6KazaPo
fbTmVdneNWuOF7GAHsYP2A6d9pyTjTA7ZsJpq8gBHFzPJnAWlKH2dN5cCwLVQ9qF
zTbCeyMnk0RjJ87z9HozFc8Y86kJxVnJk8WL91NX7vy0W3YQYGvc10mzuuD9Ojve
WZ/rEvl2deUbBxEkgFJtnKdMElDGDDhPShPBMDAXOCMUQldFvCfKt3KV3Kr3W1z/
CHPcU7zNgeYU8GTSmvCE+wcgIK3MQaQrqoRxc526STYl9ULwoO+Kg2lHhJaO1vMK
qycQZCj3AzKOk8gO2Mkebb26LG2P1Z1Bk84vCTc49vTdQ3drGp71+uLDYRMMVyRL
Tld2AludTeBKv2753Ay2IslF5v5NQ/ov6lDx/mdBxB5jdJocqxUYhTKRrZM0EpaJ
84F9NsibhdF5PtTwQYENh5PA24XmPjH19cCc1vO09GbIori7BGigCqkPR/IS6r2R
sdnaP4DLX9iDNILAksQ8Kyq4/kSYIjoINqHeslSl9nImLSFwUwedXJP5pRrECHXd
TnnY8/VCuFbOJSP2siuCpk54EdMLx1wj+YYtJl8hMVUQNEmN54nItykCMwd6dOfy
vODpgLDdf4YIdop7YyTQgzHwLpbh23v7zpO0xfdQvLARez4uYQN6HuuKrnlzrZCi
kRAA00U9QBQiQPpsKeJhmbxdFj+BSSzpPtbHcUV22G3RcnGvb0yqkchO3zjOSpO4
wwIdpycjeJDVpjG8n9IYBMC3d+LC/0ddhAp8J0xw/0HF+Bp0Jiy4p6eYNdRBDwyL
NQ6I2gm2OLsD/oF68lI9aDDqcBAX7kxqV09qNhQM19/dS+HEIYlyKnPU/nVZTHyD
pjroR5ZGS2mokHqpuXE1Byi+GlFDJFEUp3SkFco0qH9R0Ldd92YHrjtjvUCLB2o1
1TiVpdA7U1o4fe7EbxP27EwvU1PVdzRkug16NXD6hngKwB+NscRLqL/HbfXbbKiI
vsQ2QL0CVBY8QLoIS67Wekw8GdmftxQNVWt0H2AzOA/L38+WMxw4eJW97S8ErpcK
KOC3Hy4/JfHSOnyl2djMBU0lFI5zX9i/8nSVHCjvc4kqzRuIuE4XWoXFb6o3uyS6
Kd0MF0jKc1alKme2ZD+KAsMUjkgItSioxT7LVHGegISbL1dU2YG7aNLtvqC1y9m0
xc63NakvPGUqf8Q4Aj4/38M2VH2F/QCHwiiMm9+TvGhLbxqH94nlb1kVec0qMVIn
xoJdiNB/4Wblj3nSzWr4nY7JvciBldHD7FPxGehTznUejqp/fSAHZFRBVYD+lnv6
dHJytEju4KxrmTE1g5j3TNYThB9j2LZ3DnJQ4lBr1zEC00AThgjN+hhXUkn0NYPA
T0EbQ75GwVVKqmBgqIgDKgpfsvuBXBi5r3NlUTkxifaMixD8MewT77R4nYPVfN+6
1bjBehaLuMyNs02CtcMi4aNBxcLjZ/NkSZHx8+KjQoyNjFAK7WeTor7qgcYdljSL
b7rWrHdgaslkKXu0IVG7wafWdgvVf+FbVSpT0XgHWKItaaIE/kJkuaU2ruXIw6Ay
D1NWl7VScGXKyuwDEQearh/mHCWoIEGCdTQ/sexn4VTVBVw5vh8TWhK9q6xj62UQ
Q/fvVSvs/GHhBY9IaHzOe+rQXzL0BKKYbGrKj/rIrsBk8XTsHhs24HN86WQY9JSd
HZqwUN6wQtbN0wiB4xFm8GT4JYLCj11+xyBsEZW3Xh6SPbviIM0AeiVQWTLgJS5C
jdZ9s9ioYLrWulQXeD5jrIA5lUu/p//c4Cp3LtaYwx5GzEFWDkbO0HpKNlPBDYhU
j5gV+nTH+y1kQgQ8yj6tijSN1i8lacoWpxsyf9X715vTWBRV3llHnf4Cu71DiIcN
9/XdEIVs3Frv9pZ4NeWjo3loa8J4JsilnWzf6CinEZhN6Q4sNCDBCbhf+i+7+Gn5
A4FYc7UU455gU6jMVltIm9WhF9gcXO907bPDJzWDV5cGcT8kL1isMddTy87Wt8Vd
VbJMEUn2BWwP0oOpDpB7JaawmPFrxd/1iTH4ADxRXZJ+PXP8v/YAWXJqXkoQ+pCV
TCU8A9ADIr99g617ODM86bm9hEx549epCOsZXwaQdrDG0xxNQjzegzQF1auUxCbT
1u+i+TvCOryaHOSceD5TbLH1kPdcjXXjozS32A/nzV5lhHtc+PZw7gcejvRmgg+v
7hCObU4sTfL1bZ4D5RRA7wYV0AYbS13SXdLkvtc4yuqBZpBV5rL6cvqj6MdiPSkv
brw7JjKz2ZQ79UOtE37ew8ryAqXgL/Yh6iXrolkyt039aYB0P5IIgjMVU1w6BXmj
FGgNUuSwX8qPVErXCyxGitW6X0l/YyCDO8XUTaBzqHsOsKRa0HmH3zRr6IbF03NF
mivzkf7SDEzbn2FhlHxisP2j2djhjXhHu4V36mIcdAS+VODWeJ/Kuc8D6qhLN/Ob
hds0e0Pr2wH28wwYxyhg/ZrroZgASa1DjuwjU//qQ/SbeAlT23JKrc7jizb7x+Ll
NwE0sHA0HLxJkYi3x0hOWmQeCwLYobn118yvZ+Z0bNdHbrNTSD/MBq65+yFme5xi
zh0gQNVonEM8FdUJ25x9G7iKCBq+qkBTIUrDxgQxQml0xa/Tpqj7YaBelkH0u9fL
MIWPWiWanykrovqQlXv6/LwjnHjoTY0GwFjjEYHBq9f/PmDnju5SLunV/35FJkJz
cvUv4mRDRsop4LT+S4fh6Z1Ug+LTRBl5bD1bW8XOUBFIC/uZJcLwdnKJZnCGxM4/
qGcEfJkVTEwhHhkn4ZbBUMVjGiiODTPzqpDzhCm4MqlnmKKx8pUzzNuecMIG0RWJ
xE36CkzNdrQmSbRsToDaahUflgiAXNksD1cj92PLBPyyBogupduVD+a0tA7/5DLF
0GJy/yvgEkjZMnBYpODDYT/Z47B81gXzZaT8cPeJKlme1aO1K+XBHnXbWrPyNtQZ
FxeFvbsMONPP3G9MJ6mNi1hjqtPQsgGUbWQnpq4Mxfrv6lvz9WNTeGss2yWsQ+fz
Oxn+mtFusrAPVogz96ygcKRqkM3QtB3/nvX/gSC8Xb82iEtO2vOaC2iZqpIm432p
I6pOJUlV1uuZcH8v4hhZetFv7WPsjUlcsbbkmevvyC7btrbuo8JFFFVCmP9l+J/a
BystAPmyr/Esd9PLaFz5Squdr/JWKKtDD6dojvnO4NxcHbZTh/ju3HXrZE8u0bsX
2N9E/EaFVB4HCM5jNI50eNlt2Q/GX+cMiRt6taSGlHrUcCpc6IriCaw736mEZ8w0
3uDhdXY5pT1f8bEqKV4cscfnhO4SDh73SyM/nNTOL9vpz+SRnrQylm8mOVyw8RW0
gxz30Ku/obetDBEt3Jzvz7LDcZMP5yxl4vcMzZUEGENASlAtmZzlv9YNl7rwgylc
yqEZIWvsnLJuWaxadSGe3nq9F7VO2mBQtbezycKXYNk/H/sA0rXRaw8lFUJ41Jao
cjqJiC/QtT1PLciuANyYKPLwZCCK22br92D4aOYjU+YsOkYKNX/1Pw7uXGPd9pk3
QWnxlyQ8lfaqFauiPK0E1k86IOJCxg3Fv3DFdRI41OqbCopP6bxUn0GFHpJQj82q
c+xf6/q1acXNGiMNkQ3KNPxyiTUT5y5x6czTGMyC12/H0tWnVX1xlxKnGNziUesw
lNuBxv9ESw/aprnmWfuDmXRS6CBARd5HPYMnngmb3hfh8yspltA4qUK7U6Y/6Mzh
ChNUvZdZ2qy8VmyZuTOZF08011mpatkPuN6UBDerYyJo2gM/pI+bHjTxrmAR1Zzr
pQOxsdWgUZSY7cna6+v9M/v51hnpTQWsXfBdE809cIMBI60NUUVRUhiPY5zC4Xzd
IzAdVIvqDFVq26JB8rYtXYMyzOfVJBsL+9twt2k5cTK3KoC5X8iIxQQJUdtfzRSj
pRNVUk5Ew2ftEERjhjWu9/Tgd8E4+CXR6yAi/mMkM6V+gL/F0TQ0i272YOw7qNZH
xC9SffdMxX5qzX0zKPPrMkPd1Z8j9V3e1EaMkiK6QFTbQFucnplL4imnv1yUJmuh
shdbA6XnsAC8jXIsJqdo5pPhO+k+MBJsafqb7Wg1sC9jYiMrzIJef7QFixVwE3Bw
z47SilZ+XqaeGdlv/iANGYN+odfWb22JFnhm3MVk+43Rn4N4hmQNi5N2xk3YX50J
D8hwqo2uWqrq3fE7I5j2NPErOs3COzVnQRkOCOkhQSmI0XPe7Chc+ubrHsssm9J/
/2tMGHBqawvJju10YR1s9QTBXDvPfLLyCTAuLqYIEpqVRykTeDep5jthQaPA3/Tu
1TzF9przmFEmjLhS931QafRma+t6S/XiAs+klhnespS85th45Al6iilvwHzZOL2o
hW4XUeRjBb4wzSsiGPSCWPlaBnAPOyBXscTfRM61vpwqKAurDPpwGQI3PvOlcUCi
4hzMX+WjpeB9a8KkQTQu6++dahRASxzYjBjVCTFbKZDtWWWDMKzy6rssWtyxwTRx
N95xccRq7kAab4aNBLGpmiEgTf6myNSq2kfBEoxmBgv7s0blJ4GCTddASAsW8k7j
HIHQk3vhxS7KSj8u8TGSbMxbxZVtXGeSglvg23x/YAhd5AzIQ3tNTox6dMM9KHXA
s1hkXnV1cSodKtRztZLsNpAZkVKvOpY3gc0iNCTsONqjk729MM+3IoBVjj+rgxlG
NO2sAS3exjqGDMpZmBGJRgBTGlcEwmHaGjttxKymKnu+VJkOagqJZnTEEsZlCqhv
4nM1ojePoKqnJ652ZkQPYA1z4Sjz1xqg2YgbDn81vpTI+Z0kDTKm7QDm+ou5p3xj
dCksPbiyS45KCW2A079jvWZasHMslGinEnhAraxMUiPm3PG+yRzaDCwKuP2YAOHn
Y7mNBNi/wpA27WRQO+XZxCcwAQ+3aIDx2fznNtnSJfkkM+on0EtwmbvZrjwgi/zr
1Rls8u7UWR4uSHj00z2qMQCHnPeW+Z8lJM1DUaRejyBE3hREvo2nVV3sXhNhclqQ
Qi05m4tMQSSWVUZbXAHBVGe10QGOtdskWSIIcThZDwQlAiSRZHZHI/8YItLD6/h/
lpuPpfm1yGv2uuKra0lmRX5J6fqOAAmAy8m9xbUgw2o6K5uCtwvo6BYKmle6x7Rh
bd6wywJnWyYzE7rftR3yEd0tnGxI4Ka4hpEEZ3I6UuEC7+v4LFUFRFfYTBPlEGlU
sb101VpoXbHme17b/uJekqOOcQysXImB7AfZEFxNZo8LqXCKdXYW+1cyykpLhDF4
PU9ekJpueDkGEMc4A8qdHebMFczGiBO8ojwlnr6XzcGgvCurk34Iz+0GQ6hFnw2J
MuL3W89D16cTPZ0aaLqUiiXP/03+TS9kRLfzpIdt7nphMzDXLypG5Ec6vXKPGvt8
tbMuu0KdPMzElPEJQKlWEKfmDQt8dRq4EnQT3SP/838KjxBeWcO8g6uwjxCGxOT5
Qs9znwwNWAIBDr7mSlRq+jRizdJikIvuaTnrgDyFGMiVn+mNG9XXFjVgRz6IZRSH
GHxvza3fGpXW1jOZgXXahestg6kYsmmSPloNksgjBWhptIO3T01uvwDPjIKKj9Un
+JcIShWPw3ucv5jVmvZ+k8QMsw5WPmfKNl0JcKXi5vlkUlxoylyvXUdhJYHw35E7
DXjchPbQ8jnkJi636jOTjytM4+ayINppsQRvFV6fOpr1HRYaZqfemDXFL0srFIlv
zhahadxOWBw9RjpQcjN0Xie9qXEV9ftVzXH2JfcBNSRo6JaAsjFqA1vdOc1tGAG3
gKo9yACbpvOmHp5GvAEvTyhIHBH90k/klQ7ojtgkP6F05Gb1+cLm4ZBVSg9VBnM3
moNx2OXt76wQNVtsQ7Xt31kvqZSnScvTKWwMhOpK77hrIF5zUMLwIwK9yaf4cCOM
rIz6qUPnIHgJpH9dDQjiT/O8HzrlnD7nZ23wRaRAsw4zL3EAbtuRra0qFhTTulxR
0pCmpRDy30YdOtu1SBVRhtax2SNmP1y51x1NriMr0ljJH0nhZIFyTN/VEyzEyOT3
AqSHEGNxRwkBiZAh1FCoJURg0d7oJ5wmUL1TKPZvyYzfsJyZq87IoymQPVc0jLLZ
xJC+NS2bU+MBh35xe4tdRyZHD5x5Zel9Ou3zSdLib7xVJqhblfm/RVMzi1nv13u9
0u6GxXN1pNLPcekAjkQD8p/7T7JsnDvpFrzwJtQlsprXcfk/gQkzFF4DZYJfATUb
jxBluR/zUufv/6L7F3Cg3ogyH3ByZe5PZJI7lhLgozxdJfOBlemSefA+Q/t4/h1U
okMCKHqPizJKuKi6bIuLPYiEuY1FJce9eLYAcHvaJ03zbXq/CM3DzQssdiiJL2zp
egiFkaoyl+UNRMMQLnwqm5vPyrOSl8G51sdx915KrAMWJctLNCDPaT06ITw1b7T2
+Dz9HbowvsFsfq4cglb4q4yPeyzLzSiLGLN6DNfJiUcHD19MDGBet8zXlMIV6RyQ
gmEIi/5XYao/b1wMU3G1SqzxN8aJNlcSUwmaQYxBH+5FB9L4zDLdXmUPNNVjuvwU
fOlfvk0igyNUwQGjR4GmfbgGkCNehfFGNJNBqkNqdfuhK6mBi+YnqeRA1/LzIXcP
Htz4SYhjJ4FedxWXYXUlIwE9pYVk+M6zX6HkAuHk/+UgqgKO7OzePPJ6rpC8U6FX
l3MpechIY9yrbzz2kDvxiq3fqQd9yDMzS9r4la4PBLIDTCMca/YW6jrvhcEwY4FZ
4UfuvVPOb7uaL9nnAwAr+dNcuXS/Xld8lqGzI59tXSegJRGoxapNJTsFW3Fk2BfU
KGLy9CQ6eGvjWsPhAg+Nxkq7k1cLkTDXvWkb+6JkjBHxWG1yaKwMPkS/w2ejoqXZ
wz0CT2z4iTQA2AA3FQGn2jXxv0th56Eyw8ZyWvuIQ/FtCu0aBcO2KZN2fkAzENHY
zl4JtVo0RlSMaZcrhqWrqUDsHRnRcavyn0Rg9sytHUnmHRgVOYw47F3v68tV8kDM
LoVro9ag5V+gmN3/gr3TGNZKNF3YqXMAV50vPEeE3LXJqkfPivCWIVFs6r0MLG5D
QgomB4xFLbtcAEcfskB0/BpSxJpVZYQYBakmnB2vL/6BtdpfjVbxKnjZk3NAjtD8
WGNZfg5bTW5z/QcO7TCodmRZH050sIeoa1BNaBjkUfiV8iToIxPWYIqHvORWR0tL
0Une6KCOV/+BxWuByAaWNlMypuLfvJhZPAFxfWcuVkNVdnbt0nkJmrEgbQPGe+d0
EjbwdPsQQ0Icq44eLixwSLSNSYMesoGVyzOsnXlPqesFMeXYDYCmyS3XlAOHifqv
5VnSGUtGTFhiK8LjFclITIlmoV5NXW4hMo9tNFUjDt6GUgjmpMNnedALMDlJSPPs
Kd3btlPV7NVn2SaRQcf5sZSGyEGPP2mf+/Db/S4KIIDHsTOwtIzXayjRrzqETnFE
zIIYQXhnFEJJXPKaoDjbg0sSJdh3rq6Wv5bbf/oB4zzinGEHTbPxisEUkvof5JRQ
25cuwId76HYTOMyAKIKvo6d4GT2wvwR2pW1gCpPjBG2L+UWtRGQt56RalmW0xWVx
S50J+Be+GQqWxGEh5N6MsmmBFtYTwZJQRigsm+4hBlO0tdQIkd9kEwKsDZFJo1xf
LCo0ftjyZZNn+mr+5/mi7RdbMRaxOLHqproMNoEoUJlw4//EgDenG4NjLXNOLUT9
G/FmM/E869e8l48AY3acaTGTjmR696paBEW8uwcZCE2PxH4KI0bKcs6MM6r2uLRe
hvXgLnPJ2NTCO780wU8ZtMHPlKb1tjnP2/Xn7I4K6+JPhP5Rl11QatLUWu573ebs
5/fAqwJWXs/jGZCCFNj7gxNrTy39jLh+ZiOxLS1pG453bCtbWv2QG7QJhGqIzTCJ
RJPEl2VKdj3lvaxFg7MaoDk+jpWMfv37BhrU1Jqs6cfs0b7OcLpk0tKJZRVlFDtg
84pvTiKtn3tQpqjY2K04zPlFi///1X/Ux8BeqHHQpY+6oUGDnHAySGG3TS1Ymb0O
rK7f1/CsngzEsWFYpgWb9QFs6L0Fj271DLswTWRJtXW3rFcU6FSXjei/Wflp0jE+
uSGJ6M8cYUBmkBTWg4AiUxhocibzgAdMyT4lfL82LQY6TH7twJzR8J0qbJScS0IT
wHj7e3mPSjSmU4YWaJXdp/QvttAJkTKkZ0/jrO/HSvkUcsAMev1BcD0zuoQC/zEU
ZDNZp9qtkGjbK1RvBMB2RQQzbYUpoj3erhxpuaVs0YC+izoMhQKvhnng70bCRsCN
VGXL1dJxSR32RM+6W4tAtRNwflRjhp6FDaeo/NNIxRfiy8CLdU0kQL1JN2rGswPm
di1WGuhsowS+k1p5eFvKwJVKkxsB6lNLYZnDD7l6aL5fKC065EIWlnIVXJvFKJnc
nT/tRCvuOWcbG4D6buktal3YuEQ4Lbzj88lmCCOr+PbQcZHzxF3sYnLnRVdroeUQ
CXa+X4nR5yRktrT7OzrTdDES8TuXHBl50K9TsUeAnzRjFoKdlnorHVEiqj125rdL
eBxD+BaOVOYY96QmP2SJF0v1IoF6rj2yxrj2OzXhntlsEGEwOmF/g3lhBOR9HGDL
B2IKnIIfVP+AUT7Emf19nh6uJlB61OHhFLdK5RtrzCfHgZ0o3o+n4KuTK7ujjgmP
BPkzXa1NJ5Hn/sGxXRenAfPaAY6+1+z2ZCtSf8y/c3t1F7fNK4Q8T0azsfy7UzAx
1c/M+qoodcLA3KR8sc07qatQI2NUM4Bx/13/zgarRYAajG0MmwL6fkwyIIVCk+3U
SiTvEVsWlPmbRnr+Oig0n4ADi6pMYw39tpe6Eu584ZN9gWqWunUZl4/FVlhF/ARA
Iq3Dp/kP0JprGO9ROIeaLXl8yuw3CqGHTXwwFZFhkrOCxD3NuyR9ZzP6lyYLDp+0
I/sOy75zlUS/SDK0ysMcEuqT2+e3+n4hnlPlwQmrGW9oOtIeFmXXzikcM/Et2Vey
0b2p40ZA+cZSfxEpe0P4PbnO7bEmm2pYqfh8qKaGBg+G9hrUJ0pdvi0wUlWWlXpH
88AK6B1xB7dPWMfBGhOCrVwoPd/pi5B/MrFZcEGhoPb+2n1D1I/OV3lpIWveRwRb
5pxCpN2baGVR7M6ER7QK5Xa78AaZKOjH4Bi/FGsNbJMOaXcI4jcbGdZByHUIoPbe
aGpTHjs3K6FTYHgDqftkw5um2biJbejwiNHeAFS5ECYJSnHDFHklsWpeX1xxKNVu
j0+drMsVdlFwZh9rPWkFDwFx+IE+vBCvMZcbALiMRmqA+NJ/BIgI3460vhI2Lxn/
qgsSLPCro4ssBx5y/VHUYSjLhwd3+/5ch1Ov47shRng/CvOmIKDPc3XNaYgKyB1t
OW6E1/FIQSGNTAqfe2vuYUCxDNN5l5RWe+ZnsPmpVkcl0HTr/e0yRfxHBGjKZosq
6B5RuS/VNz7OeFgH3fm5+S7he+QvoJwPp/n2AqQ5EcWKFGh3ljRF16M0TNdeFKnp
fXcL/mIv6ucF9UFYF+SZRtdN7sX5jcPlvCA0mzhcev5b2XuQ8SqCynkrzj9MiOUj
E56SZLWi4PuNL+slsaAOM1koC2XY37bJNrGdeXlLEx7oa+dIcHAZV1mxQoNQCw2D
SyeWls4AufvEFSw6tmAyBlx6z4nnVCBjPnbCAlDP2eeyv6ohxVx/xVbAMpQta1an
roWr8nS9xIaRUtv1xWE6/QPFLmO8GeZh5c4Qb/sntf2Bofos7Yy5aTO5CeN8W6MG
9f6L9cRHsbfZrol5PvmrTXDZNlQLSltnjHCad93dpEPVMOL8x0HMCxjDu3jtgLAl
OXhLZCL8kR/C6WLuWeDPWyjz+sfHQkw5kyvo8ddah/ERcws7QGRuNd7Xxda2MlVy
0T9nylsob3EXFKXfGfVb+6HioS68bz6q+QuJ2rKp9DO2Ynfi76DLZ7Xyt7K61fOC
bYyFX/ETJzazc1qFyTPE685e9qvFq5Wzg5TbAoCPNL0XOLP1QBrIie+AN2wKeClV
BuBiJRBePxn4t1GSD1QK4JlsUkFjzDkO6Ns1F8t2gRz/AxchdeV3+bWYS9hgygZO
unIh6CXeGc7fJ2ee2rRSSoICL9rWRu+4s9PZwWevLQcOHWocGe96FeSBnCOASr2E
N9vihNknJxI/q76d3XL5BkjEMxl58uZ5jJ5LPoTQCA9+gQ9WeGzDpkiYyTR77V/o
V08J1KlQreCFQgkwXiWJTI569O+2S1XuHM7RkxkZ3fmObTF5nEWC7vY7e/pP7iuv
gmHdu421I/RAj6F9tN62n6YKOeCEy+CRQfdoID1TZ68oySsShF3XtMI5SznPo3nF
jaVsVRbBQCC9/l29GXKFp4AnDbd7sjEgRHoGPxTVRWnGBOKXlJh8/5IOObSZe0F+
fXGYIGo5xNRGiJhKZRHeY27M2duxh4kxMXpyT95TdG664ifdxHecS6Q0whrgjYQE
CUsuCpVldF60jc0GNJJHW6BWF8TB99dYeTCLogMFTA1bjaeZjvHQLjOwjdpXKmq0
0GPKUzSyoQpobSZtrcYjinF6sL+X0vGZEVZRDRQ1aAvxGSIqp7pp2FChUhTzBB/G
z4VsV/LUAhJvL9V+J/HulOvGeUB5rSqduZ7nEzFLpHFstD5KR4u+XnajhGYHHtOU
ZxVkahdGqzwdOWgQjZEiV3IfyR99XFgMs6H02Jg1c5W7hbdcNvAHAZvetCMtWhzD
YgXgzx/sWzZ9SccjyYrta/AMIKHmu2SomkNxQvTWT3PEKJjbo6TCXvxst59lxotL
5MTz0zMfPnlIYCUqBsGer+iFQUiXbS4z0VdpwNv0s+0TdKlnayCR0v4gT3xVc7M9
XbpqBBfi2E5wfuzJuwhCKhN4bsXoykfsyRMu0UrHr1/BdgpHCSB7H3cke+RgPpAn
/RjAoBej91pxb+M3V8eaLu2X2ULOgadvwwMmeZga2QYAmEFCKrzMzX3NQGxed13w
/8VySe3DLP++gn54EkjZx13O4fooOcUdVxCw1MxNlWSq2LmGVXOCh6ezdOoGvYUJ
WGapgFqqOd+2tv8sKoE/ya+TEft2D2cVFnSofn6bn6ipkg4PpMTk666bqfntJcID
0wVIAiN3GOGGSu8CcERMwhpjHHpc6IIeIHk+VlLOkLMvswCCdiaN7sncwOOcq7kU
yd4eLr6tzdUhBTccs71eXozEjTC7wBx2+08r03iP1OriKCqM97IShJbQysbazqu9
43aID8lPLlJFq9u98ElQFrX6f0PovBfgo+hSyRjj2wyMcrG2zay8qab6KLrRX/pp
ThRgD3B02Yq6IslDg2hsOA2DUFicgiM0cCBtpnS6vR8b4J5L8aP7W+9ilLAMd0hR
lor1QBHqz1Jh/Cr4+C6MXwPfvf4CVNswVU867iajW85nqMdGR7WXjZ3Gi2Wnu1S3
GWgMyrnR/+rxk/8lUR/sCjK0C058LcHEMrlzuQkh0TGB3pGtQqat6NzWNJqG08GR
QsRBantUJ45geAG1Q8Fo3etyPEE35YOWoFm7RgD/IPVD8778lIZavC7a/TO0hCNy
rG0rbtird/Je6K9th+iRkhaqyNfmsgWFkq8l8yAqGIUzMB68Us6OQHYgtc19v7nC
iG+FbtwEmwCNo3qWm/1EqDbVyzDAkKBylCANGiiAHwTS4F83g4v4NnQtWxzZJTay
z5t99RqQxqQCWnsKo/LmCF7u6GWmkbPGBk5ZjxsQkwsm/j9xZcp1Dy1TDLHPMyp+
KsPGLfKYE0vLZYe/EO6DJ2NYoOGwW1BBP2jKfCiDsaGFvsYcl17m13Osehd98j6c
z0N4SzjkOyWXwyK3CIcNry3lcrlk2Rc8JEROxMwsFigDe9kgggLOkkCV6ZEp3Zy4
yRiXMk6HyMy3ekn/ME0oHyy9+++zl72qLh175caodGYDWnsnMGbmOIbe5WBuJg6o
AWC21rcUnnERU922pnQfcKS/ndo6V8n8nx2HgZJW3482sAjh3pmJ/I/hCcs9QW25
Iebgu3YWbP0KifP6SIGop5xhfVl9XF7Y+wiiCqWK/K0tMrcH3dNERTaIKvIqVylG
D8QUCSCyctedBb6WBruSxiXMMnrJjD6gRF6XfFbgfyi0cj9xjGm7/vb1FPZR/NlJ
on+TqM6+LOtqsJ+ChV3x4aiDBeBGB+Z0g689kDE0FpQtjHJEzcFfbdQU63QUYNH3
NuVqHKmiWOidcYXPKzzQ2vMt5L+EnVLqZqkmZZXYNT3f1e3ql5gnImZIScrk6Txk
R/LbIOrnIC0ISX5Pke1FbMd7qo/+ziVV70QhR6CzdKBrXhkYzrndxkLo8mWxjfL9
+aY4nmbgyqqxnlkvvPvH+tDU6vvddMhYxbH7r+3NlD04wQt3COi4iKtoAWj2rN3O
/CbRQS+3d8fOYdfklUVCkPKAF7/C0NFDoWAioOBy+mliSM4MCAYsGScNQSYotzqp
/uYTcTnVVnCwbLCJfI0mX/mEKb/afYv3h9jYrBEbBCb0WuqgBIIu6mEqXgOxOE7y
cHW9Mq/DIfdpeq92ihWbn8gvmwvRHoUPhGtF434DBWNucoWOkffxiMWe/hgJ4oOH
n24SvM5MncckZgLNkkSc38TaB6rROQ+S3RHf4zoeblPDs44Ch8/ksu9HGRnFkwiT
WYnhDfhFs7VscOZP6tlGjatqsRIEQZz6vgd/8jUUkAFUzxm1R10cwWPeZ8Cp7eEI
hpIEBkvngGsyYeowbXZccaV8q1zEGRnjQ2BfoZBt6pRcGVR9ZicE1/5ZNrtSeaAL
nOJ/dINUyYTzNm/3pDW3luTtPFW/n/vA7ySPVVrqiss9JDfiDdVF8aW24Zrcriez
1KYodUvl3fSCsJi8xuNX/NmfifRkI+PLvNjfnme1ujuS1DOLuM09qFdLou+1n4ry
B1QOC4GL1GXc0QLgeByz6b7qjewtKRx+EFh6XxQ9JeclvodS5Z6hX1kBMvf1dIWJ
Tt90ZOqfo2OVKrnfMbDQT2gWLijz3+UDe/PR7rfVIHOKIceKItxiIfB69rEpxgGq
D/qbkDvG7VfbcUvPHLPyBYayWa9Yc5DWjp72mOEIT8O2vmMoiQIMMw6t/1VqTcWD
zmrT+v5soUKEzDjQ8fWhK58VonNm+Ft+4Mhbe70g9bAoC7zhSW7vTZoyy6pHmR8O
6UTvVWxb8Jc1sx8OMDsE1FiI18CmKgj7Okutv0eboPbBLkt+ikyNftvk7GonhFjc
ytQFX+ko+MoQpcgjwUn5BzutnABEwvyr6Ltpylz8fmrg88zDNmh3kXNnhQaoN1bA
Qdf+iKiMX9futvsQNIQMo86CzI0E7j+8rawOOp+LkoT8XOVcONvp9FmblD8dYY4x
Ny+IcD81Zgg/dKHhNV0RfRDznJ1UcNLbXjX6VMaWtTlVOCGRypcCutO0hWKU3BXH
RWii4EGEyFHwywgYjjpSK5szZiqX5BL7paQwwdgabI2IvkZFL2aQNG7p15s9sEeY
HhkSo2fioF+ikNr6Vdoggsiaz4d1T2owEwfOfwgM7+37HvD+nuGAca/p1yrReEUf
90Mk4zDYYkDjUeQE4UAh0BL9pEfhg5pP43iL51EJbTUNDGnCtxMZz1oz+2JQNEsP
MUydXOeo+emOrDMinD13OfXkTu2n2cLOy3S0bgzZnJRJp8jxYkA6Q58V9m3GtfyS
d/lN6B66uiHFLluJClJ57eYsxJsrjMqmJg09N0rb2teBGBQSYanmLE8yxbjVSl/g
d7ibLgyBqiZkFt9DEX2QJ8oBd/gQA2RItXUmwHxgEQJsAo491Gk+4cnTynnZv0HC
sRioxUwtawwT2rUxpTUU4zp+5UDhX+CZYjOVXnRDVMkpw1bCNJdjJhqRYKeNNyB3
D8qqqMS7Mmu65k2vJoOilAlOn+Vwl5RpvTCUvahy/9zRSDNJDFT2ZGzSql9Dampn
NU8N8tzsXSfi2us73zzgBUsBkl8BrIssondia88ZSJ2WaRJ+KBF0p8nw2tsFxOKY
U1aPz06hGxLHf+96QMrrh6vsnNJb4x4mfdTD9beLnmomEAfUJ8h9PDDCJbGbXl4t
DT1y0I6s81zg2qlOvfbeaGO+5fJcfnCNDJmLJCeHq+1NFQKXY6etVpO322uYROfp
zhggpZbBZRPAV5uo1XnaLf4toHMUxZXTfr7mCUY/J4Giqqgv7dmPwFwEK/JMKJAd
PpmLZMABqL0RT4pUy5Mzt5xLMFYNWsFTrDIDjyD/YEq1u2SLBz1yLPO980NxDj2q
kCOMx13UpiVDGoKiKrIbw0jay2TZYOqOkwQtlfcbzwHvBtITpC2lGqX/mIwDh1mu
KaZCpRO6QTf9kf3mgQo7RqhYrgfjXlB7RWpcjHm11aNM3aYiBLZ+j4JNFrydv1E2
ClG8mkZFRKbt6FCq8bxeCRXe8drSBFu1D2m6nawcDTUauf9L0b5KhHSS/ZoGj1EV
KkZFkt1TqRfEeqDSqDVcnRmxYz4Fy323tyPEO5qkDtlb4K0XlpOF7QpT82sAUbay
EcgsqCxcmV5CKyQ4TyBKaTUyOSMS1ERem99YBX1xNMedCC4c0A0DaK6mlIJXBuit
oilm6NvIBc4hbdb4KT17EfCE3a/pz6t3Y1JLNIjzkly/RiYVfLLcRgF2MzxTpBfK
RNiuHlIis9eAZG/4U44eb3K3BjF9LUpXIWaCaCxFOhWDhe/8eotvDkfb4OC5Iisv
J4wppBbuZRINJrazcCEhHdDKEGSobYRS2M1FfEBO76g9nbIMBWFn7Y3mqLS+/UJ6
CWJkJdHtmWyN7AS8+m2nhREy8XXmB+8EbDMIzQ4+XQWrlmU8SUFvoLUP3sWJhKi4
rCh83POnJSN17yPxMWYr6yT6J/ZLoGOjjIwbrjPJm4f043WY/X1AC6H2RQFUyKtj
JgS77Km3PfmxrXyCRoTLRlXq5bR6DKVpDMAEcABdxc5FQacJBAzbYjZxpWB/3hmL
7pGDFWUwlxs0O+ddryex0vvIVAMNNwvW3y+BDEvMkydrEx86HaiIg5zlamgZbbuI
61iNUXiVapLUaSE0Gnl1PYNuX64FaSCSyCqR6kjf98yncdIpbyQR5Hw+eLPcVGGC
tZ+J5pgCWHfjf2lBu7LhxIvUERq2jMrZ5k0hJRTL5Wmpu+5C+SnFMU3OdDFMHWhM
sST50vKn7GlKIDpKibtYL/fegoyVtkZ0r+/0d4G4rlqbhwNA+ezRX/zQfSp0IELQ
sjaUtzPsn+brrcQqPADF9LdYFaQWAEVrBtl/LWsh1kOJ1Hnaf7NpuiEWIUOPgDGL
k0U7vgvM3nw5KOTiayXzAYobfVg7iRNXAYuIdWpdL9vLAcYXQZuzgsk0rsgME9+G
liiEb3yGBFf/p2ON/4rt8c5XUl8NyYVqXT0JapiEBWdi2u/wgerrmHjAZTLvVMAY
eiPhPBiegvp9l9hi0ZkwsEAMyXDUvLAB894Twe+SUoXx9ITRnq4oOhoU+U/f0LIO
pjuZMP34i88l+4i8AE91UcqYgR3ekpa7Gl4myWU9McTQz+1w3KBtASOv3nEx2OKb
urSgoYRwtQchXd2IQsvBu38S6coO9yx98Ib8HzOotqWEDYDc0rZvfn4iNck1/y5k
4V1K/rCXSjx34641zaNvfZN8c3EkGFvO32BCsNw9fREmEiq6FDoeIUYpHHOyElHW
DdBT2pC8O/2addrrUi+4xavKKRvDqy4l0UyDBpAik+Gbae9VwTgW0aXf6RvMV/hl
/z2AGpTr9pigxhl2arWP0sYby5g6HaQJ+ObLoICpp3poq3rLqOFTUVRSwYrhZSS3
EDLXOvr+GxY/JVPvAAoBxznDKpRI8UY7E7tkpefgBLbNBUYOrPCf4qzc3oxIEaYi
Vas85FwPl0PEcROjNt05tfe034UWA6lrzOJHCPTV/AfxdZ4PCaqq+J1i/lLdXT6H
4t7bvNnXDii0CeXVMCWDEu8XsfIjLXoOOiFbT1xNfz+ZwRAafwN2itiECVLtNQI5
AZ2qqSNLoHwMP5NKskL+1BS77wPz4wXG0QBRAs8BPRZFVf3WoSJyNhke9Aq3f5mI
vhhzpoCNBtOzKy57Ye5VZjjlq7FX/8dMW6OXzzVAWTmpAkyenNnYANCAXUUu98S4
btPPJjHnzQiMuG2fAn/PgErrn7GtmOFKs97J/D9O84JvgdnIgKly0IgpM4TuHcFh
KoEJZ1QQO0gMITZ/1cntiEVdbLIiAjoDDAWLhptf2DrrBuPsP+S4qfTIH6f5UA/Q
/4K29aikaiiA7NXXDcEeU69LFNd/DfdNIC+0MX7r7rJR9mGY20NvhQ9SuwygFDHa
9Wv3cuFTl40B88iVDSnfWPJylAp06gOWGMcChyJFxnhnLOy3W4xa7BdYnF0u2/Am
R5NbmiJx985ywNBuBLZF+WHrKeDekHq5WjBu7U/WUq2DP7phxaxLTnfzZKsA4Ca9
J8y5HzNUFGqtQmfsuMMr/IMXGiAIyOqnopchxPVHQozM26kNr6QCJ8RikQpM0Bn2
y4zZEDGdRtzDNk94W25q8fJb6F0WRLi4ks178Ld3y/enyqlasc4vx0bsfBewDCTh
ARx+F2FmqyBqoMDm07W2Io+c/5Y+2eho4psIkLQPWLio5o1w3LhCQJqNzcFh3aKX
Jf71Y+C05/kFTspjK6MzPapoxbIvzUsO5jGNPRUdmHy2WQz/32wYFK76i0RElj4w
AYVv5L8oYlxJ8yn+yrnnXEvhTvMhMg0WD+KTEblOfcIfV6loNv7sy7nvY6+jbdQb
EsPTUEsA07VxAw2+HB9MD/2BDad0GaPeuPgYV6Daf/HezS08UTyO76iyUJ/ch9T8
C0aMoawX9Xt16gWOJAe8W5O/bp0D7NyQ9StOJ1U5joCOonen+XfXF8yEOj5K2FX3
bSS9mG/MA1mzBgOI9W98MnsYPHQKtc8O1BOQ0KMwj6QdzH0pAQbdZH1/BxYf4VFj
zTJF9vq9+B1CHNfrZNqYCk6bhjnSUFbELYlFE7Nv/TI1ZAF+KceEdABFMiyZ8v+L
J9cSqx1vWyhUdWb4krJXo/kBVbEIfZpDqGsu9HdaH/i+oAfVw/ZRbrEiqXEZr+ry
Iwz1XLH/ZgiMk96TCSTj5BcrY8ylmtpxf1Mn+vmYM+0Zz/pPGYikbXoCjXm4TW4y
XUx4bBbXGSBCq0w3Sup/P/GE9FYGgEsqWagzWKBmzkpV43tJFtc0vp6aZs66+6vf
WXxOZalyPMUCIYm/lo8MiX5MMx/L6GsqHiwT22+UQrsFhL7LBf3QkMED3j2OtE9W
/LV6lhMLUMZb6E/1yj2PxP90eaZvZOhg4iCh7h69tX9pLxakYkuruTJhXtd55D7H
e6KBpW3Rkwn/MtiwqtbtAmGsZD3vORRzbXhujViRGkPO0DHmJooNZMV+z+O9RnZS
EE93coCZve9N7q0F5rqVQjYmpRSnEKTn1K1nEQkkEYjBH0zfEA7eFhwDIXiX8ISg
krtoIKF8RBr0NcNJrsTLGWBq8GVT6GosToLKHGCZV2/Qnmf7JSF8o6OrBOwzHwv+
3iTlPcn1v3gLcNCKwq8479aYgg+S/frm95vFJVk/HXBUriqMFQ5pl4Hpmj1VyscO
4cNM6Ls6eCNKTHiYNYJAeeIj84xvmLE0B96VYuYHzliPkTs7+Og6pm1gwj4C9mhq
7WeJYceQZeuApAHGRTJ1TKa95u7mDgc+IciyRDANRRAnDlwNXWHQlW+Uiag/NES4
14mZx+8YTBCVumTj9fL2mGqxTygQ1bdZY0digRlw4li+sbNQcfAAow9YbeJtCVag
Z2bSmUQkzAylCPXDsBfhe3Wdiq0Fy1q9SLRWuXgTSWsR9HnLh5dO8I57cFpak+5W
Wds6R9GDHgzjcOU7ibNtZJlLHqoh0SQbIIY4okEqHP/oRCQC6+/WbtaCMsXN839u
QyhpY+Iy7BV8YTlNXbragOoku1b/ckTS2JhkDBQ7CL232jpe02fF4Z6ogD8Htf8L
OctBgTGJtfE5y/RqLDbWk+xjYzoLuGO20v58WO2XG1bugYTqjXFix3AnlXKhAvWH
ma3Jd1ci7hnLLvAiaseIHuALBI+9QT9KPORiPObVH+NhQRpJ3SpnT0Fc3pjtujUP
KV+DXYZo+uSHrQqLCxH6RIOJVECWEq/WMAnZ0JP5W+YH3gaLZdwR+oRY0fc4/cEP
392niM7iU+Cf34Sl+fNUeJV6DvGGWqX3+Vvn4KSk+BcUfdEzKOkNymr6caawfk2R
WsBaAOKcQmKbV0OHuYDYpSfZ6qrqeTWlVhCcceK31gMnX6jvWnNQSouFLA8QC3sl
itEF3w+EfG+D/MCpk5KzIPf4JlxZ6nOctnX7/V9fgSPcB6jQjuT57yNds/flndZz
zsUfTc/TyH2MQQm7Ww/RDskEIzTJVoIBnRQerAIgiy0XqcN4l0Mfsul54t+i1XDm
RAE4RjhTd03KFPaymwQvtDSV54qS/X0A//nGNi41PFm3UwDG92x734hiQVunl3Jt
3eUZOLAuYY+srXlULTigke+h2fn5I2A/6YoYY3VA0VuOGy2TjgX0S3GG2LnOtNkK
Z+honP6q/c0ljT1ZieBnotjvhnrfwkGKxA2cV8nZvvIoleK7chZB0trak3uLw4x7
VGpcAp6YkGGrF/fCfeO6FR9F3tAbPh9YUaTNXac8PHDSEE6h8JDrWEbWeK/MVu9H
rQ6B00XKAkx/CgmFyn9bp4oyNJ1xngDb0/wsNtZKl7v+F/ShFGbJ/g5yN+UQJfLR
dHkywjtwVhzc6ejUaxWnZPe9unSP2pawcb46Va0maMiFzBp638H9DB9UHgXdweyL
G6xyrX+TDQ42mxaTGcl6+hvpw73kHYzQ1R/8WrVBQMA+Oxey81vzQWbKdMJC/8Mz
j7cKYnmNAnxfHVLiWmjk5nfBfrgZoHSzJHtiS6ec8prVsNUh07DuBvBq25jG3cz5
1U8++J/ci8Q0yQFlZCLzKm7NWgKUPNEkjiCNpbklbyPPKprnvyb9GViiVA0KjEKp
3davNKib+9naBVrI/a6BUighV5UYXNMVTdx/Uiyd0pr7RJOx3YhWVSYFdc8W6bgP
Tubb4TGQpaP/IBa5roTNj14tt5341siv1dIr26gyz0lXqbHs+vKfFiEMe3BGdFpG
klT7DAIEsNWFy+3lnQSgWuahud9R/iLmK1GgnGExBYRzPdZ1AvEDjMiE+lkydyOs
sUPi/DbrE5SZObkMRSrc+KArqYrLCAc2zSFVA0si3f18Kgz8WflKG09bUoqqbuWC
T9LzVU+CpdzaqPgCtmfsw5aMvDwMOVo1znteqCdvoCwK2B5UxlFSnvLkevr3TCny
OIM3WPRM6mHgeO8HpIVa0X1iaDd3KQk1gd/zjc4tsIG2d8Hgff7jbDoDvnqFIM3m
2M4gMNRW/SJQcYd1WbYweTJZuYjIJg1XKW8a5+uoafByYbE53Fo9J49Oku2cO1L2
LxaC2ASXicZxfo14OgQ074GxA/r3xsHv5ITTUbCYpVopkOzU91ZcpC8avjMO+IIg
yK8Is9/1wK6lTkXcGjM9FWXo4c1QOFWV6QIM8P1qwafHxf2yg6fyxVbS9H66SzQo
ps4SnDdK94cflCA6CsZeAwOg9I4QxVqSJJncWnF5rgroLfldcU0pFN2dmdHn5CvS
jyc8FOYteWWwgjUdI1j08teh/BbprV1AKWeanraa+BzQp4QugAoWO5mSxf20htnc
yCMBZNyKGu5TcMJh8ZtWv0pP5hsZZau2N/cB5fQQFTfo+UUPzmuwkh+pYj+fdvGS
uOL166aFkwRaRwveA+hsm3Oo/rcdqAOBskOJop7ANfOxP3YxhD5EHKdJMI8Chs5I
ttkKTsGykD715ZbcmbB1Dl9HYjOxDxLsBX1HE+I+hXNeEXJhmR/2zjst2KJ4jhq3
bZ7HhqYi55YViDS/FzziNFuNPzCO0sq9Y3s0r16Y2x3w36fxtHYyVoLdEAemCjen
7PRaaSOClWXhudBAZNZqxxLXj9i3wxjVAjslDB85X8CHkbB8Ios86BcsX1zbtnQJ
K635rdq7FvOovUa/zEQb3wUFK/Ul/THAGr9IjPQ68F7DAFHOZRbw5VS7PNHy/1sf
JwWFdPs0eMfTQw3b2UJ5UlitdMavJLEku5rOJgZ3Q47PpwZw9cJiM0FRexdJjGQL
x9cv0sx062O4+wDk+RPUyQXCJGnvG+Z9ljIBgRJvoCpEYeA4caWtWUvdt6rKMGkF
67yMhilK7b/btN3j4D5lsEAX72tGbPjJc6gpIl/kREwAZ/6lHeuUtvXxkKYbvhs9
7TgBk2ggkEhsR535ZhurUkC/hnmuwNsrDfH1MzvSDA+r/0rHCvV/VaAYXVbDya95
YTPQhVKKZEOApdWBEFAV8imZeWk60ic2lKVlLgh8XdC56j8yLwBp5e119bAqWVf8
HOPqWYwTwcCKYBQjUHRcE10H3x6LHhOi+Gz54YJH4m4617e17gtauE9HN9OdIkHQ
wG25x+uA+YsIH592/VDUuTn8/5oQmYCb/BiHMoSHE7KsaA1muURCuB1AexXHHl9a
XBH5OghUgyH6UBcEEWdjZABB4Tn9voE1RLaIwP1oQ0D57XrYaTx5+JBQvO/E+B7V
oTToSOw3IQ37Ga00PtNboRTkfUlw6vriZMnt1SlXEGGJtnlU94Zpp83EBqqGzIfD
hBjY9wq9dD8avvzqd561KvupMWXCe1tFNNo3ridz/2Ca7HoTGwyQ3kmoBAO3fyt3
/KWkIuyycONaY81McJXOSJbQu4gKXtLc+ugjIHhI/067MkgH7AcLofqabw5gF7Fb
imdw4U1VphjCPpJVbJROliLZ9WGndDUjyMk8KF3BcTfSTh2m9OO9FE6iki5jjrTL
otlePre+DnwpR/gQ0oX9lxQiLWD9N4utKIKGrcBod5bG6ngjHIDhhNsbkRdSqr2b
tAd6D+5mgDg+7dwa6RJuzi1C/D1k75k1djF9Z/1yqvtCHMa8VhRoGZh0Ney6dMKV
9jfyVWSDOWL8W6RDF6KFcj20nyOJNN5I7r6KG9t07Cv1cwPk2SKQphcu9h3NPkyK
+NBr8K4fAB/ElYd8DEa3l5vUQNbwu6628Dc0INJqkagVBMoiEhC37FertfH4V6FD
ywtQ1Qb9kcbXmIpbJDFeVCJNRfJ3nxA+v3bIdht31mhrxoWfkOZtqFSKnfPqaUKY
EuxJofH1gUHWHVdjb1uQX/cYiUb434PtwAZOF//YiAlYtoayzT3SOS6vw/d54rfy
CmFaG8Z4FJ8Vqd3jPcdFz7aQ0a/BhZ3n4PkDCP/Efoetma9buAi1tcxtqtv8Kf9B
cM26IbjmM/5jsDxxEHY6lI1ndIoY91fNw3Ep/zuUx31yw72mYzE51Pd1Sha6KeBe
aMnrqHCWvpFXx6xEd/PrNO/yu/IDYSPXT7L1xILr0H9lpTA3gGz4dtMAzxFT05TU
OHCWqPpwHEvCAZ+gxe0vs8TQfn7cs4kZ4pjxWm9I6sGqE208cufsetniZiMWUQ/s
YDmNnKokhbjZPQRjjbc+zzfW/1KWyiBTIuymp3s7G/pS4SMJiEwCTo87+XnkEddo
Mt2g318p0mErcko3dmPDZKkkLEwHd5LPTitalz5+GiborwB7uTFaRWYi0yEmgDgg
3bFh7km96+xs3AUFBDN2HGE/f5/Sw8pxJM0oNpQ+ofYdI4rE4fdAmNU9Uc+EMzzw
D7IY3UUZWang6dtShwZxVqXIlDpWB//epzJbWFArtuRl8B2biZkM8ePHXMbU8eUa
mruUoLh5wd+0E1ZmNaKUVBeKDewqRbSXoOjhfZ3yjXrCYHr8vGI1kaGLBhx5sG3A
V8RUsGkrXrdk6aG2grgWu28cyAQUEFT1CretGaQ7r3DhruOATyPazhxYpQX/iun8
HX3BOrKgKNE6IhbE6LaMm+Lav0teoKZvFpDCNoDGqYkGptzw9Og+4KRz4fUpdTOU
Xosen2EPkYagJDG6PcsNlJDEi57riJOOemtlZwBGG+E0f+TskB1gE4pxmaMPXaUq
S6WFtUW1AsBMFCSETuDE+IiUz3spG+aHrtGYIHS92aRwxg3oqTTBybBKNKDH7FhC
2MDxg1dVcyA84ZwVEbcTvDuxqunOyPLZg0dvK6rXb42P9jRG6YaA2YvXQcZm1une
Hx0eCnmEeDhEb1jO26YeoAzjEa5jyROGDw9csuMw2mso6Tvwl02NAt6IyWnOq0/4
LXX+nqyYGrU2jWCutjj2FX4WrBJS69KIDO1IBge41HEC/FK/ThGftrB/4XbAU6EG
HGWvVW7/jvy+ZjG4G2koEdO5jb16CF8AvgBvccucmGUTK4nqbnYP+kAI5ovfjrvw
oenTIdoO9jdIdEjNcrddsSZklqYSjZhGPVi2XjMzTGzocV9j/5IL4RAs4vBykczX
8tsDN6ETYjp/07ZIPd13ZNZeH9J3ItiNPYn7dknsz2KXMH97buHu98tjtciJze7m
MwbSapoLrh8ZGRT1/zi1S+HAHuUUV7ueJl+9kAcbff+DLX/vDM9CY/hlKc/4h09f
D1ffcgy+Cz6tqEeBWVQf0qYu859m8mRVxYFqnl8UmoHPp5U7wwpEpnmok7QkqADl
NOkkk+3od/SDa/h/mQx3vS0hClTFcOEpJeFrNtQmlEn6tZJMWuqoiycJ91qJJS/Y
0BTCMvgvnWmxSCnhQz6KBKiNBUcz0RxlR5zxs/1YvV7ZixElonF72Hy7URUlXVSq
taMXEBbM7Lapj+ElsxqiGLFRZLkbB6QPLAmK16JEM5jKfPJOZ25rBT9r8tnAqUR+
wgXr3w0hoyrjCerEAn3C9WOhVPrRalZ+hyOUGenh0zP5wSpEh2G3mVuugVdLl7Gp
PugnBJO032/AaZQi2FUSZ/HMeHDKIo/96fzOsqFTNal/37RSTEI6PngQSxKC9UPt
kzn2m1q6oI9u0lekkcaofq14h9lm2o69YrI2za8dk4jwuubLrsAqbvm2otlzsfgq
qDWL7bwhnLxTpJn+hlQNyZ7Lssxuh7yKHvUQrZttYsI2Q6q55eJlb4WrB9/l4Mfx
6/d4fc2E8LjyMajcMHywdvNUoEz8jXg+tCrKUmhqPieMBEabkdgK6U6vHQYG1DOU
20YlULc8+eQMJFWqmWLeRAxk49GdRQbzSEwv1iST+7WszaAEfXK1+gXsBS1zqZna
GRyvPuPhAlsjibUebGBzwWgw3SQgazVevAZ+bigpJZWNGJ6bJfJAUsrrGlx9CJYF
m08gVqtsvHenh1j3ssB3uyKHpM3xgMpxgMQSqAYCElbKENtpWPdyub7m8pnqH2iO
MD9As5cpAznne5vnanuNbarrWVIp12yKkW0eZQRO5jmh/tLYhEVbAz2wYub9OU/k
ySJDuPKR/OkDZMtS8p6FDqlGj83HrOrFpP4OiD03xJjv/EDXKGz0ydWIoVyccVw2
m8y1ON637HkBFEs7wNgs5Tby2uDiiLHl5wwmltLmrP8APkwM1xq2omLsgXQd0uue
4prP6zgmE7D6llKyEO5Q9J2HbKCPHAgQ3nQezfmU/stT4Sgp0d4/92K5Nmb2uKd9
808XX+IbNIG2laD2Ay7rVg4hh1pWnoRhv8TX6tEjfHSUOWoRMken7R8SToTEBFtl
6GIf4ZpDqgMkF+7m/tNb4TcwIBO4mzJdsriKQsxh6P5Mm0jEH7C4TmDfA3MxgeJj
aLuDTQxs1nXn0CyXDm2xCKzKgA/+jJzSQqKE0Se0U1h/ajFfKg72kL7XaIISDsm3
p5fNbWG/TH45XrWlYLU5LcUB8mytpNhZThTzbB+qCheRLuu84oyoDr9bR18ADuHP
L+ISZuc2gLzbUZWMzzieQo0boWJIgFJnfQEtICeYzCmTPuG8ut9Ynq1N9XObCXcj
xd1/p5CMMUxHViz1J2Dt3Aq8WsqyWmsmVtOzxcDlPO3OoAI6P3CPMwNfp/TzkmC2
cKUVKs+EbasWZi//U5Xq8H8BjW3oWF7IlHwzebYVPVI3iyhrKguakgGr/HFHPfwa
SZp/i9IUsB5XfUNZNAXGLB6zOhipf2xxB/p8zizxOIR2f7R/KOAaE9dD+qB88j13
Y/iW7jAP/A3Kd0c7eh/6hoHCK9feW0gEU5yB1tE2nCEOJY8iypR5ldyWZwCnsaJE
R218/JlVCd7XUJct87wuqisyzvM1tNgQ6FTm1nkGPhwDOvxRB4Z3S3G5NzTogRTF
fMAJcseDrgjqb+FN5B6OtlNA4olI0YAd6JVhjwlJLQKXt3xbr6Qa1hi4iYuZ7Alb
0cjc0PSFrFsmC5lNBa7iJm6ZzpUSKODhLlLWYW2+kTkzSphYNB4DB6Ef3xLLGF3g
FWFaCJ0u8CvydBQG5tbRpyUATC+OnzPSRvehaqDD72L46xrcHrjo2y9NzcI3DRs6
/VMMuN3YNov8e2u9zCTtWF92eUZaaZyrx6oNxGYc8tYInJ4lXiAo8m3K5Glxqp8v
rbU2+lwopHN35GGVJrzrbYeZTLQgN1rc6HmHxfvjjEAtbSuYhXqS1vxb4Bq2JjNV
zrJEUR+AfAArkUQMY2LmXrJNvu/bJWGJWTvxCca08i4vsYZIHIlTd2RfgjRZnViG
OVSTYMdRIIr5Qw1KQfZQ7me8/oxcL2LULPrPD5UeNwo8d/pGuOVdkhSA3S4soMI9
6LzSbMSygywU3RfRrJY5T6q8vNV9pShK32OMR4EoJLEymnux1tJpVX7Y/ceZZbKp
FD615UeZQA5pB+FblaOI8yBAruQADc4ay9UUxvl305EHoX0sQuWZrrPJJGKbXixd
FruJKO0rD47aLfGtQftXa5wITNe4MDD3B+tPBSztHPZ3z34zXiUZWXVbba39csu7
BKFHZx+hOlMMFXzMFc4fjdHYAgq1uWxmeII7Bj25Pe7eLVrz0qWw8mOEerLk1jSA
zj8a1APH/LLaxVqLhO81QLmqBez5IOjAY1P+5wgf6NTjj9cw1BBbp5SlbstK4aCI
xfnbK8m5b2ClClAhbk6BZtM7489Mf077d8fvdXyvN8jsh6sOKRPhcT005K9bv3CG
xveRVfgqcbBMfwxYbBPmG31Nf4QEUke+p7tzxT4LvKAu4lEFAtQHZAr87I4bWImn
X4LjrRtAcLbM0d43X1GASLwHJL3klFDPhAxetSIB8Q9RiKvnRQXXFKE9/bjCNwDP
Rn3ReYBY/+1GhCoEZfAtnsmpjdD3w1rKRod8Ang2nfT5YaDgSjcoM/yXnQzUWqyM
t20ZLsXAd54KI3mz1KJdKgkyzT8EeaNxRdpgf4T8Sx6c9FyzQbv8kYuRjgU+SJax
Y6aeE9jX64Ll6edeyufaF2gUwHnuuVG1jWck9vGbhfjB3h1va4PfE6YyF/37JBs+
7C7TGr4N+dWi1P75ydm36o4v3gEVnJwH/2LkqKcY5AF2X/Gpb5fgH2Q2d1TrBTAX
1o0cs+HrfXUy6lw1nLEwbgZipRm0d3bKyRGWycRMu4KzWg5SsT7dNpCGytKYK9pL
T5kB9/Llqh/IunaUee9t3lYos7rBMd6qSr2VFDj2d43M5bBAwWjzP9XPqBRVz1cH
qhOMoERctxB7U53gqLbJhA1h69Ey3inMeSB9JO8W5ZqeHJPHnG3m644qBsaT+ui8
mC7YVTRkOAGzS+HM+yQhnaI8bMg9PuXqWrGvbYbPh0VR5Okc1ZYOJpU7wd+2yA+s
iXs15urD16ISvC9fYpinl8eQ/sLtl4A7lviBYnZItNrHwE18U8LzLNv4fgFgtlHu
slNuBhRUs0c+F6XW7avNfkACqJfHFuPrD2cGaT6gbhYdSay4PqxnVp4VgyHipUvO
Fh7FIjVTmsJXmFXFQN9xCOYSsn6E7Vl5In//upeFiNysEtwj0URB/stoQqws1I2j
2LYPaptljj6YYOst/kem+2PQNqAVNVAnUAL+9LLebLfdrANbWdlqEF96uaLGL8Wq
MaOpK8gqh5h307PX7MqsPgjTiDtuyqQskV7Iegf8WXgIImIVGRwSN4JlqHGf4vow
G4YzTthGIqCfiuWov0DhZlWurLDYprlmTrQQQUBOgXb/kQ7sq9wuTPkP1idyG9nr
iRcUXwPd7z2GxhcERdcuaaI/o7h14vFraUujzfQsVCrJfPiTsPyZHIjal4Aotspk
ZhxIU7sxdNG9qhBcI6od16ZOCngl9KcA8F6ZPxeEYhhl/NmbMgUJ40ZFkgIOsVdT
9Hpnaq2/NQmajuxGKNLOb2HmMMlWTMFmXvKUzhJPbG2OzEIgoFj2v12SvPih2Tg9
KiwV7zspsAUDRrfn3WMOnwmq4R+jVlQ3KcKw97z9DyfleTzzAU69caq4yaBJsPWS
a+6KoYtfzBdp6cUzShFCzdHZGovxYDId17bLiyrSA2B+MlNPDGqTkJUke8N0He3c
DB3rBiGnfVWqos1X6mxUMDwCunvYaYvMphJG5WkXA95bowHAHTcmXKRZtZgt0P51
jJGRxciMhOy5VWkxuziVyDnRC+gun57j5wchsbpnz1bhVV1Tdb8nKxAZK3hm06Gy
KVG9N+E4bCVDcGMxwJdKrAM0auHAlEG5lP4J+WpA7H+7uasIY7QAiIPWQ/8F7NxT
D9mQKFgs9WgFfmQqdMF3ME+nsuNnCp2Vhrncg5m58sDa+kOj3FegfvoaOLnVhzvO
P1vHssmhRQdre4d5xrKJGSdrXWut0k9Pmgp3fe7SRI2FF9BRfKaSfo6WWCb48v4v
BD/sFI0G6ttxgO0jGXtr28aXQBnW4suMFGpvA2+PgT8LxtvDWM9ucrUGIyJlzY6k
+RsiXx+9cBhRvU7gK+sdznh465htM+q0PU1CszLMzvMDnTBTYBZvPhF//Y6LNZaX
dEonNAfQVEO8jj5qqJDOZquO/soLeIj+UqZnipZJX/jdrDLfTiktEeYHSRIzA9Eg
JlvUm9AOh1JcMzRzKiElAurX1A0p0j1V0A4yN4OhbiH/LWsPIvOOk6aZgPgjDAWB
O7JLvLyOfDGigeuA66zIeDGX3MqOr3aRrMkBOHf+gWPaYVTCe3Jg+GA2wnurujds
o6TaHebeneAQHclnxWzPZZbXDq72Psc9toWqHd/bp6FA156veCPCecOUU1h1Z2Ax
4yX/K4Pz1f4KWP8DNL8SVqfHCRYkebh68gxR7i0Lvf563Ns3heI0dQFnhvgPGeRW
uZW4fBlVvQk7hDYycoP5aDL08YQZm+x+A5oH1FhGxu7TcwQcSCK2KXqLPPdcXd4S
mO4/Gcwzc2CaA4BY45kEVm/6DdW754iWsNanEd9aDQuXCY4P4tmUp27ChfwWj0+k
AmpP+r7gg9exBpL8iJPPauFnZS391xHCrf8FaUQjARWHDyG3g/ZZmyImPakk9k7H
+SFcWZkgF1LTiOHIlvlQ6+i+QDXTanXKjzvtocIkmv4EIsjNb50ENXWbHRQBBv8M
f+dEpnhO/gmrXMFSS5Dwp7WSaiMXmWLG0vSCjYj87sRJb5inIlvK/iCJzhJreKDn
Anu8kfroMZn/YKNQFSip3Cvnr08NjWpk+7A25payRFvQX9/BsZ1UqrjrrpBgh4Bg
X8G1aLXeoSs5RhRWdh69+diXx4M0FE3vH8Ly31OIgUYfzfe1eYxpSq7LzZ/An4cG
D94Csnd4lnhE6+syoe/QBQTeFscyY3uZc1+l1xWl0JnuQFRxqv0dqODVxm64MIK6
eTc+72bTB78md0J1K4GyDeGwUaCaeXFmLfjG9zlDAIBCNV++HnpXZCWk2kRvH9ME
iOIj8lE0iRV30kHUYFeklOiAEiK7a5GHA7bZxfJ0IJXu6h4Wnu/yXrnz5x+8j5An
tFiP3OzDLOD0uZs/stgbaX7hmSPE+TDDj6DQXvlNGyVBdEjpGLDNkxG9wh+oP0wX
Z/Pm/lyz9hBddeyqk3MTpVgMM8HPQ+CuwqTUFEltikUNvJ/UbTQYPVCwTzQmw4zU
TCe90/TYFuihLWvXpB4ZODQIM8BlhQ5a/42Q2hsfjLGAxRDaDAXHeAMdq6Py4PV5
3WAe+dlDBTyPwkC5D79W2RIj0hwbxZUbeSlvFCcdS4VTCAE3i7pUwI1MoC0/+p9z
CfLahNv8qzQujcv5eNjgQSih/TZCwrm/L+Ko7WPlpWwC/wBgalHOo71vo4Nl4JKw
GK5FYRPMWhX53iMkDWlr7fuHNKuqKJAnb4WAzD5ntgDBz6w4phSe0YsOczqWlhjB
Sb+PEcuhL9DxcI0pMEru1x7axUxhrDYVQVCHpPdRq1DWWVgenA3KT0RG9m3lINXv
sj/EaDw0TJNtkbLxRD2xMZHe4byaWexXjUtNMI2ivHoipnkSwGfqLD95OskU5YLM
0mnfqJQULxQV+1GHS78jc02ncx0rTsxtaNPuQsQ0fy82kAg8OszdMxRTjbsmF93H
z5ukJUWvnit/zrrIVVEvEbqRnuP3SWB5AI4wFEjh+UKRqlTBAOkONWaCv7P7Ue9S
t5o6zR4z6ZFCt46fDEhcw4GmaBpHxhjJBjARdnqwkSTFe13lKa2qnskOG/T7u9SJ
DbUS/YEu1AOu8g9XuokT29LBj2ozxnl/QkzQHJHUTUQb3FMteFb7iydOgCSg/and
8jpoQPlSoLSN50KktrrZXPZ4vM5UmcjXYVsk4kqxByqeXaXDxRgnitQ9s3ZXgyX6
hQwP86aCqt4knFcfSfi72SxEto1pPRq15Q36KN20j3QHRbbSYUhPjJevHyHbYAxh
Aw0yyYYcpxcqzBzOh9HkYV8FBUpbcRwrqXepScmaMJTK56R2dJs+pCv+QndpVVD+
g7ZJaMpP8kyAin30jMMEiytE4mjQ2g1ja0PUFU/NL6M/Ovn7qdH8mNrumPNA0EEj
4mANbBiXjtfJN/ObatjrsGiUL58zKCYvA7/6KYBq8+SSONUUkIkz1jYOI/ZF2UL5
Lfd+LbrJYM9wA8wm9f+44qhPrqO9QF575Kv3eIApf7v0RV25MMZGbbhmlRuJ5ZeG
cupVpTV3+B6avE2S5AXwmFGNy3ZPL3vag7ART3FseExCOJLW5bcqdm3jS2T4jzxs
OVoyGb+/YDQBjq6hIKf5OTbOQlLyHRcdssuIuuLUTNwxJHGTo9BAyHXKRvYO4Gwe
4d8/Ckr76iuzDJnRRzGxBRMZzrDoZLhbCRFKjdBXnQrFgi50+7qT2Ts+53Hlr0GH
1dpjyvbU/WSgs1CZj1itErWf0PCj3aY3ZfsdS79YcncIyjxhBLhFI08deLAclqlw
/UJdP44mUcMuWtdXUkKzRgLZuXX8BvC1bFkUCt4bz+iB/Ds4qGTDzxernVe5BlzS
ALl0wlUCyfBbHldwaWAveqRA7mOJQZklisipb7YynE2dMPtCdBatMu3o+AVQd6yN
pmPGvVRG4ekMF6P4bbCkKM+YmcxqJOVzMJ8iXyvBbWaHbr7tiRoCzZGhvn83lSdw
8EvtVqJmPNas7yr00S8CKehIK6nKTGJA4ZwQfgGbEatTb8qh4H+dq9Mv0U6mr5jq
WU37zLjDnt2lNRPWDJgnfseX3daoaeVoF9BQJxz6On5fJwnleOVU0XWuQCj2Y6f8
/LUzto0az/n3bga32bhjqgkG2f4Udl2qlSvY6bXF1ntdad7lck6Tf8XKSZB2JTXk
im00drb2lR7KgdJ7kxCPXjq4m41Tn557N5Dp4IWClPmUx5pdvRmi/Hzqx/CAximA
AoTR7as8dR+ieCmmG6RDq1m5MW9otudK2P5zmgsTGMIBFMRJ3OFJsJ2UEYgQh9kb
N18/TmPCrz4gMcJMn/LoIdyE9RTJzZeHK2LOgPR5uv1rteyF86VKd3zv2yDWQFFO
x66R86ahdbY+qPT9APAlc5NFGt9v5ppnIv2at0eV2lZ+iGcNgaSB4N2XD+i/xgXL
82V4WZbFb/4lMBByvHjzn40WKkWkO6/6CTPkLfbG9+W1vsvK5igsw2U5VrG6oUIl
pBd4vcVTh/caO9bcySc6ntgso8/xXOJCYqr+QXx4HzYTBvXvAKir0hG7MLYEFsEx
QYncaLDeMZJNezkop4s1lacQCf5Ibu4u+tZix0nIytnfEys7d7lWZuza46C0bF+p
aO+hhWdao+0d6FETQh00Xr940eZ09wgTrUGqUR3rlUZnq5TppIhZRyWQrR6XkIoJ
LDOIViQfd7/bUvpDpgprZhhovvxDnWZdKM1K5atL+M7Z4qZJUYYhETnKfygxEdHd
2jn3A4kKKsT28YocWKvrD8p5XO7+0GqtZGaOSDMY0sS/S+BYlt7AwGc3gUfqDHeO
6XMbPHJ8TbDCOYBLOHk/FyC50TSQl2pSw2Ga1IpeuPT3uv2H6i58e14PYIO5UbtC
U4pDv+t9GG7YrOHL91l6+3S21l6jGisHbAhxU+85RGRrszXeB0SSZiLbSxt1+DlP
LnMhy3PPR73BOeT8WP28tz1SsPlNkrGNfCbNuivVKq8oTB9J0sgYf6IDM9PSLAzQ
XUFHMU4KiVOn8ae0o4Fg1Obd38QIuDOgyrzXnNw1D9G/s1N0rf2GYqLchMfipAzF
0Xm205HUGTP+4m/1s5XYS7MDAec3JjjUH7bB4Ez00s/bWiurIhpT1CkJ9d12+BVQ
U02WOPgmOIws7p4PrMkto9D4LS+qoWLkExQAyoXsqnnMW5KzWcX0KHLXYZhLNB6b
ZdaKHaQLaPTvHNRNZ+j3PbtxuOvz5dEhHATCu3TVFKwncM14NaYZcZRwhrjQbOXh
Osz80X9Rf9GIa79wEm/+YaIIJE3cuAhXhfoKCxrRV1xD7VBzIqcUoeCRFhyOkHPI
aElaxQyOsbGxxRwZXrPbaF7KQN5lsISFoBbMuWkPIGx2C4x2eUt9N5Wj3epUqQUt
1nB8dhkFg2r3BWtZ6NpJGD4gp2VEY+Rnre+is/R7JP9gI6fISg86sCuZiuVYiWZk
3M6mkraoqoc+n1YwDdi9B2cJM+607GBVZxTrVMdmjN8MBY0gOoIsnmK1rdO46ZzI
Hqit0XPEj3JPqX2O3g/sAPX7XPGoNg9IGTUwlLDl/0VjDqpH1HOZEAOP+Wa3pjzt
4BaqcR2BU0mVT50pETaiSsZ4yu0BALoasHrBWJU8iC3fBrBTW1z+dNj3WWpMFhfG
lJ9RhWYIgBaQ0hMJa0tHBAtf9C9pS9mMyQaeu2zs94O0AEz/QvNR0uc7e4dcy0CZ
ohGuxn9rxktWGLcSf0/xbLR0BJbVYOE22aDrio9ZMcnFx6DV0kxnFROmXFFKdHRl
q/EN3o6PoS/MuS4Hmffob/8s+ksJD411RAIDWWtdYV6bixi5oKj03Pvj6GUrVlcf
iKqGxt7YuPN1MraWYkJEoT16Zhb82CeX65I8nnQXFWfFxtVZAK/xJcEWvE6i+MNT
2flnORvpUW5k2W6Q0SD7TTfSF1Aa3KCjCQ5sBzpK5jc+HGBgQ2m4mMzljTAuLepB
keFf7Y3phYh5UmNDEYUwcDK7UYsILRrz3Yu346zw4d9lVt6dVoDtQfiuGlEAm6ZX
76Kfd/qKECt5ZTttPEsrv/eA08QzW1NdFeMc+QmNtxdxZj7HNp7PJO60FAOgYt6n
6NvBbudnAP7B+a4rp6zP2Gz7NtwZOXNeiW6XvsJzi+Fl536QVyceTQ+weOKsWNk8
ffo/0krECb2KIl49Ra2COMiGi/FN8fJNTWlakJynrlly/MsIeUyiTGZwDpsO9qm9
oxqXyTc3CSYc1qtlmBYrl1LqFCVScmlK2cvJlhZ1DY7WqskCa7BvqqakO++HJ6Jh
KFAYnQsAcCSaMMYzcCj1oHxpvONPdSEloWMxlnRwBTUOEo//fcBdMwqGwQMJzOci
uyaYXGWJ2Yr8HjKFiRt8HlEegzeedA8LTK1ciGsMVGV+ZgjAt4YAEsM4BIjqDfN7
AW+t9zHhkUDClYxjcPtjw6IMkZ0D/X7OUGjiGOiaOBdBCc3ZgahvIFRIyllpAioT
68nuQUngqUW4ipkaDMDuNAzpyvKlw9VTNrOOiEm/DCyW53YpDl55ZYB/BwhTwgXf
Nnb7bIxvEsY2xVyQbqeuxNMSpgSCbU2OCCc0YdhL77y4RbkKrIbBMgto4MfX9slf
a3nS/PTJiXGWvMGo4jruG0BUTBr3pgeTJ5h39UULqqXJJzG5G3Sw9c5qadD8v/3k
Vqy6i+3u906cdvwQTPPxjqd9DNFdIUHvEfg/PdaFC/PdorFxGfCtX68UStVdMtnN
+N/4zgXaEYBwmuDNq4Okb5rGUTVj3bMt/mjBn4fJ48wj+s0kT/qq8U8Pnvnx3yqF
AvXx/89OPy1urO2JPuAFxLAC+y4BQnyV+Vj1YvLYr9YE/13oq5YJJkudyYpR+1ry
Zl+pIST4Zf8ZUHRc7TvUKIfq+FyQvxuZshhsPegWhJjEqkRPlDMvysv52j11K7ZF
7T/U1Hasfz9/kwsQsBamQ/faNWd3Dvd11Z2dZNPwsWlBajI+bbnp40DIvXW9rE6f
cDqBXH3uPzK0QdlfuQW5nwdVZIxBHFtYyKkIeCrczsHK+zyirDvaeNMEeUUyOGAB
tDRSooM8f4buVACLU6Q9ygpo86zSvFSz+QLnwdLtXFr6fdtTOjbkh8tmdhjRi89O
eLv50zojGULcODrjk6TGzU9HvFg8hopqVpjXiVII6yyFbx8iOyN6M2SymUIV0rSU
0hzYKopvCfiOzRfIoyWvtynN68belNH5p952ZdZBSShafUqwnQa7CPkaw6V0orZz
o2WoVmpXPMIWgc1SC4u7AxZPrx8xITAdtObomCVIuL5pqe2HMlMK5c4SrMLPf8Sb
HaTNnIloAWjDLZETfUIiRqqVBH2hd5bDaK6L/qOx29+8LZpZuThAmr9ECMessUb1
pi6IYA2klF0KGAo4s7Fw+ZJBf25U+EBDOmkqnbUirx1Av1NHh2aWeimVS0FndhwM
HGOslK7XEnfJJimpzKPs1rAS84mGG2DRSAeDFZ7f79w5hA/pP84n8p/rOI3U2MWr
VNlu+lyPKgolaAK7CDgsxDIPorii9UjGbHkWhKQygUBKsKnWcZEm3GbAYIdRDki3
vNClJMYOV2RSvDaZCsSv4s8L29ZXtpwRlQUWZ6sqNCPgnF0oQPjP/XRox8SQJX65
1SnmDbvsZ/23BQVbL4QkowzUcPbByTa+h96c65rH8J5FlrgNlCyCnEj+x0I7IDSb
CKuwxxU2hMgRR8Zxw4TYtjzOwaYf2h5PR3yN5HkIU7wrgJNeTmN+OSnA11Jh0WNS
SSEH8VAJP3ebrIR314LyNVFthgmvHC0jHjgacIo90BAX+TKqkU0NlpVyG8kC/hb5
/ejM9RML1FQVSSRUzHIDSYDT6HcslGLNievX4uMNYtjo4CXB7BCkRIBdCiqBq36m
6k+soV7Ca3QKbqxAPyb++KI7ymgw+yz0PCMPq9XGz9gSU6h2H2j1B/Sbkz/xIg0l
LKp++30xZaqQJhR8O1ckMlP6+dgnWRrkFCKN8TqM6lVgHnfR8yzd3+iTKEFCzK3n
0ZLHIXLnJh7uplTnd6EOfmmF7fWrMU8mr8IXbuKGtAXMpeeenz8ZAyMiwuUCMwP1
65Tuno+fwqHe9fDskyn8GLSMwk5efzn3ZlNjNFGqhSqUIVFGoWdLkBXozKQ/7dsf
5mKsSDh3j451t2KrBvW5Zo/OPLKxh4vM1tFGP3Z3O/N4x98P0YCV41JJ1aJlCu4s
BMnSzIl6Nf1bPRTU+sXjW1Q8vwiNMJ15kdgFbQ2YB9fwpKqyrbvT3EWuw0olDq99
SUQHFkpRkMakOzWc45BhG+JxIh+yUNg73qtHS5A3V34R21GLDA3O0kZ7A0IJpBPc
iYbPze0uVEYvwkShVGgDEqC3paBwzFO+F9FU+MP9ZBXmp+Snot0tK6UlYXvJCBdk
bbYIX7yuJ7nylPkQ/9LfmWVzp1Z8UsLUngkYz1Cz/ftbw3COfjUvANQvPZfRgRmw
B0mr04O1PV7yx1eyuwk5iP/XRBetMWWFN1dcuUQoE6X+LvIegAZStV72UlR7n/2/
Qkzmiv0cDh0vEO9I3CCnxTQ7dY9IRR5NZcUVSizK7tFPKzThV9d57mBI9tVA1p1c
9YTBZJ6kDuCWvppEgSlAPzwtx4xhc8X0NmJs0225K3qu/CGPCp9cXtMdj1xSf88Z
moFP4R/5Z6ADSJHg3b93Q3ZBmcbow69lxz5ii39W1TeL/d1FlaK5pOFHFW1ra07l
Fs3rLin6ZFVDTWWxdLJ8YA0tIDWBUoVOr44H8oNe7PcY7gNPX7jvP32j2EOLrRvl
OCckc0+1ICBmIX0ddI9WJZMK55YjGs8v1Sftni6fCn/AKC1OL/ZZY2SHJyKGoL7s
FOtMQcQwOHCEts14hQWicX5XaS5vsA1JTaqsNgmv0WgheB9QqNrNEaCkP4sh2DT8
cVYbMC5CTQ8iOIgziOJ0ooJGOHo4SmBVeOX7mrUOg67OVBd6G7sSv1usnoSZarZR
biXxsngNkosPpvtnt3eHXB3EvmKMa1vE0wMhuygOA1em3Hmv7uzFi8fydKXuCPhn
yuvmt43ILYY7JIljBy8RAiyE9i6+ekRnb0YOq610872uacpDPcrkEwSGhVQKQIbZ
aX5u3JasFgS09MemugjbIjZ1DhfiQViLqCMA3jGzjyaQh0ZYb6o517G2A4KCGRe7
yX0gY8qXL4siKmEuS4/82yd3OE2AG/+IOi7+El1muYTyBMUJECTzJD0SKKTJEKYY
v9vqrrUQihJKCrKrxHVkBPU8F9/bZ5O0E+nLecd9Qxu9JyBQxnhANH6aPJqxzD6Y
S1+7DMDbjzR/LEJ/wEGuM6LatoRhyyJmPKZqUeQxWtuep9iydf6rI11jWB17C8TF
MRsT9jPtTcBYgbCtc+CpQIbxJKHJ2EbP9ZsUMvMqKDPvN73aXZny5dsJlOuwu5Py
xisZdOu28MVZf8vdNooigamupWv802/f535Efz+v0dGCPPQbIRRS2pGB5Quc8Ui7
h5Dl27Bk2Adc/77DJ/v2s4cQGyNkfqI3fOPNXwdhe4D1dgmaF7g7/PPq0klfG5CW
CW2FUs3xshZ4gl3MKYBzbD4kUqQyBbbcMoedteSxjxaO2t6XWn/nVpdo/CI3Vfyo
6b8Cs1E+6ROzDgbDQN3FOdTfaxAfbQpooVwiXmGS7OjvEFdzGm27efCyoT+2JV8+
HR+jMaCrQfGIJHtz6W7IUy+BahYUw6seSaVMHrdGUkDvIZCYapQmegwCIZQGDZEn
NqoXXvog+jM2G7dLHXrKBoBYXHnZCJZIg+gD9+CJMRsttW5fdnvA2s2nktSknddu
aPGjuGr7uO1Cckn+kafuJx1tPs0bOhfyGSZcy+oqip7MyEjUWLsuu4ONEGWMBTZN
zhy61/eyjKXZGxEwDcnOP9q2npnda60iv7wki2PlGsUnryOZg4F/1vK/FKKfadYH
eYvtGaEwAfBGLyx1NWrKgBxu06+fY8sXR0FlEA246J8VT8qiK6NkD95uxwgtexgG
YumTuRtdjGwcSEJJlNRmxJeStRCCZ5ZSmfx9nKhWDD0w13/wqlBogoR4ngu4yCMn
WM6BFPz5epLYqryogstczgwVOdAWHhjxSz11I/IqjapwmH5egLzi7X+ALVPedOMG
RZUuq+WWZnh6AoKNDZzXaJkaB21dW6VwDmUf78obC2Wnz4Mj9EtpsZ9NmWjcgw7O
2kEpZDYw32HEU2oPXtongfYVA4w7u1Ch5LCzS08Mmk6P6+QJA+ABgi7YfvYy36Zo
RKpZfI/FTeHHLScLupiUyEDYdOiRR+5zQqoGnxwG9ByQYxCEDjIgfLhr6Gk8E0xi
dxvRu41sEpZhAOzGCwLBj71iawG67s5dNQ8GiZNzLeOpfa8B1MSyxwgaA2Ir8qpT
iG567Ga6yojEPfMygwO1Ak0WcVinhD9dSGoxHmu4d6/gGEAtJrGecKzY6MuqgT1I
pOpeE+LaQWeiqAKtt2XwHrR3zJOHxaVOgChOJgH6sOHtdfcaaefxU2c4C7xDn0AG
EyT4XsOTCvAd9mqFZ/Ndw74Sv3OMeDSdEUzQoREuypb/F+6WSqQ1TjRavepajoWt
r07g/aHEnYCOmdjZozZriAAKPDHo4DPIJBlVkyKA7AbsTFbu54ialN1K4IOoeHGh
KrYfeQoAZyLWB6V4hOt1zzCGLhSryggu2l654vs7R6urcOiQ9ZNrw7D0lay2fUx7
wJX48Yn8/2Fs9yOJl1XlBGfsBYdHPFF1m+fCAD/k1v4gDTcdsYLelauPXJfuQmGO
Ctg9VFpthlfNm7g4+7Dc5DbiSlVLkQvE8av1Ai9FlM7FNOALxF+SnjesI4EYEmqn
UymNvO9cqMcIR9DCI1bcfhQXDudi71jTIa3qvzuxtc9QqkMJeMEB38UqZgWIxROf
uzgWmzpe3EIQz2rMlpQDyEmAHV0JRJs8EK8LF+ZfGxnT5UssOAkT2bplhZFQ1lsB
nVjfRhGCJ3xZZL2k3LQ6v3su+FJDR6hvb5W/GxJY8+ZtVk+LE0pAX9ktUoZ9Z9GX
yUirWW5erb+y2hq5A0RVmSZN7yo1bxmdQOW9UfuYj2QV8AdriVwBLPmySd6xnOBK
b1HPlY0s1fmwThVrVotbyNdqkVj4q+6gtVemsadrhOXWXuDlLrmmNP2hXVxSKIuW
2gI80EVSQOS8o0W9/WSSjy1DQzQGfefIhHu/4A3VqLTUFJ9+aQv+gHqfIvpJzwO0
aVNle8VZ0LkYUNRO5raY10kCK/e4afl6JTeDQh4BoVSclb4nM4k+WaYP1DEcsD2w
JSX9qcJuWLBX+2HY72c4qxkv2X0YE0PswH4yqslcjVudwti1W1bFehthrC1LKvMo
Xh53AH9S6ocnASkgAd4f5SUuE8ugfpZkxFhmevakOcgXfUr5STYGebcfLX++O9+X
MfQktL50Jwh/kHqzy27tDcCAzCX+EL1zVsGQKN3cQepi/dlqGhOuKGDC9UT2nB1D
sfqs5Lill+5F2eApEjwhqWMQsVpqTOAX4X6qvLnYVUQPBpE+aaMGbYfRdRR2Pn65
7Bj8dmyeg5eIudIudXvD0N16eEK3jIvSHyPPpI4R2w0aId/R6AFg2Yk/FW407Gk7
V8sUVlvIhc12VMRflbD9f2Xy9fg7ABwwLVXdW6OrHuytibfR7r3oCm0d2yS+j9JX
3DEpuWcQ4stNfswfbLiUbiEgJXmUmd38UTBpwekhH+jRQVgOmR1Wgjkq57Pm5+3y
2aiv6JPD7L9HQjo0PIeMecbstyjf7KhFNDXuF6P5Kdo6HbRyDWszWbm9FJtZaCyt
wO2GZZnxrPWylHGf+O52hIh7/mIYuoi5iBnIPgdpQewrbTA8NprqzJWCDA6DZXEr
NIkH7kKCfkLEq3RJ8ppsa+Wv2QN40ODE/UV+uUz08c561Am6MKR44p4yOamddUxy
C9ObuO0d7Bxr+AxCe0Ke7Z/kykBQWH7RAy7wz9Y/CsYPYXu7WkEjUQdlyEf7fouX
mmq9+udAdx1O+9ZAbPB/XK0FCxxy04zC5rxUYLXmzw0P9FzQkrYbbrHSuxUGowGj
MhWOo3xNuO7a5gQatN3GOIbuVhbNonGFDm5FGrePqTXVSfHxp7JwZI9dp6B9V/fX
yYXewcYTFiV8MuHqO8BDMEz2nKZRLOXMhnY9MXj35viuLED9zFQTp9Ngh9KMjM5C
JNzFiNwmmFgmseRb1+3UEzTWkZ8ya688g5NmqMhbJF27Gms2Up7RGaotHgud9RJX
ZtbOR5w9/xoiD69s8928/g10OiEyrjrTsbwYHrXNlBstWpl5c2LY4+Tpcu6DtWob
k2NBHMEY8fpXDsIDYtyDP9vEk2G31xIakzQ1cxz6K6bm0EoBxbs2aUyGhGr411+L
2LUhhZpwyYaMtP3GdvthY3sCrxuIpxUAqIxMvjN/pSpViK22UqXtwN/T3ka/v0nK
6eAsRntR8IegUg9I841HNoYYX4ImI4SB8Vro3N9Si1HjUWzfp2fQTiR9Ust7enoX
ILLmxw1e1o8gOf1WFkaZwzR5rQGXQJwbor+TmJwusmMs71qLDX/eRBeg/iJRLyZP
mql0dVJQcNC8Rz8bVYTrphya7PTG5wnx0IQ1rP6inFUMvnG34+bSHbMP/TQiqJ3d
NcwOPhK80AHWNTCQ8DkdSOEwMCIC38dmhPP41pKaFkuzRvYZWdyXaAa37aFiyRkx
TTcZks0mkHN2QfLwycEZ2H6VVimYffBbPaOOGeMPp9OOnjmtB5rCoST6IWvHHKVm
0rHx62A4zWL1qCBuZuBwsfpukPE4rR4Ho0mDdcxmy1/YNGZsrz8ZJfJQotLxAUeG
Ievpd++x9vN6MPZTyk9lAEvYvNtefl+djZFbqGHEa6P6X6r/OCDEKlR/Gu0TqQHj
BSXFnxw65lEeuKXmsCc2QhcwMvWf/nvuay0jpzNajQr2Tye89hOw8H/5G02J1QBS
g8/NrooThsHTISorZy96hY9IfbNpyXqz2ag6EykDA2sbJRqwDz7hvrX9TQ2WK5As
ra9aUTXUQ1TTiDEs0/SR50vc2GFUS/9iz5HmMcHaC18pMymfFQfiikNcjiALctIj
ca1AP/1QllcW/aAx6qOgUpji6M+e+qWV00lRrpDmXmIh1pYG6SWyaTWTnSAzYW/K
zHb483OUUZHOxzSfV76Uknf9ZTeqXTlQS3fxzAbOiyb2uKsLSJ2cMfeMmmzZf3XI
hJobLBNLHqQDFHU7Pfk2vwZLeL4ObJdqAxPDzeDbLlokuVCoXUe0pN2jfSN7RF5q
bqkhToaCWMMgk7pw2wo5dzqHNmV/TmEdH03Mg0+EY67DlQckrbYa4R++hC3qSlSP
epHnJzSpsdM0pQ1Re62HPf2JIi+1Lrd1sYkQ/A6dnG468CUpTM3cKu1O6CGYSxOk
AnRCXWnD3gQn/mrwqQwcCt5MRwV2sBcrHhVDnqVFL8c5iKZRZjArtXwQRCL5B75d
Tu7DVPlT3jD8JWgADK721WQnG2S61Em3lshE0vXsvjyoHNqJxWjx4WTGKNB2iygU
UwVoWUXw9kXPCtvGLMwiGFIlRlwyecVkZUCgQscoTd9tFWAvLsdPDL+hWNq8Zjzh
/vOQn29sqEzEeCGvuyvLm59JFIU+D3z0+GtJQQHLaKk3RPsit4aw4UkbgHDEMIfN
AGYOscsAo4uyRygf1ecntH+rNdDkDvnOe/R05Rn24x0gWeDoaisKT0EjamHr5N6W
tDNsfIhxX0u/Dl2rOXF3epdPOxzq0AIoGRf9KFfN36vcb3dA5bcY01FdwthnNC0S
oYi0RekmHxjVhaoAnWNkje7mtGBQjKHfE7PJmKp0JjNPUtcZtkU5VhCzIfGtN3jJ
BxVulgvldjmqJHoejVoud4iTqO4NfLZow3+vJWzv0A7yNoSBC+6WBBoBq/C8vn9c
Ua4oXcMLXuGYYMWCwrk2FCmlJcO3s0Yabi7jYJkXkbtr7yIUrfBaATCCWAHzBh+H
UFwG7/eqMFsWtC6MZwGsNcGOPYvCk+68RaY5zaFToOiFTRvT7XoJkdqmrWb2WBKg
ptLCF2tSsN2YHAeS1ulIcslCZUmBOo0Nx/KbEVUG9GOMjHbymMDagY3LhxvMP/9U
ZroXGJHimHCOpJQKxow2wsgu/l5yKpULynN/BR51D5ote0dU0h9KN3zU1xYiVU/t
gwku0txXXqUDgkMmYUQHR2SPDI2Xai18L+h8lc9N7dv5vLSOH6CER2LA+Mgtt6xs
hyLDVUaxtDe8qr+t8jmpkRVu59Ij4PN5tt+6lnQaZJOwZJPqFf00jte97EajaPDN
49Ar/cWcVr/tr4zjJ6NtKfNxQ+Pk0lUGr1mCcVRdNhvf/mGlA6dyCIQuAuWm67ms
6p2+bQRq9ZRzA+4T7G9saTrd/hbXOuxriV2LeaLjNsRGQ3xW7+lPEc3zItrQNMVR
edINKKT18mdZPEGdw+Wq54z0ZUimfZcd+3jf+xhJzC1l+gX8WHhviVXhlXMy9S5y
xSul5TdgLauWAA+b1La2CicXXM5SYJ2BnPrE+AgmootJ8BsLhqYAIK+VhBLr8NuZ
73Dgxi1yvFkmtX30mxcGN+Rif3SUw+6nZ0xFnp3AgEhYqJcNW7Ho1HuejEfim/jT
i94GaE9FYVz3CULgmBZwChIch4vo7TjTeN+9FrX+DkfcJ+WmYPonW8GrDMKgf0aO
pLXlr8VM7OZB7F9RIz/Tr0aXxcObgrQovIfEPhAlY+6PS7Qm+P5NPYltIrIytC7G
JAh6Di0aKQr0tHT3s8UFf55GUHT7If7N5jnq3mmay2M+Nt7mCoLyrqKA5/1/m5F0
sjwOB/vDoqKCT3oYAPQfuHf+Yt/XvYPOwhwmkkKgV2GN9AJvChA7xfToCducpyQM
BnPBraJqZDVPFVMMypwqOiiBpPtvjw3utx1Nh9C8c/6IkYC+DTbvx9Hq9uD/dsUF
TlSKPD/Hbyb7pKsWSYFttk4u/RgKOBK07ZyzRE02FJ/jc8otGU1ccAgCxpRNnRnT
Y5A4UzIxfM9ZaE1HL0t/qmz5KVFYH3dbt7rY7cgxo9Fu/FRCO8U9r3UYgqMDhGuz
NQnnG/U5aOmANo3ol8pTb7qTgj7psJ358K+5nEZJ9iK8Zk30R6So/RGGlW/SZu6k
ftxsCCF1sSrNQvRETEkkPUvA76FlKz24OlK8kAetyhKYvM2resV1iyYXHlLagtL9
SMDEn6n0YaSNLeTg8SAFUG/mK2ee779xeCbUfdrNg9CEN9KINnfkXLHSbFOkC/+R
d/BijJZaeiTKIgP2YNHXuvHQ5uxBbQJ0G7Qbx0DdEPd3HzDJ+IpPvUqHUpM/sn9x
YUmqKENw7rZQO3Acnmudc/bP/GlGVQJnbiYhcjHyOzDXg/X7J2nfmcnQXaqLT71U
cg4s9hj5ckSKLNbec6UMj0N8qf90T+xMFcfwLf41kfdYWKXuU5KEdx81648FEMgM
Dwr62j8kVyMstgnVxuffcCGSh63fbPO83a2KZl3T//Bfcp7nwBFRo3WkMtMGnHVE
uSPdiL+LqtFA9LsyXNIet+IW5W9/sAvp+2PhBOlLXdMz0Qy2FitXFkW0wu22+gI9
Av3XMUf5zJANelYbKmrOyNRqaDcgwBrd7FqOA+flwFmt9CaJghHpjXdzGcd/VRA0
zy43Bj0e7bQBveoOYSKMtBhkJR2liZmqpe8nkLh1jSlfWcP2V99lEK4fe5S8maXz
gQoIS1zv5DF6lLolcGizLELR6QF2DBWezUtqY9opU0C2DFFPsHfLspBpoKvISVwD
IlBx292TE3qRZ9PgowPZiz96B4S9KUZGJ5UHHRajTO+s7pHhvzfLhk/MUwg8YOzo
dUnMaIvBvGSJvMT+vuSfVc3c3uAqXpY3rdjk/i7JRMy8DXX0BxWlnqAUNjS9oL22
mmMZBYMOf2iJLhZ+eATLZyWKXL+hUdV4TzxJZrt82lVMUChi3d3MFRvCHLbZoklO
hTsyFmPBiG1aq/Ecz9I/JqJgeJWd4H93kWuIOjYLBqzu4ur+oSDIKmbdJXJX2K0/
fO8hTxZCbxLY/JliGx76wg4kRVj4EJ9lyqmSvfiw+1IPuQNA/gTRLmxooM0imQEG
dIDSd6XUSIHjVuuZU99zfQWJuwVRaqXmHYkO552fLiFo5UscLOiL31JhW/b5p+kE
BIrqpjUUB3OtDSAVCRUHyEMpYuvouNT0nJmhAXnPdMAshp74by82l/Kb+eMAMzjJ
acsbT/BUDZGQ9qEmlEjfLms1peA/wG5ICOa8YrxD8kwDgqyPdjVQ9gGRCx3R0b++
DAYnkeCXi7KIn3ifbxjLlikkycxi+I57W6l4ZuM0ssoKG8eUdIN7nee8ceofCFR9
67QKv/TSwrVoiNi/6IAPSEfG3H26OsKjWpNGPD1QrbKp/Op6iyiQPoK08ar+a5eK
o4rOG6jdaV4HP4V8v+I1obMGoc0qWktwc4wDFGaDZKmzHdeCowapWS2tJxGHU81I
W2gJ6HOaJFz7JK2Km74wwOT+/h/pBT0gE99XTNJj8I9CaC6bn7qb4dYQxFuOS3r8
dxjhh/Isl8/r27HZOwwQY0gBV9sKZ/euAVOJ+Wc/HzlfzjZj9ongtFu/GbEwOGzU
pu0EcbyYNRoOkW8CuDrJdYzWGMwpBmcOQr+DWAbRaiojuxfZLQj/2IJgQsg31dKk
6cYlQngxCXaB1hEqxt2khzR9KRXtkShlJqwRxWQoDFe0a9bGQ11GvV3s3Z5Ad1aj
K2k8ixqai164S4XaIUNz57EddxGNuHjvwpLAtsDl9drsYNVpR8G1gdk76E4s7cHO
FzUm/FdjryrHlOLLwW3uiLr1EI+r39H6gN2JQjEybo0J5LGwCSt+0WnK8OlFi8cb
E2w97JiwQg6P322LuvNMXnAVqARE39F+wsTYL/HygakMs3zXFrE/NE0IRWukjM98
FSbb19GVCIERbf+7xN4tf49WyTsbGjryh9rF8fSJu17sWQ81969DBEfV7V/af5IP
MyBkahKYhDpuT25ycvX6ooTmQjBMiMIN68ZOuwYDtFsFbGcoOklEZ0d8kT7009UR
rlO76gMAxEH3sw1UcNHXVFEA2ZYseB8ac2uQhEkonqbcg2+7vh3SOHrJL/wmJ1QA
9WSh6BTHwNgaNMi+4zmmjpHBKvbA6OT2CgEKOTy9TUQebddBST03ZwHVJiHCljWg
kvcHt9exkmXPPhX3qnIrrM6HY2YPPG9f8j+pyMDCHQVBwdRFY6MKqce8clIsfz4s
CZq29uBhVBesmrcf3x3TqYBYuqD+S8d8iu9oipj0dyF6YLVSOu3RIno0NVwguOPu
JA/8FiTHZj7aQNCGoF9U3DvRNwFelACpOQ7zFFXBjMGwjJnp4FeVzzHqV3UX9j43
VOCj7EVX89CTzRlUDsNYJS/7brothKmFCOg50RDoetNa3rP6drrdBGtIbZv62muD
qkYLr3aQ3CkTLn5ZJ2ArnydoHAKPDjkNxza/mGbAeh16LcZZnMY2pE682gM9waIM
zjfgS9s4SYaeL62cF14aJmvy3GwUZrDCyzOVkdI636eyBCJx8pdMPWYjv/bk2XZV
LFOaucQu5A8LpeDrT7AoaFSpmHZWPdn8c+AN9zLhEXI96/l27eeiwA/9HVgoF2lX
+iB42+JyFyZY+zf2vJJpe8x+HtT9oA5cTlgH86fdfFR2HCMsAKUdFnrZ0kyGcEk/
A0DiaII0kKdzSCfz/R9GgDxiFoeYPlT1LDfhzTg/wQ0v7ojV4RWoQDeZMynn9KpV
VtZ1EAeTiR5qW9v9Mvjc21FGlMQq/Mrdr9inK4mcP4Ka28NoKxm2jqHftNNcZsiC
UPmklPcPJDoqxHSmLXeKyPJCOjWEm003UD2+WcyW0OYv4VF4Q7TzspOnB1icKkbl
PoE9jA3aIpEIggo5LlVVrTqoPVXwSsAlJq4Cs6MeKjPjCQ/1Ia5maZrh5gxIu3cJ
hbFJHc63Y6Eph9//dVyGBOo7uT+XdM+7OOsA5QoJSOG5UQhNdiYxDwcW4eZF8p8q
f0xTPJqtvTVfr+gNlfuoEYR7MKQzbFxCqlMrnrReGWuBPcT+y6R7lYtQDF56yCWx
FDdNFePS2eY0PqpFkSM/VPI8//Rpjrli1yN2F9/o4RtzC+zf/MjIAcKVmpYW3h1I
/GvkbBQrsDtmi8ae/QX1ValsR8bdUukhYNxu2daj3PcYCX4ZUQdq6sB74uvetpMM
cm81Xzm9ZnrIlJMxS8oS3sNHifyeNrohoxY4m3nFAQt3Cd17MtVg9f+kOBezYpaL
8ZJXmufQhLpgA1GyjMRKpV3HYEZ0suJSJEW/xTQRsD/EISTqYhYDVbHh+0dbWaAr
IU3gxCGopw8IHNw7YOdT//1Ga8CE8crqqX+PBDAxBOZYUyzCIxtF+GK0oKzbTi0n
9d93cvtpBOEk4xoUFSTtZMFL39whhOg8o52rM/Mw9m8aoHXIkO1XW/rqDl32xjIC
NeGgHzaXEYDxxWBpUgpOhPtC7J5hfk88uloiwcGPVQKynqyrZYgcVl1T9S12gukx
s+J8VqafYbhkNhyo6lQ2lluK09bSG4cO60I0skHy4VMx3pQVd4OSfBh3FzdyWnb3
Z7XQHLW1Ozpen1L6e7sS6+R8Gg9TynRGCM9EUOrotB5xFbqYQOkOV0lpRYM4YAJo
h25OBuDNwK+yFR3LzwyGLcaXlCGtJe+UPGmz8V1ZU3FPhMdqKXjJgMej2J8zGu2b
eoRY6pFlzmp7lIBxQTWQ17hfGyJu6SM5Is+RpYi3LtRYwJZwJAwQ6F9LumOyWRWp
xMV7r+Zh74Kamb1TjrOurbk240DYD0UVY0E056RZDm53q5FT2KkP699y8Crrb4Mq
9IdHEKzirysEg7BZzuz2pPeMmI8Td4fBvOjg0lk9JHtk04I/rszV2op6yqE0c4kd
AdwPrbcTIDXi9ATWz9/C+sp1KIX0kN35TfBCllAHq8R5Wv/flcLB8iUvLEkBV1dW
BPF+3kG/WIfwtC0NxFkLtxh0X9+Jq3QVzcd/5Z/HlYEq4XzPq9TbTpFgtbZMGxKb
a1caWpjDp9TPZjg1035NLJ8wsg/QJHQiwEasJZqHOJU/o4OL6QdJnR2p0M6+LB6p
988E8IeOmHzw1a7/RdKXyHGNzWx/0f4VtGH+k5agwvdwFkhh/Iq/h3Yue5j0dcYz
DKjx+1UX3JXAKQ/UL/cgPJq1VC3lASxcXwVVfFhK345ODPoR9wDaSIJOeajK1uwZ
p7TBPJI/rSSfCSPv92ZmHSg2ZM0WyYBtYdu+WzGHJcqsQmUHW2Bap5SsHQbSFCHF
HN+k4EBwxiau29QCl8BJD1N3t710+rjVw+CojSZmt6U1wco90ChS2b46ySCmq83o
3Z7kxEuwoxk9UDgzw6sZPI7jTcNirfWRlfEMN4OzL/0c3qd9Gk8MoTt0ZMRxV3c9
3tIFhmjnq9tmyjaE6ZTczLZwfUopsdGVYi4/WMrgH9IN3xHC6ikOOryoiDtJPN0K
YZ2KmUpQUKYb/TscUkDwslhf/qtLxCOgrPz5IJMbP8ENmJtfq2Ql/VxwSwAewFuI
KBzNneL2OWHg7yE2v9vQI3flKkfnKJZkB0JsoRCMlXVxNgKItkz9MgiJOhC1BdwH
+2N1Rs69W5zPtN5WXwM6AfDsZWvhwQFLwavdQoSNgilJcgns7pmlG5GCSC38XpLy
ei9LXIH4A41aktSP22EXewzibuAlCWygU3MqWz3FysxNklj+G/FU3p3EaZfwzxOu
e1zUp3ZbgG3ldNo0zH/SdsxKq+0svQHDUc5w7JDvwY2Ax3kiwky2MxLvQ+bdZhXg
PZ4GPBEHEFhnDRShith9h//Yu4+Xh7WRk25NkhOjgpzXQk8mMVSo5tGTOzkwYyRG
FWF3yrR1CVFME6ONrRxLj3FrSCSvOtROsas+tWUvd9LLoXyXy/b6sriI/GSaf3Eb
HdF0FDjGKJxvxMaXBzwSldSZN4P1jhjr17nUqUCcp3qVQLxgpq3zlPoetCkD4Jjt
tjb3Lo8jj3or9gxN8DTOhG3Pf7PUNvJ3RcbPoHbwUJG+Ev/WR+pAEdFqhpQlval+
URarHAmPWal3ebeZt2RKSVUb1kIrScKfl1HuttLjuTsTQgv0jQtMB0S2tx2e9S+n
+RVW45Dp/vCX8LpIFNY5hXt8nmeV0L4TNWKp+TciknlHASJSszY8XO0ZEQxUXeP6
cXLNU4IKM6vWblrbUbn0lyLmcTWKbL5Mtnn5Dh6ZMt0O2pomE2/KVRVMxR/LGNlm
99WiYPNHB4zfLtHtrnAx4S1ToxsU2IUAiRF83LtX4s0b69wXth6OhUIHMpRreIiw
vjMOQzRm2FuSMdTmTy9KTQiTS+PsvFKmU6In5kNCaLwE2dDEQHv1htEu8n9gDxRt
DUpxQ6OBGdFtOtfv/LY/IfsySuRk/WolRYlrghSeDSY6QQO1bowqGiBnht4TH6ZS
o64UFNj9IIT23KtuTtLi4S99+z6UftAsx1ErENO3DVwE2ald91TNVpFhNFay+MW/
0y13e/1Avp4VmVCbn4KNBWgT7g9wABXywKmvnG/pqL5PR4uHBj5Ma/wfP1esTnJr
diX/WP/m9r9l6VxUKkFGQzNT+sXDF2DrW1bvMVssMKcu8xR8LF/LonhwCRiKowIS
UhhW3yzo9UYJU89ky62+LQYCWcLF69HlOe6GCBYcSstOXUSmx00t1apSnu4tgIZ6
rKTnuoOoRdi4OSuap/nCdpfrDCqJWvAFcVl4OvfF5RdXr6uEOGs88ybrJ/cyhBSq
MEO43rzlD/O61Oyl4/aP9IAiHUrgMghn12smu+OdSjjS5Gcp9aGf0FSutZfqr1kr
KE+LTJn/cSMnRpLxirauDDm+XZQ+U/PI60m27S7PX41qewsFAYC5lm2wswkBrgSq
mAozIFSyjrLKP/xeD3TiVDLmVNsTblYg51ZMITirZCFm7wGTJXtpd5a5XeFFxxED
vdjyhwaKRxKXDIAT78Riaf2KaC4pUZJa0l7izBuGEzoVRnXMVFZPUW+6Bik2irr4
hGreInD4e2pM6rBx44M9knSpqccbhiRN0wsV50xmX5mNCAQZdWgrHkegpz341FPn
NjXK6nvi/Mp6pA0ZKbl4hs8unvSq8q43+QZdsydoTD3h9/AkQjEcNx+5aAg1/ZmZ
lfgLxlFtbQbSk3i7wKrYz6fP45r2hqao1RWf240qiQh5v9VKteWOvJwROKkRunOf
Kzzd+CDH4ybg0vL+xDFe46Sba5N24LFwdoH7IqbIxTxY2ivLP3BJ4nqkCKOTdXbN
HO18F3dwIYnWCEfboaTfp5wMehJpPhI1cXGFMFyDF5aeSbjKpRn5D0wCkLA6Th/e
dM9/1VW4U1XOycwAFuamRJYC72JLsGNwqUmKaoQsc/mnIEHTnbo+/TxAPNaerQ/v
ykytNt2zi5lSG2Yp/3Ll6qyFpXq1CAgxIjmG6GdsOnfG9LKVWQ2TD0Xqb/32+Bku
K4HKAUS+k/wchvz/6oNiqLiFiSRHO08cEHWVbLj65lMPBe3bpS5LoniljuRmdky5
pbiXE0mFJeaWmDiItK7e3FOnUcO93qprkUOlv11i7dTmmcPL1eFL2mVIEpuU4jGp
z8lMWtru970p3fxa8aA5Ry4RNRth4TwM8+w9pHl4i7WsZjGyxSHaRNNRqhg6mCFZ
cQgz7+0ZOd1f08wqaLkQ9sEFM7U8q53lyCyxEk+eYbYY+cLCgT/ggHIwWRtCWie6
iME8uJhhMt1PWXbJnE8Cm3mnMPdaftnVUOBOn/rAdZsjfXHdahUtyLIsyCkslBEF
NPe7S+aOkO1soSeJutypa601HIysQuQl4n1bNFMeuc2WeAPb0WmcY/n++F96qVSm
7cmZQN/0/TXVlHL9/INmV+/41QjcF2zup+6X0Q0WVSL/F9g4e3fXI/WtYyFlyou+
krNf8OPyQb9QgL2xswaOB4bx+rTY0eyQ88crMbmz2oWbpCeDJaQ3VDGtmUt8s1bK
ghkRT8K7ZmjUQXEQAdoW6zMQXVQtZYTz6lzJfYugwpXRC0aR+AZgn4DCnHWSn/4k
TU89YE5ZXmves16PYvVu48lFt8UD3NmmHA3Rk2VCxf3ULYgGZtDkS+BToe0SnRDG
H1Nmi5EsG+iHl3QUrKh+w/Q/JljA61pllaq3rXrXVKFxmO34lk2ZVw2Am4k3yxeE
2z9TWrhPFaLg/5d9bVCYnoOGuwqxKGvoVlQ+RnngVEN85oNTZ6G/wBOczv57qF9x
x4pQl2HzqV7C1fpslg+Z30UtiL34xgzbFsGNZOpTyESAF5W10yYZJG4Fuml5JoJU
ZiCynb8QcZIQStzZgXd9/zxY8KQdb5s3udEUR2r+y8+EpPNZbzvOWFWEsCrfaiRD
8opFLjfvNn5d9OD7n59SeCMa3wvrNUO3q5mN8vg3JlRb1OyPrEkZ/HpqlOPhNLiO
31g/0EthdqQX36Q9b650SltT/YyFDNIzmpKUpLijq7j9Jnbw2wIYh7MJqq6QfOu2
/adlrtJ8xLMeSuzgpjFpdAUiBCpU5NhzXufx1/A5TMJFSoH8jkT9+63Uj7LH20E2
MqaPY7k9sBNeOBEemGYEEtC4K7fHyg/koV8SX3kS4XDUR7paPgqZ8IjBOd2y9pqN
y5BNWPaRujjWf8k9Vw92Sd4MssLEIDSm91u4F+78bN24f4pGeDjuZQZjSyKy3OXC
xdtqOaIhXa+iueikG8+ykymcZqvH5J1i1hwtohnrkKtvEa4UfU27sme3e6iLtRa4
fvj90+V7DpZmb/ll3GP4nRluIcoFdSD4PPQ/vjZ1GzSTOQZiuQcvbvODs7x+HkN7
HDFwtXHj/U2urXJUV9XC8yaMtxzQG4Qibvt3ItQ24Dl1CTEnz3Qouw/IphT7JEAH
aa5J+ZIpvjv9NIt0acSKGs/XIfiPwL2vU1ft10G86TZFkK1eg2g/DvqlGaqRC9IY
znjzpsaHiTfg/EMaLMsI9e36PVEKIdkhBg60+VASM11X3xcKUZFEz/6F7SZu+8Mk
WIj3V7kjYc2fk7wx2N+2u6+b0YlDOIZId6AhbbFmIq0uks2DvM+BYuukQl+DNM5N
95zqGMtqSwt8a+i8Sl7v4aS7CP1lWUeA34b9YBqB/rGsLj4DntdCMjKypSsQjMJT
bvePP/BiQnZxqXAY9LY0dZ0/+JF944gvq9KUq9mFRYtYK0UUs1uGKugSHZho7teN
EZF6fHCi5gF1tvFnFvXGlexusx5ZVmJZsP182LWyD6EGyM0SvDHAbiLCao2HjiLz
2FHICtLEBKyEAn4scxlg4x6/2O7txcGv1n54aZJmsAuypLvXAiNj1Lx2MV6K4Ad8
Dxy4zDlOPxcDSiLOUBFSIAunY/7dLEs4F/qWtIHlLyIDmYcG9nzIL29WSGHehm5L
4GLnDo9Z5u1b1t5V+TsKplEXjZRdSzRrlCI7qjF9ig/gZe7WavH0VGWdomCvvrGn
Xh193kxm2uXQvyr4Qw6Vxeggb1x1eWM57zjZnjvtU+XJwVY1FDvVClksQONvK/0O
Ta5BG902wrUpLShhfGMUTIlmat6gMU3kqCEksBghMUmtA3KHBPfjEsCk3rDzZULU
1BPDzwwuJ2t9KJTXAzFozPJjkYI6NDxGLwnmzEcz2TBIGgT2bPfO3NRFhnyemcOT
HHVeOXmyFXmUr7w1jb2aSrlINw2PNw+O4Sp8cioBayU28Zl3UgqpDD39SwpN+UyW
yB7VTAFs1KiVjQN0HOKxs3zfdcSMBawRzH+PtxYsiGLip/nSSaCspWqdPS/zg/yr
eD1AUntDxEITpyMHReJK6RqczS6nVV1EokvyhcqdRNokZT24kpu701+ljp0h1Shm
WYKtwpja5CjgmNTHUptDqaFouE4x4coG6whrPpWMSnric/KWxQjP+ihAADO5LYAw
mzuZgpblmhL4U2QJMp1z9lpSH8lQS1FpCg6ZeTkBEDAlnyDZW0g7vgNi4QIaNcjD
4Oy3mGxrQhmvWz8ojFbUxwPpn3TOpYEcdIFbUR8bk1czt6KQuOEcxUcg7upRJpoN
tNnUEMRDVPmSgMI/g+oatW70EM/KUtSRx29bmJS4yimdV4qp7cUV88Usf8oobAiJ
Cy7LQ33rYjJRK76XXKepTW6laLLISFnK/7NkiBLsGsrWRLuFwSpw5d+3ZMiyeoS8
UnNmgUYUQZf+c2aWSER+TLIa97OcMTfL5skeWC/OR8o7CRAojVLUCPuwUDhVqrOZ
9jJ6odGyitj2W1NpHY8jGbXXM9BjrQyCyb+zN++Qsz8Ge9uJ/eFqh3+2a9xYwSxk
TLAEHhF6Oi7if765dbX1rgDe3iAvKf33FR6FQ1m1JAvhiklS/JJ3IzcDwaaRUwZT
Z7i8srS62evKnFclMgEiPw9JeSZN31yei/CZdT+N/Bh46LRQaUCWV1mrJ7e1Xhws
EjSlczhzZT00vRau9ZEgx9xPOmZr/nfu/QuZrX6mCpPQXTRhAUzvb/fbVeO8cfO2
yz+ONgw/dBrwaH57qwWuo/rGFBGkcUZULt+JxKUTESL7fcYGHYFexgFaUINJQfVb
UNTcWn4D0MJKGg3jyiJunkw2L7w2daSnx97tDBOL5C8z6v8qkT0Q3S4CIkmpLi/s
YSqdu+pIUymQXIdI+QUCN/JaRC0FUIfvjmWIeg8RpkEGZ9zOcLkzUWYXihw9VdXD
eM7P6LsC89CAHkl7rfLvE1zvZUF2hAaxlw6b/wt4cp5o2QthlQS1LHX5Q5ErfWsi
kigGYWvaeVepdzZhaQkrReCiudshLFWMFXijIqc5w75f6Ji70KMmraN8DWs1pWT+
Vk6Z102372KEc7C4B0drVK6ZrYr1PP4YqnmCgBBcsS23X1itxCU8hPtOVFmWux98
FDsoOOdX8rOMC+mkNmByllOGWg7SbndjAqiV5Z1R1J1Iet9MERv7aLJf6HkEIFwM
+suhp3M/66bIt6eFKix2drl8apWl9k9SIIf7HPBmwgtYCBNpBuXLBtABy16Jvf+c
a4WAzfe7ZF2sG64WbDCzLCtqPHjr5RnFhqu4mvvv/Q3+DFPyo6YxnNdEX27UdISA
lEXtX7oA5Qe838HvdpmJX8aUS6LAHTmvpPc5Go9fBcmDiY/Nbbl+JyirbHW6fwkX
MwDtExPgUKeXyGtH+7sLsM5FArr5x4EaBTmobmX0y+nwpr3IpapPXLEBBI8VeI9Q
2+UPIWFvO4zLd7M4Vu+8Irk8+L/Qnz60vjd2hx+yFjIqKsYh4fJ9Y4LLUWnASzxO
OXgZx7WOX1e7EHO0PxtsktqZNcTDOiJOelVnIjrG2ki5iNuePU6P/kic7ICr6sKF
lcZgJOWfcDZitbj18gsKssKYPwFAJEdJgfWIwvvHiOM0RcRb7xAH4qVTskjVmgFE
lZ06stzX3wtwPGP6OZxBOsjYAm3A1tuEOEW6PemQuI0WIls6nvz6idUEfD96zuXl
5xu0lbOyA9f0yylUGrDkrYKnBH3HCMzLHUHLxfZNTGS+WKsQEzUeP/8md43Cg4Q+
qHcXOmdf8nUIOmRBPzUCNF8vOvcBuOfOnCB5BvEGcMh0z0upsIYKKE7SvhFMGa3J
2+WVxZ8ch3cHyYPSoIkILyNKyl0/s95ieVjEehNSAvtlvOaVMFxN/uhJX5tX1hoe
Qu+PR29subnCol/OJRwbC4/lDVeopSaw3BbrKUu2bxcr/rKuaSDgq83cDiHc1UHO
pg+LAsb0QMF+G0zLn6lTeTDKvOH2t9EYP5H2qiO5xzGOsKL/j1pZVuYwaohL6UxU
IG6ITlTtj8oIFZ7JjbKjUZZxmsQ4HuCndcWEYtvC3dViCLFydxTs9EL3tXrOy4Lq
CG78WmA5XlQuB1+prc/UF1mTDj8c4M/xKeMrxxKOdcqPYn2vySsmmeXbrx1kKNag
kg32kbYFH94ySAx2aKlONbKSCkJklD3quGweWNZJ754F7rHpNdhn5CewZdeCj3WT
kCiVKdEqhre6zQSA6DbC2BA9p+gogpbfb1j5SJr9eTmiBNinOD253KNBPOMG5Ihr
y+2GfhK6v/TuxyD9F1q/jPppv5JIt6gG9e6aHNI/Y39f7bFIpAvW6oFHkmfUZJcf
00ty10mJf5O7uz8T5SruWVb9LH8NK73Qh3hVcUa8O86gCR22rqqj3E/d4yO24Bjf
eGNh2CdyPrlH1OEOaCK6OKbdP2mboiywe6tiUwvQbUTMEO5kd6csiuINcVZPmKrf
zTUVumozbMK6Kylwk+eX58rhv2izsGc2QKXlgnjLW2qChdN/LJA8g+TgmcId8gEC
L5GOQforXELq+3GkOiwJnkLmsRmEZBIySynvDKkG5y0uIk8GT6tiaicU6khuDkRI
OQQOz7GTO7nQT7w9ly6zUPBxjIWMmcACrsKZPljls8NKPxSHFfmLAnlXnX4u0A/t
ctpbl/7PusFbUys9ubPy5rTwg5nTQdbZNcAN7LYxkT0wsQdPRVCfeSnlqZLbU/8u
6JPKZ6zjr9LHyeivF6BFkf143MEQpJzr2ajUwUFAajVXHYdvZOH5IaoHfTB1Mrka
BxfSMIBPZmdAcBk54XSXBzrUmvm7p5K+BIAZe8IoXpbqpZLccek5kkfurgLf+XtU
81cGBB0FA+brDlIsiPR/URqt9M/9j3OxQxQaxab1DpcBPh+gTkLBgvqyXsWfzXv7
z/V5ILT7BPDk7VnhgKSCXbDvjT+UjSnGaL/D2Lb9spyYbRbFr/vsUVeMNV7uaamA
b16FsCMLAOnFrVbjNV+pyQVXjK4T8tHqqtvYYr94lxCQM7opRRkYzzmsiPE52bAR
xsKnnFL9yu0lW+LfXcyzqYnvQO+3j11cREKZAyaiLUU3HBRlU/s228fxp2Qvss5U
WrR9yyeWrTF/+TYDY3tzdMeaXLtx7RYN5hTXAUEOMh+IFtbOksWk0utyHl1Dn1bZ
i2JJ/uVDePmoYPaHJrULSrIkPb6prvy7Fve85ydBJqAayZp2zA58+BqTwSC4SCvv
oKnFQi3d5RYcLMe+W3y7Rxxotw/bsiHj9Ul+8HrCN8mD9OuGfoTxikzyTjpzzWOZ
Is4T0QIbqXu5GZ3Jv0mZAluFz1oRupAa91rYVKop7Ii+f2HrD+1w21VQf+AyayKo
sIdcvnPvZMFL3BUuecTDYB7whbJ1W84ccTZngu31SpHPEGm3AKm+UUP0EzzWIQtt
uKRWLYMmD4ywo8iReK6FZ77u1dlyDXpyMEOWmL1Fw+vUwPNY9cGSx3Fn65ouksC1
R8+3gVvYIlYZk8CSUX5Bqvb9sxeiTkM7VZS1slpZ6nykVPkCZRXlFyqY/RiwncRd
yPH3Y7dntmE3tK+hrAkRcUoeU18YDzt4bH8pS2obkCg1SsADBGHI99BqELenbzKa
5r4kBaGW/m8P6e4G/mNMgNeHpxVEhQiQ486J+PeTXpfY9N/gcfxuyGjnBUUssCz6
MWmdHloByWv1tG8zsdwVXi5HS4as2/F28Zm+YbUasF7Bu7Zlc+WHoKs1dEkjPfCk
EfX7pMWroC3Xar2QLREVSHgGtMfY95qq6mklzyw5JwlqzfyujI/qEZFCuvz2E1kj
dUI8epnAR3h4AEenPcrDyiC7r2SIbfrI40pNrAK8wjE2Ud+deNk4n3McMjvJHiHy
/5Hs/RQ4FFtexawT1tkpzHqi1K46XxAJea9+SQXwBbTzkLOHLUlZkty+yRGgAiFZ
2RX2OJRzNHom4JUv8nxfLAcsP8q6UNkmEsF/lW2UXj1Vm9zGg4kp/x1Rlyw0GW73
JAwaHFaHhijyAUH1TmNvpuMxxx1+WbHycZbVVoYSXkY7FAdpBjpc5yGCZ+trXxzj
ELC2dJkvaf0BIKoO2hrm+Z5f7HGKiO+hTD5bRNukr4mTsCb2lKi3qK4XJRFPNLh3
DUkt7W4LDtcnfaFoQKnCwxgStrmS6Jy+24+YK/g4VM5cWWLNarnM7DO5xUqv2EAG
WCNfSpM4bErxSR/OlYfr7XAPiyle2dfP0CHty7fuB/CnwOkikWv1rDU8+5qmzD3C
rluq3MP+RAmpJMpn7MYsUvL3IyJjoRE2ufbqBKpOfMODV7epfhlR8/7RaGA1Wfa1
88kROGocSypjayNceFXgTwnCzeKUeNM684glDJZAMM6LSuLGrg7dxljANBCLG3LT
cnHaDsBekaCMd4fK6i10xmiy73suXCTAWHDpCeAhSvGYLbrMg10u8U0kIQzZ8xhv
6/vKMkdwXHGViJfUm8X5V12uZZjGfNtk6BmJf02tYC3DdE7AXByTpPUaqFr37oJO
KcPqZbgplHS9QF3AG25sVznXP++k5mi85ZG0xax0ACqepJ/QH8m+JvlKOa1Rm4sp
pwGzZ8n98HYDgqu7UxMLP28pFzaemZf6CfdAKz0ORTNpC9Tf0v0xuJ8sgqvenJcP
MfFbGWCXjHxTnhUnuVIH9CzST54kII+T3tjG7vYX6Cg8dvCUCEEGQhw5UxUHAu8D
0+feW88QZqVTOykZ0k1XqKWUk2P3E7HVWqiWQpbggxVRRvMQLv7CrYEXKSDYLuUB
9hgmUVEM7Y7tQnbGDtOgoLT/Ux87BSaTMDjt+fkElO0xyp0gGvU8r0uymehbxVYX
x8PsyANN1Km9R+tu4f7Z1M8+J+YT/Ooo/c648iZE3IKshIgDOvutDvpg8ltz05IB
L44aujogRI4CoYyaIb2VUbRdi2VvKwkZ9DLi1oOqwwOSyrqH02qmPu1dejoKdPDj
4EAxudZrRKGaXHXEz0UvjyYN0UQyidflCwurYUm5Y/ZNFFLGwS7Ik1AL1d7MjFfn
MVCASFESIPbSV7AGffWuqQngTd12jGwuotFM+fow0nsLkDgKFgiyFS7JdMXHqBXc
OG0HB8ApD11KqRZgCSNDSF+k6k5ZdnL+4TaSKEeIVdKiQ93RcFWSyKmJl7Br5FC+
zoUC1lFKD5COo9aOgmAafHpgxQ1Wh81v7/45r5hJ8KFk0rAj9QLnIRcLgYzNuJxM
hxi5iBCqiR7WczSV0iv2RImGB+RAsPNVO26Iifx3UEwF3SfgseLW8RPWCs9lK6rv
zDs3KCmnM2B5Y2xgInVsTH6UV8gbIFo2uQ0ITffFNoFP/pY4VpRZm/hxgHWhv/Fw
2mJwWPUadJbUFIHX771rOzraJei1YFRT7EqJtnr+P2KZMu7pQfdjMe5vilplOxd2
Ak26QkGNd3u9nr3bXMty3wziJ7xAQRHtrawkfArFK24GNRhQHsf6zIzgz4Q+QQO/
hXoiJDuy5gx3LLxjW090ZogMhcIRop+xzRC4aH7Sk0+nzBvs68d9o5h5qzLxgKxu
loaW6Vf17BB+SJCoFHRz9lpEyJvI3C6VuisBvYS+oJ3T442kC78FyVnTA7AQz4OX
u6mAzRVECQNXp3UpHnKOZvw54gIsGdBHE9wGsviLVpJt92fe6HhSXBNIc0+UeVwG
lBOdUClBWB8T0EgHlTTmJhWQJZoxMJirvbZsGfWOUIuS1/cTh13ivblHJ1u1OZB1
ebbb/HgvhSG2ngl+R9NHJ01j5wRoqxiDYhhARCL2YMQvpgbGdUBLnquROJdGq5D7
R76HipV5koC9cIUGb3mtxFwOY+TkVncOpxNOllA0Q5G4FTuXxC/MChGX4IpHQupK
ZFdU4L/eHTgJjCW24IbzNwuJkHM7z9iWQMiz/5kD2o4/qbzgk2Lhh2/OPbGjGY4C
/bYl+6fSLB0KZ3zd44UitLPNYqCXhxKVKKXjblmR9rvw2NVLaNrQVB+FbpvpDBjg
OJJwcCi0Xq5acgiKTdke9AWoVW/tuhSPvcNY6yfF6durIPyRgJAZ6TYbtPb++R/X
+9+q0VOlvWm70yZTKLIz8gq0h5E4p2a/lpSy3gm9pyNOFb4NYvMl6ghsN0/dhZ3d
j34UVeAPD4GzMhwSNNevHAUgkDX/rqfYceNN6UmalWrGT+SxMR+oxMBJf30KcrXR
REMuxRmtozy2gJrpEsfvon8XvDxSBX4tF+vx1C7Kjnkf56RQJja4h6t8D4/X0VeZ
1poI/Z5NgGm6MTcdCgU13L8enkkCkh54xxbmdOB4D5bPOo9kw/2DFG/RN69IFEDH
TB+Ifp3Ms8zn/p/mTqAfObCVI0OL54CtD5aS14OgHI6KMKXyOtYrKyjOZYqQxkDG
6X10D5ISq+lFtCzxCU1cOcGnGPYpXGP235A+fL1G5HU/UfrMeem1MjFcUckFgVQT
H/DkwH+nk/ibp2GF/NVChi8CzZQBFq9TwFxqXMdXQIUuu3158equ7iSQvHJhOTDA
PMXHo+OojtEZtn2NVlkZbqz2I7AWpzBjIwMccOl+qc4Uk5ara16WqHWTKLZXsWUG
Ll6wV/yNJgCt2gnvqOnOQNofwf164miAi9GKP7VL2rQ3y62QBzKvYmrDgBKa9ra1
NN2I3yigQH9ZhdmoQ3AJQZF6hACwDPn20YYlwR/rqZqq5flBLvut5wO+yVWfu25Q
Ngh6OlcT6ZAd6SsuidLuPBW5UGwX491HjrAnSaRikuxNKVTQjugjkDsLkQ/UyReA
KSPp+9JUaxYWqE8/euQyW3F21xxBke8zex3gYNDQRHCeKQ6+z3l9O3ef9UtW0TFF
8OrvJQPYa68I7ss1Bil+MiiuB5uxVUXPKgOHNeMgXbYVgujqHz3yD8yJQq4yoSSD
MvCzc9L3qP2YpW1oQPUkagWmRxUOhWWV6cU6ICNMmiSdR+icvMX0XOlQgfojqLh7
CYcjTK/6aEtr5wqrtlYVsedNKUHxYU5gEBqB1G71cw2pIIl8G8jDxMk4Bem8YaBF
dDShjN7HqIdm/fYufNZ3GfcC4xVGQeSJBXqLwawm79Bik2v7a9nHLT4BmJQuIVI4
K3SRlkXXJ8Ggzzt8BdlNqdyEuC4TV0EqwijdSqnXWZdaGn+TmHeXtXB7pQzpyBfP
31YtEn54hmadafoQ6jGxB/J4ow5iASEwQ7fgPNq01tB/yBy8C36S4H4+xO6e4FcR
OlVlNHRr9VAnuGXX1nlVCsTMYQ9IQut9AdC0lIDr9VhZvGcZMmJUrH7bA1edWK3x
AiQO48kCHkY9sw2i0WcixSi70RMhAvEyTneAJYh/krId2k4Cix+iO35jKKVIeuet
sJb9pvBjumS3T6TICDDQVM/+CIm1d+Wx824550opkfLon9wFRIV7lXe/xK55GAGY
i13VW27ZXD5XulP4AyLYrDQALdwYZrrkpRhI7seZ4npl8ysQo5WuSC/QhjHrJiGa
a/lanEOsfWRQ4US5JGB0HOxl1bTKs2fNusQA2pmVQnKq7Og+VDQwt121DzEBCDhT
dhgkLGHKbiaP8sjj8qxKus3hyv3fSJjJXV0GsJJoot2ZCbxnB56AtHeFWJepUNVa
Zd+5MRJ2Scl2VOmtD59HlgZbilnceqjCT8UQaNC877ljC+wTgasfegH9nXeQstNk
wTSXAu6EHIbEZWHdu+vHKxH+tE41ja2f0qc1tj7LT3C+hqGmzXjdmjUvmWEFtg0n
uN6dSfVSYGZFWc4EHOoTjvlaML+PAxYPvB2uzeOMAN3OaLM80KrgbYdRfbmG6hj2
s8ytWmdTIBIzN4czPlXJg04+u56hwNjoDkWW/s1fiLQRgvzFJe5X/TZImSsJ3d3b
YSpQvszfEmv7XMSKhJhy6r1XNPm8TvSQXGHWHLcDX+PnL8ojqmhieraJ619u3UnB
dOI8/XcF9/5s5bddG6pWUPbDlbWOYOU+YxqxyqYzaPvr5NiYacyO27OHH+P/j+0m
YMGztkd7pF8uqrDAMxHsF89XBVaR/Z7INSPRPx4eg0h/Qa75k6iAZt/5AoFgOuUA
ldXt2XZtSQTF/3QM21KTYPXhToVZihLaRNT7zdfdDdB5+afRm+oenYKoji0seZfA
dc0RDI2WA8mnSz4wqP/HEVQb3Ogpmvpyp2KSZLE3LuOKb2EHuHEI8N71sqTP60UG
NsPdyapybdcHLL+Unz1cU3zZcz9nBbWPfzE+wZ0lJuB0hXZt0zfyH//ZBcLyY8JH
WIc5HQN+YMfbJgxY5am+B9wbntg0ZPFW8a7VdiKUGLy1ETm5t0Cp3IbOOaHG/1h8
oNpQD5bo4KmTvHE+SMZ2PgFIIB3wupMi4tMc7VvNwxEVkH+z5eQGz/lKzyJG0qKl
Pcv4IA6DCHPRcAruw3yfWXCSQmBoLuuJvYtmZZTHaRaoolX9PZDKQLn+DzrbRlb3
XMNo/heTuRLoLHTI6xrWwux3sxdeUZ//6RNLwiDh2ZuAZ+6xSIiBymWDp7sf6zGs
5A4p/5nqYyYZL1baXKVdnw9Th1IgIvvnvomjgXKfphGTHXcGfNptgJJkr4liuxoV
o5Wrd0/ValSxHCw2AocLMTMB1/yW3AQ4VbaINfzhaiFNMhmt4cflLGWUy9iUKMZm
GblX7WxQ9AxqNaySFqUiFsLmvP7FU4hT6EB4wY2H1zKzse+elUACmz5XUyNyMKUk
iFqSB+vGykn9B74iYfUJZGKvrruirUN6vPJR0fFVCNI7n8R1zOHEDS+/8hxdkddM
BHf7hoWODuWs3O7EtrZcO8D6ZyKR9eqbXX+q9Xjh5izaajDrJu+RKU2zKpZwIhe2
AtcxqUAFpV4jSbKSltGjQwCnjBa2DnIeiaU5x3SjfXblq/gNVzh1u5VmEb9RyeI+
aZ+q6eeu1+XQ/Lp23QD4NDEzCysZ2HQXlgil9h6axNKrZ8UnTyygaf9XoX29yLbz
APVvaeGCExmDeLOn7qSm888BVjvFRzE6D2WT2fgR/UJUFJ3sj2g0WBE4BUqax/pn
FRGXllIE0+N+7AJs/i+Mt2YRX0144d0X0ui5AzxtbKZbAPMD0dRV8qn5xVjmrvMB
MrQ5WuNQT0vgMEycOV9DDT/jOFVgqj2RP0fOYKXXgxc4t6NjQnet2Ec4S4rrl359
fC8slXiC1wZsBTyQWXkdAxncRLfpjCDCzee5r+qKMu4sycAEZZAOasRGGjZJI85h
fqFpWlSS2FLrKWi11bPn1FXXA6pgcLXfYl5fJ7QxeHraFRf+BPjHuaAN1bruDlC9
x3+AM3X5ABlkPqyeSvBukTRQPDjjW/ZpOEG+WCWCRKSAsnmXaxOyl0rw+TOBCIAP
zg6zP8drqBOu9l3m6m4Ka1HfJfd85Y/b+A5Tk/bL4vx2ekTyOvJwo7kPTT4fhC+5
bBm25zQo0fif6Uqlzbp85slKtKtY1TAP7r+IxGSDw0/soUDxfv8+wQvCf2ZsX44T
zmY7rox4eeUVeWLFHP+Vx6ijV7iyZJ87do/xJymFdJ80Q7Hm33AqzJjJj8bc/dW+
b6ccX3LXpz4FNaM0oQRLxH3SGl/CmvcF8fZcYV14gibDzsMB7iWgcn/WzQ21i0tD
x6PtEAHkbdBd7iRWIclnpV5wHJPNDS6/g7Tvn9yagP6kX+UAwcopa3iGXc095cx3
Hz9tyguN8CmiEJzRCLCJ7o1TUzFxkpR6ddMCjnL3VGq9gOGozXI3pfoKHcHxm/x0
DTUPWDDe4U+M6pq0uZR1W/YCaFLqt7xwVAetEBiIh1X7KPDwMPCP5w0/jDjBGLLu
63bhi5hCW8IjloVgERnlNU1rJ6AUqfOrDjIj+O0thh7p0i8aA8P87CPtpaaF19Xl
HdVNnzj6qFRgM08vnHhxCvQWx8zH71s1cKolFlmyZLvN6nhAF67ZcyPQvSVMPGT9
PDyZD7hdrnsuzV6mIzFtFtPkiOt8LuBsmap+zBkowFyeic1WNlYAwq4rVwcvjoUf
mBY2qziwMj1sreflXCjpGq53aB33YYW8wgnn2RqA/VdbSCBX8qPLTFrtU3tM1SCV
kdIFcRUgSfGGnyh/CvezkcL6L4TmJtf3Y8HCNkrDbIwjRMWUDKCzIN5ahKYjCKXh
Z7x9zzG1Byls6L+1+kDfLp2tyNwPZEHU83k/D/JUYB8xy66gEUbBqms5Jh6iozzf
BpCnMCYm81/jcvprLXsSH1iSOjYYh8MPMNcArpC0vITYbrTwBnuHRPwNh6Quzi42
0QUQHRgc4jDhP5wRGJ/XppOvw1UDM7qwU1mT6tf0pFTSsoinnmifW+Po1L+5s7FH
YyEFx/nVG9c23cC1VQIuJRLn12U03Ymts8Y/8n2GgJBO/Z3kvcOgKFKxFRMHUaI2
gEPdkNrZq11SCPuEU3jbdB8TdrcJzl0tgsTLx+cs7v9YkT0GQF2FpP0RsIKaGtdc
s/t2HJJwyZzZXuNAk1s5HPg8EVZQv+lpxtEaK/AVfEL/SGmrIPVRzpyDvMMj1n9U
WOlg93eSgvcANya/4OXBAqGyst3thbp+V4wT4BujsGILMolCkDYcIRFx9OI8Oifh
ZgfX7yRW4HMEuDr3i/cllrD8vU9qURkqmvYmN9OFTY47waV9EChqN1jtygKiGvkZ
MRvaF7LoYiwR70H3X4NWXalyLY/9zio13AexPR70/tryVdn77ej1F+gR+4EgRs4i
kjfmFlQL0mlY/Sn5wHli5mVrIL2qnbnuLLFRXlcFXxkmzlbE+ioHmPGn2OG/xDxK
jwe2snsCNjfz4Qa+D3/ifjJQ0qMTQULT1iYlR1RKWiSG3x5MocHWJV5tDPraMrYg
KoWLWMe40i8Vip7ZzajHgTug1A0xukcQmGeW10OlYGR4ttrbNkXZPcdCVmiJ5mry
+FXTDRpbPMaNUA8SqldaKcC3Crd5M2zlLh8s/BATBoNiKEX2ZnQYuKWmWr+mX/dW
ROJ3eWjIA1qkeWqFX5bMZnEJrrhhsfpJ7S7zNpEI2QGRmvtsTWfZ0ZPUJvD27tN8
zvMG75YAvA5b6QRQKXWpV95vUHkRFGK6H/NvUVsN5d36Hz6/EIO3Dtigq1eQYgDP
+ZSA3iZB9YFAkQ4KhqSmiHhoFnK6MDjlAfWjy3sT1McC2SUGeeRfyCUcv2JBOwlz
+tE3SYl3vXiFUmAO42/5755oc8b2lwBFemBM67oWTlnML05L1WaAVV+0BGcBz88+
wXVZhGOYcvNaIasJNXQhkCs8Ui9ZkJ+JLNyf8MMYtbpG3qoznFZNuS76fFGP5usu
gmvmA4Dtiv3RoRTCmLLLgEK6L3sOQHzss70IAY/I7d8E/+RaPUKXfcgynPfb/7Oe
AoHUzE5XVL0IeKE4dgG55gQcw1661XEzdSNGO3+LFZSW6hP3vfEmwX5QG7E49iiV
yIlIptcTbcAgThuBTyEKpUTSp0N1/qUIb4wKbEJ9yYDzpHGEUOWKsK2bnK7GSZQE
mtv3QxZHRABYyZWIOGgk794vZx6kTfKxdc9Pftf0+qRz8BY1fO3RdfsnJFKNY0eb
6ueOvpGB99jI5RKhfUjaO2RZ/KV4W7P/mbZ3lOaX+Q2aw6CTTr5FhYN4oYw8G/1B
k8IZpA/GxhffTsAr+4v2RTrqlnIaLOjERYcuMhUFKehXHUohHWHBWDipZbXXctP8
LnMOnWtE141LbufOwrnS+y2hNGh+wGHxCnN2VdD9tOPP+8vO9qTdF+ASmyuYkuWP
pn+jExxHfZ9lZhIDqFrvKLeVynxqFV3LYOxXItAVeI0S0hDzcuCyxJGn/PIiurIv
tqDlLFzll4YgQzJUlvSCrUXrM4zp8w02xYZfKLVs//Hmn81cGtXwwGkyfya2OPrg
7BDnYaU/7pzxVoI+mZCZFM5HB2tvhMz3IA2ksyDsDIQrYocN4DkO1u0SfeVB8MRK
ImoJbo+VLO+bH7LBtm0HosZteJhDhg1z3hYZ01xobnvZ6kbFA1tkxQHxEFI1gPyJ
ozufebOZnsOXqZ98cKTUnoWG/o+x95PAKbcmOtdr5eV0fC3uEizAAkXFFPk2CtWQ
ZG0b/JeOSrFmu3KHiazTNTv8hF1EA3LfYX7P6r0MeYg/C1w8WuTzU0AVNNnuJ6fg
mw4bbR4h/zrTTGEWneksYjE1I1NXxD1dxdPAwaWTt3akRRRdAxiZeJPXRMuczZf2
8HP+DT8sxXfwEkiPEZcC3RtW5X+mYKK284Jie2Ni+58LFz1FVV6nr00nLCGj+V+f
pS7Jm4qahQm0uaJIbeJnIJLcW7YsJs2wWP2anXXzA55T61XafVAKb15NG5SMPx8o
rrRZIjADxiO7yoVZ9tUgvHTS4DDUGg+zlf/3uhfFYZoPdPhj0aInyBKKcn4dK0I2
JXet3CVL1AQ5ehF2OdEWqtkwz32RTdoLqSvtFvvg71U8r7H+sFtJYhUOGwNazBBL
romxzf3EQPZiDZsVoDwcrsOjydUHibL+uyrLd8IhM0pe2tJ2DsdxVU0hvaFUjY4x
fW604TFQhein1+ECLUTFIN4hZhFtHFXY7B8OrMCULj2PtNA2SHx1+6gtionYoWS1
v69uAEtR9mt7oa8EdiGVX7Fpt9o1N8e/o4B//kvyLPAsxuZuI8kcUU4SBM6aflmU
53aeS75qXOm3BFJ8VXT2irsDd/oQRau+i+KbXU9k9GMbD08A5zCRXCH+FTHzXVl+
fzv1yiK+J3rUnoo7UaOx8wrCdo3nXVq1hhhTz2CBdgPw4/M7shJowAfxB90bHIU0
bXGQdgIVnL7D7RRboffS8E+JO3vFsHAGMY4FbP1vxSa7fDF8HloD39QhusNHT4nK
apzmfMY9cU8AsyeRscqK7wH1r2yqFCvx0AdzcJrnr6tKL5NvidmdFzTVLmO9eHVO
GyxqnWEQCbJWey4GgVedtf2z7vUuKPKuyPgsh1mjzonaz5pTolahtxuUEHFA8IR8
9GRs7z43rw7S7ft9GLbWkuISMpdadhgVTbYXnCRmrzIDVdgpu3ifT38yvwGyW+Si
jmBKQdxRBv1iq0ymeZiFFqhWNjQ5HFN0k2i/kWHxaLo+Zg3GqVH31LVcfQICfD64
uzIgfcJb7xwNUYp/At6l2umY/wTgXc9pgx1ZdRH0qg3A3cP/E+G1jxTbvOsei+J3
CfID1T7THo/WUIKEU5IS4PM2W1VYtZ7yTI0xtP6VXplBou1cNVDrXJBIn1pCFOnx
SPRARBldPfpbP/xeEeBeGJSlISWtUXqSpv/QOB53Owl626TxA+iKW9yfG0axHefS
xaZMyxP9EEB+AGin0Tf9M759WFx7Z7Gep9a1NJ1taWmtRR7mDRgNQCDUClAdUeej
f5KgT9avSxuaSDh2xvHnArI1LIPE2iER0ZpEbGA1+fBgz5xwAUuNphhOsaY9eRaq
TbbOcT6umiH+6a37Jkedp6v87lq6J2WdkDGtolfU1jFXkCOdUMQ/MOo+IdIqR1HG
l7heVNbOk/4W0ImzL4tdY3CbeU8+0bAZlwGbB5J+wLM2PrDN+yNB4569ESUde5rD
2n79Cz/9aLhdZRG7G6f2AGtIZ70japZys7SPmnFYNk+REpAJh6QrAkaXJOy+vHUe
y5Hm0BnPOjmr2xwZgTOKBB5ZRm2IJsjYJBLqIxvcVNTx1eTx5PmsffDBcYXuMLnD
cOtR6Gaz6D3lW3jYIWBf68XISuFN6QlAmbdGl2xzOifoXpA6nYOy3XlblIL4Jmyv
s7FvDk7Q2lYyB8VjJD919rEz6esee8f5SQ2w7kXo0IZDyJhm6ZVK1OvmmtjmPDGd
is7+edSm0vb3c+nXi8YlHSEVq2BCY91D4ReJIKNJeB0orfg+x9J4hHIr2GcKK00R
uh/ka2JbHkJeknsttBWL6afJ38RnRh174OGn3xUpT01+UJxxArCh0dB/ip268xyV
kzir/cbZ5QUNUOxPguIbI+HqabV3O7G9/QlgNX84BqUKA4Qxx13021yOseQtelKW
MR3F7IL2dZo215+j2Nh8wGOmTNQRl9ufIx0XCB7r7X+em6hN4PBi3lNARwXTSeMT
RDrJT7Khgcrvy1E3qEoOs8AJk9G/qClgRLYl15UvFJ3/PlyfO352HqipcC7F9coZ
YdG0AtSYiX64LnEsojHLxoc3DN8lwURIXHI4wy6uDU/hfcyqWr40ljnuMSeHQda6
7r8BBHDOvlGxYsRZxZYXxLRuOR8Bs4cfI9vnG+VgiNBqksNZoPqZKpPe9CUd56um
J+z5qXNVZW+0PIglhw0SCwW219+9YY4oz14dMumRxCbWCSAEBtHRnmOJvsPHDxS8
HU8SA7psEpVB2rgu4OzXM1m3Ijh4r8Lvxn/Miu4d1Imkl/FIuWLvT8HcFCNaGCAs
jJxyp7XHkNrULf6LvIvTKjoNB7AHeja2Xo4WPVI9xPhyFDgFubHLp3fRDldkb8KB
eDFncPDaYMC/TLa9ZRYuJ9Fl4hKHoG0J7U7MbuJTxZAY/cbzBClXQFGgcQfHRoLv
Ghaa/uyhe2RxuxUBOnya34b0mjlHYikkliPLUMzdtRmPR2bWuYmgpSn8A+XCq7SZ
DTm4EQRtb236XTzuvPNbEQ0e45dZoid7Jvk6pu2KuncgsXt5ulpbVW2wCEc+wqhh
TSDMUGvsU4WzjsigzlF8ctdzG4EZ+ljamNq1Nlh624yBE6qBz0Gs6HcaWyqRJSiZ
w0abTnP67ulkKCmWUI8Q12TsQdruHstA1dVMlD5QCYld3YlJhhRPqReSeH63rRKv
ECCWhKGsTzusKAips/0UWbaMDyWXyMCwLrgX5HAXYvXhjI8FKJLga0INcB/9ORVF
xzisESFl9jzOdLikgPKCXpMlOnVPqEovZYpRBWRYAznIiI19qNudnZUo7EU1uPsT
B2xeqiM2tmyFLqS42AQ81ACP25OOxQBVXwaPpzO0tLOYbIgTe0idXKMqNfmhEdP8
3d4DbVA6ef6gM72E4poi4mQwOmAOGOV3wadBCPJJiJQwBXYbJ6zJ6uuomgQe4OLj
e9RBr0jj1JpX9eqqDBhe9g20Pl1alAa7TKWAHcO3r6pWYIPet9/thXIzV7X42nyX
v+1do2O55HmeOuhjURDeO3vl50IZcLsn0G+QrthUjyAXbMoDcQDkXC9OC+62e93c
p+GwfMVLied7t60NFT2B/LkN8oh6CIPlXVjRfClGUcrS/nEEjIt+JijzsuoXIFFM
E5TX/jlF9PdSrFlR0eonNCGmgR8uZX7wWrpwC/RR16APS8HfklX2VGwSWWpGR92I
w5u7rGzLAynzUVJFUfSDpO1Bh+axtT+bn2emRyqSxBGBY6uluh761fyOdLIMEp/T
BGL1BhnLb2m2kwtjHDvf2uTSQhYBzwYaMR4kJYplObDU4JDrgjZDvHr5WRhTDuto
cUmWDiw1qY7+xZNJpUQ/29iskqR5i5Iqtf/mdTTj+M+isB47hK8LdR/+CWhbAkll
sCyUTU2yUiUouSo5MkUnBrfpxNa0MbmIRicAEp+aUtjBoXJhXhp8S2oRdKbExugi
P5tGP2jllZqzumNAgkQZvj8uqkFJGUFAqKeY7UhtJzrC3iPa8P1fyuCgU46i5ypR
yORA/TOwAzOKhLlMuwjKW28T9rd7qW+5LilShH5UcnF/BPj6l9ACVWu5ji/2bsIL
4t1AQy4EPENnfmWvbVwks5Yt8bSP+gtidsc6f3k2heWfSaDWnal6PEEgdglgzThm
8b9KfXuaMXt5VofTQFHVelaPl4JJJoB1ibnNXAomMgRW5MSunVtCCFLzeiS+ZduS
g9AX6pfpmhzDoxnhBmtZjF1eX8e3/gGI8g50AYgq441+CRZn+KOCkyYXWdXg6hIZ
HF3SY8XJh8DTIn27Keo5wIeaj+RjjqStONbWagvIWdJ3HcU7sorSBEad3TsB1n4k
/D25QlsFQgpFlOEcLR/vuwJhPhQFpExIGwRWZ+P50OWPFci3oBFfH6zxeT2YIfO5
OBLYeQt7UhX8Q3j67uKLYRE4drbb5PIXW9Mqk/AOCSD+4QJw29zkAVKfLN3jQMWc
6UpdY+4DDE2tcU4dSyZ7hAmrMAvc/Wn5vwF4cCDxsKxlPUjk3EYKeXjUNT3QJbV8
mpE24vyEdRPKKRWSbCY0LdKEdjowCahuXlUvY+MRM/V9PGAm803gNBBzBNX5PqSU
QTEaOMv6K0wPWFgayN+mIdfAWAL6etmolOA91YG+hzHMZNwB1NVKvde0LcL6SoFe
Y6JRA14OluUBkvE2Uggy7WvZQ8mvu9Ywe9K3F+OGnGGBGaDbPA/tfU9i5GJm0TFM
bmwryadACXRV5C2kLxA2/356YFm6FyWEvSm1+4AhdITnUHu2T9Uced5YvfKLpDND
Iw2Sr2wcH+SpmhGHYrPYtwvIwLi99kZ5ee/4jKZClXD3P97n5ra05covl1itwUDs
WsDnFq7fnw/B9D27eHnWW2P8DHVBoV+gX94KiVdavLhZVrjmXG0okUzjDgwyJsit
fN53QlMncYxl6YbGkgWqG301Izd3lQ9oviirVjOx1UqBd7NK+4o8VyafGPV1wNQg
/rba7d05g0shQ1njPUQXPG6b5Uo1wZh/CM9s6oygkAaUVtOkd3LIsOwOk+OtBScw
n9Go7tmq1yZebvUrhTns7JRY1/Ji4+jlcyrk3+McUNE1/MBQAxlGD9uXsZVU8Iem
p4UTrLA7ML2T79EWujd/+rwJEObE0QJK4rphTb3EKeWUT6llffwz7PIQCp2F+US+
fyd/f8ABA452KqHXpTLFW1MKgoGUOrMDGbT1DoSBZKC29UPUVLV1zDAaLrMdk98t
xTeGDnGmfh8kw4ZGg/GyZREyPuD3p8CnnkVtgzYAee65Rc7iNr6l27dfJvUakYOM
S7Jf5GtjcBY1fVJx48i+tfXst40h5tfLOlHxSW8aanGneTZSnDOY/D9QoHlMVwMo
r0xXURO5o79mq3lnGA5dP+xnWOd4jBkjv0Ag5RJOfHtgvYBslZjCrPaqGxSWJ6gd
s65L/GC7LZiCSau+pQ0PuphU8NGnebgWob0oF+aQ5AefGBzKp3YlTgf8sqRVpDtb
rWqPPkzHWDA/oql0HXlj7qDlfVm0Rwgn7IOk0cDMYGoKWGrEO1nKfQBEH9fwH51L
Z2APXZ2BUQ5v6NB/aodc4XddFkW8jnY6d8Bx2A1aisAWDVzk4SmSqomhNUNJ5TFn
+g+Vmq1P6KWUNK0a7uH43oUZMfcRptfgZHneIc51izjrE9heVJuD8qB245jWJDEA
zXvItczz8nPPWLTdXL84Rm7c6dGzKIAha7bVXntCfHsdSsqJmyuAkqwBuXfiTqry
1Li31EaFhMin6I9+zldy6cZGom/t08mwWyT2uECCZu1M/SOKxPTxywrOtC0BiMUK
MSAs/7Vr83NnydqSY4yUCIMQpVEcgxD3hEQximLzoSq7dyw8PhwOF/ZP850h3/bv
8XYZS7ZBy5FWn+NXU9WnaiSCThYopvsQlL7/Rqrjv0rXorMzrrhynSpLRcdvnW+B
4SGrlNRQvyg8b9Weqg4hCOG1YwUDXecy7tMxi0X2w2MQhG9MW9h/DZ9cS26FpH20
hbxejwP2kzWVOORBAe8sjTv1Krg5Ra1mxucpqJ+kawthKlcVC10faN7E8KYDE72g
7xS7ezaJbLuZOvMPzSieDPmIM66kvFGc93XYuDPZGN5Tmseo1y+qgj8v1D3IRxDr
b9U1T8/nUBRrAywQ29XV+T1TJNk259xZo3qBq1yoh6EqEI2fSeLMFvdrrenDs87n
Mrnh9GediJ92UjMMshAyMft00x1OaIH3x5b9nXENcgEkHF4WYEz6prgQ2WR0LCvo
0i6LG4w/Rgff60gzhJGfB+/O32wYiURrab/2p7pfgCxiRf+tP9l15y91r2+j0L0H
4MvqUCrhFfUje95hXRayoAIxOCZ8jmvbbOPsXMsZkczBCg8xemlh5KgtNv5IlaN/
wcTZCAMjTymiYs2wiwSYF1fOspXBDHqZtTkn1DXqDnNiAj/PHwHv38QFFmjt3bcU
2NB2jQjkvyhE6ccnRdMUQjYp5JqJugXJ4i3AqHmbtuRWbmqnUSBtSpRm7ykMC/o8
8TurS/mDa7CjqWGkDvuF9r+SFr/GlLXLyGovqtcNAmB1CbStp11TFFw0cVU5TMg4
+gMYk0RSIDXJRn5Udo34QG4qseuzTqxmnS7B5tuGMQlLSH2+v2u+i8jIbAx9DXHS
HPCh+hVqiubStoqSLl/TqTpowojrNIw8xibLFnv0cIs3O72i46Ef+ZxyYxQwa+MQ
11oQjs8Hzkx3nWcfid+LxsRJpzlvvezGVql8wwl1Ok1rUqGmq5x7IbjMdrMbDAjb
jmNwRdm3iXFY+Qfb7aSgb7TpknjuKBZEBiPrSrLY0Stjee1ckxNdAgdK4cS1kNCr
wwBycwIz119CN35MJBAICZwT7QiJv2RUq2HM5COykcnbu+oXBkabuQbOusS0a5iz
aKTheZt8muZeqH9iqSZYuLisGB5bcL/+SYNJMXsWXrbpmjspM5LTHN+jj8i8jl8P
0yzCPadlMqL+9Jv2itcHxa0C5Zn4BgMPl1S0oMmP/awpL4c40LpXRDjEED1YJon4
bUopgnfk86B9WSoPJ4o0Va3lhohITYE1medQNIn3VfrXOVBCaiB8OkTUOkxbe1WI
GH96f9hIm/Dp8Bq444x+MwKnS6L9WlxkGxj7pn/JmywNGVQ0A1k30DmkN/GUWdvE
2Pf54S7Q4vLNXADEw8SweuwMwQN8MC7LFcJji/iWYXaD8KxufF+sEUF2C5cbPg0O
9GblRF+Pun96/+tuznjCr2vpR9Th8U0u7b7xHi4Oy1oW79u0pDFUz/OTW1hTazAP
kIJNyQ6S9tXkkKlRK7pUaZBHRMSg6gEZyZPV1aoIXq+9LpbeIADGz/06qvnWWHY8
708eLdtJ7C5BDu8jEbeXkWO0MBc3NQ4C9AdvpkCz9sFrMEgv7qwgfkcyNzW5YSr4
Oi2y6esrXVhSwQLOZsOJA3/78NkRY1MKjJicm/mm84wTFaVrnK24vwRHQAuYFpMx
jyNucq78UiunsjAyHb8NeMHSUvrzs88qnubKA0vb3kaelocpq7ka0A7jsrk3GcYu
rpnF+8bpl5q8VkovINpCU/npax1JNy533I0tfpQWeU4s7pSIYblC11AezR6c/rXU
YCTEeBw7cF7/Z2Qc9tZNQRHxKTM5qWQKK1DcVKuKoecsjqHee5/VIoKOM0iMks+c
88804Z+LJ3avqkYXdKrHxCpuH6/S/r1skGBRzlHtXCbXgLOCmL6QseWQ7pmjtdn6
1SoEXWxh4zy2YdJumhY1f8v9lY/AfB2FzXGvgBWgHpzJJXFqw54Jf7gDblGtjmwJ
wQjcFX7pi0REPvoptfVcu16kgimPqC4e7LWsUEJTj6E1QhaCARz9YKLwNYXr8ZGa
gT4fGkpDOKa07B87GurDVpo/jh4nsmuDZlq0PlxtrjeskBUUdT+8yy50OdlJW8o9
E1HW4zzzHn+XxJ/Gj7YueN0us0gXG1BqB8nADuN6FJcoWSexCjIEZCrtm/h7E61E
I3FulA+WV8e6r4+mhU1ZP3dHwtlCJjm4wqtQmc9yhxd7wbJJemqvcOewKM06BnDY
rAT94/HdepI4zu9ripl7rBramEhdLJqH29PqgrzB9F/GPrjDUwbTzh/SbIwb6LW/
TTzaceJ+L0B1feeM1gkEbT2F/wxI7q9SmWUma24BiEMSRgtueNzdOLf7Otio8Br+
d+KVxd9ZvSIo+bsYOprN5BZ5WufCprKCNg2Vq55LXNS5Vk3gc698k/rlh65Ggh2r
pukgCFNCHTX0r/Ul92XXwnQd43NfIrxgamF6a20EXO3b/6VK2Xz6Q+CQf0mZIP/7
emhjLwHxig0D5TR3hT0Oae+XaG1GXgAbw+ahbDFh9Zoe7BPAMdaKtoMfUO6spm8s
GHMTcMup8OlausMz4JpnLK1kftaFSNuDwTDWm7DcNn/4g2yMRSkSkzQsvmt6AZnL
yzyA14i3sbf4FtbLUL7whw5sHlZ/ax7sMBY1pIGWsbjk45r9w6cCOXoDVGdiL7Aj
Vvt0E13ZKBohn58f5eyRbeM31gKpb7ftEr8vxsj0MM0gD462VWoS9uZoPpRtKVIA
hDLD/yH1+Tc57hwkIpUfRk9DHNbo3gOEOus92mdRv1D8shXxc003kJtzjNxdES73
jD5VRmJGJR/fLaDRAWE2t3co20wO527wOPjv3TzrVeybPC01gampTs+FFgS+SB3y
9XfMI+Akzc36mm26rQik5Wp9GSLILnaKoqFOwkZuB1btUegRZO3H5KFyhfaByRwf
ZFf0WAPTZSiVzp74x6pt5KwP6+ExRfRfOrvRmdxjJ6saDTAYHL3dckx0QSuVmkBP
CUgs25n/90Xn669z7hr4k5Xtef0pvSkQPdh7GxLkQ/LcE+Mf9EYNfpkmUd7V1Z4K
MeiPt6V2Z/qZzyf55kl738eo1YWTzO1R8frU2P8F5d4h5BThsDHSEPK4clBm4RC2
2Vw/q9J2jWb9Bc1AWIJZKZxhPbDPWe6KMXbDrz4kQ4Vswk8vyG8Enwtszsky3qLQ
jt1a/M4LgTJdVNxl7hCrRir0xwVnz0+Kkq3lzoR1WU4ktOERHEZSpoK87ci2PpiW
cjO6njsEfg5GpELkMz6zbJPSNKB3e5qJGLEKl8pGy7wwT/BoprQTgdQ7lRyRmkNb
jktm9ATGwIT5eDEJ2iOCopTlU9ClD4zY3xdcuPCgBhnHrnED7AI8k6/45lWCkpg/
ssfO6cPNBixVCd7P/9yCcDOherA0HegYULNOq8nLHqbkoD8ssc5qQHyR7lQbY2rR
ozLey85VLDxOSlGbZAFx1AsbhIIoAXfBpOwizALp+8LlkrwmrrkLy9pHlmnkSryj
mFoisPVoPOaQt7wM4VDltweAKR6H0lGvAxLO4q1+6dnGagEHjah1wM0r9HO/eYz7
NjRusNKf1K86gbruY/Eenl3cCRUSAXD0ozq6cX3M5doghdZc1UmRXMoTVueVJFl6
xmuTsI4tuA0B3Hu+j3SQJPqXUtvxKHrahaGnFMIiJ6AOaiOSQeLugRGeIyGmXvTU
x88jDVMpkWnpfcBVXdgfpLWBiHWclD3m1xnwG6t0sqxfh/8S29quXpAhoiwXWnu9
wuv9dz0p1cY/MX7K+hKZYNBAjHMj/DuPX6h/TagBC2J1rBjBdeBqTpHZjFGkWWm/
lPU3cGuKQJ0FxOjLtfspxLrVTwF5ASXDmsmP7zgVklCDmbAb/5ge/NtFKGpazQYH
7epiF/lo1hKUQrPsCVTe20kehN80+9lTpfP8ySmNPkuxCulq15S9rWcCQDrTvojU
RqKvPWp7PJPcuDvxd57VtXdREL+c2WtlMjiopt7T/qTvpvd2ahJA16qFzdAOKaQP
u0gzqVtm37TohF2rRd56SRjy8tdoNJ341IUwp3VGgOwjVbvAxmJ7Bs7Vz8t7xt7r
Ze6tvc0pqSB7HCvHa57dNpQm4OhOMA3PS2rnyB6IWrfGkzZmQ5LS8gVrT6H1J5vY
Sklc0DOy+W1nfEr5gSwuSY7/ekD20wJCKp4XuahJB/iFN1zqzNKgR/YBOBtmky58
3tSDaZEay8F8gsDtPRsmzo9RDZmGFqy+P8Cexf6DRL0pA2VAAvs8dhwMvYcp+cMT
6Lkw5InoVdLYYZ+1nzpnwx8ZcjlTtz9ADYnoDyuZREvMEY/3hEnb6W3NhpuHvSN3
KGf8R50gXArLg6JghhINffbJUHOgEkKchLUgU1KMyqC9utb3NOv9DpKkuRzEEI2N
28OwR/4AmABj2SNE5ppSXLQFpMqzvRo4Q2TgcLIGFSO3201AKWNEFtfT4oYOzPgR
lT7L2bcFxj92zG3aikHY/mZg5os3smowwrSGn04k1IX4i/71f6lB9lhrEwVuC8g7
gCPLDcGVpq9uTEzNrw5BhOOi8nQCDDiYWVj4KfE3WXD8fOGCc1iu/br4KAgl9ZBf
2t6rFFKIS/v4+5oamhI0lxc1YaDVUlPHCzl1pP5Nr82hsAAQ03Wi2dJds4603Lnm
qb0mHJ2hfe8UQEVUKclnAQKAGFsLnk5havgOHlUMIlT71Qyo00BTOY3VypOgZkPv
+27wNuwp/1NeuZW9XTLtIwfEhmQ7LuSohzmpZrBuGmsJ6YFQ+uPA63vKjIL7k6Bs
8p1aPyZLC45s8KKGREr0X0yIAyWzXACVybPGlUth549ky12V09eZFOO+zJHXBMim
oQruMJ44rmzOXWr1hfrZE1CAqPSoJQNCpMKCdkvWk+SHw/VQBiKHlip+yP+iZRp7
g/vQLpWovCduIHCMExOSicwciZLHNrlYIbvi4Ykq0RX+WX8MJ0FXXu2gVEeW0s/J
LJPJow5XkaiqQAVne97vspMhatWA9cmaI9+8wrA9B0dC7/W0hY2MvqtWcdzbeYAI
6a30xJHpLwY9wQ5E3F71tRcb9iuD7HqigdDpNYT/hkPpIZDSmIa+98W9yFn/lkj7
luF9KoH7e9vV/7aOvobM6jt9driXCpCYIcVjzGzOON2tXdfIOd6kCGExuBhG4NTm
Uukf3OQtp9njb8CtqticHIlrVcK/0BFFPN7yPaJk0+leJc1Pvew/VsUsGcGdtuzO
3bp6DRwz4A1THW3Z9EjSy1vClORwzj8gT0Frk6xNOHbNUyV6P9BSPERhTNkj2aSJ
NKSq+mEba8wNvONv1/7DUlDmkpu6c2I2qteMLJhWYP8CbIRO3zrinzmALbA2ejWV
1QhkrQeTq8gIkGDlHo42gNiRa+6zs/3gX7b38lirGoi+95LdAA42dvpjquetjm4E
hCeS4JePrHTkd9AHnZScCvcjwQTTeSL5ytICdW4qH0z0/fQYxxPKAxacprNp92II
I+mDMOIGCZDWat0XxjXjLC0UHTUrh6OkiWRRxjHVTl9UfBqt6DiVhSIBS5WONpxp
YZLL9xdsLIJYfjGfvBxHgjkRBxkGnoFfJIa4ENBGs6XvA5Sb+czTeEwzJKY2HKY3
d9k8TvipzAszJAMLrHfIjv2GPx9uYLJbAirkUWzFOPWF8JYOmd7IUijnwGPipK0r
YSiXBx/sGtJJHDRgA4F+24WZnxkuBy0lOd8Xv6L7FBQJ84JWy42nwVsbWUWWwftt
2BBQ4CCuuWp8v3I+ZUaubWzjZkb9gE2A3201piImowXpEkQFETwh63q8UFoK82Nw
+xYfF44MhwZnTkl9Y+F9mizmmXZ7GuXBlSSWDMpikqrorxfLTa90lto8zYaNp29B
0E/dpHzHJJcXNEVd4vhV9+W50XYK/YFNBCBSolnMIRlwJH5847nwpU8s8jzxKLux
YlNOtOEDECCJLjyxrLursFwXXBu5P9BKNt6IQMu3TORVOM/cyNKZ/yYeYCWaiKNI
YK2a2MVVqAiiSazDcOWT0R4675VWXybc1rL7VjK8jV5TxvfT/fbe+tQ+nZdRp+ba
6sg3+n5p/R5/T2fBqOMlZj1TA9xn2x0xDeVtvq5F0BaLBf9rCufc35Wlx8mCPi3P
olWthdfoaG3Z89S1sofInWaxoF9//M4K3wS+ewFoLmVZrnZ4jw8YJv9ZbIHlzQmi
3ucD44jYXFD0zDENCHMWOEjkQTRJsi2PmBiAhW0tcA7w0PHvpou4A4ILgLWuR10L
1pXneMjVtqWiYCr5CXziCEocBDPC4sfgKh5JsMvftsmxJFMgPTDepPQph9n4wKDp
an0Nu+PKY1Xq2BR8TjwXP51URAc1j5Q39N2qhrAPjGzxO9nXV5PR3jgSxGb+yjZj
X6a323ytHzuWXu8MfrPQ1IhQ0RqdZXcPz0cW2M3Ffo0SZJNYIj9B1bL6Kn0C1MKY
K1/FltmlwnXv45kK0/tOTfiHwYjhZriLforucd03aahY0Oo76EtxiORniFFuc0Bj
YN4WyJQB5ixd4LV41FFZC7Vq72yvfqOXN4qR+SoJlVuq3gRhMFeM8gY1cOA1JWyX
iBHce9DwnzG71n0cze1Lp5DzzwNjKP9UjE5FHW+z17O6hTYJ4L8cKuRNp4jJIqnb
2J5lfjRO22KEQ38VTxS3XM8S0n33qHcLSQpfdCyjELuXIcA3aYqzBVjEb6AD9xmM
YfdF2jRXfr9CQP1THgQAIpylzX4Om2XuiAWIbcs0tYC827JhGbKjICssfBU+g78/
FnM+Qyr3DgR62wpkRPeRQ8Z7HBQe4BcnSkjTKcBqXvXpdePCAPkV9zGsBNCknBu0
poURtoNVDvLlLQbjxDh9880S2tFw94Nlczc+WJYAX/N5FSQ9oIfRdvIVqoUiWQO0
pzkYGFcQXCVVhtwaE3OdFfWK0A53sWM8MZTrOL7I21j+dQMd0iSteR4qTHhkzAcd
nLx38EbQCzRB5cQFgq6gmKglocEXiSxD7LfSXQHuOWp8DLWNDzKtD+3UhCBnvAWl
R2MnSuWdOHRuYPbQOCMnuPUmIsGlHQegHxem3u2rI7JhrhR1JEoKY8RX40su5/tt
FMkFGTsy4vbJqi2R3tuRECLSs7BFYCFXYTCnQGTG1KL8CvwkQtpnhxZhx65gjL2Q
hY//zHEXLM+zPVmz/32PA/7eRsnuDz+4ptkKg6x+VkBQTDtE+3SKV7C50x3yRrND
J8SB3XFuladiRjcQfh4p3hITZMcAEI252fJVpx5LHUBxnXolkHoJtb4eptYw4yWD
S26yDd9MFal6xJ3rvmJI1ELMGd9L/fF8l0rB0cL+/rvR7vv9Yu2Zkr6TZG5df4Vt
vANu2Caav5ecWzrLQ22MezVzY1lXTeabzUU5F0d0H2TgS+FKAZ5sG9tzrmzwjavt
mK4uJg2reod4S2KioVMzsB8eZpSPW0I/ukdI62PG664EfKlC2UyCKgYNmcZMvymt
77YXypNSJ4KYMq/3g05C1uK73cTWBgwaLRkpavS2x80qlQZNKjy2xsI5t+xkK0Xy
2kvAwuNnFjtTPBetW843Rg9PdCWVqfRVoXmIxwHejq+0102w2x0zKL1XzD91qFEv
uk6VJZCqfwv9ypLGLyXdHKf3ZI/2WZ1dSpIXXIW52D09njTj3tz3cfU0LRuRwNIB
SGfQkdZwq8wGsKpDcoL7+XIoDg2K6x+Qwk2Gq5YLFAFu8jHqyj1Sak9hrDUMhvsJ
QVz4W7t9SIUCO5/f3qMajEvx7qdGyFqNq0b0rNt1PtyxxVudCAShqQaz5YRbOdrb
cOWHZOmKzIHgK109r8xwuiunBtGn/K8bJIkXCRyFu8oUS69LhJGP16NHr+lf4h+v
OlrU5Hok8nrbmE3tuQeNQbwzs4QMUv3je4fHXIHV1RoL1UrkjM6TFXWZ/sEOzmoH
neOiH+pnrKIWun3dT6aGZ3I2xmCOmPtxjoEk6eMjgHool5EyEe1UVPfJC//+/QLj
mEG8omwlN49Z8vKxGmSux/rE0VUoN3Y8HdY2QVhTRidPzfNtF8x1CKjdTfY59BAq
9r7UVMFuOQwULK86wfs3BGQHbyfoF22LnMZQ46RPd0SN2aqykAcFZ2/Bc5Od3/x/
FOMLbFvqczK8ZqrbMVsSKOK0QXnC+wgMRDN5TZfooTwAluf4u+vMykzQFrEFXzoY
jbh+neeg01ptflfQuRE/95JkFd0rSTPHRzDbZAeqQed5c3Ajn7CS2PWNMmiOC2Eo
N0V1ivfRXE9nKVyQZ/AyFzDy3myzJXuKHv36drz4kOFmkBaDHGuFQ7vtMDDNeHnY
sBAIBgCM5cFXzgUkLEosHXIWj6Cpovu387UXEVx34hcX0cNdgj4je10KYauEWsUw
vnfcxhGd+dekWuEYCTH0lbR0gOmYdPj5+HV325fjGG2zH1gq9QdYAEDEc5GP8yv6
4b7r8jHJj4g3OZH7s5hKQ9IaVFYXQXbuALGEveKpD9v+9EIQwHncN7rCdUQyyxvZ
SsL8c3KV/kfpJgRf92WVUwMWLskkzTJvlD0vjOBeA+JuYqubj2S+3GHyBuwB0THk
14hUU+ivRMMp7ZO9Dq3QwvpJw9Sy+6+VHy/Ru6tpVNgLGxmZwNH7zAngd5mLTkFs
G4XQQD/B6cPRBljDbjtlSGeRqrPRtfhaqrXjb1gRM4chO9EFP6rzQXCzkYjJwobz
blbAbJlwxxdd05GGSLM8/DDn9OChVRoXsttJoFnoaTWRbj78jccU74pyrf7ddfxt
u+Z2y6bDuc/PHrvDYJhZ6bZyeZI/bLlUKdbKKCJJa4gC6ujPNOFHu/n6Gc+XvpVc
ouSuDSAq0JBHBbdf5GyCgROf1lCLRIcelRZOxtDdXehjd9xYpqDEAxdWosLTurwS
M0RCsseekvEIJxbubY2efd02P3NhGEnrtuMHDOk6Lo73UJvAQSwiRN3qsfHyC/lc
9nJ1yQuATV4A+aXWjqIVIMF2aUSD48s9LsHDgIj9IZbMT6uUSo9dQzJd8t0qfges
SKMe9KqUPdUkOHPM8fy81YM1OHWlT2lhRSqpiZuzOGkMEgbqPGNTQJrbazd92Cqe
6DNioO409X3HOIIX4py6mETv6hGut4eVImerZsjKdVJeaN8ZeLoUTIT1n3dIjbea
RRjsq/JxEU97ssvS+XgmadKptvqpCA5FGB6s4GuaKc3L3KH+MQ5akx3xyYhZLsWg
T9y8iM7URUkx7cP5sGjzrQk5y4SjDPo+F62O2qA9sliUOTB7xPHXImpMlegB94/l
93T/3p6zp0420/pHZrHBoUMw8lP0cgIeaWp1OkgtBai1xurb8U1vEDEOlwIhpDI0
oeXD3BXZZAImnpf0wf4aTu6t9WbYJ9P4kbgp3ypRJPCGLl+AjVfI8kVuygxTagME
cYVb7K4h+h4DNzojuaJBN6Fzc0JJje0f5lQYmeRUiD5zbykYAgoQBCrk3spL8Btn
mmP84/M7YgwQ1zVE5/grMmQE8kqJNLAMjzOzTjuGIaY9KdEcLMLMXZ3avDb57CIv
4W8A059fi6owx3+I+AvbiB9YGE7VRYdK1SStBfdpiB8e5F5fBrRaXNQ45WPxXWfo
MXmr02pav39Mn9lTglC64tIaTbfuQMOPz0AtuEICnfAANi+FIckzOSY5MI+Qmk4G
7qrwQd2kO3bMfBf9+ZubulvahF/mx7qtrvRghQa0Fkquupeh/d36t1yFxloSXQRx
Cdo7A3mWNo7tkUfarLi3vIXUG8DFj5R3whO+ii9jeBIyGWyJ8u7pMd2sSREqjLdI
alkDCbvij/QIk4COOm7xnIywmWF8D1hw//gdoLHoBm8WJ7sJfYcfVy/a/TtKOjIC
qUntYMXyg5S9/IpD4kZrDSq3Mn4wDQuee+LygO627f4bbPd1g6p9HLg2g+MJPFPD
OaBYIa9VUSAsrSxJeycXeL2Wc6lBUg2h/sxH7BI2F5t+8MsCQQepVWLY4nWCz9aH
WymB2+Xq/lv4DsGL3bany0ZOUQ7q/Om3d7z8AihWkMKeerd0M/ozNleinJbioZgc
Toz9MG9geVl8VjQw1evYimohc5GvV02tICWfMmZWXvEtAIXm+yaT8mB++0xHhpc1
rO+Jdb1rRj71skCDIbCNLZYOVw8EBiIuZfizHJJWRrByEdEajJhIUh61O03TPUAS
lE6HJsDsMffawpnKblORZ/D6HUJ5/aDyQ4tdxDs7LPhCAIwdI9C3t9MFnV10PqG8
Krzws0hE0HVGCsm5OIr00I3n/5qAH7e9pgCfw6m9+vO3f+BjP8jDZ/7syAaXLNSr
myFmGIfGCwU/yrLC0XF/K10ak/FRRKdJ6P5GVagI492+Phexr9a2ArzEV52OcpNc
gAQ6+D7x7rI4PeqOlc8UL/hDgmTCRPC5udy4QV6Pd72chCs/Ullqn8OBzksk/+Fk
ijQwdFlCbcDJTqYKz6oGr5SBLJc1IYSNV94L3DscItlhc1cCUV93pRPEAl+tv5Nm
rkd7xssiku/QLE5xkkvT9afrG66/zHI08X4v74rOehCnJq9Wjo+/+3XFfJkIok4B
ErvCjp0La+AAsrH26Ya+ATmh3wNyLlCP6K7aBOpTR/jLnL+KxsUQ0iQm/6SWOKlL
nYAZWEhiSYDzdXsLbQBkd/ZWHOqtjvLLp/wSonC4OcrwlkQYTW6EuiondFcK2O3S
nJhewB/1SdE7T1uKEEyax9NoiV9hn9+3IoPTPJ88djrbsMaw251uiJAxc1NzlAJZ
IjuzFX4BXzQ2eNG2l5W2Z/rFaginw35PjaXkb4Bu9rvpLKYUyhXdetNta1nvNGIh
On4sHa2k3v4TtEXdxEphz66NSV02PjK5Atcjcq2FYU0l4JJp7r0MUXjUH5Wcu2Qm
ss7/r5Rm4QBkUPsN08K7XKFcQcwVNri+kqnTXOlx63AmhMCwHMaN0nLghtskIeRV
O37tBAloZSo0cHyqafSRbyKk8oO25syb1rvgRefOXyp/aJZWOGuG1sTE1KaF3HeJ
3guIpXrx2BU/8utyGL2bTw17mMmDbkyJLBEbu5nfYiN4f9FuAvEmvhbOs33O1iEE
BFbK07I2gTB2V6gQGT2G1tfHPWQg2b+NugCIiOZvXVRLFZLSqJ0lFcCQpp8Sz6QT
bQx7oJNJeKWfadIcTtUj5xSdoBf7ge60LrtzGXz7bG03EjDXKwC6q/G8lE6htwOO
Kq/voayQukVQVSEvb1xMReMonqnuz3dAk7zNrYmMEyQcuKkNkFavCtif7IS4mdQn
6LrlT5dulWqUCbe6qxwEAp9s4DuGS1T8DtFBf59FEWR1qgg1qBsM2KP6W4gIPCFd
2VeYwgt+Rrh5Sn/vwR4r+ge7MI+K8rjlfcvKFEZEIR8MToqLU29yLly2MdclVjwk
aaf8o3wAyGWld3JA1tVi6aLqio/tey7Z2QnUyUQnIsVp01rv5G6cYPPg3ySwbiYZ
a6LVkAPAKBk55HofnRyNCX21Gsvs4zNp8kyXugtPrXysYG+bOZszGsWxrzJYejai
kKIB1D/9BLuI9E6flCIAKLBS5FIZvySAGhp1tM2ZmMcpE7FnUFd0AZs8y95gcPsp
2WlxxaUt/+fsHA0zaAvkYNQnqDJ4f38a2TWOl/JguG/S/fd+UHkYXxFLRw5t3dZy
WWsSV25ziA8kXLwix3c5QNn4ZuXIxxXaU5JWT7aP5BlKs4DIcCOc/8X0JbF5jk9T
3+0luVKUiPNkNrig/bdenLW+VSS+WFqWmf/1VWu93UI2X0G4jvgd9vsGKrc2zuHH
pn575XVwyPR02XFq2ep6xY3C0PDk2+HugUZc7l/OIIk4SGJ5LLCJoW0PW0AePKhI
A/5IQfpdwItG7z5/OHzW7BP4quphkHEL+ZB+PsOZgnBaY2qVu/im7RIT1Gdp0BFQ
ltz/xtb77GFHg9UPigfmoTvk0mWJxx9oySeqbjGxGuZa2u1gPtvdDslFJoWimeVW
NT+ACBDQWuDcS0vJRAFwl8WkNy1yLLCoO8sHAYNtlDiGhAg6YIy6ikqftx/dI5vv
Mw/JoxJHHwZgjn06uL4980jCd9U7HcyxoJYIjiaSa9nCN4mMYv6+lgtK3eP/6sDk
rfOvmiVvFCv6HaMNiFRTiDUCBOMWBIvwVZG0zwY5r60rQwHwyH8Esy032KFHKwqq
ajOXlAFND22noasG5Va2+/Ua+bC9H3wpL8vAAwjxa+2xZgH7ki9qCn0JteHJ8rLH
q+KBLra9uiBCzgBzeurFU8YtwJR0Ksuh7aLyvVhGnwle97ZOS+lrTh0Tawb/KmNR
s1Vh7R4HYmbfuE8ukBHH+CnaPE/bp/lZuDd9on9ivyPKhL4fvU3fKRly2prrgW3m
5gFcSJp8Vgb8mMDeqtBbEnn7tVjg866r9MtBUSudGReVnd3whQoQ9MR0orsBAyxr
LzOi/OL17+VEVh2sy3Qtd0xb8lCRGsdwsj6Pz5W+nZzGPJvJWIjbrWm448bqca1n
HvvFGsa7Qmlx0VTuxBuy7yEeUgkJgK33uYq4q7LigNzgVCUcL6Gsj/WdceJykMlz
nimDImci6fwkpw1cMSpUFNGi0LeilUScCP52KQ4IqDxTWh8Y8+lANpgzYlRk6Q8o
if2y0lewWZCKLrg7T75XPHQb/mDQFitZPAuzgMjwjnuShjuK5rQKChDR9eU41Er8
kaiU5ZZCDFs3RlFHR9+fxRq3XNXOvn1j7J0n87hRfYulXbKuyPdX54P8TaOs7SdY
HAAQLJgEaN5YguT/TnsACZyN40bDA7JpwxRybH03narBJVVmJsM3uvca2PNAVFsu
IDSSm2+JeGHMfazkpdadG+91EYjUeZiJDUBq/NvhX5lSJ3FJ5bM0IYFY5didedM+
uZ15hceE9PIBUhxfhqACrFSd9c5C5IAz2zLaLQz55jM0vCZvNfRJWlpsFd9bLX24
XZwROO3Mt0UME5f3Xhw6GnsO1s/astw4fsKXbqrqyG7fxieuqCYiMJjRrKanvlRY
L6PnEuxVcpVfegZOzHKtpkFTZ/0v+Ykc6HFE/81XQKc2KTejwqgaZO+E69EYZWNH
J4I/aS/hUdVgxu3w2rnqF3IgJs2qM3B77PZqh4gP9f1WX0wNAzsJzyQyxTepeiP3
otoju+WEBVBc4psFsdlfAc/VfLQMR13iU4sYiPavrzQdj6imO12kzkfPzp3N+j0F
qtVO9futtXq6SFnppZwgv4l34zOIGTLsUCun5TPBXoP2kU8u4DsR2e5tsk/tOSj7
K2ZPjLNCSVQBQSxq6sM3E8cAz0S7irXgX550HtSvB/ruJUy150xBpD5yk6gtTV1t
Mbm7WSJtD//jUesEyFnsreeMDDbGE+F6EDKZiA8rtVvqDSjvjnyLNI5QRMgfYqEF
Z+bB1RBnT6ISykjN0lDF70bPN68xz6f2eXWcoaAVDsOyD+5c4PeO3hOD+/JI1jGa
0wLvXKGA+g7h6UjJjBaJboPvqR6C2n4KGdtxZHoN3jT/seOg4WAzT5C+6hKN+WsF
/Ln0vsg5dA9H/tyWEkiO6YxpDygJ2ueFH0aVXTPwWiGBJnxu0VirqaKOe58kVZRW
sv/iwGTAIPX0tyjhhdgxzPYFiRGvNAQKPCaz0ErH0i+CNs14/iMZ4rPLo2bQ9lpT
x+sKezpath0oAcWQyMhkWPECaWR70edjXwa3mV0wLbF1iYopgO1PVzDSfzxvgJbQ
69Gv3MgixV/64RMazbnVBibuGVMWN0m3F32YTCrk+1lY2Ie/hUsHnQgKnAatByrR
k9s+5Nz3TXQX91wGFCttfYq5SNwkc/g9qbom66A1F2/TrG7vv21FfII3xqxpgS2v
tMBwDXBgyTx+jyFsjs+TApF61kLqXl/pqlb9BZyOMQm80ZdTWK/VWEX7cMAeVgv9
NZnjO7rY84BiJ12hxEjNlbaQ2XD1M8bs7fTtTS2NQ4AyY0P0gevMSlV6gfZRB2id
TYCowAHISuSlYzaVUeECiMvRS5GjcCqWuLiE0wYyyxPmVXiiGW/dJuCti0NNAL5c
pXrJyI5pXfTJanyKpvQPI074ZBla7V0zMof44b8RsWE5clUP1tApmHYyPI8aN5Xl
u3toKRGW66iQNMX7X8lFPGwSSHKe59435NNfnzdaJZLI21PLdb/WlvqHk/u9OXwp
kb48k4koEHOnyacvNuavjYHNx3bGhs/X1o6LVOwYqDcVNiIZsad7uHJtmevyn+T3
yyztyrc6cnLa81rXU8+FpbsQ/4NCuwXF5KDuy58AwdQ+IeVZRZXUzZ+lqgXqB70O
O4zb9GJHWvpvj7BbnpbZqn8BocXLzF6y2Z1ehkfmzDW6xzK061H6QZlz60VGcTyJ
Z4oUexk6fsBNcmJFwzALsH7GfY0B6xLEvpKotss6U0a7LiBpFW4aL1vrEqjUgTuW
eDsWu4ZlT1U9cuJQ4DUMDQZkYuuZ/lIF3r6fxPOQKt18a04P9VPW4+WdAz/5dSep
oC5wSiqixN7DyxOzbxJS2kBWWp0WilW68sLe4W8IGDvtGDrfGBnP4sJtSKPgDOFi
jDNr8mBU+/8rGl5nYLgrTddUicHCVSu4j1NN+zeqTUNX9gfjeFn0wccC3J/PjcUb
skRCvYPE7kVq+GeEk2kWtYtMRGU6l57bcnfTxJOmVkmd74eYbNfw5Xo2nS2DYMow
xIf0lcxSyn9/61oinStVXZCP961NFBhHD0qjxspQrQsYbv0W7AQwBsOjg2eUYLG8
KQ0KvaT0Q76KBTJiiUMEE3/ms+mhv2VHrP5F8QIGUaRdyCWvsJB9pofhIrazzOl/
+HF1LPbRnf1E+okC24REzquaLv7kVIQ6xMZYyo9zzYlmOA0+tFPJI/aqfNkQBVml
nV4KkLL7PvKmYFW5TOTw0H4JLAIos90iZleZVwqotNYkyHbtjVp4CvJ0pfVH6BYo
R9dKgKFJQKKfv8jOKw9B6gM1Jx2W7SXZ9BPghn0fs++xl/iIa+qXSqeN1kneYUir
m3CO4phxlZM4kz9UYdrUpIopDKHKS3vZ+c5I3IHUBCP4m7RJpiP6AoMDO2nDuGN9
YdQ7o+wInDNz6SNeLq/kFwfxOe0aM1lNYtjuQPnwyVFUYPBLnEXkM8aUD9Azv1nz
EkkKy4D+fhymgvxCxwOFr6R/LoHac3j+IzVbpmxrlkDw1xZ5kODBZNfT7kRcu0TF
21v41C06szKVQ9oZ9msZX2jNqtc/NuF2Te6OAOfG6EtNYvdfQBo8BtAutiUioYu2
Odsfh/2yS9rUvPschY8BprHZ9wXf5RbDJE+uncBUodgvg3EGvZM6hWeDkoqX9qov
DHs7O9d9GCfZfgKCUJZioIbO5UWvUJyb7UIJLAkGcXfFvchfBvlmKdEGVUiSEOQ6
N4yqIbEa701yStZt3ESP5lg93yVdU9esRm7DgB3Ljv01JnysB8IVzVl12grRjT7Y
vxEMLN0hkLahXlJ5zBJ04CEeuT1OeOn7RFmmmTFwDwVXbzG9uR3FFr1CaenqZGAU
ZPYtxBcicNQ6V99hyatGiMTesdm0BHg3popOt048VY+fCSCNEQ0qjAJ9T2T9YReB
vZAiZWnniNys0uHCQS0bUmHruuMcRVrHmSWXgkt28d2kBr9Et1EKj+xFQwIME2eO
8rtZpwEi1E+SlZBfhPBD3YPRc+MMSDZ3FPw8zSPC41tFiRHSWxRgzO6Sg/CS7nEy
Ev+WxAH5nK077JgbdmwRH7WxtbACVAlG2ywtHiXeoeb+xWfZcAU3Y21Dad1wtTDD
3ZZ7Va+y+5mT0bBbTdFwBKW8k8U/Fe5Ftwb0QSMUPuoXfJP2YCf4xx5CygviJCwm
ZRSemk/BQ6YQxEvDFUzb3vvEkqSkJ81KPB308GAG5eDkUj1RLjAAE1jyeVQfq0CV
1TC7ZWI+u/A+sz/hUy4knv4ddnXCFJHBohyjndGsBtAatSX8oa5OGdqOpcy7ZMfa
fDIHcT/LaPJ+uYVF0cG9y3dcHNRXTPjvdJqYGAe+aM6rOMn3SxZOqCXxfI+YPQiJ
cj8OogHjdm9vl8YggtZBeFZy2zqt1jXZ+qH0U2kW/dahaQIS6Td7StzJl/pcm0Q2
R5NfnppPuFgrE0MDYiInr86APiKM23pFOAMhMn9LYIuUb+Kv9s7JT5RHWIyOU5C9
KiRHr/2NDjTwDsKYOGTXCrLTNwyPbd3roofW7Zyvg2x+6f9Bvcqs4K6lkIZLl2Jd
TPPXug3kYc8BpChEVWRT0eRTjiKD7WvkILDWkfPcNCsdMXsYHmLE+S68HwvrxgJ5
RbVCJkWW2sP1hk3c+8X1bIvOcqhZ00S+qJKJ3YWet9Np/eweK83FjbspsDYA297E
6xfl5kesEzWrGDQeiIEKpy1ahf+2emvsxT9deHvHQpZPa+zSgnv61pJHhmdMdwBg
RV2vxUENSuLbTufrgb6Iu7GDV+oAdV3K9JmcUVwmRmlU2Y3AAyoF2H+cQh5qZi5w
rDPsx8V8OUSr0aJfHVKIiBcSXgwTbt/NzMOg2eOuTolsnueFcA8O8IE69QT9IMkv
ml+T40p+o7kjXbnSAnv11PKDEi2etLES9nBeOySQtISAbVdEF8+fNASGw6KKhSpV
YHeKXuFPasTOxebhtuVazGFuj+nKuv497tDYJhq9GZa1IL8fph/lRTT86xY64fKC
x9ODIYpmB+YShjO2BAMJ2ofXHejqhXZHGUx1+SSGqrvAVlgcP5eeLJj8Q9SFEzqZ
dXvhrVR7rT2NdQicfMNiKnVKT9TcI9swMlkXB/iD2nLGpbJpli+5jcgZyhrKYO9N
CIbkQddJpMXUWuGvJnXc02F8UBS74Na/JCLbFDbePEnOVl4rD1q8xnN+R5B2PJ0c
iFawlTotf/6JjIXkvVK0SDNgYBFDaGad1QW0GUzqOmGAfBPd3kese/m0ckyzxdiT
uM5RbQ6OToLNV1pxeXkTd6pKQdSTvSjpSn9DR7XWfma3fp/1L14olgBDwcRxVug+
s01RTaJMXyrtiClWqy+x/fPwmZjrNrIlcSwatB7Flf9yTyTa7IHRuEu5/tHwuu2F
09VJ4ylPXkCVreDI0IxFrrF/RugAMft0KF+pHvpoej7MxEM1mcqKXGLU1ytQOUuW
oEqPRSu5AAm/mNw8n21GaO4aBYAoy9zZrZx3xp3JQaYs8NTGMNor6c1maLg1LqcF
OiPioLTBTfPFI1+RhMlC0cD6F6G28gFWWfotq5hXHiV7tK3x+lIpi5nQ9b1KWGQ+
OOCRDAstq2vhrcewKxAKbccp+1319Mm8C9uBhWJIpUoe+9np5nnMrlka4ILEEgVA
V4J6JvRLmdDqXSuKti5Kn/nfEnv9iQGPzAS4jpMUCyMbmevn8BnrQ0akrJMAiyoF
S/MXOpKJY1O+K6vNWE97GJz6f9tzhqIkN0dBlotZnLx4PsokBX1kpq6JEOwru2gb
D8RhQNkXt395CXOcpSlbFUI2HFVVYZf1tEUaQDDQPjNYsUqbtrgsRS4vvM0mzyKC
FTOiupwOqg4oGaH8VymBIIxEhdCHGjM+HX2vOffxjN0tCS8l/CoUXkCymD1dpPUV
wDJ5KmdaVimWtu4qHwh5CmNOYzR867vDvyj8LVaroAy8g2VaEYOfjozCeRTHX8Li
BH9qqCiTZFQNJxGAftEVQvz5ou1KQH3wi3tm75nCoxBGhsD8iHiFUQ4Fq/gXoZXb
MYOesa73+ksvHu1OpzPRXJDLOoyNknaNe3eSomWbA02p3+aHcTrnMDLyvZ0HId7r
gZ0xSS59/4IAIfUFbW7XIUD+VN7XEdmYm9XgLhPGtFLBy5Uq8bmZqY1Cafh13p1M
YhJ2X+qSe9vuS52N4vRYilIZkzB582F5qMq9AHpHZZNyN9ozpUZe528c/pJV1hiF
wvvL7VSEnpvVt8dvI118+P2/LkhwUjYPZ3Islrbgz0l4ToMQMkFRoDq2F2lHRY5E
owVbb1wJ4zxKUaV8AM4iExNQdT1mXMc/WrfZzFE+Hzv638fX7Q3RknbI6AqX6tXv
3MKLHhiZ9YddVQHn3wwkpfoqThNIm9hjio7vLwI+FjNvmg4+FcunLTi7RfnSPRXi
67Xn5k1SA6g7QKkOzKLsgIMHXbBWszZFJY70qUbZhwpPNWywcC82qQ73hoVcLWBF
f2C3xDM4CczLeFuD3fHF/5TyOl1XZKJLKvmqkzoI03/qf8vlWFC74yRkBgRxnjTo
Cm7YPCgcwQ736HABg3dgIeWGQHus0lzQMl+1Faadj+8T3n4TRvbKBpp8BBrS7UAQ
2C2zhYsxD+/NPI2mQlgoD/771IgZMApFk1dm1zjNPgKrV37SVbW7mzcVOcnGohB2
p+ztzgWfOHrP9FJScSdhWnODceDP/DW86rQvUsUP95qxwPdNimDDWMMzc6aP2mOf
ZZM9LnKw04F68WrR97CERKPew/c4yKsRCbSdYO/NEbFVJWzRwSfBOWDgggXezlle
u0/auLJuvRXqsHp6BnAfOvF7N/Ur/NC9SDB54DszDF4f66DTrXUP3TOk4fAPXtMV
PB3mnn4yYOHbIgcS4xJyG6XPkJzzN6g1VPqgp5jFRacQdNGoA2Uf3nn+OKjyuELs
WEjtOy/T3kYCNlW79tnFZiM74f7dJfGrT2uueTs92WNvWenyGukP5BMT8mBWGFd2
c2wJRo4UiWMT2LLrHAMfPBVzlKwjMl8rKIXaOYofPLH3PaEpC7diggyDbxz3nfwV
B6jjDrjafv3ksHZBv/wupJdQT+0zl67oj7mteAu6ukQEcr/86KtwmGOkOK93ztO/
D0cg2bmkLkZQUtkEdoKx2iD1r+uySoBdvv6kV0Xb6rP2139fv0uUZstjOL0myJ6U
CZex59MHtSDM4jV6Y65NfaGggAgo0F8aftyG4QT4SvE83MMEwUgxHoRMRENJaHfE
0u3bB4HVJfUqXijyBGDN8HFLEJ41yUmUou+62aLDs24Ix3TrfLs8nU6j2ITIAWsG
yFyBEhvK0nFYQX7SoR326dReLtL+g/i4EbawPcgS4qf99X0OC7eQYEnYInKCsCKi
cZMkCLB+M8R+6VzOT7XQ7+vFiRPPxd0NcWWmbZwC3juzaPpAPVWcpsGebkhz9bTu
n8aVOerFws63usJMB30yFEoa0KZEsJv+llz548IeTTAMqw7zkd/GHGna/5lZAaJr
wxlYb8PWRmkbkk5mOPf8Xx2S4GbAlCc71aDbk/Sg1b3kbTCK/ql20GuNumuM3n/V
wqC0lzJFMVmzOSlAyVLjK3qXejR/qn6ZkB6De9zNKST4HydZDLJrhOwISJSphoi4
O3R69d0RbZeTFFcZmbU7Ag3C8cpecKHOF1TodrApiKskgynhaylehAqkw1KFke73
Fo+h6cXNyy/3eDmmdCWjuLpihqvkUBd/88q4rM6QZ6e3Kq7S6N5HQliB0Y8awTUZ
GX7tz0RznbMQhYhJieN6l3A9j/oJ53UQt+alB08j0ql+stnCrwSWc+A5G/TnLrs4
bZIc8HmeZNbB+2VwA+eLBOSfG9QwuUbqjXw9V+qaMJtdqEoACFj71+vXcBOBAJKV
1grSl4KtpxITAmTGi8jao5AuC4+B9Lvi6rhEFKYlvhn0yp1iBhMzVnJeyqGv5oif
LqfYPD6PCsVqbntRNG8Ab42Pkjr43phWq0mC8Q6+nMKsVVQOqghnRdsh0ST4VX61
o8SgLW3NPc7yoelgko9rRZSf2G3ejigaKK/R3+nZwIQ04sdgDMZ9EjSBQgYloDIK
g5tGBjVxU4QRwHzUbWYpLGYNZcFRWJQekIDG1csvY5S2zjTxTmIUJo8zETHGCuga
CyzB68oMCl8eMmJA/d7zlHsRjEQiMLWGdEVrj/WzTd8nFLSb74pZNlDMbdCLBAhv
F/2Pux8C5g9MOgWd/tlTgGrf9hki+MH/aISa6JS3Ypz4GbxvSHQ1JU6G8ut8G3H7
MdFZlVipnI/4m3LyWMJ9eSGEp1p/7u56ns0Pg/ZIrDw+L1SV69eQvkGK6Z98+ftJ
NiNjt6Ef/PWyCQEDxElaSUo1kPPN0K1ttYG6TpFxkJtTwKRyN95mDGpe6D0I0AIw
WXK5zqvGrTgJsKmriFZHxpobzWwdvW992DFEMIBq3la/LFvU73ZTJBABL4b8lPpe
uJbnl093nkBvaSvxrXpSfLnX+j2JXZoubFhpHSkwf48AGd3yK/1JH99X5L7GAqzv
CS5xj1uVH3cksPnGhEdnsPtupOXpotCapGUi6uiqQhRI9jw8y1F94ZVIgaIpn+nr
+sKRisF4M0r6NBU+MlBk5UEnZas41ic9zYMs1D+y1ggxx8JrMQp6WAN1QoBARCdo
xfjJtLJE4y61JpX0VPTLrXJdQAHbpA9W0oYeNnoDlv9ISr4PzmFXT2EisI21+9JH
vg/03hCRUcKz3Rwxehuo/0aecSex7106NarHqcZlXIZgXJRXjmhNU8u+nNfl75Le
xm5mcq7HAxNUbtkrAn7RbZT8lAvyMVR6lHe9pdpadhYp92oce5qjOUxV/hr8Mz4J
yRPZ03iOWMnXMJMBU3/vJZgrzMGOKlXoWtodHzYj+tsr2bOT7+5dqTrb5deDgy73
kJP4oL7W9adL/1ZxMiBCW2Cp3SsjfvsE2NOllUuFAVcX9UquZDGizYJ+NOYd8PUK
j+taanpbE1orFbjxRq++IvSyceJX6ru2CYAqyAv+Oft4X5rqsnrUUE4BC8Fyqifh
nRoY0fsdlsCIKRLzE09RL/bUreUbiT9yEbwZjPJe/uczDPBaSjMVFB+ZVyuj3XpQ
B5LRdnn8cHImYgr8QaxGhKmnu3PCk7XUxkQAB0ppsyugGtHc6zYDXoMOQU1nWIO6
mzn+noesKUqpo72Pm6Rw380nFV4JtzYfUNht/el6/CiMSnH06U1xBVneD81mktoC
e6UzjEdIMrqFR9lM/oTn386lzb3rFamSvYbhYiiAOwLbMCATRGcv0hREzMIlwqPc
QBGdHbb/ggpmYwbPntCNsqUzX3ljqdQCyb8jYB7cW3BkSUK3S2I8sEVL244ZHkww
i0TW9Rc3F9cevVFs0WOQGaBUWxtPRPbYoNm46rxVajHIIBqwtWhNuBd4rDmtAZY7
QOOkB6qGsj71fvVldW2ebnjm81C89N3LGO/XhJEF6jSfQEpS3P7AHKi+p04qB7Hc
u3ImoCaqNzHmlDZ9/FKbjoR2Vkhq19ailGSWc4oEkwQp+aQTvZ086ygmsNCpVxjD
F40wRBu/0qQ2+p8hD4Ei/yn+Mu08LkiiqhTBJmD22s992s6GjBdwNmP0hZcswQxe
Q8xpaD0uWvvOH5JclmCRabIACvCqYlOmN9bxO5hW8g9dYmFEnOcUhz6nOTHuYE9M
uaDbj+rAlWJ4o6+ZKL7woX3tshBWTL/rvsi3yxcrrPa4PsJruxVrySReL+CHq8T/
lB3Qvyg5v542XdlYPVsuoJi/lNq2wN3PIq0v9wduCeqbZdlbNpqA7hdmLqYGGIIy
O4xIbqfzn7KYqeBVhPgqJYZFVC48hjRTARnO7YpltTAx6W/cjRi7VgjRgpnh5rEj
6zsWZk7j6xCX9EEVpMQ+jw/iinrSv4XNuW3Jz22aRDg2cZd5dbQR8E7YrLbo9oAO
oIXX8f4PRMSZ04zYImX9EwgLpNvrKxlihbC03LKhi1XpqvmC3Te/yxtOS/03XCi/
KlfkJzK6SlqrPLgdMV/Q0ayBSdJbgB/VkV6oXO7xQqwLukuKbtSLNKqCrcjbrVxK
ogqZNq8nZ2EFuW5q1PVArK074QeUcnE404+7MdZN4dwdNfL9DNhKvms7SC6wMHmH
JvFeqp8shAbmXCH2O/QBh9UjQ/OcJRLg3i7xzXe2gulcQ7KM8ZCxsIPxmum+mbhC
lfA9WU2c2g6hUJV8ZKqLd70klPtBzZ1EDXF2rrZgTzIVpE30Z6p8dBiJD7T6eSN/
Ur7sgOSOM4A824uWbbBXwcFIJU1JNkZlke/DvGLBu6AFbE1Q59l54Pby9GE3laIC
A0gXe7fDMfW913sl83uF/hWLRhsakTtXPH+n9EIKrZlu9qa+gYY5HM5P86LOOVEw
FNR8ZQ0AUsNvMLfDNRjCrEfg9vo3kTWAvsHUOCJ3gpSFfThS5xUBj3x2tSoNtOK1
f6XQ930vsLPkmTwR0OJB5RMpyi4HBYpW81cJxABTtcbdDEsWmATzKAZWLKuyP0lG
biT49s8UCnCjTJ1EpImW/5haOI4uY39AexYnOD1GFaqJm12HyEGqAHWJctdGgNQj
y5UWtDwxvr/torGDNiTQ7FmhywlLMPWlkLC0cDiNKjpl2kjO/kzzVxDyCkDjutmo
eCOHHIvCVbnVZYM0bwag+Pj8mahv0DEUWJaY+WXFKAVMAKZuzqyy8ygthtHKLosN
n5HDUgEFWoEWrL5Ky2ZZTyEuITTWNEzeWjK+V/x6rbZ3MfvBPK28cbrUNH00jsct
D2ka7q+Fin/53AYsl6u07gfxe8sMhJw4SgRqs45n4GcQowV47Gv/R3LvbU8xLMLb
YnUhWnrN9dOm9fY+uX4xCkQqYagzwlA3rVmnu+aLc/kbwEJuyUlZDQ871F2AKfj9
bafZhKvvdKFGc39fiO6Ntgpw5s8l5k4xyrzPwU/UzZ+WDfFXyZ51Bsfl3HO7R/GL
w7OgMoTCW7fhINvqNK3HnP2xFmokSqQ5XCaZ3IdCWhHrsPylRMwMaGVhGd+GNvWN
FpfDGLZRApHQG0IVPf/yD8ZcBxL8Cl+aL/fhmcQ/oIgEhRJGE2BjcdvC/iSyx5xg
zptIqSZH4LRYt9o92xm3BFJiz+BUZNv+rg8GzrpuWyvHQl1Q5U4ZbUKt+yAd3EXM
wAGjFz4wBxHknrZA2bElzMMjCaxWxt9bgd3OpzceWFLJN5uqqtKenRkD6kyeE8dc
KpgmJ5STikqkQVrf3gWOCgxel3Sy+wmPzmcDODT3UeSRy+/OQgnx25HtCxOJDyeA
XjMliUcIfWOXQhHSiFU5YqPXn/nZl6L6oa1xaASeJzfKvN7Xmye+zF6PO/x1SKC7
rMyUW6ZzSKpXU8ZfnaNOdulpNGBDmUFBfHMDjtXJMOyhc/4s/aSDW0toT64a9FsD
c8po9deudA1WDyQ33k9+GBikcteFZ7NooyqzWnPMoDuZKdsqQ4mSz54FMig/tJzm
TMwuvi2kvEaVaXP/dh8QWYJ3AUTMT3zExAuaZ7TZ5pptXGpEAdJCp87MfgAo+a6S
Zm0Z+MAYrQ8dugUq+4iFPEEFkyCoAbMx4ZnmykBLEDMOSLJdSqP5kD8VpCwocFpH
P8CemHY8mJAzoO9CydIlIKC1xvo5+8BZk1WS0CZ3jEB7YGT3P6nYdeZw36uOfiw1
aaXJn7ic2Ny0a6Hvw/0m/4n/XfGRJoK2ydxb4Of9n9czlBs8eH/9BnGZ3kwkOtxK
7bC4glQGdq26ERZuDY4Bca+b3LPctPcx6ikAo7EUWMDymMH6uykr8DM5VwxTY5DU
3QdI4ZT5sjMwgRVMqMYaXYfePeN/v8Toq03uWm7Vu4aunrAMAqahwoVS98k3O1Pt
q39MIJhXcJ7nrvv0SfdLgBwST7nrw+l8YV7ZeS26xRt3tKIWZk9txV5dgCaN5GCu
AbN9EPrei4ce0G5nMLnK34GNAzhhy1/QRNf/2nrbVDz3MQiJSuf2nWbHB4wKFsVe
5CiCQEemsfp69vO/F5oHvrmFP9bDC0HNFcIx1SuqiwIKTEytnKv1YQk5uVAtCgv9
xsFxDRslDtoohaPIDSOG72YYS+MkOyIboEtDu7HQPo5nrSVRucj0xUFSLMYXYbNg
HK9rd1YxOCh1lWxZ6rFbF/jo5e270ozMx7/5j0VAjv1pCLkRbslwBG7+NohwbXIc
UVRol3jo3om7a86GV29ccyD1yPR37nC5aC/1b3IAW1T1jE02H7RT1N5W3AuemsMo
Yuyjqg169fQD/SK386WkHuSdrpiYN5P5tUyF/IiYyDplcB9U7D5Qulp0dd8Yqtse
IoDfpWawXmikOCg2omjL9ez3evgsFigfjkJgt8bmKYLH5hHd5EwS6mzF9b7e1RlM
Xd4JJ16qm1DLyGN0iBdNZegGrCASd202OHUgFUOxOY+8jC8HoeMMXmgUEw2Q0/z0
NkfYGbs/jrqK6dLvYUPH6Wk/J3R3P1W6pjPu4EvDhvxfNa6vHiTDZfuCOLP7kuZl
/zi9N7+egdXa4ywiniqCprQLm+m0G7smDeMCezKcGIX0PxHT0R9gwcDKlbWEbtuJ
g69gKL6Dq9TDG12d7D7TFtWAsMPr5ZQubD7yb64GODlXU0vJ/CL5XjOlodXq3Sph
itKHBmmRSo4nTDevBcfkZKcAODwSsXM9e5airsVB6VcjeddkZyuikHbdD5wM2cSs
7X+zu8rEdwN79WjigyhV41LxLCvx+k5QMqciwo+VWxlUsc/7rXPR5F0r/bJQx8aH
eTghxF+zfmGY1A/brlJbmvO1XVeru4aYRDOW8/NUejC0H2rIThqRYz0l0AY6s4/l
C8U4UaGkdcJnW30JoCLGzzj52oslYKWcYzwmM+Xb4AzeGE72b27c5w0doE16EU4s
EFIitvT+hEh6wbZkHrZhqD5KePSnkGxckUpgkA5Qgi0sHPI1eAK6Lv5Jz/+gM1id
zjZdyAqsy+uAIiDm8nwuLPFZPR7GmzzEY3b+I306D7ZGcPQ5rqH1BfydUE804V7t
WbY2XbnpUStp/OWj2QcI06hwK3Wg0ryOv1UT80EHz3eoMnDaERWnXAUZs8ubpU7i
Qu4eQTDprMU258XtLNHS44s+yIj8Lf0ZN/o/dktZxcBhy+3rPfIAO0/3C/152uSi
kUGHe7ptf5FahuxU3qq5Qb/qvpdeWg/ILYTh0ENPpKp/VSbvrD5q5BFmcJVwUgV4
FwSqazRnQG2QH1bgUFSO5miqdyhVPzSHrFiCKJblZS3It0c2fhiAbPYRMC+oTpVv
sT0huf9hcubIXJtr8ZHan+sarA40l2JOjAdBjKM45Tw56kueaLEw7oqvT2P1qz62
UWSb5NDPThyO0Ty+HBURT5a4Qv5kqNEw8diUiVHY3F1mZOZBQ8XIbt4VBqMPUBTc
FFLfsSP0aGSHJowzVOtRJzQhzq30Ge4cVWUcaDKk628fK93PMBo2IgVXG0IEnDBn
aBcUQO7Mc+lJGkL6nIqg9SYDmmD7YDV/ffnnOHST76QqVnDU/qrA7G6MaD3vyba1
k/XgeoxY8/WFgmg78PkqSGewmIxsL43pMOjDzJEPkOX9nkftwQs3W+imC5Y3t1fT
ZLgHOxDPOqa2S2sTHR435KXbbMxgtzoADoMlJEYYAqWD0tOpDRrZQHFH6RfW+VxN
kup36IowKaeUdRnbWzSxljg13EouJnsyYI0hhmTbVE/B38CBzNeQs1NG9p1zCino
FYbOhgDK1Spd56knWxz3IXMtr731r0UTdb3ISPwa1uR00yUdCTO1v0MhLzo5k00w
pC+ey9XiUFwkxa3tgOOmFWgZ9YrLtz5XRJIUvJgWIcc1Qg4L0vilXAs8qnLvJcEW
IAZVx0WtKLPs+CyQnfDMU4xXaofB0i66WctYv8UupEwhgVnu0WxPwreMysKnCflb
szDEtL1pQFGFxLZKywrKd7XhhPhK7F67MNjBGJGDYYpNQCXEJWZt8OgLy679WIRW
Z8GOLhNHTR7p2gXP8Fd3WMD9+BRd+LSJICPmkpi/9q7Pi8tBae67uXIqvLwreo8u
o6Uri15oucF0DxF8xeSCpaMKXh7ONuWayOLqArwCPxIBuQXw8IPhLkmZmsk8EgLX
iRGfsHz9UTFANuHarrZHyaNgq04V8EUWVPig+m6++/kGOtKIj2f8AeEKf4Yyy/hD
cHREDuw9dKBd1lON872S4MwmtXsc1j/DWaiK6MAjMVz+hy00zjds5sVnSubV0SWS
QDWTMerQf+qbt321/xSZuLYsiERNeqi8I7DlKxaEV5HooMQEgqvFp+U64KYZSHqZ
F63jy+as9V19xlI38zfZPIX+ShNObOkqcM5M4BQEHHQcISIkT8t1ibomfix1Nqxa
U6xnew4lY6W0IAvDkRVBNctCv7nHFnJxQ9BK3yKkj0xHoo6rFe4Osp2lCMRrxt90
Uxqyat3ghnwz5tpbcA9ZpkzpPF0wKvIuljvx+KAeujZCmyIar7zjl+3ufD9lSwyF
zXGkw6mNLNMKIJYAU+ziXSuSfBTx5eJIoBjy8A3wlRSmd8sSHnifBHPhnqFhE9T7
nSWMVVAdLZ2MC0VeKvaU2qElfJ9n8M00+nHpLqm7H25G3j8dLgYZADTrOXBwQCSn
JRbJCzHSijp8/H4kwUOX4wHSKLKO+pD9uTyv65FLDvdsaHIhlFgb4pLhm4udHbKt
TDQLalEdez1fdZ0BOfhxqrIkk6alVie8gZYbFVcRs7xxIHAQA9crj0+x20Km8iLI
x+obgfh4UW5zeVicfIRSvbJNr7lblu5L45sSTZdqFNstkq09hflu77FpWx9Edshe
luunsOBa+YAIFzQ11nTjrh9YuHMuC3m17iwPpQXR59XqEPPIQYto4x5UxY/ZYz1M
beh6y4XTM8ww5mdiSuDL32QtuABNzvVhN7vWqAnRwxA9fIuGWUBo0P2TnfPTA9Qd
HXG9imM5CGVP0emhBuHlnpRVtmtqWEtuB1dj5GfEcPNZxC8OCCn95GiLjA1u66WL
3LQO82yxGq472uR/gjWBYUEz5LeahRTVgyxqjjlandOSkFrWNPl5nNJOLgwKjuhT
kOfrNQj8x48UunGq5Ptw02DUQL2ROvtAdybwx60OEZaWEE6lJ+uyJRc6a+kO6mKe
o83T1fReAmcmbrIwW1XwAssHIvRelA20Mw4xBSgRt3RH3s4QE1owb0esIb9pzg5l
z4KyQ9rhS4oLM94scNJi9smkcMCeMY8qLM+Cn40PuEGuGcHs1k2y6RsE1bWxCUEV
QlEkWkuaxRNX/qfU0ip3jPZbP5HtS5VajLjZUnzcjoy86y2rmE+YqYh+RVfJfZEN
ZGNZLqi36GMy3KYRgfd2VsVdfozQgpq7Ax1/pIhAX5wOZjx2ebm+MCFJeUlF03mR
IrEymsNWcFAskibd566ndY3sdbAWdsVsvJl6pu+d1xTUcw2jQYs7MJ5+2EGgUo33
odV/Bp26kgpetKezi/DPLbcHiCuCjQurgpFSk+pqZNdyMcFB9C24HdPYl5umBxnY
JW5+MS52ig2ad7iYGrj5ISmE+PLoWWrr1KNoTnbhN1bqOQzWehB/GIoR4ze6QXtq
FAeJT+lfqVbZPbGdMwRMyUt2FyTORNOz3AlWpfFMdzT+zjtEspkRh2DrD0ylrs0L
aJpSjyR/FopFwZXuUo4IasRKrFqk885YPygS+eJnyDBlhCbakbKW/5J3W/z3Y6b4
8xbT1HjCTqYmhSNssKHv5fmXwIyCXCcyvKoMnFjNHrcj2l2E+3oLyoYADvveWTLH
BGD8XkRoihAkS0sWfSJ8yyWIQoK8HStiVFDuBBbMHLFFgz2b0HedNU4pDprFGh8w
c1ZO984N0N9alqZPuxCboTMcQF+WTa8zoscWb9cc+KRaWy1m6eYNzk/JljrqPuCg
YosZTjS7kNSLrhPKpxlGNPaSrDNoITWj0B6EpPOi6njwffSJW4It3CtZFHLjK/A1
2qVkGG0Pu5NE3o6XNLzqp45FIOlmLk5fcj1Hd+j1hesnaNJOz/5TUqJvvbPqtIfP
vnA18uonhyEZP4qaONQ/cgi5u+576xBG+m0PiGm4deIvXS1+tnZOl7Bn6YgP3JXq
pk3yUdO5wXV13N0z2/Lyf/aJVtfRFGFfVS8ka21+eoGyMBn+iQ8BijCnuw32ApfG
2s8dev2nkfTW36BdDuGmqGyG/xyN7djGDQiAeLoKtKvffh8LoZdIoCJW+QOewnkL
xSs4CQGWV94UNrSKByp7w3zQjkyULXc3b1grr6uT78G7Mpp1gddVonACnoBGk5wO
Pd2TDB6IhMh8upv8lgdK5KVs/70uMDzYhHlapxzfiHRzyLsR4ah98nghWKU/hjxS
K57mELsAPXBFmO52YZIRsaBwyvhnys4LdaMgc7DHE6lbKgdv3+zc3fmkmW93WcgO
GRb2XRRrfPDqia3ElJ1Xhk8ErJ8f4i+2tllmWp3beau7fIk8QP0bkDS7qWhMlimM
lMTTqgrqQpO6GMjLaA9uMjvrsAYNISiihcp3NiV2+tSPynTzmnpeOYqpNtKJncHF
xEqkvclpWo+cWPPgf2iFFgKBu/leYqdlmkvpDVORTxZ3/bEc1TV2V/c4DAHCYWOg
9vOghtXDLNsN1YM05matQ8TSxcD1NXU0t0TDuXP9Pg7GlR22Cps6uG/RKhcTAw6B
u+4VJ9gVqUWT6yz6OkJVeEWPLWcKZSdEYbno2qILPqb1/JmTyXraR1uUwEED1V+6
ZZpIeL+L0BNuZeSVuJebbO5gzcMXBPt5heoiXyA3R7dOu27FP/G9c6iFnK9GOGr4
3lPWz1g1hZhkgCw0I25Gxdbuy6odRTsDSMMTKeRzd19+XZ5A1VOAm8VB2r1M7jee
aYq9X1OFdJeBe4Az1ACdTdnuVALrafmkBavHy7+u0OantQc5x/N/xBqZ5UlNWHOp
vRC0GFk992+Z5ItFCgzsU7kJK/nvjWE5aHyVOY3McdQ6YpKPpdTIOSYtaGWC5Oxt
5DnUM6P/jmMeFNuZ0KbRB+euL2E3L8bx3T4TkxZdoLI+GfylWj5hIrzh5SVnSFuC
34eanX46VpK8YO6G3WQvodXgtI4NNpNhdJj80Eh0z/qgG+E2AStVYhBXxMBA90pP
DN81EVNgzWt0bA0ISdxIMRcIThZX+uxFQ3vkiO+mOw1UtB1mSks7Pjl+sT2yOOYq
ozW0hGeP0V7RkoZN8k1TMw860TzYOzn33bo2iZ61I85FVs9ycS1SOWLp2USW2Mva
oQxmPrwD3QA+KtEGwonR0bh/d/E5VllbBPzRcYRK0HC/fzlMNyKhInKMOOIbq77q
yQr0M/kX7hczs3r1d4/2yyv8ZQG358mVqeAs91xJieNm+M1vUNIcIFEtLqmM2fL/
QSQm5d3+/4czjQt7PXt53CrgFY/dH9vUOWA0dsulfk369hvTzI1npxht0TEM27GQ
In9H8Eg0sxlDDlYq64uwdjN/ZwreMKFf3wD1UXcjmRsWjPVUhaxggVieqLUKuFVy
KBFLKRK65+f9rb4cb40zmYmYnmo77ogTPBkoT9a/LAQYjkXrehGPfWILQbbkZcsx
T9ZgAie2vR/ciRCp1TdPxl3G2ejYXPJ9UGBnkiGw4QFlgyl44q0CkTv+3tNbrHeb
G5GdKti8Poqx1U7uHVKIO1Thp8IOpZvZ1mz+5Z5qCNgDfyCSU9XwxHT3XWDSH8EM
d91fLPl/kK7FRM1Gm3ppgyDEocltoGBpNcntRdU4yvlM+gGRpXqGazGmXFPIt0DG
6mEtIcium5Cpd2ONkK04ogjy1TY1TKTRQdkbMsxZZd3nE8j3xT40TjUR6GPoK7bL
iorupegomcAzQki72UKjD7C1JGhxnFd975+goHhajNYEmV7FUF7spInukv8/PKwS
o9k6lx+VYXfrCyuMQUExT8CdiEuDcUAImzOArTr2CTOuSThNX/0nMTAoMpzPvspM
vMwc2/JxNTRXFt02BTETbHHGK7Wexyu2FR3JIQFraJBxiHKlzB5LGqri7cyqbO/v
E/CZfVEIujpFV4XyOv4oOKHj2/opi+MkMyqsKg4YCwWvoQtXXA1O3OnAeCrpyFM0
JDjs77O4YW+6O/4Tl0ukRQH7lnCCF30aFr4DOT26gydUaWXLj6RXlMCSThfU+vIE
/7rUGuSGcbimWudP7NsFqOohfLOJ9maYPuu1KqS//Vsqx165QFkCK+9fEqQc6HYd
rk9RkUY864XJsciLMalbBtHGtfG542b8rgHVlU71zC0SNQ6SgPPzKK137ym0c2fw
1KEZEFXoNY8ommQAaIi5jQITbh30wK0jTq7ZdsfAMYaGOYwWmmF6y0MGyX82NXaK
38S2J4NNJd97XWbGAXA6W8DuvgAFqxXWmtfajUAdrInrKO62zqSOHtdq9Ht5HMcQ
/6FUt22l1llmwe3r+6bt9DwY2wEyH/Rq1+wJjfFGZ5xIoBp/gM5NLK4VcAlLlNaK
qJ7Bs0qMMPf+Vla+g3bDTFGstBIRn6ofHWLPYWCGxXXE3sKc8vPrWe/njIt6Xs2K
WmuVHLaB0bCS+UDmTNIhzZXgS/JwJHp/qtAOhdvjKFynAH1uvmV3joAux5uIQg06
9nuSzyNqdITv77TfjGUMWQlCKR1yhrlKxi73sI1xiz6ay4pQuJ2Om4936jOx6kZe
Q1dX/zei/urvgbYLaJgF0uNTrfRY009HVhiDVWNZqEaRtbdgzHF9J/g6mEleC8wx
uxWVvCEhy0Mz+RudywA/QvNHmskXvTiY31N6Yn2MXBp4XFRTHOAe+bS/w07bDnYG
5CCZMely6REZ2lG6cewuVnR9kGNLZfRwDqT2IFrOqkeClBDK8kNwkz8h3UYytxek
9/TzXGIqAnoYkBwu4H3XW9j+FNeuthLKWgb6d6a1BLvV+bKpfz4SX0qzxFbu1oWw
7+bRCdDeYdTxilt4BzQtXYeMsx/jSaj1OvQmD6SYbMn9M8a5m6NgPT0vBG1ethra
ZpayWkSzYuWQpZISHT3uYwDDVPVYp3ZlBFv6Z2aphUgPcc32UldyJy4u2EbmJd73
qOfGukqTkI1riTpo6755ccqhnWSSR24BqyGrTHyPjeQ5rIjGHxlp6RYsOV+p6fyg
Em8dluIFsz8/jrEDn2MGKAI6FPpIvFtq1MxhwJ5RPAedVuMa6mH44aCvIKGCbcZx
8H2PANDWcE4dQGgF74pWAkzRFPkDcNUuys6BXU6K/Zt6zPysaDJRY/Jcr9LVdNvv
ip0s0oBt9mnXsmJmBuSFUkkqFoeh1+YLh38LZYME42d1ywkK/0fJugW9TvgMQONw
/sMvGac3lU7ajEgzMCKj66sGhUZUqZpk+HcqQI8oFG/q8CXObKQFQlmWoLOYfIKy
KWxWgezXATDR0HIWQKlW5LMIn7SigB4oqu/JxiYHexzCBd38B63S64JAoEBWuG/j
Y6fz4AbGIsRzDKB9R4mi4YyWw0RRE4O7mPE7OsvDLhTol24axgrGjEt1C8Iivox1
oHMx8JbMaDaoLjLlmPO5tInjYIxUodWOuYRFielg2f97L3Vv6+IDweZ4tN6xi0eS
Z5eHSI/QfMfMRvizl0pyVvXrGBYYmOriEetdA7fTqfXCZ6raXAWx+Arg/+R9Emj/
VKwaM1krnNrPG4UCUvNFwG8bOfoWp2eYobX9bkdedoIOIU/gc+HnCm/A/iGoQiJq
O+momXp8xRCRIWshpyWLZeiRjU7H0ujlR4oVYfM9c455Q5Vayzl6wJnlkwDinfgw
WFZHKauUbtUgw+dxiAU5LHjQj2r0TyaFHORREbAsERXrSH+ZpCX6tX6wCKhELyEV
ZYwRWOSJQ4IlOHpqMes9MK4K7h5F58yrdaKs0SnJw38VzdO415EmTuh3t9UWHfbR
Z/FHkjdshe6NoYCm7SG4KyVVGeF/d9GNz8lV0R8OASEJ9qdOmg5GGO+mZEySjC5J
+DPiEmkqjBIN+DVGebRfCRxtFE1hX42tOD4Uy+3D0bpXwgkRzFLvVDIuNCmxNLd+
KyJNncXQf6iU07XFAhOF6S+q5gr14fMQjkNoQBJ4MwB+JF1myRjRrGy1BgLQdXyK
5utSqg6wLed3R3cOZVHLRsPcHRJPsOF4++hdaxP0Vrf5B/MgBy+GZTML4bU8BiXv
QOUAZAd0j8de0LOWA719RALnRCu0bhUg6AzJnvPIX5a9FmJ6nSoZDb9ZH453rVHO
mawlKwft1Dx3GLcrucpJ61P7I/ixBf1V4lSjKi70IJ88MRPHTB10VlSxhUCxhB6X
5ibMU5ISFfMHXafbeiIEEJncZ2toplvHd2CfytMbRofR/4xaDt/EiiC5I+c/pwgw
NnHoQ4siawFLJrZbwy0vS/N25B3mBUBO49L/EnGXnPPPke+8JXYVknlK2GNfTSMt
Um4PUc9TtznjVnoKJ3skDmofsqVWqbTi7vZ4KyMyOQbhJOAzEPCdwRqcmHuVUUQ5
T03dJfKKmSW4kddYhScUkVon9mn071TQs5YdJaS8KV1wA/0in8c/3F/emJ+rIJXL
uVupvtLWjZEeQ08u6wwNYue4LjDzVjWmKcHRjxQ2UhtD180N1C3o4YUdQ/6tUW01
8ojHoHdeqBSBd4uXRNDog6M1fWvehNN1Lhz9fPoC3Yk4zyry7qBduVBXYeHu4Q3V
yhAUZK4ewmwWyVattlm3VFZv5slvNyaEQ7tbQosq8qB+PZ1tnUBYXuQcyZKnv4Rz
uULk2fhZgGQHuPhlJKs8zYWjrLuwqUq4m8opSExLeoxUvVdYtOUQCW7O68zT9OoG
YGXP3D7MIQh9E598mSFExoIKYPsksGrRHB3VjSUJV1I97V3MTBKwCTTzQZpzNqxD
zWaZKO1N2gegYeXseasVzHTxd1R/y/KYREIrotGOZ1Qm9yQPkN7SrYDOcIM6RUv+
cK48kqJHzOzPB04670q/gogMfmKTpDcYP3FhGgTABCWgvFq7qawxjiq5kno/d5eW
ua1I9AE1Cx7nwsRRpp3qxTf+yb/O2vZNNvJe4Sh0hZ3RoF4ku+X6RpvIFsmTaNnv
kZqaLs1HkmrJV8ZGc3g6gmEt55QUpZ2+/5frQ+F0SLUEoRsIlJnfVjlB1c+L6gAZ
ZK+rXAp3SCp7xYZt7781PZBZVTVNmkEyXoa2+fZNMUiZfSGS0YtcHlrJahPFoNdH
MWaugtq0mmQ0e6ZEyK+9mNWcfM9IromzTLFztagPpjVQdAk4O+Ls2I1H1TNnyt9n
zy5l9ENcxIwTFWHd2JkC020ez0sUnk1k02nrNF6dSLr0CQJxqVCIHKZlTIcCpUzY
X/zcrmY2PGbCErD8RZIEZsjBNVODAZwgWNeD87L3JjJUYf+p1gONQK7tgTcarf3m
FhIbGs0MmqmBH/q6ATBefL4HLXTK0HWalpNjdQujc/EODQH8CwWIpM3pyx8Mt4Xy
2v+YjxESoz3GOuxc2WcDu5K/IngD0g+2gdymLsTIqbHPVy+RS39YjxUyEBUaD3If
2jW1mq2JOEj1H2bps1qv79ILjJhlxm0Yi1q9NaPWWQ/daUyG/q4Phl9oq29CWUAy
78G5FenBowW5tIQOQ687hbTXChzPOrG5yVhw2BYdiyzezvXUReNhj7Aripu9UUWI
TZ33HFuqwMSc9Hqq3V3YOfWdJigo4G1f5Tlhr+eBd761Keb2sL6MhUiUthIr89Cg
thKn5n3gxz9Rt/WL730cW4r4kNa12EYTHv+GDc0tBYmYTEKEgYgs0xYuD0V90R8H
xP2ioz3EWLBlVzw366OQaUD9qP6/+ZJHFzBMRh1ZC7/UQpWdiADq9yEXJBJxjLBG
cB4gMCWunEGDe+0jHWAs6MvTDClduECNmxjEsgYop7MJGlDZCTEOakIZiblbmZet
xEQq03M6nwFQWeN61LyHBYOyvISXHSDMeMZ7qD91L2QF1fdQdqPWKmFi4dnYMjmz
HkwVRisoo2rFLUf9wdk9OgIrB9EQsyOuFXdWrhgBVuX/KKtAU+0ONR2RU4rRKE+K
qeNfw/Ov39bYNM3I6USHNBR4EodtrzEQIEEN8LJuT/ElBomzX/t5bfuKQnFJiIj/
a90gDqf8sEYhxy8xzsgBhEgW/SKkaeUV6wpbAlYom2NzYfO/Gr4v0Z8uF0NGnnSu
Ze0dFFrPTfWDsKe1fOsZZbeGsAD65vL6GtJzYCEolE5jIfnyVS0TfQU9mUZRU7TV
2FVDFp9krqhIkqaXLGgf7P0uuCcXuGo6SmP77JMKBaP8+P2iii/DMDmPcEskUdeC
E44AbQS10tqDc3M/OlQpnXw7Ypf8kvBVBc7Kl8utCMkEwfvflmcBCIXu6H9WuzXh
Y5/EWHu6RnU+yeB63U+zazxDtVH8aEnz3ptznXC7klfU4ufwwRfhBgOHs5dbOwmS
qJWcRTM5S2yD+l0RdcFCiRzkQgp6RoIgCFBht8Zuoub2bp7EKdTU9yU+Kp9lAFmt
bv/UXDNOyagj/ldOD59NwxCx4fvCi7NQObg9WDs8853Zdk90dOafGZDPUMrOI4L4
vcEgWCAAN8lCqDzLimlpnji6WccfWgtAqFPr889+WRrHzZ3+SgEK4ZNcqzgSIV+/
6kRjY/3HGs3zCkzHTvp85TvOe5e1PpRX83omtYCInLzmz0sI09+2bouHSkum7m8H
vzCQJ2Oth084/aFLJ57X8Td0aBGtIVxuDZ6vwigpZPdJYG4u1Nb/k3CBhGlnpynj
jly2AFagBmngiGeO/9Sfgu5vTECDfcLkfDvVOfQZdkpzWSnNJQCuqWKSzeN4yzzq
dTQ//7aYg9EV6BbRIoT3gEVh11IJU1B/CWKYExRJtVEY/pvVrm7nYgJJGmw9ivzv
j9fzZFXrCrXjgkCuadvnSJBFdmGoYcQ15czuYvSQmSXspdxo2weQKGzXbdHjPotu
MHuJr6BAJXKGmSpVJFHGAF9q9W4wcXvOC/dPS7HCGs5rmqyevp9/zF27sIFnkPIU
jS1hgAmeVXh1IXGgBWSjGhPU0VU4qUy/ps831zpX1SqBJE5O3IG53ugCdo0aPKAA
Z+Bm0CwkYm2rnpdRS/IbbG4FTLjmVM8ye2Wy9K6l9ZjEXb72FYLPlF8NCwZV+BpI
uIBrqSBvanFsZu9s02NPq1N3uVzhAm0nuFdbd7AqXmvmAU2X6n4/GPIyJ2NLMpfp
pX9ToFu6NW8E/El6uBTyC3t6EbU0GpGcWq6gR+mx4eCgzdHaocD5zSMN5bhNIE/L
0XTzQtGYgYeiYqwH6VU5X5V0v+uiRQn3YEexsQj61QRJ9YdcRUk4W/4BNev0X5oK
Y0+b1A1omj5Fz9ByuJxUEgZDzg1TYKiorAmz1uMN3U6AdFykMCCukc1lVzxHVsiT
izLjtnHkmQxRdo3WzgfT5iADKgHXVA2x73CJT1zEQvDEZNngG7vePrb2WB1NQiAB
U1inJ2FRz4+B4TFM1Vx4zmrkpmVU5n+lpEVZEGjJHp6YPsQoL5ItE7MvkBSIJfMH
1bICA/HSUAts1Sosk0/y73GMNuQ96FfhX/mslDJ2VWfOIkuxSqiN0KmeYlgFkY77
31SFig89Wvliq9M+6OJMwmm+CGL7YBGyX+qDPi9jh3FzmoWtU/JzxyFh20Wl/uOc
XNNQMBCIm2vG0H4z4QXDH/KAmhxEchmo0Y7BAQW0nhqBj51kBqwZY1ZNDuBY+985
HXAL3io8WTTeu9IJK3DzJUdrQfulTEUUrTcrWT/3cq5fosfSiHRnTurXzCJ1+9OA
w8JMuQIeCCVWlzSMJ4J8aT3TXiIeuaQszGly7A0JNZ4K42qg5IW/4YsFYsSWy6Iv
LDJXLDKRaQU25Gq76Z0jGGGs61+mh8PdNEHhtvQEI39MkLElVf9u5Zzez7DW0o8z
1GC+fPIK6Z4MnyGovREXAfv8n78zZTxjxQez1Q1vUFQkplRM0Xgg370ojkHePq/o
AKggJ8b03in1bONUQaaSCHk17H2GwW3ruJQ54WmgFciEvVbigzrWC20a+GzRHw0a
/rndLmO0LT0Gp1+i0QfSHG+GbhCCz08OiGe7uDwo5ZdzYFgkndt8zxkkeog1yQVv
kqdp03NXYkKsj1Uk7pAIKMcrDi/4UHQa7jsz81wvJLVw9CPCdCJjLwZiNRoCWWlS
UL8JEciRxE8RQW7GgqNabFUNUY5VeVvCt9nzdwC8IxAuN/gZVjeH5RIc4SIgihgw
dONpyQh4IWPagv5wjGDKuVdDlXIAGJmyf4vWQTjIt3SQqzXAmo06uYv6QOC7BKcA
yJg7TRRDNQpynmllR4wWzg00o/miRq6MFJp/U4BOIX+JavN34TuSvRJO4Y7Pt1L4
H2oRpuemEFiAx3c+mJQAEJrj331hbjyjT7bWpEnUXA+ircVZDisBB9+DNqqPDoor
nLHRAMugqmOCFocK3DVuXByykn2Hy2JcBeTtO4F90JVUzhRtZQiCX8nm8gEDg8Ye
blyXUhFEXJmGbwCLQGLvv9VcBOqp4lHICbzEj8KQ4LCqkByCyF0tRxaCskt/1+ko
ITBEkXfVickL+z7S6t0IHGR/4BvpqDTDS8a5m7WK6IeVQhfXCSmg2ugzoRNBIqoh
hgCo5AU0OctRlFx3OglpIMmbfSMdCXAC0MY70fRDyvjTT5qpekezsxepvDzrvqLp
N+d6gsUrWE2x1nd166RKOqRsBtlrbUrTk9YjguXdjiwHPE2duy4lexy8uieLWofL
HiDwyiKXrEdmm7RTHWqOfHjxpuHQl7hzu9GBMBuJEqxx1j2cWGDbGLxXs4J1Cbp8
/EAH1FMqL0WIHedl61ydIT/v434WEDTVMNvTHYuOpNqbvoLFdxYR+SWF1lE78uBu
ZKdEgLeTr0zLI+0QmWnhgBSx4AzKUzAoFS5rL1jKga16BoGJPlnggI/zQEOI21JJ
yY1sxGKcAkFGgl8BaeS1RsYIoWWQgQhq1VaLyfSnPa4dqzGWyXpcuMCFjlSsiBLQ
2iRQMHfLMfkx+ho2vBH37PJyy6kri3RBYXwcIJayL+8qL+9eYi7XpTHCYm6cYvU9
Npn4OpometmEIIWcdJupLulcoDgOPbLZFLC9U0W7hFc9aR229BGi06jVakOqNrE1
02PNNvAzSRFYT4ek/YXQlrFwE5wUgM3a5Mi2reqQHZ8h9fnu8K+C9hg1Xlan4qy8
ofb6dCjuItiUAqd3XV2HM8pIMlXTkMB7LFWBBe5FplwntQYcQCT36zIz7AuBDdaO
7eNWYC7Wq+tO6XZHPxs2FUTflsyrOQEc7Hh/scDPIoT624c3i4YnABus6yOAWZzR
xMSCVBzLGl8mHDGKcZz5bVzdyigt7tj1CW9ihdHsC9YKFrD4O3YawNeVk4JmUc43
J8fiJDh8MDy8YfW58ZFn7/7Z8XwmzMlxLVyQpOAzAg/z4BTAzLehJGathD7STaeA
sARih8rvTcTLAUUxh8T5Ga+SpbhruAW3Io1sZuJjJIqPr+VYO8dDOHlczvyD9oGI
rRebtmJ2OZx130qZk4e2nG0U35ksvcudauEqI53jWncQ2VHIOfMIXa58ObRn+b97
OdwHwNFVfE9VGBhurTV5YGMPoQKUCWqVBPS+75kZRG80SU0QGE4RlWaMVRu4qSLC
je+0IMPXBJQNZM2GjbQwScmVlPwtUFs1PhnyMkqA2justB3NyWpF6GUTfqegyyAV
VDlL6XgNlamntYQuPgvGT64ToyOCdx1sT2tbY6XqX72W66X5TohOKmAmsNxRZJ8B
3URSzY6WTtwJzoQcoLnBbhKkdDRZRFARCNi2Yx0ZMILBMjtSmxG/K6IgOmvpPFxr
rsQdQ8khVxtX9njTFZ4beY7aNB4SYbKu6Afpknby5bgu6a6mXo6YVOayMxgGQQWo
k44zwqzTJ8fMiw2YinG0ZiBQakm8D0undamOrzzCtyRodVArHPiVm84AAcwo1Szx
hmaESgZZ6n2rQ5W6K7ygW8MkIaap/Wqkc6b9MTgS6HjwAnUsKXoOQ8+w1C/bNWhO
FnckrDXKvIeoX3oa7hKSOSeDBnNJDfq/U8O3B5ISSIkni1MIx6EVXLmScfd9hJ0w
K3TUNXEyFWjCuBfDMkeg4+djRG9l1CG3XK6LLRipqCeqQdkSrnUCa80yXCd81lWn
vLJ267JyL70cHa2cZAORqh/UnWqXmRiSXJKjScQRbb6KMqHHoj3Mval7T9aMLiGh
5pajXgZtJg2Gfw/Og3PtvzrJgKGZDk0pEmgVjzrgOiT4dEzkRGd25ct0anxTc4ZV
IhjNJa6YNIH9uz1IPX8S8+gWiwWE181s0sMT3VkyJxWLLio4CIPZb0rali1vjP/2
reaB+RNLWGepKf0l5fYcRefOoXIrxAqlPObONoZZ3nVFKUGmdkrrhXOT/azB0yZ0
U4cnWkirvKRRLa7KeWOdjlTMpY5Fh+rSJ/wCTOp7TOKWbhDBSE4JRrquDo047RIK
M0eRorct/1cq2ZOXjx9b6UAKeE8U2tFYKOMy4ctboQK1ryZ0DA2VHu8Ov7qYxxAg
GG63D9te6tLkBY35JcoAnpki37HELuVq9WtMl1zzemcFEIrflVe8yPv5KaCxU3GY
JMYAHo/2Z3sTpckHpbyAcIDq28ZNeCYCcgEpWML0yzgMcgWClo/qAvl4uVIbzHEV
ZoMqbXucPHAjyORQvyWqrILeLZdPAA91rROfU8DcrYU7SIwn2onvz3WqG1ZnLXpA
PVTaJpayoIgk21yvEsTRZpGDX6SQWfuLeY1Y+XTL/NhkrYUyuFrfWoVQI7oky2Pt
ySTHExHB9Ir0Bf+xqE6rWb39y9amxrXRMXLkHFuqh6NOMQ6kB5VgzHKbQRiYozcL
4v+AI7u8um+BU8Q85OHK5sO7ylAdWtTMdB1ou6EAQzme+qAP13Lft14RZuhi0jyX
zM/AIuC8Jrg0nB2qNeuJMDpBl3VNyBoHpa0L3BrzWsNZGt+vVag2k/RTBMZJ5UGK
+Zx/P6uW1k4JYF9pkT1/tKHDer1bM6zeh9AxqxZ7Je4zvlF4WZG6NauXvMkTNGDM
3MszkLZe8P2CMHVpnw/7k+J7TbHIGaPaBaxEY7XYo1W3X0hzxquqE8sbwp7cnUQV
xvSSg3EsRCXaeBymDwwZOl5cR2rJGJlUUYmMiawpV/XpJkGZp7mqcQ0ybGDQX64y
PM6sPVV689SRkEI5+oJ2l1swfd48qt0iGbVtpOvwR7MGmZrKFQMOvE4Y7abQfwhT
5B8rA27qP0kY5l7GFtBK78xqorLR19B/Kq7YyyJtNTvBHUqTIdBWAShc3EKo74Xp
a7M5Eqv0wU4LnqVm4Gar8shRocXCGy8h29EtCtvWEpi7I9MDLYYEfl/DKXyIdvLU
NISMR6CIVDyYEO0PN9MkkJYzDlrNnEC57NG/X7AHnBq5y5NMsRzuE2q8h0UWsbcC
CWS8Y/GaExsxNUrpYL6zIWokKd/2k6625mEMseKbMANyLDlnOyp97j4gB2t2ZWmq
V1A9+BqgjXj8ZnTTgAybB+aHVPG2D857rfxP/av/87t/twno5cfB/uTScpQgWbAb
azO8SzELLS2hENJklcpN66xssdIhtWqPYU4KMXzFlP87jKL3ZuCFNQJTWRhWJk4b
cfPELPeQxYzX1uKp6NA0Dc3jFxvX98DMxG7yYRNOKbI+ro+Ftr3vns89es7XS7v4
NhkalrI4Vu6IrTzFi0xbBeOjrfoz16mwaDzPY9uoy87jewGh5XPW3P3qvslVlzBC
08CnXeh5m9Ls8abJ3Ww18H/n8I9eHlizYJ+Y+XO+R8x5W5RgXOjeI7k/86obP88l
sq1k84/FSEYyZ+SIaVBZ6Iwtk9Wd+dEdSfSCebFXHE9BuSbzuY+vwidNL8kv6uDc
i83gcJ3vXWkJOB3N8UHrde1++80M1WbUWSPG5GhPFSyq650uQQkFWj8B0L/BNJ1G
kreNLSWLfCJC21FESaBZXalY1JdfXMYfzvuJcqriPjcSn7/sIWRFCfyxwz/H6NgL
SDiz5XMBs65NQRJ49ncS3dVjE0ZEQXi3F+ypNYIPS0F4artu7O3rp2aPKdX/mM7W
uS2JPvyTZxBd3anW/A2QUkoAWYnB2MirE65mURngDFQY2u5KjLEXDftkDrRy8vlH
ROYhrJtWQefMSLYS04rfKmjCzATcL0ZCsAWwTy8v9Ppl+6bS3oafDTe916u037SY
iTChccj4nS4npm1l99ShRx6rPFLx+FzHIwb/0zK9hAz+ITJO37h1WcLcqb52YL/f
1QwUWCSqsJ4UG4gMqD8+L26FmRBXNp3vOclRrXv9UHiPpsbqujZxLr+Wrc40bYco
4hufJiwH0K1RBR1vrOL/ajxr3lLzsD83/kIhzAsPfbXAHAff1n1R6k74dp0Z2XiQ
VG1pkvRgkp2mSjjvWEpyH8ThXiACnuorVHHJ33dWn/dP/p5Chfzoh7UOurAiwFFg
LoeiHqr9QJ4HV/YlqjQeTHNQovgmXqlKxleAbLyvJ4vd3EgATr2XF32lPqZydGWk
iK8J2KI76MOSaa9/2+ozbZ3eJ1fL1ayegAYckr+o3zkgxFCurrv30su7F8RfVL5Y
pZaTIRyMT0FBHoBxcQUq/n1L8BhSTC7erSDVCVFMnZsKCB0NiJd72ctFu4t7ap7s
d8veEFZeJOpqAv/WdX4OqlAesvdRcnvNyqVaaP6uytLJYYMyvr1cRRILPwTXjjBC
Ht+AljwVoYEHvmaKwu8k2oQGnllpBIDlOMginCPfhNIndcKAuDiZrXaz5O429Jsp
3wHg3jAi7lAy+aTmPKwbqze6H5tfkJHSx7edRv5xrCddX9PNQ2tqFrdSAnw2k6ue
cvwQiybjIf6TUrGgig/cj2Xyjl/lUMxozoaLCAnzb5s/Fga6A87F6KujX78sTfdw
+lQMpGUZSdNYrTCixKWcXmeJznvPPZJrRv10+6cAdqlH5vWvMHhn/XZYH8Qv17OR
77oMTHlKKnhfBBUzRTCVhJAFZNNJOODisTHzD0a9l/HLHyYki+DoG/FggvN9Y8fe
tFkMR0ugNkwJpWkR/PIeeJLio+XrRzBpHib12jPmyg7V0eQyWP0Ou/Qru/nYCWe4
/ApHqQT/WA8lQeftbhR4MfiLP4t6YibetLn0MfVT927XegvDtDKb+/dWe28JT292
5vCcVbFgV4k24BFaJ5gRrH9y+iK61dMK/SXJQNz4zwGQNhIggJ2H1HIRNeEDswXe
bMon6aHJ/4bXteHSd+1SSUl+VPqtlx7fegYvlvvlpT64Jcb6sms9KfL+bHRaJHJJ
zxh8m/KZA/GyrG116ell9pPygYler4rvFwO0R682LPf25I05xo46dD6HNFVpsOdr
Ccfj0aPstCqJtyLYkV3xA7Uweo7XMA1NKhPRRjS/4tuhcQM3pafHbEIo6QXUX4ux
NdSnOgfumbuPeUw2WlDOE1qVJpGfqjv4x8tairgzd03IESRjPWpa2m1oEpe0gjUD
2sapzAiK29uS8NAcSWnfwEWD86jW9OqE+2j6jCA2JA1LQXClnFz5GiKw/klMirTB
mqguBp3CyyF0Z7GpBJSury1+7s3jZsi0xN05VytyyOvX8WEPMMhqxubvN4VqJWe8
2Y9W1DpBdXnEB3R2npCAZkEnMZsbwXAm01ZBAN3a5yMkM2Qif1OflIxYZraFkD0D
jmKaNv5eOFy3xFIZMVhQWnVc4/i36mPj0n7iDjUGcjqc5l4wN8uYE42oVNmRloLu
urfZyYkl9tq8ZlvISaeRZwH7BGfJ+ydsW3aYcqD6dlq3hKGY7UhSNglVadBr/VHe
ZJqFCh83pnzpGh99WPbJSlmutMqBOQTH4MDchLSJ/RWwR0taccMiw/VPvhUAj13t
HyFb8g2HO9OBO22zjvAU+tzBAEn7WkTbnkTriZRx2fEi8egN10VtAjR+dfP4yFmh
XRBA6SIngzHt8tW6SloMbMTbXY334i34L6304FALxNNBwa26kJ9MjEN0P8Eu71h2
3xF1cM7O/J6lFf/zE3ZwtY4zOzxDiWCpJ+zN33jYUa0sPr/FKY0uJJgcMqJVI2Vh
t8HHZRm7+xJV/Ggl/SG3Gy82hI1gadI4DFZSwarwn2U07KF2UudCkmay1bVunAJx
zZGRDve6rRKf+8/PKIS3XC1YbQcsrsJQGljEczhNn/zWObIlOr3F/ock9PCRc7RI
wD3fmmGJCQzqY754En/V3NwXLQ6QuFFDQqAGIvvuHx5hoequx+Z3ZIhqOcv/mqMt
DHFh0zIcKjcZ71OukXNpertZjBUKmCnhIkxsGkmHNFr1K1fn5kXMORKgweFx3zS7
n28lsZgCq8zWWAeDtLLUjREL8r6wsz29sKa9cNuFLHBdLoVZ+TQOIj7z6G7Ru6BH
zt9oa3y0NLsvDOI3VfR8MnWElJ3ZGfaTCSAZfUBTYCDfwSSvdSqcKkpcOMlAg3wP
13ljIMbMSG7uBDpd0LcGi5lj/rzdX91CcbITbFuwENjP1NJ6wCWooFqWwwH6W6nd
mcudWTvErp+cPad1rrIZPMgmXOPZDGJ1Rpq7ns9hrbFoRrIQAcHPHreyTwigutH8
TcseVnaf3o4UxWrVsnfoj6+OEDANps+vIHtrhgkUxFp4phK9Jpc/zQpLupiqiD6V
amdYy1TEyJfQbWh2HyqGbz/WjRnbgO5ljX8EcbhKhwhvOHpqjhfQxCXixneN577c
mehbAPxuOH2owmt21Paax0Mn2T9NIHXZwhzNzgeTgKTKwh17O6NRfpSPac0YEhTJ
Rh/gIwJIGcE+5Jevg1TjzCjla7yGiVEkmazmhg+gGtTU2VZk2NbZnogbCvLB6+xe
CAvb0LcBYyRKS6m9UCQsEN6PUCNtXAY4hzAU17qnmc54rpsLf/dAsMPSwp8Yf4a2
oZEUBtGkHDUec34wIWmEal05wYsThZLdFwhroZqn04Tekg/lMYCzIcsmPoAjOJqU
ACFAikqPBNz4tLOCqb2yLZ03oGeEtIN1jGFblSRLZLgGK7HCYWbaEqKLu2fw444Z
a/+2mtf7Uqr5nHeKYlvjOLNsutnBJ2YxFPpSMEeB2wgpet1+wltuedwyOi/g0djG
HUoTqka7Mf+pyV7xUwqX001NDyt0wE4BiOwFhnqURgRVQ6Hrs4kIWLWCAfe8rSze
cy3GwiUJQL+rkrNxYlNSSUFgtbjlxAFWHgWYMQTF7f567DnUljTQbrLmf1ZiBnxG
B7NkOVVY2AZyxO7bdU/sds/5Kh1Gp4NhV9gqr9NN1ow5VLjtaGumjg649H/vjJVR
EtfAUsckicC3dSfz7FrwortrsQQrH6FK0I3OaT1rhnq6wYy1dAOoq+KpTu4uTY7v
cQsA7kgaNr5jZ8n/ohM5nnbQT95RCn3eOOSXIFi5TtbgiTdAMHnn3FDAFk3Zk9Qq
rd/MzIB3ovX6k90JqDOZ6iVS9UuZm2CbCyIg82cupr35SAUftldHoIwaDis/L4mY
jj4VDNTgnjQNyAjczwul40eShsW5HmTBEBET9av+9ESmFkAtOz0t00jX/B/fNBdx
lBGmS+ZHQlNkU+1MERgOqHtJKJ6sXNnDsG/C+Qbge418quAhn4uzlhdVGZJA7TyZ
TkAmWSxa23DdXLuDrgYbGgBD1j0dMOgc0WhClxX0mhv1okbzM6cH/yoLY9iJOV62
0WtQZuU5W3PboRvz8EaZr69/q9AnPZigDCwL1zyStM4c3qNQLDekoXgo925cIu8i
EhbGIqaIOmqbBPQq8yH1GOaQ4I8JBr6I7fGhBJKmu+hEQusV9sXm6h+8NUr4zWmP
FR/yZ8U3EOkesxd5RgIdN/MTwjf1vrO4TYjDEbCh+GFhohxVbJGk1F9yAdKYnqGI
0QliQo5Kag4SqQ8cGmk7glB8AjPoiWCI+GbQhd0HapSxu/KIOPy8X3ZK8+cJwsA0
Ekbi88Z5ERAfH1Suz7dghYo2OVDfpXjoaqQmfSj1lv2m1Im0KM0G8EixvUKQ8r8X
KPnW42T0Jj5xRrdT3PAzkIc1Y6fNgG3p7aF/RAjthvQBJzcPIEFIyzYpy62q1rbn
lWI6YYdOPEiwJL8zWdQ9Qp33XYbX3tOKAFCx4KEywHlbDMmr9/QYwZSNcP+YXv8T
O4Lghz/EldrPKsIRU2fit58SnElFJWWeXEceltdoz5/TdYJeD8UnmAQXvysKylM1
x2r17NCSBRsB07fdso05oEKVCBRd11o5tCOd2/7kA3DppPYeWl0zkU0Kx4Kymizs
LuWlGrihyMWmKnou43lIqlmTaaGTIQ3jxJ7JMAtbfx/MWA0hdgXJKxT4afqFp1T7
qL/4U7N3vjyaJfeKS845r3lRbeLqO5m8Leha5rCCtBLvdJ3Jat5WTjGpDkhMFa4G
BFrPe8o4Lsldd77FPUyOb2jG3ehfBj7MUP1v9DOmevHPuBapWCyAOcin1KLZkwB5
P0cj1ylAlx0jo7am+LlHHK2oURDAAznNcfgqsnFOO1dhxwyPM0qmgTqVlGvIZ9o2
6/C0Unz6E+uiIHm7zsQX2uqr+oN/DbBrsUGMopqHZD1V4v3Ilx/EQhHtN44h8Lxd
KAgHYm1Eo4NuxeGDRUgEV7ZH8yxPTcoPP6gfl+zif/hLcH4PAjFGGAy0Vq5m8Jwf
wT33KZ7BJaafMwWK6HgcnHjh6UDahHqfUzJO0YztIcO5fNuTr0MIllcWUDvA6g8q
07UJeAtyxI5ujAfvxAWp/GjhmidnVFFIqAWs2CQn0g5vqfI7pC8yeKLd9V3eV8cN
Fcw9HKh6T//KJ0jvHAclQlO86oyZOhu1Y6D8xEZkktedWXLOvkYq5ySbb4FM7DiG
hL8o7id9quzqRoOlN4kLNNWe/U7yqK0UNl/lR/oimPp6fuK4cRA8kSEZUoF2fj3N
6B5Vs8Oh3ralYS2qggp82OkIrrt4gkdqFu3LaEB3fxXjG4gCqGIeE2GIWXJzKfvC
Zu1c56YGx/+rjPlz44GNyVu52CC5V5ewzgazG/fN4JLqwh3sjfRHkRuRRxblfSEf
RCmTcVK7Fyd+nxQ57AL5G4Zvol0yoTWQzT4HC+Znp+SGFPbVwtKB0YHCupkxTjyk
5c9axngsRNf/FtPP9j60n1bw9ZQGMxKxrDm8MXe1xf1mq7sY0/mXo3yrNh6EyXqJ
g0GSDClO9Ci8u59I1KWIw0rur8u5iW3iI7cpTtaNerwAlwKuXpc7jf6Wg1oVliEy
cdD1lcAyisc0y6GlOGrKiar51dkl6x93ALI0zj0OEFhjc+Xit+ESh9wI8jJJlfrp
OsuQjdm4XG7ZGrWa97w1yzYHiHV3pe3zQ/BhHTya/wQrQqwTN/4naEuq3Spjfy3K
sblSBN1Ja/tI5Fuk8at0epNupFUw6MMJJmTRQIbCjTASvyONxFSyTL40yEAYFoWz
OM8vlStvFO7DD/DMAiFQZSgdzY9k+A0C8sCBt6r2yUECL/+Vsyo1HXY/pbq0noCs
d4StMhlC9TQrI9u4uQ1l6FnIY1DzSKWXWz+sqyOwAFFR7g1sSoPgoZhiFvpgUE7F
pXx3bu68oxOdo4NciUv245AG5ZEzGvH21/5IOF8oW9wCbE2IirS8D1affawjrE6/
jGcycs2bNN5f9IQTuiCSM9TG+mEuyNv1QnljvwRx3kHPz9Jz0Qh2lyRIYa27N9Ha
SJCu5bq+yGDqvqv8wt8C0iQRX2RAuqxkoGTptZzKk21EhXgHztBhinlyecVjL+B5
9TbMDo9+7jM1AcCOYUBhfpEb23MbqcAdnd2guFKveDaGB4WNCWpesukBUR6czniY
yMtXtBighseFtkXjyPlmWFEkaHe5NUXLfyUTEsO1EW9f9GWuCjhWUXoS5Bab7EMc
I+3Bx6R64HMIcvBkj1j8dCQzDNz2amdr73/xlgXVc28a2jH8jm3ZDk84zTMa4tqQ
VdNfAbTSuORumsSU6+W+v7bsfIvlCmtWn5Dy0oPJXRM8zKnHyRB7Zb+2QSJC/VZf
GQQDkTHdDJbfTdISh2XdZ1142R53c83t28L1uNo0cqdtR9u/6d9KiFfhUl/E6Oia
QEk3o5nYkA+CbQAwslq9h60zQjCo44awbfOWysWhDr64VMRA4h0M145ddxsBx11/
3qF2J0gueIei4OoLymUjjf5jOnm4HC5B6jpbIeBmoT7rYxHsvqpmj1WnEJFT+SnM
x7DnFrXv3SPT150M29nbLk5V6n1hmWHCUIMbLTmmdjt/Yd+xhPaLZ28znMY+rvHG
SUyaYvKtKL7MR46c1d0l4hKaTyVrOR1eHhdJbiWV70w8V5OoL3XqvO3xxb7y8Imz
QLlOapQt2H+sl5KWivEdipxHZpUF5aiAeErXfFkIWVnOUtUNyioeLDs+/jktUy/e
uzk9EkEqG6S6XZ/g6ek+wFcexiGdoShVTphkttzkoHXGfWuGUZynWOsQWVgKauLy
7VO2nAlkYiQazBRgduYE9QVfUXBrD1I4PeIUg69JPbt1/rs30hnmNbyiTP2PMBpN
gE25Vc/a6mKyoW3awhyj4QEZUQuxDSaKWWOCTRlmuD6cJhWzdLUdcLGa3iy9ifZS
zlWN6poFBwhBf4dVakJUzSy6li1YsSnRMWf8geznGT3uC0aWbnrKWMExKB/JvMoD
IBy8iUnL8fH9B8NENU2a0ysykJpfwkLVi/RTBVZ5lgrFPcmE2WOCW8ErafS9vlwx
CDAhy1cMfhPmcTWl1QjYf9IzZccfRTQFRMUdjWo98NVlFiLJywZzDf2n3yyRdJQC
+TAv2gEZQTJb7dLy4s5wbz7O0Sj3vYF5foeA6iR767aId1J+cbcG1QDFTB2d6bS2
kbvQBiWUF8eX46b1xLPpe7HFqSxWpr9psQ/IcgiFCbTmHaNN9J3dIjneywreQLw5
7fjbOmUzC55DphjD0s4Oryt0WuMj3HP58Uc83+LeltKsXAofJfhtmzxaqMp6SELa
voPMkMRLcRGY6LQc5dQd+ZeKQgwKlYPXzWhoY3G5JoC234jjoKazaeDIOra+SSyL
nBfhjOx0JXhVDXG+OO9Rkbq2rGROUrA6CwsFahQ3Rw0RlYnbGFFdsbkfiwS0uVSY
DZ/wN6jIKo9kb7klmHAM7MbFXz1Zpacf1TwtN3n67mJ7kyZCbS5FsDVXYNNK+qbB
14VJW3OJX/y+ZeIb2NH5pMqSMLXMgSiikZLe2XQQB+j7ts4dNss5MyurPnfyvzzP
YKDXCJz6jZPCRo6ctXTP/dYsXQ8NL1yBRtonUYHvT+1NRt0JLxAKszoGvwLXzJmm
mLjH0MqPhNjv+T1Wd+6VI8Qv/g3cLEBEuzqViaT4/F7OQM1ZAuM6D9YKtdxBLKQc
2/8V9j6wBfHObdDrNjHDdnCRUYfQzuRrisiPhY+AXo62OD4Cxzzl5D9DXouCUt68
8UI5pkyhknv+0KZZL7ciiiHRCdg9JhAaJWgfFRBI1p4Sg0MpZULNvEf1zzIOUdNz
K9nPTsEyc0zBH3s0Lvvoy0HhNJAj6kPtObzQHAllReJqeoRf+Qo6dpPXOV03PyLE
KgaL8IXMSNZaL9dOahZ5LH82lE9Q9GceTWh4uVmhqdAdk1Ir8wk5inKhLPEXsBCG
LuwmfeEepZi53gGmVPMQshAIvvdapxKlxuflRyxDsLNh+XRpJsIXMunyPNJE0x/6
HJdewUlTXOMhtk59ArCjeOlPtBtticm5yT/X0y9CtXal3vcDLTkxfU+vIaIMgWb4
MuE7im2+dPLn+kcF8Jvfplr30VWrw0Hn6P+qcCAspsBpUBVwPE6JJ+IN59wmdXG4
RoST443Gl1+HiK707SUzXMbYtekhxvOdgIMXqaZiQzHOpuI3mzUKufFR4ds/GTbq
sSzTXKu/GBBweYntuD1XaCZo57J7S8YbxdOeqT/5X3W9oH2/nmgCJts0G0FL0wEa
p++Nj9qBP7I4075ZgrB4D9QGvhrWoQ1Ut/s6ub9Cw9Eeji8Hm1AbSLeROb9xYIBS
HO0jyquz7jySXs0vuxNLl2cWBKC8UEHup41cf9cK5gal0NjmwZvI5qt9/G2Ab6ou
qV/hqQJatgeatRrOnxmHiGobGZmRMydqzFfL2Sdzw+kilCubPhTG9mbZY/rrhuWW
Cuzm0C97OSU/CpuyYA+tTtq1U2OY+x4y+hmOMX0KpF5lEu9VIQNrtL9HgKaGJ0r1
nM9xLF0vCuF1eXKdvOt68d3Xfr2zYepSYzRCy9c4VBT2ksctBasRPuqjFeWdgKMW
81G74tsfU7NgySlig6oMi2EIiPj2lHI8YlOIuXIaSIw5S9yDjbsuH+Pkskzt454K
GwFmngiKIDKivSrbKdmYcMLIVJM2UdTxCB7u8qBTNnKyKhIcUeeWS/85Ek3U2ImA
GpMwWAO/Ppz1gnDePwLla4PQkJAdluSnI6+zaTFGFwcilrlBgNf36XEhZ201pxzz
9U/WvrGoHRMK+IndXheA8Dv6nsf99O3kGZJVXsoTOzDfedD8Ur4BvqFwzU2XM3UT
bNqi03uqIBAxtQ1O1P2Rqie53pqZKSavbYOgy+pXwb8Fwwf0xZwfKUzL20o6RUoL
VLbhtPLNhJlI+AcEz9t7PmJtBDqyI8H5Ts7dNZG1jcM+EXI3f57vO58SIoxwplyo
dkLstz9RzILHbQxAHAEdQ6wibnz6yxhzFtQ+TRE6rGA73bR43ZHsYpbTsTv0fHsS
tkoj0UDp3tW+/QAyXPMoZH0vf7gaZTHirnnxLSGjSVx/dPwI9uEw8CeAV9x5ToYk
ECQUYfyDUeIWp8heEz1xGur6ALx5faBbopCcbmiBcgUkH/FyF8C03hqNraoWuyum
J8EBA6g5GXZiH4U8A008Q07UgZgHWz2jnxIVD+teClznxrcZ0iakbADcNvDW0stC
ihQnQFAMDsH1I/H6WsjnpLS7ITzmdbo4seAeNj1FvHbJdDmWjZNDGbCKMwdeU8mJ
YMkBlDDN6Vd0Rj0WYe/MQ9DqTCMRhtpJA+b7TTuBNqHfTkQ3IMRc3ufoQ8ErEv/x
DTDHQEMvc0wKTx5cgQiBu55wIHwvGS0jVAiqasUibAl/3ISwF68f/aM38Zi71t7x
HV1GaO2bJfIFbacEwQP5z8RW/T3OOrVtXFeXH6QlyhJX3KV8/F8pIEhL1g8wJ9sA
8ScTMA/Au5axbL6FlmHP6BZpbLDPl3CK4iIkcgCIw9uc+UoNwGM9/x8z4rhADiXL
/3FRiqO60xykJ3aVohU6ymZSCVpZ6+SdkRPfq33YS+QvsykbXhDh9zAUQqrkvA8n
NNk9va9iWkPBdJbu5D/kptPOGqCK/2jDfQhrIPj0fSQ8SNbvFagkNLbVDWH4+ccv
V0C9Q56T7g6tNCNhqwE430Fid+h0vDDFuLG0J+G760Bxw6LJFhVxNufPt3zRzLfz
ruQgSH+y49MLDKj+UrRS5W+bWwVNIOVkVYcrC3bfzxgyVFCzkEFFTe2Q98os9rmG
DtHOdpJJIy8lYB27VpbG09WmUCiGIHk/oWFg3IXlUtHhSj7VDb+GSVInD6Fu2IWz
CGjobFBkizveKgmv2MY5Hr5CXVp3my29LrqCz/7ImsoRpjbDrkVKsEdWnSRrJ3GG
75crQosNEx5U82ynXVJg54kVOy0cmV/F1vxryqRkDONc45Ur0XZ0XEZfML0kcuqH
HNHaV/h+XR39DUlHjTi+zdsAvOxVa1B5XD2N0mzG5fPtMtBVoGb9z7+yHCs1OvmF
f5/EtyblgKvW7uH71Kj6KjSLgazktQKntG2kMWfD2sW4JkBwQm94s/mz9NM7X4UL
SfoAK6wdr2V9d3FnBa7onAuXkZTW+inHqyS08kv5xp5XXSs1Z2of8tsWSdakkPOR
ITZcIh7jx7TJlQ2F5cE/ovbe0Sqt0nvsQansnwEzgYz9ePmjcpugRYEqymrqLhiI
HlYeGUopyAJNfhfC8BZvXp5Ik4Y15oAllZgtzMJMVOiSsC3dxPXNB53CMWgIrwQY
cTpswCyRdF1g6oUByECB9iCy/P0lkGrgN3m63lEbIAtvd5zNy8m4HnnuIdz/KW0G
kFEhuKlz/ak2HTYzHZXM4P0p9V86UCAaBfv1TmoUr9J87gSVNxu1yqYhqUh7k96U
cMuhVVMrhwY9e74yPUjJWhcTKBYo7GkvHV5G3Ya55ojqdJTCDuQ0lBC7kd3qKoKP
6quSVk8fvH+vwkLpWx0Mg0I1Rr+IBaJc3/xUta5PdpeDp0zUCJSYlPfSjb1XR5TU
IuDCl07JohmnIQzvbyG90JgU2DQjp+uOgqK4poDp0ACocJAoa7YU1jC7g0EFyA7K
rOlJV5BZBK7g/gA9UDoUKSoYcW1UiKZL8pJDfej3jUbshCgJ6Jif76t3NtoRDb2T
QE2DsKnu/IS9MDYiTiy8AenWfYqTv3DYH96vmARelLApJVBbrBkDS8a149p/dfrK
oGTPiMSQrud30a5xusB/7+wJtlzyifb1dz3fv5EMEYL+r3yIa7FGi6VnDPP9bX7z
ZGF4eox1my3KBCLPS0ff7BZkJ8lQAY5XyE/2K5wOBOMQtfnMXg/sGKAeWhRabz0o
pxJSo0hvYLL3heVhHb9cxzQnGwrnLyZbMcqT8dc2TwdNJk448MZs/n1G3tJrvt2a
xqcML4mVSuvnVc7JC7A+/zktckpL5+YFV6vEC4+uncALAp5vequyXmRb6PjPhc5M
CGS/BgLp/WX1jTz/LXA3sp1L398ImTLCT72H8Q1DOFyfkKudry9MM2DqMxRNJR0J
jQ7XuzcVWoC8bOL6iT3TtsFpAr+FFvvgdho4SbxFPH1vtv3xvCLQcmxY83s50bWj
RQM0erYacHmc6rATyG1vlgXeY5Cr/Mvw+06IvqxUV4pAy1S6BTeVILi3JNYR9gH+
WvWtyFFg+hgQeeqKSet83ZvZI3NeKKCdrHaRMPJ+4nvcvHfl/iqrUhgUYvvMV9x3
k+ecZpl5qh7yt+ImbHqB3tdFbs9HrpP6bPF0Rfk1zrvkhh+fVFbN9g3BNcyEaG6v
wB/+wxS4crCMdd+ngKnaypYB6JNB8uBDAy6b+omhA1VWmql8ljsqeOf9T9H6x4HV
NWWQTDD6WZO8XEeVyOi8gZn0adH5Pc/RtH+kRtRFInXgCf84wRlCanYeL8+9vRum
zCwpK2eeAhgIG2JRqd2Wu24SGxn3Vg5IrvebE3P4drI6H+mFlnV2BB/cFzVzcjl1
SbaPMpXbpoUihRdJM2ZBJc8B+rMwU4qC9aprjhZhyxjmAKN8tDSR/Wc33HzyG7nD
/vGjWDybfoeglVRpLfiQZ3szW1vFinynIzqNK/ZCHoK1KnOwJlL6E7brDd6i7Prf
z8nYAXlO6bb4LmgacYE1uO8Y5yxiN71JW3Y9BZWk9bqtSnngmjohDwnQDE9IbeBG
Usvpw0zzWh6kgVsdQlp6Hba6GYWFyP7huGGWDN/zIRJPaSwcSorRk1Lo0zE8goZW
l1+ArVhprVwDS1ndT1FHSKg5llynrxI6AfMGF3CC7DbHGtnf06xXVktrBl9px0Yu
4zVFlFs4DJpsCaS8BJ8h3E8OwBhm76WAf7Q7ONcpBDGuhidhGa/EkSqt+G4bt1mo
aZAFAJmVDdqe78uw+CIeTZ0dbiEgs5oSx84CfKqAKswhzTsuTM6WbZk1Rb9qBwyr
4GA2Y2EU0N8OakMT+Fz1nAMuw2TH/WqGYnlYZZY2M1e5ZDW+a5qsNQMy80Z5X5W5
FgJhSCHLmtxkJqFVrdfJ6FZq5OmRPrgpIseXkOH+jHbhtvkrtQbnYP1LgiEYQLqC
jKaFNnDVa4Q5k2alLbbUPXvbNOvQwIQlTbxOo2kROXSBlJznJ4mV+lnvBkDLqiiC
Li9vr2XPsnRxCfU65FbAxbxlqAo8m8llPIUale9/mFg3T3RX+9OE2siar+kEMb/v
2dBaj1NiqPwrfU2BJ2XifVA3exd2zljFCLYpjlmpkPasn1CCM35n4g9h27RfI0da
vL0foFdUnK18nm8D0jj4H8OqXCzP7N/S1Vp9Q0qTkyVp9vtzH0HCwDPzm/T8tu6H
PE+Ux2m3UWjyFTkVMZhMcNqsDsVsJE7kryfTzGczYYupjzsl1Te/1K0pQOxvMVGa
VbIHnjyA0QDrsDNBUudDevYaGlrz+lRoRRnCt8tq+ceRzKSOOVXd9diKr2Bqbkvn
CdjbKA/VsLYp6KIkNwkAdX54zgQlX92qQOuAovQj0M3QI34y5HL4NOFizh7TNhDQ
EzcVeLhoSvipVrv/U8XBvik6oiQ9g8Eeu8GlloeNVzaB0yak4q4s49smgzwU1Xwb
lwsSh+/HHs9ZenW39UxuWM5f32Ccnu/W9H6MajDdFil9XXIJLQ2dfOcc9IHNLHrR
zLmfZw74I5IphZ7aNMI0zdx6QlGyLpFkTjQNYMh2RQo6bEWeRhCd4plVxM9xYxjO
NA4Hi8c1NyTU74RNj+ZppS/AGsUpQAue22kFwGmYNlLsBT0jDkiR0CiYP4PMQmc5
e/vfjb9bssEBy3V4oI+0Wsmyuum2fojseghz4DCEesaDdEKoh9M1p4GJyHbrmSFn
dDTMVixenXtyoY8O94VMxygd3HtATz60aQJTd2hc3NuNg/Ehf3sUIXBHro8ryAq/
itKX3xe+BHT4p5nxKznIuBZEpOg6u/i71VoSxySytvF0/H1f+qQdISgNj3YKDV5q
AC+qegsmW/iXe7bmHDWtmkQ8WuegMzX8BLAfElcEX0Zs4CYbph72omhr+jeu+Qkq
vGWgzDSJLiiq3hUSgJXBNtILYm1ndCXgXgRhm9HS823Sfu+kyITg6YjBxZXEmUe7
j1xLPa4z8EhlxgG+bgHtirIS+zXPWwZqJa+twH3137BJAmVBAf3hpjVhzBOIjbOD
WHuISZj+q6tQCAnYSfagvL3chx/HMGhGFL4qiUbRmrZWsmsH6qD3Qj333Hw2WNJg
7/J83htKs6WRWwjUfYNH0hVe1B3K+oOtII6KyQtAq3FpeTaGcwdnwUXmQN9BG6+6
6YOiVJ2h5sun9IE/1Tm++C4aFx6ACTgjKuW0/vE8kWm6nKKZ/aJqgjdGeYcjTDL5
NIY8Ob4dQaD6SDvW164W9cDwa1GNBX37P4h5/aHZi7mSZYPsRn6Ay4ce50+7+F/6
ErFTWTsyxy8EKreeWO/N8HtTc8xCHGyHobdCvokVGWOGk5q4y2WibwfY+Xw9lS64
V8bOyIdMibRAaswPK4rWFRCWclgOfXucuY/JWqhGvuLYlb+VRyCvriujGVG5ndUg
O8ANDOe6GoGIiIcjJDvcIadIqfrr9GhrrVxf0yEps4IlJXRYvSFsE2bkHRJJQPj8
v1Q+sbk3Bi5o02TnN0y/cIKBjcrWiOoKyBZa4KDIxWKYbi2cLM2m/QBGT5E3OzLp
xTB6b4pKnF/ifJsr5C10mdMbE+/6jZuoX+VWcMwZqufEarNJaQiBiHtwCK1oriON
o42titEnrgeohEVtB0WjYKpSkEkUohu2R/t7WVoyN+tNCaQks2xVhHw8gIK69Jma
bCSjtZ2kaGEcZt2yIl2J+M46/W/f7zTq4B9o4bw4RIpLfFhCe/IT2kJAY/iLM4PT
Eiks5nmh6IbOoKlOBxbiBr6y7U3qH5kTSp2aVVv29pX/WpYK3J9h3B4P+2G6vHqO
RY5REfo+8oALC22CB4aqy2iz+jb8yYHH8DwrPbsEtGOjOn25CIGQWRuXeR0wdp3b
0tHearywxImFBu0MqsHO8pwAJmFm01XtYEQgEKR18ZbPH9MfYmOiOdGY3Bahf6zl
mlCz5KYm8sy3WrwmpMC2hd3eDwEMycNSeZL4j1GGEJogeaTzu2+hG62SpYLI0jZE
dv5VDhZZElrURioVOkMOvNcgL5mEagMsPlkwbLxw/jwjAoZ7RN8ECuT1PGEw68Oi
xBHmktGRgaZomnB9rQkJ3ZMgu5ONVN3Mm09G7tiTWGjUtsdMN7kGdvFbBnb9JDx7
WO/iT2RmT7yRuYY7iOsvJGBrZ01cAMGu84MLX+HRH1FHcQtDplJhuurp3TeAQiU2
URCK5/Xms6TjaXSeDD1QGkeSuYAgXm2WUzv74gPfYbgP4D3aydaY3hmrd47a2RjT
TkQEIAAnTxNlzGnCP9B5Aukq0avq+Gn/u6OW+zCeNK63JTRG765DqSOKFl40wCLl
k4mxh5+GIGoCddjPFSviHGZCRXHmzwtftiKbP0PhFdDg95ncBLW/GWAmpp/IU2TD
RjAm4uodRa/VEXy2S2HRaImP8FGvx4FBoEUZ972nroZppbzkumv7PQ7b+aDaw/wF
crMjpHLrpBIobKi4QEKGKb1liw5G4I98+wAonbeIbkJecJ8wLQEXHvVWtcgKd5Yo
EOkaAQwM7zbd3xh4hPSWjhCCsC+/IwhIZczUwNKd/mFS1qavNbpOZ7HDq0Vr3s5A
chhne4poIT7HfR4QNFzuKmV/vVEtNkVCly3hpLLYrr8SnxuqmTwujqTk/Mpm7JcN
Ark3H2Rnd+vTWyY+svA6MZlff4XrEwaA3s0VNGgc5KeVWp09Usag9npLHllzF4Du
10lBF4pUSxNt9xGsZv7hiRvrFIfp/fg+l8iomsDK8Xt9JKQDjhgJxfhUnls9CClY
MUlFfFaFZZTTlzedPTUsEvvNa15b+uV0nQIU8M6RWwgXZMpkjgudrN6zC0xRAv+c
9/AkZizWcYe0BFvuqhk5wKphJwtaVfyG1d0Phm8fdb9KVtjpnRVxbmMIZU52FF8d
E7y13qWjtlDCuZszs6/hXwYbqwsP1XC6GtDkUte4VM//+ataI9XGHlZ/enxFBe9R
MSu9yn/3spSdMYp/fm7WhDp4P/Aaunz9bf44lW07GQxO1lhffTJcXQpQaWrdcZ3i
nie8Eu8pYmLt1GfnUJxa+E11IizaUEwW53rO0zXExkE1NcyYTdSfGU02D7s/UEAR
4LNRNDM4eP1mHwf4Z5b9ldJnhsso9wwyELt52i8zBfwyQw4QXnX/ZU+60H8iSyUE
eQtG93ZGfNxa8AdIglClKQ8L0QeMRvDtZXkdlrpd4fyiVCAvALUpxFmSWlR+Dgkh
deH4S2uFLTFh3JiZueVCRC+UduhIZKAgTYwWHzxkNmlIX6zAxOINZxGvsbi3eeA9
e+BGT0I5tA809FxW71Z59JcQckPs6IKNTJUw1zt2mxWx9NKD/t3iEptEhdo2jXB/
LSqMCPG75dHdwWfzRaijwZ2YjQAXBNk3LoeV4ym5ww6yAR3Crlz0NcCuonC1h9x5
9jfP3o1nyjuNWSAvOn4+yYj5wY1hLBX92XP7D6EQ+y54tXy45m3jh3BYA6RWaY1Y
N9EhGKSGRd2rlgInzF+axrk5TGSvnco+esol27TesXZcx0Qrj8619uRxZ//8P7GQ
hdga6hGy7f7Xqc8QtsfBe7BHYXhR40up0t7o/L6ZX1TMXXt4SDfIn5c+LF6dCMe8
y3emW69J57fxh5NtijF279i1IUwQAT6SYV+HVY822Tfots0KWOwmGo4B5Asec8Mw
39jUcvpX3+UGice2/Ybb0cApmk4AReiA90SR2jupLBRzue3F6SkhWH18sBIliwgW
ucbV6rg0UAksrxou67X2GPs7D4+mtEzxrkxRbPMclMRUNZ1Ox2ACUEwuR2lRvTYv
TYooBY2swJ/ggyl4Uvvkv6VfFYcBfXjpqybpWktb3K+d2MbK0HXJvM+YNGWrApFI
8dtQYtI0o+62K8c9pEoVSV9zWY4LSeEW+hY7i4c7zPqhAIGYCVIQu8SKbPeYjDBj
meF3PHZQwDzm0z2nDEfS6VkumhFFJ9S1lk+h2UFJVfMUfcZVtQ7FAcdK0+c6CRf3
QrKtS/K+FLhsVghQ4435uYiNxUSr63GrHJa5lfYaaEoGvZBmmMgglDFvVI6BPz7H
f9klDkyxTasFJ1xQsh2U/Du9NLGUlEmDW/JvceA5g7mfun5V5J1naRtVYh0ecwaA
l2l1vu1LBzcHsEh9YXnlvCzkwWYWP48GJMf2JP8La73KKOe8J3PFXQtZ3TAxIwq0
5eF+1zbawVZK/tFsCpfQc8IW7jmctVxzuroRPBLBEpy1qoubnLhZRTe33yJFelux
pTo39NYahAmHPUA2dMf4Q1PiCAVAF1vkbjEiy/06sPf0OMfhuOR3jZxjEx7cV6aW
n8h7kDRsGFs0W1S3mYeCRvotRTVBLplAcwV7TsC2bFsIOK+u+mBiJqkof8yxkFNo
K5yMmE3vp4FqZChoJqjEgaZnPc4MfVqlbsa/xGoW6jSkrqkFdnvKXP73Gyhe35JU
jc1Wi9SMkm2THlwxfkHIIiCdZXLTn7/FfsZVPN69uMrj8Bij9r8cTwFPV7VuQwA2
v5XaiEgbc6+dkP7Nmx948CCRfyshkz8zd0go1AlB6xJCHLjsQFq+zgfsOZI15l4k
2JKo0hbyRJCOzeN7DCbV7KzCj0c72moFX0G/FpXGWazWTl/TQV6QKCmqecocZkwL
qOApzyjdXBep6FZVzP5wpDmFbpn978akRK9eAc6OVk/k7yqZ77jYRR8Ik4tyKP7f
IshRnl946Erc1hU28MDCb2ZhcDTOWawhSrFYMJAjUwEC1jMtj4Q55drvqONYw/4v
H89C/Bqb0yXmwZh0JA+SbOqlFBdgU2zDDroPpwglrvZBavMAgiRc1+j4yKLyQahZ
6fAL0VaBOydPmnW+iwEJRvXVBgvQxNvqUs7k/WlC+ImqafHrpyLinV4R4xLZ3gGl
ajXZoynNWloXJP469dwtgJiUbvenJG5xIGdPacZ1uobyfRcPjnta8OxqQJHU66Zb
Y9ek7TyVLGDgImwdJqunkFkkM5QG+SvorcLMz55LgYQl0XG1zgwnW5XZtn0qbwJh
Slmij3NyuvVKURD7nDb1rGVENOU/vRCExwDrMOkK0aegQYboqVovmr73K6TxvAbO
KwtXoFyh5lce/SSd7DYMJndN5fHXkEZeVkRZF/8cQzdKWcizEpy5xold4+CpyLnP
3PmH30wj1KXnZpndANm8hc17ZJVJQxnEgPjZjzrGVxs0jN3aKrv1xPgViMyNzTpk
203lAl0PzethFpSgzIZJniY5s5XDmMimapLQURIV5RFdDbH4Ej2X4CHcj0i9PKlM
xyhTHJ8r4GrfNA33cfyO6Yce6yblBAQ02yHljLZCUwf4tRuiwYEwcinjDQFS4jTI
oHemU6binQt2/gr0NhabVfUILx8npjLlBsMdqVYcP+9R5DltOVJAlmSp5pfrrmOq
EVFa1kuBWKezzjlBk0WK0ghEIqVPm6pojxfneP77SH6kHWkBidtYahXXwSkeP6Fw
tlmO9C3p5LXeA+fchvJc/sLmvyCTBdmEYA2/LrLikyDhVz77qsQXp9uBGuNaE4KW
VravBFaJO2xyaR6EviNJ7V/txiQxWfcMB2QPy7nqfH1D470kTqFv+fcZjsAzSGTl
0BGvwizk+SQkP0qpz/wWm+mWd2kdS847zsm+QGuDY0PYQP6BbFF3uFxyT8P5eY8v
lAR033EkNopNv70d06s3ZLJBeBYVkTLvjUIyDYmJJW16XtQmKdDU+bIOOBMIGcEw
U2xfoNb86np9D/fGRWDLX+XuAfZDzUN/86K8CfAQNA2faIxCPH/p5Doo0wAsh/p4
qgXPKtTzgDBFAn8goQO1bDwjqt+/e1xTBvQ0il+rhkMmzEqVmYddN/mrI/Wo85GK
hw8810+Y0NJd/NHg/a/CbjVZogiNTzCxiCtq+ZvgwRj3MF2zQ6wKvFqc2n5I+7Fj
eomGJQlqmv8P1TwGuJyoweZ+ZhnvjeItK08NBDSWmXTHgjKFZ7WXCUWBY0DxBNrJ
UlGRtQjnSij1vCOaZ7qHECZOscWmoEVF51V6qv3En9OsLvl4LcDx6478H8fZYrdG
mT8D2ShK12Li+hX0c6oFe7d84BAynX0jNDIBOR3M+SAi+2TLUPfpv+ch+mRFyYra
ElrR6dGY3f45J8o7IFhl5X+wPe6LtL3oKTZqEh7cXTsRs4PbQ6I/2HoLX21tcdHP
Tkcd3Y+ZXwvCrrhiI5f8o6S1EXWYjRaKuNoXjiE+W/HMKSRM76LgE2FXNKXXVxgc
5tSlw1oto8kMZ7cpi2RjnaLFR1nQtpfQA8DE/qZJtHjGEzVejNtBaLg+DUIPojNF
yJQNRgID6EC478ajCQ8c/vu029kzT7HhXb0bbGgmutR/JT8S7OLmP8A/IKNGWtmJ
PDUcDw6FMBl0IfyW8yhjebZZ9HlF5Ux2iOgoCLg6iVOlL5JMR+PIw4MOrqXlz4WX
QzaxI+zkQV4b1Q8jKhy2lbWvpn83h6xk60iUrchtDRkFdET0Ty7c9mWNrNV3wkcE
/RtAp8whFENiOGf3n5dDG+ZRjEzrvGma/U6ik1vl/0qhY0frShSaVZeausKx95Xl
4rsSbdTOdEJMuhpwIVM1kkMGvjVkhkLRpI7V1GB+aMq9KeTzbgj8EbLk9ff80Ojx
kEXNDmu0zLz9quZ+ylyx2gyLqHdhfatyLx3+JQ13CnDRvM8VTNEWrY5tlEFxHLtc
4m+S40Jel8KhQXIMnWFipO9xSB+KLD5RNtqg3nDnE9EhZE5UsSaKib5oslrjSDtv
tahsaZ89PIHeYa5a5kj+j348GzUFqIiUAz/YwBh5ZxVNuJhozA2gu2sdUlZW6hHz
QOGb01yzvDhVmdbxKPtemCy66+E64X0Ovm28DlTsxOWIZ9rIUB8C9o9ExT5em3Ts
HaJFt32bOiPddlTXLFSlwehiNBNfluml5RxwFcrKOsIfLCqhVIEZxRE98AFwnNO1
Ur3ltdZsq5vgtxPiAok68e1Y163RxBMj+Q0IfiCHcHGidJZyare5RcgH0hRvcHwK
mhTRv2MArEZ2XbMkYA8/Hh7xMMu8IfI9e+q1ikC80vI9zdFLRDHh5bfCoOm/FGGi
bqB+KHkDohhfloBovnGwsB9gq2Dlc2kSGjFDcRLLiKkt25BLnhxRl7OjZID2QRhh
cE7LzLl43T+5/YC8TPoRE0s/Uviyth5FxovnK2G1FQ4hD22Evzwb2JxqEwSo9Pi7
fdsQzRtdl39VUCvIMjSx10zqqW9EvaCteIeEHqs7jefCQTlZYHO11PSECw9b59Uv
l7O1o8+ALF+XpPfWikPGYgGCnZqHPI5JDv4KcHioV95nntWVQvkMQb5wDlFQ7lUe
13+aNp5GKZk0MBatIJtjKfvXBa1FInH7cf/riXS8Xc38VccosYA6O9lyEFvyz1XD
4IijaNwOZLpVBlJrqbtjeARvVrfHJEuKXjFin2F/o+izDmFHv66pPdzUxgO8x68k
KW93dXYZFzYIla7V+kBpBgG2iTTDfsJx3v9njV6HxK9brDmXSrOiT7QaxJUafII0
hD0Z+84p3farHB7q7NU3IZAmX2xDfcKtOggB4pkQV/ZWTR2kloumrbnrFNCd/b9P
KDK+KIxXI8lBIeoSh+sjX5oKmSw3b8J3VvMJJcI8HQyRc7+g6YMbWJSC4aRL8Dvy
VHRMpn0CLaEuif2CGc89WCFi13GFGUBJOUxC+33+ArR+ydqagxY0KPPyQNZsAQ6l
1pEjEga5fdVSZ6TMPiT2swYrv2wKSOh9qbKRBH4ZvZMILGH+4O6J8aH1LQe1jrbl
CooPpqzmHLoG1l4jedWCPZBYJR4bttPDjjnwFRuXZ9vm9U+GyVPsFKi6vecjM8bm
y0aSsuSgtylW3v1/JOnSGa3We5bY4O3TUTJ+NmCS6x4V0j/MQS6B1gKpO98vq409
pdQfW32iCWcDYIr5/jklndObSBS/bsY+rtCaSy8/oVYKYlL7uo/H/aYdQ/o3OtUz
dcV3NdIzkDYYmuCuTEc6ldXv23cugKnxPGt9OPIotxoGkkF6chxKou9RlnMafLhk
ngWKNoRJuqudx97dinh9TmtAQEOnMTG7uE6ieK+w12aErUvMHYe6vPpbSfZOhu27
kIuVeB3J28aJnYvs+oaObB4W9EwZKEDoVEuCqtskpM18bXg6Eap/qH99eXmrvPWz
apK6K2HHxhpMDFg5koZT7nboBGKXBwu5/JuFU0F8Hro8egLtpG2FQYE5oCKPxRTY
4pLc4CKKxT0Q4g6dz6VLB8CUE/1QyUtS/3uHxF/K/Rgc2w+DlXTD/vDAs8MVI4Tt
t3PCsXcbxtRgMiTEFUaxwlNfEHWUze1uDBz6nwEurBY4f5Y+V0aMcuYcQ5i92AaW
ane9iog11/D6mCi8YFQ8WhfGv8tjuY8D7i7ix7+lM/VD5EccZvUGuNpA8U9DsuN+
NAw1WrOWEpK+lFLohQfr9jO9+Y1ce7pontAJpSfJ/QNVzPWBAAaKK6PeyXC9zV7X
ku8JtrMWq0qpbU2et6DPg/7jMxQ6hogyezgQh1kbEK+FG4j2kJIJhpzU07HeaGcd
5EkIckd+PoVfxZ+cZ7EpfEFeL3ORayR1x/yLjm36LxSXp7JgwfJut7BOoJVY5sLH
3qrgcvfukweEUXyf/2ZoKkFsbJOA4yoeKKrhACdSR1zJPTob+Cw/uuj6i+GIUQo+
WxVbbqu09D/cvCkjLJIIqeGcAVjRsDOkK3VZKzkCyWZQWBO9lukrUUuNtMejzzeS
sLwYOSlR89IaC3ImXIOhDfVjLDgViC1IMgK6DR4voCuhzLj/akTwpMuTgGGrGnd0
5XgeUTzp64fO3iO8X4BLtca6FYiGMZnrf5CBp7oaJfIBJWdNRU2Uhm+n3b4f9vQO
9W40NLXeKADnOLTWF/GRz9h/LHRg9DSYSSaGLyoIwzOWrMYeWcRPB+wqh4eiTLHN
DDUNToPXsUXtl5V98OYj/KsNQydmn3xsn6jpqXIoX7ynEL3Gm5LPEJWbaWubxe4U
+yePfTE5s1YZOBKt0PkY/BNEatE+PQ/AZ8VxgscJdanISRWiy+205DUvR77qm7Pb
tK7J3ly+sqWz/LXLucZbMs5jcJviqzj1wAurkWgSCw5RjQj4cUCQhHpveH1ubfRH
gIlMEUvzecjMCHPaRsP/4vPV2suTn6DtvTMXEhUEVHyMWL0tziCBo1XeDSV70I1O
Jpm9HYcvCAFr8zjKojmT2QFgNbRT+V39hvkTDXpZYad7LuOmCrVCFI+QFXQ0AbBZ
+0JJ0PIxSbZ3t+h+t8xzG/3vTskBKycVOVV0xaEa1Yirx6lL8YApLiNtnn9yYOGL
4LwH7645iNwDOdUeSEkGTGyDRZWykpKTOPbRC9hk2b5gc2JuWLgSxkfiYbPX85hv
nrH/PGQtnByci4V120qD5gTkGWM6XwAhYOqCK3f0bMO9s1ki4mtJTcTEOPNB1Sw7
4HaigZ0UaAwhI+LoCEi6B0rDFe5mR8tiZCfwKSRrVukfsCq/rA/YZu939S5RYVWx
N0H1GMr+c6+AiUZpuc6S2VL7/j6FrlpBbngvG7dSmBjGkyu4QVD3esHE8dytL+5Z
Qd0Fq76LQpedk+D1hhkJUf/AZOmA4d7GMbFy8AyKCfNWV+rqFUgC2xsWhrlQ0FKw
AudnFXEOCCkEUublrbAPn1aEdDwFMl2lFzJ+oYjk3YcQPPwrtLkZeqiKqcykC7Jy
S77Vh7Q72KcBrjh0emibxUW7EUmNrU7Ir0AKYOakZRrUCf7IDeC9EuUJK9hiSa5m
WuKZRKk6LurYP5S2JPn7gB8LOV9TmRfMQBrpWx+zTVhtlPSxzbOuJkzyJj8im2RA
SwPZKWJ38fMGOxk99t9Ui1pw5H8BI3zLEUfuT5vjmGMKLgC2wyPdzeuqwJBPOYtq
pbombt1SiR4TbI6iu59gme9N2h2KFVSTvi2JfF+dvQSTQyS9BnRP8WeZQA2j3y4A
YTx9SR6R2LrJj4IfZXZ6piwGQdso+AGhiid7PN9Gis2a2Ha7W8UouYtOMbQCblco
72VFe4cM9nrQwOmKqD800IwcAQZNtXDebBDIw0KBmOZSqykOAKH7pNMTy8Tv1DDC
G+NRObvm1w85+HdKTAUf4yyWnGgzZBXvMUNSReTdGxpSiAARQpG0fB/ffW0imQCp
zl+9eFBIlNDTRHxSHAcvjQ2bIEfmsN2qB//dVtYGhk+UH1pGwKg7CWDb9rCtwoH2
i3UBwtOynspVa9prXCfvEWUH1s40H/toKmQAB5pNVXUP42vosgGSZ+qxWZo8RY97
kYZtAw9R9br414Z+pTSFxir543Kx6gyQd2NGplm+0KN0Nepaq62I1Hk3OPK3WSi9
xeXn476nBpLjVkMfAcjHJlfOz/9sC5TX9Qw+Ydi7HVaudnjC3ZEi7pc9wGk6aQtO
gRJ1VNrmBfEUz2ucPwISGwWNTlNKwfrn/KDESf64ptHsHNlY2teDlaHcaC1ASXPE
0PdD35za4m4Suh+/zTYH1qopnFbdAGwJo3O7c5WpJ/S1oDv0Gfh3Mw1lPw8fAyxm
6mpwkl+1xluW8xkaiknRqCA8tFU5UEiPxsTSDSlQCD5pAaTQOe2eZcEaj8cnL62j
nhC8gpR8/oK1C9eb2945LBU6kIX/vdfyCTzlDqMSysbYkp39smZAVGhlE5wrNWkx
4u9q0azJhlXUHnvqFR950PuMaM2M9PZMeH/MCDgAsJI7XblsevStelm8B04mMH4r
KwppmcMVHmFNAFpbsgEniAgO1uqcNhPab9K76HDbCAJkNpq8dOZpCtcqcS84HFhg
2OEKxlHSQMlUiBhdt3WM1l8fYM5Yt3jicmGLlfYmialKZml8bAuLYvgMPL0xjfRG
7xAjzAMyMxekyecOOoMxI/VerHRVO1j0+DYNrMrAlVtGNJs4EknnPU9gch10d1Fn
TaG9x6vy6Lshk2wIzsn4WjVRTNTMarYC0dx7CPrQcYXl9xIy9NbKuabWeIM+TugI
C1rfFgnDA9YjEyLG31U1dR8UoQyqto/GCs3LBYY1Dqqk1nFTaTbo2bbUBxdV6tNz
peXSzhdfTBPmBfgnsOsngLU/WUbTAw5wfMdqKfUf8oswcVZcpkr2vs/1rSQ5/+aS
DKQKscJVJeWU2IIC5kecDOOBVDTV79Oo/FctjSeBLzwGhwAzYK6VPd/RyAfRhv/B
qd38/ufDckJFdlSvzlyPMQmm198P0zsWzg15rvQHLXfJsPpwcDLhGiJXhZ2wuZSP
/6pO5WbfmVB+Zw3b6OQvZGxVeJPsi2PVOAuYqbUXwJG23L83U3FrwkybGaboMqEk
1WK4H9Qh1mL8M4ThUIgl5AhDy6hyABY3rzSU5RStpiNsxNRUJ09vp/f0zQgSm0CJ
5eBgb/tOlQTg1xOSXrb+c54Z3K9030id8S6XAIP6fn53T59Nh6O2ag60DcZfM12f
9LrK0o/b+q7r/62ONCQuPr6GpQR2xMG+JmaZzy7OZwJkZXDCyGVSxJd7qB6/37wC
2G/CPmpg2CHYpF1APo6X/4kfwSLX/q7KFoe2x8PjlZ88l8J1PQDOrAv3VKkj6GPn
kYEAGtzwtejIIaXHge7odmY1V7fGteScLH1O1nZcefzwDztk6ZAnmraMHpYn+i4N
hh6ceAuoZuO+Foq5dl9Bf29ESl6fDM2/4/4UAIT+QzL845UPDfGFM9i+MO/DTt1S
DfNXlMIN1RhvlSp84U1CFdht8mIoAmtdP9B8CEtkEPuFqAhdND6G8ZzszYO2C5F2
8hehau54vJgVMVuInCY2MZuMMZBAgFAEHOH7LprbcTMycs0xrojfZ+tGYQsCWeCR
RyZQp2B7s+0IroyTyM9ce0Al/Mks1i1vYc1cpsnmYCP6CTIMZ8DTqttZJBd6e3nD
lglMBInQ04hGlUefGD3+xi3q3+b0QOuM6ikWWfhOSIpqUE4yN3nsjtF+rf8lp0yL
NlzaJJsLnvoE8pY9keybGqOOeKkJkt9qloOlnJ7sQ5ct0K2xziTCUhQY8ByC1ZK3
mQbzgy6fsHbt2zkGhDh4I5YPPsi5tCPLV953Ageo7HUZZHdvXH0bpzZkMt1pthkS
oWGuqiuJLSzb5LCtTjxW3nct1soRSN+MwyeiyqwBOLkWKAMP1jd3rZAMU+kM4Pzs
48Kp9iHvcsjiubpqMQU6Pe809WQ9lXZizEz4DwpoNN870CDBThJ20nPATxbd3MJ0
P5dzQQWluXDHVd6jgAqdnjwpMUFx0WjkFgrepKqhgNtVase4rLJuUarRhC8TfCLj
CQtN7KJ39aWjE95vpvrce9LssX7onjquLIs9Xmgt70m+bLzyzdzU9gonzNINEx7M
HiJzKQxrFCxrfiC9skiPW9c/4TeUxzDLoK7x0X5bLUEhUPEYKREdtQiEnbx++G5/
WdvBzMrbZVuYAG6v+wQJAoCLc3wP/U5AX9grbGp4uO20FQewOBYCA/bfHZ3e7SZa
quZLTXQqenlfSyYJ83I5U5yVQJte0drwc6+c0lnfpI7UWobxXWDMKE4x08sYa7wp
JoeESXdAJfiM2MUHESsojj8/ujLewxtYEcNCETF8lXy/vW6pQRrdlwWsVYWfrII1
v8SL74wGituchOyrsdsGo3QCjXsBGXNHT0au/4HJLqKQc5z287bCJKsTi4h6o51h
qS1/ylFprB0OeZLmTZaDrRF/zvwddfVcHRfUO0LHi++2+oiLBfijDVEPPE/VUY9J
oY+FBhlGnjipVqluExHKotUJNqgv3XBQIqAfRnYd21APekcaMRLN7wz3KvIB0aFl
3FtLbIMVxoZ7knfYfdZZQtYDDJRl6nDqfcraEhHyZh9gGupejAv7rdqD4dVvYDWR
iw3krjQ5YimkTC+bqgFWR1J19W5n8fkyvBtxJH4Qod7cJzD4Yk29EjCayvV+U+pc
nlfKHg7Vlp9a9OYMblen6ZAy6cCOZ3XplgRYMFwC/De+wNoxvjkJg1NTwk8r3dgF
uqV4ht+VzPqT2p/dHIvkPwGom9OH9kA0kahqGD89xmpLx9awSEYmqWLLuut+UHA+
xvqWqaE9QQtGTVAIIZivkTWzYadL2ju10acYDkQwGzU/KqgiWs0gIrhf9168SdaM
8MW00emkcqIPNHA8Sv1jQYCqcwYyOWkVh+E6/q3UOkmQxv+lg5cOeY1hWxehlExQ
vYi2rvhd46xlE9o92MhQ4JBU52nd46YpxVkbKFxYO/M+AC4ID0jkwzOVt91YnygI
8UMjAksPs1n2S7QDpppwGiOb0gFyn6C9zUx1ZK9FsXyf3dNpvM9D7IcihxsGAqKN
+SuIQTwOg9nz6wcR2+QEAugF9YuKQFVW16mmeJOqJ/SMzfegwFOO3XEJOD7Y+ByW
BriDUSD63IlfxKxWw2bi4pS0wS1LVGRqWN9cqAoRTyR9uAEbop6odN2rZMUd9RJF
soE7viVLauR7GyHz8OvQIYW7SJ0eXoMvUK+4kNq0AxpdnXOrdi37DtgWye7B+GI+
q/f72d5/+ASK5jqM8Vaza7Q15DtqVuFw5L5wDod0S0JwDHcukcurqZ1bbZz3jUcB
v1R2CscBaL08tHt0B8rIotmRsKCxe2fpqJMHFWbvf/jQK5SqNmiK6KcdqjmZBbq8
Nzdz2goeazAGmylR6IAK1hlHYzYkDYQasizMhiGzCjw2twq3tSjgF/cc3Xw2lRdE
d0OgSs13jbXwXsPvR2Yx/GJ0BRlMXoWh7RfTJVNIsXb6PeD1ndE3iMQDIR1pkTMK
aXwppHQOBCqNoijQawoxaEKHLS6A/F79OBUb5Dto1lMBGCuLBftPRkPTgSvZ3Rtx
SwBk32ZALUqz6uxv+DCVBoXKuPHziW6JDoDiPx2DJe2AK1h5YfG6r84y8DuYU51g
kAWF9IPui2n3MyLou+ywDXyCYAvpoSZvFlCRxL7GeIfHSwnqKWtJ2JvCN7pQxNIh
W5igsSPkqtjzr/BcGOPVOaTOt+uJH+uaOKgYdq10YY8GfuOEeaQJL55tEut2l391
ekuVAyqCOhFcSaeHhi8smN/O4ZC51z9BSv8ATCr+QaUmWSYQVbyRcJxFatrBtB+2
RjHTn252I3ZN/IKRNkDuaW+Wf9RX+s3y9AxzQ5O6ce/j9XCKc4tgO48HNnFnrP+b
Rlkxp9NQfHiCSb4g9awFs2PTetAmt7z53XkU3i4bbwb5W9bkElquyhXNl3sX3xlZ
PGSc1oJtr9pcDPiLhMUjMKGxc7vJZjee2xrFEjT2y96SYO5gO9EpLPqE3cgEqm2Z
Fn6H9GJM6i0XIhJOyuAeKcl+pUouKXBpex+AXTevedWZUGioBRIDzH5JmtMqfI1Q
vv1xOdib0XyQdCQsXTX9DiA2/aPd/0p3Hk8Iw+r0pRorDOz7sIRqYGEbHXItiMaX
E0SA8JKtYw4AUjKCWG6/bXopuo0X5yqmFOn6Q7SgTrONe5rrWSUhys4ClzhBsmtH
mzaupE1Q+x9YXaUuL9kI8rHqfwXiRQ5RwRmtV1hQRC8eUStmWbfHBlZ7nvHXhCkZ
rEAPvcAcHdKJj6ZuBQxWVIFj/kKVmEEY3undHPQBUk4vl3VmfGOG4ZZUcGjYK4tI
nlELIL12oY/Ro/aXOzg+R2XWC2mFl+TS8iCKbK43ch3VyaCeLjnwHgOBa2pxM4dJ
mbd+liScEtWR0KlG2dnPOHBsBQsheJU5SjU81Pmdyz6XcsjSDZwutTMGvwEtDB2v
02ryhPDGulbqxt8xpOiEN2STlJsYjeZxmPrRvG3sj6EbkqTHW5HUvvQOgYjEStKZ
dt2U8xPW+XPXVxHtEtiuCJWxTYW9nGSxIdVPMqB8XOwFraYt0F0PLpRhhDQkQvsf
OgeH1Z78nuGzYPqbpP1V+yQGKXVpJsVtHvBRL3Ii58Ezmhl8bXklcEjYJjWndLdQ
40JGc0sM51EgFlnafZkEPHzhNqRtSZNcuRImJ26cZdSBvcCyAb5rKQTmenqiDlyI
0kCW9RutM5pyIWQsRirWklE5/lQJRHKrGQHrvMwCwMW6AoCoR6yFIFXUQ28Hg9sc
w5XnFSkLEMewI/r8i0hRzigeyhzKKru/TtUDPu0yXkozphCXf/TZ3ZMUCRGVInZF
+S1qLuEc23kPij/xEKTShVQdehyoCoe22Iw57gDXWjxQm+LbK9rpMqpDDEbJCmv1
JXzWjpvIrxtEhEdBTy444rBZB8HHCLRkgz3437wAPZjXSIJ3540Y9sdyHF/nhdd9
szM6htbW2/TnbqwzMZqi3bctd8gtL6fZRCZkzM/YBPmbJKHDCB+KKa2kWghHdyBe
/5LjoHns6APq/PS18STEq1hL50l270ZzBUxn+GdpYhKgSlfLFnHBvA9YhO+r2TZ5
NtZiNlf2pefiTdZFfcb6AjKzWDKzhffUP4ZoVgj1LeG754XWbfdlr6rVmwQQpc3n
UV7/F8vk86BmJGzW/FVprPciMyY50HLFSgI77w+DqnFjQG6dxp+dZ5ZPPRMvowav
smhGcss7EdarbLmLuL9I/GBLn4kYORrP53ONZsnNQEdru0E4bz7ceVZ8X5tX0pk+
KIReFGmaIXCtdZYLk/A5XTQjzqEW+lF1d6fB50PR5vnHio5SeEN+yU/s+tGFktEA
N/ZwD2ZVmzehNSnCm6UQPpZvojDRd34EYi4n2CGwjCmlaHVkAr5H+lO+pl2KryXj
pM/Aj0nQwVDnERflWh7/c60HR7jzkp0gkT/PtqTb766R0Y3Bxx1YZ3G2ViCmFD39
vR55x+Aj8kLzp3zzwHzGI8VgfXE4ZOs32jkBSYEdRUklEe4Hr13xGQU9HC9Lq/vo
kjVADxxPVoh1KxmeWAQEdLCtEmse/mBO+TWwyXGHKheJJGHFJ/F23CmapMBxIm/V
1qehDVWvXBSWoC4uqKG4/GYkRQG2gPdkUzn24sOuwp6jLqbh0HFm7TB58Af3escE
6G7+h8tT3adszQiWl+0+2aL99YpGMxNDonEMVAbAP1cYk5yaijB9RlnfGZ4O3ZMu
o7bIHYZNH2Fg73hLAawVzKsPmslU/RXdCSoUOIEBvy7io232sfaAit7RaXqnsZlK
HlRG03nDE3r46oiIxB//QwoI4wVCa5YXdHR3i2M0/QwGukblGfkcrUWNlXDNjxVn
wxocnO+SM8kFEexzUVjd+e0TPQCjyd5533Y04UXVQ/HRbTC2ya4XBu6nDWJ8YF0k
VBNz3NhCSETvJ/m6Yc1l60oNDNJ8Eevr4CgKnkNzYCuFc16ad/UbgWdsI4B3ovlH
pA4Sa97jA7YOgeNvWHGmUVMPTFZt6PvnY6/BlBCjJetOwqVrBeuN+L8ubZZrK0u6
nUYXdX1uHSuKWhyqJ9KamMeT+tRjf4vV8hpfGzqZ9ny5nmvgLzz/vK1U66wmbneY
M0xHt3hx7bs2WExAPFfOFT3mson21llfSgQ+8aAABQpTRV03YSnSYts9HwBzagwt
cDb/cL0d+0oe6p6qUp5oevlJbwE26YkO5swWJCIItc0gaIE0NcTRT5MVU+A4hW0t
KM5lpc36+piz7pZgF1rmaIAPRK2TKfI3fb6siSGX3lT7mjXp0jlQ7RddKcjv1t5s
sbB738LHETaiRICkqiSRh/Hr2m4KVwxlxv+6S4Jw+V4iCu1jMO5rhaqC1IE5SKeu
UhlLko6h5QzuCQa/lkJGMaDD5RqnJzJrH9n+VbmXZpn9cSrtbTimh2WDjx+w/ERI
tfogmDHwoVixoiGdo3FQ8r9/WFqAhH1fIWwMjDRGViyvrkiPxVzviHE8jRohpGVa
hIs3PYI3e0CQ5CTVlvhMhTByVJA+YEIVJGSvp+aC4vXmmVhKWM1pvkicpHgQ8FAc
RyeB2j049DniYW97n3VH7m+tnXvuvZoWo9rO44RPWd3nFB4A7+3dSNJmQZfMfpP6
ynGT3TbidjSQ9eaEVkLwRXF2DiO1FgOKBBWJkJ8gBtaGfY2xL0T1lkp+ix3CttN4
Q/bPXgkjfXUibJOIJdzn7UdrVmnB2IhaFh1d8prF86/ESerxLSRk1as1GVXFeKm4
o/CZV/pEo7q9MkOPteqMCWRkrlMGjzVNzlzTIL6TVWTIVsZquT7zRycYI3C53vju
TVmKokzi1fSWxJpmPGSysmlY+AM7kmuKXAv3lubF+aiei99GJ5E5uK5+4ucfmPCi
nx0WUjDLcf2Cmd04adMmLtvKACbQaRdUQnUL9tNrULMnuHIsfdPlzWo7T0HueEps
YZfdQQoPCWYhPa4sRThMki8EbtpBRKUIKR9rQYsISeDwn+h1E7QHda7x2YfrGufk
w0oFY5VdAexlicBWhTq81eKPx2wib1gB5/WJVdD0j3aF3VhHwErSTP7YIHTJJBd1
6p8HkCjjZoPy7OLvA+2+ZHt/q+L/LHdLhvf2jg0ndLPnEdPjcdZg+7NcWip7s+he
4fMbb1fYfMYFRVbInSXAvcq8E8/jKev5/SGmVOLyewGvO/lLtJ/uFVlXnEtQI3Gn
tXUJQk/tVLwjmT2s4tbm+9qogWtKt3tx0Q1itWaqU0pmRTeZgJILSIh74zaIqShg
bG3TOPUlbA55NnZ5Bd2dJ2gKqwaqH/efM5RCZdP8rXlBTogfb3HoMCCD1Kht0DqO
bkD5LtLyQb8fn/Xt9PIJORXMijwXVeml5uQnbUGN3r1b6r/pRqHxkpnm0Y9pqmTC
fGvGY2gu4u7bGZHMgUVq24jbhlwk2N/eukxAmfiU2o2QmoOVFqXChii1h8Nbrcex
2IiBIrBvRAZ7zdtnz+9r0TY184SSJAgXkydJQe4aP2MwEaOGNv9WqKVxzG8ANoRc
xo+wxO39aBgOcgTI1+0Ye0cpRpkiWl+ufuNeNUibgQRtnXE9mSuVSMQaTJinUpW1
ABiIcdVoO3qKkm4cuvq3j2CvlnxbQOohOFa5kPjO0ibAmrqqlXJ4dJBN7kMSZorc
aedZZ5zuQ9RbhvevaBg7sTCt1vrjnMTZd5XvfpmcbjhBxuTgXZCuKOtx6VVupl36
IsBVsu10D4Lv3B9H45Zh9gMi8QXrz6t3Hwr0lCCIVjMbVQIdieJkRAneXfYYs3CW
INqCQJkSE8Lx+I+LmQJ58U0rAmspM0P6Wmjzx5o0nIReGf2r3eZnGF5/PBHCE4xm
uyhY6uxSTr7V62MPxGiO+zYlSetikmSRkNY9K25ZogiVvMP7b6BjCb31VpTyaGvL
xrt0kENZfQ01LAYtNsWJ2Dng743t3JWn+m4+z74Bs+A/QCxM+j0W8qW2v9iQxkVY
9HOi/tSUO1kC+NT8o6WZwArnOhRIvoPrIQLG1TFwlBG2QeW0Fsiw9yCYv2IW77gA
qyI60+brvY6lJwgWmUUqByPQlQlKfE0eYs5nNDBZZNhIpZhTKucaQjVihDhry7CF
fPX+izp46OjvS62SvMqpzbdMTmIRwq5a9yMaxPHeA/72NcEU9o1pCmMnDaSptSXZ
EDZJCRO087MHZ8Q7TlhPXLZmQRB6JDATlcYj8+AI3VQ7zWWYN6Gt2t2EGPRxI8/D
xTbiFJwJIZr5rkQ7/f+UMkqaT60UUw70ua3C97hp/CsVKA+tHN5dpKeIqHYfqFxa
C9ZfoBwHbovMs0rFJnoLJhTWA8AuiPDYgF44BiSZYGNs2PTXoM1NCQjYGDr1d18A
LYVbu52SPI6nQ5Llk0ZuPf4aeoS4bIhs5AMCI+Po+D07ApFY80w8ntqFYX/Qe6Se
CZIKU5+Na+poMKHdrhoIgCL2j5g5P9Dz1sl3ReMVTl+hP+I+oiwiYKre+1UkRuYN
C+7vb9GaPCZiCh0pOTnhPneP8UjFBszuo6K+M0Cf9I7yc7f8/v/LniX7ZSExKgbq
a8iJTP7pddqwRRy9MZw+Z53WqmOZXWjXCXbytD/pBzSCW2/y4vyoOiCXSSdlhvS+
tPUaYmDdwXtqEHVo96uMnjlxSCgjdthzRDgRqzxUQ2vpHWjhXkJuIncRYJX35p0E
ZzCgL4lvCcZleiZ9ksUVFStLixGf8XJdf+zRavKTlZf0HV9m5XQvGWyJCssAIshS
kPmM+lNDhuSJ8ws2WDTPa22g1gNjD+IRlvpVg9qf9BIDx8lGVAIsTtkWJp9MJdZt
lVngbQGzP7vfvouUQqHMrGwXX0OQnhzgrvPXvqircO3Edv7drsR8jRjIhM67lZIF
jHkShLC52H3S6kKKCyPNajQ05n/nKGIYCTYrIFkH620eOG/MIDlUOd4O1J8AhOpV
QuIQI7Q+iTGX9xRIwznDl9M5qhDEkX1n+ESJZC/+R9ySH6V4bDXtIZuY5S0tYWdG
PzlXcgRTgPWowjLixt40LTgBhExCKfe0Aum7vryk6HCjlHLSUVfHvke1fNSMlQ9P
I4X+0U3mR839CxmMC28hZE/6voVuHFdrqgU+a8zpaLq51dWOwSF33MyExPAy1ELs
o0aJ2lgVD6kLOBHgtQggcpMRBRpahYjEsbKVVcXjmXg6A/LsLqQyT+mEa+6VHyf6
lNJ1NFq7zUX43S+ZWqZ4fZP0lGItN+Diyi+4tsbeWLf4KyvrCHzVQSQFDo4uMB5g
5oSgkS0l4X1mWloHv0bAEM/X9aTruPIJQabgq7ToA0Qk3vo5rMhDh57vQZujOzjZ
7ttA4W3T9L2VkgTVwYcyWHsqQ7vn2hRBSsOBXvvA/MoCFMRhR5O2BDLrv4hODXJV
EMXzJ1MDzhAiX6XlTyUNe1HEponQSa/c1JombvafOFAcBz1moxmtrZdrlqR3jrPb
zWEj/QQRN9hggZ6yqHhLO+KnysurJBgL4v0Iom2ZlsF5XlnddYdnxP8conIwcl4Y
e63ku6WF8NOxWjWXfvpf9wRf+Z2cyG8TItMLnGLkn3c+8taicBzN8596mL2uOM9j
sytzLhxuonO6g3ZXpDulbBtmIgtEPV5LFRTGDoqSN3L6Q0zRkdN1D4cTNnakijkg
Pd1+pMxKsbq06mvCmG8Ru/I6ocge/ofbgs14UoQOoLBV8mfyY/KrBCMKVIThsn5z
zjxOKHJjwg7+/tzl99ZkOu0B69ZTM/UFPrUGocF6bAss58UyN5g4b2d9WfK9gp7K
vjfxhUdDBAEm6vgYY0KWFlY8OeV6VU6Kd8nkoGnu+CqeOqPuCIf5Okt8RFNbM5Et
k5gz3SA1pTHPf7a0dCShmhoMZZi7ATyrvbWZ6DcyFqdwd3HTuiYPpJW34c/TlEYs
bjWJQZK9qxUrG1+Ae+E4PU2Trjzu7kFlnZ5kBV0l7moYqR0SogOxBoBTvGfa/xII
hWkNseFbz/nSZM/BD4yNBaxIhP4uR4LuQjUzZTEJGVAZtBSfUVxMYkfDq8Jup6Gw
Q8/UZkHkzRtLriAqWJIAvZEiJ2fDe90Tor22DEfrJvr/PPyLPZ0jexvh55H1r6sq
srQ4dmKM+daQR5pjO3VYV000xHoGmxfKJRSzoq45Ds8RJbRlbldmye8AywsrmBs3
Ka8hdlAM5OqPTLQ/C2J9G9WDGqP02KdidGzU1rNZm1n+6F80eRjinHKvIy1SUHC/
QDAWaCdIq2e6eNiv116WABz8HFkmS7bSY8R9b5d9U+fBTAHM3661vsxBMk4T/VOv
5iQ10MoMfco6V3++PMXfbOM3SRV+qQ/ixgsZLhkT6xAs9V8pST6oNScjrluXFvkN
DUa2ytbZCi8Tgzkk7is+nrPvZQHWBnqdzWIlGlLLTh7Qlkb+Nxp6nXCRmSwbG45a
vN2zoqFFYOJtyQbpMtY6iSP5pfwoK9P57aLBlYfP8/4X2QH0To2Ti+giClzRyUlu
vuoNHmRtsccCimOlLMhR5+Erjvnv8Pyhzyi4iumqWuxJY4DQXwJhewptF3FFyvXU
5Xee18nylqnm/40McZXbO+06eXZsJCkjtq0qiNhandG+W5jeF+80riugvKFvMdFl
Ual3PEfrhyzqAdipuEmKmJMAeHIBPKRss6xXAV0AlGaeOc52DErRrqWr1j6+pKG6
qD36n23gAL2dahSz1oS/yrH90WFnnuJ8p+W2Wxd5I1M57DzHV5v+V5G8CMLIjK3P
SQrQxRzMiUpGTLOOZ1iKbkANUf/0iFs3E6qFbkKPJC7FzaK2vljfkOhpSuKMXr5U
08KGW73bCq1GUprWpVRfKiOdekL1fxAgt7zbwRTmeufzR0DiFdO0Wqi8jwkcV8p3
LkqeAh+sxwh/Lfoj2iZke+YfhDDvhfPfbVPxoDNT7p6QmN/tGXsGwWxckMruYSZ6
1U+rvGpFVtDHEtKMVl5KP9iQqQPQhZv7uVHnLCQCIxXvLO2p6CXJK6KoJXxH1RTh
Z3kvfZq7IWhlQYEUGJZucTWDnHx706DogREwgFYDZ0aura+UUIA62JJhMQFwJgdb
ps1HxtAnfMUwJgj4xN0lHnUdDkNH+PBi93PcypAS/1MwrE8DVPJONkjptYAojs+/
UgwxhKRi4x1jbtL1xa8b/OoXdwLX5giPZmxKcX0FSmJoIDRCJL6ubnNxMuNF+aHd
Zx3dsZG0BR5QptTNxM6rXdkztJjI5AobFcFvWOxtGlRiYH5dZPDrP4OV+Th7flAW
os0MYuBAO98tyiXsRtI5UK2EXeeXhpxxx71TWEWBAW0dYKYOpKG+hA6CTfd3KFnW
SaTXcC4u1H5T949u1injtMywiQjjW4dFcNugbA5Qsbfsg8tNcmBVju4nhv5NSZ3s
bzprLyfzcKeiIeo/BwBuKZtlzAcEBwpEJwpUyCkMKDq7fbUpCEnKHMpB8yIsD8AR
xRhmvu6XBfnuXznjjJC9ZFqb5PdNDK7/gpSh/rsblCQsDV1NPCW1yu7KPhVgCPD/
6rQWo8viBuENe26FdzTo0dj8xSkFqDKaxqagkTp1xl0m/r2CsMi7psuqv6vtk3Ci
ImEqzb65W/6Ngaiwjhm+qBzLSqsviYqQ1t4Tla8TWu9r8SXl+Bbe7LO6AmqdNP54
23f+kwP77pKSO7y44LuTzWkzx77KqDSIWGIup5q2j6uuJbi5BP+eDZ19FgrAhtLs
yu1DdrksgiEjnA21rGKKNV/EQclEoBskFYgegMCWT8m9nIgB2uKR7H55MYtM01y4
OGNZudYJ9V+VdufcU4q1vujqb9SUOR1KfAwIHr+eDiDlXCSRl7YplrJAl6nN2/On
jdQezAdq6D3z3MTtWFC8oiYh9GgDzYuYCH4dPuuhQ+ZZ89t0b+Rga2qzm+DW0/F5
mLLQDmdQhKXE3nkB+2ZXGMoWsijopfcQ0YP409ck5HeNz+3Eakwfk4KUOI43qW6z
U/ZX564sHAFGtJ0dGjMoxbwpg40pTltoVQkw5bDldgf0287Xf4PHAnlUnAqFuPuN
/q2rdQPACnJS+6ZWNOxAq29OIrb9GUW2Uji9z3NKKQH9oWhyhRhpfvEJ8eDrV7d/
UXqxBRimTPxtanonJgXNdb/8oYmfS5rjJjshRD527KmIV++4yTad97pAClwBwA3I
iEo8eWu4FZWCFhb/OC6mOA8qsoUd1PP0RLqwZH/GmsUd+XwcsNspHdD17jJU4Tcg
5re4h87GFpMuanFXXn/POQiRFqwRf3TYpgu/SgHhi1YBLwRnJAPu61a3B9Sj5JnM
5h4nbMfOZaFrGW+IFWT2kHcO3piLO8iM4cAUUcrvvHbfB1oXsoQKMMaKlp686KBa
5pSaUCqRzfCstFEgaWhcutxoRvlh9L6PNDUUaAyiMxk6bJ41FFnOjmInK10W3aVA
QhwNJCTSoO/sDJH18o9N/f/cboGBlU7eOMURYxFMY8vRDEdu6VKctTpGXZMn/EcR
yfC6NpMR8fYHb30A2HCqvLQ5uNn7Zb7uBaGNtgdjAopb+PEfFg4UMbdKJ6Vqs0v8
HbvfnwzxPy7vkEVDgBx5ESh8FaWEwVFs7i8PFU8XWeFwCI97pbGYP8L4iqqat8ND
VWl4wo+8lQ35TVRk0Pp/XROiNAXkfwErP+WzG/9Vq79dLO1KEh/lww5AgjG4wD9X
WuZBU+xJK/aQ02/mSutQFP5XE94KkNY/oZ/CYPCpvgy1jSEjlatLxjggAYL6f1ds
kd8pzW5ainZTnmITxw8C3RW+dEGfTo2SzvmkAjXIYd/0dbqd1UI7VSMF5J8uXn5/
QAV7D+1eGWCHkUZ7qU7hWbxdvAvEmtREbu8nK6HLIWYjc6aPVOIJfN+OwP+2VJo+
2O6gVWSve6jkAXOA/TUalU8deVH+cB4WN0NQ9arbqhx+p5Y/3Jn67ZAwUHQZKX9W
6qbWJHI3owSmdNrSVpECFywmkqicQHWgYxi1X1jjZvAUa8mFnKdfGuR+A/TsX169
jUQsKMDJtWdbs9KFm8Uyq9OfMOBAU8sTFDgtYKbfLEXszjk9joSCNkdwy10W2XqS
AauVCBSiGPxyfFtDtKxiOTkYQ23g4iw862O0/tFgQbAPxc9Aug2O4RPp9hg7vUni
rsmJMiVCDvzBDsUzr9LwSrlt/9dmunI71iQkNV310aMWWYLKO5omiam8p4StANRq
qiz7lZmM0tgzI9DQ3sk9MW+Gsl9HI5deP6IBxjffw+rEmMdkWOUW00E/Yf1E5Zcv
mZp6j6DreXrwI9u0rezK2GlpYrWHtiSHJoRfgngNzvvOGTaZoMbjUMphHGOpjNbW
WR4lmSmBITWw1JPfh1K7cJHnp6x7COvP6WTJyARS57K9lx6Nl2EzSM5E5nqyPlwd
aC3DE9YY4OAf/LXLm6ecjXxZRASk3QdH1Ak8bbEzsneioGKHZnSPEuzhmFTEN8us
vS44k43rXLZ4Dd2HuE81E1gwUAf/y9gOh0usP5RxrVzNaNGd+AFuCdLt0VbIJE8C
apaEIiTxpjjCI/eT0KrrdRx+12/3xgWUsvF20nO5NI1hvd+XlKcNV/Ok3tSOPzBh
ZyEUnYF4Rn/kb396JWX9j/H6iIxSh4es65FOkUwdx5+UDlwvptxFw+p+yh9GCx3l
nnsyu+bOopzAMhAoItLF2rwOPzFaX/IfrBrc+qtgBEfKShdoHZnPT75f6/oAFeem
oCSlPGiXdUQAxhCWcnG3Wr1rXvqNjpZRXDZshk9J0ruqPFOGCyY47jWPbADa4kqr
p5OlNEvCLD3cCkBqP1Z4QUjKrc9OVqdYNPsxevHLzs9pedP61pr26MQ/jkHxpZ4Q
Xr/cejfzfpqs7EceCV1TTUckJR3GbcCpBijL1YykasePADWNdd79E9mKMmCVFjHk
so5h2SpIxdU2S2VWzSCqMXU96I8tY7uxEkAk+R+z9TeIOUa9qaB7DsJ3GVsyv3ib
18qstgH4CJoweo7QNBdeHOaxJrBv7lGucLHzFDhjmWSlcLwgGD/kXrdYW5LcW4l2
DM9C0eG2pMGBzZM8K/PlPB/vzc973pY7cwCQ7ht32XYxUYe6JoyVpi4COe0jzUQ4
ZkSqAm8dKZ4IDMsTH5kbWTZC3yCQHSSr4kMWh8y/dSNDRx3MB42/PcMtmKOvcXF7
KwVYZRTS2lk1RnMN81g7roHy63h+tf34Sfht7pP5Amd2CL9dAxvt4IqtxMnd/OUz
hG2RjfCKceA65A41pfzLc0bbPx4cIrevbb0CE1mtxsehtdeweKLG41ums4piS9rJ
s7wT8pQHQ8WPQAjJeX7wnxDQ6TitTohoEVbiEW+4BfnycMqRZwZlmQcZmtj0anms
SBbw/E75zSnKARY9TZ37hiFn4gZtRPRDIWP6DQuXfSebBHI2Ic4zIm1WnjbRn3Fv
QUHFbz+Iux27Rz1abey9jsahJlY9U3rlEJqAnoEu2MXpHD3dhz3FofhSmB8+GqTz
1NFnFgFuQ7C3aYH9W8vTvBPWqxaiotfLe2hdIz+pP/j+OCa7kHE2TO2ANLdKQhlE
sG4pxLB2aIeEuJF/bzTDr9/uAAweEzUD2PaH4Xl8KMI7KpJRyHjDd8tLNVdC+aJk
DKJweYCIIJKpVp6RqUH06ePCtoonZ5DZUzHzm1CtdChMFTacKLMUgkWBeoi1FyjY
GdpI2eK2IRot94QFX1yfthCNWerbNtgn91FK5Hr1Z/cYLCCqVUhz45EPW1Z3kF/A
kwkUuPsXxCzqayCe0Y0aw57cLrSBA63bko4jRSFT++6Q2Cvy/H9RowdDd/IAfE5X
v+2OGXj7fZ7IUFUZEYk/XIXXVtAemfTmX5zZhs3FQBwRjp9B0qYWUzT/jZ6dlFMu
58dzACkeo+1k3msUvUZLwpJAUGfhrvjpIJBVr7/xm3RBZh/qT+1Grjlw0aDda/YO
VJlTPA4jzFnAHgrYvvUvM++qdNnUl/zAvRF4uoeAJ9HADzWE2W+W5dAhw7OYGyGg
y8zebgXMX9lKKDl8zAxu1S/0TbFPjOgJ15GSbkLkH47LngEesFyGKP462GBpXpGP
UO3CG4m2LkQwxXR+BHwD5AHVnK7s6O6vi82lU4La4wvmBxfjpoqdILpL8r5vvxgy
3AWzJQ7LlGXdERaxRk2NBlvaQuHtMg0NZc5Y+bQWplgVlgXbZJdl82l4H8+3zppR
06C82bhv5+b5KH1dh50mJJzXV7zR2aHWg2oSjhLSSiXqLqycv2eSnzxRQzTThSgj
vM8GXUJz6kWUpCyVCns74S/TfFy4yvYtDHlG4M0BH8QbzjYsIdva8rrFcXIwmiJc
kabh8UaTGSlkzQz5LtW1b6pk3bL2cb6AziVfvOAANB8SlzhVIkFUsAQJqrdLXYts
kvXR6znk7OD5ppT6uRjIVx4752nOCFAQLLWdUdEFYSq4fsmxYJZQoFvyzKbFx0pw
bgVsVCMFANshmVLOG/TFhZfYOBlOxHoyr4PHnqX+uC4Z0iiILiKCPfeH2bFhXwCf
elIrMiJqIRvjkck8Sic8FiHzs/FeMcTZfjvWenPaDw1/vOQEOPC3zdcSIOX8/Dmx
phzci+pU0oXWViyelYdVwwwup1GgKf7RTzIVeYUhVsv5/PC8j91MHKFpsL2O/mW1
VZLbYr+nP1KseZ6HLwBkTFTSpJ/hKcMEyDZ+OnmzB8ARKoRLuFF2qyc2DIpFoKSd
o34hz4z2JO6HGogv68Hpc3ZTogBosJDIXpI+pjSNcRzvm1ANTgm2GETPzHIQ9s2H
ezxxEdFINc8YAquzQglscNDXVP0zqx8+pwcffT6cpb/oJWTJhuqhL7HuliqdY9u3
fAgz4NetwoJwlD9F96Ny6F5Z3hDggFfxvzQ/I+/S2B1SgF65bd6sh+EUWHPRjyMl
c/ny7sCKJud5l9fDqItlH5YMEo3LrMgWRKXlC600Nku+yvoOD7Fk8rWdowpYZ4MJ
xtSonVQam/OozZHQBlbIUJQ4XHs/2pfs6zEfIIh4xBxG58OlOVfSbnV3Vd9TqvGz
kDYJGEEn7CvATjc/tVm+mRzvdHY3neaF/jqjAgJk1ngIGlFAFC0d67L9rdM0OD1w
94hczBV3AOxGY2IKDLgMemddoW5hiOl3yHed4smzw0jePpH17Atqwov1xbUqNm20
HJccgUhavBPebBmfzh3nKGZkthJGrLcolGaMb67Xrp5gYzlYaqQitpRkIIhjPfNt
yxcUByF3WBTihIm+9c393lDe6dqF+byP7/7jQ7PL0rMYBSlts0hnqiX//1W8v21x
iTT/c5kEmKMRE3rYzFsWXZhj6GaZekcMA0YdKunhOmAPkJZsKMAQqikAZu0mloYh
08MlAahKbVgmUrNLB33LcbWxhlC+bayOxDvuI9hW4DQQJH4nxW2csgwQ6Vj8F8ty
5mSEqryBQz6BD3V8IVfiJv8UudmS5HOYv4CkWx1+otGVuDaKvllaSChxHKZFBiey
AP5x8+kZFAQc6QgRY77bEJlBnXXDgHhC9so5rlkhE95yPMoZO0ynpxwdPWFqoL7o
F2mXA5o2YkkRrN90C5xXMFZzdztmcgyaYg8Yrj1OQfOeXAPu/WJrI9eQDSoa4h/A
XHeKXiIEUJfNhpluVHUhwecBURT9fzE6a63t0mb+vndnUaMKNcDrY2NNw4X+GixT
0Dgh1CPeGn3+JkjCT/uHEM8E/yEiF085NwYIIfO2PVTMWhwST0cxe7OgH48SOCGO
ioY6kAFYyQ4KrefAuK5svRNpn/hoo/fEyoAYWiRVwXyB3JMvPIcp+ucpfX5r4jk1
JTagzN7bJ7BI9WV+xnzpjZgieHsCAkvVnQHpPjiZB/dAhuXpXw8rd9im3fOLeKbe
VFMXCeN7sTjAjER1bpTOjpsXHvhGIK6mxeP8HaiG8JbcSr2h6PHegy/tV0QvOLRm
X6w5GJJgD/V/lsUMvJ0XfUrEgO8Zkyrdigv5ZsCm/dftzeJ79vGlCwVWUvPChELt
BpPgAB/IQRInm06klcBUP1YQFGR6rCI/XwF2ZUljVTp6cNAbSG/doQCLM0DjQLW0
k2aEKhi8bUZjNzx7ETrwdDcjl3yrU05HUOtNzhLHyrs2lQdqa4d0WqvmE4uEFguR
i2++48VmlB33MxTgVmJLrOHLwKwt1G4QAriJ//6YIsysz8du5Sbqi20MfgzmBami
SBGJav+FhESeoEEYE7ESGL8WlBUABIayjG3FBn+I7MTMIzy7jWUfMCwReBWR72qn
POSHnymqyh/jaXOIBkHkLY23yYqzPyGEWVM40Ih0oFH1CUlim55NV76ogRXYLpvK
p12qgWNJTAI7KtLhHDwl6flZmMVOj7FTzhFtElFJMtqkreMgLr+Qwo3ktJypF+52
grtShinYR+FYD8R3VhKrEK3TuMpB7BKnIsBaSs5KBILWzj09fF2Qk5qk/Q4D9yn8
97g11McmKYrXDOiUP+PRAPI46pmohOvFZ6E+1JNzH57pLYU2K5KZYAhD4RQEmI9w
F7667Z1gEd+9cKjb4FsE/47641/mg4FVL+J4vKris7ByHlMqT90VMhVCZVzgK/N8
M1DUaKkzvagfi/Rd1wVyZAMzB9kLRJVs6yz79/7wMNUjeil+TacQPGsA2DcKuUyS
vER6Y2aJBvDI+zZf9yKjT6Bc5irdJo9CJMsRgc8hi6fLalVLHOWacy1Ly72ZEzEA
f9Ks5rLfCnwqIEc3L4Qu1kfut0KL2ERufGLetCfdJGWxaISs++BiWiVrzOOCYlEr
SO6xq8bAjwZ19RbAHSR1qWQ5ymUZ9QoDuM9FJBrM/2BPl3kyuLnKqRen4v2rdtev
LV4ocYX82/ObskOGgEeljs+Lwug9f7bWHP5/V5/etA5s6UjMDh7c5gcIpA288MZB
v8x8NJhK+ihJxPY7DTCbrAUcTwIuK/K5bY9odVEZNDb5QVgD9GISVRd4mW1W5mua
ERhmnNWiEUpxyYFEalwnSvbAtITkcVZNOOt40UR/hrdfcodm/pSkTaJkZHJNGylw
77dCVM6H6I41ieLBdOXgxPorfeqMhDY2DI25l5BrL4LWjI3Os3tC05WdjW+AFEpQ
xbTGKQq5oFNBCqE6DyjQ4SPx3G/By8hfeHBHJK9fwdDykXyWbxVgCt1lpYTBNGfk
DMOHJHovTEepNEsVqXocEVbkFeSU/FgV5D/7c4TT5qMlpbabcC+PJFgLjzTgqdCZ
/JuoszbZmJRNh/tovQcjutLGrSnMfSGKQKGFBvdWaofvj3fKkUXPYzJTfx0pYFFH
+rUvjJzlHe5pae05X+TAq/uJYYucFSObhxWvW/19lIhc+irUw3dcsbKsbOmvCQoL
mdT4cu5fDp9wGw06zHTbJtf4Jmcx3gWuRsF8+6VA/UOScziTYhZAcIHGyV8606C3
y4tr5KRpij8r1qLRjbMTJQcHf+YOmUnTT5Bq/xHIJfy2afRdhbAGR2R5RJ6lM0tx
xhoCfPcVDp44nTJP8qsVMKqvetIdku7sCryWRtHMw20J+AeWOWW59hngji0Wf7Xp
ixvY8o+wMIkOzxAYU/OzDkUMnYg6BVtdKSRvPFtm5lHJRWxSVxjc0H/GtI6XHv2o
HNFXqzyE5YPGJN8jygS/0v1febvxifdCyB7zzHjb/ETnceYc0xFy1Uma1fTw5lGS
cx7oLAZuopaef2iLphC3dz60YILb4Fi/Vcy4yM9ebuGoBFZWe/Y7amyqSTvq/gsK
JjbwEANQd8pPE2g3b4l3lw8qqKQw+ljZgjUvXQz8dViDH7BIHlXemr4jjPv78CyZ
IWcsG21KSzl324UnGCeVhpeN8mRCdD718I5Q+rKEtycXZNwO7At8+9usenTKvQ76
sTnFQoFd2xke3DR76lFSs6S6jlqYpPma2ahpQTh78559BXDxAuKXOajmqTmLAjbj
Yv3D1sxEhk3653FMSK9xy7YFuQwFwIrfV985pjlzhN6rFYNhZICoyuWLswTHmoua
GHb0dm93k25luaSKTT/O8vQCXPO2DT6mTF2BEy6IEFJV/7KW7snXXed/3ir2MeWR
d8l9EpDbchUpFUzzmxxQqJR/1/bhkMkrThDR31OeRKwafFek3/1MWK/Et9JYiyr6
8n/qFEBO88mUi76UT8hEiYveB/79N8tI3FnMYcs+MT2d2coTeuLZ+d3RLKIgdY1b
UYX5UCZ0H+HPFuz//EewJVgrltt5QTuH47DH0oXFZ1yWqXL+IA05+iE++1tcWVB6
T6lxa/ORqDUZs4AihmBEL9a9z1UEdkPDJebT6Fag1w3glLl6bjP0ztwfdSSPCgK0
LLinvwhPFo86NUT5iS+GDh/Am3UFTyaqqhvjbYEc4p990jJoNU33Qu7aTokPPXC6
qjKwBu61/yeJEh/9CdcySwYwfRFpcCoJ7I+TAeVcRYhtBYOx6tbe28KpkPzSjjGR
9WCar7cyOYTkMcSBtUFan12NhDkNXeeWW/CXBDODLrtC69wM30TCsGmBBC4owpqW
TlEleudthxcDskf0g0gGnkHAQhq+jn5Dw/1mOJ5dxFBQsk465ELkDqW8GpqEdwAv
3WnVv3+bgmzXwQWbJgv/iHT38KYQFPw0mlpyuj7t99x1omv2BDU1qeOw2wKvYDTg
lVaK3rmHTMW7HeVxyfXprPvPIPvwcYrXdmOE7nh+MHivtnjlADUtVeOhmkyeX/OA
NMusZyczIiidSiy+hCiomYFP9MYuosekDrZYxVMdU5L4vKiuK6TRyJJh/39jW6gS
WwlDs8581JA8y43pVB6K53FYKZn765LTg4igXJBhx0WT+nOQL/79kHZtV/x5CH8T
NbRLO9wgY9nMwdGueVGGC9wrMwnBU4R3cf+wqZO3ierwRcV0o7Xqr729LJrrdr/R
z+8Jm+fWOAw/yRuXfA7pz9/52gQTu4GvApIwb7LXVgGJzX7WR3nUo9Psew1bFaNx
qUARK4nDFD96axXl84tNttlWRJwqMuBFdGMW3wd68zuG+gdpmR6jQNgUaEZWaghX
pDZ1Rf3dHppE1I56OUZvG6eBwEDTFic7LDTyKgC7gsL1esI2hkN/iM9hAL/9HTH5
F6OQBbFPE09OdI1LcMehnjxYjmKLixeCTmobQPgZyDYoNaIDSSlF9N70f/LkcYHc
4s4PR0sNmwGfgIlZkGdtH+RHY5m4XwusxHcfnmdQTvEcUK9CtfgmaYZFxEanwosQ
p6yGLpCGeiNm+gkmBjTP/deDBXX4/yLmTDNmmfHAdklR8Pu15kF7VGoQ8XJsM0RB
We0/+xZetEQ/O8Pgft2g+2pMpEww9FjeY5doOIrqHkdGxrDivW+rN8WkgTxspbin
we2FRm3JX/2QSfI1hQwna/fOBoH8kW3pr3GiUotVrsLgagLcvde4pMfFhjFUGy+T
N4Gj4cFOgStsP2qgpl+BISconPciO00HFB6Rur6njwxoPNm6wxgDsQ661abBJr1N
x1w9Df2+Qcu3SYJBODGXFIA4upoyprVnr/2tGsR3RC7NvmDkov9rGbRZiq1JK4Fb
ipqBgc+acEib8IIb5mSScZAdV4/54aWrdoDhxKfJjFnd+wwdmtGLnYTrEwsbk77z
xzvt+I3kcPazDVUTuURe0szVnDuFxyA0olhZyndhKtW5S3uRCmJACIYULDGnOVSS
FHU3r3d/g/rtMq3nuGCsA5MFV9qvW4IQ8PZi2wCRkMZGhuof7khsoC77IEanzFUG
ST47o9rZ+GLKOqKrpFSd3B8hM5aT4Al0Ky7LyxPEz2vWKlRJKaWdCMaUYf2oYqjm
jtmXqlYjzkDuMJxgv1nh4w79w9uaLWBzFf6UWrZz+SabkEnCYPF9PrASJYpLFP4K
ZvO5cYWWquiFx8S4k4MYvaqonkvYTqxQTSn1GJBMAH83EQxKTZhG+Tp9DkQ39ZcY
9EaOUHcGE875sM8iFvqiHP8DIkLPSZZTgxNZKqPbHxUJwbbjetaj4Z46RENDKlTz
tQcnf0cvyCOsejibYCSVsn/9q+l7mFzbrYcdBipQrUZsv1Wi9jmPBMEG7nlk3oVd
8yxo9saN2ENpBQniuB+bH+hUGgw4YodsCnwn7PkSbSkZnGlfHgJMl2l68YujhkWd
5kHEhKUzXe9Ty9MBf3NNX7HTCu43513BXAfNTFVQpb05gK3gikiKtWokeTw6hU10
iZhJ1q1aU4tPDnwE8ff+z1uPFkpc5PMCY41Xz6K9QqvFdStNPFR30X/a2o2uF0sY
B7e0/LTfnIXFWq7upXB5Dssk8M01rI1X/m253JUHKzABfav6ieogqvHYG9jEU1ul
xGh+caeJpJHuktI4bS0PoHZ8ZlApA7HycnUFCBpay/wfN+Kfqy6wHoeJp+PTzA62
ySWVgGNmQ3TTc8SgCq9SHkYXrRWruJtPUvvg1dKOU9g6G6/he1aH75khGlNY/alb
F2zIf84IZgpOWu6ShD7hlNhdJfdM7YAPfn0GAU7Vaw0zBgw1b8r1nwIVL9ff9HI5
whuPWt3Gb04pYdjOlzZPk7neIwZVRd9Um/l89BL0+8nAg7kfkls9bU1OYDbklE45
Iabt1b35vp0CN0qP1Bx/4SuyhAenSPVWJt6TUwDTH53zrtXRkgqNNVZfY8u5hQK6
f+u0f2/i7N3v9u7XJk1f4XRAf4GEjytlJprEbr6K/LjBjOcaLO3dtFkgv4w83weC
1n8XxBiYb7yqkvTPymdCLD58GD0D/dQK229a4kmpgN73vd1pKQVA+pB1Fr5YwDFK
GiBCLgWWLcD+druUH5+6ZpTEVxItGd0v1o+I4UgXpgIK7w+GGVrPS8VTKPM1griU
L9foVMTY/3U3f6P9O/dAnpJ+vbSjP1PhlKWjEuJZfEuLUKjz4oCaQtsaFYcHk/jh
t1afa21Imh4fmvGjQJE6qOKWOoKYIf/c9AAhOlyi6X5X/LrmedKMYozjfYSecv4w
ti33YozQb3zsqGBfo9e2UvhuahEuxtncbieN/Imfw2/3idG+rB3OGUfQzKLKTHEY
/MKXKp6hMM1RcO8CB806SRzhSLS8xrYP3EhjT7hneIwoDSjDRwUXQoONFtD/2OA9
Q0iHe07cL7Ev89/Zg27/JHWk+atPd9KhAmM1x93rFXBFV9tSUGNUdGp9GOmge4Qt
jYePBrrsT6e8vmmkxeQAmxEPt1N3JW1Fi7CLprOdEWrqvHtUc1RHDSNsmDe5fvHd
KnmtoHkvY5lgua04bGm7p1C6csdl8G7iF/vqrR3bXCHAzNGMl0hPkx2eDWQapkOW
J9ntGp4zbD4sF6jmGHKqGmYc6dCDBlfqy6kXG6m4JCiFxY5iOY0Ff3DIggycW3Op
Kt0dATq3lSTxyTmrtusQeg45EcFgUgzAy1MnOgzwVTW64qk6M/DWWU65ULnHL7iy
nufWB2s54qMLlLCDpvKyDG4tJh6R4ARHMyma/SxdnFx1Emz+qluioy0kDmG6dk00
OU5Qee4HzZLfCew0tXs4m//KBwG/55WkQ0IsEOsQB2Zn7FKXY/OC1VvokpvvZ0oX
h/bzfI5fQlLCGtRNo+G6Tme+qPjr5/qOTjREyRFikcHjm4Y5oCGJ0K26plb/BiBm
48IQCojPB4mQV1S5DChVbvCHSPuExJ9vBYxhdu6oYVzUlwjhtfnUFtQqc+1r8m6W
SD0Iu1j96RZQedCoYSdnuKUeTxlaO+uW42leMz9Y3VCv53Q3SN4iiytMrz5udfD7
YPe13CpoptZ7EwYXSI1y64U5+SUPLZ7pxoYl1VZHaqq8zULC5oTdOHP27Cp6UP2C
/AiSphWm7ud2z/1uH3OTtNRdACqjkVBpEpYre18/nyfc0C5RGtDyE8UDdJvO8B9f
CZWBieoEBKLOG/4vgvozClVxDkcNKjwVstaMAFDb/1xM2K/tCP6eZ1+3pyxf7PsZ
IIASmF9GTWoE61IjuFvKlmQULVNm1fO7vXOE0Bj6fGzN4nmYXzn3f/HTrBhSxBZ/
MBPKJYDx1cxodOn8DsiadZiqmiQJWx9oGxwFqXXbob9x6Qy0YaCHPgxI2Lb6YIG6
BHSaxtdOy5AJyg1IETpgGMVK6PYYWbn5GrlnIKXnapwSvdjJfLNGL8WQZU8MAf2D
tm8Q/TQ8y654Q88dle4+t31P5PbqecW35vRtOju3MuSZQfGW6GenULa5lG7KKLCN
G9HOKq6764hUcGFzeQ21fbx0XrzKK9ta5dEInva3tp2vrTWZUbSyEauBRxIaIzYJ
P6aMI5mU9Hb4KSmi4Cf4mQgJNYBWS8tMP5RxbJ0Ua4yXnfIz6H8/7MxDcJD2KdJK
YTqEei7G0IuPdj2KQRBtk2uSPxVe92T3nMhH1Nr1bq6QOPp0rouv9Obcb3eIfwax
igd8uwoOOSI2tseuH8RNYkucsphJb/Sdi9qQnANklbgtSSPBdW84UwAqb0yo8p/2
7tJbCqgKydT9/MtBMbANAXvdDCfkwPRckixVlkvCIsPEXg516g5YhUaF+JmZOBjk
lgiwa9GqixAZADGkBU0i2CKZczbHhnyW8VkqWM6KRd2iJiR2ZaGk5JW2WFQRkmkB
yksQ24flhhTceVbS4UtfpjVZ0z9TCMbXj8pGnmM+77Ya0ouMbAvtmzS5tzl9NG37
a+oJkgC23NnMBjlNDOhMFysnBHf4tyEwFU+ZRgZYRyCDZ1KaffEcaBWtiGlILhBt
4dCF+5nwfR2eqU9LzaI/7Jwuo7WloJ2pO7GzfUv7LVhkM/+ZSHFQhgHC85dnfzLh
RYbDUWLDlKndZlQILTQCPpJrty58P3ITfk7JEHIbH/n/Wufwlx/HgbfKiVTdrL3U
pNA2NPFn3OHLfA2QCKhPyNgwXpedFlVINP7+FdSB6h/BwobHVPYZu1DaSJFKT1Gp
yfDo3aJfXQNe9t8oA/D6ykwVvhj5/CuCS4axuajU44rq5W8OfBpN6mBfxu4o9CzH
wd7Xfcv0MrjyBtxhSxJqFGiV1puY4bJF205MwqjvFRUy6FDg+y3cwKhwDAC+yFdw
RLJNHMbqruARq0rIEzHNuMp487RN4/BC9rOmclg22X+nMl5zMJym0HKvyPWDFdTo
UoCDqQBBBBAx3Y+8RuwWhJ8+haZvmjBOvsUWuhnd7FWXTa/yqWSHLV9iUWMVOkBT
gBTPgsdbF1TXYAmrmuKhnPATF039TzjSVHJsMRyDYA+2xYBogTAUDI6BBnBwm2Pi
j9hlXwoVpMQh0uXePeFCUFsWH8ijxik1wmw7XhiWa8PNOBVchntf7zSg4SH7PH4Z
jl8vrvJ1vC8QGmrG7LSUFMSqaS1OUlE+gJr9uNUej5Vk04R6570YUQ8H2aUQVSAq
9I8B9mA/qYnSTnXiaBmlED782dN2ftZ2bg6At82VENqb3+3CmCwdHxg9NarJb8We
AsrIivFyXoOUIpe8x1pFfiYyo9WjT4yqGAZ46rXqZH2AatCSai45Rg3FBWffYuXZ
GCBZMxEtzSINlwiQh8bP3fEskHPJmXUsYNvQfJ8NQEwOcvLhsxObaJK3ezutz5yF
diZcgQnl7Dj0bSxjodSg57g7vhTt8i3NVtJBixZIECiemX8hGUMB31p2gHxVaWaT
kTWyf4cH3JljImMpbtdmVdycAkQR42IXIr9PIAGaMmVWKJLI4CbI/Pd3fylLpQ6r
hmmXymOHCKQpCQddS+XIyOYOuq95wYlg/1djFvtLAv03/bkSZdezwGOcMm5NZNqX
SGyPN5pLXy3Ef4KI7GRyQ4Gid5LYdLcancsTG+jAmpcW6z5E6rd1lOs2tNHTKACk
SIVYo6HYe4MOL9UlcN1leiLcw60lNFsXdEFPrga0eYnAC8rMW1fiETMkkWfbrXD5
S0+OVIlS54yNwyiaoHhIFjrS4cSWQPVDcc0XmBDr3GLrUW+DithB4LjiniPddIdk
UJSolOiEJuYVdkRW9VyMpqt74LRo3QhxEkPKBbmkZK0Q1Znk14gGuDGTuGvFs/4U
DWHHj+Yh0iPYGf44L83r2vZTXaztExYcthah440klHUIuuKnLYN7PFNemEeA9Fi/
3QFVgpgSWkSvB6OjicJkwgrR4xzWuIAJSZQ7FD8DSsdrf6w5W+ebDQyuJpU8FYD3
A48cbl+UlrcHabsawGnDdpduxSHhyAOfuLNuUIioMWYmnNim8UyMoPmqT1WKkmGF
21/814vcNGD5znIPGmB+eqRAMfU7d1eiX/f8CHOnPwPMacgih981Aw6sF034CfB/
M7qm/+9E6p+GtuQeR+XpTsu5Zqk+iSs0K2KUGOkL2/LOvpQzdaoiIYWOerPRxW+j
yp1VvUt4xpQwFpkurZp1YRYCYcsmd4iJxzbRy/gYjtYGUMRG35IBermfFjDbohf+
YW1br/a1kLsu2ROwVMjf4F4+MxJP0K3tluy3/WsLteEh2Bf8F0W7yzreCfS0rjbF
ecsbrumVItM/uhRWMxaRaE8EqMTvjEXAQH0K87irhRbGuiD0+yCDr2FbJJB9TiLQ
LwB2F1tIdRK9tstLB/vi/kCcn928B6WJUUDnMaC/JrdwjqLoabORjLPW3d/Im378
YyUyg985cg7pbW/cvLUVY7qHV3lTWjIrXRQ8yEspcwVEdf5SmeGKeArqV2p47C0+
GzTcTXuhWMF0qbm6DoKulBbKKtI7HZ7HpM+2ynNcCSedywrbzhuQRE8AOxNsNtw1
NYKqA1W4/9ZrGXbiMB2I7hdCAdnFgpnsR+RdvNW0K7KWHKz6mi7yQHO5oXYmmlYZ
3747LtOBp9QZ69VPfEFgvmHRUfPe96BYWWUuxGC6NE5bOmdXOzLkkmYwjGqTI6fd
h/1tuRWLqNiMt2k56tkqIkbWCv/OTSKb34i4dTuwg0EtOlv1xX8+/dJAGG/s8C7+
hQ2gGFA92G9X5WI8EY4HEbarNd63AnEazOh1pRXA9atiGwKfeRbp3ZU/BxbklHYf
lDgwJdPmKGEBfAwtnTVA59kX0XB7wwnmZubsNOM+d33Z9DD5hC7oC7bJNVJtc7Yj
g+fFGbgvYSfN6S3TAR9azVm058Rk0fCzIEYCXdcx3tM8ZoTTCQKaacf3tPS5Gkty
fN/fnHaziLAXmt0qu0AX0MeIG1dysKSquD6nDAQPPo+y5JyawkU3r1+fIr/Vd2RO
hSHeLelxr2TvFe4aIuIQcMBbmN9YmSNTcW2Ufx5y0fQKIMwMD9kM1cN+1Nq5ZIag
6bWwEPS6ofiLZ6Y4pg1ORnJYkgc9zxInMkQ7WxhUxcWrb/p7lgpySCtqDBmyDObJ
9ix49UONmiLJ1chylQvlAY+Hrh5xcRx2RR7+Fzjm2gVRaEc5/hBUbS8ckvYHTJMV
5Wr68769yhVXGf2C/uDHyKqwzUyK5xnqqOW+i3Ngyssosp9LfOiZXfqiVjJE0Lk5
plY/BJsBd63u+2L5amQ1WK2KWiEl6WJseA0fIrCMBPWQk+XAT375g6GR5ch1g/+W
fHjIsiVdOq6nplrI+hmAQd71srRk7RtrNgWq9AjyNW02Q4dDJ4fYgt163y+zckXV
UtJIxhL+fyZb8wlH9ESY9AnZeqGU37B5Y0INUFbd+cDDyaIoEHTyDwb93b7tAK/r
3MX0ixxgmc1t3LGzMSzP/8M1MqoYP0b6RJAgKIwUzYi7bSMBC3yp44/PYX0p07bu
vwUBxbd8WftqCgS+u1EKTAZHEf/Bb73unLtFxZRmBLxSMo2rHCz2gVt+PgaXbE65
k4XrfDe0WbyA+U0ls9CATwUzn8CGUkSqbsZkLpaTrp0qtBYYz6iHqxa/UPDEFZeK
9eDS9TKdUWoDwNYhdm5K8JP8cn/CLAfUet1DFAl6UwEFyE9KFf38kbLDkV7zLLLd
dCMCgQ0XbYQMfSRGDqpIfZAjD6cbXnfqMp7sAaEl4ysNf21+u7+g0l+tHy70rMxz
g1cjaXhjo2f4OyEyr8zHDhrKvkb20s9n+V8uBRb8pc8PtdVVjOvuNhSgpX7VAMPM
HRKnm78RjNER0cKAPLA/ibOWXCSYrlENQSWBwE/9RzgHw8O1tDCCc62JqdPbpZZN
/c7O8Ee5NHMPi4gKjMTtT1Qbgah/9kY4iI4XvQZzuZkphKuSbgBogWYoau7VpSQ1
uUbqQRClKwAFgFqbsy8CsmEvAzXpnO7Z0b2FkKvUQeWCvBiZy3C9KpBogSixDjzG
SDGbNwzy0v6I16koTRFG2VZa65cI1nHRTLCRmx41z4dOhtQVKhWYp/wOA90vdnWK
P1vbYAL5VrJiSRoRZ10Lj78DTMbf+lCRwdPts53OHKyUKLHTdjf66MCtho4eO/hD
wQUPfQFR4KnFbwZpZv5l7HIN+wrayRUxEsq/FkwhnZpyFjiUpyyPbq8vpWS8s/ev
AO05XZ9JwdOKDlXcvHwH8yMaBFpq93pGKRhlHUKXXsptV/rMOilrd8Veh/7QCIko
Vq+EaA8t/42ywj4bnAemTJmyUcysfq/BXJ4QKudBQRa3MgRXAJ9DQTxcy4Lej0iV
GvA2Wga/D5zvg3aSFhDmGjC14O4qBji3pWhEPD1P2vBUppFxwnVVfx5nbMUCe4S4
mnc9fs/34Ll1Umngf24RQTmOCYfGNfh/v/iNF0uIo3/io9ytAc7I+HWHbJqmOUch
tk1ZDxWDSNQHlgY/84M6z+AKwaNDgv3C2a0VWDhmv0W1ofSPHNRXmQi+mmkW/FtV
q+NEn0gTEhhpa/ETlEhbN4tGx5ffwdWm0MtzsJZAvX9dqSW6j8toqcH3Qp/4eoAg
mDWU1YYzniICaqnmmO3t1QAwNT8NN5sXqVJOQxLLj7ymLOO1zF/5DwlFEFj1jh2D
5n8Bn6FkQk4+U6YWwY9Xu7N+7X9/EQ1QIAcZ2ZV898xo5SDMcEswyHqHXjNY74CN
LOuXDVzqg+vbf8Gqin5KQvAyDf5IHL76zL5O/tzD6NuqHQLVjx0X7Tu0n9U9Hk5P
K6w75t3iqtP+do2eyRZ8BwWH51PsNtbolP1zBJiUdEXik3uWAog6ocB+EtGaq5GW
HN1KJ8Cu5+dVEZTw9B4zkzyXCwjS7h/xpbzz5IXGzWCW2bBn3gCWXnpp71A+Fcyw
h2GZfYSReCmFrHOswKRFca1TTX8IUA/ODhI77GRFzHoLXW1tVTo2CrzVysDcuW6x
V0xzuEsm78P/0zB5YbMJUGX2t6RN37Tdw1q+nUub7fNMKneMUDesK/Ne/K5itWiF
+R64vAWZVYwy6oX6gS0MTdh7xF/5wna2F/7qS0ZddFnaIwcc6QbqsSresFFhWsne
3Xd7fzZIhs1fQFMKMpMmDtwd+QvUVJ5v7E0fZlCv/FMk2vEiEQx1EVOe1b2j/TPY
sn3DHHOyRl1DznC6EPVblZN1Zfs0U9ifxxh43Lpl6KBAlW9HLJMxTo+uLi52zgGL
bKHAEZ324DjP/g5qcGb2TbO5v164iaf0/sx/SVhi/6rzZkLyhD2O5VJ3Ngb6BZBl
uTeLVVnIy1mDuYeEtpO2uMQQdliHplKRM2lO3UzQk2E1b+6/LT9oZ1wxQgmmyk+7
vknwgfifdxiTmT9e1RTSOkdCiYXmpI3nvnn/eA5rCU/HQETnMyGLpxlRjhpsY95Z
ui7DQaM3zH9sJNdiM58S6iJ0lKm95dQbSRRu28g7b7Rf90XEmuJ4oQAKg3Z7NRkk
tHc87mFuAhxgCSbVZHUpe8qPnyTlQRBseLSyxHIyCH0S3kaa9CwCY+/f37DsrYZY
33MrH9rEr0lIZQNqGCy/EM8En3aop0i2JEvAd+fHOPAbgSbR6MASvKAXNggagnuB
Yoy0ih2w2kN2tVU237+OcO1ccgqMnc0E/Ndyzn/ziKiLjjyEtrQWOCCvHY8EPkN3
TLdkHG/WNo6gdS8NO8WTrLUe0MM0Paf+GJ0HhmoP9elMfjlrn1ynWhgSHrsx9FiB
A+/5/HNYEQW/yURrAW7bxgEqPmkDWGJ3Ck45OENVWWSj7KA/9wlPjtejBBFDmTVF
2DFfkDdVXo4DzHm0bmZ/ri2IyEI3ABz6KHfgO1lnQF+xmI9jwru1T5GdloptY+Gg
jX+NAqkqnAyieeaCDJeUVswaUdNeCE88ORUpmJnja2LEx5HZg/29auO+NRbt9Hfx
TpQipTMbtvbIfoREzcEuXrjrMiQ8t3lT9b77KRnc/9KkMFdjnC/MkgegLP2TKFVx
RAfBxpVna/hv75pCnnR1Nd6lihU0Sr/Xief0MOHilFpC77hMDt84pW4IraavFTXp
+JJ6sQxcpKLlNePXnu+BK2f+r3fqNfkWIcVZVbPRbJcTJf3owZB/3/hJZLrQuMV4
bAgRZpJRKBXYPNPmYYHCoj/FiwNJE+HcLxerUytZNfKs5Xs1Z92OfTYllRcc1pwN
6rVNbBchfHWiyauyH1OiM/ahWaLEoIaRTmRErxvYlBnC9nPQisBxTO+GyzC9f8vV
W4aF9rOVZHmoHauooGIVKN94m3pcse9hYI7lXa32IAw2aJq+jFYFNKgHxGCC0yc0
JXbeClXbWl/tk8zH7yzZMAObCLXcczrroNYDHMcJKygIk+n1ODWEE36q7WU7e9vk
JXIiZ9NCXHLRM9yYA5nPZF2ujjLU0fT4KVU/pMn3/5Jg3Y8HgQRZeJ/KHt40DVv1
U4HjL4Y2aCsMs1zhyFBLcqPrHGq2oFYAHI1KUJOJqi0EL/5hhJzA3rAhZvazFlFO
5aMGpMDn7vq9a5wy8tIzu+pp4tVs1FfvJYXlFENDaDFON17h+faqebFuQo7WrOAD
mMnnzkFkffKMqyhYcpDVMvpjVxrSSyu5p4swlNPkrzVzuZKTc3IQqNyoiDntat65
Djb7lsE3cEXeXN1Oi/5o5h8NpHnylc+b4hvGCx1Y61lyPtAho9TfVUC2TwoEgsY1
7Zr8X1Q3UyNspwYEFidGK+FHoPTz+qW8lLvQOR5UCPTQMqfKEvKfa3mx3xDP3/sQ
T7ITDlkqEgNlIJkw2pes6ukf2jX3cM5vO7zDt2nqbCgrHnmBJXA48Gn9ndRHEScA
tUOl1ipSAa/I9KQVqF2fkwpcHsxSfJUgtYM1KZzuxJr9AnoKzp+LVsnWhvhyRf0a
qDk6G/r4SsfJ+L88efnCxlwqffJ1da6FZm9LDu3I6vIqH6ELF7sEnfQlbSXn+jrX
fUZdEr51ZXyHD7/iyneb3sOSO93WAd9U88d7aNREOkKvbeGfypsb/KREj7Rw7xb6
1LyihP0X5q9KQ7sV2NSTmFmSXVP/JxWlzD38QDXmMPdtwxXrEpddvHagdKjg8p+v
QXAUfgpVc2g8I7wIdxc1lyTbuqkNW1bZryNTq7HJqqzzHv5oipmsJOs2tmxIfj9S
ofQlAVI5bmC3OHtTiaqKfyUg8N3Vv6g9Z/YmIi3Az+yvbLQsHYlrmo5EbQaNYPtC
/l6Nx5Q5rdi2pZWGrlg2U4dd0GNdy5ZdLSYWh49E05Us+ZONi1g4eu5FHbg/UE47
0wKHuyRyQsKoiveeketi5u+SzSIReRGCgRo2kMomJ1hTfCz5T9lnwsOKBjO8FvEf
8mDZ8dluJ0dh+LvsryY6dE+vK3DxqzcHaN3B7c0VrfkP41n42wnLFDNZe/lGQpis
VGjb02p74JQ6ODSrOZ739OtbErqNaL0fVDqXL+eXD8FdbEpeTP3fhfnvHeaCJgGd
zjJ5tj5G1MvcVH1942pBDmYiDEAbabyQZgD/n1BT4HsftRe0Wmb3WVhNVp1vSFdw
nKdxaNXXgMP7fUUz3MsAhbY8tPMymQsMDz/AWt6Bti35V6G/MQMlTQdy0+KHBwgP
2Ho8J6On/HV+t8oWNdCFwmCW0rtPNbob6RNnBTDuo1C9TtfhiCmDuayCDyw6RrDj
TWLO2doac8dBDMZCP4ZqJYCDs88BL8eQWeW0jVln5mDsE26kItyZxvw+/+WOy0WD
hFYJz0BXmDKQIFIB7lpzQI2vP6ZigAcCDndZxYBxGGNVbeRYMJn4aV1A+GPADcE9
sreQ15B9PsYAKxTkpxewJwxowlfpqcRYaCnYqdefYaIk7kzugSPq91/o36GGaaZP
DOIxZaCNKsaiNzxKb6B4tsQsPyr0VB8aQYIrWNEwPML5OEoRhKhWl7nR2Qt/rRf2
XOmJCtB1UEIKlsB5eBneHBTai+egAzU3sWO9eKDCLYXiduJ9baSH5kF6gBwkJcUs
PO2HzfNqAL+fznrIn1UwoRTZvnGbP6UCipdunFzSlFxPOrIL284gsxUz0srSW8bT
+h10kyGl5lPuwJzpfVjFmZgmxoV4prLq0OnYMsElBVgzzJgv3uxMU7iasatHg23o
BXjYz88iH58/iIi2Vj/HQWoQlaDcA1AUcZN74VSHy9OyB0xWAjba3csvnjkO9PAn
yT5jZQkAJxxDn28KesexBy8V4ZWgmvFFk03f5InFzTEkiEYKQ7d09UNbe5lDG6rP
wAQ8y3ZhXH6zF9QHUKbOz6tbX7hiHHzYtSHz49UTbwGdI+Gll248s7+a/5hwBtku
qSkf/Ibdh96FIOkrqoAGn33qeMSEjD9PrEAT+lClm1GogKLPMY3EIbaDSMWGFTDQ
cEpf3NkNr0hF0JZeaimLc+SSMLUf6liH6o37LiXjx0DttF0l4bWUwDl2IWMeh4A6
9T9SIeSr3etpL7Lc6j5c/by7Z00ix7pNgI/qkDcp8E8uSvXZNX75lNV5nPy2pTO7
XRIW4VLjsrmb8cKHC/ZtaxL06mjdvojvF+jJ+CVkteIMb+3uPAqEeDD1u63DAT2X
/0bRwW0Kl5dY8UMGxB549S22hsSqz+KNy0Jmku6WKkyLKMbmncNB5CIFLGELnCNK
OtBsPlOCrvONVcWCx22/xw9i+fCKoDscH3hGIbHeY46Gjq8kUv0Nud6clodu2YN6
5R6cU+m/rxXk3IGzQwrZiR4XWFSFaK+ST+ExDHkGKrnXyp8JcGAjat0ZBnb/fYKT
esr+6L6WMoizDr2IN5izoWyEAuYEcSDAOcTKtttR+6XdFg8ntEvTR9kRyXXA4xW1
LpYjhd+CGdiXWFNuxuCoknAKhh/SSWJl4GyfilWRlceP2X6Tn9AQ98U08vVwGrov
n7BfdMoOJ2Ca/Icil/0FwlcjKUU5hveM+MmhiE6cIZZ1ca8N6Lq4UWOfvH0jm51z
jTv9SD0dWDDHb5qgP2PWgOTETdiTXi+pJYZ7/+mBsuEJpqPPPWr40CoE80WcWHal
rOdeiUJgAp0eIscIlmtKC9dmMECLrEB9Y0X20a9x/y2z2ddY2N+AvLHt4z6G+gUI
UA8QM3B49xs6/qLY/lRg01eTMKVq4EHFz0GmnZeGTpHq70qadVwoz2bDUCBzSmL1
LDvx/5yijtL+YaVp/aGroCXxumnz5NYx7ncanmgY9pSZAvImf/NEVwMHEUibgy5n
cY1FJTtAqp++/PwXple6kPDqAhCj/zsZ4UDnuTKKSjyGpDwH32L2bTXXkP2tC/RK
NlgOiyksxx+3mZGjV++OKUsYhc+/DjhTjA66vtxUDkxvWxu2yYS/xiJzgrk0IRJ5
5W6TqbOOCMBGCmX9yzUBtNsE7Jb+pWbUuXH/v7eP/iY5g0FcljCMmgO0PpsQRjFd
yNFREIm1q53EFhjNw3wPyO6djQ4mm99v5Er7I53NG4OJjw2b2cszN0RDQ/S1zDjR
WlCdTB1YzesQxTJvLR44v+FrS0WBI8ZfRrIl8L4wXjDY2GWQMTCUGl4WQ3+J1XJP
CzoWd67jBHBCJitMn9xtsFhS/mSyHC+wbDBbYU0yfvuSYCnwjNWLV8FIbbbQcCNd
irYNm7cpRmdDZxduq07G6HDQvT7PwAuIrnhUusnNAr/wyyBhmXVjUU7pfFyrQjPV
P7cK+WRl0oIiR9pAPTMdiDGmxMCbatlL3sKbjVlJTfcsnhP6uH5xDZBx/aFe4j0F
0PgcgTzBdmtnlAS+yeo3SYx9iSL0SGycoogmgtpBcVKtwVZGc7pa9/job8zOIPNQ
Jg16j4S6gSOkfqNIfxra7sLUteERvDo5ye8WYaUkdkAx3y/nC8WAIRwwThqyL40+
XXqwgdmZAlYU9i+SREop2XcZK07hkzqFMOK8D+hxFm832vt5eC9u0WQmB1/GeKhQ
c9iB+uaLzHCBqoP/EWozwLD/yZUe7c13B4Q8FpPkdzCx58po++5M9XGAgYvYCHyE
w29Bylpi2TEStR3fYnhLPeCGuJeVPHDb3mXdW044kmg52Mhj9S/ZEsSx+hQqdOxL
KUndTpQUd1zjjdP7sGvoPNB3/ftA7nnCYVTDZo6omOZI+tVeltZ9NYgkAMjyPZf7
NlBP9m9f12cYrn93sdkJtvhvbl7GZe82KgOuBazYQFX41N0u2p/F64OU4BzGLMeU
n64J/T3QgtLC6aeiaa0p5yQbgCJBVTHwCEmwz0D0PWHVO1ZBgTDB6kmW1LNzy0kT
xDB6M5YRa61BNAvj737HYKiFfIvs8NjABHdcKupnHjXLLEaJT6x57UhzBzZvI2jL
g9odAkrKXtQYvpOVq1OiBjJD2tgwJ9Nw9YsP63xgbE0zpqhVlmw+LAom5mDambhK
X+z76IiYEA3cCW7ROivqYgx2teyy9F/feK0O557yJKt+l2jjJPxvPXCxw7zdHTq0
n6n2uJ6QBQ5Dr+zIWqCtyeucDnB2xtZ2gZHEXBXcpCevMrNsxgIOIXxKO5vfJvk2
K/iepFyZe8pApkokj5nszKqb56CGC90QgB7VEbRCw+ODvcbfe7cxNhCFk/WCI74P
kdtrZ2qPGBjcpVyxgdwZwDSebqnyGsxGxS61ZfD7UMDHI9Xw6gaSHmmaU8jG5X6Y
9RzfjVQIoS+QqQ1AxLPmu1OZf/GVapTga41Ig07Z116gpv8AszRXVJ00kD3LOp9J
XkVIv69vlwiDB+IypcSIkwsTacX/zxj5IwxJojU7AYWP3LV2YaIYMjO4Bn5KKxXf
44pN4pVa4aTGCpf6HKI8u2i3QnD4quRZXCimeqtb50Y1EfQJDAv8p6ueZzt7wMfq
+ZHjQ+/SoDvj2+KUdgVRtSIlA7tI2zII7yHxCHphFk/7VNNk7/wA6PkAjeKYprJx
EmRFLjZEeKT2pPCtz02DUsejq8o28rw7Ptpyuef0BFpB0I3X96bmr1QahLuGu65c
5HBecEfX3mKUsWc8x8lzaU4R7NuOamBD8jdHa3k4bzZlapytZBdR6UiiLv1wM1pU
MSsqpuhs/ieH8DRUrZpZkQzXj24UqeROkwU9Rm4/IyxmZmTDDb0yCdCvXd6J7TGW
UA5XySxZj7xLc/egT1fC1hNMxkkXBsGd4PajjW9J9xCD0PA2GVpAql3vVgJsqBk2
xBkva8iTYZYHUOnQPQnu+0r6j2ohzV+sPn8cSKF5M2dWmrzr0X4+Y5ksJNoTqDUI
D0uFDoagreFV3lqvpAorRBHb4QMfryacXNLBZaDLJaiLZ7aeI+FW4fIKCzv72kNq
qMVsGPrZUl5qbPHR0Sq0GvX4Y0XZbJ8duoTNMRL/acWyTDSnI2n0DDTRMl+g1guF
urYpesE1b0HEJ2VGcbB533INpRliZJlTmWB9S4RNN7rN+0t4EO+Poe1ilgOkoJsm
bRZl1D6Ad/X4p/2AuI+Pz47mWvRnhyVLqPM1lpTR9sayC5Wu6Gjevca76pg0ZsUM
sV4dy7L2f3ZcJOCi6HuvRCV+Lcvnah9VsquKpkQmJPZMP6MzYNPjDAtqJtINTMQi
IKmFTMCJL+nWKgz+Gxdvq2VLVzdmWX0xNt/bvlJ+PUU4GtHn29t+vxgIAQzUQR7a
ZjjQRgjc2m1MnDnXqvZr0ozkntj+X6cCf3B0D8xUWz0z1jS6M0w1XA/Ncrlytze/
KUKzPZB0iiopuslownLM+BBZkZljNKUB/CSodYCBaxenv2PPAddGvaGQWYJ4G3zP
W/vjNR1mHVnhaAdbJQN2JRJ+cBcqkDSV+08AO7pmzLELnvQfWS3fBgYJZNBIx7Pc
4b2JM0/PBAH7i4huOBb+bAH1L5IZFZ4cmrnlDp5VROfV8XDioHaQ4JzqMqA+EbCG
n5MLgSnM6cXn8sVLTZ/zGLTCKsrAq9vZVyFl46UaWBUKVtTzaI/OPMcRjScfIgem
I5SOSMLIQ1TehEeaofP+YOoL185VIRpI5WUS8gQweRPoWgAsJRwL6m9E14Ed9HZO
weDG8lgyeWj1LKcmxajLBbjSHZkbqSMl8kdlK+cFicZjuIQGf7K3MBAfu+alfvsI
xV6Xq069RexU9jqAUNxirg6rgPNROEvV4+qDOdHnh8VDt4MWS2sUpjgt/oCyJV59
e4Fa0HAE8by1L74DaBzKWmjfr1Fw/rUwbIQCnZdx82GmAQrT26DoFI8AKDz3A7DX
fZvMVMFk+3sX/zFPZLVN5ZLjAQSSFP2obmybwdLJd2aPL+mId8HpgSecV5h3HFP8
vR6BypNNe+gHfJeQkferebDumVWI/IqgQI0LZCm4J6Ub6xtc9vjYTZK/OVREos4p
RBWuE5Y1mgWIUELMYpPu1pDvq2SrR+gGhVw3PxEzd2wun/7enbu5qr+afRDaG4sP
s0krYS6Vp5g18VHtffmhOoM64CLaDnndQCIqUbIYBYbctd7tJj1joCFoMAKyhDcR
pFOIUMvx51B4c2QG8Ij9WSbok4pC/svfHvTstpcJNTW9tNmqCO1cTsMIp2+trcY8
ow5p/xwli6hoB3BO8v2H5G6vgVEbQ/8t0xoAjVMvs1mdhU7RLwv8vuBmdIifUByG
cCNjkf0TcIGVQDGlBJNwWE2EXaIn/R+e6OWWJh+wFVYnkX6v6W/YXiR9Il+1/0Xd
qMIpUmLzdf0/zbgYhFyy7WfzHIx5bj6FrTbPOsVNECqyzmWN9AwvU0BAkd1LT/hS
c0ktG9LrJ6SzVLTRvPteLcogpEGqFE1WSFsB+DAEXQRfcP8EhvBvtRD+8hfk38tv
Poen8iKTvhKU4TqWbneljYa2qBjbDHt0CF1TOQcozPtUo6fxHThkOHKPtU9ie1l8
SsJf+KAm38KjbW0d12dZN7bpTrCDTDR/vr1Os5QO2yyGArPwZQV8ag4zoTi3CECe
kSkwmhwD6sb5wxOqFM4PIJAXlkTWLpXg1/nrAf2e3ZnTimFq/fAcl1xVdGmfjlc8
j+Y6tgw+s4RchWW4blVqjJJt4eIHvOuS+lVO60mE00KFqVnWHFd0AJFSIz2DsOqk
xuS/Xo6eYBHLZ1CSWz2+Yzn0GsazDHwnEMU34A8yg/OG74afgH6mSHf7kceP2Vqk
bygUFAlWbMtdztVwrvyld2BSxJRGxZvSNWIJsbTTRz+fiYf4uCRupxt9HPjkL4Nv
9H2MdwLQ4Fuz8XjyKMh940dzbxNHR9ygCL0hLF0w7QtwQnn5btUkzMrxsh3y5a2y
Y/ve3mafv84ZNG0WlQtm/QbzDaXPp7rzPh/yMh9hgEu5aVP3ohdcwy1TnorlPxXZ
z2OAJwA9/UN+4emS5N1PaoQa8HcvOfou50ZPaA8dkwzTJhj0TInSa5FjGesyMmjH
Ed/t52c6CDSyfquyvNtKUuWuSYkEnW4RkZWU5LjPXca8mreDwiy9kFY6pT+MqWG3
8AIs2jqt4ecpHlx6pSjbzJZi8jEVlLphYRk6A3xaInlZuTEU3OLgdwnLel8XGTwB
evt9UkS1OEzDErgHltwQxUZ2V7m9PybfZxasXA96+OxyLONBPkRxDIcn93gHmx5c
afQPhH61OrMrrIaJ8C8Gg4iU4P2qPup6KyP5kqpnUM8v7paVYLsdoP25zcRSWUC5
qkpGcnFe6fCad6zEgRqs7H7XTC3PMFtq/xDnVr4NRw9WJosNHQQY1F/h/rUbwcRI
mXUV6iWtzarNH/pZRBxy4Fe8rcH40Hm7+cNVPMWj+oB7nhAOJiN2+vQS9XLYozMC
qcsKgEqcM3G9g+SLzxyk3LquS0+GQ0LDFNddWAdlSki/paaxF/EUYWwlkP5BdLVR
ASxetrLDHhR1pPp+QFUXTiQnEo4YnYe0pBYmPOcIkHzWkdJ/6CoHAFwjyxgIYCM0
SSFE3CgV1Jf8cfyHUeKoj6ByJ4Mxjf1hQYwEJ+P3xF/Z5tZVU9eblwELGzEvHB3p
KIGTcKBfEnK+WiiYW606GmmP9q4y/kx1pkLmtwTfyfruLMBVnBK+MsQKJWRz2yvV
rwM5Pgd2mB3ZRbZEU94+GknPuo2fOhGpY+Rv4MDHXtZ1tLB4C18ZybRyJyN/Y70q
57OWn/D+lpQkv6RI0YYdpooiGhw2z7qbTjm0UZo4ofgZziCVPblRDS2xfeZdbN7c
gajW2VIHLjiwydSUbQR9VbxkDun1zC2yZMiRVFCx54ruKN1Ptfitk1m4VQZYJu0/
KMxlAFJu/g5inIdYUqmBzrN3QFyfJQT1O8kKcyJBvlA52wLaAvMOBGKBQ81qwoPE
/FCiohe6LlakrbY+FoQ/tYD8nb0xTJi2V4Y8pX3xpk7anGq75dW0UllCuhAXpbev
xa1f16AfROpXfjtLY6aGUhbrW3PCGXsZWv7EfTBeaqPL3trcjF+7eauPoNsp5P97
uryIAk9DePODJcPk3w06IkXqmqqhb8fPM/l8l9d/tfgaFfqCUZDXafSY+NebBBBE
GMYaY9fAWWWM0jhjiS3ZivbKKDDei6HL3FuhdnT+KD7y9RK88JMvLzJTk2o8mITv
2IDNF6cM2skbmQO2FplQwCZcGMHJpBdywHdSKBoT0mv0x7MklWUWrJlkZrDF0EJ1
UIWsZj7OuJuSguErOIkPGCNJwYadfpLyoUjVElt1JWL6whFX2kVeT7uG9oM6HNwV
EVdkuRFg17+kpQaOhQAU7xfG6B+F3K3aaU12prg2eUkEaXNsv9BTOQ6kDGs0bzeL
hkHnWnbcQW3ms3BfmrrqXnN9XnvUqTZqCdKiOK7M7otgst77/eZUGZUF9AROSESl
Z7KmJAOs8N1q4I09t9qWnLmU6uoHZPA+t2VocN74mXcYxUkderhn2zFJoTMcQbKM
883o75s3MAD8Ol4Sc8rdC2+kgnnVDgA54O8Mpqk6x6zR0xOXJjesYUq+bd8+6bjO
LU9ulXmCRAH61LSogTAuhuwD6NeMM5WKzLjEcxZPGIxFjUo8EIm3cFSy0C6K04fk
G5Vxn+gYiuCkw6zP9/ITLLFXBeMmxKIB0UcVlNsjZI4pAVFQEXNugv0AFBTVb1T6
aSCoqGWZA70PFG7BP20E49D8sXOG4+UFcrABGgmh9F9ewp+n6L1bIw4iu31cHAVG
Z2VLWBYiL5lPNgiBA/EAo4b7866yFg5WaIzxDKi4gYtK2A5Rty0jDye8VV8EkJnc
/FPHBuCDMjsC/S2NVmJx3nXmsR0UyGQ59S1AC870UES7NFhZKo/nowFzJXPomV/D
GOJLO6O4m/PND9+YlNxmMfrzQh3JnQMJIjB5u62e3Ib8mitH0TOmo04q/XxsLS9A
us95zHg7zh7AP6q7k4M16j9zA13OmbtNRZ2TVnNVqHlfuTEs6YwcJ1Vdjt3gJxIM
EWkExQmqOqCLQAoDuY75+NF3Z40HNxGf3sTr9NdSeRYO5GWUv8+BGFGfvTm+BM1G
UgZomMH/JxHtmxiwtGdhmuCh4djBs8WxH2/YYlpgk9bTxrNOjaw5ojTyK19J/6ir
9kiFlSX4NfoPPVAUj9F3lhnlI7W//NqT9pi0HOycili7U6daWRr5I7mBUBsJ62F8
+m0LXvOcWCluHogKBawt1QP6Ei1nE5iJzRsk3gkqBrIYKefuZ4I8Xzj138Pqn2Bl
YAgNp/ak988aZCiOQ8jONqaRZi1cB04wQb0RhwQswB0SYBppcj+Y5V+tUzx9dlnM
ilXLtgpMgxhP917OpN9aXu5LMSWQ89JYfCHjKEYInhWmeJbyrQUvCPR7ZBjuvYVq
CVODWPvRY0RteKodJ7RfczTgG/TB4Sy6P633TTn2EYu1Q15I0MFWVVau5w8WbQoc
0JnTuVHVI90AgLR6P8j15pIvMmBd1vQDsCBUZ1afkdNcomHKIMwrLpkP5Wa4j3lj
Bk131rnDCfyZrCUQo+uZN/gj4pTA0NfvnnqjIdT/nrFCOk2ecX7FpG5ilD3IvlfF
ogXE/wMTN9TJNrcPe6Tknt0Bg7ywGbeJPnJHAJO9jX5IoqWoJ52vwCfBpsXzQcD6
oEYdc3Ip1coS+XIFr4oyQUKZDx8JSduOISp9jrr5s00lN6saYQyz6oGIve7jnP6X
wxQCFFYp2epFqEPcxt9adIWaRl8pDxBD+zfqKuvklb0BgF+ILvo/Wa+mlkOQmDZv
zYGsw9LJyM6Fm+mShRT5mz7IYOqNXEMLDywoMeEHlNTMaD82HlZ9p/Js8FuxYOhM
oic9dctB+4tsVPdooaAlh02jgdZGUytLtMXtFCpiCy0RBmahyqgCQCoO4SrluubC
ISxZ9xAk1NCQEzWU7ambPDT4eThhwjb8S8CE5MSSahZLHOr/YLcPqO+q7gV0CdaD
p/CbEEGHbTykOvpYhHVQs/JNmUNTOlVzeRfPTEk2MW4ef7EnJaWw/DrEMtAg1DsN
DmBv7YyzoG3jDZ4pfTrLmebCx3L/5KMzh505L3jFWrUboe61w539MstE8YawwG8j
grmSzh9oEMMntGudIJifkYtmthvTB1keo/E/NNZOcwT1mIlJOZWYrv9pRUxFGecB
IaGEZu9uorlKX9O77s26iwe0HDPHvn3xj/RtEjpJ36CvL7lYUrytHiB4iVt0nMyx
yQb6KHe+8be5DnkQYXmDEILURg18rVfcM6S59vANpfTmH1Zs1y6LZb8OI+f+rlvo
ULqFdRppBvKK36rpHP5QM3R7IxpFi098ZG5slv6WZEYwCpsJ3rdauWbqsWR1uIho
HjVRa0joTTG07p2TiHfAcBPI7G42AOEvTN9OgaR09XlfzEKJA232Lt5Nf+jAv/cm
q6A9wK0/ODL8voVPqCJfP3IYn2jwxQdjOgArKjT5dNgHah/93elKMaRX+DF4ZEYg
/vDQez7GX1Dk6+Yj5UHFSG+ErDYikK8y9K+uEQ+aaYi/S35hcs8NOSAiwlUsaw+g
cKnbuIa1CtLvVJAPHobSXLgWKI/FJ3PwwQ0/a3jnWcxzjKyNFghJ9Uv+IviAPMPe
j/BTcxNkvkVXNcFdGr8zN8WPzELeIswkViHYKdDtajT+T4+69ur7rhSZM3Xf/jNO
hsVMszyDAANUWnBOXFOFNDmOD8O7WCg9+c598M6pzenHMA7baQscDP4bGbj3tS7v
FnKPEDZMzH75hhw6LBQWiXLLPrPAR+Msv7cNt5cShyW2e2XqQeCeUB8kaXjZ8pAn
mpMVU1D/tRThgXWRZrLQns/liiq4PVqhXVDF3yNvrS24kr3xtH9f/E/9WgtI/X9t
ZkUMk7NDaOWs71BjcUmTkbeyQASmomqDqWFmNvyZk0xwKk2kuYPot3ojySESyx3q
BnkFsEQdz0kAXDUZP3tUQJa5uW3iq+j3zWt5APeT1Du1P6QHd9mitzLTBkPYb5qs
Ck2Od9KsAHLE/GDyDrv6D9FCl1nO7vahZGrSodpMoCMXUOFNTt5PJeJ4YqZQoAsf
lkgsH/6gz/9UjLhz5B/xx9cn8mFBNYqThuawmPY9jQgQWW7/R2Wn8/kIS8qZBrBG
LHWnZKlwfR+2Yq1UXodandztTuhSfGPR1y4F1ZiMxlGXc/vzFQmZAmaoTf2XRze0
Zg5BMu5p8wDd//+NKh1slR72vTleqDT+qM/7BKSHwQe/xWF8Tg50vdNFFjBV+eS/
iL/arIXmhI8yTSgdqT+Pd5w82toXBGVTEjtndOGt45ICahMFvD2Iz4xEgonSn+hJ
P2Am0DLAdLKu/6PLl6d+em9B4IJFF2sS7UPvCMB8iE+racgWoR6Pg+6y7D/NNJYS
aD1B8Oy4RmXeombLM2TPQ/nKPwGbCfU4wEY03Kj7htWJe20hBuMFavouZh+P6qze
q7kaPJHZhq7BIa35kbnJpD/Hp6X3owauxaXH1PuS+kBcQ6LijLDmnwpaSDs8ba96
EunRxV4/wm3IAuA42I3+9TEeaI2IgzBxA7/pgdSdI8w5hdtGQK0pUNleUEY6Wa95
C5LxlqYURnMrGl+MHlheVxhjSoGLRF2BSK72pJjjkwgXtpSuKY6mvbnZGBZ6O+Ek
hdO840t5ziMxf27XL9+UZkc2gYcj5UxMy9anJ6mchoRJAzCGP+/I/ZcU1z4xVmQR
rr+7rzig1g8xh17QLeo1kQd6zj4m+hrCBvk8PaU9Tbs04Uk7Dur6DeFflZsAJgtN
tMMU5VXqsLd4Htu5Jl/NpZyHrKCLwheZ2OPvIfadPrwecoMIo/DyunBQNOVCaam5
6Sd78lmzUeZZLPHAqxG/INu6mAukPy0WHbr5g+YLC9+/UrZGdN4cvEIKsy1zvfU2
3f+xj4WR9Bgj+J3Be8McX+wOgdMOmfxmvEDMMdelnI98wtkSXPXf5azSsruCaqzD
PQbb2D4S1t4AJfx3HMToGK+IGH2GrRNIZSpYKHAQjjfMB5T6QS+KibSOz8bbfvST
42DzzFR4pxfUVH42Ee6oWrGh2jtv0a/fBc58tNhnEVBkiZkBwUj7ikhtNKKLR3EZ
APC0hxwIEPFDu2As8RgzD45Q2ueAlyYnPL7crWPRbPH92bpvb+7feYIx0ws+rrZw
Js4ZCgH1k32y6ZJER21SXesN7IJQ0tfNW1P6ljc8AXJYsQJsUVkfTOf8g5by939n
x3vr6V+XsKmP2MSTaAowxQP8dvKKYuYaG2blUsbIGeAZ7f2LihR7A/pv1UTGypxr
0xMrBThf/dzIajoUCgCvnlF5AYSLNt2yFqL5qQsVgOgY1XTuMUbeCahuthQ14CuS
6g775HNOSKFJ+oZR5tX6UK6Hp8K5lp19xbjbocVPqF6r0Wt86Euba1xP+nJsLB15
xGMcRTA46SpCTXETXeTjfI7h/IHHZ0v5J5IsoUehtWSzi8MIiPHlboHLxJD7zvPl
Te3kl+c283leZUA/TG6ApMXarA8Bt4dYKjOL1BdxNNIfkHnaW1kNAQJ4WCjxiH9m
IxvHTY5ZgrW1VBk+/wp5cbWK0tHnRgIRC5g8b+FNm5AkOruAP9eOKSoD5x45ssge
FLBuflDd+GAqH5lxYzfT2cU5Y/kJk/QV16hWFIU5ZK2D1hlCdrNZ6PDNyCn40tHn
0H3QCkMxqnZ6rD6/u0ofzlO6tkkI/XX1bTBxT1gprGEQ01b8TQICi29QwiDp7Zi7
HQZHgDdFDhjK+wz5pxY4qOtLtZfXfpqekvpLmjKm2w5stZHOAqjp2RhcIlsvgMup
MomomCSLHuJfz0IzXO9VA+v8Wty1DSEJBqGTbYVAoH2wwFRyYrAsyi4nk+gbXcL+
2TxpXyMfg0Q1f1uVjRA7T9GYN5sUqCUf8hmadEmYKcpAdL2hLrdig3oCSCGKRNSr
T88VApENC4QviW55WOEAGSfsCUp8emfxpVUfEns5MihFWba0ru+1Al8e8IV2/ZiN
FUspKfHty8H1VT8aln9lWZEZi74+29lyK0x3+3BGki1nHem+Ki4PU7VsFo7j0KNJ
rTkzVgynBrHRsroKM6JMu+f9NNzWktSgexYBbcpke7ZcxqBvsiIrQtAWp2dG3FGO
2f6J6SjXj32qCY2QR8cEPbW+TkZDHAbtC6lNBBHgA9nrAXXQ+wEOJV0MHBYhjtNp
guMcREelPRi3viZF3OH3aDcImO3euFS4xHwco5KBQ2G3qdA1u8VwPttF5UfhNG45
lSoF7gU6pWYsbOjDZwoshAx2L3764ntMIhIog9Zbxo7/mklGmAPQLSPHQ0DxajhM
EgV8OoiBX3Hib1xr9PGubaOamwXfptZ9ATwFmjR3Fr2tjEnGdMIeMJF+zA1lKZo3
LwxW+Wz7KSa+xseyMvGgxkX2tuV4NMlDsTy2JhRFg6PoUN9zB7/wILviEaBrpMop
kB2d6ivuYD6Gkggkfy67biKDSJep9qNWkguGfSAf8IO8KgfFoqQYMbftdri8WLiZ
lA3UuplS2sDEXRcW/lPKvdStEMNqsAxmINn+gtu4/igfxr1bEeMgO0JfQ7wXD9Yj
l20MQu19Sao0cHMycsvbw3m3nxvB/NzcFoGCEVqf2DFFhCxTcrJ9OuxgvAor66wN
IXU3sQXGzvm7xguhOLawITfPnI7ig363FmOyIZGKEeeRS2VBMAyekTFojrG1zG6u
J81yJfMzyk/8J4+M0qE3jq6twa+eEbrHYH+qNt3FU9VPu+HuBy0rUgfRAzN85xT8
U4dqRDtWXLSMOPZvJenFdDck8mVGWmezb1M8TC8JR4ygMOB9fpy2sb9qn3LJ6BYv
tJ/w/RIgVv+X+MLq/2RGv7/LvIjeRgBkKm90uwB/6ew3Dwjl1/Emtisom8eB1iuk
2Q6gpcrujNkbFrzvwc7oYMc5ROpsalITwOOZPk9i/1vrf6vQquwLCpynJ46jctS8
Wy2g6JpA0R5/4b6WZjELoYqYwSAvIo/n6lSclRUVv5EQy873wooU/wT1pZ8VhcAg
CIRJJQmxjHbipCHfYtXOQMBEJHP2kcnQZTDdZa5vYNHGZ7eYkY8TUks7vxDrNUU1
fEQyjMZ3oDVTBvlQfGXeQ5nQVcXdM8sfx/7Tn4LFYXL2VVqkl6R6Kx8WWmJ531e3
sOJpHWDlZpi9IqD5HoKFzaINV+K2Fw3hfPDPGQZjExiYe9lsDylYOIqYjpuaF12P
t11NQ2inWfAgfTjhTzK0nn5VCAyC8HLGmel3pcVEIx80OdQV5iF7qq4JG2pscLJy
/xPWLPP1ILLHydst+5H5cY9SbaaTyXE2eYnEJphfsO6ghhPtPoI/o++hZ4/IDPKo
hKtE7aO6gPpJEM880iMcCLOi4LfCmtal/qs/eIBb2yk2PvN6W/olz+q931PfvNDv
Nmfb8KPUmV6tLG1gDdq7km0cslGZ4RigipyKM4ZbyL3IGUVJapzhasq1crnOwyGb
X//QxFQ3c79xqUetLunIMvSsd/rVOebqsKdAdOoxcbTWXPzxhIzkijRWMofb9+NY
+B/F30TRYzvrw4af32XMdkF3k9JzNWIgtS+PpdxvmwT/bhz6E8YRHj6s49yY98yS
Zbgvyl+MicpV0+qz2ALHYe5f3g4xYPCvQu50UcQt+pScDOKedPYi6oZk2XQk5mc/
3ooqfxuauY75jxmBbXhFl2kLbMRxca8+3ulGZB0xQmYhot7/sAHsQcDIilQ4B5uk
bWjMnly8XFC3EOHu/lClOOKwNJncfgfLo+ay1a2xszWFSlb/ApOXGFrJJw2fZaHh
kONdj8YjazacjdZ5VH7MIUz1FDJHporj8qdCkI53u5HSRLHXziAjaoKNDo61w4H9
ieWhGeb23yUDPWQwug1BSRKcYPua8TMrZ22kcfPTlajYAqm8hsDl94KkYbB8MW3B
6b6aK/oohF/etf5saApom1cCnde2xstv3d0X3Ex0+V63XHN7JdjyWSLOTNJ9whpL
tWE88ZiPAQfUtr0Winghz1rEYiNdOnpY9YZT6A9xS8COivV8SwuCWLaHonPixy6w
rgxoxYTTewDnSL+5FTlYB0kGtalRD6Bf0+cUYdRP5R+OiE3w4L/4c3G+MfB0YOwd
6wV3zl7WWOuwulyUzp751FihOI4JQEZNm9BTJHSAv7V5UjkFN84L8R75qLSeYljs
VgN4U+laOZ5TyFgpIFw4EZyw0O6xE6bRIdVTtGsXAI3ni+vgvURcgsixBP2gV9ld
qqDXnzUW+dohLi9BW2Wa0dCrutlN2VZO5vxPlkP6VNijjbvcYbqIs/9gLk0xU1X7
Ta9wdkil83rEOEIVVluNhaGQf6xJsfiL5cRtlmJBL+nGiQY8NwpFC7kK/CnUA0ws
xKbzWhbuAXv4f9OsKof40VgIf5kghf5LnLCB4myElamfQaqKfTPU4+jjPPLGJFic
xpRfFXXZbK3PhFkJPy0zFUT3FbjvN0E+MGnI49AHOY8EHjVKo7eI9wsqCOMSHZGz
iem45OZCUVIghJxJvkVawUjAZRZoVyofWuY2jNq2JgU6o3fZZLlOQjcL+jFJJtS0
miU9K0t8jtw0CxFmYePeGhqbcCsfl87D9NYXc1i2M0dUPUHJ6MKKwJogtXHUt1ML
OZXb0ShJRKDzv87C3wtF7hEJ3dsHmSRK0C6DBn1pO49hsExjkXN0dMefxgHbsUHi
zGlpCsJ4k6VGY2BZnpgE/B14j85hJS79OWP41/D5b71XzhZkSncMv1ScIpHHekVm
d2GqBmQ7LKRgEgcnT/d4Qa+TLQIP5F2TfqZOKCBa9aTZgPI2H+Ieb1exsCQom9mN
Jf1EUu32Uv37oMrYUzUHMlLs9/gOywWm5qxuPlCxcNRQNrdBbTLU1SBY2uvx6u/x
wKPOEvryC6aw+FVzwZU6I+0Xxexir8foOC8EiJ1X/L463jZ5Zd6ckJ5hJjuG41JF
97B0htHN5/EALCOfhatha9s4CxbQApT90wVk6nWJUkDjwjwUGpyXgF7oVYLL7ATc
7+fhxzet5f2wQFa0W1urNtgV5/yAx4CyezzBfiwyPDkH0H1JYWTrP85BvZpzu7G0
CHd8oyzKooQ1HTdd3WkrFcxtU0u3TcF8QlfNfgmfgy1n6vkanPLtAzAfT3Vn793j
OPU7KYsBbYP+0b1cvrFrkNd17idHwO37tieSwD6tip2RWPKBJjWu6Jkw8kSel6Ff
0JzAT5TWVYSanRDiC2rklh9wemWLrfKlGF5yhsRAQaoyNHu+7xQltOP9HBcySOEp
igxve50ck6zrc0VqkWXICZ9ukfmpjq/EZnAPrRVt57nTUBdP+nEfhqnqsgxmVICf
7PIZ/6MLzw7H7vJQjTDfWywFrHBATOr2H996gw6gRMTq4ZIqtYoAOkngHoXfkDv8
JdgKP3xwMTJm33FW7j7O0X+KE4zkZiLyNVAac6UKwkOcLgBN1fA6/oKQI09ltMek
BcoJHe1HjrRL8wubY91T6QkEbDwEvFfQXDyOcFuqI9h/6E+7RKNQ50gUi22Zn0Nu
7RFsCzHDWfP1829RMdjqt/OGryP+MHtBpyOd9dOV6IaC8MkifqEcJAR0Ez4Fl5ru
9lsQ5xdX1sMQ2YpaybzHjJGloselcAnbHYNju0vB9Rk9TEK2NEnurMi6yVRzrZ6x
kYKha/8IcRa4PDGjZPKOX5h2jrGl4b/X+ya8r9ey6VQDMfS4dMo23/Y/KmmuUhWf
kmsnfvZwibETozVXSlxZ+1BDNJTicwQO6ckJAEJ6xne3c/A6zSnvZ1X1/ZfYsMMW
iyF+d+a45WFPijjaJoSkKtGO0xYAd78cS1uM0IUrJtkR1tHHl2YE7w47+hTFxZkF
DMiPF8/I6WUr9TvGgOloZCPbX4xAqy44j9Mk4Gxy0z88UjW2xfax3EEzw/s+KHKS
9Kf6NnZzM5uyoObvDXoH37IfGXDSu3cXHDuQtjwNcL+WJzUTjGHXdTb/sNIIGW5K
LwOrmbe0/EG1TzgpT2c0j5CUkvcaIuP1MPp/2QzIPARDLvS5G0OoYjSgu4PNn/XX
IMOoulcU5I38N6OUX0YVsTiMbV3eY/nMhbfZVnXOeRT9atwuM/24Sv5IMYLFUMGR
AFta+4B9xBtGhf9PT8iCNBt4keLvSifjaoXOw2HHo1L9sp8ewZHKzQIonGpfJzVs
AdMyxEfbmOJos2gx+OqMW0+aoMEvsBtDjTcxfC8Gdmeo03xeTbYdoZRZy/EqgIle
jjezwiUignON0bf+SWhBKvYabOOP19+iWC9VnoiVf3Pehn8jKLddLk2+kFKi3jpo
4HWO9rxJ1Ym56as1Bh6CIPvUr0oDOZYDMZrKthSIgeyKzYWZj3vJnEQwvi+MNZbp
sX3YLEPm8nej5DFDk0dOPFMgHYtbavhxdcsQKRJrILfnjgDT8W6EefY653L/7bjX
8o4Q94ro+CXw+7E2JY+k35MtCI88Xn2WclV6jOHo+rN87Oq0kqZhXHir3omrGEwz
SJeE4wCIEno4ua3Xpj3DeQg3gu+OzaVk/oH9FdJ9/8DvNSYUgQrF32a0ycyQ1aBM
QN/f4zMioe1x1C8CRrpV2KhcUyi6RaqdKvWr3ILLe4H+MPPyIGv/Nko3QBh1GYtY
8ytgmNO96DiS48pquZ9iplopWpWzjGFxXDrruBOvehBwv0lzLcwZIJN9Sqk7LjQK
IZ/Dw0xB74ubpcv71Ntpmg2NRiIqw3b5Exilzj25rAd+QVyDyTdaLXDJGUTLCVAC
5sanOHfEkuUD7/MAI42twRHgS0hKZakKDnpOups/bg4p0iJ7npD+Nw7GGm7QMu5f
MWRr93ELN2TyfdvzV+OICkdI+uGeAccynQj3lUCi8SySOYCRmvAKyZlwPhfy0ccI
5LBadsojHKaBA2vo13LItHAl9KXYSYPkEC8TR6bi3ko0PymqwwssbJo0LmVExIfg
HJpHjFK1jhQR05TrEKBO+LjdxJ7o3KBizy3DgESuTK9UUaVKX+phlXy8I/mG5Nfe
SeTHqzdQM9Fluy8o7eU4zkX3yivX1jFW3yUovr7+Ysuq4Cesu7E7+JX3Z0JLntVD
X/3PsRhTOxt74QM5a4kdsPWVhmTYgo2Mi1h0s6WIhkzdO4fssai4qBo+eCkhJspi
7MWl0oFlvf0GmY8tmaqTZ5m5vxPOU0fLUoZCf8GZkLULcRB4yOHSutwElooG8j2t
KI1l8s6f2UgJjmciLsUDFagmVPQCchyTxkkVyCCbngV0Nw9RoRdJAvpIkF1gLNWE
JA8lFVO7Oru9rtRcaXBEsybFcaZFI4aPtUPhgQiWak3PuSW869xvAXlvDceuPv5i
aoir5JnbEkccadf1ZmbHV52GYifcXHW5OTkdEKJVdK0cvOQTVx5nwE4Io4aeGVCE
qcTwcL2j/DHoSxfLDjTXr8TgR1RQlvcIVg7EyJajPIPfyvHGFPosGyqkUbsVG4oI
5z34cTKiErJEPMCkRf8OaiGuCSxQqlqLg77K7KhCgYlJQ12ZPsSZ6OwI2daZ9bUj
F7hYvCUKjm1VKtZa7wvWqU3g4EbuhPCwjqW1UiFvrVhDPoZjvc577P1t0Vzw/0Sl
HSzcljC8sWfGQZyx5Sijb9VQeI7FBEc+W/62CvtsD5SEn97/KjhyvX5D8HDdgxl8
Ymxr9UQ4dPut/jIOURpJUx1xDuJ75vo+l4bi87iXnOqNZOUNMQ8wkzqJQkPZ8Jz/
Gwh7Jr65SM8Hw5VkKeMSdx7HjP8rWsYiTxAGDld4d4zRNS/blLWIyYSTd8WmW33z
2qI2If79Gvv1hRT0sydKI5wJY6PcZ6QiieLg2X+K2bOSDZAGzzABUNYHXMRtDtkk
H4flPrKlPIrQMEu3kIhngql45+7kejXjULuLkjfYzylkARkI+PG3eBZunI5xjvQv
yCpOBO49F/+8RIocYG+gFxemdEIsa8v3IYGSPHahttGXcuxDP6tw9YBFNXAH8Sk0
bzUy0CbTcH4ibsQANsWEt++SewJtXyZVL423KBEnBfeU3INEOlBHFYHU1O0zOlON
y3mXbUudSXNt0f3KXURvfIC+WAIBtnrCsjjZKgBkQWLHklmr0hsEA22fU1wTLyZi
JaeRr+4u8r1mss5cKPQou8JmWYoyPtceCehqfBT+ElgspJO5Rvt5M6YWHB8nudXT
4g5TOLIWQfvbsl7LnJhAQByFHS4BUfvzTAs00buTK9MsEXzi7v810wWYCUiZ+Y2p
/cBvqZv1CLkGnp7AzMNhKaC3jWCKk5fmrm/RQYGO8MJvMMBfrD5oJr07UW9E5YZC
FV4TNwgTU+YuUQETypfKmcbDd+gM4OStyezwtyuiTqVC1U//fxVFBm21OXGA2+YT
LpohyBX2dh+MSQIwxCqqBj9rC8zut3YH/xTJ08tQO3G75PWijjRwwQPvbBgYw3Aj
ww/EzcYMVTGF+PrwEJin4Js1q6QopkBHpHXnNTUl1QyhSHj+LQeHJlQrqd7B64Do
XMOIx3aniCqtwgcvyViPfh6lMLyIQUPrmVn20gcRhxnjDFTq8Qr0ggJx2BaMUP6l
NQjo0S2KJx8gN78aza3ztkLCAbgFJvytK+gaB43Z/FVF0YABCl5W9b41nWQYQ3zm
xm3ddUVZWZNW0ouwRLXycLYK4ujuBWYcj+OVfg67oS5RvVJ3k5YoHo6luSX//6pQ
o50Ns7YggyN+HAo2ExvHvqf2IypVdvGPFEhvJdI/S/zjMniTgsxkq3Epcjp/z+KJ
SZksuHqqmc9heJQ6GR4mfIC8ut+4LJ77R3vioaQMKvulpP6JxJm29GuFw9bjHpmh
kEz3skBo8HskCIwQirlgmuFLXbCipdYbdJcyy5jXsW5MXS+2qOFUCbPPehm6FLNW
w1f912ETy2ofG2zHF8KHlwdYmxJqfoQG401oWUE3q3upMfx0aHL6XwiPaWF5/5h/
hFk+aROExV8uFfGwnjWfRy5dBdAGNWDB6WUlrZPyD7hXtmOrKMQMbo7VocU9Jrgx
GZEJ+QSWvzhywlrhdv8mEIN1x6B7eetKa1R/2fMeBilZbT+qlAI1pgyakGurMHBH
AZmBC+nF67X/iuUOJ7OfQRyrE9NK41G6CNsTUSvjiKYsR33IvShWzLGkOuArUjaW
Di0A2V/iDumv0oZI7u5C6+V4nfxqAHid9T1RH7rHq100s40XXX8gWp+w0+lwJpLm
BK23GflupjL0iMkUwaShf5hnTHV9lkK7VKAAcGp/PsNAEdO372GcVsI6fLW1Xvoj
BseFgyDWHfiaf7Ss9SJJHd0qPyqEPVO3nygFx4/eTOgmUB+XY8TLOjK661XnBapm
+ffQdl8KDLKu9N8RlsOeJA0rt0bNHRPrJ1AuSqWt0d6putcaXmSBojs9fo79VcaJ
lje0gmji+zfAj/OUO2QRtqtJsYQuBKxGl0S5MnxbHYDB2Zo2SObbGA1PlpJqX6jf
xJL0jnmB0CKXzti/GECQcJJxbBmKSlkR/xY6koIDUeVwKbZk30cqlEYhh1fVQ0CB
joB0Jy3WeezO+hB0iCpJuFXoZZhgAkWCLBCjStNd95FB3ynkDFn4Fu5mdD9Saa0x
kljYRKY/LRUkNB9RnnPD+r/ygKGB/Bm3JVwFyStt3fNwRpyN9xy3H6IsZBwKN7VJ
X37fADXwrvAjo48oSJTa5ns9FT4oUbdotpqa9UUGvdr1MoQ7nW9ku0twF3RAF4+p
9P5oRKacQ46ttXcsKgE62yxV8k9J+4WtY1SAWAtB5zm9ZJbSoe1tFi4xaByAtUwu
KcEKT6IOksplH1Tq6QqPbbUIzSAZJd9Ao2l/WMgqinOrXCbsRWpXzB0isbTVd2o8
MAYZifwsMd3W2KvqgyEU8MvMYlurEPJapw8/SZahvjNc0v7QtGma7vSR/n2w/98U
5ABomy2+viQwA6UL3EoGohliI0wqHAk749C9UwXp0JRBcHUxctqKi7UBpHZTACqB
258zDYTNs+ZgpxIMFcX2KvtVGwTknj5HJILwEQMctB+t6JX4ZGlbZE1jPkvUqeam
z15sBz+tlHp4l0cvQdc9BJvds0BP1yfvIup6MARQ8ZvIoqSArPdcIfgIhnmnE0al
ku20ue9eHWslWNs53j9wum0RsOW/Tm2BGB7V66ng6IPf3CtX7mFnMr25OOIPcSqG
rJiXFq/oqBfgY5XXve9YKI1pJ0NuMAkQG1mns4DTITbaabZznYxCQSlHYZ4AXwFq
ybGDe2h4jjMWjvL0bThzj9nOOOo/umHcb+THgU9gciuadVZDb/AX3aFbDRMP0sbn
xb2L9GQHUzF4xkweEaal66jf9l513EecJrTuVVRijn1v1Ul3sq6BjW5Vt0JCXA4a
ITrNT61Q0JaISZxM11hPXsAl8r2a2R2ZpDFK6ciCuD+VqmNA/ueK7JsTal8pc5+d
vIze8uwktJcXfC/kXvIrgtGqSJTQLNFcIVvYDb+xEPE4yFCe7HYR9DFxWjSizr9M
j6Gv9Swg5l8MPsU5tQ0xN+7/cIdtpOBVx0cDr4Q33v+cN05mPNb9Xbdiy97OjtbF
lprsSdYgNvVc9agGSnd75USrYXP+yDUwWo9m/yB6zfu/FNvaqSoKrBdd6u9b/hlq
b7PD6s8Q688aeJ6KMbLH3RVfjVRZO4kKvFwoc94RNlrpOoznzR0nexK8Sxxy0c1d
gg0k6gqwVSWgKQjy3KmCnesvwo43NrMN3JYqIfZMptJK6wbjBX0sceuqCTJ4idjT
blJtpqrGraANI1RXXWc1il4Fh3DD/Sdv6VkQHjuREESkOMX7WjgigDYyvkd4jjG/
NsoZ/FwUd70hrMXu4eT3RGz/SMCXd0iwIsynqXo5hSOeS3CyEBjO5Q4DnrSxbPJP
bk4Lnl8KbbzMKxTEtV7MROUFZdK3hacLQfw8AAmSnXqLu0cCpiSo7Or94VK9qjD+
wEICrLUwVN8+63IXZIdArNwvLoFa6YzKik48gQclMT6QGTC3jYnfgVLmYQE4t3es
fOnlZIYhmfjDP67FapMGqmY4iT4u1OJYVzYQMj01caK4QzCNN71hs57HbqKsuRje
SLZ5h3BF+8//DjArCvklMpYbEWuILlh4f8WZjws4X6JTbjfUR3hHV5m9x2jt01m5
QsGe3uV76dpwDihvC0bQjuMSG/bAJpE2E2NpUafb0yW5HVvKTaskk+nf34ibsqzm
UREa4StZ8EUOWr7mTwz+3rs52ZCy5K7Y523rzEx7cOdDb5PQkxjgs+8aNZwxIm7i
j0myNV4kpa0olSQ+2/a4UDTXXNt65/DbwrxhPvZzGS0Bh9FCo86zQvvyKd0aICcS
QiMyN/RiXIyn/mYRXrbQyXKlR3O0JPQoU+QDqxqSnRU00eVeBE8HDDgeBgQkHEbW
N5YDvOqPvkIyjAlu1j4KpeNZTzwb0kedVVBUHVJDqttABoNey4V/h6g2sXhBgR7p
OsE73XqJfmwgWyzofvkRU8BXbZsNF7J2OyZmZJ2YjaX3bn/CiSp00iZGJxLpCEaz
r3ubZ/9GNP00DFxnLv3fMU4rzm+UnaxTG0qa5Isrca3NHxZa937kBZ4LbnDFV7fr
SwEpQHNtJVIvg+PHx+gaS2+CdPo6biAQFAeZPVOypKaW7meOvroIzM6rmApTgeUU
7/gtaXdBbtWyYEXejAMgTJwAfnD1bUxOG9wR1q/qsRwyvwRN0NiBLu/AkJUrdD5o
cJaRAyIy5v1oZkqpaMl3giZQepiYLQ7SOLC8hkmk1dhavuy2RwYpNAtm9Xtu5pD1
cEG1ZNRRxRgT/74g3AbZQzlXRnjLL7wuChGBjeBVQ8/1967ZTZu6dTe9/vI254DG
VsWBQYKC/KWxUmy4DXbYO2QClTmzF/+Utve3+DU2HW8xiKTswbs/efrq4E11Ie7t
DtBGTyLEtVk7Qeg4ANY/oe9U3nv8O6S7xl8W4kvdg2HERPbjR9uD6cAbgF1oVif3
hu149ukg3dCcOuMzftah0Xx+06tl0PYnXyq/r0HXXmIJV/eCRAX77jqUf2K+8xQv
IuHUkTXXpVfxdrCkvHC1PBxRS0GeNlXqRsua2ASIOAFoHFvN0CI2hhEJqhgbhuvW
/zq8li+Ar80wPPybA4iLng6kekwaJRzsYinkttCjAIK6cyygF40aW0aykrtGFg64
jeZtKFHn+phkzFAKBTNNMwWyV6usLTc/aimb3k43P16SUv36Rdbk2CgJprt4d6NN
B6qasEjpy8INPLKVyncz95D5Qc4BJk0INzJCIOt7nwLnTa+O//rdlQabpBlrPh73
niHu7iXRzPTLKDzrx7ohNi7YS/9djH+seOQRQwrw/c698zWdiNR9NVWQlW0Y70tq
qWy/N76buEixxKUWTHi31Gbr97xssFIq+dOpKq12k/vcxp3iaIkxnaTc1MsvuzNQ
IlkmQ0TJ+rou8F+ZJRrlwipkNiBgQPCdmSdHnSDtxoMBzMNQITceDtEiGIMUcRjk
Ygd7Qr9HGwSoZTklrAvQC+abIyTtheLHFZcsGqWh04Ne4nlJm+/huZ+MtTuxwdg+
/3qEo2Dy0finD9Ylsp6+3bHYBalQLOMww5YPMJdw3OrB4L75Yxj8PHhJm2qDh4iU
E1AeTFL4/1Z5VViaGylxVR50W1t+Nj5P7w6tibxRpxhJgWaIYeWGDXNsaXEIez1h
7RVH6hK1/bh2Daxy+PyfLCt72t+dN81qOj8omEfa7p//jDq5TqUr/MvNXM99a5vP
Ba7ImpvXf6T6vkzphrrzMApLGGx4xlyMPjYLdBSNewn8Z3/eSwQzXErYsa31OllY
EQjxMGwTcubTET0m9NM7TapUlCtQy/P9JCPfu3ZLZ+5ehAu5JS+3TAO4AhKYUYlc
J+738r7LO+L4zdDfpKKLSvixFQ6k+3/W51C7i59VzaNfUYfsSy03U3H8vBdknBFt
PJOc24LeA2IilC9/CGRLcnJJnSX/K9k22WvpITgHN03Td0NJ09tIWR/FjFWBfh0g
TvhIilWGfDrUpKjqDkM19suGYxZEz0lRqDmC7H0YBM5MWnP3cvJzV+ohz9RyOCKM
4ekq+tDhNFHxVCblv68d7VBmiINp/fky7ownW7nHTaePnsbmBovkKj/gyUY8/+Lr
NLJV9W28qVkzKUA3w5WuEuvWMDLrQIS34e29PFMG8AIEUR4VCsCPk794CYmcXuXS
F2Hq7Y58Sgs4IpVkR/9sjC/5BUxYHKL+BC+0ngqbDeXUmDcK84vYqdc6fNyYaY0J
OBemE751MsqmQnhw5OheMaQDtAhvTNLQU9aiSt9gnW/Al033pLycJdE1qa7xuT07
xEAaNljUrKjkT7qzbCmumv2r8Xe32Swu8/PTylkTRb9bn9y7JgneQfwnEjaNg6ce
OfUx6wDYMpZum6PukXlagRAhaphyrlWjKGHyqaI6PjitcYhDOTv0+8LIa/Rb7zaP
v3brnc3loUKOmUv7KdYIq7q95g1oX05WYvyZiLmXzNt0bPMl9s5YoRXgu3Zrx0S5
D0Xipy3Zcuce81wzgzElDmMD6tQAcr/TuMSnVEF4ZtofQ8UUemGrZJvt3ID0seW+
AJs89lLNslBkdiY/jVPlXppk5JR4rXqEsNvnX6QeuGA0ITp6cWQKPU2lcm5Iavtb
vGzzh3BaMNO1XrY+Wmu14vUVSM1akStDPdAImIktW3WUbQIMX1svkQEI+C6tgK8T
KtUTmmuuyHNmfM89AaIIe+zbNIVQrOTcw0h8x9sdkfYv3LEKuSs6CoF2m/B1Khg6
IRVBP5cFQHeCa5CEanOgsPBd7IwXjpRq+1CF39WHOxmIS0Rrsb3hog90o7IAuubM
II19uPCOnAvPzqZEBuyoa0nCT+yotWdJRoQivN8+WyAaJDa+MJhydbM7OFZ/jNNx
ahHqpqgWReoKjmgKr3Udbien2CcRBBkKv23Bw2QHclJWBI9Gq2ndzyriNMWepNMV
CSah6ucP/Y2Cd1zQhMjTlSuA+DGf4EFVEPoeLidoYu3iTH+3b+zO2fy7wBAZD8XY
axRnmhS25K4zM6uuor19c0/Ls+qtFjHedLICb7gJObvRBX7T/FGJ3kjRz24sEchR
uanj4VuWkpVTtuvmgJXXhXbBj5bYkQ0x3wGj/L7F1MuhrMpWxP42yLF6z/OJGsrm
IUCO8yrrj419bCZbAlNdHZ+Eda5k/uLXZlK0orJXdoDfljujx8jhogrEatl/XYkv
FdwqWSutNTe1dS7vhgrR/Kglk/LQ4kI7vCnFjDBRI0x5YgEghTxHpdengXGMwxHt
IwfF073FOgivJQW1Haj4VoqFjnw/y7RjLvbHOk9CG2Usf+W+dqxOj9F+E69BFzXM
C8PeucTTkL+cs5tK6jFqHi46ek08e98nuvWsfxpN26smSFeqT6khYm1NuHZ7jdFh
oHaon5bzmhRmwriA9aV/ZrxDEaihMEhT0dqgx//T/1oo5HqH2ei3t/vO/lq9e4Xe
VWbXqWrcyvu2SVjtQwaoKjKHs/pYTf2CscH3P4g9Q6rD0eJQdzTS5qJwxnmFyO+N
tu7A8uM+gfGdVEWQCSDIsJRLCicsNVqwGUAkM+H0Szg05f5/J+Sy0nbL0T2WTSoO
+CS69aspVS9bPjxLu/2ByvKNmphgSuKGXcOH5BNEiLsSvTLu1gYDGPQ73vTp7cRR
QPkChZylOj6c/FBaphLFDQr4XOwNZ+kreI6zPpyMTHt7PwspxRspnSNUNVCAitEv
bhHiZIao0YAe3QBVgvezmzXL3r5haTyIeUcVFtpJfc7jPPhc6tT5AO5R5+ekcura
1ZaLpJi0L5cLa4BdvGbx2y4EkqUDyD5tW0JS++lNZnXlmdAzXrI5SDWrVuO/n96o
1gJJrUW8ucuOxUxDy2GnE1SeOczchnzaqDZ1iwqJys6COyYrQX7lGYSeaSFpNGw7
WVJbBLnk7vBrgyG+LpMbCnzSbHf+FeDRTzOBxy22FsyUWSWbPzVPUWav59MtQgmU
WF18jhpq4FVn/aes0x01RJvFHFbikOJPo8EcC9y0moyCFAlhTIyQ5fzd9Ax4P0B/
XIqzXormIeRFVElSAw9RQ26yKE/DqTFxVBXGwQO4RIqnzx2yN5tlgNFL83iDMVeu
FQcBbuziuwHqUlNr1kBl6IM8hAEVpbLvEa77i+1Oj60JLYEZ+GFIz8jIWcR8YSXB
TGZosno6s9eQLPcD8P3FfzeFHFG9qRhE7ZtHkEle+JQ4yL7LAcs6M6Klyqfnpf/d
oWvccVs7ebTr2xyWwGt3pBn6y6t39j/PheTTORHhII/ZM8EaH5DVPcnlVR3V239O
hoAjUzEONUGbgaokip4abTVk/QQlflC2UJBloLng+pmXZSi25xsCv32GpWTWEiTQ
5pYcDOEkVmDs8teGPkah0si1xsaejwEHBA9Q+7TIi/J0yw+USpbNCYAtZw9lBfho
rLx/1G1MFElkQL5Da6lhhwTrfyiz2R4fbRyY/5hyw3pCDgqTysPBLz9nMD4rt9hN
kX3Ypvoy4ZU/mKhlh4qdRZTd49SFbulntwFw1tJzcciG6LAGBy/wD+qvST+OyDam
B//ZqFZwLCn/d+A+HhSeKgvpTDivj68yfsJVz2R5xoDYXvU1tgDlBI/FrY0OpAux
yZAKMtfG14iNaZ0/GBMxaULHuQ5uGZZCI+MA231siJMc7LOHT3mr3CG5LMlqtyT2
UMeqzUPl8VAugLfdafjMkETHssOGzSJoNSr3BWXt4V0vTMQlr7fngOv+rWMb0diu
rgAUjPL214Lfd+8SbZ2AMiWyK/wyBFXrxxk6Vc25mnLIiWFKbSD++v21icGsdVfa
t8nIQfc3UU68V1qzJZIazGKOjy9atL/yWt8bqed+biNFNajVFQqlI8LmMGLv1Whn
dALjWT/4jraYEDsRlEfntthRZQomqCK/EWaymPzZDHGbOvLQPp8Y/dc3+ytv5nAw
QMuvH2YrhGAMsVzxsTtnmjBOXv388VKmiXEj3BH+ARXoY8zbnPESS4/VR1k3jO9j
pZykZfeyUy0eozhkGDdW4pYGP3aWw9Rw0mKMHsPLjNuRAhoPRI8i9nhwGyf83X9W
oHs7ZY9KrfkApNa0s1Av7RStrFj08u9F6t+keS8ZaNpLy88hJFseBSZGPvztUqg/
vOs/pkCOYQsJGppch8hXa0pzqKhCjNd68Ysbk2q5ul6RqjLMxUBlmlYEq3EL74Du
VT17dXjp6EkmOHWppCedBHxI9BRR5jqTFjs3luPeyoPYqUw5/QwKc37dEfViN0yc
FXD6c5EXcmzR7LR5PC8n5SpxXsCsNEisb07mroqcRPmc/I59HIWizgm+XDqf4RB8
HKdeTsRrjlePJnBIPfqSkycAhgl0UWlpl8+5qeu2PXVbw2rDnEqmyNw8fZm3Iu5I
HfiEm6vC/sOmjDyc0yZruS68oNVjsHpAC9C2jONyEYaiVWmlcaKOd6D6J6mjNNsK
cuE3MqkRaUSaZTDd66za3Dtl8zZuJ5RqPZGDAby8d/kyOjJ5mGc6apOcPAzTVATF
TZ2us8dQG1tUwZuTbZjYyIHJnBmwL6TNxaXv4yaKqiP7xCJ/4Jshmtt95CvRW6ay
nqbBFrQAwWlzchJzrXOwseCNi86NKQcfLnxNWZ8WCIfpv7zH1z9GYz5AY2LFCnth
Qg0UdK1JrXM6DlLRuOvBDRSv3klBumiU7LBq7jo9XTR0fq6J5e74p4fppAxgVTjZ
kCELi4DVvThYXODcgsSIFV4lzrLV/Rvlv/gWhZ1rXpxKj73MQ9t/qVxGI05yiDUD
PhMBVeK4LLLjlsY2AfWTnhdqUElkcsyseIho/iMxPY0bq7tUf1+EsG7GfdGlvR7B
TmIRkb7uJDwfTXR3Coy6zgLAAshhfXzZt/7uIRQMUVtTU6aJcJVbmDQOAvsk5Q9X
NHHDTQolMSUg8fC7QOXPXtF/qhNWf12ytAj8Cucw3zGBSsqx2HHArh2XoJBa73yZ
JcJp883fML8A8BzKpPJKQdn5EVYpCdj5zZ/W0oNZXsS4xuFniC0393KlnidZCFqM
CL3oD8Am/zFVHru83u+3qXx60GLJCV9CHTYjuO0jFhpC5XDaqhHVvBJ/DAZL4OG5
EV+YsJC+vMDpButkNYXhhHUKJDDWJggJCyqcGqmvenayjY+jcrdaNO91tAI8xKoY
NoQhCcKFDq/yqWDdxg/zbx958S22FESMvcWinhLJplAmGegulwqU25JalixcMJqg
FTuiy6dlYjiro0ar9iZcGW+HJxMQ9bb1SnCZ8WOTx5quyh2MhHwZ8BZ3Ua5XhXso
acFOjXwbT54JnmNbs4oLHNJ3ovtOrHZ1zAfQpLtYHiMHPAGDinVuvuq1bJacmFYW
toENQG7cAibTjNMRzL7oodB33tNTzfaPJbO4KURFx7LMH6Orz+onYYy7f5BbP6eA
VeY+bpdNqN04x9OY7wksEbJrUHx00Uou5afrg8RHqZYcfDPpDY9j62qdlU7FwPZn
zCxvIx+s1FOeF5BQ+6Ed/EVAd4xyJY+vM8MUQ0IU+63nwZOcgAJ4E/JkQxomFt7y
mNuVqseg+H36+OYFdw3W66xSeErqrqHOQoZ+yjtx624rEEFLoOZGG29WwnB9cevK
McOym4NyEX9S1bayMHTEGc9GxEhle54zFb4AImQGLvkxmGHPKydORyaf9aMuSX4V
E0jttH6twKZd2dYzBvc+RAlqjn9xAsaeI5eGqGJErVHRIEO7ekxNcV8Ir/bXyhhd
PEMOvWteGTdCYTR/e0dcu++CijNA+0gZqVVqa2pZDLGUPV/3lXqraAN1FD+4cjoj
BuxMrRtdDDMXiv/i1NcYy8zptzuPTZPzynDh0dYfVfbQfeogKd7JclPJeSHwq80F
soMv6vQLNmXaOdpqoA8Daa7mD7OTM100O/p/z/SNHJ6KQd1PV0lygj8KR5d74nDu
0fvsj7BrJAJIVXvlgloAF/EZZzbKuo60ZlnIeRFsCMCj2g2xwDisOuKkra0GCISm
/RSH91Bn0WwGmh0SADjmPX+AUvb2YK6EFLmm5pmWmw5qg61xem3Vs+2cl1Tn/EC4
HO0+YU2yZUFOlAX7LmpxRPRMo6PuPKyHU3msZPkgQVqgyTKRYqZBjvfI5z4JWiik
p8WHnBygebMXDMzjwvIUZ2kicpU7cNMWkfFPDkh2ObyIyVdptkITsashgAFgEvAX
tWyQXAzwi46dEGXAUmuICiagzq4EtjdjglITxKJHUFQK7L8U2FlrGR3YFheHEXSb
2Xti9DP8QwQz/7rV7Sk9TGlu1bBWguP55zUJvdTbd5WOZAKGb746GQCB94QQ83/k
esnoQR4Rd5uighOFks1cmGxWsEQrdrtBqszvv6J7MtLjHVLzap3np7dcMftjOuX4
81zpL3CqqB2caSJLC56tPEw0uSPdvyxGmhL/zBiX54FkTYjQGp9PwaJZrv7Nx/Dt
LXnAjqZAvD8oTKxQh0ARjLcwzVOXzmqIrsqAlYUzaXvZkBn4f3vNJbFanpP3RdEC
N/pa4qwIh96jWZCzmyjhxvdk7VjqGgLzB/+3BFXdRJGbu4JxjcrmeB14Lh/XIHiE
0tyUlOh6kXtKrOFxYEYBPZvWWgX90rmie5rYdcXIUAW2OiDOfN3heMw8ZvlOpKwF
xCHfoJavNaNuStWe6iZhidrY33lLZqtBo9yIYq9nNNc0Zgozj0A6qiBagv5oHvTl
srojA6sqSdJ6IsXR1t2/FQevllEtsO+oJvIBudmPX+koc2y2lfgIpHgT5R16BqS5
yb9dGpLXukNTDygon9ESrPz2HUShDkiW3XUeFGx0AtH9k5piJLaqNdJGNMKPFz1r
Yh9+gD/infxrinicF84bKQsYSZ0AJuo5Pqs5R1uIRu4n2W4g+QplduceXXhmWotx
ZNusflatnVR+QYGFWAUEfnv3ZhvM/U1oS4m6PmCbczERnMOhRSESZwR/UeSTg6ru
Pv5ZN8QBnBAK7ZZC8RriCcypCe7VQnm293L1bLbrsJPGCSblBrRduptXC4z6riB5
UT298W/Gp1zX24DfUhCOketMo8L5xsqyU0aT6ueg5NS/05lMTKxSULXVeypIBSXP
ipN30ypB9HAB5BdgReg6fmxJ3jallBleo80Hqb7tEe04y3vTVQWtCtVX18vOr3Ql
miQGQvrvKIhPSio0RY2vNlaw0orlMgxZ34k8Ojt5wBtc9NA2CnbFdiCeraGre26h
RFgBCMSH52qPMwDqhpWSb1wXNF/uvEFvZWK9xeG0GCdIZBoMILQVqbOuNBYEq3TB
6z/iDrTKpP7o6ZvQZy6Cd048hQ1DEZ9bQcxvWnUJcsnBtggU1P1aR2zrA6mATwkk
S/9O9nKReVMnyHYXFPxtle0/GY2cJc+xv/H+hOAWif1HO4GoEbKuC6Ci0KoqqL6I
0TdwPafaQzpohTxW+AkQlg5qLLoxqf+L0inrmPq8wdcJZnQuIXfdWYVIuZqm0oNx
E3vECoqNlh1eka1XxXeNTgFt6tvGDGfOu+3wA38VPDllWLPzzCMjG7hXWoyunu0z
FPEgGUqeYezF16RKm1czIqrQ0bhabtlfzair0hBhrlCGEy6yvMwwQxNz6kSsEWmJ
O9HKVZ85mQEhbFxUpz3nmPFEq99q6vnfm/cKoCCCl09fXqzxiMqUisrR5ED4Ds/f
9WrBTFU3803S4ZrpPqZXSsmhqxqod2FMNSliI7oR04KyR2morespZsM573rd+EME
C/AUBuqhgpVfsabMM1PjvX/XGGwXklRbCYXM85NjmQw5IggpNCW7VZsoITLwo4D3
Eolx7r6jCqSQCyY0QmQsm3O+dskk0kFNcWTpKTQPvdA2SRzVK1f1+kI4BL2CVFLr
BWpz0jK9MjbG9iLZySex0OwMHLx9wjmYFzSqmV3deNexzpTdWArzrd3zfbERhKkG
G8KckgkZejLo9L0k54Gh5JGkM/3DR/H5EJ8uAs+TcyVqaZIAGWnr6vpq5bQl5KLP
bLnLvo4hQpdwlCqdUu/mlidXEbeEKPSUiORqXJf8tGBAc4ouob2vL3fb/4wPkSB+
+/VQMO1QCYg/pSmkXtFSEKzG87tCxUrdb649X1fWKN1uGWp8kF0RX5zcY48rKvIv
XbCYq7eg5MpZXSpus8FlRjYY1wcA4X658OASw7NjyAsAWdi1+xL2/SCrXitKaAfs
xrJSyH84qQ7DkFN49O5vt83AUOwybaHgcaFyWtLMnhVzIrOL/nXvvASM4INt2Oyj
Uvq+iegentypLROnhrO9WXpwoOhjpeKDMbhny2zeDD4S3lckKvbbgjrK3dZEEQMY
1T2JWiC69OnPdsWNMNnI5vuNnddVfv0u5dbUmxck05cls0BfPLfMwalYQRaNO+o0
wVEhV/JsnCVkhiQfgu/l2RVN2yCchfuQZ0/i0GRERbWMqC7skW61d/w5qQzNwZUY
vEsy/1g7iWWlRg5O/F5xruGKMeyafnnAhZKBSKlyKKaYy/JpZX3h1EEUQC+GqW7k
zmegjvvcQ/xhe0IKhN7gdINqGd9JTHeyCKCCNaOFtl5JFD0DyYUSSuobAdhLhiwr
dVBM5sH5jfidceSq7K7ht17YjBRnx6SQkD4VQLh6RwHrk+5XhZVklJbOqcvNexR7
3wcAlIY4D/G2/B+w98SOqenureMiCVrbDIF07S/ZoPZiwen+pz/uDBK2ccpTrdHE
Uuez2otQQ+jnr4rBNptIf6Chp/5jnY1i3I5q/F/x25mgh3GkD3GO5Bevh8ABqTJy
9DYullc81GIiIX33dgEnV4+qNaJCRbkefFkiw+hG/HtV5tP1K34Rfv8FUXcElTq+
fe5WncxFZGGT2GcPjGIXNVQ5Za4quZl4MWdykeLw3Z6H9uI/OBxmvphd1cbV6YLL
FRdyHTvYzZAYNFma2IfaecLfN6/yzyVF8dPDUVfZVgw8wriaxrPzRDWKI18HMDz4
2wdbJFv4hjSJ4g6iRMwU+QGDkeN+4WzZmC2xD6N3LBINssilJhd1UnVxJd34YX0j
LiP+Mz3wmD9/X935aUFDbSgMlXzfOhYhkslY0+ohQsuzI4YV9Ms2L8WLofOA3pjq
toQ3TgfJyUkfklWBoD63CM0UbxVHSA6gT3PZnl3vNXf9tXcj//Zhve+07DoE5oZX
DpEcnYCfvnUMCJXazcExiKmXyvZwg3BdCCf+UolVwnwb03qtIZam6IFn1fwMjv7+
xx9l95EKxwCna/P1Fy6lEuwYk19eGBn2ApbuHUf1XNRZlKG+tNtsbzL7oFyannn2
epChCOhxwOOuM0z5uRvPJFEMEFdW15x+VYRO9wXbf+W0VzOtPmEVtqM8YWGN/xkg
94p3eJ/dS+dCuC9DiMJ3TNPKoBAMLFyhjTRvuMN2eRs15HgTr4CIW22FLKQFt80T
ccmMU7VWWJIprBTUANfDZ7b0HS8pBiEBfcKIvwiaNMGrtoXySbWg0PBB+NN037el
9bKmAAWvbpc1rt04TCpkldEUViYaUqEIagjJJ0oi0f/eUsQ8uul0s9jd6dkU2/e3
P68xH6OzaekHK+6d21ufn7WGPBCobZVORl/n7bUmnQRaJx/dWW/ve5+6MA+65tOT
tg6QWdrSkOZYKYnS8E4TQiRvVvxkqUB4J6coD0scZENRCOzs5ya/NSwJgreUOTZI
QFzDw8RM1FbpTWgrq+K2lt7xlmvBa7sbE7RMxNKw6u8QUYeMMjiW+geOsVm6fHJP
azNS9SqrRUhcHq/+T/utgUi5PmxnKuabqy3IxmVX82t02Ns+apIGXZJmq48fpEZg
Oa8KYvfyxEN7A76gQputm0RdgCiAzUH/kHSvolWdGlxSS+NXrcKkjOogTOrNvOt6
7dnA6+VMkK6VbzIYuhZs6HZeRrEJJjPqi06cBXl92xblJk41rC77Ooppuk4PRO4A
lukyBmRteP5hyx15t3GO3S6YnxITtnT+GGqwoQzAldIOxIh8BEqYc3gtOrj2Qi9B
xod47UC8m+VNo+Y0SgwL/O6mj+uU6q3N18L+xIbkmVyy1IRtvsT6oXeKbGQoJi1W
ohOvF4hVTHxKATXMw9hqXdvld0mXhsHp7cmmeRHQKBcGGDYH9LU1DLRFaNQapd3B
nb9xSj04Bb/qoGXiH6MBCPq8ogC+xpV7SaqJevApe9kG+fkFYRautO0VrEit04+u
Bw1r0qtXIk5N/OZjhJFFNYeBVC1AWRkaoA4JLFpGQ4mxKLLNQDxh1y7MvfRYp8Fk
NhrNfm3Qx9mTszqVo2hX4QZ6yraEFJxYsFylqv9zMjU5wdX6Gu8JFO5i56FQB0Cm
tqRehqAnqJFuvLvXBk3Cs13bt63ZzES0EU5+aifCLBTtat+Mu6cIQDUJZLh/XvRo
ONgxZLL+aM6f+dSXRjZ/t8jM6XU53YBGapt3XkIal/iRTbA5asFQVS0XVe8Bg44/
OJjGcERHGuQ9xjr+P2N5WSn0HnmVvGheBnph5qdlepu15iormF/vgoe0fuDtd/qU
r89k6Xl1ArvmWi08a7ZIpCJuXU3hd5uA0Kg66RPrP2zZXD6aLzfoSn59oYYboQ8h
wu6cf2jEspkW5GU5o6kTGyHXaFlea2OWlYIoOSSd23SilraA0ur9c6WROwFj2OAU
1EU/jhqHfLhfzu8WftQG2zMIYRlzI2bx3/7DWAkS4J1Oq+B015heBAVvoNjS818p
Rm9qXmBGuJfe5UFlxz4EOlvJlV/3OQpZmZxCcJVfVE/lLRMCAgrzozfKIKM0FFPk
2KmvkDd12kFG94sitd2ctELdEbnw3MbFfWU4Pa33ZFka5FinCgpgmWdLxlMTVtK6
IQNjwveg9SjvrJgYBwadIjNJJIZvU0D1cVenEUTFqQBtYnynJDOWE7+KI4vMalRn
c6UbH3jwa0XbIx1NQrr/P0O3vAjY0Us7tNeIGUQO5eUMc9Yy/UJvasuov7lbko8g
c9kx3wb+kkx2hL4jaJcLMruKUUvIxEWyoM8fXCkstH51dFcTSDX0aWzYNCWFCicq
tpZFjjjVnxFWBZc9wk/ajYrpbleuNJFzLpSRNZAqL2EOEJDoJEUS+VNL7YdbXsP5
+DFf3FMh+RaQQP9gC+8BzV8m5Euc41ZUN3eK+Qm4fLJrv24OCzdlKVD/UvfaJciZ
SAlE340E5ZitK6u6Vw2RmSZ108kvKgo7+x4mmOB1lQQe/aUQYyEIipf31jsHtQK0
6ynKFeSMGlu8TiY/6HgTZnbxy+rSzp2W7B9b8X0NFiopTkXB2MF5lI4tHw6uMd7c
Xv8FcI3QP+0W0fyiokqqRVOxzZmPldpQsIjYN6z1pBkMpJyXP+Qse3LSULeXqVrQ
8UOCiacPbNYd6DzhplKU/A9Nv5DKC7ymJONMFlrFflDJy6dz7P/EznsCffOaJ7w0
v2h69VVA4UpXoCdLtrqkgxK7VirzM9a8sfXCOsdGgdgajhKl/D4KyXUOqGSuxus2
fznZhX1TAxZ4wvWZFXwB5qzuPu8CAq/I/Bf8rUAtXbx6+30nw2NNYFVMHV9C2DxL
BPNndS1Dxgy9F+WvC3pkFIFic/rPft6xSaqcpug4L8PfI+nKFgboAXWBXOPnJM3c
qA25GwVbUCgW8EXjusrY8cnxOEONgByXQpmgqJ5jynSk54C12EOY2GCJc3xw1+4z
V5tzi3COXEngc+ENMi/gR7pKCRG799JcZVVfcqWKVndGxQI/As/GRAVQGh6ShZbl
TxOXMMwsSqlTg18U0WqXRN0JBj2OTVBJxVfImlt2HzqEAhcqtKJXw6bnSXAJza8U
ht1RJEY/tORgRzu/bHuvZ7n73XWw6fnQ9tvqttkyRyZK1v7qrXEmwxr41OO6nJbN
hO+slrGgGS8KJ9dLzIlunA5+5g2cnDChupv8vY6oKWpgJpvBV9FC2zgIuVlQpxYR
MMaT293qI/iV1Ne9MLQWYJyiDA/Xag3rulmfGjqpn/PFjig+xIPD1L/ulAGIs3Rz
JJpe7xVRiGFJDWi85s/QiDRARsxeApKHO3tG8DG/j7dL+xGxGarwSeMzX5+Q0agj
M9RSs8v3dWrvqpHLwtV0YPvEQWfPh1E9WeAn70eq9E0yRsz9ptqVM6YSNWlTJt+p
NQCqvQvU9jaRPEloTtQYH22nMTSkwvkVo8/s5CRwvYytQ0+qI2cvgS1jHpbh9uQN
Ga+qTk1Gx7fyEqjxfQ250Ib76D9xui3Ro1iCM2P95daCLIE+/uCyIisF0tct25yk
vXRSWEKPquS3upCmcHObVXMN1IgbrRKZ1+1/eh9FsY1Dg7ozkAzFqbmp/SP6VH+W
M9r5usWjksQgUn6QpJOlbDc5BvVJ3baBLQuYOrAF+2aT6ta+PCRq4et53CJIMHUN
1iJ/vgxa0BgKf/R59esJM7l4hdyRPg4ZTG5q0+fZL1p645w1L71cR8J1aIt75UQi
H5g6JEYlGnTZqzIjgWk66xdKGSNaIr01r3brF8meegrWgdy+NzWvE1Oxexw+8SP3
33sFZKJkwpZD0wZo0YpEdtfp2VfPT87qg8aGgyB2ANMZo474baSMiZGeUuYK+T6S
96iUqjy7P/nfW+76ZyDPybIyNtol/UWOIb46bdld/HsXdIOKVkRdRHjhL0F0VhPX
X3qi4mXzLr/Mbc4rtLmAFnL2Kphq7d3vc99aIvjRTaUTY4XNn8DU1FmfVDBQRJ/O
sis6XWQb63DfHvDsTnRaxK8RN//4zABXQgm5sBYyUBj7qSO0mKXNvV+GI83+RSYB
2RtybDiE6Wo9k3Ctuy6ZV9wtXbR0RbAxxwBKChMlG3Gz8T+QAUimNm8TCow5EnyY
QY/PSRv6QKrfRqPRuJa2DCpke1t6uPgzIEw8OmCd5+x/fpRp/d7XPHQJqsm0qF5c
9LN8PzCkq9arXLgVMK0/jz2jCgCVaBtQ6QW8G/A9hq/Nz1Lwrw9LhQRZtp+Z9SmM
aa20YHfbwfqZVgFQqoY2e8jtwNtIRWEPV7flW/XnWyQGsWG+2Xt9gNNoOytnnoKD
Ne7UlxPglS5bewIzgYI7aBXJD4DAYf9MlxP9iavAQq1/IPdYA4CSlOqIDXnlT/zw
mS3B7CDKjoMoo7DyF9+dHaZ9Ke+FsCd/SVdeJ1ZVaxvwcfofOVDRAPkJh2vfXxP9
KbtYr+zaLxNc9pEJ+DOS+sNSuPFnbH+apzuJBfMPTP/Z+trNVVnziI0zuIBwK7fn
CCj1ux1PXVgjq23BxkGWrohZn2gaIFWhL/843SzTNb/x8G+LMC6MV42I/vJ8kjhO
Q/5MUJ+JXCSEjHB/lJP0TDArD+dGuXodBG3OmRfNfnydW2WTVGlDeaQ4b+l4F9oV
r3La1YKxTEKg60/Y6rWixPgiehMYSlSg/Y8XI9nrX/EwBkJzVutFVgZxvHMTxVCn
uFWsG6zTUbeoVj7M3n0jj2aTe3L4NwMloyJoauP5NiYbUMpir9EJwGFj7YcsUr2i
f3QerYAovzXX7NqAsvIL1/YIVArABg51Ujw9QYO8sq/alIZ1t0bIDTKpaCd3VX9S
QX0pJzA0w+UrTmigmXGToAZPoerkQRf1aEn0o3AwfsTGD9N1Tc3x6aNqoQ48Px4x
DQsb7hSyqUjgaFTmckJRveTOrltY6+R5t+UOtPIdohnpAytGvl1dtX2I5r/u1pVQ
mwM66g4MQgq5C0c8aZ8fRicuWf3y2+E5SbQo/4RBieRySaZGZ1e4Bs5UZJzR5P+d
dIaH3VEzbJj8Xk7yOyQyyagEklFYqX6Ic4Fr7v9qL2JwqtG1YWj/XciYjUE2ODzT
xW+VoV8AlDHLheyX59PCOkbFVLlnX2YhfJgIZnMsKT0MKPeGHIUG1Xmm6KHGIZHC
hAQBcZPxniZnHQRweml4yldhlYIwyBsqtvDpZVyBnBlCCvhtWhNzvLHCUEB88jFT
V7DS2Din3brRQjCgJNhjGNpCAQUDL4ptB7hLT2gMlSfA/mk+pqqr6h1p6e9mDMPY
ugopQ5eTA+9aGr5ZL5pENA6C/rOKtz2xsrEZmXrdJ52Klprsbn4B3Fy5+ldnU0ot
nqhHj6DV5pKuyD8jMQ+NWG7NrNdky64srOo7g3JMd8ZZxXw9V14CluhzLgGrftea
3cBl8MHocPKMO0yccYw3wcKkYoLwA2m6eqwMuDHZUb48ArneJzpLKDvvgRrKQELl
TnqaLDghuFVadykuaiO7IcFfVPrXw2KAekyocJQ45HgAkFf47fl64iZG2k2Kq/nv
4GtD6wXoEluzBTrmwRwo/rkX+URecubktP8wsKJ0aX5LSqZdOslgKJzd7WFvbMec
eJ0KinkEoANe06irB+IHJuI9CseFmaVv8EKkpvJi9/0lm+AXPyiPzc7W/gWN1gqS
kIZPZpSmIIMgFw3bBmsAYXo7BlSB/YNbOwYUJz9MLtYT88BXx3EVLJe3IhIxRTJb
u4KUqnqUsT52jdapSLldIxW6i5NwN0w4UiZMoHO88pC0YTx33tzctHb66YEYxqSw
ljSM4lrIOzI6/G7SEqfHb8DZ5t6lqc+54QT7Ezf2ozd2ecbL7e9ChjNy1NO3rA9J
2nrCgWJ1MS5xT/4S+291qou9sw50/TiauoUAp/0NygvRAjhnXak4aIG/CDn/duX0
BqInjqvUAQzy2a/RxOzUF8o//3Op0iOj8fkLNZy/yDNDmMoEZWlDV9qBaKvS54BN
Y2yrDAqKLlH4BPSP2V2JPzZrmfwQjImdL8YVYpWkkcHup1Qqaxdet9uW10K451M7
AfAcWb+wKsP7xgHF0CAkzUsuIc0k+I2WcUqUrCKqARbXmyRFqVUGcBxN4QvrfpGq
+SyMVgDJ5WGEQZBuwN90RAEfVuM0kMxoKdD5zxoJPDviMPl6xZdo1DgpDHDnvPVc
IFZeetDYB6CVB9Ve/+z0oyFDdlvi+UspzsFGJngX7m3TXuu2wkaiy7nxUqgQJmLe
piH1mlCjUNAO2/i18SDopGb2tKNn4bguN7IyJpR2I2GJqjaIdxRMgU6D6UAMJqJp
z+pedD6Tf95tdcg+LGcFnMaY1/jjDSaOyDLpcwYfeCU2ZwSE8lf/OqQfFYunE5Js
coD1stFYSodQMalFqeOOr7LXXvWO0nbQj/a5GJw+uIoiGXPl5h1OgHmMjtbOKiu9
c//UXGGycWs0dpKL7fKbtLS+IRM5b6qMAvUyamu+dmcuzvQr4RO/bq4d0VRSUacF
O9c0ww9lLUBiwcQKAtp+qznuhXoeOU4r+LaMakGPo4W6fMLUhpdIquCQKpjj0YSS
3DHb/E+RTE0I7FHnT5SPXyn4SfkZ/JftkcyYvqiSluFbQjJ8YGA+l4b6Swyanuyv
1pArgBG6LNSCqUFkFI9vUn6Yj8safsjMXIk4AOshEMTZlcECBedEg9BgPkIknbzp
vMNGpkpRdtKwbnU56UbVWAN9ZAeAQqis5kW5m7jqF6aSPu5sK1MEMulrXbzJditW
PsDbhzOrNOSEVxYCsJbfx6SXTY+JyocZORSiyS94QkwFA4PbmbpGLnPrY1bI1aZ3
UJwnSee6oTbSaIEQ3CpTNmBi1PdJaWKYWoX80hdHtnL8SnYdt5KopA8DypkRHSkS
wEjzMuspUAGN67tdqEc3WDW1/9FqS3mruFMLihThR3HWRSlpLvVkWsy1QmsVsl6/
eTdgV1/BNWITGPZ+NPsrXkzPnK7WVlFhz8NaezCkwuIXRyiV67sfLuqjUAbK0v/w
xAWCj8Ky6/A9QMWqbnTyM5Z7JV31Qkv1JwVHbksQXZKa7RJplaNEIcVi6AIo5zmV
9/upL46KHTj5GD/iZgHEA6nDK7CI2mvX2c0viG2n7DhJqyz7KKexqrqMNOZyT72Z
5E8+y2ZJMYMgkHRIt6Y6jM2H9rlbbgYShBJMnbLxSmDxH/qP/bGPhooBDXuBRj9y
dFfg97AmIA1bWm3guULUECCruXW+GVl5jNqoPrSbJ4ofDb1hFbH13tEEogPdbkKw
o6Aj0mZjZckrqFTSs2cT5vosgKzr8f1Jb1tGoN8Hh57SPwexvw90avfxQjDQ2Jnk
NsBaRCy2WoOHHEwf9E2qE0DFbZlaf+XpxmrUuXnAsS5K8JjUifCSRZb+bFWFQfaq
1xhHHrsoPu6xY4DCQyulYV7Cq+5imO76K9ZBezHy7HgmfcXF23Gxo4ndO/ll90M3
5bJt5GdKdK3ofMG5nmNbpC+LCEg8GOlRFBF+EyOhFYYcntsCQanZu9zQ2kkQt7KY
OOI74jBJkyTejdu0stbMw8mznmCDkX/R5MGR7I1JlPcZZoCmqisYZgY9OAH+p0/l
2CHCa0y6fdZIXwRciG403fonUjZQa4xG5rUL+F/3iCWhdV7vswBbxoZa1LcQ6kUd
O1Sk/qOM1pJcyQ1oQAG2qYp3qYE9YlZHX47+tZhPySJ3CawzNBjW8DX8iJsFdtkB
Fml77VmPKC6f5HgL8LY1hA/p3gq0RmgDb/sV4jTPg5jRVD/5W9yszKyfsK0C8dgm
T5GB3/SPS1xvOYAcQSxk9Z//7QjpRHfWKjaMFc6WC7epUvWbkwAcWKcACRoH6dD/
i1KeBGa/7MLoXukOjCb2jxLrweecKi2o9M1zqQr1mBtOElbnDRqg+DzUJVtpsH6p
8+TM+e6QBA1Ze6WyhRKRwUxzz4MD+6nCYzkXPY1agYa9SnqFpHuIEjmSfYeFkBcR
Ze8e9GpB0aCaJ6RgPFZyA3jdDYL0xqbFNAqrA4OnwmCB/t9pxywvV2QX/DcrW4Cn
tjELF5wO1URVEgvxR6P0URpVEqW0YmNVeF6bvny3dTSEgvJl4qFdH5vrkZSq57Jv
c3tcnnaDyXOZh0o3+GNRL4zkYuoqS+FzNN7R7u7HPR8tVqgkE6IoT/IeHrwWe+fh
+0Iny4s1b1bt1VO686YNNTRPKk5TNLc5XNYktHwIjHg92geByR5d6OXTvdvmzkUu
NL4QMyh6/7HHcxlDdW3+k0Aqj7wyw5FCTq6qn6H9pgvUDDM3Q7pHcToiNYibC1vw
x0ub9qD3AztkPCQqRVO2DEF3VUeGfdK2/qWWDCjZn2Bk8wdGUe/v/e5suouBTqvQ
ucigtfJ/B3oOpWOFZHb0jAQT0p1L6px9zKH2gYblvW9S2eu85gKPQ/+w7aJGF/qW
BUKqmm40Iepzh2RxcweH3c9FbEWR91WKskVuFBF00OMuwvpz64t+fYwk0nwivgHV
LxadQqL93qS7W+plisme+b1NTLMiI+xUctT3OOarD7M7j7Ebq/LEyHxAQeCCl3z7
j2Rcq31BAwq8sQ37FaeqFYL18xCVga/+AYGSuCIESq/JSIGgIOnki2+i4PXE7SNW
TYollJIwGQBeD9utIg2X4q5clx9AiIKsNbKxWW3LR6vdDhrEpU4lFuNkm8DToDyj
aMyhyjBBdoiY9nZzHkusg85yTBAC3Zl5d8c7d6Oi09iVRFyZGdYhp2o3XThfGtXV
bzX5ya/t1YFh1w3v6z8rxgm8aM0Atutt4Jr6N7Ajm3lSCEBTFnU3LZcZOw8FVD6Z
y8+25f+cW1XLhpnBgdo81it1QLx9U7vwnJt+cV2cNvafJDoIR/IYli2WBcAtpqdu
G/L1DGi7e6DPk4Irhbup52/m9vJOfnf/kZXTRjWd3cV5Qb1BZr4dVQl0lNU7Ycpw
Ql5M3uqGdve14Q/pEx7iDcksXmXLH2GtxUzhZms2rYUuxnenMqbjez3sInBhIaDy
kQti6W+i4bxO3LOoffHOwlH5b9YM+Lb3nLLxJqSX9nkp77Ig9qrrlo9VxXlYuULB
0UbpSexMxmb5Xi4Se9YEZTtijly79PonUJB1jwxSJn+OJmaixdwKxFdF7y1NbEFc
xhnykuzy+vZj29v40nFtCOW58p23rh4PNx2N4SrLCNU2WyQvFxgO+3rnEaAQ4cDg
FQT2sa2g5w6PgjtjR7fQebsAXoRF0pjpndNy3vVQQjH2OcRUx5RqW+zIEb+TgW+o
9zjmaMoux49H6F7Ef0vLSIQ87GyFdb/lj6VWiX38Pmg2+aF3QXq+nFAE73MxlQNp
0sOAqX5yXP+YEHH39UJb/M9uvp+fBtpAlVuPYQRXr6O+efaItjXdz0yhtC18y+8C
ndp08h9pO+ichumhs38jIDsj5nT5hVR9x0R2A7HQgnk5VybTisqgrmkD9VjHgqSi
ZMlVnmZ78Cywed+wn0i7zspx7SKpgrSiwXlbVrk8DzPh3n8tITNRDOCc97/VweuZ
w1fvhBo8GSDiid07xpdCO+rdZs64NGnIdQwuDBDfTfAheBUxD4JekfDx698UBg0i
z+CpeRWclJX1C//Qhx9bnJyZClYChyxNMZakmhHiJZBxK2Sqirmjws7FxbK/TPT2
rV8QCLUC3cf0NjAOrclPEVIgRDpxgn/FDN4+sUYNIhvyoLTa06pBhOY4gV1zd48M
sS/gIdtdAhjpYEU2x+YI+7whLYG8pgJ/dlXS7P033YDpKgoRLBF3tJFEH+SXN31n
XUypL7gJW9KiSHKXF4sA4CYVwzGe+xDOcOYeexIokmFxl7iM6sPlY5pN0K6WCpFo
1TtJ39pZP0ADwOc87t97EZQv9EtBZe1EXqv9GexATi0KGWnrZh3QQvusX1VcnQxM
DnV0UYnvKtEQkJga+v1zJyPtCTGgCRlqfuD+MeShzAB2d1QUjhmfXFU4fPI2wLND
LNRbjLXpEGLRIMfn4yLoL8J6xzP+h2n3pJdebByjGiZdUrGGZVsx743EX8uSPc60
Pd+jR2//etop4uYam1mOJBXF1L1PvpWyqdLrB9uozzMvXZVyHSxP466sejw2xy2s
iR2TGSL9bYNuKndQ7pTS6zs1rk3TC0z3Jg8PYa4CC/LfnjhZO6IVWTP1UWxJqTK4
qfMtGxJzdEdtx9VoIVPh/pX98NrZmFrdPtpKGjpOEKM6Cz4O5mjL6F99r5kOJgju
E+or4KBjOXkOXzTsiHLN/uY1OL89FwH8IZ+h7Lo9JrDpP8mv1SiKiNXenTTvOXbB
BOGC2zM8WknRGuwzRW1ENMlHLdU5FqQf83+Dae7Cq6VWfRO234Kmh0EIviJNhbnp
EYhRIZFPwYPDGV1LsXMlXcOjTKF7HnAEeLMFUwUElvmmzdf/mx4w+6wYwOcnaNHm
kqkMd3pLNyXT+ECjCt0ErjAqzR/Hxt1nQozj1M7hiEQvsVFtNkKLEL383q6Rarjy
Nwx8XMZOOEQH0PKg1glTfVswbHmNc0wcNZFBE0Evc237Fkk88owQPKsQd51yoD0M
CJJBFGHj/LiM02L0HDzoMIx/sTmebV5yyYtsGjL+KfQFv3GEB77uk/XPUsaAh5BV
C84CQwLtZZy7acjQ1/uEwueNHrpQtlThkL0OyiLJzOZtreM8Dz8zl0cocrLId65b
AI7VhmYK6EG5FRSaj6eyfUlS5IY7+jUwn5TngK7grNj14Gw6rWvXRprt1dDnCXsB
XNqKU+7uI2Pqw6Q7AivA5C5lOQWsYzWKjIoa21rtx0QaZGbnX7hO/UTJpfzGtXLq
Kk9XbVyhr9TuwlCK3Uylc2aG1bGoUv5hURcPytPjrvb/Ds59xeE7m5QyNE6qAAR4
MYEY+Dcvc+89hVmsjWAyrkVNFbM/uJAG6mKoGngi9ux5XAy7S1NQyMwjxCq71e98
rQZf8V5g6AcYhxm9eUyyyGWlscsmmM57WzKBFI6BzI2HW6oPR7xEOEfrcOqklqMW
W6juO9iUHTdPw1FdTZXTHABrczN2rL3AXcQMb+g0ctFDzsMfSqR2wIyDg6edMPP0
QVlntuD9EoW+rhLFA3EPEV+gPavrdw6CB+tPViK7TU/JgOYmJRBdXMLqNrP1EeOW
ez1YjFFlNEWIXd8VT1EFpCt0QAqYERt5N9X8uE0u8vpje23xC1IxKGAfUYVvA63o
4TFc9Y/EcJvZ0QZSz1oeyxfe3GarjZyzlXFykCTaizkVhy0ijXDyRYS8Gf6qkzja
dEstSrH/BC/LNsmSAYkwm2ux9p4a2kbTpKUBGnvitnnzbcE1WRq+5O6NSe0kPKqD
ZV5Q+0XiXEsWcdYhujXhpd+5xiUX6BQjx/rsgNEKF3FvaQqSqzU5cydhdJiE/K3B
L6J/fH+u5CoBSqNChyBpby/vIlKR4TECmHolxZaewsgb4rjmQ8z8lHNNaBO/gTAY
bqBGpDNvQ3X0OcKt7AyT8vWOulV190JU/N7yMdLwy+KttdYj3XLKzVf5BnqviGax
B3vuFD9IvPak/uFgwmZPXi+ge9lkO7SQRMa1d7gTkx3VHMeK2s3GbE1Es75zjrLt
6omsp62gw0w0SHSG3pX0BAa5nEWJY/0xWLVq5+bpDxdZB02gyMhQhvSgkuAzzOai
ukwRmMuuyfiFzlESFUcs8+SC9wcIdaJfGR+b6NYHgXeXKAv21KVXfW8iiBh1gaYw
8pgDNG9MhWwrYzxnGe/tqMs7aIUeLDUAOKtdBts4pnYHAJ5s+BTSQPhJD2wkQqWb
PErpoLk6Y5Hh+SLvfpQf/Hg1h/+aSOg6pMEaVIjik6nu5ra/29vy2JBP3RPhtCBe
Pj25bdx7myvf3clCMBIp6yKI0XT+DhAFJWny+wdnW4tplM+RmaZDTCu/i5y8FTWG
nAUQ5SwxvNgbDDw/EcfZkyDkbWpbKEPT0JMMdn/dDQQ/7xj1Pe6SCrkRKvzcy/Zt
iKmWrg7h+D1KYLJgout09nwS6bnRTHz6wNoOuQSjUTflw0mWLW/COjtpWyJoVnve
74BoKYCf3kTFbXqXbyXvrXnaTq1A6dN6Ut+detEfijxeTDJECtrE6OV2XjAcbZky
tjw+TvYIh53CKDMoF1GZvR0G9+t1QDHdlA3zzuL9/K78S/fgT2WymlSj2isQ2oFb
g6duzBUIqyVwY02YzQqa0f92z1qrREeC0xka8MT+iI7HLF9jeweFoG8dSYE1j2ue
kHkqw5rNHZE9cctNg0/7RL4wMYnvEfNQo7iCOL3+nJksvUmX8LVVQVTUOTkl+9QC
zbX9RPWynYxeDhKRXRMeErJHWnTZWHOZAghwkZW2gYWxOraQqoIn6iIe+N1nEepp
kweJbpmpi7uYnJoMSrVphsRHt7uiz4ABnK7kzoIdhv9Uv/crYsmkUQMZQah6EtgO
GAZWSrb14MHrFA5E9/QhYKwr+auihCRmC4DR+kY2XFzdqu0gs3aHWPSEmB6vxG8R
xnqP0JF5DBu0ZQGLmb3q4hIqQbQWyqiq6HoUxLPKih8OGx6UJWcbWwbPyt42pc1d
i8vCEIN9mMGDvO/Hpx9LVsGQl2TBWdUjn+49q8GCARXZxHvIjshfOkVDFe0g/IS/
sSfYOLlA9y8+xy2ef3bQyAyuGPT8RKr5+wpvelJ8qVdpOYQe+GX0SPQyRuylUgHz
vTWQdowrXRdkzgQlNdJbuZp4X/xCU8ct+EVzgbntbiPEaZXMgHP69Pe8KMcLC7g8
1Gugj9sc6X3HPylDvYgzyeY4yRxmlNs6V1KwVZk8A/UdbvDrq4sHG5+1i0VeK2Fl
wnHLZQHXNedKS02yen2k6cYKbwGyrdmVWccWyH9zPLQjy69tufwWPGRPEAB0H9UO
lgBEsUTU59f7q/M/v/W6n/jchD7a4nt0MZUxBSW+Sis+cx7zUlTkbXrlHLNF82TH
4HV4ogfGo0qhdeKNy8Uv8b33nlx8GvZL2iO/MUeMu+E+g82umiRp1byRb6wD0aOL
KBOMwdjzGK/p2EqaJPIDXPER4mihOLLlyHko0quhASi+5kKiefIJMYedCAeaWkvS
ttifGgMh6CrJtrngfwrKBTQ6sedTWXhH9xOPCIg6K/HzLel3qclcq+dNPka0E2eZ
9rNZ5rdfVcwXmtIsA5wlf6T4YCFRw7vCwIDNv16S4sKRTlH1ESE7GHssfRUp0+Hi
RD/nd/Nz5/MMVh1ZXSEznOwOjXD2hBBAxtGaufW6oqgTAwhIwJpONmpi6SoWdeqa
WCvOmUUeW+AaKf2xEjvN88eCXPFF2hQMdzJHjFy++5W46tgJeJVZg7kb0jjhrGSL
yQerlqWzfMSB8Ua4dusOK5NRNAH50Ymfa2AS+q0uVaX5w4bsxkk1JWCR8tms5BaX
CtVQGTaYV4ftcn544ycaky4imxy7GTK2kUhfIBBlSbLdTrsXpH39ZqOtAk27Lifz
emRNxkjEClU2UIqncOcXlUnZAeW6/JIrNUdWVonSa5C95ye8VpzDuiQ6PI6ByNt/
BrtOy4MVc6+QjQP7n7A5f0a5KEBmAq/DnDyKX9eVk7hgDEExWmlJ0EZCPlXjdC2N
msfpgws7pUrkQCEnT4ic/Q4b1zCaEUFaQFVHIQFKlg3cJFZ180JYhF8dfQ7Fvs0G
TuwEYCvy+OHkhFqMbaPzO+dVTAB1+gGVdfKEt2ZxyxajOUNrV69LM0PqsfN23I6T
sWiKw7v1mN/RHaFlH18firzEKwYcjPuWQU2VV0wAXO6gjFawJXkBMot5gDwgpH0h
jSThRT10gD06I3vIsL35zEXPJJC8bq4rXm73v2v66oLS3KnoUNo2pF5EfFLJ5cm/
4fLUXjuP862t0Z8lS5zs6CYri/fL8AKQysvCKFtvUhddC8gECjGVNtyRKhfbd9e/
OtxjcoZcMmD0SlWQcGIWeBQpDhHGfoyktSJ8Cq9RswjjwP8afxFFWaNRLvotNM/L
elOJBaO+ROswxfJFLEnK4cAcPBaMelsY8EuTrf40BfI2yEDoihmfjUmiOeXU5VM/
wldQ0Iv5D5XfWdv8i7USAYtnFCDGaJm0H1uGWrgf+bPtKiFfARHUP/JKyFxE9hU9
vo7y2wekaiRlx2gW6dkMMkR1SNw8NF7fx6puYnjC44WvTJHPRn+coNEeShct2NTG
ebnmxxWvv+ZXYq95RO9G1arjSc5bY2dBMO/i0C+OqTzBzGxCK0eCm7/pQIsvABYV
tglpWFfn+irnS6kJSZdMw1A1Rvk2Se7nX25c3BirekJkeeZdAotjTXTyZmGcsd2Q
qTgN5TDcuCJ97XolkJVP2sbZT/Mdr2sZM5R2plkGjmxQnpy4vyHfDYRPx73vYLpn
DliEV14MCiNPnV/idC1wQBYP2dAICRkhz/CKe3suZXRdWgHDgHF7WXkVpVAHPp/5
0GYY1aNKsxc22+rgWG9BHruisrSQ3q8WEeq083ltZHcQVAYocXvY0yar26M3JXHM
2X6Cl0L6PszCMh4nPmGc+XUjEVe5Mh6cKJ9DR7DeAKAnKNok+PLG16TIZ3PQvtb0
w+Oi5bC4DFIQfW+PwD5xYTXzLeeb0q0ugbtqDPVG/LjGuzEUfnK5p+XuKlxa9KNk
iRjZ2JZK4Z51awsI5kGKHeB5LJKPoGpocm4GtzY3vtfMhxOptGNnegNv6+zlWfCT
u9zH5mNO79caRCfF8kzZlE5YmOuxWycxqeDmvtu37ghhQlchGvKVVzlCGMpHkLGA
0IOjwQRh6GP8g6zrXTVuuCPvXIsziYRkbrAZLGfTUD6LH3F0/mH6VJc4+nckFzEW
LxEgHl2nVfpR1XuybYuIRJk8KGBVPR+DGtUeAV5/K6zyLvzhFZCmpQZnZHga4e3n
w/4Ty3/np6o8UCL7FQ1CWLXEkMVLSV2i4oJqggqUwZ7qMAXrPVIJUEtvq5I+mLFA
u4dD9PH3P0+aAF6Jhe/6PQFlEx+0bHL/O2vfv2B430aESpHOwNniuypDgZQrgYc7
NT7ZSWcdbOw4pvzmi+o7B7G0ff/kBlnkHE3m9T1Sw6sN0sRRIYY+6tJivVDxpuT8
oOGEVipFSC2bTCv4m8fWAypEv2KKq4/YUiXkj6O7cueN7qW8VkpmZ3c4lTQkqoRe
/h0IWexkuUbW5hE57M0AwsfhHN8pV1SYWkJ4BEM7lvfp/Z8eq+e7NQZTz1TadQnT
JJwtfPMLi7TLqk2swHRHVfozYJhPmsRLClwcDVCa+XJj3DW1s1YMpZhBIS57/asq
lPEa2E/Nd8LytBURgCu4ueGNXsi0patVvvPf+ulPxsUFxtcXbTYjZkj6FE6k/sgf
MTs2izkdqmzS2ak1DJ6Ud2Uz0D6oSNncwLcZBKpsfNddoWsTMCxEL7qS3NzcsjcA
EoGuEMiIHWoWoddyTjAMWW3qixxgL9niy05gPYmxnmdPDeX9jRCt5BgMvRX4uXRz
UKb1Kh9yY/1HOacWDJlTxTPZsPqrH3GvOFPxGop72rfsI81ozLnNxXu3MXaXrBk7
v7OzjPv1YL/0OKlF3Jg8I/EdL+f+RskUdUzzPRK0Iyysm7hSyCBIRoAnyoRnGN/6
4T2WSVW2iZRcLFTFgYVHLaaaqj1BaXHbWVECsyykuMb1uLVc5WUJGLvWfwGVuiF4
8ep6FiN46OV5xttxttUlxXwZvrH3CBlLEH0BcfUU3q3Jh6JeUQKF+Zz82fwFVLhN
ykufWwDalF3ybY649EBUMcNRi79Io7eMkAXsZmpsH3r14XxsSwn/EGOZFxq8hdDT
i4Im8Dvhg9q+WpBJ7f5o8NDeLkL8VI1RW8merVZf4NNZDQeZgvdi6Y3wqdJvlfhq
i/uDYANhzKsA+H/pa++j0nf2St+cB441rElRhFKIeg2vJ+l2a3YfnsSXoBsp7McW
4s9PT0yr+RxV099gxFldadFUdOOPQXzk0qTja5TYuQQpbpv8iQiUYb/2DozubbTE
Zjzl+BwQsMYr88sYkY1iDTp8Jch/+aeoilX7wWH+2Z5G8BJ3D+/kHORSf3RCRM7R
xLAJ68pD5RO80CYtHC3r8PLbDZh800Bm/TOVqEtPIC3nwupQrVHSu/Dtd/FSxpGV
S/yA4QkKR55TLtPsuyt6Iw6OkwWNdG08tYjsHpgZqdHtiuRIS21cp70R4n9PdoYZ
mpz3esF2ENSlvsEgu+xs/zvULAcKx0kdap6OCvXjA3hqR3YxsmJ124m0f1zkdVSt
xVIxGXnXDrpOrYVdN3xyPoPFQcrxd+v1CCTlqgRu9IvH8MoDLrkdkmS48wYj0le2
pKjDxeV9kePPwZkETWsjGDR0CHIa5DqRwJRI6NnRc97JQfkNFqoyLMq6Op7m9Xwp
kwbu7roJmBZ1gQm11OeFlwP4HNeAqtpxXpqCNpguX5g00BKsNbqA8B1tHEqZQlLn
GXpUPLkCcC3LXdKfu5dlZRUO+rzRL84ebKFBftVulqJJZiMCQNWKIBo5Vgw7BZXD
AzZy4FjNnlydqv3SIaNN4cIWlcz8ddS77R5iMuRh4vPZQeTVGasFPLjW/J/Za9yP
hs44jRuqfZAGVu8tkNLRXQ0BYGzlB5EOgs2OV4oT94QZ/phcerzL6MiIXiesBZ/Z
R0zwDDpe4eGu7XbvcOzd9KfhS6XIRTWSOCF9prh5+nV0HQ/n0cvmCNUlzbkOU34S
7oYR88hjoRakZubXl7yln0wjXBW9AGqXT7/QpkYVB6Jddk/uNQt9Fre9rGq3kTa0
LJGnZK9cDu4ydBogqbE+7hcjAFpto1nqUpYS7XamlEm4EJxGg84PkS1LWeb1i/4j
oW0eTkZAgfQbpmvPG4WTDAn9BUZ65fBB4D7GvuyF5rq/7Zy2TR8skE1x4Y4gkW17
9NZgG5VJw+5Mu0GNka63VlRKYuQ+e5OGbp0/jczozHYxybyid4ubabT0tR2dfG/R
HYZ+akrCtyRQHTm+Dy71Tr/N6KqAlJIOo4TvMjA+xBXoQzEkxY0WqvYo344F9Q+W
WS9e3n1Loo+romfbOLc8w+OlqOOODXHVhylWTlRcy3s16OzHxYKKX74OOhh3kHRB
h+/N+WjeSfH2zFeFhU2L14CsMWxlJycYjiUtnl4HiC+rkjF4p/1DDaw8BhbFTDbi
JNQKJea/Q1LlRgJOPpvyc7Sy5WBYk2+pRgNpt0sZctXTzhiDDaJz7Gx1IJK0SqvL
0Dz6xyUEIhZMdScuGrXeVDaIsHRu+ISRBpz8EXSVTfx3vHNXZDmpzgASKB6V7bNF
iRZZjfu1A/05Hp2W30N/8poE013ZF/7XGHxmydPgrIXGzctdLYSsbSTqv7LR2siv
DxYWyIMzkqepQpK+3butA1ITF2+2LA1Vbusf2Kn8NTH4gA8L7NHPcpmD9V38L6eO
kOb9sRlNZ9Ki5UbRZ1RG7dxYW7UFYTyVonl3Ck4Y5YDLmEJb2hAivwyk18fCUwBa
uw0CVaYhd3FQ6tgrK0FN4jU0cT4eoPyoHfMn+sUFoueceRy7vz/lLGF9bLBeeyje
BJ4J0v9hOPHqIcBaGDoYoj8zn7LfC3NZFJ+pi4INcpXDTqYdqg1Po32vpvU52gV7
8TjO/x3HjUYYIHmM8TNVUuF1KKqa3z9tlRWmXNGLkSX4wXX+P1En41uUHYEg+WjC
SjLvPPJVqORW68DPsIQu0k2fUy+XWnNVt20oD3d+G6vQ6Ekm2csMoye3WDpkI+l1
7KyaoQuQpVtTPJ44b1RJcAGsX6zN7aunHRwKdbmHTZdVI83P5lhoHIHi4Wp6NjgE
Q/r8LWJkAYS0w+pcJl5VpeRSxLQI7Eh5r0QGo1mHkGT70DSbIhaydJG6j/5QdJ7C
4s1k/OCYel/ZgktLvz9/Ba4+OPMe6Km5XfkTvfDsKoZFNKM5lUqlo1TRSKKrQPZL
WHj4n/yGqil7/mmw/nXVW+QNujH/n+hM+I/TL/rIR2z/KOcDuxYOevDA8TSxsFv7
6c0fD7pAKEPfzB76x1ZEeMHtGZO8GRc9TxTu9YXHXav37jNczFuGL4XjstCznird
UIHkMtFsPJ9Ifezods5G6iVvq7t+wYBZYPEAwxQHdEH+Jw4sybLuhgXp/RtbM07q
Cffk/l+bxdq5DG+Xq/ZukYWSSj/gxqAxedR9f3nwvi/Ktm/6srzipTR6e5ov3eJE
MTjjZfXocSYw1jSlIh4zRWq5i2Wqww2TPqghQ3Yy6UXoAmWuWs/N5yZcOS7ol1nr
8GrAb9GKI38Xv6a1/ij4RJAMGgMlgPOFu/7Kk6fKspsiI6D2kr4zhp1Ii4S6Gp/b
ejihzlp5dt0j9AvpRVDG8XjMiool7/Xk6zNpvj/xuF47yuiUqKg0Pi/bDkZ9tplq
csE1uOPdce3ugTsOdvHDz4qeqqJQ2Vh2pZV62iqYi0xNNBAEmocsu2vXOQViNNYV
4A3u8s+4/DJEnueHQVuxxTJUbHtb4E3iQOpPJOA/ivAnbUQrPuNDFVMuxO+4RstK
7D0UciMoB/aGhddERfY3YR0WWw9H6SvkVDy4prIS+2uYAuRIqDZ0NJi9lxicfRgv
K9NGcSohofEpriCV5J4SXTl8ZztjAHKwC/nZoP8bmvn2bRBZUfs9nw2ySCTg9E32
KDt2PZ8k3759ldNorpEiSXmkAGZyoR0WtzUqQgqf/wqSW66wfUXkiZA9BJyAZOur
Pkx3z4gY8WRj7cjkmniIvKZaSLDulA3m2+nqVk+U24MvJdYagbFdI2s3iqUNIfYX
7QbxjP/ZnDH0HVs+mVszyp+Omwhzk8Jdoeslxu5Za4NF7ZRwY53e0B9mHdfsJRmK
vwuLHuIgFMC4U9RdR8APg5p9ckvJ+qZsNzRmuzBUOwqoHoKSoAwR0yioj9geolku
XSPR3XfqppClCowADeLS0slzo+SD1c4c76m5kKai4gh4X9nn4DiNdXI3u3aZeaNp
Wqd87kfz4aKj4Z/ndqiqAhnnDmydMYd6VzCU77anBJUfivuiiG+9yW8XiIsgdRAC
ugG1YZcX1oJi3IkD7u03CU5+nS3KzyMNo+PzvQWJsutQZ3ztV2DM8rb3k8bVmDBu
eLWLSsnVydhlx4ce+wDFGPGk2WTlyMry8GJMBMgRYL1BwazrOHeIYyt/9uPvAwNz
Z8BZUOQowe4BaMSEVnsoCNtPpTpv2I6JFkzAC1PBYhTtrhPQfON3aNPIpQG6mJsL
NstoGhIR0//bE3rFHWEs9FQmFMEbz8ob/81STrWVtzLYhTjrDPecGGBgrFPek4Ts
UnDB0tXLHt8rkBWDDLFhP6NAVc3zyohsK3T/9qyXvB83fRLm+CzT7zZv5j3KsaEL
hj3rw7Gn3BCsa9bDJAGRuwagHGtVFMsvTBFSwHtRsBgeBTXZV+LYfa0qfoOHDeVK
Ordvx2c5vf6QVYjOXz6q3hCUHoDdDZqSWLsRuvwDUXF+0TRkJhAbRKjEQ8mamm0e
xl+Bugm5J9EWxBK79tQrR3+yNQTZit02VHYRurL5BkTWzVSf9OkJ1DWnXhejRNOT
RGcW+Y6G1G1P1tyIW1XUp9ggpCbaNUgWII444wtZkSuEE/RApZf29/4TSARaEuA8
PNObbVKEjTetSbaZu+Yqiw7EAR+8DJdzcjDt42xopqreRizVFV7PoB36n4Q0iaS6
cupTHCIIWX7mqObTGcaXrk/XYJtu57/Zcg6dFfBUSWTRA0pZo1iEAySwhkuVhvGE
eCLREptjHHUXjfXIRQrS42Xz9hF05CoXtdb/qVYt/EIGztVtEnzEsxVgWrtL92EM
pJhW094EYuIWPlo7dk1MW8unZCROuESrROLx2cE/lZgIDE5bQZUtHBjE/SJwFHi9
cYbebMORcjLhiIGuZqTL9LPeZnbzS5fXU0Rrl4BsLlu2Uyye4IJTxLBgBaAbLsEV
/Sek7vVNDVS4e1u9m1D3V2Cc3wpGqYzKSsM1QTmAoQsdRuxQ/0J7jnD6K1WECs7a
FkMh15dftY1e+Gx9yLizVW1sQclFX/tQxhvfwGCnxwOS6jPoWb7ZBDGvciy70Q4W
Wc0OJOOLtjb7Xc3Oyb/jDMd6Ht18pDwavC/p2UjLEOq466MKEf7p1oRGVpR9sUqe
otX9cI+WPIWTkPiK5iak3gWR4KKyj6nAWQ2X/oDQryD0ZzufjCUfX+V9cg5VX+6G
tpn68LheE40nyetPjN/Hbm8oO0PJuh5A7VzFtFHM9Kj+zW+Sw0T5u3V+xTLYwyLO
nJccE7uMpM8Ncu0SGuqg7J5Mo3hJazbtrzHxP/BAul1PB3QENBgl1qfS58SHu7jW
lPakLvTa9zJjN3f2xAQ+FXbKhJtYfUrxVuERMY0hfLlvF5BoM8t4aceROaHSU7xq
FZQe/d2HgH4JOKzSlDyv+lyoZWlZFAEi9lfisJVJd0CSv6n4QI5lCZakTFAXlq7G
+I0FFj84LMOupWd9c+jhHLU2J8/NDPiB0YFVgP/KsxjZBwd42sr3OlS+x2HrQrxp
qtvaoliKPHEq3th4CLjCjBmVYFPUE2Si6exLmB7ioaXI0VhbdAZMT8igZYyXWMAU
Dz/J76p8FLz6dfgKqzJzJE5tnJJpgGzZcuEyeesYNbAIt60jL4F46ghb8CavryKA
1FzDucBF6hDKNZik0CHmR15doxxX9Nqi0WRKezI7nV4gawXuEXixJKewKZkLK0Du
qqZtlWqIErY9t1VhqDeIgjDm0czEX/jZ/A63cqSbuhbVeK0MVFw0ymMPB0NTL4YD
nGUYleH+CHmH3iR2/QMmTHwg/cUREnEpCPnvf31w1QXkzHM1KwWeswHnWoXJKl7M
GJXpZgUrPGHXu+JKid/RwT0+NciKDVhSebcOYNPm9aMM0ywVxbpNFVY+op+g07L3
lW8WMwhtoYMlleAUIDhtUQMoQI1QjufXwFdVW6umqUBK2Qn1cnbe090fgsKkFTim
8Jkvi1r1BmyPWPa1qyuOgPRK6MOqW4xrILy4JfhTGacdUJE98V6A8hQsjuRV/2jk
cYkcv0ReaeLEc/lUYtGVfYCd/hM4CeE8ZCvmyjFnPJks2o/fvrYjXfdsCJ9YW2MT
PwSi4dbFyeZxZ+yZFBpsXJpM2eUkEOIaZUte0CeiV1HoZ/q6YIf4uk+Uiz8hbPYU
3FVdOlEM9cCYC1L0Ow5B0odzR03zCbsL945ME0D1BYO7NJBhjMmmy/gNxuPuBOzH
z1UrOYOZ8p7pQaFm+TOXJyiTjQ2fSxeUjo986MyBKUc5H8n21RaG531BxvS6IuO+
O3Dm9nZ5nd61FAdBt5wVsA211UqsoIOh8Kw4xJ8lhi50qvqwRuKuTDOTxa+FetJO
+PBHPEAM7yL0AeyklkimiUGpwbAegrHF3zVSZ6BEDa74XbNID7jweODKkJjyhkEH
FmlShqpXLZBm/RGwEQr2YZnn2VDR5pEziWpQd6NrDtKefp5sxuwoKxXFWCxLrVd+
XP5EiZI6CVSmVHlysG+zSOPbM6XtA/q/VswCzev1TtF/ItHLGkyk3B1yhQxVmOGI
8kLAlZxbyEglFuZCt+jURM7tratnHNkEzxpoM8IV0/pHjEYl0gzIFK2W0k4fpgnn
Dzc34bY4Y46PM9yh0/eVk0g/37OkG56KAxte+F8/XvVNTFh3btQn7tsioisE2rTJ
AtyP9IXdXde/GalkyXT/wFA/ryjDQEX+E5n7g9yEWInipDhKyGHRI6elOQGD/5Cr
xFyalCe3I8sjEvbWD9FZkgBSwqrnB5TUnkyAk42m44coJyHaJBYzvXb2+a+mg8fL
FZwgqyQkbQ4ECPBkSTtX53GrXyD0pUZ9lybdSrHIQ6lipkT+yY4AUQHQYR2Dc7Zk
bzhmUsfdQFrNaY44nuVMeByNqY07Hp4/0GAT4nBHiC8gY8wIf/siuj9t+IEMgRSM
BHHEvCmk1DZUCx+6qABbXu2GE7w9vONch8PKBKHaN6Il5o61Xgs9Aj7pUkI65By+
k9eShat5+vxY/J6jlFZz2kpwLuXEBDM9DW6hzoa0W5WeoJXw48hDa+rYoUji16Nw
TIp+5K8ukAtX9jUSWBC2PD8EWzgPT1wYRTXjlZzH+a6ARSpu0H4jXQtl9NIa33Yy
Y90ksHz4UCWOC8KqmgBXC2pf8gwl+XihdsReGWcH61T6bI/n8v/Z2JIvic6xor76
Cm7xvY2VRpeFRtXnmhBaMtYiUfogazmyh0qVBuDkCTBdSyE5LZfkNgXKrkvBDy7D
Re2S6+CsbDgP1qZS/RLWd1EqXqek91tbuoyOrkAkQTbtmpXGow0EzxOH/RxgarFX
JAsBzD2FHt2WdNilyIG1OdWeCiqFRCW7t3kLVafz4+Mvr//uM4epTsk5EcMyJkcy
prU3QXF/BnBh4g0wqen3a+GtehECXSZ/1ijoRbxwWT3X7WEvjyzoJ9YYf8NdL+JQ
fWSh6xvFxoiGPQYwNW4Y7O2le+BOJ1DJFExVybNdreRPfmJOQ8JaU34EW+XC0T4y
q4vnj3qAVaW+9FmQJoI+DLe+0X1yTgJ7+AarVfuszjfzw+B9VRtuIMYedyhgyE3y
gxhtXGhsJ53/IXJsQXCEvVtRhqbFG1xlAcOyr1+SRrOxcvQHBYKxoGX9kswkUyyy
BBRCJUz7QjBJWRfjHDhTw7pS2CgTzrm1lLJJzPLfegxea1VFfDJ02vx7qUw0R8hF
A3q581s4TwBLIJYajeBD+jxTch2rOn4PTLN4k4mxk92k6dpLYyfIkmOKv9/aKx38
SzRb1feKPihwil+b9/3INUSEc9519OcuHhEgQGRyJNTJpzWiNebWgM/SL3GJnfig
LjHLEuIisNhBtbwFAoraLdgLiK5qbRiBbnzadr2P4/yYrHn2ANntOkpt4Y7z5CvN
mDQwgNKKuGAWYsM0oB/13O8xzbkc78RbUiXo90EmZrp02UiJPGnAC8CyBUSvt80Q
VKALFFZ1lMNEi7K+KTHyu5aGcDgqhhOzssVAgbLmKgVgor99fb3NKjFumRgw0opW
pkbEFOIKhYVnk0aILj9tNA4CPNqRRpQ9NjIkmkOPgCRwTfmmoKh2WRWQdhErC2M4
whRBk0/sL3yBUOcJ6YmBkVO9RWvvwt5DMM73ug55GAquI8WLXvcAM1vZ1v5blt6q
B4C/QQEd8dovM3UlXZuewR8SqWpeY3cws4voaDRxE1517H/A3aqYpSz+QTcnVU5/
A0YNxNRJWFcRXz97gj7QoTcJkRQEu/yfiHuk49zpOhJSMqse798N9Fg7waFXfmU4
21zOXN+c61Ev/DBvuEdRbOGIAExa1bwVTRD+GoXb2UWKHlPh2tp6fL9SyE7VvChT
doWICh0QHC/EsbU5DuhDZ0+yBwO3cEV2CuMXmc+SoS8KEO/OyLPrrLeL26JdLCqE
OrAjf6HkxXo3qvWPzdfnEzSxv26kyxNS5Pg0OtDig+BOWBYJPo4DUm+u3C7I4Li4
NKXaz42QVFfrY0PGJCGsj9ZH8OSBcrKyThB4QJREJLsYHPvn83CqNfcf62vHWPO3
h5hjbdKogVV9elxt3gyjyRE87j9N3o5tXjsxTtfOLfhcffWsJ0yKXgv2NxRbwQ3f
qRhdhnmeCumOoJKm2mD/N/CyyirZmQHfvGgv3Ssxmg+UM+p4fVunT9DdOYojeVxF
YZSm29o+Q0dz0nLcn3MdtEZdnOw6u0ShIxUegzbi2jdSuHHlszUDNluUNRlBATay
B+EUquzFwtkohiKnRGNWNKQ6CSkmq3XQNwveT5PXAoEWV3nG3E67mblSKYJhKeok
s7EG+RVQRynQAxxS7990biKNifEme7O6wQCY/shIp8GtdojnLEL3GN59sLgL54lR
Wob1s5dCj8k8ZwY68yBl8RBza6xjGxEFX4g3/25E2teXDW+BR2Lovc0eHj1K4p1f
RCBbO3s6pGbthObXs8SorZSZQDb7ZyeFscFz8MV91uleknFs4+ldg0m3TiRwFlFL
yj7z0WabefFVbovrN9gdJm51y9VZWzZP9oSdMV6ZRE4u//59jdf9MtTu9hwBv93C
dtbFRM6GOyQJhy06W2fD+fF1KQj21LweJdQ/+XK6x5egehHOencsoUbRBa8Y9vCd
pWdE8NgxGEeVchF9SUATe2KAORrKXDzR9tidaHoVgZbUpOqWGj4AWiuUDtniEuUQ
9+0wK5Rwkyfrv4xRObSgIwSva/gUErrCxNCVpGnCHCO6Xq0oG6kkXrnkV38NzTz7
0s0+tPmaS/Sg+RNBwovaa/RITwdW+NcFjTsWyG5D3zvFRH6IEashNVeQii+3dTdZ
PPov5zKa+WV6pnT8reH4/HJum1u5MbGTHgRU+eRpFD+nQCqdDOF/y6r7hlbY5can
kYiUln0OsEkmQ3dO24C6XBL6n8Ln7KLQL7bKoYs70XOZgQCiqwsOgY8Vmf1Qt2Mi
JJ1tXrInVyh02DenP24FQesJ72qTuwlpgYpaRmWPjzq3SLaKyoZO3BGKbh74oUgp
6trm/GQFDumnlDm1BhOyCiaGQTZFFU0sd5OSoj5tH7PLpXOPMUSj76sPFOZu8qzx
j4Mti8b9QMZjcA/x6Y3PZR0cReBzVUyQ0Y9QqIchjlZqIbhkGonv1T52jGycwCnk
zJ5uEFjAzshMdOHTdgrV30R7xmCYB3GKg/abGLDRFKrCW9RSRadNheazszlh2jqN
belS4YoDcXwwTmvABtYiD2V+Rwippw4GDAUjab13vLdohlJgrm9euxODbDZpC3sm
W+zOp0Bn5drdk02u79+jCRItCT1YqSzXpN1YJEus5VsaJ39q65gXytOgQBZgG9Pb
VPqhcjPIEMZjhjJrbbaRhB0DM9FiJJ2OkPmg52DP2sUmjjwfTuvXF8KG9ZYhwn3G
5IxP02g6gylHet54EvemmqsRKpNEUgBuMtTs1n7T6FeiFz4Kf8NnS6cewBn5SEi6
6cO9SiQ04sJG30G5NMjRaC2TYn81ACPivF1oa+pZULslYv1xELqyPckgRKgw7nxz
G3EhebfJ63rPlm0lpqShwjf3mOoXlOs7Bs0fjlTwI9N5rCwaq5srDj8ISliJoIqZ
5jtwax/vYi07dgwl6yn3Z6Sci5MHJOCLbXTZluDCKsZND/r9jWB6O7kmI1iL/+L6
ynIIlD3PNT9IufPl+pHO+NhR6il1IclSv1JpA8bDjNZ04NHbXAkmHUhNbti30Jrx
fm2Ex9G9RP1+8aY0upyH7B6tP+jAfdA4uZV4ERZso5Y1YEOprNbIzqDyGBxzGAPi
C5Cr6zaV0dNoyC01MGVTNg8/hh2ERIRpRxvTnukUlnW0JOekQK3KFHD+p2rmI9e+
wAnHJ8QhqA1zaEcZDgEoQLfgUJp3YpJvj/X7Rgpg0u2BiDdhArHTwjsUN5MOJtNZ
5BS1rTiAD7soY0yqrSHfvzSvChggYQXtllKihyWDFLXWNN6qpBCWVq9rUfXU9gmH
4JO53tBtqt/kAijRQWn3yOiXRFhLM3hyrkTc48PogwF0kKx2AQusjlPCE8gANjJh
8VhWJpIJ6o0otJP24X0KwObXsf+d+z7M3hQP8hN/LSX+RZ0U9T0kFIbqMAunwYwM
v1nC/rlOp/IqsDpJJa80PSdZsShTPg+RHu1M43wkUUwDrBJi54Oheb6F1NRfycTX
E01RrJmbprWhLkFGu1P7Y+/N/oEbR+5Ck6nW3GOfltbuU5C3sVKf3zd5mrz4C9ud
G9ZoPRKMH65MAFFR8L09BspCHpcEVJr1t8TH2sRnkDUVhm5cfwdO3nq+nEi0hjKY
0TL4KuquBQdtFxmWouGJ2VjoOYtszL1aDR1MFwmXgl8MErGcwvt5heGI7X/3+sFd
cLEQ2ALiz2qdE8K6N8RNQ/H2wYy+vpTVeQVyHAqFwVmSykrQDdgOMvoDn8SocAoO
PJtaK6IMtrXAicF8bO93D8WSFq8VShuQbjSZxp8oT/AukuevGd9yEVzSXCNHb62h
mlIrMn0/zZBCAGPh9MWvA5X6HqmiAKw7MxL3ONhx+XjcKgxXf4hdS8GkPk9Gnf1p
vakXJNWvvjtjuL8GN1hed8DmOeowAsJmER0EiW36pE55lQtadob4Bkf+czi00io6
+pCCNUsm3smqDOIgZSw7ruw85ntd510YaZYu8xKNdlkCQ1zn4aENEkWdCxQZICmy
NdCUF9Mx7keiQ4QnORKfUFANT324ijO/q2Js3fBt7LEt8TnJiO9Z4o/OhMn4JuPQ
EzQuSxDtK6fy0uV3E06006up79z0iEmQOak8aM8HCLeRmH31QxzUrXJtitzstDRB
8WaC4vSNlVmhbJQJDd0Xr5Y8t2f5L5LSnzY1owq9a/UmclyBNHNgNo/TayNOWY80
l7DNwgZAGH7U7+YIvixXs44QkqhlBgTNGtWH8SgaJrWVbkBe8ElBp8VfiLSgMaSZ
yy0sQW67/uiRblEYK3Jb4kLveusx1iJyhWdCSox9plvMvht38R/NQlBx8O2wRU3y
Wvj8x2bSCPATyQ7EWCwVSSg8C+Z0nTReFafUH7asusib4LxpwBaJBDEc9mz+gJyg
Hd1F4OIgc8kRiTr4yeXOHAF9qyBivgifx2lT/N2wS9WqZAmZJnb/wDt+tG/BqcaZ
IsvwZ0gax47Oybq+Rxt43UWshPqcO2fA9DDBIsuoR4oa+zdpjPBvdjiF+VULkWPK
i9HnMgm24KBXb63YZobU4R3qTwvpzz7e9qImjXt1qYP2IqtY0e5KEX8ZLS6VKRkI
cqL5dhq1N+odexaxBXhGY2UqDtWMPZ17dWthKBbADq8b6by7/rxBRpp7Rf9bj1Qo
Ovjdo43WRulxYhyb6Ez3aZkMWkoqGq4rA4SRpABy8mEHTOpoJdfhjTIvY20B0XPK
vNwkW0HsGoyEarqUnuQ7Cz66iVuWDnToQDYCmGekD+jzcplNvWwFwHNVv504jgpJ
yQmgDFuadCTWUSjCMDT3Sb8frV9AQSBmjmYgP1zau5VkXr41vVctO+UsWI4FgGgR
IQBapBU+FKvqtVO6EsNZgPe7BeT4pDFx2WS14ReMgJqRfFM3bU9C6Dy2SVM6qvQm
sYL/OZHw6Lk1KG4mXtiCsr3eSQAmWqZgc9FYHTYzrgaia+IgF6jEtgsa+gNUtx5K
7ZcY9g/JCf/eXLb0nGKVSs1FvY6rrV3bZ7LdVMVtyxUULYdwQIqb+WMKkd0dfMD2
ImvVTWbGALf1EwnKE0nzkan6euyrg81VCS+mEpG3kMsgdAZbHnpj/Bg0ciQAhGDA
QqWPnkxLVg/Q6e6XTo2FUcd8AzWINtwHX/JYyYhU23vAVJGaXngSyd6ZvxAMlPkR
ywtPJfOBlc8O3wl502JkTcmKzn1enwgsOstBrItGZGvt9o5OkaMe9NuqXWtOryRA
hhdc4zSpQKep3O8h8fUlUxM5rypUlj1QgaRW+MIRJ9t7ase3WVNjcALe+nVEv3NU
jsI5Fb/D9dhfRFw3lsZMDA81ZF/BXnfRizcJ9K2tqw/UiUORTeeaDr9q507iIKY4
LJS9HFVk70dZA34W+TW9sQsEuUTFmYtQZDfwCwUWh/hCMoHoo8syIfwcOOqeQ4ov
9qwfIrphB9VHcB9ACYFdZCnvw1zZPB4j/pRiSUehnF8fr5wI0qbCxXBQmYM91j/U
PMRyYo44gjC+eZclV4XYV31W1uiuehmY455jDHSJ7yUyMdLt+G6qBm+f+CGrMJPC
cW2kNQf/roTXmgUxT6gdkx6OCKwpBL30pyDGr8dZ+SD/AU6ilya00k3gl4REZj5R
C8hAz5LVBRZxEhXFxCatIy/vocvkmTP4w+OXBaCyqM8PkJnS5hv+3oXXQ+i6WJSz
v91F8AR93wgMkUZ3KAWdVCp8mn/27E3PLQMq3UlY1Iy778Fz7DW+ujUx05/cGl9q
h9kOeTLxWF3uPKodQViVcYopowLPPyEQdecH8PQtNaTO8tR7FlLOf8240H8ndNEc
iHyO5VaX15kGV3DWU7sQvcbAgNqjOYMrFVqB4cy0b0sVBgN6doAid1eOcZv6MkEo
OVjm4Ib1/zM0LHVP6mo5BNiXGWssZANsi9MC3of/7Go6rCy0EkVmXBrNQ1LyJ74I
KLe9AsGXWCILkXh7Sb17WGPFheG2m0ZVq6xzTiQTm663NF5CaS2SHG7fZPtXFP/a
ajyiy3v5QN+qcpS2+2dyc67+efM+b9I/aAe1b7FbXXTh0qLk225MT9ZYfH3xfsJk
N98JrftiKG9XuToAwEKGasFaikSybhBUxpCVHC+yUkma3UbHgxNn/JrJSbl8fUak
9jrfhrNeHnTrIQuNkoOnB6lba6zF54pHoF9TdnoVQ8O4LiJYS9qrY4t9GEctDIRI
Sae2S72xIHEEP/jGdEJzYuOjHB7zsrajwWBOI3TDMHC+H1Il2gpFzF/xkoG3s7pZ
kTyBW6N79Ath5IVrwNJYc6rWg+oHjdFI0j6ROqqknZr22sR4b+7QB/ckiIuNV7fC
QYqLw8w/vxwNliLEs5u40PWnoGwjbjPttyOCqBkeGN4w2/WvBRmbJo4KpXq9t1ni
+Vqr2wyBDDCKd1P5A+sP50ixChX/0p3R85zinzh1WMF4xSRuyj9iMdp5CpkJKtcH
wrOcd0P+aQENl7zbb3JH/ZrEHsOGl7HbWEk54MaJqpJ1NU61KQ16Uh4FN92C3MKh
n+7uOGK94eEbAlmvLHeDNvLmYbONMyACVYzyuXRtSuC5LsN2gnfMIFQ9RrwwpaB9
7Mo1BtobvXJf5K6+yZcXbfFJCSAfQYKrIASybHD1ZwFf/e5Whhxpk8XPfWcF5u3x
B/rnlSkqOudXsdbGOLT5SgInEREpqQLulaUzak1WqcVoyqT4Uqr5S+dwDqvO5FGv
XT5xBIM7syLS0dRZkiT9bSJiD0+mcCwser5IhyxbwOClxkOugCCnm9WyzEZc7mKJ
FDtujqRSVuqP6kFIRmzZe8HCmOtf3WkhwT4hkcBg0dbtYxYGr7n3kW7WH2kEtpoy
HqVacGN7il++nkfXYR9Eco9mj2RPftjBoFXRXjM62ytBAFo/CAxtZZejCjvyFLIX
hLFzM7xYXs9At+u9AaLF+vmWI+DfqfNLw40jB0ezNmYjWTAnq52Wz7wcAlDufLz/
z++cfiWucQ2Sw1bHG0T/D0RImNd9mY23ejUez72gzoT333b6H5yxKnlwv4wtbpAT
YOfj9nEnU2bRz9F7cU9m6df2KfL1EMUFQdbbeZqchcqORmwcspHribCiJkBbj+o2
ubKQllhpXByv8Z/DO9t4xznRzmB+Wd0PAVM1cNMk67nid5KKiqrlaQmRi7B/g+/c
C1BIAfp3l1+DNxsjZ65thc3vP3kZzskR/kKl4735fVU9XSjRd38oh8wL6FTcsbe6
iPuaIfvFbncXTSe+L54Ha8FjbpX0cI2zyTu4sqtzAHMsiy+SfwQ65+M0lf6IS06z
w52Xr5IRDXRy3safK614A+Zsq91zhpWWWAL6+zZHkpVn80Kr7fQTl4a+B99eIJTr
/5GPITTay1tgquZrHS9btPodRaAv1H52ZjFwE1PM1SH027+cyO1omNPBfcr9TM8l
Tsl9Ot4wP2tAmWuScK7f3ncGDFEdXCaMbmQVKOVCHbysew+MjGLzbk3gmmmY41vd
BHof35sd8tCY6EWwjItzJdi6YSFeYNf0yWg9+D0XYcFwCiGXbHVCRsfoLIQc49HA
cQteKyUkQG6WmIE0MGTBOF6/q3oKbkNtzNPpOUx2IZ6JCFgMfZJLK+npkqG1TQaA
l4Jxe8SXzLTxdYle+NdsBzw+rM/GhjQa3jrWzQWNWD/0q92pO4EDTzRnrAYQigls
LpdCZTPFRMg6nURVqRI1SMLlKefZHLjybM7iohgFcir43EoeXz3JcER3Rug67rGq
F0xDA8xzYTwaMTfsk5pZjofyh0hGd1vMH+U4JnebmCNBJAjmUsQpcbKD7vwb4uSP
6ubz5zmqmLigGxuB5ps6aCp6E4kBI+/B6rthcTEjVBikTvecUwDeSOWqOUxowyd9
P+t3goXkbMKknVjUuRVaD4WEJiujpICcaTWp0Me9oj64xLOOZVAarwEp704k8v5U
Lf9zPnz1KkjB1p/MWgRjlRMp+C8cV/05pVvy0EVSMGXIrl+WT860xbOjHdAN31vF
PgpuE3z7rYYynWvQda4klU3IBThTKIcOwFfLcLmw6mo7M+ehbu9/fk1N4q5NgAbu
w4PyKldwrGlHXMGCbUgYyNFwWqpWi3lyshK+7YjQZT6oyZGWRAa4fs/UNyOssjoe
BOI51EEGQ1aWFvtmCUxJ92feommAcVYWcPmMdqXLGEK53ZpN+eFV7GfF4wirtdDg
gP7EnZH4oPCwGHruygNvpllLChPF2CggFUK21g3xAgE7aw8k7vqNtIZ/wAXtdn8x
jIVcRLPyhMMG0SJCnszL4yr1bXopvD2y6IeuNEqckF4SG+4Yxos8VNWcyfuUn1Mu
BPzJ52ndEQRCJJtMMGKDre4/9QV5yaKRkWyshB7UULkhSjdk/rE/UbPSphHtNlV8
WhFSlLELfE54J2UZLKzP6vgq+ZyV7nCOK4IpXjDtHGA1T9pR2zxZA6lQ6HHxCHVV
qBqpajeHggsxHHk1nZZn+8csABfCorLfLot1DugqYdH5b8zmQl6d5PFI9sIYPd0x
wiM72txjCJsIS/lFvEQ4HHJrjeAmMdG045hCVKUPKmqCZjAA0ybLhLlp9NlCYwLY
bx5KCmYP5g+xhQ5D4MvV6fqv7/wUjj5Imyjw5lWcRVSwJmKyGLyIpzDM2zBLvLfZ
ruwhdgANXetNUCFQ0w1CbwcdXiQmDDanUBXzGuAbvnwtoYtg8wnROg0UvuiSp5ws
qHZj/irS96rCFkeX58a9XBcDdeh03e3Yn2xNaBcz3Q9F4CTQMEI2LiqQjB8TFG7V
hrU6h1JYX/ZEtJWTbwsGi6BzdYacP+fWJZa5aSaiyuFZgfyagajjuO2Y/HEc6uXP
HULWrBWzjBaFjjgTz9hduoa7sUjfTsD2cnQv5ykTqCOgrt1iSSyqFalusaRGpGfe
sv3U0tyqh+28/0Sa3kw12Sz618scT/dfGx/ccSta6/LKr9Q8+Xh+CMZdZns24H7F
rTPCstAyF2nkfPaZb8aR+fuj/HwZIHriINH4oSADyLcQ+dwyvJUGb24v0WdY9/Ho
TgI3plzNA3PDZU0JgAgjxDdSR/q2t/YpI98XNdJDme1GkcYjYDWAVAPj5O4mRlBg
cikwM/5eLOckz96uQFam3ALJesjjcYaqGdUFzEanbrHNcIip6kWet+Nrxq0vHAti
t1RdM3bcsoGEXkMgjXD83G/M9ohjvGI6/XSy5GHr6ktnLa9/frQG8+Wv2toryNj3
BFye8zIZL6RligWSAVRQbo8QpJVThsFLQ2ZuzjEtGu1Xirv1Dcflx7QroNWXNhRd
txy7jfYqCvwhQbU5u8VIupxMh+gx/FRpts6B5JwgEYnI4KsO9mWnDG4dPeFDIv4o
DfnuOGCS/GmAh08jn4rXTI9g+wLNaYX784/HW+RvVWXWKJQ/QPuTyUwzYD9dS13l
qwBx2WQzvT0JjLMecnQ97K5Yucqf9d/g7v96FfE8tGsJPalEfAa/pN9WFawQPVPy
A5JazQBeoFcjAPP1YzhMZCSLOfhJBJ3yRaWC5MXOtU/+F9MU4U9X5dhBiKia6Qw/
ETZDsEa+Kd/kabbLpeDq90TM36y3ymti4NjNR+rUxm6iqLIhEDuMTeLeB2SkGGWQ
dbFiKJ//RXn8iTPMs/bJ2BQ3JxGcaNRLal1YFixfbNZugwSFhnNkd2nEE9X2l9oA
y6A7mqtE0N5JVS6jGy1PVLnzRObB+40DogRpnFqTvXQBl9TMEQPoZ6oa9JuJNeik
FGvRQXub/kcQ7/dRP9sGemns+Y7pNFhyWW17McrRBxAMqersDTXz1deY/w27Jm1a
+Vwu3NKOwVS45bFX42CyRg9gMdMivggEh+Yrk9dcd8vVdNioudsEpgPlzS2B+rrX
TnPcqkZoCPTEn9jeg4ELyx+MslDwgeg65eri/6hdJUbdNMqgybM+pqS/SVyl54KW
qCXNPJFr7VglSeGgSu0lkiECHpMiI1XGmwAPRTuKxqbjRzAFf2oCiyDGkfg/4WiO
A2B+hB2gBVgThuNYkAP/IAhqXqxHdks8Q8b3oySjjm24QekvRicxjTGJL0pTl4Vi
jtT2a7GeTKKk43bfmezMYTfFIZatIKutS6isJ9r12kvhf8l4hUhBlHpzh+nCSozC
iIsmnj45G+H3ytKwdhN1PP1jRJeuacZea4ZLKl8/RtBUm7c3S7Q/E0PlfyJPwkwS
2cocg5Y/LPZKNmVWmdLMO1GQ5DixJEuJUqBH0oY9W/+HcYGEUcjAR1dc/SScaLnt
NcBJEd4S7ZlAp/697bvLirVHJstFtw7vet9E/lzvmYsInZw48mqEHr7zTzMZjAnA
tQMfHQddgc8j3VFpAlqwVxSZpET7mOgZd78TEidOLv1MESSyG9BFdu9DWjkEnGud
YX4GfjpT/2t6EB4VSmFVGBDimgrgPoCSXw0RdDbPhVm8y6RJuyHufRum7wlJa7QU
YfwJ7WqF11Mh0bAVwvGOvjQ44NN/C+wOVeTyGXNzuWq4OZ9Q7vrlSzEcVwf8vmmI
3eUEqPDJd054yva648WuD9DVNbxeKk11WXdIzzC3+J+2kB0rXZa6xPYmfMquAZDg
J+3p4JTL9VkcPK6HdJhSlGMqAIRLKvkZ1FgJmTHsi+Z4SIwylfD0K5cgwuqnrHiR
GRsTbRVefytcyWmTEPYZCP4Ju2BAK4T9XzRC747B1lNklviWhvmmekLDTofjbiE3
usfsFRtaGuZlUVy9bnFPyadN1BjhZU+5/0LxmsLHqRjaDkNn31KM5fetjguCkOYg
m3eV0UL0+FdgHV/wKb4beEo/VZq9qXkXq7oxpklkDP9MIahwqpHBj5B3vGHQckYO
pKsYR0XngsbXPVuMEQy82Q+f5YFgiZP0B/sxgJyHhyZxd+OoeqzabnbQwJuvweVk
Oh7ZbuovMWf4cHzJf09keQLLtHHoEXLRyf7VqeqqKjanBFSkEpJeWgthIrAoUsU/
NpyrlMRbkG/8ywsVqJpz6pNTvLtRjcWE4sDqj7JmbokjKlt8lKgHemmQ2MuewLpO
swzXjEUojt3bmUKA077/6gtyspNZ6ichz9XyIXMBxSq4Majt4yVtl3oZWJxaBH2u
hNmg/oOBNVNkQT4cj6GKkZwN8kCaZj8fmdB5dPvjymYZQkL7mNIRqvmpp0GLlwOO
5iMVD0lTanpmuUv926Pne6t2tByPixUwSCjHz0AdH2rV+NbfezjbLTmb3ZQ+VGx5
HISs7GMD8D273aF/AbwzX/T5uToJ44sJv7uSIzsHR40AVAkGOAyF1VyBLuLQ9uh/
oDiFKvcbRbfUB5ZwjKA/TztQUbN7FL2gr5CwYjVbqb8PCZjvmhhxgn/7pLPsLFh0
HJb5qjZ1rnPyxPjopprdS9VvBP9spEghxqfWu2W6RIdmcvsCm8YRkTJ5t/0sV5gp
ZgmJx8UIWm6UIi3iUSY4Wtv2OZX/fGF4/Da1euNZxiMKS43E+48L0YCOyYjh4rcn
8ayFGTZybKVEEZPQ2uk4QhBJGKtySkxFbaAx0IGLStu5vBin/MEJDTbu9ISSORwo
g7f8PDAMvgK4G5koS20pe330KAvPcQnazgpWoqP6LDht89AFMBD+u6dXQn9llPlK
RruQN0ks8slB+Nr1PHSBDhDsfFzMw3zpPp5pMuhbWS16XS6/fWU5trwnMsCinckp
lmN/3Abc0H5ALJWPAbGCrmnEzuOj19ib9FZ2wp4L00vCDx8p7Ifvo2cCntm8P78I
wuDBtHhI5XBTNnDTY68yG7QfrZkpxUXeBq7VM7899E62gCCJo+M+zyRwSBjZ5ttk
mKEGqtpHs6JzxOiCPW8FfV16aNZGSE+oepMrgXeB2scl3JSngGDQQUXG0v9EYOZk
KoodgvUPBX1cbuz2IzHrf7nWthz6hKYZ7N6X3OSbs15hIRfzlFrSP4ysylX8BN83
AMTN/Xbdl1jVOoOIDqUHv/5JBLRcU8T1O2lrEhhFK6ILu0pmKMgyLcC4/ZfRDUgl
iOo/L5owEmN1eqaHYkM6MK7zQL5uTZf6AEnaa8e4Ma/R/kZJgGbJoaNbYXGyDPMc
0fvgbRHYcdzBDvnsC2wwEuDc/7AO/xnREJ5m6uk96knYoOCVLDyuJ6kYUVMehAhl
a/wz/yi1GtMi6sYWfkScyg7tPvOJqS+NHuHoqFAg4+iobnDQjpYDj4GWhQcUMNKu
zfdKhngL+wekVZHRbiFxc5AAZXRnjBma3Z+PqD/Flm8mWr4Zur0V8ZirRt9x+yuw
zPRI+QG863lzXtTnagCbud37fV5zNix1z08UiEfAVh+VipQpAhU2zWWuOc7RY3ac
Q+xQ35HDDiEdtMGPaIi5JJKUFN8uTRG7vw6mZXRNUSu+XZeeoUPmOcR23qowIcbi
Of7zvs81QgblyZQijkx2KAHaYRs08BRgvhMNSuWy1ExAUHPU1wOKS66H2j8Fm+na
YuO1LuiVtqs+oA/QNfY0gBdlEO9Ke+4Yr0Y+MmItpn40SJIlRyTQ65RXw3wjuGRJ
YwHnLcOidF0IVpiuOcYLd6q/apJ7jDoKHZdWXQguVMcFFe3mkLIZKJfroKsoDmCP
wdp5yN3rt+SVf4oGgHVj1jQ7HCXHHSSwraQKGyHu6VoZnnQ4OrzdiP8mnCybga0H
PWqwVeQ7/SeC7UqvXhUrz+7VbMmv292vb8wswnh4xKYcKJ8Hh0O2Z2PtNF0XXEXy
p+rmFp6XW01AFLJ/PSwgLUeZ++24/6mWbNL3BsUEEgZ/LQlvU5OiXfKcfxBOSzqB
YoH2tbSwJVU50A3n1Aaup2aubkJvI1520YBYSNUze+xMP55OuFBz7xToB9p5JOTf
J3kG1Ld1hax2PqGdaP0QR81bXWgx3rHM6WKGDa6UmVD9LPtXfkMAIMyWOLbKB7bQ
cR6sa7ebZ0Su4URAMMhofwTmjtWW08SNIgV6XGyhuT95VxXG/pCs9JoOhAKCwWjR
ecMkPmEHWHwlJUpI/BfoWxDWamQUQyHmanIflxBP/79pGpM+9+6aopV2FW9Q81Za
/oaP/W+9UMmLehtw2eDKHUV85kqYFuSQv+A4CrVKwzkEXZCQDZ7+HgBW3hlhz/9c
8AI1G7fj9jkXAK9hUHRXLy/bJrIshaqpbaUslMELcoHrDr6xjVPWDXmijr+1RIhS
W/39yvbKx9dvkMrCuvUvvu6Kk/HVP/551Oz4Q/z+JbKQUXTx86pBqbgVLp7TMaBR
DIrzk1P7QTyBLG4bibJ4VzxWDDP5WvQrmSe0RzPdDz80PyjT6pQlkXXMO/oYtWVv
mjmpzbRYRnSr8+DpBYE961ZvwtSYo1TQ778jp6G6usMbreUVkA26KrpUYtrxr83Y
j2YaPVp/V0Ju/5huHTHYL7V/Q1o/1vjj6EB8zj5J1Lu/zZWj7HpEKGbiwbeJhoTE
kA6ffpStu2re0+8SUV6uvwEeOG1U2bP2rQPE05OZbwb5e38p33nmoB1nwmQSfNV2
v2oshLDxuZ8A1arfFnBi5laNX1/0VrhofNsUugWwd4I09SGr0XCa93pkYtFqU8vv
/l5riimdH+e//5q99UXEZevXAqUIStYmPN81NPt+/aeUBemoDvbfAPeyOCLbrepD
P8KOGb4T5pdInJRoEdHY1C3ScHBZRbYfTn9mDUdjI5W1rd21DXhrcXV26T+UHRGX
8MXiqLGTjGVd98rKnHqA5EU0ukebOQs9riycAgqNLQBFe/5oqT47cxheNFTOxW46
APUwv336LDUhZI44B/KhWs4QhR42k2fFOINkZ+MiGXWe4ZzAesStbkWmU+RizKsM
FIuzkOo7L4IyQL+N/LLLerPu3D23Z9ldh0pEkxcet8cRKVuU8kFU9wq6nhe7w6fO
hjh4nY+8Amn6Z5Qv+fZX2r+z3UtB9l7PqoYECf4YkDLAxYyRiUQrggQhuoGWFfP2
bi92jvypFQXRIT9SRYt6nC+CoIdVF5WVHzcmBBe0rLa/iQT5EzB7+73e3A4bDhez
GHlGBirXTBMa6K2BoF2h5xunvkBo9rra7AJV01+5YeRL7rt0t6rCjH+l4YdNRM+e
W/GwYsSxR1VZhskoyOS317g30h//CwFwFo3jQsAsJp8ucgnIra7/D+kf0/wTcI8u
H7/zzZG9u1OoRzoHjdWbcO8rw581GEvemzl6B7JIDN786gpzX89sw2GmZJf/1t0C
kZ0S94fIm9lknq0GLdDn2geWXtK/9Xdti7WuXu2ej0zyhdT9MTHPMOTtfMOd3d0x
pgBz44dO/7KyhQSteS9AymjGlSUDrDkpuREVXw8Vqh1uOheiv2Ufpe9aXqXgltA4
FcglGEpf2Kva92ZtxGCpNVKvx45cxe8BS6Wg964T8EkISZwTDBhz//cmgPrbOXB1
/6EjgRSVVBmzY0be2OdnGhoa/CASaCGrSQAC6LIW4d922NN6yUOPRHHcJmOmrx+n
Qj6pZH/zwUtwcEaq+SDDeHmlzeHGEtSHXl8jtbwQnz3ikIniTHlfSEOSx9KIQcSN
q0osMR0T1E1wr2LZupZBk2W4ticp6vUkuH5hNX65kZaruQVHJpbezwoOE5i4EZs6
3xtSc3rCX5/pf4T4PVs/QYa3q16ecoj+a4cj94H0lDnVy4DuaXZtXCEId8G5/vDk
m9KLSYJS2kA+nupUFSWbUWNLfNhwBcrkg9LzgImu9xtlaGDjSUqyuKhOpm7KHQ8A
0SctiW6AmbLMpbQGEsH3wGSW9/l2LfGpB2sKZeRMN2kq6KQeHSM09ss3sOQcXgA2
cv0ta6bzycnLkjH+ag2KRDpIhTmqysD35kb1yrC3BnqeMSXSAwvFQlcqkkt9AaF5
OswAllEY1WSa0LrthX/IuFp6Ywppv5OJxGcZFYzCSpBL5hFurfcmGHvM9aRPVt8h
EUoxFpQVAkc2oXOMGTfyk0t48XMe/IfAOmgugQLfRGOXLu1mr4KhTweq0F+Af19H
awA91G9bipTzQkZItcZ3nc8tkar5YYSqjLKgIftHtZzafR5Hg6bVuzr7jS6bK7HC
TNqks7ReleHKMU7mMnP61d2C0Fa0eisViHOhIh4tvudxQxim6PbquLrH4JrQvl2p
VMfedn49FxRzWR+6INhjN+cHIk7azfs2DP3J4272DvM4WEmVn+60msHnydgmSk74
mI9CUHKUol89kHTEUuEScSvX1dHXkicKg5lTEAaYQ125yjJq/LbU0rbmVoWIaNWe
MbJPTkA/Ln7XEYaEjmjaw/z1+UZEfo5vs7crGYcA1U893A2GjrrX/lvONt9OzIB/
nlaqu+m7LLkO7+pPoJadhk7aO75pQHnkeHzS8nzAZ1Pp4S8kA45v7kSRhkoptN9b
NbqGinAX2R6wRClq4eCiJKK9v5DTztbj/ftsP4/ZBwRrk1RBLreD6ABvOy4k0hzL
Il28p9N3UmNxTmUZ8wt0+t8VDWd3xRVmqKa337HlLi0PipKegsSSfpTMMmYXaGvY
TNS0WSUVyvR9FCdVEr8GpEy+TvBxJKWNlJ1cFGLj/SdBQOESCjHGqLSClLeA9r1I
a3ZhhjJf8PV/frpg1IUZsxpXqoyI/jZqZFCwnzEiDuUHhjjE7qdfWg8gBkemV82n
WDssOtI5Tam0poQv+GvCkELer92eHk6VxETxFxq0UM1QGkoPu/JZ1dBsJI9qZ/Pd
TicD9A4kDf5PBeT+fb3xeoCQR3jzUUOQjrnTg3192ZvFjzorVcJ7CKWausZ6C9I8
B1E1JVhItKxNezpTpTQto5aGtpfZRUK2m9x1VOw5t7bqsRscBlzFPhPpWXUQwNZd
3FDjVMcrZJLRa4eCyroALyLeqQwpuFJLz10xSBTR4/Na2cXSxWROT5w3uZuq/Jc/
676PyYir14gSjBVD+UzuMS9xuS+hHlx7tIVMETLNbsQRjXPSV0FmovnsYdAve2Iz
b+fwQVRnPxB+Cd/yRoBN9qDL8Vl2/dvxlrKNt9LK2dtA4Pet2+h+Ca/KDWOxi+m5
qf24cjStAwgrlWdkQnOHoyYyhQB4FE4lMhE6Zf0lv49FbIL/G8BJiYjNY7GFYUGD
S/h6SpDdRUjwMVP0Mm6PJ9vZbKCx94xWy7rvovhccBpH5Ni6btIep5brI1Ws0fTi
Vi/G1ZGUhEJqxLIBehLp17IpkKt7J1eXKs1VflIQZZ728gq/QsM3NEoe8VTBDExK
jwgElfcHvJGyLtw1SuylKbFf61CY1A8MKv1QJZcne9kUZdjBN5rS5kDDrRwp4Jlr
UwObKtHgaC7jVtOGN+3CO0O8xxNqo2jG/TtWfLsNp8KU/jLAMSL0fjZmMG61MEKt
AnrQWwNsY0OKeZgPJYhtQIK69qGP2s1FNEsJNZ+r8+yIwiowWBbcPbjska2tJwow
Pxi+pdwlLB8mRqzR0DNikqEwAA7LQpZIlGDCrlbczspZJG7oEvTfPTafksEzb6Iy
Mk8Hn2AI9m1j9nStunLB2FUT19jg8p56HyNh9ZIQo8SyHoC1yjc6ySI/VW/D2Z95
OwjgSnYwu3Wy28fh/MfYf5gZGexEGkd6lMPWS55bXY3PHURq+QvF0cTX9YILpR+V
iFKIM+IDjnKjv/Gk9vPZNYFDyFSGIjBQXyw97OKy3vBibR8dSPNQ8OUomazU7067
nFkUM8CxmEEH5bp/88jpQ1M4mNTjJ7sYssDnRotlLX7sUqI/An3eIFDnroljpkwn
5VYs8BSD5CKs+LXvz2DJ873uK7rVz8z03tf/AhHSCLQZPky7DGOS0GvAxmRxJY8P
ravCUbUhicenCrdd3C4zkWDNRGgXLMqmY6PaIVlYhnmrAJS8ogBYx1Jy/Uxa7bN5
w6p7eXZaX4her9wpIql1OQYOemt42Cew+dJ+oV7kguwnLl3oi3apbSyI4XEtVQ0h
y+0gQgAQYhSK1+uR7tVI2brKh7i+66jkwxTKCaBh076ArII2uwBIINKOvcdgUSsv
m1esAf8saG6zhrCTk4HSZxC8U0UXfd1yXzSR/g/sSBsDQB/i8j2ocVcxYrHDK7ez
j0tsr1lQE8d+c/67lE1kUIw8a7kzb79nBX8uTNlreRUyusO54/RYmLuO+28YzRmX
KgbhsX3T3JXfrYHFwBpICnq6FkTU1QzLPbuExnrJWvPhbGTQA2zNvNzRrFHgi+/D
JojojF9clxTD1DEdvIM+fICrOSWnxHdhLnHnU5hWs9uBOh1xFwjip05HsOeipdN2
0u1qaeRObiKUdr+I6TLTLriCqQNlbILyI5jrjyzYo+IQ8Rq3h+beojkWHMDz69/S
hhVjnt0VM02HFHbQtwtzY1hnvH93o1KZ3bYiSXMPedu7HaSTfyiCIBOfdHkBjhGt
S+h3qCQOnn42jGuLothafqWkd8N9A2H0bvYbFucdw6ZAkkSB+uizMN9Vf/Ach69B
fzLRUQgvBq5dyV4AqS7HZZpWKRqci2noBuVz/qYHhQ9SiqzLoLDwbygkcyHRNwcm
FtI/A1WIt1iNBCEHccgZ0DKGEU2t7Wccngqzm0DDeBrzctW8fkrUWGKJiPJpA2Jf
gZUs0QtZkuW/ystu1URa5UL3Wa2bC9zPiinetwG+ybu5JbynokijfHHZSH62f93h
bc4MBgYHi9yveGN4kPLEE3TzVpqg8tFMdwkJMD3y50wRMNhBBXwAzV4I5C678rJ+
eKWTYq4GQWw104N3E8tBLfKoMOz99bAZ5Kwoc+pek9pV7h0K5Awh394uNSNQq7je
Baxf9Q+biNwHe1jfQMXbr05h/7VcfhInNUhwl6bfoxFi+7FSwmi5DbHs+E9vPIW6
BoDx34sO5/6czrmPlezj+DCYZp9rtahk6wZSgGchYieonYelkCVgxf8TUNqSOqiT
pELQZgYgBgvleQ3V7BV0ttFsS4qK2dAstWXrJ2p55RZtSCD1rq9AyyM+UJPcwerY
S/RalKCPQFFfPHKnjUf/8JPoa5pp7X1CF4SneDq91ng8iCI/VZZNf5DYolZYHf31
/n9SO+rKb9+NCQqrByTOn+jrl6Eub838b/6SC/A3/vhelI3XWG3HGzYCVRPgpqEd
8rKewXoJ+bS7KNn57epMM/Qbq3MTeqYbtyeTTdH4D18SAm5IBC2au6Zz3iNB+7Ja
I1Ic1+MoBddZotz7cYy4lkKlfTxFtG9JgGsH5sRWefhyzVpeKsdmw09V56lm0L8L
Yx+Ai7JeOQ2ytNL3u+vE0cY0SquRJ91AwXNhtDQw6Jjm+OYODz4fKXP88LdMyGPz
catBVGcNB9kTmpxt1aGDuHoLIxm6vBHORxOjsiKe7awv6SBcdKuK3ZmI0UJlXq6W
I/irSsI5ixZ+kBEQeXKV+/GtmER1KE8zGkZvN6gABrTDTyPUi+DVuEagslL0mNav
juIZ0GGKl3GQQybw+Ks0HXTR6k0ZtkF+jFoGkLxH0BxrwC2Tuk2kKw8xlJCKsAHE
vY6MczpPa6GpeNwhRxIIOzw9foMXeZ9pQgDEuBL9dupPMwjBels2+8864cEO/jf0
b4t3lMQsIKBNtqQGeZ7PaDJpzzh7HOuffmTeJVa8kvRXhavukrXPR30iOL2G+J4c
f/JS+7E+l26OWLb0D26R8efxA15E0Rn0Xy+MTQcfIhXlqT1X4BgRmfcFe97cZCko
VDNqtvdO2AP/l/uhYOKDDdwxi4PJyEp1o9ylF5I0YEiqd+IPzlQ5nEJYhdI7RerT
aIGPwWWxoLgPBGIkZ5AOKLbcSX9EkXdYySkDcPWVvDJfG0UP9mz2gSmq1wLp4uPA
8jeqF/Od5P91POVaaktMBEVOtlBhc1vp6BXqHtL+2SnedAvlJonpK0XPOv1+SHdy
LZW73j+fCK0esl5Bd+RJf4+NECoWhmkkolnCbFK72Ue3Y/056nUps3jz2Zl8LRCO
wjWh8XvEyJWSdeVE4TmqHaxHKr5DZ8jPUWpJcIEV99l9DVpfM1dFkILu1WDk6Un6
51NBrSN7fQszWXZ6uX84dN4SQtyz6Ra40qQ6oWMeU0eHl+g1318Q21CqTgwccuaJ
pA0jGrlcD9HMTnq70nnwsYsDcSzQzTAErVutUWh8boa8Xl9ts40m3tIQ6U7DJ/E7
ZT6ObSaOWm2UseLuzGXMnH5mAGEmoFxl6ZQE8lZUk+pjTTqJ0HAH/IvBGDOrP2L4
YHrFa8U2Xo23dR3q1eT1jP5bKR0ymHXE74qwyfvUV/+V+c0Xto6y5VopXDzXySE/
5UrkGjrnxZr+8UMrVh3rLe6RGNJ9N4DvCCtRCQ51oPBNO1EDwiilgSxrSyXI/mWo
PF26uqQJetBNBO+Jsqu7UBGkHyqb/aAgXgF3nLRaGxvrXog/3t1Tm/qf7EPRgcM1
slQe5Kv22PBByDLyFKLypnn1bSXLE58KWKQ4YrpluMKwgdHw6RSdwHUwlXywkUc8
3ux541DIJsdpjmhvDF5in7LQaiYZe4CYc3XZpkv6dOrMl3hDjWhWU6UWei6lqepQ
TpBA1ZfgvSQqWw+hwz1jJiA/Jn8P3najtMSXQYLQPn0xIJ5fduWqXfNaprGlRTPy
aKPBNVvsvu6ZJlz7N5mnDgs2A78lpxeGNV94FiJjXvVNCAFxDgL5urzGaLEx/3Qg
8FRpE6yqedpuzUsbsffTQRf6YKmGjCPp6XvdoRyBfOLwzKUboX6x6EsazheSj+Xp
LXTGOHZjwHNc/S8u7IKsep11tU7qfru+wnQGa0+Bsf2KxAS4PmwZbeswigA0nPHF
O2Z7rxRIv4GSo6Cbi1siMm8yL2aE6S/rghkXG4uk0zpac5X6vkFrmHX5IySHmqor
SgsV+tz1Ov0hlC0V6Ph0m+wdVPvjvOJ33PBMlbhfPlejoXQPGcF0l3Tlcn3qUC2M
dsh8BG9pTIITFl/tMBPZkLN5o1TPadzav5V7IOsfl6C4VDcSXF6xv7nPAT7XJviv
V+U8LIGypNF0spekmO4P226Ee7hsmWmdk+C9v9D4q8aAqZAt6j4h/+1uyxdClflZ
VThiVeCqanFqDeeE4dHHmM9BbyMqLPAQBVvfVH+JBgQqaO9ryYt/Tj+oMmT1rYSj
gh24/AhLVcMGTIhOyPNbQTBtTPpQfeDt4IfJuq/pcsHLpy30aDh1cgT9PqZDQjPF
gwHrOVWAMGkcIRsfEzGBqou1JUnnQajvSEqh6uUsT2qEya8uA89GW9cOGRtApllk
RHmRfMzzKC1y/SngbbCXhw/Mg0HwfyNJyCm+ODNNPxpX7dpessxt2rowVT8N1Rsh
aZ0h22Y3FpeXAhXIaawwflQvfBc/eL2g/jKM3CNuiBRvTuejXalkXFLm794Euc4K
R4vN1aTnP98faIPRfrMq61SvcQYHsm72efu/TlPxu/fHARctYHFH78j3Ew+LMn66
ORekPBuqC7xW540uBjRID0EmlKr3Dn6VFJUOimSgZHY/FmFlsOO95QUt1bIECai7
Ew+WJXcS5/KBsYqT3QMh1Qz1c1HZGXKuw40Zcnd+SmaI1deUw6+4IJ5nWTAw4dNI
Lx40R+a3ZLHjqxG6yXkbn9rdV2MH2o/fxdWf5FC0ZKfmDyyDSgL2G4GFGAQaPIwy
OE+PshrGtY6JmJOGybZ6M+6RqriGjzKjx10Ol6t8orDKz/k8ubse1xZHFZe1A9Cp
5xBur3KA+g975cQuTxxPHqS+jypCQAUJk5xjiH7SJgMV00jmmSj3+53Ju3LZIjlQ
9hQmaGCuopflHfloJ92UE3pqjlgazW9opJ0ge0RxhFnIn2RW8p9aUJp8dJcs5TDf
SgsHst1mGfdCGOWVCa/WZUJGMAutUdygFy/I+PlaLzJs/NV6ep2orrQfizWmpZBm
l+gFedBUmIBRL9/Fsdps+NMycCgj4Yp8s6t6QgWlMF3IT/9QB+HD/6BjscAZJ9A5
fFFcuiGurzS/NzCk48dWR/4no9RYSvaM9+PLG6egD8GHDDSZZNVHnj/EsrT6fod9
JBMWO6uNEVmNqCaR85P9j1DP+Mgj2uItIeioUgG0ZcxkbdNN6V5NCqqWqQIC/pQI
w74P0f5X/Vc5Mny+DrjcwEgF8/QVPz8CDAtFHx4j9TxQI9MJw/OlKUqxAM7cywhM
tt2K6uEj1vz8CHEthI2s4yxUZzFQM2pxeJetNXNHSiY0KSBwjEMr1AhsCg1eTY2R
ipC3FN9PqPqOEYWd7RNGESwJnQaoUgKmXhL8RS+0LDJTP31aiXIauUU2D4nYRiUE
kO6DUhzzu5/PLHgZTVH/WmCf5jFA9OVqxkm+T4vxL4g7pIiAEAlG525+w505aX6r
69GrqH1bU2lKUmD8kLR9H1hDyq2W8QGvLGa6DOe2hTnPPcsrQmKbR6GYJCcjfXT5
zz+0SwJSHmMFf7rPzLyDNl/mXpgaqKgGaczpevFEbkzxGX0k6N96NGLRqyk2D3RJ
dreRbykWGruyobg6HuyryQo4lHXiA7xtgWvzpk0t1soCj/5Sermk3yxr0Bs1430S
4hwVO5KXMqKAhdT80MHKzQn9kUDJoGUWrwinzoZN+MbLLwGohMTbqVP/cFdKxSFY
HC2NEoZUsLoyM41SeC/0+YWxuyLADcDH6WT0XfrawZW7DU3IKPj5nT+Trp+7zYll
eOBcrLWFS5dsu8NSDclxFpAENQZr8kH9P8dPB3YFgg1+AHpD/kQ1ay8CTx+msKWv
ac9Zdu9eWXfsdsXqilrvu549Xgd8/68taIZgWHVcPM06j8xc7qgWaz5nOPb1Fj1B
vP7RefSRX8KuwdIvqccsHCsUYo25ZNdd7ixwq21/L6rXCj8e/T+hBAoGbt06CrYt
Or2+7ogxpz2K+QZ2dy3ZY7DHfJdeI69X15f2ZRs4OMNyCi78ZnbBAWyjw7RTWrjP
XggoCoOPHpjrS467qezskxHIhk7Chq0+5IlNOx1AzrVog0kbbWomAfOPPAQjIPb9
YhRDYcCWtt7kMn1JaNPNMOQ/I23FbckoatYm7BNjBnkPjS+XwbbIXhZJJSh458K0
OMJTjmxh3YBw0MAj6qsZBgJecAC5kZ4TjxmOj6VZ2Rm1QTLbmikjKZZLhUutz/k7
HeUgTebCxHgrOc+yVBzEtdCBqzle66BCguRs/zPvw+otQgWQwKkAffSS8eidH9MA
fGeyKpZ/qUpfCoM0DoFZ8Fcd3cCTh5fnsA9q7xo2ji8pWX+oeDL1exFzzQ2Rcxsf
C3AJ9c/1S6r1tudxVatS7ffd5caB5htwifZoqwBwgTc1muTfpCQo0SuLSyaQ9nqh
sXjOk8o972oFPp1L4UGErrcGtALvrIluWt1jXjLAetQ6u+Py172FcUm0Rx3bBurl
gQLUZpUaUSkvYFwTF28/38GahiaVU08rau1zbI85tOp/NgO9UaIFF1KFoto/TVmi
3/rT4vU4eV+YtKwxni02+kNGFGAkkuzpHTsjEOsp+oEkUzoxLhG1lJw9a1CzawUW
OgoAAsRubEqkngcbtEihvUoHPIltbw8TLXIMuoxfjGy487KZ3eze8ySWqnPCAgZ9
inYWviZpvyyd51lDvmvKos3ckIpf/dzxKY1JqCsmc01aVxXS2QESh0AYFNgws+pq
oyCesSRd3DIMPJ8K2rQl/HYsmO8EKozOyob4kAKHp6ldGy6S7Tuv4mxwy/QIs4hF
kPzk+7zR64NCMOD9HZBC85H3yFV9fvZpG7DUjrN2pilby5Y4fxCtSs5YcYCKd6T7
PE2ltrJlRJotp23LF9lyGv2gesP7WypjL1YnwT/Ivcnc61nct1iyUK+lO3vesWsz
907oGXdaUBIbtFW0vinRL678QMCzcbdFMy8OrFD/kg1rTj/3hF/A+BtWvzuJ4c3/
ZmE5zl3qhTrhQsuSOGPYBhrOFZnRNG+T0t1Fei0iC/+siDBtKbIdmUFPZykhJ/SS
HmbyMhQ3wbR/qzEcWH7d5QB7c3/PMWXzn5HLzoTJKRKsSmKWwMjwgOXAr5e+7F2p
0T/1YIMW/w5fv/rEARilf5on9t3spzhwtJLIREZFJSdU4FcbFv0t6abgbzAQ4OPi
M+hOTdFMkUSU8vJ08y9oePtGFfYwLforZkH5WZ68XV0P/xhGo+2mXjD1us/5bcG5
bfEXtWs+vEpx2coYTWBA5YGgMgFZfzC5V7XZsXma/DUN5oGQyPjYnwS8t6JK8oUy
sHZG9f7dQA3H7LeIzVRggDPOkFKgbLl44xHvNe+BZ8hDS5tRg68iFRKBTDOJfb9p
LVhlchKFm0l12tsTj25hcCFnOR7apZQhjV2lb4GzIj+70T5vwxV4QfHugS1gCY4e
CH7N0PBDZ41HU6X0IJ6rwdJf6X4JghvZQ72cJTZu4JNiy/ZjTvkCAXUPrF4kIYMs
N/w/RwynaSyrz4uW8B6R68n8XEMSE3rxNS7WkfWj8hyjyli3aP4W2dIyqBHjKfEP
iW8unHkxmvyjTGlMyjHgXf0Bx7vaauaj2lFmKmDjhBPJEvfbrwLiNXO7z6A2zX3l
ALMdla/ZRDcU8mZfTv2EB5kZB8ZRvKyXomx8dL3eFW1YZgf/Edn+iGE2Ysc5tAFf
9sm444qHY2D4yoPTlEQQ/0CrKyNDrIN6esKe2s/9/X1x+Pm0H0sgpLVXhtMvjC2B
qA05QtrM8xofrFG3DqhSsm53ciC/8LFEnR9f7h5q+uY/Rld05lgNphGhh9FgGaY9
cbY5LI4uof7vz1QDydK+kh6JkUlV1N3RYTjMgD+5L4yRlh9ZnfzsAwRLG66ao6x3
uZQPZGY+4gveMGV2EtJAZw0+mfYQ8kyZk/TTQQzPV/URBkCWAk2h/0YrWcwY796N
GbnSOgzUabvEzYqUCBgJGHrLnfZrjBMOSnotkIRstnsPUFVVWc9ALdunwn9ZPSGQ
8eBx7dbn4YmiY8AY4v3soBBklwmmsEpbYWZT+rjYpX5LhvXsN1ZTBkfe5YdU/ZAS
y4cjSzDiIJi0HzTi0p3wfG1lquo6/0uIh3bwF3CIGN//dmGv9k2/JjI6Gf/PwVZM
4uUpJaACMkFL74jq6KgFVFLnwW9ZZOgpt3jsRNMyV8FkCVDg8HzjOSlcxhcbtGFr
Ag0e/LZKhud8AOZuA5SZCjldLo8U1l7ClWVqxFc85VVsaMtPcuaJdFaIlPzf8tPS
wvNOVKiK+Df01XwzWkm5JB0uyVFY3MBpCFCi91To6RdL8r3VyOYpDxWfJUbxDlAO
ATUJIwzM7wRf2hA37zYn7I0RsPxaIwVlggiPah3Ta+fI0IQ1g4RfjNaNmogQF0ja
USpzJVl4AaGpcPqHUQP3RVqV7V2D1xwln1UIRvercTzrypuUM74XW2fYCZBT0fer
u15Jua9pXiW/v8mUoQW1+eybQRZ003vAfWBSs32Q6WXpeU4vp+jevKtVmdqFJnP+
OLyd0mRbsidtRBlhcT+bZpDVkFqA9yhGBAaT6Yug88118hgU0eFwHNlPpDIC8z2q
xTZzOTH/4FYY4+O7tRzBwQKXek6rDXNMRvrU9dadl4o/0oCb05mzcwIJgT3B+Au2
8QTcaJ6/So3UPuJPOEg3F6+AUv8PySweO0snQCTep2ngUAuI7ffCNM1SrVQ/gLbP
1bjYDAuhVPy0DxOixpPgFVXkbz9OzVlnccmeAE6PYigzWFlusvO+xwBdci9yXM/C
rVKtpoqaR6vhVREw0HhReadKjuIrsY6jZ8ekkWApAS8MFErFd9JCzTvA8dhjNpik
I8wUSJvKtAGLl9OorAHO5q9ou1SGXVx5oL544qNF3LBIcyzY+JSR3LG0sKQTpsNO
y/L1zLDrueczFWlUc2Pkr/uxbR0wQXPs2mSvLdBQ1YJF8xzBNab98zUqQqfNv478
HmhzhLog1zLuaL8VjHVMhmkPmJDIaSB2IzpD0sIoSKt+e1xLgTTGzGuaAkUadrIz
qj+HCHTtaHuiPoT9QKWrKsM789hiMLJAuEPJk9LQo3hEhyJkGywrf8pqz7vDPmQT
oVOeExfK/39iwwZtWxWyHIvr5j9iS3c+1JPZ+5vw1nKllAPLzGnJcziTjOIo9Ycl
r6Zayms9dGfIgszrdPu01Lu9etp18XSBZJ9h+1xpOkkjTfW/ovuJbwYz/53zGVYV
GvvHi6YkByBx0RokC/MtconiCRtY0mL0gUA6vkwIgnFtIkp2tS4eNEAPwpo5sRef
JYF9zr9Cye1t+JCm1fjgQoU1aXfYjOoVgGjMBM6m7/fOOs2tvKlYUoRiyvrvQvIC
WmwwsmzryBV297HDoAxtKNeWrsz+HuXc8of6yVdf44sw6U+q8RZ6awRGkGO/o95F
QJEVcO5dJSwjTv3BWvyj1Egurkzrn5aKQY7vhkSwBLz+6JbuiLy59+OI5c3MwVdm
BEVmfUlhPAegWoMvLCTzG00O0mVnKY3wmRo9YlbqIPVe7l10ArWBJJloBq2pxsBe
lYiqwwSVcGfsuElIHm3WNo70rUMeJJS8bBA1OfauFPgYsO1xFUX3KZfdW/AASPr+
DaT1mdmO0j/aP5B0vKdzncMxFuJ+eXywc5hrA7f0vi2CpVW2v2e3JOsbH+4ckbQw
7bZP9kM939y2TPqM1TKRUpRVO0Ku55pVLqOJBS6Z9G8BgnouDuE5QKFyKsX4U4ic
yCt7ln9sRFaSYztX94fRRP6bw8DYyRy3rRKf8gw7gaIjV7BrMyI2nWgo+Dc3J8Ay
x993UaDg0ktoo4ujqvCTE3Sfuw5z/YlKnMeFTP6CtwuDJ7dplS800YtS3uq37FDf
3+UsoDUazpxLv14EzqNKKctzoohPwzoaRDJhZhxG1rSPq+hIVVlsvVbYLqz0RTRN
wAzvMPnKHfdnQIsmvoMYwL4/PtX0550wW6zhAGrZSfcjIRY17oWLRXUE0K1YTCbD
w8Ko88zVb6aUD/vP7wHvIl5W6xEOuWeMdk4M0odNDtVf9zxZN1Wb0abNagWp40zp
uN4SH8L5cGhgTCPqKDrfelsgzTqh4/AQaYgrUsi9zhhGddu8NSns+MGZazZALRx3
n0PyBJyuDC4hm8Pqbd2GBlYMXQHnsBRykt04CGAhOA5kF62Xo8OrMObtSdDl1DKH
UHPDsE8ezTlHYKqDj/ZF8/CT2csqqk0yZeGlfAv6omACEFf8w3yqp6tvbNuDiv70
IldPeMkDdNP2NRkiE/eUwqT2xHtEPsOrrecBHXJk4AmaS6+mgmtuQLl1sbUjFaYe
yA0qebjyQxEapXxLO2zp0Q2ZyWmZ2BnUjhJ8gX1+KJNT+/+b91KFJWJrDFTUVQIk
s9Fa52XsZoNZ0glAoNKPBJcT+kmyhu9ybu9O0RzRT3YttlSAXfV379229mhdzmx1
TcKmX5Ir0eU1vzOlEGhZBgKIul+oDsKq357YiCe3Oo0WtJ8KUqOx85llDC0QTu+h
EbAD4kbP17WSEjcOLovpJ9SmPeZKB+rfIk5o6/d3Z1s4WsRTmJ7rwka4u1jKUK69
xyUXlKg3CZgTNpAwdEBak3W1PlyFvDpqllZuO10i486gTF3u5ay3mWfO3jMYhqi0
P4ue1/1cA1YPsD0EP1bAcmVuCAf4xGyk17Hp4ZaP09z7Pb+n6VbPdVqyCkEWYSWE
RyFwOYfwInIBgPfT/u8OymvGW3Y/ch7V7KOSK9kXeUOUyAIHINItxhGuyddo9tGU
V2U5siCNakgxSsb8kqUvQeWc58nXBOlJoLQuvzZ0LyXXO0bZMmcyVjO5Z826LROV
FJ3q9vGffUJC2o63Eg46HxisJM+NqQuhokoJwUxQ+z8wS6T85sHv83vOV56Yf3f+
wgn9H3Kj7EJ+jkJdDHpQJLTR8xCRv27UROiiUeM0HKXMYWzfmhXr0UepSmPCuCKV
qdcGzMwnIXHoilMRXnw6UHZ6fgicnrgOIB39jci7Z6VHY08Ow2VIG0TJK2gYhVv4
Ffw/vjQ7xap83/QEQ/9qLlfLVrsD3O8wn8MrFggeMIJM/1uERIuTbUs+UcRP89Lq
G7dYZYSfHtzfAXGD9DYk+Ex41oPoSXde9bvKOQ5Z0oSDnfVUVBoshSOMmPcZq1u1
OUe8nA/0jvdDFy13uPKdr+48CZTB9E0vrXLdwvlIJnpT/0BJE7VK4LHDXnxvdjo0
pYCaXjWSHKBHK09dOMKxcQ/+7IzfP4GcA4AaWy1q11hMl7P5/TkDd2qwg+xMv6x4
ONyqq8siBucRpCHN3efDShZHV13g7+X+me3ubBeHkOgdDmUCM2aJ3bMuaHOCX/6e
RjhaR6KtW69+TiUGQhOeEy5tlkbPocap2pjosso2yzZfRWASRxbknbFjt9AKvXw0
1xGRcVqozf2SN27FwUw8ztdri5GWrgXn11XgyWKgpp9aBuPwjMTkMSg7iqGIyjNy
zmWkqnIumJ5YZnCiIwI3D6YN2EA0szKc+D7naC/4QvGKi8wVEbKfo/gSgZueMbY7
AftdGy0YI+9rYT7/RuQUc6xao5irrlZaWyvnBY+JELJJEvQ79XlHOrE1McolqKA1
joaoOlYh81Y3+cyWbVQkAPgMmUDBkG1EN7qbHhcSOSgXh9AfKz4IrWZCebUEEcp/
9fSi0qGwWtK+jXxkR2+rr5evnexqVlzXpAY8pyAAw6COuIBonmvcAkkBDNwLR3/P
Ycg4IHUCfpMvVJX158QQ2i5mXOZ8sCIg5U6LwToD8i7RrRn82op38pkpWJh3vsLs
VsLmE/Y6Gypcokt/TJ+7VDysPDLGRq8Rn+mJxqyusVVs+N/oG9a5mrtGmTZ6o6Gi
pDpyaMrCMqR96R966XlzzO+I5h68BGL4zP25YjpIoPuE+vBA4p5rkDxBsHPvQ/FD
GOIvX6SKxtlWkBgSOGTkwukVU9eAZ6PbSgupL6eNKAwC+bZ0gZXELrlWS4/EOZn8
ZCMtRhojsojzE+7dDrSIRK1lSpFjf3WkU1qz6ndjIcfjPtjh2tG0Or2SpoAEyT0O
LQePWK2wvj7JxuvAqwB7q9vmwp+z+JGn9NNDZdWDmg6kln8X6cZjGHJ5wRdZyVlg
ZtnXDytOhtIhSmcxKeLCmIt+Q+RnR1H/pXSbPEIuxf6mFKUnu4beNi1EBd0dTQ+o
8QLvdJx2C/uAqer2RmXrnr8pS2JciatzFNlE4iKOAWb/5gATsyzqhdIbOrFW3J+d
B0WRib/Z/0gbnPkTGBMJ1tRkA60dCMSOcOAZ775hmv4NTuXycmZIDyF1QWzTq2AN
sfltmg+PYWTuwmLK53ir0a0BDpMsJA6eKxVHtRZANuSbF/+5MQXNR+5SEoIl+Hlb
WmGeB35fJU0FGyRhdxR3IghO8+tvhLeHeq5yC2ligTaceeTJa2dmiBINkfi5K7zr
7kpNM0SE9KiMFJxbrw97kXpWn3d/bndAojjimNubJzhBqnWZoSApwFFn5bRvPRwM
kH+lTAMqbnVhe0QlUalcDxV0rPgTFBeaCDYKmdGseGxzqjkgokhhXFSUKDWlufyC
yivrFRjZBy8zWIFgBMy6UopKIOc0vy/QGwj/mOaPqMTdJqJ1w7iu5UMx1OYSNTYx
3aTGAEr5ML9My8UhF3Rt+Zm5PLN3rQB6NVY7vj1iUYnWwf2gwb0UtwWiSvJVV8k+
Pce8QQ/k/fQOgxulCJSfLRAz41QzDO8B4+251Herh1RktKV4vADXyP4Nybi03ra6
Xu6dFWP+g/xk5frNJdHXdeoyAH2srMpOXpZBwyYzKZuEmRAKC47QxEuV1clbK0hK
ouvjNkaPlp0xzKmFFXZfyFFdJ+lo8wmq04OQa3MCIjE+WIsvSEYjCIey5wwIfMwW
CLm+vV3CVLAf0V3b9UAt1DhnoFICaXI7nXyth1bPenruRgJVOkanEtZ3t9Tf8M7/
NBUrC46jedUf8ZWJDVf+2omAjUXHAJYmfdiuGTbtGL5e6PRVtKnxZcm91cm+4amv
FuiG0+RNxAtvvBhsfhtqxkvgH/EIh76EGk6FOE6uO4tPqUCNsASCUt4j+COa0KVg
UnT6I6L84/WtGZ4K0eMYLmKYcUMOnqG4YMjnKQMlVk79ySPtRQtdh1WSYqX4U5m2
iInEKt1WbOeIkkSd0nhp65SDQsVnrcP+n987nizN8NFNEsjN8K8jBn/RJnezddee
aiPaF/8vEmtgJXBUj7es3SI9W+HpiTp72n8LfTxWO3FRVe1J7fgccT4tN/TawxU7
Yz/tkDshuK9luIEk+/kxx8u7dxBO7dKI1uxLun9NL3dhDjMWQk/+97hyfhKzzDfr
LA+qr8PmYZDVuzCWIH770iRmCscyvwfe5FSwKHQOVTwhLusvR7drgWOOsHjHj8sj
jy7olGLFOgqQyDSnNkOJ5Cm1RvJ4lkKCFu7VOk7kiNzFYLKx79zuNSXr1HA3ykf5
Y4TB965+3oqJ49n4BTRXSuKje84jAHmcOhR6sfrBkLpIIEPPKkuXAmA8dLiUrIdt
13TJ+nKCufPzcymqksHEpYxbU01LHfwL8tHUragQsNlah3lZONHtCwnwZnvWkEKN
qq0x17uibLGkweSIOLY6XNLeFbWJo7DY6BoXZOdigkiXuq/ZyXPQR4E+RaafrFae
Kq4wyqtPDUtJXKb68spPk/VRMNLC2+EF84bhXHaUIr7k0Kohc7LepNt+PHET/TcE
kS1pwdOtSaohwikHj9mHt3MlbZLSuztntnEeEiJi+/gf9Fr+s2SJ9Am9oO4X2+fb
1fVCEoxLBPMvvuxG+JYlhUnhYnn9k1lJk9iJpz3P/LydEL/QlPHYy6K8+p/ULCas
HQXmX+vgL/aUJimzudgiO/zW1meeKS2PDPhX4NAmO82l4hLOKECeKGP6rg9KNq8w
5QFle/MrRjeNosJxeIVEqDi4YobvJTZMddivGpH8j+qekF6ZIR1tr9fse3hHx6PT
SmlhbU2ZeNVy3vNAHvdrsHgqrjVcKW5e+VBbPgFxMoa5WfCEjY03AmkEBAU2qUKO
aAPny4jw6FHsSgLbN/WV9yS0L8xC/Y++D4Z0dxflv2dNnPmWtIWjdJFcnForHM5R
MEDio+mOtmY1cuB/ivyg3lRR84rAVGYE/SFzpoOfxp4CFod+LoUezhMiUQtznpGO
61lEckAZ3SlDPPdtXUTl7XeRDBMA32LA9xT1KIY9zVml2Pbr/9qllm47zpt4IwIa
stOWvja4+5n0sgaHylgP/HpRpOOSLLvpPKI+Va1ILqQppGngYRiWo2LP8eQ8kjmi
ZSLvZqiNM2M6Y3a/YCYfRzWOFgPA+zcolkgcYUR+jGz7zQHicTVU6eH/e/NpyBt2
QmCIrM8klIis5mQ6kMFkPknxV4noBbOrBFyV6IqDf1Tyj/kbcjTAXVMCpn/8Rx9v
oWy4V7faweRwNhNwmnZx/KkpTtFUG4wJ6yZ7/Fw5L3wTeAEEPd6QAiYSdOJtQ9T/
T5o2gh1Tk/W3AvtSAHWpp5LgHMiX36eCFd9cpSbmcFzrjFX1GTE1nj2xyQfB8nz1
qPGXz5j3thUZ7tI9NEHj8EpxSittw5A7NBg2PzEtVI00BM5nwl9hDjYTSA+N7F3A
uttSki82UX81iL1tiRtzc80monJNDhwprItEEEGqNu6a50AAC098haZj6y0vX2My
RxiO/nkWStvp0oEniFosVdthnyXf+aQ0ZuTucYI1zTzFqRy1rTEYz/NC+YQnBqaP
wworrgu4l6QkUBydkOUm3iAMn0Umx/PcvxqcKRArpHkLl/eD/UJOa3cVZxHx3udt
ew0PoFJRri0PzEoPGEZIjpm4+MIXFsCXKIXe8ZMru7EWvA4LuilMsYiedVxFkliR
vroVqR2mcyz6//hLC6ipiW9WWz9D3V2ItiOMUgjDUvhiOZJfCQchTx2bW44OTUvL
F/BsuEKAFHEk27IhzZL9jnHgvfF7MopWJnmZxlYR6xltbmEfSoAcqn1YZsnKlhe1
CDwq2FfbwmHO3CQ2U++AXOxD0dBGL/2ccgojvTQaW4WHWwcqOkuvjTU+jWnpm2dP
8oPOcWqjMsUaEKpC3dttb0Jg0YFd82OOPKQp/Ay1JIt1VogPealcGpYINgXLMm7J
M6L0NYysQF5kNmsBm5dSWI/K0pnKsX3qSHiDsibwRBvvitwNfJYwLetPOnSVmnjd
6R3EReYV04yDBwrupYEpLA35EuVP35zGMC10lLeW1mqitqJ9UtSBdG1NxiDlKoEx
lMy22/l8XvXu0oV3j1b2Yk64aR3Z+buJ7tFA04jVlo7QO0WTICYmjihiTF+OKgro
ulEtSa5bm9jv/cnd4BJncZnIWgPuErGTWCj/SWrNYKsQBofnvmFcxFSKY9N3RJ8u
PJ/f+PilM6oHUZN8ddpmlK85ap+/NQNg2KrTqboSmpuQaHeEZUxkORWV4F3TUmRB
OIaXz+QM62LWLLL9pZDOpYGbgMkmSdEBcB28nBqkEdx14h4rSJMB6n841RwJhadm
WJECkvCy/BRCNuuI7Uv2IKX6SzmgYN387a8iK2pLfoN2tlXAO8IKbdvymjBc3aeJ
RDQIALDezurQK/K/s4WapAOwmQNWDADJr8H7cDBG9P1kjZ0rLBGxlc+6GwZtHUTC
Y0XetfcT4yn3ay9Ae/d5+X07Sjd2b8HEvm1ukvUr3Ur66RKaZf0hNkCz4QnhCVBG
+w75gV1Tqr42Zc6s+squvrKLdxHlvA2r8dG7sSewuutRzRpL3bLEj7JBq6HBknSp
9wng7sSma3JZX//fKU7/a4YbovEfFd1Qm7MPVUJAVvi6l/Fx9trtRjZDGN12vzuR
J+LkNnl7VdFNtbQ0qxi5eJjwVwD5jbhWkU7LpiGKrP884UTYtwj5xjd1prOYVkPb
OM0gImhSdZhvSJO5Lu2TRTktbReLy8N7+7PAMlVoevtsoxBRP8DjEMplAP6FwFJN
ltTxUZeKJKdA81yHyEA6YziGmi8eEk2bA6bjl6kG8Uw+ggkscDWyoalk78MptpMz
c8O42tjFY3vyWaD31iqfcaUBdfXDJvzuYvYPfAul3N8POWoB3XwM2j9YzsSMW59o
YRDlkU9wqVfROu8Lmorq4sD3Xb5xKP4UiNGpxUsYnDXGzHDjJUGq88cUmBse2nFV
i8t4LzZ4imtkpdhChzgAoIpqW8fvbb5NmDLes80v5hFRXfVqMyEhjWHCdUjFkh0j
9HAluuBUBlajd8ySmfmqrHsoHPAWnKilbvouceD4KjBn+R6Xpm5LrcW5Xs6R0w1X
rijAYu2FQGSOuxm+gMpZq2k6IjfqLSrZ1LJ4mCI4GMqgWlB9+hk+fW4U/d2XmpVx
KKy0Ds8C/EmRo0/hrs2DxKSlgH5pfTMM6PjzwRZ7LlD+uRBsco7eYiK/rH2h+zDl
/Kp6km1dDQ0/8NYUpFPWq6RIOzCyp9ILh4vuM2nbVJdpfaWyOzOdSNWX8zpSmxIX
jGbhfSvMBTLf1Y/vdYFl54NNVpAkg6ddebqGUqB5uTWkk1epIreXPj8Y2kasv19Q
8IValOlwKlH5vKuE7QxWST/bhpD3pUM+yuO7XjZ4FJmAgPxhXLsgEk0IfTRqKB2R
TlOVgSpGfz02mE532qAVySseNh/XCH5tLNakdI6vEEhsDNCM7M1ZPyT1EFoHkl1K
kFjm9xzpJg1g55PwKExAof7a4anaMwC9gTGiyhNJIgLLpUE2pTpM4KHIYFsjiBgj
YxCwtEUtuDDhsT1L7cY6G4yO9Jrl4gCEdVHWbNSoYlKlSX7BXGySDjFfRzmaT3Y/
5flVpU/gKuMflFu5sr9QBgVC7EbfTm2cFTUpVZ6CTc0H00qL64JFdnStLHsfW3TK
5sJRft62oNiCaLdgL0z92eCxwQbgz0wsIDTJXWqHwjZD9bRCsqwA05oANjtFevww
rdbhkHDW6e6Jq4bRLC7K4OjK7dTyoP3jZiwdQXmOpylMDaEHinqHUpq9mHoUxSyR
umHoYXIreX2o7ouWsBoI/0S/3ll+vvmiToLPinhr/jNC5v1lBRrycuccHUwuIwe/
RDYRdIJ0CyTNok3bxsETLnIQDayuxhYJghJm18KtN+tQ7F242tws089zjPuXkJ9a
bh7sSTy0oeKVTcaVsZtjFJkPHYqWWXgFOMXOT4jD8hQ8aSsJJakjkrZOrPQu3TVv
ZW9AjDwyE9cLi4aKy54saH6bNxQQUN2o+f/20imAeIMRCbR+Ljbwk16VYLU6Vxdz
OytVlJl6x5xPB5uR2r3FDmPWNHAtGVqw511k2gVZyz68nkrSdx79z+ZKldTb1xYh
SZpAz7gtuU0GHyNofKFKazGBRx65J0UsR7LBvT8Hj5/agRf0sAgInXqE4CrH47Y/
qhtqaDKQuLZUDQ4cH3kQKDYgkD0BTQEzxdCVSsDMtIHohadDNU1Oof4g2cr/7yz0
c5iv6ciPiwNoQmt1EICX2lodsFC8W8uzL4Q1thCj+FOpMA8aMkUEOlkodA72gqx9
7rdvbR4X+hSrtUQyfDmmtGQ/eU4i7+16WJ/u6ZklE99ybfvRshv449ggSNEkVYpD
ixJKKmNFiNa6kqKpwuEv7EB5ZdEib5Fw7qex1XZI/v/gNJTMstfMSuR9Pyrt/7yR
3+Vt2qBWEHzgNUVSW2nKUHva3GgYWSiSbzlFb+efTHLSlmuzrvV2/a9WYesBTNcd
wW1NXau23IS1qv+NPrKO/hp0LWeElcwdwo0eJGAg/fMeFjfi7lHGiQjMgS8pTnAK
IgLIbtM//lxNiCVyeHaE9RAcUbsQQDgzDUsdDXvlrdN/ozI5Ldd8MEv3jOFlb2/N
TN8gV8IW7sCwRnOv/EZk1Oz7E+PskxNtCgkx7hXBcaYAe8Mv8iuvIpRZ84WaIc8X
wzf0AAOvfNscR3u3/d9q5UsFsXbaLjK07A+78uCiwAvxcXKpuivYIgaSaO1EidnZ
U8G91Xus2wR3sqYE2MqVP9yUXlss88uYpwGF0NtJnBh/RtDNflntUuw/BmDfDDri
RM+1agxyZFqtJ75Gxg+40WPGUwOwzSt2jFuvAl//1QPg46oHhjmaAa3XL4/ZAGqs
C7bTWPC+r1/XXBUfi+RMsgPlGcNZcjCpMSNuwHFEjCxogIoLPRChC5xXkLkzsXHA
isAf4s9H5juJsGEEwN91aFeLlNCxqgn9wl2KoLqpmR2i3neU68YOb6nUl1fEakkj
tjye9KAe4Uzo+pSXGnmV1Pb5jSUBgLxIYjUktLdz8Hh11Vm8DNkpAMdnULOYze1x
Ba+r8a9BcB1+Sk9Vwl3Bn9DXrGxrLGkkRJlnJ0x3giCxwIj2EppebEuUYAfQfwkP
13cm+ebvh6EAtfV2K7N0s6Jd6V7EpIlIR3EaDT5ylDzUMwEMSENjWAIJNo12AuIu
HcZSHkPmVR2n0vSzp3ohP5RF90pWbBr6J7rRKIpY9JrRxNnJNcSIOXmomMvmB6RQ
GOaR1k+L4IUPh6oBzqOzzidjtIbix9d5qaObE1JMOBMfyTFM8Cj/6ecSum0SUFrD
6hZAOFmC4L6vDCNZgRYrfuuob6vgosnRwxKsLouqxQQ8hvSkBeq0JdQ7peQeDst/
lnYErwhyOy5E82v9FBKlOXiLqP29RaunsU6Pb8xisQI4Rfk/LbIIjXuOCJ0et/f7
uuLtbBRj1SyDgAiWYAOLWybfoY16fj0Obw3qWNKSDiQ7dYkts2b9JuIK3+sp5koG
hYF8A8HsCIxAqdmvJziD3e0eK2WW8IZPcTUqP7aTvf23vVzEkj0WzPFA9GFJt/Au
EkRDWSo14xEnxYGWoQnjWIwFjCTXD8QZk+5VrXxH62RJOfaADmpJUlS+7fWcEmsO
PNvH9JgUsOem9+6g0aKbcJVsLYfMgjSAZNoGtEm1OW3PmhbGpxYscFNrTMIWNV98
hLnVNOidtmgAg3rDkzXEdM5c4onmtqwDpRyn9mkWcki0hKhLJqgKxq0uRhYr/tOH
/ABBL/lo5GO0AvSN85csbZ6EDrwOhYcy5IftEyLEH6s12Y/OzZxkyaNJe4yG/bua
s/IJ8bAKYT+S/nxDFBkw3ILcUi9Ene7cb+50KhDE6IJ7715hfQYSQnt91PbkBXyi
QLY4bx/9A+PzNM6U5dEqDay2h2t1x/xuKbve23tlC3EdngVDY1Yi1pEzIfxtrO8L
OqkMEEH+UqXllM9HG4dDPW9yrUWxYTm0IXmM26jB0Vku5L6DcLlzKx3aaft3oj74
dH+Lbjv5NvD+9Kb9PAlIdfd1aXbhMqcZpEOAayyl7SEXEw3wkUQuNB7BbThWsk1F
Q0d3zayTPJ82jHuWoiTfdKMB07JUORW4PgtG27pdYXL7Q2ZN5IyzL8ICOQ8gKQuJ
nRfTfA6/pdOxBrnwVNL+E9mdMoFfO8WwZaalYBRmlMkccvoA7Y0kU+msRW57pRfw
6phdFK8FeCCUICE3zHUbpRnjTxBnJJG5LVqeSSfB5uVltTvNJREeOVEfw88E8XNZ
4hfHIZDPhFfkq64MRPRYrRvNnS5g3HRRa5ZxnmTH4SjT0UeMGDXmBh1VhukKAW6g
1FZIpqoW3unvP/8cKSO9+UgvxW6SyCSNdISsUK2icHlJu589gW8lTolZ+3NmfvCr
QS0Y/hlp1Vprenfmqc1CFABJDL0zcWfUm76CiMRLCdx8MqgS7HKkUK4lQQOlhhPX
rFN0YoHeirWmmV3EX2q7qhouSkPdfFFlRkcV9wUUPyhbnvjJ9r5cFi8fyvLBoQQ2
ZQQZnFSexhjqOcyNuewCam703LhzKcCIyQdlbx0n8+xa8E5Lvd48vjvnA2m9E8Go
fCGLXhpE11GWIl1K6xLD68gVCp2OSwCLSIFioSkQEBtTUmi2Bcg9ml+2ahsaBCxw
2k8ldxQ2nUpR3FaTIhLgebullps7T+9feRcNRqfpEkcNwvTqKpJhKJszr1Wo7XFx
IPWi/aDmReyxZ/wJ95BsJE5z9NG3iIzJYoQ5zak37jJxbxsn79OvoTI/cuEVW3hO
/z4oDUgJ7Rti19472CpfrQQDItwBboUUNHz9FbXIEF4rEQdJwTkBgJ9RgUE2v4mL
fa3403Niv3u6q7buYy8Z6ROoIPN5KPcKvPK8OqgR4j3WPJna44RwU38P4Gya+VGb
cDDLZsqAM/0iCMNClzIZsEmBrcD4rnXiHgO8jv1pcBtdDoR3GC8EA/JBNsOo82cz
o/v3n2t1UoFLVvXz29mMpc1aRBq7oVX5CzwKF9Cc2Q3WKLRuE1bglfTPBYbGB4ya
XNWsuXDvXul7yYWsMcLFCfwq/Ktzi71dJ4ZDir/0/lZZA+OUjXuZir/z8Pmu/1/o
vdWd2yWiXJsNFd28GUj73J02kAAbo0byK7zFJ8wGrcHJgkqeTYNNQmKbnjQDy+mZ
SNen70TidxUM+vXYfMYzWmf0xw3q/m1FmvxVJXftHApe9i6QcRssFA9zaB5AlzwI
lt3ftQ1409sxo+uU6gReWUFzzxrqOu919NaIlAmlE+sS9dqMWtLvVW+DsMnd6iL/
kXAI8SCMxpbaqLm475kUy/u/IPAzNTjsiZhnPxuAgEGhblnaKoyJpTGDKL+ejNXs
57aV0i3uSzXESr+/MIbX1rUbftQKvGS90dvxQCm8HxsI0M1N7uB4Ybn85pgvLgux
Q1cWh8IBPnlwBpAPnx1XEuYFoqtPgrFyWalaS/cIpaNyFSJB50hwv23gIUXP1bHF
QGzACiPojWdKIIyJyZAciCydAXY78HtDwaPAezHfMeoWKveDuNtS3alxxXi3ErUT
FKDCtDJShYmBU6C3hIqfkNlhkm7yyVxdSvlLO+b6s7w0Jl7yFcVguTujWk4mv7Gb
eMYz/raoNBFG9jJ1X123bVMTQol8VXOcUaeKrVVyyF8ALfsq7EzEgFwxXcv9PnMG
sk8xAQ7vpHu55y1T6+1O9acNBkbOf4joce0U3svBgHQmO9Xp4/xMPH6dIb7tElgG
Gx6dbkdjjF27yC6dkBRhDeKOaZhZWs1sEp56Iq8Xrw5j74yMRYGpTa+UJF8Jh6x1
9es4JquLYMGpn7i0hOF60YEFJYBx7xPvl1SiDmBJYrJlTr+qxm/SowQYABPFyeHE
+AFoi87H2D09HqLO+tyB9GvCn7I1DgmX4dFt0DMPiPrlyvHYgJWrf25Lr8WCZKNY
zUoTvDNY7x/YYO+sRRiLln8t6UaEMoGWqu+FVe77Md1yh6bKXP8/kQcg/3N44T6C
nBqunK012CXv6h2+At6Gz7l8Yl+Gf0PosombDoafUgrgzjNq+reNhj3fmC4D0ffW
Er+qYSq9BANUCL1I2rdHZk4cj+7ATkkq76GXYh9jlCJIXjtdWPn8gAEKJQlYoDBI
bsny6CYKcYrVYvHqtYnHJQtDIOjJkQM96ONXkyUDmJkFqaZUS5wSaOUyAzqhlZMV
Qx/WFhlHBsFyMZ+5Im2P+ozWys+waOsxP1/lnqs0ZCnCY9dczl6WIChmUnjTGKB2
O8pt4QywVC1UCB02mBegV1ndE0bMXoUS7VyXjgRBbHiGuYDuv+5T+OcjEAlmCCSC
emKYJzcdZnXy5nnInvHFVW87SbXIqqIUddTPpFc1t7m4YUWiOtpdi1hynD0q6Xyz
t5nv302N6Xl1BhRLvSncvNezmJheLgdUU2uBdipdXQJgLhiPcKJXifwLT5aCQQ9y
lCpKXi1SZQCWRURfqij6JhTWU738L+98vD0p3YcB/hAumM7hudNr5yNI8UBg/OBe
mqk/GwTid+PlaBA8MfmEpehnLYiPhMYR/vecz/2TZ7UYIDjtOvybaDnM+O4S7M0B
KyTjTBBLvu3SA7yWhaSGIXCgwycjD802cjIEjMX/bHxmDCqvuYs24PuZ7TRfZVYA
pUQJ5qeGzBPYT2tTtrqIBdaJlq7fP12hcCOnQBwMAceRUfZ3uq5IwcDEz8KLTUJh
snoz7akNsmwEDUvyx5roOqaLOcI20UcGeDtJ7b8fPHJME8ojD90TYSxGNzhUZxZI
k4AAdoKzp2oRsDyDofQPAahfsbB+sFmjqUcK6onZpX8op6f1Z3qVLY0AzSfTaSWb
AKbaZS89FEUMtqhuc/xt+bWCxg1jqQngN8q5sESJytcdwu6JCNkC0UyhGZDfy5J9
XxGpWXvnrw1vDoC6s5zeNHUfPV3ka/tlvxXmg2pxyjnPvaLZ+KP+a7EVJ5romi0I
j581xGguxvqu0//tRZIeEk4xn2QhLYcdcWMk6mmjn+nEKoJsrGKpDf1RDGas+2Z4
2gSB8kTrztbeyVtpHob1nzemjoeJ6zDY+iv8SyqmkbcbAtv58VRuSNlqGSti1Dm1
wMlV5WTBhyvafK+S5qdPSSBpaaGCJmt9pBg+0S6h9+mTMJ2Ff29p9FiVwc27Tkv8
pK8qNH6gDdJdmEgb3UhPpO12rqtYQSXUAWgkLda2TS94aiz4T1B/L4/I9riphLGB
gbqrxwuKNHfGaKG+ScS4hphTqkdSlRSMcwhUYyeuRr5UPlKjAK4qnrq5tqCRLjPO
8TlXsrrGbmeIIkVieayF7+wwEiVchPn9dKZDgOd2LuwpMrJpHdMOt3dyRpZR6bqp
Xq+yqhWxEqnwwr7PyNBA9eKw1nz6Bq1/AhhMkOH8Q15PYRcUryNASw6YOmAK8g6L
BQDlRGbbF9j0YHOV974bKCLba18SrhRenwGt0jDHsdSl5G00d1u7QfI8s2eu53D5
aQHQdEuO4J2IBVihmZ0X5t9RGbvEhIGrLt/SLIJ2NWWwqQVngAysA8Z7jfRp3V6N
MeXUQJXiN4egWotGDVSmXLE/E+/wDF8p9QfvT4FK+k5tqBHs/u9T8YPb6zgOtcpQ
ZfjkouRy4rzQRO7lyUncRB5YgK/oH13l9aGZ0QEbApK0czK9kdk+3WUju1RlKRFl
ryI8V1C01jMcMMDZxrgrodb6A3HEFzb/psMos/YKSiDWTEIxeWD3A0LUq4z0xcfx
+vjJuxvVPUeIgpsa11yPwKNx9MZ14RtX9k27Xszq32poye9PhmQJNiGJLvU6006P
S9WrSPs9WMtkcLGqDKkY22N1nJIInu8fZstiMvypkWjgHOgUt3BVlq1jFK5MsngO
Acj+qn96NQNPzfRd/haIArIZFvTZjACnBh6ccLtszueyqhYvgv/V/51ISlvnNqgM
l4Xt8px87ZHuPPLfUbueOte4MwnDliZh5zBU0Uxoy/CH+3QtvEL5Zu6dg3uGvfQ1
rllVt4o+3W2XLj6pP++fWemmthUlSoyOGiOah6z3f+imQzvaEc7t+O6DOdd9GQNk
GbPacu4bj84YD0CtsoIBtLrT3JKSkTjEzU7wpT3CSVxmxwnB4xXNurZo4EwdMUm3
OPHThhJY60kI/C5VRTMNwl2F4U86O6q4/F/UrEARcEgIru5l8cY0gw5H1qQ8aoEP
WHb1DHi7vP/wtcpD0cpKlcN9K+SJYvIUL6L48/hoG4Ue85buEkj+xUjXmVp5hNV/
TuyGMSZklSaHZ5U7HUimXbP3AkZ6DHEWbQIaIsLTDjfKm1M5g3sX1z5bDAqhdFQ0
S9u0DSekx+yzY3ipFNwzQS9G8aOId/adlGQ5TRme0/iHZmH9zLedmEsCMXBm5l8C
bZ/1tkuyOkRLq0s56MPB3BTOSGB/xfwugtSdaHpXtWfgMawFN5rqO0WdvcwWTmPb
nfc/lSHviAsT9mezZ3xWlP0qI4uGxgAnUE9lPzzdOfI/XxraeSeQclyeQ/5jUap7
CicMTQkZld1vNuhnWXFR05YJYmGu5WmG3+T6gRTU7ockBe03Q24Kzo+9FVas1UGU
Ygmd4S3rnaIwBcmVQ07FzHWW5JHeuRKZo8RaN6Bnf5ULG2bUEZbTTpsuG7LPHPxf
+ltFBO9xT4XcWg+n6sDvEeiJeRWuI3umkno8EJZOhP3aqAFBzz1rTPKD+LM6wG5A
6deEEdGe+qwM0cF4L919PAqTCDbbRnFFaLNQSaclvMHGPne3SD6irphW2lBlAyJc
pz5V/pVpS7Y4YxKabbE0dzqffcYrVV+VGbjCQiqtqEmiScUWv+4WWOE4Hof26Czn
/n+CA2cX16kxJsBgvUIOD7jwj4zLxMTwImzZuBYtCgdSAowQ3zW1AeUiCV9ONZc4
f/LCRvZpjplZlBf8MeriHjHZEU8vWFg7lDYGbmpntSUFmaaXFvrtuQc3jvezgVzF
2bwG+WlOJWSgM+NmfAdZJUhR10pF23j+wtf8JVCYdG8FzlZktDdCJGEZamjBQ3oJ
FCHQIr9vGeM00IX0DplVQjZLDUr9Nu+9Gig0AfC1SQb8LzPhXuwKfChGLDfKv34d
VToeMjkx6a0v5D9T0KSQa38nt/2mfxlu4wjrztKysnNFmyED9ApLL6/6nxcF/CZ7
6c4ooydiurVNsG1NbZ7OfLSVrWFr/wwwOiRik40fDdFEy/9242VD4j9mu1/3W2mz
22516ZqKfCi3FTBgFPuGeYbDOs20J5tMeFN+JM6T5Ar4i788Rp1LfD35mjZL+eVP
JuM38F8sa9pTWnEc6dyOCLjmHqTONYMKdeT5B74U5j17DfzCZ39ZOIX4KX8oqBaX
IkvRnXaa3zL+4/hykYk4eNOWq4IGm06kcaWImWTecOiP24UFrTXz7VnbyNMzsXJc
oTXCo+TO3cKc7RwuYzzmQ3HYv+xCQelwRE7OLXM2Yu4lY0JPVn9kZvC4wmtyQl37
ncRYWnc0yfZECpyGW0QwVSisvVZboQdrvvZDapIhW30b9b5tTqzD/JDpWS0j4bPx
uKEQrEc8gZUMmtcwWrbAE2449r4ts0NCTf1HdfZdq9ThF983eUDggaHoEiEDaiB4
+KC4edf9qebkUdQ3jrMMNq9OOJODAs/tnKfPhA6kZXluSU+N4Rs/34CxWwKqNgUb
CJYecr/KYHk9ND52ylSiixSKvJdbuxaHuTUAKEbh4wa08Efzm9q9duFhYoyaCDKR
f9KPBImXNjZy5qTW3FqNmjSTonIV7ZzLhkuCijRhCX50YXBjA5GWXHI1pM/AZR66
YuvjERHn/sOJ4yVfq9IlWNIY5y9yo8WUSzh2C+/7d7aPVoa1jdjCPKlSHQHMzVJc
+Ar55VaMet66jgwuW310ABKLpmbW8lMf42DjFeJfpfcUv40bV0vCMVp/4LHaq4FA
H7GrgphMVgdI6KTLFHjZoU/EoZVkoxdqBj0iURaSfm9mf0aHAhLfoGc/Zmtd/A6o
+DMaCJlL6dH84bmE4w0g2a+wIlembV8Fa2efyx4cBxM7MWS3pa2Nt6QOj+cbPUVG
mXL0OqyejTZfkN/VT5jZJEimBoBNrsK/Sx19SwreFWY9yjkIKqLn/W4+EDMmwS54
9zd1P1KXbHfb+ItvoQg3ijcRr6r0xOZ7BikhUGFTrMWfoW3bli7jYQ1T/oa5rg+w
dXnFYkCCmTH7y/e+WAXNVprvt9J1brZqIskPducQaComOFEAJOwRVHXLQ+4iKyXR
aXlbNPR1nL+j8k7HSL1JtmCIGkwyAvzD+EB4NW7Iad5PLlPery7pL4KbkZ8R1oa+
iwXlmP2cBPPbe5RFvznjDyfotkDywSWsmwwOssgSxRrC1Gk3N67MAYDTYX7b5x9f
QZUXt4ZGSiJRjv6bMCk6PKaNqPLi2zR/34yx1I8vtHMWXwW2UWSSjBXVQRMpcNtD
2cMnxDbCYfAv0q/H6dCrc/iyPlpvDsYprnsx6lgG8qseMH/E6ZcaP9Lu3m5c9Ot2
T3hELthYKoL6P6oHTaPLGsNAUPGAes68Z878NyQZGx9Ui72ll7CX+AlptJvwBTVH
qYGAt2b80ZDTkBC47I7ixz9pfXYiJfaJS/sGlrXcBuO9OxYGIbTiulgHnll0BLA1
KbvU+m91jIaOM5C+yhpqlPHGDAT2jvZbsIEAdSTxVJ/RPpBySNXA5h5HhViikzMd
eSYW3+evGgVVhyg9mi2KcNeQweYybeqmoPP9BrZ9nEcEiMfrfNQa6tVgFpDsrf+V
Idna4nhFno7NxOgUejg0mxJdq0sJWsGOn7aRGisdV2MhDT6sNiLctJuJRl6yNlaQ
y2uaTIy62I7XvVmdYInsain8HIya8nlHy5aUVv8ffvFIztq9QZwGfR2X7nOlsl+s
Zc4xMO4t9obSs3ftH+IRsNyr0juVqlVaNRU3AeRrrQjtLHWEOQa7W+Bbe2xbnOxN
H9p3Jzj3wGucCyZIUZliMmA08whailOiS4wEXjY5AeGeOC8d07auKwfQBqMLFcz4
PuqODoThhDkZ6kvkhmjToEqLDO3CC5DPYX6RqQRoC3jsHGyvlSdiPkmZHMT6P5ur
kY0K4+QzvEumoqTiwik8xcxRUeiGf0k2AklAG9Oqhii/GRrhs/s10Z0jhJPKp4TA
lcokN7guTaNAhDA8s8l4hlg26B9wwWhjElaXsGOSrSewoMTPDccZ9F9/XrtJBI7q
NREa/Em66Sg6Aasni5U3J+w2fykjwCHm9GLWwImc8D6U0mYn+NgUZAUblfiHcf2E
u+3VM/HD+ISoTruMW2mrtnHZdbyXXkdVN5s8LyPGHmMtUrHY+hS02E2qdCM9oSkS
hOU5Coxe3vUiggj8INxMCAK1a1kcpmhcYOUMpTe5mhEHPzFToACkYhOy8PXDx0iS
HvujZqmkHxG3PyMAzG+HhXNk7+T18CqQFUGmrjqluKd9CXVo4OUIMQdJRthcpKE0
vfYUgis4c0CiJIkRjXf8t6x2etGSUVn7+cXrZ4qSggCNppjcXDWFFFo88t8WOhL9
R1SVFXk4KSZHJXCY5OlHdYPcuGon+809hm/7mAT38shYKajHVBDwD5YYxWA/EiIN
9svxcpvC7EOjy5Ix9lqqNiQkkeei7qZ3wIBnDnmTUw/3nNOCiL3qDyy1CkvE+NrA
2Mzs7WO7bpYuv7wruWK7CSJ4PHtXSNoJgz8LSgnEDsgf0GvwG/cLUrtb7D4CPJtT
WlVUx7Jg4OeVzomKNVz/Ept5xZAL7N38pe+3TwXqzzuF+c+Gb0hMO5Z7q/6uLqyU
+6xO5oWOAbVKkazcE6G8dUKYxGOrmWP1CSG60XaJ1rH8Hbal1wtFAE/pCPHweRoP
DmUxoXwZh3EDWp3UeD4zXjwpOFRH47ScL8KRLbpROj01utZZr8DFHn7a9VO/T1jZ
MMiHL+eZ5ohisIKgKmwvpvp0TwhDLWeJq/yUWlVSou4ErDfgRHSKDKO5ISmyL83B
NskfJcqXkwN7MNdc+Ez0P51EPG0CC3nDyVlIZO+4TaRM+VoPn+dznfJq8NKlOMsj
p5aUEjL0UgCSTbWHbisOHxXiDSjOvea5qRdv4T4Hg9wJscqrWWuGVxXb5rUbJiKM
p5gwLXJ2f5dipjOvHYsuLbjvYyGCMkRgeF0okxx9b5eDk4gxIIKYc0KHnn5bW8pW
YTujXdnGn5AiE8SKHk6l7hr1uaqAP8DiSxRP4C7nj4x2P4Ymhu8n10knR706d+6+
BlV0YssjNpkKJ3GDpFuWQJ/WTmn+u3wxiqHOQmEZMzf0SKey8Pj96YNh+/A3bK5V
kmeSKnZ8RMIbnENM0zLlPKXdvsquvIyyknn+7wBbfGigVq7gX+U8A2Bl+3y2oAI+
ddWDPU/sAqmzhOHK/1cbk5tmuF+gyMVtHCMLw2EzSuhB0uDSXXG0Gs31+VQgysup
o8ZWG/q4YDwfUJR5ZJaNC30K9YYRa6kYcJJoIXz7JGpDvqcXTQlp0GfP5++VRYh2
LopJgn0GFVuDNbVf0eIYwEAKrAe7LmHWPst3lIIn+R3X9xmRGWGD71VKgrD3EnxQ
48aEbjx4G2ANVk4c2wWhCvjNyiBMbHQuNTcDld71krlE8JahUJF8VGn8EF7t+yq9
VWdHvUmo6T1OoTrtNuywBa989wXHLMhOfimYpejgtvXqWBoQ7dDRoQvSdMOEVWbL
a7aNzntKWaEzihRorAPiCoAY7f8qx7JRJ2ReFFUVP8h/VSZcdDTjwBk5XXnsN0tN
TXwm8JeJf1JexB67uneFqGmhH+4dGHX05h7sCYTGty4PEZZZ6arEOlH3isWUMekY
+iHejBNHxhlcf48N9SkeC+NklEB8MMs5CvNU65m4rZjMqY5QOYBIyH9ao2nLakJk
MRL++0CREli/h6Nm0D3iJqnh2CUfUL3Y25PfItxQb0vRAvTEdvRPpDqd4RQnVqtg
oNiO21VGTvVEOAT4BcM1JWE749oCMB497mK1F8MsO0/FjKe1FZ4rJfYhpmqboNB4
6b5iMIeLWJZTaa/Ns0zvXkGTkvdgRKpjubdBvifCzTCZTe+3KpaBpmb+fumx3Hqn
whq3oylfeajbkS3L+bdgFSZ8pGvQxACsmQ6JH7OUT1df8DUTya9LANpyDAl/QRJ6
gYSI2oXF9MvVX5PmkBXyzcelQ9nBX5RLcKeP2DzrQKeTjvh7t2XsHNoDDCYnqs7o
JU16dpUeZHSq+85C8l47xVJgOZKxPUF/WF790zBuDbhjRokEoExk3b1+gS7gICPG
Y573idHNlIecWp1wviRgbspxzGPD5d+/gN1dILOzBy1/+lqugcOaUbBZzCtfMRKj
uZvCNvwkvN5lMG0Lxz6s5z4FG3wl22qEfwuYq534EFDmF+hD6PxEqlZIDOIitLfR
rX4sKtnxPmgOsAMObqG1r+0BcGJV/PrYTiO3SX4PhU1dKUqMLU7T8kKqIMYw//MS
cS5yp8EZdF+pt6KGeznE76L1ecZlh8o3a13xeD4BDM7T7rR5GNPYIluBhioHjzVV
tacdQJ8BlUqFhdlqq70QHDJLW8kkIZgjf8yc0DxaXadJBUzYyELAZFh2ZX+qqdym
kUbo0BS15e3SquVapVqFDjESQUjzAhbldg9ntcXTOyv0h+bASM/DSRzTAwFEn/vr
ZjX9chIkLA6n/mzs7tYb5CPEbtdVoY0AJ++FGMeULfBY2BOH4hx/D7VeaZtJcW23
uHHFc46WO8EcFmBHEy2hRXqDlS238BSvs0tyriIxGoF61MpC5jognHC2NBjc5wa0
7e77gmYWWPQq+ZtDvs5EnsKRq5FOkzHaT0FyQXn0t59TKjslYNIEuKITDyiha3qO
o3zZyuV/slSxH/UGwPj4LeSGCvBDfJHYwYyMebhNqTkQfMZwNgZJYZIEInh8dQnO
PDkIFQtfVqXNjWZLKtyY/JvIBe2RNw2DN578oCXUJIxA/Hdi+OaiOIftuggMYBsZ
OOKyXrrZPq7NJhwXwVuaUtBKVWDaIbZYucWCxG4V6t6cdHURhWgNpDUCU0Q1Rcby
9WaTbEdtLyaYaQE63F7t+bLOn+5hKotZGNzVvcr1opEsFVe26oG0o4bJPQCrQjGB
V7ABZhi2HMoi32E7sfyIWOOwEyG/Qm0A6gYK0K9igc0mGg1Y/zhZztFc1f5i3M8B
1kxk9t5a1FJIPtr6KeMW1AtXsPyGScUfO1kqa58qXGfss9rOfSfa54r0M7YB+u6+
QZBYKyFC5zkauWi5bYhdnBRPTAPyPs6oCapNjOlumxQjElId8aM7J6nntq4sLoxW
cAyo0YFWBwY9DcH8/cAX5wlozYAspTzWO2hsQFNmRvHiK9sQChRXBHpxPuU+1k0X
EluMLoyBtjQqlYTs/iqxC/Miy5w7eBMOlodmbxDMEsSyrLlGuCAABt+CcDBE7w1z
LKZzAZK0iJf60YCPKDGWvK3nBNZbT52PaCrhea1o7m/TMYiE1Ip0j9kI+jUSG5Uw
10mhNQE29m7I2D6hiDH920djmme7vRKc6oidUi+LyVgfmnyOmfcqIaTw8pixyEf6
eP0x/FiAlcrF/gpWjNpL4mKwk2bbWRCp9//vOZL4OhxC3vh+o2oNyyhlsVvgBFQm
M3DmjY7TbLl9qEG+3Kq5j5EqE0StiV9pIlKTSbG7PbGcFAKXI47IXJ814vMabSfj
nv/hwn6rRHAetkXSB05pe+oMMUM+yX1teXkhqz4E3y9Bf7HNSTFzYCTmA1k5Kuo9
qO9Zby73Vc06N5OVyg3fjdEUMytFINTLASpCL9f8eCcB7qO2xy8lSyKCVA99HQTh
M4MI6HHrGsyvPWqyfL01HitIT4dNiCg+d6+IrYjEoT8EVLCpZZCdZGSoZTSx50dJ
x0D30gFejJMcqPrvpVvhvOvbeRumqqLPgjYQIV1bIF1IqFzAvMCIvvNu3xo0EZJm
inHzB7CtmUTmGfDPkQGxcpuI9k7IAEMPG/cLUTYkM/ZzjyflMU1Va9zN7il16uxK
BLxg0+DlitHisrOvoRcTE5+7pE1UeVAsrIhj8KIFmIzC4otPoGyL/hw20zK6AJ4o
D3tOaDLaFFtxYNzrTCmyBUDEbQgRPkkmwV7C9oh98MXLAxef2wy+l2E6X4Vpeq0S
l52cvGdqxDs81Dn/oEt+DIXzIoX/Cs4v8ByDmVCGajp3NtTBaAs2BO5nbFQQxljB
svMuO0hdoLoG13IfktRarBNQGjzQ3p6aHZPdtxgwMoQW2+7VpxX+uuejo/p2aRWX
FJbNoQPAxLYo+B2H69jA0XGQOUHtvCkC6l5TN3EMB9AyXx1HQtHASV4by1wfiaED
0/CQUppRPDsqCfHEIT7eTib/9GK4+PDeXlBG8Tw4i++IxAGaocrRo9lWi9WYT0A6
HqAScoj6YtFuyarYDSXljWmD3Uawh0u7geZY4OoX6zMigY9ZQlTb2KVPDc5xlUxm
KyrJ0LSbWr4hvlcVV46uffqj943Lwr+oLe8vTVYjKgWk4VEu1yqEkO+rGPhbQ7C9
JEqmHpsBraF3wu55pLhOzPMPMMe5pLsVPxZZhqekylBrwzsWitfpt5Gbnx8GELtV
HM9XXzesFp69Zpc2wiFmIP+N+JWxlN/FU8QWUptLeSBHDf177uxvb+uLubXaehO2
9yJzqmTTKtsrCsCExechMo4AatwAGBvfTDieApr7R6aJRZbSaPhxyvl2puyOa2a6
lwmAEriOJXZA2+m4jZd8U7Oam+G/DwcMxrRttZ0t+ARCn/cMqSEPcaKk5Y6BB+f2
gqgDFMTGhF13wGDHEYYGd6sIvrSQIkjJIMW4CAHzAumM6AXXpYqcOG60/+y1niem
fRDawv8wUDjls5iAWTG6qijVXOQsAGa9SCGwKu3LYvNtrvhr+gbZf0tYijd4Zr/6
dYXRLfZFmeO63I6CvTBTB1HBvR402RsZG5yp6OdIU2kt38Bev8OSh2LTNnPMHRAN
UgrxEZcZOPJjUuRQBDJ/7lmv2JbKsUEJ4os8nf3lsrEIxvfLTW2jYVrmxWp3SYm7
8y5brqceVg0MkIW5bkMZTwGtPcvalkb5GJBt3w2Fc0iYbuja1sq060W+uHdgiD4F
YdeBwZ7FKYpedwz25TfsJH5GF/6uwcuFvIj45exH7vVRLmFBw6TVxQgVsBG00QG7
Fmv/7GEzylmq2E6OHK1pX8chQuAi0dd6yuMbnd3M3xqQHY8qnPk/L5t0D1k1aP6H
AZ7CNMf2Ds2KlzOM7sTztDsyxkHVzS1BJeTGycWtlUjQJv3dJzuFbVvMs1Tcvp2c
GOUsJWCTShZLbQEquvvEX5LtszO8TPu0TNM9rmLsA/HVAQFjYK/ZXutT+u2I7kXV
KA+m0sS5sW8y6HsfeSrAyKNHTs3vemHku8OG1+PddYISnEKLDqduSZ43kykFXFvq
C5c59T3mdXXPwABY2YH5fjqMmoaJPYZunog+DJDgcnLkuQuYP5IdAod16V5jpwVR
p4I5PPWe2oWAnCB0DY1OEvkKdMbVftmUfNk9OFMLI5j03CuauYPAb3ugdhO/r+sf
mf6R8zVfgKBXqeTCaqal3j0GML3herhh/ITy9N5kyBJuCE6hKWDJU+9zUzXMYjLc
LYtEQmIjfBjN7k8Je63pezCK+x2nFO/BSJoMOa8xP8eKXiFN0D8Vi7ng7nsYYhWS
HTh1Dn662d3EWWCPWqMm0+n+sSXQMA11w5eEwTcCkzEE4/m7Eoxq+XIlHm18C0zw
GV9+ylIAWUI9aAMR47l/RG4nqFKRlcuFGlX2Ny0FgsDcR4vbCqUgEWkmxior0KYR
OWJO8pqeaSA27QPaS1cVN5LaYOVCRzibBxvW1mNj8ezYehZi39+BTTtir3dABLv8
1tcUFT0eZg6B3H3Rq1ygzAoszW6D0aIEuk5tT0fsKb00NtdM2xe07SPH+3s6OCg3
iP/1UujBJlLDLo1zDgYZPBdsbDieVcw/X1J7Ra75d+AvPKHa4aynY/ujdxcL3gOP
eBMPBEONTPJSiJzG018e8O23n8sRekcDS8729uhxwV7RgcaeoFl6mOxLIfAV0n7F
VHn7KFstTUD6XCbvqzg45SuPkruvmAk1Lz46FYy7LSRra7BBDRXgUaPMpUGJVxeW
p6nXM7CBzZcrIn+PCMY9uabXbF1XkctfxHH86zi/gG17j8ZOsqxIFxA2MymMt4r7
wklKBHRC/n/T2IlgWHyDZMhvgWu/zB6KjsnbKUdDWXjTV86ESDtcJOhUgtV7i++m
gJY9cpE/QrbAormNShFQq/tZAGiFJDFb1gA+LfJzh/kOlYTuebRkzOrG6Z+uRZ3p
l5YRF2ZaHWoEOtro9ojvu9Wmcge3Hvk2niU7pqye7nfvLSrHqL6CCFgOofs6wZe9
rEEomhR7LuVN2vKX4r008lVy75PBDzrlYX/tYynTaeLyS5H6Wxy4ZP1vPhS6quuo
26XoDikQeSpgcV22C7a+e12xWV0uG7ucXEofKVeijmlSnKAF0JF/FSEBMa2/l8Az
fNcCcibqQiBQZiDm0rpnIisRmPRBz8OEFBtqcyppfyfT9opUDnRnZzXlzrqYwyj8
ZSDC3DzKvvZbbHsyYUc1V/A2yfWxbCCc5OwLRgmPKPbf4gOCaaHwf+FlNyBzEas/
V9vpPF/b0F+uNGFr4zkOdZBqQfAyrdbSAcTkBvfLsP4mKU2qn82IN4TvTZXPkdgF
qMOIyzB9B4MSLS7gfkvhCgIcFdHU6pvUHq0rmstghI8EAbGbS5odJmQhUSW0u9TZ
6yDRxMqa/vKevGrpFmWJF6A2725oVFBjHs694c9St9+Hikvcf3CKJXFJeTOF+8uA
2zkbhU1p4TQJaHB5+PmASgKcfzUmvzl/c13auyzPp1ZpWlR3M2SeMA3yPDM1KOZ5
orWtZrqdIY+AJh+5xsup19bnIcsf9KgKQF6wRYd5e9NcVv7I6DvYPwQ07bLDjee4
z8P0eTA8xywQF8qihrnERLZhPWAiIwAyQCoe5uxzhDugboyu2TaZMx2lhoKLGqme
c8Xkd0assKxgApFFziEpVubLVqh+iJrgKbKRDKrkNfvjdIXukyt0iggAV+7mgvQb
kgwBAPoi9RVkTu5uW+KpWB4HDhB7x7BRoDrspMf0GGEvsdSgAHcyBxDatTX//siI
9FTK9WsfglKAHV1noyviucO4Y/UlmgL4gcICy8FrzsmceIviU0j+aeOjgRcbb3Kj
JOpYO28obON5AfxDMcIwiRUwuPlfGYRsgEgXexSEBiXYW14nPNIGQGUveoxT1lfP
JmyWzvaiZLkSCjYHqHzAaI4SdBRXVASsRowhsCqmWnJFRGnOK6+CwgAlF3IibYdT
OWyRNVvCw87qOb9+t9wmNcM/KAwBaV8SQySLp1KwaGzzKe3ZRbWxSWCKqXEyw0hQ
Xssv6y+23yoTbz7kB9zluK6cl85/JXJZ0qw75MXk9/knvEZRy/qdqKO0iTy9yTqO
Wmqvf6WbP8eHiLtXaRb6T5kUAQ72Hi6oV5C73lT+ux8pnznZVAKSbScJiGe2xqwl
3oZU7+tSblLqGs2q1qUbgxhVSz9KpGtJWhqk50qtKojZMyhOhMb8JVy9TXye8myj
a7H7UQm2OsGUsgyJivY4SqHy67JjW4blaNkFR2MMtkfFZaXpe3nErdhhWz2ZyXO4
Oe2FcyAuv91avHHgDUZHg+SJLwg48nD4IHiRCnIgY30NYNij/xCjXr/d3fKFsbFg
2LBvoCEZHvwqrD8BggLd7hENviyEBdrTtW6NyAhRSg9o01VgR1YLjJWYvTda5GYJ
F2QM3wA2EImImIBT4LqGllQ786P+SyuE9lkgjBzDkuSyVjzEETTPWaRy+Cw50evj
9ya2GTOpD7aK92GYRiV38UmJ9ym2OChTCIoIiCTXHrBDx4Gn65IuSapF/a31SqSq
4H2/r246fT+gTAP74RwgS1NYk0+tnGN2pkFKl8//pY34wk5lwRHWGj846IjMiFJ5
v+3JYKpkM40zVfpk0KCdO7ryHHGa82Hlvfs9ansiqNT0Xl9odMeLiZfCFMUotbth
NA8KNcYEPebUZRpGAlWqx4PzyxNJ4L7T0Zf2Ff4OZrqtGgzFm9jGyIanFqV+5BKB
OFYHaHG8VykRsfnIe2envntVADal1EkDYr9ltr9sFfELqx+uF2Lju11EHyo9wiNa
Dppp085TXQHXdvsvOuswgrRa4F+DcKRULUuRGW+BCj8BjnXvC1wVbxSJkvh38TyO
daZSFEyDWuu9bjh4sSmzRxvKNL8j1FhbXg4oeYNcfcyx9AxHNt5JnCHkWqZUXJPL
39gKxf8BOFr8OSe6Nsli/HrBVyk/x02ldrUyd+FwA3Qn++Ily/pTN//HjuHnPItj
KDjVwRx7AFWiC4gtNn57iR5kWEPMAgeu/eEMUxaQkHz0q1vSKy68lx5qv0N8wpQA
j18mMeZux3GMIxVvXFuBkk77I0vItQtQHiZDJY0zaUMG1DNGm/OfsRMFOgAdLDPZ
7mDceJ6T1DlYKud5TPZlWpJdffKR1oH02YVR/z+tiTh4Cr7RriWcgL1yhxaxmDkh
DhI0zvSZLdqoKeSGAoitTKJ+MPZglbOM3AdHL3g2gl8nkh0Fjo0AMAITqIf7m/jP
qCQj4sH+p0ELhEfU0HFqdyg6sxRSjDVZ5ku3iU0FtMMVZyP0+BaRdacE8YK3BOGs
e/2gTDLJGcdG8bg3N2IoGjx0+HxfjjmxqqEIH1KdKHCjcVuMtVZ4MjY9mrdXvaHc
omqm+v/lYVPwFsbkivUwmWNcqb4wKEmzaQPrSeJ7pE597QkO4yeEvqxLCSDJUH6T
FNxQiGfxxSn8YHhAA+XuuhYBkbFV2PjYYRFm/Ie79C8TfmcAeADNKPKls2wIBmEJ
mLfTIqyAJ7gTMF/Bz58pEoC6Yv/GHwyLcW1QXXY+OP/gV7+oSjrtuPOzDnFe4iR9
yX9ODLwWcB1szE+ds9qaOqKBVP8j55JHD3Yk951tdWS2JcP+6Lai/uzIxuhyFxCj
KU39ZV6kwjQEgBrEVwCCkNZNCub3sEWHPkPqE2QEkaYeoQrftCLQXGnUnNmcFNmd
WXDn9F7kSGZi6UanAUI3taqsWk6PnHdjiasTLkxIw8/ZtO8jvypfaz4PyD5kgPBD
6ywEUiscXU80rJ75kiPWYZ7CXgk5Pq+gSNuG3WyL3SmHhsP3cn6KAUNmFsB2yQYQ
ZdHY1bdxTy+xaCxctXqIW+QigXOA6vC3so+AlIwZqaQI5VscLvHKNhJVbmirvKFN
OVT5ALdDQY02PKcPqzIcebOUNjvrjpcwWUFMBYAl7hWuVyprTfilOagdT+03nWpI
LyUHi82Ntgg8mv2zBZzaeuWBH+orizp/yGnZhLftVYjeTo5+RI+H4R2e8kgy2J9P
7+xDBUGHhdgxbHrEBYq7NV1WYhxuMnfN8x/rJsNuCcAKVjCEFRsordRxUAqZlpPE
ke+WTRttoFAsdmNlDP8UV7UCtEq4CJVh7oVGTTCxaCasr3I10NKUpbmh4jDTGd7I
WrfaKN/53O+7w5lNs1s+3Y4wc0x9lCDI1oHnjzfowszXKuVrhqLli6Aq1EdQz3bO
6uYCugM2/8f4spn2tzHn9i73xJM7FOA8yx1g0bPL8M+CllaEE52cKHcimJO6hq1g
ZmrVf/JkQ/U2tNeUx32EcrU8fJ9hB3VrCS/aHjqYJt5eAnS9f0OJ/r9iY33cZ4MP
6UCUy8TWcsl9Iw1LIhjsE5DvoWpWk6qx90tclaJZmLmBaVhkkMiwXh3HJ7Ie5gFN
pzjz6H2CYLqWltzf/dHpK8ZCkCHuyZNwvPZozAYzkUu0XO/lcbBawTA5e69/Mxvl
tLmBUeuOS34RSc9Wxt77eLBDTkNFDNduSwUecPK8aBzbPP2TYy5cRSTKIIGTnkxe
xrpYqiT6FpB2x3vXffxlmxegridSKlYOuDXKjPi6p6ZmsEGvEOkjQhs1HWjo92jG
GKKCD3trY6p+dgp9VU3xZuNUPBFhlfiddd/mVh/WtDYwvlb2PNjt7gU5AUUcOBGw
Li5dHeTWOhToRWMpoSDRCojmzd6xs00NfrX/TkdH8Uj5Ep+VII9Ii389DmvyjV8P
+R0VyXIBWzHJhjCEY/Ki+8Ot1nMnekESDCaMRkOgqJIS41qfUeMTE+jwClb6joTu
xcHz8ti6e6oCfQCcXCqsqeG1LZHdYZRviiVoCFaxqjmP7FDudaS3s2s6BsoaZOba
9UBuyfGznNREZfEyOJmplkgSKb3L/4WT22CzBkcqf+m/D8ti0bvcQ/TagBNvsuPw
3bn5uKWfh+Dnlizf/cuxwKtQZ6XBJ8QQqpxDucJ1s9H8ibddDlpS5rQAsElW0ihw
qrq9PZyeplx6siGCaQMwEcubB3zttWuZVQBxP6/LXWOD9SogTyFiEpYglCTuj+TV
a2zfVLWKwvx/uuxxypSuygmDBbB4c47mQ9YLjo+L0yyHQeYRNTqcCFgxtp7ptgeE
PRbXMGsTQn98frE2bY9LxJBQ5uweiHOwBdW7R79FqHSwLoNrggNTfBtacFZ8z3yq
lNeXE4vN2txoLPm9jO0qb/GlQXie4YTjViaGPcAxLjPRwYS59HZNaN1bBG8YNP/e
zJ8WOlVPMpd9Ysruso13HwG9JbSqwkKwIf3xsMthH177MDP4tgKU0w5SBrvkdOU8
c2ysiqRr/4ImuAXfhKpmMzVYUqmJgcvctiCx1Xbt2ZhGcmDcgUCQoqyBzm9K0LcK
CKXnG37Z9U+SrQ7Vh3xJAatzocClz9pRQ2BXwkegVzsrIdmA70pGtaRP88NMA0PO
QEkHpjROIJpna/g6YFTjkWthhrorSS7UShiO/qRKkcmjPAQkQvei7/SzM45WDbXq
QaygkeClgqnU5k7qrko28v4qcYQPRMTOBWZ0ZH9lFPV14/bhywTJTVNzb8YkLkFt
Qesd7dby+Kvh2VC1QbSTIUqkkz0a9qUENA+D/NqTzgYABmeBtcKaorMtsimNvwO8
kEDWStUxB4Hdlt+zbja7koprZOzH88bJG64uSY3D3u0kD+7k5SqB4nd5ED9wmwpH
q/4xj6Dd6y52cRS0XStBM4xlNDyjcQLRuoJs/OdRwMaN2ZcAX74WaTNHWTet/F7I
IDle9lOFf26H4LjxSkOS18mVaXHEO7k9uwY7z1thDYVKK/v4SWMPF2p8wHbbbukt
ziKIeci6rgMvaYZRR5XyFMUI35w6+kAD0lyT2NQjC3D32sN+Wqfk6hU1IyG9mDvu
MMe1DoPJaEY28H/14JiYp88FqitNkkfXXTb+fOey2N/lEIcELxEJJa+ydFn3fpHA
iPhNNGINJH5wpMVakRK8wtjvttDUSzk0nE1mMXJs4Xd4GxqpNSfY1X/MuarxgpGl
Nkp5oTFHAEZ9RnwWfem9Am15PY65+6GTkXUCUWRDs3ml7i9JLx6vodxZd32yHBnQ
C3ZFlZLOTolko0yrM5IVCCfItDT8LTw0hKD1hKzIV/f6qJyzQvI2vlce4E8xouGg
dCzLST9oLZrDY8GicAGGaWFPvtYdcH6Q9utlgz5pkynlaR8X0k3kdx4jzs/QqyfE
DtEjg07Ff/4VwmVfaZCgnsRSv/NRjsnYhFIsqwes348Rnym3fQzVXlWoPvS9Cw+j
IXXdZUuxZNR7D3BOZtZi33hajTTPcTd1cqmvPuRf6W0+wKrQvMnCmJNd1ogkZD37
EMogdld4ft/2rCs8dXDDW1f7ySLMo/7jMjHQdCZ4azMxVqG1UQN/x86Z3dxYMk0G
3HaYy6kOzZXfPKdBJo1LoL0K9NlJzAFwhgMxCCnxR/sFIOUt9oB04p9XYF9RkE8h
rr+lk+8MCk0SPp+6nRF8NQi5SU0h2Bhl1Q/I40HWC1Eeyal/kbawPuBM9kpjCYT/
JJSdurj8ZHC13HwCmHpYnP3NVq+YRT9PxpqHc8UMdL9kHzJLBinO0SS5X96IcKjD
bpfmB9uracn/1hVLfoC6Vm//j1juuFhVUuIJFu5w5olRsp/N8LBiKp9O3zoH5seP
0i6dz10s84tggpQ/hhGa2T8jwcmHf9AHIDNpSnFbfjkX49ivl/gJ/OuoZUUi8omw
JnvCnBuQx0uFQ8JWIYrVcXS5pfiMU2w/z3g9D2x+5bo9R25IEYjNONFLyR+QgZsY
VUFza8gg2enyjTg64+5YoPzR41UqacW12LkZxoo5ftvQUl/sCmEVsZg7oIKEWjIp
T3iPuLr4Sjf5UxBw3A+J6bmW5iSVq7den5yd/UdjsAjNeicWAQrJLQIDVNdr3zuP
iCpAjCOVI6O6wLKgXdwi6ewXKRZKYNMOviVyWrsd6hlNUrnRW16F1rlE3i6GxPRg
U04bFsV8tmfzhAti2HQQRdrH4EIE8+wpRxLMa1mpeGl8DJ64rXtDSSmMYvaQLNv9
XkbQu/oqQDbIxSN4EdaGPAbvPMpSaK2H7jk9UPjGuuqbGKSyhYpjj6v+x3xu/7i9
54wwv6+EijnQI3Gc5g899nCHwdwYGzcW46+20pgPPp5iogA2qPxBT9E3X/zZJtd0
Zz+PrXFiN6+493n5A818JT+VafHt0faOF89Q6XJ8cKPmEtkH0gron6CRPPv7LRhf
Y+LNQsRLW8D6UA5nbqAbi3ktLvui/R1GDo/XuMd0YnGfx78Tn6CYruDKlZN9+39H
Dudoiwn5daVy41qqISGRnPSbDeF39MsPYyXYgjxcfwfsbMxV0Bd/WUcTpq6U+7fg
E+PjHQxYux/5kMHavtuoLHTsFRL7zj0PxwjGd5/eYbjmJ+LIjRCYbos3Qvg2vBPZ
o3Vo6Dw8wiI0VeJBQNMWD+iTz55JyiE3idLTmMm2lYQlbo8niqXP4OM4+A1cJ+zr
3D8DD1b6yW0yeeq3MkakQ9O7+6Ryy4jPlCaKegdkX1yiyJwyGyA/FOyIxF/xojjs
NoukI1HK5jVKhjUhVKzM2lepXqKN37qy1S7sYoX3NwgShUq04IzkjwIXSHqrqiA6
4qyTpk7DmORzwZ1Uc0IB0NkvHvvy71nzGCIhbD6iC1xYMfLccAMCxDuTgaKy7hPK
YNhv2ikeWpYyPZwac8+n85IxRTbwPnc9QfV3kCno08dFOTgee+ci8e9TDHlQZus4
96sOGLMfSL3IzwHLOqvZ2hNY6yHKlBRUap15sdxRStXwzX3h+gRS4aRPwtWJDnNq
dDYVxQ6gB/HcyLPyu6MalA5Yscs3ut0uaDnBc45oaOz+StZEU/G/waMX/p3w3A2U
xIOZU7yytnpayRSLbWPYRRmGkZzCz7vfyRb7MHMm7X1d3ZkNf2f4tMRMONS9PTp8
bvN3EA1wB+i6vYYOKm0DmGpqFni+PdW+sF2DuahUAJEhW6DKA5lywRC8zJGtBZhv
KcXsx8ZEZqhlLPTypMVy956cGpcA0FzF7PxYemmBUqGAsoupkLqQS+hNFFe7Z9DY
l2meOfejX6ePr1Tx//c1EUkeXRPXnpC8QGdgV2DGn2RJ3HX+xt/mT4SbjkeGVbOR
JOzoCCHgadnr1VIAyqzqIzQbzgrddyWRja72BiteImdclY0GshETRxWKAjdkwZey
YhBEXJuR2YbujYG/rJOYbgdl/2cAuXy3omuRKqFlg8uMcn7fytl2R/g5v3gcefml
ZtGJGHZszMoeix8iohFq7+2XuvihHhNM0tYmX41saazK5kLLoq8TeixkLsfN+5s1
YzM9NLvkF2jF8wzY4C+B9q7pPHWXHhNTMUNfwNVruqAd7RcavXvvMtdz2fqjfpd+
ldfIfLX326JM8rJctIp3IN0XaOoLhmeDVXu9h9v+hf6CHIRgBD0QmAfZKqGUc8Pv
c0AUz35uwRIuEaeOjfrS8WuOoVSYn0kEJmSRO2TeciMCBnI/Ultbw5iQDFf/vvFk
qg9qp8smp8YEsf07ms5EUWSLWwk1FgOKjbp/8r4VWNLttqGLjcf3HLBfkY2GExna
8vYLv9LToNCa2tDU0wDX1aT1dud5ySGDuVUVCjrJFzMgoB4kG9bTVIT6oyn3lUEt
VcMjS7H8+2ACiQWF7+/aTuvs2i18+fZ/eZNkIKwfiticTQhxIyyzxC4a/8ujwc7B
4d9os9GwcgnQwPm7LZQIc/WTxetPxMerr8ngPI6aHRjzRJPbPE8Im10ztoIEc7UD
tIRffaIua82Hz+P5VRQKpCIO6ECihfID3qA/H1D7QCCAH2rlmdotIAJlF7sdtlDL
D0vQGmIpxJmjgXj4RaIZ/f4i+HFSU7fWmy9aGoYt/oHnemMjcAup04XImKkgS7wG
fivfYfq/ixgBNf7u8R4lq+cSFv5yC5mB3TS3HQr8/vYGITqmtW3tbAN/p36gwh8N
EcFgnIoD9fh61LtvsgUO3ks5ghXyE7l5VFrRwMZ6/utF/bUq5zr1wVtp3nb5bq10
Y7ohePTSMmH+WhbdBawxFEYCuZKLqtYiceSr31G2n9e8RR9EeNZ5feszQXrAVmV8
FWJxJ4EXXMht8XPfFeuGNP0EDS4y076FNZkOmlFLM1xuuq2MIC73Szpy4APLtyLI
vI0Zlb0QXjoJCKaIwIXQLkWSvvv4fvKt7Jip5U0yd+N2mci7MTcnGBFuE746Am0p
PNCnoq0jlc7J7mNb29T2+HxO4+l9apwrv/5Bl87NdNQQRjqcVVP7cZJJMwZ2L1T6
siHAxwZxAs/APA5xlQZMtE8AJ5ZMbkkTJCotSWPZ/Deu+O35dWMg9ZiEHWPx7sIC
wT0MnRW4NuAMyLdu7SDUng9qensn5f5xrcnqjXDOuz+JFW3z93m5lvkbX3EqxT+Q
IRnBEo91OwrAQn/gidPU4EUSiXnA//TcZqulcoyUop6ireDx9xqcduxdMPQ9rWmI
LoM4k7WLwIi5y6WN1xSI3KL+ekV4IhpU3t4XHUmZkS50tKSmY45cmkz7wKP1Jl00
V7rlt51KRQvbj7eacLilEb7lD/4T/D5nqd0pE+kDzPWi6E1wYa6anu1SpxZbOmC9
+ziVcbUENK0ibadRPGf5qxstXac72uJ4Puf58naNrjQVOeV0BjlX47R34S4ML5uN
15GYnZiI65V7RuYhK0fNOyHJRK8uqa+6Mf76lhX5uKsbQ3GDJrYnrbW03qy4EIW6
8To+Oeqbx906H3O/P7JzabjZ1+weMNqbXVur2l4Q5igrt11llgbM8GoXARPx5DTc
Hr6UbARUVEHzuWmy9Oe1xu37I6pOUAbwiHgePkwVHdp0Ofv13cPj7pYywuCRrdYT
khQldcX1u3qoaXcV3vOofPK+AGiVDWCp9wSP5HtVNlhNCwlXj9CTd1PUrgfF25z7
sUdirNwL8iO7rS2xfqIZk6R1cyiiZwlAs8UUzHFn3t+Q54Drxm4gl9k0soTvj81T
AB5DkemIIePEGt+J7AAp1fX1ZW6UyCztk5ZqEmaoY+tumQBEKfzDPPaTYDw79YHy
emaT/ne+9ZZH2ox8V9WtV/1AFXOcfE+rSg7WP0Zy2S7a8Ew13SSg654qcfX4yiHj
lPumrHTUnta+qcci1Q8yDdiCLfgypAjPr1rjrgexYSmMAzJ+FncdOp5RG8AsW230
JEpD9Yxx4h3KMGUqTEhT07RB6tjI4cpRUqJ+b8iUE6sft1AtSB6IR/yzAtFjG7js
s+mkK/V8n5O17+caYzEkiyEaE3LOLe/BEP2YJ789xfYnGBxA1wZJuUrk/JEni/7E
EQ28XgkPkWYE+Uo7K6dIOUiDc9sGxk3Fkjn+b5wbTOFSziPWAt+5SjqrhgcIJXao
CJ18n9gjaZFc/nBsGaZ0Vz+EgErN/HqEZiFZ7rI5v9kfMcE0pJZLn+Zh4rRkeTm/
QLlFpm9nRv4bn1JT9V9kymwZu5+WnrTm3WDBxNVT4AreDuhX56NOgNzrgNGc1a5z
g7ICimKY8xc9jxxxpOUisgV7qLOyzf1VB6yY71vUbKyWp8j6Ui5haQwtrt78+XI5
bEzqCtFzw/ifqbj53AO9boiR1B51SB6IS7NtQ1FMa32x37qD8S17PXjlWhU4DAWU
2HbVzyUNCa2OgqVHuaOVLJTSyYhkeUgJzyuaRJMdplExOC3cyV5uo1UePMtGP/Lv
zbfrDZ7ztkXtDCM8pKHR6xJhfQfcen6P1i/FnWjRGfSABQAZ1XD7h8mlIpsi+3qu
IjinpGvR+8C6elWesUxWTCt8X/Cq3XQ5+/W57EiWwPlvVeRILogAEVyC+pMQYT2A
mMtYTNsP/CbeyjiTf4jHuoS+7Go8tKEzEdU9OT9cU5CvQezxso+MCbsg+C7CMs7s
+Ueu4FfIKr8zYIu4PECgXGg/Nf2vNJJSpc/teQBO5hpzswKzj5Du+jKeZnx+FC/V
Pn9pgmr86TLxEtIrEUqnCSRvW5OcqW/r9y0u7OguBYgY31VFDxb24T1nBEj31t3n
1NdzlyIiPvpv0TqlpH8OcFsy/eb6OM67cxapGNkteaG2cJLYmrlsbW59V7RP0orF
NIcNZrB17ZezWWouyQMmQnY/ZOSg2ThTfDZ5cWGMj/cBvyblKV3ao2A5MMqP1Sum
DlUT+MKv9la5y0vkokxmMc7A7wy7T8J/9g8S2PDwet+jV5abc05vf64SEOvuOUw4
I88qDBRmxR92PeQlz4yBZ1VspVCgtGrWZJFBt754QOWOdvIJqRG4H/ok9+JsKgf9
3ulAJD78Pgmcu9pX84Dj7Ehie0gb12RCSRB/DNTVa6/TgOCVkTuyB0RGO0iXJkg5
3vBtN+bkTsVcXsFO2Sm/LLdl/TIPJw4d7WrCaXJjc5YAP3SUeiPVUmPapkQ0MaJr
SO0iNbET9EixXllnWNkjKCJK2nNKf2pHycrigr/eNbXBOZv+o0gWgkCybfHbaZU7
vX56s1w4wI+d9CUwz+56j89E48MZuSvsr6kAiQXKCtX5aNlFLhD2KugH3/dPksTb
Uew9rLjSSpCHy8PLB0Kcs2luLj9XuMCSD08V6nIkMrVMPMVK1oXvv5t3A3Q2MscO
3ec4ayIyoExtOdLh+zRlbaow6hZJqRmrMqN4WD9kaJP2wCy5eNFee7WZiq/KN+He
lWoMRxOKHD0bPIQPRgAHgkQYuwMiLs8Sr5l5Dmu5KGSrHKNK4wQ/dM0TuwpTyTLi
eZ83d6QRpGMCojC+ETwl5vioUcPGkQ9SweVrpjFi+A2uFPcMIXTL/5HuMMD819jN
hcGoEng2Cc9GInSZKRYnLZcqYUpC+84TsrUHs15UZ8Wb8PySeFNMzEyzvGz557BJ
jhp9kd2HZDDNMrz6MA4tEbYVmqf84t0n7qLUrYGJ2vmAUmr4hmRA6812DWNjQAts
uHwPCBfz3pgsRm+mhzgc7WQFYBt/MEqovCzw/Jw5ki0G/7nZxWTolqE3iHkAikHW
usKykI2q4LZsubntklnLCpvGz3k/pGCOM3wTPZxh9KELmI38GuH+7uVpGnCivaik
9Hjs6aGClRR7BlXH4kbt9IczuECf4AMhLiuIwJJSzbbRaQOBvckvRQySSzyrnPoi
dvBSsPs/0wF8+f5pqn9qWYAz3VXuUemC6Mh5Gy1C3atEkL7qkSsNgzLhRm6h7vFC
W6fm3RvtrhoDqZtAYlK3FnAZZ2V1Pn5FyEc38NVDnmcxLzUyuWzGEBbfLU0+xeHi
h1uHIQwbOHJ5qnkfaO6pruQL9XpFs2VbkAR3B6czPZIAsdjxjgUXwcPwzhzcZosH
MSLdAbFAtaWoJ1PHSr2DArWXHwkyqMklc/LcCXxWkIUHzQ2H+MOCTW5q6e+c3xBN
vXADstkTRH0AJqUwVWLzJrOeHrkOmH77WvQy5XY/Cr6ce0fueryDcM5wyzXHopPm
7oRwRngOK0W5Khj4cVwVXTX2JW5AFrsnAvDjtLpLZC3S0M0NqwaLkYywcvUkDokd
iFittr9oIWldMETm+KmAycCCOu+Wvj/HbF0p+qy6i0tiuK24JETM36XxB53apzBR
5htytyArdJq/DE6GDexoPqdTEpa1KMUKiC5uwhpmlsyOzi6lTf8sqJlcfzvja4YR
uKnXkF6CJBhU5RNUWt/7cywCh69UU92wetxHibxjqV+mdK0oUPdyqmziel0tFli3
xSHOJ6eXftj+0FKdhKt2B2+i6FMqLddw191CJLbyIIXD5g/khwGIWxX9+ZiJEhI1
rp2Kcq2aKHnF5zN9fQrgXZ5Xbnfvnws8SJk05roOOce/tkCnBmLKgHicZ/v9zFoS
poMi/M8dmNZ/X7tw+aCpxkZohkXCjWUfnadNMLA6Vbhe5IGklpCngD9rjfzlzeFl
ml2Rvd6y1qOpn9Uhtzpwl8tx1dhzYA//M9lgRFmNkuj8lmyqy6019uocQjtTmr3x
0+pXkw6nDOQw81WWJ3nM/zK42mA5pklKuAslTDdQhFpcX0b2jCx0gPY3zPrsp60H
AhSSX4YHHjIjtR3lYVX5i55Wajvw8nOMsxF4AldSthOmZPCRK+qT929jaDnmyBeg
GIlx9qhUeTJHo1pKBf8bGvt4Tcxqf5xV/5Il/lUzWfcUXbQZacJ26PB6kyMvtshs
NAeRgOtCG+eam8KNcyNuD9qzfiq1T1ZVrkV0dUbD08ECFxqr3Abfz8Uw9e4+ofHh
dYRqLaj3FMCTEYz1rq8pxfaSBFkVnUklHTYfsq4MmoaCWlKJMabzrGfJwXPd045n
dG5+YcHW9uxrUGAlj2JBFNa2LSX54VDHZsmbFbTJMUjk3dhiog/Yh7kIGWd4/d2I
tBZ9z195y/uTkoyxzFtWyiWAgMtyeQKD+qa4KPyOEkbwmq9pB7ekMG2LR/8Frl/V
d4ahQafPDdgpyoS4ppyFLC1s+uXvxTBU9sz+JAk0Pf6V2LT/ZgF1YGjv58k91ZZP
9NLWCY0Y4oRrJviuAMd3ba5M1odJjcRxmc9crsG1f7hJKF2QsnCdItGVtmLw0Irv
PfoE6fXbGaOYy3gXlYHm26BwZKu6xELI/YTX9RpWROUNGzCnm/yYMdIQMIcfIjoy
idsQg/IDN0XjegkV/uyImIwQtF9S0PYz7267oyY8GiGnA6qfwaqu8IlDagb/9Y6a
s97bVIYJwk4iH0t7yzuGHZ+CQtojWdtJEXrZPdXP9CaUYgDce9M4yGj0JlINMqds
GOo+vBJIY8uwBHv70QRLmXjWAvYlzbwoAIuuIJ6gq1QbXICXdFD4p1lS8NapstzI
w+KEtvoiErZgSHV2O6pqaHtz9/qq/O2nKTmN0H8iyxremUCRz+tnPAmk98T68kkK
L/HjEEdnybWpIdaBoMKhyo42zpcrYaVOnTU3wJ2x7uaprKbnchcaHQMUAKxAv2YU
dp5DM1PEqrTpaaKcmuJmY2nLua+cjFFFaQuAD2T6aFFrpVJ/mNUaYyzqQl1OiUvT
o8K2LRNoAe5BpLPp0aK07Mh97IPgXnuzvzqhZenCzwflg8ZwqO4/jEmyK1Zyd+/o
FTY+lc4A34h4TpqaVJtBunpRCXH4iLTQ6vWlwdVTM2veAJuE315ia9ca0NokvS69
b2DZ2dtnq6kmiQlHIxnyCek7z9EkuOA4NQSRfFxs92uYWHbqGTYo57ug/YAVONcG
kc6lpSGv3JWHConmHq8pnCmnyq8zUTwg3zUclpzlGZkaKzxpC/woV7zULg/1II/2
LiaSSujigHWETX8/YC2VZJjoc/W9y0ERK+joOrKiXFh4sUaD7f+uHjNLr4bw4U9A
E0iGOxAlNmLoyaKQ1bf+bOAGlzVGZ90+Hpma1K2WsQ7WCOJ6ikJ+oEsVqdAhlkDb
4nYtDSCXI50YjSaVp/ssmGByYdo5RMYdpc/gug2oy+SxiWK2XNx8Z5iK6Rqn1GM3
awXsYcRuDpmXQph8+RczkAapylXLfHfMBjqAiFSOQWP7NzWFUrmqmpBjxguy60S2
Xw0dKLl25d2GOG1e2N+LMh39/y90cnFaukaBQ1T1iUIepwmnLJXJAGe4WQTuAkZH
bA016s967iwH1YweKq0C4964U8qDXrfXKbstpRw8Ex2AfXhUBiWTVWdY4koogY6y
1Ttzak+D4efAg+P8HGjK4CBZbzWZXiPriZkdnUhKJkKsG+1PyIgzIt7uHHInov6n
ihQh+7WgP/k8UlsIwMK9GbVqkqT0MPDqsrCaRqDvN5sEdWXa/LHSIVgvmu/36PzL
3Pno9EV43Ixnob6Ozp3wA5QGM2F+7hq0IwdgspD0tYJPMId5C4bVgurg+Vha3uOz
MY9yRp6BynoiGWIlSiBhuvdT9HScPm45HU1M8I2lY6dAViU9Fovp3bw82KR5IYeR
qPtnwFm8F3d6qLe57DQjeON/lvctubGC6EcPti0Lpu0O0VRPoA6A3Tu/DPwyfZH7
/smVmbCkLj67jMQdSRN1YAk5JenEjREeYjD6CIPFrDDE2uQ4XmFH1jtS3E66hI9y
Q1Og0z0E9O7k6DHDWNLhCwSJe55N762uMNWWgtNHta7pGL3o46jLYQEdZicQuGKS
w2LXwhOhvcZfl0TMxX0Vp1c7cuXd/M3iXEa+mvl2e+gJmJUNyny4BdKkA2xBNTyk
tv/9FJJez7Rb24t5YM2efrp3xvgKt6u26xMIavwLmjXAYcafIHMDtspLc5YrY5Sb
tKx4v2MlTiOMpD5djwazHhGidjy7hln0cziNl1ccHhaaTwm9SCDSp+94DbxhzK+I
5giq211l6gkPkwO4PTkJ8tg/Dhfo6rF4Mhq6cI7Zh2Hs22F9/4rvjVUYwwMXJbs1
ymfYi/AsIE+VwRrmKSzKb6hPa5fYf+V8ruBZuUl1XGxjfQ+tuXaRV2ZtvpPGxQdj
+OD+H6R06xK/STjQg9fI9IYrJwJhzGZG4znYyq/UmO2KyDM3qA79Kl0fSHmuy6eO
k7ipByrPExV5yfTXC+NpHFDZRhJ0aKX40nNWnnwE7iDnjS0ESD7Fizq57+Qhpxvc
VunLkgTwHVVgQG6u/3bVSJo24iss/t3YEwr3V3QJl7vPb8faxkckqZI/h/CBJ5uo
4gBME/8b9xm5JTGGzFFtYYv0ThCF5QY5E37XMpm/P8gUJeMo5pJyB9HUwRa12BrA
7WKBo+5L4XMpjYCulmIgLEfaKwZQdowWoZkaBedtCfFcjjtxl5nCdN/YswT7c3kQ
RrGL7x/ximyTeNqoFWHzyP+/KqkfD7z93kmy3oVYmWYkmVji5DG+XojZpGFfx12M
0IeDLuNGv+NprVPbx68GR2IE/gNp4i12MQrYEn9FsOr6WoWjo/ABfmzEmbT4TBU4
UyNJywFIHvcfbui0n/itfPoeq9lMs0dHzrgyYlY33j9pGJuvDbmZ7f0D+sj6PeUr
u12/nzK5O/ulT11SVB6hJ2Ae4EYDjz8+dPqvep795GTQE4XJAT+NhiDH80K2h0le
dfpLld+LkLOlC9hub1X1wqZRIUJMEfNuSbU2Hay8zl9e7EsNd3+aDpBIQona1plf
h589wwArFzMX6tWofR4DDje9MSrnFnAAAYfR5mzMC1RQmhRMVU7T5n8JZ01vuuKx
NL9CvqcXa72We945PNZS+oZYRY7OV4pyB9E7l6eokxG0q4OYdF0prjczMkFS+Tsu
qQ6jkmWjMsuoOPzhBKE8/8dm9JA6czfqUbAhYW2sJsfMY3zq2KmHgZ/WeeRweiHT
+qEcE8TiOGgQG0NQZ4KwJUnmg7h4MXwCvE1nqAo7J/L5yOOPvpeCa5KTUPXn9r7T
OolUXYy/x74ezjbmzfi3dz6U4hfO/Yqe7sTdL8AtkxefVmYB39mwCuiclO1p8ReA
L+GP3inaY5+JNFKgn7yKd9H+6YDMjtcJqzEsCXlDYHJLB92gBMmmF5v05Es6HjNm
PTmQZ+1u9FKAsXF/MuACXcQ4s4od0m1OHrHczwbFeaKTstm9hnSADcvZurind099
+cjl3IrWDcVv5y71eAkXeUkq5FsOo0WSx0H4Fylb5EUnjWbTb+b2ZEep+ANlqYAV
csTC/qJwKchDyP1bYrbAz1h+JKpBbrG9f9EIgV1srrWTaE8X1kCMh8MjDhDAb+0X
LpBw98zHdPNEzTGM0qq7nMbdGyl/s33GsqGVdz9PeDwexXWlt0mkZ0LeXjxW0AS1
8j6Mp1GDHoJInMyr6DtBKDkZEbumySSXs8n5gMPe/kVMZ+MJfMZZ/HKbYuoQBubm
dfNBPLUQxm33HzoSeceCUV7kfTdabUkQ4oTuPo9Dyo+p8WiUMBtsjL4yijjfDj8/
ng522mSqJVgROrFsfzVWy5aK7EyeeJDB0UOYETSWuHqRYZy2P+iPFIPjDmCdnxJE
iO/4rXjpyWrjytjV78SxDo58GtUGm3qz2w01XzZoTzYVuH5ylnZP3SrqLje5II2E
4bXmlNT9hd46i+WQ8hHec91rCpm82mbkQazdeA5HAmcbzyLHP4skQWJ6vJHzWkjS
mTcfzthhtGpgmc6BjA4b/wST8GcSDswJQhfPtoNQUd6dy5fvGeEEmalNu1dGijkC
7hX/bN1MfEny+NeIoOqUQlvNYa2DnDn28OkyPs0AemwRVjMHGtj109CPcqRz1yR3
Bh5VAfLMQPLrBSFbqsLqFnVyE60hoBdceO5SGwRPoh8GcnJ+/y1wZKUZdLkf5DHt
Au/F+BRyjbfhAQQk5fn9u8l1DcEdxUepliVGQD2jcCiolbT63Slh4IJAxmOn6jnP
iRumVK8dRlgSNBUyQgzs1hKCFVyPdqwZ6pu0BVHswNqiZh8ChU6TFIg3pq/lyneX
/vqnuQBqzvYF07U0JUkE1rXDXbNyCfHSCn3M/0UvM1jh+B2aV8nZQq3D1/Y59mQT
YPFiqDDhiVsKXtVXpJ7rKSjmXOLoYk+uF6+sNa7FFbOslLOgan4EY9/aeLNlvEH/
7+aOuWFvqPc8F4ZyxTApuCM6iKTc7EfqLBmEO37zfTCsIJRblwZOiew0KwTNaUP8
ls++f3wmWHMTFBcx3tB9NV+0/D3Gl+EMwfg7N+aGzx6Ro9s2dEhvULe1AvD5AJKU
ZNvdDOfaal5zj25ZL+FphHjnMaPQ1SKuoQiLGrBM8GedwTZH+VYY3zYHMKdqOZfm
jmQRDNKmHlE3W+C701lDMnkkUwLawf56oBBsHUW1w/CoMd9WRPosEVEHPMfdXHcY
3qcSbb/R8J9ZfMWwcEc4grbRdFmUdNEKTNT1LWghM5qr8az24QMKlo/V18ZM5RN/
aADs35Uk0RxJlqJNfIooldt/kMHO860zapmPJ9mYvJDox3eEPDuLvfVsvQey7NP1
F6sTM/HLTQUbMV8YYzBtfpAJ2pDz7F0lqDR4IwoZOSPDHHTVJgmVrn/j0omVO1WB
5Fpt56BGzJ32aUXNoAsf+eZHOU1DMF4nsuKyf00JNtYrcKLp6W2Nd8Czb4Dgky10
tshwbGidfJi59ngGAVq0i+hI9rzyVb+fa0ydv/rZl+3ax9ctVsm30HyM0hPAwe38
GfyPhr911698LbCKlXjFJOuf1iK+SVeIGWXQVByxqF383egRpd1i7wkSTGlOBoxW
6SPDPi8Nf3zLJ87WBDqvmMzg7RyGWG1BatamoYMsg/061NxqGJ6jvQ+nCgHA7/Fr
Y1kh6qSI7OifrkZJCpk3t6OXFYxE+3S8W+sQit7fZIC0jMd2X/dLhX6h2outzBzq
nn1Ts8neakMWNjr8Q59D4zpwo8qhHLXyJsYiLJKGs2HjXWn6KKNVbvRV0SFfjSCl
uK/D2UAxxBTSd8KimlYu3ZFgl75DdWxLOgFKZjmFT7DZycJTqDS+m1K0GK1MXP0n
DKZEDdGnEbHM8RJbII1EUIWvluoHuxAQM++2YvkYWzJrbX/OV43SUS8bIJjC/uFe
bawU7Smk9w50KKtJoKx/suU0BLZ6nSmCO/jSgPicEQsRsXpOTnvuwZwUcQ64Xo/E
5jzdoAouay3FcyifqIMI7JPdWChVc3KkKc4jmfbJzd1KQLLClhmtyruBxuCdzLS2
rVxXjP0RkaDxW3oDNVva7hd5zaNzaVkck2CYWphHoaBm/MoWeDLyOpxlb4bwuo/i
mvBKb0sPTxBhioCapVdByVoWceO0L4eeEfQKL+p8VcAYvBnLFAkIt7nKoKCCzzFb
wCbCFesFQ0qIDkyHz2coMKN6RAy6b4sw0gE+KcS+ClHRb4fB7JSRFZFBWDJlMklM
F1tLLxEhYoldAocHdUXg+zatKesLCPDNxtM3N8wvi5FPubByUtGoslTbRNT0IyP6
Kpu6CKy+c5KR5iO7n/7kem4D8R/CUil8WnCLxuWOm0WHWHYdVMYAXYAYTIbg+FNp
cAeSwUtasy731q631r8pw24tCJmM/JjMRFoSv4hHUqaCQa6SFnTuCjY5xomhqf4U
M0gsyjUkZdQRdVVcrzcIUB5CKMn/XLwHjPkhZATLxshypP7731nUkjFdNekFsztg
gUgqG0iLbnLMgs0ppjrK3OMdss8+TsMQ48PWsKJ1c2keT2owtDUlT55yIRKO3XFS
A2SZxZks6AxTSQkM0m5Fa+aJg7fo0knLG2V909s+0NSjafrEDndhn0sMUMJMuMI7
HBNTdc1fAvObsh2U8MDXpctl0Gh/yCPPIDCQJFy7qXxBsbtAMGZSVFnSp+MyaMb7
KCM2K+pxo15fP8oKr0tJNxKQfzf5TtPiTrPr0vb99bJ69lPXdcXt67juM63QG7h9
0TsIK109WDzgrG7wb3ZOXgh1nbjzVJ21NeFoAm2jFqkd71ZrCbZeux58kJq8TSDZ
LPLw5TvegEPDsn1KoEB2qkYcTsq3LtyJ7+iSdHMRxymoVFqTtSi8E1Q0iR4qGaRY
PUw7chfLZR7UhCr2NcFe5MFWuWVu7+1lOErNJgJJYj7r1bLtafA4WOt8tCYSucHF
KypPklmWWTQVIprTfCX6RyYpWY7wvide/1yXoAnBotnxc8fnNSECNH21yBCkIWnS
tDrGplWOyf8XLEHVsg/66yM/UCsGZTEoeIuSHch5WcoPcwW7vfJYaCFkQtSgSkrS
tV+I8lYqkUEHRoWeHXShw34hrOLicGDHzaHO8z1+lF7RgZLf4IDbQVQKWo9GBpwz
SkHJETdTMIzd3tU5p0HW+7dPbQiH3wmjCuFq9Zdgpsm70NSgXk2E987KqX2TUyc6
BQ1CesVyZ8QE02uuP3Ew19bV+QlC3WuDfa8co/fyy+qbIPAYznnimpT4fR1jf6uI
Xn3onYdIF5MLLKArbo+PN0vWpKC6cFB1yHtXSSA2sm7JeHRySlPlr/JBJa1L+Qg1
ZfpLJvjPnloAweULEDMcG/cWC/BFPYE6Dcs3gloDG+pxX1A8m7wpW7pmlv2TNBhu
ktP8YsvHbVewZGo68qQSwtX91tXOeG3J+1WDnliVoLkP73uNk+dDlaXkzxH4GFqA
4EKoS4rXr2C/JaCgoF/M6JwM7T7S9WgX1y/bQiE4xfGZ/2/j88ePKfWhK7ylHwU9
VFR1EjITmiOjA+9OcDmAJXHlXpsz35AoYVDf25tZDf0oNhPmPa39v2Rgel3K1QTq
dfnJvpvx8++BWWihoowzh+MrORSaZStQV+pFD8QzAx9EUa4Khv6DaApqXrOhxYfu
v0kbxtiYFfVy0+l6YAGshngx/sggEn+aE6DiJfbKs5u6vumd7ATlsvgktTbxRfn9
HHCOvhSoQ99CA4lKsyShLolaUrCEz/1mxSXzL5gnbtZzrvna7cVVW1j17ygk7JJJ
n/sByMuVTwWcHJbwf8R9DbJBaouZZzkPSG6udbJ5ITjqoHclibcvMMmhmWCe0VFV
kBO0+8p5vcmE4vU3uevJjn6+JWT8EN/BTW/Bh6Lr1JPcuSZARk1nzk/uZ0jwHR1q
DjfzAd4sYbI4oiXiM7fELE4qmX0Q/KmP+CbbSMvQLeLQs4pFIRPdITLKJZ4zqBhE
RhTvWkvti0tmWCsoqxBgOB9XflF5PQbHu7WCXzFaQT+Z3DOaLht6cWBzmD3efnBn
jMr6VjPNTMaZGJ+aGD71T4tuR47nJtSrnwW+W7LrRu86GWYOuolL06aqcdJjUqiI
n0vcYhjF+katAucomg1P0wAITuifFEplcnEdPP9YeFdct8Jc0zvhRqAlfHdI40a/
/iJQ+Lwxda3yVvPbQ/El2JscSP/DGU/anUTvr90f8AQ2QNBZnCLbSAznLmjqtdHu
zPkkicgEOC3uT5JK+gj0xcQ1Vhf+/OzIT5eRdJ5rWpRmnB1k8NYVuWf/QvfCqaIi
Unw6RKs9KPUde/N8vl63DKS3u6B1VBktixsHo3vHRxSqrZ3kL6pPmw6IrTSxAviU
Q6w3WXWKALdLuSklr4yxYXyl+3u/FUuBYMGZWElHgecabKubLVqOgIC2NmGHP+d3
puexAZ/hTBffCLaty7+h0mxiZz//+jq0qKt5KuTkQAkg+a4XKd+3o0BAWE1+LvQ9
cbd8V4FhyDCdpAnR8/BHPKWux3OERZBVVf0d+KDVx0jUjHU2g5/fPdjgI+/R46Ea
/TCGiWaFVesQo6InXoHgSpa2AIaA3OaTay7qiQjPj1Iff6h9+ahKv/ORBkISakrD
sLKYu3hN6ByCBMyD8LMEktOv1Nr3NIVy/MAq0mFcwnsaDua7Tz0XSrFI+RVue2Yt
3YJU+Q69sC4rOmyezBpj+zmbqUbLhFQ2Llk6rb46cpb9sG7s5SuMfzSf3xazgx+G
QwvnojqB0wr5r+1HEv41NDxI2ZiJHB2T7L/kn5h9VFbFhDM1Sw8QUp7XNK2f5vw6
yiWt6XUU0vMJgtTWKFqOdcWM7RQIQPsoGhBTQ2TwInrNlWZKpqkqltMkhgC51Yv1
SC7eYUm1R4SH1rE18R2JS/lffV+2x8pD0bRBuSTX5RlqPhjdvPjJGGsKgNKnu6ft
lrNOBAkpPZNTXucU2cLOEWz544LazsuXBQP5z0DfaNwyK6JY5x7WubxHRCZUyuXv
0tdGwRRiVsuNZEkLKyitZ6dKhyGC6STmE8HxNNiz8jEYLgRnTIhFhKw9njjDTpxO
fnApCtRT674a8yKJp+qlGG39GdkY4e8ZiNsJIXRqlDe+bd8P92/AsJlsIT8jSs62
POu+DmTiW3AhikMhkUPDpbCSExBBeOOJwN+srIsB7r9XCeY0XFNBXsp03patwvLg
lQou5fojf4ibZVzZbBRrRoLR5Ddh4EKbvoCcvUFkt4amc4G48C0Y3lRW8v8t7hiA
CF6Zcd9EfCHWy92H+e6TU/izvRFxkwIrysnYhif1w6lOBLuOK8W/TJ0OX7CgpSmS
s4NGy3O9W7ECvvq9I1kM7ldto9D8AbJ63MN3hpdHTqg+oWZ7m5rMQclSJ2Ov+1rK
hn8VIgjTLBPtLuQHg1kCVyYR1sJcgyZwkDpdxQ7KzFnC0SqdxsMcbz81v3WqGUKW
NlLqYU3+04G7QOOLnu3D1tTGhTSZ8OvHNcNdy8SrxtbalDI6ewKj4UBoNMrEUfnJ
5yhxa+DajI/HhqdBxM5NWyXRA2TwMrRIZzAz4scKgzAs8pLjx17/g7+8UbsIiRsC
fejw4LOHzzzrr7T8P0YRMLdaoN9KS3pqXlltPOx5DpknyE+D41ol1WB2g/nhtTuW
5B1yqpG2RNNMoXi8wytsVjKsMJtjC+iPqMHb6dwj1FZB4FNsBpTiNaDaNzoXCfjV
U01qObQC20HIH60DPwKHRd2Mzc/FB8277UOjz0yQOHnj4dd1pFQ2aHpuvI0/JVc9
8Hl7isvsAD4/yPh2Lo3rdPr4FpEIfLdueifEW+FSAQY5Ger2xf/hBNNBw6JhiW9N
RAoxz0FXkmE0SOWSbmK+7SbjSLTZwcVrZPM4gLgVwLW4W7g3mFr8ek5fm4e93Uyc
LNOs/hSp5Uv5UuW3PvLJVXmoETSOryOZXm5QEBZGALQDerWlpqqmGLmTVzKbBe/j
v/em2KRNPOGJlmxar5Zt/Sv6gpmll68KwHYG3F8vpzsh5T2Kn1hwaSgqIZMe476g
CaQAZoY/MGcNiBxog96k/N7XGiqr82MCumW69emwALhJJv91r8udZcZO02WmIrrt
lXhXL9i/CPQcnctbH6QO/8HSg9/9prCK4OIxcVsSqfqiEiJsCNeQgCq1z1c4fnjc
GvpKFwpnFN3Y6ZCLJ4la8f1el/JcC++eU0zoNeKiWlu48NYidxgptflkBsv8dvVL
sM/y7A7DbfA5rh6ev0HG+8ITCpooXPUxUP36ryq3NRPrEWUEkc4gtbq/xyV25Re0
ZkAm5qXPBj2BfOPB3ReXNUbxs4NIDJMFM4XjbbtjSXtgPLAVGTebshgdqQSnuG2L
F9GWBTiOVyfzIrEHSa4vzWlL1rBHot/MdQMXHEKUThEmJ7R46JqEstLMvMVaRjpt
9ORpGcWA860W+BU7YbZ1wIZNNyRBIyq0C+e9zFqt2+HvOcnceS7tMgPMA4nrqUJn
NQamdRCmQlC98WYpu1GnKl+9mj6Oe0r5z2XeVbogQV/vo3jHGXBGlI2Lb1SMyiAw
ezRkkplwFPdRTNVN3CuZ9BwLw7wEcwhNVbPJZkSBxyFZRCFijibY56+nmijWbUU3
xupCY7BVLHGzE55W1KDAwHDby6u1xUakTaq/QKJyCUaRXZh0vmWgKcDwERzQ24AO
lTneUnKtLWtEJAnM3PJ54+RF2YephiyqD2h/aZ71O9hwKADe6NctoHqY4yNI+UGC
hgfAKXpLzFYVpCV0Cplj+SzG1o5z2DlSVYx+am3OYukCFI8hx5eeCkLXT2f1ALbs
wEV0o/mkGjC5Bc7EFGjdbMt5kN+W/vBnF0/CMBLawWf2z6vvJI4f+wPiZm/WAK5a
y/EaMek+sBZVdTyAbvHhGlyRH3plhgCZsRgm6+1NJehkI2scJOq1JcfR8u/VZem4
6hX1kLq9IwoMF9wYL3Er7Uq7RuBdxeikImj4FK9cuRZOir/VUd3h2t66srVbhcJQ
1UCKTNCpg8tZ21Yteibc9f24xU9BUXssskzNGSeMGg4fw32cxXvnqgoY6fRNEE8E
zUvdNI1PeqnBl8Ha3SLQb2nTkOkKxLKzz43ORcaXBDYVeCR0HrouoVn3zQKs/Y5A
NzNHlwlHpMIQWieXMvL+HdMD+ovZqzx/vmuzxQ8qKmQiX+NXyr6XarbiwWGMcPi8
zIpctBAM4un6Vn6xHMwplAY7ovvNMLp8sFqTpbuiFkZ52CFLbvW2mwXIrutbTSY8
aolpfshyYxAUDr9SDPnvAhmLYjyvnhqvmbqq8278RMpU2wt/MCJc52Z9I35EDQet
0VA8Cm9kDkPteyEgouGXkMI7ePhXjKsUL2NPnQP0UZocLhtKA4Y1JO+6x28BBvir
iNXC4IfcTEcDUw0yCr7nUfgLAlSwhBmNDBBNMnK/N0uHyjFP+Z2KbvY+iakjHDJk
C4rahtuTa5lUQpbFzH6tCECKnEahQ3OvQWGKYHJMj+IvHrcHUjeuX37ne/Ta4aQs
aahef3IqfTsVsrF60atYWITC+vrFE7cBVWeorv6Gn94429alPrvdXOGsEt7YBbjZ
2+Lm6uxVzNJvGj651rEz540j24HfzOz/mfIb1Q0r1iG0jwY7uyuhGjb4Wtxq6AFY
caH4+u7WwPLwrWOnT+dVOG1mMhAqFMwLlL5VIJN73T7f1mATPF3qMCZEX2irQ38m
FX2ubDtedu+I6C+bvaRHhjVLUWfgeUMBp3km0GyDB38CTm6K2eSC0zqj3GK/Ru73
fbfkvzh3em48vXiFFgpnqGRKgIEPPdqhSxLVJgQND0yF20+4gea2+GErwO+99Ge9
OWFFQI6lFJpOk0HgQRwAAKojRWL3NOp4iAnBRuLwvgRqENd4CfzzfY3SeS3OIJoP
2xUeiJ9pguVvUn2aqEwGzHwEKpNsyNgOsx0mYHPuLP1QQGXrzzKu1mQGl93DhLiB
xVaR059cavkDINcwaSfq3/qkUHzL9MZLbuy+H3+ZaixTpCZK77xw1sACO3qeblp1
rXor8afN8aVxi6vtP0jwjWs4MK7Ve1Q0l4V2DwGnrIu7XdDSCT9XnUJoyt5yqS5d
LCU47nn0Wc+Ir/C23KgjchOrKcBioIRFGRFCHdSMtzmLwti+0GX1yJzZp9GS/PRZ
oA3w5G/EvwgJyFMJgK006lg7T4DMIg7JwJqC4Dmj2BpVthyVZdzKZekERR+42jp2
V/WEgOfsNeful/vKRd14jr7yG8/C1YwF5fuhzDSgrUnWor3/+NzWlDryLXZvYxOg
7JAkdjFKyD+RyeRLXTgUfUGjuL/Qh7DlIGF2OYKBSoziV22Tl61SqnSB9nxuE/Tg
/IFmnFxHvzG3smyM3Wjv4ABG1nXXy5vBzWREKqi0NY7huzwMcvLreiR2krEXBGUz
73jz6qfnwx+7gn+G8A8ZeJGtsafK8yPnoZPI8BjtugAeQnCDS6nQaznDPDhLJk7i
lm+rlAiihqs1AtqBFu/zYwdO/COW2rPWakhNX6lr0rYfIIIvSnz58vVk2rc6faxP
HKW35VuTMTkpwwbqVVhXo6iTFUdfKlNoiUIzSFoPgz78iDItVOF6ERTsgnU6godR
Mpi+oOc4DiX1lgOqXXjKUp3swXG+vEjat2w6W43l7b7muG/DsrCTCUnLcgwwreEV
fYbS6UQODK7ru0Hjs0oB89M8vZcJFeUE43Ui28cFFd74ptb5y0dY82LFGYjn0gv5
8Dh/LWP6g08JtYNjrWTIqGgjCAawKAk6Sh9Um0H3jhbrAmeP2q5kuygKN1Km+IK2
Rm+1/P1ER90MD+Pdv4ObZ4NGO7aavztct3unC2i0MpN4dSEEecvpF22Xj+ASDDEP
QmiVkWw2m/AsUU1BcX+AQAb6S6xNj/LVQau/xmx3lBd1C7G1qog5Fj+D58ge0U4G
t5qknoAZ/XeC7oztv8VvRNUjKNY5VSqQYqpjbJlmuJn6knwH8qfBlKqzs6ohfylf
NzC2TXKAxeOFVVyo2AI6tMY7G3limD0X0K/8c9rrHi+m/pnd9vE/cSX0kb4vcJ3I
lI1ub+UDDJ0Q2hVA5h/G+cJyuK89ACeKA1qSWyi5Xen4Ih5KRprf3iD264gAnFEy
1SPRFISOBarWK38FFVSacpoBhUV3yoxVHP1lZCwnbg1230utqGtdpywKqXlk6ZVs
YYrH22tLaO4StGGnsHsVSO+Wqqe4TDtdm5lPlNmFOLOY3x0ABrmWU7XnIqWztdnU
XTb6JLbTGyMybh1QS5DzoqrgcWONld3xF0fw/dkj7wGmKrg2vPDkgCzg2S2Va/qe
L3dTVE8Ufd5e5W8VMWWODv9dlxSv6mt8UKU7dhTT6Jr0QOZE+6EPqJbP6hwBfcp+
VxDu3MnL1+Qq3TzQ/OEqlWRe57qFf3d6yn4RX8uMyl8+3v/FZMXDvn/ZG/wY04cq
6cL4gCnGVkut63gJasgDC7yWSHDq5KlDMoLnB0VEtug67+hV1fYunjfxI3eNURq9
QJ+hGQjOuY/NDO+CzFzgvAAxhCJt9FNVZpA4TFTfikmlqmajrHL6YYzQInrGQrHn
bCbVAyLdCCDBeYBCbNmC60qS7y2WkdrccREBaMVZ5rxFS7hlxqJjmVaW1RW+SZIQ
Ytmv5QBjOuVWfl50kbgYM8CfkEVU0SshmWn+h19YTbs0LhVWJFSTy88vC7MkZrz7
1gsFbREqJwu+lANdxB+gjlTtpmVaC4eAwYM6DTD3vLSuACrUtvIxlL4BkZS+jmpY
jFBJgBDisBYF6ywZaTRosEBtqiIyC5o9Xf1lSXfLXLXuwOr6emxAYVIQUNX8ljVh
mkHinfiZ25vdBoPfVxk2uENYhxOW4uU05utbEsEjYNTeKzUbgBvmXm/230eMHCf4
D9LDJ5fDvXNhpqoSIkxgXlRBRrepI5hB16B2abvxP32eyLzGNoovNbcquRGcGWG2
LtT375iqPtzpin1Az583dFqTt6tIVVwx2Kp8UB/KD0npFK3IviZE7NJrQIDT4wcw
B24jKCiS9Rhv1bIE8HyVTMoG4r4flu9SL3TOR///RJq3IVxXYRSAb+/FiHQFZ3E0
RKFqlxYD8qXXjqMJo9i5QEuDQd3c0PW0sqkqhpQi/nKWMvHhZBmS1CDWPbNphBGB
5937U/YdI6UBA61Lyh8zd33kX9lPLFFgKiVwTwg2M2BL2xbUexDKah5cZEjBEoxi
dS6AmtMlVCrFsGrETjMblc7p+YyNjKxcMI6RMnUB535xK3tUX1ZbiJQNutfvQuB8
x7RFTB7GSdCtYMQFSJ8Agsll/1KTcZsZdlkM7mzSO6hceFnFc3bQ3q+x+kpqSrxQ
Bl/jhwgnfkY1VA/Y9hYYRH8dc4s4hNPPh/8hou5J3HgktsLnDajwYI1ULhW+MwBC
rObLTELaQopgDUTxQCeCchXm75rRLxM18+Kf/EmHngMV+pSJaVqqOyTHQDBFefnj
7YyQc0V41uVmQeB55gZ34AIBEidqj9FoGvcdkkWwMfOcOS1jBwbIYuzUMI5eLAp4
4yOaaRDyYeN/AkWKUFIhHE1HlQmZIgdka+Vv78QHmCKVA6NsbVZLfKWbmqbGlzWk
UeSq7rmQe2XOybNzKwctwxK6QYxFsqaLddI6pIy5d4kdY/pePZ8775He4PbVuAuS
8zGLPAq9sR3LfWES0NW/t5X0MOLZZbKUyQ55CDBBtgJOWweR61Nrsq0pMu5rptd5
V0DvzUTClBYsBRFpgbO7PfgzQ2sgoSTgf4x8Ow3Zmnq/HmesEXAgdmDPnKy1XI/b
sGoIV0myUVUyylpFYEp0r2erSs3wHRErdbqP9vibh+q+TZXPtjFgv8fzNctt43gw
8Q+g2Hx92FWxQPvX61tH3XqxNxpWs74bbdn1B0eFiK7YzgC1VAbz4vHouluCiRW0
Bp6r8APO0xQwQoZwHkI07Hbcx4+7aiX3uoiulE+iCL1g7HccpvNeOKl5Yf2xZNSw
Qa0wvtHeFAsN1R1DogqlPxMd6O4OBEdd3lJE0CfeKQuSfjAVJz5/ZAfzc9Pisjsn
hwb6L3zLkkKmu+wleKDWAdEUdovfi4rIUR+f23/8G1kxndEtyoBjQQGHMqh1sQ7I
RNhGtFafZPKL+HH8nDZ+/1aKAj0iYQjngWM8u3/jXEthQaAVS53sjK+6gR7oLZ60
36p0ScZVlG5GtnvaIKEUdz38bfCG2ScHw0B+XNsS9atqEJAnzBPWJmZ+NS7KaABk
CzzGV2OPh9sY8daD/JDZFeIveeQvbtXsN28xB7EACw+F8HWoIsKH7YiZew8I8IRk
njE/or1sk+7fabWU8fp/BV0wGVebL6tDQMcet1aRwo46lV1s8VvPvl3ExuaSmywH
RfYjqS5/beLDTXyakL6lzQh4SfWZ46pPR/UskVAdoKSxsxbkZ2xOa/9EB+yhNKw9
ToKO8LEB4pJQmHA5rXPTo9GUhdEVsdT6m2CPse8/lNLSDXZm6wsESuHkMEdJGuUm
erBbepOkGnVhhq+moJL2ZdJy0o/XM+392Zx9peqtJUMkJl1nET3UdGWk2Ds0n7au
K3LS8piLBeUwvDYarN/ZXa4NWpxXefX/Zq50oDXcb+52jdbYpRVpFrKP5cY12ItB
KqNNRxquzslMCp7fDn6cHtpH7FaeHZhTncPdljFE0775yaK7lfpSN8wB7XvbepY8
h7P3iqdQvwP0MtBV0trqwEQpnD/99cqtwxM3oBcyviGshBNvA675zRfvYO1BWnnf
Myqfs4vh0AhpOUnES8erwxyWn0CiElJYN5H++55JLiJSZbeT5oNv0Cw64tWm0Cdw
RwkzuKr1qC08ghxziV0DkaS0TBIGFkak50aFQE1qziDAg4+S9q9+oc/y6zE8FHrN
z2GnhebRyPN8hjyCCuOiNw/Txuvb/cE1Lltq9YjXKUG93pgP9sAfdzYPMsOzL681
fxrP6z6vf8FmyBJupu8uY9i+XQdnigQtOGvsYioTQshyiNe7eQpe5RLwXAbtQv/T
Xp3+o0vPmHEcnEpzBRpYyTWWKHebw8uByojxGuQ0WWyuTK73QcYnlFe+hbvabJvK
3zEZwjz8UbHWmAGoGmkkO54fNblG1D+EB+Ca3gnE+K0ld0s8mSosgMf4hiJdiYaU
ZivWwj+ymG300HHK5/dcb29E8jwD2AsSbrWQMvC8GylHTJC8OgOPqnfWCaar/0fX
b7YhW6CK5IPZUIa9O4kVco125uZfJC22Pe5+I+rCSyY5dcEfTcoQDgS8JEtuvaGo
u/Sf7MoiW4WGx4nYiKkWGJpyJT/R28AYUp4PED3j+fHgM70LqgmUwwVXYDjLL57u
EgJQbem6nI6LxGedp//p/y4GMrvu5l4kZ45MSCJDYCra2YsfYdAME95wQlbERig5
epCWrgu6iLDNAacHBYdsKK+fDfAN34n4LbphTeomDQhANT+kUCRqhlsVmSQW9MX/
mWC89WhHxRuX7eF0phZsK3WOFs6aHwvpqhrhv0nV1iNISpKW7hgyb7p6BnPpk7Vk
zPQ6fk871GCQOhcgaQG5pM67VFEz7JVM3a9mx0FJ7O1otHMOL1WLN4QVBJGYU1aE
IrTgjsdGA5fSo8iH5WkmIDIi5AzeOcGdN5tSH0uSy5KVu+msuj3GGVj3hUSqAij4
v/Uq5Gc52+1R+H1ZiHZeTGmYmQ0OWD8bqmnzPo6I8Z11Nc/HqUfm9UlUbWQU6DRT
yNziWfAZIy7hY72B7M5KgpPIiX6mOR26aDKY5MrQqnd9awvoqJI5OlmTez1PYaOY
HZVK9HLJLCSYHf4KgHa0DTLk9myF0zngFw/9qHR2Obfaki6qIYVF2lppTjVjtbSY
xf8IQavIVaxEJ2cKibIY7tifL+IaviTSViaG8dYCbOizX6fxmdf+QAuZMjLJwc84
pMshSH33ADSvBbpuV1OwQM01mK5c1LYh42ViRPiPsYOdaWncsowacFZHkt/Y8TTT
Se0yUS2p7X4Lj30621RO7Ry6ac72wLrhmad7RTYk0Ju1QVi1EA5tenDFh1VToPDY
pFctvuf8istaVcrBD6cYyb0ddxp7EM47JLoTAHkEBHnb8tw95xuFXFoE5pyMOlyA
v+V2Knku4L8h1v1Wu3K4cjwj9IrOtHOFqUpy6XDP9e4rnK/OePmrH/KOD3m9yndV
zihJma6FKV8N3NfUb4jtHiLeZaXX1G7nYNed9kYwtoakP+ZHQifo66qsj4EM7HLg
sD9z1U2mIeIsSot/aUv/1LBYnYQ9BVy+MBbouh7b1jID/NsxAhT9EHO7zAMPFZgI
3ikTV6lEId2ZfAshJapVZP0Quup4yT/tsR8/42VpwPCIwnjUpeE0Av0IeKwH/WJw
u8UtSlpVpSUKXAUONN5tD7a/tno4rHXhPBuUj7BAarlgvIybS7LGl1XHhSb+tjw1
fBHQg4rkdwj/KnyhXTyFfi0bBwQKyIx/EEJf3HbBPpXXA+ZBLO5q8CwLNX/EDAxR
UecLzV+Rh30wAz9rUwtVnQP0zcil+5QP2fGvR7l/gCfeFRZXm69OkZDPvDL+d7tz
IGJuXv4bNggCz5QA4qGnVJYZ0LC4ug3jBmL47ld/5wWq9mMtbWSSIS1edNbSFJXS
ZmoHFF/9QWSUDk7ZX9Xuuk/CHbrJfFbe4JuTLm6Bv4WrYk1vwY7aUU5velQEk83+
vZJSC5qUSSXl3Kk2tfH7HrqwzlHMbDcY1Qmg8neUuzdmnFNX2ah2emeyxpycnlpu
teeQzdA6KMkZrXTMcGT1wOgmj567mm4ZhSZ6JWSPTR67uzTTdtpHut3sfuynFm5r
ag6GDlLN2kAhykX4V2tifQORBlxbpPak1sXc5NfCZLIiZlBvFRfqdrk+5k+xighf
EpSuWPuRJkjU4mwsZIdK6GTNpaZbzClWY7IYKgMu/bboqjmfjJYFC3xB9G1SDCMt
CC40aVpWmhi6O7pzL7dJxMnmkP17Ug+4nZ0GqXacIK19EQ/3lB7oSvvpxQtS77Mi
lzM0Yn3aEXwR+knzglPUU+wZuvaprEC1SOh64aGzhC+ea3S3xJMLOLRi+DLkBKeY
oXfsKG0lg1UprtW+lzsHnYXZVRh29vsJ0pZOM9gh7JfcGs8mKfk6iWtzSxPzc5tf
nTb+nhAOVSEreDPmLISspvowRrO/J93K5teqt3UM/1T8daUEFBfTG2KyuMlYYnYv
pK0Tof6N0JX9YfZ6SdCJDlSuQ0IIPmeINqdmJ4X/RiuXPnjkLG/zVCiVAYorybPW
LL8xD4WwFp9DlBchXoLMcJMQ3rcAy2z75IchnFYoeYgM3Q6kcA5/ATYjFi22BOsp
kJKK5W7dItm/TzmWy0BFRl3okeQuwCt7jOCqQ+8DlQI0WNkzB3w4fC33G8gEN6gw
ld5b/NJIhnpoNQb9hVXlwD05zLSje+qItRR6soPHiQzivw/bQG3T73mviv4VphZL
9HVljdoxLBTd1QWvhb7He3tN1KpBKuJl6l4yEEjq8yXnubDOCaATmtxXMXwixa4d
dWZJ3B0BWKBqPGUA8K7tA7WAvVASvduwleqQshTf6TnoOzdJ0XsKi/h4ZGj/JdHd
o0qAwQLWbl9+9+ks1RSGt10f/HUHMju+jiqatqlxTPmaxFiXp61oYjfkv3LwuEG6
7uxorbyORMenQBV3YvGBkfivevbp1pFfHskgqSSbgiM7awkM5ug5M683+vSQIlLL
h2AlIdmP/SNBHWsNwwINNvhw5i0JPkrntNiqn4s9E3irI/xZGHC6yiGHhyz5UsRL
tQ8S5Ny/8u6aR2VAfmbMDRBCqKmR512vJXTmqgGangA56Y9QYaB0m1yZDODfQ0w9
AvTlkJ5u5T9MELAmyu/d6qNe5QHxnP9xVfrFXBlgHuzjByEpe3htuLqKsvApUsd4
tJ+uhnbvQ1G1S1FhDJf55DuHp0mE6zCjDmPQ4ZpgeWGlY9MBvHFAJ8+fuoPTrkRs
jrvwzJl7lIe8iX3m15a/7bi+EKKAjbgMrUSSKshJSwhd+8Kr2oYEXQtfunBLRJ/Z
KfwkbzLdGOM/L3DaefwD70oAo71xpfC/VxXocRLYnvCUvKThdIVWYi43uyoEFFvH
eGkv1pNBzZu440QDu37YBrgmq7gTG4RmBOlg0f1PK/X4QqdYkmvZh9xVOg8MVUKn
8PqQmcnULVvTbxnn5dS0E2fDJwdVJN9xYKrvLkg2wQUrJrA+lks8W9FTerAKMJ5u
lzMQ7S1KoukJ1IzDNQfJnNLwtuaJqJpGcuyhU4CmSFzUimyGqtIM3Zr83RNTz9a/
OZN/MuxCDxEsB3gNZgh7sbWgCtUWTnp/hZ91/tb9RBXNy+4HbPa4M4kr0LCs+nKl
lbk6bmdIi5JgzE4FdBC5xNoZ3m4rZw9VMp9JyWsvYzkfV9EkF5/YEBL23+Z6VD6o
QUoO3cBexxhyLHTLHgdhhNnzi0lcgVLlr4Hu7R9/prfh2lhVSev85GtyzN0e+ear
ZbD2XoQ7PEX0FU1jttKBUBz1W8wYYc3zb/kC2POXbYqdj3nUxwRfi4ayySWcxWUm
megkCegYEapmq+GN8HAquj+6z0V3VoUehBD8OOg9SM4OccckIsLAJ+vK9PPzeGfN
WBZ+cLGbq8ujJTs+qMQqlq0ACzX0XltJa2slyUL0GpCbLhFqgvh45bqsFqmdHDA9
cpVoXigJmam47NOvpT/Rxcsbqiu7pawEoQcKnhBoc6b5hkYlgmJnqJYP80Aeps6i
j4lwZVNBcHR/OVqs1xa510RJuPxQ0hbNB8ZCjQ9qt7yHhjICXng7wR+Oqw6z/1SB
BjDzNFeya5RYkfY9qBwL/0iU+eSMCEkSVS2kmTt7Ix/x7SgHHNEvvZkycN05vHYZ
frYkjT52ImMNAfxH4iwoU8NA7FPBI8mYeVqEwSc0Jewqkst9VBbTSgtJ6sZQ7BSD
BGW+kF95WuO+3QWAOLOyZvqtotT/Pb3GZYSoXks7rxj/O0cHF+GoOYn3ZNJEEzrj
ehpriLV9os5pi3g5P1qWifNqCAvVlVUktZXOgVHidf+UZhe9f/8eONYftiEHqylL
Hr6ySXKBeE/VKH+SM9ipcT8Nz3riHDxlmQS0PasrIhFHgpMaB6+5LRd/ygvpKTh1
sp6ED3M5FNBXf0Y1ZS7IIclV1EHVR6p86nSfIXjJn52wL4whjt/BGr9nFP0OLuD7
qYBtTJ75VZiBFqNRMFVKCCucdFGUK2XWEdVwtIsqqFWEYszhzFZW8fis0q97m6es
DRY6nwo+rcsEBdoobP4BbFKyTN26ilkbqPe7s0EAQS2kVHeCjFdSYgOgRqotmPM4
EmobXsVgyZV6m1lGhMb1318JnjEMf2pfHQVnw3NoAWKYXcg7oIvNNwRnrpe8gynO
lLuTnky6UmD86MwnQY9IHHGfElYF5zlFmkT/M/CGVyuPpfOZ4nIkiTlkSCKrToEH
iD8iB9yX5BIiTrYGjpScJ/AcSaSo/2lGOTKQpzcLaZ5WDAK/A9kQfhHuzWfgq2xk
w9hay57N5Y/pT4hHZWLTkoDvEdWJl2S2UIa8Dcvef/aeVyuOxbPzhWyy2eQUXS/L
AzESiXPM6x3sIpGx+DQO7FInDw1Tuov+EDvzNlW1hbjCmjN3fh+q1p43pmVuFehz
MKawO1GHAH/QJ+HbaKv6qIRV7iN2d3OuvFxJoSgX71xFrp70bOhoSW67f2fGSIgG
pxfyqHUIpIdn7bc/PIPvUpfIX2/CBfNkt9xuBdP8eMh03Vh6j1Q8chZBrwYPjkBN
87UqJqGwoUE/UziJw7ZQlwj/xX9NINOvzcCgBcT7eC4rllIT2ad8a0EpXOnbh6ln
xnA01W0O4X9ulGybUDrUY4gxc/JZi/sCBYDh40owTNtrzQuE0HMeBPWnNIqXpzfl
Vl9DfQGyctgSuUFyPzq8L8ifXOYA9g0iKS5/nr3Y6+n2bFCCViWj3VlmUFLrFzEE
8C4BXVxXh+bH/vBfBDMjlT+2TcyYL7lvfUBQaE1npt5HNGZ9w6hCECEOsl5fhEO0
UHsjT7ZyWgPE1wkwtvHpQxzEaJGUaPMobmQPMRdp7xwIT0tJUcfEDsqCI1LDtZvk
eKeBJ4fYlr19NttsyCviIvqcPYNCqssJsKB+jekSsfRbbbsdKUFydhCurUR9Iov6
vC6+Fqmtxmk51ogJoEhjPc5/Bs+2Z9tGAiuU1NCQ75CDm0JVakW6Kffo+/M/J642
tDfeyTHKtInfqYynIs6xkqn6cUBtZlW0ZvQiMTs1CGQGvPGYIlYTi4nx6cYFBN2g
GnM7OZ+d5VWvzFVr8rG33OKRBRr4gPlgONAlDD0KBbgIvDr9E5iQas1VBni8hSbL
a8KOOYpxdKIfFilGKxBeDyhnSx7hWjDqWuBSodMbYwLokodgLS+SWUIiELzFuBGN
pi88pOdN2eRmJiSwJGeALUdHXPHr6WvmLM5krKmYbsCHcMWd1YNSiecQpvkeDYyD
U0GZ6qatZfylrGAjJYhzfcfpp/mS7c4t+m270UonRZF7TgYX1RQA8X8uY9o8yI1o
TxoNY2gOIipUgHyuVGnNVcpav9zpDhvKPrjM1cYEN2XUwtTfZ5vVZOF+0okkbtGW
rL9xPo5kKtaFTwi0PImIAS8yblSrDAHZJGiVBG0wcPYMTFovzbFy5tmw/aHGmiFS
7rTMvJyUAqDIdTvrABE6/xtPcwF9lDqm37mfOj2Sz3kzCoXxJD9mYXP88GChzhMv
6owNZjAJ7Jox3BfiuroMZNUQVPTpnqE726iEZq7drz+spg95/pxN/8Egk7TBFbtb
/6Ok7r2a4TJstfe+TlMxI0rdktZRILbL9otVlzEtcsyAD9tjDaLmMZF95Xy8QTiZ
k2RTg1Ah50OKglIkDVQNAUJRcGrdDG+S4zQablmjNxpzlE9oJ62fK+fi0KeakYwh
Rs0E5BIGZL6MEbXNU3tdx6IYDTE8T7HJl3e28e3pKSQXJw51t6EP422BKDgcOkcQ
YKZeVBnPDxbQn+9GCU+8N0aEsak7Y6w7TcCHwtJlgvuKhGNSMTpB8kooKJ6UUMww
S6qdvTpAEgq47lfaZc0iB5zsUmP1mQPZi8T/6yf+BP2UaEWpIMWZUnpJ4cLAJQjo
VnvooAyGgMqrxUd26KnDfeSqRtd6qIoXVJzQNl4V6eUObrRZtHemgBCtvR5KD0GJ
dATgwpT0Jw4n+dowYpgEo61x3WvKwlpe81VFNC8lkYKfzxW/7lQwvspZPJ+NurCs
P15qFTovYo/+HXwCIpRL6MGpdXzcK0gljT3d3uT/kVJj9wMBvnEfyNYdM4Svv5EA
+/Fnc51IEdEeE5S3oroMHsbkhlQdF3z4J20foaZFDZD8LlorprFARBBwHMHGGYI3
/HSs8xyFJWrlgW4CTUBu4EARPQP4HywLrau/jQ2vu4SWKT8Rl19UUWbgBTE5MMmv
LUSfPa64b98xgDrmd/fEUnvLgNgGl2Q6QPogtDCsShsZIPUkaEPSJ7YgdKwVhse1
oLTqXN2g6TGMb/1MFDzf3255TgUg/YpnROJIt7Wjl43j9nLD5cXLlVqBlcFDXnx0
Ap5Lg8Cvmty3yOAbvR8g8ZeO29GtwB9Y/WkiR4BrHAMutPNFDzCKEEvFrOkCltg2
OlbTKS9KE8OMf44Wgxz+RlVowrPxBtuwE80beKRMOPWs3L/dS3oRm4zx/Dszb7pe
RoW2jhXQHda18s+Oz/BPYNW2tsWyrqH8uQBuEuMk8jWkhKVw3iMpg1YkM9Ot97CS
qdg6K5CG6Nf35BvUfBo9CJZrpZ7kKu9aZJ6dAJVxxMfeocSbOaARH4d19G/ddNAM
9M+ihBMvVJYNDPjqP2x79ahdP/QooFHDuqNxlhAmXdNs8vvO/9IgLOrQSoqO1tzY
CwWZf+B+J2LfPwH4YUiPnghnVhvBlUs9ooHK9il2gDvJ76ioYWRZWaaLtQST6Kng
4YW/m123sDK8REJ/WBstlk5hsSLEFpJZjZ+EwuNxYU/+EYOX05lzklsjaRHPUxz9
wcEGoGA8tQFxgon6gPtBoBZQRJnUnfntKy3VfQzFD3xlIUYejBO8O36fYfPKuFEo
WkhVVBJoKiOms2wZVgzWirLQniC0Sbmzq9iNTjH1aEFkT/o93ForRbeRFXI868IV
ZsQ7Y3/s/wVWM+TJNfv9SPM9n4U4RAs7pKvtADCsWY4gGCfpiyWF9sjECtjrz6s7
VTDJ1eArHe7ZjCdQuMyo098Z3eBW4376OFkXCfj0oGhoMKhRBN9yZm7CGDwT/Jvc
i/42SFKuuTpBFdyvgplJ7JghaRGX+UdHSuPDNPYoBmEZU0vMdweRQsBiqj0rvd/K
3j8kTogylLNuW+EWmD9Qrtl8jNgaXJxjID9TFyETaJfIkz7/ZPMzwkv7GyP6bEea
+lGS0EuehRFkoRhzheyXEda1lHHLood6+HrkClTbvzCk3IJtgNJ9Gv9lyfpuEQEx
ckcvU/YRo1iG/nrFg0g4BtyEDSIo0XeLqU82pa8DNi8o8ArvJ8k1ixOkfGkgjppY
6pGy0glu1FX6veghRHBiFNw42Xf/peMwIDqO6NtIWvWj6zk93XXO0IVgtHu31UvF
yKlQ8V/odQ60BVo3saASNynOLgvzdM7PSouUVG4gqGDJwTJmsprIlgq7xju2R8wX
PCNca3LoXeBtnApgtOKYNuOee28hWJRudane9YhZPOa6uWuWNOYi/rFLNrPWhcaX
uok6fMfYVC2WFfKH6QhpCK7dyYchd3hY9C1fecg5Wi2iUV2RZCkv4o3orGIbRI/M
VR9yJTvG6dvHNCVE6TUzOB2gUZX1Jo0+EngOcfOsL4qQluLBo7Pz8vUsA9AW+9ye
215COpj00aYvX1eZjjPZOT+97MhW5q82AlfTiRNjlJAG3/B6ii49CopDoGWlucyu
Ji8LhuMpV2EJbjLmQddfmV2ob7dFHvPYgNUqI9Xkp/MZvjr1+RcQGS+JIMyRDBzK
KhZQuou0afs4nN8JsQ1u/5dzUIF3Mc3CCJM97bAA6MB+q3xUxpNU4Tbv9Bfc5PmG
CzJyOnQqERg3JRaV398/cYea3uL4KGVeddjM0qumOpdlWtH3BFuJgPJBkD1mtGe0
+8o4PhbXlIO+GHRdTx6/EgDD9r2QZIeKnOJpLp8v/wjXo56s5jKSwSwGa860LsWA
jwxvZaZKVdFWLQVTi4fgP926+dPYjA4JmHPZEUsdTLswHLjd4R7S+bNe+wnKrx4S
uZD14X07YtwSK6L5k//gHwj/gIhdNDumBqa3KYY0amPkMyuMrhBm4bgv5lg5FgiL
fOkWCqMxsa/1MzH+0vwXPx/X0YWUOhYg5i0p97mHlzEee/xoJJtYlbWc+TwOwBEe
AI6MW2uVYsiIDzHwFyd1ALlXO5lYzmPM753VVhhVdqHtJWi+qDSydrceXWovl7m7
jSXhmQMqkmLTX5R9x+EmtBpu3lmgK1EOtotpowrXhQ89864yf7KdRmcinfh73uXw
vGSBAct2UyxiCvKMMyTPxkvLXj1xvJ6Mqxc1kwFthWjry+Jyj/WOqwAp1bYewyJt
0f+632ld9FvL+C52qPVA3LMKZ9jR+ixIvPDv+5KpPZ8eRm1Y9C2Zge5hJWRodadV
0+KxzQIVeziVipih1a8Rj9PozpkP89CKpQ1+u6brFV/o/MyMs9PuJV+T48+yDACX
YoA+UM+EeNYDJby75vbNULI8CU13SrM6Mj7/kV9l9q9Nb+Hs/btd4evBu4LZjhll
pSH/1D+8fHNuh8D6zZz2EAe4+ILr7hXOohvA2trmVDFrpnYNZrVVod05uaQ2GY3R
/WM+y+w7CjBneuJaJI911R82C5pDPnqxeBzW4FLdsadMPNahuaHoKfk5LyA6Oyo1
0dt99Ccuz9FMT8o3BUJsJK1yyjAgItCM3Q7jbAOWEDcmi+QxFzcYDk6wx3DjRf4+
frrbDq4cukOf3fypcWSJLg3bH+c/HQbD2lysoOfQW0LgJfEmWzqyVATZ2fFGL3ay
WkNlcq6zIWODGzvG8jodeLP+miPKn0XIT3WTyRzVeARk2ht+9aPNgbPRgso7wYBD
Pzh9SnD8Fw4Zs7nqNofY2BW1gCojDnfHPxkMbnW5xGVxnGw0zFZpbhet9T+asRqw
LKhZmc8B+DkNUhLWVwrsRZttrnuK89frSdwQfGdsWCNHAuRBgSL4RauI5qRMXggX
iVjGCnKhdN8866hVtPyYmDvMmqKAc2Oy+NurFh6NSaYfa8dBZixec+Jj9Tb+vZ9E
z8Eq3+vNagLTIWocIhzmPed3EDIzBZmlNTuD7hrFDbhOMKU8XOlICj+FlcpWQpXC
lW08dLYNjSHCThfV0L5WQH+ibvCU0jfgpZ9K2eM8CHNzknkzMG3WQRBg3CFMyPJ1
DXcA1xMIpCAypC3NgSGbr1PQ/9REB5aiK7203/ZCHeZDpXRq2J0I4ClM2WLsB07x
lr4Yx+REdCmyUi7fbVRGYZMH0pdzpr5fVwo6qL99JHgjHOiOt68MoLXGrjlUFiTb
viC9396UBnxlaVMhh+0e/S/D1WzfP3L3+0ZkhPSS/ZDMZBF05p8fUCHIwc+2qZW8
4WUvQ3Fv6RPEquhNGBgi1Xzy9VpZxPTmfZ3j8UDvsltwHAYv45pnEhYCrUNlRIIH
+pBrjuEMHPxD1zFgFcOAxmfHx05rrWh4W7vMOJXgCjAKzn6ajNmNmCg1vYsGgFYg
U8sAkb5FgHN5HmYvFAtS0Sii03Rcl5aMfja0IdTlSEWp+UKjureY7VjgYRVGoKjh
hV+aQKZS/yTGCbikgyTYUdSHaf5IFiZ+XnsSWO9eMh5sDkDaVbkRuYCuhbsC6RNC
LgNVJ3qJUH4BqKkr56MVjwOmQcNuoUKELXHeT13x0WjjYJCycGmiwQNFUSvWYLB9
IgU/yfQZeSeL4sZF4bHTeM2j4bzVALzIDgeb4KqsUn25Ee1q0hIgOQkstGQHRz0L
/HY77CQ7eJHaS/l0MUu40PxOwD2z3tANok6U5WwgbVkB5J3YpVV1A9JOpB3bx8Rs
af8oxqd+xoG9ob+GRks2+dWnkyfgeCGGuGmcEaTii2AA9s74PQOUkS/W1xKJ+sqU
B/MlDVZ1+o0jMVoxySibpBkJ05D2z72qvgfYiKMJgRWXdYMuyGTSo4OYbDiVTrJO
+XdP8/25pt8ju4YSbnfSlxtykB5ssI65Xa6eH8lGO8b7j5TMyhl+5Dq8kjdeOyWW
q0JHJf/TlelyFVFKEFaZJdf3OgoAm6uXe+D5k22ExaiqBWWGsAajg+7XCvfbRgS3
eXZ/j5mC9HMQCu2V+fmZhjRZIbCEctP7kLnKXFLKxzxCEqiC2mLberciUuj4kH/b
UehDi95n3vkR+VzRyzckmUMuOF+y2uItPXpH29qTSOaUm6s3nXMqbT7Qxpjhv3Bs
Oz7RxL+AP4Kdmv36MPdjduAg0eSfmdEHZ5fLCiCs2omUlcfnpkvGkrCosp6iOAys
z1KigEQyEHZ9xkSy+ZaWw3lOXecxZXWrDxnHiE1wAWepX7y0bRooA+pOjQU4u+yA
dBsfFZDx0/MySwWbtIo4FLW8ZN+Yc/WSE+bd91FV7QHp7wZVy0UxYveyLZ3ijyvr
dMV91g1dJ5RT0nRoB9chIzNqURN7oEtpWGzc9Yyr4lbiWmpykp7/z72oY1E2onZO
fmxYptd8rpEjlB+ExfuCnDhLIQnorj5x+Pu6YOqX50MOH9shXdMcaVWGiocjsosB
EGkXpu0T0P0DGjn2FvYdHw3AiEnx4zwU8R+AjkD0niRTtRd1Z5AU+/qe9GaYV9Fo
oZlLxfpAs7XNo0URyWkQtyC8m1auWJMyywqpMGMjADbAcaQA45qu5yFOv6DG5Cyu
RHyATsNDx9GNqs86l2jaAvh+7+e7O5wbZEdpkWuwn15QZ1KSJljC5WTdP2gkRrQV
OWX3fSWnPPZ/A+NG0H7iXd20peqScMtFzHbZFrLEiyJ1jh+mzQxQxiCJ+voVmflw
Wt9HVOflQMBPcxjATglHz4pzr5YbayOz+o5NOm5DDs4k8I3NOxExrsbzvqE6bi6R
uBSZCzEnuR0+Kma512dPSqXz8fKv/HrB2WcbjbjaNyDcbEOo3vK2RhJEnlMxzs04
EJs38eIMKDX5eaKIqQsIAMA3Kin/TTVPYK3HLkVsNss4IGcwEbCmtwe1PCQfIsVi
wopuUDcwxpxU3RMHDtTa1ItUm/HPwmZJ6G/F0Z6BR9+piVQS0rTFu9YHgu0igHHw
KktzwREjEMgUreaxQuhj+tQvbYcSBI+qG0ula0H4YIokvGNyDhe9PANVmw85RBVE
pm960LqaT+ynNLdB2sIn+V+cHTkaUnLO6ygg7H4mnBkkq5OnDGv+m2K9Zx9prTUK
DJxDCj+mxCDjVuLn1zhLOBPF9xDboLzV9pG8cZGfaafsExD3zAoeWiEWIS/u9BmY
JarE1NdYmpdLR0BKnI4Hb7mc88FCJhcWFlaDge6t8UW8c6wFZCTopq24I/HeyCiA
l2fpkPCrPjxJLLk/EYIrte44wqPD/ns+9nDDfCYZkEt+V2Nfm+6zcJB5uRhvtfcw
93CYeL4RLaUqKgTj2gybQtWm/QNDO3uqfdwlEqn4rYawEKNCc7tMA1GbGPXm4XSB
61l1zeCf+aSCqv0fYhhJCWcFsXhuNY0sSZ1PneCoyIdvA8TdryIVw724ZJkgqjok
RAFduhVsaBRPD3grSkZSQPBK+ls/xqdZsBKcDZ21V9tQU+I+G10xWJLlN84wOCwS
rUDg761tuy1ked+K0ZsCWW/CkdgDF8OPittE8Ju0J4JYlyjBmpG4kGcw/AjhgYQ7
3CQNP6DDIe5bAqVZnVPwuDChpx3lhXrKa8tLcmxQ4DmggJdKBnyRTifu3U3l8GBV
7ZbCKCDnCYoPrz0iJ7cZAD0nRAia2nu4XHrN0Sww5C1FpipgS1mYjhGvxn6sTTVs
OgiT7sVK5kBVtSYCiPyRVMV5f8U5SNBLyC7VVcnsovS/gIKeEiZK56bYoN5PWB7s
7YHenuR0HQWBxZsOOXDLzoQoNMt4Bz4NcTGJw8cSXk4RWBM3Ez7ZOIebfJOtw6/H
j1pFONoIpoyf3UxBKwaKpz/HGTeYsnUTI1iVBwmf7Tb93DTyTz+RKzZl8Hx+WHly
mOINVstVEUhI779A/me2cBiuMloKHdSBnZjlPAbmINNh72iXDKdRMENedpo8sM6A
Cp5ctWTrWkiFsMRD8i2uXTdeAQIrzlcyJ8H/CaaZTbNEH4eHnnG2NASK6PFIyP4Z
twZ9uPbgFzEBRPB06MOIQ6UfGNkOdcxdNxoFeTTHlfbHi1Dw6oR0bU01MX1Mw87Q
pONw+QtdELGOOwGFXEz65+ejDrtg6F3d4DcEITNzFkPbjswNy86r9H9HAiySh7vv
0Fb7ScPMZetYJRoS3Y8itRA0puFayLg01ZahnxUO4hu5o/p7k01s3QnMpDTOW0xH
HNgA2eLdrDfO1XNj7WZYo7HQc9fAFR5n6CyiYSqAdwP2u3Ti469vRnoHpE8N6Zdy
Fz+a+l2+g/FiSm4DrKCO8fSHRdLsl1p3CMD7ezEPN3xIYSIiCkXw2UjIMP1OJ6/z
+iSYGpeO2wMXIiSjphwn6P2jns7/SOY7aB4a2HpbqQdaZRO1paVNsQkCULStVFpE
+IUl2R7KRN1tB8IQsC7Ypz5exBn5JjZ0eM1r+Gozo1G160LC5o47lKMhSqrQCZUB
hAAHRxQSE8AyPXgESS8ExJu7fXT+Av5qt450t6G2vr7kPN76GKInjlE6COddnXBd
XNjg8eQIS/Hh0QYWFh0OUf/lunH86GssVh4VNPUaFJxnTR4GQD5ah9P9AKSr6CKo
BRfqog+iISMSk7cPsxcA2k7a6cV1qOTQZrW4Xh5Lf/VU2Mza5QvUaUa4gjgHRUfL
HcSQzj0CjBPBx0Cc3KOmE6N61CthhgNhDuAF++TTXyhKb6S53+NN5yBRRTr0bsI2
/LLFBn6wlUq+dyKSSojTIzaKj2H1+8wttPG4iH0ArNdHe4wTJqPZ4TMSMF6UIZXa
BiFbvCY/aSEC5EUUm0rAIruDYi5IOWMak7DdSMBg1z3Nkie+cO4vZJcp+tHxLGbg
0wZQkXVwj2JfKUmRpifl2UW29ShaeUp+2OSdP9Dk2Gvz15cs8RrfkoKnKgLL08FA
JOEdJtHd7RGgKMVl6AUg2P5Ye8QzvCpT4EDklSIUuJURXIHpHzCmCnk2fuo7fZLJ
pXcBS9jUl+JM8t/Cz6G7fek33/7kdi1Aoy2UXWr9z9MTaI6Ms6BsnAZvLPQrLoBb
HajSVGr9nlnWAocN8b1VE/bh1sfo282HOKDxxHRFZlXsn46QvFASc6gW+uu2yZdP
6Vvv6LAqLv8SpUkeOEdhn1nN8LUFEmVNpAdAFZ1izibbXreXfssoc2KAbeMl16tn
jdVz/BXT0hgB6ikik3IpdLD68q1WZLCP9ORfXamuaPyEIcQ1q1tskxzFzClnpBOP
fkjN2kmshHywReRrqxz/g+olAnLrSdbfT/UDlrWJ93YxSFfr32ys2nE4hhKLrQNW
GaWO2wU0VaQ86x32yES+5Af2zO3dk/ob5YihuEKwEdh87rKe17dQ5K80uTFTb9Yd
m45V3iGi5JbcU0arUw/FXEBPH8hRV863kf35UqU5pjl6xuXl7oxtDmq5K4seaWwi
KUEmBeh2cCh+s/2DYmajWll6D3CeQqsDuvxa4LdfqYvCL82jEXfxD+1bmHv1D2kg
aEFw0JlK/+UMUGS2zJj2RjVp/Sj79vKDcVj7aTEZOz+NaRO3z8FsRbrG70viGsw9
Mu7AwPlDya6kroVlB5lM5yGbYC/rhalNNsYWt5CltzOeMCkA4Sx3ZCuVMFm6Pn3/
FUW/VXM86xPT89SMF8qF3zuh2Dt98TmuesGM0C1v4GNZ+5JEKOxEH5dX9gzXkybM
K/ND76hTwkTfzIOHljpWwPuwOejRIUPiUgUbqJKjS2rJQWnCwliIlvLP+iWN4qKN
bx9C8KVK93oD8fGDqK4cOVidUmHE5D4iBVwq/chB0Olox1IpH+ts/df2uNqbnn7X
urMJh3L15cSZ9nH49ZBHdh2jTZU5gUDqZhvi+OXIvz04x6Hl9D9k8xQPHvGqm5/+
MKeKWJXMRdGhH+y3XBdnTat0tM4TiJyBLXw0VV51r9XlH1QNv+TBHwEJ6uOP8aUv
hZXteu/qVPAe2cw+Dth6Peh+/oYKC/uHr87ilpZ+LmgPiUSyW5U1yLPHaoBxzeEP
aEk+rJNHs7KDwOOGyIpo1VNlIfQI/ACwIlCnyfV2ik8wOPKfmY3WnFjqmGMRSAK8
UihbQky6A1ZO4MrA8/T9Z0S6qqFK4QbQ26mGOHF8hzGiclyQsfP//3w3EF91Kg87
Vh6ZVkKlZDKTp8mtn2oG3wm8UbE45qtzuVbT4ndz4sQnr3YCk77+nTDCWhRs7ifj
vws7u/FgZYisI2v7YDw5DDVvj2WGz5AfEn8UKh6n40RLw6F3fUY2NOJ1gOR3k93F
h0n08mVceiF1hHoKFF9nCJLk8ZDQoFSeBpvrvJEyfIL/7xVhhhTLTQKxKK6Nf8/X
9aaTXVWNZ5sDmc0xLf/1E+AJ0473mTg6Xn0RJWS2anYhoRD+GqxxmD6KrjQz5Kk5
dV/X5y/4G+fDsqZYbF3zTd0/oVnS51HNz9vGEaYCfmh+wGdzd1jmV5BKBcym0BNP
EpYtwxjvf3e07+lnyIEny9xljCaWms81AwSbix3LO1Ar/ObS1pEYdgcn3gUL2y4I
Uow/UtQVKd5bwJiKtR/REjxzy7VMF9RRwBnHvwQ9NMX11JXKm9d5J40tsj7Af/PE
3HE1Gwm9GDKQZ63RTmGCECQkbXU3MYoyHOWHtA2Ca7VOCn3DT0af24rSqyyxuZj/
UN51by8a5hJCWqSfZnAe7kP7BAOL5m95x3hIe4Eg0G0gYaB2BWxp3TB5fsuzBdTi
w3jz4oKEcN3KlQ8t+GaFwMieIhfN6G3mwq0kp3HCGf8+mwTuo7DwSCJZqjHH6F57
FrgQ4h4ZSalgIWnKpg3/Q8SU2RHqVdZ/ewowzS9E3BflhJVghtZn5bTgjQdiZwjD
PmVNXkfKNeZZ+LPxD8wgR176fDN2eQ0Ql/GIQaRfom6p5GRqlYGKhKfswkOmCf7Q
NycFjnp8qPZi0Yz8AKRQip9oWolEFywnylly8jwNMFEUMH2gLl8fiYpuFIVHDvvT
fQ6xQIZMpXVDysvLTpHdKFN1ZffUcBrksiLe33M4+JEiTGgsis9IzYiiblY5dsll
JB5VE6tx/9L0AUeQwvZpoS2aZjJFMTN+7qJblXk9A0eMOT+9an+mjRjUYI2d0OQC
BCVkJdSB2IvSIqEvbpoTTC3mfl9cx3ogm5wK50OI4ybIP92q+WvKeM05+S0FDaAC
PU3ftHLpv/eIFzij55PDNdbCv+26/79bEiwU/BBinuaceBu95Yasxq47Dy11AyCs
/UCAmrdLxJD/QwNviv61EZb0eZR/e30XMOD9mJV/m9JIlvcidHkelOldrFBFcn1q
5sjwxQYbm7qJTRMXwx8wT6GoBJKFKS67HxNIanUZ0vaCtpRTalHYYBgwQRu6eLgr
wfFhwqzw9YD7Ig0SLm4kqZD+ETAvYuia/d/myLKE47F+fbXLeYNapCROQm+CqJM+
9YVuxCsMHB4uyHmmPEt4+h+oLvexKQkiUBPx18vlP8Mn8K6ax3MtpA4kmzW2mUFq
Xu7WMwAdexEtP8bJLOAX1OZJ17JndgqMi+YtC9BBWx+Sx3Y/JO1FLwUOImZ6IQU+
I21WTMGYrNFUhPoB3t0o+J/jAjPLsDUN9WlzAAxX4u3aJoRpwdiCCGf16kIfqIAh
fTPJ7U6x1uNodsdU1Pj14n9TN3o0hAygNSrvFKBxTfL22fFjh/3CWTYu+gQC2q9+
tFwDYhulJcvFnguuIUarr8WKLrIADJYxviIaAn96ZWh/XwXXpnk2s9s8NrcvxY5S
3iBWgzOwVxbNUqRh49qv3t70SRlcqiDm8CBcLAT7VK9I6rmT8nmmpRN/K2gtzwd8
I0YQyneM2ukwQ2+4iIpviJZ6P85sEZrXkgrivME+ZukHgRXdqHzkCtGab59Lq7+L
tNeilRb1683AjMhucH3jPd7dmAxkcZIM4PqFZBrbCGkNQCeThMCI5n+chkDE9Ar/
ca52ImjqLE7o7Yp3hp3KSTQ3ov+VnjjvXZZYCC7hOu0XkAL8W38CBcA1paix+TLO
6UoqlXUTFn1iRs0Z7P++eX9hMP27iQzFA6DOtcX0LUhS/BOfGuDhN00ZcByEfngg
B+XRgUZIT4875GFgv6s9J4FfctmvixxGr6CIHG0f/f1dm5q1wernMeYea62nYHTI
AXLWhRNc3d0Z/VqEK9lu65b+KNkDh7HHMBKTp/pqEtbLPQyEB+mFRdkIAiHQVXoE
m5Mkedc+Fde48wMm/GWwot+ILHwMKFjPlsbPQc3JkXaEJ/hTRgwPaN50DIso+AKo
++RrLnLbxSV3M67D8rOVx9n9Yj0c4zd6HjFm23jHOr5rTDZe76q/Z5guC4ezGjze
vZInZYMmH0xDjQ9jSnjA6/mtbqO6BMbEIVSCsT8Onq/JMzkUDLDaA2HiNQPLcdVa
V0aiQitGewJYFq2E7lxz5QdBwQUkCuQ5UkTrjjmilRSVl3T/X8AjjTaZEAUQGnDa
ZgC1JkaNVkj1qEMseU916zuYjETPHJDfTP1VNkTJFW66gvPIzHySvovSPQuZM6z/
ze8LFAbR7H0Z7AB37Gpo2g8GxsMgMJ9q0/yvyDcO2Xv72N0tzxZoe61Lr9lEB2Jm
blBpEK2tTRSkmoqiRzJb5cx/jCF4KCgXkmk0GzbS5v9Dy+RlQDlH8NkRoMAGe7my
koDdfmlkwHPghIoqG0vT0fjn4PvGLnNti3Ub7QCDhi8PQ0BYfRX/6tGTZ/qVx2Up
nXlPJt7MnGwhaetErePltbLadb8m+vmf05ehZhZSsNPmV0h/AQmTlDyRIM2I4NkU
Bo0o496ObDZ+HKi9rCb+y2IvU9tjlIW3jDereMMOc8N8fvzxIYO99Rs62gkHVfhs
ZwB1Ji9EBnpgW71EKFvCIeE/PYiHodUdK1es/cTVRNlziKPR4dbQpjiZEVmNHM3m
ueNyuLqDgX7TVbRF8ONke+PTRg9FzSSdkyTmePGmsIAv8SsNB+LpSSC/FnphrAKF
fbYJNWa6l/3I/+c1CjVHZW5aIjFnNe1t/nl2dbt8F6XTNizkSuS3rehpyqmVnpQz
kNPW+vSDU84wgNw00vE2xPbKhhjl9PTfcuvA5++Hsr4jwLMQN8ClC6lZ01d2F+cw
vnRIS1Kbi/O7BWeZNXepRWTItJ7U5hjE+I9vkGddknL44YJNcTnL3E0QKbySw3Ig
CpvAOcRQDOP3xgZsLXBeEUBDSdLWOrn+A7ak7G6Zq5thDieMdDv7Y/AxYGHdaU/e
NFSOijmxmzNKlqHurRvZmisJ8jL8bHSeNdsJQJuxJz9jrMchRS2kgOJ0D4ljtCPi
tT/TbbkPAauvt0iN08SoHxVsdFY6CDFCab9WvJ+jztZJ+45gqXs9dJRia99Mtl0y
5z+SuictiVoC4VQCV6aADMaWKL9tricJwzG15qfTSLy/kIRkC7YzHUywza1bxmhI
NAzuB2NoseE/aW3+FUZ1EQ+rfwzEIDqNNPDqwFdfvu9civAgaEx++81Qbi/E75zg
8q6KADniPnIBGHDSp7x2pQfrnAuxZlyp1E1VbBMm1yv5+9IT2jArZrKGAFtQD+9n
o2VXWNe6JyM/4h1ZgxTuGSy2QizvwwUKvkEJB1vhf5qUJJ52P2339aPpCblOI1Ak
zGlA/l9BnNANXS9iKgcUdfC1Tdpu/LcxCjK6m/jodafn0TQ2lPByF7HMgzQaFDud
sP0YO2Ok+89KqHlwMAg153jzyl338LDhESEcjz1fFzQDsXof6o8XYIgQ4Upy5I5R
0/fqyrnDU0sr/cCOWw8NszxVhrKmiV1C73Y9BqYFfIas62+pVAqpZ4p4CnigQF1b
JKJruC8XzFub3AUweWheRzqzOlqjU3RxuHiAj7RYsN/KMRqWzz+LjCnqbSuAH5Ek
Hwk8vENYxcBoGhFUni1h5omcvA1fRHilo3wCSvqQSOq7JS+jhDcIvKRa+V5wmzwN
v0ETWSrwy5uAF1GX7hynU5AQVl9yEvi4/IX6lN6WsId0+v9sCoUm61o6VGNUaD/x
0N0SIpxJiFikHKGcLPmn7kWO3RpwTZLoafjDa23a+EiuLACuUwBn3Gd5FPAo2q8G
cEzofxqW0ClkcPyQshmZTL+EAj9gQfC+gWD7g3vsK9TDRkWCu54orP6A786QQN9y
ySfwn8MDqwjWyXADMl+O2HglBE5hoyyrDKA1+5MfMhk3TFEOcXBgydg0Lw6xZ/1M
YBRT+ErFSQpQZnmlb88AcaQ/hAsfxtSEuTB9iJw++Udh21EZIfgoVDcWeUA69Yya
BQkK3cXGdObo6bFDbc7OgVnemjzPLFcz2dLIdwIOXsrcwMW7IMKsZF1J6haeqsDj
/idaFAbxcW9d+O6x8uaJLbCcrN2QFAibxlfaPd6R7xjRLvKKh6o31FEkes+/Umfw
SBynyi/MtikLNWxaWlM84ZofA71fCgTWnVEBFExJGvkcYDFI5Be9hOtOkpzkOTdx
5w0/kojXbeotXS3/MH4GSYmHqBs7oxueL/SWTFRv1wZBSFvEvjEpR3myjhiGHFxu
Dcs85HWVnZskmEPAzD8MZHBbmgOkJ3oGIMfPpZw5KK+s7d5cld/ql+P60TwLAXl1
SlVT18N9AMW1KtIFS9ZNCkR9vB1osjXyPcsTvbQ1HIDd0d8wNCKNq14cSyAXTsTE
EgzJsq0tmhDATskHqGgzHuY4+gQl1AddyspNHIhBPSRBEWAuiNge1MvM2hHZoNdg
h0nAFc73X7oAUMuCvTAmtDeWwS7fr93R/1KM6t2lkRuhufBFxmnG3v5zOYwHmIm3
XMAgdebhlZvtnJshntWglQ+BlvrgfvqjqPw2b9BKGoTadDgHMQrIIBiddkvC29mX
S+KcZUzss5ZHA49vCpY+9pJiHW8D/7vRdqMtF5u3uG3795tYAtIl0cJVUOu3lk3g
c8EKGKJg25Bhm9jTTDE8bIfePWch+WpVms6NIVXQUzeGXL5hC2Y2E5uO9i+x2Bz6
KX0feOQTwujC8GVDLXPDG7kcWq8vkpQxFKLIhPKYdP1i7uP3LA78KYugOFj2nHbf
jhafC8BZyACA9uWSBiYM1O9SHCUNck4j+/wZmbD62OF2qtGP5W2fBqDLvOngVeo2
2LzjfpCcshQQS3OAT0IdRQRy0SNO8MbPPTBx+0DcuvYmO7xEvZxvW9ZkbnKImoCa
5vd5h+RkfjOy4wla9CXp8Yhqn3roLYUAQslPrV5XKmt+cSwgT4PO493A6H4vRuO0
/eilLCb8Y7fzzjb2EC5pgn/9IEMsmNRCqO/OBxpw02pv54lkeFpV5OjRLVjw20Ty
M1bR2Zq/KAR44KM1mYGaWwUpmuG/4h3iz/w7xGSD6dAdB5mNc87ZNx0iC6vdWvUY
1vW8cNvTYZrbiBZko4Qt2GgoiAbodOU2OOeKJ7OvkU39yugYr2ru6LcOcmBCvjx9
WJU5wHghFDbjiiV+dCLbMnml7TECaQLxd1QlmJ1nvcgzS8u60nyVQvQAMD1tyt7Y
uqZukgNiApGONAGDTAIVi3xlPOOSHzz6jRbVADgC+5jZ5Y61vW+VFosEZ3FottQJ
fR82dqMqDstp/K3Eklh2A1xNQ/80hB5tyzxzRACBuR9ihlZns5fdu0w8zNyAu1bT
tqBr8f+P+i3k1BgqP1z1XrhbmA53NHN0V5Lx0LDHtwMInvpT+k44p8BDK2g2bl9c
v0HNdbQ23NRfMykGiObCdw9UweYFurKxjtoNOVEl+InQxFBZxbIq0RE53FzAG+fs
c8veavug0ho2lXnqyu5ev1YFKvjqbpQOR3cx8kDqMdj+n1Q7UJrpywDbITjo4RYL
eySxGjlrqt/REBtfTVexznMRwL554zVs8QLSQ5xIBUXnbuIkqIrviKy+2RM/xugG
hd5H8SK5Vb1LrqSp7HdnmgFH8IT+O8WETvYDy/I3Mo8sHWh2jv4SrQ/02cEqSS35
YQomWV6RPFdeQC62veoCJ9+kIOsBmf3Bewvd8JckqV0PImp/n8Iu0w8gf/om2CAz
MbBWbAbGurLuFrxtx1CD6wXi/c1brpEAXQTFv6LV5HMDdfgl6ywVVm1NGHBD8h97
ld/ZWuXOTSDoE50ILPKaQsFzZP9qloVyGdM5+lq2uNX3vMLVswWAdlOqjqS7aoKq
8eThmUNacE8piCNUGELloPK9l9lkfbJ8VdnOFBn+jc+PMJxwT4qBCFA5eRp8K1oK
3wJwlXU3teQM26vkAhDGE/usGM+De9k7qOiGLqSEu8xpZDEWFFWUsCZyv1sb8f8k
QM9OtEX3P+FperAjYWhBJnjxcz1NBjrPRQ2FbBMwTjx/TEyzg68/pAGICOgxinLy
Vym5AO+wnt6ftv0CZkSjBHOGD0QBTb+WnFbuXWTvL8NHF3bWtDxpqk05PNNVh88P
G+oezB4rRaCtrXJ6+ufI2Ee6hgEwC2PwBaU5KDSDlzobZmbljp0nlMmhQ0vqAo59
/q/BFWaZSlI2HmHdnboAYuXf4UAeHr93USk+ML0LE1E37V4SkvhcPrqQBUCRW+rC
qIIFcHjVT3sX7/lsMbsUZUAmNQGopnNsfRX6e63MYOJDakgjnqRZinWPvsI081RC
3r/Gi6brFmpupBo50TEmiRh5zLTFMIpJpGg//OilOxMhiqLQknzSUy2pU3CuZZLT
1Zj3xzGnHMtyd16wVi2hgPlyRnUjCLuZZwMsrVWILwLRKeD1CEYUGIM7MuQKnxfQ
m0cQn4eaW4THxVbvO2BKY4JyyA+8F79dAQX3xyvhgfRu7AZSni7XBKjNAJ/uSTXz
PFsB7xnEy2wLW0pDpU/TpRuFp80Iq06sBTazBr+Uc/tSYmtqzIjPBdEYbejq7JVE
0lO07xSkLQHR68I1XCZyZ8hslFYv5STHNOCUv/xlaJe+e5Q9JLLQLf3J7vd7DkdT
h6LjFHUEUKtkPcPdDGyFsqCsmsEFx9ZFnc0gUdVtdBaeeluF9T123IRnYCm/FbmB
hU8azCyZNCW4cjGThsc/sHGQihgevrmaRgFFHZLzUzOVkaoJ0oS52WAnw4Ooa/ge
UNU0ZgmxByqSojeXJFvVjp1F22Ax8Iy+OrWOWEIbI07/0LDhFiE++e4GR/iGCJ5j
H7pvpShH70OMo2OIh0s/Et2DqPFnDp/rWZn3KjYPs6hvzS+fGbm6J3ETF+rOMU59
AEBfP3/bZJGKE3Lv8mCsDYS5JIOEiJjqKQtRKjoJg99wjvAdglSB7LXWoy6mURb5
rdV0KnWgrZBGxUEKR9rImcETNcCzRVwC5R2MHg4qnQMQZXEly2F5hcXEGCJV7/1o
/AX1O6Zb+eriUDd9WMh0rl3MNH89JcLNJ6tqx6g5eHaEZfg8uJsUdIrHzpdw57sM
nrzRQ+Ufcd6atOP0pFw/BSV1w17WfD78I4RPgXB5maZldj0iX0bp4oikp2roHklu
r1Y1URCuzb37Spz1gS5XgPFC4MpGoVF95jCZpoDRz8QCCpNhBv1lIgfcD51ZXg/r
XK6bCGhZ2fWGc4jkCOct16qvGEuBw22AGHYMUEBm9Omagq+cAF8CQ87MzBoJ770a
/MYZM0ONbKucjngIE664Th847B8y9cMQNGMyrVcgnPyTijYB2KMblsswgr3IUsEz
/D5lg7cJBIC8+Uu8gOMo323NFmVsYboieUEfpnjWK6Df0Jf30pArgQl+jEtUMAZh
5TMQ4NYjmYb9klXU7/z1VE9bHHCLQ+3j1LFrw+vZMVVn24y2P9/E2YKjgJkygT7K
5CiRBZegeKhuGDQJWbKrakznD3uWbk+4ArdxkH25sbddn+wXNMTV1490mw+3hxmr
pL46WnIZwmyCs+rD6MbbPyUYYvD9KAkJJMv0p3ga3OouhraR2L1i0HcEeLph9avW
FEnOPXpjy11m0V+ve5M0gfzPxFWbO0F9oaP0xMdj/RmL7snbogHVkwWMjPJyS+5a
qwkrMcDky8YYYu6Tll3V1t6CqK2hYaODLtzLAfvRgp2QYODsb8ou+VHO7Q0DQICq
yfOOOGcSkdi4haEqK4d8KY65ThJRMPBzd9cKOKSK3uCQM4kwtJEJAH6WnPSei9+n
69zKODMlEbHQez3hzh6Wh3Ga4gEWpVoU4T19al+1yIombr80BL5U3Us735+tGoPJ
taZrIjANEr/vnUvjcCH1m834txGRqoNXiV6DICywULvE0p5JDXOy+acMXkQu7hBh
dHVLkUlF3alFFPQGzAVpt2nd2yTyu28Dk8m80LuTMKyIZd++8RZL4pTA1dp5h4YA
MlAGdo/7B5nFIgPN3ronInQ5kDj/FvpAXFJaOCsuhvleT/MlekSHMjEXwXcmxZnW
F17+OEy7K5Wz7xd4rGdJmhIVNQDzwrrXzav30oeOSVs1k7yST1XZ7q88Egvz0is0
h/YAeaVUhJBZrfCZvCWsaaSYbvvl5uhJmnaMWdA5P3endxSa9AfVJqykgTaAhCu1
qzPka4Tc/5TMZxQRxsGLHSihrUrr/eRI3subAGkjrrWStX7RIg73OfGZsmbN+u6T
e9gz/dZsv0iE1i7DQ87E7YorFCX2LvBvdF9Q0vaaylOXys8jKQjXkRhgX6QKx4Dk
+3lAdyR+tewENWaK5YRCt05cGpnfLPz6rfhGuNiFygnzpa4wLEa2oGxcpcQWR8fC
bVbCYGyP9h8U0kFY/+tyuVzWAgiiGBA0EgezsE1uQ+/q+96Gus4jpszIF3IAh0GR
MoNfzbww+0itYrAeDVDaa+ZXZYJ7e6db+WyhjZ/r0VjgmkZShQRn1FGF36TCcZEu
SNXRdSCFHimzPDLRuMw65GrKgKOyKqJllNPhSBhwNtG3+ImV9LHqfsenbI7RvgJs
ydSkZK8OLMVzlmD3RLQkYo2pDEuCyd9D/N3JobhDPxySO9JRC3pVhl4FUkFzEM84
05UtkePwKXM2ZeeRW6cgjtvU+pSSJGSqaUVHJhq7B5QXMd1Vha/liRfTT8aOj+uw
P6y7AQ/KZsoHXhGgVBSrK30iACiqPFALuIS/yS2YZAb8bJKxysrF8OO69+5l4u9R
Jujd1MJ2VcnxmBTRB00Oilr2yTLsrKwHAKX5QoSjDzRadMSamreIYTCgr/4g8EpA
IjOdDSI3pD+bABADvM2KInWH7D1r86Nc0Dr8Oz8A1k4oOXzpybM8pHgYNpbRU9+P
ORfRYbKOUaA8Nztg51RhNZdByvOePc90ZvDiszx6SGMOdl5JTzOyrxZL25L0inPI
XqVToCrfjF/S+guVD+B77SzXX9pI9hX9EmB/iqKd1BGH5R1OmexJlomyxd9usyOr
4vRcxnZiydFQzF9c9MQkP4vIpxuj0q3LJb8eYbDQMPuzfn24kelKEevhp6dS6eN8
b16KJfweQtVns1o/XL+9O2eDzBphdSbaDUlBKn40/KEgiNqxdYoPgAvN0usb9RU5
7Kv+q/BB1se1ESMQiutojbL213nYR/v9hjnn8VcXcsCOIgA+iKdTw79LjLfKFhlT
pEJ+3aGj+366OWu6YyTH+AXe7QunnRYRj36RiRaaMMVeFdArjGh4Ddgt4NF4Ug+L
TWTsOdOvd3sHmGR8YteYqdhM/7B2e9M45I9O2OrrBq1PDziJr/9TQuOlFzWjNTVz
c2z/A353LG88x2lyA1/Jt381u40Jox/+ZYPXc2fxNNZzl+gx1c35X1aqOKX1/Hww
a5shNqnwDYO7mcCepHx9iK8jKp/lBfMHCSbXkMpYroytu8VwQsx6ArCH/z2miLIA
TCYxRjis3lVDtMe4y2J5IZ1r+ZsJ+IC0n2SHVYYimryeuSH9wm/7HYE6rgqLz3fU
Q7QNbEGsZMkVepQEgF+HaUjNKtkjE1UmAFpRRDodL0N9saHlBD5U7H88z6f3eqHg
Q0z1N62hD1GiOtk/pJW3q7U1j0L0qDk5TZgMflLDEpYTiSm9mDB8Bkkic3aVg7fZ
d8FTSVfTDIEHuMQ+xbQjtnZ4dgpxoiZIwNNLeqM8sIivrAh4ydukvoyhTfgo/j4+
btAZh9FvDr7PLlxNs0jVhw9nGIUGXCbFfRSgxOhW4b5RWT6hKXImamRpPSiOwB8z
PTdT0u2NHLcNbmxWUCWVqTsysK/lyEDAXnEdFH+qEC2naLiZtIOO5cEK521loHwI
NbxY3tav1FU/TpCWS6rfNOFl93u7KUoUsXflVfm6Gyw/Pj1UH1YM07Ye2uyhyoCJ
XKykhJ7C/JupJd+Y4LCR6GVFYUbAy4lNS50/BqO4rUQdeQDLb+xobus4wcvewsjq
I21vGR5nEDa9R3Kbv2RQljDPXTKSF5IPggfxaLJRPAaXUVCUgEcD9cg+UveoJxbv
XPxozrHv7a2MVaQc0kxDeIHzVep4JOtR+z4hg1X/ffl6G+2UOq4Xl5v0MT0gMlxo
lp7TD1VPMBU8mHZpZFCCldwlweDHrsFpMItBIeHJwOaaBfqx8VWuNNu3adgdaFEP
tMHBGfj90ZmlkmNvJPMBPsXedb75d5TJeyVnKqNXiGEX6PXpcJ17VHaU5NOtVXem
QduNmiK2q+iKkpL8K3MG/ps+t8f+CjN0txe0qHbV0LOF1rTcmvMmqUztABxtDLYh
+I3fiTu/cQ1RWvzK8utBrHMYYPmj1O2/gyfNkXrUyXCk/f4ftrqKBhSeqb8omu8V
eMCI2W3VhfSoxXh23MKNuQdHkiiIBlpSCllPRTztePUBHEwk75giacMPVR5R2c8D
HPlLEp6dIbGgKvoLfuS5R/UEC0TBAj6Apl/s3T+3PHlcCB1ipPywGKlBmAMbheHT
8n6vETropwMPTgk92uQU2oAGuarRz/kTrAaHZzCo2EB/tGxH16Pl55jojbmUXsd4
aPw45487Yzm1Jj0y9+dhJhdhomgQo/7yNYAW9jPZSrwMrqw5GXdkt/44e5l0zKj7
UEoM4RexqABLTONUNHOBir8EMDZRgeLmeJcCgnZ628P5QGVZpYM+BVrO99dI3b1B
GoQfTLdMwtLzKpTk22hjsNKylwG3n7wCiZ0+NVElVqNJDOo4FmQ0DMJ6B5hW8c7i
nKsRO3B2I8MvCqJQesn9fO7Ov4dFrrz0Ixh5joqwjDSxy6I3ws2Ft/atwfLTeKZ8
xI/jU9cBeTEgXLgBK+NzTzKV/fFY+qdxT+Ln/DelX5oP9XUPCDhaHCTKNX87N8tk
JAS/HYM/9kUj8P8BD+Y9g6+9t3V/ClSfPUOgrOOk+iCg1lqhy2k25FPQAfJiFbX3
D/g3zuAxQReqcNA97oWQGS+F2O84ALd7VvwF7TeqggTlb3O/nyMm6WYnvPL6lS4h
ZXWQTl4DalVH43Ao4EQunBSEiQxGns7iB6km8fizqfXdc1EemglEvyMorYwS7EY5
Nm1Na45HtbPcVX0B5B8ze86x9RovpyjjVpWyw7oEbphkmxXASII+eviig5JF8hfs
nXoVXCVCi/KpyY9H0NT1Fyae/cOIN9QoB/asASnblpVEnO6HJ48tHtxCTHz0ZBrg
iKbUNHY4gP28Olk7xuOm05YHZFih6zpR2bAyHuR4nEOIG+ueWcsSKTyuo6Yj43g3
0sJBaSb4IBiEoq8A2AlgjHUS+DEcQzh3ml6pzEFZl3ZqCjobksF1czXr621pzbP2
8F3xTcKq7yxSHR0HaAADPUxE5Cxfk6WjwJvl1yK/D9ZxkzCSI6fNjn6GnuYrR7Ni
OleE0M8CHV8T5EBkqLxKmqUdf29q20/GQXCt+vNNkbKAE7tp+uMZZUdd85nUh0pG
9bUMPKG7ok6eejq0IzjxVTorUJfn58qBvbamSusmBmfTjnsUDqRgCXhlBjNBhceo
2A8LLi3QLfwb+dU73aLkBXQrQy60fLWkxhFOumCLG5e0CVdhppFsIQMa42Y4VdUe
UuGL52BmwYWh0c8c6FJ3He0TyyQAD8TK3W/Cbz4ksdYXfQCsM5p17EaF17oB4hrb
G8ks8CUZc9YTTt6F5WExphh1xSIJz2w5C3zyIOoDQcetrFxpbShMWHt7U1NdrVMe
G7m6+ZKxSXUzCx7ZP+8nBlwOHLDn9yRb3AdOQ7NlyrVMKKIZdbRcrB+3WLMO41hv
2ZE4quNwK0wCENpDVUhn+sT6/coZeOLd92DufxzaAoYaHGPYg8j1mPjgjyuupqJw
D+ZZUhlyzEEIKKHJYhw4Pu6onruKIBSbPJNWaUVZGrII8uPN6K9W73SemGKcmGyv
hVK1JeKIeLhiUoO7TOZ6X8yW1Gt5aF/R+XwJpRLCBKJ55x0Jt4ogeSVn025L1MHi
90MEvrVMga/zfp2XzkIoZWYLLBBLAwHm8ECL8bqhfivHtm15XXZ3693/Ie9K6KcR
tn2YCiLI1wzLoGGhtOzZZIaIBVeq34AtA9tQJ7Sk2nXLeOwUvBXNjgK6UH02B9H9
lkc3iF0ysBCRrahX72hWKSREs8YJ3FIpKdnFPL6OSvEkWR+IYNLJkWCo+uDSHNho
qHv+3n4yLelvqhORkZkYoHQ0QQnNs//8yIZlw+Sn0ePIOzbDS3+0YIMsgABnJFjd
7ZdtGq7Vj5Lr1gV9C8ytfZEgyTEfhD5dA8CoY3+LYopzbQT2MCaDW/9QRNX/HodK
Rr0nDe6ugw8jwHGFF3jSlw0pAA4AF20ncNONfA8EFs4tBCRMXY4xDkmH4oXMRSEx
VyC1+7C6/bhSGl3GS6vIwF54W80Rqwkmxvb6v+iBqvjAHk0Z4W1GVNVBVnB51NJ5
yXVzAvP+eY1Qfu+bm7jWeJdb1RgSfqhwSB0uOGqXsl/vusuFFY4CaZbDtDKjCzkh
EzFDHl72LuUGOHN3a/DEXN/LqI9zU3VTeVIomRs3gelZFuIJwZ/ocXCK/D3MGAYd
AVmrWQF/e/rPUQEJn6mRd8lcgcebuVuxe+9qwn7Nz9c3+eMn7RAaeTUHzL1Pa+8S
wibahDCHsiO8PwkpHMjQyjqzFrsfAQloTsqZZjPMCkvF1dGI4bpFGrWVpoArO11F
aXOrgwJqjcs83Ff0AEZ9T0XZP+7bkaFGoqzgA0+LC7YGQ92wiEQYKgq9SNzzEGxj
7ckAkcIh1M/sEpUXD3y39S+p/9DI8pJ55xMcP6m0roq836+b0Aaecs5mxXFMrhuD
aUWdMdiCQ055/E2GVxGOxbSDKkUsVUQg4SbmnKeQaCblOPrwTGNKpn3wFYQE0JMm
/IBqfNYISsjxymM21mOc5SQuYbQbcwAVrsypXm5sHsogqInRROZCMbZ3DJ2QRnsx
lhGs15tC/ipJQ9Wrto8WN2hJ+TLx1TvhcXf+cbev4QGG7/WZzNTFqcVr0S1Al1Ut
nGPMr66g9miGXIVROI75JdpudjL389DkVVGxT8BXVOSCqyUIH9B1I0+rsEwETioM
cwiCGxiXKj9eMgkW5NYormgASpPz9w2iII/K8e9VkeiJaK5AcqJWTBGW4yhgyQUf
b8BLzZDqRhJK3uNEhQ6EP9C/qYb7sGhysW7b8TJe3VnoXYFdAQ+ijVPI42ExyzKF
4Pys4WPXsQCBXV4ymyj+AqzGEqVq91OkvdsrWKj5p5gGjiEKQ/XqkiNEQJtR9B37
6WMhBzOOR5elbs+IxJZPDQPVyp/8bXe8VYgpoAQYFnbOBevrBkr3HhbqEhOrLA0u
VIMFYK9GheQVVyApdwmU5K3uswi0ulfrEGVFIqLsfsBGidYsEg8wzFjyqeVWydF4
Si4M6uvJ/bgvXaKWSw61yNz3tc0A9buHyTH4AaPBACSx85N9SBSXl5/0Kue7/gNK
QTMlBRGWJCd6RFvMiJTem1qhscBQu2u5LeshmxZ71GMMLBdLuTmpDq0UO1D7VInj
abfm5OthOM+AoDd7ibINux/fgk1ZgloZvuMbpGxaK84X2x4TKJV/S+Sc4bBJxF3j
e1e23N9qbkHS3nEhFqdTYBcYxkO9AP4G8FiYtswCKEc4tmGXb0kacvF9Y4F59y50
jtFrW781J3QCjtzDOZErlhGrUy8qyjADLsl3ssQ05nPFdYKxUZ+saYinUfV8z0xO
iTSV4x5TSG03yV62UBfJ3GQZXgQ+om0AZFGPT/lYBXgnKcsgsFMJ/kSHvpTdayWJ
iY5PSbpdi1LelZKEeLhkRTpPkxzpQyENX8mdUzTPPy6gHP08m+Uoa7B1588WbUyR
PKvj6MZDduO4QtRfccSxzLeqT33ZanQl2zYTTy7Vjy6jsuVoMIxV7UFY71TYg4VU
ZDMNFqJrOTrZtNANgf710bYeHPhFhvqVf2vl+nhkVbZWLXHDNnl2OTrVCt4fpvDM
/ZPKj6FDDlKC4IDyuphzf9LeTJXtUB/Uw+eI5kxgXFxBDtrE1g+4qamkjbIsw/sF
EnKH4tf5nVCKJaoJT7JYXnjf/geuzU+h3z0vqCkP+bnHqdLVpLU6f4ScvC2rBvIB
bbWf7CW8ukD+pse6+cyJG7Ev62rJAes09ioothaOdLGsOk5ItPzvd2c0zBbmefeW
U/02aW4IVdwTmsqMP551gXlzLGdZzn5UdsKU4AiwRUlQwSw3uw6QViHwmV8npgNZ
zF9NX1+fbvb+X56VwL3Fg2VA0qWOVB3Q0v/DhLHxxppF3diKxfVGBu0owrco4MuI
g5GremGt8VyuJGa1z6XYwZpryrVjozkTMdsruXFS6N3kk0clf/U6kfAyJl9zrIwu
6KbMkWrOzHMAE99x8i0mB0Urcn72tH7kUp3lQlGqD6pX258isAOfm8BUw8L1SoT8
u3rTMP9RZiX0QoDzal/hAeT1IFsUIOgv4YJQ6bNUsGCMiNW9lrkZgTNq7uUpEDb8
5nj2NYbjPP2hKiqPOqciIl+RljVQyD9hUDmFUZR9OzsABAt6x6CNw8UgfnnGswC4
pYfVba0P7MQx19k5ycH8AWuOYSkzqAUXJ9XdCtDwn21WB8indwMVZ8Hof7am1h3R
kkRtxw331Ws4dAlb87uqnKRiKyk3NnuY/Hkr9rVrrF1QTICqvnpzUtUtrZcXcbbX
F/mlkkf8FX9XAhSRbBZvH7RFWWOIn5/HDM5i45fXc3mK7ZOh5/xGYsu2J5vQMK4/
PSRVixcAzs5Zh8SyYxWmoBVtZG8bBmBsHZFo4akZ5kJF1fUvgY4Q0+17laCHHhwh
cY4WsiDGZn9hvuvIwDRnyzolg/YfTjFwRYKYibZZsDjddGP8wtQyqJ+uA5exXAIp
i4Bj+S2cmDLscL+JyW7CHLPwcgD46xNymo6o3ucunDfaXteyQ93YiA7uOZCp9yfM
PUBtL8A2jYMpSwTj3vZ2+D/4TtQ/NahlwYehQO4nc1SU9jOYjLgRRtfrS388DYhI
i/ohM7zP0NV19hJkWB+w+l0SnWBR71fP3gFOgXbo5XQAl0AO/Skl7q1zl+/3sBMR
pkG2nLL8YKw6aRG08vQUhrvH9FLFNoaffBrcj/Xaz5PEygrWxWz7AzC8JOo/hAto
xeiXqQy9hHFB9QIKKvozcmWv6OD9RTI4KsaNdYAtXor6fncndh03ix+mn4YIhBJt
3dWoRHqv/l6McHfVBPwDDRAdIOV4VeS/4PYtJviFQg4KGXM3sZUqT6ZIIz2YkI7P
JBTlRyEZSqD1lZNyCLH2Qb/x28WBK0qVoPFvLa9Zi3vdUiy6uFCMoQAx09ut1d60
l/yntx3Mh4GobUtB55FygDcPlhqH/Z4xbsetqfPEvGgNIOkNZZyuXok/mHe2OsFw
vks/wyIyL/OAJq/wC8mzo2Svb7fhZt8/Tj3frO7Cjj6FrbuzcE2WoSh0jUE3w46p
eMRyekwuRRuy9q4SpKanB16yb+UjOlksjnOJSHmaMnt8ZeC2NjYl0ao+oBrR0uvj
u0ultAGUOnhK6TAmb4J2DlLvT5hpelqvORKeLNAHArP4LDw9EjTt5wRUJKqvM7i7
XpN5v4PP8Ly2FlAW3Ce6dZakL+08qpoRRbP+WhlH2tIF7syAg7KS7ij63tFjSuPl
XP+vIL6DUZtPsgnuqYj3CcDjuBsMuWTo9pPXGagcE1FvOf2he0ftTavcl47NCO6D
dJqbf6hpeFveby2t5f4/bN4dStgH5h9zHLzRNo0quwgG9ULwYdg3zALKQYyfNhbh
x7wrJXEDMR+tnvw54b0gI90gK1dDgNMNdfCZ5AKTdmAGxBA1jBYVwVIt13H6YSMC
khy+QahMZSbMpm89jYgtzoKSocLHrWsXMvQ/qLG70yChaTx+HP0kg9EaPedhimi7
K7va8YbIi2rzbdOnOJTWMnqlfKli3h9Sj0shVqnn8Yypn7hD4s1U4zRyN7MaT7mG
hn2RtKL/0srOXv2sthSsesoTlQyKy5EC9RTP6VoIeFfQBDmU+jIChrySXcT1Rn2e
VsnzbwsHJg55TPwkHhum3PHIIqtuLyj0x+pZn1JKkWmH2sC/7fYFuMzS1jsRAJWp
P16rjLwS2ByNSSNxVfOijYY8FbXx/8G5j7lmLR4WhsYrtl9ffzaVsREY/PJUBZN1
+0jHQjj9xNcQyya2QfcxTNU4PWh9reSnLYOyCaWgPtHLwwsRE+lWrPA6oM7+RxGP
rCj1gWG+ypLWrNjgecVE/MDYtzbqCGI8SONBET66E3wqkBWsoDDFEKn+BsVGQT33
4ft96piTDNrNI3GxRk6pbnPJ8mVl1eypxv8ncv8fldMJ0zq2mxlP0Zy0J1m5YBJh
nzrAsHvyf+Meoep8vLNaQ8pBKsUekcBrt8zPw6yK+mmlU5fe5VD5Vg0UipIzAHw6
krbygiiXWZ6VxoNnKzGlDHbSrZ+d7V9+3bF9AhhEnTGxhAXZa49r+BUM/5BMKo1A
TQKcWQtuLZtta+5xwJxR8Q1eSlr1j9qojNRWmiZmexUKvn647S2DijjapXn8Mx13
bG8PFCTfjajy7XAPHueBsw4HRBq5mm5PHbAfCFJ5Ic4+RgdxNnlrxRRaENi/Z5Oq
uMaypwHjXt8MCZs78BU1RuM0BVU5Xbvy4/9XNyXjGiJh8Xu+ndJNI+ESjPnNSFOq
QTJdDVWXDi8nVuqiOiPCIIf6QrB6wKZovejhy/zTfVZw5ILCvwRm4x7CS/XTXxTX
SXXs3YKJG9wefi+rh9hG9jTR6as0D19kNH3k1jPguoks76ZMwoMIgfC9T4OJ6mus
+Vj1FUQSdU/Nf6vFhOBPt5jdoWky6aSb9zkvHZ+WmJlMYrTm9M/mqjh/e5EGvGrc
/4FOGco1GHS/ukca2y+pN53/b4T+KiB1JnZEHPoSCGo+HDj5xKqZKOJW8GCNMark
kTjDp5Mtd6qZ1tFgZy7CUy48T5dJRDQx8IM9a02uWEcPuHq+/4l5jz/YwxrQZ+wv
PdNBQwBjO1JfxAPvdFnugCcXvg59l/Ubp7A5Zuf+m65btm/XOEDBjpl/UgmrBz5Q
yNIXRpgYoTRuONgDZEoE+Rvmuy9OeRFs9nLmJuw818jVxid8s4dOcIAqArXrKaWZ
Z47xYq3FN/Z9V1SLXpshUw2RsEpukSSX1t2EVZH+N2XY6N9H6zXZleviEff7M4dh
c56I+nmx/Yd7f/vDxxlZYWB4dEJbuabwZ3YoDbh/yooyQ6I+wpnLYJLcpZDkE4yT
LOGKoRATAQsIX9qt0lHMTc2V/EPnS3g6xA/4/v6G6BcxjSh2aOHy69vuKjmpmZ7W
m40CWjphTB49YUDx3Pss28i7YAFnOokEW5o8s4jwigX4wCcgonxWxRvdFxuKFTfy
vA8MeBEhGLjnGQbAeTjcUEaWHsWANIf9ZuR9q9SVhbX8PniKbBcgm6357QzBn85j
PJudPgF03ru/5rCqylIHdi3PNEsj2KN/Zh6lxfcBKnnrXkrzFsl9ri4gfF6KpfVs
EcKVrybtWznEXkhQSHYiM6YlvUlVYRo+qsXexQfuWhoIviK5wMPyZpTiKWUuwqDj
ycu9IR4/JXcrKu3PV82WYV/J3mPrpFLRnM9CVKSt6eV8cCU9867ON7yo97PTNbVT
OZUaXbc06mDHHltQmO6UiMRVqODoZO6sbfuQOHKC0IDbQC2Y2D58+7eNtojjatJO
+5UREv7WzQ2Vfee/PPgz1yjRbUZWZgF70rj1v//f7L7vj4ZSU7QNgz9dQq55acnG
n4o7PtJDn+w8QvzJ7rjTCHf4zAvFMnA20jABae2KM1Xa/d5aBi3XRpaPWMBzpfSH
vVpNF5a3Im5twqfrW2NMSh1LdWTleyrUMcaMU6LNhOfbGIJT5iXHGrtCksNL8cEt
AwByTx4M9fZavcRlKdUWp3Zk/EYzhtqPsB0tMYfMkoQjQN+7f34tGKTYSKay0kUm
g1BZ2Mv/8qcyhSETIqgsMc+smb4bEtsfSFOcuLvtnVl7DZtN4wUybMwPQhJ6Zt9V
ixXaEDAPtu6fuWzmkDJock0gAmIhTJiyTD33W5QcnTaHsFsEj3w7z5UpZ/Rglmif
5cCVt3a3I5r/28Pils5arf51Rf987epYWOUg+JiJYCE0IzukgRvef5aljy73OAoB
vVwUEmeW46VEOVTR5N4dhbqM7p/ChTvfBm+CBFmkA/qnLwGqrFoowlhEpieoczvx
njgxE5jSgDz8l2wx3kssu4oTdC4cByiyUANlf9imHHyPB96NWal1BW8cfQ4y7T5t
AP+Pk9Xhg0ndq9AzKRpE1oW/O48e4oV1OdY0O0s7vwQnb/b3IfVP27S7ThrgtFKJ
VAuc/IfsWRc5goldpoqAtOIHq4jhpt3rDM/2BmJsTLC99ZujCUrZAcxZe7/1AOje
29doPtQ24MERjdqp2JtmOagrypbnaveRUuNCmLL38KpuZYAcy+z7/v7OOOdUK68y
cddAwzuoUANny/CVdMWg/Q9kMJ/JbCz4zGp7eqxdb60q7HveYCuq0nPFERr/y2p1
it2ISd57Rw5NniWgIo0GxM7Uv9u/63NM5KHI4ikZ+dVZOv5qbS2R1E8/9mPQV3DD
VMmF8qB5hkGSC4acOKR7nX2drYdXKQ1ZHUdq4iH1w5f6svUIw20zT3WnQqW2Df8j
4au9Dz56swObcfgWhuokFxh/m+X7iUeuVkhGBEOhoiGB+NsVweTIYYpE9MpA2vru
RYnA4xR4mz5056U8YEpS5asj1gO/sVu3u40c3JYBPWNu4Bz875hFsoD4Fn0/IWRZ
BK0sgMkR6VKvafHMcvVXcNehbpUcwsEOJc0qGjlL9tjla2bCLp1JaEJftVYLEGtR
0uH0C/SujSh3ZGs49ydkwBYV9TBaITZsVWgEaYkAo/yXzOHXh6kP/jKEiXKi1xlQ
2NH15frgtU7rVmAaDz0GoSEE5BksjkVqhdOpMYac/vFLT/bYBjaKfBLiDzckXhUI
RJ/SZ4gmrmWccN+Ou+bazN/dgr6GMpgjp4bfhtnlSzG7AqSB1aCVxSCLYi7DtJgB
5UBU6zVJs1bAulULq4868KAio3fETuFQc4qTy7azJ2fBpTwwtjr/NZISWGCOqWZ/
GeXc/zDcvArMeiHuw3O9et/wkwRXHEqlATTHl5XxsrJj0ss8amER5mGwCJSmPSAw
pVa1j0l5P4MQmA5mPrKyWN81Ax2Av1nR0PF2fBgNwe/ZlRXJ+y0KmBo2sE0UwOgh
INd6ktcOIb5AwlpS9UmvmyMQ8hvStCXojBV9blJfUbD/+aj8CzH5QHFGdyowkRK7
F7VcCLeRlHRnuWEpNNDlNF+reGxyuwLMM+Akhi9X8fIWjeZpEw4dMNJldH+hIaGR
Gjrlo5+VTLHc7+SdAEezyTMteY/I5v66Srow5MC87MX4FnUvT9LM6oRvnlDgymYa
9+aTIHmbBD4wbXXpvxjaS+oM2nPuPByxdIcKeQ36aIlFCcy76bfITUn6MY4Dht7J
00WNhKdp4DUC+qi/WD+C4RZg+sTw8OTACjuXbP7gJvLNUbQ19VvkHXDyYRg3fyV7
vzKuMkT0pNHfUCQTh88bipb4N7EB+URgGssydj0C2yyTG1aMAPYYngWU+exIcdvN
9J18QZ4/LD5WCPSZgn1sOlD8kwN5aYoZyxGREmURmfEaUci07iwKUCbjCKuE6yrj
1lccc0FVqea2Ghk8BIDU0RIQfvkD8D9OhB6lKNIVdXdnSussL8OGGWAJ1CL1Czz4
CLQdTRBLZfR7Ac+Vfi9bR/D6Eg56FlOq/581zKXauJeyO8kbId7CxoJ+a/44tPAL
7CejQDsBoCWk/agYHnq05eWwcwIBzgd7NXHIrtt8ZfWe9TIskEfK10VAmJfTNNbe
zi6o/Bho84Ql1AthE2F4+XaAj5qyhWhFPSZ1Xm1O8PZthfeqYjs26fv8mrXBZtdQ
0D7RfJpkezfYxdbhd2QiP2aYfVJf8edXjE8RaFpfsSOkug2dgF2jsPEQHKXOyMWR
JcNj1g5cdN8BOzCh4/L/iQttiPRr7Bw6t3socn9P5H5hPkhpNb2NtV3n3uq6IGcy
Ib+tarIDoOfCjGUCXfi4Zs4QfHYyyl34W2WZpMiTG/RZg2nvwnpM6Xcq+YjqbtbF
qZX3DIZbNyui27MjkhAbz9uRB9eAn4P+qMpyBwtNDFsMnce1PtMZdz3rPMdNw4VX
287vf9bHlexsTI8kMbYLGPI3ZmwY4loY2/ZFuk7ow1oJDrPxicytK6u1MKFCz/10
1oF4vTiXjKWPm4xgHT13FgSHLPh0JLrsiifboGmWJB/xK4LO8EdEnTnVOX6WNrLd
5j3ETiEyDpQFnMr3XtbdSAt/KzvnZxPTL4z5ddGCnvJ/oGYxx11LgQWShMb4USZo
meRp4U0kCcMTdl53OZ8Yzyj7RuCpoj9FKBkwsEJsr319hGCqXawXCu0ag0xz9R4u
zctTZobSimu9E5HnUSnVQikMU8skbHbta3aSXu6H+Z+8/eZ7YL5VOG4eRqwxuaft
0im1b3zLMcWddpFYcplEX/FTvVBSalBsA0gTzZGo/OW5kJLucSiI03cxwMC6e5Cv
xI1tE5bw/L+UZiKrfIVdQ84Z+VxHuplfXBZ8VALqbtZyuOkk8zjNOuZy3nRPpPZq
WdQYhc9kOjNQop0SMub7TOrQK30Va1XVFUo+rM4h6NknktNMkR8iwYUiFe0IOflb
F6j5ThY7vnSm1XnTkMxdF9TZZSqxKts2wszLf7Bj8qmskDBRBHgZKpeCyjboaB1k
UVlODeubCeR8o71ue4tgCSJ+csFsavv7mNhI7TYCFCQwK/K58d/f6qgKJV6H6EMV
hG1cGRHhWVMGcwyr+MDIdOZJuc0Mb6yNu3XxCf7QVSh3VTTkci2xw+jAys6kFEDP
tvDNoaCU6K0LnNVGDI2G7HgoGsjVxm0C+vdq0eqlCwfO1BMm1GN0v+JhFD+sNaVJ
A3Xu/6UWh/8EwYs59tiyOOHBEHWJiSuU7k30zjXonrWuKkzglU8iAng/8nUYwuge
r3wlWVDuU5Zr2UvO8LocvEEwP/1f0QBYKu2/2txmIfI2QKmbubZxGntHlBbtgpXq
bJYsY6Kr2uTuMIMrT7gll4hVIa66MtIK3smNPI0P7PDCfyh4i9l3RAKSbdpifHeI
Rn2MKv3ziruiK6OzTYxNOLh2Xf6tbB8225ReJJ4q04d0aRJjJ9SjtRdvTrLVqOTd
sZ8U0aN/+/1qBPe5vitDE9axtp8NHjMBgKLR5Y91x+8lBUsFSpgs1vmfFw+OOqit
s8sy3lv13N3byhLDNAFK/lS70+YKijiGOSMlt8aIcfg9m5/U9R4Mrr6iZvlhgDfF
vmaUs8F6TzlP76xAwQKh1l0zYfBVQC68neHyi1D3iH9C94zepTmu2BZ7fdiy4+4c
UjYuLPObBUidA8qGLOnwimTbp9vzxNp0hohcofKKjeSL15u/43CD7k8xCGODKmX0
WXk0AIf1ZcKTHXuL0yh4eRWutRzIlFu1HM2NnMWigJFKdKCf9hqpymyzRF+Sb1FD
0rvVp6/ZfbM23kks0gxyajTwbOPo45m6g7PE3w37Q90XQbGzHV9A6a6CtdjOutZ4
wq/wjRmq4qd1qsGhPLwOlfWAr16bcovAj+7w/qyxUfUSvBC8fN0PuOr4NnrVo32k
F5ASB2BDEXcz9FiXKIv4R47E3N1gbNQBAjKf1HCxG1z3dikJ0brLiQxLH7RbcayL
+W9I9CWkoL3bRy9aRaWNyXkzuXN2Cngv//XP3+bbcXKxnxVL0ENJLhgk1lgPsp13
2iDGymuT/7wYjJyX1PvuWvQDiosDj6sjEJx/Vb6yeR9eHQADo1bt/RCPDOChBp14
szjMr0SqpowRPYTK2l8PtHlPa9sYxHJjeAs4pRyFa1Ht8LZ+liPC3NaePqpo3uFw
6uCNrm9IXUBMnZefH5+e/hTgc1rgnmBHQ/gRtmD9lP6LnWMty3/UeZ+eLP4mCdR4
qkmPBZu2u0/wFGgLTrZqW8RhAtLaV+TFfRbmYv9uCKDNiQvROVj6dz0OwBmSefby
dRESGjn670nAANC8C/JSm9TDvsRdkliLoMRxS88MOjg6QZ+CXfF7xBj+FspZ7+6s
dUEvui9sQ0PpcusQIstHYVIkxguMmOn+2tY3ev7q6evGgo+f0FgWO5MGgWNIFb3m
dVFjtISUnIH3U4+6NbXhKiNktgtudVZxZxO65OZJyDs2TmH5AJiJrFAVn2YoXdjC
PGGd/3lFHbqiHkrwjM/w+iO8IPmGB0BDTJ5Y0cV0rRkIOoKWoYHvyEXgwKuu3kO1
gHbIRNJngXYnQfqGWDS68Rz3qaUOMAF22wB2cOOd/HwfIJ63YLnYqbKHDtmEZ72l
S5wG/j5YM+7vShwuh9l2HrGiMvyRp6zfG6I7GQgwf9YgF0oyFtRh56+6+oKVcZaT
nmmkkFNm2+Aj6zPk1SeXm91ug53BjorP87sq8Xyaz8WRrYT8NbeGbw80duYQCTSy
5YatHM6N9e6yTMLfqHBAelnVdUZTvcU0ppUzA8hHoP4kDacrxL0YqQvIGoyFn+vE
BZ2dnJXoocLRRdXsFDn67w3xz3zm8t7rzfO8h/yBL7uP5g5O+9KUo0vA31ecSIfI
u8epP2ugfowWup3i679Nr/dXrnpvme3Iar+otw57S07U9BjLlKmBBa6x5p8rcOHN
x6qW3OSslwtb337W0NiMNHu2szRXESAT3HTEJqGv/86IRFYjuTeQB6vmGcRK3Z+n
lyapV+xJajVevqUVkADyZmQMvTQXbCR4gFlg/6Rbaw7MoZ/Y7qTUjcW2h/7N2ZRt
yLzAPYn46EhAGc8NdJ2rdwltYRpqIr3nZZapt2Yv24tL8bxS+4T1EgtNrEfQzl92
OOle5nzwbaSswtRMIMKrazqNosVaFFtGVo0Xc7fI+rfV77kxbUFGohIJvfwUSKV1
eMppayf7a89i/RAmaU88iiMIa0pN8J/g9fUMTfXSvlVBi0WhR04IbMAgomcGjPLI
2f2oTbygQ9f6Jazr7Avs/Kjh1q7k5Taz+W2U2Ln5PziH46101J3WrR+JYrhF5gPq
G+rwnEh93rRApeTxfW5lqYIuXoebMLaS80ENh2lTrK+qD2EjFbQ4p0Ssr7fYEbQD
Eq3zQtqTdbrjA//3MPxgcQ1bTr7ckdJQgt6JG4RENCuTPOz42+46jE4wvGfd/DD+
I98pl1IIFxW9mdGVTYqZp/8XRzV9hh/XMK/sKIk08VMNpiF8PfloyyyKledwUPLo
eUFVWTdDMpytpawM0vF85lSqI6LwyDSbYyiHwpqpAB5Pyu81UWk8w4tiVmKq305Y
1ROPAqnctKaCDRNtML8HlUuNXANEtBOKgw6BjnzpsIVX5tq4E4ocwnXmfGiQDmmd
3qOmhSQb7MFUkb8oqro3hxpjS+q8avFrSyNhpCQFjJGpJPaS8YihKPhrcTPe6Sg4
UiVZ+YK/d+2NqJnUqhHA0DSKtPy0uKXF5giynSy1C6bSrm5ZeM4txDkBSKq30zVH
JP9sBEBngHztILlmcZtPNCZ5fSw67PzB1BMcDuki+J591MbdTslNq1jab7GvbMf/
JAKnwG49sFdOuqtiYlQR/Nl6Oi/Z/Ox2vwr6itQBWddeRhd6+LzAe/gG33Eijh5Q
3L2Pndd9Cz179BSJjQFQEmwNNUiQMi4LUHv/d5HoNJMPAdKk1h6frryV5rVL6YVN
AcDCNHKACxNjtjFtPbjPw8U9Lsn+13JaHC+Jbupo4YyTeG9hEQHJmH/xC5MxBcGw
haWkQ8Jn1Yi6NsYvN214cgQRlzK9AUwW9VtbRRyDiRxpEb0W7pF0v51PBN0pXg7z
n1+5Z8R4Lz1b2e+/6ugFlJN/w4nnooa+RNG5Zz/13cyhhpAeW89xrI5NvLFxSbz6
hGEm0arQlSGa0pNuwyFTPGIrwOsWTJr9p3aYccTsnUVO0h/6n1ykuZpK1ZulRhhF
BcAc6QYdQX78ift9YM1ySjf3BV/9b+mdYI2gbEGjaEYwo+dsz3qKE/xDPqIYEBHN
qjGZm6iYd5qdowTMGAX52xgCLXoZCDBDrl72HEqnTFjzYHtATAIYsL9+4wwcJcMs
o7XAkL/RVe7wUKkE5/TFVALZ91BLL6WNHB+KaJO6OMRkQC48Vpt4W/oDmv1CAXds
MjshTdPDrXdy1An6a/giS2FrkiO4ErPui3duZ+8Yc3jTIg5CGn1/w4mZ3mFk3kA3
keLLna7ujbroFgGjDn17x1UUaLSPySGd08bEQs4aF7wNTgCq56HMx2IfyL+1JM0T
wlpQImPl3+QwUVOUEwzaEkNd6zWGdOpMbrzfwmUu3iDrg8qc4mI+qIhmND8/7AHx
CkyuDRgi6ouReWe/fkxquDYYOZtY2RWAPqFLGyQQAxN50J/8730XdPcIX/zH+b7w
e7zgeIQTjLM/4P5G3J2YRMzZEHerRWEpZVDSiIyY1vfUcFbag6HctOgAXuD3F6sQ
AscON5RRqRZnyzYuSwRv94LKhtylxN9bIaHyLIujKAIsvSBgMiVcDTBhftD7rze+
ZVe+qKX78zhvQHLYVmpDznHjU1ItNo0C0Md4Nkfm+Bu/jgrKbKwPMWviuSEUkCAk
V5KBwBhgJ5QGq1SXPBRhmsZtUVhPNT01u1gcQQDuZxoM0qiXs+X7/OFVvEbIg4Mz
OpUj/pwfra/dGnIkcwwnFLvynMC9eqOw22lH8y0B5Sof5mFwabg5k+AhaYtMakRY
yqryBcd3gjxnZphUzkxPMegkHreLL7g5KCH7asmff9CzeMcLB9Wgfq4axnt7pIMC
u2OwfwKQS4lgCGpsJSpipFygNAYv4CsgzXGCk4A34AW0WP01YpmWuQe8jgOwfDTx
nVQovDnTX6bC/jmJTxE9IoFwC8u6AX8rZ2VOFUXbWDq40zk4TBzz5tpzFG3ORdpA
WrypNFy0jtP6y3aAA17ejYMWWJbFg2jAzfmpfFnMMFMyH0nI8cNFXIOi6sWiC/pN
HnaUKfjudQvve3nLmDabn1EZWwvKpjFtFgPZOHjkjgdsOSn9bcYThN7s8jhv42ge
/9cOKKNtwvP4nfdDCoqqNFopSuK7z89Lu0oWLhTt6sZUtfXSQsaHMyh/tIDK5THL
6e8bGGhziFWXNpiVbxY125VuBqNXPxdfY8XjAlYY0X2ISer9u7f6M66Xqaj3fQjl
yVBgGHZX/v1SZFXlhb9MFW74fsQhz6tKhFzj21Ieeew9EDN2G8QKfjMjux1kws/0
MgHBOfObA4iwU/jtFcNbZTdIVl5x01UsNtE5y/z/2oADvXvIhITZfYJifxwyscBz
U76VU0PIxrsNONSJ6SripPKxqqSj/MWOgAtuMUHby9TDrr7GH1x3HRpKDF/k/shK
UDIB7KegX7q1bRdAnUY2TXS5Y/fN6iNsdFOTKhbPUZuv0Ys3RaDteV4yj1hLCpr7
7lRkzwqHjZGGbme3OwATSoxgwWO/S31CeOp8Vzz74KkR04QVeKV/W2FP+XuaaTJU
sS7L4cURa5rUrq7KuB5rFiz1nngAHxK88238WErVELEnglxWZk2EYjP8/hfje7mF
+mDLsZAdzQHjymux3OoksD+qOXZswlwxMByAWMBBnjoT3bh57koWppLMHqrN0XBh
yZhcYdVOR1Q7Z9iz+r+hTlsVTyVg2OvR+CzY2i2wMUb24XXxlqxvKBwq7lPhoONC
g2bBUqKgclTw1VFwDQIOMLWnYKF4MdzFxJKpQOXxB92cllB8yhOrSnCNFkTxIDd4
8HPZY10sEsc1NfHglOLiM7Uc9jcovjkroHrvYGDvFiIF+A7re4Q3gw88x5gCN6Oo
qB/kmW6Py1nvUkVr96csmEE2vyGXGbgRIYGXhYRWG1UTIIFI+AKLUpIqOIuwCk5U
kEqyYimhEAAEbv2grBHmRTPbYrtKCTbH0uRhdP6qZf9pzpvPbHnv+iCXZt0MUiHa
UjOw4TLCNiVC6wwBuh20dsvAR9+p+4+yid30doOtc6GNO1/+0Alf0E/oj3N9CqP3
HySWfh/PSXmvn0o3OqGJIgDPjZrs83NDnApTE3f/nFPh/LZZVSa8wO6iUNZAdfOA
+MDAWCluFMa5zPMWzGOhEUrtUYca+st6iiWUp7E/LMF0AIiYi+3ed5emYROaYAbV
Oysx5wKOJFfuA71Gsgw5nkDcqE77eKBJD1YncJf4rHHjWf0Hl1c17lulhY6YPgYC
8iC26BKlJip0qvOeZX8qWWVsPmHM59MnBNJMHJZiRTjTKAEIax6GTgJi2f1FD3e7
b4TYNweRmeOBwp7XAWFf3Q8Fyq3fRPru1xBOnww//zWp1SW5ukHMPnCDWOvzg417
ttlkKzK9bXHzFoYrqd/83RrwszJ92SRQTtoyQYC7KGa/J8/WSslN6z71WFApRGw7
vzHhk3/VYgrC6vdqncEtai+0ZqEwA4ve44kDNEo8azELI8B5rg1U4UXA4BAFXez9
IX6IVw63Pxdj+csunkYHnELYaICqvTOEiZBc+NG0wCzxSvSBgdH8x8mEHA6F4PzA
CAOdwxmFCi4BW/XMi60a07fz9+KC2ASu2leJ/LdDz1NVq2gQ2F8GOz0Z+Qi8tL+2
Iw9X8IQxSlAr/a7SHlTgMiyqSezouFn3r8qp/4rkuZAwzrzv+EUmLnTNpfMw5JUH
PxptiUPGMZFo2l9r21v7+c6Zo+w1MXa02CY4CVZii5OCxEE0SAKnDyDuOOuA8j1m
LfPiVv3MnwvEEHxu4CUuMF3xknogFV7fveKtPlHIjy2P7+8CVf+hAbmhuFc0W3AN
3ApYQetrFuVx+eUIQv9V0aQHeN5SDMjKRcqiT+BJVZ7dgLg+0WkXL9hUF0FvG9ag
hp/Xv+XPE+j25hOrLqOlgHvEsP1dtoALw8yFN92McLngvpubg423MJbQB8T70y7H
5tMGEVNnYLuTwjlfhyuAhfBCZXLM5mAkUreqlOYJd1Nek4wy8HO61rvh9PpnRd5J
R7YIXD43BRkxgtAxnOiy2oI5N1XM2zppeurmNfhLEolhL33krGLGsU1npuyBhK3E
tmxa7pZFroe3Hd1FDUsleJ9xalklZ14WdoXYF/qR29uKPXzrKjbCXSs6qloxem6/
+lxhu8pifAVUTNFKnJ4jtDwUsHobQwZoGmuGF0mn9g8Ob/Smle8B6KN0g1ex0bE/
jYw45ABIdL3eeQ49ZVRbvTYyMgf5K6mjO8qhUyWJ75zk4VhEH7HABtMb4Ruyu5S9
sQwi50ozNh8R+PANYNWBCpfsSaNinQIlG/i8ehsmxInpyrqjxsfEXXhAoDAydUlk
PWuJRlY7zgQT+lwe2s0LnA18ryldIVwwLll5ZpKqCtEkA+RWMKPj+rRBayfLezjY
AgzgznWiBMKWJCDI3zfOVXOf4bVNNTUmCXu2YFtB2VXRmPpsy/9hFza0Nnk534Lw
UbMTxB3s/YNTrwwOlf51YW9THQUgCNqbM3MpYQY9hBTEcBm5MJyh4ySGQcj+Vt9r
bzzL7/ZmEd3g3melE0Q8BCVY82H9YsgjYy8KfXic28waWLNT+wqrtbDs1M3SF80k
dC045JE2PLDExVumgiKPhmAAY11/eQU/bL2g8wwy4c5eUzSzGep/84xaGWqPJW00
arz4cCdaz59DI3tDBiTNWUZgrMgHQsOJZvvN0oHA2qiblrwymhjgu7HoCYtDfv+b
tHalmqLVHWsiSe1QPHP4V2MAk+iwcSJ8/BD+vyMJaSLG27dC9SsNbC/7hX8BzIti
9sIbM6jfvMlxqcywvvRdoZwW4raIRPUSXOV8Ql4XmzA3K1PfZxVwKpbS/ZWZXYR/
9drIZEvN6c32O+m88Tx3v/0ylABUHR3NKr2hGOgJagF9II1bOHR/FOgmGbovgbFY
vdGhWJqsgW9ZfcRp98Xc3ghVYKzsWVHeD9dNzEP0x01KCYbC/V9ILbMS4hH5tDaF
PGsKqBhny57zzXe5IlOtuAAbJqAB1Hp68d295hQDt6SmGrWGUwFlXMJXnZq57dzx
DSWWY2AV4Ih0SgErc1nRcpVFUAQm0aV+oI4LsreaRGy2IZmpnEqI4DrmqT9PMdst
Vcy/ZWWeND2vg0fZcnIgaGaUzP2PqQHXEOgPdDu9UPV7n/k0B9RUFP0Mp7UZQ05L
piJa6aH835VZdd+7Z1GmG1DpLk+pMY2uL/dNqNMiEZI9fyuNsvNFQmvu7l8MLR6y
pcSESblcUTj9OK1PWO1xqh7GQ8oAB7s/fbmubp4/VM3xseOt2qctnyuyiUZJjpqQ
aEVHMgpw1xGVGUjLrrdfiCFY326DLYKrin3XzN4yukg4scYYcLQsgmDg0rUxyS5L
by49TduBa4Las1KIip4EehIehH8D9G3LzaV4vlF3Ks2IZ8bjT1+Ldb5TQywWndkV
LfYV41AXmMyB6mK/JkYXoig9va2mxm7dW+jiecYM+8Xi+eFShoHA2btwQJaX2Ey1
d0QSO3h4BXmgNE7RWEJccJEFCK2zUJBDmXj/u5CzwKkNEvfR25x3A1Yx8Wg2nINw
+lB3oNWu2LUvn2n+ig2jyiODWW2ve+V3HokO5CFbSpPm+CPKPConIcWetIgdSbrX
ZqMg90if+McKHkHVoLf7VGpKlzkwaVFH1Vz6jqrWsK0h4onU4znlSXgoG1guH34F
UZMj8R/8iSN0nTdXZjoO/1okTe7vtxHFmRDF/b88Mw0fs97b81RcO6XHdDJdQbfc
t3zWtzt7KjGXzx8Zh4Ay9VGYAyrq0cXL2KdMOIroJTgggPXaeo/lPk78/Pot+ZGt
bbKoPqeMPKDxcp0AO8Ji1b3sbYz/bYLJT87YFVE2bUkI+IcuNkleiwahNKeBZ4XM
8Z0r0Q1ikh+XImu0QW7qUlkVipaNF8x9lztcUh0H4W0dRRCvEjnvehKtc1dFsnh/
umxlwG+MYGFaTGn2F3qfinhM06iSzVT2w5m62akG6z27OnySZx5rgCodoqf0Bppi
GNQlvN6T6N/kSybUV+ShZUy6dmiaKAtzOchGwprJjYNA3873KkeN2RWJ12jxDBK4
LHDDxJja68mDa/4BwYir4zmdJqI5pNpBL6TpgqxMtRjQXSelS5VTAkzt2wvDrft2
DCvUH0biuBjx5yD1MMc4i/xqAHKlWYorEQCvmpMoYJx8VOK2MZWoDGeUam3K7Hvj
LCHESOEMipVF6S2BPCIAMZckyE+ArO4XtcDEijYJWG1qJZpQnDXmn/BCbiCPHErx
LBomDQ0LNbRs8N56Bk0sdme4Yc6Qpr2WIfy8db7zott2nYh1xCYDmiMmj3WjKE4P
3MxzRho8WysSTBGviS6ck0m8O27amCh6KBmiJUrcRq64szbHMnN/9Uraa6vnH9Zz
MmHKDa9w7OapOJxorLjDkZDAFV566HjLHZ2odcRcvJ7AwtZiors50dxVF2dfnKzA
Npo1Op14WYYypPBzIza8X8SGfv2g1OLkZj3R5UXLlV6H38vh9+UytbIQiWwKwFnn
1hpm944GrBBwfAh0V3+q41+ZYgY4aQyVm1v32EDKyqJVNi8RDGpF26JcZciKfIbw
VUPzOA1HE69/xY1fJu3c0b2B/rhzqZlY6luRGCeMNaz7LjwsUVZQ8XOc9rfuPqsr
GBEJt37cuGZGO4VOT7/F78ksmLHrAPeUOs/p7SeNI1RY+0M1pAHaY9A2LAeQWBVF
J10Haiky+6Acl72qPx1BUEOmAqGSIA/XsNs3KmfigG8M2/ssNZO7FeTB3GnTeBFV
JAh2KQ8vY3UtnsbZOGwCuPNq8CoJcmDAAwBSCvpb+DW8YtN7g0eb+dWrmONjxGxz
PERf0r+GMwF6B7rRnsEUeOSv3jmY9+KVytUNn0dCMQdxjAhI/8kJpYIblT6w2NeW
TxZL3bw7OKGmicnrp/mjzDt73Axcld3B3NcgcDVqJ0Wl6ZvdwXcQ40l0WEX/porn
Y8CIJRZ8yBJgIww3nXaQ3ilmp3gf9aXWldkachhAXsXEakywqwZ/GhMpy19y+Nkd
DoMyUh0cg72MVs9zu02YvpKHhBEfxlc08gm8HCZz5SkCzJFH0AbZYextY/uKZd2+
sVt/x9c9QzcHTIyAujdCS5fRVYcsg5jP2uKUjYtdVS3/V45KoKrtSkqzmbAYAB/F
4QunhrwDKByl1Rx0lEroKQLhh5AjuHXJYPGCvRgEs7uwt2yhsvz6cOqLTxroYX37
y3+U5OXA5k5FeUP2R8IgU5B0rqqnhcDFQC+ThIrku7IxXqEwaaz9cNhws/Ve+c1t
ww2hxZZG8si0IehynTOrPFxkOiAe4LjPbEEQMVBBHGLFd5L4YiQhvMnjI+y2I0fJ
EdAQzzGMa4odKs1LTVD6CkkTJ5jNFod3/CmIEpPaMfKGBMEcSbgI6Xbzsa0T58X5
R7iVblcqxo1aJaFvbAZQKi4SBjbQVrtkYyzknOYpTI10tcUeODQBhVvuw2eJAEqf
QQUYQLxwYvKb7DyVngje4A1jxyjVzU5x9gXnyJrTjn8yg0hPBzM4eQ56Q0ufYT2e
CWfhqrwrIcPCEkw9pHAFLe5UAaAPopBZm+Cyghmgax0uuMsLmP09cuCk6qcKtTVF
zI5ZzrunLoZ5HmSkxzMPUA4UeYUT9VxMtIxzE+KhNJ2HgaHUizeloomISt01pZoj
TGR4XQrK0cMmUFJJnM2r+9kqOy7AALqkt0WdmiqDXqhEVfmerTkX5C2jOBhkoeW1
rpXjhr/Js4Sgrk9wUGHJZWlFxTLmm/aOgnkbr6tdcMpmGghVhevLFarNkVtgicPo
SQPNdzuV/ZESfErUQqHjbvzbgvR3Iz5Od+mICkVIwraa2bieYnYIitAi9ugippS+
IuYC+g6tg+t9ESFVOeBpvdVUTe0sI5qrgfjYadyDVcR7w5+zQKCLqqPxlD+xxZm1
m7CjXnVbL5T4Vzf3zVgbPw4l9y20AfnjweweeEB4E5aj699h1SEHBA/WEUzlBdB3
tySPzcCFBoloH3TTZaYFdaqDdjkYihWJs3n+OTtgl8055bJk1b0YuByFOYS5JZuH
lfTSzQNVDqkltrZIZLBDuBvHDAPetRkoXEERzESuKx0YoqfMVmMcn0l34Vii/SC5
2sNJY088m/TvBHWTlJvxUswwUmm4EZ6OU8uovFelRBD0UTC3hs+2BoB3FaGGe5gt
x/SMGDOyKUMjuScW7KicPBgTqCCRM52Cug7LxqFSUe9MkqEtnCCg71EYhOTWbmgB
b7TAKxCbhkR9Is6yXPGKo+uDVciS9PRtAvggOV6ziQnnikhox7m1/NpqhsYjI9s+
5SE6VpL7x8TZ23rVxtDhhxuMeZE3FuUw6bEofHofpGUz77Ia5SSrWzSOVXX0xO6w
ixKpLezKAPZoHMy0q35rY8sJ6HcMVfQN2PiODqrnGY5xg486OLKjsEQigvvn+vpZ
WpGq3/q6Fz1EXx1JVGaa67T3AiHEnsleRUqO0NaynPejFhncynLe4DvaawZfBfH3
CvgC5w9a1PQQJTZU876FFEeH6Bweqca+WoFH1KD7cgzgg9hpssLmAOXpzTo/QuB4
inUulKaUXFHgjva1e2sg46ylKTNJ/L6BFhwg6h6TtoML8AdhyPb8MjP07QZnn7Jn
1NGQN61HXpmPNOHn46IfB9v+eb0yaEli9F4zFfYaTE1jILY+7BOKzMwE7rnao7zE
OWqvhFximlAN/5PqmSIVbzJVClJ08AALREX0N8bUNgt0QBYrhAHzdMxvBicsIC9X
sbtbC0jpwCrBofmY8YhaPo3xI0k5FF+WdaECzbiOSR5Hy5TJhpLcLCJisweMSARP
uWFosZuK0rVtxID4UEjVQby8p977BwowzQfJaoi7uvfD1sBQsUIuqhv5iqxqHKVa
8RSfbvVux8KmYjvep2VjOPuvNk60Hmvc4kP3PrvXoLo6wBemNar1U18LtIIR+uZ1
y54jh1jbfW4nCxNsdwruwGcN8+6EMeU+PI/gn4TbSLTtIOB04Nttivj8wvujDYvC
vuSDdpN2spO4pxs5P4OgRClLaRhbSe53mFrkg602GaMfmIQrBaJ3k6scfv5oYKpm
DE56GcKURNC3CSSSyCoivYGIpqCZ4TdpPLBaVaiU+sJ9z2hfLQYbwMyhkrHOxPdv
JSeXfJCxQ8DpJgD+2BW+TEBgp3qs4mfdj7vQ2aaOH+WC7GRKFBVU0nUapCNmMKH6
PNnvDADhXx+HN1T6KFtFisuEfUsN88kmBGzXYQ451ws9PyvEjMIDiHk3RLjkVKYG
/jiTo/ljxUasCq8Q0DDOiWK58gph95nSOJmYb7SmL8LbW36PBaselY8KUWW/9Him
mUOBHDyRGndiQiPzGJqVZA1byuZTT/8wpW0iPkaeP2GfsRXUz/4BRwN2y2tkOuSK
Eu96QRFbqRU+87tkTqKc1x6vXViZ6YZInXl+DheGGAXMXfphUuil3bW1OhB24NuS
9/HmP71fraiCdqW0d4G9rZHzFmIF1R2YzUSfydkeTEXqYJrd/iVjQ9ET0xXOZixQ
uvm5tdF9LiKYiZzDLHXdQa3HBcWFZL7pfBwOpeTwKJPlQ8JIGk7xxnIbaXPu5uDo
SqXwlX3AQcAml9awyla/nAeHTl/NDLK67gKO272taqbA4ZMODzFOiwx4W88un/yr
kWjbfG91LYYehFzTUXWzmUwIbNM5HgF0KS8cG1NOEGTwDeiJai8pfDhFBNv+CRZ7
3WF62/UhTzL7CdtZ449ez8FeBhZxWj+bgEP7+VJXhvQcneOcfA7icQjOyZoeR4uM
s3jGLymCQ69xrfUKh5+eUoBrC7mdv+8MhJfz91D2ggzWVIcE/DXUu/4nkYyuMqCg
5HHWQop8sPeCIJK+DlXjAqloZhXxryAwSfDa9ghJvWpCUBGVLYSSQxB1GQ4Ubf/P
UPT44MgN1EU6ZPVlOPz6svitUh0+FdzhPALztQGALVBcBkqHXtyfVC936mBGlnoM
vyHLaCz8KG1KTPHQ7t+AS1FBW4N1yK9BWOPsvDm7mAfleNhIn57ZROHCYKv6Pi0f
DuVvcTuVQcGk9whs3cczotpEcgMzeKtI1AjrSypjuNg9aHgtaM4VVyzA8pTBtA6k
UhGD4PF57E84DNMkIaK0svfOyYU3v6GFHBY1yy+BQkO0HIuLxuMGQW+CEc1GM8g+
jZUK6w2ykrRAKgBkcRrOxKTpERAYpXjnU0hQDCBgccOCwkSk1JJSbXZEQ/St6g33
bdYwIh4WOB7+TSM7Z9Kt8fdoYOWSkFptp7CLeetxgxlGF75a0Kd9Yzk7srpgzoCA
VhvTDqwCcrz9Hf3Djn5tuyisL8FD01jvtEgpe4+QBcFbuRKA7CpC9dG5joVanec5
h6UHT43G0AERZ4TNfA4YwTDh4MQKjiginNZL8giTj0Vu7EmpxZHQHsOoTboeHv4+
ldw+ITpjUFSUDhEBAI7bWRRmF2Imh3Mh0fnQ8YZBnUjwdXmf6PwaCnhSOJLR+jyv
ZMD2Eu3FXhqrqToX2qOxM5wEqCBV1RKEm1/+Piz8SjsFwYbuwTT5CKPOyDOWUuJD
pIXebnqkXez32Hv4AE3tMUFlHqmhvby7eI6CDrOUOunbJ0utAkBYRyiDsvdvCj14
Nkod1SKT1UgTDyxSgHFy7kkUIZPVJ4ZLLptafKRSTaHleJGGQR50rnUr8TgVfYvX
AaugCI514crKYjrZgKuen6DT7TNCpBPI7cZcCiMN7a7XCk2leciFLLirSv48RsnN
ni1qC6oVt3th/oFVlKsSoCpDCAL4inAgFD6KVDRKzylVq9IhsDxBdObMqUPiQoyG
egWTORq5ePOV8CgYwr23EOscHLd/sKfynZHNVpPKyUiQ8iSagEORWbw2FEttBDap
xQxQgFlguCDXC2cqmE67aKo4ivr1+g+UCUX/3OR1pax9oaSLNLybP9/QqhqzdH68
UlbJxkjGcBj8ZE6U9bQ8V9IFJ84qtWdVPgQ0T25qubihiLygCxa2+Gd4EX6GqDMe
x6HvV5fnNmHUQDlAODRQzvVD4pmhl3JNYdzCsRejf49izIXB2Ci3koGk9O1QBRRU
NdEq+NZimjaIdqZ6ZQMLqx9oiPUOYywtmeMDPwAbXAST9Igtl1GuVoBX1X64c6Jv
06WD3EIixr93B2kODfVO/nXB1D0nDqOMlHwTENpzZ4DdWF4B1b56VxCgBohvJWIl
RRDmbI9nLJSF5ISuBBJEiPxrnU+YmSCSSRhvAa9T4uWZGo9puzlmH2lJtYHRmxLu
0CnKUE/W2AmZyuztH8eAxb+LpqC3wy54pKpZGYeM+fyd21PnLiCOaRnWLrTy87Ry
h0i7QMG4bk+hyw+TQmV2IjE+NIJsfYko9iTHYXU2sMea7dRYZvYhpIir3aYBMBmn
L4YP1nm87E0CbmcXtk28U0BaIh9DaN6ncGZ0Bo8dzVXGh0iY0Xq7v6C+5y00mnVK
TPrSTexf65pQjmS9mTnyw5PN6GqA6ISsewflJeEDaxzQRwRjSQ+sALIMc9WAuhh/
XymWXxRpRb0YTa4yRXa9af5dyLqnA4iw+u3e7nTp2RlN49zq9mpB324ivvCLJCyY
CWw9SS4yYR60jMLZqRRx1hWEDSRfJs+CugVL9ejjofYjJ613frXUrQqsGr+BD+8K
G0JNoAaPSdOWEDymHoijNcQ9LYpFbOIvOooZDyIGYCzCbSSe/aPu8oahPtJj76Fq
e6m3XJofW0W9C/19xxfCLwzE3JVf7KgyN6InSoewe/HlKiyPUPapXrYTjRmwL0fG
7s38VUgohSDreu8MktprSu8jeE4RBIvntN3arFFiIPZaTsTWEpKrw3ksxOKhSgUc
CkJKCO/P66pyqbsISrV0XA6fLtzuaVIlmrEsoUANONP859yrO0sFZc3Y9rhPGO5V
jRoHp0S7UPLNbm7GJxN2sjv7yOUw/5nNKSnNdc1hZaA84uENMPCzFN6668v73P7F
sU/8JOu8Mh3zwokGJVKfzCvvF8m1OmWkR2PmZI1SXVP2rv3C4gOb4xhiHtOAp86R
xK38lnF1+Onjsd5PBtCpLpRU6LaHNYGqVznyBZUefsxHrQs0nxWMKyo7lr/SgXvc
B4Z+j7X5JWxowmBbTYgF5bGf2NIhfPWtgLroIhOTJw7f/Msv3Y9wG87Jn1WtOkhc
XuZ+0abxSXyp9jvXRGxPf5tnqNE1UVQSvlAVBCd/i86SaMnZ1OJUyXFdrE88Ot3p
lBcDwWYzM0NdAeEiAYtgDZH9C7mFwms3Anj86JYtoGzsOmnKv8VSgw2ASbIllcvH
t6A/daP4gm9Ur9WsPM2GggQbmGiuFRsE17X1sn3UdCUQu7t49nkCYd76bvE9oi1l
dqDsrT/pq6++kxYwQov5QfBbqISsNe8SAyb0iPMw0yKcTA1Vao0GliNKUFr40UsR
fo658qGtUsXgB2P/rYanLjnSXuPk0+VvpkbMoMMzmBeue1QlLy3NPdRHVVojtMlG
fD9lHainjDQsDDsWrxCO/9cIgDnTosV2r43wXmB5BcEz/j2/9M4FiPOcYn2za4Z1
Xe23Fjy2wOLx54Pb843b36KSYYgdVH0AYBqZAy3m7CFqniB1Lpwuf5hopcGQmyjK
1u8qZR90RUYBMU+5vtoTbTW2/Gzq8TtGhtJvv8j/MSo83+rzJUTiZkxtLXWTA5X8
scvenwA4fk2jCEomguavflgn2yYDuhC2nkUpJu6aQULr+hHVfRu1jpMF+bRlW4kM
REIXu6DbY9vgSy/QMsXYN+0GyQxu+ubmZ1GpTPwqSJPPJBTwPi0EvBd7Dkliw50L
d0bkmXuss6Plsc6ZtYoK8q28CwQ/VHObT4eBqgFKHrk5N4OXL/cLjWMzZwdeoP4R
ddgw2yqnVEMTues2R3PncSqgGx8FhwORJ3iU8TbP/oP0hJWkDmTfd6W99+/AXKPM
SC5PQjWdaeWrG8au9N+e55g7QHElL4BLMyn7p9Se9fYa9suH2REmPpTMGg3zs56u
XpbRPyLQO/IkUF2m9e31r3s7agf9pRvs+vQ8WjtcLp2+aQyCxRrkponggm866drn
HFOvUSL41jqzvEh1wafGkNxOv5O2KonNZt3E9P6u97as7nNuA04QBx0r9Jc43jc1
j6CelGpAdqy+IJwaxaBozUcHS4XlAD0hEECsq9T6cgrSM7hHzPq1gs8/7h2y7OD2
LoKQPJgzVV2u/URL9nqkBOxhI4SZWO2gQ890GBFUih44Hipyh+egSly/8NxCoQ6t
sj8vJSz4iUH3Bedq3brF01czPnNBT1rZmaQgtEiGAOHN7eMs0DI1OBoHSwjt+aSx
dSt5mn91V4tULVO3asLcp7C5dgMoWvnl9GuD4KZPWAUb/Y9hapkjQiufSau0ytbK
VWFxnHWf+3suwTF5dsas0fxdX3aFiIIbW8UjKINf1OOLSV5PLFTjHrZ5s3hscv5r
rnvh5Kiz8ENkrLOt3I8CIIFTrXgJiwYXTHPqhEr9e3Xpu+dGX+Xmtr1j/VK3UEgB
YTSjftUboShvZj3Y4Qoiic/dHO4xDPLS98ZsaP4IO+tNQ0EW8sgezqPYfHbHr63g
mcMD2rKxpq8UgywmDfeVTfjp9sson3j37wMEsPKRbc1klPAMKrLpN5I4C/WB0bvj
23D/b6PU4AudvLx12Tvk6AOK24k/wmhTGdBTBGES/+DKAzaEGa3HV7beR7fkqKnx
ceIk88qmHZFt3GAGzfhpx4fNQSVJ5X1pMYsGB+GTg+5Fws/5B6PnTe2gBM0TmikB
NCIf/u0ScZhEW3HAFLGeTYiF8GmtM+u45ur3T4hYnUApOrIsbAtrLi53pjj6MolV
Io5A4iS5EUU8KK/KHAdryAb6wo0xr+56qRVcOsl++pKXFMoAdy1mRitPU3ykkbyL
AhXVI+5eBanj6A0PowQJhoobl6L1+CBp8HZ134fnuytr70P7B+GG3lvu9cEvVKv+
hJHwDQHflmcIORjXyI0KVj62OS7PN6zmPrvI5y+9y1m5yZ1OstQH4Tr0snvCOsFY
y72jZzlaSAwNHly39AfXnLrVH2gZzhC95lIvCBHTKtTr53fK9CdbrNJTxXcL3UkS
TWtJP256FpvceRMrLbqKF7A6drhKC/6nsYTFEqmhYzXrMXkr2sJ2SnziO/t0+4og
zeHFVECBoRUzoASqxR62c/XMvDjnbnaymSn9GzMVSJxD10qyAeB3obq/pCPNi48g
s0S6BwYDPV2CdJi96DcdKHbFcryBKvULEOKM9OVdNZaFyOh6pwHWi1B4w9pY/3x+
7PWRkv2gnf+J2QPZfPlqPloamPRaV5BngZRKjB/50kDkrhFAwDZEdjEj4ztjXayL
SVhJcSFWYgx7fHrJDQc78mKUI6x0pq5Io86yC+1pVhJr6FpY8SGVl+2KveLUkzlZ
6W+05F1arc3URtXnX+Ns32siRRyp8PUzE0YULYNhLVR4SMHF1Dgn4aZgtbwSCANT
ae0+huMl2+KV8SrEL39NfeluIqCDINnzf9xCMgG65tqZ6kaGxPfvMkCv8gzhiNeF
3EXQtrnV95xzZI4maAoHlw2em7+OC33G66dbKQEq3z9PpxnhDFZk4Z5ujOj+oc/8
Z9w2n/GNE3sNpC2dUCpJPbRDnEi1u3+skyWKCokF/5z0sRqmGI9hnBdVzO5Sd29o
6X2rxiJT7upXN7tVcIK2aD5gy0S9anbOrkp3jtaHBoIRK4O+uZs9x7mX924Baz4n
p0oll4KV1JZnCYgRRESqb8XZaL9iit6fSfhD+RdprCuU6Hs3r/llFPIZZWZXtfJp
8WVn92kzfvQjFMD3QM6Bp1bzmYS7WTCtXJmRDpv5hnDCcR8rqDRwt9lomoXXQTw5
+c8vSXtQ9VVcpzxUz9OO4N6LWwtM3wUDZl73OOAY9B5sM07yLtBMESbROs17SC1U
YFRbObWG12Xo5vLhXoCTZQp0nq2PaBsc+qA1h2oZaCJ5YpswnnE/l+/FEkTDaI0o
mFhp5s0dX1IyR5xQCIOz6NJsjdr/buLn5nyp6wFfFSWtXT0f9mVsOLb4md7vj/Np
x3472GRSCWgVt0tspjNcPoi13G1DIhhuA3Fj/a0sTuzm+Jfw/+F8XL3zsN5scpG2
bvz1ehcJGavPVlTU2c50hAUUpdaVQw/RVm1KSjUgNC7AmhrWZ2qy/Um0iZ2BeqF3
W6Fbb5h2EL3Fa1Y21jAJMzQKSA8GFpOiGjjJ+QGx9HtDtqYMR9AwYvnD1u14QzUc
1JF0Hj7WqX5lk1sDjlul5r19zNva+cQ2Aq1FzWcZ+588suQMJ4R4UOAbTLVdGM6e
1LCGSCaLzQOorVnDr/B5vu/kx+LRTHT88GcC1Y5LaQp80CtTT/FLmX9Bp+l5kCNN
1UwPhTDBkuc2jRfGmUBKK70u84wT9EN1DBlRVaHsSoW3zLVqgxECHkdkQn9fAgBb
t2fQ8gTzRkranJKQ86ZtBgCOvdfmWgbEQOvLCwsVKnpVl62fssvypGu8VRSUN1nz
lET3oIF67Fu7dkW5hBXYEprstU5dMVkE+KM6e+RaUzvay6UhBqNIVcuJVmnlKxOe
sLF+zUFCuKy3NGlMGDclI5f/CanVhLPJZHfcvszg2hsuFB97KAiSkkRzYqLS0fM2
E07mGyGlG+DBfylP0B/odge27fYRJE7IdCbTz7OCer+0Mfgw8dOApKwAKItc2CFf
xsmB2bcRyRcqviq8va/Q2VnwpuFm7CA0+7ovkVe9wJhLu+32rfUAmhzrcqm7+fRe
pfWiQ1AaV5Khbns15/xcp6I8kpYnj7EmC62YKVcEahyHK7dgITrOG48oAgcyrRv1
y7ghOW4pa0ii31zQQoFD5xVW2Oxh94BaJLtZBjD5pOh25MBmHcMUCYeBnxUBPeEI
fxmqup15ctDS/jRQcZLmHGhuxpIldr924sPSvjJadVtuxVMV+6lwYqeAV5pVtj7S
EszbD3qynPAQRzskVduNQFz4aDoliAz4qwDrSWkVfkuE4ZWx2O1mI2F+fWpAWV70
qcloTG6b8IN3XxYDEHD+8E6smTle9YihMCH+H+X/LJu7RBazhxzaf9b9UxE72+sf
CZPijHHh7Ur4pv2Sf8XW/5OYFXWdEL4MB+ZuD9yqhNMoZqcI5gVUurMhnCa4+5dw
2dWCL2muy7m1PAwNWW3Ph58yHziZ4cegIUYWaRUdfrJ4ujOliSM423K3MYYLpmRT
BGY0DvmSz6pK7Df7AoRmTYjHzpLeBIWfIJN5opgFSMJ0iPKbvXJK+b1nNtjo3wcF
7R43Y2/ZBYQA8gHLfbprSpj4ixcyOm6Kpxn+TPTpBY0F9saB2RG/uG5hLuQHIcYx
PnByblR5EgIgoCSvzv1iCdFf3pISyNgsMl45EM0ki62No61skymRdA/Qt6XFVZsy
H8Dyn8SUB3pHudcjKj/zJQ8+WVjnwfGzaUEeYs5Ipzk5xCywLmDgCl6Ceojrtx0f
eU6iOp7MIZSWFha/8Q5UlN0m6zrehPPok8FG7352j0rcwGeyN6cyr6o4YP/gzw3X
t33xEWiCJ4WQoLpFbE1JvD06o1j79z77Cd0y5AsALKVKBq4oPiJIBIYq1iJ7Se7/
OqPEKExPTUgYJmhDeMGshELC78YBa/xMbJ6pL+5vAv0tNbkXvLf6+VrLasZqYTD0
61QTXXcSr8JaY2Gjob4ZRdXTVmbjRD819q0LCE5HIgrF0ypnqIavNZwDOORL3fUg
ZWt/Ov5YeDOriXjeroKgwlC20A2lJ915K5U/sqIi6bC7bBVyxD0an1S5+ctNTCh2
Ezi/zAkuE2itxVxABD+cR2ElTcDPCBBiH5IQ2i7WM5gNRdzFY1u4dPArNkYpO9jz
nCfB2VVFJPgmBZ/OmFiTGpjQZKYSaHydi8Zfi+H8k+eVKquQANPUtmJHSgmUEn+e
gUR55o4QnQtSRG4JKhdlW+k00LLupXXbyPx2LRYEK6rv082J4ogJL5qzSJ/evo2p
1nEa4+4HPxsWMSfKuysR/RydSt3WM7cAp1Hus8e2/7zeqpAg7ZhR2U5hmC2zifyM
E7EpKCLD/hCKvFimFp0JjU3xdmTtn0ut8nxCl1Xlp2Sax5urmUS/6jzLSExex84f
JF2N5W7vCq7luQLZluEAOcS+569SjrapWKwCYq/Dkw9oxiGFT7Sjg5y1nh9Wa45t
i6ogpm/8UkGkJ8pPq7pzNEyVeMkVoMJYtenjMtkCP8dgeJNL5n5/tN/3fF/XYG7S
N2pHFH5XntuXIDrYvkImMqbcDL3kSXupBNgqqdIqb7ZMA+Aa0IAV1woU2TJKTg8e
4x+3mE64yJPMEvew/798GIHx2i0PyrUkAUtPcI3tJPqQ0O4plfN4nF4p1oWxRt7j
Ae2bR+nMPmqmVeCOixFwkyA1fvwpngkbLXrB8EIIVBKb5KMbC3iFkAacwHaCmY0L
3yE7ITDDOT76hW/yFCloYi6o5DT3pQrdKNUfsOcl6J7DIxYRni30XlK6Vgc0ZamZ
q8GI9OaazedaF3AE1LefAp5H2LNi5ejmUiC2gVyi7wna5zleF/uk4h7kH7iQRKZh
lRdCYjgqZkUXwyIV/mPBPSCAXOjThvNFUDiQP+fCB/IGpuoe8VgiUAx6sW6jdiI0
j+NwdkKMT24Ohb9R961nJTK3YKPuS49PdggH3LKUx3bDwFuXyy5wJh2m4xCMAPGg
+RgEMmPvUDIcY41qQx7oe7HWAFPba9DVlIQTWKib+dJF6XlTpibuLZm2ENRb7iBb
4RAepB46iciUyPRhldGXJ/3CN4RLoEMmS19dnKMHo6oILazpANKKI4EpsQLPE5uP
VcthSonyumIX+IZHl4nxItNStieyW72ORRVGXOrW5i1cTP1aQ+2s5GI2LLl4Jyae
dqpjBJ1PuwhOlqzxbxFnpubc5TOUOLmjBwdefOKvt4Kdxk6cYLYWP4hJqO+N7KqS
TCWMLbrZmxNViQx3mG7nzq3MWtKqnJPHNdU5q4AYatlorYCKuPR8BldDtz8YdZ0Z
FawyQXCr9f+WCgnZSu3/T3CIhKnrmoGjNw5jwMKlbfLoWP+sYt7WDLyvlpkbxeTF
AtPf8O93w2qiQtIZ0HXLpp8TFlV579Sy6IXg9NS/SJHatbH6R10HrLO+6HZsWbSR
60VO7jdBReS9zNs0LVVOeoSQRxwWPyHI1zXz2XGaeFnRbMbu4YEInMqCnDhBTIu1
W0ZwPgUbJdzFzm0H2LAbVl4h8Z/YsqBlxw1qo8nKa+Bl4nPNDtsarIZXurowL7mr
Peowu5ZGY9jjFNltm9nH/vnY1SVzKWJJZa8feE/7i+6FG+Q3myZ9Y8CW1bvFeGYo
Gw8IOjLcgKU7WbKq+lsJzcPCgLF6ifrn9HCD+/8bHG03ipNRSV5zqP2P0nVW2fLu
9NkKcKH1YFyi6vDFLX66Mb9md7ZlkdZl7P8wQ6kYpbdVme7R0WgyQDXMuScibQkC
5OlKe5XezidiaTr2lLrScVQu7VOoMVIQr8oJ3DNCJ6nF52NPKCZcywfJIO7uSA2+
bJWMxM9mMAIgL2rNbuO4QqmeiDkZiIYB5VVHr43roozmmtBRIm/3vWGfGMHgH53G
EGLcHkzno6T0Q9PoUuCgSPXPnMQQXw8b2xCcCMmpfs2OJHPkCAudXiyClzoMPsCE
4Y9IZYb9l771VFgkHq6PMqIP9HiXF6EQdIzMiE7mDVV80vf8dVa5vkqPKYv9h4fE
DD84T5N6rQzcvjdSHjvuBoIUpYDvxadjJVROUA90fqXlUdyyhhCbPBMsVnhPY2l1
W1LdV6nOcYsqQInmGUUtWxIcTDIEm5tbHkv8f1yuPKySaQfqoIBQqMQbffVy1O5W
vPU3wlbez5PcrT6LaJ2EDjDNj5ijnTtBZMtJsClIslf6qW/1NTLN2X+Mo8smE9qO
E02H5V2Fl4NaR3lsquy4jlmkmfnxcoOyB7tkS9eBLs9RtXqMbzDHu94Q/becqi75
isaVYNQ+SZq1NkWXUZY6TmgQPtNnhEEGIelmJ7NomyExgE9NWpvDA+U/DzjjRLs9
1xg72251+eQxYnR8PRxB3vh1WlZdsgkolXt4W0C3a9YjNGwF8Sv9wx3zzXw9jtRz
PmwZzvk7CZOWm5CFQclhdLMojlN7ttdNS9FCjt+up+AqLzIO+MvEeST3CR3z+D8U
vYkOG2Mrg94YZ6cpzUM6xtnluXN8Z6hn0BlZmic5/RzaCCXt5gS5O5SINOnbrkxA
HjXuTV+Zdd+E/KPRdWEIk0pJPj6H3CV80QvaSiNIak+H9mgP8KQF5lBEh30SJhP1
9EkojVtMaj9Kv7Cm8R4Z0YsQIM5OQTy0HOzEOoP8LOaDLBORGsQSo0+9YKfDOOcG
IBiAncQSeOEEj7dgiKUvu8iP7J4Z+siJ+Xv6vyq8qpM6vz+3nEdFoCnA8Ocee4sO
Sy9RfJf+YVChRdITqdjoK1GI/Xb45hilSZ1XgHf2lDsbXxD3pwMjIy2Wh3mjcTPN
kaHN/p+gUr7mrSxODj4Nq63wqOFe271qe3B7lApogIiWW+wq6F7rAv1vnWzEUFl0
qW1NZqTH6weNqSeVU4bUJjRkxcw74PCkEvtNDMvOr0iw+3M6QKJDyr9PME6g1+Lg
QwtlDptlVbKoLYnxU9ZRAZN70YZn30FwQkaHnyyaTqxLPJwBfiMEjlL81A2a45as
Lg6hOqN57mO+sC2fFWqNcDZu3IiGV2YZX6UQ6eUHY3kVYBDFy1LBERLteDP62/df
s50cvgVe1POXuENJA+aMTCRRcbJQcj5nETmQieoxrqVjtBCwqmMPc1tfMPvSduB1
NAShSCnGvYqnik1/rmGCCIypViEenLT91VV0GJj5+C2VbZ1Ynwvqi8gZiJ/zMPRf
ZuH2AfqFDa5VnGRqw67l69qLUR/CSraPktN9OWtQNoxKwbYXRZ6Eb+VEPCr92h5M
MiGUfZi0rf2Urp+0iv4PYBSeXsL/Tnd9cXFwSz3JyR3fkpUtM0bPI9mFzhZF1ZYH
w1fHi4wQrzIUoSoGdX1Mnf6WnUq+K50DsmKj0ao1+dpQ0JEr/aMiGBrv1cM7wAy0
RzB2KvfnobAzdkrAJ5QEaHRWzdeDEflunDDgrwkFWuP7IrUm+B0r5mv6LGbhqrn+
9tkL94EuRgmQoGxZWK7LCdnXnXqbc8EgIbimQjHSFR16DTk6rBfY7znOKvlV5/8u
LHLhvajRRw+bUal/4Oi3s8I00BCJdQj+l3YjSWr/s+D1/2Ed22hDmrBjpo5mphQl
z9a6Cs/Q624FUXT+s0aQuQX1XxdWZgB1SMasZX2UMM1dOJiscUA8oIm39TwRvWKW
r9ZPx7fbrIsr32zPBKtaJgpeAPJw06F7BsFBgBnvzuFEEAmzo4mgf3ADuEcmijVR
GcjkozsuI8tTWYF3upjHqfuN6/Cg5wYBSXLMVAxEcA1ezxCCP/Oc84kgRYF0qH2s
56iOcwitsxP7RGM0ui2Yr+53gNHh0L/uHyY7p+otd84meFJ/SUlCHnxl0BWNoUsI
8pUBjW1uJvVBUE3HW5L+K9m8eUNez6XC2HLh72xaDKNWDH1OTR4PNJx6JDgvWkxM
vNcaGW16simunRipU/hoYk8kwCuDwEpLoGSDRQp/2iCbP6kjveiacPU4FkZO9KZ9
jzQWuQXFpjHnR/WoVTu36HLrjaooVJHccqqZ2gsrRD6WOU8ZGQdHQM7uZc+57VwT
/DiMEuYxJR/6x65xGTCgRnPPxerzBbD6yoD+S2TkTt4v5mZdZx86+xY+cgy4Sf/t
lGD7u+sVRDednUlzGn4TIbxuCOXgXvbUq3USN2UumigVrR8ohlI9Gp/gMG0TG4Pq
qyVMASQphJUhPELtC72ptl4aTHB9Izz5h7QPPv758Tg95c0JTML/RnrsNjSxVeC7
87VzJN/o7PH3Og3Xr4ZcYAruiBdWaalPG2OSvEeSdMSg03Sf2vuB7nNcSEzyWiDl
Y4OmNsXGggWbomwvGAnDy0Yk4s8xn24tjhDtN7SPOuC7chxi7GKwe116o/PZNUe6
zGBDdTwojJb70U1Gtnglt4xTW7IJLWam4phZtnyhoAR5qYoL1fJaLlWcB6Tk9RmO
bfBvCJ3n7s2vHCAlVTz867nWAYwoY0lCNBzWPma9Mir3TNlIds0rGztuzufDvoGW
/LCtRSP05WdCHyECoHSkcEcOOoIf9eQRCg4Vk4UnoaRoFJn+gTkqli0TET2gzaLL
gzxb1r6J+8feTvQcKou+ok1l0/GGdpNGHehs5vWkP6hz3xXOWlk+1XQi0f6tRDen
gN3VJaxGxsQ1b04lAd3LYKg66p8Yj1BK46g2zMClZ0ejXcb7GHdqTcEw3ejMdnDn
Ces8z1XIFnOgozh60qPeK12Mm7Iq+zp/VxEbBD4MH8dgSWX70XCFWa08B8SMg5iM
UfUSF97NtkejVGKPeYMqUQgRKkEp7Uk3fprt4Myxj1HX+2ysj7qzZiI64JZDK7bq
ff/Y5fa8cggxVly7wPBP8VqK8sEmtQ+NiOhrqxF7vGziFvdgii/1XAXLF3Tyxzsv
/zHJnF1Ix83Ef8tcSU1EQGwp32xwn0aSrW8g1uuCOH4jY1G82JzahQ8mAK5PW8L9
xZnxkfc2onYFGe5pYM3X9/54E0KxVJPPAOQeDVS2Yxsy9TmzIXLWk3qeD09oUksT
e3BztGK8RtyIYCrRgNZqX51nKzoejQJ/VBs6gUhZuOsH4GP1ZEiO5fPq//kKF1oW
ztSRrbAxlwWh8wdZC2EiA7JTE+916OzaeXTiqEL3B4AzUTTEHTkGGlaY59IAza0G
bjvSJhQ5HhkbpB7qjknZdBUS+N4f12+n1UtBW4Oa2FEqDZc1TXUyUCy8b3jLZ7Lm
2CubwPfY1SJ+6c7Xbp07uTMVyD19dKYvOuLTC4ai5a0Qsxbna3rR0ZehHvCogBXC
KZdRgXF8yAEZURWiZEY934mGjN4uUNz27g1cwoqMVU9m2Vwd4q0D6jVlDzY9Y8X/
/GeX1zGyezsJXuXO+wy0EYYV5z9tjNGNAoTsdPu76J+52nu3Zpim8V3qS/S1Q5mS
RDaQ6YnGAPsZbJ2aGqRQeNwI+9X8iCmmFRJQqM64UHpnHkZ5l8hyagqcg/Yiwn8y
LK+f6/R0YbF24BV1paE6Uk7KwOvsaEJm39yGrMGEMB4CANpPzXkgOyWpRmrWx0Q1
iDReUv5ySqbsjPsChEgYRpmDlS1PIjfsnd3jmI/2mYSJi+9UfvG4YF8OuZpB/aYX
aKq+VhokbOoFemEF7zTWj2vaPbS2qUjeGLZ3FLN6NCsELvQ/iQ9gnaUw6zpp8Y7F
Gc0rMJHDlzENbtSGPSym/urGf17U49kyIZ1931ZgITNXn292K9+ZgwXtu8NijYBO
6S4mNMP9vVSZ13Pk50PrZOsb+/X7XJEe2+JmCMYreuG7ECj0LHbuA2WCuRB3u4IN
/QYWlqTEslJvBmkM2HFZnaT2pNSKr3/rifRBFwMZMDXZEJR97S8RD/SjbtLV5Gqn
vhFJjHQNAcbA+6psyFGKRgPmkGMpAB3SmM35MugURUMK+QWAt68paT0eIFWgXLSg
9/PRkXBPlIpiMCU6pjRIIiRduYp5HrTJ8PUv3fFmnEGrsoaTgSqoDQvJXMBOC4Dl
NFdj0tBQpdDGVhgK83PN9DXOwenqsoTxrwQYE3y3M6tVwOde7i7TE9JO6N7HaUVT
FkI6kz2yQC6uf2CNR4zYr/aIGIlj1/jOw6dKo0tT86GIGJ/PhAAFkGLG3/HLnJsI
B9zVZeLIrjQRX5nGFdZC54XGIje8U+25qcjGFgi65x6N7P6ylr5gnWfVASk2Uj/B
PigzhFlimeoprYTMvm/dFGcwIWsvq9HXEmqtLGE+tF/VpMfZyYd83bEEfUuSRYk1
cpzYRVvwkT2HU/I574QhAssdFvg67ih7vFSBfRFixt6uVAAIxLtb/yWuXeDBEboo
evLxdyEFyZZUICOK4rzW+pH2Tm9dIyRh3fhFCAPOgSMFGciYhoukkeET08/08wvj
WNITzVdw0Tg1YUx438mIUUjLjb4H9zaDMqYJmESCxIwi+Z9T3DGkCQKJVaiu1Pbq
yQguunotk7HCYN5xjU6pVpZJm2id+vm4NksMCY83Xr/Dhjn21IabzaiAyaKQZCo9
9hg9qXnyv4oBSnI8i+1zn9Fpck2YZwm/s/zEMg8u/f2VM3bS6Ojz1XCvZWWSTBYg
M6ghOeGLHydxf2V/ooDUQD8urzHm8+aow6NdsfzOyKW0DugZQd42jfDrJMGuBWdI
08R1Jk25oYVd4/Ev9TxHLZAJU5I8W+R04Erd/6MJ8+nr+P1ISrOA/xtn3yTyEBFq
E8okVaI7tlulU9jQGjrGnQdhv7IPt7CH3FpY/zoDru49SKwl1m0Vi6CD5/ca+X7H
9pnf/4f1Y4cDhrz8TBoxX8vI1m5zkXNhIdZ2mdabwRWeRL2q2iDdBsZ/5zNV+Md3
UOVeMlfruBlwsOd1K9QEb2BO/QslrX8Xp3825nE+IjO0OrOjfoSMiaX8UFyMXwAF
6U/kVInt9ln7IsRHY5II5CQY0RW1cA7B9FE8XcoUcmPWA0WG6kFDbT/bQI7A9C9v
HFh3mEdnu7VwMqp/05TGDGMrI/2S9hpjpsw8kTdU8lPjeigil+Bki1fu7ZPq/5m9
+tYT7uv9ciBd2hPQoM976ld6VXHks3h0o7lvwNaLoV4VBh9v45G+X7jMPYKk99bn
hg8ejz7AB8QsmXINpqIwG28aPPC7kPcU5SH6QCghijWFNK+KwKUtMbWHoBi47lPr
5uLIToS8fXWEJrYwl2JFHvnnbPnjXT0A1v5g7ITbBmVQveLgsmLwSCoukqWdCp76
MCNz/bNFJ+Qym/M/AlDbEK8EK4rQ8DPgJ3ozf1xRC3XnqNC8f7bxvOZsQAnWJjzp
0Sq6SZTUTLosaIKVZBEbtRZNsRzKD8dQYPE3ttwbDZqk6x44/wOM6u3pZX/qFbyn
Jaz4O230GEtRLfqsQxz1oVo+N0n5sbUukn4599u2XfF8LVaEMfXhbtuHGVIincqM
fIrxqZ7M4ebjaV2XE+xIJIMlrNdRRbRUZWVtiqv2oaQFGe9HtQ3HBSYYxKv83Hab
JbXWOERLvLsYHF/PpJQyiFYdddp52OvNmAZD3lrOqFsEA/XD/urm5PTwCTbcHhE2
jFX7XFM6jvimh1qJxakR5p6X9WPrMU544c6IF8VUYWdXlJwxokJW2/1rmYLhgaBL
IvNCyipzhCqlGT6oeqTaLx1uzofnvtuspaRdrEqjT5TeYgz6C8Nuz0S7BHCXh5ic
iZLh5Sr5ERjKLnX7C2WQBx4dz1+wykEN0+hOvu5kPNpkT2qwoeVct4bF461zieS2
iv9m5uzFfZERwRAMjCpH1/F+3Jehs9zTmlozH6wuzPGJ74zLWK8uhgJQOVaCPOLV
E3PWdlHTk1ivym4RjcLzBNvSpf+P9AMqAKuJFlD9ck/lDDDk5rBL4NNlyZlzMI5Y
2XQNsUi6ztRDzlQt/U0JHXeZlKuAtZfOt8sillk9Nm7s0XQjfG+y4eRPENT2RA3f
oABBUwapnXPBJvb/1SDBQa/yMRgf9MEacur16WhoZiVmvr2c7+DNrlcN3toQSo4Y
TrzG+ekksgkeuKx7CJ1OzjK6EMzLcKm3m+FXGgY6KyqnVB8gW/+LnvCkgg06EHTY
EsA2BG8HgSQnxc0ITNcghK0Qtb8zO3O/2C0T6H4ZMXZYXo0xt7QOKALXtuFkfO+5
ZyPoA1ETIxuB26iXM4x895P4t2nhBW0y5u6igbVQ/PokBepo72u119pN9ZTCLduF
OqMnaVTcPcc+lU2Z/pkr8IlMvOB5K7hGJM6My0AJCJK3uuKBYB5JAIrqdQnL1yQP
ixJ+0I7kaOxj9e20dNvS9+A4scJVKQRHm+kbm7iULcgCnXTDAavlm5C1kVD1L2e9
f95Mqn6J/Dl+8DOUPQOlLTu2k232zmSdrPjCxr5x/Bu07iRF4wtldRsYdDTjgisc
DUR/KX4hff2A+SVVLu5FW5lFJTxlp1bzckkl/YxFsB2arr4q3bmKo8iTJlXSJvON
sTcoIps6GdVzKMAJu23chzl8FHsZZbo2ivb8pyBi7XjnQMsrPnQyajNLqyeyNx7o
50pYif7BbJ7BM51GirF772ONqmZQ94n1Y2qllBo1IUrmeTlu4ZlHYjiEwGjWjYX0
PC/zV5NOwVJcncQ0l6IIxEvXA3z0qefmJd+dZZXFABiovHUUiSQIK3swUpNSZcGF
SsjsLoW15XytmgRzEaICLGDM6teGv9MrPn1cRed8VMmKVhLjR5PkR4O/HlEk3+fD
i4bOt4gV8K8tuMOa41txnUb27e35qBAln7qPPoCA6k/+G6f3YdINKDdVxaZ1wcBl
bGHohLe1FQHUQBVa78AAzjPg476JJ7y698eCgy1bugD4IM6zAuurDkaALPiguAB7
WvFudP8zH+m6tj5As8Z1pL4Gh+EOkQDZebtSfzPiU4ttpT/orQIOPMj5m2CyIe1Q
R0/aGRFSPUIAMwdzUo4k3U/UNHR6rgfy6D0IWNf9R+8E9IZxzhx+drnOd1ra23iG
0A0r4cpawJylnxPey++j6jamIoM64xR7v2Op/ccY0151Nqb5FWgZBvu6vj862S1e
IhD21hHPH2863tvCxGeAUlTVhCXQdEVriqzRiV6NoiSiDy/KKCFvBVK+ay3tkuZx
loaswwO6StDQ3pse6QlkRbYDdOSRV/OA9rNgJLhMsZcyNh0a71FXkyxqYJlFd65n
tPogPkNKmF2agI64pgI0LXmPGpeZgDEaza54zug7gGakuArblgOwFOSfzrMHghQm
v/goXno/dzGk0copyY+ewaCULRwWF1y18O1SbIgZCaAzMXCBRfulN7LVkVl7pU5g
mXei1e/wSHvh9W2fYgaBOQDlvslcaAa/UcQNF2/KoDw+KMzk5WktvOoJfeSnYhY7
qiwuw/5tfXoVQ2tlmrCMHcIKTIr6NLZ0NV6p1J69KaohruBqiOWrMH3iSFeu2dJY
hzjGeU/bGU6w/s5FwCkynBjNIUatbe5+yXaTlsSXTA2OjHucKUsFhrW3ZbK5/+JS
GuhcEJfDuDfj/dBWVgbNSCHe1BrYF62vml8y0DX7kc8fyt4FwqMp2ifA+4RJ25ke
X9sF7YL9pKFkogqlFtw3wa9320EvBLCTQlaDKwzsaeKZbD9lC9NJFlvA3fc4jGwd
njU0CzlKbEVHinGdgnWlqkeGmBwWCqOsW6hxWpm3qNxVvZk8lbcAVec5JKQAO77u
XrOnLjiP3ycVX/hg0zTAU4A/suU+Ck0OYyV9bW8/NRbJIyc/lph3mCL21JcITo3Z
JtR/xhvn5Q/rgGr54BnBgzfZ9b1HKLaBQUS3avnjidkvAZEfhn18wfdITdYFzf6j
EURQFapn8um66mseCuHkPH7e27Zctn2BudDiVYJyYqvSZhV1hLwJJ5hO6ZvXUIx7
rvf7wYWTf39kgwfeh31btQelKJ7fJmT+F4/2HTchSzjtmPB52Ep8bWGc76Bl4pFG
rLyievgHMQlM0fEfxq94WwzQOX5K/F7fTisbR36ZNoRpDiDrpEZI26hO4L79QAVI
4x4E2XDRXOuBSl0C4Uvrt6/xzbZyW317Ba/ZSYOuqLOq+0d4QPpVkk9QemiizorZ
lID3jTtQbown2ADKYvdzAKSbBVObxJwGCkCSW2XHlY75Gj/2KZtFptf7pbGpKl88
kMEAAxnhLYmgXUMqIaBZ7EDq5CtnwO/X8tD1Tu4Hx8zHVVKlqQvW2zoUSJEfYB9O
4rw9CUyKjqYe1CUF9qGLYc52WHgr3GOQOybO9mCAQF+mr3Hc01CdJkZAzIQf73aC
SNKaohZJBV68pQ7gkqr/Hb/Lgn9WH5dmLv6EH35e1o2Eq5P9QKLdrNre4nVO4Z/y
bEUPS6/TJEAj2vpFGeVIMh+2kePx9AgINsXBC6m6mFDR5HWqyOddw3xB2uZzeadv
9zwcTUDB46Of27dyZq8QGTPHnklIBpQ5yj+2dMy2bFJVrGrWkEQgmK7VkWfCsZzh
Hbf8LGROwifgeCbRFPT+94YFF2JjXnuMPsNxQPUquXwDssxz9FOBXY8f751YYEiu
4c3h3RWjafMBRx6mB882ZDi3OLPahC2B/9g5hhM/36kZvtzv3Tu2ZSfaUeU7xTyy
38FzijJThq+W09FOuZJLfNWPiGKHkOrDv/xlkCJKYK1w3fwo7UKUHBXMRxwhWxi0
O3c2fc3sNclNFa9YTp9qYZ1cLrRr1hDIcrU0fjDd3zMm2pWuB5gh64fVpsjb0rxM
aYYjHLR0TmqmE+Wh1L7e2E1Zsph7Sg5zhht1HDNKSDegtmmvzJ5hNtOK5den6e+a
15rs7ephjHfSIZAGomKxS0M6eNp55VLhfPCn+HF5fn14yUvDpffOZ0lAqi72MVq8
i7Q3WiamwSn1pRe9FDpLn1nREM4alBhHEwX3/4du3aPGV/vG/nv0aBJ7Z6MrNPtA
U9K2Rzo3vNOTuxnBUC78/tl67pcf6Hz9RWHRsIztZT8k5wAjRxUL/UPZ6EyCTOfs
qEtkerUaipbFxetf70tCWijSXN80PtqGR6bC8g+g5l3s4+L3n5wOFfJQF0f/63gT
jOJiYQftbt1dJOfL66TbMMLCA+0z4NmtcNmD8wYpvWk5pJeczfR/ojw29VREatZH
ba972Cu9LNt3h+skYCcXjUqLCw/qKgmubXdatZ4LzTrzy8d8nYmeNNdfx50fTt1A
Bgs3G3qZWhtydMsSD8xDJODZN9zv9lGdfJCYQc4lvE6ZvpwQZp5GQXU+PH0mXwhe
644kmjeahk87Gur/azdIAWsa2m5uEF71ZD5lhEPGjdopIZVnEnwSiN3h883tQNij
N6rk4QPVUXTQ0ChTkaPD04CfFtGSy90Ja+J+DzVtGpmRRIgwLQ2SVStVXb3eH6N7
Re3uliyo6bTiusR8GlEh0SPLRC4QhPOSvOHB4OXLmgTTbyPs6G9qdciPmwn1HADz
4+a65Iuff4BM7KTHfnoTi99dz6Smad8fadDGz5EvLK1mWayEjTPQhXml+EZEn+xU
RKIHb/m578wugyXUZny/O9yW5hgikWgaf1L1l5UMiTWS82c/bB8W9D3K1geUnxSn
sPTjZ4wJtDJqqgUvgdKjX3GJBA9RMEwopE3pw4NfL0Es1lTzWdCxEEt/Ej8nVRLW
0e8Oy83YMfLDfx8poZacs1fZ4FOQ9hynyN7PN1tpg2sf2ekHPkk2F0HMFKcoJwGa
sKGnVnw6gX5Rd6B0j2WIrakBGYcidFKIlTFyYk/OTqEG5yY/ud+kM7YnYaYql5vg
cIoUoUpYMvZ7lLKvEC26KdHinkxICe1EGr+gaAW9FIhhDCADsIvwFkIeyZf1YHSL
7kQBJdAo48eh004ItqGFJMTbC0o4TzbLKoGgLHYfCh3LN1U26ppwNkbeOpX+gcI6
ebjsJZbM4xROH7N8v+PQ1oapOGtHd3v+XIAghYZp2pDT0s1E4v6u8kOmRaL5BuwS
GL6gvFbnu1cKPAoE6P+4fW67Qj64QzqZ6ryCr9EO7RW0kbJSTnQZs/5ZoxTyjZ3w
EJg7u6jhTsRVv3jIbDc0CoUKP7zVR8BLe9iCB28ELOGKSrMlmjiYw/yKJrBOPu7w
adOZFlx7gEqQKCnSjtADj9wCQSZHQt3Mz78vOC8SK4qvl9Iy4aDcdJIx8vt+vgq2
/tVNwx1NOPufKBoI5ehgf5JkJnlADlLdqjn9BjWvcbsJ7X5QzRe0bLcrV+WfFhWR
AmSjwjR157I8TTB61l91vWuAqvyCTKtWBo1gHzh5AOTNilkddF9/3OLvY2qVnG+I
w8EEIeXPj2w1sToNSVY4fpTe8/sRNYr2wWqkDKljndWd4jFrPbtnIKETG4rvuQVA
vC6ucjhRWKiuneijIaaBmd5I7jaMCKk+L7OkOPngVc/KCGGpGqBCniwqukBhU5ea
9hVXeW4WjLAiU7nF5ZqLaar5e9jIt4MpT+hHTDqsMdrDiFrTnJZa3kfw0lr9ZfYg
18Wt9T/qDeTy/qKwZwF87/zKPV9Wj4kt42qqXN3uxMlAfXnU6FQ0jpponJKGsGLZ
9FYRI21VWp2FN3N/MpvyJDnXY7xPHmRVQja4mcIjQSxNswhM+h00YcD55uw45CoR
FrE4xtRybaoUoXcmCs/EPGiDSPrspkG3Cl0A9QyN/10wdwZwFqOw5NFQHesdCSYo
2dHuD39/AcN+ZfupKMNZVz85P3BXIc++TyI9CLR/uP5JT06f2Ru/bM7O8C39qgQ+
xXNYpOslWDGfOuC8hr4vYWLrIdBJ48voIQsgp46KwgL34SGtU1bukxhKZimU9OM7
CBimgNPst4q6dyAgyT38GER3M34FQRF88WVXB/A9Yerxw+GBMWYkQ+h19QrZZpRL
u6LSVZTBpEQ0oMgrU/OLeJljXfxU7qwLFCyWDZVzZ1vMXwPzAqBNNlO8vdQ1/QuT
K+8wKkT+8mumMx5tuzpyJKKZsAW0q7Moqg+wxeUTMYM0XTQBN9FYvVnTeIGf9GSk
PWumhxadLxbpHxxDS6uRoyjvbJGcehpPbF4Bj9IC4HSOs/vvDDEXc3/OPFtPmNNK
hTiqByvc+jhkvpcvoKL5Oek8NcT8lBPB/P72fH+fz6dgqbiv4spTctByGwVAHhvH
DgSIaL7TDNooEkimQhGr+wtIkScBQw+silW9Pub/ZAgBdnIFLp/yur8RJaInLczs
jnd+0ujvDfETWDvqycNrsyJvuMHKqACRr0mCLidCMWzCWHf4b1cJe+h1a4zVbUR1
3QAKmkdh8Xc0YYxyxcW1cJeop+G5flVMuQTD8b0TijzBoz1Pgw3y6vfTvIb6MHQ3
NN90aCy006c2h0pvxOGA/TOWOFghTeLxSMBGKJIoIgpS836WcdAZqZ0WQaN1OB9+
nLdBAZg+CMLHyGR+Q/ui91MxGAR7HtgJHZGbmM9pARZMZJgLejXfJG5ZcAxLi12n
3P4RXqHapOlCcv+Pngf68z60aKMi2pOHIqk80xggy/R94/jdRffqEi8yj5GJpVvr
DaX+LHAUF0c9RdAkcCFRBlNRH9MRWRfsR8EZTcMv/XuCFjNi2tTER2QkPIQnMbv9
R42nfcmuDBf62ybukvfg5PY+6sV1gXTbKtrUZtVNzTJDGVLLrXPnZJ0C4dC1h9TC
TxgZl5ToQVcrWGrcyTQQVCpke61UqIC9zLRetLSSMLzAbw9pHlN2+VS9MapJPdpB
65l3wGZsiDYjSfH6+E6DkWxBSAKFMV9cOC2fFOPofYA16DnzASdWWPmIBY3w3P5M
qBrFIuoY4W5td56/P6OmHrVGCCytbHm/7EvQKiyX5DJALjrZdUSsvfVVfdI/7V3q
LDwluh+v7ORJPQjUdeQ4T5tzsEYoCvaDzBlpTCTim85We01Nb/ORfEPwr3fdjf9s
JV9eKl/cbDyAG/7ygEnoQ3wj7ZsmtzoAXsGQOz1U2fpHhgWOtrjgbWiKe3GDre77
u6ofBLftZAdskg1Gi7z1aFDAaejWqN2/z6xFZsv4Yvd9nWYlVoflm7qYTG4sJHlj
79SE/W8+HMbqmC6cMmXxls638qf7dMFFreVrsPudv6hVmxTnzQ6WpimrL3p4tNSu
aXPTfRw7fSFj8CgvHXzODSK+vBc+4r8iMbF1jTvTFl9LmFomZI5WBcDYslS7GEdl
XXz+x4YL/zGI+U1/MtV78C1qbvNWrDCb8JlVFTZPI7R3j1t5QgrlTk0vq1jRNs3W
MPhKIrNpEuKj2SWUnrUFmGoUcR0qyERKbg85ArDMdznllMfLeisVOn3tr5LAWr4X
o22e49RrXp8++7sLicCTEBlVmahdRdSmeR6Lqdz/iV+3nrC3zdCbE0aEQfdwrC7s
zP5ujpQUqFzMxlbnsVG+M14Vd8+FJ3ZpDQa0UNW5J/MH30ziofvYev5N7k7I5mxV
LQqMxcJ0ygxiQkzRk6gk7GYsODAHdzIXPxOsQOZV1fyLooCE7CVLlZTEM7R0OTsS
qjtrEnnLQhz2+OlN1sTs2jItcJiGCxwpCWZ1Z+gtsfEJp/TV3Lyep0VxH+talW29
iT/xChfX+WHh4dakcDrEsX62YfkwdzYj9miLioTbeetIKCF/JXzlQiB/QHACvyRB
KN3Kcc4Khe3zBFH/Qmtvo6SU8YtNkg7BFN22+7+F8UrTTlg0Cu1csvti/hFUo7Ir
6EdFTScLTVzK6BGHT2/FhirQ15ZP59JodGptNpdgHUQt1O+ZI4busLH/HYRpx18s
2eqMKiUWmxL2uXJwit9pKFLkefvAZ5G/XI+w0YkDqdy1wovtOs0LCgfV/uq1H+cd
kEkz3X78Q6I/GSG3WzwME85XHwjgyuvAwgOQ1oO4tJ9G6AfBqxgl+cCduIyT6j0V
b9HpT+2Um1rhFATA0aYRpwTrq1ylKOd5URVHJ0z3N3vmmpmaumEW4kJbjBGnic81
BtFHgluARGcK5RM9Ulu1B59XR3Wu8dwglwk9akG8jwCH2gwH7MC5Rmtn+yQlHZYU
ZTBXfzLIMjn+6/OrjmQLnBWOVrzKv4pS4xILPXraV8rtKbNrEoi4p+54INNsYT82
BrGHh0ijd0XFOGuIAeGrrEWGHuheZmC0nASmxajY94DviGjjKJL0tgaLU0dGtDfy
xfXarQO6+oXXXt8QVvwkGAbwBnpl1Udv8fq4Ndj0L+lYAB99p3o7OfPWbQYQWIwD
d3YEZHHBj0qG+EdBMi26/iMEVk1fgL1SYJTpIEGJEd5lyUEHtJMIS+N0a6Dd81H5
Vx6FRxy+rnwhqi0eHmLhyH8nTqRuxFIYF7vXERCHsQE64Zv8Zyn3bPOO+YhJsQsG
OkG44MVUZbYpgAt+gnPtp/fe896zGn+ew6l3/6ZlAJpUyUsMCCBdDAHw4JYKgpJ6
6BTCfGCxCt69yP1Ai2vYhH13Dow5Wg9Q4CsbCu7NinLLSI9qPCOiVbYXVx5l2NjS
1oymQwisvj5aX2/zGUH6d65+RGouRIH0ufWxC7T525gpnJp82jHY/yNIHopn4DVO
gd5+mRvniczh80TXI+4nKPkth9DQ80HpwT8W/kUeC1seMDdmLNglJOsZwCpcNWcv
/U/8/f/WvzCfhcX6ICoIKQXww/ki+jMT5P1VWIktQFhpyV9RtoQq0TUmUOVfiaRO
woTolWMbb6/Uu+LBbfixNyPt9/RGpTnpfCReL8xcD2GPqhrS+b9vgVWVncIBqt0L
d4hHEOXn8iobpF7ySLNwwkLGz5UVpatuCDf6/JFUIPHnihH3l+z6yfBP7e9KoO2a
gB7qH6mXTbJYGw2Ct3Uuggggo97N3iOsjFxdV+WfM7pp4ilTLeHs5rBdW0sCryXz
6mtENbKqn70X5wTNLV2kWZbpH0By+oqdwoGWICs2MCYvrQAYKqJDUNVK0YWx98ms
gwFQnKeGJFVXlMnhiPZcHXlkjAdy7hFHlVsgyAFUBaucltGrKwfQs5j81O5jsmN5
rqzoU1/O8ih/j+s41ek9l3p34IkQ5U4OfSo0ecaArX79GMD+l/7+1O/B9AXhSYiD
IOmQjApJG+kg8QhuRqBVj4ajG3SFjP+5w4ZBAEs3PhwuKyengm8ljb3HSU4IX285
sz0F9CWrseD+TID5SYyoOxfZgJJJDGZ7GFj4DhQeDlUxWIK3uQ1Ys2U7zfsZ/ZjU
AXGZnRVaLygXj4OElPg28EE1oo4XAHifWxxZVsCNY7E6+pWtQFNDC+BQTFwgCycQ
EMt/0LVSb8oEHcLpcUcYPplHqeI1wumCiLlJbqg4PmeCcURl36OCHAwa2dqvi12o
94GjYe+cCedsPLdXJeh3qovno4B8wYnbPUrhxfO8s26dHJChNVNaf/+ZZQXURd+W
Bd3lZnWUV6TxojPDFrrxxOaCisY34tSgBRIdzaLIAZ93oO719t7hYRcRgO0oNrMw
iEfkTaSFqobb4OkuxBPayS1pq8AxDYegoMeFUhK0k7GCme76cDaDLzAavPw7SdIx
S1OC+AKbTtiyUw9sLYp6hyOFH1iKyWySnWrcgSjLuudF9lpA237VsxBTtWYhkCK+
tBifR4zix2fBq8tiX+UBAK4e3SS32fKYLtzY8ftEQHhlrzqwpybH4G4vgduOc7/1
Nphqoes/XL/XixkmZawKP+noNzDJcYTogndm/3JXs5hMG8wtt/Mzpv/u9no92X2U
eXIhsXOm+BfMoSX/uu89ooH5G2fb5qh54tbl1BtfRo04ZYUF/Q1GR+68liWJjjEq
CY30lOVkwvyZmseC1h4/pyvCbkB7QnPzM/1q8cY/tQ3idlZhJeTTfwo7k2MPFMO9
0xRnRqL1tgZ+9MCq+tRipvpb3rg4KhHIvK9uaN8I5t/MtjcQa7X7MMTKsPzJWD0C
j+mBz4xOeoVgGx5UiIxxrh8oWA9+iUEYzrpx1jQy9V3l+aIRXWXJo4txi739qB67
cQqArbemyii9aHVD6QJM0iPRu2Cjx37K0uikbI7rHeryU3eYn2w9sdOyEZaKXpYM
dNr3XJqbXTmByXGwKKAoFxJIJNxwioJDVHCvJxrZFtYHb/7OdQjSZYTWyJm0pD34
kbQWvNgvLwhDqFDerWfSNsMeWJMopds9N0FJBjnKM6/R9+dgqQ6H25Kx8wBLjJA9
G0xhqzekogpGdVM247l7rfQIexBRw+o/FoqOrCumC8J05Tfb0oBD5JPXPTe+Q60R
1J8mvEImh+W0eHxehNWCGVI84DCnqp8KkG3pWfehZn9N14qhY/HWfv3FwfulQaZE
Z1lZZ19FRD/Fa98BYx3n7SYoFTcKgfFDoCTIrRoCwdqH83ibiD13FsAr7SfpDXOB
cwuN2fj4Tg8lbgg/hrROXIQGJLKEhQenYoja2SkvyrtMiGJtgRWChcW9Ra53gk/r
auqyloj7R9kfxMzZKO362uDr52Jo3/Dbh1qs8FlemZcxYpVDIxCvNDTuu7gqBwaV
ZyIjB7GAv7cycr7eiB6jQpQHdVp+LJ3V+lFJXAWKJiB4h/HjKv9HOlJ3WlvOetCA
sirit6icx+8VX+AUtWNAhlou45olsXy9nmDQfdmCasdSwugDlFIPsRc5xOCrqLed
PSKk8CGNdSUT4iALQ8nMTl3Iu29C0Mvr0vQLga32PGHu71nSF3zeVopCVcdLOKjt
pqaf5DcAGMPiQUJSbMTgJalW6y0IgD3RNLE7w6eQMEcn0PPRei9Itd8Cq097EUgo
ckO/QoqX0BiouddX0WC/5OpheSDb6ARm2zIJlypwlOpzKggkzypR3RQVaSsFBeMu
i+zemoEycygPuBtlAjREaP/h3QffJOGMdIV0QYeCZH1zge/9V9+QVUO3Mv4HbWGr
amXDgOZo5gXmS0oTWucIOw5MLUpmZwgx5wTGH2sLRq9MKtFvD+sEV2a3qXnYjNQN
Np0vJURcIPJf141XVb7pHYUwxzrsszn899XG6JzI8sFri7fOB0uPjucd3rJL9NkM
HddyXtVZ74mM30CmFQLBGwKj0bWYy81zZChiKnWU7/+ygHKKVPnIr4v0T4upAV0p
HJPLb+OFeXXWSOFATeEDdMRNtslDAPIvGYROZB5hHA5+D7flNdd/4sqvrJfDX/6m
JIvUNXhQ6CmtytADyRFOsK5dk2TdoB5EQVsbMxKRr1wf/kK1SNz4iQYfw28ZSVxs
X8xOTmvcHJ3XAsDt5EryeHsuA1nGjjffxs4urV20zukiWFuwSAgoLO7/ANtdegvl
lOF2L0FlPL/XFrMRZftUOLRTopNIyxqbjlYM0L6OHFVuAOHXjpl3D7I2HEnivL9x
x8ofM73xGuTYoLHvcAH5jsUFK0biMrVihtFvZEmfdrV2zcUuOLlqibsW4UPYsXSY
uy6XunWMtSHRpXOggYaVpip0vRYWGF0ocDcNREGFXTXccgtMJDCQgg8pv+SqLonY
CEvarLaPb4j9XKmR45cVtIifULF2UMcXRai6WBNwkmdEH86FbQk8KMOd8zXvITpj
M3LCtcspYn6aQUbK3vtqU8g8mhUG2D/Tcg6ZX/Ag0MOqW7JhO9a+WMgoCHBUan/e
G+DjlaXxNZ/o8mIehHRmw84feSmy08Tm05IOOPMtm0mZd1oFFpHGbHEGUOWrkLZV
E90fZ1f2ZyKwikbva3dOVFf7+NE9iMeos/iKsGTddEfPuYMfGO9DDwqT2EHlMnNM
qd5/K7Cgiy04U7+1IQS5SA+ld6zkwcbFmNoIvwAAPPWOM0v+ibumwizl/rwqpLz4
OdI31+WaGniXU5RTTrXpyPJC3T5vpFNPJRdO/Fohvco9F0fA6uA6P8i7K5ZjxEA+
JDnblggqC4n7+tlAZ0dbttWjSTN0YoedPR1HfebeLvp6Vl6TW9jQVCLRSx23lJAg
2FvAyTIjwILnKWC9BXuEnDU6nvwyznmgH95d1HK2cqFPtaCaHeSAE5wX4Auhqicb
Tz8xFifDOnN1YBfPYYToa/simGOoshbi4eRGy2T6XQCFISHw8yc7/yzN37kDrKDR
bzVXRO2Ut2+dDpGUHVt3k3NXvsiwVx8d4peX1Tz8xfqI5AhZCGPIZ9VaB0L6rTKq
bpDXJbkKQkgxhAfjrFgooq97/TK5RWGA5j5St2w+pYaNQ0kxq70+bEHY66obyoav
2SWGBNDC4FSY75Z1ibqHGX45sc6947izEt7E/6LGXLg8apJnld7gU2bi3IuRIlzK
dihEY9CnTF+0ZdofYh6d3Zf72H9r/cwWB/BOm+g0gK7v91siewKiFnjmJK5tvxHN
/Kb94R+ElOR79nxRkmb/jeU5OrnB8WBUruUKsIHuuslJ0S7dIuOwThW5qEwvyt7t
kf1ldzZDnhTTYGJ9BwcI5xeiyveQz5Oa050nqRvmbuyQCk3mLdxRwsWhslMOGqu0
Z2/rigf3tbyxwSzwyk9R2e9EZIsVYh1YnN2ezTRLcR4KWeheqQxqQosU/fHrX47G
Vi1lZdrj0Qa4Tu2Z9kE5hak6SxvvqsAvj+hbLA4+Edth2l2sgHlJL2eEslndzUYi
fq1RRwnl/Te2nZxFCXVzEErk39r/VwX6ZXctymhtOWdsAZCtDK+3YScCMLG3ky4M
Rqa9XlMa3c8o5NKQi/Ipw+dg9Cb5cI4BsfdQ9Vt2gZRaMMseQEmDat2jCJYVQN+j
L0/D75EoPVcQJxAuagQ2KMLgD7x739/9HA3vBRmEoZpFOjFx8emkvTThoudGYU5r
qwC0pvnaYVmYgKrME0bS1XsbjLHstJi17+TFMcNNKHhU6DOrPuzCV0f5gdvS5CiI
+SABn2NmK/2woUL1Icc9PKISZzMm2Fwk8Jkwb7XaX5nVHtHw3ruQ7Ly3rhG8RME+
sFMD0yr8R0atfLintCr7DJCgVglZlhOAty86wO+dGiGtk1jNPe/JC9vCnDvoAGaB
qgjCoRLqfbSE32qvqlc1hGYLtiXqzi+WYow/kq4QoNV7CVwX5xaiO3/E3Tluz/f8
EnOJ/b6h5OlAJ8hereVPO3IJ+HRcyAWK0BDIn4P+BJr6Ip0g/jO8bCNyChMO5n61
goRD4/k4yfVai8zpkxhOjn2E0f10o2rrf7vXJw78Gum2OEMNGdLr5bRFpaxLbf8W
0J7U3fI/EFJKUWgAZp27zmPHMP3Fk8ZL2AKAl9uHeyi+b0+HabJlB9jeHHbBjtjx
RkyjkD/HVy7gkas2dY5q1em94kBLdq9Xq6FByXJ4lVDh8Ftmlsxzn/Z3RB/O0NFM
uV40Fx02IPKBxj/AUXPCo3qcrPwGqqgpqZ6T1KnrfvRcrJXKyatnorMFF3gSkRW/
F7cOoZAS/1+YV8dGECk3PlVg+KDFsiay6zPbsZmw1bLq5mnfg7CzZeeazvY88Sfa
tzd6vRSzTtz7LfpqzAi8wVOME1YA5y5AnvIUoCdHWlSZ3pr5Q/hg0X6GIx15mywH
gMMKXksrj7scOKxQ48Mw1Tftk55x2SpC9SetPQJg8l6PoAWu0n/eCt543vhHGvUV
bNFGJvjhOuJVpfgaOB5N+S3YEvQZJNYTUnyIkHH9lc4XakS6jjzxVbkeO/NFtpyk
uAWM/fFktAJHCEWErKGJCJzSTNKndJyXWw/DyAjWhAajaaTOgewoilp1OVc4tNlH
j8DL/1tw47xux88v4eDNclhK4OXE2PfG0ch8PqrqU47ynI4qygET2q06z0H4259Q
0vHIPUmGbyyMcBx/y0kVMTQvIi0AGSiUimANuVHWoiOCozK3DeI4qOA1gbNkWxiE
2xvsnHrzZNoIjFd5DYEb3ftqMrxcgri66McFmPuS0gaBP9ETaMngN7yleWx0QcNY
75znv4ET9Rm5FM1Wgo3owOZu86CESi823U5NuoQ0M3vRlSXyuogXC0k2e6xhrE52
u5L+pGuGcCfW05BJ/BD5mhFxAGHNSWOE7TVzxF+iQvvMkLQQ0fHIwPMQV3fqWFd8
QFjuuaAaVnJL3d67eqehVvZ+AaCHMsbtAH/x78DTVtl2cYGrixXRbf64a+je4DPs
igE8jqPvrzq+9ZGYbY3Hp6kbQIozhiVPMMWW5oJ7cq7NiDWEvcoFBR8PEXjLHEkZ
M8HJoF1jezPzILE/gnJkZ4hWSDqV8XYZ/Qhxb6sSZeoNqWbGreuc1C8rxHyB5MoE
eYQ7KHkSfWlmecoZlp9BdnbJqGXuRYUNMZhDK7t2N3T92kpTSmu/XbEZYXappbQ0
AbAERBAK8AE+uGvO1gP0ktblYAxAMKmd0Yz1UNr+N9TM39zww2ibTwIftBIS7/Od
uJ5nx/XYgGe4bBADe/j9fiMbHLW4DGeeaJ2x1frkuf2B4AMkWYwndoxOn4vMOSxI
73Klah2vpj5J9g8yKWAiZGA+hoiJQcswqgu5QOWOYJw9C6aZEXDfDykxVRVsWmL+
sFeWQRgPr/mc/9WvKobXJypKTd6pzdXmK3+4OY72IanOGDgSgypSD6K8OzK/h+ZD
WKOikSiqfPdA+w8wOfa75b682eGSCAFcf/NZB8HvJTIoPB6iUlY2pQyqbi3A9/JO
tXUSwOuh+Yo/YnRpMQ9qjK77ZOCqoIGzz2TK/X3w/gHqVFBPvZSfVjkGae8/HFFg
9vO0o3//BJHHk8EmJftz/lkB9fbO6rkrREH2BXpLtzjNcT6NIZzrgHmfA16Ulc/2
ActV6JGDRuHed76NImyQd0dosr7iB0qLOtjDx7l0aCo3BfBzTilYs6eTL79WLGng
AkvA39ZF39zmEjRaaaf3adAtfnGgPLWg24mCl5hDMK/sVOT9tgak0rp+DMjqnWBK
6lpLV3DNWnmzda33Ehzb+m6dxiBl9iEFvFLm4ty9nX86VTpBk2hNqVtVBX7H07T4
TsR43rqQ7dfQnwWXopyBNiO7qmjSfznRBG4yd8zoCcZXot5hwiH3scfcMp1yR/w3
yNi6ZSDTpeUbce9D/LSuSpVdsJmfcPCJin5y7HDgFuhFHYs6wXzwVXbrBCqXRe8B
Kj0mo1U2q/McGh0gJSRf7CQNw9xBOfwodVnFZGcpyGojdFSJh9ldK0VoNcgnAYDk
2XxcDU5r3lAaRbpaYD/MBjyN9trXAK/uBdi/IHopg7GljWAsNZXcAvwJBJgnU30h
QOZSIbSNa3nX+zV7zLo6cc4MtoQb1cufEHhHRvFommJL3D+lLTZ+ucZgJxztbvfX
y/v7sab9wT+r0bDqI+PGLlB4end0ZBIt5+JrydI3twasXH3q0FbydVIUBbZryqDd
9XyZRYfrRF7YaiEHTxbUxL6LVK+bWQ+icQuyAtm3nzJWieOCeWuhY0pENxRmMPDk
gH5YhdtvBzKOvFBhiiCC6OTmcOBZGWoMcKnJS1btyCgaAYnVUuV3U8HjVByhkPAz
pOs0FObFSSj63TuRx0Nc6i0SIKEIP+XEKSBO6C39ZZEYtwz1AdhS5yfULpksdfG+
8tW0PzOO/DE9DIyh2ox+oFm/UfABie+Fs/ireJSZtOGxzKXbvcqHTmjXRRuJREAV
C+JmLCBNHm8iFD6qve3DAyxA/wWND7CJALXZWJreaXqDxg55M4X44xV4orjslDWS
mTx/p0aeUEa730faP3ptHjrSCo1a60C2ZIQsC1F3fd4xn3PdlNgpcRGoG2dGhqfs
fzQ4fzrkZ0d6lM0/dKoORXAcOeObWfe25GJePqvAA9yhCIcpjN3NSeP/gmQysi0C
UJUTvoUY8WC+HvTXcWg/D+S6wg4OSRN+OwCNdQAnSaJtpACOtC59FpP2yIKqDL+j
QctN+U1GRt0MKedDJ0NnTacMnVONVmcvNLHmEGZ1ZqwRT4nrF7Pr9HKTzIpHT6eV
nLFSF7w+f2Bu7tHv0bULUzPQvv7cW3/yPxURg2C5J8dNiKlhgWI/eVqo8Mr/DF7P
eY1hZI4ntHqj2D+Z8TPMnOMLReIMlQH8OT6kSgS0evufim0AjE5jP0WXJPd5gl9x
fzuADz4yEgrpFMRuoS/JyI0Ou6XNvPtQ/3BDHFZwI78caXkx2k92OshPm+sGRi22
PCau/9Rz1Qf4EedJZ3hMhl4/LVGLYYiP7MMebt3/GeVMaN75L5D2HwwWJC9ha6Fi
xWPlY5tZk3gOC7Dtm0cFIt47lRwI6rXSOjQ0xvKD9ue/g5othmC50Glls1baKzUs
tCE/LOXlc058eyae6aobieNxSMuVvvQHznBkTblLIbJLKDj5upwuEY2xm7bx8Psw
h01NDEaKIk9UFXVRt42ZprxEaeOaOSPvXvMz43A2VouMPLnOkJIDbGzY4iuu+B/T
K/ACfzVlY5FYAmlhv82xdvueRqXvIFnc1lz2A+vtZtrfF8Tt/0MPImT1m5wyvR9s
150semv06uOsHOIAMf2Ggc8fofOIDwPuNgXOQi7bSpGRxdAHmnooGS87p8dB+OsD
QmFfKXk6oM3eAnT+HFX0BE2BOwlFtnuKlCphkRXcJxJ+nh2BpaEFGUl7NqXw+1MC
XkX3bcXYHcWW1RdbNMTDglyfEh5AliJVT6LrWzGcJiBKuiJrvh2dzz00b3G/hTpd
9w/cH0DylVGvkCJ+bDEUjR42Df2U1V2pohSABtKz5jQWOa1PtdUWUWtR0LBOfjCh
+wo6KfIR7UnuvV8oPwN3e64cRcQqAjWIkRpG7450XAzH6dfjfGSjMwdbVqtRwxjQ
UdCtYtMV5fHHP4ZvPEjK2+CFo9Yf5FE3/pyKD9/x5piwNyvGS4ThBvZ9s8V56MqF
eNgeUJuF0aHUIXnO2LQPX+bPiX5JhuUfw5Zvl0h4jCNcKiTWzDect17+plEHNHRc
9lzwGM+/2JER9IE8/uESQlEFVAFEolmhpdGSn3Hg3DRLjfuYXDQTU6Rc7eiaOy6s
KZS3ocCFSLwwuNs8rmhwAa2sTwiUnibTQys66tlaTTy1AmuaVAIzwmV6xRdDL/Nn
DjuSU5d2yCaNQvCzmYbxZTec83MDYdZpipOir7XaA+j1d/tGoKLsjczCQSnQ8qXd
pxp9DlzDWRTv/GC8LHdlT2SVSa8yfu1RNAllWMmOWjvfzT+zHxsS6s9XKWGKduaC
NfokYHJQf2166Z7/f2oiy4lbEehBQUqk6J593+mEmcLFcrXuNtPKEVXLBrO0dZN2
brSnbUReAuLJrURZK+wslPbV9Y7Ge62kz9sUMH7SIUGfxfV50K3dOt68c74Ohufq
65AxBd4LrjKm5/Wk8Jl5yFYxD5RkPWaaKAzfDDYKozPeJCDPlpzi9kZs4zOFydWd
AjV/h/V2ymO+kDDrorHi7kf228K++KLdMvfogQtGFcFDJGXUYIMXZSWs7G4s42P4
V4iuDR7AQ/YP/pi7TmCfVvkqki1RiKolwC1hrwSPTzvpt/bwhE63NbRD2WyCiqMr
GufB65SG280g4KoEdnVzLGnbc4MbouZbp6MXLbYlA1r6pMj1KJ2ijFNdhWCfO54G
7v47uOmnccrvEmJ5OV/i90NGWgrUs+awFBm3MroYEVpICA7CAQL6BouECPPUjOme
v45sIFhAyfuSLyY5yZkHvtQg6hA7BuLytSofdilAtifnL1W7E454xi1D8uw/2ntX
vdQwHXEWKfyaAncftvq3WExaH7FSbzxZgdLSLK3D3eQfPAeNp4GBEOxAYoiMHJE6
S2cz28bVNrLnjqLOHnXlt8qZc1qBH6MyHjq4j6fTaeEzdf+ATgdoPg58sH1WA/vY
tvyZz5BAsCAenilMdHZd+EsXGHSJm83zBEndyuUidWlF4Kv9Qhwe2RdIuxpNLwgX
klZokCEDGoXhUSQLwsqVh8Vv/lf5tbE0igRWMbJsV2i/wQ1La3nGg42suDT9UTCn
Sfj+3QGFxDqBBAoYaqYChzt3xbLTmXjasZeT3pw7rHUlDqCpCV8dM7Y9AW5LBXR1
YPMBfO/KdBbsMG72WEuYEHy952D27ylVLshUrHLtgHtG21eoUhZvmMdabwnHbkpd
n1/3hgLvSIGdqWAa+qEcYrxH61ZuJcYz4jKLq1NtmzuczTzTENPDGV717KUod+Hj
PqzTXbwbkU2eE9NKbw4oVMyKb+FZBnmnVdvZzK+A5+9cbtPO+xDD29fW8iWJNdNM
xG4+SAuw1sNSab7hjZRH6/eVbAhNypepLq63uYQqXqBcTrl1HlgdeDekWeorV3sI
QqvO4Ri5CnrWXhCa5epW7gQCSCEfUs8HmJRRdyF1B5wKdYWpiq7OYCkZmOMSAWn8
DfprSD1i9xzJZ4HuzyDkqdHTj3mNetOhWDg7OTg1zXMzWM6Y8bOraHMtc4jbVi9G
K+ldzq3s54Ng+LoRE/9i8J0L6nKgA3lnyaUY9PWlmxh/ySb3B7THwjGVxytSJ11E
4CA4vqs9bsDcR2LEjge2b/Gr3FYQZRHcFpxad0/REXP8DfYRl/WGm1oXkyd+qwb9
gFe0FPpczo6TszFoFB6ki1CjB8NkRFNkrwiXcOhuH6CMpXjStb0xKxy2ecUNWNlq
KGFvjhDfcQaANr47s1VX2xluB6ZDiAKi/p2IbcfOEEFf7woisT3FbFCUCi169uRz
uTk564rbQMszyWOB05d3QkRGzZo2zG198vDzoEKJZvRjKatN3zOPc4hwxhy87tBd
BvCF/oY3/iFHXM6Q7QP5Ox3xnjwBGen1MaOcxZVfK7nsRlfz7VxiGfOQm2Zg/50a
hzHJlkKv6dKpM8DIMYSQTZoUE6uTz+1WKR+O67ZLSKpwupohFq6xJqZZOV3dEQp/
kgNJZKU0qQVsHwhiEEzU5YGu1k6E7AcV6Xr8P7+yf6C9vQCvNtQ8YJlGFOsOTTzk
bu30Xt8yd8RvETzxnaq2IsEwYpWG2bUefJ5e3V8CIgTZpKK9Aag2HHhmm4ese1gM
QQhte2z1v+nvf4QgQ20PNv+ifv9A6nA0tV2XPVcegOMCuDTAoAzJBaJjJQRlFhy6
h748QYu90gKKZckDMQ5+xl4k22Qh/S+7OxlOZRoXKVRW3d6FZvxJu4el7AoQNXUm
rpQoqUQf4P3MRHThTNHfB+Ch+vELcdX6nZUNsrsTRaDDzhmhYpd6+Zh5Mn5h8XL7
NNGruJUmNyoc1CgSO7svNgHbaECP3O46GT0I3/pNI37gBB5lMzho08GPiOT5oiGa
LH0Ul1+aB4zSj5GX99I8CdidGhaq0Dhi/kS4HwOR6K0l5/xn4ld4PS6QUaK1y9sZ
aCpn39XOkPbVLhsMoRwTMxwjMWIOK7cU9mWy1eVEX7vBhOjwICzzztb2uPFGK4ji
KyzXRfkufzmpfXsi0GGiP+y3KfYx+rxqSms7Rb8eQhg/VJQpQjfETadpYCQuutRB
CNsPmj10EloLVlNUngP9itaGBSqg3tTFcXsN2BBvRFb1P3r7EKdjQVJ4aGbkY95G
5C3sw1l9GHUFdCYBa0DNHrQJgAyxJblBLTj0n23Er/S5FaLjb08cbFk9lYJvXAni
LWrhQdIhJ3QatnG3UKmzZo+0YJZtNRHCoIz72uOUEgrKqFFh3WtuVik/3vA/Kn1j
YIQYUwRuNs0osS7YQYYNiTNDmiBsl4jm1fWULIRNdbC0HSWUdde9loMhlnxV2sOb
b26SqdDC1NF81+N48S9lejb1S9a0FPKDGJUPanrZF39wtTNPb1+6bXlLFbpKpGQn
LsTmi3AYOYGGGqcUkPZfbralaNvWwZ3Lh5rDPNKtd5rzUmzx7GR6/yJI/Dqo5oXb
lbkus7bvJK9SzU0k/MTDBiVykUGanKYFv/VtHLwrRwJE+KIMtCgHeaMyaRb2shpR
mr7TAcswjV8HRPKS/M0poxXUUVPBIYfiS2yyU6Psc76eb07EFTl0CP3GfnxbR/cM
zxJdPcMcU/AZUChjiuFs8ZiDZ6DYVNSyzVAOBy0v+p7XMxYMn2bxzHaYPpwRVw0S
dSCXr8l/dgoLChYH8p0BmytEqBcc1SSieiMe9yth4DbQTv1Jn66BGG7tvholoF3f
0WzTwuTXN5Pnza/3Ivi91GBJvQ/XvYLrSAgcSC3vXmEZEZP999rRdpTVxf9NMQ4m
n5csNSotcGL/x/2ae7RAT6fgiCU9mWOswFsLDANRkEcV78BjDRWFbEiMggze5GU0
ytlCiyB0kt/PPV2khvv9yzuA9L5aKnvhGo1o0TkRJOW+z0ya7ONvsoekso9Hm7AN
K8f3alk9c1oq+ZwA0ckE8FLW8mYgeDTxxmAn3fF2kL6spuIq+O2TNij6aVdRrjKv
atm4/0bpPU42VKAE2O9w0DEr56+xTa89FxlcGRBigWx6hpXfS2yl3t/rzTRcuLIv
N0txcQly2En8mn8tCIsS/P5w4upBOzjYBpRXl5misy8w3tT0N33Y513xHH9BOIYe
dLJThF3p+JjepCp45iA9i89/dSCHadPRwEddGRCw2hK10KhGIY9r5DXHY6fidw/W
L55lRRQ7jhyDZAAI+mawMcGWui5pKKdecxeTulHYT4D4dAL9bk4wS2GiWHf7j9O4
MS3+27PA8Yi4JOZu7FRn+x6N3h1iARqHhGpUhaBY7P3wbD1598HSHcg3TTEJ7+Uk
RVfZpS2C6ILX7+KZ+Ui6j2i/BK/brmj9gc6ipYTUAjOMFSk+oo8WQpTDbYse8V98
lZNnSKnc9tV0pbzNwLAm244bkiBDEfsSsjFe0fI/dueKWmMt28UX646JvdtXsSpg
P8HF9RyxvNjhqngGg4mll7GG1W2xOtHc3j8i4CPb4uUTqoN+HEUnjhuSPrEKurT6
m8lFgyYTPfoNgBS66hfXqr5+s0oUto5CT7MprU/BC+ETzZpIp6vqTrxWd4QnnWua
wn+gQ66FwlQ2t/Bph6QXmhzc4OYJD9ix3bT2LU3Hi83UXJMuUGcn/RfslnX4JNH+
BeEsbtvR3L1XAjgMhaDVk6AUBIeeoGeb4RQ2pKqNlSGG1F5T9NaqR8aZD2VFwx48
bVOZc6nq03GHdfEoYz3cvjMVTL/R4qOvlqDtHKIB/JonNjLQQESi9Mzd0DQy9/Ww
cZdsxqimWgED5vZiCDhEyBoHn6UFFh2xXpTvMLQ7rIB2RVX1Y0NVmlPe8K3iAAwP
rSsNxKHKUDnRkVLMbAiZ7rno6ss3awhuXuJGxunjt5OP4SsLUTrGGW/ir1yQyfEs
kTdTupvazU2dJbvar3dV4f6i3G+OaXVy7mjWOAW7cMfqO6JkmGmbUagPoUi7sL2K
Awz4jfBFCXZ/JbPPNTEzn7ZDMjv74satyMmb6m0UFv0J6AWyoEmxLN/gBJHb4A0u
pDmgJGpFqK2vkSI07iZJlv4R2ZoBJGxRoM0iRHwjopxQgqPWsGs9Ul1ZyCdIlUpn
aAV3LjkVOE6E6d1N8Z6QgzUuv2GUitXWzaNgh7lD78yK7jXyp4QCCTBrchMXbfh6
zUDnReLnv7PexwRDxc9Vt6HXMFET30SzP7jv4lmQ5Q/OupZg7gDbawvhz1h4AmWi
3jUVCpQ206kQmb9+TisxRzF26Hz88QxuqMD/qIPJL1PCVD11fV+F+lUUimhUOh/a
R8P5OCyVGrW1uY8t5O4XVArSpNerfN/BVfuZaVWUqFUUwRjtqadPbjByJNJsl1xb
LjyoephJx/fbbtJfUQNt0/Qq3wFrjA6SW1TL0yNoSwtXs2Yk84SGSCyLCdYoKTHv
Bv7pszChA+L/jeuCbQLXWSK62jCtKJMA+Dr7k1cS/t5bxgRPJ3uPeR6H/BLw2GNP
x8gfPfQ4/Bn5GoB/GdaMJuRKK8EVfZYpa2IW2t2WjJEKN8TvAN0HRImVXtqx3f5l
YH0nz5TLiXEamcVHkt+M0lhZF6EzSm+JEYFLgvl5yAZXyg89UBlriNVh81qFN6pI
IznAWTh5dCVWxeldYpdUd9dZf78QeSCJdqjkmeEZjOt499h3q9BH7+tyi0naQvtz
eA4ELMa9U0wtnWbh9knlflBfE5kvjRS3LLdY9IMHq1ZWgfIGGwXqUp4FTnWE7oqJ
r/CNwDOMqlZt7RKDWmMW1rI8cPuQTaGNKXJwzqIfzD42E1qaa9C2ntpk+rXDiGfE
vpRXRxFLM7XVTk+8QhhnhE8NGdmclgGMKSGDF0fPc8/s+Xvd/lULD2umMc9QJLaS
zrgGEo+iWpRt0iWzS9MwdQeF+btDQVhPcarrdWxfTRRILOLnvGmQx0DhwD4qPIYV
hy/uSn5ZwvCr/rchmROzY+Yn1yMsbWMRqSqr4D/mwRqsb+tYCOpGrC8Baidsv5Lx
kzmKcmx57HtRsAoB9+fpIfGsNAp70rUrtP8V2DJyGoJFEfXHX07xCdInlSbfedz6
XVUdGtHr5QvPWPgOjJuKvKuV96Cox4j6EJMJKhX+t/ho6zvwINfe2npp5sN0Hwy/
y2E/oLTzgpH6YEGUDljIkSEmATdnjJAZdKipfMtEGGI+efvMsIyf0NicmafBq8W8
hmMmPe4c9XOh/TXURJjDWrZLK4murayuHftiMMo+P2A5qIeG02+byY/PCqKBSLEN
vVo3rGrAluBHtvsm3fg5Kg/1bFjiGWU8KZNG3PSuaz2qUdCCVQNdCSwOh0HD8KlL
pnDjmoZEiyJFBCBX1CjlsMA75L1c0geCgI1WM8CXgSGcQcgH6rVohFymGPxMJZrl
PYmb0ZJwWY10L591Hm4B3UuKUT25jo6PRpThmGNyhym8qsRIG0waZBmfNyTgW3zE
s0bUsae2PntHZsA3IYEYF54C4E4UNcfVP6TaAU0bmAB2Gm28QD4igQBz41mV9M8A
wff8LWtUo9fGVY7KkbIx9N8MedkCnIRPzV5OUWDlI0Oo8qO49ZreOudjC7wWvcKH
tJWHNJtoKY+GRMG1BigKZThk5RuhFjgUzvK+EFzVZkKfQSzYl8f2WT9QxVu9hSGJ
3cISgAvMRRbosA8Qi5pqxIkcTtaZEjHoy9Kxqonsi/tnfaYHBpAybe3gKPxa09ad
j+M6MUVRpa5XJaLNC0nCKSzUaKml7laFsyccx/XtIhtO7Lt2YDUKcNj5ra4ikS34
IvWZqH0vsueDI7sGGXBN1FaHIUWUYlLmqdCvHIP63xnbV3VKBPKOeSnJuh6hduI5
988BpN+EHnEDi1XZQzbEBPBRXwZuUyEFeNwv8sfhcdj/9r+nI7FrsIUiL91lkd3R
2EIZE8UNZQRWjFo3rA5cYuAtiTJll1ioGKHKA9JIucGjjI87CXuMaFjJx1Nxro+F
qvjcUKQLOBIsFx/ee3YC99NpbNrkWb2K/1Qza3eskFHourwEqRtF/eYAG4x5slsJ
fo0C8p6KcUkp4sSAaVoWPjrbm2hKUQz2YoclYKAj1BsOm3exKVzoyiZJpx70LCdn
rGcHYYfMD5nDQAMEKe4u4xhghnAYW4ZsGXvRXSX3kejLHZcphDCoyOseCEAMhzdV
BKod6w5jbYSreFccKCoQNDz9NbysUHCKhCoxxaJKMB8CwuVhJTL2gZm6ZtcF7oJY
eWVi6l5JpOl5w5ezE54arbs82o46S/8oRPCW4UeFxeFPH9c9+FDwnS6GsDaIAhkJ
ARs652RxbeHgtqu8zRnwB5TqzFgpLukYYo4gAl0q0pgV82dE2VkA6VkDEFlbgeDg
Q5bUwhQ9DnIHjDzzQwRzM64rP0XRZitvZFG9zH1PEZNUM9dVKCoDhjUHpDOGjhtr
/AlUKMTLT2+Xj9xr6+V4UHiEgnxLT+nO4XVfrqIBf6Dk3GW34i9jT9gE6l8Llm9m
lz7ivlPh1/EZ8Z+U9KjsXIHXqC97ctg7gTdg71K+2/f8tTzlVeXuxLwWslqEaxO+
hEkNLzFY6ufzRaLqE8Kx8AZgk7vO08nm36wBy/60w4uk2vL9RuuL0YzYqYf2+srg
JDW/NoQFgCSY28+d0S+s/HMqZIKAQ7E3EcK1Tp0Dd8g0MoEYBlaprICdVk++B6+k
EB6fO9rQmoldDxXioxDopcY4F7WcrFKyxYpuJv5Mr9CWhX4/wK2bYCr+pP7CqYpF
yfpXQw6tI1296SbVMMje8V+4eUJ9AOc+U7eXqagHQ1mxsoBoR7l3w7KrlQtaDRB6
yX9F/vNAbW9rdBGt/gmwc83imyTkaWVx24ZQJWqxCKQBfkJPM+Qt4szLOTI30P5y
iR3miG6WH/kNkzcLej3Bgf2fHO/3aBahw6KM4s7KhX8AkUPTRlqsYAALDzmKYkur
81nS+D+3ZeVXILqJV4+pgyiJoDi7n4GZFr9T31EgNOJYpp3L7acwCWQaV2vr0H8G
DOKJUNLNxnifwFCCx4rgcOXZx3ubbyJfgUEawotS+1xWDoG49Xdr4N/kN3usK07s
5Vgz+13odVwNdV8rnrR6osYBnTjkmeduzgWq6rOiH4UQHBgV/IzVI4mEsrBnFD44
kLpReJ2fnR43/zxDWWydYGjMx70UznbUjaoaUq9HRwsYWxDWfHLWqgxKDfU9ByfQ
WGZgIq+fCU3QNvulJNJD6oFd75pecgaqfSja8zTwR09HBV+GCQLIjRZochI+c7Vp
svuk1fpw1YSNVMOXh7gCj3vSAV9UG0WxRKodR9jTwLuQ7I9zsC4Glwe4zEuiBNUd
M4gjzJXg4avkKVSsAwQ5+EcDq/Nrb3CzRqAcrH/hshHURpWYGN4GIq9Jr+Buqj0K
Wk8r1110Z3ik1+sQaxOZ9WcYDkGrl6LQ1/Ia8BYve8ze5fLzUonvd1os2P6TpnSi
C0buPmsBwhWow2cgwf3nFzwGgYnS81p43bbbzcoqvwn1lrh5ZKCDdNTtYJHHdzEX
wHQP9eIQtcpBBILIRubdK5pB5NC4ufSbYgTDO7kd/OlZpJxjqvdZL7Cnpb/omaeY
aAMZkp+ldEaU5C/pY5+njjv6W5tTuyk1fVTb6ZZVMLbqakFuPAoQVPlOMjzYu4rj
D5MVU4eZGOXta1XWmeLAGJ89BZeFhStSUy/DlEeBBgaEWcKdAhq9C96BJ/3A0k6F
C5NdZ+EceZcyjBPLVcN7nHFu0zYmh0Jkp5qvJTXANbmxl993mcnv3ZLrIQoKOaAI
1ITXMzyHBxrDhgop3wCh2lhPgFTFn2Jwjqegk9ZiOsX1PpW7JF45Z4avi63LF9sq
ouUvqLKZuJZ7ZeUoDGVMTxMRJ+reb5s/w9jzPh+VEaPKDQo5u/bHkdETWJ1Zhrhs
u8DVEms3l0xa5Ecr+bAa8xjgsRLWz194R/1PxOpjsrI8VS0uc9ogqCAUCZrY7zeD
1vABIBkofj/O/Ev6UyCiqh2kLoepVWhoG6LpaKQpfdgzWd4agNpB/erqCOuft2KG
jqjBSrvsMwuNKml/rEw8cOQBdEMrkAQHVSqMog2AFplVfO/yTCEvElvFCu1I1jg2
kGM/jYFHBIltHpKPQHxr/OtxkhZaDypssziCuaHTyzz8oB+zJnTU8R1EgyPem0/J
rskqvAspSuz0Nqk6Z4FD/7Z/A1madkUKrRONyQfuA0NhxWUNzHQH3eYvqIbR22C9
RGp9xxMpOOq7/DkZszVuITQ6aFexx72cvp7Ytk6vJiE3JJl+xCRYNCn42rWSyp9q
kFKhHdKvyAPPC/Ox9YvuuLZht5gaa1rcDILP6G0A+8PcVsLd5U/EEqfrc6h/eRIU
MYlr0VNElHt07OMYgAV6h8milBzcXQW17dQJttA/LzGCXrK9eXE0qIe4+8ld1vtO
n5o57v5t9aeiTvzuHfVhgyRxMwixIpcDuluZsHvjCnhzuNfwfrPmPk5HLEVuszvs
jM17/yJETyIArNaAK6Fxi1UeShhzcm4j/2seJk90AVnkmL/ITO7lo0d5CG4cdmjs
/a6WL9tGmjfSFayYN1i1rGYOjiz0hR/IBH7Hrs0ZSFkb7sIzWZhZqmzsuZpyv8kZ
zs5C/MbTmrUzXecfVgjlBm8l9mTS1gmGc/szzKqdlCI9T3/rk7QsDZ7sKIDEBrAO
qxa6c1PfkNMc1AjBgGnGbhsCb6nUfBonxnHwYgYVRXRjdg9mkhrJjbwggySLZQ04
PMEBwf1NvC87hXaqs/i8wugYkUSDoz0q4yCeS2P12Ti7/1TLps9fQUMQl+5anaxX
+1yzjovqcje8h6L8T5HnaD9tuKRPtv56auJnFXffsybh3fxpKiobqUcf3yiZOSWi
KUHzQyoc/81RyU7tTgUalLf6co8x9yFkqWvBDtiA9Wm9TvdVgVnw6wUkdgrIhPVo
mH8HJE4FWqgnoHQ7xkJi99XnXs37gQ3syylz9PkXggLoEHeIpxndRU41cAMx5Fun
CfjHrCRVgrwmqM1Aa1bQxBWY53uhK0NxE+1zcxlVI/QCAvGd9j7pZ710lXIhSDTj
+Qj48ABfC+27fugQ1iOjJRmSwR/hpP4awDvacpkFmgyKPTt4s1MBug7LAfoITbsU
vFYfK16N0Oii62gMbyPaMRcEaOxXcfj2e0gzwKHv5+FSAmUWwF/bSY4x+f9GwYsM
/8mcd+G9977EQXWZ6g3OrNDvM8+dcW8Xgbp3B2jEzvPibZGQD3NKaH74C/xNjmmc
oV/Q2kBiNqvxfRBevDavMWxPChpM5/8m7LLRx6gUpQIB5DUhj3cRgfs9UR7W01ZO
arZ7D1EiL37xsm0tnMBhIXXdfT1+TqGzTms9KAgoJXrCqRCs+IYCUU1tTxcBeQLZ
C1rZyCmyPj7XlWDc6dtTTMxACC6CdKjO72mRzjn2LQ+/p6iVn9w6XVFCHXYVIM5s
VxnxLogDp6G2hGNWTmRbjCqe6pXFFa71oKim6M4JRLMbLTHvLpxwcGh+fjTyGCD2
K+VtoP3N/vG7FD3oFaZrUwgRslJk6uKq7fl7moIn9qvRI28jiIvaVft58GJ6Siq5
bE63g0b1EiEbKYIy5rgtocxy10SZ30Bmr/7sLpXK+FoQKFlM4rwL7j+9HPUyMKjN
jGO/Tinjf28k/+hnNRzlaql0+7ZS/9ZdeQtCadgbfFZLieybDxPw4RiAsNcV+34N
Yle3+EdX8v/0mB6rem+N557wrHeEMMAyZLyq5FKZcBbZ59FKQ9F7TRkjcrB1z849
lxxc4o06DwTgAOZDLW6RMiWEooNODTwu+wH8uj4kUqOMEzwmMygEmw3eXnxD0Omy
qmzx5eht9rd/5aQhFMxwthtnjM0ohk31uWLnBZ0CeqHY1NeTcj9fBh3ABBMUGvkJ
68rO31+yc/eH7D4+5qRlyDUSuPTap4BR3i3cP7/Ka3YGJriN4SCvi5SPQozVg6Ij
hQVtRdnAJi8ja5AQC3Lw7nD8+RTXFGikzGweRzLB8EHYOYIlgWUMsIQNi6X9/G/r
dZoVCdLWp/Fzlv0XORDRYa0TChu0JxQ1fK+s6ftEX5QHTBkzCWFjH8R+LdBt7EaA
KOp9KdJJJpSXZvQvN+oXIgzLzLNdERdW0tRvGr918AowTBHABh+P/xE4l1l1+3uq
pVI8I89p160MyVWwZtJnTJ68T2UB3aWF28vVDSswmjafyd+oxwCmtZj1s4rFJadN
G0MDs0HWy+PGx7Lyodq0m5lg0w8QDflwMYMdTFkm3HLdNWUdETKwuPcc/H2DEyJa
C6pTW7rhNLXRliNgH7XPHB981gbwmLjHvvIg0Z+piVTGHDxHWyhvNuQstBBwstOz
7i9k2suN1VHwmTOjpM0nXYww501mCPPdlTgPGTqte13usfPalYHO9pTLpZHSYWRr
vek1GJbX/1b5u0hzvkPcyqary0OYqEtOCYkq2R5b3tEiKiJpDdTlxYNUTRGd5HnN
URVzhdCQvTGnReNfEkyNQb7NWVrPKWIoQq31MBQEvk7Dcj9B6GTkPV40SrRSbOwq
HR/A2GSrQ6YfQLKdrMdUCfolHBRoGrjsKfd2fxojQs4naJ92bskwtfn8l496vq7J
ITWwx2nC7hAdhetXl3i5D9dfPNWyHegxDnSP47tbDmy9Ms28evA3tbp3yY8D9Lik
vWb8QykILJP9qME5+SAOEdUNMcRxhmPhQ0FYnbuxQOXjBqV0FxwYJsK+bMI6r2F9
cFmqT+zkDQTYchGxgyGUhFcIKDKbyUfYV7+Rs4IjB1WMVtnog1xIMQqvnmZ/t5qy
B2xK4zMaNtoNdhn8fvSpkszIFGNcbrzu5VOITh5xZ0sjshgZsLmhj51ssBUzAiKU
bSl/XDHsIiDq7NZ5Z7PfMZRzri3QXW8kIgXinWlfTmBx/3EbZcZchREOEfgJsD+p
SKlJ2J5T55IxRpnKMOzEIpq1yJwd4+GX14Ecfis72Q8bypHPm2JACgzcwStouoyT
XvBlLK310ZHbCrP3B16rA8IUsF//Knadm4n4bwyBJu0XyRS1CSTBx/vtD86fhOUn
4+FNiITaCR2S4D5PK3xn8twpKroThWgwvBeA3GlWulpHAxBNUp+tu3uDbvWG35+O
Sdm2Bnw0Ugk+ZYxSc8mYhIqji87Z9XTCLwtXS5b4Gkovql9JOK4BitZunXwDmGAr
idC3vly+De5alkFB3/eoKG1hifti2H61NFkovgI5YplhTkQ4+ApU1xMG3r+7y4iC
/lIKLcAssvp8WV+H9Ue/nPrsVRCFcYi8oAW78K3S/PxfACZ05ym246iAo0XC2EHe
4J8d6LEkSDyQSFiyuxGGl3w4CjOD+ZHMeqZ6Wlf2VdmlODaej2pkyw5nH5ExXirl
ohs2JVBz2WSJVYuY36k+GgfgWTffk3iiCnrqLU0mQNAtDS+ZSdKykdwjPtTqoyPS
wUKdSyK1S9ntYnt0B9zJo5KensLPKPeq9ZP3gsMmFWcmBgYCydXP3LhofogmRYxI
jmSZxGV0HqhU2oR5SybpOcWVO+EvXXJQ/LDb8rRYxCEv+3YcByHfXlFZDUy2qxJq
HJ6BOumaHrP2l+TdEtDXheJ/vhc6B1Nap+yxQdpUXM+g+NDKrzLvxYgXNktfIat4
LZ+sRRTcsmBQn55WVoHoRE+qEJw1jbBkcnA+aM1mwbo1nSfHXh++v4aOreDCiCak
HBHkh9Fcyq2h2tV0zm3noJMpjdDWBhwtubQzTpcPpUQEZYPQOI6rPP5laNZn8J1Z
Xydd4IAuhp5ae49RBvLSkFk63RFeJZCM7ATaqqyianQ3rYqBY+oV9O151cTMqJcW
2krVm9e5HS92MAuRHGAVZTitIdfKRU7CI2V4PttuQBrd/rloez2WbSQYWRUiG+L+
WIe6Av7bVG+TOkQsi1v/9297PZWMx3wZCeP8+xo2Junyarcb5aESbVuUzvTyMkct
AybEa9Zgh13Lm4fBOnXip5nevFuTPFyOA7n9lgCsjpZ1K2muinTiUWof/zHi9FwS
wiXc8tIyFkPyzddLwVGsuNkVdZUAM7b5SRDJtbwUKzk/eHMiXO4Y0QNvY5PFsi0U
FHXQxgRFk33Nc+cCU+JuZwFToBKnUxGz6AQaq6w4hTeJUGaEZ9UTDHp1y04ptnkh
r5MPjK9SfnpU3t+mfEy5z1Vcq/nkIuQxrIP59QED3JoOxysMViEm+6U7m/pK8djz
guEr8f00IdtHGGADP845hiTe+UrX2zYr97Rag08zw6La1kFQ23CSysfNTTEj+qpv
bOtt85rdc8egAGgfDOGTMdZZY6lsQKRf6hzenIf+Sfx0wpnkYD5AoBzyPTi1u2D+
UHcdmHY/calr3Jz+MEpW85FcV0r+F44Ofi5qWQgh8jHLjoNhIhShfH01jCnZH1mw
gOzmqzbbVwtYt1nufTAT3iSksexJKTC9ihIlm/H9coVMK8riNMitnoCma6Z+MoQH
g4tT3CCYDeBU8rIC4QGGiNbxmoZZGa9sTqFDS8hVUMPdXxDsTCKUC9tPstJNtBsk
l9xADmVRRU71X0zJ8bOKVx3uEaywfhWubVPPxdFBUHk3I5YhDmtZ9wtaupDSQlfu
6debrbv9nPGuqGNhxZlYx0B2F5hIT4nd4AcVzGuzTc3zqpwtUIXMI8I2YcTlZWu2
LTLFHfAaGGEPS0Qui8Vww9DMbUJrDxNYS1QVjVR+p+KZJOa6eNLr4ZuweDjjYEic
b6AhdMslHkDFchlI9YnLmK/gecEWO9/vlAfSXNP8HRq1KJWvXHUujw8gAJWnoLTt
rDp4CSLJbNPjN/yVzBTJjnYNsDDeoMkAyjjVVRRt8s/Cy3/Pc1lS4vxyJ3hmc5j3
UtNISxryXoL6ce+4XC73QoXaze0rIH53cV9qb7hf15Np31ZpovCtacSbx1H21sK6
5h91X6hYjxmgDVVEDqoCDk/Bkcp0TI0uw9eRKV1Y1rzBmzUvOjzOpWiM4NzgVISA
tUnYZpHxqncmijciajvQXRCaT+vvrjHXuF5V4dTdnrXyQqdhk8Qj7sbLXRW4/G1C
jVbl/rbuFS85+IUg/7twitEFv5k1BtAhmEeSa+WgPeJ/1g/LoAyzvsGHzYKtMZrc
S02OV6aFF4xSWiEPT6IvxIC8RK9sGBqiE8dvwPv2tgCMv0EKmqtjFBe+kzm4cC1h
tk4dblhO/byguYx46GaLt81iial4PTbQiVp0W+SGodByLAvJDRnxp3nRzWmQ5ZB5
nwvPYE1z3U3unf3Rq+sCZ6K79BidZCD8d1y0IrMgYc+FUxGZcux/ZQyhpnNDNCgS
uV07lNcw5BLvsemGGoNVv9tLT9kf/EbY9nt5SVO7ImAYp0/yNSo8JJEnPG3TTK7T
wc7RqN2LBZiTEmxZ3A2JvwnWwT0OgQIpltFnkfga7DpbGQX3n7Fo5KfI/k4DjbPp
S4Ey3FEcBMBWiAyqUwTw42hTS3RzqWKNZN4oPwUNaa8v/b2nZZuBH8ATXzYkZYm7
4RrJdN8z8NLeK3t8VIiYI9snN3eWgm1IoQN5e8kNy2USzHy4T+nV/M9M0m/6Ir8D
seDwobsuz1gsv1x3eZMtLBnrYlyJtPhgxUVT2sKyyN6tPGesqGMqSy9/PimhUDAU
xJKM2wJgmUUY8TiGhIxv1wnJ7zKqhwcbfgHeVMKECRYd86Zi9mVuL+WI6PS6yJyr
OvwQNYuobAMV0x3KjE7wp69goL++3LyyjKSBaLQWrpq4bTLFp5XnVQRYKqidBLFC
WmaAmDras1rmfBrAXXK+BQAw+GwkIef1NPFMIooxh2XfGPrao8kQ9YzMKX0CsScY
Bg8G7sS/+mr+ATTUGywfa8JUJvXvYrpEgJYajOj03nLeosi/fyaF4xSITtmzY9Go
/qPuK95bV7z84lxjQlzlqHOxSpSX+V0io6fSHWfev4DeJjvqOLAUmELb2JpIwxrF
pvcMMHhoX+0U4Hl1phEN/6wW+HIW7DX6dSyj4vx2Oo5saCrPVex4gByoeKD7iScJ
VFqXKgwsmb5f7cE0zoAELSjmN0kZeUQDwsZT0aciRx0pWLEzK9IQzxC6sd2Pws1a
l+RerXRQsnDSZb6tDD8jyGlWiFj4LsAGkgxU3y9lvDrMCOTA8Pm34EL/TK8uQ53R
vhVn9mjbQHleI0KCJ//9gABKG3TuKeAnIF8OSb42Qrf92kCu7B2wRFQbofMg/OK5
Wopwy8i9HF6AnY0r1KOBx0s+PaMnaEeE2nQa9F/fDDCurlPjqeUc6YzlP6fIxjNJ
5tsa4V4fwBWAAoboTOC5YZw05mM4ScN4AgBQrGt/tXFFBeiFA1Ca8YNRZFzYFh2x
SFzo+uYNpFPrA0nvBQLP5vGc/ArARu/rduyvm/PAkcCWnCHdpwuX4pAARHDR1g3x
rl+y2fiPA+Ccto9Y9J5fyFno7d66cG/lREuDyiSekvwkN9lysV9sxdhzoWw0QcBW
0qI/GQ3rG38aIBDELLYibECH+ZSKcP2B8dgjx3pUL1gp7roXk2IhRZyQDBp2czev
X6attRMK+lOp5elzbl10gOgLGEWo6s9qn6TGHr1o6yhVzy3+Qb6sGiyti3Yjhi65
nR+fvJ18FMmfWuTHPuPpbu/Mg33xMkI0pnUVF/D9X9jnEMMpMT05p7DfjfNsuru2
i23d8CqHQerIe5QiNQrrEOkKGTe+h/RL9lLYdVk0nN2CqaoPQSuHsw/Sb5yX5LJw
QPpFDuxVvVrcMb5IbeuCUegWCiuhwUsjpCO8H82C2CthQst83d9g/xTO+HsXOXZI
ldev41nGA4zBehK+u8WHT6/Yz55m0AmCBYzaBY3qNMjJVRDqV+Hy5bKbyM/c5E6n
FGPbAAG1ocJujaIsRkbXlcuWI79LwyLON8tgCEKkb9Yb5ytIeojayhioISO9JEBq
fbuGLQU2A3CKj5hvPOyk5JUyGxDaaeniNmrqUti/imGyZubMxmcFCOZgeWu/KZXk
7VrHylQAkhhihHJjkmVaJod04zY25KO9P3JYosD2sy81WuCN/D771ocT+j7Es8AS
MWld8u4nDAO47e4txeBblIRbXgN7j2VQu1HcxV+BeolCdsioEpYh6vpOql0Nl/vi
2rQv/uOwPra4WLZPmdxTWBthPmubxd8mTs1LVj+Bg9yJT6is2NldVO4IO34WmOvS
LHkDsprq77gzpHlZDDL8QQAhz8cX//WUkvgCrHn/GstXaCYpTbBiGcDf4YiaLzl5
jRutV00DTKq7tq95VvPP15CpidlagSUENvJYCnQxgnC3fd7wK101JzxBn1TmpCEY
sqJVISHlDuBycxFLKYqwh3U/Mqtab0uIYC6UHFliMLHH9tJeFhCuNvwKG79A0iaR
O1H4csngVIm+3lCmcZdsG1sbobcYsfZbrXkV+Xk/AVaRFNi2cr7QjAh6azDHCujU
Oh2E9KoKKOOEWa/CpgjEZLqmZmVWPOqe8bxKl2/11DCzWgGxlp/k6k1preHgnwYD
r+yh54laXj9Raj4HCIdeuPwPuhn6w0agUQXuaJ0jzOFy8ahtUQrPN46TcjCa3I4V
pNH9vX0zbB05594qjhJ82sLNaWm6zwrwU8fOBc1FUIOvmgGVCkkmEBWZiqZvQ00W
hAEh6QtFZMGZqKi3KoG5T2ve3EKDjg5o6tWrCAJ4AOePY24EsN91B9J1AU60DORL
jvpFKVq7KQVB+6qhQIhKDd5ConMOwPVedivBvBTpwGTOI5v2+FcRLrrO64a7zEAf
yEWhBOd1CZjJKn8xZ6dHpOjqiUCFjkZ/b3C/ccOTWZj/YPuNAYgtX8KQ9NPsQLdr
ECTI34/lj5UnTtuqG9lQMKCndysOq9WQyGTQPsU23HC/vC+B/cqYFA+huqig+X1O
l3EgjIx662IDM8160r/K4DxV9suaiHR2/ZyErk5bskCAeOfj23bkHAX9tSAflzwr
oOac5Ce4+CTxqbZIx65LzDoo7bejD1Kdu0Giq7O6KmS4PFdvwEoti7zBzqAzph42
IkWr8HgH0asZol5OeckZr8L4wgIHtnc8fXSnYEG8knU+2FGl7redR1DMDpnQcjbt
11NEDms1nF15eLciSd+McwUPa+9VoJPAOzAsSlULLEQ74piobxOZXyqL8+1tyvLy
FUhHSuLeS5rvvUAAeYSNK4wxNNLa1dgzqniZHOPHzqplADryQd7lvIbw8gGRODx9
j3Qcw9h0K9sxdetgYSSxZU/nbxFDNsO51v8z4MVOGuSyHRP9EhT43GAh5qcZSdRp
uh01Ng0p+ONbZDLX1EWifakBaODKdeGdHecuoehT/xETaLs2gIOlTpLHGmVStXQC
mSXf+d3u0c8J6NL6l+reS9kyGb7QmomDkjuQyR2r4zthiHPbc5QYG8WCdBZpnuwY
NjPvO+Xc+9KNXwwxh3yPkYWadNcTmbmKOdRew9GOCpeyTw6nbBq4JiabT2HkxNXW
e8Q2qbS1Xy0aVDUb7MVvLoqMwz1Qkk67b/k1TBUEhIoAnqwb0x7aIpa8vTu4xudt
6IqtGNVkyG8fFWN2cFvV2eygVTxsjlG0EAUH2Hg6ZcH7XLNRL5phCir/In3btoyK
hfcaR8WDY92nSFzn/dsirDUJaBlKmAm6GZnw/n2cUHf2SZlMCQ9tEukUMxpnvtYc
LH2MfeMTNB1BmCCTjwe1nMUmZ800tHjfu6TyjFCK6/fvRc9QbOkx/+JomORE/cbt
EXX5D4vuXJOdq3YRPi7dGlUJ789C+dsEnBp2M8h4sZcksbuSSg36DVh/cBVir83m
oaE9GtK5EfiH756g59JrUJnPprCpKlGGmHjCxcZy27347QUYkCdkCuC8a2yfQxC4
bappy8Qi/sRayKoqIbnNgLZU8GbU4awpBmnzWG16qQdr7HXuuuGZ+/C1SINIFgow
UBq3WbQ6dVpbaMq2mQpktzHmLBgMzpnF53oEogen5vGXOst/GF1Zc7ryGnYZhNiF
Fx39V4+/jMgfaz7YiLLZu017+zwM640XntpRRzggPPjNblQJxo7g5io9WXxMPKxo
czC+daLDxd1YTg8bcxT9P6o4uHnZM80knH0pYjyL3YH+Qmr/g0uIJ+ypoZDtnXzp
QbrWo51iuWF/UjLLwF1DmXhuVrgwesSqMqDSorwNbiz3rpew1jmd9Vw4rYzNGoSW
L1ifiEJ+uanZ1lmHO9fGz02MxeZ9PMvCBVkg8YssUJOthScFs79kpPZtYAu28C4O
sHca9NkQHtYS6eU27nB7WPR9iDiqrqQDd77dflCwuyCCIlAHC/a0gKVrzlRImrlZ
IwrcdaAUjG3oNEDFWJnQm23ImeglM7iYZ7Vsc8aziEGhl60OeoPDOWyrKhw+b5nM
TvedSngmbJYVesYqE0chpUK79iUS9EcbzsNpp4HNz/Zh9rth+36iCVb5LlInwptQ
vm92zXVeLRSsGIOagpFT2mr0ZgEJtosbur5UeJ6YnIMRxUA8YYVfbZ1GdGlY2Trr
UgDb0ZjtnJIkS7bTImw6Pltkddg/+ab1eSbmVk9BdDaXx7DIzOnXilijkrl09ilK
nPzja3sBe+HvdR3ADtn6f1gnj3n+8fqccZMc2iVKWbcvr7JQesY7adlohorDIh0W
ws1hCC3oJA/uqG8xQI+mF3ls7WhO9XFmnZGn+4nCN9mpI2isnmt9tQEeS33JYPgz
r9zgmqyJhyeomPg2FzYia3VvXYcmZ3XH9h0hIkdvl6mr5G1eEIBDQZvj8m+/T1W1
nJ/wCRRDR/y3Rsco2EADUSK+2cSCMh6jUfbikhF9OgrH/2115+wfbtK/gKpdxRQv
YXJi6R6PpS/oIx4PAus7PCOIlMZai9y5+MoF+8b/RwAduuBMF7TlpzcmowGgATfG
+0cRxQHSXVFekYVvWtRMlWiR2VJyKiDTVKdFbp4U+J8LEGo/IzTFqVs/m2QSFa5c
YN8C5CNz/deGIJoQGStPCd6Qc5I2emGUp+i9H5VE1/vZXxIBZO/FXxEopY58+6Nv
8AsOzNlDhGFNaQsbs/IWYqEbATVRiNN5FC3toMVjI4xmM6p4LW2xkDaXU9v3Ok4r
+FTLuFxJTAnTlkLkaY3vOkcTxfbr/NNqIEhBdsmEuIrEjpsVTYjNmQ25j7n2c88a
kEa5lJAQMfuICI8MWqeo3SW5LKfj1TlRRkhGiCTsoemt14Oaj0z0FutMPDP3PcCS
EXcJ6YjiEi7y+NChVf4PARlfXL8u/oiSjNxqJQC/ASQIrqlmnhoYpQreIyNMQ4eg
HcNAUMdUw8rAtZuv/n2WlZw6+v50AwTqnvUiEXf9/4V5XyCB2Xpbnzc8cvSdMPAm
PNaq51ToQCEqJyrMFUarMOsY17eily0xpn1SRJ5h0O5H9mg2lH7BbZMkSGY6w3/U
UT5IUUGOET/IdGROEMKefEw9XLdr5HyUW+6CLbFzS4+RNJyLlTLaU1Vv1SXjK65o
MwZBHkOxDJ3O86QYmd1hUUDlkC/EcTN2N/F8dvkP3kxXoqHHP81GFrGBrS2Z8+0i
4QoK784oig30KCvXGD8FVgtxA0LjSyfbUEcpPQTB8gd5jq+y8b8wor3Irm9TqN5e
m+PkvlX2dJD38exYQ2yLHGcQaMaXEArTg4TO3rB1elZ8zoVId+LDzhdEJR4Z55Kq
VvLLyVEaIhJuyq75a0Q6HwO+sWZs6qESl3qwURhl/YImXogr0IoeC7yGMg9LMjkW
yXHJuMKSYJvg9cRp6hX8R4b9eaoDbL06Y+X9h/iNSDjNddh6+7yaw0kBDRLIvFEK
SigDaUN4/BjOdjt4Vw8ms52DCsV1D7dvKvH4FmS2qSpF/VdOPy2jiHOEVZ3TLHOs
Ilpck+eW1OHJ05J5IE0WoF2wOotA40DasrsS4OOi8ImMENkL2VCSPNMCfAh+59Tg
vqVhDTg48xNaxsWXpqxVtbEac73QNNeZn7PqKAY7jEdgvScqQeRrKN9bUHVV0OIG
Vxz3Eo70WoPZDD0x7DnwcYAXmwvIn36Ix8yllvHkq7jui+HCxT7PSfDEqZnY1R44
8CPOdqyHmuVO8ihpxy/4pW9PKxx7MUOAMrH6EzGpQnNHzeuMEdWxY7uwcoFfj8hi
d2gduus8k5CxJvh0ziyIO9FJLls/JjLDJH+pytHfCPmpyPDZ8IOBSJ+ugsK9i4Md
jtBY9MrjiJqkvh7n9diAqO5y8DZi3fEFzlWMMcUrC4khflZYzphHB6lLxS+MpSIq
D6qehAwG6MHC8fIzg7xyxk+Oy00FLuNxHHRu4VB6/Y9vyUsxmSS7Tx/r6mrUQe9m
mQedDhkQlc5P5AIn9XI/47hKTbX4AVUJM8q+hPwELWEOnbiNNX+cyJZQtW0IxPgH
HFkmI8MTvBZPviZ+x8bpRHpFaHWh2rX/HTVogf0rK1ookAojvT7nuRZ8VJ85/8FA
WVWo1m40ccbHKGYSpZms6aZ+42g41ybkFHm43isWe4SLytkM3NJZqe8DhfrkzHzJ
aGgu1vP5fa3/DiqLP2IrR7G9irpVW2uzA+BeZwrwOuV8nnKFJyVyIN/jm/W7HDw+
V4f9mvtetyjyAKNmllNzXVAR7q0EXJR+LSOyjBDSdbsgiKlbiiWoiGVzR3w4KeA/
cS+iyOUWVgZsrD38XeY8aZ292iZl86jncYCyUxaxOm6oeMZrns6cP3ehFllVR0+l
Z318dLxxQUKvxwT5eNWeMbmwPVbspZGJsXQVcvgtB8ams62S4C7LNsF2t3TeeZNA
o3g3IUqwOdfnh4NeEbTukza+gfFLnu4h4IJUbDZh859GXR9qyectxDEebyTZUX4h
h8CSyp+XEf+giZhDVT0TanXh9/D7kPnhCL5vR1i8CKI0rVW9aF1KYqDn7PTAh/6c
bwLpjLgxdUsCGlvy5pWpQL8+5ZwVdu+mOM/HP8noMaMx5mpBZuXhYCB/osFWIhHs
WAbOgPClF96PY4+Nvcao407bJk0+31zVfz5UBZ620Bbq52inm6UA05TcfJ6Ww3GV
LtZrOrB3GzDxD4vB5atSatnrIokILbserFBQXuK07TkP3s4gy4OvEzc7Bsc+kCee
uvyP8qAVplYFgcxtQlPv1yA/9tcp9auBVKgxjVHqBOqRkmnrArRfBY/VU36b6REu
1Y+dPFv3zccgRpKGvqVxEqivdKON73NqjSzoNqrX1J/D4IEsT5S8R1C7GsbSObE6
FcUQmYuuoPw4kEbcvbByL93GAk+2p7/W9zbx8BV+9WUu4YrtmsrLFiJ1pMAK5HN5
EXPvxcKlfAaCXJRCI7EZYtfMceW8IWLu6z2/EvwoT5ilsdszIRtRFakX+Nv4EVec
/ZCdIQEbhcerK+A+KPZVh9wkcf6nUaGPhQeuito5DaDBlXRzx5rbW0/fXgN/K4u5
4HXt85RH+XCAfNiaRRu4H1f9QsvmusSaHOE/LOif/H3dc2gHjAdlaBKfldJKIjmH
Sgf+9pUsw7aad/7hIKImP91S0L5UqZVMkkJOASpHnYMtRot8hHVSIBpZz8J8iaUD
sjpHSglUxCcV6Eo8f33hZ9ztIcrPdlst9IyTqat9UBrjrQRET+D3js/fJCrroJcS
XyIH6wkqpHBq6GSG9af9lnax4WYnl+KHAhr8cV7YDtd2w6N5JKzRo97EbJTxRQAr
aQ60WZ6HrY4zszHUrDLxFC7s8eEOV3U+ubV+vp4r+kwgXj/jQiiaRdrHhHPfJtQm
hWVO4Ti0EYLYDPUOmw9ZEzCl6tm9xBvhW8fK/v+1vLu7x/BYq+KLUBKZ3sWVTwAr
HKuHqI6FfkOKb464eUTRRnTtkUR6wigIHf10AkOzEvp+i1latzXiF303pUz+lzQx
I+p3hGb9q5CRwFQHKTBPPLl00xYGmg5529IvOHqtZ18p98ZcMx96qmzeTPRIh7Wq
0IAc8fPtESWxpL6DYmkzbE+e7+zbwkS1NYQqFdkqvEwFV/HiPMTeze+HBshOXqvN
UpKAG6Ivu1XOEofATrjxubMws0aeLrf5PaZfnyoUbY89wVKY3UuQynLehS/musMY
GZKYxhw/qCDmDBovn/pOkLw2IvRhGiVL/yTJ8Xb59fU6kyL+fDR0nP1i04jhJvwQ
jR+OYm4DKKP1vFApYaRATs22MbCDP2ciHFMkWZ++G4M32WHpS5e7xY84lNsG1Ttc
m4T+dbAkMfkgvO2n6vhgt+/idgg8lTmEzo+vrAeHE2B0A+Y7azWoEVI1q7e9NZgI
LyOIE2BqjFWQUfR+tKaTsw/Jorgm8FEsjyqgBIRti/xyXd9gsdDRrpBP1BF1D6VJ
0wvDriH7vz0IBfJKBWmF4ZTVCsBeIEUEFMmqopqsFEtxFhRaq/ADJ7TM49/Fcyfg
YpNsBGKKJlDzsoP+aqiDnbYwd2yohCsW6mjgXkESCFAatPMnBsMaokdYQStw6Hfj
5sWOTbMtja7i9jRcaCG7bQ+Dj8qBQLSWrJ4Klrcr9s6vteZvoMTcuQsfiKi+Liwg
zY30BPcZq66VP9FHyOfOTFK8US/+PBS0HJKDGmW02umaujooTdjwAPuC+7R5QDai
Fnigmf0FC3HVfxcVD6BJFj+qbNY5UuubexIdnocPZ8n4FIQPE2ihDlFRS0sLoRXV
0NnWWRAASu4iLnLqA7Qp+nDbZprkqKxNjz05lRipk+C/9X8KhsGnkoKIBjQyxxl8
u3AfTmFyHONX3Bjc9AW988B4mgy13qS0iMfKxLtissoB3SSeTmMusAc5+T1vGlc3
uGuH33QNBMDlGCU4Yk5mXVbSEDKdPsl2V0VKxmKxsrHUx0yeeT42409nxES6QAOy
Sx5SfqFfFPZ4TCD6KpwFwLmzu/bVoGlxLxC/teAZ3VsQsEIW+AtSuFEvhMhg9+Jr
LpplNpCfgU5Te6EhtiBgZAH1eS/wOCXSXoS2XFonj3/JCzJTu2J7jruVegI9lfPg
VlJVgVZigjGx6gv775x46/nwKI4Ia6Bi/BrR8gWA9Oe/hJmcW+v706R4hXyQdqor
WshsxxYmUuvRpglWxh8afDstCmdyjjgUFHum356OsM5kXKeJV3za483/l0hFOGfa
u5MMnbzFmDDBIhvjV151kh6oSqidNFjiyBDnbbY+9KFLfZsyAUdmSFtBAGqqX0Vj
DNb+KE0F83lZC36EDYmcbTOVXSXhzhR4vNCvhA3SbIv6JPEkAH4YlIfgbzVMitkU
jYdJfmmNdGXj+wS1yryRCobj1mAtR0MTh9Lrztx9BV78XM6e66WdKACa4S25CQNo
Mkk8uBqRscvi5wGGL5MaMZm6cjoIFDYlNsSjLq9DHqd6QJIMIRK/ImTEg7nAzV46
oZVw/7PpXyRy07kB1xhVUo1/fwF8/aM9v9FsxfcdHfISdsaWhB9JY7t5Sf/pgycF
/7/P7ws78qPFGWIgpMM+S/ROEJiyH4LINMQ9VI4UvkcmMcgPhj0ANdqqVXWqIC6d
QUPRkHTFrp+uqJGuxrZd5Wij2c+59WVt+kdgHMOW8/3EcmfT8P6auxfqXKt6GgDV
LHciFaCLI4ytNDejLVT76PMDkyCPD6QrUfLSpdsiXdTV/O/mfWDwO+uP392zHznX
oYcjli+vF7cNbPlBoBRH+0kPDvVmTc0KO3ujMzNTqqrP8F1ndJ2kamVPbL5/4jFi
i9sQCgdp528mmEIyNQdjLzvG8Gl0UqZ4wZu4zVUzOrwt3ZTtNxcKI5HfhOJH35Ya
eoiDhSfSCTvlCEBwFfeZgxb2nhOebCy3tpVm6/Euo0PgSc73QtrVaSPjkzPgVELT
FNficT0okNNfiSgS3vg+oBBKHLULfMmG6VF9FiFqrJSnsDbfkIQ/7jr4iVdpxnb5
Fx+eHMYtx0kSjCEUzITKyj/bVkwkKRYABfWfgkrQNFwNdfnDAtv1o/zawJ6GHNre
BzFBi173lLwoFxhUw97EnrF/g42S3qAY4DYJbqSbMDxGCwFR4DgjJg0RAJ4YiHU3
rGCns5/1SgrNYKnl+qOCEgOvZxil/M8fKvjq9s+JqDkie32y9IjKpJGyPUJJnBJG
nsvHdfvW8KeubjLhN9bPjoDfHOrEFjwXamzpP6aU7V/W1iln4z3j76FUmHybkCaC
gVvnRvGaNBPXkBZcCcEJtjTk05Av4iT6ZXGYAXXhOvJwFsenyR3xryc4u6f1+EhB
UipIRs6txcv6yi7ktBycGCMkMfoenbESiBu6zaIKmf7x666ot0VSEmt57zSPICY8
qnREPj33lPgxGmDv1ke2RRYGM0y16DoqGxrWjU4DV8zrRgRP86eNJQtJvpm8iRrk
Oq9YV/axYaPUvCUlJeF+cq6lpqPvHksowWmoUCQ03GtiESrWARi5oYWXOCoPzs2S
KVZb2wFFoQqzg2IHo6Teh15mxRFVJPiH9JaQBZOBZtu/6sMGBdo8dqESC85WSsJX
LoMYfci2Pv8qTH3rG0+h7vRhRap42JYcG/fxLronWaL2LSSR0YP1SsnGzj+DjXQH
9yMOe6n1pQZ0jK3/iB9WtAdqTe0XssjnPwkQAA96UZtvL6+OVl7DcOi9QS2tUwNz
XUJzfV2qhnoN6KZh5ELsSggITqfacyxc3gQ4OFrJIpywbfEVJ64iB+rhmq38q27o
5D0rHkVCgr8gilUhWZZd/aCNCqSdczolLad0tq9GwAvE5pTkH1jPGw1SEywZH02y
ghlRAwYVeOSdi9FYDbzzsJmSbz+/5jH92P02kRdWraL2VXWB7pUFoWxUsj5FFwne
XhBQ5b60xnwV4MSV8d/lpzfxt5IKRr4ZEpWZSFiLlGjh1AyqZOqCe8tMK42olG7f
aXCgwBS/tdQxMZCa0qmBKWdAW0/1odQ6n1HxTMmG0q6GvyNMcNc8EOyN8WSYlk6b
MZiX5ntLWOM4ur/lm64xd+yJoIOT4VTnjeJmTlLqbA8W7u7WhY+hb7f7HYX5FROY
U/PFISLJ0Miq7YhCHEgxsxUlKtfb3c4VlMjnTxAxucABr/pbI26lpxy02btAMiHS
Rf448FSjILZcS92YkLH9V7DowSra3DUd3Qxr532MhFrpB3Rxn/Dn9KzEPh0LLKrR
0/WyvyIj5B1wGq+Z7gkSSdpjf8JBA2j8GGVC0Mu8bpIEKQNpv5w3/ktmi4tF0Rku
t82W1oiFBih3AJS6ez8X0bv47mWNBr/nOuY2TM6YpHK0gI75pLEdD+Vzk36vsgiW
T5NYoFgA2aCDmMjjtSOtyD0kL0kFnZ3sBD2wkStKAtOWXFXXvRE8sYT0nCz7FL2H
tnmMIM7iI5ZBbTwjUcowpEncJuOJDXyZseUpsi0QJfyRmasQGkR+3P1jds0HecCx
CDSfyknTenrhvNuX6I+IVfjJci0Uva3OanCEV3y3wyUUlGuJo3RJkjKGqrHYGCVZ
nFHrrv/TQOJlhyc4VdJ917XXnp9/vIvZksiOMOBthOvRn23CM2HJukKq/SvGm60B
0k1NeBdRLeqFtYySQ16TyOA18XWq0/Wb2yIF5RRB4OuTue2k2f6ae81E7xUDkPal
WdBLFdb3dTg3KFdHMx4uB3s74Fv8oGlLWAU1RHYzpNgqC0ngwdiTjpnXjfOe4luB
6qJ0PSG2h2k436cjyNawcjGLJmBSmO+wZwu+kTsFHn2Ke7ZN8KJKxVnTQguIknkt
utjemdKOIEqHpf2PTFUbsDj8TQ5wBgDZtX9rZXzkugLuQsalXRrZSSChFwAW5thw
6r/9HmMzPoUoRRNneHJbgQ4oXejsIpmWJO2FDltQc+AUaYgpFY5XAJkgXBFBlcs8
fa1GMwohwMjDP4wfUv/YnBJo32tqtZmotLOQ25wyT/vbvIceYXMgGKfzE4uTT0CJ
hYGL3thPeBNGT3HEFVCi4es7OXoxP5O/m1MyhYRxNeEmxC/zk8SEP16jBx3v2jFv
D4KXNyT9esJ7NS3CW9na00GXhcSub+0HfmhFbtrXdYadK+VBb7g8GWhH+yeSkMd8
L/S7DMu9g776A0UwaptzKRPqtXzknqrBUV72jO+g/bI5KOUJPSEDgq0Z3HaEYrJy
CgneoIh9fzcdHVtM+xAYJDRndsa11jLq0n0wgb27JOHz+jugrmweBre34oV3FHtc
mBDApVIhpuU6b8Ga4+FD4mlW5h2o6QnmMI+ggK276mPUnhhHUEM1inURP/Djs2/t
mmjp4GV+XIVuG98raAA9cq5L6+0Syw70D4cSAanj4O+2WX2TvSrvHNoQOBTqoxSL
oGrexKlg+MMbLVeJtsf4DspiHCsR6wsexCOTFJsN/esRAObRhwQbpffYr4Xl4AnF
NzsfxuByAhgozz3YYVeIZRlzf7iORX9OzDPlioOkI0BzSai6uy2qEv6QzYm/sBmR
K3nP7cN6hrwDUIhzv1SGqjwVDOGBpfn1Npr1lK0CzXZghmjWHUc3ClA4fK8u7vhE
PaGTN6xH5WnhH+2cMuZBDg5UhxHOoVTsWJ6c2dKPhYBjy9rTZUHprPF8q4We8WtU
Agj1zSLBVbFB+w+8Hv+mNjR9+/hKrjxzAXcYE+BJdpousfgTtzXsA3w4IxZ/BiiT
iueoXPZvzbxZ9DtlDvQbbJO3xSb23IeC31kzr8UkwOy/FqpXFWIwSzLht+QchFWI
ukKf7MhmFSkqBgoINNbv6syxBVIq35h0V6m9E4BuAnHatZnhfBQRO5jYSj2NrbkH
8tETRcuIHNgEtIjFsREfomWoM94fsQ9+2Em5U0SxbBxLK2iHd85gFsXR3z33Sdba
fBMbvgg7NNCUXAzh00boef5gG2YKYwj/Z7LLwV7JD7cScd0U5+QjYVRhYVsnCldJ
wjIjAAgnAJ/V4CsvZx2ngVIujq+cXEJZqPXAWnU7ZE/YxeYaL1nX3OTkDZD2oEze
WW76T+7QNxMsTCsw59xkFEUyvB6OmKM2ASqk9qpUV2sH4kbXvVgU726g9FHnz9Gj
Nqunol0pLNgPNzVyxt0hdoJT0XMg5b7DUBp5+ti8Uls9+4Bhk02dSEmHS9bb/0Ow
RJFtdgIcw7GkDoZA1C0igqUR2inbN8aLGohe0uU6Vj7/ur1C/gsrEzLONIwN3TbP
EIRmh2bHkVPNFzHTxtZwE8hUN20tz0B+YhmrKRqzwMYm6kk85Cn1vgAjeFNRv75p
FPi2YkZBpDQpfkVFkuWcqJrPUJ/jdp9W7UFqzEQPv3EGdEYiZnWK76k+l4Ljs+bg
HrkJZbIfLkXd0WEeEE5p6OftSKZiVQr/nQ38BuoH8SJAM1XrmoNyq2WEu31si7qc
ME7HYqQA/6iQyaQM04l27sPYCrMrRdUbKORQeS2b0+EwjL1OTx9hS8ePrQtzs2Lq
h6lbCs3jhGzQnnWq4Wt2VI1Y4s9o9LQYA7MKCNlYULSy9Z3uH3CnxZrgSvqhlShN
swN5Y72g2Oi00NIoDghObbmJV5BwqksbRO3oNMTzLm6cBr1vlYwWsFtKcUzhM3bK
PAPdlO414DUqg5BclWgn2ZECqCio3h01xOr/4hP9JnlxKIKFWcaC7KjWIT7vdH97
ezUuiEY20sJi1dtx1rwm74dehyMRFDETC9He5ajOFMt1VYnShS5g9py5ZJcXzlEv
hIBW1Y3ddk5HV1plEhQ9m+IILN1jra9nZj4KkL6Ctiu63rkfqYcR+HU+5dFOA/Dt
2nlf0Q+bTUGYL6QAIhFrzJ+F+uhuWE3gdTKysogxBuQVaZ2m1SwfXBOrMoMck20p
sD3xOqf2OQP8ejDHs37j9mBYFVOOKbn3sC/cUIBLbleyzE5rzmAsOM50GUQPt0UN
HT7b2IXRX4KYwRmbgow/eeS+tSC8LpPp73fv0Bsjekr2YjiQyVFVVvT+U1e/nr0q
EXSzWTwAo7CVO7IhDtnhgsTDVcwZm1UDUsCwj+RttLGS+Szxekkv+IaBvlZcGXG0
M7XitVX0VF/2+6ZfcaLbag267uHXSokhpkP092u8TVXiGZnfil5dAVcT/JTx7OPh
oTR114kvc8G76ukfMmYyEgV/1adfvrzjRNHpH6d75SFUKItcEBsF2HF5jG5I+A1b
ybyjPWoeE4JbmsC4IOGsTgUrADf6NFOtxfRUWrJja8Z1mdsIi2ePRCGlKSjW6MKS
E+zJK/4iI3UbWhbkbLiIkgEMzk7yZosl3tNutBPXyXH1SSDyc4mhsFTlBoiIpREn
9k9NXw4llZrLWRLJdhre/BHPDk3V92r84f9xmOzCViSBXXEdCw+srQj6AB92ocT/
RT+mSma/3a6MR9CRcAdUXFpeiszWnxb+5ZSMjVT7tdfoOQdBgNNxtEvmFA5TlIKQ
dfNEEL6noCaeiRnlDhBQzO3aGZCSwKjyc1akHdS8Pj5U3V39Dp24zDsxSwcyVXkY
XREVc6eo9wLVCoqTnmAE18X57mNd5txgX6vd9dyRYfkO7rvMRAyj+cBVoNZ7kPkR
HC3L92W9FajvODos1VpeQNIw9VFR5IVSCjLAzhGorId4UrgKhjBXhc7t+Axx3z4J
12ufGd3kK2tn36Agm2woAayZ2KFyIK19NM0dudtjo0qjrCPcbhMLjXxk7AP+DRXK
Ifz9xaXhJBIdz6vNFaHPiA1PjmvTuUsztIp0AB7K5fhzgUFk2xfmm719mB9AzOF7
nBhNFkuDBGqEpj7mAuZhQpJWIcEkv1/rvnfGbJHjg5IPvLSmz7eHHnVIGzaEkYGO
jshy2xDcOkeySFd1UDEeV7V1yRDUgwPvBaL8yYbE3UPwVScRmXLgX9BWTmVc1RwB
pTpkBm/lWIE6xOHDejjFwOBXvH/ffNcd1PgOQ4jN0TSwDVmUXLXj8bwMu1Pvn1CG
pM6XXONzjKrO+GT8Lqs1aWMZ2inaP19nOg8I5QxUXhLZBO9jgCP6zxwz5Ob2d+K8
w4fVpDz8aGvxSdMezF32qNOuSc48wwHW0MnN/z+W3J28s4ippGNczbOwM3ihctF3
UuhC7j7050NWAeNpam671cAeogxeL6OUG09GliTHUPnu/Dzs7VS5bmdJE4r9vNih
mcPZzE0aeQzZFxePVqRZGKKyoHmFmire6+l7hKn/dBcO9TQytdSCn1GL6sN51QGF
RSnUNyQJJyyFI+0RPbRE6wS9fbGyAcAwHdpYvisep5RTCGLX+BCIMJJvd83fH79/
rQ4ERgcXonrAPPXRChTvXezDIuMj+RQII7TsNqLr9qroL/qNrRl67qrX9ZiMhrB6
b6ZMe6nKv+4bGa+7s1/nUhwb7hfijuYj3u69srhGZvo1RH408cX4P5V4+YvKomH+
yg03nd6vg2PoDIARZxd/78bqTSTAoVJIofG3RkscLOFxK+7+rFDi1DSyBWUTOqhI
mXE7ItNQbS5iqNX5ttAUrpw8MPOHzNuHYf0TsYTP4zOeFjTdNYG1iTIByS4QZ81L
hXHTLdSZ/vodTU1VvHqw5GSwONiZuO3oLS+0xOR1s7nBZoOgjerOaNua9CX61Sm2
Zj60b3nQSa9Ygot+f2DL4GL5wCaL4d2ZKXlBqOmv686Fiwvi+gxVfb1bTASu38LC
U/VpVAsmtif0ttU3mvsBhph8XXimwqpExhtHQ8mXq277w3QiVjmbJ6KxRiU5c9Gr
XAuK4gPs4F217i4nJA/zDS6ixnu0HrbanIU2tuHJSHpyVx0QaeazNDuthhBpKP0S
O2FmxfWq6nP+61U2M2vPfHJSR8dIrplrn4JrFFbt5E0SgAUgAh3HrRmVXX1tbqs7
x0MzpR7o0RFXEFsaXykt78F64gPkqgz6THnTj6PL19yW9KAx2OVH+DhJ2WiOPFFr
3hwZV2OcH0dvGy4qceDr0N9vRecYR6japTs5hSNIrSOwY0MhC42Dtp9tzdHCt2HV
oV954O51eWrvhB1cpJW9EQjFyAOpITXsRuCDRYZX3gAUY9LMcKSF73Vodxnw8fEJ
UjDHYGWCnhRc8+R7dsodEau45Zzjju4IjRhWZZobCHIoSSqjVzpgIbls49m5dtka
nHSbVxTL29yPnjNMJGunrKzl/VQTTj0+AVfxFXqLRZXWEiYfxNQz5gLFgq11DGz+
gBbjgGx964yVwEF9IaVzae+GIqzyAfVl/ZHR5mU7apkODelwVASWRL1+v4kKsU5a
8fw3SgBC+7RkbJnQtFeqeXpcYo+HZg7iYFkoHXVBK4E8tqBWIZRjOLlzJFyOhahW
/JrrajXGmyGaK9+O3CGv9jTaYsNfXVotKp7WXYE+luYyqFunnEAyacEjyjp2PYAp
6/aqFK1vVssjL8te2MGBUMqrKzVNueI7GwbFuxbwoVN/t/cUbz3ef6kjzbW9XW9s
GRZdmCsNZbQe2BQ7vv4hhhh65lKVCQX+SCQ2tx4N3tqunJUQOpBruhd3CA0VMBnx
EOAJi0xDosmbcMkKxsZ8Birt+ar5qubqdkW24TX1nA2S6Y7Ft95BvUgniBkwT/Ze
epIGrI+O5BI6wMW1B5gGpoOOJjvAFKuGaCh+3VWfZsyoUFPX+GFZU7D4Ax0n0X7a
KKM6ph1bC8mu36ZdbfAah/HU9vaAiellL38QPOY/hKLgulGZYxaqkFRvO7WKKyZ8
4JKqt+Vg/GSimmmfbAyNjsIj3GmzpzllnmodSySllCPxVbxfmABXvwIBoSdZOlXy
YUu1dPErjWqFj7jH/h5iRRHMIaxgjlj7tODldkRCXqr+uQtuiMQDjbzOdzYBwbjm
EWrvUUEKQReGfWb+OUwmcHZfxqqHk5/kkwiDqAKBmqZYNuorHY0kZ7kwQPNgqi6c
qTB53kQPAZHohgo8YqU3/kgiS9Z+8Vx4/8Xs0mKwRnuSMUSNtFWQQjCEQnrYSNvl
DlokDvac0L4nlmAQ/o6HnsWp/VOlW/q0pbP14gw+XBz/FJJx3I81EMgEUCg8Ap6b
iDHYn09GAqcMkfbzAW0+yb9C1VnV9L5YtuwPFUQEnljx8XeQ6k0K6+VDEbicn3RD
DF9GwUWG5bvQdMynfltBrovmzuZHrqlZ+qR28/p0oA2M8O4xTGfBSPYBf7rGFvEf
pa3tTsDLOxjEzs1b21OIZizWSmF9KLrW0tygbK/H7WNNmaujEt8O0Im2oOmxgt5h
5cwW3YMgYXUrEscKbZfSHzDTr/YUL9Xvhxw4X4XcIbAV1+FkqTa3q/QQXRYN5Lnb
ysNAV/tvafBNAXoHI/W3pHe7qRoV/LUa4VYJWRx0Ep0negCe2r2ue0Fq+Sf74LLb
6oQSpwbX458WrG4Pr5KF068L5ZJELGDHLhscnVAz2Zkdfz/YKqW/BsWNiYcyFg33
0yKaB3F5x91OAMITL8RexolEdK02ZflcnRIR8/XfON5/nVtfEWRwbuwhpM5HLpiP
KYjA9xBBTLfeH9SrmeoeqkX6iJmTBaNWfn8fX1i+TZjl6XoDMVPgJxF5VisImp6/
n98/OHWNRge7qrG8WTqX5aMTcUUFbkpayvEr6cyY23HweYRJuIGFVAPlFz+FF4sp
vXQIFST5i5b7GwykW2z4/2yFQdL52+sBo0p+VqpmvCchrcjqwPPN8PusNCxYvEEB
SfiWXTlecENRsLetYhYI9XKdqo3/zr6cWpbe0rMZtYl7eR6jkU/NnYaSDSIPUOKA
RJe8UBZn4xibVurCAQAUlCAXO4Xp1tCPCGBItJQnH19mqX+hwNi5jWZGACaOT4Ep
sjFLPq1T6exqHPRIlDTFWzohStJwghtq6Ryvv3V06lqNd+IMVr//B190diJYeYHL
RWTaaX44SmAAX86LfUudeo1vXxmVKKIslRPIskRho2aSnvRrqyBMBdqFi47mckpJ
VHmVlB5umaLKCh4nJc8f6HD2psXrLwW5DJjLf5XoLJKcdCV7W5IcEB06LTPzJ55q
y0lr9R9xORsmrsJsFiEfbICZvo9Ao5edEeJuDN4+epSKSPVDXvCLmleX5FjOAu7x
OYTwIjghMnTDtkl1Enm3oORWz00ZdofXvkwzRtsejqk40Rtn9vmolGdDYNBU4xvk
jGzzINQHo7SPHViNEDLhnK3uByi/jSff/Ehctcb7FdME6fXm0ydGRcmU5G5xlddS
X/eWK4XzRgK1rd84LKzATYgRqj5UK2zs4ED95cNuyWAXsucuYr7uEW0iyg65X56S
DjMvJhi6WMn4kRDFdjTnI5xmEWEuJcnJyZ2EKOxYVD8T2/+qRny//xhKVdggIAks
A5U4yRU8YEgtLY1iiN9ebpktSxZcE9iuDCvwj/n+jtY9yxE35QC5Y2p7EEFYMxVv
HDot41Rx4cYThIvxFZFE+WOdQKeauLO3jUR9J+om/D0m4D+edHgvG+tn2rUDNOPY
KeBMVlGlNsC361JK7hZac/HpFLwzPKbrLGlHip/3VpElScwveKbOB5de9zzl7F55
0zIqOHauMlAmEq3Z/v3cM6D5lOKkdbUkrxWDRysXSmEqD+LNP7ZsFsgf10RSButQ
pT956hKCyvwKbVSicURKAgUYypFFOQiW91UmjNzSrY5gKIEwQITTKiJ0NIzvyKXt
o1BjKbGtR9q6kcS1g3S/mg6Q5zuCxZM9jPT9W1sd3f+L/VZs4uNMoqT8tZqljjzz
vpOLpFPv3QWjsjJcv7GupQszp5sKjGjGX0fXhQS9i9Wd9enxxhacJ2034NYbPZzj
AUU9SWK31KO9MXpxPc9CcVjYRNWyUd471baJQi7gD7WL1l8zi/kuXyPNqkdVQOZ/
jxRVCx/4H94IlFVuTGv02c2sWaQM6xDN1fH6uuyPa+PB91K1cvE8NEqDODCEIvQq
P5kaudQxVD+3hEGVe/iVrxwt/dBLJ5pENlxy0jh3raNT0012wdGoZRPZcjvS53eX
52gYv1FcXSO6jLeBkGI6j+bhXNl7qTaLdkTN2UpGf9DO1k+wvKMQS+QX9Bzy67QP
bVmVMyJK7/Jcl8va5+Ymu6p4HiCKrTdwgC1lp/Ahwo0n7EWtfa1EOEPBhcihrMln
Ve3N5eMZGcQSMua7VZW3LbJZjZiXhirgkNnSzCsys8SHX5u3/GtSKmEXHdkjwiLR
bUj9cbt6KTlHEQlo/MPC2fBnMhSVAUp7gUYuKNVwyEA+J8V5eRk72OPbAj/CtQx7
b99b2g7YiRXcPNfBRfYOdqeQUR3v3aDaf0pc3LSoMdSyhgY9dPnoifpSPKskIJpf
o85Yq+jx5ZByf+IPxtVt+qvMtibchOZkjtYK/sQw4Ibz+vDotVeCeAaLqVnY2cpd
Hme5uqNxuWSGJPMCybZqciFWN+MEdez3Bczgo5khtROQEG5o2XyFPyVhlurBvQsw
m338uGdPD0qj/gsK+KR5p4eSjeE5FxTNYHxrQja1A4pMS05MvHQSnLo+D9skhB7o
Mtmx4Y5J/dj4O8Z/1lsxw2u40lnNPtF5lrjhCl+CeDIUZmIlgwggQQB97TAiKarQ
EH/uHJPHOVgXaXGSM429CEQUSqQsWr9p3cftphaoGXDRtwlHuYvN2rDqHLhANzzl
yJxByR5EUItCSr6loubc6TJEf9N0zK2F8Eor4KvOSgQEuwXagbDKIokRSSjk7Ffq
+d9Ko/lNgbgqfPEZRXvy5rV9u7tWCyN4Owt0eLlVQM15LmufxojB+8I6orvupPGs
QbGap9KAp4YNAd3F9BzWxvSK/N9G8h/vebtT1CpHBE0Qf5FuP588oCpPIoBqIkTs
GFAWliDOkyg1m6f33V0IAdUBzeNaX/E4JvkhWA+TqtVHDIoqad5z0nhCWyJeEpp6
Fef/XlNJIjuRNBhz6lvXbpiuV1F35egFuPC2fRyboYiukAN2B3jO7xY0FvzZcCW9
AjBsHK8DPxtXHNDyV/TElVqomJTxDjv0L2YKImMjopkaQSvWUkOZNIkEVVq1UYp+
/F0jujAXcPqA5I908vspcQthPDpMx5ZKC1MEyNMaLqGgdk8wdgiyhYGhSGIKJDAT
nvOJVkSYyGAH5E/byuHOf+q69eazRaOpEJYd6cLhR5F6L0pQzQp0Q1MhOPUqgE/N
qsYfm245+0ke84q7OHsgh8XCOq7KhYOZo+foFLTcHcYW5KCcGA9YQ/2qZ1EO+oUX
RZuI9jyetJBBz6+Uir1HE3GXc7df+pr42yeqguR4tH46DVioV00MwAr9jGF7udy4
nzRA2ypd8a1vRFzEIh4wyVz0GKI1A8Qpu57+BMg5jqWviD1Sxo0VI0PAlFJdERFa
LiDDpVeeceUXIEi+v9O6KRLKh9TOQT1KNya6tMbtRoCKYa9ZeBJyKv8VJT0B8RJy
dSt+K96XYFQSX004/NAye1P/QHhugmbDsvE0ebmyboZND1gHJfTPpbHibxFlexCo
a0ixVas37ES7Jn1qWyVnU+1/kCAYeznEWGL3elmvu4XifMTwltjBXzeLvt3VAN0f
7PweU/vmidVAooyS8AIJpOOZAEmBxnJBygil2HQDXNZe5CPUzAgeA3IYh3IYB4AH
PmyU76wo38rdRWu75YDjNG0+WfUPmLdDCuII0duz12N3+cfGUAU1CRyarPgNHsnY
re5pTn5cZl0nxFDrc1ZfMJ/8VuW8CikhrhEe6BxZIwrGSEAsbkX/ZWgQ1ubYZkmU
YBYoyS1rLyPqGp9XDd2i64/ZtH64ZM0yMEduRCp/L8m8spn8hkliRWwhwwhXfUny
/0rajEjnnVPTdFVMrzLGCKFVOmqc4ectwWHFU4+1ZHN7a1Gmhxo9y/JZuXM5PRtv
AQNHnus+ZsGh0ILrHRoPqrDipwGOYNBAOp0h7fqFC2aKMgPccviI9s5bZao0T9JG
DrDI7Bo6L39sfzBKJuderZ+cSrn/xl9jAIbEANeg3jn6/wAIyrUC/glGisKIlMJg
DDBtyILzKOpU7To3g8Rt8ti7VjSzjde4F/M/KExJqlm0uihwVbTFx7WaNRoxhHs+
qDRszH9mCIB66VCW1QlO0cnjmOVggQELsexVglrcixH+1ZYrXklVXuyWX/7kZWog
UxfclzLeYei2Sar8liZDTNiTexCZXUSaahB3yxsJYu9d1CU3QUwrfqrSRNkRIhm/
ZjAHkg/xhxTj8z1Q2Bv4DWAfcQCDc1y5mcWJEAyT6xBuZhISVEHfZnrQtNbasaHm
JG6FGThufqLfLcsIa035KJ2MKLt6RiiP93Df/59tdFdKIFVjXWqB7vLGPEzfcX6V
2qUo6SEJQCeR1z3zd/xo1Ttzj9e+amLCd7DXRbo019rp5KkGyfq0uoyaEpZEx3tP
2a7nr0WDbZmoHtvLbQacs+DTwu/kPEEABlIo3Gi05nePgE3OgkZXp+oNe8u/X680
BcQAsex1EXAdo8t1M0stpemSpPi0EylOECO5aNnAd+oNpIzHKSPFsj7unmEjdHd4
KQoFUBRJuusXmBJhBxMoxyayFBd0GzbyBEpuYN9rOqMw0Ulczl/17peAkFj7rwQ9
kkvGmGJrcikB5Dx3SZCMAi5I81nJU3/UJv+sMi+KKkxDpa4OnHIPq7/hw5yufLir
uRGWQPz95BqeJK9fRA9E94Mlw6oBHd8suAxOLZRtOKpVyE9sas1wugsBBNUm9UHK
ZF1olJvHT+bbJljbcSrsljAIOr+8Hn9AhzeQVvT0Phr25aiBJi1SrZQKSsw26XbD
vOZemXlGqNqeQ63KCdfeNuymZ6IwVpu415t1dFF7l/DebwoECfm6OYT9rmozV/wn
fURvRKILt7GnPg4b3IsmdNgPCgyYBELGpgv+mLYmqZzbJwZc2IYNo+z60sKC4O26
ASpIXHQBtHIySUXZGiKPG0dgfZqj1qskpUpswUCm39KnMoZu0I7RwuTJ2FdEcpY9
ULPRyKMimdjAqQULeFankkEULILacVFETfFh8XOnzGYZZsgltrTeZaBHovaDW7gl
beLvvGyiIbYDpNMA10Gmja06bUvb6cx3TMQeMS3IdHzoIWfSBfHPouYIK/gnc2y6
3m1du9/zbERMLrzU5vJ0Kvil91fBK9VGuOZPFzjGVBlbrlZVjpia+uYV0qL8Yyll
lTBLmPxFwkFMjIRWPgeSo9NKSRKXKDgojYltV/cznR+MgzxeCoK+3TS31VCf4cf+
E/vC4kvii0NzYlnwdSN1/JnsRsgGtN5BWoUNpqbG2FXZsxRB2PFS6hVWNl0t7ycR
hZ+3DUSOGMxHh8Q6A05TRvfsSJgHnom3C8mrUNq814tnN/cFw/SP9DBAOXhnZQMr
AMI0hacd3It8l9hHtiUdJIjWOyftyyJknJ8cSDk/qn2mcus8SB/dd4TMCW8cBAKQ
TZwihkYtWiUmjJzCJwQxg8vJ7a17U4OZWBN2zanHvYGZD7evijKX4GZL6VWDhYZn
QQD7chKcescAySjvlYRfR+PmXzOQv55u716QFbXdC67559yXo6ld4mnM3O279h1S
iuieGnLzd1JBCd8SEUDl+GwJ5zKVneApvbiXnl0Es4Pk1EzLxjWB7vPnn/M4ckU6
rP5w6kzDwcI8roLaHICz1Nd0Mpo2REeIaNoJQcw+/oNnbTb7lZ3CmhR8qxtYDTJ3
SXdHBYH/Sk4S4UZN5uQxfJupL9JlJIGFyF3xhk9N3YAIKLpb/ZqPOUS0cM6VaquP
vw2/xy+cBzE//4KzIo8eeZS/z5RjbYggMJkIXTuE9oJjUs0PnC8q9IoLQB8LryKx
iAl/uIvJYf6jqjoqXzHektWOUh2oPw1pkh22JCLfljplT8JT35eCJyV3MPx+GTCK
Qmul9+K7Q/9/Sui+jfhHP5memMb/XEXg98/2svSEkWSYWc2e4/SKHib7fc1DOORo
U6rSJkDmbqfFMftZwO75axEp/IzU+5EC/FMeq0BU5j1MbCGiP4TJKdI/Y9eps8Bf
ebNikagRBtsYwArAhc9gmoc6Rey77vHRO460plz0IzfAKB3S6ufTO4ZZTtJsFtzG
tNZrL3012h5lCLfdaPA7UTsF0w4+/eITCcug40MS1BWw9iFRsnZC3moqc6OjdzGK
fS812DHX/+AMQqL45DNToqsxIMY+JhCh3LumF9vOlS8HilbCyR3iwF1NAafNI9XP
m4UyIpTJCGfXpkAlilIAo9H9z+ZCmb8Yi91O4kqh8QbDbZ0M2NFHTUiE1/Kh7vGR
dKkQLDDvXb2vL1bJMDe/5po8AGTNxCxwYCNnaa3BpkEPq0eny9E7SQq3hKHVVEYf
2smt36kFzUKi5Y0kdlF7ifUGm7WBMoKL8mqq8W4AeG8hyJjeQomIEeIsBDO+j9bl
noj1Ug/nhuDcN5hgE6UwSuY++UFGs+bspwgsezYB5GmUF3L6UaceZpVVOyz7KnIP
4oEzJutAMAKdXmbEetBJsgMFi6B+Xz8PD4hcZMmAfWXUY+0ZS47cXF795MNwvcwI
uIJKInndr2QcQMRRkxxuLYd0SNiNE6mwLNwgFVKPihBm00fNXeAbZLCd4kyHBCn3
FJ7z0vC4EJqDzPkufL1WpM+FprtTLn7B6a7slS/wcRl+4QV8qyvK5LapXlqL/16Q
kHmaoFWsRmO/YkMeXpVqI7eGAzlZ9bbMS9A9s3y+mxH4VZzWMf3WLqQHFH4xkXdn
210PrAW/v9bSYBoBN8xSskNTQq1JgYnjS0GJszHe7fCnp9C/fp53pLyu10h3CJKe
zADgwvWB1/g9jM+lpONTPluzFIEOMzBOeQ4eHY4jGr8s38M6tL9U3bgunD7Vf/PM
GVipEbeD2GiD8kxQ8esqjw5ROrBfM024BLGsl8AsBz6Md+WGX3g2mbdmfhQlRAxb
ifjDXjtrqK4GLt1m/5zb6ku7KCmyXD1fQWrPWHQbrTkFh/1gG3cp/P4uZO3SHiK8
IUylvMfCOhwvlwdJ57Rf12L8/F6rOI3f64dR3GAm7WPsediZqavOxlhdXnlBWhzl
hjwRFrisd89g0m0NPgIQcQP9qEQyNSzdCHj1JcYebYYMeLOWlhjQEbzgiRDR8j6o
zxmWqjMNUvqzEVy63M6LZJxOyM+H+3wGd+08qs7OFuIqej+Gh02kPQtci3SfMkNW
0z4OwW+f761bq7vs78gcsbm1Yht/JZoOAQInKa+K+IDugjxANMA/atIg2a9SxPly
I/sFcBFAkcSr7Bae2eM0N0dGQNG0xwDvsKvGbBiZcI79Yys01JdXrQMyU0E9uH9t
HWapMt30jfjQN0aO79sIBKG6/xCTO9H8+proMCf4folz29iu3fjFHx/r9+G2zwHi
h7ikabPWk1Ym3klgk/udmJiJHvta72KglxESVgGa/ejBMQz6Csiws+g2c9qnhqNH
soDU+7CgcLG0UU2CN8r/rZm0CaCuW86AT7iiOeLxrTmVcNeBE+GOzEeBG4JLoUcc
Z2JEPu+oNpGBjVqSsJ6v7E27RjnuRAMn7wxRLJVOtJXYvUry9RKrkCaV0xfpg81g
fLuZx8O96yZBtuG6FH+j/RvuKxzeAaFckod60ihLJvKj+9ig3DGM8DfzS9BC+/Bt
TVm8/Wf4RbTvt0VNGbwb+yiacOFAt+KB9zH0RLNNmceZTeddiqr06sd6CxtACuOL
EG+oE88TZ80PGBO2WGwRSPuA9OsLCCLMeEffrkybVp2atjX6Vmpw/C4164LJdjSJ
yEfY2TpywlD2P3wn5mP0TSgvX+x2UEWsvR9Aqt8Ytgr7yvu0jaGe42LvQSyjVGIr
4SeXl7k6vmkKNITpGcMuupJmktcKkqbW4PgMu6oZy3TYLWJGJfPn0A8txmKxmigq
hU28Re1nPf2ALTkYsa+nWMGh8QKetI8NqsqXKF6z5R1MG/8Q7wa/i9etCeumj8LN
xsPzybuDMD0WHCDNoOTIl0Ij6WAcu6RW5jtJETXupEbYhxmeYdn1rIFL1V6ZwzmB
KuZKFYc7kn2f5HEZR7vbtWV1ZK1OFWR4gt/u5pF4Ozj31uyeKx5gPkoQarpl/Tb+
ntqzoR9XNMJxZqJhpt/G6xKbg7MBmHtIx2kTa+98kRiptlWfp//RzXwUS4w+3jiP
cl5TpKrW0fUwj70VR2hEqlM2/YgghL/OyzSY1XcI/ax1nun65XvfK5CHUQD6o8yl
ux1RU17WLrT8lw0sTVR91XLtZhkNjhHXIa92EeF5kKCX/cbaJ+Wsp8vIdUhz4S41
CPcKOTlosJl55hFA723zImiFaaL3eyQNNeyoMUsebI4wSS/kz+Mzgl2f6UVgq7r7
jOUc0/WeoyCxIDbr/lpN5WTnb0NwIdJ8wKSi179K9jAo3L9YVmBo6s5R25rtTFe4
7bea3qRdr3RsL7nfjUDx/bzvUaPRDunOGJNz9FNV8e5eXjUItQX9sXyBRHeHgCM9
aUiNHHzPOo/D5GoRiKgi5ukdl01cWOWmXy6a+2aLFjsVyY90x48n+SjiXzOCABrZ
MuyvirIAX4yux+ZydQmhfz1HcadbbGUYcOcs/AQCmbC7KCfLnsP9oVP+IupB4oAl
cvpvEY+9JTa+3WA07NcXHv6wv5BzCC/Vt/Xyg0qqclCEt1tpgjHO3Z0HJISHSJSm
Hnmp1MJGNphvrh5733p6IPc4CWShK2V52Jc4suNiiQSZ6I1nVikdFpxVp2LOiKCN
ZT6u2wC0wsgto1pHsZGoXwXy2Nv1TVRV4XVlozZMMe++bI+8DQKp++4LuHjjksXX
bk7l3avxEawErKlZiCVkRbz8lz6XSpqaVpGtbHuQ5qocJHQEZn2ALa7/kbhQQzvO
I71iZy3cPezfi8tjJtqShCF4+u8iK081hPhIFUojU1UbJEjXO2YSnxhJ0zRj+R8l
DWIlq69yAJgFHb4TGNhkQj2duiGPzo0h1zsyQdKOVCDOKaacPqJVJM/fjSsYLHqe
ks0D+VRFzABPUfZh1bFjaQiCt6uJUxdLiatmIDKM7rqSK6K4rMX8ZiAeacQ37Bfj
6o80+qcITaSCRW8djswWMpIVn2RQRr/8e7dOZD15k6Rjrg+FAEZGWCgKY9jrKTAB
NhCHCdW5u/R2w/MvnOxe0ILgxApVPY1cOyYinC1L1NJVGulY8Xz0tzHBAdhyN5k8
FtxT2hGdSyMuuW99iqSyirVrTSAbEh/9iaw28mZ2c5ZJKycd1OymQF2QeS0R+pyb
L5OzNEymQNaKOh/nXqErQnaHGELmoSpiWWkjko5RwzvI3agugVIgCE8c7662WS7f
S6pHnw2OcFrZf1u6zqJLhO3yuER5hCd+HKUeVZbA/wLa4B/ygkCeKTCBG0pd7nPP
AUmyFJWv7pTcvPhdatUQCEduOZLuXBARRsQT6u1lVchCcAw9dg8MG6vvOuiJYU+r
+Qf/tiG8oILlshUTfla4viJx/MBeTaMWpuctXAJYj3Udqvmtqo7P8pA9HN07emmy
IMwzcrJWUAbodwzjO+/xFfQfODadRRR/5HDELTzYrGkwju0zrtdeF7ZzfPNJhmfl
+4Yk67QhR2D2bMyovaNryj4GpjJeu/OHG0ogLf76JTRaxAVKLhdpxUWAdA9WY14Q
+8wK7qHFrpAAKh+jDOWQrSrXytFmou+pDQdqoM2hmtonfgNEz7HlIm3cf2N8WcWK
mHjqjr8OKDud55xTpqVOPc+LC680dQaY3aAtwshAkwNLDbtCQJDUBvfepzta//9T
/2GZirfuxaj3YQIH3BlaYVi9u+xUn0TIlhtVKlF+QTFpJmKEwQbwmgkI44ts/c9D
qfmbI6CtiMnsFD67x360ccEE56TGeOHkYaUu2EtXrCMCthruozANpJo0JZEAOjYX
ilvlXSQfT6wewDf8210Vhe7fZlVtnMQDNMFJDXAVzfFwczs30x+WNAyT56K6G1BE
yPmvvboxkPS8IsSdRiWS+PNu8j69at1BMZW1FebjnUobEc3Wsv/F+kXNyood6JYh
Jt8Yvu8zZpYDfkAL8QyyeV/fbD1Zuol6qABUFI2a2gh2hjaXewhw5GU3RpHYaXIA
I9Nm4PxKMRZ6hIfKgb/Punv1J6tO+7x6yR890/KOCs6g5yKWb9IcYazNztmd6PhS
hP1bw1YCQhPfOj+MIRkqszJ4agsKE+/ZYbw5Lh4ql9H7cmm1LNzcqBccKfsURJ5B
RY7iOS+Jd9zEChPPE4jfjaM+OkeoVZpOAggQXa9JUxfydD0zDDfoMLGa745f7kRF
OMohG2dHGKsaqw3na2G5lCagQL8axx3oqvoKYtRzWWEwcsyrIcTrMEsTW8PWNebw
noyw9jYcvqNdTig/kSVlsnIzWE1i7jlWeixS/uWI5XZYReFEGnFL3QsIQCO97KiX
yDWSz6kM22bF5kSGQHDixklDEi/Yq9dMTfwKq/lMD9Dm5nBgeLeb1PwnN4IhoQ3u
9UHW2z6LpVTozF2Yw2ktFabrQTFpbyK2TlM99VBivq0g/YJC7uIswpLhfv+rg1kr
U9Xb0sWOevo6Xmosv7lms5tAxHIhRXAsNtU84fEP9C0LY7Pge2c2aut+662wjsS+
4AG4TOksDuuwQ9rz1tKyuEt4VtW7RMiCYsdkDApyCWlWsDB20V77RtRF3LojXRaO
i3ZnzjNNXrAEwlV9mC9MWOU93887d1+tEhrhJkmXa+BXEJxNK1mKzQW2D9aJBJzv
UdALc6Fkyxx+o465oP1E5+EyIkh3YvnRXgh2foxx+2XR7z624QjFGt2gsAw16J0d
+9bpgmqZZrMy4rMO4+UWjSjytM1nwOHHMB/Ow4YJb/XsE7WJ9grHiDEOW4SdZWXu
7VfVfgv0aUHlP8wUXQIkqNlbbaMpan9KZVuYWzTc0KFgleDsPC4fOYYO82b6vGG5
sYLjphvZWYxCJj50jpgsu97+h7hV1vwUl0UNd54nsKoZrrTgFnOKbrf/7z0m1D5W
R+jHwOPkCGpAoPMYMMv/51lmqbyZ65qMS+21k6SEI2w0nCFKPGik8GggOLp6X27y
dYO+laAvgfydhe45dlWysL+sFB0/tG1h+BtX9MhPKn2siFtl7PrRk25vL8VzTi4e
kQD4VLUjmGkvNNUHjX6MQQFJDO6Zc6tlJYteGBd+qPMTAa8y9cLiRgS1OnNAT4c3
TnjvL72AFNw0UNvMUmC5JjgHL/nB+569RNfJjKTEQstQuEFvsjgrAPThyBRC/B+J
1mLEaNq7cHsxLBEoTA3XRSbUz8h+QusrNpyE/uIDicsYeHdDY4HKtJM+mRITlLoW
ePEdIUvBMzci32adY5+ghjfctzLA1oxhC06Kh0Yirwt65/lH7CCSNIuEEbDjDDIi
KhF3fhK/KkmIdngzetpmEIR2eLgNMJwZxjfyJGOk+I0TM8X0SLb3jco1i+Uzey5N
+SZ8qmNR77DhtynGE1imv6PbNOpUGhOzg6BabWDOlxrEE/7HO2N6dTOuyPkdwFV3
i36vcocmeqT/SeorRnlCUQEkOivwhH8MRfgdIpzqPoJExWv6LqelaJKEnc2HgcM/
PSAIppJDtV5mIB8Octl8oa9Ab27Lclhay8JPxiElofcbDiEjgvjoOU+J8iLL/ShZ
4EEzqHbww/nfdxcwu4kPHpmU8a04DBG8LhtQvK6p8kkv089JDlqxvoeAVFjQ9h6/
Vh7VyCGW5Uu5VWARCXGMMYuPrQHCOTHD8b5GBG9xwmcSh11hiJMMXKK/juQwS3gt
vph4RV73hl9ihqqFbFFjI0kgLa2rR6SaE9wjuncXyI+6K6/wgvL+AnivP5LRVsSa
KHhrHUPuN6MQcXBvcpeWTMa0W0kXw+vFMGQ0zuw3i4eCQpHldrZ0XQLwNZLL/O1C
bugHrTAwxnObjE5u+fYpMoxkggI7vknqXoc8WTmRXrxhpT5v0cVS0tZa5gHOjLeE
jLwonC0tm4855mU1SFxvzWwDCWOgyKkx2kyi0P1aVhkhOY3Sc47dn/7kXktRFh7p
h6FkGMEUDek0xgl/phH3uAP20tgdBLlRpGiwxnhar9aNsiKhBwu+bi7i7CvCXe16
qcN8f0AwGRAfWmcmksmzW01IgEl75d5j9EfV7M5WpXfQ41mw4ovb/sAFOO395488
C1QFd8gstVdviqKUst2/qF6SlAvPzHmF/MGpRzLCg18FzuxRj6j5z+JcGyt95lLr
lIcWbmIWEc0RZSkhhPpmpFfy/GHIBQepdHddiKLEBY7x8KjkANTC96ZBxVL8tKX3
OyrmmtuskAijp3bWfYn9tmEYocPdZA/vJjbwSX0i15nDgsM1QKkEGELgdsNSP/OL
fWlbq0SiJXLCvRgZLh83J50J1OsxumVNz3Gkt6c9RAZYXzQ56QuMNnNgEZ2hnQuB
/NwumOydEJvNNgM9EFStXk+wXdWlwVKK9k/Az9FuC4Adbn7zfFoBOVnWQ9VZt+FY
NrI4bGcMXtQRYbzRQUTKmHQE5jMZWJjpCRUW6vfgBXibbUYh/H6RRzLgbaR5bQ2I
mt7TQVgTAMTyUB3e65FbzGNtwx5+8fOI99zzqUrQ0s5IW+S0BhGe2+R3eT16bvtc
lSlsMtTPcDHKCry18v2Er6ITHWk7yyyiCtQRNOzqyNonXmFQtmBa27S4JSBwouEL
EmA1sttJIHPTf1PncT4ESceb+2seiWIgjV1POeL0YnDW9LNaRL+waBOyGaLXnuxA
L4kWMx27qDt+bcbMh+HsmA2yOD9FTHGAuJYkqVnvcELkb7B9kBzoBHosGMLUpi5Y
s+SLuNsEFCa7YEGE4p4d1rI0kLWiA5AT6Ak9NKzOlBArXjpF0VOFUKwZyo7u6bNS
fzDGrTph11kKpyVtBwTaQn4jwh8Otb6mO7ZPA8vIAafEWOnWHETzl00QVkY+TpCp
dc+GCekNywsNfEdVF6BmJjbvMBPOnDTD4TbRHO0QqVrTxPG/N1myn7Edx8OXF9hf
9PXpNgRakFWNfTTMgmgihzd1YI7Zgqf+bE0YzpXoKKltOIasvq9zGXvh+UriEwdY
buSK/errfjlBsRyxDlF71frRH7VBGEM6zj0Tg7d0Sikwj/rdaed1DHudQZ9m8zG3
OherZKmRI1xKYhZBn+3r7Um4V4iTKTk1C0hCkFxeZ3JbW2r0Vl938gqOA4GCJV3+
uxXiakQ3m5HRCv/qvkv3b8C0RNaGzr9a55PSrh5nWuup9V1RcSP9eNZ3/d3gBJa2
aWAI92Me51vYmUiKOwuyRKmj09mdHtsJepN/d5DL/HcEoA0MuDwzA356MmYSV7oG
ClZADJmF7Ay9N6xw92c8172hSKJacnpUqSWCW/0NDHnOkbFP+9yfI/a38ANwSTSt
+zDRbU9NCIQugbgEqCLKhhQ2HVMGceAHfXmFdr1Ow0A9jQ5FYPumohUwWp4KoxCb
5w0l8fwaDIkDj4Tn+YGCPWOpGtbQHjMvkOkJ1eW1HfpSQiYNNjxRAilxQIxQ1zFY
mvHR4TrZ95G0Wj+4bE1CdhZRprNHLS+qS/3904nQG/6ydXaW+g8WZ7ejKD5hOFS/
ssQv/MtLi+6YAXutrZukdXpzUDsTJ2ILqfWHKeY0pjC4uIB/HZfSGMxuDdYZGEG9
lwD0Ju+EBf13kOSeQ1oyCUQEyhflJ04zUfkURkeryE8YuATsvIX3LhTkiQyuOYdv
HjIoLgP34D7YHl1Hm+4k2RTCPHQI75hbPBaUcqpJdqUA41k7rcL5HL4SZH5P3wHd
UDB1M2B6GOGXQNdgQ0vu1kQg8p20XLWC8bcogFzDniy0iF1KEwkYgYO1sBTVJCSa
ybSm2ydQEuE+XtzIktrm3NO4ZSjyhv/8aSSIJMUnphhvZ9POS/fMCngLPsQpM63f
TGaqPUAhsN5dNTl67TUaDwzvZviMK2j+FbaNPcdZp/Su2Od+urGT/gV8EMrFAgoK
+nZcjMcyBF7ApYvs0Kcin2PTtrMWxhjfIxN/gaB6SvACsD/hYEgLypDUawNCoM7L
EVzIvRo21tl2AUJI/67BVwsTu8waHQVbakCJjYp3ut53YzOSqqrWXy2rBZ/yxRkN
sNA2fLipUQZjpAbs9xMCWS2gkw9ebzEbsxRGDPcJjg1iA3QmdBE6OcNH1g5niEWM
a6xdgSPeCfPpcovxQIq5HqYm5KMMzlK60OP8CC/5R6howUnmETCxlHksCJIUguhP
6u8LaLwbWyJDXZjlnTzVfB4q/a1/dCTIDJzJNRToX9TzNPxls42GLElaDY1Bl12G
3Zelr/du9y1XyuVoxpJjsufyQd2BvgAKdg5UtJ9BGulz2FdpF47WFF+yEK6NfZEP
nHL+gcKwA0NHG4/zu4rWaHvFO22jt1Cpy3dzfhLnO6iiq83CDDVD+WZFr9RYW8tf
E+PJ7l7dvwXi1M9vEA5T38wN/yadRQV5yrcW1NE8CJ9SoALjJVqBxSHmvmpyPzOV
iSQL8re9mPFGVmzotLNlgZxM8wHcyErokHrCq0LvKhLj1+Vs3N0Pn7co4QA0joio
UCktNIClcJEga4Rsw8aF5mDhPzurIHtpDaWdIjTBKn6vQM9pqNDW4mpDnCNmQEIF
LOS0QZGTx7Do+pNZOp0WMvd9Cx8TlimJ5WiH5IKMgXdYR7gr1ye1fYos4qsxjI2a
qVdFkaMRhV6OLlyzaaIWG9BupkxvJ6nN8hj5IR6qTEFr+SuukADl6gpQXMMXrd7m
/VWa3mgvPQjlefgRoYwKZHuqoFuq/F9PJa61Mgkj5J5e0xot0lol5A+tsP7nUU8X
13WhtTfV6rC2fqejqfY7/FxM48V6xgUYtq77A0F5scN4GhhA/52y36PReJSK6u/e
Q9/c3oDG7KoEi3+5LEzNKyK0fJyCCQK4CzeLvsgKBZ615zZqmCkchNzQ12qd9An/
qPC7fRfE0S9DBxk0wkoE9z93yC8tJ3PjsG1GJe90at5jrWrXiGx6X0GyGCyhD7//
N3SCvjiLL93I40BUJh6hd8nsJstBZabhuXzI6e+csX6NOSQnmDxwcmevkNPRIeOL
2SX3xH0fptMi7gyUxltoIAHFX8Wun0bjo4MHovhym7ISuxJ7qK8ozmg/6QUxOEt7
Vlam5irARVpi1S5w6BXaLYirlcJGrkmEsG0OLf1R6FGU7HbMY6hiEBVNk3IqLLKR
o8/2zaewfnGF2kTtv3lK5KpkbHMB0OScU/4Kv6lXAiTOsBbC2NNj9CmN54xWbakG
pyofM7UtBgyo2eolW559KyJVpKckgCxdk4S0fZwjJ4BFVvbRd7y9gcfIRJgzZ5Jq
7hY0l6gHb2VZIRjziKxNlNzcrse+ns+fjA3wwJP8sn69/VVB2fXA68nSYPZHuSjN
0BYJ7BCHn9A4Iyeao7vF53GCcwM/0UmAvNUWZIKJKVdgqO4Ig+SiHnDnn6w3iaY+
gKa8j9EDQAMSJsv1KZIc21flCB2FR3FUMAZg2czANmAClfaqJl5uL0qH+O8GTOby
zTKCpNZoy9Mv7MxxDU/Kg64bbX3/1s+GUGB0qKQHF+scEMVrAGh1wgy35cb/IEq4
5gwawunuuNHw01rjiTupu35W/Z8KidmaRuf/lmhRIJJxhk849Nqlt4JhfbqTNs9D
REPCuX2Tzauz6ToxkXou+PM4MCN8yNWieQXQ8rm/zIvaub72qG5lW3wvXKQVJERe
XfSfbaxiPIu/pajfTEmB8f/fmouCSGrQrM7Hft8yBQLWwgJHP4EoP8spTuxzoer3
j1Kat1SmeUCVgGfqcb2/tj2YVa0ofdFhyhxwJjERQlKMQxu0HdytQ8iA/RJE9cCB
b2Ug51dn0/x8BmWxm1oiPxxBb5plEBRYKHGlNfoH7xjVr4E2YllGsG1F09jdz75t
zgoKD1Y+bMclH/II4FSJ5jv2KuWi+kr4CTRvFxJ46KNfebftYk7fAxlj4Vp1l372
zAcZ/dma6+a+oIIaN0xFsd2yx+yDAJjPLwza6lleRxv0w6zg4bnzAa2b8c+K3yLV
T88rx4pZaffXKox5/AMlyKbDXoB57RQD+vdWHxDsf6d9K3Itvz7vB5gMPxvAR5PZ
pl5vjUzMXvOrnIu7tIZzypbZZHJZp8uN8OdOTR7nNn0caqQ0z41gwYHVxLGrbA+z
qcKPVFRg6ewhfMScqxiy18j6lU3zjwbur68Dpe+n6+YFT+cBiraw5LwTIsOLleJ/
7aXDVE2uIjRZvzltKNoOWUZ2+d82i8b88LBrC7cGZffwCrGYZLxi+o1/tese/lkp
K9v+nVZLKJJKNumIdahhrI6hXjr5f0mX6enEtTc7bGZHbhwDsRcvwh2n7hmImt0C
BDtywfvwZ5ZOQBdi2oidR4AOtUYNqCSVwG3V3jLdtJfrkV184d8xTrJlGPw43yVe
aYr1+9OMJlV7kvQWp8SgWDgQUfPIvfzkB4ZlT3HSPblDM1ZZLurpL+gm4KA1RKmx
SGxljwTL8DS/t0BznXVsFtshjP1YKRuF1SQMcznMh+EjSaT5QC7SDkwViaTl5ifj
tzkzfw8my8NjqM0tINvfBi2XKWtKTGe0ws42QdcaM1qRgI10PIF0Bw0ks0j8Lhll
/riSlmuSn3XZkP1pgeljPI+8wuFifiskZTCo40JTkur/F2iE2XZlnrThxcxl4kGd
Pd+JplO9kX16ang/t3HRhYsUKIpgXtxUVsQyvVJ6Iz3doMZG6ADBswwuBzlWuRSJ
FIFSF2XujW5vEslyO+booMtamNTi5c8LRI+P1kxjmiGryWI8cKW50BFcQi4Z2aJ3
NhF5Ip17R1I9LvY/T5bkBqiZFiAZQ4gKz4tD+N1TiaBm+R3AxZC+mYZvogpc6eEH
HzToH7OBvsSk0EGUZMcclbZ7FXbxdNZlLvc4llE5U4FMvmNEGZpwIgrgwLDsfzNz
Y0IpHiMkuaF3pGgk1l583zL06/RGBapInOrxLhk6y90yvn/iHUYyidhaSlAQXXYL
n0cxC5TxVN8X5Zkcu6P/B33a0fDXDAA/6NgAbGBkEfO5iTgF7a/n/3Z8FsUFtPWS
XcvcJnOQmGKDxQaLt+f0Vt5ljGYG2NfR/K01twizgV8cidwQudU5ZLcf/iF4RHs4
06XCMhD9a9OIJ8gkRUJ7V9MP6rxWwPuVycvox+CrTfzaTeU2IAXMCDkG3+0To+zX
JKp5T9wCDojiv51C4rUvKXhRlqAFSkIs3yG0O96qSBTYOi3rgbfo0vJf+R2ETxr6
752e4Acqp/ixF7+Ly7C9ID4SQzj34ZfBy8xHugnENvzyVV5TL7xKtlyztNWGNLhI
9etxWgxCjA1I/r5fMg67UvazN2Ayt61P1fB/JxV1T35DxzXo9tbraqOO4RfMST/o
7OionJUns+COiF+2KdmmJdg189LE9aVs3tHdBCkOS68aRqRbBLjYUT/CX91ciS8K
V522KXIGiia3MxnVOy44Oz4Zyh5TO9qS1GjtU0f+rLay81uBBCQHMzEJ8WEHIS+a
oEnusIJE4UuRgpbpN83AU0brs4b7LBlVp0/gwFZkDTyx7DVbJ+S9q/fIOkHXtstk
W5sUufDUorBwzSPTROJ0t9vlpe6EPBcm7rAQj/T8RZlM4c/i7sR8S7V1UpFAi2ol
HDXhI072fEVmBQhdpTzOweLN2RyxAgiZVm3iDDAcLvEuJg0JO8gF3exzENXWWTrF
fAkB3jx0SmpiYpGd1PKq4/pRs0SlJU/rkJBTCgLjbvzfT903Xe7hjcxycz+1DLGc
EhG48dIZCHLvNEU5mCnV90f0bpwX6AQD2/x1pSIuK8QHAkJKj0qkaej6bGC+L/IM
Y5co+4WOPtE8IbD1WuVvdZlYsMSg5guK4HhkwZ6ONplfiTh2vOI23JhQG8p/nfyB
JbySTPp5CTIUzn99H1QKPZC+HLxpvRgym5yWbQtkyhFsS0xEqyWVRlklCM3CswCR
YPjnnZ/PM/3U9rbs1+jV0mAjZZ78GUGQEf60v5jERNjCVyRB96jZqneTZ5tROt7x
oFDy5pmttWH6IXz+cQNB8KlM2HF6xqi1RAUWSUmkkGxM4u1ZTj2m4GmX2BVrCsT9
A9TVuO8yxZxpAinPSXZWrBA+U5cb5aBZf2tz0H4Ag671crf/d0oPWKdXvp3Ixd7O
yvhv5SjzBLx1YYvqZAb9Aksn2AC4cKmDC0XGxwQl+Ex4u15VjmfR73oCquzeEJRv
cTGSa6uN6RIiUra7hKD5JgLd9pUPijG6UKQTlsRT1rhW6vtB2Oojk8JzOaLZ7vKa
RPSSnws45PhYO/IGpxFsKIxwjCCUlgevRuZr13biLtrHBleHIks7V9VQQ6k9Q71l
VoNO5LF/bXU/x9JAuzKE1aeFjRThcHuOTxfL/IDNv8uFW1GJdZrOiZyBtcalZ+LI
xk8DHPc4Mpbls3i1qOiyPwk2Bqj2xsQ7Q4R+qC8Zka1M/ef58W/RIQcLVu7tTLOd
v2DX7r2WRkjDMfe3Jn97nXprQcehXJX1HiENWJ55rl6hP3ZsgoI9UpNuPcWdAB7c
Bi78AYnPuqXD086IMhTx6D9xhOaDakPEotCOhXx7j/9XEnbSINKDKMoGl32iXEOB
jUhb9HlszMIv3SERHtK1Yxc6eC6E0XQ9yNDhNjZ4kTjpOmnGU5ytKfcVb3D3Nqn+
uHQuFQCLmtnZBtE/tW0RF+7BcQrx56j3R5iRE+bUcO6m1gGF7Ls1XD9zDeyMRIvt
iZaTvWxwjPXGvNgCG2DawDZGwOZuP0Wxe/p2+SNudz9U/S7s/haKxkd40qBThfWt
fXuTMnMvw8gO/sarBDMa3ia6CbUdNFnY8lxHgweE+F7h3hfXq3n1TeAOrDzSsI6F
jorFCkfeo3PV2NmVL5UjAIBoWrf/OEqRPnlfLFLbvW//E0PBkQJWLhzMW/PJjyJ8
nJmeVs2RUoWRtN+38WN4O2sv5hBUetfx+QlG+cW5WnuaPJxw8eNJs8YOxkEruwV3
VSQnUyEpiF2X9+Ig0ISg401mCoTqnqeat3E+1dZXEcdVlRA5QnGOA7H4d8IsFpF2
Hfi8l3nnHtvrCwGVY4bkSmzaX75Pv8k8KmAWna4TMu2/PlE9a0WvuSGbW4sYSFu9
KJGpNdclxB9WdxZRh6yOtYL+gEui5jIDHiThk3/JHqwAXDJ7rKVGHcQhxiihWunI
Lj7JjPvTnqM557tgju1mPeMfAzhCGbxVR5LIDLerIFHSO9eeR1Hj7S5/BgJ2a8tZ
8ij2/UHIHjcKcSYzfkvE4Vp0Vot9tv8eM4iQhlMSrq1hiyblrys6/cO+xyKJ2XXG
vcCUTvORXWV4N7vtoMsFdt/xivt6Rxzm2yJgeB+CoGcKmK5Yx9S725Vd8MjKWbgg
uUJ3XldTAuqLmSlLCe5eBsKsoFgOdMompV5pdanwDqvIegVGI9Sv743lag8lYjV6
QyMhU1CwGAUfO1g1w8/48vQbstVtADOU9dF5bXT6s34B5PLswzRVk/gdYaj5OBlz
/XhgoRxLdAr/j30C/ZUk+a0P7yQyBQcNYrVUM2EAt01Jjt3jp43m6tlCy5d9NUvs
NDtQDlFCtHAqzQ9zGTlfXKmUw1E1DrNT3TLRxCnwULo00jMjkl+NPXNrc2jg6xhz
K6CRHIUg2dFEvT8XFnBQJ7TXLFOSM7GUjTw0c0aA6FtyIPGofXR/GYnysW5MVUPz
zMk298P4m7F3m90pgM03E224FbJqX1oa32xHy0vPgwb6FWUktHUNb8D61E6v2Sq8
XV4bYJDSOWw8TVW5F88OBFOk11eERBSl7gpZR/3fx6/K+fhGSBRZS/CqLJ6aeqMV
L6nyJO1+Bm2AwuTLLnMLNRQPb/8g3OuceGzLZEIuT78G3r6CfJqgURjPTo/kYkiW
6Ly1DUfCoDOMHTwQtWTapuKwxd+VQDyvnm5ilPxodCL2qDXUwU7L299EWSbqiq9o
kfi+j6OHh6RP2ekTmBQPlJwN6JbUBHnLg0jQe1wAJQnhreR9kyl3IcMD7/eaUEsG
LOrouuU8SBkTdJCiihpGsyiKAOHZWrUmkhi3jbMnS9KalDHoxWNFeuua5F+/gmCw
AzZGuTPTVu1S8CgyVSaCR40TWwAP8CE6uFnUZFocVn2RuvAC2tlbqx59XaFj/9Rv
jEoLVDM0O81Y8Ebn8DMd0FCcQSofHn0Dz7+RGbN/z56WQhHhtRgwuJZNPY/p/9BU
A576c6G2l8eEXo/QkHNekn0HwOOHJF5hi7ZIsKyfBwF5dPAlZUVZ2h+fi1TU8xPs
LcK4yqjUmSVQOEvAWWTaLIjTD/gnEaDdv54vCcP2uZ0WyDXmIJjxf+iIMacnLY7b
o58vW6YX/w8AfBfccqEQ0lrKTvSK1ubSJJVZVGi1Uva03wQGWqT/Utc9mEAq2ye0
DVnIdOF7FDsaKsDAVSmuLEloPyyPV1GYngKCpkGuXSvS45jppnSM5GaoV5pm7i1J
DHYTUN8euz5P6dzRVlIuDmPRBHwPGFVetez0MWZJYwopw1PQIfg8Hs3HVSTd/jHj
tMcEo7fKaMDZNOEn1Dls4Zk9lYklX/RgXgLLM5rzz79YuHFLH83MO2gInNvfaZRj
YKqDaV4D0JajriUJ/KUVvHILbRzodmCnfDWzFLqoaHknkq6gROpXyw6ybRaTmn6C
mPQc1VOt/4e7x2sUW4GSmfrv94sR2kLJFbcNIeufGOuATBg0B22OKMljDdWh/gAg
+ZY0dlMMy/YmQBlvY3Kc0ND6jc9ioUxN0oZ/mvLVmQfKaMwIf2w6MOQOHMBQ0zJu
Pd/B3nv+y+Ba6MbtoYahSoHip+GZd8XKvTBu5e6KPplkX9po30+cCc36WVSo4uSt
K+z71Id1ti1nUbTHFQxnuV0bNWy7UKIjIVgywTZ/6jseiEyQzkltqV5qT1dVe8TF
DXC5eWT8eSSHfOreihDFTouucC/ZCn5gCXx+C8J8UqD0bT8+0mrRpa59HoA2rJHT
q19aZVpYuMIMF7e7XDClH1UdEtbEhCyhs7/F63t3sa3dSl1wjw/BxXmRnwK1cl/M
dp/B95iJymlzT33eG7p+e8SqR/sjBTZv25Pq9l78Z756HRCLrf3ul2yDNH/fbtN8
bTcoQX1kGFueLvxGS4QudDI+mq8Lxrjosa789ervOaxEOWksQVkjKbgQr6DVFq+F
egNskPxW44t4l7Jqz5iWOEyavaYg36shSbVCnL2OLTOl5pQVH3YKumgltgycFjFf
EVhP4zvBB1y5VpPTdHnhm8pZ4p5A78sfnJXW41e8QLGIKuoXRLYllJNSwrQEpNYy
jh8IiWWOpLE1URJZ/J9q4SZ/8V35CViLZqjaI9Av1OZTTxI0rol6r3aYEDjKt4ce
XyquQQi4qpz86tPE+fyaB/gtMzI83Un5BycOk/44kefr4m+/wzil67uBwbngbNdN
3iAZNSc9AglpsS47w5v+9c3hDufcLB3sVAHKOGBJJjNSj5vV920iJ8ABrsN+E6yi
XnKx6ArlS+SiSeGBZ5HKg1Sz63KQDIFrOyscAbkVb/6LswXcgShNyLvYdP7k+2yE
umOVpDoy8N6/W8aJvx+Shw11mvTm5SYMxmRpAcQrNX85NpcsEfcZkGHE/WckEYRY
5aHUsJ0SqowgYCz8oELUKJD82aslBKm2JIFihYFkkhFcXlnIaTTOXmEdKGJaO09w
IjrgpFvBEgvIVHfA8+PPNNMbzRAtKE/hJIjbnUq9CdwHn+OERLKtt5Z2rdlY9W12
NybNDFEMFpsqcxRla54hF0rODqfyt8f/RnkjXf6QSBp2mT7TVaaZmD34Ogbqtkhi
pGpRfgs7wJRwmWAwTOFb3ZQdENP6rVH1Hf3jEHTFOePS2L1an/gmkzTbnTw9VebP
+uE3u8eTQKTvsacu6M6YWscpILJem7DB/IlgqT5pIknFh+RzrmJZeg/tw242c8qg
ezgQtNGlp24kw87Z9nHlZZ0JI58v1qAer+0VAUhkk0bo2o7J4Q3YETyddhav7Wq/
DQF71/GplFfvO0pX+M2K2rsnGE2DkgdW22+aiHxE8DeomfMiwlJFAID0rdu1KmGh
ZppUZ8ypirELo8aYZSP5nKXEDuscEYqtLlIrN+s8u7K/Ym0To/qxACw37Stroiro
90puXiINsS/hTjuMd7+V1VyBZYlR5S+ZMwR0fHIT9iSlt2PTQbwS5sjav+M6OZWd
pLRm71LDWHl5fBJm1pMkZCcobFXq+DrOIxGc7UGbGN1gFLQIpf0ZaZMd2IH6k3gw
3VfrlzgeC5nnlg+xnXn3Lx8zDBq682xb+YzYSg+fdh0nsm3nKtKPwbvyolXA5CVw
qGlfjZXVHbl8f4ftq0tU019a+hvfPP7Ih7wQSkzUpbmeOTjeMfO64+fChSQYZh8Z
Gn9XwCrhw1V5IhGAGlxxQCoCTflDFmBQEB83qD+lr2b/81PMAH915BRRbm+i7VBK
N2gPyJ5PR78WSJKZSAiEIFQJrdB3EvRilk3ykWQy7Vm8KzfZZ6hLn9LNAKc16QsF
yLsBoXWDly6ocD239xI1LibHgCH6Dp2fZXV1XC9Ohq8SC7o0wXoYhrHHufziAQjW
FyTg7mwb3PzNk4ju7TVr/pT9imxvZzGll4EKnVEiGBQszLvt9XDL7QUtWorXb7Dp
bGPhL+zN7jFBgPmo3CWMA09j53jWFUvst0ptxyWsTevy28V5s8gvRfe//TwT9Kmp
PvCcpdv0LnCR3kphPtCgtykh8w1I2XhsDXtaG0RMAfDjCmIraoZJ+UYQfiozvzS8
cBNqRNw5sdhcwajogfznFUeqSHKJyvtU4wdqCxStFixrjWRk4UCu8nFaghX0zObc
le2vFdmyef998E7fBT1dl4pnBar0z4d+SId38yQ2Jq7NlA4JO910w3PQrKUM+Fxf
nNKpEyHFWN4zzJKJpdcj9rRIcXBkRDxkjwBCUkplBR6vRjQsjjsX+XMZvkDIhQGW
29RHfFu+0n5fbcJ3qnKwdgPq+66dziEUy91luM+ogR0KU7SXQqX/0O/KG9IlobfM
wEqqjyFkL4N16G47D1YuNY7CH5e9oEGohJV48RQCqIJX2Xv+6DgW+yJai1B9aqbn
tk1UJ06b3LtcoZ0MoWw4IrvOGb/qSr+ZdhGsdXSD1GxK6OC5SpsWPsQ32g7mHEMw
y+S4zDpg8VnVZcGOPGmXMmeKkvDu0oI7WVOlyFKA0pHD3l4rbxrVGPT3AhHGBYfD
kFQuIcwJsqQjFtKv9soMi8/OuXqgzMOpUZUvpsMaU8u7UUZN8X6etZd31lk8lqqh
Ipr2Nw7ZW+HwdyJI7zBJcN4FfzYLrr8HlaVNDhnYF/Rt/x9cxvXZiHjYTeg0fFH8
NL0cbLG+v3j+Oa58m/Abtr7Us5RIg5eivsSyw90VInhzt3k5m2jmn+SbYRmKHE5o
wCvwp7dObdM2VWuDT4iA+tK9bokphE84p/KJYKIYPeUngRHqujoKelaXR/Qd8LnY
ytda8yeePqr/JOss6EpbboVj3pRFeGeHcG4osdeSXrljqowim6ZnkWwWxEzHdhc2
6p+KHziYaFbR+fLioXYDLHIJ4KLpkhvI0n9VSIR5WhVyvcLeVWRRr4JfVs6G9pBa
guzumWvaVCHzyYAIwu6z7tjmcgpkfgE/hOnjl5nGGoFnzr8cK/ZGR9fq+VAWrwdA
8UQaAjFp0Eaym1XUfmY3PbJ8N/+PntCd+0A4omRkWjRlSN1bEZm4xHYkJtTgDQCa
Hj+Px+xI5iPtZpx4Uy03KxC68jDwOhJnK4nco15nFg+E8zUuU6yRNiVOx8qOXLJY
ZbNBgwWlu9w92SxdD/0xHcZ/aJHnuEef4ModrSGbzuA8c83My2oa+ffJW4tOgjfY
pPuKWssQbQr1ppDj4N/T1xNFfee6J/Ha5/yv7O0GV5CNpp5aYjavtSR2Ff0Mhosq
TXQzyQJUu73PtAz0iCYTSIBLXxjXjrFWGzlyv78ZO4aUlO/gwW62GkelRI6su8Jz
clenqyLQTeisn3/MIHbualgSZkvSQjGaJ90kpexosmeutR/FU0FQJVlemr1Z6gft
YmZ7fm2G8rGTop5qdp469cU50K0loM0NTeE3XZtKUX2OHPbd2nJoYpatgyx5xG9d
rymkUeQ1JRjtI09zSX7COKcRQH2YLvdXMIR27ZZCXFG7pJLNzga9+0YtfUV3zeNF
RbAzbhqWQ6u5JJ7d9mkg10Sh9lyVAzaYFTFWYj9EWqb2JvdNFldaKDrI7E1ZbS3e
VIzTfdUHFb1evU8wpIH7q1+Tvpwmw9SnF606L8Vw/8sud84LeyZ6IqAdCyPKiPUS
xBxO4szk9YPvpfvjXUjaFMoYvKCgGFMpeBrGSdXpL1Ljo+UowUJNuFrOaO7R+rcS
QVcJ8MzQ8bQVR7OLhcCHwEnOTZxwYN5fvCWQW66vibGU5r2hR+O593nH9OTFQC4a
2ZizAFJI2wbdMXfx/sjSnEUd/1PILlRaFmultkIRnj5t9nZrVjUSoQEiqjtUPb3H
0o4YxnJSB6UK/kbhteMGXJdqCrEJsS8rLSmIl7rKFYXsuICyGKNdMv+IO6chH7Ky
o1SJLdhSi4AGgIaCkDhWw2y12O7EQ1wS9c6ZZoXQqj8JjF10MCtRImbvrpJKHLev
nFaqqKtmG7LOceX4u8K6RZWv31Y8E1kqB17wHe6pVdeBE6iczgygoIC748832ePh
esuDQG+RR5egLbDvF0as0O+r7jV0cdpqOviQOzrPa8rxUvYY2/qQWaIrWobD8HJ5
jJoYOnOTS25p2DbhY87SeLe6NCE07WOskKImmobdsFRtg/jtB5h9CgSotd6Dc0hp
jydgR+YJTvAW8YK9tsqx64h/GBE1cpSrKC7uaGqRmlWhg5rSlit97gQDik2z6qlI
LTvYiJNXVPXD7y7hcPRpiOZ1KjIMaolbso9A11x+9D4woUhhX6hqEoaFD0GzOK0E
fXHf5vx86w3dFlrNBR161cfQbA8VVX/8oVyeKcbKDsARe9UF/5a6P7t0EPO42Yhl
ZFx4wUwvr8IsFsGcSyoFzQ9CN8LzFFdDKLpJD+d7bj2pJjseSG/k0+pzu1cjkZ0f
GCww719C9hyLj9TdJJMAI2JHNaKM2F5JXHJBw141vY5rSiF8Ex8VoSAvUrtgi5Uk
6hMRdBKG7EgvanOrxYL3ovHj0YSt4FgHs1pMg+wlsQrhg8uz/XjMrY7e39db1l9W
VW8QBvS891K4MysmpYRJGvilvZ1FpQ2rGHo2j+wcakzrQzjvme+ejVJiE2f+AimA
FyZI+M8filolyRKTaMErp476x79mTIdNlqEY1Z0ciuFV6ypfrtGn2t630+0ZFuqB
Yq3HrtbPpm3SdlHbQCBXIbFqphmRMmeanhmfXQZXLZBF8BtkH1wZH+nofsHm4lyZ
bxxAfmsDlF4V0ynYcGdFrqRcdBOpbljSGXp5HkCJ7bYWQtz1hHNXyo7fBLXOyJEZ
975VWt0zDdL4GY+xDjhOn5Y26M2Wrka/pnUGAAeHWdyavEd1CWFI+Zrasq319fOu
P3uVOJWdlg1gD6eOv95X5zKYUrQq5m96aWsQHTLuWpE2WDRSzpEFd0GUd1Ky4lcK
sfFTrKDQ5UZdvS9j+aODGdvXam9s12FQSw/PwD+VhydFrtWzFdULi6j6Lq/Ps6L2
mpYO0+kFQGu9Il2oxYTRxHmhtwTF5u309aDwNp1PHb43NP0hxmaKFWnxIRlITfwk
RWGSZtQOWSIZNrXLjlYcs1ujKCXLdOxarPyARz/2ARxcY1fn6Do22aDBfCCj40ov
Lsq9vhObOoGs4+ypXi5hZDLvJw5+e7zqnNELP2bGstRNZAD4PX/q3m1hxN7ktdMd
zxwQzbliIEMAhG/DH01DvtOWhfDrs3Iwey7rnw5P4khsb9y1Pwbwla221oJSjCV3
+9FQQpjsPdP6DnrgDKHxPfcmaTpXzpWTBfrNb9Dyfhas951GwIJNblfugaWgE6j/
e6Hd6Wu/8RIxPBp8GIzKCQ2YuxN4RKGDQs0ncH6vKpI7dPYpp4XZ9JrwAJLr77dH
vEt9NKXf4DnhkUYWx22XqglLu3a5Q5w4bR9z3A3Xcc8sRUlfn35tVwDjy8nXzSu8
zaCv+dSs42s/UpC552TeycgxTSFT6l71UtX+UIZpKsjJh35R6/qVBUNg+00I5kSv
P2EsIUfH3JEcvIcxMxm7089ZR7hEY3pwUL9royNEJSV4ZSBMUUtw058+1INgXPJi
MxCQW8+wgKSgyBbn4ltetlG7tYZuRVlRB99dcvow9TWEfAmxk8CBHz10ZC24K6c8
TmYurTCY8UUcadOQJnMOicz/t+68FFJKsN1KFyg6HnR1NYNwO2o6EbT2WifEs/pr
04ZLl0Bkh89H4Ca9fwFPIS6Y4+AKGBsp0fXmbMIhhI63PlutUxKvjnoj8Cw5Nevx
6GR+VpTqNJYWFVPi1p7pWuRj1VXvJ/36IJTCs17JIoVKjwCuE85B2lXZ2Yufm5DV
a+oE/1GfN1lYhMtJ8/L4/frKpfRPwrtgeNvLFfXNYTpJaCqqNHwsSdrGmyAS72x+
RtbsgJVef4JI7pxfDwUiNVgVBN7XjmU4iE3DCDrj56Mutmk9zHZ0tuSlKoYGrQkJ
PEKepLrlCWAq1NAZAenFVg+YAjnjnePIISP7VWF6OBkQdZAPTbdpPQIh/pPSN4ZW
xqv+811mlFVbp6ZmoZ+sDv5+EHgbdEEUoMwHlPa4KiX+vArxXTJzpseTlqtrdkrk
GphLyJ/TlwxZgwtmQIQXa4pHf/0pMqKJWPUHEeOwcfwu3Ke3KOtYzkdnEBEATFYW
/xiOzcJORtblA30eEA0Wcu9qSokFUtO9YiIFL2ULZXwyJsev48l7XxtSA4Z2Wx4d
huN3p8rbcsiHO1+i671FgoTh/YAXbk2pA11h4W8xsOME/2PwmLYqROCfcB/pnEiN
hmKm3wkW/erslPDuNzbGKmnj0rfkDO5VLnWVCeypNknVVGyDwsnO1OMaHJ0peaIy
/MM5PQ06CNIzij2HqfE2GiHkwFlCor/NX5ZYhHBjrKi0z0Cm0EzZw54TlqRKjgKI
p/1BqU3NG1CCc5/+e1s6mqrUw7TBYYWcV5vW4NGz7x0Wf4/F83bPJ0f7iKyTMy9Y
zebdeE4dITemIjWUyQAfUTz48UAFUJz0bx2YCA8c9EOoxhBspUHApfzkJrD0tMiX
/O+LeoiwYWw9fn+6J7TLShuBPyyhzdbYH7bqADNVrvCzsuybTsjYoXprul3QbFAO
NollHKjKWAK1vxXL13z2IXaXudGFvnwdRQsuN9T1Dx3FPc2sFJGCARYylY/Py3oG
2JmBR5N7qXqSM0zE+/A7NzbR4foaBhEral2UDAfupRTWkydYgtl4MDXJ09BkJm0e
cR+Nn9h+M+0SSq4+SGURLnhbK2lf0ixIXUo7eKuVdEh4ZIFFnvhWOdmjP0R3Neu9
uk6bnP+wXX/NtxBGwu0UGadpcfk6hPnULmiTOutjenSIjgQQDB/DAFtldfsO34i7
gVybT4eO8oHfXi/4kjUFWfGua6727mfrsZ/i6Bf9JlbblMy6DHvSD4u084OgN8wz
IwuzpRnHhAGN0GrNUhbO5aD8B6FL7QzQcQzdMQA21I90U5OYZsRN2ap2+stJdeY2
yMkqIiKHfHzaONs6D/AnH6eCBDOlhwNwtzJP+qbvmjTzEkH3wlEnFDSPcb6iCe7z
WPk0AlkenJxeq/i4zYhqLt/r1ynKy58rcauRzvVbjzOXmEqcNg7BKZ5w28bidi06
NWTc2L0yoh+gaVOj/4AqIec0PoVLaUW0Zaq81XUbqq6pNpjeZLBOgUfihsQ7d5Yu
MSLF3ZcagSRl2TnTuhpZiscirVwE68vjXqcLNHUWxtU6hz636p4S0bbwj+XRfblP
TZE158p0ZM03fmMdPlhizpNre8Xd+yyqxC0j+LnAtVUZvdFYlnG5z3uzDJcgeYh6
eTUngA97EFZc0qgLsEmdvzPklMslJ5Udj4ZUk7BQtyoaHpTuygU3IVcyzPCLh2U1
SgdrJ1OaynlUU0X06Yrd8yTbLtaIYDHBhReQH0OrVEvDqpYNgFcxdcT04uNpfOkt
to4pLkL/twYf0TZuSJIMaG5Bmwlu7nBFyo3B1lw0CsoO8eRqtBph9grI+puAb4AW
0/Hh2DG93/ekFne60yP5/hAFhNiJTWPcTyaXUQLaG3RW9DsrwKDcC8gORbFlj3tl
DqiIOdmaEGrLw3Mq+W3Rue2IHLeTXUboRRLeJeHqPsfMX7zzMLvtQfGQe6zG7Blt
eY1J9ng/q4MdKGo5XvTH+8/OyRgvcTrBe3nYWIS+0vbnDlfnnHBo1UQ0eH+ChsFl
MxeH8JRPmbc3t5FGUGnl25YKt9QbzF5qnYpVRzVFPgduS38gKW+Pb9qEtK/J+Tdt
O+3ITMRaPyqwFmwG2796Jotgd1RGSX9RH16U0Qj5GKhmRvqID0GX5STYNhKhhpR/
x1KhNk0c2M/t6XDsUOEaRj8iol1wELGT9X/qX5t6XysPqBZYTB+O6ruic16+qECL
xW4d6a+1rPrgqe55u6F50F5Tvf+5rhlqemsfoyDnRAsA8kQA+qzhVwVc2LqvPDGS
q1htM2gxWkS+siKPqtQ2ZYp66vsG0k+KYurDvLMv6JcZBfW9mIoXaVx4lDn2pmIx
kJjuw5wBnHzl+TDiYzaMfdKJSG/aFf65MHzmEPoTRvcv4tVrmWJeYwRYfkzXs56i
NcSopR90TyEbM0AHHdm+oEsVrCX3WRk+Vszpuso4aYz/s9K06zpEr45TSNOPxouN
Ix6SQDFzxxnEOTria4DS75xxTofv9CM0p2JTwzNgxcgRLmSQwOOKjMn97v047cUM
gsFGcl9rY1k0Y9diFQlFfco2dniPs4H2sMv7zkQIc/W5qH2hNuC6GqJ2kJ2/82nc
D8PdJJf+rIEFRis1jl+qYA2MSWA0kgB5l5vLSglnesOC6ZXFNkK/5wWVcnU26xk6
g+4Ru8TKT3ahitR7SaNk16cIMwssVI8/74ZODDBo/hMsv6hPa/4uILXnj/PpzVMv
ILF/hHSJTxvBeGaSwCuFRA2XhYRdUjPN4Wq+ts60Ig7GNJOtQbD5rwLHtfqFmmOg
PwZPTMkKrDleg47xeozFBtLMU823HWK7oILKKKXPSxBjO8QeLyNI7BIG+v37B9fU
6/1A03aShht00u+0FCT+F2fG1d0ndlLF403CMpPrYu1fMwhLw67zEZKhppWTMxVA
p3WSSMilzRR6jQMW1iDWyODBRGIM8BGHm0YfJWDBL+u/59f75iguQD2l4rAGbZnt
9Lc9vbCXcDP2sGAJMD+CZShP5S6eDPrVGEOjMzTUIktfp+H4R+0wCsmp6akW5SBR
8ddbFfkmfFQ0m4o3naN+o5EJd0it7E2G9DQcCl1xciKEo9so0aHQ62O4wbULLbSS
CuDC2aPQplFMsY3lX2ndQRCPt0PNK02ucHRJQH8oI71oUsDyin3FSZ5uF2bVvYMC
rfItrQy8oYB15s6CeJ2amVkUbah2GT0K2h6UIWx6fYFvSTLUFvkmyLqiSTlZNdoV
N1GyDZYTIrBH7/CJEaaFFH04NC5rvSuxB9XmnrRJw0eP+ox6O8RmaAomqoaz34SL
hwkruH+DCNkcwxY+EUUo1PTWSGvFY03LMHnLGL1JQA3H3R+uXrz0FEiYfypF3iqZ
HdAqJUxmJp6C/N7zPD6HDlvy9N/nONaVHRXfP3/amf6GYW6gVdeQk1XulWGx0gQE
2vRKIjNggimXnOtpS9gIRAowcMyEkqveyLnzk0jqisF+DL/v1Y7uCGVO3HnIMN36
/YZi+3sBVXkwK9wuoNdHoCyAIvyo4UIdzcYI4ZXYIMFUj19rhC1LO5eScbTGG7mY
EyQAWkUn7/SK64RFsI+o8lKdOwYpFhPvbHiah99wlv+e+dQONn02LOnLI9KR0JPU
zGLDRcya/2rbJD9DmGUgkO/Bo3yGMcME3eu1pGQeeYNbXdK/c9Fb3ztrXqSUkysn
6cjxhNdx9BZtLOB34xOEptA+VwsIyKXGfvqEhF1pbDxpIp9qQlh/5r2O61vZPTLf
O2NJDrFigzWFi5t1IMOTqqaNKE4PWba5wX0SrWBujDhCc3QBOA/miTrhQ128njps
y6UfU2lG5myr2zBM/Fr+/+3BrN2It8z6majiWln0xS0gafhgynzzs0C0b2Vvtr+w
6JXacA5zohiC8gwLKbZ5cXwzDMKdZFFVZiyw23wE109TCb7A228p5AGSZFtsVNX5
RhvO57kGmTQvlvtkJ1kXO45jRnsaZWKePXCN58mMAQ+opS9DRXL+dZl0E4eER6RO
Y1qx2a7FmuFEcXi0fCLhtRXst5ZHH37wCuDE2e0cbYdKzPZYmwMLxSX33XKGaON+
39OgfmgtVhCVe3e+MNXosdOAzwC892kg0JiaPOyLU/5jY0NoEUz8265Z5HaMGjUX
II0PRjl6WRqNARmcktaUMcMhwEaVoW6n6ODw187x4i6AMUBkkUGGQ95AupBat+UK
WRZCHfNbC6Ogr1DkUaW6EGicsw5jTtQw7vbAjRDPlzhBvO1dwjFo11P6yCeD8pRm
Z5MbpomG9fuRauQ2SyJQtALJY0oN7dfr15ZQH3fCYNBR573rhsAipXpB7fBNdzNl
aYpoKfTcUz+BOEgnZVsXxRkij54JX+R4zMqk6ye6LP4B1LpbOnFhb+no2Azz4E4L
2zXlgIY7Q3MayhfsQ0sOvQlM3uyjwaVIgy5cfuvC14aFG44HYdJ7R5l510ra/HKl
zpDdDMx00Ncl+wpYkYbZ8ZEjVdr/cGzDZBFEbjSb1Eguij9WSuUBPRq+AldJr1eK
ANc+54V5UebeSFc62YEzoVN94tr9EaZFJX7SHYUQ3SkROV+Ie0DBUSEeTtkslLzm
uK859xRsvI2LeJHhj+MVHIO8dOrkaw1WfMsGki9YzPUHoafv1p8TRzI7wMP75bAu
/RKKAJEn+/7zcXYIVXS2CNyBXaedLmgIo4nRtEdOG9iKWQsJmsQCjvvZR4/bjiqi
69l9xouDTA01J8k2USIMryJB0QEievFfpqV+KWe9rwvbYtOQ7DdAvCLol14pYoN7
+YR9HgADg9l5jzCGzE04J+JO+HdyVUZcbvvSWE3eBwizbq6LhxGiKkqLKDl/rOha
H7ZgptNM+PRkgIrcgZLaSszmwWG4zSs/kzUrpHlz9cxFZZ1PejBcX70wg5PoFR6B
TareeLiONNyz+Rj9ZsW8fOMzf02/8DlDwsxe6FsBhJe8v/BJdfaLBL+Sq6nLxrj9
HgG7xnciGOQMd6SdRo5p/FOgCZsR8v39sTAgub2K8E0bPxFd0jYmYZC0D/4U8MJA
8tVwz/JbvOO2j8Jt9Uw1Cl/MZENMkVionUjlb9hBpHFTMveuXa5HkR1ouLmd7w+b
5FWPlv1xQu+BHjNiGFaOmh22MVhHYBhJ3cDkBnytxJM5nWi6qU+z+lqwiNNOHZSR
YO1PqHCWLG+uN2bIgzw0Eg3dZlJUE2o4NGzh/9yKpPePtciZ5c8x2u0uPBz4fNn1
ieaySYqwSY/zscwdn9M6LMeR+sq9nQGQGah+hKr0JmeCIzP+8B/y+/tztjxqqMVX
DAVp2HraMw0Sqx0Jm5pgvplqZD5vxwg9PLa2Ijx3+lx/U6u6ODSxtZHBC7gvphkY
iLQwNfOnOiC6FklVn5TIxTIRrrtn8bzg02TJJa0VIHH8wFHnUYrSPZ5biWn6740w
QahjwwJdwwg/zpeyXVtGC0Lr5HI2xF2R8ZB2BgqAWqQHu+MCE3Uh0QAAHe2gl8dt
T1GDL1r1YaAqNsByXTDZmlYwKrgAOV5dEFmoHTM4ue3ym318rWI+9Tlo2VM+tmIj
3hCbeSgRxvL01ZSJpHON4Dl/IEkX8H8Bh0XX+KJb8J2iFuVlM8mzKgzpLAKVFyLi
oC406Y2R8l1XR1o4tDEDVrm4FrzBm5M22CFJXoi5LPQcYz8/RC62YyLZVpHkUs61
hpJXWC6qXELqtw5XRqwGtj3+ge9q5HDzfFObMPd6mjDxCuylqMC4/yYaj7L9N1uy
X9YO2RlOwH1huX62dHuYePP036pxdieFz2Cl0MbuPAKJJl3SjjXStAIUiCPFKjjO
oYs+Y5Ns5oZOe7fB1J9ksYanNaMVF2pZcF7oHJiSN4q37LdRJc1nD/zEkU4M/hPP
nETjH8WacO8VssLpeM+h8DVTKhhNkYotrFt+w9dYfQyfxZ21FSDYmfMlFucoC3bs
glQDy2rfoCPc/e6vWLBz4ZLlAlzzVchLMoTJtZx1axdkFMl3tmMFdtzLjxaV80Eq
ZrrMPw/7l2rQEFulr0Ck2SQF1k++nzuoRUpx/bn665hnUWgx0jOZKFzU37rE12v6
hY8NrD5xuiwE9MLnamVkp72sbRd/FC7Vf6mWd+4j0lybvF1EQr6NPYXuPptPc89m
Oqt20gnaNm50kI+uDlwL34e6f2LIrAVhMswOI+bF8QOufABCmKndrH6sfZhUVQ5C
KCOWelbrUdAEgRh5W8ZbLkLa9Iz/0llRMOosbDIjIu+UGSc+YzghgPl0LGNP8Oy8
CBJuhcCP8eCiFIRb4xFSEJt0Maoh2IWm+JcSfS05fxvcgn8a0U2/XR8CZ/TDBCPV
2rKJnDEWmNJBy7sAcr0NsTn2EJuckdredOxxk2gtf+Z0VuCGn6K/53nm3U9Zo8a3
ZJyc4LCMJdx4I03g/ZY1utn/t+TX9//71Qj5JCtzyakUrsrTiISgMN2GX+YAzkbl
GHss47QVVitKCfTDy1aBsvpIFSrodsXy+GyuZr06Fdt2Kb0z3hIBslRQLDWFFkKF
iquGg+5IB/RqZ4TH4zRmLDgoaZArobXcGaGUQUwEXXUYjFpy6D5FLUhMCKjWJA9G
+b0eze5PSICN/DHxCG9ngFGZ9l/AYu1kW7OUndo0nUcWAxEfqyES+Auo5JSfv/6N
og+fE/XISBE5fXn9cm8OvZEIcE3qdRWUkvPfCNf2cgFyFywszyhAVAOSYABq1EDA
L8Onc8FUH5H3SNY5OIwrISY7VKmFDpIMfsJv/hDE2P0vslOP3qQHvvu6Nuwj+SkI
MY9Mi+6AbcTcS4qq9ckcfsG6MORpzfnsaBJbskB9OET24u90vcGlYDY8Wb85ReWU
1pj0U0xzZCdqbHLsMxHCWowW3csdTz6pKV0YYJ4ZIbBcnBUhWb7cyjR8K2qV9XmJ
Hkd83sabiAVDiJqfjXtDx+Kvwa0ntAWlGWEqETiPfDaUFa4U4utEKXhf2fIBt29e
uqQogxuhS5BIackdkxP0w9HFdiK1Sr1jCQixdRNA2297fukUnVpCVC5Z+LKIX8t7
sgcgfPUhuO+5tGstFm3/SfJLHkLgfD5lBHJHloKw/IRLUCLch6iIp6teSDqogbcU
/87Yl8AJTv6kqHVvvrw/Yc6il3Es4SpiO1ICcIoqhDHOqXZhouzMMpBDBKpljd2k
pkeXGJ+JD1eI33/O8QlnlgAZYD7DhKnZhfpzIkUzdNJp3oIrAnrEiBtjcYtdeLIa
xOgSUD2uQC+cOsO/emlYJLzXxmTYtv5BuQyRlVKww7YiFm0T3vlBn1r+PdBX+Dwo
h6iKADpfxkxPqo8aeQxLy8V6987pybn9LZdIE6c9hXzZgvaELW3m4fBHA674S9lm
7FkbtmCrY0b3yUrrk11CwYUGYS4Q1w330hmHhd6Y9tiOl2N1XdHtgzxr7VG+sAbj
rcbE1/5mPL+Z0yWBsE6AUJzUzYai3Uhh5kmLuA2koRqpgeltb+XoxjRc7xYjDKrx
/VWoIFnMX3xBoPSvqt0AUM1Vts+JcTJcLn7qDb1hg3MXH0ld9YCJQGAAVCD6vEo5
UvsdqvdByw/Rz6kwZK/usQ1nkEKuPLRkG3UrIOWR5JxsYCudjs5Fma2Ypk0gQOYd
fpGIkdj13GdtI+J2nHuxzQIJTbmeRrW2bFiiUTqnXP/gE8JXbXRc9utzC/J7LJ+4
fOhSgYLvavO8HG5eX2tHYijUPIx/6TNHnDiBxyEOv1Us9WL35bFQwD03LpBkca8Y
pUQtT9LX6wOP+ujtgop8QIiCeNR6wcB43N8c18VgZpQITCx3aPROusME9XW5BX8+
BOE/UrSQmug5Ax+nzP5pG1CEK7pRaMmuDYspSKCgQ9l++9v5cBfvlkGJYHx/c+n0
PGycpwgMgkHRTbnawVSWjJNZwfEYJG1nebeg++HVn7JqUOBaWysKcGkZrZwe29YU
AwLCUZf73anlfX2OPo0R0tQa64hGkKpmf0Q4y0ZDm2PV9yFbqe1x+E8vuNZT8i9P
XOKhbzIOk5Q6ceWjr1bfgLLIKSeBXO//CAECKmX4CJLKQhoVnW2AnprHwx5OFTYd
pp71F92ZlW+q68WTppiiCeuZaa6jRyvilFJwT/wld82uwOLCt0jEQHu5pIYU7znl
q1RHeIJw1ZUiCwuTOjZUK1121edCp1B3+104QkFvyp7vGsJ2y3nfiFd2juwCJyCv
ddBDvjOHfOsqsOcqvmmL/WPv2hua2FpqOTkLXPOqZRAVwsxHoNgVdEKOvotzsrKD
hHgqB/PNjluB+XhoeSV92SC1HrzghNy27MVSyBC/aCkL6Bp9pDxomaEWCsXDJWwo
lZ2cuSEsNvD7qfvefDJLlZCh3q7701lcgLGRLWK4yqIvUrvc5YS2Iowdij7BJ3QL
PE5dJtaqDKFbebDcnhplHk9WSftDr/gFpzWicgQzE3TvJjA97sMtSWBIsLUBv2I+
qrSahGzhevrVNIiC8L/GCyKijh0gWKCSX9S9Xte5kQKGOUiv6CpUNMgKw9BQXc8c
ehNnvi+xawK2LmqPp7ljmCu4XJJmo8zVTKs4MlROB/IolPgZEYsRDqjbR6v+3lH9
7Dyx6peH1NflbWQv8Qah6MCYm7PWWXvzclJJXPtRRDchZ6qAiUyIzJbfgcYzJcco
QPCS8RyGKHjqttSj/zlXf+7lRpPPno3PCj7XRf5+P27DvvEDcvBXuvIm6TcI7ujE
h1YjVH/KkAIjc80JuRbY+Wuk3RoCfzIoQOF3zi/WrLd9N9LhT/1L8JbSDFfhaLpC
kA40iSP6BmtA3oJNzh746PLfrlMrgayz/H0RuboO/7RHBAH8HHvaX4yxzFEBd9rg
YmXDnp+pOs+z3kJqdneUkmwgA+n+YhGjAvWoX1RAggT6g0jxtX2NZ6qNQ3I/DU9m
iqZFF589AfJUu/cWiTbJ1icTxK2hfV+zITgsGDLYB133V0D9yVGu7BRhAykXTkEa
z237IABf2vBUxqK2lA7X58puQGFdNF0Tyszd4gV1gWSyAJGFxYSa8TG0lzG/qSIC
jBZvNyJuCLvik5T+aWI7Y2PgTdDTkotTUbRou8NUmmhXgWSVN8Dysggrt9kllkBt
1yP0cylll8+vXqdcRDwyq6Xo3uy93h4jmTxZXEnfNSDjLNZCudTUYLb/lkpauzrH
vue9cHhwxvS0fuQp7+C46vk51qblz/PuQ31q+HyYNMFQSau+eJ1/+pUMfxHwEbhV
PgNCzfOa1zmvquDYpyrgMb6k8BEG6asJKOImfghcyDU/agtBsiKzTUHw1KwK4Kyh
0b48zT70PAkY3UXu98/CdiaN8TTwsd+6ZVOsVSq08xvoPi3nKidaiqd4FwWALXDL
KCXihmvTQxJtKHWqmAbU6UsFhQFnoHvFJcSobnEmRRRD+rsfpiNacAQBp1Y7Q+/z
gR+3nnsusjingyDYQpzJ1Ap9f69dpxlMxS9xTpmfxxtzRNhptR+pG88QhiDQB7jc
acyh01VZNuxa326o/5fgZr24w7AUlytB248E6mYN6YgdumJ/XImsMZc1Ql6qS84m
FJFLDYtVM0kaNs24/I3gAaz673uleFIoOLro/MbqhhqOm7p3/WYuRByYZmY88ylx
4ClVNEN+Y2SaBIGqzHnkVP4qMVcqtvIY5i+Lc0vHNjl1D/891dSo1nDmuuUQlL2G
edRE4P8G/q7iSbgT2EYyg8Y+sBMQbaQYLUFt0I02w8E/vnUhsxUJwrriHYMbtF2U
FMBvF7xzlZkV7zPHZdWCrXFKBr0I9cJC8Ne3nCXPzsuT6CzmKf55R9vM5HSwI/mr
ALX0HTJZWRnwSWB7hCxf9zRRb2BeYOXuFs5LS7BLFbC8qBMCoXaFviZtIXJkwbl1
9VxXnSNC8pfAb9AlFnSaWoJRWmjZavPHVkE4JXuUYXuxX5oZY34fBQthpuzQtn7O
rPewqG451dbJ8TmZKy191VDbZLINuSI9jpA4UbuG6AjIXg4I6fRL9adTc1ZegxIY
ogh0YYiBGrcvZTS1/CbG7v03BtIj6I4R1CrZ2mSHrXs44WgFe0jfd16CgrUJOG1L
ainJbM+iduyDwEmyjtBpec2oZmWCdKs7NLznBnIXMIzgHJpR9eBzeo4t49t7C6py
bs38sjRnZpSIdzlSHiuMqUN+0GmqoLr4LupwTWPXduyVG713DhTx6KMGv93cuQtr
cFMjI/bOtVIogzDdDXj7wCDWg94B4WHv6KGk696+lFGTZH6n1eUCtQ8k3bImAKAk
DkBrdSvGfBkLF6tvvrNb0qDHIl1QdLM50VDrZRQQTNiUzv1p3Wi/FqamAUQFrHBT
mtr6MW7Jq3TcA70YurvJUHJMYJcbxOE+UKso6Q3LBQ0JRuKdNo8despKnGf8AVFu
qgj2q3DQw+Rc1Qb9PmYeyOh/lrwh1weqwtMZqVAUtsNVtWBJGHq0a/m3Vchgr2Bo
UGE7ULcMJ5vP433YZXQUgueAGx1XoMJ+nKRn2OVD+WbfsSj3B20C0+vVnHklFr+e
VGMDyoCYegsgRKvGlXar0c7wys4h/jPYTc4z432hRdprdIJ0MwcdBvHqmn4LK6hj
EmhjEqkf+4eTCto0WBDvytUZMYiYxmJ5lvKmjxLio1J2VAcHZW1TZx6a6RBjJ9EV
gg98TnQORntyHhlm8RB1dOvT5uE4bmYi+MkS5LuVJrLEUcYx7/GMeCrcf5X4DK8i
i5MkJCeBlfZFlOFXD5JcoA2tP7XA75xIiT0wily+zsdX/S/7bWf2eYi/6FJZCol6
Nzoy44BuwNeQGGcawVbehjJ9W53pQjAweMvFGF7pj7iuGCq3uV66j5E06WFAfcfk
sMovSnvwEWaa3ql9bfgtb3VTQuYqAvDVEjszNJa4WuFOkRqoF48DDQu12ux7DiJu
aFnE722U+qnIDud82AS1pG9EN9q8UHPQC1QoSP1cOnDVTkIuijjZwd728hFJgv4x
BSGJ0inyQo7sCmJxb4ApC6lrEPvzxL3fDqfRWvhHNKI21L6VOGQV21gdZFtTYOgq
c4XIznGs87Ge8ztjteezXOC/c6xVwLbtQ9yaM7FzksUmGdiAOeEalu1rsP8ojyAy
wvvCfSOGupyIIaADQvBq5jSmtcPoaMUGWelT+IoFbGWwVhNX63bjabFj3p4rVFGo
w2BRl6R4p56iiH5L8bOa2pBfTAtKvupHpla2eqw2UMBBfCN6Sn+LqMbNenYrTSFh
SjspiMIjuAQVUR4Y/pE8lJkK1zG7hDz/Bpr3rPl3rvsFICD22WOI5r7xIxID4PWU
9uTxzJfsZBIyS4OoNTw/I9A5Ihe7nI3IOvZauhnJB/PSb3hYY70M0CA6fB97AyOo
pByPrpBER0diDHHAT3h6pySk9lrci8euYx9VuuZC3o6xX1cVEC8weISRYd68+T+Y
UVN71nMeIizWLEvWO1D8AJY2ZAcAIA/pI0wXYWFsgRpattUT1Kcnjk3iuq4n5/Lp
z4jl+aEYB6GD7VjV55Wb3AaiD2b8LUENrV82JGxfVqUO6jCqkHUrAyyjlINWjKVM
jLBwBuKhvNFIqNnAutcU50IEzt+Sa3drgwTx59uGK6k5xL4DdSvlI+EmvQqBwlVj
PNGeuWsEw7hLGWfZtBqlsanLci1agUGFNNAfJ6Iz5DMR/qLB8InToG/eLcBJ5vOj
ajqlrpjeDV5nStU92fHKu5+SNZc1jlxuD4G3CTiuFG8Tjh2N4llr+zDecWv5yZY3
q47BaAbWR9XzttROH/+8W/BPRDcfbbBMNmMqFYKfeJ8qhOH/tRW53RqpeWZaQ+Ni
+WMmkTDOjRR/B2SAfKQldAtsD7/roRVLghcAvr2mQcZ8eae5lEwnM1hyXhayUnvf
601bXclf5YefZlqfv8CReAOwg+/bjJdR87j3KxAeQjDGaSBmbvFvKT9OQ35tYGgD
r4kc06K8a0no6S5wWJJ6JZPYbFYtFuR4XUfrcdBXrBUuCxZSdLN2Do++EkjnLkQW
QTzMjUO53mUzk1W894v8Z0Esr9kwl1XJjy1md3sYJzDBCwjHNcuv4d9gn8vboAbg
J6EBs/C4PtBRNaCr9bPXCo0rCNj/vaaZJ1BTaGSv/3Vvv16wFPo3Qc33DP8yEewf
yw/GRrkE9EDpYbYeJDqzrRFz3nqyhnjgv3hBGVqj3Z/saJB0dCH4j1+vEc//KTst
xIEr6n7od9s7jCnQQHyBSkLja17NoXvXNZlWcxPZtZ8NkdWK9UMsxcMjVM//HwU7
RgDBOrl/KoRvdz/VikVbcN0+xSWUX5ErRDUl1hm9IC/ZBcUFF0xy72YJ25bTKzYq
QDFcxtGK6R+yV/OkQ7JujMJYG2kVAjB7tpv/Jn2rCQ/R7TaqY2/MjIDeCVknQXlp
BOv34e4EeUBRjMDgF9aG3KOlcFQlKcZQH+Tv2pyLltGaQl4s2ApdEbysHcGxQAYa
HK5R8PAl/BWjyZpWn94G2NhspStg1s+juV6RMxgeCZPqmNs2FtYTeTpJF8EkbT0f
5nBYLCLkuexrdz6uVjgCLx4sMpvbcZkXj5u9KDWt/onGM/l7bsjQI1ut64Ov7Brl
R0dZbvzhRYV+felVYmAzz7xF/qwinJtjaAsS2ah8PNT3olnSUTpW8IIqL97Be9e4
yELFB3drA928sXWDCLC4SyQEZHLsQ9kTJcLwnBZR0H2iq14MqWiX6DPOmwg2o4hr
b6E+z1Tsk+sef3lzW+Pt4U0GHf/5cOpwmjQj+BsQ9PGZMHm3CzqbXR0WuU+drCBD
lfUovsa+1RlpnCEIE514llsC4LT8k1iBCChU1vy+rlvQQujnLFkJH4gbTlG2u6Qe
8U5VGgWHwLn123MT74Jpjb6vBdFod3GM1JvYjsgbJifhgYt+7A0Ydoo61+r/b2v2
yLCBeWi0haETxN9ckj1I6Mn44CF17BPW6YzGeL0FAa5YyJ/f+j+4XePv4yWYCoaj
8Fm57OpmVIUWd6XFZbGLocEVvmuxH7i+CZ0JVmE4QQfA7/l9j5pWmJF9EnYmpwgA
8YlcrmNxa/EHc0Rx9qUYgtN6jR0ztNVTgxZht7RL3Mi0nLlIxTugyrCGtR6umVji
z8WG28A1kemnVabpK/NIZfZtW9gvxCh5xpKe6m5GutjSUeT3anDLepTvullmpVwH
FsoXEk3TY9RVgU7aQ+l/uLVFq/BsKiGbeoi5gK94cc0uzvC6XNdy/7NVTmFPUcvk
/3odWp1SxUnBPt0opOgCMBnWiWDN4eoVNfH0nPNJrp5kW4l2ZjFqhmCTE3MEdIUg
uPXAp1OVIupXYwhRK7Sv4/APe+uPLEzSIZ5V+eWKKl2jPaM0jgNHZmdL0OmyLZKi
KupQkVp3ZQzdhdZmAllJFKngprMXTqn3evb4LcfkthBx43itynNcGVaskHunb6h9
a88PbREeB2rjWsEzAK/FiYl5UfDankNZBdJaCUVy67s5kAIbkT7TQkob2UPGh5iF
ey66NQj50/n8OxqZJ1FNE96MHtaIjOUmckev2Rk+XUAbZHRJfW2liYiUYnZHdhRt
oVL3Cldnn1ejBO7f6F/yqHOwptbINlhIgzfCcAG2cKGHeNaF5RJjbxxsIjceqIpG
cWcPvqkijoqFxmvMlOEqZqo2Q6YR0dh0BJpOEFDvT/69TAw8s7gO3YC6nKI5Rdn6
vjFUSxXVMywjB9T8I7Qr7ap+2n0TUyAh1+1chDJ/pNQSFFH9i2QhGvKxu2AyKLpF
0qJ0PaG74aeH4NCfktVnTGwV0nfVwAwzTKbv5mtiSLHklbVGZCx49ExNbe3jWKIC
rSr+04cOyE7i1HcPlOIs7f8DMViZKR5jGSWvVuzvWXZODf6XUHBFaHd1Vf8ziM+D
XIspjfcjl/DgvBc6c7nkejG8cuqAFRse53jub5kUtYyunCGvqnNi7IokKuWu0VFC
R7sdjSd4pA0JspTFyQfVtdJhQFxYVFxZ7WvvSr428qMuOINE/gXbcRJIssQzTqlo
uAb2ZtHWk+1PbmvYl5W42G/CL6CqRsUEkxbDOdd4TAVgzxuyBUceQmBZTjv55q24
lcfJ8Rqs8O3g8e3nMtxfzSLaDYDjKAaflHriyTW1TNU9HW3vbimTfeBv0rW4Gih+
fXOVHK+aIup/NM+PmI5Vp22r+WlustJmsub1Iy6EhHGkeOcDxsJYje3W9yw2+qUc
MVcF0Ka/D5uyrLFYCzAkFrQVqCfFon3aCAjPKpDpFJQnXpAyvhzCBoSAPk4lj/SK
stcqckKL7rqVit9fBkS7S5HzTG1rhJCsu2VYtGIuTL1N3fpcyFTbW6AANs7vC83B
foWTUXco7+i9n2TmYQF24pUy86Wv47lNGdzsuHf1uFktjMlPr+TpRwAphZ52c+UN
fOLqV+YyikfbeiIAJPRBKokTuuhRHLm988Zu0BF8uGtTEAxH7f8m7gJuqrdbsX1u
rzrKhbRIBT5LZ/bnBNmOPmlVX1wOJFXcoic2LaC4PQI2vmpzQWPwbDYnX5ptyTZk
ws35i8T795e3gjPvPqjnaDrQuXGI+AsY4pnE8snkMo5W91Lrkfp2vKZaRhrlXLBn
cpVRfsAV1WCzYzDuRyyVhFIniEo88KPIp/svE0gdaTpaXcKHLYcnGSHWSJYAOgVV
Mk4hzEmP6ivm1bfy7QpNWR/hFe/BY/feU9nXjMDx7++bg/EhiRYOr0QFzZKbPcCc
t2owrIbkUVgnPfma2LLc/8REJxB18Z5uVCznMc04/dabNPWV5+Hv9eaHFfU04jBo
lWA4gW2DKyW6Ww/Lk7IGp8VvZdIEBhGQcPMOqXIipuygv1g3QmnC/enQUo33Cet8
R+34Pu3o85GsBBTDCNJah7NZvyqv0B03TXi3hxgzudTX4OLJQbjkGTSL8lZh/4rU
k+yli2gR4LevZHDOrZbd1E0re7FGso5swj6FUY00cSWY1iHBDmm4CQoxpcaKhnJ1
SuC3MJsEw6XGyMQTBq/y7M7vkIBGU8BTMOIxMJAyUkWucS9D6AlgHxXHDjiti9J2
ee/4GApvcZmLDH2t4H2uaRBxiz0hAR0hhiEoDE17eWXxoz6lp4Bo6MGRunBPb5/x
fk7gLUVlor8c6kjKdOoabaOx7vpWNAPf1ZamzP0zPH6SdqnjJ/9KE9Q1q7x4j02v
ElLbc4xlddj7f1h5qydxa+BQKYz83ER4olSb3MApE8RwbN6Ln48ZkUiVMc7peA/F
nlRcltUNTtNmXyQL0auvuy+4qXXkbu+GU1OarDGz5CZMZkEV/05CsnV3PWlW3imd
HnwzVszvJyMuMfMb/+hoMVSgbIzZ+kD5hP2PiStOA5xPr2BG6aWW8exPfUuNRjbS
l1MICaZzJzJF1cNKHcutPtKFUa0UGyGhweI/s/VZq5ee3/CSaG/7FrM4IKqDNc5r
7yO/HdduK0PUxrLAAV4diQOsYMH8ghcHCl4gtpnodbp51boi7K15SFFCP7Zd4mmv
0J/I3lohyU3kdLjSyuFRJmOY+uMxaOTts6Kq8LFnjijWqO+9FDJ2BiyTm7pSn0hf
ap5ShSvFVB6jXeiphlAcqPTjJh3KLkW/f2rKPtH7EQafTONtQTEJeTq6zc0xBm4T
+dM2Jtq3MBIioMtMQq2FZGPkky47bMmOd/f4ffDV/nGExX6MBaA0NRMtBG3HyDL/
qt8/y0ohMcv+jw12tAmc+wAcAz8O6Bg94zsihpP9eNXRa74wUba1BULxnC/JIwcT
FY4pbKorRLW7rgw5Gv+VbXf9ErEIllaTvEmpsC4kBibnPY2fe+Rh4yKyYGdSAaCQ
gHhV6rdivjSwdLUogRXOqEqsqXwxh4QHRQBezH137jnYTh1clRDhNenyVfxYcbMy
ZBkTDFMwzmjFPE9NZvJH+VGvkeTn6Pj/NxsVeJ6KUphDy7o4ESdqvc8mSmO6J+Z3
MTeCouvOMEHlsRcmf5abLWWYq0SqQeAnBCmaIXWXI5TcXIw8pDeQq9QHJGFY3vG3
kHPMccUwzFEQBOCoqHW6KjDh4GFOXmnhv1xzjw/VQKCrliv/x6cu6o4xAM4kZGWX
HNSnW3RyIGhNbzrr7AsGZHGgSf2X1tTpQMc63yj5q0aE0lKKVyob/1D3ucR3VqbU
T5bRrwuvoZ3KerTYhaRZA4DmgJ33hgRG7zuVH53S0RyiQ/rXj1m4GTu0Uvl/BSIH
bI83IzmqBosQ5xu6S1H4CcdpAiKpNB+3Ct+z5sr9sGvVnKmxEL2/CK7VAgK8gNWR
VgflgNqQD0Ojmf/31PCF+uTumzy5XdJXiq0N7udr7dE+FRZqwm76DVHqFc657jgc
KnTBlz2uMkd3EmLfxzCVKkIaHbVThpxAI1g8kO32eboqhOTvPPDibp8rrJ4Od9+7
0iUJO/D167e6xEB55cEpYhiPreO/c5i2uyv9OOJPF6pbOwdvbYbqrOsmJHVGnkZn
EfCMkU9l9ORKcE6j7+DNTQVTcMAwwMphOBLLjUBwn1GoJNRb9Lru/QV2vGqMPzfV
iW7a/LOfiBlzkPfWnG4o3cf6/oOom/YwAc+70HVkirn+WftYa4q7cqWwVxSKf/3n
ZbGxdBFiEplyEukk6Ue9F7GwS7N0Wy0qcCsAk7ioThEMfZ9J0lBX+15h4aOfcBoO
Oa+eKljKAFv7K0fYO8hOsidnekutnjHCcnv/fbS/atDmb5kBqsVg/4j1zPcsc+h7
625bYvAPpXhgzU158Xj4AuO5P7wUGjOOwX4yD0ej2Ov65WLJ9oqIbCIpJQ31/P6T
AFKOSa093pHG0uft9NYYwtsR63RHlonpeNKxqcutr2wJTavog24iYZcFQHy7/NbO
H7M08E4dTgE+3Uf6qQkzXQ7shxFpmZZKQccb4DqyKWLfdIgz3wpxUYQus/QwFQTm
SUVZcyqaK2fJSe8shmcjsQDsTRGmeS7T4j+LI5LLJNMOsdjRj61KhAud9L3IoPxK
06VSZnUeHcdXcptxCqcTdn3xN5z+JNL17AnS+DPMorU6GekFXGpDdvLxq1Bf5Z/c
EuL9tegvK0zVoQmsHxwI74A/3fbwnTBR0ZsRHESwS5uUdh8Hyy8dxivOOKj7f8pZ
7SYD7hLkGAt1RCqk9YN4EztM32uIgp5pU8yskhqseYjk4EBBdSRayU5SGPoHbrbQ
yuJ5W3qzW/9tzEoCSR2ffVRBjRG8jFBmGHE6/AqSsuQwL/0QgNDeyA2GFcxBPzpz
3QVZ9UFE3v51oW89gNY9VpPTF4TAAP9pVbbr+7DmeUrgZ1G4fpb3QhJLSTnfwxuf
/9CS0lle/xNDsBwcZUctVZtYEYRpLsG/SSpS9Mh6DnfcjBV3oj+0VAFcJq0HumyC
WzoffQYMzH4+9YmQSYU4wszNg+qn2e9lUSX4BSMmBkNOA2OPZmLPKu4fksrHIcQ7
Q/IkbLZv8JCQ7afypCWiHNIJJS4PpE6CUn+z81dy89Ca6s05wHTDXyJB9PrIOD3W
BUaksEMpYcggfLIHooQ4ZywjBqq5h2pSruhzC6tyz1nClJDZyl/0iamGTMOdnHe0
G+DrgQI98BWI6CkWCr3nddS+LhS9L4hMNL/NE5glyw/ziltSwKZPGiTrK4LvYt+C
yEw8w9s3OTvnoZJlnx6xohzDmSaqJ0xfNq0NO4gzie6OAmyORnotBSbW7lxSPUGE
aA/YCTOekDn+H7EnD+xmfxXo9yUywZiZ/izey9W/wT7Msrp18/R/KCXnRaIo+Z+k
g8fU9j6Xq4oU4EyaKwfBzRO5yTObsreK9cOcV6r3E9Jp5L8COFZMz/vT+v6mAUXE
bgNQxj32Jfp2FKjFC7gjsJAK9Lw1NbMJbjAuiRXI6eJiCcWZvYJkCylMqc8f5uau
sPVHt4EuxfH6JOZX81SCCYwnUfarLgCA0m7brJpd1Ls836QOS1szy0qpzUoGyEnb
uqf6juORLE9gwFbFMNTBAQqdh0ZufV74TXNT+Wl8dnvEzPzLQhb9eXosQ05Dr5JW
dR1RYWe7wztQzxwvxAKPR6uggpJfT07S8L1JbQoQG68q9PkeWY39VUUiXygcnBi8
48jrGs+YZmOzJeLlOIs4ZiUW9/OeBntKcsw/i8D9kWKEj0lUrktYB/bBqpTauTk6
xnOcsL3XQC7k9XMijh1PmY1v98JBUcQUdSz0qApyPQhf+s3cdVuIExyF7FN7jHsO
Qt4BD2bd6bmTOGsVRL1JMAtnGMq478IUuMvBbh3ANW16/xD0z1u9LzYTRuqqa1Yi
G7e+9gJFUzjHo3FcvanYg2a/CDoMhg+z8YAyJCs3hVbqCIRG/QJlVFf90J2z5/lw
9K6F4jnSeJ19q99JS9V8HyaATTv0RJ3+Bgz6bCZE/CvWtPE1zymihuNch+dRifay
qEjuUiDihB6nZLfeQz7LJpcEa1SUcWQkZd7FG0xQby7VdUKuelnGhKQIGL0DmrkO
X27wS0bUISMDrR9OzNPobSybm5UZlRpcRkLr+W61UwrIMmQadRe05n6sDaabWQ7N
MCEub9Y34JO3Iyn+1TqNvTotch2rwYeA5TXB0RyCHN0nlsX07ZqzRuHSWMA+Bhtt
rcB+1HQyCBS51+qc1/t5S00GUaI1Ps/5iXTlROLkr50Bsm4fjs9y2hv++CW4AZcK
z63iWdBAuhAsx45o/ENpx1Cngq0IQAp6rWG8gDQY3vB1ACd8vRZh280JUeAxIET5
NvjbRl8Cm99VZczh+QhmNIqTDZ1aBHW3PhD3Z/Q6fBN8FQzhKSjhAURwZB0o/qN2
c3NXigbQfsSu77rp03dxWvMRgkm5YZIUJD+TU1zW1KNO86TgeTGKSWMycf2CZvHT
S4Y0K3RU/I2lTUlkyQdI7It95UKBkPDWB6CKoyNoZz6gcfYxR5my+0oiLI3xuCD1
hz9YJ1MbgaMKgpalWzfRWAwmL10hXe/E1DcIeGkW/gJW/+BPzDE3wxHDw1DYMgyt
DDSoHtPtHjixS0G32d2+dOtKJ/2UzQgbKkETpRSLHcPDejQRikwY61Ea/RQmAaVA
U/sYCkz0Lw0vDve7O9k9DkjqN9LmbNCSemBPSqcEYLBDv2KNMxvewxkPijDuPNUf
GKnRPbkVfyFFvFrORJiFRJUYzOl8TnVbKUbinVeokf8xS/C3AekUxnNArxkYw2nf
zCa+MS8WdyBXzCFYy7e0j6FgJK64Q6kVfaCsQqATfrMXHWZMglYgUBDYTGIZIEmM
0sVMhJzRNOeDzckOUkWeFQwMTswacQAYukund7+E8FGJYG6usLwsWXA0qiTnfu9g
TKAxW8UtRx/83MNM7seDMg0Pb5LXGYnF2D8pCdcPsVfsMkRnUTr2y3PAPwtjASiC
ulQ5hnHzCV+RkBrJidiZzf0hgSEKWl9XpujHSxkSCCSSI8nd5FF+uRxNJg/qZbpM
6jYlr1lcqC4Hzx1OujJVGVcLzmhz9c5QfibvjoHV5yEfX3WXdbZArMBp8oPV0Ynx
wg3n50WfflA1gQPG7ajRzV8+fyBGvN+Kb2qOR5OlX0+n/buHp8xsMlXK7Mahd57p
4z0BeKAjp6dHm3OW9E9Bprwq6dtGq9W1QvLepkTuq3UfFYRF9xYdO6hnuDNwj8yk
wQuQVpR9zIaGb/rsbqPLFR5zK5xb6pZd72gROFbK459Sr1QVxNFGYVwrM7SyTVvO
G8uaXywW/IUXC2r2RWj+Ku+2d9pL94XC5cRPoCHJkjXfxy6Gx2H+CO0veaUehFWC
uDTAAyEJecvAkCc/7KxyWK6noS+s7fWErCRTTs32tjzqygfS13qOAP14TQDCjQWr
8GdqH2G5XGeS7fWcgpXiPYTPUkQHRBTO7r08Ffu4rnAIYO0+bylQIsSOUN2LkF2j
4KpGYQ2R9nefP1csoDGH3ThUNgGEPdClPp6vh1S/q40xNq3d44BoJPXpFwszS9Lm
skCfpgMjJw7jePCX7EkM6dpW6jX8tQXX1Q4tI3zcpKJGXTStvlIhykagAFiAWXBJ
tiXfY+42EtVcAa5DBX0Q/+52ihtC2FBy4u2IEXnWsiZb/fRquYwIAD2j+SYHCCrs
OLd+wsSRWBpdCnEMkQd/2aq5tA86lL3FtsFrtwk5NoqSpdNdOgko4j549KwyPFfV
wuEifrTLOn9NRGOq8Q+U671KnqOxy0f13QQF8r+fbuIj9DiSTl/gnr/aVaeKjWtk
8p8gj7XCKpwxeZX+2GAJn9xY0n/fQcSX+pkfXh9aRoe7618RTj0/xpDwYrOlYCL7
A+VXZXJfT1oN2QeZCgZeX1CTuLuxO51aazkBJuUVtCC1NOHPX7X6mmxBsMV/01ir
7+Bzzq8X/w70YAJJDAUuS2Of/jYQwQZKazazMox7GyoTBHNEg13K0SU54sdk5BIS
pbc5bFrKEWT+Zk3UxHuB4FtEqY7Sk/C2ym/UBBhJmaPaN3ZR05L+R9d/sl6NpiEa
fjYB/IYPKGQlJykZnRJYb1amq6jdc7kpDPWcq0d2d5V2UbaSWgp86+XahJ4ppUjk
N3clySVqOdxN9HCL8BY4HMma3+JfamZtuG7Ycc+e5Df4HvRwSjWpsWWXxcLmjbU6
4JzSV2Xsf3X0qOq5meAPWlK9bb6iCy+7A+6GIENx1z7C/NW4hEz6WCtuzDHAHgZA
tSoog/5TUhhGI3//P79sYIst9xT8KymmR0Xg//GGdoQegXCrMitFz1nhvfTYJ6KD
lyYpHO1tSyAkM76zMYZDBzJ8scMfQbZQvi5ppiaar6+4ZgNxyKI29E7GE8bix3e3
l1E4i2iTmK3m2GqKnxaGRf88s+4TMQzys6q44g2YO839dkZ9PqrvwqsiYKK2YUHL
3ueqA8bsPv9MTcpXGIcYQzEKhAJJ0PSSq+C3JHcejBiuT7HUSIT3Xyl57VpiSowQ
izzVgfQrytUjfaqs0dk1/K8QCRRhfpzIxl//czFJ9TMxYhVER+2sphwg5Kbh+zt+
LKrH1g1HXiZe9BQysXT9rVQi9bsoASLLmIWzGh98v0foo2lHNJLw74Ji4W/OsmwF
XGSQSXi59E7HaGwNiJ80qLG1WQV2+Ju+p1evQbILSqTXcw6Z5pxLgmDAk5EtTUgZ
vR9XMhBhHNbq0oL1ObOr2KTZ8CFTG23K/2WPa1okSIJrtAcoenDL8VTQhHf1vgHw
goH6ikxBCJvq+EmWVcImeLZDMk6KSz+GBzX48IrE17RC+Kg/XxltOwisJQF7AVKY
BNEXB/RLSNqk/2Jo5Oxk0D15bIpmathO1B4qIirO1EOHCej3zqkDHhHnewCEY/7c
spFYc4EdudoO60Rg0GFWP48hrlOiebNJKHXDhJNiuRdI4K1Bkl/2GgfP8NouhAV1
94/jWPytvC/NnG/z4qrqGy/iDPK+lZ6tvEHQIpsYVzSlIHOsskX0w+OENh7OM95W
pLHtqwWjo4BWJ7HYDpSBKD/eJ63H5Y0gBTmpW8JlMqFA7Ktz5e0btkGA2kkYJxFT
rp1N0k/yEGn5S4ivwMZdf+hWeUw/IwuTBDitOM0o4GRK5UMrl//bQD3k1rCxdvJK
8dBI36D9HhVH3+7PsWbZAKP21ty1PnmkRqorRP2pIcc9LHOeeRPLNnJKbAKm1BxO
rzbiKPOV+EWNQtzpVQLtxer+iXkiKWvLXBVPzLL9qgQxON73XTiLEkAq5gKEKgPT
JiRh91U+lm6pF7XGLQAdBvng1SEFloMximTsYkvxqQvEw2iQHiC7IzcYnUwgLE58
hv8DFIuoBq1Gx6wasQUXGCDlQBKj7U79YlCLESjv4kuRN8s6sYPVySD3R54u/hX2
RNW0Qlh+GQRx5JQTGxg1gzFTBUuQNR19wx2iwoazMK7zXuRarAMlAn6koaMu3mJb
CH12Z3uT/qrR4BIFayGNXJGbYHg5Mx2KjknTfD2dewrQ3ReZx2tVBiFjYNL+iU8V
WqeTLm6soswZPY1CFlXxfUgoOw8qJlVFYVPtKbW9g7sltML+t2DRSW46F2fiIqaL
Gst0UW+MVgqXNSvuUrNHD9shy58LMR0sD3DI/zczfzz8rfa69I4h5T0vzn7Qxd01
SN1e30RykjgG2MiRUjhyPdpmelLbx+5fgWRPmD55+9HXQteudcgV4mjLvWlYVgA5
9qOusCFIy4QBBqGNh41itXohL4mP73k4FgFkZkIx2eISKVfCMHsqkw8V69t+3Ml3
Zx0yB+CH423odHu6zdCJ5Gm4wW7UUtobKSH8P1neu+X7kK2jX0lfgqa4khFzRwfS
z8DAm/PmPtIYK5Jc9WYzkFNJGZe1m/hZ2s8tG87EZZBDc27MkdntXTJym8zhQjkU
yfZMJwDIFSdZqpy8UER42ZQflYvJ3v6wLv4BC4JsWxdpqH+uz06svZ2vQavnpH0j
nmqD5G6TTRppvU0Xgp8oqXSvLIUJr5h92mk5mz1JqPezguOhboOnTYTmzmH97BKx
VdJz/CjRaGHIMEaeVbC/1au+czdrI31lhOdpoeFN/VKjVrR3jgiUOh2Ovao8RRz6
PFB1bCAEDhJNE5nma3uTlRQu1dPFp6bj9J8t0BWG8Aj0j0Xzq+Xf4BXdJK1Wc1k5
fyZL53gMB9vbNcjgu5iF8b0nXd6dWsipJZphF37vT9Jwnkd8QWoVKsOVezoY8ay5
bEPRAn+wQhCug/1sTS2vAIoDC9GBUmfVKrUMqjO5Yivc0RWfPdhNY+SCJRZt2y7N
A11e2Z9ptP/u//4XVHeEhRZaniHGjrxBDFXWdPa00qTid0jIAELyr4wbJhhOK4hM
IZ/B/qRQVwrwC0iXpoiSuMyM9I56ViJKqKhux2FkI8xEQAjVuYeiEI6Lquq3k/pv
/iUIKj15cJh2F5q6AcU3ipiIcegiut4IzJRKhXcsx85La+ypNZVte+kcIVpNjshE
4FV/r4Aay48PAmUw/JNUSGuJmVC9MVS7ZZhyVfgkV/KRX19963o2MXZ6OFVGLvbP
IF4Ca0Vth39hCSTdk3Qs75S1J/RZ7JnwxnRThNUAeZ/IVkzBYx6NJD11qeFgdfA5
lnsJ35j+M06GMCOgif85j7hfrd7Mo8wjq1a1RZfOKy3of00OZDj9BRHww5UUT2CD
E3MRzlZ+mKo3g/+eO1hOL1+UUpr12D32Zs5ZAWoCpcELg0rTspysR1y3ooHoll9V
HPIKjlttCCxZuMPXCbFka8FzCJMdKnLXgQzZYtOpjVP7o1RM4TnO712bqU2mfW9K
qygFMQQMgQvJ9NUXXCQ5nKN4yoZQq/8j9u6pxwWHE5qTiyjWU80I3Kb52DJ9s0Bg
6yYOIdDuG2G0AGnF2Sscme0PZYZfFYXSiWW8dewJItKIFMxzLFdx87DXE9bNfLYe
9hP7ldy8EcEdCqgvAZdk0DNrIR8lFlYl0JcJfDzZJB0l0k8UP7idnZDoUe5ghh7Q
NsqL0CrE5fl9q3LOl7pqp4jlVdTqdwspJK8CIVAG8DFXJLrjV4bphJI2DAsVyjjg
vTnzieDu22/itKPIMoL8+Fg6WT0rnhpLDDNUrLQgQ0MdkBtVfqRphoAzXBfofZci
98YKd7LBXDbyo4IpIWnjy2GZ7RwdPDiueoXal1SmYT/vSxU3lOO28jrGinmgQLgR
AISiy85W92+jFSeEt4ZMY0bPidk2eI8/UMrPPU2jAl88MXq6rwPi3YaQ+miyV71I
6L4GB3GVuasl031aWyE6Qc40o9XgCrUvMnX5qfSRq81cKCW//A83OltBh5ds0BxN
+ngwzEUVaYuJDL9f1ELcTJkeQMIXV4dj1BW124ei/egYuZ9lLuuKe/BD9boVj0zh
TR+becPFxBRmIrSRdYeKg6XHVccB793gWXVxHfKcX4mlfyJBUjLOfOQMCVVQcuRc
st67HU7cMAyMiXwqAyJNsTJ/o2c7eiHD1JA52Kz16v49AzWxK28/mlD6VbqEsYaW
+/zsiHe0HC0pILMpy4Au+7F7lWS7yoqSv+HlaGe6L+JvBllp7wtgHqRDEcGDWVAt
XmqKuTdyoqzXpmw15bwE4zHqwR2I6LORqJsvXzLstMZjXD0Pbfg9lctezMxoubtq
t0vBNXhtK/+mYOq8+zBXoe2lTQbXVDaBft9/vRK88GT5RDeO3/FFBatczf9Tt8ep
x2Ush6oOO24Vp8GHOTJoV63/o8DcTWePbz7RYwaT3iIQ7OsoqWVaJ453UBIcIJTQ
Kvh4n7GpuXzZ6w3GsxEtxK0frBES+LLCt/pOoJ3hr5V0RVXhrvG1X5Ik577XlC5j
nt2aOSgS7eiuJmuZ099FXoE3o6w6cdn+z4Jul2HZbK7yvCFhivADzsFREovjEagE
HVie6k7g9c5N1LMcfF7mmBhvVxKcK53YalnTtZpZRVQCF+NmuTdQRX2QH3J/sjIh
GXukqQUEVDGFsyVUfq3OxDlwuifDAoMfsmaZ6HYuTkyyVvx2N2fY3Lk8RB/7+ML3
AHpVi58C8r2GUXkRKujrDMMyKzL9Q52chfVXGeMMeW7+xcmV68OBiCJXHBdAJ08l
456SNzTlQEu11W8qsyWM7VtdLkrI3+PLCRnnSi63ArrUJ0IGdiAmS8WpPsSxODdU
kxdVjJH30hRmmOqr59pp+whtF+r+sc3nhKPAwphsu959ENHyap63VoNTu2ueh7a/
OQYchCHPr+Tgwkhv0gWs+Z/1T4S+ApIkg9UtjnxxAVNFmsvnKlYWyuLC0ZDpUA9O
wLsGF98WjzGB8M/vUNXfzYSOgCQZViNRIa3KT2ILfCfJ1IBbBNGGT5f6OrqiPlvP
0UE6iawtfIf6TuLveB8bn9A/usktNh3x/qLfZJpZJsXeZdbcC2YanZLQj8TR12V4
7qEOfgITxi+Wkynaa+hE62KH2y/lWW/ZaxzkNYyPkG3Brc/Fc3dtM7YheguDAX3j
Apcx3EfU6hFR9MNgYRMTLcxVgquPqtCQn0gtBhil8gKiuITxgYKMZTTml2XqVIVe
uFI6UPUl4T7MkEyxbdLryf3IUuto/Qsa50Sf1xPTG5jTGU63678GduTnW6yuhG7C
c/1dsxYVECis3Nu21RxTyMLawVzE0SumMWSXHfX/oBsiypdJJ3li/Uea8Vs9FWcv
DoeH3MTl+STaWJhFZmhTqYHsXMmIjSrrQRmstX6kacRBfzDgd5MuMnm1SkgwvhjA
GaQUfI94VDfpN4c6LrIj5aiaYOgho74WwsH55uCLUsA1F2HFI6RLyhmo11DlI9b/
g/FZJ6EaacgdaHqKT7d5KlVkhz8ZLAfZ3EevOy2jSbgL3mEHJpbdrdMUo627WHPh
cbDdvtNhiQ2rmt+SdtfRcVbdOMxsJhnDMO46OZgRZkzdPTCvbttcE7drv3A0Raeu
JhLuplzBwV8vyWUpOHQm98w8TZlM5xFjKqm0SwyEFiqgWZx1vM+z6fH0FqdO360C
dryinSzgIwa7kAi9LyABqcBIphQp2bKkCBKq3ngq6aPRC3iR+WxTimdj5QzSn9wj
TNZXZ0WBFNd3o5ouWJnBOmLL8sZp0VN4CaeXCpdX3SWtX931gAamnd4l+L0yt90z
Qb6E+MtRmZ9yPUEwsZX1HlcigPcKCKFhldcr4nTZDbmz/8tIBNtBXcC6UZBgWkyP
ekERQ/8OvYxe/z5lUDcjKvVg8t1DRUDBZb+YrZ0O4t1mlu9DZpxzavmBsSh1DQ8L
y2kDjb3R77K/mNGrJ4x1cICoE7/mbntaCBV1G/WP/m3rQh5u0m4R2kC2VOIH20ZO
3w2uKzqNGHctjBT/g2wC6QUOvlWVX24v8b7Z9Zh1btiMpsTxLIS8xPrU809kJx4O
ekrTuYr9uJecEyJuQFJMCvEHlmsPqZalSsqEHgCgeRiViW/Te/IhKlDJhfVsutww
ETPp4i1z7q6NaLLs6IXa/zDAnooVcORu4lo2CuSk7SRG5miNCFaE0eVQR4sgO562
gbdfnfv6IL0MBMH67MkGfcNaWn8VRYHxCee7eThvbPPbQWpFeqrS4UlWe2LdiqiR
paZvmogkGpjLb8/uNh/uPHqVUVWE9EvSsj+nxfzRlNF9OTvpjd04l8P1AHeK6DKV
x3VWgHCOBv/85xHI7xSh9CiZUiGv6fHUiwCjXYDIQdzj0uqJbzbZsb/8mtm93wH0
lvhrPuT5X0MeI1Dj4+LGsnOioyWB8J/z6YlJk7azu/ZOV9lUqxQn+XYZuqNS3ntt
8vP4JwC5zhAOGAAnY2Zli4pA8NS4Q/5b1dDQhb35NXs6VKl4mm5ya+QGAew654w3
qXWhIan0ElK7Y3ypzePBBszgHLoWbVaAHlqVUgyFFrKW9A32Wr2z2tCjofxFs4Jw
eg97TQBr5SqGynxX5VlzEuUyZQTplcFMj48Uhs0B+yyiW28texsMtKpKcIR/uPcV
aqSBqo5GVvjyc0+zmjRraDUXfPosduiv4Xjo1XCyXIK91IxAPAZQda5nAa9YZJga
AozgvDstqvFncdUqChoyvIl2hRIgE6H1FNypXa520BCaV3w6OYk4IZac/NzBCXxZ
sTg0Cn7idCwL6yf79UDxD8srq5I6e4yL2KwNFgvatuvSt2XmbJyLM4a039BHEWJf
op5T1tvA0+EcwjPdZzCYQm+AAGpnbZ47CJDbvA2R6PMtxtRNcXvMk0QcktggUxqp
tXyo5rTHxhQRl9wz9a6CEwoL8qm2wqz241zf8fIUGz9xqO25osCqftIxIv0AGrqK
ymQz6znnIXs1MKWAJpGuOpdgh0jTWdByewL7Wz0/S3LwBToWYq6lzKpD+WdS3HZM
Qd/wx8Gd2g1JdayCQl/NAUGhvX4/RmHJNWcWJOGmv3c5ncVeR4yuXSWyOtm3oiVJ
3PpRb5/6R3pSdSAmjMt2JLc91iy10lfebfqhYHC6Mo/i9pbX8Qt8xIU5oYD6i4qF
08Er25fFxFoYJo20rL8SZsgmTJVwEvBESwIU4sz/RUekH6gkfP1cZdIIq/0OV7VD
8DGzvE8fiepM3+uoj8y66PT7+RLlJCzsU1rp9VuV6b92/MIidcPDZNHx5Wi+S/MF
eLEel0lrRXPWJTXOhYxVlUxS1ajtn9oh2PAK5X9dym4DOFteTJeqJ12FhCl775dg
4uJMBPnd5uXkGJcwNTLIRlVtwVQ9Ov6t3EJw0l4Vorgp+h6VE4OYiA8Sgzntjc4r
2C1UvSjtXsPclZjvICMSAWYtvySPBXfOqRrxDIx3lnnl1fJhtU2R/TWrk0gs5poO
6M9uFTtT8S4g3UsTd0bJ5OQxLyqeJbgwxbrjoFAlPYvop3ELeCWJf/qqeVJc8Etw
UxTrbQ9PsVJS6dJ4QQRmyxHm7aOc7hFGLoB6T0PnOyrQ73RJoYP72rrSo+CEZgvM
OHK+GUFQBR2cLd9BznzeoE9cGtyGAXr+J3vFPPuE3t+InlTVgZqF8gwYYG086SZJ
/dUo7gxop/RfpVq4y6T6ZG6KH+dZ9BLWUpiJUOn2UZBuqEa5kGKRQcsTve7rXv19
B4+cal0Uett5+yjr7KprIeqbT6A/QZhcGHbf2FbRBsSRcAfXNMKWjQq+zH5Xq09I
wzshpfKPl/WLWl1KWr1OpVibT3u5LiGcuOPGRZb+syUYNPX2eZdvgnrOaedzjVoT
9CqZPh954Fxf3U4A8hl7+kNN0ZYwL9aogtgXjRQhisHwh86CFsKdbe5Jne19aE33
MJOOGKnc+9mySQLDxXYhTZwTpZagFsoQ/5SSQBH/mc9o6+GktbofKgT64T/vr39q
CQJRD5rM6T78H5XGjAmzkzAjPmxRzUBBDsMeQliHqi0g9sBPdQ2eClb6MC33z36t
H4yowcrLPjOjTYvM20sWS60t3hUZ2MKU3iYEzmY7mVu3CuN1Zn58SPSFlUDIZ4Kd
XeMxuMajbwb+hBdxYj3CyGWv9tAxQEc/aQQRjV+XHlJKv2ovzZpSwsGfo3rbaDot
lDwsnaLhKR4qHbD50EZVERO25+3wXWUG1anYOxcDNpr7b8DXNq7sSUJKKvE1MfCo
VdSPGWNIb/GEOL9BIpzrYtyokFAj+spPx1CaNH+RFEkWNI8Wm98pExQguCqidPG8
6GK5kpC43zXFdwiY2eop3oTGJcSVQd0/o27FYqcTZKcFJTQCJZOnZ7nFzx6rbmYT
xYLOk447NZcuqtP/iN5HGVPpXjhpfedb34FMkWi1GYU7mapS+30tS/3Y1KHntd37
8e/3tVhqAEXHUrHdYSzfY46CSC2+GRoOqrOn9XOc32hsOxkjv6U2UAy6trNd+E6d
mjdIHJ8aedJ+xNmT6kAxqfzIHdg2WVXe/TU7s0Rf6lhuJYBUS7wbRvuu6WzTQ+vF
9TeF9R3qxAbxk9+Dbk1WzpfngUI+j4MConq0GIuYtBGcFknBugPYe67It3bg2CYk
PDLSQCWyyGcdME3ugjYN2s7FLo9JcRbk4rm78LrINK+peAb1fY1avuPWrd1yXK4z
l5kt0EZHhGIxbhvDkLz3jtcoR5rHHj1QGgu3W/tBxcmZDh++YdvE1CEOdsL96kPV
BvQ9EY91I8oxTm5S40z2QrM4wg/MqtdmJpX9SxPpH6td0cMA00qIJ6metqx0I5/T
Qmxq7+j0lgjYHmhRs7h7suw3OyjYITQCIjJZQXNCXkfPyuDSr9KqAzjnUX456LCc
jF8W6KDtncHlKXxkr+Jolv9azkYOjH/+OyJsFHJ2GqjWjTn5DUGnY/zqGM2ADeN/
v5gyAsjf4YOlgpjfcO8EMZEKcphX7mDPczpUhX+dHWDaJ4gbyMJIKayBMG5MKc5H
iQv0dng/H4ofjT9S05mDUlTftnORYFgv0/TjdAZ93oUe/TYZ6bl3ftYqtfSUZ3ZI
JSvJMOJtoD9gCp+vVKcvmDTeaa8Ap4CFdTUdq/22ypC9MyT9feU98hIN5k5ajhH9
ew95SXfeM6pTCAdyP4xycaKu4ve7bK5PFDuVrisfZC9hQDNq0z50z+PphtpS0rV8
HJM4WmGivu2IZNjwAaO4jSMFYUt08Vq0QYi2zYW7i6kPRMhK/nkloLBBpYP4jd9y
oKh/PkUeoA4AIl8+RdzhKypnQ7/567wzhKlOQpmCCXRf4ee1ANCTtf9UohL8jCkK
6swT/WZ7ql/XnVp/PtXlLtYYsQhh9hpvhpmGIPydxHbybvaYh5UYLXuQo1X0Vpao
Karg43JvNQ49VDFwqlKyqJp/Vs96bwNzLHk9o23i6oT6f6TOyDqgCxXbx/pp2I7m
jK/zkMBcMop83cLzwuNRPa2DvKo7tKlhSbM/gpY4dPc3H1S+I5kESMyB8ocuD/DX
CxVkxjPcpnGoXzyeQcP0QwOCF00IhX802wlmUh8pI/3DFzM4NR/E4/nNQYY3e8Ug
KziKVJUpZ8T9E37aBmw/DnA3tkJWrshDUn5tJPVybzIl6FtADUsniHhYNJX3QQ34
cNzhoRvxJX7I1nDyA/juyyqZxnTFIoeD++WqiZabnsAyUnCmXfi111xe9C4Cz1yv
shyOw/GDc4TD1QFphg1xJx2GnphTUpMbx2g4hI3+EiEv2Pt4o1ufPVSH/od4Z/am
Jj2ji7aU5vwNsW29YUmR74PvOP+C5mZWWqsWX1KhGd/CaHd/5g/N9X4L7g/10Wt8
ouuf07ZcZzd3WKVVU4299CEsyeqB/kuT70fAdwSmDI8D+KhCFjBtk2kAy5MkJhtY
36gNUla63sJBWAN7qzkeQv3PzrZGdD3IgSeO3xkY7yOGeJLzKC7oa1KQmuiagmae
H7xPDb5Sjrkuk0h6Mvobxg6wVE2aSSY/UL1FByjUIPngGEuqrVdtHfL3LquCn0rA
rMjAY+ZNNxF/0pZl19xnSkS2h9d0mdlTap2AfCOYJMUbQJRdtKSyU8fm+XoSaYrt
lOiUmCEBProvu+JxbRh/ZErlRNQopxjd215XIPOmY4uUtVroacGcyJCBaq68Cpq9
GSvKPcUo8+nVLyVecQhrIJ9R5NTlrwsR+1RneOnIgDxzn+58upndjlKiPMxzKkWn
Gf/C4ixM4OrfRi+AVDAokqVcTHwfbTwXt0PaomddWupSS6x7OQ70NZK6BxG2wawr
SUSKLEVuuC7CjJeXJJGSz0mSYw0xF++7UHsWGsnUdk1POuaGdgKFaaV22X2af+8j
tXXuA0clKT6CaFJiqSLMomjpN2abN2iC7WRkPTsPpsDaZoN8dJ6UpW3vRgdgTF9z
lxCDNPedNu7hBYNZ7vlQxqHcWZZuDomYtep1gLAAOYWdy+Sloa2mMubehv68oejD
W7H1P6ba6W3lfuUI7POe4/arro/KBVdNvtHexshbBMB2TdCrLgaE4ZDhFGgHxDP5
kmzFCw0vhW7BOnC3AV0Fzo3uj75Bn923hGPAdzX7H7LyJ9wdePqLWUTHgXQk4XDj
H9dVs9DywBk/6SgM5rvuW5hJ6Mr5W4W8Uj/ktMgddXkYw9vtph1glMwclzETtnbV
YpWlkHikMXUOQbyW+vdTOjRZ93nf669rXJnpYYxhoSAYxzDBxDFUdFLWBKx55/Ma
BptDLbl6UEkGaHNtUsSO4Kad1c6y9QBv86rIgR8Nro7T6lmUnBzQItBs9WlYOU/R
eb/3KIc/4raO+g++2APM14GoLS4w0XngpZeHnHhjE2qAokirzGpopzjfGHK4MOmu
Fv1fQlh0I/LCJsXMILohrvy7cR1MhIID4eUvAIRp+hQ4URuHRpY7p+v9s29lCwHD
sdPw3Jnnt0+bdoNRskvGGWQ1PvfFQyAoGhd804qb/eiYSGo4hBMW0v39Ve5y8six
hhGSrpucoATSKdhELWXLf2giyg1o4CUQEOY1Sfjwb/cpyHAk9f8QL3e2X3z/Fd4V
eFYY3pg2S3CvheXoG5VdFiPk64KmdPZKKwxSjCp3Ef73s/bX3ATMsfTJfXH2dRiR
gyDyx+7Ae+QObUWCEVBEeYPcGpucmrJ7jKOkr/yYkE2n04AwdI9NKni6aTxKIdvH
21HTXDDo2SSp6lT9WlRjdFn8hhS6GCEinAMl0CsCnUkt+LxHnx97Lf/OvbdxtZ8N
o4Q3ZkdEbz/Hu+6roDYb+HXfBNzdP2NmQn9wNCHN14BZ+zJkZSZ6pPmb14cByuch
hD79cAefYZZ9cVE9Xu8L8RBceZz/TdKaWBXk+dwx6uzgwFJgIchFehtRrcIABMhv
XIf7GKRfDxgtXcNIKZOwVj12AXBJgBfcltVTyBWx75KwkDx1EQrrXBraiYedjq6U
BGqIAKmJldk6zwCqV9bJZ4bVx8gFK6HYaogqbCBl4epOJOnfU9Z/fQuiY5icTlIW
Xhxht9sjIkLG0lRh4HVSdWwLqCUb/gaBi5EJAT/K5hHRBQZb/uoYuIla2c9JH+uI
IWxEwgYMZPLnYw0i+oOBRuSIefspO3FgnPP6IZ+owDG5QUEZSICdVLihsHgxkhjI
Hs6uI5L5ZzZCOb+1tqiJhIaMgHY4nTLq+eNiTmV580YAqLydgLzuIl+4z5w9dv92
cM8LvNp3fU7Vy6tXrpz1kcImoVNTyen6xHQHq1lNd7cZ7r9KzW/rJHGDwRzM5GB+
Lei5h4HZr0iyikxLLWq9tbvi3Ssjw+n35sSTPJNLi1JCT+V41EX+n/fu+a/4Dm+b
JmXKJtQbe8wsP7At1XCcsSu4anW2GS6FCPV8fxRUwJ2R5eihdjzjENmRlDQtGGft
L41BtfvqOXUUtpiO4v1IIwcwUs4iEO4ZaCpiJc2/t1a6paQiTxArrEh7x5iqy3cQ
VwoP9j7QnHJWxN/ajAy6iEMpBWL2b/h/1bOkYIKYUxcWhlWeJlvev2nfPkrrezre
mGaVeQxqJHlUb8l5MAKZJw0unleSH36XmvtyIm3ByIxrvvDbEJdOIWtbnF8Zk2Lx
nkKulVrFTENmbzysPlI2kxfky9S7bOp48YWaZ91vU1Ry8dupuq46QZCNqUAbtIWy
BB+1mGqH2ZTxjryJySi1+gkY29R5Pjs9/Lcy/hSGajw7nti0Hk1AgyxInCkKatDd
hMDtebIUcEIBFLFbk/V1iLMjnVVEDcKiXzzLxlCpGG6sCixtJYMwe7Q+DAVT0Gs8
VnEyfUuULx7BRffxEp9Yc5PFvxfKg2S3w/UNtvT8fM9L7SGDZrMlkmSdsOKPzEYU
jBDC6sRb+pbQbLt2pCN0OFhWD4MaAPPVbioHxva3hJOINdqk0a00j6nAyzCLS+Fx
BoE0rL+b5cyu3WxQiJ4+0g0jsXigzjBAXYCdrl1HE1L5uwsaAOYbXsSQQ6cE9BUa
+IrechEpPp4jC+ryFHDJXFJyfOpuQQG/WUf1iK9cXlreo+bBk5UTy1mkuJuxa5KB
ao1BmizGU4Pkrp6CdoQrC1ze7orYcl0zO+UGJSu59UfW7PObayzTvM5PfsqpaEoT
8u23pBw4Xp42XUADBeGZ87lDsPljiK97KZaO4vkSFBLWMuFsQf2IWri2zGX3yrm1
p4E+SblGMRdr/CNp80fkO8jSQG8o6iYrCxY1MdMkOOAc1ch+Vi+Q5cUQ4+3yqYtW
hZEYAXMXFMH4dMQpX5PZqnKFjDu9WZ6mP36RZQfd4f5UhUW/Trn7a/Tt11dybaEO
9Z+0M2fDAjaNfpFwgqSk5xDcCMMl0yqSYTGnNadM+vGThvZf3GZNGjCeg57Oe9xm
ll8ecQ8KGj0IHo9JEtFAEt6qwVQuvZcghHqV7pUQd0rrdn4OEBjrY93zuuppUsrR
kP05J2xxrJNUQ9ZspA19v8dvrEJFHD5l5/oqNlOjKzFxp/8jxrvTViNISRGLJuwh
by58QVlS9pqnU7fu3RFIs9mIuBTwU+Oqt6EAzw6YG/+SApLvY+//I8ZgNS74ZCXV
0h9DuSlUvQIIdd1+4NglhlQ7n6YHNusu5oiOJH52DL1jUJtSRWyGaTfC2XNCi5Bd
u8tXdsz8iCYd5Vh2h7x5Ybi/YctF0vPAGaW1InJvzijEQiY7zDaEm3RbEPDNc8bR
WOLA4W9ggEPZlNiMwgWc99Cl9yyZCEpaJXcnVxdhxrvbvBEBt2IFHD1cHlK8OFp2
ZFDOhFdbEyOYT47oGsIl6C4cGDKofppMgaPBnHZy5TL20WO0M4ddJ4oFA8k62mwq
QMws91+rX/Ennwa6/gnoZnScNCUDTyR+bXiqq5GTs5wEO4k2xOE9PPH6heQcxW/Y
weZk/Ou1OdkCOtvUNWCeFHPEm/PdJp5ION1XFcGzLxcqtAQH2wxn56w3sQ4HKZlw
gnT4rpINM2Mmz+isj8sdXmUP5o2W+dSsiJ+5AAZHEQ9B2guXVWTeU7RxicOudzTw
Dy4SomD7gLQKm7qClaLAo7giCZY6op5++hmA05CnEmpIEHLNeduJDOCDOEiJ6sxf
bQv9D3qVzW9ICUSqtDwmntVk6dAJXqoozyHwunYF4V8c+3O8IB5QFmT1dk3A+APj
32nKqDiuqKL23Esngm5jN1YsCE21TgiL/aoOR3PjHg2iBnt8nwvdtPboHcW/FDf8
mH6gBDt/I963anT+BNLEfc9S3g9iHzFusNbeBsFYIN9oGMLzAurRQ2uuGFWtcVUc
LAQyUzqvBQZzfxNa3D6UV/vTvV6Nb1rePes0732xy3mMVqFQ1I5OJzgnsGagImNH
AmmdTyG+66vMOxwyFvUVejmTVF8L0ZiVRu4uUbSCwV4scORkD3t1JpHwKdDqjK0i
sgkqUwNsyGjcV5z+OyQndoEl/OQuHsIqcqEx/raHIhQ3/XcEjFedoajDfJso7HVO
rkJtIbrPq1AejGckkya+JahKtOJ3TtFkVbPbxoZxDFuTmfOBVVeWxTtNnTqnbp81
5o9aDV+VV9EnqV0cdtu24UQgUirbnGZImT8eCTHiMlTCtYPsXvVJKbFPu95mblF+
tST+NVHG7IDKH4UcrzR/HtuUUlFHpZOKiN2H7BCfIxSt2wxs02sW4pnVJ21Jiamg
QeLUcgl3qXVrL7B23zRtl1y5EY64jTn59wb0RDvL2GbaL3KhoUyNrpgU754+BmZJ
UnW4FkRUxg6doB9QpBFhWJALlGMEeZKxEiIEZrYERjxqsmiu2MzluE8Mw8uuWwHL
BOtxo2/XQwvq+LwTCl7oRjA40fwF17BaZTHUZyUz9LoNAqexsMiThL89KKntOZqc
4LiMUnyhlsHbVhpe9PfAJ9XLupukE2xarv8HgT9W4MzW02pcZbMPBnx+5b4dFFoa
48zw7R1EFG7egdJ+fgPWRXVmt/wzVW7V6rVr+lQpfT5euphp05IyBvm/niPU/mRK
T4rzWVCjopyDjfI1fJKMahqAg1PLDBrP6YHj16llo5ON7/9aIPHg7861M78cD0eG
6SXDsdXGCAcVucQVmx4oYAGTYyDP7O59faFyngzSLdsF8rbdVtH/M61KTMkOXDQ4
VDQqkiYI3ZY/XQ18K7Gr2Hbi2zBBxA2NWLnEZo/uqtk0RaVpHvwgUxy/iDmdjGG5
fW4xkomoISqQj8jaoZ20zZR9mKcueeFXUsqwVB010rdtXURbuw58x1stWFPCZOdK
1HwRe+JWz//nVeRLMVJv6G02JTQzVJsW27L5d7Un3KtTTDB0qIn2cqb4OiKGo80c
+jY72rIy4ku3jE0USopBz+Zx09q/nHCTaVMok3ZLtDTSD/kUML6ong9Rq8xcWPUK
qiBN4CFAFWUxaN6+mwhQleBuDjhtU3K/nTI+cifD+ZNGb2MKyUM7SWiruQrDkKg4
4Hwbn48FCZuUz355HE9DWst7jNkuQU9QednIYLTymppjOPrfPsCN8EIdxuDr0pUw
QQOUx7GM3uwaUi3pzBGzCV8Pd0r+2BDeR7qJvsU/+S/gjAMnoAmQXA2iHAb/QZR7
sbaQxULCDl+t7HzYkMDU1MBhjXr189Ug+lCiFouF7YW8kZyPPPiPCkwSr+ZBH/jT
aTQyhjDHMc1/6PPY+ErvWeGbGVfaAX6TfnhykHWxzfS0AX+DacAmXAOZLADsggW8
I0iLw9htJOHikkjAAU+3C9KM6bS3B7y8Mn2T+tWnFThhxBZy7roBwRXFKavKNlWN
LRFout4XZPw2xE8jOCdwl8VPWMq+IDYf/7p7hifq6WuKv5bWbfX0LmsbfpML9q6M
4jvOf+UzJjdPO8pM0AATXx9NTEhVopvq1VTl9lfzBN6O1Usp6EJR3FY44IdDIzKt
kL0731GOeXqrRYJWxJ7kPhpyc1L+z21ui1YvnSAIpBXrcD2DEe7sXujv6CoO4cDR
qhyPJhj3PNFGMzzI7Q2NSX2k15uoZClMszhIzBGSilJbZ1L9i6eswI9pOq6wid4d
LK6UnJ+DCbADToca/L24X2cIDfESFvr6HibZjXqr0pPMxrbMKEVPZrscByr9Qbje
3nOtnc2nYnxIuYIRS5DdPJ7lmDpHOYLj7aT13MjfCVbHGcwg0o4SrXf20/RG99T4
g25MTn0RoWClxfzLiY8B7nueWMJhFizWWkdviNl/NRqXKgw41PqrwlAS4S018Vty
ukRvg000B9MmgK2pwr7gfdR6tvqTfKdxD6R4KdlO25k/N3JaRu6e92bnncoULXKK
84a4vjPD7cMx54nN3n8VAkNXhP7WxoWZF78AvbrRUIh7aiGzyddwyZ53Cl/4JbIH
qpzLDLZqxGIgIK9gYYfmgL04MRaqWJScVbGnmmlSerJqqftV0vE1hCukE31nrNZV
f+KWVaKK6CALR7FHcI6aSnWlSA+iEycHCIJohKe973pJ/cEgHhxIWkE4uKQHnYOr
1kl0hLo2VVfKENIjzWfQwWZx+ZY1XLfkNgTq41l3Ol4/y93KTOi6HWSDjyzieswq
FRKaGha6Y4BAQ/reAJVlyaLhjdHIIgQ36JMFpjNWnRLaare/9d0qFe5Z2tnyUgf0
WZy6quGKIhX6UJzzOceBeoltnaC7Tfpv05hj40lp/OrPjtl1suQ23ijTW9soSkH/
pHmCWolr/4I1hRCtPDM/416hKSA3+aZ047JA09SBYcbUSB19peJDahVuZryXKpyN
G5IcanU7LH/6P5x7kYzkN4gcIb/RrizWbQ95P4Rwm+xBwcYMk1z9D/IHJWjoi9Wj
TQU6KhuBcNLH+DmZzzG/sZqyqzSk/RQtcICEWe0rn5rz0nRlsAKn8AsWO/FofogL
HQcAvXrA/INGTkQBM2yFeUdYesIdR/LdXSl9SOoRqKpM/RBUX6sZ2GrLY0uAOnJf
xJwpm8yeBYykU9FmbcsAFSrUR0csowIRqxMQYMV/kD/qHvpwBmgiJjLORAxhqyUN
2d5OS1Flu3WakAkaK3DTLJeQoYJvhV0z1zPzU22K59Vjn/PeXKqSFOlVERYpyA2r
9g2ypx69yV+ItIBZ1r9YAnkIHAdbDnhyVS9VxvRsXSi7TIb40KxKhR7ILtiGqtG1
/pAFSVXxaQTOTtyBlZYtf1tiK60VusZGe7rpgt2TxNLzVBSoGXuaHo0+9T/GYsku
rqfqM4nem8GjZOedTVomY1zS6tp34ytbUHLc6hN15sQrPG9xxjK/7p1EpoewMSPc
wZYC6YXl3Yh40SPcW+SfpoT5IT6joIPOTLSF772GC9MVaR/qn8vVXNKrQxSutTDz
4zJPtypuK8rEXCq8ZWSdLzNYO3PPInXDmpEr9YA6Vz5AEpIx0AZnQaTTtFWx3orn
I/aX/0sqwHkGP/rlqGq8BD3nmv2PRcvVU2q7m+6iczNtXZqo9cxUUzvjqAaxDQiR
nwbXP9SdfQeYkegz3W6MoCfBFsRckAELBUl0mpzsk2komnRY7EAc7E48wwocK81a
XNV6d+GEEtqMzz7TCG1M4HtD002E4OKVfdN/ip02E0wq6mRoTTeU2DY3wUUh1XYd
6y1tHR7lLQ5Axxua6G70/3R6gyETEkagX2V9jXRom37GJr7Hz4myl1Jz9E0gtwLF
KFzRDKbfkUKhEg717aUqVbKQvMgv7Sb3wnwgdDsU6BI4wH32zaOz5uLzCSgDlYvj
h3GtjD2YmZyw2QsNosXwf1ykpdf35xzX/4Wq9jfRC3KYAo34TC+Khou2JXbuJVqY
opG6Z/GoyfzrbBff9EtgTmkuYHznG3kgXadt5sP4JggL1P2zsD8M/OGH/0R3gJ+t
HAaeLQzppZihLnGXeYjhXb/c2R881IQ2dOVXXFpIZFX9K1wk2U7kXOMl9Ycaz05l
lUMAmvxv7eJ1ARmYSinyd+XnZ9iSHJIcT4/HkDVxjn+nzRcKAfeLehbd58W6OXQv
qXey63j1xpw6k2Tla0SMiklQHYhDRVBTFdDoFYiJ3Z2Xx/d9jXmDl8TpdWoaXNte
h7lpGPwhEfyn+1r++/bdA8CiuXL/L5iLQxNtNgwLjU56A/X4E02YWNjdqAXQvCVC
vNlVkXSmbQYb6BDceVfvwZtcrin5xfZWbOuGt8SXMvSndF5RWr1KHeH/7C8ktui0
X2BM6tcw66SD/3oUuDqfgvnPqQkGa81wEQxy3PRiS/2W70W8CPhB4puCy37MCGna
jknWTZEWVyGun85wRfGT0Ly03FXTxEj3fiyUUn0LJKTkBPD/Pwk51MZqaN3wcJ9N
uByUejzd0UizTx2NKIbvRza+g7UAdl9wE5IPu3qZQ1S2BqfFumQOYBaBaw6we5HL
QLVwCY6MvYnxaSIyQT+td7lt3/ApojNdEP5kN+x++cOpQExogW0+SM+43FF2CYUV
jxGaWVfzwo/WrVav+7VVm4b7+6AYJuv/u2338WIy++N3F3Y9nrJrwAf4PPcPnImA
pwWiTPM/CDT2D41bM4tXigYzZXdkjXPX2XLcGfcifHtqMlg44RCEO9QN24FqUOcN
LTrK5xt8D26J160ogbe9r41mkGQ1GOavaNBuRzZ5p5KX5V640tJUnTNGktJcc+0p
K20gi2riij6Wveb03P32ECy2joUPkyvDQFCimoDfia8RBdv153YAi3kaR+oAjz7h
2Xu7ZXE+m+PiAlR9RXHBCCs1FRcv5woR9yEOL0k7Sbasy8i6aSDV+uvFPnlgTK+B
Qw/OuDD3x4/xA67Nl20YVAavcpPZ3WnTcKR0tgNj1oh/AV6GzCoIfmBo3lampWeP
RKPfGgo/f8Q/XUsIMFNm7B8bRwFA7LVs+NPpaiSbPfWJWbg1x0gYmmJ97SWAXvqe
M4nMG+tYnf1445KF/xno7vQbtCtDZswPJcwsBGkvasje6rDxfloy97MCpQBU5LmI
ATAGFRW06GqviEt/z7KLyw7d36/zoZrpwVej1P2hECJTdFFY1wksM8tT/NL9N2KM
/g4rnD+9evlI0/D7L4CSIEEXkqcNOxbhqUIjweBFradagn4nO+kkQwIeDo6WvXyR
NrnWylgeMBeqiNFFI5hJ7nc7touRkM4DJLzKUfpnVpAAFXMqf2Ey4vgZ9amd0a8v
er7rV2dfPl2F2dbbkSRAj61a5EJYC37Omwgx78GEUeGBtv1QNqQt8/W8vkGxKGJA
DJcVvyyEyN9SQ+RdE+zRubDit7WbY/hVssTHwt/by2gU9ekKs0qMRWsCW04rAWJ3
1N2QM7+JVz0ZV/A5n//poOemQcD1ThivP5W/INzuaA4fyLDXb0R/2D/3XDo0hWC/
2RKd0pp9kyz/lj7eZj4K8jEDuRzhrrRUTMAZl5wr7hwwfMEbmxeSVFJsxR4fBhFf
nsPh0jsE4ryADDsfoZn5QYo9IwjabFzQ15mT8wZEXAsHO2ezs2Ikmm/xtXkZ1ODv
i1KK/BkHwR3iMNOF4Fi2gw54pmedNRUWmPu/e5stIvZU8ha8S8BaULmJNYeUsGgA
cK6R7/KRx3KyCLcnDOZtWszJOQ8fQO2/teyAUL8qJUvVbrkuPYIbV2thF2CwzxVK
+poT0aQxagkS+jj8VYk5JcdmfHuuaEwmK4SI/zEBd9tGgWTvYLE7glWrK8iJfZuo
XbyRXYggT2PYBjpPb0vpmRpkUInIMrXOM5iLkvrtaGA05tS4zU39eEfxn4nAkzuz
zT1/pcW6mTPlSkhP8Mg+bGdxxV1hbslw2YNgYo4iLoDvSSHjt9lf1scvwyISUE/Y
ZpXRuJmU/ipbes+2lTl8Z0UmSd6w3ITztjS2nldZxTiyUImqYpA4QTMfPSVYP1A5
jN6wh0mKSBlRDZDjkyC5dYi+65bJiKySSIz2YFCa6deQq1Vl7zGItiauQOraEWgh
5AmfHYGzOPblBq9zBSK0NZoSL1cv7DL3XYUIyw+Exw9mmsUuY6id5PTfXs5PxF1l
bAGOs/nyipq6np/HTqcwaCBCMBlwPWnsDTpghRVs0ezaZLe9jDQK1nno9DBTA99v
ZjS834QPq1+7rCzM8GMY7Oy245SN4F60jVg9Mk41yNOjnnd7m05Zwpe3eY7TuE+h
CBsC365w6DwqZhqu6U/iSKhSvFrVOSZq9Yf2YUU4/ArDoC9VMOW+T2JrIoVRZKsi
5G+pMhha8SZNqN3Mdtcvia7Lvgv+GxDN3Hyd1AheWar2kaVsvgLBPL8mwkbFfHcl
jr8ZtBBS2wQohimfEhno5MYPp8/lvgAC1JgG/HjwecYr1jRg78RD1sf41U5z5ZOq
uxIsTpAKFkMjKRn6VfSpkvUDbd/ZHIGs/ce4huaHNt2NIAliCrfHQfG1rPwJjnP1
9CYsk7zvbWZyWydtDmPVfbpC008k28idjFffUlRXW4e8UgMDIfoiGmRFXjFQIVZH
GHdDEtHonTisTjiIgPumCm3TTFM3dplORY2EUbLPl9GNlHpsHkXxvT6Qnircp+tH
Bzw8jWjgfT7WGCMp/oN7/z5aFGFr29M8QBhNOAuKdez1ycRtgzTPdS/3DtWR3alB
r3hC2EaVrpUFHSGaQDjCXk/faAz9KlVJ6m30IBO9EDUVM9+CMA4mP+Kj7JJ3WjSa
if5ULcWpHdCLzoHKMrdwlKv5KQppkmG4YeEqnbMNY2/HQQ7jjoSA4WHr0oi17AB6
h56QKLfaTu1cru4PdDarGmuN8XS823mE2pZ/K1CWhfoNOI70Bc+oxj80hjlvBgA5
vdPAdSXakWw/aqNhNiJrBZJAwoJB/t38hhIhUX11i1Kb4uwP+IOxPoxacZMFGUCR
kmcM5WHE2+ajjYaZoG5PRgn92uyPtHf1+0VHHgrFPVUG7AffmdV7T5TTMfXDEJZv
gqSk6GT4nN+0Rxle876tiW2AC67eSBKt/KVY0QzLN513LJ4zsjZ6CrSPAJCmMN1U
diemXfgPIOAdC/GZYWw9iFVUNl30gVrCVtc7w+g/v/iDEq1SdFD/Q/Oxo+7k6yOi
lhRBbkEvBsoFpFv1+bwJdXrmhKqtBLbc2oFBBI+D86FPnPOB56x+/TnZO48A9UmB
E1MiQo8AwnYonZxj5++utE8MiGhQaMhHTK9735gSRxoSVWfXW4Jf6eQ+jtKY5CJM
NHaNQLsNy8Fz9OP8rmm/zoJs9DJyW1EJWLLAP/M9LOtr15pmow0HnkFsJ5s0Cs8u
sxC2DE6imCuVr8nh/SzwUDz5VsaYucsehozzKEdZJE7EfygGKjRy/T5yLB4+Wvj8
/V33OndUQnwCJQAujMzCphp5tHplaSfWTrrnIwn2LDL+m9HoF+fBzWhUho3Ik8J1
2dCdGIL4FiI5pKOGkFWtBRuGp1Y1lxBG/YzUzOmqHnUDowdb8khv2V/RrDo0xl2d
peLWj8LFq6ojiVziFkcxElQfPgG6Ba8x7OYU/k245TEmXKYoWTKurAK9/SkJkAqh
LOkgVyo1XxRErZEX6uW0S1LkM6DvFSlQojK7F3rSeFvFWPLtfKLgWCOHzVD3HhQ6
+JvAKUkfC5gqIDc6FkFa+r9MYWLxhH7mD91TkHyjU/G9ybSui4R6NejZlTxMYo1q
Ex8CYvZSgl5oyEQgRSnZFL15PTBD+lEGBGdhMSAtC0gVYhaLH2vFdDMWQ0WzX3Pg
wQbZPqEaIOrHL/MxpnlPCPuHrrRzSZGYvXbEB/6vMl2QPRQxVPx3sPw+Sjf6uJeh
QL4XSKdryVLTdByVGQtaIQGZ8oS1W9Ddrs+02DnmG7m5NxOyXmiBemQsbY/RoB5W
RitCXqxld7zVkeR1poCRlGoArmVb1CjFuLBAWzdzxm0TuUoBwF3Ss9WFuZjM0xMI
MOJMWbnioco/YVIHEQRjC0YdFeDbOcmJUAvFDUTK5MC71TuJB7DIzIDJ+s+acP6G
ml4yZ9v1+vHrJVvykW0zOzZKxLcoDwHr6GvZGru8S/hNIgANN8tiNscDyTZ2J4Fr
qzebheAFvtJ5IVd5OehVYZDZyWolzBiF2OoFSTdzMf3VAlO+vjQeaRkmDPPDEjsQ
+pywqaAwdhFlAwPAbdB0jTPw1i3EDM3w8AzFCRU6PTscVw+j4kOyUL7ndLSjTj7X
42D39SIDdchp5bEzkboFlTpSODO5/Tlu94imzo6kvpdQb2iAmKjalOVMFflGFvn+
bDGldCpqPfzUAqL3cHeD/zPkJ4e4HudO970WUjPxg2SSwbzG65RK2zAd4GtJW52A
/QMfD/OSO+tP91gfx6ANIlwtASums5gNXqjCGzklTgC9YJcFBUrR140y9fwTr9uZ
q2QTOm9OeKd9Nbi5LRUyH1h0SD78r8Uje+u+RbbK9og7pFi0Ws1olxXxoWpXmqnt
DvVsI2TbeoAaZ2z8syx95PvP/qZmCsKdwMjQyT/t+22SYAR48U/KzEZD/IpcCNnV
0Y9s6HiRwo53zE1VNIMFCwNLhThTl3J/4df1L7UV+J3l2s9YupNl1zxvWvgn7Y5C
+LrJrJbXFmFMTeUjvtm2HMIr4uteUqGaN1wVSScgl/RbML0uJCtQQtAJznVZGLuq
fUzCTqzhDr7u58byzFE+1AZRC6BOYlJtUh+MjsBDo/ZZk/F4iwgFl88n8H4xLAxI
UOQhQxnYYu1NckAoL/HcH4PJZuv3Q8NFMByR7vBGDCtpNelVh0T+jdeGihkLXQMQ
ZVc9guK7SrD8QjpgSlrv/4hEVnc5LADyDb8w9qFgz505bMbDPLx/5PwjKa7PkajK
kGg/G8q7tkfhN/jskE1Eo1psdZCjrwHy3JmJHmpX3wQiJYW+mv5ghWtIub9Bk/lJ
HLPgjjDzy/WyrqhbOAO0UBfXiZevzDSINO7qzqjoKN82RdwK7qlpIwPBadDYrLXA
+WXAdHUatUtYVUMzyYiyKAACUT6bKkdyAMT/ooMDQ5oWHJbRz89PiASSSkHaYbe7
XYoH6MVN+q4mSdv4YtyOwCeRUqFKqwfighYk/1JoFBJ4UC1orcpjP8Tw4N7a7SIY
itpLJMERMkZMGf83xr7uik+LuBD2n0eeypTQX+2diNv6rSdLKfAdGBHGnl4OyWeZ
guV5ulRV9nylDzInavyZWu0wkw1XcnTtRbwiaRjdKCYbbfx5QwIbgBmtw6gch/bV
oOQqMe6ZyK7Hxp42OxZxA0UmtxQLk11TXAIa+ent2oXnpCwsKz/rFzkoNzbBQ2AL
CmDayFPNNDLGnkNsnHV8ZaVAvy2HUkua+1DXqS46/jXHaf4IPmHWB9Xm1OqQ3Wp7
DsUR4knZhooZ1ks2gj1TyTr8aKPtkcTJ3YeHp20CUOgb6dKD9dntrey1jjh59KoQ
kie50YBjQXRcnRST5Gk7aJP4zlw26bxhooscEy3FBHyTxa/vGirm2/3iGpJXtBxg
/EaJBZ7grKHlglhTCKjXabr13DL3wuxfFg9wq7X2NRc1d4pMYDXvN3rmj7vioilR
oLotfi8nD3wBC+RuV3Y2AE9kSFn4vSSICYN3t6GFoEcMqMJ/L4vJlFpHmRzNGFOO
lXSvlBMRAqUqGBlO9+gSPHbpWC/zaR1BqGMBASNQi2YJMVhXxgC8vIMi576Fvu7V
wrJnr3g5yAe3RKjzr+nijwiTaC9679yQEFZ5PzgsmxxwhuQu3CzOAXViq0x39S+4
zPp4nNjmCCD5r1dBhZO7HIJjXsOYlfj9AZ7bCDG74tes2a+pHTnEeNJfMOO4CjGq
PaWfs8RpaM2bZcvOLvya2rJ/NKtnn6qviNm3I9V11HJuOC0GX/7lCxkJdAlx/FWD
FBMqO5TOskk+3yvb/7gebsts9xt5U4DqNF0ACYQWQLn1b1Xj/p9Rk4LBa4Cv/8iK
i3wqh8eM5vtzWGSZrWciFRhhPFPafnanEw4r6+yI68yYqofCLLXC0MWRKIV3Yvm4
VapnxrxHcbxftPDDMoWoAyvt1vwkOVLsz5OgDS4L1ISysttomfxTNxHRQ5XggClE
hMY9KUrn9wCT1xqUOw2McMQ8lHvrMWQoLro8gmVG+mr8kn8EkvSfu+veS4NLRrPa
aaKUbO5Q3vcutPFZxw7EKiDxYonHQAkPiz9tvW43+RUilWjFhmWMytK6ePewPCLI
1CaAltWKtEznfjSYU0DaUt3tpSe/CSZUQxDSgz28+nTcIK985+p3zvEPAey7ECkH
MO4XNdRvfY+xwzjYJWrPgkGqrw5ic/PWHJM+VZ4k03avmaV18QMN3lwodYjjM99k
y6a5gj57GYmnd2RM9Z9svuGzSMNQJOiKtzW8XtHJhxjukrN7dcM8lQL3HldaB/rB
s6UFg0+t+8hzQAQqHjM4s/ygyJb9tdVxatO2LLNTgxYWm8Z6ZA+TRgiJSm+Qe7jW
YEi72yYO35KX+J8HLK3MwpLPEfdlfMIu81qzLgyt3HjGekPrDejYAz2KiFDSYcBH
u/FBiEAeQudqSOxoV5brdA4Ze7R1VKOdthUyVzUwXBx5hZ83/9Q1ekW9G7mw8nZN
0gOhg4mHf+S/0Bei6+/0Gg4vA7m2ijalxqO/MBgOP0T77IXHVrEWqqr2BIO1UEus
jVW0tagYPXbyvlCnReG6oQ7kAqKMJyt2TMKgb0ld+fOPGKb/B8iM7hqwaUG4PPQh
n5GyEosemlYYfPQ0b4UOG60xPHIWsrcEPb07K7LW37caoJzaueVD4m2DwwiUeapR
JPNw0O0Kz2/kSkgXPxJUqYB3SkCxn6Uo5rF8BrfQ3Cgfkj2l0nVg6Ap6URcNKu9L
l1wGSxt3n96EmhOlRPjpHv0aLCYclF1HprwXoCtz5C1sHa1QCk8XY5NzTmZr5tKJ
2Ke4MOE2rPY3p3I9lFe91jOF01LESpIK7nPZtL+aOeih7ClpNvHhzkIxYbPq3MKM
lHxV8k0PsKgAH8o/I8FiXWRxpWKr1jLeZfpnhWccqJalXx7MqcN6guRMHnywf7br
YcXlnWLKb88CI+nFnxTpio4iQpyg5KItAyaaKPust9F3PsfuUy5p07EsoRhzO/CI
pQltLv+9N8K8xQfXqom8fj46ZCkqelVVUBbTBYbyaO5Ot3v611gHlatKrlLR5556
M6J9k16HQyCdK6FU9JKd+W4vzt6YmU61K+R3GqWRFeequu7dE6hCJ/AoPe7+I0ag
TpqgAsztWSsCr/MNpGM79IqwdQMWmd/tpcpL6aXiq+XpnEQEFVu472muTUa3YHZk
ZDVHnVJcNAgYPFJlKqDgbZnqDl7HbN0TlNKDnWPe+8fn5QGGSqpY0ulCyf/6yW0E
6GWi7UqB89+i2wZO5ZVEffaG4vvPJxI/BiXSRhUabKx+f4EDAUp75aflZsNSQyE7
8ww7tDcVeM4VtOKc6urufFggcLYK59T9/wBUtI25eJPx9hmR5TGSH1PMNSE6w959
EFJYpGZ4YEL+GwexHtiWKw/J701defoVXMgZPFCm1c65aYjm0Vsd4gc2E6RkzI2f
Z3cgqSpG5TWmB1ougvnlXF6DfLNMv7mXF8w6+rv8RmOXgBxD0UbHjYDquJihCDU8
/vtptPvWEktYN5pHCURzgPTDgHLAEl6CvqRyxT19GPBpY6es+8W8E/7C3/b4U++j
83zs/oC94UUFZC8buu7UHEbdj4RKr8NcnCJcZnkDPAvnwdowXg6D3NJypHxExLoL
ouA5JyZ6JAG/3T4nJxDUla85nVzQtbfWBfUR/ulQaWqlqn9FsCJHJ0L+MM3IP77x
uz/p4b/rVu2I6ans683m7ePkh14uW3S12retpq6FyElsLZVPAVQR9BJV10DLcjW0
ui44WuFuOM3gXGK2IqOUbss0+tdn3Cx1tfOdnEAI/XEQX1Sku9cmKUjCeaFfRY6v
hf1lBlI3HoSn4DAMdwWlCcwN0xoPFJk0cSqyR3MlH31o/8nPPOyYaUJNiI+kUBER
vWuy4XJEzgSGWlEUrk8YSD8gS0kWKhVJTWZ4q2Vtq5yuMd3vjcFbg8iM1fsoLofK
vwe5SL8LQ3HK3n0GiKh4TY45qNVqa0ZuCIrwVN5QivCnkXlkxlcymle2RdjIFTvk
PLfxE/+Af85i2FhtKRbG224O/82VhGPvb4H3ySK4tlVGh+vKFBzCe4XT2/aaBsdJ
FUxtOVQ14i1ymyGZjYesLAPXUi2szUlEN0Ly33pYL/7OVAtKon37uoqsdg6yzVkF
84M5ftE3UTeHJVDqX+KcdedY7g3tH2sJqwsKG0LmV94pDHtVaZ+bfYSNyBPu9cuy
tWUG2PJsmWrAGcbap3qIJpN4a2yHxHx37bP1zSnprzzfgX+/4CxMnpIhRzuCfRr/
IQZRDUpDq5FJqiaAJGFd4d1QyAXqtzO7HdoNv4mdZ0bUWInya/xIrwIwwpOxzoZu
rYezRj0OVSkAc3eZOY2OYwKyp16qU4JuXZW4TWSWwcwhhWXOCbyZ3Ej9PoSLLdP6
Y9V2abBNSs2DoTaia7NuPsYg/bKeHriDDzOCzx2Hm1bHQucn3IgRTL7nFjGtzVSI
/AxkY3ro+ZfLnbGeQtJdM85UpfETa4PLLerg914YKm2T8C1FztUIWPeZhb4tCwUY
PW1scMSSeTXkgHpJcyxjPIQTtUO3z5B8LR3PFbpSuPXPsyKJveCj7eXuKRh6tEYY
Y2PTcOg6KTUIfU55c+qfwdGep6+3hOFElI0eDVFvHURXZyE10/767p7H0b7KU3VZ
YcVvhtT0MY6WhxkoYCZEjbGH0UTVLnczSiZrpWgcOGOz2Pxr+AAt4NBg6iaGViIK
qbPTqyb6xXs7EYaCnddXw9szvbHhliVi1lU4DNAy+xK6G3HiWuHVfo28IB/OM7TM
aoUJJhKOd8xb/iVSw5CelCoABl49zbxcN6pu1bxtJQzUqvi/cX5qaaHQtU6IHiOK
Sej8S2baQ+uysbmvbnAqLNr02aq1DN6LCa4s7N1N4Eo5T5MCNTwI4zdRo+3pSnn2
jXQAiNaa65xUELCjom6esyEmwrpT39lwZIxM1KS4/IqSP/OoX7IF5VNICU3cTpJL
nI5bTl1wB5ZUFbBk5rJf2vorEccesoq3KCuCopzDz7YyeASLzT1bGASAQm28cpVF
bARWXqeQhUFIg6NoNzYkT3yzLVycIzqBG328FCUEdKp3P+hAGQ0btfN1mdgEjEY3
s1Lei9/3UBvtvd+PTP0j471CoHw5J6XElJ5Wqjj171d03ZVyRYsRAbswgMKTsW2I
BbLdwFfkrElgGMFbuGmDuL3DQ2yydil69rAKbrsMY5wEZYMT9oOBCmF1eFCRugOo
SAQj8AlNUZq93mP9kznBz5D2+F0gP/oXsqYVFgMFuF9Joe7gf3MV4NkrBQ8YLcSw
gYTVcgcR0w9Xj9B4i4hHFfmdZK2m6WvRc+VD+w+giWVmuQp0okVeFHmuKSKXbLIw
+Taczt9LjM6GkDwDOWL1ckVMAxY6v1HapM+2sM+bjdPMbCEMNnnSTiRF2rTHbbEW
f2UTNurI15gzUPekR/P+rIi247uMNEYo0KcM4YSXCmkUbS4ZrXvd3CIcLhHNPaqF
IdSWbl8h3USOT8pOD9qsCqHZEAdvRLWUlOoumlnfY0Eyx6pmvanpfzMnvO3lfvUr
NQYkzhdwesHmqWSRGO6FrVWy9bdFyhyyIBBSVlJ16E1yuBuNCqgC9BNfZSBZG4U1
2G1goishT4UdpyJ5Xr4/sNP/Db1JWxVxvTk1TXf6j5/fQcNrrvp5om+Faj5oy0JB
xgrPSxZJvuNbTzdhFqS7yuq6oGZWRZVP4/Upg1nAtr6F9gL5FeTVucn+Knd3IgTp
uA6eMPcdDNEpHb7DLAz34fa/wwltEyCVtdVsUR346wjKHACT0wHB/un2uV0YqGjq
TKBZ6fznG5rkslFrgr0pOrDOl42srb95C3smKC8oiYoWBQVbeVC9YDxWQ+e2ZR8F
3hzsZAmd7LwHE32OQEtVLpXRQ9BjBAVBGtS4rP0VaeUE8KL4CFR4W2RDiCb+0GOt
1G+mCw/lgO5eilr2D3El9+4/CSSsfUGzGNfwPdXdTqAyq/Fy/j1CGirZ/gJ3xAsj
PWTamkzhn+Cn5jgQGKjIPBCkkkjHFrONo3tIEf6Yqwtv0441NAmCQyp6uW8jGMHL
0+lKh4G6I9USJQ6ejVjhwVtagV1iC9iRwcc6MUnux1r8JkBbapgX+fhW9+S3P1aI
1Cqj6QDSLQje9PtKKwSSLxw31k8ck6LTxelwXyZzc18TmqPeTl/V+1YKVPUN1gsS
Pw5uXmvf3tE72m+Zqq5mnuWlNviiz17sKFJhW2Fzyk5Knv3bSUEZmFANqrOz1Tqx
4EgXVc7/qMS+g/aDE1REyN7K9DmAV3VZvJejhs8cZkyHK1QVc7bn338HuQWiQ/CG
mj9//NUJSp98un7P93DHk4uBTk2zkc6gbYgMNnpZmm7XU+nlrCn9UQ4RMcat5w1P
vzP78ewHHg7i+je11MrBooZI8TYMPwihgK/Jidi0ZffoNCBTGkY/BjxlKJj9MF4Y
XNrQsSOhdiLBRJ0BmrzQWgHWQ9w4jIn09pNrAq/6j9WSn/ZtY41a6VEdGvUL3rtT
huP3Hsb8ODqb3O/9Z3YCUS++PNjidflFYQk+kZocPaqgo02KOppYraSvDQOHFav6
t8BbgUre0VZQnaWTHed1kT4VJSSBql2U4SBEqbzXrg9oiO56ixs5saOskAvviuVr
5/Nn/yK3L9duvJcljIbxfBPFlss0EEz1lsfXMjxRg/Jb7aI7ylWsSooIB/LF7MI8
PkbcpJloHWhxKyAbbWiH4Re/08rcKPPNthO8OyDZStJlJv1aHQNobmoXhgWezog/
hHSR/QS29LuZN63IYcMS0gh4bgNaWgftgKYb/1bpobyqdeXypHGQYnXJd2eoM22M
GBQjhB8M/DKs18TvVM5zYfL3L8P+31ohDJafW7TgIxZWCDDmlZiW2meamOruKuuB
cjHR5Awvmjp7MK7qp86ztxvpDE5jmFgIcURIITrLs40invc8atyikAKOBhn7H4zv
M6M4P9NJcN8bwyFK9emOreL+5nFfsvCaBbsUi6zEpj6/9alx1NGnRFmNLoWESqBp
8AvHpuDJl6WZvHc6gE1P3WxM80skpVaA4/trTInYksviR1EYOyrkfBg7NPilzODT
8M+dRKjrK1dlw30MNrq/qJnBXctlp5H6wKXFL5CBZJ97Yu8BFj1soe+int/GeqSb
Yqphq6y210wPUVWfnKQhLAQeVkI2bI7jQaIi4M4aMjlwWdFG18yo+sQ+0lZicn66
9m1hneZkA7+XYgLH1D1ZLzp0SLzEC+/rvS+s0jwNVR/zJw3khJeJK8DDDn/l5aFn
7Rn4QLj8RILI3yGQ9qxbQftaneQzS0G3uBDNR9B/p3Z3Ls/CqzPe3HqUh7yMzGjK
+tlSuVqM/ITaMVIw6rFN6kiDCL4qk11VDpKBVNxZD9O7J7QUarHUYqRsCAZWfNqw
lnBKefGy6Qo15V95SDSqyDEro8SQz5hdK2L6181Ie+kHnWESRkjZlE+tr32PsBZg
0IpzaPNpV+/DHd4BeGar0rpy39tioc1DIgRZvThZoLYpRk6n1+odOPo6Okm+2yiD
31eF9oIu5r9disi2DNIiFKTSq0CUXOTm02tzva3jjxzR9YWxk6hC9/VfYMUsdQUF
5kYi00iEt8mhR9Yafwn6dKW3yVvlqQa1NQap7jF60qQo+KF3IZkB182fM11zakvu
AprAexKR1mL/ETJ6NTUTWcv/ShNYuwTdHeFm3Pu7LvZFMQfb6VkWq3eM1Zyz6iTW
FLnHFhzhgDEBccYuMIHauneu7iIgKWTxBQ2lGwLMo7HTt9c8EALH5NCSea+7R5nd
OTJSZ7zGl5IwVSnTx90VOF0RbysgFQY4brHFD2s58g+dPD5eIjbblX6uXfzBZT43
gm6erF/u5VdXGN+zsO2sHxsD492EKLVY83UvKpQYfLz4DxXgX1YmFaRI/2d8oVPp
ItnrrIjKPmhS7/Zq0RRuUiReQfTdwQkXRuzqhOGS8SMocNmJmoyJLduC2U6Zs/VK
dtm0qYvwXPGfmaAg7txOvSqZx8I2UTAtYg9pHcICAZqcKQTXDirgFmVITOSTcQMz
obUJqB3zy+u/zSsKSn6u0W1nMldlvfqwnX5lluLcseJU5PprxxwAX/oukZgfjd1q
/iivARl/U5NLXIqS+UOXGr0yn0kx4YeQ99uT3IjxEPcLOVIl1Z2RDdDPg3PHQpjP
ddd0aq0KIhUXNruEU246v+itmokMlcOclTI3bPVSNJQaF3J9veNkSjLEmtpkXknZ
G1qInEXXzTplhrXpKvzbzfS3rDYofHop7bdT5e1Djv7g51MZGbwc3d2hqZ2spHke
5s/TnQmCCNCd8Y8lFqeewtetSEFmyoDMksyTFxesUpiFtTyc+1QgK4G0nYY57Kjr
u0d5sk1rz4t/K1Kqm2PrDoGF7EuoyhqyDMf7c19XiGI1rkf5mRFIP6G5KvQk2tGv
bhtNa396lvPQAxagbPmVHHaon8acWc+G9mlzrNk15e3A1SC0Uy0D6xztuoidNay4
9fUoV+yzmDvWbgTaPRO5fZyK6f5HtbGlaC0/ux+4cr40Qgqt/nCSNDrHoMqK9ajc
SAkZnhImb2TcoNeFCLTzHGGxLR/hPpzyV+6Etg7OkFkydu7msxwYfats7s8hrkn2
Li94MXvBgLnnntviPV3xGRt4OODx9QOeBYyTj/YoFXHaZeJtLMA5ecoLk/llJCGT
KTAHApzyIag4GnsK3tpE7Qx3Omp91NLeM8oySoTcS93T8eZOeYJSBpeuIV2jHHOG
XHI8ojNCf/D0sUwexKJuFxzyDBx/TmwUH//iKCZraosfRjVDQmLc8hZBTxQCTq/M
5tMVSXWgn3SFsZ4Fuq8KGycvKGFIg7H5+l+vF9wIZ1Sj1sr9Am2BhhKXMDn/fF4B
OA86zJJ06wrTkiWXZVI8Cx6WZxQR5B+cvztP9XDtV9qmogRjnX4v11VhngAuIVG3
B8vy+GDY3bNcTy4cX3pHiJRvUY9wBm0wmagSsOfs5MKtVZhlxSwHloDepdnLb8a1
RIR/1x3ij12VrdfWaMQkUUr09V2G9UWSApwgTmPex/RTdQN3IK9t5/f63wCE1hnQ
Hj7ZxTRFpK5udJ4ornTvk+Jvu78CGByJc8EINLVngENnbg9eQWJlONA0UzW2cpuL
QOOtftCmZGp6MCnSbcO7NBZGpH7rWEiaexqXeyVOOcZ8UdNSZ4GdrG9vWlbtCyg7
EeWm62PMPIOAoUwtFRt+rHk/ohfO5QrTBta3+Zpbj/oGus0pLV4OTtuvdoLWbDHQ
BKC9JYNB6BHAAXnmQYQoUt72rkS6KOfHTeNF2lqQZgqA6iiL99cMHT3Kwa8k+Dc2
+Mt73GAI7EtwMoKVMrjHLcyAc6jIJm4QmrmTwRMEiJuNMommsf/SqZYEHSbHkpDL
z0MsRtswx8R9bvl1PVDCKq179a6sPcoCJzQ/mMpfRPDry0yHWNnbROGTUAIpTWuF
frqCVZtCG+a8i4IUBiqJmt7j63Cg4VeJl3vYUWXNOq1PTdKDlhDSgw4UDWWpjUYL
8qThkjq+BFuxnnoefQczAe/2FxYoXsko0Oo2EY9WR4B20cS4DzXmB2p30/ShdSOG
rUZXt9A6/qgaG6gupxCyENLjDsKXYri7e1e9yBedIzH5MKO1MILfcZuEn1HtfqmZ
FEQWHPPuv9BDa+rWS5hPAYTR+vQIVqE6bO1t1SSqoY43b6+9TqWwuOzLhJVFXVIz
6w0hla0Uh7jUUzjTr+nt2E83gfwrR66pJAL1a06ceoyWl9GC2frZLWGnZ7kPN9+d
3n/wHjz8pap1MtJjFz3vpCzO//Vm+8BPdQh/fWrkBCmU3Z+CVnQkg2yv1EbNDH4/
Y7V1WCrHrYgAhx9qx+GwQc3I2Ub2/MujjFiHpNczB481YU942RYvhHdjqOxybnvN
qkGV+XfX4uO8JP8Pg5eSuk2HiyqACrD9q/C0coClqDWsRd9oxe1WIqCjIOyviX+I
jV8pqqdBuh4rKquEuwpF4pqDR4WRPqrScUEnddCFb80EQrKy15SKBaQ+fevg/hZF
j1gwmuII4OrPCbVNSeIsMNocdm7kDqoXM0kR/750JSgrn3MTmSzrM4FLmmRl4U71
Q5bEmbVrF4ZiYZ70JO5DJnkGkLeU0mw4u68fL3lKHTezUjoIxGy1btSJRb2GSqs/
JopGyAMG215pia0TFqW2hyttzWhkDOF497UF+zoPBxbkzSGNhNcCY/TS2CpPwgj0
USy9lS5wn9TNyPy4ZBxIQq6YCNkYO5y576lUMGyiC9L2vs/oECa2lv0Pn1Fk3kzO
IezbT/uerQOwaq+ZXUN+A4V87h6KYB8A6qLvN4MEiG6QcHdZh6Yat+P9w/BuNx85
9SarvNtjnXyQxicAgv2jpeysAzkkdBYfX38dYj8YKzel7n9eoz5wf2xZ9pDo9ada
UWZGR5CK9hK7l0zsL+u4heBpflBDbfDeS5VRYOeBW9GLcVzTGPL3NHz6l4iojOiO
DTUenxQY+QSZFMnO+D/Do9rBAPvVP5HODFvxQh71GObXq0I26GDUnAmfRseaklhN
renTRuEHv1AiTgmrtU7sYf63VAsce9oFgO56ScbnhYi5prnvnfui7eZp39KZacOG
qVhi5NEahAYU7FYsabqsRYhLANggiokXvpLh2e3hk9YayaV2kLVdEwFaliNr8yuZ
vmXv3eAZVZjXUaltAmaOkn/Fpcyp16fYrWa+wXrkBKM8Pzu1mg2A2dAOaPkxHN4N
KfmEWS1kwL34b85IlfRA1S+XNriI2nO0p82+wEeIycyAHcK2wX/x3+TIW0SxadoM
AiR5hhKSzTYCYgqS5l/k6fJ3pU+eYKGgGTLDXVvgEyC5IJOnWbPTte2+o303KBhZ
nCFZcb5Tk7EG6cYroLaE0QNLibaan3uCbxRM8daxQmqNGtasqeHT04dpa5cfFxnJ
F8rd58s5RRxAQRwGh8QXQElkAw6UrDMTG7bxsWSo+aGAHP08jzFY8tkrRdRn/7SM
EkZOBF+FQ49ckm3qgmRIlw22nGXObiNXPe30576QlTniRZysnIQleg6YRs7nIeI4
ZvZEKtkBHKO+piZ6k+G7rpYNFuts0Ufb+9d2uWSJ3PKukxaMSy4wKG3pedf82rHi
Mr279ZE+gTbT4TNd2n1L/IvRcub7ERUdznV18xR1EE+9V8nWLsLjbEE49K/Mhkl4
TFTei8QbcoyUL5Z9lsbj6xpcyDLMPqLBgB9b1sKVHcjM7g3z3/mPxM1zOGzjCkKH
LnciEjAe0OhhkmxZk/3AUnd1NbrcJqgOLb3IOgnuEaaruZYKIoS1PJ2N2eFsar6e
nf/wx2m+T+lNlfknkiJ4YSONuDrVJVJPNB8hVVAo1II95gUtHauLIUZJZpO5Te9Z
ppjCA8V58zntsHUyG7Hr0Kn9RdQ9Uf07qvA7LTnU5XQXwG+3VOITzlGtqi6ut2WF
cuYVktSFGKR3QqH5WTIZsMeiAisIhOCPztCBz6V65dbnCHmPn0w9y43cu3oVYMsz
tKEDL0MYd9x/7TwuF3YV7osGniXprmAXxfnILFAqZ9Is/gTH+vxWpoAFFrg9NE5u
UDb1GZfzIuioAc2A2AIz2AU4viyCMN3sUHqEJbyOGOUMgRH/T7pesm5juuzRj1uk
ZWXAJRy5J4deOQR82rUDI5ahVE700H+fFd2WjBKcyL61YFak8piKYyLfupmPkY5f
RDZhEAfp54tFvFPLG/zfdpNPAIkIsSvXD2OcpUnWSJjiClIlbCLWmV3Hfx8Bbmu4
RU7RjUDNrnV0llxPn0FO10KABu+RvcNYBgaXBDqe3SgnhBET0Wt0/YUpFfarJ7fl
x0NSk9Tgl5BFDhBDwDQylqVLEn+pVULs4F9sarJ1OjnQnpKZvp2Nbq7boui/KK2V
kPYfdIHAuLRkiBlzkbSSfW7Sbv/4edippU2Ox4sRCP347CsEv6GoDpPCUicPPw5a
6OrCwIeZtSylu3mxoPkoEN8m7lrJU6Ju+3XUaXyjFlb5E2jdUdE/EFGgVVeW8kuU
ig8+YCoNnhMnhxA6MYjm/3nPcc6to5undrWkInybp4AHHQlHBOTRhhDFAgXvZ1Xe
jJbfkDPzJXRA7iAnTLQWNvC9QRzwyrmamjk38GgTj7mYu4DPj4QF2dEsnQz8MtgU
XX/BdWDoBkL5CTiO2xObjzshihxVeR6NMlksjUOLppKVqzZ8I10KZY9gpoYBEVJg
et7m2zBG1ug0rZ0yGGlsxFWyblrZBdZfXxEQ+sFax/gA3kc+KAzAg6MriSAvfgMF
6p52Vq+IJjy9gcivE3Umo7pM3tSCh93lX2k2d4xqLWju1HwrxVHDqnHMuHWHbjDC
oCuzlryXtoza2RZCVt2urIlPsPn5bzjk55Lzgz3VS14s8UCKmw0Op13uyh7n/Rwa
e7zFiDK/QImbtUEYpUtdcse7alPhYC7qpP7S480c3PNtX6kUBLiDYIzmUOF3gjSy
SR1oa8ZJoTy9qyPQnq2EceO3jeWZasqHpI56rFMvCrumN1dFk791CJSPM2Ca+pJO
ZzPIV0xSrOT6GS58r18XOuVs6u4l/29AeZqn4ADbvJqtXh/OCCXMa3v6KDFx/vew
GcCumwlXBZ1NkXUMtnQt/ng4o33NZRbtDcNu8bg6VyTCWwYL5Si7gpxD5Ot9iq3v
HCeTC3+f5v4uhr1B+AIwTObu1NuvsIInk0Tix9JlpAUCQHJ2u49PVPr/Oj5JFbO8
MKN7i+qQ0X+PmyaasRdB0wIUdOGv903bJk8s+HdOaMEfXmjwCisubkVVFopVsKGx
9DrU3/a31F/eTrIt0iv2C5yJF85ZGsLqJUV0SQPuSw7hXBfDjI7Nh3oBWrhGCnjI
dIB91dofunNrlS8g4+XltRN5IogEiQG9ds03q/w0R3U0thRSNh0T4tpYFqS1er6Z
f4J8WgFAcTejkkFSrCz7PLHJlVRbTi3dtiRC4dIhIKUltxF5Zmh47pymebA7PTVH
tpe4u/1ZMhIVIU1KfYIWzLIEjxE26yfJ+2Bv9y5pqF+tPNyn/JtOR2zIoRxm8kOE
51VxJllApHTJpp04jRdLggAxkqfDl3OJ2v5/JuDebG57OnHlpMKDRc5+iJ/eQ4tQ
zwknQi/lWKeK5PflZO707EmQTwnF6YaIrNeHYe9eodlCPhAMuYlcRnB3VAuiCsMx
kkadIYl6jPv3hMFFzzsmmgd5G7fycPlKFouIgvOsjOGM/T/BBntKinSJWiUJCxYz
fzmEyjO3QX+q9wwUGoa5isTInh4H34BnbnYI82tcCEcfB/eKvYFDBYHEyMCK4rqC
X84bC2WTrXTwhVAmLjGbYSsFwthqcCt7+0xCBoDNGZ0AKmBZ+A7Wu4PFFUo9cciF
bQjg95P+FQB1SfunfG2MBew0GOjGjS8dlFb2zYBuamA5oFS6gh43td15xA0fDrfs
sWGfrMZIKJNcKdz7q99j69Ki+QEs7qgnrVTPpcfolmCQk1g9rFB4SeCroqZXHZur
x1IEjMvW8ibdyJbekuhgp6cufjXsjWdWarOJc1O4SSZmPcQoERke3kxA0QD56nUf
bDQGgYBCdkYTIU2IgEuRZUny5/dqBtivRSEdO7WCeSocOcy1k6KY+l0SFacpqJzu
QO157HBnJq4/nEIEVAr8xq8Jh+nrEwvFh+BvuP0jNdm9vX7JVQLJX9ghjkC9TZnc
fOy4uISISdWlu4W3S1OwpDg4gYAU2X0mx5IR6LKFn+pMwXLN/2zDziHjvKhXWEJK
LkwFOmEE2jmBwXpBIV0YyF4pXEhvmQLMKfIMq4fjzIKUaUlxkX/sGh8BBhXkw4A2
iF3dyea+Aiyyu2o4/D3os/DBH+H9oeMGXsNfkaC4PCnIay+KkVefxeDlTOJCRbPJ
p40dqjTc1JlDtffMl1ZwAfnPdHXJJ7SNhx4BE47wQ48R8Bq/50hdMh6KbxDN5M4C
7Z6rKQb5SVcD9Ybt+9lBJZr4vYa4Zfe8MUDqzPjYFQCrh28J/b7SE1i1MNl1yx3J
Z/DjO0opfWgBZQbtE6Qz3uezRe2M/ChbW8OUefpawRXxwEhz0RiRM0X2JS+x6MvL
fYDpuxneEcT2TH3YnjlProRuPUBSo0uHvnJR0Zb4CgVoPb0DPkrsyipNLQi1swKN
4OKhA82EWfQw+VTOi+C2k7A76aWKgeIa5LMMQKHoOjjJhZSqoiz403ptuoSOKOk+
2OEaUIw5TtYyCIsNGsMSTfoglH7dW+ZHE15btsnMt1NMKk9coAO+qtxBj4hFgj3J
Nw6qfe8kBaO8ZI75VHQ4JZi8fET1WZmb44BUp6+JDX3fTUo0YMloR97EtAfsY8mk
ZNAcSdyZ96Oh8n4tzCiWEvCWXeygeEcDayeL4YizDy3ia7bz/nwWT2xasuGa0dqA
K95qMxGkWRTMbny+seQSv24SPNfCnw8OTroBO46594ThxG9ggNbn9EFw82l8XD3H
+6qIDS2jrKmx+q1/YcSwQdYgMWi37FCYk7anuI/qSq1l/BGicdAySd0CKTPUH1Cb
uIRwgFGDn26Bqa6uM2rKCQE4yzuLlDNqF47UtpZU1mYagpTmV0XaHfhlnn3YDqnh
Doay90YPR+UwJI9dt3U2ttH8zaFeX+FUVmZVKtB9steu/zgcnyYh5X5PTt5G/x6S
3vp5euYw10bZTGdZb3+FCKmcIz6iapb84FvsnVxaPmlDAeyvTNTsf4rijeprtV5W
+lkyWPKSpEW0syrkcYn81nMvd4OBjjfJqFkxILMaItmn60tkaKW7MgEnlgv/wEmT
GJbgdw4+ORI5h6yDT2DD8kuo1/cfKoOuc/dzdUu2Jamm4e3Sj7YWmA45MmJr6Nmm
6D3Wp3X7j6hHHGkcK3AP4wjNjwSWF+LRA+2MhVre9CYUoHr88XjyL6olxkSw/dN+
A+sruBpJLDTo7sthFRkOPsSNZTUIkH666TZ9W/JCl1wZHewDieoqga9XtgF74I7j
33YcLUfRbj9kKXzWDsibtMRWaDlgdtcXlUTWnSMa9fjj3MnOgAMU9BU0yNVP+d7R
GTKcrmdRubhSb4P/gHsf8eGg385BxvW4MxgKYRogL4XzcELu+L82ZnoROMTgUe7N
ASEozdaBuW73xzvDZIhMDraTV8gv0pssICxuo1X3AME22d1ddw/k7quL/3yyJtFg
nFbRswy30XrTP5ILelrfWN+yjaSfsriOhH7qT8E0HPZpGoZv3A/unZpaUMcxM1Rh
kXKlRG6BG1coDPhgQmzoFVT3Yu0e9bQ94Ls02W5FjKBEfGnBk/xRoS7VhvnDosaw
sx6nmwnTWcLyWRsW/HyIWL9HK8M049gvcG/R1wfW0ZQ4eBvJk0TM+xqF3V9YP4zm
Ez47FM6XLMYPiRd/f24mUBEgC/vQRv6G2Kvfa5N2ek/o2nvivW17F7JYW7RIl3G8
9MHUpI6x2YpHe60+7ikqyqJED56W1zK2fudCbUh69EsiMKDhmodNwA8GKzFnLZhg
Ez4nSbHyQx4N2ip1EtvV1DTzThgbY05DJySmNi+v2mcjkRV1O655Ddviiub1/eLc
PzeBGz+8ZrhMjDzgU4qUquv7KthIXdNxwQcCfeZCzKe+MAk4mACA2mRcs88vgYLg
O3oVJHP3AJLtmc/O/RBhxibtNjp1ullEnZ3V6eGC7PyTw66+3v0vA2wtP0RfxvfP
mk4eXXMQhk1SM4sYjkr9ymTmWwcrGozKaDt/Cku4wme883XBMesJiRCa8KOo+A7n
DMKp9hJseG9bfOAXtKDxooJyLoeLceppa52Kwb7bfJckjVRCe37EZMGJ95ahdohu
S86mW2gg2K9l8ZbTz/H32K+yij/5Q7A+1nR3DTkwDY8VMENM/q3ot+DY0XZkRey1
Ynlk9P2qtn9z8YTA0CtJEdttf1+2VW63C4K7PdqxG3ZGWahTYV8txUGgl4AR2yPc
qug2/ipEXeGFIjBVdyPTIYTK2a4nAQnszvZF/bLxZdARIh7DsvlXE9jwDZSdkwxd
R6wv1osptdvL8Ux2hqpE9qymd5Fm+891J/SyDVyCTEbVZddQvKw819CPjj2IuUGm
MFh6N0lEqMqQSqNonk+VvPFgRdFbEVy11xOvbzU7ZyUcBliU6SWp9RAXoOFcdFZo
OFjfgTEElQ/WNmyOoCoifo0UPQXL3wEcywIrGcq8PBC3bYTwFk+disMMRte5Hfpf
bWyMVOqL6b00wiI6R0lMMpGIaTc9GQX+Sbkn3KmgsohV4ATmWv939LhHi15a/yHv
u4ritTI+F6hJNLdCV+FFMUduhHQdX1tUj1ZoZPB/ZvoQ25agLB9FCsAqMRIxvCNE
LoeMlAXF/sE11ihYWtYUv9nNOMjDPOI8um0Shs/UepXLcyZrB16quEIy1x/RqDx0
8sUq2FTieMka1UOSWbGr4LSJVgL9uwDHFMWzyn3/w09RS3/S9kSSX0GOk4OUi2cK
YLsyCgZbxED4tqVYEWHPYpdQtRFPWBIf+gZ+tB+tFsjN5lZlvmaqx9RmzrCITE7E
uZrSNSMryOs3ivYL5cGdb489Rlv0CObA2YdHBPN6F0Frylqm38LMgQaLWXOwtZpl
XpEjE7TrRPCpFpgVWq5G1Uxe8w9/ruSYO/zelniD7Ir9CtYS9Ole4gcv3JVJGn+z
Okxg7baTunEsG/jLtgbx5kn6FH8TC+TpN77n7AOT1GkdG5pIcp+GhMqPk4qWoi27
HFppGliTxv+Fu5396ZUNou4smdXW3I0df2Uw3nBLxFyU90ozLRI6H2aW9pFTOimu
8Yf+cRxYfVEpx6MyFkKW0H14krvcCt08jo+4JPG4wwGV+AXR3wswRrIC3g9NKWOU
NJGswwZiTEG3grRj8W/Zh7cDnDTb4FGApQHdxnvMVolC53Rxp8loKZSMgeAN3brC
BZ0SI3/21kf/WucN7L/JqecgRBRy98dqdDx+TD0GxoFPopzDzaixTxGQ0DUmcJ8M
/peNGJxG3IMfysHynCNxaXMUl9vr3VkwWiNUWNfzHASlWPpkiIduFMiDklMiOq/W
bMM0im6/GtQZt6C7bsXHVo5FTORywtK+1vBOS/WwYnAkhPM63eKT8KQtQxTkpaUC
EWGlblkqQZIQ43VJ33RtL5MsvD8YyTGDwdJ0lK12Uoi1CUEsjGHUof9h/c6R8Toc
LGiSQ6mF8+/WVC5lMpFH+tmYjVgbP32mn7U8Hvy/16KLN+xT2jxnhAeTDA0ySxP2
deWSZfu5MfpqYlVpprG3QPN5yvmHsxFBZuEkiS4UP5oT7CdgTbKV7RcGKeutzghC
rgGQWG/MY7qz+K5MPD/rN0xbRjKtvMo/esrd8kY5e20tufNl+XE/dAnr6On20q+/
G9T5FuHeH8NHSIXSj3HEPCgbunC8pncxZHHB3hEVGCqOFn6reyX2Z09H6uGJ7QTu
dSIvTRCdKjWyBN0a2mKhPHqglTaPs4epqsjMsSfPwtA7WmodiKuf1GnVaJfIPTj1
tiXlt/9z7Jm/sillWkb8BfhQtSc0EMuxuAK3USbSkkOAg6i9STrSBbfKvEXSVvzE
ySwQ/i1EtAVVAaFu0lUTchcyHHdbH4g32olh+7/nmmtD5GMnfDC3ihZXt5NniWYP
WLNFbH9vEv5HupUdscy1Ks2cqIe+kASCXG3ZaClNzGR7aR5BD+NXxGQX7hYr3Mm8
qqwHciF7lNVXLTaxBmoZPVFdyPSzaKkZ/iKuD3voCg0m2bfoXotp7Ou+0JJghywZ
hFCNHfd1HGfpRpkmXQT3k/A10GzV6ZJS4eYXEtaKTVBQcr9ME0lQEDooX//cF7ob
axEDe1hZ1eBuMrJwShFOBmz754Go3zjAOLfLTAl2ZJ6fSQHbeWk8BLXy2wi4EFSG
hXtARfgL1WjUqPB+vwsQj457h6tN8d0Xbg7ilZDJC+sv5Ce6h5qomgvaPPqZtQBM
vr6RpxLufewTgrlLqnMNANeJthbkkEdkYsE0oFg9Ki2qAsSN6rFJt63R95WftChT
UVFvQq7TWqKwlFR5ZhL0Zzi/xac918DlY7P+iUCHbFzbQQG5OC4oToGQtzAlsPpJ
1B9vS9ulpmATTOQypkzC/EsfDrarXGQPIlcytan/kPjNvabqTHUCKq3K2MrrWZTN
FLs3LUON7kHp813Okfq4oiEu0xEwO7M/1E1ptR5COJvR23PBUM89wlyx0obBsZQ7
OXCD7Dh31wG0sS2fFvlEfRFfxmgpkUS848mCJeM90PvmExWzMraXByxRfvGLVX9m
gC8FiHs58Zo/BdFfVRy+HWDB91N03fVqtPEu5KMGX7Ve9x2MUNlT0oUUC5aSVdKt
EHnfsW6+9O7qNtC1qwLimlNQam2MtciQLPTqi1Nn5u7pmlZR18xDmEWF6ByIi4Q0
qO9zuaNE9yEUkQxIP6Ye4Odb9sQxFd2gKH39keccwyqvui8fWoXrY4mhmLBCbCg2
cxofqt4DLsW7/PbZdZ1cWtek/8mNgzgzPtQ2w9/EpTyWQoq7Qc8gN0yR+uNKZ31/
ppyIrKUh6FOEttipGNkqgjtqh+TIbKkR+lC6GmkAGxLOcUJCUEyEYjav4CY0pXPj
E8nCh60XN8CrlIVXPpav1MHRIr6z1IeDIMzU0m9jab8fjNmfx5uyaKF/oblq+CVL
4xlzt27O/HBXc3T1ZzPiSAxuyJSaZYhXgXKwzO/paiEHSuoaMS+YYK7KDZwxQ4zL
3s1CtLdIgFGcThtmYfU0dcFYv4bliFCNnnkJhmR2WyG1TmxgM7sto+4SZCbq7Yag
/VlSfdMXCBAtKQ0Vrh5cspGZBnkFnz0kQF+c6gRJTDjeNZsYYXqmk+3W9oOsT3cu
1TOMnKc8lZG49zXy1tdiLk5hSPAmCtC9xi4iVMy6pG3b+34BDaiWOknq3GFYhMYA
u2qDnMslGbS/puh9kel03uiw96JKVQ7ByNOKv8t+h9FKvlud3twFt+EciizvYrjj
HPrnV/R33nEQ6T6Vle7/LFuGF9kkKpiIsN2ELna2oHSHWDFm+PPZyiJDebJ/biat
x/64Tc8mmhWSPgsJ0eqoMTXtyp5tuu6H4ls4klq1jD/UoLd7mj8mW2L8sCeoKrYD
c3mrWFB+mQlA5+kMSMQ8GIg7I/Dic/EWJiWG9LtqtzpyzfuOZZbljKPfOjr/v3n+
rUdD+Vwm/WmyNMSilLuN1ki5kfh3GphC9MaDQmMsjnqwpLafodfA53U+HYXmj+XX
1wNe7fwQqG+pi6HMSWHqkatIE+v7E4V0mBiQ96oRBAF3Enu+gOTIZo/iZ5IGBOKq
YTk+KXQ+WcRGVrBG7QeP4WWMWW41+WK6m/T+yQSwgYDrfhZHAZUMgIdMYcNrwkFs
lWZA0HY1fA6xvfMRv1pod/l2Cu3wQxxwcBuY/rGkx/KQvgnPLBjbwQSII7I21UUB
i131HpMmM8BDktWDffx/k1Jsr6eX8nOzHXMhntsE5qDEK/EtrVxVyCEdjQ/LUdY/
ALerJJPXxAj5QdTT7zVoFQu3R4CyvYCLXZrpu9IW2NaJMvETpOsc6pgJjAUYMbda
XkVrGy0/N6E9Xg+8G8hTsd5/PH9P3NNpwK1DKyeWR+eyN2Wi66mhSOqxvDYoTDXY
k0WrggtOvx3EFlG2HKeKsen5FQlsNt5HOgMP1mA0yCQ2e2nTEW9H0d/EuVdN3uCL
f5s26YD8O3bKn7RVXjM7bkxXCmSeTol3mbUZKb5JU3HmrnkyQrBT/XbURKNm18P8
EcYHD730Gwe+tirMBHDuTuGg56fDwISbBFuzmcg0zZS3gXPyE9dJE+AmEs0bTgwe
bCRQ3ckGfvn6CaHqonc9VlW/N+a2ODI+Rrww8iCMwViLRibFGl3aI93D+ah0322B
8jzTF81fvgYizx0Uvef07QySlN9N9fzc04x1tXDPiYN//55Jy5pNieOzOLbIhniR
6HGy+yXIUE0NFtCZppvSHpDcJayE6Sku8K2jvrOUfp39AdcZLSxmHGCb0spG5XoC
G7SB9BM5y+SMdutL8bAQONTPgEq7AwnhYNjPX/V5pNw4xJQl51OpzqAacIPSk2Ce
soEoNrLoispjEnAHEHq4kKptSGDiBQXM09WOMZKhyjpcNO5RdjD/FwTU7Y0lB6gU
cZ9NDmZzr/US33B2TSrNrhamy3WEAw2BlJyiwfm1HcjEUa2wMY/NX+O3I2/nf6BN
il+/p8CAjC1aQOTb0mMfFLhCe3hm6M6AXzAH5rfBPpDodt3dyylZaZbRpSoejyVU
HB6urYYe8FulvfFWp9oNz+pXtQxiVmH61zCG3yZSziitiWV9yryVeYrNKn4LAC+/
3GPDGgYmIRmrR4GUzngN4nHv0fbrUU+iwnMupdCuJwmxKLe7/r/qdySl5ZtO2D28
MQ+idJVnBNCwk4Zt+JThxk8QDoioxQA/Ymlg/+z4v5S//YyM1bXHh1PrGI3I6CRd
RHpk2vNb41YKrrwxdSxH7p+iqAqj9QVULwDKEMYWK/vWAnEYj9Ohihutkobre5BA
vxM4rgukaLx9DEml9WOX2kKq53tM/RMxf6zVJIjnTV28ftBKdnF2eoBNegM/mr+V
aBXPpIvnwRIhYp5LDrY3k0dKTVhXgwKFaIgoceGalH6sLhLOC5QnKS57syzWpGGI
268XuBx/xhdaljRO+8rK1VPP97KX3zFKbuRjwaakuAXhI8cn+uIZ9OfnKmFtE/Ik
4OPgCqImW6bA1IeP/9MBjipyjVMxNfSJXRoTYp66bBPrSp49wTJ30ayOl3gIh7z8
hT2ikdFO4gjW8wVXB+nUQdxRGjl/DtOrea7h3zWtBit2I4AozyNRC0zpadfK2RWA
g4N9wOQz/FUz91IX+elxM8Cv+F25RueKMA+i/EOd2C6xaztZsdjuIAwR+5RcX1Ii
q3wi+Ra7ssxkqgS9UDbX1psAGG4ZJZlztK6io0xRA1JF+TicDTZgwi+LOpsPn1Ug
dMy9/+b1GWDYzf7XIKQkhd96ipdYdmnAtl+Nne+t1uU+2tCugkyYPsMCN6nRt4I0
k+PVzddapBrrQFJ6HmoyI/sUHuBDUEU+JgLs6VrwmXI8YfgHCchK+2LT69vpdVuL
3ACPhS5rcBWDBt7+qBHWQClAewrcPJlZmT74fUourGi+EFJIeL1N2G//D1GA+ASa
IXEXJZVcyss5giEkHE4a6Xw6K83E/7gloyWH/Q7lgC0GgUKGfSlDqptY+b/rqJKu
sd5yZMWD1YWdvAfHje1P1ZV4pB2Obrm7pDbNRwDvf/W8raqH4bTNZEkmEFihw/fO
yOLyUrUA9ALQ7tMgSm2IwCVS/j+YmiUpMzDiLD0WPJ696P1BkX0WNnyB4qMiVb2w
/Cw6cGhSwRZ6ifs06caaba7+OXoJo9a+8N70P8Bk9z6ooacOfBo9l6Vi275N2CTJ
Z9jQK7eH089FyvdATi6xuXemHzqieQRjF0ySqx5DbjJz/oC/RpgI9K+tEO/HgbZp
SPm8294SwdUXpSi5ab62tYwLL9wmtcHUNT6vpCfh36M9DlBMPfuUFMaZlAA4zr9j
IKQuknsU8Vd1yOC7CWaIxTONDio3+3eEWFbkapQ/bkiWxhzkZ3tCpGYqpdY3G4ij
U3wdFff7bxvKYUYsC5XkPaLZFO/J1vP/UO0WythZBAaWRFbjoDZERaPPvMldP5wO
fMIL0HP0uzdOfKf4riMZ7leRGV0OGVmFcZqBXfiziYS7ezwysrPwRiJgvmVyS1rG
O66wpmZNhtQq+8kG22+NskV1wiSIQ7jC0+wMhQBVanBK7tQFtF5j8N/MbBtsURBx
uYtKk4pFP/VlVXZxeuzAUvXuKq7SlPO1B63tRri6WplYlxU3A8bkWextlOJfZ906
9+YgkK7AzopPtrbwhxFdEb0FFb20J7t1o8JG7vtMvenP9TQcYq+VkBdPRmy6cJnR
T2OTEniMfhtQwJzvUYlH1LueSAEOMASmqoBuNUHH9KyLuD1OX7ZQiJqdRSYPNs5l
wjD9oljyJQl2cAN65AXIOcek+Y41lGe2WGLdpMzVccefIDYmon6Z8IKP/mVg2k+k
yOIXGW7ocY8LRTK2PU8CjRGTG5xZdCnVOlNEtom8fG/WlpV+YTrHT5bn5jLSAwDA
rWHxv8Q6XuXc7zaSJy4UDF7FNPSdVX6kDKIpTC6OdmvqO+aSRmkK2P1fyDJpD/kb
mVyW2Y5BP72YbDStgvaPdVOFFGMHnl1TGU2GG7U2LwRH6ohG3mR0KLOoMZ4oQ/Pw
ut8ucnuOZtTj+8qTHBi+ww74fqMOVdv4Sybrgm1w/ZqjP9qy9PqllSeINAjdZs0x
ith84yvRu5vr09wNRUq106FX1+/XZNOwRrwzppaTWk1bVjInTS0uruz6Ni+sVorO
Zj18EeN6gtNMW90KN7Soj8qBUExSVR/OqewplYMDkOUOmS6JfNdazJVGYQxxmYNg
VTr3OPYnPETK+XJVGtF/CfrOR/8F0kTNCVoOkbfGEPRkg5M3rFiGajwIZBvNaumm
6TvLYIQ1PjyumnpYfJ4TgShwngieExDobK/qvC2zlkt+5g+k25F7CjDcPHj4GGxk
MMDvIEp8ezFKfsTbyXxnOLDy4gMKH3blhbGP1UgOzyVxguPKnxQwbSLDTlla6aCl
A6I5S6Xfb8hSgAp2xds3Zk9fzBTl3alV4yOCbBivRoD+ODUqjhSIHyxRfMQEFItw
O55BGt+42wP1ZjbVzmx5PvfOPTESKM3YKoVo+Eif3MAAlOnkgqbMMz/N+FC4UEhC
yF50BEMukB2muKADNoVl4EBqw7mcoecQOYxnOJQzH5MKaC15vMj4Zs1T0ScozyUF
p10T0C2/0wHHWIfOm1IoBTIh6Lx821C207bcZN2FafYVo7VECa1fUIUxwMW1nzXA
LynlRdh7vI6Qir6WHvd4NYIy9yZXxJO1sOVgnQBLqm6o6vWX0FZevQMoy4uKSDUT
nw8VMHKesTOmmcwe48UElN/zeLT27lxdx4+o+qC4fOCWkbgM72jKJNvU95LyOqPF
by7nPk7PO3x4DruT5Bp2DjL1arIrGr6ZVZJQ5KLLZNSGuKR2HM+dyyC+Ew+uNT8m
jcrBUSDSpzfFI6jNSsvXWluaD5nFx0RmOMtOi63AZ5kLv72fw4gTtYLbrv5djnIz
qw78ZUKbpVxYQm8WYkb1a2+RIsi4AR6vKhcngxleYGO8i+dT174Z3+ldJY6wrN8I
emyuUykH77KrY/cZYqnlY1o8C7e0wECybrnRJGilxCmsPxao12SRzHOgDNE+NPTZ
ZL2SY8CwWTFNMKK776VLxUWVX1tkyN3zYmvSxaBBv2u/jFN7MkyEfvahmFw0QJqg
MonuEXMgOxOJpwrWCdFG2W+8B8Jl6EKMCxQvsMZ68DS3xj6WPPMavRK973/21i50
dH4x9oIJCFEKQcGKn6rypU8FkaEQ94Ki3aqpRY9sosui9cWxolAL8xTESfXp44EB
sWEFSccMiQFX6izlpV0tSNXIHnlFcsggcon37CourHMLGGEMHjav597RwldMNSJh
MxjnbiLfpmyLiaw2qDcAHyN5rWq/MBiS9mlX3odl4fN7YvDjUYmTXPudl/5Yyxne
4Cg7fxX/NYbvDhCcsXk/uFy3Cuk5tpqrGtEmoxR9GkNzckhiWVWhzKBoKdSSMEQI
dkNTpPX5aiskW6FZV3QOUrZuOlywjzewdWA+uoOc3UwhbEmrLcakwVO2cW16eRGP
Z6L+krdqGkteQdf3v3r98bb+6etR3b60ySHAlDd8udSzGhCw+GRBAW/bNV2Jc9v+
xlsKTjUh9HyCoG7ZEUS41U/7dgc3dfAZr++/8Yb8NomGMqzyYrhXLZfk3WXAqqG3
stt+Ng4VJgXcbhyuHNSjkNNFxci2BzVA15Jo8vVqBf5vX7z15FNOSCw94ryiYakn
XJVJ7q3E3/kPbMCQsnTD66eGSvUkSFVQeLU3hEPGOIQQ9Acffatzi4B1q4EUQY7J
0Ue9goClU5AfYvC1oQrmlYkutRlVfxVXzmZ0k1Nba9zCKQp2zSxY7uJiCgXb0LwA
bmts4tlHnLvcJwbPmu6VP2vJCUT2UH2lt1qxDp8vcaMv+O+5DU1dzZZChhkh0+Td
FvgqgesuU7h7Wyqkcfjbz9taqNJr7ucDFdEjcNINmlyWr5zOfUpWIhPQ2OFKUaL8
E6fCPqkgHJU/MImZZUXmfAiL3u3Wraren8wT9LK4ygGAvjyEs6PrT/mp33UVemfP
ToaFqO8RrtoNyn6mZnI2aeG+gTITF2yXsrXniUgChMQELzdF0y6JsdvB3h/xrNMG
CPkbmsb+YmNsuq2KRoy+gte0sYZoc3vfg+ZiJcrWb2UF7HF6Q49i3SjFDiJ14+y5
uwIx1uvA7K1sScNIzPg/+BnFPB0Tw1GSKKp7svvptngHatYc1YhrNFzix7IYDNtm
dPxaSM8PtEoG6k6r9PX3KpLBHmIGvdQil2tEQzQhpCoQNBDN0m3ihBJMxD6W2n/9
/qI2FJxR3pEVNBW//hkMuNocYF4y8dqzl9Y0O2Kfc8YTphQ8mdYGuzznTAaKSxdZ
dUdopwmQR0vtFRM6D498TYmFtNdbQHTEuBbK7ShYM7bh5/wHjeRQP0Pv+MTYNB4e
iBKPjQ2QKakgLBidfNW4DunFJN4DxJ/dVy4UvllyQjfiHJPDJBPojaOtT48LjH3f
qgSOsJnDI5niQXqbCOr/8P56Crcc8vNlffKTe+qo3sOHaho4X4YOzZQPr94Dmbte
iJIj1GZXKgqZ70k9OkNvejElAr2jbbOmDZ9A6USs7ZDnO0mfITobjjGUi07tUCO8
Ik6AZbPSjNeajvDi4JmcBBWIMLOdcKOYEq4zFlyMn5uMVSoawKgkQHzRqqKAsLQD
szvz2GVksUBZNmOPlUB8tnJYGBgTCvvI4c+dw1KoqsX3eKDtN1BF5nUEjGgFakV7
+K+QFKPY+6nJ34Y517TdX6f/1xHtllMBzJVu7TRLefw8iht+ZT/rDIKiO4nXZwY7
DQrkMuTsOjzO0d7hHgOfnPFI7+p9RM24WA70efR53kTrCm6IRvVw0ULguCMKQlEF
bC6dJoD0NBZeibe+zmQ8YnBrFF0KtM/Kig8cvqiCiaFxZYL4B7qfmr3XivqLyY+m
W8gFqSxcp2r4b3Ma+acTJNHn2CnN87F7W7xjdDY+HZeyYN/e+JQM8soz0q8cIpOH
+KKcG0K4VNDln15Th5X/HgVusHDDefrNUc04UFyMF4nb5yY3LV7DrRak9MnsTBAc
sFFaAm5OlilaeZkJa5t2Yy+Z6DsdjpmMTzOsVZdIcK/HdKVWMbbytJTWaxNyQqSM
t6fqc0IEtfoiePGwLLQnA7kU7w7iHE6QCYRgkCupzdJKdcf7F740ygPrVefhvRER
Kb+fqCKUDrcrNhQAdynWuvX0PfFUQnIfYrBIUbXoMiYvQXC+J9zqv1OzGuwNLcha
GooIadK+3+/Du8ZAJ0Mhwvf04tkLGup1uH1YCIVkMICMbNkdvEwBq7w1X2LxXNdv
WPeANUY6ybmF6byKXd7pSaz8D0bcMVbY43KlDUKWqGJwLfEW/Ub731nL0cs2mAWl
ZRiSbzwNH54MqKMzB/LsSgb+zxY6d79NqLcGRkx0ZDinjJ4+TSJKADYrUhKN9293
ZRQSc48RwG0+9c9fOnusyTOv7G+P5miRT/UjnOY3e/W6PeJUmfzO184fQLlM2xg7
kTZ+O6BpElkjGW89E4ok4uBYVsSyYl8WkdpOUuPYk0i26s3UiR3p1BJhvQBftrVn
81RV+ReTJ6relwF7/32+saDD+cd1/+tjspXTW19QHzBDfMWtPS+o+3Ts+53t9rF3
5mmQm+w9+5xofKtvCDnodtf25O1qUDsjqS+dPrwDiwZ/ka6+4BkFtSKB2MPql5V0
Ng8fwM7PvxxMOazDCyg/Ae/jlH+O8kaxKGb5ADgxMHuzj2ePoR2I8S76ji0gSlC3
hZy+ANEwJ71VctLNeLNkBd1UJrZyGWuVXmfewDjRppa058OvwpkW50AlP4rPOB2Z
E5B0Z3S8tjZqEa87B5NeH7Ipar/2CGHIrlN9rCwLuOSPLx63SUBagpzwBKgs2NIf
gkKJzkxCCYlGyhOyr2BoDMoOc/rYFYgAunC0bbSjwelMtTEQKItgeOne7zLQO/Ae
YqQ2JwGFdFAjq9XyFtSxvRvUUE9L41CaaFDUL6kMi8+s4w5qNLRYw7W7h/uN8A2B
4iJyamkff6XQ5ozFG9DE0jPoYRohTfPGjjOEzlX6fijbvefhqeQPsLKvF1pu48Kp
VH4cZBdtWh1DojDHFTYSuriTig9B92h0i0eQlapktY6H0lyOhjpyepLGDhCSX/1J
gT47hiFW3szjTwZhpA5fKySeTG6t/3hN1EBA48AT8d5Sd/UoZ+q+EQadL4Uklzum
Ogd6rKjinDaxzMdE2l5mG2B0Z8krlzVB9fR1IMqS5HaveXDZLzq7ZbBu3s+06iLs
xh/rMGCzrkNAgrrqOt3f3vWd9eTA6sV0HlThZeYeKG5M9qyVc/C+Xneo6lfJa3yt
Z9QEAa7/+87JfbuoXbJM6ggH9Wl4BdvqwDgADccxxCRgo1x9QZLmRQIBsYDS2OYb
9weWFxhF5TBCwy+mWeVmxiqX4wLjGwKWG8D+9vPbheQ+RJZYNNtm+l89f/sW4pNI
nN6cNaEAbSTXuIvjK1zhge8whQwCRj7uFPuo74P8wJRRmdGxO2djoSObp6VmP0xF
KNK5XJZS6psm3gyrL/cRwE9wku7bc24Q++MYrXcwPrkorVhSPG0TLfvhyERq8dSK
NMUAU2pTov0L/gjGM+E39h4/gczhcU2Ka83K01a6d7x0iNVI+pv6I7StuXh+v8SD
QxY2OmlAFUnfORiSf4qucV+lE7ego8qFFnWCGuefGq9p5wjiPv8k81+F48xcZgp1
HSujpKWNaoA0+Vdxkxsx4McNxGrTMiUZD1W7HuGfaDXVqNEWUoLx9L1i4l4PeoV3
ZbZvKy+3xUF0/zyI1Xj48MBu1IRnsWOr4LEANvdBB4V4tP/U6a9VWGte1TBdVcR/
HEdU/ZtFTl17mSo5kmDZQfOsLHhAQeIcqmx3sDiFHQ25KbgoU2tmcpZC6DubE9+R
vIGx4VgRc9WiORHVQPHiTOiypoIwnHrmgFtm4BfZtMHpWMd/Z6uPpOgGj16IHjLY
aEzSe9WzG+mLgwr97mpAjHrP9Rq+thchraDfBSAI0ixbF2G0+uiYwNjaNkjtCxgy
R+ELteHx7NwlAhkM/BQeTUtxFBXiinTmT/J1tfh/d7m/1995p3u/kvAnPLsRSQqZ
qC5lbKnHPristDP1hHm5GZAmYrIPeaFsYyqgIMw9BtTtQQSI72QKz1XPCmh4R86e
uAanbb07HPhfcaSAMNaMa2Kj/UhbBsjoJRgfxFWtuznqmExIFSLITG+Jp5mdJfX0
aTuRMAERRSxy7CD+X1SywzN83W4IXI2kNW8kda8/Jdr8Gb9Z+yL/SpkO5x82UDJy
mJH0LfqjuavzEj2bs9ahSQ55Rx53USxrpuI5pdcjsm3iqD3yV9D61iY7UGnfI1U7
L0oQiM90M3vkM/vrhGVTi4/tbsOICgKefR7MSUTG+H47tjv2VRVHWU2PmZ2D9TOW
lZsZBGg/IPiX7s4O/e3+qRHziWwDBwGrO/SEsazghr39CSt2Ncb9SXTsJqZvDKYC
7ksSJIr9AX7VJh0y+bUgXuj5guooJthMwGFZc00SfholaVXnPMbvq6ms8f8cd6Db
Dgx6RMIV40NQuRDyHv73wQ1nXBIveIt2YNiLGaShzbBOv1gi/3mPBsQ6Bf1+sO4H
mHkRwwVIGwlXLdH//4xmgbXERiYCPKcdr9eXPyOhwp1jnBGghRsvhBIfIz0bOSmp
T+HO4mHbVUqRMeHMENP89nkCTCVMe9qqhq58ysGLxfwmjeRGk5MOgsYTRB2Uv6Cx
+5D9KF7NqxNn9lbgVCLd9fYaMP05xVwIdB75QMQZPoAkvO7quaCKm7Mbohk288PM
MhpRZ1TeuP6pxyzWBgtwti0UG2qJypRFa5CWPFbKNz8tXdgQIrBeKDHFuy3oBslL
S6xVveTu8B32T+0gcVHMlJs0G2PfSXsRlUZ4qmjhXakHr/cIvv3wdIDCa1wH0gYu
q5PwR65npSDov9/oNLIP033a0O6Yft+Jws37JFmX0XvAN8C/ZBMCYd6KNThzeSUd
2/MJnqWaQWWnD41l7dBNQd2tBjmczOQILln4KxrmQ5uS2l61UoKybv5IuSIdYd0S
lcbxFqVU4muNVlHdY955SBRw0hsSA4uOknrz/6IcgmTVq1GQ7RguuYBV2VRsECbN
Ixxy0Jnx6lm3GFYTgGiedSEF5fwREj43ptkjuzmh+Xi3c6WHVQjSJjz0IgSM2qnf
DvVriRWPzWjDJPFNG30Zo8k9i3t+VDNWUFZm76qOrAsw1iRpXAkCnCG/03+P/GSy
/RSNpj3RaxuEHAbnvWWKScCkevkHbTX2nfljKktghbrOJKYGBHmyfajW5nXOk7nr
YtQ7sdqYXIRV/mqd2fGM1gbrQi7RBpaUqWWI7W0MP45sVvcRjqHMhIN7K6An2X3j
AMC39QS7bqQCfdpn/vmCUSjbrc/yzkne3bszyYOPIYxl5qgAdPSPyv4bSdR7RNXI
LYko9dAC3WQJP4Qp8NfWu+fG96i82l0zeGBwo71lVrNNM21C5LCwJ+WZPIYOakmY
ZDJECerAHxVnXTfnCXJmEEqtb0zS0bAojl2e/1lClXvw484e/1er698J/yOzQ99r
nop2bnW5RnF5yq4CBwz/rk2ZiX/iQwtwOOF1tFgjsMs6AQU7YCJqqUTbe3PMsaHR
zDDsAmlMe6YN4y4TGnUMak1QkJHo85IE/ZKSDIiobPsJSs2/fbOuFaAVZYXKTK16
AY9+vw1+eUI0H16IFy4r8P45NnmtvI0qnVp+h0Xyeo3h74qsWRIb1g+cq85BcixY
KjefhO6tdJyeoeGcHnYqs1m1KQgdt7XEVliDx07US5/lt4ZsYsNFmBsEO4D/paIE
58exIxnDoZFfCz3ht84ei19oGkHtGlljFUPHlC5ymOJhDgeyZ95kJYNK0iZemeL3
zRC9COuhbpRvCpOwHx1pLYo3KGOJSl4d2xbS9F0SAm9kN0eBWsYP3Rm2RLMmpgx5
ou4yR8BT/XN04greacQU2KoUkSV+lqKWjaGwEJ41SmyWFBnhZUy54wkiZkWcWQJR
pB5yvpog8RgD9UJ4UPLGDZf/knkFA8Vmp2KIbyz22/27EVJsjahJeSYZ6nZnUfl0
tLCzP37InaHTKWB8cOoEXJaIMARgDrlSGLID7g6mMMf9DY4IJyN3ScBESPjnRbYm
bvihcIHWkLGMX/z4Fvia+IXh1/UfSWiHVYeEw9ipBxfDIoCzOTGYxWFsgFh9sT4p
gLXQdFzf5eOxVNtvwdD2rcqVwpJ5DsqFTdfF5e87HRF5uLlZ0BddB1hW8vUXcEd+
S+JT/nH/Lds/SqhWa7Cq26AYEejcuEo/lDJ3G9wIaoNIbTa1Js1oPBD4Se9FqYfV
owh80kH0Jxk0TtA1H1rPXkSyIB00c9+DyiOEefk5v4iEHG3g878f0ToEopqSAUAf
oeSYKvfMhjaWMUmtY2l4lLL6y3h+EpaUohv9HL5kq9vigWGabXb0qGOZzxOFT7A4
LVnQk/lFEec66cGCgikW1LKSzn1gG04weUtlv4Yzvh5rg5lfvKsunEDYnGQOIAsz
Tb+HkHdmETa6xRUo7MCjaHPYO1cBIXzHoaQUgQ5esFqmBEfKd6W4v67B/a8aDZ3T
AxpIRiQzrbEQvydmUx3tJM7gsgwVpvvbHsYoWDNdZmxjI5DvkfzotXCxNsTa+YW3
oHtct4Z9s/VyHI6JG35l3LLqxHq6S5Qm0HfidMiy+SHbHEYL+sGPqsAQm0gbqdif
WZitZgWiYNh23lydN8Rdyl9wtKejkC8xHmUlpbNSgAR+06kLqOGQz/yP5cKWLam7
v/sVbvvOH76wmhB4krs5TLQMvM/D0gZOjx1BTNTx96iuGbNkljDUwYit2nrOA+lO
1Yc1AI77MM8TbNKajEJAbKx2jXewQvFYfHK+Pw9IRO1csxzuukzhtKBz61vXRm7o
Yi6U23fMHLk+LZIjGooiMFgkfX3RGe7y7OPi8XBSKKOmZRLe3EhId/U1nLAwfe1K
DYHr+fFr3De6NuA35GBTVc428DY/ergUmmEamzCzlyfZeOlr3KgJir8a0vRSd2y+
26ozL0O2i+ob139MNAR9FUDNas+vYtx5yl8JC/AmDH6qLFu1Yr27DaH2vgqlH/Th
/v9noSdMDoMAC9a9j3qaxU4bo+AeNymOYMLVEBu6OggEw3HDLbP66HWUl/u8UqLu
AYr+y1FKc31dDL6nphEoVPcLak4zkogpnKJHqtEBxIePC1L8FBK8amzrQ52nIN0T
+xsEIePH7xKNdpkSDN4x83WgXrAPvpam5uCydF/sb6t8IXl4SGrvJ0MOAb4TlRvR
mo1MYcnhO7BZgAFnHP8fSFSRaB511LCsJFhQtudxknbObSjf1n4aykO1bF337TQJ
/ojdqfOVPi+PAVjd45Qi77eU1Baupn1WeoYE1tCmQaVFYtmCQwlBHTrsmybN3w0I
bFZU4s1JSyT5I6sER7k8zT4zKq4eOU4gXSlF0YfVKgrVODU40QvdIzlsOeD/HGyt
dIivoLc4SdjBeHh4SQbW+EwDq6ZfPvwDKsnMtSJWAOv7QfCj0SIcCJmEYI0pOFsO
9Sn9RxrPEchrMFW5ClwwZxcqMLOSvcWnz8GlpZzUGVVxgsemaroTL8wU5Rl+bn1M
bZoszmqiPWKywf12/MhlEqFrVT0G/6fXhV+2TW9eglMD/p2XmXzAJgIB4EYravS+
hQ5cj75lk/FBG69rOkVViH9jormjSVwW2ibP1A4vRw5zKaxN/z8ANXa9FNKLUZbx
xdbXHVT8i6Xv9hMwr7hqG+2Ug3EJN1F63WQi/KLgt1X6s/+I/aPS6zrX38l8XiwW
Zx4LOAMbrD8Aj0MDpIdi5OMglNNtMS7DG2cJOeSRIgDEZ71xKMfobLGr2b6gJwRk
sPfi9uvXNZdpLuNZnD/qh+P49cRp/SX3lje5od2bGKWkWfKTCFuq5cM9dg4nIkoo
b6z1/ftr+GcbclFKpkn84gJkgrfAys+yMHDZUDmgzbjqG9h5QX94srfflx0fiPh+
5qjQYRjyseJHuBp16Dl7O4QjFgFSFI4NnKUo4q/PkUbdCmy406/0NWxdeuTjWHSF
dtV+8qi6jXvfOpI0cIXMSY0W/uFw+/k5uPFDoX79T5mqBbidIx6umoFf8CszxdiT
NhcT/Ict3My876iLQKnTAz/OhirwgAQ0uqC387T+q/5GcIRG/Jhfy7rEVpnADetD
7yL2LiGVXs1OG4FrHpa/bT196rXLmEPlOnm0f/NvBgZ4qx/GxElVvVEK87k13FxA
wN57hJocqsI2hNcrn2LG37Qc0lMVN0aKRv5W7j9GMms26LcyAJVRjXoBYb5I1pXi
IoRKEBHAFvX+1ysKH40dvn7z4NAPQCyaYkZkc4DmSVgqkxbmy8QjuYoaGtotgvNp
NZhseGDhG++JHvVM3UmCBaZiqOrr0He8yh5cfj1QHWi+e01As4Iuy2BqN23Msj3g
nZSfMzpjyCprXmFc0f0bpzGoho0xfEZGBNF/7X2/3VeNhvwijtfgL/UklHyXJGEg
zlfWjs3pPVyXb1jeoNA+slxbpP1KGF+4C5htjlJAMF/KM9bfjz5vaRtTDhDnx/cf
fjidrDCQba0VtbexhFpUtFvGI0e4UNP5tVRvKYTF1sFA1ZJxtKcctvLLZKa03+lO
VGVpWjVj7PcPqMr+JQV1RP+z56v7v4TztFk7PDUSTh9XIqFvbdUJFYf9uY7CoyJf
DtB0AURVPfvffVctQ6alzvtnCCWGL/ZcSs5llsgAtaxUfXTqn3tBM/bLUYlPZjBX
+bbnJfpm7UTwnQWshWUJA8UqqcBCMgW9OwuHIGHbDtPxXo6DKYTKJkzCzs/8UN3S
/4SUVRyCMc3f809PTPig9hNMBOuZThBXKLIFqXYM9BAnBRT21HF4h1N1B8KxONy1
EG3Q+fydSgA1kI1DP8hdlz4ECgVomgqw04z5Zw15tesR72XzAFsLJWpKKz8pTfpH
tw3uQqabJt1Kp2ot9zFxqOwNE1/P8HG/0A2YKxhUFE0rftcsJTEhRkxt9msFRYMr
2pRSwRBK422+T9iy+uCawN9uFqrJIgcPgG793eLYgaKylAbgsjPV/frgPCZQbjmt
mYCuyDwNyGi9yG9Y6ElH7fNVjzIR/1do8+QOxlZ0OSoyFfa8HJ5oYZlU+D1yZV0k
RjnhypBr51ezP/Hmb3eGAMlTMd4s+4QlQ2Zl20/xl6Mrk+rE8Q/zmRw34OAN575z
OX+ch85mNlxqPoEUD0yrCMZhTchlVD1kA7z8FXB7DNpqf5hwXWgttBjf2/z56ou7
IPnzdxGoavSzvu9AuD7DnhI+0Dh8Cx6JdKBvKiQaKWPcNsKZPnyQcykNEnYOlP/s
6J0G59dxs1ue0mVVa5p0uE+TeBqQV+Y6BrpwuMwCG701J0arjg7NMZOoGaoXKHmf
DFiZhnorTdoFEksjYsYoL7xyu5INbhayR7bh6W+WxFvYJs3eURghLYhMkQkExPai
TjH1nY303izC+PyUs2ovFPGXJx5Vlwysb6czd4YLUir/hTRs0zoUq4WOTtiUWEgS
LhzIC1+e2mlsgbuKyYtKVwLGe/elbVahf+Pj3Ovk9y4gdx2L3P6c5Xc3F9zLTt+W
p8nBeFQN/h1JsMaPp3gzYXI4nAnWRVxB37LfDYuzUurTmWcpDIs7ePAlHmjzMtrZ
0s8eHcE2a2baMCHo5GXmPoP/qM2SFozc19pSKiohSF+H3LQ4bqOD5QH9t0TdbAyZ
p9wVrSAwbr4vOXH0aOIPalJzV56dsFARED7deiYwoyM6lhdNPzCWjuJBUOgxZ7aQ
sJTbPBgTJqdGmlSMc23H5jreIMu5FR/KF9Oj/InkTFdrzVO9AbPLkk5EmuljOg+l
u9ufRwk1MyJKuRDYh4+ZhINGyoljRIfccakUgTQt25VnSKQJRnKAVUNWPQx+lQrt
Xiv5ReSentufTrw71P7Qk5w0AYPreCmNC+dY/GPUduvSJ7CROxmR+cKVigYK7DZ6
28yDfUyWZ3sYiP0yVb7QnCDG1ieF6588MmqDyzsRRm1VbWSz2g8rp1KpaUu4Prwb
2Ca/vv8GwGW4DvaVD7rZPwvc90nGvvBmXv4tNCq8gbXWzHfZDyBVBMLkO39Q8K3V
KIXwhPgzuYaAwrBixxvJoAneaIlrtQOrmvMV5l//2Gk3VjIH+U+fMpvhGA66BkU0
r2NlrgvBfvfYHzAXbGVJFMlfqPA8KJrV6K/FKwJ5Mt5zHn+Rpi91Q+S1/QMFqDbI
YVk1BmFfURcP6HuO3ImMS90IrgGdoD5WlqV46cK1eYvtq4lBNV8orzr2JEDycr7t
ACt4c3EZ+mzsM9j0W4XOUlHgHMsPg2WE3D4uETD0PJkZ6uPCNwqgCJ2H0HWNilBS
JOnIqPZbOlinvFB0otV55xcNL6vbJ8XGUZKZiBktkKstv6kEHiNafs1FRj/Ssdfk
CYy6Fh35CuDc3Ne2l03s1FqpunPSE3DKrtJs0u0d+ZYHWVkdqchPu84QooyFHwYN
8o1vdhe9jnK0Li/2c8nUQBQnt8haua7X0q9GM2FX2zuKIFX8Pxc7GVyjr8asgnDV
DVrPwdQ/EAGDbqLgs1qWqERdy6j6gytWdsyY+cJYOktGHVPXUEJMFNaaIQczQoRo
H5//tMAc5A3OfDqr/tQDlNzFsVN/cRqQB+k0jh4U8cxFdD3W7acfsagUsGTfo13l
x9uGFZHir6HACFwJxrAUvCrBR7KTGyEKQLaGeBcZpZxJb9qiH4K23n9pbCgs0dXO
req/VGxj2NpT35hlZxsL1XVLRiJazLCzBaXLM+WfBtPfWq8CoKSN41hTFWsbU9ll
BKpq11chz3Wg74+l4L3RornBs2vrjM3Z3Iq6DymIoInAYDR5NlrXz/yV2LlQHBVf
epKVYjKdSemO0RQRLh4Jp0wg6Jp7H8a9UUjLoet2kC9sWWMAdAS/PBkZJ5bmxK1r
HxqM8OxRNOA+b7So1G0brAT+EnXWdqN2rn9DpILrkPruNlG2IUXJ59e2aYDMZV+G
IJWoq8NUmYPOqPqz5RvoCWfag4dranaWMX43MIK/pyL+XrB33MHlUz1RNohA3PRu
anisJnTIFXL3AB9m0KaKpKF/ASQu9Km7h+6uxcRbGsa68EqdgNPqOxxQ2uH+OLfu
Ulv11RR6HBQ0JmkCtnoKUDa6lMtbLE/MnjlNuNbFCvv12wRGeLnlYIjSPsnWK/HN
I5VG+IbdhNJoOK3dsx+tl8p/Qos90GV4EmCDLtUjIAWYmBxYWxpukDSthmJ9bcH+
MvyNWVgvpg8wpOh+wyK4SStXDzxc9Hcj8fmdhdhZjVVkvG4NA6Eh4DZQpF4TrbMm
ztnH+p88uYmCyd4CpblSfw2YT0V7fDZ2NXj/JD+0bv4w8Cf3IDVJtNZ8ZZxCgGQq
Fm2g0bQWWhiivGnlVzZLQHfrufeiDuVZCNajGYWlMPMsUk0zJAJ05BwQbyOZRkCg
Q8EriSD/wAIt2FzzEKFL5UurpmIbPCtylUacIkwChnRcRHkC5QukvpcGFtLPIlfX
fgscbbgWo8TYpJd0CwD2jSBrfktz1sZtdimyNvfyTBUS/2HfHr5p3MBMOGz6vGPP
a2AbijeEmLFHHZe3Msm4HOwoDxG/LvAZJR0AKwHMZYepBPpsZyAYUihkZ3jqip3a
n2D9IgfC7rqHTsQQE49jIxlH6LnZR1WZZHV+7Xjg4Lzd1XwVSfuPPRPytHk18qdI
hQYvufoKuYtXbbusssF2uYQVKiDNcRAZFs4x4ZUvlrC+Pm4Yw9Q3r1l96zWplbI0
dSQ/yuG7pa1cS9kWrhg17GDBHfMsk8pQEHOhs+UsiyP7oP8Dji6LcnDvI0VYc92E
BWFFjHcFScr3kZCY5Rra8v3GAWDP9SSClpQUyKbiXBG1z2TT2GGwm6pPSoRy6Ij1
ob7DqWU8FNIy7u3RXeUv/a+Cn9mJ1v4YgFfKDCCEEhaK2HtEzkHEqnXCV+Ric+qr
bX8+3NWElz/NJXj/ocTZ2Xnt4bgKGEpYxO77nmxePZvCiGibsl+SrVGx2eUsiXX+
Fh2ZZzMHkxu9NKXK6absqyhdfZh7i6ErnVDAvAAlHnP3BnjPedTd+hu/nEOXh9or
J2j62lRxcfIagWyBUUt4mAriD3OJKUxZYzvpN0MlwjaCE3UlahpCbXpqIDHVL+fC
lUaL5/PZcKMzd9IdtPVFL5v5+BoDMVzt+3rD2N3lUQEwkM9suZpihYkVZctYvLIG
c4HhoFCH1t3+5RXhcknxJTnwFiIWI5gvyFNoICNK8DaAW4klmIlpOoyeWxalJrQp
fG5OZvcopPGFOnENRItHUB+5T9Mx+ZI36hh1+WMXozg1kT8D4no5wEVqXScnUnMD
n1sFvQXS4yu6N90V4JXh6mVbgKjgAKSQQDxZHX6nuENCj0W9tERYt/bESprns+mE
lf9wNSxZ2TkfxCpFgviSHCE62ncU4doalUxnBYlsGxvzZu62czQNo3EeL14HwqiE
FG/Xgz6Xm50+XHHTJ9ERDrhQpq0BgjN7bocBIuhfN7JW7qRPQ/Zlm+M4RtmbeHWe
9gokFUArIBV3JJtXmosAZgNPCoC0DgksuJcP/yo5B5Obh3Z2wg1B+4oAXrXcrhdP
AZ34FRg3CyXZVpRuH55LtUoP1b0dwZT50Ykll5JrfQJ0TKaXuixbLeDgjjJ60QlX
W9ZRwfEHLs12efZEE7pwK1c7T7S6nDXzIqm60WhoPLM/qWf+A3zwT1e0Fz9BVSrQ
/o8N1P75uTB4Drv/gIln/BqqZQTwEE/6wH9gyGh/T8MeEQMFR/UyZ357ASsFjGDw
wThQYZsXIbb1CMw/iDwbjoverDF/fngMUfckZ8lON84HlNcfRiCtNxDFew4IXDyv
1LHwMKNsjXN5Lr2i9bsnRaZA08jxlRabEgkbsv/vzG75LOTJBODd3Kx4GjW9Jd/L
SCizBtbZ4T5+4XEHxRCx3HODP3K2kxboMevA/nJ3xe+jqSm14rxV+lxPYMI4JeEY
5fEXu2lGnu7OBbU9Qu60ouuz5Kerek9gzr14cjre7Sqbw11rAEaTLJuCP293FmA1
5Qpn6LnHa5OSo648EVAnFISMD/PAZx7sQl1ngzbJ4uREk1K6l7ercNgx1iq4f5c3
+00ZkJ60TUrXtrx3q76p8q9ydcbZ441qZUzC10q16iNhe8BIno0HObTFNarEBgdm
1spcINSP7O+lhb/E+4CD4T6ZTNOI7aJA8NEgR0xBBmWJk1z+4hUq7JLNqwtoMwFy
Gpbi2FzO307hpRcHaGi+38DiltuGncCTDRonK9NxQ86u2/PrtJlwmtjmqxFFXz3l
aQISrSS3OOMaYnZSwmteG/93bgvN9n3n5mSxm+PlRiv2V5FmHnqEEsiEa0MHrsNk
wXl3y3/k4xT9/Oyh70dEe2+gDFShlKjL0QQvlgyHVU6o4a+J9DNvbNTlrjUMhHPf
DfSGa82kGcvT2vLhU58ZNObv1tsuEiapnMEMK09khkM0x+CN0IQk+Ax6GcJlLxJO
a2VlcsA6B5PsC3XAdiImiGLs4HcQ8OyI1Ngb4Ziei7OlbYWil7qEdfLbjxsHLhPC
O72YaujMOx8ev6E3m52JWbSlgg3lXMwrd0MwO6G6Y75IXW1R2Sof8dKl+t/v+HFi
Dpd2AAZg3a3KiEvB16WNZezzY1TOmLjmrmFvg0tHx6SljSItQOMzSLSoqIMivpfg
pL5TYzJz0vPa3H/0m9yPRu9j3J1NHX93bOdv0WRGCpvrvJORcBK+Al6qpWLkw31N
w8ZmxaDfj5XUzuAb4UDyTqWngNN4k/2UWRH+m3lG6uiOCNfN3KHpBOn+6gc1DZMw
ln5dAp4yjhxqUY6lH3OLI4LzwWIR5nYo1U4O/XxSJeB0JSh1rUbsFR9pSddXwJiy
GiG76f8FLcq58spHMsfjoVXNbpoPFOhXmG5iHxmWEcKEJoKXh+p82uOmXqmSxPTM
fJ1+211vP5jhpvE6XweH32OtsN0x1N5a7rI5Zb1FlfFoIEroKlUiLHfOkMiQYPws
ijAMD6/YNuWeSJu7vm3SSKntQ1OD3XP+MqfJ8TLt90kAtiqDWq60dq6/62+Kj7qP
9TXAg49QrpSTUu/zhUo9hJ3/3Bl4hyRgH7W4O39tpBMoQdxrmsvK42VTTIEU5qMf
aDFqJK72pjsdB7dHGJVlzCn0kziL7OaXvRIeCar+ke5DSdxMLwaTErKgKRbI2mJZ
EhdbssnO8X3qn4sPdB1Z33561a+hvJGGSFTyzpXgi93/5SHnyrRkl1bor4YygXNb
ciUb6cP2gOCJqBv5T+iP0lewS313imowo5go6q44MkUz4QXKK92avhSnvz/NaVaH
TlGaFzM+az1hAWNrSvPpgsiPfMYDnuWKMLcTYwSdfk0bgQaXkbGmGEEmj66H5jCy
BvJxuNz4RbRqpQ9dUyAcOPYHG97p/pgvALQu9fZDenbAGk7B0DtsqJDQFES4mytW
Ph2VkHMlX0AcLHbpzo0rco5wgxBpOpHTrtBEeInYx5m5Iv29WvTt0B2tpd82bpHG
28mQm78KyoyXlpAUfhnOKv1tM0VRZqcnUD9WCxycuzTluPTZaqLd63O1yqcghbQK
9wKYwAHDzT02R2Or+mnQuIPdytEKHYzHCcdmb8jNKiJd+hbyktxAmlBk9+o98roL
8rkz+Hw6S9vJHfE05DF6sepFXVWQSRYbsVtrvkBwX2Czudg7wRQHbVFhzD1wy9qO
7lq4hq0AeFmoyPjRvRZ278hXkQ4uclBUEUJ0iVmyr3feDDMVyfzk4Ql7QwUUWLsy
hHMuLI+snc9g43Hz7IU5nxfH/lJvQWMts0qBjrMydkK+yzJua6gmukI9sCzPWDTP
bvy1XTstcUmi/nwLARC5NjAFeg9+D8drSHqIzT6piet0UiXUX7LVuKFViE/7J3kW
XrV30k9r6c1EXVuf9oBN5sVaXQiGvCd/ia83nrqkxDvDGwWvkKxwgeTsq/EJ/Ja9
K8Utv6WgypFRCEFIOOcUDUajc8fNScT6S5HRRGvAyiLo6dVDoLlgWNjPE/fozIUK
CfN154MeayurrWBx/wsM+JuMBCUMxRi7HVrqjo2UhdE+aoAy7HfGkE2vqWLVcQx7
Ajksr3b+ISfLdR13zYCMrn+IsHxOHZpKrMAiNa5Vod48BGlAUhl3nFUNEugHdISi
Y+R0c2VokGLN0680IK4vTcy5c9g2s6P8ngCR4nG1PYPuQ4UsjRWdEv+ESe6lCclT
e4WrG72iImqxE7BVg66k4UO6miHOi02MALSkCQ53QcHPMH3SllPYXJBSJSm3E+4e
KS1wMAd/SOGHdXuHGy/Qmr8frPP6rmy7kRXY2mymwiAlsBgG3LLhuwcBh7FhZ4hW
3n51t2K4UB8cRSYO2Z2FOfY+qnRLm2dR0WmClkGtHBWZPAs4qdFUnat15EjaeLwG
xVZtO9JZPP2/eEA/4bTzwyKVd7SlfISZp/7ErRp8DboxB9PyZIS8kzNgCU8kSCe+
x8RSn/zDRi7rBr9XMeJK3L9YGY7ClintOP0qbISLdqcUGS9WimUe7cudByvvzNKv
m+oJo0kHKIWs+AMJlym0T2UUZr2vIqVrxuGDZmrYMuSLru+gFJ2r90/UWPbrT9IQ
hLdb+8p9iiICEI9mInh/KBqDdrwTV1+SuDi9fWAErU1cU0sdo6HWj4OEOGSTEg4C
hCfVP4FhkwAXnH001T2hXa/Tu6Lfo3OjL/qNRlJN/hFLMaEThfk5VFmveSy8RxR7
RvqLk952hmP/mTzQFl0JpHw1aLIEwV5pp5TGBbFNUNHD676UObfjCFGoOD0y5MxX
UQpuP7AH2sHq/CEKu75gCGvdubmUJPIEU45i/lMdAx/dhDtQnkFE8tc+MrkEUszT
ep4DRlUdRNo+5D4LQZKCDYQNp8r2FSdPyOkqhJ92SMjUpXtX2mnofiBaBW7OFUct
Yr65EAzyziXLIqm9BWG0HkfDWN4dLxA11aCv6LzDm6xq5LU2hy4oZttojA/ZZNPN
IkDdS1mu8kwmePKhvQZTNtllb5rWrcLlDsphGggptZVmRKxHyPgHzuP0LsBvlsbA
RBH9Od+z9QrI5uWJw/QPd5R/wXgftn2qFFeVHjVREFZgAy9xtkvVXCP8NpSa9v2C
PsxAcfMhhwNnkZEHzhmTbSt2S0GqZxHr7dnA+SdkXuZAkn63cBggojMk7FhTX46z
3r8GfnINXPlpNtPyANMZT2DKwOuy69/yXsIPNrYW8BjAmeakVy1YPDrUXJnuyzTj
l0UegntPDs2wilnu5X9KlJ9MCtx9zczJ4ORYkhFj6X3RlmLNVDpc8qyjo545jcED
+ToOBxCxRrRmyP4KvEskrHfZ2a7O2GkQEcR0KrB6OwUn7NFa/Fe7CgRsAQ4WsLbI
tWoGfuwCSGT0HL14YEJ89h+nXZKLiDJAbkNWQennOZ4FfKieoNRUhxMM6Ag955/W
KdmdENtF02mY3/W8kqpmVfpU+pYtJnPwDUUOEakgVnqJO3zn6zv0bIA+OsTvEp8v
t4JH79Ks6lq2TfS/Uz8if1kzcEx4ZZFEZwTPJLKy8hTZRowfESuke5JrQMOj68VA
zOARjmDYoLoVSLPS9pH8V1IZc4Ravwsc+VC6YrBqQanLONwd9SS2kB8sFS7Qa42Z
gyO1h8DntLkGoh0mOC2uVTafCb0Y/mWX+kFBpiISyuNVrna9xkbCH9tonShJfvaM
uHKZ0s8DBUcJ9IgkOpmZD+5jM7+ApAgdoZ5FIgl6MMSgbWcWqqgUw29TRMpom8Xe
ZWpMtR047tsfmhKVqUKEhUex4jL2bkSf/uaBzccsXDTMr9KL9mN33YHh7E4ZPPHQ
0kPKzqg8vssY+lIUDCMoUGEifYDrOX3eJ8x8Tk4brTmkL8QD2pE9Xx12JuObianq
tc9I99tZXKMYTt+6kjxKMvn6lEKXr5aJvX8RL+gDHE8VnETVS3OU8JE5Gq9khoMw
dZ8N+Q70IcjTLb6xuYfKUD+6VV2PbJMy3dR8TLC6HJnnnUNkR8LDpdZ2DV4WIjmZ
DSt0yw1cnIlP9m0haoF4GdlDQ8HT27Y3vFOCc1gzXZMHBb2iZNKIHzfh7soPaRWQ
s8a2pp5k+7f9gDVsHKT85ve4tMmE2z2jTfY8I85dz+P/yoQ+N0GBSxZ1rwj0sxua
ssBXzDC0PnYZOvOO62ipkxaYtWPj8AkiGM3ulSLs0EjY3x4ckG9DyZdoAjB7jUWp
bung2a7IKH8gAAKrTJcHdqdqeh7J8MmXU4I+MTLnNQGtl8mMc3WrLVXBzTZyhQ7c
Zl2Q7oT751dOngnvotW7K1a7BiOrOQak96nh3gpDX0d06rxtny4K7gcx0Q2okIRO
Cdbbx5XCKBckjea3XsOD8YJ0lfqYi6JYPHcIqp6rUomy6oV2Nl7Bf9vILCTRAzJu
QUkvKZmwMDdssvQK8AWZgv1+QPeEzIBFCTUHRCjGZurGL4La5PS4w8OdqnlSa7Bz
1yk7dZw7oa8L8xRoHaSOJ2W3PNGO4czx0AwVpZmV+qjZj/2x0lq7iehivkmSdWjh
EEPJMtOAEtXuCM61y0NtYZC6Yj0umv90jlQDjXA10R2uBS7PmSJBKXp+aB1oE1dn
L3xVCnXhcs2P8DG3I9cQPpBYsocy/JnE1MaOukt0nCJDX9NS7FFT+IGmhYHrzzrl
v66rGbJq6X2vSgWn0Jl6C5t+Hbsvu/Yihjc0PGxEuStxjOpItbAdcfxOj1EoHae3
VTjiwAJ/pnIEJ5qLm1J7/AZN7FUgqcG+faQtFoqZSK2gKgVZ5bL6h8D6rlGLlmIg
23h0njtDN/Pn7Ryg9rXYmPxY3QwpwfSiMiwPYjSogOeRJrly8hZUhviaQPKTG8Mg
DZ9a73/PN9JH77cf7rJM7Q6ag+V9JmykafQ4iL4pyZcGJmZsEVyw6DfD7aY9dVpZ
5v3fhKyEQykJKc+YVqeUz+CdzYGCSGkeLvCUSXZfQ8Vir66TUn7IcTm2y0xL8bmq
M8Y5w8w3WsXwZxALVtkSeAXzj3WOmxDcZ6jlkC1ESTKnQnmWSFDDVQJLt50+Nbko
73/TdLvA4i7Thd+eiZue/1pnaDLNtW8VKdVedJma/DKT7xq/DssgmrxuLIWMvcIY
ihMsc/VXzzKT3JYzUCJVjPm9/Y/oNDx1VNBHDYO6VihU401BBLWBVpvRoGtyZkiZ
HHAPGWuFKt0UYhtRJ37D1d2n6nBsFoapQE9MIrAx8ZDeKJxeIRbqsJqM+FTnWfQ0
OZrKYlvak0Hg2+ObPqYGmlyKwiMndY9eqFdj3hdQ1NIM/5JlXdW5IraHAKwyxMh6
zNoOzx0461E61O3U1lJAzOSJME2Jj3BR/RIzEgeb12/7m4JmnR9k7naZSpT3Qd/g
Y+2tZN0hfxs/FOoo+3fS7ic9Ebup28MsQ7B5C115RIjH8J+FboV+XPVJNGxnONwN
wA4SscA/vlDwmYgPOFC8rbA7lhREYmGlwrF6tSk9AMsl0ku5JRPDCyIuWxNa8sDC
OI9a1B6zEclDWOV9oI/2TZz5UYuD4U0W4wKka/4bhMpWwcSvfNEQMSUI03Uc01SF
2oUbrJIB8mzNFufhT8NRkbyCSSiGP4AUF5bMoRaU8v9+vQ3MT7ifAxMNedcRc86E
QIHJRdZWK/hUESlLcsLFihHeNN6fZ5Q/Lbl4NanxKP74c0/wg5zm+0XZ+ISNXfA6
dPXzuOlva4D4nHbX2+NtUfvkpusdz/sAKcUUUyq9ZXbOAACh+3j/CT5GWfaKGKJL
W+wWl1xhQ1+tOjJT7wrTcCHQe8sBW6fsyeQCn7Dnze+CmA4j0kAUsw32YkBXWW1E
/FHokExEIMwlA2a4YBWgM5ZH8baGbiV7JpxRgsNpLIgOs+dCJEoiX8KNBVAmqdOq
5CC2OhZfFXIE33UmtL2oA1+xFZGt3TKmWuDMSeBxuViWtLQR0+3tgBbS8RYYlzmt
Y1e/x4FKH40uzQkbV+XPiSFjsZuEApkqpcxR9/strkwHagYEqLAvbGs0scwUi92H
cVh0q3MaMxszGBl69an6lwYccxwhojIXFhSqAolmk6isBHuP3od6NFxPSDokhJTf
p8vekSAkRImfbB/pbQA41YAmma31sLmOWNYV+YzoK4pIBa/qbR9DOZo42gHZEPdQ
htniAgIsGosM5CmP6FjUlnDIBZGSkK3S8e+tBXlNDWBtbo9Lt1LxpOceR0PHYY08
9QT36SPJCdTqvpOMZ3FouQgbx4X0noktkKgZrG+GCwwPdIyiAepLcTTl1FK0BsXX
7lQumF9pWqjaHNMQdVZW9KIvB5U+mH62JO1ATrwjf4E7QdsHAHMfUODp5cLz0fX2
SMcApGampNAGHXMjqEzYYPl1jKVtMXH9a5mt9MFsRZ2Cxw0iG8FaG2Rb/wsHsLBl
JBGoruMHGesWfDpBM4buU+F0sx5ib1CInBZ+WisTvIaO1t8+XrpR+qAe2gw+I+rz
iIjkI6GmHG0WkTXoayFRubLA02J2EyCUObhK7AEPuOv91k0nxVIOI9wNDiOtp3Vq
NHKQngypfPkQHCYT2Cbofk2HfI3+c0CZ4hGLGNDGEkSVDgKahB8BN1svZbXDDYnm
gQuuWQqN571hEP7QH2SQIxbOAjqqcA3PLcFFm2ecEtVlth4WlEnSq77mWmaby332
5+Qy9+8DnAYGdi8LkXkTWh5r7/5TSZv7K0m3ilaxr5YWhGdyypH3GS/2LwGlxyvJ
s96MzRMdR6ttGXOSued5B4F1qX7C0BYIqgkRGyV6euUorylZCFhXilP4afELlXf0
CuXN+uSzQAwTVUprZypoPU+b6W3h6kM70d5/YWWnQ29PlwVekOdgttCzb5v4bGUH
ubogJvPhS55wlTcTgyMyz7uis6OzvfP9PFjtEDyqhPh6/BfwFvEIUe+yBMPiSfQC
5eP1yCXvpHASmVUid7L0XBL1lyzbNrT5/rouZKXlxWdDmB3PG+y6ELiFu7zaZJq6
iYRtcLPDUfZOrSm0uY8Ehxd6iiMPu/W5NcFfjI0gVwpZ+naVyKoAdpgRSTkzxNX8
9rpkBibdfre9bJ4j266BPaSJe4R3zqXZkpN8vdmj75fSvg1PcvbWUStpVT0q7WrU
r4riP7P+F0lT5FKKQbS7C2Vi0oKp4ekWPzBRBOfQT/DH6g5ocp82dolqmO7vnSRZ
UFY4Gfq1oMJEs3dfq2sYWq8Y6X/4z3SVrp6kMiqZdtRSUbcOjSuVWmVnBGBkmfwX
XKfOX6uEIgZSKIajUf+NrIgWn48nHRbIVqV1fvbcj/mp4BVpvt3oQZPo9umz206z
nj2yq+l3cKEMJ521Gs4gIC+xGBDBc+W2QxSFMceFf+kQ58mCt2IwuI7LdML/olS3
sWyuxvGNwGd13xKPeFIjzXO26vMUmELxQmwNVdF7qpqg31QO6XQ9/zLeN0KVXPH1
ZZ9nmZEr2qmaw0eLX2HBe7zhTv6xXW5yMCQQNp4pQmGMiCQva54y48m7OEJV5BFK
+WDVXAqUQPUtLXCcm/CCuLrQSpT032+b8keucAXnK3/U+N0vZr9GsxTvzJirtcEb
yxXabiZEOtB9TYPDQkr2gMnDBPasQBCxZEowzNPCvmMtW9RU2l68BebyCAqoBYwv
/cfocw3ybJsTElMp78fHW1rWAAxdkFQPIUjbBRZAYfE1EJe5Pi3vGVyUihPLa00P
fJlfCoiKxfT1dEM11Aw+Ind2pxkCYoLTCUd2m3/HbQL+PUk3NGh++DfeZUOSn17O
ddCuHRD9JqhHrOFKmrqU1WiAra1I4d9Ot49wctOV53Iuetm0sE+t0svZ7u37d1Zl
pCYcGd2UaB8nEaumu1YhoxhBz56C7PfAQe6u00N07HdWLGuCdDxfJ7ALin97usX3
GtHK9RqHwbV1kbvrCPwxcbiMERDjonJIyY/nJOsWG7JCDzttE8CYPY9ENI6bFadk
zA2VLRsw4FLcmgwbKXbFnMw4glpd21QtSnKGkjqJBLKIRThynaszjThjbO+E9FDY
wMIaMqaYuxKXPDocQ5H0ql39XuFGJGb3bS5OyISfkFck147L8NvNpc4V902UZuK5
1Bz1vLCEeqi9VHxVYyXN66lZnFunCf5KQQWRDlBVv2tjVkV66Azhmxz56Y38K9/e
u9AI09Qj8qxnhbMIJNKmIKw980qLVXnUBvnWFDsU44o7x5f3E4voQQlZj7nlvjYl
JDvtfkM3RaLXHZcXlds7wdUe3aRfiUnVwQsqd+WNvs+sZWJEc1TKD1IaJM5vLYe8
dZHudVnvapShqMK0QFAOQXFZ/rJfNLln393FfQbeSE8+acBz1BJ2EK0e69XjH8Yl
zLFlEmXsuRzRIRQzqu0hTOjVJv38Sg3O0IoUiMv8f0igR3jzvDCOL1IqELwWltPk
YxYrmBXML99k80jDeBhr98DCTDZc/Ug018MyozcO1DtAYX3oNveXhCnvKj1PQ3lm
E27CGvZY3aar56bNdciBUvUQ0ewenS2QSEXVCTkhz6lNhPE3RRwMQfOof+pGOpA4
xCWl6cj0Vpqx17Xm27CtFlYqObbES/zLOb/Cz/JomeIJvMVP4d+901EdR9utxeHk
64d2a85CwTj0lP3pN68LjK+FG0hz2ymoWvpjzWw4WjrqfLEIS8sY6vhf0/fRBg8e
0vrWiyoG9qNENK0Xzu2LdSEhk0Jcaidc7oImaUvLx107RL2y+g85uS+yQ87pS2QU
RidopbBp/gShftZSw8DAV2zSdb97aSjASv330g104efGfUET6/XnnaMcFkoDseRq
q81gsI8GpheJpk1Ua2afeYiCGqyvjyYM4sk5NiPo78Nqit6+C00exjauPMIkg9/8
JXHLLHDA/hurMlIvge5i4gVJwBIlqUx3AU6uZ5L9tAJPTWCCoAZLgMFv2t6a2HaO
/1XenA+/2PpPpvKUmKjoUxOuJc6e0sy7IRvoeIBnc9MAiHBPp3qR7DD6WGFIJeaq
mtJOsjK3dHNKstQJd9O1HqVHgh0BxsVc9Dwf7zsk5l2v3Ob6mTBgzzkwPpO/5WiP
2F07Z6+/c08Djdgk8qsR2GF2AKbLBDrcq8/Oryl6nNt3rxpkJBnnIKNHTraITwJC
GhRDL+0SlCHc/U0kAcUAVFJ8jwN9koOMmH7XqPmookfLFdM4oRTs25wK47HDROOC
NzL64ouV4JMUxLByq+d5sX5hBxMkvZW82t8aCdOteBi229v+BPTsb3oLnEJ4vaZb
7Ry1kaosxz4y2OANzQWOs3uMhV6W6F1BWLvDwTAwNcbt6u5sgUXTC08/n4LCV2DE
yjua900T+Ff4UdhbT77I9G3VYFCMZW1aGwYyLu0BtSL/0u7SV9N4fqkJPaUxwLs0
5RK1YgIN+XFpuK2eEYAhTIz+XmdUCm+dmnlBJxuMmvYZU6rspz84xs7lhbPZRDQC
864p827DPCPoedfchNU9UU+3HQSZ+djMvSyeXLV54iiJu2+qs5QfPcfCw4FRyCU6
lCGGfvA8Cs+RWaFlFUBo7C8244tsbCX6bk2XU+et3pWQIkH47vdu8upkBDaht8ea
zeoIvY1HXfPaOYCN2P32vCilMh34svifOHlhvkzD2hyVu7fDtbjyQR/bX9sIZMi/
TXu9Hx5vO1VqDJP5mMGWUf4GUwB+jvRuUawxVdlNxD0+VZXhZsCWEs1LSmwsg54J
kdL2OxRiB1vMtL/EwHtjxGT7TawFN56un8giEidFZ2DH9jmuFn+sWgS9J55llMJf
2U+RBSZDypZEhcoBV3eV4lI4jjGZHo5QqQWT9yxAlXyr9bzmUqjGHP+Nfo01GFKv
1UKvCCrZU6OX02Jzjepe8KTbzqgB1X36ZBwwRP2owSUlXMg5kqpVw3l/dPNvh2kT
hkW/X5tHjzVMBUaV2DKTY35pMZZDyLoWJLbFD8bT5bPn9WIoM9X845/NAdZMmHAA
oavPC71PJ21TTFAMZk6/mq/Wy5zyVRH2vqqk/DZ1R9X8ylIv4BToSPV9r3U/EdL9
09IiYruC30ut+Etr9L9BqdGFS1NnEW/tYnT2Qy91RVTWo5XGmKEn1tzvNv26GdRl
HSaepDquC/6nd1Cznx9GDhHspFKkPFlhWYf3c0sqKQNpyBCnSHTbiBn67lnd3SLI
id6EbV1nB3WV5fVmM1UsfSreTNuhJuaKwc2l0tghMgCfJ5Z9QqFnNKXjnwJjfhgi
9YadUP3wliHOI4uU25qfrcqxjCf+fYBjT2Pf/lxKfxz7rkxoGScoK7P9tD9CB3Fr
BKUJ8V1JbSpGvgXr/7397UCxoW/qrV85GV5IFq+8zbwKQincVdoSjtm0N97NQfwH
pXmo2R0VG92N8ZSFFp5TCgSxzSSGeNtYqBVzYmumz5eqeu4I9bNWduDch97/8Za1
8rXBIcVc5LwlmARqr258PIs36vbd7LYtJAAsl40v1IOjc84YBeViYZWLVUusDkxC
q+Ke7YD7t+bCEH6aajesz3ID3rUX/RXQmDqfE+11+k+3kuPDK5kmnqE0RMbVmTUv
TIuc8oCMzxkYyIeeC3q3KKCRLagYs2n7MrlV2pfUWgnjZ2tfJheNu23NqHDbp6dV
Ywrq5I7jZ9WEW8ob+5YbXp1anKDWV4iNo4j4n20XUTRUjb1jvSt1E9F+cGSsTVBN
ahet90BgLPOqm+NXGbuHSt3xN/y12INEof/pPR7I3oesRd0nroGGlZefCyxM4nie
FjAGOvbVTlT4GMNqyTB7gG04qWPEalS4P+5anUWTiOXwZH8hU7+IFO2X4d4xvCAR
5EhOy+C47MG9H+C8rs5sDchtwxYD77qcTlEcjrJrsWGt2L3hvHyCoSTo+jZ9MFCQ
b0EIEhyMk7mkbOoXCYH8dKzAgtjfFucAgqOth+k2Xki+BnC5jAUbOcaNXYl8lDEC
eHhtc35qf3/+rNOJP7iI/h8biQ3WwY3wAPuW+EtJ3oQWFjU1BHnO3n7f6jVn8yx1
GpG76nGY0sV70tCl2YDQc7edtxR73Lb4fHddA/AIL7jrKlMkPEzDiyxR1DoVycPo
ola+zTRadtSQZz91sW48oVj0+K3vJ2LypS8JXQvQmKAvSlqamRZf4CBGMKRmrMid
VqJZ0mZUoHViOIipz0AemQ7/6kETkbUuRw4WbNe6uJeQpYGA51X8TKhZVMAMLpT3
t6+Bos3wANNSIoTA0JzYgBKO+ACB5njISVlxFtSNElSp7QbeT1SbxMQKK1doBh6D
NvFofaLyyAkHTAkE+ox1nYT/OpxeXrfWPx+3xbFB/gHD+MQccpozVq3XpFIc+MAp
IAyp5RtQdPMSz7570z4DXOTWHQ4gTGwJLAh7ksSODKCkjZzRW7kr4VeVt0BUGw1c
rvExnxcBg0WXcGbNHuIXtGepk+Uvh6EO2NMXNt6ScETdL8Ltj9ugoZ+BRWNeios0
SFrgTIsN+tyj2tZ+9Mnr5XBDt697h/ux0+toI7Qo+0rAjkkvey53sAspo61O7M9I
mQpYeUz6VM0BOlWPGBsy+mYZpeRf+LVbMfuVIUCvy6vnQCpKhrgfVA+ciBgjBw5h
NiHM46jauVpWwWvlfJbHKHZ3BCF5XiyHbCOB4+KysKRIFp+lo6sjNNODwInlL4pM
Dj2zNks3R89VZVkiUxGKzWsMa0erPgxpZicpQ6hewlmPHankCIbnPTZFqI8lhrCN
xnmTjgzOgDrSX7oggfM3/ffZKlM1DZs2/JCabS+bYhdUAnoy+axuD6x72vpPKV7Q
bkOtU7HtH4m/l3+64GcoibhlfM/xCG1tKLH3pKsgHtKBj5x/luk1l7XqTBIf2nB/
Mnu359OAVV+I4mfxgdAAPiGj+wtdLkpkW7ADsAqY7Pv3ksVKCHmFs2Ks5u45myKC
s/QEobX9q/XGczsjbxolacHSnUA4xuY9ls7U0XPYA54ZOUDXHhJU81DcptBX1/1x
wsYcaOLvSasI+Z+lZ7A1dbl/PeBtljabuRb9mJjmEiyXz8CvZTM6Jfk3DbmU/uw1
ZvtVNIWiyz0qRHvdoK8E6qnDuKTDoHZWx4sTzyieIHi2XcvU8XawdDNoaID4+rJ8
Cd0L3afzaauIZglOSaYrHwONSnJUQamzvedUZIR9k+Rg2s+3X/Aaj9Gs707vIHgM
9pKXgrplNzgH1/cy4S0s20TaLZBjETXTFcVF35MunIGu9XL/4G8L5SqSA47L5I2K
kC0h2yuTb+HYx6Inmn8VER5Mq2LqWQMrnbzRJJHV7urlfqyZwWF8lirg04xjcUco
0ZoE3VXgyhY9xz3f2TsQ16QXgCqAsj0ZApAxN0jX15aGd/RUUamY7/3CT1ZMBbJi
gLdo0jAXQiFr8H5v3A2aPtfqmqkxcgWO7G2/SAOn17FPRs+L34rG1oYHQeOoIhGr
ueQ6CMrKPCrFSgDnhwjObN6azhCwgV0aTO1UcmhookKSzsl6ZJzZfpVFvJ9QQH9s
I0/6L4qKGXeqtQZJOn1NBNREfkM1N/QVYy2+gq3fm8wAiCs4K43Pe8vCuHmxiIB4
95Fvx29LCogQnfNyrhOQIKB151R1d+A+OYTTdj20ONN5/443CkI9pAalS826VixT
dkJ8lACO64sOLLiyYE/5W/8NBv84HpFK2fUBWvEBgTGcTMelhpPn/V+QG71FOtLA
yGheQ/ZMDk/qCAKwJOJd1wHpTzDAdL+q5e+ZpMAqikgrEjQoP5FfjdH2ZPOs3ej/
g7Zf/GWF0/p9yN5XxvuBsZO3mvPZ6vGF3juUDACUPCkLIl+bmkmM57Th/pRsuVm7
DzKWLyvBDxgE0G7AV+9SCnaSaZnl+CXOZaQQZgcuaUM61Qki8LtSz3UtLWB+WWYD
CrM8o8cUKITxwaTS54Axrz1kWPHGlv3prXjdgmtsqr6IkbA3wNBh2ZlzCviNXWCO
bKVU9URKt8mbn9uuxAanQiM442l5f8fgU8SOkHJN/r2dr6vxMem/YYwC+58wwgE1
xescFPZsAWGQfkE5NgDguPC/C8W6OA9bss1KD0+RfLdJfiokYr/MefGXZr1AmgoG
QFnMi46jWKzSJmTtQml5/m81GEYSlrYeUm3Mp9KOC/2u8C5QFc2mUuU5xznl/pw6
Y6a9xkNYIWrRwbW2dpFUMJWGS2LCLwhnOGkP3VF8tCgjoPMcmBgh43fpi5pU1/Ly
WHXgX0Y2tgGHSs118NNHFsnDeAOBDKHg7FHcWW8N+5GD/iwLsNTwj9bMCRxUT4fu
UhaRWibVzQ1nSmN2U+XTef5vhBEsTV8eWXtCHUQRKK0GlJRw7AL2ucFBnEu3QPDA
Na+zmj50dVWojfll3jYlQpaDVAhNpdLxe0pMKskC1i6BdUhBYnrX26t/lAf5rFj1
jo28l8I5f4eeVzS552fPwk/hRrRAqv8Q1FxcHJ789U5OcSU05c75cA7EssR5IOSZ
OSD/AuCCGmQHFMTYzIshMyBIuW8lsukOzhvwcv8dtsPZ3y3BUUBNnb+nzJlpMp8g
6yQ1XLHtfFGLmPFNsBCxU4p8Z+xj7YHkPvM9ZiVA33qGsuC2abBqBmgsrCymUODp
4WIdZmx1uWt/WBebYsAB6ASc83KSvhjW9aC0osz/zz1qu89D3ePUWstvolG4+crC
JKvcLhtaeIkzrD7Vzm3D+ntA1G1HCbnZQgbIuhHWD10Frb6qaKW+QmQjdAL892aZ
nDxqQ0bDts1p8JWm2TjY69Eejs6b2GG9mEMaMonRTRThqiLOtp2mYkUw31KqkkUe
XhcuBd92T2JFSHpLvb2X/ZQa9J9+ui0iRBr9l1EHzpeRnKqSCSmBRYVWaW5Pigsz
T+VogNW/DEzhkEDXRvH0bZBFSvMmy++y2q22rRLyaK4BpJ+9yAs9nSMZYNcaAfnj
D9xVwTSNiJxiXwU92zw3yztB1gPZaGSwVLVXXsWJdFAtoauUnetNrDx3EsfGEIsB
r/PK8SS3KPZtVFAIy8FUbtXmC1FbB9nqS128igmAl+qYI/epm4RPrLHUBf5n79oH
xcuN+1mduvYE+wKfHsIotaGTyUiwI9xDXxitJXc2Sl64bHaJIy3IcIhp6jw8YZg7
B/gC2h7fsb60EYABE1CRNqHVus8CyO65xRc1klrDrrqT8b8r++fIqixbv+M2pKUd
el2l54sH4a8fU13FUf6P8RM0ErG0krW1QawmGltGQwcrC1DlG0rpBdr2djh6rT1K
7OeqfbrkRtDL7nCTPbk8pQGdGmBvov72/aWz2F5SR1oyAdPkTVs7rW8UooR290RU
GRif2tl76f+ofdrgoRAsT/cgATuAtba6sVm2t3gPGYGDdwMW4cwHIWLa+hqDTl4S
sltNRV6hy9hvhbPmafpRo60HODyJ9nI/UtG1mW9sPuma6sHS/ZFI2T1h+G8QvJ1M
P8MhaMXWjHZVPFylTnzfyzHeOOtU8up0yUFfq9MNhWP0ACPdKloTN8Gl9vsBkBkd
L75dIgBNcijfDwwS6FUM0Et3XnOMs/Ri4OnaNU2fdKPizyq8IRNEsnYgH9hlbRFU
X9gyS7xZyrcvrn4O071quAWyggQI/2/8Ie6XNGUWv0EZEABNP13xQN9P4SNs4fbC
lSWyXvxpbkLfMKssFQGp5rHlVlOvHTaUIrWx+Ivz8efWjqUJaw/cPw0YX3WhklO9
Zu7IyhQ1tfVlA1cizO/rM0TY+vUNpnhz8bGjLyUdd7TcjPDyEewsnSyvm5hZ+Zvt
Ty9aGdy1xlyGodB2vtRyzEg2sLtnWLm3HbTUtPVooRjVU8h6eVeEOjhWvNsS06Qg
TzdchRODVKdoUT0bKJ+4VIjZA/JD/zo7G90y1musLGS2L6wrmd8+KxhgeOYaw0iQ
KTtzgoqPFjzb8y6GBVOyPOGwiKgei+5S2CqCwuTDobAatmWfY0dBa/FDbXhYawhz
ct3pqH0eE6a8AiG6I1skpP3dKS7pVVyaD/VBXnjmv3+8mNcjSG8k71qXGiQyqLM6
gLoqMk1tWuP8iffHSnKwpTpSMGn714lcDALh75GXOcrMSi/VxqCekhBdIYsWALhT
2x+UjKxAgc2yEn1rMlPY3rRysHReuixkiL/GZuvbMO/Z01daa3iqvzO1JpWqBjMJ
N6JAsXMDbd5Dpv/TnWaFXzev4xlUA8+oUvvetXF/0LFdopDzu9b4LWVEgjTfZz3M
2u4doxmJyBbKNPIiXTWpptM1hQvKfhoGLJU35JXUEazqIg5ru/dsUHQFlY7R77th
nnDCKu5CEnn6XMBH29Rfk+R9Kc9dj5H3KAJ1sCano1JvJb8MzBwQ13mPPVgqaHFF
tUJMWM7YqPs6Am30iGaDJbUsfotFMGAZ+uAre7Gjr7iMsics9qIeafp+AXAaJJyk
twAYFKD5Ui8SXX+bNZP/0rlXyQ/xCeEfgUt2667Te9yJTkNKtXADkoCQNZIGCWx+
uL+dI7NAs/h1xhQ4bFLZDT9mbP6OKzZZthkpuYah2K1LGn7lRMtzvtF/e8DOmZhQ
Ts5ar+KOQDSFEPIM4Xm2xDQ9kNLkp/XAEHSHWzgC8/yu3xOrSZI6ZUrw7tne/KmY
gcfYF/TFnFvQNq9n32gbirDKL1OWaElnDxcNeWPQ2VnRELiF7jpqugCnm8EhzoEa
RXstt8lAgbOnRzxFKhhzUaP78sqOwwvKtKMThUUf49q68JM2rOqL9jYnbinj7SQm
M3tJPgjDPfwUFqghTFhdZjV+VHsNBPvNq00EhvesWXPO1S2IvnJZWjjeUccXTY3i
HOyULxF+Ej0EFszOEZ2jIDEERtrTdFBl7zFBIWOda8OaaaL0OjlbFVvqapgL7WIU
OVH37i7P8UmFpmenwV+sI/qlDSwxlWGor3zDPMnIgBlRu8/dwEfSwfila39TJZxd
prtDf7BsgtNin8obFEeoWbPc6pwk8sRXphMl2YAKbYn5PdaZL6ioRNLEim2OISVM
oGkEWAmZNqw1XIY0MW4aLBW2Ea8H6zoCg7vvTIXkNVBJTW6FCdKNZ2u53nVEqw8z
RJGRMXMHez8BxNcFegYwi5AEl/zCgtrGQ55NSMm0y2HgN00j2XQXcqFn3j4Bup8W
FWxLVgVRiij1bc7R4amu6uPzkLQxVtiGyq/TelDlA4KTDDTQvXOZp40bKzVsXqUI
0gMgxnW/0tleYtbZSFWvJ8fJ5IUWacf/G6rY0mBny0xgDyYYo8cdCKtBRrIdLdp3
r+2EoaT6jGYO3Wx/Re8iEn4HJXyGg7qyHso5VkOJTTtLDLFvnlQEDzBzXpeuDEND
nlNE2Yg0oIzYzdmXide7SVJ+GSrzTj6Zxn/LYSFvPAweMxUkupFDchYMX0M3IWLP
e9d5so4WuAnFq8KnFPT0tZ3qeUVzX7E3+o7UOfhXB+fddxRxu5V+SaGrS0TKJqDU
cNn/+PZ1Y0muvqHGp3FjrIhVdP9+cY0LA5mtdu5xsxec8iQNOwszU/Ik2AGOK/X5
7Gj2hWZXkgUsNVKk/nxH/3PKOxZZvQn14mG7B1rXzk1mR5u8PEET5VbCHoxxKW6H
Rj6fKWoYYq6pBgAWZO1jcylwi+KRhLZXmusgr+4owrkNoTiX2UKgDGkIYZXc8+z5
ZEi7D8gRwcsGsk2dniPNUzAgQb0KpDI8DDJsAn3vOAt2QvDDQ55aQlYZY35/F6DC
S2oHKpoRxynHV276o52YZ2KhFTnNlSiLYs5Jrbj6rD+4lv6AfR6prX7DAH+P/UgY
xK6wy9H0OFbDR52JHYyEtMzwkgLtK8Da7vXYRVWN6L5ByUb/Uj1yd0PYcSh91dCP
y15P2505ds7Mh3yYMxZMHu+vMewSZ9FXK5xdrRBfml/y/I78EcwfcYAUg0u4RK4B
LH4GyJqu+4Q363F1e+rknPJVnbGlkUvVze4G8gPfsX3UrxCrd6pewB5J4nUiCSmA
r0hiZxbkX537zunZc8WMmuBib1dTfg/XZcJMYtnYbPonZbX642auL595Wpme3ALq
sdaxHajovoPoAnWG/TVijWIonotXkxTxQa+fOZPCnLoO6dzyr/gJgeueJBPar2WT
zc22IpSbbwLmToGFIFRzfVl8ZMZNTbAuvmfYB6jFGoEK4TOUu+1uREA2qbgevMFi
kiAo/Lmn2YUEDvkQyDOOc2bnuiGx9kftdKPtYL/DLJITe9IiNupUHIEEUxOknDbl
NL6m8HHxRTSqgQXniII5ai/9D7Bi20oRkkyDetgrj/u5oEt2MP5dHOeBMagv0PEg
NIEHIkldjR7NQ5lpX1AdovwAwm8pgqrrOHsqZSdlP0BRiJ/+o8rOurbA9MaMyvYr
+jZZVVifWY/7ArJiQPuhJX8kAbp9CXU8g+K0Fyd+H/6y+bm1yp7HV++rQNQMl0yX
2aPjVWEKmFXJtgaqu1sT744tb/ORDgJvTZTXO7QclB1l9IGYzl+2PiBpFy3pyW8K
ux2IcWol69jwMts/VxT1BiafqFZmYxuWta2TgV9QpTzABP5Qnl8r333pi1+Qi4O5
HqI8b6tQpTqwGNp6tpboaz0ZMeDWFSQ5zPnyApMzw201GhcIhWKJf9qgdjDdYjZd
wxKzBlVyrcwJih6JS3MpZy/E85sOdddBLgIHkeP8hQt3yAbeWfRJK5BmSVTwuf8+
+IheOncy/pKtgDDQ4yaXadd9u4Ygz6FdkXI3G/jf/Jm637NGtERND/RNu6dHWTs3
7dpqdCliv7bzZECECZo7tQYQDdQ6xk8kDR4p8ZEDjAD+zOjCfsmFuVVERAxvEl+M
Yccvqf3vvBZZgizwz555h8KYDt0UZmyO+96WjaASQxYlonQ4nnxJ2KSg5ADuaHYc
rfa3oOylLXf7mwEP/OQ6/7bYXSINrILDPyrgka/KxnAwlvJAW0hPZZkNoMiVrAmw
7HTHAv8G81rGyBpvQAtLUkRCMGjQESgAHXEGcXqRG52IFsS3Q290/ibxnabmWLjw
1D4OV1xaqtcw0SVJlPvjl4PgjJdeMVh99xXoWEbg+fZ6KgZkR05AUK47SY+mILG4
oX9rHktlDVnrH+o/2Hm8hptJxDH1j9MEFGQJhPIEs42mUjZ+WAzp7fC4sV/iJLhX
og5stTF8HW5VVUDbZmj8PcRLirgQfyZBHypaVNzS2TGjlASRPDeXgGiG3e3luBhZ
c21gTikK45ba0O+/1yvacpsFjre1C9ckcF1G8FVUJtcGdHt+a0hvM0j12kUjp7f9
JoPOVRQk1aJIrB7Mz1VQR9Rd96adQhR7fSV1eKRLbKWoSKqFYs8No7u64XTJHs6A
CGCYlxBAMnbII2UA9QIuOHIGDnrxHo54XjEOGqdRpaqzD78G5lbS4e0QZNvttdEf
0x8V86jcvxa8gyeh9hOB9mAJi+v8dN/WMG37glErPISS2iV/3F9qvWYBjs6m4pfd
RQLEgm2a7/g/4HpCFViRYxBVQSe52JZapw1c8/rZ3YLL3E4Lx5NYbnB4KdWJ++8s
kq7jjdbRkT2YDBH4VvfPigondVQYGiB1RFJPVp3ugKBsieDpCiMuyI7nNGS33hwM
Q3d7F2RuhglxkaE3BpECLO3QnNA7+pKGbbjeJkEmHe/viSLLXmglBhM1JY/NahFT
MGwZUE0Kdhx+vOGR/d0ivadK1Qk4gzFSq+X9KYxQF6TplwUOikmdKx8OW4IKee3i
w7U2rJ3JAkpLFMScNv+svK/ZNoqiNbPiCS5yh50DmkrjUsuL7Z1FZITZtb4xEwoH
WkXAUKecWdRs4BcAYEpsuNTY0NNQaxZYj/9ArRMzjie2SAoa0pi1dnGwj/h8X9GV
TXySRfi2kCjR1G7OSOA+EWhnjE7CzG9q5PCwKyd/+3zPn7x5rds73/143z7oUTcZ
Z1O3mz6bVJI4/80ZSUOuuI33swbkghKjfz4GAA8nEuaNIWL+DeWH0nGp0gI+33OZ
RCPHFAnJ85lYruDWTAbsN/NT2GL6YUJjam4SyZ+6//MrPrK4Fg3KPoEXcOVBhghW
htPuu0LkAxYSEGxu/P6EFUJPBJwBBoRBKkEiuhY3qw3UoNUpOx15tyetvyljAksH
Q9bY9Tl39UnUPmHnaSkGoCgRha1DX/h0/KvUMurJI82LGRzWxVQpHv7euoYBhxSS
QB9t775EY50Rs2qLJ5eyfkuwokZ+srB//bjr8cI/3teXYl7s61/bXkQLJdczFM0s
bPt8MbzltIa9on1V1/jy18qfPaq+Gl19HUjGk/bdTZT6239dVFrsBz4YucDxYuXq
CK7M/mHjg34sik7MokBzHAvtv2x9kkqYSbu7/0Qd0PEdT4MpWagTfag5yr7I0XzE
gQakyMP9DH3M/hUI1/LoVAP58dmKVlI7Ay3vaIp9DHZFf/RNObePfhh8NSyR3Q7k
JtygIPLUafi9+X8LFPJLjkffTxIVZgNCUJSy++NgbORYSSqq575EflWQLVJqCBcE
TE3aVCgCvTWzyASVN41Ymn2k3sdOvyL/I/m3iY1LSLRoWvKCwG1Un8JitC8514d4
uUcz3RMvDsuPwWcMAIKJuKTRvpLwQWuz6Esc4KPFPZt0X4NcA66osj9jagN4Ruxn
b47Wty4ex/Ue+qh0jhQ91iZBHcZSoJ+/KyhwwFoFnfG7bpjTH8uLI6xDxPU/sKi+
PO1Z2/7VdpPGKgARBSR+hToxkYH2AFU/aMKSeyDGFMs/Pmz43xwt1xj3EMbTtNXf
NKMGWiwXxf5JJXoQYp9G0ziP+xqdoIUQ8MUIbEoiE1/TaVarQL/IDZMrSCDiBcAY
Wq9GuEfLIB7A2pzyEAo4VwbHqTduUgm73uReij7/v1TQyI6QOOnp1qLAo3dWoonk
1MObOxNlt0pp/+g93Kdee/pk3FWLJSTfdc6zDF3baiJ4HYJ7woiERjgVfDY8DzJ1
9CZ8mFDdfJh3QVsvYcOvOUJ/9Q5nke63b3IRG1jJBohx3Vm61D/vDvhWLp9jGDEe
Xp4KiDaPYYk95E197TD6DPs5QOr8VTRymIpowuZVL04Jr0ikYS59JtAVCp6xmEON
65DjR+Ca18H4GZXfKJiBKPGUO6tm7L0LZqJBLPP9aE6cIC4mlpSIazKw3tAcwty+
18ovp/gqKfMv1nkxTM2E4hCfe8gEnEPccq954dfFqbxX7T7G7PPMsMeloWhPLSs2
hZE5zSdo+vZZRUn7sHsyDRLhr4dqJyQkilMd0Hvj7mp5DG2MjEVQLyn2da4muFbI
G1Uvc/RkJeCGHhs91jjvm0aNkJ8cFlV1NfDnI3niuHb+n7cQDMTGXldkRRE46/bd
ShWSmZ3oN66TL3oXK/7rPYsvw6MkjEi+kPKqcxi83ujYidXqt0jhAs0KsK5n6Ji9
cisPybfEJ4+BxukRn7+H2j8dhD4ybp5Xxkt3Jxq67FuY4TrqdJuQs2UyXqNaEotk
QDZYyklnoLJwyh/VH1RmC8455qJKUhxTUKl1PtzoscmHjLqu1rhQSNXKKg+Ykm6C
5E65qo1rB3WMKrwEXO7WHB6EA/sbhgk0ZBlepm8WpM0sRe+PRQlrqPISxmqV+AZu
tOBCdrRUitsHqmxstDU0JvM4F7jDlSouvJny2ul7JERCRYZGtP9Na9JeKEeUAC+y
kAb7T2pnFCLknWVI5JiVc2YaZbOZkGIeZcUWo+tntm4pCWI+3vlJ55p1YdvNme0d
FA3ym4XQuk+KMmDQeEUqzV1UWqmfjKilHxiTLCFeWZXWOAInHT+Sch+MmZCYwMC8
FaGCdFYDGdHci0NkSxDaBlI/7VibDpVYi2dycTyqshoraesIDvIx0MNW/kdz8pNT
HT/cwURyi+d7YUGUih8Q+L2VUOaNy6L4/dmhfv2GnGSUNvRduPCbmD4DIMoPaXt+
4CQppSbYbLoktvVjoBpG2PH7KFMj2lh5BF2jplasvY1J5iKqnNu8ikMC9xNKFpYk
5OU5o8snk5upJtzcyGQHe5OfrYIFctgKptICwUOEGIe0om/YHaCVG7q8WHDEr9tx
SlkJ0zD5tc66df7P/2jYtTHNt4Zo/AWtaQ/dDo/vf/c63U6NIgUYqyIe37Xuf0U4
4U3KslbyrQdUX4bCPFxTmrcUPEEIBd+/k197CfHNE3iaQKW6UST8j/ck4EHxdU6g
bNrgc7Qloq9ZFHcCgANYkSvuyky2+fwh3Tep9wJfxLpMgjJIEwdgz+x/0i2aAKCU
LYm3ny/4oJHoDw2WHX19emde7dogCdvNcYbKCJbLUlT3nBe/niv8WdUUIeY9F6M2
0I4bfVGE9c7187V1g7EwGN1aSgwVg1Q8pj9UrDIIVgpV4O7EUZDuVokLP1kvpXKX
01QDiy1xh34CYq9cyyUTfea1oJy3WfXiRGs5BNa8j5DVIiLKly25tlXSQaqL1jA3
c7+mHOhq2p1IlxRwNMboA6UuzqRC9yIVi+gJNSkDJXUa1FNLPChBW9mLCQGwhkiZ
ZWB7u+PUhQapEx9SVOE8YxRdLy9Y6m54/MgF5JSkj60Kp1/ojvHq4jNyezYNi4cU
lr6xQQzXkHWdmzkhb3wGlOn2iuciRVU17HViWAQsP8fKIOTivTV55CKJxleDDddG
/dWQJYfM82SWOQEkCgzUue3LydK5M67r3a6GxIV8UMdwSYvWqb9o2/hltBndS23T
qPYb86lYlX9WL8iPGQPv3zzgvr04yWfpU462Qwzlar8SDodEQ6uz8yaoMuqOgjZW
/T0WkhdgjS3Ds4VWxkTPKJHKEgp+g7U7RDmWGdIyvwJBiIIxjhkBsvNxYfe7IK2L
ps3w7bcVzq0B8cMnp4o6o0xC783hl+ecT9BWvl9bWpC/FpfrlZBF+1mgSZOFQzCN
jHAJ4kJ90xk6aU9ibeXm57otM70yxfGtdFjktfSJrv0WZau74jDXvCfEd3OFnitW
gFz9ri7VmsxMNbmVXiCzIVc0ihmg/25PKR+qEUvBkQv+/DvGraYKcYZ3CweFuuI1
rhq1Alfb655zem90dqMLrtsR1VoVPKRTCR4IZsYcpQN9PnJzrOiAo0avUUQR6pN1
dSLf/jjTsYzBuV+5HHproohwX0pkyu/DNng4gIu3FNYY2QeKqvBnh32l0jUo7kwn
kDNlsDUXqy1T8+MQ34upzTvyF1EpsPgbvLFHQk79iNG+U7Nv6fUdS0dS3Ozz5yLX
zbRlDpMUZ4XlsKo1TX7UW9d6DDjXT2tD4qIZXR2SVm1NiR7jyLox0uviaXRBRCSM
ouaMAvJAXrzM+FkaxKzsGr19a4KGfJG4KoyZUTdk2UpEs2baEAp8Qxf1AVEQV8ra
ygJKEBO7kE90OqBF6dPKhQYWOW8vkGfKEBDucZ173MDqegRd+/l6fdokQtgoxDKt
QGixSCtV8GrDlOQmYLSkQuxSGhpwye96w5ZXHc6Tuf/LB1uDxUOHxZVzS2RLywK2
YBTXoRXVyxqB/tddqO41UnUmEnehe7xe/X0e0opozEJJM2HB+IEa1hDqCo7FV2Fh
TM4fC6azwGDCbM2d12UIMSSMeB1f6hL0zjYa2CiXFmNuGv3O+E7i5ac/5/DtGpWL
YyAh/YhTaXadkMociYcFTuHt8AtrixG7T3DEOyawCh3u2k0HfjomWDltvoVFTYxa
Ef73u0Y+y+eNNiElROfhcpnOn7mQB9dgS+npwWoC+MaabEuYyBQMOl6sUwIHQV9R
8aiNML3YddEmA5gXJRML+nSQw6+hQ5LDEXoMtRi99Sd05tlVk6P+ChIeQHZvbsX+
fjURY1LIp9QMVt3iizMnsHpzhamEfEcq75wRhN7tgW7sERNnBCVGc1io8Snm2IuF
mXlz6PbiCoNN9l7TRcuQcFnHW/FnAPDgGKIpRIvs9BS0vcCKzNW+Ki5PMgB3fRfl
qr4GhIxnzP7iHbVBW1qNWd9VVehfYIHXONtF5fi3NSSJQZHoOIMxUCsfXvj7u96o
0ObyT/LS2Yhr4+ciDPPOxGlBpQs7mFJ9wkS7efPRJSq9UXTQv7P+6ql2wYLsHok0
vK7XlGF7eWY6BmZpES1fcaY0iHhGHx5t3kF1OsNQmTbKqfVhzw/ASgHus4ciB9sd
S3HshPe4KYYLnGLTQoXzin2Soa4FEzdsCHIQKFjd8Be1pBTcbnsCskn1jlTrIw9L
lcIt+WZBzmqJvZeHyN5jlgLEHpe3f31qMm1UrcW1th7fEftne/3wPyLFrmeQzLV4
xkD9ZeDzabGzqvHtZhu+28PVoObFtDnns68UiNt55T8yAYhevBd5VXQ9Di3Us6Fh
tm+8b9QT2Mc4FcXaZlmpGRFfi9ci8KiHYUUu6M0rjDdWIIQt36BPI1+tMyH6Zl3X
SzF3XWqayUbO1qSBMzk0rafWj+uOCtXMr6wDtO/9nupYjqFElF6dN1FVxFF+8txR
BjAjX5SNv/5uoy/Or35rsK5h6HHieRKhbul1JAcEeO9Ubkm4DwCxqPaoCsdAlUMh
bKY4KvWKEbJdf9+PPzXZ8pJWyui0s/YJEGMLYN27M86Mk0Ok8adqcelKg5ZQAEEw
B/hY4yIQMuXGT6SqlinYk1yOO6VjwSPkeMRJ5jVn28Mas7z38v3Am60kwErVxceK
QwXfqu3OUxrC4CY0g0/efej+MiiCNn/OOydLLp+yYJARM9ePrAYI8OCUl3YFv4qq
ZpnEbc0S4OAgZ0tSBE2G9ZZrSKkUuSa/ltuw8X1JE0TZgLBGHQLEU6F5+FKOOnMX
N5hXyxHL8E1PawafSZsXcG3WE4yMGmPIfzwZEDnJBA9ZiqDLQ9l0ZtfKCsv6M1XO
fZ31tnsNkWJF3m2WQeANqR814SuqARl22h5K/XEG70etgqxPJ9Yrp6Xx82EO578t
0vlX/YFG31m6r/kMvw0NEJAxU3iB2neVqenNgw4dfkkpTQnmR2UUIfE+qVUTvWbc
Pk0KnbWtmrXe2Ow4/l1gJ3VyvwzQantOTFLd0t5Jp+t11CsfjHwTq1Uh9KkJv3Kw
e53KnZmaWP10fv6SOTJ9/HPqkgESVSmhmcumdNZ+wLgVbvecmvtI33W9uQl2+qZN
ThQ1hmaPbFR24Ps6hEn8PwPTWMyMVjVzjBhn0CjsZQCpFAGhGKplL5kRpCvZH2/+
NCDt4UwzPD10IxXUriQHbS8m71ZjXVE3PIwaJrnM+BN7Kct2XzXa93SXUw76zKrh
Bbpd9AEundCq3E72DlVUeBDF15usMjKC7lFKagkI48xl7o055/haMwRdxnKBzBs/
cdXqliAb0ymIrdxCKuKF/RZLFn4qH931JsWnc+uyMUHkoUieValOToa6kOXKrb3T
ecDMkJj/ObJO9g2pUTECb/c1hg3GzVyxuVuInsUEZFgudYOf9UKKjMPnXraYpicQ
YSiSP2aI/0HE/BI81bKiLWd/HTXf5gTv7p8FusDSHsBIYAglJ6LonzeUg4SvkHb8
pFjkodZseQ/oIpp5OogMlTCtaJbrM7OLMOQhhf6NtcObROO6T0Qf5yEGfCGRRt5k
aXGgb503CcwUDYujMKWSQ7bIZ2fSUSGyXxcRh/0YNw3zZtICR1CjgoXJbFQsODth
v4ttrISOr/PwU61SoiRwRI/bDVzmZi30JogwmdQhJ2RYSd44mxLcWZVKjJg2jExy
XZ1mRPWJ3wDNLhPeOtgZdCc2NapBlZtz0ore2HrE7nzbq7xIqzURVP54MOeXpnPI
siAuFSMLtsxTCaV6yGW0z3R5aQUbk3nHZUA/rTMX0k8SML/nZSCqpKh72L1ejReM
6+CBCcjEJHZt/nv/6JlDHKnPEaw/NwxsZ1urmmeioRSMR3ZOcnOh+ORQJnpqANmn
/MK0/aKSN9zarwhpDHRZmQOaTDZaQYBUBl7edrKvp0Ra+Sk1QWHMBvgPv6iIy3V6
6DJ4qXrQ7ov9OZ6rtnAdzHeEN7wX28BoN8dF0OaPmY7zhJYwcFfvAKCoLxNAPrLq
twRbD+ud/giuXDqir5xQLKQeoUp4IE2v2LmRdpvzOCE8MxeARwfsuSs9afEy/W/l
DTbIvS8WCj0pv4Hh2yT22vnf+2FwsFE/bw0wrY+F/7B1iBiVV5pMUsjTCZFvlzWv
rfV8X/M6pFFDyEPC5uIER5etV08sLV3FtC+LhbfCsHlS8fW8fdTq39rdVnqcP3IA
bALsCNTv5B7/SJ1G7tgoPFXJU8ZKFsOEfe7BbrZGwZF/ZVSLfuoBthJuskgB+9Gs
U+B9rpsvHS37SuoqDRSIN0XnyfQ9+9JuT2nMHVn0dHn+PFCwr10fmiizZgQpRSak
LTzsH6/vVVWnHWR1GktNlMI+UvPwKQLIzpPRf4+u8f8PNwSpeOqyV9i/cFHpQJzI
d2YljWJLP9bIn8c+4aBhEQ9N/uAa0NaSy9cE2ny7whQrS1ZKioowTtoxLpRw1JYY
aDfQ6b3XKB4+wepAOg/Gw5Ip4zl8NypQRGvj5s7k4h4nK+pYm6TK8FJtXo4Nmf+j
eEdOB61mPFdUyIeCj7/zdv5GWnT0P9fbQjBIn9NF40RR5mqi2oCKPPkC3mRfDjCx
/uAqD8M034LDhCpZV//7zBeivzIvDygttBDymwXW47qKKbD28JFTtwQ50xiQ7b3S
cpbLDUaPT9AGwMJHoksQ6dhdGNmpmqBMfuMf8wRpzzEyLO3b+ocI1tRGJ5C2oWrD
c2eBQk1InBiCVdKdw5I+tS0eabkDJiiBVamYGilE8BHuD4FUzV88OKxDifXy45nH
0tGdg0soqyKDNAl4w0IeFKd08XKqEv/AbbalZzNWbD2k+ox4BuYIXOsb5w2+aPjj
zJfrmJvc1R8PTXX6u0HnIU9r9O/PtvkUEJ2em4ZGQJuGNIQqOYAJMgwLCZIaW9YE
y9Ubp2aTAbsZJ+RSsdTLz1rqkV9QjqVEX58nBS86PufLKivgeKIp59U76rDmeq0G
CkmGgcJohDntU/Tkb8a6O5b0Utp6lE0YRzKHNWd3LYP3KGBJ2MLaabkN4rorFPbq
22vxrqySumUFQSRwr4aNchIfwwRgePOnE3hnw1pubgRIYNS8kToSAwmORtv0rRpC
rL5khmTiipFXFJZMRpravAULoDlXkgAQ1kt0o/hSMb7xuIuIKEm1wuMgvlhw5Iqe
YSp0VsS9uOfLNNErJg8qxjLD9Gx75K4JseIxlEP9EXKAFknxlRp3E0gggowP8ZsS
S9pBi+LmCgbo+IIyIRnz5MryJqCSiOCxiMAA/eZ0JwpDst3BqAwwGYS926AyfRkp
CEzLAjKUfF6LRaMThUlvxK4olXl5jcLu3iq2WyBZst0gruBqtepoEr+xhhuYwdDJ
qdzTPAxLIQ7Xstq8TjZZVNPl3771l2lAVX+mt5q7zO4pk20gao6LMBg5OYecU09B
gaYJrn1qU51s6kndr/7MOCgDh1SgIXsimIoaho61DwNC9iXzJ1JkTBYRXhhXvWCC
3LEWA28JwdUXcV7nGb/6HZAGhjEtgEspYI4ReLzuzndWaAr6+h+orNscGkuT+RWe
bIyo0xusCzB8EAdMa8W/0maPJnFOtSPPOviFeS/ixY2Y5W0G2Mnz2SUw2WK4scNL
i/mpvAvqGr85fXtO/Opdbs6Lhj2hlFHSxulXPD49gmSkwbyqlxoPcKc4MRIRCAk0
pnQT8YPVr1/CAPQvZbAT76/p/Rc0sxNytWs9UrOT3u0uLaLOykZCUpoStE7Pzk9/
imtfiRspHLeZvys5Ak0zEkEhg8qlk7savvC1nmbioZQgRqABYu2QAWiPuLigBNjn
2ItG3v237weK6LyVDSGLFmQDTg4tho6/PeUZHTSkloKMHbllNkW0O1ce2JRvMbhX
Um1kO9dDJR6dZl9EaZx28ITulFuhr6MO7rxP0GsVdRAONXtpgDkhMisx/ijHGAlg
X2xpyIYcBE94nHW+LGEvESu2e47qCkTwf4Yruwg12EXAravCAwNz40KseTLAQGHa
kDGhGPDJM/shQ02QtFW+D4gmVF0QYtGPSU4ZXfB6EDTHDRCfctuOB4XINBwa5Qp+
EZjOByv+jVF+dEGoL1r8pIX0fEjGnpmvfrNJ8EQ3cYkZCj1ZUuSfIjD2v1vVzcfV
fGrux7WMaFaH3hSpGGhgROK0GlpM2+H5aT46oe/Ojhncg46yy0/z7f3/8Z3GWz2G
pHUCRNvCXm8C32gtcFuDa+Ev2EZhZUDK5a4NRHImrvh6T2ur0sL7kTmqMOwTiTzf
TndvplHuR2ZJvW3kAgBUUlfSQi9yy6vlPI327XCZH0yehsrFOa6ftiasNDmdKAop
FVIW3nU/WlV1z+fK9s0BEZjG71LRgR50dGPqUDPLs9omJOYe+jKTGWjPOqQE9plM
P3tvf1p6eZIZXY+pVNPssWJEWW/J8llmKoeZgObpRJn0fGewgqIkXuujalN8cCMt
nQ4AJeoXt9KjtbooxJ/idt8qHvLIlm+lG1yqYyu7Ei3QIAHla7oCGBd4ZOY1g2Mf
1cMSowQ2B0iuFwb70npnWxhw1A6sh4nBm/l0D2k5TjulXNq4p9wOrdWHOKvEwWZm
80dApBrG6xo/umwSuXS1ovvsIIzO9FTcdTYHJYqWoP7KwiNx8FzHkiGOuUF7miUq
GmHSOm5vLQmJEYznXaz5yr50M9BhndcMXcmwE2AXPWWkWuyX7LtZNT8/WAzyWVOk
7SmJMej0LKaH+pI5smbYjMGllKeGWQanexBIjKr61FI5O/+zZc5UndpvFQI8/+1t
6lsa8fgPIXLI3I7NpWlsC7BAxOFXuGOJhqxFxUeXiPfODCWytvFQkkVVsQamk/rl
J003wuXwumfmOzw1+0yIgQDn7aOZlpwv16QU7ijKdOgaPAuWQo+moPQhJqFYSgBm
WHTdSEHvfj3w2R+oCTSb/450wiD6H7oRIIhYDIYi377vY2uVn8MY7rJTF2zOUijN
YJJvk+B9bHG03nmWPAEn6D8Oe4C7wUuQnEE0sWuFnU7BlT12tDT842QGutNKwhRT
27DyK/iFhmHpq4pW59zanJHC/wV6jAP6KxpNPq6X96FyjP2MrrlyB+RegPE2ig/x
6LIqfi6dYD+SFmVc2InFxvs2jEGeHute+9Q2ZcRP/p0tMCoJgZBCMuZLVbTTWYd3
6GP/MRtBxB8JM9+gsGQP1SYtMZcUJjtBWhuQtVmN+RRyIqDdD1oTbCEnF+waR8l5
KfmY+zUsY5HKXbIjieSGC88bmX0AusI6ImbQnAqYA10LaHhrWOdIzbjtnR2tLVJG
IKjAPYRifZl3xnuTBT14BM930KojUX/KBtBdqLuu1/M0ipJFAiUZkgzWDLo3UzTF
hdfk8h2Lsag4HCXE4baTXqpqx4FIE2b8v9oMa5j1YBRethcJzGO/hwsn86X8sCa4
vGvikw6QXqVkR2Ik1Ua/DdsBkakWL6R8JGPVh++1ymHK4on61eU/AdlHO3GhcCUD
oij1LcLDhaHxlt3Q/yqmQOJ/Wkir1kaU8oIbt/Hd10MmD0y4TF6hJ8yCsWdErOjT
SYebB7lZhufGgE5WIJCSEY7TDobeaKaIPXOL+WNROe6rZUJDKpMokitQx9BV182f
IUDOjbeSZr4VTHCo8XjhpB6j2zEoGbFtBXkzpNL8wjudiCB80hw2rTewX+1I/q9j
PvvLElcRfzTtNeYunCmJmuxVseia6ZO+Z67hMqzPuDVwaBQnXMWiaNSbNrC+W6D1
kNawRLZWEV88qovuy9JL8kBgcgb/evRtiq+6+9YCN9aplACHVkvzAKnlN3cYGJpT
tYsZMX0AcqmfJqyuoqtIHKBx/HSFprI/DgmPV5IvjwN8cscRTpQ1kb/s8q3qlmqQ
GYxiRZMRtlNoyb8AScqgmUAFY6zJVx2rlUMZVkKB8bkGdTAkEW9eVCIQenyCiTzb
HhTKFWpE8xVevDM7JU5CBKE7/wVASdRoFX1OnVGCU/Va30A3T1alnXtLzhYBJrzI
sMYfLohcuxN9B+uIgex7jf58S/jfM8okLP9Kp+7ktplOv8rwXhyYQRfYqabsl2iS
DWRGKV5ysm6rPDgTL8iwQsBYelvVr1U4CO/IQB8ntBI2mOp81AV9yddnTninEmen
684NGSFu+A0AuPEzA57B8kusXPn3deBq9eD/R6Vh6RtCYTZSN8SSVX9Gjdelkpon
C7IV1byFaJd2DP+5TaDTy+nKBB2QWs83iOfG8kxOfcBk6yA4J43rAWaawnAAXRBO
mc4YY4e1DuLyuQn97XQtoWQiSKBacx4CYDR4AUiCjv7C7i7b43zZkQmh4otPgqKi
+5OqPRCwwpupq5XI64xCl/JijOKLVB316HX3AxVyZ2OO3lXzf5YmezttugN3HmoS
q7uyxvMTJ6ZLjcCiNIUTLYeMonZdCJbUTxBarESW208frRKmccs98knZSRCLr225
h3Ej3JZezcqmver+NkylkOV7NEFnL614SJHm5pwWEE42PO66FlZOFnjqzdyM2Mzw
x8AbcUKkG/+mPqlByxQXRlayuyAYQJR8MdsNuCA9a041QtvcIDfxczSwGngvp3RY
gR1i8PleavdGoI8FLCSf0/SNz++8JHUm0Mllaxk7lYkeMwNOpoch5uuB8KBlo2wm
4Y9atvGz3R2lcReUDRH0NiKeBTZ29Inu6KLdTAkZFUHHejjdsD8T8h9j3UGFaE6s
iwLRLbafHhsH4EWzi47gd3Xlpy3o7XwMz5wOxFwsGaDfOz5WIiWqTjOy6oRGHSsM
reA8kfBB4OFQla4Aaq0iCKbOKpp3iZy+MneDKdKBwncGh24PlkVbBVS4VWsNi7UM
jih9KQpuPGvt4DQv8y7GHhDLe3Gqb9h+3NhSR7vs8AGg2qTiQQ0ciFJ8xWE9Gj3N
C3x5kx77b6mwmIHBDMqHskkOyXYt6KSqxrf6g+X413N95GnadEI8Q/O3fXMcww6V
DOWMZ5VX1XGf4MKh1A0evkhaup7lnnFvQEQyocCYt8yivJ2DBUdP35M/FIrKvDJZ
JrMQy9ocS4UzZQRcuxGTNbcQ5yG/fNd1CfxYjTf8VR9ANSyqiqLUADxrDsV//tOC
nbxFaw0bzOnfjM/aFD30mukJh4t23gxJ72YYWj3jPO8VM9O0RsW3DcYevefFlS+f
VVm+WL3QDtWQ8eUStdaMkBv1C1oyyI+GqZ69JrsCLaS9g1a/8YkpBROxPDGIHyoz
G7BcDL3ob2PD9owI8z/uPXL3AFiYrNvX3vQ4cNap9oNSFs7B77yk+xYPNLsyaz8Y
/x2Cmd4sPymJiq6nOA1qCcELRXVmD8KG82S3cCsVtcu45B43EUl3KXbRWul4AP0b
PqtrvWCpUkMb9evXZ3W4jZmSXxst3cJU9GxOszwxqGRvO3ejug9Fzbjzwc6FoCg5
gztBUhIpveQwtjMatVslFIoCCGJxVUACTcic97M0ITDjqjx4nReOBeSInCy942dl
VuEgC44RVEn6qVp5xskG2PTyhavTYelkBKeEL/hyx0DC3a+SfK0FxVzpoKI1o99c
cMgBbGDI0x7+iaO8IW3YCgiIl+mbwIpCtFv7ri09yQASE0OD3v1avmqM/gaRI5Os
Or+S1vuY6P0F3L7abw9CzyFA9PkdXhulA2K2M2QidxYiE9Vyjv9PTOM/43E/hRdI
AmeJ5DM37j4cFhy/uBoXqQriBiV99Zl6d69Ngajkv0SgfM1BSGtgoAyvVsK/Z9yf
kWX2Z7fPyVnCdYCKbjyqwFpvuY3YqTl8K+fYs01a8bx15tTaPXWNAJYfFQc26W6b
dN3dyMHVxL6042L1QI1aZJhPao3ynIhdEu1l4nokogMZFWg6G9nhh+vd9AjKtjif
9Kt2W8gpS3TSMkO9p5sIBywiUR1MqbyFdZbKqTP3eMDZBgOEPKuZJnH+AhvpUgpK
eoZhvsMFMSbTPgjPkjjqeVzwJDSy+VxCSneJDkdfHJ50MNO8IkIfi41TtzI1pOOT
CVKagN5jtrzcGEvFuNoi4py/BM//JtkOaQyk5u6DIPRBS5nKBv6odYpQb7FuSZiV
imu18mgJ3BtAL9BR7pCy/jBezxXLMHP/DTKKmOubk/To+DrQK23XeiUYt8YOrbGS
UEBJiGSE17bYnsj7ahpQRwAFDlmXWONgGhgEVsRC5dCvTaBnaSGv6rB0Vu9Y5EyB
iYiSkpKltIBFSVQ+Vg8AsznHFBMOZ9Af2uWCqsPgJ9OaKZfD5aDKPm+pR2qKDabH
oSAF0Lho60CtzZZh7jf6/cSpQj2ycJgh8d3RXuRqrL46LdIEUIgy/laRKyEZCjiX
tACEgJg5SrQq01AQX0hU4rDg09PzGOwd4xabrg5NGyT3rMKGfW9tPs6UenZsAy1l
cm4GmaYYaiw58QkUBNTQHBTG7L/PZ5t1kfcroGd0FEfSb9L+gNizdbvY2oDPy3aX
3mWsZ5xOT5EGNkcevLzYO7PbSDIpMFQ9NMNJq5Dhpo5J1q+PhPwW2WmMP6JYcXLL
qJDrYbOOlYRz0fk8CTj9N3UBm5ZHiTIgp/Z1SPm/OOL6Dd56Vgiwa4wZ/mzNV6WV
JhbguC1nGNIpfASJaeRylpv6mFWRH3gSpRcdG8th1ELO0ho1yiHNRuEIe55zjsYE
8ukneZ+JwL/LyWgFIu/IbbvkLtny6t+5eSQuzDYAe/L8sEUeDonjsbKq4x2ZFYUZ
xKQuZWNqGkBarh21nbbW4MBMY8nFwOVWGdTzyzxY2MgH7ekksYVvjBQpuqClxsAK
v8EG7yZqpsC7ZCRFeQ3PBdckfCmZDfAeSfJD3mi6V6dor9s+gTHEOiNe0+QN32lx
AkgYjoQ679owmLf+e3lTPdj0t5gsUtbSGLbnpvh9SLQhWfJ+O6zHY1OKmZtZEcV2
aPx6WyHdAXLuN39448ponr+3ngURZgFJE9cq/E2sfmfdcgihUYfT7I2FctAiuMuS
VgPsOJ4F3u/t9ZRq5tVNAPv8albyhPJZw5ycFGqEPF0MR+N2rZa6MHGNM+I8QFhJ
6kWWEDFYIWk9jKoAcY3+Cudv3/c2Zlzkc3t6lllC69fTk0IUFaEYrZTIuqGBYNQi
qBq4Qp3inLCRzysaL+LHC8BQG6sIl4UHPmBeRn9Pl2UIT5YPQ8U+7JA5EQpT500q
Cz9I0obBgT6IPMamp50KlVrEZGyuEjB08s6aVSbzqN1Sy6edTrpP3rTgk9VyvKwO
l0PPNjLIqgHpuY1jkNutQiCJyxFb8mJMWnilEdnPhEbk8uxOy9YdyBjJLYWoF4LK
5gNL3PJSgXjrwgOowsIR/XPvLh5ZbbiIZNC7UFssuakPlNg0rEFMzqh1EXTTPnrT
vfBxu6gJW2U7jJeeWQ8cVOqKHYZNcszk70nabXEYzPU4Hh3xENJ6r18NDYrAx8SC
7YnewFMwfcNf6E+sd5fXZebjFOKmOmXUVo5E0aqrZl8ekGMTZ7S54+k/EcBaWm8H
TGhivFGDk7ARXZTNlTcBz1p+rqjNckJ9if5mZDdTMZ3qjPq62s3PE9edSG96p48S
4SGnwjg7u/3WCjhQ6y/KD9H2WiE70vYXWKHvI94LwJWxxbYiWLWYjGN6arYyUT1P
54Dk9Wg6LxnHal97LjDGNhrkt4RHMMnkY17ef4xWewfMYR0N+Rh9Czi5hXiTONsM
T6QKmC1QGt9MPws+fjBdZMf1K6Q+BEKwL6MJQNnTTeW6ZWLYDc/tbhgntLob1R1s
D+9DAwNUgZL78xZw0vShFUaMgswqWbQTyfiLDv88D5gEcBcV47OiWWCkKnLkMxZW
7dmCDG2zrEYD9UbW6SGd5DL56VLBhOY+o0xMA0KlP/ljJF6b5pGnvG483tBtiVCc
l2+5adnRdJLt2j4cFxLla65gjf1NlawU6VD6fYg08XxI/G+M0/1r+NuHtH0iobJM
CKH3v1yUTn6IUZynkfh6S/f38EomIZd3Dh8wxdHfyB3uNdD/R/eJwGNoKnb6Z8rN
/uPp+eRQPOKgZnyfOr0vF6HU/tHkXROt2H0NyVu/avOWt13IURPXmcOIuUzctK1U
BBPMWco7nBWSJjzziMY2BYFT74V+TTMgRBtY9h4HjhnrwBkXQPqeVYZx7MNkfoFj
UVRdKv1FeDc0A+/iFN8w6RG8tjT6sRAQFJmoPcaBd9gE22+ngUt1kHv0GckJJ3AW
s1gy0vyTE2oyIjxPfAZ3p7RGIh9tMVlstMufHf6RAg814HBnjBpNdsGrzaP83cz2
qdZciBRma07jxVkUCwy+aIOcKhiHgPVAqGdBvG8Bzsjzd+X57eehPSiqGcmGJbjx
/X+AB9vls+sG4/2w6yKTvZb2WyGDjw5AXn7PSK7jgQkPoc9DxGyVRPcRJ0hCHxBR
6hd1EqKfjCOZetPIREm8CQojmGSTN0sUEcmqHycvN3dTcvHfdG6BXxBNB+qAmHWp
0MQP+T1WkCl8ZOsXXF61wrl39Rz2UE6LC36kVsarDaS+rvGTtVF12xenXNu+FsYW
99PrS9fWbEyKyPXlRH28/GFbSoZq9DmGm4d6cu0mF+gVi3UXpbI5jwtajVC85NNF
LIel+PXjiVUJfun/HsxpX1co9ZJGoif6O0IvlzqUdkRCVD0jQANSC7RVY8Yac8Rg
8mV6Viq6m/xaOZFz5KI7/qtWQ9zrUgQyqSV9AxciFk5MRW0IgkgBBCjKmZQCMcjQ
YbLaLFnJvXRPojbannoIWk3OlRvEtg52TO+aay1IZvJu6WbkWMx9DgCFhiyGtvak
GhiGqXRQL0XuB0m3V3u6qhsazs6RcZyibVshxCOpdY8cHTGEgIK2tuDBNr0scpij
7AJIG441dNO4uNmzAjcIX0Dz3M8tQiNvcjirjVS2i37KerelrjIv+yF6B6Oy1YlI
xO5AjfR+lCg+QhbuGyIVwNkPWF9dzMsFRXRAvG7EvxA3BorF7odlrDFvz6xBA4dq
hqCCQRg+ODpuwQnJCbQJ5B000tYkNGBSwDtFq4aJumU3Nehw3k7+shpDWIlqco2I
DG4GOKM0nlbcMwdbE8Qqx1jXNfw+u1SsqzwqPcjysiyWb13fkCdxNmMr6eSnSRy+
w/GC5RL22N3900SkidRr8xHeMykX5nTjKXnczoRs8FvCS3yVvg1L2UX2OTjMeEuI
RZP8PGvB4s3cXD9OlpBgg/dbaThOl4DF6ebeB+YALG0JvVoxgCy61ZsFsqQxDvPd
Ld+xYJ/T2lkxVvEL3m3mJFj4BkSOSVP+sHG++3q+uTFFAPe7Ekb3TrE5EJ5BLAEu
yC20Vqo87n6u0hTNF+oR+v+gwXyZw+TIYiYfRkFGwefpRA6MK7DUoSfNqk1x+xAm
R3vueCOUN9SM03BeZ/tqQlblzP04M9XQo9Gf3Qo8qWhk3I28chu3AcTdxqe/du9Q
Z0fn+MYMtI9yO4egVd1Q0sCcBlW525B2E3WIgSOC4BX1BFIfs3wWurpUUCx6KY/j
JuD1YmjqXbZMA8h7i+KbvGKF2eJe7NOAF3eQYSCS0f/DWcsTt21/Kh5j8lUr1mHH
wjERCO5fRwRkLXykrdvmKy+XO1yEhFncBsPLJIdGnv8Ee1pVffCU+PjXe5aGBjnZ
YMC4YvSESwY2BXjKzRXSjpprKnbFaNuama79RwTjetVwNcOkY/4Nq81nmmmrRrbN
8Ht7eCfxFOG6sDk+wwS15Y0wEsaaLRqbmMnb4+pb1nJrUiaxOEGOx0/sE838orvw
FQX7gak3mIvMs/eUXq8tY6+wKNa2xFbSXh6zApugJpkw81E9AbM5lnHTfku1nqPw
dNPiaqxuispacqnSK5oIEDhF6zRJ+aW/bFee1LaLCCM2DB08xkD41X+AKJ+KJfV1
q7iaJiiWcrN6S1P47OIC1rXljh849uhucWAXQXihyhb9Gmmh+ejc+PP1FT8RpnOA
Fm1wnBNCLyGJSNjYhLMHA782NqJS3rdYT8XEm5rt8vhNTwQAZHT9W5gw7fvCmwsC
xCMBMEQ6+oXk7h9vFo9/56lFI8cbQtI1jaSQr/M2ftqd6u4+wqUmUx/+9jNMC6RY
DHUEV4E+kdnx35cqsZzZdQZEcUwnQlEnEcOUE8K98dhi9W4w3YFxO5BhtXIMr7Hg
pl+u2cidsLv23sfpOtn1NZn6A7q98bIrLK1FpBrelfXxOg7smgvijIDIiT8TMcfm
DMgKWwDc5BkHqiQ7uL8ykRz9q9fLjhRdvwK6OeMZ/NWB2o0v9bDA3ctFnmx3prnq
a/+D8balCdKUG69/jKAVHuJlOLafQvne6hA1F+/eJi8EZMVZn/axqbbDw04Y67SC
/QywgJyl8HhO8kxrro8JWcmoJaD/TTe5xnBZ1YrhevN1/JjSaL1TQjmRnsJplTjl
IS6LL883annjmzgBQNCidJUnecLmaVr/B5mNqNFv0iZoZYgyhVnyWu2CJbUQ3hB7
qQg2D4jatzXlE6X2Dni5cITEJCnKoqFPkgGQEpyCTpjHvZmd0/YF1k+nMQ3xTU93
dXXZSMZLhpE2WJY7RNPB85VANKNnWO2syVyR2SanVJgnQXdD6TJ4AL+XPAmi40Bo
2Z5cKn6itK1MOcTXsVcP05Uh6HOO3k2tC9zAdT9uea3J6bYtXo5VYH7PRFMDPlMV
C2ip7tfmSRFrM9JPw2jUqtYK4cps0/NSYxM95rFhyy+i2x6Pt+mxck0UcXrA5lvv
n0diMfL9G5K56AqnKzQbiQE3vYqW/5RgUfD8WP+k9Fp0sqo1noLm9jxv6WTmk15S
7ImH7W/s0XxmgHnZlazqL1M1HTRxzB3niKsP2XUUIyenNYL52WVt1HGfwusPTrm/
MCYhHbug9lebCj7BYqGP8YDbghxBGtePBhOv+9csS3j+GyflMFXktpFiD747aHJ+
X9zSTH8vzOC4SlEqc/OJo3Fl3qPfO9ohBZyjiMTfgt8c2Vcl4KssBLnWDmwdOoRv
9UZ6y2ludS1JzECSQaIDL5KWz+buSnh8JaTLNqAlXpis5hVJTbHWs6pUH8+4vRLa
bx248yY0Znug3+YMwIqZ4Yt+lUBVFwH/GSEc+BU0lsNfrN7jqQ3G/73+YeN4wz2v
z0+Q7D8R/EANAe9YAMQeHLQe7NkyRt6gsXc/tqEJPGJOjoBulXpOPHv0zpF1VzSK
FqEdn3fsk08fzzx1rXFJCA6Q0YCLuK1nzn/BEsloFj4XvpAcXRcjo9XGhQAqNagJ
OU4Yvl2Ftmx+Sq9I4HhzEHCueHpstwWkkhZCrbhvrLUCQ0U4MDY2im0FtxBs9We4
FP7ET2b1Zuk65nGD+UXSuJTX4Qj7EuIidiRg6KIO5dHLuevf9jbqGRYsH+Wms1tv
jigbSO+hlFcllHtdyNTqNtXQ9CA4SIoVdSe5xoUhJwfxls/BF5lObWoAMYChoUkM
ZbmgrrRfWZwkkcP5C05/OhU0d8uyXqZ/GJIBmH0m4uIQukhwJUqDHJfc4fRut6Ix
fIY0WFds8MNx6X1mbEDgPpgGkO0MdY6ErkHENWXmL+6tvcOgERwOW7vDhJenytY/
2S2s82gfg0gxWxDUrQ5BKx9q95yxXEeJ8LIQOE8k43+/bDDyJhrT8vKdkvG3eiQ1
1SXjWigMXQ+33XNnil0z40rAbPLjtuBcbOQN2I2bxRLc8dBmCLbLM+BJAmC4uSfl
9bCP9jcu9zOpaZvCkVBxYDcJMjHAODWVZCep5+k+HzUcNLIfTqsIuMGnF1gU7KDU
ySKqIH/ooGmKi+l1degjnDz5LeB0BZ2p2ymFsSkuTaJhTUolRIHS0ruo2azIQKA3
IteE7JDyDRbQL8zqjy8wucDlz4KifObfwtUjqbjD1DqGNS9J4FrmrZHv/Bt9UqD+
xRSnTPwRHgmXpSni5nC92zBMISEndrwApoJnuR3cHKz2CTzCsib+GkEWXU3YFyWv
ULUR8v152rJubejMospU4eY6bv+5/H17wEJUyiG7J+xhUMVfZPVmxzXwowR/8K/d
SOPrmKlkvB+YqIZ1BNHcSBVdMVsC9r8wz8oNmMt4iN/b3CeEI9JD1NZ5IFRxb/vC
IIVf/WmNHLOY5ANeFJQnXXu8sESLNrP7ETtO3i7A0F28t5vh7jYhJZyWHmr6fVlB
83dhcwBOxFrIDFDKyWtXOMeAg98BsMrjyTq4E92ajnwU4ArUaPiMmG8MSjCTAIhK
2XKrbpWBncvnJFK7W536omBIjibdQuOcnCrP2SNLDB9FmJfnq/uhlWJZ8B9sjEXx
bBYeCW5fFmNSyvTai/eDQ0r/2rU2Eb8Be0ZjbRiiiPQV4ynVFEbOQOL44BccwjU8
U4sA7oQFq6N4NeFSN8N3WV3M6RnqQdclLowJc2UP0yQvTf5eg2tq+7h6RvZ/zqKB
HBTrLEMKHzaG/siPaOY3X273FqOFAovT0yA4xD+irOd5Hu0RRxXPq24JYFxevrJr
MK1E3jHFNe5oWM6Ojr1VTt+9lGgI7WmSwtDJKUWazCrcoPu+EYGVyGdnv1TS7Ygc
Y/5ZS6gpDAp8YKO/41Mp9AY2d3yfsZivulAXGvYhkIO+I3mjZ6RYdw8g+PrjnmgS
htO3oJ6a+hrgkFjC7RE7E1sjEM/5OUPvWMjGpoa6/l13mm5ZEk+e4b+0Fk4mmIpi
dTooSTS5dcAjZgeZWwncX3uLqo4chyJK7w8K0GIjORaeo1JRYfgm2m45exbfAk9h
qcaK1SMNEHVVxw9DDVHNRPIqruTJ2oOJ/Hfl3NQtGACftyAGyoNRkmUjGtuLsjxY
iP3EMr41AoJEJFCMltbq8yWr/oESgJQUV3vKf/J0rlmU+kar+3fozif8bksHni58
aKBACEp9AEPUm096aupNPLGQMXgc5bfpTzfZvkzf/zy5RVGFllkk4NQgSmUFtoRj
QVPg8ejZpRirotyjZwf9ZLpc1yDhsw3Q7cwkXxSqBvfRwanXWlgI/Ed2jDArurG3
5BCcIs/0TDfRF5njj5gAjEixGwsKsyx/v6yl3cpL8Z2yDFv9FMlIchNOwaDCcU1b
o6Y0rgxxIkMsswuqBArpojvG8g87z7TUtbCXQ9tOd8WWysl81eWP0p/UteSxnlaK
ebuyXfQmY65W5itzQDQFyt2XcZmekwoHKj22/yXHXbM3/nH8+OZ1USAJndiqhjiF
6MaeRyG1lGFHZrEPPfW8VUQp7R33qDNEnkqiy03eIVgU9RPGyd9SGXoMdO5dS6V/
rFtrmje2jJr9k+DadvNEGykh3evAZnxv5Q6215TPl6dRs5tsyLIf57ZrjBtxwtM7
LG5AmXVUUTgY43c9J/LsyhRdHGaCLWS/v0tGytsZCs7ftDOiuA3aSLPrUjns7BM7
+gbj3ev0gkAcltYgbv8WohA1kA91fZkidVMj4KVIVwaQck+FifNhcDaDHEQF/xiU
Cz4wY7jW1oGaagBgRfQlojDRwkkHma0UWJPkfD1jo6qjyfVpC2QpJh1oDvjKHES8
go724DzMHut5W0blF7xHml69q9Rm9RtjoDi4erMvH8hpp5A/vcvYnyTYe7TENlpT
Xmm7L7dnnszng+J1Tjr3IEn9R78rxb2m5Qtr13uJ34glyBHuAYBesUmXo6bkZ2cF
GtYkNXawqTmTyAt4r7TDV0bi4E6QFY9w/wFKtr1P1+HMs4EtBckoNNb8PeKvddKJ
PRFloFhCeVxzuA7W6Rj3ytuOFDJI/tfYfEWi5V/q4KnpTmH98PEnUoJk4klyjUUl
8RcZ7qmQUG+i4wB+NJBL7HpirOEAhCdGrl6eCu7ubTQamwjbEhW9Fyku0uCTjqjd
bG2OVOQa7f7ZOJXNDca8iZlQj6CcUD/6a1rI2srh19Ey6pwhfC7kpznobxNL2Z2B
BSmnZ4cpF8+Y1SwxKqbEQi6uDs3OmKfIhXEWizeC+1vsPSShqcrsV6zP+zZGHIAe
M/hQ4upq0Qxne27irzG6EDX4GvIFTVqma7Gg1rqlz2terDqaUxeKB3IS71k3n8eE
myLcyMs55mXDggA20LliLS9nZvCr3o0Ey1rOfflnJ79r/L9CneDB9bJRSoGZCS2U
73rxrXA1j7MCrsXi2bSKOc+XrHPGW6XMlVbwbPvNL9JdpVsn5QjRaZ0bHvsjR5zq
+MlHltiBok0fbDHVkEIDG5M6lr1Noro9aeMy2Cbi/jRWufnwVfXSn714lYR4LYN7
yJJZMfoVFKpK/oClFLml3yHuhqJPS7CjxE1fVuZOiFFtoSkpIteRc8j51eBpUH0a
I01/3qe5+wWB4Sp7H7saQuAInojXsHl4f4aJ9hxM/zPktZ1eald+Il6u9xu2TWLf
w7TQSsz9GqnsqcTspivrvDIozukD8Qv+lGxTDg3K8tUNSmRCElGi2RultJWJsoD8
HUMzDaBoEd4Su1Q0qoasZv+dC3fOuQy7UVy13Wq/eQJuxVrBP9YzYjV243KfQEYO
8kMmPoqiSbhhVZU0xvqsTBPiKf6w2knQ4q3+m/srYaF4V46vsg7GRP7D0JotJhyP
HuvG86uHNAG70rcgFil0b6sLh9gt+AeKzJHQp1cnas8xhzdF6rjccp37BsiDpxWJ
OmO6xZU8giMY0nKZc6jvm/6ECrGESZAdmje0hsMTM4L6apoJcNfePKUl7i3VwTE3
4iUfr8V48r/4H8cHi593/AqTdhZ1TdNijc5VncPGUxiYx9MyJv3ZGHpRCFQJfmcM
gxWjRnGDlIUCbgyoHPIFKKGdLCtMGHkD+jaYxSYlMz72hvKUdDx+VNsSfyoaE5gc
s9w9GIqKPb9W3BHVWpVQRuAGHsFJg/TQxRRmNvD8OFDwMM06XtdhsRag6CGhDdzR
EqkbrmVwOVU898FM8ZR6zPEVcQ3e0DV/nLsI0NWR+pv9P/AQFtoqxuamvHq6Fk70
wOtJjIhP4INXboDi0A527z91Si1K/Zzurl4jVLXch5uvboFo/MDCBdf6fUNnd2LS
CKi2SNWZPAA7FIpkGkcLECpmLWxknXdBVzfkuK1yos3VXE1VsTyRozETwtGYlHpK
J54IuTWFhJ4Q0peVEGu5LKZlQXe1yDJn9lR9b5l1GcbNf/uY7pv3p2BTA5drm4JM
0tCsfn2IsKLmT5duPUM4OfeWVgwR0MhM8D20TMC7bRruTAVXHUSjXy4wqvnd0Ib2
m/ANCBrzBrgltptJeRpDcMhkfVOEJTS7h8NNv819b+wKjtSygw816Sh+wrRy7IIh
fRIkvsry357pwBl5uXP8ZFovH3zDaD696nt1P2q7yIPS24oGL3QerQhcvvwFP4Tj
yCT12Ve1zOmFAYtFtgIY2wNTOjZEX2/aGcDwZrDkMd2C2SDbQJ7JEBRbBJ/xtwMD
8Ol2OQ1SNUxAtrKndWYzlFTx2/MzyDVPZyjeZQ8OQ63yyGVnPtCgCM7FiaOEyb1F
aSgS4hk8PlqVJzUnzoxJYQKx5eQ6tX2DsA01SWLlfclqSUe76k9tBBqIsy7Lt0p+
6SeeBSA7FJC6z/PIvbgOz8yBp03J/zqY8Y5qVP7gK43PMAFyMNEV579oCYOb12TK
gwY76GKAmrzRXEzHywrucTDHsdTcSbzeck1fGMWixtwh8fsQMJCkxp+6q1/2DxpY
ge5WrNxMtJK9GkuTldu44d5S2DNAmU96GNr3RdKk4S9Oxej8GqA7KHZa71PR4j9k
59Kss9SU6/vvrolzOkfDZgFwu6KdAceJldVY90jSxgzfzN/GWC9AnxcwQSpRzLHK
SXwtkXlqomih2Rvyhg3GXrCT9S9RDtTWg77cdjznchETDlA/5ppojAVnXm2aGHRC
6sk+2hi4Y3rRCO+YDXVK861vxYqI3teXGyzPPQsIxPH91v3oDw41BgHc1rDKZAwe
sCk6865LgIYNB7jVYg0ZOlGu5/kJ1tQL00eCG4xLmNrSiU9XilY0YsTDU06VfB3L
3epG4TQuM6rq50oUFadxXyQVur6HuJKBJGjwTTqE6KFtFj9vrisv4SoT863dZWMo
ngHO1+IyDO0ieYIxDS/TWFbVOymUHqnPmo/penxROdu+/D13686WB5DkU2eYGPWZ
L3Sr63oRr6EgLVqL2XZ8WI+ChrEfN4kwYMQ2YH9Va38JQ7oHgBIt/aZpfRgbd5+7
/2ZpD917jVqA2g4x9DFPKdWgsRGvuRxscshP+VLhDUyhQoCSk4NeTqlLWEgXftB2
0zkeAHGh34OzYQKzjTKVkbRIbtiwQQCVBF20FYG7AYovHUgWSoQVhOSgBN1WzfjG
efusgHexgavXEEAvQlsklrynDr7oG0mQJSZyFTlYcX1TGnwDn2fGcUJIM1rxIVCt
25ufEh068TVnfRmf/z9Q4Tfckufp372mwNRtw4WF2CTQgtkh5ZSKl64l0N47rYa3
0K02cRSfdo1kN84bPa8oQiWgsKTgU/aWukmlNhhg8heU/kB5aeZHmSYfNmh1pBNl
TASsUy0RRmOW8v2RhW6vnCOe7FyYzH7W35EsIA2CCJyj8t2O9DwDI5nJJQwYAsri
b6H9/qGyjXsPwlgq8L/9IM9sU+LfEAjuUHbVdMI9KZ4QD9O+V3PpWCj+GQ+8vRwV
aKGnllQ8b1HjFt66L1w+Z9+/ZG40Lotfo2YZYesh7Xy3oD/Vypb3g5ROQGy2Qz3w
ku+/1UNgGlcy/iWJvcoaoh4HsiNOfFQitQ9xxCQRVywOuRcIZX2+co+ECGq/kbWw
a1iP3SvsK2o/SXxh8d9kqnQhbnk1MTMOyCeBwI/LXSvJAORCCv3hM8NBlHB7QcvY
IvPImUe6v4T0+McLifvWVUGC+3Oov7aEFi4lF4THXxJsggXe4eWJi8uZ9u6P2g9L
HvI7h0kDFXlCyt/liPcJTP1Foa3erbGWIKeGJnqm9DaOikc/+o/wLNkM/76g+S1S
fOix+cPVluO6Wte5gp0lrdHOiUzwK4th+Gbg2sV5h4XvfeeBwOFsMHngfKF3J0iG
CyGpdfmXoB1vBMl1yflgqMIumac03Msni75GkRUbtwLlSeYQ8xlEVpyjeK87MDvk
uMiJFju2uHHgKJhqt0oTOa5pCZCLAqRw5sfafhpX7L9bs+CTpTT1KBXzvb98KgaH
Jvg2QVyAVWC1PMS4LkJJOKytFBlGNymq5Tquo1zq8ZT8QKDLIqxEolkJ8qd9zs3I
0rsTB5rnxtnDyewrh9shVGSuT1wjmjMu10k5zJTO+z2wfttWYYNvdCdl0+svQO13
MCZOy2saYWBfNdRY7rJhlojffQTUV9MBUR4SFhPZfe5mgCXDbET/59KLevR6D2xW
S+6zTUK+7qx4+xNg8G+fld8HF834XOaxU0Vx/XzJaSP9wYfsRm/B3XXlQN7mmghv
asrKY55FZw9awSZ4NBpEvq/Gg5B9Ma5urG+eMwja9J3604dR9fih9zy/1chrnUX+
Q8LkgJt4r0nPmzGutdWTevMc7mw1GeaXOYHdNuxvBPv+zY43+WmPvc5OowOUc7ni
gBaxFARcnEkDMHVrF4cL1N5nBOOG7Bx8NTaWtgOqDT6bFXq44XZxNnAyyR4UbFM1
0/5WKXUdQ/WHokayrywwskAXJrblwyqNzgXiarG7K3oTF60AhF7D7135TqBQ5dQQ
yivk8TtbOyR+2Hjh5bb1uZx7U84kkzaLVrivsvRU7FEMC/W+6Ae6Fv3f4v98i4Zn
Lw74MuMnMcY6q+srT9QjCqr7Ew7xp/G7fbkEGWi0zURua8of9U44c7MsktVPlXna
RNG/MudN3+oH28fMycKJzqR6tDSa4LCLBrLCBWt3PoLBZTF1N9zGZOdENnF4pzyt
ay+gO4x9U/niYCuLX0wwE5oKofP3TJ0MsRMGv1J4nzQYYUR5XBbIIqNC1JKcMr9I
H7DQpemUXFzPGXClgQfvAJzBpvFq5vlfVviVH4STuhq9oPN9HZ+bIH1xmOL2lLaR
t7et2DGBrY2rGSNmfGX2hItcEA6ojnubdthgMlrC0yijcYVDdq8y1oO3NhfQCu0C
feBN3oe+FepFKLjlw3YEnyBVbGsmGrXqybGzoVesqPeI9Jn0a/AvrXM/AuhWNeI1
13a01pxaffwsv+RwTgYpvQ3XIQwx5+5/+Pjcug2jqvAvhQ33ImgM2JI8VwgekMQj
wGBG25Rad1cuZBtcanFkWMcmykeC5zSw4ma0bStgsP29pQFxceLpeej6FYjG8Dkd
p4HKGawWMpURbAf790hClZMZdXJEMKEYmBJCy2DuYzMjTczH8Y0dBJ1kR3moyFcc
JU13ghztQMd31xOa+A2AR0hhgYcFYxzA/BlbhYrQungJoGfBGpMGr/N3/v3AnnIW
wc34+8J6TAY1A13kb87t17oh/xxQvNexYrZzxsAx0vdqtEo3fZKqR7LL3XHGBcA3
jHBQ9zlUR4Ao88PpMtYwyo41Wb96kOrswJSGiSESrxBgy2Q2w25te5N8zXK8byk7
VeMJuNDy0pw67OarrfQ3TkGtDEIlkW3DgjfC5HMyc1BRAF2Y501jV1s2yVQ0kiMT
SnQXKMP/0Zz3p2GmA+3rCKcdsYnQeMZArDqhAfeI8UOC6ZNDoTHrD7jSGrqqldOX
rNrbnqwcjChL2w6BwP2EgrGf1bS7sqhhRssFvneWEaWdesWUBoLg6oQNpNy5j0KE
IewTOgYanneynP3fquGxRNfYIGkdFTZt2yXFUC4YMHRUDkb2q0oI1jo75W92AIFa
cG/LQEQL9LWRFskPAk+9E0qwvgxh4h0zQxuoFrCMC2Cm3M/SReNzCG3Yc4CTgXIw
QtcZLLLICAvHgVZDAApqgZ8s8qDfz5fkJMdmt8jGQV/nEeeUCkvDucsZEJT4qLvM
YsPabMOxXcvL03/3s/9hcn0MYNYKcODcwMUSwOchY+xXq0avX+WotvbC98HMv+0V
4TpCGgQ+7KOOO8kplY0qLOQDYBBvgKqvevH34zqDdaYtZ42HGWycMszx0TdJaqRn
9V1+awZJoq926PxXjghMsEMiSXJdy0RDuJPMTBpDI5I2FVF6FKa/LlQ/mPSOSdPF
Rjn3byahqA+gVkpS92SqBTXfgxu9wArMngMhwE0x644HnzZzvqMud2z1IYYIAlG7
GKdsZnZ0uHwMVe61AOr7C3dtp9bxmvew/xmEjcaJWGexlcPuV2txK6NgvhZty+Q7
A9/vr++xV8e9And+V+tZULuFSvtsIgVJ130gQAriiAwNSh7E8MTgKhm8fqekYr7g
AmKhBDgzJ+4qVZAEdDU/uS048Oi5sKAhLaQLV7MGyZnUMs3cNkMS/1MwYnLlJMAS
FyQxrMVuQLcZwh+1RWWeMmcrYQF3uIBRdEl0j+kQaG3zp6B7FetBH91OOJs3sVYh
evjyapEJBpyUECs4zjYWMQkqTU3gH+ZoehMEK2f2nfJTB/8FtUX55LwVNFu41oqA
UtnkxrdAAbp3qwns9nlkFk8haTzYxHLYdSJar0CMjXbD8L4xzSP1W7jRPUH13++Y
doLvgWYzKlaHnAKqeNWaXXIigxVWczMyxfu8diJoO37E5tgx9t/nYAB+YMcyqc5B
TdUsMsHq1cFXKPRIxhPI4cNW01qCFX9xucD8DPHUB/rE6nh6rKM8JSCrwC0NxpP5
0s7rL4E6dmMlkbd2+KTusD8M+Ls5DVrMyL1fG9r27FfnOAhmC2rBDUOQ0Uw9KuNN
0rCQYa3wU++anug9RWalG63+fJDuHZrcTYHjvoR0seK11jF8E1DF8QcQYNkK72tA
J1dY/f447G1FOwHdAtNo4q1bcMH+0mpr1llBePBI9Vr4Ei8THSdT0mhJTAm+ZGZw
Z8elX8qRZXf1umjDabvYsYr9MNNBKHjVXpkwCIHNyWH4QOtLJOQVMZ2GUUGlzzoj
FDC7T9NB3JA0EMWdJTiAa4sU88xyi7BDkG92bcdtdfLkxhH4PTKkakrfB4Hv+tnm
ReM0La3o00iPpb6IWGdAGPfyG3XlEPMHFG43oXF8qXSPPV0svSiaxnSwVWS1iGgO
1FZoN2n48PW/qlz0K+/ANlcziU8VHmGD8AGlag/7KCM7Uu9TJSHpetNtZFalGztT
/eOTssddUuIwiD76K+kVvuOrzAmuUEBF/O6dSk9scyTWZm7wFW/diOfQYaErO+sD
OAbQGtzGFGgtgevlYDU5PcvqgSC9+nlSrAsUXzqUYmo+J1/n/BeuqQFGVfYOv5aL
aEUOcTe6bfcoc9fJQQ7n/G/gQ1PbzDYkavzrX0QkqTSapT4SH86a6HH44Xmnc6QW
mIEG2izy+eYzlEPuNngrvIZjdVxA9jr5JnTNjOzhAW8rqf772ysEFYQWXSJCG8AY
CrUuRfNa4Yo5zJZlJu5VdrRANylexqcUOTS+nj4DhUtyQHCYTEgPxRgUi1IHLrhY
r6fO8mHoqHRUatshshz7U+B5/DgrOBRbkSm1GjhXtzORpcB0ntzHeOeWT86nxgVM
n8990wtvxvTC5EtEScG3BDtznYtMkDtKhMpcoojC2O2B2VgpCP2rCxruuTJS2VEE
LAIgE1cbROkndySRhMYg2hMd4scIKLpoHkoWuDB0HiVp9wrifVpPhuvfjWkEkip/
Wy1KbdImcp5prJAg8C3OjBybF0aCENxeUlJx0f/VnJa0d5VwU3ZNvUy17hsPhcu3
ieA2Iyvmjrrxi5A6om8oqDMCcFQg679O+S5ffvAsnJi/FDt1m0E/FCfPZWjHxvTP
UiLW/IN8o1cy8bNRrF31gv/BLfEhUxVTxOWQSI+2EMjpYLzLzT2id9fyiWaC2+/K
9R0zEtpFmXMzDUIi7wZKCUu3zgDMY8smUZ7w6FYIkMJs8nCJ0HMKMXBM0Qh0RDkh
fR1Ij5eObGD/I59DPGe/AhitNojlleyvevunHpn9Tp/Q9Qm9f7D3FKyf4mfxrTVk
5S5EXIaiyTTrIEaZ4ETsEfEgOX7n+kR/Et6pwzea7VwzOmbkg/6SCZQGo/wUrmPh
2bdq4nPGJ8U+uhUjv9es3gLEeArrKuM/TFKmZ4r4ACtkx3vDe2RzRBNFlndcQ0F3
6kuAhPduKmAT+4x8yLxYDIAt7KmJATASAu1CwSqJfVdzWygKUBY3CA8rvtwJq23V
Jwtoe1WbKpRpZz+oEld+ESaRttR2lNAPEH+4Fzum0gPiuK/L8+X6EvLXRaLn5G0k
wROoXnGYwm3ymNPiWtLwdMnZvYd/DSbPKreT2G0KAfdD0aIWsQoGk2uBBPgekgv2
gvuSx35xA/U+q2DFhnTia6lf1OMVKoZALucWaY8yfl3NEDxZ4SRyjqSSpnONwzxy
sDZLTvCX5MzjzjFR0bVyg77zTDN/HY33txNn5vXmrb05DL8TybceVDWPnJoUkKSh
GfZspmHzMcCIN/CI0Fzcj6nkkYXJOFKbj8mzByjTPHFktCH4cFcaIhQfJro4Z7Oi
ghnMpqFaDWsg7VRHZVhK1U5RbdFDUfThrOmIcYnoFZ+/xqffmWA52NbjrfnXfNsD
3WIbh/Vr5bsgE7dYJgn0/7XI4V5oGOfPkXOXc48xAznkUdURXL9iwDrL6o+AkMFl
zsX1MWHtfkHGZTwUiNU1JMAjNDXXuKwvBf+ZSaAH8WmsdFaAvuegqqxhyjYfPYrs
RK9vvmoU0YWBIwOzEKberLrbSjg8DAjLk4Y5iZE7cM62PVqkM+LWSujKjk+4KM5+
abRy1V+fHGrQ14e5fmQjMQNWwh/ZzLtMgttd0ny3TzYsDxBI/ULdAIOAStMjtZT0
wlXH5P4tUrVjCC5eMxv+6mFhYt+swu+iB3VfZUvqVeW/af71tOQjH2JEgz+aKhbD
FncYWGhg90Z8MtezoajfbHr4ASV9Pi9es1z0Gag2kNI+T2SvJ5Tw/KUcKjqKRr5b
B24QtPT+PAecVtPVlVEv6ur0XurDyl1pk3eeIQ/HfuW29YFLtTniMP+4arone6Ch
DIeDdRzYG6j5jC+qCa7aQW9Lq34Tl2qcmLXUvNuwYPYUg0FtdE/MA0tRtnQpHsuD
i23Ed5YOOU+eMJjl7ivfd7kuOkD7dYoNDKtptePUVSvqJXBmx7WxgnRjALAeCSxI
MOvCfjYbU606E8cwFnrxnkhlxzF4GJmInnNhrCvWMcuCNXNnPnigAOEPF3Gstp3u
y/JzXXwJ5PCAliRs69iMCIrcExBo9hm1vZ6op1/NsUJyA9v9YvxYs6iy27RXwDXG
ih6tghoCY7Pb6R12ZfTCb4k89eaLFL8SFdSYJylTZ8mG47Nci//DLu97+ojr2UIU
BsAzoJ9EocC1adhLaJWyaIU5NRjg/OS2tLbJkhVn+LqG2Ij4ZGufee+wnbeBDYbM
XoyHHxYXAfIIWSdcp2AAPBlBVxeilc9xS0kaZZAhoaLjYAq6u3QlRl9AWc/tCtAC
sTyotSyVRLegUGSJfBdZc3l8ei6NK/vHhRxv7h5QN42NtuzUh/sMngyr/Bw8XJRt
+JWuP11r/MPiaxmkEBlVAt5aBNxxoL/71b81A1k871IhI8LqSzgyx7St8y8XnVSq
sQZEZJ7kFwa2vDrZeYpd3jGy3/qE+lBxB1zkTPLW0CfuobYD+DhgpQFLABjzuW8R
kkFFaZ3is43DNXSDFA5HaHe+HOF3sT9NcTIVIWsYRNZeUeMPLTYIuj1goJ0Mo/+S
v3hMBEQ5EQZI/jcxM+7Y6CzaVKxwu1j2MRA0DvjGqYI8Cfpb6IUQH0xKDhS6AP8M
xVrwhhAUO1Wy3ERTVY+b/zXig4Cmyg+tKjg/az5Mspms1esWo7p0LlaYm+nkT89L
s1jyRWIt/soFFtGYJPnAAMxPuRwn+Su3WKUCJHDHRsSozlHomTUJVGUO2AKZTNzr
GLxga5S1V8IIkhSqrEKFjkh+4jRiKVbTwOqTDc6g4tK807+qOFzWN/ytDW9WcUtQ
hLNWDHNWmoo//3m5507s8sDwEVMX2MJA/PJ0iKAjhDFhOWDUVPHvmxyK4Xbn3u6E
4ijBnuAH/eVmDFqwS8gJdgMOuXRiTg5RcnP13mL7CmtGr1W+W5dMuG+Zxa+WVpK3
d0Z2BdIjh+b50x+nLQkfqdhjvRlnhJ5JOx+p1o2x9Kf9CXhrUUsHEo6lBRfzTvUQ
TfQAbsmQyGLSwj5LUSMwFtUC2y1SI3E/DonsBcV+56HZeyUk27OGnT5Cmrx2tY24
hFh0EyktCpOqMClBAmjiwnTzRIN/0KsV+x5lcdYl2WfZ8YjArQTWpASgYcstnGAR
oPEF+K5mcDTnl9kHdZ3VFsq8lB4k9eguGpWquS7VhUzal+wiqmw/meQJXy68ilzb
daJmjaDbuRhElDxCcaqikI4G117XKS7GKmc/VlPnNhRC4R6BtDJRhVOgyFS1D7NZ
0ZhpPHnFl6PwuUpXKx1nBM18pUgV1TpT+U0hvCgC/0+W9miW8JyGfsgbgYGfM3tc
Elm8YcnMGZG6BS63ZVd57bBf2Olp/2nhHr9EVvhIXwgaZJ0vsMpD0WRtsolKAhKc
OCyGYsa/BEDP4a4DMOR5u6Pg8vRtqMvYulZQnla7OVEb22IbHimQQqHb27eoMM7B
Jh6zPKTYNFgGez7ml5TI7xk7GF83wZ7MgJxu+/WmL/9TkA2nKNrSIlZOIqEf88IZ
VOtE8Exs2LHrAqA8o5Y95HdVcPOyGnKm8lYSGpOB4Yh/CZZ7N07s2sWwXLQpZpyZ
/6j3b2cks/LDvxiz/kO4J/OlKXMjvUZb1qJyXR/2eplNqtq6mSxGYrNA8YNKa9FF
/A5hOrrb/0w3vCsPFoSkLlBKzOwAmQVOdrsMX3QSAGcFXhrjLFREpBT2Rj+j4pIQ
xOK2U/qDxxhkOH8xGwYWyQYdzZP9EaCXXVwEQ+rcWM2Ae3Ijbh4ibX+IX64x9pXh
sAj0ZZc8dp9sGwxJ0gi440BSeDCFy5bgQCOcWjSm+a75KPn+m51lXOR+VSTccopV
JUWVgxkzydgfLzIcSHFG6L4JLfdzNEfpYWrxgSqsTdiJGFaDuFP2IiOoqa7xdsIT
LvpWBUPKXF21eHZy7EwqwM3N/HDGeCq1bZHorWDMCkgYRYBfV71nqgePkIGgrUvd
qircNLW5EqKQZQEA7aXWZhYn5YOHkxPDmiedJt7MuEo6bcGYSqRf1lPUdPz8+2JL
5fVBoI9z/z0lyRTA4ID7Df74RQB7/vzlSc9H5yziDe94ew0c10mqY+RtAbe1KM8b
wIDoik4RcO+vZIhzLi5ioAv0vkFnS+XiTeGo07uPCT62VQn0U0UqQcfAeTjZI3eU
qPh9N9px3HjDGHPKoVz3LgtDR50p1tjUxIl9w0+r3VgdaWRN42L0I9EavzgkXi7F
WxF57ReIs9r+pmJtNutGitbau2ATjnemuixekp54gNLmHb9d861aGEzOJFYPQblS
9y8iWUAI3QPPsCQldgikw+zETTadCRSzgxcmFGI+ELhFD/JRBwzKJqC1zsFmJ/6k
XVnoRTXfijh5nd8E3o8ERTzBLhJHUfcy2yz0TKlEFLHTNe28eD9eUyXgaKUL7E/I
vD5W90YihSej0l1liz0zjn1H7ZKAjYp1c15zbE/+CXLc3SvzaNbuc5DvZlUmzokz
RLFxQpaTWvelzddrq0sH47dV5r4m1UWl8EAktskCTVEbSDVW3P3kSHhD6zIJWXx9
4jDzfXgcze6UVHVhIpVpIWfm3CD148usXAzkHOb+q8tz2cipO2fh14omvhkjQr11
NI9xlESEk4+e3DNKBp1S5ah5SCruvt6eBPIh0PdT9zXsv8bPjXPFB6cnAtE61y9J
B0e1OKWQCJ+cnHZ6pcYQtWxyFHO0UKymrfr9wLMtVCTnPoWPQMyw4lGiP0TXNr3w
zNK4TPnSN3HF6VG1Po7laYE5lAGplb5cNSvcB5l0AmrU4OoHCq0mLzWiHvVWJTQb
zIbEqGpcqij15VRj87WgrajRlihxe5TNuMFTrUSpBiwfCrX3gH7r+C4hkmO4Hnsy
kdHJJ6AIjPg6jiuSVAVSuZQTWsp7UeM6Adp6Xd4n/l4y61mAzJ55q3x/vODIKPRI
KphPTEkLIjce3dn6Zb/F3yB1C9n8Bn9NTZ60mltqQyPDFhRCAWV5YilW6/4lxTfi
8WvJkenH6UqnSeM+Y5fBT2WZ5zC8fFc3myWFoCq8CT9zhgg2hSnmFikPVLeBFHZd
0W5KogZzt3N5HERTeuumkX9PWR7MKQIoqoYW1wOOJQnz7lhKsjdjnjLUOEnijGsF
hJobIdEtBtaBKhkrpScPA56G5OvfeDtRRPZ2hDT7QErbHewm7A+8xe1yfTZ+smF+
HNbaLYd6acEFaqNQ9NnvdenCaP91ZYtafoutGDrvI7kCXSAZ401VkPs2/bQAmp8k
yuKQrsMdOLgfw15Muxc5eUdF0TeEtb5OuAiDvDCC/ateFOCWi3QN4sMFJiY4b/JB
ZjAPToBEghgz5bcCfGItwgOgs509+FUQJv0hoKnzzX/sigPTM2+Wl+P9Yw607m3n
urwETPF+A02tYegHVhJYnteWbw620w+NDycd5aJjsLjgIXhYBQXEI2OFlnuvgBKW
CG2qZioJjEYOVoaO8WRLtGmGGBkKEBJMiJ4xhtWPjPf46G3Cq8Ev7U5UZidRbGz7
fs/iawjn4bElZDC4DVer6a5B1UHAG3LrYidL27Dc0oKYIqATBY73eBRImJGLoVw5
Y4sRnUxsZh91EJtDvOcllZdJc7s+tUmzCn8Clugr9WwHy4YKSKrXk/QSYgnvKLo9
OMQGu6SUCtsvBLPedCJx6AX3jzfQG9cgDcVierWFBwO7StFHKCx/S5x+pQ+bW+vz
sOMhV4CaY+o3aV5sPl5pzqLhEg6VUwhm66FChDbgXmBKjcvSdkZ6CIulWFFIxmkf
S/UL7QL7seqcQt6d11djJGYSvwr+MOrUkaJPXywCCDIdOOKoFhj7S+bikQdJQ8VN
GpfN7ijCIFpuZNsRqXoklj6xGOSC4zC/gqAzd2W8cw7lX8gXQ99lf2iyV5PHKB6u
yJN3AhsvxzMlbwfAMPpXfEdvGE+4Abv+5osmyHojmz4wzyRQpPclqlZoh+pGLVwg
lwstzt/+aHui8p4nm3xj0y9uBWgApplk4804F1WBCrdOONMx2AWj6qQTGz51DGOu
SuMW10sVDzvCps0hLlfSb0EH590TBpEMaY5ZmEqxfzK3GVlQA28iyH0zuoc5oLqH
TMA2PGBisPl9TZOJvi+dFJzs0pcSid1FNM2lA3SccYgJAB5GyDp/heXjfW8NsL2D
8Tmg+WPDBWvntcqVwkOhKIU8YM8QVK0v1uuR1hpagzShzhjX3rHx5XqPrdQHIHTS
msWMpWGLJv5itawlSdB2fxy8nx74SJMVoconz5v+QX7jl19k3ASURCS1uQSgXZ1J
lD12QKQxd2aszdg+GpUbfpcYjYML7TC/5XXCHniui7Tjh0/ija1T/F/cMwnFZ69e
d3cZDfBfGShT2ks8gWukv0bsef3cLn0CZbuvjwOW7XLyxXmEabIEkBNSA7UBSVPO
KKZoJXO96GQ5MdEJHbCQ1QaXkAlSeMJKxOIKd8s+hm5L2iGm2FHS44npFEgNE8VI
NDkt6EHM1Snjso/VbnANUbsszByVJfIWKCMUDhYWnvH2QBsmmilBvyE++82jHhKe
TU9xYzSuqOkCqDq+YtoYzldEb0idhWiDMJEF/SEZGLbHCL03EMYLblpyMTA+qiKW
tTByS7UZExxv5R7HZx4JL3kszxRwTtq5MpSHFpnDz2E6O7WsyP66PeviBJyFXOza
THL7i8zXjIlosgEaMeDwZVRKSWawR13yHuQQzd/RnCA8m4WQVqZa27kNQfzNA/iB
2Ose/JlnkvyE6AO/8zdX4C/kVPTzLVJhD3nruCPClPAqzs2hevUQCNkz0QCs7jui
eH1MaSdLzHOvuvjyNS7/7cqvZ54Ioh8NeSyAxjQqTWU7mnxfrBzk104PNjVhOIIA
az/5CBxDQL8F8AcL8u3zExjF/d059tAYtQiBDGNsFzaF+OS1g1HTiNqwD5i/k00B
HEiNro6iNqJVXHCDHL6RaV9nF6pRSBQGSwatO84LhpnjBbWKFtOCvYVpIqECfuPT
gPqK/fRLticfEordmbKe6le74T7LbPc1cxXU/udY+OO0RW0zYy4uFNuKSxhT/cRD
3akWWaCJpzCXDGdg1zwYMPwi+/pbXhBDg4gwqW0IsiS84x8j4SyHtUUXDDMnFzqP
SOGGWIygrsRTqc+Xd9iHRABkwyNCkGG4h3ArpLv9bdEf8KDEZBRvizIjbQfzKS8q
lkkT6fw+x5W9qtwJNvSxSB8ue2Nzr7bvaRswXK3aek7BmhTmKZh0BNfz5TYi58BX
FPBXc7x/f381UovWRmL7HrKG9IeovKSe4g1k3730UMjOzH94+YvrFmEfN5w0wuYJ
etyhkXrk6t+gdOYWJgPpZmMUrA8mxgp5AlrE2bRhg6+FxwQXOFopp6gYHIUQoIKp
9i27I8J17qNOITHU93ObsuMDZpbtpO1RCTuz1gGZuvkcssrdOuNVmq1LxDqlN3N4
MtD/Sr0wUVrIIcDPk2/6cZDbYpZFgYwsomg4qnKOhKaAfiQFoQngQS9GCe0pEZSa
p2CF4Rm4AZ2JVv7gRs0kx+Oit8Z/tbUXg+OKQk0ZyFbu45UcgTMdrdp5NGPbyPlE
QZjfsO627nWeNGJJHv4WWVq4oFy/K0hqeER+qSKoc8xaa2VRj5zVI474JgAFrkRn
gqumsSB5WT+9ttTDp4YRA0EWHqhOtrNurtnXuo7rVwnibKPWpIUYwskbnOSTeWUy
fkm169LomeUXXUWEXeG+rtxZKjnZrEHUMwYzEPf/nnfjxhguJPLTGKCaWuy284iX
m7+oPsLPxX+AF7ZKIUc94ztgraM65CqkZFGQk9AXnUGmJFXvK5k9AqUHI4DPiXCZ
MmCo9TRu/jteWLW0SfnmYxHi94hRv5pCA2JecY+xHqDYSdASmx6BpljxB9Sn2669
uGqtLCcQjbqnae81KXQmWimF1tyWPq3/28ywo4JNBzDypixJSMgNRFjQErqvWQ2Z
pe8jkyofgtoHfJ+h1BgsFT06B1la9YhCSRkehvbXVCpBBiisbBHLtyCw6OzvxrWH
Kk8h11lekEewQWWLd/x9xe8nlX/2ihgrxWsnNuZjrPDKVqnc5V7L13Vqveh6tJ9d
i9GecPYMscm7shC0azSn79m30fGcrXTZKFlVojb0B6RyXSG9yCy9RZWV5HPQCIM7
WweCJbN9hCZJJBkseZ2Tt/G9o1VNXK0TSlqz2GC8daGSsMRcXciRJPKFP6j9OaAT
/l7/NhNf0RJMJqqGOfFm66v0DMXbYR4CToY/7HQI3EPwTqnD7AxWs4cU3bmXx0KL
AxgymasNHJpWlTFZAz7Xjt/BP8EHuo9DmVDO8H7uoZgN1zrVaNDX5ULJRrFWKfX5
xQ6JfYHMuqkg+XADyUnpBmaNu7dpRlbrkIcfDGIyshRvDMEgN8lhxfoBNQG9ggcd
tKaklSNSfqIZ49LnD9eqt+a5Jx3EmKH2BxOS2nfcFXshzTr7V9n03xpCRA/EEEMy
yRKKAtIofE8wZNiv6y7F+aYpCXIdgbAzZ7o2EaEXEOGmxcQC2r4TWxqHBgb0xNwQ
3s4Mo0b240hfedtdnfnuz7cVMDakq4SNlBACCWRrcu24SzGvf6pfUj7eV/PbivNf
qbEMVeqvIDiJ7EK9cgz3VlsnSz7nim21NpG6tGrlwEAFoFBqC+SKLMEZ4sSKP34b
JH47NS22wsfetuYfc5cSdaUIjWh1I5AF+oUQSLN0RFAI1WmI9VouBNcnpjutfURv
EANLCVXqAUk+aLunkhstcbW9wa5LzU9fLVdEmwZPN8GQq4RJynPgwKPgx5QU+5vc
1XsF9/7zcbNYu8KzMl4FqE/xgf+L51VbLU0988NpNk96phKUgaE5HNSmMHMUFwAi
ZsVsyD31WPljv1SDjEpG/+qJi1ZYs64Crai3Mdhac2uMTE3dnSkOtzfQzWtF/SZD
Hz4PoeGRPJ1hZoQP2eyMAWQsEDFRpAbUh7REn1qe9rMhKLL0MDjw73VlwJTaMYX5
WuIIQZNoRMSrSs/vJFgQ3cHSHNLfTHB2svuuF4Z0CoFrwvQ6BO3iCk7BH7lm8HMT
WBH3MkR7e7L6BPgiyFbCuv1XlQJ3tVROuxVzNUaGxjsYsXmhsGHV/Ariy9R3cTsF
QpsO2FoYUoVN/YFoCzWJLn8mAhNOFoNRuKULeDuWHJZYF4FmW1z19w2D91E7Wa+F
sGK4SCJ67rru9IwPQfDOJbncyIvSP9QBvUVcT5BxumJVAAUlPPPU5PcCXFXAZ0NC
LZwHf23byqJO8Go0csUA0FWr85TxU6H3EJYNL4a4k4aUq4PtLih+5H5T8MLb/Tk7
WVPIJCrvq10UmdfKfbYbBbFQqx9yzrJwnFbrDFK2cA3+fJCMRGRCS3oWtfeoU28E
Gxu5fSF2TOMKCkRe5MRkH7HVQvsdCUjVn2bK/B0AMBLT8UThTKfe2v0ZUnmLHuwj
h4gM72bKssbVRfHAs6CH4IQL9QS/kPVFpt+DRzD9CUXvkgtQb6IHbR4FqkVDEdSL
/DA4DaNq/Fxiv8cV7+j7I6COFfCLwFdgyZbmZGstzCZbBqd7aU6XfMdIrPgsaVqa
gdsluI2nfQgc2pZOkfIg+Ez+aCCmKnbHTR/GsWIt5qaCZkq6ob1hgMsPmOwVh1Cd
fZs8L+dF822OljjY9U57P6kHY1Dbj2NFMzHtmKj0NceMh4oDTk2pCJxxropWfd8c
V/CwopowmcyjkL0FEVumZomj/5kUQc+11Up7x6MCS8Zy+JH89thDG/N6HZWWtdkV
Mho3fK2Xb/VrI1bwWGVIOxo1VP0PexRqulGnM2w6QXJjsDGPNDPJYC4R43oxuTwJ
adFp9NkPH+Ome34YI8yI1jISosXxHuIp9dd15/gZAGYS0ISwOGOjF8zMpdFja7PE
Iax+Y0pnN+BFYDAq72TceM7D1zncNHeVwluuVFWNn8di2ZKwuT2HP0hGknghPq8z
7tuHVHq8XdRO2Dr0JxL6KxBuExoKgdOzEeDjjNkzolxjKc3rPyM7vSrqppaA3VT6
4oyZ2X1cax5wH8YSINLkG7A+a5AmIz5WhC5643if/HVZ5eekInVeBUxF9ZynbLBp
L2V3xZ5d/CWjbPzrL5JSxIzJCtXgXjPe3LSRmdGqSPScnmbx0iAioiY0OPhhn5Q/
3XKhjvMUNvmaPOQYASABrT8rv5WX/HiYEdnOUEAhRT0xTrcE+6MTak0U8CxIl48s
Ax4LzEMfeTaVh0r01RvmdLdcb9VD59cx3A14c8groqRiy4K8OxOaFZQcVgBZKh0r
2WOZQCOHmLp5GLrHEU8pKZ5ivIijTdAghRd06xb69oI8ViqLcOAy7JvfPRYIFUct
MUzmP4j3v9zIq4qLYHKHEARhNkuu5hxS1Gu10YRKjFa6Tx5DNuPBI5pB0TDWsllx
OqbbAx1h8va6xjCusQ6SV3Rh82LjVg5KHEe/GFAPv08VT4MTos/coabbRNOx6UNL
yJFf3uJdbWqKVX9AjeBLeMyxO2t0VP6tq6RfgjYmseFfyInCRuTp39AB3WU78AMK
EgcGiHcv7YQu/pg8rMq7Im9mOWmGQ6J0sEDb5ifaGV3oREmXKgnar9BQ+em30Jxh
79cz37JRQFzoVKXofgQSPjdLRorh2h+jzK4kxrsDMM3nXgffb8oDz34+9LzSe315
hOV4/LN551Dvvfxw0bGMqwoYKZ9xRqqo8Flr7+WCMXaFh2fFrOMIUMQMyfmQ3oqk
HIDXMdTMQ5Dpdb16gDK2W8eHhTnEFQJaHwdayfCY+nNweOCfUcA4H5w3aBUPmYLS
8hb0Es8hhy1PkxwyL42bmm+4R+0UshLNxa7ORSR2rYz9jM3RV/6EbFI8sTfNKdyn
mPoCCeFka/gCJO/re+v7JXJOc9P4oOw8k6BnhmZhihv4PXP191lQp+1y/ZjsfaU5
kt841TbS4HLSP39835Ta6G+tW+xRtUyMHV2NT0Zxl3wO10Q+/B2KUpF01GFSqohY
kk2c+3qrxcBcAr6HP0qWMUphcl9vRhwmngS48eUXfwVyRxtKA+/Eu/8QsACukwqs
tpCbIy1lk0wxoO6Dg1sQHFn28YhACJ1LuZjsMNLwDz1e/uOrYxXB+XHeUl4O+K+J
JAZbP2+g94ivopPJMnI09uyMv0G+du02bGVnMrP6igRxU6WArrn1ZAszA9St9SST
qz3pLAjHZavXq8BD+yrA57ry+nD037j+tdalvoJeFbrnc2t4y7Rs1HQUBpC+wo/Z
/tQ2rNmziKht0gziK7aJfKWokV36g5yKk5P4kxbJ3DeIXvlv6L9GdmxzSTE+TdtE
dmRTmve7B61DZBfoQCv+ze9yYJH64CFLxI2rYRuAOn+6gB58iw7BgloX79JbjFiP
7VQyOTmE//sseZ3tXNoD3JCyvTsfc4n7yK6SNsvGPU6mt1QzivnLsQvZZ/BRvbZ3
z0uNvePLz1FlbAQCLZnnN9+4jvPV3FSSld8OyMFN4b7bWK+yiPbjcjUMt+wqijZ7
q7nbbAnQqEDEo3O3IYJLFbbkolxu5vpyk8jhsaRaP1UQFl2JgByVAdy7mBY6xXc7
CJgDcM9Ke6x+o5vGjYu31cmRax5qgEz4mBZVy57utTk4mHNUfZla5fHe940cONNG
K52s6DDxwDxNLwD+WwIOSSW15I1hWsjJqpCuuQW0jHOpT9ctr3AxWg9WftaXMmwV
hEO+j0YBqe3fqwsn7bezhJV+Q8J6zh9UWivqjuGIsyjyl+s6cOrafqsnDWkW1yip
8k5ixupMZkL1PDI9d4qXmonGEU3lNaYnEK9cyAOnExYZzYRQJSPuSDxQ2K2YhX/m
/I4H6XBLV/ZkaIwHkfxjB3+ZDWRMS/1qoBfOyX6e2/9AvDzMIsCzWcdOzHa6vPJo
BxI0YL5P/4eK1RAZzAJGPbeMcKR31Hu25O7N3XvfoqJmOKJUd24QKJwHi3puOjSn
/t1bfYKbPJ38htjck1VRbl+M0uprp9qHl087UFaf7PDLrh70tIncJvVsFPs35sTT
Mp21lU/UDqqyg0bZpTJIB3qlRJoQxmt8lyxFk6rGcMbK5h1QySSSziga1gR6MPqq
LBdNXbPC7zS3upf9yzI/luPbSbgWfzvU5w2DGGQUmu/pL1QQSVnqFx1smgAtFDVc
3m0hWIM2B8qdlSqMdP/CW2EUS+kSqp2H4slnAxD7NGofQHLRpwBRY0zhQULSuPZQ
aNiaO4TRdrZlIn/A8POAsP01N9PEq6l3RQb0StxE0D33TWrITNqaOsTvYGc77cXE
ku889FPZXxwolRQ5Rd8buHZ450DUZwWvjlr6ah09oClj0zQVGYsMuGURFaRa5Y0r
2uxsBtTK4tYJbmbN1dQG2cf2XhuN4KJh4kE++rax+Rck3Zo0UOJk7esMJteOSDWX
Gt/6/JuInHG4XL1k/cNF89tKO918tx2XjVmWeBcy8aKGP7jFSMDXdK5/inAZwsvQ
WVtN0rFGsr9EOGUxIFSGqxx6XjL+al7AtEhRBLnpDNIeJhw5Zh6LgwRnPZ8yEzNX
xn2mXgLYhr5dEKqxVB9p11hBH3QF9fVmrhY2Um7UvZjNfesNgmjc3+nIirn1S5dc
P9JvivYhvKxF4vyeWcVFwb5BwsvEA1Pgdl/fx9omsYk48TV/ey6ZKZ/3rNCtt9d/
9t30mQoFLc5tZQlicXsLzdGYR5uCz4zgZ+zWTJHKhWitOhpS73qWTWBCPpWO+Wtj
jSgllUcjbOD9IY/FUGIHLog7f8Kj5Wj8a46kVGWD5xzdyLo7HxEgjPomuLQm/Pbf
1ttsgLD2RmrtTp2vo7VbBKqowL5hnvPFMNQcaiW6xdwHncWhtKHYAJVREq7/E/Xy
7EvPVilDmLery5TjwtNGRo/dULb8Ljotx0VRtYWol5O+cp7m2EpKgzVFu5df3LP0
d3Ct9R8SVYZUYurhzX0syeGGgeuKbXgYrbP2EaxE5IazRhcOXYlbGXPRX881Q1ok
NkQ79o/PANV+fF6LQy6o5H57FvhIav4IYgD9aqrnsywHt3JxQGchbEPg9/An1Uij
qepKPHt31RLvDtPAMTCNHYVM9Wq+cN+gZv8zRLa3d/3LUDo+6v8qUr18lZj8UiLM
7GMqnbmN3cHOHPli0scfhDko4RcFpU+h2k2weRKyFVgJgye8gxj9WtnpW9X/mULf
6CabC2yfUYBQNyGNr53jB/+bGVR1bdXjLsYIqlxfZfSRh5CXEn6aFXAV4CBxAAQx
9t/OPdPe7M+LKyQeOFeyaagHJeC9slVDHBAnCdUcbIMuzc0iUhKNhdVQiH2voMpv
1GogXQswI28p73AdLzamxkycZ8HCm8eLvsSsnYJZmr6gA5vuawL5JPB5eRT+HGWY
T3pv2E+/4AXOUpD0X8SC6UE3hQnvQBz2R5cVYeVR0Q9/6G9EZzOlKn8j6wUZgkvb
EHdWIu72gsfb8IDti4MD9JtfkcSFLv8RHbaLYDiz3kVX70JDZ1k8f6y9vEp12Yc+
/nIUOyiCcRYgHIZQgCLghsQFE7DK60hdFlWB9pePUecMq1w2gPuYloTlZ0lbCs0Q
xQsnUw0K7MuftvMMJNXIWfwJd5GeKVK20sH9OjbbWJqXO9C25Oe/fgwYGW6eoUxE
tWOYpRT4HPd7rQ+w+yrmYz38da1O2GdDXVqPFqacUB3FGDne68eQEGjvthZSnGjA
r6HOpgoX5i/jOX7YV5rpqoCgCPRwrv4Bf81egoIjET+cE5mxq9uzpLEaZipENQPD
dpZgdSBOmoKxuHYtpuR/qjOHUrhnziKyTnV1+69CdYEKsJO5eWjmzYkN/lTl4sJL
LckxyArdGsbXPLJeV4d7vwO4/fUsUPuj9F+4NVOTt/g4AZzEHaFOvAK51cK+cnVX
Z+IioTPqPoW9ygGs+LyJJdNnNNNFsEB9UO1HUL3ucJuMmJ6NVHnVDSTaoBSHX/px
65DvYuE9TjxlJcqT3whaPxnef2ALD82vOXT10ckBxLcCGfXKJF431sAtuOwYLqBX
sqevmlD0Pa+JdfhysWJVNq83C1XbjhO/q0taW9wZ7hVL9sRN33IACCNZAFyIKK2n
3HNPsI/o2t0pIKfmDVeXh3B2/Uwu7kr2rWdOaAiWVTAsnfgYiBe0iYHjnGQEO4mi
5bdxsj/k8BwtQiE23f+RWXW7132A2PJiPm2DZfD4r9Y3u2sLaA0LRpG8O1dI2FzV
Q8VRaDMRtPlj/Pg75n1RT+yGkMhKXsR1sbbeD5lS129Z+ejPFGv0ces6JF4u2z9K
HUQ/o+RDILyPGNEViZLZ8QMsZ+j2UQp1rGDJwBh93p7Jk7e2k1KGuo4M54GOeWia
Pfw1N8scWeGc8VXBgg5wfn/cFSCmOtyc1TAVM1zhmmZowA8Afqm6/jc51Aj5ebQo
geTcjA+iLFsf69ptLZ5T+nF0TsV9s9ErRekraNc9aAJnLBJhinm5050PKzNJ2gyr
lsXU0OttKTAjGgUSChz9/Cc60J06SKFLmXjGlNkEp0iXn4cI8mQRKW9eIwq7tjjH
rLt4RJf0K7THnxShtODU11peVVGtTuMwO/FDBV2V2TUEhRWqd/DL+AZJaj7QK+ap
fscqHZlxpyGYquZr+oY6OUQZ+i4MJqtDS5wRgKyqPHeyehvK9wkkwoySZGByfnj8
0ZSsMmm8eJzzPJG1VB7ty/XqBSW7IYqhDxuAguGgnpRAGvIdd1V3FoswzPmsZn7w
en/hnvDvhakjqPSTbVoyZwvm0ELFcM03ycVjMec3eXQI0UW22D5ptEURWAP4qoJS
Hm0ycmJDXaBGbk9AXVIjLZlqsKlRGV3e3YNqGg2k5BtxhLdzzUW3UNyKcAhXdOra
cIcKLkFvPaOklepa9j6kE3XIBNgDUOBDhAbStRyfO67+w33fcAgutb7cYehuFfZs
PACuVDMRUMPtKuaEuty3O7Hc9yBxdOem5P4cAFC3Ca83r5MXlgJ3S/KUh2IlSYTi
XydvOP+mULiVk0vmTbyV5Xt52nh1i3IJIA3GwIuDg5Z3THmyvugV9qpawnGatI/I
n7WyJg/Q5HEhebpICJg7YYcd5zKYXGm5Wlw3uTVLoc+PlrXWhLoB5QRoddJ67w6h
FflSJzbZXQkSLkT6HhFKraOaQ0n4cuDqdt+i8C1Y9UWBIiA6A1VsArqZZOHCxiuF
26YMH+AFF4glfXJ+R4YVDMGGeuVJMe7zeoLvCUBwk2h9cFMQtOrj50xWw55s7U93
sRGCbsFV541wZcLS3j8NgjXYPtXqG0TWZhhxKuNjIE0Qx6b/iN8gOe5ebRkVzPzT
gRI0w3mc7OBWrmiZlEU61ADoE9X136ZzFHtbICZ5FtbxcffH4gSkGQlzbff63M/k
SlJeiIRl0fq7iAQ9vA9wanTlmwFu3Pd2u99D3RV/x9bjbNZsDsjKooKDGS6F5hZl
cZ0nNPhh5xkQn5yBacQ5GAr186f2/qsl84FXj9EUqYsnhOjryaSURH/XATMkroS5
O1oBP+3GuMYrwYy+Vq0QIfw1cuiaNaV2ymM1ePOPRarQjcOTQMrph84PkJ/5ykag
Ojkn7kebn2xYbKekJdPeZ1MJVpeRHLzBRScka+H2u1aPtSY/QCQ+i1GJvu0s6lF9
INWsI/dK57lgbXctbivtQYoWqQhoCdTfPpDG25G8RTQq5JVoykm8EJuYVLIsQwJo
3sNRoL5KimKrYy7WsedQSURYzcTWT2iCEa9wIO6tX0NOEkJ4DosBNrwOD+HPcNCg
EO18kHDTP+ZgMlj6icfe3pdf9aE8LNGv1G6bS6uw7T6kKFcEv/DmZsjlTuRm/JL9
jvUwTH1jGsIsKcoQUuB6306d0rQtAZMi8llQl3wCsBP0mo4SdGf4mKJbVJ0SR+hm
q+FWQRG/IiKL7hTUMIlqhHLC3HLyDY0g7gMrEPVm0NOkWrOXh7/v342wAt8FZj8T
96F32xnwTb4FJJmzb3eokND3y/pl+Bk+7FH/0X478u+45WbZHz3nY8/xlhiwmv8I
aTWrxFBcnKn/oupJyVUtNqCIczwV962lGWGdjuuEqupC25GG0Dfi5lnF9hlsTkfW
0gepTC/S95F8DKbdqrIrlHPQE6PxucW05Yxygmg1eKDJRDEmA82pzZkoMEUfMlLV
EWNd3F/FYlBcg6Iqy3qgRnON+gs8N3wkUxKtIP898C8Bc4SV9ymKDmuzEKaRRdT8
rgZZi2WnX0irfWG3Sa4TKJHyFlzs0+HWVoabLD4S68f4WqkcmIqKAM7JFD5p/8rt
qnGdzgVn3e3PvMOMR85YHvVDFdFt/xAI25sAIMp+w8FtBti5HpM/jK3GdATF+hwL
Wu6eAYw0ZYa9JohCTdhMpKGoJfAbWyvG61QijUFj24bybrgTM/ozC91xNxZL2Nuy
te3XQ/ZojnYv/dGVkgx6de9N+2d40Yiwcx+rSuJBzgwO6UapJKYmn0MuH4tnGzdb
Y8c2/4nv2cj5RwTItCisulmzujsbCc5AiXCyKaxo1S/KVdh2yAGVOnr6j6ii2oB0
0ZM6qU2yybODpy13gg5rpBBIlG2IAhJOExmBOkuoH10C1CGB80tCOKk0tjD+dR5I
ZtQ55EZMvYFW0TTGwi3ku+QuCaqcIeZZSorOzBq8eZ6uhqdDmpIdIeVwP6aOtEqC
3T0mpivIm5B97QTeB7yYpoo5W01hxxRHo5x4EYNOW1MMDbKBwBn3GlKskNR0UDLO
KjXbKn300b06ziqAIk4GuaCAbpmKL3c99zMZJYIwxQpwEth1dyB6JLwYpjXXgPWf
j/5j1FqGnDOebJA2KlbF01aaW4QtWCotKFGSWjPlEBhfcc1dlHmnzlXgYPzp4UZ/
Ev4LvpwtT5eEMIi2jTeLI1UvOW+/lEOvpKeIAjUWAeS7H8PD+Kp8TBWyAzVhkJMa
um/kL/fAgJe+kbXhqAUGz+6bqYbZfW8puxK0UB6Hi2GAwVACxmlg9OoZQPO8IjGQ
Dp+ii+a2VsnkPVQ874mOnIYqCb9gfyaUt493u0UJBIs3LRvXxkjUOCXXOc0F9MZj
pOlygNWQT6//0kfbxC3CrIYJZe+GBKiu3+M7i3qE4NuHpmHFdtpMu6hnw08s2p/2
9tJF/XcXZw0K1T5Fg++xE4GqxwV6evb3kKJ5IE8OqR4vbV4FGJ5+G7ZxfUDzhKrQ
lCVOJflc82MWndNr8daGDVb9o+AytbQdfzwhPiJqXwmSHceSfVZiYQUHHeYsu+i7
bCD3e6HTf+0TR4VH4kZeiCFgnnKsub4ylspIaQMxxGy6BJ97d1ytK9Lo2iDolLFx
+Tb8wceAwQfDIGaqV7nVA5dW2lBhuH5FbDaeKyhV5sEtAgMKeVjlm1wuOU3zBH6j
oMIaGE96Y+G4FJEsqnOMm39fhUartkLwHpwIzv3o2GKWPkpUuBZcc36fa8SG9I1/
MOlCi3UJf8ewTJqvks2v9QL6jWnf2lcorCH9Vn3m36POL7GEi43XpghTbyVQrX/p
+3tTHXzwC+XB6bF3nhlko2fOdPuNOpD/qQlygdIBj/nhZ5RS/PA/RO9hXlylT3sO
EzkiBoj8Mn3pgf89sqQ3Fjo3+FSBy3zcLyGCsDuyfzoNWOh6e0p8rSZMvyZwGZwq
QW4FhMBIkOomis3lu4VlY5P5aDwu14dpbu3CCfvv0tJMDl8+/LFaqFOLjrI15pdd
0MhSfTaTAwg08hNapGiQ0NPxainy/W/aPpNAbN5ae4quZ5bpPtajfnJZK1lTCLO2
VPh/vajidlDQmJuDeBYEDZpwaxha7BBWDYW1N7y+St5mcwKhgOy5F0CI0YZpg+4c
WhcYWDB90w2T7x9d38NWm7QsgGuir+A7iX5BXSKFjecPflSejdZn6xLIsJBGNahc
10uqSlIXekCEWiOKSXKQLjlUspfjShZUwECorGdUemuU1QNfgDt7Gn4ueNyABYoN
3YaZ+bYw9J6itvpxr22sZehgiYrGRyV2gyxILdBa+MK8JZyX98izadWGmGb4beQm
UaYB3tX+4uu8QWrzM4jSwd+XX10V8xDfzKbjSK7pUmetKcJIcTr/mYzABux5zJTL
ZxAneCPmhg4+zPa6JvxSnwDmkydt+xhCQazeetlMImyzsc23a5AkNL6KQtNlqvSa
0N2ppqOxgkhpCnGZ2pz3FTAmN6OSMEDOsnYCoUbLRshTilJN0cZfEaQ68HIa0pLr
RDmVG7iE1x4XjD/D1LnhWaF3JQLbkIOC6tHAjzmuQkoEg5LiuZvUbZaQQEbhWNyW
/Yh0RAXtr2WFq0IiSIufiFvh25h7MVN0AgaOPa1wE2Jp4zSkWcC18cyTw+y32FZ5
POM6zQnhCtIUveDrM+TRlGEB6SgMlOtdnhgOeFfVnLGYBLknQKSnW9rrfnqx6YUZ
QChYOwtNwHLjx90Sdg/eD48YvIemOBHi9dGS0L0A+s8Iy0kOC4f54qTv4AtPtToZ
QEkaX2VsPHpUhcc/MGtUwOlPNiMtQTOyl9Dk3/lpz/4GNL3pu72+LDmTd76dtMHz
E2M52yFNeyH1M4UyXG/v/rYwbY04nrGCg05Z31F6ROUIWRhmLATJry7SzM6UMile
CIocEJn9WmU+1kUljCMiw6JiaH6re+FjcYNVE9/cKuuU+U848w5XN72N3rXy1aky
NqseoRjpYgH+jbtG2gf/XGNjeIyOyr1QZGrizUWBLA/3nOOdU/hyceL/4thDCz0c
xqwx2/BkbkqS8dI/U34CM2+tcycxAp3Djo5+Zi43nT7ZrJc9pkT6fj6C+LC8+92r
DoTUtQYfEsMqxc9nHVlniiJMqE1qUnK9J3MitGOY6hK4Seen8WaJTHMLDMvFm7Jr
8NnwVjEroT/WFXAlzgIsrAKJgXmevfT6lkdcibKwE2zJG7KG3c67x8pkMQr9zcS9
LvbkMxq7g+s5AsSgIvcqsZVyJ2YSbo8VzxNd8KvDRab58aNU4Sz7Ij2HCXkl2NBa
a6xGEz50i+Vc+FH0fAXUBLjxk93EK+T5g908phmX9lks+sM3yGq0B5K3CiGSbvXb
u9EEQ0Aogi6slgVCY8D71acCDhhJRsfcsD/sxgGS6FADyPGq2Sro/FYrAkxN4rSv
RZeQPf6WM+stm6LUyPDrb5VEGZiZMNe6nyLEi+7fdxImQ6Xdj1w0budAXFZc1yU3
YydCv/8M+PRLBA3GDvz+yz5L5sZ9TAxbpvXbiqLReP+8jueN3Zwvy2n0VlOFU1HP
sJbjfdTihUoNCVfmB81mvxlBw4DgJ5c+9vMiNeSlTgi0Pk+5/nXknvWhuD+diOXA
UQm8KXvC7NtdjNIo5aRNfuYtN1MnJ8kNnmShhohGOv0DTflwVv/ttDjh0KlArN2a
Splnh2pD2+eBLqv5hWTEHixRMcOnHrW4Eu8D7MhgAAvMcNfns2D8m3YoCO6OlggU
jFZpo/ZojsaMBszmH/Uj12n/hTm+UVOxqpu7MifN6noFS/TxfW3WtQEhd0vHh5lm
frO3thGjd80JvQdauBj1C4tDrUsR8yRUqWjSXwO32HttMtDMPuuREGnT+RHWAl0t
Rk8BRmn6RP5ACO7//bPHKBlxZpNL40p+LcjSv3knFGmTyRmlmCP4wDVcyAFWvd+P
HW1KbIM+fM/N5QHlQTZ3QK8i7rsD/zxyn/bYuQyzwfaizItYJpo7QSHUz9KhhgFV
NyCa5z1cRpSmMtSt5RrzbeWVMor9Ox7XwiSXHbjoOBfq60lTsfQPTMMoREHl615i
dwXUh0nft4dyONdhEfI+KoQkaZkiA74RwDumgGF5u3TNoOY9l7kNYMec8RkOJzI5
KZJZueCNDsD6jDLPHo4uAvWEJ8VIB4ySzAZBT6U5LGXr3bNBewdEt3N9nCysbvaS
E5QznWJb9xDu4G9bU6blxTW7zR+Ov1eq5WbpiBXU95gxlEY/NeJKFIXXqx3HB6Nh
mwv+tyPMKVOXFyDz7KIench28CA0lyiiEBCivEaIyMXI1fXkB5x5F6jWZFIhLTRa
fSOw+A9mli+2bhaVKApTT8aiE+TyerhnGBFxvm1CggyPmW1FXP48KyPOAJ5gcL1A
3yjxBGiWpuxeNGK+kLSTa2dNPuLpDmbRTodxpbDMhB2kWh1JddyKafxFchD0strj
ofLSYVNOE2+HMOduEpIWw62TMzd4ljec2IT036CI/dOST90y6Tw5F3WCLcvHAHAg
x8VjWZlSauHTbL2cK0j/00RHKFz92AOkgeLsmKvPv0u1EnBW6UTdCoxppDV3SKui
RnKNP8SWppEvjm6SBwmFK7+X0AahCadHSbWFLGfh6GOx4A0dYcjP6Z8ythM1TPej
oJ0W54JyFd6bcwajGMfW38JTlfgtaiDFfz/nBLE5DiIP/jPOyGRp41rpgKmiqNTI
sJOgEJ2fbDZ2FXeanYxABmCXEoKMFj6RcWqv2nrEFIuYfD8+8312xNAAz0jZLloy
ZiczCTUSf4ubPGdLkLGUaItXkAcz1vFi9GxrOalqywedxCFm5vVyvRIFjSmnQ+uX
v6qvTZrGpJ5SnG/LE33KXvt5UT7O90MMruPDReAdwkGkdpg/XwyQkqckm9YrRYs+
KpFEdZ8XRQly/2lUr2IAF5b8XAcibx6wijd7mor7bqmUrA7HGeIhenRnvDvcSESh
PTlc8zNae7wOer6fbV7XjFat+06mrxsi8FbeepYRUzqSsjlhlkNNV+CValxzrrW0
Ab+onATV+V5LZOhNh51QVCXIlN0Fjw7xzloIicc59e3TQ5PROsQY4NVyboYpyO6T
vmbCp03quxNuPicQpKJ8uwjjiTbmIgCeKiYoQymWDDrtAIbylEJCv/Yg5jBTdZrN
gVaKvFMUL+aadC97MGis07/Z+aG0ynxmEH/BOW+BMH6Ezf4ow2pUpnmIxi3tBzsY
Rw68wVngIpMe97Le3QAdIetfIcCnfx/R9tGFFWmtspjasLfFnlEN2z/KPm02NHF2
Egv4pOSX4+xBuLBurvgCSxJCLpNJkb3jT+lVE+23i9RyDx1aCVzlzctPnyOGb26p
eFDwtSR4kY/bd/KtZXemYTx+bNaXoQk7K+jEntflqnrEqfPMnuIjn0XX+fFJc5wu
MjszDyRKv1xtRP7r3sxSv4Qvldvsgpn7+b7iDIxcwAXL3zPI0Isugm6OIStpBYss
RY1J+fYyjcZzs58mnlEHAOF4xfbjHJTyKsFZ2kz7QZ8gAINkrfi4K6go3Sm5AQac
nFR9ODuf4S7dMQoMdYjS3dwibMjiZPIhVLgTP0+tEqh7gd2HBcn2kpYr3X3JKPG2
YX/0CowHzOSLhLVWPEr5UbWNTmtJLHk1uWiRbI+QmEnZ0f3zIxBR8eetg8MgRWXg
Zepspu9NPg3QyjKDP56MSWQVmyT/OYaZx6ZwaV9Xg1yTvQbYqASbqObTUrTQrQ4n
b17QXDhKAHTUBQ4sC3KXCdkRXxJfz6CkAXD4Qb0CH/KNwShbdMNRVHbGcIPQ/w7N
ayt+qkLC5hb3i59UDB3DFMjSiLW/ELB1TsUqHn3Ext9mm8toNLfzbrgtKvQ/3+Zb
YSIkieLKqZYZ1F9vG/WefHM6UUq+JPekc3B5BAbb8grlUDzoVC6FKCqmCxhrqJzE
/4pMFEOOtBViZWjKqtHCNZfFD+FeKVYSIZBG8p0UtU+ibbMJ9XhvrOOUn3zs6JLu
AnTM6Gy/xXh2xqx8DWZ6JhG8PdeHZvfvBlyOM8sONOO4RVI/KB033agMgAt8ckbD
wcWdKPFQPPQegrc8oElDoPY+3YB/Xko0kxhnJcSyVPj9fsQp2SznaonnSsMCQwwn
CbI+CwJ48lmsw5bw6xYRw5e2JAGf9iI/Mup592xu1LBkkcfMWC7bVxeuENUdihzu
BSBj40j3jDdwqfSw33JJIVP8FRsxa9pWTzGopGwI0xF656NiypS/Rg/f6mg3NltV
XetLJ+1NtYX/FoOr3cZWAmA6XRT0XDzYk9IPQfPAp4QKUjHPcCDrK+O9xj/u+rFW
TAWkb1YtfRzCzoQ+1xDPYPl2jTjFuIh0G/2rcem+tCjl+PWctWsdz/YhgMD1dBSM
luqbDzU6V2R9ZCKxGTrlFFB/qoosvGoFSCpU5OLQFBwJT8v2bkh1jZizSXAoMUDM
e2zidBkdAwSlKNgIE26vkPVcFTJCL20IOuD1Lfk8ynydSeoGpC3xCrYWGipdQ5qh
fvGoGvgflRFUbx20kiK1Eva3dJKolPiQZ6Oq+SZvXiStLbzXd1XyRGxbYGtIxbbP
Mt3+NeV8tIylDdB6c2GibGfedsv0Vmr9posAau2myA3Dba/zSj1UT8a6VM0W9K/L
2eN6Qvlsqyx8mOEC0IDHM3Yuuf6gs/QJ9dF6mJ8FW+WdKdx/2QIAjmx6/c5GKymT
pGNUWsMng2bLqfMZSxcCQZfkzbpkfw3X4ukIwzp2to3sCWXdUVid0njQsWGN520+
oLNIB9VnBesO0BJeoNBKr0Z0vK5kxJo/xzQNYqD97V5adCSyinGpqbV8FK7EwZoS
AnSI9+c/CoHAdzzc7VTp7BPMbxwbRFjqOfjyWWQ98Gnozg4fg9muEqNzo50pXyl7
ORsviEBYQxpsiEpLPSCSjRO3DlIeIdbnRdSLf9y13laPwPU6mF7E9/hoVgKOTlfa
1J1a/ayeu6uUMW+BrksM1cYqGLU6lsrN9RcUZlLLBUTjExY/glLvnrJ1MinO5dIo
MtCMC0Cw5mlV7eAXzbEK/BO6eq4z0yCmXhhkl0sIhTmWmxN5ZjKJiCtWi6197dTY
GGSM9jTwRlhaKra+0XBTgxguQvIOmAQrqWY0NYHI9AAg707KDTnNTOeTD85WCDtk
hvpKuT7S+GZ7Ka0zihIy8eDksjSG5GgmQwZkBpe/T0PU+7AuXjGXsgZ9KJZfvYP7
0pd/WVZ9VrrUUep5wcxnlOI313/otT8Btr+3KSagBL8EdRSV19l6l2vdm5joyiG4
TJxzPpVi+tfrJ90mfuxf7je+rbuffd/4LQRo9m64gEO0r8IrzCI5J2V86brub4QH
aoa/12FIqYuLNmieo3d4eo6smdwlgzsG95QdVpOfGe4nebf4cmmt6DW8DHFJY/Xw
5fvPpwtHfPkZrODk3cm1UeURICtODKdO1914ryJx/7epXn/GGWpM90HNeb1l1v2W
LwouvgxUidTHudrNSOApTaTObanTUEMgdH1QyYp3MatMAr1glxFIsT0w0xfSqAA1
tqv60iyViqzPRP0Nk6bPE8qdgsw4RMbTEi+gpWQabNQArdox0qnbv+Hw9h53btii
tMJEo9foJou/9Vv1ZZ4XbLUI6wAtW7PYJVCXjxg65cGXpHMUwcjfyZCrtWGqNho9
TpcX8K5EEYvmTc7mNY5EmOgIbEtNc9IjG1o5NcNOolLF2MnDwdnv/j6QvNiIHBW1
wbGcwAN5czFIsNd8BFTqtFA2TNVNnjO4OAzcEh+u9BMJ6PXqflw7uJ+lriPGfm6/
Z70y7lHFpj4eNeIRP7LGT/iHQW7tzTOxAtSm53BnfsXdmy5W6LV2vqWB4EvSHTlW
olJBrIdozar000YX5vWf+V3wUXnN82P62jJRjdvwfvJd7ITUXTnBZ+53s4VkRiW9
2mNn18SYFjC9zK213MKsN6eA1fRfPxq7tykUUTiejwKUs+ebKypW/A5GxjEMboy1
2O/2C/H+M2qWTsyZiXE3N11yaoiSu4C7h9LH4ekCVZ4hqW8dZJzOzMbaO0irVwgU
ZspxEPgu3n3xTQL3mWmYxK/zojoCkouJCxhT1AmW+FpK87dGHTmQyHs2ybu4zVDM
s6HZ8VSbh+/GtJ2KMiFVvILFiGatTDwPkbLpkbkpCDJC5e/kUFqFZiKqgY3wvK3p
8DojpUnUnHsK60alqgxcQprAzIyWlXoLnjgpbSGnRcO7QI12SInAat+YPPKo363T
4yb2UijHZ9pcRUKPDwuONso40lyxhlIfikK5ampEpvxqjStUUBOfTpvJgnjWZlP6
/GQVc9sho/eVj2t2XnK5PO9f0aomdVixaZqZt/3CMkow3mdnC0Y36tPogmMhtz75
ws0LZQYgFBbyA0AfSKHGnqAbCrZPtyzpKGxPrb9gQINHir3A93dWWtnci6RzfQqK
Fbdw2yMXsMemP3DSZuHsJtD4tsMNVAO5Cg0QgdgYiZe+xwvzxmGpcwilzyauW8Rh
b+bJ0uJwCbZCgbrm9l4uuR4Yt/xdmxbcJVJ4jMWCChOWNvy5uz9OoGXWKAXa6dxR
UxhEx3Zxh5H9WpN/fcWQh0asckJaI1tNkTzt0cz+vJHQr43YO/+mLQ0rl/r+RShX
Ce9P7B9kMaTRnJXE+vS4PAs71M4FI6QhtxzuzTqh0ylbnKFCChGiJG64nxRE9kfL
wqNVjHDt0KqIhPZ62w6Un1OFOliFCBaJjM88SPwLrwQdFqvIRM6QE8XpBv09qpdi
sD3mL2zGTix+Icp2ou8eTO3CY/ilnwObzFsDGGip9d+UAmz3yrtZg7dOD3mtQPkg
Vc+caJ13EL8IoB9HM4/llxElAu+l/YjJfm3jKrRkG93GCZOg3Mu92XAulqdewvzl
jt90P7IkC85aRLjnVqX35+A9ttzr4ceQ8gkPbWXUcVxmk7Ug85n+0IEMxf0YyCs6
qGQ9CpVmI+YRxoAkB/9h94+yDp2xn5mX04fjtHmUzTVPDpBEVIEt/VUaD54rpTl0
oCEMWasdpyoSDtpy1Q8NoL6+F8gpwcwZzEPdF4VADd9vLkZgJyKw/A9RD1thgaSm
vUFEtdGKfld4N32PDmVPY5Wb8mzf/AeTsbVcRlvC3UaSC4icWsLozskSNNZde0SY
p/WOu2Vs7NltXDT9pvoCjzPmsHAYcmi7xwDEQQrkVhTkeq68tQCGXI3HzZbK6QQb
70NJ86cnzxNz/4sbA8EuDcdwFNWZWqSfiYhCzvrFsdsCB5L9YBuPVRDmv/f/ICmm
1FkN7kpWrqh1RUtUngZE9oUFYC8aCpas+YBcZ1MsYQAMKcUJyDV1ClYychHSukOS
UYk+5M6PjMAMSu6A0HGBaCDFHtNE1KDQS08p7jxZAdDzILcq/QCXGpTwqTw8HcrW
rrsPp9qChhtyN9i1ybA5HtW+Nk4tJUIumLVo7cx+279ogfomAJaonbPinvEnNqpu
HzVyGbxgUf7s2eS/KhwKkzAkIwVSe0GxuR3YutwZuYSRDmKqbo5tYeSkVbioT5eX
pBh0NlopJgCB20hP5+0UvorTSeBC78zT0MSMp4oez3mA6vPehVikHwcDDuLuZXdY
C+dAZNywl4qDIFCQmAaKVEnK9dikAGtDijBqu1HFNVZvlCbyZ8DKGHfVhKdTDlIY
yQ5bYXpLIuIZv5To/ZUsgcbzbl3QJWLl/gnTOhLA4DjPqVSHfUVcIaxR5PKCY7ZX
w2srbvniXaU47QuZb2zZog0kj0YBTtAztRfddYlbkI0Cd41gYSxnsTCYB1vJ1Wqj
W24Rf47Bx2zI9dlFj5BtmP2X9SMubi9k2SYC3O7Rzg0T+ECfvqWJ2iDG0s9ooM35
8hFF6dlR4yj+5O+XkddcRKvAlEquVphnECWL5/LjcL2jT2tOsKa/ufDVd9pBkJ7F
Cd7i/lIsj76iMCYO6vLkZgFUubWdVjyTcsAamsLia/QiDVuVtzaIb7lRod7oLEtB
2b7n1CNUVh3VhTlhpGhf5Xg1hgoIEQc/60q5ip6LJ/PfkLAgYK02K51u31w5s2WA
vhmrEKvzBzse2Nbjk817vFY+e7WxxbTLVCy60O7fcPbP+tOWCuHE85EkwQMibtL0
uWOJPVMDhNva69UqWE9zivHv7x6kwKs1/9T43Mq/JzWzdfgPXbtxPXFIAfVOVcLx
NCPV+LDNg0MU3Wx52kAe+DXmJeRe5EGVHqRwRyAy6OYBQ/62jh6n2rRefwAnOZd2
VzLIhqtnEVy101/0A17uiF73Cgoe4JkkNYPuBTP25CITxfpjN5GA0hZUSpK3O+aF
3YDU4wByfdDy2CtJiKVAU5GMjk/fmhTssA0NjZrhaV8+K8t4/yCJUINHPQzLYxNN
zwJOyRwWVgvrtRJbHyTyTMWjtW73RGEYv4pCHSpcLuMg4Q6mwN4BJtZFKyx7j87y
F/rDHEwT4D/9EIqwmu4+H7fuctswOpxVVbOtb6bjLJXqZ47w4mgVyX24wQWWasz6
7Xx+XULBEtvbenNlc5taL5puspI01K5wFpNz10JRjsh79B3faa+fOvDCxq689gyH
kCc35Nj9A+jA/jJAZwo6wnis0I26dD1qkP6nslawmSZw/nIBidt/5x57QnaPbZlg
dsmvJ9eoy83h2UO1y3XZHeeSvJfm/2pJBHneohtWWOWruIYBJA5GFzNpxIESFblv
ZcMKH3AIdk+k6EyM3WL8+f+6x2/2M6KMAn12SygJh13yLsCAnDcBCaRq3ZvDqWZE
SdkW5U41uRXjtmMx2cqIKAyGwQFXeDDsIwy8pgch7bqlOSlOc1mJ3W6uN0fHemKK
NF8lXv0J3OJBLqx7g9uo+KO64mjupzn/Va4nzBbgfKeeQYb6Vc4Co6HFL9RJ40fc
LRNZxgLdITsye+FIxalvlsOzOb4aDGa4LM+ZS9n0RrG4qfCIDIqOiKejxAR9+o+s
l+X8g+xaq/uMeAaRAn6XnnWc+ru1qOAXIV9P58I6GM9UBsmcm3V2my9FUylntNJq
qN3WzVmEhonW0U/B86vZtYSEuvUQ1w5x1TnOJGS5tEzzvHtpGh2NtvXYzZOwCp3Q
UARt+Yal44Efe1H0SVS7UXktE3ZVxqT8eLTOyTcRNVBelopUUpZ7YKCqK9cZhjoV
bdeXRXtGXEKqo2sv29+ZzTLueZu8AP3iZKhhkMcKnMM2wqEfNXwxAH4Hze3e3f18
6fZhCjltz2ni5ltFQErnE+LR6BRG6XGBopyBKdewWiY1oMjNLLJqzkE0DpDbr8gT
NVU10LqfqvlxznSRssv0z1pD5D/DwCKBwtFkI3pLF3CVksrvxK3ilJGdg80sBgYM
JBnfOzLTDU6khCgHR1OScocDUqsMHVvXG590KoQb7ulTzhptH/MBcq+x36Y9RF56
7Y1PPCaidAV8Kzi43QquRqH11HQRG0v2PC6Z1bmEIrRI/cvrzIc6IzHOqEFJrUtw
4swSGilrUHxRjTMXVRwmsjjhSJcZ+2DdArHxHSdnJsDmlBZ5T2yUnbsJFs7ZCA39
GitOHp6LMG/qPdfzz0lojoQD5cZj9TUhMK4up5lzDEqbaQZk7F91zUijqw5rWT7U
wd5rLxr8mNHfahsyzNSgWcoBoJxAdNmdMiCiQZuGC6/iXEwWJc4DNc1X4o0G4vYw
E/YzV4XtODNXxequ0lkEzp7PrmYHNkW6j0YHyS4Xjtdsn5Ww8/uTZttiDjZ9M7/Z
aidAkDMDv9Z28cO5J8R8XAcWwOrhY+NZU7T4PzxFxTxykMD9vu71lCpNYlvaEkkc
MMbpS/oV8r2GvwFSDlnyXCSuzxOX6Oq8w9LN7OP0SkcSxEF4YpCF2e+ewYRnLQKn
VX2jrI/S38pSlzt2xy7wWyES7J7e1BogwbuCIv07yW7tMtp+9Ts7HIH9NUAbOwSN
HKBGF49ETXSKQsx7h+OjArLLe3TQdmX+SAKLA3Gz381kz5ks2o8eP+3kwXWD/SCZ
ORi75L4NKbBKFyjZg01F3rqDP6oftMO+bSHolqu805KuooKBuPD3nVvSaD8aXlSH
3q1TjT3gUn736Qio/an4Eqm6k0uxnRAZPqcHGSSMwICK1IIZmz23Islbv8aD1QhU
LvsN9CAL7lZXQ8cWkGZaz5o/D3KlBTVTT9Qyzu6L09GNOFh+EG4AczVShA3eFxbB
7hmP1yPOCZOmnnjSdlkzwfV+VVs5vuwFj5Jt29aH5kvsgA5h7wU1wm5wBhA1L5ua
+jZ3HLv6tGBWySdUWvYXB0+/amVa7jW+2QQT6q4EXWyA9PNFA6Q4dmeJSmIaDVJe
7+qr2elX2IU16PUtjW6GSfrDJhBlP0G30cOizbP368bzrAOds+FBm4TsP9rM/cLZ
+/R0r2XvU+vxg4rA/nYWV+OL0cbrnFMvFpiMAJz50k6Bg9LCdBYLD86k4ngveTTK
x0JFxkH344zxt6RrnWavo08Erg3YGCG6ANX6tYO0NPNbyrSRet+k9fyI3gk62joN
jpisr9PXPTF5EfSUkKyB4FwPzUOQSv0V4m2UZoPjF1C3cd8UNLmsgUDRqJ46abYx
vY8+ZiNodpCX8Axr9ogE5AS1Ackr6pA/+GsRTzwnOw1DlOtHqRuovOsFLUNIcGac
EbMR8QlW9VkeLzf8TQOpcDSBN7ScUccpvBprWLjV17ymclQBdplCme2bJBC4YBLk
XHRQJsJKlbpG3I5V/1wUCf2aza3TYOOlRpDiSkW4P9HOkU7QNBbl/wa85gXUHPnJ
rMOPILUYbg+KxbKO1yFpdkMn+LDtAsOVh8yOIYnSWRX4z6WniL661WOVXF0Cl8t/
I7NEputnTaCJg2tH0Ar1rKgyyXStftLjs8WsF24MND5eFEEabldZew4USucAkF16
+/gE+YxaELmG40NYJNRjTUMM/pEwvHHPC2g7EVCVFBLRspbY818djfJvLycmhBQE
PdFh5vxH7TyX4gZKB9Ya6vkj978oP2LqwveGPPywiw9xlP5cjemrDf1FJIdKRFUY
TUQvG3pFBxVKUdpsbm14jseW+jHGOb/ALg29iTP36SHJWFagYm6iX3SPY9byuZ2a
s9/ShBziMRDeLVD/A+ekmTPg4Dg4eqr7H/lCmpIZ4dwK/Z50vesmz8EA2n9vPupU
7HgweeMfF5WPP50scJODfsyXPPLfuR8qN4Vn5mNrSji+MdHI3hOK6WodCaW4uL31
oDPq6KNGcRQGmmNVyK5MAsqf+E/+v44BVT/w3IYh4mGNUyMKZGyWBOwOSnbEdLu9
kek+pwC2y9A08d1fwjWVkNerFqI4ouZbp1fmws/0VQYXsHqrYTUrqXij7aI0vp/a
HiR7I90WHLD2lsz1sOequwtFamJCxwCBYqYdtdmGGgcCQjJd184QdoGEh7cN7Ihl
UE/PLClTkclwwi+0GYdTkjTJS93ovUKiW0ifJBwGm9EIuEt/YFVR1kBhJWbop8ys
G9sW2xE4wsywdTC5DhzZzitneqKhX7HcDr/KlGeUkI3Z+VUvQla+U24LX2tPVY1g
vyDbxjnuo2lbO/MCBYGR6d9ZkF27cW/qTp5YOoTjFeh+Lj5MZLtjCrrQ7tiNUJ/9
flT2pdSBRAA2KPq4CZIvixJyB5vriiE7fydXVGICaOXdeVdBSEG4S49SiEbOu96P
iy8y6EI3r4mNnzuIhYEK2KU+co99ozkwF0NAnxZINXXJ6vyeMncYc1HHAIryM4Gt
NJKImAKFIkFQ1GJXYMh3u2ng8ezMjkBb2fVwG6lgYEvpJclleqq7zDqQu7fH1mI1
hG6QHrBWoR3FiWVN3+D54jLEZ7LsNH+FXl1fL1h45CokH8diIlxTJr5VkYeSnLZ0
msFEEoC9x8XvOa4gNZDiyFfeyXW09Wq01v2+3lGiONqMokDs5RqPFfrUUw/F1Rfd
dABwk81ShvTGQ1mEpY34vKUndME5N3WNw7BN68GElrB0QjwKqCiH6+ncbe/+eTTV
lTFFUG/NyIcr28Un5XflTXgddSoJt5Y7luhA+26JJRi1VYdizi2IffCTs57Ll6UK
7JvkQ46hZqBCogvsUpkeivwnX8+YWG9RhQOB1PJTdcp3Gds2wwkPqL2XyrPB3ocQ
9JCGS9xpoAAn69H973HyJocUMxJLdXO3l7HNUNWZJF29G+Ir11v8g3/jjl/qQA+d
c4pljjDbfDBMvGV+kmQXOeUSWSpBpT1YRJV96wVYklmcCWF8Mp/ahOCBHg9i2y8L
THEpamACmAu22Sa93uXAz13cAgxaDx17yNcZOb4PNoewBOea+UvbRI96KnwdIQFP
5HsA5MIXrrkVyP2yk6RPksDjcYeLw0SUL18QtMBEqPPQExVLFzcJg9kE9ZiWfFTV
NVpp+xY9GiDfqUzbfUx2lWiLmPB9F1PRTDo5wepzTNNsr+zvgVbTCfbNH8cmaeNO
Wm/iuKoSg6nBhl/XmWkwgpFnHLOwodsjrNyqXr8xKXNxkjf38ilEDb0znorUnCd9
+FUte1miuJ/r6Iq6bX4tUi12mjmWpW1K9gyZJSV12n8+cN0xh2L0ocY6mFy2h3Xc
rBAscaMGWpVOyP5bRBaOSP7LZR/Bq3mDtPh4q/LTD9KFRRVIvEZfamwE3PUzAqVH
6/qPXAkNqnPsP3PhTr4lQMDAq6KBOpO+qhk7a6nfbj2gqZGdTUeLeSWpyo/0QStB
ytZBDrMumqTiZk8owoiVrATloe7OrXAnezG4u4KPzkEAhot5IqldWmQGObQo+SWd
XNJ7UXm47ZsR71Q9UXjBrq1mWQxptl7RVrErp3FW3v03WmNi4awl2pR268OML5XL
trQIDy8IF01zaRsaa031iiRNGVK2NhKXKjuxOBIuCEaFruI8pfmZCWs5kTSZ88I+
4BGSmZK3IwTz7qt7oWwAMTy8uhJ8aPTbCKzaJNViFgXRUFaI1i6WGM/s2N3gHQxE
J2UTUinD1KxeYbjqa61GgfvTACMK4xrx8Fx1R2uU0seTHIDd+3dALrETC6McS1md
FXrlB6dL2/hxOQrGy8iwUPJSjTJs0YHyFF2JZi3dVXs04WSnrHCqpYqjvd3Fc8tW
/ytXT7HkyY1dW8lr8NKpBfW66hFxUG9IJ66CXPIYTSiO/tIQTnwlAVjECzAxektX
ViszIM4VzC42mX1cMjdj9bx6eZWelYLe9w0yyV2hMx91mKGokMJog13P2V1XGIJk
gFfmR19jd4q7ALAOr4KZAtX775mxwE9xjzwiLd83S43/b6T0+gYGGE9jrPahUuQf
ZhVrS75hJgxuRNVabKzH11fRCrVWf37FHdgAMiVu7bNOAC8sRw+OAdm1pHTcGKQG
MZwCfINuafKXH9i+HdoOsHmA01UcqJgO2x9cnlm4Ot9r2qKHM9HCJ7ui09x1FV3y
KJc1S9MuPJbO7epRbe4ZwNCHwTmtYX3TmddO+uoO9iNBPIu8meJOGeZ0BXezhbUr
ez4bBEZKTTrKfUJQUYyogvwOrXtXxR0Srn/y5Sv1BJsHXJDZKbmv5ExtWYMvLLhP
y/ou5t8W8ej/0PjyDcgEa80GQB0tx5wRHjxsKOpoK5rD1TGanePcNyhHq7bAD15d
36N1TaNdjaStj6qOgp08KZWhBpGrrur8WBirl+cfX/6gSKzEntFJ4MMvTPjB5qB5
wvJPuWX3PRft4+4p8OhvkxnWupTjUVSLU4BZdbKVN2Wmf2at2rKONU8wRyroRo1e
uUVmtN5Xmc+NJY8cvjNYhghMAJWlSYJ4HpaXSEysGUIMOGLXxcI02EZJRZGrJ6W5
QBFIhCTz2cCEMflXW1/RXP/ns3l5ZmCzaNTaYfPy1KjCppku5/Wyjs2gRYUiaysP
RRlW2yR+vMO0s4u8cV1aI3gIRlMW3LwHnV5g+fHx92S8LmWx+dkxhMpxrLYIB9GP
W5r6HzI8mmqbP/DzTNgwNf3nL2FKsnhOfJSx4r59bYOsnj7y8ZFlF23loq9TycRR
+nqx26nfAx058zZmKfNqkYFN2KlzJqCiH+xQL5ZtTuO+Tz6MfT0UWBYcnO+C6U06
qGxcCdyxGIxTxNmnhxs3nxSQ1YMbuYLLah/jNRghFwZ3Z04MaNynXaP1xvHFr5B9
Am+M0hiJp52UotTAgdlkuWP73TchQUQRW2a0ooTYPMZ0dOyIDTARcQtkGC+TK47A
R2iWoNJe6prGvYhJLTjenbcRUll/SaDR8lGDpEjygddpimpGnO4pM92vINzW5VSK
QX7LAAO/Q35jv9HfwWqmJ4TrcIKt9urqBlSYRC5h1JJwS7wVUkR1h+fibxRMM16A
A8gIgcCiVi0Dm6UCv+TMWEAMWXpledbjMVmcXkxI3zNkLjTBB9TRYBTHKe17AfKj
lNkHR0YAgAOmAAz9OvP4ckbI+NL5dgXFS8rRemDtYIpLQKBkpgUn/l4D/z9/yjAz
L8AEzBccueIHC7ThO5x8dReNS39QrHk5eCKmuxId2ygqzKMYqJ4ReycSQlHLlwFi
rBpecdAxjVH4qpjhz06+/5i+I0qzZiGw2oCmArrJrdq+t9ClIROhocTbyjhamy2f
ba2LqbmTTOFYDdBtBKlMZPD5Ywrru6iK+C/YV9FNnlD9ZJvkCz2S2cycRnDtAsi3
2qE6C/u+IK0C9qa1gz3munAjQf+OJQ+kF0rNOGvvo7FSjAJ7qvuY8Fe4Ii/BPwLS
KQFGptPnXeKoJ5bG+LbyYHCmpx+LfYPxWq9b0xF00REO5In88HhJUea3+yMwBGUn
98GxZ70FCdhhVt/w3LvXxLXPpoCKMEua/6sXFiPrWjcPbcBRpzTZE+KysO4wL1pC
rPRGIUoQsxfulN86Z8Q25vR2y1J4fQk07l5e5Bnv9O1TkeqEtV/iz7M687f4L/Ir
Wdiaz1VqqkQuNcd7a7N80SFMwIYDYfXnWTZ9UcgSEqDafkmWJjCXD8G0ntJ1MmEN
sn/BqF9PABlNIQ+lrcAaBmJthjff2HMnRagiRfjGIy4eeHjVkBjRqkaifUw83JA5
4DZOcRxvYjJCYHppMUvjWsT/A3sIzDAXaoYoHw0a/oLcH1xk6QZgskwcmL3+vbIN
5SOJIWpHLDgm8PIsev6RIz8HNb0eCzxEPkGOS/XOnYAYdL6lpwW/bcdNfjb0t8TC
5e4OKw6o5JJWDJXWoE7ctp1KRozEi5kYSPXoab8bTWIe9zIjdWQtPlPRQtlPnjCb
qvdiWwyd5cdADs4RjRjAAhqp6V27W+5IV7N9HNfr4SgN5uUQKJIfTnRCiPZVsyEy
YPu3yKjMB69YfH3rqXX9voM/+Hil+SfVAQKpYkEudS286Y26Ls+wMFs1xOYr6S0r
3SOxZR5F+lDm5q16utZ+S2UanlH7F36YK4IDOZGofmQc2xqGtm3nYLpRumuct2El
Xw8E7GxRoOhuiH2y/BoJCwZD/j2gTLNo5itL1LKo3KUs50La5JzTXAVl0bFxHv0a
MkobMWbd1/NzN0nIeF+NxpFmzQ7EgiplrLT0jReuVtKfA6gE4L36Cvkc2PyCV5TT
qN7Qy/7uYU3IsFMrocZsQgObmced7k7lLC5sBtlBpRt5o+hXU2JH9UxmoBDil/5J
6sr4u/XSAJITMYBXmzTiNnZ1O9GgZKoWF8UqsWMDBamvoz2F/FRfITvjpabCd/At
MNLjSX8qHI+mxmbAgKMIMd6BseL94rN02sycotEm87k9qySk2qIvDXOQOw2QMCzy
+CcjtWqIMfE+Lv/XGVdueOPW3f9icOMxkPCfjXc4uV3HeeIf7wqa+zcGQ2EZdU5z
eASYOWMIg4gRt83Gyn4U1pgQmtJOPEEljxTXmqUQqlz3vo8cbdIA2KwoiVkrdAxa
XkNqfm5PjjFF8EY9G0CYHlJMmjKsPcqGL1LgwuBtFJVOgl3fhbE1JjgMYucC7azK
EodFpMxz5JehSBvTyKbl57MGuMmekcVbCCZr3t+V1RqYR2g7Oi/Ilhn1cq+77EQE
Bf/YI0EJ5s014CkyoUs5qvAGTrQsCve5aaDFE4ISjqo0ha1U/2B+egrY5Y/it4WW
ihWsXrgnsuBVz0T70pTKqAOnENb4/WejXXidnf6GHag6pPfEhsnjZoevFXSGWPxq
k8y87BLyKVrDrZSx4/YYtn8pOcJ6JCZqCvsw1e6Utn54Le2W3q3za01OzvqmQ4PT
pisOEnMxo85s160xyStAy9dMnvyA2mA7PcdCgGg0oqx+CdPNAHbEXhM2nqG0a63B
TSVkPV2/NTmW9lyLBv0/rzwVtZD40LhbR3OuDE/lPfB8j2pr5hzvbxFdiTJyYxU+
gq1dJjoVgp4muRv67cpq3iAlynrFp2DZhKoxDJV8A/bSsylAfwjqMhusE7he8ost
Od5wDzlsa4F1RsBQvfQq8qFxa/QjyHPcvddJX1HqODuBFY9XcQ2aMSZhlWmydLHa
1rgA4hUzb6cCpFqp7Ch1mBqqzRA2PZ1+JGg4flJY2IGZ9KuTW2FzXSraOG1Z4XIb
noLS2Q9JcZELutnkMy5SndeUrCUZREwiLxgl9L+J2Cd8rxWR+C7UjPN6zfFcZihV
yCrITP4pP0Q7qKA9ivQGDUDOe/PrIavWACNoNlHOEPEqprmreO+e4plSNqUlo+eC
sRBRyCfgj+tUxGxHMAfdwVziu37lZYxgPMGxZ3zZjtvz5Ixsbp8cPUyCg5XUpFwK
ftvRCQoJZJerjkrjUAvk6M2i70owSxHV19eq9SjwRRCp2CxUPuO+YXZkNpEXNAkO
EB0Z04EHu3OnB+66zUH0C4J5TfOHlEbtFBJOr+DaUg9/PLu1feapyy389iY4ncnr
TTkk3uDIbe+OTno6S0E7MtpjVFUmuAgwOZXnGBITvOmcyNF8/lvHDhuhksGk51Cx
muoNwmiq5dRV25wz8SlMtmEcKIkUNbeTe0UDwJbKfqB37U1jkBKqPn7S7grSV+Mg
JwyaJ2w4Zzm0FVgcbqkcsgDo+dl7bLnM6pfIsvw0kEVJlqkglc2MwH/SdiuxJgDw
VXeH4z5+9jM8h3bq3BE4i8bgXBWEvhMGg4/Q5XKkeL/AsTqsZiDrz3zNRFsSxyYR
TpSRuwkCnIxkgy69z98k88DqIdiwBGSIIOUiRLR8OsGmhEgvW+Fzuz8Z7Nujwvoq
f7xMburH4h3Q9id6VjF4AGCNl10aGsb0SOjyi46R53bivCQZ1gQK09CLJGBXMs1J
45yL56MDlORJ2Medtz5boZusxvipW8b+U3S16xdguDKy8fxMPzr1GNrh8RhZsWys
+PgnSPZBH+fQqgigqASmxeEt5MTSWFSurwVSa9hhM8tEjIniZ0wN5yAXcZ/OLC0q
vt8MPDlYPGu6bMpM6N0P34tQnKVo0JHPMbihSddUPLLp0TcULGfcsgEPd1D05+Co
RaBJ1zCqfdFDFEGxq5R/5n27ogSGHQvNj42fqmfEfIWQQk1Nk3+b/WL+rxkYw4Ye
wcxHmiABy09DFXxvXfziXAilDk+x9tE97db4g1CBRnCR3t0I2EL+vhJ6K/aIkO/j
daRFaz+ElXsoebHjb918opz4TGKNw+wC/9rR471J0ONtqkwQNlMDl3SFVzwJjknY
BaHojWknZ6WfCtudohR4gnP+8yh2RuJuyH2hDZtVVsS6O5UCMLOB0aEppvExoiqC
t8+j3ht8plb0FUTLWtLn+29NAd76YOROo8Fcn4I+msFcQ+uGmZ7KdkdrZNdn7Yy8
Qq1bdeAgyiPc5EG+tWXsfvQV1WvIYuxtAHLz+sGrUs1T1LN2VFhQrXBCtwKF8rgx
5Anro9qDG9VIiDCvAjMGKvgc3bFC1SdPQxZfRugJiw4DOFeOEgerhoKZBn8Ok9Cy
p4vnZMivNAnFXHmeRuinbmYLaz+M6nY7ocUQcpvB74MS/qYs1+fitq9usuVQdVdg
KkTu5HPVX7ovTltfDjfhuQ3UeY6JUUtAuNvdgKP68GC1Vcj89wzdjQr99m+IjXKl
hJEHiKBb7QX//8Yd+PfWJmVzNW1YFjcE5VNDCwj6XJAQBHuGw/3bcmgwvy5szg5+
M19BmqbA0vQbTSDyVgbpkWmUAvnguXfqLKlvL/jc3LGtBQDsqTpDiNrfSu+FslM9
lzcIfwQjlzQB7/tel/OHmHcsli2EnUpB9HbSjaI+EMPL93jDXotwjuRDUkzae6m9
nuKbyOaZka6Pc6tA4yJDyq6DYCiox1GzDWeksHUhMp8wBGT2BDLLNskL3lQNrv1Q
YFGRiToKQbeKDhBseF7PsHD8LlNTpLJcYfM0/AviLgCADk8Xd6BY5DUhG15Lv3Yu
aPuBCFlHSJiKpI+LDl/mmoa8aYPzPtq9NcAR85Mx9EbTMt5tT/u5VFlUrS02OYZC
vJn/P5CZcaqGATUHtuFuKjMlge982kyOjcpfo4zXWFwxnl3soav1OO4S18fhhHGT
g8bam1h/pvkJqGZUWsRgxmSRkEh9b5TvMco5M/vZNQU+2bvpPlh2uc8u87MWm+Zt
EcUKi7O/o1Jv4tVGZpPCRc7C0lImd2ZLae1Dbs/Xus0lWxsbRUDkT83Uf8PYaylV
e8yPiynQ25LtTtEpmOh4cP8FAY5UoiGqRq6NbRLvmqcaRWTnXEBI3LwoacTlc3K7
JedCmul/V3zP9SsMbz3ECtt9kCd79rMy6cRwjB/6s6Gbgh+CjcYOt5r4T8pfjvxC
CH21+cXJJyQ3KOafq/+VcnG0uPlLqy9/GDC/KC5AC3GzpqJMsEVbWalbYysLVHuP
UI3Q58euKIDGMiQAD0AoiW8CtCZ33t8s8LzydQhz9MOsSEVOlQ9kiy3JySUPvQgB
ONz1LAoLUryKRRXNeJprZi5pOF9t0HzxfW/ZtWz10Be7pZClW+a2W+W01vjmrtMR
8Jmsv6sEuYX3OfyupX2s1FjBf9wruYMuLbD268Y5ZE0tVr9zH+1cFUDph7CzcZwM
hj+xd1S7/REy28AHDkbDzQaDiccxO0yw5PBIsCW9dPZIKGLssr+y6QBA9kvZyWKy
8hPc0tmYGRHT/pezOilT/03ZthO2aUESpUPiVZiY8+8r7sBgqK2Io4XtuQLpqc2l
T2X3pkOpxIXKZ/wSgbexoyRAa5SrSbBTP/07N+fKfoMq0HDlH9/ZE2xNNlf8Pxu2
LRlvXs5S6M4K/EEolPdXcxClY6qJLBjxT8jGBugbl87R9c0WabsqbnESxS/z2x7e
a8dMUyOHIFDJ+wl6I6uThzjCwzgBTUOD+MHf0xRqqZoMXXBHfIqQesHtktFqnnoT
ZF4kwEeRDt7Kq5tJKH13xV/0wgG1MLobJxbvgT15MS9UOTSq/y3ld9ykfpzIu39D
xbooDwqMvAF1rpFi9vrsgVZKktcsrgNv93jp/qVnOwnwzKDhYSzFuy19pQU2grQa
CIP0kSAVHa5kHWoxwArkdd7tbyRYJ9q7bwNzAXIyc+mBNSVyAGw0U/wha+ZnuEru
BE78fHKr7CWCxwxnUDpwUNKIiIsDAAVd5Pae9DJn5nJKdhd0Ox/jbPAUkFA4rpUn
NAuoKcfP/eNlITVpWgSUotC5MrCDZujZfuAbwkoAbazO5A7LzPwd96gYQJAWn6AK
Dxa5iW3/qs7bcLkERvnrIsTgf0mgX0Lnv+I+MyL5ChWVejRT9LN2ldxBvQ9oxcK6
QsRCb5FEWwPPo6t92CeiCrFxCArRO4aKVcZNiy88YC5Pmy181BwS16EX5e3XUAlX
vawhFOvGLhKbh5wKRhinnkzZVspVrOHAcQBOgBwhdkXs+LDuHhw+AJX9os3wEZBR
N8dzA6mjWmQULsgj4IRyZV6+cG3xhtIuBbGfsP8129CEDzmZo39m4h6fuQrCDqH1
dMq82tzcYB8ibHkxbyjpNBO9s1ID87++HssHOb3RriLqLcO9H9uyjsfVqbt9/QCD
oI8hF/cz+XK5daeDdtY22AWSspsa/oV+AvfIsKBY9HyTrvrvi8O9uqqkR/o3BE2b
zI+AvaY6lUbA12hnz7faHyjoM+6dO4YvxDGQlPNlir3x6x1FuUJ8mxP+BFPJY8Kq
pm4mdxypoYvQ3rSJc5Y0ySNclDjmPfSHKJ1fS6BHOJMwYu6T5ZGNJzZ0KRp4v7ia
RPQ1TLeDEVrtFqs3/62LjXWzzLhU8tKlBrrg+H7XpBDDlS0S0bGTAtKqclfUIOcG
D1lsT/Bj4cQXfUByrPnIDde9UXisMcdqcoCIVOPo8/oaa9SIxpHR/gcyYYt7PS/m
BcgPilgjB5Z6638Zq6qxwl1EFiwVWhpVWFiXO4WplJxAX2i/oUZsK38/B9OxQLhj
yFwsycaFLAJm5E6YnyMXEMdRaHR+pQJr93/kFJZCMLXcrJuYkeZptFp1v6ssYmSB
p6bdKIix/9TLjl9rgYKYHxRao+KQo1B7E3dJrI9B6ocezdAQ+lk5Gxy6COcdXPmp
RtwtweK4YukrEaILsBhTuD58F6zbiWTRIoTC4WHzJc2Eua/Ci1JoC0Y0aMJgZZJ1
hvfAMLXEgEl9ek6GY5cqMbUG/CgRVZ9nhLG+LUPAUrLAMe0+XzC3i664e5ULYwLK
5SIK6+zP56r8F3oX5jO1a5YFcZZEfIOQ+T4LQhuJprPJmRkxSnGXJapne1m7Glp9
SNRgiYqL/+w7m2n9Lf837ZMHLnMJFuQz7qoA0XUYjnjTCLZdmpOndMpr0vSAuMzt
YIJJMG6QXxm1nnWbj/ErzCjFVS+vU80RZ+/dBkpDuozcxp1JSfCnHzpBVfUaBZDX
xh0kBXpo6J+HLm34D+W8iTAYLVzgnY0+WIo5gdiZ1SKNUTeSgF5JDq1RFmJy1bls
7mor/+/8si/JtDGAad/W2W523t4ng11Yq+UVpbn8gfk8bDO98JQLZjW65d5Dsd2Q
oE3Qp9sdg34FotBFtA5rpymLZIUz5RtIQQCyNzxI4taldQYB+E5SS5GCF6T7mpTP
tlvtrqd2Xq8plTnOSuLKL2c7oi/LE5WneRQ7nrwiyrqcX+bxMJpZxQ/DXE90kqTw
MhxhX2mqUzJ9kHsTNSMHF4DBNP3HIKSTUaFkCQiq/sX8xOeGkQqeMLYVKbivHLYO
28B9MEnZAk4n/rczh2JTRrz6aPZQjrPn2+SdxbscqCbYHaMLl3AsE3Qra2oCP5tK
2rgKhbnB9vNVm62rB6XmpuT5+66wQ2jkNuc4q9iWxeTs7D5CJa8RUNaTKRGolEE2
ib5oovip+t8NZ8XJGE3CF/yEjMXQygXegV6m8Ywq3blsSCM2Vd5tKdCdPcif5Tos
ilotr3uHD87/tcjJQ7gMuZ/ob45CFvHWOh25j0MuSrwsM7/tVY3R8Eh600PDjsZ6
4D+zthdDyyADfq7ipk3lfWGGa+6FnNruwq2h8BG8Tt3KmNe2C+nJlunp+zremsVq
imzWMIA3EkJZRHPERvLJ7i5OZvNqHiEscHqSK9DtXTnN9CYyHWO7u4e1xdgH2gIx
v7ItkoumkiX7g+ZhVvKPNTl4tpnHk9F90VKLFRJ21pC+U4bMEWlK3SDJ2ZRGo8Sj
WsItDjaxL5pT5X39pLJt08BCudzeU/E1RMh0/5k7fIB/G7lJ/fvR+cgHw5L2H0vk
N8ftA+w3gFvUMIA4gWnf4Bs01NXVgJ3i6xzqhYnUZtPAPw9G3ZdiDct7DIrK5P9v
9E+604WzScJpEJp/24JInMVu2AgYVZqmFIuTc6tN8bLIf0mZhF/YnlJqV+dYB3c/
OB8eD0HwjPvN5aDJf2V+blcjSl8aiinqy9UJlsX3dxGrwymZSUJd5VyCBeOvYuld
rTIpFOlUUWhKL4lNgXISf9vjJNyijO6Yw8XznBJXdq9zCcSCjDYPj/cMJ8pwwbyS
8mZ47rL+lzyVL2AuCMhGX+dIQ++Lf0O4dyypGy5/oU3C8XL/Kvt0Y/+LlaSqFJFh
QjNkQLyRrVR4zXTEQnsp2zT7zj8pS31y7mwociGnp9nHSJNRgfHi9fKbcsce+Mai
0Q/MyzYTtw0LsihqRaLUewgBy35XI2RowpWJdRALLvne5GBeIPNH9ieJ4fKDAOU7
TLZuEjcSYcuYpNlZJblBQ3kAox2sJxvN581YLBlSQ+R5BCTD+/7ruOHZ5Ngb5xrU
4yVSKC+UKq6T0oi5ZEQfTmHSzDUUmhM96dV8EjvgQCXncKx+wtCvh9DHNQnPwbhc
SDSE8oNLz5iBmZhjT52yvq9FJmzESYCYAuXxgmsfBYzijsggh486j87fmaV3ojaH
btt+svnyggGZVCOltQeP5dxm9fzINdlJ+whhQlTB2QFx4CZzvV2wflPINFC5EA8K
GaunR2EhzzwcLGhP6snu/51taKOyWdBsPye3sh7ljUTDYR7yCth+8vTEHMx0v6EM
uXjqxg5M++ROiBjNiVcadv+S9GQhXdlyQdnzjX83KJ64B2nQrbDYKFEW1ING0flF
bRL9QSv2spAooMcPa0DLLq49GGJpmk9tyVpejo4uztncYhlSjv+Hh+7igT3ZfPvr
EKtnM4MDog7FhNAgkW1DQoj3u9kJp9GiCGEz4b1iq5aEZSIAXh9LDPqauGjs3Iul
4rOX/loNAVFT0nLiZGFNatelRGzrGv3yoGVvkRzkxdn7LbdCN8KPmR1eb1XPJpoT
ZocqICFjmLE2BKRg843mP8bzmepULwgi62229DHG/swiPzYRmZb4LZ5cINCCMTJv
ymoJ+EGoxR73BXDic+xnK3TyEyMavioK3TtWehpUd9zQNrbnEVim6NzYeKNiGWgC
0kwu/9xC2DDlyQt45PxuEQOFMayVlUwdOvcwEpw5I/8na7DD1hy2fY+JQYqldUmW
V0K714t4n8Sg6xrqqN7G7EJbywtUv9QSSbn0aNO3khgOo4p9k+7IeVKeOPoszpIR
D40G49zTTlsr4ICQqmJCvbw0if817oxrvwcotQwpiUGgckn+ALu5Vpzwu9t1rHEv
CSk224DlN9gOpfyxkWUksTHzmhxUZ9qTWHjtXKujgUSOzpq0QFG2DnlY1Lk8FDY+
6tfXRn3dSr+JkZAYna4jgSG+zDMqPBNh6ZzOoklNdWbtPck6mLDJ3UkmD63FY46D
Ikeu1PqQvN0Ue/MhbNMUuIIjkX2j0KbB6u9LrsmngXtSGCm+lYLnnCaNvYCP6e5I
X5hYB/tye+KBL2zf5TbQDyOzBTQxfakKrMU22zw/NLNQ6L6ru4S1pqAigxu+ubJp
6w1tFXeU2rs6NjZw/x/WOXglnJt/RedgUxZHDBYQBLIG0foV5C9geiCP6wHlfkZi
jIh9hDW5hbvFg2PcU9Z20tbsOqhQwy7JL7XRRz520nwlKz4ATFdffl7j2/Ti3JYJ
Y1KwDD+wzXWlT8wL62vcQu7xiNab+SJtvf3bww7a9pA2O4aPD+yfdZeVhqlJ8mlY
gt0qkxAY0AExpmby8Li2mX2QRj85l3/xcHfNWq1v7O+Y3hnTtLnHxqpZMmIMupiv
Az8UvOTD5it6m2Wy2tIHql36xz2mVT9lsterzdSdyTWg7F/OzIqU68AOPjCs6BBa
tkL5J/wgDk+eyCEPTW3+T1S/NzcTvr2LKp//v4c+MsVBnabgMSpCkqHpRANhhE2d
AnRHy3z/Sn7yLg/MbhvVq+H/TBRHFZqPDTwSIEc9N5Xu0ZNhM7J54X/aMXHO6lFZ
hdN4MbSIkKS7x5sxPMPHHpmDu8FOWJBli0n/eWdkhalio+ZMmM/BYvXTB7CvxKkA
XkYvdBwm8+tXCgkieed9Hj2NFv5lPfw8TeTAglmqsq70/oiWrmG5trqfags/4WAF
Kj3gNghq9P5OteA6fHdzd4UWIuzRvMMjY8yE9pQn6BYkXLbu1Fw0MaTq5ecbYB/8
XCM1QHamu/Id3DojVx3bGD/kGisD6glE+7FpgXeY+7iPEujkxGSi/vaX/bEc7tfQ
/apKW6DN/BqB7F5QicrEYnnR//cLTwXRIgRckpcfr8FINFSFENmzqmI6+OY29yT9
zumHQgIjOiNnBZgOYgG/eYuS0KbxDjZ44AFYvb0ad2S8dwAC0omkhsbSyw8kKWyO
+kZWhQ10rWXwbufAVeG655WG3UJJGYTk4TI2aOrPCh3Im/GDc4NE+dsZYQqgZ7jT
gAObb7Y2mqYUDavS0Q9SFEkxzG0YQUBE2+DA9s8Se7Sa/CGPZvLXfijmveE7N7PF
OIVO+gjtOhHMUekwcP63eHC+ggktweu3VzC/LJOcU4fI74M/MtDvvmZqONZi3y+T
SEdz8uoS/KfAYGkAtIWVIVUrvuZUpp4pKPdZi4WhMsQSAnQv/7C8eHBWuzD3WOSs
ybKQpb4PaHKBC075wWhtBWD2lBWWFisCr3RR3YAFQM+Roxa5pTkOnTWLtq/grWl1
tdScLEk9NcAibLoodfNcKYgneRcmk4DCMsIKqIps5LCFaFcr8wuOPyjOc6BchMu9
aUZgneodKLc659EgKHPArRXHTjWzHfofgYUo8dYhJHiABsSa12uM7uT2EwAz73WR
yID8NJE2uNMo3eSkFZ2gsuHnFHao6nEDepOOVBGmnzPiuzsSFx/MeeoHv0H2mrLu
p/VD0gQSoNCkF9hvovl8c5QLzvxxXYcKpl48s2k3SJKUXoO7MAD/yGE/bSwmo6Cg
nzz70xizbHxojslUtMXTv7Pkz0Rh/yCyS7pFzTH2S3jVN2pbyKqvPiFgQLuNj91B
KzPhvmMnXMjwVSx+2KS9M8q+8RMsDb8fi8XG2ewDMftw3YxZ/8zCMB/a8WfFFajT
u2r2ITwfOEBxRsDwwbRbb6AlCMP9cVexTOZFAlVJlznFiBy6MLz2Km4WS/RBtGxQ
zArtZKD5Tx9TYfCLkKsmhUAx/3eczJplnf4OruV9QVO/U4YQJxfSxjtbLRN8dpSt
cUJbnPfMt2wC2bZ3hBEpzgTPB6ew02b7Jb+s66csTOydXbFh2Y8bBJPxCbKZHc+a
NRbz/pevCsVWv8CdyTsOqxJVEU9RjcA4/N4rhsIhTGabT6N56/jrfbcLoq5j8lqF
5nQSEq3Bhze3ojWUgrDiJ3Qc4IPaiWb0amkoLjjYmjaKrddCBTICwSuuQFwxrF3X
1Z96K8zQ+jegZa0XLiPiCT/aJlnW6quAYzSSjbwdzyJSfoDHZATfFYdRmI2t7NCo
slfDZvlbBgWr/EzDk+r3/cwl7yt9niK7dT3pTjAnkCV3lXGho/ETIyDc9v0GsIVI
hkkzlgU9n33DVjWAmak+pvmoi8IY4iLgNz+lUDNHWNjGdtj+vkwe3oTBCysaCvbG
wwqb/APiNah3mmezdS4RXmxnpewWRPJQ0BgyKyMSr/R2DK8bSd73wukZegQL+ZRo
/hu3OVxd2hwW0t78EsGZqlXhHtr+IJQ70DQZQy8Ig8OZxvrmCe3sr87zc6j5E2Xh
znBM/TXcPp1OAY4LkCGT3JxbnQAaysjXU5R9ptH6k5cuLwVacxzt7h/t+Kj7xVCt
mpx5vTcu6YpB3nGEa1mTE7aukfpcaTf2h34vEJijClorDO6b4bnORPhkNzxC+PvL
ilUtSWFNIhQi35nYv8tpV9hdiBq0lPCOfhW6YBBFniQDRM1Il4fmPR233/72vgbE
kORDqBLIviCgO7qK8wXgsFL9VePD0UbPt68RXgUnw3itTtNpPEWwSU89Wk2YPZCY
splPobAi09ffbgf3cd8bgs2xW0MbgzT9N1iiod1qBs6Kwyj1TcKOxwj53kCK/dXB
baSAbC0Cap5oeU6ds8BrbM8hCzF0XIkvpOGKX31weUFCIxuhYNUlotUtvQ0EMgqI
Lg1iGy74+Uxl9K+lnzXVl94XNsKLkYwKdbETmrbq1ivI8WHJ8VUepfTeCVsNnKId
XWzBK63HDGKnUzDGpNrL0+jnlf4hRSK9EuQ8Q+99wXj0S0BWuNT71rcGus3Fagjd
1xbF0Mg8qvQdvugha/IQHha1Tj5Q4/z/Pz4BgJ1hlzRK8OTwVWDhLXgTrKK7FHuf
xYuplSKO6GeHhihsTLrzfEoKB2QRjViSKcRHXJy4ulnaWFnpYuQZPEjvIugMvn6G
fuA37gJW8hNrRgaoZkYEb62xzVF1RCV50yRE8+QAhZYLV69fb0z+hLDPQYTGCFAn
jfa4zLvghiqdTOUct9TrIh/7+KkLqr/RMW2tdaUdBgHORvUXFOogplJtoSkd7+Q3
lpuDWF1A3zWlKag46uSS/f0xz5g5h9DMUcX/Abzh3ZsXi/AOSlTOmCEoH5hUxrJC
9uiLTOSyznEgQ/t/JWYcZ+c1mKl628JM4yHHzQUNKzKcfstGVkEMiXJfSutZFdB9
K0jPG5CrFQBNirPtEcX5YSAWviWmU2bqbfPFBdFjxdU/LU6inknTmYjKxrs1qeah
k3Z7LK1lNIwZ4st2OD8YLiS7cGrgQ33/UM+chKBlCB4MF3MKaF95MafeuS3M1w/H
OcDa5XNyK6fFfzVONkjJ0N+N4LJ6pfg+bmW0dUkZOSFr9yse9cXkMQtLJ095TC3x
tuMw/HwiLy55hjUMzFvAtv4jlsSh2MpOini4WLJvYNBAMAdKTXXCK9weTD+58Hfl
sKnfKb9X5hNO91hrDSyA8l9Px2YZron59EJ6EmmZUdzp2qszziB9aqQ9BN4KSmMU
hUOlqwedKdQ9Z3tFa+w3TXR/nIdCIEPKJJxTtHn4hHe6xEPnAKQlUcA0jb6KCQDN
CHUxxTMb1dmga9Zxupnw/0if3IlIUE+MJLMROK2jaiMXpwSvXL52rT7nwYY0Xwzu
aPiBPt0BJsdoOF7lyQ69sGi/b4x0Ttz+WxoDtDZ0op5ktF+N2drAT6gAokT2zPax
5xnLFIgZiCyT94T+y7VzvnPWgyfME0r8B67bORoQVpjn58Hq2dqbJOwyKkJwDmC8
k2uJu5BzWZj1Tq2IihkiEaNYIkSU/SC32ilGTj7kVDpjjl7IQ3HkPOGuxgUXWJPl
DXpzQMja/+Z+uzPOP/1Hf/lAZUdok6EipUto7tcKUTHQ1z0rwTqFEdY//WjhZFg7
0p4zzkJlsunRw1nZLHlwj5t1s5Mj+dwwI+w1D+fQddLjpAAtSfTCofn62h0D2NzP
Dir986pzuVvgDVK+rDE6mNY+hP5FQ18aS7NEYbHgjcXMy6MWXrdPbylxhoovz56i
lWYgarBmEUGc5CtBm5xAjXw6QSe9+jDxPjSpI0BFq/OX2+WGYo8Iywd+RUA44fam
wc0MelQ2G/ZejN+7QK3Hyg1TIm5EzkvbRx90ilt0qubTTrDFSmnf9kiTWqxZp3+W
tk/gz4ZiQeiYS5YDC9OHDauwBrKFaW3ZYQMRV49GQQDDfFiWqp8kjL8dXtWv5/gB
8G4snJqMauXKcZpp6ZWnX+sKTkCDmZ8YO6Kma052t2yli/X04vklZUg8fksmZ3hb
lCxssKDjgpKlVzYXSfd559bmZYHC8ysV79dBsL31pttAfFwVsjUtcp4uTgNxqUA9
Ctp/Ah0WxB+8xcFavMYr5an7vKVQFCfZtPUQsEFSbd+ScXGIgIyFRvmDICJFabQI
/Ee3wNAX7aNzbyrt47uiEQW5s3GpoINf3lB1H9SiQ78iM1YDjQRc+8z7OVR9n31j
7geTpGFDAOcJxK/t917C1Q37HCmZKjmBjpQ8BNYPjyFIUhGa0tmTjklJZsN1bSfY
8QYw3rvii8RU3mTYaezHCLwpAnIJbGbTEtyfmWIjgRui9Q74GNojGam31Ld/TkdY
CLIFOOHIYXOQkdVK10HERh6UcAXY46dHMllwyZKATiy05uUfu3NGhVa6/dAdTI0M
2A+VDCJFoQNQuAtqHELVcPjlO3/uOQ45t1QTxVbMEeLh4KBY0Q8cS+fuKp231ZFH
x6X01mWYmFPtqWTA7eoh/bgnr0WniRwCyb48qykbAV0U89czKiwUA7r6eSx3C92r
P6hELmwqA7l/A0f37LOS0180NEaPGO2OVITALzWFQlzjkks19spjK9rhWllpkm52
N9cGDEE3oR2n/8yT2qloo3Wtd7O1SQNfnjUVoxCJ+lR2FGdYLDYnahyBhd4iIHdu
YrhyWfPrYymcpUZGE9TA+lmqLleVBAMZrFqzKMMulmLMJYUJ8iaMQ7U6HKMmFh2A
rCbRjQ1IrzSxZ+Kp8fE5iGJbE0STzB6dlSFfxRXY2ut+zNKB203AGc/Ycu1E/xQM
fM9CzzhffgMU6n9sZjlJXwzNgA8ozIx7RLx3hQloE2QXNYoG5OFDJ2nybsKzV0UR
DQa1Se5nq2ckaPwWMwx066p01Vtw23mYzubSSlrubdHASaPzH4rstopTguMBwmc0
spWkdFAa5RXkGsS8ZePvVo+FJPahaIGtWYP2VQKfLCLlz2FL4DM3dQ7rr0DsUF6Q
tRdBrGHSZH5paEqy0QjSzMgQViOIaism7UPv0Od4ogUhRva2qZ1eGl2174nymwjG
BmyH2Pi/uLthaKhRgDCLhXbvTGyOpGewolwnTGo8OV2GdwjVwMIFG1NfWIfKk6xw
bYu5Q9oE1tQzDsrI0ECDVzNajk7OJek19v+B6YoXz+C9Rg89AibcgyIN2N0rcO6m
0AHldfjqXXmkiMj4ExBqRmarRCwO1i+UxaMeutclBIxxKKmpl4YdcP+dBSJT+zlW
SDy7Ki/rX58puAaqwWc3Q+4VCfOTVD+GFyGKuBJoqpN9HodRg9zkCRKKtH5wt3Zy
brqYT9YYIiIvcFPFGGeyjsXxp/ffdnSHNZBNXOtZjhPsEvmcsDi2h8esR/4P9MCZ
O9nMhih/SwL6qFOb7IcryvO+1KZnDemrOe1uUAk+e1YgCubx0CZtGFpr8XIMouZW
ajVJHrOozqGl+IwOpiw5gD/er+At5whm9i5bZ1EaG/Svvewx3JEoJ/efnJD88dYD
9gE263bWMhNvPAYudOYQfW3o/kWez4C5THwtGvkST82lYI9A51o+D5E4IQ16QkUO
9lLnNbK2qB9gweXWuZUFAcTBVq/o3c89j4nCwyucbDJ8TyGsOyPhm3dCHNJv1uAc
liBmGbQYfmaFGUnBd0za86EaelaYnUkXTtt2WxYXFFWTlW27mnoVLb810J4cOwt9
BuKkKWXi7i1Hrzb89AQqpH8SZIAywduQvW898CMVyz9FgkjnVOZp7QpB2HX7folA
obcQhUCvUWPIF1TsIMDOjVjnfTh7qGWuAUU5/gemLehgbS5w+xA9fcgBPQfsL9xo
AJaf7mPqKP30kPwQvbh30H/QePz5wwENVbQRgNemdzPQ0lPoObJCV8FWXHSjXA3z
h8QQHmYcB8P0EJEOqiYfg6y5BbLmSkPIou8dfZeR5l01td914iO/xAewxUI/Rf64
zWmDcbJxtyXuiRN8KIgxHwgo4l1hFigzDxfwIwZ0qH/WfMQvfUwAPQ33W+M5btZA
kS/FXfoAs3j/vh7K36aXQupJN/lHG2QX3qq7Dwik1QTY9xUZoEeAh3npXpjttPDx
5BiLFbl4N6Iuol4fx3g086V7shHEX/OgS0+GE+F2kOGlTH1toWldHAjbU6kckaEr
0zhOBOmIC2ta7qOi3wasRM0Xns68G9hbYYRr6ZU5X4V2mp9e+5VObzmK55/WSwtv
iojdrih8uPv41RudQ+78RdFjC3WWG5sK5plwFRg5eweGq71bHmAYpccu07W/XRsZ
ieLYRtLVGoN8CqFStWfahd0haij6MyysVA4tztvhfTrgGU75Gynqv1I+AEiT7UfY
50XnMTZObmkgdKEuhLPct3WtSI235Slupy2rZiqcugoDAbjoVoTpmoFpAsod4YTm
sU1+G4QFw50N22y52iXJZHroi0RGtOBDt9gJqhIpYLHFQm+yjWg3UG2WdfZnWuqp
VzgJs0XTH/pdnxh1fOxyAWl2anOnGRczBQ0C4ogcDa3nakz20eHxvIBq55xFS9I5
cC3xOdIRJCY5BOZdkbaizMMjuIsI1/Bso95CyEsIamTvKzuPHZW5K8JGGsFVrrCE
h5t/F54cfh7+pUnrbdS0GqAyRPP7rxk2zk4uIUHP5g+ExQJC5H91yC8OKlj3xYkU
lp/0NA2smiUppkBAIc7RysJIDEwWrCznoO86NS22yYM8SeyZvCOaUx+PZYoDCW9e
fSpg5mXaKHYZKgpBvkfx0lIACUZXmthMPEF4O7iNn/48G/TIN/fnxJqmv8nEHJNv
0ee//QNLBk6PX4/XC6Cvos5HqNB3rFDecMGvB6lpNw9ObLpAyM/hi0C43WMJFakb
6bdGLRBKFMEB1JSdYntlpmbMq7ZxTmMPugf+WTy77h2ZbmFaWU+g5nymCkzcTWOS
LmILSzOzm9EE+2LE3vz3oGabvSwutAtN8CHrWEpHLSYr6Wt98i3HOErHREjbysdH
dajmWriE6TeBrXoB7EjzH7hH9mt71EyIWE9Exa4gI3efDmfXUB/bnxqithOgXW1U
9+Ze2PwlKdR/8P+6eif7SC8pLXFGfD4mtKpW4eFnvq6WuvPquk99byUWFS9F1KTF
kXBC1XzWa4cjmj3rEPJVGcCAkDS/ejh+WLmINUUmb0eyc7/gBFbStSWNmyDa+o/E
deU/Kh84eTc5x4ACXFUkvkekP53BO69K0nbdEt70ElmL8eH1kMxzr+Q9VNsXDNN3
e375mDLymsRnqDwGHr+jeM1pPQkfMP9Lc57JkQ1dwPqSwYZ3ILTCAuZsK1uQxbEI
UsoNitKY/98OFfVzb/5Wbs+e90TcpvSq0ebUjSNMR8vG1WJCpXZIT4efYMk5qpFu
DLZ+/kshWzA6HzqJK1cZhk9LUTf4R3pHCJ0IYZetLjYFoBY0B+fvLYwgCfQDcoGF
DT0DL0fvI+Zse5gqKA3rairhRBB10pSAPnhV4EZUisWueD5JKmhI7PdeEb/dC3DF
WTCRUitOHns0mv00dABsYzds+H/RjyhoduflVkkEb0J/IU5r/u44AB89/jsqW+pf
NzA0Pjt0mPgukyzv35AeLz6agP/0S6gBvDB7+g//Iu920TQRePAGuEdsdQOP1X2Q
YK67JLIiK45dXrReNMVaLL/0kEScD0TYDS7D5i+QIy5hB+SmngxYvkJzsrQceWOK
WUiuFMSh5DnfUDbhpAdSMbV7LJXhSiFGtc8V2Va4pI0Y3DeaRVGwTzlR9+8grfA0
tLDOOVQe2QsDW7YSHx6Ai8Fjcawuky6xWqtdWY5YSJmyiHjm9VCUiS1OTG8RRYax
Jl6D0ZypBuyz+bwawxlb1/T1h1ZBM3SjOdRBZOSNbcXA4ASakMVIX9sX52PodGBF
z/99HNUwM8P2xUlQBPBC7gXooRqEc2rSTSEIqUDJKS9qBoZ4ZBD4i4SX3daZUjvD
cuIu1YY0hjiRJSwEcoKIXwSDUPY2RntSVM474bpTtSlOUFj5hSaU4rJDXI+GDLQk
E5N8qdBPweSzMQSx7jMHzx5rE1jfGW0M2wyZmwTsq/qykrQJvKor5xOeldBtqWwL
V+/jL0g+ValEm/eB64Aj0LcQgDa99ZvYTZztdZRHvBou68td3k94L3H3BGkUQKoh
5JHlTKYKSqjpZ1tuPABF6kasTN6ebJDk9C6mNKOVCXP++B7XoP5JC0eIZbhSf+DU
2h5M6dI5TWWIprM/vXMQKCbcJRUr3MK0XqxYHgQsgncxqJWCKpN16D1+IPRfHBbV
Sz8y7rczP1t5OzcmZs1Y6QT4ettWxEtXN9ZS4UKJstNq/dTlYo9ZMfujQgQV7yl8
EVTD+Ky4Q30O59oHwFXsfxRfonGS6ceuOY0MTn53+kB6Al8jjFIAOfo6nYOvpg4s
rxRBgU87yeNZFDvvJ+jRxqzENl0vJxeoUrMQzBmqTQopQLONoMCZ3F7YWvW8ahaT
jlrUdMTiqcznpbz24emFf1UA0s32raEh9pRccrzUg15h1UcIEo0ycaV/F/hbrcbH
Kj+AaPvVPXRd1OQw6UyGf7tXC5Upd6buFCTp7o6c1g+U+x848ZCsvsWJaBMJgOcx
HG4HycecVwKQ2cTG8NlH627fzUubVmBU9DtVcjpx/a8NMecLQ9DGaoSh7250aAv7
rUQ49QVj1BVjkXroeX+azcJNx+hHr/c3G64tNztkd9eDZYPKYmlz1RNDsCArcqub
MZaLymELBpQ1fwIU9KtQ/oaMKCkvuhnldblofbvN7G6WCgW/thAykiM0cWbWwFNX
69VbmjN2opCI9TSlP774WVHZAgU0KRlBeCjY5jEcAir+J7YhNyHKaqWiBriBdXt0
1e/rGnEVwTGV7LPkDk8ss9Qe4Fv/zqp1CcDBQR70XzGxnA4Z8Rf3MrJw2oiI4Cic
2q4obq0cUpslve3uVPDrvomGhlOigkQWK5F0qwYg1KgZW0KsC7/NU5wndT5bvj4j
O3c36+dvUlST5OE+LC9fjVz1Xlyvnn/j9mVGeITDEPl8LxtxTrrXyltMsCEUjzSD
bG+zf0XReT8zVdi/+8dMtdNDCCxs2bGVB6KCht+RBg5QcjkgLw5HkOTvnXVr+Y0E
MMdxfVBWNUWwfkBKy6w37vtk6B3gK7k/f7+HQyj8Q6okbq33lvYSIYJ23NPkT79S
W29aPsAahgBu2A+tIjeDyRIV+FGadsAlVXaTYcGSBrejkate7dm0WAZ9ejJEH1Vc
F/aYRLGzkklrwvNTnEB81FX3tJezg7FvmDSfQ+vY+tZJMhTemSbogq2z+ocXTXqb
mzSU7T5u7LFQaBhtYccc0GC3FOGyuuGFjQdtcoUM1/eucQCwTJqI6RFo+S3ilV7r
KBTkpg3TZslHA1Szn9J48fowpHOTHXm8N6pcO0nCjOF/kUfvXmhTAaRTheWVxNol
kMz50ui+fdJAYbAChR9a9QqTOd7TcqUDr2ujx6dccGrWRkCx1o38HWNz57BIUgEH
go+cXrKll8TCmldJ+cUOst1AAf6MUjMuX41UjCkhTn6qg4xlmOX3OJyqlgE4PjXc
toHrw7hLNgXVkcMiOPf4hcz+34oIYA/p4ZlWWh3u/7OYl/vUdiqcFf3F2KdyYh+l
bqGVYAyFPqL1sotbBU3ITgtCXW6yCUY5lMVa+c+6jwrPGh1Gn++SfSMIZItnKkD+
72OJD4vP56bg9gd72B/oCf1YyTT63x5Ffh56siCqMaMPVe4PjVIePRFg60sWworF
tPacQiaZ9Afdfgkt4HTBYH7HgjV3iMBLsyH3kCwiacH+2CnPzjjbQodtAuKAAXIG
MLeZwJEmSoRS5soBd6alZVJKZJMCGCWZoS2/Us5T+f4DXN3+gOg1XzlQPikcJW97
cFyPy45pfR+pSVJzrrUKPk9JuPc+wtUYM0ilGJRYpcdtBMI4bMBaN/JgT8/8pujM
e5kxEUw+sUiWM+Jr9zfzD/jMI8hxSeszw7f4gVqr4+4PSnB3awaANZtswIv11Yv6
VRrh8cYHw8zvEQc+WO3+YHm9Pz3Ily+V1fN4F33hoEnfaYzs1eQMYQLQsLzKUD62
kVBtygMUjplExO8hOpmi6c28HUgyeLw3fALoGMz0Pk+tWJdi32vOzW8fVIsRLUvs
J+L7+u3DEmlwtpW6P2Ki1+ionD4Pyni+7eC9l7+ZApX86lQlhq77PSXo5xMhZDz5
shE5i2KjK5s2Xkz/I7M+kgZ1oQrwluMyHUHKCuhiirDbI6llseoF+zvnxL7ywBPo
DNptTMrJF5Q6acq7b4GObFBIoDLUIMF4Yh6yBPZZyp4TZyp6Qikx67SdnHeSjxwV
5I9WzXKaiMBrnREzmgO7z1jVDImjVhNtaZ/qHHIen/LfvZIBYL0GI09P63s1I+S/
P/2OoSilC/hyNWn2gEAuwO/wc8Vkif74Qs4pDuv6YpSFKIYC0iGACXSFDjnAQA7e
d5FF5L/8Z8sJj7OYMYa6GT3HjhH29gQmQsqh6B4CIahsdnuitixx+3OELYqQklqM
Pn2zFssGusEzbfHCtHxFIrBO4/DKSXSuGEvLlEKHizylkkfmOcsywjrsrqWu53G2
zOPl+OOwyq+vKc0oqLggBRp1f/TgwJI+xWwxYWGY8tDCVE/VIKJW/FbMrM2+foQi
+w0XXMqYRhvOkwFCnGMHuPyEXvaSA6i27M/rNe+xmaD/50LqRvKiisePMZ7CyDaC
e/1i+5f7AIVhdN9DcYlCsbnflECbIOIDywvttUeXXx/j4T0pgb2WubU7Vxz96IqW
4/rMZSt+1oHHf+npD32ekj4ZiIxCWCm9PQBsrLBmBc9kswgnMLaMKNpcQ8TQHQ+u
LrsBmRdCbDCy2BSnxp/SfNLIRXqszEjTfswD5F3ytq4m2Ir2VQO1f/8YSNho7f2A
EWlAeJo6x02gLQQwxlC5ixXdBLHw0fpCNtOHnlHuZLK2iV5C9blEkz0Imja+QhCS
WvMfLscoxZHpyt64FItB6J1W/UTFbxA2NRMhI+pPb+GLkfAE6pXI1r3ZybYczit2
RBrtw0F0DP7PleSKKrTtV0fBcyCJD870LNu8BFIbTAWeD2JykRXXwyaNCieQPdwy
mPcaX/pzhehNDBILj8yJ+5FDxi2cTd7wi1TjeSvoP3fsrlOnYqvB+LVGmQLrKANp
MIGXpWq9tvSkGyhivOaIh45G30yLMoJI+7K/j8gVfX8c9A/+UnJb8vaJdm+3RRsO
X/U0OLyQjx7g9eRDEK7+bMTPerxX6jeJKgyNrsi+hJ2l3pi3VGtlp1HRcpvRJ+ta
HodDxRQylGD5NPV7YRnHIDL3KCmE63D9djVI2MPz1CDYsRD0NIYdDqlqntjTA+Vq
IiQjF56AiGaVWbG3DalIa4Hkk3PYTPNwM4kedJIp7XJn+HlLVRNIAeGlSTPj/slG
D4Zppsm77Q30VESqDyNrXwqOzc/9+6/Lp3u/ASklGwcffbHNI95sdRGuD3o3fWH6
bqrRBnWtNNpYFA9h3mckbhX0lY1+OaS5TCytU3l2XEwGEH4+IJIfoSX02Mfox4CP
YkCDPS3pttcgIMM6nZCx3Cjc/0/nOFnKNIgAEgnqrN8angIK2ajcRE4grKGDX3GW
peFhU35HC5C5eukb6MZhremNHBH1ipRF0hO2/wFjRaPmvsbBtv6GFnStPV4QrhJQ
siPyudDcq6oOnM+pwbGzDOp9xEv5w0bFzVshZkzJF3kyEtJDAMnXGpE493hYCzZb
KsgyPIJHvAdJWX9xD4zBvZ05NEKfLZYwuJVBbwcVc7oDSQno5NTr6xYtdXZNaY1S
iGyBGYhgGG5rOe54My9ifszETfENkdtfinHTFyFvdLxA+Qt1IA1GXme1sI/AXMXW
+SjyiwG9cPIB4tbxqIhoAmZKiO4oKlkaDn0UAPvAditB7Y2M6jnwEvbIWkP5jYP4
xBK39mGksOnv5RudssiV9MHOat8I28J9HTVlMtZAOPA4seLp0b/2TerQOfk6T1S9
jzvBJnUsa7+vKPqZTnMknQ8yzF/RjZWFO6wMSyDLwB7RmMSENv4VdQBGOjhbwUxu
t+MpzZBlAUBZqbGyAmype5tUbC/2DI3vNL9/6+ZEBBpP/siLUZNEN2FxpqTjZA03
M2Pwt2vCiKtjlKoaJmaqGIdJTcESClC/8bsl+c+NZfd/pDStVLu3OdxhEDMaLmfR
Qb37xgD71r6W0FeURuN1+HY9xPhjrezYAc5S2UKIZu9dVY8lt+QTjKA3USy4NIG5
l4jo2AvziV1qR9uabmb6k5DYPRgdugQmY2NL25uJ199dHcz2tvihSP1YRi3YarNs
INcPP8ghE0KzyKcXKb4wG1E0PcK8lW0KulwBqMh79hcX40JEj8XthoHlNPitjRBx
zI94mRNk+hXmYub/f9E7NlV4XehC76g6BK+bszPnVGskZiYx9Y1S7/ZNdcnh5/Av
38FaPRKQIKe9ulV/ubjh8/cP5BqH5YpbNxdXqL4jV8wFyF6jtZ64luLEYjflOlAT
Wc93og7VOYB6Izak3EkcmiD+txBS1BIxId69P1z9Zqao8MIutFi2Qxxu2OAxks4b
dQoRh26hjD4TP+H0Yy+ZOXfcIOk5OFtx9TmRjyy0wbejsZS+HfTEUWHFCFDvx2lZ
mZnXlpsO7UgfqPB7EfsqWnJm6XFgdPQDJo8FOxIStmsBgu3nUuTJLBQn1L1vjol4
ZsXLHo1csu1hU0o894GeQfkdh6HWgHY4eJOE1XCwrSjlUcDOMsojtDqjFAA1Lrvd
QS6n/1c3ZeWBd2QS9vIxWjC2bY3yfZxBJyacaWsR/5RcKA/EgxDEQTTKLvCUsgr+
oP+FnByN81PTVUrUdjT1kqWxHPBkqXSS7H+pdYl/oAA8TevFc/BF/6ElLAIDrFd/
dQ71EwgLWRvT9TRaYSmWhJKbeoGqZ5sOl7KnA/fItkDhdW5qrBW4zHSWIXKF46xQ
ftJR1FJ1D0wbBENJQz8Nrai2dPfefzoL+ZGRlXbsS9cV2S36XIQ/1AdXpMU9mO1X
nZgJNINVW1g5/YxIhimF7Dz+U2ttJuJxto+Ujm3J495Gq4vLIAz8K4Gq4FUkGzH2
WVfB4WaqxUKY+wcYZJAUvX/rTCmkcpcsu7oa29naH4SFzVzWwGRdUmNiuEMpEQxH
0bT5OSsM0D3GJP5v3rBXiV1EHgA4MQ4r56v8qbbiYLGohqKjbgSl6fzglA+hTLhI
pv9y+RRfe49unj5blaDMOvZ7cxC95cXjUSS3fbTy3DAk4P6yvamO33ZOjRQrG5HP
m0qnAZVUSNARxR/LZwI+Xkd7SO9uuIfqc4mrMqkO+SIy2mxP6mE2ljoPVome9PWL
7KKS9CfbLIxj6d5bAks7eumwjzcmcdazRdkSZGn+p2N6zUwqIGYsRU/cN5nlpsEj
YiZIctMbLofM8un6S9fWvBkrDMHZzd9Ef7itjElozXxNdgqxlRFGYvBQiDxF2qvc
0ZJv76knN4fXExl42fVZr4TNpNpBrnN41ykqzxL1eYGUceNe0+arZntDHWSO3X+V
prvKbE5HDdfso99o4T5aNQMu1zPZXgrDADWbr05BPuSlzgaIyx2MbD/HkloVsWRX
Ryt7AmvJ+D7rI4Zc/fEk9dnmH2jIjqWl7wBZaQ8OPv89r1qliJZGZ8OO+RjKRNds
lK65uxDwke0VT6KNmxyAuZDT7qiBXtaI5fNe7NqerjDv5pAnl8lK0Uk/5+vt35Fz
rvwUecuDRznXNhUicsFuPrUPtPp50c4WFC/DlU3lxIhp+zNIsGtdREAbGFMrc6nH
uLoONy0+uVBymYtKFwMjHwHH/FNXJPvuG03245cBqL58L7YYR6VCgEi9P52pySG1
FW6cKa9wCOTHMs8l6IW4YOvSPymO0wDp+CfaELZnQwhuMfJr43HvzkAMvQ4c47PR
MEVu08lI+8fc+UxkTNal/MvkVXcf7bYNz9dpyJiWL3bdWiy0R9NQIayFobbvb0gB
dNFMTSOvuk9hY/Hgbcpd+QQOdUw0SSeoFr57UMJIOz4IA0nl33GSFEHXwz/BmRri
LL9US1j7nv7G4sspEKtxTF5HREPy9NVVuWMSmUAj0eRIf6eyzJrCiJotThhr66wX
LX8seWNK6u73TPwM3SzD5q0aESBFrsq2fixLK12E8Ghu74K+apJnKGdbcTdPQyYd
7z7yM3+WS4ZBTX1kg1KFRSsUwUxogSB/vi9vztXZpHzACV83tGCwtVFTaOiFXoD1
OgyDQjxAx6FLCpw0c804wJfmTN21B6dSrZ8/4W8qwCRLVcG+BNMOJFic9zwVLE0R
rjVRa0MGpuehIaFrJNkaUxn4/O5VTYtK1NO90b4GeHACYA1SEfnUspgFitSdEEkn
ZRG9+Us5jHwUTZmOpcfPmgjMAC4Pidol3YqJawUTCAstGUle41xmz75W/HT3ewg4
NQoxqAjkmwxVHvc+XJMJie3iSjusPgUoGx6vNeEOlyViXsZrtoKQIQE2GPjE6iBE
YtcVXfY+1HN8TOjSYAvM+nP3eAEoJotIZuvkRajvOapJkLgk2+N6STmxeZAaBQVa
BN0Zale3XC8ofQv8M/HQfDwgjcN333snN5nkcmpUVvsJuviC4DsArZEuSktr9nI3
696U1kMRo30lYG4JK4RuD4Zu9MISs3HgxGILBxsv2WDgKrqZRb80Ndw3LbVpd1zm
Pb4uBolbiXx1HpoJiUSIWbmBzdPX9Ks6SA5sxIjO7QvvDeoV9Mhvu1HjjYBQZfGe
c2oIdccu4ia/o7OQPNu6h7xtR9oiB5QP55EzA+C3HaOcBiyhmvc4v/QwCI4HAMmQ
9HVHf9D2UousgJeoYNASd2WAVznM9fpUhBP63K/w9+hSJ8j4ireVuYuv2vwhD6fj
gkyLwQhG8j2jyCTuH86JqDaMISakysMA6uAP7GOUkK/Y37PCSIk1D854ak0pE5gY
jQLdYacum4MADPU1oNzBNKxuWQUAjEZ9IVlAtt0Z0DjyfNSsLowzI02LB6DKoOjn
vefGZQRtPNGum7WBlPN5ngCR8XW6m0lqwEet+QTWG2xidv6y9GTypb5c9ZuZUBMV
f6zGQi0eADLJkBRnE8VE2Vs2+S5nsoWoWCzq044ecV5aGbBzibfSM0+XYDE0MudG
CBrrRqkb3dJ/YLsoCdO6xjiwRKQOSbdiegognWt0Dc4MQ8i0qoU81QwuexVtoHgn
2lBc0yeWsSdheGVZn1iA6qTe8HjRzs7RLj72klY0iY2F2ZOMOujUPxVXqLUozUBS
yWrx7oZkB7BO9Cg9D1V7eRacG63uh+METUiuqVMV3JmY7MedeSg4R1h6hN3axAJH
pcMlGSp9YuIxOf8RVsVV6eVda52dZ3zexF/x2Eq18kKBhj9Du+FIdl+S7YkF15qz
h75oWe1M7XZfPAZJhVI3Sb1gzGkMCc+stufX7aC3mZHA8j2kYl3MqOsQJj3urGMe
ImwKApdB67WGpW8yIMqYFUwNGjgBDxBSw0gJPFQCDTKPbqamZvqFNDCWp986P2DN
EGXhyjIhIuuKVKpecxmcc33+oMJkN9gGWH6uShWtmZsAAKvYvH2UWCbTNMiPwZB9
TSMsmbR6D+NTg+l/fcnmu6uy6/y/T3ytnydJ63uQwIs5P3XVfnLi13RLTFMKPNhf
DI/VZr8B4+Y9ba0YILDgJMx3HtEXWYtuCMHV1/xq8+IGzahd12rYaxrPzyjf8H4c
KeKBoyrbOsu8Fexb08iKkecAtg4BQ50I0ACMajGeghtGT4cDPeVlYLj8WqJQtRAG
ogGXHUYWp3jpy7fm1sgsGyHdaWZHMt/QZDRRxSPLJhrSNHcMFEYCcg0DPNDqJhJz
qAsJJMBmC6Fly2MLPa7tgzwToOIu7kuIAPivdVWhfs+Vdx/libD+ZquJ4chq6Sqc
Hrb4TRI7LziNVzp0Likg80qRS5dIN9+IzITMbyUMPVcU/tymV5USjaVDFiBqVSCQ
qnos0s6WoH6H5jSP1X+ookII+DoiKbJjF/QuIXW2RPd85piPCnk2Km2A6h1yarql
0Ha9V7zkIxzuhE9OeEEPGDso2AFVWBEC5IUgcpxMKgwA3xOacJqkJHDgxmCLn5n+
772Vn/SMnPIv2RAfEBiw0IY5/eteA+syh/FevZiw0q1lHsN9J6JSEL3L8wIpj1a9
47PogULR4ub9ysm8CTCL+1TOC7ggQLlGjnD3YFkXH2nhJOixvPua3WCfpjWD2PI5
j9+/EfyuwSpViMfyF/sWWUmRPdyU0vodfA7/l88a1vYPB8qSYbI9C80d6m1nOW2h
yV1kqzIJtcGF3Sh5qsJi02/NOZg0254PohXHQBicxEyAe7xJdsd9zOTkPUuRqHzM
BHkOVTPI2Jp66Lce4gHys9tgxCcbt2iCaZqRgFO/Gc+5Tqo8v9fmgT0yClLAbMTU
08P3sFeBO1Vj85Ihgk40ODS56dgIbG/mMCgYjkDlS9fpf9uCBWyP8pd7Xorq9NdV
96p9+IRW+xnCv3AJdHeot2QMTtXyaqYb1D2cdeaw3JZTJZ3Shu1X2OOdL4j1DXSH
0cv6XN4QiryNKaNxTVf5KOO43S2ceRcW7GcTDmUxllBlq6beWDjaN8mEKhM5ZA5j
zyozCORRnv2ATAxG+C0uTIo6KyJVO+GxEcqnb5UzllhStrwgSgyWMS3gqC67hJHE
Ic1oXpy++flmJxEvlSkC0mcjwX5k5Qi1ufgSmavREkiOrrT84iUNuEmqZctqvEE+
7iAcKhVqV1wPXGsgDMkTjRNALses88QjwzQ9rUuuW1lECCU1e2Pb6FLTeecA50z/
A83Qs4nCbdq+98CNzqZKimXGi4Se+Tl8FVw1i22lxLnR3R7V/eNjwHKKdNWtHjW+
83lCAlqkbtKXHn/KKsnFmJOi3TjjQ3xQdWeOOzIp2nL1z56lHHlGjYRo5F727X6i
TPVJZQBJDgX3ryno5a7lcJjugGZ7NVAkNUdsePvZbyHTbjTW5O/ywMBxZZyq/Dzi
cIArw2lC17dlTJxoY2Wb4JJKTOCX8yu2nqjaGyiscKhcZrlIIFJAKO9r0zBnxMbA
bVgGSzfSsftoiWjely4CELNrZR0a+4LyjvCLLDyG9tSpYNrcAApBPAAp8uQGA+yp
Ud7iD3aHvuFapKrN3jTWavs5JuZ3tqksHiPu4XbgVdiOhtGAv/Ik/Ik3JsYjdwGY
7olJ+QSlVpO2/97mo8Hwm6/U5hN1gN8qJEBtfRdz7XROyz99ytvo+cZq1IV9ATJd
Un0KVS6l1Gp9gHa0Xk58gIWo5SZQafAawi761F/yfMcc+I5msbM33QmnoZOIR+Zz
OQ+xrB0hEzJkLWvbNr/CCQ5LflPaIN61bGhflKoFiBWtuTLM4e+bc4+sg0oRb50G
3JzO6CtLT1SNCqYsoZhGvrjEzAcjeYvUqneynwEIywGwg6nSHL3DIKAgt2fW92+Y
a9rKZe39juuHDLpJAY9NzwK5+eefhb6gP7Az54rvmWMdrk2zgAHxP1ds02G834BL
e+pQjVAMBkofZRbt+ntoFt5ppBTBURn/MDW8jzRujfc9uRH77nSVJPaRgf7Bf+3S
yvwa9nLxTTpLStpHQ9FoWEWziznRhhuq09cz8fNpL7cNuEe9aBxsoNsLGvhEO1J1
Zwx3WeNc9njSIhvjisTxK3L6R6pVeRA5Mr0sybKKTCQmnkUQl4ZxuVPKi6/eNKo5
yi9cCBeDTOyjtE0owCppPthD25ZevxkU2jx6v7r85EnNwpiZeveAC02HX6U4kq7F
W9awDA7vr3qyywLX5I1gWPsVNBG3IGkK7h8ijqokJQO/W9tc+GzrBN3ZuKCM5H1W
HQJllBNfkgYM5mfkwA5w332drqLlpTJbTpE2n40WiFPT1jGPqBb1P0CtzOfH0Az9
ll/aQz7Mxn4FOOtTVRMtjZU1Y48QaLFwqzWnE0ZvNHoQUA+snr5nk4trHaTpNkB9
WsCpjGMfM9w5WGFOJqLSPSYwFkpXR73c+maXFAPeolmYHd+mFqdz1tP7HyfXbJcS
e5fA0U56AC/ySz2QSxhi3oOQePOScoEp9U6ZyNo8qAQggdcz+mcJNGWebRZw5wxI
MB4zJCoUy8yjYF2+cV+su9OiDbliEf0WhZ/EQ8qn51noczJn445sBjmOZnnFlA3g
IKpSgOFYTNY6mntcCYhN6GMwwKTk+9T+NMToPpoNZngeBHZpkrBJ9260te7eZxdq
MPzr2g68HSrY5ZKE00sdVuZJu5bRWE1+YmnriyMw6eDlQrFVExHdhdF/9UsHXA62
Xw9tHF41FhyslnUQJYOJifAhfZFSxuvCcuwq3rhfT5eDpMdNAc8dwCznt+N17OII
uE1/2byahDZOubq+zYE9OxSrmzXCSjJuwvPC3z9CpIwAb3ljY9z9oxteVEFKOP3U
4gRITU0uOtP4LKFKO/PTAd+vGoyp9RiRzjsNW6+dxbBNspB8rZWRYjA14hgKAwMo
ka9WHd4YNIaAH/3Qp4FPvnDzMWq8ikPu9K8eqgI0nihBJjm+aecye9GSbUEggVPz
nMbpS+wwEBacxl1Aj/uUBrIc1wKJngS638vApxhlZ0V0c9OSHxdEWOLKgjp7r7ct
mPyTTvlJp9mqaNLJKo+5lfnJYIikEOMKeHHCShsoTCewOtKx4citMWrRR1qgPtGX
6iS4gcVMT6Yyu7sQEJDPItnig8udT0kS/+I9+xQ65Tug+/7ZxUvO7rG/s2/UZc6c
p5izPjRY40xVs4v5iDrTXpZsf2Ja61iVz5mIU4nWefNbxr0uRA/NDyvUChcDo3/n
fePbrwfdkGdEb52bMQjxpBSmJ33GSR9OjRTpwG6oYDskpvpnm2xET/JlltGr5KUY
B+2Rjs6mWJnuinhUXQYaOIbFW5Xp29fGm3mp9dWsct4ED4UYQls/ZKk0sxftGu8t
xJiZT7b+PwAzwS9xPoC+PIYJArYBYOQD72Ee/yibzbJDF8y6rV/KJQNTlyMY/q/d
sHoZqazsf6GF0+vep+Z6l5M+iwA6i63Yy+xCARDIoIEmUNdOk9paeDoax7LCdOVY
jHaaeCg9AS9cZFp/hmCleJEJIISSgeQMT3swCZirBovZXjJ/yPv8Bs0QTxr+w9F5
3U00w2iDepI0JYMbZ0Qw2DlRE11NeJhs2nAvNK5kVWBFGg71Z45NxQLzxTST2Er5
PB7uAYJFGCeg8rQFd84hexXELvS9mmP3J1hSO7cvjBSHvl1gDEnHvSWWWMVb18Bv
m2amkRtxkFvbohS5a0Iw76ooEbv7bhSdyb94lIOfezihIJnlgjKFW56gy5m9qm1N
W1ABb7WOIME87ugH9VkdV2jozyfaYGz6HsKy8NadY5b35iY1b/83DHzVmAtilH3O
Nf4QPhcT3lVeboiaWWLoPJc+s/vmtyE3V0wNv8CDeexFK++kFDz2wzQB0ZZp70KT
CHJx+IxqJxA1WcVGj1k5zoehSEHE+ixImyLH7dQlK4Xq32cdwmrRpXFitK3PGw02
u7n1BnP11duxsIsOJoqd5HS0wG2Yo+1aPYRrpgphRRlUjeFQF+JK4AF5ol6/Syeq
/bFyy4BHBrjbjNYHt3rPzZMQGGHOthQ/f3ETp6W8R5UjS0BTEDjA4toEd2m4wqGy
iwkflSe0oUY99qabkMqBG9R2NpMOl47zaGEO2InS/8WmR4MfnRM1EB1TJfPVjG2i
j4ehbbYU7cLkE20rmxuSdpLbn+TAKR0XCttRemYOxc9XquDMSMZabu7kASz5JNaN
MwxZ07kwADyWgbijhTUq5P4LVPr6K2kGPrx91ykM6ERdZRHx1Qin2LXgiO2y57hE
n45bc5G+OTYQa04odhDaWXHdeCw/Htf+UtAm0ckzAjY50gm+lEFVowvjQxkcjLo4
Q7LDw0fpeHwuzp5RuAojhbtBsbl7DKMBGEu323EooKOz4uR5deCWszXaiBx6/cT8
ahL73CoOjctq/OFm9P2s0E/gCGQIYL+ZuMLWBI6xEHuPksnKVvVlVZ8H8f3pbekH
X+xcPNKqLSuc+tijUmlJ+Gwx5GnbFCJ/Fs7sKElhebBR37AqKzUJFI/xFttzX7ju
utc1YlNdsVu6WvnPIb8fT80LGYXDibHCYDaRVS5iZohwsHceYRRpNUzPv/JE5CVt
5hhVu/Z6+mpTAAh5saTzuz7JNoPTEs4YQbUK6pOwoYD/isaCIGRU6sC/1k85mhvW
H8S/2W/wQIZShknGkSmfhMRRs0cpHV1VD5WZRX0nalIqD5CSGultr1QGKQ9pLkkb
8js3iHn0DLhA36o75UMyEZj4EUb21YNjzfwehV2dMqiykAaTbBeg8LbcFnVRNvxJ
/KvLK5APbzkE6LIVR+tw/9xSuAsqaB498iLA9zNlExZMo3dlqGxmuSgmjBb5HB7i
RbS73guEWkw8y3zoI9Db/5/Wbz/1ecwAnsJ+grhjS7tsgaRaoZ+47NjPlCbuled0
89q9qZn5nJ1QY1yoDobyeehJuzOwuA5ur082vFnp2UJwtfvS87V8t61h4Bf2EdRM
a0Ut5YO/JOP36eHTX1oTunwLJ3EH/sZqAG+0rzxyi49L/G5Zb82P3rnI8HSQw1Og
3DzU0bOJTPysK0StqsR1XypN9gnloZt//zPWZtb0NFtpg68/mACZBu7d5XdetC50
Q7OskdljQ1fu9Qy2WVPS387LWL1s2J+dAWphYeEMgsdkZKrwK/OoevgafSqq5zy+
2kgz1TkoykgzRjlEnFbuPVnpY0iBhHhPhOmKD3BySu9U2cwOslF5dyMCrBeezbPc
dZsVcqE5h8Q33qYvDAaw33iIE7Xyi8JcP/ppfM+bqgpyE5p6zYKq4zXQeURE7XRw
8lNro9Ub34HMaMV1edPE2ZIvit6t45CZtLcSYqnFFMxsYwdIvzvc4g4iLchtv4Zo
pQxWl5X5kAlu+IAqIF1Z0ts7Hk3brY3UQsCSlKHHlufq+TbN4Jxy6GhXPw5gP5NS
deHYDULyV5l9Avy3/VL7olE2p37P6YjBpQLZ/92so16CtyPrBHSjy9qlEnJEPCe7
zOCBgdIqwnlnK3uWwptlxLedzMGspIxeSUBZYujSEeifawGxcuxpaw/AafyutyG8
khSW5zN40Hksvsyx4bxD09V1MmIr9Tbi22y+weRLlto85X2U98YmTm8niShhmz6n
TDempaZFCM7LggNPZO0XWzKetVb07CpBIWFINvYezQ8FlK9qPAyhAJ5cnJkFvTHc
PRDW5W/WgN82xn3EU57z41iDa8gRwarEcp93RiGgdAYvRVlu/PnlB9WSNl3nmWyw
A1YhDrcdErItfJhyAKStA4UVPAiFhpKA99V2y772nYojC3K9Or6tL5X/o9rGwlXI
GTNRybqFRc/3qGTEAGPuwyMbAvypiogxez/WMF6xs1Oks5Jy9ibwaRjbrc0UXGZA
qPZz/TbxtRC/3ggfdGvD5kDPJwUCkIe7c47qTG/Z6whm2cvZl1DCPFMvV5FFJ5/D
KJyHT0M9dIXzLLOefi+/m58gTbkHrznIsG+EHSsX4EY3H3Yjf+x27KX1NRZuSzsc
BwhbIaILHYdB0m4QpVQMXh0ClBas7bLlMr6SNNxXxcdGkcSNJcQALaohULPh6irL
P/793g1aOvxcBkI9mQCvrHZQ+aUOt5o7S6dAdnIZYlFy1Pq0aIDUZm1bTbnY80CU
R29Joj87btcsNd1hCO1+VbKf2bWAH6WRGRlHRJYCRL7EihDjuVyyhbTNhl4dFtQ2
8BPQKT4ajgWjse8OB4JIKIyKhwVKODqbgX6FsDjfvbFeOh4odpzFdTPVrFZrOsJd
YjvDxgkdf26FbmZNpvJMLBt9iUDL1HlIDe7oHqpgAWxdJ7aCeIuQbsYX7WSLmCgb
aGEPROGDqQtbq7HOIgYz0VGoJoTe7lVW3QQnx/Zc8qQ4glvQ3VIklLPUCYICD15w
dCjCUqy4kD+gG7qntkUO5QKogTDx0JpXejVGDuht1tWLiZJG+yF614mK9b8yD4HA
KUKlgQG6SkKHWQfq+uECzCxc1H9RZEN0o1SxaLkXjE8ASJUkm/kwQPqk7sBEjBmW
XZv9tFrXTMw6B6KDdU3EWabJJ0/Ov4xFCO9kmbjFk7sDuQL9mcbp2eMnYe1EIBls
W4g13d+pKgYJeiTvwBW7vS13jr8dgyH3DBus1F5ruMwET0MMngeeGL5+RSbdgbSG
GQ0gHWkfoNxDITYVphvScWLlqRV1Kk70SfW5Yxxevu6k6+/4Nbo4/MYV7/O6ycCr
Rw4UtnLh5cjLoqtsNIq+USMBkuLUj6iaRB/6uoahhzFYKX0ahVPZ5Z2kIljJS//b
5OegXBj65R4zka6ej+pdpoK7RUUBq9WTYJ0Nfmv1UTROiKwrIh4rLd4qDwVmstkU
xHdqYmPsMQ/yFKKReJ57htaveQOp+yZXfV0G05B0FQftZmynP3K/WgZyMO2OiCuA
zr4FL2jAgfKCvowQPswspZ9svlfcAHUPJjrDE09L8R8Caw/UCDtlkJ8WoXB2pdlF
hYKteySfI9wrVI+NOcDtOGI4OMj13v1IqfNLa6Te3jbYXNJLhLt0zrztx+oiew0I
4w1WTaur2fWkMjJHY/4OijlGTtgFQcumhrK4GUr6Zc+tmD40k087puWejqbm3NY5
GllgdzCOVRDEi9q0ThcYN06HK0zQY7r+Ny1vTCl8LzlUaohqfH3CSy/xyWIuwDRH
ikgYO+2WSMw9CW3hLf1rlRloO0xcRstNNxmgHxdBlyEe61SuiMtpQjLArgWBs5WI
/pvayTB9bI7QzQlDoVF0RU82cNmAOpqWaEIxdRdb8ucS4u/9vKC1XXnBdkeosheR
VetYPot00y4fZj/PIO6BRqXaWjkj99jaV8h17jQQkr2VRt6K+vG/vM5H+veH4av8
I8tAWSvR2+99Xpa/qmoRuXfDwGDbcSbx5o6spXlPUx2EIDE2cAodRPhxM9L/bnq4
Bmn021grNQgwsF64/ZYOUSr7CYNaEuPBaaTUYjMNuov5FH4dqCwu/c1i+/OPrelb
7FXyyWvSM15RZBCvq43NJuW3LNXCQgwymx7EqXXcEVgeurwrk5nP/cXecxVcNbkK
AHqnlqVX5ZyU83Xwg6QoOkZ5YmE/mzQNlgaqmf86i2J6onKwiPcrKClSk9oT9B2E
clJ0ap+XGlMPSJd8OzRCE99haWhPWr57vNtI7qUqoxieW/9GL9DPzUdmYN76mp1w
0dh1wVm423dQIBWDsttVLa5TEmKjPeUNrJ5/0wGSPs27IlNHyMPgliQ5Wb5b8cqV
g+TgZK4mqdaiizpSHALAircU8pliNFw2gChKurNvMq3ryEXlKta5fEghY/WCz6xg
PGBWKNqDcVjuSKp+KOonpRHsgKK05KQ3BTBK3NMyI2wWZJAsBxy/uvPj1DYYwed7
qFKsnjzYj0d2jEajqv9ONVqGgzcSgzfG6xvLqCSIN25TgDkvbunVnV648w0uP+gu
wbIASyR/Rdggh/aYEh4VdkEoCfmy8Zo2uWbw9j8DdjQ14/PC5RHAUKr8piroseZO
34/Hzz6SEYRqqDj7t0Dpwp0MJOKzRfx2nR5lLfeWWPuIgiAujNlqhZ1fbCYdCowM
RKJ4jrvDgiQg1SnPdpz584GbVaOy/XLhIL6E+nhZpl+y6hbdo7oQLUaj6J54pUWK
vHHmwP6P41jSgQsYXKYcYnwiXwRb5iFgRr2iYOLM3FahnHFmAMW2l32yugdDjb7j
hIOb3oPCfh+sIjDG2TA16dIJVSWqRo4diRJ5wv0kHrz0KXji5OMsWPsGG16O9+42
wxA1OaFNh4AAyw6tRhHLtiHIwUa5bhxyzdAL0cuMT2NGbFIu1orV7DPv7ySrmHlf
EYGAJuO8borUm8xU9Sxh5GTncMmyL4G+4nqhqOR5vcZngisaZsZLOlEuZp+gXekH
XOeOxP2ptA5IUz7SveSrWHaOf7Fe0a6CKwyn3+turlEmW4NZ8+Gu9O5JwcpyGQ8g
4Cx+8e+zBe9e0+YEE+p6ilYHoj1JuCAT1zUmT1gtJFvMszMn8ThUoX0OB0lAlD7C
Ch2SFIocq9dPRYqP+oFcEUjzgw10vcyYwiE+nqPeB/3Lz7XOgPWnBN5XuWu+h7DW
GwxQv6R4izb1VuHlXgg94V9FPRmFKza536P7NnTWUF2FpZR2D4FVzDEVL6C0tCyj
5l/s8GLUkXP8fImB8Cawyy8F1UOZvQTS5xzqfmzAZCB/ykCQv+u9Cf0j4eyv/8iX
J1pkpL2s7woxKuzlH/oa7LJf5T96te8R3caQw+LL26s2Gn2kbePYKufU/1FCZcq6
Azu92Ezgk0LtUEtelgc1PzBqZI+dnKyWcLNM8gzfhfor7wSGD7Ox/j/HgcN3djUJ
Y4TFl2yHBr9twC4UZAOtN7+pMWulAZyEj4UqiJii63xw4c9cDn6nFP3aY/nOhWeo
fAQdd3WPuXmsCYSq4l6mrUFaw2TtvGv0/RiX/t67OqGBLgMfrvk4jr8oC5ywk+2N
1GRWyMkN327nf696HStznq8f+kwGTMTWgRmiKO2XnMraRlHwsjfZYOXXF8Qz2FRa
HW6dQZyGmhKP46DNZMZNOqegyyg7U17pync8TGNfg4wibq0V4v89tYNYwh7RSo+o
HRvSuJ4Yxnu9c8Lv0ly0wVx1mppHqU2UD/ph+lyU3x8Wpkupax1Tf4qumHJZnoi3
RApJV6LtPzNTF3f8DOEcO0s/w1cwIelhQT0skvqzegDFuGzzF+8o4oSUPINz5VMe
NfLbFrN2ZdjOfaLrM+1jmtFqoYA4XPwafoM4uQVKij2YODLz9EmS/olysvMibcsP
U/rgtWmfH0AV0D1IvMW4w9c+CbU1OF9XFeY6Fx41kNNNuyDUXNkIXDTnf/9DUOtd
PeOT4xVm4xtGDsa/iQMYebtAsIJMeprEeKBMa16og8OfLVixjubutBx1hdhBd1g7
xiy+uGMiiTmCqYwFhRbxBrIKebtuwUvr9zMZZ5nZ2/TNTVGLNqOuxIzbc39IY418
TbNxpcqc9+p+kys+a3UJGRhxPhdb7TuEeqTIwchoAyHNHjVN+99eoCcGJ6YRA41t
de4wHiosrCK1fUC/mm2++uDaWyptg2rn/vfWqGkjAlW2NWrWuCZN+3RxNqF6ICzs
SPlRoYBl4e/OuCXRlZyUPAGMBJFVtmI5wl9BLLx5ddr6OF6IRRayfej4wY+Pl2ib
BlynrnUfPRYDxv9lbnC0imrT80KHTZOJOHFwMHOtclrBlEn9/Xy7J+GRnYu7BxRi
yePXQX0pQ0u3FFXe4Bk5PLhFzSyUUJcYgFYm/cjBL9Fw52eNdap1PxqCgS+O9SDp
5TgfIE3zk8Us6LeGKzrVe4gR6JKuVEZrYXpduDNaL9XnvZKbEUYDw9d4bJiWsCHP
hG0aSBKXAPmjSjfTB6p77wY9qw6PxdR/fLCeL6xfJr3chTi1SlE23wtPM09rUn27
BuG6MZ1mm3sckmoQXoes4hHwIHNtp0kOWb5kzdsAq1zePmQ0AdlrqjKncKOQJtYP
R5gw6oErdB94TUElLiHx0cJIpQcfB3wM3RGWR98WOQoCdpLmQpxYnTbFAQwYOcAf
nS34Mvw5BL8qoy3ikpCx7fL7w0vUvhSNWTZAmtxOOlEkRlCpk2snhNbYZiPwVZd4
c10MsAqRE0P9d/POovScABULllYdonpZ61PPXInmg+LU35vI9lF2Yevs1cj+imWh
5dE4EX6SPBGmmsz+B5meIe43xz9dtBtDHuYVH7BIKAu6GIiyZUSWaNEolK2pPNS/
ETWE/5fTyDQytHGoHNZ0WBUXY3TyhRrx0j1u+CxPbqlZ+h+cfUgDPX3GojGV0Myn
1qcjbRGJR3bjHdf0FxQkDeyurlY88NAmCHB+9peDWukEif/9iaR3kYV0lTtb2eBk
BvaI2HAeVoMIVoMcJRyuuyU8ZzThmU3Ru9VZnDTKJWfKqKBVXhLs/jeBXIYrcDsX
JyChQa0xd+sNpMNSFV/tB4tAWbrTXmREGkDcdqWWvR7P0zptGMoNMD0earJZIRb/
r1yngPAIPsuXDVby0oBTMWtUYvHCJ1HLQKEDOdKTsxwrVc7BW133qVhS/b2L3fbP
cr9osC0/29gdjT2XwKWbOmVkJXabgiG2T9LDhejTRt0yQya7ERKINA703PibYNNb
6gmz4JWpGIPHhAbL0LgE2VH4Mq4groGhp5AJnE04kzccHpiWSroz8JLYek2fUrxV
wBAffKgJWMiR7+p0/wnThuZBGeEiGySqo8lZzq0DwITUBVD1bntaZvUJwsyR/dSA
b79aKCH/A/FN7Iq2TONeZjM0M6ZgxzVQulyk++J1bZdBwE4B0apDrH9jZdmbAMbp
yD8bqlcCQtXRHroXakArVINiCZBjmHLBt7tRCbeunYp/qV06gf+JFNG28sW0/czA
QTdyVgFm9RNVsMsULFhelZIxs5KwTke5stFl8SV3sl/jLHcLXz/k+zUXpEDNDxIT
4AtNDZdGMZMiOaLLxbJqINW/y2YKXPeRpXcrLv2pqIvMCCKsHsQJJ4VoZ5LHEuK9
wE7ZhrDjf3wjSbIYQKusznawLNpZA8yxAChMBhOj5fvtKg49l4OZG0oVIAq3pfpR
A8sOugydt7TgxmXlLw/S1LSAKMlh9NbYbgR0llTHBv2YZ1TvYbdDUGckhGVMdByc
WoGc1SuLjtGwyud+B5nagQ+fseKBWICjEz5nY2wteE0BAsau9yzSz12TlqRNQMI3
mOjHNul4ev/8yebCQTEjPeLA2xJXGaIOpy8xXorEpRaSQFzq63u2lkEk3K+Ul7e/
r5+iyPv/26P3fwDp+aClNVbqG6F7j6bGn4QRp7LXClu13E7iD81DbaKOnoGcOuUG
LPlEJ7NG3O0XL2KgSzEsqQDuVsSxttBV7+2JhzF5+7cyZW8foNUQLB/WcxcXwNE3
n9wP686B5ioIfwVbE5BsxwViph/1OWKODwNpHyhxoEbRizB6KvD/OFbDFeH9qSKF
fGyQye6ZZgilV1mPncPg7D4lpLMdliHJtpPFYw4Tp2HfgybmumetoR8BX9ElwNvA
y5os+QsVtkIZGuTb9yQFfRSsSSuhnCdiSJHKz1KMV1v6kuG+3/FOjmRhsxNCv68S
z1gVL1bVi2iX+tz4TCGZACSqwVnN46lpRdGSHSYS+JJixQip1DvB3RsMjOHMUA5H
BVrkVl2EQhXfbfmOFuyEyE0l5pWPbTh1FHJSYkF0qIDvPEr8YkzsLIrwV0k7dv6J
0qZBh4vSGTv4Pq/ldzIE2cy3OzlNOZBVDDdfmjQ6yfM4wJ1IATe7zuvv18KqOupo
s3ocEKfYtPNbx+bOv4BixIgwdoNv2rhRHK6mzLjy29Q18kGx4yEJtYyrWWgjyGy+
tnKvZI/r/uTPFjH/cFGSMcEeQ48dRRiIZKv195lT1rI7M5uxiH92cxUn3bFfYfmG
BjBJpdp3l5IsZUZvb0h2FK8xpCerXSnKMhfifdj7VYiFi6fQu4finzvqiiAQEsfT
GZOj5pNZuIZGswKkGV8Q9c68Uk3oVTC9tYZjcktsZTH0Xz0luiVZWFLpeYL0UbLU
AgPkyA3AmG8OASk/22ru38bPmfT60ac5h/ZytchqTeqFLtSja5ls8JlfJVbjPknX
GM9lLGE1zOHd4H8UH23ApgzwcffxkBO0qR45i+M1Y4Cs9FZwg7unShWX5WHjYcf7
uHrK92U8wRbiZT0ueR7MXziGcdsuOWdkNH5KunHhogWpOK5ALg9X/L/urIRM33W3
fv6pldzHhkCuD1uaSTJ8QZJZUbMVCliSzsRP/hMYG2zwAyhvwQFgCflwqif/VQKD
BWQsAwESHXq1V3yaej0AZ9+5wbNzx/5D4lBMzeTZ+VAmsIRw/5ZbCiDdA00xrOW5
6OrBKpuAA8Fbwxs221GbMv6OtoZ7QXTrq9VtEu4m9TAQQKFEeMoVHzOamSgZmnwk
BNnU6Jef5CqL3bfVLjoJ+nu3+6THxLeYC1AelwTZOjcfdnqeFf14uooUZ5CzHrd1
TmQvZGJM+cHmOZmSzHwOmulfTx3pmVt6N1FjeoVQU2hxpqTocnp/4LeShGPBbPJq
8+3k4Oy3AZTlHDT3YesmwxejuotY6lJunbBNoX4nYZriGL0e/U6WX2I+CUouZ/67
d8bB3jbX8PnoJrDwFkeAF+uAKXcCH/rzIaOxyzXYo9xkFxIXPSaCjgS0PCk+Lt9r
FjzvCIvYROqNWNEBWgHBBRoZSYaxixlfffaa5mTAodGZxDmda7Ok7TLrDUyHGSYD
RONwBGuwXzqhha/L2RwByznIizqHwJ5zFoAfva3x/jTI42XnZmcH7qoWAeDtOAPi
ftKQ8LOTOgcV9wTKqej1L/6YZCWMAHaemCd6ZjQVGR/9iirzOwnQwsW8VibN8rk2
BonDJ86Rn6qf4jeZaoTyAnD881CEjLnGh6yzoX6GIU9EAm0KZIUrG79Cpq182Gcy
o6zZ/m2dsUIey4UA0H+c076/s9w0euqVjILmQ0l8atqIvsGnqsW5EqydrI6zDyHW
mXVhRmT6Io0JgiOnqDNQgpuajcGPudIqIs8hpzSbPlcyTflQXv6IQ1go1pnkLE/6
ocdFfqj+Cu3B09JgW034yPsNbzkq6gwUIADGv0P0XWNtw2ZiFXuoACp8Srl3S0C1
aOQVUPQ3BA8PzC8cg20Nd889MXFfdWO3a4+P4bObd4dgqlRq7jbXqGB8YZbmFYER
YQResA3aEjKXs9wUb//D1/sV/xJ9JmOv6qzl7n1DyC7BLa0GcCw8Qpw5kdPkmBGV
u6jN8sR4qbLwDrsaq3zLFwL0rs1RCACv+7tZ5Oe2MFou+1S2ELzU2l7IHtDlRyXB
k3jXoos8r2nfLwwi5C91sTYMhqRA3oaJMI2sNcJneHa3yCQxkchiyxnrZszvLePA
H2SopoWCsoJwIgf3hlF+5lxyw1OMYvN9OIehjaS26pIuL7iPbYmWO4ZlOoJ+xRl0
iNLhRQYXTktdzSmu6b2tUo/9iRLTIXLaKz//YQDa0Dm8v8OBZaVoQ1R+jZYlZlTW
wPZIcneEQCVaN+tW12YcuufLulAT7R5wkyk7C4/Rxyeu5CN44yYMkXqt1m7OQaFg
o89X/hlc+DnBUlSJ1r4O386q7FhCjBiEc2PVw8zMuiZ9qu9mzxloISnnXUsTqaHV
PqWP84tEAA94xED/yIlbD/148k2bjXia+e+4V8B3HIwt1pYWiMnp1pWqBw3rikOv
z8k3Dq1maI2/0n0SORGkqe+vCJACl/osV807D6u02iokBDtCZWLpcB3kTE4mT9vD
V3TROwwAf7wqCegQYYvPhXXySRYpMLjw5fF1mjkePWOgcgd2WRRDLiT5FK9swJC8
aDaoH3We+Jb6b+Zl3eHPIJeNJuE52tlu+iJxw+Yc6qpUSVnbbSDm/4p8crOzzBbS
wrVCOZ6pNg7reU/A0IluccdeZjstHXZqbPQwP18zVriTiRdQAduFpQrBrfa53F4H
1Ze//Fe6johKb+hgaqTSpZ+Z7fqwloDZNAIBKziXqc2ZC7QEvv8G7/fE8QTv/Dcf
f5eatgGzUY1oE+ZIx9WIxMK59rvH/Be77ITakA81JnD9bLWvtLjpWVieXAS51Usp
uT99V+iJ25Yyy7wvltJnFm+jgWzq257vUujSEcW44iy47g9yiEjc07JgEU+rCIyb
xyU9hXNBd5BB3P0BttDraz0BEy+jBhrFybTQDZ40vKgnH2oIFeExYGEnjUEX+UP3
glOU+jy+yYiTKGv/wAWLHxljBOCA/LAe2xRJK0elFmtNa5j8vMMS/bm4PMP5LFjU
vrRsvqPSlaAbk2s47u1jtotxSZO2XO+75daOeFXc8pOCoCteOy9/C3gwolKCDVje
nn1cmvykweQmzOuHC+SP5eHUrP0ek6iB1DxRGnpNlIMEHvUpLNO4yWv4RW1/AkEC
J4wUigtp1Vd85UgwuQlkkS4hDgULU05Xl8i3gvalFwFRlQAkZszG4t3Bs+NU6CEd
RAy3p0jsud8ZcYEei5Oy45WTZLTeAkCcsSe5OtywScysbz2B4XTu6NwV+F8gOLPt
io35AdJxncqov9fVHeKETfHFZ+gnmKS3D9jTr/lEyJrfWhPCSt9KNekXWXW/lSto
psIljM6KcLHh6sk2920/OXGrsXHnn9ShkQ6i8FX5asD9M6H+rMDE6q1Od1mMHnjM
k7QaFu/xqY1aEquYeoEAIfmz+OzsAEepce4v7iLmSd26zBXzmMFQ0DR/Dy1XcRpk
SxGYBlN2kGUPzxfwkIIRBKKLT2sUN3ScUB3wW3Ab9ROan8Vh/7OwNC/V2IUYMOWa
O17cB/3wdg8JWk46c2Qk7ahyVsuNtuuYLLivVEQxyyrBIHu6ZFjvcywj4DaZYlIW
iIOmCuj6rAHewUCW32bse6zpvsKAKfn0tA5mdDU1FB5KLMWfYied6L0ugQS8x3Qc
U4PaBphsHUgWbffhv+fcUvUgj3LJtGOPKaHn+L9eNLpVdSLBsGH7NmAFmQT840rH
lDvMFLFggxFCYWLRcdOESNzJkuSSnrHV466RodETOl4nv3XhveUkuCPhesUlfV6V
qecaGTtqeS7eGl9u89++MFAY0jxEeiqC/qYb8JT1UaqLETrKMOMG9jiuSLc1jIGg
siVap8ip5JIJ+nPqkZW+1R9e6+SzHRBAiVt9yZNSk/TxBIqPY1p4hNRnZ+GAEPFB
NRZPXdtUim/5g76QpZl+380ez4nz9lbfORbNSt1s4E/2EYZStzqMnx0WS1FLObKN
OOrrbBi5PonP9GTepJglkeA7tC1f67TzPY3nQkdjFYATrRwdAZwEB+7XyD2haPnX
vyYQyiy0izfxFUAwb/6jQAYLXEQ5NjfZ10S6PbMGRvB79t2eA0wSu9ivLcN0TVfc
AgdzLtmAA8p799xQwh1wbHNjoXItBrxaDbvWL0QQ93sBDBSzcwGHWwIm1n47SCMo
qlLbLtKfhGjvbw4fCJ/3V35OZ5/6kDjbqSRtGyESJIlMCEZKzI2TfCUFTAx6GUYz
6Ewzic+Ac5Ds6zYVhcJWzCqF79jck+KX+1iKeswR+aX23AJzY6FHURA3BV6Lw0Jr
UeKFczXMLPrulVnQuBUpk6LohfekjQZVXuuX8GDeDKQYX+H0wdjirpx8clDL0Ttl
ejY+wEMmL1wRWjvm8kCe2jGyUwiLkW9yob9Xnz7HIgeztMRGrM72XuZ1wSGtFt0s
jstIj0YyhQeCCy2xh9zbkybbSHLTkweXAxzcURoSkZRM2X58lKASpagQuvyKQBRe
6endzRVeaWFYOak8yuVostYUu8l0o3blRdrr7lZtT9ggSHcUSsntyXH2TVp8j7Ki
zaxmJo6lg3RxWhz7zyt+j2adddH+NsiOrQpwHGavB6jR+mYbrLSswlh9ML2CoETj
Q3oK9KQT3uvjx6c+4Q18LpZP2RWBBC+PzfmntUK8H+jutqJ6ZZ0g9a5rpD2B5qN0
aEaEk5/rBj88mgzTuQlWVGcbiHsA9ZVXgjb3tGPRWPBq0BzqAwSjcBqBtPmqj7Mo
0w6mB6vYLvp4thUAD/lvunyBjQf20QNTb+QT99VL8OWDiRtRFMXIAIc6qblaHuJK
IsVlF7oxn1lyRRbUT4+E0BNn8vTitdG+uSy6o3ZUiOFr55uNv3LfwlhmVXXk7Eo+
TLh8fQmWAxMy1d9PzDhM+xi5waU0aoe0T0ZTTzJydljnBGJ7rQUNb4tUsnz/SQkc
jO8M99C7/RnGsmTW7sjMIk3MmO0H31dpYfHDgOkX/NQFLwOgAPKbMXAy3mrkqw+P
xLipleB9h/fzasTa0b8PcOWkUFBDr+q5/N2ncmncYAMd/ns3LjPLUKNcnnQG0e6Q
JwWagipsy/9WNnnTUEFP1J92AnBfqozKxxDuIZdbFjW07ZvAMuQM2jHqvP1T2oz4
Pst8Mll3jnw9x4cqYE4FNXnsFZkSrrlUeb0Y5Qnau3/oIhyOF9RjoxZsNsKyskV7
d2CFUsUDQdkzKjZVmkhT+qF0m27flG9UNJeHJKiAj028/klu3fCoIWF8BMNWM4nD
xUeFryO1Uxllu0BALghmmK2UQomxz4DGhUy1aalDUARrBbqJ7RO9S9dYyXnqG33E
eLH2nDvRj8o4irlzTnOMmY/xGK7vcO2xuKrEHs+eZlXf510AvO64AjsA9zS6rsOV
3a6CfzCxg2m50fuXgMToO4YzN/Qw3uVK/+N7CckrpMC/dLMMQU4wm2eZpNuw0M5W
nra5m/c2bGRyL3naOg3Yw2PRo9ZG7EQHGPRUNPUiGhEyBZDvUb8gzYjnrBT+249r
ySn8BZb1/f078g+8kc626Idcy/pnVj2d3ULNnhBObPiQ39r2X4RqS51e5ablwuDp
CaLmWNQiNN+5eybunRYg1ZtiL3qvsu+qzu/lViQydvtNkLUm21iDxkM6aPqSfDd7
+2fB5GsoFFQ9pRrPItJc2uairu2X3Q6zEJtgxA1P0eekdGX2Eewl1ik7wJ+QzkJM
IMV+fkq4K+0d90fKvLgEQ5XzN9aD4J2ct8LHL+uSX+7n4DQLdfnyM1zN6xGnabJ5
E1xMAjDCiKNtxQWoJPuc79XDc0RhOdUQXYSV7j2LNY5Zl+9AW9Za/dV4p9UMJ5c9
WdEfu9gj5SCiglgAy3CISR0zQDu+ugVJaKy/QHyrdGzQMCbQ69fm+XQB/KI68dKB
JnMcy2qZ8CKWtBemIsL2niANr27w9ocmzqATDFJCbt2RJR+oMmNb8ottVyZ+yRTb
s4EudOtOd083pRNdyhInik+rB/OHZuaZ6MIHP2fg7SJsipIcLVdpHRHrceHFFcdA
Mo73xPScH7p0kXqr6m6YRnqZNHrbPFoWEC7Zoj2KGQsqI+mZlKacilJIxKgvxsOJ
T2niyBAFOLEsZwqCO0OASIt1KVswTcjQFc2jKOKfpcIwkBjlfPXAzYofEspyd5g1
phHi1O1wrVyhZp+losRacS5FyOwArf2vJY4PyqKIM6bM95R4MIJl4Tmg8I+r/9VY
YDRs9AWID82ngHqe5f9N03pMPCzTLv/Ub/ynbpFP3GnkQgbj6VqZ6X+AlE28jRng
3ws+/pXRXbTHtHV/Ou0FWpk6HFgu7wo+LwhnmN3+kIKsAEO+ZFpoXQuR1XJgUkow
F+1pdzPBPHE7DazLwLpM+xM5KZnhYM88kJQFv4krgr8mt68YQUvQH267pBKia7Fw
cUNcEAGUwCd/V8UG6IXd19jvztWGMVxx4pxS8Dsnwdvd1jzRuucWYaDwq/2h7guo
wBZ6IdeW7cVzwcfplPcvJ4gjS5IuYEeFCOrkl2yC7vG5yA46tznOaHP5077E5jjt
tNqOSKe5V3N8x3eLZUfWaQOK5bMNHUdzuHWCjguniTAKGxFKoRjnsyDPdePtFASg
Haaf0KOIjoiplngDviAdL/vbcOcw0Pkkc5ybnp+ddv8P7S7nKDjbRyaztDbanTER
0StMhUF0TPK+iARnmbRHMH36JZoHSnGZSrUhrFK7gA/N7YMEE6VCmDwLyL/iejkv
VU/jIUgShaG9baw1sFyA8jwegneESCuFByXlkE9PGTh8B6GRUypMrhd9wkFxyJ8m
IVnQQUUrcKQY2MXJEGEX0rw54d8YOf6DxvrfM7thEqzM9BxXMeR+V4lmCf48XW8U
Jj8GL9pQqNH/ijPmjn88dg+zxADAlNI00xIRCC4h/DRQGaTFJhejF/Qm2kshfjk7
pgY1UF15+0lDjb+qnXsqfd/ih+4MT2IpLo9s4fCv9Uj0nwvy4p3QPqC6KjiN0oW8
HEBJDTE0fb5CJKKrvwjEEtREsobwcmjRVIIn1BF/3+MiTqiuPsuF48+ehI6kVcMW
8/VU0NzchJnhKvMclaL9mksgvSeQ4ej7GgW2dDGbWiFyRXO3LSgpyDhD8uttstit
ui3x+dopBOtWC70SR5jB7xkBQdNAat0J2qr48HfwVc8CFs6fd5NAtte8eYD2TlYh
1NRQsVf54bIzw3I6yPWSQgZJXTLC3O7s/EB2XFniTlTPiLfo4ran8ubYI6RkEOj2
HmA4fPj2Ctmxr/6mvvchrqjZmCwqOiLmQKMCGlyJMJh4xdM6pAMFLPLKNegn+taI
1clGmGRiZQczMY722rhviTB4zJ9G+XCOXSghXSu2B1QBsiD8ZSuVSYaOHdA+1CTV
QB2k8KsL1eaiWNwHFpANFXH0PQPDlSy+e6g1M/tCYSmzUxrgZprRkhQoZZQ+nIUX
R/5keqBnz5ylA7oYn9e4CvBpO5PU5L6VjesQeiB9ghLQRQ/VSEXU/9arhEgt94Ol
JpKruZANz/3f0Mlk9mCNECCOtj1wYRlrsXbbmuxk0mBX57dZMoh56CHmTCLAAlav
pN37tbD1KVAdjpIaCq9tpSa8dQCwBZCI8t+juJJ+lgXkKI2vBbixRhD/6qzZySoV
xjluH4pGIt1HD7mtw9ZkmO/NDrj9AlwdQ1+cE0dRMhwgt0YX8RPVxN3AOn2OytZR
8BGJSC9n9QDWIFQi12Bk8HDikEtohepHNiFgkAtO7GjQTPrXPPJ3An5glwRHPayr
xX5wqMfMvz5cm3dALxZ1beNFCByNRBAiStOczheEL4pHA0Lnmf+6QsHNgigcUNrh
g81YlVsWj+zWTXlsZTvvsAuw9T9KtxueWiDN1mINc9tmZJS6Ioa/73ofQEANbw2B
xXRV6ArwH9In4MzNuTHeZoWocaB4rHw+kDGmZEWlEUhHXEMNQyrX+dHoOEQ6OOmH
KSKlctnMx6HbzFMZ/Vx5MgDvkpGU/VSjJgaECbo2WbNlVh0s17tP8rIMCq5437yZ
DKp8/elpn5P0FJW8MJzk1OPaobxREr7PzNA5QExltCMJ3BTe/HA0mKzjsm2y0nzD
DJW4my9AdH/wYCTqzRWo0fnYI/SA5MZV9RffhVLrmjD0A7CoEp2oIp8lzqX3+toH
paWnhyGEaTOR8bOAn5mujjZafAuosND8fSWg00vJn9+df8nxuO11VvfnWKwhRpii
R4w/ecpy8ZzMnGeALHp4fyIExbljlmGLfmyd10/GWd+q+i0yh4tkz4j+dIYb5w07
lbfH/LlTT35MCQGSKC5CvXW76b2PctJ+lZFGrpu1lBJ6gabEwbeOz09pS3TQ2Ulz
Rhszd4TZr5uxjvRzF/tdeHNteVeJhBS2eb5ENise+c3b37XDJFjtAOCP9Bc71REL
AdlRhWCvHhXTNcFTEOID+4yl+9ZPumPGgfBFb0kh8JdbHj4T+0k2yB6ImqGDIieT
fWrCtuJTaCSG2KT18v3xAGcyF48W2sLVLG0sdq87wgDbLVG43Oi1sD1YBdWeg+Pi
4bT9KzH3uD/Cazeb+MpHXt6mjNdffbVxhO+8Pyow1XAh4qZraFqynVjNsIgPsgnZ
ktv5tP69IHlYfovi93MpnoGyqVdANt6u+ttwSn3GWWUxLA/gRnyMEL3rTNRm2Lti
+6x30qkTRGg4WAonFM5fehDHJMPp+0js9Ey1hNE6AZH5rXCtuuxF2/D7nF0DEYL/
i6WvJVe+jl63TppEEsHtHgXJdZZnYl69wSFu4Q8eFu1HayOESr0/WoOHGBFTtOW3
wKmpoC2AxFYGy/nJOYoY+Ef/eF9OVM8ZFt/8NRCsNrztoeD63xb1NvX/vfNDM2d5
m14IQ9xqfl/jKe2uGfBjQ/tkdzfkhV2YgOge8xNgIY6wgtHQTHnrluXaS1eciWPp
0us1Bjp3TeXESO8AsNVegM342yYOIt02RVVl/LH+xH44ZsyyHlAl1TYtXWVJnSvZ
gUKdwav+nMLTuLqaaBFfIdSn9Q3VbzVJ/uG6vEXb8xcbtdmGkwVduXvjYpBHumle
E4mkyl01xTq4Rz7VWlK4VwT2Wqm1Lak/+32CKZvLehmK1fU15jNXEqkFAv7NbHxX
4FFiaIAPzGL/tj2g30hTH6uwAx30aPCYb1m8NkzGP/6F9KC51wtDtD4QQn+Ngx6s
NEY2JlWGvdnnstDbX8I/9YRxnep9eJ7+KP8VVnko5YUzixusCYA19qfDwkJjkBR/
auREHRZaNuOODFuY4Hh5bKZU9dTxrLKfe2NQKbkuuVoFtELIHu7eSmSBEecblD08
83zC+wGmfGzdmIhafNQeE9EPIo1+RZ2KusBB6J09KEWYe+EkqH1TC+GB1ofJbqJW
T+aq/LSL6aR6vIBJ0NvhAu5DmAxgqGljhP3ZoP1u11HKWyZvtr+kHVMKrJ9+bH2t
HXuDeUZn3QgDo8C/hXEpklP9XTAIi3COmtd+dRpOw/o/UvihYWOz37RPCfy7j4HZ
+DAE11hdrLOgcJHStkw5jYCWEFgkoiV2h5iy8T6eL7IP/eFU/U+2X+zrhoa+Vj2d
cmVG5x4D3+fZxRuQ54SQCa+8iC+wg0PyX5J9v8aZbm9dgp/z9S94HqzHF3X6eeiQ
XEXU4wZQuVgm9ikboxqY9LPmCaWn6RxhtYltZSuv9m8isveyR/zV+m/3AeOmCR/A
1Vgj6tJIHhov50gkkv8XN9XlaN7LuDCnQZGdwIT6BNtHrc3wJCs9NfbtVnwsrIHm
Pr9oaTFFphUNO7siUCB+Ktq7bsUe2dPy6c8gqP8CbyB3cRtPFigh5h+sNMwJKFck
cPzIxgj5uBVYS36D+mvWx3WoPTr8Yhp2Grt6y3ZJrbAYzi1RThGV7AnUCploHu0y
QLFKcvyKoo7J//qXmEys4CXjHo1g4Gh9K7sI/+ZcEDV2X7aL3l/uPTgRVnGCfacs
yyoJw1c3vai/fFZZDrzxNYJFBdcOOzVjyFRV6arcZs737D3n7ANncNZ1h3o9+uGd
W4Ojm5y9jaIL24XcAvZ456AhW7OWHioG30LXn4Y0jmNwvrEKpDKVfmEETlTw07PL
ot6Jzo03j1NrLMtKMOHne9ohfCjI8sFwnfvdLYDDiQlw7p9c4WlwYdWzBKSSObN6
VlnY0Onco7NVrL1LO+oNt+cg/goTOIa5FzX4T99VCvp9JAYF7lP7VYjXl82QQDMY
DI0Nrk849WYoXFXm3WlKhTa+Rl3ff/F4stzcY2qH14/t1AfJ5w/xSrBfWZ+3OFWg
heyGP1hXGEpTjfTK3iNAHX2cTRLuFgVN03m7OMTbqfTNK1lpfotLSO24x5rrLRXJ
bheY5imyslLJGhFAGYK+zdzqv5OdBtxj+6qMjiZ2MOw4IBvxZr8vCnQkKNfDawMj
KeVCtZXd2fbJuvMp+jk0qTxpwIopEDpGCevqLaDscFsq8ZRTy0YcvJQo+bKyrOng
RJLaYoztIVKILmxR6d4p+GtJeA+xA5G+Ka+9FIZSPPRWeE5XzfnKqwVezFrrteuI
byRxMO1uFhBBFGZxs1ev9Ef+CIrb5ppvBwQcRA2Gek320NFVYGbojdD6Gb8dPBPM
z605eZNqkAn7PnpZb0RrtVcTic3Fbp/chBLRjObccLVqDDMzSJ5UHgR5DEC+2EfE
2NOVdjSGlXCdD6+uHRHN2XWn9ZagbvMwvUV1ADvtdsa3J4h5OJP+sjl6KCwf/x7I
u+alN8PkMDZ7xDj0lCEVjIbvWebjYsvcE/KrLUjSNtlZzqFB/kp21NRxs9rw8pP3
NgaNhhHbQHGV2htl7XrGWpFvv/QbCBc3EfPTYoLYDWa1HunfE5zrHJyOecPIKFEp
1O7KF/0qcIY8Za1XckYepeftnJYvt8Q0OS8HKkUvlmCpynQlXlQ9q4GzY3vofgfd
3LHavjDqlwqj+xGICt3AbxSjBUMm7/xgp7RssphSOqxK9XdLqPlzlyUWBqeMctM/
nDBlrED4jqVEjSlMt3wqCGAioenkncs7Vvu4U0bLdhRex+jHyUd1KXHrHev7Bbcz
7+X7cwmqWrst3fLpBX/p9GNnRPAdo/ctj+JdmUHcKcQE7laZGH/DWGWIvccrh4mM
AClmVS6bXLaYq47R9TmfOK5jaefoAiIAS7P80hYrg+8MMaHROmbBRbroy82ymTz+
erMpyCA1FDehuBc6DhjewPsXTNnFXkvJXTKNO49BuH9bX7fo/Mb3vfMoSycq3Fgx
gZVxSR/A22VJemJgCLJWYwvnBmpIGItRq/JFgj0h1zEsiIYNatbjcAWOND2XMrfI
WBL3/XUUvbv2+w4mBqElGaxm+NhVEghQZWwEkViuz+3znEVei5IYaDxvNsk4DSYD
DZvnwBgs+7GnKuDg1Hg8SGllqxmTu310i/CYBm/Fr7CPDFvdBzuGiXJoL6BL0nHr
f7yHIgWqNQO2Fm6RcHE6t+U7VWg67VOwd6DlL06KAgE+c3OmjiZgYnWEnq//nF6X
oSway5onZ48zdTklLW3T9aeKhqeEZ6ITSj+evc76C1SPkDsXO9uT/UxD5GGs+mbf
AceLOdqxUT/kcvnVIZK/zdyKTdf1/poUeks3krxd9x5qw6Y48AwHSIwfX1/hpCQ1
zauQihXQXnsk6Sx5aPft6Nn0t7sJyzOlzQpZmDmVpTAhBwFwKpx3n0aDsSyWSRC7
aU0EhxVfY2UwQBRa8Jd8mJuKCyGhPXx4phXjLmdfdgicbB/Jxs7uJ2opefFKWCBc
/MI/QRlUuJhbT5aH5iUru59At3Lk62prug0yZ7725J0OcsqnGpWkR5Jp9TNvtO3W
txVb3KkZ5pjZjXZIc3yB//zjYJeLyhove8bG7juhF5xkz/fUidb4xdSE/jdLL+8p
shCiH9oLTJJyyM3doAHi6+z1rn85hmVpKplQ/5snsdsBnxJKxIEl6y+lGP48VPWo
A7ieymsQJR6oOh1R2f7NLbSow7FMhCyRIsqkJOkIpJ6gRQ5S4L0SlJ14ZHm51Yte
kEIbn8wALjc9e51gccfh3dXYUop5Np99rDVw98n2YgJ3BJ1O1NG2OCmfb7qqKdb4
nuGMm0s76ikPDUFL1PaR4jXPlyJIW6hGaUzY+Kt7IVGJJgYg6NVulbi67yfWnqBV
tgw8JQv01+Is/caxfmqY3u4dCbLCbrszgMKz1xf4hrrXkNnPqv+UlTq7hjqaJ2Ki
J5SD1SxecKHyF7xezSyMx4n4oMc6gzkk7i5We5DsyDmX0x7z82R3pCHTpcryyHxi
RhWnrF2smZBg9xgMI7hs33NpHDVLddMlrpdIvpiSqh7Ag/WJv3XH9NV48FI1jyDp
i8VLskOWm73mqKlkH8MHDcbgdVoqDTrlZlbwHOLEn1voA1zSO7SDz4u2d5ShURSR
KXdeXFYSuFJvoiWZvPnKJO/2wfA/MtppyOWTXUpZkPHsRv8LXZ3COIVX9ngCWD8l
KPyvKys6JsIu/qKBaolrY2uXwLRGWrMWa/jmHoybQZPme6uCQJOipJjqBuD+6wtK
T8PMCcy6GEtsSYE40UP22zmlW3LZPzJRfo1ED2V3KO8LWAAf+odrdu5eGs9H+PD5
aQ4SKhAIT3eGcMbHOXsEjCMKqPQoFDHitNMTLFxZsgotRInWwVRgWXbxLgN23YUL
MAUBYbBc9HTm/ByvTYXJq7Cqj+/cUgIuo3Pj5Mbi+ldla6v+dQknRzuwBlgJF5N5
kup+wHfCEVsmYGOHQbdBS1lvwj8mguspIF37ufUrMF4KEbq74agQZuBnsolmqt9T
gThydFzEF+aUuLUmbj2aR+R0Jwn2A/s5aq6wheswUFG4TOawGejzwkzddy1WXKNt
2aX0lJMaqimudS+V6vOz/FOwS5lv10jRTbJqs6YjDV6+12t2DOw8b1mSTuERWpHA
cClE7Cf9TgF/F9vaKtEZAKQ1M4FYc8iDjH5rgK4+Sl4ug7RJVGllq7fwBxKCysTv
KkK7dwcnE5Zsb7JBhnZRiCw5xDyvB5DQsGs0FaVzKegCNab93WJ42nTuqCCX0iN0
ZdgXFXXPtc2BxWMyVvBBBUevrR3huwNqt5TxavgmPtW7rJdpk9DwultArwUqyimo
K6uy8LRwWm+vXX12uLljuGDdFX4cPeTyAk7jO27w0xNOFayybYxY3O8JEkpk5j0x
N1JkSPhV9f5sNO23Cva8E9Ks1SQF38F/Zqbf/eg1DucYoJ5QO5FkJpz+tv/av+NB
kO96uKmiI9MwxXKHli6i3kn7mVD16h9iLfohiwiyV8v+Yn/jiPa0kfBssDN+1Iau
HNg4dVfciXTEW+Df04xOwu0VFI7MmLS86Zb5A8Zf1sFW60cN7Px0rABXIDd0106A
KsWR1wsGiWvV//6teTdXRqw6OsiqYkfLLQ59H4MAHnwREDAdk5ED2XY+w0QQawZm
DSFkYcrSZFI6Oarq/e0nJ02lRKqcK6eHbrZNYXwD3Bj363fhYn1mxtdOctULnWja
mxchXtFpaprhxPciKmmuPL2LfTNQRJM3L527hRxvHEc1bokCIPX9CAjYZEc6KOB6
HAJqIPtqrIh411pyssLOPSP+sbAstraV1wFNk+F+rjd9LqepWnhkizRysZo/ImIJ
rer0On8FQY/QU+CxdBE4yHtlzwjArkCoLa4vpEDCkCsffJ0xMzODHeGuB9CJoYcN
BFfPceIR9rzLOEwIHoNUAsqG5NPrNipsrS7k4qckBOOWsS9zYNtwnbyk2e2ylwgQ
T0azdm9G9LvUwE4dwkpjQTRRdZckX8fSmyakeGx5h9SCSLu6sF0W4nj5Fh7aUa1n
uyg/6CvZx/9S9CUBeMwBb+VRhB00txf427PvvmUzihbfUDnWBpTA/Y9/4LRUge0S
/iEAvSkax8eb5FS+J1bA6plA4OI0xz94+xmtMd8aCqOQpDxx63q5XOFGSRlKL/G0
GQVFGl5mpBsdXd7+3jDl/7qge/ubSZMEKGnljeyX8UrvR5AdhUvK2WX6TGqFyaqC
l2Ta9Hr4dsC9CiAQLGaGUP1GX7ZinqFRa9D9NUplCDZqBLv9JyoCwZUKY8cnA4op
MNneJFivqJIJUuT0Nm+yMwcIrXpz3//jqIAkhIKoMHGPx4J4W+WMeVLCUXUxxFWp
K3qTSvpDBoW1eoYzV2Ca/rzMnVbERi/SB8l8UHEkT1tjDqtr0kmyll8C5SX3WoRY
g25CE+0BG8Uqj/JFJmP54L2evzb5plzb5oGRLPO9jQ96eg9ixgDRxznnzuVPwp/R
m5V2OwwpuNPZQVv3X16KQNiqBz4LIB3bF6y46PpAiFJdQa8RE+O9A9NOxvurso/V
++baZqju3xbQEFRjvrPxFTYaeHNcI10FG55JmzrbCkj6cOBBGS2XYMXlZLLjqfgP
CPE0s/VZCbsx3BHm2kRz2PYRbOhUBNYshwgOqHuaQehDPrsBzlLndCQ4SunWPQp5
gZxO/sDWt6ooJSimTxVWUcEInp152U+BrgM372ZUi3yFdrWOMC/T6bUP+1pUsHkj
uuHFF//SBGCOjesbkvCVqoELok3B+Qguoyq/0MCoVtjec7Mm2mvSh+2Us70YYZ1j
z1FYy0Zc5UhHy3SDJB/R4ATKzyE1nJeRkO4xuOu6a7PPCFp2jxNAHpFSlS5ftJsC
erjwF68k0f554UwUlDto0YjZmHxZhCc9Sa38JZU2XEgkzwtfkqDGeQIN4CX3rJ66
qjON+udprQ/Y70wMZcTVvjddCYEQg59yeBLnHFHWTIiLviLOFee+QAtjiW1+x6O5
1BsJ18ueuy4v9AKfKkiPYIrsXMFUx2VpA+022uILjMt2GtUyAonx0Z+sXHV5dt08
x8p49QVN/loRYUSkCvK/kFSav6V9VTiga4AMPnCaaVuiZQ3B+hjEBZIvhCzJZP2+
w933O92AeZ5N5lrvM0wmnm3uN4Gwm5iZ+kRVgW4IoFSBOPcmuAOg1HbehJ9m/ymU
5DLWqcAwxZm/RuAmUrb2EDtX1OyKbduOhgvtIVbDS7LIyIapYAsODMyCh44SIAi+
aoMaOkYRdWicHlw8pH3GCMoHLaicxg1SpWEhSzQd7LyuRzg2WEHeMXmOuDYycfpW
xgXU3n8hxCDmMf4ZdSv56boTrFdndDsf0t7k8NT79iNWvDsi/PJ5NggmfCN8bKw1
7Y7bpOxgRzFVTqyDXlTNZaLhb3iaGFi/RW8ni8jGI2SV+V0I2Mk4K5B08z++xeJh
FWmdJ0kiAbbYWBXzE0NeJxCOjGK6XbQxoVsvUt28xd4LYLiNOojr5f7Ipjzz2h97
+sUKhf9Hab8XHe+Yo/ChkVLyNkWdiaRvtsfNTggvLcDRUMUP6b8WMVZZJluSkiVK
5+/Yb+gxe1XF/O5iuOkJXDFTRydtUAgXp907M6KnxRringCK/I/+fB7nU39TUQhW
wNfe/ZN8Nnyidllx3jDx39tCwjUEwpGAgM4IOtftpmU7NYpdu8cJQyGGZMUUR++b
/9D0bDEZ0zcApx/OixfNTws3ORGaaR5nif2P1Z90ZviFwq4bVurP85BcrN+4IQd4
A+eb8ZD6UbwsJ3zp4h5gTVTobYZ/tnf1NqkmUlzZFBI7kmyaye/z9uTPZlOCZTjN
OWmmLCfMNM/je3UCb5zDOwVjxvdWNOpK3x4K3F6ba+Xrz/ObIGtylLvrV7H4RtpW
PO784OyYcM8d+lQLAEi18+07NZfxx32t38ARiYW4oJJsyoLHD1IpB89/wbkpLpLp
SVB+Anv2kb1v6GSm2h0lXzBX6iaFwKfQz8lnQ+W+0lU9c5m9Abk1x13KKeG2k5Cx
qgmgq3HhH3t7RPu/t35VR1L9XdO1Yl21Oxud/pZg6AF/3DYOLnPapWqQX8csxt1G
+SQk0pTUWGDgl8L6mf+EeaP6x7qWrNgZWBdVgQs6Av9xAVI7/kzMVXKW+ShHsCRs
X5nLLA9W/z82/yRfOpPh7kP4B55M7M3hS9cto4evJRd2g5l0pzMqqwOqwahqL7sp
9FkXSILfsoOFq7c+8cGr8jAn25gyyD7kFVc9b4fKoJexU1S7vnpfM40WVrZNe6FA
4A9s0GpwCoGnWBAMJNJOM47JKy7C6YvpkBLJbQrVGr+eS0cm8oaZWHCvFgZAYyf8
8TwXVGPAi7s6EOI1FOo64XdjqGT2aCAPDX79JtCRZIs/CAfCSChhYUG9GqU/cAGM
EVQBffHRMUm5oDhvvq+vCuHL/MhY0hsDxT0O2CQ+uhkerJ8s0P5d1f11gKEA1tPy
p9sO/BMB+7r3W9uVOFLrmjKyLZoAZXaz7nxwta3fxDfnN0kc5ToxPN8+w0MbeI7V
fgBIsDaTphfco5uFgto0XFD7nAJrlgHOXlWK7MInQrwGH3+4fEywFt2ARArZkKgp
3VBkaEJ1z7LVplCUeaTLgfiB1zguM8rc5UcL2Z4Jzq4KSHwpGO0vczagkNcHZ0wL
zkwXATjsi10lr3jeM3bjWRgLaPyS8HMRcpwMJWkj1kh/cKoJZYPyCd4Q3gd8u3FN
EIOo6sRgvKE7Ru5fi5EdvqkjzBA9Xhhvh72V2lbnvU4Zqn+Z3jQ1SVemIM7qLEd6
XfkDx2Ze1tybVoAX4ItuyERule7hx050ipE6Qfysw1vT05u7Fu7/+U8gjHF8NcFP
TpOC+6+manj44vOVnSqFlmBKEM3Q5qpWkNvya+YUM6cE9FdbhKSBxrWhaz1IdeIy
W2Yw0uxy+0c72aUEwGFyZ/204beJ0Oy3AT32yBhlzA+WvJ74dG9xkd4X3Ip2mJBG
tyZLUGztELRZKcwsRsKU5NE9Ar532IgVIPZ7NAYt38oI06g1KThydnGBQn6U0XdA
PCk+QQL+Ynegl3E3igjvGsTD99m9ICGDTjP6ZM7TkebPkzVecvEYaJa0wSOIiXDJ
ttnpWFhgwmduIM5AbMe2JW281LG8PBbKGMjsABbgY0bq+6Lse6958BCxSvdWGGaD
dmK75KpAlt5EDSzX4HikVQFT1dzjflaWtH9eHSu7w1JnCdqpn9FbjVUTmdcITdXM
73CXiJKzZ28CpWofeeXrGy+lx5tJhyxY9q5Ea2r545p+aFK7CJpi99dQINUjGRNu
wDRggr2kset9NFAxoML8TgB4VYzuuemBm+J2i1GvBDXgZ2S4jQBBH1rlu7A3p7SI
0uoGiQWJSnV0/dUTPRuwv5A4MrL3LgfJPdsAEJ9t/q13CKRoJFi1p3GDf4j3ZO/2
PtSHmvcTGJY0BoMH4pTHIvhRzLQRdv2KzZjhoDyN2sbbi/8t0nqcSq5u1Nbm+WOS
g98HGbTSWZ/vFGm15m/vjWYlmLVIjnAUrnvCvMUsXA19lu1NUUJMshvhYmaoUSU/
Zg0l/9bgvpNQEuJDyRbS6wSF4gj7cuuk+CkMryqHW8A+Pdjdb/xFzgK7sP/Cg6/2
n6+FvjeNegl6uMo5J7/hcL3ogqV7pcXhBqoHdHnMUCZkBjmDooIVaC9teLioMnDn
riwbSZh9MckWrOt3BcC1rZgQL8OhN0LJQaIXrYRP6gzMKS40V524Hnb8b4BeSsNE
z2NL74+JlaFIfRJN+5Ye5SiQYSpDp37VS/QzUscZjq6iHWF2JiA8kd1iYOoJ81NG
2U40b/ew0uC5UAk9rxbrN3erylRzDvbmvjoAA7P1Jd/e1q1ewNibo1mxE6WTzHiw
GeiYGrLQaDadJynW/uO3BjrjmKULLVEGx9WnesLSK7g6lRpatywyUfmMDswE2DjM
6pOO4tZQgCB84v5NuuW0clKpL+DPrL3qQo90gHV2svRdnqV90uDF8qR9XvZYtf/I
StM+8ujMRACSCtfzEdpl23ydC9CnX3VdC8LLnOvx5pxzW9739gv4riolGS4k1RTf
lFRYahQMXZIoG6lY3957yZK1QW5A+w+msFnR7VdwUITVigyzm735BgbY6j6oX2vo
6+FFFPTkk5bG115hk+kSQLEWBDJmzdZqKRAUrt8p7ghBSmGcm3sBuPaVL/L5LrSS
/kENzKntaoxdvysi1yG3E+c3DEW3XeSx73ezCWg/h+OW0WVWYLGBccQAw5sq6Nka
q8zb2gpMuAA8jpBtIjl8iPC3WVBC9w7ataWwc8s92yuYuG67jlJ+dNoXvgF+SxkB
aIfJ1qMFwCL1e1JLJ9quwL6mp/80+AB0Wj4E5uICDup0SXvJSi3tycYK3kf4OzZM
ksuSaYmX1rAu7zRXpd0fJP1lk96bDZWfz9gkpaBuHKONjO3pEGMip+vS7OB6WYBV
NvkVFq9/InmSPGHAEFDH86Blxp7BzOLde9N7OTAe6qXuzMbHklINR3ODUwWd28gh
X10CLBe/KIQxEmHo9dIo5vmTLcYbmwueS0b75rOaG34sUhRYbcmMgqKqpyPDMroG
gzW+aQx0bdpzuFyFBty+22gKhpvgpZV2vEcib78l7RgeT8sQ8rOlRGuoXfXuZ34Z
qPwNntP0pdjMqhcdA8UQYO2cmlpnrk8adJJawYZn/4i3YL2JXwWMFtllbim4Nv2g
PbQBykR5JKruqtT8U+TB0NUVKrqU+mBPyJi/OGt4MMFUMcbs7plTGtpLAFO7owYy
qs0y1ZQs0uR2997fMDGKCHAL7f3Q30VHvbDyKIHPPV7xsEUHHsmsTZvhGg2tf2Vt
8sX3MEwFRn3Leu4fDHK76r6rJnUXSPQCaUgibUskEC1sgRrYyXstHIjvY16x4Cri
ocT6vftrV0CHKTJeium7F9ros7yvy7NkXkpK9SQoI7wsoWx7LOgPdd146Q3qF20l
F8SEj3MlbIapzw2QNwGqWXqVrv+3zxvTU9u3gWrPuyql3NAqYEo5zY9D+a2hbj/h
68xL1zT39W/jXYYDM/Y0/Nk0s4qtKv6dNH22f3D4hlWhgEr6vCmoBkeLvGjnGWo2
CZLXJerfnaBrmuPj/tE5HiSaxI2j9tVw0+BD1rrqvWYnvn/fgDf1af0i5ieJyLBL
gItga/s9+jRXZYpb8XRr8Ric+JsUVUXemMWcI4zfimmuNP1H8ysiVqH3J+TzMbH+
md/R9YgTrD2NYy2AqPJtC+9Z8RFepQncOb7rVs0+NWHP7YzpnD9nVvF7ftAnpF1K
i9ZYN357uDDdxC3pNg2ge/Hc33TDOWUMebF6ta6MGL7+y/XkCfUrh00+dRAOZmBn
RvM/emvoHNfLJ2r6UFABBOaM51N/s7YJd0zy62WZ00c3SfOH6Kzsn6Jvv4RqJtiw
Wkiu7LXiyRGu0C/oWykBXmks83/Rb7Gx4orb7vEsQOguJUbuOPl2yyOxq1BbXV4H
M3pjH5wuEb3z94b/IwaPblQU9/q/fEQS5MDWDN+ChmGhs4+zh5asWch20yVg/aBZ
7Py9EOzWjJ4a3QFzU04LGYR3v3IyeQSVtHYDWH0/+djQngrn+rZFLswNVMAzeAYw
MP4IzdGzftVdzlFuR6klyZd6r48z70jYUmFoZafGxo3MNBKvFilahySfVq8iNHi2
is5/EtLa0aKjCedfXa98EcFCWhWx8HQVLUdADtacjzBnUkEN37erQMvxU4pTCOCK
Be/RTPOH7UPpEP9XEZpnTm7uCFZAR24MM1pfJUteohI6ZMOMhbe+2wF771hA/Wll
plUDQjPxStL4pxjFZbeNwbp95coFmEkst2kWTCb6+v8FOxf3TSmQ0qhkbeweilg4
ADdtKxS5SHE8L1wTF+XOeHG1G+kewCOGFwsJgBqB1EqzB4A+Y+G9dOI9/ZY8K7Rf
EereXlHmkPMQUIlQamktVDxhRo5cv1nAclUKj23GHd2qmFRpDtkv70UuMBdVweb9
sylxxeCMKf6MeOxktA2OyVy1i01a4kDhgSpDHDVmLl0QzmXYnPsjLwsrpp4jYyL8
Iy1ywi5D04lqAUQaM+Xy9fmsYJ2/o4Kdqko+Eq8f8W4Kyrepb+mQRSkla73I6neS
pW/sLq0tgtEv56stL1EU5Qsb05m5PrCMDrslmgJ7SkKOFuEI8rXn6yEMzp7DSMp9
O9Vh42CHrIkIuJEAQ3O5TghvoCdH6/oGqL/0kWR5/4MHJTiaRBpFyqr6TqxB0h7c
DRSy2baXPbuBLDxFRI8ZNA5btEOaxeKeQ3OFR6v26hqRGNQFoK0GZaD695goklRL
g7vZg5/CMfijZ7TZnGgQidKE0tkUiG2GW0o5PFtRRY6xeme5dy1x7a0paMhkxdnA
yD0aWINKobLJE+f7bxlHg11FljnUlfsgRGzQVfW8AVYQSWsIRwvJlYFv8isfM/10
zdMnQurvM4ykTG1mvLOnCKTrerZMgZmK9MjXL32hERDjbMcnRFEpWSpArRyzqJup
BBC8UkVnWM4mOMlja/MM6vdIr3BZtdAy6IGgSYEgrHH3872ypEsCkw590I2bfjKt
rZcyN6WQ2wR9MXweK2lCKqPmYpb/BhVHkVet5+lR7z4W/QPJLNozsXrYGh+BdxbH
qyeTs5+uhrOEPskA2Ghdkh/RNm0JKVMzinJvTvaL/IA2f26QExj/MH+r50ypWbzJ
Nb/NGFT0N/VGBlGEO4yb463474isYaVuDjaVYFcGMz7WxLQbFa/kJlYQIEkXHxX1
JrKDuqca4hfZVZ41KYw/oGPF7a6VjqhYLLFfw8WBfxYB9TSUspeyOz3qPo+mD0cS
wWE5YOEgIWf4c6m+LclHxlC8fXkA7EEL58uBLpIND/UlahV5BxO/mBHAcr9KhnPJ
pwASsgwEi/xdTmNJQEnHAobK/ErwGJUFcK2U+/B7qH5Cn6i5wfknhMU6iOXDMukC
fwtP2UeeqVaj07fSIm+V366+vhvzW4acV2GbEb+BPiaGyjjEUIbidiDFTbV+Ba/Z
YAu67DSAAw1LXMA+apAjq7tuSyWIsuJpPhKKkhEG+pwQGQCZr4iuumHQNiEJkTdi
qs7yKN+w1CJdDPhPhhdmWgMmItFTovMuCfLrGprHthrgppunPs7XbXsD90Fa62jU
6d/4DcWyL61bwvdyp0GewG5+eOX274NsWn9lwxK6JWDvcp3t0Yk9bdeOkbG0hUmK
kBfBbZzCQ8IAszqqwZ+iwoyF/CKCjl5PjIwLNsTteh1HMkx1yQLI0niBve67+DcA
dXnusxygI90+M03ZvnbTPwnqx45YmMU3IMKhi5mz+GBdrpTun4lddBi7Sew1yEZq
22Qn34t2tugO4i+iYBcC5vySgvp7XPZJmP1q3so+m0JGfmtWqcWXQuNv1ITJsCCz
Ctdv0Gir+vF2QRFjhAohzB335QhRPfah/7Zqfv+N/sV9KZ4V39UDXOjwQVrnFpgp
QVREVMcZAQ+RsUnohseo/F+MHYLMQC0lbf7MT9I2cqpGHr199W84thusantRVx1z
wd0FwoNXyobyTHyqVQK9Y0zGkSmB5XfQYTHRJ0n/cqjN9Udw4yzk4hHk4DP3CLfM
ZjiUwnObMaV34MBWv7vtTxwNO7XINOVn0s8Vji7yXDO9BvMrWTzughXhgYW43wn1
BwuME/2aib5dN1plmGIqPjG7xxG7/gDgnOtbs412lmKrwHdlNS2w0MfZdK9Dqud8
R5lpb9DpN9Gg6y0TxocvdvLYfeG122VGYkkrpcaV6e09gu4cpJ9uiU/jfD3oyglJ
+bXEttNCMNyRLpwNJFFHSk+CsrmAWvNGWVSArctvBUreIMcrNDUsF5EVkC7X1EKh
mMxaZkpgWXD0Fqxl2kr9LjHK4cPu9MIK3LyFhCoYYGSQs3XAYu4VVMIRAi+o7VCj
opAr4mwrIG/O9X3Qz80JkUH3k6TG1+vmoUEq4iC1NS0VT1/bVMyq664OVcQg+4EF
lsEBpHlhgU8bcTEZcBW9ljRBAxBbhR7nIcOyEA9pGBjDp33YmcvMK8yc+fu68BSz
iZxd9SV8gSStKurVG+xz5ruzh/VAqHLkz/kmmwc2se6En870ezoIl2Zmmv1FpNZW
A6glpFYZvBUpZ0XghxzCFKpvmJF2nmgFYhKFHEkPjSpWX5T1/+S3vBg37IcoA8EJ
kA0VscR+/kOBUWr/dUPZgASQ6qVyg9LksYQNs2VzGgyJfVcgKgsveUN83oPp2Wq9
eK/VgF5vsjY2GaJ9loXiggXGjfs6WAJe/7YqUwNXEcAdTtL2+ElWiln2Eyuq+QQ/
f/tlj4ukidY/u+IZOZUHGanhMirWFR8yQgTzXZu0vXAl0H/KkQLFuTz/Aqejjpb3
IknablBhJNGERYnHXA/3V9VQjZP4FK5s40E6dfHJUsnt4yicNORMRvq13UjbNO7n
fgXHxdcJKdLeMr9ayjgBMRXrR+6NWFyvkdHDsaobMSBBrsZadib2fw/Mp7/LtQg1
u0FWoOplCnBFOTcIp4C1ZPBkrDp18C0eGPj7/5XhjNsRa5pKYVF8kgblntRmUWm1
sQ6DhQQR+nR/35inVO/UcKUPwyZythbkG4gTzjSYnBbj9/BJ/cv9JYB6A+43MdkR
H/OhJ+D+aUsDXTopumzCIDfa/y8tAD71F6J376sn0P5L8sZP6aV+YDHBtcCpIX6d
g8x79iht01r9Ow6mDBXqy0kHH3lh0FUMi9pfSvqwt+UWfHHKK22oG0SDmzus46tN
Neciu0VS/MRFi+3rJppiDgESK5/nQb2qGJcFdF0BEcKQzf2tuQGxDcskPhWm+k04
LahgGF5O7qsNWEPM34B0K5ydpUwOYG69T/FRO1RA//+X3FoMIaqPoq5nJbbUshxq
0nrKcrLB1Eo9V7fg/O966pUZVZuWbyaY52d5IcRljt6mZEifVy1/lFRQFv70A2+j
9pLpjR7dOwfkSaWy2jT1ac5euXQGFwT9SI9WoPaH7B5qCUbdMjupslLpVKA+M58R
y7TNnht0P/R7jdGsFilifrjCVzTxblU+KsAUsD0jGr6Wrn07ZN4dM78eBBtSkxcB
ec2STiVC22L0JEio17lhZuk6siwMih+EvEJjru9tSyPhztIALOYJWKFBnoG6lN4T
miZp40fhNL9z6gfHgxl4X6zj2f4vd0ETRSjgrtqOYvRfF7wUNWdOcaD4ZRIXP8co
GvDTvUAWHiw7XIMiRH1FlBc7/Ril5xHUizon8sz5YMq/ZJykuUh8a3pyMSrk+WVb
zILGxuGH0Hcr2+mAg0WWwqriIKEPp2/cF5EgU/x9Ak5yXa4lzcFThsuUKvxEf7Vy
/ryQlLNGDlitWw9WnLCaK9AhF4HM/QNFDKnJvka1+vWALEXV5fhZ57NM0voiM5Kj
aLKHyIgFUiZmsylS2Z1TgOMJEiWSmhSSNBajwfBxXtH2IgUrtO+EHIKLW1Q0H5s+
Jv/eaqNBJsWoTfg4avjvj10yF+nms1Iq6D3M9tsyi0Kj40XCNvBWte+OAIVCbReJ
Js01s8D5QShMc0Fea9UWcYChhv1OUw3+IHTmPvrNGX1/stbJY43yUxRSlDSEMK1V
6OXQKsCXwQ7xPZ4LEKsZiKRExylQN/1PvDEHHenNnvEWrr5OqN/oUpNFoSa5jGjb
ZK1jlH7MxTZG3dpCFxj91Mx8v2eHyvMTseZTbPXnJ/xraSREkJ+12hzkeJV2V7Ga
nUFEdrF9nw01OLbFMVdjwHKLmkAEt5hmb25HVAzWE5ahsfOmOfVHG7Qx9DNVUK9O
yDUX2fdNwoxrhIF/90+jSDZ4BpD4NnrAopphSWCtJI7pw5myozc2dNCkDIHOTACX
vDLlFElYAy2eYdgzDLsWq0mvvw+NosfpIjdIpoYSvIWA7K4gPZU4FH90p2DVyMKf
6y9ZtRLChIiTz30Hnv0YuMzAEKnD9KwtIO8kQDhtPvS0ORZ9RVtuve1EWB+YKa8m
YDVf4xUiV1FJ0D/rE9zf82udfyuUGkNXgLvhaDs7ttoTeYVQ15JcAwCi7NKXrtlP
kUOuhtgjoICbKaPGqK7WC81obJlp2WuP6QNETZ6ZAsbs7n+pmxn09u4xiXvTFR7J
AnfKdOS/OEzC32S7erK5GSpZxAEVckMC66LMmAiEdUZNEs3WWK7GN+Dl5mx4qM6o
Yg7yO5Xi7mOactVnQcbGGADHQXWQXQCL7xQkCks73AgzFPfDrMXs7A/D33PhTU7C
orKVMv0fKmb9c/Yp29UNkDQyToHXFQd0mciZ2/njTaObXZ8q8H1GaapQoPKK/+GG
w1+J7eY0V9TALgHgzRguvgvxdb2Q3VPkEqPIC905EacPAvCbBwvTyk+hgFoU+bYO
MpkEAQbn5HimPKKplXVNjtpFJKM5FuD7rHbLKgXUiAGDC9AoZBdRbHpak2rnwsk6
wKQo6nPKw1P/zm0S1REm5vpaFljfm7VuEHTVdPdjwVpQQFtaMPUwGrMKR66E5vV0
N4MMZviZPsjA560LVuFeeO7Zb5SHPtxc9iv3EwDAgiBPlIakfR1Is/4VS3g7Ga6u
XyGo+cnwuVpDjSUhOveV3Y7xFyHiVkiIBQmbKQMtsK7oTF8gH/dMDEDnKGpYR8Yj
c1I/sbwRaCiKUbbvkS+GY0D5mnq6h3bp2HgCFtiG8iXrdi93KQA9KX36QcCnAVeT
Y9gvJR1dCnptlWY+tVU6RUbJDuUEx5p1CL0ecNFlkTtkiuJ8hlo2FW1ozqjg/RLB
fbutT1O8uJ5a2xwApd1Ge4q8kOoUOXWOuq3Qdy5J/juDdgLS+yl7OGhH7FLT8XHr
l8p87zMN7abzQAIRUNLw/WPf57reJNQRQmDJ7koHlqG5brYDaunCVMw0dE4Xuenj
6SyhqWlqAf2Ad0ILLPQ233IH2TEnCjmF8VAhBQbpIsQsjNiAI4ZCa6PFOt79xYst
+zIbiCxaqrZRpKGpQZzNtnCGz+sTU+h6yBPqMiSeKLqsMkgS7VWYSP4v0q1OblZl
ZwfB4Znd9TXbaTmX2LwsiPKeTosjEbbOYB9cBntilVAGnUNrRLgkxlHIYGX6DeqF
L9WM1CorGo8LKDsg3Wi1WlG4jw2mmmrCk0FqBURISas/vWs8HGhZJZELBr1qTvLD
HZZGSue4cWj5rF1Sq1NXDy7YzVkP8VsrU9ocwbLsZw4GvvPpuRMqcpT6m1y+IzSI
P3ZYFp20BVDpUSTftBrLvYAITl52MLVpr7uIPHP+mceZZW/vx70RpuSV7V92GtN0
LH+dHlec/bvZt9xxJ4Mx9IkPAgzVyGXwDM+WwnteeCdEyqNhCfW2KyUx+1IS4Af1
FjBXyAX0p2o9T2y1ohavyyqCM+5DRoOfhvFxqs7VgE/lsEQ/yrEWfBk6DpE3/yrP
+hwR5xqRHX8up9Jzh+Fbh0TyUTmGa8/EO3ugQu4ub0o+bD+24qKBRkPK9ETmMMM6
P/OReL3Nt7u1GdMZzDrJOgSV8XxG5YjugO6cTQLZeSCYHZEtzmYQjnQD0jvGMmxT
9xgprLks+O06bdP7XyjHNFVwncPRRyj7gXKCOjD2ryDzi+8EWQB1zzqa4cHtJX9J
+YthysxKpkx31fZxtSxQAj97/UxKcjGYvsFLOxAxTXSm4g/5NjwWlOiN0+FF5SDC
JH6HQFdCi/nJYUcgtdJTlz5jxYC9ODpE+bhWtTvHcPOZjn/cJhRn3TeV7zf1eCHK
0Jp+thlUfo7YTTkMsqvypSbQBBj3ft1FEOxT/Esb15+rp7I8kFDgm9h03+Vi6FMq
1PA0Ix2j60T4TW5N2UtoDEXFlcyhHL/r9NEDuTBamNkyIM4K6vok6j5o9aN0pA+w
0eBUvQy5vDiEqO/ZRyaAA1dzY7b5omT8WikC3+/Oe6QK/DBlMP9+DMeUad0qyct0
gO6eqZsx4MG2JskSlxVvrlpjfQnxiD6uoBZZa9qdJBe/bUErEJwDjn18H9RejECx
FB1gN1jUbnEiB7o/E5rbhrEqoDwMv+lnJNFU3V1AurIlYYQeRQeKZqSBo7hVTXgX
a+8XaP/5CIFgRLmjCXF+0paIN/L+zh9i98Dy8wca6nmFZxw54GzMvKSlryvTCVt0
/vCFQcPlObkNsIb0bwkNkkDKbZ4G3l1U++IYGQNcV1Fz5kMPvyVwsKtMQA/N/MnK
8GXjrzpcJ8N58YgV5jwWnPKXjpz1HZQnLYEkMoYfRBLYEtL/GrBZ1zfgcQh08fOy
fUMB0jtaAtEJBqbzNd1Reib31s9Nr5efCK86pn0TReUEvtbVjdvdWey/GaL3omAT
D+9zpVzrNVCQiyCVXPrWxYd226SlMmeYClh/Xr+bJuCQg+gCgz3a+jEUW6HjLRDM
ZiC5DFO9SWY1op0m3Oc6CQFZnefHJvH/SmGpgpNqUTTsDFVD5JnKXO1SB9EABi/s
YAir7lIAWX3QCjswxFaKBA0DHieNkM0cA+bJp1hmzZ+u7IIHeFkxCkvYZy5gsH3U
GTWA9XkgnUy+SgHSuxf9Zv91/rBfOrxpIguTN1Dc/ljsrGziiF7pNpAyw5n6ba90
lFMTQN0srHhdjZxwB6BnizPn95vK+q/e/BgnhCm1qNeViNSWiLte/YB0eaJWNCnM
s/s5hC8XPGfPHtvDS6yAEBbaZl6u2wPN555kqjl7tiTAdgsS4SRBdR7l74iIwCmp
Aie8M6f5gdYUJx5maLnSdwk0RXRpISHoTm3JPg4OraDGwtUINBpmXtBthDHqhDqe
/i3HMB3y10aUg99ioqHUYE47WRgLO1AWtJlQeXLSqlIGvitp+cDpMlj2ioZOr+WS
44TcPdWx550xrj/YT/Ii/zGIjMeTLlj8FnmUE/kEF3RKtq26a/VfxAw1IrP4Ol9c
I9T7P21Ya/9rAU0nL97B//zm251WxPi/NTtA1iJ6rcr6AttsZtdaqF/tekUH/+H2
ocKdDQbvQeBYacNDW1vlk8YQttNfVodYCAdVJe6flnTjcqzvwjtekRXd1By8Nc0L
PyOz1mfXVmxahNpjhHetPSxAu2UOG0/K0QK9t1ErtM6g86cuo6/6S4XXlkatrM8L
9tP5hA9TQGbjx5W1QK+uSIMnJJ7kvH5xOhKrzxD9mH0M4xlYckdD1C9o0JAftUZU
P9QBktCz+73GAYt5TT2NJOVRBD8S/WS17NzR9jtoR1UL5WHOajdxixv36f1yaCW8
LoLzNHhUNTUuIyxUZxaF4oC7j7c6UoNFyxmKFo9bMiKgZGbz1Sy2zP4ipfEBflVW
S93tQaYovfWd/OzloS6/I/tocGrBw1QLFKAINYbonsLmOYrzepxgV1KpKQcTfnmp
X42pIQbV7IN86dOUsqAdMIRB37JOxdaiD6Zk2vK1cwGR9c20dlHtVn3+dqEpMBFq
BI4dn7izrlp23Wn738yCgr17F9FwS0eCbsFfVXboWjbGoQ2ZU/ouKgfSYk9yyMcc
cZE1MGsGnITBbVTx/nkJQsnjIoszMor+dEgzNtUYOhRxEofxlppjT6K/Mv+lbAe6
7zANXE6S57J9STb27gcDHbdvmUkeM2Kjsrmu+OfFgNlwc1q2n3VwMHSMQ4l1o9mT
LZScl0fantwoEfiEK3Vm/UrXx7wFryjweNYl8aQ0BwrJji8NrnD/TZ0elWewc/ih
UnmCTcrQhf36/+RnNY5qjF2X5OzmYCr+UqFb+AD819AjicS9u6Tb8y6NslH0z5EO
QCM64+a6mmFPVRgVZLs/Kf8YoIkKT41WiSMzIKG+0xwrj+wlqaLzgVFW1aCVTEm8
kTtl0U0IFtrKlbSKO2RebnV+41PJlYULoKZELgIEcTxxotG2nIuIep9ws9dXSBSx
JXFPU/KF/ABK9w14EnzhprErFA+DBPlik86wNQ5iW1WVpTpzYhVTZEXnGVHFrTVk
g0aTRmVA+aOuLJgG4ETO98cF2Bc82aGNHWSun1qSCxx4qxn68g9JpBcpGZ8kekXZ
aUc45S9UyF0ckXbws2eq69AsYvVIkQoqiRR/dNRmCDPC6OW4j20ovqYws3VxxeO9
Jw2yGhAIaI5kPpSbSJYnyhn12Z2YFPOY2D9a9GI7LYkfLAVkFcHdR6pOTqsszW1l
YlBS6Ebd73+Z8EXcCQ0JbkzG4msn25O90WiTNPa0OZ5NFaaKQwRoN7fJYeD0HFhw
OI9BDLlMzzx+zA4Ws0SepP55UVVEWsZlkz4iqy5o8CF9gRWHKiYp1dpjbOiuPXYQ
qVPhMh12qXEG2AADuxEmMz2Xy0gXqd71beJSc9qqpKLH5ilWMS+nytTt/JRu0wVJ
SwO/NLcwcgjlswmYstUIz+/P/iozMpL5eatgmY9mORcwrvxuUlQtrWHi0i1LGDSe
P/rzoNxB03kTRO2D9N7wjRJuc88PcAJQLEsbUeUzKGY/UeYZ6K5DiA7PNVeJIM77
oS2XAHkW55/T4BqCkB19GGp12j20lfLgeZVfbiwLfXwGtxDu2uKgFsRRQ+XaqjHI
12L1Y+Sjg1A4dxbQDwh81zi7YbKLuFTEcLYwDThpP2/co+/RQvWcY3CgY1FLqfgB
Lsulcbks6fbmZBwCKIj4fEbRv5WPMWjDWby2W6vu58BHmJwlfajrGHSO6JTNM3sl
ofvN5pDIfa3I5nLhRFwTyxsL0D63xHe4y/IGnCi+77Y3HgV9QiT5fnz+rcRBhxM1
TCcznfOHhPXcQKs4d7D+hv+GEtmEB3T9/88orG8bNSUPcxUQ0seK4Imtzy7hK79Z
Okq8Q4CLLCYqUDkQEQEHkC6Q16wJK7wiKCsAOnClbDUaD5/1HLWTz7USIN5Yft1C
NZ91vnKWD000r2oiWniMVDwqEwszVYkzsjtKBKxkclaptI0CHr4ldcJTb+f6Xtim
wR77aq4IgtqvzHGgx5LEIxEaF8JpUcOpfyz9ZMfHro8fjetscdzF0ixPbjXVUyJr
+0WAGhdMUtI+RepDYBJ94EIuty740ZKYhp2VMei4yZI4v7AqBQpjU8UiM4KcFl9Y
WJQvy/7/QvNnQNc7jIboNMXp6yeomqHBUN2G7APbWtGy/qHNg8AlblgzIw6V8/Gc
Us9Z/wht4uT77/FVWANmeoh8gQeHycWbvCv0zJxWG/audx/+Gdg9fjyzMy1xfMBE
Q4fgi2ul6TInTuglz6YR/IOY0Yi/vVrLiywIrIxrq7EMEsmyO8oDdvkRe1WnU/Lw
KCCe9ZV0KjjT4my0EQdwiYm06bqZEY/XxGXIVqaKF7GTu/HkmqCuYV4VSQ0K3MLx
9+V994/MZtM1IorbkEQfpo6C3r3qXd0cLg5AZcO9q9WK851PUsrCwoK3AlGtXRQT
y8dkpuG0tVUs3NFp9KvZSLY9xK6SxcWTcL6Vcdc5D575FIb9zijpSziwEGK2yKGy
RFuOT9WO+pCV1cEIQnP1y/eE3Y9TDplgMb0hhHpswlwJ0v6OyqJunl8BCBZGzHWb
KRcuqxhHEFCR4aCBMJlwXo8LzOwasIn44Ef3FY/HHOi00hj713acJAjurBQxgAbU
Elxrcvzo4p7Pj/iD3KUAr95wHyyFjRjaoOfcXb1o+T3vhQ9ncnbAURvZaRz8+eHO
1eG+5BYm17oIWr7+CGsOClUGVWauSlZ+gAP7ZSzAYQd3Og9mBWMty6/TMatXPQxX
3be/bEDSvbNXh5lE5RkkDov97yL3EC/WYlbp1FftINql12A2t4vH4UfZ7JzfcO8g
cf/ISzUX4ibHvjnbHWIspAxyVLNgKT1Gi5d+/j5reHpHGc8hJMue7rwhkGrk+R1t
bzLfpt3Qs/KpPtr8ijluyVIiCvo7Fp68hrdpSHTRCOdGLJ7joR6mitI9fr98/dOf
JFsVBMxp0m49dHHMzEpR5zEbF0ibJ/Rz5TPgpotD6a6HSTX5hT75h/HxYo2N8BqS
LusGSJCa/OpT6+ojl7RPwSjx5YNGRwc52dg6k3QtUxl3Pqjx40LqAHL+PlJR5BFS
p0rYNFC/dx56k+6xMd4ZSar3rn3W7q5xEFylWgGz+ij7rcjp1YuxL8T2CrVfM42v
zn5XTMy4x6yzD0ppw3Gy2/XlLm5vp9Qu/uqaa8iVzLLYDZm+sA4W69T+QVQfE4d3
6E7nMsKETbgs4bdzUkU6iIRbSLWoN6IKtnqHw8FYV2qTa4Kx1iHzAnYqHUBHMpln
cqDnZWigJTYcw8Hppq+YElwAHzQcCEpkVmVkosc+QcoGyZ/e9KxOg/Z0y/TUMVfT
bd+ryzThJrfyWGtMiwWwqbmdV5xTdDkuWEK+55uLAs5NaM0dpuB3wrY6YQeF4n+A
F5kV4M0FvcHqED5MuZ5Y7+yBfKPNbqoE1YQDwNwVuQMVrra/0epSUSiFWY8Wj6oI
Cv/8Ik7qpUXavlhAbj3CbNtKyrG9IlTcF3Z8ocr4zXQlWcg04KxeL7QlK1+2/ppV
SC7rthFQF1sh2CR0KbQJ2IF5rOolt9IgJyJARAtwyKZ7o2xqTEqWg44Q7GVUPh0g
EzzXYIdQXlv4X44hGhQ3Q5chZXyTZ9QXafNUFHzo+PQQgdj6LXzcSRIySJ+6fE0i
BEOe6Lhoca8ca9LXRZBvLD6Uj/b6agsnz2Yt7eVYEeP+KgDR+76GBGuFCxaUEEAM
ruOO2y/WAQcAzRMS1BOvKxJDlvkMTdJhF5xpe06xNq7Nz96LAHsgOg0mp/ATw9I6
ogbJiRjF9sHO0OUz/YsZzFdff6mWe8X92YXskm9M7OeIkl2I3NQVGdP/mGyOTo9S
qlMDhNzFtTkmBzPCZI4cF786yEGcHuean4LCFTnwTJSf1AageDfJhJyLf2Lr9Ksq
N3y4fdf/TWPT9UtxHJjzzj5vVhLwT7rSdJX7b7clYWCMguLZgebPSw/2nUrh+vgB
gKVMLcQWaxQt4xLavkzzSJSKOiDuwJ6BuFqetLAViwRrxMx0Lv5bXGIGIGDJ0hYM
mR0LId+QCQdQGw7Xy0iCmhMiTlFwcC/xERwMhefKxxSs5tz6MtsLcaraU9HBwNFl
8jIHxgwVl/XPh2ePS4gJcaYXsPnr77vYF8YtZQWkx1BzNJKru/wf27s6zHM+PHtJ
8HFVuY14SQIJKN7sfRUFEy2Szq2v8zcOfiPB2aI6mBLWEoKRjrAhe7LLr1dqR41p
SV79+yfzbTOF8bgGwGtPpr7K++9/zL5lF5ZVtllMlwM4/lg5i7ULxUCYEzapIn7w
pbnEDfw+8x5fCTOZSwgR7zyikKVhdyQX0j907oQ7lhsyH9oTpprmgPNTfaiWSYFK
Y4bJajsqQkXx5qAohNlseTYOMaH6IJKu4Y5hrnyapuv/fhCi5hdDXAIHHQzflnp0
xw+3ad3ipH5xUvS91V6YibVt64NIIUkxDRnh9gF5HWHe91ozpH2kPQEM7vezYKlU
p+zBHCJGIpKL5l4gzO2o53bVrmnjZCNhl97kNAPiyuuiSfCDPQoEPDsxCLjFtCr0
M7rumVUAE1t6VlN2gg6ckPgDqlrcrYni5kJcudnpVPLmitqNtdUWQyerrXM2CThS
M4BQdi3/QFcPNVPxad0tQb+Z1f7iMBjNOvRhJqiDbkxXcZek1rbffydX5PTci51l
dgLdBPDcqLgzH0ZS0tvWusPUZABlkrNbHG5Y8ndJUwGmpMXEIKOevjTODSTUq9BZ
widVzjNXQXlERFt7HesydX//bWUM3s/T6ExHoFUgeHdXE15hB6NxHFs8sIt/M6c0
prba2/mP49L8kJxL5BwJFy6/h8qasC+woxhpW3X2A0XBnBjaRGu6arasS5P7ciog
H0J+U/a7udoaYHyqrvBnN61uOnp0aZRcGc41TAbjzwkF8c2DCdJpH2r0iBgPeyva
m8Q0OdEBSST8WeGA+uo0HYk1MUKuzpqMyRZh9D2KHrXXBbJVmcjeVYAk+ngSfGGw
y+k43btcM8b8u3OF8lygYFkcey9pi7vg2jWPCpJ3p2p9C/lh5nPNlfmeRfhTRKl6
+tSC41CsgHWlX97VMIsVmpIsw+IqZu0Da6WhxVEEbv04Aii4KV6H/Pby6ydO5IPZ
lZXrffsjiHsmGkZCwBE9U8Wg7e+y33KAOl98oAHyIb9tLvvvpkHuYYVobtjnaEvz
1hj0StN89qFqj5D0+QIcoL4iswbsnxfvOqVM9oBm36R3/XYipm5e7wwrCu9vKM1I
KXMMLLGH6U/zw80MjLFAIwzHCOYL9pHJ7ge3wKkwuKfoIgLLlKXUILnxatHeDEPw
J5Cqpg/Igsy9r98wp2sYCB3wlxLaspvwTpe28FyEZjMo7Qzy9yBIhmqpfKvSDFuu
t9c737fw9yPSYpkHgQ4csksf7z0JkYs6W/09PY7uP/yfrlAJWCR1UAFx0/qBvuad
CNsKHn4hQ5ILwyfPWZPrE/08U/ZuzDex3tklpzDy3a3yz6X7uegRTrwg9z7eA5IS
tZIp1tgQIFvuJo+rG/cgHcFPpBZ631yovQFltoIdZdNbyIB5Ap+flHF2AAwQdaAD
CIywmGzm6WqBeMlsCMpXCu9JZ/cMlPYmG/+o1JnDHFGeEDr3aPNjz98hkillg5Ac
TvZF9RPKXG2DFV/xQCBfRme2Q9NHwtrgGlD7rEgbblVb+9Lax96xMb0Dmq51wRJL
EnYUkmXDyyuNP3v9SVRuTSW/54aqpqYn1eDfFccarKY9ISlee4KTkcwJ0LyCZihW
2KvG7b14mLA7rC8xgrMB8ZkphLtv0qAMXfdumJnvqWUMm/YAO0t6G9zyaFK2+VvI
DHk+0NAsUDpfh4AzXh0YOnyyj/OdU6xaffR0+Ql7QyGDVvCMJ7VEYqcqVQuXdSju
ILoSFfL1TsZ7CnKZ7l9XQmY4Se/x2yDNOmnRL1R8aELf8WyCzedjyHKnDSEU3E7N
gffaX1yvdcsxBrSe0ZDVe8/F43q2kgQHGAov4VAPnUzP/DRp+SNDqZQaP0qeeewl
trtAZ+tK/lfSPx4w9Bd4bKH+bFC/DR7z4jjWdb6aKph9ODMX5EM2AK1EDMBsBbYA
h8KYge3Qj/GoqnccLCPlmXiC11AW3CryqdUEHOp+3AUKJdApsKB796BIqXXT+vOU
YOwTZv9OlbP+Nm8wcwG9xG3GD2JWVLXddciz1bVcACQBc5aGF9W7UHkq2JlnkjqN
c8RDkTyL8ZFq1fJaNL7huqpPitlL6/SX1oH1tg7jmGujygCPLmV0JrMM/nvf+Vo4
SYy/l/QGHWHUv1cBaN1N2EAIEBkpP8S/KlYXjGByBAeeIW5GZPfWE5jNlzrcVCRX
lYhFk7fz3h40s0tU7pryPSC1KUINUJwnmSzP6A62+wbnSOwKABKyVnSsB842FqOq
+F/7Q48DTFVKoyX8TYftn6yd3+5lwFJ4ii59rvBogEjFqh22G6t5zXbhksQ/d6s1
Vt+pQLW9gz9238DU9HN8dYZdyrCKtrqjx721k3qmqG26SMAOTzWz0oeM9BlKmVPU
OOqSeS1B5ni8M8acnQknjbtQKFPC6FzSDHAMXmH2rkv1fhlIilb730GsYhk2OpIA
iOad+K6Z9e7/OnzTsid58LugzYKeOG2LxKAecITWkw4gYJzUmZjr40lQgJLlsi/K
b5fPOXe5Bx3LKnl4c80s247J25JV5EK5dSqWMGznBzMz2dpzRWHxpvHtCWKx1i7/
Xqp44hxx842cFR/1spkovAzFU4/nBgxB9MFPMAp5UBl6DPpBDp0wDUpbOuaM13rs
APZ6vSMfQ0O/ocHxbpUbgER0c3JQs2uJEW+wMGc21racqhPcOuP+fB+C+3nSLFNZ
m8rnDlRX5YvyQ67DuHBtemn/71Dg8SGgb7osbtsAGWr6LmDTyJ8N3d9gJ1FrAVbA
OIrfGgqQJI/kKNAZ1UmhNIqp0woLfDzc7wZ55+Fyi2zDyfk8E+mW2b2NbfHhknPa
Lwye8VRjtJCNOP5G6a5sUcfHIFa2bhMDl19Po2L3s92rXtNihOivim+oeS0Gl1pz
AMzJanNrIF9kZeE0nVwZyO8mjKfjkt9kaoj8PND8+1ia8qYnrb7MkyyEoy4jMtuL
jAbwp+pXXIhs3lldz2PET725CZHTMqxxU6yclCamwbtFrZsZX0wwFSsLBQRFsE4C
mRdczTKrNw0/LtmHkCZUBtm5mqZFvexBCAxImrZiShB+ndE330Q5t+LsBla+ERX9
Ml+uaUUChnDXQ/TJKim46yF/bYoW8+IPz8sCIFECuOOH36QrT7kM0wAY4sgK1ysL
dEKe8eAwGHbBCvDwvN//XCGrPSTg53+9vvsaWmS7eT5ylQyRwLh2it6U8SIMnQv2
0wMCGZT6VPN6Jswb5iqhufbgwTAbZVz7BiSViPUVxlL16EZh6NjMgNCSio5uUUYk
i1g7TYwHJQDwHuwpMY6YyLyTDcCtw+evQEa7uUY00zYJ5RgQXZNl7Naazops3zbJ
7SMJsh2LVQH3qXbren3YHUoclm3MuCYd6FY4S89FvRzejK29L8aIEQnyV6jkHasv
xVPxoCHfcIG2fwsehHaI67AXa0rW9LNYZKJB80wwkxZsbPXBlRvJF5nxE9eygd1z
JxyC8gZALnnEDO+67RNC2POv/WZ3iRIpCgxkqsIpxcz7IMYD10cjJDdW+rIUYpOy
jgFeB64HWbFsypCFZbSTkYwKwhMBCFJTyehqtzGNZglLe/x17FZzIRvGGaI5OiH2
naDQ/mI0gEsJx7HlzuP2MJ0+Wq6Jkwe3+l1zoAW26/iov1QmH2i/pGepdF8ZfxzB
uU6pRvjah0wfRb87pFkj5ZiV8Aoop9DrwXJe+HRH5IFK9zJ9yVHMNgONe6/0UsLg
FCH7APJPG1kIuUwWOKSNFQ+0R3buSIKRRcWATruHar6ab2XeUgntpOlXuEZ25PbK
YRUKVq+6KIJ8tQVKVPC1qxYnLHRXe1Kqtbf4gX1sy5PMtpqrn0O507jJFZZgOKpP
XP60siPus+TZoQWlzXs562H791DEc0T+igAS7TLg1gYgStoYNPNFiS3aIOvrvPxN
LLEnwryLtgnD69DPPE/k8c9dA9yPdM1r6DIckk+2TlHHCeTWS6aPU3nBi7fBCpPf
vejDVs8rcm+jOfsBVj5k5Nx0q7NOvAtaiQpYKiiCXQ3zrmUCx+zGXAscnyKXipC7
/wbfVy+m7fMuGCb4OkOBLkYYC48nef36zb3wUkQiKCmgTijE9meDti9gSjgqzAVk
fnUGZMcfzbER+R5bXhbJvVwxopw5yPmOr+I8ij+HZW4rKFzgnKDr09OHJaXARnO3
gejQlznV4uCXXIEIk4uuedpcamfZLku98YtmP7it+knTQ9z+a76MsJJFBKcNXwIT
gML6JWDSBgLnm+HXwIUdA1ysbTRLAXcRCMoS9/yJKLYxd45FKU9DUrIJXzzEjQrn
YfM1PEq4WGCV6RQHWMY5qDHs8C7BQhynZxrAjrluyLds8FyUC4WOo7lUu8z3GgZ5
08me2pemjx9WIvKu/IAaqNJDDmR+cirBqOIfwfYbe+dR77awz3xAZ2f54LIucYQk
X9+P42uaVPtQZhYR5Fk6urPpl+0kLUir7yW6oZv4cSVnA0Y/SbT69ElOUj6x+j3c
GNjEHUsQSb9kLYgxtEFfcYU11fyaxn+7osmD5ChvfdX6CKZulT6nkOEIC12Oij/n
gVwjlBpGECHYp/GCFMwfEBf4Nv+E2vg5NYjyGeEewyTIIyIo6G5WXbJ1AdJitrXU
gS6Tjd9sATzk9bSkm6zPN7WuAy+caKRsJcdk0tvdSccwIaOPmeRBxS/yvwpl7tVc
+iVKX102CoSkEpnHHe78jjStHofx9y0jcXZ/00x3R43WVlqE2tuhquEL5+SS1/Sp
C56Gug/gnGdDUlihQ7gf60kE0FBljqDdTJZhycVoKbHX79k18kbww1eKBuEpwgFw
NF7fuSKLpmJ2LAE9bkHFkTu2+8/5ysgI31PI4R867sbVx+4mT1/gQZICFSS43lnZ
qUAcHha+hIM5NrmWRh04smSgkopFeoiBaXcq2RDaGyVRaJpRA2e0+JGp/bvIpAx1
cU97d1+qtR9AP9FW4WF2Z5HfSW6shOcHkyH/4l7/v7AVm5O4oLOqkubyeM3B4Ijc
4+rHCB9VhKhKZN0WZzE+DuaME/tSaxoVGehaB31zpT7gLbgEAcpFlR7xWpwuYFxv
L7W8uKNFsTVaVTRWDFIQywjskEyBSsXNoLOZeRM+fONn/tP1CMqp7LA6m/k3PuRz
Ap+eZ2fLAD9Ui59kvBvaKI4RUdPpU8P0TTrFcNPgcbGfC8SrwEi+VtJweFq+1x+F
1glkVTGpKqE3uE7ltfNLDsWE1NwTqqiFRo+AdDrJmWtj0ghQPTJEM0KchhzgEgE4
5ru+he0v+mEByYdXZ6L0PU4vX7Huq8/Wj19e/kWYkCX4pM1wDR6Afo5LVFV+SljQ
FlN83G9eZ4lGN4Lw4qBSugfhfMLhXC0KL/DkL8+R0AS/Y/G+F1ooXmwFcQjL6xk4
UZaEotGN/NneTWkdvCJdvRyItkMmqEJLHzWDWrtZtmb3haFi1fAYzCDBfFiilPyi
1RR8lelRq4TgDPNbMJJ2m/80FfgpTvi/7CNpAYbQ+eAGRTpqB8CNLvnnhftJue5Q
eK5zj1wp0V7HmRS9CZI01xz6GAvXgpq8lhY2brjTuV7RgKR5UOTqh8jvsTwaUIkn
QQnvbTFsRQ19yQPSyyHGCT6X2j3HRPRxWwI0mz5aE4FJeKZ6FRgquEy+olRTgPew
4mSBerhNKIFlAPzV0jjkwN+tRYtp35WbaveZwg/qjoZjByc7Gni2ks1wPgr4p1vp
bE4Shvwham3GviYIZlu/i6xWfz4D2x95koAlFXW+ftADtuT4t2aLJOpsSUnkwxpf
i4GyRqW1pXRJAPYrlhGtWwwnibFonzzFg/tnd0tbs8/Q9RLjljWt7qcVhAUdMwwu
ijMefmtVoMfO48YgbPm+7gU93aWvLo7GIySZ+KPMkb75j9cVE55bNtKc2hx0ay4+
6inmNGDyIj0oFOlYmQtaxlDy+oM1ZmYPwuNN5o2AA5FXuTkv8bWVnUxF988lxbCe
WjjMIg0Jz6TQrwvJLimne6MmcROVu6X0nYarWnN92YJ8zAjdONJW0AxTEJUre49C
QRnWINZasAdSROjBQ+R6ehad8uQUZj+odxKF0EC5nLjcxIAbcvdlTxy55hBYbYZc
nQ4rKJhKn6fAZcw8Jg2rXUFlaodhr4r2re964w+clQVFDSSdB4DgO/qwRTJ3EDDk
YNDdmMMkZb+5BK58DvWX4hO0XlM/BU50/R3SyVmV/fWSIXN7OdlHWlxwZOpoofqR
4mrLsNaOJbL5e2Za+N9FvK0Vcs77jOwASR5XapUg8ZO6gotsPoKUx38k8Cq168+W
4Z/xN431w6Mf1iw5XG7l5PILAFmVYyt0OTi2rrJ4ymNhS4NnuJiFZDw97I9Jngeq
iFMDTbNovwBKfXw9op2+OaGzkG7pMDul8ZqMP1czSCVALJUtVAYnq6thzMvRzqVG
3F/HAAY6+jztJUqxvUYS5023P0ILmc9odzWOW/4P118akYYM18gTK1hmCr4X2Xsq
VrLEgrIuQ7MAe1lvOABJGF6j1mUpSb1b5yPeYU0HrJnNEsaKz0nuxn8fDAFzv0qA
ww4WjQTnUy5cKnAKDmIyxAvSlbY3VO3F7d1aNF9r5q758J9EpCyjF75bbdsVrC68
gVMHJr6Q5dhV+nC0gK09Cnz1RQWu+Ud/vhQ5EgrDhtQTsxkoX1+5zfU20H4D8k1v
xWc82HT5nUIZ0khyFNgsfDr/SLGAfK/853RGy+CastbMFVvVVkb31cxXpTTP0IoF
0gVx62fn5d9KcpDzwkedVIQ0g2WQFJobq1RVo5llkbsbA6XTHKymlgzBOAIn/zpV
296MSaaBA/K2hpqEE98d+pou3ZpB0vNhQ0npt6BdkvZS6xNuA1r10qa1ecY3Iepk
xd/a6o3KwZy507POUxB4MKPZDaBr7OVNyox+oPjKnsUNjI3jdZActhlOjh3LZtrA
lbqhHxveSg04r2VyMCWjNGSH8izVqx1e2qc0bPUfcZAXmXv3JoM4ZoyFB1O0fQjZ
L2Oz/qTBmesBLxVxZNYkl2xz/k9jCYZbsID6IK+u8yXZF3dZzaoOfO8OOAe6CEI1
XEjaz5p/7l7B8NPDEG/CTGYNj/n6XlRaK654RVrj18144H1MWveI7fQH6IPh3e1k
M+BxyWopnE/k70O4+gtH4wFZkY6jAnhbKjRXy2Vx81/NZy8pSSJNMgwEixkrJDrJ
0VvKx5geKopVNKf1x1RhgjPZ1NpTqVlARn+q9iudvhKJtVWI+b1B8kswP4BsMEWh
oOaPZJBihT07C83+iZDZUcdoyxUS/IfcZK2qSNlPUeky05j/GZHwqAJtBf//TE8z
7JS4FvdGuQ8q0Ao/DkG9ESiabskUMNXhXGBeklMiYkyOGRwljth61mXAGMm/SggD
hZXDQpqWgkinBzPm/1/SeXo93xl3jMQgqh3vjVVerJY5KHrgDPHs65s+xOFQsww9
8qFqaYfnNU2pcLki9xk04KTVqv7DUSDjN/lOx2srp26zm8TYMDkSzIavrKXz/db+
0mmVynbykbUcwmYTlSwkPr8fSeEoxrVNKwUopf4aczRftW0E3Dfo4aLOaWR/rQf7
ero7AORw6MuyMqQXtZ7Us2vtS0tUN8pmChNG0AWfzwtlpkiWs7aB1eCNotxEzoMK
WknwOGpIORCHHd5zYu9lBrVp1S7oGRoctjqvAmUsxQ1Kb0h29dBoEM5Pi6ehW0jS
agY26RwXfEXrDbSQ68DPmyIBmk6J0kG2GXvKzAWGs7R1TNQGrFdjmafIiLXwOP/v
vatMhRX9dYKFUbeOQAYwkH7G3SIt7oXHqHzhEYfmezfZ/b62Pv6jMiCIkGrZQpiE
wyOLV7HprwAelBdylR5+rzPdI0TatYdQ2QrnghPM0b18oBcS5P4Cd8uXq5dmjGBj
QD8h5BXGNHFEfSZ+DATzFdrxy9mNRsTSQvssHb6JNZLwcX9UaY06PT3JgEXx8pIw
d0YUcq0aKTLfr81o4sHKPVHMXyzj1FkHG3ruosvtHIZ8bD8gRy7c//Mx2mmIOfxb
gsMnB6DtOOVdVFWaWCC5bmawFD5WeyORa1QhCqDyEK7YwcC43TLLGLsZrIU7kPMA
SyzRNHAgV8QuI9oqGZS+e80blFwH7k/yyoFLeY6VGZtqpF27KPEvywpPtM0Smyuf
FReAFVXnmmna6a3iiEGevf4Yb7ntqauDdKt0LcMC9cFK8i2CGY3DVcea/A5Qw1hk
wzj7sSxnPIHY0O34/qah6/Vy4cnTKCP8rkBmFkAJmwjaKwzpkj9TiUH1tSGKVOI7
9OYaqgZnSV7dUNNU4ElopES+U0KBr9JkWJR7/gZTZWyrq65fWRdHBBKb6kde2NMB
RYZR5slAsXS3QIvWELFGVSeCn5XeUfsf1GZPM2gnVaoulstl40rAQMoWsX28q+dH
SOxk9FKwbtFpTliDjVCfL72ERsH5yOfDpXaLeeoJ3suvTvV0Npv+qxbgegsZvFpB
kLBK9RIYlx1s/H/AFfaYVQxOrQGT75g825eq2px87GKLl4TAlMoBUDlqq2QCJ95Z
cOkHpRHj1O49wErBZsgp/gK5+srWcWMeYyR6gXA7coCUXi7sgqE/w/+RXgXrSIe5
yt45IwBFKeRCPP0zNF95EjEX6GnxtcFOdYIu/juEw6jcBwBDryRdjxiIzVesQisX
1HuNsQsSMXUE+e+NrcvC6b/kYvGHR5+BupqUAIn9k7aashGNZtsqOZsr+rbccS3j
whm3jarDNa8EFtYwHYWj9NZCNGJJ5BSsFNqRs4UZwdkplvauDrY17rFONkFhW0nr
6o/F0Bz21qzQLQkIQxVBj8fhQ6zRVEOwa09cDft6nA+tFIoZvLff0SGrvzfkHZPN
p/q1YaOcg/bK3DmgQSAaez/9SGvGXJLuCp5kDHoXVAlreI/HAtWmPc0NX49D8Dxs
2zB9tRToJ3zihmAFG+U6geyUJ9dFY8rRdyfx1wVobhLfcQmCZNE2Smb2q6eivPJz
2vuQ03jnplL8T9Pg5jZ+gWNUIedBgt5x8cn+rrVjb/VNhdXHvVcuurW0Om7XfsbB
UfxFLTCDwuGL5OAKuo8z0PhA/zyNDZL44OO27IUlmXf7Q2jfSQqeoGu9/MkPmaZK
T1bu4y7Xbz3EYOYoMZyLQNxHqiDIa/r3YczikqPCMWHwpaXdopyBU/uVwFofuO6+
6bLlZEIm7s86GtEMLUQK0zUx4zEOaox5WZkJjng7noM0redHepZQNG09nlEKv1OI
qDk1xz7QpfW4JHq6oCvj41WAFpgpw7uCQkyczzy3rsatzSDWCv7sivIUsMmrwUxU
lHoRX0mZmq7mQPGz/z4ELmfnmWDuuDzdL2N6AI6BOnh5zRZAxCncJ8br5R+OI+5x
JDwpskDXnq3+CnFUgAOBA4m8A0SmqwOrpLoCMfOyUJ0FNApgAEpsOZbNA9AP722y
CNI8rILO8TaisZxJaCCQq7P3lVwYvRWMdG1D7BCu/eeBW49jkQyuLreArHTqwe0d
2S/bZ1giNbE+DAWPfQyvFquvFS1+Zir6TZPFATvFJqwOUg98Q/QaWrEXaIOcTk2y
tgwJtQAgdxti5J8uKAEXTZOOZrkLqj1cGBc8QydF0odrDOPO6PyCkNU9ysmLyybS
HR9TzSk9MWyWugjew9gHYhmldeBvCY2g/GqjKLe/DM0HreuZ4DPclW314CwlgKfi
iZKpJPuOOg37xyt/4IedRfnp+9RtdKQbAxoIoeVy/XkN+kcMB9ya6W53miIh/uLv
8BMEyJMcHPdX6eHd49LkAznbODxiEYHZn75S9m/sdUsSplFjLVjSGgUZRbnwQquT
G5/o7W1Pwooq82wNEKLdZqzj8abOAgjgxMu/VZKKYhvW9mXVG079QE1LGMNJjuDV
AAg76cAWaHzKcX0p5FvCcsYaN5fPiMIzKuaS9sUSG370ADQ8l5OuPTlK/oDp4sBw
kmGhia449YrrgzkwC16HuYjc1zkizAKmCwWnQABLFt5HIomHxPew2UyafzDmo/FV
RrJpwmmapnZp5YMBF0cEhurvWnA6afuGV+RrTIy/TFs5xxO9d8ZN+Ywy9njpa/LY
kzMuo7E5X9fq7hLolpHS74xY6EIc+eBfLYLrlQ0THSCtTll4AociDjXj1E06NZqV
IRTjF/9r+X3nEM0KPk4ZS5sjeFrCCmt5nLxA5kbuz5G0gTJk1jrz9AJTBcLOZHMc
niBXQmig5OFasUukH0kWKjLzTbnftQeml7lsHuUdHfxRJcPwcGNvXiLq8bs/H8g9
7ape/Pmi6izbt2KXTcSAyCzzkzUKRaQodA7g9mVAsCMDzotILeqa+K02QILT9PJV
rN/j8Fq4XfMRiG9DLjp/y48EWZNRSe2cqbOhpVrKMN9z5VoBUB4QYCEopVh8PNK3
vw1n+582XkIbof3T0RxdqF5AlG/Alj8+F2nzrT9bDThl+ldRU9eq95ynteKTtiUb
n8h67POJT+MBLVwKeYzWZi1aVrOQC9+AbEgdB3ddAD+QUnVSPdm0zm5c54yjrfb6
7RzBjCW52zO+gNC5hyxQJWBTJjcDkjgWXS74FfHB2e2Ak0ygCrw52lXmibfauoen
daYZd/FjkscKqWvR+BPK6BUhNdbuUICl7gJd4hEucAgIFTH7I+TgrfRD+OuZ9uYm
eV13+XTRo93NnBNv9dkmp4OsD36Tr+2IEwhK7XMS08HhvUBZF0GBWZznbk9W6h5S
iUzY0mfxoqR/dT9zk2obiCQo5sR4p3gYDP724AGFnVsulSIwJBb/E0zjtWtru0jF
SabwKpn4yAbmlNmPXn8g3nClrhkcu4io3NUb0o18ZQsu7RkfRGaOFBZDN+dN0eth
IPNuv9qaqyHHUs1qqtpxLs7PCu2frz7meX8vUsXNPQHYfl5PdSfF/7C13ioVhKhI
1tsINLACykuLihIj6FPnVE309vCqAAvKgfDJnVQKDOqO0rMYJQOY0YnE30zs0AY9
/Euk5V+fwBjUjiAS9J4nqUJ50qxL17YCmEnbTaYjMC9GcxTEjKqX9X0Z5aKdj9+h
artmH209YzJ/qvCy64eOayvWDE/2mTX9um8zBMNkeNDb+b/l2FekZwBf5fbZtC+n
p5V2M2IXldVhd42iI66r6N54oVwqrndMVEEKw4dMXwhtLnVwWVm6ECuKgRyRUJ82
FrWuZtuYF5AhwcL1O7AMmIstGeOBANas/uhuSoTWhTmbKHfx96n5k1avkc7ffgbS
MVpBRv/usSkasikmeJ5T6m1JVD1PgaCvgNp5XbwFGSnmfQDLWUqT7zdthPnFtwne
5alg41HbYeI0CZO1LwDJQFU++cpFvrbu3Y8qykST2Gw/nScx+Ktta3M9PCrcci5x
BNwhZJeYnU5jBgA36ghi4fgfnRVVo114MZsb1Ctdl6I7UYPP63yuI5sz31hql7Yv
SC92mSyX/L9F/IJ0tQRPohqmDrSOOA487v0L/SPoKWa5w8wpNo5vbOEn+ysu72A1
LNJG78Cv80cS5vVlfdUJR33AYSx9ynoOhi+9e5MQHlx5slvCBERcvlvIl8AMWTQy
KYAc98RoWmxia1MdNxLLBRTX9P9hujWxLUy7mEgtaG2S6jURVLJk79F+i8d1KGgq
uVCPR/rCozD7x7Gomx01RK2p3A7ZpKR3rYRKLJN3RDSEcjo8eKjehbmSrtpMgGjS
VXbKfx9jb49RXB96fW3zO4IXYazoTCVv8GJWzxF0fEX1HRzDzsqVItyHRpsFEBwD
QxRgogHRh5SGNqE8xr44MDH0/iBs7tRL0GcKEqFI+JfJgflj62hP3Cmwrg1Qgjbp
0hJgfEsp1qaqys6ibTnrlLntB9qBu+QzKN1X+fTENSqUO8F846ZA+8Aq8V9fiES+
fKguCXLaNIV9hwqW7ns2cLvQaXR6Nn99DT2fV/ZGGFJIo54yVYvTREGXaEfEFnS/
ZOVTXG9hYh7p7rU6GhCsJoAY5P7fUYwHgQTqJt3SmLeh3LbEp8pNFmEsRU8jgJwH
S/eTE3+DaGsMsfRyfp8o8R2S/xRsxuTlOoDUflPT6qx9RAtqzpctXNmTaRl5bvcw
tidNvWXEmAkqOC5LKidSj5F5dXY0TA03I1rlsOC47gaO6+jJixWkMWsbblKuFtPB
5mbqRdoHvp+ULIoAbmaz5zW+HN+r013xnyM8JZ76NcWh95kJLLdkmhCU67nxbXrZ
CcGm6hkwaMF2cVzl9U026ZGLRX3dLK/yH3WoaRILAnxlb6ROCCarTiztEbkxYIFR
wj/nGaV1ckxHGB3G+vnUlp0etVjKhmhy+OL4xjJsldpOvaSmjdFYzAHc9CZATXVW
Pps4OKe79kjoFq7KqCibD3QOcEaTvz7PD3CadHctjSoeX7VtncpU2JlIezdMPE6z
Cxk21lMV5Wza3l8p3e9fGWeSBlZAnIoP+rCxWSEkoZIqt2SQI4+btmXWTfhGS17Q
LuXxSLXgktyl8sNtEeW6n0P+7cH3Jx2VuFRtkYyjyMZlsyhX7pNBSe/ULeejr4b+
EeTscq5TrlZWmn79Af5Wv+ZlZWUff3prMEibB2V/VmNliEmhxDORt08tDYgHwxG4
rIa8qaUuu2wUywhZZvlxZmKHQfdII+mx3ZyiDZWaVylQnQS8hjqcFhx4ASBkqZ2D
AUbdOIaUE9p5MxPFJ40uvQqCqiuGSFc8xxt9MT0ROw8yXacSHZtai3wFXi0OC504
/tf7CblELCw9hzluRbCJ3alUqYAN1igs9LH6z+EW3OeWDBuWmist0p4yxXeyRzSq
ot8pnS024jtlQakOBJ/75T86baGoFA8PdRn33tZH+p3aGbg4TBD0iZzj0m5/UHhy
OCOoTgK6MAns9c4Y7A9oShjCS5QVrRrJL6FM9lTRusO2g706ylh83FnDxey9rBkQ
Wq5YOWAs4oO0SR+cKmbWuIkD8RqsGaywuclvD8wheLm3Alw0WHjtJyLq/TIipvHI
ZPZ8jOvg85yqdwX6g50PMAeOBL5EJvesVKZ3RmJvey5ieNJ/4CKiz4B5iDnof2Bw
tpb7CytuJwdbATXfxKVE6JtjvgQhfNaP7W8ec0z0rEIx1BLsPQYV7L206Davalzf
ZqsuEtnL0SxIT9b59vihFwaW6Dp7IvuPZHqNUMFe6WBqxmCb/RQ3dwZCHEgbuzwI
eh4113JuV5Glgzq5LNLJhs0csxltVTJzsBVoebJx7Kca/juJGs5dHfqldrKQW6Tk
by6ZY5Xu46eOWa22022zKYV5nh62/rv3WpMcIVgXmD2jTU9UFrs8yrjNhPM1rhzU
8jD3qPut1wNsmQ36QcTm0THGpDouMpFDBpPMD1NLZTqJkP4Cy3Y2bqPJEMKPK5D0
qAkVIekfRwxplxN1iYnyKwbXYtxrlCVEhzZ35Brclmbd3UOtd7yHM3H2EKk0bEpG
yaeqbu8IocLZjUfFLo2Zv/oFRNOU7pZs4MZu5NFlnhLvnw4uvFUs2no4MUDO0vwW
i/2I5dCbkvsswbqf5F0AjIw8q2k5HBoPtPdNvTNYew+rHodJs85xSECjQ8A+gq8n
M6zEMQEgD1jsFOZCBIVIO6/lVLpMdKZzk8WJy6J99YP3sC5hGSxC3Oj/NBkxlucI
aCDd2pE4JDtuXAnTpRVGtMqYJd4yrdFk9mKYLt4ACGIn2zgw8pLpE3H57Elk//nb
uvLkiit+y6cK+Q80JjXSkjuMgQ+fXB02pZvuc+pJ98V3X8J3DccjlTCf4wrm7rTt
GkdYIjJ45mIPLfXQ9vNqZxEjdl2xBWYY57URmnj+ORrl1QLFgpLx5DuZvzk8OOnf
qoSCz4UKeZqnV6bJETGZavy8nUsWFx80px4pu/FuGQaTAxpUJ3Qr1crZhShTd6Ul
S4HHQr99jpNz5j2gllUFL+KKqw6TZR8hvLNdit7U3uYXwqXGC692M7D8LEgfe0us
JSyVFCztEvvFDrd5eogOgXYoVkPV13ntPuS9icjsgcwEIo+m8fqcTDfIfzOZnV9p
VJt+46TgGaEB+W+SlVBF7i9UXeZ0hVDzFoBL5TF5j2MvqsrUTK9jIU87xTxywHI9
uOO7WyyTiuIjfEgIfqieaKB4igKJvWZrZy/c4c+sEiP6uQxDXmXFvdqSesFHr+XA
m7JjNehEot+vHz/N4PZZwnEPPuJaMHIYayuYOiWxT2dD3FT4F2WP9ylIgELMb0x8
FMfKl5meofFJ8mYDdqDIeklXvlWwB+Kyi85XiHOpT8cFvo9GUSPWbVVmQWtnlmDG
P0MxBQmUbiyZH7a9/a9V3lpGjkj59x595/N3P6lKSaE2F7u+Lkl7/CEyr8CjmDWE
uqTYBO2YnJRbzm1VkocSigzEYxAAuZs4WyApdDFMamxkVG0WPlYusuXWagUdXu3K
W85CaflQCv0h9FfuZLUy7LTNBnavhcEQgIqZT9HUpFUrFPdycOv6r42WWIQIRByr
gHc6iTsFxwqvsv7UHrc99KvbmooXhdkpfMMUh7BgHBVzlOjtROEKJILW6ToDfCqZ
cFuQ48PVJr6IziMs5/+5/jmOlRrXuB2f7IG9Ze2NcJ1dsedBPhOCEyUtDgTTfFUS
YuX/mDmthJTEz/7qaAQG6O2GTP7UIuTEYQJolvkp1vjnOo9tUCir0DKnuduCEDBJ
zue6uCv6lbvLdXT4LQ2ngOf4FferXenLQEnAFSQ+auT1rF2fP+TKHXnRkglzFVf/
pFH3Xm1CaI9Gv1eXS01bVhFocHPXwDNSW9IZV0SuGNZJ7XLU8PA+1a82tU+PAFcY
SpyryUxftN+UU8ctu8zFOnapm+h3mbOtLi+QGoBgxDtyRR63DCDcy1/KhMqQVNFL
iAwBIyrIbAJa7OBWhEHv68wqTYsjf7igBGc0b/MaswzCquIs8BqVY1ohCThKKTIb
BHa0IabE2rRa+dh8o/o+OBxkr9uOwEOjG0Otn7E3U8LiSrc1r99HPwTOIzLcNqDA
1NJghJSmUzqbWgtmNOVXJbQSPfB/287iuvZ4e/knrcksZ2BpaK3U1U30lgRmMFJ4
oSYWEBCeg9gAfC0sUrapXqO2gddyCNJgG3D69VojVUk6mAUHWiZFQET9QQwv+ZSY
3qqUIBOKFLUAQnxYwP9SgSQGqKrR6hqfFunhTc3ESZf/opVDVvrjKEua+nmWxui9
ywcwutvL09IR3eLDi2PrcV8lsp4LVp4GUU1Agl08MPLOE8ExckBmCEjDun6jlwAs
68ZfQOVi/nCgNEhbfegwte+LKWp+VMY3Ondkt6mBKq/cV7iH2sCzjOD7AcxW2Hl3
CYtR2X0bJakMU4zK+l0DIJZgpORY53O1NJ3PiyGa3rJeKz5El7Hrz2Ld1Za+HSZi
e/RdaI6bMwRRiEdIISsD6j38HOUNyj5v3GVGZCU3ddJWE7pCM58PdmGUbqZC+bRE
Pg3F8LBGvDUGQdcNY3JEgOzwQ+zhoB2u6tZ15L11Zl7sczLG9iuLH8utZb1uLo3d
0gKKcnSuclmOAlJGMdssgyOgUNtUPGLlmNH4U3CqJwMPWSfGlcc864QeVo85gpQs
NlARtgTGMTM7rW0EGR50grJnZ2Q0U/l9JaXY1sgQcAkYiNH2YWqv860Yx2TLm188
GRONYCi2GWI5h3CKiUe5hHJnD8lvK4BJjVkP7TIjGkZXbHio4syOOUtR7qdLeNkW
03TpSFzg7PtUVv3heisb2a600e1zYxTpxqaMjA/GK4OdBfcH0jZlQgf2Tk/AnGA9
Wn0StJ1UwRmojskqsx/FkIGc4FQI44qGeD92tbIxyGmNH7NrDE/6OHrqlt4ICNTV
KXoHHe+P+sM7iSNUwilHr99TL5mOnx0yM1ng4fkEhPevMD4t7sHs+Z+QAbjRiyKH
5J3wFDU3KjrnziNUHO7SNZ7WBuz/O4w0ss2j3p1MFGMDUwYaL5FhRGFcYuX+fLT2
HCZuf1MP/3H4d420OtMtVgsV3kwqcxgw0TBUhxMHpj92mjOhV6CvM+LEowr/O5NI
m0gOeSp47pFMTGVFgJm1S3tsGZ+vNk6+IaGitni4FQYLbpcwtcepWt1GHGNpRr+j
Ky7O47EE0zT5V6lY5dC3sNysstza0VghyscD+XJN5u9jhhMexF63qzOCF4dugauq
uTpvD1XvYd6fJWx5Cp9ewM85/jNTrWIDWf7Gldo3DpOn70EsEjU2WDpS6MpkxQVz
VBmo6NVxlyeDC/vl8Xd8QXPvyG2yhAKh0+LcOZTePsmxNyC+N9wWj947uN+k9hXH
t095217dJ+C33OTXAzOmJvS+8RWZD5bECZYdlmO4JGy5qIjA0q5gWNCBr0LnQGok
0KXh/ltwfmvXVprt8ES9VqlOj81E63Llh8Wl3kQXTNujD6WwzIjv/k0/Z9jYmnae
8WrFE/FPLg0UC0Hr6727vc0697eAEvpi7bC8XwodOiaUzU+HvKHYQnB/XUtopxWM
TLp6/qBjUfXy88K01nz5PWWscU9DP11ikCMCXx2ItJyt6Vl3+doqtxP2mG/YqGrQ
+t3m8BOiqdgw6jdGa5MEX3vYjzyOi33RhdNGqmA+QI1WAUK5EU/M6gSUtuDROh5p
Z7THUWgQ7ezClVGaUYUpZ36LHqdCqLVGcb0ktaS2V7tfUSl2Q4ygPVIW0qCn2pcO
yjdN+zPVjQlFki4iPBd5nWps5ZocTdRfXsoN0bMfr92bgmpi+syS5a5cHY3IysR6
mCn3P2ASFqpeSX3+O3/Yh16J2dEfpu2qHlA99mC7fq2qvc+6ju126fkFQXDnkVzG
cLfyqMtwcmeJhpn0oY6zsSf0AsVHMKU6ptZJfJ2BXKOfjsHOvqGPPz4/Sd4i2jmK
ZQseId0hb1VQWffv8rb45w7y8b8b2rsOE78M2gTvYR+60cCkXYs69crU/AGXmU0c
r6D3zLpil9BpFzLJixZhf57/oliPkHLehoZG8IOkvas8l8mz0uRHUMMRodQ6LGSV
lhcxVHAuSQOz1uC83+fXXLw2ufwRxj+1xCRnm9GN823/wBvNPoxNJqrQAfeoZDjN
eIfvbYaS0Me8BNoTNVzwB/LJc9j/FOFkftV+hvWi77k+Au2DW1yBV92M1HPJYwoI
qs7v2W8UUXqASp2bks+tA5oOXMmlGv2EmPr5SkVCu6djFTPi42q0d2wI2Jp47Ref
4651aIZxsW/V0vW79qNd7sP01CyRiWcMmS1JBl6nwg+kkFMYDJ7Y0lVtYM/0Omab
dVR8l9i9B0IUEolQk1ySE+NwrbWuvUhbyLku8oyF8eJPVDaN40bI4hncyeZa+xBY
ne5pRrREdEpUAJGSsYjhktm/plhX+1g5eiYvIJXUGELSifAxYrpMns1Lo6R9FQYO
mkvt/vBtpsBs1SYaA/ZzKdYlwsZwj62XYROuYFJ+nTSlcvQtGgaaBWZBWSxJCSdx
HWvKyQ6seiPuM63lUIO9zYiTVwSLr+8zyBBg+fK+/8yK98EU56ibKAU8IIZbC8Gl
wkVYaV0WfDNE3b2uyDCbBw2gP6sP9XG/IwTqwEbzL2LssXLfSGtlSffaHAkgb/9r
ZusO54oTOa74Qj8r0ib8RXaPqdkBhrZnwEOKsUhdXZ/lrUdRZe4YnwovwoAb2IHr
NhoG6JkpfFf1Fxrw83Xz/pUoLYT+5Wuy45KXseUfFEhSSnxeR7YoPv9JfSqWk/8I
eFB2CkJaOqXhjVlroQ4xF6mnMc4QJ57Biji3McRJJpfGjZPpAB08pcgvxA+LLOJ7
f5Ry/OyvmP5klTLjzA1bhWPu76Kf2FuQtIlFaQPYiwympDadnEc46Au1cSEuHmJI
0wFlBwxX1Yye+ntv8mlADRD1sTdcWsUran0KJRz6M+UPs+Td8pkDZbs5jTLyv26Z
O3Z7gCpCyHMSnkcczne+3RdNH4gr7dKGZ8/aM1KZzLUodgeONOfb1XX76DoSiPps
HjS1szKGcxv+ukEIJA/TIj7/Hn5BPCCdXAl2NsUEtTfz9ggvmBFPecpMQnCg3VGc
WCqXW7zqLpWa8WJghcqf5hE1N0wE/KdOQJACwClfax7HRxXeACSzg+uJm4KnVCna
aVsZ3hozZagRfdohtL3eDw0KMhlas1kcOsgeEi6d6sI0lH0GTTd27DW9+wL35+6V
pTOZlxJVIniZgswZ5Ghp5IP8GaFqWRhW/VSEoTyxax3gEn7frpWiDFeogkIiwfpz
27mWP51GDoKbo+7ae9XgeiyIL9TJ82tNKPYsPgojmM0gvL+rrvIdoBLEKiQbK+CT
RtCg656A6q0Do9jtu6OZb4Xpabz9kQY36IdgBVnCCXbyoNhbF4InkrSQpUvvN+Nb
z57ZbfW+sGSozG/hPv+ewPO45JmnSG8cYXBiRNVGWMZqOpZrRHVy1SbbMsenM5jY
OgHp4rgYaSLPuNDo00vLbn1HUePzqsuCkrUmWAXpcxiaTmSXzMmEf3ffZ3fswDxv
ZfuA5LHu+biRQbFGkor85k8Qfz4Py/OJWx2ykraQMx0mlm4iXzde0fJkR9HM2FDR
lzgFd+/TBXQ8M9DQkrzTYA9CQySWrM7t6UWKmlo+8CUiOtuJeFtrSvitr0WdGDjV
svDd8YIJS4mjiizQreexHoKHc1J9sUKjyKc+JOplAxtORI9otMTTLc3dTnt09wr4
WQEAxuGlhjoTQhedRddLXwQgjLL0qSHf6wFXwMfr6likDJRN5+X0SjI7VtYwO86M
ZVNSqjCplH66A4Jr95bbh0bCIP6ORFhmZwoTbRS5OIpTLxWiM6kALYR1W7IOfek0
5zSZU/EP7E8xzpdTxlLHR7Vzeqz72oQyYW8FcKG7GTBPnvbbiz4iGSfw89gwbGmT
j0qvRsgTbDFpJoKGhW8pXT9RPJCKtVV2350c4jb84EQ+D0MDeNUFeXAJX+NO/wkh
4kg6LiwwAYUD17H1kU1BBs6IIg6WCmclExlf9aQ+YdlSasuTqo6kF78hFUaUtYVX
awaNdGn//1RhnoW/gRVwoPX8pnhQgeRgZ8T5/LMCSCVanbH9wI8GF0jRh6rVSR2a
fpFQjxcxybqf6w67kpO5FnhNOMhNBPZEUt3mZRKcDDipMua/a+ho03Vs28pdSPmx
EIUPCelvwKCSY2kyuht8/ir5r3BnlpkzDyV6mOj0ECFBOSQWbpYb+3z5RsCx4m/e
yzZG5Aoh7FrFrlqQkosOvynlFtY7f6A0gLhnlapRmYOD4Uvw41oiDAOykf9qFe18
qtJHy1aHaaAFCcqjpHb1Jvey4tklrruM5JCvyL3zXy2aeRUDgs3tE+d6H+tIhUHI
ezsSvTIQB6EMxrno7BWPTzofVKbxc3fIwsRM3RPQWAyC0zfMH8VPxEqdlAI+GR4T
gXonVIu0PquNcmUAAjBscGwT0/aOWkdAqXTDzgCrvpcCMt4uqgXVMYOAHvSo3b2A
xwS/zVUtIAmaIysai+qhOmJ2nw0SIVNO0Op4VkND0oP0kuP5wZhyEg1TYqdI3CeR
Gq2v5U/jNgxmFxaambYYjDaaxIyQs5d+VD2xF+jG+aQIR2L7hsOmI/Znn6ZeN+4V
YmkQgmSmDQkufifCP7VvgRqt74n0lj2FZyII7gMu+qH9IqSN/48IJF/dhWpNRvyS
Wys7b92d6ZdRU1Q7gtCuejn3f8a9eeOp31WGlKcxa+6baeiEo5VVPrkoLfqtiykr
A4FdMjohuZXwuwkHLbZp9NQjRdBWp748HTY4y/wSccgnbYl/tmQ5iYnQeIJLTaM1
pcARSKz6pshDZT0Aim1vDWzMrUj6Dn0FIOF6vkrZbbWelaQBqbAvlV5MfvNjuYMI
cxt19dajG1Ou1EfVjp6/zOP2Ar9YadL7niQaHjn3whRNzdv4DMEuDF07ckPuo9F4
jYzwxm7RXdfqMjR5BnyBAGNqOn9MhKv6P+3LdPT/I4rDYmPL8BUOBChnSSgPK4AH
pf9mMfWMObBm9CeJlM6EoLJT8+ubytfHTL9NA6w/67E1EzNuY8mPAUwgoxvof8wM
V/HVCbmZfgzg7h9bDVmYNJTe/R2YNAhyDYu1Qj1fv/qsxd7anItnK/fAefca0gxb
nSzDrA1aaliNVGHHgb+2AEkz+gHeBvLbdU0qt1eqTY93K2L6L60lvi5Rnway4D8t
1E9Jga+5V9QAaShJQGa0DRmzlFTNDpnlr4Imf3j7iXsUXL+TvaiYsKT6PODm/9GB
oo3So9RAv0Coqs8U703r2q2XZo1o13jVVwIiNCt+hDwcLBp+q2EIsfaFhy0osUWx
19NIv8rqw7OU/SZ0hglYgdmrAcoRorkK4JZZgdsQGsib0k2YnoM6a1zFFZMv2SNI
wodsMvZoN23Hv5GyiqXZhqOTKKINgGMj2zGe5Smysdz17dUVuIkKZGbSkKA5Do3o
wtxMJnm88ocH8GxGrQ6AHCc+wcRFDK4FIEg01xh9RCOWc2dIdWeBsXJGgmZdDn8s
eWf65sOh7mqH/DgaE7NI2LXb9A4sToVPH15xd7BYkYQEPUPtDBrZFge+QtCNp+ts
32J6G7rElgsDQqKifARnRcJqiSXYQkVQpxnNIMxbjg/WQ4d4iMG0x61AaQ1U0SkM
6l+vMM7cogVzdMhwGLwifZZ3UnpS/pq0qHfl687reTgUSHAwXioROt723Z69k8BQ
2RzOoRdf/IM/9dKL//FMuAe+TDEfIDwsCdiHuomkcvd9MrHUMSPj+XueBaChyH9z
RguguVCIQiXSN8wI4Ii8RtTd+8qMAlySKpXdQWO4bco6pMt66whKztAnTqJ1CRjw
LUm6Uzdrxa1y6rCqzq+wv/YI2lphI59661pB9YWsSpQvXgYmiSrHBzNgCmmjquQ0
ZYVF2NHeQjxGojy/c+NC33QMru2JVCjVe45E6/WKYDiTOSIr/9H6Le/mxotnCnYT
n9TmIfl9qBuFXB4+ZmY3wCFHzxFYcnkLDqxqxEHpKETTfkEIwigoPxJ0cLW4vrrO
q7AJkFOXX3QUijB2PSDK7PItV6lAX8XEtm8nmFcXtRkdkKIzjnu+8a/D3zFjEXr5
4laqb024TrdhHS7iQgJDIEW5Amh2ukHJjToh4c+bMGTb0YPp+t3YUc6N/8ckxMHR
q7+ORYEdIW34t6IY0r2aBKJ1R1amiSAI9LLtZ1FMbkE/u1kGbLXrq37EFC2VElGo
xd9yNBrND0HmvjyLDhe0orJGEGVg6rUSi1i08Ge9HA8KMt9pq3PyyuOUgg3wVWLp
6vm3KV04bEd+TzZEgnWi6uSbNzo0qeaHBys2gp6PF3oEGz7ahXq7LR9pEDXVk+my
qmOIDFaW8yBiz8t1smjQOYE2AOyoE+FKX7jigGnvqx4avBKJcfQE6OBs/vnfBIaj
VtQN0ryH9ZA72o8HCslKdrr/db13r1Tp+HQVgqRpyyxxe6qAuf86hLEnfnnTeYkR
s5i9aGbUVHxM5TIbFLCekEdQHr0XtsZnoRU/SBeQmpOZIthHqKt5Laow5RKK3aPJ
tUEsHplKnKW/bwDgAkOz2RB0jPYADulLiX7Prs3qwZED66fYhvByPUl/yikiMTen
QgM8lM+1Aj7IXcnKbkdk+Lyk5Yy189qaxrsDQLZI9ms4/3dSOphaANED0s36L9uw
96KUq3Wl6/CHERRGl6V4sfOqdm5mCpN1JsrmUpL/m1CwIYOEy0qT7k27khOsIQM3
TIB6qyJvUWnteEGzSXmRnSe+PsrV5Yv/8bTGbeH2KHPdhIbf7jnKFuciCyWvyAwT
vAYaDwsY/EuMKW8YWtsULimmqujj8LW2pBxocu1UIHFitKrz7pnw/qbiG9AZ6wQg
gWbvP2x2vWC9yRGN5JivYf5yWa4Jf8uaK41zNPR/9hZtOc4BdBDaEfZnuGaSkqJm
ZI6ojZeuYhTar4Vak9GrSOGCeKBiGqKit4ufx6OXDkblPqgR7KIm+fa0OSAJ1GUH
nE1IPUnpqZVzBCYvC/cP0Yt7BpFFou5A79vsyqYeqOQPqI06MD+kfB4/uaqcT72O
L1i+6pLTPjJ+j0VgPm5RBnjMNK4LsAPbaMUUPrQRzTNCatGG3a8lmzpo3SCpzhLk
Vbs1OVx2DsAgwzL0G6KR2cyGbQHWLNLwQKHHCG/I2ULcBjIi9HhtOdqtkW2o2dON
i9JiZzF09KPrQXDd6HUPmj3ueYkqOalT8E2MwWdwmED3oeRhAO8p2dFTYGb8MA4O
c5DQR3ckA1z8ueQcHhhTWyg5CObEiNPgY8/qUJlLZLHeQZGpE/5wOMWPhzRnwITJ
bt7hClUh6UG+mYlgRZlW/Rn9cKb5t9LKAVxFfYI75UtjnIgcRm4zG8Tv+OScWx+e
YduAvsSPWaudmWr9H/tV2KwqnRUw6NA4K4KDOFWGDo6OBKxxDR90DCsb8iT1sPPd
FuljfIXQvhCaJX/NNmeDS6teBWgdTnNztoHO5W1d/kybobi7ea7dDAhFiyLGczbh
9nqtGJhKAdFoFmYP9uGKF//b3Qt9pLlr+wcpa4aR6kliWLUPzV6SrG0k33jz5BIW
snBK8H+8j0uVL1cmsvZdo7fNo5iEl2QT7nGdrpeBBBiOtdM0EOP53HNYTGepSY8I
G1XCjaCy3/tp7/RTV+0yhDSh0tfzFdBb1EhJQY/D0WaqD9hfXdApkTPgrrZyF4P/
fpL4tVr8lKmdVi6DGiEpdeFXs7gWom9q6o7SFAUE0s/1rpk/N1kcC4CxAqKPfocb
u39+AQwwJy0wcQx6o+BDYMJxTK0bWcrX3QnNPhuJRe7yshmn9gBA4I0BNsn3dSU3
9E469XPaDpJIoMdj4bunjdTnxWOSBTLMLNN5qJ7dvgtbSwCyp9ABt9ZxADhfXTdD
IDi03HchK+AG/TGob+z7UcbEzm+P26Hb6NLRJqFrDbnC9B6EK7ygeN7N95wzwBAl
vaqmycO1QpEbxUy7hykiNxVonqdaPeaZrayp9B4jzUtKszMBWduMLcjP94VLdlLj
jr+5g+k4mY/xPmmXIujIqAA4cAnfmWYqlzxUXSRCH6l1oA72yyYEIHkk+B6WYF1g
Lz7HIBRxIsOqHRwG/68grpsJfRdWTr9Mprcw1pQprZCsZuQmcFo1ndtG0P61zoLv
k5svezSwNMLP1JVBdRm7pkz4Bq+3H0CDIt66HhbMlSdiF1WEi5TFeSyHOyMRFiF3
wpKq99ay1Vc20iVtU9AaQoKNB7LACEAZHhS8YVYvvNztKVYCxM769/IzzmIsloEt
HViL3kyclBHvO6m/JPoA+llAHmFk5x9ebSqAvHkXdbJP1d0si64MOu9pi6gRjrbQ
dmIntAaEWIFSY08VVPbuqb4e38/vPrXezC1eeoQK23+nbpMqMpvzrv1K+NpLuiFB
rlAv+wCkBYvsX66D7U+kRPBRr47hWhycWmB2cKs9DCpJMRViJbKBlZBvsHuZU2S7
RzXtU/FpxtDscjzlMyHSwNZ1eW8y5dV4URuGnY4Als4vec+s3mBkNYJmcpajOQtD
UW55j+p03ijx+aQMyS1mRnZEUEfGN9hxckjNh3WWp8RHxvTgHHV1LzTrSEJg/1om
vvh36u1PYOMvpy0hMRNIiOxtgSy6qJmfvBmrFKukoCiBdz+aWTveyCy0pqVi2xfK
urw3UIrP5TPgHChWemYgpbtELTBb9Yy/PQsklAYEAr8RlgwZGp8uUBTPhnMvEJXn
BmBdrG/MsxWlqa4WcJWf5QsEpZmAQbQjuw0xg6cIJuDE2YaBRTX37D/+xYFkwxtD
dQh/8Wfi8RUnxgVzFFZGVxIPdwqpZmSeFSrTW8fhxGX/4KF49P1PgASfY3JSZyPv
OZgrMLVbp2/WYgYy01P/mgT7V4jNlY+a3yKpxP3RZZdExc5Q5Wga9oIaBgHQ+5eN
v5BOXz7tujJtgesiTHjlznPeKCxHAIQ9GovGxfJS6ANLH5G+ZcNA4eNJjHv28ZDv
4EiYr4CkqggH3ju3oq9RJxdMAhVsIeeM4rR6w7vJJzOJGNp0ToQT3+omSycdtPWH
snNUhcQvY/kzaAebbWDSaxFnRvDVvBFEML55EFnsuXS9ShHQjNkrz+0A3cwIeORj
IP3s02EzWe0gszgk4utk9J/+QP0kxT7qcjhN0m3KGdqoKwLcfCzVmbeC+h68HSh9
RV0Ot054y+j8bj2lc5FBrKVs3MpQuqIxt2RTHwFA+02gi5LPPLp3ugfiapgSpX9F
8e4vHV0nZs0eHW+PShTVOxlOAjcwXL4n6wHOtlbbcyHoY6jATMDxvHiKVVLz4C8e
dvHr5okeOEz7OcBLtBMtCdfylA8wCZ6o0qnlPCzG6Sqw3Z9qdEJvkjd9qpejUGgd
+V4WBlmFqZP1IfrPVJFAgAIYNlCmdJyETN9J2Me6dvtFtGifGlrxvi5ushwibNEt
tUHRoaGHhZjdIVtKmKVTrVVGG9DVrnp0c9VeTTuvq2VXN9shdZbgTy+rGaw3+xnP
DBSBjHZqpIv35YwOfO9YMT16mzrZzWuYFRqksVzyvpWdtd479ZtYoBhJy7nybrsM
RqSBBTCQ2OKmpcJb0es9jMXDwl8eHNS1gi3OLpIgeceMXTvdPopY/zqXaFuGk97U
oXNj5+HpZHqPiiBISG8hFPsehssMbh2LNFiCNzmMOg3DQhcIDDUHf0SsmYVQviih
CuWxQEA6bQyGDabes7isujaHmpE0jWxoCCrMHoV5kA20WrboKG6AvQxPOCMOt57/
h+dSM9dTGpoT8zseCLeBXr4GCAAaEs5wif5KVGrLuwHAMiFQiii+tAAxj8ZbCsG5
7pzb5aHcB5uSfF1BANIDDhyWwEDmA5ls9wylSQRQJx35Eh8lI5UEG8ImA1+su6X8
EM1lZqgZZq5n8Kjovd0Jz5jqO+NwgmyKF7ZmjGafwK4II1FNpWX14fGtIfnn+OLe
/3CyhXiDOxu/9J9mzqUTmxGcGc+bjORiYI4NoyP+nRAwJcLGxiwuCoinn3XuY8Ap
m9KnJN4HA+PeIChhs5PWzgeGFhOhAVYqo1f2j+ktOezS6PfyotZ/DvOe/RhCUwiP
ODAQeS3Bdhm7l7o3ZwFvj9ZiQrLfDIDexG66SotYqRawcG7+8pVrfqI7jb1325j4
VqfBznCNjVKdIZlBssbm1jQnBSNMobIQGrgJfA9AONTHcPgWsW2zWeGOs2MvFUg4
YAdjV/QfEXf8dDHbCURX0a5PdO6K0GCfEYlHs/T39vXlBlMVf3033Mv8A4Kr+9yE
C3mMomVAMwW8v5F3FEAUR6W6AsK9R5qpjbvYLYIfsTWkIgLHTrOPad3ql0hggXZF
/BX5uT1wEPrq8LltFnpd0LvnTWbC+0mLLvkguLf70XAgk1x0xOEVDlsJWJT8b9w3
UU8BAmjS6OR9o8tuHtEnBvOL5wI/BS7Tyt56YZyXVAnbV+sZhVgX0iJ4W8kSV8lI
syZ4PcOXif3TFoH5eJR856dfHefTz9tAlvOg/cu+pBJ6dxDAQZgta/Mcmtomhqv4
XzCyEa1kZxoX9JRHuKQWQz6Q7A+z+pkJ3xvYHmNgaq04gYREp51RP0bM/utxI8Xq
P4kP3lZoHPCh+LKecCOsOmTSzKogTB8qwCx8d/VP2jnajWoRJ5B0sbQAJKq+mMur
hnVXZvmAyAptBoBgcUjrnWInJzfoHRPPedSrAeA54hynxkVY4bIhFSj7sf0fc3Ja
bbpi4Na22hiIsiMAeb4P13bez4IVdzdOPc37Y+JR55zlYjp6D/GQo3KDWl5MmMlB
o2J+fm3lgqZii3Xqg72H6YjCDKn4FWJHWVLv5LwF6Yh0vcQDfNuL0cMp0sepmGNO
6ipGPBU8btN6dGIg4I9M9VhE3zqoXD3vDCAJExeOSfWyat/kH/Dcpw6nwNz9sru+
bHWnTqS8CNCWtGslMeL0NIHB392oKAx2C6S9MvpXnfDSraiC93i3voSM/x8kdgtZ
2ytIy9lYewiL4rgunoqOPJSEQH/kIBIkHoXiUN9ECorAOsFcIgvtwUJJi0zQ+5ym
WMnWE8OzrQuvIZd25XhYHj5VHMg4e0xY637rBhoJ5WWK6C6mVfMzJgBf2ZSa3+4Y
DKYMQ1wIu5jO+YiB8tGUGivNltWRBOpheGBt1rM2xa+ZOnRWrlEYnsd9Ar2x1nIR
XcM1G18WjIryV+9VgXHcY/J8uvspKHyJReyI4NmIj+uawNZC74tVae8gOySDdP/C
/ENuERciXAjP9GDYM4/xjhRRwf94j6HrV+if86dkT8dEspvAkfW334aK42BOwgCP
hFIZdlh6L1ah0/2QIw+oBx9e7T0xtcF7JkXmfs/5tW+xIh3G9uy1UXK6GEP7QLy4
iPRVEERH+NyU9a0DW70f9dCseKiojGNsBCp/BrMDn4UwRsRLe8wtsb9YX6Y3kpiv
7ATMnjla6vU6gtDaxU+GK3Gi+LlY6g3yEaSaB3en00M5LF0uIw1kFwbW0DTKJQCy
2phUi/bkC4XhXxHM6pemuaDuyvRmTUs/u1nKVmgn3J6/xZuPzFWnGC/4/aEo0+UM
9xskvXsVBSicX0ynuV5P0mOyWuXjHYBAtWDhM/ATqlx/QYdR0xe356MYrUeig8/o
v0tnINfGXJPKGPTY8I1mpHRQ1nEJ1Uz1iW8v2B2tFzUEzGg6l5QTWR0fyDaOUFK8
DAPfDkD/CDp5Z7gWY5n43xIopYPy+vS2iKDyhedhRCnhHjjTxvJ3a4hHLfgi+9aM
rX3I3VTOIr4L0AhXks/Pn3T9BL68eL0ncPUF+Rhh9Kmzekz7wCVX5E5mPQ+WoJEj
J9wzRkJRw8mlloPjJyrn0xJuTlZZUhlu0PzELUvrTTh7nyob26YH3bf4nlFZ2mN0
/eR4l8ckbZ+Cs3BPAsa9Txk2hge92w1MyqO7+NF+GFsOnVq/emByL6LQ2rVEZdXv
5qwq5cyqVV9Vq/w0eZr2+BG8iGNCEWNwg/2Vjt6qS2+7xpGV/DXD5aOfhsTRjIxI
yA6vyTQEjEDfpcVAZHL1EwZfdP6Gl3prNS5nzS1aLCyD7V+cgc2HDT4iB2ng/TBh
ZQrF3G0uqB4PvZuw1OWuoCKjN52W/89y/3Fp/Rk05PMzw9xfr+81hVATH7LV3vl0
VPUmzFIFwt1XoowTNxdEpxtMA5ITSMTRy12ELYZdZf9R5hMDzY3icRiEXtgFVNXC
Njkqzf4GAkCOIhNkPu37r3sahcExzHKGP0QQF0o9a7Okx242C91nV/QN81MAbnx1
ZGB/CkB3kW5IrUWCsV2n4cmExU6pwzZhns4FELiJkAS1JV6Mb1G3BKP5a6V5WuUJ
CLB05+gUpTZYSCOe18MXUiwDCQZisqeLwnEVp07KWlS+hjUMrYlDfy8dZrxIMsR0
A3s4e2jXcCZ1NrTEH9LXWY+Vmu/jO8xoCqy+b09bN7bIwHZatTlsiIuhSmm1jx1m
VnjrkyffVo2E/RpZLJ5oszhvs/ID/LyQCAjesT8Iy7cECUYrOhS4DnQaTwHDSdgK
lXOGasZFQaGZ9FfVbV8coI5P4kuHJL1+xkVEicUJ3JsHINwyhOmyotC88Lp6PNcp
vDlbhqoEAbQKaQjqLCM0iJ8C1rXJQuHSABAfljktKXmTzNOy6sEHcYGtNmXGdKB1
aIDRee+A799faB3Pj/qp0b/pDhfMMD9HS5P+PeFJmTdClOPByZ+GeSvyOiy+fFyn
xTFgxZwaHGAmdvFRSpFOKIfOfZBSZLneM+o4tqpypd2frbozfFeMsK6hZyrkSTnH
qKi5j1DBVGvTWAYtt5fNgW+nhQeFTb8Rbafd3nZF3qig3xxVFdTFnpJ9y2iSaCJG
NNQxeYIg/hbXXvJ2G+5WoJhMqfhwg0837Fto3XmH/2UUbj7scHUMDrSyqvj20xsd
YTqMBw90CVDrBcla/cVYKpbTRpymxgHIN74yAUyXdrPWr+f4rHsrLwiBXbOhSHLq
UQgra+0dEAL1tlk+h1wVHLxPwdN318NvUNOBmZ1vWjWM1XOYJTy67rPm2fL5l7vq
ijkiwJJZmhFoZ9oMZ0SvD1l29JT5wVaM8I+iJCXWpAjJAV9QWYAhS3O43Po1+pBX
7ygW0UeEE+cH6DtgHUBtkEEwqxh1zMUF07gzAed0fkTviYUuifOQR2ifT6lytsFb
2y0Pvtpx2DLc9SLxYc5dWE28Gq8HHGXX4ZpY/btwMj39MqD0V7z/zRMWXgY1t1qg
Dst/bGVQOqZ6qppkbx72N1fifKTqS0AzWXlRw9q/YhohRfebYwV62V6wfhTD9bcx
t8gWBGePqaOhKsZLOQ4VG22WF7dL4sYmbeMhCj2T3yB2+aNXVHVhts6EY8tVkk93
+4IP3r6brycdcZPv7utAbRy774uGQruHVsXDQSxw8bP0+8a6T1yN0XFCp+bsbkFo
LKY+X+2vQG+fbxD68mx/LErQr9AygPR4TPoOkGg4umHygZIoT41FkmSNaZ5FhhbG
CDYcFZudHSWfssVsocJNDSrTJFnTw3LVDw1tEb75na+KSPkx1QwLCZsBV/ZF1aOA
7jNwijJcqHX/1JxYyXXfnyF/i4pV44kJNsqQllgeDQYmDyf3+PyPVmZaRtWlUI6n
4SMu+HlDHDVFmIE27BpHzZO4ziLn2tR9IHGnrIZdiS3xRZtXFesFKkI0Alo1mkD0
yHXhE1JHP+u2bjsZyOWcscCcgbsb62v3wquP9P6PJTKOQcw2723oS00HUzbIRfji
j/aXw4k+BB2128liwcc414rf/Y7s9WPQE9/fhFHqRVn+TBnLGTCPJk58/ponJBEH
OyLV4tv/rNbImxVTkFORGJwYmx832IyQdbvjNogtWGZZeank1ig7td3IznIA8C+K
rcOVuqnz05RoUgPYgk/z9ZKNOl4H91wURGyS5j9ndneKqX8YxzFsIn+/rvM3qiQi
H2FRERFMUO7I9fvVyKaNjcDq81tOh3TVibh3v5q5KX4QDcwcCBRyKiFhcP0PXxIr
o2DC6V8Pz+RNc4puR14wFJFQj5tQZ8mjIEKhxCkZ24Dmw1Rd/hUrfP4/XEwsMBGe
cQtJacXljcMpyJVUAWFkX1SRFUWHb2MDh5WNO+w5+F/AY9pkwgJCR7xkN8+DkiZi
Zr7TedwiZaZ2rwpuJInVXgGP6DV3CDuff3o7uQmhwOvmexpuJGHEIs/+a3DvRvvU
lG4IgzoXknHtf9plwKT01llonThWtKSE8uKeTykq87mlBvLVv3NUGaiZoz16HuWp
rdhNN1TdxCmZ7CjXzeXzTlLfRmLJ8b+kEVHHcXsdk9gghCN0f+1IVXvkCLVvgHQu
ApLa4bR2ke2fOWkHzoUZroDfULCMDCrksMMmlfdDbLfKAzx5smnFEGOVjzP/KDbF
jHf4cQDXFVxsNC+qQ19XA9IQeqnQ38zI72K/PEPBpx2UtncPtA/9WyEnfN0KnjAv
0j7MEhPxFv9JzkeoDu9x8rJQlwWUuv0snQHoQL2NMHzMSaA7iwT6hkmbWNhihXrj
QhBjbI04XPE32nLkuxPTCKnrK2uq0QUGmyVeuj5sr+fr6mH1yoGdp+Gyd1ZJVWVh
yP58nR6jNE5CknDFab13A8KWNpf23yxDLGPEkdkJzlGH0+xt+9UhWrsW8vefxxDm
RB1LiFL0R/YIhST6tag8e6vC6VEYxqvFFIpYowPqiDvwRbhDkC+Mfxjv7NncrEtR
OtqHNdzdeGe7Df5Va5cK9t62ZdAbwI7OZq82KSYHpeARF1+pms5SAz8E1+A8Ty/5
uwszbPvNtINFVvyrKwOphbJiEQ9nKYzPsedgDje//+WCrtS3x2mNNsO54sf0OL59
BRDJZHB7tpQ6w+W4u+PJ6JbvREa2KF2XlnlY2s0vvJfk95FbdxHsJsBvUZggeKtb
OpHRhIO/nLfdaGAUmlH05dVYn56XXoHcDxvGhu7sbcx+fBs1n8rZsesMprDHRfXq
x3n5q597LsAk/gRu252fG+sqrB+rPneob31F3LHT4WAGPOXTvUbPndjB/Stad1Zz
eC+2xiKr4/z2pXQwaaKmjx/WKHeYITlDukj66Sm6AXdXVJAKSmpZB6w7dO62fqgz
eLIzS+WzBGFiaGQcMS6Fu6lhhJF0gvLhcjJrEZmfk5SXvav5rPpl9+C1N4wE0UcH
6PHCtJRnrIhjXknZVHbkr9USJK10xQ1q/ArbyvbBp6iIB2qLnWeKq7KhZ0RW7iZG
GUYFKAf7asA7h9j2tDW7GqAoO0a1yXwoZdlg3R2d1r26pGSx+ds44UHakVxIJrWd
csyTWgMaKp18X3OitOUUmF1ATdYPaILZaWjc/s43k/qKbEowNDSkiTTSxNvaOkcK
3bVMs9mOV8voav4GY/IybDJ3j3u927RbeSjVkzrpHPBVbsrRBc/50fx+pjzqOnu4
Dc/vdmQzITad19h+HFrObmnLdFXpJCZOti0NhhNl8nIEdTMNq1Sc51ao+CiG3eAu
9kAXDdiKCGbtTAoEg3Z+340SIQ0/rywTtSKpg3AvCNC2nycA1RUMjcIgDOLUg7sS
JeXwcRROKkz5gQYEVa4hMgRrl7Jxqx9xPKPDMxFZF16AoDQBj8NvDIKygOFQGQ5g
ikZKMpl63G5YE5vbB+6GLz1AITylP+iG2F3WKfo2AAgyzVuF+vGEFIjhSrIxUTp9
nRmUdS1ANBAl7D5AF47Ms7SYVXsRc+gQqJkG+wxt/6btoQ8MJbD5ocP2HxZlyFNm
Bex/Puq4uBItAVpdKh715J0NunBcLP/2L41wdJllBNBginxRg2hgk6+ijMdAV/um
6IcaJUEJSajDtw0uZSNgiJgQ/Tj+vpqhkY+30uK6j+E00UkB6/e3zKJygZky/07g
RlslO5iFEjfnBhuWAelvOyXK0geEdzGypwcFuhzXH4Y2Ey4ChwqXcbR8uL9GDDmD
O/5NxkPopfCVKQeQNXBGFUM9QxZJBhaTbp8JrRc0j+PpU27w2FnLKuAhPvzLoLey
5TOKJuB+vqqYi8UdXKRtPi3vyEkaT+zmzmaX4ZWkmtaoUs6XatNmQk0yiba8wJhJ
w8CPUwyLeP63bOvKnEWZhN3yYujwZvjJitEQvUwHvXijv2dxtw4qaCnBfNj5HZ/q
ZsAbhni9soloW3A+I6jTRAwDf9SRgJ7cWnFzZl4zq9PeCpwB8s8LTamkD5vBbeei
xixXrK7br/ibWwhgMqWXCVJgCsr6muQF703N7ciimduKpTXqxF9ORFFVwLu+C4tM
6DlfAhitZW5cIsqB1x5w1U06vXwzCp0NyApzpKyMK1cNICbU65unnj/xQlaTveRh
KNLVvkyYvv+oEXG7NBaMazNaiW2x4lq9kavp/dwn6nOwJbwUCJwVcx2dJooXJiPU
BYopQSWwtnLM7Gi1emPSf34W7Riq/dbQJJ+dBLSAphLFM+99XuKfulAOXL1Q6ETl
y/JriM14JACYdLrAhCgO+wnXhBP3B90qDyXCGnkvcHAsu7xy3sBUUZcsa18+Jd9H
RRokhpQRg0pqAmJ7krLZeqdUV8KMYrWM0YscPqt/wOVDmISjRxBZGiGUEG5g9LoY
yttrMDkwTTLGh91faYC1bNouD0IUIQFIlwpF210/SInAFqcGWpol025QRtu1A0Xm
RiNglVJheNvZ78iDlkbsYep0zR+bycIL7PEbaRI4SK9OG8bbQD5tTqqpY4wHJeKG
RmXamGqFnQs/l05zp1RsePVm2QVn2O/n6I0++p1NHBdV2WSY7NqiwCOENwuQLIND
/XfRpU/Y2h8BLxqRlsXA1oixB4d932mc0k2M+cvDSI1gRwzPzMgehAmwXZJ92TO+
SakoMlfw4ep4hiH2wgV6LSsBjdhFWKnn78RSMBpouiaArO9+LoKeDxz7DT4lVcLP
VVpGewQENnTk31HYBdKp06ve7AQqfHF3/6gQo4JR8ZWE98/Xqd3tjhMiFBhNXRBv
zBMlxnqfAmIaN0hz5Xg+z73gOEM4RUxHj9gpVDTbwvEuqNJ209AWFGWaCunZdXWX
jLkVJeHOk/kibZSzZCM1po1CiTFvvAPh62Gigi2rzvUdrtBbZH7S/cfkQIM+xe3A
7f4tGt0o+COCE4bMmFbkbK7iqgm67sV/ACrXGTGnDPWsvd0XE5SOLHSujuGA44bu
tzg+HLcYFAtPvpGPamJ1o3M600CT5iz9m0gubOy+3hoSJ8Enqshl3tbA9KreAG5F
Ka6mBKrIe/Ti850FZT6PehY3I/eWzLxLZ7R/tq5ZR0H1hYw6zzUadFzuyoK5VgYO
7jnkiPDat7tZhc2C/Rwod5ebm3ZFkfPXtEBEaHUu9qfLlnC2209eb/nphezoCwF4
5+ZcScbTX7+R8JM2OtmEiHwQMALpuYzg1iGuiT77ibmEqJnpzK8oY6wBae81fqOC
84ZKZo4uFAKCj2HHEsfOmgsFx1A7AA/me1rUTpUivmPxeJwDzK5IQi5o+60H/ed1
XPNUWXKC3FleJLlXikC1Yecd5zADH/K9ubUOu5X21eOJT/rzXXwxPe/rvpuSrhX5
IWvd4dskzFgL1ey6I+yWyojFy6x5xY2+IHC0vyCrKl6CbT3nwxkYxZFs7lvNyp/b
Wn6YOMxOXTorKVQKx4M2gNYqmaMXq5oRJYTwISul8lfveUwT7yvICBCGDGseBDHZ
nsYiOtJP8uBDdcmjUxRke6CsOnfylcW6Xuz1qXO5jtSwFXvLtfcnJ/52sKzSZyLU
xTCIfsDKAAjv1cJLz2Dcg/eWEEFAovbmT9+9Flbl91FaG3XYzqF+fo8nRa1DWWLx
o928rwGTug4Ditao5GjgdS+5cmZwymA6np83pyTxOi1jjsJjFoWBG0oqAeuS/rvv
0p2Ak+TKYaCZ++bqO7M/xKycKDZ0uDd3AZqe+YBeSjBQQH5qwhKgun2sIGyQK6Pd
dvMNIBUPT8cc7BwwrliPJAU5MnEpBTTZFjPmiFf3RJ4wHfKV8Mob5wjuBRpsbkpp
zhcZxKFfqYw1vZLuZq0qYlXe1kVlQtqnDLKOQkI2RS4PznYdi2gn/F3+wAy9b3lJ
1RDCemUWC4Q6HsTjEN9xc4jRBlYAYAYG2RlJxt9+KpqIHj3EwE3WvceLWU+/92n8
ybYqoyg/cYx+acJmRzdX6p5DJzIVXqy5RPBacv3Ynu5j9Z26pKyEDxTh9/p+vzJx
z2j6OqXOpR3Yu4qN3bV0cu9O92YmjHHc5OcKEx4OvFlUJA/ViTYtNGEpd1nDcekX
UefFd9I1rlQShJkh9gaxyJFKiwdjWlqa5I6uCRxqrZZaRnpMmDQXcvwgtF1LoY1U
eQ8f/9iJExEUPC+VdY3rTw8UB2kzLnzKCG8rHiQeNH7SJ9auK2miROKiO9rXHySb
2QNNVWrP1yB+pgGutjurL9+XCTHwvJB38f3tTw7AgQa3iAiCD8OuAMjQ4eZgXjq7
mnNJ4tg5zNiCdPNLhlNgxaZLfhy+LskkOxdnFHCV1UWeSPQ2ePkvg1INR/UnNShL
2gOa6w8Mh9NzS2hb8B11ZkFes0V5OcFebgkbnB6joKXe6PVkgZYUFUPI9/spkTCw
K2muW+BOZ7gOaadbFUJ6qqf0bgNSUwE/JusKKN+WtigirwbwRVjDyIRKCQ5leLV9
nxQCwcSX0jNFTlIaVfcl4eumhuEwOmkufYeBWV5Y9d1XKoZCErtrwxfqrlfVoA++
3nzaOT2el920zBQKNazaJclrDwUoKNvT0BCo4kgD1LM882sOanuqQwyw2S+QKJUv
CW9NUz/FLYn8F+IuHxuxhuuaz8fWBDXVoSzJbt1T8g0dkiZ7IGsZvJqunrr4x/kz
85Oh6PXHx60a3DTXKtNXQ6htMXU40x4cI76wyEskEagmnXiY+81lQ8xW8sT6Al/V
4l1Uwgx0Fundu07OjOh8CO2qKMSUfY1SLOJr0vK6bb8Q/Dh80vjwMruusrlJSfuH
pQ9+70k7ipx9nBG1nIinnsaPh7wjMug1zKQeBliw1QDeoLsqKd6XOn4Hf7NAle30
bF4Xi7DXdKKpe4H/TA30NhjR31DVGjWK0eGloguV+zVKvDV0j87JpetXSxd2+AlC
lYpJvwVpsBlsMHfwUjczI1zygPMZH4XZDZSHVb2hxxPtgm377TVJnDUep/HQ8x66
c84NIul6aYZwciknoojBWQ+JrR1rgI31corfxs1dvIF3Nu7sTNhwJCy+FRN85HWo
KsDaNSsA1gXSH4SzDQA6uFoKqgx77EFdmdslk84Kabl7wGPPBZnADALtU/aiUJF6
inkUNIqfJWfWwV15jTIvNcM9HgoPgHBrHLZv4ZhQQAaTYxYAUePAhQG14cjDwLfU
yBW6XqJ/en18vQsByG/YqdefXZSXcLjAIgtmoFmKtEkhN2poo1hIemCCye7/k9G3
NlAWSS03BZpJQFXTRz9VA8jmzVsf1QJ2R9DzSpyesd0jNUg83R2eB1Tjf6i5kwDF
z6ugFZVZu8Q0Jm6iJ6jfT0roskF/UKqy9za24yetzR2rZc7U4FQM4WnjdF4P3Y2a
8109GVY/oGheZVqiITznhSNzBDX23OOsqkneAmzN4v4RaO0F7lv39sj5MhlXTtbo
HXf1X0afMyNbMql92pK/R0byKELmFfHYKFsolWnCacq+9vR6QABj1zw9xUGhOMzi
y+n57TajNIXnxOLoy2S7gOM2/wnM7Wgpo9p3OlM73FZZN/K8jqsxJBkzv3LoAjWc
QdbISr6Gh95jOj/olkZceIW/rhrmt+kKYnLl6CH7CcXaprj/L96ckMp5rvZtIbax
lSG8az3U7rwmFnf+ddpzvqBzCXmYmazhTsHVxUrnORYibUJ28i7jZ1BLZphmcln1
SajB3X/U8Z9bVLlHtjfyk3HzLqwOWez122qFzLEK4UWU3+a4BHAHui3gKqOyRMoe
Bm/xISKyqUPKTev1iXW/JLZ2pOYaCDlpwQoU4FMlAQxz2BpxRyAaCBvvZm2J6yN8
pxmuAX1owiKSD1iP+9tskJfKRi7OAxpRZFa3Z3aZBw55fWQMQXV+KomF81ZBFiIR
tWZn/vZg4Gr8JSryQZ8cLS/zZr4X/XqtO1SnKlbP+j9k7veWGC/dqW2IP9xGo1WQ
Hwcu31O5xhUGdKh65WiqzwUwQJoBEn2atIN+vEiW4cpshqTlKYSpB2vJUwvqyYhU
ZQkCPflxCWLZuWP5oRbhUXPwjyC515JzcQIxBCD27aslhPEgNoRKjv74AxTK9zFA
cMm1aDU2jRLpTVIL7rRmOIRoDe+ih/3k0NffWSp402K/6UOVia3ErPFPK11+EJ1Y
5R824VpCNdkEMf0TW/ooZUOH2ea5bGuL7cQ9s+E7iFKCykOeLxKvt1FQ41zXZW9c
8ExTt0z1N+qauz68PLKVyDeVdFIR408pnvtu2DBJc2x1bNna8xigO7v5YTmhWB5m
vW6ATUEPg86Zc2knAaR83OmdgIBoxkhqqq3buv4EJUX+4qcPe69ovbYpXCvh+foZ
1Sx23GnCyQH85O4ruwlw1qc/+YavrjMTLTB4oaPktgP/0bh+d0Ldtgqj294U04MP
9Zp3xJH1LGqzz2iAZTHzt/8FBSVMLWFlitoS+UX09RhEr2XMR675atZhbx+04S1s
KS89kYD7W3sdWXNQYbMK0JUCf2lyz0S26KjcKXdzXYEiO4jxL5Zj8JFcDln3qPYS
gjMnb6KjJKa3IoOnCqWFagGJ2EnRwQWnXR09RbXPg2gaZcPg1Zg9lJ/+JsrYCpA5
e0QWpE4bT9U4woDXah1Yi9MueGjTqJcbHBg5fxdG1XOBZVNTAVuOWVvGL+f6DLui
xMpQz8l5xP5EZnM/IBijHGhPwnVIyQsgrfCh6U46L36AAtM2ZvWKgGyHX6MexxnV
ndGvq+/IbXBS3nXBZzgSj3Cwg3z+g7d1tZUktIfpDo/qB+U+Gp7jQ/Ogr/xyY7LO
74L/vzWZE4Dy64aabpJWoiULkiHs4ZQ2Dtq1rLDbwDMHVVJzFkoQ64iHhHh3MlHh
E1+k33Ln/1L+R7gADGqZs1bwp3YsmlVK1PbaEpJsaLFJ10SN77yNkCTMeYxkDiqf
I/elv+XOpRYQ1+/+fxCxjtSy6uFpVGm/tMXu5zprpT1RRAlYe/A/lFxP8R38HXFb
7NkM1Z+2NP7u7jf43LdJzIZd+toSsf+QZQHwRHZhJ1Vy5tDojQuhrxyirvaQ/+bA
mRQy7gCzQxptGVauKoPBa5OPya6m8yKJE5kUMspKm/VLr+zpuhHOvl0SR5npB1nk
SKknFqxVyRp6RHfMDO6cZ2HHL47GYmO6pDN1Y9+ke92GJbon6KA/Zh/RBCtMMGrV
91PVSZN/j/H8cruzcDkER8uY9nRtFnqIzzN+k6SQV4QAcHrGRvY+VgYWsjzEsi6Q
F4eLKb9uNhLfL1L7wxmQ3DsFmSFX0TvuosVJPlOhpC/OBg9D2UgZuk6baXI+y6Oe
WEb1EJ0laT3VAMfnm9HK8p2ijA02uAeLmdEiATXk5Aq5Sbw4ovpJGyhxbHlnGO+g
nUijr9BPqpOKXK4KZExVF5R/QrVzUX/ZgpLUBVKPW4H4tQYYMqAP0ttAEvk5651L
T6yuK/M283qvmpcx2BhZrCC47upwe+g2xOlbCWYKHuIs+sbbCFNbLq0DWL6eGbLW
aaiHifhwB6ISq9ssIc0krrIYYWiAl6ukcTj/f/XV9rY7j5knL0eSdiTSTuId0SNU
UQ/h9yOMabImE4bzSIGglnOgsevfbR6lTSXo+qK/eEvyQV36exqYEe66doy0BP8L
o6hF+rIHGgwI1n+S/GgslWl41/3N+BlZ4VGhqXbCm9V2ID/UPcVRDH8k/Pxt9rcI
HMwffn/aCDGUbv23wH2p4BtaKe63qNhcysV9NC58Xrx0nmL0Vi9cUSY5OHUE/39R
Wo2vz6EV6aqIRF9NNIHu8gDJqEtrNJ9uv+HzkMILbHm1LtDU/QrBDvXTE3mZVnDL
2fOQAgl1HXBowSCuWwmpqa3zHN0GS6+FtIOBj2bx95nxJgLHm0KjkIkUSxkEwPrJ
TR6dhsUk+LcfhDwrpJSPYQr74eIZiv9w+qbLz3YZ1RjdjWbrVflGyPh5QqY+t25e
uHHQgPSQQhWI6hPneQPzDgtDegEeibRRznVtyzJdCRahCo1iUk2by0Fd7q1Q7xSb
SvO6tszFnIAMzw4qQGqD6auuPb0OzkaiWStY/1SL8lgUJeK3qLvl+zdj0eoo2t8v
S1l7JCu9P5eZtDV79cdqwg5H7g4BrzOhMexbskU6yybtRp0nTtrwvQwxDhpFOCbH
G6G0RZVbDUrbd6NA9LBc45ateJLnfRCyTyg7M2r6xkVnKWW2flp+VTGV2GjhxUzI
SDCrbLlAnOYDYaZkKG89wr3VE5pmKVBh1gPN1jMhZgygZKQShZmwQGTzbFsYnJXW
qULF1oM0Tu+9mQLjUwBxgUVlRfTZjnjfNkrK43SQihS6OUwmwnw2CGsKZNOFw3dJ
aMFja/wRQfgPlVgcDuVWfcxoSp6ePpZDdBBmbgUlt3tItYSCXXCXnj8r8UqIbe51
bogKni4MMLPH/ae7Ad62mNPIQBV5bldZNlm4qlpZ8nOuOvnnYsrVD6JSfiRi5HVa
50XKnZcPhXqRZe91+OU1BvBtRIIeS5EEk0NOMNnKnUvXcZdHeX0430ojEUlAMZhO
Z8J5JeGKzmxwuo7GKIeVHIf/2aMqb0q8LSC/Jbe1/oUODSRLhMn/PILUdYQA0pUB
mBZFsGPvyZ1Bk+ZDMfGLwfEFKsSosBfPKMhtLqswIK8b6aW+DzrGv0Mnx1n/WtvL
BC8gGidR1JvHGFaPEgKeZ3E7YMgBdBdU3WoDOXBOhjoXOEzXqWL4I6kl9ICmncaI
QNmwX+Ofb5Hy3zrVCsIHEgoQjBiDIpV+4XYb0D4T9nIk8I5wBcRN4H+WM4fnW8dM
tGiD3UvGIUNthpUNM4tYNa5jVD6R6TlAoVDoOHsTL8Gsv8LnI8TgAnI/KKijnXJR
z/Q7tz+vp0XsuNVeb9YlM56wRHmo4V+d9rgfSHuVtRajfUtMFb5/mBzKZUxyEsit
QbhfFgDId7FbpEzdKxJ+yB39O6z2mGiXSbG4qLwIzCz0gR0UhbubmUpMDwI4kEsv
9fuB5zrc25iWl9pPyH5Ui0WBZg0gUmn0x7pZUvj8lqdCj7pMA7mYhGxeVylvo7EL
/JxjwGE3IP7pJsq7RFhh9ByUfl+iCIEzoIFawFUUZNPinFaf5Uw4BpdowvUp+PgN
fOGC/VmholKb4mhGGtLYRfWg0XGegD3soTZ+ejBi1VtzG/7D8Qg81Dj0NsJXIe+A
friXTBQ+4m85olCGynomHT7TnRm9+V8kMpPdSCkAD1PyIkF5Fj4EvndcSV/drg/G
u8vYE6zcmvQ2Nyqk6x5k9X3aU68mr7cUl2oZXkXFZDE1W1W6aqJjsrlFxQYjYhTn
iNt9At1jPVKUsEUgv6L05FRF840lBz9TKLZpvLhnNktdkgd53vkTppD8xvxrVBUd
OQ6S43ILKDGLzEBof7/1GxN7CAY7bhb+jZ9mazQMtYvs9oeANQ3CHa9d+9iXgXj1
C3QBTWxDN6tiENwRrvF5PI4piGYzquvNp/KEaxfoWTCdOhG5+S/k4FlR8oTS3efg
FpjAZT+TE2fz7LPH0icO3w6FPHDXx5fplKGCgBKIbz/q594yUjMZMndPR+PxT8ud
5Kb/mdM7vJUbBwLvAOaPeo7KCrrf3yOp77dsCKg7AfA7hR1Uwn/sIcaRivCH0bmr
CAWjqh+a6xJjCzAj9ePbKHA85w+wlB8uX9cyL9SZRYG6AY4vncA7GpX4BgjNLpbl
cOMAnsPNi29G5Z8hnWJ7HSVjBU3kNq5H1AoDWgscEyB1f7/b2MCQv+yiFw99PUWb
wsZqeMW7qoLkJrmkORbZ/XRj4EanU1Eucynk+kvwHJRTREPSXhu5yaT8XiWXR/IE
tduWwGD9b93fnaKKV9rGtRG9HXiGuWyHXzM2+2frbPvv7ADP8ltfYh9j30O+Tk0h
0U0JCe3n1QiTtIhL0rH+1lP/PhdUh2DMthKZf9qPFXeAzLZ2Oe/aPWc1TDM8fEQ+
fdl9JGTIquX44vciWc9w34k8lrf9STiAyzZlRQ98QXEV2LQmo3ZnqAs9IdOtfXnQ
w9Glb4DayaSkXZdzQykb3Q2xfitsshtmnCZD8P7+9HpX5niiHETiIn1IXUXi40pW
8N4DiwG8Uq3qEYXLa/O0U3nwKXuGltvfCs5YBW0gM8n7socHmlLovxoSYkVpx+I5
oKL2zR0ENcRrkT2L+GShYy2yOYVsb9BQD+RpRz0pagUfI7p/kZTV9AKsc11gs/Nm
/dp1jj/UVZq4Vs1WeWgak4yRNmL+Qd4Xyq+9RCulBy5+zybns79zzJfPs0mPTYQV
WWvj3juCk5eFZp2NU6PayqxHus1kwJISHhS279bS14V7k9qd68FHNABmkXJJQUSK
cp1eUeBUroYQk99h22uKLRSJigLcxTxAL0e68rhOO5uppaMVtxhe2QprCx/CA2je
Qle3d1S3q2N/DthojB4t6Bk5UDhISm5xrO0rPpffXbl550ef+ZJg/vCkauN9wwTW
D5aBroXpUY7TJjp3f4MCWUqNnNF4L8+mZCYUko0EM6qX3cc+xTKkbngLfDl05S9w
UQcSQt2bTCk9yfTzqPfb5ZMZBUn51gCeRYAXV41BOF6tFoqINanc5j3dfz9d8s4K
7QHxVXpfqS7owWYskvbho/+jtoSwdB0FDijNCPXhuu7my/HsveDPxPec/G1IHGzH
Glk4YhICtoOBaaDcUUhScFMjNhtGSFK8+VV+QLgF9wtPk1oPLgDg82WY+4t/XR4l
5vq5U9QWzOc2mVZb4dTMK37BWsvkukA4GWQg5cXKZ8d0UPCw5x6x3QnuLgtx0G7g
3Ay9oLGhV9cP71akcq9KJnJhXQ58riP/LxnZpop47AMIMwnjho9hf+O5tJxixYnu
fCpT3EzE8pxFRYe0abLyqfrdmsTX6iny0ot/Tgml4rmjxoBJOVbNzpRNaROk0LQk
bj/nPEZXf19zpE41oPRCzNDopJqfmyrOg9xsIZL41qvsmNgnSMMZWPl9zBgQaorA
43jxAiYrNgtoOzVtfVkjXkQWNqPx6EziDJkGOY5OumXri13DxcRtIoTNZ2uqLJ5b
IVtR7lwEU/EiVq7fBRSvFiMId9Fhsfr9kig8pvLYjlFHKkadY+nz8IIGyAJs7hjx
wJMbPx2yXAbgc7gdjSuCdtI7eRvlOftUHMmfvRRfOT8Klyqx1O0HhegP7JbfLWBa
jRZu2Bm2Te5jdo2e3Tkl6WR38p+JvyHYEl3cb0C9WSkdOfemVVzVJy1nl/V+JvAW
WxyQ417lTsdb496wzcNAgaDhOQTRH5hYREtubOY+SNFAPNGLfckTvyeL68I5jeeL
XHabevlZQVjna+iFRet0d1yXyotVLlgfuqlJW2tVqjiUyfkfIqWciLxeQsFbGO7B
j5lS0h1HGB/91+rfYV5FI+ykvAgFKndYqS50LY0EdHZegSjYb5Nco+j0kVkYqe2b
TfI9272DCb8mR1PaB///ypWrgncOPmRtd02iByke7wlVDYZ93BV7/+AS4pHfv+CO
dTPXwwr/ulNKHlrc6uuo7G0/cyQoK93oTDFB+xIg4jc/yBFCfw6X4XOLzrTqCmsp
Ryxy7swi1t4wz2hG9HUfUI8gx9zQ56WSy3tx5twLeHQBwLF7RUbgZf1A+zndZlrb
ErafrojpmxJFOr2pCURT3fg2wIdccOGQRoTjr9joG8mV3xjldirodBFfnnIpnmm/
9zorqoo5HRtzQvw2L32iVxrsDB1jeRV/10i/RkaUdAqkIMJSz0vOaReWlgQlAZVL
q0kFC/Wp+eBilx+8Xbj5RgPw1j6Ks4XIzqDCzyNhwzL0fZQzawDfoaehNDtFSWVU
cKs3hhHC/NeCGlT3qX26CyUlhWZoh3xv6EdEx0B9WkxgCnjOfPHRV+qSknXcY7+n
yVLttjf3/KX7pf5HzgMN4D04iY7QLUWJS+p3XB6ixooc4fj3Ue3arLDGucAFvPAB
zLP1CKHNCUSbIqV8fvveelmsN95DsS0n6Dww54krM/G8PUzfeto593TaqQEyU2rb
BFPTYnBWVW0dIp4oWYNhww4ey5ybHkKO9v9BHvsLCJxeVdcFo0YTjLeeXq173lcN
MlUGe9XumllfWFEwLANyFKiUu13ZsQ+iQDM9Z3Lxbbq9BjVgWuKWE4jRFtXx5j50
PwOgb682WtZ2lxpwreLqlZr7Tiqr+1w1tvnGpgUrzdWtcs4Ko+ymWS2hjnsem0Et
gzlacZSGyPZVMHJzW4yBYvPHP1KyYr5M+QXb3wLfg+Nu71BEBgsQXNkPvGHUylWc
HqVlq4Cxro+4vevrGbIkrTFWFqaKXEJjUiCRp2j8OtqHqfqdzG+9cxIgm7FchoDr
Je4xmQhJ8ogbWm+Oc5txPUCVzhVVhu7MHSmr5Al2rkQBfC7h6Ybh1kUy3CKU39IP
tBNEDuVhLL6WgT1q8/3DgdTLnEmAAdu5yRRyULaBpa4okPAeOZpjg3sX9RlpzFWS
Ui3WkRXpx4XiHordJj72fPxWjN+TnLn9J1f2nAKyJKFeJh4o4Lwt3QiqR/ruWR8p
xh280kbnXGIKcZIl1VVdGWuqxD99iKC6r9u4+j8GjoDHnk2Su/Q0b5GKpLcRnclL
QFs+coGbW5shxS8T5csKNHMkoEfRaUG/DHA9Njc2r4DS2PUwZa33fiVxd6LjjkZE
+ph1FdfRonqFwZXmdJEHgVb7YH1Z1xWkBNriCRujusW8ewE0Kk2kLLEZtYs/C5es
fCuDoT8I1WItB9GgDecGmlkfD80fHQNZieECpoaXIVO1gelg79ouIhHar5ewSKre
NMjJuAiSUhyb058GKg2bC/7bKq3bY+jTd8hkr2uk+wzxiQNeC4pwOk0EQ8/aMSrS
zcMBzoxUxResGZA3eMgBAUTq0sX+pOLNLBUsTfg+qd08QmDE5VfAjmL5uzjh8yZ6
n8Nw/RW2t0fmx1pctSjK2OO2h4ayNYttWmtgLkaWww0iaAtibikbmfjDQz4D5XCU
KDafpO+iKm6WyUGF9nkrh6T2sJPwLd+nTIdY18d80Zn7m7L1hRt8uuqguW7zDrnK
yjumDmTl5Y3+/cXTHkvd4h3j+ACDxrcUTl3nJkkwPdTYUJk3kLV9sKqYbthxyozB
CtrUW3gNZR00DHsEZQknUaqgKxmXwLOjqchWLg25K+6ZihSNCKcLkopze9ywJ3uo
eGwr/7lNuYvrNzl8VkBBWgxnWnKunCTIUo06w0yIEelK7FOSrEN6O4IsRt16kofY
A9Px5owyhHQEnrY9y6q1X9stIECNgG4og1YTylauAHiCYgowT0S0Iy4Klz48h2Wg
af+U90ydIaZPZehLG0EFJ6yq+R8A5LsRIzWw/v1O0dBs8V+S5PwzPoh5pn1py8TC
BZ1sWDn1XXL1T7ZEii45PB8i+JI2MGulQkhVwwA7SK6HFRyh2AaAKgoE0tLwtZSc
BP3RAgOwfezv6UpgX8nczwFNWHMzCCM9Yfd2dHeqTE3WUbRJuxeSfVGX22yWAoyN
AinkMzZTp57YXHgfNUCNBh81OBd6pLmskAX42RaOWGxZPNHDpcaGjZpo8BXh+1H1
matpXguZk72KOsH6Qh6Ir3nKXKWF9uJ0pPlPjO34luS1id+rRagveDQvlPaKDXlY
VOxB99DAs5bb5KR5qoRtfI42FyMR48o727NOe/5Cc+6S0/7ou01OijdFaxSr43Q4
UsbHzGLae1Qc9+SE+gh9nvAo+9wUeK2h2pp3ibRlEP6awTw8ZjFyFdHXMvkeHM3n
8APJZU0TI67RwVB/CDFu+lju3o+Lj9JPPOnt86PWNEc7HcT+9kvcAFt4HnWInTHc
NFxfu1GBYEXEqdTrhENtgxd5WMTtgX3CjSI77GIB5aW2qSIbjzyA4a4V3NeaByOK
qI6GbIy1ziesmTeJX+CK1d5/R/um1xDH5rlogK3ZeuM6lj9jQzIe2nErRDq7V/vP
iDcxp+2+aycaRNTBaCSCXoZbD/ItjWkvm0snz9oEQwHZSKdd4frqI8ep4M4AU+pI
agrOhl16tgEDB4OOyRCj8sAj3odGL4SVm/hG3fqVh8DVWlWaJQecqj7G1qc+v7T5
zAG2NhssxGQHDQvcuIv2OwtYo4cV32qWTJwMMqIYmNjfadA8rejT5VOiwEXn2PoR
fd9QcQlbqXcy5+LgMIlF5zUQy+Aa9GXTlCHDpWkmu8SgYcgrpO3pVC6bkB/kjSwV
78qvEI/jbGEvufe9uZteu7gxMZIBSNMyHp3A2GvA84HhMC1whJQKh+EIX3SFLOmc
IcTy0etcM6WAG3/p9Jkn29I8VPj57AZJpx70z8QMOnl+yD3znIvqk6CAmVFpPEud
9ZZ7z2qqUTzbZqN1z0MdHlPFO7SRbPoDJO6QtaZFUSmlAWyCmdSRrh0Wod/IZt0E
EKD6w57Ok4MgmHVwIiq4bA/BytFevA/ROfQam9ERVetnqZGTYx3oKic8d2cgugQm
YTuZ9j7GGFQ8TBLurL8rA2bmEBfJ2kb8Bj+4/NAP9DvYup71yA3PYeYwCZHA1fGq
65ThWBBv7cIa2KlnbHJzMaZLb51fPTztr/hBf6MqEOelarz2hlGJPHRgdBKsi7jG
0m7nRYqkUM2P+mb3OyMzwuTdTS4SW2Jl3rfMmyvUEFAe2WRavnKhN2DIDF92jBEx
+d9BOxjrpUyOgsle/nNt1dqvgql2hZWreTIzFIfY9f/8ZQ14RV75iLDptwlUtl9q
xQ99ZI/MGEcw1x5CiPWoxrY2pS4vDcG0BlLCxMDMYi6efjDrJV8Xua8ZPUHepCos
URWnv2hTz8D5OUPwoKfzmr6rxxbcUi7spuEzY+a04xJEy3zCg1cGwfuU8Xo7Fwzb
4/NIJWtzhxSAa2IOcPvRzTfFCmpwhoIVStp50mHuM8L95UhHzl7NYzvSwLWVOHV1
CAJRXWkOVGBSqwuQsfmMuxUd+5tfGACOBbYtdDWFLQd7b3CwPWN5CyIFTWAZ6PYc
RDCyeab2QE0LnfrokIyexIEUW85OkhcwiLddCGGIIsLSCJRVCoQLu3h5bez1cAXE
CeFOsCcI/63Wb+gh9tESo2RpDFVnF4RuWu/hnfNWQt6aI21xXQmtc41Q4wH3D+A3
F9xQsDSO881nEQ5kucOKZiDSEmGLXJCJv76L2S2fnIHpOmgMPpOZIVYiMFZl3zfF
orYV2Cc1RWh5kmJo9iPQtaysS/cUIwXg3Gl5frgJmdEqka6n0fKfmc7czTmwiIkp
pa441uwXAard//tcdvHkHr+6e4BiSDmsuCvvHdoMUYemftGzgl/3kbSK6wWjZzZX
+3JIVD7Fp0TfMgs1a5inhD1PloOOT6APuRooS2BxjcPAxe2TAF11cR+BR04gBDS1
sZQup9WiqLTtMZ5vzRmx+Y39tkajfkn1aTi0xh0e6ue8hA7BSf4mY/L3Q2Uagfh3
0VNqmhN5gzYoZFptsnuxpLNJ8WtYLceAbPyEhmwiLRDj5kbiikGEOmXFDVluaYig
448b6mgV1szSv6yqHAsJWTOzAITUPpYLGl3HuBERwOTDic0laqDSUgDY4XBJokUR
SS6hQuCWEtqx8msNALzSgY2JizgrJa1Sm7U8cTb7bCkRty4lpgUiWZzalhUi2dBT
lID7VbrXl5GtWCzr8t5bjRiwaXjQuhmthO5ZkmQsSKT7KHpnr4pSY++lPKm5ARIu
iU7rJXJUdTKaNRUi7JNPRxxWB7SLdbyVp4nS+KrkH5ow9fn7xQ0OcQp1u6CyqPjT
w0bpz4vLaGmq3GUTbl0k60ZJ12VaYfJud5uAPWSx54VbnjGw+0Zm4dibwHbihDkd
lqA/9iK7YGUWiuJTE80EbrD+lxFAnsHmIvTIt64/mDpL02zWc7D1aEvlwRHmFWqR
AYzG21w6hLExYLHdqN+rIFSMfQurzBn96qlSydR/M57yXe2/tT/kg+276p04beLH
z2bB28sfWwc82/iOWLXSDvIyhJJCyXOIzMEIevLx9NnL3vBN5kvDQpYPAoJ+b+dz
oTK9B8yGpHAbkDL5X7QH9u3WgGKsMIh+iiC0OiNVLYHLxQ/zzHqYgTu51x+PwSCR
UcBsOlFNRXbqo9eguJW1QTEbXlAmnkfc6v56XVIbkldKsl7HfIsBb3C6IOsWRuvZ
2yEbj0eWU5vesQ/jKuvCk/8keuM+YsNcReviRKnElxMBUg3kpINsXd6scNC9kWwN
wJqPkcx1FrBza1Hi98BQmkLeQla8/4fB30o4ynvIbYIuwt5YblQXgCO4YlN11b6I
H+0R2nHps/etFUlf6VJg7r14eubDcnmafuGrVxwKpu6TWHP2Q/uE8Cx0wmkoKUfO
twxErNy4pkMpnj3YaoJiFaxHkXiJHo2O/W+J0ZWdARRckIoUMorrKI/7hsII727x
Gyx2NoKI0cm6+yqWwHQDeH69PZ6KxAzN/pRomxlYvcvcCiKoNIw07vBe0N6B1km2
vume1FjB7G0fyqV80SakGCJAC/5vS86jLRuW8V9su+gmu8DqNUtoU0km5SL5C4k/
jRiF/fM4vYCN8ie9gXOJx7v5j/hPg0TCNgccp/vqs9tMnQ/IZQtVk3KMt4zgcSJk
lbbQqp/2YcUMbNI5bicgPv3T5gyXM9A0GVTt5jvPYJwEUuJafg+b38ThqhwGgVke
OF/2zElA392gYxcO63yByvg21ce8udqq2bzGy9NMKuQXxdW+0WJQvSUcQwVVZXzG
0mGc31TAXeYRYv/0hIA8fEylbZ4+Ac3AETsNcCsdBObBcQk4ts3b+FUngG8QwUX8
niAoa8x0W0vJOhwCVOgHetX4h3dVBoH1otfshy2HJ0os/Nud7a94znvEc9+Z5fkn
7aepAezF6WTS7pHvu4CaWEptereEwrNadIICuyiwK80J3/t4eVhlX8Eksq+QtCNg
veN0G4gLgz9y2g4QdAc2Fn3vJVWpidcyW56koXu+PF1Nq/qlkxy8V0kC0ClSoXjb
iRqk5/1nq201anJce2GpfAV1NBScHrOK0ZFYC52QHJ321cIDHELJAgWiRudya1fM
jNIEzRfax+OoiMBO1D18dCxDIoDi6NnIjgMvIvz2kNGNGpyOEtG5YZzpbyf3+j1y
WqpkCkS59ZX5ImgTvksCqRMC3gtwNWJzKA13f7+jFZcAUyAzeXuddll8eYmK2Pnk
C9TclWaWvCz+INjJviYAOski8JDM4Xm0KOmPUvFXoK9CAYwIuKxUK+hvHesvFJRW
H/p+v7Q4dVcXWFUvpvytmA5XAOYxkA8eZg2ya2STGibCuJQSdgzyDzndP4cSuLd+
74k6xQsSRzHdHwIyOGhw7lDQ/GydwVTW+1+IZY2YScusx3aZ+vcft/Wb4YEsdoK0
af9cHYI5M/FyKYSS9cw+vCYOd4+GlcuDapS+ahzZuCb/AY9r9GUMvz9Bu8Uiuaoc
KrhoTX8TFVAzVPPTvfGq/YFYV1xzWdGX1sZcuZLwWElnUOT0vXd2qPwchPKQn10Z
n7XuMtL7bFSzKx7O8MWOB1CA2rF2goj/EE+AcnS4WfU9eTWUWPVXd34+f5kMFWA+
tBtKVEO1En/mf6Svs9A4aG7X8fDdfA2r292POHoxTeorNhhdJ6wPkw5JCUexLqUX
8zNwF7MKjmP9b0y+Trh+W9PJwDrAeSrU7cSkfI3PpU7EWP2XlnsOAszapJTFT+pK
L6kykL2/00qR3E4o/9EghnInfeCOBdzUNvHvZ6YJYZROqqEBAuo4rsn4ozAQcd/r
gVqlPqY7jxl0weVmxr5/GXKrSDaFv8aMkTW8zIivfEHqA+FuSY7ovzxcZC/8wfgh
j7F/PeebwPbik8FjVhNa3JPIOV64pJ0fPXzXhSqITCDOLSrceuoLWnagiu2HiupJ
l75yVZs/J6cdJpeQ+E2hfYh3w/LYpQqr611JXMRRowTDUCHU2iCbRepmrxhwXYgQ
QeR4r4NSAdEA4r8n/53VgVW5POxYmIJJWDXniIRAQVQyJmi2LINLn6kuqoHDPxCy
VbFBorwC2gi9tRJE6suEd/rb/CCTSYJPApUVRvyPSU+SQ6gt8UzZ070XZ1SybesK
lH2ku/mJvRmgKq9BqKdVj2sdKtQLXsx2gg2RFNy9kqgzTf8ANZf3X8H+unFVVGPi
EaUv2LmUU2ed64E+1tvCN0otEC76kkgWK2H88OseBygiWfKXTVeW3fT3go+4LQXD
bHpObv3+o7M81AkR0K1h9qxGTwpeIi4/OWdNxiX98YqCB0WPBF29pdxFQSjHBWPh
iYBM2HFI2Awy/Q5nMWKfCZofMiZ0YF2MIzf4hHu548R2PNokega+p5h6tirzPmMt
CvcdUTrWWaHVc3tJLCyj1ex1U3wBKGvfSaTAcnGyFbvvj0wK8DjLAGdj+XoibWSD
q+bHLp+nlpBanmCRcb9PhlJqrXKH64dwPhwLNcxs07p7oOU/lUkaW7GxZYfB6y3l
Gzd3vQ5ZYKGVJ67luOqiFtZ4tr4VxouWRSiQjXAvaSI+5Jk0fBddGRLBRqKhgA5o
1SbrjnLJyRK1vz1mxefAHonGOsdYc0jdbJ7SQZZO0gkQnN736sS2cXkyOhEJGoca
JHAdihl3cfEhqfWCEN/olvyNnERstP2e5rvWYBiCmy+hT/8lzoUOn4FmH9bVBWJj
hQBqRJ/FcQSmpyEIrA8Q93OEx6gVfqbDAH/wLKZ03qzsAJV+NiJxejn/OBOFrTp8
qnhKGyWe6icOBwibkIPpxZ4bRLJRBjKQ1xMj9V/U83z0O6XsMWzhriGddF1WoIOq
34n2W3Pom1Pk1Cj1OoQU2ZmqH5vasDXBEoQzVZhNHLaQcOy0hwHsLhiNk5jwlKJ1
Or4CbKuMhzzmn+a3aq0GHS7W9lPVE07PcKRcOJD5Q93T7DkM6mL5ShhOY50qVLfG
zV4L92fbEOhGuzEN2e6WhsN7krCtqFci0NV3blANZMYgtlQbaZtZTbxbP9iIa2pr
RXZtaPG4D/9A5CTllpa+woFaUQjW22JGjTT5zI6YE69LjLCMYmF394dmJFaiDTCg
z4t2yA5DBPkTauCDZwnzqcgTWynmoPkDh1mUPju3Q+3wVlNbUdYAZhEsbIgQkzra
Xc6e81c+CI/CBf0VgfPgM/MKt73yZHLM1zv9fZee35OHbBeHq2M0JL9tQEzhd3Kj
cn+YVnI6t2NxklfQHX1g8XjdS55lar2IpVv5VgYqCJslLwPAPRf+d7l6IyIC3sdz
cegdjEdVd/P9T8VnijLMbxgebmR7e42YkjAX4wKNQydNZhyxbZa+TlHZkFzxyP4c
PbRxpCzRsS3i2O6VIxq55LlX2u7b/r7Kzj34u8vaEtJK/kZD8s/IXDPR8tzvg/1j
vrNAUhrl6dStb/jyxTlX6gGCn4tMvLTz7cgZ/xuoB/XYIMGJ7JLySX7FIyLpgWT1
xp2888K5t4yIggqm90Emj7rp2GGkWw+QdRZB8QHsDKuSbDChVPpX1hzSCLKpGVLR
rhJy6h0Sdy6Y/8J0ulY5kH6IKb8AnxnxUGddpsdhQzH+qe8wZyHZXstlHhsvPR7/
kMM5IOq1BHTtTWqYcTlJw6F/we8jjPfT89aZgc4JWJahDjh4Z7lnXKA5ij6pykRN
H5Ah/0+W5oSU/nMojHrlOlxJfwVXmt1GMsTjzntKr1O3OAI/xGO/xDS6SfZAF+YX
nSloKZ3SsuaUbZdHDRhkffLgEMDZW0e5xEGiXZiBEQfKTPaJB+czO0ds8Luw4Zud
MUvT8SSRr2FeXQpZ/QMlVje2nZOUyZrLp8HcvwpZ9UpiaREsqm46U7zv0UPSTvMd
ymGYGY7/2cDb/DeBMAh1tPuqw0E/1Hy5nMat4AlTylvFzpgLdgErboBZkNpvsr+V
RYa2YzzDZGlRUZk/UcOLf5QsV13zN1c7tqlyxVm3/m0aVVdthm/fP4Plg5Cz+lba
akjkOQ5/f+cNOe5mr/JHn9poHwLZGqiZwVdvA3WP5po1JzsGFKNQLCGGVCaIyboX
BfnY7ZUvuK/SdJ6YpJwgF+OSHkRcBuJSzyZ9EJTKVPNIqxTCc7iegZS1X/IelLzW
dD3Gw8IFmA0vZYTdaT+XLz5p7L0h5XTMRUUecfrmqndaoHcuCIdWJ7KtN0KhrH+5
OPcPxLKE7ByzTKOVMswtQRkeg21IJPUMy/GsiCkT1fx/Gt7iblxUsZJLMCh+jhHT
caTctD2RxjzJntgq/5UB3Cz1RL6bWCLh7axvxhDLyL/jFuZRV43YhSwLtJ7/Dazh
eXb1SJfVoI3EgjikMhDRzaPSvYRr/pFNHxhNP5eccsIUd7Zh5TRY5C1SkhSEH32r
n8M8F6zva5BcRh9qPSafLBYK/ESp/j+XzZHCeucPLJ4N6fJg48tXyVrSUYUYYmoP
cOiHfV6pj4X+fr0MK9JczxfL3tLdCiY8tgxrREOd183DzVR1M9ReTafYN7WSFP6N
Y7416RDzb8WPzEFZr5EAa/H7qc5+UGkp9KDLDVsY98P5wz2ZTslReHEvo8YgxVat
+SgZwd5H5l+gmpnaYcsNAKMZqdXmbiC643wG3CxwMae92GV68MNnHSoHsU91V9Tn
WQ0Vm9f0zjlRUeNQcognQj0AkBAHae+HwZUoSiqoXJd4r4fPc+8zqHZrz2MWBDmh
3T8NwQVn3utGj3vvWGp2alebQI3wLh79yWE4b9STFqjUuys0RK7YP+H1WokACg64
wJf/sJhW+Kl3xBj9btY8H8YT4z5qzZE55xj1QUDFMhBfWpEnXaBChyhMhLaWDF/H
8bnDR+JlQckepOtLePm3C3dDJ+LWJJOsmCGB3gmVdytzl0LbUIbRvtwIF+p43Gpy
5ca3gRGlIrdH1S0iM4vA5cJS3FeHKlKRlIgF3N02GjBnFNEmZOjoYDrhrnhursd4
WBJqqiYHrfIes7kSeGmWr5+Gl1hs7P5L/h4p1JUtbAlxKG5ZUdTselZ4iHNjB09E
4TRdrIdh5EB8w/lU/vq5u0nudCo3/bTEM4pNVkx7imVPmv2IVesIybU2I1EDv4xg
yvzGk1/OZnMrriF+b7lnt5eVTwzngAw/QGbx7fSJ9VztDE+iQhwxXfazc0SKeAJ2
yQjoxjigHzj5A6MqgoQ2SbEkWoda/rBFYomWX89gctg5ydRjSQzmN2KfNmYvNxp6
ACJib9Mk988LY4BZnidY3CONq5+pfLn/0dY8ViOOADcVp3CJduzFmW6yO0UgPRCo
wIBOj122Q1ly054JQ4eGgIpRg3sH1nHk4Jajs5RavMf8llXqESjP1DhsD7bYZiuX
BNsv9hCq2Zh0qoxRcUeZJPKmQhCyoKR3Y4hieGsIwbDp3Elo/OrfOBpL0vET6b8j
/xPHQVN7sS4+o668QFgEkEHBOgJC9QEFebcFkAB6a+HJh1OjwUzcHzXcvStx8aXb
uyG8ort51mf5djm8MUlj25Zzpz55X3L+5nVECz+ld5vOXa/o5EKBQSx5wNTubqZJ
0CZsEsjablb0HtxO0ZedL63twA+S3MDznfTEcpLzf9AivHKIQ4Ll1PQaRR/LV/pc
4ixEJgkl71mo2miJsgKKindYTVtUrNpLSe5SYvbPqUsfTEntMthls9HJnDAv8wl4
DUnDpSHGJFfXbHXlhPObxGgJt7vDDfUvG74yAHdNjxJzLyl9yL3CY76H6E3rPRvC
pCnamUXPCIOr0Q39Cr5gJgjfIo2zmoSMMuedoaVzIQKoDFM5alR1DhCMCjIXGndJ
Xcr389mX/f0BUkEg+WdkGmH6MlBNgP7AEtshDb/NjgWL//jnTOuuan/ONsdLLLLH
ehopBaDBeo3xTioYD+1OE3gsv4JmPfhAv1EOaBi3pSum51EKt9Hk276e4O9qDiug
44ixsMqc8abO8kX5+h84TFKBeqM7Zhef43MwhtRNee8yot7rS56cDAP/cvqVxFfh
SyjJsy5lL9BilqhHa7yHduWoUI2eY4vYlwkR3y8crL2PRe8gsLl/PpyMldnzhwzY
k+ze+LQfFeLhBjzpx045lzMC+XB0e2deZbLS+NMGiq7SeraEeGUBUNpn9osguaHb
16o97UKAQirpM0vkPq0ZEc8JJfhBWQYvSLNvx3yrT0S+A4YGhz/JoQcBkIlDQdq3
Ge8/L5yzQvsFH28+v2SU7UKoZKcN9VbckA4C/laAcTOmqeVHPJZ3xmFtorJIyO5W
z34wE6A0wcIsP72vJt+OOlR/A0mKDLBSBkSP5QRIrZoSjtqCBHElf82KpZOcxnY3
xWSmXoKKrrDH1Dr5vpkN1DLfKb34fg9agYZ91GhFWBTVmlUnYDxFCZI25wsY9/CX
hz23LhS2hvHHXxAq5Rb8dxuE8jibUsVm+OZ7snRmv6HOI11E2ODSEId/vziu1zR+
1DypJFhIhXx8nFIJSlPOJRVsaOE30my3a9O4j7X7MtiyCrnShu9+VDBD1MKk5HSY
xr4pELrpYxMUQWIPhw9KZYHJG0ZmBnH3u7JWt8MTy5hDfTbUf+ZVE+lCsFdZ0j5E
/32s57Gq3iPzMRKNpcmQS38pnTFF46ksEJMqohzaQWP5Yn7Ufu+ORSWilrRA0aUc
D5XnioskZvtY32s/WicEeEsjKNgXcfMeGQkl1b6UkLCmUtrwZ15NulUsw+uuh01C
4067YQzU94A6oO7yC+w520E9rQcScars9zi/OmUpJCJOwie/Tm0uA6mFsT5PsuBS
cfy/HPxaE15zIt+OVsCUDxwn01uRshso6Hz8Enw7Jlv+pVPdE0XhffbZolf54TcI
6DN1fGFSavCwO2PARaeMjNWabPIjq32Wn7z3Y78RWwaphW4MlZWIiAFhcv3Az6ro
Hgf39PBrkF6d2c11/y7wP/yOvpgNXXTbuF1Hm3TplzUHSXw8JMAGG2vvwCNHe/Kx
+yYcrf51Zt20zvZVl2mGBZwUJaY4xHSow/co0pkTdLKVnJUVeGhK7HEC4VKQBWvi
L+jclQFKgsPT2P1959EjWXcYXJJcBfe0ZospvllS8qObQRwAzdOomsfipAEhqYzU
Sn9B5uvrjKhTEGcCs0EQasyJ3mNJE3pxEAfrCEkeINdCYtP3fiu/Jy5s8XRxQpXV
yFkDPerZ2IYv2l8kvG6Qss+S7yafah8dlESdxYsWxf7hNx9nLS1DO2sN4av0JzGO
AqcHz04kd9fIeM8QgAvYvHQxvFUWXAjpxCrLk7zJlWnhkFyvjA/eTrLeHKfYKH54
iR81DFjJCLIpkvR5FtuCt63sxaDteGjEZfudBlQu/99LYGaE7olYTMTtHYGfgzDI
vzTNgblpJYxQjfQ7HzXKD8KahxkOW4505aXrLvcGBXfdBmeQtr8bB+8kwxz6H91/
yElTV+3O4ldpc0MV7gEQTgCjB7k3pNo/JXymS8jGNFvlR31xnbGubSc9/uAIQFFR
KZx4/vAstoUm95S9gjKgVmvryLIvV/L0NFkEaAwICnWZivYtOHGI+zlD5qpShTEa
KinWymLA0lN+T2NpDd1r+ZHenLupAiP+NvxaX9JuMD7kQ6IhNqYoQn4+WWzNQisd
fZEy1bPY8jBYLMAm5gFFMEQ3bvGJMy5VCQR/TO3EG7bMWfB3RdyQR1uB04RYWTTU
ElifbeMRFloC1+UopcaJt/E9Nq1sPqTxMHJHh20Jj6LRkbc6mOEs684wFfqjeF6F
avc1Wux4oYXliQQYJtAiF44Ar3rEG70quKyeib7VItN130w0GAqUAK48KVdxBYtt
IID7BMLrPnM1lR8vNKnOJolHD2cs3Yl8Qdk7tW7Nyipj2iVQjnuH7MZ/auXquOE7
OIOq8amEbFTsyFfblcwVNxgiAKmEVdhh3k4aNRlG4W1nIFmOSXDfcUHEQLtLlJGi
e5Erw6uAle829Zc47uzEpCATutCCGmNrvqF6AKrl4JZUz3yoNg15RB88UsJVY8lH
6VVkV5HqVfP+8L+uZ3D1/Iw/RhseDumow1jJo5Oas5k7jEcvZhV1ZFPU7u2y8Aou
ocZT6kDRhNdKHMqISctLjxO+9gjUEpeAcDnm7HBxuzuln8FlD4LJjFfEVnRuD+DE
4JKAqqNsEp86qEUNwY1lUyohFJaHtxcjrBrXeZH6NOooxY8B0dX0cUoYyrKCvZT4
8ml5wWhSJMCEpT7AOk326c2d9VVQu1+APq+gaLUaFIp4eMfTX2PxuLdmYnQGT+qB
Gsi80iA78tgrALGDjGi+Cf05Y5LCeMD5XHxBEpmfPVlPfE43qI0dMge65gfJHnuv
2aQdALxmFeKYmw83XR7qFKeXmAsPIkuBHCG+SWVWPkii7ZTGaSPvakFmegsXUuRI
drq0k/tJPyKwKzfy27O8ivksa598Q2HYn2m6YkDOXBP5BZGenYpw1GkhNoKwl1eL
yUIjaj547fLtrNM3LQub5Awn2et5Yz9SLslDbCHvqTpIrMlYVUYyK+tmOzGDqqHX
doPFhAuF5t1lMaHpQsbd2puBcNQAy/eedOlrXtQ+p/7o0mKcZaCOsK7uWcPvghuQ
3UmQjFI2i57WMRrn0XIVnA9J9D7nXeo6AZ9sBrcvrNqhnCJ8SmB/dvNdmIL51jKg
GB32tDvw0xePsnEWfzZ26JcrR7siIBLrHC+ap6p18Zi48Qubsxk/umm3zj1PRf/2
nKTzj5cZKdqmljn5KyuxsescF3DgfO679pjQWNSbisqNICXcCMVRs3bspp+3MoIb
A6ZuYoz445P71MHdLi+GLQ8qBXnBQ/xxMU0qEDM1RcWYb3ToXQwcbfJCGar3Fh6T
Somwco6DuOyHLoyzHRcfPdrUXXldopQ01E1sCfe7AFvZLOYErQdQfInbPVk0kxZ9
upGOY/fxAkbvtypTOB9/GhlRMk9zovcibN6laFPHg7dH3ga8RIOJjQAkK9/AHxxT
KJZeRHTbvsIVatQ44oOHzoYh/J9IIXLS2XoAKtCCg3r8RSIEys57Hu+jU54UYBw1
sjb4tYWpO5NfWqvUEHjo+86lCme9hKr94BhvU0bhB+oI99dbtH/9W3ZTaiw5Ih6k
ch4ojb+EjEwTT9Q1Uh1RyTi6+8ybHETGkbGYgHvdQDiHzSdFUsVZ7XWNZ51HH/8x
tUvgBEJZ2vBgnjKsiqiO77lR+nRHecCIk1qBg2ytG5tHQ48fUT8tZhlUu3YvcCZ0
B0mvhCtXdYAjBk2NQ3y6P0XQioqZUD2S+845GFMaLrYt0Ug8VtL1uulmqBFhUlv3
vD49Sr3jw83HSL2UfEKDXYiCz8f7Cw+dghziEbTgkW2vtWXl+IPEGf97iJXsOL5w
FtM8Bz3xCg2EALIxLvCnnu3vMwAGv9+t3M1t2GqLg0uC3y7GE9GwXcfPenM8loYd
VqyZW3hSrjDcO6EhtiwGm8yYVYgIQvwAuKeMI9zOmfeDQWh1VmXHPJMAMboxh11e
esbWUgnDShDOCZRFR0pG5K6oGO/LJ7cb3ZAgIbI7NARw7XFN6WB1RZpDrxIVRTp0
40Wd3xcXo/Ln0k6G9xv/6o5qL1Qq5Hregisdj8JG5T4yt+32IDQ03I3kVNz0ElQ/
0qtniowSFaO8+rT6Ewkcbh/HY63G/fbr1r0VnJJ0UgYKJ7NRhlJUkS5l4cbWpRPw
gjYgH7JpYUsB1yLhtDQGCzdEn2lNMuu8Awaq8tAV73miCdqZOYVIMwPO0ts5/1ka
aPF2NcDocCaWMkX4IoNLp6vgV/+YC+xsv+1R680CW/SdcDl5Ji98E2s2AhNRNs6S
UP02bHr3rAjkKUjy5qbRF8hy1S1pS0ggiZRuxfeP5fUzqLcztIuNxHq1zPXHE9pb
VvRYLq3TpzNI66NU4zqUepkSsKqidQ4vX2nzETJPGXQRcrHr1koOIPdq1EPRX4kk
El2TYH9SJ6O4H6exKu8rT27rI7jsv6Z2I2Ndv/jBq0WZuumgQW4JKgzQjmtP+GNM
dmZ+1ijsC2aWCXcYXKyaph9HlNI8+7eXIMdASE4hoGDeIp6ANJcvUvLMcAIeIlYD
8MDXpFrDj6/SqzUDdaBz6hybDA4dcnxyHNaXRYEEXz3s0bi0vAGi+hGxDmlIQnJh
aE3iV7yHYID1AXvbPpfL1/Eg2KVZs0ZV4JB9OZJRD56PtmDI52cBmqyfrZ2Dx632
KKV6sOl0FfpgefpCzLEHiNQaQwmgqGK2O2s0iW8bL2sAyP2Xu/ZJynUBAPbxMoSN
afQUhuzzjlCEJbXmETl1HQaoYYhO4cU7u8pzo0KUs4aabJSbYrhKthwXuR2iXHlo
tjKcobxJGjHVIUWQsEW3jbqYB1lS+rgXKgJ7iL7knKm9/2YnNCYkLmJ3wqyjyX6j
SBA+xrff3uObki/QBd9+JXl6vJZltH7aykBxskMMswSn5YmUv4Lr5Y2DQObmoh9v
txK4SFQzm3aa1bBzKus8v8gOVNmI+nDkzvQbgy7ifNtMb8mx7kXIU2xO/yZyzP3N
xCmEq3ZpOKJCSvFFgEllnlzL90EssEq5VdTrW0YFpdhnXuQUt+SGcEug011cI1SG
hdLf3A+saV1ad9rHdGrB8QZvc/1P78DCzb5JYwz+2YnMddrrIjjpYbqt8qMdkuzG
DID98EkiZUMvqCyekQpMaCXFuI9e3HO/TrLAqsboVS8zdi6NpXItTTlRRwdiboCY
ZsAYkPcgWwZXiBaHiH3D4nO5vPXl+luDYOPtudwHync/ihVo3ty843AuYa0heSkk
HNUkWI+KMonl7Git9ErkTH9al6glT8wvG+kHhpWr7gAaJaLNF6O2AehuVHD4+hfI
Pi3eQPrisLspLKjPd7k88s55apvpiF7ANGwpSbxtYFkMk3Qc6dl1vWW6eJ0YL5E3
ZS0yU/5UoluWVWmIjLmfNsdKW3PRk5GvhljJ9XQ0gv7rzoxwdGU7w3xPn+iEPVZG
vc33kI/iAk+nSMv72ifHmSTx3yNaYe6MRRd97UslA7S1WgmLMZN/CO0Iu0sw+vZl
jTLRyAm6IWpq7wqctONaTK4nayHEPX/J18F4UEQy+TD981ipeSp7qPEUErBoZILK
qLBiRnHhNjy3bvu6AOf49rFWupJ7LJsRexGtCFgD5GVpxVVWlkYqzBALMuEoasD1
br18HR9SjopBvOwSdBlA/FfG1/fnpb3IwbNPBp7RKWx1H0JWaPAb+0P/yNT733tC
ArLbT0QSsiaoJroiqM6SBJAlZBeK4FhS16lUPY/hDaEdMVXA3oGeKipEuukYUONa
3tpEfmaT45vHH1mtS7MKDkQGZEX7g+b31uwcJFf/o8hfTCI6SmKxEV8/n3sJHhbU
kjGqRZVP/4in7nYCOgr6QnV6NoX2QXOVgdkLmD3H7CmSwyUDMR0mgrEobzmbfuYq
VyqIi+TMthUNtBXjSPowCzQoOb67VxzQsHmpFsjt3X5EusPlZEfSJxHr4FG3Vxfc
t0HFgBhueu21wucog7P203fZIZ/xgbdOEjdV1K273wQS7PtTfhP6icL4WL8M8Cp+
V685NGEaiWOwhCMZ5Qute8dDchDsyz1i69WU6iNeiLq1z803i4lDYSdsgAbuwLQv
MhvWAs4riC7jvLfrBE4q8xRXfJjhNjcovqbHL0Z612OSmB2W5j1rOo15AwRAjFRb
+T1Pdqf9367d3tRZbEfGGa3OZ14/2lkLOP4OVsCc4/YuFsnnKbqtAY7wggCkRvV0
XxeKFMqy32X8nqjitCyWH3f6CeBUOXS8v7YhcQ6oedqK7b5Nl+/7e9gXyTdAFqwU
+rouCIF7khD89ueOD2LnYe9bfTK9N6J9iyZdg8lfetw92aRXq6MaG2Z3eo7Oqzn6
Ha6mfh71VVCu7/FMgreTly+FzlYHWkj/eIAKinPM+Xxes/G2X/Cn26D9mRLukEso
Y9VrJ1p7V2Hc30YQDqRXIt1ai/AbThXlBfw9Ul71+BshYgF8Z0R8KeDgZbuHA7X0
IyM4pRTT2VlBWn9w8iiMU2b1+k+t4xsSKAF3vtZD1FsUuaR5+LqTR9VpAyYNQ6Ek
YxBf2d6rKP3kNGVMY+jnkebq+5t9VIdyVNUrICXYPl9PO5pOIAu49VyXA2VtI+Le
ZRxnbhmdshVLE5akaawh5q7xM44GxYBD2XL+lZqMw3Ok6qbF77Hpzf1w6zrqjvJ5
2GH4iogVF6Zk858v4snQJUwNJAeRv275EVJEpuFFgdsKBgKuh6jEhdBCHAIUs28I
+VpxMmkeCmPkxknX6+ypoBBAroTn2ymfJuiA4ZJPakTjq32Xdy7HIakeddmVsP6k
MITSbYSyzMW4/XtL944BLeAUNUhqgaMESz0zPfYtQ4KEl/ZHw48aeaWuZ1NbidhB
PCDjnjQ2HGdGKP5DaOndoUEPNMW12jc4uetTKofyTkCkG3AKfqs4FCbcJDaS8D6S
/b+f5VU+tqwlkrSrrFc9tv1chN8s9fMmTQhcChvZhfmZNvTmCJHQSdhIqK02WZhc
+Lu8yitIwH3qW6JhXDa917DZTyEKoeL7AkQK/FK25YHYoWwol61/C0hObXdvPi7M
CDfyEJh7K/J6P1ycLigl+R8Va0JxHdUwQXEfmqnbxaVvcUpjUVAZKIGhmbxI1elk
lhttePd1AOY1QYkruf9pUwfxOCEgqFS8sTDKprOdbNWbue49uqWJW3LCV3XlrqRo
ORhPFeTAX3ZkZ81AG9l5PQEwOgXaAtCYpmS87HCEC4iQZn6Orn9FCXEnKzsxL/Ac
7NhmOpMMsnO4hNdDvXTQkdIZGKNH5F5L/Qeu4iWcLrl1y9350Jj2Jy3EVC0xeK7A
M00tMYiDVvN/a33mZ3gHcU/Kh+614Fbw5jke0pa5KH9GIG/uIVLq3tUy7skZhBhs
j5IZKQ1JictnDLpiwcGVTPOj3mduWRmf3WG1r+K9fa+ApWMz4niSqVr7/xuM+G8W
VD6PEnqFfXBrbu2bXPgRDB4D9ldcohQPuX6/Z1gv29t616wi7GncBxWI4ecQs72N
mcvBG3zXRrjMqRFD/l6LJiACsm9TwlXOXPzlTYPsD7Nvl1m/qKe4K0KhLYmkpyUZ
cx205nzDR6dbaectw394hgbbOGtpEDw0Bg9YEuZe954kHbJHF6ZICSZePZQMcrAj
P3wnxRRqx09rr66iwSReUCkdE+2yBUW5vt3/GYjXxemPA+n720XSeypQJuVt8PBy
dbtLFXwSDRwag2TwqOLLhDO9+ASD5K0RcXAMKipDoDhGZzDRFRytbg6nKE58a+Lo
j91Z2jGaEk8gXqp9C28RCWdlgesnL4lrPE6SiRItdZzaFxoki1dZxBgNGrcqW0wh
bdLxj0RCISo+curWSuGko2O3cTvJwbGuClck2rvTsf1opW7W+Cm9mKyNXM0HND26
qwB2mhr75O9sICdOsCGh7OLdX6goeScVezvLJ/u5edutYKlxv37SZZSmrJ6duaJt
aJ8tR9ruJLZUxs5QQirurjBaNTZFg3FTHl19Oh/hikxeT+uQEEXc8QSpeMhfvr8H
TLYuUaYDK4X13E55eenB2XC3eottMExCjPqIISAl6Yn5Ll0L4K36OXi57xXnfuYn
x6LLKw/X1LRQ2s7analPJiue4UZibbRHqW3ufFlcSnBJ29XoHDjRhWiQWYG4qf+J
Fsy5d1+Dh65MjH0jbLwJJw85bW6AvS0yYAJ8OmmtCC74MCeV3Wsnf8wyxAJlg8+f
ILm2DBzII4ka/8Q7Xqb9Sr7pyhPD+/R7Z/iCiOcK+kAErTxKat6PREd7drHYxXez
X0U/IyXMZjNN01hZCohJO90Saixtt7gvp6pY6ffOXHbTHSqeP8a2SCFDt9+S2njJ
fer9kPd1AOqp2yZzOvp/DuF5/fYDr/8KbfYmjZoxP5LncTsQ+sjjIyxPXPjrUL5f
yQ00OJcfmFEhVCk/oyY4XuLGOO34/Psg7PBEnkYAbgQEfb61s2XrZevqc/rJP3na
1GLd24EfQ+p7C1QAfqupDjqM5tX+gZAnqVU1Y2UoCUE9pOUGxyhhcpX8OfxpIJHj
VT2U4BAdJkkHF1+FKCs1fd5izQ87W1SE98u5SAOEvjvdgD4LZu6x0TOEYOu4oObh
JZd+cvEbsfhq95G9jxC6ajKvC2/CEO9nxrdfBl+GCJEls3OhRool8EtLVg7BJDPN
Omas8EH+Oczz1VlczLzKYPbAO/iZOY+575xc6lOJRPtA5e4i15VikDrOJbI6Vyng
Hrt9AW8Dpk7u+SKEyWrqZV05gHKbdUlkCsH0GLEdBGLnRTjAYhDyD7+sz5LhM2oB
0U8n4ZN+PFkSxOrpEWh9rY+dGW4gG+fH72xqD3hC+jMDhkRULULfZTPJMwThTCzm
wk/ISpJIHrSFWUAmzfJ0AExBJyDziah0UR4e1siPVnHA3w5XrDinPlR6dPhOrFYT
pK2d8XWx+/k3XO+/2xuz4f8EYheZayq6Z86eTM/IlizvO/eC/XKGimYp+5UyZpHh
R+fkDR0rfOYuzuri1r6HERCf0cUlGrs1kqauZo1K4hqLietCU21rUs1me2HerDkw
/Q19hiKXPGt7s0uIIrgHAnL6owjPnKLL947jGOuGT3iCwsng2dqiQUvkLw9767Od
DYG1iINvNPscvasDfZxKTHu6LUCpeaAfI39fHlYAzB2Ff1QHgz/9t9IxEXdqr92V
llkT3NnXXM77UYZE5IKdvXVcTOGDLWbU3ZQX4aXoYmoHw+9thcyWA3uEqHTKvV3i
07DQb5w15AIR1mGJ3+kAuEXKgwozgcl+HKFtZ8YXleK5jmQ8OTTVLDLlWaj8399b
PAxSeQ7ipeL2pNXnv8iBYDvGs8d3uiIbJAe2PINhXBEY74t4nVqrxembq37KwwlZ
KkabPfYKwFHzo4DPB7Hi8wTjTNOvsYE0hyMPWNJgS7FJyHq8fXPxlRwYzlzSVDyv
zdNBArhcuehWVURBHMc52UtLFRETFF9HXztjmhFkhXlr9LFqaqr1Fa5hm2ZRwEoy
GOqUiuvg828Zk0Qx9wbMS6RtxOjuyT0wPd9ZAvZfWiyND50wGwPaLlnnOiNm/Hmn
pw65xk+1G7YGIXl8mdJXXnpKJLHd46SvuRKie1x9oriq38oBGO1r2Xxeg8uD2f14
xLLPm5g7avDZ3PKohxmi6fSSZJSWemQV5elqVtV+xPYY84AxlZ2iqHcD84IBOIeY
z6SjDc93wI+mM7e/fWZP0pHc3TseEKqDyzYdYfsWL3+R/5jniJ/cX83ttQf4PfwZ
Bkqk/w6/J8tsaAbycEsggmpRTRF0eaD31b/QlDupgGzzzKb5tU3yqTgwtZM5dReV
vTXylLmCdBvvG5zjHp6PyHkD4wgFKRaxL6RRPq3SEqu9J4V0Rf87w1dcHDyJvP8H
tCX0zDn6AT1KkDK/zQkOSj9Lb85obMp9e7lsMN7hY30u+qMRziAgL4hXI+Hdg5qC
3iVdik+Wmjuz3twsEZqHbck4gWeIoS9vD8aPquviZ1fsEC1qJxYAGY/mQkVVk8Vl
/98wf4n9p+Yxmf5b9zmwWlrR3ov8QWnsyf0XljmsT4NclZy8i/5o4IL0x8xPbOUi
FEQw58gIjJa1KcTOcb0gx7HmyUmOHjT2+qJW533b/yprfLzm/Jr9ZCuT2qJagOSS
kaaCTMu+V2gvQM7rCvqMozu6Q2R2LOw7ozVHPWMqJmntmCqzb8tft4Gzzml6qP20
h2S7UTMIsJXBFmV6omYveM7ZNoDCwIxOuVzuyxNj2H5uyOFF74pdWtWpzwUGoP3C
Q/oDihDgyZVCuTvmohW04goHTkmpnWoktpl7lRCDFVNhQna/sHOb02BEVztcFj05
976fq/ZQ26OJtkJQM3IN8BSNE++rdajZppB34R1QjdqZ/HKWwVa7OgWvKo2VgoDM
EmwInXdJ8ew2Xwe+dAcX1ATp06DGNREQLKxQjdHNOc0KGRjZZ6VV2qjEXfxc8VkH
MfyJRIUfRBJ/xjtfFsTUSDEYNnlpvJyj3kaCOpngQJfrAFPJKW8ZU1OPnqx9bd8W
iuUufIKAWNOrHlhHczjVLO4e57l6+xX7mq+D1O/QO/efnkMl5COWu39lzf4PHt6V
tlcFozHn/Zhw8ETavU2uNJLIUZUamJIeBPksDmIL1iWGL9Zs7wi/p5UpAN9P76YR
D9dGV/0vwde98bR4YQccbJqJqUG0XCwta3apE24I2oYANYO1ZuV0ixgkNUObs4Ud
8FGTIgEoyDgE+g54L2TiDHv+aAB17jg+be7ld1rSl/NYJRFi16ii3twoFVWwZ5mm
lqa+He17NiZ/d5v7RIoc4wpgNnU4SKM3Qz+0JgWorBTcZGlrq3rLyTqcG4jxx2qC
oXt11ZmWRRw+2OSMuIkBzKZIhdFaR5KqPwZSOMYjusiveM7Z+VcXSzSo7XRqUL80
2svIB7J8fOeQZtD2Rx/LtxN4dgLrN3OMR7RSnz+YI3rPy27bZgeLqptehWHJXslu
YOchS8L2Y1IXmfpysMe+sh8RoPe3xbzWuXe9LusampkDwZEZvV0gI6O6YC2BzZLi
qNtoqbvJGv7dtNNEkR11LqKfcBPyIiOOOsD50FGASAQIOoVM5TGq8FbctZL+9FDb
TkE+f5R9P2N0ugLpcTXYdFC0VifvQcSo1kGJDrrvsn1cDC6casnbSwoUydjm1pRu
wiEHmmfqC94IyHC00qU0CZr3f1+Sh16d/kZz96CJ0S+OOG5Ofi/bL3uBsIrFvKZr
ltVvlwRXfOAoQXqE9Dn1ikQT11fPGFIDFuQvj+nJ+nFiY0HEDTgHq9cGoekcaE6D
P2E9SS7pLY7oc3hb72z8gfywWeVCyCzkPy47vy547BQUe3HMbUdgfI0WPte+6/6Q
7qjBMS7SPZDfz0dmHVbHZKf1/LCRDNqgWMX+e8yZZ042ixbXQ9IR8JyN8ujnARcR
xGxTpxt4nlfanR/8D36zDBKqLsWHyboG2k1De/XyKNCv2CEqgRHRmbApOUb0o386
U5BZOVlu3ofN08IMMUfPBZvstieGo5Ka9FRfL3dyaOYozINwkUythL0O2w9DZbs/
hP+aETDT+672NRllkf1mYFmrPHzXwoZ8TOGnGfqj0TLKNfzYMgRiTJP2ghGla5Ry
iS2D+0AdrkpiPzWTNVWusG4Fap6MfHtjVfBgFRuEzBmyukkcwKTdvxJyCr5znGd4
5lM/OWs34Szjs4rjs+SqWgnlddLhpgzqtu3VkL95/d5o6f8cq1GSx3YVqIL2iouA
HVwkyMRRmC1JSfF1QqrDjX4MDpq356AS+/M3Nta63TpL/6efxDglTaKlWve8bfWA
Yt1qgGvttAQJAn7SmjSJ+2QwaGsS8onkqeL9Y5qUMvfmn5ZEZ7dhULB7tIYSyOcI
3RqdSfDGQVMXuo7tEFoz4VIShOuvGJ0V+6VCAcl6mLDdSc2u0mBgJ03hp6gJOChk
Qsq/0YrBNBuL6/X8OY50TS+rd1AtVUMrMsDFm3gdIiPQA61gZw39fz+jmhxOdkif
Z3D09twuf6QHd1AYenI3VDSA19reuwz4pP19tnq0gYePIx1LEnNBbKPV15Q7pZdy
LiNXQizvsVZAW2PS6F3xNf3Ai0v0bQF+S1dReQ/5AK0C7KRjqkW1H/DqxSDATaCr
f/faJ+emcE6U3s8gDoE/Q7NByies4kiD9cx+tXCRF8kc6h4JiGE2WKM0a+4ABLP6
6c5Em9SsFbgHs6gcdEH1iM9/8C51EmTtxE6rTIt0yxdd9hqLi9VXVMPPEKoHNfn3
Clhqwxls65c9kYD5fu+lx7CN+TXoEFqRfY/c3T31VMEREOSYafAl/9FtUY0Zv+6b
+/9EVmdPN+cgHWd+yPNGwxxdSHriEZu3S0eHksJPsUWf1fdE6MENXcAoUcAecrC9
G6wXySfUkv1R2islZEYKOzqrhO/xzFKxDKSMJcfultL+TLWTKhBTXsY1LLWLJyP2
9tayicIXqUGgkU5+HTEKQRdKkFzFWvWDdglo3EQ6Icar2f4nA64fqxtQCsuHLbMp
PEdLe2lRHHmdwrN/aF0hnIsVmqESNifGnsrb46Nruj2ZQazq0C8n7IarVxhnNgDL
JFttUISI+Ot+YHixrxuDw86lCaW7luEKYeftSVvQNjc1SFdhPoTJCDTW20YlFLPN
TleTG0hiHTRLdLomcAThlb20PNAfNKTS8CgGxAXy7asa5phbeDFJfMrVuvYhMB6E
zdEScWfzqQ+wU7JFsP3IGh3z8xIrkg89zvlndC+HREyXczYJEPcMWlXqW5dPO1Zk
2w/e1bNj/V/RYc4IeJU00qQyW3g57q+23YlrTSLek8lySIRGgEfMp/oBNvoGt6R2
DKtfzR2AsfMc+xVmN0MKSMqUpMnV5iDhgS+PZTFCBd5+AKZeozIaedaw/9CdL0q0
W+4Aa0Q6UzY7GI0ag3xeQb6S4ZQYExSiW3en5IJIor4C4m7onPYgGT+tgt34H7+m
qQ/MDkhJd74H4INyTXhm5RqVIUePANYtO/rHK6X0BZtqvPN60bndUmWSbobUZfru
wFY056wwSdiaF1d1x1/zHBEp9Q1hGiu0doS4FnYQSBdJ0tRe2jNKt6WEhNCrw5Fy
AgMAMKh+xYsMkZzc1G+C8yI1jCAl+0amOLsPHTnmY0ta/CsSKcA26IStp3GBPRqq
7FInvD7c1qeT4jHx3/jnK/3P400kcxL9pIe3h9VNf9M2mpA+ZJI6KLd5alc2wQcR
ftHGnOJv2QsBymCSCEYTVYfPaBedbzd9gVeuS+L+eNrigzVpi+OVPZjczW5e1aOD
+ewyDyiplsENv6G4a1FHdDKR2Rdx+FTYEV0ELl+kIg5QgBbecm71kQE/LpV4sMon
vFbFa1vOA75aSwVjViQegBMrvZYeT73ihnRGz0CLp6f12k4BeOYU6lyOHPbdJmGS
RC/xqXXqRQoJbg14pYefboaPPf2Jp9ssY9mzr9HdZwqsIf4hG1KTRIptsqxTzITk
Q4B5RstDyER3cAL1GjjS7J+HoHdUtP+5WSfDqW9/ksUvWISqIAxntIwSF+WO2SkQ
69YVQEadmRK+aUdMVVsWTGWM5VZJo/hCVOKUkmfbFFxGjgFlxeFgJz0tAC4wFLSp
q7tyuZR4UZxt1EOEtPnxsPzbX5MYTDXPb0mKxzDz4NBhGiG5WUsGlXF54/QGeNO/
Hp5JdtL7fA9yHoG5inJmFVaAPaOo/15+pD1rIKLQABw+prRow8tLiPgRAgK61YXW
XpiD30RfFcuzgNw4L9+sKN/c7waEsQLXhvb7MWqoS/8bInF37IUcSJdKs2Psy1KA
Z6+U+PHnt2XSx0m0tU8p0+QDgXAQKJssdhejfsTFK5WKfOS4FzYTsLbbXqy3KxG8
aes9W+NnjjIROPfq2+fQRZW2BZq/dfn4Y3Cxofa4MtmYJIAh4IOGM8fUqPLKAc1a
H2wIrk+v+6cacsMearJXDyhyxaJcJ5BRn8eCo3yK6PsyA/ryFXJ1xiJEbzDHJrp/
yt6tks/4udCgKRn3PdmvPTZJfRukntkgmJB02085NeoGonXeKFxHOeyi71vcyXQv
oGncLYIni0KNpzcxGdR7FA4G+evRbRv3A6iDDmD1544twtf6RBR8jglUKAIjXRFd
BwPbNxeMcgEKPa+jnroRzRnKSj9tK6mYNE3IXPNOagYd57NEqEB9Tf6vUcSeYbeO
XLzBnx4HLtfS1dCu+LkRW2nR82ESwKTf6zwwrw1ETdQtKW0rXm4OWIM5NzYhniWV
wzp4rtCyl6DXInX7nA8IsrqJrdPSXWfS0E6oQmsuQhssnRtklfGAbwEa5jJ0QUpu
c1tEBxVpRav3WOFjVHeD9G0foVYYSa2Gqfd+l0OQfJTDYYO4XIbYXDhTRvGfaWoH
7IeuO8GONymD1EmsjaIFaiSBF8gii+Y3k2b15vR+0S+/aoZi08VpVpEzreM8pq9y
URkSgeEKoVtIe/zPyI//YAnwsrIyn5or/mRrQQNQ2r/Y4Z5MYTKF8WVEfEpADe/N
He007AvbVfHyYgByS4zdmX32j5Gnqrujem6PXm60VmTFx4XuBGS7RUsxnfsO9N7R
U6HCThxB02xdTmw0C/JZn+9sZY8VoLYlcJX149m8wTbrMd3CuHtLDXBbjxPjzKQf
iNNiE+TYQoqV4uk96e8OCD2mVlZZV/kLMiPf3O75XHnOi6w0kzc1equzbdIzDRSm
S7OgfL4sn0I+Qql29M+/xGX/9b/0vlsoMknBXh3TKY1/KqI98uHpLug1q1g69iLl
eFMbIzQqGBy6ApxjrJ/00IvUZ0skfNonujYJB8bBCnWytu1RZIPuTeXZbCXWe+X/
BbK+GIAGdit/HJWvuloqRa74/DGN7ncIuXltyiFGBXrEn0g0wJXu+tZhb+G7qg5A
AeMU9whgWCTniLKUE3x4DuKpUavpAkYo5CcGhLjeDxEMri+DUqLeSI/+TnCoqrOt
6Y1ER18x8WtY3Yv448izqgN4KPDuoJ5gnMdRoSMSBw7vizwz0QnwkRTBtM6nzzC5
ruYnzqdLIFFWm8D8e8/n0Ah6E2FpOEav+a/uQZAU+XnzrKuYTb25AujNozT8WH7E
UTR+/gcwm99JwILUeSgsNVQ/jeOoLVxzoNRprYdSznd389sNMKOYa3R/4pqQ0CDQ
o1dHrB1MsFWQhqF8r0Ww99vHEVjh2y0SmL/lJygGNOYeKYsdRp82y6BsmlvGQxwJ
Mg/G1cRB8T9cJGWyqbr8MNWpEcaHp8cLD2h4QPh27kM8E0809FXPouP4AeqCs28X
Ca3iOdLcJi2lyltlb8SLM8jWoIqXQ1USOoMyxGHZtDls6A+Od14bzjiuf3iQ6/np
6MR+QRtS2ubPJU6171NEem9Pd9tR5zHl+3GwSTPLgWtPd96SLJkz0reNKouIw4kx
yFiha+pxRrhOhL5EmClqqYSMC+rS6dMW8KdDhkVOBht4KUtjK9arHiUkKPMr9aqG
FSqKgyYVF6aZTZBW6UF9yS6ZXVoaRe3jooXAOfvVz0yLU11j2KxLJ+04h3K0Yb1m
eW/v1Mm+MYDsmpbNckD3g4iYAV4UhSFfHtpTqmZA3fALS+qk6UzFkFrKhQSk5Rud
1/SBCX01khg+e67BaanF4V9sMLHBZroJzY1MtCgzQ8k5OyjpJir/byyBDNHPk+HN
ATl7vxYVZe/x0uQiYp9iDTTEHiUC5G3v5ulIsJ+PGoXAu6FGC6X5mKXbxlTOuJf3
jYunHotfYVP09JL9Va23vC6bT9ms0mp5StZ0o+/cZc4ab/ollgTPbUtxFm+5pFp7
+MxYRl78+q3VUILbYNeW2qr1ZdI18EjvlkVy9wSjwk3E6Rbg4RYaj6L4qbvkQzPt
nVnoxiMZSgwF0QfXEGPp/1YKcuLF1st1fzJUz1xMJgbTij9C/jNar+HpkrSgpuFP
Nu9N1umRWtThlY99W5RHR1KZqEnYJoqsowiVyyTPhWutVeE2dGoJGfAw4kiv/X6L
Jv60gSGE3guGfa1VQzXKE95+GXj0xDYjmgKtfiLF7obsYNl6BrddQAjC3JOCE2UE
5KvCP6ZS2DUqEu9l2MBxPnn0XtDtVZQQXz0IWi/+eW7x433FIyhxRzviuM/0nS2S
rBgye7vgJlJZdyIu2eYDRM4CAQCNTEV+VDHhKvCeC7Bcj8CfxNHGnLdMpA3kqjw+
UH8qdhe5PCGXVilVIHGWRQMlkR+XMrBoWRsgp2L77jy451GRtVfhzwvugoMim09z
Cj1uzbdAn/29qN6ZHTblpcWfOWUvsJuOxKcW2riKx6tQGnhZsKWUenBnOnGY0HHx
15g0rmjhwB6ALeOGmareMLlko/sRKYjwd04VjQwsa3SoI9rjtzBO4ZkbTEEfaIT5
ZbYRhr4Qp5ZqHxkBHFIhjVsuJUVPrmLmHnaVuPVIusvydr5VzdX44qEKfFsfyt9Z
BY1hgRG89z0IXFD4VpQW18lS5KFUirIOcr6kmrIiB0CBeHX/3UGW0I/5aGNAfDpp
bhk3IA1XUJ5fAfxZ0A3FY+9TcQBqMuzI7tECXBsFyMTQW5nzqh/C572DadiRbu3S
9eZQQEiNH/Hnql31yx5+3EAGhvO7geKTnlSWoHJHQEFeYeG8f70OhS0eeyoYv07l
BX+TLatf20N07+xibglMXgt4jI/gSnjWtr10DdfumFce8BJoRPS53B/3dr+D/neI
E3+u8vJ2xqK8axlE6CVUFNje0qfKhsAjBvHffu+83XJ8upf/HcF2RglK0jusYIdj
uwIXDryze0EU7BUhQu0YpMonL65yDTfjsQKB2clCdvSYaPQFHooetRs9l/SZU8/u
ouJkLQshAVhG+bubrdBEkyTShg/hBAl2N8fSg5zkVC1UsL9hyv2uHUHlT7AjMwiV
kgKlyF4SktNOTNH2ns/G9bBQGEhx4o8/g+m/smFUEnopYxOu5x6ntnESfJPFUttN
gN8z2qbBdQjCFenAaQwqPkc/utVQPpn4g9Fk0KXjU4nnZ4JXbVA4RPfexL16CovV
ATadm0KuuiijCks0tUSiakLmgDfbANA+B8m0cK8TNNvqD4mxiObLBxYRV9hMmTXE
H+vyOP+NGzM1dRGQyKBt1ZikW2tFTMmb4reMw6t7J7qcshyO+OJpi93D29M+NB9i
zr8eMBfxrPcyErI1jHyT95J/bRbZn8GrDdzSf/WS7maYIOqnAy4znYsZiHPw5oak
AFeBm318l1MZpNOdRnZe/oUrE3/QllhwHVY77fbkhsxZUfIbl4671EtgDeBtZ/rl
ZQ3InScMUSZ5zrfgzTfWiSeuG0TVwrbLW7ghXD33sUa+5EyaZglBU+EfVZnMjTVY
GbQ4Cbm32CFFeSm75+8nx0OdH+01jWSCNAFN+fp1Ilmu+t0kmv/APlMc2etCTDXJ
+IEd3MDuxgz6hqqsRpkJ8UNt4HHmAXts+hbyvan5sfpJZEdXBQCNjZeazkRqvuQY
MSd8hxbq/BzRgMsJg6UWNHpZtseiCE718jSqT3G4ZikowvbPXOBtNayOWfdvxllQ
18qVHjp6ELDINT7Wj9M11qQor/Um8jVvy6GJyqWXTjV3hdn2IHcGQq6VN3C7dmxe
8NQHaix6/vDqBf9CBZeVV/VHndDhpJ+usbgDOBJFrER8ZP7JJzqvMJX8JoBL70nG
YR2ybhi2pMpNdpVpJC0ybsj9rkgiMSDKuCVOO5lbL6ojhsqz6x9H3ByJAM1yUQqv
+JE2D7yLkEedCNVgm9RFcdjJxL6u1ChwK9uAkt5GoFsFNx4Lqdh8ozQ1vqjwpFR9
Wltr/8F+uArcGB36LPCs9nmU2BeZAt5D1wNSpVVMbT+OqpjS0zSBf4rTucG2tXAX
v0ANccHR/gxkECMJLQXrNutrZLYvclF2Lx+MHiQM6P8RMEfkkcoA9Rq+XeODBk1/
QeLaM+D4jbQHU9NUl5CwcRkiyhqTXx0kLC2Xgf8QIsKjfa07N8agCI5LPMJzNuOX
gcB+VTxqwIGXzSxOxEV7I3BBT0RTXPFNrRGpXcevFroXalG3GYTkrhdKyBr4o4yj
ZoOO/TKZzd4sNxEHXqw4ZhDDegP7M77jSewErJPIZ04JlkmYBKGuQL5sy9ACnNP+
iQbmSgUkZ0nsv6lNsYh5Wv5gILuXrlprWKSbshSYIxLiTKGcLT2j0wp45Hvaa3xL
MDZEYm2bRBlaKAUPMSNw7gdbfVk6QC9fHgHjPxPCEEl+EwNWqMQAbDD/ZwlYZR+4
7Poy5vgAVmYaW3VvHNb2Be2bxuZteXZTGsuiNEB0VZEFfT9NwG4At7AM0c4jseXT
ig2OgTOsQAw3PX8HZpCvJhnkhM7B5NgJo/VP72ZwSGJ+WFoOQ8CmORRvvoYHC5SG
BFmJceolpj1/sM8qaSsqmH3IUeNV4S26nLy6ety9lPUbDePS0swVjPmmXlCxQo8l
9vhOQL25BlN+yeCtpjwrz0uTlhWH32BH0sRCHPHe39q9AAOZ9eWInvg1nGXxqiuq
AwH6Cdtu1GNwPPGm5OPLK6kD6Ot3mvrtNclmUJ07xalnMZ16gVTQxXBGcnQ9/TVI
zEgisYpJujevxIPWe0wEbh91LZUe7qNPRBu94bKiob85Vg8Pd737Oy+91So4DW3i
VRNABe/SvwX8pCEVfaz0NB3FfOEYc57cl20lt1vaiJJr8hb7NAB8tkx5Nr7Bn3TU
Hxi5U7PhCjYw4ItXNlY6jq9iXtHvyeUo375ksHQGy0VPpX8UG5PQJUwWBCrhqcHK
u4SYKwzCJzXBkyvP1PrJY1GvdsAI1GiWaMf0xJyALQ8Wi322LMkjgf6EoJfFCf6c
VPfPPb7r5E0G0eSWnjMQsy7Wiwuz2hHEQfmLEM41RRGbG1A8aZxaRWDijd3ypOCh
jsdZhqrhX0epTIiJUyk90L5J4N4W4Q7vUb6cp3JXCUVE9u106N0gw1QpWXkUaeXV
I5mqNE2fMxaJEPxErtoeezPKYSRFFFKMSjf7hjZxIdtXY2qU3jKP9hALI0EeqYSn
6E6MeFKFi9QoCZoK1D9N3fn4oiE1dk6MsDRzdQwLRFVYnsqmc1kPC8ok91w5sfUZ
rXjyhUIcAm//vAQInhqRsekAWb4vQx/BYpPmn5Tcys9i9axu+hg59pFsR0vafeQ6
tuzll4oTznD65MCe/psZCUZ8qz7Ot0JrgdchbfEfo2UKRYcqDjUnD6xe3hNN9p/D
zNRKXU/G8mwp9jJbug35PBV+tjhsrRDw5hDuo4O8GHyC/dIugemo1J5NcMjLrheQ
maQqJu8ZtLXkA7HItHBhU2eTm1/NoLj4E8cTBGZNR7Y81WzdU8h//uCCuge45J3I
H4VjkOqcT/jLxPJDXFU+pfeeaf4T2e+fnUTt++twKfOAna6L3TlLTEikLEEX1jQh
Ag9/p43y0EgVbXuT/P2ntPL7YrEMScGYlRz4em0CUtHKP67kLJftP8Z65KZw0TVN
I92VGjOK3QDMHy2TG1qP0q8oiDjlfZA3ekeGPd+EFp62fSf21n+mrdtprBVEeKRs
EV21iTvSYHPpYFhcy6v167ztjrLLkpEP/aMeVpx8itYoKVaaXGed1g1BrFy8OdHp
SQhVbZxyDSUgU1urQSa4Fb+sD9FnWzpslMYhdkPwtN8xcIv9Y8SS7TwvvBDTdVUZ
+M6mE0KsFwK6CaQqAnIZFx0m6lSLB9twcDqGBjmGxPNUApjAtPTl7vsWwTPJJGdi
Ckgl3/IsFtOCn4RlofmrgV5EHoVQrmy0D9m9HR5naTld/VRWlF+zmhvCmdCfT7hc
VMFLzh17kj4hsRkWHiUyuJx6D/9GKZu/eAoVDOc73cTPSm33OxFDxu6QZCgf3xUT
azz2raMhudIMOxeyvYilcaBkVK3P4NZ5hPTtdRYoJD9+7kr+fdzh/DMGcJPJtOgR
aKyUc1B8zf2r9vps2YaQCLPyVP7VwOb36q0TJa7m0gX8GDSMRY2Hp8i4FWrFbdmD
hYK7UpLkbHxaF3NLcHw46tNLDQ6iNDI2SYrIOBo74/syFPsB+A7wK3CgBXEYsYyV
25O/5W3KiKtM6oO2Vjg+ftZ9Ck7THZzubdwsQdubtlezL7er0NoifpEF5KFXgMS5
8/w2/WyCF9vSc1FErU8+nwYSk/JTawISFRnlzEKgbOiBIkbbBZMcF6xvgK0QKhU8
mZc46v2dq265Zj5ydgNsZeQadepogG4MGAZfsbqh5WGtN0A4mLKrqnXSCt0RUOjf
ZfONGEjfQ7jQOupcJPOy9Wr6rkO/USW3rBqMd8vmV9h9InYwBwOxBz6LccCIyyHN
GF+beyUN+U6IBrJZihlstUn+iCxY5yDu5sMWpdZexZ45/2v8qf6CAfyyi6wMow2I
jVs68J0DKZengKxf8H6XRXeSZVaN9pFTcEJvXbVbgtuUZz3QbBkFo7KkYrZwB8nL
40dyJ4sp8e0lf2st0X/zhO/bTsjX0Z3QsFQ/NCzdKgcP+tzW4aOHF1MPZnskwJqu
xJNuklhE0SB6biugThM0ckbYG1OWz4pQ6GDoa2h2uMPovZfagLKe2PPYy9CKYcIf
ewt9vIyntN+s7nHi9hcDg93kG4UcO+IrlDzcEjYMexezboiQdo7BzXMTQs1M4YMc
wbRnoJT5chzYCT/2aBv0mUvJ2Hda1YjlckQf8MlepzUT3MHLQNoxe9HDRKLr11Y9
ELBWRCRlWdVYJUMdqxFvv1esbVkY2qkXKGwrGw9puB+mYAeOrWuQgv93iwPxzbI3
n4qUCp2doSIg53mICiTDVrHZmdzjtbij5WQmBodhDB7mhWZB6LJlZO8fxoE4rsDK
cZol1SlePQnyjEaHJLGbksncYVVT+M6bxYJPZuO/OVCpt017AeMGxrt4tbmKjyO9
f1lAGObM5rFapo8foztuo1eCrhDlfJYMuBLAxRlz5Tno+ET8lHXj57JzzLFKH8pO
geGSVp50flJM+0LyV356rctZ9+A4nNLSPSD0GRiNaJehhq+BAuqU0d0M6Y5OvMGv
r+lQGKcjDUvjtQvsHer0aP4tu81MwBeqnG7apecNGwGku6VTHvpH5i4FyZCai+IO
5B3Y/MbFGntSIILOkKBG+aIBCQZEhdaJG49Nu0v4KKRXPj0DEq2VG0M0rED3vy8U
33ui0CgnTlnlEhAMHdhs17yQ+4rN0xBGJQIMLveBn1G11CnUoysN69RBAoyx7fsi
BO/MPPxtKzfSrw5YSzh5PliTM91e8VWdkQcaWffZP8sTSWu4nWtyIOaFWFN+qqWc
YfM4bYnNAXtZp7v0lASjTc8/bPeB00onabVzbmiCtWVARQxurxYiRGyBBdt/Qb+L
XpcqMFzsaZxGF/fBD+ryvVdLN8w5wcS/wJ+THI4SiDg7S2U6SPCJZDdCvrYjPia6
RxB26gZjnMBpo66Jj2bGwOYlhNUsyClxp/rNTqWBrOpJRXh1OO8if4/6KLHNeMnM
NZFY6J25P4q70x5A4paghx8VZMN0OssxOnC+v2VkhBffTWsPWN90G3VkZ5H8Og0P
JtGBx5lVsFot6jPsK22bD1/qZeQDj7hpM2Ex6m7BDZmIBAACSRb+WPz0vjiNIIOX
VyLey041urYTT6xvNRKvUndXroJQ2AnwD1325gxbiOzTjNEW5k0UUR9ahduCu6HF
hy8b7ZKVuULrAG2606iU489cJSb0sPJplr9A3/dgcnGyVEBIOZg/tU5roMSYr4Nq
xkdSCd7Wg8P7Zm22Z0bH0WkUyhZVoBUyvqOsU1ixZ24nAPTDC1IgLklnCFgdCtxM
Z1r2npc78tzfTlVyAa8kvef8kD1ctjy2Vca4iGAmo9E6X+qlhkkreV3e3fftIndF
y5nsrdqnrA6VSe/9ueaGvhkBHsxYDxrZ1N9CMhU4fbSlTHXh5Pskud6c9mYhM/Wy
H1RmHj2u6Mm/4Af8sIiNynR453l2yEwjVCPOju95jg7LFLMOyjcagKLaUPdCoIGP
PPSSd91ffSXHtx0T2xIx8bv2F6fX5Xd7B770ORYY3/8TKN1r4ch2jyKIAziPHyWb
b6858UeN231h/mk/curVl498tz1v/vd+eGCXJWBklObjHSgfiOLjWZVjbmw5yDbV
TMy5DPn/7NQBQXLNpW8xW50+UYV5tsBSeFd6dfsfAwp7HCfukAIy79hlbh5wrvOY
VMttZMskULD2UnNegzsJ2hkPTJto/WwkQiMdMMxogfc9XAUblcPsec0oXny5XVIP
oigZwlGhoNA0u3V1mXNMT/MojlqAeRNd/SlP5H/0d+XuH9MSaUG8Qz54bEViFVi0
ZuWqAfoUF8YA1mNHrsXG67e9ovPytYrVPXTKqXPExvuWHHDQWdpoEzOj400hhJIx
EEknvQjYZAk3Y4qfXZTNAzLibHiFuBnEx9wzDcqTkLy1YgEWGjkgxu+Ynp9NP2YX
4nMcf+R9qeGnJcrZB77zT76mGXbXskx6TVGIFOopIAtRULBiHHtT88ieCS1aVlrd
dhExjOZqWk9uM7E0MU93sPbed7UFmpc7Z6UUCL2cuu/LWMNxhBlK4/ZOsEJmIyF2
xcr9AG00q3ExbN101zAUSCWFdLSK9+bcRQbe7I08KWT4D7KpuMX70kxjAO9351fe
G4PJ794mJRGnFFlTVYAnbHYBo4Yi5LJA+uXro9xpOHMcSZgde2FW6Psq5aUPM8J1
ZTOTzU3sjNCWHpi8BTJajEIe/xX5Yh+wC4uYovFL3AMhxdwBbjLUwIdMJKr3oFbP
u2JxfWFr7gRMyAZaIf6SIvx95alWUtFQVIF+qkLhb9u8kdkrlhFKOMWRN/ZFEWWG
KBO1TnemYWPoWH5BhNWyhaYTfAPSAqXo5/Yh1l8p8TbVDQ//8cQXruzQihdYAO0/
mGLlza7RdqnoqPVrzWEjGcM70PbPxCuNYNZs77HNZQ/s9bcI5WnRmJGnpZlD8L4K
X1a7hLT4N50tkpsAUoQ5ZMNOHFNRI/6Ooej9W0w3nsdnIwVuTNuSTcY6XA0zeeCo
Xbhkeh9WpzD1QrhYtMTBHF8FFg4nmPlDndgcI/HhEC+Bw+qbzpf+3b8zRSWYlnMJ
2g4UMH3GEdyB9WUr9I5sdRtj0tmPF4wRxJ3RIhMr4VOUy2Cxev3ji8TG1JNLCMYf
uVV8Q6UCU5lOSzfIOVeV4S9/mkPXtsf2TLecflQ1GLVi2QKjeX7q1RSrilwOrKiO
PsZw2Sxfm2e7DPUasY6MGsmttEpZlpP8Bhk9B/DjMljVxf4nDPI6Pe/BVwE5+wSF
4jXePot2U8KRA4+s+Y+3xxQxfr+uRONhTUNwkCBFjSDbRQYKBPjUGteMBvL/gokh
yA2eW31Fmb9fLamhX0mJuMZ3dY9cuYQNcCKvnN+NON9Cpn04IXrlOfR54hO/74+N
tTgaRrGFZZvrwOm33fwijpiW1411ewBWVcPilasboyD0IuYlwXkE3BWR+BJToFAh
mQa+iyd1VBBizofoykB4fg54IQz0pATsj/QRySNu0+RV6hDe6mLhifqlmOanCq7B
aUaUs79wQleE4bV1C7QTrCpfZE7S2qZ4V7FcCRgTfB79r/LeGf0FBn7WHNDEpzqV
2fo6TQSSQ0an6CPR54hi48s3Xb47vnOZqcMSOJv8wypjr7Fg2mR9C8FQvg1oqOVg
fr4IwalUeaugIxq+/2NjqUQlAkZKpoiZ/K5FCLq3PFlSIBDq07yYF6CWFaYzxj6g
13Hnv31KhAOjR7eYIOc8xN5hbed+HplKxc2jh+KutKGomSrcb8kS4mJ/M/nBA0OQ
LR5vslc0oywxi+08oeeCflfif+Z83oqZdfXKirMewnOTuggUacsowLWdT7rrAFKI
WmnRAjASVu9RG7WNfDFgkDoRqWYFQgAh1DwYluMHAKjVd5ORmRGLtJdPGh6uMfKX
N6AWJwGCBp7E5ZtMhQ/S3rmo0U+T5EYhFXh54x5teHhPxdPFqurFqNXERrjBIxHl
dOVVUXwBEpa6sevuTqY51N0VdvPnlDVsSQ0r8azXoTj44/o1xwk2TNJzCTK1vTnN
rENFAiVc1q5as26RMNNgkjD9J7FhFeOON5Caz1axkezrbg+1ofLlDN2PxZtKbgUD
dAWXVR4YtI+SivHY3H2n4W/vRtIoIlGazCWX4CuTrHu7qd28p0udMl2CMTGjtFs/
E8hhFe1y75fLXxQ2n3EHjE9YxCoDv1jLTnRrhYlDs4Y0rCCO6V7QzX/MdlIAqkdw
DP76Ekid6cV0LDOObdI7sZuVYupB8j2Imn3pgqKeQ4SxkGK+DnjLJkZRcpXZFdyn
WTmEa60gXFv6MHKKuQbyY87N+1+he/HIFhjbPkwxTnGG2mmeJSZ4jVQMaDg3IQfk
xUhb8Z3OF+B7N/sy+/hyxFvPGpv3aA3WmFl2uJkOQJBIBjINrX9RO1pi8pZPfzZ8
d8cmbQXNZsCy5H1PNMKEjT6FBB7ggDQci2PydU1g/SaAHyIbl5Ykhaty+ijzrgxx
U/smsxUbkSe+04BtnTDyz3i2MtrCVJniD2UWZBF4JeENDz7POmg16zCSN02+iBmO
xchHY0lWNbw3g9iX02+ZlGgj3TnKpeDAAgP7K5Mn496cSM2NRPwfaVWWB4XayB5u
UxKXpXCGnCViC1E0or9+HvZA3TOVt9FsXewQ0tNI/Ofg5EMfNjmMutZVkTweqwsO
Yshls+1rwB2yDVvP1uVgdggIfVrklPrhwh2EMs3TBXM7kZHxjnk5kYqHO8s2cKtt
GgbxdmRkkaAc76RwQUFzysHOVx9hvrMosR0qCduCU+lJ1Kjq+jOuWY7k7n7MXy/n
+pgUI71qrWFFhmzd+L+D7vwwBKoo0dVx0E1m0zbiohCO+l0/r68PVQUzun5DRFZm
ELeIGeQNFchWyXxdj8czf3g94xm3blX1smv9UyZLJGwChwWgMk5dEImxf6IFrPUR
bg1Hpn92Zwf/QUAVuwbZbeqjLZuhMIHPiuVk9Sq4Ov7HM+5crshwzfvQ7XfctrCB
qauHWf/HnlkZypoZc/08dGPkEvG8xjaDXZL/MxRGoYVyBDjj5c5FuTNVvE2oTE82
qtA6hwckS7TsoUZ40KPNNmQL4M0y0C85CWHT8WNfX89Am/tX6hYRkHyJiFX+dx5c
F62Ex1/TTeHPMeLo0vJEq+bQdqJDhRkEr1jxPQO0Ozrf7+8Jq91dX3we5nV4AZ6Q
85FNaxE1+T6KP+SjLLec1gwz5RNiMurlBqxEz8QGr8D8K46Y4dkMb0RWWS98xmAj
cIDK/iB50i2pvb2+qFX5wTFoukKhPZX0nfFLyYZGS3dxlbQwdGCjytZhtK+FvHmh
hMYk5Z4vwyakYhTJ2wNCdo0K+6bYbtCGOwyO5IUemFaF7LCLak35ACbPSlvbgnUh
jG9RheOAtWeFdfMzeq6KqpdI6w3KK+EmBd3bpimuZMO37LfTYKwcx45BAWJ9MBuE
CHs9SN2N5MdGgabdLqxAZIr8rDFXsn8VQRqwnJs3oGWVthYlxzvUlrHCZHX1Fugt
Av5wZ4hxrHYlC+yh5MUHIsGM5/XaG8RPBgpjoGpnch9CNz9x8NDV6sj19KGyNacl
zzdJ0T3xg/yXVe2HydhP9iaE97xWQsWfGmJHaz7GazTCJwFxZHedRYTBMmeOUSig
B9pUXG4XLB9cc3Q+R9ysUK5zfQEfiuzpekOP87W+WIfI0yJuGk7XKEG6BScXKc5v
HRu3KD+QtBgnRo7BtOMDQbAtVKR+USZ2xWRdiCwfnXbVRAb5HwQh0++RGK1G3+Fl
l25heuimkm9GQkBobN0YtwXCwo2RF7LzfCgljN3Dp/bSQQj80LBThdw3uncwm/S8
QycUkFTBlalxasJKwXgcMMsRoit8sIzv9UEsYiPJskt3N7kD4G2Q2C0yipafYffM
75Xg0XHtAnh0i3NQxZ03wDpsWBx9mBaNVrlzQyLHuDuW/fwzCZ2/4Ave4MeryfAa
GFNBaMXfHdyq8XLJY6+S12SGAMh7mPUwF5OQNz2ptOyWhElG3q1Sq30rFko+3XPR
xEW/xbgTAhpS8N7g4h5eX8iA2wHKWM2kuUeqY/QCBm88rtz7/cP11ggX6JdyHgVw
MP1IS9+JkTjnMCbLnjEFO9r/TRhtkJtMf+L1XScTJl/fJG6TXDPbeQJ12zGhDR/F
LJlvmYhizwuG98SetJ8CVNFBfMDTYqwZKFI+eD9igZBJg3f+ag5oL//y5lgrBVli
bQQ2iQIpfK3jl8/ukVWFtlmZtjzndBJj3mnCj6UljAWZE72y3zfYilkthXiLGryr
tYRgcWBOk6ovEXUbISXXqW5AOLe7ZJiN32K2nkD7B2v851GUvR6DtdYlbiljmWrC
6/K2g/tx72VdqgBvgDWfIA+9MVpOCm9N0nvyTA0sQsbQS/Qi5B9YskmHUyxe3K99
1zkdihz0DnzJghT5nG4ok28V/9/622+YcT9ZHihXpb/Lot+F0mPgs4FUTw2YJJCA
qTjV3u6NIHS1bFKWHIZ7pIpQiklQjZG6lCpvfly5rng5nPPXvy5rxGloO8l51yiO
u9TChPKApWho3OqCGeQonUA0lTU/CsS7Lpq6L3Cl4b40ZIN+4pYXco/JUFVHpet1
9W5pvKGmjVwpldOyuuXKWLJ81st6YXtivnuJ6nzox46RhaQYRZIJ+4wElbc2A2Kz
CVGJpTnKvG0vnh/ySx3X/p14TqukLOYoydVIp6o7Buexo1McOA0ZZmd+vMtkdnat
bLkdPEwBgPhw6I14zxizuuQCKLUnv7u/kel3SU8HSh8i4edUDQW1kPNVVD9usM1u
ZlGTa2EeqS1fWDDyaYHFWdj+9h9g/0doOR0z12hhAxzeExsyILq524YcBuWfl18f
g09yQob8FKY+atK5uwboYF/hxSmFAfJL1PI22V27TSTvhVgBBlLCBHVEPhNtklGD
UGnTrb3hhXgD7AcU1HTYT555ggrFKRQCAJAjMO4mZf+Vlh4/CtHWJLPd2VNdQtOw
SjNAR9jS274ojpq0ikQM6joGDEJbw742wso75H8+EoJubPH8pOTJiLWHB7s+Pek/
NYk3U8xj55rokvTVwu7eNAGNQfvOV7Tcxu9XmEgYMulCeDgrV8cbLgtWMEAs450j
eZZjSRXhoSZO0Njw0meza1mbzmLnMrZSTazJXLhozuwGO3Kee1ikEik3EpKKylIA
AYO96zLdufoFMNhzWYxHuhB9LxZwhjYimt2Ti3h+9huev8dn78x4Te6xNwF7cll0
wTqxc7Eg+//kh8Ggb2/LUS9VzogliyRJU6bp5Bw2dR3uZcGl32G2eF0q87bvl6en
vaNZRw+W0xcz58Ug/Zxl5jjx2iRfOLK1ztXedHuqXKTxSooedyIE6CDYPCHKOv6E
TtdccCyZ3i/3EJY/wRNxkYCnrMaRzPVosVGH86ChS3SFzRXegzp0PAZYrhGXFt5P
OWf8B2U54i9bFBMWS8h4k7bEFRwBhWkqodyMXfh77x2LEre17JGz8F16NLDIWI8c
JLCp0RVfREZoLfqCx2uhrIVf56i2cnuu+DAERRHn78fji9lA51JbOhvcfHRJeJPg
fySoe6YfJlcaEryOpX+CDwQo+u6mw25m8OYRphQWXbTwI6sKu3jqEtVtNN8CYdLb
ktDpuCiEqc3SuemlTJhzs4hbedmYy6KDRESsDS4YxjVPbJKExtjY/Nrd/bNFL4Fn
WuSwPETeHGhBhnIP2kJPD4VcSmjjyCl4FTpHzlUMwegKO8uJ7MmQ8WJXQdR4V463
9u92bP+zu+ky1+/W6GyoL2Z+pITg1OxfXx52njwHwxEkiFkv5YKKL59gOlTBssHy
GuSzxoklapNq/ktIG11RrVsHsMzN7r5FJUvcrZ0nlYkK2pTKBM5V4Y4TRNL+Ik6r
vegb21GnXS5D6puH4ZG+0/WiTk+RSpYdmwA/fdVNQYhGLt0UYhKiGMyAwzN1ZV3U
K5NPMXzg34aJ85IqCrzTZRrhPuWCW/8sWWSBzTDRsZ5xhVHmC0yTgouZFHHcLgT1
DNAVwhABCYrnbssjEEMMUUksUbkQ9MghoqdSndP7F4SeS6Yw2tHOBxOmibP/pdx9
URYCj9PyDLRfN33JPVNVU4PgLTb3KmZhovIe0w6MkEwlZijPPmTX9N00ZEts0hSW
QaPPPOIuqugzhWrqMgIVYknLWVoMRzgfn3FPF76B/fMQPPOrf9UEqykQLApCxujK
xVXWmvsiSxkQ7O/4CEjYuZQOphUf8yWqPCQE611ZOhYctQl2ZJZ4CeqylN5iNKC5
n49uup3Z86sxP0/3i1csX4uMO1bSfnWe8n8qpYubLYoSKbHsDdB2EpmuCK96u5mw
KY2OpuEmHZIpVdMP6bodfb9cuYgrCKbki3Xx2ECsPhhg2aS44RBF9hvtyqQqJ4Dn
U3PqtbGlALnMD7BTLDSCLp0Wxcs9cnuBZizuszc3w7uUxuXqYJ6C8JUcCz/Nwjmq
JGc3iSCt8UB0mGntWfH6f7apGYTr5ZAo2MrXszUrGSGOinrm/DrxdpSToTdR8AhX
/2jXOl+JWJe1WpZHty4IqGY1D1h9Ls4/tRp1Ja6hRgwhlkq2fDogc0r8VAxJ3KHk
kbu31tW8u1pKb7xWrkChbxPqQsEGVXE/YMkQZ6S09BjuNpoUA2xJdyX2AQWLySAF
THEj0N4U3NTL/ygGK8Qw/9uNpatlQ6vicu5E3PNn1UCMPBFYBmZHlVRTpK3L6tCC
jI3mgHqVykpDUUp6ZxSfYUcnlDJMOOeS21V0C1T3APeqVIE7efioxP0hXnHwI3J6
Ra4hvUv45jch//H8qKdfG8dOyyzwDlIYdHi80jPrQVGU+2NHe+GuA9kSuuOhBLWJ
dzxJO0DiKCNPpKYCZPMywaiLQusIwvNPFi1qxyugdHCJFWcHGAEmPpYIoVQNSaQO
W6fq8jrC1GrECDjYADYanzm3hxxx0vUzifYnZ3Rtujih/tk15zK3IypC1nyeLD2i
yu5KiYPcAjLTKMIRUxcRAP7FqKWHFPfdd5VOMpvQjjtuFZLI1h0QoH/WqzRxbDaX
Y1GEKWFIH9iUo8N2nMTXgTKQvr5ap0KrGFdoXBBCxlVlxI7LQQZmsi+/AaZnKpEs
Z2YYsNq9Z7HkPTsH4w+vcLU++0pmtjS+JNX8ewNJSCmA/Wg6BtrEAJP+y/23DPLP
lprcOVbWXacq5Sve94dNYl50tBexCVFaZlLo7uV4CHFNAc01yF+FAIFAC+kuVgLL
UQYNkgFtvPj0twUgsXstWSUoE1OedqjFbPn3C1pIPPuQYzF5vWODt+53x4q9ToEH
zfz8J276dDJE+EC9iC34TX9871GQvdDkBY3VuuEIqOwX1IfR6QMXR85AhGZieQTk
KaehLL+Ks+Gk416ptgu2ywQ62ZTXfm5LheVnoMxwcaBQCcF0qbGy+VfnIWdPsBJy
l70rL0DEM0IEIKJwH69mNnPMfZPWdsjLwa/cBySLSvAMQX76XQSgKbi12Q20i8Vv
atEwq+jqQ+fH2ejxFM1/76jnwMOLnnEeEWi5XhYmeZWBwSsRzmTpBHg0CZDptaSK
7slJ+vrHk6ux+ZN+pbHLulwY2pBXNX9Pv7uBM9GEHeJuCVyOzXlXMaab/3NdddoN
kYJbjAU8kPsUR5Vcg+YQwXcLqQ6SYxDikf5kd/ZsjORApaXfbaxiy5Skp55b+zWk
/KfPQTX5qPb6tn1S7URT2DqhhQ/Dg1ThkGSDXpEf6h8Yt9k/cOYRxkbvOrqUMEHJ
Y5Car8aNh3nYLxl0dINBoqLRnWREknzZY4ACgaQqNokayNx4nVXzoI/Kcj597B2D
DA4J0rDuEhQgMccmcNbKpbX2XJo6TK4kpLa4duWjK7qeNV8caZuSNytLvtf7W6j5
2MIH98IFnwRztZ4F7/+zBHmSY6NzsxT0ncgQm4F09qIhEVTXgom0fGMY41L1GWqL
5uG4S/Ln+1EXY02CdQVACVe9E0qkYMweAgLCI1kioV8MXrCgTl4BgiqARgHD+vSy
x9LnZJ5j6ccllXYPA09IZ7xbTlLtkcswNKKvAZ+0UccCf0BMCPurwGhGcXzsAblH
9T/7e5fRjeTvumJz1Bra8RWdpCeCFFAUgnjubbcG8ofF0GawBcGLHj1zDiSjFVtN
7SDFkg64z019Z1tLgsRbjLLXt5/CWBnz8UzlSjvcZDsan9tOsO0lvcSXugtd3kpC
ki5eRnt5Ud6USgTyu3gDJUww2Jm0JQrCkKRA+z29unCuLjWX2aek8efUyOqAOn8c
5OG26Zx+Nj2e1xq0oPkSvAx+EyslKXDyKVG1mX7ESm6rKFVw4u/g61Z1SvPe1vwm
Qbt9nrqoO9DeCQXtyZVQhk4APEOWtXexfRK7c4/8jjd9LLJHIN+vTb2wAd6sWxOU
v1isvlJUu9hIqzSOowvMwa+AAdsfliUgCTcBBZBhaCQ5ANj73Yjo2RocTSOv6wJg
lSxZKN7BTH+LtxzKJzTfabo2cgi0XpLl30r+ier7C3c21AF/a4qRTl5PuhzdoVub
IQGuifbcX1z+jguRR4MFamepHC5J4ru8xnqngac8gKrJ5gukZRa6/QIa2/QlKlgR
OPEogwP89ct/n2s1LKKV3kpq3kqgIzJ3xOw2fXpWzWAsRHYg+pgBdho8ycIZpMk4
EceXEwNJxUkWY02QDP5xFdhhmHrVfH2XCgy9UtsBuJMtISqx4kx/hjL6938EYmo0
iQFo4TwMA3sNJkUXSBnVXW81/8bdzfOHm7q+W8k1CSjjcM07AJVmaNs48ej15Qhw
PX5YoeZ/phkhAAyOd/OqbzPvKmob5eKn2anYBUsxYzrx6p3kxTeAbJvyG6iMsgA0
lwZBFUQreicF9iXMckKlts9QkovjKE68P99ytDORvD917IV3u9wL/ZAsF30EKn/O
1GJXJqDu2GohWkdpghskCXzTGfWqhxS2BFk9Tjaacl9Mhfu3SSBIoONUCWStVNXq
kLS7sI91EoYvSXQdwS9J5HNFkbi8hvSWseuGORDnfzms70ZCCVVXnUvJ7AWBlRNe
PrnBJnTzTNT3q+WIL39QE6zo2dps4oKgyEV9LdvVy5To9McyVPApRlV1JwTh9JDQ
UeufcgQ8maEbDKauoYZZ6Mgp5nuhjk8Z/DwetQPl5vBrV9b3Rb48qsVW4oCavqHO
8OqJ8goj7OjySiyayfeyCGOShbnmbt2s9fmLo6Uy2KXXcrebrUdwfFkRQvni3g9U
xgl9NMrjYf9okJz/jgy/m6S+HVxpw1OsBrQF3pZ4eVA/oBxLaLCFbewIRZgrTmUg
4P8GekhmNuE+orMQm180Cu/dQ2MWsTDKQq9ev4gs1jI1/dLi6xSFXi7KDB23oXH8
k3vjtM49KIfvuZ9pneVLMxlaWcqwYoVfDyODh80jgiHDtETry8Ss+LOG0F2OliWm
8vwdc1esrazRGehFXMQXj6NvlIfpSrDyqwg3RerT1ViJv/t+zQv0NxDXtwqW9uiU
gxmgbb2Y4iO6IMS9qw+8xTGpSph8fWL7uMCXI6mHafsFuZa6QmUCZyqzl5SzrD2x
nkqpEzKxL3TkJMHhLc9gmnztFpE1bFCi5jc5nRHLWoHue3M7vxeUKKl1/DS/EJqy
gbWHI6IKgtZUk7rvvPh3T8PrWlZ3HM1IVyETcYGhBkjMmoYQSUjBZYvl+lK8E2rv
qWIohfDVkkrm9cjuORPQiqcZw8BzdI3uV6vdulxP3HbhH5KhzWcm2ZBc0GElsY4V
VPU6YIVZdx1cUEiZd3lfloirmmfkNQ6js42O7JnaeYFUEe8UwLT97JnBtqzu0U/K
qZnfnjAVNjWtJMwcc0W0gZ/APNu8Hhvv1xKFosx32CJdeBBWCvXJniYJgl58MjUj
lg8hqPnII6m5tU7QNJsFA9yK5R19x/z42QO62t3k0150GQK2yThS736wjaDGvH/0
8aPPUzJKjHfTUGVRtvjOhwRB2nRKuEEEdsUcw6pIvBqh00A3Dcv5/qO7OZ5R8KJi
QKNCE/LjtfLXUwEl2j8jwKZIxaGD/JaC7E33N61BUWN1Pwh8wRPoe0LALDgCmtsi
fGEzdTmQIQBQlGlWhwNuBJCg6FaoOrdhra88o7wA50NDs6H1qJ9iaUVvGALs1pM2
dMwkNhMA5ZwhBLlljBCB2kB5m048BBb2w/vVG8S6bLjq8zm8KJtt6f9zBobCaGaF
OrLm5GAf8Mwyh8tbsmfSRtx0V7cWRls2NsH2fBFTJXuazTE0z1KKVmx0W0GOsNT/
pHr0GNfclXyENgoFqNONp1jSAVZRtLoEYzRfoaKim9Ts/ut/49X41SmbV7bkQsuU
3RB9iXy/OFz2a5wpCyBEL/Do0+xgNvpAhMpfgdia8LtlJSjdEZfb/mUla6+Kz/M9
zhe29yVPPaU9PCtqESqGFFC/eFDAZn5FygkGGZX6T3Q/hLoJrL65rTJYEmo7T1PR
8fUv+bvnHNiWXklUN6TOgaGwQrbxezttaxgcJFhlWGOBY5d/b/QtQh6LARBiFeIz
NUes5bJ1tgM1nZaFTq9ZQJZx7eaRtwwIXqyWGkKi0w2+25MFSCT6K+ZkfcaUkJRd
IhGNQIJ42YmjppKVcEtmvQNcyXryL4AaHq9I6BhLy1Ah1Gb74ZnSg7muQBhcAYAr
vYvmkQUFxmNJles2KsjB/Mb5Mx1P7PkmgQy7wD+eGD6kjBNNu570zE6+s2pnNz+d
twUGyQpZ5VbXw3tiGvzm+HMttsLYJvhKtAjBvwuBdrCWqBfSfahuSxTJLFwe6GLB
rAQobbUErlq080MkMv5FJRilrBU8ijqFw2bPRSoQStKs9QhzjhQ8vcQXtdYLOIyP
yK9257nQHmspaEHQl1ZwF57NfKcWPFzdKm8wCENlzVH16sFbCK0YKQhHRo4TQTy4
yoMDatZrutwOwkuoKzrjtr6QeDffUnx+OJbk15dELMtXiX1yE1YTo6hJ6LKs13cX
lbpnk0FKpRFrmmu9WQMNI8yfkgJkpwVMiFjezr0RxdjSAVbwpaaz30LG8B/a6Yek
EvyYEkc6IeVLxJGsCFKqgCrOyIQE1IVUu98Krsf2oqwZ03m4TODXVGkASfFbeS+R
zT/tLxs5Fr+2QXYpXe2dxYhkG1VWFvtaBGCxy67TCEdnxj7ZXtPVk17bEvTB27EX
HbEaiDkxYpCwyWMNHhyhJc20jA83N5r0LO4Cte6Pdv5r8JLVJUK9WbgOWkOChzqS
KhDz460ELMF5B0Y6ah2nSkJuMsI5WJo9FlvFUwWbri1f77/YN0Jl7qDs/1/e04Wk
Jw6g5B+DMekUiDLU9fHP6RBHj3zdUob+u6AplG6veB7wAC5z2rhge1talw8Gyv5S
XHZ0YKXR+/i6LzCrBPcz3M9h6B5cMvTe3J9VsQ7Bv52z+uz0xjyjnkrEUzScZUvA
EpPpH+bzzOfo4rMHONJU8RXc8DdVaBDUCF6VQMCFIZ2FUbNILF9fBbQePodMZ1gS
BvEYl/U98mfhKiaP5ZwsiNSYZ0aGC264ATL7NAynRR+46Gy7YcQbvmilZqV3cfmG
MU+SM/QMMhZlMzXafLUPQaq3vzBqUX9jYrxA+dDZINl1EiAwGR9x3O4JtwgGF9Vw
9rxgXLUNtUXsDmrquweSkq34/cZTs4Y9vrYeup24cX7WSuCd+787AkSvvnSI9m+C
D9Y8N0cHIpIb+LR7vFgTebbA06MhvEaeEKvWpiouts30k/1IwoNQPf6udW+59rGU
42cB8WHt52pGYbLXpnZWwLvkpvGTq0acegPWCyCrUynPy9piH1ZA5/AOoozONxoF
NPoiuWnDVkvKpFVy8qZOXYgSGL3uH76pvLTfsRHSzVknT1MeoSh0kyi7XVWqcVQm
tYiHWWCYwtC3+7V1o4W+ZXUmTvZJDL0F3rZFzqa2B7OGqmM4GAOYCeFyYEy0tsRK
dSVNFNNn57DRcwyoeuJSpCeS56XDqJvwjkoD3ybFAIcR8tTqsfXylfL88vmFyTpB
w14bf/k/ZV9JhL5fNcBXOzkYLpWtyoqzmCtKXJi2wyg5oq9QSTVnB4ufy3qH9Ixc
v9L2RUZueQswMp5HQL3hZlmoPcNdKzRuEJDNI2/rWSMn+dR2zdxx7n23kJhpmsMH
QZ0X14OILlePM520mPR17OIqDfe4PvuwoSoWuDAeNCHLsTLlPwHj0kqkgkz0c8Sf
ne3O1gRGHaocgMohqHOzvoy+SesfQhi7/HNQNyTH0snlcW2XkmWx6hQA4WIVQqSl
LvCVBK9vMF8xl20xECOqh/kk9NB3xP7/RH20yUdHS2n8noyd7ldFF6voDG4EQOxU
iXl2Aey4ia7kjRUngSw4+G3iE7A4Fy65bWhudmXXiqTaphQAMjgQ4tJFbQ30OhOO
CuH/+5tlzIDaQ7cc4WyriNG5hFaI9esddWmhgxim+wG84wqvv9PbWKZdfGH/949u
D9lVflx1sTNoUi2EKbUqL/eP6YvkxE6w6seGiHg8nn9GCpDQXseOv3YVWNNmeoHN
VI5HCEMnZHdK5SZCl1dGSax5pMTg7RrnB+gKvBWCDTxtlY55l9prvsIuFJh1BkB6
BBt416kpRgAOanHrZdJPRDIqcLpvEYJEir924hSOwVfFKGx+HNo5H14e1O4vrllM
vkZ1Dh5NWp6uG12x9uRcgHPTZM5d8FvRWykuEitAb2sagefZWtNV3imzNorAlWqm
3ai6oEldQ47OKXbtIwWD/2eNvz2HBI2MW4Qk0Lyi55aiFRSEeuK4k3mgvYHSiuuJ
1qTywBwVe0Fsl1RfKCfCmezb6TpK8GJoKRv6SM47auSlZW3tUdCjlNctwRTsFLqk
sFjbTT2rJyocz/3vJMdgt5MgC57B+nDBmcvAybByHe3TTFGyLx7hjIpGP1efrEr2
+oAy1VxUicd8+T2Y8RgHo6CSSTbrO2gpNB3YD9VjFVF5P6LkMhyRVjQSpqXUMu3D
DQ6nsswRNxJQXRYd86v/5QWvK5qWb8FvdclReMgaMuEwxP3Fa+CBHhEMYBSQXk7Z
sa/tWq3vhYlmuTgAGQ99YKsx4TGcITRnpwvQdYApK8LgoGLm1GwlWe+z65BbWBcv
+Hr0qbPfLPkiWA5cYNjoSEzDvpV743W/xtB50nJKhadabZbp/ZddNHhSVI1pbUsi
HHeCHh48gofMFJOvCluk4Cq6xKMvUuU2n5qg+JI1aiFsldnmJlpRaCCCDadWVYso
fyaSwDpoYJ6aND6ZhoFYF7Q/5phVMU5pOaKYQxc9QHsm3oqOyyvHouQsCG/LtpXu
0nF8rVoL61t5PfWEnpVwPOma9vQaNjy7+JFYXeb3FXtKJjEsZS6/nHQ4A4gpB0ZU
J4QgqCxpOKu3ZrK/n/Odg7oQ2jaEPwa9nQ3sJ4rN4wT4RYXbdbcYqikEc7Ys4FCf
FQKRQHRUjLUGGM1DAYcJCb7CfO17FiPwq6j64irY1549mVGbJ4q7XcoUJm+YcSb7
2V1Ugs/Ag7uQhd8HGPY7IBZRhT50WgRmwPBX+2iijLM0+gT8no/27UoFw+N1HwrK
G7spzSpswBaX4sAWvrcE+MQWydq+j/THP6EurjvvWksofSXVlJQiy77Ui3kmqG4L
FFgNwDBAmY9161ZrtShqZiqpminyPI/6+6ZfqLKEH3r/gpH6Nd9lE2lmy4ipQ/Op
fXs5u4MionJK6B5UoUgB4ChZoiFn1CRAimj04dzsPJ4R4F74Voh60wI0xqYt5T7N
3C5SxFEHvO67BqDEgBCOjOQ0QEQtc+Xlwh/sot8Zo8veupGQozIupOCN1CN1svlb
fEbhalHfKNGBdXtMy+F64iaE8qBrawW0KBxxvtkn38+oZHtSK6oqjaEHTZURIYjF
5eN/EFnD58KbJ13GQwtQ1+WNVRNrLYXs+Jja3jGwhWTF42aPmSBzD1ULdYi2jYcz
xJ33pZx3XfsDpNMoQlzRk3LFi5MUZyYE4x8qY/ZOTGxcTnuMJ14V/u6n403PIQo/
nTHNeUmosuFdAnJIOGOsz3VoTFnI7Th++h7gKSq1kZJ176Bw2oKb9/d5flHM14ep
DafPGajjX8koDPnk+UUJQPbqFItYwCLS6ydA+khNVes7bqv003vTXENHXWWn9RSR
1AfjefL0Jc2X/5m71g0Mvuvs7ZH16KXTXjKYyaItatZuGoJsRLMCgJywvejw4QP2
IdKSYNEmRzWz4GNKIU8k8i+Zl+nLj/9Hc2rS514vYeWgUjMPv5ZEczq4XuTkZg0X
dPPnZJxhm/1+YIqrhNA1WPlmrwQTj6V+XhVRA6FFgg6jHDwg9Cq5n8kGCF5+iyuX
DKbLvJSMLnH4f1vaLuZId+OdBrrQxYtmB7fNm/FpdECaWW3oMoDIl68RH0RsSUAQ
0JE9D2cgQkF511I7gB9/wwPz+PfeNVYZ/KTt0K6WmfCk2M2JF6AF/7KJZc9YztPk
xmqGetVg4D1vJjtk/n8wZgQ6bNp5IDIBUe1WWYrctJKWPJtTO1hXOQHwA0xvZmYD
2ydWdrAy/tFs331AzDfDslKZFS8sFy5xtdL6z7yA6BEnFtH6ZRajHlT985vlGH4I
YGN2B3HXpiGWby/5J9X7ayRoJfSLUyObTNzSPtEJxcIUbCBwrBOLKkNxw4QZG21B
R1ZXlDjW24WfdvCRA0bR84J8mR0UfYeOJPocOnTBubHWCEEPoiZ5t3cZ/c0/yvCs
ZFgqVldrytEHoW8mxNSSy8C4SQqeVlFQBP1mLhAkpD8vhDLN3UM3MBpndzAl3wp5
7s7r3z7FXPA4xn2Tw+nvkTUpYlPKL/pE2dGHXGET6LcYUNYagslySCjNuY8hBgI7
iQ/NvNiu5rQXbpJX9oxAHpHdp2VrH4qWddPAv/4mPYDFyPp4126jajahKpk6w96e
i1aU/oLNBOcx1w2S8a7SW2G6YWQWm7iM+CXAuSArJrBEAlekdCKdfX1tC7kQ7yBq
ztDMxV/Y+lQfquh/qpl+1qfGhQaNFM71HJeOdISmqG4g6tBJzf+iOd40u5aEpJRv
kSafyJh5/wi3pboVN8dYvmfkHLrjiJjjJAbeVUpVaHFG5LFD4WbI8r8yJj1jikh+
1h+lEc2N2DmrPLeHr1CLPFJ3eZSoZUbDawC1anflon4JkPK7HqKG2CVySPTTaLal
j81UwbhFrjBEMmLvjX2FLenry8vNW+SS46COJ12jxUotdrFDPpKhgqhhZqZKZNIF
XfzSEHufBxzJDQgdfXDldQJ71eNJQGBTkPccAGqFqTqn+Rjh87fnAt5CQe9FaUac
yxRNDKUhK8y43W0v5rc7pzXo42O6R8uAECG9N4OHjdE7gdjVdChMZXjVDnNHQ1/2
Jefszguus9xLnR8wwMNGnlP/DzjU5AiocOVOcUI2tDmqMmhRqxjmGFJlCz5t1CN0
YhR/qeC2amFmKHvmQKicK2JCrl8T/wNJR9svqiKXUuzVJB0IIQbwwaln5k1U3AgC
3ZL0HNZwIz4fMGZ60u4o3TBT/kuWqwLx3vqqibliSv/szlQ553QiBvKkWgvOpEwn
mMJrghsELNnxY7RJ3MFiBccF9IoCPLDEIuXnQ7HYO4EOwEjIPHZwY32qQUFrldav
C8bqaiRyWWmgY8cxD7pRIXb+opC9lzEAH5RjAmyK2ZKINfNKxFuKBMumzDazawJH
GF5cxopVD+qQlsbZXaxOnlE3K7uvFbg0kgAbjtqzr5dm5ZwPYiTDuUfj1VC3KRrb
kSspXjzmFgnjZkhC/hXiDAAwsjEyhzCB1f2bWefjsBAnnEsCB0yM4HOJY9Auc+R5
gXRw6xgG1SILDbVA/wHDGZ5+38IK9/rdwdH5pZriEQfpMideBMYN8SKb/8zL/sA5
gTZyFzBD+tamSnmbDvj7suTPjsAFut/OFF63L+3hLLVltiGSzQLiMJaJpIqkRbtO
RMZPpDuQHVVQdZr/2jdwSQIAjbO6NXCA2gCbL7bZCi7W+8BNc/2kaJrrOBKySq8T
b49xBh1EOglNa/juDcG8Jly+EFate3L66fBxhwnhuydfAaS92ysJruMNE9r0HEvi
LPqGl8MXxrfiPxQ1uwqBlvVxed4aTYel2dLtBXYG+LhHbEFSA/fX63u9QIOghDMv
E7hbVEEBl7kozaP7UUH1k6TlR5i5085VYpL4lG/3hjulEiuAVZLxy0SDjjGUqomp
wLc08eYSN5OH+ChKofpM2aPAo3NOYpvLaXsZUOW6LwK6CDJcK2Be5Ym3ZtkGuPjw
ROGqw+5MJX4joNSKbFvGxBTadT2Cw8QDNEwHAGl8gKgXk62tprSICQ3VCHr5deYc
tgl9KkKsNwnCrqaSk+lqoOojRPmf+DQ36aZkKPQUWDdIkxb19KmTiNyx7DJeWqXl
pagAxH1K5Sv7/iBa+ecZN9O2wMeJN/LGoFZDSeBijFHXQL5xsoiOQ5yzfgAqgLII
BYj3Kg0RZs//WUk+uITYwkMmEh0WrV/rRQMb+hoGSldHC1ueA7T8d6M1LDsQRyW2
hScmFLEBGgeebGwrdMMpnIxkoRdZ+dcb1QmngnFkM57zyIqK3EwvdgFKVEPDM6UE
7HUWStkwEssLAuUhdqhXHkPS/BYpjIZ4WHYhojdn4FlUuT9yvCtNPRR7z71Kk2P7
gob47O+/7ROWu2ih5ALeG53+jXK/W+cJUp8Dhj4OEmqkdqTXXj/dfhEKSRe3GETU
NaC6uxPEXx3lQTuCaYXIhWtCwSQrC0yEv7/XUNa7vnTuBqSog+tXeW3GOKYVX7Te
1BZO0OVZF6CygsD9gx5/TwXKhgNR7+R5NVLSczua59UilTzm+dVwUVhbSLtjGo0R
MyPYUeLKUprDeiByJGY/GucJWDCC9scAKSu6H5KXS58VLUvngMCD/Qs8OlsJ0ynu
RqsPyLa2Q2w4wWQ5jp506vh+OL4haE4JSydQCVlwQGyHvLXlLs9o971Oy9QZ5Imq
rK7zSbQhHWdLwZrCugq/98jRFWTK0RyQ1X5p3O+JUEd17etSS/LXT8cDzgP7D81W
DkqfpzMHgwAAgQ2W0XWc7CCTc6qfvSvYODLNNZyEoSAEm1b2POR6S9tr9i6M4wnR
3hh70HtXTH/1sdueMuE2jm8J+v2Uc8MFhOdOaYUb0+goHvAI09LnY4Dh+OKZRp32
tEpifTEq/I2Zla1OAceP8WSNFlrMU+zqV/zuD1GwZ8hy6sBF7b55Jah7ezgiglG8
YYc1YkKcOMSdtDneRdd1yJPjsnWLq8H+OCMwg/7V+DZxmqt52RGeiYtbCnb0++VC
XX3d0X8Y1gCA4gWNVik2lqKsK5XKL8KLrfDhAuhXQzW18gNKew2Xd+5RsOiHgrjw
h/QLNEBAr9pbJAt/TvRQQmA9Q78LOR9ZUXJ3YVz+KAi1csXTjhieViODJNOTe8XK
gVl0Ei8GVCpp0FMvZYYDGS101i3QtzLh5mhXWx78Sfic6LgM/58NuDPNBM5uBqA5
sXXx3T2wDY+xCbJVdMNJ5krg9k0o0hhcmEOvoG3OvBVqQPaKXgLW3Srhg0glWYBK
WK5bL4eD+XhRUaeuwt9cgPeBQ95jusyrtM6Zj2vX/Yfmo3N7GKnvcZ62JBnyfgZF
BWe8ZK4tLWBF109nIdfqBO6welGG5r7t9D4Mu0Nartr1PF1l575wLzyDHKUatSSS
WpeieZlpNRvbSeG5eD0bcOMIF88+DGrvuMbHg5I2cKaBhURBIR3brnWKdOmpLGyO
vSeB80BDedEzfqiZKP+sQv9q37oUQVxAu8PZB8vueu2TFv87unXl/LiPnRdSvROJ
MVVTGZ+Nvn0kWuj3vIi9KULxV4mKi8VFPx1iFFc7qTrE+98qKnCSHRnnWXK5JSoV
vnfQwh4HGsvrpHVsX/Pl1EEO+KUD6FpepiEcyA0j/pOIoCFJWNRrzsiQ1RSvrTdC
Ms/Oikf8t6szohCuXbfF9PHph5fjaGsW5g6S7kpR8I66qfWiPOzxNYDo18OxKxD4
5VpQ7EDrvTVvTx4pNFS9wtG622hbM9BmgrjuG666nRmmGmKwywS0B/JKt1Mbw7zW
/CGu76fpW964YZvCM1+TsUr2921n+ZONuPBPtDxFgROfzRyTSHFfaaB1iRhbUotN
CLCdIyXSbomOtPu33ZkkySDpY03JiIryW9IPylI29rrwP1EcWg5SMFM7cnfnlahl
OLT6xzIZn6B4t2XkoKICY9MVruzuqCof4nYsXXXQdpXpYst863DT6FeA7ITgkSqf
36wJG0RZpQjsddnKCFRr38mGT3en03+ENtxn26mPpxXQ2RoT7K/Cdev6uAlWUyy+
IfOpRn2zn3/wKkwn86V7Lp4Gd+NK0UPFwZMpqV+TCcrtpuN/M9tUBb3I3qHvPXYQ
L9E1gD7tzyjvW/xu23ZZaMHlixRJcdEfG5VFyBtv9yMUMTEb2BHCjxACxbvOiWHx
k3fJcHdEBCYq9dl09zDHYkltauH9i8ZuQQcg6MMWpd3kmsHDrp8KJ/LW7kn/KrBA
Y/ZRFaavn4z0OoGt1atu+LakIRjOfsXOycaLGF2ek39VaC5aCwSKna3b/wuOGk2e
n6baVBFFGNcK0w04a6W2nsh5xmPHqgjuk23EuU2SNGp2VFrHPLWWUnr9kHV8ed5g
rYDcOsgW3nNqpWXStjSMWQmGvR9Fb92GfbovlgvGENji4wkNBCKbICP1xoUECrbJ
q2cGdrwfbhWJIW6CNFWgMdzTMab7t0fKT2NnVgkic5lm+wSdfATjVBCdJAEqQVaK
U/ijeL5cOxcSc1yjCw+g4mC1+WFMjoAhRmuV4pBU8jF7Pf7ZQQZbC3KhR6d5djYh
WnjHUtdrsOMZMffSwGZkQh+10t0v3HD1UY4qBhkeEca3tqeUCXDQTXZUzZG81/nj
mNJOtrO9kK294PgRGW1fa4PFhShwW9gJc4SGKTXEmbR4mBfiWHkR5NOywlvjWbXE
oXXeHpcvHmuSZc7xOh44G8jRGKy58a5dCKoUMhb1gM/bp+rftbm91GqnXfN6L7lE
TnM2YhAgaIG815ZfjQe9vxmugUHGiVgZbtN2I0Ywj5ze4NuKC420uZG4Xyp2j7Y2
bfZ4o3iUR5DLVBj6+XCEQMQoeO8cvJhfj3tbC3kcsp7dgEBpeAS289FDA3y3DDMp
DiSflk0w91Dho52oA8eBVBraux/3tkfgyJZH4ox5YjEWfMdQ1g5aPKOHozrvgH8A
/BgZiXWjq/HZju2c/MtF7cWv5XmYa5QsF7rrsdSxZrmP7njGMZ3hxGKBL9Xuw9+O
7aT5cpnVNVb4160kWeRAzVbLkgEQGgS61pgmDjYAEF/zuTinpM5zaSy+mp5eSHYU
StonlJkBTEKsXXVOq50k5GPhNz2ICkscTpt7hvMkpB1Rl7F491Csf8f2TipWc/Ib
lJVaLogAMu5KCWNlWhyM7ceHSmrZR5o8D7ss5lDHmpGKG1d1Lf4LJHuuowcqIkDN
izzASjWVyPCkNdYe836BoSq/WVvTc7RCDgqiSn+izmOFmx9Pv4e1Jd+10TqyFkqp
UFci2hkBn6NrCR2TzTzjsXzHaSympuKk9Epe/gHhflyub5FOUgDXpeEcmK1ynkab
5rz5OVYodrNF+G36PvTWyNNAR6TTaEt8FNi+AWZ8FTihe53dsLhkVWbDPEpH0We8
5PmuP3+rZNTAnO6wpNk66ODzEKCq43SLkjTBWAZREPB3ZryIzMB3ItD/FHpWaBlb
Aq6yy6+Z87NTNuBgqqb5HKbXfxLzJdeqDtKifduTIORFgjWkJ+EnWI/cxVFD2HMK
OTufyjcf+rTWDvGQvxcelvy4IvXvQM209YUgPZOq0Z788A2DUs21ED2bunoCZlRa
0CSRqyta2p/ld7jVhaflxT6XM0OBx9SIfvDCcpHeXNHJcZqKhigT3OGZ3C/U7N40
YUayeNF1sFDDwKJpEUbFDqwQYjl2BXQZZTLep8KLOg3+n/TN/hsCELYgzKRdcg4j
p40Jjduh1QDGQzjd6fM2DFlco2xcFgUGMmbTa/rLv5I1Thww3fk4uUrR+8ZlxW/e
1tI42F9WRO4SOicxXoSM0Qm21JIH7s9B2dyYPwcEPLqi7WLlfLuFOHw3ZkzUhAxY
GlGyCU6te6bSWnasyjXx7zfHjWo+qLYTuRZzrFQiNmkQuwhyWZxFV35rr7na3QLR
sqcCv5zRJjmJ4oXcPPgJYiTmlHc8ho00MMxYQKoa0GzZzH6PXw6zMFelPDZnl5wT
HEWkWu1HUdcUn32Z6lX9mxhpK8fKsq5AbdqnpThDAoy/ZY49tJaAU6ZCG2YRIglk
YlrjE8Edr1PezOAyJ9sCvRObi83iN2zcrMpJDsCecl2Ged5j8GYLFMMrUJRY2jXL
WBku+pnZ/1THFQ3vWoyEuB2qASCu3fYiK4uNjPyNwb0Hr82BqrV1zB/CBNFpzgLl
nVZg+goWl7+ul3QyaK+mJy++vPZz6MF8+Ir9TJqUbUYSzBeODTws5wR2suUaprLX
Fp/GVqq2KBNyCFt/ga1W6dVZw0FHC1nVKQWRMOIE4zunQhBJxpTdKm5PFG0DBHpj
8YWExlW7+w/bjpGhOVyeV7PpEEfwz2Csh2qmIgqV6UGplfob45xBT47oqxx2wNRs
rUPL+gJwiJEz1YgiATnC2bBaALvtJBEBZGD3AVK9yfRQ9/Cqri7NruF9T9Q7NMtq
qc4tcOAqMUxCb2bFQCII6MqY/0bYcApBO44P5sSFFMyfwKjuO/LMJjPJYDsw7tFF
+COd+CM0DzHrpQIIHGcrZGApT5aZm51s5WSbPffpOEW2nF+l9ZOA9C4Xn6ZtHuPH
rIF/Kq0ObgM2vs4ZDGx7Gmdr4G9zu/oZZjfv3sxqEKNABtWPU/vOQXiaYX0lVT2S
UWNaNyozNCeOyvwgNPtChUUToAUB4WLqmRpws68uJ0tpGEPCxWA0dnIzlXClQkW4
5wKugMLlL/pWgi5O0BEnl5C/mqUYe/7wbyhw9abP3NhEvrR/J86EHYHGGtHfx0XL
b0dGVDnIS0l3aKL2RtRjnaa79QB7tXj6ED5RImePbhAsihLyQjPcvVpLqZAevp2H
Jt+b7cF62K1aj8rfglTLfxQU6H3e31FdvJtqbFjagnysVEDra9LSv3mr0RmY27o4
bOVXJQlqcyhKUpJ4fwCPnaoFlxbAQ0d3Fbx+L97m9l3w4FKfAnXxPas4p4X3y41H
U+yJnPjGR0McZk/qQhZKPP9EYSN/U/5BIEtkTcEESmQXLXjNal8ZjSt7bryHQx2G
4EdnK+QH3cQKnh9stn7CHOXz/feanqZ8CBOHoKgLVscGsT+Q/TO/4zQr7KHaEkhk
UMW0xk8Iyl65nGScGnIDt9coahJ9q1Ag9bCj2tJY0TilG70hpGYopqIqzBBGT2FP
mdMvrfdgGuY1nDIbjWOLmKXWfIKwiFIczXyxBWW4lcLw0FQ1rc35OWIEMKMwZeXO
+mLum6t0IT0eltHAgVzyn+8wMjKuyi5E/8y1URlqkdGlG+hCA83y/pgvETuJylwR
BXGpWFRX+Kl6i/BSHN+HaDzcY8mhRuXNouQtRgsR2xxteuAx5aKvUYe+X/2tmz8y
zxCw+BuB2clQFICeTLjS3aajg2jJPOQCtLpFWMPVUNU4BkS09n0h8ac+ROoe19IM
JVyi0lsq3aAJKWJUx0JlrYBoMasUsnX25GZG8Z1c+GAHdQ0JH+ENpVCEYxjemczN
1zPyvt7ApAuuFXAgXfFFo2x3Q0w23eRThc9Z57RRFqSx/ENmO153j5k5v7pSb1SQ
pfFly3FTQjIEMOohLf9xu9Z/Cf7OfxwU1N+62u+EiLIlAssgtusMLeFCQQ29VDpp
b6KTPSNgTZggQA1jPCd7zqOjHW2vm7FCAH3dcQDDOg6fP+62w0+6GFHWIF9B+0Y+
su2r+fy2ytvJQbIiOkNbN4ZFbkWtR6lrbZzWfnrGhm8ShD2YYEBloRG/kN6wVW+G
bdlw1na+JnqdDR8WBPT4CJLAnLkSWMljuocWR4SiMFuE5IKlL5aPek5t7eP1BL5H
kkXjE/+HaPTBzeCMEuRoHUzWUdDDqH4KG/aaiubIjL5Y37Gk//0aqsa3BpqkXVtA
Te/BWPYaYtNAghXapo72HBFrDOlUV94+zGoc/VqBAIAiO8ymlzllaOdI9Ld9reHn
rTmvT5LvEzxovjxWUDzhEk4BozxDRKo9mrqsRgsonJ5hRi+rbQVk5N+3sHjJuw+t
RUGn3/d8G4n+4Wa0+0rnQgqsfPByK/DT3BrFwVum+woPORjINI7Z06H6YrwSaZzn
JfS3hwAygxpEAgAk5JXQbruUX2IRsVWI5FJm/3GO+YxvIwsdAubFrDmf1oqbdlb+
tBEp2HhF7ESswW7DxbQeMoEpmaK6JIayui2xOK7ymtH4DYzNfW00NomMPu/o6JLR
Nblp6dpgB2lp1dDa80PWuE08Xu53O2YAOfDptFhgxlHEHn/Bc/QKp0ltX4agv1Fj
uelf+zD87gEy0ZvIH+uI6GiAWpjQhgg0ligqOEaZGXe7sWR+NTtF2YoOyZaWyQ1i
zNvQJDSVTx0jD96JBIZykLJHxcTPDYb3i3vMp1DVA3z2JaYV3OV5uIyK8qbHIpJj
a0/B89cRJSTtuz+r4DK80G4JZiwZLFXZJJQK60jDjWT79uJQ6ee0edc/dnhzK3vB
ZKzo7qGjieozj7odxaljhmC58DA4vYyk7mb991hUrXNlq++5M7UUWWiaNGh8HRDO
RTqs4pm/qticvRevy+JR0kHQeQfasHZA9AK8TpR7LLsTvHccOjEABHEONySNIYcL
L7VhjQwpKh9jKMa/cdgPEdIRIbR6JugmDn5dACnXfd1xRYByYKopWkNHAwAE2O3A
37PSzp+hyK+Sj6ghxQrbKafXJos7IcrahtK8DJRmOJ6w1ZVeO9z7lXi2jKKgwG60
N9gBnPg18JP2HcQ8FGnixmvoK3+jgghnrsQ2AwijArHYYnitj+6u9iBHNqG7dK2X
PRX3OijoqI7ZtCGBqBc9uZSChiWxe2wm8JsZr1fzPh/gR+jOsQ/Fk0zyhhSRUlls
UZ1FAPC3rjbDt3svL6h17r71STW5UHXaMmfFpVrZOSN2b4Rfe+MPw523tjx0c39N
16g0liWriGHC7Ajb2H0RQqlTlPquoJ32Rz0VblqvpXZmL5f9y+wUzIEbcXOP2866
fJmkBD9rdXXVSIkYfgbJhSpIHgB8pj1f0UgLFi4mgHXpOMxzX7Dukjah4mYQgidZ
RWDsvE9fhOfjhUA7fyWPAuJXwKALBcGD80kxqzRxAloVEapO/lyW3/ZwnJhH8gla
aUxa8zDDoc1idX8Djx/OVww34h+89INViTX/v6FBdbzKZlTM9psYxyEQ41IAihvh
DogdWObrBeKrXHd/eU0tU+hsqNg5uFtH7yB6MKbMPQIdahJbwH4+gLhA64oUT0V0
2fIgypLoYpk4v925E6rD7Oa9teI0zNSVmCDQzb0iREsEsDw0a/ZhiMZFoAS4h5xz
e4TUJESZmQO+SdOj46TsNyimTXuUki5uymBXgyYUA/49qafw18yFhVnsdAxBL2fW
UkQ2ADM0Bd9tb6lKNYkhNt7ZAnarKU8vQvHFG3W+wNMZZ75aI7MADifKI7uTYHEL
q3Q/g/OzsLM41DJjeol3JJwbpM1GUUTu0jp4sogjcJdpzFCIPazUV8B7MHcGvSaU
VmZ3G73JPEzqjQmwq+EBSjXAp6pUBmIWDFpXaJrRuHJeL9kI9vXGGKLor1FS10vX
rlxd/ruk7IfHrZKY3k5FcNEcyahWyZtJ8iBxL0ieoRlTXTFamrmoV7lFHWrs2q8w
Za8YyWK4hsFhazmAFtXga0DjunjIERMh+5XhnB78l3whwONW7HZ+Jjr80kvdfHLW
4JnKeJOxoSZVlpRVivUB/zYs2e0SZ0xnrmO/D2o0Febj/eE/o7wR8hcpL5tlI3aq
VV3HuSzIRU/UiGkxgIzFjsb2tspmvsAaJWW9cR/Z89oRai8v+pINAbFXpIO2Z8Jf
R/NKFJc3dQ3YCGT8+yFIwKq8OHsX65+Lhq2y7xOhf0gNddZCfpVPgySaWxD8e8oL
nO7GTO6DVW/+28I+SUSmpXpjwZnAK29Soo+Y5bkirPZCqRyU5cp+B9yxcHJaz6tA
LZMJ4CWqOukufQERTVk2auqO96JTRWGtxOQKEFp9gGr1eyhDSGFUfVwcmAOenrxW
IfffK00pzNrnY0EEf+4lOu/1rubn/PzHpCM482MJ1Cn4XrKygvF+ETT7/AGik+wW
iVuaA/H2jT7DkL4U5f0ca2EdnoUICS9SETvOMtwTquT8sfSzSDptpgokDcR38LeN
jOsU0sSCFlewTVYT65r2O8fZCu8XOjhFMkpPka5uLLelhwWqK0ipGlGnpHbDhtBH
jgPMTpM1eyIoysLTsbTdtKZKz7BNBV3KicaGCD6YMzq7hCC/RflvF/z4gOqhGX9I
/nfDLKMkt2X85nMkOVrB3MWHnfkJVfIXCZ8elLq62MrpJxfsJ717shcc8N9wYHLP
iKYYU2in8W1RDxWjmSosW9kNXuIMPLxQj6xWwlTETygWGMAFJzArsJC44cRvhLh7
BcC1hkRFUSVkikFGHMKm+P0KsP9zktiII3/dvdV9+W/xVKMwU+TydB54jPsvJW97
dIT6AMgsyheboYijRJbCqWP5sZPGJP4hsVdkuniUMbGQ9hSTFf0iJown7MNYJi/g
XgKcmPZTZn5yXdG+d3i9gGcyPJc5Til1aPfNCwvHcbg+f7Au+tDBWtbsae+NzW/9
EoNXgZvE5K2Wsy1rhsheSquwDvnTJoTxuUwDW8V1H3EF97LWYuyp/XO7upbgbT55
Y/BZQNqYkp/WlS1Qja4D28++1MAhIrNq/s8ccIAz/ZmtqIw3cDXyE0fvqecGNJPD
vXDaREZWo4Oh0TOq1o5awFzaEyZLo9xXPtP6ztXzqK/llDPOCGP0YH+Oh5CEM64o
TYn3HqjR/fxw2Jk/HSBYWfGtsMtQryFyO8av6pTDWMg59GuCOQ8tsaPVqXqHN/bd
rKoBT1uGZdi9l8W2oARa+sfT0lJhXdxccoyuULZRxFPpiYUfuUDtEGSZJ+YtBSa9
7lua3ue1pOrM54RxE3H6t6BJfvlicpNT6sQCK4xIXbehL4VdBD73Rc4O2/QXmN5O
pMxT5WhPuR2onFLoshcRvNgD9I2u28jTwSNBCKkMJYEejqpIco6KRhlLkauLnMza
7KeKZlMEbU1gkcyb0CvvM2JrCJVkyhVCzEkCAoDFcLlefIVuevtjyJKz9Szqvs8o
fxsH5NR7QpLNK1+6wRlu1Ad8lcFP3iLqxER4i3r1cwu2D5uU3Geg+/d1gZKk/Lk0
IeXZviTQKMwKb8wKsC/PgXUBYXeqFrFg6ORVJtRAWDg8HP7fGFBQMuqViEiZ66D0
sN2TERvsXA2eqwIDIxDrFGQM3f0lJwcEDQ4XSXDntN6Tk7OIbkmqfopzzK0779eQ
5BhTMGoa+4Jn7TD7yEB/Mjv6F0AJ7FWPkdQHZjnfE5zdD2nDHHrBzJmF8j+9cR7f
mv7XtKl8T72Y4KYxEEgldVR2AssfFn8IF2x3S97a5iT0XVMHh0afP25PlGlyCCti
+ovJHQ8aDjfKaPgXPnHDlBej9LA/Gj9fisjyfgxNyVQ8e15bkbAcCaEHz+cpCojg
nIltxS9jrBFm2DFLzjYHPRqVBCDyNinNgKIzoio+yCB4+6jDwIVIfxcbtsYDVyVj
pNVEucTUuv9cCjbXWDr9RTk4OpAwxpYvx9WZ/rZtS1my1xOilW6ALphBVXflCcDR
+rGSTYZjLmL5lhGcCosy4NDd8LFpYKs7B03qlm8LpZw/ZY75DwINbQVFzv2pr2G/
uha4nLjUaECu/lQ9Mp/zmbOKv4JrUJ1ts2ZGwyATM0+AAzYU0qmItUXjxlfpHUZy
rfiKwDriHBdC+7AfU9lztiPOAHkqUtu+prGfnoYrd3pT9rbjk02ZLH6IPVlBjwcc
x3VUumh6hgT8QvBaaDTjR56pHmIwe2Cp29PjJjwkXjgXwrQ1iUemhAJZVGDayKhi
zORe7VEe5qhurphvWNAgN7QwRWGXheHXUN8UHVphx/teyRABHFGZ/gsWy1sE0xX4
O5t0pZWV7cCXrDmJboj/LuQ5jS+EtsCygVNcScI/ZzEAcTH7x5eHDDPS7BA0el74
wJytYpNDW8xw8lBWCXOcf5+X9XWOPVA9gCvHF75Bwy+rfkvwz202Tv4lG1pdBSGk
+sIQR2Ga1gKy1BGn+MSS2ctjXkQ45tEtsoQIhMmOeJwfR6zazMoAuA87EcskqgDX
OAjKLCLXZ9fkC9BhUKJb26qK+XAFZfpwbqH2EQEp7VfyGjiwyITZfAGDGOidjgVe
xtU0evtJHIxFLD+ur6hNH7LjN7et6wMTT2BAqqirV/+ZwhtNLu1UrsKM/5JsUhnR
HPKZrABzWxMP6hzXdKojh0138unYUN5dbkVRax2E0dXrIR4tVZjI+rE1pfsP3kYF
aL93W9KjzIeHtI8fSLuGyhIz/GtSCnYLmiL38GSfWDHUUIt4ZsQh/O8nXTeVunT9
IfxCEbNV0lUuEy9zW5p87AZjFbJO4Mx73ppNxNbYX3aETRenw4C7NaStcoRNiMuC
gNp8bzwZBCNA6DNaC6aITO9vha2trO1IHshPq2PnfgLnp1FVxIv87VbE7vO3sfwV
feFHQvuxZdX+AFFvmqnZfMZjQtBCC9bTNW1jWeYv1Imt1KftbFeqEy/n+BwC9ujA
pGs4yg88jgNu1alCJFYSSIJ7Lw4USh8BdXlXtY1jM7P8o1+uygUca+PeHFNZ+YLq
HgdU3bzaSFEbdAXJuXdtV7hzZevGo8KlPQ3vIvstBwii8WkSTyQ/nQaX0Kz8wIf9
UGdA/noNOwv8yeMuUPqR3GRMswFNba8dXwr1vhzho/3rfdKtjtIQZ7MnpodEvRlg
2zf4QkrsHDwvAfWknomzVkbqmeAP/6iAodEeTp6AXwT4tbybKKQy+omeMsY4dpGk
MoN8cgnaD+aD8ZwbgJCyF8puzaHPTgpGDzaJ4d5z+Oo0dDlCmIeElF64b8UMAjuO
F0FYfdK09bVufP/OO9npI2lju9QlRvElqp5/sN46QQJNgfL8PvNBfb6nIhTSJg/j
Z+PWB80iFoLPI4ue1XZcpNvn57T3A9EZumPrH72Fe9Rt+tdS2PjNas8MOl0Jkho3
jMtU9bANY9mT5yJS/PDryU4RidfkvrIbS+yMq2TMDPwyiS9tneq56hzHGQV4Vi2O
Pb8s35BLdFQZHQRMvOhS2Y+OpuN4SqA+e6dy4L+UduYHh5Bkkj7nKAea3OBKk24L
h3noRH80EfBP/DFiWY8sHjmL0LJUtop37Rjr0oAN34aL2ep97gCr69BsUV58S9jt
dMUhqRs8ClHOCluxwL2DFUPQGbypG9wRJaKfLSPSev9/RDnEUK3/70A4sZgeP1X6
xxJaUOiSMPxxMn8yP/bR7AvTPFCvOuNzHdXQU/71MCJELhKOLVazl8Yb8Pzf9Hia
w6C2tamGGnchLGweRS/MEWQTY83GmYa2SxC5bdspipIKbvjLf4JyjxYvMF9rVdiE
pPH3Ngd8KSgJ6QCtJzDM1f+F/AEx7G8ItZjG2v2BkEgmMUbcqyzngkjVSuc+5YT+
Yycn+n11yjzsrIY2/Iy4c7PzH+fBVs33JJVYmVnBO5hPyjZ5NgNldvjLMtQ56w6/
kyDtr/NJsOS9I66HMIpdJjVOfgk+5d1xppfhEkcxrv5KzD025ZaBeMPcu7+7dH6J
HbPv0Rta6R+58vinGJhWPDp/UBpkxLK6mV483awrRAgeVdBwPkhe8pchBj5l/lkY
qvt7ihC1dmONNJWm6ZwCNYAX5dVuvaW5y52WXFLRzUM0XEEftDjf1VvSuLDnursh
qSp+pGYaELIftWYp53H3ciLubAoh5imi35pMBCqxK12WBG1QQemUaU8aZuRUk51/
x6C2Y/hLS9VsHT3GB0nRNBAmGLwcKT4jFpMSSG3Dhhl7YjnW2YSgUycrt8c9LsvE
m+cv4wdZhDhnlFBqhS570Foosz2EEsxdOVl5r5aeGOOc/Cx6a0yGx8dOTZdxcWUC
n3M5OJ20oQbTE2Xj2EGMH6qhPBU3sLgEE/mTUbSjCxpcC+CnGceGW+88YN/6E8fA
yIIfFGDUzQ92XBTgaHQN94okMwAW1HN+wf582BMumLrVBxPcQnghVw05lNiSTnvz
17XAYfaNDtHEV2tZhq4H9hdaP9mKPVppLm6do5hg9gdZLBr7G9pXzN5W5yuBIgNc
zqSaF2yEm1MsOzIdaNIyRgXyhBCsxacavd1CsN1ahKPehFTs3kovxhfgdmddvLSb
iFCMIhhrIxzPiY8bHX2hT6h2Rnr7f78hQ05K6D1fgd6UXerKnm7txemlEQmzNGPc
KhMHr1uV/TqCOoGSx9w4IliWJxGyvBpKVNgnCA/0MEZhV1v24jLJt53tXEnLJKrx
Zg/u9YNKs1ITEYJ7rz76CuzCkua7uTXB78yxp+pnI/jyUCCv6vmUYDfYFh7dyuTp
SSniMeKP4HuO3/iPhIizXo9gsZvW65okEs/tooaYwXCwzQgpv7xNq5FJBAYqe+aC
0gGXkBJKL1gfD6wYNT09LUd+9V/eURqZIAvPyDW2+wv0teP6jCYUp7TLfwf8LLhH
GDm7zPDnQV32cb8fsZF97d/nECZGXLfOyrUfmykO6brxnEpyfNCTM6yNKNr54Tic
ioJmox9mPyyWPReW3x6/f9P9weW8d7xzi7lGm3i4o4MVKxsKRxd551Us0YXdcH3N
vlvDpYE8Uosh48SjlUAWCxHF12Cj/5kL+QC3WwE/pwJGusW/3dYB6u3K0bwUR4Fh
1lEBp4pKwJJUt9XXS5IQnfsP06Jc+AmAASf7v24LJcryCT0dsyiueRbdio1/unY+
NJe/m6XE6h/nvswZTHQEFuNjon/arugRLo9bKSxXHJSMJm/0zG/3q6oui9XgILhs
omlGqlLUVOhyFdW6hy7SvO7g23wp1xUNOSLl+AJQcyU5brni5NOoEFrExWu7xTp5
bB7v1k2AbxQvtk1aklSJq1joEs6sTHbxagryoCP/AMkmPujwfCpSl0HiH3oCiOEa
8tmuURhNOQCd3kYOp7ao28vKhcApP/P2YcYnscvkWj95Tf3qs/5oTg1lAECtf0nG
w6hmECbpEce8oFVLLdLtttCPPeGSabrq4FCv5eRsKyn1X/fSqJebYRVCoz6Cmaiu
hT+QZfOLMqcn9m0ztKTuMoPEWjaOwOJWZAbaS+wpiJ0YmrCxO5yrSQCGdhXPodr9
7SHBk2MbDcKuVqpR/SWFraSc6h1Cr1mh40Uj7XTHxtr24f/MYPFBmaPp/YtzazEl
f0oCOt0+fBiF9kynNya7YhzR1ExaEA+Zb31Hd/Ztqc+GnFqWKP+ZpOFnJ6TYPIP0
IaSps/WkP+Amwv2xeSfOu+y1bd8jN+MR/QHKIaB4lG96Syn855y0aoNIsTClsnUQ
pEOJVjUR6GAeCMoUqoxl4ce5HTxSE7fRuoGfJZxbWXYiaLSunV191UVdq/pYno7k
1dNhzC2JF2g/GJwNAvIt73kqm0gBgi7yNO7D5ILB5JdpiubxiGhRdpxsNljmwvoj
fMa/UwHq3wGjFvnbMp6SWi3u5ZIzTOFySkPnY/5qYDLf0IvCakYB8I4QX7GGL9hr
QtW3GUkGiuat7XzketDWuiPegIrHse/yJR6ExKAnJmPpKdZDgz2F8C704P2F8BAe
MHJ82FXPfsouM9Mm4Db8TzaDpblzILpah+50emraTm9Ix4Xhy7qHYIBp95YBv5NN
voMi5SY7PwKPCPoXs0MHzQCxuqfwDX8HEFqBSn8dr5TjJD13CjC1bYZp1Mc13OmH
OJfjcTB0yjT1dzFwfnUQfonOVyQMM9HFnUPw9gsnS9DHYCABoTSbp/gT9hBXDa7x
hcBm9L5WUHpn6oLi2vnnR582L/Jhw7xxpw3RGwzVpaYiCIVIdaUAHkD3QMaHn6We
6ppWlFt3Ct/LVNQJdQ+B1/HpY3xQzzrI1m6qWQoBMhjYSWEB67DMZAOQTAbACblR
Hy/woEQ5v7mcPBrc3dG/Id/t2Hc7yAB1lZ3cP8nLOv2dnXU7AWJFEKPRp9droGIS
IzzMFbmVVsVKKN6xFu+FSoZYNjnPqf5hJ8edGdSqcCSlb9Qi/4spK1jjJxRXEAYa
Fk94PM28xv6D0TZi/qf18qwOP1N9wDUU493pkhKV5RHc5J072Os+dkR9aUTwUd3o
7rYfniJO8s6hEwdh+Y9a+IFmw245LiR3qVfSCCMlY9ieEn5FDsLmM1FyHBUGLelN
hViv52PqrbYzZUGkswV7Nc2dbvHrn7JyYx2PN3XlqdsGlcdIiRrkb3ZSKuvWHcZL
WIwSSddwpltKlvbDlqlW89ofZFW9BZn4tfZzVwpVOKnj51lxkZsE8x/aDwc+Ua9t
lMfT7AL2JtXG/p8PyBQ0Aky6c08xTYwGULidc4aQPifvExXb4qvArgtSlysDsm9H
EFSdNNyN35/4es0o5bhHjtCjpKa9nbzhQEI+N6yC026IBi+VtaGtDzRbu+S5i4pp
IpsbpEJc0GVRo/2Ll0XkkdhbvCrvt0UJ2TAXYvUyAbNG+8Uk+1LiBmxUTHUF+x+q
u/ilcshmx+W59Kx3Ga/kIl+Z79sId0uFtZLNm+5vynnTmL1XkwjlIuq44utgqYA3
jH80LKNobGJt5n3baGZJ7lB3AGXtnvOGkIxSpF0Xj+AKG/b28TPgi70pr4PbPwm3
psJzMpIkbN8PJYz93I5TXRsIAd1fAv3zFPsICbFUnUQb5OTqE6lWJvsTuO8lteTp
O5QNMpum9f8K1vC+d6+/PT51ghLdpi0QGjA3O6p8jAE+brHixf7cUvKuJiOMu6nr
WAoyB6TJi9oLpBaq3GIo2NUOv4mUxmlgrGKiM3vTbX5eLJYAiCzRRHrU2dI48Mws
+qVDKes0ABJTOO9ryT3exrxaKAwEnc1/QupXnajTSTT0WhK0zE93WD0NRDYvNrx2
Vc0+0aew6vyh1qSkds8iCepTnsmiXPmxNT89SjjtQgOZM0DHxPt7Km/n3c9iIRX9
Q2KqQOMI/P09mUqfcK+7WcQVdPFMJr8pgRI1wjKA3HRyDrk0MikhE/uZSqKNvcTz
A18xAtJVUyQgzJHKwi1242CZ7jqZCMGz05Nxj2rM93mwRq6TpdQaP4U0VutQnCgZ
aE03L720nhxPKFWaUc6LC9TpnJATDndffWZq/HQjU89exzUPKw9eG/iBuTrYtFuz
kry2Dqc5p77NG0PES8w0Yf26XT4W7Ac9ImnQfMgYJVkw9Uep48RlcZ5CUimAsI98
cM/Swmcz+KxenCBTY7s1WHAyPecZA/BBEfinHCe4wEqEu140JB2CVaTaMoXwRKeC
cXcOpqHOv2N503pSsuh3qqdzGaPnO5nawupiDOrVrWXOKCQtzKj5saisOds3R0fp
HOTkq7UzyUG0BrN0jniekmdJR1CmXr2EM1rrBnFQzAgrZqc5XkwOQoxYwhs/ye86
v4XoOIdFd3J3fUpg57PWwxD9noJIBovvD149hncDxRq7zAPGfXkliB8mfY3Oq+7V
8DzgD6OIIJnePgK1ev+w30kwYPxVhVv1HopbBV9gEwr4tSyO0chtqTFE8pfNIyhe
401+aInqG63OVGSc/sDcbo8Gjlqq81pDUEwfyDyhEAHIT6p5T8Dyj0ixg5aAjLHN
aMtQZC9WpKUmIibho9GMlIE9tAQbO0sQH+WI+jPR7HcANpPs/gMma+WoFYJA7hWK
SxaF7rZf/0IKVUmiPYNReZqz4oRlv1sWW/YcHWmsEgLWhxZvkB/VFjcJPwuJ9n+S
qXhAuQDQGAa3avZlRW8hwgdIj31G0vOkaVTaTu3a4V0JpZi3czYiOEeYhPEhBjnL
yHUnC+yKBi5vNeQlR+H5j1zDi68aQH3sx4WrPh27VmSLm3JittQH4g6dhWHgvalE
3m7fH5II090O+Rx8M0PF3Ym7AxVNqsI38o6H5IuNP5YaciVWkO532d7BBTMCPZFz
qbRHfnptLlFFi7LnAowqmPO+egypdaLEa0cm3x6WRDCA4/DIBc0s57si4gLavCYs
ox4ymfCyEMLkzCTTIIAC+dOli2JY/ggQiblPCwvY/RLxXqKpsl/yAVLtlYHUSLHt
LisbK6a9yDgozAxEUPMjZJHSlSznoFgh//TdJLMukUWieaeI+BaliROU1IXLQAIc
Qismof0jNU4dIwoSzmf5DsC70E/7cFOZYlzR7ZtkYidml7K3wcjn14b6/EiQPKC6
3UZSZ+pmvCfz7lednLeyJfHqTU8OI8gIssbjWagHT95rIrPbiZFFk9L+ZRhM+EVy
geqgVP7PnwngjpM39mJ4q817wtt0LtzMSeE9wQWxG2mE7pfsLootFLvIvGuUG4PK
Xm4KFcClZor8QT0lR2enix4LzihIJmDr3k011rU6exnEU9ezT1btrRq0UiSaKSpa
gPYLNs7cl3PH0VDuuwht1EXJyop3kKA8/aaLh+D0KXivBdUlAv5GfjVSTVv0YYQ8
LvOMyCm/5sXJ8pc4KNFLRCsm3ngDcIyDdfSsBeG2cYk0CngE7DrY+ZEmdXcE6sTc
22FYdQt6k69XSjzL9WL2a74/VLqnKZWwBUNAcdt7kifx0jbJ7BENbUBGGjy8uFct
wsZT2UDSFn5fNgK+1XYtRrvar21/SChNtm8XFVJwqhXQdkRMtnVU5G7XI3cthAno
NE5hfHjJyzQOZEjpfmzCtfeOqXwSXtMpSKSbSbYSXGu57N+prj6L09Wg8gToeATC
nAEAxPxYOJhG4Qbj2UMpibJBS05917BHioJqqAT8g/YhNYpUnPvFg+6cmYMxH5ZY
CA8vri80cyqr+Xw8khR2X9ktJEmCwnupxQyld1idZvY9ctl+zEOH6dPESapMN1rc
v8A0RMn2aYK+Lmnw65caZXhPtUUr1NcHgHFedO5wwkd5/BwqBukYuu1OmQGG4/ie
YmtfJpXasenQtsA7AoxgzHqTfblcdGGIJ3KgCIaeY6wms45vSEtw5AMQNm5SB1Xw
YLrmF+B6/hX1ESFkT8GLpaDJNjVRlCRgmr0lNoG9JsqzJ9CyMF3/ca5DqfWaszGW
LSqzHZIxSqhGoOZ+xQ+5Cng44byyKJ/X0PY61X/lI0AQHNwx1rzJF4PFKw1eUcuk
HOHTLRrpAvssTwSVeOevVmzYpyxqPQROh5mFehwUeQPd3ND+8WZKxqKB3RzyAfob
F8DOUKimcFhMD5UznRyT+/+wE7rITTiJfJKnY0kOUGZo2soX3yOcflL2LwWkluh/
RdXVMEMOLzCMHNxxU22uN9u0ju1pP38IiE565k/Z5VUQKcRBOoclwaH8X81mtRG1
9SBgN19EQipyXjgxh0cIAloWl/sKZVnbjZ/oaKI+w+GP437pcp3SwksKobl0W4AI
K2cHNFS/E78QvU6d95EyP03IArb/IKef7WydRoYK3FfMXkdiLgIHtE3A6MlkrIvt
65KGdeYePV0hS9sAHyuHLt7Gq1Payw7qc27XNyQ52lvXrb8ASiBE2bTTlZ6gC6cA
1qsaVbH4m21ipWYFeZ8rh+GvLvzucdjzOXsI7ICl3355zq/wMPftIp8TjEOa8Wiq
r4lJLsjCSex+dfUjpi8qC3ZzA4gtBeg1WA64W5SjoQvh0Stu3m3Q4Z2VlLuybVEx
nXGWLKKFLGsmHoFi6eTrGx9zkUqs6W93XP+TOF/gnq4fmnFPAT7WVTijBm8XG9u7
4KUpu6ag7lrN4EKXmTOSaY6t8HO4Gk/yKpgLXo5zh3BJX0qK3V/pXJ+63h8gz7E0
6Sft0hohr7hGNx0s/hcRfNkr9oV7SbdSxHE0lz+MyXDSMN6sMdVIBUPUHeYo3Eq3
t8CvHQvaFtSuL4SRR0yK8mevpbpUtY0TmSbRDVrXM60ZtcruTBAxaPUd9ZqZxAKz
Wju/VEH2b0hWq9jpjOV8MiO4rIJD3pQa0GBwUlVN/sb+u7sPwDqSJ4BGQ5QZ1IVN
IJQUkrv8SoUvEjzqBwbDcFA9eCn+pan40l6IwSFQCuBr40F4bdbl7jieT6jVSZ3d
Xs81JNFIeO6tskBEHmqHDDlV7t7sJNxxQc2Df+KDKSZ4dSRtHmpnGApU4QzC93LF
TSVKQpgRyXnPh7bMomDG2PG+NglT2sl27tA86qFr7B3pvdpf82/O5SySd3tCqXH9
AG/bTrJ2OjOUTf6XtINgTnbPxWpo0fExCMXxywoU5EjLANAtGt2DpH3N0XSLN/zs
c8QvIyiNZJ3LhljYFWja0KG+r+SmkewjyMPA880TZCF7X0uq/jbFuu+2cUw9BL96
O+9Gnv3auIqvh2f+a2hjaOrKqeUchIpMqycLZsKLeMoFvDt/aYJzoaiwTdtz21Hs
xmJGSN4DQDzxkxs+ANtL9vKNdkiUuqYJ2HyhiraoAWlwuNJxcHazTjrAnS9CLczO
4Az06MwYuUbEsboUKY8d5D9+NV3bVMLh9n+QqHSB6D+fJPrvJiqIsi4VtVXdOvB5
bvUSL9iRaqqx3EXiGVHE+HT/iHSZ1FYZKCw7ePWiSXVcUYnYtPN/bbkDASfEU9ed
fTz8VfAo8Mb7cWOrJoT3gFpWhUdR/ot96dDPVm5u80GZ+0H1bQLJ3gyEL45hJLbS
M6MjTjxgZG0rDELMAIrBM+D3nhbImUMEJzw4htv8OoPzAka2O+8tYxlOI6FM+OHY
3tUNkyia37vS6TetKF5SF396p+qC3TGJ6VMRgQORI1wgcdlWzcaftUNP/vzft7mn
cp71tn9FJeb6m7fYCxV3LSot37J0+S4ligm058C2oOSUV4X1cGU80SLA+yz0+3qk
AigpfDyRViLnzE1xj4VkHxgZ5B7kLlu8KK0COZRw5/LpWLPt4zonMHvUV0PBY4TU
GtDuf7bY3yHGo9t9VDG02nDOFaC8ltOezE1+owQT7CkuoYyCPS0syU4xHcu5R+W5
7iS5+/YPW1R1+IjFfvRgeBatc2ExepgM+UnJJ2VCF2E1eKjroCs9latl8gQbyTd+
tAD6XqrXgTKjywJcBPnU0phoVyvHWx6C8e65gSoqgZW9BhPLdFeLpFGEuYpc1h9w
FWZhAVRmdkMsS2wJ5M08NFPAjEHJk7K0Or9YSeGZgWYSOyGP1kqsgwMoSjkQubfX
IUQ/kYZgJpQ4e9UnAR7j304Ajn9MUaxV8r6rSy9fxEM4dmpBndUpewBLOyEE8D9O
K1bSRbvd56dfQrip6/f8Uq1jasVjF37EtrEcVemknAPnRs9669fVEY6zl+6JnHZ0
nI8txqY85gJbrYwG0oL6kVV9wG0ZbUNLdg69vJer3nQnhpSm4zs/WdwRtTD7qSRU
2yW92xTgAYbzTPIVU4bBNMFzGnLPwoRRzPuKT/ONjLvACy2YMunnmoBB+IrE0hLY
oZkB8Bp0RzgYmpKrqk2I3Umbf4C58k+fIFa4AD4r89iOMukL9g5N7MjsykRiofwH
eDRvqXs7iVCcJsZUYO7iTGonk5PPIDn4MPRz4CU2vQnhqJPmz2PJHyCfaJqbtFSy
kRqln3SzqqSW+ehFKAF3YZS7zfBbsYqC2PbIu9xOwPXgbWQRApP/pl2XUN80/9Ue
FJHOFCd1cVahuaHi+YWKwNtkaErjwaYqDHPJD5JJAfrxGoV/QMcZHkW8rz5Vc+kS
d8ehoX/DHanCUNyXitFy3dr8rBOR07G1di7un59h+MYRcOe4420Rrr45n8GzJRzX
h0LLqGOwqx6HsBPz4OxBPIzzDv88wHMzoeRrRrItnqpl5KVpQl64xU35KhDdOknR
KHQdQbbLAmlUpX+q6DPZJWIbtLCyiHyTAJkMwnHQo5yahlb1SEgksGwt+4/gGU4B
0DWsMfPnjyCE7/ODELIcI4a8cMR/BXmmo0JdfwpTyG15YWwlyHYNxkUu6869Gyis
Evw+ES87SCt7j/qqagx/+xUCsa4B5IxIj72iC8FDbJpM8ECFRKF/BGqATv7EOs7R
5m6xcBr4GSYD2/pHGngbLc1x8wdkPhz9DdL8dKJNZhAMvuxMTJRwTyjWeMY2Curm
beYYfQolmArNoXfV4ZGowH6pwfsWB19jBHUyyll1S0qYq81MZwUDWmHR6jnMja8z
cqo5s/cwgIsRJ+tkJX7ISIiTjQNexr9fH11xKCw2pnU0S/VTE+ABbnmXsOAjom19
ld3jFoDaR9y6zVbUbFhQlvVmGiy8hRsZJHuL9rHgQAFFeI56ZOhQHgUBrNmJEl+Z
gAeIMyqqmE0p+Yg+5igmlsIR2Qo58AOuOtYzVcl6o9eJU+ZRGpkVcmEngwPs0aOW
Gjnx15fpLw1Qx3szcU5r9haTIcJd13eNQB6b/wek/3edA4OEycPWIhcxnGnXp9IG
JoCqrtIJL/9sYrAAfLOWHOf0m1eDKR5ssJEzp6YCyl+evmmldsb/kHlB8al/SS+L
2G9li4NnTr5gg6+7FIVpgY/ECnM+s4icpIC5zyhoYanJ68+TinFG9VXbw5cyHGja
KaY4+3fvRG63ete0UTb0PJbZ578lIEd3twp7L9Wrzb7RDg6BnjUAsFUzRDW2Iwd8
Qo5C6rcsL+mgiayJb5aq7ZbNenb0Ww07CEgiyrltR1JCP6mY06EyyEbtt4+oDnFF
xJJ5JgtSU17oQiaLSaZstbli/bVfyD2Z6gkjfkkBX7AX/sETYnThIecnrYOtcF6f
BQrUuf7jSxXYky0FNEiO8UiylxMiNxbUskeGmkOMsa0ce2mG/GjLilDKD5b4XaRt
T5BnK9q7hAiIEkusOWtX0JII680/9AiHyYo6oJbuu0Zaoo/8rP8pX4m3c6fZI5rj
Tduj3yyV9K4F6nu+yTHXuXGiDCVA3IZFJep5K4wi5bkKV5aNo2kSIf0q887T01SJ
GlyzZ1NYGaXzX8EEnP6n1lbaKJQYs5Hi6saxNXvDCO/pFyJ+1g5v3vkB3v7R5Kau
M2+xOvj5UcDhDeGxKbr2T6b+jyoSo7MqxFcT3uFtx5rbI/9WiHMEiAOE8bQk5JMM
MUFt0O92E4iCear7OeHdKBpEBYgh3ShemCp/tiXb6RD/K2NNQ7Am7Yg8lVjYschJ
z1tSKE34+clGMreQw5FL866Mxg7tkeIpKEtZsQdpJpymBxpT9QNdlOOzOYvA0Gim
heoaQZctv/Ku37HqhUUo/t8JatzOneO7fBGowPdVxA1KCEY+BbCFPBkTZn3sQawz
wwMKmTpdOcHkXEZkiV0hs+JNvYugvjoS9c68jT4J1WlDHmNgH2Dthq1nnILfjS4E
b/4XHJO5MITlOf6SmM0ABjOCMhtP3zqk6QOyC0FpyVyLjVWldZen/DZ5ASg5hKAA
7xMB9c5LYKEzpbX7srRsaFZgpG19raTlLia8a8kq2aRNy7F7ky30LTiQR5Za0oDa
3l+2YHrsai9VVR6p8Gz8FxgzUKxXth/t7fOzzkfig/qeZjg38+g6M4kDt4NKsQLy
ly7Qo49QX10NJhBv2f8+4Bn3KpPqsrh0kcHUtAYA3lV1qSiD3WULtXLYg1A0ejAY
hbtlwYhRw7AsoK8PrH2zHdcm6N2MCb7AFJNBbfLtpohO/NH8L7jiO9xzr4iC7jfX
CkD4L/xgj8RycFNxWJYDdcWN90TYplT/g6f6MajlW8jQokT6mxZ/k4nnN7e0jXmB
7VCqJJIU4DB1hyP3s3Z4ztNjFh+RSIMl+ESceayt2F8Fyri3jWuiY+TDjnfa8Zlx
Gh6EYiWHbdfjJ9RbZuLhLdwMkAAF3dToW+M3rYOo/8ohaxWrc3MZSXmJrr9ZNvjy
n/gjXWI1vG9gLiehYFf1UT+2EybKCCpJEKb4zaQs+jfnTRFrxhfM60aIr9zNxxaS
2Hmo+LCR+RNspndBM6k0eDde4DaGiFDTBICgNV0l8pTcbynodpySTcTPLI/3N8iX
38hg0kwEcaNlxuewm3oryp95/j8k6wFlIjVE/cXqBgGfMtpdVIurPRiD0iTRUo2l
h6yak5g2sXVsyuCjuCxOBQ+WqlME7Py+ljFFcp8aZnMKcJBJlcOjs5jVu33y7P2C
x1taNK3xFFLnTHJvJTjiDr33RBP8i7sTwgZGgmVml7KDjfN8sofwlimc1ewnMzi9
ggm9hwE0JchVknO+3OY+0Hza6vm8wOBKXu4oREinoSM+DEqOZPFaAGLKNcm4enng
RYomkiAAemG/OKvvJcI4fcal7Z6PWdnIwSnXGFZOG+G6zpBbRQ7uc64RWjLox9C1
vvcodaQcZ4UQsG4dNOCkTl1Scw0ijaQ/w26dl4Ov4OMbRjNqiBtLZf/PrX8aeBI8
oOA0oie9LoVrirBe0roJGWPF0VW9/p1HZdjvGXcOGny+HQnZZ5l9NustX9TiQ9jl
z8xgaYp9ii2rSmLmdngxS+0HXDnJBsIMJmTbDsf4CnYtVCJvlHJOy5q9Zi3q7dZS
DZrYcAxpI7nxMPGY63WL+8wBhz27ZLMdALgYQQ4T5L9U32Md1wk+zV50z9yIJW7M
GDjIy8MgUFK9gMLffjuV8wOEhyBnf6fFTWH9veTwmKcC6CplcfzDh6KVC8zwQfKY
IZ4MqEKsdPXs/o7PNc9wgr+2vXQvOh2Is0Tj8rPJl3jCwv2xRvloqDtse2/Upa7o
GABv4ldYWY1Ns5eukCnwfy++rUddLy5CbHUF1OHny+Dx/bFQ79HYRPok56jTnnhO
m1wvR+c1Zk6HgQBl+vyX3cQzVYD0SPK9GBdQTdb2/OJPiXNWQYFIMlQ5rBYgOV4+
ExubZu/1FBa1JmBH+tg+/Lpq1LQkbFalRgCXm0QXf/4ieQS7nyS3Yf2N+SRxomwE
mJoGCZqA83vzBtw4jL4q79ERi9MatztmUsohtaQr/NM8qXtysF6Qxbwgm0r5Zxzm
YYSgj7ySfuZhcb6XpYkjWdwwy0m9c4wU8XHPe0bS4+cmnnJy6dL7stPrj6aca533
rpSL/uiegTorDLsBfE39Fj4+vUNq1bzURrEDi+W6ICHgMTIewH/fOE9GfnREk6tA
P7rvnLtOV0EfQj4eaJhRf/C/BD/eSUXbj3yKRrIrO40KYZquJSgfPPQYsizutDAp
SpFwJwAiRTesz71y4fHDIz9azRC5K+xRY/RyYhxf1yBnriU1SWuCIk2KDgPQjfA7
CAKemr42WmiGcYd/1PYSKaiLEKIAoMqL3O69fRsYd9yiKFKHVO6kRYxHg+pzAArW
y9FGJaUnsCa5rfBEHuIJnjMGZTgBEynD6ooGzLZTwQUXjP/YAJ98G5cWuqu0ooOA
roCGg4Y6Isv1LzfRXWAkxJeefptkfpXQbdVBpF+Te9UqptYV+MdH7W6LvVJGibcQ
C93yEpviF3jRfiR1N2qgwl59Gwfn+p0s+KjF5wmn6vVuuxli58TVwFGANxOIkr63
54k1luqSsNybad9T+l7eIN1RZYOoGJiAhveHQ/BTnvAIVi3C1v9kEG4NXQ4RUZZ8
/7ihbhlDQSl3Ii8yu6ER0AqIzXffbTmDlPXCXwAWUEHJ+GK6rKFQLRx71KJLLGDh
vvnE7ioPZkcpWOvgloBTjmRBiMJzPTosaKHzuYmSUAI8e9aPva0X7FxOQgKTrxkz
6TRjUXSR1LCLcHb2kt/c9SR4VIB3/eKWDbg0WXw2EQzr/wLo4j9FWO3x3NUjpes5
9lgr5i34ECR9wM7T8n/CSxl64EFL45TLLJVvh/dQn3vi3dw4IW9SAvYwaFsJL5xx
VPrb9AuUEH3zb6TRqXwScQhZQqhn7A711qJQw9JD3pDSDbZ2wCsLF+LJsRVbM5Mp
s1ooDmNWdV312Tk5Be5xUN2BjxtG6a/4tBMuNFNqPRn1Nh5yyoDD/tC2FM50FU1V
T+VgtYBN2YGMuzBUnjtiGi96yXQI+UqHh2MeK7c8D2EOdRQrelx1cC4phoDNfNoS
1zuPXiSsCij8Y3slQveOedeUqJUcqk7IMLGTNkk9mhgM8xj2qAVT6YGUUcz2Bs24
u+ypPUqY8Iq51V08oREwxIKP3XMMGj81wxjyLWqdiCM0hWYl7HZrzOwmln4Qrv+R
PHDvEVMwiZTiOQdm/thKD82C1+56Ab0XWfGvLu0gjipofs7XRi7kRSgeIQGRN3xu
9zfKRlLlVUm6iIkXg4ycf1CqK+vgA4IM7g+IJuVwIdkGOm8EagCgHjSCYnTtooxh
DJfs040Dfz3abFXhx9rikN70ZwJvZUOKkqfgpweEmActFEsWD7450497Y6+weDQ/
JWMjaW/Eu1g82vkeC8jw/eICJAIrmS/5JtKX69EdQ8l+AsSky8N9Pm+/KboMBLOM
TjKC/mqr/xDKO3sY8GPYIJYdS1GOl3VP41rL08u0W+QvwNZ9Lm8B5KQ/lD976Lsj
87iUn3CCkw61N1WeYvvZsEpG4/wBqnNIx6DSXRM6Sy/4t2VwFaR/uGMPrLp2Ok7F
scQmQ5l6iSMBHaUIfNvbjm3J235PARrrEp8wsRpkRV0P8qL3YbPWwiaV1zi6G6Hr
dWk/aVzKi1u8eIFKV2TXHlQEOcxdw5qiLp5+hXuqs5vt9ZT1nHh47wB331R7oMQm
TEKVTFMIgm6aJXnLx7cVCgBUvxyMzH2QfXUFuEZ/qhbwn2txEUgkgfsUc3FzRFOo
OTViqAv8wx39M54g0r5HqX7A8+obQp9E1N94seXR2hfAo76q/U97rI4/tVRHu9Rk
tlFm2vZEglY+M9OX6TkBg8w5blHJVpfj/GeWmW002zP+JBX3OHvh9nOrBJGiMpdj
xlPg7ELEMeU30YRF0AIaBb5ZPF3Z1NhvdqS/z68KmWNdz/3pxKuvdU1d5IASUo18
tzB0L7Yo6LBlglWSuljSLzjr5HBuisB0vKHli3+R9xRUDY/6OXvfVTURY8Ox4Pmo
djsj81EvJEUKfFjv6Q1IMzrdut5JScWSrc5WUrgcUQhiZQ+nM+MT1jbQVp0C95Dc
bJPRufctU2gWkr+WcWe742SjwJO00Abg0OyuQHkz2x2K5J1QcEAoP1nxxK2nlq/v
Al1OkM1fqGHagnbY/MP8/hHHyZctNg7/UTiZYKFTUd4TUUbomi5s3pOMpfKbPBJL
ZYKIU141+RanhiSD6kzdQPp3FUO8mxDMreurSoM3jxayE56z6hssoaeMMvBIpY4L
J+wq3Uj7iOECoESfYfLehqeNGWp8i274aTE60zgE7wp2nRBxzHVPMj2a/nGo51Bk
Ky46JD37BZKJ2d3GQlU8xCVJ9P5aShZbAZSfm7DWvghzHYzk3Wto281/M0Oi8rAG
I7Cz84K+y//2cZosbJq2ncV4Oq/DW+f6U75uB51IfvubqaJZPMpQ3gI4whK+39ZP
Y/PjrtR3qWW8QQWj0IJ5X39QkQDk6HhFh96wABPXvjjwVc637eOSphtm8dM6hJHS
Q3zH4TLmOG3mPrCY0fpFsVml9hAwN8OYDf32rcsyljZCCWMOSGDPMILQ9NL8JnRA
vZrhrdL+WS0fyDZXN0sNDqhmPKmK8n1KbnLFwF8gmlDXrzaWt0eOhKKL2A+6Xe0V
lqUac/GC8ZKxEgfbYOVR326xBH+P6yXoTDgpvnLfgS7vLOwZ8pYItfggMtAHxtui
vjfBeyN0fDSGEBFv0h4mKtxLLB6OZleZWZSJyZaldsx+oJPkk9m8wLdHUUDicuhn
/sLjvSx0/dJ1NBwFLFJXT4s4cxa+h/x7U0r8hT/DaHJwvEkKLj7acMtoG4oyPGyd
k9WVcOEBJeOEEHH2JAHuGUQuEY9VWb0W/Vm0PIgX4dj4klJTC7cuCOm46fekvHLH
h4p0+NGMh2VZ0YkCltfaaXxJVLjHQIP2EaYpABseKYlnKr52gCwp1vOZR5hl9KnR
0hAiT5OvPj9KYJRJyts38mmQ5FSlkJVAW8pbsC0tM/bbaLq4MV2FWMliX+QBrI//
3ErfxpqsjkJAX35V959gUku1Q2F2aJactzF7ahemYXbk/BJ+lyYnq4/VmHwkPiUd
hR9rXYPin7dE6knYk36bqfSRmAGz8M3pOQO8SVuYwiOKznWIrmL+BdMZdgdbdEVd
Ej0s2E2RTSJDBDvvwIjFejSKUgH8i9JEiLi4r9aunk86VgqNzYzG0Tc2/ag+Hp6c
LeypfDf5NNpv9o9wGMPxZ06M68BCm8NJy0N3B/YpQmWAi8cwpQ4sOkkPADW9haBP
ZXXqOOG9c1SEJUrK6q1C3RPcV5ZDkJo7SH+Jgo9poiF6K+tQg/IX2F+3aZRhm7ZW
N40aeuBZKINaqb2BbRfSXwF/2ZQ2HLzO3cDgDSyVl2pmMwb4VHCVf9seUE21oS3s
Dytci41nxI3r8X+qQLZOgMLKetdM9cuZt69ItN3cRCdgLFBQr25Wm3oNqZk2Id8J
3tj8V89sx6yEZfbX7oYRahsqzvQBDJYhvv9DY/e6lCCM8YIOS2JHs/AsbwluEmH5
g8GnLpS0poMFP+Qkv2hnR5rF62iZ/BDkNxaxeqECBxfWRqKRuydoDqwZf9ZKUOWD
3R/mWqPpyuAQ31XgMSjmwYuHFeeLxSMjNRR7+9lgz0aILXlifHUcI4h9BRTwDBK9
TWdspLV29BMA36TdTZojV6kfh831k1vFcnXnClUbpliV5QLXux2ZF0x5Va4JJa3b
NlKjbC7g/MaBWHhu/MsMKZnD0gQaKRFDhTjLtRLbNBoI3gcWQ+kffQ/SnXHjtcWr
mwb8Tkb43er2KzsTvXVuK/zo0r/ZVHqUFpKcP0YQXkG7D/QXKCizayJi8U64fDJO
jfjIxXyDfaLVavw+zp7WA5PNRTvnJ6kAM/185ZGgJBTrwbt/qXL3Vd5AwdzbzmM5
ITyZm1olqe9BI8LaRo+TgoT35/oDiCq8TaNTBYm6yvOkk9NKRZc0FlG/zST5Tx6a
31i6gZOFYzqUIziCFKUHCjsYa99K3+N/QTYG8b/V86HdAGlFs5Tfb++8OJBObfbZ
IU4fM12EQGQSQdqbZdMTofbxKBppUg/h3DUIl8dfJ6n6lORrQI1dy43kw+vbjRmW
0FpjcD2LoZB/8kp6E72qSQNoaHaQFNs0F+uIBxr6QFqxLaS1fkxB9+Awqz02vY4a
KAxWmDvGyWo1xpI2BdTqL5QuTNynAUHQCuwciHpGVCCd28y3sarbOCLhyLP8PM9t
awZV0iRrEFXzBo+D2XslZpVY8vo8aPQY5TPzdc458k9oj7a6fGIKnVi1ZsQ5QzM3
lO6/PVGvP6LDksGlteHMrHqwX7aasxpge1MHHb7TdkEt+ujpPE7qYGvj0gPnbtX0
eAj4P6/6UmwQzKYgDFiqarpl/qJQHKQ64wpSGWz95hllRrNzgw5ctEkeqhwAZJZL
5y2v6peQ0vUezKy7y6kfiRe/8N2h/iJ7sjczNvzUC3jUh3oWd9rDVNKyuiInFed1
3DMNIMfAO2K5LDkp07dC3YaKYVUBrEoRyReSi7MxBYkVYPTZyWR8fVMJdgJNVnA7
CRLBeQGBwVSDmPO1gXBjf0Vqc8AVx5YBnnCEx8EcX1oXuJAcYHlckD0uN/d2tQ+r
5SRUm3/r7a0TTfPasDskFlYPAiWZWY0DApdVI7SBFgEncImh6KYRYkvrTJKN3KM/
hvOFTMxnD5+dDe1YzekB3Ny7zYR70byHAS8P7V/U6SG/LpLI5VQbmjBvOoYEHnKT
DsogREU9KjGK5pWpojmxzNq0NgPAEBBGLbdKq/HbVldXbmB5cjOYJ16x6CCG3va/
slmjNWrKJ5rd92xLflVTW+mZk7xWsGrdGVt6DLnj6JtBwFrdv1bIenE5HsEy1Cqz
GkSIzcPlM0Z2eDzhCoMewKOSFk3ePGc+OzAPwD99d4dheqmyA/WCdwsRJ489iJnu
TCO1uD1xQCq+LorvIDq71Ejfg6RGhiN1faqQIeJTzqFa0kFr7iE8IRXiGAuiY8M6
MMFj2Shce4/Ott+d0Zq1z0ZZN+pbJDWhnHWpLk6jxs45CDzpjHQDSvVQtroUPrlH
84L2BsQ6fgKF+ur2DXNO22Jto4F6itX/e3Ga+mFF2Vx85kqCtVmkGK1ylTghErmE
5V2thYo2x70eHCEsnr1NbuBCtm4Z/48cM3ZZzQQRKtby7lSy9PvLDW5suGNk3uIi
b/GdK1q2++J3ahG2zevlSBAc5oEJU3qCvAnRkE08uNZMwu4HcIhSUldJMpoQdmw0
4JF3DdUC5ozrEjWRFXq4hgEfAHYmLJ91DwGqLUsZwmur1fijzlxXob9DC3EbtpIm
PnxpQKjsAHjwbWDwmJGk5l7ai8aRUg727YaxpNXqQdDxn3IGc1EYRF6iYYX46l8U
WPKEkPQ9VkaEhtfpe1vlCagaPzmHBnWDKHAIRvWRkuj1N7TN4Wi4MZRrprKhkcxG
MJERU+sQx3asFWPcKhgVS+58qgIAOw00b9HTK21oUePvIE9V1a41cg2k/5+mUGLq
kpW0iM88MEV0du2i9YoQURD+e0MtsyU+fYuF3s1KvytfIFHd04VryEGx5OCS8S1g
KRiMjgtgZ3p3we/ECaKjgw2EhBiEpmgroOa+BIad/JffA5q6vVtHH4RCJIpsPpkE
duJmnKXB2RP9Qj/D8wClsw3nQk9aZaUCWtphYK3G+I8xPIMsiNjPQbG5f67dIKQb
gdLhP5ZXBSAHuLEj2/tG8MlFFMswoi6hWJFCcxreG4BA61hToK2B54mBKdqjZUz6
cZagx4hyA3sc13gfRLFpOpAZ9skj/kgnuYLw2O0/s/c1UhAgrn/IHtJr0SxtSdV/
T74yugL/OygkFhdWjFmw/c6shnwpGSPGI0dPrsKJ4vXMk5yunBwuOmcJDWbnQd1Y
f6x4LH226vluCNnPS7inIZ587/OXtdWznw24uy7jIXQb6Wjt7WwBm6DvRAHH0NTQ
2PwSfWOqR2mN9B/rPXr9zURFmiGR2BtRvV3uArvV6uJJltq8muIDGcEeP+1Sc3Dh
4GmY31JJNo2XjjnJ2xMz6WXqQsd+ibORa7AFqypOkvIgCH17TpiwHsj827h/b7Ij
FmtmNytn88BOygMz5w8bjPTS1ku9CH8jO+4rBQpO76DTvviwaA/IzM9cVk8QAFsv
KCbnotFYWpe1vWRY6CNWIGcIfeHYmC/bSTtXB3lG1lyesXqR1xhUHp0RVdxq0V+M
CtFBTpNIeR+THlLu/Xqbwdj5zWpIymUz9oMsAeKCqIF9pPffUTtoU+TK32SVabsw
Dn85oTTYiiMZrCmNLM3j6l0JosYzwclmRDOKvNV8oxGpfOtuhNEeh586n+lNhIPs
XKs5cDSrcpaC3TZOesIQ8Uo4kyKNaml6QgOzyOVp9urGOke2vsimJmoMohEV42Bm
H3C8vo7g/XcoroJfBq4zEGoDuKiWF3jfBM0svcrSukmZ3Zx5xAgMXd/KuaEn6Dua
FKWrZ79mHrcxtREwA6MgljjlWnJujzQLxXGwsAtO0wXG1DaWHtnH9pFl6KEvmGsP
7IJse3qsGtGzGSNCzGQomD7zT0Xon77QG7ufGxDKINJHzP4obMcwIHfHNdAQQs2X
ed551mGvrtFeHpXs+UxfEUlJdrq4jqqFNDwQrj/O9bI63q5D4ZybzsNAxu2zdh86
aswvy1zCIJXCLN5nqwd3rJqOTUJziCxZwdt6t1TztX0W9W2o/6/cpRVzJQ49QqZl
ZFKWpPTnTGiIqYdXWlcdUs/nUWRycT2DfyrBPE2C/gxlly+wb3p1S0OeS60U6o/B
l6nufuyxeFAEhLz1E/IE6CT4BILNQfuDhh8QxpG35OlAzR8X53pezNyDtQleYdoD
SDBdNcwu8Q6UTbTLQ7dShjdV31jZCnh6Ap7JrIdBgPlmHq66T1m/Wvnd4alQrArg
ZZhmASUm5Kjf6qRv8C65MgJ0I997Rvjlx17w74CkeLK7PO+HBCLuBqtOPc8ncSs7
KN8+WKTx2k27c55xdjD3ClyJYI6wnlZxKj0KpNFUNU27OgY1Y7hSqfgIiVMx4CQl
gRlZ+7ccJ8v9WSeBKEte1EoUO8+7URT1wTJg2s2OP3JJbceikPnBwhiMM3c3noeK
7LDQjUEDu4P4elGkSanyyE8nZlNzVw1wLqKWXPlFF0ehHGKhNUPC2Uf+AZGLShKI
Q217gBSVUhKnGqLg+u3+jiWwcbzbs1rcrWsdf9NbPEynikpzXuHQjj1lSAFFQsG3
ipYKq9icFCZi25q1rqSq7pnZT++8vDgJHV6Uxk20rXxq04KPZC84n5muNsMK8Sps
v/AK1p/2rh+rsluJV2prWBAr/mnLFMWbYljKdEKvsvbJxlCgj9grCXgU1Yw9nEg0
ZBhAa0AQ98uduJDBng5orcDSkc215/i0L5cT+oVGx9ZQ4tCtVUBNA/EmyBZ8WL5e
xaiYB3mKubxX/MDBTO9fHhosBIC3cJqh3MwHlnqMkAKK+CcUKxNNxTLytonpjdLy
zSPtrqd2JHDtWhpTDYeBvvII8k5t0nf0JpHJ3w9wz02IIpJh4ANA9cnfd6+R3fQh
4y249Tlia5OrU1+nXtYX95dLytLIooA+j7pEY7veFqsgezfcFxS637Zq6Vt3EMQg
PRnjKAxvhgckU6iuhlXU/5mbotdPEgUZwjVFgMnXp/gxJZqdw5tmVt8bfY3HfyVl
YbDpIKFD4+8J7Njb6INLOFLKNXKXw7ypMXBiy56bTPSJtidIdqWV6TecfQHxMCgv
6xqpOLs2O+KeLU01zs4hLl5fjDDdD9f4BWKEIDDvEpctBZFCRyw9RqqhUPTMIai5
0+he6xcLYjPr7BqaitmgVdfdPXEy4WE+QuxygbR6RemMOGC6lcdR4QmlPjdqzkr1
G1QDVrf7Vr302yVvq2q6QJKBfcWIgS0aLibCu+OBb/uj4gFM3Yf86GWM7d4ovYzM
hTPrpyB0k22EaGOiFW6alKn6dizB3/Hi1EX6b4MTdd31Yb6rvNFOW1BulTgz94Pp
qp8JJ6bYRuQ+0i4OpOYikpbLnBvXhYanG5TD89K1JLobOrIf6HXMTG0emVnrYx1w
36AsJclOpBMnIO4o6miO7OhhxKJEVd+4t4oUdZWjg1WkxFRwwX2gzUtTcbzNXgW/
BNI/2A6pBL13hpktj8ZHlRytIy2hPaLYbXLHIrjGw15oftPsVLQdCLYcsAmRsu2M
pjg05heNO/ADvrN9LdvefcgyNWbJkclZn5G8eiOKPKobgSrgpZQtRTNUFHTRQfZr
EfbnBWq0hWPOEm0aVVwhMxdTMVPIJuXntraFWBl9+tE/PiLRkLLJBmYfYhAOoMTK
fG8s1oNijEgxVHK/lspYooNNFfhgctJfanHWV8V3bF+L9cADpYN1DP0gX7YjJbrD
dyD5A2mimBSCAqLmzjug4Ube4ORu+KA+8+Y7BnFhlycJlJ2Whb4vN0Gm9miNCy+m
nUhHA8GGaH51T0lQ6lCus9PiA9Ds7dQzsJe8Gazx9SE69Cmp1wWfW5+UgPM4huor
8hXQGNcFcCy+u1j7SYT3O34gyHCG7jn+wECr7O/a8w2J6F2pgchVxHilDJPMeIDN
Hp3SgyjJeeYmO8GoLg69XGF2r6G4YrqQTXdY+yvRvARohR7VNHwuOG5JlE1FugEb
NvS6JAtrK8Yyk2lwq34XNqWOiWCE8JxunRYZcrRqhprGkWRVxZua3YloOCBCUQJZ
I5yHFhf8ZiBT1Cvx0G0qVJAFKOE1Uf1V3CF1H4Jvd9QDbP70VwFFHgyHjzbSecm3
XwuJZ9xaoOF1HdOKhQjNK4WJ86RuEJyWgL00feUT8LppAIld90mthnXZLsJrXH4J
5bnXtFrY9fU5gelAMOLJZ5RXHrWiJqiZV3BZjMR3cgZ4ZcM65UaWa3So8z3Io/nH
3deI3l6EFH0ygHfUHzrdrPCDvWQyxo3WTsFauWwylSsMyhgmARCAPeJW0JqyPK7Q
IuAFV/d1z56DvhOnpWx7uFuklwZYxF5ktAfF7s+IyMiSP3Vx0OFwDbTN6RIVbTNe
OUZ+0NY9wCz9Jl/o2BdqKtgi4+TMTSpDGNiFjkrSj+uo56ovFH1bUrrO/QqlxNOF
mcZBNWHZEJ5577LupuakC/USbRdj2cHUUTbYhf4erayH18RBl3w+ivNW2FrnTWwH
j7sgXakOLA3nwnc6N6evTNCXq8XsqRvy2QjnmTpyqb1668e1tExRjvns01EW8n7T
R3MD8onB+dO03lJiqMZxw1GnQ71muaV7pihqQ0JO9213Dd0yhomVuXMmQmx0ZeQE
OjjvNh3P9I2PDo3kA0zco80t3bivCCsx9kOZRgj0HgpefpfEaj1bc0ahcW1bkJII
OITF8S5wVp9HfAcFUff0Vp+6Gq8R1ACeAgQeyWn0YS95MAkmHJxzNm1FRHAQc6c8
tDrDk7diRA00V6rJWB+CzagghbqMzvxpBVObGc45qGibOvDk8w5dW9GpPB9NkMGV
4ceuKgsFdTKAZ0sqcv9YOmFnQBx2AvM507j7Q8gOf1WEWvJ/LYyQY5CPf0ASrf8X
g3y0tPgX+u6h/VeVBRoJFnQkMvKt3ObE/TO03gjaIERPWzvBAtltYB3h4uxwzRZP
FOOD4VvWI10tZuldLyljnpUPu9mQM9ifNXTl1IfICuRQOAMet7jOGTD7r30DAn3n
JepZzC6H8+yPxDQdMOPFyLH5CznLZFRfViLSPiJKbrhSYwyo+pmJ9xs+xuxftp0P
ZGwAR6ClcGuT/W5SJccCT1a+6genIYK8DyAdMW7D0m43L5cmSYorYBx72vo0W+S/
x23MsmwuAXCq9dIBY2Wzd7e5XyL/TIW1QdEWXWCUMoB9ek0NPvhTvkdaLo3fYFY5
mFiGoh/HCYwelB+mr2eOY+2ULVfakKFcxEaQkpDiJuQYHu18LStDgaW9WFoPN3Ct
f5MeUD+AxNPRKS+LW31RxmJgKvKJOQj+zeuU+zba7269bi6SIy/tbOtioSr2OjYZ
I/nkMUXGcgY39Ep/fwGMVTVVIDIXce79NuFCr9YcX6eUXjYqMpOLaR1xb8hF05ra
sbhV9RsR5ngMNd52JhvUaK2coI9HXv49ZqmbR9jJ6RQUrvPxDF9ykSIfJadmLyOW
J1lC6Sc+Bv7KeTmpY2knWGwgj80w7q8oVyE5EJmgMMu5XMQ2/bfEh5N6QWUDODr5
wtGMcJwipLXzkUBqJ9T0fk0VnDmhlDItxtcr8rIUnlUzkfiNcTxsMshLXqrbVi0g
RU5bM+nVCFWg7PcPBQ+k52wEwm9kj6jfLMhr5hTVfs8FBxrOQt5cDXtio25r2RGZ
SLs28H9SU3kBtYQ8s5Q0T8Oj1rYprU2zHxQnHsjmzsruv7zlklOCQvlyuKkrj29l
wbSTAW1JvagJMOpvPjI8vcsL/nJMX3J5VAdCgp5EVA8l81lFkVz+qfrojzAQ1w8q
mYTkr2dPirGk5fHonT6XsHz82EavrNQCfD9JmVOv0TdlfPl5/CZXg5MRpenQk0rc
Frh4xnbSQbMlPjtneFOfWh3QPcbh5ENPA1gyQlTLVNvLllh13jen2ptJA5Ivqgrz
QjZI5vgPJxJiPR27MO43V9JN+EkUVn+nMZoSjvown5WYaNxYz9wSO7ojmm4ZkTFt
JOgJJMMTMZBT27uQjYxSVA+bFUoL11rQonoHbHPorBSApA6fk3aQtn/Om77DOYb2
pns854B+C1EmfHxqP1RKTX9Xy1C4kulN57JVr88jH8PziWg5isfJZ4vV/cJFz/Xx
Zo7/3ozc6UHWSa4ySaws8an7bly6iodkXWACP/in+Mmfy2L6yly35piyJShQFn1n
+prhwXNBO/BLiD58rU5CbBKyudT/64EnzOsNEF7wtvRBUQQAcqw4osVk+a4/2o+j
UJHdlzCP3Ca8BWWCS5A2pOOszvk7K2QgzRr57m+M3rGmLvmmTnDI+rgp5Lp9Rv81
b+v7mhUg52Kd70GyfN1LauwdlNqOpg4EGe845YsE6lvAuguwzpgNefgl4ST+dwAb
7VCd+Vt4tWIidCXIpal0Ml0UaUw6NHuyfGTF0MfOEq+sy8ZebUql2a6JQ2QvHN2k
NK3OmcBDIv/uuo+6YLRlHL0tkaNsoEqTdLB8nbus+yfYkWV2HxHxQcapn7reXMU8
JwDgsYMprxCkb92wcfVW6JlNfQBMz0oCkOiAZ52kKQ8ZT2N9MmaT8XM0BS4cpSI7
CnLCKVUcD3ur4plRCqmhrWmliXzE6MiywldxTuBnjPqbpkmwTeU3Q7Y+676RVo30
N9b2w6b8CxRa1Q1+qaJeInlN5Ws4ysiQ1Vx5FMRtAEy/IB17KQ9L0zGQQlCKs/La
Ngirk/wpWdZ+Ec0OziV/8VHW5+igdmKkzsJ4OAa9WpTbRAV577ecvVCPJ4eACM9Y
yGoAnkQPpBiH5IXZgp37clm+NXDBJVfzb+YdS35Ezrd6U1Zm2DV4HZaMztaKsF54
i0PlGGApaZX/a7aBaXSFa6E89nBxw9L7SLqod3hYlRbJ1jVxqeecr9MkC1x5wjks
iKzxMFJzZE47fQRblQDZsCTcqrFPPJdogn0ly1fzPb8aMnaqqgzAr1v1htZbXev1
seM9CIcombFKRMxNvguoIQU69z1MlZkpYaF1s7OC2NmA2rzcu3LD9C7frLLLlvgB
vSRFWszCR1kfCFdEwCA08fkiZrADCrl6P1pHc51g5H7Q0FUAdQnsuahbrVLQ7KAM
D9cEjiMVPptUX03FHyRg1LUqbpNCrIVRz8UUwutgySUNXm5IBgfD9eQkGLn/nhGw
XimdGjE05bP+lpEMQ62S6JLGRYDrLIEEANoU6JsGm9DrDLs9yNlLFU3aKGleDsma
Il5O44q71Sd5hqhQWlIr9OaswX8aTVPoBJmhSNqRh1am/PuryQPzqMy6EcoaDRH8
Q3wpwlpIkxj4UtIVOrv5kBjqnlPaIQyuRuhwk5afUMJZDOTNGXJhTGZ4G8oJQzIW
quz+/ruqE2hIRW2vZ/Oj9ixqJAdQDynC1wALr5z40GQbkH062cKyzBYoD5jcuxBA
S4ADfpc3I0DFaVsiYemFL3KOQfHk0iDC2sFjwe4ciKxwZj9dpqMok5+Lw4Hvfit3
IxbPdadskzGHXN2e3O5iWbNVoGrQzPWAgUrVGAd9tgPKVaRfRvikdRChJg2SfA7i
d5E96O6BgS9pjqIo2vjsyahtHo/JWYWiZ9LKTyUMNZjR8jGRNAUVvlkx6IzsCKPS
4yNtUfEH7Jkp6o8Hv9K0aHvDj+dkjfcGSDWhOB5rUR0fpQ+mlARJAbStBjs4c1gq
ip76LcSV1vYNqOLggVT46ww0XqC+3d/NOQECmULBC473T61xgPBUvAQmnbPFD+5V
+rKD2irUd8tZEODC4/9Nh7RYgblXoSgLjDT/RVakyXgSSJpblmFmoxNXNKdIdIMZ
WZwfn6XLNlUYznhTQwhNRFpd41zFRC1llo8IAvmOwnvpI0LmPmliXkzGMfcX7+IM
y1IklEr65+02OGj2CtVMR9SNgvK/FZgI46PBJ9AR4v/CfMw11u+cIL0Nq4ORmwle
N8BqDvCIgNJgm7KisBHUyrpH5k626gkenkZgHTydlG0EY1sa6J7edRXIzS8WS4ML
BePsOm8K/f576TRwzvCS0c4r3WbASIwcCblAD5wX+uydA+PHGfmVMG2gzVdq4ZKi
KLadziUfaquHYYw6YRv9qomf2TJMA1dNffPwaONxJaRedSaFhTMKxfeYkjag6eYp
FWOv8TtKSX3M2Yzst6wUMabWTgSqa+qTLxItl6rzCYUOcheocGJHeIOjsHAJYlje
9VrwA6u7RVyGFLZ4TvRRSXhtBcAZwNMiGXF3ibzDCT4rbpfN1N/hHHSD/XzAc3MO
xHkW0J2UhR7hABv2LPtlSPQukJDQGdRbnVEie1r4a5f0etTAmOSD/oSImuEomKuM
TbqNuUEK0SqE3Kg4P5g2GxCPjn7IypkSsoaTHewcWU6jxDjFDu7RTsLuC9XdSuSt
Qp2dZ9pmvKrxxinXVI+V4HQFUq7QfnLzK71ypJVuCyFBvlM8QT17lJZVunffNxGb
2FVhMMAzL/EymmdzECxy8ZALdWqxWRy1bCEs9iAdkF2Vclgeq/vugupLmS9VQ4hk
cG+CeHaZWIwfbPzTKPZzEbC2q82GXpmaorPT1ZtGa6au6Ti+R2FQxLDTxh3PCNUp
E934uxy+SI26DWQSWv4UzRlJxpp0F0044iYDHlvOLkgGK3p3YwpK0JjCTQtdoZoG
Eay9iiINd05wLYpuELOXi1rUAhxIhZYmgQMtXtdAIXWvNj+wLOUWhlUiuOWdr+uR
q4PIqegm33vG4Dk6Wxe82St6f5ZMPperSYuTmNRw32RhEZl/vi8fSrjkvcFr1s45
8J+E1BL2DUzKhT1lLMTKGru/IRLh2rJRMZB2QwNe0sf15XGXSniWzzR8gLBrBs+L
nZFIy0pIkHvn1jfdw3y11S31/a4OhtYsPzVX6D1GpG9i1C8akudqZCM3N7G0kmPf
UsZQoecxjDcQfIodWjoO/jxFJ6iwSzmDxSyUyTdJJkoaxIXEXMxxlETKBImqgUiZ
R04nWD5JWqTwxBhheSG5Bqdd6JWpYYC3jSaIzoCw/HGhd7FVlPURPAWJ1+1x5APW
iCceyqB9S3436sAuk0L019Bbp6OvRlUKJALoM/QTnMc3N7imgIUHTnmcxWdYECCN
go6t9OTp101PqqH35G0FW83lExTUzjlURg4wK4rhyfXL7iTaoksDk4JJV53uqL50
DnIns+IEpJqUcz+iG+inH1nX+oZuJkanSxosvrgo3Kkhn+k4JGESBSYN9Nq0ZHFf
/5zBfLt9WWMcWL3ID35hyfbuaomow3QMiGIX0/qQFtvf4QN2Y9FSI3g3qaton2KC
9zS94hls7CdaV/vyXMlLrJMz/cH+sQosR45UCfAzMMwMG7GN2Qajv+8QwH2GjwaB
al9micZfItuNBh7K05rKNabH7THvLE2txDo4cPLW8P3NsookWpv0od0KWl0ZsOlG
TJGrG5rcBuBpuDTLWWTodL1qA3PCrACRsJ+X29O4NaaDiZxUooFyWRRjJO7s1pg5
O96LCtmYrUWrdlgJNVpL0Ev5fgKxsHWncoWrZ7/fUXky0Gm6z5ajyd0k0lpPugmq
4qLeZdnHvPqwfDbKmF/fgTjqjAGBUh9l/DFTVtuhGBX4LQboi7YhEFuOJbjkwe19
yNgld/bRhUOwtw9Xor8ORUi26r3SoS16HGe9bWCBuVvFlhfhCi3A/4HbI0drX0gu
8UcbtnkahYWA0lv1565rym1oTmzx0t6PL6esZcFt/4OAhktmAZUFswY5E0eU2Wla
Nt0GEHdz9I4vIrfx+8d5ddSzSb7E3F6xjr/35AbHV1E/mOli168nOsQ+7hwoNlNp
llcJ+s7a05Vg6ApitkNZPpZfhj5z78i8JlGVDSOHbhYCKpMI5iKhtV9vv25htCBh
PaAAXEAaOQpUPfBogFU/L8xRmoEMGyYYMZnma5Kbwr85IpHl+KPLUtd6ba3UqjsK
6Pr+y8Oct58bpfKxzaXZIQHq10TiI5ELlghR7lFIPzsAJh/tUR92+goLG+RPF2CZ
SXM3uNBDF6mGsEW/PAz9Bd4RKh8hmis7CSlQ+7pRdqQJva0d3ZfcHQ9OsdE+51e3
Ihqxy3qGnH8I/SuAOaAOSpSXQ85DcYJ50v5zT1sO3eLKkE9FYjsyhwhpUd/+noyo
tJaPq5QitP/VZd6ikyQhayXHnJPV/L3MRRQn3U2IqLGiLpuOnPz9EGEBqCTBvDos
yJAosKj+kcHAWN6sh/zGKwn5tYEXQ3auVW9X93ZVswOPNI98+F6EPgVpPl/7cF9V
+KgQNYdF9icwfaibFMMuDutr09hvo3i9i6QIOnop7AM0N8Uypacov5LT+h9Fhu6n
g3ySWxqgsBMYXamuNcmVXq9X204gGK7c2zsrah10SqA5uVBDnAcks+4jY275jArM
hGIdcV4XWS+A/xZBofz8KbFKXcK1+dN7HqPn/nJ2mAb6MJ8eaIE1L+DG1XRARtpK
eyPG1+ot1zXLLF/RwNqgcu7Hp06fFKkZOdqZRYyk42TchrJB07DpNksWpCZxU1WA
GY4/q/T0X5yyBMoQGUMrFF9qtQy26+SG96pRqKQW9sq3nqICLoRobTrNL3LgBMRG
JUVkVbIoNre8SEzuuaR1IEz1xzO/4jvFWXzoaHxlOCJW7zS+kapaUlJvbt88X+ym
HI/ip9SHzBVyiljhkXR5qgoqAw8z+CNO/KxuzOfQuLnB1RkDHzk8QZtCqJtqElx4
kpOUQn8hM2m5m3MDy85dIt4TTKcIzSThHXIp7Jlj6kw0hGVj902RSp2X7SQSI3ia
/Vo1ldEhgbw/BtYzpxxSqgYYtzgLyZ+EOY3x6q7lGJzcBVH9+nYroVq1tJ25CuMH
oB7mWL4j7J9EFhjCJBxkmit9szSPGi7y7PnyTr2ftFbHx6iRRumvvve8fDaI9riF
8pUBbsKdOp8Y1o4MJ1vKTMX8nYyqpKUAslAxwd6Zd8woTK3W/6DxzKX4wIKKdV5s
J1lKjQQi09ApzXptmbT5VIKw+T4kRERj1CmZWE//yep5GZCUpjd1KYYCSZ6n1rKu
moz0gxxfDCJCpuHX3fl5nqHCWDIaLQvELqf0wzztSGgjLZPxLpHh7ns5A7B+8Q+b
XI5cJoW3Kx/eEZhyNDhr0j6pPTi6UcdCQM5eV7T35EN4dmozcGFStZNooS56QkKB
LwSNauHlo+819IbPL1eHkLnx/f6vsq5EOMNkR9sgKe8fKLMFG56D5F0ALKM4aCLF
FcaRnFYLGM01CY3PbqjUGhTkKWxQqD2dqOLaOjgR1vrOrXWYoz2gR1MlgbrH7CrY
Clym/Hp4yGKNHagCbrq2jKUPmlCQaejTfDyLJYw1tJ55AwQ/XLvh5Uduk92mKHLC
wKmxVm18KY0AvAhGo+l6J786I12YN0Y8gaZdecCuEBBuLVTYJOwbQ7GprrMmg4Q/
4egDbflxHPE/L3EzOiwARkhQh+nc0cvDKnvTJaxPJBMutY16R3y60GJjOvZH3Tu2
12ZyoeZsYz5Bli5qcBEb/+Gv/Cmv+4i+yBA0MlYujadQiGxbM/togDI/0z1DJMBe
M8IdCGv0npbi8jY0SxzSXCs1DMI7afgGnexzh1GI92B1v37NOyxuiVOo2hi8Rd2a
Jfdni8rb7ACmriGYH6Hi5J1d8vdnCCfeQvKUipQZPMqa+jnklPzLBp5clbjqt9Gt
A3jz1tYEzLLrlS7FfBNr8M6Jh5Myk/foTvwfrK1lNZOB5ucCx/WLw1DyWe9GePKA
b8BL0RZGUyjsdf/h/TFD6lFD0RiP7fCekNJuI50IjL2v9XXRsrZ0dQDdkh36mkWv
nSJK4N8mJROf2GfVmYXdsDKL8/J25Z8vtAtgBGbstKclPsFWTUq/yzDG1Riq1O0s
ai6Tj7O7k03WjbTKyqKvrBQ85B911zcjo3HSIi/QrDIWDYPUVwYxQe0zrXppSnwn
0a/guC7rPPdRIneTbMobcfu91QO1VlqU83aRh2YL2U9J0wAsxb1PAh9567KV7ggP
mvDAok/ywrheu/OOxXKpU0VTsE/mJy6sEptnPNZDPI2NomtpPd85eIlT6PLlkp4O
qRUyKyT1epxrygYs44a0ddzg6fu50OtpfXNYGoygRQcHfzoTBagK6Gq84aCWTy9S
lpWLm7qx1KLCqQTxfSTcEUylqLtaB3su/0yZkkrONOHNSa7mCbCSTf/IC65Xhd1S
ZsgOaAKBSyFCKJQPjTv0FQ4uJIg0RQkF7YEXqaOTiaUhhvqqGT0woRVIGiek0Ovz
WS7q6UYUfwJgY6MtSSTt2TD5YOMv/2v+tBiYrRQbehecnXhSVn/bqStpMkEY6QjM
uRQH20dcobkUxCoIJ6gqAbLmVNFMEnByUAIgvyqVbidyuOCctji/N5aEGKxARK4t
UbmSGALnnxj/wbTt/CKNgO/cCyLM7fUay7AjGwya9gUb2W/rMRQzQmjQpjliwb68
n75V7e/VB+h6ATjs7id4s9pC7u43cNHz9W94qoil7QD0IyWTDyg2/lF0f8sbNUrc
Ss4z4yOV5QypO0mN5N1zwENuPgI6TVeSngUr0sYj3biaw0DCVsbl4NV83g17Y8Tq
r9W/5dXT6ZxdS/MeyleHHoPeiX4BIiZ0tEpTUDF3JT8rZKGVSlYZw460aQyO56uu
bsjkv5VEjG8oH/iku/3mb5jtq8ZJevOrETLldv7SO42Qhr0xYY1+qRE2BGFJ3avI
OK3ZbhIY7tbwiPGqLzuD/dDVIIMKJ2/VhpRyE16czXS/ooYroaPK/CNWdj3yrtd2
n7P0016hdzEVzaD3XKYlkq+DbfBBCJnpYAmaM8f99koCxKRZyQs0spZYs+4GgbPC
ejsMqanMxgInNw10yzBKrvOws85bW5h2pASWCX/oPEGldR6C7OnAtry+AdB87i1R
e2j+MUBsikLDbzAiYOFA7+wfF2zaRU+/7GoTC0iNOmoYas2and283wBc16Zaxe8L
SEzWhsaOTEXuzYWOtpoz0pIbr904Gslg6tta/rCjD6TUZz+IQK0nlITH4IU9qcUy
3xF8vx7rST7Eg5V36slnPSZCkvfQ8EkXaMI5KvkUiefyfT0MrhScqRldj1Hol/tc
EGXViD1zObxlum1T8rze1+MnwpvDoCrW6Zi6+bzWgf5M5ccF213o+ZWBlZTdEFzQ
FDmUYmnCoNZa/6fA6a7N6bx+PSZr2S81/k4BIEnATvRW/UzjNrUkq+1chj0PtjqI
V3Tvgrb63OGEBmTQCfOaTqH+7igSAPymAZYuM+VEby+SKVgdI8WVVdYfUNKxkRmV
HvaINn2gx/1nWvhRyQn01A6CFnDpN9vPoeU7NIewWhU8AJYC7RTHHSpO0elvdtKz
Vw3Dvi/tJLR3qV256insS2yndavfUQx9sziJB/fM4mlEcMVdhB92yBG/qIChxvqw
KVmekRLydwq/Tj5TQuHyR7biMyvbq6K+I+b7VfYFuPSTVb7z6PKKSxmjJaEWUdvy
Pt51QL+mddu0zpivMG1C7JNIIXBa66nltNiqs0G90ZclSl9TXhHz3S5MsdcTb4ek
LPF3KwrwCX+WhSKsq/7J1sm0ubOyPXvmPSSqcDL9XsynkPEXjKNwvCEQteqpjHb6
/lYhqzSdk5gDjgy3gux5aV3NET390H2F9NpT8f/v637tsX5r7u1due6kgsGvgG95
2iDge2gUhVS+Pe70eszHmDa5CYyIB6OxWWVLuqtun/lAqQNrMrHoLTySBQzkEy6z
YQuy4wl9/p3ARqVBdKGN+WIBTn+4oHkhuZBbmY6LYYVhZxMPIGAJLbLA7SK0lz2R
XvQRYCDxu1OxYZDpb6X/NqllrzW3NXErovZvisnL7TzKvfJGlFo/AXIWX8FwvRtJ
9JhlgbVHTAFUP26ZOvfnfBcCaERO9n/PeIGWuySi3KbNL7+v4GND6t/MPn8O5x2i
VThlRPKCLq7UXbEljgkiggW4FmhRCWRvACl0fuAX93O4cMKEmlIuhd4qzc2NQRvU
6qgumcO5Sr05cqScocATZt828kDFhbR3n65iNBm9OWiI1H7MM/nM61VPe3fA9Dnz
5jJgp6Y7iDwGYVZhnnfY14/PQI75mNraoUn/hc/DkigDxL6gx5DzUcMcd5DLGijs
YcmDUnp0fegnGUz47hoYyUgsvkqoR7ZUC+rcJLpoPm3svtBi8T3jBhCkcQ1qL0Ha
y3moejqk8jGSQBAp9fPel9Lv8o6NlvchwHJ0BYyfyNItwd4jNWaEb9+gm8sm1Eni
xmtPj4DJzm5G1/7eUthB0+iqTo55I0BSTmJxBn4D2XiiDqw31SM3SMJ4IAkBJUP+
sHz1D4ukBfLwpLUY6MrZ801OGNAC0l7rj9WKyfvl7U0qO6f3wzEMcqow4gGJXQ2+
5XZjMbz4STr0N7ly/zopgmr/X2R72i7ocYJMpSkNHtvpzs/eJYVLX+jkYuAnVwgC
ttZ3sTsMmTV5wWJPpq/ishjkeVrbB3K1rSlifGeXNo7eG9n+KRmInGH02l5/RshP
kQK00TAAOpH8aQFx5irWljGvikpba7nYGoJxGoZeQVSzrMN/i86TfDT6Vy+wr/86
CVYDIOX7XWJBxk3k7V/7QfurkU0lsOGqMZivq44ABaNAlGAj0iNgouYGA+c+jeO2
S5qAIMwYPZWdz8/eLkREmVlVFiPsTsf1O217tT8vwtES7exmxZ4Km+Mqv7kMbpW3
33gQTPDbw3WLZzOPrkFONKr9hID2ayfG0NPUgPtF+tSbOxk8ubDBkYZvt/I21zLh
lVZmn0V2/oiDGV55STn5QcKkHGbhOHSt8hzIw/jlftb4ZW+y7SSdPDcickeIY/iy
h1yUgk+0qENjyVgyX5Vfw330Ph0Dw2eHcdvrayHtTuq0AMVGqX3QpwCbxDtqrGSp
VNFSBKbLDdStsN7bMTh1bJd2ueHhBhyNaCebHqKwX/StSFf21y5+BE+koneusBtX
vV2AjYiIC1XRfz9pRXo7OsiqY+aqscosNDbPCkn/nfujzx1ExEZ1TpWPuoZ3miss
pA0CX0Snxzd+UXqWfW2c5MyK/Z8rVZstHIXxIV3djXxEfxq1I1HjsoCAKCg1fPfJ
4yU+XatOvi0pD10bGguDDOH/V2pW2ENr/lpONQ1S3Y1YpWvuuummHrbKMJgvoWrg
zbQjXWMJrqUJT2mfoLWm8INhSH7gFM36NI2WwtIgbl+wSN7PdE+OU2rBid42tCnW
/IXoK8B1OlO+PF814+mVrDmFxFpSvpMbH+8GuZqeEbkqtC+q5VNzt3GDyKY1de/B
T1yzCKEO3gcl064Ea78uBKqLWCVWr0KYWL4VTlsEZl5U/WCBKsK1gE+p0DbfKMnp
KKvEiW5EzhxsFSHhq88rDG8RdFzC3XgUHV4BbOoZkeUpEiHA5uYJwv9HaXHlLRnn
8FWgkyOzucrCdlBfOAPcK0FXtCjF6tPAG/olM+LJnqM5kdEzXxLSQvJHI3UWlyo/
DjbeEcnCAXcmWoV8ARKkAjLB+zSPE1Ij8vXxsiF9I2b93VBYbtvOnJlTEbRhYA2F
XEEw/WfIRPiopDI0Uk7NxdIfQMf/l0mMV9pFIf3cb2Ut/L36a+m9RThnA7ggTLFc
y/76l5+2Pnp9nOKQoGM7iQtnkSeRMKyF9z8uobViaZjo4ssgo5Tj7bi/2vBaV/Gx
dpf69bnwvh0O0ritmKMnl2o9QHfr9XGm6DaFBAyRCgtk+dzb/zA/HaJrqH7yEaZS
6q7ZbVsEqkpKrDtkWsXUI4EjWCaptfotTPoTStVw125rLS8+Ol7aFx6RUmS8rc0U
zgYTZp4EndMxCjfFUBiuS4iA4KIvsYRC7SGRx2d21egUa6SgHjxwLCmV3XmilI4i
Rc6HrtsGsrTM08WAAJThDsQkfLT08C2cfCUQarDWgG8e2tRItz9DP22O78kO6taV
SW9Ca2FyL/r3SyNUxPySMuGpqCM9F2G6cv1G/io7Ev4woayJEHY8ANSjySJQ9wSp
MswI6e6GVGnbyaIP2ypok4zE88Zk6hhTnv1c6PuYeNORvqZweGoJJ2IiJzal0Yzf
eCZJRx8Qa0Z9RiY1tMgC+BVyeV8bH6235H4Ts3fyU6Ede0hB3dRQjTEWddDD7Har
s/JWj+OWp8BudALMDblvpy0Ml3Nkkf/IRAYDNV53YCCbxDeA2uEiKJtjnLp9gR+B
byuN1WU9i8EDNQyZrzL+O1kq326RBijggRvttrfJo7Gk0+Vwev9v+dUYVL7XzD0f
MVkY68HH/k1yG6jVr1gvA+v5f83guodVzhEImmo3+yLL6tOnEktdYVj9UkchNiJ0
WbSdxEm6ezJ7LjOd0hWOO2w4igFk52kbqAmJgBY5OmdNtvsAhaw9C2edbAvrk1wL
95fefTgimGHsR/nyEDSLYwg3VhRhFihzwFZiRhHdgsU+tm6iiZ3XsAtw9s6KIslp
+8c+WKVLKYCRr0G6nuH9LkysDOqY9rCGu/jP4cLKbKIpFrInbwwNfpSDq2uGw4Ec
+cKhV4QOITPHRCHEw+VNuSW3dGwkx1JfSk4gUpHUb9g7MsEKGgRcKGhEMGMze7Q2
BKjjv2BgyD7lKhbujhLfrJm/R7i3FMzPOX1/s7Uw4utTAj/mSVWS8pzCoPFabjgC
FL/Rjn4dsmPg4lndOBzAp/QNzfsWCIt8lFj/sl0nGRI4YfaJVMbaZUhN6mb2DV+u
M5IvFK84QmwlF3MEfP9CVCEsVa1rMysmR69kWvhECIFF6oOEK144di9yeSxAAxHK
Ghubx41pPMDpq0g2jQbppdBB8x19ve281muAZ+M6pkqvL0FebQd36fLHVt7s08rY
iItpDqV57ngMK1vfn4d4fBrbschDXXYGcCZhZw6c5HebqC9SWSD2BrJ4a2j3IB4A
tDY8DMp6G5LWbJzhzv1B6f0UUnPcXKbBVUuPXCfTwVhlIMiRg3ZW6VkFOgJg8M+D
tloZd3tJqsnGQUKPTOTZphLFeYnfG1i0npDFUOhBZu2hSaoyx9vY1WAdLWoNi4De
CuYrggmrNtfGioeqkZCjjwht7q0UY9ONKnPOCZ9jeYgb/9+gvnU4n1m/CjwTXZnT
9hmCK0LtdKXG65zJkxotl+BLBDi8TbqjphFdUDvzjLj0td1b3bPEQ6D3tqaiH0zH
RgiZZrzeRFQkdA2VHcB4MCd3KQU/xq0cjsNOJdvhSnk7tTkLWEMVt1yITZHRLHjP
HHhu5lPfskMFao7nusLHraCHn3rhRFVnZQCK3LUjpG4OemsG6PTcNkwmzLZvKbDG
CcUO9ZY2caALaD0NRspR7AKKBRkqid8gk9henfD78Pz8cCswT7laB1Cyno3tFhBB
4M7PtbVHWelEVBe3wc8Q7I2RAZeAqw9IOP58ssQhYdJnIxAyCsofRtQFHvwdV9dF
ZHCrROUXtUx3lV8XM1rWh/6ZnwayexH4UJBH1FAYxvGKceIBbGac/mPpd1q9Q+z+
Zr9vlzJKmMZoo4RVHRFRNsrei6toUG9iGN2xb83uuqa0DtSMTFUeZSCehc/ZilBL
M9VDTrua6ITdkBP23E15XELVQ62XG+6FPS03fIFUVfX5q0JtRlGicd+4P+vVt1c1
lgjhS6wjHp1dtyjL946H7ehvvI7kkWMmhqWe+tCyRqrMeykMVT2wfvp2HY8FhY1g
j1CNH8bsswsZ33gLuOufXHvRzRJjbpspNJVA3B3XAqjvVM6nUNwlH9SARODRSny5
kOezw7zbikiTDH9VyeI1FclEsHx3VcAShcKA+KpBg/GJlnlALktP22r3JKGsHE51
BveYbRhcjcCmHSP2wChGXmj7fRlqkJ1bLsSZmKGH3n99t5EDocDZWNUI8Q9Nuz+2
zdhWJHmcBw31tMGuFsZTPYbqHt4Gcg5X4hV8Lc1/aV88+aVeRigISeW94EIEg0Ys
QUHFODqqIFBCMzgnZmWoS2UpWUtVf7Hg0j0HvY7SbsSJ1duo05/uyU1k4z6RXG17
I/uNwi8Zb7SviKAYF1lhFrXCJRrdJxdXwcjXTfugKtB+B1skyrTBIy3BdGBc5obQ
jgBqVVFyxAkmrxFmitN4jpG3Jw4kD8vmlzu2NoeuiIz0B2pDZCjnekH2Wjw/6d9R
M/3IswFUKIGUlNaak6eTNx6J8tK8aY32BnHEr90nxcujyVcqd/JKXk+UftCY1NU1
kcuCdoEWtAqp0IR7z7iUHjC4mTWSp7Ot8pQkZl7yJ/pHMt1AGcaREIjNc5Oaayd9
ejfWO7dpGiajjXTPpdeHbqGDV15WuYMIC9+q1lcpIXJfrcvlpK+qiYb3atiomgw1
Tr5Ku3A4wISsT8tqui3a/Pfa/t36zqeJ+7ZbZpy/JEZZMZkXdfhxdE/7dn8KSj77
oRhScnlAek1W/44Y1zbyUBFqe/LS+94ooZgRgTxvSIHGIggKEClGDRvKNWNBsdUD
f9Rs/4SGxqXtULSg1U3yQyAjmztsgoiliYlUd8iAbiU5oRqbinxUBgaSIYPSvGFS
qfBb4hBR9IpWZCaJQDQUpEWf/+SG6FPjcw0o+3WEBzPcNCrYDyV9MBY+y+sGt8OO
FrriG2FtNrvRBNTuR5U2694MUa0YYXmGGXSLsbJp2fLBEiWY/EdSK6lAhdZvdfN5
udnNKsiZt4MMQqNXHrpAfTWuBtKehEJxtzQ7CXlNrs3y8srD0ij2NNeANMyebQMp
fEZx3czlJcuj71tkuk3+Sk0avV/XQ4DSOoft+0UjC7P6Hyk7XIaFD/fMXx3RW2/w
KV9AM4nF3GFU71KiF1dfRiIyrf9VIlWHmzl2QgwgXGljnrWY6uhENR6bTLrAbOeu
rL0ZVm25fscD1ig/gYJye4VOd7dYrKTf4SaFA/UgL9KHPsa6tx+2S+8940Qso/Eu
JqLzEkuFp5CWN/whXRbitOQTMtl1YO33YehNNfiX4SfhvNZDnneKztXcRd50bSPA
R0HSAxPkSHx599JFmIbxQRI3+Uu5jsQbuYOcgzCdjS1BUhuRDNzhB+n5K4Md0mt4
MwWg5akaH/ReGFvikKi882sysCkuPeSolS7NZZ4NN6cFKREYiTSWahXd/MJg28+V
B8CdZpxBDNwtJolbCvGSRi0tZ7zcPidiC2K1knEzAwJ4ENjCCw6j+XuQao/lVeAr
LCBtXsDPlb+1li6hjN7tCZEYhVYVBGWlx/J/xFmX55KedchA1VdVrDo119AadNW8
mUjF+59eGOH6wnp2DcBkku5nYW/E3tH9TiSc5wk0b45HDiQo9Z6YMkO+8g4get6r
ORKYdKdqWO7EqF5FrtJHYf7jyw2Cu4ahQuzcdfqDCOXZQ0TSi1vg0OsDb0Y1WvyZ
H1QIF1GwBmVXRzJoAM6pR1mSWDhKU+ObDU5j2W7IGobjVvFoNgPe10eq7Kf3egyL
lDZ7AGOrOkkUf96dC8vbwDCjSK4Uqav7GMbWe8Pa5yfJPvCnodEpDJqR1X0VNzgI
YdrszrSMh8DGZ/EDRL6gcnIXmWUV/gZi/o055xbodkxiRusuroJu7xmkZBUmnxez
dkuTI0gVuGrbhJnpfbllIe9psBR32+Bb3lI4pA//9pbL5w9ZXQgJ8ZRBDkUfVwdA
PRHPHwYPUEFhj9qi/m1nBOS49Dj13Ywc1WtcapuA334aMen3ahYpbsCcRIx+ZRIl
o3NLawobwzAmOD1AJmqX86Df/0FjjfrUVp5LPy+XBLjDk175Ml9EZ7t/cNKS9ift
FMNUzqYyfooiFh56T18GQw+qkphaTCtq9H+hx79kxMs9mvUDJl/u9NRdY12QKiB5
GYoNUKN8MtdJ0+XQLdHIk2imHxIg/iMXQ5y5hUTJxDBTV5cVD27LDwrdgKDRtWC4
SzcoL67b44Hx1HphaTTY8EeChYchq2ESOd+10Cg3V4R6/FlaJAZ97Ij0CV2PcRym
a0UvoWJrNJyyuhelWqMPC88+0qIdC5lLcSplhGxDxBCwWmKxwDfCbrXldyi7fUlK
w9zQbb+IUbsEreRrDD1byauJHzJECNt6k+pM5uGfVRpoBDpLyFpb0ErxuprvKjPc
7hP2prpxo6sDMx4IO3W+eREHrY3mtF1o4HtGznEB1iXaiqEul50Bk3PUgk8j245F
vnZKaGIgQQsZ88j+Gt9xZd2sUI+6T5+r2Y6PO4xBErwkwK+cwrAuRrV9MjNgZU1X
Y3G7ivD5iHVqD3u4dcdgWm2xei04O4aAZ22tP+nWx/tToaMk0lizsAH68kCrSg8g
ESDWx88Xl35QN28xUk+BMBwFSLDcgLgaBG5dg89vR6ctR6wssca8QKZhC8hic0lb
/2iVJOz4g5D5a6VtmcdyLBgM2NmKKLrmKLt0x8jQaSX2DMTrMU6fwgXiuSqRck7C
gh/A7DQtWVG8tJZDDZ8c2ZM9UvgTEUFw7uUyvCb4CsPG3JbcL7QwBY9gSGUf4Nr2
Fpp7cfZaNjK2F149trguftZL7ayLqHVu8e/8MZ3nK+kFUnVkGoVvEOSx1ewYZOZw
4aFo5Skixn+g8hw/lphaH6NdU0s7Y70ZDkzECAOhJtEzDNgSBtPnFlNJ/XtrVLq9
ekkq2q4uiPBcBPI2DQL68Vtc8hxzHMrqGpvbVMrETMceQHYq+26sT5h9aq+X1c3x
NAUkojZXnYTT7Fmarpwgj4zkOOqy4BC3F86LrPu79aFismO9YHJiE+2cPhsVZ+2h
Py5ctpiXi8X+Yn6NpGL0sKnPH1r2fT/Ro2FdRBil0e2EuJopx0whfkN5xvyweFxz
djY/Y/OBW8iHJ6mQbJQ4x4aZaPn6eEftK9jOZ0F/WQcOG0jgsHItNS0gEb5r0CiP
fw7Hw4l7dobPazdDCYZ6cAt9cuat8YqzRmCjICS08iqtoecOnVu5fndDFFHBFUTR
SoYi40tRIolzqHSLynBbeggWLMH7rxlj7nQAmtAcUKTKVu3II1ly5I1pMm2+qmaE
9ZBRgVPICo5m1IeBc8w1jIC9a9bLNtVOBtd4sLFL645YgMb8oXQqGyt8kvRFfGYl
oNKXFrglu9Tu8pOdUqbtgUtC9HA2QwXVkrPS/3R+WTLVf42Jre2Wr5FdSOwRsaUB
Zaos+x2z5dihvV/5uwDINOf8wwJpenhRqDw8tjfCn3QBGX4v/fIFuySs11FXKMvX
qkAveLb7NUgDhRedwPsPhcxiX2mYlbfi7G48UfvoLjaUAsKtIMskIgDjyAFVupQU
TI00mbNgD5De/6U80W7FRCSyW2bDtqmWnrU9bygj5yQDCVxODR057r62bCWladJo
Z/rtBR6Dvgo4R19kHgO/9Oili4cMy33SI9E4VtZuwF4/SM3avejIgsz0L8Orf5G/
DsNmpiR2bHrhsEepQPM5GA3IRM10h+XnZR8Nk1v0sQbeMPSEIK6fQ+vQe4QHdDwY
vzpdGWUxIuyXUZrSIkN9YoDTzsEPjUj2MOc5k5MnsqbckVLXWmahowCoHLGtXaA+
UDtDN26XlpeBF+L5QXsmdcexufi1GPJK/IM4NsOiYHwO5je+ZkwEgObCb5yDk5Bj
NB2Y4EIlfo/5tvrSa4Q7z6XxBwagMqDOGtLutSNq8FYN0i3KDu8xIlKIFyIaT0Dm
kycQO893XfIc2kTwUs26/qOGmkoPvQ/JzV4mjUKxkItfp0xlfSwYSA/5zoSe07+Y
Kn4XpB9kQRmesuzpZUY7C+Xg8wJ9r6I/cl3hLgVIz3VAiSPClSW4laibQKhKcdNq
OmefddGkSyqivHKXT2gZLC52qoihXLmhGIguJk57V4WWUglsVf0QAIP/JmcWwtKS
Yy1z+wLtUahsMJVwE1mh/JnxQU6SrUxlMz444Fx4upKPFNVuPaR6jzhsp94hMlfU
fb/8GS3aNquu61pRUim7bMbNKC7oBaTYsz39Jqa5scXTVnCWdK5hfAYWbCkQiWU8
dFbqcBPIC3c52aByr6Y8qOC3EUxV//zZLkD8GH2Onh70qzyQtwJI13QmcRWrl8mh
6pyxK1/5/a1ltIesHWJnXAHm8QrOSyuylySK7G+fWy2IT27fNEv5HYVv9xRI+BCq
RJRbV40XTPDgbGQLdZouw4fZ85OstGwowj0da/eoqHWNPd/b7nEydjqeCcRjNEe6
xDGypib5KcURPJNNU584Hi82lloDLXcuHH3ACDJcDcW4mQQVM9mKap+zKyE9F73p
W+ncSV8iCQ54aqsdcf3C76WNnnl6j9rc16bZ7rJe2moxTVEOTioBSBrqMr7l+sAF
SOg/G1bu/bCDIueNj6bZulFi46BElhqPYYlCISjlHucsFPeCnLHvhTPwgJrANVfA
VHrYBf9uR516z14gPw25z0Mbt0ESw32g8So1pNhxIx1QS6ISn18jmPWUm1k/8i13
7ql2wvoAsWpPcp0rpr9KjBEYvWB/thB1pZYEy6OtCp612fMJsi/w19nXQ8fTi4eQ
kzv02embZiK6rArbplLqt14yCcrL6od6wsgfRtLFHFHtkAzsUa2Ej2wfqLYXlWiS
yv0EQKaD93/2TIMHv1I2sS5JEDraxn5oUOZvHE6uhYe5zNkC5/tqEWhCHnHngi8y
clJY0oKBA/ZSVn1LwckRSWoXStG+D713xCgO0w7E9x/Q/fWUdFocSUejxSZck8lh
Ela4Fd49H3HlFdewzGZhk8f2QxfGtg3/LwDlY11ynpsIvg4++kfdOi8aFh7W1LkL
zW28/Vda6AyRMg9si7NGlMkuQCCsOqS+3l0pw5e3mO1olzwrs1JOc6QaBqX/UvGl
+l2MBY0iMbowFnGqm1VD8OQj15k0OtvS/gItvrTr1JeJb/2tIKnFckT5qsRzzKxZ
PnoESc6RQC2OoxbDwU+ni6Np3Iwo2IIBFebtCuVmiRv4WCF6k3w9RZ2XADLSki/V
pLrqfrelWzDYNL5KNsfkvUbfVY1IptPvgeKFH20LZjTKV+JoG57SlsUcHwfc7TVa
HtBL9QY5DpoTz6CSjdGATc7uCFUgQkXr2wunQ9gxoyYkzH3CgW1lmZdgzxJL3u3f
2d/Pqx5anau4SPl8thL1RRJnMdFghIrsMUOgbk6Gd95FKxKsiJQ7ZMFLe/7R85z2
OjHcLaIBSe1yYiPEg+oX5FLDKtd+NlBPbHAT4NGHMKSRYgQMxUq8H1iPw+40qPgC
V4D8hEmiJ0by+EU4FFdwgvTaCrfVYNnEEUwU8INYDBoJExgMYn6WZbeiEbtg8d9E
dbakVxzr8Edor/sMzV4MZF0V60tBC7oRitflMITSwET3LXcMTKjDeGZPd+aiKrXa
idvTUgYHToUhlM+0wdFe8DB6Fs5RqUR8wA6/tacMpm882sQd+DIlo7gRDlNqifwx
bbHY7rwFUgvA88Tz9FQEo/SCU4mHTpmuSKBF33MendZsZoPhEaqOQ7ZjopS1mjEd
pT90UzceaWZk9Pc/ip0FBznS6RoHtiFZHh8qMfW8VEiLQ+q4aiquNPwwM5s5tnhb
0lGmUJiGATEL8OdYJ5kEkYUs17hH3Ah+MdTIMfBkXPcsFYb4i9cEYZTb5lwgECxl
7saduznZv5Xim7X57KjdRDXHB7Djb/+/S9Pj2erIh0ecnebzE7EN41vBYleHpbS6
v+gcSDVjrEpJvqwfulzuwLLswP7xi0+14J53kil3KS9yAjlb12mTDdKbCVH3XQY5
M9MJIF/yymbQKT6HAV0RzI0RZgrHkckXZcFp2CAwMpZ9vErZ9twZ54N1Zne0OCFf
MptUh62TScw/DhbauWxWwpcuXeGvzxOMR/qI4gBrn2Gkim84TKeSW+nlO3i1EsUA
VN3sP13r/PHHzp9YGs5DQFnXeUCcS98+Ir7z/StDP16jiF/IvVJORhwnRiBTlXC0
a+wY1dHAoUwNLSsmmOA89gZtmB9ArX7fIgkW51K1Wqg2FpOOEnAaTn9MYt1vQi2G
cvMJnmiKzap30YOdyJqLBluKGmWMPrVF6e62aJdJbzaeAFJmRN5enVtjTfw8FVA7
T2RdJr1RCpi8XgRDjy8fV1+dr+XXebLHwUF0W+ngkhHwyBedg6S3C2rT8til4Xcp
yNY9Vq4Zs25GxO6+5/onkjGUs+aw+DuOamwqV3K7+g5/+6cCmfIshFigmju9XfC0
BQf5SGyXC5sR5tjSkHaYBtu5pm1tSaY0fL0Xq3sE373KDy50xdfGoIMLwNn1Twx2
YMQW9Jn6r1WjqR8bRDmlNYakY5VBc+4QPXjUc+3dhTX9Hlt3Fj98N5KzHG6oox7Y
K3W736wuEaJH7INWSgGxu8ss3Pz62uPjBUiNVHAOjFkdyYUQmS3U9sNBESEhNAOb
Lqwi+QDcSs0qydwgI08VP3BXlAE/dc+Z6m0/HMUcWnvAfnabr9uqkoOonKKR5+Ym
2xUTN5VM9X/2Onb3j5OyWuZFV/URYFtIs3dUOHUG6JQ87Sh89KEje4KTcdnKxCMp
7Y/jPXMq/k45X4yXlYzD8mJa2LvVidg1bHg88qGZXX8I0bTDCIncFAblRDOp2BjJ
jCTnQvydPNnbSvWdvpandoMlUuiTtFMQ0jZUm2Hzym3HAYBwnBrUH1AOZnI3Oeis
BH/hMLXfrTEJNxnPZnarGmzFDcaYIHt7NfkBgKfsA3EhG0unwq+ybeQZ4eXaXUxZ
+5nILtZW13kR52tuKhOiIxLXR2RSTMEXNJ9WShns4QMQWWXWJMXxUus5UV6HXkbG
WP4qt3DZcH7036re+nB8+7JA7Lnr7cYCZ2YamKqCua1yAlvX0pQj0TeyJOgMDYfe
iYu1gR2bCUuzVR9eh9byI5zRsOi5sG9hilu30V1zhGIxqqfaBr49eyC3R00T4/Ck
ogEDe+zp1C5ZNkP3QOWCTCd7JWk4A2lpELiKbQ7VKNqC3yiuLQAEl1f4gc1e/gEU
abXTNZjOdOngsYEGtqeCK9lnPrcxb8LPlOXQ7RHetELB56MPLyetYYjl6KOYf5YF
4sig8KYz7B9rD4xF66opZUtOSv5d6mWHoPDZVSSCsa+6/TzsR8+edbanbLNdUbma
pE+OOq91HHvpEsmIj477DToJ5uV5eFdnZbL0cqlC+1i/f+mjnn9jWFvYgG8hv5/Q
l0cXOLpfJCIgyxse98UlYf1z2SyCLeGeB0Fz+aVelTPTJhEFsDJsvFWoKeJhhw6b
2wC5q4tE+0tRkiy9yp42yx/C2AoudNKEYL66I/GkOBwWZMRs0+pBeEqT1j5X/PWt
htgcEQ+RR5NSuBu16qgFfQ8mXPYzISLvo/3n+YGQFzr0uu1Db0PKGwwO4YiX18te
uwnA3IwL8ob7zUyemXnekFIg2rcx2ldADBcKli5fACmPRYvL63ElHFNnI09VAOA4
NkK5uhpVTG1cUBqRC3O9vSDM+uM+H8eTLYQ4vyrls+6YGMhmzcQSSWs77Htho0Uv
Ri2gRblkwa48eoX5TzT9fkkwtcAVVuCtTSw1g7jYPlRQb5FFOb5Oxvq29OqN/kZ5
CxNUTu0TFXfjt1dqz10Y2hrG9pfE6CHfmlhBKeRMW4loubAL8NdDcAmnMQ9Cyh3P
fIskIO0HDrMIaw6vuTCPLqdSrzXCS+He8hhOya+4aRgO6s+ym3SML7oJ9tjmQ9Wt
unlLxrX1o0VTdaQI++SF8tPhmLB2g7jwAjjRpxLjpLdcdeHlUZiNG9afQ/ndVcuY
T1t6HW12GDNJNOX51VIouy9RDYfvWcu+PS4S8oCylyHFUefFjdGUPuMPlml1SH+i
LgHliK6LCMq+OiiKFd8lPph/XcaR30wFdM2mdirQbX38Fc5MBRMrl9BTpO7r9TSO
isg8Ivs6C62dwnmD8STB2mdNxQ8CbSR+Q91+cZF7Z/pKp4NHq76wbN5ojUBp1VUE
3U5DAasNYAHMy5kohzPVX/C+yDwFdsQS9/nM4DJ0tgNKgSMc8xPbwvZxTtf+j1Vl
qCgmWiOtXVzlxtlbfP2ximD5VD8picJpo5fsEwMx/jGycJ/nH88BIeBfsZdlPxSw
8aJnGYdn3XdZW3GAJMLls8WxfqodkUFdYrqHzLhRDA/C1GgN1fePB5RI++OrDRlY
Ck6XkqhqotIAhqH57F0vK54X3CPGILC7ARz1eAcwoWVUaRr8e+yBjoeaW19p/6nh
3rijTZow2HtEeniNSQlgkgSSXtk/OE54vR9T8LoELGcHnB22N84reJzvv6ZIP5eD
IyWcZFxPWMtnRP7S+D64dE3Xn7minSCXlY1CMiqEjrTobgtN90vjVq8Bnq77hhbr
2DTQy2Z6G2Ixl+qkj9Nux8Xnt+wb9U5kMf3pZpEqq94+U7uHvb2d3Ry5jbB1Pf2v
7iolNCgEQE2M+ORuLZC95dreJGeehzkbennO74H23ec7lrm2UGTAJVMQF+8L5sAY
9qwBap6EzvgzoHUVwiOu5MPDknzOT0hhimQEaeWxOtT9cVe31KZygr+y/7VBcHSm
ey6cWZKRBs2W/ioEBuTL5IejMJnr+H7hl9UK5644Z6l4jFkL7NEMAtBaOuFEDxZx
AzlKebwS92/4IR1Js+B6W3ENMZFIPoy4XYIgxzsf6foJB383GhU0r5sYz4bddmtx
yqT/pBfaG59QDFeKIC6/l1xC6VFGmEm1Rj/ePn8v/DgF5mBkLo7UJ5phPu6Cvpk1
dvKyoJLeeiZ2bquw1lOIqeQA0smcKEjgHIbvklu2f5rnWpohtOGIzLJq9ngwwrOg
7ogupO1GyBdJ8H0dgiKhd2Kio1hlUd0aKiKgCeJFa9J/niUN/eO7PZtETwf7j66q
o6KZ7nzb6TOZNDNgbzaLNbIz9UvGc9pkJkwC0ElRq1WqpZ5ffZjnACoe8Jnwa6SG
t9uhtaA+GGaPVS1zrBW8qSeiBNDtnqh6hcSuuQns1deXzlXlyjNFfdr8Neefvfin
XheuRG+W8qX1cUkeslRJrCo5WDSZk9tEFTbGhfomUcThcB1dlEZkG5vbj1OVSUqj
3J6eCaDmUSD9tr+jcu5tPmZ1b4vAdMbbkuExu+2VLTwQgedOHFgkUwaDldKcd8IJ
ciTb0Wvs4FS1WscW+Czbqc2eME5b7+23Ltyc6jgKSfSYzger2aWxsyy5+sHmonsD
eZ4ztSehE8kKYfjJ0xOKWOeKafn6sup8w8akR35hat1b2EBipNHNO9rEx7aTIoOa
fAbNsjHfniwR4Kp628vmlMaAGTwfybOmGeEsMKL0KZbR6GYlQlFRyU494afrQUli
ZmhqDYBj5k+SjBbOSq0M1Plm8wcTMV4iAgD+ec5IDxsl9QvQy4e2k2tweBOaUHWV
KiIhGH+uuGV3BmZrntfcYbAQpyq0jW8AwMJqVs1Rc3nSBktYiAv3NRhwuV4kFl8R
sDQBw29pL4QFPWYKA2W+SCBhqJT0Cxc+W+p0zxTCGmiuGU6F/TRQ5Ip6G7iHSpFD
g5DNf+P9SPc3Fng+7NbFnABy5T2CicXjzUrN9bY6GCXXmHl6+dsGQ6y0rVYaLj7N
V9fENplPIdLIxdtifUPQKDSxF/HAuhUIpMdzsi58p3VBcZ/mBWppkt97TJt2N0jw
P1GEeY/KFjpGpginOTKlPB57Y2I+JkVVK0t4Pct+ZmLHmA5NGLONtcnV19QR+tpB
YSKPpFpAy6o4x0Cp+eSq9xrMzyF3PYur3bjs+BR5rbgRr+dcM6LFSWcqTFyKtJKS
RLhNPTf33ny8Zg5kk0G/UkTpzOKour9SuY9Dcd+XeyIXUXz83SywowFzo57yj0+e
GEMd7qPWCXGfd2de2e3UyWB4dKy+gGX+YwKObtuxKOVFjDJbdKLCyLge4irny2aM
P+vMYDQcXlsy09TxfTA30fYX8/iLtGyZddb738HG6o+i9YyD87Nws1AFDbPGpeyz
isy8AZ0/SGs+XjhXtPcViLq7XzBTObmsHgK3wJLru+sb9CQxUvZawy7aOo2AlZHT
bE4iyIxAN+gTSmErIIjcWNTvHZiricvfgvfGZgzp7IBwtUOmCNu3sPO5G6im3upr
8+YXai07ZoqWoQeZpys75LoiUwzkcWvOtzilduE11k3tP+RuJwONbjKSebxFXNl2
JmiFBWSBbUQtJ8tmDeFG4L5lHT26fWEutMRnHjlLJt9ud8hJ+piM9CkgDxzbfCj8
w7GYHkfHupTnJFvIEKGkW+V4zMiLlge66y/D812tC1JkEAI9KhyW3nUFFDTQFB4W
yDlPWOPFqGizD3A3VKZh2SLm4ZBMWr4/RkDvYAC8Cb6ClkOmbecsMmp+RdorysxH
jN40gnArzDEgARSsWWy8DSYOSbOgnBtDaYAugkCY4+IoeVEEW9tEbtwkNLWanVeA
+I9d5aRcXMLByFmNO0atd5zz8t2KHPGxskL73EzuFQD6ZBwM6wsUKNJ/UrtgXt2c
jDknBS4cmVS54yAl7HZQWM1ZlOjdGATeYpGwjK4GByASKgSfe7cPHf32HkILwaaX
419sASRUpoLvFaFa9vRn7v13moP36Trgf9Ia6k4YdAkMWKMq75JImwY58YruL+iK
oXea5/wFFWMdRukxgMUteAqVN9nRIvz8sKbO+Pn7UqOuQ1Ij7gYeqLxnVtCYt2MT
5u6u77XyxTDZbtUhoMWw++w7FWxLcSlSZma+wyYdVLFE7rlHOUHCp0DgGNHbPhpQ
ORfHNvQsN6hC5cmlzV3xEWKWCiVz5g+O87jXzJbtKoN2ilYDMeuA85Y3wjYPXv1X
DnvSUb4i771oiiZZgMpj6qFoS3XEkN/2nlZE/FdBW4zJiH7EhcCGSQW1pT4WpUqL
MU/DhHqJxceA/1/mUazbrI0p33SLjXOfuFS8LqJvh/dZlMYrPEYOIJjhMo/uA/dj
MWzqLzc/6jOWTuSuqJ9fz+n09H3LCqOXQZkloi0RCwjnzrx+kR2FAnp3HZ1e6LL8
FEw6AdG7ZqeoulwqXEBTshZWAF6ucQ2C/s1My+00kaIMpT1PkvdQdmGXF4KVh4lP
DelkU8EsSUO2DJfu3+QcR3ZrHTy67sQcrSisvANfn58aDbrt/8zSNMWMlpkuYmRp
nEPS5rSxfpukUpog9QWdR7gJLakEgTy7HcbkQ6Zw/8jy6z1UlLueGH3N7Bwy8ktw
Lb1Yrmpnky0WO3PgQvp4G7pkXv5MHym+WicWRGv51tY5BQuUzc08mTtCMJul66ln
9cqFxz+NktbPhibsj37Kza6buVru88KMBxM90e9aee5nvo6QPn+SnNNG0icjk/Fk
CQVVrRrjQl2cGlUv/xhxYqbcffpCW9/0ioKxBZUVEg7/M3ejmTOd5z0TpvbtHODh
WrIYMMpkDSBbO+30fI+Le+ZdKHcncA1jI0yNJOxwSx07kG4Ov+LciAinkYH29S/l
h/YeP0nJ9c6pKwLr5Hm7ve1I3z7GOQfeEABXNC5uS52pSa5NZGUtmlezGnrruUO+
ZGF789cwn48xc4gafV/4dT5TkMRZ6+Gq9LMArUvHDXk7QeKKVIAu/HFVTFDsGDXS
LuAbN4ydJSDY3n8olAHoEgkfI4A3oNo8H1+jglFNGOiknD595boPLMB+Wz6t0lxG
eOAxSAln7Wx88K9wM5jSkF0dcUBa1qBqIO8xXu0sfi44stYKEZ8ClEB5QUh7jEw5
frfPn9HsOKGOcSOz4y27B/iPJUJnZmMIHVviJXcXfJrzgWdmLaGSRkyKdqO897DS
+LLZaC6f9IiXpFbKkInXlglbStKc1+YamDpzdBI8bFgHrEEpQJf6eHqHaHvZGtwt
GN+po47X+u8Kd1OyH+Zjc5EVD0aAccqpo/pROnbZxPfkXuQRY2jzAZBXUyGJ9Mue
VwDQQzHjVyGAdtEi/Q44vWAFkSCxlxoLpjNZZrZZDmYBrm1gMy0RiAS3iZZy2fuE
tkB294TJPADHyeXCNpAvqvKn1kPAipMoUDqEIBHlWxRY84SfkirD9ackCSDxxSQ0
m/7sF9s7t0HTx+F5kmVhWFkjjJZaoxo+PWexkIE7ciCZ4ogq0vAw4bQxWE9u/mdt
Ytarb60vGPNp79ap2x7KmxKLPqHxIVfuSNZbAncD3ABRoHf/9y38BEOv1x4Tgj96
xTd7Y+gt6/G+4sOEIjCnBQaV1NtIJKabKnenGGAKESPgNFmiSBZy58M7VGx4xVL2
BzIKoN8MS3pKHQytb05DEh6T2R5FSZJM0P43dra8tfLM6yB/tqi4iHXXSnPN1bwI
0fq99hRD8uQv6qD3065tpmOnhxtKjwp8DkBhJ01VcfAo2VDTzm/+xEBbmH/4H3jD
B3l8e5MSr8ghAHMEXIgIxr/PCVoY4wlQJrfJKbbdMh2GhfgYvrJJ9zVAj4Bgp7+Z
Gdmfd1CdLWFN04KOGsaoJa345TZGh7essUagP49/1HfoZvs+cpaCOmQWhMEQnNCA
Z5xW0BQMMCT8aLYilGjme6SFBuERaRJUZ1QRnbMGXIf+42pCPdfkyrP0q4FtG28h
Z7QuSjgWwpxt1xG7lNva04tseO3QAwKOeQqASzAm8u+A7V7V/+7/V9atB/sgmFHf
qR1LgThaDz/Wdb0+LsbyEhfuJRjaXrcqaC1YLP2rioCMZAC5VMypsBmBWf766+PQ
+p9LWq06/iq/t2uRyq9bjwEqSMoXjS0qH4b8HZaE0iY+Pglk8T2TFvtI2YMrsNwn
iqLx2P1Wj3GqN8pbN0mz5O20pH29DtUU/jS8IkSTEyYSw3ssILmuWUmuh3ApIhRI
NsRkJRSuG0ebycPaksYzwgJMU+X74lVG1t/MRQJVrDbt80yjkBCyq838fZPO4JIg
wfY89z8vrPIeSxOV13ZQeDIrf5U3JEtJTH+5Evn0YQbbPzW29VAezLrOx0gSPpSm
f4ezD6lexI4j4jhcJ3YDFAqqvKytkqBpRVEZTQi0/AWBvKIZiz4W+0PIliNc5/5M
fgiVaVXgyVcKNVvbg60IOgvJMri/rCqZ98CNds9zykB+eTAsgwEs221Fss1cajtn
CNi6pkytyI/1zmw/HgHRg9L94awa5j/l179GEbPyqLSgcsGpElphqk0cqlxXynp7
8iarKFiRu9DO026v2M0EcmhFR0ov9dCXYDrcfyGU04pxn7Ts1FFFTYIwMbKzhhmE
pT9Gt8BHud/kLpF+ed08LQFLwvl3veKAXPrSQMy+izPEG8dwSMmzTEzncn8FInJ+
Afm+G8c7uOaWzyzSuBUPuuYyThNiTuUvZK0iy8qabGFUb6HEgrXWsFgfTOG8qN8j
qpBuc6yUabhUfpNGbciuT5CM3mAzIosP8rpJUnhauGG+yW4bVDBSBfXmiW7scy7H
glAkd0LN07JbolNd22r2AskBcc8xbzBCHAqYi2nC4aHrBWl9U5xPIRWpjoy7iwmc
Hb2Yj1TUBZonxX/svmmmy9RfkiPDLVs7id//CGytHI+vivehZG3rrdfKlQQ4n8g5
wU81/TVCPYcQ7DmL5BVdNx04hNPpDGSGB0r3ER/wGz0UDrQaUt+msSpfGgPHwlA/
woqQ4mtHN0BYzZWlLuF4OC0j31/a5WfqeyO3clQof5Bt/x+Op8iy9lQmOcbx9pXS
zWPiM5TzXZ3XI86tiHpbv4czoE+LuRVcge/8hve0U0E2LoiukZQzPKv9AxpgMllI
ZYsku08QJlIDI0s3YQZ4i43j92jYKkAdKM3KPLBRM1TRCZDnhjce/hgMdL61jbI/
U4IlqTd59HZyctXLQ/CYbsEW5ZsbXlCtA5mVhvqUjzYaWJJv+aVlNqiZlu4xA7am
ytxo0qhjg48ZY22nk/rKZy1Kbb75AI9H6tw+tTVZ0Us2it5K9mgaokTi0V7ojm1f
KjnOfKsxBsG7K7fQZd2G2VljzEfA6dLZOidIkIYrA9Ay//8NACJC31zzCxliQ2M3
LgYFHBrnlEqhJPLluuuCOEj3RLhX+3neMukaQkG6W/OSMz/lqW3oF4W8Iy8CCc1E
O0+MU9RrETmAMjEJH49tgdpT2Ab8pOMv4nnxAXvre9LtbCc5kilng9GyF40wuQSS
u1X04w81jENF4eISMq733p222rBE5JexB72NIe+uAHjeouL5mlXjFAhZKTokJi3W
Idh/HxUwQtUaaGH+8w7rR44FdiAdBV4g9N6SGjyU/Je7wkaiXsOowgQacaWTTv8s
kremndHI9xoQuNJyZIDb/w6HnIsBiQ5sW1veOn8Qv5VUuXPIiGJfwD2M8BIJX4tq
XaXpMS1263jAE/Swuw4l7SbmgSi7mV21QD+kdfnot763cJNwsVUmrEPF4ZQy8wrO
o5goDNuh+TZt6P1GZM8DecwMVH8W8/cam7v7GUmL8taCZJn0YmviTcPsaQUt+H/J
/OVzYf+e5LN2zr+V10cLpQ/YPEoofXg+I0uXgp+IktYLYt9sPuzKqZV6WETTxKRP
OS+T8qQCtBzmvX6IonquvfvK9kRsr+5318wGJgeU8aULA5+Hyajp7YdtR/fDpRK0
/sZdZ6nP8zodc7DbX7KQuFnK42rTnh9fDzV0hr1QljhcE4lpzsrPUUkeS+YUGyNW
xaTk2AmqKcXRGRofkuCL/Znaey8h9lDnBwKyF5Vk8Z7KPK6bt0YVHSRivuM1NHDq
oEDS2n0qG51YGDAyvnGcnZmAWCxOHg03bkEfQLpv5yCG3j8Fj4tXzx6pKF58VMs+
22BWGVnA9+HXK4858z1l5GH9cP3fJoiioIpPrOUDPgmL2AxUnbdkfvOL/UfvYoIu
J+rrQWvBrQTyaWUlXaPvhQqxgIYVrRNc1H7pTFFEqON0nv/mzpkcnycHSuS0mfzh
zv2BQwSmXCwaZpoz34iJD76LSHCpUiNAZ/3spoArsBkLl4HQR6nnAX4fBy+oTF6S
7pKnEA98WvpjsO78o6KGdkDZZCB5JPp1wCF9YJ1xM3xBTN/aM02O+A3pwbDu+92E
FG6KiWoqciOD7pLrjrqjUhBrWCLF1Yi1uj3a+UbwSDuZcD7R8yvFF1zXzbTjs0zR
4lZ4waqn1+7buKt6E8ySCrWqsAcOGdsStG3bw0RHQuWwBaZQR9Vk0eU8FsjOZp30
0JN7OAwd6G9mMMuoewwBDZbbq9LwKD6nBYGD3opcUx59TfVOUAvEStI3puTFwQPd
HTWd1e9PfhRm6VqfV9SRtXsdnSkpKi2vHCztdKFC4PyWmgnruxC6aFb6hJS4Oes4
6QAhm76SQvFSUxY+A2/aXKt0HRHSbTDBaLzqE6Blb0UyHl84rhfuD5qqTpjeDFTs
uhoQsDrp+9zLFwoV/C/l/snijDCYfeAzyKfWyRYSAjpcUbvwfYPt7jf/t/2iexSR
WKwBKw5xT/TaGlivDEkp7Z5KgDQZDXYr+XUFVWv7ITuopNPVzi8fviahqmFo4ALp
TS9bBI+w8PEAy5tij13xlWlXLR1K3fesNc0Gcydwf9uYO8Ma7Jmly8SKW3jEgQdO
ZwYIWhDRWiRJz8nj51plMk98D/5kbHfVxiSd1mCI0y4VRvdCipaBHMPJQzhN/eCZ
poSSzRqwLxn6v4sGCOAzWehADgR+kuXBKVniAAzujJ9fujd8j89lsddpCzuBURC1
nQEHSqL8htpeKLG/mSBgyiWq4jHnoRsafITbaLn8HeeQ9b71VtuQMfw9hTveJ8DJ
kZOxP3uNFS1ttHBIVBztQMAqz0M4EQAlmjNC0jIzrdObPR9Rrx6kD/Ut+ho26xIu
CUIOnBLORkcc+MgeA0BNntC0zaN3gkfw6v3CBOF5sFyFA4FzVtfy8xA8Agitm7/C
NleDO3fbMAW2YrmzURI5RKFySEEeEwYg4XZRI0qrjCe1W+qz0dAVZFpT1GTq7g/3
O8s+BTVKUveu7MhQ/0C76vRfCgns3Ixhqayr39AfbFREvPjdJcSFRbJg7BfDQ0fB
xl7pjfY+N/0HC5K/dRSOf/UZmDTL2tQ2Q19C3rMglBIJfMuqO+FfphfcwYKhUqtK
fVTsYZLjG+2mJVLsaFdWoEchwRCnhaS/NyJQqxwipw6i0AFXjytVEzkldJHcn3e6
HAbHBtCp5S3ff502bQ4+ohkTG1n2IoLXJbtH+qPVfLvqEQIXRtNO94CiwDQAi26w
bGqY4aNU01A9SgmUzFQe/Lx01ojDkZSDYjwk3afQUjupwEIYG1fC+UGNIBxhes4V
ui2GFdLiLKfs5MbIHT/tDySFBIIY3BlPQkGDvozBiZ9PpxuMHaw31zjKi/Japeis
xDLYW7gkVijGOApXe8UJyfDJ7gMKkg4Ls6USoZ7ZV3hkI6S74jmDlorHZ1+V3naH
VRro1KB1TaJ1rUNzAh03J5AMtoDlsEiLyrF9qfPzIjO8ontDPJFdF1J6+A5me2VU
OtKzuN7b3s4LqwJEHw+mG4IzOc7V9N3lAaz1b8MlTSlkyLh5b5ZefWiOKriu7db4
hRcBv1cGmO6ip5kf1Bq5xn0Rm2+TvlnNdFhy70bpStdZ5D3IJjrdvX01+kARwdWv
O6pLmsMB+JlCuCQyIDl93Wu9r14+/2xQZoHxUKUKGC0jpAH90PB/JjhAoGzkQ8zP
UaEi2QP8EKeTIYQTd9IhaIlOblsp4cgbqlyepQ1UHf8nF/Hvk+803dm+vfbYZU+C
XXxYdJPc2ajH6AsvElmVrrwVsWvnDZFTRCpyT9Kay5V74OlgSpQo+iqJQMlRwEqD
dxsgBf/WW8AkI01QzFDNQSljPdAYarK/vsVco8ZBJrz24bTIgLn1w72raf00OjjD
8EDQF2LbTbxV+lM0r0P+J7arlav3lzhQ0x04ooxLXs/VGeZHbEvXepQP0OIUYUJR
AZtz/admwR3YO2qVYfrOUL5WyfFuW3jkDeBvhs0aNm8MaDiiNkxHbkYGMBcpDnU9
W0ocT1t14LgnKT+eC/1psljNsK1kZBf8hH3WDCI9TNOmgojBBd1FeUlXHmooeudF
RoHziSGBqx08M8kQk3tQlnwwsHFgjUzwW2r8KfEApOnkC6VTc6V9Ry8K/nh6BojI
7aA3MLx589bTwXSvMShAtT148gubIIsbWf1Gc+utcZtmHLsoXLZaDLqDD+3DQN6c
O8Up4BFz3FoEWR6TBSgdsKUGRrWFVLSR7JRFGleMPOB+IQxfZf2+4NY1g9VTJ+GP
NEGDCCBsDes42w/7oGdmGA9OoLsJi1GQdWaeLhYFSkiEC7v0X//ngyA0VaNs9dgm
xE0UtSEUrSkR4oDyeyOSdWBTweZf6sGS6pZFYHlfG/6a6qP/Bsaw0OXVpeDSP0JJ
mcq9mPz3Uz2H/Kz/ywtujJltJa4GYkHkTT5/nwfi7kIZvqce7dCHOEVbez6Adfdq
AXbbKqCLxUgFOEd3Vu0Xq/lcb/AXSpDs9A70N+kHKvcXJC/6HKmXaLo26FhSSd/W
Gq7a/ENDjWuLCWPkGcOz36L0Ehw6csdnBuuATn8ydkRGD4agLDdjB0DIo51z4W2g
6pKDFWTTuyJjviQkHEd1KeHkNvFtvQGC4yUKgidbG6PO0+Kn8pdEme08TkWkjy/+
68pFnOX2lNyZp3g0x/Ym8X+LC6Hv3Ap/DzHD0svkTyEVwwMewC90xk50SZd1aaw4
50Z07PzIn9USowgJ/K1BJJn3ShARaGsL58mYh9O4gCLeTxmw/moPPWZDeeKIxgYH
R4T3ct7EB6R4xlvbCkBawmQdCHjs0zQ7JGdyanMv/KtTskGFOeUfq0+q4bStc+uP
YULva6/oywipllDOhWmvQaHmEl65FVOU5PbckOmoRhuJwAr2b0HLnEhiJF7MJuXP
joZvI9bZ+p69DkE5NaM3ZLeRh2lfCJm8vlndW8Sqyfg2ej7daSTSW64WA2PipCyB
1/aOhiZumRndTofs8M+ohM6ViT2Mjmm7FBlleWMp5uB3DvNYHog3tsbyUDTETp/u
gOTSvXGCmS6QmmRA/Q3HVOJkdUuHz2sZBtJZ5EF4WGnVhubVYkx7m1cnerr02fhJ
32QJAk3+Ozh9BYayG4yPMxyDZgUofLgxcmGNOOcdvBvWNu0CIxu582lRFQeeRPRn
iHpYSfOmwVJTsgZYMepx4MNrdp11IB3SN9MeEQBP6R7xb262ns5h4FlfEEsxPcUD
S1SEZgzoXrleuqOJN7PQQPsQ5jqXaYhxgeZPgYZs5k3yvoljUGZoLsWitJxuWN8n
4u0NU6oMFeK8tybMDP6T6DOZgG778z77yIQYIizlz2ucL8t6mC1X8EChVc4zxM9r
JyS+0ClygulqMPlG//KK/m06rCMFH3FtoNpM56JqGUmJtmAgOmNfN34WwnKlKfkj
uhsvUN6AZ8GSsIVc1gLtM5hM5OTnzugdAeAHASD2bZcGJUhDuvuQAB6H6qwSZv2K
Fnt2gNLzn7DDym/SROFtZyAP4iusjOPGrp91pKWKlqOqB4OW8JUbUUZV6xVKxjY3
Yd4IkevzuumsvXXFq2WNPuvYQ4m/JcclbLtyG3rn0hnpoKTZv5Oo1uXEh3oe5J4i
Dy0CYxyYQlsHcpeW84+XDNe+HtUJKr3rPdNF6tejsgdU8kTAOtjAeaDhA3MTb0bn
f5VL1HZfPFVA4zFixLwiwEJehUi3OUlbp3eTIbqSzH2MRIUQ62oOEHhPJUTaVrAQ
T3S0gqHcO3S8Si7wAuy/vsdISyRgpCs0fidtXYLjaqA7RWpk8mUFMkerOhfg/RqN
PGPMQrCkvzSY8DPD/mNOceEui1q/8wjEnwS8H+RfrJKwVOIepnP4tFyWEJIbEPW8
+npZB6N6IsHYsQvsoWUNj8s+n+1f4WLhmZj4xPUSCPQGmwHhKPPSmnBMbbobjOjQ
HD/63/+shve9iH1o2mx/yTpNWSu0AX/VYtwAI52BL9sndMsdJ+Dr3WSGOZOb82Ug
Gr0ZktiY9wWz1ea365FFwaum0C8B0YIMbO9DQ+m3gDbrXwgUbQnx7F0DRfMrk1S+
Vjnq3E6DxJvzM7JEhrdTicOte5Kw+C/5ourYypq4ClL/bX6IcSVEg6oEO126LBPo
pXGQbTciOHEIF8Pgrz/M/y6RRz1C9VXY9MpsO5+w9Ccnhrb9xmTVBmTnnzuGCbpW
CVq1vsC5rJJIqMH4Po0zhWW53oE37G0jSkELxE/dXZSl0G8WtYY/shVCwTFYxVPc
VKgoKonbbXUWAvHBuaFJlkEE+aT/PgrNr0iKJFTDuZVwZIy/seIO082T2q6Klcu4
vZc5zkp//8g8xw0ICt+mf/1u8Dgsz9XyKgNgAEImjxPQKY68Y2fSbe98vd9omPyA
GiI0Y51s7XPjJyw0l9Dv2mVGEgdVX1c0Wh1CKJQroR4mmuM/VayoWs5O3HMb/u9P
RRK/lEpBKildqwgUj8o5bEwHCywTu8K4FBHPgMc8GzAAPLN822vqfeF/fImvhE3O
LqJOJIS8pJ8AIXcLiM5frOR77miyxnzRTUfB2bIH7hyve0kP5MtiZ9kJCaOF0HGQ
WSZ8rMVsKEckhHgAaJvhzFUy9MK7DDeAHQuqiUgSzhblKTxf2FxJGOJooNOIRsi4
Kpkg4boPWpMZi6yfdiW8AYJLh1CHRT8pzncW03N8CY8Wj1TkMgW8hukbKEgO4nvq
z38sbmZPgiB5QH5G3rteKhWoOHBpR9hh2rfkDs7mbMEhctYwnKFYYbNtOD254yvY
TX3fbMZU8iwHNmZm7JQyidROOy7Dpj+nVYMi6e0IfTlorALDah6Slws+Jc+MIJdq
TpotGilEnuCCO6qGhMfauS0aIWjKMUPE8D29OlaD6fSBUhlm9wL5QopWDYsylRVK
2WDqU36m6KEERzG+sWHv7QbsbiJRuevhXvX3F3SXaTrq+chxGdd4v9A+EJtZvXW6
zTXbhBnHrHZM2UHSRIeiYSQGNAckxi8PByAMQo3gdlTj9mraODu62vxWcPQq4X0Z
7Hfv1DcPg2j3TQhd23aMW5IIQ3VTPO4S/qbv9YkYrbhzGO8F5UEgmp+siY8d56Oj
sOrBiC/MVKYLOQz+Ty/yF6vJPuEo+ukmQqcomNII9PHL2hVTGJqvifpRedyhrSEo
9ybu+/KqMpF4l4IA+nLBnr23feMv0mNYdn7GJuAR7U81iEJaspdAQQdJzgx8bw6P
dicxi8JHNF94Rcrs9Luads+mIbsurwGxlIBTYt3TCH9aDE02+YPdfwqWl/UKJy6f
RtdheQygphenOJKGEeodYE7UC9IpANWKwIjPHtshWY+W6BpFH9w6MUjcfjP63dbb
EQdNnljJikZdQiXqo05nGg0F7xjvmE5jcfiAvyzJVYr+4sQnmdIlkbR+C0wupH1M
87Dojy9qd+4wJ6dDOc4AIoK77sxD8aKTElZOo9RDXybcYSvRwjU70BAMUp0JzXsN
m0lryDiQpygoKchaijUVpO461wA5yAtSxcQ8lY9Rim2opeLwEGHOlFyLY+Zh8Tdu
HDSEieNgLGXD/h/9bEMKNZlXNudU6V75rZjVnBv5hCsK87UsZ5yLzFjFwijlrkwr
7mGXSyyHB+5HiH2+lJV7fxXwONIm7DDUvywXPbUOakOwsrthWG/Qw0pHROp2B3+H
67oyg33PJkHUbHo3EbRJrRg4Nz1WdkPdiv0wW9GyRQBO0Bkx+hcp5kqagZWFGOms
rHkjzaMaMEiv2DlV+LkeuCfuJJUYKQAN5/kMbMIPHFZb7BSgaZrP/E5fuqSUnKKn
YLrOnwWS3D3q+dB9L9M8CaWqgnOCA1CH9I/eAJccMcQuEsKRAUexJzGM5K0CkNWO
+2/WOVnaFNWC51NcuGoj/6XE1jWQw1Ow3P6+31R7FoyUlftijDd+raFE3xYdDFRl
pXOExzpab/W9W/iiPAetmHl4HG/LHqkhgaBDxjrh5JNvYMAaNNWIasb0bIuSLqrP
U2XbRI367lGROenP4TfkJ2BYGjCnOv6MRkmxRIZhKvPi2pyxRcCh1vjCti9IGZJV
YK5VM+A43gqA4wspOzXxth2Up+v3OadxTbWwO1lwrhb8L4+ASHw/U/SGlq8F9FCR
oFaRUx8gUpme8EnR7MR07IhgNtL5KIoN5tPqbda4dIYYgaQpZ4/3gnFLdxmAJrYi
q3G0oFb7vDhlMXqgS3p17c50oCpS2jYThffN/dlMkbs3C0XwCWEuOoHl0bnVfkDN
dCrRqNnjAX2McmyY72b4J8zW0eUe5DevdX9GhTmfeC6ByNnJHSEysEQlbemiB3Wv
Ni117n87jKFZ4DwBdfamDkE7Hu61oe4C1oadbQaDYC8l9kM6kvIl0c5cfer90i/E
IFfPZ/fuznMyH8LOvWVcUmB43LixEuF7ub7tPDsxij7goKeNRo1x+UlzUFDWdBB9
UYPMGk9l8eULbq++MZT7safS9eAXwRSlowcKYz9HG/b3hSr+XedPQhiZW5dEDaQZ
fN+0pqXSwe8w7Syr1X61hO2Sa5eQE3PR6Nzs2ZfOeUCFlMdLY0jX2z39rEeenXrU
X54A59vqlO+fNw5Lq4Wlsbw9PzWN3E0SQqa4cZ6sQ4dMUGWS6unXTrZo+dI3uSTg
CmSF+/Fx1aI0zz/tYmMx0RUOPwDES4apfdXfYwCNVN9x03dcCqrG2JAENp1ttF1B
JJeF7sg9haLjuDEUGlMp7wpfvE2wdW8+DrSIDHBKec/8meEDUgwV6Z5YvzHuglEb
74aLLqizMxr7NP51RDGrdYrj9c7jS1F+rhkPvVThkaJdSLMNcjaxhqWbX8dcc7Jg
nRAFrKTXZBbk2RQFAgLrypK5staXEIEYQCqL9eOjaVQCMQIvV3ECkW3vV9Ha8Jpz
Wg7ZbOKH1+yzyMgTUus9xs96/RxIV5RFDv20PThtxTWXbzn9nXGCrOpM3n/IOqPo
QFRF0rOWLzItYDQIr8NJaKe64chXwtbwDTe2JWRZGNVjaMYgZz8oBcxJ+NNU2kYg
7RSyBigLkLOa2U88mlxTJuYMHXC7YsJmPgzLtSod384SMzkQMUUQW/HE9ec73SPP
CKhjcJxPv14ga1aTwpmhbekUcaE17nOR7Uk9nlLiZ61XVb0uNjyVJ/ksBdVNTZao
YXhRl+T38XeHerhDD2MZDcfKEpl80LTitnKPYmHCnL8hBJnWlF1Fmt8IhsJCtnZz
4rwiM8MZq+kNbdHn1T0hSmMJUOYsoeBqaaX3TS9Yb+K94Sc1weX0KbqFSrw5PbMW
KpZgtf8YtkCMH0H63u7Uc3GirplXZ3Dt/7eBIaTgNUBaeSf4nj+vlHOS35ZkT9D7
Xuo6e+e4QEdJyttG0DXYV52FP3BWkwyymCWydTXxAdUBdBLWOP7ZtxhRFbxS7wPf
MRKxgJ+NsW8ei4KHs8SpgFX/4PROtU5GC3z3LOENlLnhRnnNT2gE/lAIsdNytrVj
UybTaD4zerZ3vO+T4Qp4+xMf73+0rB3au1fXmbicGBDj9oMNnFeCAzTzVGCAVeSk
JMxvPBPe/A5AJYUzUj6uD4tGPjBCkwsI81Sr1uFoX3Wb7Z5tyJFy+epQEpMk+6en
oMxLmrzxUtepwADr8s+/4jrYcn7WrxcQDdNF1/BJPXPbG53QkhSI7LuWxob2GCJy
WbbA8wpoXKo6qrivrHNy+7apEBt7M5T6OQpGnQ3s6Ua+yQvqXjswsf8uYy4cGjJl
aNA1OXOR9LiWTVj81XGKUvc9ndFhA43dZSzCB8K996n+8Qbi65Tja3D0OPgCgU63
yfisvSiwdy7BXPolTo8gryz8bi1Qoqv673h6PQlgCGQh8OdqgK7S2oE+j2FgH6jq
yGR+i/7QAuAFOyDSFuhcb8/WgFiJ4ZusPWtRLdqswz8xKEz14Ae1cEiYkBHg7H2R
+vfb9yPfC0omLb9tRxx2/DKO+Iwp4tH7m/86BHaYw73oc7ZVKIWQvojxs66dfAFv
es6jkBwi2Cr9hB7bOMfY25dhSq9VfmMuenyaBOdhSutX31+a3S+2bcu+KOoCLmr1
u/RHqgtpzlhj7mFgfUWk/Gs78lHkyHuaFAa3P3L6hkMuu5fV6xi4Cn4yDMU00O/6
0L7uB/OkS02JOY71XJberDsojaw6rA3m9xyOvQG/cExr6nSYmlG5D25GlR2ZCMt+
jf0bwFdjXqbU3bXeidLHQLXvWp06zvLd7nMxXesZGeG0AGDbooe0B8pzcIYafs0C
yjWzgNZK1enYM5z2so/eG3rK4x5ftX4dGPJ6AeKR7nNwpyxV/BmwUR7D0TBXMs0+
1nRm/3/YApKo/OWF2X6vykiPMDIWBdAUPsejX/UMqVi7tcxWDP3QeHw2fejNqwBr
MMYy/tur8evmT5BUbjo0gj6ZX2gXyJJ8dpM5bfF15RSIjVsP4IJSdjUR1ugeTAXa
Q3W1q7gVufCo030qcUCHKSP3yNx2wM8R9dmKSapjXdLJy6TMQf8DVJqvjMeh10+J
6tCaeY6mZjjGn1A0iX4Toi/iDvNqc7BdbztogqgmRTyy3JRuTQ4M6l5ihDBs0fVQ
BEWU5NsEr3j9HW1X/91Ue2uXD+KgQpZSaBrNwDgsLyh+PD2veFBNM0xRiwXLAELj
Lrd+MUASnZyMaHj3fvDD6WkwPW6qNzo3M82C2M23feFNGjGODaAHaha5eOUOTWKE
bLLCy1RYzSjUSDOOnnWn5/pEPmplEanYXb7++wGECWMhG37YIe6QZ4NkqA8u5rXM
ZrmTuo1DWrxKcDzWkU3tOIe5GYbzqB9uzr1ojo5dOSfQohrmA0JQWUVowPb2AmSx
e/bcGzSB797FABWPgRtcXA1oXM5Wz2jfZoA3UBXFDQSVJEY3dSdQ4zJ/7DHzyZJw
zX+MJgcccCLOfyQbO8gXBpspTUKT+Bfq2vX3NHO0u41NmNnhGixRl/jnbGADE6rW
CezRiimZxJ77p3z/0cBCx0cfjEqqYgsmNhOJUI1HrFLP7sSc1+uEgk5T/+vL9RCJ
Q1dde/1Pf4f85WhBfp3IzQ4VDMJj6Nekha80ApMUyXZX5XsetmiQL4qFk6gWmKoW
SRNKTQkSXCzj0bxU7aJdtBplukOpRRIoH5AhO9NiSqcCepo08s+PX720Tj6g2JXC
grr5RTRvv84+dZf48IbQZOCtZD7FUWc1CU1mHY117jiu1qzLCcR/q/zmQQzKGZWs
arxEP0wh6NqtVKmE7gmyw6aCItwk/x/QXKpq61GwoGX7Yw+KfEXk/pasZ0l8t7/8
H6gsBC8qV9kqVcYEN0DBbev84HvsoWUgvrA4fwUzxaStsxbsYtzF5N7bRi2hYWyx
Yf2IVCko7ZKufjxh4NlMCzmyy9D2uVZVnILFjq2I88P88ndorPDunLu7SmPyTO+k
mwXFIWLgP0hQEi8GiQ2S5+CudRzDe0kk3D6ReNNahkV/8fF6oiv/lWBRhcH9915l
RnZVcCQlUAnkh3oR2o4yLr3i/V7rvYFKmPQb3Wh1NMa6avUCp+ooVcjAddeJlV7E
9OiiGtYiRUEVx/61NWIDQll9e6zd1GpIVuS9uzq8zzvIOcxRZj1aSclg/8xJyWd/
Ahz8N4GM0h925XH3KjaKRrxXL1aeOC81yn/uwzTVakIcx7e6MRBdlOpV62omeG3A
lCMm5uPu4hIDANLYpkH/v0SphK55dFprA1+ohu0ChAWlZs52Ok1fzmcICZuy5Xap
B4FSyW5+qDBhFBDMbCGNV16Bj0yz7KWPj34j6vionspanYU8Ik1/bhMiLzgV+0iI
UTH6VfHUL6+dIvLTRv5UohXB/QwavqCYpKdPDZuOXNSd4tIngZxajVro9/FTveHd
ZL+C2FshH6kkXd/ZqZ4nKAmoJGJ9lG6/SUbSgKO4Hom0279C3KAPBM4uwepXaKSQ
3OT0p+964IEPDp8UbWWbMGNejBbcP0bFNWxKyOilRPRnFFwB++iW9VpfK4Pb/AFY
Voc2v6u7JQx4kYvdkEN9P17lv7yM9zoIlXwLRK9JGxZ0CemN05l5WC9ntVVX6yyA
yrkLcIASJGOURzu0hO2vNmNk65/eq65bni/NmmTTiMH6lERIDXAMGwSdbAcvN7sE
4mNunroBxD0V2TMo9xI2yDaABitTr88rNts072/ZgwHa+GAPWdmnwI+uNyH+ig42
Au1TQCaYUrjDfsv9l9qJ3PM0d6PyZhDbMkFYPzcz1qoalbAWjszetZMMSgG0AjVE
WAnRyRNWdOqdlAVFe+BTepNhIihpZDLzmUgyP7qtObeSboKLKB/GvEEBbAV4C/8b
uDE2MNElsNQyQHNd73xVMvGeuq4CAZskHdO+6pW5L7+Gk0kYACu1+J3Ts7yhBX8s
AiDTohXlpMgB0DS9IP5xBjbG4G/RHa3wZWJ2nGhgKFeh2293/JO8bQJ8s64p2PZa
UYegC4GWIwdTatYzgjDB75ihxlmkaBrUqp8D71oz79KghF03xZ6mQqiLIgV2Tuzf
eftuNlxi5pzeiH7omJ+SgTpgrMX0oHbPW452YGasSAxj30ovZMaatKI5giOu6TuM
DuNVnqhUngchTy79N/DFiKaOWn0IbuvYL7UcUIQBifSOWhwxdYjH1poXSFFEy1Ot
9Yd1rFGRn5OWA0Ige6FmJ+dxuwr58ZY/L43KAktbt5WzCh4Ur7Wy33z0MgXs4eAv
zQp06a+/dEGGoMUmA59fmj20fmeyMqFCsWr0XATPW4A2IhCglGSe/srLXRq8RUhm
BGFCduCCZaqZ1Lx/+HVo1Wnb39Hu29CG+gweB8/gWlQvOnukWB0OESyF7PNCCdMR
wUc0d+TJ5FRS3I2daTKsLnjfNsMYNev8h5IviSeD/tm6k+hMksSo+H/gkDTbqJmc
scN2PgDWZzl/zwPchcHHRn9IGlsTdXbWtVYvqxT9ANZm2XtWoZDQtdmmSu2YSlLH
3OfDm5S+GdRKtCguZQfdPgT0TZWjE3UXormz4Mfmjqz35BqexH9X9EaGj9NChAXP
LdrX66WSf5VNbg9fignLJ5POwuhPVuyjXOiiOB6WluOkIKuVmbYmaUC/dfqKhxlR
hK1EjcvXOi2+D4d6gSEXBpxDq5ZEfFUjyoTu2fhAXsYdR+MV357rC014nxSVUo11
3kzveLoHDE27pZhBgH7CnnmjFfxiE0gtNFFvyXOmi4eYhoecoa2H+YUiV+DgHe19
dSq9nFvSpagzT51GW6GMa6Qm5TgZyk8wk9OQRtThEFbzpgEvXg6554WK8WWRNl34
Zc1xVHc6xU1qpMNGrUHmysTJw5mxFKSY58qWIDCh+AF9bY3J6CouCaC2fC0IoT3i
E2mXbit1NKbrxqhTcF8eevKYJWOftKuqgBNVjptcL4Q+Y+NflJtLkzbKCkIlq0pL
eFyux99uxA6jGoEgcX8DSDlSpTGj1tTaugJ/Yeq3FzQIiaQlqnKgWcczwXYdr1uj
u+6FAyzCeJduDNic1gg+mUykDZTqYf8OemD+vVtKh6gZDJrr3cVRaNyyf33OWitd
RlIMD1vx9NgFLO0FArl2I3tdKcM+6oJH3O5crI5jxAgH4SzH8WWk80KElYXIgD5g
eS2S9CAfo/fzBZOpGSDs6yt//FjzUG2Ncd5HiMMbhs8jXuCfZLgD63f/pJ0K4Uhw
GWzV8MFhuuC5Xx1W2SOxqQ0PMQeid/B5/WZmxCjLLIkRRO7hoZiTdu6TVSJ8HnDd
2e6vv7o3+dyk5gOfwaQvKSkxCC9CYNckmKYKbgkwFmYTJs77M4kRstDiQT21zUFH
Frwf5j5uGSmb5t2yZMZgyJCiUjWg6qhuXLKQNFVLc9bbxUy/gPUI4FhQtWo8Xqi/
hwLD4+GjzO2ki3cN+51j53TZ8BlZDDk+Sce6uKGuRGDEF4T07csVHIyT45g+D8Ds
bpduCajDixsMfUqX/aFPdrxG1eGKb/njGuxAGMMDGgu6drQduKy7xTOippfM6YPi
TKMmqWvoBwDNLPAIulODMUdoMq0wRC4AKrG/isMBgWbdH0J8G2+qcHDh5TDkqPM+
nHLOtic8WWr0SBiMUq6w/XoIiqQNw2nDPS6K8k0lAZ4wOdf2I4MTxWbO9TP3UDbZ
L+inByOVy6IoGY60yVE/GY7wE2Z1b2Y+Rb/6uUWSXc88qZgx+FoWZp9nUi24SdbY
ZGDVQ/iCi2MOi8wJxVtahOEl+kc4dWE977Pvbtv1pcJljUtsJRGJy4s87Mc562lS
V34sN9BkRq5092z0vk9wno88NbEvgj1llDs8eP4H2X7p/P5zmfni2DyuDxnuy+EH
qkad3pSaQOQUPaXEJWEXoLqfATjExZ5nLKMkVq0WAcTVcEccXomkI6B4WnRMYluP
lBBdwMH8QhFhpfiubZeNL8rUhBn0cJpdZF3zosUzlF6IhSMrX9MpO39lSgy05Lew
EEOwhMdL8+t87kBXx7Ocr3O2KkuHWxoMWJhGtmec6YnDRh2aNN47qOj8rL5Z3zub
V9ie1vpcMImW5J7vd/090Ysu0ATUfSO7F71aoDhk+2Eeepaq+KPW0uCeg+eH2rlc
1ArgE0eOQLA3xlu6ntOusG5cbCUO4JyVpve5Z53LXfJJ889kNpNcTYYvV0KmTLQv
2plt81x9rdlnZoZ/mfz0+OxIdQUEsj+HYlBAaDjJMM4MQj+7TaMdo3hQZSssdhZf
wwQURbi63TGfEGxVibhAgrlpRwgqCxJLgnDyWbf6K9KTI7awnoQNgbaUBr5ATcR6
Jpc2xPIcqS+aDlU+7KDVJhrLjbZ7WbqRHjoKmipyaG0+3WfEqwoJDjurEKL6gMta
l3x4DDGpXUmmKVpVDqQYQJz6Y08aP8n7wPnsZpLaqpLk9IEC0LIJgFWa0neaUtHr
7u5b8t/olilSpWIKa7D8xyTQWR0V889QfNCr9CPcutBnw9VMWngn2cjY9WgZrQLB
Gbt3S597KQXaMlTpCyCCOQU4QUfqq4LJOeoDNNjKUqRV+UNURrpDNq+sVyNpT8eb
A1PecctIZtFcSq9fYBSSC479FPbrvnjOD+Mu7oBkkLGKIxr5o74vajOhzWEF3MCD
GXErC/BYwbJvNeUKiECy4t1zNmI0xT3RlxGMxI1Ovx5a3t48kAMrPcpE+dlTvcuS
084i8mBsxyW1TLzS8UzpcwDCHcD8uls2BbM5jXNFZXVt1TVrQ/Da1rL+eQ+R1CML
SSIBG9EzDzJ3x4m0s8/3P3cLPwGAW5YZDsVFSVYPXiK5kYgX+mHb3NbSnFg8say5
BwcudwT7eqOuXc7vvLceCPNGIU1XJuH7AtRf065GgIbKt0VjUhMIixJ7hwzryVx3
OTCfx09JBnB/hjBYMSrYCLR4v+Jpj3nD3Y9YMcsXR8CSSjJDRDPzCpNnWCmpx2QU
ma9qmAWIu1WF5zIJpwzjbDRXXjMcJ91DcmJQNtBiHb1YW31ZRQVZCrAv9p+D5b4t
BWZfZGUZpKjXIXc8eGANtWjSnOmAAX+JXIwLKkYAgbTcDjSCSD6A0PX9mj3cfB19
iXa1KbJ0L6eqLf2qYFcIiz2t+sOfQ1gIueJEKxeCPEWlSEr1K10bqZMzDU0o7dbG
IZSL29qRRKh6aCEbc4iWIgKNCg0U0plrmADfbplhUqCEwQf4hUWrlAXkk9Umm6Xb
4hrXL9nXjbXsOTj25i5PPApSeXiCYGl+l8lcdcNuirQSLGtsXjL0vVTV8+H8pJKf
e3w2iMYDhghf3XC64tnKG3EPcs18hP4IzhhRi6NdkxvHOypb5WoPg/wTBsbHhb/m
ohhpjmjKiD932JJQJ+BkVi9FXE7l9bBv17wk9bk3mW103JGi32fGwuch9brM3CIo
+VkX/K2Ee1wGSrd25eqDOEf35ZTxen++Bz+Stl9CiP4OddCSrgV+k/uUE5SYMeLG
5VgcnLxOxlKG8RJmrDESO3SpETLVcKxVxKFWCvM5CAnC3SBNlMpwAgT2vSzy+cUI
eVsc3JTee/h3ijFTUAwqWO5fmSgtTzEEeF2F4mE0m50sA6UTwcgrrLk42psvRbUz
LdhsTsy7PVplJ1pgngnHqwg2Vgwg//UmbCZMplVSwQO78JWk0OKSt//QJriqHqPH
k0hqS44ghXOuM8y15a/6zDNHfAtVebDhcDR0IWwcblYTrHYAIPCRBvIcXJz1ebbD
Fx1KD2+YP+HK9Jr8Cv2IFijgsI2b0bNk0/gg/iELJnPC0JJ89TxeIY46wmrRD9tD
tkYA+fR24oAvAH999uvsKJjttLI87PmXWbiZLe6+H3qTKMD1JR+z+SBiY4VRnisK
gceIvpjfZgP3ZxbIQtLq82MXqWYBbOddZl2JhTKwg+ds5j/p4U4NJKvLyRKbiBaG
XrB2qp46vKJ8QPDSfpwtWROb3H0i5etAzCn/m97vL2e4qDeC54xSg9bXMK3hHgTU
mIJ8q7kvpc30lC18LsWhGsDm5ai41EQfTt9neFq9mmSnwzDPsEHoNRbjM3RlmhDR
Im5w0VZAFsjzlEOTxUug2erZiGFrxxxikcSy406S9e6T8DKBJONuMl0aaLS4SMHs
Tava5FDoe0aoPpYGM5VC5XqFgWjtYgW7+qJ2NBr3vrsNfbr4YqqxLD+KX39tZFnh
obH6x4WUjMT//gQEurFk+9LcSPvfZKH054n7ALCtQHNEHzZmKeEf9QxQc6Np+FsX
VqGZRYwplVCagJUS74X0reGJ8a1ri7RW03Y27+6OlDj3A2NqO12DgPL9sAU6eJTr
g8fE4SKkPYP/2MdScJ3jpPVAF27ljQK+HtoLohuG3fZuyP8oM11eryS5QmgS1N/2
Bwz40ZRcY6XqyPeOs+SzGBOyJi6SDsfus4XFFO5u16EUBDruoTCKVCussUriAaxe
j6Y5fZVyi0OtWI0WXHgcspeuEM9wPgbja7jGjm1OFLjK2TKgjRuQpfbsQY5cjQcA
wf96zpqAIpI7f+kL/fMi7TGhQkEC2On6SE3vWbi1lAEiB7Mhwz9sFLkBUI+4K7LV
DAy4SB/Jd7F4z6mIbaWWKUOJWvJwEG9968o27w5GsG6xwTHDC4YtO181oZhjtIK4
RKuJo7aX+QB/kqxsg/2+PL3qIjMiy+hSXcuu/Pb16gkK6By3gpZs3J4BU1MtcHV9
6ZMkxC9qp6Kh+PQTZ34jzbUJbD7jtMUNDBt4jigvRhd9F4jrNVjyoNOXZetLXrMo
VItkbJJ8ZLXjooTfBeCWotlfpvbBTkf7yTseeFYzO3hLS7LD6JwFsqrVRmvWdhsZ
uzlUtGQqbeYba80P2xj9oW9M/J5WZ9yEH0ZxXcLZGoFHwSkqJo5SjNm62WngiUUm
TxDPIDDX2OTA72GdADrBZammrMotyt5ivGmix0XDh2R2+52SIpaEGkZ1xWyabQu7
dx77OU+xI9R1ZzUokV73TbzPGc/XWIDbbDqB6uraBbdg71OUeBV6DQ1zvRt0B8D4
CP+FW8BzBekaWHc3oihNzp5LG2VYI6e/hFFWDDPBoONivYP3OK8Qm7/RsZRyl+os
tXAWw0k1uTBxbrfmDVDCbUT7YXp9zCwpJ5+gUEyK/QiFuVP7kdmNNYsrE4ujR5P7
zo/l5Z57aXrzlVSAhUlCXDbFACLhgs4zpXpd01etu0y3tT3sM5Mms0FzEYX7x4YZ
+Se4+A1eI+n4freSSsoT2ztCq1dEp0CRRJbSmyvkBvFuAcGNv6dX6l9CSSD4MOSF
y+8TDWyJXf9BeFUiqLUm2F0NGBA2I1U7LV1phJk3GyptwTqWfECm9dg851tkV3qj
JifEuA/v38aVNYv8d35a511DFIuqvrT+lo9bJB+9ickfR3pUrrY9/TTnKI39kpSw
/G2E70TDlmFATeAlBy8TRt2YFH8/BRIjBDxovTcW37mF96HJDzpzsPfC6a6cm2Jx
+jqn0Ul+ZtJjfFPnjdS9IPgKD6lF5Rcjq5XH1lg8cRv+Mo1vB3mylZcBz3zZYtwE
IHpj0sRR6Me2KdCl3Jm6co1ayqwN41HtZSa78fxKFRbQOJX5DWbp0+RD/k9cpGQH
iozfNJxH8YV0p3BhFgktqZZiAcpR3rXduI27l5usTnOuHD6tYoPgCWMGLfiifIEj
O5pVEQet1XzWvjhl07JqNswfGUoekag+gWbysdxqaowG3ntjizwHSRU3lUHAqgfG
tnOVHL//2h/uotOOXNv4FQhe3aXHuKnhVR3oxz29EUlWzokB/zmRECTdY1mqkyja
UFBbTxANrj85di60CwOztSVFACrVYlKwLjyCqHfGmk58wAHnvl446ZH/VZF6T1hc
QGwJW4KlgtcugdBswYPP+z6+uxWltOUp7iQIqr0YM0TV7iw9OVmyBzgHSPnxx8n4
UvuwYRJawq3ve/qc4a3kvdm6FfkEQ5STSzI70Tb3N4+KZmbqLRjh1P8/XEoG6avA
bJe71gq6eD34hUqCPwrVeojNa/H1P40P1WUENkh2J1Z03DqNOr7xud5UZ7GUJkfJ
pMPy+aiyMXOkj+873MnQSxQ/KtaMcQtGMhS+ccDDpREkWDdHKdGHFPp9S3qI1vw7
EgOwYHArV49PLR550FGW6756Ndowsz+swJy5fN5sF/CF5Q5y5qbCZtkalCkxnOQu
BLFPg1wGrnlOLO0eKrxsYY5plYRILJGO6i+oCAd8NyfCpyEm5H7SaNLz2xkLl8nf
6ALCJvrLI0v+i7bmX/0HdLT3dwI+7ig+z+beNyJAD2S1RasXBxrtmisBfTNvH0yW
MFI+LrzP9lLR3elgzUaKiVwiHS66xBllkb3rP/xznBC7cAq8mByUbU6eDsroXq3i
+NxnZUyChg3ng0eo0i9Q1OMeT4QXeDVd8bI0PQSJwlNJNKTQ5M8QLVQP5rEHp8nv
n2B3wOZLgoJjc2zOVthaVCyFZJCDPFSpO77uVTzXmwMJuLaHp2hjsTxEQ949NMKO
IEoTdhhUOAJUq62Pq+iqf8cvxEgjQIsB/AY9wOQcQl08/EIVGampwqczB7eSBrL2
KJXcpPNc5K4GUKqR1f/Ij4OOLJ2w47bk47wjF1wvJrDuaHbgK3CqNK0SS1mn/QkW
8erY76+fzR5eOFPfSZYB8SL1otn7lZSe302ysNwICi4EqIaCNy6O0w4iEwRE1ZAu
/+F6T9L7ObttOwnMDt1OsaPXqRMdpPCcZlpZ2dE+HikZApz8EbBxF31b+TCa+18Z
m+Yi3mCwV+rLxqsOzmHDht8xZWLVnYegjOHfyd2+2ufknQSaiJqb9IRcGvdmBFP/
HqU/oWLaq7xX3ocsskwhv3vb09vWDOMI095ti0Pt3+OlqMk9hz+cym54ddgIWEW/
Y8RDiR33Xl/9y9s0bteRVSgH3vMBgAvJrvTESIyaYYmGx75aZuy4zJkP0sigu+qP
JJhH9LY43e3ZG5WE36yO1T4JpguMKq/V8vfFoAN0TvQHHnjfkdb5PZv7zIuASzJa
B5QztEb8lxPj0Ccv2cFM4+5pptlAh5qubouI9g9YjqKOgS3Y537i7Wih/zE9hfN9
4ZQ4zk14tsi+eFX1od36FS7xVcua69pgzDwrCOiuEbtlLyIa4scDeqC2JfS1dlnz
KraakNkzl6u6LeqXxX4j1LMcq/3luL0wGVBv5obx3d05m7WqO8xbmlQaMb5btHbs
GoxnGc5d0xEXq1/Is5fsdxswJQt8mKz8HLm/5FEMnklnp75Dx1hL6cqZNZA7jTAJ
ucHoHfuposd/McwDwXn1KS9bNq9I8WDIxf9mBXZA87SySQQcbXEYlkFognsY6jZg
VhUKTdAR7zXD5Povc1HjQB6iA6O1Rr57ARY1k33LayIfHmwBQd70UXSz1A0PQfcA
Id23RKVM7zWgNqjzg8bTD569dHYPhJk3dUtPDVVYGthU6eHQKpsckrHGKPgI/cCG
7RjhlFiL8hNq8TIXdZTLkNqYf6QEzXkS8/P9OSKM483a9nH08X9syoXRxCkfTExy
8R6YVWgOJJlJxZHsihdoNIDXvy/72RlsTPinUxQ30ll/JxpNfPjYql52XTbFAv5h
TzE82dQ040l7slKq6//Ne6h6dl5lQ3Ogi0h55+9rVptweGZfFMezk8efEt+epA4r
XypEtBJDWY+90BHSPCnX0GuPJZvFxCMKBNkqQyFBK3PVySTdMiEeZQ9Phcyjmu61
6W4volgM68N8bIBYAlgS6Vmm1Isp1+BuFLywzSs8a+hFiGbVVjUmXLV4klBFj2IX
ZX4+GCNzNbQRqczIJk7+sdCpyjjt4b6bbrNikHFJ7HcXIqEXEF0QuMrTiDgSMKGb
T4eyz9L2/AbrREiLt8ORGqGlPZaqjTxQK37MF7wq4VIKyjwWhWzsteFc5LqvSdeg
cDsGrdIL+Fb/ME635+vSfOxNzUijMOAAVLFO40lZaEYttxQ83Fes1T1juB6h2PvX
PMJLqpXxqVYl6Cxpb2gRpxJUZHiUeDadGvTr4AvnDd+nugzdVu6kX5qRS/YRosKy
gFLS744xu/6F8C+E9k8g9ARnwojidbKUFpcLsvWWDVX2QBYmcdaZhHr0a5ldzxJp
dj9QqGdTzr6bYel0y2jCIwK4T8T2Siin4ypFTpkOgZoqBMMtTZrWNkvxH7RwM9Ip
OfUSva4zHeUtODYcTjGHLkmJJfFiNSLnVxJn60GvjcmuBvsbfvTfkooSv7PLfU52
T2uPXGk/FcixldalB/F1YUOM7LroNy2NgmbisBl+B3q7OMz4og5vBnGpdiRvnD7m
YTAF4DFh5+jbQDOT9dX7QQ37uNeiCww67RK/qZ8PIghYfbD1q02sntfEhRVrAAF3
6+MU2r95xkKrF3z4SeqfWdyv/Pge6DfiDIVPDWzapVkO+YysdzIGeJZKwtz7dJMG
IuQ2IGk/reY2OXpqkMTzod4v320hemPCDzi9rZqxa0UeCgJVlAJde/qz0n4mE7HB
pi88X12ky8NItweztMDaqlRjWXjZl0Hm3w9GvvWAUHV8JKuFrukYUHHRI2/eG/xP
0NR/GhmFCxbD1z3inHUnoHizphQk+ExRCZdoPigoQHl7DNlgWb5soh2xVcneMyJD
jkFMc7y6JVX7TkslIQc+2Kg6fJhNdeOdVcc4dqDJWMVJLRmQSnZKqjbbXQFt0piy
F+5R7VWXwyJxCIqlwo0wrBv1AriF4RUydyq3QDpPvZQe/u4rJLWedN76K6mHMa1F
DUOb73TpYdFyBrORyAG9UkCSfQ91ylMmujkCstAr5OHS1QpVyybSNQVYkzS0aHeH
/dZnE8XjQgEa2Fs4F1b9APJNLsYeOyTsRC9/axyjciSfFS2Q2vrQG7jSz+kCzxu+
2VRm8JaiA0UrQIR4mn5y2HtByXulPvyWbkO2tjKxauCVgYYzaN7Ymrf05iS5yAEc
flV/ZZqCArHJh2MxETbTD+4NvG9tB/VEm+/l827pm5c65xg1Z4EbRBRjW2vGcmU0
5olkUGmRoAAzTRbwDYAdQWIXNyEHOaV2MHvGoKV92EBWcyo+g1L9tVxZI2SDIoRI
32zphR9NiNTDwC9gvXDb9WfkJ0P5uWYP4KjfhxgmsgZO+D91P1Zbi62LZMWeVfAN
XB8yAUS0TnEDNV9W7mcyFucpk2N7ULQhjTAdFjoQFf3WEzouu0ZA4T+Br03dhAMd
qD4enV6Wjrwj5qgpqGnLo/PMkC8HV3SKto4m+gXYKihrY8V9WHiCEx2doHd8btfN
PTfZoaHuffe645D40JDINWO4hfXSmh97f+Sk3ezIPgPlDc11W9vMToqLtTMPr6dF
G/AaqeelYqQhFgKMqdP6yUJOnWMtngfWQzR9fR6/Rkphva4aBh/gvBjFaMAGoPNN
Im7NjVp/4AR6ShPeZ6Wqke/PVzg0R6b2Ad50mIHLIO6YhgavlaBXhrE/6UXLVUfw
Hm/eVzk9IBmv/Ab1YVPJJEkB8+N6cFey5LtFkdMtaffUvqYpbsDLr6A3t/z6C6YA
Gs+Vs4SmvYnXGVVb3oLkAcI3rjbrT0zXYGZvYH9E6qMAXPx+5fsgO9qdb21kShlQ
F2WPjvN2lnQW0/uM85SaZd/DO7ndv+fJ+koDJ6LZqe/E0+F7gBhvSP7b6d+5bi+l
vobDxucmBC7/+GkRgF/lDUaUyYFvxRcDgpNvJTL+W4cos27tDLOg7od+NR0MApd9
rQP1eUBzumytn02d/Kvqa4murna8Npy7Xfwt8T/xzDe0K/O4PTxDPFhXmK5vjyHc
WuWqtuzD1fLj24Yw/wabzVmRmVhaZ5qO7NZUL1qmNK9FSas5WIsk6pcV74dk0BID
qjz4y0tvut/3vu4HUQCFhld5yE0lcyZrBAyjmWpReohEZc9DxuzrVw7YAcRwHz2T
6kMsCp9tmVr5wI9yozVLLBxFKYtwrFeQI3DnC07K1auh30Ian/5eJF468IbtGeQa
Sh9ax0vC3gaBZdoeoy7TOkMm/phKR9VSclBw4PF4JnxuvW2/n9G8uk67t1M4Npbk
K8/O5RjTDLd3nuzzwuzZmcTUKnLIyilw5qGqui3DSHtymXP8bgOaIPuGrZbOVuAI
rIn5T13StU+oBHeY4XC1mt1px/kR5mHTcn1AYbmOsTGvZqS/zEIkROtHpq9oDdY/
kL5Zc7oVmuzoTdACke58Q6aYeYIvWLm5M/N1m2hw6S8hegSyIRlhHkc3cHdBhVRP
fSOsPTvJSnDpaDxisdK1BzmPj8bOJj88uDEaJeaILD7OIpnzgUORRrUmR6EvdYWv
qBkhJ2RaSf3fdCBoPUjzVR0DfHQYXIAxDvnAi/8fGJlGKc5HMs4nN9/Xjz13S2Re
KT+BzgqK7iI7P92YuVWO5+xk4+8p6+atBRcOMsawFUwo0Uq0oQ46i+qd4UGXe6Ck
o24F2lQ5KWLyzN+pHqlr8vkqLNS9MIjjk5Gld+kR9fMhLxBrh2CR7KHHxyKOGuuJ
VySrGSlfReEUlGA4wMY8ZZwbWDUWQQfUVl1OO0UzapNIGeLcE8drWa5AW/sW/2Ga
PaKzyBI+XecRWnB4h04AbHk7297cuq0Miw9DHAKc9ezuyBLrVY9jKCpcCsoi8P5j
lPUk1BsJVIOokID42MoaGws5fdCn7/ZqH29a/prJiyezP8Vt1OHjtaNlAG60VdkU
eqVRFv54IYjtheHYvuY0E/gP/K9uyVngAvI3CeAaIM+XwHPf/imWHarE8QPIJbij
RTq9hfriz82JJqSPoZld415mdlR4nfk82iMn2I2rDN0YoJCsFK+o34goBUsVjR1T
mDv3zIR81aT0eefdIjSIqvE2C4bB7UhDAwx7fXIfV4ZUvor2URJl7yw7vurr0Hd/
psGgnvjM+ZZo4/NaDl59bPLt8xtlcRV1F9aQUNsQvH7PSAoJBLdga0X+F8VYAhj/
C8ndUiamfPUxG9G77eAHO/yIqaYBCABgo5FyOfM0aXGDtqh3rCGXfvHCE9ucEviw
wpLC9CidmO1SrLBiWygbtbD066Tqf3JDMO04UZ0NQeDw5a+rtCMUeK3bcuW9SrLf
ClOWgsxkmj6BKVhJGPr+oE1GFqQ0VemNXBrghhZnJpJcdO6YqP466n5qEzElyEBP
NTAlxqyC+CVPsb9W513hUShlqPjarL1ReE2kXEXQomKBddcdhyjC5yqJMNgFy/t1
dlUu03o+0NomhZ+RyCMnnxrpFZ0PqqUN29wFkXYK8Z//qo1jYZFt9uLoWDNI5gEV
NtS87jTvuOnV7sYdG+rrLXr4ESKrh+SsVJxasmYzBR9UDRazjnWjX8Rk5AKlKgrj
Y4EgIf2LrdfjLnNRNLEEahEvjLKQZ4XLMusgF6nfKJ/phdvm7lKPTGt63FkG0/z/
BHMzTxRAvdZZ6WbRr1e19pfuVLd1ZV4UjbOZErrKn0THrjk8WeHh7gdozNw4d6re
WhokR54oBEjv/wpaO1L7TAt8ERMPRm98nKNZgJ+wt7RgEqwduuOOsBueIssEIMsc
S8NxfG1ezdcCUUaUJHKYOOEwwjx7f2iGQ7QG1yXyEhBzPB5awhnLID427nzLiKVc
T+K7jpjFF0kb6NY4pV2wi+YN/CROsWb37O7K5uOwHmaj3C7gUOC8zLaHUuLyoa8e
6j8qG6WthLTFJ3/rb1gSx5ubxv3CViSV46Ves4Es32sdhjHfPsZxgRhbmGW8Ab7z
8YYH9zbZsEEU7WZZCB1d3U0sWgmOr5DFZcR5NhI5rXvmkwJ4Rj20MQ1J1uGYS8me
Y6rgcCE0ajNCf8bIDnmCwzd2GPs4uZX3Imv4U1XA56fPC+HzOnGh733RRrGLzn++
ywr+7TXdEBfQZXNrcNMbb3awQcZwvT5K0qhecLNQx6whFTnHRp/gzsUaKPrg3Q8h
kUp78JbcsdQr47AwP/nGCBs/6Apei+8wgFhCsbWMTJmyXYIsIT+utBM+VxsOWOT1
1GPjk9ak2pZgaENeqR9Qz8BQodGZ/F9fYRRAytY9J608QMjyrXdojZx0TWNdblN2
bUf4WlaLJrVzd0sM/sBsaoxdkWsJsu0FcB2ZhprqCgjRQcTfUXjaEGiylD21x4NO
zWGeouQXsDHVb0Iu4LoicrZb9EWsfOdDm+fgK/kJpgfL7Wh0SliR6jDcUF2VMLNi
vwBB6jqKBiSWHJMbDLPT0q/mSfzcqXdv7BCXqtaLNGbQeuH0h3IVMhCwYi5mxVLT
gQuD7/h1C5L71DqDNfEgofjqC/L3NJvykcRFMXANVrpxVPOCzlJlhHgJgiLZTq0Z
Jl9+vr68Eq8TDAY77mo7BBIYbtKmbiEUkUDi915+7h8aCNNeStFpGBM9wWjkNi80
RqRMl3Zybj1H134qG2dB2tKlydUlpWK7eQhk6vCs+TlN8P5+/YZpf0UNkAlGabcl
Co9mn+fBtA0YTpX/cyNc+ggytI5GLcSu7vBjz+cRky9xsPoGtV/dvceT7ajOJAQw
4sOC37SJhRuvvZIndEXCGSNxGQgn9hQYKuqstKe4XP4ybz4wK/gS+SjoJ5Ioui8e
NI/QGKWHSjSxmeJhhBusOY16IL5QlYfm8WFk/cRfYW68kdmYmoZyMnXpAWbrhTyN
3Z+23e7HIZ2Wo9fXGdsOlViPQ5t+zpqjRaLKAApFJP9/A2JiMbRXisYg8/iAf5Rw
RQi2WpaUOX/tfEP5hq4MnLlwEseB/ismBaie7kLVF7eKFn1Ea2J2tOJ3M4ZLGKKS
1PBWx9c1I5+R1C8UdMw7tuk6qf7hmP2ZY6nZL7cd8sCV1DGNCR5dGj7nJJiusbq2
K4ZLwyHKuTo3jfVw9ObR7jabevNWLwWLhjKtLmcKb7RwDfUgaswfn9FckvD0Wnoo
QFCUCZSee/a3QjvhySJxu1mIi4GYnp+v8nNWi9JhlDMHPOhLlzzBbS8dak1HS38d
AsHK56aRn8uW+k6Sey88W1iFbk8Ogz57SGzDnQjy5qoDjRDOzQg9JIL1Rx0IVlp6
6RS3PlRXB3DyzATVpzT+7XsofkGfdcTQES3YOtRGw0y+R2b3mlmrNTblxxctZViD
a/zx5K9B3jON1aQO0wSLELFWemkLSkc0bXDNxi8QVtvR8hoaIr6S+4CHyapqs7Lu
wKh8m9BXhjZE4imCKai1gbIP1jVEZ4XV8f0hyXOzxuERyfnFWPqu/pE9o+dURhci
aLBo90exACKygQEBCjTc9GBUFxQdMhRchiR+75okWmNDQYjBxDNbvP3NH7sU3afP
eOn4ytNaHaY2ecaHyItb613RjIGWhAkayHfIB9kWnNFSxP2aqiOuN5hwXgH2FcoM
HELxoEWc+M3UKQ0O9cRfBxZwDPOwctadQqDoMgMjEWclmcBe99ftLN5Dy8RyCk12
qp071lUXbNPCYfpSMczm0GeN9jYOLAZRUBV/9j8mUx6mXlNmFDtPuFw+He5BYSNI
OZ/Vm5AwtfHJVcHOc+PMTK9YUw9lWy3KEu5JqU3cSAItQD6IR+lNzhKAknn6HLrA
Kc6MBWF1/TbrJGUbCFblktriXP+syns6JHe8pY8rC9IDrVwj8Ng0sJlN75j8nQv3
h83/tD01/yTu20rURpUXMO3foY0sD+HgBfscpy5gpCqtgumdyCUZaCdet3g/Gz3a
JT7m+SLn+alKGm5GRQyTrDXHHIHo0X9SqfT/txiN1v8GrHEr3hVI+F8TWEB9Ygwd
LkHsFPoEajVBIl9RT2gHHlwyyeLkXoKAdfRcMd9mnIfNmB1R0BFF5scWXLO3f8db
kzQOmbNDrHV8AXgz/cjz5Cmiw25uivrLFC6Vyfmobi1EITLZ4NuyQcCdHswLP2aP
7gB5wY3KG8I2LRE4g2KvXl9AmCcWGJpwMQDLKCAlB7c+1lrsaoagogKTaKsJ2hhb
XCkiR7X1Q/limroc51AThv2ae5ymxXEdlIWtuBqAxCkDjMFc73Tq1ykxE4ynx7Mi
zdK2RSoXrtWH43KC/Cj1LcXAahmfzG/N8BmzpH1OxT8giA4uA4Tt7lgwq8QiAxq8
e8D3xTukl7IDxRcpmSTuAT3aErbA3fWLMPyvD8kKDG3RZ2eXLPY3zoNKphpxs/sv
G9wUwwxcifSs6Z7Q9iJsiDw7VkgGUhJMe3GQF0aMgCzaaRU/IYSnXym9lZ4J5d8Y
Bot7tcdQorqJeWGPl38bgiqnw3MjQr5DDjhuSigKZpLxGNLJtbEtSYRY+/+71ahU
uH+C/hqHvOXZln3MXGTiJ4/nXlOTZFoY8ut2bzq2aXu7xKjXpasrJZcMgtz9BISQ
1d2aDxZvGdLSnrcZlA0txI6xEe/TuwBIxgUV3GCvPfKvaBmRwpaEsjfHzUp1SOQV
DQX1uMqa/OFuNea5miEQYjwmHpZ52E2Zlof+/TmKn1bCNwnF8bNTuz4/7CGpO054
HJJ6P1nXqJDifRqikhDBdrpsog6mZv165+8VJCooGPyu5ESZ31nw2L/CAUM3mcCf
svxVnfG3ItehQloB3lPclf88KIQBqlv/9zSWYTEYQ2njd7B6fFk/BY+RnllutIUi
THlZbH3rKNO9yghowcxh7q27HFnb/ZkaExX0GahTUSoCT69nbhuiMb8HciXk10on
YQKvC8fAZmfdNQ+xFrCzACv1cnyJokIzMaJk/sXWos9XQlPRT6G1FPrz2Raro1kh
tX9EJxwZrbELtv+BvpmwoSJYxXRDl0s8LnnU5WyIpcoZWeNefqrjl3DGEmSGbH/z
QrmDLtQAstELV+4ypkvzkhhZm014I75Am29qXg7k98FreJNnSmlm8uNcQi+jq4hl
SKXH5BZqRY/2tW/qoB5mcxaIFt2sPsjsT1ldzIaKI8OG2dWx9Zb2E5hcB32CI7Le
7sZ1EoeFpfQZAMiNWEp3DlUWWsUFCDDqZp3JNXCM4G3p0GPSDqHdv7zJKS18giAR
b75zTgywvw8XUteVGklWwDwq8ztdc7A7dYZz1vFi8yFgoT+2m+rThEDcwBpSW+1S
184Z309CEjT6W2tXiFh3BsjTDIxA4rJhKTvSCwls97jMAle2bUkeuqHAQ9FUZQ1h
ARGThuNYca+MNzVMX6R2hX7bmwGtamtmFVd5RetyEOqBsU2NoVBJCpxVLzATTDhF
qRI/JfgZ/PXCYFiMnJ75Xw97PuLhLNtv9GgenrAYKC+28iwuyymfpFefEVZNKZwd
M2XR+0i8vqQYb2DKGDyV7GBfKKm0tvvnZhdSbY3lb6q76sjvwBKIvRfRSCG9nxGv
V7l8BVsEVIi0rmfSd71yoMf83g1o9CW5UmyfGeWavzUupIll2Hkyfn4CoOCkjW91
UmvWEhyeufOEqZL3+LGd4AdXNz43t6o8CHudhdE4o5ZC3phXzf/C1LFRNvap7TX7
59dZQ30hT5goP285R9kFAAPkN8UqIsoWiKPM6kJ0hCfpAJfd6PfpFZzIfT408l7g
tjrF5XuUsNdgPEQR1Icxqp6oKv589F1+M16IfZXdSmdJj1KaxTW3ScZgtp+evRgC
zxe6y9zgdwXLryohG4vXhoiCSln9f/wPLvu4f6Q5bycChYq/yRUP8V9H+A62039A
TnC3rSE9r+pe9pHmc2Y3m8XAS5gT84x8MYmKjvO6NDYn0oIdfTD6lFkvpvik21P3
VqiYnIBn1lLym2/qsu5iEPiVxzvYwkvWpd3XeGTJfFUlMoQGSOeMdLFh/A/MipjC
vMSkx+NN+QONKMfGDK1Njc6iG7ebV9z1euRIa8RIM160L4SJ/0dCgzvEVjkZP/9x
VI+8r0JWnPfVo7vybxUR9tLe1rYZ1jejMFWxzj3DWNkEH8w4cpjpD4UJWPZNhxea
0FMCFpR/k6wbi2Sk6RHoQrMAoDa7gAxsW22gaxk+sToLTrjuF+o6i6Uxh8xSSWGR
Vh1+FAK7vHWwN1JGwQbHJRzD4G8mBX3aqHPWoXLI3PCW1esUsrk76j/z+3xLgPGV
ICocdvzt0ZXEg+qMJZ8/8v/uh2kUZ5weixWy++1/mCx0c4seMxS35plfA7f1ORex
zFKNKM+fAyEiLS4ehFinu6LEdMMBliuFY2KOjgU4xtRxQA1TR3pEHrEIphgJoAQK
XrqiRhP3KFsGu+084X/BCvwrm8/Hi+U5oAYAL0KuGHr1vCWGvISK5sD4ZoChWzI8
iKPgW5H0EGUmzlPpt8RGBxAADlqdGeUWd+X8BV8vtU7xgTw5LtorpIuXUQKHh/2+
J3y3LcPQnTAieyFoVQGSlasaNdUo+5RgOvqy+EKyObvvxnOZLv7yzaLNXXAcCWZx
5w+5WU/Wb/no8T55aGqpbLtCMSooAwipb6HMbNB3b31TL+anafemKui65zWBczhn
NIMUYaiT3NWrKUWL6QyHXFXA6NKBdZMpOqwkasXsmDULky9xwQFwePRqgXWKqE/1
Ufwho9fsrTVkUVcKKSmE/NhYHM9VCeLh38hKe2+zRrT0IDsGUGsNK8AHB3bntUYI
rNu5OwcQ9bLqqUdD3vAu5/UNbYLWxMlIoZrsQuw+0s/FPz7zo8t6dT60ndyUxngB
AjLH+XDrLlrQeZA+xTIvBCWnMvB6yAZNWokUKyL+HVjRXny5CfBISUTU5DFSmfza
ZdkW8mWkuBNGNALAKlfytcdxSw34XT2AaVnUs+06igJxQ1yGmHDFqo0+cKuM6+bs
7mgJmOf+eDOnoWQHzDzuzA5/8dNzyNx7XoYDYHYdNNrn1bmIPojVIUyiz00OseX7
VJGpH1VhNvB8arkJMxPQeAwqNzmp+S6NW6EAkXGa79YvuuGU80Rk7KlWLqbC1ZH1
bPG1x4H8UH4768yyFdklZxKJob1AM326hz49xGrM3nw61aDK3rEdmiBI41GukWsv
VDJPO9VcsWwsB4rWEWCDAkI4cPpgFg6kOpVDV2te0SiscOJOt6VeTPFbEhNhrBA7
sBPP+FIkvh3VG5TP962ifrQEOpWZMKOesEDZNmE8UulItVwXGVuehG7fvvUR9Rf2
FGluFjKOh9IO7HOGQU3NviYuNXN+yeAEtOFr9Etp6REfomKTpe6VjGgG//W9wwnn
iDLGKRvamj3PgZkRjdXY14xwHp4uw3moUkdpfHQWu1FcpIfjEovZb2RqzDkj1Cbv
lOdyONe+W7NAKcXBhvsAkyg7n5X2Ja3a6NS9LCOXSiw0Pb9qPb2sQxVZDIo5mBQR
v8aZ3RuMnKei1i9fKr95FPX2gUIXMudJg+bI4n0TgqrP/0evJC8IkGgHAxCbxEkU
vE94A0wZTWlrrz0d+wENVHTVlmPJS3aQT05DcNAp5q6Rylh5I6h1DZwcMqQVvvdv
frEFyogNEKQ5CV/RjV0XSMupO7e57giCQ++wqPzrnHMuyVbL3E0drD+WvLBOW4+U
teaxzh8y10wOzH+uJMwF6scaYMM69BedvOGOD2KD1L7Z6RcI+BRxuEYaOaXZd65m
gMSlWZZ+gKHMrR0oTCRWfnGLKBx/UEsBcVn4+BaxtgS3dWrtFQSWM9Rbg/4QlWiC
aML6uLUh7f8gs1+Y17CHpxQM14DD/SLws09lss8rF9IXHexh2NaI4E3TEV2L0s9C
osOVsRKbKczo59546zE3yQUJ2Lhke2biwHerDfRlp8rmLGLybmftoBR8/X5AMmZn
qZcDCpMD34mNpiW2cn6qtav7kB8vnMEZ5jA+CiUE757duZy4DF97o8h3YgnJZzk/
/2eaERgh9qKvXeYhzRqoclNA04mxU0Way5xmyauME+yd+JAkwGz+Qxrw2Ll4HG1D
1T6AEUTULvrJRJoQ7v+yjuZIoLReela5LAPyurn5SWfNLIc+/nR6l5Jvl1XS4MuE
yQ9SJ9IH6yj99sE6LSL1lFdKAVxg0xPKFlBAEcafznY9cQwR17VXxpNFrMzxAhAT
9jXVtGnAWwtSvtPx4knT700It88sIdFJJcYUaR3jAWH7/53Lvk6gfc2TDboAJQYY
ygiu0gziLGONl70qUA+ToLA0XKtclsB39Eq8qdGmUm+HwmMdpA2joHlpGpUEeojZ
ej/vOGy6UrhphlKPFVK9lgrS/To8HU9jeX5yaK6+SnOMCxV99RLfVROELYr4tQAP
7OVkZvqibpDniyP1HnGnBYeV8ak8SDgyV2fbB1MROjnYAci47S6eNRNf7F+0f9r8
oZabpMSiqeuJsY9+kmdxDB2NWedhalLkcw6NpR6OtMb61j+InfINlMPNf2sd+66Y
+g2+sjNDQ44ce/fd8phPieKOVhm2pCGJSnZJmlKvFoHsc+/TguLrgUIYl3orbtWc
ECTgLOhZ6/ZUYwAmELZ0nGOS8CIIqugBQ0OuQ4juG8zQVytpWjOm6XDY0bOL06XE
jSoCfqrzvs5KlzrAbtV4HoP0QAJTC53i6PT+lZIX0jeTRoISGMn2XEKMcDhHeL+C
Fvi30odAtsdSf6HnSOd4bvbNN92mZSaN+mZvMV6mfTrG//tV6XLDRfrnOeHGcBUm
2KELSkSy4zvCMMIlQwdfjvmMnLjOwdjqaS/JEGSZllHVS1AAFf8GNvBEyob9p36w
DAuHAeoeel3Yj/nsCkrhJOBkV6etXiqk6cyJkk5zcD47W8/BJJuixBJnaov/iCbN
7iGGekYua7y0YUzryZs8p9yUqSFn1+EJ9qWUsZ5pTy+qidFhPPrFfhTJHrfPVuAL
FkpgJG5z9g0oGixvpML0qHgjU2rhCUH+e3Ko8mbq2NoSVuWZw5rF8D2oMrCgR1WO
smjL6BUYVJgk5GIQP+aA7BOb8cxCLYqZDsVSKy148ZHTAq+Lj4jQIuX0yzFfbmjS
9ErsmNPEQrEt0vLQwVpGubZGl/GXvAZ3xecOXiDsaphEnT3vkNxnDuFIMKg7jA7i
A0dtqgRlvjJ+gpKkhADJZ1AP98AgB15DYSK/rJDBl/3isWvlX6XYHxdRVX/b3ORz
NPqATcskz6R24X7AZeT6rep9gaH1v4rRRmsFBmfxKcISh9BsHjfK6JCYc/LovVgi
6XbgSFkTwnF+ZaiE8dHuhe4bJ67R/d15ZPZ7RkJ5LyMotwzUgx8H9az9SNyigh9X
DGBVgyyyJ2zgy9MHRel9x5Ll+CxxrWI75ldThqjxA+EvUmvGdCBw/Ghg0AQGfoNc
NtUlznfplD0WyIiU/Usgl0KZK6Fu458n1jA8W2fO6jtYa5vPW8pi7W8FpFKvo2Nm
2gsYX1WpdAV/sOYl15RUhwGeaUnM46Rpm6mHzrPpmtGmy5cjcWfPuSpE2j7Nuk4x
dTDKEXMC8/wDb7ozjhHlLqU1G8NsqLBFKTWREAket17LXo/AouiO3eD/Gvxc94oP
TfJD+WdWoZqeB8MtO7qgyT2yXk1nWTJeLGEjHTkePl19PCenW9VSHjqz9rOxaqb9
vv6ztgmw0KWIWWnjArNC1BbCnH3zT8KTWNcihr8fEwXyGYhKegfCSFUjwBAi4Mnb
vz5UtZPjvFN8CV2NTr3ay8hoscShRXtEbVnOe0jbxCrafWY+4K3o5mZ3bJCMTAjn
m+TmEJmt5QshCtLioxIxQQ3vTfOEnihxB6QpGhTRHS8QUOLJXnN0z8g+d3yHo3jI
yDgt0JdfL9ZjFiFXF9CPZHp82xKIB/dcRSdqvMcbAZcg9W9VQvVakRGX7FSoTUPs
zJ7YqRTPbMkvSMdLVM4z8SUJx725ONcLU/ipRuPd2+ERPozFvCWqs4T7YcDRBPqC
lMgE+1uQZqE2MfooDRCvaxuWgvh2y+ADlqn8ShtQ9Z5JK98ozltG2qTDtjjYfFRD
SiAU+Fipr6fMrLwiR5XoVQzs86AhwCFFw0s60KdMBhtl2pmjEa/N+Cjxu8GF3DmT
nc8FaLtVmXZ9m+f4HKK+BmaLBQjsMc1E/iQegSRo/TKIC3OYJzQaAMZ6v+Bulnlq
p9xMD0q2vWgZojh/uf4X0GxM04HnKj2PzW7c52nPGGIB0d3bcQB1J+yIfQfNJ/ec
f1bCsuHIuhALii3rDCpaQlKFve9LHh9L31rCdD1chvrgRXK1w9JA02719vq/LQ+j
e2fqirAld6aLZ8cNZhfSetuolhcZziLyz4ECgnUCeZR2tFQqoh0wlxXPViLETkT+
lTG/O2V5wwXdTbxZfLIOphEANXCUy+sokctPIq2yRX/lcA6D7n750GuCRbnyC7oF
VDvI6B98hcE6LgCG4oNbp5XkMG+a4hIt8Q8ftJhCQTQM1SoxxuUhojC6tkTiq6e6
UmSnU7NZdbH5NhrxH32i7uEbC7EaaBxRcEA/q3h8EZC+J1WMff3a+XBdaa5WMqvM
lPoKn4LTNTYQLVkx1U4KCIjZrSMMds7WbYFW/xFbTWOaFv6YoSkbWt92j9Ai/Koe
8c5kuRiG+Gfl7O/yourpK73n8dpZ7JwTICzjjOqiS+53bxT5J/rGm8yWSC62JBKG
FP0DY9r7lE3j9YIDQUeL6PPeOcB7urFjellcH1/CgEeGejqGI9hSob4qs9TOHni0
Hkh9mPCbgzxm9eiAdnuZCe6hoSLU+hYwv8PzoynZeFQp6dPMfAPkFLL//ZRR5Sg0
APjx2S8qjG11bODgDHoDSSrW6t5qN+glPafnNf7wQebEeuWCCxS4EN7iOJaNS3P5
ElMmEsRbhIOUSPgFGRSlk+TsURjwVHzvDdf8oKH9aFEH+0GTlS12G9I8LQbEfRtg
t8ofpklpLGblWfQUPe/EsqxT6KtaZXg1iakV77YSfb4FkqGvHUHRHf8vuN0z1Ej9
SWWj1n7oIKKV0KwthVG/w7P899qeOdNmtzOYtawUKbLhlD3jTJMwnfY1fOvEzkFO
iXLEME6jls95QEo9oDWedoHe5ZIYN74ZlLo9QVLWFdoxdbtY4V7ty2eqKygeIzFs
xKIiIsTttqrNsh+dhOU0jmldvn+ocZiGL+tuePCgfwZDXCyMncLHTDbfsRdHb9hB
Sgknn7Gc5CFWWazgG05ffzUZiQxwfGZJ63QMsoMwo1sWLRZsvz9MxZQbs3DIL8Rz
NrjFQ/5yHOEvIiGUh5YRyjARd1MHELba5+JbNjT+Y+YKJuX4V4GBBZmZ/zml7bbp
yZkoKT6PXTpfpbQ1Wa6w+Agfl2lkNL5fLJElvvQbPpTGv+ZiCND9NV0N5oJrJFsi
X+aMx1s73gAfA1EQJ20JKwP1FThELT+ihlOjIJ+u/W3ef1WjficsFJO6YeMc1lfd
G5rhIHRQnpAotpljTo4mPD1znx+KZtj5C8+vOj6k/WJy27hmp4FVoaFy6qLKWlzt
CxZkflQTvpPGM6OXm9+pQwafxsTf5vyF1su2EI21QH7ftPRSWD2Sy9sN5EFykZmm
bl09Yx6vohECTZ9ElfsZrJz3MWy0xw6t4tWDzAdRJ/imMwLrcjJxewE4zSRG35RJ
FqzPAbACcT2qO7YkFkm6zy8ReRjrBFmicMEjVBk1FTF1FOAOf5ZSXcZJOKDZvE53
AWHM74ujI+zJYan3YUowm9X2cukyItoyCpftaKrc1kE38LxhubEiE2ZdiB7wN3tr
crBCauUveKjg2ymxsxL1u2F/ndOL7WQI0xjTf2Ekjhc8s5M7h0kcDVz1+3EtYNLg
BGtVLPd5DlAOsriNZbQFN2sUw9Bc3C0Vrvua9YBom726/XoM80E3Sv0t6B069jxB
YanIesNzMsNZ3kLzCUbwemC22V27zrtmD+zdpChR0OL1FzgQ7xu7yATvuSOtZ8P+
sMrSjI8OlyCkgMQOjXQjlGI9Z0HynCVl4bcvLdSFAEakLk4MDJvQ3KTzXz2P493O
YPrMhEaTw9wg76VAYZEFLGlB5NSQhwJqmz+j6ae/OKb9VPr56oem9u4uv9g79iyv
EjQJN9pUb+uwVoTmVd3HBPTnHSd07M74bZrbpn1TUytBLUM5K1HdDdJ4Jy7ZIK/q
ckTM0sjIVBcLAkSIiu5rScuT7h/G04QQ08wc4+mlcJ/0RAFwbqfmGqqrrjxayWuE
aSlEip8evpa9ofpuKCJQT2n40gLUv47p/vl8cmFWJ0HyPYLthohQS6iswrSeBTyA
Dg4Z/kdAjmpAuPsepHltscqHxKTa8o06sJwqYYoVh/MCMQ5a99GnuuQktVCAs29k
y+gvQobjC2NBioW4J0W3V6q4zviA7boCJUcswKojH9olhGPXl/XuUBAJ7ZGF6Lxf
sgv9NxAEsKf1neKiUVQuDjvMg2JAllNiStRSZ7RcdBhQQXqexiWlePMHFvz1ZrWY
v3yyN23WxpbctQfwrsCMwSgRWONWsoJ7cOLPuDtQ2V3O8VTSthGgtOWpJZEUa1JZ
Qbpk76qqeLhfhnH69kh4u9pkjNtKf66OvuhXzgmOsF9ovVtl3Ua02GnGaOomeCKy
KoD62YS8xdKWo7uEoRofgS/7OSty6X3oomNd6VIaI2WMvtP94ZMMTN360NMsM49d
rWmhD3QSdeGSeF6V2CpmDCTevz+UWMEhKs9Q0qW8lP49mWGTUfGuEyMNzWLh4K5j
6Jta1/WZRZcDKgHfHiQztTL8949pmX13DKZn74JEARvTYKUIQVkDH1QbuQnnsusP
OP7e9oEVS0LNLJUHPhSF0DUyF8xB5dufQfNdT/GvKp8mABZZX8FdQBkXUy9jvrx3
eZF5K8RH6hcj6daH45N5YmloD5YpIzcd7y5J/EN2N9gKTE6dY5YLVio6g/qd7FyN
dNSr+spEKcqE8tg8g6g7OVIRm+oUCt0D7dWSl00AzyPoB/cGcQoGcQ0FTg2rdnlP
yHAiAOzzTrX9noXf0p4+TDNj9kqP09SPLPxDVxMezcodiiHYOaTwkbl/72Vm4h83
SZb+KYC0ICzMhkqFi14Qu4tta6dqwilWTUfTzLjDdcVYbkQCyqkprjReR6t7Z/mD
Ofa82aDmu0Eg6CIcbz3enR5MNdC+e4BFPBIV3ltmzzmYPa3CVnwnwqt6Kr2CUEeL
+dBokbZBPAHDCkYhayQBS5qNz/XR9F2Z1no5G+eZAJukHbzrQnCMcPBdhbyexbPr
0IwB0ry1W5FNzylqxw5bER4aBbtvskXbFpvYSgswao3bzn9Q6y1vxPyd3zPfhYGE
U7URC9VlFp+3zEp4kuzt0cbVWeUX+srPDP1Bwvyp262Ehbqg62uucRTB6TgH2W9o
f+5Lvjj1bjQSUYrXcOi/0CoqexxCbjPX3W9Ol04fDTyb6JS7EKBHsQuRMwKX0DlL
iEipJU10dDFwuY0WJ6Bb6YpCTV37RbG4vWgSsQotq5u0xpspz0Ej9aBEGNun9+BE
+24pLh6hHFy5HhkFcWVc62CFr/z5nsy4Rem684V2WluacSZ251Dxma3zJl7jNnAk
FMsmjWCG4cd1c3TJMFd83ohfXjuxH5IGCiIPIwQCIKUaq0hDBx2T0hsQAQCExvy8
WFY34wNhAlTpUiq/is/bpD/0l4n62H69TUQYcyseN6XK9kXiF8AKkCTuaVAFY1B6
IpicrL3oZeUgEtQQvBbLnRsx+eWafQnC2CLoJlIOGLHxnwPY7C/R1IJ14rcy9OvL
bXnQEs2tk3OWswGVcUbQohPCpXsuDAW9fxEn+9dZUsoKbITusd6MKijhO374vrPX
mAqusIYXI21JSBbDBn1hMJNDiYgYyW1xHPJa0Ydq4SDuvD0aN0pE96FzoOJsu2fH
uuBYhowpE5uNB0s5O0zRkboOhv5C3oemO9HzArgGKasQE7jvlp4m5aEaERklwcp7
EHkY6C3xsIRf1cLXlEDKy+a1EocceGs02JsG9f4sYWRNal9j6Z9aSrLf1aJF08ME
nCS1ALO3joYBcoYUs5D+tXfZkZkqOHzSZNP5CR8zQT6NHSk3AtZTtsc6OcLYNl0t
lYGshaE0xFPFAXKYLk2arVO+L+npZcbrOR8y3viwsYL3x7htfatAo+E2yxRvLA2S
+G1Grh2Y4bBcT2/6jVQi7ED7LBDawpR4kKLbpHYaZj/rG1bkdgDhL+OpATYYUctO
LlgoON6GmRnPURhp030nE9rztAfZ0vZxTs8BdaKpmi74qIi8rPSu6kbegqU89HS/
2QAzwpZTmW6Jd9pQEVae17EWniXvsVs7apa6TilhdVFqFDJR8TQ1E0+9FyfAFh7q
L4UxZzg+HVD6fEGxkxhUv9fBYHf4ZQ334aAwCM0UlqpByfqXzKztNYP5t6UPjP+N
tzhrXI29WheaQHbBCqMmkZ9oerGPC7jCgFso+/PHIoyLmpZyk3vAwxYaQ6lHJqPt
hTpQRT9frIgN3XpPWFtBsFe/x5y430M9LRHmulymUzxBsKfyYVd1Q+OEWDGyGkh+
buRl6qv1mb+nLc5V6cYbzY8vx5CRtiIjcYcUvDvF7DaG5/WSP9TfZS+YYGi4TtzG
vf5B9mGATtwXenvtvV/8DTa95+D+MM5x9/aUXWm+sqtKVzust7MTwSp/K5GpL1du
NJ8tnlskdeRATw5ptgWHTuVV8iFFI3lt8cwqWylNey84kOG4U6TJ1FCHUBQqCj8i
3XJi+mEVxbcXtVJ3K58PfAKUmXE1aJI/ZJI880WYgaCmN4adn1roR/bdb7YospI+
Y3TZedPP4BnNTVqLO8TX/5ybg07wBM6vaixmVYAJV+z0W2VADVvUa8xXCTNWNNAS
aqe1QqSg5D5ku8PC86e2JqMeq72zBpwjI/1aVlqZcr24AeAw1MswlYkpS16jEJus
mn1dWyDqLuccW4tQqM2QrrUp9EzHCZlnO4UgylkJSBx1nc3WByLsbfirynGHTYQP
6fOfpz6eliORRQm1zs03JR97jFMlGnUw/iQDE+74XGc9uSE3o6bUuq1bL/+JAPjf
QANcFAJChB57dTU30mLloE7cUBgk5FlBv5ih4MjGIDfX1atsYoeRhZWbFBeBuNVX
fJlHTmRHFuijrl19OQdUAGBeajX1JzlrRaGj7x9weqLJ5ozEAPMFkv9+hC1vsoTM
uj3APbHUVK3Mby8KrtrKad1as385caokmNlVo5DemYu/hFJF6CzCUuBTBdlhdsAh
amjVtRIqV/3Q2S/WT3MLGPr/veoVGjvXuU1EnT15kf8+LdosfBP/7fADSmvBISQh
YbDTFUbZuCpsIbCaMf0kqVW8Xgf+p4quh7uYq9yUvCcKnJALtN4T6wU04bJsHs/T
LqLdaBFLoJ9+5CutSGruKhmdDS/MVutAQ1thb1MiMQ/sWFVcIJv8ap5huDbCB85X
iUCIKtyDX5Rfv3ZZYLFuogSWjpW0Bp3nJkPAh4aQtdtRMX2Ev43xnXlAfnDcUUHk
pqwmazxqknDSi98lWLeP30p8zt2gjZretWkq3Ek1ikR5d7WlfhEWgFODsNMLmGyM
QhAmq2E7WOyzFhj93Mwg1si3F3VoRoJWoZlv4Xvgb/vpBLrOLrgf8jchq7V6zEgF
4toEks/ZNIgJ8bircfT0MqpNfpQ1s4OQJE3f/ik4wGrilOHKl93XPCvsHdWSNmpP
WtTcDL14GG5kHAC1pNFkakmLec9srlLHciDEoCC7eD+rxq+rWidGY6Q5gW5o4/0C
aq8aq9mdR0jifjE5HyPEEZGM5k5k4v1KJY2+nVIAaLTVOXt5dF97fEyCMnPvOUMd
NzhqZlmRn1n7b5aRFaRbvASxO6G/+snPUanC71WGMyRfVxMKk44xpVlKnZ0YP1WG
jdFCfPcz+UBpBwT2ZDndVXdF03uYTNV2qiHnpUhfrZx5gu37KbZcI9dW5wjiFUu+
RkUAsIEnSwTj1pTbFpglZBFKC8aCKFjYoJqjbokIGCSZuVq5n2a4bhdWnZ+KbvtA
d2czlIXmWvkOyrpLuwLSD0J71PCHhx4njF174S5mVm39DN0tB5j2lSZFBvZhNEi7
fb/Iy2z1Ne9Fxgu798Mc1EUkVvuUuhQOmKDt8B03OReCW/e1CDRHnkx2aknfwFq2
xS6I8TnhIl5Ps40OZcMb0HXhYbwvWH9RPu9MXXtG2r5UxMV6kARbvinekEqT3QfF
LQ8/1GfE6b2KZMAW/A8eaUNG0EyXX9NETVgO9a56kCJnosxfg4gCLURycB4XKPlL
ytKUls+DheO6wr56/PcZsFERxv9RfEDWh7JhqeUJDvCoVNndzDLAmjG6cOOKZrT9
gLHe74J5gU2T5aL1RfGAO5PsXk281B35BIQteKvXlMiPq8VwU1wrEL2PCA7l/sJP
AT1EYRpQyn1IoLf3ypPLDKWRZTwB1NSMuxcMOUBY1fK55Swu4qNDIAKu+XLgRT41
uauomXz23/L+xVaDMhCrGdYpyqaWcbjOyxKCweQ1gqYldC4ueXIJ7qaHHuo9t3Ps
89+QWDLZsmkpLAl7nyiC2DatWpzmHpqOwzL/VBJENKf/6rUDgjL6tC5H5SwEg381
H5gQFBL9gzeL+u7dp52GR7csbXNbkt3/2Ja9EItXEG/8HHDLHpJVOJPKRZ+5/zG/
DBV81ilHQwYp+hWyU1P5WZaoL+rSc/eJadqCvPwml3HXmL+Klgy8D0mLK+Hl9b0b
G+pcEyhJy4qhPbWZbZtLUMRfJEvJV2qAdwErFjmd4uoJnseqFwsnMxCyF+qJ5Lqz
ZxqYz9cz8Sic+YMCakoWvi6NcuYGWD7ITEEkP6WcjxcuTL8HVXdpno46JEGmTiSL
J2E2AOanWVBw4ijY98/NLMgBXhVpAu6qkDBV0v1lrgSE+JdeO1DkzrCpQpTFDfIx
gIrpGMfwZav2yc2SikycwyzMgygTW+WLflt3qi2ZOInS2IiZj+5PH01ZuMrFVmxP
DWZL3upyduFMCnG9/fmqZM7J0c3oYy2hXfjyRaXFv9FEbmn1t+3VoTIaUxHqM3UE
O2xN3JaT5U1ogXpr7TSE4L8XY7G2SZMAGuyra6UMecUZ8FqJ6yXpOIy9CQXHfysE
UhTKw5f2LyWEXVXYV49TxcoR+j8LGxiaf27jUG7UcaJnBpA6GuX3zQyvcNlkewC8
S+G4QAx1AcdTkMECY8RGLD+pe+AufYHzHn8ZdogAojbHlAs8gWbPfnyJWX7l5bSt
/crb/+BlCyZDl2sNNpFxlE7coG00M6GbAcgWuqZmLHrOrFIPx2ubBxAyYyXP4mAt
5NtqLW2tqwUVt0r7FeEFh4B6WkxdashRdB1RnGlUQ3TUV7mMV/+pYH2Fn0JkAenl
EVIzM/r1pJ+3e9vtFRW2ism8IaaJOC9LJBpvC3ruk3Zt7SP/gZjVaWsCeixYI+Y9
xPKGTQNly5f6kM+UoY96ioo1ghtgH8bSzrc2pyhRXlTQgtgOMbADF2ZGhTJDlKaG
CvsG2Jwc5+zixLb/XyiRptfLCrko+SagMnMb0yWkgkOrXPCNikDea3CiLgA1eX+S
MUM+UHcEfp5Uy5kcobXAeHLvDSQ7gLFK+5pLR/n4JeYyyKWSVqMUUjUckCYVldxQ
4lWqBm0QjyFLM7oAu0m+vVRxW4TqUataUgpCLkPl0z9QdCZ+u/hNjyMhzWX9/jYu
bSv6/0zDForuFH/MJbiEqFJsSB4tqx3wdW6/eIi8keHx+YwkpWDRBCHxD158H1dq
xvMTnlc4mREVqw7GvkbszA9OPsqGS1KIWuTOiCBDJQFuIY+Q/jcpgB7crvxU4UkN
TKNFe80/0S0tPqKTl2QNi9Ji38kClN0usa6JiSqk6sKIHOb1U0oB44RjKVnXHO3a
gGLRr2dUlwuea/7PvdK4lvXA6iQDVT5qsd7wc9rxjPC16eiELKzDxit6gwvza9eG
fI1byuZ65C45vYgaav+aub2WRH/fnRGRoVyHHw2TDBpjhOuLmKqkNHOe5oWc9ftH
fRijmC+zdnsxIGEuNtW/gbn0yockcDdizAWMNIN4DU5JVwbhECY7MHvGyTCOnoUz
bnyVyWw2btUAckM2ap2eeKflXek4ySYFAk0bIVgFbiIgjO/h9bBXtWHopwjAx64e
Ok7SXlSYUte3P0aXaQKZQYVweCzbPQGoC9AYXObSABIW0amRZUl7Y/OMc/Ij+Wxo
ANJUSGCKZUEwTUC98Z+1C1ZD4IF7PEwmngYMoG95/zEyIywNgTAyp91Ov4Qf3E+u
WzQNbdzw03nbSveyO8TiP4BPY0oc0cm/EmULXdEaGuTVUgdArcqrP+ujsadGC6F1
0T/dTScXvQgd82QX25M/upKoVbGMC8KgG0h7ayapIBl2Fepo1S8DXKo3sDM6D4X6
WBbWTs1EeA6LbJtD2HfWgHh+ljTZcwhsvZxvmo1K2wDkXAI62g0JIHwksi4kLHbj
/VTHM2aLS0NdTbhLKaFc0DyrfwVymeKQJrY0HU0vTLPwz/oUXYBQgyTF7e2BqY9S
TBu5HexW9xpP1GUap5tycGv7+vA2Pqtms6fAlwLEm06rx58utCdr9oIrwVn6m0WJ
rcoHH86aCKJVEAzIyA5Dq/EKZSt8V9icsCWehfAo+YLzWlfj9eJ+25KrTSIdjbBq
7KwJIWn7k5JgdG9lUEsGmTL89LJa99bBvIaCV5vuoBopJDHTXmOJlaT9U9/N+raN
WUjve/kEsrX1lcMMdPdcZueqXYgs3wNLDDDPcFtVoE3iJ2NDZ+pDkTsBdZuan1CQ
nttGb8BsprzCpXJ6T6Y7lroAb5u4loyS9k0VdSjuU3XE6cTbJw2MkG9DJdyblvem
vXHJuYUSbgxXd47r4OGZeFjv4arnllFW0dHBt3A4+9JeCkx4Lda16j7+Utk7uJfD
YQGZB3lWjJN+w7LnrIGB7PupGTDBxyXT3kkVWxo9+zzZ1qNziSxa94WDD+EMPd3f
oRH3W6Bo9en88SVzcZLzErVCxbGxhopGYsFVjIVtg59c2hVPm7Ebj33czVgMnhtH
zTW+aRW+1gJm7KHqRNfOrvZGkHoZpuRtOcSDnDSkfT7Gotj9a9bWZNk2pV8iAzW4
PyhA8ZtaYOFao9tBe5tR86I+kIhDm5wEmHiq+1vLUmFIhuPez/GInOMeIQ2gufqW
TnTkdpw+6Z9lTK5CtIxNCY/H1eIoCjVyG4/B9lUtJnLRnsriHBaQpd7ay8PaAXIe
CUaEPi2oQEmmli1n/B6aCq0Nwx1N1doGLTJnH1XpzRUPfxNd6tC+QN7/TUJ+TEAS
PJ0HkONeDM9P1jTfkwEgS5Heqs1x7dz2UxR88KJB/bS+RnDT4yplXRG7mM0qmnXz
0sFLZQXgP2MyBvfoU5VeKfaaZLjlk5F1Bah1Mj8fxrNKwHAvQkMUbyFZAw6dpGXI
xaId2eQR7x+PN+/UPsHe1j/9IypvfnBq31slbFRV0z08aHDwNQD9dyr9wWfp+Sbv
mGcUx1tQrEtnHNj+QHHN/NkfoX1FyxjjzIy1oJtcthnqQDB1o4rh7k6tnUlDfjlM
z6zk+7nGGA/AYlmDYvMHdS/yNq8yOmiI1rEzXEXD4WE8JA9zaPQEk/g9NlPveVcK
njiMp1hcxQQPw+iygYrzUtxoVHqRMJxKrR+aaOKG/dTWZi6+9DXU5hBhjkqZE0Ca
G3i9fF7ecuPQzeyeXucZnnSayF1OdW9SmCfUQuPjrUavhwj9FNyBpswlNycDgg+y
GPwvo25tAi01qdiZo5CXuwmGJsRD7touhe4oKXCw6hxb+oj4liCraJN0QFtD/ooH
afUPKHmpBVxN4CzhkO/TcQ++pjr35R+zf8XjMbKGrj3gYK42cURlGd+03HpjXkNz
jhWnsMEd/MSUs1fnwKTZ2NarZWrbb9sjX0fDRQFJHB8mJ/ns7Hj0li6vL/xSOjEX
+6bbxGAprnyF1LL3E6ww9a067Ulht+FZk0MUXl+tHJNDKArDtKf4VYcfNEcwHYx1
c1MRzPE0JQAyJsIh/gxe3hwng48MV9nHHRDMCOQCkh1gn4cyBYM1tqSscFtGojoR
chde/LB/VgGYDxy6D1DxiZEOirOSsyInQuqXiw+8Dz+acjlXsHLCSVoqCZw9G3T8
ZcIUPL4Agf1Z66pExSs0uj6bMRoFj0fR9oMTvjkgXMteCDQyKnDp0xEH9pLyUJCg
kJaCQlt+rjFivEHwAWpNgPlybNI6637c6j3S8xAglO4Sm3pUGoa5Ybx+wxRAE+hk
8ERHPo6YE/daaqzo86mSUHizVmlHGhM+hNLP/TlRzhi6YUMGnhfrOcxgFdx0VA3C
Y/JZN9bodiVuwDuKQN9A/syQEMN4z4sEaAzV66QvyvmEtTxzv8WMnv3pYO2hY+AA
orU97up9oh4ZLP8ftAC9n2otHSR9X0k9O/V3JL7N7IsXTlDv72xk/BDuodlkQXsO
r+buctDQ782IjCfxzDt6ipsooHaUtNrpM568VfjkZifPhVz7m4xJl9rXPnQrtCY2
9p7ITC5AwF4ne8wN37RXQJxduvhuARk9Kxf5EBy7Dv2WeEb6RTzTZeexe5Taasbj
fb0HjVUikBc46w6I4Zw62Wyn/CQXhBptuXNMMJ6Mo7Te2wIqRrBW+lMsf/5c2sN9
yXTUeDDReHC9dmVGa4FU7DWR3IBYj9ukrW1aKH1K1AbrrUdmoixQ0FHYzysW1q+8
Ua3sioukZQNbG+rVVEV0D6ppyuhzaEUEqMHS3irtXPBqGRuv0hLmipZdVOZqFfw6
x+jS+uNUFGzrm/BfjJbQAJpi17+VtHoneEVAAJU50JN868DIpCILqZ9nDU0ECXnA
U1Q8ARaylV7UKBxrBDTbBpfk4K0G57nSHQVXhQJaAa3gK+ey+cCJ+HX/fMP8ZlTN
o2RLd/xHEODReKQ4qhDw6yjtSfx+dyCOvpIem2uq1DNgkQHlI5XXdjxlBY7RAk4M
xlBX7E0d1Hi+gbVu7rZ/ETK/Onmo6SfiDsKozB11ZbC+xo1ZU+cFX/UHqQLNkSYD
dn2tWfMSYtqFZK6Ap3zbu6JXtFIS2qUI3lQYZdyTuA8v604/4vOH5z58wNRK/8k/
6jFm4a2li2TkCq6+sgoifAGGE9Um/tztaDLGLRfv8c0sDC61brYtW8iXtJHRIdja
2CDRGM7uNuKENiAjy96S72ZdZtQ6XlXHR1E1Jfasx/6OX24/pbvyva55A+AnMBDn
XTNmhRjojpcNhaDuRiwuTG81vDHyMnuhIJRSf0xJ1JI58gd67MxHFZllVsBD5ab3
qFp7Og/qGxxCaSTmyLcMxob7IPwLz4fvUu8sznfjRCAADtWqL0EEDwQ0HFgNp9R+
LGXvSJNUiwmekQqeM8z9zjAZQaBA2JzJ6K3u2dsDGllis0Hzj16QnaRbT4qvBnG+
JHMY4xxuMY/bBg0GXyCXJ2KIOkIdlpKGLtb2UmC8ILdojpAwrdEBq9daCN8TdCgu
GWAas8lc09588YZjOO/ICQ1e3IG1dTJHS8JO5Ja5+2sbE1DwV6c53WD0bX4QPitU
1VuD+SwV7uSPyIjPCiNsz81C4dL3o7L6f/KVmUuIHfoB8pn46+2p9uCiyQzy0rfS
KNDmUfK3nl/hqb+aOi7LGcCHCXEIOnmBdHdWghI7rliYVRGFDrH0pLFOSa8udjPU
Ppxnq/UjIg0pSyv2+/vO64DBu1zYpBoRpgH0hgnEkDBdgcrazn+WGGV1uHkdXwPd
WCehDNEfxY2+8+oeh05cKo9i4mYsZ7t+UqAmFhoREX35Xpshw0bO+/FE/l2PyIJQ
2rWxUD91BqUAJW5Bo39lvQVDiT2XPPKj2jiaVLG+R22wBhoPrjGJSbDLJjuixUZU
/y60VdEykPLF42+VMP2BPiO4UnF6MF9ppME4r3S/psuBEsYGE2LmVgPGeQ9tfCej
Gx+BSMZ9wCQztKIi9Vsw513CL+ho9Fi6Yw4mELMIQnkWC/ic/atssrfasbuLZ1oe
pvBZI9RN2o0jNDPlwD3xpY2yQ7PTTSMzd6Oihld1h+Yfge+2ysVJZNf8Y83SLOiO
8fuqiNkYiezRTsxBULLiuWZ1QIQ9S0wiVwog3kQAlxLvcU139N5SvJ9Blj5jg068
p+C4l2wFk9zT9t49ZNv6elr4RctpZGvV+1eO0iXXXqdPZJPb5066alP3IZHMyum9
plQimuhYGkuwLkrMeb4v2H+WCMcErfJ9DBmaUUwb1RTHgNHaHewjlqLSHMJd086P
Q0u/U6hpbXNJUahTQlC0bb4EyCik3mAsa2dHgvVQoKz/CWzWYltjrPdUO+DUJ6mv
FLnKpcyZAiYgGz888p4wqmr00ezJVEAv6CR3w6nxy8wwzU3USvKlVWQQ6KFOIakM
GGz5NYfS8IMzElQ0DSQCXMeY+SsJ+WWdJgfRDfO5e6qF3Yp0gT7P3F7HLOYX1Zdi
CmY8SC9HZ1YwjVAONS019DUy7o0Bkth6Qmty7rMUgMMLiKAbbppuj51mJl8Jjszc
CNq0aDrtNzyKiuFzK688Y1BzRWUTXgVTnBl7OanjaKFSKGHNWVlX08TaURCalt/f
A/t7xIIZOvUiSMWuQ47RZeAQEf45lmVBVeQSoObaAzH6+Kdix3r345CcBVm1C7zt
RiS0SvVC6/wk63kw1UBKvc6pH8KlnZhad0ma8nnFkke1VBPM0kkrHBEjglv63Yjg
Te7bW2zXzfEyPCmWTwoS3m1D/fGsDnPvfp/ymeV1juER7CkasKQgo/+Pqm0gGOgj
cTHeEGjAhbpIF5PtehcOJSnTk9isgzGFydpfiAt3MCNzh1CfKWCYG26H9jAfx9ic
V5UoqQBdDz/N1JnN8Qz5VpmdEZtwIjWbYtePy9FEXPoABkef4PqjIn/29wplXKp4
PE33aSKE5PcLGt7qwi3Yed5I0tasVS+GHXVQRsjD7L3lfLzlOPmQWifKzlIbjpZW
hSakz2tB+OtHimNI5y3mkLwFtcucLtOcSC9QeepBWN+urhIXnsw29OR+JqsKTzJz
pYShUBBIDXPonzOWXvuLNnaMYCtp4ssvMpe6pX0Nu3BzmivZKN5RVieF7UiGE+wy
HCprHW5cubELQTLChGnM9OVo2lwHU0yUyAQJgUpC+Qx+KpeCy5KCREsNQgvsTUyE
SfXpcadqhcC+RGQB2VkUtsD4wt9JEE41wvfAzBpco7Ah6MwobkVL995OZUlicJzR
OGsxrwKmpDnF1scqIA3W+0ykgQFI9pzUyfL6a1EjGc9jDAttxezcKM5y/XM1iK8F
jCvy+g0zgWtXZPZ/XnB1cch0G+W/tTDpWaF7QpMor/KiiDsEVlFfSUhnhWNMB9W3
Y0l/ByeH03AjdtSZOnL/+mW80PjVs0lWGaDUFgqnZwtvBxP7G5ZkCx73gCIuHRgL
cU6vdnrUuxmpAa0V1TAITGYNUgjQKr1gnBgzCDPKmrrOxN+8HnN8FEELpwcf8q+P
Ft1YE2aW2+vGF3S8wKk3LtQy2xCSy7p9gT1H+l94YCBjrfnYPbGcqvX5cIdDfvAr
UdZVyptWh/oJEXjuV58nphj70eZTrTzR2SfQIfEQNMzPXPe2Le1jNeifyYaA0dO7
WQzJM/Jp44VFIYsV+GV7CDlPWEo/p7+gM4hxi0lxOPzv+2kY50P1H1gJlVyCITEO
TLt3u4o2lNqt8MZHcqHtEoeos1kJuGrkJwsbGVelr84CXHVRHcq4sDv9xBLNvFBi
hAWrIEtm/xmG0OTfa2RxmMEDlOzCdZAcLosmawNRQBL3GBIGny0rGOJCUihHQQf3
+fCSUGUmEmlomCfB0ob+Ta+534Vlr1pYjibgBqfey0Si9gvv/NPlfJG3V9t2+YIg
k90agabSgnjdBMH9AfOzmhMpLajbib5Ez+Souxuy5cPE/ggLvRShQUERh0TAVpjh
fIE7UDLDQy4+TcD25MLlwkdfp9ti5rVrq8Uoa5/AEPceIrUDSlKMbkWrXwjujH/D
A9TgWczAVaXDwgjwRZbMmeUIuDB5F4CmP6xpBHNvCUAU078t89wFHSHFTovYCW8B
fGk3Q1ugJCrADuHlwLUsr14RQX4mHWdEGvi+jKMuanBDEg5NM+sRCyuR8OFdE51T
xiRrMu7Qa8YRQeD45TObAfktHljQrXgXBS9Exh7lnDsTdBz+TSfPCdvG7eQVhqWm
Dkmq4LpGmTGclJgxrtt5ko49Rzv6Gj+dNj6W6Uyr5eK+LuCsAVvmWPdVMgrkKRF8
1juuCB3IqkX+iE58S6h9BmgPr/PnGE70zIq25V117t14jPqq++FU/g0btgAkNSgx
TS9MX6dO2KuoYsxcFkX8qxh7eJCbaC9YFobYA5l22hUW/jdUwpmlv+r+7eakrXoS
Q7Zp6mmwBET8SbowDalh1WYCf5r+8njjf7h/z3P7+bD9E88/OoQgIos30h/bK+Z/
21a1mdQ/muJvHGmjTZR9s7VsqjQtQjllanoj/OWkAWv+T5889QH2TWgsyXGSo+MV
rOqDZVH+CbHcGE98JlnPQTPDvE1j/knLWIKZth1gpyXNY7jhqZ0XoF2zTkZLRghi
SZgbebifWeHEq4cWRBATm9rj1IAwF/E9seA+kyyRFGZu2n5k3u+i9SPwAdwv5Idg
0crC4Tp6lfKnar76lnJZ6F7VmzklUFulYBfWZ44MDNzeteGECmPgBZqBF44CcXAN
xi3D/6N4pid5mDgOdtiO74KP4pYt7SCStgO1d2h+HHInFBME8uTtlLAAtGolz3Vq
p9rXdoQV5cPLOz6m4bcv/vWGVr9g3PFu+mlJ4mFriUkQoAOuc9lDuSdGAAqk5qks
BuMHi6vQAMSNDLSx5EJkh8DqvrAn8NSKEMOhWGCGjQUE3/Hx04+/XZWBjHLgvO7i
/u/KtKyPj8dEUEejRzWLJuHKagLmekEmftkw1KDmr1LVF3nT6AG2HGWdz1a6BQ6G
fLb5WOaOAYXZiaWgtjaoMNgi0XtRL28f6x8jRz7Ey56A7E+/asObZ79mmuMd9CD0
yFp5Du1qvO7If74r4pGTORpwItkMwBRXZbWFEhLywWVZTf2SPmOk9z29uLENWr9r
fYjkuxUso/LcTN/RwYii1wSdDVxoYrO8ZWGm+jdHw28nBtY+Zawr7KYfUAZgE2M6
161aCDT+VCVeaCBx00fQ3UbwJM+Jha7vtsZ4s6I3rWp9hGCcmhYl2moRxni3xvm3
TvIOe9XbmMLfUToQj1d+fhgh1T7RP0cWKeH0+LmG61R5woJJu7So1J14oVkx7DID
7JG4Y8UTThr3F4acpG9noc1wzaHpOn9Ru/oc0oYnSm7eiA36/K/6xP8ZjHrgyDt1
20XSFaF1N4e+N1CX1PDoAH0umwW119wcROTagzXpveLn8kgfGiJIOkS6BX8CT0NY
8/3aQX4KtU0d3bm8+Ku9Vk/++tGVx0yjpohK0jgGJGATBBDOk+QJSuBaL9NGfu/v
H5uDqIhQ4xHBD4GeCEDNJoW3XofKXxOFNyjP5cl6ad6mpZxuJe/rYDM61kW08PvT
2sYdG9mmT/3yd/e8UIdam8H1KaQvhETM7M3gzTGd7kZQ27jNJAyn27efB5XkWGMQ
UK68efYARAce2GF5SxNWqpYq27JzrIfpnd1qQSdKnrF0czmwE6+bh6Fwf4sDjtdR
aqqyHAJ1LZyekXE/SM/aIt7C/RI5iA/RKSWJAkYjEQf0rPaYY4/4n2BX/D+bjruz
nKzc89cuvXtVfucAiAqkd2dEfdyK4e5g1AiVGwVPUENi+wNHMiGQ4uJHgunqIOwe
PZYP5Lfy1yb87bvqaTiJATd2tDLZIednnPG0Pb5vlfJ+W0v7PMNX9snqsqR/exzV
O5vZ97KqnhwM6ILdzxkdYdJa+LVIWSA+sf4URD+q4xenfLDT1JjBmQP5t+ASaNd5
Ue79ME8O+c2ijwnvfEJmP2caxp521x1azvDZgofztCYCW+T2wpPFwKk8vvUsUCv7
+icZU92clPoLfvpnIC2mvSm9+CVnJPQg9sI53XihCki3/2xSGsNvLrrb235Bre+X
we0BGPf+La51/Gao5zZL1Ux7uQdsoorHWOqlVU3IaxkKuqrg7kpua+jpgUTnMRoO
zlNlXXDS/Ee8EDvVasdocNB5k4k7NIBzpS7Ij7Vdi4Tuy3D+DYTCU6er9kCdpccJ
kqQIaVf0KhLZBVwqPi969xYdQIaGJyJEHyV4tk9k95Y2Kn12X2qRXa0A8nCEJ/PK
kCehTA0qvMi4bDNCovd7MZckWRRudC66j8On3e7HoIym9Ks9vIKrpe/mblGcLdyj
tCapXREyKZn/qYJE822YGS+lndkGabofJ+DfB26CNcG4sLfWUnVptYalkmE6XPXj
Q2eU3ds0tYVBfZNeaky297RVk7tAQw1nTigknpQEBcTkbmy3POIgYdhQLH9cDAVL
RloVzL9xKCSXz0oIukC3nqA7hIrCq2WuAFVvrLzoc5ype/A+2gfbbSXmoKRdSefo
aNuCNBaDzDPnTstjbrHYvWQBRM4B4rOBSJXteOAKRAhYI+/NpXPM//BiCZ3mKRFV
oXA/iHNq9ApLVdr7WUSmWQgmw4INGCj0JNHsZluAkVGY4uzGCIVSWB70MzR9LKet
sArlevAihgz3B1ja+Joh2jo11PfVsbhl67sF/ow4BubkDbOXBRgGC2m5GrJ/lggM
Yvgn3Ykgm04eK1SIHwj5hrKccShR7GDWM4JHsqBDP4VQg05zq7yH10EtxDpbdPX1
n8cwEXJhq0cKRzlJElVSsw4H+PxMTzPqRBtjL6auatFLpNeLuD9u0yKzqVhWlcAK
0AqEC1eYpf7LhedaqxYwne5N3OrMAhbotIi66tQZLRiL45QDCS+FLT247jN5blS2
QdJOHV/XBi2/3JwtQzqVSuHqTiOuIdVo+0fZ9UvS6kz1u9KIj+BFK1uVae0RrzJt
Ubyiha3K7UxhHk2VbSvsIVzb8a2kLj2xBDbI5pgMnCE6uc4PTCSEaL1UE6lANWyl
xuUR5ybuy6UWWbEBgnCzG+aCJBrer/AHaYoTXTB7qJc40rygs7ZuC1HDctXMoX9u
N+prcig2bI5wG0NU5ykB1LF5Y4dZWpgGEQr33oeDsfFAgtXC0U81aauksEBcgOa3
O4eWeQqBW6Obl+UhJBzjckTkVy9U6k+HLkVKEJuW9cwhbC9FnznFqp1ncDN8Jg38
Whrj9wSdYrxjENfhzDJW5HSPWvxKE4DXReJGqPLqkZYdNrUogd6Sy5flKn2DPqi2
3qs1HtlSHOislzzbr7naALKbWkKiEwNm1sjGXwaMtTHycj/CEcUUP1PSv4BP223w
64cHKVY+Mqip6G+qkp1U3UD3MzwuXkQy8kQhcsHN2k4pwrVSNT1pjkMoyvsEGdEy
duWaqCGO7RyjCmYABCVtzmfFcqn67SKC9OyA7/S8aHSszMQmAaF97X57D4z9om9/
N/ISuuRpAYvKlJL0DV7SxBhefjZ7J8lJJemGRRr4JXa1WgpIu7m+YI8/FnYiWd11
OP52/LJAr685FNmjsopnnYY5UqRp1B5pIROsizsYjj4sEvbek28QCh/6kS81TDT3
X1biNrSIKZIFbKczpIdzHDu+NOen2EzsR54gRtgA1Lpm/gQ7ixMKktv3lBU3fNS7
fQR386A/UNDgzKIHhDtixCzY3Bs/zVMPTnDWGmA5rhcvobMUak/36G+QNl6zqoPS
pnjSy1rMYY4glplzXcmxUh4JClrIjq6tqQPkcSGkxHLrytJZ2QP+TQVEVlaKzWt2
NCwIDpCfN8gbMHDiyjv85sTu0LJsbNEi4qMVCTX+bF4znHR1byGHWuWHGqZoLp0R
OAjHFdfMjP0/+eZeUZgzs+LaTrPQM17FauHVccRk3TbTI7Ek80zrI8nbwNP9oJxo
bTqeYIsQGSULYB6EkoQqz1P5iBKgmWybsEjxbM6ykkmQIaq71GDqwnhpwLLT4rvS
LylSmnvUleQaT7FuvGtg9jYn11VUwMXIIb2JiRjly2GL1hRdVIkd7b3nbTP93HFg
+zTStHRl3isknIxh41HPoBwdUxpiW6rhMOKvEDft2gI1LBO8QBEgcXm00+GrM33B
FgdPIGYlbDAIXFZpTK1I5N20DvP6HWbImc6EGXe6ccPhu/djew7gwpvbA34XfS3C
2FMMVZ6rEA2TVSog56JT2rwHmeOYHvcfEFFp7jmCIaufRRl4Y9t7g8KN6Rge9DnK
TD3ga6RcsKqsaURaPapLY8S9pqm3Mq9DTjjwr9173TDpRhoY0y8AatAQ/MUCeWEV
D3fvRsrEi217OT+Bfywoq75dH+w0W+fHwwZpydVWQOUIAYmjMDNC35iXMRAEuX8P
odjDrDowEYQWNzVDYcwDaKHuwZDo/YFgHUXt4VCycmMmIyHCw64lMey2Yf8mG/a4
hNhZuHDRwhIAfuskK+kJZinYkJZCy4Op6II2xFciyz9mI8t5ZUCxpwJcOjRX/VzR
pg5Nz+En4bMN0CMI79el6w+Fed7ZM4RnLNEoLUJorX2/ENf2i+qgfet3AMX+0FTx
99jf1v/i0jP9AhTMaDLydNOn42tmrKdMNIIwZUK0P4B8Mcl2Pj3E1Mzqx4GdBQb0
ilw4jEXo46qT50v14j1JN3cQnyAPYP/EdtN+HKOWSQbT/T9ZQQSzl3nyXi/ZmEVp
n1Hu1sCYCYT4KH1sy4ucZjQkRLUq1emqz3tLuSGoMVEbSRWFYyHY0Sj64yw5Mc/c
PFSANOPtK6dPdbtYII4SOT6OTJARpvkff2jdNuPJ5MtHsKxYPXOyGIgG2Wyn0bF0
LRyca+lDvhopuTd+j8tRw6B5nPcw3L/zqYJ4/+fh5frZ65nIWarJdbJAE5GPF2rZ
8HJaY/e7J3pRw4BoBtma55Z97vV1Uuj8puEB3DSS7At1GMvm922rpcJ47qbG8U11
mb3ILZYbJgiHYBSm9uudFRSHb2bJ3iZbUw9zZA9WDS5+8gTRUExqv5f+pP/39fm0
OG7fVwxAt5NJx70cEvh+23ZFyToHHB2FRv/aA4AFoEVsTR6JOtbtE4EuLCWZp54L
QkQ8w2F71v9EST+ZlA41AarGlRrOAnzpgDXdF5dBeed49ub1Co5hSwcC6dyoXq7y
dsdRomjitho3lV/ER3PwWExxOQMISNV7fgKpooZ0IhefA2WCsfehfJfdRUdE13Xy
yG4Q5oB32dGaRyLrxB069AMwEqp84Mkj5AIb3miiyZTarPOFeOTuEPd/fKygSoE9
/QrSFzxEs4g5IxH4XPR6s4woNRe8UnJrn9/ny4oWUUKHXuGOJpKg7l7iPmrDOq4x
9aiKLXhDVDsI+DL76TWMbzYPx0LR3EbUvlGH8CIZwc4SPYIkgefytn1U+FK/B2qs
kKIf9QR5P/Ua5xbi+bJFx81d8UuNTNNzgHXBnMtsDDTc7SBTqwOo41ac/Ye++YyC
HkAo7bhL3SHWlhIwhQ7dWln0P2vSVOhgzoVJgel8F9wXyLKEdRHYtfNufNL73I1e
No7zUXomRn+JCQrvO2T2QNX5tjZWgPZQDSqiJkQhPOByk5FmYOaFVaCykgKEjPTK
HDvQPr+m6OJgjeE3+meBic05lbK2wRk24slZhJXV1sXUmsZWbbh12zm5SpSJfySp
Rk1AlO1XytSPsHz5oaYhUZh85TNeBFEd2EhuUuOgjhs41CV+RPrlLSR+is9KPDKh
Ht+BrZDoNq2Ck0NiTkpmy8DFpZ1jDypsCr4lNY0/TNShrwlRyXY9yvUoZiEvhsCD
DgXKXMowsqfK8gV7PdRV7kgxzyW9U7qoQtXGQi3zQAucvB3SMuZ7JvF70+emHQvM
Y0VZBaWVI3D7ERnzZEOdD4cbfvQvnm17O7GXUtj5O/aN6K4rFjWXlao1jgAwAN3L
UY3KDhXS7KQq8LF4u2tfbMNwk3MFfECxUugbN02idfvULpHE6x8qKSwbrqAcSnJG
Ekr7xKrcz0bwdFPhC5gdFjL5zrn0HimfkoOQZbWg+KZmJ0PecWyQUQBYb3vWV7km
1C3V1UeHCp7Gg5SdzAPqmkj7yPnFejj0EyDEbw1siZaTqcdK05WUBU64DbPUlIkz
jLojm1VX1wkqVnySIv8p+X4ZfJ0jrSYX+pYvwm9qGBy6HqrSTD/iBQqfwMDCs7Pn
Y/oqr7D13sGgxFTrRQuy9K0gNqnE53OJRiCs2agaUX5bfmDOllsR6NcntwbizIMq
y/aXLJBciyjQvjmY5YyJdia+9G6i7QdGYRY3wTqsn/6W2YDHIZVisxjQkr9mY0lY
KS/czBFjIxeIitURf5fuTDidzxN89VkmJH4FGctSQODGWpUSdgIq2fX+3RAex/Dd
UvD4CQoo6lM0j8kc71LdCikQEAuLsT6MeEBsrLYFkNmrdzsu8+I+ZbNehHs/ovuM
hrIupOaeduH1x2HwKK+AsEn0XsOEweyUqxnaf5dXy3O+EZm4RIBhILjpdSMNBZoJ
3XF5SD8oUNufJ3o3O6sPmntLvCunaEgzIorGMKELIuPpiZlm1gqP+4E7PJVfKi1e
XB++333305vd6O3sP/4Mi3CvI7tg/1KBBtppU6wWsqF5BPKGYyolSt/Bu7mlbBRl
uCgDR91iFNNhx5QDrhwEXTy7s/lBXEv+fILhqN57KpB81IDmEW7gacqddjbj17PU
B0pmHU4dai8hUEgm5OMy2vaR7TAMW5hXnqzeh/8BQE5XrQZAE9paWn1v7CEWqMfl
ngNfalhT6X2myfM4j4eMJB4+rE+IhwK8JBsisGlMI7wxvg9E+l5FX+5/ajy1DQjP
+6jaZhnjdSr7uPVmV0SuZrN2bL+N2XPP3XPKaRTNBeg/ly+kLrZsz8E5DaaXalqw
MbwmZRq/7jBU9VuCVJFrNJ6BeCg2d3X1s9dsxKA6+Pynn+9DQPlvfSAzBbLts7NM
e7cNYb4atnthvNOB1SdJXUHpdZMP6PxWYoMDFhFCaj/QcKKrUpsyqekyg1GA+O9L
gLihqMb7TfIdd3z7+pqgZBMXnQZDcnEBF1xCN7qEeQ+EGOO1xtTTjfp+iq8ddUvL
KWJAPR3aoql6bgiGo07jyCMWU3HGIXrl+v4ZwPWXzVUm6g4zM2eaP7aC5p2S4y2H
zowIA92uaCe8/hyAXnQ1e0+5IwjCWdK2FY8aplsZWhb+C6frwtpXdHwdoJWYpeOJ
1iNmdZdstbchuZyr6wgPUl2CzuTAT2yFZyBYGHdoM3cexkCZaecCo/lybFQsqXyW
lIHq26jc2LFK5NgB0K2v4J7iLMsKUIn32AwlPLVO5BpwxV90tEBGaodQdABd0LgD
oE5oyGc8bTihIGNDkPRs7jwJKqqR5pNOvfokx155VJHYcc+y/ARTs4Din+n0R4rK
W2ePNAeyB/Qc9ImxuW43ZLQrzSa88eZfo2XKWSwk/FeHiTXFHAYpTHg+ofeqsF4X
yyyWdIEYZ23wyw+ZxUWAk2YJsc1q9QEtGjEE28OGl+VdyHiRVgIXzZucJgDYb0qE
0rr27qGHXzofDhLd4zrfpByHl0sBKZP35ahKzDnMUrCrvPiC+TdISobTURLDhoKC
dVKgGqZxmIdzx3lFHDwE/3vPAvrLWXq9dOec7cDE204sqUuWHHhhV6RVtjX5yeZh
l3MFEGPXZJmn+3P46XMCuzYKxlONoe2nurfpCU4e5ddub9yg4XitPgH343z2GkTP
NM8mJVN2dU6T5EWEPvNenUk0dzw4JnjE7rwy94nlh6IgwunoG5J+MJy79b+bfVvp
IOeU9Qt/9ZZOhEq/tpcm+AncGMp7b+prVmvuuylL6wrXvy8PO8nChZSV/wHj1/xX
92/0kbjpkUys+uLQ0M/drw14LSCGTAsGhMBODYwFWSXOWxuWu0/IGPSeyAJFcGQP
G9Jv9qYDs4hh8BbcTZkdNEbE8ephRjWv8fUyYL1jkTtbtPkgZ7dAZWTcOYZOEZmn
VjwA65qq6LDf2UaQ7WdcA709y/xf5P80Z9H4LfAJ6/oP3teLr0kif58TpJ9E8Qdc
6nKRvnqIgGn924OrtvZBB7op0lcjiTVQmmg0HQZjN++vyvYEMoudRuEBTmiF4oj+
JOWMUEeZ0/86Eq1MxA0Y8czeKcat3fHK2D68yTLGf33Vu+prx8+SUF9DgUo+GPex
9BLh7tiuO+FliXR1Nwi9lkrGyg4yyKK/ugBmdgLp9p8hjmcaA+WevZkFHbhQrgal
ljgh8jkvmZ4gLxZX118fnbTfZBRQ12G3OnZnV6EK/Zqsc0J19HTW1JyoPQSdkvUQ
qYosOg4UxigPLCNZKUc+8nHK+gg2dIivzbLFRfnJ0zUQFqRBP4x0SBhtcGD7z5qD
SeAtbV1Wxw+l91BBSqPjfZDD50w2uombQ2rzYyZOF3abDnn9yHidTsxbSHK6DuCU
VEdK9Hkl9NkWB2dlquCY3UBJ32MmI1eJtN6qLLKsx6sbt6ro0YzeLjZa9kBIx6dO
IserP8+GoyQLSQzXndsWaF7tglLcsDW7OZ9+zj7wEywHaaBpBNhu74wVregE3y6p
ucXFXeX/8CKHSp4D8scPr+Y1F97RbCEVOUhDTYHBS/J8+Y8eEl0kUsc4zvXq+8iq
s/m04BF3vN4HGQxMYfJmjPm59HdUSg1AldNYOr93gMH1GondMgwdcPjVa5Are6Ng
jrjc1xOSivPHeN5GID3pKftpvKwUS1HV+tDoMlr9/ow6HkBARnyyOvfFhtEweM1Y
JjPxHzikWdDsMFDludDsNPINYRknYEnJYTq0gjnrRkORmZ3dc81/Iygy3piJkvfI
L13zAn5v2FdZPIe+21wrOQJoPjibw/43J9NfdbsgbLYZJdCkU1Z9KVVHNGGWdbLt
4q2Uayw++A7bglJPTZBCGYAyIh7oZGRlZ14C15RNdtvwDyNr9Byj5KR26WHbFiVb
1jSqYZQ6l1ebG7yGzJc8l+mIozPRse0HFlPASLJXbribZrofjTJ/4vX9lanR4BWb
jSLFII7B0MTi0/IwUXYg8iwKyFBci1tpo+7mCH2+fMK+sRtvaXdkcgf7i8sMZo3J
7mXH1WeYhg2kYB/Ztv6Z89+NGslncieUznNcvfnyE3UOU0HnWWC/K3yiX8LTSq/+
6uyIigCR/+SNXBgJ/w3KJEL1BgCK0QxXtdSH9SlQwobVkwFcr+3SgWu1lI7gayjR
5x8g/drWD9iXiad5e8MeD8hJQfHsLZObuttm7RLDERo6UEfKcvRtJfbDMbby4U+e
G6YcZrKCOUmqdI8WEwM3fPTfhXRqoytMZjdel/ttUrxEitO4d07BWbebEWf6dKA5
nePWr8xrglVbvYl2iSvXzH3DnKRMOO4vFZ+3QkZksI5tdK2xXzDlyLGKXKQ0iuxd
L5R5up0HB/XMB8s3JYRRAzOk8tDxUXmPLhL86btDnh2pXxjoZnU9vlV8N33ghDf/
l0JD/Q5rHJdKaIHfAOmsT8NcReWeft3UGy2Z1fnSRyeut4BUhsYEsz1lPfSi1nv7
DY3hvGxsJC+p55Ybdngc8atGaGNJiA3U7H5G08Xk92+NBbbCrPSIK9r94uSA/5u6
w4t+74OZ+L4NFmM5LK+gqRGyFIBpmEEoRGe2ILyfKSqC9Ks4L0JDPFIAgA33W1r9
dlYutLDPfLVjrMNdurNuQVMf3sfy4A7X1dQpCuti9CeeQa7CXzQLarJa/tBqcATP
eBG1ntDnyH2lmp7EaI2UPNgVMds+Z0RujIKk40NyA2zZQ+6SfARSVjaHyuxlS6CD
YuLIGfWa6a1beToRyuJxAUDDlZ70pDWdJXfuCGAObMQq6B7X7Iml9dbOE1+I70oy
Oj8zNOOJ2LKc8k03ofCVfr+6JXCbdD54Z8qb0/YJ++BNj2HR4yAHMyZ0HOjaDZaz
WPWtJbe1ZUf/O337Uleuw0NyZvKef5ERnA3D3LFOZPf+800nDm+RZoGXI0gp3aJ1
r60z/1tWIt0l5G6dFhgSgf/fmQRcpnEIUQTPpULQdmFQI3cNVPOLoJCUaK7PhsCW
e5njaRG1cN56mUck138ay0vJyIlJX+7AWtnqMtTjsml4Kz7PaFP0gcEQQU0LNUio
7udLoOjpYjVmSLv44x4abyGcRCMFtIJSh8ksGB/B29g96Uj+f/rWxRerS09EqGDH
hcVp8QHFI5fp4h5XmgifEhszcdpMjMNVZnAi8SXX0K2sXR6rvVddLj5tIicMDYwR
VorTmUHHX8u9twN7et649k9IT75W3GMJiHFHhVR6dLSAVrnGeQ6MDK7M1tprENWj
FdYJJVgpkvGQSkkD4rEJD0QxXqgs1jB+9Iq/tQ8R5O2qpW21/bQ99WKhXc23wNZn
wr5NSFz0r/hfYKW0SgQyVUplZCJHXRaDbCecZe/NK8KnXSZIndqytNCNHU/3aPIy
naPqnN73VI5XGF1dWBLR0f7Rp9gXXS513KZdF5aWCCrOj8DKmkyVXdhz5NfxJxEE
SyuT7JRU0qjjdHkaaozRVgyjdF9xA+Fe/UOkOwfpgjAx2PnMEvcFCLTcksoe33Fz
wy/3lwxAb1mveqy24/y0/ucRfmOWqsZiYFFTMCVEZu0e1WUW6hzxzoLV1f5qUBQ9
ckPFqEtlkGXLt2dvIL9fdShdnNkbMMBsAcwMvvr+Pk6Oc2ntF2+A75KC3l3qgaT+
UcZ7cVIW8zd4gIPJvqJUJowdAONP5GQe3RmRXEI3aaAXNoDrJOylNHWLmLmYk/2Q
JQVhO25Un4jXEJ2VragRo6nh2dFOdNQ4mXqWV27MAAGiJd+ECV3mCDm0Muv1mGQc
SIy1xACSd8RI2nmzOHMFRWMdWjaoEOiuvd8ip75EXvKUZe/4ydf1APUgo+sCB9Qz
Sd9d0hzaoIRJ+3GmGgAuKzx581SZgf2boykuFdQHUFO4HgaPVPjmjSxV57r8rSme
Uo5rAuq+ujQrxoA1LJo8y5YAhP6usEy0b+UTNpp7FdfZlQldtjY85bofJBR1/Xaz
I4nHWxzElH0NapRnRymgvjVTaIRi4+y2ipqZWK+1c31vkN1O21Ftd2Pt0OVywb1p
GwPeG7He1ocVceVAqZYNhBtAzhyaFrbI8wJAgcrKXheZvTiAMYMI12yU0cI61ad8
M7bfbZA8GVPmiqkNESZm7rv2QzQY4R4CIf7fsYynfPEKg9FYSMzQmrJZhSA0YbDL
0Vf2Rp8alPtltDexEfnW/IUrhnqFoUA4g3V9FllXtPHEMtvKzia7CD9NgL/AmZnA
Kqrt/lAY8nj//0/3utyquZXX8TCUUUDFlJ/haL9QNjMr2ghrdKWu6kVL6gtuOmsL
In8WJvCNqCVFMAaty/iGpNj7jHkhs6rwuvrIpsGU2Yy6NwQUbPKVGqkQb20usA2i
j9phopqiXYTGP6cYX2KZWRGQ9VBOfHAbKRvHE7Y7cjcQ/1i0TBFV451nNoQs800b
Q3X9DG15uYrwkbxjsA1W1rDFUnhRn5ql+09G8Ug1WTQhWkaacGh1LR+zOsXu1dOF
awGBQizOTT4zOezvxuet0NIITvtryj6TnqWwV64f2szkKRJkAJRqNSUI75tdKlBe
i0Q5CHKwOn92fUQ68EZiYUwMQ1ZMkyRXhkT96asEiBddk7AM3F5Y6gTBsQPvZvbP
AQhKJgtFmgbTz/3Xbwpbv63gKHvGtRWHTMsqpI5fUEOoTLSXBmRSROc/6N0uDZhS
AqVcZffdXkYkLNv/5zad4erGagUFBDI/QjPEPY/5kg9AexHUuFB1Wq41ml6TRUWZ
o/WVv6hqgWdFxOAzusuOIX2/ea8QF683EPBKgSp+Ilatfzp8H/QNZq87mP5hYzOX
1HZ44HF1qcH5p64yUgibu0ZwRvHdYWd2uUPMO1G3RI5GGc0UpJ0SPHUrk1pdAOgL
NpsnAl1saZZ+vueNFPZCP1x3Q0d77PsVGjs/+ku7/12ejGo3juqhhLUDwAFlE/8g
KafCmZGY3Uz+W6725YLPPwC/UDLdZ2YVV55wbHk0X6bEr5Yyvtdm8DZb2y6qvaux
gRISGqCzx5EqgxUhe4n4Ac805PTzPH+/HmDDtyLOoGUHXfncbLrhuuFv4lSVTQpY
BWtDr6BklM3wNlIrvT8fvMre1iwZYDxcoH8OwZkzPH0ts5sL1e44k0xIXx2EL4Y4
fephDLYOOLn3HHD4QDYARjeO+c0A69TRFrPwTaVsa1pTUGTe0BGuqk2M+1hXQX0e
hB9napBO780c9gCjgZMBFkvOKJIX7WKA29JEJ/IUxWlotPU/OV8XYQeggJZrrnZn
1QgzwWgYwa/4M5CV7y6c3PHAmJtIHgG/JubDen4TJcrNrcnuDBMHl7Gno4cOw8Jb
oCldMs+KZyKxLJ0/W5OwrNmUSioh13lFfGrM0pjMvwcJztVhZjhaeqQHPQQRqKET
NQz1wJVlkxv++8vLtk+n4S6bqsgbigx8MuJ9+dKVqqxe6Fqj0n7ChdBbghsjXwMT
M6QFtTd+eQoz24vRvQQXZnMwEE/tCAMTL3fAB3HOUi10d82xJ8kCuariZ41dIPG5
kbqmgqBCJKejNHBWZoG0TqWx63dIR9xUov+S1BQv/LO+XXJqaTJbb0ehlYlcbJkj
j6PlChrJ5Y7zDWtbLAAJU9hSv57LdE+O3pqKaaskZhfJicThIGNLfe6ZckLxzYks
X5SAy30+DU8koE+ev2V/ti0rLjLM/7g9JP0iWBdugqgq3kzusiHGembuMhSfChOb
t8yP2uZKz2mIcEP3LuaY18kH9OYxHGdr6bCxUS5abV//pwQXMwzozv7PJi54Oebj
9YQSf0Sir4BEXPGsyxSKSzW2DfTrMiyUuWexKmGWQXMZjahe/yNYhrHsfThgD6JZ
dH3EWAp+8oxfsAXIG6ne5KFWShOWUcIhoBo1U54WQqbl8QD0xfqrwjYqKl7KzyYn
ypDDLJuZuAc81q3H/z7D3jRCfSQAYQQvN40nn+zgo8ltI9FWFOGWsQpDaG030YTt
AnSHdugB7nwuSlhfJIiv+PkrCMPy2NgdFOBPFJufUqiO0EhwNGMkUXNaGO6Cw4H9
r+NRzcaMUVAF8euyuVGAKV8dzUrnRQtihwqcJzXpjw2AFqRiEph0/cXpev5A5fNX
+wf0XhJMyFTxM/oDdManUjOyDk7zxgLQnqsHQV7KWAA1pnMrD+ZDvePSuz13N9ZQ
r/K9lA9eE0JFrl8h+wcgJNyWwhX98BgZ+iZWiVE0jlj95YWcBNQpZjhg638TJPfr
dxefNBmffEZqArGRavBHzWS71fWzDCCFVwspSgA+jPP9UvVgV3JUNMCTheO+UgQY
+QiHnr/N65u3WzItOxRIZ/mvl/stj8AY3Sm+bL2jcj0l55OvpJ3gDOELjwtPoMYg
DpHBmq1KOM0h63l/dbTdN3m0yLaXGM7kdPyqoujRbwocRRyge/0ygDXeRDKMvEHR
YTJwVe0fSgz+GOW/1S9wsy/dD6lwDsdnwAbjBI5NM5DI2ch05IZebwqb4ICtO2gh
wF+cSmyx3z1tLFlrjLa/vT/S6B+G+WPtcZHf/qFfu9jp/bcfGFN2jlq5+AzheAr1
ij1cFctFzvROKlisYtKwEi2VKXbMPWryF35crKY+J1gOquenxXLyz2LXjJfjm8fp
8SmqEhgFdwk9hbH+D2rrzws0luyLiRzkFwFXiMm449aOEZgE6QeyFrtbfiSLAiTh
0gbFB1qrFiSoW9E1BLYq803QLf89DsDBsomG41pNi8Qt6CK/ME8EFnXNhxSgk4IB
k4DEIslrmvoiX2+2I/w7WuqbPtHt5fThXHEsfKmjTAXQQ4ngbX+A1+mhJJF/X1Fk
OnLgJFYxEUMexl7XCZGDCEI3nNGiGxvH0vK9UBaA2Bb629LQ6blMPRUnxl0eQ7sN
7IOeznrl8CZNRc683IQUp49kjBw/AOEg+phmL6hvcBDh2m0HN7Ww1ohA9rQ/IvHh
RCQ900IBGeJUt4l91mJR8e7VEpNsSxYvcmM2zJpFQXQXBpgBHaND+6h42776zsIo
RYJqmmuO1yXM+bKUkbQ8PKoSvfnuYwo6QTJXcLigioMs07o7Sg/iIhyPAu0yBBRS
z3OngDQdKA0yYWqvstjrwHVAYUFUOP1wpGx4p8/YNaLFM4w/vzjK+E5T0AZlcwEA
4+zHH9fFVsz8ME5xkcK6WvGBV8j8rWq7Qdw6Er2+mB3YN78K6FtTBgzUVQKTKC2c
f61VfFN3YOxP8jjAGKM6Lh1t5WYBp+6EmbROR6KBSUgi5etK4MUXviW66GYgMAWL
banPuyXf9ck2qKb9Hb6UaxCDZCT+rmbtZfgdkfokhKNPn4a2owpMA26oZMFfO+9z
Sa7+LFBF1e+XPLP0liLs16TEiT98SFzuv8ux5TA2AM8vO45b1tKujflgqfP6+3CU
9aOsqigxe3pLMEjYbVyoJr9K530Kh8HkhIdToBchZV5pda9GSIhVR3cLyWiijR0l
xfzq99VNK4GoIesGBUKcB+t1Md+k6O0bMvx4zXJaaPXstLN4UtGaFEUQzN21CI1v
mfgMVVZpluuCJ2K8EZrUDVtiSpINMhejDE6NMrc92nw4cq/2Ggf3NF9kcIt1JzTn
EYGx0gf64VfSjhrFmtti2AtFB6EgjEWbTvpBpv9iKuN34NYkjb1eRwHu0F25/Rto
nl86W4DBZugG/g5lY119LyKttgU22Tm8UX8u/mk4+8TAVn8k+oUDmxxQ6/aSd+aG
ijTESQOfl6CIXM1ooNOIsY9YHCUMpWZBp5QbGpXMcAo7bq1L3u7jZFK7kjASE0G6
0LXodp7p3v78jwzmcjhCJyGPFbmbzSwNaEJWDkZfY8hfFGXhRCLmnKFZ9NugpDUz
qqniD5fet5OPxfinqaJ5H5xMoDYIQeIA9zNvkvIViAY1SnizdRKiB+n8gpiZHu2T
MP/JnUdRnP6GMdN9zA4UVgp8DTobweEibcfAyjyg/wtE63oloiREmYZkrzlRElda
aNH79lsHaXsj6j1CQlcEx1Dr6oRU1P81XN/i3HA2IJIqEdFaInm5g2XNuxpSKoZr
hyeiEYTmqYd+cLTBB0q/yvp2EZRASj0J/Z8iyqVLtfuXMcce1AZQDqv/bi+r9hXq
00d+LBRZcq7txan1C8twTMj805gmcU5dp456JDdcjKr64RurP+viUwQqLc8ycqOU
e3+fl2QoOTkj21hWGZ1IX0QhbOe/IfGdOO8y1+h0Z5U7bdZJP59ZcySFcOtT2bEq
cfiQQNXvYGfziOOS2wglNRJx0miVm19p7ly88qs9ZFjSLfAcxwYcXiVBjh+Ilz2c
fGiwH2mOHmLWxd+VRqcLNHgfldreEChrVwnEtPs164treeGV4iEv2FN1YnahhEz/
Q2KKgDB6eDaaP5oXGeSzSS7l5j53waOBgEZofMN6NcX5vLbEAuniy+BOLM6rr48W
c44Okt1E0lXQR22n6PzQ0/2iHh5l+3IFOUh3hAS1Q9OhTxRA/t+Me8TW4wGRnUmk
r9MBWe8cl7dPbOQKUJAcPT5Y3NMhMGGIp4YhY33tJGUzEMa7F49kwU7xLOpicH1Z
oqNkksr6hfWo4noL7Pv7ifLTTsmutW41Tbq5jn1KYiZS4CgVk0ZtP2ySUfqLhzBc
LeQLQTyigsEUCd8h9uGhUyJfiQCCo+4rpSA+ZBUDBZDZ/IguuWJKORtyZlzwidtA
7HVi2gX+qqoDYEEMBwgOgdK9Zb0TXl8Qbas67D5WPHl3y4j27XogOHnPO5u81VQW
jeKW8B/hZ5h9cRhDzhx/C/pSecO5xQzvCHYmAJLhvtO7bjnN87rB2HHD9dDj16Yq
7LfDyz83/MYOLT3sbGOsDoXV6sIJ2q0BJW07MuDY2W2mgW9lrVdhCdLMWV6v30Xn
G4kRQ04WPRbRHaOw751PrGIjX9ZnBdzHpfDYMwrNwW5IpLZ6hd9ekRVHsPW4lHI2
V1j5gXxhNIO4735nmKRQvO206GsPhmLlOA4WsxzebHFLw/3a/jnMh29Hd+ehqrbJ
/nWiKrfz0lejiL5/C8OVDDT6GNZ3sUF5GqIt056zXNRXKiRvESvrZzuVzQS+bgel
LobEsIa5kR48ZF9hernH8rvfPcXD2ctrMItCpXYv7BiVCGtAY3ag8laOXNWI2tZX
3c1E6m2kWbhlEEsw0AVltkm36nV76xbKgQaU4NGaaHoUcvtMsCyZ6y/TOxyUom3b
I9mbeavOL2goWkSOWPHy2ioBx3t0RXgbIDVUQqbnTv/N8daCp+5JRYBxuTEVqUJc
cUZK8iBO1NzkSh4HU46Mc1xJBbvF0krkZGmUwn3d5DPoQbvmdto+QrKVnQ4vWOr3
1MJ96hzCzk5I27IzTJDfntScFa4drdQQWXcHWLG9yAEc5iB9gxGznkSNjnG97Pag
/9UA/95UNGc+7lBFIGr+oZmHHJl1S7nRwb68xxjSgPJLdm9fQjgXJQTy/MqRTml5
y+yQNRvay7hU7Hb11M3RPDVm3WUirz4WLWX9kRHvODTWBt/CNhi6U1rQPibFz9Bh
3LqbtVF6RXEw8EuXd7JvDetOdoyvt2joHzaS4Ov4dcZgL7fiou+POjSZRB1kF9RK
qGTrD1aVdajoM3u7RJ5NkckaPuDG1ZGwM9KVRU4c8rCfFD3voIWo0E80zsTRIDAx
Av5lo5l6naskEp+qJ836h9fgTbR7ZUxwijaIozIRToS6NbdMqB0ZU8NGhf24mhtt
cNRvO9yPQ5AKyIfdxDXBnP/0NTq+9uzgenwAKxy+APgrEL9xiTCAKJT0yQvCJZna
xO9WfvZ0xd7NV5uDmQ2f17kYfNGtepes4XACrIv0iPPjXPCWLkPGo6Qe3xC7zD68
1YwmoBjf2aS9qakSlxUacV+m85GfbI38B3zRYME19lKaZewVpOvUUIuCoDaBA2Sg
e8J6YxX9sexQGiin6QSy9NM/443EwC2rIbu3xzwAc2ymZOFnHm+lQx3mB0CAK3ll
exWzU28P7b1/PNko7N36846BJnHf7N962g/rxp+0JIZSwV4gyQIa45wA24INeMxO
+a7dYYPvF6AkPl7NDuHyPh1vYuL2XimFijAduLQ7vRPaEUn+4544nfuKmjFSRfuT
6ZiZeDhxgDxHMtuTjtuOUfdmbSdu/GLpMvvoYkGAUe3pJLiYM3dELI10nuS77YxW
bX6t3mjd9XTW6G4JfZNI6o0tFhL0VIuCME7Bj8il5iYoz399oNDYUSUHJ5HZBV6u
2WIT7g7xsIKvEA8J6/EANA62RFE6AVurlRDyRBPNySlFUly5Sh1/k2o6y+2J8mBn
MF/wIo2GJYGfxROi8qlN11r7rCKGKIAHKlw/Owd6hPd1bSw2dUl444SEhB0kyIY+
p+r3hLoxmQ9Ssb+lnr87b4Wt1li3gbWlAKwIXRg3VjJnU0Izp9EVCHEhYl4HcXJW
MZwpX3x85/KrLMPRjFViV/RL1KBV6YizjbRbEynMJQyFbJAbazvyQHQA2bNWKcdJ
0qG9QGMHBndKw5liU2f4flCO2sGN3tMA8d75tMPqPdORjztaMtNu1CvgJoeG0gNI
3PMQhmdK6qB7/HPizV5tMMQA3FJ3kAXG2fYRKhXnwNNvacPeVuTHZ2Z2ek90I/0f
VOAEyZamv0VqMfoiIO7W9qbUONUCwTXvShJ6UWEWSY13UBGT66R05Dmlk2yYwDnt
91MqMxgWjlgXu4unKYriWidNUQXx9jfj3jf0ZitEgcwQnWfmEztknRFB0IlNONco
QpNhj0a+xj23kLcJVju+BIrpdLP1Dq96f8enhkfwNX3f2T1sXr83c4wqQdlq6tnf
CTz+qlvXFyd9Kb4NWy6HRHFiCX4XCkhE0EMsWgkjtZ1jgUNuQHvXLTujHpgNr0GI
2OocrNIpZBHEqbJ970SWYbzG7jnFrKZC22LnMo/x5CVhMOVf6MOzYrkwnzrYJpg6
pTNk2uoK7t+UEZqyBHUql/YXoCTx+GRDGZAMfPbhHBPwQCM8p4vd+l7rYE1IqXWr
/BNNWKCj49E3rmEofpSXllhTM8fW0+G10I6hqUOuhVsHKCu4Gk8cNV/PkxNcFmuK
Km9k3VgX1V+kfVNXUOt/nw0EMrwxG98QSyddEYKuwXiDcsOdHgeTGrQZbtU8hQVP
WoAgo0RyciF0OjVGp3YXmHRGaf9W6b7/a2OjHKoEw3l0PYrBlTtEhT6GcRCONjGm
cbtY91cs4y3AVHqL8gBBTL2xOAb9c9qZyhHOjTp3XmQNeLbaV6stxP1ieUESTbGD
86yPelyjWQbiSFoXZPuDph8+aN9hDdWH8b8eDTDlpJh4dJ+uXCUKTsLRnSDMnDXw
9N17ij9HalmAglgrmFalzrOZWiGmGIKxOT3oGPzzX0wh9EKtNb4c+ZDXXwKrS52R
bqQdWQqPXLmZgR7fI2cgYmsKpD6XCNB/PbDdU0XVIk7qGow+UtcdzY0+1lZap/GT
bgXgH2LSUtO4aC0nye+svTx/PD+zX88UZFnY5CSeOgA99xwWxNOhNjNdX7Dn+EdN
BgpDduEq0mUobxA4zL9GJaIxERH3Ct+SZuHRT/aO1s8cy3ge0OWdOuVKGgARLNpm
1BJCAS6qudogmMyb5bri/RFQRifmse+lhHdjtOdN+gt2xkSozszjyVhsIaeKmkjV
QKDlrtxf06YuEAfbPYyZhFM4d0tI66SuWKbUl3uiSv6yFDSeEAE0B3MWokHDW9Ez
17QhCmirN+NzFgF/roqj7wWntMyO4PSLu6EJmGzuwQ+ULeQrnKZx2htDTslRWwRh
1lzUIW32GRH9n1Bd6rwCA7bAvzeFXk1nTWf7BpzrV2Xj/Zmjt6W5Q/V57ZsWaGoS
ESK8V2A0cbDkP1FdGk0S3Ys/EccjxswZhxiYg/10bXm/kSi6JLbVl0U7k3ac6qmx
gXokacT/4o0DgMyQ+iaVp8QzHiIdEPkHmOxCvUVtcoQkyiLTYJCr8WnGrvTLh53w
hVQC5UAVwHhlTK+yHhKTOI3ivvQiokYoET1nGad6PUgRLy36R0XCav+lsvPhmdhw
1uVbIKSxB3cPGyBKI/EebrRGkirhgZBwZzEFSEWv+kce9Ps5rJkJmZ7V+5Z4MQ85
xquc1VNZNlRUta+IyGk28AlGpZ8g/RQBYeFaNuNtaoLeofXrCY21hh5wjrF4PNjt
7mVL4WKaEsTwq1jpGhE/5A4C7pdyg7gB6yxG0/nIur0MxLt4cLV9bCaGWcmtxkLW
r1jt9Jn3FN7ehNzYQwSKY8V2Md0FPyhD88PNk3D7lVEa43hEJmWwnxHNWA3dAzVx
XRop5eN8xsBOoyiI3wKz9e7d4b7w5b4EB940sN1ZHuLt46VDJEcSMGA3a+zWochX
NebtTneXPp0OygjHB/LZgr9k5divLgqezDwUYkdeUeefYjBaXcOmKiQ1u/UteEVC
7x4x6ZwWY9yjkDTxXDOo9V1d1dO5JzRUJNTuqBJ1ZX8twi7OqfEEzMPGXd0l08Cl
lBWw9NtgAmWu0+oBBW0W1zqN9taVFyJN9VZZsV2N/SkL6PbhRzY0boAQE65suZYx
ogjKvvFhRuukvEl//Hpv18S1RqM6V2Oi9Dztkcau6td18yHFsgxSp5pFtKXaK6d8
vy7y4IgQ3FOfyh03eFwfcTnwCFjw+ZDzST5JYDF3m32EMsIOqCGVynXLxd1HnSvS
TH2II8SI4aw1qJooD+MgTJQmJRRvJuoHJRSp/M4rtvnPbd6/3xUMpKyYqZnp5oCP
X0+WCIPhP6hyjyX+sEdVaVE8BU/50jQ4QbthxJP9w2uZHsDwd0I89T/ex4FXzNuf
MVkufXdQE277GvubL+zh6maZW6LK8jvU4lkhrC50V9bArBiduFg1Ho2W0rETB4LA
oLuCgKu3ld2vsYwmUXwGM2uj50x9BQ7WBV3iDkVY1aRofvI1dp5NIBfgVDpW8cHk
iWgMirT7eHVBXZey8Rxum0sFcSjB1UZzSpC2jnygvJb1QMtDpwhDNA5I22zXLqh/
ymzV3kZiSosStc7epSNCiaEZTcqFcCZ6Bd+Hc+ltGdWvTY2BmbRznHNGrs0FXzF6
+8mN7jW0DvMz9olcEBksYtO4t6EMaJ+BpLhKjnBHq8Dl1t3yj9mjYKTmwsWEv2nf
Iw1vz2AC5AOtAg/ulwo/3omOwqYpZ9sp3WCbIXJ1InV1pL1U2QYHrqSxRAJtww+1
x4dhA7YEl+oJ5TdYVc5hqqlef/Ecfjp/P0rAOOnaaLxvDwsZeRxPMi485HtPirbT
x8UavutUNLF0BivRoGTnnXKcW9ihdjZ3T5OEqF3Fn7ACSWkcEAVFDMK1By9hgoqv
rr4rkqy0ArswKd0CM9+NUjPFTpkeKrAiACXdWFmcI/cWciAQei6IiXdnOssFfQxZ
vIWvecKVVX9uSexmANyntWYgy0Fqr+Lo7EXnGiixpJ4MdniAkGkcOn/7nl8qE2lQ
ROSU3eZdBJ6mxuh8HzyF+oZcw2r9afsLg0pqe7wz4foHA/HSVBCEtGyFmWSqDKBl
WHqxzRBFo/idv3xbpWBBKJv/OH3dwEjP/NNT58ESzU+g+9TrMjl/6rx1uXI6B0xh
q+XNS4XHMTR06sPgU2FhVvWhzEWxgEwe9djNHxgI3oWjVWh9b76t6OsjOcgdXJuF
rM3F0I3orCzWiMDnf1CqhUEH90d49J5Bsk21AciPgl+sV1cnTZNBfn+YmDEgLLkJ
XCRgLZWhzDjZBbXuzSRvFsGXOgkXytlyEwDNGy0cNXhkCZDkg9ogPkLXaevqySIo
G2CeyWKI4pdr33Y3EUjQJGO1KPo4T0thcfhaNoT5bMILby8eavSZ3VEhx2pj+xFy
Qz4jIt/ALM5dvSLLS0zE7/s70Ur2iP5782vtuMGLZe6uVuQBokNU/3hEgm+yP5ZF
3sRFBb6GFiZsMCO2PFOTEMsEvZ8N+3BovZKEwl2q1LeNA/BKlY8NlsBPWUahw8cT
RBPkzzmwU4r0I4xBGwnvj/l4czBPINA59oU86elMLdxyfBgmJI24KdPM2TJ7RKMD
VJSvGBi7lnNArO2UigqTB1RImEa7KYQbQy1GaO0tLHXB0Kg1OPWMdkEmKEdQeOge
HK2cnKm4qqMWKWWCS+3Z037OjDPi8fPyWcObyOZSe3ttdEoE5Ahf8RdcQIqTJeSf
umJJR8YX10YnF2w6WO5nLBEBQVQjXZOBwjPbTRa1mje7u78qbwAWPIv7vmmByFFv
lcGI5fR9koVJlTpBzqzI7NP6LQhXMKf5NUQG/YvaCmg4eZd4Owjm5+c826FFIT6q
WRIGlEM5jO15d+F4HfTmIwuMlgfb68kq90wtG9dd0/R4knuKe4Wxue9VveUId7yA
jD0nqXD797L16sVKY5LZpOMszfTtQJz1BjBu+tkWPNuSb0s+eLbO3C7u+URsw/Zq
EZ9jPyBDYheGdWT9hrd1jJH0yVvKK8DZJbxlLTU9xd1SVr8CBmsoYfM2hRwk2mAK
LHI0eKjXFnVNLxu8L/phurFA7iphv/JDWSHIJkikP7QFSUXC71TjKuiJCMa2LHpO
aItdI8cFGE+BIqYiZDk8bki4Qy/GHLxEvFQYID/1xMuPVK/HipDzkFBluziGXb3N
Ov2T4Pdjx1N5Bv/zFR6YN7Twcq2Xjezd7cjQxaT6KDNQJNLLb5aCuokbECS7MUml
/EqhRAqpiUyDoeGC199tvXHVGFe/K4OmYPwJrHVYwPcjBPF+epSQ1Llre6zmM2HJ
Q35XjxzJNz1965JTrdVZKg4FPtK3I2n8xskq6fAukfeKysOJieVXE33xCy2F4QAC
3jaJUoG4qngqBAcVXmNueO3JBZh9dNIO7bjBfPdgpwuaX8+0UyFVK0U1UCAWfO58
wqjXm3lmHn0DX+g8vr+ngd5ERb0whlTQy43mzsQY1DOu8Rky0i0NtiTDaheED4Mz
O3rdVc40uJ78rGd0D+Lc7KwYnJ+zIo+x718BbY4mSMdp+9cWA6KN/ifwMadOKqFW
vjmYNy6WgMRnrZIYpmnMhoZ6LYVmmz3y/2OMUO5FhKOIuxMAclwc2OnyEP1HxTg+
Tv3WNxM1rm2dMudXXAznI1PhMR/rq/2+hsIPISxvfjb+w8ESbL89Vg76chc80wVB
UGjmcyJxWgK10nvQogqWI/dVNeBqa7L3gm8ic/W/D10zbaxXiz3CplKUfBD9GKMJ
pKgNj+fiC3cXOHIz7JIN3K0zOJrRZhwsEq4StZWqfu0JFP2a0cC6ewZag33O1FZo
OYw3w27+ukmLbOADqOLB07KX8pyVZpCxLjK7o2Q2n4s2HAS3xMPqJhgk5sskRzdO
oS8l+xbPlkvwszoHiaNVCltLNKgyXaiTIeCw3bF8ffBx7MxJIvoA0JoPFHRYu2Hz
JkQJ5ICK3l1FKx0JjRT79xdvCcJLvlZ/ZOad1W4KATUCvHlNB5mmqXYn0bJiCLap
ApoMUoC1u/ePAT6G7cGhIvxtz2Y9rZfJVXoKlSeES7YPnAGr4/eK1m0y5g1kK4A9
y4xcspOTq5Xnhrz3stHHubd0+PFNkILKdFhxM7tRKEHeTEYFnCSHZ6v7Siqag4gf
rjOPMycfG1QBjJIJeYFcn8af58o/n0l1sAw3isQxO0y1SEmGgt7s/duQRE1aK7yN
4ch7yTOOtqKhGEfV4vex3HQGY9JzMLeC7n7CBAJUZHpUuYI4kGPKAQhGgPCs1fTL
hdDXwQPE+udP651d5vwnskywN0z8pmRYRyyrpJL/EIWMMkMn5b4/TmU7j3lOweLz
cMD0MM+R+caxKPV+Xd6CahoReaQQW/p+gtWUuviNEQstX5GHaA1KC/ItMm6Cc97/
NGyLOWEqEXU5LSRMXCwi5lcMG9qzoXtZ5P8uB2THrnI27l+i4B1H8TIAeop4AUGh
fzprZi0Bcv0ZklLtJT68WjTUi88BWJqEetTCNx7snev49E2w6UcXeariudMV/dzv
19Yfl32uMZksT6M7xud9j92kgsvbiyFHvrpcU1hkC+VFrozR6+CVMf53ogkO9P+R
D75/bdEI8tkr4MQ8e+Z6EQ0nj6b2bpQ60S8ik0kG50p3T4XhHGM3eFla1VKq0tG8
odVl3yqjRT2utnU0aHn0LazUN+y2a3xdhqn4u24NE4rZHEMkyUPIXQvaTR2dST7D
0LFg067GZQ5lDMQ1WPBmmJJmvhKlz16ekQmaPq0hIcsCjBIPB5mxx28vg31LNAZz
yCh4somY4irngH6Ajg8+HrromNFMEslKZbhBaNjNQ6ufk1XkxBRiQuUWNlYJCNZl
PyRbfH6BBAcAfCSuBOGLTqTxUA42XXkilkJo8gbcyoFxFEVxxO5e+kn7hsjInvEx
AYvJ6oNhXf8zsNtsYFpadUfhhIybnfAzcYisPAJsS1yM7ntw9/xybrgixLJZV3Ho
XdTyexqe7g/bMLjoO+U7bRNnh7n5HkQB8FgEH/2jMtkK/GNXGAvnSzUYgzeTzrnb
ck6cf7zEYYystDWzHrbyurkOyAkkHYPUEuUUFF0l2YamZIUYfDWgaZRagw9S3hF9
7ntOccgubhla7wqvn6d+LcpPudReaumzhtMHDV/pXm6h8P7fwfvBOGDUD4c5BTZl
YQs/RzBs+Wyj4UqcuW/j8Cj2ln2Hflb19wD7/wJ3Sbr3fcqUtOmx3drla/1AiUVt
wIbXfGG0t229x5QsFQLFfj/rOQd48FZdQ+OxsVic3CKcsxJSZ6guQ0uQ4xHe8ZxE
ZGnFMy1vULGuQ2cIiD+CTqDwhD2iuh3nkCmDosytfsy2+zkEZlZ9DNehfPiMibdb
TZxGqrMy0Mh9Pbyr286s0H9GOmBbhYdwnuZXjqkIp5L1a+TRyr2HKi5ihTJTqQ9P
ScPTSkZEHxordg0QoxbIU1ic2Irg2qtiKhcrDV1JpBUKYffPlRqdUkqf8nUH2yUG
Zq5mgg8+s00AoO5pwmcu5jH6P0B1REqztVwFO/qgi7vC87cAltXIcyjV/AcX5sag
zQ9Lnse3H6ykUM8rQgHI7KfCU+GfwFIFuzLGn5n5IJ9mMehSzkhOHQ0Re14DR7zp
gHJpnHDDvnVBBU8fW7EMELB3VSTsSefeWLReLKqo8rO8Tl+vVwE1e3NcSU/IN30M
vwRlNsYqwd/+ik2FXeCML4l6UlU2Opo1Re/fbCx9DPIPkoFIaw4YUD0GRGpDgxxL
il4sYOPvbEwdvr69Jxt93bHDNq1XE1vf3VIwid+sOegS4w+kzVc+HanzWQ0PU8zo
WfkYq9NIRnlhr/8T4Kc5f0cpBt1pSgzjprsnAamXMNmDByCW8NBk5vsQ3zZdSr6Y
WPlFcHREdYeQKqU5nY5WsFZ30Q2sBhyo/oN3y+msQ6IdYlVkUc+GE/+fqCFZJQAI
YDwIyguz1DE2sy2nO/DmYVxU+4qWFTNTET/c7iN1RpcKl5LhGbFwoFnpnM6204fA
O27f85cB0UYByU1Q8QTCsgTOuWG9ivIXI5wF3YzaTopsZ+uSZSEd64J7xuNzYK/S
mx1PMwXte4LEde2hnLOTOgLwn2iEP0kfyu0RlGlaYXWKFbx02ndr/evEobK7CKHq
ktdJOGwsDVwfYR+fpclmaI9S+ypDFtQGIJJee8uPGag7f+SShsKmubfGq1wkCgWi
I0RJmYxmXYm5qMM0o/2pDXmtvj5ofYLE/sAoG+2b6xH+/8d5T84J2Mhc7Ef4HQWS
sRYIzMh+KsSoJPSDQzJ8kPTxM5foZVgEP0Uz7w30ziefffbJd6ENPOQs1wHYqqdF
XWoWoS8tTnTeshVfCqMOHIsIR+uczO9yKKZRUDUOAgEB2a+VnVTYTp4xz4e94u44
gs/ivnmRwko6+Rkv6Zup8oSE1srar1DJD66d3ebQ4t9Ep9/q9EQabwZgBNtZQm6L
mDZ4/jFx5oWxtSCPHpCcNItq+vbIS4GSKPQzG4LzfPyXA5l9yPgvi/KhZ+49I0Q0
+DwUv1QrUPcmH12h0RTgc/eXpmm2Hk5eAmSYEgeZIVQCvg9D7CngMsmyWvZBrHm6
HcCYVbcVPcZ3XtgCJJ6If6LEOu4z7aR7enyVtpaOnkB6Iak9u3tIJomS8f7KD/Z4
oWqP2apLOFWui1V2sMI72LIE1q1TdrpDSYZz8ymqWtPT+Jl2ummSuxMiLDR1Qm9v
KFmMNqYIBAJVHZYZoDKUyXRepCNx8rqJ2TK/6VfiPhY2BN8k2knCqDdTSYoKT6Fy
opLz/usBpB6dAOlwNOzvsd5lc4ucgflQAJkCz2/JlwLqIBT+AxBNEWuwUKWVl1Vu
si6ZgSsROmpv62qVpOhJeft+lnHsnkywiWUbxiOzTdLvTkoooQwoz+cOcWrAOWRJ
WXzTBRZy4g1RznNtxiiFVofnDbPe6KLqQgaWLu0e3qI5QU4nQ1rF6nFIPpukQ7dN
qxs8940ctyN4I4TjDCN1hI30NLLbi1seKoQ4Qem2cfApmeZ+Vhfwcz0iw5R4kY8F
6TA7TSCS/5c1UVCVviSXQ1VwEA9S6A6mYFk2vOlNeFfidsYipSChGmrBlcbNwIbc
vAr+4Fdyhh2aDwdjXdx2ZwtwethGUbvfIjnbjBrGfVQ3PKhxMOTIGy5iDju6eker
1MkzfXyt+XZ9tR/zYx0RffemjTw4iYsWLpJRJIDae8eV0dlOQaq3mYP+JOFl3RqF
idlMQbh9ZvpQX4bBWOX3eF3HWjrrTk1JbUPv1oLOgDUQOM39qMOMIrxYIgOtAj0O
+xVA3mFl6xUskDF3wrXJ5vuoNpWKh1nhb/zdx2aoAipREA7LiIQtZ0lQGtvnh4Ha
C2nUJDczOorEtahYIcmvlgxVepKYFt3sY+hhr45xjFX5Wuh3Am3xJemxfCD0avsS
s4VDXJONxLaG0XVytmEPgnZE2YUVKm/DBvoQdcVVdnM/hXAXObDZAwJYq4tBzCj/
0FPoO1b1jLb/QDWAJtaA+rUU52Sd8AYfwwctDT6Vt2gM2DFahN6xYA3CBVsv8LdQ
uAMvWgICkQBm0l+f3lyrraljmelJvzbronu8mAUtsZhBhVT1Nx150Zua4fOEtxCZ
ry5fri5T47XNRB0hMmpNNRjQH74kTjiAIWH+jfaxIBstdqVU1u/qp9+VgOQmmiQd
UfHe5+DRy8hD2Mmwx0psT9S5ZRf+uxQsdtpUFNqjeleJCfSaW9CHJoa9Z18qDu4I
xjzHaH4BC1wDb5weO87OKh47K8qHf3FfQ8OEQJawXJ1pHQQ4je/uf7nHA/AiaoEe
sjUMIy6JcfVtw9LHbFMm7pj0DlHwWOEqKFb8XZQJnvVM++PtqcHRJ+kq77lGW43G
bKBmXChNjo+wFp6ys+PjdIYy6KlEARxNr/CTzQHxATwT9ZFfwhDzDiB5qzEbdD/P
LV1CE4mHX/ODrnNEMQj31aaRwnSZwW6fVCjPn3gQRViVHav104khaMqcwu4FOQ3p
ouS4YIeK947N7v3UdKpJQj4e47RCtEwgcg2xeaH7P39U3gY/Tc3OUqwEfTYRB2Ar
LaJ3AZyLViS15ZB92uCfFwOqMxEvJNEcHs9B2M22WxBrUhjdnbZ0e0OYWwQ0jWMv
zH/D5TqzmDqRkaMaHcdUKzXqbgdaXciYPdB/uyw5onAyvwvqFD5YrEZqu9BL3FO9
ROrTdLczDozkQHkDQnESxtcqKKVE5yZWgaR18eMiFeQKpDGb47hkd62yZr3qD9KW
HNTBsPs5sVp8volLOEIYb4fbZgRRmJJDaQkVTwpW8gBsGauUD9yT76GGSdOWP2Wi
0Psa5Cfe5DLuN9cDPmC2cJs75SDO7VPSJj7FTVWxWr1uSpC+ImPmuyJBvWCbqxA8
1Hky0+In3+CK+k7eGODivi/NNNxwQzgiDdZkLybSdTysnK5zpiBT0PYo6+v8rc4R
7m/nwDaXVvOzgb3PsjZWvLGyOykZomlL6hBBFYlpAGVNnW2A0HguPA4CtEG8FPJy
2brSrfvKwJ8HBBJhs3k/9YbAF+kbwiwpPPrdfup0GzC7eGFvdpJyiEx7RgwunBFW
4pFrfk8iQOhiiKJnEXwJzKf9IhUvlh4CiviZoke4maqbl/gSx2thedrW1IR11tEo
66LjDMXHjG4VRXEupSdjP+e1KmuPO3x1FLdN28kzbeot+snMUT7a94cc832zEVs8
m1JwnhMaPSPz6yvS2XXZW6NkTFxwYoCnMqEXxV7LQMirs4Btr1xyh6VCgC+r9eNX
U1lbDHnFdPULCqu28heQHkdkuPEoDIvbNcHNVLN8k4Iv9hD6yzP2NDHE9Sd2oUDz
xK8hV4FAagqvXw1CDQ50Uo/kYgEAESnMPXFotatvziRHf8hc2JSJtmcJiH6DVZ8a
viaRMf1euGbuAOLZmtU6MAlDxjkf3S5l55Ur5jiuYzxKmgwg00kuU9RqpyuhtEHk
NvdyQopR+gGCY/9OXQEzb5vG+pndi0ReclbLWu5fTu0/QamTmrKFan3yLUghBzGL
n9JBNbA+RXCu7oL046yZq0aEhVoS+fvDbtfBgVik0EJvPZFrjbh5d/yvYOuZBA2o
rRidm5nGJLuTUCMIi0PIY7djLWYg5Cd7USTFcpfqR3e6vbWXDLdjo8cNT55zvs3E
JBe4cNmsvaligS0k5woSV37kOAnO/+6sGX8wZTUUV4gFwanPLxLqo0CWt6S/NFsz
omAtmevTEl/NlCQ7qIadf5N8TAFaPdQAzNY+M0dsAkY+ZDcUI4oSbYwqWlPb4I0a
x/ZZFSOFUjZ0Me1CXXCLq4BS/SYkcPWegHRPewoJxJf3VN1HZkeSDh17CIeM4KZU
qwWdZh7gGBBJ9uQ8+JdtCwI69mxc/r18d5qDBHH2wnR4ar3rmAJSx8V0+OkXJG+P
X/WbgNS/P8NAXnL4NvfeERwGdzb752OVnNvbFxQSxXjBxIkIH6beEJH+oZ0B4S2q
H5rOXC1sZBuSLKloLidXuk/mJdyCL5L9Ggk9p8BXCj00oXohNk3ctgnnz0LTb3sF
9i537pRY/46Vid0VUqw6VzNYkdedF7rESuk9emaZfTxzLJzawRqHeAuDT026rX8d
UZFekkLJz1PE0cDWUWKadb4cFkwth0RmNMrbcoEvOFBfPMCAC3uN2lRVqSIUdAGl
/GsU0FLpN2IjOTgMalPKvu/dGOvAPD0xjdw1zbE4lstUszsJKHoGoV4RSPwjkST6
g7VWZx2n7VDpi9ozske82PIoLLS3TejSRoSbbAZmr92SRR1Ed2oJI0odEjqeiTM3
IwqGda1P7xai5c5cc3BYZQU7PPfzU+iR8KSjSjKBZjSoPbFg9dghZbtKP10y8rJv
wIaKQeWUF2O8bvLb58B69hRpsB9vLAE4B1YHogNDLV3QwiD1MW/wR+q9qJGimtWd
9Ls69vWV2bzfJqk+TiTBFHtKNYb/jAmW1+/cvQ57Fg+ed4pnqKKnqB/2lJQMXDLw
SHf2jdv716bWgpPBilD00Rd2kC8Qk8R7DYQ82pp3zj2iU+EQ5UJUUbv8MlcZIlvN
tgV1IRKGbyBwwFEl4XwhMh1d1oqIkxtLeFyafO9QnqwrmowV1UFHgaj7tDVbE4Si
NQqAywWacmkC3/upmklVKQcA4JGm/DAMNybg4qV31H0nYluGHMPeKDMYOau3jh0s
F5BKgfkpzt0QpiXF7on682n4rLY9YpBKCuH8XO6aJXHPrhivjuF3yJxOrmK+UhW0
kXVcpKdQYuPkWkS3fGBke4WV1bjKIbiZVFYD/0MCQBv8npfnIYdlVZ6RrFpAq3q6
iRay0tcXpwmOIEmwNne90yHP66YBNTNINtFj6oLaJduzIex1RkRo0ZHnWnxkmlJU
HS3byjO7mREad/c00c69pskdxjsNSYThncg62+PT5AunGzBXuOVyKtEnL42EPKIu
uB/xsKgqShimtD0HSbwEhA//oayVAjvaCtPJaL0qCjBMn0FQjRSPYuWbJkaWjj0m
VhKUYMNU7F1wkofwTyXpFdTwrkhr3vsMpvZxTm2ppcPi5XlxCoyRURrSSrcf0EmN
Yveq4VtjkI8zkCcwnNsBotOh4j/oUsXJ9xSaMk3pyOF4rCYxb0Oi6CFOjJjcY2sn
WRpk7hmjtIqiY8lc1/52RzFyDjdjV4W43+T8zTymUy11Sr0Wb+8+NA01ZBaqWH9y
wPvfoqqSXSfd1hurgGK0dMZcIU489AmaWNfpc0efXsVHQG2emvR3RTK8zmz4xpm6
4xPdUQFGMuvCOLN3kDFwcG/p9YzrKP6PY2GCYUv09mYEgFTRwX8d6W2A+Y+zad1/
cOjEhu9/85rWlmOonC9nNxpKRNgJvQb7B/rnfu/1XI3Mdk4YN1tc9us4DQuX7O9y
TP2wCKH6XPIWEZWqPdqPUu0RljrPp8nVMwSW3BGCc22C8Cpj8r4Am6mqYqIkZDYO
8fLqJ1rS7up7WwRFENt/fkKMZ/t0UWzdEJ6wgvW1J/Dzm6qfntmQZNwoaZIyFmWG
P3t/opRZr/zFAYY3szWlNExkxHEfQbmjYnQ7GzKJLyWqM/IJbnK6VXf8Cz9fGCpz
t4wy53meQ45DbeeI7O7QGvYb3qCWr8XAwkivDAWHDyEDEYmc+M0C9NHAN4OIe/0n
uPNTFrEmI+U5p8pJ5zkVpiQ3hkQVUj7u6N4IF3Djz+7gyh1ASDy9HNi7Z0eIhgvd
WfC33FiB2/1mXYiag2oi0UWUs77w8FN6vWfzu5iTOH7w0RolMxS/LpNbtX8cYJ4b
vlySlGs1Dlf2Eb85OUia4+dQfyTve2Upkrf2XyyFdFVv1KgDwkdFZPycmbNsvnBp
FKAQ/Sz5kcZbJVuNnwC2kNTcXFgSqQSFnf4x/Dqm7ONBQVWSwprDKdQmJx65Lisv
a3b+gu6cCTIi+Z4nXcQoxwSV+45KigpZ2hjm5EcAxa1S7yAynauzr/IiexSA6xoS
3Gc9BjQSB0jQKOMHhoqIFhpWjQmfa8zxe0OlUeOn+bpiGj3DeERlL0EchvpjeFXB
itWJCd2/vNMHrBaGkFLNIfNFCsD5OQ0d9EfFcsbfrg1P2tTL6vFC6yGP8kFIUxj1
9s2hhxdNjll7blKTbovpofRxoOu5FEC4QCfsYpu5jAKtKvs8lkW0V6zQiMl83xTm
jSXR7l46WkvyiAnfd+7RBvjBNBwGEwOr/i8zxWLF306CgXpyXfAY4IZ3fEBQt8ol
M5L4Lk2Mi8VBE7vLlgG22ODFpRZXiSIqhV22x/VMTf7x3JDm3dry60h7j65bS4Rq
hemZ9UAXab1esWQb8uNnY0Pz0AZWNB5a2tAYC5Y0Rma7VYWTX8pSqQwOGLanwu/R
fp6AO4yC2XdPt2OOa4AyoOtnpIV1A1UAuGgqFqLC6VGnSHA2VCQ+6/TC24N8oqSH
ptuslKFG8MZ8tEq1DrNGRvLOL6TD0JjjVPcgZTbwUguyOA5dnPqkdHAQKggmwROg
XQj1ObhJgSfXYbSEoq5MLANsxXdVLTIQi+MAnPITWlHr8i9oByrW16sfPkgvnWmm
VLjyzmGzW0l+7QePbvSYvOHZSVyTjFSGCpFn/yTrnz+bQqIlc8RSJDOJrVB4Gbgb
YeMWeU9npWcQR1Xw+cbv+WmomuISXf0CmbFKDvkklW2d6/uZgg41hnfmc0MFd0/u
Sl9Uvx7tWnosQ6OxIgLr48umhWwMXbdDzSOHF/Qr8mgqpe7Dy3pd45Mvc64DdpXD
GkYlpeEFhZHsP6XjWOI6wDwhjyrNeEanZznfDsr4KDYVbw3ZW2mBHJ1iWTNzW7Bl
aGLvXtg355AqUqTod+MjWi65p/bvuut3nxhzh2Hr214UiiS49LCZDTlBBe6dMTHG
ionZ1In6mrOS6N16OHtq2aNQATw2pDUFx0+gZjwIzUpjNipCN2EdY+OEAmEhfWua
bHANItoIlp4Nz1g+FU39J44zWV5gcxZel7XsgcHgRBG5aUNURhhtMa7poPz1P5FC
VQednh1qEQgnir3X3fVDojNTXrtA56/rg26QDnoIjzGecf9dtEeM3bZuWcVbdvhw
WwvStyZ2iI46PJCk5PS8P3M1GERFjo5u3w51xLTgWhd4zIdQGA/BahmPyaS16svc
t0WC9Ri9cfT+YUEZEu4tLEfrDAxX7zArOkuevftYbNSB5M1OvUEFqtQ/oPvh6nkG
o6Sm6j1kUJEQvdFDZHAJKDskX9Z5NUlqMQPa2G4a166LFUvqXjNqb1bPF/8SqcEM
d0Dg5yMbXUL3gwIalFrrNVH3DjX3sdqGCF7JhNK6qaXDVCRRREMhCzrWgq9oxlu3
yWVmsU1gUhOVIgSt19MNvhPptfmScwBDGKNCz9XTMY1guma4M/1yZYI6AH7caeZD
ejttiJr9MQ6IvgB0/QiPh2i4SGNlZFPniUvEGzOVdcCJJhxiV3QXobUsjWuBL8rg
Xy8r9WWPfcGYCM/KD6z79HsyL4qOeBcLiJZmMHlSObnRaD/gD0ntZl9R1A9waifs
BmrszZTG8N3T/pS9jYSIYrhQO3oHDzG0fJ/zzd+vDFC0Byymh8ZcuzU8N1jHbjhl
IkE8MHiVn/pcn/66oskesIc4KLoE8FiMNguc69LobFpQZ02LEpNIkcOa8UIl4n9c
ppIjFdb5zUTNrYQfeNna5gty6Yqd/OQZduBdLibx6uwC7/BY6H5Mkzh/L4faDnrR
poe3CNjrSD5ixCG+R9FmJUcaTV/Yujtd8tr9a7F92MG2dyYx/JWoK5qLnVOrsmEj
1U6bX1FZCAklzrxOhjtfi9ZUiM8YHFAAbtB3ptrehB37VSWCeuP3nMBN2t2ywANn
Ojb6Wylwggk8WU18ke8AxWkJdQxJrz7ksYv6zwpC8XXRZGyY6mweIQRIyu2ssTNK
A2lOrsaQZXckR+jHvtnJhGO46gatXxfHM3duVTE7RRuAWhpjLhVgTR5O/Zn9PBzf
D15/JZttIsvrCR9HMTOvtmV8DcgC1raP1IR24xROVBqeuAkuC4Eo1MxEs5vVaW36
hT+t64g1V6GQVW0LDN8iouHGwQaXcLKT2vydYbKZXZU4iQkjDgH4LMK/XOWkutK8
zwA3ypmwzO7d4DTpDeZ0rSxUjPY/guwlFHiDx1rsiACEYysAcCkF3c5GFcwB7Eyd
LSyWQnLbSASC088Q0//Nmmsemw1/bwD3V+CvuRRWutHFWv+sTywFj5Lf1UV2HTHA
WP6oks37Cmm8spnrDGw5aF+ETmZ/6qKofLBa1PujYT2ai5fHUkbgIS+YraSTJlka
jVv2rhmtb87emWenThLIpUO3FV28Vmd3hnKhOzaHBGFCDCAEjKeyhw4ad+fosHaD
j5U5Ni1d8MQlwj4IiPcbo6ZwWmLpr3f4KQpk/Xc6EB9qtvQu1VMAgOWliB8BDhDP
Rjx5wysJ8paiHwUOp+VzW2Kk9AglSDnnZ0jUQQA+vAck4hw9D+r8TDdOJSyqXxXB
WfO8SAtgyTuCAacd+b0mxrI+XudGcNsD+jxkGlD08qlNZuXEeD75mTNRHJ/muPs5
kp8hx7aIz43CdywCi4gkvp9K9Kxrl1BnuU4b+CoOpZUguGEZpUb1xtltq4A+hsmC
ilXmOuqXsv+chaEJDBiF+AbFhXYroOlHeVT3TI79dz19M/wtJhu9sWQjIY1X+96u
CO4NDsJRbesJdfsffA4xgsW54rzMXSKkHmlamK9tGselmitQ34L7QVShiwSwrvXm
Yb8Zqz8mGkFkrWT4INCGVutY3y80Kz4nn239aToK9HejrLKYXFywl5sPGfrV/l0v
JRuEO+uGNmEMsNlCjA1nEmtm8wJI4ZQS49dCen2Cej5/aESDteLvad4a/o45Nsqq
jjZpKv4XTYuyKLWFO+k1EoCOhlTv1hFwZ+zVCdsEcMP+QpQvoWlqbNu7XW32RNwZ
vwwsFRxTesJT6HZP1boy09/oGtQ5/YUiwvJNWri3qFihmbodW06TId1CSbwqAD26
wL7ZC7mGNIaCWiz4A7GDK1yCX/eYhbKsGrdgRAmp8tZJw+9+atn35NNfci7/xFAm
HUmzjCf5LwW8fx/tH6SrzVW+GPgTJ2/6m8BcOeF0NdE58BovkKDDQgqjEf9MHukf
lXAwfwMKbGxjegMZJXKhzqfCrGUmmXlPBK5BtdiwE4SswJnmHAC5U/fJEZi/NVtW
CQ4SRHPtp3oBc0rXclckAckT5vnaI5lNtMRXK28zwF2QPZcv6XpYDx3AqSLwjfuP
izzr4pyZPbFi5VBZpy5zBGwlPdIrbIqNYI6NnGb+zBNrpYxPbhLUjwpmNvDR9p/F
CSxs+DBnFZzhs07XrSrJkyHz6ahOasU6Vlk1hkZPGa+1e/P5IP+mT0o3v3huT2xn
Yw5+nwyS01flqIQdyB2g51zu6kB5RRWm9ZwtPVgzS+cZpQ221so5h3NOOCPLCfrQ
w8rFUPI0Uc3xzdNlo0cIJV16zdBktp/oRTJ2FZQIeQsGOK0nq/QbVih7f4v+tlvT
olMGGbFSh6JS71fuwEZGxpGeuthpqf1+weAw+efoJE24BFnLO22aIP8IqQNoFaCn
XEZs6eE/STsFr1p4wYwf8m8dcGmnvHtRdhKiQv3XiE2P1YzGG/0nq06XCYYm6Yy4
obGgp/vjlwgXZ9NEgW//DiPDvW6cU6ckWC/eac3BoVFLtZYC23Bfjg76oGXXA3qa
duvXrIzteX0gXyblbUq9Eh5Nz87Ol5iBIJoIqrtXOoI68JaTeci0DWP88faTwGDN
mCkkaBziH37sajQMeqleecCtNADNvPcNV2tyBuhIp+kd6VwAu92YS3wZDgkw3R+9
McgNUpb8tBl+Q+AX8VGtgUJFqWlCtVp/e200Fu1WMb+gD+SyrPlyEcujYVpIsDLJ
6p/JW+E49dIbrKbySWDCSo7GV5k0vni33eNGjSfZFO4Y86/+Tmx72e4esWIt0PyW
fDAD91Ks3uMvN3zQ2pI+NhlkXiljPFOs4keI9OMUKJZAV/6GVJiA7aqm2gCV3Tqq
OhJFakLuUObolsCsJx1lW6mCAAtoYl4YICZO7e9e+9LLXTVjiwNvf3r4eoQiCG2p
vjAX4nDWXsjj3m6s0+S/MSMesUNCs22g/qRW26pxvJlGs3Y3PDXJtnnf1+xlOjQA
QxuoyO3Uo4wp1/cKV1St4aKBLcmrUykx5vsQjhybZ0vTdiXH1/HnFwcSDjAUS2fy
yXtrvh3pVnPUIeW6nXrGoFCHchpecZCnUaZ2D76dew0NaeYuw92wPReiDeCvbYOk
t8fMa8yWcMU+AUe51gDQZfdViFRg3jn0Qfus7sY6ATo7ZbjkcgJI7T9qhou5aEzW
/HPor+8nGzf1d1nVs3uAPKPJ31j0wAjEWxFXBZadXDHdNADEJRLbToDIcknX/elq
cPEUoXmRu8EGaNeMIqJoIoND28vSgnaXFy5l0jG7R7nv4goGyYrRgavY3TON6eeG
VtqjlDdjT1O2uq0C6oBElFlAOaBpbEuQnKIBs15Fy8MAUkUVbGR0a/f0en14ecG2
GHvliSsUJCwVUjcHyX4sswYp1iCLemiuY+MQ/O5dLoe59HFMnIGUcfMnOrRATBV/
6+fuRxeh3EM5fj09yu20/8+1TQ2TYtWh6pR9NEwAKS14qKkY0exY9tnGPyw+ZAcQ
xybuFOaXD+tbf/YwBbpdrfMD3QNJzzCwRGbEkLXcAgtHCjRBvA2S9niYtIsIFipB
O6/7WPEZ5FOuBJ5trmvUfkybnQM+p1ca2kOAP66Gttoxh/twuhCSR/DZL4Dp3EEK
EhCwqs/25ExF6UyrNHwQzqpomRXkUMoynu4d0Fmf0UYW/8N2zrJwMPoRzM1GV1kC
q24v2uFZ+hFgCt8LPsCq5r4/EPm9hRpfSMvYlUeTinoKBLw7gnHjTPNwfIwwUVA5
3/Fh81Kh5VDLZ8wCRKabN3m0KxYG3ma/K7NkBbiAnckLXwLwHt8ZtrHPJCi4pz5Z
SQEKUvUhzcSyeox90PXilz9jBMBPDrCfj+EoRTgmMWF2cxpk2+5LOOAz1ixpJog9
A+cHSUuWAkP6g0vTuRF8OH8yY0XUfVYKDKvymV7VlKDb4sZ3/ShM2D0vYgIZ4ehH
ycMVgLqzgxd+8nDaOmmyHv2Pqs6jy39/ATG/u7t4e96mAeoAvbCuLEuvegocawQ1
TTflR7Zx6fpcAhq3vngTciv+J7GJXrAPROcgJoE3JHZKHPtAYyjW3EX6+RnpmaAs
zwz9eL0Ltcpw0yW8Yl0m9jN9cYVTrbjCDfOUht1Vf/6UKW+Rd31fMLp7RKZaqlAy
5e3/kczDYiM5SBLSbNjVHl8Ne92fa3vGB6mWJVJsPOoIdP+UGil9n0Ko4rIx4wtL
77zH4FeZ5lAE7qIMFPrCNUVlrKOezHUwoVeU+F9Rql4Xe5tAf4pYh81Pp1WVOXdS
Gb4G8PhwrVjVFmV35XTXHWFJGcKVc89Aw8EFxZV3nxgbAuqrSImBZ/dJT3Rjx8Zd
NrImuKfdPa/Q/aXSXNcxWD+Jw5FajvuM91egjNdR1T3FBDzlxKleK0pTr6HjtMY/
XCO0wXk1bsiG4mYcRsJrT2PDtNElBq6aUIlw1gdIP1b4AzIltdEsi3oEKMjZyebu
6evXrmm0O1+JFfdc66WyBGJmEk/TC8NmdqXlzBo4q2QHnHJkW37RU5B2ew32M4Pb
fivkF7zlruGcuAgusjXInosl77AGRNfSH16nkIy2sPibsid1kqbHcwQOb8rQ0Cf6
dPte2t9nZS14cBqylZ1+YSrnnWDgrS3wDpCQPJgD8llTRlaOJiDceDgHTf29UFjk
FEbcWiSxN/aruXWZpjuOYOMV58lxH8IhaJqYrEOel/nG1wljx8onY97f2pLo7vRp
QyTDDACKi97w2U17/IwtNJFyl5eXCMVh51NLF5xzyf60CoBLkiwZO2zt0u/a12GV
f3ilSiMLHlr8UMY9lkA1RGU5W7/1GJ+la6/hWJn+/Bz0H0Yy1sO3cBxVCfiQSN2+
Jyu1FtmgNwXIsdlJTl7zL5cBfjgqCh4RKCCL1iGgg76dZgDLhfBj3nbP9DS2FU8F
Vuiv4rpmA4G7q1vgkEOTBG9z1UvjcL9RIB1rFf1xPBvT8KfJAhbFhiTodHlZzTS3
o4nE3UdseO0yapBtnyfzLVpODncQdzpqKnvZqjoj9JVjFQL2FGHLCl/LuAx+mAcv
jzxbyivUlkr5G8vY2T4VKi3YHq9IXu7+VJxzOipQS/1fOw3Zf0tNUiODk5cz2Zoo
pCkAaWBoI8j/0lJUxtpEIfRZeQe1+nUQIzXJDg5/DAKXuGYjKBCi680TvyszG03f
9M0o/9yGNRxuSQ82OYu85gVr72NpWJUZ4+r8X1ghRRYd/glo+8Sn9SavPEXRaLm7
cu5I5fz/UBx0Qde/UtUeaP2JU17935n/vTwTW2Q3JqhO9x1DiyHwYxhZFRrfeRw+
kuHsfAUjTeTXOjstNHz3pX35BB5OVr+oE5icPsLythf1aVM3LnZJjOtzjPVYSfrI
+DNYC1Aq5TqMbyt7boUjiU1p9hn/vPhOklQ+0MnoUma1YJb6uaEBTs7Xd/3L3omB
YBXFVZQ7DTLVQXg8M+pMVUIaQkzEA3Iw9YP97pu2IxkZvYLaXKF7vfv8yUpnj0nu
jqrxOXfGY3K6LmMgE3+F/XZRXDRPe7ktvImkGT5W6V73uxtgBjrk7YnTr9K0S9H0
NtcvnpzcsYy/JfBZPAce6tzL4OZsehX12pzBANsUCS/YzIUEYQTZEZjpMiniwL2A
FvbfJQ45QS1Au7UZ0Kcnv8DyuaVDJppNI0XFziOrhe35tXA7bWHLI+K9Z+yp9eqe
tQA3Dyt2UjpX4ZiSXYs89j0h5OVJSOJWchrZATNGGN8i1QsCZUfAdHjTG9YC9rrT
9qbvUiZfK4MiV2pgstyOZy82iItsa5GJu1tjQolz0nxu7c7WqHxaVLqe9pxu/5fa
1exM0Zg2/lss3+lmxXqF0Nric2WY+pJBtdO5BCx79KUsInvz7L6JuyXbSSTcR8y7
W9z97HX4nzWfcMMXbTJF9Iixrr0O6HoODEwkmIySvy17JENG33q7iqghvDrmkXXY
FN7iHSHfBTmfV3KUAfj24C7O8no6SCYZESumhPybox6WMxeOVpjmznADoXQZ1MO4
e/j9lSulDL/xblqxiQ7yRMpL4iJe7I8uoTC4QvatNEs4/RFlhKv+YSVFbo5DxHky
gr3JFSBrOdOGLWIvKyXhBVAN9oQnwJKrrF8wE775QSWdqUVTzcXuR2sfCa2FOIas
kTD7rdLKDO8jX5dP4ib9IxmetvB8r2t1AOALuaa49Efw5YsnWohs3xyImtmHUbfC
Y/rtmC1KE4XcbLrVhEucAV9J/4lT1eKD7JybytmgcRKTxfpQ/dFMfHqzvVcHi5Tp
wOHF9C417+6ljD4HsQnk84BsvXZXqy+VlKwUymN1AokxVk7AJSP8+yy0NEGNpCuW
togJ4e85M4haj1/rDnBqRdf4UH/WtDak9CpI+9uiR+GUhzN9dxHeKKyOav6MbkBI
wO98HuXQs/kKMvmne95cPPP7zAOLKF2h2PfCs2W/9l5nd/fom1eerK70gSpf2KP9
Vws5zoJDeNJw8FSiYQ+0KEYneFbyqRPvmuk5IZynOBt7J91LWDjbxjFixZqCc/qK
aZ0CjOHX769LRCIzt1DB0UHtvJ4WAZ5yNdqInxw3ZXkKXZyTgF9HcT7Bj1ZCkDZm
j1wAfv53/bli8LdWw5ZYSU821dPxQf+b7WwmBgoWh3rMVlrdaW5nvqwhj4kRm7sT
7rc1+TPsCtThehrIWDYuNrq5bRwiczCGa5qk0IIUpCLm9kGvYD29aiPk4pwBWMmU
ObOIdlwB4cruRzdlIAO+L/anMfwbXS3yP+K5ZIDrqaGk1pEwJsAhmgsexhKj+1ge
poxgOWyaHQp2xTZ5IuwGKWY1Hai4qmJ9Yne40lfPcJ6uMIU+E0N9JHQHNCFAwRZQ
MCJUVIGWOQlaFukyEOuini4YZI3EDMG09wkN72ZJxDS9fSsMOBXJXKI+2AofrP1D
9vMsnwrZ0LucTeTgOl/D7RhP5Jy9hNehTuG4smnjMN2xbAZ1ZmnlfL6kBp8A2g7O
+MMNmrSpmE+VJvTaSd5gST/R8kmXE11Y5G0gOlvz4HMGBgJr0OerNarngX19BTfV
nJWTvtTuDsRKZZrgIyNvF5uh26ViGSNjZ+NoQKmtT8eBJ27OxHRD2/AkhxUYWCV1
Ug0gQsaJdZ8TTC8TnMiHRNeWUXN2ckehcOPyNPopdVp0kwZDdOXX3ixo+pnHvIui
HbYCRbnts1pRqUz+sP5NVz/Uc1Jwb/GmpJoyXY9CTBEHmARlAJUpWSHzpqLKnYQQ
fFwL5AYnYHTzBvfOJwbuU+IDQrtXhT7p9vTpTdgULxN04xBlj4tb6qNEm1KlV4SZ
7dRlWHBWMRlnivVuBL1zcVVCxS78z6xfJO/kmODtp0YYOqRox1hT9V/NA8R6Dci+
kLgHXd6BX82i+WchcVKc9xPqLo6vCuaLfDzDI1A9M3tulR0u8YxDF17G8T+kHDbL
Vyv4YdUzv9XkVIjoAvninYBKgmftjyiFE5lR4iuvJBxBl6nEEbEoyiakv5gmSa3e
bhHz41cnCsX0JApB9Nzp7jgLYSKRgpXspRLHjGwaYShv5zmITDuxzbh0Pa1HI+7h
QmOKqpESh1269kVQCIOxvbliQW3pzD4w8u/nA2hkQRdagFATcuWwhsDWk8+EG46k
2HNuPcqUagmcj9BuoewXC3Xj82hTSIdMoWRh0XIggpAaZIPqG5EUDHfm2Uoxq1an
z0rbIFelz7U6x4yGk3v+blmmU4JPhKNClYqvagNVL85XYwjIy1v5FV5A6TyiXVX2
GI6HOndsE4x74ebjrUobZWN1QSu91PQk8P22jAihG5Zqb0I7ImFw2sNNCEZMvKVj
vfH1Oz1AfMMncmj+TuS0UTY1wUPWaoqdBEsbGf+C4P+63NbTDAjY1JMT0EDsdhqD
O5rKtLQTcbWcyeKdw01am89bG6FNmXYuffBPQzYNBfJsk5voZoeWZVS1e6Q96Ps9
xFAzcfqzFuZDV4L7TsvNGIeYyZ9i5+jjk4hnGDnT5hT8VXfeseHJmxjHLgPrbAi+
bsyJzsOkaj9fhSgiRVoC2SPWGsTWgOlHty4lpgtP7I0T7h9i9hBd/VgCL9Yaebmn
groAuQ22HkUJJjS7aYlfq5rxs03nMiHTZdCRSVDAwHmxbWdKaZgQ100eQ4IFD/XI
486gVQihCTl1plQq2Ca+HWG9zGcPo4Ug6Wy2+8SIK8Tfa4p16KRwWovKNCP+H/sK
rx4BtPnejjvyYRJph2OK4GvI9RnckxG+HgZeNii2g+2PecDEiHeNV7MyU55aK1PA
Zwy2TCA6UDdx4BVK3PRuDfOEXjXyU7aJugCFuMYqs6Pd/jIsOamLlcq3V+SFsz1+
XPTApK/Lcgc9sJTztHQ9ughZ7KkzhSz7ZZh4uMlg647lRfu1/MQviHezepO7TmdU
1Hu7x/AmGgH9RT0L6+xBioPdcTi5mGGuZXDboOgXJKMAc2B9XT/+yFgjGxLzREoh
abOnaI/x2x3b6LxTssMw2fxO00qWqC78WgsrnWKaDiCtl7dqmHgmP3vlboSdLl3I
CNgKu9SwW3tSFZ2cj9yXz6EP5hXk53DkRaEwFBs0JQOwRoarUVOYLAaneRg/65FA
8eLKdHd45vzGfUh9mfshYp99DqKccRRyJunqPxItWXQxSKxU2wz6Ajr/abVF8B0q
oBd569trwig/oVDqx4vZkI/td2mOgb2CufXPTi77IYlcz8tr9QXhZ3fC8396jDBe
PAOq2oKmxf00ItyVbGWS3G1klb2gUORckj59x5u9Qa2MQP9oE6MJiQXeile1f5l7
j+VAZdY2xTUwvRXCvY7W6tknObNCJjIhXUxwYAkKN/U8QQYgBKYy5p3oIFdsQBns
sy4ujW/txZbO+r5aMzK3BRWXqlembLW7CJkT79UUmKjyYmpNzWCdHUDaUBfeqNJl
hKqj5tAby5rM2Qr7WAlKh4vErnkh95tmHNDxkm3iNDz+MCOtYxeXD39hVq4mSooQ
oHFaumhyEzUB36dZe07VaK1Neg2wtiAVdSdbotDUFnIvRkLrYjFusY9/DJUsBFgY
tO3tXNGkzdmpQelTvDhYEYel0THVjhc5PyNPihqUGIftH6o0ewiEi5KHJzL+iny6
gbTjLN5PRcCGguPGzYgS8kkxny6FmfI1UA5OqeFczR0Vic/oKLKEbCFzQU0XjDwr
XVDBCk+4yiQRUWgI29E2Mdx+iM+yH5d5Kr+7euxxhhiXdxBXVHzEHTm6YskLs+9r
ug1Ey2nbKm0fhZspvfbXTL6afY6wz+g+/pngpj6cDKrosswPA3HRS6b1b/3mabGR
GlzUYjEBuJnzT7eUj5jrtSLADKRDDTtjDGaQ68HrluT9NJi+t7akvJd7ek8CdlZu
D33aw31Gz+PT+nrST3Ql6ubsDVHC1ul43+dtKTZen96Kb6mfLlMmsO86iG5o09Pu
FfkHgkZbnuXWPNGAyvKg06FWE6WAzgQQPvzTh2dgI5yZgJlmy6hxN/96A+bwikQr
OstVIoBQIlF8LVoDipTiKyLgaZIcZc7Nuyyq4pCU6rn+mWkmYtmb24s6lpiHWyy3
RCxd7mYfq62O6OgsGXsxudL3dhpzCrlFDE5JE/KrrL9uy7n3QW2dfN0z/zGn+dXk
M1eCJ0VtFbR1koc5s+x2YW7BIUKQQvfe01rK8z4ogGODarXXvpP03uqzHDDn6oKu
cIxE3j896q3X/zN2HyMIcgpqArtMK3RQpaM+hTJYnuem0058F7RYUTQk3/Jdyd58
QdVy0tYLcLo5p3CKkXou0wXbpyZ8SOZ9dKvMZ6DZOF4olyveAUbOtENqmq5JRJA+
zb6SydMgBJnW7hgNgZv0+n6QndhqUEk7/x9zOPUrzSB7/CMF8yukt8guZCDmi21f
zKI3GzTcHzT9d2khaJRSkAGIpBEiqv7TkQlN5BGFHIj6+r8oV/UUZ88Bt/5X0WAf
aILdhjDaHz8gFYFawpsKR0wAQY7cijGXWvDW7d50xKz9+ze2UrZxFZ/6C6FM7AZ5
AbOw4VUyYuVLsDMo/aymYV1HSitPvUyygjyu2ew78z9O3ngN56mKYsrtU4xh1LhC
8pb+YZtkcxMEsRHQv5tGAcdTU/5iIKAUyyMKtKXXAr3qeBs3AQTEFzHjG11U7Cwo
XfrZIrfPIjlZAW8i14HW0hvODed9AJ/rVwbt5qGk1Wf8jLM2U9ak/kBC+VWmPXmX
A3WB6dFcUjZ6CMRVX/xaS9A5zUh086VomAz/PpjP4XS+vqcf8ShnUKPbkoDyvxna
UxIbYuF77kGeQP0o/ZLnoZQ5kmrqw2Wo09Q8XCgByyNOkOuYnDFVX7w1fWiQHMeu
ajYq0D9a/p2N5y44H4PzKh5PLJPor0lWOlDegZM/EUPFHGO3jVQ/hBYHcWwJJOuq
vFz6Yfn4qE+MonBDVI44MhQlFh/YegTPVlofu7Fmt9l2SJQ218QFn5xUj7WET3Dj
HA+d42vRoh+3IEaU2W2URq5/C8IaoIwWt8WKX+xPikEAEosfwBMpj6ZUXaMfH4eA
AHyi6JKYdo22hG558ZFVNIJR5skx97S8LRnszEcBuIBP9c6QqJpN99yyZ3ceL1uj
BGzUs7Xdce/q445XVLQWO/as74dLyE7PVXw5WnDuxtNCsfLVE2+B6WuijIbjQVBe
B8hGzmjiRptFCMSQXc43x4Fowhs5QXLXzv38vCWyMa4z/aguDbOrb7GHi729Efr1
N9Dy8cZu6hqyAKGEHPnrwdalFmGwUz+x3AYYy8uInwil/2Slb/hOBQZNJYYrQq2X
RPKsO5iBfNEL7BSUusJEJHgRmzpcGrHrBwoWe3+YKYKXGmgJlBs6GU7nKkfB7HsC
9Dr/afGNB/l62mzjBLkCd/kik4btSGbd024vwWfh2DDaG0MOBEB1e4rkTB7UKdrw
JajSKCciHDIJKKjYjp9TzVyQQ3ySakourdvft5e5TxU0VqxXVye1ZlJniPc17pjI
ewxWzF0HTUwIxp3krVtvl47pHWLLZu2qojErG9Vg+Hk1W7G4UIi7KiPf6LnAtYhl
DtzQ4I4maCsSK92T7/6cFiFXZdIDbEyQhiOgA7Ca3SWc05dU4kyAvXu3N3WrpcBt
0Ca2cW+8Lu/Vp7d6EpU5AhTn1UIJqw+6TjpaMvQpuJECIdcsulQtVk4d26bxhGYh
JJCx7tKSCAmMLIE55ID2MMBqmXbkL9uPi7Himtvc6ZSbu/WzkHO9eAtta9g3jNFO
mi6qd96hPXB+xMooBUND1lvR89s7agCwjUu5vjzrXApDzGK3t6BtXykBUuEW3uiV
+afZ5Q3J4HnkNEm/0yRlSwv59FJIPb1FVnNZ8wSzRAzM+auUb8zZJZ6/E+RNbjKz
U+2lzNUMtpvfylG8AZbmyYacC9upDJtn184R1m3dKROctpCRd9ybX7Rhcilb+nkr
coVankCil0jOb+73lvNxi/i+42JOhwBaAiQVdJFtYFySJNmQ3/Oow5exN47iLKn2
nvYzMTTopXWPnZLiQU1wQ34pqusCFNCyEDQZ0utPgnLicHX/BW2imAWHH7RFMilI
OihRWzhqHnpG3e7i4HoBVsygS7uI/adAk+BMSRMY5aipH+CD9E51tDPnF4ZqEuQ4
c8zocy+W8/6f6LaxkH51Ot0hmdg2zlI82BTzwnzzte9RZG13YMlglBwxw+RRfF1B
czKSywrxOttiGng2r11Ef0J1QVhGmLXRN4TJOPgOjw9nfT/tsQ3aQSZiebEGqMsC
y1axKWxSEYj/ao7CYvUMERLpvxWvk+4BbrnrE+/8bXRs4TzJRYv+hasOUrK58nUV
x4gSGBnQWmX/MBjGcHLybP0fjaDPcmjtNmTLLbGZXLlKLDmehajwsW5piOLqs5Qn
ssa8SVnJvR6x3M7CwY6dBmoBnFLIYL/oAdXQ0rLOAzJswF8pB3Ih+5s9wrAse6WB
00N044EAaLZ88ZV5BOwK8cxsL3ea+pt9JKmUzvSm6SUbRe0ugyzlSeQAyLOpo02i
LveM4taXBnLpMhGCpJiiU2vE+4KLQTkSm1Cqbj+rzD3JPscUCm92F9WxmD7xjWcl
xK9xHUcgOZMaSq3EqEyN6Up3pqJqcchbx8kfOGZ6y+9MbMldsN3fIso7v8pza2cc
8WenXLvwe2sO6+AZt7GsNC31u/+IERb7scJjlz9LrUnrYA/ZqclTMRUyS/ShGTp3
LtROrYkwimAWdDfoESAqb9jnhfeyw6G1GgdcuPe7rmavQ9Py69bEz2qDtTGb98RP
uwpqEn9cHd71l4ttBTc1/S7oWOdwCsTJhlEGeQH+cpHwDGnCn+GSOv+thLPO/TPu
XRK6peNCqKeKeVxf7wMClju6Ck6YNMygl+8vtDrpqw14veeu0p0fHpC3ePu6cPPU
kg42Qb8p0a9JYojJjHW8DwzVTrk778HUY8hm4IvS7yALiNqv+jjMOHpp2TrcuehB
Eg9PTAMs1mhY6U6ZF3jY0UUFSU6Q+Tu1AetGW6O0Ge1BSQsWePNmC+3C3eUH0xu9
XTsbXLj+W/B5v187bn+o81vnakIMRBbAiUNQ1GMr4iuw67f9Bw39aWJ7/BLPFHIE
0AnCgz4MV/9FSVwYRzb5sXtny1fRoQuC0EqK3myAbOEC+8kJj471YTKVasfif5i9
qZPuCSZgwqtf5m+/+OcwbYcNRC2VKOIDrl4Hg+nub7k3S2n0uSuuDZHmoJRG767N
zAqz9DDFGQEJSwU3z9019++5wSPVSkQnXA6Hisrk9UlcQL/DuUcO0hUNqDrCsHBw
LhHT5pDnJoIOSAvamjMJT5Js/8Wy70eE1sPZhE7jEY/HcHTRLYVTlMzl16tfRCeK
KBVIr74aLx16cve59KH7kD49gCmpJSV9xNALEBERm+Q6BCsSji3AhySSN6EuieyV
WtOhxSkBJT1YTB94ghfTMjTMnabrRXJTsiXuV9AqicsuFr3Iv6Nnos3nuDp+ul3z
auj8ioXU7nwfMDj0NYFf8Iahau9ZRmk80mUfsDfVNqUDuD/P4RaHwGYwVZCjlShA
4H1QC3N0JBnAPlhAzgssZRFOi6EppgFLhuYLoTsfcxdSY5StfCdZxy6YAiRaZzBC
M50e32WdZMOgNO/cIazz2Si2sY0FZfhIuiRawZ/pmF3Mu8Mu007E2Qgh6om5PDz4
jDUn4+rKdOXlPxw5ShQyQGXM0BIFRu1X6AxAGDfHYH7eZuhLOAqtSCFJ0Ed5ak4x
cJOD3gafCzqqFpBe6ZzSqCdPSFx5zBo89ZN2ZdriPK37N/VK7YBH44H7vzMA8lME
AUEgekMU8c/8W4DlDwnmaSnMOnGJKXGLJpIBaKpDyGk2mkRpz+7Z9Y1DkX7UkXlK
JY7jG1TX6DnejmO8Ehs7DxYZlB2S1csNGsqndzJLYWJMiOb826zO4iHKNszmBcwl
IFrcvPnopu2vkP6dwqeTh4ONTMUF38WegzAPqzi7ZFzf32bqrt/kqGf6HTXTQYf+
UEnprZ3pIq9zYyd+FyXcqT6aM8brA3YsvJJBHIbnF2KmEz7KgKhqGU5JzFisM2eT
HjeUhr/Vi0b4qLDeg6CkJN6Jk47Gpk8QVO5rlfdyC+qOwUZfISctVvJ0iJ7O81Ph
jJUkGLNYPu921rVR9gqLTzh6roBbs6PD1OVt+eqsQTwVFBdvqe6ihV13Xf4NUH0h
bzJr9W9BLAA/mQ+E4adXvBPI6vQc3DNUjAbA1WNKHsiQGB4Bvyd4wyzzCIPdvmGl
6LfGHlW27owDd0GzBAdWlr6AGoGihMcHC96OAz3Mu1qdiyrbn9Qfy2kAcS/s8rvl
kZInQ6rWbvZbvHNpqsekRaOSluoAN9Zs/k/jl47mhuAlhhGyx8HL4X/Yl/w6MabC
Fxbpok1lTB+dPI55QkpKasmDdJcn145+V8R3UQGdNaIMsJT8nDp7khs+H8vA7n5I
psJKq1U+aYZl3PLGrZ6beDnswB/lL7vMb5qd8oadoDykFHBBnp9AXcnxipY0dDqX
zLapKQX8cSg/e7h+/z3vcDv7WGpGVYharI7Q9wwxIKxhcymMAtZ8dOoLSXRAyjrv
ThOUUwRE7sAzEa9yCnjCnynjOKPhqTMZCZzf9H1gKr/eSaZTzcvCPvx95q9Kq5ne
/m06TQ6KhuCue7jrNYgfJTqelLavxhl8IEnMdGBLYnAqK44w8Bq4/HiCU1+2FDM7
qSytbJa+EnwilQppUAgc8LAG6D/d4kLWAMR5MhwQuZeTcQEZUL5JsEV8pjazHApc
oItc4BqWMbel3T1H/ujL21A2qHhwbngM+tm1hIp+VwwLdH4ZOlOnMPLoHEiOgKIf
5C8kK4Qe21TEgbcwhOwRqJBl9D3kyHZj01ZdcdnI+ip4b/kmMooWvdiHkM1cskSq
ZM+deQ691uzOANnAoJAmy2sY6B8+Sk0wlqxJ4Rvy8ZynVW1BXdVDyYT8HFNmOBLz
Lcxe0C77WsXDWY1NuUMkeoM/t7En1u5uijj9C6jIGUwk1fbp3+l9LmyiXfCo6+ug
V6JLVUwQJ63jQ41JH1YOrURwEoWflRunqf1r/5POp9NrfDpOYPpjYa9N237sEW+W
ToVDjPj64jpZcUFAn/4C81E0snzzJnV4CcJPnwH/gyrL7RSVeGD/ltP549hw0fDm
WZ8yvdmLviGjMtREC2hZDwqm+xz7MHaT9jjw4pXbufBTOF3L3CkXwDaR4xar3Fzx
fZ5ysuABa0IPskgnKyGEFPDUKTWW5pVRGa8rpzXCze+MRQ+TVZJDbXMG4mj+G++X
1fBWMTW+WM4p1QbSeKS9TG2sGT0hqmjIWTwlMLm64uuxZd5TZfFpxEPGIHj6s3up
uuB1susZt13NWBw3cvyemtJpXg/bK93EeqrFrnRQCR55D4lJpeRmZiEk81FNKpN4
FF3MPyEbNeaar41Rj5EELF2sDylb74WLy4ZUcY9PPFOyR8OHWwUIpYyqzDIXYFt2
MJa3gXypcYO6d/pkRL9h/wehYrS7W4rCRqkbcqLiQekeOa9f2HlIhhfixi6QhpPQ
o8K56vwNRTo3XsdnR35Wndks+6/TtdEy3HI66Agyg1yz9TVBjWAVHO6R7BTBmPMc
kjBGRW8Tf5vRe3ROcYQVtELaq1c9aMJ9KjsE459Dgt5pJUzIlcQYC9dnd3udeoAn
XJyw2rNWWs8ZPFLyMNaF/L0M1y22220S/1VX6wE1gvFZVoAKMV2uk1l45vO4Zs1l
2A0urrFa14fcRDpCdsH28KVlMKcm+xI8HhroNYRUuBo+mHeZqHO58wke6BiKWF9B
ZuoxOLxYQ0xsbepN6kTDi0YnqQl8tXZrLnuPS8F/DDAvZyaVxcg6Vs0TEmEnZ35Y
k44kyYRUqcv01sh9yKA1My1TWJ2bBXSiGCXmWLtn42bVBNYqB8nM90KEIPxVwVtx
UT8Mkp3gNyVAmruf40604dtS8dzLzJP+e5dJ91U+eMKsiuC6t2ZCRCmvbJUflByD
PKGCdr58JbniRwuuVaHo1w1ukHsttT//mhbb8lVxR84OetdjFOmA2yyg1yeumlWL
rlaZ50fvafXS5cn1JeLdVgez+fnRq+f7oUrc84qZs2+UdhE+nA07fXn2T0AFdudD
wru55mKwawONTy3UUraKklv65N0Og/KwMllC4UOLoT5Ay0VzkQbU/ngn8GN4Sg50
07THB1fO8XkZoKj0WZMfcs527alIv7GXB2EVkwnGZDlqCSnZ7wU7uBcfaSOjyuY+
6oKfprGgUwv+8c9CwKXiYN9TWFA1q+a8VZ8oU7CfQe1wyDFi4GySUecgQLmne4fy
Kim1d34K4n4wL7cLI41hZ/Oyg4cKu2R8O8/eC76r0fRrWs9yXQDZvJPuSAHGxQRp
XqbZcRvs8GbuQeKLIvvxWLiGRudB7Nt/tcMpx0U1qUNB+8QTDEuvyjPxrNjXZrpP
KarlBPEkxGmsb5LZnHXENpsTIV2fBzdLBZRnapgtWasUFDlnkbLU0M6T/S8RbbVp
HCe4s9qbafA4pJ9L3Jz/2smTzT/1bgjWxOPjihbbGEc09hCIYU23f26kuNMLjoFF
X7Vex3afhX2ZrMs+6W+fxOJS4ZfUs001Xj7YMqAKSaPZc2wgDQ6tPEatxWEkjTDz
QEoqRL87RfR7BrpPMTaGj75FWeDHgYLWaZ8xLtRU5ZIbvWUVsrqu8Jf3A8c9U5ij
Nyj97scoT74z4hKN9CIQd5iiqLUmA5myB80Zai+xI36i/RUzumpxKkfMtHkf64+j
er8RBLxCEME+JeJdqEfrV4R2UUJjMh5jRAQcFbD1YIO51cV36f/hfHCCdjgVeLQW
ucfRUGETlbc008KhrnbR24oss4dw2N6eBKzxE4b8JtcmQCH5Ib9i2w6BKIV3WzWr
Z+LYB+K1+p+BU11cwy186RDcbUwctp0QpMczLshZ0EGiKDfkSblJe++D04//A0mN
Q4ENOooDAVeG5ZmdzmoKutQHc/IcV/aCRB8sDi/IKiLRmI6vIa0n7ntgGs0P71jG
KAzYmt6kPsK2bG8xXiuvfpk998AW7Zfv1dmPg/M7MQkNgLVfEnKTQnFJ+EfG+OHE
3lVpkagLXUM+Fi6+ssTD3xpX4JfUarTpX35MuwID1xEihsQ5j0V+affrKp9H6d7U
cwQWs7IY6iAV6sgtSMjzOEGwEOmT8MK5BK8EJY+1wgTt4R4zczBbpk3d2Pm14M0z
LsZ+W3+YmhPmg1ZkL1hpgKFduAd2IgvggxLyI3TkocR8i47wapaqNhITTBtr//mJ
Mm5+pe+RgKsyCBtXBazJC06uGmLzlnDt23YkDvn1joQx/FLBBzHzT/axs5Xc0Kxu
Un+bU8wxaeZSXIktwOBgHenluoq626B1pC4Wr+c7QgXixtOae9katE0RJgFNot8A
XiTeWXiURyXSBiqQST1zpwRrJfAVvmz4JfeizvfzP1Xu5fQ92fnwboeFcmic7wMd
kmOsP3+40o54t8lkgtq+Axp5m+prE3CxMR7yBhBbGzAiNjRk4MtWO4krSrU1sHH+
NOOq2913UATfDdJxjJsNT74PfvY9fPv8QDswpNAIK6hExfW0sNxCAhhruNQ+KOLk
iXXAZ15FnJ//FHHh9KuvZNhlqYUEdoSyLzNQ2O3iHUbQvh9nE6u0XYIqPIFZGp7Q
GzxcYMUP0RIY2X8qMcY3//bAOMQz7pQGR5HeqygSfBBzGKi9p5LdMWyKaCX7ue+v
fRJTIZPZC/GURjzbUXZDybTAJXmCb69TVm2/WDzJe0qZ+5tW3wQmBq38SDU2Edsp
0ulQ24PkSVN2KT76kuAgcfgM+ldXuRFlVgOKogb5h4yiwAkgXo7ZOjbn4SFp5SbI
wy+yfYg85xl0EmgeT7+Bn8fmYgqCv+ztcdR6zVV91oHkRqGZjcW2x/jMvAXIHg71
ieDMzowW/0Urg1uExJW1F06FmZ5rfQ/3cZE90rIwqxEPErso8UvC1kbng+Z5ZBf6
OdsRaRR9zM617xD+7Wbh5JN6Lsdzkz9LBIRhsO/pkZDmHZu6Ynj2ZxIunam10lqN
gje+JQ2P7RcB5IARAuc6gDHLPOMUBdmVvVPyxZ8R6M8hagYYQX1LTNhNyAls50Qa
d2n1kI/aQM9zRwG9Xj0N5hTJIG+WYxTgzMArKAO50dcikwzX/USGTz5CjCV1JMME
ebwNy0EAnhi/8u+bXeGVQifNySfjPXW+qWZb0GJ8h0Zx24NcIL6V2YvvX62YX8u6
R6cbIcKIj2J5YdPTBF8g/fV2RSVtICGEe57AfsMfY533pEhRuBWiIqoUqBkoGyJn
sHfledkt4i6T8QrcnTEYgS4N4iDYEamzV2zTm0QzqC1y/TcHldGsEvbGJ4qqHYfO
mfUZDCaeCYgoXmDgwR17sfHhkVM5c+oBRCYcTnSz/EuYfNVGUHUl3jTqFcec6IIn
Gs2b9fM2hKnM0ZoushKnEEHQgBWTxIco6Lg/0Apn8fYYsHndKC/KJQeBXRVLMiaD
QimSyYRVar4FU7VfR1rP9ERtXbezgW5WxPHxHLiN/4LnTsY70VDJUpmB4InYGXl5
e0lKxNM1C5vYG3/F8Kgbl7cE5SLmiOBDkBuouWnjv0CFMsWvfS6YEr2QikRxMJM+
YgpAL/uDAmJnwkHFHTUR37uiB5ZNnfCIhJec31LEubMjHj7AjPkPCkqYcP9SSCpn
m7CpbtA2Jduu/23qJ52/xMhE7uG2msAQQxK8Yhc3X+R7kwTZ3C36ydyq9IlBz822
JY9YVacH8rTq2S0wZqZxuNTWn/coRY7qXek/cZZOoyJ8n9WQvn2v3wp9znGGLdju
0r1OltTm0I6HQ8He5TIBC78rz/3B97ml29ONNmopWOogEIMoh8isaK6TySKGeq+f
M/pQflHnBvJDyTiG0HJIrugGTDmYiukAgH/8UjVI6jTZtt+QF0aMqtDFsJvfd+ER
/gH9AzfTzSN0bNRNoZv4afWXpoW9qNz9PB5xfj5tZKtK3hMWHxIOmmrCsPrIb7fS
1uCOIK6NHfrT3yFuvIY2kdgnW8vjYR547g2z3i355mbCQ/2GmEtsN0SL4/IGdWlW
YssPLoJvzo/PnFSu29222M5vcIaDWBcdy9BsJha1nZ314oUOybWG5P88DJhhaSUr
sZjftkStXAON9acaYNrWXDuUVV1wmTYvM9A3ePk7ncxUDBJLkiwqv3ylCtGsjvJ9
sq2vk+x7cvzd9TG1oaaFr9rQta8ySFQN8kQWDD8kHGGGcQcrxqDalsIpLc7DIF5R
JwaOnYrE2OfQPeXT1d4jtoIyjUJjs7i5cqLtyIXpvhz8oDys+5tZjz4ftzfLNiXC
Xz3Zwz2Grz5rKtBo8LlEQBNN8xmBC6af8gJzp/sm6kWu8Z/urPXM3FWzkoOL+6Hf
C0A2fOZLRSKlVPVsvl7wJJtvRNKCgtFNwv6mryFvodDib04hY43oCkPvSioO9iUU
F143DMX6LiPhhNbYa57EpDnBB8n0arSj6UflDz/E8KUtvL0mq+ynbbhN44k22eFr
L3FnHtjePLlHwQruSjZFiL5wn2IBr+xyKMUJ/LHC5N54pEA2YRbcHPSwLQ6atL6g
OX9N8pZnxizRDOQt0cIQOydTRWMpqPSbtfBCeTNws5FZkw+eP8zZofIM3zZkyYGV
YcSZN/Q9mtEPznL6QQ5iSGQYILLdam/jFNUNdGnx521XfW2dxJP8eVtA2CELazrb
0wbXEpbhUau6nZ77bDSO//9j/QgkPfbJpTDHesrsBnTKOln2RTlAYba4y0VTn6zc
+CKWWqVKYIowy8+Cr+tSDMS1oi4EzJTOWOqJSIJWqWTdSpWUbbCpGLN7SnPeHsbD
3XM3bmIQhNa52E9IC+CzwyjSeoh0LtmUsV3VzqF4NiDkuTEbNU2oKEiHDplaUw6+
27QiCSwgFxcH404bCBEXesoisA3gFGdFPwbBWu+doOdn/GrUqoOvY1ecT91HS6An
oFAG03QcpuhE4V702EIyCcQnah2HWSGpuiclgqMdfxsgmnigZb7j02BjGNX89jkw
gepQ5MWVAjw7WDWKw2Abp3wVp+r20YJlfGHcw4r19spKzS++0s9iJsXYOHZPJ5IR
2MRb6dKb2P2FpuPVYTmZgBUxhebukAfoBnukX65YND2Yt8kNJrGJRNCuJ/NNpDHL
vxh11NV2PkuN1/Ly/xYnoJPWidwzKRgj1FX7nwWIfTIx9Gj3vHdt1yGj2W/YWHwY
6iJWdFrWgaViCIvBhK5nvx0FrRk5xN+RjjFEmpVK+yXda4pJcpHiX624uS8GbNZB
r3eVAy5kfr+HAKOWStOAw3QlKJERJdyPyqQEkFQD1YzDKy/ynQTJOBXR0Z3bAeB1
oTdHZIf5WLvk0c2Tc67C4fl/utRwUTQUbDgW7CxkzCt/z74m4OpuWSNHq/jpr073
YxWlxMvqDGCLycuJjq4QLin8VcvjYLCV4VGW8rbly+JOxYiOVRaFfgNfMvSp3Mkr
jbBmcO9ZKxsKmS2FMItR9Cbm2Z6zc2oKMuBunTKM7+0gza8glHcTvtJZtzIwD3lm
rLSQdu8dCjzhuYxPV7QTd7OJpP/GnH4MMaFUTT6MGVn1kRy8DqImsXk9CToxYonE
8sG3/ZuQ8k+O6ikRwIdV/U2RtfDaPG+jM3p+aMq5Q9wGKFt+2FjYtyNtAJ1f64EO
V6N+UBF0iTLrAZcJCG2G8hTmTk7RtepSd6ECGIrtjSzGSKbBVRbTIbRaR5XVWPTQ
GKq82pyGBkm9PZkHeGW1HrY5KZw4NnWYyyd1OLc+brL+sshRnM0liOq+QmrVUVDS
8TXMRFqyEzjgHVFd58WcPJXRO+T0XAmqdaLZWz/MHrDefV+6cRhFGUplJ+Qhg41c
XrNDhGThxqyjJiQeZWeWgVpT+e9EOLeaqyF/BVDO9gUQemhki6b7lz0q0lOWbChq
StRgVAssYQvV1sxholz/Y/83nuvNaTVgZ1yK0eko8bArZwcJEAmb0Y5aASbnLI9I
vEqE4Elg7rsu7uF/q3h4UnO8FdJ1xfa/szfTTZgsVZL50RsQap3ua5HAQ+2Z5vlV
LtZ8nmA1ikXSh5EJZHEkhypDDNJiKoDXDmRxSVvCE9Sg+LM3T85mXNOGVbFNCmMw
FHNMlyTSiYJ8P+TDObxyB+uODIKPDvew5EitHpI0l7oPtQP7QRP/CcX998PN26i6
OpFjZAll5dwjOSH2+rUBYzA841kEIDhfaNvLXf0hKuO5ZEcVbtGBH1F5b/XwohRP
YlC0qipJZ+FupuKBH4pEXZHnf+E08ZMAqQwW0/p6NhNnfTWY8iFcQ8Ql9AxMNfaY
kwoObwY1WVcIoKQBjYZKV1UmnoihTwG1eKuuzbTKPOeTgp7c7/j8kyg7Ven9x3Ne
d/QwBHnDuyugpE+CZRCXsV5bHk2VIyu5AuYm8Vjs56bVup6HDqGtYag2BtKg3kpV
IEBXh44MmCIFDuTrqN2bW0B8M7pEcn2RV51+PtMORjMw/J9HquomgSy/exoqld1q
DqxPb9iJr0kltaBe+3/BCt/ccoh6msOvZHlj4iDS6CRC4hDkdOq20wqSNk1WCHaL
XhV6lMELvu/xeQbeBQVzMSo7ERiVcLMOJ+8AhHIzIg8/f3vGsGITuQkmqqFkZanT
6uHsWqvrTk/WOR8QbXPBe/IVV8Bed3jEX0b+GUKddOj9uR7k8nlN9r4L4zvqbJrr
y2hi6XBJFoyVBOzy5ZTBLkDJ9R6FBXEh8oJMw6m2QIO2IcSxHmCELYRprsR8lo98
YDFFnM0urhPVINAVqGS2Vvo2Weo0ymBUuNTO/5Ywai9k/Wq3wAyIn6v0gjsCTdXJ
lTiSP5xue6H4pbwjkf0an97FU3YMBF7zx1r7wyDScoueWc2iyFqskJwV5Pe6E0tG
EI1gQk/nVc0bgtx4pLzhAP0dA93vbfj7NQ0FthKPiB3LCzgr+RmqBAbVapcJKUAe
bJvgd8Hua0I4EJStNRpeIK6ossex1Qb1ABikYaDKoAt9zuDKjaQf2ZfsVlzOLOXx
bz/IH1a3TI08pxINtXT/iboNAos/MZU/o8lJgOMYWf8lTgoF6GGW1EqaAr+k2Yjh
kEQw6Jcuyuq+1lk3CLgXJo6c6d4Z1du41ENnuDQuE3PwhF8wc3IxfcfhQQsD/a5n
GN3npUMDsQ2m1SieCjuSEiODna4pFTCXlljhh6d8z3iVISwPzASnp/nXJcvqEJ4L
Tu/vtIJHU1n1WdclKQsPkUjGKYU86AEEjoElHKVPvT4vdC811XWKKF80zL6+UQXS
qBa8D0XGVfN1C4TSsYkD2oSpDMfJ/sknUYrgwUlunkiQ3Zesve4CPdisZO283r/m
jBZeCCgV9xhq+8ntcdIWYoeACc6uJJ1kAUjEVvtdRzkCrECdoaVsB/f+UacLTZw9
+c34TQnMfMgjQEC58VTUSNdR6hSbhp9iVyGZsvbHMWWdbzzi1SCiT7jRO1PetvSu
XPC4JIqYlPRbWCdFI9zaTjPnYeH4cCre7zo9e+lUfAOvICpts2Yc3XHVHK15giA3
BRf9BtlKpNtoRv0YHuwdhXk/WNEwXjV/G3TUOhKc96RGRhNv5aLhMZMVnwJ+LPr1
F6oWQ7H7cG6HW4BWrH4MUhvv5vAcbnu7PyEmGTR71Rf5ldtDndC+zBV7pVlajyWm
fKusDw1iqkvtZizJFDWJ0rnw74rfkOKdwmh68uH4SriOkVBniidWIU3XR1DLM1af
4kOYDL3OeRD2b3XMGuRBXsB8uFifhwujLylA5RlUqa1SvXAJwYNnkX+JeI13fxrp
wL/AK7RgNJ0H90LtVdkwlyidUEnnozUgYMlS8fafwb3sFyRnLnQdvtiB7V6Qprvo
rb0TOUnvGa9NNprVlcQMfizQsHrnSswKwLTnVdV/LMshObM8qdrn4VFpeDnDx+vt
aGR+s/B61zz+1hgy4oWVCZwsov2r926qKSjnA50T1DkutuuFbCYn9JEGWXJavSnw
S9Sc9uchCZKwQ/jOSjQ2hhHJcYrZs/X9Y4t4OsCyNo2H05jqPNQLprIm+jTlY+JS
Rik3H5xvcbadhpG4TGqKNROt3LrMp6se1I8F/+Rkt6j2allfUluKtH/iuvdJrfvu
Z52Kpc3XvP8cKhBiYhjmIMbo5NArRChHOVMMPt+H+BKcfylz7VtZisiMKdXkYcM4
67i4WP0C4Z8yXQ7JOJGu3qDK896ry2Ta4B/UC5xHiINpGqoxGhn8C7vGOQjmMK+r
LUsXn9JDqrWq6RVRqsrB2f/WMcFY6BN22SlzwvU7OVJb2fOXY+l9j78gw6ko8aPy
cqeVDm7nN/PoJ+czgWNl4GMjiGZSa4ONw4r+4PEuSZjTi4EcAiAygB7giSSVVRmE
SPddBCLohh2a0YAIPTVrKdEY/7txmDgwCaKwxI+w+e0v5d2DR8/vElgfKTRMTVqQ
M57yUvLUTsFrP41zlBF4Q25y3CKVuzczwVph0FCJUR54eKJHetrspLk70G6CDMCB
tT8btNB9Wn4Dh+Okavi+2WEsHD5fnBYJIkyCBLBkjYTMFaCGEHtdm9oZBLXkrm/O
Xqcmyp+6ek9oCjAHqC8r1Uxk0UiAXkOMqFfnCX8qkOXGZC6HADUSvIHJ6maljHIx
a83r6Kd0Z/hDdKituWoMsYWvPtgxyPkQf96UoK5hcN6amPJAvE7m27Z0WM4SVo36
bNUAWRdk6AMtxBTOMaVTOWQhApo0nmWusvkhluKPOV7JGwvdQQ2Law/wntezKWBJ
g/eI38CVeaQxSBFjDYXZgfmnJ3CfqOjSCEJYyd2syP/B1tguy87fSPqI2o29hGaY
1bZpotAFOGyDhChrW9wSw1TEaPbQR2EOcT8C+K2aMMdPlDqEk3qp/gwiShdAy6oe
khsCcVRmJvBI1E1n8haiF9aOAX/bHHkzygMXBd7ko6gRGQcVB1jN8ZNRL8CH2IJP
rjnehkacnS401n7v+bk6EHCEJMnHuyg1aDiDPwUGsTckld+ulETuJOAlYPfhbk4P
sS291uSd1C/1kmjSiufQBR4Esdwy5aaoxFK0rd9Qwyjk+ut/nbzm2yaBNpAZKOKu
GVFSDWUsC93qnUEi9icd+bU8WygRbCX946gF1YUfN7gPqsuVOJTRVoEQmh1gnX46
uPrspV5xuBSNdbDiz+zovBqmGiqDTXnRUEEoOZg9rB7ae5W9a/XWFm+hitRZ7wvH
ph7DZrDmANQTEz2wUqpwk+EWWc6Ee6nzWBvcZbF/nI4/gC7mZw8w6dQ3G2fZjFTY
Rp9alZlvGmPROAnvIdg1HJ8sQctOrimtMsnUnboLNcWl8RoNJ7rfhuTDahTSrqmM
sB5LVlF3DBdRxPZk7KG6UZMgyvCH+eFNhvDtg0nAoHGeRcam4Vx8h9BE3YAhDALS
e4fMOvMn+U5ShPLEJuhw406p7VpClbzw2hHs5xjNob0Rh/dRwFB6tTY3KWO44acG
PAd4IduuEFo2k8siuW/gfA4P3A0Ut/oPyzW4DQ28E1ofS0ym7Jg9NOBugmrAFW58
fZYoKDPRX+85uW22xBqB1GtkdvqZztBuR+/bTREan5C0dTYMubdLi5ntA5HqpQIi
Wm5JOhm8DB1WS8/Y0s7iuo6hoDE+LFShq3xgxhrpe4nd/6RomXJK1WQ+rH/H1Beo
9gZ/41q263B6aG3qMep8HRYOXH8h+24BZG9uKEIwI3AoK7Im2ikFaXGvJIcZrlOG
Y/ots8PRsDJBKfEf368o19KYbLV3+8p4H0kD/lPZEjgaBWF7GFAweQnBGlzrgxUz
aAjJS/bruV6uh6JpKqtgMmwgVeVUyxpPFvnp7JY33fhnPiMvp61OyQbVkj8V38ZT
ZAMeRmdJEQx+PH8GsSL3EUe4+yUMPnBdECZPFi4nPIgNAX2Nvw6adcVKBEkm0KZ+
UbYxsDs5IRb7AVwOjp5w550M/wf/J+3EfpUGJtpbsGYYhNEy6TSCNNSBlaTJSMyu
8HSwBiR1askkMgR4M9Ueb+NVyTz/lql0stSY2t+yR7QIi1HySjTEPsVXw1WhE9VD
lz92jbxcumJF5Up2Kn5FYW1MtmNmp8zuwOJCcXsNYEKhWrmICFEyHbwtyMlh4/il
SY1rIpy+VcQeLCZk/cl4eW3VDMm+bRjRgtaMFHhjuSx43nzGuOTLeuG3Sx9mHL+B
X7+UJWZ6mm454pXN+fMY2FsA9Li8aqQ55iRwQltm27xsF0mSXZ3Eoj3SS5txEtF/
E2cblWhbSr17LFBHNS+/N5Cu4gWdrHROrmj1O/H5vZcSUB/Gs/blpfnI+B7acRdu
Fjq9VmKM197gNFRU/KPoTvyPJnuNr+VcuzlzW01068ErSGJVE16gB7OPj5OFO0jp
7RDahCZpJIRMpaRe8lxdfU/mJ7/gfBPjthRa5k73J6J507bcprhc+BB9uAPGDGSl
Fv+b4oRRycVuAx7v3iaGYnh3Sk1XfehJ4JvzuMmAxEo/Wrs6Rf1gndwb0y27w72Z
Gu8WrS/zyBzDeEskQKou+sGWtf4UoSqPFdTqSIo7a34HY+KEpGTAHFrX2dvVwsOj
9HwNha+WOx27daIfVF8BbWY4Lgq7Xk0GubpLgBPMQPBWxDbhNzAsR8cZGgdjv1Xz
ee6muhqzKZUhokhTN0hgjOV2A+T54R4PyQ8Zg6hIJtl4rY2JiSsBC1LYQmJqsZZV
nF3CuLny5tA8D5Bq/M/qJXEReq1iw28FBXcRqJ+CTNBNvF6lIACqHiOuo2yeNbf8
NAGDhusJYuRT8YSrZG25S1dF/4qtXfILjo50nBCIbWIMEU4Y2+FST8zYUxoRtsQc
AWtdJKlRzOM+TAtzKWRifJb2ptauMvNj59LmF0eqJyld8fEbLZuY14OQzRNqRgSt
qIzbplzqj4hJ+4cQdI1PYX3vXMcpiz59H8ra7sdVTNLVB7qjZydTWxHm+BeJ7hl3
m79WNtdzyTtxhYYpx8tumKjA9VD7EJnfKCgAz5CR1/zxLq/nI/wJX8/Zs1TUroQv
y5qvKsS4Udt4GUnLJmx1XFz027fhtrDiAnAz90cTa3lmGONt9LjY3p/RZR822oKP
SFTKbmfPk2L77TQgxVPQIecbLsq5tjWb6ZVJM624DqLaJS9Ji15P62rPY8QGo4p8
lO4E6Vcnolon0SiqNvfYEyDWSxT8g00ujfkdH+iN7f8fwl6qsxmHJqG1/1+IMTik
QUxb0YoaqL6xEbR2K1//zYCc0tKKJE9xHTFGVhB9Qqgsya0KYo+uiFtdq6xNaC3q
iCYNKhHIaheixNv7X33TEm39vI4/8dtXDg5ffhKs5MTi2edX0/8R2OC2xizQgt01
OCmuTfGaDi0GfeyVxpj9QtakoBK0LSELTJl0dW0KuA/bk5qgNEZ46MiQWcECmXbv
B0oYBG2GJ0IJyu4+qPRM/NE1DbmyfyGmKzSls17tNNKHDWvb6qUc4M6diw3ty4zN
U9ymI8Q3A+zV0GRg4QFycHTLsRtvp6Dsj08CIuc4DKDkUfGd2zH2KI+lU4r+CfUL
SEWGNkmBq3/Wnr7FUb+cn179g1nVUEyVFMHvSSccm04tx13byWCWrK2u8tMlLouU
QnzvGVsPXMvrryFdGWHpmVj0Ron2dNX9ibkXdNlzR+HmVoiyjczeeyc3iq5YO3al
oJyv+k0C+LeI5zc2/EaAwrpfbnR6MHYw6mK/YscDetNVi+o50rh84uKJKbSoXjE+
k37eKWArqAmrY7DgURWXeczQaq5C/cTMf1sn3CiOj1eekgiSjfl5fMFLLFtyDuXF
HQ0SjzD6TAks0qKDcfW/4o4X6DHcrWCp2pUSnIdBi9dL9EUzd5opQ/vy/p8AWyQL
J3QlnlPmQTaSpnzfuL3feei+mJBPUvttdjt83bThlFi0jsN/3J6yAsJoNlFunO4o
93lMcdTkHSqTHgPD37m/IzwPto5F16I8/3Wtc6dvd5vGySS8m1ZxMEUtwTMCSug3
W8D4UUMdsRBeoycWpGBsnIXP/QkaDffX9WdvGgSRq3Ljd9guH5nSgxOS4OC35rBY
e5FSyo8I4GPaAVXIPkh06TpldCgn/NyvpMaj1sfNKpCXv32J2Rzrf30rrm8XYQke
33CXb6pq3mPARohbJyLyN5Tpf0FXE9yAor9BLPFPvHxFlBRIOcm0xGFDmt2bLZCs
RiksOQf68QkUZP99mXnXV2joEhwdxPa5qAfNve4h0fRBCstbwtxkCoSQkwkgOyD0
dJibhqYrIGQXISk1YAc98Up1KDgrAd/EbltXe/NWrIUTp7Io6pWVifl+3A2liZFg
jS+axckqF9Ol/6ZZawL4i4uJz+7Sa0s9XaHXyMhJn9at88+LSHFXZ3QA2/I8Srg6
QLqFGh2ziXYEOWZkPdJ4wmICnFAWXsJCho4au9kDJXdqPD7dxTBLSo3CofAyua8M
bCNyjeDD5ILJdt96LduJQnfdQukxlyoJ/NElXB9gED58rY3Qd2k+D/bbefiSJFHH
1B0Hea9z9CfebYhQaN25tFO2gNkBUS5nfHxV1wjK9AbEt33WI1zwHEuWJDlbf+lK
rYkJ6+44u8YwHIkkdopLJrD39pwUq8t9ZPsYa5f60jNeepiMqBY/v1IVLwv09tWh
iWn6VBAKvEUiX6tQv1MvUGpPrNKrP1KzNIXnBcO3vlWZFLJ4/cBUEbuqdZxWFPD0
XgK3UQkJo8BjsSDPWaJCv7tpA0RaOBfASS8r1C4rren35ufDlLkvwkBbU2JV90YJ
Yl1rki1RsCPeUoWL4CQ9Qwb14AmyZTbmGEsjqW90+iZJJCrzXnrKcwzUXLUDBSmF
oxc14oZt8EUv0rQa0+9P2Ju3qU/OrOnnfUVZWa6+xOHh97NwC4/9tyuLMiBr5jDj
ZKxkPFnGSdmhR7KAJ82AWUXnSRBRwovSLix+2lHwlo5essA3UH/d8vVFJI1HUi4/
PFyAIQnTKiTDx6W7GSOMBjOn1/i8cw2epai3dRxheQwGBhsjYjPz4WmS3GiAn4Bs
KZF2nRsthAFB1UMHrY5HhG1H238pem3WGFwNDRCWq+F4bQ7mXuQpu6NFF6rB+Ecu
xXSjVKBUe3JFAHtRZbbVxAkiCn76+E1qem5jCR7ORGU1ue0iHSZWsdJoMwaVVFrR
S3d5goQGWCQOjKC3oAOBQygZR9sz+KUTr7X1V4fdLd11xQ0hB/eSFQ5V7kWQ3xG9
VukaE1t8kbTY5uXObzgz7Vqgw1/nAd7qXsh06bMus/dn+Wmq4GkYmfFRH7us4dJ5
Sna6chnJkmenWbBZG5m0kiYyTm4LRCju+9mjQF4qOthQNlIxl9UON4imwoBZZqKi
H3doSdwSCelLupxSAwOLsFt1VsDRQYLGX3e3O3vgJrqzeRHzM0KsfSCYNxFU7Yfz
c7jCQ6I8/p0ara8V1jj8oFhMtL25v7Tj276SgI52sPljRaIAc/6D02mzrRYejLcX
O5rpFd9BYrg7OMB6HT1AC/usqNglqYS8JcC6vMXi0ZotSqcEj9tA587LPrbewM4N
k+Qo6vzEQOqhfokja1rrtF/ivG4Y85xxkpi/fSoqOX1GkU01voFTOHKOf78mR5Dx
0TCegZBpeOCgUQUtXnPazUcC/390JoQt5zMsothnxmpKPczfa6r9H4jyYTY2renT
lPJ022O8DsAM60PP4CHiUejaRfer32WmVD7GytedWnPGtU/yHuAZ0Ej8NC0Z5MpE
Z7JqnmNQW4spYeLTbV+lTyUY81qC16gXtBIc5+Ddj1jMGC4D5eoI8xzWUBAmUNvu
C9uf11Z8VPo/vel0enVfpEIxV4rxWoRME8qallgXoTRUSgbYuS3KVWI/TCM/7qZV
o6jwd/vxlxhMoyz/rEqqEBvAahCICFbZm4ioGAhSJvf35qUMG6uNv7f2M5XLWNky
bm2ErXuve6nQQgxJcimYZLhmsk2QXjZlQabzqJtFLRTBoz7TzWy5jRbQrEyam4Yb
LKKn/UCOnpzxTkV832aJeOpKabumJpBaT8z8oZ1gcPIMPMvGZTUbnWXug0p2oYrf
ZJFQo7yaVJBHCcwwqw9ZJEz+7rC+W2Lx2Pw07QSbKCWcC5rqMABKKSUj5Myr4Fx1
h2eqIcnhrdY5F0X4LWy+W7F3xBLutRMiIs37+wUFZCeToqLDypkiAlOofZ3LytEU
Z4oGfxi5FTKRpzb0yMKH9gpE68whzHJA+VkGloL66FnEkcEGbvt0FyPLOyPHu6S2
6DO0p97QZSKyB035W0VoFtLC04SoE2i5DsTUVxZPBy4Iczmqj6C6qQ4wr0iFxNmr
VzPvswa0rs/eC8ZmhOa+AlaZb2hlC5Ev3DfdSYGdHn0s75o+QzfC9UbD9uOFf4aZ
SwRFmZxHhdkeGAzAD9X1rD9WgF/+rCdELa/vTB7JEQ04f8mvP+h3ur/53ODbRTpa
nPw9nBOKAN7Z9m+pNAk6q1ubQsdXCbXp+AekZfRzKe3HhOPMGcadEXSKaJ/C1Myw
lAc2oiRZmgH9/ShHfsMH/Sxle16opU1W1Kjf3ZmsLgtMYjVN/Z+V2i5WqLcFf7uW
7fACY0zPKYOAo5CZoyLWD/YfDQ49SRP45F2ppUnAi6PPPb6Qux1jxX8UR+IMGH0h
4ZpLgycrYffiiOetOhgkuL/Rh0jronD/moEqKmy+13DNRSmpm4KKaaOSAOlnQv5+
fbwn1lYXNXY8vN7swMwxI7gijFdeSGfnFUTLW5/GyDVG8GEB7wi8SJBlmiCopb1e
uAFVQvU7gQkV6GKNFQx7cLIC7+MCknQ7ai2kG6h7cGESN2WxVkDb/pFzqe5VNvas
ZFWyIM3yAdqREIwmCkAYox9kWIscXHVgNKxq0OOpmJOdiJJNgCFMEiTKRjDJ4y2s
45bdDmaBchchcRxCPseSB/Epc9r5WM7j98cib4tgEX5b7gdneEc9kEXHq3/y8x6G
UTashpYC0cU0fD4l66bRoZeQc62ALierDldHxMR26FwKtXGUDDvofAfRmCDSkhqd
EkQzKN3uBQ/kNHDaJz+wsG0qK6jTQObUt+wOoaEYxIRrCsLyabuKCqs1b4YF6ZNK
uqh/+7/myHSIbyuwhKxFIaZvHB14WMzcx7zuUVCchF0mc+6WHfiqUTMJ4qjDNn3p
6q9w9f5o7l4FNXwEswP1VowOt/BVgERdgXJK7Jzhh8uGJmjo2pmgUYZqWz9lGhGO
wEYnGOcaWCONXdzcDzbeinVTjMBjHWaCE2iPRDCxhPwIQ8eEzrfk4EJoY+WN6QXo
CCPr8WiBztT72pbT4BG7SmEEOoXHiq0dr4LiO9h661uKD/qhY9Wl6s/ZR7fln1GU
Ymuy+I4wHZIu2z1jR6U5LNU+jtZhVcfQl2BuZuZMOtIC+azMQVlA5WENo8qFVRid
BO2aa5nUQUMykygZz74JCL33WYF0gQR8aJBkXcMhA5GEBiAXv6VQHTeuEGBYHOD8
J/OBGYLao/lPMHjbZnmYfXJaMs6rSXdgo8xHAKo9gm8f3GIGW6fjfx1zNIvP+GmZ
akxudT7gvFr+e1KNi8JVu7yeEPG4G9QvWJjxVZhBabnrKdKs9yzwUanLJNwNtYER
yVSt7VAKE9oyel3s4JUwKEkUC8noS6DTErOVqSuoq6UQNOd+tVpPAPHPGiSH5iv4
Klg7poXE7f2pVhKFdTp78bRv8yfm1jusl0EtmHTYHPA4keOo6R4K1x6oJBKPa7VM
V1QNo3nyd2PeekpUJBIOPn/ZsToz+ROCHuubbZC088ArcRolteWIYFsJp45xX3Fi
c88owIWy8bc9tq6E810riSCIWIq+TrlXI+SN3k4Fc9z1ORylmfvuVxPPrjAxUut0
Ia7ZfqzSy5lI1/8b9lG1tf2r/ADLG1P9TNufF3U6h0Z6GZrXdBHSL/A7utUo6cJ/
lzsnG0N/+YvAkSWyBppy2cVsc23VSXQJ4TentVdSIqNcq6mJ0kJLS21RZT02EsK4
6cOKPJjpVYpttbsdTqWuzQuGzt87MXBejYzA9E72gfhebWztWpPkYCYrQgSNufsn
Z4eqq8mPGQ/q1FaX+NU1M5mbzXsX6VKrzoC4cxnZzF8DogkNrZhokSV07f5wgdCy
a5ptFwFVy0tGZ1FkN8fM9dBVAMSoHkAdouZ30qp3ecX4eShWn8s0/EZY8NIuE78V
EzhaGpiNxUmmd2LLbv1sLtvCV+62AVj+CHCGz4gdnmQXZiNxBLXHgx/w6RGiP6tI
ptngtWf+PNf7pgqN/myZQ4Ag3hv6XN5SbwahuXymfTk2rbIGeQBF2BoduZyCNeaK
zyJVeDEpjufBW+/fcuhV2IP3GEgLzNDbSIaRClhPO66Sc4Lfrhn+Co7kOfYLg04M
95KUdBKG04NaIqkL6jk2kNcWoVy5eP2c7oCSVAgtbSJ/pj+OWSygfKUgPWmg6QjC
Or7nOWDarA6DgZ9D2xs6fQ4jfK82Vhoh+NNpaQpfOuEovmXFKYjsg5pw21QFVnOl
UmT7v1QMmV55yoX+pbtmapTOIuXnonXz6iL4n1s742Ig+L6+oXtBzdhOIS3TMrDO
8ZBiVoAVp9qb/6RaVP6m0OW53JXANVUuLr04F68yiY8JyCw5suoqJU1dLypnAPfx
igq8idLx8fBUimSAnGYY0kOs096tTbA0MCa32fdJxcoC+oQxMvX4JRy6U0Co65rJ
Nx5bfQfldNsb3+DqsXZI8LlDbyQ1CFeCAAWzEeTxkCBTynX8xFEVnTkJ58EBYKlv
VTtlodKdB29sCDnNDOal856cPGeiF6rqgbpwke2FLPmkEuouF7PqgOLnR7Sc8J8j
L/Vqk+v8LN50v0CiOBOARi7hWLS/0WT2hUl2lbbyA/HN3mPaNwFXD1SxCB1vm1RS
6Jx7UrDhyo8KVvZcXXVDs+OlWFOkDSEwhlx3X0Y7FsgwY8wT1YccdUe7+cBXHoaF
Y2GZN99yxjVdpvocKLVErxvnEAgrcCBFqpzqXTyiarugTJMzDfSn0aa+i2lz0a6Q
zDfldmDZoYZRnaAcm3Sv4Zvx0uDHiP+16/niqgVFD7rQrbF6v9Fawtr1oiCm/Kdr
PkxbffdILy7Kmg2TEFXZSuSyKGicRBY1DUTMHlgNZ0v9HabsDWR1AMvzF13gBitO
RE3//1a4X+2jTmBEBOE/fhMPuNjUv542ZfPGRWHs4FDOi7/HQYyLdrzzUl+dyWvG
9P2Am9A09V/s4x9ZA+wrtqfa19bxk0vxVA5HVdXpqQLIrKyTBwEZabsl9BCF8coP
ddjjNKK3DHeeGOjGRx0379Qcs/abSRUKf7vXGbxHifEEQa+a/hMo4GmxyPlpUwok
Pra3STvEro1JP8GcD5JwFMzm+9NpMM1V6NYvKbnpa49ZaC7M00QdZ7GdP8fVb5yc
OOPrK6AjcjYIVLyWt9QqWmnrh5tBr/bhP2nEp0ELro/Ex5iVg7B7aXlHPfPFA3/z
me2RnIRW78UslV7FmFIruqIVNO+h/oIVV8i+0Q133m4yWYA920YK7fxp+lP9sDnM
Q8V7sEwMcE/9n4AO5CITLd/gKoQKnwhXv+QU3NjJj8dDhCYBnXhuXWAdHdhC1iy9
AJlCPkHYIvrbY3DP6C6OF5uOWsMzjS0PfpTIkZ3Z7mUSd5wo6oSD21yKsOBGUxzJ
6XV5vm7EKHe20AEeB8wZnS6zr3vPTpU+veUfP1U8M2fKlTvhnLPlPMxyakQJ7eSX
/33bI25N28PlgKqPpsheg60/n/2BAvWfUECfgGn+4oJu2UKAclKXoJ/50iqRgZqL
a2Qb5tUp3mtZsdPwb2PG06ZAv9bKhu4L7xQ3j08gLvDd7I1uiCG0FJOUuauqeYtr
kJ+Nf5sdQ6YBZi5hQ4Cm+l207FLkpAWsGEjxZVOi9P2kyD7KHsoPsFsLLNb0gYzN
JBeQ7GZIcie0R5Mv71XV8FNLhg0H2MKJP6es2QpCAfcWIu8SLxbInbm9CuBM8Ted
waK2RkvfVxOScGvPBlZF1zPFs4USYMBykoEaeq5s5Q8Y1i6IAPd8KHB+Pp5BRF6i
p29gCeUeCrbxofRZjOg8KG9WnJVwT7XSbqN0B9Mp07h2RR1LzDI416eHG1ySrWo8
c95NGEjYrXkVtjPZa+G/M3yHZy7uFGfJehfg+vJmmfbN6L3JPgwE7QTtFbonQkk2
wXmyx2PNvHYCQRT+qI1NHIxzpeMqX4mH42QrXdjUsHxFHlHk+NaXgFW471Rqr1Z1
D0MV2KEqUXU5fde9GkdSm1wo5PH3bxg1iQZOUb5lDJW/G/PsBXROntNX+ccAPAly
Qq62U/Yl0JkeJXxLvizO+fAgB9unKTDAzIgDjmUEg7E+KDU8EIx+RThmRlXywA1x
x2XhmEiaE0J8EaRogxopzsIs3WGZsguvf5/9oJBpBJUBP2s9sDn8lmSZIjOBdJMt
VvhQDesdFi0x2unNkvdqIMn9eVrXeq9asS6tDcso2CKVvfq3dBSwwWBsN0oQJANu
KL2nFXbmBylK1KgGWFkRG7t4wc8xQO/5rKvmZO8qkcunKSBvH9CrH0xccczqZQn0
wCsiq3EPeUqHLL3a6iZfdu/G8fB0ndrlyx3aUDW4bykkOxjxjx6jR6hYGmJfMiU+
Pc09XL9jHf3fgU9oe5rgzp78iX4RD1Nk5jzx9uTOtFNlWfQS+tUbVYpfw/gcqA9T
iG4I9qWiM8u9zqz5/jGjGcucKs+GCJo24h7/nCkMe66dDQBxhxuUVOeCfNp6vZYW
D4Vt0pt+gnIg8Sa+j2o8Fzos+Skyl5/ITsb5JDwZiwB059QSONiRKklX1VnIJi5M
eMs5lDGNPHIEzlLjYxEymNP0p4mmw5WP7pb8+aiscQShma50MXgDXmW+hBJiSxNO
Di/GYFn2MyiMZAwZ09eH1xxKZxH/hEau9330LW8urejImoqAbwv2P+ta4UNBisCb
+hpwcExwjUGgmh9kY2dQ+HWg4rHxszer6GTwKuQZ1oJbqqTdq/WJoboWOspPQs66
Nqn8beC/BqT9meQ/4K0Xo9M5xTzhVPFunenUwrG7rBNGGcteXRkrxcZm2D1uIKTg
0mKdAQ3Ou8JVPZe94Vaivl8MaokvLK2TkLz8Cr05QdoRlxt/yvYht6J7OOjQyjGj
B5Dgi1ZhFQa0ya7g8K+QZ3n9jVG2WorkJbe23/WJrXbAe53GG8HEuEejLgnJdkzM
n4P4rohMxzQPW8yH3V4xxnfjNxF5NtrnY2zVvVrqbHFqjEAdSHf0h6uPwGIE+Bza
VnuohZiwpjAa0EkHOQ5n/It3e6SVamkD6cF0JlaMZXO2tohr7z5nxfI3qS/b8R1R
Ep2WoQ0dq9Y7vsYwXQxeSk+VTNhxjOFp2Q7rx0drNUqn7A7t3xaP7ns6JwJ46HqL
ZhhTrzgjkXbEzI3lBpG2k0nR6SEjDyA6HCdVoYwXCVKUAbT/gJ9eTv/7LNQpGtRy
emjYpBkATCcsCLCVMOLxfKWpSzCElV5kBvZDqIVfTSv30N6YTX/nWFB9mO8Sixv0
s9yS4KjcNt6hd5QnLQV6uS+ZY/4O7t4vU/fSFqn8Nkknnf0Av+GPsobm58pujsss
DX3gWdEjz4UheuM2nEtiDbvSPbN9iH5vwUsbg0f6IDYLaJxl8Jyw5VlpGKhbup+q
RdScmCn5T3gBwtElgygkUtY4ei2pLJV709J3Ql2ias6wxGKSCUVeLogCTKiWpTv4
aVVJsPDZ/AKT6Bs4ggavZkdOlNxk+5NfO+xGNit7Xgsyfc10jnm986eD27gDtTKd
UiYrf+V04TL98Ep62UEDhZpcGYNORxZJjS7LRlBGi8T9KcG4EfLrM6sEILLHjFK/
2zwUo+NF34R2HqTMZly7FQ9U1bATSM2mRoSXQKXmkOG8qF3WCF+ZaMRHYGNLIULw
ng9axdaD+wiOzuUNdqeq/M2gzHYxasI21nE8d2eBgC1GlDtAwk/wNCUqEp+U7KUK
Jd+1lMcVUdNjhB1eLVo8bnAbiVltr4x4Luo4U3Ed6BNoqIiNVAazhoRxcB5+1PR8
Y5WHQ/09HQ4LaBt/6n9fNWm4xdZxffDNcArKddg6vBdgHqxP4z8IWtZSjvmvhzK/
o9QRhu3LxWJb7+9LBxdPPtLEC/mzmcwQjOYVX0QYxCmrUphn5zA7FtDOh+Ep5fkY
SLArcrQoQLa//QuxQFqUUlODQfpGnx9pTsiVuXp8OXSpq8cyU/ElvjapdoVIrdLz
C6Urr7N/LqcQu5PmCu0HOztqZ0nzMAd7j10/7rI2FbhmTBRTw5oFFJ+qm9XRfkby
gvsp3EZhBPnIznUkYOU9Z0XVeaQ8kf8iQHs/fUs7Ygkbf1zEby7A5Ql6WJYiAx4H
D36KkjKtIheJQZ3qqes/4l6nGdAIobirDUt8816ev9CcMC7KVWHMDTe7ZrvOr94g
FKggTxNn9elmpD2MKVqzw36JWhjcAL+Dn5D4FSrpEI7hr5LOq17mxr17/4ca7vlX
pnnjnLHpXrj56LGdD6eYUVU/PSkTqL/lEBvP5uaU29Zf8FE3TdX4fgfjORH28Dw9
3qZAZnpCEQk56l2vkr0iMrVKrX9VQIcpNT0lS/WHLd+yBt6xBvPQ+UfA2aJ+gJHb
EFFnsH/sEfOlRO0b1VDfpoVV2h+nv7H+arDvtTd8xOFmEaETDp2EdpCTGnd62u3W
zmfdQF1rl/forV6s5i3UWMNjgSpKiFTCJS0A5T4al/RanWY1oYjLvNaVnlWyGz6Q
wqMyg7rnzuyvIciJBBQ4sTi5DZ6S2Az2klhh3AoR0BnU0XhF9gySksdcspcPbHx/
+Ky3rl6Ktj92YinwK7N8k/ZXM+9g+N2XilxooY2aWgiyZIJN5JVdg7NoNfL8Ejnj
xu6dL4s31/5UYuQZFyK7tYH7S+/PZ2IhEti5OVIUdPfP2JO0aKU3WxZeUH0DNQuY
k3KlQb1t40wY+Sl8lliq7yHRD39kFvqzx4vc5MdTGsAhbkGPnbYJlJezSj811JC4
sKq6bvv98IMtV7nOAQtc/p3n8CmL0wPFVggMDJ20Gf9ZnIT6q/v+mxkFYlPfeYMG
A5t1LLDCeSsDXxLKBhvQH8PSsgxNdnf1LChuielu2QV7nmSKxYHHG1AxqwtbKhIJ
r1lge5cV4Vmh9rhLi9p0HxPtZDcAf7dJgfot6cRjLdhBzFDxxA8yQY3HfC6klPcX
wdVO0g9HOLLBxrNqdai1oreM7JkdBnxJvWxys1++yYYgzHRb0HDrDZCyDAIAcYug
4d9LD0oXVWOUsrQUseqjEf8X4KDbJgRoa4Ej7xlH4JB9ohRxA+Hly7hLDGSw2Rhy
tt+iUKBGNWaAMmgFuJrM8LjqzV2MB/EtZ1PvhjR4YujgMwICl+X/nVg1FdKE1ROn
EeMbiPpVoWmJMD4oOT6TnwsGasZd863HD/ZAbUKcsyfnvLaMvmEu3ovy6SyFk6M1
eWt55EzcfdPTSJ2xnhLisV5IpQOeg4cnKv80izFn29BIgj3cyNy3SUTuS34d4gye
21m69mrDKXA1rmXQWcdFR0ADOXjG0h2rSXDrs5jyehPBuLomAnFt37b2Pgyj/ZM3
DdykL+Q95vIEeKsDT81vX0HhN7Jx0A5lhgJWJC7a0fV60zjtpTFDBeyIpEzV3Zt0
3AQ7XQWfsiblAZG0NqB3dA03aj7/6SVk1/M6uwKpE/BsphRdpZshgdv67nDIiAK1
NKwLqejWxVAwTe12fl0QMdoBzSOjs6B2MxvjBT4GXE/AgFESsktv8BhcVNCkaKWY
47lDyfzi/jhkLfYaeFJbVJgrVzBJfnuW7TnJY4ka60rZC+4JiqOcoDg8jHm3tMq3
RBkVt86Fq3kbolT6Mw6JeCpvfX2jJ+2DO1RjwFoPPMTrpWttyQiGKaE6nScnvwIA
F5AeHrjtmbJ8ixmnnIPf1Nzjq4mjcJ9J283caA9q+90YxcyINMBRTz3JhfMgEkPL
VK6gG77mUuPqSWj1s1Zm/FCfr0kXXstYGxDcK9RhVG9GBYh3tah8nUi0AoppJ9/Y
QMphmNPzhWLcb9GsnEQDRQFydePd/xaulNZgRSMgMkXEW67iQSiUGa5Hi8pGf+L5
e0I2OcwnQtQruZNt6kRUuchwgYswteAr8qycP0QIq4pF1wunKQXz7YxZnlQIsP+4
zt0/l7jfnifmJOHvu3WSnw6BwiISca+v4qCDac7kAsC6ZRnfS0M2haXe/v2jXtLu
bW7wT7IB9wNcYJ5pgNHgGibUul19YCBUfBC2KzBVpYvyK5EZrCQK9lNSeH3WVAiT
5QZ/GVIBQFjQp6qN4038Ea13qmywYAfF4Hiu2FhfSKhq85dLS1wGWx1N8TxVtTeM
7FfoUCzHi2X2IFd13m3oxuzH0Sb08YmZ4RBmvzjWX1oUSl6yIFQyk6tPgZd+dwIR
UrMGdaAb9Cv1WGfhRyu3uwoxo08xib6zKToVdpNDb5Y2zO3eff9gXE/97k4qGaYI
DgSXQwpSRQH2sEtn9jn3aggPsUjagehMlXHTa4yQXASWgS/mj1R72GAGbE99Wqmq
zs5qV6vL667/7JdRCXc/V4nIzZOwQfhH/3l2Bs7QnqDU8VjiJgkyrZfCwdYj0Tkg
YfpBDVw7HKlRIjwhhdK2o2Xfiak1iWUdBIgJAHSR7tGf3Akb9iTV/8SWBNo9vE78
wTQJRCU2rEV69mMD36FIcPUAVgpyU/9Eo2Ut+hBeRYWgvEcqNwiLD3LDjMZMfrA7
cTOw+3yuW5uPzbmtlEVjCA2Rei4Ag1fE05BBfasiveF8R3L8GFl84Vu7WU25fgl+
+zz14im6uX4rMyXpkZ1NAatMiwYBAUraurjwix96oV0EK0G1m/0RXAoYU3Cb6TvW
mjmufpqSF3fcykMnFBOAYDpbhitQn9QGlaXBNz/UiENtme/rpE9n72QmdGybVIBQ
fGgFAtpQjwbW2aLxv3VEvTIQvKcWB/4NNM1mDR5XMtMo6ZjrjAfikUlXesIMVI7A
ieIfR/x0cBXTlZqs1ru/4eC9jGwC7Hz/HMvZEv5/2Relr7bJoAEOkBA7qzRdbT51
PhEkZF0shQ9CFZWm/0J9HkLLv5CQlLIDcagEd+0PKb1nHpwmax/1f8THhcfEJoJG
09pdvkHwuuKDZTF7x0gz8/RlmMuHEowRtTKQO4Uw/Inl7l+JQDhSp4kaR8ZLPDFF
pFd0/5EeI7e34wZSbolUt5oz3V6NGK/zkhLut7C0vf6e5HkBgq9x3uygwXlOlvAK
0vGB3WirHIEEJobe0NSarEv7tiKXCN6V27pz2tkwelUM1fq7rLbyxQP5gnp03BT5
+Rd6Cn/2LZzB7KpSc47N6Oj/r48r1KuC8D+8dO6t2Ed9rT2efknmuLGpSTxec83B
yELlUSdWhC+tAeVwY+RY47np4o+Wb/VVkFkG+gOE1Y7YrNRoIJFLxXfykJip5be2
ygb+cbmex2xXn4mC5D+XHBe05O1EY/8aenOfu2XjBux2+BNuANLQI4ZBpbbE6P9I
a+6Nr9uYy1NXIpyVWnygZkcc2qhHHzHu07h6XG0cBQCGETAo7i+FqH7v6ZVeBP2+
9+mJdDfo2tQX5B4XIaYyAYV8GFyv65afaMxPghetrfvmcTbLCSrtMvyDKWKcvJYP
LMqpBEVKMYisoAkTrM0pXtAVtvWHu++c3DTBS9PyUHCBVKADOOkYhEJ6N4wbWmWt
hMmNw2U5gAu0QESW0kj2L/w/GdYXRi4Z99yQnWiaUFNxsX0Sc8gAcZyLNj3byZ9L
HER3aTLj7eDb5rCqplJjGjCF+iO6xBEUS+MKGcAhfXe0z8lwpDD4lsoAOuyewDu4
7iZtZzjO5y7lHefhtazlalORd4tidMsEpzo+q2CTYU0tXjiZp6e7QkrAFdJbsFcx
RPloYQd3IaAzwJbcmRUN9TbnQr9Fze8AguH9VvMzqzFAeaMdjQg1MqeSMrtF25RP
VCy1th9s/OTeMuite2evSMYR1t8q0eFJRbPuUtVzQVDC+fvDZlrJ+N0lENp9MtfC
Xa8Q9oClUWSuFWlAnEVO+BwW+gYJN6DSuFWoW63ZKOLg9ije75yIQZOHbqww/Ba2
W9ixba0MEx27HUWY4ukWpmkRmASsctB0BYdve5M6Oato3wFQjdPBHn8Lw85xImen
l6cbAl9yGCPCUixQ2sHwQhpKkTvFF10Mait1E9sXFMEMPu6e1nJw9M5jXJrAaPgK
aDwYrgRrDuyPWPAOo8vb9GWwONp3klk0m/I+vWCg27FTCgb0SP9fXwskrS41TN7y
2H162AX7XcXiAAmBhla9Mfy+z7p8t9eQuQHvu8jqgo2zA09MI4+R8Hq0JUjrLB7A
fMYyt3+fCdZxugZ8xEaqkeJNk5ihGY8+Tgwg5cQYReTYVNEnftYEzNqgIvo8w9Iq
EPg7jJ070S/2jnrz03LSJ3QzzRDm2rQJUKl2Scz5QI/wi2XFLvFGuXlykQHPjzR/
mYO21JK1Df62vHGX2ZAdf9M/RW+zJLWW7JlKkZMg23PQEN2tTxB7eAavWPBgdwxF
sYXgbBSWlWyzzT4q/4hRxKU9WQaTrsORqD/w06F7k/6va0sdoZdRgVWGWKDUCK8f
hp6gsW7Lzi8xgnGH2ELDr7MlFPg7PJnAQJV/zHg+jBgY3ujlK9IMrwHT18BTynN0
jIu5oxcfkZQcTyjbUcOg9zEnfpRINsq2hb9jp/hAhBlyXGDsqkh7ZYm+Aa+H41iL
11U9OtjrhaQuB88LCWappW1Mt72hDB+0W7ZT59zw5FQzyy4yM73CrGB6kgpuop2D
UySipJhuUDwSQa7KJgoxQiKAXMNUtEB+lskaLNCHK5pRbFH7Jvd6g6adVCVcxy/9
Uoywuo9bCHjVCBxKDQJYZNUjZGpk3HbPb6C6XVMST1IVGrod5aO+Qj1DvN2XMoS2
Zy8D9Et89/SlaOzSXgFz9HpEQ4Vzd+dOG0FueT576rZW1Y8pqf+XJpjxqK12znlm
3/Ul8H1pt0KKVQexN7Yl+qSdKRTuQy1XCLnbLuphuUa030nwSF7H/5QdXWfilCGl
rPXOg7U0Dm2WkHQdfinOFVD85m96bAhYBEkcHXw7zFN6zKxErBcIU2WJyuTVBwXr
aXbXnZSbfwrL4qw5ytHdf3VCcPoV42wGyZn44g5R8KUqH/KG3i9LSwkyJtun/Nb0
GFlu31cpyhUS51DbmWkjGqPyTYUu60pjV0GVI47ilfeioFI0ikbGySa6AEyucTRG
xdbakdsS8pNDO8IA2mKNVSRDYiVO2sWm+dJ8stQSRaAX+TosiHDNciBEIjWNdn90
nbjw7AARNtJ8TwLVAm4L5gsRIxYqDh3hEHeHUSUDYTP47hgKqbi546yFU3wvGsqv
w1VaMSrcHwKelDEjD7NGLtzXOPS89PqGT0Xw1EjMROxkVclVv25Gr3l2Ap34OKeb
Lf/cFSYY1MlZu9ObsCno636EqEEn5OHE6tg/DJQVFcAqLZDO+fyc1ea1VFP/Z54h
MoWIIR8Eo0MkQLsjG/k0d9AssHFMY0V286hBjj2sMdrcXkVNd98cFVnKd12zPore
hOFstUosONwKnSrp6wtSniGe/UV4qkjuNrUGZCQFZzUQMZFrNiMD1XvYUYWCxjze
HCNBJ6ohxR4LNTEDP+Lf+0zgoe6+4v63s2+FOpn7fZ0TKcFXHsw5+kF3Qe+KqGxL
8sPrNiUcxgwdrhnZJYFk7UhQn/cpxQDhDOXIoKen0IeMyoWjhr9KAH/ITHcvEsq1
y4N7fwP1N5laaDJQFuQ1fnD9yFSXABRZj76v0uQra87JdUi8eJ9OTy/qZU4TD1Aj
eP8AyJk4tJJKmqWN0fZqERH4dKnFt1aFd27SKSjQU4wK+kaTVm87JuUoEXPZcLm5
fYhZYloAG6z+1SkBhT00HAGU/GpM4QJe+PD0fN8LVQ7tymnbCD1Qrw7lICvV0k9c
iF3N5kvmOlW3wvDsWbqRUio7Fzpn4CrJL82x0FpiCvGLhzZFzuIY45sTOyXutpIf
7AB3Tjxp0xOGXFsk6mxQ/exkYbWC/bJxqG2Ro294bDHxLqwkmbsyjKd9W/dQqU4V
uhebtD6NhGYS2RIkYpXb+T9Vg7Wt8z5MVtQlm/xdWWyX9DlQS+O1KyWW8D66kJzT
g1HcdB0nBWZV1PRwWGgS6Fcac3MhDBVoMxEhNbOcoxNkHFUg+aT/7kXpXf7Pq4mL
xhYJvb0qjtQrDHUEENe3Wzj9qqxY1hKDA9dXieK6UVQz13HHIf5hSZFe/8VCmCSL
TV7ZouT4qiz5ZvlYtj1CpXz8TaF8E4cW/U0UgwocktuGQzYkuVEDarJUrCT6BtsF
jHiMqmUX57dgPjFCbbjdMPQT53+56YInvSnwt/xdyw9IJ1wGJyKF583HqbBx8cmj
Srjz+aCRDjvu6ZazGIS+mE5wc+kXOfGCTMQKmTPQRP6LLCKr+C/UrX82S6niKSf5
hu7VBCvZOvM+cXxGpUx+foAskYHxFpj+6mnqLi1q4XYxKpg58Tp0fGjQsTPdHrZc
C9OO4PFypJIWIvZl+ok/o/dC8Sp63zwGWUnD2HsD1WD9UBGDNp3MQBit4Ze/MVcy
I7mF7Zql3LnOznii+LTOc8WFpIDaw/l7Cwm6zaQHz3G41kHjoORGfBKZ9CuVXOuG
vY8bwKVSW7pDn/hBZmf+0Fu2kCQmkxsxATlVlhh8GCdkqWdeXZw7ij4e9HJOkZlN
FlAUcdfN4IAQNfB3bEcTP5a8o5tC0WLQ/f5kRq0dA7oA0gRN/qXkL/XGHr+DzINy
tLVAmqxiIIH/NjxeidPvHx0aw/y5HMpSU3e/TevWI5FGejceWDaSvpZ0iUWNv+OS
t3QO4oUUsp5gGUvrAdxRr6e1/acswTVDiEZTa0EbnDumSxwA4IBZyymkjS4cyNlL
Z0bmcUWj/B5QoYHpme/11VHZdSToNr853rjB9A2nW9hvJi7N+vhfexxH5llP8fJ9
5R9UBjhGQ484t0D7x9tNhTZ8172urvElALBfnPU9SHHh2frvPuEtnW61QWq2uYP3
o66V7sQt9Dwum2CpUVEPW09+V4KEHZcpoPfk7XG37WIbtL8RUFK8jo3x7Fj/dv1e
bXv4OkVvBSQiTq0T4UgFnHLZ7mHKa1L8PHB/HoAX0KR+C3pEkXsUNMzSKWSU09P6
80ocbyHX33TRmQBNMbc4SJa7TnpjQLnvS/yKHcwvIDH8zLYgjXQiDywOhb01zKE0
SQMfB+azCi+xU4/nTo1Q8hGethJgNAmKdSCbz6zSVTkajM6owt1F2njmfzHeKywl
XRea352YFPhlN3Sk0BWE4KW7lXtiHJ8TQjRXksGD5XgJTnt0+XLW5csRbu6KyAGV
3nzr2QAZ1zsk1zsvcYShHhWtIp0ZfAL0EQHeiBy0PZfDRPxVmAarvmfGtOtPwYxJ
SFPaE2kLF27Xv1DxMSiMBgsNPAhDzQP79L/xxTMvkWE5eA7wItvbQNBF4/cupQGM
VuXKr2Ft2gbl8uTu4GADDIconDKGWvpjSMj26Xj6A0l+AWVaQ8HqrkipeIwLMDlX
6/Oz74K9NySMbdaQlrw04cq4337rnEg1ZDgCuiMNirfX+wMsrnGVDFuPEMUj49K4
KBNOBz54HYr4eCLcrQtsGWqOtXFexihPVU6Wdc+tOf47hXM6EqKZkjrmZbbSZFSN
jB76LUMYKhLoQ9QvjCEZW2hm9lrekKm5KtaZ7kw7GMDk+JZD/n1jq5UO+i7xYCCz
ApcHWrN/iIR4V4edBqBMCiXWotqa9R02/Q1d3QP90kcxCZJKgX6fGDYxykcNde/u
ZQOA5j9YV0etUy7FM6TJVV44ZB0mljE+cOxghxmxY+Cmz3SO48z4blF4ScPLtrOl
NtyEmK3QYDfvXJ8DJznwV6MDOfcF5hZ4P8ZsFDmwb/1RgHI6G+uL7Y0ZS0KGBslY
RxUraoPsoncQSTkPc5rSEY8uwP7u/CDkgH0Lwjt2AvkfN1lyATQIqkIpz2VfoEeW
NecGGZPBsqbRRwPYuElS30D8FdSxnQZInsMLKNJOwQb03ecq/Uo5yCSUCdX8qAGC
u5Dr9oF4vIvpfZuBiNW5TDHceFi/sf7wL1Tx9XKHpCn7TE3ulMj4UvZ3PeEtvLYV
a/+0+QKlv0y8becG8Imwywy4NWubNwK5aojvGoLGby1STn9+y0NbAp0cOpo5UYzs
AF4dn5ewQrNq62ar3NxZVAlNsf0/ACmaoedoY9uVuKGQyQ17R+aUg60sKdgRbA0T
bC8xGjT6IW/cI3Vgh+ctZ3UlVObzpNkeg+wK5TKq1iD0aG9DUzaF6ge4n+By2gDY
I3YNGIds/ffHBnIFXjn5uByilvkQ8TqHcuSvSy+Tc8DGDrLGj2Q20OCBoUMTJMWR
mSMKvWBVphXORLXPwizhdKXcUHVZ0YArt8wHNf+JQD+1qY9bmGMGpCrDYLRXhZR5
ZMHJpW/bAFn/0gKwqbPggn1fOukcm+VEGTOj+T+7Zy20QaY6Ih0ghQhrIkizwfXw
bAWx2fiAN1JBOQg3sUz3MmfFEhV3dkcbK4O3SxGQGt85bVjPYfQ4xsEOmrfUNRVQ
QcuC9Wk1cC+vDS6yuK4zAreY2sWo3OCSbv/zvFt+md/V0usZgfPttkWQ0LtI4v7u
Da/Jaqlwfbhh3g7fBhAFKJVjZiNnr2EwrKnnVayPpBcvl5wngW0aF+VPA3xHTQ6q
y3MFN4GuZIB7Dr55Jp+7YEFdqhu/Qe+nM9cTtK55gv/6fYCMjNeP3ePFJFn4zLME
DyfEi/DWyhSXjeaRdqXHVawkisrOSwoWIHKqdnxNu/yv9/EI7NekdJ6jBBEIeKEi
4mJF/HIcup1lapviSYUvZRhftQLDe9bYYzNqw7LVynmb1vCiclF/HvXJvxz4cT7l
O7zD+1rA6dN6tAnxWb4XpeOlfFpMSSgLN9zJL+Wol+70cX31HM7nlz9u1OolJ9eI
AdoT6IKX2QU0PsM5Z+wbGwpZL1+S5QaH6hkJr66SyFVp06uiCGYcEcucJubnJEV1
AyKpbxsOrH3JNGjssfP6wZn+tBq0HZqxCBO9sxGjUX+lyYXk6WSWSEyU1l6ifHd3
f6oiPWLfwtHTziu0rl9YJcSguTzPfuEfnJy2kXueU3z0r/q5Y0i744meVzi5gZjV
xCwnzLghiAtbyAODcsyzCQKyDUrfXbjx66ZWchpmIXgZjEmMspyMObKwaR4F6K0j
lw8L/LoFm0sUSN3iF9SBqyQJoP/Dkhe/QikknLzd6wxS8YeI0PX99ATarbpq7i1C
RBIF7ITOuBphsA9/k6Z+PPVaCiasyJSGhwcfOOeRR9EhlitPU85DzaGgoUyfj1eT
483k/10x4E2VV7N82wa+zcuUA1iCUvkF5ugwJkecWhjiaTF8v4kj6XBOWHSA+I3c
VelY+DLAGNgR44YV4WWww7pM2DJiRqU6ITQTjbsvA1tCdQ18pIUHKu18CiUaVgT1
+Q1dX4Dy+YqlPwPXLou07hq5gAWIJBuu1E0oGa0KbK65ZEFIzJsHRO4JwnbfuCZB
TWSXl5rstJsD/z5DTi1NUHcG87LnfE30QdnoOkvs4r6xDORbttQtkx99OzXI2DY2
5lTfgonlqjCmXnvdiQogyDwrdeUwTLxGWiXh+hEcP5UwAg61zanTaz+vEZaN9god
LycpI4T0PPltLl7wOyKJGdH2mVrAp5Hq9jojeL3FpSpUiDaos8zoOzXMYpouWeTa
k36SlfjAlIH1T5Xx9Vz5mYHiBAPKpcfSGSfsGtUqbchb+gPx9eX4qoG0uOxz3A9p
BM3H+gjLdqtwSdO0MgsbukCGaPAcd6ONsl7ETThPFpxhnoyIdTiCd6RRgsyNQ+67
RUSKNUxmH2Vi5af4TdJdYBiHHLi5EAO12HjoRyhkiAH/QpXs/uG13ht17w4gFqoq
dGb6yrlMfTaUGSfV7HVMhau/hb0ejJJh/NJ1DpJUG26dOrZnbmc6OTjrOYI/vz2p
rSVNnpmDsvrIgnxugGvN3zr9dOq5Ont2PNw/kMwifi6TZ9hD2yduzkAB/gWbaRtb
r7lNZohB60XFyA2kURjIutkYT3m9SaMSLh3U+1o8MhcxVdJc3EF8+4mNCPdT4W09
tnY3HQathdYvj43/KmObugiz0ZFJJ+ajidbhTjCnhbqKhqLlPlLVsQp8dypoaiOs
zOfITrNgx6U5j2jaPvN1yUNq+3PVbQ7u13RXVwsJqKy6ftxH+PP0XnYv21ukos4V
Zd62zCXWeBzLB85ZT8cvstUwYToJT6UKvPucVi7M49GIJPZbOnXoF6C2yb8r4yGJ
kqb4SnMfv5oPhC5ulEQtokKwirA5vPttMy0rUcvTToC/fPiDD5QUjSYaG/7IX2GJ
UZPaEAjPm+JUAxGP5wJKMM/mUP/G2Cabl0gxlY/1dgt6IEw5CmsN0lDaso3aTZyk
w1In97+QL63QyjmMc/0fqwYOG//JPnu7vQiGikcDsdckKz86hYVKYiHvwRb2nm5M
BadJqFP0PYXiV8OUDM56GLqQ/Yu0jejhXoDuqLzXCSNiD2BchBCLRbk3eWZud8xg
Jdvx1n/PG50cQMFP/L8l1+Z6Zh+20ULnZ+JqQiJK2xYJfxdDAE1eOB+AJNsshagy
skwsZ7wIPOhzckggI8xgHl7uo3pF9WQuJDDVujELeCXHJX6MVpK5TKSdyDGWOB0h
8HeZzBZ6TTA+1TFPBsym8uMTetoEqO4KFP7x9mbOQoLSoZt1hudxsJbbgl0ZM7gT
6Yeo2YLS9oyPmjecbC9FSZwpvRkHqAVS9QNWkI4iW7J+5jVuiREphF2ZOeEPXoxU
MVMAj10bLPeTUdsJSH61eUNuvAvHXI5AUVGoIRRpcRzHQiMyQjWEl7hbTYeLtOL5
Su9SiPArMuSMbygSliMT/G1VonHEsLygXvgbH+pj+zKPIvLBe4VrqjKLxAPNURNu
hlDr/vnVxO+2EtRgcAj8gwZw/IP8veYfllTgUx0v8cyWYHRLGZzwfg2MWEzbgD0A
SQOf+6eBL4tbiKatcKEzH4PsjuL6umo3psW2E6lRFN0EIJJyFNtRZxVcnO+Wabqc
q5lMx/ZFNBLcQIbaNyaTGKEaJyLNdhLwLdEseGxt5sx0KiI1nPXPowsEIYGKDBPH
jNouugUs5x1G//46Eu26inOK91k3NH0hUuW8fGLuBGYxG1HyOiAZuqjDo+boSprs
LacF4arr0kEtrX5SXrgUauDfh+oIPbTuLsyRC4SU2CBI8pnkA/FbUuc10RAoCiz9
nHx0U25OaeX+EGWDVf0UpLMc6AoMc2W4n8bWe25bKy3ov6jjIosrvk7EFptB2iST
+KSHsQ54ruzbaMjeBPZACYa6Yqqw1Gf7X8JZgR0gz0/Sz6FmaLBJGd13O1I7Q/XL
8oIThlPoPMYps7cvhfRlFEXLKWSfLXzCpq3sRq1qZYyjBJNEWCcEE18MbnxPsT8c
LtqECXtxPabHrdNSlQnrf/bs5uqmPWfXn1NNMKigR8i+6jnCTHe8YkG7gI0yhZyT
cTqnbo1k8atRThQJmCpjns7LIcj/R1UZa6U7oKEgySoAEnbZBNkZsnSKDjui4DcN
YAy0Pob2CoBKm40Ny+ODDTmvBGbmdlbBm9zBzuVmW7jXh1ybs330Xv+Tach7b+AY
bkcx1NMq4RZXDFxUaVso+d9wzdkEDDP18kHJ5agm7dr4EEYdOwHFWqSXDI/jbEST
Ee3Y3pq2gp3LjxVzBZd6uUwztrWok/WSKJtBloK/l+euCf4P3cvEBfKDd3lVtnzO
HB5kZkttK0xmIz+kRoI7738JIJDeolePoscXDtNfpK+xk58wzl8lsilYlkw1l553
36Lzj4LQASe38IQTDDCSmzTxnR8uUOLA/phFYluKSyUS2H/6sU81vZgIygJQv5rV
t5y5Sg7JgFhCeM7EkBPg+GNO4ynnfAdznRDR9vCZh5hay4WYGeidKj9vUHYNob+c
TIgQYmu1iCu/TJHMF65hrGYoue4WY251vj1kSXg59jlfnBw0nMJVLAkiQZiozNVe
FnO+AfmOG2vPWTyBrlJzh/QSBSeXUvnwKerjdmggsF0pxXlnjDaXNwHyd4j2zTTi
r4cLeZ+0f4So+oMPkVFdgzqR5C6rfkCu34DYjdUr8wVJQ2l24LmB8wlTUajkqGPO
SoWSzKFPLhyvBfAm80dLdr5LxlY0hZjL6CM8gW2NoFNkfDp8CMyICEkRDH/5WzRa
7QU1CBGAIc5pouHIOv1Q4/dYW5wsBAccMMh7LPhn3tIrhgxmOxn22WrJd0eTJV6l
DsmzASr1IcrQGSsrRaLy9IZYeuny7nDFnAluIieVBiAmgbplnZS0cR0IF5whn0Jw
5BW8xHlAfXgR9HDBNUDn9NsQavLzlsFfRjFVJEqUryj+qEkxgNjOSplJfSnESa/9
Tv+1O2n/umu2OPPpFAKpjZNw6YkbPd+KiX8EMH2xCK4cbeRtbP1SjXQ9+znt5zHG
1mq2aAZ0sD3ioBNE6xoi8r+kzzF7JTnscs8+atQkGKLvyD7WvKKpymYJh9CElVys
yppPfmwP0tX5ZyB2xRBjLdC0lbGuquG0uf2pdoPhMit4SK3BqJNC0REZ6vnJBJml
QPS4ub7LVtU9F19iKrJJxOsIyQyj2o8PaIZflFPzmKF638TqHJdqeWZM5tJbnoxb
Inkygaf7mJyjIuXJBWfKhdNzvT3Bj+5wwoycEWa6U0ivLnbJMndrlA5UfYYeMXnH
ocgUY+XW/yFMYdKqLLySwgaDWva9ydBZpxn17jmzJBQdwdZT/KcsxOMZZqKYvIrd
PrYrSWt0bZxHVsxIKdy/MUhQHovcCRKPsyLfSVfeiZhLbQxRz/Qh4aTtDPk3DqD0
9yC+NgmdQpbQrjwbyDoen7xj3xrqWPsO7ls76RB+dyDVsq5AuT7N/de+DrFE8IO3
KgPQV2ug3hYZeS3Ew35YzUosbZzKCP3s+e8xwjtMf1gplihidmzdePRXeINcnryy
+JwjrRsYZV9gy3tzqHVrfrWYgQ5MGikgrFAFX1LaM/BZ11QMDEE5DinZyp0ILe/K
vLYoOVyjNwdxD1EiT8IJoMCZzlUf8WwJ2ghf3DJ8wMnR4D+HlBLvXy52y6GqbWNK
t6QflrDETiyG2/MtvI1HQzAZ+Hjtsw1hwIOVchLZMVJ7iE89HqLsS0vOVOLdGb3n
mqP9IP5EWohrNhEjJl7lcvVnNSStXN7Ucn6A0Vy8k0k/QcB3wcNI0ykLpDBZbchc
npKK4dyEAPBBL+S4Xke356fbNyxyua1LK7k8NIM6yPjTvGbKLjy8Ib1/IJdA1A2K
qMs3KUo3c3WMRI94DdYNbuFM0PkvAeCt+ifQrLMhpEY6OHd0FqbrhGhJe8ncIDGW
k/afLP6UuyPZbIbgynAe+nw5vs2jVKlRBbxn9Qj6C8cWayaf2GDHra2zYvXAkXer
WHB4PKjmYzK87hvBequsykCvhRtDMgPRfPDw4+W18VYPcxzS3v21FY90SHuoC657
OSoBn4vex2tL1UfKJsUTQYxQZEA92OIl8Bb5LEPSj58Blvrz1XAYxpPaK1YxDY6o
VycMjhvx1iXWUC5dNIDnGQqfLHV57rIwdF7huZJwti7FKPEaf1+9tUI35XZEHt69
Dt/8iD+Vlo75X7tVjn51hrEag9e3wOT8uEfwNWpk3+bOCa8dfIWldkf1jWgipjfo
49YstNqKeNa/wgdOSHffdG5OViYL12/+WLGAH+3ncQv/oZIL+79QQsJsenapdWjH
v4+uWEdPuqrmsB+hhs08xxd3jMq1gUudkQEe4NYH5G5/vXHyHby2atod9oMNgj4C
/v0ufmUiS0sPYjv2ZlkDb76GYmoK6QbS3TUabhcCTxE4v1y8lBlxcKUh7TtBxbnB
i3kVmZjtwOR+nFCrITVRPs9LPmYn+OMIiWsMh3hXocqin8pUlJrVA600gQVqvnZh
QKthL++Rojrq2v4yNFVcwiKW4jgpCSJWlcx20fHgysXkvPXGj+yCgRxRN0JTcPeg
ZyPn+qj8CqmB2rAGGLHzLR8VMbhEeTa7YJRlPywvkl//5azvvUkH7K9oSit9Nv5c
FdwcrmZGYlEa8fHAV9fsrKwQjuhFufteG1SuDF+lMZo698adO+dt7C7mYHVYvWCm
9w4wzU7qpWgAr1CFHG8xTWgXJ9dCi1Yg62GY1VpAIWZWrX1eGt9VcqIEVrIKQqUo
k29SShnIoN1TXJlX63cxZVa3BzqeXFN77BG3IJr4tmar17SUc3NfOZfngYMZtfFy
LKLdvZYF+Y4iAluLkp/MdHzAKv+1Hxt+fjsi11ga3T//p+Mjrv46JKl7fZJNciQx
9VAtuCk3nVVMJt6hVk4VHweH9C3RXFfj7DOEYtRJwaD4fG9CwkaLut4j9PFfPx+F
89brQy9Bnbh9T1sRHGFoTbR9L5+1xSWY4li+RS9duArtrX3dfTT4xnOjAh8Kwyw2
SOmmgOEzTjPQFUEieMpKCMFwsFzCcF+mCx3oZICJnnIRIVQKn18tIbFbDu7B9HC6
py2ivC56TwvQafDjnb587KmjESj3irpI0A7tfcreudbalPBBQcenGExxNvO7vWem
5iFrL5lj7W4Tk96ILREQgTlkQzuq3+BZYW2v7PSU0X3iAYFqbpM3o01BZs0uoedb
tr3MJEUunNU6c/TZ6Fg/tv1VCOju/GEKd6YTroFf9eRYeubJEEAXxTRFOpsLHI5k
iKSP7uDROJvkLWvxPzVdq0YczBjhaXfVGPvZw9NCUOivzz3zW7+d9zwXxy5kp+oT
miIYhn4oCWIXxXWE1u3E/0bJc4er9/3Qx1DELlBy12H8NnGa70Lt/XUYXoJ+w1LY
wD7TGPi5Y+39FYuGK4/QWfY9CGs45yjt1IOckBa2PVBGe2zB2zYqz4B2hdtUH+wM
wONJ4V2v3QBmJCVLZFcccTK8nE6a2xqWMCoYRUhyeVdBhYKeNuGqz2bst2Jrz0dT
p4S2CG05vcxeUQNYVIHnFOi9L8Lr99+nLj72Bleiu5HNsDkkD6Jv/g09CfjFcsRz
PAHTmImP+THqf6hh0iZ9rPEfjIR2IXcTZBQWJ1xvwHYcmy2Age0wjH8c7Rf3QW13
BizDQCy/0fgHZMpwWOs49V/Gj5mG9FE1igeADCrz4D+ZpeY/xWEy5MZJtVHdC9jq
idwhW0kbr+rs0XWMNwR6WfcnuFm61bXMOc8/sUwkPAScEbn4sK3YBu7SE5KEJ+J7
cCkmAeqZ/iCBn/lm8PlS7a/PP3Pi2MhD3YIuGo/m6aAVWT226Y+tfIyjbYI7di/G
95v+QIopk+k/v+4ABpnIxlTTHfR0q8VHgZR4Vyp7jBP8IIytU+0Qoa6AVQt9Pavz
6GIIvct8qfcU3qxGQShFGBzOVAcr3M29iQKJGjWYoEPk5oJns7qUP0KNS6hCUVkY
IFadHp8JigXMul2vdmRkZZz2TyxRpHZIzlztmIFIasB+vDA0SByzDdwzvTKzDA5I
+fGkYOfUn4FN2ImjYYLY1b6ygkX5xIZBXr7QzpMcjBedJ7QIJheKfQ4uXWwX+mDS
OKsrUmK+N2obaeYS6EFkpBQFFbESBCSWjU1CdiaM4LaarjEJgKXSW1WBXba32JP0
cZSC7akBUOGXTaiQ3OWthSwWSXF6zgb2ZxpXDrrdhDHU/hCxK6uoeWyKlU0NC88T
mcsSgYyF8hZiBjbctkrL7vZyF+EMhZrhJ8YS32/qBhKnVeKaMnHI+vfgoOeH23Nh
jlnusEJS4KDab3B8Jn5jhpygTbWijf50hHoHwStl1Z+uLLfMfIK00wnmvIIro3GV
uKe9P1ew+RHM2Qonsu/pbxJdd77eXaMryIuTrOMQDSXar+SZUOglAikptr5GBU9N
dxtC9V0UyC29gVL8fc7VaG1gn+PS3hGi2udX9T66VpfkcVuQnaLNMVl0qmqQUg3q
Spl4iEFKg8HgXr5F2GcsWADe43UGXCvn02OemFKAC29ZIkxxtRZDgw2+Li6zKzTv
b0mxylPfH4aINuy7VDtXBtcgDNFPchN0pDut4wkdQZWWoK2D1MS+VEbo7Q0RU1O0
k5nZXW9QjDN9LXS9XcaELyP6icgrRTsy/ZlIzG1weMcoQ7cAkY6sqUYXj24TK+3W
Ro7FuhUvny7lf3XdMmFXSB9z4u3+TsZRluKgC31c0T3ZMdzWqMJGk+bdSaK34dhd
+o+td8pXus/G+OXGwUSvbYLezeoP++R7poFEKuzQu/LlZyVTgAZcgNIwJeYsoP5v
RTd+Xewhuf8AtObBV9phmUgOQmU/3bpP8lpI6AII9gIO2WSxpk0Ej0jcAjDe+QaE
TvlxXiiNi0USa+h4YJp1fvOuxECnfrdltgv42PoGCa29rqdXCCo+CvLPZwk4yADc
D3JFM2P5kDJoI3NNg4h7XgHGEtrQywZSrqTvmrMYUeBoQhYkvseR4R1pL4z+zHFG
z9QCVnZLjroarKxX/GjMieW4qJCE4Pi2kVr7kpsx4qVjFAz/2YTRPkqikQ/n/qZb
QDCMNscKvig5rAxfZi8rmDqg9XF/+Xp5ewwmgC5ATVHkXiCtW39Vfml0Wrm4b7K+
11ovXhY6WECrkVvLHvie87svf08JnsIaSU9XzwTAwR+xmqzwds8UWa1VXnlTKRyC
Azax7li+dB/ASYJPccYL2tCibqecDP/IHmekP4F3iF17X0LfLYDIH3S7vMX+s32o
gXDbkuSEdExYrbSVeM6r7ql0xm9kKZphRavqzyJKSL0EGoS3LYmK2oH6lk08j1Jy
JElMhBBCCK5odQ0fn5GtkH6YiMTZTTnYZXNyaYeFumBYn+4Mjm4eAdlzu5Ye6voc
qNBhkc4SDqCBnQNGDiVIMJcJ/rzARmePvAz0V64/RdCiV1vrIp4eGsmxu/jhpYS8
8xIgFwwNfUpzNA4wuxIRNXePT02MQw65rvfKOUKv8sQOhY7PB/HheVaETq+4Ca66
pP5tA6+dEbrK2i5qI1djMgOCihx/8Z5PclDLmhIQfM3UT8ynloGdCNxfv/FFKXik
FEV/Ah0WVHD9XLKin2JaMCW8cZvo047jiM4bmuQ1S6kgwP6VUJatAwSjaLkV1DPE
1HGUZtzLkm2Tvn0IeHmK0CH+EHCcVjwPI8/u6uDJuKnkaOYgdrMUfwyDd78evW11
R4KGZtqRZXiUttHSaTfUYpKaHonfON4ElYmVftYdLP1h/EKJvzMdRDNs1e+Y2Xe6
g7Ixi2YmWH6yYEd4PrUCn28rdtbLeMvYyDCewPsnx00SPAl2wqleVRnclttYShor
sUXdkpxsRHXNiOc3SWC73CEQswgAg5pKEFis+gnYxlIkwE5zZm9B7OA/o06hPlC5
ki4IK+/9oo3xa2LaScUW6gbn6hDFCRibfbzTYu6SJr7/N/IfhWbfdzfb3V1CwUgV
BN7uPWRAMoJ0+QFNd9mELxH/AdQknZQ9kwrJV4hzjis3lX8b3nBntG3omle5gwew
SQqfEAEdPgPBJzwv0SVCDLAcilfhkacxTVCQRYbJ8z+qne0hIq9DcV5nz+j3Vt17
W9eJ+kH93/1X467h93ihPQNVuDS6Z4qDY7M5DMfhYs2L0rt8LZCUMS9viPZ8Qw9P
XmK2rdM75IKdMHC2VoJ75PQqYL1B3Eji6MEGiBXxXkb5mBGObQJDujPI9DXqh8Jo
hKAlCOu+XoIA2mFAvRflYNkAzpFYtg7tt4BVpksRuVuG69FdmVVSbPObRrNEQtYX
Gp1n82MkKom74vMF67XUT/Rn5GlQw+BaG4MOeCDu1xFU9z/7vTCpjnw2Bgmqh/yO
BhvmB9mqfo4ztXp3/LNVutwTkGzyGp7Qdpry42UJ+Y7sAewEzF3jSeRpWpPSXjxL
chOO2lemBfj85OUZ0tdarAf0IY4rA/nGM61dYgawG6YEdbLhdJ3So7EZGb0ZQmAR
iD2K1dbeuAcull7WhvPTbtJpCWhkI19H4jpPGHN3c99gXnpCTXosC8Hm0oljzi+A
xT9MWeXomHQKZulpa/Pw9d9MXOGIbsMPYB1n5cP2on+XttsXiyWRHDk05rnG/XPV
2uz/HgB03xx8Qe1oyGrJ/nFu6fRL5o+n8b8FLUaA63nDwueQSIVmePYMJatmnkKI
Sh03bZywMahk04VS/lc+Xet50s5j+p1/M9z+bhkpYOBfJXCXJiNy2G58QV623Jl8
+CwCYcou7G4oOuc8JIaSaMCh+e9nXJGARaT9+0uHx0q99fg/I8ckwozBRHyu+lBD
uu3V8/Nqj8xE5nKaeGPzrKx16L7Awyir3JIN1WSr5x/ZPeLj9DzH6tSbWIXABez6
ktiwia6nyKNaQbyt1m6Zue/rz7VZPkUDzj5IWnmZu6CbhWk4LRxEyKzOFUm0zk++
oNFXnSRpd86vOS89bhybcBOP6fsaYczUT8ws5Qoo+D/Vn+wmZeU9twA/F9WPU8x5
v6On6y6E3NhOrr7MZRss+Gt/XJADKKe6QdpT0Hq28rOjjFJJb4p/uQnxRblG0Fx2
BvpfYwW0JVVJ3RPTq8gZWd/XjdaZKXcPkAIZBgTa2FYF4+oaSajnGNHGaTQGvNro
LaUT3NfxMbjH/cAR+1Dn7ZSzM5QQTFHQv49tZECQa/McCGfXuj06gf0zV0lydVEU
qdD8I9IfpifYiffbdOhebfkBR0+2hqUVDA5ywlXG0tvKyZHddyaFLHTO+018J8mH
NicSKieq/LRc5HMGjbPZOnLho7Lg66mfYNVXOGREzRpf8nMFk9UopZU59Kalu0uN
e7vnSttG3nXj3gS542tGCcfW+9PBHdt2Hg0B4YLVmCMeKk17Y/34R9JTDqY9EaKQ
3h9E+QMTso3lYlqGzM7Q/AOos+YiGcOQZ3wCzJ7ki8TS8PIv+Q6SUW4yKs6pQk2o
94U1tn7ToJiaQA9oGwiUOKMGC9bjs7uP/M9ABUfCG1Lyh3GAGlcR3vG1k+gPHLNJ
/y05NqY75PzWtVpPcnn6RssU1tROysWgeCksiVIctSe0z5iBQtnn53P5EL1M96kc
GoR7c2gdWbc8379EoZsMLF2hM98byj+c3uI9Ejhx20U4JIuQywtt3mtzBu7Ity0k
YFohhpDIaDCMJEsQJ7Kq15WsexwRQP3psW8zM94brJe1lN1/bpOofUbPFV/b3Xla
AX0KJsaGE1c3NnQWvIHawTGYNWRzjLVOzgcoEZQyRYK82UOT+/VE5MSR1/bMHUPH
K9dbZCzYaQSkEpf7NrBxsTW/REeX2CIFHiZWaowbNZb5enJGegvrODToiT/7IV85
z2+FfBPsbAdDBS2PvnS4Syy5jBF1/4tfAwcO+2i1cZVz3O/Kkpsbv7T2YMfTX8Lg
BsaLzO+6B46IDnzT9eVEEbN4cUs5Z2OopOSdQXIKPakjtAR9KjYk8oWr37GKYNKX
sIUsAsnfWxH8h9j28YW8yYk6RAaKy92/kf3uLoqTBGI0R+9NMED2LP0MpJ/3+7E/
nIPQMGr9bK+n3IfFiMzMloBAlOsjd3vTH8ZSkR30nviRi/0+J96bQDj6Cluz78l2
H/NBoFtWQwb2lyzAdJeKG8aZ8qTfJrGtaM2DtejFG5I+e+XCKYjrMx82IGV9WSP5
cpOP20l+B1/uKJgEkLrDsffGmB1uChLBYldnVq9a768Rw5ARuxk/td/lzYG9tY9T
Prh5KFOF2LiWE33O/hveFhPaAe/jclQMMNxnpQCO3vW/dAf0vqkqrcV/Ch7jR3/L
pag6eqRjdzKm7IIiZwrR4v9yLNSlEUhOJjJY7n/m4eaW5LO1pJ2l7nRG+QcywrBu
2iZqVRx736AlQklw6TjbBhptGnJa/R+zxV68bRnEbTT0QhcnWW0axqiB9DgfohCs
AG2EETeIlv3dQzb9xpLzT/yyoyswTppRR8BPGxvYDh2IGlDtHfhddVYDH2GTQ1ad
bJf7OH9FQJ/unCocohF1+h3oadc6pwgERZ1ksgK7NOdjBC3B6DKBfJI1jqz5vefB
D9bl0TJgCCwRvr3/gcQPeNPsCU09QIRQgcrpMjefpT15Yswgq4dd78CB9c/apmi7
IigBtMzmFvCkudOnmuFgZTjtvyuRBWc6JsSEwMabkU+uABWegammxoLcGqFHlMiE
56Mb4L4ZRaHJr8PUKimUjbL0atpW+zimMLp8sIz/1l6TO6JSiQChFFbZvicu0yYF
E74nVnUEH6Zcre+D1Jw9A6I1uf4TGYdf8AZ7pH7fX81LdpziK8i3fYcY1F6UDRXK
aA12OzJ0NHnpwgMiHjKjFgzvnivRiGYGa1TS7jTMQJkHb2yD/22JLPTTlZuZxq0z
4Zo7BWMzJbGyikq89Bc1lXZRAmrzS7EVy7y9sgDEKug6lBfhqmQZMg76Z6AIWasc
1QG9TLpuYb4WrTsYtBHRS9lj5voGhYGW0Gbs0pUTx4mfg2uUymEZeSG/eOyTAxln
3v/TxpRSkkt2Dk/er47rlKKz4+enwEajIDDyfC61i0bZCw+VqHbXKmYjcrrBVqN+
8i62+DuUJE9RBDO3EVQciIVnsldssuEK4DHJGEQFCqAAxvh/i+XB3Dv37b0HaZmS
KLlhsEEvFUYXAdXYBGX5ciz8pDV4pF5SKYgK4laN4jL68Py6KM9zDA9xfDTiibXt
1/eWFW2vCCuAwhuGpEEzzsSUZNjTlYgQXTfjQVxFuJ507UqEb8+vttKk/ww1Z2VD
AOdahDKewHfuqm0P6Bd4M5f/zxC8DHEbTH3SXPnQYXA3X25ApuYVsx2seuLEKt+6
MQDbCF9Vpm2hSRUQ8nxJuZ7KER/U8hFkOro4gbQOpyhMYiit4EuEQOCAjlLYtCW5
p7jnwzJSQy8HjnqcbAk5uv7Ti4hhm7s5/AN3cqo1E2cwYXuBKpx5AwS8ENbxbIg2
S6vsNlkuMrTc3ipUA2n7AuifsbGsMHh/U6MBkdd9NpqVmgsKXhiMtRqB+zqxet5n
XzDwu3TadWMe13efECdc9UzgG9yNq3M3Zn8mGmzBn3TtzMAY1PsKx9SAUqYa3QDf
4Eofx0eBFM4EhuuL+gk/oRmtgwzdl/k0ANb5XgDxfa7xOfRFWipBXXUHpw1pjXcS
Zq2v8YtoY3rGm9ayI8k2tWV+kdt80CpydZMrTvQLN0fZq1twe5X1NJKgQ3Pflsj7
JGP7efo1/manlFN3mqLGRSsdYVWGpl7XyN8BtckNqa7dMWvqfkz6sxCDXLix+uCL
Ex7/DjkwJptTLtUdS8OCeCSRzrQ6H2RygbcJQKoyynhlTf1lc87LjtUdh2/LqaaI
Ad6bgoxncuipWpQzPqje3/vFPmnfIDk2Pljh7kKEVRm88JuCIsvqfQn7IvGwMHMr
VvUiqPtg0Jp5a7yXHbngKN9+pztKRvuGiAmU75pasRt2OeOXNUqB1NK+U+pXLx4m
QiCz1LZD5DWKS+NJlMzOuoFEy+EMLHVWB/QfqujadMzkKIi0CpWm+qUBIt6HgxjO
RiKcsK367uouBBgLI2iK5C0xSiWho2NokpLTXCM5wnJUAVrxdorrest+EOaUlyO5
IYYr5MExKrs7QkpJ30TUymRWEl7Qecwaap7mmnHAsFiFa3xJqPiKBHJxG8Cjj8p0
oq8lbB7qiI1I+RkSjOKngkqr2md/oHlhJ9TRRmD/pt6CZOYydSLOfsglMfKxkgax
uHYbSke+qUtF5fLDUoWOuD81TI5yprisFqF7Q00FEUuxoDLgSsry4SvGHHX/+ZBm
5Lmf/rlHqAyG3uFxHNHA4vAdyKfTMONrv4hoR7/ohTMW7A1wuNHL5du7eOWR+HTK
sw/SOSc7cvA2xOhMChSBJKGkSi53a7hgGP9SllI9LiGT9Iqnx7USp9QsH6+W+4NZ
t6YzVTpzhxpI99he/4LVCX+uyqdaLo+03FUKCRp1W5P4KyUS42mRHywNM6UTaq8B
RKfdPbudW49oYdyKbRoMq2YxCqZ40sJq5n519/STV6v/7imzA0kB6xvRsIhYqAWS
zkOphSXf2//IejDHXeQNw3hOK1bdCvWWq8vkVG4EWrVgbAhdAwD0qXgJkyD4JRmT
+bWugBNig+WcVIYrWz+yR/oi3WvsfW+ng+XEyJ9YvcG66yBlSRfDLvVOhP2kQzFu
nZ5XW+uw+dHqmt8T4pVLgcL94h1ngz8EAmy+RNYu+jQVRWrE+jmOIQzR9ReaMuk3
pd5Z4Is1jn+ClyAVhs9ds2KiyBMeoU2XKUMyE9YHkM4QyrPJUsjd1gqXUtFSyv4V
A5Q5lfACD8ZylgInN4qI9SROQYW1N+eeDccTld5p27EjxwkJe836n9NgaiNcYFYE
7DOQ5X/w0VrylroCP0cV81cFNW9Vk/HjaynuvNvBxshMAMebhNBguXM+td8mv050
ZDDku9eFHLiGDDZM3+sL6dplOAXC+iDs+ItvOz8c4pDECGgiJ4EJecDeDocjQBEX
HhedZ3xNmpWkHYQA6KIMfw1lRDC+sT3Mp2EuOmgKcDYiEDELmvt5henKHEG30TR0
WuhIG9qZFjRv+ce4rpSNk2oxgASwVu8mvS76yjBIoQH/awUkGwu0K6HvXxM52A3I
84KlW1eDjOHG4ae8lGUxvNQbanIPeIKkCXjwKuwELZ2N4bNhWjR0GLcGiKlWyQnS
l1T/lGu8Mlj4NE17IoCQzQfU8pnfKbjpGqf+v0+8E9bhI9W+LoaGUvRp08jIS/mJ
JvSu+QMCP/y7gI+qf1V8jFJIVDriTgfGrzA7IvLRCyh3TALhZKC5pr+Etz12/sqd
YVEpcGBLDDJuK8lBH5I8jG1hTuyIh24OFPTCsdsB74Gmf9szvd0EbA+uP//s+f+J
DzEy1Gsk+pVLsdg+U5jq+ubhzoO0vSfGM/FzMmGYWE3NbXFs9bi5N7oEZrW1565a
uzsw2FyKOc40kawuuSzJ14hpDedls5OdsT8DOJhweJ3gvMeCdJ3+rtHrWvB0L4J9
ohgVvfugpVchWAHbIe+fGLqiZI0Xdzwm0AMw1XVoYqJNWmTjr8+MZFcCbeq5gveP
sK+FoYF4kDL/Mn9t0b0M2PmK0/rdesP5vsTB5YxlF5o4PGfe8np3vw6XjGpsBj+t
hRuJmM1BK900+0ZK5MHac+n+Ka/83Q6hr4ar6Mg3lKj176Rqoe/LyD25h750SrYQ
PizyN7oxxu18cBxRbfYQ6pnY706ThXeq83TvTZYSHy6c9nrVKp5sv2bFWuDTuheI
ZUkYZZagUJvm9py20n8PE6TdqEMB2c1CwdsoSlVORX8SoHaeS/XYFPvva7Juuodo
hSkkvFB6tXpUUlcMI2+9h+Bw7vcN8vMJ5qWHNJi9pfYXF4FrB2NW49VCeb6pMQYL
EBl6p88yow4VXLFoUy4Tr/P8R2jkPzJbakelkr8ZBYQZ3nFVQJWS4eZPxl1NASrj
+I8yRq5HrWM/QpPuupE6dpEZkrj2N8Xc+n2XYpGiNsXPYK4p0Sa2iOSC5lmLuFdI
8H0jUsChzLQTVyIdCCkA9nwLzKdASAF6gadKJdWF7wRWUhZD0DJ+bOoZQ8Oeizft
raZVpA7LjnfKb47V1y30aSLTm2imkIuxuKIhegAlIVET8XAur3S23VS+dE+lwnPj
Eb1bmiDyM+rL0xVO3pKluEuub9OJlAYbQ3t7VFfD7VxBxZ94u71n4sc8bnqRu0N3
i8x1hz0b6E/FmNocz3ybdGAC1n/+gQBliKfzS7dF98VbCYfqMybC8ZgGz9642DLS
cy2UMZymix9NI1BIGtTjmhP/CovDaqONhW4Jyzr+iYO8yOZ6YaipsbhnNSIQClXt
JO/l/O/KLNJY786vUc6toxmBQa7/YLIgqvSTbatVAmwE0yDk7urvMh1xmhe5HKcJ
0XPqVd0oOPDq/t02P0as2tJXnO+6zaTcp2VkgFk1wn7+hlIP+nhFyPSdkyJuOG47
Yqr3ybU2vHy9kB5yK91zTlvk3Hvkg4ENk5QayFFL5CI+8JtDPnPolGFb2nXEv6iz
OB7vR/06nOMoEl+ADPA6tBvxQpUMxDxT55tHjvGz9I4YY7T3CdOW6unvULvbZxiU
ndOsnbn9Z6C1Vqi07/MfkPWHHo76vldWt8tmsXZcnVHUOMJbRAi+b5ZgfAFHto4C
z1zL2smiIgW3t1cflPKsue0M9O1+3B+Yf5VG+dM0QSpO38uliA6aigmqOaINSqtg
BsWtTaUZFvbDBWVDvXdRiwFqqbwOMkJw+7U8dPk146zWbjFcjuNdvY/G+EWQ3D8M
mExgLuE9B30joMecTA1z+93Ijox5dqLlVASrRAR168x6D76FfCnQWN72NWoa923Q
J8KnGyfGuQvnMu5LGrZZVizsGMAtcg4saf8VkZIWVKcvh++84vXOni+4Apibn594
DpNzFSPruKVcMFSiVSBu9szEFycwNTooYCxBnSxdYY38fsAYqj4ly0dPdQwtjrRM
FcQtWTnBoAMd2k+cL91yahIauLWPJnK8UmhmYG5t6+MFQKsRqJvdiKAg7if0I6Hv
1st0IpjfuUjXG0V91VlpBvMj+edVIrqc2slYwEzs1odBksSsUX6DBHxZzJ7Tjhf1
0ago6krCmlue9yKhmGU1wUNSrjXU83Yl+9uMUJErrm4RMeUzt3fkaCaqnkTkRZQQ
36N+AC0llN6xjX6Roj09vdH3iSY00mXjEMAM0HX4ZbCjK1r5/ptaGArE2qlda+JP
x2SIkUB/+10qO1KS/OYsy8eqpmk2EW+C2UlGpxOnLUIl9+fl3fMITMlJpC6XetaC
u2ghinmndQ09mCbSGtbu+/hpakz6X4lw+bl7hJWbhMztU9xZQEgAFCNA4NKQ6+rj
6D52Aa4Mx2FnxlB/C0qt3PtJwfdoGOel7a/ryi3n2YLp3BQk4inIaEhtehK631yS
jfyPlbY/WJqJOu5fyvEOCnsuK3LwtT8TwEymR3uVbHdJ06/J13Ih3aUkSs4p6YgD
s2As1PC1EkyTTxE3muGk44+PclZnipXq95VDNAWPzknLl/1Ab4fEuKiRJco3RNUV
luB4dyDUP4XQ5TgwRnedfmiSqwP5DCYxlUJayHIeFVr6bHaV5gVfEnzEp8/XRQQk
iXC36+k80/QOiF6YsKUZEYVd6qXhrb8311YEEmD/E3IBvaEofTkk4/g7ItvOMErS
TZTyG95ZTfBd4EIbWLld9l17Ln1KEFhZHEQlXrGT7+Q5Jzk594PhxE7LbZF5OSSi
nsuLraMd2uwQtU0XBUzfoqLys2k4WR1VoisxhOcvLtXSzAx7GKr42zjYU8W87Gm9
AeoPdoAr+alSi6O6bgNFTAcYhEEm/HdKjeAbqrUdq+KFjiulVy+O5U8mUCRCwt+q
p5cHPb5DC4mkbfXEm7Y6R0f5YjbC29GvDKIl3CenoesGmwchAx+3ZjDAejQ0mPCx
uZSttrDjUx8jKZNPqY7nfRkSY/pI4j994VBttEZYN0MfAYZI6IVpHbjtBHsDa9he
+Yna0IqE/Hr4EfXMcvpHed4IvD8e4XSRM4slZ9+eA6QoLH2FU9xqItO+p2IFnUsj
8XwC3JBW/vFG6T9ylpXQ7lz96iCxk762fz9tnew0KYOaJmUfREkMFCRRzCJfyxUu
7+QFIJpe5LIYPpNRUgu6+Ozf2Ogd+h0kTl4O25E21wJMVbMnU9zW9q++5TV14Jnq
892cKnOj2i6fu5gjzOguQUToj9kxPq6cUSwj2nnspayTCcbULEeq/a4t5J8fZM69
K9fhF2WpYNZO0pohupy2GWX6gVgMWGQ4S87T3J4YxxD29aRZO48geOZxzYEw+rxz
IDL2mYp+toKqCZr+MJSwTA0QDEUqOhDsPgowrfDIN6m3i8LvUn5uulkRYZDcCTrZ
+O49O7+jtXLNeP+4+8p/qCC5w0xjAYnCCmqEpKzaKe3tic2V+Lg7grWJ4hq3Pmud
g+KVNX6hoZ0bn8TJzB/+MXhPgLIrHkix0H9RWZxfbbb45bqbdTWx33hrQDBVn+QN
RhBBTEB+Ugl7nqplBRStRAUmNLpivMo8vS8dFd7z6FcxHISd2omcnlv3A4GepySv
aDej0yeePHT6Wwwvvg1IkmQGz6ej/xNLbyj2EVZZvOWfQGyCGMTCCL1/pe0V4RyO
WEljx0rzgx3iVwZ+dlMgfL7myiGXBlLscHekOuVVT/dZk1kUEHE0KIyYQugjZjg4
9eYmxh0E+k2e5sMFXkQYp6mQEGgRWjxvjKvvpi2MjQMOFwlnZnvB9jSuNCd3BPwM
z7fOA6CDNPIEKfOmLesLtAjWbyxp4DzqpKf0VAy0i6wbrCC5mU4xRga9zQgODI4e
FQsJNFwcS8GFXmT+vzadb+29+8ejGzTVyWvOHwZ9D+E5FVfQjKGjCbxAhiu1BabE
BF1EoXKd3jOyAePjXVnHwkcGNHqBXOJSrn/B4BCZ5ZMlLj1TO+LTwyrzexWr6dZ4
VTJu1tTE8S9JmPhG5HvnXK2tks+5X7Lxpfe2S3EUqxY9uuQSII0Qv4TZ7h60DDrZ
ZGIPZpIn35g2/FZKv8o57MhNiiZPdb8azCgamGsOfwQyiMkAPhR9zKGKKAedZYjj
2kLgVrNQCLT/dLpqjcRg/O6zL1/oE5a1vduiyvvY92197RvmA/4GCTW4Qh/DjXgy
O80bJsLMJ/gCuPi/hkOH9+XCk2zPIzgMSUalbVdg2BE+LUsjaeMwfD1fKCfGB9+f
kAj4zi9n3MpEWZHi9A3ZxlDnFgglQnrfNJEk3fajy7lMOZ5pVq9L8DtGoEFJZ3qV
sXZc8hf+43t1A1IVnFEri5Opne5k/XRKAdOI07iVtwIxLHqlwbT/GpTsNysR/CO/
Ti6E1NUq6WdG/KYxRTIMCHsDPaZGHlYW5FMuovLarfaMd/JAZ0w22fMAxQV24CTY
bHtpak1LPIqPogGGHo1xgunhimz1E6i2oPnLF9+7BnSPe/19JXP1gy7hZgu5kEEK
0Gq0NItTAzADhodpLphWoBsbXaHyzsIp7z4SiZQIWJV0DHgxE3c6g73eoeyqd2L6
8QwzGhGK5qrt4yNz01MC7a81qcTLCnQEuGry2kyHGec/oyZkCZuiYEBEQoxRPbiQ
wTreIispKYz7QfpukOc2l7+Q5GFz28/s1gvM00oQBw6a8APYUrVliwAGWSEYLH4a
4fjhxkwPJrvXjTiZVhPcCivv8Ik9iS2tb2UZprFEOataDZq92Kt9rzWqQz20mK6n
hjsHX8haidxoTzTfstuSsIIjQ+xP07B/0CW/lceIUGsoKtowc65Dmn69kbMm2yok
BHmojuXvLltQy+yCbgzkHvUQ6AEJen8v8tiBdSlqScvj2nhnMjBMl8OoGNje6xx6
LjNGNB6KsGPhROo56ViQ4Nfr/rASsKVN6j4hLpjVWTqyn7E7GWkjOG4IWr13kmey
tWEvABCxiBPOe7msg6NBUEBYM6PbBJb5L2u1p5knV1IrVnP2oOcVBbK1RxaQ4Gux
CQ7e2NFSALRlLqlR+RO+VzMwurHmbfT4NL9+ZizvT9NKLky2IreidPhc1+/qtByA
HEQEW1eS/4f5oWx8J+inRBJzQj5LjPLvs1s3OsCrhKpkblfJCrLsBc/ik3kvoQCx
ehOQxar3r7rifND0loFhEUfxXnrNJFEQd2ssG+QgoyMd9hJ8N0F1lo7ImlHWMly0
WmUeO3wMXK1xWPANS8HraUOLUvFi6EIP4IlBjXktC3RD5CWbvJPfcitG10wZ9NZQ
fehQW+6vlmRQ3FKkX6eM8PtXdlORS54/93yIDD6cZEWbWCeEcENK6w62RxLm4YKy
+Rg8Wpl+VMVUHmAk/nnzQnAmeymFcSx7O0vE2XYc0JOhYu/w0LJoAgnFNC9M3w6b
A8rfhaBs98hq10BKRBhETO2XlrhfUkRf8VuCvST/0D67o477j5xS7ReR5T+AT8z5
Z/ZskYK1osKaBcZgClHoVtY2NXOVzN0fiurJ0fMw0LvF95ZEU586WUSMLh4H+dbC
//jDEVmr+hS9LrvWNEuZ9eBNf1k8ib6CWKaW3TWcQXUiJaqqq3pCeK4cP/1Ayk4V
tbG4xrCb4mOvgXCmytB6I7ilc2MYCcmUPk+wu9d1ao4ZpLRMdLoxLLmwrtnpKvW9
Xa+gRW4fzptyxBTKMaoWx8VrsX+8/bHb3f4k/2YMCSfmR8STXuCqMMI6sTa6Hn+d
Zo3QqIroobOZch+fCFm9JUuneNb9vDq6r6yJTHfEoG4p00Yz+3Yj2Efd3eKdNoS2
SqdNoFZdkS3knG30V3VkPWNeejVVXvmCwhRy+oLPc2uM75gVgMi8CElaufy+s4dZ
xF0w9D3bzjDBfuhe/hQZi4ouiRfPw6qXmFN/uXqwBgUI9cAl8OtLlcCABdMBFySN
qHu36fkwt5ETcoQdaic3RQiKom1VvcsDeqCmBBe7D1uAELGM8yafhAaacm0BaLJT
+bJ4psrSJ4UwWZ3SbNa71VMRKQnpau2nWRAc6WCjQuNw8AD0JzuKunfviAnH9czY
ur18vXViHZlHvaGMWLbMWNWS7Kf48sB6EEh5Qngg+OVNjcaJk8gjWQlnsBDi7mZr
RqZ0FuMDHDeL2iIZ87+VvfPEQwWyY1IrKRmZVqkdOmWcdZ9S64/TlTDRtdcQCX/8
QPmbH7BsxfIbvyWutTaZWqp796Ok1uQF7pU+uC4s8xgyl5j73mL1pW/PassZP51F
IR2ipVSGT9+ebqpLzXx0q/+Ve7zCy2iyBInl8a5SsFDRb41sHQ5qKOvGVwYRZXN7
GZwuQ78IfupkfVHVNQneZMr3NtzWnDSqnsQ39DyJ0ybSJhAINRekiLpLj23A2jE0
OIh43Edbn8yyNxWgay7uTN+xlEquEUfnBaeVKXoZGKS0T07zHUsZfDbLrnXzU6kt
NnlbeMcfhZPKP9SzfhyKtWjE+ReuPxEcmF1tMKiHMj2zmfKvje2ifhNAFCJvmyvi
0JOwJYIokilYhTrr9RPWrgd/kBzRr7gekcMDhrCJsANSojsRdwhLA2TnZXD9LIwQ
5hBC1WTdywQZlojcdPfSYt1E50kc/DVxukt2nK/RaALbWkILIh+xi4ykrs/Ioubl
DD2VAFNmHI3qF3qUfzCW5KkPMPM5iCpTf4yYfpr8BlNt8kp/5I9M4BZe1icSwwx/
qZjHWoApQlj7woGbLu8WeDNLgrwx7E0l8YjfWVQ5rBh2I+AJ+CU2DxumRfHXqVCU
u4EINXxmXxZNQx8yTZ2AqjNRgHRDodpkGO2yOYOeZc8SgAdluqilgPKgqV24KjcZ
MCRT9oG8iI7Z1R7ta1pkFt39acQddL08kj1E+EtK3selx/Vw9id3xz0RXtDLaEjD
e2tvuln2Htrpl7Vo2/1ZR1CS7eeFvDfepx0pwxVg4Sj4ULsQCdXY7LuarpkAAtOH
vY8YiniHl/JQIHaB+a93qFEDKYRzvUEtYb0gV8Q+bvGxAqk6fz6TjORNNbqFRIqD
ZMHcVnOsMywXMfKE8EMdpnzSCUhncw2VmT4seSl+dN39crFU9EodOTcC/Cd4oF7l
YBPEG/491LS0hyNhWTgsDhzapFV6lJDPZPWwYg/WvzASrpgKAXTN/x3lWaUuUzZ7
xvFa8u4U1Yhu59ktbvGgCDYj3Vf2HY+e1BNIcJdxkUz0RPgBwlHOURm3XOXqu0Te
Tji53Je38SnguouavY/tiHdnZ8Jol3frN/j43n3JwqflD+3zCMOaxcYfGxIQrmq7
Pk3IgJWyeJOBe5aZtQxhJ2o1rMU0W0w47nmm284/N+bNru3mCrOCpQTGwdmIUQQn
Y6ESTathHiSLvD//wZ/HkY9Z9jNu5kev9IsHjvY7+x4k3x/FQwNfYAFqDRBUVJoe
yxSZAJV9Gh2LoOUhWO7SDnvIbljf6n8yTMn+dp9Ke9RO+ZAwbW+DjOJN52T8NeLp
vaxVMLpKKB+Ozd0FziMORQ2N/Azs6yOIDufVFgs47XeY6fb0Mtl0fjQX2qLCRfEf
MY/K+rpn0IV4Ccz8d5wjBNCrQsoIiOBS6bLdHr63dxLr44IMoypKY8IryHKDJfwo
D1pRjrW/ZHYj8+bZbvQSuv1uWQyhZ+CIivjQmDgTHcCLID2CrDDokoPhDZ5Lm7hU
PCOqVO9k+gnvrSdx4REJcO4m/p4HXMotRlyVE14mldE19EUbF0EuXPZ67jtEHdio
pPQxeKD7BFW4T/Vzk4ETNmLTIZO5SXPsTvB+4BttlNXmS/yqqaZ4bl25SpxlpeUn
vcAP6RDO2Vc6+Nt7Xe9E8WzcsN2UW9oH9nAYzc5NwGOQNpqY5s7U8iouuuMW4zdG
KtDsWmts4KBDYVZTUVbr8LD70OqTIMkUw8z264FTrQClKbUikKlaBhoJzgGSrNYI
R62fm1miPf+AOqxhK0qRQHNPuO0JAJh+DhMmLIQcZVYi6v613W1uZ/33Nx0FbWno
HQxEf4jJkrRXzJ/BrN9UfscOZ4Nm2/BpqXV5jk72wyVgssWfwv04shxvrDqY5ZQn
4bE8gbRolpspJu/VhsmE9tOCQcXS1ZHcCWUkOEVoUq9wzx5tuCJIuwGFHP+D0m5d
TZUE3uKWi1jqDZLxOgC4O4zi25G/2UtoX7WVxVbHvzKS3ICfnr0iKZKjqcoEEri/
p2W2R56izzeA5vK4wK+jI8pxO2ZWDpkQ+mRSxPtdqF3g6lWug5A7tEjOHRdWt0so
VKwIJRE6WoaygkmOeaPqxGzSQuNLlQBYJUa5rzjMdIikP43YsIohU2pGBDhxtNUi
iC4Yk6qcTV3huV2f+Da5bP7vTYNXMMb8EvheBIWrSaEQLPZG1VuZLRN5mPdojwqq
Dr3UXISSwz01dECTdnb8Zrv77kMK+42qvfY+01v7oiHQxMpI1UPMHr3ZwKNXFIZu
JTgwSE1aEqod9PQ/lzF/ZquvR1ISdHjZqX4noTkODZxKI5jW/NV3KDQokLidv1Mb
PDkq//TiFEFCA5udGXE3wCB8/XfsL2kRXTs9v6oACjm5ZTUCT+XNmtFnG60gr0y0
olVKlg6hFm7g+dnJcqjntmVv5vxKF4criPyQb+tpKcCQpooUWsmK5WIsh1hrGDfP
kqnEzow3LrZD2VWcURQNOsel/mR/YotXMYKLeLnX/Aycq2f/h7DMFkAD3uy0CzAH
rj9wQ3fYUrOZuUEXfVzgBp21RZuxEKURllnRxG3lL4ef0Q2ea7cW1xJwf5Nn7Us3
Sa4mSaipKl7Fmr+2hgLwbIGWUnIfnz3c4j6oPFMwY+QAE6afDn4hFFu/aldQZv2M
Kgienyyvbs4VW8pb5Mw9sZcw4hy/2Wd/MP1gz0sHZhSnMR3nDHijAbXF9w65cJ1C
mAVQKzeakhuEFWjKYVcAZAanaJXNoBFnaRAj1aq6DOpnhtI/IWuHt8X/mI79b4Bi
r9jqR4JsgZ9cK6gzUDE8xL7Iw8raH26ymeQEZGTXprUr9aKXfD18hswUarVL8vEb
HgQC2uxCX9I8pbQBhNZpDRK3PDWgQ9reGxTk9cDq/GOBwh46Vkaz4fiXfWuQZNWw
5knfHTG5rcsZeQ0jL68t8+ztrNkYYlnfjApVkH4Cep14vS2BYrBv71uJHVYZD/Js
SfLk6HororEuOu8oMqJv2J/RSz1db7L+JqDQXMUOwhRXq9eVD/0vp3HAMe+PXKx+
d/OL8k5mtY56iGPeQtAQ4YFWOnE5x1ujuM4fj6LW89zCPIw0m0Sz4SwI/GWMv8Zf
vx5JlrpPwFqIrH9iEMID0d6Bmg1mDxgi2s76K+XoVI5EHcr4aVH5/cbKvNaHAPkH
isV+jazOhzOfT7sPAdqkAflC7dn1mwrI/0eMyJDZlJgr2dGnXUw7pOmTrkJ4vCn3
zhC0u5k4lVBh67LplY3EGQbU8z63L7MGDt+sPnVQVUuTXvGJhim8V0XAtTb1fXxf
zEaKiBwCx7+wgIc3UOgV1c/90mGou0H/+lr7ADt4xdwAE0jnWRCBfdoA6d9ZRsxx
bsdeutvpX9gTnaAqV5G9sDqTTspYJ7n1sOXd+SFLNiG+qh+SPEpLgzIfjPuGCo/j
PRfS7+gg+1/+T+UFre7ZlpUw/n2tIaxTwN3vgiKAMUei7cz8y1JYT4ogn4BHoGrM
WQpeGccQmVpKArULJWlryWK891YiqJy2Z/gMjsX8tIRA6gilj2z8SJfHpH7ruyRQ
3uWQS3mm4s5PWMyCq5WbPxt8tXc3Z0gWawuW+sdZ0Vv8V/2Q7NrNf1HWaiuoDRig
fglvTsssrVo68M/n6mWikykk8RmBPP0fcFbobPsTjAcsZw87ccoXZaz919+hvOx1
5K926R/gEDS4Q0GWHBYc9IiZSu+jycI77q5AfpfqG4p0NVKKHpsRUnCPz+8QqeHm
KYaf5BNQVYXDHN9roWiZMPzxCOhBnMmgWjlockkKPNyDbdhOp1bZ3MlJiv7gQvDk
nACKBqkmeboMxNYVb7PuXx+lv+RmNSwCgXPeEoNZeq5K5ZEgnRDJWDKrrNkFJE4c
y/GpAfQCNnzhc65KQfMj0HU5AzZrEgtLhMWW9Qq94DjXsz0j5wHFLyusFgC6va4k
wdpYKMp4jIxD1RURoVCR9gxDQ7TWzxjJ9yHO16vi1JMSYD516cBvgo4NYSZa+i/n
JnNgKLqMpocPJXqs/liya3fSwxachHXQpmSlNa977vb88HQ6kpNVogcBR0UPhnz3
y+k+cTqnILpyDAXUxqFGEA9ARz18CUeI051QxkVRwE2GKBPB7ultO6vQl76usCBy
aY1S7ydglNqIfCupFn9kiLWXLh1iNCsktSH90stV39qts39rXcvAZeVprSBXUHk9
hyrLEbGiUUsZo/dHFwZbNWZMi8X33XOn8mWwgAwb48hgMU32ijNR0k10WLBkOhn0
T1Od00PX5r6flyPvI32XiZjmeNiNs1MSVehGI/z5O37Ce2N174z8M55Al8pZGTXM
mZ3xHTuct2AtAS+/qWC0IiJ3AfLRLbJ2hK6qRQJaRmUuA+VlvCPVbp96c0uONh1e
WXIf73G+WNrthJkKeLWcZ3U7vR33cVt9r2acQCa/tWzhfHGWkzerE7tBrH3rgokT
D2UQ4guZIdZ7Q6fgX1AekT+ngRt2JQlu9s42AqWCHkPrGMmiDn2BLE399gvPDmpe
XJgwVcG1dNrrUOT3Diiv8mXnqKdWz1jb4hCANhwV/FTI9e88B9EfJANx2fTD2zVb
ny4KF9L2te2osKaI2bwz1JPn9+LwofyOTlZRPDDP3jlh7M7ZG6R+9OAvAS9Ru8W+
wFEx9prNuSdrPN3APAqUoKMGmanUSt9YZQu/rQ+1N5FZkD7bcMx3mSwpJuH4T/SD
uHRpAHBTiQLKtpmnt291cspo9ef9A0LPyON8D7lhCEyqZ5d2cURPnr5VFuqG6c1b
kJhjCXw1MNXcR19KHtGEUQOmpNKKl4z6xGkYTWiyQQyTnHI+6pHhibQ8ZzTUrIA4
lbVzl0L/H5VaEOlKatNa1ykgbx4jouBO/NUDOMaSXKXzYK+n/F3BE5miO8Q3cpj2
pVohF9vXQ1lpDjkyLAKB+FjKZ1/98X5tdJi3g6hniTCa3kxfE0MXbZ4EUp4Fn11k
/4UaKP8SczQRO4FPx/S6vT/PjJP+5Y6RclK0rlIjybYd64nhGgGndRN9BqkKiKYq
+7kfAgYXmReJ2ThZCPd6w5usbf5f0TjGZ8hGJuijDyksFBnNukR762IGEO/R2GaZ
xxW6NoBaQeL9AQ/AuIjzHhh2E/P/5ntgQHYePUFXi+VSYsuAg4UaJPsg7f+iJPGL
VXEsRd1j5ZVPUdYWPrAlVtZpTesL7vOkK+l/NZKUGbX/aWJbYWYUCJUMdxhtMhDD
8OTrRLtlBPBirq+rKgH+H+Cc754vS9bG3Ftgq6m54R3UO1A1KJEC94iBBYGLXUqg
Ae1A/slW5F+H1zKorrsrmsLniwEbLq4yNrohemaMMWUzJ4qAjA9frDG4LkjwQDEn
BlZYienqEplKdwDKCSVbjd21JtO6Z4hn7W+uzpc6H1jGNEUwzJOA8DUlp56kz+jO
iRHZDdTOyYmvVDX2bfS1lgo1bD9ynSheLzzTGMHjdpi+UXwCRPPsRAc8zYj+7EgI
rOdkxuXr5AZ6j9fOdtfvjMuZzI0EKc7wN9I+CBW3VXM63rglIqup2wIpFu/Ypi7d
/2UTyqPZouPouaSRVmpe4edHNNir0+YRV24HhSNMdz1M1iYKmEclT9KZjRsjEQpu
NTjJt9qxaXuIFYNdrTRyby8/Jt8Cpz7a7bgJwziyEZJzEE7emsJwj/4YoB0oRIxc
J93oa4AGD/8LQT/CTGPNNMXdD1kZdM6/DbqSif+EJb5oGcfglP36fwdXYNaRedjQ
lSfrGBI1ec20LB7WFyXKhBGAn3C0Sd43u2TvoUaUcLzIwBkjaADPFLnH2kv+ZwvK
8KI2/QPr545ZZYLwG/wqz82MWmRkAatgwWUFdmeQ6CLLQ5zc3GcOij2NX18HzIIi
5FA1j7lAA3Cb7v7Vfxm5BOSR34cZhbJlol2chx/hPEIaIq4gEyzPQ/HYxHRP5o4b
m98kXOx1FAH2zbqXp8oXt8m0twDdAlyYd7YNMzcQcCpIJDXCXuEssZdb9qmx69Dc
xit1dHs5FziatA50mXknRfI2JkYrBmG1u+9OnZf5c3Zpigy+ibi44F+ND50CWzqY
Qw2HzSe3QvZ52JIy9dBgXK+MXKpD04NBzJpwZW7NEjU6TAAHNRfRhB3sqMzs66PU
TFP0VqtAM1z+D8ACVc9HmpDsdNVjZCCEM59sSk1Nif48hG+blffJ13wMTeDFJ7qr
8iRzAisgFm9SU6XXFCG/OpPrs5sGQ7vBPHJQPmpFQUD+OSRWgPAOcyYO1TCStOb2
9ZRm1UsYTBRwVzKlEHXeV1wjX4JgzSXBkTKjQQLVTi4fKDxhdxnqgZjoKsdhozPR
FAlTvgwBzxTnbAZ/+KMJPWc03h+ZzrP6gc0xTkWn/TQCYUePSN+ufSe0dsEcxrSe
DBH5Xk8obYvMSGy3ujaTgJyexqqGy0AcW5aGTpAzpod5cH35Ru0t68KJ7fyf1L6z
ElDUHJvxh5l5TDxKtWe0bEbV2lEyf5Lud48JG2tomTkd8qLTn+fmDMC/bsm7Y3av
O8bbGBlyHy3kZTC1n3lvAJ0BD62iWt7DePZsqXNzf4rEKHE0TvUn+MzAhRQv6N4q
0QTYZTlR2buogYVCpu4Sq79nbMNwm/ElK0Xd7LAtyLxO711pJOXMhTaInp1CBLT/
pylfm8MnlJ3f9N3sAwXrxsXp/KSOv2/uRakScDUz2sHrTve4SFx0J48zazsSxZez
2/vxrWRXZxU0UKfMjwif8kBrXiRZUS/PhpBXV1tjYQFikmG/aZ+39pGmG1AARVCa
tWCQwY44CtBgyUZeP/KQy7RgmZy95kFc6pSTyEiR+ybV1DGGqNpjIpu/3lIhIgXs
VpLPbsuaGo6uRjJY09JbkO9I8jlAI5TqVhVh4gTqBVf4AKztcshozUwtV8PCV76Q
9r2nkkp1OclwJU9NE4JCdUFRft8oEgbFYnVbYowSaH5EJLh/d4csya+BppL8CN3U
LTTOHwfxSgWlbbRtYEu7W+3r1oAmHjPjezTv2YuJZMaqM/l0XaG6LIseVbGADgzO
eGZBFGMDi5BSdTYAtyWMYKAZAFhsVhO54Yqh6LtwVXMjvrNKAXlYIdQxXW27eL4Z
hbsR6MVxhXTAeELMoYfe9c6+NGvvnhLhHgcQxrzaf2XeCeW8EAbUNbj1sBoBNJpW
IjNxgQeb9SudyVTJEIVrC0F6b6qCDd18YK3oZkhpepLcRWLhZRJwG8ZjBQypoFSk
JMh83A6OuZYLiKfmTrFgzeWOSdrS9WyLPcbfO3eTc2QpXclUOPxRMZnjMmwTOz3z
tdGXnOwTasc/CJON2W47OxzMd4tQiWcu9FhZx5yeQ7xvdj8zXPgHyWumJhRcd+F6
PTIJkX6Xxg/tJeGQhQGH3TJ/DL3iv+ik9n7NBWb+3H/ZfAVkxFqhmmhcc7dfLSG4
5K5h81pEONRFcI+5nsgqczZSyiwnSA/3nf9ElJLLlm1z8bytLmpWRIjh9wPWK46e
CeAe5WuQ8MaiIJFqztR/BZp24MyzaQB4AbY8IUHTORAw0U4VaytPNdKcHhGYDGtQ
lMWuQ+BK420Zcsgslgu10DsYaeNre36dsIcMogpXcYOsYqqzDhev4HjHV7mOfDkS
iU0T85DOoG7zsfaKC4WF5yYULqHT5COrrwYt8aeIAZAA6R/TNmu8X1hH++ZLwiSq
Gw5fFjFIxV8f1YH64hFg87543D3lLXC97GLomuNX2Ht+xVkarKY6xk2BGVXhKqKj
YXODaiXknlH6IpPscHsgKrF43kuZcz9omJdmtd4JMTth4ZU1eQ0XVTNaY+viiDnW
prl4AbYgT18gGYMBTkkQ136CmIFg3GhxroFCp6GPQgVpUUhw0js84ySnFHpEvsz2
TajM6ZR6huVQfoaqBUvv+wvpGLMt6XLXHwxAEp4dzoW/wSvJQdL1B78CvFNHRQ0O
dVGAR+zcqlQ2JJojrmadWrm/btn/NMWOPy3ss1EXBfQ00uDdxiEEZ46Ya34j8w5F
ldXzonPFDeXtpJ304lEivGHBbhlPuQAa9TivvsdH80HlgeGN1zpGATMGGQHPWReO
8tmON6l0HGApXQF7doG5FWK3FiD6DMNCGBUfkAxytreOSh+qzuLkE/pyNcZ6RbfB
9b1UYn1mR27ufa0V2zeCgOH3It3dw9lCHgqaVg+z0tRxO1LEHjWMzRUfdsIQ9bqn
wc0CZ9HP72H1uUQS8PrgFfD55/xKooRcnDqo8CvCK/wrWVSP8LySTbdqEmzMHou3
CWMIFtMGAxRoGE2LeY0Axv2U5DxxoXpNDGzBU1fdZsK/ql1se6XXtoEpWwStBCYO
FbZUqGHKeALq6WPLdcarMHzA8SqMHkFA2h4aauKCh8RldUveYu64yD6NigX7j7Rz
40KDZsfF7tCB/24tRosOziWGypOobS6XeZMziLYWgaCtQyz6p9oPWrmc+bNJ4jFi
lypIncXbGFiiI4jXNH7JJY2u+oE63ebDPhYkueI2WH1cfEi5GnfbUxAKeeHTPWWW
4EbtZ1zI7oIrfE8ySkxM4cj0XlwqlPjKb58V5dH5tKwNe5gv+8bT7vK+kP6iZ/e5
/cHgSM/LEAGsz4SxLslqi1vJC2R9P4Pw9Hit+7Y3X3RUb/BgjTH4wKFgeTu52XER
otOwNC4jwhbfxasR7miOUS4WYCg5cGMXBTGLcZzPmbFUi5arOavvq+8txMUJ1joo
3e6pzVvO8xLc2X/zlIHFhZP4u7DUKTCbI/8kD4asGnt9VqTYY+0mgX+u3vk8YQVs
FGNmuxlbBL++dQRN1pNQ8omaqFqTgfufjJ/iskloosnB0hqRKT81sjmSc4UcZzb3
e2BctchmYFGy3PCdb9NULL/7j4CKtDmDyixVKt5lctvc4rfEGzGHdPGairvsmVjF
Rs0M14R+tfvfakqsIsqc2qEiGyhWUOHoTtqCcDwYw0eqAOiZx9pR17IbyN5idrlW
RqGODvL1tngYg8FGKWiUeCepzsIJoKcDV33DOhOivd2mSnz6amoaSi/od5h8z+iM
gWtsYxMgTSDYoDqz4tWp6Tx7hgf7B7DOMWWCtyuL+8EIZZQrrLF9KBty3+ef+fwq
4JOkywcyQkfDynNwlMmE/q9soF4iHWiFSAz8qtApNXw3M/wfJjulT6kii8K97ztM
JOviZIZUeqvDunRwmvtVhMGBqhsn30sXjLSFwol/Ym8Dkh9JjSVZkRPUueY838PE
8S9DuQ/wtVbQo4mSzOIq4rvbJFEGOXljUsfu2NUaCHRPKZxukJ0sbnSKHZHgQR0A
Emxo0l4OAVaCdg1yiswlVONTo0SFYlMgjiApPiJCuor64BP0dVX9wHwP7ltrOf1t
D/4QWcYPrr92k8nibHsxS8uKF/T+fHoR95ir+jgzK/RRsr3yPJRGKdkUlOREC2UN
tlvi2ba1Jj18Hhz/0JvCzZZcjTXY7G3gZF/4dy5VJWl0jYQ+4DDE8ZVKciL/7k5K
s6EbRl95HO8cnFIlhlgHfwi17powHh+GSmSU95EOSq15T8uhqKgmKV8lwoA+Pruv
Llm0cm7rZnRH+7jF0+SDO6d/YlcjbMbNlMIpBOi+w7Y4+eQZ1eKDM1k+Z0+lhzgf
1qTOOz6a9A3eRi7Kx/I9yvSXkn4y7kwSXj3UZPNsh5LQjlH2Q2/49ns5Uj4Db6Z1
zgAoUt6B56qpwkJ5sL957qVfi/jEzq48UqeRvb0KhXCsNlyVD2Vmnk6lZz++1cRS
HUja/ZSlOKRuymJDQ+ifTYPawcYdn+38T0kjHwKp0++G7b3X2qpDzBVupq9961R7
IC+kAj8byCIkGhIc4ITFyfPQMe1Eyt3y3IGsZ8Ik67weSPrHVUCw2aygNLDRTGGQ
JvB7elEmzDC+Pex18aoTUffbrt8kT55hL61ET3DHHuojkadEOsvkyQ3HmBSLzfmz
svaZpzIeT2deTFqd5EUOOXtMZdjR9GnMClfISS1PRGyW5siQ6pWRGDTa+fSiW77q
9H/E2h1uze/Whc37YHjft9LV/NmXQhhOcP/SKmS44mdmdqpumKGXuub9wd6fzIbb
Jccf4p2ADA/CP63AHqeaYJ6mS8jK9S0cv+jQcAEqTDqH1cYWtl9Xh3tkvo2oXTo0
yqC+4pt3ZRnPzTZgCJeXYNKREi/Zti69qFcvxw5wdeoL46+YYSz17ZKvKvpcciEi
QEJx3xkenddsPFSGLOUBMnE6nREz9LlpXkur4K+H6NsI31vC/GxqZws+bolGLC1a
EG5ytxfQSe8wfoTzt9IgqkwWAUQde8NYdmz+4WpMXvgVaAFUca4oDo/QrkpMkuBr
2KWPauHj3MZ/AhW1Ro69P9F8QvB0Lo6xc1sQZ5xV+YeAfgUlcQ0qhzm3u+OJlNj3
/KzyXBxIFH+5Rawydt+UO0LOznxFS/8uK3y8PwpfU1dsyfFe80ABigJJgysQ/lVC
zDvtNFlCN7q5jZwNwnsrTdwPKihyIzQHC+0aQFg89bPMzu7ponrNolwl6cysrXzd
PymVCf8T4u+DgUBgj6e0GpNSOroR/b6x4aNCwHwiwlppQYeS+R2GrIytmGvUrYlT
OkLX8ynhiEoo2hdiOe71H0rSKbcurgfuH6aHXBbvKTnu7CVVBCFMSvDDEDOA5jAA
9VDJFuwvSd5+5MCPl5VkSDTAFI/ndmVOmGB+SqK2Wni+aGNxhPg+cKJ44ta2UU5D
vWfPxVs6U2aaCU22kYzaYAbLWok7KA3PKATwBMvDw/NdaUnQh0uNmAzf6KqO+8IO
3Vn1O4ebWh1A/QHnTPLPg4GblJsd+NAUDrccIRYI0H8LTXLKyL20Q0W3VLGTPM9/
yYJcS1kEEOYp/B+loLGcuEklHMqvQoC3OT7FtcGoRahmjY7siKRbNJPjhDdfJB8A
IkXYjsfwl0mdcCFggtlv1U+3XkIbqATXAn4pQIbd41sYUHaf7lb/MGGbmwXxY8/y
VaKVcqb6VbQnYV7hdePgxCD4An7yjpDqhBugJr82hCj/QaNFQMD7JhvJ/6zh8Yz1
E1t30KM9Wpw1DyjcAp98AlzVDb45VK9UyKtmLLEisKXWiWYX4aEMhAQ6NhpjQVtU
fQTj/9HJbE1xzMS8Fa+K8loRK+JTfzN/U9hgHFAmy9RbNA0r0vUqpTdhnOxNExfo
7l1of4YxhsOUJ6O4WkKeK7Q1KJYoMoFuo9u1kt4UFzzSUvmtzHxYi98acaqdoQb3
OeDSepRJk0KlS9cZIjA8W/NAr0tn26BrK1a0HHD+niS+9r4ct3Lv1YwmLwoQNyjv
shZCwVwNxbSoEKuYaimkTbnhItGB7JSfqLqQcmmXUJdamftNyI2d7F7G6S69kBOm
84hWa4qWEIp2hvzYFAXG6qOTNdt7sh6jjY/Gx3qKv3/L2sJjvj5jIfbnsBlp3Z+k
v8vDK7nWI2PulSVVwBU/9vW/jQE37+euZ8t2sNRyajv/7rfW69OdVY0DYMF7h7q0
2qds4Mda/2/6cihntl0okA3MT1VZKtoyly0JWDZxezZnDxQVTkmv92sJwuc2T7kj
dYBXg9/wRf//vDey8lBVFt333eOOy8a5nGCl7nBujW6Uq+IzOIvTvribWvOopcFQ
FPt3tridnMRe/mxVOsIT20UQg9n5pdBoqizrwdVmAJohg1Ol5WOk3WjdoC4D23Y4
macC2quMPUsZNDco4u762eJJuxhwVgL8zKkEZM0P9JpVgozA8J6xzdDEhQIsD2P3
hfm9mYSliaCY/p5mt7qCKF/3nTzAhbLaVaT+wzbOmZ4q0LSFrLwN/YEh5tRFpOCJ
fGyD3Xc7P1LozWVxqr9XecCap32JeaWplZLCOvf/0wEjokr823gBTRn9KziF2LiK
Boj5ajmptAy1EzLnmUD0EAyHyDrcJu9urmm/CI9kCt0R+GV66fxgFeLkGcRMkPeD
TLdII5awJw1mWQc46Ii+QX8WCHvxncd7diqyI7qjSydK57V58Ngy3go59C+Zu1io
QFgM2ErHvo9vwhkmh3FwU+DpSrWtDay5cvzWH3soEHB5a9/pF2DxCVxds41v4P3W
aJI5cz8S2psnJ0jtWrPKsYJzKVfzJsfCu8359kAsMiLQd48vSaGt+EbUxAoI2tZB
cG3je0ze+R3z2f5BJMbm42Yzb3f0CO3P0HLNR68XV4xLDrjMn+yoVsauO5WG0AaN
++jGV4dr7vaIGTTSQKE3ZCt+o4agarViX3fcInLX7h/5pvOEdJypT/MmHUO1Z+L7
ghMqxbA0u9Dlw9sWNmmF1e/AhkpTvrAEirDcZo7RWZeChtG0O7NBbRurOQVN00qo
Nj7MuVKyp1XR7eCFQpvBHgDueqXVZC/FB3zl+4hLoJ/492c1npQTrugcKkSSOIf/
lpXs5c7LN2b8a2QcEcotXNnmo1/NnAZqLdBSmNRxAG0NX9VdJ9AYtZ0FvOxBYJPK
Z3IyNuwhTpsYaByLlOkhlUkCCO3ie9yxeyRyFB+uAivwkXE39jBFAnnR7ArPtGXo
YOO2tREYhtOTyfWSJvCnM9RjdmipEBlXyd/uablD0nJjMxZMKmF97vuQLR+TqP9g
/tAjUq3aAOfT+UNzy9kyNOtP1KwFPLgm+2SF24U4K+JhzJ2HoreCaWUJ/OwpfNlf
jNkMk32SwPx7qmKABXktC/7L5lRFN5AUJ1AgpWOHTzSS7I/Rh6/GAMFelU1NGquB
VlGmYX+rT/9g7PQ8LnC/y6ShqufagPFJleWaPUx7L7DRxbW+Mcg86SyzrNsdV5Xw
dWVEj+EXDON5sCtVMTflK8p7lYZPeKmALHTFCLEcvSTjPjnx3GULoWi7G4wGKESS
TP1TyMHIffx2MxBz04w9xigTdkS0NPkZdcsv1wohPEhWXAPdTa+F5vIN92eQJRxF
lp6loFk9xumYh3UoQ8p1Oar+bC0IHzUqt3ZuCT9zZx21Zl7nj+MNAo8XxtFfFgjW
6YsaCGfSQpqGkfMOiYOVEXvjq1x39XAlchQ1dbtS++vnjKOQ4FqAQbMrtPN2Kt3L
7aV8mY2n5DrVhSIhmEucHEeMtuTdKjmWMA2nPCXFZcEmwF1ass43um6S/pQVP6S4
v6oZ1wfSVroTn3LTKbxvw2/JviMKrp2eGnE15bfazAbauWDwac9A/ISSH8BWqglC
a3mxoDjM01jef0aJYRFaWibfe2bjGpleeXiXDG+AweG1LpBiRQIWKYjYOh4K3kkV
OR4b9zQwfT8MXi4+GHmpGKo6RJ932luzG2ZJ8QHQydH/+BJDAw3L/RCl2Z4XmmQz
So82Rna+Ai5YfFO2VRD9T/rByOdt5XUyxaC7Ff6VrsWKNKQimyUC8nUgOODiq3cq
IIySCkJu/K4kqzzat0J63WAqPg74M2RGeGogiZx86FphUFu8+rJTkFgr4sl9A/qn
YdQLT9IoRRV65GhVk0jfAdG3gvMVOTWT804WRbm7YsVGoA1aYJms9xrxEetkeqfS
A3SX1xK4a/kqeE7H+ebNP/s3EzDW62stcwXEfLMVvgyTfI2x3vuFfdQIW4rVyqDI
d/sFuCEZIbLr2jnwlLzpfaYDxake6reDE8UHDuTVuMMgM/2C5HbbAuYVRpk4Z7cT
ue08uiEpbOO5DMsSzINqZuTchOX8MkifYGTsHWgwauo9C+nVSKL3hDntXLo7Slah
Xrhj9TBdyOMD9z8dqfOivUwTUZowNtLpV/WF71Fw9wnM8oKXM1DoXnHev7zULBu7
QgjzRpV7JN2rDiLi8a3hK4S1HkJh9ZLFBXpBJmGiBYjC9DXn4Vl/iZPZqzWknrnH
MGuPyS0OchliAvt9Xk4GgpEPige9HYVpHvuw90HlSGwu9CeeO91Q1e+dWW3sCZoq
b5H05qMvYHucrJBRIJ97H+uiF4V3dPJFbbEqq2ZXx6Cn0TiYVxGVLqBmus69fXwp
58P/MOkO1tP4GuMv0hmd1iypIe5lqNNg6dWnQkM1J0+N84QxxdzeisjrC4pxjRLX
OPKJLchVxQqKsLWCEvRQ2MtQMQXiNO+Lg1PYubm0gZwmeL0ydiSa32BbTSckW+AL
5DBFW6w3unKm6Y/Cr8ZdE9j1bpCoCupdwSs62gafoezW7zG9HAevNa33iOQMt4qt
IpPa0ehn7j6YnfcKyEyGMg7GT7hkHGyew0bSTcnuAV7aIVAVF0s3OjRabmCsr7fQ
NXMI6ivC976rt/s7LGlghlbDojS2EtjkqXkjtehajN6w7mhvTSLOp6mKlNQO+/1+
U1pTMr1WgB00S96t1gTXz5ZrCrRLWN8Eg4cKo/tb1LqaTXG3WCvF4EqZh3V/ln8h
htjSzyje4sOHysBn9oTsnlmxoPFwOvEiU+HOWEIWt0Rvkmb34vmnp/z//7a6U37M
iz+mKfN9LB2Xc2jHKlXso3w06L4xQqvlTPsradFAJunDQsVG411pZcdLn2iaHIlJ
XBpdmxGyoAF5QBVstClM7BpPv4TrLNaUgYPpeXsDWtg0e5CH0XmVh3JP9xNl4Cr6
DWzxJcy4T4wdtSD+Sirem7gSyE/MEgcTbgoLkOcJuSbmqsnF8Sfte4UI5uLhD+/o
QwazwpFlB9wEQAhWHQm1SSRSuJS1poudC3CSiq2Tuaalfj6abSE48ny76tOhGar/
xuQWZTQBmswjT/aV2yFyGUOl1wsIKo+uH+h8LEc+ydcB3xSKUXQho0CppE7H9c1f
BUWEs3heML5ggJePMtKAEOOT1AfNfIyPmPbmhEOQKPeIJASGwFk7nWywZXI2qXHY
e89EcKSDFoEWD07O7Kahiea8aOs/GFyxEiZVfdI2J6UHY0e5XXDb3S5gKAVXC/v3
ptzoEhitQAHVSzRJ8Okou++4VBj1IH8UH25ywuDCSdiPMZtE21+f9LiRFlIsOwMQ
LVL6OdfrikI7CTi6WBu5ZKLjsQfF9zv5/F8BRLrOpRaWLULinzaHxk86c253pBDT
bLPp+7TL9kHdP51jWbDM+e+R4BQYVKL4E6w8RRZt8La/zNlNBQMav9tjqaVEnpDC
6+XQiXRmi8PWiH2XED9UaIgY4ULhG2QCzWV9IgDKrN3bYCct+FIqziuPVScjFY+d
26jiNzLZl9oP/kYD5RsyK1f/BP00DL4dR/9XAdUGswCuQVdiMh0LrdUZItlNag1E
s7FpD3eHp4Y8xoidpLtGgDSS+svLkRNbi1AM46v6Q3TxU+k3Vsg/ysbGvw39FR3/
Vq1IValR86nbKOomZhNUtF2tIPpeYA5WceOu3J7LM7EmXUBrae896hYXTmJBUfB8
chAB3ls1TdWWuuY6rBqP8afkTpwIamxQj6CNb1BNyVXkbZx8qTHsPw4EiIP1tR4/
O1hSIwX2HscqOpaEs7NDtjyhDehZTCmPGavmAd6PJmmSOC9kvfXfsNHeFn1SjTfS
1y1d11jLN9lu9MRje222bP5R7+e0z+JiFpv0UKn1j/PkugUz7ZrGIn15WzdFdBHw
zngxaZcrfhZXVc1E+4FjVbtJfnOO+k87dTy83gpDlsCOEHFso0P1g1h8DUx1hWXn
vJMnE2hxZ7z4z15yZTh07pauomSnNrcxElML6m7p6J7ZDMF5hERusIWNtVCldKwV
J850sxb9lIINVlUn9JE8ty4rwOXMtPJdC2uXmAE1DY/hxdNxIMXS4wXijIzpviW1
AiqG5RKBwoZR0dcW222RWcFrnwwKTvRZWIFD5ksXxkbDIF/l2hrufwJZfAH3MZE0
bGvO7ieJKkpMBX9m/S/543omADDq3j+gaKesfJ8At89llRayW7pwNFLP27ll1fvF
Ha9sPJ3yv4aTIG2B3q7325oD/NaKbvOP0KLhPk9Gu7bRqnGd3/GFgm5TihlRcUO6
kcpMbVMtKO/vNhBjiuUEOrlF4T1rff1q4YwHDJO3rcRnQhLdyQAv1pbx3NqNa9/m
v4E4DVFlpSh1KcAvLpBqEXJQBTuzDxFce20Z7fwGlGK29S4C22ahX/GfgZfcawiM
o21Mbm01NOMzQCIRsS/rjLixEX/3Jc+0cDM4rXfN0eV323VxnI4EHop3JiiuKUqT
mY8Y7Z+89pjWWCm9KY8HKYiPaueeYKAZZsb/VdguNoQX30jdzYACbN44WDfIpQK0
urwCFlAz3Zarxp2L2SkrDN0bg3coWLcvXMBYcWjeebvZfOD9SRwN/+o9rkh3N3yk
EnkCbk/2Apif8ZfZDZywY/Ip3QRVdSuDQDRFJsNRi8+yZG4znBnQG9/iyV1rGn0p
/FvGEnpzMmDwMPct11JXoHZp01moF7PDYUwVOBRmBohMb4mbZBj1Qd2lOWfX5j54
TEsAFHnyJWNBkJ2xbtn8cwRMtWwR5a2hKAO/6R7w4eaG05kH2xMQUh3nhgmS5P3p
sC7Mn4Zt3k4blMZBSztq/Tdmp3RUIJ0+Psw4pqJTxlBcM4GWAwii31y+N85PUe+G
yXeqqAgCj/agbW6G/GVtUtf5fUbzdMab2b2Vi32qjUjeNt4VTfkIsGg5FiFal3mc
ggNvh2QbUtSr00aK6mYL7ZSeAemUot/1rjpMeft+3RqXcM556RtXGHECxGwzS2q0
xoq1vw2iPSKwLyvib+eJyk4bXY5OgZ/2WMy5nWFRiu5GDagtCIoUPYzRNs4A3TWD
W8uKzctO1SdUy805s0EgI0st/s3k+FNbMJN1X94+j8AXpgyh3RFH34IiuO8jDXfs
mlLQFUBlz++snMVYzPbnj1Xu2+NF8zTY3f6emMAsXKyQh2Gyuy/pyi7eMJAQVBKb
zuHM+Rl7nTqri7AywKMFWsQpxojDfOXfFJqmvokN6/52EFxZKCGeg7/o6UJC81Wk
CJpsUzxDzMuu40ru7b61TLek97j9DXmf1q/kPavyxa3rPFEvgPc0aKpfmQMej8Z6
2e5O9twtqau7UhWrJ/rws2iS1pCsu+nVugyi5B7m9ze5LB6OINU7oMozJ2E1WNWR
sUhHC56p/89dA3rZ33LhnlGdsfj8sWQpB3ByE/OvsWDMXcpP54M21z7J5T09U9EG
y2DqlLJnB9ngdu034Y/PmnqSkYU3YwHOfd4tJUbIwrJGOGOZ39Q3T3IRgCLGVouv
eLXu4mcYsmkbQK3sNyc0KvUAw9okk2oxlaeTBaC+tmSM8Z9yXnOxhzoWom+THM6t
YQwHTAhX8BDxfmxLQ7JUQQ4xfk4e7iyslo4ENeAlNWPEauK3REV5ALMBzTLf6azJ
tuSdfGgcdT9207v6pxLMuBF6piO+VGw57+q9Rd8BqbRuV3dE6XxsHu7fX992RRFG
h/8kyefdBeSCXM+UxmF+l/nFf6iW1LYiQUExN7IB7MNy0RCiYp/8fbTcLGj/oQPH
CV6Y090weT1ph2ZKRDnWFPsUxdWyN7lkZEjA9EyK+5Jrd3kJnr82zYd+wkbj8NYt
MMh3tfo7QnRCj6kmCv5Rm6I+143UZjNqA9YKd8heIr3vjAff0ZwZLL9UdaAFUyTr
Bm9G4Qm8WwfmR8YlyZ4sfanuTHYaJuxCmg2XKgrKdmVpDuvDpsvUxfTwwATNPKWB
1TlIRY3U7nGHAsDMs3TIeSICp+JBvYykZ7AGIq/GhPY1kP5aB0QYlyY3qx7IfZ2+
w8csRySCaYmBhTL8xSjEc5nEZEZ8ZJigtNjQMp0cqNwD7uxF1ng69gmQ8E6Y6l1G
yc7c9e2C/tPQerPGH16vjJ0xDIA1TXn61k+DhP32pxC4yYkiUSEawUVXjzXzKFE1
nUeActMv+fB59Paeqr+/GWgsPbXyuSkffATXed/nsgE1V5zj+xl93GyNm/GynpYo
zeQXg9FpdHTHrJ2TI0FVOhbjvhm9WXiqBiVx3qaQFM+XDI90woLNLIPO6L2fon6F
Kpw/8ATW+clwtOehsjdNngBj6O5t9B6Ys0YRmTz/Va7+LMmvXDCESltfpGwzpZ//
ciLzQYz8aNf3fucU5IacKrFuSVl2vJUF0HhvfvRHP38FbMUW/uCFUP8DuC9AzZtC
pLsjvE1YTFC+L+qNMsixc3arvj5oDr6Az5tLhrOkrahVlgNp8GEJnly7XgAQ/tbg
+OOK8VWuLQGNTzvehsxj6dy86PN68K/DKNX/AxfRdVc8d1sem4vMTi6NnRkrVx8Z
TCD0ovU4V45PtfFmH9XZU63WAPQSExJnFEfJboebVJEmRUsA55O+dCCteOg6iHvi
OkAkfOuoWv8fbQJq6V6cjv9uibKgpVgD2OknStg6PuBqKsBoK7b66JnmVzBTmDBy
7Mhq1JNvPNcpkr4V7LBoXzR9p2B/dNvxHbY8yBiPLnuEGASyZbOAO15E1eChdDWu
OsO2jEZTpHLsqSYIzk2FUk89HKmxERJ9htvMFiypbXImPHS8M2VkKRoSRWRR22Sx
/hiC5c75hAb4C9qN4sayUVyCZ3TBFvf4ou7gjjmK+ZFXwLftaLI2Wkc5j6GLzsrU
n1IFMh++twYTNYtcSAiJAJR9QGZHphqd36fyQJifHrRxBi9qu8wESm4EUB5CQEJc
4AV7JSie5a3K7S9dPsp3DS8r2SVE7EGOd2evZLwXyY0TwbwZQYXFFXUWMkZbdaWQ
KblgRJ+yJQssPDvFOaRntM8zJn32nHShJgIfd59auSyXmdiIAPYTm+mJgSe3MFa5
u/vPn6aVSVo2KWuTLrBgsgh5IRQUZOMm6++Ii+hVZjAupcEbTtCSdALc33AzhxY+
aA7qJNZe8tt+4p9SA7e90KkvW8AvaQ6ZqJMIQRVL8lJ3TdfH41K/v7tx90WQUCe1
QASx2qpn5WCwNm9/73d7sX82XGtIoKDE9+LvahU9DTOKl0sx5wqHvrmYPbwWdZej
KAVn0ksptxs4ubpcWpSVK0mLzQ/mbQsLYSgefL39j5whdWncZqgp0D8yzIyNqktd
x+YAidhVkguWF6xFg84gaq+yN1Lr4HZJrH9odeCNlAZV99jDLzdN+zQVdKs/wD5J
2Pprxcj3Ta5R+asj67ShIetDo1mV9BZo+FGMJazeN2hCLpb1Q0P9dn+2A5f1uUxi
Pe39GFtXI8du+oVTBfBxZOu50GpeRM152oNGOCZLMg1y2LMnbRdJUbq9VkHXOwy4
b8kA60LxauqX8mZls2/HbELp1+TPeLa+3fPAr0l5gwSkxRKT0KtG/j7d9nXW1Ytk
xdzRM7yxinqqV6LtSaVY8fpDBMbsM/sKs+1u1BJ1LG6XlAPyxg0C5AbdYPF444EV
yCQ8hR9k2gGhXDQQrvv9BJCFsPn0ce20BZaBoAltHbpiAX7IqbH8NeaMxkZlsZzU
mis6bxRGZhaV+CvbUC6HGQuIxxavieCyPy1bf8e9Giw6fP8akhG9bQ2MVYntrjT0
jgFfiArvsYRccWveceBgaqoK2Jad+g9pnUkOS2Mi0R4g5JC1fxlkc6JBi9SSgnqc
TeBILohLuF0GL2WuGe8PikUVFbFN5orvyS+ocPx8uZKXp67NcTZ6CXiX7Jx8HJQi
vZGZLW1otU0ShCSJs1qStIM2RzCNcaCvbfG48Z2K7dniirQCwkhs7QbGK+j6TcmO
tjGkysQOgwcDwV6vGSgETlotDIFKguxGzFBugFdtUBNBHe7CoLuxM/4hjJ4LJ42g
qDoNB/RaaCsW0qSI7AIZ/z7nqMDpd1FhH/aA3eK8AFxlpdpBx1z57VXePhHHsHp/
2E58vJJivGhV6FS7q6YlagYJ9BKAlpyR8cis9mA4fEUjYsrVFJ3bfqYxIvXFJ6Xo
HvbmmAGL4SUSfV+opUfrqXeattlKo5vKGyhBDYPrY933vhrCRQ5mY3NJHlTJlEO6
c2pmMD0FQbQ6WaRnQt+8QuR7AZYlll3Qao5HYfjxjKMTpuR+y/vv09S2ClNDwWgj
JzNrWWPKp/YZG+VqSlaJxG7LU5/xieu4WhV5RpCqkd/gbjI2G2PFWl3JybLdcDxx
trEkj7JjOJy2QyAotyr6sZEpVtThUv5SAKzOkhRwS9h9RvLzSA9SnXEhKTf8d3G3
9UgVBh1TzuBH8d3+jaiBxVPQ0ideaxi71p2DqPYN6lc9rWz6o5gQrRvbkFxllwYM
tVtYu5TVFixZODtDBSVZAAIPMaHQwiAC7WxdinNVXikMZrTuiRaiStMz6kC1cAID
tZQmHOj5gyr0sRkpXeKNWw1b93nyn6NibemsNtTYb/zv++NCQ7kLNw5nw861rhB4
rDZANcAFajlfjwwmMmO+Ydjnr2MUZMW+GedtOLaQxa1/FqvHBxFczi9BH60ehPTV
X1r1b/S80GXe3L3axofSirbocjD3X/mMm9+Y2Ajs9aQfyO0FIKbSPXRphSXbZV3Z
0B6TpJH8srDEXZq5RTwdBuruVg+ygv6Pp9YQxm4ysS/MW2weF6noXuGlphV63QDn
cZdqja02SzVhzsGo+2GO52H2OyHP6thg8epLMudWW3+SJ2wp/iBk4MZLyIbACN4j
rUy+zPo+A5YYID4hXG2/TezYjBqSnR2uth1S6fy4H4Y+Zkanjs6piksROpCes2l4
dMpwD/LvjaPkD0maBtgzqSW0hy6Fon1ZXhv3v1KVIlNeyawgd4fhL5UNDkG5OuAi
v8aYqR+QJWFgmm8l1lgF5sf3Jfb4LLCY81MXv+f8GUas+zARZ4XgQaLBdZQrw2kq
+CnxfOeyAtcIGGatdk6z5ls4vKwJ6muLjxglUT6VtRLRq6pYxQMRGZQkkwm9aVAm
iq+TO9nHCgbQ4iVDG819exANvaOm8xgRuVWbjAENul4rz3sBd6C5m5lKqaL3U970
Q0XbBnlIhUxhMrq0NNyjZxwwy2OSTs94xYK0mQcPmN4MxgaTh5iKGDot63aAbQ0N
7etLNnXMJqthtQWyRpgHzKKPkAj6IIstdFXNiNNzRsZ3eOylGXmMI81zctD1N3fw
Qkhe2nc5Pfh+nAsdNFtqfr9K8p/enGo42e0pBp5mLMwjJvPcgwCWZQ/4frUku9VE
fsC+yMRISnf2+9d16DXomBm8fw19QsB8KDjLQiz6+uMhSV9hoRMhSYUhFwm7yv0y
+p43qYfsG5DgXssyVf+WivfHfT7mFMHLHRZVeO8LSU2IN3CVIbOHcss6MCuafO/g
WytHH5XekkJNYtYxsriZYphGc85JqZKbxziN+Y2v3eGM2eqD91Xn5X9sWjhQBoMI
qzxD6zdhpiGNP/uZ4PADy7SbkSq7puMwuR25mAV3mJomf+/cCHhczc15PZQAZTGR
se6za9OOq0VwE0jGTbPKnIoz1NQ3ITdyLY2vkI28K/bP7cBw2hp8PnFN7IIMpGZC
Mwz8abSVavJVvPFFfX1rFcu+wkt2pkuXU6Sueu4dQmysINMZN9tVyYQTn213L9p9
s2QkipPXjtysQGEOZaNsvvE1itvW9CC+FQz/1iQWOYO+mCuYQvsiJAXLtGveAigr
cvoBcsUxkkvr3gKLO9JHdtQ2+ikzJ8UFijANkiFYV+hnNymM+735DudmYIN2coEw
XVgwEAGyczRcphuGexEAr6yslYDpnYgtmFcx+jZOUE30i669fYF04syD8XLgt9kV
pdMGIjDd1EXtQbYEIcut9iTU+XvCtTaaaM2ypOaAVwIol7POrgGtwgNgWXco87sT
R3Crq99BiNqhsgQ5+jXG4pHaXZ7mR7DiG06KeU4Dq3COhfzTqLgcCXGtF9jtqTa2
PWXQhz1YBa+/N9ZfS0MDLwJiiNaDXjfeRKXZeo2pJSE67iYYGpc8lCGm4r6LkOhG
uj8Dn0LHKwSztiFQy7hM3ghgg7OrfX7xtHnjQxe/6xwSZXWjnIaKBa++1ah9eVmx
VxmqIp/TPE+60wnpKBtvgeQ/QkoL0DG9ObdtD+j4q9PWTQIQpFVhLQ6sbOt0HjC+
VBKFhrvBBN5jWIutN8q8uTVtjiZGl7RjpNKJ/YATa9kx1+m1AJZGMzsCxGcQmnlr
I5r7Tg1O+F9zVPZ8/xRxapVzTe/0+3ANAJiz0jsKamZNK5zbjxmok4MJ39eWu+KC
aTIqCI5BR980XxaBwuc1H0ys72IrVMnuwOBUgAvKxZbNcqZ/uX3V5PNcJ8sGVWXo
tA3Huj4kGF8vdBgyXCCgN1OxAX185l2gWzSOH44vk0Wr1aLNVN7gL6f2bUDkT0ZN
8K8hCx0tG4WxR3ZVBhpZthYGjrpdSLkaQxHQZJWBDy0vZAhwfuS5l1Kb4zRLfHIn
9jCQhZhKJiQZiKKWeocL/zZ/XZv7/Go+Q+ks+EvqCPL0Inng8W0r+4PTTblsXjuk
8bE31zDk75QjyQrklr1u6QHK1NEuoCdepL3V+3qQEnqUeQj9UOGmDgBsGcx+88rF
Zg6AJAqkfsdErbpPq7yZVH6fqfyENYOzkeu3CL+u2a6A5/iBZmDuIWgAQ0PiqgK6
qhZy2bM+9/xG/tFQwRVi7RklCNKDCFwDoe+UfZZ1B37PHoP17PcdGu2lAXVroCQm
lurH+zscJIToKcQ951FCVtTR14i1k2LjGkytFhsHiYp05PVtUZJ8C1QzWvgJg7dD
CBZ+utGQ5CXauO64BRaSaSMRLuKEtD/W03uwCSgWCqjVKY/OsXqtKCqtk5MsuOdS
wvEkdT0BMtWCU/s+/S0uA45cXu3wqkyhT/zfGx51rGAqa3QM3NaQUHwbI61czUtM
7sLjOCUBtqR0TJ14QpoitBM2+oGJZGD49YQEIwXVy/MHIo5WG4TZ7XnedkIZpGOq
3VLsu9e99eWa5xSmT7HOzAG7isY4ulAUdNPQFhSnFsYJ1keSUphM603/ky6fvviX
HW1LU8K+Qp5/U6+KT+9xkzdvWXKl1RKlR5UI3FZpEBsCt7WKfmWQVJ11qrZs0my5
ECiZjpjX2CFRiK3Vx8R6z6a7oIgWs6fGOthJQ1KxbVqh+ZdEPZWpYojMZuse4sCm
AGkM4Wro21qjrbuJ++CqY5kVlbojVvlS8p3biA4o2fZpvrPLz0cdTUSpQRIcF7gX
l2GPXdv+wLjC7+2IWFDAM7Y9/hzisGCc3jD2Fhor03/foTqC097N5lgJyqm+pO60
8YP+FEsjoSPODVFN9Xftvjrea2HqOBs3lupVZAh6azwyWnraD6ky4KQtxhlldpqy
luqozEV0F9HPzrOvAORbDpWwfgcqqxF5ILKWrfKM4aBcDFmp9VqJaYgRUxdum5ZL
MmwmGsPAbGfbgl3xUAcKvOEPTZeEcxTnKkIyZDhBysB5xDoOaFrSLtL/IAssO7Ld
hqxye7B779sC4CLZcY/mQMw3iUqbakYIzM5sGGzD6yErOU61tbGv9rv/SecKgEep
9nJq6D+bUkd0SawkEZ+NgbsRH8jIodOxF6iESFU+JGAfLssQ8/Dt18dJZ+oVAoDX
+BeXutuqomccbdH7qjAXW+CF+m9ruT/D2o4LaylXKHglG/w5HXpPpSXQNjLJeYAk
USRx7kUxtZSKfzPQE3kpLy0pl4j0IeI6wNLuXmp3+qsYu2/mC6jaSCddHcW2rT6E
jkBnx+e7+JZWmfhXFolIvwIJf1SjRYU3rQMHkDX6H1VAa994QYYPdSJYek6S+/ed
FQBsFILoAio5slgbvLOvknb7ldseHV3EKs1xPhNGcjGuGuq2Vxi0irz+Gsi/1Zd2
ShBDRUl7/wqoLxYOD9OkHgmAc9SAYtdzLwFPkWhDDWuFv0aZ4ollZwhpQvPxogo7
lAjADoRTwl7w1wfzfGKdGOgjZ3RGoRr/8gcRkmg9ZAbZlf/PjrCPGBhruzi09aJi
xChEtZ74/DC/YPLFqsDl4+GTGMPcDr8TQ5nk7dHRQTLa4ncuuga25cuvuroAHOKs
a3HJl6eiH6sZ24zw8L4YCxxOutobCjYcEZG6UKNjQXONmW4j3bcimbxLl/N0HFEw
X/d2dEIR/DqqEqLlCYPrDMfSSrCjEor0cOPEZLI18neX1VYIyAln0rRq6bRsQRIf
haDRbq3DTeZBsHFBYsQo6sN/Yr0eL5d+Mnr+4+DBnUeKjUlpmb3ctl/9egDWliUU
TLgwAvLxLydC/DBcfjcmjYnTgp8gYKsphSc+fwXgg0JV406rd36Hebqj+tQ+VTmE
6o6jQ8yZGVDuk7gfoaStr0g6A6Uo3J1Ujg6f9GHJpkBqW/kRv8dUXeuxyhTpAb/4
7MMIS7YIMXeVFwuy5WtRgeXSPwt4dRE9UtlSU7aYi7Fa4jEsIGbNyM0/En49h1v6
i+HC9KTL3ylNe+z0shfpdGIkF4313QT0yc2wymYHZNLyI/pbzybdAPBBQdJvioEI
IwM0WX1fyqp4y0KQSJxojR3lva47WNxj5RESkiFMTLclPYI8n7UthNUxxMRjPPfE
kVPIquhqMHhw3nwIXLSO4DG10AS0O8x7yWN9ueO4LjzEOsLVTeE2x5sDE7qp4bHx
vVEnH9QXJfcjHgc2+FTUX/iPElml4l8g4fY832Svpbugz2dMghyYUcRExAPHDWp8
LfRGNO41OKQPuihqJrnblfqFFpRfdz5RBG25kOsRh1mCptcauCzEHwARku67F5KX
y85sAdMxmKDT5+9jHE4vk1AJhMTRdOpBS4v7DEEbJkxZ9Q32+KXgftixh3fLaVO+
wufMAIMQZj/9i98TCU5h9Xv+ZEcfVCpOT3y4dRjlHHkHD8c8NeVyk6xFxQRII7gV
F8/CPHqVjZKQsB+rRT+VVv28FBcGmqfjoH4law+ALRolAi9dQvZsdafqBuGiVrQ5
Oy//kCFVcUYmXMHcX/Fp2kZJVRqDfKGwA3s23nAWy3QcRgkW6gldZB1A21Ort3ep
COMcgptmsg65pkX7ZxfY2fmQjee5pJo/B3SDzqsXrVznSLbze+9fBRi/eBDVEAq7
RjHr8xGbb2n46c7CCe8u7gzyuUdhLGSuUAzco5DUxq2pNHDmD6chTP9i64oNtJss
2a+W8n13uO/o0/UvcA1b1KzBwdmSWmvEJrlRoXtb76fKF3MIDVI29cDpCUjS0NwR
lbAWIxhQRT9FHlzjeHYXv4vansep7AUekc/XEbT79eZ1Fs64SRMSkTaSyQwdimrI
+CoeWtC/y93vD7nlDpL7cXfP8YZDp2YhCjzbVeiMmsKs3m/LKqqgqI04H7ZjHKo9
mmkvMioZxmjNe+ucZA9bYkTu2Wb57i8p9B5mZLtg8gCBycIu/TaYa56bQjkXwngP
WHQH/lrYlI2xY0BzHFGEJg2mAbKNMjpw/sF2AeP8viJ2NdxpJ88+Ge4fEm0nQCOb
R4DhZRpcG4E4x4e1z56Hon4Tsm0cYcK0xxNdMt1XhZumV9j5EBQcn/RK7BXj7ECc
4R4jD4cap/XRob4V4WiAkANWJylJ2bH5paC8d7G9uJMuGg32rZTbViqQLmU7kmge
wwrzcKePNCiJWGwQjgZAO0XE/Of3ZsJGOtKWyPi7LS9dHHtXle1NkI7xcpQC3nfI
qRdortkRM6T9qfakokQhJsth5S4X7tzSM1DG+IXNe/3W5uxUiKAsZWSjzl+nK8ap
bIWAdCGHPTnEblJ21WNhBHY0Limsez0yYfSwceCdcyeiQAISgmA0id6qjfWAT/J6
WU27sofcm7P4JgJpD0gpKA3opV4xCIBudPsCyx8nVV14Uuej0f6GZnm/WqTk4ocH
68g5Go/a5HPALwXnthewg2jYmofRxA7qRAr4Aj7HCP/nJv5VqmdA9zQttAL6Kive
oZUAEFNdieLuDyT/2bOIpuT40OlVHs+Zb6SDE3rd52D+2nY+LyApOuuuGr1T7H84
faJNXAdGtOjadSvhjigOud4WaEoZEpSx2kEn/kc2z23+0enceEKLxemVp0b1zdFs
4fT4rxCfjBusdksFgfc/zUr1fBjNrIxzpKY6CAEzq6x0yqCGdEwIxL7Z7HBl7GGP
FVwg+jlvqm+btWYiVDwG+XdIQj6ErklkjqFi1dTjkoQ2GipEjFma2wfelqZYKHbS
EdJZUUXJaT+1j6frQCMFa0DS1mwEQdQBOt7hNmRiEY9tfpEjq3UMJarEVXaHbWqR
G4MzkMaLrIkQSVC+p4zi+dKndeBDVDTGtPNEM4Z49o+diXt7V/GmI4p17hHoSRYT
B5MLYlHW94sJqaJN/uW7YtiE4+wzNXkIORZuWPEtHpPT4uHF5p9ESdDdfCeBUNGX
wAdXtrDararmjbS7N91IOfLLJp+DBnk2VK9Z5DV/uMy/DV8tuQs8tIIjaV9eC4f9
596Sm8ds4eZokxvsFXeYOyBvy70QDrbDFeErvCSEoHK3sA9HWCebMhf09eDUpAvP
NmrvB4pL5kNc9xxWKpdZm03qJzmz6P2BvZ2629m4xBAUAcxQDMESvI2E4m/gty7j
xQViWZp9EWk/ZdOZlyubxt3SpgVJjuXlMZlt4/YBijLvGo+vmrIiPa2QOp6+dgd4
vY4j3eecSV2RQwQpi8KRIeUlp0UbitQ2GuXqyoQZaMWHmfAnSsYeCpCPO4dg3IlW
iRhV/7mtzBqcDDzCO2jjiw1ETqUPS5V8vX9pU2nEYbYERPf8qnRhJeaZb3v+DfpH
zV49wB3Mk9M78Su1hV+9Hf8P70sBzdhiBaK2HnFXj3Pkee9W85FEcx/N5IB5IA7w
Rny5Q0SUzNKY5Pftmti9fpEc6aHbLmNjt2qtmcBLq6hjuyoNGygUUVw7+CPQ09zQ
iWuF0b1ECHkv1fLg2+ZC0z/l8jRHhyztPKKiHpEAHSEL+//0IC1bSYPSJ2TTHiLS
WXrYKD3//IpiGHNsRGHJuxZ203Z4XCyiKN1jIR8vtt6Msl3gdYc+mN7GYiLNctqR
RF+9Q4LmhOX+tYFNKJXnp1hM6Vm/KyORt9Fl5dW8/OM4oTjoeeC4bUlhJODNtDHD
cR9+AbMTYFTrMXDlUuTpTCQ5Vp0PO0mvF9PbvzFU8IyHdbMrTMIhvoDsnK2Bd84s
7PPYwqBPJs29MrL6pWF5bpR6k9mD+geK5n+eJI/SpO7aY1pqXqa6WpfnpO4VnwNb
aICOPEB+kjakzZzq4tTfOlEG6ewkpVeqVmLD3AlYW+wXN+gEU5aXgZxrUrwCVqmo
CawgZWdtWEAaumCLqU8lF4BCFbhegAkb5dZBtYnm9MrtCFHJbr3f/Vxy0PqR8Bm0
9h5gtcr6MO/Z47PYODs+TwwB3ojJnf0EDZd4jVfXHoqn1n5oNOqZk23N5PpRi5KY
te1/pm4EcIfdUTxFXtImEZ8v/4se0wxVNTguFUYgNisG3yDPRsVcc8wm+j19ZaHy
CObXa5OKp9efO5P6pcGruKjyk+6KHfoRQNE8NtfChiPaOiZafkL+cL3fJdMnbbBg
CjLL+z7kbFHfYiiuSN79SwXUc9WqCHfGBO8Tu8zk7WqM/cMzz7v+FsqBnTZwdAx8
p7xRl510FhqNyZJIapZd3HAQZMwHtpPMsXDqIX49shv7vhsn2yFx15cPVId7v28y
OKjARGx/KJImV7zRveB3ThNDhPkJihHcaiL1BHeeGXwvAuQJUNICudSAC0cdWUVd
toRl2eK+VfIKxB+U2hMh4L6aFm3WcRfRLKkXhdzaMUmQvrn4+EleAF+CVoCP11NG
LiwCTUZwaPYqRVqaXldzLWHe9SpHATXKoqBrI7L5tNYJm0l55oq7/r0C7hRCZcLU
8vBXhE6JZns0rJIDxybxtNi9BxYPkz44nRO960STWwJNqyxZ0h8kuvZfXNwAoH1T
sXxf7t9kVf+D/TaR4LIIbFXT0mopbf2cKCFhctwlj4PpvFhLLQbAZXqDSh4KFzMB
sn3uInbZGYwatZ2JeBLuL9t5/1jgY/9yCB73uz1/WyQdIwBzviyVLhZYvG6gICqu
Vla1Vn4p3sA9P4AR3Zxu/0WPJNjhfIHOxEh3UvdXdMjFbb0JKmsRdmQRnaB8InCN
kZMoS55l9ABdjEaVDVyzvVdV7R7nElSqvSv+tH8R9xpCUW4opo51rDHeRnsLJaMW
Lv48qh6jdjB2tbbzPuZ8LkFdRmh1biIEYS2AazJGrAJy3NJLLcfzF5TyilO54STG
U2tEedZdnx4sQi8jr8zwKFd2grWrRw/F9JBnnJ4FA4JsizUoXj+Q311bOIXrFLaX
jmoRqU0+1GpVZhGATC0StLcsZmXJ0S4kriBKnNkqUxzI7AmbrH4/UoQ42orEjHv8
t6QPWwTZZXm+vjm8KNKkGaZ5ZpAEX1HEnQDYpGZJnqSB0QlEJCDwYE43zrV2Kl/T
xaCLsSc8yjxnQED3wauc/J+5eMU/bw+57FBdSZu5zS5/EGjAdF+OWTewmUGi48nw
8Qe15YI/LdNUNfb+ZPpl/nYD/13l6kY4Zln6in6BcePqfJZpAVeV3WsLd8ErdQB6
JIxbrrjpPeZGsUSd075NxLhTVOYH8R1AIltNeBp6QdiRyKjwl8JRr1kFeW+c2pIK
siYygJBB53q4SGfnBeQCKHhYhfIcahh7Tp0NtQU7dUFoAnezI5vZ4+ft3X0I++pv
L4TfUVPNDxfUlYJQcX4WRZk4u5USbDpr0TDDPX0NRsN8a5TITs81ufHyUg7VLiFh
PFY9untJdV3h75R7L7YgfvA1AvrMBLEb/8pDqBQ4H+gXEgBPAli5ynnOgQnuh0by
/b1yTP/qud302XJ0krlrTsyIIN0lqaCdl37RkM2XypxQL66i4vSwFnq9/nsONUjo
VRNDRtJUAcIHXyCKrSyXQsiriPEV5/ssA5a0hznZk85f3Yq0ivocY1eUNXcfqufv
FdrOP2aipBVJpUr2nbYV20jpzfviyfwHIhsvxu136AG3nvPElBAjaPbI4VUICVsN
6UdOoPqDZNKd+KyRGFh3s+dDfQ9s0rIqBTxUXAcKV8vPuv6Rpos//XyglULoy2Dy
WYP2S7icaze2d3h3VpMjIxlSRbGhc0k5xT3E8UrZw263erycIFl1J/4H5kZ97YTW
sSnoAAU4Kb+eMqILzaWOfXa+am4vTd9PdotIUE17Eh15t67OTIKcrvwIytecLazU
I7iSzWa9k0t1NwOp6NqdyCP1d76MOXCiIxAr+Bl1EVefClZVfVD7TqOT5uqw0pCK
qVjeybzRmk4+KX6FUhtS+fi5EMJVpLGSjff8p3Bxnd6gvze2eaQDYwmbNNG3JCdA
Zw0UrUkrvdomg3HFBfCbr9yFqFGtjbJgZDFl7kUoM9Wn6BqfBPlkwfAOWYiTfSKY
FhVu2igbY4YUeMAgHaaDOep5IcdjWJFeC/edOEYbrVGTDJawjQE3fxA5zbBTKRBR
qpgD/TfEymBptZJVa0eemFF3/d5x20+jJqIDxK+8ALjy3UX5d9kCHCb4vg2gYuBu
ILfEUPoZNRoO2wQpQlH5Pb2ERzkMY1sjCkVnNnR/vGXBDPNBu33ZyJpTxTvGvH4e
Gr/rat9gvYFLrAQDWZ1kqmrb3mXSgGcV1w/7jS9gDTkiE4T2jV12/gC8UQEKXuZs
3v2gxrEyZ8tAXZ8Z9lstzb90mBlAdy39OXHgQir+jMqOZJcjXxH3E7LVpNeYK13L
pwOl8o8gRYs5rbq21fl104fSqzDyMBYJuKboZoPcE2LMfYKRGDE7I5XezkaGfaxW
b2Alp/3adABB+qUrPLhrgkdYBzOypNXlgHYgu9A/5MGbcQ2YWtfIiATV2s0JtVqM
216xBHuAxdjJ+GFNpGN4iXxWPKaOJxiMnJBi1Fck+bv/3RzM+KzNXvz2GqDij6zl
DFw6ePMQw5BEDtllxIe86f//PD5PH36q6ABiOk3DvCJ9iTNVv5MTLB/kqAKL326Y
pJq4HeJ9wdgbwX8muVMDtmS5NlZfFWgx5HeqtI0KoV+ARdMFB8GXsBPX3t2/X9l4
1CusINsQfT5vFUzZWA2JhwjmmlVauHCXEXRp75AfDSSiipaXdvwyYbE7k2hW8OA1
/Mg7iTlP7u45aCFssyoJs6YP+V9E2puLGX+WA9qfu9ha7UpYztE/JhAvUjV80LVn
7hBjxzMlO8FMlFGKwb4MI+SE+gaONYvfrLeyhQe3HMuYQBEhIZ1T+R3ArJvqmQ8A
xQ1guFrIUe8dI7yr9hkiU4I7W/AC84yFoRvR/6p5/fNtjtdrMII8aTRibHXY+Tbe
+C0nq4mdzmlU5NjjnBIGD3kKlk/h9m0YUjTWd8BO5uUgfCYYou7vBM9ZfvWJ8+i9
YxuDwrUBz1y1dGhvL9AF8CAOeFL8dxoezRBOSziDj96dgAeldabtdkjcgOc9atdg
bF86UGd1ZkkHRbWecmcnRB/wctsvoRZ1rxNA8zL4ZJQCuLxqsJ1bs8fhi1ll1nPS
j9V50gWJUnH6kSKs6fpixrLEmUBekYbATb/p9mSrt3sS/IH0JNb+AEIvwVFf6w6B
2WGz5rR+4vz/X/lo2dvAILqx9drVeUsa6aDbRkNaK8KnaVr6WshT28rhTiWT5svg
2pPKda9hRQD6vedhtm2IvQCtFqnW1pwFMtSGUfb9TdHIQ9KxlYdu2agoxVOQSUj7
IoVXC3qDvhbET/5ADOA9DNJlU8lss7DY0wr0YziFQ896kMQrRosxWDWebu6QmHHB
/b2jPcs7vSuVTwlqGH8OA/Xm9/wS+Lo6oTY6gxGabkwTV9cryta+Pmv0kc0xL7Fx
JwMpBEmPr3T+Byc4/m9IIRI4VTytAIz8xuG6mEeIdV+PXt52yR2QSI4cnDhXMBsx
RzXMPc9EK6NOkJcV9Vs3oCvsnXcodF1jrGjnVY760756q8NVYLcoeAUEUlWccFh7
qzGMAKeRIz4MWkLb6BC1Wc6owaZat7hFC/Oy5/1b+vfJZL1WR1ZlEdjUFLpegAJQ
VjEkMhYRhTuxJO8b5DTt+eEfCWulKGBbJA3b4q+YLOdY4ZvwCrhIHwRQOLPg3jT1
HyfRIKarl+VbGQFz9CK2qqrdI6RowaRF+aaUA16nhdr/D7MQVdNnxtyjNdYAs646
Qohnw8rZBQEc/oogdgCFR8A9Yor1uz0bLqFvWCcletgk0uWLNmCt8kWek84DWZM5
DGlFh7jxO2fEKsJL8Dft/OhHVlUeKZHuRceKXQ2sZEbQ3Di1zi/Rx93w+xLAoQ+v
ztKGyvDaqSuQXh68w4Nkp9Lm9aSeJXixlr72P58Lnsi9AgotsgPdj5fb9hptJicN
Q03ZQ9VcyNHNe82qqzXuABqgo/eTG9Wlxn5Ti85dl1+eWtOonZCamR3+4HA3CT2v
hXUUQQ+9oAGAd9DH3d9PjoYip2rIBFckTJDF2gv/psq5sn3vyPLJif3RQnegLydZ
M3FWjft/X7uY91OMsJFRthZp9RtcfwQ0cydqKMj5ke1u2hDD+BQgP6OtBu9duObw
V2PkP4fZAH/3Yh5izPwEJUVsW7ofDFoQb3X7TIdq1eWSSVuoq9VFyF02Te/MDkHg
TYhYNgKFTdAXMs2UwSGIevYgidJudlEH2BJk2Cher1CTD7Bj3u3VOlt8f+tibYik
FP0SttfGCPfWVzi3U96FeTiaxhYLuHcM1q6n3nzh93VSFD4A3UkseF6uGWXMvVLL
rDN8LmOdmp8Dp9apAltMhKz/e/XpGuqNVboWV5BQ3bCdwkN5BMnHLcvEZPW6Op5p
WAfbe8pfXK6fjdROs5s/KEFmsaAtCGXz4vCSduNAJgtcO4SIwiEIwgPpIq6TAb7G
CFfnJ9I4dFTj2NOtk82a6SN14/B2CKgEiVoAk9uOoy8qNZRInjhWHOa7vHMoXm2O
fOD/hH91LCesFzLP+3bxriHdMuTGlezGmcVsRkgucp7yzJdGoxl3MpfkgDnDj6Ot
leuaI/kGA4EGqW7amCbMs05e1E4inoWKiUmd42hw9ZmC/MMpl4s9IVJi5OBtLg3o
pZuw3mlt/0ZHWqg64UQFOfqVuwiVVsJdhVcEL6egnYIeyd8PJ0k2JbDd6H6TbJ4E
gbgIf3sScMMUIPYU5gfUiYzHvj74mm6AVZGpwLXG9uoWpVNGWyKmvI38fLP6eDo7
6JjW/yBwYlFapLPpWlx3xP+BbizRqPn4v8ohnK+lNqoZyfTM/cHkZ9cIkTvhTqQ6
oS0Q7S/5V3BOJ95IV5zNfASwIhyrWXEBzywQxppytrO5SNkdmUPVJaOwSzfnjP0D
sQHTwdosFTx+KXuE+ZCCYsm12tfBncdiD2fQOxuEFlXZxlc1P3YEOJTSlp2Hzrea
RBgF+TIH8SF86AGEjB0EiDLqQmU4kXJm7Rd5tBH5FhtWfrvh26mX+AEKQ2M+eDD+
jrPynW87vcilAd4MoH+Bx5F1Y8rL++UJhCoHRoeL4EtCPLTRod0Diyhryd74r7G8
ZMqujbfJF0nLO9jQ0NzteQ3eIN+KHl5DLSn8t/u0JVxaFVF1bpOZttqA3D04G+ip
QSqJ+oV5eV9QyIctaX9YmlS4O8gVINbetK3No3XJNwA21AwYHccMLIXoZ+PUNLyq
ceJqFal7wr8PeSnF9fzrc8JWwEXhymR0byFcBmG2TesbU6GWWHfe2qLuseP1Lqiy
OUHJdL0CbfON2Itya40eIp/8Q63ApE7vPYA+yxUbcy66TMmZbtHnsGcx0is8NjS6
uJpDtQ4/KmHwURmc5ZoiMVgnVAA1K7LPhmH6mpTHmgPr0Yux4jhszZ8enPbWgDou
bqq8RHQwzLdVM+YTYjvXkQbi87TnpDa4qcMk4DOkqAO48q0+rp3n+8NEwORVT0Pq
wSiUjRQ5iP48oa1E+JlSw0LKbdC8HGsIdr72uZo22DFTxZUpCiO8fO9bV6jha840
+VF9Juxi+eFDOUvoesoBiIaxbpW4D1yJn4U8Q9uawsIrSZOMZM95gBs79fNGFFBS
+xtJ2t+1HNgWUpqGDS5vhAKHA2hFvzVenOPY12AkWuD0o6sLMMyHC118/QRwjAFe
ua8t7QAFOtN43VOryFfSQ+Ig7VlvJtdKbdWUuNVPut4xloKjHO+Hz+3rHgjUmCri
JHqoTET/qXJs0C6yIzdw42bMh0xedRA6Tr+04OhB/vC5OOKacmYbV31g7Vd0g/N4
Ml02rf3oi0rzZrZm8NpWOfLPBoHmMvXIaY1zu5RrRFqwRGmhGw7vrPjpQ/lMEiZi
ZeF8IgdjvJtfGoCZIjvoiwgevsIU8KZydT8bHoirr2nYTjWdy23PZwLpF7bJoRXT
xGsi0OnLevuXz9m1XZVo4J64UTgMRvfAl7CmtAOgPUfS6hHK2GtkPRB8B/MjDsQ0
rfupjlWMjvM9dgmGEC8EZJjFPHC3Tn86ryZlqqZ6kUg9rIPEBQTgYHMbQSm/nUPS
m/CjGI1QxkJ/+3U+lYrIBlYrrxIut602quV61mnpBcWEAsekY3wutJLQtTaXWjEA
6hHKD2iLQ0SGasRIS2IsjG7jf3SFtBTVhw/3vR58M85zodSaB9j/DPyu+tw+/Bup
7hLc0URXjOnhNdaCh/G4SzERUuTjJE6L/khkXk+Gr8viKCUTh66gEGgMMqnrlGPn
YceU+w9VBfpoFxEYF49MNEToVsy0NuEGfNlQvr4seo16mI7ZyIZfLFfZmpRz2l7D
M98KnYZOp/nUj3zSQaZfOWDQqweE86/lN5FcA8Q0oZzrAKGGMgaAODC9nQVN5zuJ
3tJGdaAmgQlw8bW862C5cNMC8eA5zWz5VYlCUVv2z+pvGuYz8hZUtiML+XckEQDr
qez3YEDUqXVDiPkBQ3FpLSawzMw2jT7Ds5nP0oRh20+kHKCqqFhtIkO1/E0Iufdd
i1JrhTpUdZjhsg/V7bT6khqbM/SlgJS+kV154V8C1VLWJbvBkvWCiOvZk9CmZ8kd
PsCvgdLRpH2wMgdWyVyz9DDxkHOClVn6NGOBGy2zqmFC1LLHAYr0CGn+RiqnpCba
+2EZmVWRIHs/TwzAuvDHh+71t1gvAP89VGK5VS8kYjWim3JHIRMI4714YKXHex/e
WVIsaD83oPmjaKM1Zd9HaFggOgzOf+KS/nJm+BAUVtGc+gMriwIX9fu1fz/Skva+
irHIBCMGOv3t9Ka7OC/z1VLEb/rMVup4SSa8fcuLdSn6vpWVv3rXfUg9bOZGv24D
MmlnPJl8q/9d7ahoeCQQOh0PkkeRLRZp32UfZCxN3dYLX3l/D1cLdyAWKU2Fq5+D
UoaSYE7goYlZFIcciW1kknH2YiQ4aRullHiZ7f3426b++NwwZ4F4LfIcWLxhm1WJ
3X+VU/wR2kjCrBPRYP4VfwGLTfxAUIzWEqGaq/gWFFcioW097HcoWB40b8JNLFYt
lqqD+Xmc0f2P4JgMjmI0/ETs5ZdFbmCoVx0xBwmQiVX/bNvKlZyC25I9U2EDk9Nd
WornEydk6wQrd9Haih2QUA1Lfi+JVAv8GKPPUeUIKpupTXMcQLw4Bc/9E6gNaKl1
SjwY6kSwu8etgzT3t5SWQcdwpuC+TwlYeyVxWmMFm3TQtvYM5Pw0QC40gkDJgxlV
DrLuRPxkMmvcva2aZ2dAF9e81utnmjCXESz8omoP57SSTnXFOp6Owv+MMjb2w5ZF
ar7Gdf7TtYGevCyGIJw7FJzuRgKyTUEieWbyxzsSdUqD7E4l1zcByvVfkVd+7Xjc
lIuyYlks72lpZqiTYhLtWtiMDOnzF7V0pDwIDav20aN0Dq22eRBdzFq/Qv++N431
mfgZmmSMQLexzk/eTcMeRwjRwA6w+wWnWg2GjM2H8MBtExlQJVxbtJq91ohnJ81m
489TIhhqw1y3pemQafLdVKPN06JSsbhET6RrlzFqy3Kl4ljj/pl1duPxjbuYq/FX
GE6Yv4zFW9EydvTRx3kntc/GDOuAYCDBpPzGEzHX1fDmGRoUOfCAIYeA4GZeiNDB
xAswDam+x0r60ejbZIyX3pbkJSJxidn6d5wdnHG3hNKdv6dAzVXmLgK3JFicCpyz
vnKt8nac/Y/Tefwi5972JG+Xms/a9pbKfEeR+69qZOI1RpqzsjmVd2fbwf4ojET4
GcEB6akJl+qfXjg7EDfbshUwjXdVWx6775HN0TPC75krkyoQKkNzNrl0B99e4ucj
dYXWAxLe20QBMdxUObTsGPXBNlpCMvr1hkOfgd5HqVKrGOjlBQeKm0xDso//4jDx
s30qcDn1dBaudJT1ADmBoadsnv+oRAOmYv5GsvWNFvNxfbnPQUeWqtHyX9ktSxZP
r0/P9dbIA5WdnHfoft3R2opijnEFtISQfz/ryvo/zHWOY4LpRVWoHBe3PXItMFbO
uDUvlrzFe9vtY1C5jXLotdq6oHPcAX54aIitZqtn0u87mI3QzXfPFR/fG7hbmv/A
m/ln3CpWYmeXRhZKZ40lB/QcqtSoCszajkpz/MGdE1gdhpbjJq5OHPhuR6F4uOZN
rsp5ReCf1hzU+sYdhA/2A07IBUZDH8K42E4XAH3bymQHpIZzGzFn+jr4VrWM0yFw
uflkuFiCuGP/QMW2U7pQtc3o6asi11HSL0AU+n1nN2UfJQg1pH0gK4onCMRkhUVJ
A1DKtA1H0h5b2QXkIHQ5qu2gi7dsT9RMH7n099ENHFMiJTRtiEvGrKuUMZ/ZIWdG
ZGK7SJuI3cUO7HodFVQH1YddG/jzCGZeYu2tqdDxlkjvXMjYJn5I+FxMRaa+ugOv
3Zs7U0U8/VY5WmQ9XJ5sY0RUnZOlqTAPUHke3B9JIhE/QJpXITEHdd+vN5JIOMXB
uMkBWv38rq66JsuKgrlzz6cFWI04afJgFHw2rh6I/yOOjxBEhpVk45at0dIMmQRT
R3UUCYYG5sAfawVetsxShfD/d4KwvFOztvxLSRRd/IsGN/C4bGeuDdoXTvYXuUbU
Yj19/ZqPlXRD5ShzgUZIJoH1gQ2MahMX88k+QXKhN5covHEE2fAH8G/YimVjNgqh
NaJuf8K4rA5SSF1Pk9KOCuV3BR7AP4AR5hJHr/2ydxrHoRItYLscBLU0BqSpkEym
TtV1coEGAosY1C3QCKV7Okb7IXoF7+HHPJMEVkCj0XyZxU4s80rL8RAbX5F/ac58
3cDwPrFTy8qia6JD9JBAefvgoxow6GAma54LrTswElGb0BBartzMMIbkNBw8lYNm
/FQrpVP25OOOtn9AoTLBmxUEcaqcEwXLCDZWg2oSfsDuour4wzK59NCxu9yUS/vK
7g0f+w0qsVcYJtti60aKPje4fEjOCTropUHJz0A/OLB1stAOzS/jh7IFYAQb1CcI
2MaVgEJhQTduWifI45s2WqDIu4IBKWIO5DSqOwg1/jZ1SqfSD6K3k3eDYpUK0W3k
HosDqzycZoUvl1biHkSCxBQEc9tyEyhL6T1t5/UivUc0WtsMgC47QXcuqV75WaZc
qRXCVFEI2uA5oih48yPpg8qo+o9i5rFR8Wqp50UqMAcU7wKyDpEkJvOPs3VH4guT
HQ5hrzGMaWn3/5mETwFXnGhLbT81fOMNCMP//OqGX+Rl5npB1fwSjmf+msS/+8c3
k1AqsyoJsVM/XKD/zbDk9d+uzSUeLnfq3f7+8RJgH9WAgQ8fXfXB1YIW48dMckYR
CteF/aLE1yCsYy2U5G6cNDAvOItkGpWqLJC92TGgVNiV+V7eb5o42JeMe7HuXyOx
NPOTDlxLg8GhpngUPbtQeub7xG2hrxQCc9mGEgKkMFIcH2a4zGzYEs0xVHvs4VJk
/I4TtAXU4gbYilJSyxVqvScFZ/YAnE2G5hkkH+UF43PsQujTjQNhaxTxUUmkXDos
geS7oPO6iFHOH20gahq9c2+JKrLyYfO9pnKJwjpJdkN5uJBo3d9lquwhWZ5+BZ2j
gIuSYCnSM8xLr3hHNFfgoFJd17AbZgNqz3XalqcW2pma9fx4laIqMiFAsmN3cFgr
SQ4TsQKeGOFahQ1SQ9597uLD3N0IcpxaSaQhiVbGhdT621WWBPASAFBgZnrGO0n0
iEtBm0Tx83IY2hdZRyUP6bFmxDQrCRc0KhMXuZuLXMniceMk5spHLJLEc34DwFRL
UgIav5P4vp+vbDWgwT5AA1ywavSmLGPs19Px3O5x6BwfuN87ZA7v046opA9UwswY
ydTDs4HYBqxeJ7y+79pgK3lLUZetc7IUShDGSrWYZuJ6yxoNzrPWkkvVdyfdlb4D
4e5OAYLjC8vqnsNRbyUfiwHnxu0EcOLiK6DPqT7UgZBQFZL6kEvJ3SaSrnVO+Ro/
SfxNpjh6v8Xgz66VgXXi8tZoSvEYN5rZNlrEYCcRSDycpqj1GELDZOqA/nuTuab1
x3QdICSgsm3icIjjSzD7VUU2502tHFES72Y//L6Q2P3OQj7U3FuAnlFtWLuaCGpa
iY3eadu3LkN8D7rV6U+WndDr7YUnanj8d0JkPzoSv9ISTAu2auJbuw/jc0IvLwAe
NVON8K0ArlqmQMzENgVSROCorbe3YfgtanTkkyZN0lIGuVoF2uhC7kwI9doIho3B
bmFEJlQrQrOYvYG62TU2mZEbmp5J9PXB87zdIAVcwapjH6LB2XLSDqaIgmrFxwre
8C9a+89yeXvH8bb73wLZeSz0VE1kZVVUX56s8YA23tZCkCZh68uE3LjQHCfttZ2C
ZIdBfQnk+0YxIYA3DZVAMjmnYwxk5fnh/oHsTzwzjLIk/BtehuCuIWwLlackJ2b4
JTIdYe8tFBioL0sxzlxe9qXBtVdU4tMqviHgrjUKURKi8kt4ZYJ2ko2KuyePKrtn
KBLv1VCGlFBFDlEEQHnUztaOjMcoozqSsYo/CSsK47EEvZVj2uEiFvjVpt87TwyP
b6su38wQi9d33MbWhvl4na2/+cYO2Zb1GtyzxxkRSmnpidki6Bw4ZwzVVB22GQ5+
uKz3fhZgE3twj27RWLyjzsWXuNWPLQRN95eIsFd8nRcF7EHZzacaQOPxPPWc6rMx
AKJo8WHBZEdRWerA8pJYZxWom+8+ysPg1Wvb8aS78D5Xmmz6cwPmgvcp3D5h4siE
rUASdo7PnNEON4Gk1i7tjRWreISjp7BWWrXegBp+356lYKqS1XewDPtxxnK+SqKy
g3ereItSOenLfhKM38ooxHl0CsvSZY/IxWMsNDN4kclLK6LvBtpTW0Qzr+AnumCH
KOVvLX5WPqbxweClnLpmyMfVDvua+y9qoSAjMNgLupXjcOLRGjcMobdaulbi2uN2
166EbNn2+vQpijBWNkbryfsUvnuFKoLAoRNfBe/GzaYlQzAHarrgIZWj0f2+E7Az
xl4Sh291xt66pWh31v03elWn3YPpxtPXkQOGpDq1vUbuDFU2CsXJpKljGXySRmMj
ryWNL5TvnO5ODUxaJno5UyIUqESlEvMb1XvGEe+i6twuhfJCu8I2HxH07hWk+gzw
IFeW0hFPaTyJeW4/gNNUOUXcJd9TiUJuuU6iTZkW42AmWEpaG6Q2/o157+pqp9Zc
ji4dCoRSWg+FKLcV/UDq28RSbd0Cy55MwtPL8mEuXeMLBxtUWfM89HOd2fyNRWfb
whyEvOe0Y3YFZMUIOtvR4t3GDVdhYK8Zacxtu2fOJhsfpY6N41J6MLemldxc9XQM
VS9KIa4Oc+m/zlt+31M2gU+ZbLCNuqt6W0RK8w4Km5hWnL10z1y+mq3xUc0z9Sje
kqbA4Dgtcg+IzRtfJW4STIfpSFJ/O/6HIejVK2QRo5Syessdgtew3pJDqI9dc0E8
HJTVRWamhKDMkcrFGXyGp1mC5XBv/gARAFK0hsC4UOVbHf5+klxFo8Mo5EKaY63d
mr1SoPbMKxq9UguWp5rDFcUq1MRH1gw1fg3zWDXusEKJbyWME6Fu/xE/UJy+Av72
R0PVHQ8zU0Ecm0PNJCCG6P/8ca3POWbaIYAX9uP49BTaFdqJXnvWoUfYB382/rUD
ToX6VUsFnJX2LI2/LfzCIy/aIEFu1EtfXbpjU6b+MNQKE3t8tvsf/F8GBscxaAQn
n6hqSWYZyo7udwVdHqlJEQiPEBN5HavRylJ9iM8pFGzWYY7X+NVqkzHUxx58nsXX
LAX5ofq4ev24R3JGvZlW8BgdBSKAsVRmtLlHAbt0C/aYYcJoIhe4EHD9IJ/xRLtH
kjB5YLz2/KBdDigaes1tkDgqDR5BJnr4PKibJHGeOXQU005lZeg9bgK6l8U1hJ1v
Ge+OVrPS+/0zAR4Xetk1Z8qMf/7pVXZV8jC2XdFxETNSZJ/ssjORYOB9aBT2/M8C
hjTeh/ibdp8YPAVFpOOy6SBW45Oid3/JfAu5rz0efpB7sD1yilfKppbHHi+qlrBi
U/y68hcbSXqQ7BO59gAmswe8fvV2JDPSfDMp5zhucJMTvQeqUqI70KNkRfaU8eJ/
hLT73fi/NVqtnnr/G6uV9yukX5Aqslp8V01d+BFFVVVcyW/uxs/TOFhI9Rg4ug6O
UpRI2D2aYR5qRZYD5AeHVhYkgjbQYawt0Y4H7ojKA1CeElQyYMC5moK2kStWJTJC
OE4ozqdks17i4vQZ257aHQjT68UVqhcQbVDUUE2O/Y6bODoNlsad4tF+fajI3kIf
e9yQ7S0JiyIJnDMKRHnrAOp0EwQTiAwbvfwPC1MOfrOeviLgn6kmFL1iu8+ysBgx
W2C1MR8zFFbiPIbzMVlNkXs3zKO8MIto0mh+uGsNNWcRHrXybbZrePlJbrpXn6+G
oHETEbbl/nZkCVdamMnYUSpKZTFJILe1r2wk70T2RQ+gei4r5WRII89xdZ08ilZH
t5DYoMcerfyVG+YlScTK/MGX8n7wGFzHgy0Gy+NAE4S5m7mztIXaDL6OZpOppeZS
n2Ef49mqbcA64De8H+TL0RX0fOiOJcGN4+MQVRYthpWczxpH3QB2KIkCbXkQt/zu
39szyjbJJtpTy/lPJV/vSc1BUsspbRgCJSZ0Gp8ev+spgjZLHQymrGfKlpHN/JUF
DaHWQ3h/YAqs4AW+Bqh0UsDJYekE6E0I2BFQaNg8fqLF1DmLvZs5LFcSWTvhGQ/x
0V2DJVPs5io3lNWn8OYplW2UyA6OAN2bRdBN/BmnbgHsAtyCngUnxrwmQPSv7LjX
Y20B+uQaG248IugKvpVemih3qBdVYut6AdB/fENmbbR57mPH1m1UNr/QYMm6C4PB
CzVCyRmvd2FtrRLCeU15QuWVQZiUhm6EcxFksKYwoAMmiCRsUD9DpkRTkaMdGeu2
F9UoZJ1M4xMGJ1hf5gySjpZ8/GzXnXsb3XIiZ8aKgjjVagYpdfvPAlE904SyShYv
ManL4b2TPMJC0anRjnDT/h1s6zV0gDSaoVs+92v2hp395/LmQdatAh1WdK4vlSuA
8FozZ8D5OKQjlFZiyqNbqMK5PkoEayut8GztsTLjgjKNz9bLquP+s6lpZ37LZkrN
FbFh1xwMo3pp+FQM5m1k+QnOCNlWhXRZr9VZZyGojSxa+83FUjQ8PJbVQ96abMGc
y+2zHRXrvbKHGjWyOHJwO8QPYMAb2lZRPQywd5xZKQXbxfIIhGcqTUP7mGGhELcT
vx6mPVteOInW6F+2Ag7Lo2g+iDxJ3/KY7rrBlTzWPEcTbZh49NV2SUJgci6of9Ha
ysh2XW9q7QnMHhkZ+Zapzrru2szF5Vp9vnGnsNpCiViX+IP5Ho3MdW0RkGR1nsJ9
59FtJXuEbrk3dZiqP8PamEkmDu2SMSR8SycKgUZPnc1oqiwjzjydm9VeTssHBi6j
V2wl0dtm/skoo/rm8HO9KyhQAeK4AuWHO3IhTIQpu/IpNADCDzeiBbjCwCojbDMh
fb39pHL6UG1/tkF2EE2WdNqm5R/WDSHIIbR+bVDS9AZAakg6SutOJniixJPoboBb
uLch3qxDq3593kVbZ6Xy0gcXhyjai8KEWKs6q0UiyFKrn9n0DyXqyyVS1zh0H+vZ
hY1AZgqUSGUfhn06FhxMIpEpxIY7g19nDpIjr8fEIgzmfdJyJwIGM48kteckj8Df
e4VTi9u6d3DQ/c8ddjIQXwsc5wipz1K3ZRC4hyYcya/wDIGFfBSfQRkf14nHDVEB
oH5lZmDvqSSn8qVYkcKEOHCw3hy1EZPF6DoOpLEJhYJA6KoMnO2DovuYkS0cZTaj
W2RhwxKb4xBWVhbyif4YhGWIMqRkIJqlwiyTY39CSEBGVUl85Jq3GTsivQzWoDml
t1TVzIVvxcQokEuee7I5/Rhaa5SnPhudAEvdiV22ZZUelppgoVO1IvNymLPToVvM
ed2SToCSqYkdk/NSdNnkjF1/d9eW8Sgi69ho49+QOdEKvebxhhF9ISuOWf4Pfc8L
7jZyNSXzJepTnR+2K30Ma3UNQb8aC0i4WwCP8mY5bh88gkA6T/9Wf9xoxvN09Vyh
G7OnfKH9IWbn7ukuygjS+6qKeLMxIfzcRDab58izZ2lAh0qRbwt+EdScAqUQm0fu
VykjyCCl3pP5ALSWMtlZL2eCv+87tJS0B/3UpRFLiY3Lm/MefqLgzk0RtOMLG8TX
aZegrycmbR3dujCs6Luc6nsHZNWSuzix7xAi4kUmVWw3yaAS2Gy2keb0a8Ee9h4I
iA5i9vrJKub4qjmDxhhJjOGBD9GHbTZyoUm5M18b1tNpyiB5hFBm9f6nqNZ3miA4
uxkl+0SGJ/IwikDJtt9i9zAS1cEa06znsqxhuqZ6feL5/aIqIjNYSQyqWDBWgHHI
1Z2XiJR2v1ofHO4J4S6lO+6mLiJbKZ8QF103Bu7CGFkwMQdS4VDXeathFoj/ipxu
pLCRPNk5Q0fJQojCajUwMTYNHBVzIhE7hu1bI2OJZK5bs1BZW5jGpH7sVms9JqpV
9BBDfrV6xydC/G2t8kxttNTFaeT5DRJJ6VbrW5p5JFJCzC5+0Q0xrROSaxSDk5iL
JeE2/WFI/xm0xwdTDV9mVaBd70oAEBxIqvBAlDM+eDz3NUJy9zSIHY67lBkf/7yd
S0y7MUy0hQvfkCbOgBm1HJi1CDWt9QJpS7zeHULPrNEFpDU7dJCWZ5s+5ZtZawlr
aA2zKy/AiAii3n/rK6pu+rs0wh2pd4WEE+hrwVbrdHdKjo3AMbMFFoYJSSJ8t6ax
ASJepYMz/unIGsrEMBcCuVxHUbEK1Wr+t5AOa78xGQbX4UYfkTAOYdpb3Xq/xlFZ
8o4gA888tb3f4LkDWhkIRrPGjEZM/0z83PpCO4FCS8hopusjtFjyHPKWwRbyMkDR
BuFEmFSRdGob+iigfPYyaWKakf6bV+P/UnZpzOU15zGSn/56H+mQ3b0OqKezgf/g
shB4WOORMRaKBjHKzDIuaOLGaB4KpcI01XUBi+ar/gKhkAOpRzY0kbNzGfZ/HxM3
OINJEriRDHa5BblX4fv22oBGBw9LAioGUk52ZhxwkEVpC9UMxAOzqkIxXVK6tVKX
nGkL/5jw2tfFbXoP9PRlqwB6DrFFJkbuv2CwB9Kx5yTHJjeh2XQHTlNkbu0Uzvon
uW6d75m0kRE0qfZp0FpVfL+enXIt3dhSAchvKqI7fanJC8VRk8VNo7s8OrbNFFNo
PDhGJzOpoC7Rlnr+ETuwfqKrsEkVIPVluuw6vCsjqPZrwty4/0L46VSCCtztLXAw
nM4Jcuy85RRVO54q+q2x/ApbqgOVTRAl3cV1xGu4bRK6Xi6tgtyi4ZaLIEmpVL39
GjQyR/6AmYOJmiQT/p09dMyo/60ovPe14ixHE8IdZ80Q9qYbO4WYrLTIg3zuHA60
2+5c0refU2Kweu7YDNNNhKcQbk8Kl10oJxFFcXuLxc4yG/TQChK3tlb2na0z2CmQ
FbP8hy1d3CT/76Eh3nJy20YYgL5kyDEpYIxGV3zbgED2ssDRXkoWgLs/2x0uiG43
dQIXlimYCp+A4WlOwV/DcLMzQnCci1mEeZTEAeBfDmHrhVoLPwrUaQabMpBnZvmA
cxZyHv5xpLfQhCqIx2TsfuUn6uxGHCBwipK8bJODei8PFUmtMjeDvsxlmVufnPkv
tW+8AOSvyBWTVjL+x27oDNEBy8JaKHh+9sJW+ym0HY/O/TVI0WHro6QsR9gSSZh7
JDE5eLWkvv8BqL1pRuxccxFqpTVA4rk82+aTrcBKyfziQsthGlZJsAcmMd1dfRv1
7KDNOlFKeHnB4RqBqldFc0Iz2H8jRQ97YuakIZq0IJUZ6t4TDPLrd/kPT0amUixq
M8M9P5PsoGqIXFh3/C34Ip6QuMQnj01dSMn1rhWXsjO/FcluGgUg7VUqbm7Su225
4RtWxWDCyzrMI6k7d+M1nJDQtbPdz2QL23oh10xsoUdDg9wiTg0VVdbWQAuDu1g4
fl2zKMNLLoZEDuIvk3F35Gk1R8W27c87aTDjZNOJ3ylu/KdDX+T/QA5AUrNsD2S1
0hER9QtpHAbaBEwX0ZrashfE4MVnTbQteZ+BR/4YOL92U7HX4oKjPKki5M2wJ8l7
ZukOJDUeaDezHOeAo6o8/3CioFKqeBlFnPDwdmagVEF0kA4FUaHmNl+AsGg4ZpDk
akk+e5kfbv+Q9uaxUEIOnKfjNcBkKALQEKOxNUTA8dCkTUYITDZzwtbFLf4k8+SW
9JkF/Igu4++874eFx6p44REtkwBKXaPtxS2WeY/JcwwKPTDGcxIzb5jeTSmA9H22
DW6GrWaOVl4isci1A5FBDfXXIEWaLD7sKbOkw9YpjEF6ViGl4QJZCWiFGEcOdH7R
qJTbSp/GLqt2yqsithW6kxMeuj/F9uAONAQzyKRzMMnzmrWPdlhHT/ImBNJ4dtQL
t4Z14N/6b5/s++GdtwR8hGlSE5dPrD3fCw1dd7/kNUqAoQGOv/JzjlVZeRucASMN
m5zFR5ZD0mLMmqbtve2gs2V1PZRQInWA4DUP5GpiBhLFz7DwxFO1V02mqmMsX+lr
oLMNQd2jijLpWP4FoLapltPMW7J6beGo/uCb4XeG/6TiMODQ4p5SX3pgvs+YOm47
rBS0lKD9n5sdq5gYFPWqvQAxM0FH+J4SFqZquLRjz/O/xnK1f9BS2PEfZmTjUJyM
IDIqrL+KXQSnit3z2bgmYrJkPfbTj0S1/snAdsxNBEYs/OHhfef7onndxUgLKUTO
b5NefxukOhj+HmUhJnr8rvX4HTMljVOMlnBphlGSXX4tVsSB1i9H16bXJ4S38vlO
zrNyjzxEdx6YROHuI/rcZIBHL3ThLFgHepYTOhUJhDtiHDU+0jo8oWz1ujfEZePe
OnjdbtVwTNlj/HJ2Ew97AnY3xfm6KrmmoclSRm3FO+jtXlO21wjO5Qh85LgiT6/F
F7wWGE2kgsWDWC+wuRDiRPRr+VaedxKCZYDN8arUB9FW/rsgpeUlv/bN7+sp8Rcg
W+ht4ki3jJa6XbEHAPiDUfhXxQnmUXcO33IwzSGBCjSqwZ+sSYN9VcqBcfwz/SJ4
4le+zYANDid2mo3lyXsZgW2wfvwRFV09frNEB+FLP20GlOk+NqkyR722cNnNOkwK
7Mm0x1kWTdLlSGHSGYw/1Ag9h9VOglFZ2XyyzoH5mCdsdmFyZs94Xqk6heryockK
JsKqf3JxkCsQB+izb88tklOBqa50BcQedrp8GSqEnoyh/1/edof6wL1mfHJKspq5
yarWH62P4mhMKWib/g0z9Wd0UP+/aeYTJkj0O0TeQ5/J8duwStURzU93H688Q24F
Za0YPCmAOIK/4iHJtKtVHnnqjkP161oNcVen/9oFosHP8buAnkuBNHRsY1B3pmfs
31VDSHSFBt8PG7Z94M/FwHSHEhpNZ67mykffV795Jp2j5NFSuWV8p03hLrKfBqJF
j5g58uAb9ScCIovy8gEJx9/EBwrMmfPMrCMybF8adVMP0CvXWs0OUzBX4LL0p8Xx
gZYsrxoss4dMPwNK84Cs4NutGoJFNowdzbxySk7PKbISwNc1C2xygmZImrH9JELf
YbyiOpcHCTUCYaHm+Ty1LstpuAEZPrAMc2fqS/I/mGgPdztaLYVQpZAtBRPtFLq9
bID9pPnqvQtOw2DLG2YQtEW73FvPR1U65hdR9OwgMLWsLPA2JF3jA/AWgHXr5wox
dWKk0/o+DTiRHhvDgJP4b3dAEuawh+d2B0NLbUJiDGZHKnu2GN5V06XCrZtNkQAm
H7ZY2ZRW7xtqHhMQpGLvoC5rDh4TGnB4dbJ0wWRgFzd118pgIdwdvrIxKMBD8QrB
I/sOiIaIW5pFISF8D6Cq13Y22S2ng2F3cr1zO291mAb0J0Jl4IM7bNEQ3ygqk5t4
MTpU4VyGDmBz0mrwOWkmPT9h+pN77ivqnIITCKJ7F8qwhmianzLEQVMNBCtwxbwR
en+o/hW1DXfMnc2KEJTF+eBKl9ex3s6SsSXHc6Ld7ns0BnGykqspzq9DhdCE1Gfr
aMCPKMyxM3jm3aM0dXrv577OdEOCOUvjE9hT5tGvSmW+lXXbMaRuLi7Ux96YWyGE
fhdNYifSNSw9hbHoeebrrGBo3ODJdrtBLpPqXt+vDjMzy7KHupfUfxllgrLrRfiF
FAbUTesTYL4R/oIbFC74TkAEbJyCr+KziV5+Pmf9h8HkcUj2OD5k/gwYl2Qa8pLq
fKvq+4gy174oGI1nZDdL7ALZmhAlHmq7W3e1z0LvS4k5KnI5dLHobDys8ddGZLsA
Fl0xuGTe6ift2UiZsaNZqvLGeTtvHj6+RUoFXq1qAB9nTno1czBwlhBf3dAspFum
0pC/lvheuisXjRg6PCPxY99u8yhoBingBQ9j3LBZkOyZqqZ4dE/e/Aa95oY33AL8
+nrzrDts9buLlPPXGo90mzv/dZ2MrU1tx5IdgTAbEShLTmi7IV7fIgkEj3EeaBIy
WPbVMaMHA4wY17xzBH7Pt2jTQvfEDpcdUDnLvAqOzJLlVQiBmU6FqGDtPx/2Am1N
zFVzpuZ937UevSjQILMF/rEziY3I3qbo5sPr+uICb4N20h3cVLWpvTvsbUOCewaG
JWe971g5q1vdsTu+5oHDKx+7rR8fIOt4oHv1aT4SZnUZyx26EvQ6NQlFKuxcec+B
93jBpYRnMn32dTddJAVdysjI7fNPFwrR/RCZOk2pO86SPqNLzO+j2GHIC/re7HP5
2sflapsN2pyVg+6rFuWVatGfrloQGimDCJuDb1yoSAeBMia8SU5q3Dbxx/NknLO0
r8fuo4Ievd7PHQHOQG/ljRmUdMMHtrxe2ADIxnZq51yaK+CPjGeRChqoiCqsGtLX
dmqInuWjIOM7OOKjA4q6Qazm4QseeXnFprCrc15F5/tknjPR1fx+zMQh2jQmHm52
trmvrkdHEt71FXZ9hiIzTAqmqrlXUT4sSZLQVuXvZnOTNaq/CXrvgWBQDdZhLiUm
10iTdh/5KPY72huXCmwdXewu3QHJFuaR8QryhgfcRw2vaTUJBAZtUcrtJUyFHeEu
gmteKrWZRQ/qHmI+ChcJUfQi3J6KKzhEtevNc7XoI74P9vY7j5O20gPOnF4B8Lh2
pNvOdhXID8lRUsYCCuR0B5ymJ8QhmzTVvKAOcnkgWMFIrtrhr2cmWstb7T4s8hyE
cF6TY8VT6Tozw06xzUDytkeHlUz+mlakyl2NcL5ag2OUbRm7VppbIivl+v6UeFqN
pDoAgvvt8MntcItfSNgChcFhzWZOeiJZ4M2A49qpsjwxkm5wOCpj2AHPxYDbYmjT
fjFYkHfl9rZBMD2j9m+Q7ToEbyITPmQBUpmXkxsFZmVGEuB1jRdbXcgnD55aNRHa
D8wy8/vG6X1Wp7oEkM4QaqOYRNZ0uwGBJBztr/24zIxT2LTBy1Xfejq2eeaer8O0
QHGaG95cia8aMbWWGzllztJ2DI02AfqU1sX/NBf7VU90vYtISboen1B7zCfoj3AT
GfqsgbFmh22klYaWzRwfxHw0NZYLvX/DV6qXoieAaatTmX8lF7Qdf8RGIzJuj1G2
9YFkZREv/Dp8bnVgwnlRbBM2hoRzGvvcuKbrgQwPavSTFBZwpBdup3uZEr2B7mqK
l+D4F3MV+m2eFO1MynWIAKd4eSKgpmpbVVuvH6s+mpWjDBmAWTovLiiGGTfsffj1
F7Yc5kYzQXLb3lVpRITOJvDyivLSfnSawiPa51TjaZykAyP1LuDItMdtRvTtvKxY
xesAUZAGFnpZVtjmo0dE4Frf2OM/ZsboVv4KSUPl1xwGXqLnvNTcmoMWkPXA+Qka
xNT6KlXsaOULn74CSk5gwP8/x3LuX5S0m8JV6chG6OdsiWxYBdSJzSkydhb8F23e
F2Dca2v1GqALdda0DSJQRwNMimXfwX5b3iFwMwRfyiTIT2H+2Ike8dPlCEpGjHdB
L5fbqVSfQrksg9s4uKi8TOL+pVVo4nDFDXhiAstwSGhE2fKJs2UH30TREhRaVqRz
bGNiz5IC5oryqeCNm3+reJgWS6KSIbKJ31RGxaqSB42J4aaP9CbT69qoSJbS5Pnm
fVSiG36AJ6BqKy6kwUpfr8dckwhLu2U8xg/x28Q2lHzcdMmcuGkgTEoUUc+F2+ld
RgZzkSNB5Q5gV92M74w6BAnmAuDBc6DqKbCMkxgF1cHoNP1EjEg6Kf7TCDHKgtTJ
WF+CGwYsEF9BJfrgJGm8ldfOqEiBSy0ghTINPN9F9iIkdwg5vgDpJlgh0iU+QNfx
yvHvSU8ZCV9Vnm6emPpmxWhaEAt4lxFtOz0ruy5eYtkw54E4C+GqUMMklwpt0Exo
eKqNLUb2RpIIdwwKKqH6MqJTsHsWfjkVFg2/6PdhldYlUckGtJT3cmW9HXCGt2q1
UwVHt5LQmjRrKcGYHzIzM/J8hWKSA5G7i/qAwAidu2LE/8XdAkyBzTp4hYXAdr1v
3/brppRYgp11rO8FX9cfMScbwju2bgC2tQ++rKK5gcp8RN/V6T4ibBG1wD8LozD6
/M94pILnJ4BhS4ujhmMiowSOK17gGDWk83rtDBm4gIHp7WTSYDRrn2yT6gbXq3px
2JuZhWw/KKO+b+mFmdu/+XkzKu5aXrn0FbQPWHLBEuU+dyHa+9lr7kPKInryKA9J
ZcjvSwqsvQ0RhM6bAyeE7isZIhJ8kZtthiS0H0si28mPbCPnDqyXdY+WtZrwmU21
bBgokdTxo5b9wzquubNzbz5AoL0Dt7EndLGd8rg9+3Tk42UpaNvIn3bh/7Fv3917
FVHnutV8XrPjLvrJOVoPGMTKX1YQ6mdMeR4RH7o8Bhp48ayDIyTTTqR/Nk2L8llg
nLyft3o6EHtE3b/ceiruJoIT7jTIpLzAPQxKQYbggJmTghGKfWgh91gElRAZsysB
K6W3mYGWWzBzKO7YIEYjSNSolvzaE/cmrDaN+KcAnEnDV+m+BbJLhQSRLoCReQ65
gx1iHGf5XfNAcQt3lGWayKqYuI2oQUeXn8ja6eOJmhon9E3GVHBZQiJClsJEQf46
Ae27PQrY+L0rEH2+AywLjeUNoRVYvVyFvoRPcL+DdIy3Ba9O+3ZRJEbrdjj3EhdB
nftex7E8eoglLozayqGW9EJiBOsuusbVYS5Uhxm1VrVYGSMwcb+HVgAEWmLf8JDi
SQMXTGIjUpNnRfNHLWdoKo+2hoqzWHOq9o9cmnq0ofj9sGtIYy0Vn/d+OtcGeZBw
+Zz7EUQObFAEB9WfjtLbExM/tm9BkV8zVTseAfPcXfQgT51xSck1sc/vQa0wcjKv
+gnxGYnGgdvqS1634s1AN1PUD6RZyAZy7vBbAPAupGDlbfI3WAy3ErkMgoD5KSUh
encfvuRvy27atpMjkKJTUxmDXkI54JIr6k6EM5bTIsO7QmAVfitpze8SLZkmKu3U
kt6kHUrRDJAyQJKv9cgwY/421xbA6eowc9qkYxmBaP9ih2NPsfen9hDETwsqjMUI
OiBawjbgs7P5tbaNI61CSClEiq4+Ogv/6LEtxSqgspBWuzapd5wykcbzqKn+ViKK
UOr36B+Mi0L11zPp0zGN8xqLEkdg7N7ur2/QvmSQVVUq8ReiUrXGMww3xjhFQJ6I
bFxotXYgb+8td6JyZLGTUDIS7ukyKy+/6YJpXzY+nv0LgaqR0OxJqnyKQc65iYU0
alCbJ/b1fseMA5+/t00MoKAzkA6RuTfNEgZH353nYf/rYDocZvDc4BwBBp5/s3TG
fR5DL+/49E25/UohMpLG+G6UQbMlHuy/JqWUMFqjy+djdqYwK6A3//0rhn/a7yPR
vJp8TR7qVXVIC0H3pFHt3xQuZgJRv3GSEKIcHfW5ssvpsY5RwC2bMDvtZuRy1zIs
iiRZs8KH+qabZzVyVU4erFqr0pMEBDUxcfrd1GD1ETcOiyKXrozCFrAaZh1qh7r5
fgn/pST2882X8fKS2XoW0ptc5BiArEG27bCARKS4JRH1JR1GZO8l8yQ1zhVzIFwu
NurWr2UcpRJRKquN1HX/nbpRN3RaW3K5tH1ddrJyGt1gvWhJcDDUyVHDnVOn+FHq
I7XguUd4zMQd1EZkFFwtl2/iacNR19aYpz1/P1lpBwTQ0x2TFoqlsT8Q6Ah4XE+P
w59EKE6iUgObD8+dbeYbKkxm9+N+9lcZqQ105JiUjwQGLq4xAkrGgheNOFEr6tK5
snk5MFrLfYHLeq6acWn8NnRJI0eAF67Ht0wTR8NPbmpYPTz3RspYNLebTvPEUMdG
nzihCYq4xzi9A8X1v8mF7CY4y3DadtmnobL6+MLmDNQdzLtyaPEg2XukU8ZTIPQS
RAoILV+OUAuzhp4HipbFmA0cMIZOPnNy5lFiA/BmLfoJCKV2DpMJXSXHGONJKEMx
WEBRNcULrHnsUlzngRnFc2XHiZJ8Zedh1LArLRW2+z21psd2uOCwQ/7ULxDhrtRY
YZ4gdTPCY8ouqHdSef9ucK5EhRWcDe0wZymsM7tgBHkOA7vau58eXY8TSnnL1+gm
nX0Ym96Z/r0mM0qPOPGOcr+K/fZIE0oRGk95nvOWwUHG7Zx5BFzKO1ECpz3QaMFl
nOtRPzte6oqhfAGE5UsNvgY4n67ByE9WegV1XUObacabF+JEwXIgkqfmoEzubEtG
8YZDk7Cpyj+duSJnPCSVwQ1PFPIJx5XpUZxLOfZFVb5K8VIinRDMHm3lzc5j/8pD
e2E14d0GVH1Utcydh8agGQxy9vi5fZpecpvOkvT3sHPHC7Dh5Hka2oBkG6tuI1Aa
N2ymmLPc79Xix2zIwZWeJAlDIiuKcGOT/tC3hURkgOUDgeyrOvnW/LVAnPc7VCr5
UDyXnIs5ypfa1Qnsn5V5krby/imf53O7o9Hdv5uViuG+MCjf9Xe6crswQlziRFU0
zGzajNL2fBn0czSWPzQNe0HNwHz4EKyqpart3RuoLfVW9AggvsgMoNkWNheYsN8E
25hM/eN+ZuMR/OXCfUuo42Y1IjjbpaS2S5iMUlldVlBpwbIavzWZEq9S56Zn9By+
wgJrZ2luhEMIBIy8UzbRE5g7byDwrpIrnnks++tcAMPZ7rPK/9zs9rmxjrrMk7ev
RvBQiqn5MKNYqfp8VkDKL0n4HYrl7uWGTo79liXiWaVzHvLups0FdEGIpleIoiRd
1WdMXNM3q4ONkg7gaOzlQ4KEB13NHdNSai0qpWNIQuFL2IPuDnM6LeeG9W4rN9eD
x4yrWY2W10gKXQAJWX3aFJ13ssHUpJi5stkF2yNn/CBN5zNivDX07CLLHd6QpzgP
siVBE/CMARkgT2K30qcyASkgyOvuZLWX1a4ssSszkOIWQ2MTD3LrM48zcExl/b1M
ajJwe4bsajaHWxjOfzwp8wG2n4OHYNO1/nXYG5Alj39OP/mrzAotGYqZ18UXCmR+
MzfyqEyRJCIay7B+C8jEOa2+MplGEydYijX6WGZsHq+/eX/JJ+KIrJTqvyzdMOCH
YEDD6F1CJ0aiBGJT0dqobNC+MUPWkVj6IIURSapfWMDuVyRU4SZPn2PDw8wpwmPo
7qGXo1kRCCHzv8l+XwYFqqggslPj/P2RBzkyOO8on7K+AYreGzIk0+H8sAbqZ8bT
ndylyuPOqZX3mG9GlyD2UhKociZDbmGkLi2CHSIal3hPfEshxJcsE0sgKzbFCE03
F9py5+GwextIwm/iPK1U6Z8pAcgelFvGtrnbMWpoaxp49HEBMQBlxFGSYbCbW42p
7NN6owfXcO9Kr7nk0eYla/JeKHRKt/dYZQMoQw0JDqu0N+Kev3ieun7VZMwEA0ZT
F8N6Td59vOQkEc+yjbnXmXG+a85UQ3bgQm7NR/k+ZK0RtoRVdzQIpRDCW+yJtk/i
PnbF+NW6L/hp29XLdFSWdTCo08u84tta2BIbtIrN81cZfuTryXwp4rWJZoUg1kjw
o4nyWKtlPmlYa2xmrJwVRjUdIbMvmRGzb/so+ix+cJjwzzq+3VudYbNPB4ou/E/h
Ki24fvjSvfH7lj4H/qOWVv/VqwWMxfsqn2i9zqYURT4ySEIAHA6CdBWXpne8EUim
WGrZ+widxeK0cy1oHqtJIHS9qQa5V9GrrVtfzLWo3KU96kzzmWpBNGE2i+r1LZIj
ChT2oleGmY1qYphojSV5WoW7kI6YXbJT4Q8vU+G4KfZX8ZIWzuR9AT+7hzHT8S0C
AyaoXQTeNebhE+ALnNGf5zTaRUlfmzMX7SLetZ8ARmpLfurQtF38x4fgOVrAynHn
hKnSyqoMtpJIQTKLht+s7+cEl22OgqsQYKzSOe5OxfKGhAEsdzS5bMTmUyd8CIG0
8VfsxQxxV6oNtp6W3UoR4bX6Qt55VRNDhVeW9HLmFINrw7Yj9vMCV9w1LCHYvdEM
4HbfcUMpTVXduu5kOVvuUbnRE1UXj3bunXZ3/sa+xsAxZ5lrP8/sKyzeuUKdPHNX
fu2/ZVp0TBI5oEEGuWxgmPlhbjl2hUxqrPrA/VGHpsmSgg7j+kQRRH9AgBDGyYYB
KH4b6rfHvVv8gdOTbGw2rvwmPwYYM3GnSRrRIiGBo5kdk+2BybYL83oAUsQtAyhW
IpklIlIc1RApzNp00I8qoWC+Vp+UgZ1XvhY7siM1jlCKJfaN4gjRoZlXpDgBby/8
mVObhuPEOoWqNw1TbXzTHB9ihwKIA4x2Ww+KJ3D/EMI+lZtW3zHM34HTMrlPQlRK
ucKfjrB5IQjmEBWpzjp2k5+YipyyyYr9wbpgjYxp3A+tPKhbxCABt+v/B7EcZkA3
RmA59AnXvX6UiL6M91xo6psqbljQtbyBCCQBCv4BbTBJXQVOO7SuavG7iE9DqFgI
jDEjYEESzdnbs2T3z380abAMXwLCu5u/i7IeeUHDFfSLWFeXXeouZrT7V1UugSbu
Q8m0ij9s1BE7gYBaXskLRxUVz6uEzPMK7FPiCgUzs1fcT3Vhteo1DxDwlu/LDplE
RdfPQWJRZprlA1f/0br7gl2BS9eREceCOuSh5AF7V+b3nxUXIsTJ5sGHlIea6sbv
+kNSV2LkjA7hpo4+56qwKL+7LpXwy3jx7iQ4wuhX+oRVd5g+cQ9zBFOkb/tV7MVt
+nmHU0VEbz+WNKy1ftqnEGiO53M3mZUgIvXQZhrTewRMi0DLfn1Acqw6wh7pz+i0
IDhgVLqGb448oZQFe41MZNMoyZyUXP5DV3sZsOCunwOloQI3ZlUBxqwqL9Hz89zP
uk50IaiM892oUAQKeqRw9ag/yyxvDYhnqOMHZwk3hNkLdUGsv1d/QtnqFnqLSuvf
J9lvvrRHumFOcdu25nuSqCuliUvsahWxTUVMcpPjFTRX2R7EiIbUflU2U5kMJ8Mf
l87pDhAqZ9kYKL4jj8sSGigcoXBTAp90x5bF7BdfPko0makeKPFg9uiTbGOXk8Qf
E+NxplXFFnBAUXYzLO0EakbmPXuGN4fd0vMBLTAwhnhSAmuhCqzGfFggATtEDGY8
Ib1rBs3ZbPtkz3Bibl/iVlwrSUxZm7TzHDIpsFnQKdfFV+tD5AAWZeWvsiwLUQ39
MkXd8TanuQ9RXMrcix02CFQ4fBu+7z3Ph08JCx2zThiUaH0INw3bZbezF2YpoytW
QAoZwrQo7onuGxGCQ1FKWortIWr9YILgb3oQtN2nrGHxgja/IaXbdOX2VCL7cl9G
FPUdEqlch6Mshz5okwAUDTurTTnIe/mFQTWJnY4wgnsD1G8S6dpg3HWNCS9gfGgM
KKe3NVQ6y7CQWLT++KlXXshq71xptXKT5V/1WxkVgSMdvWd1JNA8VqwUgOAQHORp
gXgUxqjZuCShKZBVWx8sICJbyq3G+08kwUk7qDEGHBbXJHBen46eX6HBx55RgjP5
+5Rxp2WV6+beq3h3WFEb80y5yLeDuaIQeckhn9koP7kJVgSlMnVqbFgzdym1wt/j
WFG3ef8i+dP+KKYgWRSYv9nS5u6DhzwYh9EZaSVIJDYnRpa2c8bLpwHCrgltxchu
5BNN3iVh8fZmtzNIgZi3dtgf3Z2YCHdbBLYPX/wFdMkd4V14l3ZqhfvgtYO1EX2m
AT/hKW0Lq1vF1wOm5MW2cedgvf2ynbGvHb7B1fWxuMLJXSn0MG19aAeAgHOWVrqd
tHzAqRfNBnHIN3QBw110d9xvOuOho+lRKbgOsKLi1KyKhgJ8pmI/W2M3ylousP7I
zMzQgsyIerbQmS6mRKg+ZPdygU5OaNLN33ANIEqp3Yw3wKwoy0TDAD2iI8h4zLzN
FRHKlehLV1qYiruUe0Emk335rRGvRzSxTJdFU75gM4Y8zKTOjtxeKRR/tOFAMo+i
VOzhGghaRskbWnBIKH9uiVf208gnzDO+tI2ZhPoLY4RSYQvp1wNWn/UHa/tQvdwQ
4EIgkhJKugr4cXJiMwOlAXmJEdzFimNP8K45H+ulGDEfpxZZKDsSEKTC8rM75SyO
b+1N7WiQZUMryiDIeKrujoj/pYnhYfv2M+wB+MFff3nSSlUGmiSL996UQAqmogRN
ItijCn1T0kzVxbVbBRfssRWJQYZHUazK6Yj0YuqNePqofjd9NaYeao4rRS1UXmyJ
pHUOiL5PFkvW26uBJ2bqAD9bj6y3ZKwMYNWcRnbs8XErBRyu715lgZqosnkJ+Zr0
d/xtL+FtGzbRWTurvYZ2wLXGKp+Pbk7f1hnHx5QKFQ8tYUhy84Yk17RYcYwOCi2+
EqsYxcezXiQSwhtoIC0laFJr8EtyV3f/h4DxNq0loxkSPwMvs45xh/NbrwaGgVoY
2aWPtBzBH9dUKpbwMeRRv9d1mn6dc7uNXPTqkCeqbSwl/CHBb7lEhP7i5bYB/PYE
tijOenZ8ccnKYQfOQJJU6oLFwQeGBwpmRu/88qTwzWnHJetwx0A5DlcNE8g8CkMR
jyBaTtR37POdWYrPn9n3uik6tNw5Jiqr62gqEt4rLpQqHXcOD2tql2JW1aDp9szX
ZdkuS+qnXGmwcIYYhtb36lR+46pT4GNDwpG9qrzSM9moU0N58Vr592B0pg/k1tUt
2h+3XQTcqN9L0VCYvLlxvfozXz2MtFg8hfA2r/M576lYvM7958eNxvABtSjlcii9
++hsu6S8QT933vmEKillMKw7UoHvT8sDAIOECL/kGYbmJBbwrVmJOrfSbTOg8gK9
Wf9sIAlzDDNgaZmBxUfCVCJkRA1Ie1+S2Ie0yr5wF6tcHe3ua8CDmMKJ7+emxtzA
WKCPizu2u95ONrLLPz7ztGfyZ/Xb3bhzeuKM6baWVYvoorvvxg4ZXVaZ6Et57BAQ
9tuQd5pwX3LnaZMoU4CNYlpoTaVqLtbeqx35pBJcAt2VkGwQibEwIuTJcZ8CUgep
xzfFDrLzeY2tqZ7WwY4MyQf8F+lKszeIayd5T9MLz0e1ylVEn/j8WUYACGYYtT6Z
6lZzbKflhq4HY4muukA4Fpo2H7aouPpGFsiZ5XqrVKSUVVZKyj8gIAaVPx8+QGFW
a027dGL853jSRxHgypeQ9Q0VuCAYOKevx2MwLwkrDAVNSgr8g5oLDdhd6Gfhd6al
LkqFkF4FaHNhVfku2+vagLTcO00S7VcpHWBfdCx/kaYRbMgJxDPZE3ojLLA3Nt97
av/qjugqbbx6tvdtgvJs+OVgMwtkzkk4FtB8BJr6/iZjOL8liDZFOF9NqvZk2zW1
2NW4BFuWEKqjmHCS1g6m4Gtksu87D0V9kFcRWqxx1+AYVFxkooDLnW8kkW083tN6
TMWlbbhFlI0pppdmiRrYMEbopefjfZVTIT9xLupAg51jj9m+cSSibXB8fuMrLx11
vwQDSv4KOBTB5F52pXxz08JvgvJEI8BlnNvLs4paX3KdiAKTdOwU/pCItVag2JG+
NjjKAc+FF6ZpisgHZmTAOPORqZt4+X7ytFviv6GKibIRHUneYSXS0+d5bAQm4cRP
KrOLuPHC9MDSqn63rE35RioCvg25qOvYCaotIv5ZMq0ImaSuSdrDdG0981l+rKB2
2U8cl3pyQuo2RHKcboA+5fkaIzIZ5aNIvnQMK7Qz/ztdUOtNoaxONUPIDTpFja5C
5/iv05eByfj3oK43hU2ldI+/7aTZFpdFhnrr4yDb1FIibHKDBzy1GlWT/pODjW8x
jYt1py5WNYNBZt7TCMpg+PCnMCYWdH1yMpwplasrPs9MYcI+AUH9CRmDPBC0i5no
1WQSciWLbSyk5IS1FMrwBiJ8pWs7Defe149dlnWHsVmPlKuq/kbuF3BqBqK/PrIT
to1jPQ6bPMSLGovpgTdVNCLVqerLx95otx4OMdKAur/tFaR6x9kx3AGkq6DFupAA
bxg28hb8qduGvJ7YDoKRq4p9/mds8bUilsD+vybVuuZzXyFdbbu3dAkqsRXK3j7T
3ERFER7DMdP9wk1jiXCOIbdFOf1UZjpKvcelkRDuKrEEGUtykKb79j/JhHi8JVid
JBdDaO9A+UkcdzZawZnlSPO+P00IJRPeagO/EdXXYtR3WQW3tb++rAv5NbGRJzvn
3AEaB5vKqFG3oiNZba0bE2zyrNMQbGgnoX9S3eXkd7iYSwaEjvgEmBmYpPBiJCFZ
kpy2BpFnHvX+7EClKDU/G1M6yCszNoF7BXrrzd/gCAeOQyDfMmzXRDLVUoh53GG7
VDwDwdrdoJKOtzlXjkGrIdAKfwvHDnYnxMrYuNcUzi8ZiTRMt9HD8MvHFj6CMAtP
EQ281aaGB37k1mN818Ks0dNdF4xDjYbj3eaSSjNp3ZvHPmYbKUxX3tPO0OFIzMgV
D/QwF8ZI0YcejpBc0aC3eGWkb0aWRHXjodufkKUzRdTgxcO2bdfR6JI1FDdnVhiH
yfII2UYEgOa+q2GfJpqicO5VDauScLpOtdFRL352b0GxfsLDlpSu7+s5X/dBVdAv
LbdgTrt4P5whIKaMq+hi+Gd2COuiy1BKg9aT5kTmkppPK4yqQ5OWv9bf67eFBfID
esbV8iHX7Z5jJdWwmH4eST/d1DLa/uDfvtUEQlJy9ARqXy//Izt8Puz2LbF+w0PM
7a1ZYa91+uQFSV3UiVcWW3hmyih4YMECygyXx4p7Se+8ru1DZ5+XCu29d6n71RuT
qYZJczEDrwPSVf2h78iC+sJ3Zy02rRdl7Yz9YvC4rBTKeOlJsr0ZTKa1kmg6QN2Q
INIRK0nx5wOtHQcyCbRX1WElBM2vDDoGSfgpQ5HOyKdYvYqAcoUWmfV77IbmlmC3
LMJeTCQVnFppY5SGyKGjG6JX/sgYEhzSCpy2TdXMJve1nRII9v4p/+ypHo/58YaO
emL+DrSlSf48N3bsWw0YYSHJEzzSSJzWSwugckZNTaSXnIgHKDo3wEQ/VPmyf4NW
R16lglPx7AWpMJacMd/vS53EcecTFW2VXGfQqV589EPlRmgr9Hv1M/AIwwYD7zAR
UOjVKlgQ0V4MDYM1kFV8vXepTN3ZelFbZ/kfOm1wF0QdZMP68+Y31fQLqT6FLgRr
zLTOMMjri6v7le87xNCtUu6hq+d9VK4wE2whEVPgqWw/AdQCn9LIDKjr9keBsnV4
NbEjmm6idTg1A2Xx5xL18l9yuR4oVmgSBzyM20gF3uYPLH1NLWsutiU+K7Li+cGo
t3zo9GXdmEMsMs9k5VY9WVooj3k4J0U4jIiIeZEB293d/rQEnlY7CTJiji4rsFLI
EBWv+ZnhXodbjjx9LZTF/rXI8iUz2CC8GpEGmct6WNArsDdD0Fqv6rAXdn0O5nk8
JIaSBWsZQ0FoDQaLlCz7NHX7idPhgwLJ3d/hgvAEp+HgsHHVo2FaKeAEexEt6Aow
2pt1gKkol0wkSnMKuvbrvCqBeVnWId7KqVDpIGFERL7uyMalKdiO9P73HNrktHbQ
PfDTNWlDxQd+25ganR9g+74cN//6SuKdtj16DSEE/WI3b2tkC+/mzCah2j6QcWqk
k/TrsIJ9ThPsrlnzWB5GnITHzEM9CVZ/SCajTvZEpKiN/6A76rBu5vRzsR2Tmyg9
QgcOWPWNLxOyHpYGW3mVeQ9FKe29aHnnQRznUIM72DyoteNE4kmWgxfkVB7ueM/1
ArfGnIrdC80s7yHleLqCKsJ7RyVsy5L4gyfSlEUN62sJV4VubcfQp+6KoiF9apfM
OSFS8Hhow71K187HiYXf+bW33I1oCdjrVdVF40Jh1Pk+4WFSg04gE4htoF/Uu9sY
oSDGqpt39B2nxlMKZxvfQQbue9aJeOrOrhK6/5OfW8SqWN4Rzxkd/rkGHwgOcZPl
QHhh7K4UEePLErSeew4nOagVOubkk64+0et1V8JyezoLWaoKVK2uv54jsyOhZ7bt
S6uOD0OxmTJY7+dxiHhxAbvkeXtPNsjsraV9+Gk8NlYobhhDb6cPFQ8ee57CBYy3
bwSv2wSBxES2q3kzjO/LYLax+vYKSlHBDL4nmYdKKuWF8BqxeaIrxrqbKhzlwwmF
DDtwrv8A8qnnJTBSeGLGSdHr5RYH7BCaWIPRn7Tt61O4jqaIwGHR/PAeHCcAK8wJ
XoCFV0ktHjpzMfntCWFmi2odsCh0q9Cp42X9swgJugUf8ntiH44lulIanCzdfdII
Gem7DVZnCqYT6K0qgBY/+jqXddpthSUvkRaOiOkN7FY9q5OQvL1K4jNb0A61Nz4T
+iz6Bpf8nrfsOZpAqo3xHMVKoYwgKuDLyo5R54gYi9+esg6GgYv70sonQwlQ4zJn
+Rybb2ZPVAKCWMCqQ9DHePEQunvzXMxWNW7hTHfNJhSzqSajHQ1CVe5WvFDjrOmJ
3RD3Zm1tjAG2UvBpmdQx85fapHUuEeAJJblwVEvSPXCf/oN7W9Ws6dAPi0+Bn/JW
xKdqHKU/oy+y5YFIxfEU2JazDRPYYQ78k12SmfF5CnlVMmdEhhuKbf6Zc1q741RZ
VWU5IZP28qnTm+blYkAKXqWAdzUZEArEwC2Q8g54D/cUm7ZrEQkmWLHEyzRkqLiw
FULi3+i3lBo6V1DtdnQugeY0OD3K9YW9Xeak1c7/YNrOYT2j4fhU/zb12ruXozxZ
5GpUnQ2jYZwDVrgKU6m9DnX0o+Zx9WpeCWrOkHUkMOY3d5LjYNxuDQXTGUpeavgy
FcYch4F1Y52Q8d19y1Z+YyRdk6JUv3iAGtmtU5/TV2Ll4EitVt+9ZAZvNWpZvnow
HGiGxFVsTWv0mCKhHxOTeY7/45yYcjji6UnRqd2OM4nRMWV+vkZQygB98IWXrj2t
C69XJo6hOBbuiPN0n/VNIAYBAZYu/ihFYEbjHBlHiAKPLot8lQi9MTxnlyFeL9Aw
s/Ym7t5f71MKILyHhxO9+2HWMakSjzs3f7w6L+1ol2AsiyG5QQ+Hmb3ToTGNVmN/
89SxsQXX1U607+h86FjNEabJ3hrKUqNWHygYV/NEFZqi9xfDtYC+atpihWdQLTTZ
ievsmW0Dh9XbKaPCz6jFVx9xOA+F9PJfKBsX6W8MlLXAnNEstLk0YTlwW+PvPc0m
uVNRvoIAVb6YkFH+9ktKZ+JBmYZ4WRPsyuLOljxhFH1Q6/I0nisTU9scy4df8fDT
AoXz7SngjuDwkMRiGeXickxWrUEbhFULZC0tQGSc5NpAxrZ1NL9oiWFkUm2W7zNe
rLDZs25xFR1O9h8yfBVV3od7/cBwieDVXE+kWIvuT3m7Wnbo/gkX1uIT6rOi9NH4
FqdZaB1JVmHNJysc6fB4HrsgDdIYyvaTYEnvR8fAjTuERtTENQOlEhqkBU+Iyl8c
p+XITfum9cqrX9kxLYWnyoo/l0tMgwswW+7ZVYQEp0tqTmHLA+rQySYRwcjgobTp
koe+KhinE+Iw9UbSG0SfTv7NK0xTXWnid4q95VAXPojJkE+nuuBDJfY0+giHZzpT
NH4ABF9i4lOidir5VCD6MKN7hb4gYzstMEmgJsOwXrtzDHXKEIIG0M4+gm9NOWP+
Bz38PrlngLE1m4LnaEQTa8ylM6pXWYpnZoEKKAFSdoyml5ciuzB4m4RxSWcuaywg
9mYcnU5hqRldsfdOp998ZNXDyr0JVgnuPztvPH9HhnY9scGam/Urfn/f9AtYgOx7
B/5qeYrycvtrAlcjItCIyEvkdlKLk/nWW6NGii/pRFznJAKJeQggjMiU/csQES0Y
NJWhzvwO8VZhXIO5P3jQHBmckMLmGAnw/6D9v5n0UqMBy7WKbVbJLxT4CQ27/dAp
FVFLPlRJtAvm2jz70hlilpOGwuX7jhsnulJ3fn37vyf2ssl9olNGHxh4vYIeJ7xx
z8PmZm5LTsuUy0kXD3zsrqWGnlq1xyTGAWCQFmupp20LCfawAEobg7EZ1ruPIYXg
yU1GFyTE5j5oPsLgGQ/z6FLyLdS1bTflmEz/nrAqqa86zRdXjwo8rTqYu5PonjU6
UgyxfNTVD4ZrGynq56mKiZXQGN4/T3UB49hjZFwMkWg2yG0P8aAEpwypsKigNhis
rf7/TmeHmzvAQQlE8XPdMpwtEuD1lRhOMOtuPc5qjQ471KnC5Qzn+Ex9fIqDSpdM
zQsDirHhykqSyfvBpoRCLEwRYHXzeNIjxTMi1FidG1V+WEAUlIVyj9rD9kNQ2Jvr
+deDmHyZB9jOEsShUhsMmY7r7FPQ2iGa1vU3Kh3PoXl49z4O6rq65CX4mN/QvMCA
/BXi+6KFWGvKW1ZUgwSw31FCe7twq4J5EqA8C0ymOFXFFDv3hk6BwPcWP6ty8+uY
2/SiipUCL2YAAaL7//QM5M0/3Rcy5adnuYmI4ZNpinCzQltuGbeMZFdNRtZIPd8L
e2WfAqQyRIs4PEA0kTC6TNGPWjWTAim3AtfAQK25c1aZS4OuaUZA8OxImre5JdbX
O2g+BK7u0P5qiakg5UU5WwLffhe3UM4mPv7kBqLuPJBapEv5G+BHokUNvsUq5WRK
vzRCXzje7me4Hcfxl38HjdkLTyEv2fjsLcL84A7WCawkR6Oc2zaBTqOnIxJbniEg
z7eekKkFTh1s+2gUvjPlSIUTwti3UQYLqR3Y+At62ZIIBB9I/ekSGi7/5kLnwGE7
FabsnOzAxMDR+9pDmK0Qunq105s0+NSECTntPCF7/nY26x9luu9Jcvh5RTP6rFXM
LdPCQB9k44kJIXBTHY74mbg4pC/3yuKcrDilG3mw48g3VT78YOCiIbYyIxcoTmEY
ZEm08lC5Csvce4a2NX6bssrhn6EZPft619l5m63AIm2szjacu4W+XsL+eosWYl+S
wZCQa1qOZdq0MyaSs+v9r7lP1mjTQZrHAg61v7I39G6Zgap7V64xVQ0qPNd3vsuo
zV8Y58tFkTgvyhFgDnrc1UnEU/3zEWrasNc87lqvMIQA7WkCTY1MgkRgoLcp4ho+
DXrnNZO6+vM9YYx7eI9Jw6wyPWisNuMGAqrvoYW+DA7nhaoZUs9vtJlPQKs5xjJ8
MRyLTthO5N1faer6IjkdisSneAlwN4tATCSyprlSvObab7ZxgFikjC1lYzBA2xKi
Plq2VBxcJ4hH0SXekucxIKtl4Owbk725u07J6MQsX5r09l8DJSwHb+Y/1XZN9p/I
UFOCsH1zcW+rIPzZf0BcRZqtjhg0dGPJOxxHVKn0ye84gRxW3kcEH2r7nMDURcTP
UwPV0EzcqydK8RWSfOeFhCk34i7KNi5a+5hU7mGmjKQ0QZWPoWp/u2e5PPXFCneR
+58RkMKuexrIc/BafgxwpY3bpI8eXVY0GUJSOCLfk2MT5aJxKLX0eLMyhBmv/ueQ
zINHS4i8qHOUUeZ8+6Ub2V0zaOaoqYZUhy2ufk1XV84pNdnED61AejuRFGSy4q20
GPhLWZn8JmjrUEo+UJoNocuLgIk+Z1aGtTDkzhC7zSBtGCBePxeNFKtFOxOwSgNH
pNORMa4XbrkUJqGf630FiYKuNFEnQbiJhwO/TIoCNZENcOsDn+ZN9ZKWDWtHFCVs
Twx9+2mD4+J85grRppM0IPjLNsJhFEjgpLLtVkWO/uT5RL8cEhoww9/KhsRsiic+
63bkH3ip4X99cuB8Fh5P6yTXLr/dVjI6HjoUbwKx38erYyNrv/kCARAD2YSbHkN6
mmic8+U0l5UdJtDqJfOz9fw/CbiJpulUlMuNmSiruQuQcBCRUfl7brv7vrpUjNf6
tTlV+IQV3OGbwP6daQm27TjDjICB6SMtGnwTrIiTaAGlqoTim10+LAvVoxe3DQPr
P0eHFxlAs4Zk6lfsV5gbkFh78qqRxt5vjU+zHJSXRMyl4x+mdYB+lvVFp60wW1dy
mmpdX3oSJKmGLQPkMU9BB39VHpgItHBsvgEVdpen6HcZuB1lj/T2hwdCCyKpT+Kl
uHbvXWO5kP5Dez+91GPHJGDgU22CywT67kP3a4rRptqsdUMK/+bRYSAoMmqVd1Oh
XbjAs3SEUwXSTx2/tqNa+0Oub26zenSl5tyy9Z/xXSYd3Xt5qw6UoTcWfXaaRtGc
r5SS2G/vNiOzR09NdkihBZLYhVv1X1pQ6R2YY1BizMXQRVW/iE0CSqMO4GXtdMwf
B+1sF0+saZJGQPyot/vmR90fdGERPSr0jHa+FKphkxuZlwV8TsPMpNr5hkoHa3Il
7gw1jDqJOZxi8gIGC4w5SUwe5aPFaufiXxt+RfVocBVOMgUA3foDvaKUO1r4lSrW
LKQku3MOzQTjUypg8iSrbPwcIgdriVK+nUOPCgosl+4rknyt3pYSDgZASMZiF+Ll
LIo+g93grYrljhCIlaDZacO0NTgP8ImiQHVk9K0YUR73Q46k/euN1m2KHmfh+Bh9
hm6wYzKiSEGseCJFOB7FwgseqmLgdrD0F/3vDeGeT5FgQDSRFl+sf2S3kHavzQO0
3TVcOmy3XUSH6itfNine+EHVMx+R5GJ8QK9LeGiNOtjiEoS/h1FuwbskAhEhPSH+
h/vYHpKFMWMMHKW4WvT3ZjVEnYuuICQEJKx257BYdRV3qh7DXRof8xc5yCnca41m
9/deD05/sydWbNslOQ+iBWTPRzpAucJ4S9tbtW4fMideWGy77+Rsv6c3hM65aypQ
PnspK1GOfKHW0HvWs98eRdM1vOfx8FTTWtohcRwH99oa0dPUVX9mPYumg9FK44F7
li1U2E09b/5LzuqpsgRUm5aC03msvN1BuXpRb03eBKOs/GGQbmeNjhlcpkRUhjB2
AZerJhcoLZIvped2ugHCYh4xqLussQZ2xJ4bmhAKwNpeHiKbfX02E28OOM7V2NAc
htkz1b6UyJy1zg+1UXaMJRRKWLdbT1x19DKuqpx1sX984f15LH6EL7oio5gU1UYt
TSiwHBiXmchmJDA/35H1LY+xgkK9I93SEPgjjLXUoK3mwqSiL2PDkK9fZfCQJU5O
bhqHZIACXj+++f2ieyexy/6SOM9Kj0FMzgtv3BZF8ZKp+VrUVWrgWkhlwI6wUoUQ
xqEbwwjWYkj/XA5YuOeu4ayf4zBSOq6q2ZKcjUhJ8DUkViDQJt12DRcO37hfuEkV
GJMcxC6VohF8yJKRYk85nkpL8KvU+USbYviJ7euiJe8Uakd0bFmc/63w10tnUiMR
V8lB/zaxGxbkTd8BCa3Fn0Z9pHT50fxk/Jl1RhylFBus7XNwgIgI3q5D08276dPC
mBZdYzJbUvI9AioY9bpT1R8BGYJ2cckfkEOxJj5A28iL3cAbY45+v5J2CzuGGQHS
y8tcxL9fIPiZaTql+KTTTzbce+FMh66sRszYZURb8Nohf2AyLHXLjksDbsWYxKHr
4pdcT9wUyPJyl5aVDFqjxMbSlGSQZbfpXVuwzMp3FaHWQTG5OOcfLteXqWqtpX8s
XG+WwBakZs7+ESpJ9HLMWTWbpsDbtgmyw8NV3hfyn65DltmY6Ocl5f8eSotFvYMF
8U7MH/j1wUOwqD6xwK6c+viJzUiz1NhqKbyIe2FuQRqe0CNb0p0jSC/r+8WKpEui
/etXyKlwO5vz4konywBuuP7ODXkyY18s27wpzkDGRglMBmLqruoz8Hsg1dVCR/In
85dWZmG+caH64w42aN8NZCKnS3ohfAwxgLD/nmAU7b00rJGUbrH5ttqUCO0xTyGe
sm98mml9H4PamEBzHKdq3zLhdw7BAbgWp/4klVOSvIgeATcpwM+bPFiI2osQP3lV
qR64G8D9QtWXORBIPBlPG67Pdh47LpC35AbWdYpXPWah92lGK0GvzE4UKFoi+S4p
cxjNo5IBDibKcUq0mimsAsbtubjy45Hg0jtD8UQ506Gop9jChSGHVLlWdHg5HtNT
YmqIIBRcssn6Hi1Zbgb/i26yiCe3LB9AYySH9icUNKujv451X5Sm+g7coVwMEJ84
P6z6UnbV5TsM03uUWva7vPEJ0TuELjwTZiQTGglsOo17PC9qgwmLthNE96epHT6o
oMoe3ZqXTPQa7t6sBBKJAKCVLEzy11GfABoqaHASASeJdqEBU6/74sn6izlmaU/Y
NjSkNRWWGGVaEPtk3XnIMJv0LfqEF42um6aP6JaVtQaTXvQaRLRR9/Y3ADtGJuZr
tnSfwQ9a3j6LBQdgcejMnFTZ8nYtgYp9qkpBrxBaa12eJo5k0PdiZvFKNsKjff5C
3iJGtPfD4Ils+wg4BZGE1LeHZV/medWXKcSBbde9zrJUbvrNVmYOHkB9ecKO5AK7
dQVvqCQ5SCX6UjOI6yuCbZmib4SOvos5i+2BYGyUMH6zJL1k1T0J4k3YipM0oJ8Q
ECBEhl0kPfEYNoEwjLauh79EuBI0ncplykCU2DYbRHa2EmuNn4qQRaDg21nVxUYZ
KV8B2HJUXtLBqxRfUYjlnbO25iOKSCY+hvLtgxrwvVQTEheL8Uken2YWMLT/HvL6
ipdW6Bm9NN9jDQMHijPT09q0PfIq4oy8BsKLD8r7HalQU6GNNr+r/jwRXdC2fmeE
v109qvsNQe0xKk1nCcxGYwOFJj2HGh/pRm+g3yPnrLc0NQkWYiCubnM3tS7K3hR1
unkD6kLV5sNxxptNls7xjk15fbQNJFEgFvIPZSUgIFFCsbqQvaNPLDwvDC2Ye0Br
qp042tWMQZF0eU3/RI6LQ6lJCNdzYlwdY811H/5v4LrMzRsH/03XVsz4u4Tt3U2j
vTe9Fh3NR38hUCaDwTCNgzoN/J3CY+lnNt4K13mF6lx5Ua1bcxwIPXE18p/J0+s+
/TE7BGsYetmjsmEde5oK6anbsQKZa5v3C9HR0vVbiAurn3gPTv0L+zVFhiF3+pS/
1hXOxlLwSRZSGmlZddqrrHeU9ESZtwvV+LiuozhmNh80ngjG/Z69BFQgBizgELJ+
JooqJO0kuxEuKb8jQ374mqgzPvM2nTkQSTNz2t6kSGp2x23NJSjGH1XjyEDgYUwG
rV3WpkOE+4+sV5OGOwEQ2zAhexd+uhN798ksU2KhY2jnpNYGYptTxTsHX4zhXPO4
gR76w1gCvO3oFOJAD45XjV9Oi7n212nEr/h6XGT5z2sRqugozBo556JOfdqDEpG3
PIfhdthy1JmH3S0vqvJlNDDkxFTz5vFte/XMCwoxDZm7pMSIajo8dXBhIw4CO+Jc
oGXRYNYVuFHRmAbsJ39+Xbrr7wSFgbozC99LNqurLWi2XfLTOPZuJHbXccDy5VTv
j/L0WQxPLFJYKawhWp81GWMB9RT4FlSgMQNqArwoNp6dK1crH632pCqfvsG96aSt
rYlbBurfdMV1IAsADfB2zbticBZxxrN+lrXaVANULMPNpMUaAx4c+yxsMc7UB8BK
BcC9GTClv2MPxUdpLe38vvw/ZPhUBVSg5vz4LV6IREr1ydZvn0p8eKwrsHUc/JW5
WkloGo1ZxP5wHPln8ohUzk6zzU+WTf/HEuPZ0ubGAyTp/cX5AWOVqVcgpUAo5tvz
Z3KMnQMUdlFSa57FnUKsBxWHQtwFT0U0GvW1EH2MLPeRZNLj7Bh2J6DUM8skrune
fjBH7nNsqgBWyvR0B54Xmjb9tLO4SjUmlSgDq5MlolACKLYi30gHJ+Ic3OQJm4wz
ToD/xixFldmYqa+808UAqt2/gQWrD9007Vo9/PVEVdvO0JFLLcL7M3z0RtJI7odw
4KzHLW6E5s5sbfYeiIYcGLUyGImHPtb0R1nOkNWYYxwpkMor73+sSFhfpmehJALI
zTJNKBNe2Q9stNc6o6L9uH3ay1yEIEr+Iff6rFYpEzMGiz+G86Y7T0IUjP9NL79u
8o6fKMBbv7bWA8CRlrke80DWKEQ6iWX3ahwdVxGHIEYOiDLFkTlsqOAUKFI7pk8y
72Te31LOEARAsDEs/U7IHGAuNzQ8dYf0G5hl8BNx8NPwMZ1VxZmSCZ+Zr9qh+yYy
s44TtfT3pIBnfQIEPhuCDFWWEplwMLWRbRkXjZYmezaG7NTRtHUc110alf1FFpdr
4R4eRRtmXiUDdJoxyaN324HG58xabIgKq6FibpRu3hYmKDP5PVsdkE0+kGdvTy6Z
v+Ic82dqC5hWQLAgehUf5jIk/em2apsLut9/3bHKXVfNp185G+6ebaPlPawB72Zt
FjjkNyl/ZagB+DatKzQtbclfBdn0f4m6zVBoc/YeULvnN7qXxnUCd+dIY471yBZ4
ztVbCFyagvjC5sFdqHzoJdALycvszNNURyzTMcC754ckMOtRNdie0dOE8yIancdC
rH3IenM/szqSWwoeOdS7bRkmWbW87UroF1PA03idYKMtHzKwztSyie2VmZwnzDq5
f+5Vk7rQpGaUYxMR2CzJS4z+npQpSP26l8WxIcgSzJqcF7m0xy4Px6DPniO4Q181
aqNKE5scURNCMTh6ZuIN7rFwXowWgx1GLFH3aMOCKxhH2vXXEAFxqC44ZUvFvViZ
wp9isylUJqo7AxTKjv4kIZCWo73dblRtKdCA7S+AOgwhV+Mm1u4ZauvHD8doYSsx
S1UN5WAkt0Uh101nQS0Gn9eCoZyY+VhryavE6ErDfKza4W/9A9P5gcg9f8qMiVjE
PpMtHZ+EnmDux4urWjYC/EYN/0o4u8bsGj4q0oYsPopu9mfb9hJZhbRMWp3oziQl
udAVuieGQrNZa3nXwbttlX1TLFc5nkq4AoftgVvgXTUo26AjK40e0rtlbf7c7arn
NYT/qzPNryBYmpBFghMpzAQjj6bTVIqwTz7C2Pmy/tPajOl1KmNCVYOJM+pax1f1
Gr6ODBGRKyDky6ZsWXXl5JwpuWxGU7JLqpOzLvifXaaZ4S/fDrdTy1mcZb7XAhA0
gk7pa3ZPuP/XRDNdAEsm/sRixll+PcVrHH8Po1b3mptsl6GzI2NB8hjc1kb/4lb0
T7ixv+5nqg+IqVTNddn5dNdlt7AE6egtNiawJUOHoO+KNMzNpwRYyeZgsktafps0
2jBt5iHj64tSr/nHJr+KpfSL7M8b8otuHeGr/6gTHaJJwewlyndRZQuNP763w09v
K7aedNv4l8tY4v9PKMChVzqAXKCY0n3YfuaXFx6p+97v3Ygoi0QcB6wWTw4UfG5J
PY2QxvgbgEhU8OvbPIPqsTkeI0gmUFE36qJrhx4gdQRUmBZ0y46kUMv/8kRrE0uA
yZYcoHsqlnPmLbPClDrHoY0h9uR9G64C7oQM64WAuL/uo8dUL7fBZedobaNpYsvV
deJ0q4rwyMFZHlFBNfRzU63tsXWEdOZYIf64J9XVwcdNYTEaoZbyXtKPd6XXSYQA
TQEwrHZsyEKNMLb0A3PQcxJvI7Mxq19CEPmiQGu3tQBrIJ1zSBQTuxYLcNo3vk2o
3zUOX0Zq5r0l0tPLSpp2UNQIvKC2HUm4n9pcPyU30FVjg/xTEjq/42fA/btRVtvZ
8LlRE2dnbt+Vfv4s+xolCD17S8ghh6ak7EHejo+6zpBTa5Wp5AybJSBWL9dCWCSx
0/dttMJIuVGUk6v5ZjbyqoCdZaDasRUzVpC7jYPxbqnNOdmedFmGKSZfRP5Kb8n+
T3zoyKt9GH2LEJEP+P1zytJ9hkhkiKscXaMw1qtIycNQI5YhUBKzNv6aLZs3Wddt
lpy+yikngKMN8pc+Fs6vDeVHd4SN5YI5MX96WErtLFekwy3u3pkwpEOwGy/yQLI1
Gg8dyfI8QPtcKyai2h92F0IZRBDPh8nxdBlvO0r81qPc93+DnDoPwSgpN8lBHcht
qdjjsTy1Al04xEnXImK77KzZexC4r/HA7Mwt8ycyp5OIRFrIuv6dnoEF2rrcml0Y
euurhAOm7V4pm3wtrRgzwmqYe+EL1FvlnA6HRK/t+FpG24hncwptu6ymfmbH4WFc
kAfDEdBpqy7IC4WP5uTFiHVVNd1s6xuEJ/ZTP762472ftRMpiyqn9SVxzJzSiiSc
lUsNoBS+HD7EgqlPVxOM1Kl97/nBnUAfqUNHU+DqDoG9op31kVFJRJ2jGr3ZoXtJ
z2sDUJD2ahn4ltSNTfh2s5DkdLGY8+JeKz2Nbs/KLD+pwq3O0uWFnk9yBKOYV/y7
FfWUYasKQeB1ubm06Nd/4EeRqrxcHJom/bq6nIj0UeUACM12jyQXcYfd7Y89d4Bt
5SoD9R1ON+k2zkvELMBUGL+nNEV6997jxIYacZgC/tuG/O6RmAJXwmYRTrNDZqfu
Z96drhudYlOUGnQqc9DFBmcX6DKqF9ivSWyrXz1dC7PhlIltVDXGA+jrKPkvbXF1
U2NSdtgudxph+blNgz8b6NJOWHGz518d23+FEjGO0azBmIii5Jsd8tCCCnmn8sGb
fXjBtlQOLYQGjoYcYq+gACGUh+xExElfKBzSJs7U/x/aIpCqGl8vMQNB8ZAztUBe
tj4zwgnUTQdS1CLTKuaI8VC2WtdkZXc86LpzcA9KIVmRHf52lsi4zns1jmn2Wwr0
qHMz+SPa4fqZmzpQ9MuU7ePW9n9GOnaN+8lEHJslDNF4Nx0tLrLvvN2hdzm81LGw
wdyeYEGtdfIG/f+ZvKioQWatSl/TH71oneB8pXtr90o4IuGZGM86sOmL9lacCX7k
56WcUIDW/2xEGfVyP2yVx1K0juOaOR5eBrjbxV6jKuxVqsOBs3ibzmYMAV723JSs
394L7pTQ8njAcflDovcMrr9GoQ3W0AZAP6EHRG9cbWt3csG/1NQea7nifZJ02Qg8
MUa6m1OBCjcr8tLaniBO/3vG5oPnB22E+JKjgLwInp7FYXb2IDkbt0d/z30PmRGm
bdgdlsx/byOauAGd84kkv9Yxvs2y0dbDB7R7UlYcb+fN4TL47k3OYNiYPSZKNDF8
79GhcaFE4xLJYq72+FvrgX/CfY+Q/mnAGgdkQD4IuG4Odn/HwmMBUtFsFlTT8wAl
t0LbMD4ysV9c7pcQJypzFcullfsy9pHdCvqA1DG/5e9qXDDiXjoaFy4b+27DJWrS
ZHOhJvA74pabPvGz5HBwulWRKqYWTa+5XX4+O7TBMRx55fDaJ8wcUgTSl9brikrW
Qy5s+d1IYQ+6A9K7I6IBuU0M7SwoPWITqNM7jQq6Bfq7vFViX06HROAKoQRzwAuO
YioATr9qafM7qOmqin4JB/INI/CIBXdRwgUnVz379wxs8xx+0P2FSQfmKs2RlYus
skeA/X+hf/sU1IQT1VDNfc6H+3hPKE0hd/LPemHAxheWlaWMyf4JNU6PrJEidiEs
AZrQMvg/HzRtOGLqDe/SQhU1qdrv3g98nO8zc3RmVk4rwgZ29EKIw/7txHXrfJbX
fvAjGxOwzodShs0MYcNjUtGJD5FuCmugRh9RYeCsdkkpVagEjgG5DudhHYUW8apu
aqlpE2gfLwEYSPsI+gVoRTT4mHVydJVXI6gsEDcYLgC5QjN11pT3Vn5V0AZy/xOd
dFrQfHC1hKZMdT4RhTZhmu1bcLJ8hSmnHM3J1ZyTbcOTjAxfoLGzXTb281tx6p4K
Ke0YIIEVYDzch3XIEibzzUGen6BQuzfZcTOiEdJowhrDghJ9t8Yy+SlbnF53uIYD
vMmsaCy00ZmDx4tXiIbuc+yL4AtBRb2trWtN9ow/Nz6N1B8frI8xEZVb9bnAqZQZ
vMlPh3CvRpcz2idcZQ880qP+3VeqqGuXfSqoyuUtksqU2Vyn1hzqXJBk8e7/f0c2
L7Hx6vv78uk239GUPLicV+skUl/KyXPu0qKW3BesB6UkYSD1gO8+5yVUnKaNvCYv
5a5Pi7PK9pDdepo1PW2HVOOuCobnSDnj15bNTqWMv9wU5ut1b3E954Z3l9ICwmU6
UZ56f0l0Uh/hlwRaTDRqR8ebMhaeaKg+ragM8baD1PDZGw2oWiWJHjtYq+gZLXy1
N/d8VQjPN3PgtXrBxAl7FYg+8sER5C084Q+1HMrdTBbM/ZqaVmbcfqIem1BdVVKs
qvcSQC2NBiuOOtSxeNN16w6LzlHnfQP3XDQ8c4nYiCjzNj483SvVxnSp2qjB8XqB
hR7I8P8SE+75vOtEeZ0112q6AMk1BiYEvorxOzkqko2pd6RrtDUZnsZz8RM3sznU
BKmhvT5X3S3Tu73J4vXPG/BknNUc8GTxCgangU7xzb0QOaKqiFyV8YqllIy55tTw
Xl6av3Y6wwx5pI5Jn6SmCGY0Mkz7cpvVqKQiRdAq8kHJBLlwCrvTqfvMoONWV8EB
68BHiiDCtDGArSIq3Ylo32+xxdUGbGl0eUqrI6wgc9oKNJPNkQ7a1Vs5znNJflyy
bVoKJDO2/Fyx/or7BxRLg5Ot9H/OWieWYmQrfkk6coZ65Nezv3KgnbGYRaXL4kMA
ce0S3EOMc97mKVt23VXOFwE83FAQ4CcT1k2k3rzD6wcEHhQFeMqgXV954GM32lY/
ZdPpU2ULMXq1bh228dft+O/8FGSHhQHdLqOUKyso911K1OCOBlpHbmjDAnH/+yZl
xkrG/E1x3ejhSxTZ/HEZVAsH+RKPzGXO7TCdcnaeXpa++IaSsh5V6cozjormTjW3
xR6vbM9C908GYarnAM98BYXRkZbUA6BrF2lGPcjdj0V1otOHrk+xDfrNGGeEd8Fd
wFuD7o+lcOJvmuY7XErbNShM0vgohhrq3DFHqomVG9JjsBeGXbjGCuYydHUVtSyB
jsQKPGLFvlJjyUmL94mMPOSj9kYu7jN6PsevELMH/KrWgdH1PTQ/2DUTrjINfYhG
l672zCEGwTqkaSYHZpDJ94gBotq1Uv/tIwaprzcT/hm3dFOZRtnnvKYFeQ94R/Nc
4HUunLdMfkAwBmJ0VC4QF0NzS6EXldadSnirD5ZNZ7hVoPmndlfuGI8EeLKpFf+D
f7TTs6b+2MV2lc9IQaVZxMioPZNASsj5Vs2d8zcTsWSluF+J+jQbnECbdNPk7V0I
/qv1hHJWr0N4cfdNXIfqD9jp47X4x4xwvMXpfb+yMfyNjQMavnftnnazgbr6YJOO
CkYn2wpLSZiOeRqfBS3tX4PPW/OoBB3RWpfU3WX9AvnpmkfsMRYo5qnqisRyVQYe
sF6mKOJQQ5OmYaTXCbEMEe1k6oL9ToN0w/yjMpUBxoWy9PqyAhdA6ONQviODy4m4
OYYT7QoIwxp344z15j/J1qbdz4KQ5Siz4Vwn27yCt03lcqik4TXblcq/ulcjBU5l
f2q9ymLUvurorMDDMC+RM7DV+rfjrPZc+mjRr3QlCPQUgfdx4s9zn1XRF/DKJdv9
NX8CJJBCfdKyjAAy7K+zRp+7daI6hNYOgTl/HHcb4reoCb9NsyQ0gYbnA6ZTBOt0
zgN+36ddo/H90ZjMz2SHBGw8U2i5W4dMzeWwJqXDiUEziXfTvB2ZHgy6eZhZZNK0
l9k0OJWFGTTDiArTTTXMyAIWXnzMOqr1uERmQhv2cI4DBgAXAq5kWZNo+sGY19cV
BlK3BIf39C3Ki+vFyNs7dYQe4kKiLLKgQdGxKtpSd6OI3u4aGH9T/x6SAXv6L76p
oXbKvl3bXDFW1sX2OcJuSjwt0LYMfKsq8NTwBvY6EeAhKh9X/IFBlFR9r3Xt0mhc
Uqx2hctm+DyWBmcEYuGVOf88guWhui3jpJlz1T30hsNsOGwSX03GqLXSTd8U150n
v83f29tg9wn5dPERzzfsGdOof+HVEa3A+sdKz/PtS4Ei3UmFlkffgLkxepzAQVzF
FrRZmAQ3kmbqomXyJEuCVD+YuiQtyvwQePUv11ZNosocm/VS237mPdZhMqXs+xqJ
tw0tcq1ShhVKeXvcysp394b2Wln7DUKNdfP9N3Ju/TQTHWGRA64ono5qOTG10/Qo
uGrmaKqIaUZEyrKRydXfcZmFQdiloZl3blLfF8JVNapCmNSn45Md/sbTr6uX46oK
ylFxHJBBTGAgh5xoj9QMc5htulObT892DxEnlPJOWGXGVVpvJI0allTLctcssWYd
EobH/fPhzRt2he5445e/+1icg09VHg+cgxHlATOWgU0WdoONPgs8pnc7H+O4/67J
KOvBbDpX6MrqMVbHfnIDiAXvyguhWLiIZGcVLO66MeLpb4I3sVJ+8j0HPbqw++JG
BJ/jSOHK67hLJVZyT5gmgaGofN7sma6m+/VT0A53MUnncHs6YBB8l/ruF0t7EAqz
Q5ouZY5WPF7q+/tJMJ9mBA6MXH1sZ6NvHZGonEOli66FF1OnklrPSKsf5I79+0/O
Il40hqEHE1xNte91oXeAheEH2kLGUgviVLoRwUx4O57BLhUNwyFZQsxp9CgrzKy5
6NEsEb10oFLrU9DIFvqbQyI0/rAtWp4nn4W4/ieFtZ+hnTScfsOfHUp/EVHYd9xI
IWb+NKTwJeyR0KqbRokaFA+bfvZLqOAFFUk1GrYFuswJOaGwy5fW+dkvF5MWRap1
9uq3XSjDWlhwF8IuIXVlCleusWG1kSbmVs+HEA1sC47wJBetoy/8yXweY5e/2JLd
PiDv6WDo4KOGOc26fAotyy2qMCpIHmgxcDGXvxPOI+5hZpX5rhz44sdY5cCCQ5Ff
cBWOJCm4kMC21rHTaRNVaVtcCKyMnrpHMkXM/x27e7W9WMEDxXa+30slIXrRswmQ
tRvW9PLRJuz3R1n1SLMek06i4qFKYxqj3PaCpO9DyMGKv0p84dm1evFaK8y3g9Tl
4CSyW3r1zLiy58rcbbfqu/8GAgu5tEnIk9/uakU8X80kV7mLdMb3z1T4LhthRz94
1TZdATbV6jyMDGbq4bbLuhewj60/nDpT1iaxrWE6s30j1Qjl/pWacjxokCs2Hmzv
JR9AoFtIwDqzXoTMJwUXhfPTaau/M/KuE5UOiBADyS972D35Neej+Dcqu12YSDdw
zhFn4EvTSnMZWKLBIMKtRSIbVc9cM3JJTN9oMrgYGoU48Q2RI72E7Pgr4eGfBTeQ
7//1qJdPb/h0baYwwnhJEfoV9vR80jrUssSB9U51NgxZSyOdqdQGnjhQCynwBARj
My/xoM7pHXh0DWHFvFdB55s6OBUzV37gm6BRZBMngrXsjaTI3RC7fonhEa679k8l
NU6IIq3OWh/UxWtTXm2tCmgBErPzivLVvxZ8sGmowE790ZoW0XwfWeBtGxltC/PG
Yl+fiF+gPxi5klHcpoeJrrqc7iRMaaNN/It2uOFAiIXM7QW/e3Ko0wscCIMnnvq8
bJrTq1GFo5Zl8RR710OerCzEQ1EMfkVYPTb2Ye2ZnNdNMYJCjmen1yBzI4F7nEYn
XJnvWQ51EP9me/6wyDlkzLkJ36Toof5vxxJhMI0uf3NqcMkR6t83C47gwL+iGNkj
dnD6ea4eDSdcI0YNS8PYq5RJGyQsZFPQr3l7TVDAtDwDmwgFpjKgzg7fHyFTDq75
xQ9IDcSvAjjVjX2H61HO7z9EZEq9LASX0Av8k3sAo9JXfGjLaRUo1qWnvua0yN6l
mgWJ3gdnv8N3ySUccJE5mz4BBc+mj5VErBMWGQMlXq0CktxwE4ZPHZuC9tpWpvj/
BkJDmzAw9Ey97dPFUlmx2eTYSDBk6r8khK9VM9qBq175aaJ2QVZ3pzkj7fFlAmU3
f8MBu7GzeltTg/rxHqtn+asRRQxfQfNMKbgr4aYSWeDcpA1Dsxf7gO+d6Z97KKPW
zCcBtvrSdOwhhueNsp+X7O2ycHZkdU2KRCZ5nOU56TFQJOLS0ZOJeQVijCSAPM4O
sx8ljAiypvYQnWYGwxdSVd2lw2t+ZO63PhwbZJqNj3QUi5U9glOEDqFw6/Alm/uT
YgNkqvIZxFHmC+e5J5fTs1wJmh+aKkpuuKBvLnjZy3L0YV4Dh8Ph64bms37kPD7T
RQ7mHtmsZsC/taKC3yp7F6alc75jnM6W3j1MUMJs9y6AsCgab9ssxe0eHpq4c50p
PYTb8T7ll4a2wVCHbr604OY+VYoh8FGWh+5taTie/jo1PxvPOEzwqhuKwEsX3Z9K
9jToY+aGXP3lJwFt/U4IpIRj6IYa8xaTKoBQv6+VIFPFqU+s7m10ebpQGzKEXekz
HpcFifdbvyNT66kI4QKxCLjELIOowrOkbi9kJ/n7eaHZE9eKk9rLy3dPg70GdH+k
/2ww/ic7AsxjApJlPsS55maQx3r6eM4YNEVJMNE0IWDqO/HHQHM4oH3LWXJ3M54v
asxFq4QAMFJ0a70vuwjfClgRPFGweSjRogbYi6Hzk03OYqWDIvrwjNaAFHWI0XUu
kUJfHj8Eym33QTv6/wq/Q/GKG9fraEqc8pN2QuqjjLvQf69aO0x4P/p02sg1IIJU
Ub1++f/c6OBiJwnLtNdYkIRtvskMREQDCWoFeYUC35wgGBi3J+H7Q/0+x8fFXG41
0AA14p+tB8Ho1xwImKnXxOWO9vaafU6GPNNaDhKpHf91IQ0ZL+d5gZs7+YxQbiWK
iCIR66M19LkKXKN6Q6xb07vBbtg42jK1DXuJ/tQjMoviNLv4n5IGjDzEF6DoBc5N
v0utzPB1rONAnRqsc19TFvNS5y3PB6BOvfrDo7XvSjPDcyW9qkLmVT0vqe/gKGGk
ECJUx/qFdIW51+v1vvHtWlppkOQ3SWDijKIfFgPmadY+a1PB/FCBtyr/7BwUNQqf
miVIVYI/BGdJY2cfNl+a+5E4fFni9xzYeDm8SrqchXnSGSPt3sSIQKIAcjrtVVVb
K9AYf3Fb+pOjbSYY293ii9Hg2XTqLZ4o5273rKe+JZRreBABAkHRQ1QfaCosKFKa
keRZ1M6zizSdWjEZy/nuwkpslkSl6mnEJN9f/ifjjUpwJ4lsFC98XokepU6pvo4j
AMhuUHp+lpl7QlHLwFXgWpvqr000+6Mru8smKk5SaJv2h0I1CBb/Oq/iMrcRYQEi
4OAG/T40UexojS7cRYKI7ReqnFXb7HYXYrT0t2CXj47JO5/qj9V+ePHg2x/rVyVa
3QusTI8XsraUdkbl0Yk/7KgjdRONwL9rCOH87MMxnT3jz9NQvrsFB68VklZSafKb
15H00rU0pOsS3VT/VttTYibFfK6HpZFo3yFuQ7nlb/I0/C37LrDkGsNeOQmSl/Yi
NnAEmT3PW4LnIEadre04qVXJ8tjTjxmqjQ6VQ7ssj7fJ1GxMSzVSMSb5EhsBqr5A
r90ZWirDGkGIQ6cVC4YWE0/HQYnSO4dWGb184w09EDCCT60Ba+DYh2KuK4Kxasx2
yNS5QoZVuyWrVHy0uQKKiwV3YiOMGreJOttzCG+nzwNdxpvuNowW5mFY4VQRjz6G
7VnYq/I/hHgxIZdJbFNOt37f8gbCOVpvccm56TPlQ1C+Pv9iFUPUwjySfmltARYW
JlloKJJhAAG88bF7WkpxUpwlgpBAgMF1ozQDwTcB69dt+9xP7ghGTuF70AyvPilV
Q58O9oXtscd/ZKt94ZEqRpWdT+DOm1lPwWk8U8QqAJ0aHquuMxsjitzcTWUuG8aA
m2wkkDg5GioDnt+FGhmkdbx3fIWWxJwWsFmzeLRUxrkUGiyjJ8APQuxrqibNyStK
qe0bkHUEbiR8urMBigy2ZX4VTHMTzAmHOwCvqVPZu2ct0JlYDmrJkRurZ84toFx1
Rn2yWy1nGw27NT2uiR6tSVftNtuEsiiib/xpq5rK+sQh73iwm4sZM58SoWcG8wCm
Uv+ZGqmf852199bcC5SPfv7p14msK2Z3Va16d5QD8TDwCde4Sx96zWyD+/ZanLuj
qZzuj+gtLycwtNicLk6rygJnfjjJxw+LY+YuYdx6uoTezjG4wqE60OiBB/EwttLL
uqaK6d7XlaXClF5YSwGWpStpfWX/wV7zh60Yd+H4g6gQW9qaBEn/V191cyaglvc6
QVtXJ/Ea2Agseqq5n46OD15xqVssGO6myPY+qe2Bhv/QO9t41usYNuC8gvzpoam2
mGE9SmpIRq/UtyyKNTZrNwNDPH3dqzwrunaW12AZP7+7iT+TNq9iOkweRggAVfbn
qKeXy2DiF0osVZXh2S0N12gzbgxmFvUJlIOrGEtX86Du1QZGKCRScDpEfRaCJfVw
JNUAvHf4H7j6lMuXNNfSs44EbZGkdtatgcnCrK4eOV+AUdX3yQUyCnQREPRzd1Yz
Nn4g/pyDzDpS0qSvCGVdO/cJyDq/NsOdmL2DGq+jYntbM6/U4IX+ATV8J94irIp9
mEjy/vdd6LdwRQay3V1eUt1PGCGP1FUcgOHF8AwXg0Y74sjUaao+q/keilridHNo
zEmkbvwMYZ46SZmHJ/I4p456gcnJTWJUotUQ62/Q1eHw4fzu5ZrtVUgBuIQUkoA1
cxHmuJjXrVU2eiA00erbUNv6B93iintm0i4o6iEM+xelH8x3RYZSQIN4npSrO4Rm
jAl4bGq+yxqfqwONw4J+2L/gHwnlb9Z8XFLU90Ows5dkbdhSxhs2wb8s/ynWKpHy
5zUqOJuV5bUuQpz0coe68QcuDdcd8+4m8P0KFg1TfqO7fJqt+dObLQYizaKFa2Os
7oBhL8b1obz4KrfZFDDJxgyNrYnyINuuUtA8rinoZswjx4NL1W8hq0R+xjL6C3YG
UyWhl8f+TMX+hr2ftvI/05+f915juPmaT/50j+kKD2Ze8Y2IMhkSeHFUjhZuoQ7s
IeEbL91Uyu5yt6BTRIrK5XlnQH1p+KQXtjEbtfujTxZBoTORVyr45R8uZGGOjXPH
mEBQ3awx8v11ZQE88aL20uMZP7DVTopsL9YO/Of7DWWbITWb0qr8YzZXdmKduz9W
N9mHXO64oT0+8ct+4omG+uSSQaIyE5k/+7g1xDBImzbiQjU/iSK+OKserRQ9pfOB
OhnQNH7MCUaPeuXe5Jt/UQeOtss7jpOYVQZQyeZ6aVHYwswSTIR5YFeifxqefkGC
/mNn2Z689wrrid7TsX/3iju5G2W/WnjxlKzxZd3sX+6oGCnaTOeUsQdWegBz+7KX
4EKHucGmrSbcIaCx1m05Ka9qW14f8gn9eG661tsZxCkWyhKpOkg+JTQiG+fz9Wlu
mkIkaVGzzF+SG/2EsAXA4B3VDRk0QwhYloqWJNzaMAp9O851e6LR9Ewu+9+sivwT
AQVkn7AmE9sfURlD+I33UBdAxh7V0MBNxDZ+rQDGv2doD5G0LTItKOKKJUYM8vzl
d3kC/8CEvT9A6vfR9Wl9MtpfUFSuJwzZYJfF29/BfLtGDut49GwAgqNZA0LlONOP
MZuggOQa0J4kAuUW2suJUQiMaNr6jDzXPvT7n8Y9EKBV/S6AY8qTUJCb5xt/pzuI
UpuxIyPNMc9JPyyI4NS5TLa7hmuwlaX6IdFwADZrUSwuo6FV7OFLTQMi4Svm4chF
iOsfImaiWkJQMyKtRXVyMq8/t2M6aO3FrARVGUASvYQnfDljmHOHekubGcNcoIKy
FTd9DB2X36Gvl+UhdSOCOgbSNPNkY9qcFYIr2SR6owcO1R55bNU12qLt1dla6u3W
SRSHMmiSTCndB9cbxD/dZfFb9rxmK74Bzrp7BsZLwihqNdZ2bSqxasSxQfIAxHZJ
AAtH+ShMyXP/GwpoIN1J0lbGDsFP3q9audRU9WhcgetrnuOwryKd2QjZnoAqPSnW
BXiV4Jsppc8PYbfT9x8ZmHz0h8fvB7LRZ/7/IO6ZJZNZrw5Z3ielQ5gjhm+jpsmS
AH7bg8q6vR757bm71cda5z0dkMnEbO9DeQIdpOARI1hccy1x/yhdFd5niOlqYJi1
AA/AsEQI2fjNrkbu85DjRz0zqKJ/CKPi27X1m5kTNPtd/yxHzEMU1v0uQOJisAaz
I++ExYmdBUZDNvE1VkmJRguCmi6ZzC4Sn9289Qyqv42Vh7Wcbkr6lY5SpNGmqryY
3W5l/DYPaZ3sjae1fyBuQPE9hyDyZcV2NuR9JTADZVa7EKmnsSe8w666qkfzOB5i
BZA4Q0vuagbO0yMle+wbHrt4b3V19aGv0g0ODh3pMCnoIFfPktkdGXFWLAhfji+h
Uca2EH9yMqvNJ1qv4XbyxoLE0biP00LYrdUlNsCwnyW8dTqw8BI6vzGk3K/eeXOl
GPcvOJvzOEaK65LmmFHj7oMK5UMdRZMGKNKnbUgL7Ry+TklzhmIFOa2+9TYGHs5f
6mnJlGA6HaEM6vgFy/0sx87AYB54l1msbtTh1gTbjwS/wOwu2Xkq8+rYhG9oJLb8
o0PicGJTbOACaEFj/8CxmLW5rwC9mcfZnv++nlZmV/bfERM/zTjYWNRhylaQi/IL
meT3nYUtbZfMPQwM7AZm3mJ7qHKjcIyI1qnA76jYQkPYUcxCuA+WV4iJ3OEMNflz
YuuVZqq+rys50bB1MueVXDoqEUrE65Clg4hmrGw6SQYQbnp/RmwWyfx1DqKo5lkF
ij9QgkotplMMCtTJfYdScr5wVQ/DZz79EovhoSAOiLu1nOwzQwlzJGmNgDANtTT+
LLvoYFDL/vtM6u+RJem/Y2Rezy+lsuUjgalExeYgGVVDszyMIRlWh9jjXr3ywYbx
Rty+4ltmUb2/G5zXtbIf13Gi6sNRKVDZ98aNYaATiLoCZ1DyXZa6t5pPpNC/6KOY
8umUtTiQ3okSlpatrtQ5Yz3rRKiP1lNPYy4E4k3NgASVNPe3xY/nbOH0R9c+7ygp
9PNTM98RWLoWNQi1zSvXeRXwhFpd92jB8ZO5tBjQOzpwtohNW0fKm1UImJlWaduz
kUtfdFK+Br85ePL8ilyDVrl62VX7doHKlwbatel8o+5vyNGTgpzzFKEnckP75R7W
n0qqZAhVdNjcvPbn9GMrd6Yoduh25ul8lFpqfYuiIttsEGyEzuxO/3orEIlHQ/kR
YnNs9ltiZ+/+Z8ybCZ5hxz2mKL+VKFAC+QXuKaJzX30s4cr+6a2GdZHgDMs0vqpc
BDQCkQC/+ePKlZo9Xv79mSGq/Bnj3uzh/Ijy3sHixD9f50+o3atkegTzZdLOiX3E
7+kZrIwum4HOzJh4NPShhJ6bDPgxRWQs0C8lhDNXoOnoE5LSzyb+swq2KJszovut
JMI7jRU8SK14T9i/WdKXZgZGZIkddz+H6gTYU1/FuCZ/UXzsKokFt9m1BSf/W2/e
+fvUcjtFvFy44duPg9ewc6LUzoT3Hnmh2a+YDUWgNrMkPXFijQxmNSgsI/LzlmlW
NZumSHeJby1hE5axjd/PGYPPSx9EdBFb5XQlUfthPismuRmN2bLGVRkxbeTPOcHZ
YipniW9VXnp3zenOoGrGUfwxHkno/MPsMBvW+C7tPGvSlKFIcUPIjUIph+xzkREx
ocHdPkw+KWW7kjzeDeDBIh/kLWt5qrqPQHN1+9pO9KVECXz3OvG61+Ujz19Bp9bZ
k7LG4V5LwGdKt30vudsgUceO5K8lu1kjs3KWFJ5Yat33Qrd/fpk/mUT/zWW2hvDT
BZN93245dtei8uddksp2OqIujcLpRLgP/KdLu8UX7fW1fIiytf8z+tGosGnygBM7
1U5lkIkIJBmsINZ3GxaN66+xTF8oNGSZ/0o0H7uEyZMvTfzBh9cWBjRZnaNDotUP
MQDTmWSrvyWzqwZy/ElahOfNPpg3+nulhOUhRHj3ovm3H10i+LzeTQMOfx0OCs77
fOSEi5jl0Ll+/tTMXaQG2MG69DQ960GlvG4SWXYoyQCtqaVnQ5MAyx0/PMoI7Hvu
cZTYPDSZ5M/U7tMV7+S27GUpjSR0RwVmK3OYPqvBQibre+wFS2PkwdtU1EuGVmxx
q4efJOofaw99nkngieqlbWzduHnLr9zGWHzzAritWmH50ZPWzPQjVt58C41X+4JR
2+7Qjvng+xdGXaheH0HKMoik/v0pys6oHaCBCwNVi8IPwqYDLMcKCP9anwbfWQ4t
hLsfi3cIa9flbk1yFjejihcIIGkkOfTAhmAnrrodfLFexjR24KXRs3sX75IHbeKl
opySxbKWZOBACEel7I/myKvYh7fQehSqo+sytJ7G2D7BUovNiIM6ryvxsws2I7N3
rn8xMjRtGxDVmKYdLKbpBsa0kVPQcXMrQ1594Xfv6JyNRaABj8aa7Yn0LxCPFk2F
dZsSbRw36ZtQIdj3Icvq8XdAPspdvqBWTJuteqJa/ZLMkpVEwkuqbjvJcKajzCuJ
zta6czIl1CcP1QXm5KQsPDXH6G8L8+tePVnNgQ6yvYnSPSk7p2FqiurmyfYaPCCk
QYiRZ1wGru50/8nc2wrRQspDRWnF+sxj8ziJXXvVYYBJdYLggUQp4Q0/ny4Wk4P+
uxH/7hq3wtdZnlMZBELUY74ilgsjq82xeKtRWMzxtmocqzZ0wbel4YwuNbw1uTt5
AP9IzRESSEpZ3VsVBDx1vFfNSRdZRGWy89pXM9PYClTGIPVt58SEm1YBsJPAOf/g
wFpVAY3NG/siOnNDDxy8GZP1jQj6hy21QO++QnUTiNG2mNl0E2dztuAp0GWjjYur
+fl4OSSQjCsEmhxZbM0MssYDh2x2bl70kqndfGw5m1o0lBpFI3XigOwV1BCgT+an
OYWh5dDymdLkOWqRl+/KK3PfNpapXqQQJvl3uO48MrFXslrpqkrzw0AL1pqiP/JN
MSV0sRLittGts0ZwVL0xPiAyZOa9FxAO1OOirGd1LLdHnrqSxiy3o1Q1Akec9YTR
CFXY5UoLGOp8mOmNU/tdbtpyxhSsb7nCZZwP/iKzmcxAl3lYAJlCoLzQkHlV2r70
/tFDHw83jP4u9b9RYtau1xDW0VQK9ERWctDpkFiUTEkcdzV8TFQcstbGhQYz0QOf
ui4MDOcfbHI7hv/x0uTn9LOpge0eo0j0hKwqWyNNXPVvbM8YVHBxd4EtQMzyx8cC
gtgkr69e6obBKbuvtNTPgUiMffWceNiMl6whuXR2oeuwIKByjPRq8KJAt1RVWWOB
yOUuLKK18afs9LPOdBx0kDP8WS9RdQYpD8Z22YytkU8bEhIzMNUnVEkydgy+kBx8
CveuXABIRAqne1gUgy0wZVj3oJfFMRGSm6X4S9JUY0MV9hEu86Vou5F96YKbStBr
1rnT+wKui30lao6hpmVVEZgvyje4TKKSYcaf/cUKKm0zDloJYxidNjswygI09mQu
7ytpyUakOP8sAYqxaENFJVIEEuwSDniazzTvEf6+jn0Iy2rRntWj5uO8ITIO1ElT
YrZYTzI06hV06tE88I3zSw36XPU7owyuy8K34aRCub/PBItLJTAuxVNVMkzlhnQ2
Jel9ZxPIXy3kXh1lBNxxbGWHIYnEmmn/ZMMULkcJUPnHetUv+BOy4jA/EIXSwK+E
r0u0pG7Ufk3Npft092xO4Md1uZV43UK5HDICH8Csg+svK0E4TIAmDzYE3/JvhzTa
yoCV5ngRuytLPCkJoi+vwgPcfcytxV5eudrWbJCS4mJL2Sq0NJDz7/68g+A7MuoQ
zHNEbrhYywy/OFwvbKTwx2tvi4yK6T/qQTgABkwA8SLEx6Mdw/mJ+Xv4s0pXrbCe
SG5jHfkWjFMms4JtCqeaa9fIeiNapt4QeLsnf7hHJrrytpCmpF68C3+ffZ/yQ71X
sUNsAsQeYqY+pD2QpUDZcq2VTJxMIJ4ZQ0wZeZcfSMar0mf2pk0Lv5iu9J0uObER
0gQYXZMkNQs2s2VBOlM6a+Zz7yNA5H3EavYuTEXv+lEUDmAZB4WLjC09Fpo/McgN
mJyDO+2ESDY7JyybUcJsB3W8b8O+Nzu1OxBQJyiTzGnWZcoT9WSa7nEp+pXWh3bV
MIYD7bHi9vUv57SxcZ91xEH60mJR8M6Ln9Is1LM5Zq67nmTBP0tyi3WaaOhcwGj+
pGnRrYey+rIlpmIQqCLboBw9nCFKEpFghozcuusoWU6UnNf3Cr7Qb+9Tl7p1Vae4
ZnzLfg+mEIGVX6T0dbPQgCp2EpldqWXoqBbpveJTVgbiZEHFuLpojVGDGGkWcU/s
XI+TlpdWpyFGmm7Hn+3OeRTfZemNq1P8fjuhZkWwfK000A4V98xf1F7tMtwjjSgi
+ubChacevDQSAiIFvTRVHfXj0nuwmeuust6l0RfnwZfe5uhKZ1z0oYuzsZSYrnNI
A0QyXctmGWYE93eRScs5YhYhhfeeq8dNbAyBWd+RJkvi5eZyYQ39uyhW4kGCmr1z
3xSTe79OUy4XmvSdzd/vbQqwYFNMX70ZpIgYtLG17tUGWtKBEEPwi+pTec0xe7EQ
LCTpmJVhbtZrQ8DOdSC8E26FhtivaQnsj5/OY/Pdn/r/wfgjCtrMQL4s1Y0nyQTg
sZ4gDRD5KLxue9oBCP882lMhM3li5orp00EYTkVOrjjFTmhU/75U1hbUqiPoF2w0
AzIwabwrb/uxmvxKCQy0vU+uvI06wZI4rVkdRdRFV0p0V0IAGYNZSb1C4cXFGDcj
5J+KftjwTnshy2JsiR2vWPd4B4u9Ae3LN5NA6xMcThOLFxDRoHcEo4kLLCzivpK9
i/dFuzaORHyf8QvXcYMmojdNpH83Zyb4n1B2YaGKrnuckZt8cBHr6TBFr4o5bHvD
q+3ldNMZM+r597am2vmNny0M2BgPaK2MsAWsLOGkN0ZWGD07Y3OZ7rS4VsoQ3VqD
Px3OHAdpvlYuBEO2i7WK2fA2aTn+/Q2T3ysMnRwRrMPXgwahxotpjf3wI+ebLkgT
nauCl2g3LC+xcl5n3htZtgjtviMISm7tWwWAU+PyvRL4XkG7MHwvFM/UXB2pK9oo
qohnviUC2zpPhxZ71wn9xZFUTbEapJ2qgDZTum8dMMPLm/0lwXx0pV4DThkdCBVc
Dx1WJY5oZqzNbDBlYYoK8CwsXN+FJObjo7lH8TmREVuyJjTndjx9WBvz/kSnGH+D
o3m38by2jrAXXv/8EomAmlJvkdSsp4vWKvnbVx2dOVhSAbhAgq/e00MxIE8LHqNV
J8QFc+OOKDaZeaODD79IZM5UAimpxZdm7/2hIoUNDKAZFcKMEJg5PKUhVbhIOaPR
+oZofSEInpycq74iTOBacPAc9QcInvJtAFw+e776FX2ffo/c64S0KTChGORtd3Nc
eMN8QgbEXbNqbX0ZUgVW58Cl6OWYM4MFT2beO2Wk2Ry48F3nW4x2wmE4skNwUTWP
BrhGOzUTiN8Nsa2VeegmZJE7rpOn5OI/XhC++DKCM+M/A9EwUnFaXmbNMSeYNVJ8
5feF7R40l1K0Ubg2YAsv59pLRLcLt+3i+n1IHuXXOrF0Uzr6IRmOPDsj4QbT/9ty
45WkOXvxjtMQwIqn2XHlVI7Je6y9UeGH9ysubLbjjbHLyRmaInhodB+sHhe5Vig8
dg5gCCUyIz09ut7g8pOp8lkFLdzdy0mADbsfW0ZG13jDwXqOXE7FJuiB4tyDIV9E
fuYDFBf1B2R1lS5UD2eNBmEynQ2cAp7KofOgh9JExIasPpTa7llpkeDNaASmzQSn
ZVWfZ54kRD3/iYzVITK7Wc3pME77SHgg2/18jinHi9MvSLILkwYAaVbkUqL63sU6
78Pc8+6tNixcvmQkETqZgF0NmmFJDpLJ8sPS6tP9+KkBfQIZ95ASIeccudR9TOCA
AqCRwN8M/VC2xy9ikBbGpBBrnf0s5A7ww0loR1oSH1mlJJHE2h3NXzqDJ6n/Lxqc
KON2IUgG27kDAL8vOEK8p+rLUGVYLwzvzyMMa7b8d+5FWX2PAyjlZZHwsz6nkpQO
Bdaa2WxWeheu22hYv2tYkEAFVZUaKVhGyc6UGCLCcvVe3Sl8MHRF+LPs1Gy/W8fq
mduQMP4tWqBGmOlWWY2uxdDUit1IAAH+bs8Lt65YH4tN76/SLsIteFjm+zlAFGxm
/aONLV22uwlKsTtOJD7dRhAUNJqSLnD5sxzYipIRqMhwg3qQ0fIZCkepUTcg39Dx
fvukBgfquQXs7O+LDD5W6fj9To3FglCFwAJwR7mmS2lCMLoPEw3Wqpx5fxJq5aFj
Y+EmBTu5jA/13UNTKQHr2V4ZYraQmqPoLZlAgP/StGz98EeWnyzkUW+T8Z6qH3Uz
I8bR00ppEFhsJ8ZPLs2nqXuCqHYlpIusl0WHFFjRiRRdBfvZpzQ0WP5wdk61gyHc
Iz2vH1LMWmfDqSv5s91J1txXGCueBLb4l/OODSNSXUvSXRPiHJRcj9AR/FmONs+X
yocy4//me+lyJdrtncKyMMgZmy44BBPJwcn3XydpbG73RpI774e8tF2w+ELY3MQc
AtjrzDapWkoLA283yxdY9gCcWl/ftNRe+pa3lxn2DXgO1E2T3p4bjWP4V960wJCN
141499VHyz7L5djY+fzVYhq82dMLAapgVPndNoUOVAFUIjvr9i47tPIlu1yXps+A
JaNCAmyet/MiP0XwNAUPn0ZeQz1sBMEF8uDl3H7wUKAlSDfCbyHvmRcLQuhHNPaF
bWFvk2g0kSD/yykrNf3G7kjcL7wu2HIPYiQ6vWEXUNnTFZsj0zKFiBxtWOjiveH9
kbKzFY4cy1TZfq/a+1siIrQcyg76wpq020Zb5WtUVHsSRlF4n7ELekFWRQ7Q7qUJ
wve6xtX3fyrEGe5JjAxkdoQbum5BdTPUIucQSuv2nwFvocHWkx6bbn8efzPmTkCr
ir/zqYdwWZuk4Q46Wsr44emfzHYQJQvY/l6KFFTyAnxUzgc6ExEqFe0NM7GTVcxX
KfCDUuxGvI5AXBfQDbD45HBH4xIPKxi5fJDSFcX1u6xmVJYVDVGAOQ/ari5PbSyJ
P32JOtHuwMQQsJxGw9RVhrGoa4RIorg6XXFWnGGgOztQCZ0N5ASmK/HVhq90AEiC
JOFW2Tp91UJTvYHG6jzKbrdznHjwOnO+kBGgtPqirT2JtIRJ3ZQmIfpUPuyTKWRo
Z5YMKMLpKyFNkUGLNgn4ONRYPUeONH46Xi3DR+2Gcutkoyt3vRJqOYfWSIPJE2dO
lu9SBQyKVuV5epuLf/meaipdo3FPjpmvaZCr7Q71sIU106e3vdkVBX5YQ+pRLmUJ
WRRbcZ1WqbrmgG1r/duVF1cGd2k+cX5pE2toUVuBYrhMEGE+sjkqk65u6AcL7Zju
PnOa1PAnkix5iCpcIGgsAVt75vQAyH8RwZbIwQ5AHJYSLHsU9RzmwvP1LUX0Qajk
YfRo9deBxZxVeoarmYnwWqD+1cXWSQaD3wZUHOYM5RpIyAzhw1yeLPeE012YKWjA
cp6kY5jqAhNONwODtO1mQBVoJPm2aWT9UtOB1n7uw+ZtYfiXpKsKsDsM3BsufLix
Gq/6zxoXYIYDKBe0oj+wAnQhGDX2c8X31uF1iGdFtS8vLF4Fv4iAG5ilg9e6khI9
+z3V+7BjpZch4FPAxx2KTWaZ2vlP7tZmu5LdVYgxtZDMRwVkpQFEfoHvqW87rIfj
IO2mGcKTjgtVs+W7Pb3PqWqmTnNJzbsCQhjcYt4KNh2qaI+N1C8dUerkKLOAAP0R
z9F7nG8FWWEs0CWSQw30uvGE8Ra9dQWaFeEaKwPeJKKCIrxWO2SbH0Oh1/fyG08L
dZMw56VJoGfRXf9E63GQ/2q+SLSlxmqyL6jihv3WDBPpTeplGVCXqA/erQvFP1UU
Js+tfGjCQ52h3Sexd58CvJShdBg4OcWi+gA6FoEglMfHZvQ85EGINMQ4Y36Up4mB
4WO9BJh+gyEhRYNwtm1hDvCKDJujK3hwk6Rdms9Q4yISK7LZE5PeSqmo2PIhAt1U
uqyhShVEY1/HtHVQfCnuZaKCia4XsBpfFw6TQ0MOH+xrAzaqW41m9+JyXmK1bwFd
WjE+AzD3lP/rOhNA1PhjeSLhhXgRre4hNowUXIhSGm39i7SWTFDGh8bpDTlCQs34
kYeat2PsF9fJgaGrKedw2d01nJAbyPdm/NtlDkiU+G+/QjyItFBgvqXaipOoRIMe
wABrQ3EXdZQ1fC1sA3TOgfFquPd3mXYkg6rJG/R1OydOtG7dAEpzaW2ElqaPu8H7
/H8jLI+ILOGfFGmqFqcxvXuvXha6jzSYNaefcmH6OYBs7tgfl72dUqfbU/4Tt+tt
d4RFAoqakMYi/gx65Ts68vrDAtwL6D0rAffDE6JH51cVfbHjjo3zD8p58Mjxz7zq
J3B+0XTCbUSm/0Uw9dqPQmeJY4XRGqgSSLBZxij+0HscTQV3Hmy4NMBEqGnJCLLf
7q24YHM55IxOzH8ot6t2F8kNk8JRje1tK4MqeC+mWoUpQCD0/6oiAh9PooO5R84D
SPc4uWQODMkkEk/rqoUu2JvRGJpeDHHPWBsNctyHM9eNR2UXSIcQeOO0M50zwhUC
tVYi8ChKebu6gxcFNj4ZgfgHctB8X9eXD/rvlui7ynlaS5xCyamRSIW9A72o2Apn
tqm5aknSdqWzrDSQQUDhacozYdSJNBsMESwJ5q8C+4VM39mbtFR998R99bd8qLO0
E9LWithO1/EPhAC0GDya0/ym29PwtG1Yg+t9KoTmHHgi9e3XxEbspAMWZklkzStV
XNPKeT2xUlvGBNQUUhJOmXbBPhnU66umJMKsm3iNChHp4Bi8V8t1a9wxyK0om0dX
ZwSCiRzSBEnXJjJKHBFQk5qiZi/Z/J5WwzdaTGmNccmKSyACK89JNWoHlzdrPBGE
vaF3aYCbspNVJ6FNjG0AUK7d5THrcgIJ6VNc4bwp5pNt57hDj8mG/p98RlZxxWyI
kwhhOZZUr+9x6Yl95J9dM7W6S6YhNFJ2acfBICyDaRoANi5NlqmyxE7fkEipDcYx
y5QT4yJbngZAXSzpx6Ah7BLZOkHLHhffNbLnb/0dCBp8uXj+4+r33hrn/l6GMCD+
fTsh8W7c9UaLcVjmfmkkw7XDVdELJCdmMbnq08u53vAzkNE8bVHuEYFl/HenJmEm
UZZFNBOeU3tbQUDjnSxDggfRw3D32tIaOKq1t8SigMfGPk3M+xvNs6rY+Bk5Wv6l
TSfbgt6UQJ0kVsh2gg7i2KaPMaUotqMnXxXxG2rZQGKkUTbM+RWPjZ3wbPFsBA9Y
TYVyCSY0lyPNN1ktjdWTw7i+z/gq5snbSqH4XubMWVZGJ4k1fQR4q7Xpb3gugMtO
LKWm4MHqWs5exZ0UwICQYiyKaeoDvGFesv2JQBRxJHr52M38PfNmhTkDj6vEI9gq
BznYUMsaohoyeNRS8nm3mJ2E6/3xiLAJP2zyy5xO4o9euK+Z+wNEOjI2Ag3qZ0lk
+m88lTDal6JxJ6OUuVEa2uppAGRFQ9ZarwIjXr70885+au7ciIe43tODjtWlofoX
Eflc1fbWJdqrqsQMrJWf4YH+GGuqD5GkiiUO0Io/auWoyYHaOlMQrOXi3JF1Pms1
PcQgrX7KwdFbLXUtbU5yjGQvhZRSPntuxgxbuOolbSFY+LGcM5b55ceVd4uvP0Xe
DdMMNIeYikdKA8X/ybKm51jQmF9aoqYJMbVlN5RuJ6yY+LoYO19qfkbb3Eom78gR
8CuHb3OeOAo+VlfNJ9wgD4arLlactBkHe1jU27dsSus/4i8K6D+M5ePrdTZl4C75
5CAVLuEzmPMWWfw5RUjACdIzF4sQbNc+fotNZ2o6skO+ng6JTbqNHqclk8jYuRrr
EAtf7wNMmNEiu9Y9njBy7dcmO7khmD6C6R/ayhy8U+ZQuXvSmK6tliTG9CQwp39I
PaLRMnUmTIfrL1St7bPusGLGKg/4lJbOCVxaxLOFYqa7ipsG8q80RjHipyOPaPXP
JItffdLpBQ7a9qQW2pS+kccwTffwlzmjwPye2BOE3ayZ6Bz/zN/1/DduUTo3T6Py
hTEz73hODYA6CmHSvIW+Edl7bBgcu2hpUqB+mjeqLkS1E24KNxtw6zGhUSLlivaP
bGX9jXTVG8ucHrMfYKchT+E367/UL1Eh9gY9iRdI4dXaCMUlhQvHfJX9TTCQiy2+
mYNhTiJ9Kj7wBFvVni5KhvipmqwkJ0WGek6Y3EVcxuubPoxm6GvhKNI8r4+P35St
P/sxphdAfZ7Nx+1chprTcB54pVLyWxaVtjCmsG5fqBk1sOs6TrseTFCSfZ8Rf+/T
I43jJ4e4t76lvC9X1IRRWfD8eUKZ6+jrQ75rddWMUb1y2hQ5KHEIhZdz0skjWZkX
S1Sjh28pzwJyk2OPGFqRh3jv/kY9OksdLKHn7BGw6WTXH5k2VwOwPKBR2veHF5DR
IsPRTWn2xmSlBlsDRBJE6laL/vF76Mp17vH9C7DxqALYZExLdDybQCKOFKd5dStt
LrbehG5dCjEUCUAo8VI/J9YdbS74QXWW6GHBAbDMuwbISFnicqgbVw9eJwTMUOcm
AKrusE1MZ5O1HcH0Fx9eH3DTE19iKaOU3s6ujWL9yC14c7PySRLtAzdgpGVah27V
ARHIvLPx/KhIlHyiMiBrgpjVqPlnsGmNpJZwYBLBTe7J2bSPlbZP7lKWacvpyhH/
rKE0nARpEKsBiqHp9TwdenT6gJ106gGlmpznmMNGIGSuFzrrDSG2cB2uJKDeY6Vm
mEo6hDP4QNfknTToKa/cdBo8r5jC89xXT4rdirFHYew3oJxZCD0gzp9VYS2+ck1W
einXfBXCrjtogHrbdFd8uAdKaVwkuSn5ZDVXOTdyxgFBnyMqQ+8Rq+lRP/uR/kOp
nPZq++foWt/u7bMXHTQehtJTdvas/jLNOgB87fQJ+9sR9Tk9yafUC7vOlGXU/Nf0
An8/yOekfmC4Sz2cxUso2m+kF3MewG0DNaFhakpqTc2jdFh54WjyCbSH26HGrMOD
mpdLcu9JZaaheO93zLtTzEKVywFkzwMbN21ngjYN5TIKjryRqiXuTxnh2nzdzBvd
bYHXyWPfPW+byfnTBovb40EVix4s1JlPg6i0/glfj3rwMZzR3vo8aXsmXSgpjvlo
xZ8INI0rFmm+SLJBlB150wfjOZ1utmRinBuzbMSYu6XcKFSZbRMqD/zhD5cZCRyU
JgmTAej6fjxkMXN0nE59TaTCLEmGE7xaJ5Yi4PJUqxBFxLeNaD8dcqVNFOt5+Uya
X5l8X3wPtrkHa1P1GjXv+d+yD2cPOEm5ZmE6AV0FGdcGCVCEWpOCtelUHacA19eS
xR5DtLb3fuj0agrEg1yEtliAtC/38Ldrh9IGwSRghlOVKt1si1X/sgrotk94gqLU
80WOUj6OtdjTGxkz7oSQ1k7P+TfdpFsZXMB1V2ilPB/06R4zVxCDSf4W4oImjUJx
4uGueIt8VqzRAp4HKnmKdCfUg/FR/+mO1ZbFAuWVjy7jrG5qZtS4DhFWXwe/O7lC
4WwX2RVUkDtxWA7KPQTRPNuMuCpdQixeGURtWQV1CL7gpmXMi3p0YW9gclRsGCn+
CGBPjljbg3L6rLIokxEHs9PRKP2CK3PiafBAA4ajyj6+zYCOKN0Tqf1CAjpdhKG4
NGmzH6ZvGQm05KwaxARlb5Nih3jjqILzCmYkPQj843vaFtustyDBEZJrHUY5yCVr
EVIlLI/lLY5DZKpfE0nY8x53QL48hyyIt04FH3tRiOBPJbNSsHNAple04Xlad4/A
xiFLyKzK9tJu36H1tY8L1FAxDOb26U7kC+F5nt88apyqYUYc2PwfYKQV20rHZwVU
zimrEhFkBQKPE3utFi5neKqlZ5k8bP5LwDVhssDqXbd5AxUpc9i7me3PCl+JHCL/
HXS3xZe2VEoUlfSTZPuMIF7vgOXloZLhajJrDvTycRG0+ba6IJUOoHETSfDjFeDE
/j1kL3EwX7+VLLX1CGFx0h/5XiaWT5zQMyqn/ne2idx+S5yCr99c/2JUOfCDnDNS
VoiReR3tKZSC3P4W7JLHhc3jUs140wBFNE6R4klZ13wQWRE7shTXrpoPJle5LvJB
53p6tMBbB400JVows2cRtnJtMfxbvrmTghL0KuMvvYWKJC9Kg73971tgH/uowujW
UOla/jv/sfDk4KIJb811cFOzTxdhllStP9ov3r3ddesrRKmC7vuZLdQO+OejEy+k
4t96zkypUDW45CpNWmRakoA6BODx2Aa+2ZwnK4t+KZqEoqr0U2RR+HthBG8BttMJ
EYC3SE63WOC5TPcML+QrKGT2Mm6LEC+rFKSSeIg8YjP0hQOFM49fE1wufzVF+8X3
TXPnECJcCi/1PsLPMshw2rwEIq8OYF1bn8NG1KUfAfjxc1GbUqzx4BQeR96URm0o
+WS4LE7qiwDxbMf5cZWW1QzD2xGqvrFQrCdvgZa5avZ1na5oUwmBvaeBZ+KB+GYU
bl4HhQbPU58rlFpB7fTqm2UTx8mj2OXSK6ttVlU5L6JVWE7NcHRkpEXOrvgn/8PH
Jy+hPoNHhJqojfTJmvELOMr4F/AGuEhQ3eRYxJOa/luWZGexXbpi2w5Elb9OFJ69
1o1560iQZevfwzABqprMD6IAwtd146hM6LnWvHmQYAYrGlROxffJ9/P9b6r0LpSP
/i3gXAqBhGL+JFyB/KpmsHhdZkLA/c1bPLnIw4wMA6/rVTi6u3jwSsptLmgUUoHR
sUBXaHtS3CGnc5yjm5Nj8EjkrIB0ViPyGAiO3swh85KmP1elck326ULoCOQtizzX
eVAhQLPZK4OXib1wkK4ZgwYsXJ4P0nQHYBdwCx3Ov9gAg9bEiKfLIlDzKbbi6MZN
eMhZoYQgaVKrTOEJ+iir1chCT8kTHsysgATivZei+uBR7XlSscIFFFibw8mawcSU
v/3J7p98AJw+Pecejd37HxSGzJdxB2xVLO/5WC8fOSrJUqt3grQBTF+SGmCODljZ
5fuqYXL0Alh5kTq7OH7O1pFQJZLTl7TYKWag8lFvBhNp3ohOLztpjOL/IiLN8HMq
rld7yBfTDmDtM3Gr01vJhWWYvyrbzVPYk6LLxMCgX0U0i0qjh5hahw+AQQJmNs7/
hpjQagMpWxzGpCvqKPPgJcfKZkzz9GpmLDKiW+uAKLr1G4Sv8iy8osWlKtmPsllC
Bc5efCQjJIwEWcwFz/uJ3o7gQLjGOW0UNl1piJn0QLrzlqf8YnqF0FjviJyfQXb4
n5msozcX1vu91tbOM+9AA49doPqCJeLC0goz7UEykhc1pbEeNzxSjSerrQVwh9m+
NJ4WANhmdPFILlPaAH0g7bpLBa4T1I6VVs67kTy8kCV1joM0Dq69rjEWXSQuusm4
QWr2/R/Hag2TD3RRoLzXfOnouxAlDbT/54FQDNTBCZjAxKNohWhmwJOuGs7qvXBP
M69IQ6bjSLEqRz4VCzUwjORVukeGgdFYi9nh0DOLyP1fnaUFZTmbtSXp3LVZ3R4n
hZUu0xweh09/xn6QjZXbkM/pInV6vslkLWqeau1yyhBC+AVhoiB6YfFlDkXxeie1
wH6hol51klY4ruyFNyKQHgwodOtzLBeilr1mLHdz8V803W6ACUDHQ0TB3HkkLdmj
IZYNSRkqX+USEZCdEu6a+CZJHrEpyxOCybFOOepDxWqGXUMvlpqjCq93x9D3jpLd
fVsmKAxD9GPDVh/gliYfg5kmkMh+oROZj5RDvToC9nZfNRSAPHR6sOTlG0ij9ToB
AUic9ozG1fbD4r861SJzEMCbGkbWEWDrkLsZmhK9tzwQFj2+VcDiyqldmq5Tb87V
fFVH6KSUZ7zELNto+JbyWxhwdjuohSBLlaMPlerMmlUw8N0XZ6AR+1QCH8yl80sK
dhZqzOGid4XI4KkzUL95hXgR3EPvs50i0iyTBh1VisrjZgyM1jJ0Z5ArKsfqFI6U
qNZagzlXZUUutWGkQwnXSb0ERoz4UcVZB6HYWVZYDxQQgUmyvemguagzrfupBwXl
euuLR4br/NwUMPIomfs87oo10RXzF/u7zt2SV5Wz9VUG5vbDUZiDNtbFD51NVvC8
Mu6cffNPeN1UEpl5HdEH0Q0sl6DTtaGawUtD8Si6B8Uw3H+7w+5DApWyRiyyCWqQ
IR8FNKKNyWFpMmtrjwRRFqJOuej3fV2ENedPwRwr8tqAFvChG3HcjFmpDdl97Lgh
ta596vM4mSxQefeesuZW68R8ohTotPsfeQMVr0vqAXbLdHu7tNKmKGvzgGRiLlnJ
F1R7cEDRmJJXY3ouO7hylX2ouxKxUT8tZvPXhDXoW53I9Znb2N6A4kabSKA5pztc
N2+7jD2UvA0BJrglg3l29dNH53hezTa+t3Ph8/C7SnEBpxzK5V8CglPpbONMmyvo
BEmpCow89YsIQ68PL6osdQwPfru8PJXoHlFTDY992VsJ1vv1z8BLbEyh70PRrqG5
qISNv+ICLKaYRtA0M+RYVuIztksR5dc+q8q8HSOYaJDYb2cAbmbIplcdTagYmaUo
4kr3o8aEzEZNTg4YdqesBw27RTHjje46AbfN7DrXZv8LhLhSknUl1gdu6eyTA+Qc
v7fi4/ZiuWrbZWXvaa0FRGlfLkLwmpbhIfgSFZfIWTmaFLWjaMJGjFmi+kTJzoaW
tGrufNbAps6tRcKa/H+bFzb1NDFaOkM8vVUZeoodp2UJfplEwubPsu9F61wQ3jDZ
VQoVDC1t+PvT6hJRmhd8zdTFAPBnB9o82Kdk+jwEvG5uVEXFMZDNHmxD9CmOb4oS
gnpTlV0+Jt4fU/u4ecxkT9DJKpNq6P3yYjuh6D7GFH8gI16kNUcUqVEqOr6G7CBV
IJkos2X7lYwNG+QQLo0r6ZeBDpCOSnMBmQv9pxdH98XQOAVsqdZpTyo0pgWdweL1
q3lO7mWQjD9vL2xvHOxO9QbSQv3Nl1lyU9/gFeIIQjkVM53y2XKu2na8VFMPM5tz
y/2Eu0+6c6x/EsDbLd7HKhCbYOddaO0p5mXHU+Dc+ykGzzoqL4kXznv5sY4ag5Cb
glwMVe9MR6xwlRMeKUR5vm4445B8Q7FJ/dhvEv6nooO8P/w5+YmfvUO/sOMi+k5Y
DUE3xhdaw7RAEby6P29u7+L1S3HlLAluN1fgj98RNZSwr6xnJTulM1VLw3C++d6T
CcA24DcydUpkFMA1vWBpVxDkoKh0gN2RVDSKsd4OqOIDj2jXNRL4mDp3kRAozGj4
3eU7X3K0nvEF1HpwYWxdO0wMxcs+0kdXSNxJ133TDbBIDS41wlaFQZzXXp4iUXk5
GIh/StvgSCO/PrAE9+tagpet9SMUysIbDWBRhNoeC6RBLL4ISL9nPzsrI0fZdjEu
vBEZNVmpordI9MDv8G7U8crNXfxLEiZPrG1leLFLJVX/ts/Vddmrf0hqF8BjIRq5
ZRLm5x4IedEZVOLdyP45vhKF/+zNzF19YNb8ZVrvBxzFwGoUYD8G+vV+ar4UWEBf
IOx+xdHqNlkP92qZJ4IGj9XWsqHr8uIA5o9BseKXQSpFiwlopnquj5o9yvTjbndf
UMCmiW5kkJbM1xIcanSBpdh/41Z+ddfNNFggIIwPIBa+Fmv/y0r4jhkkJ42Mmqy9
OaQwGtzPVddwexwwr6GMhlF6AXjDvpfcHkcwd7/DJh/DkT/c7XGaRUDuvE1gHwn/
NxNR40HBUS9AoLkvjUwsWkZjB5rAmlzBCfuk/Yw8aVpbMy/6wVfxPP85R5xOp1u5
HOAwprfKi4m6byG3ja+w5wwNjvvjOtIblKYUaIqWhpd10oiaHfAUuSklB2NuqM3e
tXbB9+0XiaNnkQFpfYORAzXPav5zVxpV6tBxnoas9UYTZRPdt3jtcPO2Eoo5cwSl
0cyGPIq/A/NJP3hPbuPMfkJl1Y3wH51pQ3A+FOjMKthkGuq1JVNuSZxbeeeJDL1G
ZVRoclRkSBR6bd5J+GbxHhszYI7hbPUUn/J0Pq7r5FZSnav0nFRLc0LucdFuwP+z
CDG9RGbcrVmSe+UsY+34Mt3Rl5/F8JXFVPXY/4RzTqVgA6YZbFfovzJ9RTpCeAvF
Bnm5/haKVrq7w9xZDVBUT8AgeNYLvJZ4KMiiqFDGE4JdydFehLcZAEe0C1SW+GcA
m22k/HgxjmPmyHW0utyokzNkVBmnlWasE48RrigYme2XeGKHBq4hP9ZLDclBNtFn
HfhuSMmfgDN3LNud36liJHR947Do17cV4gQlT99dC1lZERMyUMd606o4NCeAMtxm
hopjM/Hn3dKjWmbVuP09gTK56XbPnspHJnt4cxcGPlndUiJ23Db4tTeMe8fqRymC
gHbWwlh/mNB/2M8cXb6v7RqED30B+CnHaUdCWUy16r6xwLNYlpwHHiIH73eVMSli
mwMgXQTVReJusRRA4im31R+XyZrvOXzAcsga5B1pR4C/pVxo+6WQe6ZhLnFzXPJ9
D4skZT6OxYAL82bfzkmwK8xrZxhfsbUaRGDlwRjGhyhd8Wex9kEGZtUdRmqCpe7k
Fvp1XDSUbbiOBAHN4b58kdNMjW8BjIo1p/uRl/+EKyAlCJOBOg4G/3Vc2llO1yhe
Z/MXcnoliiX+p4yj+7u3IAM29YpWR/iF42rfhAd40g//LH2ZJ4mn+wXpewkd7Xnd
3OZ1a9EAyCLaXmPi+IcMEKJhl9+yc5SsFA9+XG6B5Cfp5kAlcXiyEh810YEJ9z6j
GRKKyqLZV14jxTPYBVewNFHjRwErD/2lsgAcCqlqXezMZlbyNe/Pj5XZM8SCBQIs
xp07XOTosQ+bAVNJkHbsViVzb6PDncGUoHy78e70OLcvLSEfeQkLccwOAJ0dzKd7
xyrqYVWfFMta00d8GMX/glKfth625bcB9tgqOfAYQK7fjSd34uMfKs9mGmP2+w3/
4VYRf6C8TA2I9KcYq05CEM3qHApeIqxiEZ6g/fXRDeH6h04zDYKz0Hafr9p6R/5a
enydgitDBSrsGmSCmMshIf5H9XSAuuLBRKyFxQXw57QkGIeXsESAvCsJGdcwlkKV
ck+SwGFBMPpMS5UDFiRf0bNb5O8FeColCdTfRA3xMi5mZ9sIQKqgFv4OsKDMRhcl
6b4ghD47+4ozfkIunfIvg7cuCeiAeSkmN7FKAEimemJqog420DcdY2zL+E0xyJM1
J0OvzSQkapekwyx+uSPk5aPFU3ukWLU7HTujLpiEE3QAAGwo7V2U5ax1ZwhZbhES
SxdZnZrWON3DzWMy3AF6HV/q1bPwq11JLAZpnpLTvAzorMHtYV/6YVf45kcfK07z
XcX2GB1T4WJdCPndLlqCw1uhhiKL8WPMiuzwQi8x2/IdqLDwIrpkNtRxHzqffM1r
dYIitvndecuEcIu/KP2dqFThlFqTFDE4Tvs1YZP5dy0uqifcqiJSs2UbVVLa+qHU
sk1bZH9J6nkHKRSkVutGJc3bEhOuRm5xBFNlXlXjQuMWab2y+aa97QeKUvvKUWcb
V2S6SV53snJ7HnEfeEIqarea576CDirz63bAp7hrwdIlJIFVr/uIBNwc5nBVc6Km
cUC3IK6pw7d2xE2vBvl/jg38gLQcpDDqymEAMX/pm+jIC0qkaYmaQj0QJpUox4F5
WxUkIFmqU5D2KjH3dvnKMTP9JIDo5vcoAaA/tVlMgtgfoCwHsapM/jxrlq3GWD96
q1SdFuK5t3OJavNhmOiV833ubhzWIFiuKf3muK06gzA2qIUitjgBtr8uCdXK7YWd
VKjKLBwbJ3FDgHiu6ONOhc/jo1hVVCOvqC9IS0n4mcxZEs3KrOZRunpPx9FRFUai
gh76qIxMFRYf1W6JcB3dCLRmUGbGMuugjAtoxfx2hymgt8rR8lYwkmK5Nx6yH90Z
DYgD/bBh8DoQyygc6059R2YKNSzyY6gNJFdriH1dIYvJc2tUMhmJPsgiLldiPPWE
4Am+sCDmkfZqRWvmWJbYvSlRrrzVKVK89DREw5dHfFfwiKBCCtPP3u0zxbSzqW5P
7rmyD/X0uh4alAMegXXpdBbbwgDcjCzlHKlswIBzCqjA6iEVVQ7vIeLlDD4PbECm
UzuSFvqLZwpfrdUdFkYyncZQ6muAo5MMH0WJIUX/Vz5YEys7C7/bdoOqC7rEL2DJ
9bb7Pi77GKdkAfJOir/DhkRtLHft3w9wXkwxrxOeNc2rl8MLagAvDm9FGKNWSybQ
hk6p1T6/MK1dsYf9rO5I3TvoVeSU2nsqx1gATxfQCczmyev4vwTnuOqeGV0lZXdO
BHEcusTzHETFmSi3LaISr3DawxvbLWy/L7JmIRlYnSytHWeCokjm47ttBHCT3ka3
4U7ZJmR1qgM89D3tWFVIgmqEzzBKZJExMN72nhZ+WHvqqyxm4GpDwdxsGWMfKoqH
rEi1tIc3uUQSj28QW32ctp2gAiO0pBEizuB8/J7ZzY7jXEodPk1/hf5R4P3s3rpA
4LFe2nXtm4hGOuY2v0PoCIEu2IHOT1Jw1k4p/mlrdE6rSwaX9OuOgUmYvvH966zD
FxosbUo9JZ5i0Hz57xr4Q9fMJIKXnSsJ8qJmXgH/b6buBWQDX3N5v0pZse0qeYjk
oG04nfHIIIOkiGSZxD9cyQVZRs8GQixFMrIDZB641ObLkwtCk3Bs36mVIIckFxb+
875sOXCdmbIxbqdYCFph993cP1/7+HmqwXX28YNMONJHzVumNPoZhs1QjeDCRh5t
8Y5prG3WBD4JAOwExbrrfhjNe3F2AAa/TVrxgN1/+5LFtUU9SWq/PziSCjHWoz9m
0Q9iT3mAGfVTG7ZCxCK+KCYZG4Y/7lX9TemzccWMXgRUmQflj45IpetqMABWqbLx
oSMoHYeMhPerUUm7A2tdTWQrXA9edDBWgMr6/McSQPtWlFNxWuxAruyuqMXAl6fN
2U2MYG/PodjxgLH55FqzrsK0UAkvyy9tUNzp0F1KSkzfCLo/dajOpZLKEDoUIjob
P7f3T0+64Krn76GIYcAjVlWiNNslMAuJGC9Y2Vas3WVu4h/DWZoTN0Cj57bez94Z
pncTgD0oPWh4Px0Bh0ILfgi3PWZQvE4gj+EwOkiLh2KZcKYTJJ+mfQFKnkmx1+Ah
PjyyKe6ndFB9dQNDp6awleBHah581802NZ6dpG0BPgxJGwME6/jCk8HzBBnOmIOW
iJrreyowuVz+oZXY4Gj1+WcAeCTV85SetdRfupU98ArGPLQKF/+/7T7Sg4YmDPpv
iO6+EM7uY1V0kNw7CgkEqwta/zheeSw9Yf4RXJBrbVmLzMAcNL3BWRjuEUT+bTWA
PRvp39Tt94TqjDNPFrP1KegUh+Ck4eBcFImFdiV0DRtp3YeySoKt+XENFphz4H9Y
/kln4LJFjaFsp+eg2NgJG5szrf8hKuUS/EKnrVYAJUnwkI1faX3ELSk5nvfzVS91
HzvcvW8C7i21KG9JyoMhoJe9C/MTZwW+kLONUUxgL4m2Mv3yGG1oaLG9lyypIW4L
71Tz1fi5AlcwDhUpmtpXSbhz5PbD9epe9laSX2xHpAWwkU/1pvoMpcbscIP+oLln
E5gQ5kLOmbLj93Ot9a4QPguuvaPabYSuohrrl7qgKQTDqodaXJ1dagcFgqKWKUYY
WMmJziVSJK4tcti13qYbuV3D7ASGlWRcmH0C5UJRq1jTb8EXnl4IJW26To8MaKEC
45vU1hl5ouqwM7Vd7KqotPu8CpjGAGZFn6CI86WD8E2TR29Cprcd5RvzhRZdRRER
0iL7GbcMj6NuMBvUt/hNYiXR59OIEXGkVFRySYN3/K492xvdOS6H3zDoxd9gBxMp
3g0N/d5g1+1m0lL8vNTNb1t7gDmNoew0hXjei0om1PEB04I11ZEy8d39gcu0hPXB
OqEeJRpDkQUAiPo8WH0fQpm1xK+6UuzYNU9fHN5tJCcVyA9AoavlNTMIfbXCjw+f
Oh8QX6F2Q3ZEXWVbRvjTls8/PaIAXnuWFupZPf7M+MjGner3B/w2mY87hlR9dZeh
FdQCF/b8WTOq0BzLNi+D0GE8RQhPCvKdEDG8Vs/ao0fx7EWWXOkC5iSc2+Mit7Nn
c26lIP7g9aIlVFvqP6CWzBloo1QkrPiQdoHROBtkAjhujhlhmRHKbCp5q22RMhwJ
N2UTYxOUNPXbsCpeVaxJopyaERWJS3RNBQ7cPEYNgoCx1pnPTihner5rSbNB8fIr
qno0l0Sw+5EWg/9nvYoaJOnvwk9nMbf7An8AL+RT0Jbcxjek+qGVqsByrVM1vbpD
1QZQcbPmESy7cmKrM1S1k0+ZOoX2b2ywseQr3pWOuEcxnx1J7m1oDDtQFW6v5//q
A4AjTQfD7Q2OWVFoA1N8QODnYfu+fZSHdI7a9+Sa3NT9b77GomDW5FrN7vGGQlrf
FcYyWB13Uli1dMm7yc72ezpu8AFKnsmLNiheM/fy2VrOaXTcOwWKUxzEpWonhobp
kSxEK8644uJ4lbkp8dTuVM5TRLt46izfJIu7Mag0O68Y50BuO1Qa2gZ0FniyxZGn
hAyV4HLFQX3oioFkAZ7P+YIsfiWs6yi/sOh/g0Q59wsvJBi2ijF0Pypw5etKl6al
mx3HHFjoqPATltCCsu9zjFpAZ6lkX2HdvV0O/HncIEhxso82uOlH54Bg4tBFkXzd
bY/tHdfgmbFQT+un+QCEFzLalv/qXtZCI2tebjAHL0SGASV76rQVYKHByPlw5xoS
Hrq7ZCVeh8juoQp32AeOGLYUjfyil6nNjHJm7bXu1wIT7UqOzGZ3mE86MyVd2V3x
29ff+wQsZVAHkpuzQ+ap+2ds2YVc9ElXQyDB1GcaqsFXDY4tQHJGs85iF12SEb5o
U6yN/4PY6by7xpdA4n722WguPD3YB6cInoUyfi6QijpwoZbDdI/NZBWNegBNfUDW
75hu2zNFo9sQK2gTDBiCorgKV6bCxqE9xGg+e4/CJNeNGyxoUeT5WfvNjsvt4LUa
uuNo7tMnx+BWUrdBfF9K+0fiVutzPJOp9sDJtfqc1M/Man1nTAs8BxBP35722wEk
0hFh34nxszzOT46rDMzcbHwHm8slr1VHDiXOoR2ONykLDvDUjaq53hW+6WDGffQ2
hDBVlwRCV8hgOZFks0Lu0T9xwSH1Z/Qa5mSiBlk+Gr/6ipI8moMw5xA70sFgcbqY
Y3TQnhUdRMVPu6YtW0NS1hBNwzjdZFeczZfNbbEYAlN9xxCO0ct3u1CLwni+sJkH
jx7VG8qjvq/LTErbLYf0nT9ANuShb+Ro1fd6PMbDn8xEqhSgN7lxV1MLhVjbleK3
74FdD2U2D50mFyYnhfrnT3TA4dL8sc3Ccf6H1juZh42f91ecvJmHAL375Spps6yt
HoXVPnVo8rtgYjCKNHo4VE0nUl8DfZ8ELeTCb2CctWVv7VwJY696WLbA/IusQP3V
daVdUL6bJePhpdD1urxFFNpU2usDLFBi6BPh12ibEapDvQnj+ztu6Sr+FzWdzzE/
sLOzdVGTpcapW5omF+jmGUfQ8IRuFZgFPO4cL44YrKthDPakzpf8Zf60wy1sGq1/
9egT4e1YfCqfJAbt4TbOYhu+O+Xo2B/u7x9npCeaCiWqn2HZQh+mEej+/vJT3qll
UqxAGTmJFt0Q96aRV6iXhfC5CFN14/7k3sS+wTczm6O1eA93cLYRbAcmNklw6pF/
q2F3rQjLOqJuccCrkFZgcRNvi0tSO/eyM/FhpDl0R6XG2CX43l/MD87X98EhqFq2
JEJulJq6LLhBXKOzmrcF/CRl+S4pkIDa1zAquvVgbaFUvE8P5zpURa3nqVC1Nddw
vkj1rU3xdm1OWGsRfX8pW/0JKJQL9Lku1NyYiveoIWczO39xLmXF+Iv5Xuq6ElB2
NsSOVIl0AkVvy3Lq6/KrZd4xCaGRZGd0121gW+HnqoVuclk8b1FgoOR34PhZN6/s
EeMldQxNLHyl2qnaulUrztyBtHuo5SEQYFCkqib2I9Nudp9lw5ubeBctHlsJi+X6
MO31F5nqjOh2/CtTN+XIegzmzul6p85RZWcJOOOy24fQgQFgD7XNDvuZeoJBWMPM
sLBo2yuUafLILdhIYSckGuIIXRaPfnsA3h8iY1elpkhEl08k4x4vPjMbM1vSZ1B+
wf174enBL4s1kjNH3ZmoQ7GLp3pVZoVl468HRsnKdQm6DLcYMxQZQrm//aJtQPwt
mtrgL6145t6doGuiZd5bAAcQnnUQls0suDnA0qeciIR+VVn+CfoJt4SJOi1OdiI5
g1AdA2cYoqCMjMCarMPjUUD1wiUcEaT+r58kKsTJUtXO6U6ss2FeeoiKsticOI+D
ighKFc5epB5N2W8ZoGdmBIgV+h2zRZP+iTRQT3qWZKB3XzDIEYgtkgdnsZQSlWn1
HdcqADH1A2iPzTAyDpoRKKUzfgXEgjAaWiipWmBMq/2C8cAW9ORsKH2Le6abctu4
tgFkJN3xVOKjkEEJDnxfwWmOrxcBFnty/zaEJOzeuognB90i6ttCxGhDKGELNDUa
jr6qvnH3YkLEhAPMuLZTqZvFpXFewWqy9jnm4mXwpALwduvRmmkoymFU+68XU4b4
b0wpn+IVC5N+O87TWuQrJyskxA/ISK1QcVDV/VrV7TqYU3bmw3TjB2HTfd1QZCke
sK9P57MDImWBnZSf3CLPzOR168EokE4NArx/a5qd+Dqnpda/oIWeBAfugtbEVVHn
PCrr99/CkmGyS4xVwslbkszyO2D89ZrG9gBKPYA2crjlGI/6Rtz2GTwEOZ6oQiyK
kFYdwFq3yc1GBH2Y8sZFp5vfrjeo7y+P9T0qaWJhqHsVOllyuChUDzX6SFZ2pEb5
CNNtomXadkfVcOtQXbdY2tzVlQULdJ/9DFqr7yTR7UEIaPqQpl977oAjBsfWO1KP
uXTrt+6drr1yW3LoGnMwmCoBtqkPOPCskJ4+3mIG+I9CiqNOVi2eE30U4mXN/0Cp
O/nIWNvdtqG9qQrc322y7WMAJ3pFm/9wsFNa/05eJAE4s2I+ucO+LbTh/uTvHpkY
r2SYciifcxUaFWo2l+zCigcTeYirSOEFkhb2GoHXxCbt20We5f5KovATh7bzFpTJ
sUD1Frr38SR9ryls7py1K4Dh/s9IlLCi0OqeWDrDP12PQb1JlqF5Omjgt1jD/yEj
iou+pgdWLeK7qTMpAPjSPrg9xUozYtU28RM7Kw+tWPpzroCTG9R2dXgxtGuQyF0w
7zBw//AVH5TnN7jPe1KFmZPiYqlUBgLT60roTbdYrHCqk2jVGsQZ6a9X/gmWysSl
2lzS5V7Ia4YVRYaOJe9qbf8kFIh+DA4gsGiroDq/YJautJKtCkmsGbJSZnUSt1kJ
dchgriqcpBz2tFSJTONfErN0CPSzF/MqoUa12r2x4++GjqMPg5v61QIT/Q8TU8wK
1XOzOEc58IfLxKyzWd7mMnrzhRNsUZAJTCfgA/Z8JFjWH0/ylachcdGVfwLQJ1lz
rkc9xgXSj6fpZvoTXl5jlY6tPYWO5FqHjqzVAdhuUN0bnPMAQw592kIajcqEPiL/
8ElMYtXRoEq9Mf7c/U/GGP5elbpVD1dbhwiXCoo4JkY+n/zaTxNf/VoM+IxYEFOZ
npAltphTdszpt0i85ZL6hJIOl7IokLYWImGKNE6I38hprV8fMeZNtbjJZ3AW1TLy
748IF/YdqE5V+Pm/QAwJ9TjGZik2kBsbhqTTdODcm4R82faPuRrr9UwnSNBmmqYA
JCPq1SqzL0Fnb4ng/iqsBPnnHESP8njfhEANVJYYxuwzvVoMFFQDuoD/RJVz21s4
XH3BeOkZZJWB/cyKynwMKFU/A8VXBxN9ELH9wwuvyGUKK5WQmbmP9sFjkpAdmGOR
EBhoT9ByiJaSBOUo3gPheUdcV+jeGCJVGCqWnatZI/+inEaDRGtANFNPAJeNC8pN
Wf/IAoncaz+nEZEFTGwOz87dbWeqtulvDIX99vAyVu/LW2I1pjVv/O5unGpX3Z6q
CWi8ba4AV1RAKEZ57Yy86r1FYxLJIrZcML2yqpHdtO8xcKkjlkEGkqAlyveMAJ3d
loJOEyTGb8V1cdnKgP2cPSOtm2lrmSjan3Ds8pDEXtd2xm0CG6C6fCk/k/Mni3Ob
WwKfSaO6PRcU8Y5l9MHfbxwpGNkQjZ8B38ui8Y7gNoJ3NdgCNCpHknABX4G2c5G9
l1IOrztMH8fhWsANmIyl0NoyYvFXDaPdK4gBV57hgzPRE3dUxvnbu1pERX732XzY
z1Kia9OO6AU+hrDDIvfz0FphrXZInVESt/WDySxhAVcPOvzjxh6SVTzQ+pCSkjDI
cR10AmmhBNtuCDPl7YWg6mmf1t7qDGMnwUe/t2UiSPQrlZLmSE9bcDFCkp8gdNU6
MYqRBo5A0i+EieCAbZtM3eM2YUkMOvwbIC+dAFmmfVaIIfMySC6k2fozkceljVxt
2ZcwCSxIrOKH8iu+Ik0Zkm38MEfCqxM2iKIvSRtlchiBH8IlRl2bHEeKoJDv5Ee8
fwNCE8exHzW2UP6OSwzo6pa0uorDOXl8NO/uGmzImvQYjvfo9LbDSmjJlIFpOdE7
XdMSR5dz3AMDz4B9qZJ9tTzWlnDZHtKTrfaiQAsYjFyBsUe0TP+sw6++LOwZ+kgp
aU6PLGgfokPaRMnmwzC4JgPrNQnHdiQwQkxAapiLPjcvjuCJDsjDhBV3JcAuWAf8
f7nealZ6fhAxe7p4Dffm32gqNpCld6IVtT3O15Df7OUt/Z4C+VNy5hJsY3xcEeu7
BTQWZcoelQsJ3iM9IAL5tPdBtrpuT1NhIClrtI9zEWXoupLZCawrpBR42DeBA+cu
D4TFnLhagkxqEHgutRAkkykckjORiLkiesG9Txu+aegJNBLXdgyDcLxjBZWKtJYZ
czaTkD6Vu//qR19yAc6V6TdzxxXuWLJ/5hUEvMRHbZ3BNdLa3MSx6P4Hw1NsUnau
I3UkFDB7nzD0nCxEZpyq5anGLGH7DNyC6s3tnTcbj7pvPdACb2J6LtkZe2jk53in
O4N0duAbxnXVWf603n3EJvaqd3UlVqDKk6/6hVCOExtxyJ+7QhgXtx9Z7qrJRxrN
UDNrhHuMERJzLytnJsJFtyuGZzYeIy4IExaYs3zi40S0TaONyO2V5vpw6KEDIxMo
7mkrCPWb1RXiqBW9C9DmaYAL2dOooo8WUoqJc6xYb7hiZ8in0QLpAN2dQb1ij29O
VrM6V4viFyhD76EjOzz1qAGLt4A0cV+ccb9JsKCWuqBPb8sC3Ctb0SyElal+T4Tp
84qVauz8h0ZtDFaP4wTR/FoJu/N+PSIYxivbAaRlLOnEkLRNOuRCs++KPLoSn/tq
RHg2F1tDLXwArqtkvcmeOopz5C6myRYsG9G0h3a5j5O9z5V2d0py8EVJOtlgvgx0
c/7FDEzbu08hx6smNpmI4nDdUomgHBbvZBW0iXh8lUwRuta2C0lmIkOADHwLIknw
4xinOOzXd0llZ8BxDbmTpH74RxBee+bu9EaKeDQM8N33SxU3lvPlNfst9ZQgA8x7
PD0YMbWccsHQ8tsv7cpaTNdgJ0RdV4hHi8F6vOdtEzai9lYjcpYpRiPJGgGSLqbm
euzZJMkzCbEXnQy/c8XISHv+awNRd9TfnBj/MAeBJNgxOUXvc3OxVpSfqmxGAjP2
X7b6woG4Rd7QlhLSSBZQOEDfs/f8rAXSm5n9CZX8eaOh9I3A68INijasv5XsyBs7
o9B//llFZIfqzhbEKspR3ZOElPbZ8jfAd0It5GxSMPVTFz6BMEX9A8GXUvm5PYsz
L0zj6ZpuYjb078WaP1PkTMlcspS97ytvvdWvBFVaYCFvp7/L142TesSzYBgPbX4P
5br8E4Jue1CMJjlbWXpCXSCn7c8mP54QsSqu3G0k4iXY2ciB359zpPllaqOvPpnu
EylI7r4Q37ojTfVR/DPW2TgmgPJbBmxehIuQJBQ0XvhiMC/QuGLNuls9lP8tFYNF
znd4I3vJXN80CsX3sqMTHpOGZRnhz2oGXQnzorlipUSRtQY3pITxP8HtUj8avGzD
uCuzxOCrd5sO8W+GhruJzAqLo7SHdkB7K63t6iA4Q+EisgutKmplkjYKDMASlb6W
kqGQglQQsJL9isyYgaInt5D3772B1PYcvBCN7PgddIezu66Dmg7f2fkwaV6DDRTI
8S7SnmViSnc4SM/kfu+BA0S5cq/g7rsYmHd+7FZhB93xfx6wBKnfETk0QpevO3IC
SFPYpy4WBOM2qI2NXb+lB/iVIdQrHF77hSwWDwLPg9BFHo4te9qfxWOfE1h7Tusp
M3HTOwslukIpTR+zO/MMyXZxCmL7NcwkVvt+MEQKtem0UeB93AfRiTK6tBdyB0KX
kNysvGdY3KbEMFzJw5eQjgvXLL1jrVW133JrSztDiGc4H1MD2UvUVWWGoKqMekgO
IfhVHbfrPr1ZI/rZdNu2s0j01PFcuPEQi7/wXP/JwLHhUpgmGA9p19PodX3O/6RZ
jPCnAG4aDmNJ+AFVrjjXXTDzywzO1CSzCwE9O34ZFiVa0BraSmceZC/o6upQcG9D
7qxNgIOPc4gGZzPEillJc51nlvmXalKe89E2fQeMyLxpFKYl/o0QW90bPurAKTe0
XoAHHMiwTxiWa+EE4rdH/CLLy+Y/WM92YEjurljIFdHt4yg2aNZruGiZiLBeUWMh
Rl24ehaXvv4Qyug7K0ggrgDcpfQS9lKa0dXgnh7Dqq+44jQZMxmr4W9M9vNk1oos
TNgUEbpi/sGkyGfLBo32mwSXGvpLYwdcp1Izb2hVcXnUO0Wp8w9DdxU0BVAcbKfA
MY9iviRhXID4xjvRFVDyRP6ppQDURv6AgsYnHg2VdxLf1XpBba7QSN6V1Lb1jb2S
Jag+SnSJQ9c12RMivAPn9Iw8fXESgZKjMZS4YlKarwmfwrGxeLHe++FMJ7eTqf1r
Uh+WSp2UxXASgScE8xzlsSGDrTHhUxr3tblcCNp824CwzLDKG0RBshD3JpGvMsjZ
r31uV9w8UDabs9ZN8R64ElCSn106c/8+I4u1YtrHiJovn/TFInFqTU9xXt8dNnLu
ReoGm8Oy7+Z0s8zNxiZ+YEcs5jXjXjW3mP3jd48AA22yh0VLMk32fE6ATOPlRNbx
GLFUhgQNB4HLqpVGxqsKxSojUzNDlYOCroY8hspMSpL8jECTWLWPtS8CBX6ezfNy
6xud/ulD8efDCvf2ASGQjQE9hX1zKHLsCb2rL7WXKYkXobubhtBqPZUCPKAFrhMa
u9PEpwEQzT4hjp4EIDvbELzT6cz10YtEopkgWJGZMXTegoQn0rpcZBhowXHT3pe/
6OwtfVnSQVtFHMj9CsMkwbVywwFxQnM7UCFcjvi1+eiuNDtsqrolGCOM0cW7dUxe
8j+96cqZY4qzE5GUHpxxO1B92Dtl3IvfFj9bPK8l1RNCZdSPlErsRRcZ8nmnLc9B
NMqNHQOIyQLTDi0bs/iJF33e7fC8UV8K9/G78/7jDwOR7frET0Q9HBAfVPuq3YJK
IQ8NC9pGI6SavqgR/VsomEgaHjJsg63qV42Z5W31eiL7m/LYrhvEWnEK5JaKxgql
JMPrXvEZ/3aFIN+P7O2iqaCcTH069PjH5a74dG+GGrNMd0qkxAm2vDgr8SBbpWln
CIILu9MYkC9+teTaxp/8i/X3PhXrqGzSIf0BSwzIN+115i63JgfgfG8ElhbQJegl
zkuR7mtu/n52oSbdyKpNn66qE08rDwS73jnfRFAxc1MXSB7YWETK0BOc9mIvqHae
VGY6sWgfmQfe04Sq3NNPqxNoBREqr94yoKmi12nycOsddFtmDv9L15mUXTtRbyPk
6pKPE7DUFg8gGuOfpwIGhVchN3EzRzTwgKkuKL7AyY4wT3IumRwpHMMpn6/B114H
K+wniy0l8s+G33Y+8pm5i1KYFoKZcn+yU75+lSOGE53UGPB+osXhD7a7RBws3aIv
/4+gfwZHFnLfmiw32omxmvqaTUiU7DRd2hN1wsRAt6E7U/EA57fsefQ9K0eLvaJy
ON+BVO1o74iV2vdOkkFBCPWVC93b8+h+xrWRDCfUPTgQsCDGaVyv9xP+Ijiq1Efa
NGcPbd3IUgDu7lbPOp8IYPfS2quhqMOO8pGvDjdB0RaUyr5eMfXzRl5usHym+TsU
/9ebErJXrcsoBhU37QTgxjG+FNP+CEw5yQKQovMOIwjGf5y9oDo8jskGioHkmb5C
q/fgLgg82hqRnfpv6kOilpGRT1GxRsBh9FwsbRWHZSsuEBpr8awraAZb5fUZU9Db
KWHL//yLYAl42GD3pjceemaf/PCEpq5ur3CPGwOOje7lnZBaerOyhUlXxJPh1YS/
X4DSujg8jNJ+4SA1MchlLxVYO6xxYqEZ4JaEkfCQ0WprUGNtUWqjO2vrcNxmfOdb
pWA6RfCm0cnqIWRYNyOfeDUsFgQJJhrHdsMFIrpN9/w1lpYAHDSKTBsJzLFba/tt
1Bly42F0nqA480h59wxFMsl/2RU1D5el+nXovthj6wx0i6Z2pKrS1Vowx9NaXlQA
OSNZ1zgosNfQX4zd63g8lkOT2LJqe6a/2ihFy+d1xhbyPFdREeKSHuL2/1aOchda
ty9Xr3kJlFI9StPYljEryeTWYSI80CffAS60aMOEyYafILd5GUJlTH1laV+iWMK6
qUB4+aIN4QtgTxIgaxdA9Tn10C+PCTvioHzj4EnaYD2k2dNa5igcqYRPCfzyg/ng
UPWdkc1QTKeHqgnce1Q11Ypd7+2s2EIsaAYASCR58jDf449v1dMDj83Xfo7AMC3Y
gcvuN+Iw5l1YZMC7+Tu8HuNgkPAMyecfl7wKvMUHvE9BvrLjODhfams8UnItqTEn
jwKWWVNNDol68caIrd0wD44FqFQ8LG8cnvw8b+5XGEUaL6jUeud8Xcu0efIjP/ro
aUCXUvUwS7OssA/IiButfPzglpQGoXhc7Ul0my/IVOpio/htzGEcPzUy0HE5mtOf
tvyYI2grEimlNyyZim45JfiIGhqepe6uJ72QtVXwAatNOgyKFxcjTmEmJgUiAYzh
9akA3FdNzcC1JWUbuyapp76JghENuUl/i56qSVl0IDcugGb12AWa2qgW3CLdBlCm
Wf2kdpu8aMvD6XWmJ7ZaQJ6TAhwkcrj3mrUKDlcR6GjtrK1yvv46d7hSJckzuUU2
ysxFLnsxAoqXHOMihngm/MUDt/z5RIA5DoU+kPck+orDWvRt4FOZ+adNCLe2ddcJ
dDY//+GGbEUR+bPGDhR5lVzsFsJMOxMBaJ8/hYtIEMGmg+gvfh1QO5bgG0VoKjPy
jRs6s186bzp3g5jiyAP0q6H9ZgDsvkM++WA9/csbQ9CAPZoCx9sBafjmm0d+NwO8
VapreD/r5vtFqxG3k5urc2WlJwyfygh+T2MKt/Hf91a4xVIuZMgIv0bsg4YI6N5b
339Afuw5ZHaLDfMo/R5FuoKtG67CJL8rGXvMstV1GNpVQRr5ejTJU+VJKSyCgz/O
HUCrwu2F4rQZb1HJD1H9CCsEsAy97yJ7bUezRfAcEHt+a2VBwkfCYO/nrx7iLTGs
rrFFkIFiCEpwU/BFjboUipmU+ONVXsG9I25+0/ydMB1PthVJfsilr6pbhGFSNW9j
J3EDgXPqhth96dagD4iiltIS1kH2mIGEJRJzD4psjfvA/7orpVk6/RBZpENL4pm/
uuTWAetgTgZz/BkYPJ8HZ2ub5HtB0k9rELguGAO1vaKDNap2OoN22iS8htDLj889
hQgQaAX+UcJi+pgNwl6EenvbruxB1ecQMs2HB/Ps8u86wr/Zlz9A5hW7ycMFrS+4
I77FJLUfeRlzbvMpN/M79TsK3xDNfcEmCEi2Sgvni1kBO5gu79H7oxrNaBt3Iw76
Ce79N+pOWsFU8GF6I0LxSL7C3TD+rgIPiFzGNah83tR4+JQWy9rQKrzmtjAu/fT4
kpq8PnG6lRWZesX8oyyvLtf4tAQdVpcv+pTDM7ufbK6OBzqR3HG79N7lpnu3z3yt
7evi4p3BiX6CF0wyQ09/3+d5HdvHT14Z/QAemGF1TBZDZ+aBzCQMMxI5D9isbeX3
83DvYULLWCxt4zzzDXYbUJjhP4hvOemYpTkfM/Y0BG+zIDjLKXCEJbhNH12M6zhD
+9dz4UBrezdsGrMfID3fV0T1U15QZF/Rq9XXvSlKD0Qm1BBYUAdKvs+eKQGghzdF
mt00fiN8+whsg3DWl9KN/GLQsI/hP1XuIHih5SA4ofb4djohbNOacnZOhpOTNKDp
X9Sef84MOri3atlYtuLrFb+EPe6Vf+ih5wt3Xct5C8i7PSAP8ZCwJSxeXeQUAMjj
zFfvyF/AzNoq7QIAqLu4vhMx4JMOJ1Slokw2ZSuYm4yebbgIMbE1ZGS4QpXgvpP+
I7+EIVQje0gIjhTSPRHqxuQVs0K1tXHjbr7OOsdFgubjpFEYrrWuZAPWbrvbO9YU
36XD9sH2R+AB9PwLo+13H2TFl2z/A/AzQfAhQ9O2oHmOAY8q9GYnWZ2vM9ArjB88
zQHOaQIlJghIB1pDvOld+cbhTAlXj6PbFYSWcZx3O6BkVdPb1+p40ArH8bXu+4ES
usBPGDuqlGTYCQNl8EW5g1d1J5Bme6n6ypZF02g3cUG/GDRZAt2NqsBpYhqJRcia
rCEBvYo0krp7csmNj4CjRTFyhU7nZsKeVt4AnAvO0bG00myHviUa9EDnIpKRw5Pa
b+q8D37MhU0R+BN2S25Itq3fNc910BP6egIjZFh3MJyO8u7P6V6qOtZvUSmhaLxy
jt2KA9QjwGZSHiDso9HFGmiGkBPS5+yn/yRSZfRAP5QpkibaiWacAk28ggDqFJMv
hd4fea6oE48ilFMVglZAUXf8KHeBigXTSb66n/DclD3jN5GXaEOe4UV9Q59MKuIm
1U0vl3iWTnEVoAHUWlRR4p828wx0Pq8207PrR+j5qpv6ZZ/JHrInxGNnUkSNnf3/
+Lyz8m/GmhjzxDCdsN9E+L4jOY0QprFLiWKPmbDitf+fb3SgML5e0R7SXMrO68xT
5VsLOLL1PyBJMNDjhJgKEjg2cfJdC73yd5oPzqzgOt6Cco4vJylaT9UMxZufSQHe
xZAVkGzgx+RlrKt8xYczbu57PmsfZCD97+6SYBy4i21weYr75xPdbzUiVpa8TguL
Cu2avlaP8RePPvDNd8cuInZZw2AUBonATpUuzKVkt1byFH1mpoDW/JyTnV4a1nDM
rk0lTum/cpkCT5pWQLFZd1CWHbvkqCRvqdQ/FLBgkyR0WxlP3TISdRkkXz4Catk/
Hq6hmqRkqKg73+zbVsRnxIh7aCMX3BRC9ZFSeAN7zTsWlW0rS0ictPhcnbXo7Dgr
uKNR2wrL4rn+0A+Sa1+dctcV8KtGO/+0c3PLnt2d9nQOsuQKHRjn+TENzuvN1/ER
vNFfuWf8F0KEQUhO/M6tv2FIcBKhcLdARpvKkCwLghT/tu9CItDmhDzNvmYG9Zkr
D5gcL/9W71TvfALCqZUZkCKiAaHTxiDVnkOCYXbvNudCrBiy0P6aqA2e3E5+u95V
i8u4I03pE9pSBEQ9+wumxHYnTvW211qkSMtquVScQtxU5WzbOq5BIoRV+MNX0tlS
92RpJUW8Or81CwXdGPl2HCvQxka71355ubCMsHbHYpI9uCcdcZzRUw5H0LlMXzaX
ocTYmuHPWYMO6wT8t11lsHZ8npDHvt/t6uX4vCqOAUoxncDWk3s2Tmm5wln4l8PW
4gd4vuwqK6F4gtvtAPaFpprPCaFiVu9GXAW+ydhNBj+Ps91IH7F3G59eDbQ8O8hS
9aqRFnb+DQzzTrDJGEmBCtX1qo4xmwN09tOxR1ADWCVhGsWDxDzgVhUmKNBX98su
gTNM64O1KRS/o2qUOsxnh2biU7MiE0fO0LiCFuNF8P1+Sb91f/77WCoHJ/bLMTu4
q2r0S5urKfgIdwnz+LTwlFy/YJFdvb6CwWTMfrqcymNjtfPHHnYgrutRqaJ9O7+8
lzhG0vWVv++x7WTljyTuyuXIzCIi4gPsZkzjRNH5pMOqMxslJtulK95lq49jO625
Yu6ctbCaDdpOIQf0sysB8Tiv7AW1dVrgWKrIWM14tzu26uVtrRpiTsc+kjHaiv5J
n8rpnau4Ah+CT4Ta3wxfRvp8PbrfCcGVHT7izUD+YSzKfjIMvIJ63SOp7YpidIe7
Gc19nPdZb4AWl/hOqUfEuCWVxVogdHSyDiSYtlMFKm4TtWHe3PjYMLX6ZOCMpWFN
TzzyB9TE6/mM6o/KbbzI5Pqez2ZFL/OLu0qFPA6DQax7zNlvXhIbB/HgOZNH9ZgQ
P1KP665NsY65GsxjaPh0pyuYJUjeAwuw10wEmMApHYUu2U46Y155swXXgNEn/dpF
Y/jD144vFzC1P4zlLXoV2nfI0RjdPWlOQaTQjaACA0GZk7sxurS3it2cZeR6nPEr
K/lxpNpnda4trsq50b+8/TJJxfu5sWNb9SRLJq4e/I7R8JyOaoM31YlUBr+cnqAk
anx2az9EzR7Z3SNL2VD5nWV9fxoBnvPTEno+XrrknEAUNJDjDrcrNKoRaJEynuaZ
slCQTmNTFeh2Lre9y7rHnNVqmoPxW45OsU2SnPL+kmD/yknLpi2BGJjaOHhwfy8U
pqwqToEkcRIfTGf1IgZszPPC7EDYblcSvLjPJ12oS7h9FnpnxycFx2cj52a56F2O
iaeoQqa5la23hovyfiLF7YLFGDyt+edfZ0zORtGL2WYl3EYYqeSR/AQ4FvnovWL5
HHNqKIZMQGXVZqQDNEu+MnqI5Nrqr1UBpQdsbjOA7VwLtshm9H/FsHUqgdgjBRKG
vy2K2uUnIdg2WFfwbid4yxPyxozpKX1Eayfpi6eO3IUEmUQ4Uj7++cnAdVy9UDha
6TPWISBpxLLMSqlbHUEZF3UHfdRFMkYZg1DBcz6b1ba/LtxtoO30EupUUCIWDzSA
qEpczwKw2NhMm2h3bYvA1XO/9COEtqJSMf/+jwCK7A6zzd93QG/F4tvgyMy+P9RD
CDW6F6Z8bLangsO21FEgjhyfiaQrvPhMm3WuT3NYcjnlTLK7CUvab0ObAGP4AUM3
qpxovuvypN+9Yndvyn6sJFr3ScUaZH72X7EI7P8kgEzeyFY2Id+CS0fe0PNd8DNx
1pBVRpXXq2+BHCpxCbyaRRSqEvWCMvVWYro0VzCm6x0Ik4fHJD9JH3+NCSOOmfoI
Q61ye1ISSA1Ev/d8ROd5IvONQgMEeSttdYLMsOpS7Ar0ihnCIaUCDuGgZxmf2kjH
454tlZSVhTPv5qSLh0BakWASLBTU7SqgDkuqyc/7vsubqUli7kdoqArfZzQK28Po
A6nIvXXwqxA3eqgARlEEOIVi1LRCRHoksGXDvlc0mrfs139IRMcqBNtzXO2YEtC9
K4sSQfVOsEzTFrCTWklNddai5TfWYJbjtNYhytjREaiCamgoDGGsKa4BEnZ5yfOy
2FP6cKByCVxCFkW2OTO1JAePcp0agvaDtNrkAAKUyZhYFvCJQn9gtJSUKYoLeWIQ
0LfG29PQ2jJA1HJ0TNlW0vJE04w/su4oIgsfOfbeE9R4I02d13nrRr9WClG25hgd
4TQuDu/IMljQwDXaR8A/hbdLMg61qvX+4chKwzcW/52STkvFOj7Rfxtc9Bk+TfNj
Oih9IKwe4rLtg0lMszuxsSO1ZkkIVeicinhaA7FERhL3g6mbcDz9q12jFDiTmd5y
k9aeaFLNkq9AEwJzzjPdLKAt+9rcmG6RFGICPUBjoj9OISAo7nYhpJ9rWsrFAHH+
GSLhq0JYIsNobf/U4RVMWnFr11fvA+qGDgBWqfHNjX26o7Mas36ERoVD/BAJOJiO
gRD+6lMRllXPuJyJk0ksfUJQXCoSHnXOJ1GAVOtUMlLGXXK6ndYuXLt2xeZ1kLjf
279geupEFdcCvjiM5Kss7i5+eAm/xmlqf51npAC7uRGcfW5eYacOfAV0XdXtCBPM
oMm3ZH83tevmlCOuBBKdnkrBDogfhwsKsskX91pq9JsZu3C79XxZa/1qKutx8jPg
ZKCEu8/4z2l+imn5ad44fI2jjxC/Fiov/V43SXyDEqX7DdwB6NWXOkYz6sAGKbLj
K2+3OWNiOfXpryPlOVw5rm2v6sArLa6sE08dBEZdT58Asa8IY5TpZj9txB4BShjU
CA1Iux6od9BNkczvtdbBD6olVgFsgnxGzbh8osM0Sj9x6GS8oPwGE65t7Gsx1j1Z
EJwHzZwcyH/iTmjnAFTp80yOfzpIe795TYk6+rw0Cc2aef+/oaUSBl68jbHRnnRz
afhdO2qniucBld99g9FdwhAamtEPlIHZLAVZvH9OTxsIYuzGSoyQ/TDlklKms5bR
exiCZR2Wlw993uvr4iJrbTZAtW1aAvA9KNSVfK4cKSp8z1qOM0nvL0ds684l97Dx
+cPBDHMpCsjQWSkH7iKHOJiMmlk1BviZ3lRu3NMgoYTswNPLzv0RoVzJCKHtw/37
h/QncS+2RBuxnVkYG3WaNxL1Jl6Cr/8wjE0M/wnEZJvMgETwCcwo7/iv6yURbyke
UWok30OtswXt8ZRTqPBX6xUxxohBCSYNR2bNTIf+1emYDHmZZjgB/CddA8wkIOAp
7PvAhFDTuYi15+FEt1w2WnIz5qYZ1f9jjPghridSlBDBleT7aGUmZ2bPAfxXFPWL
BTBpw+KdM5xduLq4VUO47yri9Uh28ob9rIKkn+eFDTGrxz+njwsccQcZNx/6odZi
/ZwRHK82V+2/Oovmf7fz3IMQLea0pIyHydwZYa95fmV8/AG3FaC1L1m/NUa/iX1i
LA2NBvZ0s2LY6mGisNyfZ7lasl0fsxsmL9tTZNxOXyW1R9Zyudn+nlyvqRxARXOo
oxD34ddg63BxXmZ7cPEBBkjIHB+xyAXmSTPeISqEv52G7pbdppEx3Xg9/ao6FfIk
friFjHwZR/t5xbcZbfnDBK7R5NQJhgfYJOlRxKRfWp5dqHlycaC4sZa5TKqzRo/b
cKr4CclP4cZ8g82OSu51aFEGGF2XyrEyD+OwzhaXy4OtODoAJOXZ74XQJPWqM80E
Xx+UrL3bG6kW0E3gP4rMzseMLmXoPFcPM3O/d9AW4b3i5UyoozYbYmzIpUsKwRWy
ADjSfDcPOqR5v+36rUAt70isVk48UMRVM/vvevrNe0B98fMM43XFAeEVxJpkX9Ey
ocL+OUhpZ4XUQ15+U/hngUJdjpES/RhzwTSPHSf/lXzBaidF3aGchzITHrjHP4+t
oqNEOM59L+Qsm/Lm8C6GqJK32j7nOdHz+YeKDO0XarCPc+YIfAcbWCekgWJlRAKl
GAjQqdPL+CFPB0zidKcuOiTRhiomyxG9oZWw8MJwplYVXUe+BoXtGNF202YiKayF
COp1IKRIK9JHCtNdb2dxz8nDGvmm2BS216DY962M57gwz8yKD+sf5r/Z2uxRFYT/
+q9HS0C/9W3hCdNeTp4R65ms5wzj6FxM9+zmy0cIwh52YK4Wmax2xn0UiVR7BOpx
IT4sASvRb5r8qkhurWh/Vd/2VrAR49pw8KVowkCqqpSTAv3jSNPo3ppOLBsgq/7o
zUKXT4JQN+HwNEG/IvMJdfb38LEwRZM1pveCnb5rTJzgoNGGnxPA6BU1/1DSZPKg
stxt4eYStq5J3Ol6R6TT7Yk3FxByYGVmC7nD30QVhvrmoPu0HfavRmPwEkS2b/wK
oAVPy6a+Wj2095UOJxSt9BpU7Ju1osGT3dGrGDq0yvyJzhlpzYnIEgmL2+ru/ojO
AAS+XUGG5vFxd2EAKEW1eA7maBlWfiyAFtJaxRmkUQZK3JKQpeC8TUvg668vUJ4g
sLORgakuxHKGF0rS3W5kf50IsVv5K1NaqicGKpGP7K79uMqtyB2LlVtjEXsyU9Cl
RmU1StHrnTpREYUuCiKHcUyJLWx0agdTsqMAMhlMhah/MmJCshTIhQQL8dBtSudW
aaA9+keYjkhE+dwOxn99hx3Zs0th15CVGIAJqH51Edmo3OYN9vtyd3yMkPpvioGL
DwikT4+zh0FS5s/LJfOIjm1SdpJoWMvG01xU6EFZw0KXXAriW5IKeZLB6NrkMssc
OIbqMztiDBnkd9p/5igLARol9u00w1KWb8bTISAUKNXG7QMz7ih/04J+nBQdo0kI
MsF6492F16aWQmiNcy2AHLwMSlXiR65JQp6Tiqbwdc83r6lQ5/8Xvmc3/04rBvIg
7iX2sd4syFsHpZ8fMs1LtEdHfDPTJTb2QEnsYH2UnaZZFa9O0iKU3UulXQSGLadW
kYcWZxerrOjaOu2wLVBLfBIgfyZYYcSOk+p1a6cArz/MsdhQiimR2G1yWJfK5mGD
2V7TCYCfIJhcg17HUhvOoSpf/4mTTPwwKkLVn10rqnzhLvsSYrInCRvthu+EhUZQ
4/ekedAKDyBYMOGKywNgV7oymEHDl6UieJm/9KyZ1uS37Zo5gu8djeigc5c7v4ht
JQ/BSAH7So4cr2w3kBy1kNUdVhcv//Hg0l3iMwqWD4gwFvaiT1w/4gBNnS97g2M4
r12mhcbfClhPBTzJN7lRE7mBPlCS8YDMkR5fKFI5P8TBW7Rz7vqHQIdNiNC3YGRN
Uto0KGPNMtf1tk49OP+I3/Rncc1oHCc658bEuN/VJkHwmz1oqvkOJb7X3/0px4sT
GHc1nxvpTpU6/emH0WoTh9u1ilWA/+u1rw6gcPtdFQ50OTmH+TJm47/r4XrLojGM
3fJKHad+ZbQKzrimh0SDg9unEub4+SK/cYOPWBzD6NCjLNyrbzl7OgEBYN+Dx5/f
ICe/sI1KWf2UqNp1oU7EEVakhFA7nz0UH4RfqE7xs01bzYM3xns2XFyP+dOqH/sP
h7eJBy7ARCEmo8RB0YbxXp22XXieNCamm1M1JFstu60Y2UsJWeA/yQCVzFEt3drg
eO0Mv2LBw4c4jMt7oAcpjKxk7CO8vRHGQ815LZ4awtOCZblV5aM6PCL9AGMW9xqJ
n+qANOhZPV0qXLhNfzfReJSqZEkTBKtUnnqYNjMHQIXOe9LqhOsCP/VAqdnr4Fna
4AqP2uchBndygp6mtVsH0pdX4xiiD/2WhFZ1SdKCu8T3394oSPUdn+LSYdCtTL/S
mB1bvvbqvQgSEN/8MigMljzvJwy/8mIqxAHoTrHHoz73qsF/3cWLXdxYmC1uiwGk
d2X+bcgJP0+dWbVsfzN3p5/XP55aHKLkvFswcfu3xXcYzGUxkOZbp+ZHCpy1gDm5
wG9BKho3QBVfoG44Zu3TN3aY7g3ARx+CR1eWVhZBLYMkDxY7DSoQG8xGU5Vu063W
rkmD7JbpxIJnklIBzKPoaS59Zm9YY6Y6mxj6scvnriwpu+JJiUFc0sm9WvP3XIqS
g022HGtlvvkJW7OjgDyfdOFjmjkXLsMJIPE+7A1jNM8UxY3INh46ksveX1eOhGWf
GoEhmZrLIHz1ng3IAILIVLzbTuDzKXCrRxRDl+jsvDXMangVDIcmCRbFRD9L7k+2
AasowHGVhHli/9qeo+n/tPXliQ8ASbY7H4IEDCjLE+MfdyCLjJ71ByEg3432HsAX
ZD/binWPfuLKPik+psX3d7/9LvS53SsP6BFLPcmu8SwF3F01tOdPyWdbWgRmvD9e
jLyvEmt3+s2knaAPQaiaOYafxvB3PM2pEdfFB0hz4fXue40qUOtB5HzZrfiZFZXJ
DPv4skJ8KyyIkbnSJQdHEjzosCSa7kA+n54fsFDBuFJFgFIIEQu06aMc8Ci0JzVx
+rLOBBUgEMo7KcwevQJmLAeuWo7LI8wmT7+Tb9nVC1jrB3s2wvO/WPpEL7iIQtDj
SP1+QptwmTVapxNb8i9PNrMvsa5Wh/ctG3d1DTj2oJqXsZg365NwlzKH95pXQuYZ
/4jmE3xkSYKU2WvvVVBEEg/7NmAngB7cR0QjUS1IRYVJCq6NtUVnh+PGFZIqI0e2
OyC1DTpfaVp43mCUBrzpVVRZvYEcXBV4Dn2eRr8LoAXcsiLT0szpoRWF1OYq6Myy
9hx7cm0Se2dG4eRgQVrtQXYbiu7f8/DbudLRCsaZQkMc3/9Z6r5Eign6fJmgkCNo
W2pi2leOd0p0SWMvTmQtxvp3cJ60JG6+l7thOTd5KRrbu9UfjSMgocLqf+3/h6cC
ouUxB6BCAQiecVCHi8VbMYPiqL0CGTdnqibM3EhmjBOLS90C62jdVWNEjeg4TFPo
pZrJQWrwp9/u5k1JVAhpSWAmIcx5dKiVe9zY6tTB8LF9mimpaETtxpOeUvviSGXK
yVoVxQ0er/K40pF4vva2tbjcfxUCNZI9hGZAHOrawKWDyb2kaOnfPtyOTD5oX4D+
ovt/krkQxMQUUAqVHbwYKEfqK1JlQE0wsh3ZY1aSKvtrrE1TLYS/Ck96dbkGEBTB
Xfi3XOQ//vBrXYbVUjP0qtKcrfNinKBJbO7TXWNYuvWem3+Q2mvREBGAuD1keXpL
6xPvg/etT9OS+h6FkKYTK2FzTGfO+rWmL+1EHMmCP6suLt4LkmsEFO/U1cVj8uKf
7xtPevivRLNxqSiGl25xZUy23B6SwNMgeaT8k/f2uIaP3ipr2/ZSfxgIYofRcusG
9NZgz8hu56BXDGNcJrXzFDFdMPU5cUOQfB25rP7w569c0YDNWFwG/HP6lpHFR7fg
TTesjS44doyN0c/HUNBcRyNaVFAHbfa8I/J4zAxRE/nP17SrZPpesptqJaDBJbLI
8lYtZ/xp3tSgYE2aL9MLnbx0Dft+hY4mgKy9LKu7IQjtgaUe95fKNu+cmRowq5Ht
eJk9mx3IRTNcKQ02v2Ca2eD5sc9eilDZ4ur7KSMzajgqkWLJrfkXUK4GGqjW4FJv
fTnDZ+kC3wVkZgEJCoLqHxH8rR0M61DaoQYEpnA9OlcUE7Bl1ZMM9pnI1fuMrSv+
L/KvCvoZ08BiemwKEdP7abrQ4Ek3wmJHHFsXGbhlXvPmMuyuZfaaUzHeOfFJtPgZ
0XcBIAUrxsw/dR2esWmJrSuhdXfPin/7X+i5xe8tnfrsvif3j6Apzddob2kFxtrn
g4UFaGFO3wOAtuSACYnQ19e6ydgAhl79TxBlpJo6NcV6TrcC1ZBpdC86uiEMWJbb
aydgtRQztgQD4iXyNGdu8U1qRr1zT/ybfsJvmeN+JLfTb5b93SRhiaRvjZ7rwP0r
f0ffvId/bR7tMpa0WHvaeQnIvD+4/DPDjkVN/od2sPL3xpT+0pWILl1LTjqI6FQx
RIhdtKCh+xzuS3AMX1XJqotN1kH7JvTDugyu+W+RdRjT0x1fWOJAlQ0P21LrIMKf
T4Sxzhr42UCflFZLNS2jq6v3GGxBX9hbVLiShhsCVFdAfsx9DOlGRRriuSFIbbXw
Hw06PM/95rgG60rj3lrH9L3hgskq2LswU/Tw2c7Z98U4W3LcvRqesZKMjCpfeAJe
EnB8CkboE2i4OM/0tKRQ4Bi6f4uJ3LAI6O/Bhxl7PtOzsT05aT142MasQfwhvYu2
dKt1LKk8ybr1KIfTlApx99nHknfVleChw7i2krqS3uz0QXIyZgKF57N+aFeHIf8h
KzETeY/QoAUaNliJea6EMS+HEYk0qMHod+F1kj83Pj+55bHPQGtFaCw17CxXdBlK
5ngiFVHklbW8vYlnJhrV2QoCAxoV4dgPbowEBju85PQcN4G0xU4obG7LlAswaCQp
FGozrmCvk7ybhGipYloKTB1xqp/6qIV/3oqD9/8Q9scfaWpFjp42W+VNC4oGs3pv
knj5ARrYCcDKJ/5pusrotSewLDmQJjHqXXO/k42HqGGQ+3X05/5Q1BXeKex7glKO
rRJoM7Vg1wUtrUrV+NPuDakbtUjw77pQWP1RzQ+jOxKWDrrpueFxOIQqrrJOjoJY
iEU1fsdOcIUBo98sULDIWZe+v9Kc3G+/05Cd6PxIgiejGXoQIkJrTZhjs6DjNE0F
gTZUiK0PFZTNR7CZ2PrbuAnmt8j2gyUsMIyWMS8n0O9MZ2/w9C6sVGy2HgXW6QPY
HVEBmu4mzzt5xm0RGhlL+9man9lvSvCEP2AU8HzSENSk81gkWva+33ieZbNK+Zcl
ux0oEdiirtCKo2tlWQhmGLNF+pjuWuIh8dOYHNNrSGtms6sPZGFu+kJr4+7CHDdg
5Hgk9/wguYqy6lqmSLOFPwa/Oybls+9XnxB/rr1EHAvgeszV1diT5OkwN8IIQxQ+
eaLSwgzpcxdStJz/5efeZdYZ6Qx4k2IHMRdOBkfK5FGd9TWrVvbDRpWc1s3Aqy/d
ub5NlYldwd7UickVieRErw6l6feT5zBVxKOszwYWlE8LUNFKtK/bD96tFdpvevmq
7tnu3HpUi5Nw5H6NvydAaWNJx1u2y/KfSh4SfbBYP96lRa+6RPdshndKjGIr5G0c
pD1g+1p0YfkmIYrQiRHBMClBjj8A0WPjHeK7DOLEgj4pW0gpnqyj18PP4Amt1Yl0
t5+PwSyb5g/9XSfPTeyX48INS9O87ImezgB3q2FkhjTdoafqwSyVAym7TvSvXuPH
Ui9xcWnfBtWWFu1LRWoXiW4GMF4Runl3bmv+SpZ+YLPDDmt/9HfHK2mAGwNnMOXE
0Sm4uUiUFg9HRY8M/P0KxvwA+wAD461m5WA85Mbra6Yin5xjT2AqDCPAdvwanZKG
LysrPg4uRx7vo2E5eiJJXu8geS8ZS5IRvUw7WzaIPcCpJxyRz1xyupPvv4lgFegC
R2++hV9x3N1SLo9/DxCNARr9yvbxMq+YLtp+7jr/uLiFXFQyYGIf6nxTM9Z2Bb7z
pacQnd1t9OEYlKtzYDUgNm3JnnqF26Ect2MfMk1iADYBfPowyw/Sv6oy4Ymq4ktB
MBLiUvnzmIJnM+hrjb7z7OVQ2BZg9FKpok0p4xWiKZzcLaWuwQ5P92dlcsMKZRcw
EiEFhI/mKBZ7IdHoDNCJv34TwWotqT339y+oyRxOgRz7SPTyJ9HPEPzyBGKh4XK7
32sYGb0Oa/keJWJWcQZaKXXeuhtFUUat1glUh4LizzwJL3eL5nVhzL9WhdQZJD81
2C6NdpdaIca5btGjdo5bNBaZP3dHje0+YLRW5KhIHQfKA0BxPr0tJ2LGuQPhEPz3
Bk7w2oKWUclZjHi8HYS++BSZzsjzeB9RVA/9LHUec9kBBpfZtwtZCsKCeP9d/7F1
Kug0nPdKEXHxMEpQiubOjes3s46roON8avjt5gJOx0DVmjEWAKrtg6/3SNKst+LZ
8eczHwBX8Fhx+FrnZoogdBXjt0BK0HXWjyt3BpkxgeUYqAxlO0AIZACex1dwBWPl
mRt/EfTZbT8/GM76PopD556uY37572ALE4nZCo4244EM5wlcTXiscHBtgSdC9TDu
wJ+bvoZO0SmLoAO7VxjlH5+NB/cUudKc/7q58GZOJUN7E09RzZCI4ewpap3WYxBT
wiGvIR/ZFhp/T/DDEapvaAQ5tPANCcmZqjIKMMv9ovZbjiC3xcey2kDEHY4Wqn8w
4jgoFJUpayX7Vn+btCceaA9yTL2ho8DJPCZM4QO/MTHMm9Lq5aaa4IZMZHvEWGHz
RHZiJCqfAdHjGYR9aqnbsxpyxmpwu9UYcIaL1ad7puTU9PRn3LeNHNummUhVQhXY
WwlQ84d+3/d8627A1JVzSqIt8qFMJQkVDVL+bAvHKHhA9ppWGs1UUb7rLHXt6a2O
9RHU6ZRI3jF5hANeBYYTrOpTkN1iufNrw7ITjtBJpRvqkH430X8fP2F2jKFlsnWT
mkxKAiMs/VLy2yj6WqtONHfmwdnNExByZIvI1KoOZ6KcY2+P2YQzUdv73BkPdDyw
Pxz9kc+DhqRnvfWOOVQfzCxO0K5UhhqA/tIfUZsV83i++So9VwkIEu0mdpsIVqHq
Q8S5ajYJxuy9ASIqp8u66esSIEMl3qvmi0dXkwrTBRP+vIVxvSEN6nzsoesc1/m4
Tz84K+RH7A2N+M0IAmEZQdP9ff9RhQNMFQs55oQAFwB7lqD8j9auH4Okh4Ms4cyy
LfnwxTaRn6c5gpToDvJr1aJEh6Ni1CaLaOcKZjJxMPHUl0bhdb2cmC9j5Oo0kYv0
fYdgREqf9H9E8ECpY5askROKF7fKYyYEfYIo0s/abiJ26F2CmTM8ZEJvdaSmRzOV
aroCgGhQMbvbNQf5kaLIcT28if/hAv2p9esTeUN9Poy23gZalUaQNVXOdZXl+CK2
lCTuFoMbrtKPv/ApD/bcaNSJgsSirXk1OpbgEhkscYisDibp6DEMBCXg3hXlguFV
K0MkRYPpKs0ZS33SBNZzAa34Z4yopkF3WUEhQfnZ4S8csrSBZQMHCqAh6b2/yApr
6w9eXZPT1WFCj2KnWFVzQPi97XLwTvhFadj+k1fHzA8D9TmYySVI/piMWvphaHn5
u0r3Nc8rbWkOEFn7jl5O6dQ71SwRWfBsiUHwq7GujKHzPX1wG+hxcsQLY8E8tjZU
s/EGDVZzOW1TiBU8Cz2CjAyVzEwA4S35Z6JW15E1wytwnOO/aEvSU1R1uy7qzmzf
ZKU7khyB3FIQbcuRd8epKODzaumrSNxcCsO3nIgDNo5A2jddXuliaZGqIOBkf+sq
2Nma/RGkLdKH1QLRKWfT2LwofdDpBSrr1EwjhqfFVP+CCMKC9pxHMVhGkmp+DgYm
BaEKMGQnKxQeSpRXcFCFdE089BGZ5YFv4+z1CcMBO0CTlI1c8HGiA6RNoz/qDfV1
vX9WRwGXtdyNWLsZoroE14Qf+aidn8aOfe4zkkKvqbs5+GSooop3jQlvV248Nfzd
93/2i/3/N+AAjXw7lVmyO8lvYf3XXm4Qv6HVeCQfD0swhltt+iBAZyJwfxbBu3+m
/+SKIrVIYerTYGW9GfpcUAsckK+TSVFtb9y2dH9ALN9inEscI+q1o5+vUZZkk03J
ZeEyeU0c+xEEate1mbf9gHBK/o7D3dwUsz+2fP524ZXm+i0B3nm+DqKXMPGHKYnr
DTV0XSb/9E8iCI/0leUO1PDpZ6IrT+L/+Pvwt+7PY5jSxCZAe4gWimeT7vLzs6i4
mBPxleg7IoPG+dC1DiUt2Ee9sT8ATMt4z14tWFaryOhFsPvqpNajBox4tX5TIEbY
AoiTisFkvgNhx278WpC8PIGLkYohuOczM8iRKSVf85QwUwqA1YZgsBQTpX/4Ktce
T8n+h4Y1MKe00OklH6Dl4hldTygNQzc0oGGm5/jJYt+s2iZ1Y5e0u1OjIH94NdIj
KNISQZc0eC6AViBUui+MMykI5ju3EOorWJRTeWbH7bGaCYJQ2+Be2/EZx7i8CVuC
XNXOqs9/d4/hw4BCLbVwn6z7uGFzvHwBGd8mvYvOo2sD1o0luB29cJly0ocA93QE
Qr96Vp90ktrULdz6hG6KM7rUqdfI20DUSw3Qp3ggetLMRzklaDEuckcczrp5Wp6J
sc91l3H5uFAlbYoZgBCme9LdII1XZoRiajAqAwChD1gzw4QkdKkrgHQMCsKRpCXi
ifLvybrDssNssRDD0V6KIrMDPTxEmUoORf6nDbYYs1U/UGHmpnFsSy9Iy//cOWnB
DRIuj4TeT294nfLf9H10DesNxm/McLx/3Pr6rkWyAznCJpbxeV2yhYjOa3YTMUMZ
yNu+OMhDYQQ7fSD84M15fqYzvkO3ikfb5HSrdYau9xohlxhEKkU+F4xwb+am2NG7
Dab3bKE4/fDgwpBpO00cz0JBtUDMrBeK4/dBJntfR1eylfJQDQ0kSRBzf/Xz86OH
4lS6gcJy4hado+xG9gAN81281Xhc8HutZOsyZ/uln0khxsa8plfeCH7fJB0EJrUG
HWz0VMCPRrPITdIhMMYE03Sy+kcbjT8pATZJEiJbn0w7W/Aju6iciOdMYxqSPila
jaXsRWcOgG4K9SxMKh+sE8BjSWd1EdrOfjwVAYJU7zvm//ER+MSZ9iprW1h8XrbY
1VFR4cckv8JNOCzM7njdG2hpdmUh08QOcUOFvk1URNSlFO9/y2OzMN4jRxfy2DCz
miwneI1FGi2RtiBcz8FGvPLkq1NuCGh/srMKllglPEw+jH0fnGdiE2FUWGWf1Jdi
0rG2VecjWv1ehtAN+zlaA8aXbCkC0ew3hX0jbiES+wT7fF04DJGa8eH96SdEmOFe
QBXB+EoUbzNxS/l6qFBCZ7ie3GGLJu5oWvochZlVxEz6LfwUEAL2AvwR+UPzotig
7w7PDScc6vkxx4jfPjiz4Luy431QYqkqBi/gOqH7Pr82fstoH4Fpabz01jLzet/8
sFv9xDLt+GZW61Oz/XW07jRlzrPmijrmi36odjnaVlT+gaedl+ZhLoyLfDJxiMU8
W++baAjEriiCimy+3/rYuM7YPvH3rFLrHtGCxWKEI0KCUXdv8RcYVAc2EGfgJa0d
e5ZhW7Slno+Vq0WJYbYavUdUXBG0Fae89y0DNkTiPc3CFbJO3c2dOKwU6cLDQZ8b
XR3kpbIwTYsAY3QzyeavBsU6KOOinv9i389lXQ9NJdhKeSydszwF7pV4MXEh1M49
19j8ttSPbvOZsnBglw06/zBUBTJeCH3fsM7t5OBitU8q+5pAlyOF4ewKCQM/nShX
mDPlthPdNtwoIdCCwP0G3gdRnPuEBkFPKIDaEQVUMXFaIXh6CTVYCVOnW8gSNhDp
q0Kj8lOzMEJ8RBUrb1EaUrs7o5uNwkf9q/DAcXFASBlHBEgNDajVHn3vxOyDlS+N
cC+6aqDNya+RJYy1wt0SeOSd8WfPvbMQvJTYVl0mFp7IZuD24YkFyz5EVMXQoSGR
Dy9sYK3I++1Md8mw/wW7DX1PWm7CKxWkN1yZJ8QXWpNAP0se7MQbhYxtXWYX6YXL
OWu1owEQr6LW7yYLBCIDjc8Ve7iZJ8K18df4e17yNyfJpcUByZn5SyvyHUhvYVWw
HZZwuBtn2cI4GOfrCu91TMAbQ+NxmEtTbcpqK0d4bQaSQV7FGVDDeGekf0wviv/4
gG2pqI4yw4LHEZVzD9L+KE/jI7/R66z+IYkpZZ+y4PSx3ZCg3PLG73Aof/8s96gl
n0f12eRKer1RIXdOTo5vvZW/O3ue+1WBLikci/WTmVp5W84hDIo1O2mgDQVAv78z
tXS64aJNIc5RjrUrlYX1CbPZaaMY+xYZa8c7GNwEtd28DQxWDq8XCI9LNwECUP7n
HiRfxmScnQYaIu16Mr/oXCy76pNwd0bqlSEg2QoqQYGRIE6rR7vCVRDxhowdJC8N
qsp4Otlnlf+P+v9WknPycjPrwmQ+G6WAeeteV9vCAyPxVysLWfF1Mvr25jxm+49T
p01bwSzRODh0+IAdRPBynOR4hT+zVSkDkAoQgy+hKFY/pgIi9oy4/qrGYNJ5bBJ1
yt/qXPGF+fYr2tuIepFjIuhLCZcZfJiMWjyMeMag1r1bDrN/5nI/h///E7kK1N/q
G7eQf2olNeSfLDvd0DFcL/PyupulMzfa+WF954BRyGfRtQxjGXBlrPOb3eFyi1jC
ivg/4+760oc/+iv+PheCwfY9HlgRouT9WUxWWZX5c32q4CkqRaYjdag6HZiOaL8Y
M53RWZDmt5udJCKbAbbtj4Gkprq65/UPgnpmgJod4Zlb3mD6284+5aZ1aF46m89C
Mx9MycN8SjsFDEsZUigcD1FBuJkgKRZZnfylE4DTghmWCn4UeURFHF8whOs7yQcp
3H0ZEAe0Am3X2hh7K3wyaT0MwkanXj3505xmV70NDkyICIEUdjSUJTTn7IyaSxdY
rhq7+krIU37Zfit+mQU9EyAobbaSxDvmci9wozb1EfP3efuUg4h5TsriMnkikj26
nIPzeQVVlLDME8WuyNWPu0ocBrd3HFN3mB3F0RrzOWPy5Z5sGsJwi/YaY2XACBH4
Ui0qVwDZQmwNvFpeZ1PGtjXrO64YLfM3AIooTeC628MjIi4wBNwvOPiOkZUSkFTs
pgL5YdeFcBLoKY+1beb79zD9cXJVav2lEAupuFCuykyjhzNb52Awjlo1dos0F8hl
3c0HfEc5/Gxi1oWApApkHQoMYg5myHmtmiU3w+SCMal8m9LPZX/DcggKSEvlq8if
RKksdrlGEn0MTd4SxbQWXInf+VzzmJHY3PUXt1a56KhVVVCmecgAqmYZ3BRom+9J
JlWQdq2Z3Y691NcOKtvyptBMGtFOAXMHhuCj5Zhb7TZXf+5Md5/k0/RJSEMMlls2
nQlT7WOSUdSa0jlg5xdsLO2ya1yRtBuGu4Vcj4RrEAcln2ARMpMeZLgV8R5VrlvM
jYjg9w4rFBPf05IDL8gs3UukGcjB0FN9j/SWfF5dC2b0Tes2u9F3MngVscuESfhS
MK6xLaOP0+tN7119L4ohP/rDQ0r4O77Vhyd89fepzI7K6ZJ8IQLr9iN6uhPe09wP
CkJkkgwHFmoE/xUSW/2pir+aXsWl0fQOdG4rwTPjFvKUnQ8f6ohh3xTLia6TtSZr
fROkUHl9CLhxNFzftmSsiADKhoYyRJR+gek/ziJxB3aJ2HUBdEUgY3DCiafaOHZj
7vsNxOlszMr7GfEPHhSzUFT9jLJUojbSw8NgfRq22euelFu8+02R2Umoz6Ur3Zkm
kUklKNkZ6J5Qiat9QEDpEdokSX0RSmGjNT5xfuD23gzbh0T2f5I9BG8CL8jS0hiM
WKwed3z3s++CusWBi9hR8/km0uNOnAp4FnRfvFaaTZq/XTWD/jyAWJ4djleNR6VK
TTgu8R8Jzmdo38eokcAua0WD6tnjox+oX8OsmWZ24sX8uRFsd85SNy3kCioQ9awO
F7eHclXzFoEoAGkjmMaj64BwA8E612t5vJOCaql8eR4nBnq9TNA+biRU4y8ZXomT
ibFiJZel2K7MUeFBTuoSWxIer3V8zQHsYVlg3XPw0ph2o/3Gk+t7SXN61G6FOLjG
41qyubaQtYRk+zRAR6PdnYmDgeRoaPuowmJbJWE4uA/oPdRzAbIkFFutumYf//pq
btoDDpZZTATZdQgV11HEPY8LqKiYRVPeFCs+dYQXeliUU1+elOub+GkjSFA4oNHe
or15ovyJOt2WqYqCcfujL9AtogH0AtQkZaI5oTHNE/NWkabnkV4t3IMApS3jygw1
7BImsqPe2UyfSc7jsLE/jxaa2UHJcc13S0TL6Emrw/3BtZB9ntADl/ATL4Im0+1h
ICaMv5cGoodUtgty0oCAm30nCGIoXTH4wQyDvMEMQUgWGhTAiXvsUGzcuSovA8Hx
FqJVz1yf63wNfSBZjtPmdt2MJa/hDGa0Lfi5+aLbJZ8BjXx1XKI+caq0eVb7W4fp
dooIXzB9xD30wq61peUO1PIcdcM2zbynC9tyDRee4awceMaFuYFEo5YXeQ/lPDOW
KUjwK3emwVtkf9fp227I/6cIfGZUQ6uqvasemIqe7UXPQe5JVvT61nHwFN7rBWmZ
jMXlU3TJC/xdnyYlGRl4xmWypKNSIFzY8h9b2kH1n8KKzjjlTxjwIEN3X2SV8OZh
CuUu+Pf60iNbyb8i8NPaZyZgwHZL3gvwFOTsTwXlfkFA691YNrOsxeG0g0/IPNFd
9ZW836Njb3/K9sqYDCLwWnFryiriUSgMlg5m6XZDSiXpK+v41nNcIeEuuik9yPZ0
bpeGSkAKQSWB+EZiNB8Ry9kWZLgRP9iycCnlSWGoyxl+Ey9cb8nGX3pRRwQjLJcE
npYsrBwgr3qCBi3eKH6yOBqKKRXSxkWg0jfCksFbsdSZSKgwzl7V7DpGngMwOFdy
7ubQr29gcZnEA+X91vI4RY95QuP6HkMuXaNs8L/TBqvomrIk9fi7O2EQBrSkmXyQ
eKpYA2Ig6xNdAvIwTrAvaOmkn6x9JLcZSs5uZqbyHB5VNw5pAjAl9cO+0pAPpjB3
8y3B5AAMnT4dzuClbqbaAR0tM/4NNFyiFsQPEesgNYrmQNNlJ3X9OK9Jr4NK4uXR
XdxhQOHP7+k+A+f2nvkbh9QiCL98nWrzgl9fdUMDlQJahnwidrw30HCRLqaiHDOW
OTIP9JS4uVGxsG0dJWWcw2xu3ffsigc2nnyhxkb4OIZFAOUs5faRtAedcwliUaGk
K5dBE03W872qlQzwRwyWyQMsOT5Re0M2Hu86nnmAF/qqPA0swWOjw4GFd0IOOZpq
iQLp9Z9lC4YMulIJm4zW/d/09SloPgmj0oZC67L8e2g1XeYo8H5ZoCOMMKW1+bpA
1Obnug6jwnyGkz9zX5MJw14y0M5+8x/+pGjOM8XLFXp1URTS/g41xQkwKb3Ss1Qq
P98atMPMoz3MMqmaihIVEr4Y9w84yVE7ucUKKaYdpnaOU68sdVM3YuiBzj71qjYF
iomplJRMsqA8fzysaO1zshxN7jZrARAIgtMUkcQ5bjhPebRqAbdRa38Cv1uDaF/M
v29NELW/4Qg4bYfk8f9ggCNVbSKf5Dijgf8b/Zw1gHhlDMEHexSUzmJgTi5034ZV
L+ZWB2ZXLfJ3nsNYmg86fRxaflP6KVoshRa8xJZNmfGnKkTCXJ30SGqRUPeVzvNW
yx+AvGHyEijpXnz2TFEXGHerdbeb/c15NVDm8YJ9SVyWCUktUfdus7cfGlq4a760
DYjdb3cHXo9TaTt4mCydU5M63DUVBy2x5DrjvWFuQRgTbcbNzjkq197/JTx1E7VF
O7iPJdjogCif2dTP7d3p5PAplbqKBtqZ4qMb/EajOqQZBrO6oCtxbsM9rVzN8vxQ
LdtK5L2Wng8XMQ7jplvAtOzyaQgBYk3hELkaBZzU8QcIHnFTEQ8t579FNOQngcI0
orin229P1HuF6u2TVx0ltkQDmEFJoHQz7dZP/GYLklJJLHCh83SNKtoMVCiJvLez
x8KSB+Gi+9HbId2CHCJaajEp6/yCtJVpWthf26s/MvkXbdC/qEgbXHu3NkeRVZbH
/x2qz8VOiSN1y/G2uWVaxIjY8XlJzJDCZhQ3zddLShrCpnibyyqMNfNA83gay+o1
t8gC9eSRWuX3yLBs10JnnccSxeIGT67pyzAIjTj9DndfzN50n26kfmCROn8e+5QS
6pw7k/RyQq6yFsmgSugU+C7fiK2rGpNqCi1AlsBLCX8MWlX4MEh7ygjte9xQp/it
sLfn6hpw2duoan+SZMWWOkqWt69H2sKcH3rKgevhjr8r8RHvwmgT4taJ359dnlyP
2/pVRXqdOs1VVzZMkXt/7tiXMZIt0xx0/XUbfXxuGTMhk3JIchwr9eQkIxAKM9Bs
FjvI5DPIOH6hfGzWU6YQKl0Ng6RNwqrfoes2azVuQHDtEvQuKzBNdT/+NSWEzoNP
S5PaaHsjOfSnx9j+NQSKae/E7hGfG6I90DgZgSA6d5z4gfjmybXbFmneMYI7IGB5
k7J3gX0zsN8IzEXjWGceLPKbljS8wYd/6v9+/eK90zpEGAtYUlfdsG/Q/8pVk4lG
EKfEHggq3yu4X0lyALA+Jl/LlfHbAzYdxQBnt3zA4YsNeQ4lZvbAq+yekSYFXrym
2waE7Qc5/XamOai5o8SAiA0tY1dqSVdMw0Ja97AC/JJknCoc7lkomsjpl96seU2T
FGx2jpZHRPm0usFeMLRSE9djYlDmhBpBj8kk/ovmPNX61N9hJvEZgDugPvv1aHNM
/elOK+RzWYPfWlg/BxSqdA3Oz4KllbaP92HMMKdKpto3qC7CvSnsBAXbgDURAXPG
Sok/aQP/Km/BoFi1WqifWkgkTucXAWm446+btE3ScZDmm/PZ7uK9zJYa0E0868M2
S8+IhbBZrrjTAFQ2BPrOOybMZvuZI07vnEiEgWSbtfPxjcKHlAcH65f1ndserv+W
GKv9DC5qtndhI9BC+dYBEyUjR8bVnB+CjV1E1dW1JDPRIK7sE5UwfgNcxK3SznhZ
HrwbC4vbNQLuj+jAmUti4k58/nB0o1mz+HcRTSvkQ3potbU2hKifu+dA0hgOS3Y4
/Mcez7is7BIpylE04llfn+1Fvn0FJC6HvsmteiiAcuIKzdqYnQgfdpvKVWMbYH7p
aNfUHpG7JPT97eCr1sgfslqVU6ULV3gSMZ+OlX8zYDmp1V1BOmsexVMcH+xuwAwc
ul9akcDSZgnOv+KpZ/VaNgmy+JvPykaML46GGAX9aN1TvqgBnxG+v0EMevQVfCq3
7potISE9JD8EXTbBtr/0AwiG0RIL9Yy1KqwKtiPyLJkQjJ1/LQ+BFiqpQyAef42K
KYwycEfhEuu7N3Mpqws/FyGtkbU4eTIu/b7I4lkuNi8ep4S9sPM/4/btLG8iT/sj
UtN67d/8avKv0iF8pN2WXJ3CwZB7VORGn2vo2CTdrjKyXSBr63Y3/fmqW9BaNk5r
scUVBwBKHg8vx/Ezsd40SQ9x7YpHmC3B0nUeEAUnJtZEY2g9iCMC9eQXO7ePiU0X
jRdPiYcrRQgTii0rxDf9hfXnhTYXOMjE2HCAKREs0koUHqf7LS19nwf+Ip2cNM0L
Id/XSmSUUZaAS00rHeXDlUnt7d9bvl7yI6bE1anWsZOnYZUF/HCSXFy2XbpRjbXt
+ELdPXjjDjSZ+EcnCp/eFMczg3gL+YQffC/8mB4hViMdSg02x8OpXMnTzwSHQfZW
RP2NazQb5WUOxf7+GadzAZ/e0nKVdVGdigLunO5Xc39OmaDg5B3Hq923Q2gg5oh6
u1LRq6zE/XBOUzaQc6yFgqcOmyy3+9RMWOERlrFhsG90G8h0jOhD2+AqI0AtLNr5
Lljb/Mi3B22bc3+qXGiGOR/KZMTm1VDs5oz+BMdqqPKuvjAeB41OYaUDPC9wY7pE
l3vQkmoRSmFLwl1U+liUAjEFdg+3FsnUCaTfAWkN+EmVmvwPaT2p2TGEMnQ3a/Qg
BMCwxz1JMBzxIvY3VBDCveT4jTfJXeZ9k5zzSuNyY1ot6Fe0eD2dTqCbMs1394LT
AF9/z/9BzQqKx8pfWHyAryg+55hG7MzWqC3Li88lOc4u3QElBnCiIgOtQ9UtLtEM
WMomyW4DdMVwpD7wiDH0NLJXJ3Z7Lnl7DUXSAB1KIegqqoQy3LFV2WOPY21Og4oT
WWdRubiIS4y5dntjm98SR0QSDUeZz26LPLpiLwWRu5ZOmFLerW4jMLF/Sd0RH5vI
02qayudeqQin31Xt1zt6eSxblvw5XG0+UPMRT2Sshm71l/qOjckURi8PppwCwoqa
XlRH3a1iGX46V7Jxy7FAUqlWbdfSOcb+xchgxfyI5GPw1REU+hki93Xr/ad7jXz9
UGI0kDx6sC2ExoA2SCegbgf48u0u4BLYZN2o6AtqeicsUxCFezZwin8eRLDX92qC
Nea/0gCMLmHIbmmhdkTnyoHjUCzWlD0kMEc80bZYbPd2IyxPWbSx8kz+Vh6NkCoO
HAvNQii0f+Yq8OJzzWKsIt83+FqDj9aMjtXRy2p9UE/f4faVsyMkXhv41a/atjFz
Dr6EiztYeapSB/vJD6tP3RUK4xNpaojSOtCoDzd/p1qdxJDCaiBMB6F7cOQWTIqE
Bc3oeh0gCq0O9UTw3vH+ccu2pJoK9ytXUkMU80OhK+aPcCKb7KiwHVuwM0o/o0Q8
qPRo+NS1f9hv4LSV/v78NI7+rLOtF+6bUpQWU5SHEyltBMnQjrVSSycBWC+dspAo
o4eXEZiPXqTv7FKE17kZ7yiNCH673TfrhNNCM7/mZ1QVl/L0b7Byd6JdpSLiWX+1
OnYJuFJWl/EmvVU0pCqCO0fA+LLXAnxGS6npYU4gD+KbEdP+vJK+MNxscin6dll7
Xf6YfKroYQWG+L1TcQgwEqWdnL0fWC21IDR0ij964woMeHYtYXsYoxF+2JnxwJD7
YW86L2qFeJBDT2vXhutDCKMGG24k5tg7MQ2692MNXR/49FIwCKR12ljLYMFtZKQG
An5gmWYkmlxelSCNTOR7UT7tAm3QlLlUv2Rif24FpF3ZfjAS0qEu7n0wQU74E7NJ
QBm6v/AzE99roI8fdIrqczlMTKC1YBVo7TPmTvyCe8gPIyBgqqjP4WpDO8vovMVd
QJcgb39QyOTk8Gp2n6MDtPw76196oObDEQJC0J42NGepkd69+/bbwFCy6km5KD69
Q3ueanxrEXclTc+zluwjbrIseXTEQ3/u6vSMFv4Uoml6ZZh2/BKbuaDa/SsAHk/B
7kXRM2S2zpHQDusMHmjGZF6xdkhlumxUjwgN83EbQPBJnQu3v0h9OO8TiLm0Jke+
O/g9lhV1k6uf4i0hWDzZzHL24emq9CaFKJ77HYbQihtFsQWIRb/503LDEEcegRUv
VPB9b2PGmpkJSJ3qG0pBQvCD1zAV0TKyDOYqMu0wBNnMxUTyWBembNWFZ6Y31i+O
rThiljZXYKrqilaGtHols0HJeJ42MS9uPI+K7uZ+t43nUputLd39ot1aaAoIPyAC
EEaZGabvHe7VIgQCR0tVFHHwPpvcXg43wYXLNjp6naU3F3H8iCCjDEQwx4TYyy7p
W0p64J5ZVK8T8b6bNdYqvzr+nMXBcGvt7s8/XaMU85iZOi7petDk0SAlHwvLeejJ
21J0XNYfFtuGT18Sr7WXzsoQniUVUvZUzJ2F16zJFIxJVeNxuiHtNVJ9/wZjtWcW
5Uj+kfmfwh70NXPCIMQitZQPWc1ybEZHXp6p9eumvX1GHWAPp/sBWznphgxB6KBM
sbBT0IU09E6ePSMA+muiSAyqiaD+54+j8TYIrr+TD0vtB2ASVWFTpQum9qrGYNUv
ap87sELiTGcovNOv/0MBY5w8LC9eg/yRooNnUUMnGcmqYQfTJUdB36lGhbOyIjz/
6tezHubgC58ioRBHCuRpVri3NQQTzUraTEZpRKMBSekAxnHc7xo5kKyDK5Uu0whG
aFbyI3Qpcm5rgyBeKg0F+SbMkGkWKuaZojVSrdarJ1tg93ytGGzXBsWZ3V1LWawa
vGOb0SzuaT3HyBdO+066SD4/l0Bt2ZTKX9MizOR6v2hQRSnZm5+xKiYgkFlefpOO
cTnvLLPJtAo4Imco3dxnIfrfwzn4W4KkPrtOJqLZOdzRjIVvkkoy3QaHmBzmji2v
Z/R+J9dSNdzahCIJJpOBnXHWcO35KKrqEiCbtFTQGYQ1qDdfhr9nurV5zWGBeDRw
pi4Bt6P2NayuMY9IeruyYfjdc3XpPor7GxtqVs5XW2jVXUJWVyd4BEAiskOdZZQV
GvF36UV6gjb4KjYiowbBQo+zMjlc1MU6lDUQQN2/8M6X2puXlpy2qr3gGSQc5X3n
0jZXi5D6FskZsNxvrk/pQMx3o3lq5MnQeGlLK1O+9XCJsOa0SJdVh4KToaBUGZgY
gvBOkfS7qIEFBVGkRhyDyEqnQxJ63rGqoxD+TBBanJTUN6nSu6q00IKg0yDY0QUA
X4RyUh0iKTNdNqV01879m3vtfZI36mCdGqqLKAAo3JIQDc42roQ44bZ8FhTjRpSB
cB5Vid9Jidd1SDtXULwPU5SfwSWuGzcknlgS/gIiVYJdoBkZWgRt0xBVnYeLKjK/
9KNatbCA5V50pOz0Q/1iCkrjQADLKkihAq2WNOLin206LmsEuwV4vKqisPFV0QYQ
7MubTsTxFnQuA9ojAgHgNim9fBCXn9I8LYfJ8uAps+64FhLjjJyKDgZJ0RGntg1p
fokG2PZoFo9soEd3YlbKZQFUQDcXzgGD1b9rgtOglZnsuJ0LheBmK/Oy6q9f+fTF
PkZvR2YF+mizmj4eQkrgLjYg/Cg4x0RMeAe8D3EBu/NSMQlx5UmR6L51ED4BQfPE
FaAsfdaVEjVCWBGktfRYrSvuig4DDSxPETQfsoGYTiVx6hQ6ij1waYxplcJIymJ7
kr2cvKltOWblzmJMKtQUBzEc5TbZ4LWqv6TFq+6dsf3/xpGTQ6QMBY+MhbaN2gGI
53wJjbq2GZDsyDu13tt8+uGBuS0rLnr7FzI39WrzEI9gADUJAt7bPYYUNF4SvlmG
UAW+LM/PM1eSgROf3VZLFn0VBbTP21gu6GFS6rH1irKzi8UKd2JU4P+KymRbYN/b
ZAV/rtPBxnQ2FOHSRDhNHtThZyeS68dKjzW1nAxFDBGQt1EnIYfKFm8l8+L8MKT/
hmCvBFL9m1M9j3DT44w8/DwzRARHFWh6xGvRi4IC5WJa/x3TnltlHuwv4L1Z6ZDo
KgYZIEAGaps2IpBsS9blo12hmtSQSUpFWx7Veh15CMLKJReptJ2xAuuJZXJV+3Kx
wk7XQ5JyjTY0ws4JzkuMN2vPxAEVU7Dsz1hYY49d9A6DXmzU+mU7WI04p3hwKT0V
aS8zOGEna2MswEpT4p/d0hvvvj1rt1/NfYxmLPydSqTn0B4b5rB/IfC0O+YsOV2r
45uwrl/PKqrl0tHwlHNRMR7qne0QDzkSim/IzsnUts6GrjJNvjpMNgfphR8GfkvJ
7QNSiMBM5TtXmnw50d01F5o0AwJGS8TMX3xRbwKVSLo40gCE8JL2qoGeBVgXCBLQ
n2BJEIP0WAxsSzvh1I/64fWzAQZ34UHvERnale7+UNZKPOeiyCofDsuMP/aw5/dx
v/hCHOne5Ntr9mnb3qDaDUSTZtLrmbiRwoKFSxgbWF9Wy/ffVxORaL8yOhEfMbdV
rZHEsOt8BMizCgFj/cCaB2YcUexYvqw5f4/fwDrkacMIqrEdV0ti3RjwR1vCmtFV
LRlOCpbYIL7WgHwgcOFr/fmUfFYsNIc/K+QPWLOQ/ysid519bHY9zaGD2JSkUU8N
ssn9xNaPDj+lXlTFCYwlcV0lQcNINXSAhegOOl2P0jilxZm/iTFKu/juCn3+BUiT
1epzIXyXRLzsDrUlqUpoEyfV0wCbvh9yKkYYgxuwi2SsfyBUNJgJEHfj+Ed6BRdV
14w83mGSXvT8zPFfkeulHJeVWINI1tqotI59OZbm8ermv2CRHNATuyoLgdehRuXh
n6+XTd0yUaX3REsQu/FkHstdzqpn5o8flCp9qjCjQAf7C0AWDclUIq+GQK3gGY7u
UuCQJKpr0qMB9qIud6xf3/EzqM8/CuQ02+tMTUt5JJBy63v5gkJQUEjYhDI9H+jW
udSGDPPb0kDZA9qj7aK9xaHi7enZuY5stjXvy3uy6+oxj5jwh9UVa6M9LLbDw0qw
tKQaGDiHxYmcTFruX9O0ns3AzCQeSdP4Onm7cBLcuHvHkGUvaeFoyDrwPKs4ae5Z
p/rFkdpy4gKxHm0WqdTcONb2s2mPbfh5ENPxJ8ZemVVpAU3XtYx4F7dzmjcEuW/z
fSeSen90XW8W9yaRpGWpHkbUxbziYUe6x96rf8LSc7LivOgB+NUbNpUOLEr4qhXi
G4uJ0AHdKzERYHoBDiZmRdX3DLSgHzGoHNeN+CcgTAxT8rL0c4erGEaxdlQxPFuB
tKdkasVYgO3CnlXi0I7df9Ivegvx63rq/IY8xD9j3s8y6ioBo8bcr2LKf2XsJVDy
6MZemU7sBjuJpo8CITtYzie3OWF4icBVjC3z8ajA1H5N28R8uRcsA/BvGW9flYci
GawvsR6SbPCMtLPNfQle8t+7tIekW/jVbMAB0csiqUBRVolKy7Gcu0Bx0vmvgJd1
IrJqlKAQi6mriKQfMy4g7AQj+oIezmMzXOVoZCBvlPpw3HSBZ2raub/+F+u7VeD4
0uc+ggMXFER8ziFwBRZbO/KDN5eHmVZ8XlqW1THzuBJ3RjfrB6gx8gQ/ARGZ+5MY
E3jIwSGeLyG5PzmuqPW0owVT8u6td0nEKjM8/2Zpa21PYKInDLFhDc2y6sIh0jtH
3mwPE32H9MQe3Vdd7I2oPd7dH6M+ORB83ERcvcZPePDiYxEgkHs3pySCLu4LqECY
vk27oYJSBBCS1V5t4ruIIez4NthBDYbbnLzO+tYyFBChLWGDpczdfETTvzzrLWFj
BBx4jfNLYv2oWlbtAlRJ6FMeYqPJaSyDXd3/MBgiBPly/W7pXl9oPHBSK0NSAEhb
EbgsaQp6SjAie1vbLnAdy+SmkuYLkatOi+4c6P1nIShssVHy464E31OsaeCoqOMF
OsQ/Qsnel+QcWybz86wMIAr592ihP8CCYceQ8zEIYpWzLzwgyzCoahidRKbEhvWp
sYfbahi842+5K4km2voGYNVpsEGejWrCKEPV+lWhZjxpq+Kw8f8f+8UBYJC+0F0W
4FhIvHrDS5qFsh99RC/IvCAJt5DOhFT5aAhCox1akjAWC8Zpt4BK3iNlGGqL0FFQ
0KI6DYAJbFyDNAo9VxJCFGqfP3xp05kD2Kkxe9rNgm4pF9QCl34gtHBq9sRa6dXl
HJR3vXPZnc4Em8HBpkp6cmBn6r8LUHK09cMfJUL+uUhnRTli+SRtBrJWSvNvr+vp
JupJiU2rqAqLKwPz1K3B4XMlkUeVyq05WcybEtyudGjvkJA9+UbEla1ix3jGE/Dl
6jJc3WgOP2k/TlWgM249x5rjoAKSdV9gfA9m0uEbFY5QBIA3GSxtQaJkQdgV8DCM
NqkH2ftEIkWWfE7ttq8mGfKYjGbD86V+vPv968p6nUB3O+mVDd+6f6alvTl9xU2G
AHA5Wxd07QJx8V3oFAtcftHYK9InwhZSKpUrxqbX7RQblCAT5aE7RYAno2CNqKHT
Xbynq7W9ZaFpN64W2Epi9kh0NmuiWqdgsqEtLer09fhthu8rT6zlcnLwArUd1TBj
Q4Om+MOpp6KY5z6sHo5sPyo+aTQLnycM4gKBrvJVWm5u/Dz8qYBvAIcB5qQyXmeS
lRY8L8TyLFK8h5y8Ad8UeCJnCSpnIh3dFSCIGqDKPW+jRe5iK9FMmnBjSvhYNJj5
5rTIgaNj3Rg4gXfAopjChhUwEzOyqylujcEGoiCx45jJb2NQsWhZjL9mHcyrK/Yf
EqzGhjJ8xK/WZ9T6cqvZjxgh4NWz/XFRGftNrTh0na9/dEU1LzHfLSLnDlRnf+oy
mVGAUQLA79S/Xepv3PDPes854FkClHeZqrhoXQ/ntviAnJHM4iZph3uZVsC2J9bu
3wob+sHJ/+LsL2xhgNII2Vg9oJg+J5Ri5chrMzMEv97iklSHVfqW1mTTB/J5G9mU
0/wa8ulMCNHEMppFnE3JLnIpt7CPtBiMEOks2ZBvCYAgquSb5f+7oMS2GMhjh4ep
nYzz6Tkg8WPT1Lsrrlma6VMiclgcbHZrH1IZMvOKE8KdozwrUBw4aPcUKee45ovf
TTXl7yID8hR1enBRHX6b7H0GUqUSW1YrnZ8ucmIsy1loQdS5GKuq+6zkCikQW1Yz
6nlYAmecCRRjGrGgVUEn2BwLNo9CJ+t3FBrVfrr+H1FCAaSvk4OlPatNyGLTAOEk
SOhbFolVZzKeWX/AgF8vsOX2znt2uOw2ONWDHCVlMtdb4GVL31itVcmUDRHl9+QF
4dQNBNjUWzSswF166IWGEJzEfLpmC2MekFb7NQmCd2+lhtrrYCMGkgZCtC78vtIx
VDXAfxBsxWnM6qa2t3p55DcH/h6kG88b6BPk4yrQRO8bML0h8G4NxtaBG3GIbt3X
6Tcf8UGmfaT8rXZoyT1w1aphh9el6A9cgpZOaj0xm2ed9aJJ52dR5DN+lYdg1n9r
V2jCFGU5TV8mteFVfYwOMjQFYqt2HjqMo6gfFn82ziso9lqo1lJaebKfEtnzvm/z
3tf2N/DPsdtTHO5HblCCRLZR9aDH++oGLqRYExtuiBdGFwoAjYcwapN17OLbMriH
MbCERrkdjW3W2BVySAy1y0hjFichAtJi7PKHyXgS4X7UPqfFVOWzIKQ6UJ08ge5I
RNXrPMINbbznH34VOz0fRQTSdtXgV105IQ6/FW44xj5E9IqT8MdEdw1L7iI7s088
F2V5QIu0iJST3YDuYhJ4XI7+W2CaF6Pr1zjOELTYkv+u+rJ21geAzG46sahc79Gd
iffZMxwLGZpjz5QFlmLnArD2dgZeg1lOCdvcIE25FMHeMG4aH46/SODpyPFEUx4W
WVNqRNCT3Y0ssilBb/sICi0qRdEd3Jyg3qzr3WA8ImIyyoxABpi7CTGwtVdj2O4w
3q+eaEKV9p1ONtDPp+W9WTFmv99C2/I/TUAMtNOStMOl+olM5/S9XHDw5jKgaWPU
sG68BnHbuZ88d8pQftwxPGHY0y5PjGrpB/ug9EH16xEeRoEYOKtlBjavJXw5zIXb
Mg+B1+Wg2rl5n9gW1wS1UItAkY4BqZ6EkyC2/zrgyjGerPD/g/e9pK+4iK1RtsSZ
xCbQDZZNPS4jGt5f8hWq9aUOR3m7DF8GL1VWkcEWeBYiEvGSh+UiEFuf7fjiK4XM
eMkfSzxuxZXfgjZDTfyrLg8VQ3r4q1BN/iYQWVotxhsb2IO/6XwjPlkssRtH5DA+
+BYtyaWnhfDUbDJAInOfoLdlrsX0fasaQXgBz9DOevZ+Du0FfFj/HVoJDzA5rGYC
ybCFlsDUw4vULdcCxta4XC2eYHsrImtXl3YyJ+rkAirwocF3c0GIQaKvZ+DVG49M
hnyo8wBIaXVWQYWQ/FE6MTOneDz/VuE4fAOZY8pgR9i2Cwrb9mlX6cqRTJTaCC8N
F3234kn+ggEVgKPQEroj6GGSNv1JSy1EUTKutbQOjlCJb6mP1xFoLUsMgROBHyog
kojAMXK4Eoa9k8UCHfvASWKvBb/bRmoaZKnNYZY/M2HXst3C3f1fJZ81Gt9KSZZS
xrdhSlCBcWcgAerBtjYZMZQ1fCIVxZQPCfuapDZoxH1sV4Wy+yiobbfPXo8Wrx9G
5Y8jVc05LzwrYysKF+KF+GvtDJ0hcvCOWQ9Qj2iYxRtCmt9Nsuyd/Lt6g/jRGnb6
WzwyYmtL/F+swsvMQ5yifmBBfqqJ9WrUSCgto2m5b4p3jFpjUMm4MdiFLT3hKXB3
0TnVJdk5MGOepBE0b5xCvljoKMYQcyU6+y/sglBCyqxpyaAB1iovn3R76U1GbKbV
MRD2v/JSrkBdhJpsm1B6bNQ0FXjzrgxxltTp5Bb8Du1bFkYanJvqsAZCBNmLjRHl
7TbVr+MU6vWFxl7D9si8NblFwkKRp+VC+kk2r4PTQvNb08Q8aqwnE4vdFkAyfSDb
tB8yVgQ8NS5oBcBdbjsNPRXhtiKPG8jLUv9UYF+++2k0Pv02M2y8MS4TOnL1jpF8
rU2L41uB2Y5OgnGFXd0z6NUotgFTAke7e6QFzN+BPWNJXQShs7DcQBjZs4aqcaHv
M05aXsFrjap45VY0cCKRCtXYnInY1maktqta6nZRKeL5x90ez91adzFg0tW5NAK+
xmAVQbeeGT2ULSa5a1kbvFOoP/PXsUS364oVD7tje2dy5R/LtJXFlO2dWBpyLxTs
J0zwsNMNc2ZmXKcnw/xni9c7YhG7SEBdGbiDBZZ/uLCpjAeb2FKTOtRw4xZXxciv
0Jlk4nNhz/sCUoosBDBIdPFcqeR/MyLYyBcM1vnBGyVf0jYVKmXCM8KR4uI2+tqG
OaSjQEIc3a2PU/ybuya4H7Ftpkyj0CYvLf+XGpYKEt0sBjOvEtLoXgRof7i5tBCw
ImbPYLjtnMHj4Df23GEUs7qG9duzpC3aBdTF4J9L5xClAhXcDZ6HpxnlXCCP8uKV
niLGrxbeleA6hhMQIBiIN0sfit9vssoFB7ikPA5QIntn9rkAVs+iWcUWsr3DTFOE
go9wCpslUyKOfTAOzVYkigqYEnSUXtUngn+8s1zMXFhuGRBclez36Jyaraollil2
pX5A7/b+UhpXZX5MoIjdOwH2kS5txAwjcjTJahcqpCJ4QRSDRsW2YW7wcvVtHSUM
A8KLvL2GCJHbDfSqstVVQllG2WeQC4lvef4H2o+BDDW45Gp4bC/4LluFOggIEaW5
UpLgnHENrCxjkoPKjLltcyO1B5be+BduJEWnqlEFsZOcOCWTVcO3ut9qedCpFZzR
uc+6TAnrqDGvvjHRia8N6K2n8TG2+15eBUI5/jv25es7aot9M6AAKVYC8xK1r6hK
gntvMC2+MsMTQ/XmTzFl6K0JrKTrZA6/H7BgAZj0ghr338ED9CKiJ0cX/fxaPfpD
dIVVOuqXiJ8BK/uztNXfwvi+DEvV9o1gEOP0aBUB3iqdVbk9hhPkXrQHDOa0/ok9
JVvDOFhoUc6DeP/tk39ljq3aTGteCLCit2a3r9HqsfTqtL9vOIUrGkdCeC5WQdsS
PJRdBTl+PbUegIHh4tNl+r6pYUBpcJpv9d/lm+8iVWcIYV+IU1ERhByUe+vOTN8N
GgWi36zry9QNTWX36raAvB9lRcU9lFanGZ7nxRtmy01+UaXrRp1KAaAqBmxFmOSO
kQs40yO1kdIjx5fJhp8Tp9fX/B9ICqepEzdMepExdWIkfuVZnCCmyx1KeVGqLiBO
Wr6xLa3wCoC762mYoreOCXaYhST7kHTUk3BgJt+PyrxldI7WTct+If3Y/+31R+mO
kln9Of9xlNisuw/7FVczad/gZ42VgI+PChRS3AO7JAgras/c7vS9YKzOCjvIVKAw
rOp1alVP/E/ASCzqHswjlJVvb8zCNNKFEKkeGaN3ZJhEevQ9wx14R4isPRI3cX4b
oODOwcoRf58Yx/VfuaCRY9jKTAGXNfVZgcw5cLzd7LMaP5qugJYZPGZqiCLE0bQA
LtuD4gPvqqNEJwyrNw1kMOMew5gU7wr3+Za6vH2WjlQILucnOMxeqgWGykZYAdkF
lDq938Fj3Xztmon6q5qC1d3P1DSpsRQfoOzvewZhB0ajVeH0qPMx1A/5LYZSiSa3
GjR5fWl4+VE7QmSbgCvgXstVPZlH1YGreZm6gIUujsRLr1A2WewWS7vhcLxpJfvG
50JsfR01Er/hYMI8umQ74EQnLFCwFa0+ukaUt6yCuHhWh5/TEhPyZ1diaBYs55jx
je25GsctjMPlwfhFD+ngG0s/0gmi6pG6jLJQ7HdOZEAMMz+TQPTmG2jjuWV7fqTk
aM9nfskFmkF77aGv+NiJIQ7k+QeHICWn2Fo5FQ7wzQ87Hp27QbU6y1z462GlUs/i
Ma5Lf7idz3v5eADavYPwvRfgoEzYOXA+OkH4SNDblDQV5qkCSkiripoCuChmdxLE
vZM4vN0uzlbvredKx7wF1ijMWDzS784v1oFuZOanjsC3mw/S7aDe7QJ3VduvEbvH
Ag5yt3pUgH+q3SDGCWqbDVhQDiT8PXgiBNFf/uK5gIbEl1BmWC+xvcy72Tl4wgF4
yG3ZQ6/WyeAmCgzBB9Xl5UU6ICTApDGUJuf85aL8SfXJzu0sjKZN5ZBf4UGI4eAm
hGDfF9mKlvPVbbkNezxM1nt+soBamdWXgNKJWrTYEs1BvR7nsbnMyluvQFnX77V+
YuZX7ZmPHzQ0EVSdQxoXmc2Al1ojOodRIoxpDOEFT+gGS5NDaBgZVL5uA1QR/q1z
EEdex5yfJvjeuPS8DoB0CydfUPzINBHALKKOkY3MjKhgKhFlKFKXawTTcxNNqi77
kU9TrHvSRvLJv8NVmXNQy3bGy0PGXkbm/jusgVS2p+mJvHCTrfULVHFIh59rtV4H
feYUxi0DcpFDhFnThAgm7TYi7miyADACyuuhjKWtcd6T2Moi2DoDMk7P6E/A4D8w
LHpoHz9VHYxARWujFNXyO1ovingzwZvUEnB4/QhiiSrO+ZuureMXZKMbln44RGz6
etUhJ+pToO9mqCxdYAtVvYNlp+E0V6enCgBVFw66QXVCCuOPp/lpzl+UDMF0H0qz
HSJny7ShUck5JGdqiVvzKULe24/78ns/8b5OIWTUanOfw3zl1D3SUKwt+CwsO5Jg
MibZxyv7JyyrAns5HBIuH/qPm+te15louVFUgk23C62kd94FL1kZSFRV1AIrJFGH
6osn554rlnkWEu8jsfkrLSyR6G1ElrqId3RJNdu6B4mi+LQez9c154yns0PtxU87
MJneSdyj/6zaWtLu29L3WymrYVSPmpn++y6VajdcrK/QBWad+jb3CRZDOsjHFw5C
+f7p8fYh/x6G0dOZvdL2SWfcFIX+EuPvxaeNoq8FzT3G2dWp/l4klYXg472BgH9F
xnmcqNKtb9cdJGBQD7Gd75+WZvsO4vGG+CvfO6dP2DqudzWxPt2oYL8qEyfoamND
m/bkOB+hqqeHpjy0jonBSM6/aOt/ayuuU+DAe4h3KtIPBlWhSrJ13auQ7TfkQ1D2
M1dRImVE+TIdXyNa9jabYgHRwb7ar2YLjhNfwU6vI+qdoNSpoPIgMfWFFDNJpZ4K
rcifzGR8rA+52Vbg2RL4Tu48lg/ZrQtT0QrIO1wP5g0GYDhMzOWSY2sU7W1uGgoV
l6ar9itWC+29v/grdwPsxhnMoWE8kCBKIpCyyC2u6Zd9jgspFG5H1tbyp1qLm+3Q
/SDMWbZYGnToS8pcpt1jW1UZEPB+8JqXAn7Z4/MKOnwt8o0gLmODY/XkducO6gOC
s1cBWibYDivDQaLhs2Hhf461cUFmLlhWzI+1z/7pWG5UNv8vmus8DopZ73Ethtae
ts0MHJUUBsB4tAAAqaHSVcE7Xmt6RdRC5qjT7k+9TMCMV306pc4BtQW0u5J94fho
wbbVy3P+M5ogq6/Z8hNqu/E1BVaToeGs14iu+iQq1ybtyTnqjg3NFCJKYEHMZr5h
JgnTfLAIRUkXr6/L9Hwg25dNnAVORen9CBS1rA6MLdVb/aG8ugY08/bovgNN0IhK
GoNbIZhA8kZOuD9JwmtUyCZq/P0laBniZzxOHjYzcVWSMXJVl8t47KzquhF65Cr7
fQluSoOMyKVx0S9oq5AF+0FtXMOrFsUN6vYLcpXzmro9iorpcVebnCyJNe333CVb
7TN+UcSyRzvFWfgwCAxuDuwIoW2oJwYN+9YuKKfzTEpwjBHusNLbxCkOiUmcres3
Xl5ZTUP1iTx7gGz5MVQCTgg4Ldn2R5cpB+nSADsbt9sJ1hG4ICXfBFFT7Hqw67+Y
9iUJzqH2M+jJrubLDzsfKYVMZGolRV76TiISskT9KXiia7uvRGPAl6x1wP0VjgTI
gEWb3MZkoro+OAD8ANXAMzhshbQRUyu63uaY8L0D2J3ma1x+rL+UFXN1C02pJZQV
Wx7w5eUOirtxKt2OxN1so+hBj7Br+iy16TpbdK5XOifQ2nc1HPp8ckgf68ZK0YJ9
yqKVnEFodHK8Icsb5trbepMx2QLqhaUOqrE2wJYLaqRv49/qFQ5aRqabkY9IVA7c
8V6n5nFx/BnzkX/TFX2ptR8vmN6QI0aMK+Me3iTiZBqZoBavdeulYPApGKopzAau
eh4MM0nw7nD0wWLiiq63U2SIo4J+Eqhb9b804Gj5wmBRY2uxAGaqF8Ta10h+skQg
TUkghJ7Ls+fGpe03DPbW/A9vPHs9j4NZoEajCgJWrMNYJdW29j1K3T8kdUHdA3JQ
SHjo6uLqzXK8HTM/bJdopz+J48PjGv94jHZULe+wURAhuebeaCta7vO4d8cA0n+5
P6Gv33sKU9MNTA+7A1AVLuPaMukQpMNKU+/6P627Hi61HR2NTYxDzNXC2sSuIao0
+ayFq8FstgAAEEkUhzVok/qHACqkcfC4pIQ2BTsAqqg03L7gCRiH91gGONFZc7Rh
lOpkgcZYfdfvbxEmFInDmcA6iql/F/AX2D91UIvYMidPhn9zq4H3DZuon5r/BJlf
V4ttImQc6WzavqfKJ2GLz+XcUv7X/VVi/sa/5l7xO9QHCTpbxnjAFwF0UGsdxW2F
t2pKpN2EoF4ApomrsLifD5UbH6ohwLgoYzgCqBC7pFR84f1+iZoPFkslOX9dqo3Y
oY4R/38p4c4Vp8mVBAbqBWwL4mAEn5jfVMaYGq7ix3h7NIhxu6np3XR/P03fBJMh
++fWgXLbI+mCQE7ydAuYkNXY2JqRjGVf8v3MyBo7zKX8zzXOcbhsdvE+l4/VbIk8
o7q0oXbuFYXBJJTVcKtSJuSOruh8OSk7+zdJgBmRSqyLMgtTTZfcv9yHwZdBSQ0B
xjEC+qg47bUBmg9lfnGG6ibJhpUE0xEuMD6MIPCNxHJ/s4snyJNjejvSTBZc1Ibq
svUwH/RoJNN96C3SY/KR1Nr0Sdey9bEb3zhoDfd/JU5Hr3iqspsA9QJZPUTHnwKl
arSELXpYiW8Ao6RwLOov4qu4sJxez0L0Srf17NW8xjuLkPVt2MfXx0k4Q6eFuV1R
jTUFlex8U60+J3SIK+TeaLfZO6MAItlbdrty1QKZ2LT21NyjB9VEYZosRUddIVE2
GdA3OGb7BmIYAApbk33VIuMb6lMevc8LXs1Hw+gJbUsKdQykOWU7M/DQgUDdZVnc
M4qtvdDIvCnvyRZaaZ9whCFV86PUObjLlQWul90NY8iRY1ZsQ32/0O+50Syd+eEW
LA/dFqyERg7rcGgJ0oMJEW3pzQe+QPycz0WvQib53LxMh1auy6SIEGnkn1xQFfWz
4ye+b6gxVb9FWhXcqMav4y8qy4DlZe0jcK5kfv0HiQ7Wp9PB4hGHpE5JWQ90v+sx
ds7IcODjvQibrSS1mXHHsnSN1tiuR1y+jahP00mZpGa/RqxBjjQxcPmS+UKPCTvF
PbHwv2XROUfalx8uVY07/segmJnoOFbUVpfwbD1DdEfqHwuymhOw+DBButMV2BdF
qcbwxb+zcNKHE/C+H2uifOJst3N13+YvTDII+ZejfSLqUCyIs9yoHbig5ccIgspj
bfn8CybTuQAAXPV0dDWrScnHKv/lCKv+4UX5niRFOmGYu22TJW/VUlmcGthfIN+K
wjeOmqRpU0IoscWZE72ovRiIQYewHi4j9XDToo2u/mNFwZPlp633HCEOmQ4doRBw
VbaJ0FmJLIYytyM64oSwkDP8cRKOSKln9KsCUhFp1KBPpGuBWIobxdToAM1Fz+BT
cv2zY+NNegS7pi7Bd24s1PbTCNGjbO/RrmyNAB6Uu1p+ebmMwjJp70wG57yxSW1S
yPPdY/9uK9/hjNvnFBSgd5eD7sDWpgG3dOH5T9pxjMtf+i/NhXKyRnJMl4f50vES
0u1IKEbwd1XDZ+zimAIxdkwFp6s1SGV3himSWGIO9CqjpEmk3v7+YvW9KeymAU4t
1LTqhn8J0x9jpHWb6erGoO5zNw/F53R6DiiaePhfkjw+6pc2WHZy3dmtSQDoMKxQ
+vPgo/JB3sxTD2Nt94ITWLS04PyrR3gA8BMOnPDhTSyDVZDvMjKImDit2WBoWq9E
1fhgFUrMwdc7sZCF0v8+EfOHqvTtymLrYKrt8+/g+kHyFifjnuSpZ5raL9Gho9LZ
009UeUe5xWvoYGvSeAo8Rh1jWS8kd2L/KVCRgpl/YRP5L9EIsupIhnyCTXulDoog
FeyK8iNGcL81tsYUixIg2JnrWatLZfwB5LTSVuG1XJeibzcJ6q9WlpADX3hybk4G
4N6DbMackR6hEpdfFCUQ9+tRdWofhLQLqegtwR+t56tLov67D/b5QzsphVL4Tava
sSbJwU0d+eWgmYVSRqwJjq09eU5/b+bGnON4qY54iHnlesWbNYkzYG32ZxM+b/Fu
B0esvmRLHHzlNPpDI6GH8zhMZpGHFdWlvkO1XN4Zw7DkoLiISmJF/JKzoCD1IMt1
i4TblKaHICIh1mvOlSN1Djt6sjICgortXOLm0J+Wz/dj6l8nvUiz8nKt/HS4MAaz
+NMkuNIBflbFNgjPoGkOMazZf4X+m/Ecy7KEd51EmmNC6a5IDsR6i/s9H2LFEBk1
e6+ucOqAYV8K9bZOrQ2EYTt4hKNC6VJrab56Q2GjdVXPkJsdpOIx3+oR4RPo57sh
liBCyTsYT7oKn4N96RF+rbaMvQ8Eg4KE+hvhiInpsykAEPSxJw/1cwzO6F5bNBYN
00yxpnFOQjyf04k15TXB68AoRqJyVt0sMKUzhG+zS3gequToOU1A1JoCFGgbCzHl
CcoQ4YQILC28XYgsRB5rxEnN+nft/r7BO4x6xosz2jURzqiCw9IpapbGACumq5D1
uYY2+4oedJOCCUe3uWnKh+kdxc6aHbuadE4c0Jr820QoHPJa5y6/9Knwthg+vIX9
t9wpGH/wkyqtsHNk97ozpVS4XnXJr1o055ff1J9hioY0i0JdFyeAbCdSuYL+CpwR
m50JAtu0gooaUhMbU1w0FCwL59n33uA9gWGDJnbZk+IqsRim6sQEdOqO5WDwwmas
Bw9im/JRXBgdA/clBJd5q6reBSph+Sk/yF22/jt18SqlB8C8nPm0flU1/OgEPTwy
TdmYnOJOUFAvAucgLzJmIY1e2qiqepjL/+SeEhzsZRjLcep/GD2r5qEteksibyQm
2e9PmRkmKz+d8XxuSifL3vkYUx1Cq2INx7KBmlcAPYjRbcvZ2LGAhn/BZTrSjebk
egIUnMCrYVGyeQPm33RrKvuteYYnRE1l9PJ5dg/4x7nuWJyU2Uu5LJY58mgtLqFk
EBgT0VhZV4ko7gFPFWM0llhxe1venxD/qXeHNWVRddKhdRNcRWgRvsZ9rJqLxyne
8jYcKxGHAaQCZP2S2LadzT4ztHh8hK9nBFBvYQHZ84HMaNtValHNQTN+A42XX0Cv
XectKlG9/MFCLqxR21/CHX9q9rwSO7gPKsQC1JQ+1DHiV488Y9MRuJtCyYPYNuUf
EyqZTsNMtJtWgRihT2tuATkEBULV3UT6xLZ6ee5PS+4X0VSxlq4O3rcQh7hOaufh
H7bbJO3kXvL2bdY7JoFo0/VFg/l+lZYU5E+iGFT3yQKUXPDMfIH3IaQANZsyDf5Y
BaT9bOgSVRMAsrA78XD77/dm9zns2Li9aMELVc8HIJvyiI+nH2Sz8qoDJ+tqwXky
Zl3TvRLq9SOCHdBzpDDJfQHqpLZwY/fclERgPU1Llks7LPYj2nefpdZonGqC0x6h
HfQi6+wSIVi6z1f0WT7caGEGatXxfDPrFY9EKtD/4NoLPsDfSpbv1T/FdukNgWgp
LYOHvPh6braxhTy9SP5fd5n/4Ce9cg3dXPNKipO1gdycuSRiSTCsu4IPynHAXYqa
AaoRQdNxZ228cKo+2/m4Hp6fjooVMFhUStbBOVoWDGkGRmYgaq+r8ISBInX9/Y8o
L9OC9sg6I0Lhh+nbOCw4ziffDufnXb8RTdsgJWvTCssYx1YlTW36IDwzYZWXtEWv
jZG4Kjztl2IaGsjQ4+uwSiH3wu+kRYFcN8XqpSF0fVALFG7IDwNtn/HaAj2CvV3o
8eSzYeiMBollzqSXnMyjOOzsrq7DITYCn9NkXGPLFYBB8+OalhPMvzUSEAigLQAF
wyNcqaBk8WPfUWMmheyI62bmWNTIXkINZKRfikEYfdhikAEslPpkqZPfy/KDJmra
omyCa6YOe51pJHN//oPZWSP2TbhmpTSLQo5OM9lKTXOmjhd+sGkG+z9eUPgLqiu8
Fy07+2wEmg7yaqCLm1CvJTHi7dUsGvmRn3/4yPSTC+uVh1yUMXgIeVCjVmW/KtkI
3GfhwQHIVOMlDgNRH/CBZxOQe3V3VJYyi2G497MvVQhXXxww0ZVRAqg3zGgGA4jA
URYhc3vQR+YOSfpRqGHIhDraitu4UcZuy/POU5/1tbrf2vtsdV6AU0H3dAnxmxKJ
CDnse0Ih+3N+xe0rrRc8gRlKRf5TexR+Nr0dDkFIomwTqzv5MKvXuJK682v62Edk
+L/LublDfe/NzS8QERu2bXdNLjvb5Umb9U4FXOcqEb9HKA4jEmpfLmpc93jYl87N
ewiOcn8C1lBzD1uiUmBai2L7+ABp9EXZHBSrh6vJnZxRC8sTIRfYL+zjVo2L6Oc0
1qAwI73VXp/sflt6B5RbVRQmM7I36yK/en48icC0qXsbiYUbn7JxHBlEih0bVO7O
rx7tPx8WgkkNcJFyIxXa2w1Z5l8uTF/RI4YrKI7bQIFeVBL9JHr8Jmr40YHezcV9
6MBRhYEdnQrpJaDmuNJX9TEZmU+XfHxPcrH2P9A5K2R3YHRDN7F6Om/hkN3pSOuE
q8mibXzrzgqsXriaW/Gjl8yttt+u5eJcJFd4dmi7xiWRYRFhcsLhYAtV6h9n3H/C
3Uf5pjrMJgOlCSp79D8Uby5lPX+76QBQB8cGKTuEa7UnmL0mfPU10dZht6rPoSfD
mkKjpHDFh+Iz1mxXmyItahAHg4qvw583bgHOzl+1Wb9nB7Yljr735ula5Jeoylcd
6DPYCinfMx5tB3FJxQ8a5Nuv1O7nrD6VChhE68PLaLBtocdEVjGMnF1/4iEhZKm5
iLOIY/Z0jnBNpmIN+KIn1j9MSOv5NTk5Cw7g34B/JfzYSOiStNDRggI+hTZVk+nF
RSz9G1lnirZmrPc8FlW83JtxYUgLcsG3fhCBTYLtRvbVGUXa0avETYQX4yRdOynr
P1E1CkInVxJCshmnlXO/zyhQgrJcUUsgEyfoJMqqo8d819NYUCIAOQFfFoyXugBJ
whpu4shh9ebJecpAi1wCF4zss/TRv3C3TI/9mBlbqcISS15/yqIWrkTR9qr3rCIE
LLpJq8wN602AmPYLB7xJ864NSanwtfbRXNW2E9ZBN0tawHGtsLqswt0FMSo4OdLF
cqLbWe0MoGfZUgGE1H1+wasxYgYB0Qp7vBniFIzlDbKj2CqjQeV9+AvK5041Kfa1
WsBaf8Vrkzu+6LCWV5V5F9C0sQwEZRq1tMnErgnkNIop+jxf7Ma+R+eNUE0CpYu/
x4KM9avMWMemkaPW5D8zsNJEmyHt0LJa1tVjmlaQInCALDN8BtxlxhzQlWUPiMn2
LiRzz0Re9bQgMeqwfAUTTcKN9LtlmEzEMRf9T7tXWegiRniugYJa7LypPWpmo/pW
IciUx9nXThFElGpwUAFEWhLF32QF03mE+r8PhY5yTP+Eoy1Qin3SCTAxrviWoiKo
yLkc6vtdWF1cdHfiBy5qloh18v7KVDYjKxBzJWw/NJvKSIZGdl2pruZso6631SbU
YI1O0Dch0vi76IKRBraZAWOHWY6t6N6UhcNggflYY+ZNHIo4zbWSLGFwp4djjX04
mXKvJnH4dp1900a8yvqo/Mnr+Vk6PTJ0+N99Gxuq9IQw+D2MSOWULRQLRljOTAs8
wBLY0QWtsv9fVeuW0MneGDQh83+ZSTshArweO24wWTL+cr2/BRDpDGqhn0beAZs+
2vdpM04BncV4gBxqoKgRX2DJW7lSxEteTFhNoKC8ipgvc+5miJ/P7aBiSkOsbudB
uaV75xBnvOvAF7hfYNzQ6zVQjEJ1dbWI4KYIDACUqSbL4JxrEGdpawsuMSmWl5fo
5vJ0fvVdOrcB6EvZS3PBM/0luwgFVRwwJjCKf5Mw/iduL3DRrkvwXmp/1B8RDOP7
UnEbVbXI6xEBPYUyap6DZ+fFdm+2CpRwp05ecZmJFEiAw1CSbHj4WtNa867EXjTm
UQMbZGOLN0Y0MyiqNRZPzWmmmaWo3yMN2trOCaO/C7RtfIuYI2EhApYqV4xzEKOW
uD9qe+cQUNWKYurPNdvHymOjQGy9Vr6XeGFucjUCfrdcDjDQBSX7k6QXCmCtkHxZ
KewUb6ZFdo1Tgraz4aWuWx3w5CMBiTMRBKjJtlpe8kqD+DlK5PTCj3Im75fpWnYZ
wmxLL2bVUUqiGSujYc5Fitomn/yjb+UJFvcbS/7Zmde5bzbwXxsfzkNl+DzTc78N
jUBqD9TZXK3dAUnawGiRZsfHeJxI+chDhDVqRSUWwSctoAmNlFXcnjVIadvNZFxS
II4lPfyVNVpIbDOG+OE9JzxJMbMHO+ydGxmVexVMeWA+ssqswAC0MBznc0jetJQG
SPV5AAUHTwpxW/R3ColCx4BE2NRH7WJlKCLwk6YY6RkHxCIjdiQzo07ad+XLSfWU
FUOh/3oQ5t2UnRHWhqHGZvv39AAE70ZY+jl7M9YJGq4w4x14gHC5sD7h5MZ4+uRl
sYrmb1muggJnYOkHtw4na1+KAzwlVeDxldsqzuUnC8bI8tVj8ikbRzo+vV+5pIZe
JrAPWRhiQmr5H3nUzB9ROBBdJ1FS2zjMERhUSBmKdXx2cedL7FdlpOFVtwvdeLXj
ullXeXjieXWXP9di2DUe62ChaHyDcBDQ0S0ClhUkIgbffnUmTPQ2VgJM8gry/KAc
Vp5z1gExEDfh8NQfxePotgUp31C7dsY/UMqfSExSi+1XImyOpTV2SVS+WQwRj4TS
l4eafaGV0TAhte7lu8gnTLuv61Erbsl7HNTi/icP4u/QOZ9yH2ZMP4Vi/VUvGj6r
SVGaJLhBXilD/dq7X/xf+iQvmv4xGoElnnkYBdbZFoajrASoEtbBmChRL9jRJGsm
0dOcGK1OaNhTUqUyTDGjqi6ncdJ9sKf1+rJwWXSWHOi+j+YHy8QmnKWOi0+kfSTc
ZYxyRB/Zqi7rIJWQObEZ489jgJhUrDqj1GW4a0ArwZXAJ2Eo1Usx8Fnh4RYWAREE
3DO7Cbm80kR5xOOIdNbvXNcEWb+/05E59CXlB2XhpWU0tgsa8s9qETeAPtNmzNpY
bhZKGb7T5cPG3ebLJaJJ+njWrdv3Rna/ao2WfEnbFcRVKHwXMsK4M3MANyxhnU2M
BxbQBaQCITwnRsl7VImO6n2IQV22MgoUWp+Z0PXQgqzfd5s+lQSqk9/k1Bl0yJw8
NU+9+K96YvjrNo+uwLsNvTXg+AMdScYpr/C9Dp46t2Gz4XcYaTExuecyPqfmhqOG
VqB6PdHMh5YaBIIQEJnSNFx9/sA7/qF1gDHGDk7X2MApqc1ubWKmg8Nw/VNkEJAs
CzZyfX2W8HJPDtZlHDNQVfnrGGkQ2zf8eVgbtj+k1tk+bGj6KXQWD68E9iV5Eg0+
biIkBt05KBA6c0N+RvFT7MgpYsvdJ/qJnXko5W7VCQM/upisAfp4UIVo6uPRE03D
xDL45m0iyybePUd1fgYcBtZ+teAA2w00Bkkoc7Ws8DfxGgoyguyhRzEtvEnRPrIX
I2wzYRUYyM8r7lI/q+wpZMhIyybopQppgztKZf4P8clrmJzitk3TXRMJ5pAV7/LJ
KbUWVm0SMJpzlYicg6RpHdEDZLZjKce2ouGcatJd0nIkadFLLux7WNjtU2EaO6pg
prFo7xwXlDgerJs3SCncPpHxLntNfFwPAtC3TUO4Sl9Jxs7I8dDMvsUtOKOL3oRO
qVfLv7AIUiiX50OmW3f1/nxesvbLwsxkyW3BEjWY5my/IUV80n8BL5atZgte0HzJ
ecRSvkvH2yZdUFsK7uiDC3jKOzeyO+rT5hCrOLLd3c3APEvDNP9u3+RY+gXzmI0y
/y6ipmhgju+8uD8tKIMV2cHLfW+Psa3suxKMqiHQ7KSKKuMVrGsEzjNcfbmsKAXf
8+9pcYW+koFRU+x90CEU1wBeMU56yS9hx9t75l7i488dbaO8Z/Isw5Rvp3US3Mj0
NO0RtybwtxRgCnU9sgVfgzuYcKftpBooKW35ZZr1LjV/Jn40eRodLJtZ3wg2/I42
IwEQoTnWLKy7dMXhyvXnx3nP7OqmgdOaL0Qpr2TGjGqOs+rfYq6tprW+TBt3J55V
/1oaw521pZMOWH+ZBEVDwi9Y55Hkha8YlZACTAYF1UoWntW4k9IpFAhK5zdDfpXm
LGaJghWz7UQOoFJhHjXN9yyrhl0SsZ8zeT1kXquqb7fVr4yZv4ChanIQqIzExEO5
Fg4Kg4+Rx8hp63N/uaprUqcTaFImL/NOuANyr0+CXPEXvfiruwfBphfcj8pZgqeh
g+m1JNCeWSGtZMY2grTAniRbr9KfX4CX3S3aZjBeaahOFG55Us2rsvshT33d9Qzv
cwEj9rx+cxhY7a7Vj/iXZCvaedA2HBT3Hoc5bBSUWWmrwxywbwo7Yb0vGLDTILGj
a5GKgW1H+tJn+k21G251QEzLeN7uijN/ntH3SeQ7Mo9Bv9T/lJZ+u6mwRL65XGz6
jVbqme3x7vsIxhU8xKIQP5Eu7lmdwqVpKRoYRTGFkEMS3rDBvBA+R9PQoFU1/Qx4
DFPMmYAt947xYY3wb/92HzRvy211p3J6MXuRf197GS4hOFYqCDbdCjjHKuzDxPmB
7SKi1nqDwn1EjWKZnATEdP4zWPfjm2zUBeI2A0Ab7sCjPiWNdNAKHPnTX/48Gtp2
B7kPt3elG5haj29Hv+gQIS29VfCVOdboDPtBrjrn/tACoBIwIopoIK6pr3L7gX9a
vEtc35nRtCjC2RenFWPT5K29BxmiFNTeOZChs1B4j1x+irPXTZU9pn2LWOfISuq7
3icF+KQKkL4fLQTV6ghLvx9BxmVnO4JFD+0O+jYWPYNuHMOO2o9XlNfIKANPQ0S5
kAnr1yYhZIrf6rzp6yPDSYVinY1o+M/NzvEakvaOWT3Z0/A1prID4BYl3fDCA5HZ
veZQu/vV7D4YPrsN/DmmRejj/OMVC+PaxWyLV+DloTPza5KUiGI5hyDRXvdzNz7E
tPipx6L5SLSQudtXOSlK3mirAsBefzzrhojkf3XglfUDtSTcIcZicQWt9fAnljqS
4c3hb0cvptsAz12SvHnkG7nEAdD02mZfSztky+0lWb9zxAl5dBFYbL3igHeL+7Xg
V3m3PAgdyZ58zzsxwKTJQu5kS8xF3ZnaqqN88CYFIvCZ0wQRcA0+W0NnzyafJ1TR
TLIzi87Z7cAwmLLdaWkHx++HNYgeCOnIf49zKL6q4gHZQe6BzN9DLE42mw0qOGDE
RpKep9ahvz3cNvVJssS/K8Fsy7a2/OetqL14nAdD7Ef8oS/raXxOrIplhjCL421b
RoJ2G/QwYfHpVyGfE6BfBnqm8sudZ4ftIRl6iPpKrJbGEcx2usaYYXf5YiamqOHw
gPunyvQwjnSqz2EQq6ED+hBHA6U5/hq9kHG6miKtYJaLbHmV4MYdKSgzedzgI+K5
1gccJchbqPFqrxtChx0n2xE1BCvlGZPpwwzhrVXnM7xnO8eeLbPcMFUoO7eHpYzc
L2jcNAhEh4Vy0AOoER3k0Rl+P6XYnlP87+xehloJE6crvtv4jOWWgoSV1lOhSgf8
8ey/ndr+wl8K7aGVL7y0T/NO1E+8BvMiWOQ+nGoOIUY/8xYitxgagrqIxLN+ZNaA
v+hoz8yfa0o6t+0JIepRH5iWpSnkJiXFFarvOnggFIHTZFhroQdNz2z0ZOR1Czdt
Zhgf4xX/ojhHMEeU+BkmsdTsUpbpXu+VP2n5gSNT32Ce0JhzK+AqjkXUkLLaWL8H
lOdxeNjZkTZDxYPGQJakAjeCYxcPVWr68918/XxRh/0NB9DQYBQNiXd+OBViqc3e
sgR4GyxkIywPlU1aSESMqzDyVipjtG3qZhpqidoPkRS5n5j42NBnyhkcKw8pUy1a
4OBcnjp6sAtIOYIsHAtUZx/6Dnr8jKNYwbrMf1JJFVXhz0jHcrwgK9yXv7t73Syj
8E1CJVnWFayks+1UIhv/BFeWxprEc8COXwCtDq+KcqI7yUhdCtyLzBSFp0Z94lBR
tafyvVkAwY14O6CkfvnwGCs1JZ9pLNhiNgB+LxLxIZLQCuGu/iAWPrZ8wQmFi3SD
BdjZ3WrHJvepHuYPFP3xM+CnHic/2UquN5NQc4ZrMJfw80wv8+FuY0R2npt1pgtA
DYAw10ne+d91KyYyflonLGW1rRm1bph+bAKmzNBDwjuj1eKO7GuHZ8M6OZVRLkSo
Jpx/+omJzC5xcrBLmxfaUqeAaXJGy14IBfrQpVQWUqeJo+Si4j7BDyB4JIQI8RAF
vLpcojnJkhZCBEvcPgHpYg66qNetlP3jf/6uVwgsF/Sprx64ShX0+4N4IbpxW48o
v16YbaiHcrKZ93lzvHqAifXI3DSf2GhbOZPeHllQiCyvlJGR4uvBzkJpgtS12V7h
jG9K1QVHkEeg5rLiEvvbrybiqvdKEbb7x9dwoDKmgN0t11GeJWjMX9ADxWcLd8Ab
ZY9IAGyAc2bsNPyAqIizMva1SWuUUfcG6gNA9PmRx8adXzOE+xw5sDzbC98nu6aa
Zg3/MXq14mg1Hz36lrQZRVUHGlzAuHyXhrtQMKUcL0OsgQormtS35UBDXgoSebup
klMNCu7R601yHxgJKQwUq3zVACD5uqvRlRVu879Hk6Mn+PgVGflRstJftE5aHRTF
UnvuNtAvCICV1CN6Z2XxLs6FgXfjy9r49Y/kDo313lCXUdEGUvskWLy0jdzfuwmi
vXTzkgEQs4NxMGfSClZIDUX6OOUiJJ0ENonEktwfLvxDmoBGHoef6309WiGTcw85
qfL9/Wvhw9SyvJMGV0z/p3+890EaTVwyJ/pok+e0h2ppAGAjmO6gS9DKE0EYqmVI
mSORrQAHqnZvWtfw26GmyyoYt4qu1D0A8cdJUJB50l9jv1rHI9hwaj91JGMDIwOh
qByGjNYoQz6rVOAgqYHAoqN3lKwJDlJ5HRENfFXFsuA7s/H40c7u9HCIqkUpUYtC
KxixaUOJ838JRBIoLnM7M9OFy2H0221TqiBC/w20WcZ/TKVWIrr13d4fbikkat1z
9xHuXYu7D0ygQwIHhnQWmnQ2OsJtM+mf3MK7D/epxeN13hri/0HU7xHms3GWOmZe
FE28+1fQAmBLQEdORESK9/yM/kthC6qQcNGWZtSYqxT4onT+Pi+3AUHvcUHAkQ/6
p2K8F0zMFgDQ9DjF8E2OZoP6Zw9bYfRJrT6qoxLaPEH/yPXI06uWZtLyEmDPdkZG
TU8Ifakx5ohtZwP5aS2Ofes+QOcqW7RxWMD3u2EEG+NhkVGfKHFZJeN8yp3I3WK9
2mL3ke71y7IINDgTjOqTs+XiYuATee+q2NdYaNTG39j3LGoM5fZ9CaQUUSpigtHD
ISAkTQa1/jQXK5QizCIrMWkAcb4HOLX0JquQ3zIt85bPj2OGpOV8qpg2pepr/04B
vy0XLKV/Al7GoCGQwhXPhW2usZMIFfsRVhCOQoJCT++vabe6+joCjNwWCd77h3AK
EBPywFnzDRWfRrWHLUNVfZVFjSM8YjnqcY2oYDIkS8Yn+H4XZoObNo6Wbudh96ng
JvCBUFmh4OcbeFWyuHKGQfKOC6h4CFO3T7dUqe9Uu5uX0g2mUx+F52Hx6hrd6c0a
wvuWeq3PDmut5+ZCjZGbjxHeVn/v5eIjPJtx2ze8mvG4m6nu8X6LPRfvqULmJS81
Mx6YTv3YE96CjbGo/w4YWaJT3W4Q3T+bjbmjGMPPhxYeXUIqiCj960M6LwULKeO6
L59AnKOHUfsmSKL+LjJeajzaIWNnKuuzhWnyJOojymrzHt3lukVElhCCcHP43IFY
DIDwoP9i51VBTPukdgwkcmGpRSU6ynbOdVtJzrxGylzPyNxxvLIPO1dkUl4JawUZ
/dzHqFra8ULw4Pw5zL2iSyIbzTrezw3vSjkIdbjF3YnE5bkHmazqtwIOM50R6upY
ZTdCg7Dxtg5dijgNdVz9UAFxCV12FxXyWbSrHOiW3RFVqnNx++6Ws1B46MBTNdIw
XRDnCJhbQDForLuJSUhMzteLgXZOQ7cqzxmkHu88p9DoyOebv8m5OePWVPG3sgVK
Ogf53tUoyxgBHtBcUM+xOlxFjWjXsnbVLxuvaReScNPb90oOZ8Apzey4qfQcAm8V
E4h+6Gjn5QHoW3choDTp9aNGvZje77Yf0Uh8OR3qArL7anCpEEr8a1dujEy/aPLL
55PyqTBdLbbKGZbuVF+5MGz2k8fJM86L2MfBqiNX61/0KL1B/hC+vDFuiJBYuG6c
6jSfb1dCvnoNz3m8fOTY+pWSaArOUR04Z4deXkuvGqCJf5BSHg15FK0EbyKKMioX
jIqLWttITGk73Q5OFXjAHv6Qj7BILiDEOWlB0JVWPaQz/IXFiUvzIrHN9apPm0+t
iv0eNGOE3KXpmtrvwZuvA9b7kYGZfXA5sKJ4eY9UJwHLD+T6nL850mXgt63p+7ZE
xod/kPQmVFiASO6LR0vkGZVQWecG285ZLYVrbjYl5zaSZZ4Ov8K/J1OB0d0nUSEo
BoaPtC+swQjBubFbnlFyPRP+3teZR0caD/L0JALUo3zo8CrfdZ+DZ7k5nNfdomLE
ish1TeAj85zAgjS5UFoSWJbJCJ0Yarpvu+jRgmEBwT2B9tLvMP0tSlUhtUNVXICy
T3qjMpSrTVO7nLR21oN9KWSuwQu+Lx7kJv6SMCEkcoZdFc07PjnpybtLXlFl6YFT
Kmx1K2+arITwygBTLDoZ7zcnshQouUPp9syKIPbCvwRR3wAK9tifCtMbBGMVUgQa
bbnKp6KGTq/fF/9qtqcFQ2KiqPewA4KP580w/Bi7JOQ6F7IAbm7qZwe5K5ZNJXYA
uJ4Mvgyfqa0mk+9l4FOReNptCO0SLpF55RgrOW10IuzKRR6CziSzgdGmy2bLtLQ/
HKr1kLQ+ez/aHr8SEve7ztFLB7NLfNgaTesfL5RBiwL+kxNqgR8C6e1cc87THiEm
jgGahzlFzok7isWot8jXolIXxTMDUHeGWznBeUVqe/uRMAynTbPf65jH4qqhmYWv
JTvvgOahPtNMePjM4v59+61TyCnT4Wh74SOSaK0hPOqDXAAASjMghS7HaFa4jUOC
qLt2zWCetT7IWXf5++aIqQIe5M3f+K5tKsypvVw9oHUvR7sHT5z9EcDN0vCgoqoR
sxc7VreEMtnecXjUEokIKo9CZYVeJjgwpm4mW84DPlL52GNZcLIMnY/HTO3cZzsR
0rEOjhVhAEu+VeG8kmPTrY7lPnUtIcLidkglBcm4T5lEgPzl4FT9X4nXEmCR98FT
zQR0CxAmLlD0awCJ1GCkZHGDJZXVElalb5hHhm/LBTxbfPZMbI3EKMOrK8P5iJCo
SdlsMUFMmmJpUXdM33LYJlLWeh5JQqyeKO4oydm86Z9WWeWiyapkvmFAuHWkmEgo
Sl/eF5HsqGjO1dhbkoAx8fvr8970z3Q8g0vqaGYveJ+rV72pkp/G+NH8BlnVZsAa
sI27NC44bI2aFtvw6oE+hplnuw0cwnLZ2LQyChz/dYvuzK/e/1KlUsLRJF3cY+vJ
xLolnyhpNI25aLaWH/yZbG9wntjeajc6SN2E9atL2QjNlgn0nA7/cTSfqCXNxsua
df8vP5SuiI4sNu+O8WhfqMIL1pLVEtkOpHtspMsVETmMMwyc+U+IV5+qfAg/9HfQ
kGlg6pYRTO2nQ6b7tiWwGKF4PHOq8wl1KnZ0ycVNfa3yKUMpSPrPMdLatrBtJQxi
HHy7xgJGWL8RIPKhKz023QA4PeME2twEcL/KfjhJuULkbR1n+YBP4SyyJa0lB84p
Vixb04STxFq22ofVWOY3B7l62SG/ryCjVRYiWShAMmSmVCpx/WwYH2tYKU7nQgP7
ItlEyNi/bCiDrFhujH7I5Cx3fp8PR6Ks1Yj1RjyUPgQdMeSLZN60MM/bg1KrkbKz
3gQVhg87GGzd3vooJJgqMM09fJ338q/BRFdrOq3pGMOjhMIUHOXe0c0C1IHch9YB
QRQwRpI8Fbe6vh4SRT/NRps7BajhK/TDL0QidmxfjTxp52RpZ5BpH8RPa5/+HO0y
jQzauZ8WjN7KhnJjmZByL/deatw4thoB66QQBfTHHH+/sAHdN3vFKPIKpCKhZ8cy
zbFimOl4ugRO9y2WjwmAVZQrkPMYCis2c0ALm05UKHjbZQ2eZNKbHvj0Bxdt9S96
+Q/kfkEtOAQIxcbh/MJTr7J4C4GpzmnVq47LJXLTElOloROLcrPgP8zRTByCCE/0
VYIHULWS+2Ln01I7p6f3gqWMQFkX4QN1kUAcsKC5Ukc9JC2ENT8QJVRsPDd6FBw6
8c0oUA1oOYwNij9eJXRH3rTFEzTZDlVNMhW3U+fCHU8PadgpaRBH1/WRPlCUVvqK
GJ8mdOQYPlpll1vHtyESYbJzE81d92FCInddL4+qz0Has3HjMbCLcDdmN3prZekt
I2RI0x6SW9YNfl4vbVknv6TjIRlzLWDytxycAszM4IZeYpYZ8JAf44oPMIG82IS/
ThtLVDTT6C2I5OgocuQ7VK4UxcGlGMa22Usp6n8CG1uuvvDjaaMmWIPtbSHNjwo9
J8dLytI4KgODRj0v+38bpUr/d5EWuIHUcI4Fj0tJCbeKRcPcDzDzF9w3K+6vE904
N7UVCe99qDEHpMfiaemqJv1vH3T5Q8xeArEUPMxqP5ukE21OH1Apil+jyeETI9lY
vOwxie4Lx0l3jsTPFU3j4QOCN3ykgOFHDGib6Axp8AQum8B3AkvRx3StPnasJcvc
SrmInXfs7NGVHoi4JgD91oTCvS8AXddp88ka+f3YqTJIEXib3ZftQ5vgt0T2hNw7
a7oFm14v3fePXOXA7iAwFyvhiitDgjf7KgDIMDhiLTOSyBB16PmlG78imkTNq3iX
HnWSlG3O39Cku8trBb8XUL0E1t7blPx0A0oYnOoIEKoB6V8+Aa4J3Dcr/P9TdzFA
DuV7kHyivElt8NVjDjUV+UnGHkBjOt92cEd5NGl1f2th470LDkZJWOocK20ZGl50
fXtod+dHFMeDLRDOTHLq23vghTIX7a/prdT9SZS4iW6xsGa5VsYsCtZOCNZXK1Um
zfQFsYhNGpO8xKaq8WccUm1jFmRHNuAzHPr1YEC5hQExwoGOe3fjIVFP29cpJ11v
WaY1xD1v6oWSoFs6kFr4vc0YhG4A5x0lmShM+upGrNI9IzcGLOFOLnyyo0d6lAN0
OFgm/u+sQeTlm3P7ln/ORWJ4BaHp1V2SglyvTjS+fGMkeQnytPrce81jLBpkcsso
HktjbsfYJ6Zn/ihKkoKHlKbA9rUYLPJrsnoTJvdNC4HXvholAOJT5fcC128BKjEM
uZ1KL8KrsVdrPjXi6naJ7sg+gkee/MMiCkYGfwAYa6fnmbF4KDQVv/uIXnTI+ID6
AFlIwQUgz73tvpRF22vKZHYzJUEx6GBzfdl3/Ey5mPvGjXRWqZNVRLA9eMVIyfBb
RWCp39vB+kOrOhpfOsxcFZYxPDJACBAG1H0LD6Y7i/Tl5Iix+BEwa1s2xtUIrBY/
Cc9CQQBbtPMRtDlbJE45K5t/FDIo975ivuvC8GLrUZlG8zAYW/x1T31nuhXjbnv/
Xchl6OyDHh7p2lJ49lwMYPeAjmgvXoHZ2JUV65nsnBo+iN5Os8womKUAtFhSwHqD
VmjL+pTDYIl7oOllXuXHBRELsbJIuOeK8zeDsLBzb2fS6MIlxHFU1YYlbm/0aDAB
9NiOKqmSr0njabI+E02mp84isVeyJVWe7jaUUJRWhqHKO+MbUrl0hUQDfpVyrSf2
sJ/ImwEzKJKj/liiKyYIr/Us8Y0S73/5nifqWHavaUKqPD/NoMQIEk9zOtEvfhl7
CVqe8NAKXsmYq2XSLQN5bvdT8wxDj7i3LXyWSUS+xRRzH7b2h18bFRYy09B1kuy7
bHwmgEwY6PEO8rCMGxjT/fV2Lpq+W5aG6LwvWrqcXxlDWSjAVI8YC9bbhICnX7+9
H8jS2k+gtpNwZBX5tt/T7JoIMEXQGcWFM1Mn18eg5RKSf0VY9RQiHmX0G6T8sko7
Lxdvl4mESFx6RTpmdNV9wtDmp2JTbH0R6HT/F2bJsoNfSXWgM0fuqZ1xmYsjuPls
35QUX5nBDOhxemwEwzceY82tg5CHXCiksBUVT1LzV6CBNjHfL/HLNgtJXy0KtMjf
337JvC3ZW+tkm3fsCw+zZzylYuLfstRDld7n8YYVqWsBv9fmNwPkbYwERmaWPIqx
RKohA9BtLgVvAVuFHnGl1WFOAok8XVP7iKI6DNcdgLuL0bcxZ/U3/GB/z30txUdD
Wxu7KhXW8D5bk252YhgtqJ8q02LewPE22RhkOU/KWWV3ANZCPtsNdJuiNhs23az7
v946ODdCNR1NpNIeQHB+3f1mAkQS8WwDbq6K0V97JfJ59UxlE0IbKbyo1wDwDGyA
mAM8dJZc1vPrf1gZwVPbQgX+E2ZPTazDX+F6j8oIu5IY2untZgvthwlavtUX0pj7
pwRdIJ+wAU3gfGmoejKu2gx1AI18hmu3WRmQmlZqjz8dM/jGPwEJZCLo/k/eV80O
F9opliKEf6dQ4I2hw9sCQ6vO2nRgIqK4Diyeq9R/ssYI0zXyrbqQlpprNtrceTRD
ivMCjcHqDasIrTOfyZlbuLW2x0jYYY9zFTBc6GmPi0b/B7aEoLp8eOgz4AJIHKQ9
cRDUNKS9djT/hqStGslHjX9QFKcqemUEsrFbIp1cj8mLObBSL8qM16Fatg07HVTR
Q2hd83qcosy1KYA/nWSa8GkTuY+cUNT+BBfi1saHZ2zn4+BCkPoQ0pcyBpVhV46X
R26f4xsRqhOfYa5CSOyyNeHUj1A4v9AtxH0IBW2XaQIf1GjqCP3fYA5Zojs8Holx
PYFWflKLw5alb7P5USPZHe9UNY13Zb7b5biQjxeywL06KvJ22PCLv5KxmD+ZSxKQ
JqKFLI1CUl+vuzLcV2Ljt8rW6T2Juvp817nmKj4JYjIg9PW9tGt0KGjFIQdFi/Tv
Wmu7R3TFjZ00enAJ6IloA93rmBRCFYKEC68Ls2ur5RBtQNiEblk1j9ymXQUlJDBK
scHERVn2BiwX5DUNQn+ruea3+23VQURQz3+DuCDDkslNOHe+Xjng4XxXMrOekZ2l
Bxm53Jrpf3Uwt6ZyOfON2/RzaRN/ZMJIDkrfp1t6U10fnLbZtzDMXJRLv59G+sXY
z52pKsOiTiXKM4m5/MegJo1WRAJEObDyKiX9WEHC1uNMZhntbrrC1zvLI2pbcTuL
Po8hBy3Z5OMTTJ1UaugPXyqA/uWSbKrYnMmpH4jyMruX7DYfjflghMAofpNvh9yU
lsb9C5gvfwsM6H5lbzF19z9zAhbQ8+eoBaK4ueJea4Sg3uC1wUXB98x6jyAhZ6cN
zSb0LUu22ETcR6gq5DnCUi/xkPmN+N6ntjbl+oX2BuehJE/gZogataZj84SKwoCe
rcEuBVt+XriYowq/LJHZQ1jB03PtgjGQsuPXKLtzlO82jZG230WZ4Tvv/6drZFBr
ZvzgAC+sPP3EOUXXUSyKrdoxv4TP2HNhyz+wRagxXjxFjT5VLgc6AyJsfUcVhQG4
0kK5JFAdHKAJOB3oR9L5v1iNl1EPUK59e4l/qVGxx22VJoch510SQAoUwtOj0fNu
a8SdsOos8viEqIi8tZskUkQ44jrFocEdd6+AZYvJ1HdGV5mwPELx/G5dZDtvhO1y
6a9VpkbDovP6POZIPjEsGnZNGL9avaqjbaADH3cQ1fPcUKvrrUoLqAqAT2L/0oMM
6KPItm6uas6bjtg/Bnd5ZDcBzszDBYagkh/PFkit1f2w4rmSEmhAXa2WYR0zAkc+
GJ3XSMDHwOOYxdlLaozJJxg2zJpws1VnkpxIDeNh2SfM0/limqfMyTpmF4ut0j0y
n+lizFnqgEyRzZCkj5nG53ApB+Jd/OPSQ/OZTQFWw6XVtEEiBZWQFNU+++/LCrgM
/iWiGYGVD/AgEskYd5XRv/gmrYdtbzs+/ZYQBwHdYdOIr/3xfFz7Jrf8WMuO3tvn
EodWgKnyNCaMs/I1lj/ag4EENXHOshjvSeEDeIHSbALUWdbYWaoZGIbIu4/QLrXW
RjKuX9/B7O5x/08M7YEedpiEIKa8O9MWSABXDtocZAom6RlkWDQZqncX6zTvCCfU
wXstK4OBBGCwDJnSibbYxdjG3Vya8S26yDFVoVvDGD36TvJrPAEjsmHSJe3enOUr
eiCXNBmxbPEdh5ZFhq7ko0hTMXkisugSzgCz5WLkayV2pCGSouvkfWr6cz/u5vH5
jw+fqQQWMs3Fey8eEURZCzNYY6pZUC6KmgcBAXrr9LxCRP0XmXeSmJQQPC93K2Pi
qJC+EA6JL7TxLgz//2S39pjfSpbDYmYt+3uc3MLDmGpZijsRihHe2VtWTHHpS1NQ
xuX8i7kZPUhW+xni8ZUi2L7/goDkdV8JGJl+lPfqdMxaoInNpVkpA/8DcZeDWm7N
iqLHXWhuIlqlfhB28Lj8GPU5mK9IgWWiNdDC28Skx5u+0FWfC8UZlXnyG6PPc8ln
5YcsYqRKXzeuIU3vsRnOHlFoD5R7Rm9IyUZ7RmzcMw3DGROwSS+roKs+/nOiQxIJ
lE0WM70SbdxzqCBCgEuScHhnb1a28Njwvbje8M5EH+zXBeUmkWDe6ZZ2pUH+y6XL
IJcuM/JIXi5iwSFsqQai7wV6cSq9YlgwtBstG40MTmkWZTNuIWO1I3YiLqT1UgLW
cJIeU8IxbZK6Ji0MNUhmKEq3CmDgR4PyP5lfzVOA8HXfQz4foWtrEU/qrFNRsWUN
2lbUpCniBaBV5aAssPZVm78+J69UXIUl4CZ4gTdztCDOWUsEV7DWT9VCn8ovywzx
NRM1cEZ4M5imwQ7gu6WMabTYZKBebpx6H0NzM4yeL9ES7egFGA//oQqhjoZsZ2gv
aX3mUuz+jvX73nxGishUL/nKf8Y6cbGf15/jOy0MgONFrjUeX078RkzZn07TmXUo
yG7Qqt2CUSS+PNPo1ZrS91eeZgpeWpLdEqN8dk8JMN899VUsy7bht0oLXlMb0l7C
by6ztWciyLrohnET8EBDNd0+e/7V+u0ho/vuy+W4IrvVV0WRpPLrClPq4IGiq3Qk
+TipxfOaPdoFOhzX6cyT4e3wtdIyB9eB9iEFMAMMavmMZc+2NQOflJl2MXWWJOYj
+RLTFWPRqpBjq7nrjfm2LXXU1YJgz+jQUTXI2XBD4MHjxVkYtb4Lf/yyNUhcbzSo
FhFhZzgG4CkSqiYlFEKcJJ/H+Qzk5T81vIFYVY3W/AqjvVLdimy6Vy9Ko8u101H3
eLoVmKXHI/qnNp39MxeIwW4EymUSvTdMzYYH4HrfsZn6x9BTLroSxKTHfz7RhlcK
k8NokUuqk20u4wYexTW83ML6JL3gMe1aR4J6XLeGtogi1wh/cBdArYL7NbzQf3Dq
ujHQSu+t4QZAjhJrls+/nS3upQtpxPKs40ukftPJSEjTMiFVfUSKQN8HmybYacB7
MqJWWUs3Ld+uYtwMM9qvQvaupvmUv00baO7W8NhnjIw0TZOYjGY1U/7I5vwtrrG+
75Q75awPqNbnd5+Ke88cPLz+rnA0kTgfRm5265IGOMY4TPlA2PhveMFhk4Hyix/n
mnWxHqGurOZ5AJ0LpFKD1MbETr8N6ixD1R5TkuRSmoitY/BySeic+/eHbYACsH6u
KXGtVwVbBl1GBW7m2OH/iu2HpLRzzFBuSNJUghkd4XgNQNu6ivQA/Y8hY3VI2fBf
Fs58TdiPRnhbkKhL/HxG16JRlFk2TSq5BtR33GxTT24QkzdyXgvfpTa85cWNPGBy
x26kRgDNEIwZUbNtWlH2OjuBfit9d/yehkn+esLs3RumTcwdnHPt19g1mCgq+J+Q
3SH+30/e1Ap4Bl77/NRC64CTAvnwkK5u3XdvJn2D9akDADp9AWGwpNucgJzsxSd1
lv73+Y2jdn6431MXiu2sWB9UOqviTcHIVzdfBvzt38veBI4CBawb1qmZydV9aw6S
zRiv0bqYccts+TLdg2/v2YsADHHWl87eH50B8rpWoKYW8L4MPD7dIyw1VkGU/6rS
JAfwKP8ED9IcITmJMhktyYTJG0FzAXv3peBBrPzV2JtrDlerbzHcHkTtWtRB5opU
ghHDYRhxx6IC2xQDvAgA8cobYFYXyLYbwjFexQMBB6PXwAPGFPE0rfIjNbM+sqPw
idMOS/oHtv/UWjTBTe7eQj5uXRZAC6DgI5gpTKt3sCR4dYInkg1oRQLkbDNuXPkK
Ep98zooUr83gXbkvgQdvHdKuain5cSjGqkRQHA9LJ6Q1LrCpYLOl41bkEqNAYBiB
XYI0lg2WXYn6g4FUm3h6+l2v0f7rIegX/VlQ5arXuiWpmco6977uv2pX3smX8QUT
mm3gLmjzQ9Yi4mulnsqhBi2ANpfn3Ky6YiUKDHTHCYIv7zHQeUoET5TiAAyPNIMi
foeqNeE97xzIXMG+iOJSHQITJzgHjPiAr1aW7RSN2nodCnYPZ2SfsMHISNOniLGX
ughfQNPmifRJk6JHNXhpR/cdISPzTwFxGNPyrO2lFZdDFcV0zs7krkuaRzT/6us0
Qhs1n+JrCrvTlo2QTwsCaTaA1bYIdldL0H3AzkIPJObrq+NknBlVQ7xAwU2zXoRE
tYpY4Rjh4ic/f8Mak3vEPpGCNuOfD3uT/ouPU8lkhz0guylao0hgcRpohUlCyaY7
XjoxoS/k8jeIVwvRE8ZHgvq8DPWrkGrzJyZP0q90HafoGbMX7Ky0IV5bXuNs/2wC
yFaG+w3IAzo6ZX9eK91bKXlDsM9nz9U/t5NiSwYMA05nMLp3BwJVBAS+MluzFPVX
FS8WdhYPIXFu3o355cZ2jwH1hJdA21Fj9v4tjpPqMfRTVJidaocFyGr94+EMyoaW
lOu8YmG22wwhtTwhbOYq02vQyrWWMtW5en3LzldWb6LQDJA2FzhAGGt9Yta9ewIh
1gBQDGuRSFobMUWxadiAXXdS31DeOPZ+4Pn+kLAtMdn3iqgz+nyOcELFgF1DGren
OTxSbzR2g9tkdUmsPHPbosZleY7Pr9f1TAN+W6b52HhoQSeaM5vWBp7aG+haDs38
Zak7faDMc9w7dYqSPwQqqkRQ1kqRBrQcB/f8KGQlOOt8VDPB4Nt7EtP1/hHKF2gQ
4R6pSjKjqb74ibQ98g9kEEPb6qiyUgFq4F3sOF8wUQWEUiL5yVZonoRUI+2PohYk
zOJBapkqPk8JTQh2GvCwfSrhusmQ3xTtc5SB0iSAUX2hMOsqK8OiaFGc83F90pTZ
/6ait/0rxzSaTfWCL6s+1z0bmkMYZSev7bDrOlCJft43IofuJK1wxI4R5OLdWrRO
40YAlCwuEiKAN8/OQaDDwcfaxwJBiUs5HCXNBGKGvZH9YsY05nvsCiupDh4a9BnS
YkFnWnOPpts77lLzWOlQTBQ9A5AqGViCF/WVZJPb/7oKGS/03IXQLVaD0XM/DAkc
LP8YJf8AjPIBOqcwpwvlIG6tnVFf31lfClfmpxNXlxBL9w/bUw3G7BCoWPk2d6GO
LitdbkGEwbmmSVBgwcxJOdARvUYLuj6lnUFOpATXKprWXxVnvXLBKhxeGCwI0/cY
8/oxoDLi/4po5bgq7FE40VRpZaVvLqjfxqGb8Fb8Xyl70cSv3l3UXqsmfGLAhYLm
Wfxi63JFEHdBXT9ne/ehUfJ2vjk/vsBDTXjNKU05J0mGzGI8GtWhob25gL3hUYAu
UdhRAOHAQgsDub32KBytwLndE+ng/eBkMQFlhGi0rFo2yaOOrKA+HEhzH5ULVT9h
+WPGULXafngEQi8AKxa5/HNoET5YKFB5W7zlIyApVqfd6DUvkmFBkOuXZvxwGwhC
N/7DbjNsJ0RNAOCT6I6Tp3WIT4/Lfutr1kntb9mKtSYQ4rT0M5dzpFxsjv/kSk1p
1OplnnV+X1+S8CJRJ7bAeYmAsNwaNIwpiiq+B0grjeLd7CTp8KO6LuV834kAKDIc
4o36+HRzfCKrZnwG2PwkOEVfpinYXNyKYhIc3tqy/vx7+lOuoHVWjJolaQx4pToz
2jcF6zBGmvmWDlrba72Ca6cEqQHo2l4hUPupqd3z6X7Cz7PMicVyjCDKHvEnmmZa
AFPptdJM9fHYorGyOROwubWHpys0d7zGJpDdqc3UvZ9ufw7xVcrQBnV/XEjMQIUM
lK3uueE9DwHS2P5JWN2x3C1uEjIKPyaisI0GUA+brfpelPjomXs15zoZ83NMju35
nwojN88y5KE/SYMpM7mD7siTzdkH9nzaz1XIpiGyuiNQsVFpDwSJz1XHbn7iCNbv
BKIJy2MoBhzwOWWkTYXnRB4zlwaB6CnGDTZJHvvJuNYOTKM0wXdzYJLJV3dzOWXJ
r3XimXvzOXDjWW2UztRY2TNRQomwR2Tsx2bBi6Wh2DPK0X1Ouff4QXj7Un4VcNT4
fmq2ZfVh89aBmkCmgkD4uDDarXCrCuAQCiKpOa8O2nuRzK9JqGOqgWZ59eleZMYL
gfxy06qhZRc4HzUHBDszmoSV11iYlLu4FABfy1oZc2opCcY12iWmgk1ZXD8biJd9
qp3DZRS4cDBnDB4RnmtgIDSr3ILhhuRtVBIWwwkdvSVikdi8zt3thzAHIo3CDQuc
JTfBm33hQMK/mYesfpytDCGbUbmkMne4RQ1PuVZbvnehiYQSUv6xGjLWKW1/1yST
cqLxSWwAr3tUVHIT/2csJCcQtFYMUSWz0gcHdztN0rgJLLOj6pOrG01lNtRevWrC
8SFXA1skqH6LJp7QnPjjh42VM0KMhpylF4KJVFGLbX47LtoMsT3PAmJBDErcGKAg
qCxETDpgmaoUopkKXMJcMThhBZHyDX9qWSJWAd99mEWoJfbsaiLH5n7AhBs9w5gj
22A6OIMDzmCxDEmlmB4DqU9t+SariQMtymUUT1+lIiclmFGGs3jpTV8XOHmQbT9B
HfxtBlNzomvyrxLcBq3KZMRbJiQVfDOx4y14Rm1epLnxnaLh4n4yJt95rgXf4CjD
vsJL6VC8hM9/B+5/LW0+aJkLeEZ09yGqW05DaocqRzbm5AwdbbrhSFcFdk9Ruzou
iJYaSBd9DwEJpAHvnmwm80NKRiEaP+NmpfwNBeNNvMPsNLobGDRJlx4tPUe53d6M
rXJXrXN0xmm5lCAL0nm1FbUCjMSq3nDc9cjZazYljt/JCbutNHRU3+11TpVcLt3i
PNbG6Nx6xHzNncBHWNFvgFWFYUjWzhE5kDSA1FT2qSAldPDzlTcLuuHFFGY3QRPx
UmGm/X0Bibycz5+WvexCCQzXmzLJxdLSYcQNACs11Wapln4/B9x1mtQUvRQ4yOb6
EipbMqRlQaPQYrVo4M3wbJbwZoqmRcHuH7KTqVeBKIcJnaEk+OJ/O5ss5mTUxGOV
6ogT14YVMyH/VUT/0F7WieQz2eWSGpFFC1wHJ/eABPRUHpOhInG3L/ROq7qOaX3L
1gEHxTfpnxteRJ3pSYbbxPloAS2PaL2sRAUdyJX30E+5zq+LxZQSy1EBlNOZPuq7
DIfV3G2YXyrupznFhCdLExFXrkcaTfmsE1TaoFGwH25njUILp8qUZjDmLVJuN6Wr
p6BdoklSvk+U+uGfxyWZHZjG0CNQ2KEs+neiuZgBt0uTjtabssfXtfK3MVTbsrN3
/n99P1SoYsaqx8xpaLqXdWj03iISfLxQesCWe0xEsDp59+0T3EFitzrjEMAY/oDV
po+fXZEXVTAyO/nVxlXHLxOHe19GPNV8zgHZRTvSiP3YZcmmCx+IkyqYCaL8rrGY
F9pFITT7sb0fASLmoW73S7qNUNUXpilsF3OBEJ+z21RZBkEVHOq6Y7lPLVUvq1Qg
jGyj7bWj7MXor4JW5cG/eDRtttSWVVCXgOHFn0jMMUPq+uEd86hVjZ2M7Zq2jlpX
q1rleLhq5JvuH1LT8azlgCN4PrMYClmdHufdEeXdcqwc+7Hi1i13M2VIyjFls6Zv
GVV8VY1D8+2RxwjGioj3pS87vZFYA9QlbEQGbzTpIDKiAELmWz4S9wlQTesQoqQt
nTpslHdTCQm3wTHD43BPjGtMkC0/lksejEayP6+Qh4AXe9hvBiHUrw94Uee8DvA1
+plhXV0p0/PDFHQ0q6fOxPnFXDlHhM7Xdjt6JIZlkTCNkEyYiJwUg3yXJd7rdlKx
jrLGjKCvFyFaksNumxKukht6xUPHAzuyOPWE63DC/IQTuYDm1N9VPtZHjBM+7Qij
Ht4Yu21ADoZEEqVsWsnalZ00GBv5cEyOvTbxV/jOvOOvBySNYRatnS8eYTIHzBy9
qswXK8I1NRGoiupLtkR5rKmUkeTF6rxec/2vndqVCsw/reB3Ga1pQfu3b7kTh5ZM
3oO3FdmMUa2ct5zZ8XR4FGVn4fbT192woLJDNLdTN/aGMQ5s4bgvuHH/OegtIXZ1
H1syKgUtAAyfXdW+lcxEkWLDJsNP//QJA9xqRmpBMx3zN5WP/6GTpViSF0MZFfwk
fam0c91xvyP3YSJtvSocC9ekaumsC6ejnHe91Po4MY/mUduLcdmblgO5/XPYdhDJ
2GnZzaEGF+9Ma7tKFNDn0ieR1EOUpkbTni43p3XT+GOZuFm6aBm+ld8FIzqNPqMo
iwZ4cy+fI2whtZ9YrIHSJmb+OqvgxPuJaD764jv5AMA2YiCqRZMgqMHpcejQb+/i
2hs3KJpNc79/KcGmljHZivfE0GII7G9vZxa4R+HP5IGvlrqMy/xBq65243LJcz93
Egco/GiXd3/w1LX92xDx/VERHcx7eG9fLq6lunzZFGyVQkLsKTpxaOWLoy2BsLZa
LtUOmVvyiEJlMBLKLTLDbLLKIshKlsDD+2A1xhvHvmIEVFZwLTitGpIgdRGuXsb7
aqbM2l7ZC4uZg51oQms5zSNI0S22mrZmEv2zDtZat0bIxOAFG0HcBa1lT9jSJbl3
v8yWZ1wI2Tv5bdj2eXAFcNOIyP1vI2SMfXcFUXMo8s2RzHHj0mpVbAX2wyHASOZB
IYKj9/7pV3Ru/PJhypxhaV/d2EymYNWfzeCT+NXhcQbsQFm3J+vt8uEr4V7qOJAp
5zGkAHepQjGvFuqDqKj+4XFxgZXoOnQlPoLrn0IxqYyfFBQGBUnJbn5QGRf/o5BU
fcJ/puA9fJlp4NLXrwy9LsdMVeoCldxYf0xiWmaYpPqtbfeT/pwEVumoK3nQqKnJ
WU6Ga2Gq1OmvqoOXV5MMohK+vnwewO+kmU+QRXvQYILcHMv/AtzxjCpI0cHy8eE5
gX7EOrMirGrkAti9gNn1Y8Rzk5PfdNsxpGygSqQ0hzD6GrZUAVATuncv27QqoWcV
OywhL3fdxPqwXYKKXVT18wTtH3StoFvLYlaeNvGIiOZAexbqVO98eMcZDly1JvIN
Rm7WCVyFD0nafE8SFr35w7PlDuMllrWousKgM05L+5KXiGDqz/QMKl1rOuHmwoEF
AueEKlrkY6s5mM8ojIHqeXSZit0gidT2fzioMrPp50uYOdzujzuyS1PYGRwaomAQ
RqyyBivwdITh0xj44WTBqDBrOqfUjmgFEP3JhDVvlPJZrtKq4OzvSGrfKgKT5+XB
mzUtHdOX+hU6VwzZCtMgl1IvZYXYJOKaiEvAxUOtjEiskJKRAWbp/m1AD3ZXInBb
6mJP48huQiA4HSiFXXq4IIz8zrBfwL7IxFwszVv2nfPvFPrv8eVG1pqSMwJsWALv
W+2b05PP9tdJygo3LyzbVnn3XiNpt6e1vkrZCx7HfGvZrc/aCHhfA0bg70LbqbIj
YZlFLr71WcEXNk877VMVbSjTpVcnMIlBytt6p+A0ZPUwyjXxf6oI/k0iYC0Ts5At
uq3PUkMwXtOYOeojKAbMwXoCiAQAD7c4oPEYipyZQCOn5YaURmupC8E/AiC/9sLQ
7/lyvA9xIjIwRK42dGEbFUCGUQtWRATqjmqiVNeWkW8wAMfeccry0akzRRku0Dtr
luX+F42penEhTWWJFlFvq9eq/SsLZZ1PaXlmtvLkjMaBLpYDqQL/La1po1M0b86k
DBpGGAfflN8ZrnqQepKsTSj7bIRw8O8hI+12W7m833gL+xAgjQR1nqH/5BfHG8Qy
VkkN1C1oDD38mW5ibV3OSt5ftuF/NC+bgVIntyc5kZivy7YAYlgetPJ2hiyxp1Ud
LmCzWVlt2qGg2WDrdkLznKbazvBP4Vlk+oHLIOK9qvof1aOZOIeGYrfrZQ16uhaa
CRS6rMj+ULB6XPvDSST3lObD0NAewEBfNBq9Lz2E6M08mSJkruwXQuZMNldNaruk
VGsEe5R5WsEJDi+3X0GcrzGf0yKw/cq7GJ+ZHP16gZX7tkmPMnnXSTovodWgYBTR
zrZB5Ufr3NDOPqRW54QeeDq/2XX7Ft3Kyv2L0LRFOfhlTNdyK7tB/d1TDpDeDcEc
wk2TylvPE+w+TZ0zJyJ5n0yKaPv2+ozbJ0Ml7v7PuLKoO4Y4OdS+28IlKaQ8MLZC
wkrjbvsgerWwThmkEcA2/PuwwuTHyr/Dp3tzQvgFtuAe9sxK6meoh1Tlg+FyueYi
321QoczqkWNaTfiQzxBpvNFQ7VrZrhRNB+V6ZWH6d8hqU2tIs4Fgjk+La5/ZS8q1
jFJoGUQl2ilicJyc7b2ph2OpV4yx7dg7WGMPvEwzlPmdqs3J2l4DBOfbgD+LQ/mk
8lN64ZT0qgDCZ/kTu5yHL1jRdT+htGU96LSugalYCxqrONCP2Au2WkgJKVHIO0n4
DeUNoBjhIQu+XrRSww3WQcbKzUl2KXynKA3aLQvndA4oBsMgHt/uH5LE+GpwEaF0
eGQxUlfXqNEBVqe1REjsd9mqB5Fkal++mkjUH1FF5fh8asYeovOtxwoLW+7FWX9a
d5kMxGM2SzYoux6qY6TMpWpiBlAtssUDLctt3/R8My6jNljAbjx3XrNRqJJ3fZ32
qze1tB8/S2PdbNPrmjCuRie5enmVyuEJSpG2VyiINwhNLTMcluH+tPG5iUZ0q+ib
1wjUV22zUH1juaVUXQ62r4zdtcltnd9xeGKqcbHFPlQaeZeeX11JIMKVIjr9kzAh
SyzbYNc8KJwjkkatbhSQ3AKPQCo6bXjpqirZd7xNswh3Xd9nzhvdk3H4fg0m/2WF
PChLp49xKVZ6SIOYQKmRYxA0Q4xO6PZPBWz/KWB4JvZUWjVl70NBkzxrK/Ul/Z6a
2C575w2XlgiT1dknEK3ROopg8w+uh5hXCDYclwecWyeogqi+i0OWYvlZJtk6gXgR
smoqOkuo5I2qIEIXK429Ai/x51127whZ+8IC2efvYrZVXw+VTaKGPy5Apn7KPu0X
APvay/cxZf3P7DgBOabOlOriCKkMcngvmFbh20Zipy2Qb5egB7MrTPfuRIDbJX8z
qCwe5tWe0LW6CU0999dERF3xpfEdOx9OYzFVLpYjqSDCPvByiO9adfz/epCeQZaD
I3xL8hGaVgWk4J3gRCdQu38jqKNf/2r94nu0Fc+qNYWNB7ZU/Oz6FBcM+Sb8IWSz
W+vQmlyLrtO+HlP1TZ8Pvi09CCCrP5BdJx3YmOBS6PZJR+h+zp/stTQ4xp6aBxyL
ZuGL09DRPLbC0Rq1tyAdvkFn5LYi1CdtrWG6RwgMVrr6NgPMfhEfhgx9unSo2R9Z
d6a7w4IpONyira4SkdP3X6rn4wLBGnqEQzryscUuja7ZMxgXzBSyyAbZw9SVDlnB
YJLy61EZuoHeUILnod75OEc0jGOUV3KgODPF6ATEuDNhE2tNzwIoizEWZNf9EZg2
EFyimpB+o/kk4VepxdSUdHqeQpZApxwYQOx5dR9jIdRFPrELHWAe+pxQxpfHVryr
t5E4OFV0z3wp/5cvQ9v6cVLSTsf9e8C7UCjINa4USg5KDUHxct86dwXwcgBkFyA8
AGpsQtFvnxQeSXo8e8nW4FqyCqf5eLEkyc1Gx5kr5j6NJ2Zvgdgdw+mjlpfDgQNy
8T2iZuA1UlPojwanJXWmfyAMngzLNZRvnUbJOl5SdR4yJaJFpJ+Uh845bk/Kjedk
0S9styybS0nOYddajvQmbE95BugJq0s5Rj9lvePisFSF97ERuXMwLQ1PjiEgcI1d
Qcjq+iitz2dIl/5VA7BAcvq86vepMB3YVSu/K4OPABkwRl216QDzweILjVR3LTX0
uBHa/gHY/vcmoi3xXqnmdv9FP/qOupS4aAdCOgTXt16Zl445EYQ8YFayeA08RFEY
5O5mHK5sEPw+guRy52DSrD/l/9cldx6LB9hzE0gwTux0qMSTjGTiv+vNfT0FWQIP
/kejJ2hvV1Dd/VOPxgiustuoWyHayDfUZE21eCxmYyuVBfnM6AjDHb6ZuSOlpJLK
wSu6ZNUzHBDHiPnlhoBsroFs73w6TZYW1+8By3aJg5fVP6XTkJvYZ6O57bQmhiG9
2GTE/sbY0se6Zp0sT/ukj/jaeegrb/BtqnOvIktASNjgGwz4AFFTMNJ1sK5rggJ9
inKdSSMc9rLockawmNpm1rncPxM/CTA+BMPUaxAp37VIuH5kCXULgdw4Rp5iSyQD
5qZd3/0PA25GLb9p638+JZUPf3IECwrnlaNT6bx3QH9gNRGzzdZNuWI/fEQ404M4
kGCc0TvHczo9h/AONLTP+/I2+FrfdFHjOsuRIm+9V8OSZ21+/PhI9dAtj1VnYYHR
KKW81F5jPyzoot+2dPUdVXOT7Og5jqhZ4VuvJ+Pa8aLGZJ8n+vIpBFMc2xCceJZB
1neK/5r9sNSCThYLfGE+uvWCZmjr8yzaml4WuMWpOYqB+w0yETMXjbGNnLweSB8D
yEmCbW9zqiV9d8pGxehZlwa53vhuDLknGLsQs8xYJ9npEa1CQXlw0wNknc9kFIFM
QIJM4c5Ia9zzrIu7Xb/lv2pCkAiMnax+1P7WcEESsJPaeGC20Sb3avEqoEKEiCK8
ZFcIn29yUVbSJGpoIczTps40nyB3J5XxfmczPciTQr9WpqybDwDFj0VRhLjP9N04
lviKC5L6IjMTikVE3GiFe54KUjvv6SOBq4o2f9q++Qroywwag04zG9RBo86v0Rtc
OevAPm/2b7bgfVHN5EAJM3rQ0FMWL+eEolybyaadc9vz7mel92DkcrpstxEEL9wt
/jdMy4tn/pwAn+V24532ADUZUuTgJ3fFqE3TJofDnralauB4XDXe8uHDBG6zPAaZ
LmypmK7uAmbDZxZBLlq7CwDLNsuQsK0E1irXdO8DH8chwdKwB4BU6J51L23WwJ+9
I8WKNPm0L/R2fa9Vaoc92kN1Qw5wowk0U+R33I8HLei7AmsskZMthbjacTKUvITR
dP8wjPM8SOMUWRi573gwDNGj+d9+TUSKJrDlIFvjmZoglw5S5UFDAxVrzNOOMFoG
/RjxcJ3od4294BDFJWyKV2yNrzJwyKDJCACI2CLSdM5x+6b/V4FO22NLYS/X3QwX
fdS9ycP9+wO2WJ3oSZaEqOcdVBAXarDllUHxGJoGrlXnoNzyFextkYlUbhbYjBbQ
1thUF1S9qLOuix3/NX//vR9uNESFrhZRT6sdx+89EJ00g0B3QHYrMOeXBU25k6J9
GN5PTiZM7EIBnyt9QZ1yncvY3zv0Mn49rA16lpdkoDl93+h/n81qWrgnwQ6KLRhd
6NcZKX/+/lQ4vtn9KMYbX+YrISfaScn3eOCRdFUV4cJhS/hnZQs3KlaUPssYT+L/
nn6nLM4ZqQB2vJFB9IbM7m8P8DcIFMerjAsWmpXVrNhwQHHsX55E7ruai7j+uzZy
H8CJ4LgzFI2pf5Tc0fjxS77iX0UlmwANMyLqtOYzM6OhpVBnqISWIOMEKVkE4tal
/DtNZzPr11NAnD/bUHIG9mDLfziyP0kCQBjy6uwzycnDtrmbjYy0anPUBxeOjZ2J
KPH9YUrsuI+jhnHFwMXos590UYLpVhAhYGYsJTxVK6JGVJ6TKzE3JDIOyp4xDzuR
aXG7pHoiPRbx9hw1fKctHghOOFeqMOJ5jcDVJS++2HKE29Z5eg5CgigvCn+CCb03
wxEyWSDWr1kH+jgMJ5LzRlU0U/O+YICm2M0kMsm11mPa5pIvRFsJ/C7cJUFeCByK
b16SiTmGQ8kKn9QzF03cYq0FmL/HhbhN7iosHyZ4RylrBC+Wn8egMuuH46eJPWFI
9gKqHh/FDUBICcmU6WWyFhXyECCvZjiIWFgqG0BOaW4YAl/EwJuZJWKE/r6nLN8/
zykq4Y+XB9CTWcKVdYKi/Rn45jMa3TrCkKj0cBFR62Mg9MTvef0A7s3oHS6s9SZE
K6kc6ut4DcdopRjRtEKQ+vj0dd+X88vSUurMhpa1AU54DmsULXyo6wT5o5jwOebh
SJhXY5mGYkXX2UFeiOJHM+OQOifDb+QeBXI3wjxbK/8rMJ/a+Ev9TVtbPYQrpvvK
SGupQ5JrfDI7yAUhl3wkG7V2Vgu2NIX6gAqD3IsSkTxqRlU2RTsmKhZ5QRFvcNmD
twc1UOi5M21SItUlx9m2jocm04AL+LTr9615g61Gz+PUUCassRvwl/5hrbPOBhBB
Gd/I6a/2MPOX4WN4mUPEE+dmw9ZYvqpoyk4cbMByb6nJ7QwBm1Utl9wrRfu6UpLf
K+hCKksvLIzplHrPLNI/EItPjHiminJIXKPqZPu/8RKf/BpT/nDAYha5ZtyuIQGh
8gkCUIfLNULF7lgTlFVHT0MfMF2Q5DfP0MRcFDCuVorYP9T9mQuW/QZpIg+7LQgQ
yGLy4mq2GN8vBdmjj+AJZpmAZqHwcYqpdvn4/FrxWi6ZGgTw8DRLXuFAlDUF0R99
1Ho2KmB0MG6shuXB6vpPzV8hou0L/XOlz1YLWBfsF84nHivPnExZQ2rheQ9e5QOe
KpZJUILP/PgriuncZzmNdqATx/47/rOiRbBXCfGBS/YehJMiyNsEjnssTlJzSAmU
5Zb+vl4qFqbuteRtbn5qeXYZuk4gx14lzrpFUq8l2/4fFvno7Yj2NUz6Wh23NTFI
O704rZ47fcKtdEJUQ+Tqtg+/8KPVPUby983k1WIx2oryRCsv1aBWbh5m2W8Zz+wK
Ds+kfry1KQJxTM5WlOs21/ze6MwmgtfuBuwP8tNTBkXI5CONtkUDlW0h2Oc2oCvN
+OirXvZAqdWevjNHboyt/dm6uQe0F55YVK89ChoesDtBwqvpymcq2ISd8oZW2Vhv
qQD0yCMLTTveRdKRnQgqbd/+tl/fFuroO6r+n3AGqkvFNO3XoBugmMvnb/3wn7ic
IbKAvsnpSjNN3arZsTfdR551DN0r0WTQbubJHMAAYX1LxlKD3sIO6wmONqnsONmg
NlC3iGuMhCGiuDrlRSvESwgvsxQMjZ5MuWMXnA3aGeEV6NIb/AOzIpkCAO918fmK
scVth/a+0wLoqV1fKZYyOBLg+o4v4Mz93Vl54c/1BNE1ei1kLbu4TnS8hxfgg30s
yAvPBf2ce5KhHf/2exGrgp6FW3MhsMZj09oSTKVpqKHj3GT/hz0WG8Fgu/N4yOcc
pgg9wnnpTRuQBOwiBNMPKKR62+JY16ME+74/5SY9K/aXkQVMPmrhHjkWDxyk2F5s
2snUlJ4AJFMpCu9qmcPbzMkJugDNgFhbddBqzlzie/N4WJMZekDRuFWrkZPZcxRn
9mrvD2h9FaxMWOVZQREi4H9HJcugvv42Npz/hiyvdtfk3duu+qj6e3ONsGKUH3iZ
Jwllap6v6QAEw2NTJAPvYSZa5KWGRkI8f3gwsGWXs9xJZbOrWrupOBm79DUvGOM6
oNMOTiBcCMMyuIdZ170Hg8pCTL8a3Ovd+/DoCdy7gaQihPTiJGYzlKRy79cEg+Da
22anU1ls1ygHTXpiMbEy0168o5Q9h8moaEV+Vpo5IfGhCVfbD4G7p6ZnI9PZGJTy
911lI4EMyjoswePaJw032rJDc2AMz7+D/ixTq2u7Ul93jBVuoXTVPjtsIjBHjma9
QoZjATSgI6Im8ewdLaVWCH9bjcaSxJobbl6xS64MNeSYK6HzsjBbsTFgADV9ZFHE
Sud0gI1uTeRw2hQdQQCsGKn+039Wn0RS51qLeHGFXgCX2wqFpqBSGEi6KcX6dxfD
skBKCMqjKl7kNgLby5IzCr29YI4FM1aRrDkjn634ycmZV7gYJ/aHNszUAt4EXXFl
SDwqDSbTub9yiq224kilpdr6Fg8PH92A3DEu1upwz8rU+Jli/9/drNUxtYTG1clD
aZ2Mq1lKaqQ9dCL0I4Lqf/Qe9qjKrJBwEsd66QFRXQ8p2iKluGE4iTL0TvB295+L
WPI7rHOKQUEuOsoH3TTQh+8X5rHY5e0bBm6CTtq0yK9v1ZmrXW+D9NsHWktGNFyF
eRPCMHLjTt/+5ToEp+kKYaAmQTmC8BrOjxYa8wOv1KyuO4yrRa4E4lGIrnGcYnk8
XJQVWLUZ3KZFIprEKv/dU4UI2v6l2FaHzdxqsj8zc55C+hIa5Yva4w11KOm4rTPd
Lzho61mO46ZQzzDe2CKz8kudr7EPsdRIoiIh7aG0k218eTuOGs/JGzRZv/OXZGZM
lO3Ot1j3gkjiUOf+aSPKvQFksPpmJ7wO5MwSZLVuYn5NYKJA9lPh0ue0ljV6ftgi
0DegZfcERGS3WbTkSz58yn7DuqtPS57ImUfT9DkeJ+2162K/faLmPpFb0I/QWo36
C69iyfui3puIwkHOLAsHjxeFunNx8ffV7f4LlnYTDCei7JV/Y1rVjtXJ/s9SEpCd
lJXT6XvRmgAmKjqUUgs6Ck28Il1Wnj6u2J9CVh2PsswMTR4VF6/4sIShDG+7hT1u
YqCSoa4ALQQQyG5zbKMh2i+MRDsq3SefcCtx6Z/FEd4BSFUClhfauq7Y3aziH3I2
Qvlozlj52xuLSkM1F3OTpyprZ1usnQzkhfKpFHLKPLxvHWWZVXELhkDzNOdd7OL9
DLlkGvjTmpLDjH4PQkleUFSWEnUQaMui7DfyhvjVzdaRMC8iPZy2WrEYEZIhKQ5+
J6cS8+7kyfipnWqJQQFs8evp4l1wSa7oNsGh3fKXFBWUf4c1wGWUujBOACFNu8ui
MyPYNH6SEzv3Ti/FlVaoV1Lgy+gj5/yt8bGPci78q5/kFg1oi5qQfGJVuOqkpJ5d
z6zBgHnUJLkwKaUyho2VGnnyUfSVa918MA2Xo+XDA9Oh/ApCNg1Ib4O597ebCuyX
lIkzQRBD0CrnqTDfZR03zUZ+N57QVsxk/SlfmZWal6257gLB8F13rK7un9o4DD0Q
s2bR+LHPxpp5Uror5bG9OsjnanPtcELMIWSBVT4z5nDfaWbjqkaV11MmVsCi0a+u
v5XlKbxEOXECPALEILwR33rB7JS3vbY+Ja36FM5Dlqejhs4tTWZnI+2K9wY17m+0
Tl/ZipY613iPyeLvlJQlwK2yJnE9Z1p15lhQOQFPtJMAC24Pxo30ONBYRSR0DIP2
VFHFljl2Od/7cQbN9WcB9tNVDzF3sB9nBzLryGpmLXMANMYNwGwAOORRdWO6OPrq
spZzBdFNK0v4yKJ+/jPKmcTK1SNSnRWB4ocAlL/nBHgZeCzQbeQhbKcg4cJuHQiY
dBlFOOh2Mjh67A4vru4Lle+5nY9grd8NqYF7Y7bbT44j9uqKr7hR1Jd4OOnOLP2o
I7w13bpGuhovpr/kd7Svhhmhh12tLB0K+zHla4P49jO0xYgG35DU8pARS+M6bs4Q
HyN+4UFJhwVgeK4ZEQ2Fs7NsRF2Q1k9X+QWKXdzVyajtVwJu9UqbyFfncHQgEfJ/
GQ4P3AzBV1Ok7WCWYiPj+/TbuSz0PQTYD/CJ6VTIXRpWzkUcjCi/G/qAgPRmP5VE
kUORt2aIPs0AmwPG5P/zaCUWwd84Ee/Dx/dCGNGGLE8VAw4MzAAz3B6X+FnKZHGw
3jlKDgQOGPBFVMtIgo5zHOqNIDaPrrZw7Z4DilZtJTguld1YqUxuJqmBkYl2gR3v
RLcOz8cgYnf836KEXI7xR7CyEetY/cRNH9dOAhYYUGoUhzoPzQjbCFA58cKivptI
Uk6NICbRwbpz723CpFUVRScJn32QmLu15bcbIPz47SwtlOaot4SbXYCgyTRxXEyX
wC/fxmievWjuqSDCdqgdEnuYqT9JlGyvSZf8lNr7PO2Z1f+g0sYb+mBvKJeLZYDm
hNhQwQvwboF8soxXBL5+z53j+sDZVohA4dUTikyeIbFlOEoE6fOpRLkPehbWf8Wd
uQitUyES07XzVbk4oz8D2hxpCZGqlUG3ie6MX+qo+HgHw09jJSqi5oFVD8/uytM/
Y9cJBk03kA8e3gUXhDPFKmTLv2SmEsD7gbxNIV/VAd9nASAO2mYyYYxpV7hcC+pI
M32JzzvdHBVNnS8+Y8W3x8j8s+OY00n9igvegZOdROWFF8AFOtZHCo8dYt8biJlz
DRKMtKLVNekDKtD1aNY1esZBeUU3bbb20/5SK0oK1vAszNoD5KkF+LouF5y3H4Ku
zvUVCTTCbbrP6nt5pBMVcf8UEoPjEk5zy1nyijdyrwWlsme9ofnprcR6u7OBcNJs
qpOdHsSvuvuKnn08l227+MwjD+DFIFAkl9+UdlWwbQ2D4hsTHAfYe0+XgJCJZpa7
IX6Axp0tQU/8fsrTih+08tQ/47GhyDGD2ZSd5wDsi3kxtNMP0OHMMbli/wXujx2D
ejtrH5NDdWGOaluTAFsDXSq7lewxsVXkFSmWtcqX3LiL/nbSl1xZoUxSjpOor1Zf
CvYDGgWUAlxMfvenrYiNwMusWU3wEYRqeNQkUIJZQ36oiOjfk9XcF0Z4S8tQobaO
16NsRm2USkxJsYgFqxI+lsQ5bz78RcpjL3tlsYEF3ztQIJg2aHc+rs1d/hKp/Uoh
mx3H1ZSilYLgDuO/oPkNFWJeaGIm6mUVBkuVzRijHfkPMhqGLJ0PzKQi7G5T6ByS
88KZKRjCLr21UAVWP4Cg7yccmaKr/Or9zoESZumE0idRnpSGGqWj8hyzRkBuVf4Q
pvP/BJnh1FGUPmLTCOPktrcSOO4CiDY3V9JYC31Py/27aNDr07Bzh9+fI2LtiXwK
hm3gG6jz7HGl+67Me2gM+Ub7ZXG7ofBVk6BpIMllrBvYk8gM0H6j0G2jKDD/ucoK
BJ3snRE6ukorSM+7u+tpzTZrEI9iZPyD//CMoiqXCl2DqMCWqmhZcHw5ZLUgmt2R
v9S8jSLhOWGCUpStIN6wEALupQuvs3vly2QcDYWhFH7je01VfdbsGbDt7tOBG3NR
Nv6A3HrEcmvMcF0ZbsQiDhF2WN3SSqBYhDl/UtxP9p9XEJ8F08Ok9vkfL+Bko5W+
O7ObeTBp3QYvWQ5p1W9N5QkVN2FGm1B9t618qCFYGGTkxQWYTUnFwXOp5dNptT83
6WU0+NjkIP6Xz3dAFxjwh8xn46a8SqFUCdJwx9gnD8Eu0j42JiIhqUAkQh7YEE2V
ml5Bpw3VuJYwskt7averW5KHTDKNUDUJWzpCfIt3AAPGDXa00UTdmnpvW48PpVg/
4pgADmGzQd6e5XViW6zGHB88e5FyTOcqm5o/UdjiZ4L6eSE63rN3dDeSL1hqSPP1
0dfuZwemppqHqZ5ZyKz0jV/u7BWuyNXI7AIr+2TpGBeQxHQkLlUH8UCgl9ArIddT
h3vvEwlqJGMS2p/ku7YMsvW1DxM49y4oAxGqbnfbunuEOnWH194UUOd9MG7xR7cj
TErn1bLnTrwm8pNg02hINwXBUBV6R8tySQZmGcPL2L6kIdFAWhRzhBXzTKedtjQc
fLUEhNgyHVKbshTF8+ePnrHLjUKwDywrIc0pE49Bo/JJ4Fn7ADuHA6jvTmCB2NNE
aPmMkNObLvFqie1V44lbvpOJV2GrSn8ARzmIN/CNJTaEnRfeLFWLGsQjtXLLqBAS
X5chh9n8xat3hpaIMwSXJc6SIfvGHs4CiY076PQa3JS9VAdFaJKjPDTeSMmQlDFD
JDifOQYzgeETN3qBE1tDASAUEBFXH4sIwdmFJCalpcvr82ygiXZgLMwIrSX34oC1
/PgLaDs6QlwZlRRyJtwo+AW8kwPDKLuwU8ijFkZbW1JaboLZB7M0qQKSdMNcuB1P
OPFKVdyaauYTEnqHwprx3u0YFxj4WZQY3Zq40hkdtl7rzGewhw9c9+Z9b9ATDdS0
2/YdAVkJGmaiGIMwsp1PUzkTox0eNrM08E3lxt0t2EmG0FuWERpZWfGKb6o6Si1k
WVqSreVpZpQygSLAXaCxLy7DgZH8A1uOX/cMuR4yVP/RwEB7M6ynkyN9Nb/f14nO
j0d/5FzPWlX+E6LYqDFMGz/RNkF/B37IsSuhNlaSz9ZVCHyJ2DKLdf1eN+MkDY1l
N8rUuk7WrlQqf5dvFw/+pZTfLOVKfZf6SEWMePSA1ZdX52FoyjlHwZGngBWijKis
UKwEGBBkIzYxeinq6t+AosSDKPdF5SIj7RiaXdHh4RnMU9FLcFANxfLUMip+dwua
v5OxnSUOYaq1JNXB+fcu+ALOpLoS7BJTGosEn79yva8lt4zBv+Pc/su3Ub7ugMlE
f6boFinCIB7ch5MkVlnnItkr4M2Uey7cUwDo1YVFZobsXePFy/2U502jG6fY3XtF
bXQdQvzWtesKxRUsDAWlGqnfzbug5wBKF0fTdq0f9dAz01ySasSR4V2HXk5sTVwV
MVlPccLbFemZDcrKM2X1FIUMDM9cDIFJJWFZMc2PuC7MYnbGz20D2f0hsgJl7jCy
kJYXvITelMCU4dClxwxw1vcSRBAuylp6XoF0cYbUoILjzZ/iQwGGvl+3RcCE5rU5
HWLFg08I1YUOeZBlvGfa9ZRxlCy+NB5FaIVFyQKhJnh8SuM37gJuTCZTz7c1OG+5
WWwqK8QJPxKU5mhiFCw9RTuJS0QJfTaIP+MtXwjGeIkhzo+C9iOC/ZJjiJAnnfKC
KHfmwKpJsNwKmD4e6BSAMkbLeGVZJGLGZmwi1X6DKbCAKxILoJ0N4W318Syb54DE
CUwN7Kk3hyHuHZtyKRg5h0Z6pdexC8aoAN0oBZdp6PsaA9Auw6SMUK0rSotc1Hnp
nvvezRnQWVCO3fJKSQJS/zcZNSUG5Ky5x0BrzlLEnvxAujft378StIz1VTqSIN2j
83qdaNlIdItoPMj5DJ7O05pLrDnqIeMDtlb/8f6DFw60FI5i+lagKiOhAsK9wxum
f66Ik22lddODksrg3bkpv7NV27ahPrGjaUu7xeAgRr17+Ewe/mKFTcNePof8Ode9
h+0vEeDdagLUyieACyOMnlVE0Y0oSRLc2jKu0aBeGG0AuSxxiNj0Ocs6ycmU+SWe
f7wpuTD/BRW5V2/v3KDIJgHTS1kxQUgoSLqaBxSIK7fcHxuuOB4tT0Ep5KbHbSQO
aYZH4zR0/D2otNNiuq+OJclgFPqnZ/N9dafd1xLJqHurdEk/37n9AKEMLXV+x1+L
1jp2KK0/oYyfaNvAyulJm78tlSQETdf0IMzYmegi6iihWBSpT85+BM8JQNxzzoqu
NSKYp3q0fmsp9KUP1kIdEf+p32BMXBPBVXH2bJfZcOo8Jb4kMjIqymfU52dOx5lT
c9q75oQT8sK6J2wjO8083cVylFQo7SrvSd7fXPyvQk17YZ0QnRYJmmHEhU6pUB1Q
3yTYHdpmOGKmzQvzTxtnR4X/5aBGfEz1MyQbn2PmCj2911aQdjhUHcqfyndpaG1E
ZY2aDsJh3AeNnGqIUDsfVQRqPBVy8hJxf5LJy6oAB9TR4u6r1qIWiI7duXiYUyaH
KA1RBWR5thmBJnqRzXGYtTsIe0hSw/JRTuD9QdQRCD2NuzhyqfN2JPsEANqh2zWj
qJtY9hQmgyMLuGY+4QxwjwkNb5L8hRdufUmgwcBGIFWe4FafFb/TPI8isjoNqwlI
Wfwdd/3/E8meNnNNkrOopaxjsr+GYFm4hyPAhGY5X14Tds2wQQUc5KMOel63UEnt
FAcy9vi9+wEpOv47NkQAWvjxJCZRMM3dk9WJgEyGlpGkw9WNpCe5kWAh3k+5aZBE
/ggqXAUsblubIAWUq13lTAyaWR5trkXQN6hVPN3UUzVkuJyekzrBt9x78yt81QEO
Yvi+HYhVD2sa2V38ekKqVA1OAddq9n1hytjmS8rYo+sGgvEp0WVkMVYmW2uGrAwq
LxW+uOpQKmC1m91sl0kdZiSP52uf/PTzZXT5ISdSc2QxkMnncr1boY4tlmCr2nh2
rqL5RpHw8ManOkvoS5D72FtmOguvnN7VxiBwqkBOn9FA4T7ny1Qx0pAfA/z2n93c
H/1eAam5zb/wwk2oe3XvOd1Oq8TX73KZ9uB4jDkAlME3UZzV0kA9/rz06gI97zse
zkruuYXTQSkxg6sy+iAipT35NyfFf0ZwZfXhkr432D0S4/eROCjBt7vO0yP4vD6n
riatdxUJ5hQo2BK5W082mMsbuAxzpz6k4IkDtdxMWujTdVt1be6t1tw9L+6Uv7Wa
rPFXjfQz5z+F50Ko2OSVncV+6wrF98/G9a1dFCfeVrvn8jx5tbwEc+9P8J5wFhOZ
qynWLfYucDXFvTwU2Oz8/kqwsoVoQ+GG02zkWkOlo0knQIIBMOL2Z07GCJ7pWCau
8coI3YUSVTPGhxzTgn4WPxxGvsExjQwKhi5SsNTKlaRfDx28dkzRQaenc4XpI6kY
EYC+wfmmGvXDwZhqIK293xomolL07NDf9Hv6DZqz9eiIzgZ1UJYLVo/XVe7B39YC
CIylTZeruSuVh9RUwkb9nDG5lyE/XYPwduZlcm+FdUwXgaqCaZ/NdeA/ThBF1e6L
wUnMluXi9bLbMPn4oj2fNxfUiPzDt7yaMLBDoOGGsX4kd89NmFuG1WnSiIXt2v8D
iZEY5EUIjT+/FjEbmh0hAWHQNZhPsHw42vTICFF8sLDy3WIa50Z2thcb2fiQmL9N
IFtmdqAt/DJy1tBWz6h6fE+bOnrAkXq7V04FtI9g5cttG3JzgDSkoXlqNSSAKvj6
a4L/Tlu+gduINBdGaj7PhcPVx5UI8aAFPybqueyszTSFH6AIQvlfEhg4TfnDy6Mi
mRkz5x6UEfWBvdMgvEOUDqEjbAPhwXM++CNJ4O/OJUKAoRO95eJnR8ckqX6ki4TZ
/6t1vwQFLERfZ2HPcHqu4JOYfwF5AGF6QthsgTyvLDnP1ysgYvtOyOCYSm0kbvP0
z87/E5Ex+/qaihwrdT1tbQ3opCufoa6/Ds0vJZp2GncyiAegtAygRHzSWuJlzauk
0C2XTEFaDbt13YLQq0A1lwt0lVcJRWAY7cVmWqn7i643V8+3enSWzFGteTKFeLfY
zjFnRMxNKal/wsN/88z1tzaU2UlsHFkdSD68TupOzwmAOwmpFMvvjCTfgSTJM7LX
3v6lW2kmB5KVc00y4C5tIjIJuvED1bKWOvh94nuUxd07IQOGUl848FMmhldy7Dd2
4Lu1bqXQhh2+TAtQPNbKPPutMP15CtNgdFY7UOr+s8+k30Tpnjn832ybXTEVPOxu
L//Jjeh/K9VCse+S9TSlaQ/oSmokjSRMM0SxKsjwsSW/3lj8N/eS4SFSY1nBsNLP
Oab+KSpjwz5rv7V0I21zn3Qb2cHwKj+Lsbj3awH25yGP9UuYUa3ysHTi6aoZymLC
DTsJL5olnyDzOHYdGOMmM9+9x9t6lOGbbNezzV78Fgb8aOR4s7qr/ue1kmTojD9P
3Qy9t/QssOm8rmuNN7KamMgwyBCuJDBRLzKWc0pdqZJLTAhXvSgB79KF4U4asqU4
y5NFMHdHbm1nyjrQG/60J5jOe8OTp4VGDb/5/9kp9WNSkIrAUBQ9SVkhOTJH6I8K
cZBE1zmpIyW4Jlp/aYXQKQRRz1lMMf7YYEgm/Qru6fV2WVbsV76wRXI5l0wz575r
gb3OgEWusGS1kz4pvyI3jcQhk7R6CVQ3fgEm/RMXG3U80DdGbimj/hndrQLvlANF
JKGi6pLdF85kpceynlX7V4IFUkDN/Fu1TyWZWvj7J7heN10ktkvNADs5Pjy1N8dd
0gv6dJi75NgjQREhs4I2w+LhtWi7aTcyS7Rau25viu/hIMbFMMcTDVn9w1Irr2q0
xkLv10CUnIVvdznSfN8rSjfQ+5+MEAzRSFOI7CQuDbe1T5JGDdlf10/EXsCTXc0s
B4zBYZuEEownXP/5jcIGHQmkP1nZtcxV9nx3UVrbrZSwV27dBLeuD8ghPx9Kbn9K
CVtA2KH0dxL41qCYH1S2uKbPuH8d+hcbl6Hmkrc0a7N7VLbZlmLF/0BLCdAlMlFl
YLM1J4bQTk5eKTdV3QgVjqlAr3ikQBxwV99vRUlzEus8DrPFjNva2QUaLH9EFWyh
0DwaEBhOa8LmFGHpx1VuXol340rsqQsBHJZy6AH1H1lVq2z8s4AjpmMoVE+GB0SJ
RU7B1YUykw/Ck2KkadRYkUg2jCSko5w8hypTAuHtsjib1llxS27WU48LctMZfT73
rC5fRDnCDfg3Jd8xjejVT0W7b5VquMxme+//aYVZdNiNwPtmsuU984rmJfhNR7Ac
wvz0OiOzjLjddyAMtvQ9zf/dE0Y0GdeuoDsMMjj2gMhQDVVaeKfPrvcfl6U18qHn
8fKl40pIz2nEUw+b+AoOjW/n2gw9ua+OFpargUSj11dri9bYP2GYSrt3Reus5ofk
44jlDTK1bhLJL4v48ldoXQ5xdojIWiN5SQE1JVmQURwrCIuJPLhTxBs4IWGIZtt2
OXWUip+61o+kpSi3ZKdZ8wT0LgTqnKpfCuKd2hMoyZqDp24qjP0h4q0UCoYumOo8
r1a22vvv3f+sGwncTUYFxgQuOOv3r/HpNkBlSz9JjhfV6mrUxeg97rs9wG3/YTmT
VhMldrga97pEQ0sIx3RkZyM1xRLoCQWk6wr4pEvKx8PPHwKTfQ1/OqCeI7aRJJc8
l3ycn6zsCTBfM4wWZZrIvu53dtp/Mdys9d8G7pq9QX4Oy5Ab3tUQhd16wJl9JTEv
HZm6B8RnaTS0DreUho1w/PXITA4WgTgUyTlGaiNrcGd259NU+dnuTqGCXRPS+f3e
GKS5KdKFW24B8LiRIi3E1CJmEqb2PPPJhtOyW2lY39vnomuGefeN29Pn4+U988cR
TNUQheXYArw82cPVJArdbu8ycI3M22CnOnA1JQJSDW0IovNEAhXtvEN1/zjbPmkt
UqX01hiQKtGXljimEi0LAM4o02ETInC0VcGDNLUB5ELEca99WRizDcSUfqKNNR73
MNy4TmiEWMPXhCQ6uGnO0yT/jh8G1TdZB6Xb/gKbvpMs9gqMAp3S9teYmfjP6S8f
5qudftaKAj6S1cbhsJ5wQBegPb2btx5p0YjSyponXvJBq0O4iHfBHQEjFlcAKBXN
6EovoBfkk4C/8MWDNMsxLcdLN89CoMvasal56wK4+UAXbdiSx+YbY92pHslq5IIR
a23+T+QyLu9bSZKfR2kEM91WQyN4tH6lc+EKcYyR22ajLxEuJZjNKUq6I5z3cu65
2sZ4h3SuE4AYG1xpc8P4u2gxqmGJ+mPuS8dpiXDcC9dEQOzb/M24fJ4JY4mtOIo1
ZxFGsW3wM7O1DADrY7YoRL+HCF0/6oq7l1P7wJw3AEonTfY06Uyc1OiuIxaycPk3
9a9d8dXy7/qDh8y5Vz3JY331jHXWEAYWTOrDJ0WWOAR9VU+PUQm66I+rC3XPonvk
B8aMssed1MP9uoMeXBH7t1g4bnXqnqbGanDAvHdeZwuAeyLZtfBwqRxefi52oZVy
VBotIcRgJexWBXF45C/P+FBStYnxX+0aTHhkdfuNxFAamroLIQkFfPzW9jInPA1n
e4E9L605ahMw/r23aYsSQ8LXpG2FY4xJVfgmHKpbJm358hBwPIGzQw/D2fRKiemM
8upmbH5VR68mkY8KAnDMdlpI9TihRp+d4j5Q3DvR26353qJK21Uk4aRBNrOCOe8n
hJV977aeRxhm7TGFDrTNZSgkuplh/CUU2TsdqZH0wCe4I+lZmToowaLDxQ6Rk7ZR
t4kp/kRgfSSnO2NKAokrlODtWpYTP1gppYKM9J6egp8RgHwcCqcGL5+EWolk1ZpY
RzMlES+KyQfLPG3HxbBmoLqpAABFKMHqSeSybZd/h/s3XDnHc6vMGyXo+V+Kneg9
f7EnWC9k218EUlRUsPF3EInlaWLzrEzr0zc+1aThQw5VLqsxyHhRsiYPlyoRdJBv
Zcl6EXh2rpwt+udYAeYiL2bi9KPK4/E1NiLbsVxV2at1KmKAh/MP3xF3PJejzLCL
74LesxnJO8JbAo9cw0TX1i6whgoE4L76p7G5/iYtGN5QFqWhuuRokuLXWwksKley
X0TKWYm0/qwQyKlnlFQQ9+24IjP1LTOQjMHWI4DiuxSHlwcnI9yyGhLO97iCSy4N
t23yP/B2zsYUafHUyuL4YZxSN6FhlxkClrCSC+2taKID6UvBwTUVdGdQtmdBG+5F
BdODN9Esf/xY2D1RT1YFAXblN1I6Zx5tnWj0r7TgYKW5Q1US3K4EkU4Nv7SI+vh6
PFZQlfsBZvo8YRdautfEIY35ZHrpYuI6HJbJBnzOfUIt3A/QShV4+uCDQvQVsYBF
N/hFLU3d0+wJIgnhs4JD5kVIfjIZsHBEhxsrDi83W617HDpZhyLo1IvPpEl1MHix
5q/YQ28iamuYYs9g2F0F7c8I90d28FNcIWKHagsmGGJfEGwahmJrg9xcQ5LrSVVb
DF9BfKX2GFzBTSIsxYgmWjKJ4hYAvItQwTztGIf5Fcw1zBtRE8N15U52FonqN0Sy
aIzPO0wI96ud1jwBkAAqEmrU5taGT5wNQggB2yYS6KQE/RjJ50kEZuXhtPhWFEWd
uHlHrSFk/EuV7FAb7fqLyGm3BXC7b+oVjcS4IbBfJk8VMGoTL9oRKimGwNm9jNxx
cxUVayoHm5r9Y6DcnXij8oHRIHfagXDUtFutHA7C7Gn7FIqAcrKEe+uqUg4GN743
jPJaQxWtqmwhbOftmKzwuzz4f7rEtrEOr3DHLe9kRXCAwnt2Fp4DyWoz0coqq/OI
B+Li6wxGkPGHy2M3vGiNsLpG0R3TGhoi5o2GsZkvxL6zjNNWAhsK5zTWtv6TZlP0
cSnzKxYhZqZwc20hxPZdyfnPOtq72Q1fN89TN+jOYcTGlkf6DfRcgEBvqyC3iYWX
VM3dx15LAVcm15h55M1eULnrWOupHfbaZ7IQxwge6QUE+N3qYMIw7a/p8+WCi+GH
cOZ+o7IOAnynJdBYaXonJ3ki2NHRhgrtSNFJv+bnvd2NLriBh9LHywTwiP2yC6ak
UhyBWixJwJs/Tlvwjmu71TfXyVka4mMZNOD0eLA9Nf4Rg1uzILFx6mGR/2eMNixk
WKBAUVlsmxOz6zgLcTexd7ObgJNNkgyVlxrV2xQnHkcMUEGQEbbzK9WB5gi6Nt7W
peeJvMN68UpVzsULF34UNll0F+Bks/Gv6VrX427kF/q34C9k0zFHyjBBuELjzgqB
8YG7IV5kYiAVwWGPBKac4fbdKFXbWBfmzqjI9swz5Eur98swp1u/lUcFXpU67vuu
CBM7TYue/FCuX8tNfqTWrD6ddsodNXmbaMGevL6eUsJS0nPqG/b+kKrG1iV5+cNl
mrCwBiATz2Y8M32nl0FuzO/252rLPeWZOvANROaZRDoGvsTakcwh0JXEAlq03muc
m3u+mktnRLbR4CdCuo6dNptAXmqOd6gIuQHMt0mZnVJMC6tgA0G6Sc4+pCL/330Z
MUvYl+jQVLYfNz06uUqyYDylKkNXZwSzku2Lt8GmfItQu9sdvVOYDiYmN1/j7yCV
agmNC9YRHco0mw8EW5cxXsu3YURzP0hSE8MpliBCyNMqZnnTbmjJviO+6T4XnLKD
zMaAZpnujI6GPq7rOks+P/JcEwFUjkZKpqc4OIf1vepdY4QbwhRzZnqVzngzBe6E
r3vIyTfEF6YrfEvajYD186q7sVl+0WYyRqD6f3GOQWhQnK07PDsyDvucQqNWAL0C
98c3o8gdu+kD9j3enwuchFJOsQ4kXdsx1EzBWEDkqYd/f2/rXFsQril6ioMLMrZo
bnvHREjnkKc8mTCmaMf4O9goG7fsMiu1ebYi/VMn2PAW4n0l1HMlyjn1vIZxzGxu
pU5kim0/l1z8o1rsT4NS0nKSQ5jBfQ3+zqTAUixo1AlrDH1EUGqptCJomlYOWErV
aZaoHLJQD8ablm48YyNPJDI63puYLHDVDQUPFReRcK2C1oBDqUakZF6QHLMLO7en
0HZs9/Qoo80BREBtkEtdS0TinCnqzl77xDBV7UOBJQXfEcrQsH7jl8RTe88dan7n
h4kUEzhgmr39M89CXay8FB54Z5E3YApdvrjnQzHEh6GBO01bCi9UOIzT+8mQAVbv
cGhTa2xgovHckNuD4pX7YbodawDHzD2D7ezisT1bdgRdkacspN0On+ztmRDWHOaL
erpUZkCs3EaHLI8UdaM4tOij2HzU/tHgdaAK/wHudIGYmSxSlUbPFdD5a5V99VuK
zrDkGLLC0kh/7SrxneoNG7HnyD7ubwRXaLdbDpuqyYat92fOtWkwuuMir56aPm6w
FkY++PH+s1hSyBEJeyI5/g5PpzPVCPL5oj/vg+UEi4q4+mNxLAz4Qk2xYk6YG8Ez
LRMrf0WhVL00gfDmAN71n2mqDuEIiqnNtQzZkUUNBIDZoqGyHTkB4mJeZPCSA7GT
xKhjUOMT8BbNNI8Z7xdfTdTWQRiKBhhA3Xu4O0tucLt9QzcGoHfmCaX6ZxRZkQzu
ZwVQVg0QAH5JT2eseRtYRqJsm26PC96THXENxudg9fLMaly9C9RjhXmntij1ffWW
c31qsx7Oh66aLg3jZOkPymYyBhPOu3rdh9WmnaEn7672ujyUpBrV2pFmTfXVOclX
+O3O7V/0RGq/+pfJXbRyxdg3zxM2e7zog5LHfgSWWCChxmtrXakbwp+/xVMmOyYs
crIbimeLieC3e6OmyiVtTLDEb2eVnSUUQoIr6Xxdvx4f5aY5pKpJjLpR8QHhdDpz
7kcVQ7KMDqs5KQeex/6vJzw94pAqxkVlhV/9jMFWGfkYm8yL3XBZGfMfcA+25tb4
Hqgmi1ZlMaYtJI9kYTEn3MnCxuIFweIdKEQWxaI69sAeqqzH9q8AUa8t+wFpmDCq
cpHocxi9if3Ml3MS0ehjKfHRsk2TW6IaPr4tpISCNAkQ2ruH6M2ps6GPlpGdx3wr
pNbY9+NwMcwz/yo5yMbgIc3zciE2AhlUWfNn1HLvkq0CnxOk+G+kjJim4/j2lwr8
mgW0O5bre969Q4KBFdrvUXunpgz7tyYXWHI//tGLHau1G7hq9R4Sj8AattOC3AUJ
X0figi6Lr0LEZg2KQ78hI41UDbWwGcqR/ccc7MFbpKgca7CtM2y8YW93ypxBUVjH
q3h0c1xfFw+sc3Ql8y9MQPJmq27MBPc8FD/jGhCcxKFMAOeUqBntPGSxRZ74UxMZ
JEYijUm3q6ldtQoxgdBG/AHVdue2z8P06Y1HUz6TbXknwkqw2MVlsC1OnG9ZXcJB
gkhTuxRMvwTxfOgPwyBbIwL0fJfR0kjc7eL8IEUHCI4oSW8JlDbpqgjxOu5rPWIb
idPT/eY3igvH59b/mz0PPBCidjGy11KxlnJIp6roHb+p1tdYG7Pbs9w9mSSAN3Qt
KbNXqbj1oSdM6zm1krZzOQQotDrw43vuu78yORtsOJ+PaulFiMuLmW1LT0i33yed
wb097eH7hsx/JAt0IR+1xfGCu9IWICYApOzDhXx2V7T59Fwddndvo/wvMIr98d4S
jvtGzw1ifSGmJ5F8q8+OUSDXZxUDmTS11cNXKBZiitetyNC61OZjQAekZGhn0wKt
sMvMw5+Y2YCsBxSEuAeSiK/S2A7TH0c8epag4gNrgzx1AfY7ys6eaLbnL2dmpsyg
edy96XM6WUJUCxRgoOV2k8BPTiiL3piRxTV2z7bWg7bgPEvjVUhgN8Xqxt1t3k9s
KgrOWBpErjdRFhVmAcDEjPZRwGQ1wvjMWLbfHhaLHy4I2+Tp6EuvJOepeXESwWX2
QI6K1aLqNekd2q1U+Q+7mLNBWKW2hPaj5ecg0gaNNeAijBtmsXLLTed7KyZ1t/jk
we6dVNKvacJoGpN5Al5zBIVYdRaVKrpSzY1YeVZNh8UBCDWtk8TNryADQlSXdfw/
N1VweWnk442hwbAue8ojqQffoXaFZCs9bs6LShStXElWeNEFY7gWeX7JPgO2han+
L2u6GrmPvPuQwlsFm4PJiSs66Lkat3WcVuwUZfQsUcERvvQVbZsN9asFmKymObtQ
7dajCIttC1G+H1pIJBeiHfncv5mcrHqcFsd1XLlYnQEX95/MFRtMHVtQcLnzQM8x
/I0YrIFX5fzsLdN0nIKg7pWvBFbkWrInH3OPqbtTUI5fUrU9mkmTN2vwdfetQAiJ
ROInFA6HSIlgUT6PrTpIhs30NAoCniB1i/C4LswTOAtNBnTw4hdAQxaIv2ykokgU
YzHh5rZcutBp71Dc3Q5qoCcuZp81F+noULf1/B/by9UiIQ18hbcZZah3/hemPObR
64XTdrA8AbUobpjIDPLZ6sDR+7PjtT5u07aitejzOLweb9n82TpCyzFuz52vVofb
9E/uRkATyGAK8sQt4VruoEu+89l7tJ+41gxHlonUTzCoDEkhHnUsn4RfR2Eswf6K
u6RKw+lD8HYITnRjTUI7xeV+BVMxrCrIwMBf97gLDqO8pP0NBJHQeW8gs+APB14i
da7U5HiiJ5ZIsYiv9CubsK8TAtRi6yTGW0tuC3mMTSJi/R5hwpvGy64MkoBL4JDU
80u/72AJVxAREMuT81OkXIHdT90MZHUConkiDvbdfca1YWyUlYX/zmDaimXh5jQn
YkWCTvEJ1xH4BY7Ia29rFH9Y98gkHhS00MQQke7vxiPe+VJdAoJWW8uRFZlh9Og7
GJns4YI7+6qMyojwoOpUrGAsyIpOnzSKCyzVw+cYDWv4bpVsH301aLG6s1Vjs/0L
gwzvA1/qaqSDB/GMI5YRc6qbGeiGxfisqFq9eoLSXZUbiHu5miaYjsv6bp1nBiFe
S0g4J22lrpzuiMIiIjhzvw0IsPqJpwMfM+J88UYB9IPo5X+hcoloCBN8X6kG+3t/
nQCQyQIWsWbclaaWbqneVnGyowEvNDzYfiFd5xJ5yLVis6Qtab8iG0X6bP+Si1mp
HGkje1DjpeGlDFCTRyoDWsmjlW22OadOUog44MhmWFDb8bF9O/dskR3Ffnc7CYPK
tUfspAz4KcjVLO1XjjjPeY8ApJ+5n8RQV3fEvVV6R6A6WOMgc05nfUORQ6ITXdpE
LjNrh4BRa4FtIq9gO1d6osCs8pdlveu86H7hu1kw7+WKCqNQtIZmIJHD17Y8Xhiu
/YR9ftFUpJATLqsMaD/SFm7MiNrOQZa9+NJMOlt3rdClWvCRYaiTpupKvg+tb8jy
zrLVhfrMGNuQFA0V23yvaD++VIMuwB+LxDf6DjQSHpbxz4e3A8f6Pqxm9HEHDYfU
0t3LTi6fQNDD2pvI6TvP1AsZil/k7tk6DIAs7u6xh5vuxjWqvyajmSJoUQfolCmj
w0PumHagU0wH5oi44WzuM/sLNGVl39HpkZLIj6QlRbVFZ+1fY5ptuSh9r1Xx+/ct
jgVTqRohEq5qZKQbUg6kh/oXo6RUNloSPbSNp/Lyb0FL4W2j07Jshufcx9eAfHAD
sCxHHuN3I9K0IDhN/afffJ4//A13PDJBS+29Pbok4FCcAc/jTNSRPXY028+4FGu4
0JOtT4u/GN6XEwJ4tesHeCCYKJ+WcMJSA0LlP8kAuoNxQqkZcUBTtTbbOPFpnMeB
E9ZaFuoYORtPjLKx3EO0T008Nziy3ZmtnUri9FiREltmxdL+003F652+Y//DwH1v
cIaqvsRmRi5ITY6zqivcCqI3t5I/6K0lsDoG5PMB4s/wy5BqVBctxF14/Jia+gET
8EXdvjBrJ1oLpOlsHWc+1/LTz5E/TB4n2+6GqVX53Bqu0zGUVbbOpqShgsf+3kQW
DRVOxn5J7L5YooOiiA2ch6tkhLTyroZVS477iIk0Pf5otAIT3nC5404UNTAoqWCq
drJR8Y/lSLeSByTUlEBJ8Q0VHQ5qmg+6yMtOCLOHnuzJpO0I8MB/GzwHleTpIasX
tub5DotsJA77XDcMC5hmsbKt6idh+tqLgEOCt8wH8u2rr9yjVitx61jPuGXmzh2M
kbCvYs8evk1mhfccFp076JMCSxSYEZqX4Tzjcx1pPQBQjGECdkzXJOHX7ar057nr
c1YaBJaGrRUKF8hmjmWa5KmQmqVUsPkXYtP3qZaYNtFhYJxc82G+5VI6WgyDT6L4
iwSnZu0Y8tk9pvHil0zSEe+LLJT8JIctbPoS4gFGV/a//wZrPWAJZJZNGXxWtpC9
U0ln3FnZpABU4Yi3952+GCfy+wBBK7/+NZzyWd8eKmRRGXxslJZHJ7jAcBbIneDi
VUnQBL/+OnK88ojs6hKoAJiJJhneLQPHUUcREjHsWH6yKZVX5oDlPIZBOypcAgZJ
A3F8uJqQvX6QakXISPVWGEZn5Ktzoks0dFfrS5PnrCFbJ6i/uDTmqi/h02IO85I1
D8cE74ozGDl7fK1+b26jJRtuOfUvrn7tOnVPDjJfGv09e48t2yRF7LP+g7N4wbQb
IvE1yK0caFkxqX4QHcE3Go7C/GUSv+tGlrzlhlZO15O1uS/OWBlA5vHfPDNXLX+O
/znv3gaRQgWJQztZFLkiaovt5+3N0Iq8Q3ugH0RvMhe1oXASskLc7rlQxvIJ+X6K
P/gewJ557L78NP5Bl79NwTLSElAZXnLJr70G7gTFgscbM2qOLBC+7yrpQEikd5mb
ilIfAYg8OSd0W7rHogdH8mLYtRQWqfVn4+MHGJSSuS5RKFRyoAzWFNXdOaxYkjhG
UrD11Yg0JbCvbbjF3a5ZIRKb2We9DspKj988TtkFjixO1CLGKQRZaw7hllNxHUT4
Rhe3kHTS6OUYjqAeJu0o7vpRx+RjxP8dixPzPIE2jFD9iWyBhOozGz7FHnfiMCxB
ll2U33noq/XtQfs1EPnNdx4yN0AgujpTk3c2e4zAcxdaawC9XunjSEbRRHquQcxF
dbE4qZa4zGQd1WCA9VMxZJeAjix04U1x8qPnM/5NfCULabYBaTbhXKk49jyR5feJ
GVRvzqon36jYr97GORCHldpl9F8oLxiXg9hHP3Qw6TcBThoUNuxQ6K2Li6biveQc
p6pABkFOoSJKGMpDi79+asE/KrXJEhh20ZKEN/BJt8xqOiBv9Luyey6B62PIq2sN
YU6/Hmz239umivKOYDgCma+8IDoXizDL1jt9t7fLyuLW+wu/REz1PV4Rq50Iqj6m
iJFbvhroOR5hfbhUJjQQwjyYb9cOu8RYeQ+yR//E6XD7lmkd7xyAzpVdWwVgzGFu
3P3d4/nJ//RNZJ4pXJwaLCVSO765hUqKQYufo3GJ2CtPBPmMz765VqhyuvQzKU4E
zcjcNnwkFF6xmu9vN/tlG2Avvc7QtlwJQqFk4lNZbHVYPhwzY+6XrquiHwkdTPTd
HQ9/CRuP9OkJ0wQpm4MkrZeESU+bNoOqMQAbmrzGOjOS9BUI42f7YmSyxO/UNPNR
0sJedZ3pvtGzk+E4pFuTUuXYxxtAdPtn+yrrFwmmiYrSAdUmG2uaktfEhH3XJmUX
twWT3d1pF6Xg/onmrdvEv87k69QZOQCHezAN16N/USfEouX2OPkgIUqCRimWCywP
BCOJiOIB1P+CoJ/1Q7CHD6ASgxDBt7pPN5eRMRLawqXXnKdcHnAiPiOQqppNC8st
wpl24W7dwfkxyC5hMcHZ16zHZMHDFuOjCx1czUJ5SOvIg+fz1wrQ8wG5hIZJJ3Q9
TiK7wrCCbERRk2kABfbEnx/OKju4CRMVImP47JvZHHWHl830/A7XcHnC3IwdaYiv
vqMJ+1KHcM8pSPnSvQefAGd+9C2hVUknMeOrv7O31cC1stEcKu48SwFbGSYmmEJ1
5Esbx61ChMOg8giiKNY8TZDIs+MwN9JrH5TpOo0pLYmOtI4TPaoL3xXqcqeIe7dZ
FkrDGDu/iBRlvoADtGnSSA8j8fo9wV7la3f1JYuX7uEGD6rj91ObrOP+wi2vFoC4
ZreI1ZwRxrtdK/LhLGQCoQEARWEBNQ5sMtcgMgPxFjvdFNZaNDLJRZHNKVx56iV5
0/G5562zMYPR3cs9XQGAZPfn6IzOcQH2xQZ9hXBOxuoaSAuqePvsWtOR5UvwB3rD
hPcV6Z+Gk7HBOXdpkaKJPz8x3o4uidyHC0owmpiwR23+ExiOCp0nEgub8l4aEvoA
gPvW6oT7YQG0MN6BC2OabWL1Vb53u+S8ULO+CpKCQRKhIrfyTXnzdPoeimHHuPLZ
DFYvonaz+E2GTqbmNIzDaETnN92JgPgJx0g5h3U/lHVuc0pw3Frl/l8KcUHRvU2j
OC77KF/hTa2xs3Io/EFV2aFyiFD98Xl2MfTnh2428aecILl82p8+FumqIHj90foz
CDmWcZnBLwfqGvPsY4C3I3BQUvgMF7I5vxnCjyvjujDj8KRFj2MZxmPP2u2eyV7N
WJ3VPoT4ncCoIV/faVeD1UNMy+aumCcSDw71RDA7BHGZzvhwHQ6GIgSTyWyy/4yO
fjm3K/rVOTZsnrXzVyQ6vooZ6CEW0qFEBMX+mv9ZGD3gR3+JXgt23KIKfmgXvr3E
Z8C7obDaIwN8lVOVyXDqNmxUCbfI1RjPIp99zBKBdej2cj6ncet1SOgFrIjuBqOb
HxExOA3+WeiEbmeuriwwzt7sYio3j9sMJ8J0RzT2FZrM9ExSoAosU0WdGmenVd0N
RMY5bpkN3nzqOWTOH/BuZe20XimODRs4Pkmybwt7B599J9zaWc9Q5vMMNnh4l96K
yx3OAZTarnkUhQeBen5/ngDHUjWWN5IqliSRMz4auIEYOsnBKBFtItrV2kYYHcCb
OPkfhEgff+fatJcYCrNThqhADhrPzZUNWiU3qGyI2c9mVrtgibjk1g7MGbq+0enQ
FNXRiLQQr4vpo3cDEmcwaPcf8DbxgwmD4LRjVZtb4ZObppU9jfbW2GF0RRFKLsdD
dEV6hhKTtgjGxbzsHrD+YX2c8XOvuQ70tnx1DMgCvdJUXmrbBTMO8qWokyE1nrbt
2xPHzSAQzyQFkfDJXVnMNtRKvgH2OgSyARC1ctosJwxm5wHuM61BgOzf9hW0TRoH
OzMMA4nTFn9UGl1qu1vg4taD8EuRPysK51hULfiB3MXeLm4rlOAFO41CWEhUscE+
QqSBKKSnRJH1L3SC2vtLtQ031h8f7fcLfYPJH8DLwHYGz6CGZ55o66eElw6o1jXa
nMJyJrmjgr69jZNpRmnxdk9nKDnD1jJld9tiCWMXXsOif80dOo3TlJaIDryZ1mlZ
M0P8Kiob1mALIHjf5UdjqGYduBwArk1SCoApeYwMXZGKeLfFsg273AXsoOtNSdtu
Y9IY3sLykNer3ayt+IUfEeVLjgFRN+uIEj4d/81afDfbY7GhBlegWtFCkRa5GhXm
jiha06J+lmprhmuKZ4sr9Z9K3L3l7KU5bJq4XROXIdL7VQ86tOE0aZiDkW5qaSks
xgTnQw7DYwpTaSK1iz1OZkgm3V00gkGOAMN+/SZE9nisxAHsv6x7wqDV81S90hiZ
3kEuWt2qq6tEJSIqWAbFkA2ho9m0LozQq63kzpBnis0aGHj4DAw1Dk1LZRNTFKlP
4dZh++gUryHNXOUjYgI9LHhjjj4JXnKB0pRl3lt0jYcZOxhUUrKHM0EpqqAnLkej
FqDf/gVsDZGwbCsg2oCp5NmVYvtDvxT8Mc8cyxwZkTw2o2YNMsLftiPPMzIRyW54
WPc5EH2jG4vqPNVuTS40xDdSRSTMxFqcw0I0i9w5QGuxHq0SraowwONkW44j6xB1
sAdGfe5wP9tTFZtdnSc6ELaIIV1sht0jyAL5MSdXdqf/OE/U0+uV0dHv73zEsVbg
dG2O7jag4F2WCDhWl4TLv4J+o9Gm8PI5JQs0njM3sunCkw10MzHMltTCCISpnTya
3UAfuckNm3QOIO5S1kZnS7z9nosuWLDUSvrQbKrFc/NA6SpqaihSzCV7L1ngwTPf
GTsvlM9VA3r6RvxMBNdr4kyfQVyyxURDyh9vSq7I+KJyYTVycgUI9s01G3JY36WS
N00GKm9ajs5y0pRj4SSNI3olk44OzhHG+K2PAlK8Ci9q6QrLv+o4ZaYYIL4BB3AN
NIbO4nN2J2EVWQkNkyew/cbh+u6frE8QQweyeEEewPfftT8ibALnrVHCSMhowQsB
3+Kcr7QYJWHs0CVTvmOzQD2LilK+FyfhDCk0DtNaZxNktlYS/Nyo6/7oQUGWulOS
mplQj8uuuFfBxWR2a9RSXcew1kXoUJMLgsHIraxtok2ONZjBazHLIY1IzM9mwMa7
XRCRffRHAFco6BLRZbzMO+1EM23nFtRNMvqibQ+fx9IOqC6GrflQUC1WSmbEVaeQ
zMpcdrTsdbscF2ZLmh7S5NKZ995BUvGfgUvqbgelCzLSAc18AhuS47WWENyIYRbB
fy52IL9g057D/FzlCieQsOVxCoNKmaAgPG/xXYu5dcs1/9Ag7LlZpAfz9g5+nPbF
jwQpzeASkKfKRUyJ4jMWfltA1McoPbwXfsECx6quhHYlMv6szugz9mDP+rH0MvdJ
Ugzeu/NdBPvTHP62JF+YJdbbdY9ghyWnxxn1b+M5SlZoZbqxU3fOvXZJCnpSH61b
/wUMwl4nlTS0L45Ncyqct2JCAJER7joVAzqUOZvidxa3OzdDoM3Vo+/Ssz1ssDuE
Sz29m+zMDKJPWoRuxauNv6YCKd1F+dn46Uw0LHZKvp4u6N/OnYgTnTse75PwuUk8
0CtPxj7VgEx1lzjpKP+YYpvruREB4rKOaS+9euX23cQO0lxHCdd+fB9cHE+MmF2u
5zDlrYjSnb1oAGvZIVrHEPkD7EQ/nSu57azqqapsn0rspr00Slsau0HNinq3Nzlc
0te3FDuIU0MqR0mfjVx8lmYTO1Pl0oGBQBO1+XHVIwONpjpeiagDhvhGJUFxvwnR
jjv4A/nbMDMBrWi7v/ECMWrAdzdBS28menJ7kmCg8NvhQcN7n/HjTsg5INEj0O51
VWUhMcxQYM6Vuv/oEvluxCFZXaWNanrfsxiSdTKhWcfXd5i1pfP/Jpfaed7FCPua
xgKVzBVVMoxjRnnKhneUnuvNtQDjLIp7th9wIwO6mz8fVjObTQNtNM//wmtFzfGD
gH/aO8RuCx5u7UIZO2E+R924qpXmgomEzQ0cGS5L3UmjxBtp6KMhcBTcZUwwWuaH
pjcJyG+BBKH/43WDCJBzYYRU6CvXocd/3aNyow++R9flCntb0AvLnV42EP7tCth1
Ashk8Dho+2HRkahJJO+MP3BF5GzbAKgZRIq4X7tLD3IBZASvdNM1YZ4mrx2E73/R
oim64yG+HNYCvH84+Lx8Vk2vdDdjGsNnj8s4da4Occt+GtPJ8PTcmt+LIIYRB+S/
oJ739WRUhs4EZ3eZ7CBEbvTWIopm1tCoGhWU6HLGdT9PvOxqVqxkMgH1UpOvE1aW
Kcy0wkoWnutUo7vdSzjIGtJB5viT4AjmIPqQqNUjxDGeqW3UyXyqlB5IVsEWj05y
snYWpqVz5MtrZyVmhzR8Ep48ztxQD/r7QcaP9JieVCPT8IeypV4jbidQZd6KFkJe
Mo3CD0FoM0bs2OjDhuTZhtGt+ADpPHMpoHBeaoVB5nm+wUuf59NDJb2OGEQVrvN7
OIpwJnMImOIqtV9Ip2oM9kW3R/3ZJnPuoBPoMFqEOK5m8oQG5BZ7iVAKnhjHHrtT
xjJThwa/uihtSG8QiyP+FlkgKqkyjL2ebOMXp3pEvSVtQrZgfFyyxK7wOiBmpHZ5
ayMeJbcOHAcpayjHNZXVjGfWhULQNSXKCm/k6ivKDLrYM6zewSGCl8Oz5fXIMPC5
pzt7+St5YJReq5SQtvDh3ijEo/sJboswmlEs/sbA+NOLAFppHR/rU91/dbZf6WLz
0nKZ10pxjI0Afpq4JtXHjE6GFd+hAL9ATX/bEh6GXFU7bP3HG11AsMnzrVPJvgIX
HXsfx7Ya74L2qalINie6Uo21fUCGfVxUna30/w6DxD/UFD+N2iDnXeGVgv5b5GiH
Oekaol1UTMWBZ4l/W10LgMCZqfMcT+YwZMues446rBjRvGHe3H9q4N6/YFNAY2Vv
TogOKRVkJPtcRNSGmWLSaWrtpKEHC1MSRzBu1nf9TE+MgCYwcCldLqbYc9UjAF/c
V/5vAJK3cvLUFsh4a8aB66vER/ADYg6VQVJOYHu0w/pF96wAM0w42SqDchCc6Zc6
ctTTLp2faApbm7CDP9BJT97mEzsgO5dcjoGSrcfZeKKmlbetF//CetRParRbm+az
JaWJ39x1JohRd7tTZTc/7ZBoNOOiLmyZd2M8jJz4rayTvNg1MagFb3CtC778iGxw
86tCRZRiAQXViAjNz80JmJHUu0cKBlpO7xNY7ftHg/nchKDTs2194bOoO5MIT6KO
p1e6onUWhVTrjqiJv0aHjEjYPwsOzJJJoGAsE+uV8WO7776Zd5MMvTEnRKQ/NPzj
WRsn9vwaAUQZViNPnzK5OXI8l8AhuCL3WF8kQxXzDLUa3+OuL3Q7sp/dNd1wTAah
gF3AWOdLbGcAjky0p/u9PdAsxUGYy4n506jnrl4NRCh9C4j5SiGMs+n9tZCPQPqr
1w6Re9oceCDu1SfnN380OvZsWTQ+UUPxwE3QxHBiYhy9braU/cv27m9asjTPmFff
5slcxDDaZeREKSvzAHSMpBfukMroWKYxKEKICmnYKtLo2T/MN4Wfaut+Ws65S/8U
anIZ/X2EWR7oeD544fYlnEviZSVOvybyNNEoWXwnb5K0IOcHKWGAhttqW6ZAEJXL
IqvqFOb5Vj+Gr66kQbl9r/PesTiFP8Sw1f9Cd5N9FizRjlExZKXJFckDgLyI6b7r
HqH5q6XvXlZKFzmSwyE830PNM8Rg0uQSAyfK2BMUI9tOEFgdX878S+0QKgUbppkj
g72Wrsq4lyCDdvnWonRqdg5KF5pZgCmNRWf2ZTnz0WgvG5IQfBiAHu11qOLpqkVs
fNbRqYnzI8Hu6vI9t/Rwc+sfuGUb8i4D0qYd2EdCp3KLkgk5gtReYZes70knQ4Nv
3XBbLAnKWDboXTulo88Vn9u7h9ItGn33DU0owkgVY5y++TJjaqH2qIWH2zlWH3cw
o7qVar1pB+fFstlfCpjLJcWtJtp4UemTbG7k1ckDB5hRgGzq8OWDa4siThoHukSc
NWxtJRanDJKcfMCym78p8FiUiawx/sQVedQcxmcmW0t7Es54p1xdzdVysMDVrBmI
aZPL5aJH0z2tQJOZ5SoRMjDr43JI9jgBSMCgzjbqkWKq2ZQF3sajcgUNEOyKF0A4
A91wxYfj5MEqYPkwsyoRAnypmlqBjcCCgaFl2k1a/rgb7brJW046yHI2lCwNuLvG
rhFd36LVeSjIXkIhHL6YS219pOY1ncM+XhFFzq2Cv1Qzsnz7azKyWcv85X6UqvAA
i7RPPrVzD4g36+lhCMZfhsJ1NHMskKoIJBq1IbfrQWuLgwoQ6TFJhwANE0kYAYsW
td9ATWLisNGmVJCR7mSJA1g2fGkq5JvkF47qdHxVkVmo5HW9fJ6B8dXfMyLniyJ5
Zv5jZdmEIav6CUHkHzh4CYcI3TCwQ0aEy8rWl5MTMESbDTbjZX5Z2eaRn56gvZdV
kiCo2C9DuEl5NVr3brOY5M6g5vOrBDyVWPo0w1YxQQGvgq05M4rBpl/zPHk6nDgY
wRtrPONSaDQXhS1/jxCxt9T0Wdv32pIlWAGs6NPgVicQ8Hpb7Vgvj3oWjiJX+pRJ
zq34DvZAJg1hIns+q9K+K0KDqia329fexL4g3Qn4d507uUlG7k5rrN1U/kvu82VK
j78BOzL1KabZWiJIAImfqR7R9wAcIgPMSrHmc/35PTwhDD4uy96TrMc7j+WwGrZW
W7Zq7e1fYizSdusNSTecXC6uLtdeJBHZ5mVSYzT/pfOikK1HBn4yfcwrYsdKfMj9
6NUfOrojmE5PYTZsUkBD59NGWoCE+AZYzXcEnvWPWTrXAyAKw17Aj7pX+yi3jrFh
84o09UqFVXttPGN6Kemyry0CVFPEZ988Cq8vWL51v9Cva95r15KIP+bvJI6Nd8s1
C4YXWlYv443H271c0hohQ02TCRs90sv/bJ+MhF1SR703x8FnR7zM5Qqu/zitK7I6
Uko+JfZ4a7rGKc0fu28YYX0gYBmtXlteDrVTW5g3k0ccQCEQWN5TIAsLeh6WY0kI
HNL7uF7MTrOf/zbh82RpbuxckqOwRwTKIYAsImCrJgOOTuqXqZwo7gVFjF5xtCLG
5InjmSczhqu07vn2hZloOQeMNv35LXCf5fY9G1bq23ww5sLvNse+0Jd+g7RcNtF0
cv3h9pF8dTEQHhs3+B6UfGdwtJ133/wnhA9lrPpa0zqS8IpQhwLNoCfAvPs3gh8s
oMBaB89wrm21A2+wOMX67DCSv7SJdtd+l7cRL5BGpncttRoj1csCc2HevbraYDzu
qlYH8Z5z4vs42lXRcfsi+OkaEFEI29rLn/EBPHoo+avmEuw5KFotB2oWOfYmene7
RZPqZyroqKhYxjchN+08gDiDrb/TkDdlet3OHlqBh01mF4v6YbgIKWOImuO9HUX1
FikltSvLR+qP2yZucfmCDEc6Drdn5AnIMOV7tGScwTndpZ6Hy/kMYcfKpmhQiuaE
ilyC6Q6nW+Jrzga/q08oHdzI9JGv/3lwk5fy5ocLl6HGrfGIeeX772zzzSWS/+O6
badCClDZTuppl4tN3jwQK2J1b9XODZhxzo0GbuOlFcuoYbiBTYblOr5sJDYoXH5k
J2gk1V8VkGCeapYBXo7r6WxCJNDxIYqUYkGFYqfzj5yBG5Z70OqRzT85lyx+Zt8L
iflrx0Uc7sm5FY3xmkpUnMQDVz1UJe+SKJjW+wqWUFIpmlqgd9kfzAPnIEqmuY25
h5vss1u1k93+5DM+EYUqhpUGVDbaY8+AYafLbLSf+dlA3OxPGLx16qvc7Sm3H9bG
amca9KoJE8P78iYXjk8rjuSwxj3afmQhz/ZveW6PgOYk5+YaXc9E6KknfPMRQNp7
iDxmAdam4IokNMgYJxo96wU5Nicy0vdNBeHsHh5NwA6TFJdmvnJeiZxcVdwpRLGN
3ST4saNnrk95BMUWDmnWwzV9nwkxq0J9uwSqsjWzpXfbUBqhIreklO2kdStSUOGa
pSDyqYjzpuQZzk3R9y8PfEkiGgt2lEvXcyHzMCMDB4pdabft1EhrXIwmZCw2q4G3
c2WZqhGeVagD3H1F+p7UZrLZsNTEmJk/CbxKOmysoA4beAz3v3xynvN0O7A/t6Ks
Jtz9vudROySZEHx0q0+keQJ5EiilTI+fLgF6xeoAhBFfXl8o3hEPHgA/RxoVqH1o
/EFlHVPzwG4VWtozIK+lhzXTIUsW8Hmy8cxV2rgqEyqBY6uqHMIgrAv950b9Czqx
ADFRu5zB6dr17hR32NQDsGgl9lEHzy/GyLiZi4YnnC/dSid6ww29fghn9HlqXuaq
uTJJ7eFmi5Nvaj0oebyry81s132siM4pZH4RUXeMLg0StyU+xYqOdUKixdRguVbl
XIHotw6UCt+M8odf8I81q+3KHreB5UkhV/I/8H52151rMEeo6qdNpgJHy7HobVP8
YFn17cThC3KLcgU504g7aDNC12qSq9fQ+o3AMEGK3K+Et9TEL2b16pOEYaSawl5a
zbSMonoQtnyOs2sjduMfzc7nGKP3N2m3oIp2G9skUYrpPG7U0oLCIn6kneN3A55Q
/oFBys0RUaaxwtzbWQQuMSNOUWadBhztpH1DvbjMSQdI0ZZm4B7EKCtWShQ2oy5r
t0bbc/a3lNTGaIUIjnd7X4xKwR/lBef/QGzgLwN6E5fK9PbkGeVKL7q+MtMVgdt/
jAlnhdir8eqV3c7oeId6qMBf1kAC7QKhVEr1FHNiqLshBsUFdQF9uS/UEEKdKPDz
ZNnTX/dhPfmII13h+1xvxERkPbZy23Ls4i53f0jF6QduRMOOXfLcqtTeNFh5SVFF
lUb+e6Gxmjl5k4vK6BEhi8fO/9xcT1jn2CkyKvhFTCKxKFOjYbALPqlb8VJKgjx1
V2na/my6GDxjdHPUjTUMkMKZpUlpNz2F+kzkQT/KalcKXG+PYnbAQNylM6aksM6p
/xZ/ZY7rL8A3gHoogYxY4P7AZxVGESvjxNUlhlk2y+RGHAynLWJQdUyqmjHeY4FF
qY6Wl59bp18iuAs+Q0ABtX2h0y0vzrZ7uHdJTWHoTo3LJRxycIB7f7UNEqjPzjmw
03Sol+OW/BTIp41enxtDahg7IDei7FdD8C/zWp9CYsoiUWy3wxUQNqoRX2/ZiFBq
Kzt6cwSgDtYe9dL3xxcAve51nqz17mmG2JvdgejPOnn6wOqP6VbMM5b1j3V88xtT
9LOJOskEVMjGtUtdvZgDEcA7B1T5cosXlIJFed+CwqcPZ2FNYh1cLBxan6UY14lf
A6DgjADu56WzxRKJsmKrd7lkJFK8XFFxGXGu2HEh9sbgKFdPn5F89ITvGEaHCHz0
RiQ7+gZTOhq6YBSRMsLHn6H6YVn1iVqNAcBV3092NOMXNCrO/BOeUBAX9M3iZmAe
1sdzVGvoknyr0/OAuXCWmv1pRxRhY06UqH17IU/3qB0Gs8HAGxNbz7YyggGt1X5g
CYykDd9VQnVghKI+XhPlidNO6Yusk5m2/i4cXLb3CJKxDZ51EBZnzN7LEfqiFJpD
xWsjdP45dD6CBv7kcjS6iIZX3pQNRW3mhKCyXGyQkA42VcgP0nMOUOYKzlCqbCLx
Rx7tMklenE8rbfkqFyheZ0zcvpEAy11Cz4xFLpY/2pA+bqaHnxLOFUpeKgqofhDR
Awbzd8n5DhakEC+e4nSwxpYH/vQZT7CBdhGkyXbH93Kao/A5q5CcHLMUsQe16ciG
TzdWp09YET0Zndmu8BzhKlYLFC7LCbegFH+tc7Tsnd/KIt+ZX1a+Ut8iP1U7dEOJ
OHtA7pQuCFUq2244oi9aVuDp48FDa8xyIoEBjGKIQlTQLydTACxYxLU6gpx+v3o/
itFolOdDNgerf70uMPD9qIxLcz5z7ToERIf54IQbu7zaXJyju/RRoAt89dMIXZE3
EmbC3j9gn2xsFTaEovcrXKqcEZa2oJSjfWDW6Ie/I048x1A+KGVFT8Qp1m6dKIRT
ZJX3pmiLavjAdIQYU4KkrB18WZuLPGYnGy9/v9DgOQ2fvHTI5jg0y1Vmp6K501F8
D/T4N1vErsAe91a5/QiTtsWoLO60Uju5pnc2RyMSUOS9IohMWxVqwLpAFsMisZnF
P3wbvMxDkQAMc7JtDCYSApd685pvtFQXe/XT9lZxvlsNZXC2jXwd+XGcKcU52Epo
fnJFeZnVCflNbz4WFvB9owb/jKEtNHqKvJgd+UH7nRNWETSfoVCgDPFvBw+SZ9er
r7/sRbhng84QDJ3HAx0bZPkJSrYaoHlUL6hFQ3wYUpxPA6fTFfiPSsXroJsOwp8h
hR0QiyqK+YSDlHFhTWZlMdrR5o5L1/ZqkonbJQl4Paw/xraOA61G3aN4u19TfunI
EzWsTgXyzmMZGuAo3QM39XN2HbrzPYMuZAOBcvYmveQmr150mmdP9IRnSOEkIpkt
Iwi/kuLTrhW0+uc2NLksYDTIL8pUDKFLGaJN3uN82G7XRGLy9nPP1LQ3cHq9ugD6
yGUEIeMetYMmX6Esb9D3/p4mRPZM6AncWuxVF8c/mRUluWu15tSDXEat1v8PaxBl
ByPMAiVXutcQVscO5Lg63MyZDb5COFBqa8sVll7PT2Kk5IsS2nND6b/m97uAJ39u
nS7chxDlQuUyH+jzHGEXtw+3NMuCZ1zLObI/hGKEiaFVAwfoPjw3W7fm0dNK4YMI
OaThfPukz/CTnU5tu+JnTSKK9X8LQ4flir2YRimabRyJM0/nNxYgtv9sbgaCpxpE
8K7I20rnQ+QwUm2JCHTLYJISi9pilgiXbr+QY7vcFg9JvqZq+Lq3zLu6g6FUW7SL
rcacLLcDXxAtlahwW28ujMktblRX6Dt/+gW58nMoOmNR8cQ3QzRqPPckAm807rBJ
Zf3SDVMIQtzuQ9JdBUh5hB/BCj7wPEIMkH8qxiHYNVJb4jz2Qe87fejR4oENhp02
83qD+vsAhtgbkGM3g+KBz40sT4TZvTzyE5pLHr1UG4m0todDo+wGIs0dn3iJdYuT
MlnzshYp6QTHs/yCck8N+RR+x0+Y+xRuU4N/C/MyRUGHPL4YEUjAeNj3IvpuUx4j
LfeizgvjDDE7MEFLWHiwtqJ3GwlvtiFnETaGsbP0HFaDmWBmGPadW2av+4FUqYdN
YudTuooPO94cv0auZ1aUGDVTFvgqswTldm0osUJZHubYnb7aLpDbx317WrDkcK+7
MBq4kNOyc5tRbwHb4KxqvbkYpz9/8YmZGE0EJUf+pUP/8BX54i9Fp7cTj+ZULCY6
J4ED2OJ7XJ7EzgquvUFfvULE1yuJINlTbmhNBUNd274tAZaS5cxCHzHrF1xXQnhr
JJhvcww9zEcdxGA+qXSpMCY/yITIWjKhLQBc+7EHlNVMxrPGO36TCc9aZr9mhaOi
dzrlJ7O89oaUQSd4bCyejFvZgnSDAHy7v+TkuPfw3SzLKTZAeC0qTTAZdodQKv7o
ZqLO4WnGsRK2I5h0XByUYnnpLBPbGU9CcieeJ7NBB9W0EblPrns4f3l31bZ8EwTd
Zl4kBJMhhd/a5U//MXbe2fHWgh4FlVctCcuKdMXHLTWrO692G8KzhjpHmo0kE/+3
YwX1PQ0LUnEO3F+eHmpszlzRjAZvqtHNadOM4kcx28+ByGNxOQRMy5bG/9O600H7
YRfkUU5IOrui0/bEc3qtpQGodrLN6ZljsjaaFB056R6vbYpxWx7lnDxbsXsSp7Un
EIMrLf5g0IPitBzOUh8kR33P4Wn8LK+GJA1UWVEpOKK13OIPbIbvu+idwUkBXRtP
KTpwRlYg9e/Jkbw/Zmu2h+/IPdCK1IQIokE7ZqW3xrOhnf0isQGK8AfrQogzhtDb
dDW9Ef4PGVVnGuiLtcrSt6n6hGCftjjJ3qiQ4nN7VN2E+ZxiqdBq1MWGz2O+cZnE
gUy4if5rVR0JZGHd78yVa68Qh3JRBRvjIsc27R6XujRwIMhjN/hVvSiTzceOaBNT
KE/gk1RG0jrCkCi58m5REzHmH9bKLA5GSz5keg6aMdF7ryIxhfmBWwCQqpzLe1Ev
SLVk5kX9BpByjI3vynUEum2+uXh07cj19qxf9FYNDL4o3CpyNSVgXierlD6UYE3Z
IPpHjuIL7ioYlHhT8FOK0axDx7Wmt/LSjQNu6ZB13ZbwQhgbhaXK+hFviuiD7GqU
JddCFu5i4cU6AdyEwK6mQeuulWHwoWuZ3k4A2DjjgMbjy0FbLPA+Hok64VgWV+0O
tx0q+GMtCnS9GClHIWJ9E32nRzowCuFMEpBmw8PpgA9LsCrXIxOQeYRFKcxln8w4
syI70lOb2j97pYTUd7JXUh0G61RAazvAuVUjqbBmLRiJNa8Q3o1D109oRCDzyHut
++458YVoKO3v4Iy/68U5uAFl998EO8Zy2zT4qelmioG0PeBKdo1/SujCilphLpjb
LB5HmQm/N66R4SRVo+IB0oqeljsPZGLcfbEwvKWXDS+4TmdeIBJDlpR/Akg4P9Qp
r5089JbcAKdb8fBTOdmBTzLp+Xbx89JzG8TwrRr/6dwMZF+H87Xo6DYyZULUL6RA
3l5rDsy14Vr0W4+QzXq71n0bTU6uLYIp8j9lor0WNSFHI/izJSP0CO9WklsO4BAw
WulwAn/+y8F5QH3G17vE75Wz4pPgmtfZLCao41UoQrsLkpR4vm63gYurmppW8xbq
cKcZjPkgE5VC2AQgrzXI1by7KZGYYQVt+TMVqeMOK2gIWa3+tpkXtBGUMhqguW4F
h2WxHkCi/DBhyQdx4J/Mdru73xNqvhjfXmpAPZ2v2at15NIWF2NW2SMuJTJ8cytW
cbZPzbtQUAHII7GhCbV6PGrmTzeXw3ydx/XkZqyh172wlfyolv5xDtLgI+QzONiK
jroTwqF3eF0yLyJbybYt+A0jZIBEClIcRVGLefwYB4WZrTMXkmPtJ9sp3QNVTx/y
3+JhvjdBBvQf6X+l7p2aK5EGsEPoQMcFzyTPa3u+CbzoB+qfChT/VME6bOhfccZD
MlTxm2iBiaWHv3PTvsDfmKDIxcN0ckMao9Vwcv+HraKVkGCzx1ZyIYdLcEeMNQ4G
4EpmfwSHZvAwXANpU4ESqXNmQU408ZtrNOkBKb2N+MVyvIstc4EaMxZ3FbxDZAuw
v4eOTzYpFFjUGwGAFfosRSWcOBLKp36pQTgZ/9ySEbqUsiKLm5WRo5ts9+ty99iV
kcBlYQnVpRznB2/5veH54W8aqvbGM0vUJc+YHOV0bg8OZm7azBiPgTa8K07perHx
4e1uNj6eDVI2OVuB2SpauoGr/V7Gfgg+VzwZNXEJ6Nl4U+e3+uRzJF60f+TFBTP/
WHo5DrQYl5TWY8Zcl14VvOXQoZDisdrqFRCmTXen603AFLJDlUJQ5MDypbVkkRxf
NWi+CMpI8CrntvWNXYbsrC41pXGhLHI5G9I7VjcG9YLNDNSM4s9fZZywuhtRlVqd
4CDqVq+xQo5uCCd9SHrFUvp1sN+1WhMo8Rzdo91shT443u4Xt4hSxW/DeKNdeQah
9M1YZ6Qrv9kLrBWTFfkLIa7chq7Fcoj1XeO+Y4UQUMt6e5kIKFIOCAmuT0fbUzMb
yJe/BszMdLaH6TJO3gh00v/ddH0QFRzDn3UdwW04vqEjXdv6kEgz7kWQkNvuZps+
4pTJmS0+jRnbCaVxeF1FIJzsFsIjBxtQYXnsoTntvz2QPTbi7ciflfEUdKDjwDz+
gdZglT2/VzW1SGyDW1Pi1qHtZMs1KDn5wOLATN9bENzUYQ9MLw8aiOaXFQUKnCrS
mt1Yh7ZcLzp8Z7nSBGP0z8K/GmL9fNeFkocN29LbNmbMh7INZWRqcZc1VjLo5ntJ
hweGMTw5rXimpfBmP5UIorTsGC4RR7Z1nwmss+YoeKvDyTLEMGqTWksLGl3qM8Ri
qz3gerXPSWfvwHcCiwhkzumz1Qx8hiecaHIDewZNIb6K00YbvBCwRGMN0HgZBwNb
Z6KGkwr23D6EmgnNV3xJUDXXfPrujO1AnyFAF5saLD0u2TwWp5ZQD3fZVmKaKcHd
9Uz8ZDUdIpP/bfdFEDUwpdN/5yPCWMH0IJssTsM9byUhJKuGs+ow2/TcXGD/4S4l
aJ6zITmDxBLo5RE9Kc4jfQiF2SsdwaXcA3tBvRx0abCPcSEsbMiWpOWf847uAixt
7IV+gtdGUdNB9+kiaqDB6t8LfVK/67IPxei9jaGp5YHdnssCXt125s4C/gsVtOTB
TwUAZU1ZCwbOIyJoqFD/4PrEsJaCG5WkF3Cz1QV0zCJXnhSMQKYM12zRnaw4T4V5
qeJydhViBln7S5egcEXDCHB7iudh8JDYlne2R5eXJgtl23QalpojH5kIK8+YzcLA
AuDBsgN+RTtxLlhh4c5U6B/DfP0UcunzUcYAv7u8xx4TRgyWVCvU2JbWQ2wlMEWF
jrHeqwy8EbAfgqZiH17wlCF+WLlELhH+UpMkNDdaf6c2d+7lHEFpmr6Omjrj6wEL
tajgI2lOS501jScyvXQ97vTjTr0TfaW/ePcKS//so3iQyVy2oniwAKMENAthKLJ6
XHaFFSKtr5qUhc8U8xzqcOgii29i3iuvF/DincxPFXz+mVit10AC0bu/lE3gvwVm
0mi2BjRagO7aKcbxndnwO8ePwUyALmJ+siqtwTA2fgIjbUirABqBLS+i9R1bVVce
R11CN0wkMMo4EBAyZuPwNhALgjbP5QB71PYW7kmMP6EA+7t8xPM8yg1W4i8V9qko
1U7XneM/yjIcwpp3GHh4veC5NAb1pMwJ4Z4hkwWMa8caijrq1mYXe9ZggzWo70xk
w592NDOI5zzILpW1pw5uP4E9FHQgMb8l9RqX23/fXPjyPhoAeo/LSQCEg51TuYec
dTYfosSqFCAB27Pb8bZjcjyE2HurHumOP1uymJA3JJOQA6h9tqHJ5dqO2u8V2FLC
dRyU7Iltf8h4SjtUgII++g/2Wd4jEKVjOVp1b4xbAihuyEoUx1eRtw5jb0lFZU/8
PCOC5VvP7jUzRCpsYRdjOai64CyKbujL/Lr1URVntkEG20rQIaINRi3j3CZsgtVw
8LZCzq7xcIMk+AhVPAM08orvE9Jhz3PWmZBquf6alSP3B+RAIpZQRnbpm0EW37Py
TYTD8UZrY9i8wGyF1gFtMY5kPnWhAN9zRikc3EXDsed0aAB2bOWFm8cjn5UMIIqq
/aODkIdKF3eI8jkM9pW+EkcWISZgjLLo1m2nL2G93kC+c/KteKsYkE2v2nJJIheM
kgmM6XEWeUAK/RWmAoY8GMVDt0GVp6Sgia5O6l5wOYVOTlo4igpKpUipWfTxc4ma
4Mmzodmxjrs5/sX4i7ER6Q5IebhMSS/AI7MCp9fNSYM3rSX4wo5+5xaUZC9sV/o8
K5FLIZF3v6aoBAoBAKefecviquYFuJGJIuXrl+8DH98We0GjTBBqc5WPpJzSWkeX
YflQY0qRLDKBp2GHhn40ET1pbANM0u5dPpssk5Z9+xofeyzGKCr/WPbShJIxo7s+
W0YP/xm8OwFL3GjgzxXC9ikywxpUobRRovdIL0/0V9PCPJmWzwC6PYFBiidP9uJB
C9yqG0HRT/vMa1l+z5ycn1v+xWsQfGWCcHfD0CVNC1jEDsJmWPkOMOy8n7lCr3MR
Q+CE+cRjeH4GvX5DxP0L4y6uxQlACqnPX++DiLqaQp4O8sI3iV2WcCNxp9CxHL4h
SjMDoip4O0TSCBZGZC5nL+is+e9hDBfdhZ7EcGzcD/yib4kGTB5f2aaBm/0as4Yz
DRbERFDHJg4FME3bS7NBxzaS2HxbPrNWwR4sMt64XkkuMZ2trFr+vNHk4NUCvjSb
uFtptKOVeDwVLBKv0tvngpTPKMvM0iCg2CKe7sGsA1xw4pZRqklVX8+rFLmn54VQ
nWG8pxNiJaNUONAJL39VRz5XvNT9g/pCzdcf44YJIQkJl5xHYfhAV1oNZvVd5qHO
K+l/8DPKCEqglYqEu6trehHJTk8RwOACKA1pNa72BP+ITFtXxgw6jmtvMIA9Idws
M4WZNYgB3iUU0hPjqdKXlUzMaBAHaNxZv5ccSiUHT7gr3McSrNmoIcpkDjGIZkE/
hd6ayumYnKoppj4sfuMH9mGKM6MWG5z0GU1MQ7YQ3D3Ep2Wk1DG5L+QQJAlW0fcm
3q6FLvMB3+Zm4IFgsr1y4IkizjtxX1bw8CN1ubYxlW1qXOdz44/t3uwsnEkGeVjg
vQbJ7X/mN20CHTK0lxYUkNw6/YwhY9GUy2ZrhNkN3eXpliHy1tAJcc2ANSZm9V7B
BY5um43dQRvy5dpOHf85QWo993FosdKxWZWJTdPzWng9Zwiq5l8YuK6N4rzvXv1y
Cbnm6LMvIJ5KG2CcJoHWFJqdtalt2/P762+NPnzg/yHZMTrbvTRHgNa6WwXg6GCQ
ZTDEovv9mKmSdioCHq1k4c2GpggShqCa2uI/a8ko9LbkgK7LtbcVn/WJdmCn14As
sNQev5XoF+ABJAWRZDWrB6sak81T1ZjjHAWjjvdqu0yt0o21oUCg0O4ZXNgMC2Bo
vfl1Q/YU/ENajgGvpQiIVfVE2t6goDFPNEuvcD8gBV5S6tbquqSqNsqbp3YZKN0I
LfKvc5Ie61/peGSlTGdIAda02EyhhKSZ+Zme/8gaJeInWF80l0k3vzwxJesabB1w
B6lHOWV6IjIFJeInGyuVlL7NwZ9jNW7Qol50GCH1RTnz+UOjiGVr4YQ1ASjmebm9
bGymOjRdbq+56VIrFKsvcVfTWDz1laiZ4weVdb2KyX/fI3Ai5w8VLTEec19A2aBa
q0RreKXJdSdYxwn+0rZL+AYDi9LKGSmLbuhr3J07flHb6oGVnXsVxXwLm3Y5kQrH
z2KC0dpzi0p3Izw3S7bmZDHrddYFouAXS22OmM6sx4AmsHUxmlH3El2gk5vA65pT
5Nw9C6edImYmhIAoKw4/8qbW6jT4qa9Jg3NmZklaGbYobnc3+Rc2+DnN4XIbZYvk
/z6DbRWauyHKcBYt+0eXGTbvc+ARL7G+vg3p50fI/OQ1iyoDkF++sFugJmNyrlLn
/dHYd2IRvvKLDle9JjCspMUj5qpP4idNImHvP/cnas0BgOgBCNln/SqZcnVY6La8
elX05GA1JDwifc1XV1gdwaZ85wP9nPQfry5a0odMx6jYryZU/zl5ShS0YciUg7gs
5t0UV+lPgkpDHAoN3v8jLJqhtORyF92SM8ZqJulIgZousgGa/Rf2/fAa54aHH3Qk
SynYM0/s1gpqJbCjbgeKgHsoh0xr4TOUYZ9zPEv8VKM+OZWRHqOazlu8d84WqpQf
N6g8IAXayMe3YiqkCmTbFjZIKxDZvApFsQhUzpn1UcHPIFx6xRDmqBle1wsFMj2p
LxmqmKKMYb17DV/TUOBCV6mtlsU3ozWwZ0gswS2MIVqiNdJOUstjXicK7pRwA6lF
mrXP5sVZh6M3X8AGJDEYFyM4dWPCv/N9ylBB/5b1R2k9PqR493CEOf4meDKOfxdO
xsENu6e183OfNe2Cm4abl0SrkL+SRTy2OW9x7g7MObKz7Y6KNi3MuDvmO5Txze+2
suzxYKSewYJiylFHNhmdCxamgfLAm1WQ3dBotVUbHVA3acNm9zw5O1O21aeS1kWr
ezCMe74gR6kG2RXu6iH+muPG8/G53wyS8JG1Cg74eiXyby7ao6Gtd2AfTVPbJs9k
WikMPb+i3+xamtYHmZtj5wT82V7D7KkJGJBut+Wvq+X+8VCNLSCbT7wbhwO/lXDC
+qc1+FHmzB12teZODXR9n0cQ6FMYJcUu4tU+gTxscQP4P7NcJGV+Xe6BbiqoIEy0
ciopY1JumJ/tC6vXB4SIWJoAc969t0NNPhEW65ejaZ9uPTGr36wz+7U/GyoXyz+e
CqTT1+sRnQN4jJVN8AtsMZTMdn7MwWtjtehDmTeqfTEZMrz2j1YIf1hV79/OWgdx
JyajZZNmFv4DeWUDo0qrTk/lcknSUfawWGuHKu6SfcvJNVLFIYK+0YF/Z5uFkrKO
oLd7d9unAkYW1oI11A1Sv845R5qVpCtrnQT4phBcbjCiI7oSa5dzQJAhK59uw9yz
ZF1ACmQYaLoNtTbJumlWtVd95+0qwVtJmJ7AGzKDaJ+SErFkSGwA1Q1J8G08hsiX
et9RDJdUGHZSIsVLmfNkKp9W8qU9yoUa1wvc3vVqoLUIiUUJoojnlgGE3i0iXlcn
y1wDomeGqAXwPhvWGgAC7rWO3/BgnIrbZghq0nLa8wxmcBg6o/n2FLN7E1sS+s+z
zNGwybuPIuSrG7hmp4xA3959JJ64AUbTjrbcfV4uXYGF9tc9TbWKfI3w1VINUMFf
xBQfylGsE1EMTvj3RpDkvjIWz9a2E3SXT74tnQCvmP9Km//uJEKArwNsidjYIQ96
QCT04ohE+pCxL0oeGJRAowApCAL+1EifjDHZ/9XgEauwdDv2zbjRoqxM6ej4fAWk
Cch21jQ0JalWMjhPIqnZQHobn/CbsM0NjN8Z7WWGSdV15XKkpJVG063BRgpW9OQo
+t10gGBIxRSEqLM3k4k6SdpgaFLWwUhU+zLk9N200cjYtk81Zkleu0jBbws2hBwN
6g37wCRuBizH2sJlkcm+DloZycYC4Sym/+Fsqg6Y+tXb3w3+kWfqpa5AIU5cFw8V
md2buegXrHp1w4sobBi1KjyNZf0n9qBn/2zVw9twZe1NFMfwwDJN5WrUSFrZNjM3
UdlALzgwQUd/LR1hg7yfdDxIA7Sx9NQRxUTIWjv6dRSPDbN9xDkBxRlVnnBe/4WB
mq6kOuIRhCLS6UnwpNRFEbhYLJQVDnzwGZTsWkYw/RiVUj9rdADBbVUMbDzGJr5I
FrtXhz8JOfcIQUgAb4XcqWT5dlBMZOpuLfIbCR9y6X1n9WvHTTZMpb8x9KTxxegH
t1rBNzFMj/DFH7HnFauZ4kOD0ufgnZ5n9NHH+ztH3RvhgC2Kj386SMYW3IUBSnmi
m7EqNjWuEEWlT/6nNkwRJi9gKC6SUz8qboymDIwTV2qkrbJk1wn3UkHs7r9h9T58
gW9SqSHZbWoS6EWXDRrVRbyPDDeG0UU5MX2xCpJFpfK8rEXzqFL/o5/FE5mpq7uI
C6y35pUrcN8FlQHB2pFrZoIW4vKuaCH0r+Ru2l4Oixkz4UbjerTIhgm3AT/MYi2R
S3lumVVRgveVjsGu4wqyvcejPytGyqoxpCjKrRXKTWKh6NRVfY/zdtoN5/M0loID
M8KwskS5LLI12I3h0mgAXfQk+T58beEdkfQ/3CzlNq2/zWiBZ3lr5ee2t3HMCPgq
tPVB5rm+8KD72U5X5YbN303Pv4G3uH20hOKBPOZMJdgC62DU31bEesIyn9nVzVSy
VYH1OlcSJthGaiOkO3PbWgREENmFZwfmNlpJFiEx+NMXbLXXCLDH1sUEpt/69O8B
VUjcj79vD2Eoh9mRIFV40T3cRGSakFij6imj/74EQQU7T4xG8dXpGrWz6G826Eij
oylHcibEJIw5Pp6CK20iu9hWoTsR2NMplHWOBQnINCb1m3GECqfckJIgWTiLlP9+
oyZE+bALZwHHt444ikgElqy8HxJB5Yb6tuGHAXGKskY6Sjb552MFV8ccQbLPdmFe
sGFSlUN7CMONYVbLLXEV5SZWL5TQZDxoAafuOy6oQJRxMSkd/Cgh+zfVLwZOmGsZ
PLphmbxpW7JAkl1VweGFWyY/pUAmW4njMdMjWdxrcZSJwhq3L0uaiA2dSGkEZPts
5Hh/OBhWbgoPds+ywX4P77fqrAcKSOGBBCV4UsXQpt6EhUsef+2VVF3Ay3ClKybG
KXvj8xGMd2BsSnSBrz06p0kXRJVLHGVXiilLoGoXL9PuhFNsPzDREewYn2yswt8q
TyBNcit+2+5NfxIrbEQVfloFi4u9L7WTbxxTGETFLs8EkaamZscZld+OdcwMcWMx
r7CtygaeMsyXTLQzUQ3FVpEq2I3bGaJccz21cjM6RXHquAcDaPhIzgy8ps58cP6g
tVOvEbaRj/vZE8lf+p9qtM5v94l/chWKQV5rRwIqcf+txWkfnHC6m94ZpHFreDMF
esoZmQOguW0i597FzCv7L73A3JXf+5URdlr6BaaIqu1ra6KkTKF2KWJrYVhOAeqO
1k4MMT1pMrbKU0jEz79wSnw64NWkaoYoska17tI/DdQFuf4SbwXeaD8DvGFDijzZ
88AlX4L7nvRuoqZXmXcmiXklrwNYIDcVUWZ+VeyH9ONPUpjDdcpD0PR4WsFfnwJV
+2G/aPybRo786dfjiyFcxtKaYRX3AC1Nrhhhqx8kz/VuzYGhPTH809kjc6b1C2Y7
pac+fCTa78cbLm11mUweyo5uy8j+FK2EC2CgV6By0aX+CAfU7b3xPz73JqKgMPr5
nvTBAkL2TbiOt+4kWOQ8e1LFLih8eE0B/ZpsbeRO12Ayx/2QlFhC26Fxsvly6XC5
4Ikz5peZMFZoyb395AsRhxGxSFi2vfiY8YFEyCKU6ebfpVCRHMIpLS2hHKRkNtLV
TmIxHUC4/2JapjyXZ8LSoDWZejf6VzDEptONW8YFiqtELsMqbrOaWjbhQQCl0Hh9
rcpgFmgpNw+RkxXNRPUOBcAMt+inQllxnJfVDuXFxjcpOt9W3AohUK+c0b0LwTuB
F2VSD9jrwPZKC9Rr9KvBQn/uaF4Ajeb+ARx0NXEyRk78fpx+G1xzFte2PP9IKLQ+
VEl8fXgOqKfbMIlFQ/ylT1T4Ql7Qnj9QRmCgQ2M6rKUX+unNvCA5vgNAz6BSp/ac
ajc/WbIW5kfxT+u9+tZTGFDfRkv9phkiCSEycbx9mqxVUU3qaW4L9TWRCeUWJBOx
c0sZ/9393o0v5mRaScdvpUJWvDF4fVR4dl/Gp77y4yLLE863kBWH8YYsum5lyFGd
pZUCV53qHaoNg8mmeQdv7ANmL2sHUZw0lOY8AnVS1O6h+MA2OJtLUER3c//uFd1H
YhPhb0J6OmnmIBjrDhogeuRwr04TqqC4/rAJzxzvn8STzbk00uAz1nNf7jOxnqOw
iHggxvCSK1v5aqKznq5VtZc+hGwKnVPeHyb9YiuTf4P0br5nMHadrrU9TCmVcrB4
3BYyoyBws530HIEh+KjcUTquFd8wGnUzrxfEzMX8ILnkqYIgs68JqWfCkozr0iHw
iW2lWiFS+WEp2pLV7jskiJbjptBdgXfV6KHtFTk9PDXDQikeKOsSw/8ooak40O7/
I7qAsSpj+olxgvMjjsBOFD5PB6OQ9BaW7RSbYRRZMQw0+sMr47CAuyyabQ6Y558u
r4C33NLkvaQL6jDqmXnP3Bl/E0cOBrOCPs8Ogh9lhONpUXFkcQOEAO76fahN2eQG
heUl1i8LLR9CBnHdPKwQh1ae7S8lE9YjIkjLhHuIyW3GemqwdKr7X861MyrA/OWN
W8Goq7jfpT0pqkZQVPM5jnz/uKOz8fHOlnrp+lP40OkXuXCtvG3oYcCTGLoVCak5
FuyxdzKlrjJ4kQ1lZ5lHX4BqblJf7DYjn6YmRxnuTQh9mHiR3n3ECWQQnkGzd9Jl
OUg+al2uEXGmvpeYOSxs2vsqsuglFTnjPiKpmChdMwUfq+T0gN2lJtYJ0RIzOY32
LG1Z0YmpkzrwxY38d4qcnkYzypVA80k20Kbk52jQnut5fwQ+obpGhtrIDfx/cbtl
3YpG+NRbkpIuY+ZWRHRDf+EZALRpRuyVARHpjVbVkasxeKLLs3PnmHedxdeKoiWS
nOoNLqvU+JZvQE+X4JBcSPLq8Xzf/iFzTv0VJd/yT6h4MCo+45cUffZ3CWpjDFvv
P3r5V/Mvwl3D6WyjDZbxYESlaJvq8QxGgpcsLuEW9ECr5dkm3qm13LiLG2Vq0ONd
nnDICHas8JjLvOC6Bn7lEJho2kzNGNF9a6jF2VqOtwxgSq4RW0keIIhIFPJKwYLk
qT/UKtNaV8LtgZwAv7TSFd1YBUQoFxolkAuZeVMQqdAh5VwQUgwxZPL0/Xe9+ppl
BfXaR+eYlli5tnWpBcbP6mvwFSEZRQ6dh+NQor5kmFpNG58ZzNfsjdTZTPnnyzc2
2+4qLm83qMNmIZ1uWY+eX4ps1aVexNBSEXiq9jRPC/bxMwt9oniDByveVdSrvlLY
vGzRfklSb5Wg5+/A7vpX85YujfGMnP3wIw7GkZc3aGJ2X7EwTWCTYzlKBq7VJ1yg
2CMYSCg6LWsJO8rvUMNQ+MKRuxOq6L+9fQ1/0Njxnm8oIEzTx+DYzxF7QuL5Qdcd
KljhrvlwKEHEpP/rK9LTSTTCA95dSxCQ441vzse0QQhmX0QSkYFg3BST6N2YeI2L
A+uiguOkuHDDReXTIFUwxfIfp42wLDUZjy+xSzK2eT3M7K4TrzSWhxBQ2SkVcCNB
osnsoKlm5M/MhtE9sPMf1+61X34BxUEUqs0oPxDMYKCGWaiYXL0RQGREOQ4rFXUP
TIHEsT5TIzkTt3iqmKrWH6NGmK+FfQUhc4TLhrJv7IDhua7IU/cH2R8NnnXZz2S7
TnDA8aHEkJQs174QRNqtRzZvbDnSfl9NpAa1Jux13DPn9UMIr3T5Yd/x4WlSVBmd
gVetNNC/y+RX43hG6pJzMqQYVxo8DC+Y9ocpukTuUuHEj9yT/nMV9Nt8CvxVkxyX
J3qqXA8V54rXWXaYbNPx0trJEroFeu3uIJSk0ckZIrRYIYnoG2MpTSw0hIAsr4oC
9Ahy3qbo70z2ZSWLnbpo8X3alLFxRjpU+Th8iVWJRn6yx+9HZ5hHpHCjpY5OOtbD
6Zoe1zMlOJowi1l/CDUmre8OrRdA5Kk4GwToHSTmsm6QFZFL7JJnQti4CUvgH9OT
ppUEZn1k7qjy/4ug3A3mncFDw9o0WrZyGSEREmj6KaP/EHZCfFCNtFE3FoZb5qov
Qw1ha05DE9ARuO97dC3atXuRpQHC0r6pL7uEm6NNwYOvhqzvooNV/qrKjZ26YdMK
uiOjtUbQq4Koc/6c2IQ5WdA7o7r8R0RS8IQKJxwOhw1zB9uPa6i2+MKYANY4J5rC
KMPHtgcIuSxR6Zp84XBRyx+xTvkXMdY8fLWTZ0ZYijsnfLEsYI/43X/YQdxnB2Ze
vXHmmZ3XxDoKr9YaysA/pbT+87f0qflTU2mazCY9K3kxZEN1EaSBvxedrbwF7LZm
KsMVn9pUR2Rh7/jQrj5TqtFc357DGvQWtCVFV3BuD10iv0O+sP3P4wMDkRDjCYok
kdW+qngxqAKX3cbDzw0J4qHUz2OdMD0GsyaBfuNbNSmSnYHmxTDN+zi+SmfyFBhh
8AaPFTtI8xiPsd5aOpFj7mJEHwsha+xfn9HfnR1fiSSZunRpRe++pPLeCD9H3T83
TJGwcCY9rp8KmUi118C19WGYqYPaQmRKVPSt8JcwcZxvkaDJQBGOl0GxRNV9lL5U
a1Pj0r8YYty9hoKo+UdZDWGAT5QjrftGUpC1BEf2+O1/BkM3UfTVCSrW0Mm5noPB
vKntUTzlpjm0bhHf4qZ691pXN2bsYte+PRYny4TK/o7L+Rt/aecP471lG03tqw1x
4qst8Lotlq80UdSz2bTv5opAaNPekoWKlx1s4D/xGuhMeVIewDHzVYjfzO8aSGfz
g58nwaGUtib3MPl80Ph8xJxoflxd1dXuvxdzUEJiWrIlE8Qgw5SrY+7lSi5/MVio
Nhjh5An26PIPjk2dbZGQqePb8ATwDlPHDeu2pOmVbqZf5+G8WFElkCfTNe8qNZVM
ivUcKXUO5qOqeu1UurjkvrRq3ngCYB7IgUN882ZuSQV4eEAze54Yh+2Ra8W5hqiA
rPWHvqwLpZJPN7kuPuB+wfhUf0QUXU3cYf81A7MWFkIzrEsELGKQ+Pgk22UBzXWk
1ZoCUsMl9+0iioCxvfjlrql6xcriMOuK04QLzktHbo4a1kLpf7ZaSqlX/dVTyySS
MlYhI6iCIbHOq255W/bjchC3zFGb7jODGtfUbHvcnzBaiscxiThthYYWIjuwkLWb
gqHZ2ahM2H8ygp18RmmnpM24s9GEe+jRdeZMZ383vQcclvwVgGXQ9vTap4K6F5Fa
x7X06YvdIuNldlE1WpZiFvvfKSm/HUG8WalPes7Rcx1T99+K6ZfpnQQ2UO+Dt7G0
Q4zSdBAoPKBhLrlMVA81QMC7gzb0I1+xpW+gALUnILecdVF2CPiHbvqYZBue0oUb
LMmd6R7LLz3rENhXVX9g5rfJke401R+WOduRA/ZoefYxWi2ANxYK7xdAtp+b9Og9
JNYo2yEZQnbuSzcDUBZjomoHVPLhPVxHoTKZXpZE8co+eK80CwQKiBG6k+sv7VOH
aCgUyK1fF81isF82qkjsp2gfPG4iVAd+BeD0Sot+CsZDrbqj4coe03h6k2FYcMRi
vfOkESUdih3Smo9a3Q/7OWAXhSAtG62niKlC+XIaFu5eWRR84D/5DpCEVNvpSijh
s3PNR+N8A9BP0nRe7SgfV0bAZOAxbOAwXf4nuX97ILFFv49axY7lrWHczNVVI4RY
QJZkLZLPLTHT5WYUHvlbYYVO2BEhhtcJ8yWZgMlLon0M1ogHw+DCF+KcJHsuqaMh
PciCLEXpcX6HkY7BfpGUOs7Uw7Fd+tkLwbpC0Lefodc44aoZSVszADVX4LsUYUxZ
6EqCmFLpeTpJasFvooiBvj1NsJ99wyJy1sk+Ue2s6/SnWgStWjA2tMAH0rRqnk6n
ip3DDl4mBz+kuS4dSqajeYJ2Ck3ynxq7fOleL4V9YRtGNAEuzFy4L7aMom3iN+au
OYuUwQoCfxFqJLPeatwKM4QIfMApdojVnpM2GUWD5C0Mxu7T5WIF/+BcwKitA9Kg
KdOTvDF4pQODVpcHKEZRg9TvKdQZW3W3Um1Vq1fClLo2f8H5lMl01f2lAfyCe5+G
1uszoQrCxY6OyPTAY6XWXGwhgZolLuY4XXJtFNq29UAstSE7XI/H/C7/vLZEwXf4
kydhakRFyWQnctd9NJct3QCPt/9Qcps/q41HIWznbTOztq+le0FG3166Qtj1uJwx
+wsl815qoKYcbfUAL/QQH1YHTebNheYtYVRSNnf7wqC5bCau/3ZJdX9l6g+NJvGX
JPHrziicYn/PpBQpGOb1mZOEC+ahAUYygItK1NDxf0ZrI/89k3wUc4UuiQoACpjA
0netR9rlCqy38mSBIwxPefKt/NvOACVGz/Uw60HVUmuOG/xUg/cGOHapz/JKsAdU
ACjl92TARuUmkAquAl3IjLWp1xWkDctvb/CLxRPcU9sREvY4YvAIlVSfJEBTPRHn
5svbtPpeujZp4/66I+HPTkgPuo7rDsABN0CXQlqnVP9sEg7g9ErShLuhdsC2+9oO
xK+ffcHiBUi2xyTLEePN0+M1nBm9UsE1tO2KMRmt4FghdN1HJQYgA9hWfwXptniU
m2uF5wiITmUjvo5JnK1TNYGFHTQt4fdmKvHhczN/2JJ5AABYpXHGo+jzcgcLPDO1
04ic2IBrUZfDZFbK9ducjkBKjUE0SIV1B/j7K4tcYho50FkxVHp8BzLnYoLFj5JO
9YRhXhTu4/gM5UKl4jj/31/BP7cYBEaOvZncPPmK/Vu5M2m5hzTixAuS81+PLPgB
6n09hHJ2pq/Dgx9Cy/XXBezcIyzdZ2hR+oua2eU4vpozs34UCFOG4PNbV32vHlxn
otLGDaHGftoSYucqlxwRd7i4wQawjCuF60s1nPFyIu5d+huuiS+uX9obSKWeL5u2
2TUlx91uz+TocLi73E7XcVWKcIriH7mRlf64NoLO2iVjQ6J25BdjNDTXlJ+TWDpq
coWWRVNuExQRi26PbMDtJyR1jHfj5Wd6SK4EF4GOk3ppPd4y/wvLbamfvGMF2oMv
IpXG5xQGFTjEOxtYswmJY2GJFDNv4YNJ4WPj8J13bSjyNhSjyyQQlOjK9/ZS0l5X
o51drdqTeGtXlPCds3jZAefTLcuYb4ZGFiXmqjHkkqE9x1VcFyUWNHLTPMKH59eY
9PXoM4m23NuCQsnn7UPT3HJntMk3sIpPQ0fEqEWqAX6DM0VahmHhQE7c1AUdL/1A
UhfMswCArvzuVUwH4eWipZqGYCAQnM77xlckyRQPH7xCNX7sVCiBVgLgXg2jpuIu
ZsSMriP3ZGZUEcID5j5ZXDtnejMdgt335DDF+YesZHFyRmVwpKJQ2XjEhxgRMG16
+uq1+k7CaeNCbpm5IWxOA2G2Ope9Q85NHyTbt+F2DBbCAO00+jkCsO9tP+YwcKpW
L0pYJol73QzB/dpKuNHB/yC8GNLPoPxSVyOvdpLFzXJxXtkvG3+fDgcDgmxHHmg6
pokgJSCGsva/RNaP9C8/kWBBjm/kcMjmo94z/X/gfhYfg84yj5A2+q+YgbaJ/fna
dtHnVHbXAYnyKd7DsVbu3/Z+Sj2Z+P8urJ3kEY4WnafVTZMZPNjwyWADY3TRAhEu
1W6UsSkTRSzZpfP+gOX4akVdkdLkQL2wDXykgWW2DZ7wScR5MzY1KqLOCCxqpc6G
Rw+HnGGdrXfxYqBvlbRXGe7PO1i6/RHgOzjyZ2aSO9b8Gl5zJHOtfK/KZiWS4vGd
4SQaEdE7r/sy73H1SYj3SXdEebG8dWoTwThNN8qli5Xvm+rqssugpDjinCA9GnKw
0QhHKLMlP37LzJ8SB2X8XOpb7upRXSylPWkgOGohvi/coaDamFLF6Ov0xnz7jAK3
JwQ9CZWmPNE3VLzS+cSpAiy+loi+MO9y0hseQcKbKbHJJ49p0lM2SqbPBlmBrMU8
UVMXaiKY5xEeQeps5mNKjTGeBi+NyNv2bcvTUoQ/x7q92b59AXmlb1yvpsoK68k3
vkFLHFv0xWcj2caU47G8ohXlTDR6VCsdCX2RkijU992vq1/Lry8V+oQ1roz+S4iR
CGQmP4ZjX8+epvlcrLtIQ9fbo7bhBSYCuyoiwwb6KNf/dXk8nEmS5cgwyupC4ayB
ZUtGlsYQdCi7v07kI20q3RdiVV7lqMVwMqTMf5Ai/6i2MvHUtCPx82JFJkZaRbRb
TwdC1GlhhNY1+lixrNET2+AZBEsgtdRxROo2Zb1/4fHzYzZgTp8mVyl8qdhWoI59
t7bW8JO6Q69A7TLs29UwAWthqdQ5MAdc2IL5f7LAzEY+ezsLoxVJSGXnQpcP12BL
LFN5eD57zf4wlxxO7Oe5U4bJdR/sTDP1uMUfmyxgiHLdFK5siC5wkgVn+rioOcQf
PCxIp6RbD46R3lROGQIYTvm0RSJxxlcTkuaJkAO+zFM21Zl8fTFZZr97nuhddqXA
zeGFDpQ6r2NMtXn3faGreryEi3Y5MG6reBwWXSfP8Oa93YxXXWafF6+f9chBLNOI
Z3nwVdzQHbhdN5Dyj6TAyyJsxbn3Ly+tuXhjMQPvoqmGCToiyhBuP87YBHeNODxb
LFCsl9Yaf+EdQ9A6dlveyijBlxISxRIBolOTQOuBL3K3/p14R8frZCKwbM3n194a
mxeu99pTyFe0Th/wS/YglRQ8GEJYcZ7Yriw8C1bOyJ0utC7XTjH0uWY3OqRCjwBp
i91kCDhP6xQ+OeTC4BZqGqf5PnSkCaAdQs9oc4O/opTcI0nlbTI7lVHEwOt3KCy/
DHCT46CPxRyypBLNmeQkLCfD6Ca4H+s2P9hmdyKk5D6/uAisJH14DwooYQj/6eNZ
kkzePfwiN/RSMocThjdZYy/8oKp3OcjMwddoftycnU8f5+saaK9iF5hJXV7OnIR+
RyYKLnHWgwdFA/37i+4HCBOFZzLLHtvAc1NGDiIwNuNiLzh0MfDE84H4m6dIqWOE
XqsIDF3ZtmN3NbirXrQj4H18fZQeMKURbXSNXshprIHXwHLgf1et3ZcLJCnakBGg
Hj1fuljQKaY8O+wbz2D2omSyAysbFDo5I/lZtXvf8N73dBJX+kKqPfkeGpeNMu26
OwO88dH+/jYYCvn2hvQvsWxGI42sON4v8/JuCyFUufRFp7PhM4WFrdr+QA5NizlG
gCo9YC1j/n/994XZcdF1Qh8Nh6cnl6w1wnR+vMuut8/6J00j4rDL+mzoAS1bEBO6
tClhZ0t0F1ZKDJ6vvNiQzz4mLn/XM+0Qrzing7X/IfsSuNm7iVpzbXe/EpXPGwfn
hNipTSbgU61yNh8BbYQ2f2NLu8PqjhiUmq0NqfjtwyD8cDwDNWOW4AlQ3Dlp74CR
HACAIWAprza8XBLvmLyrxnRVlQhHtnITjtKUX7ygvJApRcvQxvoM5+oHCypI56XN
bNbV0Mzm9naS1UGj1eN1t7WMB+cdaxnlLgFAQ716qpIL0Q8MFGeuxRoP+bsz5tWW
0Ih903dZnoaFTGH6MOIYsnn4aq1BijMbYXC2VZu2O/Ps7HPLbSSPwUesRp4qhVXv
6w2fTe6RBv8ePqo+hVosYwDIopY8avPL8n+nkettQZuOWCUkN1WUlKy+JXwTYxCF
uhfGsT78ZNmxzICSGg6BF2A6ty15JvatliSzCJ7DE/UG0dLF16frT/Ecxv2OWxIn
MSTNuMStWTCFjz/BNa8ohhagqSQDzrxrCAcvGYEAwN3upagfDxmQbLiPPU8KFAc4
S7MDfcnycnlbWvqkbxtniaO4Q1i9qfavW2Xh7bts1skE9HREwzQBMmHs/9JY/NzC
pvTGhQHXEarIFXlfZrJptRgPLHmDBsfjs6jZTLKUXnak/8rKRdjfGLhe6gCJRMmW
aMAEXFUs0xw6cEj16tRHQ7LmbxxUG8I+LeirhgYI5n16H9F1ZffIzSfxTC2llUrm
69eyl49LdtT/GToE4bRUHBPcY7oaA1JmZePmRK0JrH89KtjlUjsy8h4ue5ace/cS
UOadwJQySfvxv2JRmjE33yCy0C2Q5x4GiiQbJ8ZHzBtCN7AEM738nBhPrl8gwolI
o+a/Ar6TWs1IlqMXYDmwlfpLBMzPjTyIapgSjx4yl1wHTpqh2h4yIP9MznRC9e5Q
HeGgSROjP2AnJeMJ0Od3EkAbGEat0BfRUmpVDQCRme9oIA+o5R6FJvPnomtTGnOA
Qp8N0cCaAGsEsfOy696I4Dkfm/qg6nuksTspvBktNot7ypZuBGSKBO6gNbEA6dmm
BCGFS89gqWBZfDYuBFre8kSU/c3sgxzXBB+VoozSHCgAsK0EHO0mtrTxotx8t+kq
UKv2Z9/OzgBpD7BcPKKeH5l3V3WmshLfU4dxWyZxvSQa1F98iCW5nNbjMu9dDA/e
6N/wyheRKVf4EDAEKPVw+j2DPSI/qBZBRM3PDl5NkhEMTi5wNIPNE7uNOot1HD2T
3vPJe1hdmkznEzPBO/EONFXnnkPJ2lHiJnKNtCPJrbEwPhHiWpCMIEHaxI9iV+F5
WsT2QllrHxPUIwQUkG8t5GXFnmzPioHPZdwTBLpBS0PJblnLeNm2v094J8UOajPe
PY1IrE5kJC14TnrcOSTtiBaEnXy4oB5lnQurdYVbU4uC2wx9HHmHGN40p329pFAU
Ppqmyd98j/Ydk8jdnWGruug0wuUbMd06MIIQGNxN9Xxu2jyaLEt9yvIeyN+UE+lm
/UfsouatAjVek/aMY5Vp25BQKeKBqCBQl6iIXENCESucR6MyKihcfNMm1nx0vrKJ
jlWFoTA7wDGic5pAyye8RKur2NMBWPAvGzigrTaHhdE/ufNRbNPxumDA/oLUYzE2
+RnoAQ0bv9DBLpTLK1e+OCdLpELDpzJ8P0CotwrPu/zGYu6C2viPiABMQazNfbAp
tCHzYnlpxv81bQbXWyJsSwgA7TGm2eBUB2fg5kLJ9hel9fL4pZvHl7+LxJgxVuic
Ro0238JHyLFykXsiwPVLrAi+0etLLOGuQcomYH39xJbGwmKENOnlgfMP+NHszfyR
8eTwvBF/QPln8TcVGaGI4uCHLULNImdTvG1HxNREno05hRhT+RwovKeVwa5ZLsrJ
comHp3Wr6tt3APRDxxzquM6i5dl9JKkwRJi0A6mUAh7QrgjaFPCmlOX8l0xXw7YW
7Ntlz3/R4Tsepz2FPJ33w4PUyi19ZIvkBNs+ruELkhY08NTl1dOk4HQWRCni2h+8
UPPzW+ICituKJ4TxDsyGlSjGvX4y974TO4mNsSnwVLRUrKs3t8b6z3fA/wyGQuWo
MOuoDpLqNp/jlo/tkJteD2MJ7M/B5HEG7ERN6p3W8CfVnMcJKzwEd9O9ukizHIra
Cg+dq0rtC6uiVpYmtN+ToQ49rZcf2yMxgVv4d1T7+amDNahVatyjllbqHEtbhuTm
zmOE2rtrDN+Ozy2ndbe6RwEgR8cdNGsstKCK+dyHP8jBWyEkJHCjc94zgNJuKQzo
JgHuL7NTb4ml3KZwST+hzOUMu59M6dt+U1Fk62Y1dprYKT6EzslspSfD/rgSJbpY
9cSz35oRX+ayZgMYWrtPVu1jlKUzJ6NESbmRJpmAEfyHNae+e0X4iQHsv25cUPBL
KYfAbmWumK6iGMnKuw41NuJBoV34y3KuLNPGnUdoiNG/D5F68mYJpd1j2OF8wrN6
jqzNuxyYXe2Jpoc42zTc7q+LLy0+2hadmlPFMWXwPHD9MK2t0eoYmfKvanXBYLGp
wtts/RhlR7fyIBAX2YV0+GH3cURPUdNaLbMAWugkt9kvn5kVO8Vloow7ykF3dAd+
i1PyziIOkGMjIgaMxwDZwzdU5i+kg5P760/4osj8TcKFwI0yzscPdE+OkkWR26gS
bIWGVo1Wxoy91DgaJl1t9y0+csuMaqxqrHAIc0VhCBOA+q/pPgKRZrLUvnILpRGP
Z/E/Wliz+wj8dZ6ilIawOUloWfqs8Ft2jnkP3nLdQuy8Q6Jceg6qWYdGriq0cUmo
OQ5UDLq32LVDFeFs/zIdX1wmhzu7EEqV41Ork2NDT0hB0p5vDLiJDbs/1/6RbLcG
iQaYkr+FLAlXmvBJsxLyRIkWBTB6CjGjckHOVVPYpxxFFWVmShgb8SDcmUJEGhwQ
h7dUVm7QonA299gZqXOrbJL8DrhIph8j2yZH0wIB1uTzhdyNxfhqraE2w3UeVCug
lSqdB+Zprgv8pi8xiu61bovu2Z/TdIwcPDjNE9eXeyjJIjNzvIR4mauuS6I3PY0t
6bUJTw39t5cnhbjk7jT7j6pF5md0YjORFaOfu3rk344gKDP/nKs0YquNPbeZHYNg
ZdZ8lw3qzcYCUtOqf0NMmXVQSrZbVb3oTXjLpydWJY/SX633b3ibQfNRzFnUk0Wd
IFrDrVJX5KCfScK7n9idotF6lBq9JKxT7DZcbm824x4C1v57GeSWXsDfXIUgDRGZ
XpHn+aaSvBmoeBeEg0JNdiG0O400zv5EAD2DFFw/kEkRnTvE9AC2eAT7eGOkCwdN
LyXeAAm0m+zwWfw8Ho+kcY1LsF/bn/ccEsjAzXD6VJ2JVmR1u3glIChDbr0lqXNs
1Ah/TpWxxpeM8Iz4br1QrdyXzl2Dim6RUKYGNq2cxAds3iCsQFZKxxKDEbIEAI26
S2CwD06F9OWzhsmts5YNtn4sbtkaruE/mSSru8oX3jNznctJ0hYgmhwyuIxoUPb0
CxYdt2gRK9JOcGoiE8dvivpMEzQsDnEKEdC8SoqhTTPzLzPtcSwbH6Y3066KvOqX
JwMQPtAOgDSpiJ7GFxF8xDsgcHFlt63APJHlXIT+Da1bZMVJXQHl1Mtsr1wPUEws
AAe1A1DYM6nBpt6BapnuCO4QdPKicKbLlNHk9Krz2sRde7DBEnRfLEsHaMKRAUla
+x8tvzj6kUGxlq4RrBehfLjI0qlUBERqyvfLYfsS4/ABmn8u9iTM/32VH2mbvNP6
/wVB6fstt8EFgGIETu1pUT9CovzcOx4/qV1G2mKOmTLHqfPU4b0demRpA5WlJ16t
iAKaRqwi4HAOhgo3PFGBzd6ODMMZseezUio+toZ+BrRumNnkL/9tjj2YuNjPGnG7
4L1AO7XvqCpzv8HXCz1zNWe6Kvci/lljGDZMTzpFWzLavEF6Mx8MVGF5h0xodMEo
mNfhiTwM1x+NkeIKB3AoyRxB8Ocltbbm21cSJsZTVBWp3KB7szO12Cf8EzIR4Dgl
0vYb0kivF6CVTbAO/oi4FfBhXFx6YB0SpvjpVbm43ec33dBxu/znwo3yDXlLkA32
gz70iRAHbhGm91438J3ItZRNSM4H3FFoArChxAVnQQPqvteo7cQg4B+dq7wLGB4M
GWk7zpdad00j4n4dioWOaIFebXDPssPLiKWBFn95M26tpmCWaFPhpozdhREg2GWn
pggdJBJoFTd5EPsFa/pqjhxiBQNEuD+89Rl26+RfxNq42PURVpwbJAMiqJBmrZQG
mMr8HDvF4AKtjoUI3Kyjx6SW72HK7EImFSawtKL7gtST18eepnBtaGERCvE6T7+C
HW+k3Ian4w6ua/U6lRmQj0IpF65W9fpHcO6pqergYMxDFRFP/fGu2iWDtTcQOttB
mWGic+lPhHOexQI6qm4r9ZtJdTqDYoqK6H+sls9Vd4aJ/IdBcM3wHJu8svMqSRxO
JlIblgbFhU8TO99GtAdB79pGogoIeoAnDfkySl2tQ3sayzQTpqUYQMm4cW+5TCOh
+wTv95NRT1DvetIH1ipPhHShMVdGhf6+sKMpQpWdEs4nb8ma7X5aXGun8t4uel0g
XKFjjx+MVI337fBYfK0BCVh1i+QYu7u0V3zMCUjNHdTNd4FawU8eCcMPPkCAzpDn
YfLTu2PQoCZCx02eib2AtBP2HedDH4E0pbNw3J0oe0/ITbCUmtNWHf4MvduEom7z
ezFzjV1ONMgC18d5uvcVYHDYf58sFxGcF6j3qzRNrlEJ/rlf0mIR6j3GyP1nGN96
Ccmk/2F4/L78DAbJBPOA4yojTRfDKemT4CNVFGH0jFYYMEB4ga2cqo64WNnGJgD9
+6BrBM1Ey+wQMBkfelhGs6wOm42ulvTXS3IPI622jknP13RXMXZmdLYj9AcCPNHL
V1UJUhmBpONtP4odmQHuGrsLBTXjwKavZ0ezguJxIz2lqZQGWLvPQlvyB+0/FWVd
9DuIDL34f5tFQeeG5IboWsRtZGjp2TyVdp+jBQ9lpnOTFR4gLVDRt7nNCkXNW0fo
udNiVjEU+vVQLHRrQl1xEQdnnmXASofZontdcFcDdnUEheEbN3d0+ZDvKkG3GYS1
QegkKn+Dvuxpa9CWQeEvrvnOotuQO7g3Y4Czz3DpKVNUsAcnVWgseJH2fHd34I4G
nocGU2dsqQqAEcTTIhgX+2YCWCpml8aEHHI6daWawtJt5PIi8wjBI/8fR3ATDu+U
n5khjhxZevY+ro7LkNrYX+wEXllNTKvHAg7967xbjft7QOsZJiLTH7HH36cpOEQW
ToB4oexwxIHDqEAAA7Ebp2hug2mCf17JhGEUGkx7nwobCjLVbS0vdnLqP3bfu5+4
HP5ScnuFEAovchxZhIe+p75EbXbwnk+bz2dDAGbp7kgHrpC38vxliY+TXqyLsUp6
OZHpqPtp7wV2SmxVsg7BIJmhZ68ICzQCO4UAM0hxxfVRDJuodv9UpCB9RY4bgVBX
2nyKF9cGYTfx+/BCua2NhxjXZFLUCaxc1LeaPDmS4AgE3qfYPyr4vOUQKZS1LU4Z
tamZ45IJCxROSI0mO7c7jz+khl8frxbhIy5QichU27kwRQBs0x8gDkJLJh41Irjd
REAPw6B7HCoMAL14sj7VJV4J1TjsQq7CntNp4c4KsGxI9z2luOoPpEfRuyD7QIUc
ZgMvW4c8p9Aklhm127d+DbaTsUU9KZB04jjkKeT+w9DcZwUiqmLOFaypudA8JVco
7/mM3hwaQb5Hn5gYhazveinstl82lsZFJQM0BPBa5jWy0Z1VIg3fnbs7YuCvRtUp
uMv4+E7h+M7A9cJIV9//+2LaHpmu+KLd0uA5HjCO9ZVThPxMSkAxg6PA5SO1+FP8
mWfHHUACsaoj7G1iiYZSFzi9A69IiSzH7OuNYjLy9fQ92foZg3k2GvOo/6+aZXBJ
/HDGfJOxHrCsbcjCB0D4AW+yUclmgXnjmPHB0BbSRe8aNPb4LqqBILJ/YnwBXWXc
Pv9E9MPcpNhGxuPq2pDhwOWEgglXWgKbFVna5eyd7PJW6ed09d2TcfqnYn0shqiY
a6+UecqudUM7GwrPb2U3S+f73viHqeNl+pZwtV4D4tjhWU4OHOYMStA4o2JfkBhH
rEsWz0rpTQABvPCnWcXHyR7+IJfyTpeTM6yg6GlHphCaJhUze3Vjh/UCDnfCpO67
e9z0N5XT18t8uAyuO7uxn6hrXqv0hfPtGZKErvuzzyW9JRIn0tqF0V1Z4Zc14hMj
9Wj7bcA9wOULrTfAXcdW4y1i0QG7gyG+qGWirdxQcwKn51HwblJqCpVnBOhZxPDu
+gzflJUryhPh+qSjMxML8Vatrq7WFQE9DgF69GqI7RosYC0TLzruhDTUZzXujAA0
mDXMK3bphHEpDb9I96Fp6rh8aE7qivkkNmuEM4czu/T2VK+1/Jxo0gEG74uJXwCW
2/Kg6s8UpVZfW2FQxVdrWf2n3Wx67/AU2WrVUX4ctNCQhaWaDb77DtLgTCrJZ0nU
PTMKWOeCO8MK/BYqE+gFOPmrajkmVoORCOV5Hxr2yNDLn8Kl5+TyKO6QRMDnLbRV
a77SQbZDQtikpJ8Ze65jFPTZeF85psm9cF/OlPXlxBYQLVeLIZe6NbZ2E1JCoylr
kZ8tdGaWO72kq5akJDw0Y2ITlmVMhXNx+ZnHuizFPVEYPazwW9P0HLPdJ8W1Nl9N
lp4KywfEh3JNk5m39vqoEGPrDh2kNYZUodu7RR0Hl1VMQcpOpHiDSLYBv6aSMhK8
sMUPp1dwxgs76ZpWWPPx+r+OI2nG9ZoUFFXjqGROobg18v6hxHa23jPuOgpKzGnR
ru0/EVpBnfCL+D1Km6KU1oz8a/0p3RYNpegz6+DkmNt5Zpvi1WqbT6pxqU2qpU2q
M6VFx3DF++/PuBoInQLsSov/XZHkGLIhC3vtrvT4mCrCwwyuHa27Kxk7mZeI1ecp
tWA4IgOFgYM48NOoHBLdSGtZAsdjyAspVrs8IGI/9mN1pV8ZBzkI4L1Z9YQRml9K
BMvzpCNxqZjkh4dpkaCKPadIVMlHDWmm/7Xp5B3v8dkLbuml98MNY8k/dtNghUMV
yb6olB/bpmvd6DZW+V41Y82Xrfzsz/spxds6pqFKTkYemldAaeUyrNz25RAF2cB3
QyjHaWuUcc/GUjFXga5hI45R/ZfYH+A2HVWs3yKyMYhuScLpJaj3a+eZLvDtH/vA
eig1KRXsNGYYZrHWfmjnapC7H9WE6sd9AK88gLTPYClQGT0zwYBlbzk/AmSGafrl
tMmei4sJ5VBwRu6WkJ8Yijw3UqDvLJkC216ospLBujyoDJ49Yqkn3fP/r0JaGTWT
ynoao+voYQqP+QhjdnIjGGKFiAVuOlJ/dKVpg44eiSOyCL5nZMBc28ukLred5Oat
Ow5ssNRN0H5/7MJaKHK8bqDuQlst4OaGanb20U0lxTrPYryWsa4dFISBPW//t5GT
m4pv+KfeeGudcvPwNOaEhh9HPSb4TETpCk1xzLe+mBYnN/xFlAUmvmpJKDPUHvm6
qpUmgStSt8wApIE+EAl9YL7GJ4K8+gMMdCK6Wd2G/7K/DruwGoLkHSfm549Jnlcq
pJAERU94evAyllE50y3Ah4zEhKHdsKlUgFSfPXAA2Fz9bWCAfN4xe+/3hiIk+CHi
2ks0rR+L7F6VL6Ai+6FDyXbWd3Vh6oXYSqGh9SP+2iZBh4dUsw8tfYRgAKf8U6Wt
9umRUP44w0fF+m43M8vYEZfyLJgERcdyHvgPH848uSjIS9Om5lBdnjK6ZY8cClDd
5eow6IxAkTBtDEYm7KfyKpOpGPh6aQXP3j/CESqMldo5q06ggUz8JyNY57FjN7nC
cOmK2hVheCZWvYDOzMgySymn6eam1xlBzatWSxq8OwF7Yltv0Zw1vTOPFrfg9Zp7
Jw+inB+kmcDaNn9xpbPkjG5HxATEei+eftVTaR22ED1Dj0XCubqhh3kMNqxuVSGt
NIjKWvAag39IWe5UWj6IAOpjWDnQ0kKTlVtfsvBgvkQP/8dEoLSGKpRkQtymhsvr
5BWKmncPxWBaHGW+eeyxt/HM9kXnUpz2z2R25X7riizbS1g/bGYB5qXzE1s4HJa7
QnLgOUiGc4wG9KF7hQh27TjEqe67AYBi7TXtiLeZyFvtk8FEQgFkTgWliB2zrg3d
XKqDEK4B8bshX8zkyvlKjdQW4x1v5QRo0R0tb5IBv9hpHn4yJcErl9asvzUGu64n
qDZNP7NOMft641dQjOftft8QaW8f+HlRSBEUfpfhn99J2fiJorDO5DtEh/VMZHfb
0RAwP9ngcGoz2wZf/U1t0laVgoaFbRgkR3lluA9nSUFvbGtpCjDaoRHvJpAU/m0u
psc8hRjeazKLh7jr/UpQrUO2gopaFEBggi/UV6obY8eAGuGzSDWE5pnb9MfOZQcx
qBioeeGwWWaixJLVbOe5f7pAu55/g1YpLY9VY77Z3F2Smg+0qUfO7dLFi21dEXo5
t7aeXxqEPz18vef8yXzgb+04vUUZtc3C9aoULp6Snxr0sCWAsEXbCsE7W6pOyScU
krFvRbPdjWXr6HUXmGPFXivaYG8hDB+XaXAWehBl8+ZdauoZ5TDIUN8xpQn0MqAm
+Lml+r4178MK5XUCFRr9o2EGl90TPj5yzbLQA35d867ONNZYcl6W2F9YFC5kd2NW
3h8h83iyheKa1gUwIW2+5RONeNJStYI9RzsuMroXiK7yA5BbB+vcgMnwFtJG/3sR
R1ANq5Z3eStWakNbTe4v3WGu06rPnMYx3Xem/xVuaBlx+idL76HrQ17g35YpfoYd
NcB1KsInHlCbM4v+fPvRL6B4wSCAKpmF8aEdBil4Sbwrv5Nluu3YDRtJ7ZkPMgSH
6J0rqzWWxd/4rxe02Nn0umezuF4GSE3GVD3zTh4z4uFznMEnQcw3+y3O/JXX8yxA
wHdYkEqXBQY4VnW6fu8wqxi1ZUtsRv91EWETZN6+erPIaMAa08APslTk2fJYZHve
LhB/u6Duilw3VWbYnitYC3wPBqmPBt3e4EIDg5WTM8NEIdWg9JMJvZUgGs8gshxj
4qMK54PvG7FG96cbM0kGQir9HcVYdDftBFfbMH7lTdlSRJAVSwQFrAf0/yROQz5G
4zq2ZMMM6jZMY7ZePPrC7KWmNpftPB0z/+IUpvV3frlr10Dj1UKjM+tAA0BVnNCJ
fIsc5N+jvJdpNFwa3G0NV/UDOzI1izOWFEDIjD2WR4t24FV2cV/MGZK7q80CFvS9
vrCS109v1lNCff8wcOd65JB8Qkq0TtJ82RtQVerai41ztV2FWeEdQjStlfqmOUZb
0ozX2/w4FyykGmJikNfh0QC4X85zdtrdjBhheabprBdxb57OQ/i3JK4P0RelA9RV
lSAv/pf1ppr5toPDb3g1bVNz43gGZHkbeCk8RyWTLMITipQvGpdjEJWT/SP7W4DI
8Q7hctY7APjybqSKNorPLvEYEEI0Qghlx1VzzzU+89/IGhpa5UxU5zpvnw/N91cy
Z5CCL4+PFQSkTApsPPXFlEeUhrg45vnanoql1rSkX4oc/cmx2QPVKLltpdRUAXmX
OHKXgSONUb3TeJQRahMPg0ZtZ+vVWBgygJxV0pX+G1qqoE7NlY9boDxCqTbaAn++
yvta6WB3WTxFdnlkPmSzN/QRkU2+BE4UfAZ5UiyHoAsx6t2pepBVglNf916SVKig
HrokJFg9WMNfizXuxyUAHiRLMmawdlBmpZi7R0wbOkns/ibT3rJs0nW52Y9KrHgH
1UMAGfS4QSKY7wbUlytCc30MFMxI8IY6SZan/3wn9qG984Ea4NfKb7p02vMPuwa9
sJ8IO9nveG1735RUlz0hLbF2v6RaHVgxjw1SWIVnbqA5nMMXUGS4n/zDsdI8JqMw
gOqkM5r7B7mG39udu/ZmufvWACtCvxza9FdWSrI8GiLAB9Du5qpG/qk6Zo3xbrci
d5rTZ67pku3JHDaiX15AhTmUETnhdVi80JfKD2yj01vB4R4O28IJ+DbZyQgt3QW+
8+denrhnwUl6udd7NZYJaCJSeydXfJz43raHfPK6H2ywQE6v6nnokrrTeGJf0T8M
qiTM4ExdzdHIfz7L46XvnVwY16Gg8KFvPJLrPOtskKeUg2uABzcI4t8GNgMTt1H7
Ro6rIOO6F7nrdsoD1Lip02daZLP3akx17euKmpbQWXlz5qk3BXRzEbxwV89v68P8
Ljc08EZLzLVuKeP4KSc1SvyNtGCj4AqRSTeOpAggM1Fv+4IVnU3o6Nwqz1Fknhei
CgrBPFQ5A0uQSaTokuqmX/K/aZe5r5+vPmD6nBTFRo9gImhXE94s8h5STDB015DP
EZPQphNiahlq1XdDDn+EiPJMDW2RELkzfUESZrA88oPJp6/o/ruXnRepB41MXt4f
DN7eszqjVT9VML6NLmnG8qdWJyWMH/TxegrxSgFMw3M9OZM86AqQL4dX/P65uaPh
zYxYkpKqtnlxAkXh+IzaMOiD7aI4U+Fw1GapXShCIQJ4bXxcAI/RbMoDxIePRiy2
9S2wx0aiCCEvXbDWCl3V1eD9LKH8UKGB3HQrLj4MEnGq/yzHL7uy/QeVGUTMAAue
EEBwcgdvD9r+r/ArZXq8+qCGu5p3QOsyPOZDC6gwJvyZuw8z9TFMTcFaA57RDHKB
CnOQ185gp8Fhihf5cpINKSbw5VqB0ThfMSiqa7SJlkDBrxS00hpJSzLraOdNf4l6
CWxmPNG3bHs5ICE/MV6M6KiSdjnTx+uMav912RQv0Njm9u2QCfqQbO3jFuTP6oaY
4rE+3KDMiurrQCtppErrmpWT7Ly4yg+ZAYCLMgQMsyak+nvjsmhfwMBa/D5AA8JF
ZL8y90JUNc/lvkUJKXPmLfiuQ9ot2masPIsS5C1X1lbFaY/C+wn7Lta5XIa29PFQ
mOddmukodRU7mDDM/Pe3LMYu6fwOD6Xg/kcdIM4iDaAgwadUwHyo5m/OgRBNNYdu
4x+W5tcV9Kt9jt+iVgfQJIP+jrleXRa3ioS1kL+cWlyCyowJuUciPZe8barNcZ+H
YhClre5NeciUKyUSkggpvUFawUQpxtq+ZNYF+FxD2h84drg2CsmGLweOo2o8IF5E
zW3lXqeBEJD4dBSumGfQaKSv2v5WRujXQ/fATV6LR4irW9T++lfy4Pu07QyrZ5Jn
ZH23MhDwNlOGyn3yhB2QMpLpx+keX4HbwOEiiyUJMmBe6jve2BRE7wn/m/sb76cx
bDacnTrLcOia6LKwMgKbhNamI92/eVy1Yq5zh9vdynsBYPIVQT+3TTwa6MPAJ7+f
TWPUePjcu4ZRKMD2i/0iljh8ZFBd3B8XfvHCq9Ld7YR7PwrI6wDy4qkt1dJVsBhU
Kuo/9PxnzdV7ri3++yi9E2HzTTmNN4yvZfW6ncfJOMgiy1zUIZx0pKLCGQuMzNpQ
x06TgwrBhseksZdIFLNE2GonqFAJ0pmdKbQddhBdmT/uHxGavfkmMC/JeCV/k41f
IEjKn/NpbOmOEjuuqTzecDOtf2AmNQ2OeKnExjApnjLMYIyPgQ/UeMOD3T/iSjk+
q7jlOkAEnyRQBwYyHE0u+a6vMniXLx8DRkhLy+fgmnHnTXIGGsue1vArYNi1bXWx
SXcLxNO3tJY6ue0/ZVyjLGr18x9ssYwfdsjpxYUJarIvjedtMGFbAWgVHDSf/1iT
aIU2CfsVTGPO41T+dNDI4f0kXPbGDSLcQrMu0J3CYM3+sJ2HBMySK64yfgGgoVRd
mkV1rSuqOrtP9JNETAPuuXP9lB4jxIwUpbt2grlggUSgOznXqfu8yWv25Uz8n+JG
GAoHC3IvZIZwSx0EDs+WESl/HyAeBaTT8Ra0Q76qKIsqTpuz7EUHisJsvKxdST8g
Sa/Af+MFV9PRpmYyCQpC3upHoPBbeY6jvvhrfs8aIs9lN/9U94LP1eAQaxPjsZlC
Pwop+orxuC+yJU6cyl14SDizqDZwofrdAq5qkw2ZI0exVXc8HryXrqUBM0DqaA8/
dSvE1RqaO4fLbpur2XsE5LcHxn1ui3vwxA/5PejnFuhjmSdHTE+K7HJs8tli9hV2
N+s5ahZgt13O0EZdz7vFz25pdrJ1L78493BKQMmkeCRFu2uHcz4EX4k9Nzj1DQps
t4Uo9krnMDkMo9pmzkEjxv5hgTDDpkpC6L/dOE/ew5ah/WfRjzeR6Dpou5BSS59m
jzQq+rv4Z1iP5rSNLJTjO3QJC1W4DGsoEi8n8LKK/huGJsqT15Ex/bjew2jcJJIo
mmOAdQptwWgf9+lAsIRPVtjugaUOzDcZFFsOQrvNEqF4kuYRkEmyHL/KGB5OcqqP
/MNgdVf857JFzYYysEuqLcrNp6j49lbid4R/gUzFG4CQxObiupE2sMYUSiR1QgER
e31IaYImP4oOj8SCqe7df9Ieiwxn3j5v0DSWbGwtI/g5ZLxqL+tydjmFShZL2sMV
ulPJKhE7pdoh2P7whPglaVn7dbq7ofKIsihI5LovffY0Mmf6qiQGACWhAKn8A2pl
Xfw9vuh8upShVUGcSMCylfbNQGDdv2ZKWGUjxy4EHXdc9I0yvbys5ABIgoh5EQ/m
SF9oPaHCEOBYu/bWDrSOnFoKEyTbxbaDlyEHEF94fdDvlQfSvfh+sZgsz/BOH2ve
Kl8IDRuUsVbXFH37WBTq10EZJZUX2O55UAAiKLjZcpL/usceCTNmcfHPLAfdWHhI
/e4Z2g7DxjNz/4eeCKG2h3N7sM5c4BHRZ2QG4q9A3PCbw6f7Sl0hkqLkdq69b2vs
Lt2ximsTbCqDYHTG+ZZdJ9Oa/8JcoZZdJtqgf7pEmHix+nhOG1JNYPJF0NHUOgs3
rKAwbYoVqqbiRT/N7BUIpcVRzaiVnWoPoSiqgq6wl4KsDMHY/QyMMHvUXZFeIqvH
FPY3zFzk0IWI+zTKUZVybWEN9B5v0nNQOp9r9kKnAJ9vPTTbkir19dQcXBbDaE6p
q5Ve0CLWLsMNtEH1PF908iEXmLRVqOK857drtQZiMZfYaPyaOT4pkggrhr4xMCT/
ihdQJCien7p9CNAbNP8eO4z/JJ1Erm0EXojR7HpMVGKDPKBtmKDkGILUhbfOlh3g
hdcVfSJ2RzKodP6K5DxAsA/8kyRaw4vPlYUwq45X/MDqvWc4MaxV0/i8vGCydeBC
XzgwukU1c2SMkwHN5DIw/0u2wxhYzXvpdPrqEeTYLR1I4FPYNkonSFb6xlkKJNJQ
Qjty+fNwEVT/KN/5o/QIjAsEaRjJPLut9zBGPfA+QzSovKT2YJphmCU4honBPsa+
2ucMbcsHgtNwtJmzk6ohD2CM6mblzQ+rBwm4Vw0ypg92bQk6b5AfnwyOg7Q285AR
95kqU1pVPNzJ73qMhg/sxbfP0LyGrFSDg6d96vCidQPoXNuZmiINAJ+AhewMjDXT
4M0cohwDmqL7AerX++ZlDTbu2gph16InbFQ4WMu3sg0NfwGhkAY26XpLt3cNzxIm
vfKNIh6vxrXgAbzZCJgbzomH0LBo446NxmjdREhcK/q48DrEfD+nUAHvyhrnvQT8
NWhl7bvnNuRJX6oMZoBpUcuuaPl8Qth84LRpVmgOfN9fl+x4ni9FtZah9xNAjqIr
bcL6oh+JIP2SR5a3zKqBzz40w8v7gjvNFVBA2K1bJmhnwX3uHmS+TT+pjDzHsdGg
sCAxn0S4pVBpCaUqzHS30PNoH9aoCvLj+xiLVNUHCOQyhl5Nd86/Hc89LRU5cASs
rEIJ9PQGCtMhtPrM3iRhkkMI+G7VbbtcZWooVaFePDz7HSXRr8Mp7AhX4d4nDNKC
wmvawPm4Ue1roDs6QDHpg0lHQkE9fIrgJJ7X0Wfurt8kMFFMYrORtmCjS/BG0bFW
yHwn5ynvl+UnmWbS2wY0FQUqHLJVihYuMmKIM6RsWHTzqDYgVvZvLYEK7g78mT3r
73t9ydq5+7miZbN+n4BdeMZszLMQMHwj5I2q0X8YmJNgf0RXqxXdDDG2NCHTw8HT
+pRAx/uuQweHZ3cSPJZkxNAGVwoXpMaG9C9YYZ44T8eeQ81sKaQ7cF7eU0GOdpcI
7Rl2fT3hggQrPPLCD/7KQA1Qaz7xP2DssPIcNfT7pAiSQ/utNY/Ju5uEkuaY//Ck
NSakrtU7Exp2gu+qL6BR4BqwgbCqQxblwDorrGvxN3lq4akINerNmBAa8QPIIfEH
SF78TB6qlu6rEEVqp0iFqdb/GXgjtrhMQurRUjxpuNXD0dogV/ktghH9wxf2OmgL
5PGI/A3h6/45DBPYgfmw5vDpNg2+Gq5siO+Op+fLjlwd81IgxuGR7JDrIjBPWPZk
oPiBRXgGHaJZIcZrw8xbRJ+mNJ7TgyTZl0VzFhZDb+WwvYsBl9i42+snLLI6YEUt
Y7zNEo6zjAWa6R2T3Amwxri3nrTS75JyfR0f4HQAsXypWEG3yz+DWKK928+WxhPP
0qbcR3ym66V6f0OL9R+aO8kTEQ3f0+AvoiRyMfHp8WWrS9+Y+SVgS+0Ub64/G/BM
r2YuDpdtvk0ddVyGwOH06TqwEb5vKPFfZYSiPG4jeDaLDXfdDadcHkYZ9h27Y2Td
ZJakK+Kp+I+BrEbL3ujf+iI81MiMSQsvpKQ8ItJ/6+j5o3i0so+kUY8L0vnBmPeN
YYLzYiOuJD/IrIBMCa2ztsYVK3WoE9z5NuoZpWaVpYI0f5duQLGd7o0mV3ElbHgE
ZYBpnN4qhIk9E78kbmPI2O8AxClEbplJocQzhIMlcsiZdtbriHTv+VoxC1pdI4ID
6YhjAHzE3IGQzL1xWXg6GWwQL+Id2uZIsR3YXxmaxe6Q8BHiaWRjKi1HW2k7U8At
dD1zVmnHQIf+YXREbTgHI11X5QAJcDqPy+FFR0yFu6JberM4KuZxbQC22GD8WLat
4PNXima3XgavPdJCZi395UopA/Jb+l04FCVAROEzA2UWCK3Hyx3aFidElfEdcdRr
xKsPqpGZ1+Lurr+OfNJ8+2RkYUZ8wyQ7LjP4KWIxOAzX1NAP/KhGteWm4L6FmXT7
yfpMr62uqYb+qwK3qt9+3S5qlxxgmRIYX7IJ7lRXNkq7PZ3gA2Q9FCNRZwBCNnoA
bSAeuHrco3LMOpLsh7AWhp835vi281TlIGB/9sMIBEa6Wkd4O7pdtI6pX7wvRl1r
r8fRELfPmA8uFHYwjfxit2Ny484Q5W6/pfDnow7xydVN7Ce/E4oFFlKkX2Olt5l9
Srvx3djkRAig73+i9usICk893urHSlTFcybIygbNOKme3Bo/0Rbej2x6YbT9n9Ht
6vPGzMFxC5wFbK23BUdxL96mB5CFBrmtF+YHE8lHeqWWqitKGAhG2g65oYK9Z7xl
5sN8kwwkmwYvGMjQEKE88diG+ehS0mOPPhrYYXSyOMGYjIEjzgp9M7UbDOFuZmSI
KtluF3r+BYSN42BfO15Undy2/iQbzin09jtX3MhBeh0bMXH6+kUhT2OsfB2CKhlS
Z2v0bpDAjgmgBiZS1HjMJzr+dN3TIPizfrfm+ZM/wgCQNLmEaF/6grMUjfLB3DUj
VRUdGtEzMRE9un/9zckf2WfOj4KF7RmuzmjJkbBWtcZs1Ce4H6kPUJgpE8k4DujA
tMr0UD4UKsqvN/OyRVNRZnDJjZwm8e92swYI5SA2ILT+KiJMDI2QMKpBH4fjKs66
f70FiN8rCyg6qP+p6mOMvCPtXyrxGIhL5aLL5FGMHz96OtJDv7gV5+xAhOe12j4b
dgw6DtcpCOfVBlX7Xs5PoXp0tsgZ7c8hNZTjUrpFwBUpxhnpe1TbjqaaCjB1RUOU
4dNY7JKBAVShrbVBv3p7lJwxQGHLIRFFco5kLw+5NbCZ4DGQpzYxRnNAuLkBABdM
xt1NmXcCbQ0MyRZl4tAxHtqqOsbXPRMwYc1+glgRuN72gqYhIqZNWTF3U6rnjmRm
jrBKoQTDCt+u2kCV/k+//Qjp8hDNRWIf9IyQcXEr5kD7SS/eXy/joBYEpINN5Vq5
p8boKk8kpYEPGv4If1xeEeQdKF87xTNYAZFD9Yu97nZq9n/ZTRLjtijHELQFY6yG
E8JUxw5qaztGauE2parKT7XYiUX0xbpJVIv/eX+FwwAi3qLBid4tE9sQ87FCmuVK
rkZvPw+AoeyNyMB69AU9sXa2QvO5w4FCJb2RDd28Uv2iN7QouxBIK97Y6d2i9wxl
Q1ZEQwnJDt3UOiEwHnsa1VGxaXLtUBvT+2ap1gqTJXVFv2y4tg4gbAw5PsGWEpz/
0o4908AFUU/3Wg8RwYNpzzDEPX5O48v2saxfPnvuG8tm5edXfGIggL2Zx8209zwl
evZHz3gDdy7I6PquPJeKAlT/NkBnIfn2ptcKVEx9LfCK8N//rRDetQZT3Hqg1KXv
6+XNBb9T2KnBtmGbosEpL1CXSBp3KK2tA5FMR8jV/HFkqWU5LgWgr9fEOoCnkrVX
R8RQTVh8qebHL7u8oEkCkAahWLyFPTP8UQIBTxeqW3oq4JcDfmvcks6FyBHVpALL
Jsw+Y+aF45bxZ1cXu6Q77rqYniXVFQdRyHpHs4DbN7EidLr1ylBlQw2G7R2PWdP7
+HHAeRXSAoN7Evb9A66GEYEAYJpx3DgVMajg7HjDYqHLO00mGv3tdu+vnXUHzmRy
MGPIP4hvRctBWPXFJXd6/brJJ0e6zNLgXYyRzZ02xlkco4FVbqrBUrc2VKS0dwDC
ytaxNSUOspDFHvNtKf0aRasq28Ttn71NXrt6X9YZ73a7hWq4PQq1m/ENDjctuW9r
ENn5EwPEHwUj3+X25pgeWibZiY9Hvtxn2067To5QVLQrFziP3gYgckgR1TVOVTc1
Iz1sMSn7iRLlOTtSGskFXpvOK1CmOY2nakx2W/ZQj3/f6+EhadHsJwmp7pelzz+M
tIivEnjRCyAMrrfF8OJunCGTU8oh0fadtslumUT173v3H8ugjdbzs/a1jQFh5Du/
zmp5ycTz/hzOU8kfOUF0bcSsMtnYHDYX8ssIhGMma3+2Tsnd388FGs8fuMj0jbmA
SguWXPerilQ4M7RBHUnj8pyi1DDiQfBWBY/w1lPm18REQCUj0ucjKC75lVorW9+A
6EqiDTSKXM7jxe27H+a9RJf0eDdvLhD4qm4C0aMUYzffogVGLezKaPKeCWbNFKBU
MXrOzaFSw77LjTj8cfvruFblsCZVWZ8fGabIW1JRgd15bYcrN6QDdkfJa/VObShQ
CK9/bTmyGL6D4HslwlJAmM/lpecjf/5l0vDdI16ISDq3/bn2ht29jb/xnJ3UFxEk
8TyuFLfskdNagQC2b9eyW/zp/M1ktO7zW7PgTheTJDUygAkd64JyQ1zwAhM6EE9w
6NmMfCFwryMz0rpvw2U+diTTopFX9ptkdWWIz1t7CxEmMFjvMMCc1zbXE9HHqKqi
s8/qDs1tgLKflfUrP3Hzo+ZpT3t+4X+ATTeW+UPrKWqNYIZlQXA1fXYZUGuN75qF
dh5OrbCk7ZvAGSQHH2JtCLrGVfTUI8hNtTc6cmf4uiqSj6k/VGKLArBiYnErmGAS
V09kgt3dsx7u+J4FfMZJJRa6leO7cuKgq6E5unIo6VhKGL++hLWd0zC+abooxMFj
GjthAZFJxqoG0+ygmFDLMcedHbykZHZyLIFno8nY+bzw0CvZQheiyewDQ39vAZyr
UXXflKp2ak30AD0mqEKE6mqKVoQhAdiRGrZEC+Z9dYArO8jbbmSJupOJBqFCwiRc
Ge6gFi4DyknM0KTRTnHi/U7lZhf53FsGoKz8z4uodZeNyuAzUPbQEYocXXuWkz7H
cq8BgBnleOy2zrgvCBArAiu/VO2Du80u+pszuksWtGGbLQRUP7/GpRRjX9+Wv1Zl
4HYplPifq6icwCtz0+nmj/lYIH4c1AqvBKAittY+3vDCmKhBZGdCwNTYnBXRQB7w
XXMaqynWTk4v5AstI6KWdjhXcWfZW96fW1lQxT1sRXBjUvClMvYNKFJYeSXGwspn
VNYqdBA8dEIlbRkIEOgahWNXnAe5KRhT2ncZryc06PC5GJI8IIGH4RKJjOMgmXgW
LScvWTbcxG3KaKaP4bYfLiOGpYlLlcXW+xpdOA5k+Z7XvVcUq9YaRNJ55lvW9Bau
orWZ9maVYokkqEf2OkTCsxT14qtOTiQzUj/yjJgAWQ8hdmxIo9LRq+FvyQlptxmw
WUJtzcl+QLYClsAvU54LfATGSURABrDGZUYMIGAqRrteXCQV72akj0pvpnjKSx0H
CyvjDTDRIBJj4RaIl0W9/0LMSqazRd5IUyh1/NAezRmKXqz5EdGWSXNfHbOODXyv
p1UcKY5vDdka+ZO2jSZEweLERD95yd/TdGe2iJrURF3MWNGAAprslT3pJcwWICrl
OwO+EVTJBrQ2yWUnyhHLqCD/heJV/3h/SZCYwXn5RJAYpqMW6iprx5uwHDbKlJjj
fr5CyFH7owv2H8rMHwxwkaorZohfXByGsVaYd4ER00CTmy0n81ygnH/lwIF8d8EV
v4AThR8t2nmtzoVT26NgjOmqjGia1S+YsWSu5b/Tb8U2loJSZ2ewJqx/QQ2XchNE
8xj0DAQZp0eHutZJEijZfqR6CB6cHiHE5jEPthwXRK3cZGt64gosw24Rw8WnoS+X
LGvK3PEI7zEbiivKaUHmKM6Kia9K/rCUxh4xezc7TRmjjqEhJA3pzYQ8PUSFGJEn
LcitNww1IUNWf2eUIHBNYg1Vx5tjJSEo4y9087vvMQUnIyD97ZIljCX8N5dA23/5
h3u7UJWuQ6yC0nwfuBhuzNfkKqri17E2BB2WWCnxOOpCJvjA0j2RM4bTNDGwAy+a
1NYBBDIh7QsA0PwjsI5yVzJyKYbvhyjhWUuqpz/hHL4P0KTKFKGTL+cT1y+Kf3AE
Mt2qove93qa7o/am+32TBaxtaRr2rxotMCN0jass/qdg6kZeTNrzU8PT3lNwDJEr
YRW2hIoA0bl1nRBZl3IJkYLZnirS8pttD3XJtolEZsds4Qr7DCXZjIjP/oRjtHgt
yH8ev7zcw54LBG65BnGtoBYXtQEHsf4OPYS5ZB96+/7Zc/xUkLOvrRgyC35Lfv3o
c5mM/gSgGBpFkcW3xcNVyEhTwsZrtdp1uPLhdffE7EOQmwzjE+epEyXtD5MZwCwO
Q60oyjLeNZyLiLdiLpsHmCeBaJjvmdd2cfyIuhTAQVqL9RlvFCKy56FmhbuvNmWk
8fr2HPc81k7TA4IWXXrREK5SZ1Uk8MAUXCndpQYjpT37zF5kiTi8LwfSrQqMtb+u
NW3uC6i0WJPwRgrH/QNomD8DPNgEEkdf/kHA5RYHpoFW2rMxVLSg/AE5G4D0ZyMu
NGgd6BO6EBeQNB6gan3xcXucdd7UfZRIc7F/c+7KGLwS+jpE1qsOaLasJtRRw/4/
v4MUDX+MPVgLAF0LHTke6X7WuA0Bvj1gEdl/p+XuB8SdUuV0Uhfr4fPUzX0ladRr
RBQ/t/aFbco7hSUcCSJaY9lTFG6lVXq0VssVpqyNKgMLOyObeMM6OGJnI/UGjLQ9
5z8pHTzIwX/4EHQE9lq+vfrAN3V6xSqYX577B2lxavJcZKcj8XO7N8uiXUv9DN2G
LXW1L5EV1OmhF3W90hmMIdlVp9Xmpuh43Vl2BqQggiiU6csE4BCAnanwdisqY7Pt
ThvGr2TWAUm3gBLqBgwZa/PFvhDeQTNOe1mkrNzzANpauJl0yIZMUImTp01eRSEG
ihCKR77kJOFHZ1xh3QTC3Yu2Spv0eOOc13b88kZGW4DB7WSDaOOf9psSPOM4TE0h
BNsZ3/01JLwWnEKBTAx7BYtu1dN0ZGZcUl/Qc5XU7t6IfUMEOowp5vY4aFDNH/21
Rrbo/f96sqjThHQ2VGbrEvXXffE0JFRsHLhZWTgMQy5Z7/sNEqS1+BHf6kZLoEY7
kOdzGOuvFWykv6w5qPZqX3jcitxlpcnR7Xnwq2vdQXRMHJ58JELz7tYrszkk2EVL
E7ip5geirvXIswwk1chdzG//Ed7MjuAHroHdSGqh2Ae4Q8ET5XMVXBqxR/hBsZK2
bIq0JjfmZdpFGoll3TI5O7E0fWi0v7kDd+OSUzbTzxyqwnXtskOG9VrfymdbX/ZD
Y2VJajjb+oHcfUsOuM2xY1nwcXH+mZsOK+RNEIe4HMdH0Kgv05tTg1uJUvm6QP6t
8Ifeb6KTcELRxy3tTJZoVJ5egqn/OVkEycCFSOxFLoNtv0TCcxeiuOIqWbjLarRy
ZuvLk/v+qmPhK1I2g8MiKWVPAZ6GuNZ2/Q8/z15OxszuX6yo19kOAmCMq32sOdUx
nHmWWXyuRVFOnS0Dng3hvq2PASJUcUrdp8IN9BNMV4MjBOiUrRAb03Q7vRN7f/ns
gApW/UHkBHwdOCs/MB8GtyWTNuBP4Ne1DN8QBoSfbSZ6A0ZIg8wIiIRb5A3Fx6E/
Fnkl9n6/J/T0kNYaakG5KmjYJ8y/7KJXNrjs5miTlKYu42UsU0as2qfrQVIr+Afh
umzuiWyqJn2VE//h+nJXV10LOfAM77oP/CXlhPh6QzH9chdbR0p8UWqNdlFt926T
SROCiDH3nofMXtZjWJ/wgispqeZm8gRnDVzMO/Qx17MuG35Vi+mPBVDYQEKB6I2z
5bOP8zVIHFqXINaNA6g2Pcc5tKnHvZXtg2kc5gbqRtVo874QEBSZCGidUG4fG0Nd
Km8uyKL1lFVsqkdHoW9kkC8/a+olm7giVBSgcIOmCmiJPQRUWeccTo3Qdivg1UUQ
OsUTX+GjCtbY+zgT/OJY+EkA+NUJvuCvOTIrE4o6G+yjFfUrN8pX3e2hIB0qE591
aRvim97aqDaBfxys5KRixbErRUt0+avn7JEfb5WTK+uSi5gG/mTXcs+dIo0X7o8j
S7YkRI8dPaDWYthe2zVeNMwc6AFB9mAKvxLa+Sp+yaLZVolsdK+CRum2kWUbV0Ur
ir35b4B0HWuj8b22S/D2RWcDpLrtot2hjU+1TmdZ/Y7DrXlLSSBgBZwaq8RGGTc3
WuzFM3DezAGYfeAt9Wl8JBvxmFfAB1g+9bit1zltsmeftY8cmsblNUa3968YYyoV
QHqtEe+I7oPukQBuc+XC6zeVUOuSFwQHoXxv7JqMaU8IWrLJbbIZZHgyYTbRuwKp
Uk7cUKMW0pYWriv2j8E7BwoMkn7OLFmKz/zmOcfupWsEM7rhief0DPrYe9EzJZYO
MLoWtnyvzUz8778M9fTVdLTh503nO5uS98vtpfvAfZN257/lB78UoVCKbkl1lTrM
UYsXGiDnO0aSwgAFfGKUexZ5FKpUJj5ryBNU10VBypxpFvwcj+mCrajzlL9RYgU/
zsgNrnuF7Olc5SCxHLuIAV1lWz9g5S93RN9t0/iFqu/wPwdZBe/bF+HByiy5TzvT
E74hAzh1aITHS1nhYHftxF7DgyR3OjMfRmfhTreD3DAqh9/3RXz6s3E1fz3bUX4t
z9rjzsdll3oSDjZV8z9I8by7ToENHaMCs61ZEC4tydxPhjEG1RzIAbRCdg0ze8KA
E+32RwMqULAkH+AUMwsiwKmxx3xj28j6nrjHCp0UzgMIJlrVkwxN2Jb/4FY877C/
dp8jXDsS2xp7L1UUYI+A8i2FvOmdiPA7Ma4mvF5tAqMCSyOm8ECs55kG5XzRubo7
OczGsdB1EfwPjI7lrdwutEV4JdknP48v0QX92EO4sYbWXg0R+nm2CjULRaHfZrSv
OaEuxTl4SVvw6BW1LQA51qbpTbDPQ9R/+LLjcQMiIO4cj/VdSo+d1Eb/RVgfrPXQ
rjhOArevC1yeH1KJab4fIHvJor4DeNzprKQLj0L7UO3akzrqNy+KyznnuTITNRXP
Adt/wHKTHgA3Si7ZnPLDBxUg6/vqsXuTShP5t8NG40mKV+ygXJcHbj0m+tpsLaxt
ZedhYAMNiyJXhDYwrlTIFQaFR3GFjqx+8ye4BA3eWuf6K0PHIVaBFb+KrGqjqv7A
NgbxjkraFuP8iH3xE5ezevcI8I7DL51Ibl/VuMJgUkvipeqrCkJ2RgK0qCnZP55M
xf51boafsWYzFmUAVsORmhAchpMRtLEHx/HBzGhGGZwb6vPVmWajdnIkjFL6G9l0
OUTKZxUk3If6BLYudR607gft96SRmVxC4WyHwmEa5g2BiUyRUKzq+AHVn1zsT2JT
t7wX8VnWvTegLWmWJKFdBJ+TSeocKyIIO8kZZuSbk2LvU8NEtw5QWVGJV0iStmly
3maEAc6bFvyPt3n+642rRs6KmxGdMxg4guFa01EsCloYW1KQjG3Y0Sw3/dg1/tsM
rTb1HQu7qD+qrMmZ5qjJGbkGew978VxEjz2Y3BCPu+2+JFtqsij6v/PWQmGtXKDW
QdJiHHhWD845DJzhLoOJVxECQV3kWvj6f/7VHck9iIKG5aXtD4koMiIJKQxrk7vg
7xovZyGNWY29IS69qBWBGlfDTu5uIMjlwZKDOp57PU9itbeUgYXQEJkD7hA51O7g
NJLCyEZqEpP5drX61w6ojuqFYzw8HTPexgvhqHOdLCJ6OU4/gGtsWZ9XtniG6K7Q
rlGzqIjyIgbnbgXTJ8DRpRBbrcpVMXDKFRQ2WLxZs5ZBJGtr4BuwnB36W5Q+M0jx
7T5HT9ryH6f2JJHbpDpEQncinqJRi6aqE8XPWALZLkobkcVtBL6UrLfdUHQr6ro2
Fo7JSeYEQR5A+RZinG6yj1Zk3ZGiwkJuGHr2BSI81tOBSYJBFv7AiKHSFhjRLRYG
nzyAiG0nKBiq0tsVfnFltfKO4fUyNwovZ4OaxdltNFjyckYCeCDUYs7E3QI9gqRR
Q4vktP9nKYKgM12cBKP4mXrTCHcnI+ZWlHhzoY0vtBjPn02qWmid64ugQRBTE+MP
yQhk7zzqhqWpjFGJ/gBCQeUsm7JRTBX/bxGHNcWeUh6G54q3zx3eAenO8JoPL8eg
sjdkHPup4V/G//FRlRxvDbtYQLLu8GoeaVys90CDaCcVzwvBlZis3Q/t4SrNLWp0
nVES5WAcHW0hfxoDh3W1u0pZhK4d1Mu0vUW7UsCrKxhrQrNf41G5h3tqqkhA947H
/cLdN7tn/AGmhq7VD2OimgICCeeMBKuJVSwNa4RB5sJPYoeZRAf9F60J+o66WyBf
xYiE3ePAOWZ1lEMsr9YT/F07vic0ZrYFnzzbrPSMXi7gqkmgqVcah6w7ZheC6+Kk
HfDBY9K5VCsbQUV+RLrkEDjilVtcQh/RrmEisYbSxbV+9Enl5QL/Hzwl0hpsnsb0
sfR7svY9Zg+N9ipXBx8dQaL08OO+Sle2NqoI2AwlXZsyd201QyH/tAuJVLWKrXpd
C2G88JvtZjxa6HL09pBEUu+S4d+lwjjju1UQirvVBs4cuDHnBa5Xp9cHOMhj9szz
OuQnd4C3eia9BfSh/jD0hBpoUCKFFbAawdUg2zkoLGb7nF53KMptSMTPXh3ol4k4
u/sv4pvzdgGRbVgKqu2i51yuICRHgIW5a9VrxbhG8V7dGx5rBAGDyYRm3Czzwm+P
iGozjCCdyjwXCu6+jkGtETlesszaHZsCas2N6O9le9kXogh4MYsXebOymbrZ7rBn
bpbZS55IvKnsK/iBR9XZZROKEfgW6zdjeEuw+3ctSF0MEQxMjNhj0Xh7faN/IcVg
AC57Zzm4PsMw0712J8HLdrZSDSOIcZmqGjfgnWARTmKvnDXmUBhWLEx/iRlS778l
GSMGM88Agz0QrT9Jh4/uYi3788+aWXLpMJH953/wyNZGZ5qCDVAYoofANG42va8b
b0dPXDWzkbS5ZuKUu2U3uRSeqpqa4nvopukZrUV4mJxjE1CGLz0PYAKm6lEuNY67
3M94q9utwWAyrpYA8LIKJJqtUTV5zuZi/+JpDk+TnfRcPjcBEXci952Y09kKyKcG
KkojzjLKBDejoSSfAilOww1pr03HAj8vhdP78AO4ZISCM6KGOMZ4++lEogagOR+p
QM11BZCCmJhC+I1LYz3OirIf2u8Gf3HSwY5mrz6TDT//F6Nb//+25RYccD5OQPoF
lVnYntWKms/9o00yKFVS3k/+4fEMQ13/jJfo8D0Tn1MTIH7FLe05Q+o49pfJMRVR
kRG7J9g4pc07eCjlcAC0dHmy8drrlYpbEODIzbWDAtw+TrSR47uYpJK41BF0gPtp
R+g+EQrOwyicRqxNg5wsvRuE4swlzSda65XkO+eL/BHNMJ/xRXrdtJre41NaDAvq
FvXv004VGXOWi5ZB6VSs/Q8sIPKTJDtMqasr9wh8oLDLBphaQmMbmMT31lLdy+0d
VCHhCD6kqwdWCLdnoiNO89baQJWw8x4F+6XI28MSWbzMx/gBpNwSuLzugRJ0KVym
OBJ8ihKk3QGlSl9qEaCPmCxLTGeEx9txAJnJNktW3/eAjUcu8xLMZa3/Er2GurUm
oRxRUMhPzHd/yYw7vWDiEJekFcTMxOAd332LrS0eoPi+I/NvNQkokcfqiJS6bySJ
CegaPkr1Z7c05e5hS3Otp0q8GFV/06h3R9XyuE57JYpL8rn/KDPa5V84YuNwjdUc
a0qbQ/jqBSvpQ8NU/0e5YgQZB+/v4rbkQqiYSNUh8OROpmN/HugcrqD+545pVFyE
f19mGTOnJnSalgYr3SAdNaFCg5FJ4yl2x1P8gmHEwRX/ZKv9m9Fzy467uKJ/GdOW
qaHNvB9nmA6n+dAX15DGuXsUywmJ8FD1+GzzidIqST9whERNlngBt8F3QFxNbqX9
P99nUkUwVVPda3VhKWX5w/lzmWGHblrTldEC7DPCZdeh4rWs5bmXdo4tY4fxj/xo
6TGjyTyiQy7ZzXl9TEZRw6wTWD53IhmKeTix+XI+ggj0d0S9PjUgXgVeS9sKP+46
RmQiSsfu1Ci2MSDlNkyhBmJTW7zvO/2jcm2CnLTd4hpf6uaOK3yhTw7ge7Rl6tNy
QeHncLXi+Qnj5NU4MfAfUQqItNEkvzAzE15A5wGVU44cZagsJizJrmNUmwiFRfjS
SL98CxusvDog+bHj1dxezvq9eWr0U4a4OqdmkL+rP2Ocl6PKIsHYB++jR+U8dzht
6JwDUuMD3+zvG/6QYhzaXAK54DOv/R/j4aIh/7Vv6kRD4eltl5hM1hPXAdTA+YfW
4kssWIbHSOZzVR6dCMCerWUkAupauF1XYtXpFk4ZnxPIBJyBRgGKs0znt6i8X82d
2YyEEGu+PMiN2zeqzTXa6BpIhBl9x7lLIeE/bT7YZtDEX0ExZvxjY7P8apHuart+
y53Yk/B6G+xj78AiC3sBZbb5Ht6XqFsAjCw2m6gKwuG5l/jL9eO7KaRlUgzWYQig
FhhDsZ1mAf3o0T5U9q012hMfiNHt0/CGjdU/jqkZBDvqmjncorhm3JbkrEBhqlQR
orXla3f+OVNsfC5ls/dttiQ64y1u2oBzw+oJHTBQnSc1oPSF4U3OgLgf+LBJqURi
ec88mbbJT9BsJkuhSd9q0trID/SQUk5z96XfJu42KY+OymgjD2tgTb7VsE28GQ7q
a+xC+xPdnAj0iWldAplGNUCrxWnW4LAWnSqw+3Zu1+KGaV6d69LJNaxXwZrzmGlY
MXQIkcHbO6ypb8ejsKV3UGYJtfb4LpbmBvMgZcrD+IDg1bgMF0Cm6TfVTaBxnd8H
qMYpjMo6DOtk1sso62nq06LeIpAKbNQc64Sjki3A61lPblNFvWH0U36b1I6o6NWM
VqP9NBaDsKqsq59JJElX473+svK/2o4AgLmG68wG6Y0PAbXssprohIoEsV/F+PSp
pdQmTTOp4sGF0b1WGpyrXXtNSzWy6q9U/Ve9d/T1BxOUlm6dAK8QCkuQ4Lb+R50W
gN5cVunUTrGjc3XB93BzA9/c9v18gSZd6+VUoQbikOOWUuRzM/NcjudGBL7PhqX6
XjZ7qHbeGGMBzoZVYqQpPAzf9QBzW0RVgbXbYBs/+0XSuGcIQqBl5+t20e9yxSPA
BF3x1bje1wMDGl63RUq2Gnt2J51jSALnmaSiGqv6aS1XwenLNy7PrspE3wypKS/X
7UXc2p2wLe2mZxyjOhY/UWtI5+mDpNWfZOG92ovthY8Ue7/04n4OZ5SqDzkv5cIG
t+y+of6XwA5MDda4uW791Dzj9cLjQSQ2DutKCeYf9KGb1JDtN5M4+evLF5LtgKUU
PYB1x5LBOVbI7XtMvm4PDbXlskxkFNacCmfOCu2DvVr0lingGQXhQk6lWaYqZK7o
LyrH/fvWOPm8tyIficFhIFEjtzDIZ4pWUJLs+RB/xUKa5oBLex40haIzSoE/yaH9
FCFIlMVdP9CSylpTwyk4B/LdIfObuk6OLvyFqh1BKZgZV15pvg7vkI8WaZoqUl57
HzF2q01kLWSEJP0Oj5IbVRxDPdNkeOjy3eT38x8lwEmKKv6NAeh8rMuSS0+PthL/
oXh2uDCd5J9PlcMtLSuBVjrM2vy+o9FPAivnbDDSLiZT8+U9QbwXK6IIy9iZUq5J
jRX8D/b/n7c7VCQqvKXpmTF0o+4fwuo/6GjeL0xhrCSB/fBxPx9omv4hdYP5RQFO
sP/Xy8Y3Moyc9hFzoFYpxEDp4BexuVR9O8zzG2rqCt00m96Vr4aUI5ab4bJ5QiTf
50ktGpg9cn5UCwXWi7aB/86a7C9uTj8AZJcS01jsGogYDbBsG6tuKVOW4Sbii4/0
9lvhI+yhSdqOxtx8Q23wTm9DUynJ0RTIT/3mnMY5fJL5xjCli4s36aoRlYfWYmIT
6NFb48q59X9b9UA6Tz5f8p1lnleAHQjAARDEsWFO0VMoi7CPTDy/fGnQpud3KdDb
xpU6WX+ywX/n9mSyEmFQmvHSS1l9RaSayiTjxmI6SpijcOQWl3pw98NokEZ5/d/c
RRYZsTvK6DDg2jSHbtqLsTYyyphiNNpkE4XGsVwCkMeUtc8ru1Od2bD/ImVBoEvj
5508C8Yomb0NcYmG97O66o4vM9gOpvqT0S/az3GJqVPXcFVXJk3xfpgm4UfePUji
VQj2YO90d2Ey5VNKYKqy4Ne8lLkM3hbNVHmRZJ4w/SEHtuHU6ilm5RC+Yphir2PR
Gp4sEmhDiWlNC6SQ8rY6IaFayd0PJr0RVGfFLRNbzC2F6WEEDbEqpZiXsdAsMImk
aR7YFbjYnw8NN6nyM2zCy86eYYm+gc5OJu5EDiRYDhlKRzEowXHB7b4UE0L6LpE3
kAe08fNircx8GbEoDCrXa+YUrCmmAMEoXM+17C4mW8TNEsXFs8prjiqb/pQ2+AMO
znGnBs3qixXybZ/+3Zj1anZiXZO7nqgDBgg2/w5fKeV88IONs/eeCQULTOS7Hges
NOvQTypZL+eQ5dGw2B1Tjug9Xgy7FkWkrEPIGgFTwvic4nH4O5/l8lOREry56nRR
cAkCfRBk8Ykl2v2w2Rq1Gx69NeeVgd0xtSRSrUaIpiOQs9wORoOp2h1MH/JtYBa2
yhuA+kX4P0uZuUzAbGOrU8fsvrO5LSJyURsL5OEabWgopLxvfJv5NTM8TNq8hHdM
Q4fqdEw7aAB5T1F2EcAnbHuzWn+Pr0AR5TB/vINxfanjLF9WCIp6SHnqkLgz/kHQ
zM2sHjElrSh59GELzfGVuX8ZeWgBC+uJs20tUne0iucQTh4i4O83eogm15yFJr7T
wIl3gAiUCDl2QbW8kL5gk9OabC2ugaqiDLF0aIv3Pj8JeDd1snWElBpds7lj8J+p
iQRwAwVQzgabBXYn9SQ/F72rDvh828umNNPDtCZDb01luIGFhigW9BeZGGtoaJuv
bXLaRBZxybTBP0IzWrPaog89ZdDcJxoQ9nL07QAWtuFUxFhs1QQYVAXHDejcyovd
EEVRgMNV4MlQbJeFBfvATS4zgydK3gDZ5V5i7Ogx404jXnVTExWRm5R6vp0ppfBn
VJ1ljGptDC7cen2vLqhxHRGv0BVhAqTNSz7QNCDW4FK/Lwj72SZ7Vbswgblo2bAN
Xy/zJ+C+zQsKcoNegZC/+iEBSzBPcJPgI08n5kdIf1dhSPOF0Do1waeAL90AeYR+
i5HKPuxUX+vrUp0CqX76hW3txemTFXC0LQZQSJl8uLtK4NVVspWksfj2QIkGRZ5E
MHXErgbu+UZyxwWw9VooW7QsT95fUQmJLOYHMD9y1nWPa4kO3Z8C5/Yhpth33l0W
rhKFb5hLxqrL1t8Fg9Fw0xhHo0w9x8LYeH/YUadYU/OnXOoxPDfaDm55IPf/yLbW
Td2ns4oTQjg9czB6YMm9QmCw3FNY9aPAKH6hgJRJqsvKjKlf4y2l/G7Sl53MGb3q
waCrTk8+WO/ocK6XSppN5keRKXpZMxCPZyIWIS6+43cCib6YrWOBaLZZBu5N/6Jn
xO4plyUbWoKTFC55rEiqVnETzAkla0wGgqn7dliiwg22bEu4Soa++M0K+ppwlP9C
mp4M6q7seBrX7o8dfReXip86PphQLA+ErOrlWE5z3PmRGkcr+op+g4Te9/B9QcuU
47PT8N/SBwFgC8ihLS0qgNllblXfrctLm+tlJs4npSwoWKxnAxf5DDV2k1qN6rW9
IPZKnypNkPIFuEIr6OpQzBU/JeB0snvSgPzaJRJyVv1u7UWVwzOVZTw3vS1mi27V
y8ZDzfjdU70ZXH8ueR3GNuTibEAVO+T7so9gLyuSs/wn6/2Vj//YgabC5q10RjUT
0WbWgpM/iDWnNHc1vjbMQ8CoRgRNssPYVm+FBJMPS+4nAQVwDe9GcopOo27pvRlD
aW/G6aUxwwjqQHkkTeui4WX8wTT4nvU+EVkBH/Y0aOpPwkilQXVrPsgU6GozAl7Q
u2iss6IW3C/OE/1ZwlNcoQDkyJDzzLrI6j+Ov4G+EyvxL8Oq98vVqFmg1t5UCcfO
4Wg0cil8QCMtlnW7X1zd19yLT7mnbonX9WhhMQVRWz+KMI4Am26C2ZaubxnvFfhE
sqielY7RSzryMH201f8hgNI6RhTzqLjlDFNtCJQUNrB5qEcwJMfG54CBeA5ALbW9
GyugIDMBsaca8+pwvQo9oOTpoEEW2e6R8csQvMbDMDeU6b+5PJ8Ps1tNYFFPyppu
xb00APJL7lE+0NHdiRIGBAo1mkdYGasWMqszpWwBE3CmfmOmBaTDTEOckpjCn0kH
xmM1GUi2XX8/FxXLkdigGcKrCjDwMwLW4jBDTVft4fm+Dvwr0EkpvU+9OULakMnk
u1jntQZ6t996SzE9vtKSeoIdGy+2JiCRo2jcvY/4ZFoAl/Lrzc3sF37ihDS8tFmq
/nCYt0q5TrDgSEHu5Il7+rWuqUuXaYZgzRd6zV5WeedWbqMfukb9a9ikGZd2tfYF
f3SeUZgQGcnvMI7V9h3WzcEQtdRvxoAcrVNGv56VK7IhidkyhBcUB9cXucfLlg6b
51kYCEejfmlgtl+ezkmrf716sy4YKVnCxVjZugHCOuGu4V5EcEN6vXOyL8hyyebF
cRR2TcKqokidyHaW2pUGeBxJqXAMl0WkerwFndf63VFYftl4Y8QcdZN6gr6O5CXt
nFgsxyn2024Tp4uHZRDz51gtkPO0XCIrpmKLTmtuvQ4yt0GuvcQL9eAXB4Hz9I7y
aKy8OsSUzGR39Vq6/knoCCfxsCHxTIkYGj1xtgx9WRjhxvcQqsDNDWKGwNs1YCUo
r6CYbVUxFO4+cj3kWk7WTNCZ/Yr5xjOocjmCaljWlBdapZuCn5WJZbCPGbQmDTTx
a481P8GqJSm9rMi2IFz9dpJJA1JUkzPgcKBHoc+ox3DrHtUpf0chA7B7rJZPEgBd
obTKP8DTvY1T+/QDcGJNXB5r8ZhTdc1q4b19Q5pOEZ1w3VeLPG6g5lND3KV7bezh
C+/LCjFnTyFPOsvHsKvKxhWdGIRcnxZKSL5rBla4qaSwkkTSEeuwDn3gbDT7d8uI
9w3yzHCIfDK9070V8oa+bem07+xvOVsdRQZ5Wmm767JaBQGQ9I+5ev0gKBoiTTZj
rDtk1a7/nLW7zgB9zyLvtNf3F1bW9SkM73vZTqFfMraui+xv2POx6Qg4bGEz5o5C
A9sWlS/TJeIrHrkJsHWw1XThXo2DZOH/3fmXYrd3UUypIbebFMH0KGqPNyFNbWuf
2V7Kio1R6Lpa+omhPYAkFFTltctOA36KdxgU/eH+20Qsk0VYa1aXFrhUtY90J2OY
Ynej38LgtNj5+b1qm3pqzOfMwhz5b60QLA0Pm/0HiUbfzjKmyqLEeK0n8qTZWoiz
JVGcpuCo0g3ABipY6GzZ8nXPUquCxSwJDV3u6NCmGRSapMOCo6LRcvuEBn69ygpU
QxSfOwcqTSMBzqXvbqjdZWCzZbCJUeoQnBvcWxrNOAXkvWQ/p3fJEkfv3S0zFvTy
C3BUKQn7Jhnr2LoNKPF+qxAsSnntH7GmPc77NUc0P7mPRvIUr8MpH6mcZU/N9rkn
kBe6fC10qOnahJs1/nUn5KXrqCwnMjh7eCPBU8AUb1BYz6rGmFRCFsdBg6oPXcSV
+NSXrjlW7aFgfk3V4Hf11yYUDypwal0/zfreJzK7f1Pa47ETi5vmNjHBGNsHQPyB
IDvI3jf8kEc6hP3liFEgGFCPzgleO0zk56MJn7jBulhm8OU39SnefVEIr1AtEWMn
FPzNnSL7sYV7Uq5IKqVLgPAahjYbUjK+gVS0eD6g2xvL/gVM6RioNC9HGhp8oYO4
BJnlDNwJMPwUBrziwHnsaLtDFHbQ2COHcJeM00/5BWoq/Z6lo6tI3G5Kh9q8Lyb6
hDyfLa507xr/pJu1vJlkmTFGA/YxUY5mBs3Ulk5q77jiaVn1FD+x1/Bc+fAU9HVb
tH7BUX1kIhDh2uOhYZev6zvYlh5ITiBIAvvbdM5rQtVCXLu9eSZwib20Lv4Mx5ys
LlJ/m3mOAaLyY0fjpmkmT61NsbJN8XPF1l1hwaIdJinRCHn0k3E5L8nlUYx1Kwvp
igutKqNNgfAaU/SrofDZ/298H7tiFeau5lF28gEYD4pTNJsTePVhVRW4gltU8L01
alLBNR7IDZrQBbU+rQrmmFCrQ0B4g71eICEZvETry/BvFDQBjKVH6E3XsuGhthSI
C1EFpSQ6IHVcAvvCXQN4Q3WW/yAO5JdzXlnuUHxTr6d4InKT7HBDW/pTZoXILJwD
oCMeons5CpY8kCwSoeMdscXJH4B/HRFrht/BOJ0E/k180blBQAiv1tVWAONWCCxW
7N61HIQBNJlqN4Aa1bY4sZAfQP3/lA/qcfH3mdgItZyqUavK4JWkdZJWbDa21ONg
Z9wOnnHi4w8YbnKY+rYolkFjIYrDUnuYR2aZuPjNYLRv5J5wLkYP5wsi1mdJuX7h
cqU2WZRhSGPbz0PvZkWeVQQNXU6CoB+hb7T/X2/1ez5uYN66v6MHL9XHYSPnVH7s
WSsvzgUTRbAspKa8bHQsjnv5cCXcLS7qR76WTl6o5AkcVFPjfmWom0sxQ1ygJeZx
wOmJghvpnZejFZaCcT9+9unCsoUE/RT7tZ2CeWMwlmlKAVbo7dg9VL6glLbqdPE7
L0rasvS7thiup+RGJL0g4wmVx/CBGQBjdzlsIbPrsqCklz7JF2Vas/WZ3tTkIqFV
7Jvne7PeGzqKahBPz75g3MTMCHc0i1tCzFw81OzWFoRHWVz/iz3i2hkbDGoPIyEA
qQapST7UyXGrHPvA1K3LwxsvtMupTbx62nN4dYKLtmp9+oZUlAVFrxE5Vt/9w5ct
Qsfm4Qmh/hFkxK+qmSJalRtlczc3G21k4rrhIM2XTuMwcX8JuyvTfKKwafmxG7lC
w79A5HFSonyPAnZQ1p5FlQaUvoWosWSSR+7z2V1bODBNmHK3rxFoDNX4xQUpArOW
vphQWXFyCVDer+QlVz1C/A8PIJk3s33pqYM1eEYUHTyLxOJ7aCwf0dwTocKu6S3Q
HDs57kNDG2g9LkuBqwSX41JKDSDUB9F5FWRXCNVCgFw9WcdCTT7dy39aJO3bmnCo
EXxWeKKBiuMpGK4gyVNyjIzijkf0T7Qlp53HLBWDJWw8neHHXlfXvvH3tQ24+rVD
iHyNpzzvRMNiU8eUxQl9nfQz8wiDyRh978UFXM05yLnwg3pKskafPptYNhdEvKu2
tZUiIYg0j2xfVpnP+JAxGAKNGwmb528luB5G0edcJ9eBY8YnNlSK1uLqW4ZhJxbD
xPlh4nvTK9jCwiNW7ropzwDF5UHZD9Ek4EdHLHTS6UM+KKE94Z2RIhKnd9Q2UNzC
rRv5CfL7MR64r8XX8Zvi6+YpxGZd2jq3kaEzFbflbOu7Dydzdf86tHIzGC/NrSZH
EJjL61/xHBbI3wYB4MVUTrLDKyjICUvlamFq8CngDTiC6kVGYSwETOeNbuWwmYH+
Rf7ABvhz8DYfQ30cgOy4NTd0ls+2sjhSfYKmzSsbMyTl+uksdLO37APXj7NHacE8
C9pUbz1TKpOmjccEFR/59dyMxiJkBQTlxXqGmDSxkNSy4CSVu+DlbTjqGNymQo/M
GcJMF0cP+4HDuWqZux1h4MsiA5KLJIvUn/1FD4fCDh0kShdNwhd0OA/S2Dm8fh+l
bNJnu/JNepR54j/JVBU7cZYnHUZDKalxMIGZGGnsSiMsE5HSEVn2oD10Jsm14+jf
ve+88ezZkAcXg28ZC5R4Vwe2ogj8lJbyEbKblnjCjqYBTikj5rdECHL3O4PKGgOq
kgTfZ6B00CvO+N0w+S9DNQW+hhLgowsZGaciIqn2Cp8he1cZvZp7eAgEtvcJFkMc
IaJp/u5JLg/t6ssWK1c4K77znLBW1kYfCh9ZCRHDQFZlDEa7dxg5Z54Hgzslos3/
sxkw4FOxzn/Xn49wu/vDE6hut4U9JAhfYu2/WHCvtAuj6+EDk2v/DtHjrwJilRBT
MQBQuOeXwrJJAfC2/yZ8l4aF1V5hYIFYiwBVZNHwctUy9y0zVEd711jlFGVoC50P
T4B8w64Em11Gkc+AYDiYCl4yOO4LvHnYsmjeryPWou2jWJJ3wx8ezUWCMpWsJhhV
C6UhyDmX4LAuvL0KZcsmxoryA7NSTkXLm1UOQ9tnXqCD+RsGgvNyOYh1Km/sUri4
cBPbYm4gmm+X/zDBmRYTKiVc3v9Ue3RnnvBIIGUwFMlnkVL91RPU7YOG66rh/wD0
h5sCz1JThufrWlhaJHfZ8htd3u2SU9B+lxET2JLvmyjo5F5pr7lIEJKoZlCTwhJO
L8Qq4l1DTywifvikyKgIp+AYZ/Bbn5Zhq/pN/WQofjkGfVKwnkw5DSJTbIejkirD
EMBhOlZeJBZSkMKuKWI0yrsQN0cCgLW30O5lECtMI6HdPrmd0yBSEaL/hyYrpxbg
wlItwhOHAfj5SBqoQjK/R72yTFoQuKsCmYg6KqfH1cxswelQEBplbhWQesAOBAsd
i+upplx8edNsF0hsHscmiS+6EjO0CaOqMvHywn4m9erDuTdR3vYimp+p/dxGWPDv
QAfL0nbpzcEI/+B1vH+OMBav9pUNwvToC7pBBRL1roEl1jyzKHYaW8pThYH9ouUv
1kevW59UuWpCv2s4IrI/zGMNPP4C8rLpEnhBW0bfx30UO3vgdfGo4/kBE5k3EPSu
e40I22Pp+oOCrS1Z+2rlh2EyyzHhyDoA21FeylWL4ePZQGk8yqUFqMJThrvqneDq
DfmcvpveVH2k/xn/djQjvQQU2nsSRLUjBOJbowbeNxTomxz8V/UsHwn4584uOihT
GidbBXhO/TKGTpPi4Frsu4z3jw/l2fA2uR8uqmCcUeyhA9nmRAhj5gsLbA9jPjaU
CnDe6z9X2tOt3dvffaHOJ4blj4WB/DGOn8qIrvg84Y7dx7cc2XsV4CI8R+7Si9dV
r4wO4lh6H+WZoQClLw2fKLpyk17PliPlW2HEXqcwdNPoa/hZST+ePZC3Oc0Iwopw
G00UXpAVF7r4Z8msb+4Eta5rZmJ9Hy3wghtJ7rs773paZZnfK/t19HQzXr1Zfw2B
I3YBfDZntDlp9FOearpPeAYhy1XkcZHSEGgXuyyVksmB280ozwNQ+vb8sIlprTTl
XV/spXilKWWHn/Y/tv7BUfs9tYjd65woZjn3eZj1O79rDijd2sz+G5OAeMlmzUjo
Q6hvmetcqxaa4jdg1gxIG1OTWAo2rDjzTwxJ0SxxR4yGo5G3GJON6w9nc0uea7sS
ldONDCNkfC3LRWsfb9fzPkwZc+yA+cPmCHmRQz7RbbPK8NPjF45I7SMXzeTEADSk
pJZ1A6EpW/GgtUJrfoJ2f84cU99KmBUZpPpooAST9gf4Z2uQ2dH9QXbSS8AJ1VsQ
4xdCBK1sJwh2G6oywZDmdwQxemEFDyBkJy/2a9YSaS1wtJT6MLKFM6alkp9QoRtN
hy8lP+xprRWywrFmrNUJlRJ3sJv9JsZH9FAsOkFoL8EVbKkqmdgpj7fPpaQFpdnt
okGNUtTc+gWpXMZBrYsK9D1chysgXyuZpTPtARk/3iqzrIBjfhz2KCodjQD0jK3k
zGUAO3D5airMUlE11xY5dU0jTn9OCTttKJ/pakNrdNHNABndn+evL9oYgCDUwbFB
ixAzE+e5Ofpl/j1YXNqZSJxDn/ZWWlqjs6cPPcQ78X4ZptWVMB1pKakZIXukyb7a
bfYp3U+UjGBat9OFWOgvH7eqdHmzVM0ulqox5ErAt9CGIVBkAit8yM6ccCvDpERH
4C3iEituEgq181AXyfa+DDHsjfTsVuQnbE6z0dWA7WAy3kq/qjB70THgWOlELSRA
n9rO0e1hMyxeYlEd95jv7s1ziTXxq4xsK16wGQorsfzfmiibH7ok1M++JSTJ3suE
5CHW/N75771as2jf5wJZLaiAzOCIcWcuKvqZzV3ibtRvgqzkm1R2S2ii04f5/6J3
SjUfz/g7/Kbc8vdcoPN+ZbDVbpNxvWkgrfqFCSE8Ckt2D5CnxcwP2c1nGrZyxyF8
BKIfkRLw66LBdpTbI8hSNULAzebNpt6uf65gwBxES9rthjSYdx3O1HIWzu+DQxlS
T4iObjatsxuL1EMNKAjDprtcgkeWfKsoUCnf8SvqZA2SuAjj/rgjq17VkFq2EwkL
Z67vk3al2LHOL2Fnak1JRuH+Gjbusbqi1K47epr1TJjfeCzGyYHMO4wzcowxZ9MK
JWef6uKuskoLD3F5v6uop6TABeXMTATk74NIbeDmWiTXs5flkJAwrWiqZ/y18ykV
335TmyR1km9jjjBbaxzDFZB3FPvxCGSMQSgzzlDZTE1ae0RkyWXJKK9HN/6Sv+v1
d1jomi2aLUON+O728ny0dB/By2UDdOy2LjR2UJoJLeXQ2rAjb3Ur7DAjYJVxBQQo
Oomb2/DGQ0m/Z8QF/npDLb/8Dtc5Fe/8PS4rEhcCcnUxYNBn4TrYGENR1Wd4TmVr
stjUQSokgprQDpzF9mgzrKebveLsIgDd0OWklGJ2FRR4Vs+3vs+blODEo7fSpi5W
qPApTAdcqM4aYxO6csc6+M/g7haIaAPxG/jfsEq7q+7th1ovCoa4ZJEWZ71rO1YC
cCd7U2u2CX+TLuUMX8tWQzISi9nFruHh2EFyOcZuIn0Fqqg1uNym2kkbVAs0/8xv
S02p/cZtJNbNV+WcahnMl/OCVx9UJ3iVyapddgIdPn6qwt6OPRmxj6wycqxs+MP4
MnAGDjLHErsu6320k91KN+z5ap2V+SpZ5GNdp7yWE+8fYkLMjgW7Mi7GpfJ2kllJ
CJSKoJsvhX8yxoN4RNrZzpa0zJ7rIOZ67hsN0OnNiUPsWpNfnHkICdag96uQarer
wdke/O9ojE4thcn1/wUYGvxV1XQg/eMg64wEfNOzkEYcOs8BZYikkmu0FAQOAz7w
qWG6Z2lSVCaF0sZYA4C8tKbqs1H/uFXEc3a7TEReIBjORkDP8hZMY12rRu4rGnj5
KKkUG5rQvKYTLzacDwm9iFVlLrhDdtZ4Ezd1iB16PB1TYt5lxa1ugFGr0TeQcOji
lJljXu8HVD/pg8jsHwV6lOIgBD5RZZXAM8rADwps2ytD5lKJWAbk1I+hriBdL/CP
0Ijc0m00qLsWOMZkPLcTiYoDzDtqSwT/mfTV4v2xkM5H0PDe8ssoUf8se1fQNX9G
fzS0LJ+ZcjGyW98Z7NAcJ8tJJb+OU+SvTIaqhwIgNXkeAk+pNKSbfus+25G7b/I6
znhxxhw4OvW10Uq1fuis3yjnJcZlfhBmeNc3sD8unCqQZyE/h+pjTAZM8B135Hcg
O1EIFqXJWlMeJQkRugAgV6Mf9lMaeEHzJEmyogizf5/8jGV1cga02Bhlm2C219cp
vRC2BUos/3N7AIMrw/+0UQLFrKa8Tq+jH/4nHZXk3CCS8HiJ33+zuxk0Baf8rsBE
OryaSRkx/wrPG8hCPVfS9xUdD3N+HyFRwKUDCeFHBpNIbr/qiuFpCjZq2t/YRrdv
DzIwrRSBSnaMeNyI/1l5CWd1fjTJMO2kYm77bqJufoPDeA/QpQYuWUhKQ3anEVRK
DnhFGI2gtyP0R8IKC+wn7wBUP4jMJVfp2XdBBy7D07hudxFCVcB0wGm8hjj9guvb
srjbcH2iNHkgALW44dl9uAHSdM2Pp5y4wtzE2Gyevh7YovAoQCLhbe17aNsffdWb
O6Lzq4GSCFeecgg9Q64w/gQoZXHOSy5L+PvHV4ekrRXWXmFAs20JJl7JpJ/Ml6hz
nj4LFeQi2lnfPuiTbhO22g0ZTOLEBl0AmRHJTX1LfwbaM7RoUg3q7gg0Ox1B/274
Ls4+i5dgjDo6/EsxAlXQNyK4DoDb77K7/+MtGdmWTzCRoZHD19q2eImYiQ0jPsRi
yyA+JHiMifZmjDi7qN3/1pL6au0szO0k/fZ8q5QJ6mNu3EfiCiStc/V+GCh7TlYj
tt6tr1aQAlFI8cjPQqETanTKjW9X23dwzGOZri8dfiG8JuEg3X8WV4TTVoFzi/5r
6Tcqbwuu0AH9RSbw21sXLkoy7LVRV/OUMQ6WlUlg/k45YCBxqjCCKfUW9Y2gR30K
CKbjkhYaajCPsg4g5r3zUC/c4CllhWchzD7k2YlFd4UQFixkYNRDSYg/WFHcdEkn
VjCOOF0UTMRt2JrPH5hQvBR8/dwi9zl0MnNGdQ3VeWTRJ8F1jn89LyUn2Mlwopax
5hqCYg1BPhyqYqWiVhONBlFGBWowMqSEUaaCDrmrVrCPUFS/buQTwshQ02qtYKu7
ZspVXAetf90f6PcQqpwlowcXnqsc9z4DLCWRl3vhvN+elu9K1DPPX8pW2etm3mwt
B8OIyUU6UN4oPlC/M5XkTU7pFbCQQ8rYK7wWcP5wkh1GDSC9VmuUxNSdMdlNnbm8
i8InT01ZyEKJBOtb4lcdATSIUq2yM5faz0rKcw1Dbsdr7NhK9UPMiAVAm3VHvv28
C7tOXngiwydHgaiuUKCioZbXilkfgoBM/Z2DYYDx1iB6pDvDWIuSuSuMVo0wUquF
TY+IlZQmyRwwYLgkeK18HhMQz0+/EfYJQpXhMqGxwNKTB03zNUHcEBsC/bPXFXHS
qVWJKAXZa5iNjTsN6/aE4bz3UTSqoI+0zExc26FTeWn6utjgWEYjCIuXN3CRcy5D
gpC8ADhTqb4K2ONn7UGJJEkYh/0hoOONdsyccrtVHI5wIDzdN66OmixmEa/UJW0u
ibF3XANY8vgn9kWO+gYxvvwf9K4O2z/h6dLb8q9Jm/Ylu0ukrr2wYrXReqW3R/ic
DCsFOixhdroji5v8s1+JsWdKYEppJROGQz/I39hwTgHGLeks5fq6L0PSgwrdAYUp
SPbBmik018PE5HmmKQzYUdexFTidedvAjGoMEmTMIkct1pFqU0v0E3geBt5aXk2I
rBHnsn4FVUGYJVLPyQtrecOQfY/VuwCd6y9ORpoV5AcDmmYRFkQQUY0z2KP4nAh3
HDeFgk0VMYGiMDMxo+lkb2ivo9tbpyi9ZnP0POQvguNXXIjdnG+foLfIGstuLvRj
hlcjkbO3DVLkx+KH/qu/53XUn3HuEgs1+wEf8NWjHOb9mNcI8FfIAHFpGXkDcQ+a
NvssnDmVpXJw6+mMq48skVWXLQwxYF6xxxRzMlb+VnDzgC/VvGhBxC1ftUhmkr2U
irEPY7BC9tci4o9GqUH/F08dWaU+W/JvQiXM289sML2TdjqFspEr6Zjd1+2iZSyM
PuOvKBHZ4qqyBmCK4w21cdDgh7yoB8wGYCzOujIHnqvtEJ/FW/W4HW7MvCoc3Lar
2FjwUVbyXEPR6VOakbDdtrm7hd/8xWCYNvBaTFrKAVXahCQ8QhlYsMG9fN5wWDjt
+k2ucN1zO4TzMZPnWX1+0ncsFLiLr8CMeeGTkeMeqvvVkgY9+fMDf376weF8lb46
G9Nb2hTzELxfCO6EVtKih20dY/GYbiZsN6d//c8oKVQ95wggPd9gSaz81Wth1Fia
V3eiz7ulW+EEkwI9bVvrH0GSqHvjRIEJsZQxJw/Op0UEyc01Cov1bHOAPXb9eFMb
CY/jiV+5q12rNAFqY+Z9jzvwKCCnzk+Pf+uMPrvcK7RymDTgGPNnFesR1/mmipXt
ZlUAlqHvZdDEouZi1gRraD+NuKCSIaE5yLQJG2lCwmdaqaNTKCxuYYPzwKqvDA55
Afyynw0MNNK8Bfj2TLJtCOegsr+7qYI/9NR6StAX+lmXEmlWuxCKAwWOO3IvUsbV
sNOtW/Z91ycGeyhFPOMy9MIz6Yscpfk4ZfBre4o9VhRaYxxn10RrZ3S+C3vdBaDS
LvQwIZKHeWqtxlTzG0388dqwNkZimLB58Hd+toO+Qkg2MmjFqmYaJlEVdk/w9RIx
bI2ofV64EUvcWYrNqyVhLLwd2WU4EzdJXdQgAdCOiRbgxe1IlSoVdOHwjLdsTcMw
ioIX7oEXu8b2iFUe7eZQdTgVlQzdK3Irqq+tKsAPgMQqAyLJAemJ1hatD+6ZtFXR
AX0AfoQdN4qjTYICbfqtj5LkcIwmi1jEbXAuEqXCh+i+fafXjhZYjAaHiSckZDCg
2JO/ytNIEOK+HhWE6d1JA/qTHYhgi+m5qOwFx3WmtvOYTkQkiivQZ/FSbasw8UnN
zsbVteA1o0rFkgra2YalyMghw/3DXav4bJggZdu4q5ma0S5RmiMKNNhYpYtIyqBV
wHC41+OWXIiyoytb4OZA80PMcqgy+Dsw50pCN3EWZ2T9XBHCspVhWGXQ0bRUcARW
Wl/3y1yG1APQngciPU3xe0yeXWTPK52OPMf/x0GQ8U02GGPyYdxBiq0hhPaienKq
+wXrMvcsUuI+v/OPQ8L9nnuU4mBsjX6D6eB4FUVvcTZhlyxks5wEJT4lhkJEg0Yt
2uHQfqF1yf8kLEV6GK27H6zJftJtaFJJD0TyQ0IXW26bNDn5VS8pey3W8McHMtF0
qLtjfyi8mLQWDnSHN4NU/A6s4855byASVwdY9W2hYHzv3hYXJ72qyfiI0ByJ8sNK
VAoNINbOO6Y+ek+h0dA5dWhnYqcAK2Urh9kIANmIZJRDv1jEQ910XGmHhUY/jvmW
sJgFlHv+QIbBK9QSb2hyGZsWyc+uxI3ci8XjzEhJm93LgrXvGIii8hhkElE4bQwL
3Dm7SfwYx4p7WxZs5eReyYa+A9/yUTZAYEqhoR1mZRNHL/9DaOwHlsl7wr0GHHk1
CySbSe4YcFF1VZ5pAdUAe+r4kxljHu6iZhVziAG2IyK2OWnIlNO48a13vVI6gYfP
0sj9LEC0+EIp6LHN5QlZPWooFyWHeiYm1i39OuNeV8xhjnAGKNvZGLQZkvGe/uA0
4wONB9GazBYkNPdZQmYqNgBuIyusl1Sbqzxzj4YuL2GKN6TWqVCY1lytmk3Ra2gW
FIR8GlJBki6RGa+AB/I4gEC0Tle8BRsFkf5FAQbskWPRkJyC6gQ1x//scj1tFZQt
hpaI9bVIOiOq/j2HHR01a4YBLHNJg5xyS+MOLSeAyR8LSoSrKdb/yJbnspE3NUGj
dC3S+V7//INzE83y2eEvI081mbj+0XgdpMcBaRBPpNeus5V2hfIQXqbmXF4gThdw
X2ZxgQQFn0GyUGOfj13tf4FB4St380d/q4QLCHx46RLh+J1uRU14uKf3UDuVBHhq
jvyW+/6+TGlsZsjtTApzxgtzpymaycDMo00ETdkG7R67Nrewmb5ymmTehzx+fYoD
HpYwKkdVlAd3HAW2e48R8xm8x2AKys3hUxreyabTnpLP5uXHFKrUkBnCDgnIeFdI
ENV8j2EcCV/GRRPKSInZcBLxax6c/7XU1LnRyvWKhaHDZNSeM+i+iv79Q5yjhUEz
VnqTzl9uJKF09JbSHM40ll4Bt59RTkoDLIGCkwTEO6vARWrTHrgsxnsSf1sYhnGS
V4yFrkFv6FsPLyoX53UOuDoJXtikpdN9Oj7ZAIvr2kyeCjWyGjkEu/FZ1ZwZLT0q
plPFerojYW/4b9Gks3dbeUt1QpPUQkbsFOF5VMT6pfQcVzNksGkuwjPQ6ngegwsN
oZeVnkGM4zpAeO4ENx1HgJOdiw3rhBPQdkb9JtJe9LeBb18TZf6mwySQnbhkWTwd
DjB0p/KcrrO877zd+cidooRHqPdOyoI4FP6jjx2nk1Lih4LFfFRtfGq5pUlnJcGR
sntsPG2+kPxWIXFgtenH+vSLddqW93uRgCW5k4anoeFw5q6l+Qa8JlgoJ118Djjj
eK9mQHGxz9kgO8QYnwEzxtTJUOub3/dQHGMijRO1ybGKfNRipCMBGfcHcvuIspYc
Br1Cxbq8jdTD9xWVOmmCvKQzvu54dg2MWRxtVy/m7F8et5MW4vBsZWPfssEi3/IK
yWsgCo2Es8JXHDvpmldPJCAGD2Zq3JjtvzmD7U+NNIXni2MA4a3WYxyqUZLc2f7M
vmcyruXJ/isj/z5zeAM9/XY6RjWOn6AXJo+PZach4ujGOfZKgk1HHFKBq9MYIMNl
QB2PD0je9gRESRHftxabd/e2ArRUYsbEjwRGnYROsugNPyVCt/7B+4HEC4ecdcgM
tLKlkMAOemHPYWqZuymyWCDWYkHLGnBtGTosPkxqXrjSyIq06XE1gWxl6oF0dzgN
X4yIXChhGGCXsdk1h9l1iEaa3GzRbG43JJ4dwQQmRdbcfYslU+DMAEJuacx0ZoR5
K503EaCCPpCjvKqQNbzB1BKwzzf8oqyo4/GjpDtIxZnPvT4DforPK9lOn5qfgAWX
DH5Tx4jxUhzB9w3iQPmNLnSYpVtR3HzSfN9KivET6qurBraVTQ3r0VeGwi0kpBuM
LBA7LrECC/0M4ASJjHBozJFfh9rpgFOnRYD9/wT8Bc0LUWvTbYnwMibtavb1krPL
5DEqUiLUQKn7ERB5OFlRixMKMmwRTK1mdupFFx/5OClyGKOcmBWSQMMDoFxuoWv9
QbTbwrS24micCtuwYvscNUnQD9UWi4e31IJ5Da+tg8t3W1hyYLLN5DdnojWnuvNs
qNnIm7eTrrzToCPAXtSdO/BA1PkG4I2rRhO4bL+k+UBLBg6eCPe1a9eGAcyAaX4W
NtJilwoZ3lEvjLZQRffkGEH549l1WpUGPTawLwXPddDt5XzSPB0CbyHX4umh/Msi
tr86jLal+wqTN4XakWNjHw2WQAdSw3t7JAbMzLWXN022x2D6K5/z70YqmqLqkrBm
4Sf17tt1pauv+qcg4vWMZTfJuOSn60xNW/fxMSYtwL0HvjGpb0N3g7yOK7VqiUPj
CQerU0h/VeN6TRuSKO+OthATY1ZidrIgspml6fGkIlN6CWSTtvhszfu468icfzmP
IukDEHv+r9Zw8rc6YYBixAQHARfweGBuhNitrdII0F0ybTmtSGCY2/hQmOM9WExZ
BNcD+WnsxZUaaP+11AuIjkoUPl51Dpsrg6dCuO5nG0Y+xWIhgDxm3jQjXqnx+Lix
qBsgaaDoGoL8BOZn1CRVHm2+/ZvTiMgmnc8xH4tp3PX0QA+3HfIY788t3riUAxaL
QuuyouOvh9NJXh/3TIXBuOoBU3qWHT6xsWrZc1YwxJcb2THCKeIbBQqInE+JYjjV
GUkZlsVX5bi70krD8J1w5J5/b/8QVbf74g1pXsqvCnSH77gq30zBKZRa73fMqnG0
2kWf7KIzK79eWYCNxNRxbadIChAegQ3WOWZk36O6M8L404cc+JtJ0Dp76ZtvN/OP
x0XmsdnR//jrRFFt44FzybhTlNaCDVXv3Kkr6F2evZn0qUyTmHcRQbwbG5+voS+3
Opm7mYMYXBeYr6E8dOe/1c3im6D9KfN+BeUP/+NUT8mAsnNdpNlYI897zv6E4AhI
wvqMSxmv846ecVRPxaPJIARe5xNb1Q+OhS/m2NlOIHQHdjYgajqvoz1QC/60kqWN
snh9bB4uhymh1s4rQr84mAHzr0U2MVHB+e14KuLu2iMAE32lgV8/FtvRrHMk9/pl
p1pDl1/zssJRuVskk7CHUwD8/1b09MfeX4iVbgYJ5mOPkHjopuyrzZ7hRJGzhG3S
XmjFJg/8+Bgq+PavjR+Q4bI1Xslq72c4JGklco4QPNfEz4GmNEivdWj2J7tXyPDx
pdHaSgqQDy64zyrSO4ckLHV6yf4BKeewMLfZuAVanQtrqyKdXCDycnedC73aSaRE
g++YxbX7LoLl11l2qJSO39+leAjGa+AdWwTx5r1sfB2miXzGkES+7apL91JJwQgJ
Ncr8cpnPCdzCSN+MItM/gjf7QEWqsetwov1gFwpXZi882NjHlPF+wUBSZKPOD1SC
ihsVmXaX3TB/MUVylgi/GUO2z/7CbAhUtYSVKjbvEjLf3VAep4yZ/KwW4RQ//1Wt
nx6t2beucv0I92ETZqs77RL14/GD7M1yud0/9ERY8oy/g8s9OvFiyUTrz5ThUi8/
Wrx9yt/uvpkKLtSC8n2dDzNbTDKhLE1gyqXp6BikLN5Dc2byWtQ9lRANztRCIcJv
aTTT1phDD2RLRM+5aXikkK3Tw1k6IAbxRuwNc+GAIGCSm+CAUveMNhQ/7uaXA12/
xDg5rHfY/kWFdosDWKNLvXNBCd3FhktZ2wTa5Vu2FXX7jXVFcOipnZt16DVAX9E6
itDseUTCMbSEHg8fAT43AesDEkhkql3ZCZz2RNt3gS8ejohBPszdY/+4D5Rxt+Tx
gJgH+FFWnBQGZ/kocHb/DUMSU1UZOBB/MH2CgfEMwGq+wQhSyrR6HYFad7LoZaJ3
V1QNZeBQNiwKLnvZGXuVkzs7wyu3oMJa6qD7s2duAzN7RpqPcmSwcM5Rv4XYBq8r
Eky/1Fu1G5TA9LoY6II/DZ+MgmgLPZURvoyTktdG9QdfLN8G1zbDMJHsvw5Es4VG
uDau/YEf24WJDYODQLB82paAtvCU6imNiW6edSns764j4cvKcwJfW0VDZdWn63sG
DitNolN2jfSonsg23oS1IOU47fq3gCjuCFTdz+UkGmI3lCJ2pSNJDgiOuNuWjMSd
iLj+PG2uWWs4w4FEYDs+B+G8EfkmCZ+bcrphyt9IiU37yNCfv4ZWikmWBT2e/frx
aePCt4z1n6Q6NKPhnZSGGBOvU9JDWyLRcTET+TYdDBgmboN1ZojzTr4JV5GYK2FC
RLN9yFZtmUi+wBGXCDKhr1zSqr9ctQicvDfqGYU1PC/bTnOid5oIr6gfOCrlldpn
fUdFQHz2n2QauD3kFKiV2nYUupW0iTF/Kp6kiXfXv+8GwO2BSSBsL4Jc6tbnGpuX
mf9hq+K5Wo2eI+fEGQ+19cQqd0bsupFf0SY3XPILnvaFMpVu++ZfkdPfQrn+W/3+
wB9LWJudp+SqyXHOJ3mjOtV1Re5VXjevnjkuHjTg590kEgbVBNjoNfKVCjFfbBn+
PJxmOk2Ccotc88TJ38JieQk7zhhV+Wk4lOfMMBlHO33/dAMehRjkTgcRG2hbY395
+J+sIgEJFWT9nb7i151xNLsLuGfzAqyQj059Eh6lGJ4+bVOrwe3TniybWz23Ro9Y
QPwj5OP7ZPa171I75SdK4eqB1+8kx/dISiqVpL3C3i2hquKO69w/fkiu1hnYxIH2
1VOfPy7c9mClO/gJ3PPkr4a8JWzm+7gSu/e4jPst0CliC9WxiFfMeseEKMFCI0uZ
8oi5Zqh8R0QZp4cz2BPEsQTteR4bOTt56yR05VUH6+2t/nLaxVdrhY8qKPXhfx9m
U5wWX1d1FL7Fg3BeeGnec/QbyO8vNBydKb/QCc7oetxdXGkHI0NMASZVIXBQqxMS
Vtnhhqzy/Q7ZoJ+lI7oGYC/Jb7Wr7ABkDmqpwb3wI7hy7PbC7dZyNMZSUkDkH7/e
04vi7c9q1cojzC0LE1eJbboaMou3L/8lwYakvYvGRsz8PVZBDer50Lv9Hqu7cVZj
sErBf4YQr/pqYwjO4wVblzrtyEn5meZg09PfMWik6abjesnMmktzre1pV4kTgr4h
FUKJBmgGFN+GXsl0zTGMxmm25tPuqGCCsaEjWdGMJ8ykZGLJjgxfQ1aceoSkTBQt
Lz0Vh+SbcsyXtL4A8e161g68NZOIkdJTNiy42wXJ5sjUAi5vEeaaHJIwoBWGltwP
3LAty3idio8CkCYAh8uVw5qzcYr+x2uuzTNkn0L8rxwoRx5QUqT/A6N4dGvc/kVf
b9dpGTxAXePT+JLXbgJLPj5Q7wxeEwRWOnG9JsTn5F+xCcTy617+DEpCwfIINk7q
BK+28Y/v/XQhjy2gFB2zN0WTaTnyYAVN2myQNWNmMknKhqPkAfGBQau2JOtiEtc6
BbVD8Wc2qsC0qNmuTChm1i5KEX0cl22rCbg1FGUcUjtelU/AfoAc54kamZ50k3Ou
9QJ6jYiWWFdCpnxOWfKPuooD4uACg9G5WqKw9a0EwUER5spwmE004DdHuHaKdU7u
hUtIEotPfzNEM+nV5s8y6PCbL1r1M/2wpOcdyFqktdF+AMNmRrnk/r7+9KxOGZWE
yizWHQMtEBtpnvYwDW+fw54UlioRi9a8uwyJuDTYibEeD75MDgONzlQbSiU/FhWs
582KdFjXfG9RuuLLIsEkSbAGtI9cjlg3T3mr7KLIcOfS/eGPkdFjHk83VnOdbH7g
jdM7wq3uZDj9yEv2eCV8YsBNSb/j8oXHTyEeBvC1DPQ6k1et2X1EgteUrpcLymlE
R7NXYC00h6UhGMr/caCgr7pXtc4eOyjpepk2wmr20X7ddZHV9fBJ+ywk8USyuJIQ
IZKWgQebr5KAtY6gRuvwwZ2iU+7vNcdrFC14ge8LO3cORh/DQ6Pr+ou2Hi4Kx6Wt
DY2Ok+cUe/GjEn2/5A3UtNZcYVWFguy5TaLmc2HFKXO3XcFz5h0fpUkZzq+vSbTp
WPwdZWyss9WZnUTGZ/MYP8Iay/nFlWhj/VkpwnLhR4YbFeNZBPaIueDWW3jKcelM
emtUWeHgGavktSkSLTSyca0IIoeTPwjLE797wV3depJdtUEqMQ7EdyZNnXjtw5SJ
BBJwtnL0VjTCyxavFtEKVGGak2w2TokpEsUVbkagJ3LhQuqoOzSfp6qgRE7A6BMG
6K4P9nnQVWjr6Juxx223kcYXJMTIh/7PKdtEPL76130tsrcxOnvks69F8C1aCu8Y
c3YODkFfFSiBjK55SssT4xqD7g1+7I62uT0EfYvuS71M7G9evV5wmkOBVa0Ola1T
sCbX49oISVLP+Q2qfC8PXq0zF+BXkrGSnWnQa8glv3CMZRQc885/TF7f/2QRPW2t
TPNwUwd1rTYBscUBkFK3z0MOcQ1UwTGuZMlOH+jybPYbycX35N4wcdKlUifhs5/J
nnKjUaRU0cNnXFsnFrTWXC4/bx2We7SJ3iF+pBMOFsng7CRhuepv1IPsBZf7WYS4
r7Z49pw9lUpkFha65TAcr5MXXVskI3rbogpNBvgqFfOzzMQibCtpYH/9k07PFUq1
75xXEkCaG9ReivF3LujvfAkYJE1Q7zhjaTZ4wXwjFPZw3rlvSHT2of79xc+JEKvN
gCTnE9in1mZy9AcDe7ZRIgMoCqnP5sE0IyI/86Zy2/sbP3z29HMojrV4LHIKlUvP
ehzWmclCOO0bwzoMFSSJYs04JOSrmkFJ3Jif11Ys46MJ4PTb+HCQTHLvSsRklQ48
HHWRXVWfDBIc2jF9ZFBOrj9VGjCPbGxEEYlGEd5sSbwIoOUD6uA+8fnJd+XR75cB
G3g8j5AgzH3NEeSSSKRdSwPUZ8jRxJhM2pIV+pYoetA32hKOsYlJMnrOkWhj0gZl
IR/QeUQuEUOrEYbfXJECE0LJ5Ka0Fd994TVWjlJZpKUsUxLoBjOhRzBtu7bRZzfN
Oareo+1cDF9dXk06/mOa3W0ikc/1UWq4GtQcA9vPRskKsY8xfpPbqugPjVvMmcl3
p5YmyHVO7DCOSzIFBN4u6tvfYoWYA/MqFD3eVtlPUhCMa6M2qnFnmBpWGficbtzL
7+ZsEdm/EKhu2xT98b/CTTO/2/7uFwR/zVElEHiaNR3vKgaBXvME08h1/q8Z6g20
QKUSH0T27Tq0tRNzGwRraRtJf8MJuo58Fif7NX+mzIa+7HaapW6fSsh55gS8NFAE
/t8Q6arZ4dY2V5YGrgSAae1V5Lz70XNsW0OOm0ZufC28umKLcDeWxJ7YaH7nly+h
LJNO/bSllEejswPoJi1F5KPD1sJrKYEpBpP0s46sHr0wwv78unQvRsMkOg4izcN9
MKm1f9YeNCg/q/+DUJErhXp/BiYmblhyNN7fkccYIsl3mvZUWsPcV7BkBg2zUDjK
ImE7yhkeD92Jo0qCdGFZwgLOVntjPePoAxDQcsviu9yO5BiCflYslbepwpAfktAb
XlNe0cGbYGkqHkYPrutg44pm9ElVvozPldzeXbFG483O2CVJ8q2mnWW12HCy18yQ
5Ac4pMiVjgxIaY1ol5F2nVZ1NibBP4yqMp2Cu6MFFEwv/Br/xuPn/+UtKFGhOUTF
iuYi/xw+bvFRriasvY/R7XAer6rFVfL8jU0csEbCoPUeMp4NjrQpaS9vjxmFXQd7
gvOdFvYCgkpvvCGOZVb1qJY/j/ASI497V1PwQqwIBD7/z0DiHD2fwSBhCOLsOl8P
7qJzsC1VeFi5f9OcWWavu/ei257mPcSIBzQIsNpxrm6H0DERg+JjWZ+Trl86KShP
N6ZMJVwF5jP5VeXPchZFTBC1xNzFpSQ9x8r+WVv11HDG/cxlFutCFCKrLCOvHsue
WGskUKuY+csNL5QWAKugj6QxCyXmNd3jhgfE/ervfWrx2L3l+eJRCjSzMfHDdVxH
bPpAZkbIRkPDj48Jw0LB+ewPkG+hY+JaGKxSysrHI/Vgp5D43qksAim2TkdTRl1Y
Zo3NcdwjRC/doyYgq3fNg6TqWPoQ3jFteBveW34D/wiz1oIRb/3EDoYWpZjz0bWH
RGzAhvqiBiG06yrNtFUoLgegxXYyHy8GAwLs+HE4O7lSdo3+rNC9sYUEUQz8CMjN
/SHJvyrKumu7CFlPa7nf8hIIp/puoC0JazBPVU+O9XumbMpjRAy3b5GFEL/AqfQZ
WihjzfWTmjreOLSpUlzWd8JtfkkND11aX0y0RHTy5CQyzDnYhP92S0qkRubwZVWw
VndCauXixG/Xy7IFP/tsug1EHT0fP5B5YtAeVpXaiiWc4VsLBp+0xdGlgqduU/px
sn0HrHI15/nzIutpY1oLxv180/f9ox+9n0X2yj+KxdctcwGrzjvhgovuDxHHRWSr
wkzlCE225Xl/npYSPS7+7aM76hrOeAvM075H0DKUtlO3F4FG/MAeVF376v7G6Uf+
Qyh9/sIr5B9EtRFts5LCb0Amwf8o/c8AXWASxyFFT2kMI3nVAGDpm35B45JUfzTy
fKSscsQy0yPWOUZzqBgtnpftki2TygLufpICO0bQsWHX2c5FkEmp6VI/vw2zsglQ
HdtZkMnTZsOtQCrYC5JZprSJ1NmY6puCgAH5CGs6Qwazc1tFI8Ut+VdJZyBfKeim
mRe5jGWIp7xGDigqT2Kp+1H6EiGiOVruDvGmbQSAgRXGwf4nrSC8eT+gF8x2qlWi
JEpfTGFXuNczc/WzcVpfvaH7kVZ7WsbKBb5b1Dwih1hibiB+FRFyjuIlFxDxLNrv
A/TBipuyHdqp2TYrWmJxJzFwxhouaABWRyillPE6FlcOyDLLmDe+Z//niHb6tPQX
GjiB5lV76vWWa6jg+bf3ORc/NSDyHrc4wyNBVCGEdvDGRf4CyvK+BZuQ67EOxcqt
c1Isoj7PWLmkg55dref0BkOeiCfljT4zKjDgI/McJHqz+4emo+s3g2SZmNJQCofZ
UqG2h87v80k0PntxYqDGp8XvHS3OeFlaXuF59I3aTUe+tdwL4jec6a7c68dPVV4k
pkp9tPLmVtML/uUsSmHWioKFVcEPonKiGPrE2giMhWoijcAaBRsPJuNepPgpZS64
eWgQGSjTtlQI7XWO5X/zpGrPdnZV6MoHRZyPCCk14INhSDx11N0ZC9Qn76cWlIKu
HipnMJeisRmHKymifNAviiiQ0FK+TMGWJrFa71JRd6+EQY/ur/fnBPxOeNIn637a
YFXRVOzEA2QUD5oOVpjniZLNRSFf+ojfwZX5PFIA1EgMxePvsqz12oP84hB9GBCb
AQjyayXnpuVLNEynm87f5Eynd+s8qxXbreY00/SDBdcpNRGG6QYarM/gGlVr4QoB
Bh7tsMqj8k82b3mIwTjgNxyVGId3cxYpSdxZwSbnk5BMnDDy7yXhGvX1YEovAlif
WgyepQqAgo6AXRq/0OCiD1BGwCTXfxS8hnvc1e7KJGV8JtAX4MpAfjv2ebpG3DK9
TJyk6Zcc0up8dUKBZEFXRZDzK29cdNyKnAiyxwN8NgdGeI76y4EqG66uPAWDNkAA
LNHhVYXGJB0Gv0sqp150EBn++D2UXa5npiutHaGXbek+YJCJuOZW8zi+gojEI6i9
J9XXLntqT5zfHP/gW1VLhgU0saDNCI5SqZSoktSzF0rO31j0SMJt79SdsLpoNy0c
IbsFpnilvdF1YCrinMx8i8DsNi4Zu2B16Hz8I0V7inEFanO5iIHxpQo4vfu7xN2U
r0oJZ9KAtk8lgUb7c749NWAtK/JhiPE2uLjmjjbyWRwr6VzGJE4oijxmpOp2GW3t
C/n012YYz68rWG6VDpI41HhikI2aOuTLwxYdurYUu83x2JRBFc8aKXvnVb93K8+D
qkcjs8iDNYUTHC5EaQNpLtcJXdFqZbiHT8+u0Fz6lyHfyY12oXyejZx6d6N7KAaz
qoc9+4CeOLwsf8MmFBocR7pTHufhF3R5OhVK7B5mYOIc3APxweQMeiGqbTvN4h9c
lOq2QKU6kAMIqFqUTH8a6oGmztB/06hSVHz5/8bMsn5EOb87NDKE2HhLN9B6WurH
89XMMF+gcIHi3Enl/BaD0FAAYW0DO/CURUWx7e42wXttFQdbbMtt+X6Tq/jPSk/m
ROX/b4eOuQnWJLgHkr69iFI/JyhMkSIxbpEG2bM+QIyIjjbYuXIPlC6cDTdCskhO
PT6R2yMPbsJ0kiQ/gO8GMr+qW/hGOS3LH3yyAuxE+eTgvM/JgD0x9gC9wZ/dFwEk
AF7g+POKL4gd/Ik2nT/4FFqe14I6hZg8XoYTMgh/yr/DJnGyC7oFJ1G5yBW3lQue
RPLtFJRgWVcFdxNoE6mW1EKa9GipIf0jz4vZRjqFJjIPYKdfbrFUARXAx/DWAcqn
30yFX0jp4ZGSe8v7kUKpc9RgRyn+07RwSgOQt0ant2gdo59HNbP7TK71PF1slX7o
95W9DBQLy/EZOQOONpigmf43i9dUroK4JLTlzCjjVYYr0rYbi9oqBk8jegsGkIc4
A2vOCImt8LDWgpI/HDw8Qdm1fhqyV83SlMwnt9nkHQMZrqF5bhRvqFVug2rvaQOw
3PJ+R+uxEy2boepBYbvvaMHO2BMzEKfi4B3HcZdBFRsEAsQ4B6bM8kVjflkT+WNr
6738nAmvlWJWDVqVoB7LsR4Xe9hM6qQceZvWG/OTbMtUR9EhJ9H9MmBFbl768/SA
Yx+ExNn5a6vNJCP64o0Zx+1V0J+T9Jgd+VkqyCKD44ZGz9b2R1C+olYAg0HQaUZT
6ZaZ/WuiMIt/ckxkPwZa6urEaSV1VHDiVTXglTcyPo1xw16l85g305grAtdPLE3g
/bw1hpGxrMDdYJgHGjlVX2zTaJAgudEYewQ8IOseBtLm1UYr/+yvzIK3A3wBY0+X
bGsid5uxh0Er5YSO+BDmgwYIMHI0Y5w+78oKQzBGNI8UbhyCqLGNAFRMWs7EUqJr
H4YpRIAx7zngvnq8wZALxfa19OTicBmo0ZGd6GF+JyQ8Z5cCM6HEg6gt755u3BTh
rAtB4CuVxFP3hGq3hsbpDmgDD8KLTYQwgNTc5ZK7iyW8Sytr9xsKggAlVHlGVyk7
G0UwKAbAjn3Wx65P+DcB1zBviN04oYiRu9q6lXgjOaF5O3tbRGZiR/5Kip063HrA
s5JGi/WjsM5IIOQOuWFejlJwIgTvZRsEUrgSVLYNrPVP2FfVS9aAmV/sGVbQHIEF
rqLbchNDUzr/MoG/vGEi5/a/p31rbrmkrJsE5WFN5nWK6QCWcsN7t3t/D3Fr9nGq
lBy1fpBP4r8fFT1/BEB1KF6pNah4YAm3VJHkxTpAO71mPl/rgBUbJEIhH2f3ug4R
XUtmrh/3IRiNp3Q+Z1FeUPsiZuDJx9zbeCVPLdGUdrk02E2HRzkT9OfFIwXV9XY5
GG0rHI1XDLz7j/iyrG+G82fWIaBo6Zm6wdrz4WTxCx1a2hPaJjCZcteS0phSiMVi
qf+RpiCj4kZoaurz21qLQDu2BU96o2hxf0UaE2zW4Ry/tuJ8iP7fWTDfGsS67mk2
Ndju0GYtsJK/fpeS0NshtLvClwSeUVGkUYiVRLJXJbkvG86tNf9KEz/sVvCe37iX
L6BSfil8IfaEyFfn3pzoEMDQVu+mKJQvleC1mjDxyj10lGaCwiLajQuDiQXY4ZyY
I3lIx3zwu6rJIE3qyRnxrFz5HlpXh5Cmc6ABrLBWSNogbLNu2ABRsHj2iln3dd7z
n3w57KtyepjkTNmvuB+31TQVTnL43VixQZ++XcMizSek63ELsc16zXHelRS2l9bc
Q/y4qrQAj2CjhzDkkr6XSp0JlBKhJ9x0K7/hV8n08LTTvH9b3ilD5Mwo5MQXJFch
jv7xq2Din58jbi5s8z/DcpLwv+1Y8hRSAIg3596gLNbULmZbr9CQoDif6hQDN3V4
u0r0ddG0Sp16Wr4894itV4OG0Gtb2vJvitV/4r1zubN3xcewRvIXz842qAafZuQb
LYQu6iLZEV+/S85h/zNd6kgUrZfgzKLNA1q0K0k96/lcjNulTfVk5ngqr56oZGEE
b4c5dMUUiiPLjego3fqU0ibi5JjEPy31o+BRSKLFznJ2a+JupXXKlW7QjOQyz0xV
s0HSCEmfHo4uYFeTZTiwMjdUnTRyYndYgSbOUC5YaRYVswM3h3Euui/jWuC3pD6W
giY6JorW1feQ/hBNk+2cyKQzbtDV6z+94l50YcCjNaOMDY6nHcWTvWQwzIfs+JJv
eQNE+pRFsihlX4r+EWjcxStkI+YPwET4joh/P3z2F2aG8HG5ibgqDFBPiX14pdNu
rE/2AVlrqR90jY+cu4p/y5SCkg6qcECu9YS0AO2gmfohE+y9YfDZjNVEYVBslZLK
KLEvIICgFEc8ssvehI1Nm3xBFpXm08cZScPp67aZbebfqxUlYFx6cyLdcfNAOk4m
83LhWMiYG3mARMWBTvc7kN6GhjXB8dmZO9t6LhJr7kRN6BjlSwafjFGBFP/fC0P4
HYLF/5VATpili4GgLzIPCGpB0lCXDFE3EGLxKABHFCK7CCzFI2axpQS4hkxGzNPM
74T5v6fATBy8NaWjGLTahMe06sho4tzKA8dwxxpDUsI1ConKE38aS2L8ntz+4z6k
hzl+qmIIeuzlk7F5pk1XHbt8cb21r32u3R2RLEa0ATBJSiZsRvkd0qA3sGOLC6fU
1R5KANX1uyefbU5g51WxNGFTU+/Oh6IYlH95mERBZLxQjS6FJAOP1YhzvAuGVvL0
yehVMz1aR8ow9o1rvF5iy+XdCwHluf4Q7C5zN3sClsMm8u9L4EwGmlXVMvQiaQaz
lOE99tM7NVwruBYVArugeb9fMoLd2Hu1PxnYvrvU9f0DagTqIiIF/I4/br0nsy6Y
bsb0Fjqh5r65ojrfrbmLtU2cgNd84qJxE+8Ib7hz3VIO9kbiMuvsYojlM2gcuzUw
mR/2Q8bTRNeAE17Id2wYobxnDr9nmxtkan6RWoWmoTNUVI3Vq1JpYYzVUdGcv8+T
cKcYKRta6l+1CPweOTmmFnc6SChswqHLS2JBa6fzW5o5ZrxiTNe8MCBVV5Tf7IFR
tOgptIYwsgPfv4zXd7xDZlb9XP1pPYr532GphX4JepgkBiLvK3Ja10y0Ejo+lxQ3
TuEi0OWYdw3Cz5ldhmLfM2Q7pE55YwXd+j/yf1YFer5YT8sR0/FUBk9S78BVUOOR
LsCwcmPao3L69xN5La5pg1FGdyj8urdwvUM201hdNQBrv62ZyoO83D6JnX/5Tbxx
3wp5ZiVl750d79o+vM6rbQ6G9RyjuEmkngF5uX/ULpZxBA53vckamwkRx3ac6k6k
BlsDxIVPCGIRPcSSGzNvr4Elki97oU/4gz5vABQwOyUTowNBQ/7JHAqTftoMwv/v
Qa6fJJJlVAw0nE6myJBnY/GxHg4lJFtkoo4BR+4KNKuyewnhuFC0hTddHDphBe7/
xSk/FzrfKzc+MP+zKtFBazlOf1fGaCjKbm6kY7GwwzrfMWRQ6K2cWXikZ7Ez4z5A
Orkbw0Y1sgCxRm5tBxxz8f4O7cQK1KXZ9QptbJhURon7pzP9+waYJJILtDuOoxLC
oJ2HWiejvII5P2eWcnFnuej0sIoFjNQVTdw3sUDhWkfFMfJWsERggtIo50vj7v9R
31qNQFLpOnSEsmFKVzzDVUchatEWhTdmU3l1K1lEK52tig6zac9veGXV63uRJ+5j
zLir/WA+YHumzZoaMY58zySpfCFvT1rOTuq21oY8yhtm53VrKyU6P6z/TwYE3WXO
mfb1C4Yti1esGLbcpNMKDyxBEsF0Btw9Ekw/zjyDQVmKOQXRBwxGmz2IDk/7QoLI
4nRVwLiSj5p25MLwaTxfxShnRoC4z/V4rW/4/JmjthbXYwCtwu31pdDLzRu7ma5l
EjB1lp17kHXhKuP29+KI4bG7hFYEV/iDZk92XMFU7czIeEhK3YJmmwS1gr1OoOkG
GYgL/TprlmKvfZsVtRVsBTPoO5KsNLLP97DUOpaeHbHDz4qZqYh/Knvhjc+YUM3V
DgEqNGg+DrXW+8qdYbPC1KprFJktBqb+d25+sfe8ejbS4fjxKHefKHEMe/5x7eU6
Ddz6+F5GxkORTsnD9vEV6MQxb7eLEsfWtFQTNzdI0okhW4zzIJp2Pl0/9dNRPIT6
NINNr8izR6lTEN429zN8bmmpuTZff1kwgyMxA1dk9a0Cm6tnAQQxoAOq7rrqF49/
+8vrt2tqrXPrZPQz4lku5MK3RIg0IXQWy8zzadXPHu2vg6tIuRgTSyYh9tmJc8Aq
QRQWf1mQJtkAUIQpiZM2aPI9b8uln5eS4UNK+NHCFy3poGuCGMuQhpydnH7RgqZQ
0xVGLW3+BVRclwtPBGhEDM2XaE97tTGVebcVUBKz8NJjwOt3nSqErsPCniql4k4D
DlZbR12bmhKQjxMT/A/3LO6+SMEsqSB/gCgPrQPjp1kTctHL3v6XAeFgvOnQWysi
Nz2/HxIWiebSUjFwNP7aTkAwgDfkB8KiXSv8P7JNmpy+OxcNHjKR9WEh9dYtBfO1
fUvro7Ylb1C5MqSX9cgKym572H5UU1th0Njn2/qANBzjOClBYmogdEwdoguU6/MS
0A00D/xD/PbzhmA6uTTDetY+q8gieJaWslva+LFw9gclVfFO6VsMKfNBi94BBcoG
RWi+vt5w9FL8HuYJwJ0OHTiaYee/fbHepZpCl1VIu7AGfgecSMFKBSvDoh8j05EO
4XzmHMwh7PvXr+dSf+zuxaqpGoPJXkHFdJJ0miMOulGxUTGJfpK3SR6x2tclUjdY
jAXUdWeUeBo9t6WmtI8fWOiAO2L52tu05pqoo4lJm5yaMBcyRG7LO+akMc9Ey8GU
1IigkHBXNcOjrIMnfaTDdZFXGMEzRxV+QBzON1ZxYAgxqJKUlI/PbFIHgw+yhHfG
NsHC/P8Ohb+/PDQ9dZR1JBT0mBQG1zNEeaY33AeN7YZzAN3hGPDuMQ9dNd89BQ67
UJXrazDYOxLCk4RDBnfCGPSZUoc/IJFMkfn/KQxwOa9CGDWz/w1WfNCQOQdBwzuD
Q5ac1riLpJB6YZL0RmrNxlgAgx3oueOQOJRDZZk6xesm25wZTPczAXUIDm9YtDjQ
h8H+WzM93grGAYTtu+UlHlsm4s5Lm8aWPdr5wrj5ci8zYzwwnBRczXHJknurFtxY
j2o8jU+pWMY6O1GKAXxR7srkvxphlTx+IzQ5FjPLLyF7TNv+/a8XCSzZIkj2jfGM
ct2ji06dIUQIljJ7gAhD0PQTGzrsrwWE7TrgT0XSjGcvQgE2V9CzzQXqOdmMF2nN
wAxJFhCL4tiVYAA3PYcWxbTr5gAkidZH9cXBPoTCTMCYN5MgfHMFYpiQUew1xLpt
JxeRUX8tmlTV4Haequv2Qc4Wohwtr2NyrFxWaixnEkNhJqakqP7H3Q2zCnAN+KhC
QaLnM5y5Js0ZoDXBRUTdhrfASzOmLhNFo1QKUXpYyzymyScSExkStt1P8FveVsVj
7TBkzJ5GtvesEIkqy3Fk626XqACdTjYWbEpJT8iYBh5pckASofuS2wRFGmszktio
wczGciT7nHDCOKoa5WhaDubCjLXf/6HPYZKMt8GfVL9NfBGpLj6xq/QIZbdrO2/D
GapFGvqmxyf6cMkfkTe5PkAPzlCglIW1gVcBgnMSWrbLa+fnPEhUgY8MioBo7QW3
DDYvMDznK1GEQ9GTAue7fBIfv3JOP1Td8agW9Jd7NGNlQs0IuVq/6Fh5m64YLPpJ
925Lwvb0ufmSH4jbX/9M4dM42osWzRqvyzlwnU+CB12U2UBxFQMRy7+h4gwUSYI8
SOow1V5995gBw96VQhSdG7VWxsKz2MnTw8ew/3t7/90DyJiHTVS4wgoG6nTvWq3+
yWTOd859hBlJ/aamiq9UqDJNxdFWMU2AFTdHmfxez/DFH9zK9HRQ6SXLsLF+OsAd
EGrHxQawGx9P5r5w51Iqxz+FLDYfnwLDa8gOthitw1cq0lgRvVOJlnD6xvha2pWC
/rwGgt3D67NnWGDSaLBnZYl4d0OCWkEU+SzVU7Krs/WAE2SjsC8NgvDCyUJ81TBW
y+phIc/5guklRocrrWPAGTAHDlITvkXnjiDIgezChdfYWU/K4DxpVi/GfQfotBOx
Jxb815bfX9xfK6jQueJF1aVp94w3Ip/avOG9u3cb5J1MPtaCDZ+kdVlyQEAhU9nx
gEhzyaRdYeuH1cvXvKWiG9Sy/6VhL4C8jcVvlZAuAJ3x3IL4nH6vo64WChU3sVi9
2fX2G5FUj/YdiOsAkf7V1UaOSOQDYVP9h8FgoTBEqDbVbgiJNvrz98snAat8GgJA
Yg4iVVNkQqz4KAxUH+zV4CeCQVeCXXAIHRB2GGiaTTCCANexjXVwZHU38rZPeenC
8MzZIJaXBDlHOfhu5b1xgUpnSiKzxUxco7TPCD/GUX8yQVwZ1MOtKNz92ntnhwgK
kFJLv6a/aPXYZO2tNUleNaubcNy+E4+GKG41EwAMaHKlib2CN661a2qFe2mGzr4f
LHERuyJUjy5uwNvSeb3D+N325lE+8rfrrdgHUZi7FeHOC6376sAFCh2hu5/KYYyZ
7cSjHgXpK0qYa12LDDTMovHeC2QRAWDYU10Bm1LAkE3qKPl8zVtZx0duox8f5B9u
hHJ2tzoTbA667AszReteUe3iUAga9kB1gTBHYIcWoVJRDQwHxDcvJO+dOwT/VG9Y
6WhOdu3o7iGH7WjNOqGsMGsPZPH7TY1BNX01vJ9GJVo8Mb31NQE96+AbO7rqf0Gn
W5ZWQqtZ0w7UpEZqPOYLkBJitaTGOfIiSQSpNd/3PkZl2rT98IeU43qAOGwpcNNy
Kc/dPUwn1pICrIwA7SLSHy3aATfTcb67apurcxpxgApunifLQtHtxsrTATl1i9Bx
pAi1wmHPWhUAeSLtLv5y+dbeDyU2qEyCYltmTrzi2G1UEoN5fQazY/7dmwEeONS0
SixIWNFCD5oJm8fav8+hbhyBuDDUIyTcI+csAz5je+VIYsMVcjIVPCwo5+axvevQ
Csu9EUxHvSMf8nBPo2evSPpaKsnOcRJd+vB/RMrTVqP8HOEByjYGwaYtQBMabNku
qST3uQims+D5JO5lX2Wt3yBmOhiMRZRAP+X6CNXXIlO07i99/HnmGJNnK36FEyFA
iGs2YFHCD/kLH8LQdUSnMsbhMvZBhEXLjCQD2qbBLRKWo7d9vyMBU5dGaoOntMPH
Bpr7QD/qdMilzkLZPooig23o73DKIiDmgMpF4GIHJV8DiYecvCcc8RUC+ecxbIti
3wHm23sjv3KF1xC/dYThWv7+KF53gjK2M7X+Dm74IHJZBVR0BcmtK/hkoVglaEh/
ZtyleJPrL0ZyToIkt40eBLEUV9V2J1+iRh83n4+QXUc2BZK90OAI91RKbwEDXp31
93Qmab/uFPtYCeihTTiEtxDYiw3YpQrhzPEI3t2EHJIf0hxX4CR3QuxIxa8VCAAX
ILoWVvwv4szyU6VZpKJQv8PndQRaI3RMN1JIMcS4kkuez4chWZOJx6yxcv1rq/lp
GqRZRyu9Wxnk2mIWuq0kk5DgyPnNMR/BHGYjtM1x/3kn3xHGoLj9iubPv6y0f/2i
UiqfkFe/n7o4iORfdf/l3x5faH5b3r7kDpsaOofNf6g7eGJa4l2T/Coo3jM7JDRD
GtWaQddO+JypkFDHxISsrMNuvnHQrNEJJk8SxLxMMmiSfEx5yCVVdFWBxxT4p+i0
sLHyN52Xi2FdueWhHs6VCzzWD7gYdf2V639gh3NkxXHL/OJzt65gdCxiNhH6VZjK
cgvP2tM2m+1WCjeJrc0h/hdDRbJck/HAseJrE74E5x0ozE2yLrNZOCAfzA1qcxaX
GTePdGxhQWAShF4fKlsdh4C/HDe7UtypgDVrnpdnWShJSTtvUuHaVMEhz1FN3yv6
zseY7t3Odajv3IO0xIeDKUx6XydULw7le2jEk67drq2SmMuJEMUX1z+7uuhZZgAU
oZxsSyOUWu0YaCJr/z9RSLv5Sw0Ue2tTcX6DoaZdKuppOEwzA0jk57+yQteVSpUy
lzShb+Do0BoqhvTK2Pm6rL7PMS7rImtGz3Sf9vD1EiqhD5D0WXi0m9OqdZEAGFGB
qqeoMiJ5Tz4ulADxdenbhLdhtsYfzhpFXoqqIqEn/00aectNO748lcxbX6hDwGml
grkwggA10D99nAIUb6B5UTqwL+E1bl1jo2PIvTw1FgNU42H27+Znv1isegNJdj0U
XY1ff0Tvuh1Jpq8Rep3R1R6ae4CgwXLWp5GsoV764BCmOx6xsnjtL/Grx7/HpN1L
7MsoMTZxVHZin7+hCffR5cPXZwq0aWmHE8mrbj4jiiudXPM87QHaEjTVmEtgYC1G
weGZU/VDPRxcjSjwl7kUaPQ5mVk7KQHgZZEI3q5ICdB9ltUoHBdb6s9QCai83X/R
feSH1YBuCr7+oYvnwg6VMKAbH5vN6MFWYANBYVmg0+nRqgGd/OxYG0c72h2RH0j0
YAELidCHnATualMG8J3M+F0xNGYnAqwmy1LwlPDpd7IAnIBa2daOkBOORZn6s+1Y
DRaeyBT/g4i22VwFHsB29NKT0OQSNLdTyrBwm3F/1e8fImFndNO9J70JcfzFAdza
/W7rIck/KdwIjhaPUOPefheWhELRs+aahT08ebgd3+yNlX3+AK2XBUDAa1I3+2oM
nRA760u8sTyFxpnLwfMDwZMpIOcmk9XibjYrsTp0Nw6zToYrkJIu7uqemVTy3C5n
Hzm/Pvi9y+sf8JXSG+Qj5IGbF7TAvkU9sXE6LWQQkuKMByUw0dI90d0R/yhdGIfZ
HZ81ya3le/VytjkAy9LdkDg+8EhQTR5jUHverJ7eMqA9rSEb3LQZ7FpMdTYnb2G5
YUjJsETvVtQRcUZebRHlceRyqfxtqrOO0jlLabkuwPcmg+mHixTkboicS7cEA2y+
NOJ/yGNmiomn8kCoFp1FE/V6o9Mcxh2lrjrTZMeKE1RWlOUHcU1zH8KJpxcTALis
kdMhJ1kl00vv4uwsub2hNdBPWzawUVW/EE318lJkKARBS1y/4qg+uuIYnTPkr8ev
Z0N2BHSUc2w0+gDqs0NkXtsuPA4dZg9UmI/Kq6pVJxib/bz4hmLwiuNMSOPDXvZl
zkwQ86VFnK57Z5U5qRzb3RFN8S8kEHsMEAqLgKWXmQSvHLkGA1Jq7ZOtoUJ5qOIu
gQj8y6iWxfH2HhavKTK3uiOndnDNELxHu2M57/KxjOBjoQlR1DtMdp8HA5TKM+by
D2DEpNDajAdI4micptZVWGqxYoXEda4SeyA1u371BA3sxxeye4zWVmMdLCnA+kIX
tOHK5HBSt6+anNjRy44qGaIg1mgtEL7kTEhnUcRgb0ftm1w3uUBLGjO1dDLTYLGW
j00WwNSWTgkkr3rB+r+RSs/oZH/P+Oo9RP8TCjEjpR+jLW5AlcTr2D3Bk6NnbpPX
+j5kIOB4gmN3AzngXV+u070+0aXngz6T+O34b3L/iz8a6/G+Y3WB1sZAqsZvEQ22
/J9soclrjkGpf90qXRjhdZgCiLH/V6AsyI4Zuo4RvaWmtE8zZITAx3/gHT6m3RaU
kUYFIJK6gxc3HCn67aAaNCjwUzpctkARar+xKK7fjfZRftCK1c1+HFiTmFyJsdTY
CTOvdRnbhilT4GF994s4EaRcIF4cY3cbSa+DLSb3TEF8v5feFoJFvSbCNP10Aqwr
Zd6bYoW0HvchR+CRFL7eifEGb7Xxs+w+YI4wjOo6I8iT52M1tZwfQl9D71dmKwqc
8aYljN24aj3CkqLCHgt194ZY+x4xj6yz4sFqY9Vbe/QWMEEqyi4LTXCwETueF3re
I8fTh/17fhWx/kjtlIX/i8r/zo/uI6gKZoQsZIBEvOG5Y1zAx4OVTbFBpfGzH+sN
5diw2uWHJ+d6PzZZ+fGqnPUYEwT6lrHGeD8+1dWSMYbrraL1jDHfAVG6biXD9W/5
w6PJ0n8KXxoJDfMbleqTLMCGXYTr1PpXSdmr9G6dCpq/o1gS6VKjoPmwdDiiJ+1j
86DOUeZ+LNEmrxoS1irAkkuLMVLlVe4MYT7O59BmNs/N9LZhRRqscJ00yk1Xn3/s
mabFDmcFmDyvf8eCyeQZjD9KOr3mKB3KzLZcjvmhpUac0kfY/inpsj8vximAe98P
cyk2OG1M+r6UOTLBzVJItwqg75iavSfQ88ItSy3jak8eno8rIePNXO2ixz6xdeLP
DxZ4Lct/N5TI6LQLbk4yAz3asfUeMoDfu7MZHGjBZ+B0H2P2KXitnbR+rOhL6K/9
FL4fCgmBvn5IwF7qMkmZjqxumFhG1lbkAbyjHkPjg3IFKLEDIH7r4QbaTeO4jifk
J3s4Fd4VaBEq/fTD6fldW0j4y5qUJfEZGiueT/TixE+92/mnqgzC98UbgS3TsdTe
NJInt7ovD1Htg1ADPxECHtJlFAjf7kF2SWaou17JZspHQEUkW/6vc+bINRx2e7Du
sMwyRfiViOcwwT97p3mhV4DhHIi34Gfe0F3Bmmm4+8lFIisANcC+M2WBm18QWuNV
+XZNN6e1PKLCUBOOOV2E19PdATLTfG1Ek4/3RXHoHzybU8wKehWXMMxW2Q65YDS/
3madyoKGrxmC6QKUdWAPa3o83xrkSoiP4MhrgvNKafUNfbO/FxEkQTHvVuTsfFnl
kMD9YHV3jBrT5f2fB3yStV+fltLbZzI5u79qVcToQctq34JkzfqMkHuiSDqSP4AY
6b1KmOIA2MWzT5NA6qviOFA0ZmTnllGCDFNBGedXfmIjec0NbSXOEK7gJUyN+HiB
8OmAAINQMCLJaFLjdkxzBWHRJMLKM4f7i5cmJl6twI627QSoK3HhYegygnZ6voWo
BaIHQM7noue+9gZ/g0QtSPtPRslzERmzgp5VWJ13lU0TS3TRL7V2Czdqd9FTORH0
/JPB4QHJiCpXQQd4mQOPJHtooPNwnHJiCHOKpqOhDtq3v8CnMH5aMqPYFb9kh6KS
em3l0RWG0w5L2NmPzXMW5BdNs2BgnWkHPqcl+yiddqxiiXI74aMHjPzsuOkh2BCS
Q7HSyINRYo8GLJiPBMIQUaSMuKS9QDTUrFYQkBmpCdFl9NV5c9R5qrQOlQG5vuZ2
zxZCmH6vzAr6ulIZh3gM3nxgPlctOuS4PaEU2NwHneelJZx4VHxLaVbjsOZqB9Nz
z2sGtLNuieR2zKmr+ZqdFCddUDH56ev3OfJMd+Kfkyjm+mD9TPFH5Bh/lBlbNVgf
W2eho4PZ1S7NO17d/fq17G/YLIUdmlMk+s24nuezhwzOf/VSwf2+BINFpqfpMCKr
tKZRKLj4AYsok609zoBCOw+SLVPRYm4uzQkM0yqgZZkICyycyDA9+0t/MzP9EqrZ
T9tTI4NDgvpqNnecsaaxa8jsNTSY+LvvwKN43h/RhDWWu5nWf/8hI6LvkmUibUUq
Cffdqask0KfJDevy5pCjfltnnEqDtg875ocarDRT3lKS5dkM8kxBBh/z0Qp9zQnD
CnrR5RPnB3FXyPTM3k+EyX5y3x5EccFwtGpQ3ZufCo7zvK6XXWA1va22mGf5hG5k
SG4+pIzVUWA/vLlGSfUbCZWl1B8tu+U50u6lrggMnAcMwp+aItpOvvGz06X5XlJv
niacHkwm97K1hcKCQaDhYeEDC/McuwWoKE2Y2D0QjodHOJK05sp2UDUIdOSbVOEm
N/4qtRcoDS5LlU8lg9XVpiaPZfg5HgUGY4O3YgIiUhDN+q8EJ6wZPSIB2QwiUv8J
0Ayi54r3H2gKhVWrCV+8s6YfyfWlz3HavG8MNaMuSTdI4E7TXuspwczIPUDsnpE3
V6p4dNKzS6Mb1HriE0Zlt4++arKn5hnrBEqe9qehdbzMbYQzFiOJ2pQlEqUeC43s
EESf+IsAfKoynD7ehD8vZ8tgZpbGJRfRf5PJqImW+oR81xOy5HnUWpq1oiZLJZZh
slFL2el2o5aM8oUdlr6JgcUk8UbPxqyavyU5bF8jLfR31vm1QbKVhvjuLyOT+Jtq
eBTpd5OcJ2vVeO0RtXpza4cQDUWk7uTQqo/e5S/+FvgP9tOSIZtAtxV4pxWCBkBd
fCwvfSefBjZVYSj8jeCasCdoUfnK80kTF/0MCktU7cBX9EMYLyvvdn1sssFpBJVX
DlEkByk2Y6X1ODlTSjccIw/UPgto6DpAyCE/20loIROLLyLQhY6GUZ5305A6QVOg
s+SL0APyLtgWDCsGTV6bc+W3mNu+ann51FT7GR++B/2HDfLSzk0uQHFAdzapJDR/
PqlfMpj7Fs2R+HU2Aynuhd1IiaqhPSEmZffO3T/sCBDdkl3IIFHrNODwilwFgd97
DJn+0OzZScScxVzIeNv0Qo3aPrBfrZnT2yGsEbY9U99wv/4uyT/SD43tycFgrD9a
5CwxxZAW/0F5Vh/0DjG2ccEDKUP47FUJsmtiKxmuJYWSSUGBbgoioPS/pf1PLOV5
w8eZqOiBeALpYFXueFBEOYxaUIrgzj0E1JdP6aPfssaPlAR7m9666yyIJbNMjUgQ
PuUQhr0Iqqb1adw4RnP9UYzmcOwq38zFImYTSrD+AT/O0tQfnCf8xPO45FUDt1iC
JQ9AnxIR0BGX4QKrLX1TkLP+5ujo1f/XSxRMUhwTVRFFqhgDu0siHqsgRl7I1bGu
PmMmxme7SYYbInLBLuP3m/EJfC2xp4JfuJ6WTb8i3vsH8LpMMOdUwh6WM4EZ4zSb
Jl1E80j/mxX399oiZ9DfkHusT+5to1tZEZY3y5ADNg7kUxDIoa7UNFi7wXJw0A3f
bSfzFr437+BTZMcKaGL7CwlEVjm2fDTvVRBJy+1kNWRaaCYvNoztG7m8gBdgx+z0
+uFSwlO4prE1JkMKtcbWShjuuZtswwN0KX3+ujUZowCiSQS6K+Scz5hdIkuOCyDV
WyqhnO3HodL6J8cpZExvzN/BFKyXfJ8UDZJ3zxEnNknndtPOPsVB/iymiiM3n4XF
EEVThSmJoulnGy9AItyg/VhYoxtZzRxb+1fi80b6JKUxP3+wmZfo47es0W/Q8tT4
3SrvH6ZcdHXpcbyiz7h/NeROrPY9WEpSgpCprbkmlHf9ShdVEJmHve+bXu9/iEWj
w1k//dVBzVyTLFl+/7By+SwZQJqc9HUqqD3T4ylA/i2kFo9TfNt/MRuNISGzm8tq
MmPpP63zZKwAfHmkREN66xDERLLmXtbpNBvlDO0ND9Pjx9UTcOUO6IRwFrMZwx87
AF2cXiBGTN8QZH8X9S/ggiIuAoh2phDUZgm06pX/yi/6ExiPB5GzmIwYG4r0uEoN
WnfrYPQgLonCnG93O1iM9rTUdx+YlMVjk1xVSogni8d3xMVClGnhAJArNLbxhyY8
M63qxliKRq++POajbUqMo+29/2P4kHVohs1/Fngbz3lshwYxl5saGZ8AHqJBYQ7q
wjUirvmXOVNGuHEzbELl4LjPWrPnafPsEhXdjQRWfnT2SRsi1I1/7Mw8oxy57V5C
H2zsJ2ss9cnh/yv22rrxlvI17HV1GUNtXLFkfPgTuRXKdNczlyGq5+4Z6WMZN2S/
p7VmOLQgVdSo7MpiEjvT9edhX9jIvxTXGAJOCS8XBjpiTZm8JTOIAQnMJTYSIhEW
PcSUyesdf+/IDxNhr9V8c7Q7pvwQZ+qeNSzRKy+uCsWFB0aLV/iKgEOi2CCVTyhz
qJopEQaI+B8xv04xozu6ZjChz6IWXwKItlcfVIbsvN8+MjEPSl2g/pIsH7PXNUD/
WwJA4FV62dLpRcz3Q+ytTdFZhNI0MkdxYZGx9i1NokYd8B8Ohos2g7yEDGLpQiAR
VKu/ggP/UEKaJuP89X+Txs+8QKllVJCsfK6FIiKKfHswGXX5eDFQu+xx4d+ueDY/
oVM4KFpV5KC3LKmpkW0Fyugh/ckN0mHPWx/pt4j4PsKasXxVND5XWth48cwhlaOp
8odhZvtLWhUyBHRHYF3ebW4gffj4D1rjC23dt7aBAFWs6yfBDAWzWDAcunezfnB0
tbYn+uEqhwozPFbWDEOfMeLCX1FNFPa5vzL2Z7MYmHbnbMTktYMQiAkwrfRsqbhP
7q3NIrPQH/BdiodlC+K8TTAp1ZfiWEGPsM//oYJE1xWTgBoarta0s6w+e3z2E2d9
6LP7prEbSftJaO9vnLUWsalr6kIkEi3XSNY87R8bRFkfxsQGhT9PlEck6wn5hRl6
Uyyeg1bUz/oOapYu/4w5/DegmToZfNKhXrmhbuLTcwmi1tcrta5/8LuhfZIS8Meg
9IBvcaIkru5W0SIjsJjqmzU5bsMVyZDGntSm/pWCbsaPh8xirJPSwc6+KgrPJn61
+n+T+0XrgPIwimLrU9cDagTcbRKQx6v6qe3HskalPKsXRQreT8utuTG5K0f29St2
HjS9fW40VYQdFm81xUNPBylldTHnmNl7FYvd7Wv46g+MGykEPsnwr5uhG0LGNV8m
JFUzy/GpibXykLLNCYmzlR7WKqJwTJs7uTkMzNrSupLvA/qExeMgqma8Q+OiTUj3
sObZthghWtAWYzmHxrd4TO8pKpaXRtE6ZxPmz1SOYgw0k96PQKPFwT1HcsrUupBM
lUK5YtYfCuhggLZgR9Pq55z3J90Qy6qrclUeMDU+wvUstJRxvhn7ulxotv3PNZfS
vV27Z9FnhOTHIemM4OLVng3gDlVDfy8meg80bfeUg1EqE5/qrNgk59wmpgmanfKW
SXacx2eNj4ESwelTQm0To4HhSrhQUah1i/Oc5SqJBzAaQoPetoEi3daBxopcP7Un
WNfQWISd0Yd4EN+geDDN5Yc9jKPNhqvjxgDxtntmdk69o/Dncw/UfrWRN5k857kq
18QK0BGmKRi95rjNlQmXoTqJVHRFUDY+2FYenGjS6A4vNcTb4fho0gSnQUrzLis+
5DcocfsPnfIrE/Q4S0Dul3mLa0vDDEA6S6U4x6OFaxinHAOM6wjW9z4+RN8jWQpA
ku4VaebxVmxKfRGSEf2HGVk9YSu8Pl/1V8gFgMPUdTAtjXnRg4jBjaiW9GYFrDlE
b5bL1N5Rmy/mRcyvkZKRrmykCM4cuUL1ot7EoVW/0OaZiMJBsY5PwkoOlisxpXfC
vWYwPnFZ11xwD6SEVv2XQV/YzVi7haF2VTScHkijvO6E6LOVfXbAuN3BF/D5AFM5
+rTHJeD1if5zqHc79qCtNSYo2YxfjjnQJ3eX0hKCcP/V2i/9QXUvaCcTWcrdIRXz
5kTVW4EDsK5SJrIAkgNOEk0INcFiBkyuIqh/p3G2IWkk2mxFsN3gu3OVjsWdtxRN
NSIGO3zi+KNAkmDWbrRRf5Br4MDCLdia+IFllWPYCSQnDxbCJtirOoJbunQnurXS
Klg3IU9SZm0mNwE0K5+2ATPxRCy3xASWXppzprLPuQ3G5ENnXdsVa431wCapd7CE
uFMuKcSqXMSt5bmcq2NDgXE1e3zIxcS7+3xcA9TrDZFJwX30hVLT3gAwD1esLTGy
5XkkKtqg18PSU87RUHtTtu8LVN7t6wDry9QA7GDO3+KWljRMo9D7zUDF04D8ro0n
U+072h6PQXDsbRVDXxY4JFJTPlM/30lzejgMKe9PLE3c7dJp2I6i86UKgIEgQivo
umK8JzK3TRF3sPTa/UgaOS8S7yWAsNnqShYrznttPPqoSIFDvHLW8qkrf/Zoavd0
OcByRw/qSCulE6E2OjUrDyxTZUmPoukCluDQuxgiTpCIF5lrgceAFO7g3qGjxEPi
7RjjlSmKeOsYnrfnQ5zG2OqkfZkBZTcaDobiF0QMxVmJQpyfZMx3rIbXc6+1gleN
QJf8a5UUKd5hky5nM8KnUZEiKCDoOstML+ZpnBKXDz/ma5DCbVSeinOIQ1jQi1lH
wWM76epjmn8IEJDwLRNf9pklJvZ9pMHjIi29HF1aM8y0NJCNNv3sr4OC/3VpH4je
kbsW3nZkQDs4/6IUtiafRJNe+/jwinkhYtsWre6YRK9TuUjx08CMHsIh0GdNFP8L
it1dfJjWQAlI3eF7jDhNP06Vl7scHvPWXOjpVqKGFlxf227kjPWtMFjMkK1sdKEK
5oxp3x0IpNaySC4QwkJnWMEQAzu308VkZPkl+pDHkQx5vdDlKIu0inUBW6f5IpSA
DQ9evycgFP9sk0oIcTeLmryXnvUbH413f2ZeEyrEY5IQDsunuTKKymh+R9IAQdW9
Pq/IR4gHDt5EPpttRFGN/SP/82VOimS3814n6fqWF+yQlcbatPFZDfxfIVUinDKW
AQbeyqJnGR06x0WMlQ8hKHYFZR22kVlPh+PFR8HNFP1j3zQa+QbfLYLadiyxR1sU
I5i/iHrDwk4bJcAa9NQ7XAqBUA/X6byZazDDlIGeg9rFXzqKGWj+u04/2yOMJ85e
llR5A9ur3JJ+XY2Uxle+aBmVgSvdFk67OLvYaUMVMPb33pGdCVGDn4A4bkGKpoaR
WEwfj0eUazxU7hb/jJh99Nannkb14rTtprsjqjgoXmHZrRUmxYfmm3mzN4KW2Q7c
e0dYT3W0BTD7fbQw1ZHp/B9BMtLfGsGsITu8oRL6OnsHG3BBE/ufSUlaTzlDb3eU
DaCUi4pPhuKNL5YnUMOfZRKhlXOACm1o3NbxCdo3AlD2JyNfXzw56oudlGZJ2Wk8
5KWiZPLwyZwTBc2aICj4nsJxKiy3CNTZ4S1yhgNcuARdplDV9rSDJN6Tmvn6I3Hc
oFM8lLKkLBKh6zFyzrVObQnkE+3RRyqDIiNjgSdpXte45jwbM4US3XM+3/XEUiI+
RUim59CdwqJ8ot5KTni2mzAJfmDyJyjFSN3h+C7kqO3pJpP8j81ZP90FBY/HRU+0
AIkJmf1WGGEscM1ovYHu5BRbaR3r1uQ6XPHf0DnRW/HsT3G4H/e33heUzTjEzZ88
Bt7oJYdY1IST6JRqITj1ZdsuQ4G8bctNVOQJCVHRnbC/GTBFldHdQVG6NNjtAs3a
cjg99M2AUlLkSYR006s/DWKKXBga8SSbuY3xpBU2FN7UVh84mN3tgUORmgDRdvAO
EruY56/FBNCA5zqQFdoQrPg59V0DjOPFHLTPMjVb11GKQYwdLHZSdHK+SXYL/nQV
PGDQXrfjikfuHzhkX2j3mLvWB8MeCPJIf+r5LOAhp9Grz4fdF4iazUpNAT/7wWjV
UwcX07BPiM2TlhIRjT+yDWojCbHFvZEWbRzigxxqMCKlFz6cqVNjYLq21L4/LLr7
fdE067npaXUIAuKtB2M+r6kD2mI4f8OtLuK40iC/cyIizct7wEOFP6+FFeKr7sUH
z3fdUe0NYZ2/41Zb8gO1qFVVeL/fZNzNOBtukRTDj6rArxCbkEhgX9uL2ITh1qfs
cY+Xm+4L8WmIIfUV21m4nxp6XpDasyV29Jb/q/C0DO9G+ApUuW6Vca3sO8vVpcx5
hTlQ2QD5FqYdOybWbwxyQCFI1dXdjMJS2IdO7imTtH2eL3nvehsW2d69z3HvjC0e
5CCbPDGiz2Mswg3vTdYPkqQoxJ6pnHBJTQHbcKl8BBaYQCOg1dudyf0e3zbgdSG+
9Hf1c+3xaiXL5xhIDq4rceBDJD1oB27/r0NYecTtynR+dFseLvYg4bqGRuFUFkXY
d02p7RzoK749AXGODYQU8OlO4n9y6x92DW0n6oztEjJHdoC909rBlt9n1iBT6npU
WEPmeSF3mQgHdFP25Ks4sH5SSBJHi0LQDj3wMC9dwPu/NDsW8ON3EwddOpIPxXFU
vklptfp+yERakgvyO70xJ9mJDkk55DF4wzpFrgqyYmfFWyyFo9v6AX3HKK8N5Ppw
X8cwhmDKdf7DNlOBWTPH7rvPTtM9jYxZf66hDqVNZjiAfE32k9HL5f5qjCul7qij
Bbgvwc2PKjzT7JPw7QNGgsxnt8n9PVMPeYuZFLnB4hb6dIEhoHg5kxY4hJbzwBnK
hwr9LA+I7N8Ru+KWcmqyGGrBuNZCCvfRyFGG696zEFgHW087PIkgLY+1Zvob0PoR
KK/E6bSQNTjphzTrHa/3Ij2s6p9mfWmmTYARcMrPCBkeYASlIt/uPiF/3UXX+eO5
BfaShfHotqMLaE5xvxp7BzQmbFcYgSfIKBfurJXuJOGmLxSrvvTEoix2B6Ekg2Lc
eT1sIXp1zw1ZY6EVuISFkkW39d/ZkDd39hTGHTNYzYEmaUreDIM5B3Vr9yCX4WdZ
CnR2qOlJZRuPa5CJRJ0EwUNrA6xl7yNKYftse//fuKe2o6L/PltTgO1tkCFlp9/b
RDeml3ubD6wNrPeGc32RsghphMUhTQxO59mwKNxt72G1cD8/FV3GYVLprotoCja0
CvMOA/TLFh17o11vw7iypzx893tXGNctXAF2Qs7X+NPUYCzV6lseiumEI1p8B844
K8c1F/3qpLO6+EW9sTj4189jwAkrheQ1502763/v6NgOQeIp0YFzYDYwi91v7p5G
RWWptylFqJR9KkqxYtNjNvTMRCGIixTOmHV6hVSbuctUVDy6lYamgy13WahNx+pO
wvHCVSBtAY+W/kD5yMBn4KPWpdA7mHWqPN29qOfaInqpidfoAaa/TwXjMmtY7vVM
mG4McE4rBUwGhouqQmw/HJ/e68i1p9ihu8Snk0ogO5TWYuJ9ktZeLwZGmHTOvMuG
OD/rZTPXA3Od9l5JkcloLdTQN8LFxwqgyYDMmrLmGJO6OdC/V+2WiuG14k49iiZ8
RsfIcC6WH/nEmflw1IMGMLoAMULEbrbPRtHoqvsWyvGsOZzs9Rb4NIMRlgE0cogi
dnjNC4xArSZAf0MQPniDCOLJjgCDVAzb5fS3l0POlkIyEpPv59Qzn2WNWrezl3pr
QRKPMqwNFV3gAXWGrrGuZuZF9H1szLSkiQgk2o8++iaIzL8QKypynZVPhm3ujnY9
Ntl5r13Hb4131NR4PR4aMYCxK8I/l12p4Qz81rQ4i6h4UMb00FPZsU8ube0yhKF5
4SgnrLZb7WBqZMCs0ydxLjb3aN10UAl1QiLwlxoBu5Uo7RghUKjhffv6T7kxNgKm
/NPq/6BBjUZk7utgtqEEx4tLivZRlyg5t/Q5m7YansM8XWehPwNFnPvuZGXomLot
HV8MAeZULnizUfGs3PK/zSrfEvxsg7sLzKYLEmIsgelUZnTX2GKzsRrLjiD4K9J4
TiGGatjV6So2FN0BHkRn8f0jCGQAP5ouYaimxDtdIsA8drgygq9N+LPiM6hdSw10
TLgEcbMm+Jz3VV5vMadldS0hUluSSyB7EPqLEThVG024H9loLdQNGBV+ySrB1N7f
GHscKuHcSJKDPI8DoyoLbGaZcixOtdpZ9H/YqL+vg7wvnVW6MTipAb2xLzR15xGn
Spz1x4NAUjRduYvIkQXHLApbrO66RCOYSxzzgXPntPBc1o43j/OzSxPGYPgYZL5J
9XA/NXVWKeDkozzGCiMxBY9vG9IUfVRiyBW+iBOb7+GnWOJ5UZXpIgYs5IPg4H+b
WKnIkhof6SMmk+3K13DdQ0sbnNONI3sKcZoMjLWVFT6Nl/DWJTs7JC7c2yR/v/WU
l+uGPAAr84YqfdnPP/3FwFnqOFkrupDNq6iMeanlsZ68Um0+m0EQNiafLWyUDPhL
Yjfapp/8DEqpfXAYXU0kvErzl3lEOmDO21/01iFch13VK7iGdGjLQ6Yo6GyC8jls
geKp4tiS6QPMNBerxaJR0D7W85WX4Sfsu9xkcwfg9HaBWLBeUP9SL8Kjlk8Zw285
19hzOcRKc30vhC9cLRLLVfbAMrNvTlYYxeWGdFZovu0qBnOc1DrQ5bbwwsF059TX
cxSzdhggkWsoTsf6owi8t8VaoZpC3ChZIEQosx0l22yDec26F2wYidkvyIawg5Ui
quluqKX13DFY99v1Y9DKWLkbJaiqH36Lc4/BBg3WR84ggAbUIEjj36CilW1oYAPx
/MPekG1YfvsFpVVuC5eMLN95cLIdkKzIYRkpM13ox3ZH/+fSjgBFzhDAVBS95fP3
M9MBho2a1Je0IFGZz6/MEwyuMQJUiMpNdjGaeLV+DqOeyJZfOaF9WS9OPWabQtnM
h5C1vGDMpjK4fcty3I3lU/QWkHofmwmL7sYOsjIj5KlvnfuFaIBDomgA+X7UCkKX
ddx5uyUCvDWKxyCGUSJ4i7HVESByGyEayJt4ale82LE7pJW8aau1twCk76nVvwnR
3ZVVxRwsTp3zt8alX94nTPtolThY2s0CRo4F+8Yvpze9TzCoqE+PxnhNhELIIF0m
yRWZ5w+u95n+TBuywzKtwqiT2grfqU4+Z7YjY91it6Tzs4sHPBGW+TSv2kLr541t
a5ohKEqceSY2lbq+U7iMNvB8dliC3gLk3Q63VqUDsG+XUudg3GcmY212e4GyKork
NZle7/Q85LK+KMEgLdfbQomaZefrqR56Hh1l76DNIOnn+3pW6P+L+xwaBkLCW4bM
2Tyt1WfQyRPcyl6pgt9GhdQYF1ubqFiGjdzO970SYprO8znGrOLgfRLWQLTAtXSA
IgcKM7atvzFxV238UOpQdyouOGEVDNDPYhqoNpoG2UbSp87W3sqTzB8sRXKxMZim
i4D7z0v/PZzTVaSf5Lhz91+25kYaRW1NOU28bF04T3gTcToo8eVsgRHo6/LsCJMt
DvCNh849Ugg9nOabHHdFgstOMBaCjgB+Y5fm4zM0Mk++GOBpya/km4xxuGO8YjvS
CVZX6NRUhDFu/1gOsOUJJ1MXqGU6TGjj8GnlfE0MQbkF+6Lr60iAGomTEJXIZvJr
X5NMwW0c7/D3FLwEeB+03O9g5GxfO4PxL4J3L95x2OmwzVmTlgm736VbDYz3S10f
bOXuE4MCN7LpSwcNg/E8aHwFMeoI2OlWlTZ1Va3hUtW/QR+u+Yd4vKvZTX5ysVzv
Eb92EG9Q/aJEvpXIop8qK/prwkIsG8QWwAxrHFtHLK87lKKFA5kL6yIX6QPChdUG
56Otj6MXUcpZYB3tnoCBLqqCAnZyIAvGtFhHlkhtflxye6QgqUq8aDGt9gJFW+pk
+eTgQfnclahbT2p6TnDU4KYZXD3aVJ/UyXqX3eMPhbDHiNW4FAtxnQctxRm7+ksj
ct4inT/ByBJrt4EzCp09PgO978IZ/DHtGY3GDhRlO8Hss1Hz1ABYdKf7Yt3zIQL6
LTqaRfrTCEmlOTaeqGDRadCj6AbazIYVOqTUQc/YHpRIoOv/TU7KRtkn7ubxRqS+
fF6x6vufHPeEeyW40v6KholfCJU3iLUprGLc8ZHwKjyWEHt2F2w8BF8SpsBftgp3
Abj7GLYiRQ5CZAd00ObBMrN8tlSlK2vP2QHWTHmiDPSvW+5X0MlPJGGYX1lO54px
PcG273NyDTXcU7nsQ20VzSj9QHhLAffTkS82yuD8LxtfEok6iMFsTi68VN2hT69I
9Gnd+kgzwGiaD+egAHSvzOG6uKzsKDuNAUaqh4LnavLpXpDstRdfF6m2l4WgS1JT
ZDanQjpk4i2OlVLVFLsDf7gJRjIAwWrB39T48Etwg3Fk6sNj54b+7LX33sQC9YAQ
Ef3QZJgdCacD12DsY8mL5nCry6HrTTwUVut0Ayvjt3Hfqs447ab3dgN6ahastGaQ
1mqrFtRxsS6L1u1AsReyWc/oR7N3sTwi1GoI8muoli7EBZLu9dfs64XQDS/HMv7v
0DBRN0Ixf1ZWm9XOHC440ELShd1buMds+98gQ1Rp9DW5omSxja3j2CL0Z2FXaRrX
llqMiYsC/HfCJYcMPwmzqWER+2DtfHShxfRJZRLla+A3yy9wKgCeBI3qSRqpcNWm
AxkXEWys4O+HwMc6sIu+tw9T2Mkpw35ersEkYuY4Tz/RSS5GpOs/lzk6VPGLdzAC
yK8ze9l1YtD96H2NwC8n/X1QiH00zuQUDwa+d8nUakojXAFVDk3w0SuZ9aOqyFqL
nAI//5fe6dgZeRTYn2aTQrjcQ7ONcYqqeHabAhqWonsZd/E/tukQjjTQ4n5dlDqx
TAEu1uzofvup3/PMsQKwOwNCPxxZtaA+4dptM3UQoteToAAqOeLD3PNrzrLw/r+y
MvwSTEE+u3DfMgW52qVPdclLCLIX99W6zmxRT2yR1qi5cuUxj5IgI+zME/QDte2x
kU2EVFErSX+INVawUkCgE4rj/RMhBRfI3PC8qqdc84aY42fdXLbNdY1+RxOP+Si0
VWvRyaBJF6Ogzf4lxWED/m7DoRfzmo7bTB5KQwZdTHpDmeaJaNwmyL4k33taAqVT
lkppmSRhKMqfPTG+5QSMFqKjeYUWK3E6WfdOr5rEfUEIRKsilg81aG8t/+4Sqe1H
FAD8sHU380RPN+H/eHI8AMQ9YUmPghnKNMx6nkS0cHVufTAJg5gCO7nXrq2sp26K
4P7Ac8CcXdryb8tgk+T2Y5GSd5+ukg/8uE0pPog0vXQVW49rZoMxFdZTbiQaEZui
+zSHmQSW5KMR4UlQL3JbFBVbHXZ3DaApiQd8MtZZ2gMHl/NF+rkFomLFNz4JPFfh
EMBEkNe3ATdhwzJwuhUd14huMt6cmO8N3OoKWDQL991q+nzQG2is2/kCwSWnlWXC
/gWDxxa8LWvIZBr+KdyEluKzMeZfeVCJmPiQnMmd7ga9I/KYD7LvJvaT/+bQ7cYT
NP7LVyO1oUdL5645BkXX+QwXsB7rJjN5ATv7jmzRu9azXWhltk/Ovo+M1uIIgeWP
N2Dr6SQoGL2dU7Q1jzPap/4QTyP93jW5eneDeia4ZMNfSavv2xWhb1ksrjBDMPpW
IFv0AMiowBo696OVVr4She5CZq+ZgeE/Ni3hg2ZrnNdCcdVEt7KqgDgRrap6Sp49
4q84EUpvook41Oq83DhSBmj+72lzfMgIU2qGJXZqtNIeGi9mjKnyAcQSJKNNDvAh
vAeuveApA3v9M6fN8uOrlq0yNO1KuKH7mzok7x6kaHSl1xjeHkLy5wDBK0UFWCiz
VUGmzgVV7gCMEENO6M40ILsE7OycORW+jKBpE/jI3ykKgkVDsHWI99jN16UW/mLU
7Orm5loWD1uxzMvrEksIsmh0Zjc3k3OzSe48AK7ZcWtinc1Iu7JzmPsu8eHal7Z8
p7QCuw6nnSleWnRM1FYJ707yUy7q88afYf9MsXPzHPh9FsNiQ0zq4lZpuwE8CTmj
bij81Ju7V4AxXYlPCDskvcfXE6HKIDvI6RIgEAk6mcmPLlEfgQPMRfVvaV0p5ZeQ
WyS5+XlxQ28N3OJhOFG+SoLhsHiAjGdVED16avQCWWs1klrsuq59zMMUH0hJoYY6
227cNBupX+1tR0qzOoFj8OGfRo6ki9tlxL4leAPKEqzDZQ9+RbmI0Wa3ZtnjlNok
9uf6TjiGKjC2H2bfJIQDTZSri29Jdk96W0zGQyRFyeL6EX1KGRb8oEzmFlltAKFf
QysIBZNDuqZ86/hGDbS3rh4cAFAjLFilIClcrWX3BsgD2ob/UE330NHRtq7EbtED
oM5ptMNkiER9cTefm2jk+0ZeShchI2NsotEeWAolg0WSMNxSpapl5jqdQ+PYwi/q
L02aqK3Z9IthdPBR+SLZiS/GEHK2ode7yFsvfgz8lPdK2DzLtRaxg3gwPqra/NUG
EJ2HwtxnjPZiNqGhbSsPLPcEeVOI2NWQ/RnsfJbGuD9bR/Np63gPyW9P/5Ws2rRT
OIQSyiWw3ZY1yP6MlurBJsTRFaFabFbO2wN0gO7Ts5CokGmHKIO461+Gus8mIpIh
2aezT6VSmgB6ri0ynykWkcNn+TxCtsT1L11WYXPcTk0vtbo3h8mEp1d+9/9a6bdH
EyizdZGRafdzhAPQBYlQ/uA9Y5yGPxHXCkjtDrD0RHbvDIE9DNShbafcpN3HCZBo
MdcknraOqhoD2zmEHdNrMx6yqOpJ8i5s4GbH+0QzqIC9naAE1jdSJgt1OmvLvVWn
Ku3fOjqYSB2BECWgNGdZOmAavLbQCbraJouDoQ9/0FYTUStWHIdmOjMjhGtmnFz6
1GkPjys2GOnPgCIPuo+CZgF9j1KKttkfvAsb9PL+DmN0I2ww8pEAsQjsAShexZ5J
x7LBsYdoibIwN6D/CQXqH+wVAR97/EJ/WyptLXvrqJ9XsSruviUUUdECImVGdsnn
yKyAWd1qMuwyeONvoeWrVGOHAZZB4lnx2yUpO+gyC8i8Mg0lSOQr+sIlEhc/2AZc
bOlZwmy1E30fauZk8LSZOxosKr4GmNtxLvAfquTYiAHkVW7cBungwjSI9kuowCLe
18Dmz82DRFexqPl37Krq6kNSk9RPKJS61u3DSSkl8/tzQY6hxTTNKW41ey8p2v4W
aJtz6XmK01QAwJxOIgMPlBOqa8EoPhfTNgsEXOuyxIREoB4YUqxuTDHOmpLi6qWA
DP9BghYE19LC8Pud0cgZPUMXrvJVl+MHcABLmF9pkJRwpjDpSxGvM51dAUO6vSi3
MnnRAMxwOEX3KkgJDdN9rlupfI8+4BtwlGfjO9ZekH7IQWLVf1AnuqnGeePQj8Qr
QMuFD3GFnPZEf7OWSbgJcx4jyKhb7SsrtITrFLoJkASVGn3ZosNYL2OqRA0ujA4E
GQLmO9O4pFQ53fSrLkJ6DonQH+eAmJzQjTviv/50n8Um/Kgq3N3LUJjVdeDgGMpo
Pe3W4vfERO8SYmM2lHYPv7ZqrvCU4eZF72wYqiM/bJOL7BKGj93Q2vvnj1iGctqQ
uHOEGS2a6CiT+jWU2KJr1hLkKRgWtJRdqenPr3n3o6I9/abLtbLb35YT2tqLC738
nS2xUJCPsmylt1LoGzBsiYiC/vxdRLndqeXMMj5vySZN/K4TAmV68xnA3vlaJB62
ha6ZKpFEHKptTtYQYZt9kkXHHMS07gG4roSMtmtQ8tVzeJn6e8he2JCw6JLBki6S
OC37uujiMeBhqpt6zWotS5KmMuecyl3hRV32faFzBTYj7p+AmL1xnuR1jrOEW6AG
jyFF5zJyShSeUVw3qGXKmG8I8tH5qkNvIVWUKlKd/4xWQOaDziW73pxWLKN+91/G
c4wQ9SMyuPjaCR5MMEZNoe55evINNfv5qW+a9fnfAzvx9Cn8mbLH7tAR4YH33LWA
9bgYUxhim8A/eksZObjyJb5sgZP3AhaKsw54zY2mkKf+bS2GNVjeS7HdCRf8Ak/T
nPB3K5nZLFnDL0wzw/alSQ3Pi0qgliZEQjV2Q54sPMgyHVDvJBhekpcazcafRjcc
KApCyDJfJ4SFGv3V4ARODsjVDrzpcaJN3rE2ZFnqN7/OT5G4uB7gwa9GeDi+0v2L
hNlGuTEbqwUTzWtmhon2BpalALHePDb90t0P7RRG0ID9YbXXX6zdaGIgwpkspGta
lYgDFkq0/zeHAFedjPL4OeWvn4JvmBUs7t1PTIru9upXud7UYh2PzLZezjgw9sJT
dQtNrDY4n0Z9uzT9HogZinqh2ckt+Q/Ku96H5DaY4BN29YqIX8klC1pVNcRJaRmW
VO0MAzxaDlRf61jS1MIsomvyHul6va3EGuB0BO1ovw/AH9yZdqyuHH8TBFv3e35b
x37i4X3lFugIw8D/fpAVuWGHDgtns/Nexq9dl6qKhbh2dSQtgZ93z2FtaaVJggNr
28IwN0+QN4fIqyLc/JHSVaoqmfebsy2nK6kqVvNMeErULGbPG6RwytQ0Ll6mvoHh
yBn8+1IRrqlI5QFMSdkJnMiSlO/c9XZ7KH+KtCqOc/vWVdMbzuU+6acGaGxEoqAI
3/KGGz7idYBCSeMsqtL3x8CjJwpR4CvI4mJKB0AOP9dhkNR8uxofS59VMeFdR0sK
n8RNIisnQnERwAM3pTcCqknNrUQz6cxTlMeu0E0msLaxWxW3nxnWGD5w4ZKZ4kx4
gkRMq/CWKWB+jHlaUnphj0/2fanz5v9BlUtdmPk10NtiKAqutJgrl9Uz5EWlo2+O
WN0ZpK/D+9bEqqPjPdK5cVXFq5lwn1skOwWWxb/ElWjDqtIGSkeplxeKDwQdd6xp
lLiDbM9q73/D55eY2fIVW+5UcDTidEmm8GEKw17SCkdTUGbkItay3yhXj5M8RyG5
y3ham06EMyAgOmVDnqgCvudJeqKrN0FEQF9xrng2w7bw1bKw1fZ970rgw6uzwmmU
vu5D/pNaXhKHtU9/0OERUkAXrLrJRQZKztsdtMcRdKYCrUsMf33mBWZIIb5dDZ4U
UsL2PVlpQdMFnIVnVCwxe4gUdV4PHvDha3ejYgzM2JOX9dNHPdzusPaPglYwQ+fZ
3Lqt/69fICS77GAUU4nULgLxT4WTRw/gVvrejjQS64ozogihoGihfXMtUUeIqk8X
8Dk2n2yrXPiWNSlQAwvCOYf/5DGRahsDC17WJqWovRtmeRSuSPjPqZJW8vu79PqU
3SuG7SIXfTmsBtK9EmMfIM8O9jQj0NPZTg9QJPR3v4u9L19mPn93NGud0bXArxIU
s+XkDDYvxQAZP7ti/Qt9An8iJSTNu1Sn+xyjczJC54rioh0/709kkFkowRPj3IPk
bGZKswQPbQAYyz43cilAgY5q3JiGOnThjU0QdTl5xVghanXUolRXCo8z+JPWgrFp
OgDDHU3pnTq7Osrjy680xzCFdDEinUD/b/W8QlpPgFqGkyUen5ynSvSAyKZbBEew
Aj5UDsdH+3uxvjLuotc1wuXiDNqCj185KQ9Mq5INIKF6oLuj2lJiFsA520reNa0/
uAvu9u0xUzRzd/lO+nPvb0MSyazp3Kdi3q658apfvevJtLZWoFaJ0cl3puCp5PEz
Rs/FU0bJ+q1YdKdnWGLf0elMLGGEuafe10+vJgLQ6A/5UV7bQKLBjaUhQJJh3qby
WcogYFbUm+zmcDulNrof8U3ukvUc4lVEvy1Ya/yZSe5xeHFMzwnT2iUiuzOwsiGR
bLHVHpYoOQcMPBHY2FAgl3LfkboQQvxTkIsqiNCwXfWVAr8UoNenWWh2DI4+MeYE
+k+OjkOyJzjYKlAtRC/ceFKs9XIbYGA1RWiE75zEWoym7cOfYKAM2E2zEUnmZkCK
a92QxcugFJMJwyRa2LehpcPVHwNc832d5oq3IfRFEW1med35kEfJ0r8gxA1Vwt1A
KXrM2tdWQ4LOCRMRheteDypiAfEXxFbBaTs0jpp4jkn1QPsnk/lzH4xj3aJEcE+Z
OZ91CY2xiXxVJ4IqpqVpiHlWWmHNnujXnS6FFAqEJOjKihyAYQR97GI8zoG8mHqy
ZAtdd0Hj86Q0r2FR6/BD3UKtIOGlWnm+Gzv/ak7tXxBSJ042UPqZ8PDuGNqm9QXt
K2NP8NSp/vZS85EOH7qliaEVIdJoEpPRlbjTCaVxxnQcBnEEnot9lgmepFMQSykT
uySGTnH6fyVYNNdA9wewpt1lDakTtoZ73oL4DGu4CUgxRdZjYs4NgrFGBNLkdg/2
nc98FqicPBVGIWcfqmehEkVV7VOmFX1l4QF9n/j6xvJ5jZQMDef7/K63jKUxRPD0
6rCvb0xlZYp7ZkQmBMErJOEUAHRNRUzvSlEkdWhGysLmYuLDruvGz6XPE2HScmRi
0pTiEclA4u77cF0wPd72vOxleQY88qW7SqAEYPDmuW5eNoD32hWETuAofsCiZ9M+
87RgSzzAEm23h7EGeqIdWNNywJlsI/QBFLBxR3cQWNZO/fUUtL0yK3M2msgDw/Uq
mrYhDnOV5m1XJSl6Iaesxul/A66y4Mj/YbSPm/RjKMjQNjdyVDK39xvW/oOIoiUu
1FIR1Yf4wHI8xPJesXuCxYjUofZkwDiyfSh8Ape9bp+kvsCu/h54oEC+1lQxWN7V
7Yr0Q0eDWXt4hl4FPhkpOoyuqoGk9PHXkW0z7naE4EhUk7TqT4UDDXctMqVTMYHz
T/+dSRV4PcvwLz2pD4NZEQHzndEsCxe8+oWhtmqkgBrkR1EaP6ejYj+IojII/+P+
+oJMyzxXH2PnCG/bk8K6k1Z8YnfP6A20PZTIZrAKTW95M/YQeTnNMGtTFZpjLbUL
fEvWi0g6UGnI7CYwyXIKv3C4mfhzGNh8Va8HlvocTdaef7t72TzL3Lx1hubmtAAf
Ujfu5by3EOVeV2svoznWtAOblXkkxLHwql/M8XYNp6hswej/pAsfTYAw9iG2qSTR
PSzofEUI4hD16/sevaowTSpnT40sq2981CmjdvGSmAWmJE1R0UjtnbNDzEyPe/lj
4d5G8qeS/C4CDQiCrTaNv9CkJYBgfu5l5epqPmqCRTrUFo03wZViibTW60+iOrUb
hfOZhB8mmHCmMSk4W7ZD5u7bvyQRwB5C0sol/hOlb7Fsv8FltSdg8HlUIU68MyHE
BlkcXVdnuGpcV8hikYdBq4gT9Pj93FP/tk4COeiFUYENBByiuuSYsfoe0A2Z0z9Z
xzWkSuGctsW4T6G8gqFxdIhywxxVX2e0PglFfo3PyS1jv39kXVS4PakkTvtk6UqF
DRmdbsGjpeRnSUPAAHePGlMxmJ0dhqFaRar1StlNqAW4g+TzuowrdEDfsCA5KzNj
Pa5OGQ0ivb5M43pzpQwAQ1vN2d0Rk0F8KqfIBqJPhqUi/wCkO0INjjeL/IOkusv/
AORkpGM86N7jyfKT0Jsi4D1g4u/KYT5Y8fEXM/55TJZ7BUtuA4pW1pVhJWA1a/4E
aH47IHGGCp0Rg9ni3AjC2hq+Z0RF677aNaMjHsHIm3+DDV0nSSrtmNYLX44tx+ln
LgHK4nYeLXDA8GtCzyGq9vvkEFuUgWitvHPawyRYgHhkrKl48ITP7D5KFc89x9E/
DRkeeBis5d0uIsIIzjS2dODAKyK8YccSGPYXU4aX/a8FAKrTYw5U/A3EHHy4RWHe
bPP00/DkfLVS+D8CDnRLJJ/iy6/4CuNBSY1n9N+EyPPAzGoPjRFtEdXod54q5zfE
v2Q45pBp+vT+K/bl/Ws5v1CXiuNerk6psVXK1qcVIYIUxrt7srQVNHwx+OgheY6P
NdLtSzX6w7e9StIVhJaMHkV20bSYVn1Yi1sw6dPHBFHyQi1Hd4iIhx8fljcsAux9
ZMSPV840QeQDkhIf5uJJ7WUYyN2OlcBmnHxMbELWXk/+tSnpRBg3vxocf6SpdR6F
V1XGK2/KddsBRbi1IWRJysGkRUsQZ4Z0jhIwu6QsGUR/izbZywzU7jzPL/NFPamz
SuMeTF9ThRhH/vuCjvYsqCZO3OXvh0x7QOXfZb/h7qignEh1xGBAymmbU0j+iOtE
8wWFuez8YO7EuSEFhjHcygvNHsW4Ngh2mhrlCtbeobWXEUetLHZNyBKGCP2fuUgw
N8f5DRjxvV+SPSIBnoRwfQuR4x/eBewjbsidqLY8D/Gu8QvoZl4gJ6QspwF1dwxs
OJsG+/LdrYx5BtWn0S4nWRzjs3aUu1bljjV/o6Sxe2bgE6tCMGl0YVamDCR2jxfQ
ojeFPvK4y85c4WdgzjFEVQUTImJGXDD+gUvc0lgtQ9JmQFTNOgdHRxJ9Gd73CCc1
HOCwP+8s3iTNVnTPjyG5Vs9ukfP0nGutHJtchDQNkUrp4dB2DopHlKaUtxmWx+uL
PVYEOmE7afJjOpcrYODVooFYBTiA0zWJqXZGkWEGKdMt5jopa0LceBVVmXmgsc+t
8XdNR6QuKzdMJTOQbX8dk4W4KrSk+JYibwuKjXxGORiGOhquVY6780vOMQo1QnyG
My1IFYwidQU5rKk28R4vfIg6InUwfKLKkwH+EtBRpBrNBssJpZ8fQE2LLU7N20YB
eFNCbXyw1IM5epEZaAHeLdj7UJ7R5ZWnqp2ni0pDJ+8lfowya/1qOn2z8K6Xh3FW
xQygNSO3SaB/p3LQ8ur40O2gN2PK4+xO7zIgLold9HW3BnAVlY1n1mW+L+ZH8tDy
etT6OHzNaUx4Qs0eI2/O7ttQ1nDKU31Pc32AmKD0jm95fY7U0MgDqYykGEuZhSg3
8vzcZusFmJ/Ub9ICZSxYMzu4hHghSWqSbJgpO8dbi6km1vjjkRkHqscWUBAqcMvX
2K9/R82nqi71B3MhO95PLhfe88g5yf2bm7J0IIUl4onO2soxtdqhFH6BupNrjRfP
3T8y/MHfmUGl4eMxu+M9yAgqtGw3UanUGjL3PWblTyVgMqFEfWtkkMhjLtGicYqg
OiM2VXnGtNtLAP5qk35uPFspRPOUOrateBdMo3IeirUEqTKXlcz4vH/a6HCL0s/G
yUaqoY2Ul9ILHmT+KQF1tsiC5+FohxxQrceQHMf8ARjyJMQOaPVw8BSjbL4VK9lr
7LhTluCnUel3egcFFIko7kSXGDeULSyfZUJAA+BDWlqdZZ8zht9gos+HpixDhoxW
8IzhYim/JZw/LODpUv7D3x5tujXlgGcOeWOvUy6kJr8w5nrBKjueSjd0NJqU/qP5
eJMECT2spU99pmCM2TDhZAIO8SxB6hmAhw4iDFpgS0gGeXW0RY7+EnrKcPXJqRYu
tdCvVnlywxLjALH/xJ17FT8+H1GrSruObuht0QP9iyZRvW9jUZ8D36RLo9ub5dfs
nq9+dbgWU7WFLlZNTR2EquKqOAa28W5ehS2X1yy7hA8QeqZLHsSWIi9fJZFgT+34
SCKVV3Rn9k1BZTAaoXB96+j65IrJLJF875Zl4Yve2/clIZkhQsgOL7km7e/mccx8
Gm6OKR6puMN8kEfDq6EPDk0RbdEbrPntBgris90HDd6RGkgfIBwO2HMFE5GQWT1/
wGAhhrzzVHxgGHDJMV2FtMLV22WBotnYeHLuCRe/B4VxTunHcV71btstR9bzP1S4
P3Qvco2Zk8dfeEsc0HT9P4vdfDoXoI0lwqWSZfqE4HRjEunfeR9NMtCaOeJGoaCW
h0hdiD2hDP29nSeorr1QbSu7By1L33edEGhL2IP/NHBjWyUU7krgmOvCQPslx6Cs
4Mv3vHedsQmwlYR77dApMwFqft3zXA/v+wFCh/TSY4oHdi3wQqv8/qbmiUFcWXej
8ATHUsFko40mF20GxrjJrm8FiQa79Sn35om0OVkRRE56JqIVRyR9+ekfbK5UZqQW
2Hc2SCcQpDaKdyRZm5lpm5Q1zjiAWk5xV0yPVYVhbOvRUz/c67voffHMSUwiHIzW
ewMGr+BYdhj36V4fvwXjULbVOci+dS9ru6MYUM/ET6MyeyEvalqJWTS1hOp+E++n
TXZE9iZ7SovVeLMCE+uLw/oUu5zhsqkERKZzIgbMEsUi2sTRT6axgO7LUVse9JmH
JsqbJOPBV+/BQ4lGwerbG/CFv0auU4ScYnHomJBPxDZYUxwfcaP0elgHBVgn+Z22
BvMbcKa/uJMejpHW7pknk/JjN7azVK+ehhSEF62eoZ00i5sAFMUyBeGEWpG9Kwho
ZveD0Y29olzC9DCAU8Ijpzd1j5iC1xPsefoMrGGHjMgkQjKlV1aZzAtiFoEQSs3H
/lvo4BAgDZp9CJoSNTNRmOgIyjZrqGYy8HTyBT6XsZPAcbV6VPh9BQ1idutp9sor
+Tw2QzsbsXBEGug7l+A3n8xgS2dQYsdsU7YgpVjWPp05yjbfO6QLbtWDavlLcv+/
C4xzKXm35a4gyZhQiBPmExg/XyXBZ6tnPzH61rDw/ZSVcvAHlgMTX4cBOaP6Gxa5
tynzOIWWc3ELc9hYMvkBXEFJtRBgOE/iGFYLbNERomzvR8VHr91e0v7JabqOg+Lj
JKJtcdhb9jkquwu3jhpboqAJPOEvqtz1Fif/BOhVkjijH9XntElC1QCtHwdFAq2r
YrN1e1qTFsZDXhbnNNjwxaqOwQ667PHSOflD3AWvAKIn8Ue44zDx+1phRvQ4qAFZ
yUkmDgcF1OEq5R9RIGYj74rNnhRXLGMAy+Zt1aGj8Q57mqKJpXUNNXirB6DurfA4
iaiQ9uvafADOGEdxRA1Ewr4PbeOoksL+eV1bsbPKuPSmwDuOqjZ8PLT2gBbvuPHm
q8G2L9AZliFLEq2sdrfIME7Y3u1KvdWIOP6H71tJPAS7I0FMmECYPY84wffHVXZF
gitsF7IybZDjyTpG7ZaaKBg5dR9xOpVtWHF0JW9qmDzFEbnBAa+ytR4eL3CitfGh
Tezr0ZkhrxUsww5e8Mfj5rOUr5KHGtRFrRqUi56fHXYVyHZqG5duoTL+AvrxNw+F
y2/W/+i8Z8yY4dg4IpefxxgWyleMsJ0Bo2Y8hJROIN6h1/7e0SW6iNKQFazmT6o7
QF6LBFWMyFo/pt30vW086+LMXO0VmfTSMC14rG0VIqYXXylfWkGj6oBplJ1xcZud
3wko3HsRPTooL2kx3aTWjlFSooqCjvsyBA/Ob4Z/CceE4zzlj3mW0eETQz4+C8ov
xkIJVwG7SdoXgeZTF06l334IFsGKqvW2xAM+PuoEfoDIA2YLRkRdjPPPdX5hURss
9pbsu1vSV6Xh4/mJCDhE10xXKJKS4T1Gej/SFuNxo0uWx7LWJ+X7ra3+mW6YCaPq
oUPw6EEm/9u6jO5vQWuuXus5KqdWRxeJsYyMkJZPm+M6h78+upObjmiaH7smvvPG
eWei6xYnek5r/wPe9b6UMw4U+LuSRQHvqB9Ruo1zGRa5uLQeuunpK7cdWfNBy8o+
Wi7ULyarYcu/tazLhmve70IPSMSGnqOUa6QbfvGD782rKzGsbuidueCZZhlMdx2G
cryGOxFbd37PrpP5X6o0CxEPuqrfhnehQ+TKp5tEztFNEMEd2w25v66uglugnuJD
OYCUaYYWctTTgHyywVAcbfAyzJWfxvxHujUqYdEbvAzCEHpGCTujquweABTa90d1
/AGQX70wL54f8PUOJRDdH2Ntdq68Nxz1nB8Eof5Bjrl9H4K3/AY64Ol2HJOSHUZF
h2e0yuc7kTKY9nnWbGvuGkTEMA48DmlJrjMVtxJXcpmcbdXawDy6GWvGAZoDt+zk
Strjgkm4IBtztRBDzd0ecOMR4W5vzsYE3tfP6xwBWSKRFufNGFPkR8e+/pnn1Jmf
aDJ4jt5I4w5gjdjLPB3tVpURVCIdyUEOWZLXchQI5nrBvjdvZveE2DvEP4rgH0+4
V4+AXLu6L6F+P3ERnhdwpnVfKkt9rpnegrhyBjx2n4o1JJZTD98uPu1Usn87kDyz
ANg9YUtuo6BHiZWsNxXOuvENKSnh7koNrGGMDXQ+3okt4m6AH0oBU0qvHzS/pIQy
mxTRFxq4ZdY8cn+hOSQOXmB7RpMlK4UtuJAITshdpJmQwGDnY3jLwBK9A5Oy3wkR
8DToiUxh23m3ofV8rnhKRf7DPfFo4JHhWmn0U30cTeyIxnU9lAHKHCVBLI6pwqVb
vplMHjR1atZnfsktACmSNCRG8Fmqh5M2NoDzgj1+raJyoKezNLh1YwX6KXSP8Ctz
au3+LPooAPpYAEb7HiPPlzkSzAfJMFejDATMts9TOJkC58vj66DiU/GcJOOl+YS6
WMC8z8SpampnXrRmZZIB21B5raoA8oqVxrRSsbLPiw7iA4wid2Y94z1PfgDYt48Z
fZDlHXOSUCm1P3R9qiP592pGyQI32iE8Vr5ZMmJMT+HVukrghgUy8Oqt/g1Opsyp
jkD4WxI+P+PqgKdP6d0qqllJ3lc1sK9IngnB5BL6trJep2d5ZjnzuCtHbxZZoUQm
IWNWWpLLakNX2oZtzeWFhyV8V7hLB841+EbQh0JSSh+rbJQaV2h/IRG79rntEAcZ
eduZxBSjfDaqzx+pFotsHHTrmPS8xWcV07YT+43Wb6qem/6fwaerNETR4oNFN5qw
L3uDdVlH7weRUVBNelyk0z1U4nOPUxIXTsQB3kW99tjb0uO5YjRvjOiblh80d3eW
Jk4bxGJHjlFQi1WBNQCH40lPy3SoKCd/bIIYH6fhhbSFn4wYcnHQWW8VolNK5ILS
smvS/V5VZJiKUY41pbOubQSxAoyffQ+Y8wWb1m3HjIfBn+9/Y5GWnTLLKdNevFv2
gx/TIkf1cMXWf6JGLo5mTg1n1sYNdjz8C64XohfD2iML29bA34qN5T4eTA2yE0Ms
S9mKQZHZ4Of1FV/6hwRbsnESp20hD60B+NRzy7p+TDFJA9zx7mY/TUZMnELMWWl5
nIqc+l5lLyp530LIt1G+m6SMqE9ECJlgTGQAlSUa2/UChqKm2XHpWHE64rIZMvCJ
iYuKVwNWivj43Uuxu5/Eo9yPzv+Pm/KPta5594fvkStLOLsCjvhFuk4FhpvIspqr
PTcXTq5HscjSi6di7vg7/0LFo466P81FNBEGJRTI8LNX6uXss6qZ2DUGOHP0JuMN
p0RJRMCSbCqbdeFVH497vEAaeCcj0HnigDSWsojrfQZ9laqWblDEh1OkBlE8A0nC
4daw/NRidUvQ0WQfVjVB+vRwxw7uN1Nz8J+HfMzOlwoHujyN4x76i/Yg1WmPSOj2
tVpkDQr/5dFT7uugN1ljS7dWSz1GvLbpQl96aF29WXUeYyHSbZ65Crricgbf41TD
+1y7JMM20oY8+bg6AA1WSWxk4wS1EjoNAYKyaMUu4tbzqvQH0THSyvNeYcAmIs5v
3Gjmyj+QqRwk00zdBisFatV/OjyziVj86Q3n0t6+8s7jDtdTeryRIRRw+vODopsC
kYw8FzWs55GRWWQXNl7KhGEtqnlvLcASq8o6/Uv1PryDxnKZMjedtgKGQzwSMOSF
yMkXnA7BhUfygGl3Kmyemz6Gy7l/bNTJ7ztBjnNnfip9cGKyL3DBfEqaZBE8pWLk
9M7oIiJFsYleW0HG0a6vGtBs1sOTz34LcV4229hG6YEmAtRRCBL+USEDFPT2hE4h
Ejpa6I1nHqhIvzpwK46+3CJe+vCHJgOdZBOBlN6aZbTEp0UO+HE3kspxJVLpm5CA
csTbO2WYuT3MKm7SebAWWJPttCKqwcgyMeio+WYUBqsSC+PDn9VNqU2J3m5NkUAZ
G7qPNuqv/lGq4lDjyGmPhwpcbCczH6ozRjZvyj/2rHEjcRS0K9YIOsXOb/hMlnma
azwlOsraRyTHvqL5Uv5YUGeIh4zhaXFyJlBCaO7ODrj5pNuxmpjmem5Eoovy2RaY
4AM7eA+SEXLW181ue21b++AXdAk9blEPg5qxfIqHL5skW0YTL33k1uCqCSIrN9vL
qI5NdauH3BEVQ8M4dmYIwoEKbPVVUy4gK2XtCIJNops2+/F6rBYghwjDNy+6M+nX
KwVnESZHqqC8EeVOLj3HAOOk31gncYyscdcO+uGaNn6kSr7ZWH8rjcfIs0iW+mq1
YWdtn+uc4E+x99BlDJljT19oDVWUhSd9GJx5+NF35W7NXH62xdLPw1Pi+1hMZfoN
zzYZkoIdoYFwFxkcBtrez5iA+oYZHbl4L4ICEv5HeaTUWfAdbdQD2exsAxFf5+Zy
325TKcF9VKaWXAmXULz2HQ+u8EKALzEEgZdmX5eUBHZev3tiZKRyeQXKY3SU5ls+
XkUVsV02fx56KUfKEa6Vxr537q9wP3y1sdmoVAa5xpuuic1KyFj7nNiHKijujz3J
x5q4iVPTQy4/2GlPq5EISBJhgSAJMJlEea5lEZplvFioAi6m8v1SRYcYNZi9BwJf
Dr7vE9Sv0IsipqDgx1zbSJxv8UdgLkwYDN8euipLKYerWGOn1775gyI15dauqpjQ
zoNeR0fTTOm4WNVm9t16WOYeNqkM4tjlf5tStw8fmeAFT6fzEFJUv7NnU6SZd1Cs
GhmfnIz7LrOAyt00ErKrP5tsPKiGdUsuveynVrf4aBVNtB0u8ix57Ca5u/4xIN/e
X1yHmkx+YB+Im/eZZR1WJPKIWA7JKuiq1M/eQ1hqUvdEcsioYJ/xPcD6nsnpymft
eFqATcfdHteJr+JP7GKcFNblNZ06I/fdgBnFRmkJp4IrQfGGQtMPIEFjIqNYYcRP
7kikLefecLDcoKYRz7p7APeu9FHqLeLCrc6fs3gknv61bSLC6AewZyy5sysKMBOy
5l6Cer860e/ZDSQIpu19W++I/CfU68CYKW3B2aolieR5tjBbU83SKYm1cVznMzWs
NBO8JQeRhR5rerXL41Z1YMuHHjA1O37eP1cHYZXzLOq1Lt2SSS5MYHzb0HubSOIX
+v0lG0F7KynoNWU1tsKaKMdqw/hyt67tnPJfvccT5Xw6GpPpUeNbK9EXOF4d0mTU
RDWRrQH8hGpNbG0HSImDtcOKcbl0+Yj5qRElFnOR7zCs4/nj26OAQIHro1phNT7u
mBbaQTCrVDrv9iH1g3kcYUHqiTpAOWZ3tus5fFw8hLESlOgvApMbXAwbQFKYipiu
j9i8yIYvYTuAYGa4qcViXG/rOMj5pNKVXzTr6zScZamP9d40xWS9JcYJRp+OFCsN
13N4bGrlLSN9n2BzsveQbBu3xoDAYxqHXL8zu+j/8ObjFncHHnWAoluu9cQLzRIJ
snjFg0efLDG4gwy97dnk0uUJ3feifWDv8bQRHHuLWzCJjQpR9yp9MgCH/IfQLQUN
GCmEX4v7H167/nAXzFUfLuqrUHy/gAPClA0Ai8qm+CEhRU+/P6sO6MKFJZXip7p1
RJtqzIi7fnxNWz+UgT0Ep5GA3QVXV9u9GbB3vX3s/o6v3jsi99Lo93kB9vhLH46T
LMeKJHOM8U8s5qLBrHifFPP1VcjNPLIatQ7D6bWK3gNmSMdC1HxPGx1U+Aqayptn
E2QLLlwIhm2C8xbLsQ25qSocy4M6F2sskAJkkW4MIVeno5ue3hLxUv7xb2vsEiCS
6I3SESCuKCQb0nIDaskEhgbXEi+u8tkov5DSFCn2k0k3mux0c24CCsi4xghNTdhN
Sn8dVoRGdDpf8HoO7zJetiKJNIdF1kxrCj4DdwN+yKyDKFl6h5ye4Lf4JuVX9ZJa
MLUbRAZ6ZRpbVfoSF2h5n0SlwVi0/S88bJS8I7JHSVZPA8lywpOD/0cTLAO1DFU3
uudvc8t4K3m6i9Gm5vHDl1QCfQjnVNEDdrjRvlIJg+yYpoOp4xUxxscJ203L0dcn
nWgssC/FgHUcWARoH12vmz6hC2S9HIK7xdK2I528Yqg8D7Ynxj8mhlgTlM4/TBIQ
sXa9lnY/ClnWTirSMhYH6m5zQVx2Owfz8BkxUCm8Fqog/csfXyGnrdVJ47X4xb8B
H6sLX9IYD2UroKK/kf6fveRiRs+vVuQXsCLAP4V5+oYCsbXG6QxeVfeW4z1y6Pky
Gfz1AXATeV5izHOYjkBMi733JX7eWAjLsHyejrQQcWwbC5zT1ucHrCglhQSeIMTL
V+W+BvDmLMzvHGBTYPUdBf6DkrHdERZLQ/JYauGo6CpRPLAV59GCAhNTTDUuCyuF
elLzdXvtCO6xVQ9Zd4NckWXe3V/4ZOU26f3k/J8g2M04ZDKemLVe2wkV5WRiS6LT
07c5VnzcZ6MxiMSwqd/UimqFx5TExLNSVGe/9k78LZsP2661P5G38YEWBLJgjXaX
8juvI4e0FLF5UHnGxWCRmVqDKwIulU9xC2XuML30HfBhJLGs1LQgXchzzOExoQ8U
jm2yJC0g9jXwYg67G2MFRte7+mi8e5ALYZpmcey5geFzIkKf1v/mHdIlEWUCSva0
f8t8DT5y6/emC5WGdE8g2zrRrmfNFA4xaZ6nPie7XqbB6dJHM2JcrLNjIZoxZwyF
Aa8yuKE7O6j3qLulEn4/JKc2LcwYZ+kIJ1ia+NYiqnNFyYc5vBNs7baWUtS6iGhy
jhgAmdAOuXFrV66ELIgL5ChH6pcuvZO5EgfEK30Q26d5QbhJHtjK9tkCL0d0AYXp
6xkh9BD4dSVpNvdPydv7C/PoI1a02n/Q8KTrdvY0F7Ex1QJCh0YOcj+QE7/m+6Wp
wcVZ1K6IvIpCShwxUDJUzRM7hLEm3KBK6c4McLuePt7Jw8mUHBOrkExj8UrsYK9m
S35q56MZopz5+VBezQKb92zDeHZN4wYbom6e8ZruLO6CBx4SAE3enKCqyJ1JTiAd
Zche8Jf8vwhQeYvHuCE57iCehApc/UiFLHo0A+y4EKel7eGiiMcawAeYcL873roq
92SQQWFGG4OwMdaWdYHJ6C5AqAiqC+7Os7zrqJyDm9Z53LV8txvm9NQtggEnSmpE
lWSM/CV7YdT7xj7nx4QFZOwicYLdVeYcW7EkrSFVrpaaYxzuqp2/uDdl2MkVg06a
kCE+tnE3AW7A0zmRlTUW8XEjRd/ZbPA1lbaYi2bm1sDqu06z3OMDI+Fn6jkI6Lbu
c6gF96RtAHLgQVmeyu/lug1W/wAEMc/fTVJ5mf5AokqSMRSOat2zBYrY7R/474Nv
zlFrjehU3jGXQ8snnl6PATkENkAl1CAdlbcq0ILf0vcZEMWO6DPFymjhUO9W6sBV
AEw0R+ocTvzhkCXZ5RBh7f+e53omitYkh0ZdmDjSSn9E0v3ahr0AucjfbJaA68xH
YgOiLGnr6Z2kci55V2kBavystBWLNMqZ3+aBwIvWRvCprmplzq7hwpAIoCY6SEjH
td7gciNWCMTIEx6lVsWoxaIaAGyJ255L6NQWVfBIHQd/PduwpXgwUX99EVh7kDv0
ScUH1Oluz6b2riawtxzdAou2RjcYJLqbGA3UQvi344K3VzWRiRVtteWWSZq7x5C0
u963iAKAffEyge9pz2o+9ny8rlmuQ8k/yYbc8N6AmXBUcwWnyitmTgYfFutdfM6t
NRpB/kiMJ2xeUUBrfMPaxPMzz0RY2Hci6v2A1x5MmDp/MfLwTNT9mK8yW23O2st/
4sJiMwpGoum1AmS4km3lSFnGqGjJZr7dShAAGdyVDe93awDR2KbzbJnIB6fRdSjv
D1b2sxCQ0+Db+Bd80/QAP69+y0Im0c7pNyp1k6UKqxdvl/LaIdVkBB0jaAKA1oW6
lCUzrWplVM3KtlDzJsqimKmsaiiGOktBGpnNgSE6Q+LGjCNFC71dDFswCikaU3vM
TFdaRizuwwvh7TQHyN34fWDi7Nr+s3tkTKuQkiu31fAQZKoZNTFNwoApk+9sgEbm
hhxN9zNfHSCqeYcoGwW1KRc8e64PouiD04uC0+l19H5wzewOUdm2H+MU9J+noRah
DgONmm8hx25IMhWE05qEtwpWk2RnGth0a+Ijtjzm/hXPWzNmOX3IFvfGOYOo2Ycv
a3uVYaN/2WHkYAby1H6VTQPnvDw0xm+RgXwRnYuPhy3r83AQyFzqyrI8t6xYXVO6
ylVh30Bz2hzYzyXVlqDHrLSmas1IkdUdaVLOsGD0ZOgCanFKFKtuHFqtw+3g16GQ
yjkP3CuuAP82tUQsaFWMexml71i9My4fpzSYNm3mWxziObMKySTo5p7QX8XLdz1y
J1oBkz3+Knl/+aJOhXPinjxswreG6DgsZoyqDiC1i0ClrZX0XUtTMXbR07yxGE4h
UxYBjX/4+uASiRfhz/XVzl7rF9zKO/SX5HhFG3LwipuK1zLY/xjU3bPNJ7ChmeYp
JUy561gCn8YFo/5xZFNPQ47DcRdchN2ShAt0sFlUHBabawJvbZDqsX6mRdrV9gTs
7V3o4Z31YW4a1Fr+FkFLT2urF/EG21i8XQZGDRXQSbxv4Jx2Tgo0dgHoa0Kinwky
ZbI2sgPDkpfPolOf30NWbzgoR+CmG5UTBms2eK9UaQ1tapn2ERS/5Tl0bC2J5xJ1
eewebEz+OMbzuDyIltu8nwclw2ZyLDiIRrVWPQWTx1E+MhgVlnzErVUAbPR96Plg
0GVEnnuivvnzlfWQfZF8dmr0kWPa08Wq6BEBVRVaAdzJeN5V9thOyRO3wcLi4kFe
sItcwNadLRGSjXoFqSNK01DSVEiwSB5Mh+azvAJq1I2pQCkkW2xUNeFmMgRF4Yk3
BcbtYzhlGluAoBuBUSnh/KGGZHBmuboPA27H04V0MvH9G/NhCV84ArRKNug9P5nF
6KyL6XvhATn0j6Zzt2UNl66OaMtYl2FiotD+5koELDSBI9fB7ENQjuPJXpXqlS6w
BJJ0D9xQDJQpM8mA/hpt313nYKl5Rha136KuNa2tV91Ky0bymB66iagceY9H7j88
JHVfowOyPbDfo/Nkti1NSc175QDFPIi1YfgXcdXSJWxP1RR+n7AAMBzBNXY2REje
hbiCAPXns8Ls2CRqGMlWcgmiiOmqKeJ6wNqqvVawnnlQYGHPlnpDBiy42u95L4sa
D3aq4Fjs7dy/sIt4pGW3emO2tlZ6sGbgmEFYeRM25HcicxyqNDsuomDsvnBeSs5W
CCx/jfpfigEuKR8E0PCP1nROfe1pEdpocbGPYfqhn/zgnUlUA2sD9DKBFX9SHZrd
J2LqwfWL2z9+4AVtbLElyjhwbmn5fu20Bnyk4DlbweQne2Nd822BTKxlr+FcCaLE
pqHDSs+fzFKG/8tUfugyqk8UOpr/wjGPZTuPhojKeJ0SJx7OIsDpZ1ExRUS1ESXG
E6jnR1TCOZ1GZfmDXno9+qAfT38mPuzBwNLYYgQd2BMRvKJvDB2J5PSVnyb2AM8j
udWxXLlIs0NUnEAPEiZoEJdj38hYtc3TsJmeOSbZZrOWV+dOf0dYWSRT7iNcZe6S
iQjHkcDwFxZiuDNOwtpiA5cuPfYMrho4+NKqpCeY9Y938nu9z3aeHw6c7vZj5JeN
lT5TSDuXCwtNAHOpGIT6AMn3pSEWo1G3OAdz+yzy1ybrE5bhRUBfGwDl6nAFvFXB
LzCkjqKS0NjAwdDUrxkZcLKz7Jm6HOpfSyU/2kwCaYrq17UqiaY425sZOJk0SBO6
VnMZECHbidb4wkw4ACL56pK1SWDHjWVqEQYmFklMvZ1xDoksPbdE7S2V5x/j+00I
dk+Z6Gktb8HAHHFUJsEWDmpHlz2RFf0bVZTKQbQEcSf+A+5FYcdCvtu38YpoWO09
uOZzBnzxolkAFVkW5Ph4Omzo1Mx9DvkbHqOGa0WhS4YvWUjJAcxt0wUlJAXtHrHi
qDf+rqMUaoGnIEqqxiDYL9K9L2aLD30WBeEV00RZXKY9dSDw7qNGD0cwT4EBm0eT
GxBQJ+Q/InwoSvqWnb4rMjTluKebX7Ovxbos5x95IfyvA7WC16EPFAAMhXN3ebJy
Qut9EfT/al973wi6ClfsrJgnm4U70TbDxwBSG4FJcfEUviSi9OBS9E597GVoDS4V
U5yguSsx3sNlCytbe5QGiJMi5bhxOPj1+UMFPDd1LWbpanRtHSVt4GGu/C1KFXfp
M4FGfPUQAmYekiwm1ahzpk71A1sMRsv8KwKUTyMH1Bh/PfPcsCjquzjgCmwCbVqQ
TJBu/xQTb7EFsxvjBdo/1ucNZxh44sBVRv8EVnayKYaI/p0eDrA8Vrs4Rw2ywrqz
Xvl46D9vT5YArquEGCu5xo4OT0768qcQ0JVPR0G+NOKCWpBLIonridKoVca0yGzD
XB6LlOjp8o9VgT0cnhsCVRcEdhlp91/gjqRAwmzw1Ur2IxUfwGa39InjaPNTtl/t
S32eIZcEC4NsNBVR7WrpNAe0EnfN3RTCOl6IYTSAbv9XerkkcajH8edhdeO35flo
OmqUSNUrcDuYnuvsICFDsgUYzhLK1HVoarwvSw6S6A9zkuzb+QvxboP4YYcrvKYB
u+5aQGi8A0AWH2Q6/luV25gC8lRT6ia8zNFYk7paR26DDqxh4ocXPtFo03AvbgTP
Y14I3SXdqCdKDV2HcwovJ1maO2KTQzEmOX6Fmd5moDVJljAlBmFqGMogd/61OQN3
jDnxTdzbs3oHBBugmzMo9uNrJ3mkMaBnWNXQQFOgKGUZ1sPR58KXpYmv6iyztJa9
dUQKxCKk0ooDOOG2noycy0a2fqhQjGvI4fFLZjMCGA31US2AJQf50oXYbw1owtKx
HyaTJCIpLTe4hFpq5RuG0b/ixUAmpprtYWahjBde1AAMy+IkwVY0K5y9IEawYc1+
h2Xymh0K4NOT+3H5P38M5127HvK2/VQ6nG7iOGH3SBgJmO13pLscU5BsLfvbaiJn
mB3yVjMPjIaFRQuyebF27GqGbQeUKrUUbDwiuoic8ZdqR5gdTmJUtJrRksxrlMSI
oQarDmOvUdf2sZFBBQvonm6kJjaX/XhMQSto9apE1bLP0KYry74ymLkYc7P3BSzr
SHVUlaNxTo1dL0caDBJLoDtOOaiL0/IMtcGipwTYCZF8FgP/bBOafBdfGjJRIjbA
TXZzDz2NUfRaYl3zgAPQRAp/FV7wsGWD73SUqQVV+eYw5c+LZCzn+wvF7kTy4LbF
f9y0ZyYU2ItL2q6T6frAH3CwWv2ZXZ6dFgEu1vPYmNWe1q0bGiQ3d/tC9s3gu/9A
kLabih0si9NS4BDKpNcjRtknn57+2F7Z/9/fJWmXa1ukC75MZhi4NzdQu355hBGc
2oVCVWw37gXaYoj1ypTKutHaLQTM/d5rTgAf0Jb6xg2yQWi+lZ7RlSN5hw/Dn6mr
D0u/W8tr6UGi9n7OqX52/vuDaxRL4DaPxibQBzZTqwa/ga3AmJAaz25uo7i65Xnf
EwL2oOR03AntOj1gb2Y2LyNcfK8VT05X+qqn4jwTzxnUAtdM1wt/z1HGN8dPthKY
qPZl3TY0AbmcZpmPEnpo+teFbzI5XRntJR5oQ5P/px9lKOvu/f95i9NWOOEfftOl
ILevbLbRzggJfiGFPEaSSj6IWdv6KLY/gSImA+M92avUXb6GX4qlnMH8hXu6LsUB
F5A1sKOjdh5n9UjG86dPhg1X6Vn8Qx8gyEI/iui/gJYhoYWOZazXaRJgAYuvoSt4
cz2gs7cxExmYfFdufUBNGBrqi5wzOtJa2UrxJuYfnjCceS9N7kLiO9iZDbLE2xGj
TZZq1g7s1SW3W2EpC/ZoDWHmuaWYMp1ehJwmmajNinHO7ThO4uIH44vpbaWEQcVn
dQwNaHztkEoPAsCbUVt/ZVBD+NGWBRcAzvUii3rh05ePRqimdUoXtFYAg+TDjXBX
urtW7DExIYW2U6wDf2lzkUnjdit1Zw/z+kpV9ttnJNvqd94Yjf1o65ym9MJs+qoi
JGK5QQ0ObXUqzgtupLjN+uZpCVkxDHpFc4JBjrObdlXsoF+lWcEAgNf7cHPklR7y
MvNxr6OVUxthwV1o3SxxwYBjP74d3MuaRVKDAXRBq+n5Zntxu3P5Z7WOSaublrOJ
lSURzKRUw7MLJkKiphgyRMAKAr9J927o3UbkDSOdJ9SQpkbWE777zzbh36nRW3d0
Ws9U1NMY9VvfYTtGiqi2fDTD6VSWoP4vKnwKLaNfhJRo6SmqMY9B/lkk36DXcPGU
wy+B6ML8HDTSaeOK/BBDvBR2t52KSNnaEE/IDzszBlNxeLK8fKu+sjKmBtG4eRhP
zvweQJo9sWVQ+diWqDYkdIPm5yCdVvgy+rcnCE1BKu9KFg1JumNRpn9oxUaDALc8
CCGjjxbmrAompvDHu2lfECDQQZjhqC/QAcSWgRiQfLkGk+pr6vofQRWhtCr08AyG
Rj0dbzducVUO1xXnk/bdJTLEvI6zDc2G0Y/9Wl7zsVJxtmkANqEJ+3VWofdBDuQ/
zF3RcQcDp3F2HlZU7B269tham1F6KgTdyH6z2zhfb1HSud3eK6eRZw+QJ6/Ybntk
R0YqOt6DHKtJzeAc/R5Mihoe126HxMuXz4Ft4ygqttJ/n+jmG+PvTFAmBaSKO5Kg
W6EcaJdmVfug59zBUs2HZBOlsYlONw+VQe8xKBN4ffr3G1IRtF/t4ON4WkGoPNkC
VTTu7fguKdpVYpfGcpitLfoFcGJrFot1uHvi7+/8kBaMPTtXYyt9Pe2NlDyBM+kq
/hFSdFMY+JVXl/hf0rm1Behif08CJARXYTE36SGv1bZbbFPFqj65aWF9Gm4aHZpY
X4TasqOFETWlNOH0k+xgyUfPtnPgm3a+t/An6ody4F3rnodSHTB3JmCKCbjBQTxw
EIHI0syG6n4LJuZj37vHooGD3PNELUcWA8r0PrOC8yDfCrwbO8CMRx3cKKaWFHxi
dmfOPpZojFdXmnrQ4pnazLQo+l0uvaEMggsw1hi+m/c+28DIg1OnTlV8+4GgZzSY
X2cxiejbGolyrTeFPZOXjpQpFf8yFuJuhQY/uqf8oWPa7k7sBFLazFu07plbU/YC
ldPhgHSbt40szoQ67Im3j2XOOpNnuC3on5R/+58n3sDJ0tf9Ra9rb9K4OXgvbEJ3
3yi03ujIlwBrqzKTYqfMsHIHgsWVuYz6fRMk9n5YY/ZqwIjP9HutkNVMhYtaDfCm
zPvk31I4LpRbCDqSSaEltGJlrEeDHc8PeRSBOSJzi33skWOvRgknjV1OloQbc0KF
H1RkgrXMRfbI6+xB5vfZTH7e5JsRPfZpukBfdy+7EqMff8O4fbNxWJU/suvE6SEe
fMNukncab8sVQNKcNVUec/JrTHw0WOlsC2X8+NsCEnj9hFbnGZhjJwLNtyRRfzv9
sU2kE3mykIbh110499+RytDQ069wa+azmyBn3zGQY4Qji6ZrEgzXlkMdeRKWyXW5
2qoHtRtTmLYhHoORL4uJADkFDwKJrrICFWRuRkAE5Kb6Oh5Bs1A16r/x1X+upU2T
9s0Fn9wSmP2j4kc+dGhXi5T6aVTAEkfIpoFmLGg6cucvzFXNeJlMMIzJCRTlMzFF
6/U4QGcA8ZPZsU857lyAkv9exKMjYC+9+ti3DSeLFnGga+ywqx+UpkqY97Ku2a4y
aZjia/nGH7ivuZkXqZaWZYgNAd6Fsnx6sRDn4feUcQYhaW75RuSYTL1eEEKhwmtJ
hFiNgWbxA+ZPayYyEf2dSu2ouxyiHN3G2yinIEReyIa5BzNnogOttPZsv+UxsgZZ
fm/70tu5yz6pJpi1vMvd798Ph/taV4vq0laZOqz54oW0tTGBY2rEs7SjLrKzORf+
KflCOEVb7RuK2ai+4nBSYNMUN7YfXZeVku4YNbCW2USjocvAt5GxXn3rduitxU0V
xfX+dJRoX+6Debn2yQQx4S4DhbyQ8KGGqlohCskTSGjiijYSUIiQZevM+enKWxZG
rTBXeMxZ3iv6u4OM2n3OtvQnpUGAS/Z4YshZ93auV+SMd0BQfDWec2BWkUby5oBL
fH4h3OSqWxCuv1EvjM7QOHyqz0tHb1bnaboWFt3ywcWFpirz2GSm/wnPZomeDqwu
U0owXqzW01UxMYgh5gXDV6tF82eQCOpmX8nRfIbLecTBJT5K10G4RxNgEFV32nNz
z53OiIS6bkAvaW/kV3E7QKvqv0ubGdrKP4lzJCGLIpS9k2SramJ7SSh3zVgwv6MX
F8bXQakIDqYVma/mpDuh2SNs9/8sKDNMpQyc5h7/ghkWwELTmH7G/aoOZ0tblqqF
2t0Yj81uHxRAjV6ULMCPYid33qg/z8MAtnmTMQQM9cXkhJWPXhrv7ZKZvqzZ3hWK
/Xb4x+Aig8SZl0XeU7bOMCPEBkij6MYrJMGfD9W5kav6gNA/BKb5LOYCWN0jHOt1
JiXiQIioB6QI9AwXcP8bA/KfgyW0F7QnAuuGFSo+lxf6e6bxyLFjhAyKmO5jKpcr
hqCvdeMUcvrtu31Bsv25soELDHqUESOp4f8ypVpak2mrrt/VEFGqA6XoeHE5Ja0T
4Ec6cL4S3VEFwpGG4P8vDL2y2PB9qK2KBz1nOvT7nI/bDmxn18FSjJAUZLmAQj7L
npz/R1Qhnp1oxGLXQie+vwXeBAsWZR6PmlCcOPENL7J+l504TNVfSaG3GSoDyqcD
mnbZbulMEzYxERKPX1q/POmmWf5o5wYWXAVZwIEMGnH5L2khVpupS/nKsS/zm3ZK
BKqBoimi67jTbpM16Qc3KuWF397GZnxch65tjbMu+pKFEghnE3tC+pYsUcHbyY4h
v4U29hV4WM+EzonYoPY9FyzEEGlf7TPsv3MKFkvHGtxkVc2bESY4DDxvNgTX2444
wyKrHmslcuIDcY9FQc1YNfVm+ToxfK/i/G/6C91OSRa6t2WCSrIRggBvj89WAAlB
7jSQv8WHrY38HVIUxZ4P8QMYTjw/rq/ZyYs98icptCjgnhulZ+Wpe8GVP6I7wv+F
TI24+JOkJNaGqRg0BKDuxzKh9TInkTv6DzhmGx9BwsnMnBdOtW2kDzNYrde4qOom
bbyqU7+DcqUbCspbD/ZIx3NvxTGJwALy4yCN3MhEIwUMoAJya2ay0FW02U1CrrEZ
id6yFTka8InccHozY3HXE1AIqBHwCddseTJJyYE2RPktWQP9x2JSjR6x+l1OhGid
KVymThz3HTHHZTda6nP3FooKC+dg7VHVl5wO1CsY1X8o2tI+F4TGA0T4OF+ckw0g
wVq9BcJ0GL0PZs8N4awRULaEGG5Old01eVGGMDq3o47UO4bdK6nRUu2JOjpmERDG
KEmmjVyktv0SzufWLD6J60T7yK8tMxRLw1ev8Msq2cvRuK+7MuktwqHZC1aI5CLK
mydRf8rmdFmnV8tEUAxL3QLwWIPs64WONIwCt8SniWvXPnHkUFywnq7ECI/IRwsE
/ZVWcfZ0Qq3MI6Eapkf9t48ySg5hWxG+wnIcLUTQOBVk1iz/6xE3YADWDDitPMU/
PZE7N6BBm1qbyd5WYqg/nieFalQojQZCKj29t5xL2AnUboZJBKC0ct44cxWdpWDR
gB5UpfgudVXeCu+xrqzAAw8s/KVu2M7d+gIv6gtSk5947z4qT0mZwf2qeFI5Nnl3
O2dZOUgo+lFwEJIEwr+dTZjpBGS6mvrcrgoIKnvAXl5U2WgJ1du4Ya3aZP5TkRp8
dJeqsqSyFXBAbR3sfff1El179icat3Eb4vAVvPZBIMHwklniCnpOoQ6qba1KfV0t
U6BBABQeyXrFEeBnqrMIUr07HXe3VNNxqnnEtY6O5cP8P2mLtL5XOJO6cIpY/vEO
+kJ9x36t96KiNGDXqV7vB37+zzjFjpA2p1ZcVSwIKeADsLGXYG3GVXB1hu1SqsKV
BjnjLROMEZdSADHvFCCQaggbX2cjWxmWZipO7txUcP9/vMP7Sc8Cu6njT8ycqT7g
hd+9twBVvBkGBqutVdYNJbQj6PzeiTCX7XdEIgaAu3ta9zG7BpJ+LBTIBgBEooz7
ZkkjctFJTyD/okf5Cg+sUpqgzg7FfP1O/Li3e4ID5yDkkXhQL+SDeuc9v0ffpVzk
TLc9cUTg2l7MjwaKL7RJ0BBWjQmJw8BKzR3Uj98Wcy99yOVO1sK1PZd2pcV6RS+1
PqDxwp4GOxkU+WwSDBoBwACT3AbFxwOsJMeV7cBAmY+l8Y2TlvYbPv5ZMQa5d6Ds
iNoJwaB1YdQq2MTn82JJWarvw2uv0ArBII5krpmRFIZQKamoQrj9pSSecXSlsfll
zJuXWwR9bCBhYQs/YLjoGH88ajqOU4OS/A1HdSaag7UmgEh3fdIzzPYfNfcW1lQQ
q1V7YHR9CxbuYpDALxwQTIp8c7fz8PdK4e08tiuHpX8E3O49lt7Igqo/g3R97OwY
2f+z0F0rs/BuQykY4qdJ8MjlbG+CwHwERVoz7gPKwUAY5DjGAJi4s9JIrMUtb+B8
s0RiELP0tNlCTXn0eyXK0K1MkLnZnookouIKKM7Hb8rwDNROlyyxvEq6Y+z1Ly+X
BpOweVC+uUEewkRbW8l4BuLmWm77xB0+RPoybiGVt2fPdxkVeUyXcDp1k9tPOGrF
hVGSmqk0bouWTJS8X7zrKw6AJqa1d1GP5y4ECsd+GMlknQPbAmUF/M4BMbICwLUx
wWzfXzOyhaH6bwv3CTDLF8j+BlH7vMwSflHnk1XTzQl2Dmsb3yYxawkWuigu3L7P
+Q+aMsShx78Ttro+gOLbEuXCavpL4G9eyGReIpIU7w8GngFaJZeRK9liKiFMqjje
fyisIdqAuX4d7RI+OLncSQUPyKLC6fL73oilfbLOIaiZn+REWiFLZJ2sFWWMctKn
8LnHNLoRen7UbUsk5WnArpbx3y/1PvT4vDcn9APJ32mKQikEF70ut3bbf64TGrhS
qH0YqxtTuyrUFrDauyEtJoGXKHA3jtDUtzTauiiTsaTdyfHVHrQytfdYAqFItk5D
PDjsUXNEnWY+Sne1iakgSmXMjBUikWxRzkTDw0emgARMh1OpXi+VNwkmoIIgtmZC
cdJF0aUOUVYlt4625KBxKYMzCAbhj8k/jRCIdMBJWXy9No/OPVMciTY9v9md95AZ
Sz4WKaYJJDv339/3VYlt4s073kOdWuJHGu3d0LQhrLXHvV0UJCYVv2xsAJmLCaeH
B62zAOUrw+hki4oSgpeUTQeoxv6TWLZm/5tLsNejx2ENhsPMh0pmRRUmEQ9CkABi
e6uUiLparf3HpmF6xky47LiiRGzXJvD5+gSjfyEJbWeevLVcyN6FYLkfgh3VNrNs
a1XMvPIluooyivtdH7o+AZRi/eevXPtDxvp9+XBGKIavme8WWLgxz3ZdHVI7VbZ7
BYFu3suHJqjXCE0A9U5FQ53QyoOj2ggEf+/6cpGhEBdB4i7fTVU+p3uZsw8sKWwG
El8YOC0HpZODUSjcZSfr6gZY0Prbw72oIKCyAk2QyXIwOp7rf9WWiphbuS3/lNQq
Hhk5xowxSqw/wSfZN2LcXrgm7+gw3XYOGswc1ey4kc9t1qj8K/rPe4+S0A9c3rcY
yclSB2Nv99NuBq0f7kRlGVr+SJbZUxTTTIwTYGv6h30KsKsUdQj/eCIxopKloIUj
fTwlgJomsinUh1gKz1p3IyL4H64lYVfzHy9s2FzuPzgIfqevWo3LoujmVZiUd4cN
9OyIxMbOgI3YUp11QTh5Isi13xapgL6NJILdnVxnagg1dEeEoHCCzQRvk3kRYBeg
V0CNe693U8yr1awPaDoH5u/EozCQmhiJ9clHnDtODQ7b1fdnHq3ncJ4qnaJ83DBx
teH3b3lAaMsKTIk0lc5VXvkLDRXE0bneI2nLZmupbeDvoLqHqx1Uh8s1h8oWSxyW
OukPnmTsCejGqcofgQtwB0KKUAlDHOyUJqPCTwKgeQYsUWLbJvRU8o4KDsaxotKm
CDlWdMSDa7E37b47ejQLovQb5uhE3jSpRzDqN7023wbp1Pq4SuTMvc82LI4FXOh7
pMySm9kgyhCiBUTlh9j6KQRuTH0lTA7MVwb2Gml2jsDTX7Z+d10LrmcTfXlUqP+f
X9aXEXg7Yigmi1nQFNg6vdVICR9bjChnLdGAIWAe/ZAAuaZQye9RGics6IybKWg6
3SnpM8U3pUS1qekiaU2YpGnbZzMjhxw4Y2hNAIb2+tfnCJDAudATBeRRK/WZS558
mTwxkPzyOSURor+3D0ia1k0q5FWQaYCKlesCZ/yFt54tJNpTWCiLxO/BmmXK1dvE
8Sxs4KLEU+rmcYgkLHqVEIMg+2rQQJ7VzLrigMLNqjXzfE2iPNB7kai8N0jbCyMT
7p+KI0FJU2Yk4GiwD+OqE40sIfnciOWIdCHTOKuR3HVNMgjTOrpYAlNTKeTeBlNJ
JqOIIi1QeV/iz4vdz9T/1xjfYPD6/G2laEExs9fahmlTPQ83wyXHvUQYT8M/lneh
NAc5kSVKTu0deykNZpRB/TZVTCroQg624mWTr8HxMTqezVPTXDJ8gTF0m21E50zF
Ckk6l2ZZMqNeREl3kQV/JS1vp5v6nsZk0rjs6SeUsPuZqOlirk60e99Uc6JjUbpg
d16UlqJx/YKVQTOybR79zTxlCk+5ev5TUt0cZqXXt7LpEeUUayCNmpMQ8WF6jfHV
910af+uyvEIq60is5vJKXG01mLTA6ouA6dEnYvhBDHho7/SDwXHgmha0mcYjRX6p
pd4w2ojJWE0lUqg5E/bkMXW0kO2zPadUNBX+lyQcFFaGEeio9Khql7b+YwJDfU79
PiwfzzX18c7x5uGbW8b0nDZupjxZHEl6fmuYKdien4ecqpXg7X3VV4ImEUgwwdjF
FWf+sCrECKEOcbn0lKpirsMXlvJOzFKIyjAHPh7989gEARaZmCVq0VEIqM1E+Cdl
1UDruOG9iIexjr6zFEhLHf4zKwySVUTDpCexxOKcdfNMeCNGL2MQAV/BdYLO0h64
wV/kerug1T3652V72Jy3Ux1AxCTbHtYLiaEX0TkjZSwFpKbbcu87labulMOr214v
WjXrf8noxsuze/JgUXPt9+aQrR3CIbR4/zqwXlD701PeosU3Q5S34BYeid/03Zre
S/hyNVYYdWKQ0Js0TS8NUQPn54NSzujkbAfinHMx85alBLqqibPysU7K5xcN9KVT
sL41SBec4XMBTesR+mxIDHOIKJ/A8TFMZsoKU4Hyl/i5L4PYQ1g0O9cjgbZf4n/b
lGFZ+adKYFpv+wgoyPAqILZDexz5bdMJoXuqrNALNzhHdnEGEYmrMFn2m5p+KalP
gJO7GlxqBkfUG1L5LCubrT+VGbR0wqV7QdrWV+vVXs8tqqCnC5liiUAf4dUX/pUa
iTlGJ1BWNihHUFcWturdLfmyZ84tsdF8JDHYWZuvMtTk6KY+pS3GnW8I6U0LGV9n
B/BMoo8cIaE7IlxOHN+4K0hs1GBdAdbymNGsJIjptdooqxF54vPK5Ulh4skVMsPd
8mrAewpGC3Mr550tZVZHC8U5NdtHu/9ivpSSAt2uVzXryevCaWtsoUSkPEnAii9Z
FtSsk5WphLaCKMw0xQrkbcM3Vn/YKI//a+SrRTU30gvJVrX8ZFurW5ymBOw2b1XG
PJjjRoZKXD2hb6My4Q0abSvB1EKKKfRYKPyQzDgcthVob4jikpx6vDOHeutteH+H
SoAVqKr8Ot+moaY0haM8Tr9z2ROOophr2GgMktYe3w8NrBDLubQodKUc09+OqGm7
Aif5lu7KhxcuchEKJljxFZuSKooWbnZz/IMrnvFOLazp6BT54lamob6EfBQhWsV0
+yI6DfuEKH86TS25YFyi3Zgs1NDVoop0QOdzaWFelm03KEvsFh7FKC5otzcfaVKN
mAd3DJAiUC7zfZZm2GplE4FpImPL0RvzAIYj2zjeXtyozzp0cKBGXej2xs+NzplE
GPM88DZwF/z390QKMKkSklGpN80DUzmvD0ypng0CS1yqn+pJQmXObEGkW/TzE+d/
gVnpbJcHiKnGYKTdwwX+LWFIUU1kouJn+57fd1SZ0+QHFvY3kuHWrvHWH+OymI7V
GC2pWicuWwk08cT8uyTY0nxbq0lRY0hTXwpu8dkLDiNO7GHw7zxkHb2RLUCyVF2P
AFfDMWT942J2QOJrIeuXCGvhoZh7l9iHyVQEXivvh0ks7OwZ9mF2klQ5vr5LiYfe
KkfoSmvIzyj0rgszStaM12cCyYVuz9H3ZOgQEsxXBQ2LESX7p3zYJIMA8eHrjb/o
32zzuZs5IZ7xaORA1eX3WakD4DG3yrKyvkAb5LP+AW/wesjusDhBrhfzssIn3k95
srArKiA+5ntWXj7F9+DoK+x+UnXDVYx2WAhtGsWl61YwCxAWXst4dvl5vGDljWez
jvC/DZTPeFAjs31ZQbElnjYy9zX12xETbGE98r1BC5IdHFd+T0J+kOyA9ceQ+hAs
WsV/+KFGtqNEv6KvO8FpntTMaB9d+lAYB6fKmj+G+ajzfLuTaejpzxMt6enxhtH3
ciSrf/gVQgFZE1E4k6yXuI2PpMatVIqMvqs+jD20RWE2dDrAUhYtFGTwqfhro+cD
eAZYfQEDSr/Z7zH3cINm++IMNDylpKs0vvMZVdpyEM16gDgMkexiCPpwc6qwnR8+
cxq1Imbe4WrUUufFqNMkAji9CLeGJgAZKsHob3at61Y4El4QUfROMgmxy3ojmoDj
j16jXXmFYsHlHWoZdgwEjkdjBz0FOyderssCY0Wim7zmxfbfx7v5KPc1dJyQpU+G
PpaCYQ45mRxiHFFFrliR3twkh+92WMJK+g00+1hgVuBv9bV7rb2vpVyaX3Ns3kHk
CTrMmLC9E6cocZDfEb42adt2dRuBnRAygQIz+BLFcfZuzi5/16/fYh6E41jsawZx
QJwsMdLO3SdoIL+4VGPJ8oDFCDz+ZRkzIxx0fAnC2QeacTLxPEbCveepl217/G0P
/an2usQKaG29OplwkGDwc3J0V/T216QTX82bUQDGCP01jYynMvPhnBjvdTiaSXcP
MXj2emw0vwuCflPRFOKTxvuQDaQxMHzf84fupUr2rNScQq6+FEheVorhxOzs/u4p
CR+c2/j0uUJaJXaNzqQHowfdslSIzA964ykJ6u5u/AnrMueyau2BhWM/W4Z0uAPZ
46d3QXE+r8Jg8BiZaLcmfsUtEnqDi63nZIDfRvtZJ0JS6FKoigDsl7o1nYQ7gQyf
LV1SHQDv2GNfmxq88hxeGt2YRoxvFwJXpjutFJZOMuCBH2DcERRiR99gcW8cAx0B
4u7XC2PsGGJAoLhYxIOYtpNCyi9pMYw9s+lK+avJSwAd5vszoN/QYmfmHquCQF0E
Us4E9XEqyYV/9ECyq8qj0jwWk1BpCnTLpJwNav6kPSYFPHoVulvnwTIBHUBNnNiK
qA/VadmwF36owVcGMqplJMFotrMvpqS5nZsP/8qLhRRFESE2XOHyMaR/2AFObV2v
xsSdAQ6q74n8tObAXQ9Gff8uxDma12NoXZfMdSItak4o617pDfYBtmd0Qzs1jWZw
dlXiK81LQ5Q4m0suIVR7S3W3OnCGPr7DYjXh4DCuWldKl0F4L4xPIHDehQsXliur
jeHnOgsTataeNw4W6BqBrn76X4kXdSEl83DGWGO3SE0JqkrEv640lsqK2Ko7wHto
uyO9GGQ/usnmcT1NFCoxoUF4zj6lTdvv001jhNbzbVyx6k/dHx9DbsDHxlReK3t/
qQWSJkeHQXIu5sMHl84Mr1/1ajhaHCtyji1NjVPBqkl6ihpKMUetrmQ/UQHljUbu
pdAXgjaNJ4SUo4k07zLNYYDuFtCGt3eDrEI/YSf6LGvhJ5Thf4JUqoVj1hOpJ+zd
R3y3f9e7lnYPYDzsKKBDoLR8+EoG6UG79eAt0Ln9RQXIAPNYOrESZAWN4zFy66ZS
Msh7GLd7cwphDSTHw2vaimkCzLttGl2Ckq5LBpp/6vqaMHa6EvLV+Mk+vP9K7Q6Z
mwXKwdGiI2vwGNhTxKDGHLnmbQROhuIuYDHFpRZDTdSjSZPHP6WB9VvYUuCijh7D
XXPsWyjTclkTA+5xw+EH26PP2pEczMXAKxNgawgg/2RTjJSwTfuOXTs83ymdoEcM
DLlko7i7O3HKv9bPuPDCP5Orvn9vAc4tgD+AN7Tquo+2ZulFZnOgGvwBtPqB48iP
kQITvIM8e3V8Ty5HMXa+gPXNZHsnQoiBK7A6mvneMrv7DYQ7CXmF9dD0Ua0phbHo
8N9/fD22uC+WTjyrTMTWiLEFe9LIpl9Wgdr2qwicP8UXImQcGWj4hasIMD4+tx5q
bZQ9FyeiHpRCLu5sQTw9R9NiACsl+LcP178wQOvHk6+CXWgZm7fFyyLy9LSLRJSW
Zqgg9u0zTH0/0Znk/snWe6Ay7z2Qo+gacXY78VV71jMZpy25ZGqmusxpyTa1vctU
yghqVeJMJn7aHA4M2eZ7ydUJQuBrqKos82Vr1bc/etrZqkcASDDf7dZySaFwWxeu
wXbBo7aXDuX57u2LKeb40vWyFl6o9p1C5zs4TxJC3NaP757RdFWycU9r3n+jw+3E
yHCMJ0yZHMDx73cEz2xZwjcaEfrS1Mob0MUL3FLwmX0Af3yZ6nZv74a49BvX2VZV
TKhtkfDIsZTdywi6R5Co7QaJOghQwkcFggTXCMNjH9lm1qOfqsG2FrMKKhm+ijbW
XPVhaChiuxNdMP0A+5QBqOJFR+f5fnMddayRbUNHyBhIbdTpy083x0kwy1W+y2tP
FC29ivdlT4m62Mz/E2KEPa/LY6QyYroHBOyYyyQzWWv2XPFf7RDRtzLM8iiKnMGl
Q8RsCiRhQlvum/TTGZaoqiqerElEX/uWOG0V1/Axwod2/e1cUjWnk5QSdT2yS42Y
6hKvoDsEIBTzj86aDKUkpR7KgrW0F1o8RLZ/pE+aV6gyGhPZ72Xohnee1I7kP+D1
dtuzcFUi2idMzyklYbJGVehSzJ9tc0+YiHXKzkiJGvT3pJtkR/2zGURm0TgCFVGN
WQoyfcd/pR8e7ex1iY3Cybx1QVrymotklLSDNTUL3Yb5v/I+tZxQ9WTFLet1GOxf
Q5ia5hQPboDYpdWP/9GVr2j1UNvj1N1FXiJL+b/s4FD4ZSqwYVCNdC7S50Ce6N5e
b6cb982fnywNuOjCu4mfKTL5efwA/IvE99+YEiGzw5V+JFN8X8+VPOxvbJxIJp37
mNhw9z9knJMk9UylSnfz2BVYzZ97epH0n9STLN+44fyqTJDXU12V/m2A8VCZ181u
SlFBGtRgGe+3wodCIPC19SLv24NkeFsyk91OmZtfoqwXAnMEJPpTwqUwY4y4e/Qz
M6k0dgjN6ffZQHefc5mheztJyHeLpXUZQJiTmlNEPwwjJUDJfcuQ4o3JwxNjYRJb
qDqKGHgsF2L7Vejf1D16jFQIt3nuLBsXsf3ICSYseHfQVF2oSxX5KreaWymIgQhK
vdgYcTcYrLtBrmNkMB8t8N1QFt3FHNBcPZKA2IfAttnY2BzURWAQbULkin1O3UP5
nD47gYdKMQ1Kjni9VaufbdJ7vcEbrfvOEx6Bs9oRizjl7iUlTPHzFUlfB8DcnEtb
XwHPhi3S9pn6yiE45wPw01LbUxHPaflwx5ovhaSeQK7xMQa6aBmjvlHWiRvEr98Y
4yIQ3OSi1TgR4pHuKt/HaWCRTaWP+AggwdNBatx78KQthULm0dxaR159N8DTZr9w
r1AGbMVhjqoHFrSHbXCYy2sxLGKFCrqwOrOnlYtT2zd/zp1K2zG8E5S8utVkOfml
jRWvN+6uGESsKRZqrhQoO6kMBybfe3JGvqK31XzVy4s+ATIIo2krw+jys+33QAdW
DQ9vQ68qSvC3TsDsrapuScFvEBnGWivA2Pq9r2lfSXPaGHAm1VVo9yM9sG3oVWw1
yt73gPDy2UvoYfqzOlQryTVrYZW/a0r3y8dn/j4081v8CZJDx8rCEEUR+DRbJk0Z
tUhyEornoRdCPlBN8yblZIa3G3ErIRFNehQZmtbILP5G8UTJ35CKjm3S1RPDJG5i
z46XavIV5IwV9HDVrP45Aqt95mCChM29l+VpSmIREERbsfR3SCiy0PI/HOzv+FsP
59BhRwhAMjiduyEtZf5/AkS2chQCshuKWPUtA7k6haASpn0/7op1IZkQQHDY8jgz
zT9RZ6ndf+RbikTwzQWZCh9dzIx3h2SyimYycWZEu9xt+yh9ahoZQx6o0ug3FeXH
wcHShhCYFk38lJVpITGeeTNxNzsTD9345ps7IsbXBn3LPP26xMWgQlfJgtINMTUc
clV+Rdj1FBV9uCfnBamzK7v0ECqjP106l9b0VxXGpzOy+w47jwPa37dM2/fk22jk
VFEwbuVB69P2dWG4E7Ia9v9khdKSLZrRRGyogrR/CtDhYXf+k2OgUfE/VFHU7CWD
vbU9mMLUyAGqK2TClsYCfzVcZqznG01LxE/FqIDlOTq5kcoVuaQhxVUunwjlMTrz
WhNP16qJ+VbDX6v8WpoFf9ztFF3PzUub67Nusd1+5KSQtdbhqY7lEtTTWqxJvlJp
vU+oZcwIlMtZu0Zg7jBC8z+5GX0cKaE+y/3ejC8xKqjGqO0XIuCbceaEhRp3bF3W
sbqtoeXKpPyKn45vsB8cyB4u2+tEiyMwv9hJ4QCDcL4H9mCAKbevZJJ+d0nIh3ep
gVcqNiKce4IPSXAoLCUy4g5KdhGpG+BOUixKFAsYSMGTmQjkYvd4Szej7Qj4PJw6
C/nWE7vlgz1rdW0hw1cxrgBuk8/660upcE+rpopYGjSIXB6wu2JExdW7wdThr9u0
Ng/DwUlByhYMEj6h6bQNSVg4PBqvapf/4a2eGxKTOnlQ59f5qL9uvGWAcd6WldBY
9zHNNIusdrEL2ecHbewkuVRKuNYU0I6qi3vnkQqCbAwOkxSkrVO1R7YtRQtOo0sV
M/Q+c3Ztz/bmnCMybu4KK8frXXhEqhup4CelLzhU3n5qgOMrK8Uw1/M0c5fD5q3S
rt4G0ytC5J17Q5TJhUiBF/khUL68EroBAEVRBcPV9daNsXSXUyaVuGvIwww5v5TW
wFbrGOk8VSLEnbT7MCwWAgH+sx6SoTmR4lzExZKMYay7H9EknBYK/uMt7HR1bpUb
k07lAw5vUennyp0XHiTrUPd1+Gl/I4ggeBbXyJjy6eBgpkWMtuf8Vod5axUBY0Kl
5wsZyxi4Ti+RvZwGnLsWKPXcP3Qt2QKJiGNhEAx2pabZ7+X1Gu+qNNIZ71qpnPIH
NUVXI7ElcFOFgYgmMFvwNL2iMU27twNh8tEo2waK5Y18s02Nex3+XhMvnq18Ry5f
dptIABnuMpV8Uv2WMRqlHNjKdIiXOhT9GsVf5TdcSpekcJDKGe/iw13Fagp7B/iK
EYIb+TtSN4yV5Wr1wXIa0bjJ3RdznOVw49G5rx6W0GX9RsOTucGLt7a7Qqp38rp7
XI2MTEtlI3kCh/WxVgt5kznSVQlb8OmYM3y74Z9fe8q49MewrsOhjNniMo4PD/Z/
mSBACJQdTzTugDgn3Is+Wgo7FhAgPmEFsZP/ux2S+V6feZRcf3z/HMpZsQFVrPzT
SSxgX8wjxOQothJX4dmUGncfsB9qxQdgYNkFm+Bx1pJW3WyPf0ehSdOgitpELV2c
8lqlOzoXzyHDD5fhnL5hJJd9aqkdDY78DWOOAM6Moq4IzIM3W1GXi6IkZD5c8Fn7
+9tI6XOg9oykDn7Wcy+ND9wFZOh343FdYBOEk6p+Oefi5QWHgfZdateq+UDN0yZK
XYWa1avMAM3UZbLGI9Dc1MRum+NHH15TqKVlxlJUhecC3ry8Xv6VFQJsGg+9Kv+/
q2mTrPfUCLq08KST+AvXfHgxZapuFO2eXL64X2mcFYpKMr3nf5S4driYZ20BJgdg
LJqstuxRuTAhFOisYHa4tUwfrffEhd7efJv71p+bwdhOX32ekb40HOdOM+m1KF9O
4xqW/nd8sAN6EqaVf5VfQTJXp6I63FWTbujoALOXfrIyloXDNpdJG8M/rP8BEW+K
KaHVX+H5aCcBYKDE8JFd2f3OE/IuXv0/LBks/D9Uw49Thpq4AU467ipf9Y9nEbNS
cr2EhZ4WlGJqq/CWhCfUrZjfBGLmBgAXEbHoy0q/mfiQU69SvmfvPxjQ9hQtkFSY
9QLa9X1+qSRHFfix9q/JA/rG73RRXELX4m8m+EJZQ9gkvmdT//zR0BgAk4vb+aw4
IeXmTygVw48OfRfw2MS282nsddLt0UvVA8ilnmUjsQHeH9O5Ly14ZYQFMGs1MzJa
DRIcr6q3HE+nOGndXPbsTgdB6jprcV0jLtS4kZORtZsPDjNK91lDqj5EhymXmKg4
mSEuPeuGAcpVhZ7Mwas0eapqMbc3aaobFnSor2sQ+o+RNSMF08OTzIXqGP3kBkUP
nO/5t/9J233uYh0P3tVqGfvyORqazYhfBRNXGRSSzuaAScCCkuIwkTBwFEvQ6ozR
6MVirxw4ulPdbT5+6ijeoft18+kWytlDiss4+lK6WDL8uHGyVqld6LVDD2mtmIzT
RqlhjBZRlP5Td0+X0mym5oD/jJpvW3i0VM+97egCE8BMeVamtR132ogOTk/czgdf
FeC49z/XlioxEJ+Qg/ej1AeioZZPenvzZa90aI3PQkn7TRFBoV7I+RXh8Dg0SxVb
qRiIquze/6Lri1KBFYkduL2kU2qBtruLxT9bAlBJmU/zAkCZO5/I1jNNY4/FJheU
M25oK8ntavA0ZOgWfjt/6oiVXg/3WwsI073/snL7IeCu/bP5egCuDWt+zQbyjuS9
/muDrX9kdGGmwZviqqUDoIM86+Ho9axf6tBvA2LHWFUcZbKsWkdwfeCkcm/p6KP9
omdPCjSKZitF+yLpXs9urACsLOfmkWBzzeS5SOamOU3K0P8L1MGG/YWCA0tlM2m2
mpjHakaHawrKXM9yqqrGx92KC0idsuxuwznCQ+9U5pNB72RAZoX+9apjLOxxPhuX
DrOgXsWLTd2X+0+Oy2yNUsztqeA+ltO/BxCzm9vXehFJCAaQzz4gYcxejhTsRGQO
y/0HdqCpkdbnT7Bv1zmLBbI4D3w3nptfny+S8Ph4pV8UF20nK0tIrLhr3szO2w4f
iIbwvuvcR8WIKZGKHI/LwpQvnFLs76+u70y4D5G8C6BAjxXV/QWQS1h6rB+aTP64
7tNYPMzua0m1ZePoaSkPGpOTc22HUN/mQFJUPMCVeXiOvVdHpIqz5PF395jWYsvB
/bR7h+ueH0LHqGpApKO42HCSe1Oe9JA24gocxAkeZsMitPwXZMV5SluOoooYMU7V
GB/8o6AXNEA7ZH1cdaf+VVq9lzlvxKiPAdcIttTtqhaUZWQR84xTUAqH8Zd5BNen
pLCOgnZvml9GZ/N6BaQgp2jW6vo8blU+JgrO4rQhsbmcl9Mksi6NhwjOCwg8Lyxg
sDP7XWUvQ8qCaz0fcHDXDehIpB47Zqa3JXJ2qhrV/CFxULSE6lE2wlb7IeAMcmWe
C0KWvMEee92nbHPJeOGZeK1tTwEk0doKX3umLNdL9Cp/GjbcOq6/ITNY/CM3Ps3j
sBwrUJ3d4vGuFvLgYSrw7A8zTmTNO/QMZQuTiL75XYifGl3u2toS+ejwrvRKngDN
Zfa/Fxh16mohCuJHeh/1/PdUFGVSZ+5THPN77O2Z59WwG625BPuGmtWKAcbT/r2N
I4rWonSBJbcjuPpwY7EHyfqmQw/honcJSbYM41cse9Y/7FrDoqHwPH91SDa+HRUJ
lhkWu9j+3lwK29xuu2FCK8qaUYQ6gG4Rc3YsUaPHz6/28MTySOo2oFtf7GfOpBGy
nGKUHrVGXxRy4idBHnZ9sX5MxGtkfFVx84h7/jE8smHUf9IYVP2dwA7NL992rovR
ld+6Ws702MJ5Ytk7GuoTO3sQigrCEd8fHsLEzN7llEeyezaim3PG5aqEIUrCXro7
zit7dZS9LyWFgEMBV9zPwRmNGa7rsjvsb13OX3l0YbEBP5Czmr+j2KLMKBbri8Qs
lTgIJ2JGL/tuoooaSdxS1eDSN+LCXJgW5y0JzGpeE2f/dlivfLSAF7/hi9RLn/X1
923aOp9dzjTZN5L/t5tlfECy/4KlYdZvNpp5l13rUK0w6DvoV/vWwYVf606yrKKK
vssJaTYZtgjqc8DKrmMrnht94I/f4hQJraueuavn9pe1NOm/Ox3sWcF1IWztnbgf
b3EBzvjTRjOrnf3dGY0Y2ZanibOi1HJFpobJNQwFdYmBXRyOWKr/UQpczGK1Vyhg
Y6uyfd/5CsM27vP+zmHn/yVQLhN6XnAVJTofvc3iM61mKlvfxdblr0I9G6RuGKB2
1s3QHduXzhKQlwAAfWclAzvi1s5/gw8HuMrZ/tfYnUqW9tXrGW5VbLIqwAwfEf46
SvGq7fvTXJPli0e26tdVDjgN6RLlrrjl+Z9Wa90RCCmC4vVzLTjS/bwfFr9bbbD/
yvDnckJrh57JNNFcuQDYsaaY+fPcD0R11QED3spKjcVPWGUiH6g9s3xhbM+PP2yF
qB88QofuJBEqYeeN8LIn3er3U7yAn7VJGMGPkdQzswQ1XDjlTfdfzn2f1aa/RMvv
wNeYOpmp1AozTvUc41pDcuJnPis2QVqK86ehuaIErYlO+dDoiBRYtiYL2LPYz4YE
wYVahko7fMyA1F+X0yxJVLeJtYuJw2KBHnoGIjqLUZJBWrZWyZkBSDOKim+ikWUY
f3VZtFWdCYZxemZ/zw9483XNOL1ZNtO4aL2enStxc6TdDSlSMLjQTUlwUfU+m/fC
aaoJUw/f4iX2Rh1g58fRDaJDxu0/bixIaj4x4VQ3AkLNS8BohN9HbWrkRaB0enYU
s5bmlpV7OnsrLA8AXcu8yorCvIOIGpl3iZKLIuXvPa6stAp9mcRfM+Ta41Wge6E5
ZUK/PpXSINfGjH6PAVx2ShQyIG1gRFJqx5xOD/VSvHgSUTytHaP8e97j1BxNAehA
xsgGzlLjJpzXNX8NfWxi3NIoIXpoxxcFGyXGiSCKGCk14XPPnxw/n1nCGUFImkwz
V+wUNL7PdgmVoIux8LAFysNOxLuLmqCTiKsL5acjwwGHwtIw7jMrVTtcoQMLp6ZQ
ElIN1y4ekokreyT33+V2mAzwGcMYWjOcinP1NC/rpSq60CIA0BG+U8DWOmYtJSsr
vXyPauzGsJKDRREwsEArxXM6IG+F+0DNEWzc+lrslh4hkE3PUAKvdHcZpIQhHGh9
IJvo2krSBlId9a1NGsxKUwO4IX4/FieWRVSlcmtj0jkf3r9WnBEcp8E3JyvbLh54
MgU4DRY9Dsl0t5QGePr0UqGc4F/4Ag+/qy53bN2tZRXgwZk1fz0VYcT0KqGGQDfA
/KdIvwAl8liL95xk8y2aMqDrgj303RuONvSC1TI5GluBHVEdDgYlV+JwS7ga8E+A
+PRRydKUjaBybDVJmZrEi902E0aC2pAumyImTXXSVT+a/AHToxjiiF9+ppvuldF1
ZyFlkDe01VqnLiJpq254nDHgLrd6RAkxymLvPL8+3zfmtWqijRoBa4NPXKFDLEhY
E6l8tKMIWJXjaRxuszhW5rGcb6ACfg/6KT7fsPomAx1J7fFiF39V1C5ASnVpthyD
dX1qIm6+YL8S0RV9TvhhCDPf6nsAXiE3aHxIkvYiPVqjLugqpRu6clfdF/aZuR9b
uKqe38xP5TNQyrhBXxhFtSKOf/Jfmyt02Ufe9plyahPBWdyXbwu+eXcFmDcRGBWI
bli+e/aMjZZNx+m68sR4bv7gI3AEK34vCnOB9RStJLD3GiFDVI/b8oYcCE65SIbZ
bOQx3RZlLPvCuHF1odnSIXSjtSvJiuRs5PKB8Uik0+U4fHvmCZKBfrhxd60/h+ix
4jpFqmIUbHoz+GmAhzBfAOi8t+5x0iAU0Ad5wzIFnS10nKifYLfrTeqd6jnpAh+O
kBveCV5vlTBfEiXrsr5Jcf/wsGWfCfP5Kn8MNz54frfapGOGbENdVzdsR5Vyn2IM
C37xrg26Ca1Af7iRSSO5M6kkhcSVKhPNOJqikjlQNaEMIq/+prZ8gsr4KSJheW4i
ID/Pwyvil+JmHvfMXiFBQFOygGSNsEWFUn80nj5vR6/ekba8Tdf3eLmOb4DCYf5J
ziEz/9AMG5lY/zUjvFBqzUhen+1hzY+xAWyIhadwOoN21oBPiuywvtGp82nxS4pn
e6BoGBxwO3KODCpLKA4bBP7isEBOCvgfuW2nmmkXcaxgcg/VEGpgOVvvLCv9h1w5
blz0nlyonpxBSROxViH17rY1GUEVlqHSwEZIKxPp0jNaLD7J7zObW62g6bSp79ki
GCJ5q6RpCc+dHFs6x385JkT+pTF3+V5aUG3D4MuYNW/PMmYEoIKzS40xdWR3WGV1
YUuiB2EhWx6FlFusUVc8em2qy1IkkAjTioMw5Evkmm7QT53wwYc5vfqycnDTgQMY
Ur2T8DtXGl5p1GJxVJjAAaX/wN0FIvD3AOFtwqvZwNOQ5SwXBHRYznOR5BmFyLip
Q7aCYGrd5ytQ6jBLnaPfbWrXQ/YHt/ReURTL98x/IzeLH7FwdYRTF4+bZDL6v2rY
muIRzi21hsRDjPRs9bqDQNdsK/jCeb20VXEUMoumbm0snTigi4enGyJWIFH+Hjhg
p7x6iMb4H3NhegwYvs5zq5fgzOPUKgleIVHpGJKIgXTa7c4Rz8zsKj2YkYyMX3Bb
6/BW6OWsu4vapg1pZv+4dZgQQ6FLty7l53+KJR9+yNnaGpVDnSZoz/E528vvrbW7
BqCLkllls7pdPfqs7EP8XsuJLOJPrfxPeZqMnQZ2zncKkQzgXxmo6o0FVWbnsR2w
q1PbcEfRCibmWDN3jfi3bQ09ZMWXPwWLPr97MBhhF7ieBV6ZURsXr5mR1wRIRAQr
b04w14xUyNk7Wo69lmKYtlTQS9ihBtBA1pxB8hxUvoNcrzwbt22Spw43cZxHO+aJ
idfEKIqV/6wq3H4D3y5iUy19jTWH8SYrdJWsohkqfsCj6EHjeJs337WblmK2NfoQ
32DEN1EMbBalaAPe07Ys0VAHZKbbRKrfOxHjUKR5WUTRCYaMspx2eXjQnsI5gmXt
5P6k5GC4cMsRvkeBHu3T0lKdWi7wnEQc+RVBTzaBXjEvZNpHkgcrmF9/pxNRX7xO
gPBbDkfLFRFOq7NHEEjdcX5ZLTDV3gw/2lAEoGbbkZWCvm6r7PIPZUKtmxcpNYa4
W7VydnLffByg1eczeAql/Rc02kxQ9BHhFWuh9YbnO5/omMNgQW8SEaZUMF5/SEn5
/hacttvBt1LOXUnm+hi3fKN6w1l1l52BIth8R3ywfYGF1/xB9fRUstVce6WZhc6o
Hygw9xZDWYuU39JIkKX0aT2drDRBUDbkeE3wUFYNDGHR+ttclHMUbUelXq8BU/dC
VO0fLjOfeRqR4gBdbE6UcUBqud1U2erTMilURP+KealLd+1va0kv5aokxfCU29tH
6yi51wXJQUqF5bfaEDLjxcCtHk/AigpdAIow0YJAjzHEpbCa4dgB15+pH26Trde3
i6iBHdb1O+k36f1VDCNWjJPFP9b8vvzKLW3XpVE5AZElMmaZmjmxsBL2eyvxphNo
tafI6lSVSc6n+48wi469gAwVCOebDGXbqy8ilMmvx+VogOv3OUNEYTJ0vzMbeRnL
FtqNQyQuoK6BGB+aWXIxJBxAk2k1sJctODmhQ4kgMqAE2zBED5OkNLCPoMYJW5uw
gXfsE3uDGBzKDNYTjV6YyxwiIthq5nNwzU0kzmTfuKa5ae4t0qlem7rry+aqZvw1
ediOXU9+SYbQCU9NuPTuZeANSE3hRLYAaz2InTs82rPb6Me2+FRnBaKZm6O7yQn8
coqEwiBV5YyJEdptzM8hsUa1GgERQDBl/wWPtW7Y44GjVly30ai1bE6MNLr/5aJ5
VJkzSqPVErq+wIJwKawsIzGP/1KNo3jjTDVVwnujGMyyR6z7pO+ZKfFFQXQekMmr
SaykSbCOQL9Bepxi1VPV+eRhsrLwZU5zssa6W37b1eZcj8JQU3zcH4RFlmlefcIP
qYYd/yA3/uzHsLVVu1MEM88TdhTEM2z6Fk2DWbxRL/twDXuQ2kQw4BeUyyY6riUf
rSS4nFFT4RbTC4ybjsLNBgmuFUok17fSCfsDVbsQXpdEsB9tHjj0eOpIoUz6HAtn
+o7t58C6HdoNUToF9OAHIGv0fs7sQVQQU7N6skuncQ1xHgq9h5WE1Hg6niussmXb
Jqzt6GZTyURTDP+yzqXBs8vdumscvLjtxnuKa15WvD6/xcvWdJygHIw1BzMlSWYb
XSkhMVwfpgtYZyE1j/PROCY/rDIVY5uI+IiNJfa06VFDwcn0/yeDJ6/ZQXW9iRsA
qBtFKjTEB8c1hG5B5b1FCc7KcESnIkhIC771zsf5Nze1aveZh23eSLF0uhVtBK9p
XCFEFrtl1YFzvV9Gs0128oyc/P1kB7AaBmYmZOOClViNEYsjjMimverpY6Q6ZVL3
J+6SHrGT2SFUgTfOBnes3Z3rUjj02+R6x5znc3xHr6B7UffC2sLDcjrjC5Y4XyoC
GVx4WIsjizmokP3qy+SrpqUEzPEm6OL2HMmbPeVRvDupbzwx8yWLLGwv1b6vdtZQ
6bpmBfXO+adqHqJR+YQYsuP5lI7K1b+afhffc3nIwLfwor91wTdoyF+f0FcpwRd0
PaDDq8fb1hgo1TW2xBqiJwpGATO7bA7vnJbODbSL7mIgUVAu+GkfW3OefluTOizZ
3NuhERYq4aVzCyxdAqLSTUzFPJh8FMbrUF7XhViDNisDXh2JIS2rSlhxgQNASAz3
MQbJmnBso/2/bVp//HE+EQlnt9MNy/WMMf9TckFkBcII0R6C8prSaBokGs3kCzaB
rMoMuhGS5ur7POL3tAUWeGH2GaFpaaAkDFlwG23PpgPdnbsaKw1bC5YuT59jY4bo
GK1cMx13qzCH2GEqRCbDZO6BjOpn9EiwLQ+Fq6i6hBW+C4De/KDrFrNZkFhZhaPZ
umuBL9j1a6tzJap5ZZMkoXQyzgPGW6GH2PXcpx3/TJ89idAiFo1KpWBNHHSABuCO
NxcAVXgYpVLoCOyd3cg9BySiZCmCnfNwqmzBfqCzQeZ0N100PMzLKB0RRMQ4nlRd
H9B3+ieKmKUpLWmf3N3RTMaqgV0Zb4xTKAkzifQ806/RUU4Q2wEZ+R5p1I6w/RzX
7ai0FTZ/eOMuJIH+zQ3Ac6Sv73dFenn2JCZUt8vmYtz3zfdPw0r+MXpeUo4pCU2f
QUQdy9mMUTfX9+X6uRyE4YrzaqmnBNeu3pACdEKXXiomrfeuXKeSOWkpAeft1ADP
5t4109rrglAxCVZaYifS2LZ0DNEkOm++5CchHNhGWMqnEF2BDSaWfZ1G17CG3DUX
GdQVq+YDQJSbnkQl97EFYp7av4D8OX7/XVIdw5Ff5KbNFVokJKXxl/oDp7ODpPnS
CJpk/kScYwNAIkGWKYdE11JZCfn2wLUkvCGzfic5TLL4xy8VmKvdEgIoJhNzPQ7X
e8vMoI91LUJTXi+HAGKHnDcSWpN7eVlMOY26LZ7REZsIuvB8VxFWOlNRuRbvKYna
YU+9bQJAZ3cnNoN6fpkuaeZyPYy8UAKzZoG7R1uLNszqRF75ybRx1cvb5hKTb65D
9BSSGI4d9ve0mYJe+nuytzqBh3JJT3/FD9uyBvh7bUigmEwKD1yaBO1/9tRFdlxA
jSX4rVXimQHF5K+Qy8DzD/Oj/DF3ihMOoCEuXSgyYgIjX+PWbgN+kAQwdEfwh6yf
CNNQvqln+IpFjzMsT3ECJUvbvXjG+7FknuZJML7KBzx7vjf+FIt7D4KCxWUABClh
75jtciEnNgJukhRPn844JOGF7sOvJQy9SZo6Xq7MEEuiQYT2k6SEUm70iQqZf+Wz
LbCvCynQkVY6xqz9Io2eLMDqDSDn0DwQCu6evsw3C9ai8xFHk1p2mFmXwApefncI
uHyOrWeoHI4mpyWGFPv7zUrl2vr+Pe7vtEzSV5nrhdUPSO3iMSSzNz3b59ERR7si
1JBS+pnUwcZDYh+vu0o/ls4hXA7+Z2gaaY4MWAiXwJXL1K/d50KGYycfjBVROANL
ykzS74v4XzDhrsbI+KyJ6v1V6tUBpwB/sOuq/LiVAoOzoj5Yo0/alx9lpSO9xIZr
gkA8Fjfw0D8kdTHT2SqD1/vwrBFEKTvSPP4om5LkbrXpnjFTobTG8aQ4ycmY6DxL
AGgg19BuZ+6TN3s6scHqzxFK6wTfVRNlopvXhcd4dCP1W5YYTIQIGMRuyoP305yP
F6mdnZ9LMlPWOWD9z0T8+u0QGcmiyx8MYyGKKq47dg1xim87wLguuRAuhOdItqTi
V72iRz+497Z6oBuvcIv6FrPV4pvYi3zia4svtOmk7G4eA1V9lLwGQl2TvMqSNr74
wp4P1O1O1DbOhCOdt9a+wLzRQih0moKqoVaK9EvobPyAdQRcgJqYFKmz7PyOWKFI
U+Zl/UIpxwDFMPoa3gKRCUcydR+UGe2SqU7Iy8en0Kq9Cqfka1Nyw6fqxWACxK6z
cP9IwtrHCukKfPlsXwpdRsYWAvvR1wXdzzk8H8uwD3s53CHJ3/cigWbgCqdNQy4u
qXAXpMw17rgzCZXhVY8Si95shz8yxc2z9860EDLaINoVVrV3SzcVUBWi+4rMqyuu
xzZ7KcThyrdbe1lNCyZtGJyYW4PVTq62AnVZ2+uHz8B0SYbmAkxyBSH0uFTouQD/
60kwsqEr915ht1p1YHnASnGJ/Ph9pU1bMc0K7yK2SQ4zBrmTOWF/XS0OXcu593ED
zFl4ecN4fV90bgRTdKSWlZQ69I/A7fG7n7/4VwTdCyRwtLYXcLFH7wWuS8wxv9xn
pdIvOKWutg57XHp5s1QJLWVF1OHUavHeHTg7GsFEnrWyzwtbT1mPYpYH/rbhMLxe
UlH187cnsSkgSWYlReMJuV4CogrcAXc6YCje6RV5crQ65ZO8h/evxHFKBZ82ospS
j/ivx7YoOrqpb+rLt0+B4lMF9yV7AQleYZKg+p455QYmwwjf7CJn76EtW4DY6h4o
PM0uMq0Xu5qeKf3R/qzb1tbFEFAjXIDsiabbP2LRqUdFkbXDrrsR1E5uQswCJr4p
iDecne3ieHPXok9ON8p3oQAGsTU0XBhIxO3FRd95YBmiTLCJA8XbEauv+A5uweNX
2lOmOqtWZZyOOFHg2EPvCJKLvWwC2IY0wiJ60b/LtFwbvF4MasK3oGBjrpn6wFrM
MUDKtUXoDh/TXZbODNJ6Xg3WB5+EyWjFr0gbjfaqwu/+n4IrkSnJIQNPECMVzkBt
KjSxwoonsNqrCaSjt8mufgRJbs7WBOCeK/ajWrNOdUPj1Z7LY40Ut5dnvK0Bm+5S
YdvTL/zn65+b2T3MMjQwqllxJL0MDwJcQYetCP3PxikvFNpy07o9oEjZRDAFqmts
pQIEIJWLZ6q4oeX3SljynDGR5nVJoKaapGVeSkQARTjXbeQrmDNyNlW9xGeg+28Q
tkXDlQTBVAqphlbf7Gfw2BpJc7CxJn8hAa0cGbkDUH+MuTptwOe8DJ5srKZx/O4X
7wV+Y5MdZU23kEWStwHdoiIZSInLV4DoqtpPfV1R5eg1Cg4qyKAFcOHMkkSKNo3S
QdVnq0XPBOH6sx4XNqOSNRjgNKRB29O8D5pxNRkjLOBsKlsdNKA1kpYH1iNPQVo3
GKBvkDlFB6KzZYpflzJEprz12aSEbZ2g1jKb69tezvd1ac2hGPxPFlB6kfyb2gDr
qT5+YuByn887ZtDXHqaPmLfLatrdfKyvz+apY5tpdR93OGj0HJPWVqR1C8wNb13i
qM+1ronl5khYk9R8TdE1LYVR11JBvRyTrH5Uoz1gnljOT98a7FFqvVSFxNJQaLUa
YzW5hDoZ/nWXdTFH9Rssz355FPPhVSefRkjd3EkFcAt378t4B+b5NFl+Au5Gy6Qg
S8uVTqZpcRmL/KUQmSasIZPaElCVXFxx+Ul+DWy0WouRt5CIlbpGvKTDf2DiR3dC
o0xMowXjuV2yg1L+VXRGgds/HBKgzoJyeSFS95/Y9OawyTtEY4nT+JhX12vWj3dE
t5JmC+fANsSUgmshbm4eJLszrYEngZ6lCI1BNVgCPm1zsXk4JvxSMgYBp2eAkcc3
pykmiSBrkb/U1NsTyxKk3CIuxmDi9V3fXCQ/UGWD2j6nGeKTpOGAe4LplGeFcuDv
wkXWSVlxwFWWwFxiBtmFqbUNTZXL6zImimijm4YQCLwACtYayj1WCBuw1limeehi
meiJLsRfRDc5NHDHiHqL08ZdSfuAioD2E2eJYuBbM9OQ1M+4wXdVhH/fo0Ae2Jlz
2qChrilLjv/UolzF2i5pFmPbkwUVufFc2nf63hP/XP4fRa2i4aGImqYDH8UUgaGk
jRnQWOMqE8q56j9IATb2GIKFj3P7S+wTQsTWXrU40G4aVDSbc3c+a/mFOfFl1kwc
QlpiVwAMkFhHPBM+zVlXPf8FcT26car1K2DMz9AXDh6jkLZtFDXI1AShE3zDmIKx
MecP2GsbXOc3mJmWXgmPuRAZRoVoY11M9FBkwcXHupB4BoEcdD1FPqgHhhSERBxo
Mji+YNV6EhzLq3OEbms5I+tS/aDE76cwhfmc1pVl3YZtJEaYM0Hf3VsGUOQW8KGs
QwBCBj1lokv5kqT/FcQhTXhdBxUiVQxhzdqlJy1pigQIOJ11dMaiTeLtb/yQg8By
hBYwAWWyNYrqyjT4saO74E7lq7RnlPLtK+cS1swSd/lg3wGCK4smtKSzhTgSLi6Q
1BihQZvbX+6mRwWqB6R903MQA9neeQABvm6wOJLFbxYsa0J+vGUDJGuFXRrPZUdk
LzaCibkBWJku+hmx16VEW68S6WPaWuyuHpW4r+DFIMr8L8z1YWsbntKgjVcaXT+U
LSkyOM6vdyurmhMVlkHTF5q7Br7j4/iKCuIjpWVMRy4vltIv3KAaWBMTIWnLfOIE
vOsecUFqbRO8NFz89KDOliFtNwjmH3Gr644uQvL+fWJLic9oGFNr76s2pX1tk3iw
gAFxF9dQ2MGU+H20W+gOrTdEoaVBq/f/jdTgI2A3DvUa9xa8awQyPT/dz9e38NC7
XpRj9fl0ayc6FK413ERKIHCL7olkwWu66YrnVliLTr624xUa3RMWPm2P/wX6zv/w
BProRYQCbBpTn3CmGG8kj7Rj1bypiZdT684wUoOmdufjzh7jaSPmpdUTHBVUCoqH
FeQQnHYAeqoA90hkVekLbYh/FTby0eztKUs4ye/CeP6Bt5R9dI5nGrGp+TdaGSBY
9T7RJO1s/yPlRlIVG89Sjwn/SYnpznleVqLFyJLtJZqgSZ+OpQeQdDfweQ3QTrfD
AlHVfi3aYIj2HC2PnJNjkKNBuyTnuX+9voBo7ZsMH6iQ7ujuBWGOtumlMFYuC6Wg
TZgD6cinoip7Gg/kr8OuWYJS0caMrSTS6rSmZ102fjsSHP2WbBLAU9R2gRd8Mui1
2aLH7CLKvZtBcVKIeKwn7IDnpzmg+LdQRtqgajaoGx20+v1uQeB4DNjCtSpAj9gM
PAYuerNqcAlLrA7gAiGqYbOGarSopAsniQxrACqaih0vmWjO04c1alXA7MFIzKAE
M+i3O/F9cIp78OxtMnpdX3M7Ix2SGs83rnOnctX+OhtK+iGkC12gdqn+DvBlYOkg
/7tI92WvTdNkJ5GZWfSHinKQVsHera3/pY+u54swUP1JUtqpF8U8Z3bhpqtczqRj
UTLFLnuNsfGzEzu0tZOzbjU4NG3si8y/1j/bMZJUl+P9Fos9TdnfAiTpqlUTggAr
D0WwybpVo/LBdt8DQcO9uStHMbpQdi3V/IgV+XRniaA3E82WtmNnwlzoG4d46UsO
MWS27TgotsZZPNm7SPmlczxl8urYipcGM70sO/Nkjq2+/nviJPLvKTWMJrbHYXnt
7Au2VsUCayq9QZQuLr3yUlClb8LMTzsuIQZTGakhTCoy8iiULRDjsyfKVBg5tIIE
wBm1RUAPZDphqMfE4WdS/IsfFOTQEp/q5DDPUDNNp2dM86cpIUOK21egTuRTj4GM
HLl5X8wbvIO+BuuGHM0ARQ7z9b8dI9NwLUL80c7R8Gm9h7+p4i6wQqJkANIygDQC
CFCqJb6XBGyHQhsygzje9sVvuyhkESRL2rSDaEil4fGUQcxp3qGbXzlCDKx16Kuv
fke9KdMPSkbYhqGuUtIuOpB0AdST2ZCkU+xBi2I4T2BVxFonSzOEkm7Dj8SeI/cQ
QX/zdim9/ioJo8AHiSsDf9W+2yQGMpWF3NKCO05eSR3p9vLXmNrjg6AW+6EAOVUt
t+lU992lgSxZ9YyVZNr1ansXY0XNjIh+j82tqCWXqAK+xfZYS1Y5JYNUiwIIVz2x
vQDzEvRH8pmG4aYrKcFwyZROwJ+d9j+U2gK58uwK+k5uWsuOUp268/NjdLUx75/K
1FyBABqDYQ2RojH7F1Dn6qB6X2nGwPYZFx1k/WNoS0dY4D1SdBITXM5BcmH9sHQZ
YG6tkOsf88hOUtJmKsSnYNpUsodHi0A4ET18yozvD4qBAbomsn0Cattj2QzfqpR0
Gb5fM5Ev/is0t+T2MTfbnjJQaUdFrQLfDVGGqyezVrgj7nvj7tCevXQiXelFuGJM
UY0M8LWWzYT3to7R6BbcDPSVrzFN4J94YXYN2Yr9bKJg43WRmzGu5UFKnSl6DE7f
z3WYVNMRPBoRgdh2/2tjJtLoHkGuH3EC4J7AtIitm5ZzGPFdbixv1m78zvPvytJs
vbTtkYTROjct687VgtbtJ1/Dj2qLcnkSsSQLKoKNWz+xkRQ8eHLOamvg89tlo/6Q
sERlyNZFnF5bDyq1o+Pl3tMjl9s06n++hwHjEud5/LTTxBoyCj2qEGz1kfp608/N
IU7NVEiCTGP5N6ZOBbDS7Rz8VNdQFnK1D4OTDgu7sppEs/lcovZ7XtczoBPwLafP
4vYmOaPEl6iEouPlu3IjP5lwkx2PaBg0oRptqSlALVBJoXcIK5gV3ZpMhJqif/KH
5xnSl1R+fvd/s2FkNQ33Ho7ZLUOqhzJVdR1bhfMmKeAyu2LdCF3LMNs8heKWQEO/
NAqEuct6rZv54iqEgmyRT5Unj/1xXmJgCiRkpDui+bgSabBTt5D+0z1KFe677H07
tpmX4Sty/IWqEtPYMdf9KVhxCzMhZJqZoqN9rlp+Va8nZmfdgwCR+OAoZA64R1hh
Sg0MNrJvB+f5LGoZGOPZK+nzAk0mRvTvWeS1Ck/35O9UqBDSK0DbrrmbmmDS2op7
ntGCkgnZgWqpmYHRPCeByzIazXdkCQgOJjjJ7VZWwZCMXg2SOr4oU+zTCmRgqH+4
OkOHuycG701rV2V7jyTrlojjnO/NX7oxjaqcDigSeLKeOiSDBBAmguzpz38d+AqG
p4wF2mV1SX5VXmjYkt6u7h/eW0IHI4r40tKBsxKDcfZI4h+sbm3FeJFVqvgVa2eV
vmJd3WyQmpTvnXtPQ3GlU1fvm0V9m06tBmfSvcOvu2dZPiKEvzevh9NmUJgPKDiz
ocruBkq6mnOZnjeUKLfwdTgp0P4chnRE4ylSuMgWhEVkewwLYievgzW6j5eB8iFn
hqt5LH9Kvkx6btgTFCRlTcutrvM7KGPMRMC6yb223TPf0leypJRuNjYojn+tHRIJ
KGWR0cT3l3TXbkOonFXPSm41Cw/m1EJCAXFDgjlEaAe6es6+dXXi//HOmbf9zoGn
qBKTMWu7aA6mlvrIKItT1yD0OFg+gDM91TNwpdbwWHq0U0VnwaRRy++/vWqtFnwc
P6zH5IXwt0GYPwsS1xgFSfMbqiztOE/J6C/q+1DanBEiCKokmloUqqksOKxEVA/j
QN4FhsbtAUOarIYwMgSvEVDnH4LEySmFNeoeJTpJ8hPQLrn76jIyTLJmyK5E7kWM
NB4FaZWuzbS5Gc1853xOciyuzv576KPWsGh/vqeWYpxB7rXKRffuhqXdWm0Zs0tC
ThFbfwCEgFNPN0PSOCubFsExPP1LtC7lqsr6fMJ42azk61gy+FsY8o9ZKVYAc2ak
BUz4qgGYg4zNwmNvmBzuRNZRdiIXb0T03QjnE2NmnilYYJP7xe57xaAnGtthwMga
o8GW7YCAe2ARkITSTu9TIQyoCen6GsmUGNYJXpTeKYKEu12MWAZlCrkXdq+uo3QR
N7KIDkfpI2izIHW2jEb8T/L8FC3jzh3hweOt1izNdeDozpANmTsz4k8e+9FZ25kz
MLeFJ3wVQcBrZIQRBw1mvtLvOgKhLzW1glDsFoZX4UJ0Nqhdcx6SZcg+9W4qaoNi
CfvPHP6rFC0ke257UiaiJITYgN/sDtG61ftcWWqt3rgs9yFmkSfw4Wv6MiabPSX2
6zTwZS0C5blQk6QwE8X0Ve78hiO6Zmxk36ECCe5n3cghNL2wMY54U0sE+R/f+2dF
hzulbMJZW44CduhvIjnnYcNQjeIjYsVRnuVWjNTalbj2XXv1DmiEcRJZtKvpoLTZ
6w7mJBxrYJxvPPI2QjVjoSNmv0ESoEyDCuoluodFa+nlRwi5VXhUuJSRoTDAji1Z
bnl5hNWFg9W3NYklvGTXk47F3LV43GJ89GjA44yWxg3JC1SFvW5bT4MzrF6UVLuk
LwJPWKvT8mgPK7LfliW1nQz0pPy2iZR4iTyUxH/7gget9hVpQT0oVripv5gJ4Zao
SfvReR4FY+Zog5Oz5BjfCh4RRUKoZKJebvykNAQRdtQsHdFVl/V1Z3jGgpdlGq9z
XN5YM1puLmRXFg8rePx0ZYLPMVqi8Vz+I9pMIkUte5mMvQmV473w8Toh6ozcgKze
u0NF0xywv5ytJymarbwxBLK45Y/PrN1gVS/saqQKNwkXq+HS7ZGI3YDoTWB5fgXh
FNtJC5bWzIyYsYjepxmIphaaQ0EH6cJjySb2cNP9w3vgWG1mWAGN9t/NSaE39AiR
D0hpFh8g/0TUdE4bEG+bO/tCsQw4tDy0Hfn5QD7xSrTZZqUeGW+YQErcyPtqp8Tr
DlrWcAA1k40PB9PpycoA0r2HkcKZJGbH+SL3pKpfeRWoeBmBnXu8tM2kdZOyelcU
va1s5bBxJNYDI/LEHgmtmtggRgcUYWHrCdVVeRZk2MDsrC8GINy9gdlya9yFNezD
LuD41nPl6BPF8od2gTqXXq1EnMFvIFMA6J/AqU+xTDI06PZLLQg8ep2nmSntttNN
Xx09klZLn8v1Da4dBceHM+iz0I4G0GcPQL8GRMoJZs4YoHsiR1R2j+6Chnopc1yz
3k0C0s1O+PrY3rWwjGmC+2fHRVaBsEpCM7EKXcKeh8zG/d75l7EhS4wphfmz8wyo
IFujaSVV+/dAT5F+WB7b43sUIvzPCu8c/2K82BVqJ8xOmFYPm5mo/2Ns9y0rrfSh
F0A3OdkTqL9PjJU7CsjWeUrGqxqIRRvWOHj5zg3HtZb2ibugUPtQ7KuRQV4VdLam
1Pa+t/ijvizKfRTSuUUIUFeQxuf4azTAIhxsbwm7ubxrkTCE8Xj8FuBjvKUbSrI6
/cs0TzofAbwq/XBDmO0527hEQw/zU7LM701cXeQLyDLyKDFlBakWaHJfl1FlgxWb
qqpzZTrzVF4LX04iCHtmrNeyyhENZKvkINoAjyMr8DQ404eQwjEhHzkg7m8GQGmU
6OoJoEvm2gNT3ZiZdAu8S8g7KO/Q9hD/AbcpwNjUMS3MBwKu5DYBBbcmfE7/5tAb
Dp0VnAqE4EqMKysigJiJ9zlJi6WFCfFPZaU1fk04Z0sp0e6oht0r+MByL1iYkNZX
BT6ZxG23/w9LJA7vb7XyfQ6dIzKzu6s/pBYRQkIxxzVMY9WJ+V1Zyx43npr67zV1
IyzDrFPDXu7+hBJyu3YvzFWseK7UX+K86xqvE9q27auvZxFRTeA1fsRKKwRu2Reb
qBA7bAOf9cTGYSOkQFnMVIGNwtfxkzNSb1np5BYB6iVBGLmPbJvrQBE2dbTJbdjg
fO2KYtoBrkSB8wAhz2Sr4At0Dqk/nVR/mPWmSWEzMPuLZfZEDzlVLKpaINxJc1DZ
1+icGAPcNQOzJewLv5fhVEGQ0jj1TIhWLjLbxPP3NRSl7+KYxqbtazNIQ/ySkSQM
z0shVrdcqeBr0GkM5IEphZAS8vHmJFwDfhFlyIgVhdbr/MdAU1twyzFWp67mVtJx
XYb5rcw2ojflWFnXdqAJ/kUKVg5A7FIC/u5wAPt93nRuxfpxbkEwFoXQ/l35JsJ8
NgqYI8yD39ak8Sz7ozlcTjYmiP7gdONrC0Y3tKj6d8iToFQHPx9hi/l811bwrW7X
3QwAO5zXWLamKPdqj34xbbk/OGJTidOnw7o4QFfVHHrUngwfJG3Mq2YNnmIeHTLH
Dty2Ti36auLvivY+9J/axBHTMxfaKZy8BsrzHNN9Qbtk06icFTpSHpD+7TvYfT/A
D29vcx4nW7t0/lSln3lWQY2Mt7uJ9NP2Bkvs4cDGNPQ32d5MPvF/f8ZmwJr74yMX
Fr0QHXbqDZoyeQo3eJaCRTZ8MSzx1bxG7/DgIwyYerDnMDP/OBthFv4Wj3G3i0yV
EsNYzYfMxLDFPEloMUjk+N0P46CHgeGODq5qEoShFRUeo/pKemxMTnZnNit+WzCU
11dHmkKCy38BkRyLNvuImPBxUUZGc1qRMkzYTEemNM0qKNptST4gApJ21MDToDx/
meBFM4PriATRyYTi8PfswOwwmDvSKGuvhis8loaM/+xMQarnH/QfUSYLml8CVUmY
Q2hrsSrQhgt/wuLv1Qx4KZeSA2ejlhIGgmSJqTcNnrRJZWqOd/TmtOd8wh0z7gfV
D5LyxN12fhHTjiCL69lXvvhabx6VpyBYgSn1qFWOak4JMwNN3oo+qHntQmzGWY0O
Pe0PRZTq516s2TaNAT670M1EfoDpDTv3mfe5uleEVAR58j+BGDpRGcOGC9QhpWQT
cqCoS4rP9cBzITqr5DFzxP84+KmavlRXH04wWg7Y5VLveO4t5jxhtZZg/wPAxbQr
WGJ+PSoNialYYze7e9d1xZza/nsEFfVkbSHzuLik2H1diyRRSEJBUV32o+v+de51
1DQDlmjdwkB+xc14k0xxdzT/LgH2eP0SrZOTfpz5sU/T3imENMoMRU86kB+nrd4U
eWjMMpMXhgDZ+ydC/XR7PYvEYeDqjZ5oMego4RKOHCxEy5XCLNEi59z4/ssU3ffk
yQwqOLSAcelGwguZeiygX0cUmRQh0+6svfkmqrz/ZKlDzPvukIesdvA45ko0X+OA
+09Urlvrs1fzzUc+FwL4RgAIros9bi3K7EIQP87yseorlrKRFtYs2aSbqmMukIrc
ZTzojlRC7GLNSKK2RQdSmoI9Bot0ygPHsGp6KGgQTSDEIgPIRKF5NJDmQ6sO5jBu
wBworouLscYnuuZoeqTojWdJQ6i/Qy6KiRYlM9NKJec9aDylDacc7LBBJaXJqdo0
UwSTOEjqc3CWNjhyqwjhOLJ8+KbZvEWx0bvldqUgk87hTtWEwwzIxP1+qlCU9Kt9
napV3gKBzgpChWdb4oWb1PLIhJ6dQyc5VM3WT2/YHJY8mACrQArCQoQWRObuD3gJ
sls3kIcORQyK0YgZ9XEI6Es40IZsbUSHP0s8GUBcegUAG8/VX9dqhCdrubUNLBNM
SpqBsMkCk3yJlWxR7Peh5k/dXqW2aGUPlEnwAgSNDrBTC3iApPJPBei6NyEWiZjk
4Rg3l4zJBOePzUmS++dXwyWcjpp3wpH34dSbM23WsSSD9Uc6Qm0CiYvWfnPlH2gy
ZxgYak6fip3B0L2bflUUuNwNQYshtWoHvCX+2W1DyhwfQpjgRKMhT9AU/5y2KkPo
z32L58w6KqOn8zkv6n7IOS50CpIifFJfe3WdoeUTR+WGiSumOeYl01W3qdBRau6q
yQHM8auozFrh6WQ6ABd+c+Lp5VGohouCy3m2HuE3dvmkzAHn7J4jzFaBWtqHAU0s
zxcNYcgVWwIFTCinGawXkqwga8zGPYb9alAIZxOGP2T8+4RTXS7bLAdw60QTtsZM
eKL/DU3a9VwVzi/jhaq5DaRI48DPZp0VabmUFALpgs9+viNjMic1PgBcnXJL2aIr
Lkig27imEGDAHLf/BQQdhREiSIrPhvpPDOKzOVVukgEqrCHDAMUilo7imUr+KJCp
o0iI8Qi+6XNjxurD88bTtGP0Qj6UNCAb9aIEpbYy5p9b7EbPMviA6v7BlIbl7YQo
Wq5at5+sJf2/Bxu7Sc2J/nmCyKv/MY60Zif0vy/sSBVX9GzS5AdenPZXogJSU+qs
nOhGYviKotaQ4eagSHxhEg77MhzYaMKOmZTtswv0TVaTjXouTV1SryZigXUjF/+/
OULkKX+hEic4UPA28jYizd7C/2swMGmYiCcARPMIQ/ZCFiRyMGgKlQGEwNJISMc5
QXpHrXGposPFsG7QBmWKwG49fZ1z6en9H5gTUH/MCWKU3eU+81HFXjwzJDbgkFHT
zHhPU7OUFMq1FhnomJd2fRZuosjLEoEtH4432V1ncxMYAPClLevueTH6ztcbaZd2
GccJmjjAGmA2kOOLXnMi/1vvK7aG51RdG5nSsAIF+NlCvL4HQTDlUQsRWHDv0xKc
VG8O1gn99xAY/zqVtUI8stRR4743rajrnu4CabtRK81k8tqzcrDUlK5p6/KAjNRW
x/zP7Hmlp9wrOc6Tv5EvwI7V3zCOPZZZPV4VtfQdctnDNywRcGSdmBDSbhUu5jRj
awjXMWSpYdcwAnAQAt2gyRKnAJizIYJ/XQ9npQE2BV7j+pj1I0odnPahQu3fzib+
rMXr5Oeyjok8PHjTWWViPWwqq5IMlHHdEtKfCNUDTwAor4nCVim9jGfWTeiaXkbg
CEjW3LMQd7u8UZxRwuVwXajFfgZN8YhhgH9ZW3Faq4t5H7b1zGmCG5qF4fqVonHE
uySsBLFM7NJGDYU5JEsmvY6jbB6G7bO4zU8/w27+PTA3uHoXhqcZjZrL/ShFD1FZ
xOVT/Ut6iPnwUWEfWVrY2vWlldsGX/ipFhYYCNaanfG5tjpjKfByF01aYgBS8N1c
EcBvoiR4bmCmB1uRYmuMnFUQdt2q9lEJxWRMNemCnbpPGMsqfFWLT4xMLFgo9h7C
6EuR0I7auTanfQRIV04qi/1moCvwcSDZm9A8tZ2rl/YEDoclJ3r6m4Y6mGw0kIRN
aleL3RxeAUgWYgiCUuqc+H9fQQ2gArx8y5Hv+NRxzb0GB6WMpuQMagDZ2rAe6L/5
8PIX/o4aQu8sdrYKeNJx1UFhqBS2iL7x+KIodCrRMoGn3dIrPZtOnecnXKmQfSvO
uTs0xcvXsSrwCNwEUzpzd0ZaZ2rT58qWqGDTpeurbKmJ9M5nKkVN7oJHvOAue3ey
NQhLQK4UcovbuIk+GhIN1ULB3cVXGiZ8bhIHr/fZRX4EGRGK93AGxsUaRkoYqHYp
ATWNukPvQ7v3AB3L6WFCj90XqfRf23WNycndWN+D+rFWMFOJSHgP3zJ+RKJvds9S
kLrMThioUJSus43ssLskVeLq4YKPJy9ZpDuW2XRnxqOgg3sBuZJh2nplzsz5wPNa
un/5aiqknTE/7yCABBQlQjs4zCAgOW+7KnVIItnPe4GS+MGy3wWRTD31T6oCTMAK
GzjjeL9P8flTY0so+UCAoUojWj53/dW/EQbee3AqtuaqgY9GiL0cRUb6nxxXc+RU
j2NqpsaAYEBNR5LHOyT5uI88tQ6kjclECP4E1XKiI66i5lte3IcMF1EoSPAjOATQ
njzSmMa5owck3/BGVERcDNDnsAExwonc29HQ3m1H9bxQfQOUBaGV8ll7dbhK9NKL
Kbye/7Vfp3hluZAL2uABVscR7keG/+Ume8piL94i/JMVtE4Q/NntGwyeCwBBvmxP
TezgwuVSidXIoTqnpsEjFQqnvN8Z0zzx9LOaVYYpF6GZdLshMh+fQwo77d3YhOFl
kH3qi6YOemb2ai6u2O2ymztPMu+sK2UShOiCh6ep3DM0Fnml8c0axV/XSwwafwdX
fueZl3aX12esqtVK+Km8RuiGZ+7nozbbaomlfz0w7+8k9I7qLYI1vFwvD85HBLqW
N4L2s6ICagq3zDL+xmZ77DdS0s1/F0J8wqfonyGO8ruYBYKf0h8qWm2NDaYzbeJM
6m9Y/Jd9MeUdFwvBvUYxLKJrnR1lpq/9caFc8lBhM71LFJhwkf95QYee8RZj/yOz
b+vNUb4ZwljX6c4KTRB2RlaDryOF8Dgip6zCkeWqWxK6yj2RdARXq4V4ezb9/WwC
2ddD5gZWIzsw1/Swuc2kKWOKRLcEYWl5vv4Sx6D32YwyEGasG8cED3cL3dxjgI3F
4z5I4ni5AdGVllrZ/ynoMqGlRJ8ItohCns88rGEWASslxizoSCwig1Uc0AKeFOY4
689LwXCDhoYny95gP01V1+Q921DgHZnijH37kkP4Vv1YuFlDpNecqJAo5jZHgQ6O
r38UQyUL0WZwmIScSzdCyYTHxqutr7MqLOGKoqld5iTOaqsIYY+jgVOmRREb0+9G
GOaWaoSQibbEB7k/CqckIDakdjXxjkW5g9FByvEQq1brsh7WP1x8giLKOIHbkfQ9
vSGmU9jKTf+gGj/PdHFYGiFmT54XdKKFcs2o/vj5+4TQ7Qi12NiMmiZW1oKPyNnx
49ZiNEU9Uuuf+3UMH+Dos/EqcPJfysApU8naI6rUJOA/T2Nfu4BvT1hjqFzXIvaf
xwxcoaZC9QN9KzycoKnvoSTHaQdebHSQYFw1kkqSDTXFvzDP6tXmVP40jmFzZjxy
fyWU0JshemqUcgY9DG9WWQlbjhejSw7+79Z8JwpgsRh1Xru/Qf2z6LyhPQIpvA+j
LpbKjrQfjICobIXfFjWdswtixNp7n6u/bw5TtqeYOqxnkNy+1rdsJQFLwf0JGexw
/OqsLi1+iQaKm8d7L4Z5z3WzvhDLmA2erS2gDGC/XFP8/LMqQc82sm1kLj2pQQwJ
GBZJjg4PJOnHrqpP3wlnrv6JokaBxSmShztr1PQPP49e5B+w2wfBZVIW+V09FUB7
rhRJDfkYLncLs9Smmsxrgk4qe5mcKRi81eX3+9pwN3y0F+XFXQFGRVrJP1rBU5Ys
1JaXtxLdN3TNkAgCkVq0nxPRQjLoFPpNoECeedzK1nfFrUBszTPnbVPpY/9dFuYN
bx8Py1dX/BvFb3lI2T+1bohgqztNlaa6oMm9L+x4aXrQMjYyiv7dNjDkLQQeL3eu
NuAZo9U+LM1vXRWPdbRhkgd4GwFxoqgxFmC1zF84OrBhzXNklDklQKTaJDyAXCW/
HP/vLqi3i+SFcl3wcDTp1nSR3X/b1EH4cZ874AYsDpYVHkCOmho7b8ipd/OunWKz
lgEdqFnhvSfIKgCUDS8MxiNh2Yu+P1AmdX6bjezUhxyFQXxF1TDV0ggEPXnP0ZPX
iqJ/iwGCFTtez9I9mL0ckgx4FaZqJhfjJvqAdEJ32S2Cg03H9gSrf9UZeydHzWpN
o12eaeeZIhBNvQ9GCt/LWwxPgR3Jtw3MzGLqaw1JTBwma4gGva+pAdSwl4IHlACr
9wBADET5Dwzen3QcOlitbmqeojhJGR1/6eRbBONgEyjGdsbm2w6BjN0MUNG1QrK0
W/WuLQ/+K9/b068DflVHpsulIsfHhLbl/6zSu7hSQPv1gzSFA9ABIr9KvSw2gQwm
n1l0lUrXNTUaW9YMLQfs5B5GMb+txsaxhZV1XHcbRXx89AIlx9Sr0xFGEuOvUfER
aw+LOjawURKHUx979O5/iaZNsSxtz/67EVji32RPOtyxQyzdqnEoS6mRgPnwYUO/
yRitSBFt2IR5NsVW6DoF4AC4aPqnzQoM+sTISEKVyQRWKOfCvTHf4EKOosBfl8Sg
1SzNJ4DmqdrtXCZGXQ7ExGVskOpi0wj9ffe48X8v/k70E62V/CW7cSaT4gQkbDU5
tu+LWSPKf3vBpoomCIh0c0DNGBdN9D7jRYoz/+WXv+tAkB2dW830MO5V2HVtLaQx
6geJAcCMbgsk6yL3EQ9s3xbcMYL2fwpJVuMRPqnJkfDci4aw/kdPnIrKTsLzrrHf
AeFpMaa1ZhpayDrJnnkMJcQEYw+94MeCyeeeeAtmSPtNgeNKnHQRl5PbalPQMfsT
1y9Lf5JHPfm3WluHI0+Mz60MfEiZ9hN2jekyETfQ0ngcsXB4QP4naNKS46/zaS2V
lsl+AJnVslTM506n4CMtId/MY4cV6RGAapanLsAF/nmVAatkymFwfvomE0WeuM3e
zkbj93aN1QS5mT80Hh4z8TLVK1Rq08KJLOs2EUPE4mhQkg/ZXFOixhH3W4NR3Af6
vrQXx+kpz94nk2utMX3LaVNVJheujsCON2+IDyeL/ScJdHG/MXyhsVrTleC5IESM
2KpDfNhAALfDXDX9+3H7F22DSU1enYelpmJVtawkn3SClyG5kH4CA3+Suh0DzDzZ
+IT0GB184EC9lBOKynpqXsuIIcY4ZDAfHn8E7UqkqtHOPfn0E1L2dOVmzrmmyQ7c
nxos9eyiHLDJ5aDdolGaFGmfNSaEKL1H0qZdijZI+D8m/9gyBMDzfajkqhjoRzn7
k4hrpVRHABEXJPnHiQQnsLu8Yf0kUQcau6PcDDFdvevEADEALfmmJ9R/EMfQRzWA
t/mvnxpm2/hSLdTZh9FVHOL4//fM8XiW1u4chYRdyh896xLBhwkx4menPM4uCuEu
N3n1Rc6r193h9dXmX2+uYqlr9OmQ7BFDC8Ilb+wMtGujEiPCiReiadZLyVbCa6Ka
1zzpGK7Q+N3MtDP6qtvBzq+KS3xA2SusaUoXNvUB1ODMUJ3mYrtVjWSZUdNELv5t
8/pmIGRYNhv3OUmIznYm+0Z3eI0/0FoZkLEIDq+hBZ1vasfVUfP4KT8QtG3A2ag8
FK8PDEo/87EoLY30TN32N0MS5YwJBdAQJVN+fiOUvA6zPQ3wO5XMaJ5Bf6Bui4Ly
9xzEwERbaonhQFexkT49B6tirH7/Zodo/2+O+rzyBhakq7mqh9KTfaJJgAgZShu+
brR9NR9IrUOeDvBMlZiUcyTjWiB0gENEe2Q719WpnKN+qz/XjsreyGXGsKHzaObF
Yvsqv0XJ/Vyu6T+SG+AiOP0h2BbJcGeZjPEhNRmJZRB77i01tCZvpF8JbyrIBmic
KoiQoC/pDmkMA11lf9mzlF5375noYtQngh1uDQ1HHuKjc4c3Fib8wkzZGVfvr8XI
plaqgINAWUvINjTCw0t8q2cTVEfRdKhC8wRyzPk+1nAiJ2sdSzNyYcer7/699q4j
X0H+3vM+2xhCNJU4RQ8JPkONYfvVFnxb3OMw3+XiISqSQIXCni2ASVRNCg9nZdQV
xMFsHn1Sbdqm1ibU12mJIypdeXd0dK24jq66XMxka4PtWvcKU3QddrsK/iK4ZF9h
Pbf4GWC9KKeXhozUYhfkeOccjTyhWlexM8Wypy+bafvR/Ujm8gs1t2+q7EY5hBLe
rGgL46++BCynvLgnqfF0cNSAhyNwXkhAMTAy9AWP3jRtPRVMaanBDGTX3QQsZgWy
osXP5F6b+gbwo63CI/KzN67bwrn6pX6LGkdfEs2CYDjin4YW5HZmTlrl1a8XZpnu
GQsfS9gMs1/3R3IQUN4XGIdkssehEMXdgTOcNMas0qMNKjSIaAezCUp+3Z6Yv7HP
inLkcAcuk9/k+WBYj7QA2RLXmIDMALQD1zP8kxiqnCF9sddT8CHgDQ9ZiTZYVNhK
B31wZtuBXgFgMJ6w806y5LidkAk6G4o5PdiHlis8Prjl/ejM4GEtTP0cnr1snr2C
giAItGxZH1BhjnlhpedoKClDwd1mx3OjhY9Y9JnOetlOyGU6HFK/hjl+ZFZVStqQ
bLkTsE6A9kzSqYvhr62YJ8xSufsci9+XgJv+mlm5pA3b8AFC/MAL0PrjBmVZHksL
AeIggShec0jdTeoeJ3U85sbdH7n9wWxg+/jarxpbhVr2vfm0VQZfDpKbeaS7XpWX
6zCiUIPNEUIE9UnkNQrZpRX5B3ZpHySY9qMYFDQsdF41MhBrkXG+/j6Db+VsVr/q
CBmdt9oOVFrM3wv+bRpbR5jKuPs8+fjrhjFkRmXBP6mQPDf2GBw3hcp/mOk1Jdis
yjnz/z36YxKyPu9fEl+EM4xBmmI8bXYqljl2CFVyFGlTpjOHG+7cKqk7/3tRlsyc
Zxhg49hVDl0f5tr1JY8vhGNV1XtngJo+OmfTJVgfvQKtz3+qmrh5mooG82ZL2M9L
zzX21CDPp3IcJlcevtJKX7K6wIneb1ixeOx/OP+RP2JWiea65dmNoobdrPUV/HlW
XFRyXO2JcVrloEUDYwEuPpnfU0nNTWPk+nkC/ixCTU6tFlSzmCkMS1hI5ke1wG2q
ck5RWLjL91G0aPA5Fk0v0OaFSre+mFButPOUKn9zwWnT9KAgLWvAntTO6RfQiFgR
bc5jQdtpT+egHN+HxARS57ZnTZ7S9oPalfyXVNJRO4pWrthkztr0vEFKFrjRlAy0
2gzMdrO+cQynSquqy8Hy3nkxrOeGt6RF5+lTihOU6t6XrQEXD7JWVfcdybAqQDQi
mWcyCexsvPuYIvH/icRtaNWDNstYJdrO6kXpx9Z5Idl49bTlmxUYQKAl8wGvz08C
fsd00lak+WAF/XQ/ukFCTHq3Y8ROU6aOQ1eyA/U1vN3yesScpvKTVsOmsJ3fU7bZ
3IAsdN3Nw7AxsuBcmcrON5FyC5KJFWw2zDM+MjxSPl+jJy1ehGfESKUUq3NiOeeW
Dvn9Ur6UFauDFooYlZLWVQiGiGuzDOH7SWPXldvizqd37pJfXtHMi9InaSLel48F
FTAhg9MMZzzMFH652N//sk9Lqs+xYJq2pVzjJgctWq5nWIlhpmikWImCr4jc5Q/8
k0RdDUKSJWWQ3XBLqK71AXgP4qVLvoppP3tzN03dvMaL583nzMWO5ZNTKe1alADR
GhdrBCLROK4lklFBJlB8RD6+J5RoNuV8zfHIf9hzlwlVAUL1lBIvBZdgLoq8cOvG
ERxb7uGFKlQLI8zEQ7wG4p/HlGzfvDOp9fUP33gkCGaOVcs7SesDlPgwFtiy4KIN
yi09JEJFq9yn+h660CMY+k09dprfiV7YP9yYV7SBHmGw3hjYsOQRi00eSpOIaeRs
2nRrAxl11bD+NsYN0apdcmofvKxkvneiLFBaZqfjgbqwO0bVvrG5SozWmSKXKayI
MiaiKrs8WOqKZ8Vc9ZftR560YMLlqZ0XsAOl82C3mzjnQZQS5HXq/5ysifckJhL/
2iIeXAnwylmZqifipsiqIOtnxjnhHJj0xGC/jkR+50wmtKQVuMWOnmkngFvdMIg3
u/RvgLUtiNJltrvOVW7bF2Au/Nq+S6zY6dkpb7pfaNyUOybh/S52nC+hftp35KMd
OIYVdy1/+380bRejgasMp2s07nyXJLs5sGtswbcmXyLsqpEGt5BYhwDtuAJjTdKQ
7L7Uws0T1DGWJCE811lfX0/P2DXyIy3xQ4b49aFOtLSm2ui9uiNyrhzXlPWV4C1v
BJGJdMzenOR9//lLoK8EJ+wOD3xzCdjnto8Ri/z4IvxNt7Ruh6zun30rA+LdJ3pJ
F4gTimx7YQ4A3+5JGb0NqGivetbJEZMHJrxwAFjP7sWg2m5udpe6gy7VtIDX7SUM
ZNb/HLeFRr8QehFHGnw/jgBzCFohrCoT50D6M+yWHUyqnNM1Aarl0aZlP/gdVw0J
zJLlsRXj9+RVhit3SQonomhvSDe0Xd13MGFjHm0cMRV4+OXUcqyaFjW8QSAHrm9A
vYP2bfdg7MvF8DSBgnEOyHT+W1NIPbCiXmEwuxgj0Q3EhC/98bLx8gmN85hnJEBu
X1FLKD02bUTBInSOuMf57/EWl+HxslEkXh4gxL2WH+9vNRcIcvD9bwqVeHi2ezBO
3LWLClMRFDUAYRZeSPy5a+V8zlGABrGKCj9WHdPKQSBklKpVjdOtPYE95pGLj8dE
YRlv3f8duWBFjbftHzRYmnBs9EAmN+PUTqXaBxoLMwtjA+/RaXIrIXR3Y+1TXBbc
hQiHPXWJNqsdDXGDJZqs/QCI0UwcbmDZ4I5UOtr/KVb16slXJOUJH/dONMRqgAaN
45ZyoBtx2bauMahg5tAWlbBodLZJ2OAuXfNcFAZdaUET4g1vUydS4Yz46QDfkyBp
8F2hG5mxqb8B2DgZS5b/ayxZKoJ2MIV+BF+ksJi7w5Lg+mYxNqfRxVPsF9raK7Ay
1AbZ7jtBbfE7pAw62wQ+yyhNcwm4AiiEf6JU2KLUHsPnM1bJ4YtsjCdp0eHVqk15
rzVf3SRBof+HCuogBKwGSANI21ZxOCuVCEalREo6yY5gdx+TssX5oIfnH5JHnyCD
gWMsJr93z91Er61xo7CA15hyXgbn9mQ0nJJDqLOweAJynOWKz+iYt1arPkT5BRy2
Bri4diGqwkp53C4Cm6XqZGiVe6PMeZ9KGlIAhKNcQSAyP1ZtydHpfXOwq9XU/6YX
1+eFhxQ4La0tthGQmbtfLsfQDuseI7jWwM3ewwjSHs06Y4r6WTR72Hyp/nj8lTJZ
76xxRnTNGH5pKzqBO8AlJzhVuWDJs4/yPljyaQGtovMupfvzUjF+tLnbq9kkQIiI
CVVdcjom6e36mFPNQUs1CHZx3f0xyWi/SKgPUDVZR10g+UcNurfrnpotWwX44Rvt
3LrOlmCMaScYYHoKllcMH+tG2inx13xc0ipkH4oAUW/4aANA0K7G9B+0Vh1abQLM
Ch5AfStvFK5fqCGXPVPQKzuypDyZA2LIfR9sVxRQOHK1ya7JpXXweAwoOc0aDlqk
1Fg+p5Jb2lVvpC89ZgECnUAXDjeL/MZzYtaSvLeYnzWTS8H0Z1CKd31La31sJQwu
DcXpW7sUwTOG5AGfaa6mncS7Y5rnRyHWQnzB2wY/SZX/zZEtJaQDQ9HGLuUC4Z+C
4Sz6jKGjfmRZsU5EDnc/e2PLzDvrqAEUtQpI9b3hwAQGE15gSuMymWdJIUbafn/B
T4FvdDw0WdEMvT1h3eBlurDacv31fTFtj4P4VWX7FjfSqHki0A2AM5kzAcMTxibG
JO/zP7Id7Padowfee9EBo5uo15+qX/lxJX4cwYlJhdjReOvtdZGEU+Ol2u9awtAJ
J5DoHZvK2A41kPwEg2v0P2C10LJndk70//Uioj95Jmt0is6VomPbEUUSW9bzJYgY
Kmu9yMmLKYDMUsJ7M6x7oYElN1jkiDFZfJytkucmddjDCXOHfExKbRXTW+f5aGBh
M0NOkkgNa0cWvg1KL4y+GupvQXjXdnxc/oZbwTP3mmGjbzQTK+3tr7l6Aymcqe1b
D82KQE8AdxFEB/K0zYEjwFHojsNhTln9KL4A9dU99m8d6UgPuBd4xD+eR1XhrmF5
NlLgJoMUa5UaUgqFyJhi13uAAUjhEjKTARdviBA1qs/Iy/Fic20AN8sgJsDn+r1Q
OYpWUVtTm6p+7WJEy2jMo/PblP9NuAPOlJU36IUSq4r8DEnaOuvdIIHbmKRqwqaN
f+6o9o1/XuzBRUC9GyTD+5pWGSvyorMhytXTET/A2TM9S6UQKRZTgefBZo2PsXp4
mwrIGRApcH58c/UrKMFCLRL4EYn07O9/ha/MAhYKeZnNG/5pBPXvILlK2ytBmspw
0vfq/n0VYshkiuSbAq8Bv6B4Qry4qYwcrDXqm86R8beWp3K1cxn2eQ3hty712I4N
5k9lZ39+xSe9ZIwH9Rj9TjuDzR8bim8ebMX5S2EmD6Ti6UnGxlqM4lh30TE5r8gF
Lg4flYEyFUAVrvHnJ6Tt8qb8km3FgH6Y/Ftoe9TgGEF2v5nBxF3Juxmmrq9SjdF3
rNNz0h16W3kAT4pU1iKehhfD2okAt0l+2XrGieDotGayhZO5ETl1g3h2cDH/a9+o
vFXs4JrBaovzBx1JO8MiXaMaELrrTTWnMO2gG3EvgHr77UJXsduGgusmp7WyF+ip
7UYEEeM57l31uB+6LRAuTCER6V/5d0TLaXQvHfboUycwUMGzrL98rP3KbNzp8c2j
wBkwW5EtnXzc3+5UvwHJMR81j5HBnlFtWyba1wVYhafp4xTC6JQ4tSsdwowUmlrz
Rt1mJpAb2PIt0NQ7irXzXAeDUUQnXL3dIx8U9mg1C/wq8IQJB3/LV+3HyQM1USXd
DiVXcYalWZ1SFqf6IVpuxpe7GVoOOwM2WPAvb3bcFagfvbZQ+XmAu73qNIEzTcrK
r/qe9aDN5ve23TrAzMqFzjtFYVqJ6QDpsNnGXbhmxEs771xzXQXBBQu5melu2/v0
ZcdqJ56Ta2pI2R7hypP0hq6N/VuMcooXusyaOML/4+NFR7z2UQWD7+tp3UN801Qc
tquhhRFT6sGCrJl8O+KzBwUwgNigHGnySrMSfNBymXJ1DY/LUXYgnCMEtw+0ni5o
R9J+CHXg+TQSmfK6Yu4HZ4A/ABrsqDhyXInR3oMkg0pSTaPQTEhbanH+dZ8dzqPa
QwDlTFZIs6qWzyoskIwAMj8dkj4TACt5gpJGuqQLVUWDrmlLcfyZk3xb7o9eVOkg
MaZH6cghPkAaLSZq7Po5OkTOq0NN5UD+Fg5CANMdMNS12A5oAksaIlNRATCqxddE
tItrLKPMhVCNOZLr9HqAdoeFJcgXfmLu9YRCUM61T8o0vsuKuT1dV6Fiem4B+dLi
nDw3W0UVVdjdnmUq8vE5rvmoEG3A7/wbHJPjY1l300shl9IPFWIMSxLAdqNKZCCW
ueQ4T5PhlxFFoucTaPKN4C/EhGVYQ3fC8ya6HtBoQyp6ElPZEooWg4+i8vnuQl2n
eVjJ6I4j1WRCWvBvwlZxbPTZP0Vn8hnLLh5f2Lss3LfA9b0tdZN7FnO7bjalhJbV
TYkpn8kbWzibQ5D5hNdvMXxqaOjVySFajLQyuueGakScNIQ/SIGtcxX/KFhFTKZN
rmWd2fA5+0c3GGu8F8Ph6VJkM39ZNNc2eCLIVZMs1Q9/2U22GnJadQia+QFS59xG
GCLX7Ef6ldzoKEgX4Q0AGBdPNMBNuzyqeOTEBFvTKcxQlRCPn2r3IurewE8a7l8r
oO2fJi3WXR5A2CtW79Hq1Kln0VddK2P/7CiSHv3rnAE013Ds01x+rh5JhXu6blNh
a2ESnpvMmkGZexd/TtWjGdq6SA1FNyz6WJoI5eqYIco3UGXH9I4oAa/mbKmRc2VE
0JNS5IAGsAuy8ppl/gy/2ZCUXQWmokF3J3sBzKaOttKnWw0QdXhkVek+J+aXiCz/
6+04ShMTSbWJOkOmV3UyEwirlrqAWbgtPQXcJLdZWFqZbDgfH7HC54SruTvaYd97
130cDGNlgI4I9vhFvPmu33wqpkDh/eVqSM/ROyQtdrfe1AsFPcx4glRWsgvoe+ue
kEHiTrdyLcj9YDr3ELbRyyWXJKK8vUu+ZtzokzekPvrwjQJWo0U4Laa64C/Iu2Pp
Hzt+2Vnm3q1mFQkMucOhYlsL8Wm8bWfVAs8ASvpH1SfTojaIO/UdyOodc7O93gqf
Ca/daIaAhCgd22Rt99JWD1bcAZzMXLRbcqGPE7s1p1KyMnKQggjMic0WulqBM1VO
TGFpL0UMgLgt3AnBhpsqkpKKKdZxhOKW9RPTEv3eZ4z07YF33M5iTHglTuQDt4G1
N3P8G3vApBZfRfUSnX/4kkObRi7JWD4mRTmZxBP4rYtHk18NYSEtFR7tCbJqVMlo
cMuferN3ywxQwuVRH6rp1LEheYItXEislDkXcIEKi39HVfCPCXeAf9B+Tp5gx9Eo
CHVGObZ/vG3VE3F6Z7oLiNekjl9qvlM7H/n6iw5AfEkMrHNZU6yGV8azIcj09Jid
KaXMrGFx3GfsDJHdEh92mPFvIDUmPhGfvDlXO7pN9Vq8t3w+caq7rCTS9oje7xxY
032PDI//R56xZ3yh4UWJ09Jufz4cnBktG5WPr9XkazwZI33GG0+YWS/cJrg2d/JI
03TdjavCuqnJmLlXXW6DNf9ADRQOXxNK8Y2xgcgWy5L87sBMlPegPimfLTjOCIhS
EX9JCzpe1I2njtfvsCcuNJIJNfsF6aLK2g3/0+Jb1Vb8gPritOsq1RHy+cxsLVon
31xEtlnmwoMWev1R0hWP/C+FkCkP4j0fl+AMfPdXCk18iUyE1+BOGErXAL5ZZU4N
/xfrw/JF17ED84dI1Oz9qzJyPBW/G8g6fIXKjI4/0Z5yUDHr37Jj71Gh4U8RbDr3
sp5hTxveWib2ISDmIdbit0Dty/YLOsrQDd0XNMqe61s34FAUGNMetc3nxCJ+KeMU
87DJiQTE0ctnitQhoXMyhxR9zFJTSFAHwuBN9/EH0u9zXiTmWLVb+DoysZ3EqnW/
JCridsXH2oUTeDR+NA4aaEryr95BUKrsmhpwAoeDT1133fukNlMbe5/BpZ8evk/1
lZuCJ5IB7SMW06HFCfNIv28p5eN5w429NbtFe2XPRflLV75bHKhi3KTPqdAhS0Nz
U91J2oqTvNIOrMxrVxY7XJOj4juYvQJEzbOCGYLG6Pub/aj0PWQEsTL7Grx44H1J
jRJzjJLkO/R208rHC9CdJvtHQIWclCDn0zx5eEeoO4iUupZARak5cTZNjrPut33u
lM4Yjog6E2XbPJdJO5NbnvkUkWckuxgIbSDsC9z4KsrvxDrdtVQDdu5fjas4V16K
QcdJPDJUoEOGdD+GAJ5gpJ1ixVLzlSPS99g1tFR6Y6XsyFI7TgOokaLdl7XTzmoa
kp0MCacPq1x1/xF52riqgmEn8opNJMt2ouUEoIheyDEajuDt86xEnh70k+9lw6mh
vcTNP/lctKxMfBB93nzAyxg/QQSr2VoLP6RyiCRR85LKBMHriv+ftaW1YV+fr+yu
QtfBUdmp7PDbRjAnzKT04BQFfdwRoFKLOj2sGjZfp9sdDQGGjr4fj3uhbyiUT4Kt
flmgRMDGt94ZcDZ/fj571kIHt6u2eYO+GOKYmAhU6+MhkaVcsuGsZMjiIdUsCv5J
oxUSf3+48HwVObRJkSyTbcPg5tYIdjDMDTUjvx4l6peqK+8NAatHs9NDX6HzOxnJ
Zv5691HpvzAjamClHr0TKFSITl8u53Kg14hHl7doSScXRxycR45TdDNSIPW0/b2J
oPoIKQfcn0dnDqWjhDTPt7/OcgeH2obYoyMKHN+J/4NGoEIlwBUfPhtgYB8G9q4o
6HkoOSsSLOZLIOVIfkLgjp9TxQsRZ+GT6Gn7BC36a1c5H/Ge8XNckfEzJrVr2+nm
1eKn2TJRkERgtBSL1C8HpnmXkXhq5Q+38OBGUftKcOF4+cvs6rBtLIlfssOBxD5I
xhjMxIdncrivnvbo13zWJOmFynZiive/ELBXYG2fyOdn55ZGOkWIvOQ3twC3koPt
LXg9ywUpMDAs3BxFLS+3KFfMcQ2bAXhMoMiExuNGeo3R/wPs7m5PVRv0S/0SaNt2
g86c/YDnh7yg2S4534rX/4MiTeMQIDO3EChDS7INwv9DxluOUK847q6K6Pe3vEd5
5Zx4DOy81DnMrPsn9HHNRDmZYxSIVTOJvnEOmidmbvfHCsK/Cx/ykcrQ/OxMinIT
qO6qFhpad6YWjDekPGihpEPW35hSrSMienVx+KzsZmpo5I4BhMN5jnlRosMFby5X
E168hOXkqFMFYNcBt9F+J0J5eV3u3Iwb1rX236QsDkdljihW+LAfeTdn16WdWO4y
gDqdfIMg3xyO7f8TVryd7V+g6je3+McNoj9qRGPJLQ7tUVQpQYERKOKvXXuuAdau
q4bUUjrEqTBQDK9xnayRa1UDdEcaj7pFtZKLj8c9hsWIH5YnvccvkS90A2BFPyYp
4FATey4nx1nTZLhiMpjrj0t4KxSUO+2ceoierqg41SgykjrlQhtRM2ECo7lh9x8f
Y5K07YoqvwwPOvRsg+PRO9Z3qCuI6DtNG72VKrp508Uh2du5NsCcf2NriTaHk8Ht
T2GZRNhFuk1UmBsSNR/gYiFXGQ1rVRkVHIMRbXPm7pWmFfO7Eb5cEp5UNOR+EYqH
Ku3CcVL5o8NZdqnxIss/CEbFkExIqt+a5lEPXSFr4bzwevidcNmmzincQ75uGHPh
rfSCaH/FB4FO0QfrU3sE8OydkOTPvLlMTJtwDn2NXi+PjdrVpy1ROpr8osfxLJ3+
MvO7wA9NFN5aBQ+aBjrakrGroI0VB7/wzgesfhckixjem+1HM/3yVf05nuyor1ns
w8uP476lU58j5v/hIEiToYUUWmtRBcrpsJcbKCQqIDXaBL8B0uIiULullKgWwzXB
dB6EJls8xMqlp7/zBh29a6tF6Lh+Zh5uhvZbJ5Tv4Qr7mY+3st6FyHotnw525V/k
Gewem+qdjCNJrmCQ+4V4UdaF2lFeQCIAb+SgOsfJd66cCIOaOTKDk+6wmifbs0IJ
qwjBEeTyENjqF5h1KSgWmpWhrG4eKpkZEr9teE1cqrplVVOreEgn0A/v0KcIWz9E
fAd2UlgdkbXem/MrrspRiV/3aykAWwabHgqoN5l523m43s2tv4fJ9rvq6kTGLyDS
AZ2Ajfw2U9+Elo+8XtwXyNJfM0X+AbA8Jz39/ewZK0JW9PzJC1RdzNllmj99tOyH
/EyRjZGh3dfi+AXci9jpyVr71No4sBCN9QKxJyRQcaBDJcFc0/rWA8E6pZf5xkDc
nUqGZScfjdFWmNRVVnM3XT8NMzkPSRMJ+H+zKjIdUWvLic7JUxBdnHVqBgtu+oW3
SHrzX0pHxYcwmO4KjNaLpPOU9O2xYhnX7IDajeS3F51qXTjdSm6PwesKGN5oqZ/C
Ka9nKroRigkB9a9kLbXC9bsNdYxPm8LOhTJzCe3jyjAdsLmdTEzvw2sxRSVsWN5e
/6voG98iHV/Duz4ijt9t14oBAJ1o7BG65KIblS3myaFp17WIcjcadSfE1qlxYWqU
0mTnyCdtLpX0an6LhaAonrv4sB34KKOXgmZwrfgVdscwBBZjJlOADpa2MMp6wgRP
hct2Zz33apf2PHS5ehBkKx1UChnG/yQt4SwvUvRiRrVhiXG90zWD+e/LokAkq6S9
+XSDfdH7Fq+35+sjI8LkXsisZ9kLrKFamCRMuqZlTNmQYi9fsuIjNlj2E01dCaHk
4O8CGgb0Zw4rX1EnTMkBcDDcwlajbhXL5d6LejY8wa+l0hGguV0uy2zYLY4DBa/W
6wVDoZHOS+OzFyvyP9Yk5ElUT2bkN8qFBEh90RH8Qt4SkxpzTGDB4TmXB+4LCCGP
p6eeOLPKoTgNMl1A/+U+X/rofJN5klnuPo3vXlV4671h1Tk9OCy7ih8QuaLIXwVA
TXtil2JxFiuMREN6sFH/+Qkgk97lKlrMCvxG7U+qHvmkCA8Q9WHDc7CisFydXL1W
byZr/99/F78TjB+8zBbihSKPn0pyypPTBL1szCXqroukNRLSKPdq5XKYxQQEOSHz
HdE9EP36Z0LdxMtd+FQg/Y6t+EHfvwZsEYI2k/tWIba4A8hTuBQ0+3EZ4nCbeOqn
gx98iqOHHEK8R6wSfnV4ErQTRRcx89u/xT/7GPBdmvjJepYIwnI+vErytiJOpDmJ
nZApj4XJg7m0HT7j1JfKR+BPZpSUrKCtORutwLqD96GInvYXYfKIi+Ufm5wohO8c
0EHclmRzMb4BefKfAL4NIskrcp5Mxpid6qC+YnFMFcYiobFAHk6d34d8/A4Lv+1P
+5r+V/edAt5KenQO7DOPoWrnF1iXn1XhbPxbC98ZP51fnBtPjouCpC4bgL+74aB/
7pAycYPQt3rFfZccY0SMunNHuFJZYyHhwZZaI/OxqqymaiTm/nNXQnsopALRT/kh
mMlrpbxv0EfJDC6DaEjPmoT3yAlL1Mmw+e/j3XyNBI0lu6z7LO1N151HJcL2eh7u
FohDdKW80/kMzyxq5FMQHPHVqBz7UkJ4KRdd0gv8l6Vnlq6IJ1B38pHp21ADh6sA
f+SSem+2mKw4fngxAVOVFRhnZMNxCZgIWvxg6u9LVxHOPs7UjksiQtywyRsfWBx4
QE0upPtHa/U9LYEotu5oUjwGL+xtq3Ht1B+LYjOOhc8R0mmD8hHcvOmhYAEG5kbB
l0cnAWJP/L56Sm4oBSSuW7lHj9JN6UsKVkm/J3Un1SABJenSY6PTLME89d4mXZt3
tbAWykKdoLbKPYVhtYvcgWkRpeAGfTsO8H6PL5OI4y2bCeDwREGa/HSwZ72Rr/E/
nW4klAjWk8YrkE4lIoREuK68v2z3cxDWXxXgKDIaqjNkUhRXwQ2caDRYt4m/ezL4
GSMd2OT4opOSy8rDSYT3LgwRO1Qp013q/mg7ZTF9R1TDSdyGJ0Zs8MnAmHJDODG8
L+o24tNV47ElfhZ4bou+NTYyRo1hNvYP2bEtXRqI1sQg9fwq9f2sORpPnMroIzWf
GJuJeRFZ3c0lkEPusNlRy4L7TmEwdhVgD1gbmB6PPav35eVcfFSuHMpVY8kdYvT+
2LIT2H5UlePXN5yuW3BYynPc1PLPvBPZ283LNAkHWX+0Hasz5deFye4YdZEBRBOp
O26JxfGY1hRp3jOK/QJOTWJmPLTq8oGTq2GUlxp0qf+8YT1FshPvnlSUNF5FIVed
hQEYGY58RXCCnmQhsSaaonmxHMRtMtGGQnw3C655T5ljYkFw/auT8uBzjzG18cfG
PnXzBtAYGT5JPxvdVDfZuPuurvpJwtmsARfu+eOAkpKWd3GCkcGItPnpusrLnQuT
4/ifIt1Nx6oTbuZ93zHrQAlE2tskYHL6KRBu71qH0+Aj5EFzGS2D1dwPyjaDlu5x
hKPCcpWsOUOcW3sOtA/I+qQ9jekihk9Nk5/s/ISwtXFMchuuA0tDQzEKZWgSt4eU
Qooi4SoGm/G14KyrsCimvAdk7LJ4Zi80kd14rocntyd4u1J53pw3JmTwXRA0vBFE
OTXzJrahORcngqlvB28j2uaP1oE9qBulYdfVvx4Vxl+Dx4rnOna402WuACFAba8W
8YxByzR4R5M3qLqn9aZ643LvBoAfVGdt7SFoiUMl8mLnIH4T8LE6L4NbX+fwvFpv
DX7xRYmQuVXQj3xRKO6XA1S545IRKol7o5WMHqx1qOCjx7oOtJcRV+OYeaNjBn1j
GIVAtfFGOMimQJuoVc5dc1qZLNTxu4czdjfM1GvSXyyPSwfmZq6LMFtTJLvzA/0N
7BzYqxqxed89gFKADXLXim1oIVIJ5Ru6GJlDyPlSV+BDZN6LcZE4VF95hzBv3RU8
H/9SGiuAAdl5GO9ahk2lSlpp9kehkTXP6H41oyiw8TATqOrHYHinewpv8CBbIb92
W3xhja88sMYv3zSanaaJhE3lXqG8UdLD4MMmETiiwtsydJhQ2X5R2xMsDVEHAS9d
0Wgxd4Xi21iqJsuyuWtoC4x53u9DjmPUqJImOjzj5orhbSxPrjQAN4VC/0ZTlhge
/9L0e8q6hpbGJTiuRWTQNOGB/YC98PMzHqLWLVAJDrmy50SkW+7vGQ65mcaxsOXV
A5olAuPbZpHMBn8dyelW1dmeyhID6WzDBZnhV4GBaATBJ3Bxjw9d18/q2jfuA/jx
kOA1+K8Nt8CV4hAefhsGCpxyAj4dqgKAXbxJhfuFixryQvd5j1qdYaszpAs+FrLr
3N1Uhh6PEGv3gK2RcRm1tJen4ddPhxVDn1mviGAdoyYFljKf+uv13ytQysO2q9sd
XZqkj794+HdbY4Cfyuqpvh0WcJ51V5rXxan3iN/KWiiNJbmV68b0tUpFinxy8rM5
+84K0hn2hF0yfdad9IonyU1BK5D3d2bzgkaS+KrxA9WVelg0Yux9V4MvFXMxZi17
pIHkyqpCjwyL5VwKPXeYlcGU1JGum1rCD1X4f1/GY0noX5wyBPYMl8FEdonDVgyQ
I2xDdCnNtfMG9zBcFckJ2LC82S9LJwCxxPs02jxpdxk3Bv9c5Q9VJx4OB1UObqYy
40JiRHhbsgvKLAvVaHnvl/A0q+v8p3UBjWTY1LmH/K9U9FZx5lur9iMt82MQIIQ4
UHnXqRY7BRFMWs8BhIb8qAN0VlPB8HnXUKnpoR6J+6YJD2snuPuHRQkongAsry1q
4GLiX6I0/ufrEA+JCCLy7zFSnBK1a25HZT6A1d7dMOFRkNMbOnMIG3SEM4iUNHDw
cP43le9d4jQ1YRM4OlMBXEADKR7sKaZtMgsExKpiH92gUKGUYus4bA11s1OgOaod
tHSwNqs107BMuvWglWTV4Ou/2yEPNIhW9S4AGqkSwlcpKHZplCNi2gbNFsn8OQzQ
OaIZmdC8YZpfZz5nGV64QbLukt2Y2gO5kEojE2V12otfMNXYawERfVTjBTmatl2w
2K5TqfxIJOStmYSlnLVkPio5BbEoXnHo8ZkcCLOKLgyqZWjOFGnGYgqsZ0prEL3I
1i8z/Wr/SUZT5nMNl+oE5lkhuTXZiA6P/MMeW5PGTKD3ewkKRLtyZ0KLnpE74oHe
TTnh2J6jDEEUy3d831uPbm7y9E5s7soXwo7mwR1H9vo+iKPB6VkJBqx8UOPbPB5l
27J6sVDozS2JGXfdaNULs1eEtkdztx++YfLk94TQ2cyZy2eCxOXVKT8V0ZeJ+jkd
v0xpQJ/kEEXbfzw6ZcKedPwIx4WNIcAjQiX89pUzQmKl7xE0qjEjHHohdU5qxGVh
sISZX3Cdm8DPPpu49Xm4T8jVZ9JwIccsd3WkjLqda7voHkG4X+/SK4701YsHbojA
/VQta8DFRKcRPgTrt1cnV+7Um+UI9o/TPHSbtHqc7oVPszYEfty9iekAN2qbBpuX
PtGfrRyS6rM0at9B1BPna/2U/GuQPEB01pbFWiCvgJx2I2km8rxa4IN3fb4BGdrY
vyWiL/7A5Vvhixw97tAzgV4aOML355kg4qWeNJbG214rNqnhp2eqP2ZI+UOm8/HX
BTGpgU7ry22jvTbSC0bhmWUktOG/ArxXhSsHGafK9HhdSJn+NFLAIz9Uh8YSzJxa
mL2CJiMwvd3pqEqJGprpQUXifiiOIE/EnDsiMGCs3pYc/qa6UQlKMMYVA/sv24WB
zjZwMWDxB1R3hFsezNfXcDDdInNUK4zFcLz6jtt2Q0mro6euWqYbmpCXiHtk0D8l
xIJb2qhntk+gAdbC5Kx9JokfyZWCRGSqPr57DNtzKoLtMrk1cDBjAqMQyJltRrSM
89e961I3cm/WnwZaCeNhsegcX5OcLRYR6i8D/uecdWt4w95xOt69sAmh7xybw9QG
0D77p4MIXZAI840i6DtKeUxZ8XVMDDMtgg7tI8aDnZFDFS5QRvJ1qE3jz2CY/tq/
x77tyqV8MrTOxWGRlUsO9Byd3eAb/wGnt7f8TFnob8/Qy73l3SjLLPOxnvOeECAt
oY3uwQ9Un+geuaF+JIfHxuIBIe2ny+ocsSnsU5fwk8z0WKzdpHAO8TjRc9J/lbj0
Isjsm9iKd1TNLWXuJI/TIKz+2ZKG8eFDD3L38opexcSKtnxCvDP1DX4H2bxP1q9p
YIMegNkxew+MLNUc+EBcwkql3knZh94ETNMmb/Nkr1BGoArw8u1WyT68WeNb2Vd5
H4kfw9Ls40wpQdg18vTZul8u2xr2zMya9jt3phYYcqJl5PtMMg3LPE1SFkn1UBwh
y3gTM2lwZNtMIJAf0A/pM4G5wBIRgt7SSovYz1xU7EdUN9Vh5U8JCXbZwej0LhvN
My460zNc+Iwt4H/mfHnq5p/FTMyeuQ0z3GnMRVWn+BfsHCreWiAYFJhmQaclfehT
q4ywkOGN4Irlx28d37jsqZ3JB4bJD8o1b8G54oRtczyCZJRSZ8/coQJUH6fU2Cc3
uZTqlj1Cf/qrrUNKhzvTp0OHXqWa/R8NPSnXzB+X3I17/fZCuUOCyLQyKdF0a9GD
4vSp/NyLPaG6rbAi9W/51DLsuFmJQu3+oinyppxUrHSPBLd7bnhOf/5i13ms+E9s
GgtRoYOl/feKyEMSaHJuQLgW661H4NnARfuCCPSBpCde9TgIH8UrjLlDo0ZLmtt3
VdgZo9hiP8HgvXeFz7jTXkoi+bkDwyJcNBPuBy8S5rHxz8cpG7t/OJGwjsgVkkUy
cR8aWoKDXKRzYSVQnsc3w+EiHL/59thsstwJRqrMFY/tAr5/yIwgQxlDwgAovsUw
1hqm4fsnb7CdazzCsB5r8cLBe1l50A5/B9IZXVod0Hy0AvLccSwFCCD9/8qR/H19
kkHrNVrLlea+ubsfKQzAsnPbsV70AgK6GcRh8N8Ky12/iTNmV893QiCg/WCgZib0
itZyl8Zf9Q9K8kG7ozHmdPrzwgdvQPO6bgEW/jzVZk0zGZRyVPtms2LvGtMedAZ/
DYNvxSzU2bki9oDIUsAlb01AMFapMV8Cwbgsl289GWWRlH0Hz8JTYSOHLZ8AjR0u
VJ9/BXHDPx2Anv4aNUkZwg2hc6eMsfStam5yDOLiUw4lvTp7Y8nvYG8jjh2nqVSn
WdKWY3lvxCsTZduBj9clm5MwO+5ERe0qD+EQ6mD8i1GYueiTJU9Wkszh2QEPjto7
EMNjFTRh42ugV8AsoWOuU6EsSpvcxvD+sotM8T+nxDFW+A4KnFXs2m7qBxOdw97C
lBOuHzg4wdi1REmgXVvWGV6aDL54BFkBqHrcj5kcsaSaYcauq7JH+e88+ZIyh+ni
4jvBK/zETJHWh0y8YH+glUxQDe3XP3B3c5PE/Kls34ZBenNhUFXC7ff7jpmA9H1w
+rTEFBZnXauwAQOzhl8a+mQanDaLaGjrn9BmaZzvCUY6/KF6RI0EGhWII4SsYJ8o
KYx15+OCdY8NN23aB+KQYwOH0xarTqUpWHB9MFEB4KZEwhr450emPrOwkQEJ5LV+
90u25Q8nsp2flfu/kr+ebp5qMaFfR3eZNZ4AaM06Z8QIlXogHqTAxF4HwLkrYnKR
chBzOx+0GZq02Xjy9HOXEmm1gHiqY5yfkoM7ofW65UW/fcJSs+dS7mkyddqYVW0D
0kbR+2fN+QzAyEVKUfV0jejRh/eIzW9Rf7zknLdu+ROSecXD56EPd3Cs9+tuJhtZ
7froaxax8Si5vyZv7vwNsg2OEm9GrKAH36daWnkmSuiGrhbJsXRUF8RWyCYYRnaP
+g/EkgHY/dodDEKXvBWD3OS3SgBTTOzmV7iKFnIpaiblXtoBzA4qVTLjmgmxHUXV
sbFA9HiTqM1kCq7/glavf2S+2P5qaxnSn88+z2mgdeMRG1O7VlQIFfsm3atykJPx
Su1W+Lgu1N66YT9RB+L/wKblDwqzM17bJufGyLZ6/84bv3PxUvTbeWuxugFmsrgj
eYjFM63ngTNCDwZ6Q+eJIMSBr/xuo3KKzRkzLIUeP+rD4pqhGwasfqyKI0AN0qhF
7KnpvZmTWzasMl9K6THDy1oDrr0O+SwwFWH3jO96IFUMNcElcd/8TKD3wvJ8smM8
5lBVU3TEff+whgnQUVHBmMxHCHHhnl7Bu+a4BYOVVKCLYbBTygcckefPJtBoUo5q
vy4XG0iCWdhEkLNoe0MJtr57uoXEz/c3oTaP0T/CoGLZSCOE4Xy0YAU5a5NSgUXS
JnxR87oP/QYnp/PZa1NTs+KcS/WVetgRwNjltnZnMfLCC2RpEyw7Npz4WBsOUge8
IG7Nux6icZBYDDJ0Bu0P3sR7Sd7ztAG6bjzV+7l9venfC1veFYBYlc5hE2wx39rU
C3RhHmYI85jME4btyg3L/rWMDc/v3t4CjgdqC/+hnRm6YqqVlLwuDj4dI0Jkg3xn
U8nBpTUkGv0MpQrLv4IBjFDZYl1qErTTO4U7CMmKTfYeNahjx+FYlREDlZgzduMo
44BvD2/wOZ/DuNS9NoG9yZhPggVIYV0yfKpchyEcFtPhyZuiznsF42r79pApFSI5
21vJSaPiLZS6eNYFef5tapQVf+XS5ogYRvb5yTa6p6PqBTzhneAGgShsGcYxi3TP
tPZhFNSTh2sNrvsPxd/jNsr1GLpTRgWIrzpWcKUq5AxVyD0bCjvGTggiR4lZ+b63
nHhViVJnuneZQU/H9zDO7+R+5gzVmPDQ/qFor6xY/XViM1dPN3NLZGr8pbivvdRk
K3MYUunJCmF6AkbiokzvHBMYzHnGs0WWOia/d7k4gLbU8LjYK5JFdqXVfelbcqOr
j9uzUH4mVaSWSFSEoSYOKXc2PVjWNKtSykNWmhja0/ZTaD5XFdqv5uH+D6oP+df7
TIgUzJKMsWHjj+woXCZDsrmvDxmej2WWCi7G7I2MNieBEaLaAW8hU80+7mba6vKz
B2oEv9jjvYIwAnmtfbTX5fI1+zP1ddqA1lhxjVV/XrHkkLpW/ipQBYFUCtaUMZOD
uioMi1YrvbNAVgEHqzWt0pDPc1MsoLBZsrQA1ZApwdfjTweK22Bp+ejfjNbz0gJ5
ELf2UBLQA/LY6fDYOGCWY816VUnPRrdi3r7Jzpa4arO7qM0xbfw7G4RnxTLieS9D
+3QRNPQVWPaxQVuLusIRNWJjgQU3GU/SGLy4544cWHMvgZleV86f1wGjjegFBDCP
Faz8e55lR/F7DDqTCTwpno7WgxeaPBweeiFt/GdY2NgPhc7wp9nniVJ+/VI5Hp3A
ayHgR1Get4qvmUSxU0vPscy/GH6CcJs/fZkh2MRzJOueB/yAPYnuskKNZC9vS5rQ
kyPgMz0ANiQfc97rP2gJtri1Xi6ynhnmNOL8yak0q29Tn5NrwWJeri3HzXyLv6tX
PbIJefYTw1f9Aavib1qh34mm60KX0ALIHEwLoqP4ocd5m4k7dFQW79s30TSSBxmS
c/Ojv/8sZmkKGz6FzAZL3BTYOVqlbufzOeB7uYewJSibo+/O4ESTw1aJWbpyvncZ
63bRud1tL5Z/bfZXAWrJ0FjX95vW5d83szUyti5/g0iP6WIdDyvKi+urFeu7oxlu
uH5iIkkAnuIw9C8gQNeR3CJ6JmweLf4OiH2rAF56vJxCyDogbMiUdhVR20mj8AlO
OlQQ9oeSQKIWQd4rmhwkvy20at8kXqYsteeIvqtEDjY2csgbJGn81IZ2tAiW+xCT
tN4KxIHuo1MgatEkn5j4fJT2FDFuQGQgD7rIcFWXoa3NP8FPC35L6e7jSMqb1Suj
7MlYS0cbMWCOVwGx5G8NFscP44XDgVhNYPox1FL6aw8OKRyiLW8ELRKnnZBdzvcY
FZMJjWHC8iOmZSwF9CWcfWgriW59snSUOQf6k8pYrTdQhFJ0RzAFVkErD4Cvpzai
KhEhe7MHyAx6NwtAD5zqhdRdCIr6g4146+CZwmsZgVT9kb7ks9orE+tICS3y6twL
XQrvj2VrmXkGwYuE+5/bvAAGYPXmVx5DPIFIs5xhXC0xJbGrfbCFe/xE/9BCftKX
20UpnSThPxSK/8adcp9emddPP5pOB8r9bUpDwkti6Ek08TQum08lbdCpxHmEMwOx
KV2n083vqU7fcvHjCuxxLK/7r68IBCiRw/BJjgPI6+VLmlwwKIxI06Ga7SHO5i7Q
pyEkVdG1eoYidiQm6mu3R26ml7GNcTwFLg/BJBM8UPtRn/iQzdkTNf0jFRXbP+1h
SFJ+O9TEpvlcl3Wz+pVRRLKlbgH9EklT0tHW4x3Nz8z1PTreWXgB1xrj/UTfahfu
hkWw7V8w0m0zlhUweFLen4XZfYsdRCb/kwZvY2N/XingmTteqkGdB1LqCtTA2c3Q
cK+z8uC1DWXRnviC0xbUsDbzjsinpmDtlQgH1kKomOYTIcO6QGxoRtElirUSmxVs
EAPxqXWwBX6BA7bF0DimGFY2SsZtB4EPxFwsHfgiYpvn8AIRkQJ5fIsAhwZjLqIq
N8XIwVZ5t2lnnCVScZm0zXTT0YbVHmKHBF2FZo967TGxv3GRd4JWnGNIae1Uzn9f
61zRTue69b16eIzE6Vnbb5YnS2pl/Bqjf15Q8wsmegbbTI3fQVKYSXsjDwn4I/rR
5qMggkeOWXNhQpZVtN8VE6hGmSVrYZrKqF9CMsm+HDOV+nN2AldghpPnyHX+frQh
fz91TdPpmrljlMYIjCoBuSHoS0szQOA9FEsPbdrFXGxtcIGbY9kz8okETADyki67
ijyZTFo3Wv4+8ClFO5r70pSk7ghh5SoXNzurnz9VfPt6j3nMZP/OOi0VOP2w+TLY
RiYcSC4dZNY86scT8TPYD5nc+j88ub/HXYiUEHBFpTfFWO99g6+P/dY2QILzPpkM
m2QHHledh3GUMhIuupCsyS5nEw/LM5vadaCgJopULUVIkPE0ZgBK6snoMGa3dBIW
f3vlUTBVMmg4dNH1Og5Jm/PEQShgJ7oOeUz3Mna+897aPKdJIDwT0o1GONBPvLYd
AkRiTJOqLKGux8JzUaiSviNo+23HnDGGCQi2nkqMK8t0lt26iXwhEwmbcDqETKXj
3ECqi3rl5Lbuc9W8xZ/EWCRgnbOntmxVR6qiZbwrixucpQDokzs3WGo1N9HSMkY9
ONFfzlqzJdpyax2Cr04TvkRjOR2cqCzn4EcFICUthhBQbLphg7evFowBtTSYD5DV
ZctIseo6Aib76JzBCWsA4kbFCGAh23nQy6taMJdOfKgD7u+bQyeGfU2PtB+lCY/p
/+osu9fW8nrMDrV88dc4aGKF8AuNUWs85ZsrqXXZem049fS25/g2D7ZxAxnBsC+U
sql+3G7Fn+Z4DP02+Q8/DKda9hzrVvfu0xs/+m2mCtgD9BPZjdGDC6XH4XGQGru7
BR83wBDX6KQFl/yXT/TGtEH1eGQQSfoIcLVaLvMUIDv1qL41UGgZNqwqtMmf6DIS
NmOs2So/DxTdhmp7rK8ZugCzndQk7iTnQXT+5N+0eQabBvpZlvO3oagiW7Q9FPOJ
gIMk4ecMYmVyOGyT55mcpnXdv7gF668UlLME2JlFRkaVdAWTX9543Krxh1N0HWc9
XZSKz53Kq8tqa5ujSaK8J6u/m9aL9zINy7hcIXevAbmt/8O6MAlt/o7DZmSXrRxV
XI1o3Nfop2XCrsB6meCpnBFY/d3maZyO1BhLlVe3rWPFY1rugN+oTSE/de926K4B
wyVEedNURTv/V4o8CHNvENmjClV2+CbNxNCeB+vKQuMlrjvjm/CDSxK+ajR52RyW
IxMPZn55B/R6EfuigBJVSdmZ08p1rWKvdoC7PLobNgZd8LOYB0J4GwNv/R3uuoyP
GcmMlDiljionNxwU+eDgNiVrJ6N9PVSfdmtB9cY5IpsqwRu7nmxAfWsvWrtsDlWG
uKkIWv5ll/cXKFERrahMFPm+8hG/pSlP7fvGizU52wbDUgzVJoZldB7i11cmj7do
JpQ/vb1664XS5AjlrevZp6DGTw4fIcysApaEDfQXROZz2lrMYe33KR60IrdIMPXr
IsGBcSzfj/crf8ej1vjkIdNYYFg3h3FlNSnhfTWZxZmXR6T8T61M775P3RQHAnHz
65gscZeLaVxW9FkaX8i8IB4jJtBXGq1fU2dQ90GncQi2EFL9zUlbIPw2XHjfuTj9
3UO/UjZSEYFM69Y/XD1sIx/bgsiHXtwyjm67tl9V8Zhzloukm1aVkA//zGwsqzNc
+MaGrIdLwIoiX2DBlzDYSNl+1LuaarMo+FXE50aYx2MwqYD4qSELbiAsMnHFroKR
dv6VSc/C6wVJ9hjZLcF+jc3/XqFZHA0FmNDCHFxYGfcGm0bXShC4YBUM2QoNc1QS
K8Y0Bbhu2+cbQEqORFlfTfsfYGjJ4bs7jOzfAvkXfqMMeklflzqYpLA5kjfv+ovb
iGcaQgZIhlDTRf/Pu6RW4vc8GdqZM3cy0Fv/PD/JvzEdzm30zjZe099j6MQiD2ib
+J6/Q+Om1DWEGe+n1ZTxB2kOVpu8YFNcq3enMfUCJx3HRNejMgx3442fizPJ96qp
XVYr7owRLW0EPNuITHUGBYUnpzphCHQPN34fFGv8z4tBvVZcTKanopU/GXr0vRpI
QxIBUOrQgEnVUXe/GVtLC4LA1FUBQLZH6leo8qbGH6SmT9xgeEarux8pI822l8ii
WP8vgf5ySvH8NCWviPcCnX7EHqlVg7n40Y1D4ok/fyGKE+FNRBWIBRXZdbkuvTXZ
AstBdhvFRstvJtqYect8c+qnLCnF3UYRLDKiwwihdF/p1MCEasQ8f5Bc3CyULTn0
DK8H0dK/ekOhe/ggyWV/itMuFD1ZWLRFky2tDpzklqzmUEyMvr8KU0k2PbSCWZ7O
wjMpXg/PbT5MgXXf/MRfvykDLS/1jALaMSbyrGHSQmzzArLvyVY45jL//+pqZHZm
A09EED7BkRK9JoEiSp2MGtQKUKhJcQxUYx2BPSoUEn6uSX9AA2xYxbmeU1TM5QJg
ibf1DoOlUVOIObaYaKXmVbhmoBV9KDV5EOd2L0W663avIW1TgfyGXglbsINXhYZL
BeUsSp7VnPaQ6lmiLyQZqpqGcbsClZwnA/jiZjIx9sWbDtUMQZXKzJazSYPIlvgI
vsjbjw09gD99xjytVbb2zEpdcHHh1v2qvVSU0aJ0Id5ZKp6J/JdqBNjvOfXPFBrR
Y/Rwr3eG5PDDEp0nfrYvFy22rEyvkfuAw83EXZJfhi0jLiwSGgZ7OzMbE30ppJIF
L+ulMWQOO/AzftXxes3oJWTb68L+8BtilQ75xMlcpDe/leOpY0nmpC1f/HY5SDO9
a0d2gfSKKBZXmzyA4i4YoneJPHQcf7RmYJjA08dTpjv4+DeyMNMhBLnjg9Z5P8J/
BS/KfNlNF1k3Lg5TEEj1Bed6M3FxKJ1F+5zKQ43jd7Kz0Kv78jxeEfi94D7CuuHx
mCdSyFjnqaTLFpn6VxYnM5M8LXCRQX1kHzwcPf/RngpP/9lLjlPcBzojkTWIrSAp
1RsHQ0zgs6DBAAuzKy4/ThCNsWXshj3JPy03GEJC1GrnJLxWocEA7SEp1cfx1oDI
HbBHIJL0+4Y5qGNsJQrfuoQ2q6W66NZP4CejSePVTTyaJLl3NZWmBcZumAqFmEfd
MSak8PpNpbI7TmDn8cJKF7xv7kDygtI7aKwz84if3siP5YKQZkWR5SLoMp7FVVK6
RKcS2derecZrF/QxOMd7XANEQuz/1f1ZOIrpbzzRQgnhI4KAqAeRwVrAv3AYW08f
6he1LqmROdFcuHBxmxhP/JzGaT09EPRMXF7j9G+m0l5kNwSGyu0kaBAv8c7vjJf1
ED0ATzyi+4VzgED+JIm5wc9+9vWb7aYQH+ucuANRZMztGUWkzJObhE5okZc1Kh8Z
vC9Zk5BuaEIGbL06RW7gdoZiXneiNusEUkj2h/p3yslSkB/qRSpaqmyvSnsgU2/P
Y4SbEd7/9OTJSLP33jSBb2QhPX63zXZ7fQVtY7uH3e1JnZXtZUQk5vQftnjM/s/O
/EgIRLNXEQp9roYU/Vy+gwgOs6bZzGpjlMvoJ8NMNcPWp0JMLeEweC+8niCqITKp
B7YsA0p4Ig60bwPZaCmrd0AObR3LaYmEWmnPOYWYZtaHMEQXK2yI7/g+x9PgZ8SH
VTJPt47ozeMlCjkp7fjLY5vYNeL1soW3WlQmCrh/cob2wiqAqZk2O2BGaexpzT+F
8kbLEL+RNYnaDWq+kIvfpfUa7ytQYc8/SyFunBRmRgpNdePTBoEghpWft6v4GiGQ
l+gEwTYtvJTbC2nRBIBbhZwQHSUyvbfWEMgisaI6Iul86evKd/TIbpzKrdaKudDd
XZHjbP6CCIa5tM5QpcSViI/9e0hPKtnXcT8O3cJeqr5BIbDW4mb3ztmpVh+wRanF
AIowVBQCxNV9HLJ940n528cKIRWIxfvVBRRHqR+8cZ0cufEuQcykClZt9tu93odR
E8CGXHS2xrE2dzUgys1nQ7WKo2vZHPQ+shbDRuWscHkS2LCVWtyKpcaJ84s6kBem
559xRgu264JUhTByRw61EmDTDsh6DbZXEmqxNxwef/Iyq9CL8pvP/dNQl4ITLV39
g+UJTmAE1ZBakIyXrnd9hiqciOQpxZdWpC60b7CNJbbiotwJ1ljcngj9ieTM8EZf
TwFy4D8A5/9E5TNJ4b4qGMibLi0MTCflkuKVi9tDmjA7wWVUGVZSCPtOGQGPkZH/
M7bb86EXDTX+ARdf1zszJ7KEgxJlXScEdADdXas4Lvhb+CbQrYLA95VExKaAuXqP
oO8djnqmQ3tCovS7LqjA9ob6QVtMWVuLzXUraIzlITjRDLBWSOYDkEpLK4eleIKa
bP5ZbwHSlTUutT/yd680ht11Ngbwrj4ae0jp6OsS/r1U1wf6nStNWQFROzok1Fph
TdTJWKthMfmCXg+LurIoKz2SrRUnazqrVsGNClcNVfudHzjcmgpaEEvYQTVLrfFZ
YsfA21vciSJfkOqVlkJD1+YE6tT3Y0czNqjHZVlmhTBuhuCZ0z/qW0xbvGfrz5vK
Z+Ydvav7w0hemX99Y9zGkskXg7aQpDOGsU92oMOti1CrGaz/JF0yW7TnlTnGvYfU
2ym6HPS/GsmZC8jFejMNrwJ/0826Pb9VIl16kFiOZBfVFfAPhRJ/LNkqNBrhCeDp
ye3SLudFqpqam8c5JCteykhsd8YL/oyHpwF9QOid3vzAT1oU5KPuhdgkjZu+XamS
DFg/mHAeXVdnsV5nXp9Vi1TmR1LJZ0JyyGueLn3aFoH1ykBCqGCSRcGLSHw6/rlY
UhyDUMRu9U8jQcXLynxA8fVyYkxdjeaPdHj2XW4hEMNzzrjJnfbWn8A+JjV7Ygdx
08VoQsnImxOpkWIKjJbRqil1Gx3/B/NcPocge/7D90gWELKIi5LWdlZJv0u5JGTg
6nf+9ekCP+//1AEa2g5/IGl27DJ42JUYrTHEdINCHWVX+gcYxKYlkYCCeY1ruw6t
VL6t3wBC99qTPDD/M5h0dZYgxjxaisQFYZejXtdoKNJTrX9PpzBbk90NJDcWezQn
5Ecf9QCQUOXS8KfEJ7OGQSdfXm6w/+jvN2L3F+cebIujIIrn9g4n92lrzTYqVG+R
s65cvup8r/0GEYUrRihVD3SJaPCZG7xrkN6CyNxNE/EDMpk0VsrwwMvfsaN0KCv0
kUqx7E4OqFt99SaZSPTpx5/NO8Gm6Kf8RfLqXqqCu5Q+cMKwLAtk+o6bCn4LxH6b
z/3/Ps7qRq8jd/AMIsZGpVVP2H3aGYrT8zEagyOyMKE5EwKprrrMGwKpVC5LTxO3
AhNDtX2VR5nyc+fKqNvblZ+RqnuNv/jUUy37HuhjJMLpb8bzuemmHjNBH2qgS0f/
PsaBGGtDB384vgGj4bOVbFfqgFkdUBUU3L24KFB0wlygwEYue9De5vkKmYx0Vvpu
qXdlYTMhpm6AnvbAncB7bux+RtM9S4X4lhGBcfcNY8g7VfM3VdWxWH6wH6Ezyh5c
I2ZmfBGi3p8MyLbd9O0siPv2d0vuJYyO1Z5OaCLM8hi0E71X4QoMFJOzkbQurQvb
UL4Il2CSIZYSWygifp8dAtdZiq9mSP7cxQirpPudWLqaQKjBX6CgpA52rLF/tZLB
SdfdDBobdfQAaFaNpPRrefN2yneim/AijQu30beh3DeXULw1sEWOaNqR7tv0mg+N
kIc/zXx1kJze0ASWRgW9E7QBp22P/yDdgBqwadhMflQSz7Jh0Auz8cnmX6MD79IJ
gbPCv8caGhwPEd58466hZY+H0e2GT08U8s1IBFoxV5ibYthNDBip+BBfB/4rRQ6k
0PfPD73my2D6fPuPh0hHrBWNjxmnDEY0ZRNnP5TrRZhQCqDMynTV+wTLvaIYFOEJ
NI7BqKyeyDeh6lZVk37a4l7Us5MJxtVU7jYx5dmIfJ8PgpAZYK83mT2pEFoHgotR
NQKzns8uCWPkhRIx1J9URoC+ePNTyuCC2IfAQ/rQtMBEP/DmProUSYHaSudvnSo5
8+lZQiISrC0XICHLSi4c3nKEDKF9//ww4nJigwWCEwdxqynQYZTqFG8J/D8i1pa/
nds5Ne8O6/JF5deOeHqdCmR5lO1iV42UWIcveSSGEWwvtirlkrTmd7nbf6uIs3Ce
IoXs5HqxZhPA0KN5XBKWtWyTq7TNAGBx8j+Or/ulN8U/AOBDmW8bZliZD9awhwoX
q2/GM/oHYltxH6Kd+VKBPkbnFpXu3fLCQlAMzUhDXS3JGv5FnqEbeggNZc+5XP3x
iGgi4ItzexWAVvHdZl52mXt9x7l3CZDvr+u/oD2lfyLU9lh7sATGqIP560PKr6DI
xyIlWkxhYttpzIIW4m7zomwZ/ZKC2+WeTBcMUZwyZW2wGG7jLr9/lMVasV+EKX0E
83vlIhQuX2yZKVUYwleGhuU3puq7uG7WoH0HUwInuFLc0iImy0lqMgFpDj4NPKqd
EMkHYpchmZopVBldhS1KsBhSnYqDPMYaum5iotpytZ9aQP5TQjgy/Apb2GELL5P5
XCf7+JzKi2v6mq/pQWiYwSPFQtYXmR1wIh7cMHIX50Qo0b1fGmW6Hewxo3GLSSEp
o4s1YVr+emtUCrS1xxpQnViOq/xaL48TMNAb4bwNzdXIHALrEYQ1NrUJbU9cZoAc
6Dh5bSI2Afmn61o1EwN9IEYtxSzL3jIZVMkuo8NkJ5MxJ/5v81NuZGO1teaytIBR
IMnolSxPK4PVNXod+BuLW2BpxgZHRnhNgtPPsstFuSz0TimwDixHWjB/R8TUBvJr
z7tWtAYwD8owk64EY87Q1r0MJR+1TNpYdhX8Nh+nMIkndGJLD2wqRPVuphMBKVk6
32qYJHNXCM2HVTzhy2IXF8f2m3KT4rKxKm6pV2fMFBNziIhlq0LsXaaXB59cg8oF
HwCfhjz8TMb2pQUiVsx7Tzi0cIRNa9cCO+at3g4yWp4+/ekTgipZpVOg/8Q7rzb7
GicPR076rZ5zajS8Z7mgxi2J+pVUaz4ggM6G0d5VHTpBplvQYbJjQnfFx6g0bjgf
uHNxZdOHy42V4FhgxLgJd9fKA/vXJGTB3S6Ag4FsOGwzS8ihSQm0W0OXM33Yc/oN
ZRVCGVKknxzVHknGbWVJ6KYxEIwr8fq9W5UoNpQr8/QKbcprxSokjxDqJazpH+pS
2NoK8qVzsz1jFnBuNtCXsHKGoKpmwbKNTshJhE6kykxJ84oUNALW+Sq2w4AO5wsv
I4AUj1Ffqx+88XnRVQtqgVJGhqWFiNpZhXGfkTKdBjFxdbSL/8FujacKZECIpDA0
hU+IEyTKXNh1yi/73IgB+90EMdHe0QIb1rI8QaraqlJvMYXnqdwVm0WVRfYOH6Nh
ltFnq9sQGmjr7YQc/dewlJs9Vt39uODoBZa6jSG108WyLEQMd+OUphQNxYuvuTUG
LWNBs4u0r32rPZpa9xofQ/SFd4Vg55s7YZ8hi5csbOK+tQkYFv86FIUvCDhY0DY9
TVT25d+scEkGt1P8RsGI0RiUfJ7qthSzMqWrL3BA8RJualPwXrawJPqmFPNdSJ+q
fpapGyEwJhzJZUIazEPIS2KhcRPXgvE+x7ABed2UgBXLru1fkfFxAgaRs7/DgkhU
qrOR9XJ/MmuvGUk+SHk70cIzPoH911AgcRLdgLPpLIM11/M7z4xnd2zFekjqvs46
nyaOCF7kbFsqzWsE8GDGhCqkZUdqU/EI5VMxgGEUIqJ3/CcuA2b0/MtpHDbl9Bzt
lWUgHH66+WO59kNVHaoL9IYQPT9/fNJDhekH719J2Snz3Gb+enGCJF69AGTmWt5Y
62aE4oOGt+zbHIX0SXka2jzsW2TsD4gldrefmZtO3H0ic+Y9Bdky9/v4PLZ14RK+
a+2MI7j+U42A2N8/+9Wm5fFhlLnQtd0ycDtpjEKAZnDJfC3itSpHl2rPF0qu/GSr
9cw568hZ1ruZbQUNF3Tf14aQP2GPBSMOXouDab9xq49MtV51xB0akK6PBapiW7R7
qS32amUDHkStkndUHf/wgnzaYJFxyIRIzrlNbySWrO/wwUHbFSEamdHNHfP5kiPr
pL4ZMRNXRnH8gnv53qZ93KrrmmQI2eJFssh0GQX8wadrPqthz6iMHs3ae2JcUdKG
n/2mrlKj52VAPbnfeqJizYp2m19EEJnAyoGfVRoia5ntvltas0h2yPrdZbu3W9C2
7Dg1w8O/kLWO2d0jMrJ1KL76Vd7Bm7BuYw0CXmO9qhLSK2Xl93//f/EBgSsN9P5c
FUNgxgaXyG2D7HNDDsDvMSdSFuwLoSYsjvclx4071lrqlHZ7n1ecm2LKdQ0Z5Ivl
pIzsf4B+hGCkrJvn1G5GWlT4gsEuteiOiGBxRlVXgxuyPA8pbyIKALjH5K82g4kW
dvHeasmk/LFl2C2VKacyCGVxw0YK4REX8i4LrqhxtO/9jKiHUx+NpxDBcG8sCEob
FJp8Ik2ac4ek7oCPC6KxstcboNrs2uAPwK5of5knnVQrw7GyabaExVUVEb7LFlxS
QF2Lm0d/oC4KPvgzaxO+Nkj3eAtg+WGcEsfaPumba15sUNssROL86wOhfKPRP/0y
pqkVazHC3Z3S5p62gfJIev9SitIX0vDRVG1IXfP3k+OC9Ch9en5v0DvDTqdsLWsQ
nifoZ0DA+jkKpkBfFVIsUXw3+wp7F61vP4CFkSlg6DMGqOigz0M+8Pw3YRGZm1Rp
3izW3hLVvWml2vzGUzlVpIugM+n7WG6iU1cZrEH79Zb8MSR3Ezj6w1aM4IA6ePzZ
WoxjqE2BaoaiFmR0/N4vFaZ6Cn+D3q4zEuPMPuMCGHxT11TiY2phKaT1XbUJEI0+
oDv2iEvDTimb7IJW389WcwBFl0S1NTOBeyU28HPR5904erphwRA53cwNkZlFOEPx
ORWwctrMfQtPrb2QX5zsuB9DNT3SsFvs+3/sOR2OwhjTl9tldAT8fl11EBwOPNT+
ZbXcC6GM2h56K/MDhyidZKV+/nF+rBMbBE4inNE6oIB6gMDOzEFcy8x4CXn60ln4
Owbu7+7BkXDUoFX6Caz8KXbuGy8iUt2EA3/Yw3cIdLNw1eVCUi/yC8zd5ObtsWsn
m3soyWKOQYt42psI4I5XdBJpGKVtrhK7j/g+Wi7S/bA0pdTe6cqmrlWoezFuOhFX
/N66uRvg12f3Rj8q8eG1tQ416mdvCJO896O/OYch0cFQRal0II2uoyqKKG5xJva1
CUQ681j59ZriUkRm4OocsLgat29pxpubq1qTG5It/R9ATe6I9d4VLqyPmANI74zS
JRhCANlgBiK9h1zhw3GeeLB+pgUQ/y4E0ObmvhnaQIVMlkzabVFcHTzzpbwQcGb3
7LEP+cg1ucxnHcuxVgfCWJKEPTo41/y5Rq8vHiuz1bddBtm1tJq4tx+IK5s+bhNg
KofwQvHone6B8xwDZo8wLmGAbEgkdaBv78NnzoS6C2BbxTfbp/graZhvLgx6zZEp
x9fKSz5M1LWANWYDj+iSP/xfWRJz4hs6lCfvZJ1bSXbegBTxWCi8GUij6o0wuTvQ
+VpUgLI+27i9GTep/2bL02RMYP3BRCHVMGGT9WFQUPWSJLWvuySdBVPLNmXLqU1S
M7VS747GuCsY9szw67icJ8DWzxSwlj46Kj53IlgjLN7J95FAEFbSq7Hn2sHcDLcn
rOXWxjCsdHXUdQUEBniOv0MNrCW3SyrX2+n16ZP8anF6CtiZ4WnH2KDA0QRFeT5m
ZLkFjPm8Ishk/KUYEsRGy7qO6to1gHm44657Ix3JOJxaRNeFnKxNc14ESaE2ad1n
p9/BR+jaZhG7ceM5mjVbCw4fl6NmKQUeX/u8OzGD99ybx14ydYBF5CXQm9LbDirT
CS9LtP+a2ywphvJkTRdo0p2SrSQZmZm9Mkd2VYaR0cLe0AmxzehQHWoviYDsUtiA
7AhFUnRqZNMWKvJS7Rf8V8ffFBCnJGw1lPozZ2HwvdF8l0npSMffNXjAa4Q1VpBE
3yGocQ/Pld/O7Y91vdDo4+iH/ChbzGURWW2yhX8NQcptt8SJEfffDbq2LaEm0keM
9Y0uhO1tMNmocM8CC1+MqHw6EOj6x9IktPHTV4SQQK9ViXv4UFvopJrpe/+UVB5e
2W87J+IGT3o6p/s1iCuUiRVq+BZ+DBtNHm4OofwIimK/xDB8uUoMklkJenXk1UVU
96zAwQ1VUiZ8jDdfwcYsuFmcV+w8vPM3/ll3LBiZBZ17cHbcaoQCo+ZCeY92y9BK
ZmcT3m8pfVbNC8MhAYR4gK3og4pP+xJiRSFXp7vhbwVM5lk5UZ8U3SrFjLXd5R/0
rrzAd6oisMc8PJxzIPuJs58Gv1ig5TbazMuSV8Dq7lnDnTPV5G1g+dfjb6LJPNiP
loN+GMOi+3MmAdKuLfD+VApA7QE78qp1W6c9q+FcFclsiSag9UwwgA4lilUuGzjb
eGOd8qzVOe2h1NiGEtSoRhSXjzxElw6jNqSAJ8dxSMnbvNN2AxEU78Rk/uRiBspQ
bMD+O5292T2ZgiZFah0hSaRtwOrreprEQ7iEnCKIYRJZZwGV0t7Q2+hVR2mYS4Iv
hRywzcrCglhWnqHSrksYj/3Pp8fKzyE8rAHKcLHcJGeaYfFTGGsIgnbI/Pqqixv3
H3kGZOd6qUr/TSiuRc6HNyjwvEnNzur1bHyKdh3prElhL6UC80P14ux6j/W4Sq9M
lUW2nY+QN9E15IwQjcvwMcTT5iKhKV/AymCIARIihegxqW+wAxB8ZVmAGPjiKBHZ
+kJENjdjwVdzDrdwnc8o1w96yj0qoPvP499cfKCYPup7zjZ8tN/saXrhGxnupzVo
uXCbnSS8rrVactMPTJSKRU6azjkb8UApiZKbKR9JIFXwC2mhV363JWuMa3VarnhX
MVcy2EuGzkls9QtUy8yqhNpx4f51mr88jz7qxLSQ5V8xE+pF2ugg34RS35u2pbkt
K1Y963mWqnZrnwhyGUMSj9ng+DHKjqMrm8zZDZ52cFE0Aog130n7zZI8JhIJyWnr
2Ptwj5+Ky5bioeDpNLneOWT3OKabnpERnYUC9Fa74vSPKumow/3CvtEyez045m17
XqUwk1EquzCNj73hZVQn0S5u+JGVPdJ4TwuPVJBOjZheAERyhdsSMmFPz9Mh7Trn
oihzyVlcm7gYgAb8c49FmxnHVq2aou2spCt5BxtbaNWtP7sFEt/6lV8+mfsmnCKt
DqV8gI3PTMqP3dmTBSc9lWPatOl2D5bfFR3r5RlIzswx6fAAvNT7RKJPgOu9GIl6
PNwD7D8MLZZ3VWafefbVotsFmJbp/Txq6CBvNHPKXsNJg+BJqY2x2umsJU5j+bxY
NYe6CjEYgdgEJfCau9AaBcy+huz7jzXmuvzG+fhAiBEMf3d2bkX+1NKRGOkpYydL
1VFjo/3xCtUSs/dnJhr+My80aVV/ow5G60S6Rqv+i6YtbYySeoa+YeDZKTh3Mln5
4c5X5tfRpMQjdnnTUZLrOt4mc/ugQdpl/DWzpi18cFPurYKQz4EOhfPxYvBZmyPh
ppVB9mux5YAFu3l+/uCXnPo26jGtwi0VKNI8miwvV5BQYcW6a5OiCftztXxyhZjK
wpIYv1HpENIIKt6l+zFjP8sjs1OEdSjS+LPv8CkYso7bqkF0tffSQDwe4LPHYJ9V
fVrqiK8DZRdkWCcjRo6HuTqHVCjR4y3l3awdZJSMs7t1ysKSB4Ux7w2Ds0GVVnQB
avM4HL9gSvJ302o5b6JDghULOMr9LDnLZ8594F/zxFdQq8yrLCJg1lBDCCNGwI/9
V/8jLEyk5DhmQx5F5w5gLfs0G09eZ/bl8pscEMOYsKnn4yMOWGW2u0aiSKrETw7w
RpXquuHhYPUkWuDUmzHLoB5w2ga0IEfjAZweC4a+xPIZ1ThyYzsshrtJGBI4US27
hc/PkU4cmUop3z/SAjStDb4qUARtRYqgI/cK23JLFMMZg6dvx3jAVZ4nUWutnNgh
axWDMBkSYKtzwdw1JASEXkAde7MIEEh/PHa2euYNH4KTb9Dp0VxL283pzIyKUwmt
L9ShmMSf++9CEu3tqJAMqA3Alq70HF4pbRLowoNotOM5nlAqKtxn1KJf8LuEmLMM
ez38I2AUoKDWCeRuuboXOSOWUUf0PW2PRImCcCqgTOQhgpN+dLOqHxAp1ELgzegf
WJdN9gvkaTlc79AU9Sf+LfHEp646WlL/bixRElo0AWB0hNU6i603wI5qDtsizsv4
aYrVw//TICqTwv0gH1KQnEdARJWAm6MISun0U64c+xw0qu/hCdAZzUcWe4LjTBWh
oYH760EjpOin68xpMDNgReKp1rsx/scJRLpQNFj2oK5+w7DI9szkw75L0x+DEHWw
37H6tfKbfbnfA+AoM04ybeny307PecCS4FdgAGfrljVOnj+Rjby8FqueQPDUrKEe
JhhMM/408mrlwa94+D1r0M5k76r0KHM8F0OwucFQwGtV0l8JVgSnTflXsjl5SdVo
RCkQ1CNuGQl0VZw5bGpOlfoqclxYVoQ1GwtOEqGLlXtmjgPCFUqRZdf1nXCfz5GM
a0oQ8Yrfa6dpAkqmam/7DAYs692sPFAEHziSi7apn3R7/Mzn3Hu1Ua4icIDXVAmw
ssJFgLdhMl5rAVh3XoGq60VJJLxrCsQZZnzApTWy92pSOU9QWZKOV+VyOMm61qyc
lsu2DmM+1IoRFMHtAe/ihOVZH3rXdtUxAHMk3DGJWW1REnZPiGJbzIne2JzFsMUc
dEGyVhYxXTfmZB5jIoAvR98WSWnlJFt2Olqi/EZTGNHdfhzprFkQmNUuYcZmSupt
3hVl/KVnSR/FRGYd4FlW7WmHzWkRPN6s1C3JSZJW+UGKptDiPAOs2g6fC3GmxuVS
VB6wjblNsBe07N5u9y0K5vUh+W4lESEzJwsYiUanOeTp93nKsJKboITXaMO2ZCct
WNW4hDWnksnncIlZmhqjz4icoiZ+6feB/JJfPYbEo7op1/tZHc6L9JI/cPpB8Y6f
8k2HcIghjIXpjOSQPtnC4XS0tDdkheV/e+xQmR4bMCqUK0HNxC2/PzCN0TAFoEsp
kI+OWLkVSgjWBnykVNux0wZ4kW6o9ukX870ugWP21FZJT6esAmpi3+XmIgMI8Bv8
ZylRM3ztF2kiQzQkSBj3TzteSWdu7251uOV8EKq8KJ1WVWwn5zTyAQJxPZbOsvoc
U8azx5NcKB9ZWZzs1Mtw07YLQYLXxRxFwX0f7BAI1XLCKLMLZYCXa/+4k3nHAnH2
+XrGirEbot8aVKLY5Im/7AaCRhiK6AB26RtXEM/zRaP92s91IMpuwhppXOIE+uiX
pGS4IyL1prYseacAdt4Fk6vim9UbX9dP5fpBTL7dE31jKnUhwvGj68sfLPEYY4kk
yX3H/bzTGqyJkvW8jYQ/qwtuHnTEJjxcmItuXKUX94GvhcygOkXQK+pOodEbeGi1
W9ZQfh2yRZRcSqzU12gEnh0mMJKmwZIxB+8cfFnGqchE2MF+m6wghn51hLFgBFM1
FVdBC4Q+QykfktVPMMMM6ATsOZlJ72YmnofALbeHeM2XUxGBggN5oUqoax1sLGOc
JFOp8Y9MV4EAvO58KbV5ekNRNe/UsWyrY1aBHZ1g8A1je1F2OnIgXFebD5EOZWYe
Us6RS2XfrUOPIruR3x5nWCrJtVhSy8XtiKLj6pRJS06LlKX0k235oasStNqkBfCu
VHUM+jXZtsgM67ChU+SsX+IRQMRhmhrKdS+DZ4jqLHZYbEHtOnLU8exAVKruhQ3X
BbFDqWSxh/h8VJ03aaEJhqTJWLWCeq0ygtOkV9bdVH3btz0/pzYHWx450dcAX45Z
CjelTyXtl44RF3RErAY89J+DoMv1vvACburlEgMiF4ZzUqOi/6+t0e73rUN6r8qR
V886bN+q9RlGgtRRlwBzm7Q1m5lcikd+W1uRvcAgHmB77KkBa6TLybRB2ME7Ob27
+1VWUW0g9RlaSEWbe5hdgTxaDpS07Xbeyxr9fz7zse+dUTKM9xqcCRvBJxJoX2Oe
KDZ/T6kJfBiHrHDdIvGoSbDSeqxskN1IVkWBLm30e50Uc9u10KYA0cO6rfOcsl7I
sZt1uTo4JRZYzefVCTxr0bF1GMDfl5yV9cwMb1f8meydjlKZufVpksy6x3ADcoHc
slWREukA/jxaNObz9fagh5/srLvEzHJucVux59CVXAHk5K4In4G+eNIuVILCSwfd
Uz9nD5Lk+Du65VKBthHBUTW1J17PxcXcG/QzaxxC5qMlihhZPT2WRXNxeXPiv7ab
EmT7iK/M3he/yOjkBMPgYM5aWooHo/Iiy8gnU5xb1v3KzEO4v+1oWJFtGHIpOSS8
UixDsno3Weh2Zyg/xJkuw71reRkeL1LuMl5MbwsGjrmrMjHt9zDcb6eYWYWqm/+l
OYTZ2tC3USxbx6sq3rSAP3qCMmovWdluGMAeae/4jXNPtM7blMXucZ8DNujCrIRj
Fbny3xN7AUOM9c7NpLPIFtVUMp4ze0kq07Nx89vI9SWdqMdrBqibDaJtpPZGJwIS
L3XGBsXAwb1BDhXaFmujz+IsP+dFiatJLLXo8WCXGcy+Y3JdDfUXhR7QwcPK8KJ6
Xl9d9Fp0vfbu9k4Cj7YHeeSoFluxZbHEW+ZbF0PRHe5+XJncqnX4VUJytMVmGY5N
E+1wQR6QvUyIr4tRZDC58ONOQ0f6KGPZ7b/okjf1cdchNCBgt7hWmrGaKcUTwTX9
vm+c7SorsP8CPzZGUt2jN8YADoXo7PAR4zrE7UQ0t86ymnLVtw2dPpSRG+ynEz73
u5aViVx/SgUcRR+qzMzUjhUz8TbFAHIxzGE+AHunqUn9uLBrvCMIElUnR1Ya+nPZ
evoUZD3jNPJgSUq73m/yZiB4x02FaYvlIrI/Z1lBu3J4Pae3xO/fiuDOIYGuCkky
WvkB/dGtV2s3NECaep3NQrX5q0gJD3j4HXDJCqdofy/etiToiBnfgHpR7AdEu5m/
aryjn+tw1fXBlisIWB5urpSVSXf3dzhp4x8/L0AhUXV7OGh0q1XrPIsbObHBCtix
pvAhJYGFm4UeHvVeh0Ta/3J/XSQpcSKWBwKgZOdBuGZS4xkNvOCkBqYff6RHMq3/
eTcDYzTDjdRj+g4YM+jn06TRypMe3ovBHTSoWg/VijFLzSjQspHvt2yCIUzHzu8P
0Xi3oQoF11ceMoUJ9lt+ItwujJu0VxULBBvSfgSMrocFy6VztcE91MxEigv/9uhw
MZctmZyMzzwozIGe90zLTPIX47AlHekr91Lp1C4ERhishZRN5LgCaPVZfd3QnlQo
LjnJMNhs12mv+KBNM3bz49v6rwSeOubtxA2Jzvmu5Rh6mu37ArGYRrwmZAgCVVkJ
TtkkfRD0fE1f1J9sN4Kyq/7/OEdkstkQqJg8CwMMLVxFNzhjeHd2vZsiIqwmS5mq
pXCTNvhpZ616EzsgAIdfwHx9j7hTuh8gI6RBSpALJNAs4Ng6imcbM5SHnpoQkaPt
PboQJLwY/AValykPnYFxPJlMZfQ4902tfu8A+i4ZOH53R220fPsWYA+U9zZfdjjo
kwcX8cW+MlVAvnRJt0i36YkMzYS3ZIcVyySm8KZJdn4h8UMZ12YMUKRv/O9ZgoXv
Iz6MzoSw6z+wpx2/IOxPCVF+KhvkkGC+AW/JWTfZ8FWyDlMTCFgPPLtOzooZsQPe
yuCWSSY+Gi/1gJLWx8j47D5SOjU3pkBWwDhxISLq3Ke48yOskk5CZKRr43CtDFsC
h0t13fuY9N8h4lUUYVwWBP/gYVLRk4Y6vNaMbg4vEp7RJ6vYpG5CGCqAi3FioJ/N
kBEVR68JVEPnA3NvkkXP6MhuOnCHtQ6btoSH/xxwoSSShcJkYt0o3e4BzAsPoKP6
SpxYSIGajxsKve/XGw+BCNWcU2jBM+Ef9g5C9ifMbqrqRRlyiQGROiD3g6TQ8b7W
gKxTZElKknTblNTsqWHAuripAN1GPbrcODLKIecjgHERbRBN9uoj5iSZjQOP83aT
VMMKXpYFMHLI7oWP1Um9GDTcoFtfSkGUbt8oBehLycIWJqjrJCnYibOwnOQS4t2d
FqtGe3aP8a7YeQZmyFprO2W11Llg7c4U0sJo6IkOnS9sNe8lqKVoKxC1BSyDrhLT
mp9I3Im5CwWDCBuuYeMrr2Q/TUI+DHKa6kFf0Z31fvOSCF0l1l59NEXFfR9p9IYn
h7b3X+M6/l0L2F+9vfxiAt+STOQYxcIgGtSGdDYWD2MRUW6lwB9Yi1N/uz1Rfl/w
LPw0/lae5Up1MLZ4PmWFRC5hw0Cx9TrYO51Ki5u/r1XusKA6+TF3ujaEl/h//wa/
2iTnjgvHTMlk5EI8kdtcJk4e34qmwadb9Lp3lePEve7a5NAbY+xkHuGmvRcoirXa
ULMYWZAQ+2GHSNvLCR1BMGYOMuJQpID+Fd5X7C9uu+KFbZ4TCjdJp6brne4FKi6Y
Wj4rS5wh53LxjUOsTcm6Hi3FwLSIQXRnddYt3udBM5ecnpqokf8gYdVWulQ3gedc
4CufBtG6FxpFUWSWCZticrKvzNyh2GwgKjIbCA0SzCwGWUvFrqDFd62MAtONQuDG
hc55ptCdj15zM9qRLF6q3Fno97H799KohgG0sMc9+ckvcf6d1MVTv/Jo6crbWA7H
iAXaFvDF/zK9owqqIVHcMkk81BZ0wVEDgGdaUlfBkbeSbiC6iXSiYJ3eU3nB25F7
28vhiZAcNUe7le5Xm8zqqnk96Zvt01tl/5n4vMrRRdgDsfBT0WWDeXLGhjGfmWvu
zcnmci2+jf/doEOKCksDZuvcWb3mk+/aL/exEy6/IOHYzOgTIWjFIiov8gnrL3Ja
SxZZ14Vx7pkKjkrOgZl61YHTLpU9w+eInG+snY06PLY0mgBe+GMkYZwwCvTpV49w
pGlKOb1fPW6JMTbX3ERm4Kn54wJkdGmTq+4eJLM3ZKgLm4EuP5gRv6u6tssQwFeO
mfSSSE5oyyWrIxSLrVpSkaAkGpZN/vxDJANbs9GtXKby+If0ApRbXYRXwoSfmY7K
F5+uiLMg3yIen6mjR/nJED2S0pMBWdODoBSqWSGH4obn1jXYVIpfMkiSza5lwUgr
VR7kbvCrNeVlr60QL8RDGtICpZTdF1zAqs1w49A9zf8XsbpoQmeQceYJ2puH+uc6
d+danYWJ4BbmapLMJYEaApgSJXQdu4prUO5+y8rDlwClMxCdWqjmHuefj/dnneE3
vDFDvhWXhMB2yMOnIZ5fNB2lQCfgUj0YXSmDO1A8Yuk50Bwjmf/tQHlWnmZUk4wj
wCZdguMYVwiHfW8sClTLytDyBzklp7uoKN7htlJa9bPaPcUDc+v4+LTpG6emn/3k
hw0+zcttupIMR2dTRZUIbyE/+aZfB0IXUhBU8/zbBlmrXpliVn7GXVIVIFYiSfeo
ryISrA0o2OaaVMO7eVTz6sjhBFDeqzwq00aO8PEZoubxl5s2k95VJNzyWNQZlzen
TPgijhRWW9n7gySNn7T2gd5oOILno478/vDxRDQH+7CGcm8Gg958sk6xE0HSKR3V
T35DPKYSXqJ9qXU4nXRpg0BoXY8ivKCW1e+2UPWinX8+kTAuZ/r2KjxeweN1EfOn
tW13/g9RdfUviSSl7sZeEBEh1EmFmGsQKI/V81IQureUt2W9gZ1/SKHU9fVP7IlK
IR5bMkQ158ApzMJur+3IF+R+D9BlbH6hbiqZ3uJpIqKUvXKQQSsSPzHtSUaV4TAJ
SaPc0bRzATAgdSK/pMLjX08bHEIgaxVtZ44XNamZ+wpKx9oDCzYeaXA1YzB/Zhyz
D58FtzSbLCGCslfi+dAAUDH3SbgcvdOjm1vFL5t7qRGu1eud2PkJXQUWRjSlxcph
/uF9xpuPuXAW6z+bamBFdPkmjTxcstE0p80lFb3ip2xXx0vDSOivZE+Pqgr1D9X2
WIR3ZhWR9iamg0RZfAyXW4UkYsz1aKWrSr2p/jBvCSjyclmbFhrEWvU6fI55vmOu
lurARGFpYSC5BJmaQ+5EpHZp5sLekxckHtMUjvrzUdPhRaS67WIMFm5yu1R7dl0d
nJ1hGgYjK8aogU1WA5dRFo76UYwH+OkfC3GZ2AKqYpqvO6jjtlaT0eJiLrf3FAvE
3+3v5r69GiFPf2X0bj8SYFDY7h4waJYT0ypXHP0KBboBq+znVxhZ4d1JBmfY4ziS
77v6ar278Dg5IaOQ6Gtg+GlkJ7lntN7Z/mk5mKFP1JsOzLahGOF7f4hVl++FgJfV
Dxn1c+4iKiUgrLTj7NNOASGlL/R7XCnuPZkqr+9qza3DTgbk84k+fqQLw5hs66cC
i5oCLosDSBs00QaA+yBQYzXKUMtEWGrPVctYBrGcOG2sc6E4OlCjix4v2MTycs7G
A3leIN9fFBSw41ZAbMYz7vJW6T8KfP1ow0MZpMy8KY6gB8hFNMKX3H86A2/9M0XW
VkcZCar0xmetHkvNHINISsCOlgBhjjNjX0AitA3j6Tf5PjgOS2oXZ9lCxjFyk6so
eLLtZIliWZpVPoUQA2XG074FmsJ/UHMfolvKrcJldCviqynoa27gHE5EMg7qb/bi
/EnMpjGLT1plOQmqF0O/Fig0MgWTgy2nZ5b/3Bv8zEX3hK+BAKVg0XQAvFKtFj6D
J9hGekEUmpVPd8hMdUilqEVwYhtxeT/n0L5Bu+z55XtiWf4336MgmJ2kRaKQnMiP
syqlKJwFqcLlIaOVPc5HCOgN4lhCJAgHwv3VqVVJtahIoVE9OuyB2fgqD1gH1CWd
QW1H+a9Iezh0QVf93/s3CX3ue5CagXkZPXyzR91Tvovg2Gl7+yfssuh4pmDo7tFJ
2esO0ftlqSretUrC9rVJUjAFPKTnD+QpIARud6wLgqIl88MYJYfHMMN7uVVene3b
OwSEza2AeYGeK+PiO3qEqWPX0f5T0v74jwOMdfllboTljAzowo1FJahHquK0nff5
xZPdozwfcpUPj/e84RW4UQ40Vq/mKoliVZXeDjNN62qeHGket0M7G91B+JHDC0Iw
5YocHB+m+yhvr1x65crYDmOTeVYsPBe5WEitgSLXAC1mdNKn3vtRqdgtSVSkKDTy
sS+0M3qYkTnlKpzulguoQzjuiGgcCP8qk+fcedYnhuFpZgjOcJHDV/jjpk2WEelP
JZUP5viuJ82lfbJ8iKSl4pV7Wf6yJbMSpyfqnlh76HspfDfT0FQQ4LIO/ETQCKpJ
lClS+JP6fM8BSgUoAHlWF3AY7S5cPugTr6o9jX9wncjU7s/3PGi2HzY7rDY82Dtc
JXguJw6xXYct19aRaQJUC9zyGMajlfosPUj4TBSJoet87IfSn3YkT37xsI0UMVYu
rlUWrS0AVtrm1pzEWxt7vqjyKhpBIRaF9+3AJzauwkPRoRTnFQRnZAY83ZgvqO8K
V+ufbVcLOY5fXE/NuTMskMPZ25z4dxqi4eIcsdiZy7JcWfhTG6QVATaihdpr8zs7
w5mo0rKdO4zLvH1umLDG7REuYRp2/Bj3Qj4SWakWtIiYzWOlZh1B6Nbj6rsI08d+
SMoWfayGSlzfIRAH/UvMYmfbxHPhM0i4F+ZwVdoJ7pgnMCcCMRxnbF3w3wy1twG0
KB68Q+sKquI8MxEcAqjqwu5pWpqgjUDysTaaLkgJTgPe42fxZ1Cge3lNGTIf5NuV
EYQ2LY2AQ4BqQM6J2xoVhK4YGqkK5CgaXbK5pmWcYx1XtUF6pFXgIkErtUtfPw67
69J637DE714bhRs20XVfbp8oXuTWFeSaN9hbdxRpSOHi/sJclFP/j71n53xsUMvf
4GTnOLC3WokKvw4TfftuZzMBFfgIkpM2yw17PiYJsaUkg+cEgft0AX+xzp1g4Kao
L1wu0Xs0178RjqAYMaGACeKnRUwyoT+NSlw4hSzM8hFLVUUf7gHVhSMZHB7XuHYA
jSNbleqU5ZcTVyplI+Vfb5ou2mtWM1trsYKDGW5IORShB7FN1mazA+nJgWu/D3kr
n5xbfARndEvL7cndzqaWyfmSoVdeFpF3Mqk4++hzgqZ27Smi6+bG51XRvqsaW07X
9QAzaar4QLa5BNNo3Q+7mymGoDUiE5lO621TmxEljLfAIgkDENk3o6Ew/ODLaYu7
X7Rdj6R7YyivY2iCmb4YaknWf+u6RUvkaSbmZ6P7PjCL161cc9rB6mPePClyXI6A
gTawwiQfikM72Rhh1xK2HbnlyyEVEqD/SLqNww/Yj+CO9cUypXRwHHBYk3qD05Co
Ws7yADtuIWoYwudOxwuEhLI3rNfXWO2+U7vwKAJIVJeBYKBLsWmd7peBQ6KcGMcw
wNWenaN+2p/cAavNlGTazVbBexqUJmgPnZCdnCQixJSxvqb1KhAPxUGsC4V/KKr+
AltHtSVL+x6AMP5ssi0JOdQ96jxL/ES8Bj2Z+QJWn9Pl0ClHwsVvEeJREJ/7Jb+F
5BRUvUhMUbE9xBvg9W/WPQWClthmoeaPKkcj+MPxK5Jzx+tiDDMEB2QKMwjNpJqS
ZfwMqpxJvho4fo4wAzDChUGCt2nQpu4wK3h1IDGx1MqQ3n2Wiysff67vkaaFybez
UllnaIAmJgCreU01XBMBC8CcHD/f8NlL+vSGk3l72RYtFOyOj7A/ds0VMCGkIdnN
3hlZgh7xnVclJby1JXmrsVCA+cgwkw9UGKqJGEgt/pgBR08sID2Ewt9w7tCmSVJN
LKaHvvhF21mbooZBtUTkEgN+S/zIrd/KhwGw5TM8S0lnB5axQRpOezuA5qR9b+oQ
jmCHDtaKAgZA/TsSMRORBlCR4HAvCKDadIAEFkw1nqZr5O+AEDuWj8WABybU0U/h
Q92aQxZk6cW+GYs5T9Ih48wNNvjnmCNY6mdNVax/DxOaG7Rknt5GWBXeE6lM0sBU
QhNOYn6qgoCjRhWp3LOLAr2bfPEULQR66VBNhT1APCHV8QOvFYmq2TrPYt9DYkj1
VKuRzajoB+ZHCjMWmjXynt7xGcHescEKiAdM09tzlNYP+ZyJTsSfJVY0rgHtbDYE
ppvEGq8/9pp64ho5F+7xPZIrpJLH8DVMOKv5leKsVxHn2s22nQbUYkeUD0yvSOXJ
5aztj21GTD+zpHM6SnG48MNF4hOF+I0U0lcXgwGZ+nLcNMol5aP6JQnXjPd+onbP
vjNrGIwFZBcfjiEgTxC5EemMX7TlfwZ/pOv4PYMQYljzUHcnw4YjDQWEbSHczewR
v+xxKnHCcBH4gbUFpUHAMsntN7eWNbv9gx7Nlft/y0jQkBnwlbN0938tDrXkNneN
KP+39cc+cB9EkjbC15cP6GGWBbWLVOzIg8LcZz7mERq+1sLbMdn5t+CYJiSBrJeE
MUG0HnecPcWHy8M0zy+PZ/+eBi7EbQjkKMjKX+4CV9mqyX4H1crawQWxarWmRKDO
o124ed3ksYTjr5GTMKxanPqq32d4tY2pLjUuY08QfZxjqvcc0GkMHsc5Wiktzfgy
FzPQFYwsH+YLS3ynZTGO3559FIlp2Heu102zPwCiXVGjN+3JUR9mmIaBGHnd3rrA
5ZBUZu4mAENho/66PsSr2x8Nn0zzRyoXDctI6X3koECc7hhQWJ2pL6nmdKLzqGBe
nSj2r0DhyIrLN1efEvqVSTjn2PZguxAtABczKmg4qq7X9pAJBnGMxyPIC6PziDlw
tnu3Z+z6Fea3SrNnaNgv1D5TEBuJmgmxCeQccMO04+OeHpuGNolZiBv17or8KslU
FCgaHpvjedbRp2nRmeE9zjJpu33G9VmAo3mjR2oGPIj56vhpfEaAoI/YGUDz8uXg
1FETi6uy6JUCvU0QEpH2p8EkVpCmU7ukZj2xJTMaYGNQ/DxC0KUu/WKqhofHgLso
U0AlY5+t6QV7HGB8dll70WVTYdGCfnYjkiJWYXCloWGGS1WDOYVSbHLrLS0PhjaI
9VWXume0r+LizGM13LemW80I4FlaknxYJjDK6GMnjzu/BauPxHqChr6AFwLp5GYH
yk5kGEabCKufaaYHM3a/dRd1CteXcqU/59KrKVHvHvUV2qe2avRksTNvA+NJ6CkH
4wZMgLsYd9MTkss7YO2T1Gh4W5SFH1KuN3VCTBCdI8qxIqHwup8k3PvZ3LkwOJfN
KvLhUr6kspX7EgpeEAffSzoMcLAFg059lv1mG437Urgi1O6+Re/4Mo6ftP1vIoDi
No+yUE72yd/yIQum4i2UVD5L2FkQYkpzzaG2evun7fCW/0IXUWlf2SbjbmGE6j08
50nBiAq8THwdiYvWvvsOy66gg/ZGP0uDCsqejPnZeQL2xgFqTfotOQyjepT9QGEJ
k6/wFCY6hVhdbHpUPefmzBvJhoMpwkWZ2B39t8xj7UwBQsQtEFjQc8gt71nNZnUF
1iS1r95h1/NmpVsQX7l/SDVV8LtqkU/Cjwf0vFmmh9U7vafeJ3PvMoVW3joAJ2mT
Wc/wqoCM0BecAFyu67IBYTNn1Mv2livVDP2D/Zt/UxE7ZiGbQE5eJOmUjzcLQtxm
F7BG39xK9lUKe6kcur9SHSchjCIYRc9cYFDA15UyjsuB8QK6h0JqAWTDEJzsFVDt
SHoZT9F3mtvoOj3sGw42Q7+1BQbeC4i8qVS/aDWc24+s9tsin1c0D1F1miymH+RA
2bAm3dpxnT3RNVk55fNjFwsM+uN4KKedwhJXenqLXWUmVDXkodYGH3U1JFjtHWNZ
V0rXK1OEmyVaNFTmWHnR+S8lDzza0tBs7H5RNFGaCjUFOZQz9pKTEsT4ldkORdqB
pSjiCU3IiPhYGu8zA3D1WVB5B1rbTwVtYtDs3uGElDndZeUT3w8qX2rmwo9LClcp
qvc0ahRV5R8W38lCbqjB1e/MzHboMfs7GMbW5N38NXnCsu4irW7tqS/4A4SaM74v
yHYepoBYZ2AM5s1+31fJbJvrhskZ9vb3DmvIXUQt2te8oxaLM6bGskfGByxuh1xh
YCteEAxNknceT5YiVYU3+pkIVQRkWxgo8O7wAUbUs+c94kdNKX2Eu/a+lP3KPXDW
19NvDVVPYQvBmPLjwTNJ/eVFRtymqIMfgRsXDStrW9zXBX0BVFRlyknkGFqmPGmx
VhYPRM3h1NhkAZNyKuyfpdCF9hTQDzC3j4olqVCJOyfxpErTI7/3ocwxIjy01+JP
tJSpCAUfR/HYRiTrZmby0fQxZUmN41naKESbEO5reCyLNUIh/+c4PYJBA/hYmXqo
f9wM2Bucfj9T3+ecL/yWiWYWEqh6d6F8oSZwbrYqLUeGkVrrWbjgp7YhAtNOYA+N
CdnAWx+19tTWSEMgWxDz4VW9HWqTn4mFIKtHKyqjFCiDIbQ0D0E07O+KyAdlpZlE
hDGNMruR7SUW5TFEiSl7joP6B5Nn2C5diuiXiFwUu/W0ZsdfLb/3oV1fBPWGaU0M
fip0KYeETf56JEqT2ieWK1dgIoI2hFYZURDxEdwIKfpcOC+NnbVEIaPTgsfVGAd+
ne7WzMudSBhI8flndACIIRACHtDzhgFmIHUgJ0YLvLX2FUS+VnHtGHnr6e7CMgLn
5V6NghcqubxbdwnHKBA3owVdkiAEGPYStiGyyfQSDpXGYfG/bBhRRiMDCtUKdgOE
wIJptVrjDgFhmDUbqMzXWxiLg3s5a6t5Jk3H9z1m/xWx0ZuNU08wb/wfOAIo5q6E
2PGE9ZOxHn0Opovt2z3YaWQ2pixsPG2bhG2uGgOoT8dutwjrkocdwtkpKtaEl8NJ
FJxn0nSZ3KbeRfJbUMtXzqc4eo/hLwfYCASvvY7huBCSGm1pAbp3S0D76Erf81Gr
giLftWO4OqNEtvjm4C/1JHWbn4Kc90x9Io1u3hEvDJV7RiU+4pk8a03H1SAPrsy5
0Y8YoY5o/cHwWE1Oi2Yc/4VjQFjsesHYx2bcf882Z3/ohMNWVtxH0jgZR6u4vV0q
p2lwk2ff3KVlfzYGopOmoJzvcxlGbdRVhk7tQfKQp1X9Gw5WOx/npD5/NMRzWcPI
hA8lspczgjDSw8wsqjPwtsk3giJ+7lTAFTnivK5V3AKCtN1yxa0ERgcMc7OJpBTr
u2KQCQTzZ26jroMQ74Hy1I4ga/KJqx5u8o7RpgYNFZ47FFbNQ9i74vm651CNJwBW
RtLHtboz0/C5VBcWkHnr/RuQNhtsgs7nk73XHLXey3oZG/2akexahtlCK9tPik/0
GrF0aeUTs11Y28IHQ+ZeZQnDatDadaUGIBZ+tzbGIJ5xOSFR18vIQuuvSK3dFTCy
iDkOwYYHue4M+jCeRlZGZ52GLl272CwYJsIX7xBkA6hQn8FfC4QfY3eI3Sgg6CFf
NPILQ4Jfa7Td8NDtdSo9GlXpXf6VgjeryRyJZpJRoWeh0KKi9D6SpRZTDnW2woXc
WSfZb8F4DG7dsSgat8WnDaBd+EAjgk6lO7MYqociSfongJleIuptmgbQ8ts55WUU
LSeobyoLK9nQZ8hI0fE5hxF0+fyOPTnbpBKUgBG/qZ0VLIbytoKIp9K0OCPJYT7B
9XiaxfgaGJlSFSgZB4KrPyMLWCO0qmCQiw3l5/OukTvEtGfO2KdCFvqzMBZ5kdRm
XZg15ieljy08oZFTrny/SgWdm8lza5+z7nVONvxE3DIeiyUMRpRL7fQ5r7IcFYme
e3sy7U+HfAi2eIcuC50kiOTMCMLqCkZ2VsqE9XOKPW7+PPqlTihrDrDG84kNSLmS
t0biKL7FkXJUoqqcBeNWkha3hzd2fgNSSvcaE+RDVTn2F0Y/1jUKWZ1/hiZXZvbB
FIfW967EX7bQVhOBm5JzkV+Bept6RA+LZ1/0o4dA2jVeV3zW0KWr/nIp383mr38Y
YjcYcS/CAOdnqKM5Bh4ZpV3rkDreiqj5AH/0MUrfYcSnAPnZ5/Z7toiwW39Kuqga
LD4m7sLMrZmx1w4lW0JRvkOpt9W1SrrIEzu6NnrEEKQ0QXuwT3i3GZcCO1tBnyDs
XdWwHAOWGVcx+2aEk1rjzWPw4p4csJdSG/4t/ZR2CHEOjCNdNo/ZVZ1Cedq3IqMF
Tkj/XqUBqklfR4M9BQwNXU/FlfeORxly7a2jU4BLQ4m8eNFYHaTXh5gFrr4g5WVx
xgz9RAXgILFCsme9X3bUJtgAWJ3ghjSAseuRkiqjIRWtvzD1MNdbrwWbuoFLEiCo
4bXMsa5ceILL4Hs0ODNdQ/F2Yd2Fg3Hs9xd3Rqv6MS7xEpdCF7Dc/FlFAcdJJojA
p9afZxRkqgfUF6R7MnCiBTFRE3c7dBYARSDl5PAjFOyOU7nsSfjYHAk66vtndIlS
MvJfzecHC2hT56663Hgq/sHdwSmQFdUI4n3x58I1DgNzqtjTuL/1Fh9IIiGd9Qgz
Gxu8ik5e7zTh00wlrfARj/4UmeoU20BgLThyIzbzX0wKZCZF7gN7QT/8pZp0V6ly
+yvsD9s80tP7qcGvsEuXblnHOyAQc/F6caWZ+c/Hc4aUr7IFFefeg6t6wEqCFTrc
2AVZQZyc6iYx9TkQBFUybsqBkfQv3mwQ6ND0QxR0sNs3qv75iJjEJ3vnIGmqNCK/
d+7VSe3gzngwIUFpxOnFFF+ba2lFzFzH/agaUiaMLYMHhPf6FdCpr3x5ICl6fOWS
ZIp75Lp7hG/dqQKgLJ4AjmbuPX9wfrPpomoBvTuqfeQq5PYvekihLzc60709bOWA
96JwgHWW0cUFsklsy5yMhOuzfvF7ZY0dWXNjbK7IdLliUeGjbyq/qZtFXDlucPwT
Dma0WSM8108+B2J5S52ivVWlMUqyWeg+C79IyV4JmAogqUofPkobgO/oii9+V+9L
UU/CgBPUtJzg5XdpEaU4OSwjXsFXO3iGt/AEYw+CsO0MLidq5slno4bFvlpVKdTT
lNcm7XNj87c/h1bIcPe8m/ZadIgGcATH/eSA905Rgk39fgIiFB8MtgTpiFU2fodn
THm1Z4uyaSJl3LLSMNMOvoDfRjlVaIz2EAZSc0RfMWtmq9+uo6Lp6u4b3YdAhpLQ
9TypcRqUAalwioKiM0IKxbDQIFkBW4AHHBkMTnapfRVOxXoYUOGtXZGrO7hHCWtr
2c7PK9nXCmRkYDYFHuT3x4yCtCoZzp7jaVWP2Xldojy+7/msrgsCUHh9KYm3cAbZ
DiPDClmaI8MTGs1L9+OtCKEvwvAi7ANuRUjrriZpujf0pIQAHv5FHLwc39kdFXPQ
Ok9QUAQxkfa4aeZ2sjln6ORomvpAKOkxOepvvx8TErgtRuJiCxFU3Hw6lexojAIR
+z/QqQcDlBPwW+GVm19nlvyzwcCtJQqpMAr4NUAoNUSAMeeHghWfJ6776Zw95BR5
Wi9yvO4w+3EpJ4cUy/7s6HtQ3vSmMpLJe1rfn+UNSyMdgn/9PlWgNDFHlp6pMrf5
wXCxOkwq257+qEAztw0ZcipGggTVh78o7RiUouoLMLq8BDU6jMWhS6XKU81Pl3qJ
rkXrNpoI5QiC8xGLP+6uZbC0yfpNOQqXaE/Afv4tVlWW4ZYhnJYJL5Ere3Rhs9KO
pkRxjkAxNvej9X8zdz6cVDfyjtKZkQqXURRlaFt/0jZRf37nnSmrxjuVxljrULnS
MWgvp84QeHZMviDFB5enNrLnDhU2adpzHa+9Lyxg/qmvbcwzdtpdCZ5PI4jdAmwk
GPsGVQLh54f3+V31H6ix1Oc6qP1Wxgr9I3/X/j+1kEPprUiQs9XqUzSdYsj8HUPb
BCEhZgSATFcjs7WbIeAqqGA8zHwNR/zLzDWujuiMubtLVlSaW+TH1ha/G41Hrpe6
P/yDPkT35iKZqxv6VJrNu1yZzWthGVbFIbGVzgDNmkIhcVl+6igJY1kXft/8FpAi
HkRYGQoNyL4xJbzz4NntpQwals5abWh24pISsk/BRaRt5/33Guzy8wSqwt5xetQ/
yq73oL3px1bBMi9GpOdQA5WGvztePHdchcndY9sfFQr7TtR3PJNb0U22tsuV1Kb0
d9Ii1lvp0kZ5hEcQ8BlImJf5wZ1tL3bNMwZ9yfzUAvUjRBVEoTsuEm/aso2x8lJq
cCJ1oNlpkUWuzIC12fgRuRFU/58pxk0io6orfqyiomOYHo3Aklue2WgNJYMbOMgv
Ajiiw2ubFUmhYwL5YP3WBvd9pWMEyinegK5lxOTDVf38jXJfrhT2Wk7ic9D4Lagi
r3JqqFyMrb/+eS4005y0B1Qy1f9glJ7gEPTlfvWkHIgiwYHPSN+bpgpx3jwXWn9i
23s5Dp3B/8YzqizQ2rLHeMcCgODNLuNh2iHONg+89thvLpUWCQx2XKaIasqD+aMS
hWOEGcsHukzixfsqGOLTGkT/bPMl4sJTvhnd1RIOpX9Hdgn4CC7StrWugd/w1stD
D1TWyTb0h2M3DnUH2IgilE48LccerTn6DCXiUrc4wSTtr7QZB11nTpJ5w0Pxd/dr
V2zPdqsmNE9SdFiVSD40gXPuzQHZ5L7oADlHCKHc5k1rMC+1JrDphOk6XRedBd+T
C3E1fZ3A6OpKCQnJAEFj4p4Q9E+lQPJOCaGFOPdswMWNH97KWD4vP2hCfIkPWOU+
5M3G7KEV3NyxmDDBulDw8LZ4c6i9MT8cBw2iAOgWI24Z8Njl/mO/KgKwTrWN7J2T
KmLkPf0uz4PyWFfaINvXTYbHNZiQFVN7hcRstLDeYx/aIbjWS0QFAH8WR9J7PRGe
3WL1OCF/u5jlymGAZYF+r5N646zObMW8ZWoNYGdukV4bMHtvomrLHTdMc1/OFnuR
gL+HpajfZPrWGaj2E5EAEqIixZXw9m0Ucc86ZOH2X/c8sazE622xOi+YdRs03Xee
qS3TAQxfujWu0gVzyR9GIJwXUdta1/PnGQhtI7A3yY5PS8eno1aKLy32+n4aJodF
tnBqWUNlwBTKATbhu5vI5L1maGkhadJMzrUS2qu3gAoZb46gRXtyktKMwGYiJRes
VAD5oDN/Ta53zPcDgwKbcVPsi6mH2K10QSsLa2agAXKpc77syMa+XKeurrJjlHFX
QG+Xy8VzB0ECXXN4/NAb/9G5bZbnvnXGRlzIpUOLmVik//iY8Vc4WUCQRp7pN/66
oA9dis6YEGEUur5LhQynXPDsIhTqO6HkZ9D9YSJLgzAEfCXFzcthRTs+Poyw+tVv
m8v5xMrOedjDtryOca1KT+YROBXrda+MN54yL+v+mpzxzX+JD8cK3VpgeTmflaP0
kM2d3zXhLbeq4m+OZMho/5W0QgvTxqXrbT+PbJ48o3bBjrohweoqDlfktUfaCNQn
YeiqmUg+MWOwllZUHgkjeB64asCC3SA6prExfPpne1KmVbGYFbQ64+qNA9hfriCb
8xBVbW24RyOm311UGWzCL38pk8+HAcJI6tBlHqdsj9bmWOdqEjzqynF/qZkT4oat
anbsiIKJkgGeoWLdU0J1408YCWYca+k3M2qHx357i9KKw0yOInl6duPjKFFC3WV5
JFAjPZiFkG1R2am97AVeCFf2pVEXSnzb0/xKKXCUL109Wg83UZnXgffeuWz3T2g3
iWWq4OC6eGR1O1YiCk3ajs4PSupZiOZfjwvB/2GAoeKaVLi+HWO9YwjbNy+nePV/
eRJyKjL6vuJJGGaZEss3LrEt44shPlOkjx51Cok4rE6TteNuASWMq7olnAqmacrh
g//htLCVIg1BaPt0sGwU5Du4M/Ay+C9FtFiLEZpAL0XMOEWPMJOUHOf0W/5vIpJa
rpDT1fjvCpbgcVvJAlWCZgzXDO8rkZxY9Zc1Kbp5Lq/DJi+XyHYvBBBzks+rG+LQ
Hq+VUe1Y4Us6OJagdixDHEYcphdz7RcD67M69jR5/6LFx4a9jXuUeekN4/69SJXk
rK30gH9x7yLObZmFIpHubsQwAvxNl7H5094Iw6Q+wEUZeA8Tru4dbb1H98sJH8UM
GJYubTwMui21QOEBDxZuTOFYSC1/dYg31X6XxH/xT2fNnH62ceGj/Qjjge4WN5Ge
uZiwj9X6Yopvyfo2BKiSuMXUbMOYwSpMt4uX4j5CcAdMjx8JeudsF+d2ax4j+5VE
7jOVrAZyCCK3Bd8PXBp7d4ePOkdjix+YvzXJqHFAC+B7D54iFAQ0Hov9TtpB0ahO
ml2r9lZlPuiuH9qSkhHZ7DBbTZ19PTTGroyTtd602Hv3FPg5B2WTBpa6zjcH+PZA
dUslS1jAjx5W1HvHyYdi96wDoBgI5No2FH9ZCi9W/4te70M9BXFoYfwSTHzmrz/I
0gWQekg0zdeUVazYiCWSKLcQZu0R/g0Xvz4RhvwVk8pW0Sd92VXWoF1xQwIQxtPT
/hdQ0C0KRXhDSxEGug8a+U4PYgwD80FZNtBtEN6VCI7JZQUb5mxghCAtHpb1biO4
cC1ujRDYghPsb6Eb7Y2oCrL3BPGoevqYEmEpjPDgjTa833DHqv3sdZjy9JJZSVQU
g5+AwvDODenyJZS29kcYU495NXdGGqwoZH+LTMsFsIvtWhjNNRkSaojXas3GtYUt
ixHoVg9zb4hclnB1IymQGKAVaZXEG0v32/koHYSgCeM9op1iCfPgm1tkQpQOwyl/
bBvAsJSH00E0K0QcLbd6qFVgZ8kuyfj4E+JzVeALMxx0M9glcvoA4Q76KP8+VaLu
ZQlKoXrfDpHr1agwdNttFlwCiGtR4hBkgm4Ns1tRoE39G3jww83aOn4wHWtZ1/lY
DbVwVu9cG3GCoKfdCtkHQ2m5vN+Old2ymWnQwyY/xWcBaB0HByAx/m6AznnpPrE8
ej6WY34A5471ThPTazMIRt/Ri7cZ+yVx8zHIdie6/2O+1hoxOpSZstFucyKP2nEI
c0TNFEHmel4rjT48EhHZToCj06H1DcdayTny/J3kkAiM5HIL0QkfiF0OuErlemV6
Utt5lZReoRTqBJTEmdPA0d8OJiAqPQeHGKWQaxTnnjX1FhaF71AIBl197mU/D+3h
yt5KW2UDeIU656VOmYpUrVfg6WFcp7Zbr5aFmxvSXWOdaDaU7gU8hUF9z5Vho6bV
y6z4je6UI92V3Dn/8tB67sFau6BXIN9yyyQuW1y71+tWe43V40BWE8rTk/ktAGzb
X318lVfrCzu3gWXuQZsUSim7VVf7HecCBuBRzlUqNloALz+J1yWq7I0u0ZHw5oJY
a+I8vSKBTB4PNNjrAMGrxJfJmppkcPyDqlsuFvGCoWTzjFQKNUDLZYJIIGwr+YVo
fTAQkZaPDqP/ew3HWhJDDHYYEUh374GTPTx7SlNc4MzGL/QeJOP23RdTwOW+usWs
5fIvqN0L82kWIeCJEcK15PQ+Cfx+Ytwdqx/Ab0niEn8t/BU68aWSJPU/VDJtsUt3
gMesxsKbPZTH2R4JgPLG4wQoXJKsb/NW+sDlvfSrdJRC8xS36+N8nePA0O1UJnPZ
s3p4dizov8eqng4SkWCwjBGzg2KA8KgPU3Kk0LHnSx1UI1s72OXWW6UTMjyK1D7a
nXk8/egLv1hRIjc4s4SyYb2FnjlAfdZwkRMpOX2p41A5KgCT1GzT4L+veN6hmFXj
kltEVN0Jga8xiMx14nh7s2HjlJo5g+W7rBrVTwBn2z5rGpvukBdFoDPJI/B5U6fb
++pdQn7atiey4LCu1bjlnTlnZMFTZ6E6p7L0uL2Zl/cOn8BK8pKhRw7OdQYKpQmA
fPSnoeMz/HKHXsqk8kcT/OjH0AMfbTwfR2TnKwM5QI4P2ichB2Rxhbcv7Ak7eeS+
BIiYwQD5CpaZ0Nj2zQRGjZCKwl+65NH9eZxa2aUfXo3G0q2SN16FbAN5dQt9oger
1pyyNZXwNRyWQiJhpMJJ4S8HZfned7PVCjWnSsDQRGCRvhaIDpOWEPexrOr37QPb
nD52c5rKdMY7OgKv5mg7kz1iU1lnpWT+zgOn6IMpEmBfDISYM5VQOyRUy8MiLEjh
ZEcZ6TSMa41phioHrhHANv6UpEYVjFARX2O+5FwruGI+FOrWX6G/wTgPpzTSLnHp
05u/uQs9Jd75w+qBs8W8yi57xBi2tlxtN21au1xCeLudwefMMfr1ly9PdjV9S/l5
Jk6izIv3OrKAurz32nshfs4cHqRjX+6AF9SmgoXUIR1EAn5tooVklUc4uNw/xaA+
sAK0ClTsmFH96/z+VdkZe99M5LWURN+hPWqDX4ekQQP2Cet2oQd9rQObC0Xr3MD7
Zb+OT/Cd+DiwHeczz5LHkaalP9VrudP5kgkkR0SieEYagceHbFmX9VdotKDoetsJ
aFyVtZNqjZsrmF7mHraHNHS5UIVztYwCKh2zjE9oQHtv5odsFfTdEeWnREh02waw
YANB5TwXZtDytNcSdoa7Ugj3HItnjW5ObFW3rCalGIExy0XAWXludhiGMI5wWvYy
G9RHlsCUzPzoYWyE+kRq3a/gKk6xiHP2JuwXkLsmda2ZBW85whsuDJG2huSMkRn/
6JOOQPyeKEB3mAcqXEk5gHxXmuS5sp5yZ12tpbDhQ2kcUSksRsh/0f7L25cTiLgq
JN/huQlYOCWana+zUxRJolge/n2rT3qBca2FjlkcZDlvby/kc0SC3QRJbUPO3F/7
JC45CCaqMdpQKl+gvTkdOXKmO88iVzeh4JTShc7n0Zf4WTkWh2iF9VqPg4gmKqE1
kTTs8eeL2T+7ORfuBthj6ghBA6Swxg2019/qa3RmAqIDeKYXhQ2ye8PCk0OId7ii
gFB5K+GdLjPUTNi18qn3ypWGqYsA+Xvs3aC2mKcyXfrVPdyCSOLxE5tQ9rvttSQ7
jtmZIq8bJEuDHr0coz1T0HP6gQOqVjiDBy2UYyrimQhAEBL/fkTs4nGPLp5Kbcqm
pWdcFqOcfTGrjvG2wnmqc+piUc9qFx/EBUrJKKdSFvY2guSMQwb6RleWQ+MibZYa
BYKIqTidIIENcKWh7x1kAleKFiQUhvKYirtRflQR7j/iTcKX6RsvjxYWCbynChmb
piB6dPkZrABlQ6muC8XnxHl69SmIoZ10e5Tb0MS1+26jqh24kuhWL9KcQAVWLeLI
HPrQKnvGQxqLPeH7znx71DbYzK98r4HU1vtSlTbwN6FUDRmuiULHJnOcOOE5S3fI
VZp+G/yN+RU7/rZnGQISiNgtOsqUufmEfjuBYWXDL6Y0+1rXIiDcEUtbqQxegyqI
gynnuztQYXjaRZIduj4xHQZtm+HLRJCZl4g9pmDt7DSSvea2JrAOvoVuptrzIkDo
ACqbQo1hV63oacBlmTKcf0dSirQYEeG4mCmLDtypkpcV1L4FY+Pdwp1VBHGTXMcg
p1v6PvHYIXY0d8nyd3uzW+c2hWoVRI3KBXL05z+gCn8tI4Vby8+ggJDqNMdDEhXB
MVluF9mQ9/hHIJ2wU8ch8P+zFOMD4NiWWAw8syeZVKct3Y8VtbkNFs7hzyc7b50V
H4qAjWrRS66OuwrnCowA2dkSJ6asAL1Na5Hc9zUHbZRV+kurvUTMS8TyOIQ+8Ead
yJIxUeOXm+eQt+ZaTd87u3u1kFUZnZHVa80omFuLnTI4brdhuyjk2kGnyhvtN/SC
z/UxmGx+J9Bx2GXv6OHY+LrcArQbfmGSQQ/FIhvN4B86e7Re95gjiDaE6HTTcCOe
ftcDxp6fLaet/0uSbFRj4UuoCcx0kYHuvkvLaZIgcJ0Z37tzmc+1O+8gG7UAJdG3
iCSP3Pd7Dx81bsL4b4h4bwPoudTWZCzP8fZYUgFPwyGNSB6hcgLxSrnJp0VBrCin
09leQLAOoP5+Ifo0ZseBX5BuJwepiWzE7ahOS/nCJgGFs0vqVaCVkgI2PBOL8yx/
QDt0b6oHfZaQ/Mz8qdBm5OcotCCQM9GYPyu38DWT/pPogSqFiyszxGhFH+1vAPqQ
JwCF57mZ9VnW/2OoRBedFDGoiOsoqLFcInBikoBI51WZ0+jXrTcwaSV6gPpe4C2H
Qzsnyqn+a0TZLTboGRvAwvoS2/u6mIDkZuJfdBPClZP03+e1QrjtyCEzlPDoO4nP
xUhy3YxuNHsTe3EuXhzFI6ayiR0nIAAELbcKQjohU64AC4tNWWCzo6orYr5LK6Lq
RAVTNWLCcJpUq59iZYyHdEZQAR6kqV0gCmXSMYtAgwkjZd7KNhqosNGQ2tAGAYnl
JyzrQ28//+OCTCPf59rZ217RFrV+BOfcbIeUXHdwezwRJsMzZi5AYxze1uMuW4ef
Z2GJoLYn1tJRNoiHTkDtf1AIl/gx+K6bTa9ja5saeMOqSLUtxheodfT0Q9qgydYX
FiGcPOWvs9+NfnBwm4LsOUVkD9I4MUUGy49+kztPO3OxiXJqGTA7buRyzM9Ni7n0
vDjt+Pb26vRpFV3Ib3MC/06Ru2RZUX4gF2dJ/GCyUb9GZkYd13wt3UXOErrjl1Vw
UrOrOBP6kF6aTUrNNDt3UsOWJAZySDS3RZ4NdC1U0V/aplVG7rOdi3AszwoW5YQB
FGXDqe8u0vT4s/muar1S8DShj7v66mb9FLFS1VOKINjNZLFCsuRAFyR4/a/ej4jS
UYPtMtVjrN+z/4Oka56ZLqtq38wI2ANA0OipJYtojSqU/1okm1YEDeVAowZJydS9
zVFBGje16MPaq6vPJfI0Wwb0Lm4YGcbbjnMOIGe1Q5uKZQbuP3pEqpq+Gy0e28BA
XmQWh7l1xKXKDfl6jk1YLgHDNWUL6vt0K0C7/Ksca9UT+PY0J4eAlEFvxt6n90LT
qf9on8kP5b8cyRbYPiT0XWbsyT8Pyt8gspX4aUznu7u4zqGvTsJa4k/+IA05EnkI
NKqj2Huiz2hSB8ZZxfCQLEhzeVLECoxGDiWepi1tXcE67Z066vKgSFhYn/BRxucg
u8xjM9htabgWcWVOHEpHk6k/E6z0xsMlKS/F8nFNJzkD95czFj6OK0GlVDi/eW4G
5KO2qsEoRWASFZGb/R7k88ST1WCKRH9Jyf0ZoaUKDPbS0zwIl8yHyVD4SY6hVoZM
ljCOOlFX8PipbqH2Jk6T3R+gCGZKuJ7srlMw1cOt2QnqKPnbqYdjPRLynR0Rtrtt
jAuMt605vNMYUZI3hT9fvgtLakQ1gj4uLVQURpWEskOcJ0Tk3ND8RVTJc5KcEo3e
v9RUsJiPvGAn7ASocWGR/IOq5hwdMrOrZkylkp8BPoUvHRGpaqV+8TqzIzt+EDXf
+C4mIsRvx00VXJ4suNgAVJXBI+8MCDZbs6NoenCpwMsH0R1ADpY2HEsAd57A6uGv
1FhYcwv1MRRavK264tUZx64VvfQhunIvAop1XVfvt+PoPk/qbar+BpbdQGTiiZ0S
93xyadHzvgjwL2mEK1w50QaWX2HAyD06StjzuwJREKKwgToUndutXtkNf2vLS1z8
YWkGkb6waud2ikvwwTzpm42Z6QlSrmJh/8uQ8X9WuB2WZ2X7T/ugEv7BIrgmrGSt
3lV7ZxlHTRBYmob7Wpn1GeXkkHiOXGvSZGX7vNCCOn+inEg3Z8SFNOdWlUah/bVJ
oVJwR7WJQsqUicCLeGlec/Sv3kKHHfhfGzYOGJBvmdaQd07FBVWx7G5UYiFqk6u0
B1rrNDNbykQ+D+dfRlQFYqLcuFBCZFzGaDbmLaTGixeCqoVcHZwGEs9z6Ok1+otR
IW8Hyc5Oi4lomcJHapqfP3+CMfcvS3Ju/chUdsit0Y+guL9aWyJ8Dcg0MOvXkqD6
ijvre3keRfl3oJYYzVRcbbGtVbDaZQWWcXsURSTHR9bhqph3uc7n6tBwkQJ374mJ
9QaXQWdhlQxpjbvQasyWH6J99ZLyxrk9Z5xlGhay0frLsPbE7zV+xdMuuqewNXbB
oMApnnDL9I78LP1v3HQuwiZH98JyAgb2BuXMxSmMZVRvtHqCGT7mrmubVsedrhWC
YeeRV3FQjcl/+MXb3XXXZ9UwscIiyhpT+wKI4OTlTgUVS7sMjYwWVX5wAebZEyec
t9L0OnvMUYT0xwa+w8ETIwZIgJqoe0trJyXadMwKNkogylSQhHJpcHX+aMOE2wPl
OkIs7pru1AS9rfWHb04q27z/duVnMr91pdaxP5Gu7/dtFjG5r7g2AL0bXGRoIDGO
GmwKKq+ovFAL0UlG6L/EeSGxMhIQvW+lxmH1cEqqG+tCRtTGckJHyCOfTJvmSnc6
lnGRbEm2YIzXk7bD25rlx1ZYK61BXIjbQd+HD0ES+EL3qx4d4rbhgzI106FtmAEx
d7QK2yhW//8rDtOSlaSfHvVxlNOIUBO76fBW8MFXHVWxrEmDkn51oF/GWooeBoAs
F7wwFU0tSJsSFYpeUNMwMKi0od5IW0WLEDHGeMOD/nlFZpnW+lS4X0ImiDckeu60
5gdKOVN90eqRhYNW8BgoZ5vKa/0InJOytvmvrkrOHRljHJQDx1Wym+nABggOJvrw
AaiUg7sKjUZF9XpNLSonvLisXLIg60h0b2kvIDi19TZOnP/5d8ZVNvIM+JiH2425
f74vCp6yL2U5y0yLNVayW5wOgiwvrlAvRqMFd+zRnml4fCuPfsnuus2iGrK6gSr0
LpRjUtswv8xeheeIBUkFpuZdpNbT5fKpUYhQz2oLWGx2/C0Qc7qmGTmDpD6Ugqck
tMSyxoLmFhXL3buC0uFeOkJb4PgHjAfLli+XX62hdWz8oic5g19gKUmc8seON4GR
NzcRQ4Z1S5uGRX3BcNe69IIqsxajCYXX9BYhmmmi+agG48xAjw0P3Ey0Ck54eLbY
Ek1Btz76pDPDxVessonLww+8wgCTi2kup+c9Yzw12DGQbqL3qFtNH2y9B6Jw9v5B
MpqHuw+A9VTwoKeS1wk1KKrQhM14YhRvjVDqn3pvulNuFh1ACREPdPbQx4CZXlVh
3CTVWUeWzGac579j377L0t4JdBr8WZtiKd/25L29pX+mtYopnyCLyK/IfNQo6lLU
CyT3IY9kOEbEecTScNJGCuN/8ZzfbvDgdd2pwvlZ/6x0H45pLQdMR4tsMd/cJNTD
d77CLrahlq4t74cjVlZACJ3P4jc4ERw/kHdXYK5L1SPWp0D9Y8TCWv9vYIzJuL7D
fdKiB10uwn5SVBMx+4YjUxzsFchPzpG/s1b/sK71IceB4PmXI/Vo+QrbpJyRbnUt
uU/HL3fqFK8EXvs+FJfYri/lR3Ub61bXMSTJCNOi626PY63Rqfe5wU9dOsJtoHe5
oGZoY5c4DEN+15lYIoxdeO0Yb2/bmochB2uHAs/qbHHaBEtIVpYS5Ef96xJ4dsP7
FRgMbtWJ8il0s/K/zpCiWA+dpAsL0/sVEU/gtsnJQmJAJDRrwFIyhIbjLCszHjQf
x4DFySzqo1e1gvLnTmcL6hYEjPyCvtiLMo8r6EZ0OOxqyZzBTNOJTy4kZgFMXeQy
fHPACt3Kg1gt8Bb3fsFX6ouHM/HiysA97PgG7oqijT7KYgG6YI0duh0nL6gFkJgw
1HFSsqZEKYgLzfnbQLgNHk8EHvp7P/NRipwH/KvNkVqIp3qxscz/aXpkRt6d+z0o
4iPRm3uT7H/qZLVHLs/lsgaeliGv6CrJvKcKscmlJku0fH8J6Be98PAzeOYEyckx
1hJOaCN3SYqO81L4h86pTOevOs+pnPp0z1Qeso1A2wFBtjE4HRi8EDhWPrx/18KS
0T81YHnODOgSMcmThMrpIlWTrosbxmXk621aLTqK1ehH8kraxaiSXRfgbqv65S2h
AtuxMMHbGxbxGIj+FcmkCLqmXTxbOWDb6gSrcNhdE9XeAcvCQu4KrDv/sfqr6OXP
d9hnS4y/148TkCKfk7ME35H8Qi0Kq4HCA4UGjZRdP0K9WKrMHQm/6usLoSbwlLj1
j6OvfvR+EAYHAFP2TryIWJs3gZ3fX016atKa1PmaIB62fepWVnjI3ZN1q0U+KjOl
1AB/zL7jb9kjlUtSbvWyg4QCRn8x8hyIzgwrX+UvrG2eZRlgoMgG/XpR4vT+QlMt
UBUG5FrUyRMWH0WT59DUejsSPJdBDuFWBH6GmUaXSojCqczR3Lc8t1GDQBJdkEvs
97YUOzepkYxcrOC6budDss0lDtpg2KoJHnjqbPvpn62RUFxLT3XbAU6wJjMmttl8
80VWdG4FrLOnt9eM0DUQ5BRn28Hrr3aVXfU15luXQ0KCMVu2GP7v/BnCNXmbmTJf
+sdHXdBF63o1pVlujZ1B5v9rte79k9bYpZQA01dcXTcA4JtjZXGYOYH3Y0YSkpjb
9fIJ0//0XEL4bL3rEvNRSONJ4nlNA4kiJTmFUOf0u/DoDxTvwVDKqRte7+9TeJMq
0gWgyDrbNFK9kquxV+72zbJNFUahLUcbYFDV9an7XdAM0TjWEH7Y82nXT1shv4p8
Qiz0hh8ypUBRPrFUZLHwNcjYWBeZDliWLF893Q+YT5cP6/ji77GIUGNqeo7LQV0H
6DcPx5gZX0Uz9rmPZvJVIdewCINbnV0fJRLKacSJbTI5n0GbrdACbfJE4AmL2IcD
ZEvjpopbBHVCABT/dEYajYplGaBHzqeVrzj8Mxbl7i3yyLxgkGPWS7W4SYBrlWia
ePmZn593crPfPBQTGd1hODZrNGTsUZylKdTadjEePXVrhp0VTfjOhLMjwwBGluhe
DpwcW4++HU9QEsti0+DJE4zrk6J9vgm0S73pzsjt1cMjNmYHL3ACaxZQURzkHv7N
JMcQqqBuDJFAYYN/tOSI6E645U61ACrhbEy7QH2ntOQGgJ6llpITjCmQBouzxlGS
/I9v4fpk3iiEIrk24S4rAYh4MMNO3eK3qVdy+Qak70DNeHEPw88Uu7VF4erwmYXH
gqF5rT/Jez3eQC5j3FHQXPnKFdBCJD35I/Ky3D4y1PWQqjs49ie1Sh23lfwmsBIO
xg3VDvkuTLi+wvXA6MAV6c1AUNK7Tc+XKW29/z15ovURIv+qEepTgLgY8mlfKS1K
Vi653+zAof8aP0z86acCYzIVDHPB21VoX/fm63PdRsKcBLD9rHz7Lttrwh2eNHcs
TmBO+4p8EXNu0ulm0SEQdp5sjJaW3IOcgdq+6QI9Q+Kh5Cnb5uhUtFPYidUEOb/t
EnGM2zwFtRc6WTDLrgeOIqO63sZnrrCbJDyY2P+xyf5DkZfjut55HKjRTaEVdOCE
7dzBcExM8EVnw6btgkjKv6XsObqgTdOXG4ejYOuD010+n2f5nZEtUY0SyAxTQScS
dx4eR+jl7Jo2A0On4QVygFRlhsE4hezTWnTIhGCmBpisNSWtJvyvq+lPwzA0Qlf0
x88sYR8QCGhjzjB2GL0NI9M1ocKvcWn6qqiB/BxcEMAEuWTTYehWtKL78AZoCL8Y
lg+bWU0dAEMXNFwengUQj9eOBVo3mQEB+vL/x1gVYq6+1a3HQVSDlZZTTvsrsPVB
UVK1ZtsJz+JR1fUQyfnxY+FOT6Xj1+IzuYH2jLWaHzncTHql7rlX8pAyWdmB4355
Bew573h1dMA7LqoUsXahilciuVBOvjDb4SyJ3BO+Q18UvWW6eaamdw5cfEHiv24H
NbyVkJjx8GklMw7VfSQD6gL8KotaM5HlvInJfIO81HR8ih6n9aogZCzPDc9D4iXU
faVG/Qns8PPufGw4bR/9HiLWuTHFWwBhL1oxC78nSJ6+HvxhK7+c5cWc2Q+u4HdM
/ZIG7IRXVADOzN0X0WgdjpqJvprTDe/YwPHsFOhGM5zUBKIovNL9x7HaOkVCBxV6
yAAujJiNIbTdOGhsirHNCx9MftBKTmBBe8QwD3ZD/P6nlg2lhrlVIT6RVEbhYXbw
y30O/4rOTc/7A0evv1Tc6Co3TRUcNZglpxUkBQ8d1j+dXiwtTIZBruSvYa5aGLUq
7rvpp+NqVGhAftcJhN+a0zPji9P1efpNsykwMlCLOUsEwqsvn3O+gUkhzyqs23AL
VymXEz8mIr1mbZsZx7JNnrnHvaVh915390VsGhLWyCGj0Z2yMmMveQvP9nXrGQna
CugzPv42a+XM8S6gEiQJJ51ru05leUh1knbFJIF0pdjUOhh82iIO+WLbZ1Ju2IoX
1b9KBQxtJMexTu7VtlO3zSlEVdPZiZfG9P4wx0SKpauJvgkejmf7PFiy7JPy10x8
tLyk6BjSqKoN3UMUi6d2sMTxZNP4P2avDvae8tARtwatN0U+tzUOWJ4A3p4zwdGb
9HDt8o+r7vzcKS17K4LzMr6LAJdIsKVh7ZI6y6bv2ayaseoQ+OCD8NlEgdd5zPjN
wbSOH9ZrSM9B5krZpYUUOvZcI7+G9XWlLlMTJZAYDujOoea7MVt0xx57vn64FaZA
F2hjZSYvvfLTsYIc//ThL54RATZuj3hn4wrWM4SzxTekIbE9WGDEvRUEFoTLqRQe
8iKVlqRhLk23VjmJXXtgI5kj/JHFeiMG1wH17OQOUaXhxrp3P9oUOsFG/SAnN5Fc
Da65fTFCX8jVMAXHQtkDxSXoH6lA+T8aPcSl8ab4H8fGEMf/arQVIk4vmzKAoaRx
JoDHWQKmU/jP4Snv4+KnABAitINdzrz69ykXtnmqkLP30wSYza8HaUxCGCSx9xDh
1kz4XUHoqTZM8cFJlMlHVB9Qq++41bY0Cdf0EKKIVKckFMrCJZtW1/3XgXwAkfgG
iXx//gqJSlNG0m6XtLgsY42jXWKwR91KE9dgw3c6fZjZq968mBgk5bM8IGfwu/0+
+46xJamzMf89OFoBHJtiX43ZRuHcV4e3R7gPxmfQTlzseCnE/H/4AMD6D2gJFp1q
JD9Ue9krYx8hmw7Sd1c2fKReNWqUYC6Io9eVyrUdtDoZAuzWLCNvz0LKqFSCXjDN
zX4ayBkM0KXzUm7SizWrHx81RLJz83gTXiEOvjn26kc6IvEEoojzRC20WnCNiN+Y
AsDXMyiCN7LftQrH0jDRywL36APDOlcFPfgbEFDyXyYsjIKspOxoP1lO/ueycv8b
Y7Z8mqAOIBLZWSjaUg2NPCr6tm+v0/WSXwCBzA+uMuAIjqHWEU4Ua4yhDL20iXhS
DqFgGMiSrsnMot0WC+EcT3mHvurh/nUG4iz5VsLkgKMZVba4rgGovYZgFyZwXsbd
ZPUDYTiG6lhtThfD8ANSaUXqsnDFwh4IQ6JhOhdfIty4/Aqp/eXF+Jhnp7spwDLK
+RaZte04OK4tmZtCxGfhJVJ7LD2dxNY9b2S1R/8g/6zuSy1wJxLsgZ1jDrS+sExS
+0+Fb+kFYW4tOnDPlPy24OciHjte9TMy/Qh8KSw2vraMzLMslYqXj08/EWPkJzsp
2GoERXLKnigjC6/HqB9FjdlY1tDuFkq8l7S8J4sRNq8URlNnqk0ItORzu0/LsmTM
+/GJTVkWyRMZ+phSkLxX3zJozv9Qj55vl8gS69u+EkfQLE8aJE0dmrRhVs0T9oXB
g9YoHyMQt/1FeI094qB0Nx6O1KZwWgpFnnwJs+S1pns72rq3hyvrtK0Aprfw0v+/
8jaOzkocVybZyH60nOf5QNeRnCAXUPBTXGKAKUtZhzb7KhwP4hu3JNCHjbWiNyQP
KSHUUKY/E/S1D5M2yeM4aO8YL1IVKPNcP+18+1JOhEGmLvPq6uxoHPD1t4feilCY
CsMOLHI1EL/4Gwb0W5e2hw2Q+q2zW3UujZ5vE1bZuJNptedYm/Gb++oFbLKFFaNe
rW+RlkyhYqfNKfkYybViB2GUaK1YTBO3yzQbxYAAZrM55lyhzPK4ZdiNZdqTalbF
zQWRF0GV3chneh2iisye0/mbuQKbYxe+i9LgmCB2Ru0PkmajdTm7y3jCdyKaeU+0
+nUkZNxMfwCkSrBmeuHcxYaNd/RET94dPTaX60dWZKqwA1V2sPTeWx++PPfw2Q61
/faK7Pxq5liIhpiqavPcIYKEi9WBgp4ueD31/IZ4cBwceB/OVsahk3opatmpmiEW
x3EtQp1Tg+m8Df/R445UAVFW0gymKWhOag9VqexbTPrxtyuYj3r8V/AXNoAlJzeG
IpfUcVzNqXLJGUoy5aFUlVXo+RqCkF75laDfvIpgE8jHYDeISCNxsCVZyJJfW/kc
ZOoKnFI01p23ybmR3KYjrnKT13yM22+pipIr9MQZxXRvQqkLLk/TIAN5i5hOmEf6
vcFLN/QlMVlXRodbwBNzKgOD4alH3s3CwLF/RRj6Dfgf5sKkNEtezhJ89DzhkuWa
TjyijlesZYH/plgz5muRfCz8JUuI8S5IBARqmN8gnDR3KvWRJPx336UUI8bpAIKb
LHg4IUmaBVzHEfyCiM9FWwHd2E1IKgmuI1BRTtG2SRgtMIlB9DWc49QhyOFj1hzz
vkjINvSQaQhnm/lmIWYA9mfWm+2I5GVaEu4rKrL/ODGz/pcL0TCMaA1RAMJPu0uX
jvbPz6o3iBLzm07Sb1cFOkt45tNKHyUkD9QfiqbrN4eNH6jiWQa0o84PHNKEfGeV
M8xLNUISPFhah3dqRL2WHlSrSBfGs2sJtBHgP7brbbAsX0L6t/sZ5e/Fvd3soKhi
RQrRFb/ZrHerDS2uBNeTVvkpsiW0AQcV1BDFQfSk+NsPU4+CIxR7Y/QQgFLyvJNy
am+g+IHWC1bBZ2gB3AgV9DHhbAzylvZDnP5z8/DwNpudprcBsWJ40RrgylnhCSu7
fqpKr6vcispE0MLQL6wcFQxpNZv682xhooi2WnQJzyOIoTK3yD33AH0MpPicGepZ
u0sChVyvKEMlVfz+PVy/yfBAkvBfFmIBndpgfbVDDgJBdhT9xCKSEmtEiJQGHEjl
j1Hwqhmsylv+aOptrsWYqBVdOdtzibY2coHGoRMuS3El3B/+myXx7yaCbW9hzi0w
GyDoHnhenRxWzvMKMfxiKZPBCkxmJ5QAZrxXi9oD19lhPs1S8gXFcmnHFa9D7voR
8zftkAbgPhC8erCBzXT+KFfVn5baLmBYLcWsqdKGyz1PZ5i8wgJ+7usg0YKeJvCj
9eSdazQI7iiFihsi5/e9vZS/ZPpiu1j5F+ReTEB3Xp7oudjTFLmUNEa7TS2xdptu
Vi2vJ4lggb2sOUyNc4j1hQtpCRQvu5RDbSN7XLaQXxDFsFABupkf6oQ4/hnphNxG
MDrcfrG9MBSq3DYYKvyNm61salJI3ge+W+7VGKH4/2y7J6mFcM7a3lUc3jZ5mkcu
iZhZI+8KBh1+O6pFJultOYigpyrh3kbk69ILNX5+N8j3pPUREIP5eqaDCemUIni+
tHTOhPvSs/Z8VelFpSLHA+wk7/lj0t/Dby7ItKrzGqJ9OpyTTEdaTJGsDdIX5994
kCBU1y4FBCan0QhB1jsNu0RwFTiDs0OuhfGugF1wP7TudNpyv9hoajVpk2UaIUW1
tyLHN2B+wJRfLGtnmI/fKkiUOn1cfy6cJM/xb+5Pl/zOv0oUzNBqbB7af2dwA3fu
1GgxI2sHcEUQ6wY4IybLmuXwYpPZ+kH5idOsx18vBZ9ytmrDFq04chtYVSj+Wy2/
MOuUOHkBjO5e3ZU7CvmpSE/EGyEwN6OcN0t3m7w670j9hW1XT3kXyzEhcUXMu5yn
YzZ5Kk1WWZAoOz832XJHtMA2nYuo/bRqt61mZOTa7pJEXbRVm0rpxVmbixrwutGD
aJKjps1AtcXNK5MvRhgmkYNoM7KlNrC3aI2Sj/sG7ucD5N79wOEt5xEqHsj9w2mR
p2wezRAofYYAfYJMA38QMjJjn19zILAzME9WfydvzYJf5WDLjze++04zbIXnV3P3
lf6uN1j+GI1IJM9LpK03Wn73ej1Kwbmhx+IdJNQPti/1Mn35J1oQvzDUeQqQvDdc
6TwrAoUMCASPeTcoSKfqVL0FUi4eixXq73LBYolGRPWkXoGggk5qgQI5OhZlmPuM
iHdfccT2EOgdV7N9r3g54q9Hfk1kG8tGyMyH5a5+GqGfERa6T3L18FsLrb8Fbr6l
/OSVMKwfL3ZmLN+FPIbSejmaMQWKnFNqRhfDnFp8jdr12tyG6K+1M3H/i9vhtM0o
xF/79hgw2oyCEI3SoToRwKX1YC+vXZwD3L0osq60A73zGwy7UBHUwGGvn0E5T/EG
9qZZjLQuynCwjRHQtTvULoUnkVf+R6CqRwMHNtGxHFR17/cnJNIBcL8LDWsFmHP/
Jfe8pfXRZqJWpVD8HuFYV0vTLfVUGxVrbYn+uVp05g22wMHuxJv9/cOhtOBc0EoO
ur0oSNm9lywvtehR/Zcm8tqWVE7WY0Fhi03h4KHT6668enkYXAVSvFUeGGzKYuZa
iY8kCVbyGvrRNt0Ts1kwfD1wY+xl+VntvynEJRCGZyBFJ9mzz8iffdaVfwZ7eo8h
eHXC6L3uGN6VLTAGbA1Bfgo9ldAxf0XEYoChNLxAcvzuc/d/i+6hZNhrPxs8EQNQ
6/iSHwYd1IDfp8Oc2Pgeq5R7g8aiYu8NyAHgOoYpO6W1pA5R4Nh7qBrhFPuBULIp
6UVMmiFn+1gQjYGQDIitZz+cr+Vqs6kvojmW4Gn0tdvD+CMJPo1x62FHhLN5MzLq
V5T5wu7GRJ6Pmo32ENAqLhKRihdUihGVsZcugTVg+nr3MomRgmWKgnCAjyRFjCG8
GItJZWUMFea3ZKiLBPXYR3IjagSmAM8H7BiQURn4YJQa9utGY2DSPa5ENr0ShUUy
3+XqKevz4iWTYioxBLojGkY3Em75fAiXgE92s/8A6l/wQQs5XhiZOzFGYo+7csB2
zIhLffSX2mrI8wvCQhtjUHKpXmR0aoC0SmlzgSCUv5iUU56EAdCP8myyoyZAy26l
ZKNgTLaUJJ7vP/HP+eIEhCNIZievx6aUefMPd2wOGAjbD8PoNTmSc0K9qcCrfp9e
bdUGdGQqsIO61pZ8tEVmWrl/pvgaSCMDdHflSXr2LBpzmOLpcczm3/N9xIxIWIXA
Ut3dxuq4RQTxJ6VhhXZCN6Lvpe7U5OsGnaBqbzCiuXRwHyGtkUGo7xJruB4LC0eA
5+wYgFn3BFu9pVKm/cVLpaisgr09CM386nHVjHpnQuN2O4Is5bDM7a+dX8wDTBFH
h/nQKTtMbyaNHXw3D6F8pZo10APyh67zIirC6IZex86fc8IzgpMWZ48mRFOtyBFT
SbWwi6xuNA+YaEQaE8AKOwtt5R5bFf95itcZ+fsFPD+xzcLRGN6NT0bYlrv/EfF8
uxC1KOHBIh7S7EOwYbQx61ji3faKcL1qA70IrPaCZCt5a4bLomWWnIaT2O4IABNZ
b9TOgdPgv0xb02DV1VzFP0clsBwc/PYq57YR3Ltg3A7L5HLUf7JZkPi3n98x7gW8
bYopbn9jH/yKCBw8WxOKZZM3vNP/voHGSIZMLngJxC6RKd22FXhVPjMUiQzCLVzs
2nzcD8+J5WAM20yxQKbqVYgRk9v5YjT3qyqofwv/x9/eIAlBMyxDvFf5gGf0sFa2
OZbgUV6+FVTgxzlBnSv1t0kEi/CsEbT8OZ1iejKRnkL2OfkZRjNBpfwc10pZeK9A
LnniKtTPY2jsRPnbdt175FosZZMz1hw30dFfYOvQaFqAiKheeoMIV+cW7hYelWwS
a/wlPxUCwTj7lw/YVmbM79qzd8c62nZ3Vq82PjK6IsTlRrWYZWgscoJRFQJZ7xdC
/D+QPlIGFnPMhAyPTQ+OPxVOutAbuxZJW7xZENNEJxZn3WwiHzFGxS1FKl+OTrFa
TwnWIR+baG7YViqePw3zUD0Th7Dm1rsCsPuU37EHhgOeEfyzcipD1w6MeJaWBqQT
/HMBVzSOr6iXCyoXDcLB+pVY90eAf7TbjYCDT9f6mIBX3FY4qUWTdsS2nAcEB28X
a8EsY2reY2bMkKYznn0bOi0I2q/ExKqp8VVhbGYaFEWmhI7hPWVXawCTCf4wkzNb
jWI6z4MsJizh6qy5FA2bSJt8+3at22uoIQL/gHJvxpfJxBVl+wucLW66uwEl5tcs
SPmn8+OwEqiQQlO38dQvqYy6UlPJ4xb69r6hKcjgE9qGYCrOoW8k6sl1lemKcoaK
ezRyrkI3YUCq7Zgi3Vrept6402qXUYami6XfDcLhd1M1G9NgZgshz2cFXm7GICm2
HR/yyJrBQaI2xSMxW01JHQnkcz0Fm6WIJcjc896ri+mbyWCzxpyujJX5yoimT2oZ
GpCpjh3iUOyqFXGtXQsquYbghdDRUvGPSpfWuNEv6aur/iW0k+yVwsxT/EYCaoNe
KNm9zx8mW/w83CwKhO72uDlR8LjXZWF3/XXAPDRyI5vxde5vzGTrMoIbb1C0BVa/
6suKgK0sMPu7QUUEiAoWVYmUeUGt2HCWXpWsmBUUoxTjhYFwxBSu55j2OLH5uvFI
MgpUpbcvB+HzCZBQ/JsnpEiyJiEgeta0Hwf19SysyZWVJKfxeU+4D52xjsshBKc+
Me+VteBGIKUw5UCWJxdWOpnDYPDeNrnR9/4LEjni5Xy/8x3rd8MNDZrF1hsVdp29
KEpyZGnP1yXcmuFybZrn0dTjiyX1uPfx+gawSVqCInFQEXkOfB7SoCuG6A8IDRxB
KHID6vG/SKJ87YL1B5UjvMbfdVow+JetnnVa29U4Ms/aHqU1WdLJZQ0SnGFNZh4v
XWJIcO8WSSe9jg4291jjgipnGc96AHWGus8r0zLQFB3Yl5xqokv/ImJpY2AjAM1K
r63v3Q7lIHqZroOIheIgnToAI03Uk1GeL1PxK7FF3CQM45XwmlEeqcctbPLYYvgp
pKEv6qjeZ6poOn/CgGQzq9gVLDWMcEL2+Cj+2syz1+HP9cWO70puExGLLbOH20Wn
OF1/0rfkHWg+VIEDScoZ6iX1FtBe1z+JvM5SwYetudvxwcbU79tXg0c42CNVNC09
RnJOEFEljRs4+9Qh0O2L9INMxMMchUeMcftnXZOaBr5sAclYrnGzZiAp8xGHbnUU
JJbh0OprroIcqXgU5S7mR5qGpXaD25mG5h0F0urDX2TwhTJY044TpxOvTmprm2sL
KP4a7oOdITGY7DfDdFhGTBvUfaccA5lXlmTpFZ0+m1fIpu1hwHPnWt5r7Qwh+VTW
NDUWB6CsUa7M+EPqnA6ViwWWR1bsPDHmDfb0p75dZ8MpNh7+En5sbpEUGzU+HNDU
GnIvbtzv2MTmLDZw9qiDChEsMhJvtAgoXo1O7LSMOV7Z5vunAR3Zw+crd3HzOkni
9igx9QC2/2AU/HVrK/kHgq8e9l7QxeVg/n7MIX/+913/ACysSvOR29RzHfVb6z5c
GE9pVM2DYP35EoUxE/8hJzxrIq1xjkr12yf2RVVT4X5zE3kjnROFddpTHAgJrV8s
cjTpwjNvKLhxp2D6fYN1xcmgTtiHWX+CPkvPQHgrmRVHJM0TgaujGiD8Ur2fCi7U
8nPfC2uXIfO71n1dULeB0XQx3fVTSJ9bltSsKdxYKZPEhGVP1zhYsXhQDbz/HuDB
H87ICAaHKTSUQgC06eJF+OLph4u8VIwVD3rqUqKe3MAJef3Yzvm/7XigrHtYy4e0
SUn2vcMeldg4VsrSF/ce6mYfJjJlMhvLV9GPG0HunxjHf4VFkQAS2T1L2w4nXriY
dA7pBfU3pWZ5L0Kn9v01gu0hSvz0YHhbhCiOob6zZg8HKnIS4uF/Hxi8u38HjjWJ
/4QpTvdk6ABIyfH5nfU9QYSqTDbNgmRsW0UVkWVeztyt0XNmJP+3V9V4mbQFUdH+
eIsY3Sz7ASDTz1xC8Di62yXGn/C/tFL2UBNBSXkrMAdsokt7QraKuUjqyojBDsIJ
l/cbbMykS92zXMn6ax3mNbgRW9FzciwDkCDQQad9C+gabjBmcfsnfVOkUNQ5wi9f
+mN3/vvSRhdnCOj1820HZvo6P8yj5GaFvYpQ4OHmeM5ivTUdortxTpPUGox2SpGO
oejMWw0HKgsprvB0nNAr1xXHtkKg3yUY+7SSlDpcIAuAhgwISmSeSZvq8YaNqnDv
wyk6Cyos5VgBYKthSet4vfjs1Iu49OVXaEbrZuma1WF95tyArqdtFlCpMe+iDwhv
lnE756P7tv6P+xtIq5XZ7rV6H9bnPe9K+I57ZF/QcUr45o9rU7yJWXbyFid7OM7l
/zA6SjNgFmN2x0BVzB33Aj/qZ7xzdVXuUD96uLNea5b1jJ4kj+tx2C5C7H/JQQ05
Z5BR1eZCNOR5wd9TZzJ7iB/BVnt51dyG9xn1B6CSM04/XQt/yYThhNKqbETI+Ae4
2l4qOiKiwwKyoVtmBf2qDQxU38/rcovMMzanRAhoHbWd/IEValdcI/pOjKEvuYmo
qpsOKaUhZY3B6ETBOS84WkjK533OqaCpBIXXLbPByo7OEhkEhzaBakgL4VGanrFO
FHg5PzlWjtDnNNW0Xax2KXNtAE2F3QQyToJdAXyHu+wiOd/FZ/U9YVnCVZIklbuA
HjSRVyErAmgRJS8ks8zXGdUpFXV+PLyDcI3W5dCrQCVogYT7pitjw3LXxX1J5v7/
hqvGt9fUs0zyN4xmaECB7I0h3rQXHyx4/4QC9f/FCAtodkchOnM2YCIvImmOnvuR
7U09txRz+9ZYtGk7JIzeLlGxkypUvHi7nR3l/IYChF7Rm/Ag6wbXjwjz86wivG4d
hUhUZh4aFlE4QQmm/lZYitCED8Ad45qlTdsT88UHtF6SyobX1xMRnt+mQ2EFy1TV
uA1K3+Wmvr0WE7UCF8dkPI4eh3ja2AO4AFRnvhBfYhw5aKTIBodCwaFGSKnFhI2L
v3pdGNM1OUwD+iMqFD6YFV3y/lGlEexU4w3MlIhUfiht4uSI4Qht+1RR6DuS/h7E
2V8byoffeK0xwLVpPvlbEw9867hkvqHYlz3ngntyCZDW0ZMvv14L170mW+wGuayD
vrel0+mun9sTi/lvGeHf4aQ4EQrr0VqgGUUyjT3GBjk8sZkh0cOArGOH+fR0fkf+
kSxuCyekYWeGeAWUorCnYTeUQRD9eDOLnN5g/Bgo/KCoWQa8gwsFgoYnCu5DHsCP
eNnBO/vy6Z9h4+0g+8NvX66V/wGHcNli7ks6l9tRsaOBZIqxA5y166jzoRyXbx1W
PsL4LXbHo5Tw+LBwUdOKwsUhtF4EY/2G/mxTcgsm7g6LzLvccxdyvMDSkjIy0G0Y
FseWhAnbiSId4ok/kSmdQ2cpJIjD/p3Wj01XuEA40NhKtii1cEJfmFNsgvcppVzd
UtnlMzEl2q3Jfpl08Cit+XCX2UZf1FScvlrH+L7mgijpgkopUnkS/DNuPCqXiL8/
35ouAitKXLvZ33/M9luQQqUEoDfa1tD77Q+nI+uy0TAFUdJghtC+NpqXorlBJoEI
8gtxOKeGZj1x7HW1XOs2tF0NIoGRBNu0watok9xd5lnM0fKgxCi8IJici4fiBLLA
g9H7x5lkUCR5ncqSHhYZ3QLxNLEiXa7wjvcWlBF20zwx17QBRg/IfDE4/nDq8Va8
aCpqPu8VVMMCBFiJMVPUvU/8D19hI5Vx7m+3WBXuddwVcyj54lBPhRs7kV4a97v/
rpwSZmKk7MaCxzG4V/VboDoAxz8etxT0dPz1ynO1EcY4EFTWUhfTX1C/So1isHDU
S+XjzgjEEpPB1UTZakm7rqYotS84+Fo/G878nAvL1lNhagZBS4LAouGnyNLOZzJJ
nPlZeuOhcF4Uyx4G06i8uqhm5ccet5rZkvnuRwCZT/dMOgR+1m2hErwYAulYv0M4
f/ausRj+3UgwHTErotZ+OvxcDPdntbX+tLm394QcD0Zv7UUiLAYwFyxxhdz94DEP
5iRnonYig+YzaliQlHicXPINyYInmZefWg9TptT8k6+9rKWinNp4rwzvvbm7hMU5
nLlaya7jtbhhLkrxO7EyHfpRu+IroSklFieXYvzakdzRAFktmtXSJQVLCNmkqeT0
F9f3NeLgTM+RLTBJHU5VkT3T6gWLp1UjP8ub+jzj8eO+bwS0n/QczdToQo+T/y+K
ILPUkLR8uB8n+BYigTeVK3Op5fUccWvqUH0Q1A9PLUfkO/saZhIbY/UYJYI/MN7d
mhaTMEZPAujgBigfI5QedykT0CEWwzcWJ3RWQAHKU97f0xHozYG85yW8dDyoDMHQ
k8ZtPLQ7TWLotDAdA+LQ4buB+cCE/XDWiDTeDrdZORlP4RQnwrvVB94UiuK1snm8
6dNSfuJNAbvyaFTaVfD/Khng6joAW3pvxnhIz1fA6SlJ45tiCl5bzgXQW4kdLOZ9
+Q9xMcg1rfbnDXTq8S+eL2Q4BzHEQrqjXw49nfrJBYV5SDLJwRmd7VSpsV/M2pl3
9pCdLtvj9R8+gJmAkTWknmTESsh6tR+TRXurqBR65Ok9qFsS7zbVbIMpxvInB9AC
SV1vktTRaSbtLBzAaK/kKNjCZc5Hrr9ShqYLtk/lwmBLuoDxtbl8u86NiO8IFlz+
Xxjc7WOM9cmgdRmR6+1XFkeSP2z/+fbGKxCwBsk2RDnzJ9wdk/DvIRPZr7Bf3Sgp
58NYwSWoLq4LlFXGXw9tQclufFATWY+5iQI6yiBJ9axVIxmPFpemSm1/t/slmN3u
qLrDx1ohUfbIcSmo8FKyin3szr58D27peHDlttNGvaew/FbpTvPMRhXKGzrKUkEv
TMXFRv0Zn+ajXAj242lIwgr5YzE6+15h26uzJPR586Qcesry40gziAie6k/slNUU
upbErOv9Y83UnI+szWkpOU4qAPecwvrcgj2YNwTDS+Qi4LC7VgMLuWaB0u7RTGRj
PskUF+C56feEDflYXr4n2wV5FdEowoX9E2cz1SCHlwBY88RVuevFMCUU2Q/AF9hy
ok/A4jed1dfcIXXP9nCHYCxjZMUYeiYHEl5d/1Y3vKLPOmGZp5EcRvC0pSlNXHis
kHelxlSZovjYGGT8Nk731sop7/QXpSytgiTOEvKftbFvbPz9aICSf10CunFqlic7
OcKOgV5jWB+Hr2CUUYwNSu1wwhBBZuT2LXZ/VmA0AYGL4p1TkVEPO75+3S2LM9k5
0cDCeGyElua8T/G3GOLAQCJaklpc2ivl2mJGoPR344VJmb/K2ZSdbPsQAjbroKVl
XFbi/OeKwoVRAoOFFUOgQ9OmgzHZwM+eK9X9ocM9CTL1x5wVPQ7nKbFI8Fwq686h
fXEJP7aZ4xlajPQ1fszbX0/gvDmVH+vA+V8v9VELm2PRPwEB0t6QtZ7gJDVcqtic
UeQOI6qfKbA+72Yjxb4XZvlWqvxgy3Bhaaykh0Xe4vMhCcRcrCBKNNEBqFo4TYu6
hgDsoq7Isoe6GPYE5SUf/aoIAtFadjCGGOCeQ4zzjkFiHvKHBqmS8HpjYWdma1r9
brXeveaPQk2C4ijWy4p3OzG78BhdAAagY1ewqamGWi6dbNlCsfDaX2sl1tF/bI9U
060PHwTUYt8ch62DxfTYevls4gzuxcMKtcbIlyqk66G4M85qprwaQzasa9oRfavF
wO/itN4c9vaaXwLDrN3G7f4/dxUBtZihBnlYBFQ/b3GcJaATW7tp2Kv6LB0TRA0N
FRjz2KvTgIwzJOFZ1WHtNAYno/dCG3A5GWpmH82rD2NvSnXAf6UndS/MQX9UX500
L4Cg4tIFihRxl/G4xAzQ83T7DQEZh5y5obLoVNkIIK2PP+ScKSpwXd0suLxEo64F
36BzlR8w7myEjMqV8byW+bpKD1EEiRB4mYhIZnX0hZcIDqxLXxhXmBkt4IPJ228n
Jt4dN7BRlVvc3/7ZK/cHZU/0kALMAmKf5eHZjqAM0mmgzmBMRchOzvmY23+nLxpB
sFJYxZgyJTTfunbmlt/qLkuEWl+oJq1gZTNXTZQJgsEfAI3IueXBwHPJlRf0yqt4
jxMwY5TVpVbqbEmgzIwoZJ6RGU+QB+x5wUWyeYpkGQ3x2Ivpg4lRDmUgaj6L1gAE
gL3ZP/3uH2Q7d0+DHFlggcurrENTsTiDq9HR+sf4l0/fPOxbV2zXIFEbpIsq+7F6
9m8qnL9DPW3mksxKlGr7W0nMl4B0kkjnIPKInTJpsfY3+4uxE7TRVUregTqDKaVD
0LaWwdB410zaN1K4LNUzP58Nsikvmc3K+N8B7gHTfLUO7QmdEE3ct4CBwS9mFcVa
+ibo0lZNjV4frgajo8fYu+tU7pI+JrqUhNL4zsoCEwY8kc6YaaP0J4vypzIeklU2
RXS5GwYC6mtAMXsbAPUPxtxTR7RrkoKYOE1f2BwCcsj1PknB3u4wK4FN6a1avMWv
8kf7lPvza6jo9VEXIE9oKiqMOO51BHWlSCMWthbu4vTqLCddXLMypD4Iw9wuMkus
DBIG9cy4QBLRCrZFLV5PVHHguHFVkJBEknRd0uKbStOSbym1NTVauOG//5XiAL3u
5Vo989AC8jnjt464G0oiGlTDK5qvFVAng7zF/d9DFtH1XmH5bZikqMIvisG3ZV3K
KqY0orqtadQ5dTVRw0wL4BRVf0cSgqDyj2UlV2bkhp5DGVRmLRKTAszc4UOp/QlN
qxy4SH55kwO8Pzgdz6GfWNGE9hkoGk3IdpUcEqyZigeb5N5Wd+Yj1tKZqIvBwp+F
aChqHURHzZfNrGzZQWUGjrrrEIr1nfmGGb2V5IRiRneHUpRe8Dnt92tv/J5cwyZ/
nZASEwgX1AnposNJPXVaYr83Zgib3VfNoi5Vs6mmIwTToQBAlr8TnFrEPwJDttXA
BUe3JEFRQ8m0Qp4gJ+61Oug3iU0pbAi8jKJ+FKnpFjFL5TZ6a0H9pWBSe7aeEdCg
kqWvfr66FO1+94SbQYhJ6u10nLCHhqhSp1+9S2/DKfpaqdZkPZ8+xCHuoLG9e0Gm
S04bp/oVXukoCCKQ01iW/J0sGnRLfxMbiG6u4rIhj2K1X7pnMOCp6uOt8YIpbFez
wxelROd3OxfoI8GvidUXpdxLWYVHbvM+lKVuCeMlrlDNFYjcRQac1IwvtGeOvYzP
NzEKXZxRO1DTeNF3Q9O4JSIeRe8TpISODCDARnGvUgrkqhKKbxhtRIGLmKDtbrPZ
IW45LSPrqOEjNv2/Cj54dWnfANU8LO+5SdF5eraPOoYqlVLlGGloQM1LWvKE3EIi
3J0+z6tS4isOlvrXukD9TLoOmCFO2yDAd5wKhuYgbu6tNN8+lOXuHSvmiQGt9bf/
sL4GO6iCHBUS8SywfhV0BVjnxTd75f1vWWdhY1CZEbuGc//DCm0nJQ8f/LNUV8XH
2iwkpIPZsdS85HLFEZPHp61PSG5FP9d5JlVsQpsGi1j2PEL18PGLCw9bk80n6LoU
WHiQ3L8R/2yNzR2fbv2fqACLMYBifubVcqsMdgNbbL8yPMJ5YoG/gApqq5wRzInl
U0dC0hFSqXaAStjslIgOX3DeiSi+SRC6Os3dFv8cFstZGXwnLQS8LBX7EwBSUpVm
Ht9NftqVtJprcOHyz7DMXWBGHQy5c6/AICe3F0EhRxUabPbsEYMkFsmvU5UDJMFV
PbK6IhRMAVreHvz1B7ytODA3PlVccT5RJ4XeWqUR0gEWInshjA5xbtIRSdxxk9R2
bS6eZ6HWgXmTGP8cT1Ma9PM7mG/fz+W2w5fY9qn5KpyjsO/y6+noqSxDBipxYaRx
tHO21kkdBkUPEhzkkaeH2N7nETksI/yYaxIdnwYa84vqDFXdd2hJ8iqM1iPZAdNy
Y4PbVYgVwHhhdnzJ8rbD/zoVEKQPCpTvkUKy4leTtrwAhxYlHjqSkgv07AtTPuqr
cUlWLn69uyUUnxOcVb5QMgytZNdqnthov3dfI2laPxN9a5qN8SpZq6fA94g7e5/6
UOPIWSc0QeA3LKYcba0f6XaAkALpalfIkxJSB9+zdagwgYiqvtrlQo4/cUP0iS27
V8+BZv1/FH2wgbs7oEEJOOA0D4M8B6XJ/UemjPQ2qUsc8d8FNqCZqH5mZxUzRNrH
k3MtZHIPKYlKx2wO6WtK+8L353/RuNMkXDnKwq+fXv7Hxm/7loUrNnmam1THLvbJ
JcYZjCvP3sdtaxfjSYtm6nkwPDl8X/JHabIciYTGHL9y5fT5KZ3LmLrRv0vwLNYB
aKd22W3QkBGZI68Ovu8tS881ACukwloEz93FxqaIYPPWM/oGFJ4Ugd5EJSrW95Ho
zPKR9mbvWKmW5IZcykbjd+hXxeSQ6kDPfrVwI2SxvoAnECwtGLtntIsIK9DubUW6
GTHeENW7lQroETZfpcW0r/5SDsDwRxa2wcpOHR4pG0eslTrlPV1aTG65JT5jHxl8
YiyFCtODPUDH6a+iyEddWw7+cm+xTV+zRSzJJJJOWXjIXKHPKS68jac+SwGY0q8p
s7B64pkNlrKNicGjp0CqOz7vv/Oy63Sa5r1/V/DcyMOMeTy//4rV7fdjNE166u8m
5jb97myq3OxGv2/hcanBENoSnWymzE3Arh6KINq31pBwLZaZ0Bv8nZFQy4EdlhO9
0GGaS7+1ZE+IgDBFlfOJNbyxGGeg9pO1EwpYsBbi0WkJLrV6ib6J4JOGu73FhoBA
0fmFIt3+kJXfEkINGHAjG7KMKWk1I/ymedFLdsNIkj4bGPT2nVv5EIFQ5FGifbvn
4PR/ZvMqxls0QZr4rTQ3wTZO1Cj7tVlsSpodvQzA/vKG+gBolhg2DUUq8dHhHS4J
+AxncKzzoUCUUtql4hK+wMDw2i/PXkUExtvCtCU7kOw9R4Zn1OY61MALgRLTSET1
0bnEx5NEn1l6HtWVLgr47UFLRAzsvFlViPYi0IrEOoOPs3MPcr4WPaLYGdIet1Ke
SJ5IORDcP1K9QQREfxmf5SVDOUBt17oISeGlSvWM5oenDtykA4RFNBUjJkQEmbYr
E8Qe4JM62xQ5N4K1Gi0wSuTZy21ztnCzm1ntBQ5bMWWvaQ1rmceYQXsNiTsCQumz
z5Ucv99uOdmq3F3ccMvviuDgSTQFEPnV8wZcioA/XKPaEiqqcyN08Us5lFHmtEfN
d0b5yZlkMyD2KIxPNMmJDluibWLB85P7/wi2bdUh3ruqvQhH5GC/2G3p6BCxsVeA
0Bi1VN2mqEUqBVofWVqfp7ngjVxMlsU6dTUeINuOXu7dRS4kEwppyrxwpZR3dCoy
1MM9PkCo+QQq/naZATZW3al7St1osnyffha1k3uBH5OyOCJHeXoY5oScKt1xZnv4
kVlMb6qjZfIpgrgvUdM/pi9mzaQww+7QivFX1J3Ziby5IP/8pGZD3kUQeyn2Kg9B
kgjeT4R3W5bUkXYNaarUI1OUBClcBS+rw1ipF3i+hFIX27MJF/jg+CEBR3Iz3rfR
ktTdUv381RmYLFojwcZhKpKwIq03iMsnw8a3Uh+XynTS19ckjrfmjfNBiTUEwgPV
DZkV6E62MBCtd5owgZxhBlGFkcMNGc9M8kiWQ6St4XVP4xU6YNEnMof50/jkdHW6
4/ZpZ8QvzMY3l/QDkMltRfwFTiVmnm2ENfRAtFBp7KeNfe4foqOBPt86jdVR3VrT
b35O7VdNFMBTgO5aoJcYemIVuVTPhwCkYT+zttAUp/sfniHj8prXhlG0XBlGe5li
NLlpXKytsU/XCCcPplAbaXpZIVwJVDmKAv+YhM7mqhQ2BdMC4pXeYtj/F2up1Q5I
vF33YqAjMvzZecCUoxVe14SU/caNmrqmWehVtKDwUoqA/lZqDF/0V875XSmUEp9B
mzajHa3tJ0+UYznwufnL2f3CpcnN7waykos+VWB/l7icAwtHY3Zppbm1foOWbzSk
viLzz+wDwkxLJMVax6vo0kLcVaQyTKeeUmDwcbxrGEiyg8OKL9vGSqBvg6lR/dsu
sFY8vbVsaXle5eYxbofe1Ebzk/pPLzzxfYTMxCJ2Qkt0pshCwGAXeC1lFMNbBeTj
AMZ7OEcLUZZFnsXuVS4Ctg0kOg5lVGtm/njO2tVL7R7dORmY93lm0QhTZt7I/RbF
sG0b7lBmdLVFqkAXPORa42vVRZ+qV+8+UGuUWQAdSMSL/kRIOMt6EcMyzTio5yKB
EpKXEXV6gDTODsxRvLEEkCMfxbBBvPrnnP5B1Vopi353Mud8q4xjNcT43Wndbfri
yaWb3hl03MFv+Awl4Q1f/snDJD2DU4c0A+tcptzqT1I4iCi5T6cJeaRlP9hJR4CE
J3St50amVetqj2qml7v1NB99G3fzY7o7rZL1y7t4Vylpt2cVNwdv0YodmbqIEw23
mGhrpj0NtamiU4XBZv3Bi2/SCf2Gn6JBaLEg6HISPQBs3aVHF4HV4x383dXHjidW
Z/1L51JSKS5CTDig6vpRK5sdY5DdnfsBdcz/Ed1kj+WhysA8IB+v5CepCHtPig2J
pC4KPOIRLTb6OK1mF0K6/OhhE6No2ViNk7hShw9UyiLB14dumuPklas7j/F4mxgH
oTK5quErQHa/KaNLwT3Yb9xYI/bJcymCPCBxuNVXenyQKC6sQSZKZjK0vjPApBTR
fwGqi1fjVmx6vZYBw6xZMH8DDtQAY90FkAgFK+7gfmdi7fVxqVZpseyInLxMQB0A
R8tcqYSx+KpTOnuJScrcc0EAE3eewA9pCNtNCfLdP9eJRg0JcbdIH/ccmOV1/RSq
lZcEJklR0JMFwXX29i/qNLzIJUiUCcJX/rPkKA5d8jCcI58YX1q56Q3QJk4RCTS+
kN87lYDEMx1hCi6z05J3gTHMV+v7v8HeJijB6UdxTrX5WhaVei7rIttWUIAWgdqj
SePY0DYS/5tBPZz+pDfAN1wLZgxbrCYerZJwettQP0DnbonbhTO34kDoNyqMugzl
ncLFiv4YPkb76mKUYSOPCj7IiTkmM0PJTP57uTKkFHMmMj7gtTrctXiE6Ds1wMeo
U8Cse3SSk6JizwrPS1KISflmoaFS5J7g4g3sZusMiFe9zvAK1Rm17PlcCyO8ATp/
N83hoFryQ3E1Kv1NFFQkEXWrJVq9GLVO6Zgj7pzntUNQ1Pe3AswFdPRFBFI7qF7c
HszROxNLN3O4eIfOu+fLRiz3qwfg6O1iH+Rl5MGzJeBii84oos6RtaH4ClwBgGfb
bSV/je88tNTtBYOYYyXMB6modmj3nj+8ve7gpQCaOwODgkND9FDGcu8ZYrv0k073
gcOM0/UKkGYBW11GTSOpCb9uq+xoZpOLQvX1pHMi7/FnXTGQ5Paic/sPdWY7eQhL
jcVLd/W/XKC9MJmNRoO1Rc3dNu6k6Ia8NU6XnYSBgrOR6NEYsqpXOMKLkMmQQmDi
rLFH0ZYAFDhu75Iw+vMoLCxIeuvFUPojntAo4ijblkA3ZtMefCycdpybjhAF7ZAZ
6LkQCnD/vxXYggAlWXPTt6Q/VmF/QDq4ce8djURN1yKbsA/LyGeuQCTUB5UymfDE
TVNFYBXRIKIMZKFk2goq9kgosg2FcJ7c4Sj6BL21SQZH7b0IpNEafjEaJbISkRzq
A1Zzrrop2Hmq7XvAFYYlTWMVH/NRXsqy5QkvhoV7Fq3h8FEdRcnrqENDJUMi88qD
m5NrWhPrHCax8T582WdjTvXMSFBYnV3UjaLOEC5+ihu7bVrfGDdSrtUKErvOapss
YnLN43x36mEAnMx6MQMiJ83NgLJiQN1OFQAiWrkerFOrDuFsVQ26FQ6gtxGP/G6R
fadR7Rt7oyNL9fmRExUMlbZnxNXPAv7xlAwq0hUjSJu3LYFlcrEYYmEO2oCVJrZR
m+INk6wHgjEBrqfYk9AzXb5hiwSCHw7/TgHV/vqkZp87jIkSaSQSj0qvBl/Xbrf+
u3lBdoHE6/vXE1TdUfmgmSuyaZBTCgXXxXhIe0AyOCiGiMr23X7f7I6lrvPsn5LS
UqcHyBPt8CRkmdDn2TEfheCTsdMIQIjnEEt0n17m8HS2Y2nK3/YV9MiDmBAKH/c9
mMgBcpFZKeMHUxUjHP1O/exWAihM1Bdw1r6AMgGQglubQPHp1gxwzCz+mVaExIDA
hx0rQe7DJQxC1oMUNclaNZqvxS2kxAoEJ8xMQEJ4gP6F5BtHIXiIIDI3sIG2HF4G
mc3TK4S4f9+lHOYaXihmK4wrADOnY9FHEFG6il8IWiuJtoPXUuGNF0G93IGiVBBR
j4mqYk39/AZ9r5+YUkDx4eLpQvkwxS+MJT0HyHcrruqkHxuMZaydzXXpr5HKf7MR
NHB1mo0KdFy577zDib7ityxXCZssN77cdDtjgwik/jIG5Bd3URB8BmjipTYv9n3F
vd+h8kKfr53SLKc/T2e/57OigE5szPzoHV3P9jgAnpgIOgCECF71QOQFZn2Kl2Va
Mtdn/RPDye4EclTMTXmRKVaaAO+P124qo7q/roAH8D8ytYEPJL2UP5k9og09YmKE
YBrei0QBPCU/0thqqjZjntPZ1dt+z6buT7O53tvWcIap8uLOP6Nx6RlOv//XZSPU
wtghC3wlgWkCJAExTPvgCGQQXc+ii/NPJeWxh9aO7Wp6TRcaasFVFU7cFdHxPWwc
RZC21fDom1pOs7fglFyB6p0C8Hhj2behVimCjb9BgssJh8V/jOfXDIdQ5HwxxWuC
XMyTc2ZXKOat2BypGsHyTIta6WbTfrojD8vhyu0LgOko9/PRm95ItRRbOPJboSJI
uophZO99sp9T5Qk1vY366dfXuJHNG17v3cSoylG8NoDAYL4t9Vq5SjCkcVSI9j+t
5p37/er4qL059Z5wL4/uQL89H70zRlE/Xz0d/MiKDcWO+lD06OCgxoUD5ippRbnu
+GpxwC79cRO9vUMLkNXrldpmFqUMNi91OBbXUqhYPQr3nSSajlLcodFdNDKi3Wna
SFj57UL/9KlZ6GQomR/1Qx7qD2eCN1rmDkP47MfPwx7lRDg/+i/1Gifp+r2mL3pd
RDZDGu7pCaYrhO8s+lGG85grGW/r5wkoltc7gV1hOPJC/GDwCVKS7W+1N+TSneiZ
41mWjl4l5887G7vQ+d/faNl1vHs87MTxnK12HiCe3ePc9lHb9d5eedU9WAs5Z9RU
BDtYD62Sks+pROhsvdHMkTJgRDrZ86+Xl7Khk1qVaxqHTj3cTB8YEWcqP4+RbXHz
u08Z8wgEbc544XZyfLd91fDm96JRLNHD6MJB5RDrYHvTjqKNUSTJ0sCFbk0Mogk1
wxy/04LD0xZVYfBrfXKtLn5SJPlmjOrx/iCINmNDSbawYcx+Jci47gJ1ZQGAR1+5
ppRH1EooIvjdhfWtP0D0QNosAqegjpR/4Wsjy/WFIjSSsMXgCa0zRxjm142S1613
RBVEAxRA9QL2IaMykUd6t7ebnlGvu+7CrGAIykGygYL3HkJSScRTzJglK13Rj6im
erbv8JIc6eFUxYse6+hfHz6U/MdAuBe6riPulZJyoQYxJLG5kaTpb9BoVJAt64ln
UN64VJSm+MTun67C32kh8cMyDchxfb29890HPHHi3zUDt8/EXHnkd9Dgiz1rTlB2
WrF+QsKJHQn0iwunDndGtxpNQSA+fQnIhX8rkzR3SL8ih6CodbzGaItuS5J2gxZi
zi8B04W1YVZqHCkJKzanNYAxPkdjtLe17K+Sm8ODtWG0RZ+XbUkF4BWdtJ8JP0zs
Tun86HVh5MNtpFfcnTiAd6JS9IXMgcs5IXTKt9V1XR/NzhEf1czJfoy0saxkztYw
2qqaTqlN/7zxjicCQJfnJTGNiHFIoRyItA1Nn6uZxg8nkp7+StyUGvMyVF7pEVVZ
wsqi3j5nT83vK4HQnFzEbL7ll0n25yfplWlG3cYGE3qkCmboWVrcLaSU3vheUzQa
d9JcyeqoH/oNe4h6JAAryR4yo0SE4rjdPHYwqf5djCyLHoR+g1OJ4/Yylw1Ti0nJ
Cwn3ko9WJUcriQ8obKC+PF+CcF5m6DsjvXNI224Ukv1QuWbT/faofIokYtF9n1QB
qDxVXMFPR+i8JvrH2oOAjXfTf1EM0wgdQP4eWDyhWi/pvplQBb+yyOGVCcN2ECJm
icK4LBLZNnnKwm2TzoOM2hBIFplyWPuU6J9xb2ma4TMhWx/+mIphcAoaBWGXwKve
37FU9gHvPD+KT8v9PeUVxf2kp6BEj6SIMkZBacr/vXEhZWkC2k3lYd84sHCIG7ze
Skny0G+kc9uFiZsPPMYv1ETdc2d/KtxD+OJlUNn5kPO8d5MSk/gEGQT/+xRjxZuH
/rHR5nf9gbDxPQ3VbFwRXpaqF/OManp/OVXGbrXZqEdyca1k/W80HnDZ1Tsxn8c9
eSvAek+VA902e5d/SKBJwHOAKqtj4O7VZy/XeCeK5T4xHSaML4rOcdMoAA7iAkS3
W6kFT+iFz6N5w2Fv7wB6g5VhUzl9k4rKxAEm9odq4huuIkKFdR/Ea2cLldcY2lKF
mtbaFeeKtlEgJYJN8Mwz/QI/Kn1b28iJkW6Rh9QcIvycnU/N0juW0dDEntjiiTss
3oJnGEcbytH3OGAp4dFTRTMJHgy1cdNROIDf7UxcAr341F+aW07nyFOtKSQnGAuP
mdtBzcHgr4NSYZ6w0yZL0OhOu0d57lm5ThyFvwfscoBI6689ExS11gw/RNCyr/bP
y76xA/+FfyyDPZnQGDSdb4w9+o72ANfvKAdsRiWEkEZ3m26pHmSqs8rRXCV4irBu
CmNE7iNIZA/B1s9bc+j9+FsAeR2XMxsr8o7lO7OfauBX91/uiV2xkTrbRMC5H/MD
FI7qBke564nzwWQuwG/cYd5A+UumqN+01Qgf2AtrsF6Ku+3OIgnuL1Z8bpbhaID4
QRW/Q1m0LukUCawqXellOCTRXDHLIG7c8ZMPpY618QRHGuZ89SDnr/TA/PvKx9xm
loWNfKAQONVmXPoCizdmd1YM6L9SPJiUoCMo6hH+r4WEXGbfQVYFUYA7YFxOL+Ti
I3zP/GvyYhJKlOmguPSK5QEhoj11rrPFpnezIBDlXDKJpG8ceoFXkOsxi7yyB0AU
V6LjTYMTElsRhwT3co3NZPbsq/6dZM5f6XTqUalt9X+OOJCtVTcB2V/cc0ZWogGN
jKuF4EU8Jmr8gIYnUvuKaNjykX5G51R7BxSfGHMOCW5BcvclaK+vP3MEoUntJxz8
/ppiX3S6OnaD0xyk8HnJAuyje00MWI72l35dDdCIteqbl2+rY6U7d+A6nGt6CYMX
MwSfGY5TR2KggX2xrnGWhwlAXX0mRwHLXZgI2mH6dbiss3zYP9SYsmZzWS9j25S7
uSZcluktsEjI+SBCC5314Ri9podBm+ov9/46ph2SUsNm3gO5jzdcEyBl1AtfO5XD
lWLrr6WuOdSGxptnRX0XzkN3m22nkxIsa2Ugkh++6TKMUysYX3mfuYoiEWVOtVgp
AJ6a7kosM4xtYfOLaeAwbDeqRB3VzFT2P7okEBFFMbgB7jVmXMoFo0AswtiwT3sK
M8jdZtvGhbIq5v6SpLAuKHRqE2rGdRyIkw58oVrERsAnG0xiGQpIaZ8tZrA7dEGu
7i8tdQVrNrjPaQ0Wylb9e5VuYn+CJgTRs3vmolWxnuw3/w4dy4bdh9OlzOldq0hL
ILyKczcDoqDNFGV2d+USZRmh/cpBkslL9N6bWKA8ulm/bnNXMJRE2W7eeMW5Y123
Wi9+5tI8dl1Ro3/O6Izb++BbBf9oipk3xPtyG4oGoHedsfLsUwumT9VpsvxrHcNv
BBbtXq+9V0cqsHkQpqDTrayFXeBekErAc92mUFfrQ7Uoyrp3UQtywGqeUyFV1sa7
OokIWIRs75bTHT3+G+eQYFoWMYxTRTiA0rbaMgR/zOW/RqPaPp03Zrag0DAinSji
HATU54/snD2r//UqlfplASs/KH+K87OjzjINdmrcSCOeVgr1y/S+hmDMeBJez6lf
4jDn/Jxe+wdH27XgLCg7qWpDcUmuyynRzNjsAfqfpSUOt56dKedXPmehWgzCjk+9
/gyuMd2GxW9H9jyPda85mG67/mSsHvlirYVcj0Pv6LYoJ+5ZNeEi+q8bJQ8EO6Ux
sTb9w0LayFOl1KO7S7v7m5lZ8GXK+LPLc0YNDasCMdgRPjhF8KUNSsZzQDe1Pkbs
77C27yHyIPl7gbnerU7QiITiIR2f4p557eCgJfGIqo8Wmv9IZBcieaXSiLizve+a
YKDaTkVEjtduw/DiMZqCBlN1eHZJZuDQMdln2Eumdk0Fz0oQmqvGC2vj7G+U752a
vrHOxgM+ZL5aY0OAVB1v38M8vzQuSxr5LhKmsARWrkpdS4dK+cyi2cxNDd3t7lwi
9744pdcejbennGIEPE+zs7v3KXy/E9+5zkh5ExVSQhrLPA87ZVxycj6uvkXv2M4P
L5dmxTyDywSqRsCpfr0nm4ECMa8VDeBeuRYCV4OjxebCq8JT+T5nffvBQl4mkq5M
VpK/ubly2bjCREJAr5wXYiHgvs5eIV3wUgc0hYD92U5LVknV1zUkrTrVIziNe6+h
IGRsHPCSgX/PGzQHViAG1+c9NLeQq/6ZvZm+KRjGssvBlpJV5GteG/98rTozlv/p
6n4NjEoIo1borYlr54T1AzAbDXfNCoF83CpbflWFxT9Tsj3uZUruhoOK+jJYllBD
8n81NQE5pibc/3LYa1yY/aIAkA1CKhanNwfvL2o4LOVwN75kmUdJMgmpxokDwjtp
lb6ap4Iwj3fVZFTqf5GK83//hDSSz1nYK745kihQ1ayYa13RUjgy65R3QJEAbKU8
bplYeR0I0q0P5hcuSS7S67DO4xWsM1Ta6hx7jXY37JahBOGyNQp74xrbk8yNDWci
Gn/W0XMnBnZqePpizZ5zEr1LHke1HS/ePaM3HIzQf8ViyjFs1F6CUIKsU15VZOFu
KYMoDJWDyqGwXmwVuX9F+//dhEb4byZuWnzSWfveB8UG58fywa+MGXZRo+uiQwpA
mSOfqce8NVjc7fmE6x3cFvAC5gQFeSjt1z93qE90EWnHGLkIeFIPc/CCcgrQ8Vam
LAlv3QmOpCf0dHEX6rolOgVGvEZXQJcwSR4+SML1KyP/ZP1+9Tyde9N/Kvr7rBLK
Q7CqUGAKsUJMimy1sjFeDdsiCIStB7ghvhXvd7oX02b7AJQ2sEkkWzKAlrypZkhb
SKtzia4zU5bLRhUGasa6JjGeaKdvOnlA8EAgBmu3+Z64O0kwRnqsdI7dxW99rFsm
9oS1xBN8Zlhk7vJqrKG2Xey1va6uoye8iqcHmlZqmV1e8rUBcfz7gzIXx2PDx8KM
Oiug4u+0iOBfg38PVSx/CN6aK/AK02V3TNBUyVFmKSROo9ENOLEKKCmP7Z5kaaRr
olNzD2LiQUKD6bBDdvgG5yrPtQzVhVQfGzd7H+rGAZ2VM4GuPN6kMmVpbwS9usZO
ZuWhsRgKE7Sx8j0fOFnIbYy/mSt7/We6I1JzSEoTaAuL/5SwfzO8mFoRA25iAywY
gfr0wMuqDCBwvwuNp7OblJm6/xZdDQ8FgtExa8es3QwD+3gIA3GKVn6ZfYYsEkFh
kVmvLBLsmhLdCUZeKkWvxO8BvLVF3PJ8eNqdil++pHJeuEiof7xd4RiZCXrAjW6t
lR0DzV0PkvoVPNZ2OUnbSvT+xZ5eCMao2c7TcMiJ3cLpZIMRUqIjH4vuEN3/wIY3
49TSD1n+RjAkXJIJGcwvNpWPUoeRalGTCQVDK4H1V0IasgVN/SHI0jjns11brBG3
drPhdkKKiJ/oIUfcU6ERYppQxM6VbLnZHy/YL5DtMPqCHeHEKp1zfjy1lK7wQQhZ
BDKwVMiWfcm3pfa/eHiAzp32EoZKQAxQlof0n4MmsUcAtyM76u+B/RCQYloH/Ppr
YEh3FwbMcNN4VbAGgEA+I/SHU0o9Ya0njQXoA34AoY/0SpEteEBkLtqUiK4cJF6R
wDLSDlIpFE7NJ4yc4bfMfmsH3WMGEgmYmB/LWk8WPpWMo1bnkx2Bk1v0b5LiFTRX
DzLHQ1JBV7uHA+JcJAF7Ctgky9iQlfpRbsS2h8jbDTRHqVQ+17aHOx08h6gnPSCp
L5fVotA44vgGMPtBYoPCiwLHCHljBSN6DtWvCf7eQzo/VE5EfVMgzesowXGG6qXj
tvJ3ruho2dasDJLSV6GObptbbAuuEsjUOMdNeSvKiUWwEEyOc8Jh/PoR9nn8D/nY
RelL2A6XIYM9tneoHBm1SCJIdRiXtJPSBbSyoOo9CIfGuS++GmKmaV8EmHLg0AyL
rv1hIYwv+dkJ3RXVMya9PUwOOpYxmp21gD2YF2LsnhkpnWhCOgq4uGgBo4M7+0CK
wOqG9h1ynMnoDCT+allfvlZ2kCHXup+IU9xqaZWJYx2kWWC70pPZcqc+CbpmUAC3
YoUjmndnO7d/YR+93hQh4iELlWEKWPKqBCJ0e+rlApb7MTS0k25r15NW4bU8CnSg
JcfcG/VaXC4ySXk6HQd3M4kbXNaXTDJRyq7d1yxPgk4nEe0Z8UTBDAGZBLmfAE22
y9c3MAZYkql9F0HmtUgkmKXCJ8Uh1wwCBDFxJl0PLPxJhIHNkkr+hfqRLhtGj7DF
BiiGnfxQqhpW9kDNH9FAHNJtrTVwOt5oCNFgHq4PYZ2FVjEST5Go+pM1YbLmv7UX
T2ZtBaAac033yFb9e7Z5hJMdAJFzzOzSoqf7FMedT2kz9I9q8DufnED1Ua4C5EBQ
ljy4kLFR0bTZwOlHGFpLfCEYW0iHhQdaDoijGVrQb4GdIxW+CracHggtC47kcnxl
8FQWq9f+m+tb+49K4TomEs4qFnIoMC8Lf4yS16jCi8gWzyh6V7DwD+uVWusgiof4
pvTfqqlVZmGkHYJkqEEk83mY+WFcIsBqFgljaNXC7t8hUoggQ3nEEiFj3tNdfZ5e
eL5qenW6RYedMfXMHmsBLJTqAWV9WMbiKk/tf24bFSav8EHq++U+ebRIDw533xaz
h6s8/ST/I7dJqPvQK/J6x88Ut5187gLquettXM9CZGpVHmoxuxK9bvLqHLLkbu5g
bv1fkDCFapkbd8Za4PD+Px2kPh8aFzEgCnXcXde3ktsOQukwyMWdTy3MB0hSmsYQ
mmLFzzztWFnqRYZnS0SBaLUI5Ao22s4rO+5YZTm/fGmf5kTE7aKhzs6csBtiHOfU
RHxcZlEIUYnEebVmAAXg13+sL5gx4r6WUo38m+bLUL6A/gua7/ImeuweZ15qbEyX
WVbJ/aR7mR9rX3db8kBFP9bOePoGyQQdGgYYjqH+8+ov1tZn7ljniwqXWzxVM2+C
05gyJNqTfT/rZf8sbImN0WZ96KQhs/ohbjEV0EgFOmeoHkmP9tYOrlvHkhp+IOJO
4/tLgZDOLumSL5tc/5BdMiZjbqfIiYkCo0lD2RodSdTQWCp95+2A6asvWQVAfMaK
tqAdXrp9ojCTMHydJTOPrCA+CR/aXkamY+oz+sSZXj+j3ru0zmZTgExignFP3bum
i3JBfgjEilq+merQswdVDsQ8mmTMytj9T1PzhhscxpuVV5SiyTT7vnAmWjzGItTD
1c7BwHmrKfCTiSmTkMUdew2aclMTZ/Rqr7hlTQ6bZf3M79sEgzfFr9NQ5YO0g0We
oOK6Oh3Mw/MkPZq0EMCGICdHAHmD2Rpg+TIuEhzT2xpgjM3uGy9+nvtT+DQrQdKU
SxQudHaUpFh+IZGwj1TC4Oo/Be/hcVQIi7PzpHhZ7suFDgjPzer2qSeNlawmxMqB
ISpwi5F9QcW3KDTbJDCvgLokCSQzGOxUJGo95MvcBn5SVS0sABj8fV82IwKHoRjY
ZveYMNe+jVIE/BB7Ig9kP+BfuLL6t7pSCDLOAXu7DkEPD4OBXlL9CKzp677XQS5D
oZUc+JSpWJhzEN7j7WFaj3C79VfIHORCW0RpGh02L0NFc7+Is8pyoV04kOIlqQJn
e8+DRhxiKq16wlvN7bHWu1U6BFE7wj10M8+HedgO/++nqAb+sL4qYwVS4gr8ImTW
wdhns9tNM0h+T045x0JWOMPoCtWDbo7DTTtnOHgzZZsv8RXOJ50Aie2gtOy0LcXN
rPWnXdztB6gMVEUP8nht51mk3VMrMOOg5U2MvMnCjVpMtWOGuhHslhdcE30aPUL0
LhMtH3v/h6F1ZTvGRrflpobHGIAZBTWBfnlIB8WiKszCEMf6vzlbLbdEkpzxq/3K
CPzMm8teQrZlGB5ClRPRKA6LBNzIJ6kNW3Ozw8TuEhNLNm3zINom2liL5r3+tLaU
f272GiKMzrHp667OvkEkM3SNfDNYdHyXPsb9UoMJo0C/4DAmpxU/Aoyim2COOHOv
AmD9ReMj0T1lWfNwzKOKPgoEEuf0sTYbhxnR2LH8n9DCfmqIbpv2j/7twNy61/4t
uCH0H9d892yz4tmfbiahrIIPMvSFMqjgIlotUWOA26lX9b45ygpd/w7dVvQ/rOv9
j1wLQhFxYHxcMzeY3GEcHx2GTfC/ypxtnbG4DcC3+bY4yNmF6etbumvTOgLGoWBi
0SCX6X9Anm+qbNucQmXBbPHnMTyGCykWRgl+bZlD+NaoSvx8oc58bTRXxWyzI/0x
znkh7vHAsfvMOu+QUVZOHx8atF0B53lpnjV37l42ldx1mhu7r8r+6Jz44CTsGNmq
AGrmStdTYmoUEHF1QCKzOxtW0gqlY7jrUBBL88wLz3BL2PVwRgNo2Twlx4HASqEj
VwfIONEpE8wGKju9+/277wrzSoxxKHuIHbVlQyVDyeb7yn8JK+iki3FZ62Dv6kzc
irFJgKmUu4ywGZ6mN3ee7YmtDEWuOIzcbx6k/H3NLWNE32TRFD4qa7H8I8ElvYcm
9foC6R9NBYTHmARXwHliW063r7CMweFaHBjixMTpf9G44Mn0lHLdE7Xrfh0AfJhJ
RFLe6BeXgJuT/K5K4Br+JXq1/LK71AC6lw8l2bbeXhaquh0FtYP04ZMBQoGRFU0Y
TyvgkBK/pLUNGkemdOOXFWoq4Spbs3lkqdYVWsp7N+tVrYN41nbuHHoX9SYSchHD
X8aZQQkfjBd0C/eccS1FkKJYSQmP/vRxvnOB5KJqZoj4qClg4HRNGXrkY2+297Z1
YCINDpIHv/LT4z5o7KlBvEedvvrxeZDFdsW/8znaYgtHaR2zAEEEUM382wBjWjIZ
g14D/H5ij0kGY6gd6sNFhjVGe82z0/L31Y3Vn5j7IUPwjYcPEVfnyP9cwddMZHts
8vZ9o2hgxctGL+7cUD6BxHfs3kVGXZlWUxDfU/3vtMvujAx61pMsM/VnK4dfMV3+
J7JvDpMV6S4mHj1+QIrddHEdpGfbGQg0xEK4kjnEZ752+P75TvH/fJA2QMWFBCfr
PYkv4XzAdyBo7vAcmClNDTh0xM1fnPY/CNfVmRnjKNJ9qP6pZjyXpLBq9jsXsViU
u1d12UXjPpeDqpnjGxs/p7wN68BDipyrdNVMAFbAMP/lBToktWJgkbAoRLVwrKsm
0gHDcM9wUXBYj3GOez7y7ffQbRG64Go9AApk8uVRauosz0itK46255X2avser6Hn
B5RGRysDMvcqS1ROLlaC4fzRvmnry+QJOryoeuD1+aTF1asdbI7EuASIk4vsH2zJ
eV77aXVZBSbxLGYSqRPkQcn7g/tMReADNcQtDtUtIo9CynzVNtWE20rfMYu6eyZF
hYWnlaN6yNnIxW/P6MyOFVk73wYVXeGdocpApYfXMkoUu31ea1oiPh3THpZ/Sebh
/U0bTavcQnuSi0UKjhnvscHxD/46w++K5SiQJdEy9bWbJeQXBCuV5RVCTIi8jDF5
29vYlbGoekBLocyhcuak9nCsSMT5lAxZw9Jkmm7r1N/jW/2EvAlVmIViNqIFtmcE
nxHhDoKSoLwtQ0l58y6lO6NrKbn/17eAip2vzWBNYKFUqPbJNztHjF83gKNTyMZJ
8BS5dsNME4R+3j7x3tz46b/OIbXvEyDvb/TwM6/5FDNU/zyHs2+4iVzhk3Hua7+b
6VtjJFEXcP+IafD0cd2qWHgBD6LlqzihW13KGdYF90zTgZDjRhI6+E1KF7zPIOwJ
34qpLQw9SkQMVegPNwE9IlDm2SDsj7XkyPIab8GqaL/iWApZ1Z/cjFBP3trc556m
i0wwWdOQaQrJJPXA3zBvNMdZxGcegmTdSa4k/w8ya95Enez/ZY1RynxrybBWS8iM
e3GVQibrD7s6xDvd4JjYkNs4upi1nIO1oGkIAVBv71GTX2DebKSOMympG/B62/UJ
QRaoI+s22SyR2L/YlRBS3HX/5bRCIYzuPTy+X0O+tciR9Z6741CV5IcdnQPhPKDO
EKFsbQKI+5UxHmnK1W4cHPUdiir+IoCnAry1UJn0X6GNMmrzV0uPnzX+00i674++
MGyD9yZlcoyBAVTD/YbRBDnkSgZVeF2kvZ1qr743fcCLTP9kzyg9jThP0B4YwcVF
7ypqupkeYuOJw73tpzugl1Ld825bYABVOCMHh0GJdilDi4vi3nhvnp7UlcpDsDQ3
tESLsMufuLcYKAcWKHHiuMWJKo2kSsnFnFJyo8GvD8r1CsW4sJ972DDRZ3W0k3tS
PEdgqi1qnhuToOu/yg1ud8M4fBXFA82E9oPggIjMNECd9XGo3/c85v9Y+tbkn0T8
Lq+fnP40oVCPooiRZHjvArbHNEu/yznf1bnHpww03DqHU0XvUDR443DsmMZV+fFI
XC0e/GoUHZ+OMDuX6DR8fblhKw9zizJoM3wvIMSIy02XqgYIR/abZSzoqbPlfm5D
/WzKtJaZJ3gstzvJFEq78l4rAHrSoUwcc/3Af81DQY4QR3AJmRE0/j4S364oRFu0
KQVYU7pzW0hi+N/zwU1iKkj4NAbBPCHVrjbhof5XPLArLcOMsR1G4NTuUWuLQol3
13uRn+JXLda3OGzm+atFOv1ZIT3m2CcWZSOwoUbzIzLWTtr/R3XHVflqhjNmhpB+
nahl6ULtOEs7Dtt7MJlBsc1mbxoIgXxCJ0Z04yH8f+kDQ5dB7PXOfzFpbrdNDsj5
qk9TFs9O8pQnQ7E0m6kbfqvQwgmKE2klLnhaPhqovRvXACu0tTnR84rbX9XMhlN2
Pl0awO9iR6Tqarwnyche1X+Fz7bS5QEiRaPZiZ931KAbxtepW20C3tVRN9Bs5OOV
OelOf4nlwGlOorLot8YRx1dnDJ9P+oFcxNUsG8c4G6KeB0qF8tKrWCYSmaOSENiw
5Nngxj2oKig3WkaFHMrbSBh7OBNzar1yhgrSvTDbXL77tPgjYN/BGRdT3jPDR5Oy
Aflxq6EQXdZSt5w3YBaZ5cqmkLxj/B0D7FlPQYSlbPOj+7GdyKG67hGbRjGqL0PO
ZVEjRsz+X+BEit9RLSHEOPxZDOyNqARhMMzv07umNky9S2h6aaQcMLTHj6Z920km
fk5re7IO5SYyqQyeHEIlGQWWo5eR+9FfWBsC4DvcbSCulIQH+n9kRU/FY/ZnYZa+
p1U8QQ1Gevy2YLlLkxeHwiKLQheEfRWCFUG6BjA77AQElyQb0jcYuACGc0sP+YYl
a49MH/npjiTFfelml+SqaMZ5BavF15mkdwjBcuDvIdsg+lxwvNarr6HahMxMoBDo
ITkiaVfIr+lnhJJujQqr1omQxSHzx3SlHE1NDsMNWgcnVmNCopY8VQ/eKMnRWTF/
PqjdEbd9gsuy3MI4fwXSDfXmhFgbEbZ1hcitoPaKbXFAw4rB/L1/VYWrQX89S1kX
bIrEsHwuuaos7VJQh9f99WFpDXQHscjalSsFKvWpY+a02bKrc5AuvkKefjbUdxE0
6Yum13oX3xb7yeEi5f75D4b2ZycZzuoWxZkzutnhNnDPIN9O3MF+J9e97mrT6myL
9fPy48k04GwPbqbPS17aAZ77wxl4NqD3JPVxgUoqb5Ack72zHNfylYPaEdSlsMbL
fQyhswjjKTNKGml7gykby2fcdzl16UYYVcqsxkO97bKLFpAHatdNtRlg76N2P5oN
Uz4GVhH9yU4s6CqHM+JaI0RirUZHuRswfcvS4NfkvrWkfM1rQEvh7Smh53gBTutx
NPCPnJz6vw2442iTAfRuZvtnKemmqHtpwDAUD4WdmYA/govkRPjHuIt6ZNWMZUJp
LiNEBS6zPR2zclpNGkePFIAG79+Hei9Q88R8Wxu6WMsWBA+ovdAJWPVjJb6SHNhS
n+GBNRxLkDxt6Ydl4RwGIOWZvm1lJhY6vBuxtVi4YMhRTBOb6awObFv7Pmh+EBSY
1dx0+W35ao/dziqnMVxDGFTAdX72fdDUsRosd/kl6hn55GvqCTX3bhjWZFiPuPWC
p6LhOZL5s8oUKfWi3MYiWL5cl5aukQmm5GTiMJqN2i2sfPOT+v1NfMIIB8L29uIc
FKziWWHKHUYDkpYFU8Lg34i2JCXVzXapZ84/696pnjh4nKf9paaV30NmQEwTOrhd
uND8CWulnYUgWrde2uhqSaJ6BBbNqKQmJ5OVMuEhslmcUCc2bgppRkiqHwPK5mQy
e5KjyXGRIuZc1DTrVJZ2rNesGL3GodGrHTd8w6Yy6+khypJtkldsSIdHf9WR2H/G
wcvuVT1iqiONGtU+kZsFuCMY/TVPah7iX11eBqVSJl5iVdy5/G7JyKBytpMO+LbQ
5SUkIrRGXpKHADN8WwD6uPbjHcvHc3AEhOHpA4B5c81eoJRyjdkJ7SNmcQF1TMlu
9QGZPEumFv+RrneRAl6ECbWJTMsVJzbp6NQ4SpnDAjC3D+5J4efbBl85JQmZ9Jo8
NHTa63/JqODTrQ3cI60NSaH59iRjg4Rj/Lh3lmk/NKvbjH6Bhfky0pQ66jbzLvA6
LXpRmMi060hVUEGk8gjDGolOxkVUXS334t1ZuGZBn1JoBKDb1JM6fStKxMSAtx6h
y7pDW+DU+F1+kybVbprgZpc3yTCBrbSZobeMB3GkvgsqDzDlYgISI5xZcSGCDhc1
rHCW4ovcEPOSHNpUytWTq6ahpYOto2BXWPe0uw3RTow55b1fOytA0GZot0hKvEe4
tsd/26y/a74SgCzcsDarK35Km7cnI8Xr3Q6jkeyU3V2CSrJRHerv5vOfHOr6quXx
CxIXscma5eq1VTRxGc+zTDwUtOvE83DUT5LYDIyhknBujYt5xEKHeYZJZdRAT2HN
UYr7u6p0Ot6sZ7uqdGAX17cLV2DUBjL3eS30mElus9o5QfSxr2xYV9SSTfp6yUgF
ERMFuTSVe8H7CBmuCEHLrWXdeFnz5V9i2QXcMBItN7IFQQovkeXjOKoDkWmkFIfF
ljQa6OBHwLV2R+vshSghQcp76BkAFiAQJGgbbvDioENKNLJrSe7e5YQlPOo1Jc41
S5a7XIqqcmxntUIAj3txYq1pFulrRnXHAhybUe/JrCwiVQcYnAwu9aMLuYoQ9K0Q
1YKOXt02umpQme3eo+BitqqZoDSZr3Gh8YweikStg5Fb4BVj1ykiZZVkmKyIGqiC
xbSdBQ6ugIs7Uvux+a6SUWFxZac5XFbdG/mTbMSw6NOhZNEhjGkrjw2CoU9vAz1J
kLqmVIBaCj+HPNYAjSUqTKXEivq+Q4uTEFyM9QVo0LXBE1q5ZdAzA7rMWvrS0dnN
w6bMrHuSr+UX3zYZnwL5cVNZn0v3upYPsYxHQ3enS7m3LqdocaKdxPxakbhC3ihb
QPF3sisvpG6X6mfos3bgi6xejtk4H6pSZuX7pj3QKoigf3k1/cPx2g1L7JfQVXlN
vTX7/hqwcy+FFti10POUDgI84sYkhscjXZZklobajp4X8a4E/i5I5ub5JEguQpOb
szu2nRK0HPX0uayXw10dZZl83oDPgy0sIOmlOaFZ/4Cw0PW5ZDu4olzHYWz4peYt
DqalwcZ7n/YinnUDG+ERWZcz9eZC25neA07Kd5xemIScA2mNKUf+GNm456ooVHog
FHVkU//hqGoDXYJdHWkPUqIy3/CexOhrSxWIw0L33IvcLtEmFJiqLZJdaxQmiVZl
c7oeYqF58EL/wojU9uTGwjKgUAXnlmsLkAmmNyjrRs+uzcopAgpZKeaObejzIf1j
3sYphFD+Ioe6d9V12IbjdYp5tRfYQHxa8MeKRRy727Bxm2RGPXUDSHQYsaZF1gu+
Bkg1npY2rmBWWxNxxzWvAyxCewYXGkxmuTiRI9HjnbVPLNxfZvg5LIxJsCfFiPx8
hnRR0rOOYV4Lxo5YjQuwpnRe2Luz2TIEGavcAXnPXxfd4qzu4ZiUux8TKTE4+q4+
cnrhphByoNBYd73jZbYTCGgWmMIGQuK0SBfpKodkApXfSSTXGy54khk1qKmH3vx5
f5me4FeO0F9e5kRAyev60LE/p/lZpRP7Urh5dRBIgdy+mwOCe1B1g8h31kXc/Am8
wH2TLAxZa9aAI02cNKNwkMP35pU93aX/VEM7lv3KTA8TLjObz85OmkdP0/7tkG5L
Y9c67QNA7qNCyBAnEy3I30YXkcL0+TNfCsEmdSV5hmvYwc9hj5kWzx7eAZzJbj2H
DTZyOCcDjPdIH+JY5zxyvqsL6NUWRqlUDTqcSd1ckgnMEuxDvcugStN1KN6L/Ogc
kJApgIC7JAWK448a/CIqD26TpB14I2/l56BCt4v/O64ufaQK707C+GveJFY0QbYb
M1KyJZp4ltCUFuKgE3qYlMvQr9fB2fHBzIpPXG3qSRBTt0elnbNKY0ujBCPWr6xu
6R7UXR1wGdKeS15eryudCQuuYLAyghLBbIwndf3MD+cDFTYWpcGlUw/VG09kXTQn
SPyKtmhIiFCeMGoAqq7nrM+gMrdNW7j5uP4eB47zwSldypno9gi+ZDNx1cs8H6BC
Ga5F+N5jTVd5JFPIBq0d/9Q46a9bOe+ezHCA2JCUkDE2Qghunte0dXcac8oa05QS
ng1HLlBmf0a96ByAd1sP2beCwRa9eRUv3sHDBQP25MOKmg6nIxeSAJWvN3Y+ms2U
ye0PefKAx2YeVVPT7U4DQ0Yts4Z3Vp8E9X2+lAkXvAHQq8CII0yUq35XykQzjNUI
IT4eW3cpDChTUETjMCOGMyElhvFvwlLw6kvpOv+EDT7bwuIj6LLM9W45wIam7H2l
4y0M1FtsJYvrDvo7V9ycEriC+7XVU0/0x430/h28XtKqjjiWbZ85sJ/TBooVbMOu
hyTPQlX+2SaDHkjmGIVb0D3IJQg8xhWDfHj6t3VA4PRn4Fuq5Z7PAZemc9lLJp5l
xbSV6sOHt/QGELZa7BtO8eT1kslpi5Nl07VSoT5Phy0rUH3XNvTTcjU4yHYNyfAd
NKEBMpJ/7QCFM2wy7MJ3hZCEbK/90Do373p7aCaTiLV4THG+8dr87dIi5p0i29cs
l9xjpMEXSkc3PoZtS4fEeij/TJY9gAiuMURT9447yjFc9u8GELaZ3Bu9q85X6+N0
bSv0ubWvKzcOLsYhBucNF6KiO8Huuq0BEFrs4LlR7SBzcuNSdeOP2CVzqr7UcoNc
5Ch4occxkTaATcqHCl/76Hf5WIzzGRBHuoH41kld8Qwfd9ZTVpe2hWO6W9zB39hK
SkrKydDTBrqDeQZlqjhba86V7FCwAwHIQxih/tFEZACRNQ9JD7MQLekmqvF1rhns
8GqJqb6WxeOdZWX90m1Ouac2EH/HxGwMrvITPuuKC5zFYMA79haZaRD0+W652kF7
K45jNngT+TQNL3FHoaLsa4ToOJC1q0IIk8hmtNHe8I/Mh9sleZQwjz7N6iCzRMiv
CzrnzBuyKnEYoOpUBsQTcyVA7jToVyMzve+SGBe7FPughIzqsAYGhhhie78P6MG1
See+G8274/lujRBrfUJsdLBVGqZGIXaINHeSfL8IW6hBkDfZUghAlZai8QWtxOgu
hOCeuY1ve1orsMBKog5jRRoYNF1QkgDsmyGoRUrkkca/Xl2fBPMkGX2IcUwidntL
yNt4C1Ll/nxG/iFUj9R0fRFbCQlfXKhLsa+zIzabZxfWM/fSMvC7+Kh5xTn0gtyx
vnEJAAaFlsRqRnBxFLC4kynWvYJstBv5Za6SDc6/HXglADi1tITJsh61lTxDW5KC
PkUpShv2woNo6trBu5w7U6ZH2deAFiLWsP29dT+rnIYaZxtE/KDfyk1gYGaayY5p
mDi1aUrfsyfj3z2Fx6FTpsf/h98zDF86YG81lVPVcPgsSCfH7nSom0hL91akyyN2
iqSdTZ7lx5JcZjwWpjg0cb33BQnO3CvNzta/YWBkmJkFUONs7h3/v2gwDZl9DDBN
EO5K+cJT8BvaY9IHLygVbMX5zWU8jigX52M5E9gHaErClVhj6LQDGU25Ws1FmBrz
h0V/JhpTTpCzAkfjCgDLokcdCEPXbR9/rALMWiORg02F2cjPyDnorQ6Dt0YES6xs
bXJje+hR6HEG55M0VrN6gG9YIE9IM4nnkHu3IIJs3jXmi+X5Y4ND+uCDkOxA8zUi
iS8nxlnykbXh5ADXi3wSxp2oNleMKkQGFKoKiv7RPT9paoKqJzX+x47pVNeIrvlk
/v4uDQEOzYPPBHABlU64OpvYAi/mbD9Z/C6HgXu7g9tWvjMShNDMN+8czeZVKnnM
PQHaL0nTNkq8ipBM3ZOLuJwLmuJ5bBv+NA6nwJqgt3IAMrFeXKI8MSUPS4cSsDLC
QSgRIJhhzbnmOigzvPgNj8FNoi4UXHsiJtmcikfmfvlG0nDXk/Ncve0alLP/ferK
F3lrKFBokLoGt+8fBV2mCjT7689Q4weym/mOAPQeUCA0uhtAqFD4l3Jkd0vyWRvV
R3wZDfS6P6FwHqSzKD2sKElHDPkgeQ8uDRxmhLQtzodiw/AcJF63Y+z6Dhfvb+Cf
vybKA/jdyMYmDJguvwGP7CD4igWWHNw2i7yXjkeFsPkq5mYySwFcMHPwtc/CHIBA
qnRfKtgAlgXdGFKG9RcqZss8sgPwY7WcopnQSAWB8r4kF/IoNPY1kxDLjLUeGm50
X8VqEBGsiSvmkkLu5SgrK8wBPgqWvfXBePN3Cow+z81/pEueJuFGD9z1a016H51N
5dJvOfgwxa7+WF+trFKL6My5KBp6dxn/hPHbBWZ8ix8Y0apwR57PjaYTHeIGN1Xc
AXQA9sepT0kKU8VqiCQOnFXK8XUnvpy57XeVf/Gq51wOqiPJqzIBPBBizfa983XK
fsYw7EgIOPleet4wY+HD8syvFHzWld1dooZDZL2CuE6iMcgQ9oMGB8fCYlKuiqWD
bsmu/wrcDL+y7eWtXP/X53yyk0PsYerYIk9B0h5sqfH5jtuUYhxi0JhXT+wWe4Bn
0SUYdNaeg8D9HjsykfuTpGP5097ewrL5oiYAtZgvW1jDRv1iLovcU+lJ1winZnan
2SsVBfMuMQtUxV5u8lLRXf28R5751qzkMWdZ4jAK1+8JC1G1MC+6IGqH+gACu70Y
DMGSf8d03r3yj0EJn1EOBviShSc6SLFNlUoGYzFp58goZgqI56Wvc1q8AqyFlmkZ
JJptcyg4mDsztA3XFLDMpfWaCltsr2PVyRET1Ue1L3ZUuG0kZW51yDq3zH60p8wY
71tPTqMtNUiHkZ7MBEfzKZdcjIClkV17jDVLy42FtAdKV9+evQVV8eplMmb4upqG
lx8iLzpvag/L/va1ev3ztdQMRsuAd1Tzp4/Zuv5ZwoT+DtXmmn24rgEC2tKfq93p
8DFuZ2VPdKivW0XdgtrsKVifDG213KRTZTyPPWuuI+7WE7LHOFVNJ8fTP/yZLNeH
NazhnvdQn1Lpag/Ot8CE0QOS5B/y5JhdisA2klCZnvDDmEYtF2oqE87WOH3ZArBA
k+/qrG+Zp94NfMXARphkZQ6BaR35l3TuPvhzVb126eemiUXyTFl0Q+TIRQCjN6Np
8dYUHpmuunmRtJdJWAMfNB+qgZYrOPvCAjVMAv4H4nhnXogVsPkResYnn7zCwDcV
HlUnCkFls+0ypnfHvUgNpy4Rs4eKZxLRX6tVkr1XOH214s54f8ELF9t6ZYQh55TA
GqPakyMEAYBEXhFWfY2PEJl5Lv9cgZFQj6J4ZceWwwGiNmCY1qgKLZfmNisjWzhl
eYEr6OQkBDYEcLGl32z49Ur0R6ehIsEEd04SPko1APLobN22rGEvunV6mQVWSh+H
gkTVmhwf8MoZpj1UPAatHveqrfoWIwIppJ58VEJ5MSTT063oQQNz1Y42vthXgQPK
NW70nItbhAC5z1KQ55EcO/FGxTu51stP3yUuPjfysmFXhp6mSM/YVSYywnkYf7+z
UegPKM8N3YcbcFiTRsmPPLhtb/PgycSu3crvld1o9mT8K75WRsvzgHx9Z4m89qvI
hJ/dmy2LwpFswSIDMPGEq8deMleM3dQDA021bbtK1yY66OdOPuejUFwD4aUzR/Vh
4ZyML15h0+NT7ycdpn1DeysPS95rdOTuZ48XXx92KKtH5wG8jMbyZsz1xohP1oHF
mhT9YEI56jwxQVbewKN2h83H4UsNQx4D8h06Jl30HOMTfG1UsqQrXz22UNArpJPh
1SnPG5NzfhojPALgevzEFMb2yJIisW7gNzejZrQO1TLTRq3Mvm+/62w7LbWliE2k
bYIXN9Q1VNVihqGarHKBcsO6R3p4qWG0DM13letxHn1oTqein/9R7PnldHcubYGk
YHyVjGlXEOZ1TEO0wsmVjt36WTG2MUkTW/BsxyfM/GEJ/tpcoiarssV/zXhXKm8D
Z523+473R5DtNuyqf5PBWJN81gDSNMfLo7/F9jBnuKzg3AENefaVco+K6hN8GzB0
fohmH9CcOjFDHEJsJZtUBYsauMGyLFLmgEIrw88qrRNFDQ3xQKI0/+27TX/n5J5d
7u7/MoxQWg4JpH7RGEf6PdiZbd1COo7g9dHX5gzYzro/rW+n3i+Bnmehneq8FygV
FJpyQq9EFFiWswRDlzqs8tvxw1sy2FwWTxPSXkujD2geyRzt9TaTCLo4am7Nj9rC
RYI85nu6bpi9rfiDgN7iAQWhanCrKEWp5gGwcVGtZ1rcMX5Q+7gB/vDRyFmH/uqY
XsOkHDAIcXiHSbES8xE0krMyJu8UgmCqPaNNUTDjoN+0kirRXVgAN7fk1Q9Wg7WK
AIUftymooxeHvUhi6U6KlBD+mua8A2+dA5CEVKqzpG4Kxr/iM4YVef1V/Sqp4w2Q
GT/k7NrqjfOKLegjdgcPD6iWL5z2WHN+tayG5yKNQ9VZgBron8uDOSJp1OTkiSNH
TKkl4B0qTcPor4oj/U1f0sdFoxF7+a4i9HPy433MVrYf14Oa03BkgFIarUkwH22o
IUPmNfqT2UdFJvpNOVf5MCmRd6nYAE0Y7wB1a2B/eaVtA71lDfBNZfXc5geWYV1i
OnG4MKuzP3HkJiLqYU0yGVLEEVGyvU11dQ9c59GN5lPd/ERbeggIPF9KU0skJoH1
flrpi1o36Pb/BorGUz59/OBaFghJIP4H4z6bhh3+Kbpw8WFQfGU1+lrkyovEBVds
xe/1gNa8d5ON7/6JXFDxzZDF/kD47HV6XRRKzCpl44zVC19GH9j9rOjTMic3NMi1
VIDlWptIbQFslQDHACu6NPX4VrPQJGfsEOoqkvdEXiSlceh6Xlh6VOT04F+HgsPh
MweVVfbIuNwpHnhE9sEC2fv2kxLnPVcYhk0xITlJaNF86TIveBomePo0Zab18IrB
7adj+1M6EOKVR7bx/njMO/D4JGRH5Kg0M2nN+Lm+9mS0kaRmfijpAyu9zzbEQTqR
eepsSYCB8JXxPvLGejZWK7gwMk3O3vdyk3WORVbNkThRiKq6eYiKrH75RAfo4itg
gEW/GLS6xh6aeA4r+abchmry2kQy9ZoRpP30OP+W+gd8lZAmOXG15qIbdLT53wKf
PB1JUjv3HWkF1/BQwxbMtDV1bFXu55iFJ6tu1zh0NP7f3FoDFhUN5BcwuYJ+REX2
vL2kt8a6UANFEGOHWfNbIjkINjQS7UfYZMnNL8ugVl27dyXhYSPNNH65PwcSPwV4
s1Obhq6Di0J7IG+RMShB+a9RRtYUsdb/vIyIqu/vNSTB0d943uuiZuOuD3GaHN8T
kDw+aLWOaDnYMKWq2/wMY7VYVI9UzrzXeRo5csgrFSnapHEes8wHpCHs+AIApoa+
45Fo8oYUvCQzKuLkxebX+CXZdHVmsD+IJt0ssNx6GOVr9u+3TceWHv3R6rig5dcQ
iWpf8avrJSEeXonu1HDzr38NyeFrWPayxzHPvJK3fx13mgVClzJzo/rGPegdLZqj
Z13eTawv22YgckuBkpFFFffFUFi5Vhc5jbqR4Y7M9jzGOVxTlybV9xVilCWH4DXJ
UnTegLBtVog3n8Or57i+MwIV763gB+8l7FxWAgQ4aeIJINFIUfQMPoc/QqpAU8b3
3qcThwQbA61YEc0G5AA4F470x/m4+tTgiaWLVNGfyPQCrQ/zSxwb9zF/0d/lbTOz
DHadqsyYPJx/tV14Kn185FXkEL6/U57CXJNaBRd8a+9BfxULBYillY3AX0/zSaSr
11nV/BAuxlPE2+pdlwBXbv0jjr5LeGebbU+XJMWWirwbRSep5Et36JH8H3PiT7N/
V+nSAQW/8Ru7xoifBcMQsK/UlpLyy6sEsxH7m1F8mePE1QDrWZLDsy99slYCbmWo
fnYQhSDPR+BC3w4N/rTaHqvt34KB4DM+B8R0HzH/OwAZZnrMMCFTR3FmD1RtCLko
F6uxNT/rENXOw4ehs914+xLMLq81j9J0TIO6cAsJ3/oSQJXn5bhh8Q59ohqlh5Kb
l8LG2GIddofSgsq9xrxGFDb5BzbreLqT85o802ybrgI7xEupvT3DyHBqqXHvlmhI
9oXAH0yLrwTNvEdxOLzQuGTKssDAkumLaLP5k4cjsXGRPWV76vCLG16zvLrV5QbI
bBYl114aD8R0SdGXgdRIO7rYa2XqS7SXQVvBv20iOrvxs1SXid9UvPIKhVYrevH/
0Gb0pbg1ehLjre28d7qRgYoD5ECKrjKgzC2M7Jy/F1emciGDaVisXsqvOWCTd3qc
iI+jJomc+ROhDmbsuj/f6e3hlxObwtoM8q/DNoxD4TwgqU5xe+H0CI+NTJR+5ZTG
hdoqw7mFll/h7YS0wxJo4FU/h9+hr38J0XL4wcnWpp5TwCU7I6dlSu6DCCAc/Zts
gdcIhJNAhkX+oXRJDIVEdteZwXidwe3mw45Tk8wG9SLCOfQQbV6fEnU2SNPcG6BO
BzYZ7+I5Vt++JC0e295vfergN3+li0owCta1c0AusZ3Wxvn1ExDcV2WeyQswy8fq
PRDAUS6ovpgXkaFPNlMbDHxkirzkX6GPAEBG3pQS53m1WAg5R8aMDesVOwdFkUDT
goP6WOBWkFUZUpgSykNHcHoOiq5GOtXXnOOBxal75zSburLgs9SA1cpBalsvGd2I
nCXHEIIKENmDrMOn2j/xzWsHNTB79VhYXf1+pqXxkKEymaoABYu3HqePxoxuMAgw
o46VzZkI5JqipRYBx64dT/QYGb57uEYBilipU7qug8yvAtQDJBoie3lgrZQI8QRQ
zFs9tRxPqx84bd2Ze/KtDluzBI5v2j3Ebny6vT5prLRB3dIfnShYAIWCey0IMMuC
qO0wx0p7s4Cf2s1+2Ng1BOUxpZUxaIiH+ApvKRJVxgd4kjevfYYHRlFJAZBs3Lwv
j+wqXPyUJ7cSbezcWLLzXYI9y3NsF3mZ10D26RovKgut9mkOoaRQrmpwY7Ydt5Pt
7rb8dscu32v2l7dpxFh9LLOnybBs7kH1TsHMDjkVBBknTWswwULYQaO87IdUlRsB
dArOPnQFzzfWB//JV3EVErPCZVw6/ABLexNjBWyKLv/UuLWNNfVsekzoRrzCqRr8
1om32pVaSuFFxCvebJSr8mOC+um20qzED2VLDgbrYxlPeq5URdQPl7ewYypl0Tox
/GHgUyx/tkVOiF/+PC6C14/UsbBuQKYBt1Bnq7YBy6V4OYPb2tMf//W3nzZRMI65
8iC8B/AcKEe5QnGrLsRuC8bYCQge9GC0EGSSEdeHEBYvV7ZKIc4K6A9DKqDcrbkO
FGGW4mVAWW0Zy5X51nCKR6ktpthT1yloKhueyGyGBEcVrRd8fPAvenJIf8hTHR7w
I4zneX2noTXH9lXxM9aQ2WYQgg7nekpNObCqgDCZyPYQBgwdD0EdGu84khdsAcN+
9pN7hdtPMVZjXBnidSEP3kJeEXW0krK6FGDopmiJmJvUGTf1Z3v/be1VC142+wsU
db/Svgj3GdgbX0F5Vykw+Lkl3E1zevJmuJewcB2n3ReVvskh8eE7uBk91bhRPfAo
xlyIo94Rg2HfOh6AnyJB9ATuXW2UTVhmDxqIHfEdBqWRnRq9qp7xBCwtP7zbUlVQ
0hNsNR3cbkRptI9m6yuhMB+EfXztxSQpeRmlk6CPVc2B2KGG1T1hv9Qtp510knAz
/mDnkmW33jhfea+oAQ6DpVt3vmo9TjfByUIIs5RPW0TzsS6S6kiW8eT3XbSZAEMQ
RwIUtUnxV+6uW+NqHFj5fqeyNwpe2eKOThAaTu65wwiAUnF6q5r527N4CZZGfG+b
ehHxNYlHrqksCeABLqXMNNJZfpTmEcrpyidIzCZ4Qk0m2EbdLWSQP/g0EMsIctG+
rihtteyPtTE5mCL+FK9OUmldqxBB7BCNPKvy4bFhIRx6p9lcQYEvLN3ckF2JMzpK
j58mnL8aqIYgrfBKh7de5liDtiUSO1OH0n2qRHziqPtiE8bRxMYUWcR27bwvKE31
31lI7cuMbFIh7ruxsZUV8nEi1AfsXJTRW/z25GixEnKR2x2aQCoUVkZs8eVYDKA5
WjwvXCdIb2iWt80H3HJztIDckjLoLSW0KU1wNry4KP8sXwXm0Sepz0XldSsvgOfc
N0LOfFtTaQwTpmlYNGSqRSHMM6PN0klz8P99Ak/geJT8ozg8gOwjYJ+Yv8/Tsng0
MYFkZ99PcvsF8vYCeoVpSOX8NsVK7O5K4EYD1yN6rCbonD2alzzp6wXYn+8zOUmL
B8Jl4BMWl+i0HIvyELsQ+NXWx+HEWJdMIp8BHNNgH0AIutLEF2i94TvZB9OWd8fe
k7BSr+FErxgQ85lEhC3IsIvP3i2aXQOJTOWeFvTGvcaquoIC4Qsq1RGzfirxHxwj
nescU25S+bRMrb5URjNIfzi1/7bxePYTSBlTbUKEjey8WXoad6kwLBrNw8cma1KQ
x+rEy6+Vhmh94SS7Z3YrzU6YMJCkw/eqrh17diwx8vQZn2RLcrp2pY6p8zlNGIeF
wWqGBWOHeu+OFsvvOrqgNLVeWQD4wA5bTXzmUIIJaY651ClVfGpCn8iJlHoV53Wb
ODMLMC9tluBqdYOWl6762oGp53s7Tt99wObE/iVWaGRkbkx71u8D/qoptUDeVf7M
6WAoqXuKEo0J688SwLRwGfgpjsBQeufwvtped3VzEfQqQDJn/BTnAbQZQxsgBtPI
BUx18/AB3p0G9Uvs1grbXvedyCyFuPJ+gLbtcmGVFwnlzMlVstkolcMyYMftnrqU
Nbl998O/6yp3qR+4H07WSy4cUY/upjWY0v/nZ7o/LQt0E3tvfJQUALkRO80m7gF7
Gg2k+XYyiOo83oc2xQzD2kTQ3MRM9lzHtiANwfxctAVvpmo6V86kztzTmyFy4Hzt
3oEBgiGl5NfFLlHSXJmX+45BhJqeO6Kajk/VTh9Rm5bW15M7WeXQ4SePcuvoQVyK
TNAHHpiqy5fxwHrMJz8Ppelv4B/CHZf8pgVndJ9I18nBtLsWYlczzV39pp0+u+7C
ZRlSYFuPHBMK3UWaEZiVEyAl7mnt5f4S56ECIkEh3Zwd2VKj8DctZ6DKk2qBmH8O
I0whRt71Sh6nv4A9bhCBzl8boKXuwb4G8UFFYjNdHr96DJKa/OOVDz2uKPnT1hsz
MtA+oqwBhIj5OsVYGAuHE0CUrJYtyYNyA1EUxNG8vh74ESzYUvFMfZersH7+pny7
dOYBi4AUme02okUhwsP8oIvRgrD72CfV9kvLKTn90iDviKtZL9qY2PWsFqrPhJqN
j4nbi2TChPTwkdlIu58RANvG7vVqXWbRC91Pb0k0bZqKgldOHj3eFUIMCg6qUTnV
0Ar0jf9EKgS0uJxx/FdGbCc6KpJCo6/XX5T2q9DylMlIidlkZ7dkl0tJ4cNpXalj
xUW1tDJ43EHi617bG23WYdHZrmKR+Oh1N1KUwaZBMzyOT78ahVCs9nCwZv2pup+x
D8vYecJ9bj3DpUwPICkVjmdkWAirbmIjvXWDGEfbkzO2AA704eoRSDGX8hqGt85S
z0jOKVpJ9+yenP+kbOfyRHYxh/k3dwboGfblL/9eSZwNGQbju3Zjn7Xcq/MPgwTE
5v0sG5JGAJTVVmd//ZS39l6Ap5iWQwN8WltC8U0sUpLkgO4JK7LZQ/Z6uPx+7fDv
bY4f72P7o9J15iZk00zbfQxkdQAKfisvA23kAhnzB+ZFo5vdzG8+rSx7WJzI7WQL
s0QOY7YSPMnjPiCM5OdOEHrysCO3Tc6xaPYwhyEnNYCMzfuvpIW7+/i44cT1F94c
kCzfY3vSiWETGDaVWthT2KGNr1J4gDrdqeHp8NWX/FTmhfVtL5D1gwGKnGO3jrsV
IN56tyZFROXKMnKuZZ0+Q2qzuArzuaNfnOGB3lB4wMivDWNyDfeYCKepCUBWdqgo
boQb8wb1KknXSdNjrjAiCpxE5VYxDMRIZF1+HXBzdH96QD3oc8yKWJQJNgDzeWHt
1nYguedczXXvGeR2sFoZZi+32NN7MHFXTTtuG7WqwHLDWUevD0RZ6l7YW9zhMEPE
rJdwJa1r+RA2RN7rSsNPJGn+OM3KsP2AbaPTT9ssenUn3bPXVeWCcmWC051KxPW0
fDGlwhAtR2fQmMubYQPAI5toifhsrT2ddhMS1OdOVLPQ8Vy13pXgWASG/IB2Mj8/
3QgAGc1+WYXRqUlKCxBXaHRjHU6eLq/wERJlrWW5oSwJQOCeU5NilzzOMsKtC7WY
+INvbv5feREK2ScIe24g4YL6ayUbDZn3smFxLMVfoDiyTZf/ZyjjLMBt+Sg2eVHL
trzxIybXoR1rCPyCbmaYxY/28ILRdSVEnH9BQyrb7Tr29WZ8AFasQB3Bj0Nce1bf
vuA6oNZ3cBVv0lSN2lRtPkzc5mDHTUovV4232JMCKAbPsT9JqqxpJvqPmzC12b8V
6vlZUtgW/9wWMQirbTbQ6MW1Ulxw2vQXAmu35isGVNRo63B+mW0VleD4p+X7iYRF
/9RYBgWiQ56VDZBS6a/k6UgW5uQZz/8byu2nzotyhTboJLyuIAK0vbrSnRIfryKo
eN7uGK07d5Y+qpuJNJhXcs5mRwMqy5r4ZxLo9uZ/5GOPWwrVbEKlq4tYUqR3G3hK
1LeOkNmnd4lDH5rar0ysl3I7yIPzLXbj/7JkbJTygzBYzlgbNclBFNxrBbS+jRos
iUplFAFoH+noznUhx5Rg0tuj811aHUZM9OaMKo2TxSp67xif3sLrdl3fF0Ols2xF
DSqAhtitdLeojS2fWojavZmYwPI3EkaKxrZk5EmXa6ZIbRaO0+SsAmOIMDoxLz86
oY5DG/tdI43HXJ+SyheENrvF8qeSKZ3bvh0j/7ZkolsYfO3Rq9tGybaxUC8qxSdH
XvJIbBOyiw7WDfyUa9EJf0zyhfil/5FJ152pS681YjV/snxtcHNRsXpGFcX3TbGw
V1y+Q2NkVlt/jJI6IfZUPTEHW99g8IscQkV0uqpV9BJHwfgM/5TlXav+KqWrMVwZ
ngqbQOD87yeiMA4L66V2JKfj0MvGY0MFWg5M0z6J/HrX/rcnrWDIiqLPnsd0Wah7
ew055dnXq3yQiYTjcSWH4hp84+UpJEaMTo0+mk5FNdVEZ7s37IUUvhBYHCrsqmIi
WC+EapjtPXcgvi1gsX9+JyEG19AggkRhscy/rMGyWbw1lsNOSmJ9VCkEGtjzTuk+
rdV1jLRERrExnsy4FERs8ENLZcJxpUy+/rSgsK7XvxuQ4Y4nd1Ao2jrwrTyt/HsW
ZbWgjcrS++pf5idWCsPSIzuvhUeTFCrc1/CTZfK8v81u+PMopxukYLNRsVI8UR71
6aP9Kv4XCdv1kWHg6YVscYjOO1JtwWsYIsR66/qLS1IIJsPqCQY20wByVCRWJY/N
jOLe3j5RA2C8CLNPrwyo97lIWDBqmchjs8nxtEVryp814i7W99f5gDnXcPCfwgRI
qgUVAiiWk5cKbvXhiyjBpd6vUxgCahoaJSAQJtCCpoMMFwb3h6H6+OW6UdFly4Vl
rHRDcXH6aUMUcO9VDzAEuoXMoNobis7X5mvVyqIpuPGBkJApTFVXl5rxNjt3WwiG
T3Gf8gvADg9gtc2Nz652zXbS0Tdupd3DYIFF1O8GG1n/9ytKd8jOqdb9HbO5SkjX
VUrHGEBGYuZutvdMp3anMFFtRKDoYLgON88UNwqn7+cOJINgbbNKL0x2ldoo+oi6
3FjGYK/7LC/a06lTM/N1od06dnWGNJywTxF+iDRei9Km1p7zBtBF8mckwtDJBayD
Wxe9Yl+anR7pwTMpIR1OjJmOViYMzElYPctL0n7OKpy9/FBbzRoPNBPzBBt7eeUW
BEtPBvhi5eclR6MhMuBAh6pq6AYY48RItOnHe9p/gC4sJqCQyHGYvL7YeBqmQR/c
yJ2r+iUq4CVOlBDeuE/WqYfwfkh8hm3hTkuYB9rLAJ9K8HMGMPh151l07r4g0D/1
HilsrvKkQb3GOuMcpJnBcAMvCPZICTHVmNFY1xO1zTFCqQFOkGBt2DBl1A0cbkiG
Zke/2aiTlhiq9NTdn4+Iw+9DDeBGrXNz1XAlojxTp442W6vNrQllSO6pJ3FojywS
/X0ACwVRZpHwZ4tm7zn9qwgLtFvsdA9pLZJ5xrMSvgO2/wPhekpXSjUGD7V+D3Gc
Lh2SFq2rJbit8UG5X2egmA7ArrxnKu/IPt4NcL6UWTBDPw29jP8O68EunvmFyegT
ctHSOIyQ2nzfZVjRgMs5rXN0F91VbQx3JKzDL9foTlgyctItl+iSltnnZ0uUSv+R
Z3cqrl6Y379hVLWdIZq/Gfw056LiHVAdaGTC2bENVziCJ8YosUJm34IQlU1HKTrb
8gnOgpA2/3JkqV/j9xsaETTqROtjZp1ZQDMolIOnWS5Ek1jxJNhpwdH959XD0U46
Ik5eMCW66BVBidaz0JUnC8pfplYmFHqYlXbsSuX5ta74bu9mdierzOXjmMK3ETgz
LpbmxPJ2ptg7AzFSxelS8FkiMuZLvaBUlphT34pIaOQDTqlDsGCi51EMloy4Luti
UQZ3HO9qVY1TQtFco7bbkJD+NuMefDbKQVLkYKle+xboJpK6FIbmU+ySD1jUtwTS
uaNn4biwP7TwUzJ7XdeW+MkE6xpJ+ik9AERua3IBKVHc8ZH/OoPi3Jijy25yTUyz
5hD3qveo28PAsSZeKUugzPutWKBA8in09GIbHArGoxImeYJgbnv/VN0YzGIuBb9R
X8otA2ewrOlKjSvfQVHjLeQCc5j3yY8n5/eV/XcH5DqwRWvV57bziD1iTnZSeecj
Q4+0Vn3skk5tgNkyya5SzsSd/vF/74rKTxr+kb1lyHF3xRgex+EuTQeJBx38XRxq
cm0b4lmiKjZr9C5Qov7b1HLUFkGeSebBaRfXvalm2FVeBzajR+dRe9H4TaknV8nH
htSrX1n26HJkdl9YVRxXrHTe2H0MKlzHpzBBppvKvNirx7QOiUcu1BmpcRQGIMMF
pNGSPf9rn6dvFmCE2x4set2ENKv9Ww0Rk+1nRBnGxkk0hye7OytNbqScIpCldybR
nV6Iqrw/0SwNZWSEkWJvHWAwNEbC0dTkihR8fPRxObLeaQrN3nnpEJ7WoIeDFK2x
OVCQB5MEOEYDcqLdzhhO7ztp5my8Hj2RzdFJY/V++IB6YwOZAw4Y9GBoWl7/VxE5
FeHwmk68Yc8V9caGmtwWTwV6gMYJQm10n4DUvmgWPDBL8ChzZCFnl5mytW/Mco/Q
ElGL0uFuA7cmkW+bHKuMtV420pOEY3I2jDgjHUPTSU6IcZELDOx4qCm5f2VuRSmq
z+7gSc6K+4LEnq6/hz9mec/QLHHW3fsZWY2aiXIabpGX9PppyUmsF7CSwbIG+/dI
wCVdNJD8GDA2eK7/g62hDq1cShg5PcJPxQc/AYFfRLcruagSCjZ8/hpn9K6OyAoZ
02VtJrCFDCzRD8VDun5j//lL8S+TuHHxGl2oNUCpFSOOTIi9Zhje3gYlY62/rT2X
CRa1LeRzapjQmdGuPSizYUQH4aDCvG61vLCkSZfM9g/EqlD3E1Su75HC67Hi1rxg
YbKrlHSBWjnuEW7T8E/vTSp5w+3xBM6YGWd3PdIyAwKCgGeo8mydtsOx6wo42JS9
Ts+TEd+OqV28yH+VlzJeMSMDYC87YPdy+ntvSsoPuLZSMFLMRVuS/OVHnjLcuwvm
vYdTj6t8wmZJJQIAgtjN+u34NCj2Gd6HM33oyvo9qGYX4CKVN0HNsMyOpnvr3lbJ
ynCAVO6YWZbP4t/YzmZ/YFZhzSn70kHVHGdg+8v75zzfPeaU3uFNnhBFmalcgCfr
7VTaMGFlSECc8pUJEy8IRlgpfdYAg/90LLRTW/HuepKOtzzabJjSFzD5IYObwibz
0TBT7SAtjlQdJLKZ0PMEXiGTY/MgCugrq8PibNodan6zMv6zyTJxrEMQFdn5Mc8w
XOnZKJWwnbxAR04xHbDAC2jVgyM8PSWqDgWhDjAKw2Fm0FOzJAAVTjG3ajm6va6F
IX/MJPSWGLLI66gmjhgeU4/XvPcuQC6SqD4SU/VCrwmKqCnrriDG1ZeZc4FYgR+p
Xd+rYGmoBtDU3DuLBirWDZGqCnUYGsgis7NstQy3VeZs8nGS9zBsQBmn+DwH6xGu
F8+aSaXH4ms2S22Lg0FGOwS3jE7FGMoeb+nqJx1TXI55LxU8MSBJD7hulk3tunK0
mOK3lNzNfI6Nd3OVgwh4Uc2H+cSxfVX+RMItQvmhu3juJ/Wq+TqIbaKlInWEbKEU
48szZLkeEjbm/luG8JTfe0EQJ/0gClmFACbYb6z2vvWz5g1WvmktxqsyCnpr/Dn/
26Ji8a1L1EnGfFkCwty14cZmjN2XjIgImAefjniJlW9XV2Miof+CWancQY6myXH4
kZdap+UhglanaGXajw1IgbyhhAtUdF7tw5NBjJvNbotiTNhSv7cc9BcN2dD1n4vW
eKXm6AGAdFHwIQuFWw6CLIkrexhGhL8HJM4VIE0Hi3pOkLoNDHD2skPUxEKEbuTs
DdgzscxX0yVA+7KkaSqSPh5aep/94QCP0wQmPliBVTKYg2Uavlv2u2IDF//nyjS+
Dj7hqcykP3/LVrUk3aMyXh125ajMg2L0chTyTSCtSVNYSvEV7eaO8guftpryF8GD
ARfCF/A3rao+NM3akbC3SIsJehVKG/nYG6TEsfy9DSBapIRvk+uTurDvggibDpr6
1gIma3HX3jPglL6t18Or5PRU23mkdFl77lwgUCgB3Rvm0g0gCn3gLqMczpI1mZ5Z
ge1DnyaNmeG/kaDKxBa3PeB8lPcfOI1MmCBSNC3kXs3GuG6DvAWtNLXmaHTrvvDo
0OaNsMRmMRTJeTd+h9bs83Fba6AYr7m1Vg/4Rv4bgPDuv1N5YAm0OpxzyFT2k8bz
X6uLwwC7dm9UkgyELhmNnLkKxadq6ZF5HSzwwxv4HiFBrziVWgHXeverv9qpeH1P
BnD3DoQ+pWqThv+/NwqNY6fECdxoh/DQBc8nDXYI11ItwqXpMDWzvMzz9gLz5f58
3v4YbnZUZLBZ+Ma8M/lJJHL6Qx2ySyVJy+Vd9PTNTdhRrs+pLsZqVPK5dIg7mBhz
P37ljIW4OK8R4topsgrHQsVUFJ/T3ypXB0Y0epSKNlQ2VJV7YyxNb1WyNYHAG0y4
mbxir90LR5+b6EZiMJ5OzfNLTjOjZ4tnihWVhfJy/QE1Q3A3QKEryntFJ9p4scDz
gzTAGgqeQ5l7Eg/mAJLVbtyfruGpw4sV+BmI1q8ccccH7GhfaX4u/lfIOC0c5Yok
KK3+OqoKn201az7mtkdQ8BMnLvSoJjOPMRXUcCmK8D2MkPGUWR/ZsGEOKtvD5KdK
xHEUVP7I/QMiWtS/5WxD1AMAI7ZdepNqz06XoDUBB2wejJiSOZ9yJeFrkQRYqFOF
EVNYKfLf8au+xn1fLVnUftGk7LYftp2zVDDaT2DbsolXsH0dXQv1LeeOb+iWSPqk
m9V/DXnYmcuF8vJZgVK4r3X2+bNm3hANeWawxdLL9v1vRA7iBO0O3xbZDuW5IbS0
Y+4JGp6pPBLQ7GTj5aD0NR41BrQLYft1cbDFHXJcRkrheVPZqGBQJo/BNJvgR6lp
6kyw+Gts8ksWpCnQoNglZXeIPTKJgmoWMKvEO/IFdYlMAFMganBCAU/k9hc0Wlx/
oJ3+vYyO3J26iupTE0ENAfg26cyzrwXk0cHeH3aXdYGDe5qmSmR1rDlZiZn+9N0P
Pv0OCb1mohCn0bwI9WKu/xAHOxA7C2CPBSUKOUDEJ5n8VW6YAyrpuYaEOfl7BJ3x
m0MpzBpAYRWc33F2dIWNVmDDQOukbWDL7/ahKCoZu2/fR0Va4ak5gp+SUpqSY+5j
TM3sqCTeqxmYN9YO8H5aLQwmVshXjuge+4ki+XNGe8jqUl2p9/lHCUcDbSb21aQX
mQaGDdwFQ1KuHOnQcHX/sUR1ypjxtH34Lwd76a4+8tBxCl57AeWMSBTcAc5CbjQ5
750BapBVkeXv4oWWNcsdVbuikTjW3uq3M3qtSHLujcSQIO47GQJot+BuhfOEZP5c
3eDZuaxz4nPVVLBPnb0YxLIpD8XPbz9kzLDyVaUc6JqloEoe43ss9mdOtJrMxsrH
+Lnw8z4NyRtCwtDinT51zPbTNNmnPuqS7G3otNgxnQ+bfOnFMmt7R9qc5b3pNKsZ
R7MpGbdbWMJusOQelsaXSHHj8gaw693z1OPMVIDnjuV/oFofJuKkLrEOKIk4Siyg
jASodQOC1qBMAjBGBIFLZWp1WY6m4bkLlaNlCPT8pNR0NHffPBMkjG+pv/l6hibZ
bKTxAEZtsG8n3y54iZsJ1usGcsq40cpFSGeG/k4Rs/ccIcEK+cWWwiqSKU4Prhu0
Y3m+TIjiMH7VCmpSgFu84hdPhCR+cFA3q+CVOnsnR52qKJRtftgFDTjTIB6q8kwm
IPkFOaHoYMnDvWqxzGUFFb+0uU3LqpfdI1FxcgS+yeYP8Po0fDzfgJCS4zxY4Vzh
bb2HGHidMXzo9kvdHz9sMG43fBK6BZJlDpRxLwaBQIPAT901KluNSyLnxY1eZfUW
V4vyWr71sCW21w5qQSclSXQ2gUx4cdyy5AJMewkQHa0kXWIsFq9c5XXmU6Gvct8o
igCI5YbAcHdu4kEXCQS3Zc343bEOP6B9XjNwE3BB4rmcuKcOCnHrZNZiaRTilax+
fsLIcgT5KYJmIKICwRcFLwDrZpynwnEKZHGwVBuH7wM7l81jiifXgHj7LN9tg8j4
m3qEPPLqr4PVTTmtGKi1Q9M4/0E38UM162fmJQUgeCPXHA7wlmaUi40ztv7S42zs
FSn0Ud+mNV+kx0mLxMcbkPvEhSCY10Mvo9WpDuzqT8XXotrXEgc0GIhL1QCgW/Ww
g7R8PzvmxHdDBNuupUDggRsX1W0HMVJCD1FOcH/lKVzIOSKl/sva/crFU9M2JomU
tFRQhxBv+TMuFbPPGyQqTkQ/8sTQdM4PPmF0ioGoiVGVSxeytttU88UJzixRaDLD
AhfGNXj9JeHiJ1UYXLHHAKxV+TjEOdTtpEGX0k2GEnXooGYX350Wd1NzrY54s6mQ
hduBlGJX4V/Rz7NQIgpyL8XX6Bpdg7f5JIg/iTWJ2Hy/b8ZGVfTW3m8PzdNZX3ho
MlIVm2JDvNenJLkWgFcXQm43924ex8VdiezwJ2y/AP8FqQiSj9R7oL2HRA8F6Q9Q
i0hs21+Dn89PZpWTsPawiFeYyaEyhPak1cNZzljq3LdSSdUeB61/c8gRIZdkIFdN
oD+vz9krIXlkfTawfZQwxoWA5zMS/U1hwzKzErd8QqWIDOPwXWcR4yws4TaRp8An
BzCmb0FI5J5bpnY+9nI1cqHHAQLvcRZcXVC41PBNeNBPzyZsD26rVq4Dt0dj8bGi
aFDIHoPoYTpjY7gS1+LLz1DGJzDnnSfV1dlqjevPPXJILTO2BLjMmFZ2Hn6/a6jM
BM+5VCWWCaW8d4KQXQt7HnR/+oviJNpD2KkgVD0AY1eqJIX5IcVLy5hfYoApyWuS
PXryBuKFJzEpfjdaaLZfVQDBPKlbi5bKzFjqP/LAAz+2TG0OJiMpM9vwwdh6EjN8
7vrjVDpZAsAMRN3+tt1V0zqOdOhAjjIkHqlk8Hoiw7nMRVwCl3JYPLh4Hz8thOio
cr/SieJaM5SzCsmX2fAd9/G/VMd9ji8Ko6mHKymThPzHfAyoeq5HJ9inHBhX19OP
5VyX2c6uniwTZia+WXBsaoqomm9iPg/ONp1ravdgrIslFecsQ9BAi3Q012Xtteg3
YTKpe9yiKpdtK3n+3XOSCLi3B7EmKL9iGeL5/stw42KtWb2bweOBSKKi3JI6z5pW
k8Szlddzev53LvIQ9v2fZ7Nh7K7h9YwThWFd3HtSHtYIoDA0ZQ57NtgksySqTleL
r99x//Do7YJ9Lm8LYt/bxR5q30lV32xT+Yql9OqUBEKb775XKbzDw50Bvvv9KCaK
foEiOlkO+q5JzvhKT+Y8CP0oiNeeOFCwDhvEws0+K5kSyiUC7FMH5wjFjCjZYzEo
kcP9zEb2Raunakg3K7WQbEDmkTsquMut22yc1/NCMyop/StlG0rdjHauRzu8Vvsd
4yQ6HJFPfKLh8k5lqP6GCgIGyngvYsZCduoS3RbdX3agrHHqjiRl7jo0lz45GTTw
2VG8M/VqhWm31PV4w18WDoYJU8OXzxDtnY+5bXKoYFSK1RVZhKOGKF8f/Bc+UQaZ
K36HKyPc4lNNiO1EQNClqKZKPvoF2T5O5kk1gJbAsgtGLR3TrDu78H/Aa5471qN2
5uZeC8I1Txm7vNyXw+xpNoFY4ytMPDg/rLoCo8lAF0y1TIdsa8k79GHRTayDpJiB
u25NL3xhq8Ijl9zGHXP8RhciI5C1OWE8lhrWs1LmYRE5J+6OZE7x0F9GKJNLwH/y
O0oR7CFlCq//SfAYXJwzRvk0ceSALJGjG2QQBfDUk54Ennk6UZ321HAMTbfPJaSJ
CqJS+hvghmhGkgK4m6FDyqLdHta5hakp9tb5Qw8YDUzYwnfOdPZxQv8fA1kw2ruQ
jHZASHT4BNZQZfX8TVYL5fJf3W6YDDj/w1YiRICgWXrc99aQsGeykjPwWgHLbwS8
V1bykTW9Rov+3g3xM3IcHbrO/FXMeCpJJEIrwbs3WFFITGT3OIsjKIZ8ZaaXLInB
uJD+L8QsXPZJ4RsHXv6CajFJqXfZZY+jcyCtRAsGFtRg2rX/hsAMl0fiLuqChJfR
E29dNCg9KklI4mLjeiFzqWwzdT+DRT06v67wbyoLGazBtiEdCMCOjwHgivL9ky3d
mzdVFLruzWqeBeTEkHNHbsHCd9hgXh1OyAK4FvriDMt8UJe9JVqAlj1H3A9ffs5t
xPlka4pi276z3u1iUcN0WakcRbWfrJxdATrCeBFS6jMYkF8Nb7zWC71mH5XSEvVx
FUXib0nfd3FWUQaSkjHgaSqXsDyzL/BmsKNSvBZpTDj3S2c/+eUqlerRb4cE7xtk
/3MpSoZFk88XknxkZEKjaWcRCUrD+KHFy9Dn5JEjzn1euUVJM8EHbdny4agQbDra
8OcKWU1doZPwxOKg6W3DiU9okcRpQba00lZz15p5UQbKKLax5WIS4PqaFM+j08vx
+pt4ETeQe/97WUfT5miTyvWnquENN1eqWzTjTZFwt2f6omdg9Dix7Kz8MstfDnKL
xJ+9MRmMlYk9q9uo4NqV75F1LJQYP3GjZhjn6vHu85MoVSXtYP+SbdQ6qsCSqXJ8
WR+sTBO68es3wVUY9G/mfQQh3ABpa6xyqMPy07+f7hTuorDO1GkXV7eizXcyuxNN
iqPH0j0g+/aDM99xilrzBjrfTSPtV/fwdPcsb7/KEmwwnRyC2pMscA7IWDVW0mXR
AcXJwMh16eILX/cx809KrCpHSAxs/ZlaOV8iPdnHgHg1u/Znv3Vy1Z9zVVlHrerH
4oOs2aGLCR1by8KC1UTwlKfKKfhV+yeeXxR0cIsmQydIBqe2L6UKCn85GB8LJUq/
PEQnY7jezdtxoT4Qo2hryIyMdMyqJjcM6nq66aLJsPGs/m7UphfHiyFtr8Cp0aAH
pfPzDS6gNLU6KG4P9nQSq/CkfeWyMkRt1xCarQiMa8ySbpEGt/8OJG0QsgdZMS29
nvW6EQg75mh+xJbe1tofJ7J+gxtA+VrBCJ1vVQX/bVG+caiRAhXBuu0WNrMYBRWk
Sbdcx+c3GK8SwTgd7uB+fbLqAyjI+T3LKs84KnanP4oh3YXhZ6Ts4/ybBWTZGCfu
8rPBeV8It8z9Zd9zcFVIkXjbHhTQqOR0Q8Qwsu/c4Spl8Y96ynXxcsnM9U7y/TEc
Bmy5tXZsjCECdfrQYRBPSEaEjKjrw+iCLb+ckkd4iWik8j8Nmk4Rir9HIl18HRef
G1rYY122VY/1t+D38Yiua6tlYa+TmmHj0iSFRBpcTH3nKpnRRG28x9te76cIr8pN
VJQnnZO8LuEFZ7QWTLzsXILVNbO5hhhpF91KHQcv9wZGInYQ0cQzGkj/ZIPgMfSM
sjGffH2osdcyPNLIkggOzOxew+PDqYZINF0aHdf5JZsidn/6zVm5DXfYh3mDWjdg
G+XEJuhAKV4twDeXiohpuCannQHojb5D8m/U1MY8hgekzVLtykFjXymWmCZkNKcU
s4hHBbsNen7d1JoZYNiunpFEXFVwX0dtEtm9jftp1MHldWIlf0GAWNe44nDTZIho
qcy+mR1aJ+WcvHPvtPEkUNpao5k1KPwd0MgKssSx+J3MyHcAShbtuB1P90BR/Ta3
KVrrGe8vQ3tcE5biy0EBXj5mG+Z5b7bO584phuRmkfkCb/dFwBdMG0TLnzipxQQ5
vevIle/lkYBIdyzwFp+F1D0wZEEM6IYgL3WaK37e7GaGZ7+JvxW4RBnV/kTQ/piK
TB7B3CEVDVm9oHFsQadz3iD7d/dU10TDJtzkoU+NVSijX/e5ihLaOBcqREDG/SgO
PI0Z9e0Zbi8jDnYExY8av+AM2w0k4ULmtCJFsCRf3LYz2dYsiaYOJQbUuzkQWlNJ
c/5gvmuXyUx91PD5u2VYa8YBqNuNtQe3Q4bJ+Yb1rfStDE6dQH4efTkrpUBVUhtM
RfFC6UkcOzWgBgTJM/p24Z520LusIEuOGW6SbN2yF4vVltrcQWLknXdQYGrDH0hx
xRkLYFlT7/o5AGN620pV3oniWYpfYAiN0R2tbx0VXe0Z5UJ3VKw88gYP09FxLvUg
efChl5zgkbnt3kDY0/dXzueFt/pY5FDyVoMgg4icIk/rKR8YEaytIEgn3l3i+RKa
NfjR0e6uSM8AardnVGs7GN4VkhSfdOVm9jKIZ8r73WZGHOuHFxYjmD5KhQWc7t1F
dwWkeIAto1baGKdK3Qn6RwPXu0q3FJAf7r/By8gdb/lcmVD66oYm4DRsVPWncmKw
i74mmlujg75tQUJ93IaKcAdv4viJnrhsUv2kT0WtxWyxu62yPAdh4lm8/JkFLt9v
+vWmGZ3UuJwRjoZlwm2eKIbBjb3D6GAvgnvIlf9T3TJ/BdGNVyfRySuAX2SGIB19
6Nq0V3Pf2gVLH8DA89oFc/oTS5I+oQJ+XJk043cfLM9pHAp63LLw33B4HtRFC+Gp
sKtIGJll4gdgjabhuOOjZgKbUy+uIUV4a4B5rtKh90RDtGHFB4Ds0xSnRfN1Pxcp
Ax09YuBGgMi75g7+SMtGGV1WNX/0NjjcICXBjrXUL0p51JXOW5d3TDMfKrexJB+k
JCqpw4qqSD275sQq3ooAazVACbB5c0FWUtX6nXFROvxaYOEsLF5xlIDntZ6qEhfl
z3xuhAY87vPYvgsmGzdLLtywRBBMGesEt9gjCM6s+lQ/MjqWkzEg1AeQ0MzS8Y2J
48zgNm1ZJVgG48ZfsswtsQmGjiW3v3e9T/VAZ/nwOQfCdtyRGoCvxJcyqWNR3ehD
WyUpfnEZ4vKDcXdc8HAkQ0NbhAwVE3n7X5A8MCn/xmyl/qN+ZK1i4HLCl/gbYvae
Qy9JJwBbozxk/Hs/L7j74/7Kgcuu39wY72wNiaNs1nAUvIvCm8dunanm+Kyy1lWW
AjP7nuOzxEiH3QeAUiWVF41SAEQ81fgAucMjv6H+i6FlRX9Q0ZEvdcfjrEY6KFJs
w0qZIRK0Z4eOCDtjtGFCbMSgiMYusut+T3iSAOCD5K1JiLxGvlPmdiaxcYOLRhiu
5LAJbI+36UbmcCBMoqAe2TH/NhCW4xBJRti4wATFrFEXdceUsGBL1EqKB9v5rWBC
SXJtU60KpLoT5iWHilT+fZEBRLV92/xzVxFwJvQsbhMgV/hMnNRSdnXIsBAndxF9
txhaY7KpUaLhU8ZVz4O8EXbL071yqMO4+QRP76n8MjLxICOWhRxgQJ6Nhu8mBimI
BfDHFlKwar7rWWJ4O+X5G02HejScCqNA8T/2uSIWbJtZcEh+1fDE2M0ZpSeRGFHz
DeVju7fYavl5S2ZiM9pO3FT3MnERyUa86AuSc2q8dl1SqyJ4S/UJ8584E3QZ1zgN
5m2mZyyFx3F6IvKF4+H6a2ZubM7/ogGejwoRutDPFmq8eJMKM3to1pXDya2NL58+
TaP/RGLHEPK8G7b3kEX1RDR9VrQB2wkytUrNB7rYqbBH/do/Lb4dgFNwvxMNuFvQ
Knb/+G7xcQIA7uBH+EFi4ygJwihpSVbtnlu2gkIrMV+QyNBNyjmJF9h2q1vkUlaO
NQm87ZLPd/J+uzuc7zUjFF9grkozsHj8auWGvpcmQKl/BGJFG/epqkPKWY9Q4G26
824ytNw3JBQTIXlL4hnqttChVjWq1nKONo3n6calmFMCdUh5nuohSnLfhaCB7G2Z
Er7ojhpjAz0bMFXbBicEPPA0JyDvhUqaCRzhW/3DObMXttiOXKGax30hbpvbguDn
OLY6qBO8QviUW7Tal95V3usKxAYLqkJ2E50M3tCALXsNj/uNe6OmO8b/KM3a7WfF
f/2Wi/c/sEo/OKR/BTya/U3PNQSGUoKd6y2bWFiVIKjPYPJrMf/TFxn89h6WDLQI
7tjSGN3g+aw8Iwf600HlmQdDaZ1iSP3+P5Z+IsL66qhUQqlTzi52AUJQnvYJjnYG
mf9WawdwEUwAXtPTnv3TUJgLYOX5hAUwMiKUaqVGk/+MhAeqD+wRi43YawOs9bW5
p7ylrf9qCAVU4mTniG4LyL7vovFAw89ffbkgPE0cgpqEcK759D/TKAp4XmSBLJQM
14Rds7qwn4VQRMjWY3pER5dQzcvYzOU27hdg9DT4KbOeI1ULNei6hXpRLwIJn1Co
OO8NGb+Hy02vsJZTIPDUFBurnAU6ctgpsbA+3O5J51zxTavieiHAvv7nx+KNRBRp
FT0EsTZyVU+afY/1UG8TXB5ESkUaJ+nqAelMfq2sT1cq5TY6QHVir3fE/Fg3xQ+u
RHjoscSv+9KALCp9vfqfl457m+8iffgyMaWJAaOCRaRQy9LM2rvf74cEbbssiZi7
VdFTMqU54Go103G/PHgpM6siKF66LYQY6r7+QHzQHfOZdtX1fNeifUSe4ClGga/r
f/VTBjapf8loAqkl798PiIQGe1FWxDhpPpvcav1UnS6pX5SlpqPRsapKUdtZH2Zs
36rQwjqh5p4oPEEC32LWgIUPgOQktzMZDZ2ocR+9RsHmZvklr486NrGJrXEwxd1j
HiNjGtb7iL3SetxJ0P8pKsy+bYwxkUw2IvNC5FzSteWYYLhjGGiMaIQFhj8LTfJh
oemdKgZZ87vS7PoLWikHCY1pqRPujhcQxA7kAp6AV30taL8InJwf19oKJ2ESUjue
kEyKk83XazFK+bMme4WWVPmsIfe9rfQyJsDb2jPcBae31VdYnFxZEcvEHDrAi9qZ
choG9E8tH5v/j/Gbe8vfkGBcwZNA3YI2gn5B93CqwlRJDJtpKPMrYtRiP+A0DSse
DZRBU041Eb4I7pq8uWtN0MKQrItsN8HRU6og4xTHrZM+5sFML0UjB/SoQ/Hbwamh
bCp4lCPUVhMLT8cjUkOWolW5F3dD6fr5IA3CJGyEgxQPOHXtvhpAB5b15TzUc6n0
ThGotEA4I61MFUFImJ6t+dXunr8NTt7ehfaOk4lTOHnpSXMvJcTR0M9oAuOByfLG
bhWltVSaaaaS7BeACFOrI+n3U8gJztQ/klK7kGL+l9DpMG3Bl22a/Hlofn0bwHiA
J74edqv+iZkluY05mjYND8zUIKBbDFMiGS2AWAVG1H1jxwUJYmhGr3U/pa03/aBg
zNEMpU+L8xFfOH7ojUsUGDa4yRkmrFDxWG7uDNCURykC+kc3Pkab9aeJ+fjKsYzx
6JnAK0j3qGCcW2ePFypJZBI9QyhiBPYuoyoDx99moTrcDaPmlncQDaJY/BYNFuOl
VONkQLIQ7R/QW2hntyWGGqAjkLfJS4zi3xq0+kXfjWinQBJGbGfsm3mRb29xarhW
TYN4qUT5UkGGoELfDuTVPIFpNZei+NXACR3TxO0OTzQDtgcEytK6AKOD6AEL7EEg
TQIX2nrHq9m5HCA0oA/3nb+yJgMXxscxlzzc/56vPKNoSdQhS4+p/jUXiTht3hiw
iJfRW7Zs/5eOQXR9kjKvYGdKc/wvxGy4mnQd7TC65s2/zWdC4mta83BiWi84709h
Qt1nj6rGGvH+/4wNM9GT5GvvttL+PsysmNcQupgJQtBDViK4HR7sBCXKzXYCltdv
sssmjSKJ1sB4o7gh59bmj36zV7UCt80S6AXZlcwP7lIBds7veJnnMoGgpHSTB759
fi7bogQcZDMnh+fzkKxLwNkFdqSBRNE1Qv8D1ZMy0n/+3ttUEkoNcjZbLd3HVt9U
q4SOuYPBEdeeW3mnbYj3oIuALE9ND17FPCiNL2CreMaSWYQq7pUL7WBn2APbZ1nq
KjiLxqCKuGCC43LErpU9b405tdScaDc/p6TSsgZqOi9MChA6nChI5GYHjwez/jbo
g5H6/mjt5Oz1EcgjIoPNu2l5FdqlamaSVIAo6kg9HQ90hRE3MHtsnrxYfR2adFZ0
opagh1bYo0RplTxg40NXrrhLhi0rYE88EfY5yAsj926yE38Ny0qviS0UNdO2tojk
5z6piNxIVDH3eoFxWIb9ifTh8LGRoUEq+6eJs4fL9dNajZmXNFJrNvPno/nLbsIP
ds0vhwI2Y3ZYPZrJgaUrMGLuA4N5CRmkV6Tz0zRZJqo1knHsYKFxi03ge87nEsBR
+W4yY7LuYdczWvgUHDRcD0RhvaGld/P113um8K0ajJdQ09KdIH5jvkRWR1DrM1Pr
QuyPKp2ApbwE0PUp6iL1Edq/v2L4F3kmyxhJi22wuTaTYe0aczUjyeeSdD4QueS3
2uSRNoXPqVmk1p5Cr7lWIqI8JTYCCjS1GxsLiRw2Bo9/h1084DxFOTf8+gKjm+2y
3+Qrdm1Q+rcAyDSgS3Vhu+WVs566fBLw0LIUVSeJuQPHFThWNkch3ImGc68aASzD
1aQ3XavsgB95OW7TYjKWg6pgpSZRcf83tnekpVK0ZWMDfGyiU7uWJ13pvO7EKZY8
P9q5SSuE8Rwrne1h4DWERFaeY3hdlcRXdhE8sMglcMKm3fzbF8wf1J9vIuZKcF9O
BSqvyKtAkKWfKEYUrKYsPR6uflU4hQCPn/MPJSYgBRdXA5fsxjj2l3s9bMql1N/0
TcpAdKOvwxT847daSW+WtRkuTV00TLR6UF4UEF9eQF/EVR3s+gnjCMaquf8AevHh
Qegi/N4WhGv+oQigZgp3OkAOp51mmrkw5km2qjiNvxFKeL16fh8seYgLGQZVVyY0
TB89DLA8ZJViGzKeTxnQUiGrh3BvLIYSWH4a7U4IHt+lc/EqvMKnakeZiRCbCNHl
go7Tx5BgiG3O/eLyroyKSTuAU2AAGSf+xDwMKfqCEA4a7lwTbqDEfSA4JrYWu9v1
UZAaQtgIomoFvK3gXZNH4mQS34skSXoBl6Vjqp7cIsAQnB1BuNkAAD7pw47lyXOi
JEEiXAu1RYo9z5hPShyMX5S2z3IRYsB4PEu9spywlP+gwqF5QefwU+j7hVXBrzAw
XOhuab/DgNbj/XRrTVXBeE5M9Arij9bB8s6mKkwRnHCKrxNFUwT8LpH0fsqYo7rB
INPXT4qmKM3xqhg7xzC2CdYNlhbyL/yy0UJvMmfbW8X5G+Ox/a7gst+tkBWINjCD
hbFvA5hBLFH+xrQGfV07AuZbzizIvL+jBs2v9frWGA0/gtvesnFFBj9cm1ebevkl
Mr1+EV7AMxnhWXgFr0E+04bL5TZ71zmFEcfw8FtwljT0afDB1PLm6g33U4MFnNKN
vWXk/uxoJX0RQyZBtPPYGY5dPYhM1iBfYmT+nQDyTD7s/mggVSG/CZj02mCE6Lb5
af3nDALVTyaoVx0rBQHJBGLzhKLaseqm0wNnopx7UOgOvnn5LbLzK/xPecwxKaro
yDFCfa3U42KYl3PhzCkMiAe6IcbwJugA6Ijo2W5t4t/pAN3jaFeKkphQqs5B1sQF
gwU+0olqiSq3KUFeNwlxz77kfqUEdDSvKV5KmTbzYyXrap1Vb2ztRgeo13//2rcM
95+qOoz95+wT/oK7Zgn2LQCC9y2JV+qR2L2DPP4eGPoPIIewvHu3QeSoBXFtNHCE
V4ffOHvoegWNAf4ES7vqAxIewidb6O2TxbvCrchqD6v9aUC+A0Gp1Sv9McrUDZ0U
JH5FC6nhkDTu0BYHTFGv/LTEJRavNuDLQPab9obeBuBFtMFZrki6uAMHficXlQiJ
1EkO+w12G3vME5UIBhNNAA8wN1FuPjY+fp60Y+jk1beAjxE6L9RZJNmwRO0rnEpY
75Fnggky4CKd8mUSSXiWhu2m0Do6GCGEr/fJa3S0WKhxLaySW4NAJ/MYDiJZPbyE
L0rv8jjKzgKeCliwx7jlqzF0NrFTi+j+4T2yfxHJcX4xbKwkTgHFoKiI5cyY4wu7
sYqdZkwQ2gGxyC+JZbryyY+FGhkFvyfeFlrs4FHMyw9g0nQ0lEDx/c0K1psFOPTP
jgG7JHQ8ib+vFcj6dKgJW+G9reDCgOW0XakqqFHZX+9RhBpzvb+jYsmzqKPzzboo
gGOFHSJZ8jPr2x/j/N276yHYnOdjRbenm8AdGWaoDXKdAwBEMAaDRuTDNvdfcZHi
6tGIp4xTp9REIcUWo3OfrlzN4FLSvm93dtWrDVafxOWI9ZaF4+SgyoswmxaVfj/J
tRnC3k00CjQXpWXHmLABcDWlWJ297SGEzRWR0/pEtBP4Ghk3NICSI8tw/v0zD06f
UnNvQlxzy1nN7umcDzkXNqYZuhCUu7QAtd3NczDQONoMH1z2/D+Am/8t8BChISDE
c6S9RgKTI3Y42WWUnuDvq0uC9SX63N6+cSKNAgrZtF9wzIXbliZx1LX47eNcuspG
8nxFaj1r87JRFmmDxNWlf6bO8XpI1viYkiykXOVf9Xx5A8A4x22EnzqS6VVy4sFA
fWaKlog57zOOaXn6PMbqCm+upJCJJLhatwPeDmts/e0ndQ2UgBIS/hoUxuiUuzvZ
Kw7WxaSYPuZVsEZWRxZlgVLYQlOth4l/rO7uKh/VIx4Muq2oEky2bh97ckCQPLL8
EDckZ9RtPoRceAM4GcyX5cJglsgO3/ItTRNg2q8JwFzppdoZMJSDxZMIbt15+V5E
b5SzG67bZ7dPj0TpDo4OHy6aurMgGdAYvKHg4DyyHHaCtk4DUzakhj6LeSI9xAYK
jSlrxNKeuBTqEAXXQ2zUmD+WrC5glTuBSi6efnDZcP4aBIGZYfrYsGomRriaPCfC
eddiZWmtwFkmFIsYkipZOXLYOXd1N5NbqKSBbJSPpWFjzAOxk9W55ztneiCYUMzg
AlJE3gaZ9cYoyqiK1jv8hmEXdvtFxhVH4HefHQg2NG6O36+Ad5rTseZeUT3iJ+eT
WqT6uG0mB5/STNDIi66BRPBkVMjpe186HldtCrYbU6qagHek1Pp/BUojk/PYI3EL
bTcI9K7RM4IqLlt8X550gNO199M0WV7YBERyf+C5+RiCpsyPIOBZDBLeTcJUxMAZ
BoFaRsz6G68seU4oDmxPoWXdatCyAGBODjTJBOxsJmN/GCar7m7DEwSi4mt3+1SP
YgP0Eu2iv7yJKTaSej70ZUZTtQZcoCWM8NagpvuLABPX9ZXyyIAhXJTEo9ooRRPj
FHaMGjZ9ak/jCtAgWgL6SXWyt/1AKFpHBTPztuP60PptveVs4TVeIakz7OslCw63
4Fl+GTwKKK5KnUtmhPcjfd2RgLikwUNn5gSyi2DujpFSQp9wIutc2RjvHFcY/v1/
sXa9OPqNP7Vr8GvkWDYlOi5n4VrkNeHbmF0NGbA5OwK6acXPwVPlunewIBy4cdjb
06u/p4lWe/aEjoDdK2vZsKrkst9TkfYwxTQuTbmoB29eL3Z+MObwkxhXI0ky1Qve
1H+ZsSyCNZ9OTrzyf01cyOuVOR0vaTemlBlYhLhWR7kXArMPyyZ2cZHrgvFXxQ3X
eecv4nALH2gYtP/iaEgHMEaGGLMZsyACwOgCZjKFxMTKq62zupKoVXjJ021kAESL
0Hey/vEveKtxgM+XoOJWPLN4Svd51e5bUpqaiYKY36ue31fJQn9iCEOZLpVtpjgG
TOgr7pk20SR5vLNY3YSLm9naZj5Bj2n43xNHZFI7DK74XdYTbMboER1/Ax+cvAOE
8P7wNqy+4C4ue5Me1Lw5HP89BcXBP/fBW/HGNLpUz/wf1+zK7tI44Zr8CyzBVnT/
IX0y+7fPzO8sCq0Yfuk4UfL2KBnxlIOVa4WMCDowq97HZZ9g909QgllkMCMaQ9Kh
fiwXpjK6mggCCGrDwxDp4rHb9VagzaBaFgKNZG0IdMQm8CHGCJW/jZKtpqhoj854
o4ob5ZfahOHWNcn32jwQAyIL1DaBt7Ooy05J7PGLXD7J827AkD2kKc4TiuN/Ogci
HzNJR78LRHsvVaRia/WXDh0gydpVytWZJx8+jmf6IJ7BRSVGith2TFp4eiVKyr1V
nIUJHDMl/MBx7yVc9VuuPViPpq60f8Sce5edqTAQLGKCFb0k69WNXqoUQa3SyxMM
7YSMNowA0hhSkevzI2An816cORiJYDFFOvkQaKOszv4nZ+TzO6aG8JjGd0/S/2Ls
mb4gzPu/gvQP6QaHHqJHGBVcSGS8hlVGZeBfVhjTaHJZF4snnlozXCEClTyFbNit
ew7kOi9UCHGtAy7lAp8HOwuDAvxWbhGQR67KSiXtFy4eL+iiYfihQhv+O1f6MmnH
ObdIXe13ah4wPDC8MJDOsZvXfwS5nsxjIBBuSsDnh9MQOaAhlPEDlj9QDoZ9gwGx
BOJOWTGJ0bEfLf8ar3qwqxVm7ZknzlW40j9pwuRpAkwH91foazvJuNFSsWbPGLfX
khNTk/byhd1zhZilFick4quapQFtiLMOUzdxhDoLmpvSC/e5wmTiTyE8k0fYBcxu
n5SDX5ITibRZvM2baGkSBihM9LCwRMPxnjZRXFHwKmchgdfYLNSXPF/zjxp+SX0n
dSJI1xdjiwHgQ4Aih0xnh24Y6lOrzC4gB3r+T5sFwcMSHWFBXdEwEc9JZ9radhC1
eZkKygEvxrup299Iu0fvPKem0ZfLRZgIatNBTZmXrrWX/fIicn4rnGclH7XmLOfN
bB0xQZtHCpL3jIgs7OBcjtEDinaT/yxOZ7goNksoCNcLHw92qS8AK1zz8JdLZG/p
AbXL+bgwDs3AE9lSr1ZVp3pN4TqOWRKvrev+c7mLbpGNPxpZ3bD710T47m0mkQBQ
/CIX1BLQ+nr9kLvBcwUxdBG7jmYORmDC6FUav5AwLu21JYW8mZAijY7Of2kxGWH3
Z48264zbTWIVJWHXIPEZNEW8uFSc/m6HzpTSeUIo50vLDXGHjiEcTBXMO9vxz3w1
ph8OEi8onxVwK5bW5We+EkYq1ZyLYI1G8gIeTRzq7MH6IOs/ePQ+E0xTacpPA0dI
ZZxRkO/C5zHI1yr/j3agknzzhL3hBKwg+stSkFCKuBx8Ti8DXv6OoWM/baqkMftU
liW6eQvtgT+Osmu29XejXS6VdMmcMt3E+AkznJACvGz6SlTPFQ/iCIVzWr+GaZ9n
ox78Vxd6Qm+jTbP6oZjE8N29xBHcIm/dgIumZtl2LmmII2EnIVMa6mo1QWRyhbUk
64w4V39OwPKbunOx36SoLNBgAvFzl9sxNXT0LeM6TYZenGinscxNwrrpz0WfymSc
ucZBuWZDywqNY23cdGkNRioShcBvAVjJsu2KFrGFZAYUjyvT0DW7ic5DxXfzv+Jr
lJ7WQAcY5d6VTQeGi2qKtrsQEhqms4kQ9HFcBiPxLvEFSczYvPoDM732+XiC8pzL
qwrO7He5QC2PKJAxH8uLben3VghG49erzguDzvHVdNG89tiLifTDPoKk28gbNRkM
JwgyOTPBZ/XHWX8a0YzXSUAJmjKyrDvLwuiA4qiFqrofmWq5CSoYtlNkBsJ1FZo1
cB0m+FWPXXLP4l0sDYGfpcTu+4YMffHBg35n6jfoVdXltt20dP6eeMehBieURCbB
lXjrGoL8nWeR+B0mB5fnZj9zQWoVkRzor7y0OjyceigT68WGXPi9bmauOdtN+Fb2
bds1v2SLEEm61hlEttlNy/IcLKQ5A2WSemmIsFiQBGKJgOXkaVkmz9IaD9VoesGO
0amEmF6itUDxmoGpqGO/CgpVyvyLtVQphoA6WLP+XE8ADIjeIfX/H14yRe+hEiuN
35NQm4MH0WK0B3cIv+iAlW4yPW0hhwUKxF0jBg/1zT/Cv7T6TuihX8I8x64Jqg+5
3v+0tmEWvQLWbdQQLrCdZGADOz+J+ZvNmwOa8RiO66e4MAOtQtvP6O+HSKeLz8j6
PETRfDWbw1GZbi6mTNlbGb1cXMN9LFqoP5GU9yyGOfGeCkQ0bT/9O+UHpDYB3cJY
x6TVAarXTFpxZK+6ft8zn7Awe5uOEtpxrhCXEDBzP9XmgM6i/6QqqgBiCpUAxD1F
lQYCIrIYQ+lptQpwEbd2wgS1k/ZsTXO3CFDlDFvmmgGfO6xrE7nelYu9J/5PGIv9
nDGNM/B3qlusVcMi6GUDPY9R/xmIYeaW+EUtQfh3bYDm7GzzKSU34R4eAdAlaxps
6ykFLkNJBtvAgJL8ixIU0OVJJhhYCm3I9+YfgdmzkeT3u4j8b27XvZHpdA5rryfU
lNU17AumQKsYGAQzXx54Wq3tcKutHZy85wsaiJOzKK1jeSkDAfxwVH4KHNWyQHf4
5EnBxaoY4g3Def7Er2O1yNbzjjqZNw5quoDctZcgRPbU2hkf/BepkawVW4CR3s1C
dQL+YJeFqIQwWJI3TvyQ65NG6hYHSYqoh97RappHznOyIS9FEctg+a0XINuRCdKb
RSSlXkH3JIDNepavIfixtP5JfWvO3Aqe7cmUj2gCSYkjsJG2kRlytoi46e4Gyax+
KmmZ+b2RailvWD99TFpu+2tVqhMlkyzCvbb0iCQxezuw5SM3bgqVLczqxtoNuHln
fUzS2TtOKsm3J6RNR+SlwmUs6dXxDWjLmVo42np5jNmVFkxYGNclkzVXZ9oQ5pw4
w0ZoQoHH2f1uJECuUvVzqvxAWlFaDcBHe5S/KzltnNGasG35enrJwqWAmhvrny5A
gcLB9St/0OJ8NL9qHxTNC1shVPPi0g75jh9iZB+4UUtEbTHtjlFW2PdDeDhflEl8
avNF6pqBcG1rMhCb4HFnCdTrts4wL3S2XZGT7wUawFDsXboJA+dKphku8iouWeMV
R12KZD5KseYhFPENE4iD6L9QoxA+dTMBVxxuA3N9FYleSwGv2RfCXMbNJ+cOasEt
TPTwJpltbB7R3DqC8kPP16eNxp22qBD935G+/SnRRUSy+GRCGphJJ5JRydjOqh5M
2I1PnBnQ4ZGo2sE+0Il/LJwF4iUA4irXBkg3FwEtL7YL4S73IgpnlRlof52Zjux0
Mu3nLbrI/XADQfgeXDvctp8PoN6XQcOagFAfcj9DG7J66vCodIRuRMeZBCicn1R2
I8W+8hnT4aOuoR2PHrZqpLMB0FhxSFG4ls8jl3jOBcOdXXSWhWdVjP6KacHwWL/n
RtGbTiUbFXzwOP+p7eI3F2AgmPKFdfC/psoU79i9duJS2+Q8TYPtW89xOIWJpPRO
+K5yBOtcm1eUo4X6YpiITpz6ApbYxNR06nBmOjyzjpWimXt5Wi7OTpVu97UE5zJG
yu5Iz6zhfD3cUnTlIDXZXAHzhZjuy1wexpMEJINnKtM+OKziU9PbC77ApAMDZkj7
wIPeqLWH5jS2Qku+WfqN383hjfhnJissi3K7bV8cd2AzjNWYZlDtG5DnUBFqeUuQ
Dv9DcCXIGnbmYUI2lBQAVUu+9kW0odFvUs8wssBsfe+lRzrvx2R6GStd8KEYtFIV
LcUJCtMbkH78ZHVfPJapDM+Lhjyll3uiPywjbvk5xWoXmMehevruSLD43Q6TmWuV
1r7dyMFkr0ataT+wVh9iKK+fW8p5YUzuHbVri68fgZUMO7lAYwCTAfBiDrYs+Aac
rYgw9m7GczVIBe9fWFKPwN2ebgQ6ER87jI/OddrkC+OrsWvTevxnnlMZ7XA4ZcUa
JQH/w0ENB9bkPPhKo8dGkSvZdCJQXOAZBrQgzWJebr08Q3HrZa7Isj/IwXWdeJ0G
9eIyKWIhgstPO9BYmGkGfx6H5ZpvQqBJwG0filRqBF3goZz29S9M/YXVgEnbRj0S
a9rwpZsaZQfKwIf/9yQith8aZZ1dE5D5Q0wu0Wi5IABjl4k6VzcguObUCr8+nvzE
iM0NX9gEz/DPN2J1ece94I/T5d7OoLkjpYEWd/4+SzT/znlHgGhSYIEHVexnRgba
CY/ZICb3rXYSWw/tXyhbtoWYe1X6wqbcccetzYML5iMI7blP2yuqd36t2xN+0vVm
jgz/TOg4egarR+tvdI0dkpY8V1e31mkOOs9lj9QlPtRnvkiawFreJL3Ost5aK7f5
5O0quBrkv46k2vLr0YtEJrGhOZ2iU37eMGq8p34SYu2iCqfv9IkgBHZNYgwI/Rtt
cCliNuBFvXwO+89bcqd95hrM6eoIi+Ho0kgr97Zkx6DV7W2Btj6pUswfPsa+e9l8
6E9KsmD+iQOm+vkZ2TfhWES6w+Icr3pF3vOWZVoECIkr+si5pEQWQuaxQwNLRTxy
3ktSP/yfSP+Gb8P+w1QT7z2p0b2hIq5/gZIw/HNlUvSnEiOM+4Lf0DpQb54mxy1J
4ngZDFZA++bQajqCepeAaT3g9RZNp/6bupAJVaE+C1ivo5HVu1hM20ys04ITiHaA
CBgUSAuTJ+I1OFXZ+XnfbL1kZq6qVH3TKhuJnM0hFQa8nrRHbp4B+p//UXxBEeDU
XkHTW9R+dq8ZeSSSm1iqavlC7NPA+8wSYB+dP8+ExZChqUZYmpOVQVxw/YEqCpcp
EEVWcqd8IoZmo3aOJItV+yjMknWSVb3UIQjLxcLZ2Nm3prFo1HRlzMgo3PT3QEcC
wFXZshQRq+dSYuOCzkg8jtLcWXZpBLacEKhjKXU52wWJ79QfUrqGrOkl3WXBaXIz
XPTG4xRffN2ZhhYJkv97Sailb4kQTEY888ecf+nrr/KMbu3AdmhibmrNkv6MbswT
SNuhsZif/Shkm96fXPTU04BBMdl06SzFERQx4B3NivzZrH5sY2PufKqrCR+UGrcP
61pZhcwkew+ivpI0GaXyJ+n0LhfKiTBRRARCMIaQNa3q/T3urVo6uT6ROUt2fVbe
PCZVGEFoCtW05mWvBxuVF0uenL/cgx/McDfzFBYe+gr7dmbWgYmtlxxse+HgF3Jp
R/pXh7M078mLEvbroNrqA5vcCnMoZfLZ7ze/QAqFR3FqG4TbMZwDdpdEVWY0bRV0
dgzh/MNAXIh8qEe4Q9UeSwqq9wkm2iZC7LxbqmcRSxKNKc+/nWAc/q2m9lYcrEEy
3Ppcim6p+ink00IXp7RBbEW1X6vXfjzNc856HwLkZ+IUc+138jWNQynpYH7sG4s2
Vx1NL1WxN+jchp8uYCT/cCYINVRFXVPfqhDMMYztXqiODjOjdryyRkeeY/qLMEPw
DO0OAE2z+8WiBAzbrVJ71IoSw0A8WCxkyhuoOqRgqVntbbULg5FR/0DjIRPXvLne
RxrWGfy/2ZmCJ+V859foU/bf3axhJSjI0yr9Mu4hImzSJt35RGORJcAboq8vdCnS
QNfOuCsattWqEjvhIdlJIdk3Y1wM/hBz1jQvkZWrwvzkT5HrdhkqPSlxKKhntlGs
TFRFh4vIgkUcn6QAu44wFUbE8Oe+0tvZ0WvXpi/C/eJ4TJG30ppZpBw+NiI/AdLi
Lilvar/T41663wYwcY0D1TfdlBfIpG+PA07IvLIYw4iYkmxUz36zk62iKHi9I5C6
hURNO2qAOIYuLKtf/jxogx9A6lru/kr70NQfc6MmzfT9bG4gfwMqNRgciG1XX8Tp
Sf4dgifwX6cPvW5RvPjPj8qdDOLAczRUTi56tMEN3pvbvo+pBsu3Q1pAlpar836p
VR+YafXdQWGiZX9a7WJxYFHiuRaP1XAFLaAjRXNW/rTdQPgFeEXMwWhIYud8U4JM
BW9uBX6hWa/jza0Vz9iIq1qBQm+AI5Y3RGEWChzaxoLBtEfp3H+WnrziQ0SicM/H
kCJJXJ7R0pWUAF/RzrC5GHbA0jaLsDsemk/OtPhqsxnJX4Wbka7fCfs67Ye2kDwH
kASjkVjOjkHkXNW8SpCdsVnANn07b+kYTjRvjDGguIXVEV0/NHlEbwSuelniYtcw
72diOMccEgay84I4w6yw7jJhHQjujsA9A9iqjh8dCx9VGENjPc99KwZ6y9RnsFg8
bFP+sXkyMcCDIeB95pRcA2oiLo503UvjmJ0Ck3+rC5QLqgne74b3A7njBYXnY7k7
Y7K50C8scugRuVL1quv8ac3tyu9dwAA7g5YYA37JhT2ipUOWFVc1+tjU0SdcK4dA
Yx36cIK1hPRMGrBuk76V6IKhmpcu1Zza6WI847j0hgYGbwAh+CVUirkYkEZKadOD
H4SMmapLZN/hHL8BEKsagkZ33KXhIJgHvy+kvgb/A/oR+9Mp2X2rmF2mRVw0g7f5
VM71abdmj6ikwWdw7bnR/JAAD2mH/TUz4qvrC9VwR3wH1VDMtX4glrF6s8cFGH7j
DBuoK2l6fm4PC9CpL6YqpJSvGjc7PV/OUcdnynsxDks7dfzvNygk5opJiZDTk99Y
jIxw3ab067KZvp9sXk7ANEk4ZRheMn/2lwBb/Pb/TNIDS9jDiC+eveyVe4o7Qsac
ZIW2f8UsIFUbbYuzacuP/DwW1HZBiM1Y3WmSJ5FrjkoijY7uMqMIqyNNigkTcssF
IlD1bQ22FgIztYG+wX9znJ7SzeXsk0gvlU/bYTXdeQLx9nQyalF9XKSjamxTqwYs
IVaOfPfEKXRSXSXeKTGgbBTDz/goG1NBP76dkYR5NfFVKdgU85j2HVi1qGK5cWen
6yI/yBbF+RQUjEMegqZANJEMSG+mm4BJrrUnCTBxlXb8BprCDQRVI9HlX0Wxus7Y
YndXyrdpFqmmNhl/GDfXbR8XW8pMAwEOTyJyG4uRXWVmO1IYWkyeM6xeOtbfFqZB
C3Z8fK8ZClg4sgQVf6u0IqSUoIc4Zw28XdFA3zrxq2skLEry5Y1og/aIdG3+N2lV
5DkUsLGS9dfKBdAkfvzsaAPohf8njJJMb2jzwJ/lUmZspxB3fJOlIuC4KyiAkBSF
s6Mvu5Tt8pCdmQaV2A+2GH6OAXkEPluxgtvNSm8hoLT7Iiu/1i1vxGZEOrF9C8jX
62L3/G5abQRzGKrdpdeJLOJwLu3gU5pS/BF/Uz7a9g2Xb/givJq/RG6DPUVYS4M0
eeZsZRO/7IbMwZEwNwmGd/rtPSD1EBGhJ0RXBeg2Ex6vv6cBsu9MhrK9P97gLpMT
gNnb8NtqTDMmkLq99g+SOMam+LZS1B/1ewD6g246imTVwrtZj2VzJhcfyD/aOAV0
xGgCgjgWjC8VVIMhzyJwdWxG1prsOpda681MANjWQFVQFg55i/DUp52Wo/YLzm5X
VSe2mtlLEnIPXntNT9JqPEQAOe9A1znPXa2uAkrc/+PDCVxgO7+YEZQmfrXaG4Jx
fvcHaU+V8Ml5va+1w2Tn3vimE6v/4d1bekAg2k/zJXZt+3N+ziBm+SSa6frArfbS
3QTqsdmAMLeVP79PB8PYDs3/ESMSK5SDfuhp2zu7gJh0yMy5lBbNLuNllJ5gLbgi
xhy1rocVM2wplTKMt/bqNyiw+HbHRqjK61f8b2qBQfzcdooMzDuXsgjJt3dNgvT+
RM7cDpr5aWXdaxgcl0k8rOnRy+2hV5AzHkHeGyM0v6utpgpYRyx2YXO2r4GdYDcy
+qkfvAp4pZqfTA23mku9PUhXoHlSzrCtAjTiMy3eAUp+2gZPFgtyTe8o/F42FeaT
pRYxSUNA1BHc4ypJ9gYICuYwm9wSrsTKKX+fgxEEcwgT+YlC1g3+mziV+czBeN7N
rXvchE2po+Wyid+tIZFSwqMeHHqWByjtVQlSFkMcqXadIkVsVo4llcaG2iSi0Phb
05YW9cwKS6vvH0Ch/hT7lkIIBIP0FsXmRctDXpQkc1YFE+9ZoObnMcb1CtS5IIg6
bV9mpStIS/l3W50O9cmHcOEuCS2sJj7Naj0tqJjcahZ1gTxidH8cR3W/FQ8sQ5Rv
3NaJmWjt8cJ8r/KUWtZVLapoYreopJEV/cHuN5xcAZWj0SOKv6MCP6477DgfV6gA
P27bEIT+nmsy/n9OvtptqP/IuB313/OEstEeZRCYUeXd7N/Ybg7G1shBEYjd1hvp
rZj5goEBxfWgwS/i1HCtaTF8bCYbqT+kegBuZjhVOVpHQZsov5ljEHdJz9aNTaOX
DKCtKPsz1p9SiX5pcepucQFnnFia5S2Ot4qFHHhz2ul6HPX1lwKXgxRre7mcB7/y
N9IT2edY4wsJd3TtGZ/gpTY1V8V8g5R9RJDiuqkat3hvhaRk8dvz9PxjYxBwq4+P
vCHPMZ4NNn77YMsw7qQ4glbm41P29+O1cc2yqnRXzveW064QYi1xqD8dDum1Fmdi
uiMXKHdXQUCWCBRbH6nBT+EPoWV7VU3z1ooQOYfFmZsS5QSNw81Lkcf0QWAvj2rY
heesPb5CKgitcH9gdOc3WcmmuBD0zDYYR7Mr5aS5WnUhCobUTYLA4Oswx5VBqaED
LC9FaJLzkaCItz7FK9PTDC2ca69wMLthzGjyMyFKxYPXLWlxfPWWByShZOhqPWw1
3SN9anc+7EB+dVMkdwtWxY5i8SMr+wNhtk2MqrIG2G/dLfh+3uA31jXv2jOQwhMT
sx2PsSRx6ls+1BT/XHkNttID+yJdjljKFaNe1oWh8mxHCM/6VjP7Yl27xeVW5TW8
qJfQ9dMZjMugXAqr5uvJhBMzHOlD1ABhaIVwCcQs4sjEwN1mES2M88OI1IxV5Iow
821UtYeAlpOl2k+3XsNUn2pd63jmNPkgVgTLRUXGmOxM1FoXjgO8R8xB75I/CFX6
pAthsuRDkrhmFRv5Ref9cKo7MxnDbXiQQNA8CVtGLzYd2zeIRFvQTUod4BUZrzgs
mPvzK9aIb6jPtGe3cKpsZxQhGmSmTGrzEPXSgj34MjFV+WZ6wFZMtGrSwIJwfkoU
8sNO7xhzQt7MhnwpX2GXpNvu0Rv+XRmiiAQLZp4auoK6JPcTNomCbtjiUrofuu3R
hed66h+f/OT11/rSLLVONyxXrNNa8UWfRwdzw3nUSmQuhyETO4K9p/auTmSJemWr
oLTXFUk9utm4bXXOuKWxVN/wKxLDFUB+DqU58Iind5vK2sopN5vJRCuJBDCwkBWW
SNUZGNxRzd9LuzWqw9ta1Hnw8w3QgBBuZYSI6ECKwhiu0VDQhBoesIsHFEBhnTcR
acixBD8dSplPvP4dlRJS9j6IKgtpnO2OzSTQp4CBzkzt4kWlXzlfVZUmErITfRpO
e0pa+ADalx72VVnVigemXEC1P2fFPDiKsj+759mrFTP0C0enCd6YqnetxDQtmND9
sWEksamLs6paN38pFETfpfTNNMuwp3bxNhOG1XIYNFb5o1pvg7/MlaO4MfVtiFiA
9Kbvjr88BJRovRarjnPIItHQu1OmHcuaPma9J5KVs890LwVv1j8SSXqFoLNxwl3F
nt0ZafQv2G11GybHURMGKcNVdl/eOWNAiBbt8WTGjy2BAy0ooDTfNBMoFuvi3iJ0
o0KfHak4TGJ+jBAOlA8VpM1vjFVseuCwImFzpWiWZa/59o0wgfE+Cxh2zMeuQkUu
WLhaF+y9rD7TDSXoN60DrYgBjwh2W5YMsGz2gk0APpMz/5j9hNecZCLLnFA2TYb7
Q11PcaRwhnMthDaVCUxbMI4maAFPQJzo+yi1BXKOXp+3+CBVC6dzPo3zyhD/MgHU
0Q96fddo+wAiaZkJgfffZkCgmtwvcdHjRyR7wm+jOCTtFfaA9tzmyHd0ucCo31K/
E/qAwm4yEXCJYjGloydZeMudNtbac/J3JsCZ3i7gjS3TUVRJoQjlapRR12G5TUig
puNYtJB0Tp/lrQ55YwwwnBLU6ARTwFBlBlFY2wvOYKD2Rd8mYGqeUIJEqxR7HvUf
Wjn3KIxSFmH+XRaxPYthN2a0G66MQIHXCSJsea6m+Ed+BrsruNDSzcSw2RNcLDdv
5SBJiavRp8amkllwhkIm56mPRz89nqDi2CPAlZBQ9IcsrLt9gYhmvQ5pc7UJTKFI
cxv7a6fcieRrcAtppRTWqceVDVmsjulGs6zt7b29xLENkPrE7T4oOFmJpAXwqX3u
P8tAbo7Qyn0H4I52yt0+WmrbES4JiA2lUY0fN9Z0LNEhnqT07Bg0fRHIw043v6Yr
LNCnIGDr9WxnkMOZA73PWctsNTNjcNu9skNP1tlbe+j3iIcXFAgxQR7nI+m6GK0k
TSC8UrmH24UxXBE3xbldvKaNXzdBCe/ncttRHrJEc1r1S29pIO6zjOE1uNMugrFy
YL9rHpUDxw7h+TD3MRgCX+q8HohMQES8Ofhm+pIP0/2HfBM1ri2Hzuow8Qji/Hr6
/AbSf/065A3RmJVWGy9WZ52en/+zJ9fnMyRlC9k5bZX6mVYqAeC/6ocykhSD3Tfz
kG30vMYK7LzLpPonjQ5zYAF1ND5d8lRUD2/w5U/yDBJ8ijX1kf1qRlSQx+jGmrXx
5DJC1Dh0MPAhZNQsm+ghVUCc0pjPToRnC5ZSmaNm0vOGaLVQjlkdGHvJji128tfd
R56jssgwZpgvTzgWo1Cevg4aSV0Cy9RpA2uzdbHFyde1kB7bzl2YpfrGK+v3WObV
tewIOUEfshjcjDjBAdo1RWr2+duUiboZtFpGXoqkqvyQIaxfPnZZUkYHyl6GpFHN
AOEYeCbf6q3Rh8thg2IOy4dWoM2ONlAsA+s58dq5/1TNS/egepZfNXEyRg193W9S
d8JpaqAA6XzdUuTiaBIMnF/2VCXaj+MsEqLWwKUKkLsR5RyNNzTvAX3EHL1bKOWR
JksE70HKExWHgrKGYr+eq18mq7kqHIyKamtS8+Nt7kXivgK6OeuGMBG34IUgVewg
LY6w0WtyUdcnHnGG2X0eZc89FUOJUZWO2/LKvL7K+XithLA7Tj+ALMcykj2ukek0
ik6lfJuw0k1/UOnfOTe5jQ2FIHEizUHGsjMAHvwvnY58I8XqLJwxGJwdLifWTOoJ
CcAmXmtmzZP7jBjIzdOtBfAuCKnZlEuWACL7CSjyQ1Ip9jviUIQZSjD3AjRWEF4z
Yt6lnZA8X1cQud+a5TIHKpMVBTseOLYPE5Yf3JpEk1EOwj1W/Q2OvtZe83ZYZJbS
lutu2U+JfCDMvPMU07bcMWmE+0ioeEPwsCtH0f8X/+Gyll8F6Y0Ack7gZB8eHpf4
ZBjs86qOAjRbk5S314WpGgULlTtovPDOqKO4gHs4BnbKL0YDn5MiAn0BA+JMsDFE
i2F5PSdsUUAx22Sb7g1Kb0rPEibAOGyp/8dHQ5gOFT4lKjBY9UZ8cGRds+qiank9
Ou32YX2RXh1v2wyW1W/7dbHeKfHthx7+V8BmIYt+RKI/fm6A+t54gSgh8CrBceEK
Yr23IyZBauJo9MCfAjP8e42KstfDR+sCEjxWNXbi0s4e4kZK1DY2bjBHMZ/dAbMq
bwLXd/ty/Ywa7bmSfimIMy+WDkE35sxtEN0maWclJeLXBvaCg91lrvGLiQYoncAZ
DoeyyxbPDtFy+1JjhfkU/Vp1k/FRc3wF8cZmioWabK98eDnftz0YbgYWfVps2yNa
DwVS9WL2rHtSc0TIfyjehP7SULU8dDRFPsxW2YkDCn8SRZBCYvhZEhlx7pBMUhwZ
61WeuWSSM5fs6TC/+U2njKPO8vYy3VTLgxLSBPE6agAzPytxSJbS4aDaQD/hNTGv
DpKZVBy+kN3C5s0noYCcXqGct49ZL4oPoB5yhNLu2+xiIHcj56GwGerBVYgHOD2K
Q5ejkzsY/nCRJYxqJnrnPwT//fxDbC1P5Luf33kV5T8EVmx0C17JCNsFlzsyL0P8
ox+va4IcA4yepAJpCFTsKM2xh8sciQMmu8DBtwcTx2pABL4QlJKb/Kzvsh/lPOCQ
HIUTNEE58zmKgDUmCZLn28FY6TmNs9/jPwHkuWyW3JRll8RCJutZyQbS/hYt5ylb
aAcrre/80lRLSEfCfxVIalJzPoeYe+/UEi6uVHlXmwrJ3WxpissKJ64DRmyTmmX3
sYC1K+JFPB/kf6xy1bbgEgn9HnGk5sI2iA74XK1B1uAOfwdwIv9pMREUQCB+hmLK
OsYdyndM7OXA5I/kDy7p1YGL1hzgiDBY25IUPc49M2kxCzSKz8sRIUQiiN/QP9zE
GhMsqXLE3o8hUu+fKEyZUT+vdLTACKvLxJzGVsM42RQQDpYfnftBtcUpnGFwKroM
ApCIotxxdrn1ZVvYPI6uaElQUGMBW5ISDmm/4xy1/H8JsqtJ3CjEhc1ZaMC5gNX8
qjSyWFuITtaq/KWlc8nL86i28T186FQtdiK01uZ6nocktcG1tgF81j5iFc3cI0Tn
oaKoUCtnOgK5blSf22uY2OUD1ITNgZgZ216EHaP+/hDGku70cx0ZolyF7gZfkrnd
/A2EQtdHWeovQAt/4AciwAZvnLT4qszABxdX87m6rFqf9UBYs0eOiCX38iPV7H+C
1kqeiq+yRXIZh3X8wOWXNqQbFywiZ+DepOhFTyeM5zA/SmqqXZMjGMERjblxMNLE
OmO3WRJPQd/KAzlYaMfg1okW3nb1GmChoag9imhe/rK5YI/9ezaudIbQ4kAh8S6c
JHnYFa1xYpRtXgAqwPeBN5O6apOMUlYSlofPx6Nj5RTQP5jDcohOcoMeJ/uQS2vM
CMFhvKvm3XdCGvmSKHzrxcpAIch4oCmk5202wdDlh0J637BdJ9G2KVYwgzpv0vIb
3i8lTgvV/Gl3IP1Xd98ak+lMYTA3SrhSqrjU0U247wsocOeqKU6BUt0Bx9Ol6Ge+
0HRNKFJDH0TUREvHAPKDgtRvvCLJWMJombmIX5XmcAQTWbA6OAylLIHmKSQU1yxA
8H9P0S/9EqdUz1QOsZzvzRWv+g+X9e039v8XTDoaqzoJ2Zdzi6wiG2HqMbIthDvM
9VF5ovyJHHYTYwBrgrj9+An6/FB3LGSDTamBFCnjjS9pto/ZUq1Ay4UC/M7T0Nji
Y3YCU3rDtyo3AFd4gQ8j1fsNVexE0wxduk355XHIASZ5hRiGs09yZMal/HIC8WnC
NStwZ9fa6BDFucbHRWLCtgwsS1TyuGkpW9sJY5SImD+C91DDcv3Zibs7CxjSaaNq
CASO4Ur66yHk7J/ewfPWUueDmrAiXw73a++FLJuEgmB5c3HMwOOo5L6jFgqUgd2G
Bg/6IGlliyK5Nv+BMKoTkjK6v7pFIdmspfSh+GuT7d/Mf4CkKymdYmBOpZh9Z6KS
tdLhgUdfigSBYppXSuuIkRG1gKiEIWuhI8xAb8IaMtfRtIWVbS++YpbvIRK+pDmY
ZF1Suh5sbkINNOnRwtmkRUp/V1gYt3U0MshOthOkNL1W9ExIems/flmKRtfSnquS
r+lGYWegEz/W1BtFkl5SnhHfIJcaf6ph9hgt06ccxf4bQOeSKStwAQgfEOehTn4o
KCUxYHI7anauqq7azDQFCwYJ1hMf5/h9mM8NxGm52wnEPYEevMKCDAlUfuIp3SQu
lH+GhekowaQhJUeeFBFzM/PrtIeNOPldiBs8ZOR0zzfTwKVPi9ZKOO+4DKTJf1gE
K2JqtzFjTLb2T+rlRDMGh4kELfKpvf1zO2YHAHD9p3F4wqlEKjt+nhVCAGX1vVQt
F0B7ap3fdnXuFOZhno+4alFepzB6WMvlstLMR4YvtlbbaeP61gO1GcvZmdN5nlZV
wkMmaZyZ4HaFP3cs88kItLJhzO52lHdj7Uje0WELLkxD3Yx2xsE039x3UWw1XBLj
rfo484FIJvUhgwRDrRilaFDH7JEBmPPHQjY9q7f92pbR3w+tPnRzc4xnxRPRA7GS
JISfyExuQ9+u8CFvGOPouFPrhte5OFIUHR5i45Sa1T3hKBV1VmE7Tj3sp4nl3a+a
aKyn4sb7TUsxMdaaw4XhB0h1i8nxxLu2yavR8GgX7RpGK470PP3d9bL0MT++ivqX
dUY/4Gp+nDElY3uNkPYbeYgFMkOAYHjUTEgEjHg9pzyW/QDUVSdnXB83SYHObCE9
SWCxdys2c2pqa/SHVLiUPecWALHFj9uPVS/yld42a0bUjjoR5CL8rnVNXjoMzP8I
8U8lDF8XX77paCrGHuwb7xWI21c6cicsDkTPsBLw1ikWq7sfF2okWrCIZ7on+KZn
Bjq/K7NUmbYOkG5HB8GRSj0X3lzNLtump66+MHweQO2eSxNMS88cnY4q5htE8nY4
w5xSz4wLfPu+wo5BIMQofcyZw+8OzmLYRTlvfsu4L57oGhJoehBDkl+5t2EVY3ua
INez0gTe4GYy3YtFNQpxS+49DiO1H+z+b9Fgq+jSDa0iqwtiMCvv2eteEhS2R/cl
gISeqTVSiSguoPwn4yymAiw0u7m00srzHGLjFd4xTd0yu8PuROy80IcX/DxIQT1d
pM0jTLBJvsbnJkw4PMan6j/pP2Ykm+zkS0eSBD1zqfSs/Q7ErsqUgE9Wii5PWART
LmBjomQU0iu5nQxJnOuoG+Dzkn98t9ZX98HPDXGr7V9Gkc3GDV5snaTb9OKQyZNr
SlTJHyNcL5OVG1qI8d4AHsQZSZQWGOO/Bgb9e01BoSTEZNn3jTXjpyM22cFVMDZE
qnh1BAOuVwLvfzfza8Pyamb6e9ZeZnE+LFbhngU8ppIDQotTf9Z1mDU29jiL+fSm
tSvVlB7SHUyQShOsfHGQXLO6faDmfr5Gntjpb8/IiMNN6HDuZdlLvnNjm7HHfquF
lEEczE5va13zL8Q2rXwCEYD6A9+LSo0/3Geo5Rbb6a0YaS17TnkmIf57paUSHBgk
zCfSlBixXCq8Mqsb0EyP88PJnaKY6I8FJO+R9bjHcDjXqKyR+qkUThJpQkrTVimP
OUdHqyOhJsljKu+lpGJTVj1UPKT9MqFX01or2J0eaHN1QI/7gGAqbil6+thJVFuR
7f8ieBdaaUV1nnHlQQXU6WViYQMc4JzNu661ZQcJNyAONdi4fm/mjbyCNvS0If/d
+ZtTjJeop7MemaKjgCcGrqYEiHaSch8SNKXo5UBlgv/hNu3Rz/hJNsT36YvdsfRy
92TbIMcIxO6ccawaw2eHLF5/kD0dJD6lAMo8Prhg07Hp9tX+D5m34jdTACk9G6Am
2tpFaxFPijVy5rnyBI3FZLTBUcot4cTfxny7Ilrg1Wv17JasJLedl9YovTE8JkFg
DWXyvu9AGbHDldWT8wJqmNBCFPjVN79qmC2ym/+9NwJ0EwO4g4f0TsnFHJpBBHqC
Ku/nb9c1CsEoEjw0nL+FEPGPV72bfBrSFlQgPx2trvWqu2NdO80d6vsbjSc93lUL
o26lKQvitrMsxMSNrtGQCk5tYsIOWe/eh2cMaPSsqa7g2qEsrnOttr7A73lBldNh
9JO/C6+B3+veV6KFxfd5H6OTk6eCFAKxKZG19+MtAcS4ySx2dLRVNpsFn4keY6fs
f95vnvY8kb1V3mLyBdHe19goIFVOA59lf3It4xjNGKyvLobVERZnOFgdSc8fusOW
a7JI0vhORIDGwOCG1DCJw0SfrgZao3xOROf1HSlhyYCQT0MqvBTbXHGSPL2C63lQ
LGvuV3aVYLBLCRpmcY9VjpY/AhI3pYnrWiNEwyZHrMJuDYLtcs+DzZLyXcrX3EBr
x8ds+vEVO5vTr8L3R46/M6OkHa7mxSmspKdJ+w0gn6xWgYPZDt66ONujpqxx2Bt8
WNaXbXJN+poulE/GMpseV3zQIDUVkVyKojZp7nWgVUHAyEMblyrSf3o4QZ7fGoc9
yCl30idvUKsjG/zo3mInXx6C2S8i1vkauQjYknROa5SYsnPSZtrF+clWrBz7UBhx
hrDJcvFC74Aeoi+t7KoKrim94pTuZvOTXwF78VZD51HnsLneMzRLnQQvmHnm1Owu
wzE8Hs60wrRLTimQjqkRlJuPJUjSEsg+I4HyZau2Ni3hZRqCS8OIsxz/D/GgKlcP
DCq9ziSb/P3JpWf1QjfpW7yEwJH6702sgqRrkJIbbnjQL6l8rY1U00eQL/PkC93i
VOolbXeD7+JLEy4+8n4V1RTF0wudoSeDOwpGmpqlc26ywrbgf2MRJf0Bq9CjYPRA
piAX0KDFfMUFonUEsxAPiTFK/YtKg4ntP1iddVsf3zUEvCoR1men9XP8ltzq2b8d
9eRWmooYHZc4H9snuSiE3M/8gsqPIyiGUas/btqq+B8Gn7bw1ZV6N2e2S9JbcYtF
QtE0GVkBMzTMqm6WEpHaiGJinSudYNPpk/lND1xCIfoXpBsk3d8jyn/JCZw6EpK1
RwZgPzLovhqixa7JiS3nNATbOS9XggwRDVEDoa2Jk7/xQ4nBNYHHWGli5ubVSEbC
/fX8Y7C6n8FCr8FTPCiKS4nn78Vlf3Io4cuvU2kUPrgouv7pdSb4KYTVP6mTQBvu
w0A84vGb1V7WWuHbjnqcWyGnm6jJuxB5sm6LSteDO0vwN7sgR9spix3TmMQdBHfm
VwBxLMKovtVyMtDkf7fmKeUZl/UJMi5nIOOHsgx/XfuWYC8P2wejIBKCNxbgEac3
jWQsq+SCbWkZO7BK/UbE5XKzw2b9Cscgye6e82oOMZxHAwcYsYBXoyQ56wGESuno
w9D2s7tJK+/Fn4mx0OKB0zrbdt93oJGXWq4SqDGa1mQTW/tYuu5q9St5ZHEJ+G1q
8rujLAOnG5nop9YT0ETmB2It4GYHHsbPVGYvnJhVigTfQvXMOn34xkQLQgkkRBSr
YozHHvOaHWQsMm+E4+cV1UQTFcvPIdT3GpLIBZWm+tro406evFUrVWkS9Pa3g7UK
jNyt6rvuAEj6omQJ4Ubze6jrLj0Ab4cZ58c0ks/4JF5UatBQqr5XxuvzySD32pX5
sCPXF/A9zdIsY1halKZXon1lHx3x+zrIQehE39LXWCVnuU78ZRiyTcYqDWHfbrps
3WuTfs1S9/wMHa6JbyCQelN9EXqrLvNsPBESiFWTCZqVilckYH9O9djBB235ticK
/laVQqF/yJHlMICUokDUAYwtIz9LQ2PwF1JBu+BkK5eQGqUhsGj30XYA6/pUe/B6
KYklj4Ou6HAUw2j9Fo0X32/c4WvfQDGYcgbLSC3Q4XSdee1oEp84ZsUxs9Wp/0lZ
EW5q3/pbKe5/HH0jzkyOor9qfdCxJrTHRtfJj3+19Haxo+QO/NZsvZow/5iQWUqQ
+O7YuRNxV9sd/R8caiD1L6iQjn7JLNdoFSmXz1rTk61o7Q/OaOIGuz3RLgRAyCNk
xkM+oZ1kmK90xrSpvpu+I5RhF3tmtSqmJYM3S2olGXopwRl27amet/vzNWFcwrAZ
1Ed0g7TAimSd9wgbX25x1yfzfw5yRggXQKnPQk4nb74nL5CbVbNQiDLKezvBDLI/
Rr8rgMKHKBAXkhFmwpyKKIoJhH92xMquyJpsFCJYQdnQNkDDPaiU78NtHxA2hk4l
mzPduNz+enMaVa/UxLChR9GSfTlRszkpK8WkM7iPFvEq9BMSvY9D8CceMK1M1UbG
im/VEc6HNyyRn1fvSeOcDxJ+vCwG0Svzile6sl33PxS/XWfV29quvZwetMREHhlz
XP5/VsbAr+iJ7JjSFlNtt/fJpVRwfRCI4tkxVk8Rvl7C4sdiCDEPVadpHd5l1qkj
BJgGj24GfKwWJ0YHTw9NjyW80EtOMiE4nlwB0W/yMIw/Q4EA1VOu1O7kLluLPdR2
iMyj2WCSlk5/Lw346KabMJZff2PCwithnqCaVyRNnohsMgxIzAWuEs0LQvPd+yML
dbgFn65j992o0nZBmAkEsfXEqp6LY9HCl6S3e6fxK9QrkFIBMEaexa1DA8YwtL7X
4C0JLpvWyyNxyh2ABg8g2TqAYhk5G/Y6s1ncL00WAzFM5sOBba6JMGW4ao702EKG
UzkYOuYo0HpV91VONuoe1XgieXuCJVV7IkUgNH+zFnEfS1jwcrTbHiz/mDVa7rx9
dwZ4NrzI2FWB1Ky0aXIJekNDb+92TxHYPk37NprWIRkhAuEUgLdNqgZhxXijcU7V
NGyTaHe2AAlRs6x6UMyfhvzlLzSI8LjyepMEWg/BQpkFx+DQUHgHIB4En/vfRIw2
FBPIULcBhHG4IAjbTTfFZ3jvTbNyAi54jHTpltpKC85J1BMcFr4ESmIJTWnF6r7a
a2V0vVwo9VR0Va7401tuhCGGmnX0V7+BbAd3keAxsqPze/2Dsg+pHIg91vW5NFhk
WWypDYFComASTfWUWpVqRIordDx1FWGD0+I0ptSL8smE609S2Iqoxn+30PV4Jx3C
+lbiqnefna7S3tq2pJ8AIQiDpQbgkGxLp7spPrFVWmrfc+AIc+dfsfhdcRERjHtS
2t7pSneopdkqVIBYqzRbiAYoNO3BtzHFSD3cqta2SgUUKaAT0KoAnOSdsWJsiIW1
9SAQwX5azQmDN5kNDy2ZbP5sZk0gyxbHksW7D7CFO0pKaezr7gFAwHnq/pLtaM9g
oMOoh9uk+jQcteWKwp3/Hqf29hGqrbvW1U27Fx3SIu7D0Q+g/lOj6zl789zSusda
SdsOIy47uUoc2IzdISHrbmN560G7RtCvyePdEyWvZkQQCCdmw6P+FxHuCq9zaTY/
Fccekg2ypL6QDKF7WMDY5EZloqGPBWsEdMxCMkCemyQC+LRnaf/rUK+GFk14/yo+
L1GOI2Ww32HHasHVNTJTRQZunQllD29SvaFi+f7jEi9xVem8Lhb6MBqCugMKTsCP
j/qfsmKOBA2jWH6iqrDoHJUkNPcvQqHlsNbGfwR6GvQnYdnHY0R/jHTZHDioQ/jS
ekaaermRSZlPYmJR+27AKuP5dxkDQ13TcZJpn9a+HPeQl7IdoFdSlbllI47bSjbA
vR6ywlZ1M7oGdqjkDpVwfDnwX3hOI8cJfYsS8OX+dFLu/NCowxBrJAxyA2r15MjM
GBo6z4B4MbpKPzT3QmCV8cplLk8eD0Y7l7F9h2wvdWK7lM4C7e4mwd+0baUK97wj
mCLLjygCiH/Q2+g5bJOcaVYqJK4ZLwgWFWC/j5VQAlY9HWWqkW8oRq0O6i5aIgN/
RC91O8Fp52EZdHEZSL5t49DMnp7bh3ednL0BMq5ch+9G1jV6fXYPm8T8Ota0hMJ2
8MgHTH7yJ7mikQ62Pp9M/XkHqOCLGbGZ4hXqv406odCV9g5dsTd2LDNuIerhVgo6
+gsZTxKV8U593/obHMSoW+Pk/Uf/990050Vy32iIvK9CAesnMG9SPLV1vvmwRxsA
gcWF4Zf53DZQK7GYDk0kqX2BvkTG40rrSO8oa2AFS95FWJwkooSQNO5jvNuOONc4
RKcZkgE9mZ9g0D5SOSsqQRd16iavhTW2eccYZrKgM7ZwBluR3+//vBmJ6Nj2qAeN
eQOWK2PRtj5JTuBvzMeeflPB3g+Prq4ThZu41qP8oD3R9rB9RVHN5jb5NQ6EqOBh
Qn7SVCZiAkYbP0RTIONUYwvorKXzwoEVGG8Wf8Zwr3Jxvuzx2e5YpzrGGfrIH8Ru
q6gfp8cXtFiebv03OKnBvVFKlBwPoGWAwCHTsyXehPHVyOQVdSUhNflZL9eR5zW/
LjDpbT7p0HYLfEBC/qCJk8w+I9ZcMUZlG8BimjibRpEF+qG8Tck9BUh+ssD4I9d3
yFymbBXInHbO35wL7xSsMaYKqUzI3sUyecSK5z4RuNIUYceMFtML1oD/Gh3DsFCY
D4uIVH5bex8P7T3+WuYDoxAJD2tQAEqr1bP37YLaTHLkWK9J98XGAljVNSgDiLl/
6njtDzzm0Cb7SRf+Xma2TiXsqFzeGuveusEX6IJwxUMYMmwZdfC2kx0IiFFRd/DA
WyNMiAtwWGsgBCJslTB9UNgFiBUMHdHUE7FOa1IPyPiq/kPwh2ySpMLk3ZShsmeG
BWhZe9hV/NtikCB+9PNrVPGMdLYDKR9xxCkfY3Th2h4arsu1ynBPpkfnRI8w4wAW
B5CYUPK7yI0zGW3p0DLghweBznaQyPZb/yNFQkeTtIboI0/wy3ulSsoMMOAPGEth
GqXUhOkUWaNpERnFTLNCmdt55L4zqyZgaJunaK+APTGC7zGGvH6yV5iNuFVTq7+N
+n/e6Go6xVTHMJZYwhTA05W6WBkvHKvxrW0w+V61uAqrQaBZMXptEKANy430f29e
/iT3/LUkuPn9V3qdD4DKnrEFpu/+QEOVJgwLqjCIoOQmCwfSNMGQLLwm0D16kNz5
IsN0fU/MPSSd6LZIWR886w9d+0EZI9YngoT9QAjly9l3H0NDHbrh2AVzRLgdpmjK
N5UTConR+XzUFO+MbCg4B2eBbC6vSCCL4zQRuBRCDxFqMk0tVKQo3bbpcwOQ4zrr
vj9dJulMiQElRJmBJBlfaxvBWCFCxZjloXmAzAFt9s+m2wbvRsgI77FY8ugSWbKD
XD+M37Upxn6l2OFkLNzHzDE/Vx/2qjy4Rn5fSehssJhfVSIT6ACjxpFGcQ6WBnNa
Akg+HeVX6i35Q2KtX9TELgrOokLX+pHZlwkwVY1sqV7aLWg6CPfNPIuT/ogH07Ka
a+xuDP0q8wzJ5e93GrXLmS1ngLFMw8PpoUflCWKz+7EWzO+oMkHqbhmDhXwVI0uX
FJfCCxCBKuRBaB/vjDcYj5NePcOUH9SIdRoNvfSyE2R414pAiMnn9YQCsn+6032v
BmFAg4wdSmjC3fe9TbmA9fh2mWvR9jFRxZyS6D7iC1nv+uCdd0l/mzMdKuhIQ3c4
efLhnGZ/h2wkfpIun3O3mkFTJqzYrCIWpeycksPJIGkNlY5J/KCSBQbO22Sog4Qr
dSFsd7RAJvEMFqL9pDBCdT6samKJhKfDP1HXylYxZm5GVKSWXu/m+OIg61wzc66P
Izi/MKEOtZ4wNKHoSJ+BIxxX2KLLHil4Y7mlI2Ozv37LTyy3vDiqv1Igh1tdcMcJ
znJK5Ft3LJ5RcXxRLKW5XpQSvCzDEuLSZUM3f4qcuDb4GA1mp0cPAHkOgWri6gWG
Qbz4yMdVlWDZrVJih7lLy7U63nqrUNP9s7IKXTZ4u0Z4paNIWczKSu1Ju+grhvs/
9+3xOezmEVqh4hgBicvhMiHyADdWQU3aYrmBim3MyfbptXH9AQdQDre/HuhUTA0t
0CDhYNUhYPyVYnrcydAMsYDHu3coTg7c+FyzlsMnY9w9jWLLcst3S33MzjurlYVt
ZWrLfSNwNTfvns80HvbzNYVEFDc77TARA2tQDxWTQiPyXJqcepAwnfjmhb4Hqmct
JCLm7hz2jL14B/nYoFwnJyxvNpqLlIJRF5R6tuSQSN3ZFYRCT2MCrWxGOp4Ks5MC
hovRRpcgITWsJWfDVkSXK0h5BIMyNeminAQ8g9F+kMI5R5DoyEkTgIkkoZDk7hgD
B9WeiTAkzzts0F+eCXqKDqdeIJpLvmAAm4QlaOX9ErFMB1KhHh7hPEEGwcXRoSpt
cXWQAGRmQ/F2O4tM1G6HiCrHBBga9PJYhE0JpvS+HSZceglyyXtM0R0lm/h/NE4Y
M5VHZPOsZNnzCHy+eLtFECyE0xwOKTrU0N+oPV259fw5/3grcnyVG5HjcYFyyWCC
WqI7TlhUJWy9N9ePlvANOIvI70KJTJZ8VhpF9usKgJlECdyJfR/ZbSexyIFzstMf
4SfhNC5EfyJRHCKimKAccarek+RDIAeNkrvdYRvBr/yg3yA7YP2GRNASeHHrRUgn
mYdGp+/4M3SOHHv1I5zEqvONcibRAIBizgg3+TsIem/PmggmV5W+tFmvn6nMkH+G
tgtWIty9grJwCkobFO9UfQoPlSC8mjW5e/7vXQhKxYUrp9B1rB+qZB7xvsYxJTxG
q6HUAU+PygIHQdwqQoJH0dwMLBQd61CBeqAnclqCnArM0XqjU4zTCNbDVFzJupNe
mE5l1c+FRUoGcHlFHRZQ9OCYN909sANjhk2UikXHSPf9D635yLo/9zLUAJT2CHK1
k8TbckrUojjlCEpCXJhYKZF+c85X720m5Ie2GY6Id07xzeAG4G1HXNXZgwy1Qm2M
/xaBpWrad0lkHrOtRTavYAwWEKHBOEEnpZ0On+popwUFIbgu0RngiN4tjPwO7blq
YyuHIIGt5DMi3ke1lNg0gEWabzlnt4+FL8KbdlT3g5va5nj10lZ1FvmXi4vwMdVg
yhFSqXyAqO0W7buwjupVNcvd8FH/hiGOrYDjaREoa3CpUqjLWbchdOydzZwBN0xj
IZZnvH1z3UBJRVT9q3eqIQ5eL5xGU/hBGLKuv15EgUKnEw7dk94+BhrjbpF6uWPk
LvaXXcXNsuYIAWnz6zrA7J1LOcGiFeZjWAxNvNSLLCMNJaeExlOKVIvbd27MzLR5
iBhQqBtieeL22Cje76lN5W9pcTctWbHHNd/mTT95RUia+6cH4u3bfPF73oobBsBE
ulUaYBqaX4lGxMNvf1IwQ8nqS5jbcCx4cKy87faLAv3ig24oRnSU7dHJKyRbktIF
kFdLIbj+/itcu+z9rAleEmuDGSp0sBzNw8sX7/HX9PqP4DakuQ6QJud/8ak75kOY
YwoIqCAerRqd4Acpmy7WkqLgw0+w9ErLIwrdtTH8oiW/q6IexQmx9wovbLax36MV
nn+nhyJq8PJCBZTnDzCnwYCrFD1dh1B3Zy4Rc232qoojtRz2FfSkzN1CMKwe72QZ
LH6EkzC2tex1+EZQViGJcgY+I/TuQE+hEyp3z7pwMDwnZTNQk2NgFioZDuTyYjFl
iO+/jDjc0T0IaPj0fjchcuyiRQckYk6RsVdzywJAHjWkVb6C395AGFXjl8aTFBcm
a0CXQ9oyVgx8Utai3wS6PlTJlU9o6RRw3HKY4wnn2hEDnrGGAUff4P5Yd+VknvOQ
VIWJZgcU+8zFZpqier3GqeyBwGiQHVPhcP3enPcO/sg/vjAq6s04YBAEg6b1/X7y
bJ0yfyfSKwdp/3Boa6dsEkxdShR4YspjWRm0ViPwKdz2evfZD67dd3ngctA4TenE
68iK7EMjl7a6+ikN0gcKks70Dr5g8FsFKS5+oNXt3pQ7fzCUwRQM+uoqgIrvLPfF
EKYwpunmnSL0a+xecip9I7Uf5LM4Uab6/fTeFEtk1ccR5fzpXMEWaFWy/M9E5ndf
X9Fh3BMbV+fEJ6sTtZVsZ2ZkZmFp77RGkSzT+07WHb++faDSZuvuHk6xinlz0Nwf
q6+Q3rNshHwhtrQFjI2mBDCMUFH57yafAuo33Er3OU3NRXx3T6ck6kTdAKWJzq6K
3tJfydGop+rxE33Sosng0J+7Cc0BVWRKiWg2mAOIIzjklYMgLawWwfw7RBzPlhBD
Xvx9lByknoIKld58tY2qwkngcfmtYi0oH6OgyRG+29pxozDYRfQ2IRAYEwdkmH1l
hw9ShQfDBHV7kvoW1zqrM2FExZ2j4qXrEtDmS86ehhaw+N2Hs0dQUQE+W3bi/M4P
Mn8nbPf7x4QQtNT8SHd/BUAZEJ6Pn0jQZQbMPB3wdFaeL0bazGL/phU0RTukcIYM
lZOOjmBR8J6WpPmnK7q7ej+TjYjFjecMM5bxgla8hSdsbbyUx/gKnEpY8hC/6bOd
stHembFWmShFnraIt4UeAivJugdOcE1CCBagdxKfBSUEHCKndIt/8FgS97slA4I3
6ZO40G+FS6ZX4gNmcka8OXLQbGpCIrc5ph+YTP7ca++/QjBdMFLLHFQlVyJxsVuQ
LBQWmIkjgAA3SAbd0Gyng1GRq6JZTT9m+CP5n5mC8ZnhJA47s19RODE3gEtZcqQ6
Jdubm54vF0duPFgf5qcNnDBS9RnVO/ZG8FIBvb0gMiq4bb5dlYGdaKFykHe+oiWq
1r3oLZnjhLbeCuZMqtxiM1wsOHFQn/2JES6TAinB5CfjOnVCxAH7yt5e7s/cpkPg
eq1XhnaJm6WP1CXnFOJYpWlPeWsdUoYTOfYKuRxyiMntNDTS7ZZiT9aQdvAQeotK
eSrtaDlbVWtyeuEotctYKBgl/qyO+Z9N6MMCJzIguvPPUkrRTrQxD398Maprpjr6
vKSOKJottT2Adi+H+ymdh0tyRtxEKrotkyllQ22Bss93pQKuT/7kx1UMYA2G3Prt
v6dJZNBTrE8zABwPUMoYOFSrUydnHhKmtFRvzZGRfWoEJ/1ImrjAUH+z+CK7z+fL
y6jTnpW4KBHWCOZBTwJkAY9gttCq53q/QxzkJXo7lmFGmhEJNMo00Vtut/5mIUBQ
cloIbjhdGm20iE6vg8Dx5wArjcwFOYSMZtnDMazvq1peoBuISw+ijwN5MINxzZ6M
4bmMYm1gpRA4xsd+WKPw0m7BxSj3axcInfNJLjLolktpw/hdIBOw7myYY8FGcCf4
i6KSC5ihGmAkGCm51oL5BB4bvP4hqukZw7La1x6eZiROVaXClUmZatvNsjK6Gv6y
c153UwKqs32WePueNdWoMTYAK9sEIgrt1KxWwpEn7KHV9YdJdmY1eRJo3Et4rs3C
XCgoXrysidLHFVvkKXF2Jn1i3MMvljWUZgWk96jwgVIoA9llmEGAhhhzCfE7sKAv
PJDEc8/GW/zJJ/zQPBosRg01Xg5rDJziC/IR3EyM6TjkfeX7M8PI+6NUY9YaxMcc
9T0vmrGVXTrr2EXgs0rxPKD9eliTP7EIlgeoaHC3xRHC4JiJe/qj1Lmx5tc9I1Nr
Kz01+in1v93D3pKQsd95QF2Xsibx+6xYnV6ps9CJjzU9Z7VuOdya8PdA0tU5BBZC
ixV1ySe3nI8K2JfSwjnB7rfsYmn6kaCb5jCie01QHYvxQbsLnS4/ouFwngoK4kLX
8RXs1jGQ4lK8JASdkTq9r+utWw4ClU8w6K2KKJ+d6cN5hdGGhElVWKVUTEqG7dpH
72rk/blnM7Qi/JobAEXAl3M112n1rD8SILvs8GXqVr96SfTXxeKWqf+dhgF18HSZ
HHmqXRKn2ApRtKMczSogYiO1oAyw+BDMHP0H93e9hPClfcZ94lH4tc7FFp7FUN6I
/8TZyqSCCrzKuWjFcOz53ekDZUnNOeTfjjfQGizO5X9/Nna7dLz2kaa6wYgTuAWw
OQGtISG+rLY9CG13G3iFPBAxNdlf8A1kS+9pUEUGFZjiBTUNBTO+f9M60kFTJhNo
xwM1lfTu9jtY8JT35uFCnBxmhwWQM2mDAPsUsoi7iByqcRcx4JB4iUANnMpJ4Rwe
JoSr8pzq5r18Pj2WA+Mbf6FvvLUzAK/mlXDfMDCBXbij20nceJSlsKWgbBQ24MZo
kCGeJoT1sfTYcZAnK+LW5IziX9BtWwegNonHEefl5Uq0WHaNALrtjPif5+oBXuaQ
LAFp19tAGusCLcww1qt7tcUbr7PvZcBordxB29fEp7YaziL41hwe28qJyBb29prN
Iuqj4OzeHqCM5sEXgRH+VR71Il2TvxmVX//8qlp+t60T4sqb58eO+j2RdHXTFP+n
FZ5InusMO7+A6a+AWFzpErCo7AgSOtHWIQzBBRnUnlDjQ89LRNXLfzERPmFiso/p
735JRyFJfzNsmuLQZbq0jpEIRxt3pqlf9cdZpd9k6ktlRsGPyY+dkuLUE4QgA3fZ
iGBzs1Y/qg7u4qv5I9RQ3s+5gF1xuCSFPkHY6GvQ3ki66oMPLdX07anYHASdgb5A
81Y9pUO9fblPZMsHKIzBSz1+sjDjGu1ZDnVjsgM4sYQQxA9PwySWZt7p/fvkGVZo
qZvg14ZFT61uPab61gUQTPW/SWGMCWt1Hxn0JP93Iawno2e+GzhMJP0OcI63ihso
I9/ZHlJr8MNjZnQaJMwXgfPjHw6clDRVXkW7wfK3W9C6uqkHIeamV8Zy9rOAxQuu
HEJwzZ7QWlyvQvGQGLsNI74i539imaIT9QhL2wn4WYcWQz9erpxY3jMeR1GRr48D
6GjsWtoQdVTQcJM3VNcGgo02Q/SSlCxxDDn2ffF7/iXJAojy6QhlVpbOAgm4HMEf
fvvsoGM05kajNe9WojPyUxPBi5IzG1E5HuNFbiZmUt3i/HJbkh6mPhsu28E6GuXv
8gZJVbVNQlM5fr6SP/H76b33ejyvtEAnzPyeyE+xMxgWMuf6CN7YjuavqVQhOzKA
6kATVWGSahIkUkVkwf1+z89uluk9h/gYHcdxsDE6JyI2hyFW7yp2Mq56EDjBN91Z
uV2s9YV3JuDaImJ3GpVtbOGbW0OwoR+B097rY3YFmXj+BFnYH7aEjHSo0gL9DKY7
4OOLze0y9v0bzLK39kxLL1QMykQKU+wRtwD6tvmmsFcS1CNK5mfK89bh8A7AnI2R
0JJPUo9+MVOhBbhao4avMebbipsHpQSYI2HLXo3sPh5wugYbQ9cYlzWB+JqLIHDx
CL2YIQFwvUwPmjOhsLG07uc5AUWHsL/+vyiRzcCr7eN47HDM4v22PhiRwhoF3LCT
2bs6Htzjy0hTjpDHaHVbwGW7OO3xdBpd2gbpIhFdW9+B6YeKqLTWhnwx+/orDbUJ
4EznKxwD7/z8byOnIJY3Qkrr+geTL/CWY/6sxZeqmq5rgtVnV8sgbfituCbqSl1H
4nfLT2g88WD+LkD6ISCAaYp7ZHRTHNNmUFCzojOMhA/wPNWcUU+GeJEKFIVrqurP
lb5zsEE0CLx7jnBbrQAr7I0DNgg3ml7Ec5vHUdAfvnY7+kiORpqa2gT6Q4J9FIw6
M6p0o94p6duuVXIYmXFqCBxz+caRmwVVqoDkVSyF6X2kySg4+wjSvlPYUcNbwY9n
CSCGfDwr/MwNMWrY7FHK1SiMSVdaoiZ3MxzoVGaE/KRWksptivMGwY1E0G5fz0HI
O/+Kai7LKs++52PWu9eni9Qi3nsNRyh8KPWJ71d+pIenlFK/QYyFU8GhsvDgmisr
+puvw3qmWEj5HUXoMDU4ELTbMPvJnRP8k0By8f0J7tciL6AEnYVN2WQfhFQrWMbD
EQRLjyiqjHyRZo9EuiLvcjo+QE9+2dGdB0TnOknpGnJA2Xu7WgDEv7pYDhf9nbeg
LMVY3Q72RVIaeYEJ4cVlEHuVnsPjsbicPVQVkJwrXYH/+Jt/rxX+zj2PFR7i+qyU
YlP9lSuoKH8U12U3jv/ljDCb3pVASPKQd26AuPucLqpm7COF2W8Gx5fHwSCwUVn6
tV5Fwzf7o7fR56YylKCyvUYOlJXISFfsjUZ6Td0AeNiDCbDAYSWoIAAh3rXKn5Ur
rY1RIBvfdsFBDiK+UPQ+RperfdpzR4xrNLjfue9YU0T4AV9g3z6KoMfKT/ZU69eA
+458LNrGGA4BaEaMCVxf5vci4368YG9ICcNQntLyTE0RB/r+spxV0q6KUAi8BSpy
JjkqJ9s/5ZYddUCC3Nu+D3jCTZ6e3fEOs29jupeGeDT+VfgkCfkilqs8aSU4J32w
s3zXTQkX8ajeG9UBnzoA0pTaV9ZOS1PyXlziCKNsc/YBERKQVcZlNwyfsssa/54Y
aQfISxIwUAjHkCQnuuTQ0NBQuKzNU4ItfkNSrP4wQKYB9c4u2W1uBEUOjU5gLkHa
jBpa1p0/Y+DTzL6fG0BxPev4+n8SiQ6bPZZcmCqdBkij/FTAriJM0ky6WLrKk3QR
ZDptSsExuHVOHUHGCWUl5j+WiBqZ+LgbyzNMZSv6pAnla+WD9U/iA72AhFVr1xWb
5NzSmLZf0B0aZlIsTwqDYD2gGznDRZPDjFtB/p4Q4yY5gZ/pjzqP/rtWs1K7sVve
ylf2dSRLYsjpFPCbANDrUQalesIwDO0vFf/WOBMt8ucQ22z95D87vPG3LnyNh+Ik
rg9bZFIH5pLV2R+spqYOT55dOznjc2DYRneoM0X5w+RMyLb4v1tPg++aJkkfxeui
XhJhF5tC8uqWkio/RxaZ5KYsSMNhz0apM7/huqEGqBg3y+TqLhYCAVkm+jDH8/sI
fv203eQ6/5/zUqaS7jYzdys3026ekbF+3pQur22XyIpGe+B7T2wy8CmrrxycCxAF
GQXtOVmrA+wYkXZsXIfYFkbjP0kS+H0JLLzskxYL4idvUX6cop92slimXKAROp1a
iRy8aq7xABuFNknohgFwXF3Ox7qxq1rNb2bX4eQ0AaSnndbRfyASoF+5muRVl1OK
x8TyA+kO+dXAJWEqUIkFPupE0pBK0qnr0A2Hr4+szFU8kS2ocw0j4VzTjqCTTN4d
+zsg7uGpOVERRiBRgctPqFQ18nU0B1N5tJ+xqD8BDa+b6fCMHR5azMkZv0ffqZZi
sY+2c7fdt4U+L5FeFR+ps5gcECIlfYosVPA+KYt9lBUkPwA3x3j9trWKDYFUOK6L
mhIvLeINkdBPRqRlKAN8LbRU3L1kQqXCMu80/ldc5UhKijJwRnliQHwg3zIrQThC
xY66P/YBM2v+PFWbDGp+YCsI/ZzxCpdrzPLO+Px22mpoL31EY5elfyWPSYt4qs+9
nV1Wak7bYEmU03TZ6A0/mFSqdhUqPGXLf2k9bvaYem4YJeuaSDFwvd+lXjvNT62L
q7CCvGcw0Y2Ffxnn7dVTsDX1pRh9VSnC70QQp1LzyJOEcyDYLLbc+mPJQ8hkKuXZ
BMyLHSWk/NF4RY/r6qjnFF2qLPUOPTZ/R99yVVxdryC13s0OxQc4tPWJx7Erupvr
WXb+0zLagXPKrK86pw6zELXf1NwiwyKq/a9mu7j7/3i0noFH0yqJk6db3IfSxffb
mHhrfA4f4wGnf7Uxo0UgBGkQ4qs0dQdokyE+v3xolXRvsQOy5eDRcMMZyx46Jby/
BjpwaySSkYwvfUlzWyOkZaAGkcNfjRREOyHspVU+9VZu6zzMAj6Xr40W4I014mJl
GHvHdB9XEag/thsZrUmIvsMT41U2mJ7a1KRa2BVuX1HBRyf+c7tP30vOoc1bwCfL
OqkyYroLAXV7hz9MZTnzW93Af9Mh690qtat2wboqoh4bTpsjbR/aeOa+Zx29lIBY
34v/Li6f8lv1bpw4oaKCOMLEx7eOxMvNjAKdTi2gNHebVpNUMocLVQKAUvRIRhCG
yyB+e4OHMeAMiC7GUJocEh6t7tJXQdadcBo6401ULeQgyiZKF6VDSS29D8w0eKkT
FDPqZP6jzILu/XBhZDkBfbgaqnTYGCtoXnwge1PkCc/9bCv5HRf9n7WS5tZgqHY3
935OBlN7/vVFpcB4epCNazUEfbgK3QoSigoe4cApycjD588Wupqaz1R2cyXmjdd+
6jv32DCKBi69BB1Fwkld1Ckk1go9bG44VpRqczhIMu43iS7Df6OLjYpiMXLLC52N
9QzDo0y1VHXZJ27luR1tquPnaZLXLzDHdiYL5lFU9PmMJvW0RMPhKIM+g40g2JWX
jlXdQpxgD39FVN3ENvNhpO9FH4/4yKnEaMAfUicURjUfnnO0WpxpODcSp2uf4hwn
Lcvv5tBBR/p24fzbH41FHiZaxXBZGFeAonu7H7h8MMXnUMap5BFqFysY/6WgVvSw
w+JBOuEhlB9UT3zelk/FKUVpi3yEy4GJHgzwpXa1mqd15Zq+Z12S8wPu1aYGmN/U
YCDjWD7YUXm+nf0nIDOzK9BpdI0aZtyEXNPRCnPDtcOaeyaNlzbKvfKe5iej5lRv
ji7MBEn4g4zbDj+eV4vMrgI8p2oRwvwd21Spb2mI4mM1i6UXVXYxfvr7QV+FrEPF
oxaM1uYsj+uy4r6UuZQgGtakWYx9LaaLQw9+qS+GIcmPYayokizta4DaY4SQAuij
vZ6IosmZQfGMel1F49PJcVljgcIpGfepadroStAGa3d4CXetFqSjtXrvpcJ3Z8vF
NE98F/VQHMrVoLa/SqkoDJA2KPmg7+MbyQtPbI6gg2vNJJN50mznB/pgdlCqmadA
HSzxELZtZXGaoBJEQagK3vq9+O5rDVaDs0elg6RZCk2BPrFgq4RXWld8zjjoMoiC
TN3ABcSa6gQZwx/lBpQpO26gqwOKk6H7ixr843V2BpqUUn53jjBEue0NpDJdm0K3
X4gwC/zndDbDzSah8/cJSrcMGfvBArLWCNivdSCW8Ab2zacJco0f5reo8MpTuJT2
dgAhZazj2zhePz3DG3335/Bh1NCcHwd2J1AM2VVgJObCqMH+Yns7/wIGc2OZtY71
g+ATonqLr6oqym/iOC2J+eU81JWXwl00FtbQ8ECk+EI8+GP7ka9BzEFJ5R72uu0g
M2xkhsI/WLzH5B6eI2qCuVlGZCxHtChccBR3UUhEvNuHHeKFNZJRe4+5ytTlW3Pu
/7loj0UO4rKEOGsSgmtZhiEMd2G7sWVGZvqud/DCc7Jy6pwcR3Umz/Bd7JWpkjXl
359AV/GXlM2Zj/NhZ8P3AwvBcCNLWV0Cezii9Vkb8KnM3ZkNlvVY5PBpvZtzQbtP
3N1M2MbmB3ir3v2FK4w7ncWPmly5XYAJkKGEt+n3TLKbDnkJ9SZRJXzVpCHtDXU3
b+/koqolDnWZhc+YU/X2Lxd/RhgdowZBjdrKWGgRhmoZYq7pYkb8Ahpgug5/tmc7
bY/v8qj6y2Bk4ywUiqCNW9Nr4Zart7/r+SJN+JkaugOpWLhwZRvKm9YL2E2HO1pD
ekQN9UxtuiQg68rKRJvQpyQdfprP6r5ih4wXYkkjQyDr8FqVTIc6FU/nw8xmQCuI
X0aNOR0Nbq7kEVuEsS4gQv8E/gERBw8hteLymopg08/Vzkk7KgVQT/pBZrMfA8wJ
cWI5mWIC0j8kugmX3jLdQeAopqE1++WE0zT/hcR9U0ypm02SOYnYd2Qsjn7pvVEp
9fvmKUMfUfiLrCDzFXNwB++dqA+dEStrzKH04mffSwLoM+lmZl00J4T+KzmJLDih
+4PlpWbLUttgTI4nqIwrk+RGn1JIHs9dAhIqVZYGaneT8ocbY9vyDM1GKHNWoOyP
un1rCa0c5OyRBQleiWhVygep0tSwFpknLKtvJ1i451whCiw7EuE1cccOrikA/PjZ
A9mY5N47yogWUL3BSRyBRyQePYY9pcOvO6exgedNYnVODB5r53G8iOW1e1+IDSlQ
y7i40Vj2i6nt0lQq8WdkbID6iJ8MoMbSA7xYP644Vt1HiweglQh4zchDltMckDVc
lXd1BqHNZ62t5hA9nRTeaXILeaT71uVcMm4i6g9mbn724SrJi9q7+BbLFxGR2Ky3
3zdYKC8NTKfyu8eRhJJgKsGNgJrlioVB1TE7VhHK8AA4DhpJ0Tv+6BaKxR3w/ooC
4e7DMXAuL3RNqiAdw59FTln31mFsIawBxnDrqeqCW+XSzPRlF7WXUqpnQaHuVKRr
TcP6cKuPXpHWF1sfLJBtOD3VtmJ+rcaTcqVsl9hQ64VJX/5Ezqexlum7ZgMgWvuw
Xosv2y7j7nZrt8sfxPxdCTA+c+jjKWWbsFrZ37OnKiStO6rtKRbmiGnnUsoh831H
PuqYUCpvmXrZVk9j41lUGXrzgVw9XpMGv+hBZrJqi2woOtUThTMTJSL3obtrKGQC
Te0e3O4S9FwI13Rr0iSLgQ9fa8m/GJC2WMtrSVpACzkOqHDQPt0CTNyREIXXThym
q8Kcgxb2wzhOayqMOQn9froG9xSfW1go07b6sE9zfR5x0GBTDKK+H9+eObFa7Aqf
QKzfcBMoTu8OtSXu6bK1snUet9I7HXdcRUaZd3aMR5RKvN+K3Xc3Ofd6udZhwVTd
l0pevvKncrtw/T+B9StKMP1Mg+z0Di5L7Jr3h97andrYfAFyJiBzCUeVsC2ZPSzK
jtm8TbaQyUamLXNHAR9Pi+vkNPKG0bUTNyu7b9fEsEIzfxkMhpbdtcXaxNeT8lTo
aaX0jUrNFA6DJDfzhjrP4+3zEg/QVudaPEG5U7DTAIgj/n4rpjUDwME+mZmxkLQG
Sl6QxYEJ5/LUjrGbwVItVehxXEjfoFgqL+F/PHGw7olx8aZGENdpCtLBHMH7f3MB
3dfBCG8J4MG8GJ2dJiTSl7z+b8LcPEYoiVrfPxKe8lGGpivkwXqJXGJRJHbXt96i
6OHrtrqGat8eeUwpmvtmLQRP5C6mUdk46uqwE4y3bo9gY69PPKO228MaZ8Gt4y3p
1fKW68MBCG4+gVbThpkn4NtxLu/EuWSXWfU84YBOEEaWSkSU+GnzJgIxYOcycc7B
UyY35qspHrRsJoNeBlPkn25vxeupYuEkiy3UZHdGa2dn0eBfuRtUVstj5+jJMIU0
5oXp60OeULwGtfEQhYeLRThB0fjwiyUnnTm+3X9y2R5lTD3xuDEQA+iCXOZM6bpn
b9uh/lj6BuG3ByEMpON1ZodEv1QX25FLFb7FzJGtYr5UhchXTfmK48BXeHkP62C8
ZzUi9t6sOYkr929JFvpUj1ge8LVP5Ra3C4B/qEINlUl8RZbKB2OVEe6hKHu0TPKt
dzN4GhCm6U/8LsT0dyngunZ6dg1m6nlYRqb+BEk6OVnsYU+fSO2SUxXtlnCSQwVx
6ORneEK3t0XrohVcYdjn4huM+JplC2Bq+yfw7r7zAARFUX0wnw5fXvf++m4p8AkW
ik1VGpI3TJBwuMBZdCY2xQ/UkgvPkzmqddEwIUB4ovGs017w3JysBrtCtTzL39Av
qV4ypl2gQj4aNe8ID2z6FDtIPQcakA8d7BCyNQl7qjns6MW+qMf98K2UFwI9bZH+
aNS2DrPQD2g+lZ0nR8wRfHpLjsuYt1f3AnVwGxFhq0EkKlJEzP2ZaeHbhUsxQ0ij
vtP8Ei+M8p991YZPfYOALDwgVsbX3ESxjzuObI0IahFcw7pTUOGyBBnCnETRTK0r
jjPNBgSZ92dfg1trsr0/joycSicIRUIxS9F+wUHzeGWfC+C12sTLyLQEhQqBJYzd
9AaS8vV10TSFqrht8tZ2aCEYDPz/14dVDRtDUjqFRnLwsJ42rCIqz8yzIOPEYtk4
G2Y45aO3zTy9HNsfWSDIKdiZIunKdZeyTiNU0n32+00KOEhcVfK7rnrZDgVhezBL
KnTEjGwj6u+QsKSkJnTJqQzuS+ahGlNwpmBsDkbxixKGvWKvOkWK8LtBNqTUdfBV
3R/BWZwbK9pr4i5WQPAiuqhV6uqSCdlb6Ar1/8CuVeWyh6F/1AXj5eNcCcILygJL
GgC2k157MFdmuWfYwC5xJm4fM16VMNK/DcCwkEAiNtD7E2rPJ8lFtRJ0K+Eg5Rf9
ot5pTK9D6EiSMSCPxI9uNQJWluPGL1UA3L46mv9+nFXFgxWtfCKxhCnLuGsTAEli
ke7ZM+Tf1ZyoG9o+sW3nDIn3ONup7oHyx9qtdaHzO7yJUEiLxML31/6GJ9nOgmZB
WVyrYe+qfH5NpcUoGzdQ6dhIwcEHK/X0RY3hoTtxPYQxWHmo5C7ZqS4kHxA+nyo2
8cjRsCKXIxefdGXROXnRyeVM4+t7G70gWmEacswkAqkiIf+IZdNO7XxANWjwY+u/
dv6amQ3IhgovdkPC03Jw2tG+E3p9Hm6sjLpraRo3mLsIfb/LgPTZEpIUBlxlWpfg
Oz23S3zPu+ibXD3hHeENrsTIjfdNdxwDdtpnjUh8OIdYUIJo9Goj8f+A8Wvnckbw
WemaEVhy1jdOww7LDDQpkZ1tqTw+mzmiJgGeI2qwRD/K/YM7ctQ5mjU8YF3Sdnlp
3kkkVKh/R+ABXHmtoWQ8hkSS4amIIwx1yX/VNqL/HCxIeGHHLOEmJuU6pGq/2Mbs
WWWUYbiBcMn0UzaMqjjm1CpfLQgIoD7pcgg/cPB4vTnl+D4neIkwPdq9ksIIX1YQ
A1dH3OgHK46Kyg18IBibFLl2LaV5JawyyBCNegqQXiMS5vqNFw4oNItyKy1/Z9c6
v8b20ofGvzLCfQBcp0pSz3yZd7Fyya3hGFscNyl9aGp9O4a3DNDwTFOhoa/3ntdR
s3O8wckTAh1rdYSc0LDKx4MdUeT82PrcQuR8rOBAj5TrPTfGNz3BTOaUvs0qS3Wf
2Bp8a4ewKOpKMCvuYdKErWngjAql704979NIXSlUoB5UxVxgus5JP3iSenSC6gvH
yQWIEfCHCZb7mcE/iZHqEMU867d5/bZWlO0McucX1iqg/sKUNZMgQ1k4kcb8adY0
+HpYUye3GBXVgA8UC2FPzqcIxlsXXaNstsTKqcll3FZt5SoopqnMDIvfUH6HM/Hw
kd81o2o2rxo9qvjUr3mrZmSU5C7ynIKFU97cY+g1URaet4iJUza78j3fQwil6UG5
YvQe8mCHh5b0KF6ZUAp1mPixCv4dPAEM9KJcFbNWVumwrSdnHImGXQ0wcoLTmmOM
XAl2wc1QkN3V8ekVkS3EOcDm+do81hTXhHhzNrBXRqozGyUEl6M8zJ4rVnWJrfET
JyXemdKipCzCXQghEESS2UwC4Zd0En5//TlOYVMQSctr4hzSafq4LunqAj7BFsTu
TtmNwcYtp6YFDT3WMWLHS57iY55+2qFNEW8WIj7SqJThgwk4NwPBOLHW4H0fJnIx
RQKWYBXFVE7YN6WV4xmjLzNcoEzwsfGyHm1mQcavdROy9ubFuSDvdBGjDBnLShvn
jmPoB0cSNBwZcIDk8lbsn2o6crd72RSqw5gJ+/NXmptGrjWqAzfPSREX8+vmDOlq
566yB+7PMblIGBkxecVJZA9OmrwYjHEObZP8cBDGMGztpxfjPSduIyAbos95+hiP
9KoFIm+blwWtxdCRUXauFNsxkOTjlCXMcOGFQZR9UXUm3ssW/I+ZyiTs5SxTjfAQ
8I40Cb/DDNAEiwcbXkyzWPlutIrX9CePnmtYFu2m9LKR8WpsUn1TUsKrpy/r2jj1
Kjbfl7yPK8KxztLu+n3pnse/lTKPbG1N4n/lNWCr/MtDhhM+zaeTlRZXpWih/IGR
yFdJj3xb+h/YWvOoa27d7WcqVMHiM5qKZ5D160GUsOAF7Ui5+/ixM+MEUD5aV+pP
wANewTB8TaAFecpz0B07G9l8h9vpqSNXbsDgaHvQFPemR3PZnMxuPM6HAV+crQIs
gLfuThHARSZ+C83VWS0yAGpuvjWAWhJxOxJf+ksRPd0XpD7rsVZ2K/2AYUKQzXU6
vGw2KZmxfkwy3ibqstUjFnTugLds9vr+11ytVaZ7u5wkGXRCl1uKeJVkTilPmLYh
RQDrwxaRJlTYu7ylSjmTUMqZEgevuvWpXuddt3MYOlscY7RIi7VMZHBJtPQ+rz0u
tqrVSOhlSiIWPQ+g1ftPUxXMRaRgoJ2MaTnFJ141wUDt1jX7iNW1oyqM1wwR+d79
wfiU/wfofZgHCdFFan4Pp3q190kmkiY5tNjyL0410GkUqqzza+VufkJ/0p8AXZMv
Od7ZHyKJYRRF3kEIKI/Oc3iMsOqNFKHmmOdomOeLsy0vexJaAxRkBBb8Q9p4q5xw
GtAAMJpqB0UgB7o5gep19VuDJui0OKrng3gfrz+5F0OOZ4zPCR9GlUXhzNd4zmaR
8iRujjBiCLblF+UpUCfIZzx3wjMNiM1ciJjhmxK1cJKjiRwOb6sEFKESawnAoZQG
XwYM8PIqK21QhhhxsRYQ7svlmuWQr6VXSJNmjlxTM44KpgLPGuSiA3gPh6DKdsrC
xStHVHUVUTdsHhEPEfhWPiFzDCHffvibxdmLl386O8HVt7mdQRMxbb/tIK+tt9K4
XtDhTXvvCvps2L633fdW1yeLCtAfyrvLyUfKGG1F7BgnmJuoIfHzwAvgFcaR5Z7+
o2KBfYVY4KSte4JRYHzYgEQNy0Eh+u9GFrtupQfj6ZycQqk/lWZ6xEKZ+/Mfwlt0
N7bc3f6AdAVN9STCy6Jracb2bii5aE/2FtYjurrOPYIu4HQyS/sNv4lMKrOnDghq
78Srugd58frUwqEg/H+2LpsucTX3COrfnD6in89GclzeYK5JORmmCx/eWZhShQ1B
FJmP3bGkM948MRqeBhm68tnYpsSqogsS3I6LoH8qxkirzfyZZKpAfvMs6r2+8EQG
jI9RjiGuzwqrLPqD63Q6g+Fw24HpEMxncuU1XO+E+xPX3YWWPeI4IukJSX6UXFVa
Aq6rLMst+d/JCG8kveg1LKQAtcRcR+aQjUL6QXXA4CB8xu+bWB3FoSaOSaiq9n6V
B7LKTsOfM8svtUnRO3HNANtbFBRq38lWHzSd0Hus7z11HY11mWvynBcRt5bQvpMS
pCGYg7TiUcLMtD5Kt7zLyggUT3mfF353TefJpQDbF88i7snFkItjl1KfCKYObLhq
KDAtH10/ZUY7WdD+B1gx3iSI8KdRTM4IZOWLWZJ85mRPvbUoOjKbW8Z97xbjEDE0
Ckp4ZgYri26HZupQBzcXaX1B/HdJDLhv4q8eBrj0sOeqj59QPPykDt58OG5eukZ9
JK3owHklwiCQBmh1DJKXJcpFryLA2Wpir4J3uzEWFnb9XMJT5fdEDJ+4V6wJf6Lj
xSw7PVzAue/B/CqDXoxTmr0tyqB7HiAjiZJdOqGn8TdO7xkYNsmIstFm/BuIxiZV
q2CychgJ2G99KnKSjJ2Rc3kZkj3E/Her+YDRfpl1O+Eqd5pQ4ryigkAgz/tw7gnI
AMPXHtcV5hjo9ChL3VQrmRhgZbkb9aC6UMbjBtF7yzFEC61y/ItlOl9W4pq64i6i
i/OevZr1VoD2fUygMxhAewX0AzVzV1rjvKKOo5MnSEqe7rhMF2bkW9HsbnWg0idl
rcGatX5jZ3908afcqOMcq5tfQI3UH9EU/LJUSkK2f/YktYEy8BXJUXFGZFw9bcJ/
7S+En+n1R5mbeaHB6F9kmooRKiD513rRNflsApaApEVnD06qyLcR1JQW6Sk5VBpL
DYJXpzzViSCSwCfo8eaMs6lkXCX/SZqmu4iEM+LiQdLPBCoznuVcyJba3Bedwk90
DmttB0PUvB24xFhQBCN8/vFVnFbMGaJ5BM0G9Bvv5y7VwKblAGTFW8IM1lr0IISJ
RTPLmQXeEFWHKt4MJ0gF68yldHVlSMJqVwWm7Pf9tdNAhp4KiHfugyTzWPkJN5IE
MRIXL73cBxwQkPboPY2f9w/5z3mG15/61X7If3gQJeD5ibV+OEGdey1xAFoJEDtu
/XmxH3EKnqRx6YzA0ih0VETA8JFPXXzlY8NzIOaWm7Yohcvk1Yn4fFQ3qSrllvsd
fDtOyJlFDx6b7BJrO05jhQ+Jh3Q5Lc5pJ28JO4qWP6G86gimxBWNW41srMGSnCWr
PZxVlUBw9nN/tbG//ZLYOFnWShxRn++/+hc6GUDCIcGkaJXEb07mMMtlAlbFm6Zk
Bi48ZyI1ZaMKbL/RRBwnVdmwJAb+Jw9O3MX45PqI4P5rgFW0B2yv2VE4YJl3CwxH
6Eeu7GpSGfcxAx16aPQU5W3Lr5alYF8TY+mVrwQ+Lgcl4KVdEzAWxaV1ntZIjoxI
ocGAaZy29IwgDK2O5NqxKES7NT7x0XT+ld5Y8VJTet2vmWl5/Ul+dpE1mivUuFfT
4CD58pqGjGFYl6p4U4aPQSexIru+9avfGI4uOuVHJP5ArPOSczKIZYp5qd7bvsR+
WKZzooE73t//T7x4XISyegTgmH9u2xzhJgZwWkyGrQVJnjPHrzDZeXvJJUJKsw7s
2h+AOE1pM3+2d+228B4J6UpA1G+yedl6LtvdhXkTrkZQ8tl1HcELjouVI8ns5Tc9
5sge5lKDUYDJJQ5Uc9DakK8VhGVdxsolXx0sV0+UGxIfRvAylBHbneMotdCpnf3T
Wa8+IOAvMRGEKpy7XwLJYJPv6mPjdW521BtvMUWgnH1b3s2nGQ+sBio2kOGqgHKs
4I5YBtPtQIMqJfHCvpLIAg3cofshxBxCcmQ3b2oZGqnt5Ypqv/Xdjo53hjgwMK4K
Ow6qNOYKd7CdF/qti4rMFl+K7Bu6GjVi3huP6Gv+OwBbNN3LOJIfEKO1Y9EKhlTQ
mdnFJmnjtfMAUGgmwcaJj24UdPPPvavK+7UD36t6CkoQY1crU7KVlBufzeojd7kB
gwC48GXVe9MIWwR+4FP4NdR0E6/6oDD2cPM6whAZ/TDh12VpUyPbLzDUtbLA4Ku9
UzjgxWyYSiQwiyjjCEhJSdMoW4kd6w993XpJiMUqrYlMhtpeyIyoQNTkQjXSK/v1
psjO8OnDLy/HSVxmDGUK5mmF3hFnyaB56XmhnZ0EZTJXTxo44flsbSrLpvOa+MF0
o4BJDOE1ANHMi/LmdjWpTutu2Ubqa0ALBeINChMcR/M5PA8BqT7lmsCnTCyNTKB2
bwCgos+x8eFiANlH2biC+fe4sBcuVYjbwhz/dQx8mKXHcL3JyHg151p8xgVVDUJ/
96hf5wzit9YrQlnPQQMXDydKqxH61x23O2nQQeP2XQv10DLMPNfYvcVM8aiw13Pp
eFIPym4eUI3ZRwqSPF1fcHkB23Rh31TAcFfPCw8bVgR56SfezFnAbBvylix9Va7M
pjNHyaIPx2bFyD9fTBh8QnzKk5udmX1RwlE7f+4Wj9yVSA7o1E7iizJ+TSQn4Pri
aJR5p9hze4c50wtc7IAB04SU38PsPULwRUUMDt6/QpgHD4M2Kkeaxx3f0vI69TSj
3x1aKxX7AXpzYgMH4CC7NXUEx8ZLJU9wy+mjhy0oSansRxt87cZfGEW5mrIuEy3h
wg94K9bWe0fGj+XF44mq5t0tei2s74k8+LaDYB556DPgbA2PMpfd3nbzH1kE6xOQ
/mpDKoXR+SIYZhyXPbdLBhhu5jJcBAkegnjduZJz6whCjz/x5QOYybhAlz9tLKQk
+/qQGnhuxWT+MQSSWgNtpJmehTcnuIRlGN8CeWvxoob3DR8SSRYF2ul1WT6/eJol
y2A1R0wClbQk4+zlK5doxKHJsscqHuzchlQST3qBZEBAZ0/3/cVlDAHvIwEHTykA
N0pBCmm6FLpBTkRMAIoQZOuZcfl1tUU9D7GRZGT5akQjpsUlQZKaPdisl3UXIeTp
//mBw4jfpsIt9Ut5FYIo6GIiQbsJflDVnbnTRzUmzP5gSAwlTgPUbhS12d4l2932
jJkV0BwI6/IMmv95ya1itcCFNKcULjIZjVSa6IrEEtfJEaihuQuHiOpvqPLGEgfI
3bY17DHD0mJc2XrYRCunHHKaRK8q1pt2OB/GSF/rUuGMd8cRSXG8O1BJmbC5aIXo
2LXHeYcoWQV0A2al4kHfW5jfMjg2+rIS+dwRdDxPQECdn55TvGgZsuaCpBYBEE/J
x1uegypxyFnlEWFV9PfRaw0bpA6j5T4MtUOfvtxJhJ/kIGdlb+pXbmCVYnlsmgLc
ibdCCqUHq6yHZM7pwKv/lcc9EuVF5Xw5ogyILlG+sH9BTzYF7jzI+Ri+xAwQjB4c
xm+rtNIN9Gkg611lmRP8sIATMXCgO28Ak8QkOK0r5lhnzc50WGXSBpLsbf1aQJFU
1lK4tUmJGBR2HCsYGRIZ+/L8pLa75vi8yMXvFG+yUU1qTg3Rft6K5MrMKl8QPoQW
qLbS0C716kb7vdOGvdLBIWz/MKBJ+jAg2zuVDvLQWc6Zc4hV6HALed2MjwV6N5jY
kXkIz21we/NMEQiq5VAvYL4jifJrsjWuEJtKtL73j+7AE8mHeHFLExcEj2xD3y/g
7PCewz7d//C/PKeFKgwzSzyle31jPgiufQettw1h1UVOoIqmu0/Fnbu1EBWDVOAi
DZAke6cDMmNXpCpOAUg53E8PK7XSDLANEuOfzJsmAkHH2q0JIhk+aSwr/TzjcYWo
muPyfIsgtPiS1wtqsz4jPPaKWzWnHxuNZH/eM3N+V9EyEIjLXXntb4E68oRLcExz
XEvL5usel2AgZ81c1JYC1jSMo4cj4kbrzE+Xl7j6IwV/EMgYD4OJkqIXgIqWnld1
24Hi5KJ0WMaRGG455t9xSqQRgjoVn+iCehFwKfqJ4ATGFNl8LunNZulD5CV2pmWn
KhUuoYA5lcQkpsoL7z0sRYxqYeX0UzPpZPLa81GE2ylch0alEjvyRRq8SVNK6lvt
FaUIGR9Npe7e3DsK+AurTIzoiLy+80McI3/d41AbGu0SW+j8c9oInWLiw9X41Ark
z52iGpjlJswXRiUCdAlHS7SYcn1el0D7cdSZUhbH3ZCc/16llNiUWSA3zzDjJ+g0
MoK1xl4XAikuW4+HqpdcprOqkMmehg/rgujDgUVHxsinw13vjOxaKqxjJ9gp8Ke0
HQXr1EqHUmX+yiUzGXd9aRJlahmYvSwLUh6k8+K/XnGiMD+h6IaC+QcAaI+JCIDt
5VnY5Om/NaSHio1FVfZx8D85o0iFLrnBeBkyUJIgaztaGq51G2nOPYPUTZ/hKX1D
KEyF3e5oCgYkMFukeJnxxiTsfJKls9U3z6FO6WI/8AbZaCzt2OS7GW2h5cEKBgnE
7Z5/AmDcMsGHI1LJX+gkigjQAvxYZaoOafyj5aG36o4Axj6V2LMDXLnEDoNrkIbh
1n/vAAeT4cqVOO1Idj7PvK5FPtVdz4Ad72aVH6knwnbgIRLZo0yonbDUrwq2Bg2l
XSuWHKo5XnXn414jmjtH8wqrZ1WRJxy0jyDMpSFd3NnGnyT42Jh6RtjFVhYrhfC3
6ncu/CHJq0+rmJIrqBNF8Tfl/8ZfFvw8hgUKGl0ql+fIojC6EScwBR7vTn1K8Dux
+95crdaNZ3LjBvb+CKEPrgdYb1uNq0QvEd6xQ0Uckl6a+y1HqEtuHsg/Q02bKiux
fCQ6QkoAWTquxmXDgnOBGSy8kVFnpneFuKTDPCxtgHEEqQ00G7O1zqp/dW9mjvEr
vVBPSOVswNbg6nWYsDDsLgD6CW0ft6mUudQiTWck/NhkqaZ6MWDWZR3WrOK+7x9L
lV/C3/D5ASh6jKTEVEbZuRX2oSfgWev876WbV6n+AB5Emwu6Ev+USxADbeohITj/
2SdlgsesE2RYJOvyjZXUViIoZi0REVTSO1aXqvVixYu0yt59WpxrEntXc8G45l/j
1ED5lbMXf0lVoEvp5nwRnqfn7kxNMsS0TjEbx6zdeGxrcHYjYOVO1KWw6QQX24QG
Hlf8G3k8uDsnBqPsgUGQ/T0H8jpDT8YTZ+bn6azhEOj+pY/j3yPww2PAlw89jAad
vQYPhUqYduBuYUvvNtWyM2AVJ7c/+nWNkQ6gnE0xCVXvOdUmptbspnAc88nRyS96
5klQCNuliKlZ0OO0ZioxMlBveXteu0BfKYn99A+n30Aix9Rh/+MaTo3K4eBGt2Ko
YfRMtQjqLR+k6AujgWIOlV2HRF+cIw7rVWAADYzbKbjIO86xHoU8WY4ok00hS6Sy
2jz3R+wwA/fKLreEQLCGHMm5HOPtrQakhNoBc/dr+byU1i9/9HVlqnu2i0WfQY6C
0nbUjBgF/DgjzFtwdJWKgDkuzn98RDy+6FnGZRgDYM+OhjsvjEDiGpF5J/FPEKwd
Lx2QXPSc2Mum1HjZhmXgYjZpZHP7ErLDnTaxlu5mcrxJYvhyssXjH4nU8zR2/12o
x2Q+LTPfFkZnff2EMawbc+ZoXvv6pSwOttOn6NXIu3zSVtv2js2/NVHXIrLtAdCg
FPgjXDqp7LssaaooKGfGdq8pF6DBXd1NzCO9bXE2+QdgHFJSVf7/cl2+HjHko8Wm
n6nTCFQx848djUDAO0mxS91TJ5bc+/hYFWwB/X1SxUDeQnTZNegBKila4d1XIhxL
XdvqtZyq6dDXk09cwvt8HZqGm2dwF5XkkV+Qh0l+RvE10ZKX1vv9q/YkOYgM2bBn
0ZECC8lGe0Q0UYXxhbaoLJVZzdvdjI0olYHw0pppHzZCONEgWAceXJEapPJrXCDp
BFgkQHCMGN+tP0tI0G6j6LGW+AKkJ9qpCemC0nJy8tjE6YH33mkj0a9wXu0kODZV
3zQw0O+pRDx9J/x2X/pH1tDeQyS6fz07Mf5f3dVSAKW5iFWzhUUe317ICZAmTf/R
r/7BVGN7PX7IVehuNymNQ9C4wOvpN5+TPVy30f8JcL/avrDVxundq9U/ob3AlNyG
jiKYh5G2MjAYLGovOlLhdyHXWcby8rIj/fwSfU3rHa2N/bWBoD4A83GZRxFoWLpy
OUYRDZwve75HQyWWX9JDSzporuTd/nKyndOobn7FMGfES8HBk2GDAngqTUgLhiPh
szUEFBJQTV9fpU6mF8dzt1vBEor8cEo9x+oVgelDIrKIi2Anmsl2Qecsl8Px/zEJ
aYPlfQFh79x9O13VLz0XDaEQ9JsMqe7FjrqKPN4zr9FyFiWwjlqsK9p9++wA7ufF
P6yO9PAXJDS58HCxr0jDbjBb5wAQn7YvZ7ZJjTcRiRa7g6/vG22reGjdFuwBlZAr
JNPo5RW6KFhmwKM0A+TZHNldwhj7QaEcF0GKbuzslVGssudb3m5DVcafROrFksXe
8kQxNc+s/AP2xZ3vwpMdOC67zmgYy/XPowl3Ftfw6lSj6jDZ+b0ZSgDw2IoB9Lkx
UBQ+HIqH4Jha4g7wOepI9x5Ma9hgaCMfny5440uDXmPFc71Al33JdmMDf3aTtTwd
7HDCCoEoPwxELcREkY+SEnOhNbK5GuTq1JAzDE53PKMFKILt8twQWMVf9JNE58Qk
+esiEl89N1vSi6/meUj+DWxYh6z7Fe8rFMHInxYQX/4MjUtYWixccotogtZGYgeh
WEVyzwn/LfGc0wdRCG2mHEHXdo8v9IuYjEdIUd1qrtMK7WUr6sL0Pn/aGLhV9LpJ
Jy+n6iMwTxUtHh3DUweLI6qfz6W+ho3TEoXWGKEoemWx71/QXKHgCOsiKvoCjZI3
/8qn0ZqZJhpBiGjz/8JNUTUbdcqMl/h3jFbaYd/QPiqgzoDwn1UnWO7rUngjpy70
tJNR2iwvku35YCiS2boHXMXDGOchVBeIokPMD5aDxhjU+mV0Fb5JSK9Mh7pNAg/S
nv2DpoFVo4tZ1el7NDjOhVJ4bPyaS4GRcf6bS4wsc4y8bTpMZcal8WRXMaCUjNhG
/njxsxKFWcDgvKUvQKios8tjnOepqjvZfaC0puV35lKsogP0wpYp/16QP0F99QYk
Ev5eQiwTXugMwig7mXCxEqIVJZlfNdT4kR1faUOvZaIl7Fr+uO7WoXO/u5tW8WD1
XJAfGZL9phy8LP1315AVPZ7VaOUpzM1rWEOjYn9jylPoIkFLlr9JvhAFXtaxF4pN
d2lCkKXNK3ZS1ZtvcZBcIWBdVgtOvCrBZi1Eecnw3xrrIS2Nfoq5+eKFbOiz0FoZ
Jm0ctvnMHEN0SaquRdg2HG4b2CSiKZwfvHQExFT4T7Qa1f8lHVRJ45fqgnH25HAJ
2hnQpDTJbumgXJuUpR0vgQUGL2a0h/eTD4PhS8sXypmao9GAA5eRQwL8LX3Vwsme
0xyNxcBMShtJVLKGuoIjNMGDHFhsBCb0VfthR90z0j7bjQlDziOaB/lFMLha9VCy
kL4b1Fi4GWHGFNQ8R3ws2/ZP5CGZIqvh55z4BqmPrHp/YEB/Shmq0Xz0lum/blpc
sT0/mYM8ggtl0pzSCQD1wDQPFWUngYiicEY7icAm4QY6wnI5IxBCnncIDq0oshXw
VyvtlMc+LWiOckB5rJ9mo/+N6jYB1myQQaETTGRIq7sj6UriGQqaW273uxIBMcav
x8kmiH68ksNzLI4ysIxuCjwm1xhSWfcqwgls8aORn+ixX+Q8SIJzhVg8EYNl565+
eHT8rPf6s6r995rUnBtedeCc2d0PmIbJqQOhQbNCT4nRIdKudDjSETvfRiYcUSaG
+uYx1IhAdfIeko1iB7/FcvO3QoiyNzuB0H+0PZ0Wa5la6gLoH8RL1R31xW2ziK2g
dJndaZR9sWLOUJ3IEaboDHZ999UuEN9dtD6HOUoB5DmEz2TvFeOTZMV12I7ht5nI
VZfJNaIhK1rJsDfM3FnHVzmDZSUxFHqHD/RUtTXZsncSXvFKN4T1IkOsyywFnmKC
OOyNIjSdL4CfJMgxABtWfe9lC5KbuSTUrNFgsHLUMCt2kHOVfIpROQ10fkCDLQDZ
lXmXMSUrdZZZCmJTwgVNmluS7+Y9e3j8bi3x7yNKlGfrRI8tJ/bnVFIYSP8rnyh2
wre7362722NOMz7Dm5EudFmqyIJZxis9TnSAb/35/6lKyk3wEElTALwPXqfPaeF7
ctQWHURrIsBN+EEDzl8+aB9wRzG5OpCC2uxyVWr9T2bD77KPm6qRFCpVoZ4A39TI
UQMRFQuvfR9s9jA9GFh+6BMStr9bXoiAVNdCYqkdRUbbwfbVtJSu4Dsa5Yrp6BKj
mwfz6FQ2+ljI+RFEcYVaCL0x76K1LE8dZs9wnZHdHtYb1vYBh8B42KtSrOjAQTA+
sdF8hkIZg55btzKEtLIWwQAsBwUMk2xx4DVpE99IvmbVcvSx48hAQmpmBy24UK6r
K9a7CAvO0xTgaaAghZzmTp/ytZ6ufkNi72LBK9QqJUfeuOcw3jKzMaf3lnmIHpel
Iqm659Qja1cajYDXij/at3ONN4lKJoj6KTzP0H8AF45WNSAt5aAv1gxYPnGNlv0Y
z2rRHGAZcws7VWo1/oil89MzUMSUE7aZxvHyYAkg6A86yJmjAN74Sl+nKFac+lk0
aYBxyL7LNKKKNYfiOkiYIEnpm2rI2KKz+115ld/mA/WeL1bQGu0VUBN0mDtc0u6n
QCsnlraPpypHHpFLcz5hWJP/+peQ3B3nt+rOv3+DY78gc2A1If9QOwJksL0OsNQW
ICo6ooFAwUBeDi+bMxF7BM4cTuNGm/OGQSoBGlaearcikd1mVLo18Og4pDLvKDif
ppl6iOq32yJRjqf6AjePztmlFjHq96nA5Gk25AdR+1lf4dNZjNMxqWLGu/p9mpXr
pNLFFdXxut5pn+WATxyv2PDXAy93JOM9vLXt+H6DxwBWVBSqxFT2yzLCR0wZLbrV
eEyIfYLoMVNz6QmOiJFG3iB5hz+bTrY3403uv3/tGY6qtpZcbvoFt0nf9C+/zEFb
KOrp/Q6gIwwoDJexBZtx9rteMmBhNgXYs6OoKc9azsa1gzB9JtmptyuO4l0/tOzA
NrZ24uP43GG7OyDR+FqH8uCrvjI5Q8NmtJwi9neGDc99BwmlWEC0NAvswQ6eXAW/
DT9ISLBm5e52QakljlKiGUV0jSFHaxZK8mYMFL6kpVrJZCSOdqwyyD1V2o57lz/y
kVQMA4kOBIRiZrPGYu/Ipt9TEizhZD7qcNYdBaRtgCJZLJotTQ9ZJ14GkODB+Z85
RdFFHRPb+sIgBaD1BR0kPfCKeuXyDnGBx+isVVuww+Rsr86ivylWqaoR2R6d23eP
QXDGywoitDqtB/3b6dsQFe/0pPEDEtk+yWAycqg9mcExhRup+bnb7bCMj9hZgr3g
xCFfB534DfE7fL7MM3QM/44XC9CZwKkFIEB8lrgdTK9cEPhv4oP+v6XLgRDt1mku
od36FNrBh5wGJDYfPV1iXzFbUYvCO60ZZkLE4RcMcj+Qk2qYHChiWMDNcQ7dnRye
weOBHMvFwaeGVhQwAc3O9yyBHNpwb6YfM5Jgo+VAh+u3cgRfDCbpF53Zcr8szSe6
bvJWx8Qt/AHT37gI5Uq5N5MkV/BniyCcEyLOfw5hZj3FbgxBaGjGvp2KFojcB88x
9yNh4YoD5EQ7iW168g5pcXLbiIdKy6Ii7DLblaqW/rKE9KlNk4FmDb9Y2KxVea2l
cGtp73qxAN7Nh8aec+wqyXx1KupBjczY6D1w/byYXd11KOKlEb8nWx9jbFmPmaT9
tKQy5ZSLB51uEvXfwO4wO7F/DJOZy7BE7NK/sNc53TMuBhh8xhNmeck1zYYKsiQg
3ap0DLhWataZ5ec/GIAEDH2DyiIPfqsVeAYHUQHf8phz34o17JrFv9yFiLDp3gbS
Eo/46eEsGntmdsgtOTFYgspoNvn1mFY9ZtjFfRvJqJ1JItp4M7p0H3PURER6dFKW
gNQ07aUp3pgjj/vkBJ3NaQHEy19ny4rjSvSx46E2VZ2igKvFjq06jPHuLindVwFm
uL8bmgBnlR9ZBL/YLp98iBzwPxN0UssC/YA0Nza54Xx1KcCQglmGccTHQL+Ehy3G
UC9ph763cNlip+W4X7u9Rcwt+CzVUQIviH7nX+AtQmKhKaOn+TjDISmvpv4RU+/F
K/dvAK4o6nINl2ha7bqd6UxLNfVIEUDottz2Gjr99be7FHOLY44L1B8WLiN/nwqB
bDLxpGS7HfCtFId1M4DzxvJK5C+Hm07en7TJNEi2J2ADnCAhCZDpw3208BO+O8wf
tSGa8DMky3KiAClq6dmQ/EvrnOwidHZ/wTMWlDqHuj4/ZwWfBxbJP3QluHMsaQhs
XO0zC/7nqLEBaAtnTK+SOXQFN3Jn902zfB2ZAgWZzZLv8MqJXMdAGFjAp13EJ90b
Z8ybyJeRnirfxi2k5BXaoUbaqpYdOiu+w6TNTCWwBnhp5NIPvfMljDtYRoPxW00v
GZUK3NiVponFJmLpxkowKHNAQz4yMvvuAxbQFhm4/6I50X8YAwn2gkPISqQEFq+5
ScSo44QnevD9mqgJDQEcRo43wFA+Dm3N5RRMkd1i4tIX2yh7AHEat5cYHuiJezsa
M6N1c+lTG7qGbBK9ynWH1fI1LF9xN4x9zCEPFmzZnis6+D0qdofk6oSPXg/f82dc
2JXErDFldLQ7wlRZ6a/RH7xbwm4vT46rrOFyifCaQ8r7wOkimVBCZ4Y40tx+KKqo
kHBtV+0X0JN9DUzkX39rq6hZ2K9Pe8r/EfxbvKN8z73yopwZ7n9HbIKBW5Z96du0
L7NZFfn17FJKwS6T/298+P9Y7tjJq1jm91HMxZAt4cP1lTuN2+GIrEdca7Sg/77c
EQzQRJm6+VdT7cGDo5aVt1B/Py9ovuQk7BoRBYvoSw/FpwHgKs+mEBFRSxGV4SDJ
lo5wV/+BBBGJ0wSL3J6jmk+ZgcxS0mVC6VB88uUt9TxQUrOHTrlxKNTkNxInOM+L
ZvXrT9qhCL3rOfN+ztl8SijNraIdXoWgtbJJDZKTY2+6DoO7X+bs7hROXI3Ahe8S
zuVXqNoLaSxjbwAUjR5VORPkp1TIn+f0hr6lLUBIkAgog7Je9PzU94bCaymXe69h
CaSRqLbOK6Y0Q/yl0FLd+NIaUnKBRDYk/KNGJvrkYu7hGABbzesBOscAAMbKo+6+
mQ4Z7vaLycA6jNXmfWY6RzgbWG6gjRSs1lwrJh0PF/UhyhzALUCq7ZzukIa4DFPb
Rem+Xwu8p7IumqQElZwdhnuKW63H3pntaVPIUAOKz1Gb5Rp3YOqOosLbR3iyFspo
4ycENmiWFCHzFomG+PGyMi+AWZLI144GbnN0IDba2CrRgN5wWtyeGm+CtHwk0Q9b
HOiWOHLfZWAGM0X8iLFiqAJJbhhTwfbEo5UAVqlOL7W9+LOVyOd6BXs+6oCRD640
8MzLE4miurLj5IHTEUugwT6JWvj5KViz8sEFpWAzfbxzB9QP3IPWkT/qEswcXeNm
MYMp9swFNlGJWQ5Siu4TxMiBU9xoCGpr6XC23dmoa7EK3Zmny/4SIFs9hM5bVK4p
DRE24WQCp4S8QHB/jPpWg+CIvwZfvkmbzZsiAsG7UkR+dsyfhKHN85PhDqc4IlbN
0AZFcCBJqkSoNFoI7DhfD9gwmM9PIwYTQZ3TCoDTguZs/NFYw0FNppPoBbYubWsZ
2Ff4APBgEjb9mFgFrpex1HvYa11KQrShOB2W/R6gYow2vXYpgumkMRbzHyQzwv27
f6Kxn9B/rbMJKvSx7hNrbCLg227bBw5fSgQlKjztxdT5KJAUGqQtxizqlccf/ylm
GLl0TLhaQ36FY1t9RxBIabebvl5VLuFx4NtkEmsFeWyWLi37mW34rQojpyiZu4aq
2ci0DVLzDJa+qyhb5yytOtetVKwiWsqD16AckDgOxVy/uTmw+a7wA0ZWsHjVEtuk
K+MokgbBSzqGwdPXB9WEiCmNNlzhqFytnO7bhkwWpQdmoeiltY912bLc8dEFdvyF
Ba6h7gKAj17+WaEaa6ZUpYcsx4k1GgXUeQcCfcd8/vC4ve783PXfIXZc7Brpyj7Q
7I2xGHSErE3H7Mb5uXlpyzJCTsRiN7LMJL7kDuAuPNNH2p32+YakY9yWh4jREult
Kf3KqIjHFTEJmfI2MJ2smAiTs1Zprc1YgAIKobp/GiI3h0loNL/GWDG1+kduqV9O
kB6eQ/3mcTkzCrUfcBywQ+xeNlgHM9DjaI8w1j4EjTlQBgchAP4zaLDYKFXHCHtS
AVeadbNKCbZndPUB1g2FI9SM3HXUg4CJV4aZHL2BJbxw58NPA3Oyt3+g6CPMxi8l
4O3noTme3zG8zovwdpOIJ/EWSOYDEZVn4/3KGF150TilCozgY3MM0whKAgl9VP8m
/I7lxa+aiXzzqjNcNKyMv9OvgoDb7/m3hPH8XzyweAmsU9Ji+Zwk8eyFDzmqYDk0
da6WlKgzkyoI5KkbilKXfWvUNl1zYPZji7ipYOdkuXO8xgL5HFGvjORwTfbT0s4a
SxnPJNlthPdslP5YhJn9is1omuDzV7E3u0kMAblcPBtaXNYPl9FDTM7Ml69y24Fc
4Znhzlsoc6qfuyo4lH7Z+ukIuAyXfsoBmCYVqWY7m3GrublTbqWhj7aPtFPRlXI3
tvwfwXympwM6l7eAgaE8PH2zWYbKhHKiaaJrMcwlZ7iWToXWe9IvCsPzyUC1vojJ
iLGaVZlCL2d7N1A8Mp4Sgl/1fUtGaOW4Oafq44KGUtJpdTKy07McgD7u7FbAsxIU
jrrt8aMHx3W10NzK+LDnOv/N9+OWQ4Rrgn0kNpkPbAfK2Kt+Vuu2ZODaRTyFSrWR
5a8PzXnA2eqYOqDc7Fu+AN/EY0PjGlXVEIGNd9xtW6gNEimxxsl10pJuxeDxRazV
3ovpKWj1UZCDCsz/Vpe+0Zv95uPjG/2JURsXzzahuuaWFR2LgWNAP/F7RGbivuIj
nZ8AXU5LJ6yPQCfpCA6PcRIODiw4Vd6LHnIroPsdDdBXww8lRml2Ney0ZCR6jR84
TQb3304/u1glSo7eQD8UW81fhu9ncvGtOIAzrD9z+ep+pQ03P7jq1K1LoJ5UIzLL
etM+ZI7OhD/rpLQSPxRtsEKqyOcZdV/LiK3+F+A1ZqPHdXFdUKHFkHS12EnxbsNZ
pcpA6+9mWHJU5f6oX/t71QLeOV2G9TddhmQSorSyFM5oZT8w/OeVQNeyu+mqBERX
yfqQEQarN9+5NwnuZtGqJcahl/N6DSTnRrU/dztjUY7QaHCL6Pdqkk9bGGV5FVhH
KVgSbkbnbkf8sgCIcuAEG+BGnnptmHkcLWIeQoUc+Qr7nwNny1OkHmC/jLnZs/Gz
qHWtblWC3Sc1gw1nvx6DCMJ6G5zq9UfNOyFJA+fESwUqSGesN0bHec5tOey9T5qC
4gTjZfSkHRAX5r/NDIEYc/bQTk3Zcd1V58+h29yrn3uAS0DaTjuzOaKZuCmLi0hC
1FjDfcxm3vN3pS/9QoEMaLW0LJIGgknOEtxx7D6KltkoBeZIHOjfcGyf5eOHfRkk
v37s2w0e12WrS0RyfZvJQn26Ll1xxTXUbsOAYTL7fvVuR57qb4JbUBYEbjrFKEAG
2mh+cj/v+W6x5Vc2f27ZObtA5Hu3svP/K250tu10qH6QJ7ESrEpCzmxkx6lTd6Cj
rhz06TFgRoxTl0FXLuCFOU/7Swu68fqYPz6qfGNgS+UI/S1WZnbtbNJlGTEqSL+b
GvF9tg1vYnfZDbKVkS3Jtc3hXR/tNzkUCmTb2tRhFbLWMOJEaWLlnn0WT34sHOOS
FGPNjWd9GSFPHE7hkpgQj9AJdl+wTYgMWjh0GIlmgYZwNz5XRi7i9xDSmZFHD3xQ
GBkfsISKKscEg7O5Gx1iXIfsBhkX9rt57HjFtQZf4154bedO43KcS2IXyZuYqG2g
BZG6/2isDvCLK4Ch2Q1eFT9kQcmDEuZ9Ih0UB3hbma+96y6HnV5MClOjlsuqBu2t
AsxguuCrLK/+EVe9MAAo930TG+kVhk7Hms+VVKa3cjWzduvPuABhoZHKig/wLtID
4jbjJy8+SzDZVGLkVq6Hxqh7nTwfTx8vpEc8ZHQY+pcR8scBA8AEx8YfgPThotpy
H6HFa+8EMQWOcxiiaa6pGRjWc/XI+Ew2AazwlFjAc2nL0khTznIsEFUuG9pVxN8I
fWqGdlFFtuj8DdcWEMoqcwV6/eEKHxt3G12T5ShU36CFXDDxmwJ+UX8wHgGhBbb4
AnxH29Q6Na4N6eBegKv6hYYsmWJS2MYJwxeLF/hLuU/cPFiPBH13PSdKtGfmotbg
1+HIAhHh/j0xEBmjF6sV0w1/+3f51r5mVbd5GwCrSJFa83q9adsTXuAqOox84MFS
4pVt35DP69UFb+CCZ5XcphbxgT0f7fOlLAk18hWXwENJCjN+HAN4j5mSD01F7spi
6cYhXLne516fFe5iPCy5vU07KXlQyincnTczqIXEFm+zD633EXwHTIlMSqic/35w
iIr3a+i9cqj9pUuNQKxhtzaO8A25XD9XcsxbqIQC0yqQiLN57EZo5AMmHPwPuMQP
ZoOM/ZUDVXInfo7Cd+2/pTirFyKGH0d6UeW8L5Mi8hvLbkFvVlmPUe1lypS4c7xV
stSljN2Ew0DK8+csvhvanxPZsmh8gyCo15yEd0YmnjG66UOBSs73wahWcOT17DVs
mHjYCbJDhPAZYybwdm3XZvUnoKtwUh1rS8jssZi3NJhg4EbGPCDzrp62Xo0Gaabe
OKrg3oaqQUrIKQmAyNW+KpyY1K2ixP5VGh9o24mSAkorHcSYKPFJ+IPg6Oz7wW8x
c7o4Icud1hcHKTZmGQAsuSGs96L5FFI6kBVaI5Ysf795obLqnvVS6rnMfkLA4wPV
QPKJ1CKAg7c7mwwK930KwkbTUHkoP8aXVl5TF7jpA+9i5kXLTjCW6Sz6ew6X/rwd
IvdWhUek++8lJpHw2FEaHkJ0TogGuvqmjw+xop/lYTchcwvRkU5G4B2UX6ZV9Fol
yyGa0gdjpSh/Vo28vFU8Mu4tcbFe8dOcAgMFh59yq9ik94AzKQRwzr78btU6zmNX
Wr7CrKyf5y/f/C51RxraDaiPY5+2Z2Q0joB9vCt+8YyKjYXTu3921EkL3p3fYkBR
L4/ogr3XB8FtKUsc9IRMFYljikD9rPKWkxXkKZmUk4e48FTpFpqsmCSefuVdGAAe
SS+Gae5FIF6aouLYZKWSZCoO42pax7OvCHdjhCX0f9JMqhtJbr4xXc6R8RJUHL6z
85HFqVDD8IOPNGVpvTge2quvxjKOS+4ima0aMxhT2je1yqojJKqginu5FHNYT5J+
reb96feYdXTRFi83NY+jw1dgDJVfhAwj5OsXK5qeQvOE5DdJTXVhvq2YSviRZks/
7nb0j+r+gwWpFSymBBGdpvqrgV6HyO3puOC8vzeL8cUTgeFvw3OnIGlAjX2+hk2Z
3pPlzT0e4KlGxIa/qIvak2ZvaWrYiVPAbOz7VV/ofnOoLkxejWWZLNGRoaUmqv1j
fQ7BZWIbToAZ9TwJ//OHXH35H7LM+pzJbAcsIKpA4fVqGK80FfCNjIvPTO+ctuHD
2VTrJLKj6pQtdPbBwyDITDR6hSjfb04cGV7q0fJ1W7NuzBWZs++YNKS9y6/eLoqp
Zi45wJLTCT/Sg/nkIzU2C/Y7PmuwqiXd4fVYB71icqs5rU41YUVXGmfdqbvV2vug
x47TOUtxcz4z9xIfNWIir356mepwWhSW95t1QY+RD9zQCJPzuO9pPbcQq20qbNGa
8kulFLQoCwyWo+mN3oTXL26XkYy8bGBFvPbNckZexWmxudG11LUZyzUndm++pfDB
d892p1Y46HLaS+sevP/ImTq4HHvTgpY3Z1LSq0ornLMgAF5pPlG7Q/2AW9qUhy+e
IhhBi54aqlh8GbeHT00KYZ4B/9pUZkTeUdngj9UShpBJoShBJPycH42Cn0HQWGTr
OTwagG+jwYfGI0T7Bbyo2pWZbfr873ghhubqPiAvHrQSav0Dtcqz44NiAlPFiCHp
Bl6zxF9b0PyZ4eIiKmBf84rHwf2HT5K3xz7hNw12XtZnCONv3oGeUCcYfNxVoLQO
w9mnnJmDItsbJ7uzMIEQn8UZCtG5vIHPd4oyU093Zw63UDEodbSNekYw1Zo+s3zP
sWV3mwT2tat9S2S6ljnCKXivYEc6zlUxQ0FZfqhyhziR46h3HCNWoRCmuAeFcehw
Uwe6ea4RXAFjyxA3FDq2MVnkuU4Nrc+mUbLdE4GjXu97SNrRMj2HjdQ9smBhvmFq
UNQuYxBGAfmGE4qp+pLgZV7HWcxwAtZ4kcQB4s2agtp9DhoUgTfCM0CJKNLpOcGA
JcSmrFb54G3KPmCwxlI4X0/r1ZZURx4TwiLStnms1JteGUW+5fVeK/jc+DfxkPR5
d49GXIDhAJXTCYdO5TB1HwHgzFtlQR6qAb9wacfqXzUrUtvAvlQ7T/NC6WQlgDUM
WTmT5odieYpoFlZT0Z9jwL5i+tmKnxiV6p+uNNtFzhsnp90vUkgxWM5euh+ui/Kq
GeaoYhplHMyhbE1wu15E6bxY7+JulNgZOC1naBjt+/X35FmzXbTDswY3knJwsBHh
7eVioFW9wDBwQMViaUk1kA+W2hr+MSZlQCaTUOtgCFaoBpTnYN9hjoMaPDFXtMMt
nk4K2Nnk3r1OBfEsZ4urPMVWJ/KyBatddxPaGt+kbQciFy4M+ksTkIEcT4ebjF7T
qoDb/BxfEfKjnD7Vl20Ph0PjftRlZqRkdgJqz3doeSX1oxy/g7UuvOSzRJB8uG4h
nPSJboXm5u0kyKAe3OCzYQEbvjydIzhhUcQjQjgwBPq7v32t/3CF1Gk4vlqNwr2R
cDDlFcNLousjyfL+yNvkA+zg4QxcEh99R6iBPSGW4v23yxhOfYWQ9Xi1c5IEc1lF
Xtm0gyQA/ai2hG8ImlgFgr4Q20t8Bjj56T6uhiJOUGl694nfuNreLMLq+UXyfwa2
PcOjnpZdVAxbLXHD46cakXug9veHbRrEVGmov4BVZkF2VQKU8TZdXO9EUY+qxTza
jD0qpUCNO9Aj0RTGhNfwLLqDt9/YXJdCcZUI7mkiKcyWjdAujHe/OyY0DZeccwKj
QlpdScOe7QaIq5KHCpMvnK2TuJX3SlpD6tjNaCBW/LVv5/E4kJVGXd3P1PuBSJhn
dknE04H6JKNmnBIOPanZYOajQIhaX7kanvDQL5DQGTfgMHR3XTkt2LRKY5VwiSsW
jrpPuxOEK4rUA6qQvWE0Vwf7o4GaldMNkCAQg60oMoE9ZD7KICYTf4vpN2kucZoZ
AtpxdbMtUtvtLHFprfZXRXwd/GtWIS5o2yeR5BXxzz5VP5cWMtb5aRtURt7E600E
rywxobA+yJ1vWrdusUbUTRmKYie7kivlZvXvxmm7A85zBas3nCWvRhq/GVjTQ9Cf
pZOAsmBSr51FSWyOybDDkaDvTG38VHxGVJ/45ShMGbU95N/sFSEh6Wxl18ZwI0Pn
JjK4kExur7yRxnxo1RNjUW5zXzkTAiNNBLKneK3LfzlWdSjVzO8/5Lm4YrRLX/ut
1PSkgRPYsHLFuBS0mfSdu0F4kBof29zELIauZsRkwg5UFOjRXcu000uCvOW7Urm0
Hs4oOuQ/0LiSMyLuJHcyJbSQhf2aXizuMGGv1+hV2NO+zyujkI013YGU1R8V+OWS
b/ozFXXI0RovsV85K26mR94MwlDuOHxR3ta0cM9frcrfwLlCCjPg17mzNLL1rKM7
HP4JWH6C9gA3aAfGvUHFNIodh5ROe2ggvQLfPNiY5i1u2Z0xJbQ2kTVUJl6dfSDW
EiiQpk3NSenslLQgWQAZnDdeGGPkU2gX0TfWXhaYdTIt2PpVylZPczj2E+LIWC9V
+0GsRduR7Zig58MWxUkETBxndBoVd9TZI7NGL9Jl2r/lzjWrfLvCVktKwLA1Lqvd
tWZXj1dXXKamE9d+4Jd2pn4DBcLoSv8mZxCb6MZklb3aPkH3XYUYNgNx7BVOXlDH
sruD9ThPcb9KZWTwoz1thd/D4Wf0mYwzIldW+eTnFx8as4CCqIgfmu+fMnjeR9QP
Q+23lnydElX5kx+C55B+BMNuKMR6z7ApOegESI5R7A60RUZaYaxKJuTlmvh/Wl5F
SMPjybg9n6RKJmdNiyMp9pu6ZmZYJfft1KI7LHIlQ8/Gx5OY/QMHLElIsa8OpOx2
MVOwmFBxhxw4RLjMAxYhX9YbVFy20mEoqp0dQAPPCSdG+53Sa8hnNYr7bLSITtL5
pVUdyup4Vr5Ekqhe/wQueUVeZ1eMkNb0u7xMK2FQb44wcuj0N+cWrk2Mtlt1DLbg
vxLAsyCUz8iFRhJ0HAxJ20/tzx+iIohVsFMIVnn5DsUrfi38OMxcYuxvYEW7XpRE
Y01bSKsBQpEWd5dgmpI/BsjRa3nlyfmoeavovftStQOD6KEwINVYmRT9pMH7+P/8
arlMlBLFpTkbI1Xjo4+8rrHFJdzW1DN2bvXZnbjuBOZXm8u5z/mccz0KZ8mAave+
EtRkFDTYStQLSz42u7hR2BvAYMUuCpLaPpWs2pxA4bUe5uZdI4zNlDrQdLueh8KE
Y2KB4TCcDP5EjpFyIZKnR5c+ne0ni3Q0ALZmJimoqGjSxqWOqy7c8bpmm5vRGZcZ
3Lfi3DiHCozuGYG+utcboH8ax+gfhdw+bmUe0LtC6RXvVLPPt0J4AzskdMaDz5SC
NhTdgAnxIpe7Rnb8yi7+J0rUa3U0qP6ywqmG4Sbqn9fhr+F8z1lagOW+mfNcQmFQ
aOsOhHo29q0zmGaDWG+ueakbDFV5hnRCR5OpigxQxC7Qn1bnqM86UQvaoIw4NqBH
JEvNdHaSVvpDx62Qou+BRtLilFOM/x67n6zpICtNelsAEJGc1uU2X2ftora8rph7
xskonfQTvRQjp0+KwI3PN+j6fg4flMPI/JNBMmm4ZIA2eAW7z6vr3LNXYHXyk/Au
880Xyg1a7e0HjLoSKTRYfwKcwo1i5JUV7fwv2HjEADqJLwrxQVHZYqbZlVwbtX+J
OOVCdHhnLop4fGPWGDq6x4mZt71ANwFNM2Owqd74Cf9wf9Uy1qjovQiieetIcDY5
LMRWQ2Dsb0fevS/M7efV6VY/y63ZNCumKVoAZ5CXJSZOJ90fUFKyhxFSirJYZFSZ
Kf+SRTbFXJhhIqxTUAoUEDAptqqRhrUJDri+nJOPstFwq7gQeU6LN3Wt8IxFGQ4K
nZQWaJPmHQBkLvOd4MA7ddesqk/CDMZLgt0QxDtaowbZeWSjyZlHv0q5lAbsRe9I
xalpdG8wgKmNpk4NLMCbyWpDkFTXNjjM9R3So7+BhqCYjHQmFTbG3vOiHwzHEs0K
9IrR5WsXO92ahoF+bXKuH0AC6QenG0znJ4LjJ2D8YSYeVFtKdbbVweP1UtwSlm7d
Hvw1PKt0iMRKGpP+riq1m7h6/rSoMCKbzMqLT2iZxSX9qzmRRK73TGTFA5qhyd/N
PK8sa9ZdIYsN1uGJN4Tv+vQnHOUGHH3jsWw1zj89uO1MV5RYl0yjUisOFe8a0POL
VY4lxPg03txfLxVBmdKb9jCqElLCPHiFaJ5GB0kjG9zhlnl0/cwCWpEi6WGxW7mV
3RpFlyZT33ndpIX0EMP0TMeLKjcoD+Hn/QBQJ4oCEI8Mhw4R8mhqywlv4jEdV0uN
vOq9i1Sb9zWLOwBbdLbfvNcAjSse3AZwOEW5zkTM7WlIwJ1LVz7LFPsVmtkBjAtG
1Pzcupk8QwlX7SlY6jpUtGfjRFV4j0kiX0JjZp/pObyo4JFIXdq5ADkdh6QpbZL7
xqH1HoawW2DnOI6AzEW+n8VcEdI3qMb6U+pdcjxTM/0BFeMQOEf6deVgmpQuePb/
ZKuR7ZPhO2wAxNFdfi/ZjDY3msg9BqwJYeAUoQVo5lTiEH9OLCYDBcoZtXqQ+7NQ
hAT/ldHcHkPXvJKnMsOB/yyIB2o/MEVTVh1rnRhvdFp4BG3HyQ/5wxXRL092Zecw
97zA7p3qRgRy7X7ywXLpa7B1N9jhstXVJzTJvLDKGJ5rnzOrn7O/+RQg9jkOAN59
HkLb6A2AhhuRehM4Lw06PEPDjA33SKh6+FGwUkpYmXlQXvpeTdwKTL6HrFF0jFxI
O0s0okZPZ4//69HMmzcASAK/0Hq/m/fNrYVeQ1om40Ajcg23zuIz/JdD9/yfMSx8
uyFh6982F7ZzQJiLJTmge8tJIyXDKyMCu1IcpdK0pczLDE28A1mwMkVrlMbeh8ie
zoeonD1Mh5vU8vKLB0U6DDe0kxs0M79TSLn5G517H8+DS8v/w+qEEuoaVPeOMsLS
to/MyHRF1IO9s3oqkSXfC4mdvtsORcBCM9En8WnjwmQJRB4Wrs5nA6WFtuUYe4D+
zUvY+EX6CDzVOh9iuEn0VdbQQ2hIbjtkxeurgf35MTglHx7OFZiMm1OJLVbQK95q
vt+m8Sde3D3kkjQM7euzEYGYL2MV3usRm60Si8H9Kv8FsNZ/0l05YvHEmzLGsgA4
BL8gLmpLpbpnk9KDHL9zVZEdD/ADe9Oaw6ycOC3OzkwqcapFkPIktLEq0fhN0d/v
c5zZsDVTQx5rdOGhnR+okfSMx8KBdg8HGCf4edisrGMqkwBv4nUBIz4Frbr2cI4Y
KnYhQd5D8kT662zI0K6OMExltHsI/d5MiwJA8PC4aokiP+RpZxnrai9q1yixzg8+
MIxPW1Yo+uWTsaGyv1FSQDYE8CO95K3L8OLAZ8rCcCvgSkREiu+TUEgU0y+vGp/L
qbJcO3n3z9mXzbunWwwrUf8sxwLiMwkZbnxDwqc+b2bOuqTHGVTHKQVtt/4P6+Mn
R1yijIc/96bNf52NYq2grEHF+KeYmumbODLyYgRY0ph9ts4XV3yHBznNJaUa0Z3K
chWOqThC/MQSvT9j0XX+Ip7rQEPqyGEHlRKZwgpNFAi+9RrCHEKI/VLaC127BY3Z
heO5H3pAeASdakcToowXpDrAupRCxAwBQWjn0bYACwwOhkdbRpd97KhK4lrI3+ki
HAaoQWBWs/kOemCy/yyLW97Gz92YrUwY1t7sSlllxsm9JuK6OdEnX5Fz9J2UjzDi
BiOvx8/PwiX5RcoQnoot4jpvMR8Ilbt7VvdCkLaI09/7btJ6IgqSmsrxFVZbLI0A
UpzRJklDncRmELNjnfVw77PHyEsSq2nzYDq5jtgnikURsHddF1AInYp2abWFgiTW
xwCjfEzRCM3Qu05pMngmBEhe1Jhu9bkdK/Ali+EF5CG6HzMtm9QeBJ4BxWh2fb2q
o2h4lyFTViT/QSFKzWs9fSjEjxG0INQbx/k3fSlxBUdjffC3YuvbSoVxT7xaIN+h
oOro+nBnZJ/6tBeBLqE4hLkfsc/u7um3Rcva4mlkXxsOOLtg69N+Yhivx0AE1cOq
A2FfVXCYpXM1e+qix5pplZOFhTZ5IRHlrynitwQnbPUlLtu5VlZgIw4MBgri5LSr
sctuqmSZcs5MxLuix49S7Y4rAWjsR05iMMvArvNZc/G9pFCd6pbs/WWeuZQiWGex
n+CKsHhM3e7NCbyjQe3q8O25GkJc9ILL3qxfFaG+az7yKkZadnj5/Hssu82+GZio
NkNBeX3J/ovIgScoTpHJNdzbgKvDfrVuFnLJoxj1S18Hc8m3XJNv73ybSdu/A1EP
HbB58d4QEKksTTGfGzoPcmJMhV2Mc/E80hvQCvxspylG63RLorhO4vk0jAqxVqge
4iD3iF37JEhXWvLrODc4ZC8ZYu5F0cIY5Xt40RgrgyJJKbwrcyeTs5xuGeyjR2TN
WaYtrF3Y6vJGSD+juqhylx4d+MR2QvGTlWTpG1C3oSU079lSJgHT9sxupKfwTp/c
EuQZzmt4GqxOHW8RQKgCaEJ5nWLllXK3k2EvozT2imNNieXC3NzkmeItSM7CmKLQ
6ScLIBPsyKinLSz8AuP7/RTA+0QetorNW7VUqTnyhhW2dZbwfI3D74S9swUI9SB8
CzPrqwO8l8xGW0PKlFLx2Hukqas/HxOheYnWw1EfWcGm+H3jymqdjwWOuOywb68x
IUL8B5q3LWGXJ6NfP1XUFt/szKKceOGit39UR/LX4GBx6S1VoAKrn5HJMVJUDYKh
FKgEE+cl957GvhYylmhVrBGYOP3r3TjcOXQfPYjWudktuZSbZmPl4sQgHvHMWZEh
zuFtasIWlznO1YvAKF37e9PI7PZA31n3w2zJA9duR1qRIO12TdGQN3oM4qP/LeMR
LEgF0dx0yHD6N3//F+aG0Eg5AKFUwC3DVugk6HYEPBvpZneHmyHIVU5DBEoN/Xla
XfuTp1Qar+AQ1LsRCjaS5AzyM68U1O8v54z163LP9LyDRx5she+sG1A7CAnHCNUH
6qtMwEPbBqsMHCpk9mSSf2Q6UNc6jvU+ADuPFuFenDrqmZaOE6vUTwAcEJ8X0ZYx
NmxCQXx7v6s4jjdFF6Xpkfy0wtdmNGDEaIvASK30CA9vtWYcFrWjf1H1x5FoOn/J
SYnes8lCez1y8IdXOkHlx64qZttN53Z6IGCbJnr/xnCMDfLoY33KybVDvAhjpEPq
1YI8dKMQGnP1RJoUwnyv2gLdAWjjdf4SidvJUWbSUYsbge5AGWxYU/teQf9NUkZE
Mo9kavTN5L4rfdbPEH235i2GYMu88TJfrsx8zPqksS6AevBLUT2NR92Y2QgDjSCd
Y+L2npkBGUVA7p1OqnsZtju0pg16ziWTovTqrdl0DOGgDtZCxyJzAgpqB7FNqK+P
PLAQICQbOFxgRozU063m8TP8huWZ249x00tRdl5y2E7Okb9AJx2n7yOlqbX0SLSb
SofvzPW57LMsQph7tkiJa1k6YVwnUU/Hl4eL5IF9ip2+WPLY0c3tkqFUHlDOERbT
kTlcUILIRFvmH6DEV1fqDLsvasw/mCaKr/BB3pd0H1MaM+uQrLvNSH77uw4GYcxe
Kmq/hzFDRoQP1HATIEAaIZZ7lPycJV7i7jJCuGvULHU9JjJMtRDJdtC40eOFP9Gl
D/xi8pu6NiJMQIHfsUHrLX5uUpzdHDU13hZYAcaGtW8lbJU0VybF7wwP54Fm2lxu
6yivcxCGahWzaGn7YTLp4GkXy5ZZU/EErPA29BNLw5Xef/oJnkULi4ap5ZdCsfP5
YnEXWAm2SKaPyId/ZSPqaHY+Om+SS4wVCMKoyvW1POP3GHJQy0FmVdws8F8Sp+QD
sNZhQIeodiedWWfQPrp7KC6+bw7V7N3RHDuBFxlVS8K3gta7U+OciDGdI027t/5b
6OnYCkO3o2/AajN3kUm2coJrEnKd52Sm8IGhlMhtn+eZ4N5c9+q5GOZwUIIbO1pt
2te87t1NDwQBvaShBeNZlBNnWVtykdfPjRvVVFZ97VaV79R8Fc2FTRmr1EQ7t4LW
ZtS2FNy6zZ9sRDMXuVfu1RhSBPuZ7vwzrxRDZ5s29p8j69RmdXxoxV0kGuU+qSq9
urCf6EYM9vZq4Lvz2240JWtXHCDqeQ05GxBf4FdHjPXJALJZ4mgvQILjoGqQ/vWW
6cc4vhdMwoiPuZN4CLZr8SFXs3Lz0YN/bl5nKyNATpvHg2+uPVKvgD2tbjYkAR8X
GmMt68k2M9NDd3XBoAySDv2D0WJ9E6W1ZtWQ5aEOPHFjUI1DpbOfVMA6mEfnQyJm
BQO+Ey+3w1fpiX2M3pFeBR2B+MG5Dd4czOPDcbAbZsIzTbNQgmBVddorZusNgXQ6
rwmba84AvwTeJtCmorWqq5O3M88EffCQR5NirfTJK2dRQgmhkdF3fuv4DdvTwJtI
3uWBAjL5Am83z8AQU4PlE9MreE1c7LRVuZMw67lvDjLG1EVZ048bVtMFL9ezneWS
rGYfgeM6xUpw0WisuVjxEhs048mJNbD99cJYeYANABw3Aluqiqu+BbE4v6DKL/lF
gBcxMBRvG4CJxkjZOPIgL2qGaiX18SDOQKdQqsZSp/uL6f+vOiM3xAq43Sg6/jAm
upnyszuS5IkPrWDO1zvVjdGUy9iyFmX/TCX6tYJ+3VWFdzs8ds3MK7ferNS0j5Bd
hU/MEujfGk1OuGYNEr9+d7ItsHyQRo5ol/o3HpjAA4AXIsRmNXfYP3FvckCO3RkJ
FNbmje06VrNo6SLrdpnltaW8e8odsq3xB6yEAWCxbulh8fqS3cWCUlUXA+yHc4dC
cfxJIMm854AXLjALrijTeysrsETeYfiREqXAzvO50x00z0zcJWzwWxX8btiKDEED
wg/RtIUzXFYiahVsM5XW+TypyH6ydkXc64SffrD7t5k4ezugm5RdBRFN1Xl1xpif
wFgOskprOK04p8PCs0cbEjsIzM9fDC5Z6PaIbdg5FdEi6shfnuPhZF9NJiCoKOvS
yS0ZpphkZQfuc5kx0ewJ0i/rrK6JeEHg0+dJ+JQ4BTpoDo5oo4LoGYPe2ZsMyRPa
QKKQMEo0o3RF6ulN8uwoQcgMFURNt8pgpmNCRYgCFvHRrfTrkvIeK+2p/WTLvW4P
WY1pqHuN75tqzzZnmm5CtEW5uq4EydfJCbAJxZd0vxuO160xx8FxN4HbDBuVD6Rf
1SSyRRxQtMNvckWyjXUUsJtOr1WVB1uumPyJBwqABbh11sd8naY4e9dyVC7ux2E8
25LaJGQp3Nej945UTTW+6Vv5RKQe8y6kJms++2hR/ycLk0q7yXnghXpgmjWHutSN
1iMqOcxeDwDjnPPbUD8Lq8yLFv75vD5kON3hyuu1kIWsRf9H6vDWDbdYV8ZcCV7e
KisiDW9533wcxtOpTmz72T3UWCCe9dI3zKOhj6p7GWfABkH0PfjgQu+UsWY1KZmQ
udNKKhRm6DG21bFoDl5zluLuFp1pXk+nwqoJvDlkLa67ZAi6oTep2JoJ8yBQfW/d
BL8oqAqI9cyOgbCyfSIJyRx6pAZ0mxA1TeG9Za1sQAP1ROzxVIKdhLsextri5bAA
RkyBR58ybMu14wfrv+oyWLUZkIo/wXHTpoTQO3wq83JiY4oZbCrx5IPKLR6KYYY+
K1XE/fdAB2h19cjyiS9aZNV95O7h8qHIqkAtJl2QQThQGFdNco1iqHu4A0bkEiiA
kt2Zzw5B0nIZZOf+lKiAK6gNZHnqnmbyEBlZqZ5iII8Qmnd/oHMShB5YvuAapoUn
ScpMoNm/DT7TwZKC3y9Bg99w4EgL9jjoBkDp82SJhBGcatHppY22QEojFPty3pdX
Bp2TxUFmLOxye46zQIMeylrBdx3rTyb1jbdczr2Jou2t8ylPZClgxx/yjIT287iV
sJ2Whj3CF5cfLwjctO24Amqyr6ETvxNV6OBvXm0RGNjOIWLi3qIF+TYn0QsaSIDg
i9g/oyW4y+dRpwd9QA4L9MVjIk4IrIq6NAqk1vm1cT+E/m3reh+BBqkakAHjujAv
7nuInNfrwXxjEGaRvvhU340zDURif0HZbRoJl5Dm7NDi/8w0spNBoOHgzRFiWtFZ
YIsSQsuFlSAX7eGkIOdZtbMMXMAdfLIOZW3Cx/NAqAkiukdBcCT3Sh3HwjjubyGQ
g3gGW1Bcmf0aszIASPce9UmSim6sPkhWzTVt5QpW1LugzJFB0ppUsth9JMgvONmc
f/pnjx3y5NKmMcejzUyL2c4z4DUqtQPBAPszlNINs8BY6P7vv+IndViXX4FNufbj
Dy0R4a5L28Ciec/vitRVaMZFemMgJ5vMypu25RbRo0/uiShqXCi6xQp47saDb6Ww
chwd2rM8o8zEw3b5tUU7hKaXXhCDuonkhblHww4Xk2XApKIGkxlKMd7ABEO6rYCg
v/m+z+fSQqQkYUr5jSGHCQrKYEvQSxhVj2Ek/w9Gb3NwWSdfJRg6BeDz5TQvBAEW
CPoy39ioUxftJSHbIPjth3iV6zztv9otiVI2T4y/LD/FtfxDLZP/xnCwgKLaXZ6M
NWW69KuHsCw4GJF/FguMiffDdGQZZnYvT7NYCGTFRU5EfAqeiYZKFqgmBzL/xf4B
tyg+8JMoH2Jts8XCVi9rEjDzbDxjMHOdQ/MuX6h/K6wanRLZw5z32nEOcZ9sMzzj
pvQYqiuM9Dgs4XIcUjyYLUP0w30bIrklCGvNDWE6crTfyTYpcCjG4b/AhtNOEzaz
o7d7rcqXtcTE1tEz6QaR1n30Utb74bO2bGXNlKUOmJTH2JBxoc98d44w5w8s3jBB
zPHH5Zvf2eXCgke5n664gUeJKjid+io2BMoUUGOqox0KY7LhgQX76ZCPUTdZk54c
/eXC0vkC+jXYycjWLVB8g5QBpmRkWxRslK5XKwSDUlvARwuKw0Dm5+OzutUcuIeD
EPvjYPKfi1wOnl/9XrMf175SAwMaN/NDEfmpYqiopo55Yt4n6vA4fh8IM4jbYe6H
LKRkg/OwEAdv5HHPa22LSsVaj3kOAeBMDBLEAEmqTjBLTALn5JN1328gaREmib8o
ItWjLQqH3CyoJrMrnAskk2K/MHQ/U16kh0zrSeJ1eN2ia+uq5V+Pd2s7Ydm+uocx
b5wvSpfd/w1IFSDgBsWyS2eipSXgKMYuEx2tBdBcGX/WGlHcMsBGUC556IyfsSgo
eOC8r4XVMGIvrNk5F9RkqSnY0H7Yqe1xGEDeUXKnoqjjulM/zDz4Ci3QAFfVOjl4
YImQDKtDmsez0T5n+jmPH4TOqp9LOiYUFDXSF4S1RzeNVFyWJhMpPSMonBhAnc/Y
1NhjsJdG3TJPqjp/RWxTbQeGKPtwLHOwatN84mAsco+TJJ70KSQ8tlr592qXEJZN
IzgKbAs3gmiqPxonjxaLBK262v06PH40ZDvfh/ZcloWbVhW9es/WXxqKwKfXo76b
Zk9aT66XzFOZ0c8kKhD3oKboeeANZuMrHpbXMYXIxhsAaRJAF9VQJBf47wZrNCCr
eJ8mhBZx4dSojAA901cLLfc57m78WV1gT6voE4fUy8T/kUKEYL+FGvIXP/Bztfta
zmZtMAG/qc9yxh6454oy4kxVW/5y53ckxZI6zB//zi4xDZS+hgoh9l/6dd1nEymW
UXpeAfydBRgHfzyCqRg1raT8+RFaylMsMq1/QNekMgBpL6EhZ3jCTEKMYrlwlFe5
fj+Ybemk7mqqsbxF1s0xcn4LKDksd7cMh+v7D2ZwlS4erUlSh5vXdypHzYBd4cOm
SyG4p842R21Yyw5GCLZVw07AGz458gAuQDoTzmzE0BB/xIU334Dvhcph65FEWGuo
3oaMeRtNph/5SPgg87h3b8/xeGQXk5PIJLRTU9vy9K/GI3qTfreNRZ78OKsg0BMW
qcxOqE+HC4gqRxwX0o3Khda+IRXyFXP2UcXKgqZf9zmBzb6N+T8PaNPxg+rW+M7u
3wlp8e3kaIoGA7yqzjt7cOUbGHK2KLYvukUOSuzBJZ3rr1zi/Nw3KLJsvXhG4iGK
D/BBr/UK7LMRHDQvEEwlCBiaw3O9XBjFqdTt+Qm0BbyF33LXU8uJVgCfO8GZne7h
JpkN0+bIncCLfZhSf+ud14zDOOoGurUzXzclChGFYgpgpMLDebtj4f70ATpK+87l
hocfadm3VdkmfAZ6F/LpQDfoQYI/JmgJTzv/Kuvrt2K2EAkgxrKmKG2OWrxl5mk2
KHmUAB1o/l1c/4YGpZnMzVIaWYs6qmy0XuXOHzz2507paGk9AYSLKJEjLiaxnEHz
glDyba+X+aX017EXElJbkWpr4y1tE71HE1TrfLARN8Croqse8tW6fIyMeOnXHl1s
VkxVxaLj9cCejLz+vUBiTJmYZN3yXn4i0iEWkukL0lV/6Z5yr9a1X9r1JOdTwiPH
DoIEQJB3hUahzTZL0HRdxOF+s4N/n7JN6kAr9HymXDIG4D31c8qwow+hJeh0DKgV
2kqGtRE8OGM6X83zRf6/gkkuUEmWGqtsbeYzWoCkNmNBjcN7MfaVB+e74whtngBw
y9CUirFgIkfr7yoYNpWLIJbs2JWSrIVRtZdhpNMUs9tGQQBnFPueRl/52yp+rKxQ
zlHGfZ6nvO/0lHRi4XWdWJhlrcFsSrMg2dZ/FwHCFenMUlbqavLI81ElatxS+vx2
qzYsclq6Wddp2gJixJxveT0hZW2Z1gzcdAH3YMXdZDv2AgtU5S9HphFDa8KiuGvd
CWZQFkVLQ3+lfYte5246ufrULvqsvEE19ory6j2YspDGABDLdNJeuqChqyLcP3L7
RrDlzFu+LhISQD54JVLC3+X9s8bmtndBUy5xPhelPUbJHR0aawKTfqx/18sUUOI7
bE7mMTo+NSDQY8FK0NvThUPw4WnB1xOZMyx5vxw7XU0zPc+8Hrkye7ljCfF2bGRA
h2ltadAgcjfVelrIKx0mpY5ldefsLzNhygfA8grQB2336U71SS0T8zzrNOBorFUD
d0jd8UjzUOOtqc7HflcvBLb+XKaXeHmXaSpdo8JEVVQ7rFO94pdeMhW8gCXiipGh
uKBOWB3wmETmn0zAh3IFjnAYWHzwA97t9I8cQQYQDx0FF5msaAsUjWFhALnn2kNe
DZhR6u0RQRD00Zy5bQOMJ4dTmyifIvKfvRzDEX7dmBgVDLRHY0HxrHy3Vj11vzPL
oE0qOT4eEafyC5mqv7lwTQHvkx08q7sAbXDljCgg2xPQKL80POCZuthgi4zqJCY6
3IUrx/5yEsQrl+ptJHA+X+6uKH64ELxL8OeA8BMyHIO1mKjld0AD691WwmnfwGfi
FRSwcNlgbXM/d6bRAFD7iLKh8AriHLbBFIVpKHzGS18j+Y0Xz77HBlXNKHA7HFKG
z04VeNKpL+dQPLrtUtBAMfcE46TN4OW47TSEclCCN0ewqW960XNWkS0FaQL+1cjR
3Mo7YHvPDgULNJaZvUrdTVQ9Yn1UdLy35Q13NorA3ZQ1njrjHrdoW7BxNQsQ6YZa
NEiz7xRow2KToDpP0POinkJFoEgSCg5jf1ITXgXuo7A//4mIqQv7Ek7t4HYVdVYg
5LdwytpAjV6+o6QyOwjJEwvgHK3nQmke8qn0rdgOoqrXHktIG0w9y6R2sC5/gvo5
X0U3m/tSfZMOdB/Y+COicjoCfqhlrC06NMYOWG1PdiDzTgskWe0NEv3S9abciBdd
8gPe6APf9hKci4v1OD1Lf5V1kr1rzizLcvajmmx0Ul46L+LSTsc2PCvOv8G2TMCo
ezX3K9vU5zoPIQyKi5mEp6GgoE8QtzSwwBGTmHvG6aXj0S/ALPwwf48/rGGBq6uL
leLPoVp4jNve/f0jfkjb3KVCXhk4bjLLBIV2sDL4o4m/qKadqojGjFCHW6oFrShe
+h+GdkDcht1aa1YJLITgPaVVxldlE26hknX5wmUxjcxtC063KO1xxJU9ALi9q0hv
yAb0krq2P0nfbYxDpeTFVZT4Uv3y+iY2V1Jq7U4nsH76cNfJTwq4xqKOZ2e9ogxG
uVvw0ipADprWIfZwVeg/CGJn5gAgpULn7CMoUP3Dg4Izs5PiQfPOUO/b+xyea9qB
CgOhJ589eR2xxzNLXl4naNIlz/Seadlf4HG2PIQtTyHMyOVF3lOobi1Onebi3dWA
RSZhK30HmnCJkKL4QQmQ8fy90H0kD3f/Mo7ap3bfHPz/iu2vZ3qiLPHQfI84fPrm
tGKeKcrszY3iMnShT/P7yKMrNpTBxedOs3X5I4v85/C4pTRWor+eaPP+YsbkZskr
rHUkwKYonm+WkCioCHSEMj7QRtxBuz4LVAR5hBtrSb/YwwXMZXQas9v2e12xWQKD
OK6ARRCbf5CxU9CrAw4tbh40GAX2XqIuqOYe6SZ/D5vIFBoGuQntGyOIF7Hf0zoM
OKDj8Sdas4sQShwvvsdF2dZjzQL1TChXFO1zNSAMBFpV7jlPPaFr4tXJaJPZ2VW/
vNxq5CiUaBiA6uLIljDMfdf37uZXwIQR5xlA6UIXyktUXGCQV4BiUMC3B6B2Fr8Z
orPflCFa3r8r/f36CmyoPU/31tkd/eQl4w7yGV560XD3R8lOoJQATQ31mNvrlJWh
vELUp+mOqq2wLjMPcB4SfwASBdHUrXXzpKUyLUrwdp+w0KvOXNk9kfPvTHjxbZa/
mjvPOSzYVFBJxTL2i8ovhVVNG7EtkIC9sM6kq8bzL6e8z0kTSR7sb9BeVlnnW12F
7iygKYOc8xH+h+M5KLZF2DZbb5+9hTul8hfE2j9XcFE4m/FxU2r8PlDrUoGxFZLF
jqj4Tmo4m8yDerRnv8XgSBh4OS1+M/+eMbr6cysqcY+L5htXUPUw06zDDbkjPmNL
fFcDtH2SkrX+H/ai0/bFDbBqcoMGnL7emL40U1P7/DoQG5MJKJrkZ3fafaZdgYva
Jf9K/1vItL/D4IumzX+3M0hlRz7/q05NrBCexYojg+sDezqoNiB7iuNZRS6dPEym
TVsUWUGvpPDhymwitnTI8DuN5vF2ZGhD0aSQtwlSYnWng3CZ3vMNh+rnzO99Y7fR
ArU+iodwjI8AwDxOXr17t6s/HmJOCA+1kxWevw2yhDPMYhso+66MAz8qTsurMZy2
a1H+oeHUcFtfLHvE4iPExEgzMxN012En3vi1liBZqZ+SEBY1jzbojJ3J6VnCqBZV
LExnroCaKXNtq5F3AZlyN3wPMdpFQ/BggUDLwFMLyzXWvhSpV79sRqiqaTgVBYCJ
13ZDa/K3oKawGoUeCgslrGe2ssJaGLX3O5O8ZCwwOGUlIaptgNaXnbvESZpP+8vQ
QhNlj2aFAY14WmUta90WIAnE2oh4bnnDzBNXajcG6tXt4LfE0OwZByhBnjT+WYwu
fOLPuIcXMmCtNQkOBTofOPEXiQ4KzyG0bVpfPtbsPzZmXpadMPgVub3aGPPClCcB
X0dFCkp4dNX+EvT/Jz3wMzAtK+VJBZ6gnccYKOwZYkCEtlIWSDrkivVW5f1edGW1
VuqXFS04QlbvsnDG2Cm/FlgqLea7okbezGTlrXH39tqOyaimK7FcLnHhCX08xtm5
GK/YMPCh5Ci1kwoxWUJGObr4i58T82ssZsX/rQEjtJEXJ1R3esBiRjIpNdx+pBfA
RAb2AQjjpecko70Vc/Aq/zhmHqWGnO7mBRzoXmgPbbmBUyoTGFh0uAHcjgJIeA2F
ZI2ZEE/1I6oJTwkrR5WUSSI2DGjsTr17RjH3ttntZKZCnCP7CDhzEVvJHnJwXBR3
KTQftfOejbz084nbFUKO5voI5HrOjuljcOL2dpyeZY17/Er9coyhw8R6wg+kP0j6
7Hxn2u0NDIw7rKOGIwamM92y/kuqTpjAAD58mLp3fcNtQ0m1qPRW5b8NQ3mn5eH3
sRyi4x2t18yF2AszbExHqUcekDyn8Yzk4OJ3d24oB7i+REkTp59vXnLTyahCq6bc
1qA0WZz4qIDQ/BgeB2B4ks4U4tfOsGXaxQtN6Lx9FI20Y2IsJd6N6EW6qlyCJOZp
PWRDTWpoS8VsUQ0vcjH6aihIfltAOS7VKviXyhfz90GD/P4/BEZfpOVg5GDxs3P1
b5mJTz5UMqQPZ5zbPDinfR5j67GaJgTBQiGSP8HRZksDXVl+4zQwe2iKGCS0QTW+
rrn1nZGI10vwMzM+sUyA9Nn0WxgOiDSjcEwQJoYzW0gGCWOeCb2vfgQ8UQ4O64wA
kbytts79KQcHe35ps/nxnz4JoKs3fxFE6hTiQXepUe7mJ78Mg3gtJ30SGndMVT82
p7Ct2wPH/5g89Rdqvonu/CGHdPTx3NiLQdAkORG7M77GcLH7hKcyCnj5b42KeaYm
IFy88z2orJWjJnpebEO0HLTaczpXZBWjNI7JJ37JczOx6xXFl5Drgk+xKWRKUw89
byel/hBm6qhAWVDs8+vsJmuAdhojWhQUsj/u1rfUQFgNS2RK25igB3SuH+Wee2qh
hY6nDWbu9fRFXGwU5f5ree7W0IX6KK3LyYR3Hj66g8q45KB9C5KPEYx6M5CQbeeo
I8kSP1tY2E0X73nn/HpC7yLbR8Db0D+ZjMiOriGOB38rB1OTK4H3eWfF5H6sjD1+
s7YquLYlFMPkyb3JazNsqujOI957ftTMchUJNlN3eZ20yq0uGaZnTa3sPaSCKKFS
MIyGNbD4sMULs5qdo79Q0rulMlSvwxC/5vvgJWHixvLNVY6C/TYsBiU2wyqThk0r
m9Wn2h66KC6TcIvyhpzv7WwYdCbdGU1jzuMIN2aRLmSeAI9htFdcQZJx36TS+hTE
uoO+fykw61lFfgbYBFoXeBd2tmQCVTHw9Yu0i3uvJqKGvmJy1Q+jvhaehoa1cdiP
N1Za0bBay2XwH5XnytYooBsRVzYqc7bgkR3PBiXjEv10fvMCi25siwr3KVQQDat0
3F5+cE+cmQDixNEPhuWKnFF2xcaioC8K9D78EqdcvZmPgsF2cbfyZ7hhfVfsMutq
U2ydouLX+AoUua0tOoqXPNj5MFUUD6qNIHK9m7VfHGzKu31ZZkEb3h5GkRUOHBgk
5nI7TidPb6BJ/D4QdftpH4sZWZ3GlJi61TeSn1IiQJ5QNd7rI79G81/zfWv7xyQL
GGGWUIP4bwxVT1u5XVa2ty+O51hW92PWq4nYXXaklAe/KcRfbXK/d3ZN5VpgJjFv
gM+0TjeJo7ZE90cnoI6PTe632CKLgy3zHtErin+SItvrDI6Z0HUYnPKM1p3iJjE+
bPbcCP6LmBRjBR+N05h8izTY7xEU7iMgLGRVbaLu5gDLB1aHlqkuIff4B0bcvMvf
UYU4yJC+0aZB2sLWAmzaY5Lgs6bHGjKiIUvwhgtNqto28sIX9kx8+D8Kosk1d3df
EX2+PeRRFk1nMxWo6WoHqhLMF+SfjzBVKr2sHSI1iBPwicYAn4GkbYjkqO37qsbb
Ddv/OJVVipe09i3rIECdHRzapM3E31gljRVikRhdhwkEiOER1jLEE19qJkekoINH
xaBkLONrsYKOzS6I5iPvl0qTxNBG3/hi4p3/6jfIUfUBO+HNmK9wWWFkQTQcZWJA
osKK5gmw+5FvEbHyMumhvChjmMmSW7DJK/fsuQU2O2YbIr5hFgYBT8UiAGw4UhmL
i/sYUNFRFjaVuE3Kj/0TPnHBbWl7ADjKzEQ7oID1zNBu1n14N82R4oycch3tRL/S
KIZWw3N1zY2WfGwV/aBK1YdOOxOuFaZnEYVPobSOjpo52HCqPIWPAbpXGG372ihd
/6DHYOqn56TycyL74isLjoqr60hX8i45aZIiD2GrIPN8S8PQ0XuAxMyngnjrAppy
WjRZsh8oly3YDRg1KWVLe0lzdYihzxrYlweKMCdGD/857QtP5n7WJOzebzpL7qLZ
FHvGgj6xhrUx4Dd1K14frQpASLyt/6XHC0SHohV3yFA5//Q/vZwF9Hj5XzO6bDIE
3i81Jb4A9ZdvrzBoSZ6kmcEbZBmfdbcEQ4EC8/n1zzIXgNoSSSDEFxMVHCcG2z6B
JVKm9l8CFkIV8V1TNU9FjPiSyPiyq2gI20lwx1PEEq7Ojs9r+VWxTk21xK2XfArG
3WCeh1eq6mMh5xNEMhVSsCA/LF8T/nVD6++ICcqdiiyhtcLW9LF1a4M4QiPooWTw
L3PxcF/+csV8b5tt+2LIoj2hh2cTxhSvQRtKxaPl/XB3dZYx1H0WfmgEsM3DKFqT
kM/INPL0aCKlXsVZQC14NiNEoGVOEFHplvYVjYSChC1JGk7qsEP7ef/maeSCsII2
Q01QXcXQgrMaPhA9vzCA0zp1WZlAHGdWeEPcrjv2HYaN20uRudvtUDhCKXe7OVHY
PNGCmM/OZE2orGHmzjU1jKn40kI8kT3okCkBgyCAs35fXDBnk7yRJleYXq/IAJyL
iVhrwA5JSPGr5X0ym1bTRJyguJXM0nZqNKEL6TVGwFL3jVkXhBn72m+4Nr++RvDm
92+mAOsRZ2RhhZc6L1lehiQuaK+WIwaBfN7k2yP8M4QyX5i8k/sdB9zK2SeVCHO6
WpQqua5wiWbT0KaoSG0XdJsOArXWZWWahh96yhKQWC4JjNsmub5OVj5VcZH1Vt43
tYDiN0HjTfIYuPgq1PvcjYgf3dYiSSfHv+HQb0VIr7PCrF3sFlolCm70swlhY353
VjBsO5iJYK4wiymZimLMuXGz9cdeq36T0+O9EcYmCGh/ja/O5SfC7rvZfdn5GZ3N
LjPKmvwOu1swbcLusjgB9G6wBNQjkvpJuq8LHL2SbV9s4gtS1MIvDSM1AV2B9HrY
xgji5PCFdlBK3NEkKVqzypiLo/db06jgQ7aLb0zk9DlEGMH5puEiYeOYNaJQc+kM
CdpPJlypbpSPpqG4GhfE4yYgYz27Va1BXV0w1SjVfc4fucJKI65nRVICg6GfTvqj
xw7IUEMeIbhLzG4HTZYWUxrBI3/IZ9UM0oWl3Vl82RROzDwKc1nI8+TyIrRXQ9h4
XlSnO+lQHbaeW6FboRji7ZNuu3506hQSp2v296lrcDGJYvvm32H+sZSBZZz302S+
jzLh0kQtGpH8Hw7G+//rA2wEu0UMfv5IxWufUBEJQHvQNoHWscWlh5O7bhJlgUwv
S2fSGzmBsNE8xLaEyi8e8sB+lkZWfGR6f0OLCzMA2VgfULx+0GtRqENsa366elsL
gUERxBxqTEGnWK5u9K16RSaPe6RjZz4ETvWJI8KOTh9HIx1RcsmPDSIBolOgM2sL
+1TSVcsH7zVk37egdYBZNONacnsh4KTPMV68zcHqcKJU0WsRGi3tIKy2ESopX8CC
J/8CFYROiRa2x+gGxlgDs45cB7GHFlgXyl4poDY1/W4Lh8XilXL/cc7JMAvuWWn9
OiSxUr/6YHNdPfZWutqrNIUVSu5LzW55y53K2bABmrv/UMHjo/NUaNGlXrlJ3njh
nX92Yi46ra4Pza0KlxYRIrKvuMA34lbL3sPK1u5GCfanRlDylg2uSftoZISIiaaZ
dnNQngwp+v2TkHWH8Jtv+y7lJD6ydm3PsH6IzJB2Ub3+onZZvgg6sj4ujWBUcLc2
KcWuy6tG6KIEMc/hEFc+MFMQMGBWHwz6IyhjdAJvHKaRKaFrwqjqO/ePIN6Gx8nr
200A/EeR0PZUjNXIcMEMS1dow5rTI9c8RxfMbve1MW/imkJ5OBr+/JD+PD87/VRf
1v/X8rbF5acZ7ou+N8XWK+WBzQA43U4/zkZ+mCJhAwTdj7/oQM99MTcl8yhpJrEU
OZWjhmF8VzxlypGNNuoPkNxvHI/xZHI/Dtp1zgyvGT2tYWEk1Udj+58CFMqbTTk/
84AmFCZGg9MgbPC96xrTo1wHRMwPRF6n9RWZEc8iV+uSTUZUgPRP57xkKd5NxvIN
4ZsjBDYstlbe0jeq0RHyHLEIk4Z2LWuTJuQhSx/y37OR7EGygQPXt9nQSngCkqBT
KwQUsRjsoBsfg+miiPsm7MjCakYSkLrcabDd0gOKvv9JwqujmzG4moUA6RXMPKwX
80wvGe0tFyyQWNHtjRrVp8EGqlKJ+qR26eHdO5rfBbT+k1wnMlW9VyrLSm3SwXPP
GNTIKDXt4I0K4Tz8ft68CUFen7B7zctjZ2AOzGQp20ueRWog7PVeZOo0kSJPhBsS
jI48znRfrFsOCxxqYpnlnENqqylm91yB5VhP8R3yNT8HrpDh7w3cN78sr1sFDn90
4Ory8W2cGu0k+Bce9J3CoFdwvUMLAn5XOjslrxuh8RIn7uNdPUKzUPBsotiGnVLV
d8+bN2bDseNfe8ULzUYH3JbGeVyrvUhOiqr5m44a0sdf2LH8dmPv1xchxfX3Czzb
5ZEvOoqF5R5TEyhu/ok90KA9QGmGh28ztGpG6SjcN/j2NwttNasTiEyrpv7olwYH
Z4tv6RhjVOXGjPb7wKyC0pJCgEXZ5RCV6TXDaVGg1ME8pki3b2EechimgQMmzTav
N+rP4Ztoh6WrIijYhYoMbtSP1SUHuUI+7CXAD5Gz0gkzDkvT+UGAZ+mfTq4mFzGM
kuLX0M8y7g48X7xkauqd/SqQkk9JrgrMo4MxOqRtswvx+JP6iepBJSeVGvQdkbWV
U8VrsbtE0M/TFY6/Fnd+ie+FGYL+YFQCae4AmM/FdEzRPFKdzUSnZhcRtoL7a+aA
NHnLfUbKZl9j1SNn1RR1sDPgis/ZsDiLdO7JOx5bAR+EeUHJ/LhEum+Ve8G/v+d2
ibiyt6gyWuRcmS6rK61hO4dezKoNdOqPXAD7mRSxp6dCtfY5bHVY9qU45GwjvKUe
uTSBdmGpF5jwuRpC7MGlvsYKpr0XnEr8ECSX/MqwDW9fvRO1z78gNkYOdd33MLsx
vB0+KgJTSZoXJ0oKz1OSvZSq8DCeMzYdAGptk/p+7x4LhCruIbjv+xfcY0k0I41e
zCOWXKkvF4oLKniNG+1asulZSUN1SpV5G/fF61cnXuJ67w1aaOVNTzUunev+StlK
HuNATPOj0th/qihuhVnycyB3GyJM9/N5xDHjXReZYAACa4hU17aWdJ0dokaeGHbE
Ce1N8U5/mfva4RqTgfYyPqpjCKkcpKHIkL0qLsDCeVHdNoI91j9zY6cniJpwGGt2
RX+e7uW91BMgqk1oT2to54f4i4DDZFGH5FwY5kZ2AtiBa0RmrfqgivOzs462Dn7y
My+4M6UGg3Fq3EZ2q9OOnOjRveRDU/AY2mREkbi24a4XJjLDNe9F6giFTURoY76h
lsMh3U9j/WtkbJkETrZ8OZN1/XM4Wg94c/iY8jhaF4qevyl15+cayK0dQEi91c++
LOxz9wQdxGtDnaim4RiMjgb1DIatUbw7ep/Dxnagr68gZ1zUHtHhCebDyJ2Z8STx
XaJ8u2FRLg5gKgGSqnuALWQfd8bS2X4fk5IBaotFWtXaXUQwmx/XOCAgL+FitL5P
ESnL1cjV/F8SZeGP8Q2ZeIqfHiiSXb3HyYmAx6m8Z9wvgOQDsIbNnwRD3Rfw2yrR
l8ZDPfUTnMA+eRyGzFVsCE1WoCBwmavcBeAY1dgSTfK8kKSIgOHP48Yva0OxIfsn
tDjI47lT6OGqDXEnExCeELcQ1uvjDwT7OvXFJkEq/SE6NVrLnbEzD4z0UhIiCnO4
ju0sVCQK3qcgg1mkzLDinOR7fPYfLZmS/XwrAZ/6hOw51hPgpt/K9WDw3PI3WOwp
SKH5aD8cljPHfIUYOhP3lUcW9strzsqFY5RRVIiOe8vnHPAX21cMf2M+E36Fnmn5
tfQtByWQpTtp0Zs2A80XI25Q5X9Kx26x8OCtYe1iDqJLdQcgVCnBp0suog7fqWYG
9tF5TqXiaKHOKzF3M4kJwDAr0ZzlDX2k8hXIYHz4I09H151eQLb16STP+p3BBkXT
uLqoy06eBQqlT+T5UjFw/OgRzYtxxIMBGK8fjcvD+ARcCKApaBkDS5jLGJPRbwu9
BN4db08ue32t/zfXsK4azD37Fk5+7faM8XSojHTHJ+73kHMUO7BIS385K4KPQBIU
oIxdVBXHE0xmNJRrSF/5DAeGWsIEuI3eZq7a5sBQS5Rtddm+mYZzzA5jCtOvtSUH
VxqPFGYge29gZGKddaSsAv+8Jrsh11cffIXsw0ZYSa0+Pf0XWppUqimo2kDnLdq5
mUecgdFQIaJm6LRQEr9rOH0Ua/9djM8KEZT0pt5OP2lSHB2IcZPjeEVVE/rqD5FQ
drnwABeiOlWfCvBCiSsr01ebc7gFJ8Zlrc/Vk9KcfQkDOaI/s1UzvCeLGEzDwCm5
p8OeHVk5KStZovMcjdvjOqlEuhH55FycNFAh/7KXOlVBG3X1Dxv9nQIj+L+XAaYI
oFJE8Rvb2FzRGHVwojbgogpKcvZYNRCML6wi9n5GH2CXuKJfG2IAh1msZU8KDY1O
m+Oqklsi/mh5Cc/DnmVI45XNRMRyGuZD4/pNFW+nA2vGZ8zDdpkCv91W2AyAtePe
00Apqz5tDOVQyYbqiOfLhkamdnFPN9CffpFJSDrn2D4M6z/VfIDYYarxBUsIZj35
RXIT/0Aw2Uoi9jDfOklQxw+GA0mZZpniahV/exhKbJNPfQutR54eofJUKUPRaAug
KNl+aPRdfEkACGbgeOCeMTWNb0Nog4PBUIkjYx96eq1lK3y1q+je+2t5Ydc+RxfJ
BapzVgObDmAlLmdXkWD6rsxXZlGWE7aErmfkKtLpdi5U5d20Ctey2u/TAQWX4ulm
nvKvhEb1WqU7IN+aY4giuUPNobRQwANx1+ABYPeorAiOYNtxg8T+62yttbEpKes2
OVPOMNreFX/EAPCnF6RyidI4wMJwu6Ax1gxM7fvkjtRUfp/H/UT9Fmq73oQriq8p
FV5kGyo5QCbqrNfYW68SJKdIRCchCiTrZSwyvA/B/IFgZeybrmZajb9VJX/tIf1+
rRWdw58wVWHbqTe9CUFKUGRC/hQp3gougk+xhcKS+yTvjpgc9ZgyDPzv8WdaqLdk
dOe2IajE52mAJZmpCU/IYXSFdsEUW0hG0Wp+dtiZ/4ut5zuyJ4HESFLcXCjkK3OW
dZmfh/33QtsZEmEgpt5XPv+em3KFV9MDGyflAk5W/U7j4imRqKiU5BEl936sNJR1
oI9pZRWMHYzBIUJybg+OqfDdKv3l3yH5Ibzgg44o0xX8DYYnK4khzoTCT3ISUqPc
fFqmY2l+CPYsHltyceaQgBbPZMt3gHLb7uhmx3LbC1lU/63RIeXNEieb24EYE5FZ
bZ5O7suk5M4/WA/JH42E1gDLrDqxuCrE6Drkg0GtrrxlFXa5qIk92y7120kQ+9Xh
UcqZXTnPwmPNce/P4SsCpjL8DngttM2QeTpaba4ddZ+liiKUAAwTIRP0z4WMxSVG
aUgS6Ykdum+ojK5GWWwBe+PQSiVW3AbXicC9/eO1cfsaw+d9PMKXhL7w60zea+WO
zck+wddmbJXNJ+1+kqymZmxAzVITxZSGK2QMxwKLWB40w8G7qHehUMCdVi1o3LNn
TVApgTDYc0o0C8HQXg7+fcHanTHBcE9jPwbXJHpNwXzVX/fwlBIHlKH/oSsvhPlc
41Rg9D/AinEQMlvGASeyH9x/Hb4FB55o0EMdEfH19qdqnnVN8EzQZn8V0d8b3M3l
a4sf+Ik+ouaT8MECuoLjiFAtEf+flXsAZGn1XtxE7NGmy8Kiq6Z21Ewb47qsMhfg
k7TBb4UmYM5HNXROvKdqs/S1os1GKjrOIdPz3kQgcFYFOenUyWWkG/kwELSmTT3B
QWe+aRD9eGNLslxVP+hFZcfgIoSNv30MOIj2B6z/S1daj/O4wUyTAyHgWPo44FTk
7KJXQvc/budJAbgW9Mx/bbcEvqnXYUfTwDoPmI/ASPbRkgLFLiuHL2NH81IMgx96
FkBsPclgMfjPNgIU7h25gfffvXkdZnObRNMqxjJEaPfOM3P6bCdM03PpX+Bcchik
mHWAKnN4SWmkvH7JgGVrCnN9YjepGdXKscYkWdK4eJ8nICsTG+dhM6HEiMRX/FiJ
25h4UtS397BD4uLY4T04LPbVDSbhPAF8DqGqrGKgRH7rvvUFFBax1GPejocmeFXJ
Fr/w8NPLEVjkpWbAKxNqzYNDjKjR99oS2kgfVQDNx72nSpKr3tIpOAV0LPxeuji6
jPZLcyF2S74uqwxNb/d2hlP4KCTfeBau7GEOqNRkJbQLokGbo6iKg7eJNsw4DDiM
btPpef8TWNJep7n7tRPa2Nx8eT9Ym29V4cT6iTa79yO0TN35DtwkTlKJVR+qVM7H
YGkciEBQyUhgEYFLLFWU9m4G/JC9H2QN4e060pQj87UfL/khO0/TgKfgX4c5+YpX
vp18enuDKI5xe5QZAn1+uweXCXeR1kmSmUz/Cn0DkYAcBDKdGe+T6mIycBaxanP3
fxNDvp0b7ILIyYfTBglUHKjUuxOmRAglve1KDHkHI3sN3CqUW3wG5SJPtriG9uvv
yPV/sUyxe2SyUcNJqzarD7jqgXcuEMKUZnQcwEvQ2R7iL4Th7LR3V9NyEdIm/1q4
8YLbSVmAuUDpP4iOnMWkDi42vTSLpGZ/FFyZCgXXOuCaXy4efGu+XAZ4V2oW+HEg
PoRMNK3zvw8oWS3LeDhq/ctqWmtLZMz7KTd+y39z8JbX2GIUWDcFXao/tZqHv9kA
GXJpUqnAWhlqhobBJby+iN75yVsbzKogO1L40M5Qd5XVBcT6Em6YTMLaM+6+XOu7
JScDzjDjwJaILmaB5IoGV6m1y9DsZd6cFteq9myyVuFo89dI1v5PoBGIf+Hu4xYQ
I8khAfw0Q1KtHMzDkidH9MwHmIkJV6LFlfTmOQSFji+LVWOeAoNHIFa0HHqyKonZ
kCVBe2VQOhjQdiWB6eSIFiG3aZpx6juryFKL9iGDk54MsVNFPgsfJQ17ec2+6Awq
JMvMA/7RDfcGrczc9dsiOUQR+i37dn4LxKs7VIJnQSodIgrwODpg9Q5eSGw9APiu
axZ4paLoKyO/0NKhfughuNu2WbrnbUlRhagsExwZFOHVKB+sfJK1OgD2jrwwybfT
R+1TrTBaMRIShpO6dtTVf01xs7Ifk7/pEViFN0081hvi70TAS6RuIn8QWVS6HUMf
lSPzKaqZ5g5Y02/NM/Gk8O0BTejYKpxaSlq4Not7LPV7iLO6nfaD2d7Cq+cDKafm
dj6zJMFgBzQYdwFcYXweKVZgz17SQIG5ikC1+91uyx8jmbVxrD87PeWS88dwQldI
yheR9JrItTP9DnAJkrdz7MgZFOniRkXOTfa6uM7OFGYzlxIaO8mGlxrhmAJw9NBN
D2retwfGkshn4uxahFIqEGZ5BMnyy6VfaWKsfcKG8qLUZJLUjZNtTlWQsYz159vg
JH0rPCIM4yoXChKLdue4GFTn7K/pwxgQkSWRZGrHeYcmpiboi5cXop5/TR/2OpH3
WOTWkIr3IFP6ZDrmanp22cJiBDXJltwj+6yWhTQqtXvhPNhDpGnI3sBI1Km0V0zJ
NDkghoUrrJ8DEKP3krilNZkafVFCCQcoaxy+ecVRTAtQNXEFwQ9wJf5m4BW8uNyr
Z1iU1l77nFwXFrinKn/OVz4E/I3vyzIq3iCnxkHKiv2TPBlKJfIbfIXbGifm367v
0aqDUCYrMAV4YpABqlwrNxN53IcYuMdaem4pym6sZjbZdzMcJmW+e+F1JIy9R6jb
Xh1juH5Q8fFXCuFtTv47+HsGxydcTzSpzFDLJJ4r29fuvMxGYQq43AYUPDPylWwG
x8/0xz78+ahj9A9apsRxujQT4lCUAVp7GeJWDo1Tj3WYsjHfVqti/EpVnclPC3/7
l7T3FAw6VKQtcDzb4MC9bdI6AqwkjO41UBWBfZIgU+YtRn38Bl4Q8tdn3tUBuwvy
FXG8i8gI9o/IF+ofFmQmLYB14IyQP0JjbYOb5+iLy75Rv8BX3n4nBbvQlk6Wx0Q5
t+vqGRb9EXgC47xru7exffNFj4duKEyPwfWIfOxwqkbT1xo1nOc9aGkNTZShcjxR
vBuJQGUFQDUWvdP1qyj4ybS9E1jk7WUdt6Wyx9feOi577Hi2ayscH5sA3Gh127xA
uGJPk/he1hPSkM2J3SKYmuHPuUL2u2VY54KFJhbNQ8MQ1Dwx+Fbl5ZyfBhSPBNjA
f32GfLhgWeLP/PAi0+FUaF3NzRdj9/Eam6mIBnMkM7jsPuMnQe6O36ej4jS3RXVU
l51bvapdVSQGBiL36Tguh0DIHfzB43mMgFfC689/7HkqbRRNjFMlXh9PO9rFnTm/
tznCkemme755Gu/O8xFKd7i93T8otG/aYHgA5KDeWHTjIpl/3wQUmRtpRS4dlx06
SKvqALWhfXz4NLmGXm/wGPhZd4osDfT1eOl42uLVKaOl/lmJ247JpsOJfh7CjQt6
v+I1GrjPNyvkZPSmin2Uh+pmWwvnzYgDmw7KFxvl9itRbeZHiQUNFgSFgCa8jJQy
AD97wUgELSubMCME+2qEaAFYbohb0UemuW6xjEdQYC6vU4VOYQOpLuIoGMucQ3t3
rHDOcjO1mG9h1nAICi7qeGrl+2kWDu3eLR6gtDIIYcrWZlA1oA6ssXM/sBBDqX/m
vPYZp7f47g/cEyW0vHyQ0SPZGivASg9EWl25f22caSIjMQlT8e0yiKO8/tlN2aY7
LGSRt1RNq6iTpPAG2JEvaYguxR6CRjB9rlYRKC/nVf3VF9BxWMK4foBKyfgiJ97s
fk1c7twDfGeunE7t0pM0ZI7N8P2mhMgGt9V2iYZ8ULBBAf9cC9r+SYRK+CYpgQ5e
nqFEg3aIFwquj1ryqrYIusEXE9E6gcEUzp+dkZcvs1uTp+x9R+0m6G2UEgPHU48U
sjMqElQ1PlbGaqvctEB6AAx7JxVxQw8NLqBCloerXMnwnowF8519suJ2GlfVAMA4
+xD39C0ush/qDq5IciL51adU6ZbroX2okiGo6kYVQbtkWPhpZ6VlA2DZ1oYf9zYB
TjtnD8bliqBrXlPkulrfFaJSlSv4TfPVrVyXvUbvvO5NdZ62r+oSGidUFbX3XrCs
YREmcSmlWcXAklBYpvN6tXDUilfIq7PuuFettFoL8OsbR38CsL+aIBHnE0CLhtyO
2VI7heTZ9zIHLHP/IXn3UGud4BMe3Uibgw9Hd1UsVFdGft+xW/k1uJre8PTlNLB+
8FwP+7d6yqJ7vz7n/ApK5zjiwrDNnZnkEwxbnmXaAnW9rb3qyOX5XcyZOSGi5wyx
0coeT7PzPjH4Dr5+gZmcX9Vv+crSXEVTNR86R7GOvIudWtOmSnHQ8RgZa/vLh/i6
fw6dmBR/OjtXoPpS0CbD9GJ1hr7SFX8xtWcf/y+tLKPdJx980+fE6VASlvKsgM2I
t/InTcHCFNfDVJb2AUFEFNddU/WVcu0ngdC4370qh8Byo9G+FjYdpfXWd1DXWnaA
6YW/1crSwVV5+9kDXuBzSb7yZ7KuSBW87WBeFSlppDtSxDiLMW8zpdS7rb1SGG81
5+LtpLptDa+l4SSdoWL2tdqmxOQtBevHVjuGYU4OBZh7070UUbWvAtcHRTrewkp5
TzfgtyxWbvfHCTfgQFzFZvJu+BWhZqHEK+pi0nvbTE8yNcy+fjk+UbFhNjIPunup
YfSQ29l4LfiZ92zKm0qKWXXuWkGSABtCRLJSs2/K3hzOgOfJmK7vzGrgTVztNTyA
ihCIXPF/WhPxHWtjK2a+f/jXaExu+ZNGRNpc4Kpr4p3hX6IDPetrwA8yIzDUH0f1
SwZ7dp4DRFLJzcXAXAjQrHemHh7uVZYZXp4k527Pr12oQ4XKtQcOo3I4+elDDxpF
nzlbrGkcXSPPeTafzPl8/Cbur8GVx+mAIDNA8MSB0UrY9T5ahqoZwIcUP+dC+kB3
GrO00VewMJsGgIw0EVJmYrTQMiUG5t+5cjyzKh9IzG1OCm+6oiU6MZ9KBxKjhqJU
kkWWXSXOlxzBPMvPkJl36xVlwkS+aC9d6ORi+Mx8F+2aLbFHjsYlWel4cZO9G5us
DTw9Z3MFzfL0PTmALMvyYyjRuYv21XUc3KFsq58bDRFF6gTS0dMDu2ektLYJ4ioE
eFQlChxEf0L7tEghyOtMfMBYUAr56udj3Fkn3Ina/iuGYMhefW0mxC822cHMR72U
QrlMA0FyVUpGFEEnOYNwkWmKcvsqp9foXJtFvCt6D+Zvz33n1CoV73EHGne2/56z
tEr68Jd/UZ8b1Tt8uN1FDkSkbKH+mmNzRai6WdyeRGCtyf5Dbxtb5ESfS41FlUqE
T1fhg/TcpzB3nLcz6I+6kMz2+82KRLmV0FGAJaCaGSwtu3MS3iireD9fWtyI3mpy
O0pSn9yhPsBotuSBVBVCvVgB4w1XqDDQmnaPYIDC0g4j5fGu6fcoVaEP9XiyiHs9
PdLYTlOtHmCzDaEtr/HankEPb0HCiLHruGJ4jkGuwVBbksRExO0+gYGt27SzFL71
l7Pn1kU+pU626SSp39TsSjfNph765s0/d3q6VZTc957vVNDt4/vBSPwdHsXiiZkf
pfvizn1pvfP1I7HEYksXSFZAdhC/2tms/Z1xUGn4Pdlx78OMinpkFeC75ZfTr/JS
s2kcguIVOzPPSm//PBLqw/IT6fTv4q6lTJ1j6UjcxscfrGrTOyCg+y+JuTnCinnj
n0rn0eNB0Ftb9aZAp/msPs+w3CxvXCuBqsK2Q9EGXGNzQ+LFJ2XZv2zBey3sw2UB
7I3RksxxS8ITEezBebnEsb+O32PjnrdD6zOtFXR4sznWzlkmedCaKMSxAWbOsVGr
Ebj8GQorUHommt/2xsq5CcmZFnGEGzDyLGU3FQLurYy26zJHyyay5I48APPeSl5I
3XZZ34FZQIS26GlH8tXHmmTFIYIldor4EA5TGrAJFdtqqo+ufi0U7D14uzqZcS19
nArBi0iPZ3Nd8vemQhbuVZZgVlW0v9SfWODaWqbGXudBSIYdSMrUl/4XNzGNR2pY
BDo3mfUlUS0BhB8faDiJTjkgO91yX8/6UADWn3vS8r7iodpnTBxgRS+A+ORTAlvk
1agxJlfIDeQ3JNDquIcwutqiOsm1vEl1LpZOjs7nVO/ljgdKojiihRRKHucidMXA
pE73pIDPVzHaThPdCGR1+KZXB7s4iuA2nyzvo3W0WAqE6WZ50WMFb735QZUUBgRu
xJMZlwwcSSpJEokHYYLe4p6jYvP0rWCaa37pww5RCTv5OJPuqYTXsjMm3rgtpA7w
B6fgnfP2G1IvF8cczC/zs2XcskVymdARrl+P9ykcgg/GXedJFX9vUj+rlXFRjVwi
vMeOoBPpRQWxFYWGaamlZ+Yfgco0NxourkhQ7437rYYwwAIExxvLZzX3wnkFo/cy
kjqBg/cdK/uRzn/0yH7BRGmGZ1lNSPpujCq4flSTSga5tVW052Pelfh5ON7qzR0b
PyktzsuBB8jo62IbEb0fKWzX6i2KW4efIs8yeB6XXNYWR7DrHBo+oj+B6QenacN2
UUq0QCCf0u6whUPIs1uwW19H/h6RMzNFZk8GgtttnDzu7olXIsYVVDePoAUeyx8n
1k9EfB6ApZDy/ddJYWnAI53rscxvKss5PlPcOOaLdjbpZUhhjaHtBK+8UJrIlDsF
hsQ1Mm9aavH4inAzZiZE5nAzszFuFjqixf4LK/9PMyUrq8UqD1FVtRmAZdeemhqQ
AIFm+RrKtThxKtItY96aBIbOlZFYGg1hJc2G0MP4NhZe4ITiXEF5Ks4Tvc4xuYDT
oKTf4CgXc19c76ilw910khdIk6Qs49QzjspKBSz+2hd6FnsYQum9djaVgwzJR2m6
iMffaTxc7KjFN1A7rNNp9IqL06q7lXJt0QY0UEudiTZOOXH/Lzb+7TgX0kNonDX2
ChE2Z8xijH3TkMtGpj0OcItHVCSvMQrqwhyDmiW4sqofqclcCX5N+c/8FnfYve5o
WnjdPreyuB6Sm8FH/hIlW8tCyXXWa3AyCM9w3Oahlv5CoTlt2XcLhd54cozrLvS9
+MNb9BYrMaCFS/YHhPVyJ28Gn9hswhmszkbcJ5czpRw1uHdYtx4y5vmS5OAey4ML
sA7aP2oNJQz03J2bhQCWO2RJeuaxO9YzEe+dZQiF+e59a4DuHMhtovST/ajjuUQx
TkTIh3GU4ICftrXeIsTzbcEm6a3+lm6gu2/0iNGGO/JNh02ti5AAqOA8ULnOdELx
lJUpcRD4L4jrOTQv3WQ4a+2dsuwUm81GgYsPxgcyqIwj/4MKXMNls6E7P4J7Bn/o
BDIrtWSBvNQnADbDVEh24KKCBKoXq7GnMNn5G65WSd5CmdpA3yEfvSxL5a3E+iCd
bknT8HuoIjVRni1UbATXIb2rY3sN4CqMwBTK+ga5Gigy8kH4TaNajmhFYW2bSCoh
aeEMlswRorTtSDK/5pbU8nH09vmIRmlIY3AA8yFQ403DLRvHanY4FgBuhLFjRY3k
yqPS4noifmxL4NruxBIwrRpyB+LT1xGVUeMla12K4CidIGK3GNOdrATA/bS9CC+u
MCHNlBqpWcYUq2KdRnpHdj/JjlSVZPWKeSoX+qjArH6m3ALEmhBka3kN77SK5/Pe
gyd2s4hV6yEPEcYTL5sZCXAr+chnqkzjzH1HnPe6qpVtKPH7e261pOD96TGVsFwF
s03hSUArJXPSQ4loBduNj9SGnp0KctJSNFa9iI3Z1vk+epVqOziFIwD03S32n7r0
DAvx+sWc/5Tj6iTFRwQa67LhByHrUNY8lcVfvTbjzuWFRcuq6I2N+9cN1+mP6OFC
dTWXtaJtDjjSMWgRCD4wuNcIL+rFHR2xEAjOZCSfwkOxIQ7Z+uEzOWAW0Nb6FdCt
1TOx5lNZrJtA92ihUBanx7ALZrcc/HZVM7Hz5L7QLPrkZieszaM1YznjXmV189Uw
X6rr66Pd2yK/8tS+3Ihpd++OKX8BFqNbD8dmYsdqLwyWygtSUoUbWkS9VoDkg8yC
On++Jrvr0HxhpnTrx6iPxFJCR17ZtfwAvdU4V2Tin6oQvsIIIkYftOasuO0pBsrU
HdZrsnrcozccrQQcwUQvRKaSZBj6A7X6AC15FoDIfEcGNd/QX+fZScvV1Qeyn6kh
MCiJC/jEWUUKsi7fcZe18ArVsrEq11I9v05NFz17ydub83L+R/eTpEvm8EQtaayk
EGARjlBB0267zZEqvdAAVzEzIl8FicA6JLzuc3VXeKWxQhyO2yTDN6+siYmanjVe
rh5SiMPlxy+FxQ5gTm5xFJraad9PcFAurrNHPc4uWjoltNUr28kHdZ/1MkJIkqAb
ZcxAIyMzNHd8aopIzLAiyHuM9ZnhJCiKN4LVcLYt3RZ2mJ91ia4LqADWcUFnBFJQ
xlKfpHZuimEXe10uElYRWq7EjTumxThcjUN2Vf0EXaMotZYKmBSqMXv8yHqZEJJq
rrOol7D3wq1buUhpCQjHMg7396LLtGPtCIQPg8ZR3C7Ya6gTgzrdemq+sZRFtthH
9liCea3iC7m7zoLWyiJ2UlrAt8peruM/t9iUzNE2GoxNFKisWTDH4L+QUR7Bl5Zn
TBmgk/EMXvIjDA36chlft0jqt7TaDh+aM2HlAtICM2ekvghq4kZp+KVt0yF6KrWK
kZH9xO5MF2k13Se0ycIaFO2M5rSNNLtM2ci6DyREoMGXc0nawSj1/bJkgMiaF8dC
LwdfS+N5H8fdQK32/OhLAyV8KjRDZO1wNRHEATHpOgZSfJf/2b/AjKPxnTCqKlKZ
q/mxiQQij8eHCUxQkMvYwQzV9GPwsAn95yQJ0zTUFr4tu9tLiMGBe8TayNTxn8Hc
Mp5Lsg/xnvfMa+UxWluke/dp10Tkg5wXMxwE5PycVq3xStJzpLY2PrPIFmX23iRM
eDtvf9yOMJwjEg9AB97w94qQU8q8aCMS+GhiNpIyz1WKmNCIjPYclUJ8z8ebh0NV
cmgSroIkqBR36vlmB/i8W4yxYpHLFGWBkfLm9/Ic5nYGPiF0f9Dl+pPRRZgFCjuJ
hN5FQRhlyj4rAScgGEzrEUejG2dZNC654qRRu5W8K4WB2pxPJUzsuTNfQpL5Hv/j
vcHZPU5NA1VR1SfnLkSpL9UtZsDzk3wbyoeN+hhINzLmHWvNKAcG369hsFDWmX5B
SM+3eSWiGXd7F3/TPzleh2Pqn5I+CJqAObf+kfH+lKfeWMfVyVzdBAOLN6/e6aoH
Vdt4DmDEvz+dDpd/hzpK3nQnvnJDuhOF+EQqmXFYSkp4aVsUY8LNtZMOK0G+eiH+
IuOPu6pGdFAphSLIti1RPdfu1qOGnxEVMJi+W+iMbFYJS7SRv0+k+XI+qXTZZfd+
olYMrYIENAZDyjYJv3ScrjM3Hwh4Ht/1cs6TRudXND4idUriBsh4Q91HIzQr5flN
bdAJG9KsmD4jN7bHOnJfFYf35doeplEwBcBgmeSM8jZMvl3g5pdbQLqF5Qxa2xFT
1eFdmCKVyfm0gA6W2KZcXHdWuZTJX33STKVRAgK9BrBLa/ntOeYU4UNPjrJWAhrY
qADrz4tz7H2GJEYlG0QzRk86KgsS0U4Qux8rBzCXA+IgmTyNtfFG00DbBiMNgT3m
b6NVD1b91R2zsXGFRHaS9mkiMkzgOzfkZg9j+ruo51ypUWGZGUq7rnoYGWHYU/4a
FjDwJwp3cLQ/6SqJi+wZbteAmvyjl4CVIqRvKSp+2Es434OPRe6OotdV13FhfqnS
bqzvIpfvcpKpPK6mMZ4Y5wux+4D37f9FRZELEUwUBc86JzrRO7LDHLoYtDl4ejuQ
fO1prMjKLKcXfyQ+rBZP7+DHC6cfKkGTEXn8fQat7bjZKKD9pdyE4dtaoR/J6A8I
nWt8SHirnNZiYbhulVMezH4lnoiOH8PbNXT3gI69MvAlbB6bcn5L2oRovYwg5PKg
t5sX/ZlkQTDhz4ksobtFcS5m8V4uv2LLv0FeBq0KzIzWxlN24PyG00kwKtAx0xBc
/HxalQOhaTEWObyBaSLup1JZjk/010sb1ka5aE64aLpdi81EP2hdJhM4zDeFqU9P
+vxlZTWMAGBoLJWm4d+36ytWmK64X811D8V8VJ3sOOemynMda7KrPggY4QgeDveL
+wdAXZ0819iguuI/XFK8ULTLLNofYNddTxA37ZaG/0LbzUIBt9jqMMA/e8po2EZ8
0aZKHGUOW7EmUXjM5tUOxQdZ/43NkyOOo+Hlb1cZEQ3MKh2Zi4BWrPkPEV2D14tB
wLJWMe9JGGUWcMFHXFACzNuYvegoL/Z8fUvc9R8NuirnrLk6xYpu8wS7TXZglaAh
ERG8gdIpyLDgd8E/6iZ/JJtFp8NNdqZ3jzqZB/xKQUirCMTCN2Dkfy5KT9gLBzvB
+UZh03u2Z3YECtpLC54GhMX8Uu74p4wFYTI6sfolTOlMnH6U2xkhqz5PpP/LaP7z
czOnk94PUflmWxDwhrhMF3eGVnO4GazUbm5it06qniw20YTYYyvUC88gpp52VkEK
Ho7ZVs/rJpYhwkfip662ebgb1v0mP6iesZ5cxLBDBwYPgBPlygdN0quqaFwlXhR2
sL1gs5IywCx6BWADw3Nl4wH6t5+MKf0Zodhk2lDR0byDqBzs1Kh0zKAnOEhbGVPE
hycyUqQlbDhXv3nCirO6io2vuIAIOmqMEc/Hns5DED5W1/aEwIbNGmwKUGZE7YVN
AW4VjsEboVw0F331A+2wPuAwgjz4Wz9+F6g6lD+1Lal5jNn/6XD1K5ut5Kl4otRt
1Hm7mDcnXrF8NSWsCgrVPxJ9YBsyCBnnar4dcnu7V/67Nedazx1nAGd0PnB2so/g
R3v8mcTLMFLIfx7KVwrgBDq7K1ik8Nv75NLkhynN6YSxF5D4gYy4ViwQ6XZAwFeD
9epQMZsaJqnSzdqN8KwkmhlaBRjrMTNP8b8ZUdUknVASm2NF5HRAOnVjWLC6XAwf
DRwYHRwa356qQdffdPabRpVH7G5SSZO5Dr3izGNg2uTHdAACHvJZMahTsxHAvVY7
dnFoaxknKkfPpJggcBALwkDppXWetMK4qJ7ACq1FDi/a4kf3uFhSghJacJ+e2lsH
GqVsCqzie7sRgKvfvf4WelKeuQkzQrGR98ssYqzWBfVmxUJ3Z7K1PZIIRJUfpYEC
GwpbyaA/mRLR3rKy2PbmKs3H+QYJydSNxGunR0PahbnfAY7w82Lf3REmLmEaYNCt
jIKNsG7cWIQ/hJtxDcA+ZELhtDX3G7s68Qc8oZIYtZCtgKnS3eJV6MAy4UhSAzKs
sgfTC2FRN4CSCDtqPQzb9EzKNbaEI3MKcfNOpCl5WkxfY7Sk0oLoK1isUJcZHSgU
CA6xYMEy3XKfbX2ZvBn8ZE1NSV0s0gpyz9/LIReSXbSbvGkoduEZzATXW/mJKpOj
ldmsg4CxRTX2tq1hjalYitOokeQD6mHHYi9rlUe3sNp3+Qapu9JJm2j/gMIoNpEM
uwsTHgd8eB5cIfXNMUbVkieMDHmT/NzkQ35nJfHEB3IfdBKDEMD391r8dFFPkzCi
VtYuvY9WjOKUoqvTn5QQIZtmM1iVprgwj3UWBZ8TqTOmesbhZMfrH2tut4NPiC4M
IV6WYfFyPHlLP3DOAJaSFfHxLbrEcTDCPbR7MjL89OqY6FOxxrpHTTWQE4AqRJqs
NOLBgoAYlkqILux7GNIJ8hX/qQgdFjhrjZhurKC37oZXnG8rjgDTinNtfkoIBuIr
EfJ+yt/K1y/MBGXYt0rqV6evs/NqLAnBzH0TR2aDntb6QmkzHZz9aBeLOPJcOknE
yY6LYZF3a5JfImuiQPk/pPYdLKLnVR9KL52Vci0O8IRTPxgbpLis8KQh3T8PM0Ey
6EBiUNB0QFa9iOkC61as4XtR74kiY1ARKWV3TJyzMo2CsoCL/yObYFwn4aJqAXu3
w0Z8cOy5HOvPKAWgoyD5WcI4x0SY2IOcM1AU2h3DLmvpT5NdvWaaX332phb3MBuN
G4gubIGMI/y9p94hc09oD3Aje2LwplZw/o4JOmnNby1ruIJv/oOmG4ihl7iu/SFP
YqpBDWmXIGMqmDupROKM8i0FmeZvGInWHLBPalxsv3hB/oZ0KSqFjADF443MsQTa
oLeCSaLsb640imlC8VDNKudyUiTpNsYQWNPgY6Zhn1ZqPGs3VdN3PqJJsTu23ifp
2vuoqu/Nl+ApUQyCmDA5DcV4NWj9p/1Q4b3106+NvmEVgsXsxrZv3XezxaUbML/q
YUOHcjfGJpJRf4p/LOXFvZAOv/XJ3rZPOSX3iGGIl0NjyeSkc9UCPwX0rvosQNac
921x71CcDH6USqKtEl8yChPDEJ9Vnrrut7V38z1Ex8fvWNrZD3QDicp3q6zDBgU1
f12VL4hrDEMw7ECyPLd9Q9p7ECnzi+Uxthl36O2mFxbK5Oku7sHrxa+eo+ldMrvw
T4uVLmypwFEI8uKqat1AjzIVyvwhVZb+cLx8DzvZ4Gt2EVE5NplwxBiUv/0VMXLg
P2RbDNZc+JLJ1UvFuAcoo/JZypKmlrpYCCfZ7hqUqhgi3JXShvhvQVYcKKWVtvVh
Q1fW343AJV17qYMOjKApCi+HjyBxogCqU8IJaPac8rc+3bTwEEs3IsjzFWARlZw2
Z5eq38nZR+NbwMU5wNqgDwFlMbQhUYbZak9kUR1e2I3z7hXOpRNSNfNZaNrqNF3Y
4YWHLHHZ6YB66cgbvLEbncQkDd+PZHSnmkTj/Ok9ZA3/MkyAXmFv/7enq8uerZ4t
I3/JHL1YRGIZZqtVrGQazGffCejczRdNi27pq5RHlsUaC2/ba9rvtPA7G8NoIGA7
ADt08HPED5kEM3dAsFVJv0FQgOQ14WQk7SWI/Dx4lyi0x6DVV9rXqiihtWwjM7tj
hhkx5NYZrePRznTKvegF03KjdGSPdJPtIyxSa/cGkyQ+U8uq5f9Leb6nZs6Kdd9d
rhfytLGgZFfrypvxa3975rlCRjXu/DXbPPEK4kd9Lh9/PEPh7sCa5OlXBXvBxN8o
lAzDoK10i7BI4wDQF1PNMVhbwdrtD47uwoN35QKXkg5QMUT6WadV266OBtMA58FJ
88I1CvyDWJS1rE53RiehztKLqhE3GM1lxWam73Tm7Dac5PbkW5tnz2xYpBB1RYcm
Eh/pOXX52zdCLSNKjLPJQLkGYh0ySNxtYIBFY19CnQprGQQamdyTJsr04etwibPf
wDGiVE7f1ZNzaPcicq6q0q7uSiMxnMO5i+C7grrOQn2K0JVwQ8f48H2Wlux3vXL5
rGokRWmMTr1YBfS9n6IJdH0/qsy4CjS3nQKFWPDR6I+6aPVM55mHW3RpPHyWhBBm
1iJRY3EsyOAR33L6WyxcbtqAkTqEx9WEP6yRmDSYforff19DSz5e4a7VeAH7QnWi
dsvG8GLkzYnqwfooUpJdfJ/jlHR6RCRDastzo9712B46O7C8wq9tUCaSq96atsiU
e4rXlwt/nDqyN98GFSc43olmUm/fRCaIN4iYhdOomUDaTKIF+Nlbo9Kprd5cJN6i
t1B6AkD77GiqkqR/6vX8zX3n3Lv4UY0SCCZ7umD1UyELdQOSE5xND3oXt7xbHPky
HZMIyBdh037dtA8z91m2AXjBsY10z6TnJg810qLNYTpTad6Y/kBeqHruc2cxJ6EV
oyA2TVQ+r2G5wGNefRHOE4LFlQO4mPdzvOtOrKELwjKy3+Nn7pJEJalXNw8UTZ/8
to3xW5G0ysKaAAhD4DiVU1Y16PKqEvusZ/PxQCad/ab4CNzsJAXw5RC2s6xZgp8W
QXmnwma+iF2JL21dcseDF0qYAUmh+mSTaoBlDuFWoR8AXgOVpmGmONhKZwEgbnjU
eCxPbWy7JLB9EXz+0HeryQK9eRemb82jqPQHzQXHd4ufqgJFbEt1dfLuIjkuyXok
S6yjU0XRkq+oRXWjzb+N+R04wvwx+l3tNk8rnwFmH8eNyDRV1pKutHaqw0qFhwgs
jrxUBgqpz3mFVwwmYQOjZWy6SnaqPW/v2HhX7VVux82XlDrPuFl8VOgOXB583Bn3
ceT3/IpL8r1VattvjjrXEhoNukia49MfMk9V0wjpvZkQqFyYEl0GukRPt1H8nGT/
xMLGmF3UOOa7yqqVQJmQEdetcry2Nfb3JAmlOR0eRYsvdZYp41cHWuSDAJbr41mU
zpNnnYhtwBCRdSrocqWEJh+6hxNaZbjBo16vhRZWtZbZSpIpnBj/J+jSVpzvLhYc
WrDwXCJtTrAocuJxynHGP/T6UyGV0izMkFTkeJctvz6RXAprEe+ktvT/EGK0Ie6d
CBBf/QfJIlXPJLChLdaRpeHo7R/7hJmugOg9R7vAXugGOlYkk/uIP+AOhCvgQvl4
tjmAPKmBdyIcZfyGWodwvRd3BckNX0+PR66z6sD0lNnhY746izf6fQhHc3d9wRqE
8/AregNC/QPZhNI8m4SX00KUFfQ399aAGnCr845ZYhsZKLjZZ7k1uMziFCfKdKhx
xcYJV5cjg6z4ckR3MqoT3zq4FNr99v20kOrmxkSYCEhUHy1RwP+/X6i3KykNVZjR
94DzxzaX7QWSndHt29iZm1X+2jdxi9YvjvzLpg1bZJjCIjTFC6kKib5Qc2Zi9+WY
vhspUEBAXxx8EFEIZvkVy4Ph7R25ttn7qq/0AZkVkhhIDwsakcTiNPg/D5fmLr7C
MW7vDxLnCCRLDx5eksW1ba7LBE1QKI9/oSlCP1hu2G+kO32QnH6a3eXXTf1GDxtE
J9i2xM2VIlfgQ6406X1mAh54F5GCMavZgPCkk42fj3DU4tNw6Zn+uuJq26CFa/uk
zQieA+mh3a8SMoHb8JmRTP5OgWn0yChrqUmUFwKBpzp3OsuovHjvdyJdJuPihvY+
rMwOl+qVfsqk6ovjXy+12xEHnfr5IhPoJiC4QXBJbSMUnhrMl0O3LphqdLaTysRj
XJfVkliDk8z2BQ9aj3cGcNWIiTX1yN8u7CWOvKxVGXNXhPGtPxD3+mZmaGmipYwM
/AFo+4vldZwQLrNzYxpzMzDQDBwdHit1EIWsMMnw9b2cYY2xxFGF+e6s/boHaGOY
HRRIUt9jW/nIhl5RpZI0nYb6xHwZERybdv8VsPXqsXgGyorJ7iSD1aDazfjWDdZy
T0u4uoAOnWjCXfceOVYPp3K6c1d6MKaQQ8YpdckWbBhPCYej0tlErAqscMCIye8t
kFnbpSM+7yMP3pLxanZFKoLUg/TkHh+ah4WvmuRkdu4QWZwAOPI/AEqbgyCrqgGA
pIbgyGz3jtiqy5PFoMp8duG1XNhkqdFNf/F2Z/J63brGckg5c63Cc6Y1dsniqawi
s1B5/ASn/VP6JL7XBNKqSzp932nOYQNgPjpuhU1WF0T01WNaA6Hz1bLOEHshm7UT
eUjy7MgTSjha4Pw1Zw6h/miaJoPQRVppX6Gt9MlYq4vFHPa08cUQAf+MPhsbCY7r
mjEul5QChFXdTCyzZWNpz21Bbn+sXIp9pb/eD3BXbmtMoXITsQ1h0Lhh/M3Az6eL
jQz8r2mTVg7inPXtngwyXD9HzJDRuIVPFgy8ITiWFfDsZtFM38yCTv4mzES3DG71
sgmGvMeE3Qhg+sNEFqrjelz5v2hbGIXQ8FORG6ezcnVcq2iXhGdMqUePwZdsKof3
oG/IS/HeUFlMvjIaCUHcnQobhy+qPMMaQg1F29SN2fHyTlLLWGEGk2lpgYJLe9bH
AKhHdMJeypkzfCxcxw+Uqpp4Qht4X8PC4k2znRdnfEPQjh76XiD+gBRqBVYqn+KJ
b5vHPYKPaIRUTEjtijWoCq1Vq1Auc5xe/VUIxD434PP1KPliqxEYQmAHzrRjlOUh
uo29WMtJEHhQf40rkLeDsupV3BYN6mizeyd5O2VRaUTBV3C/0NISEBDuS6f6dxYh
G2ltlkwDhWrWhH/fRK5mrQeMQI98kLbShz2k4/TLB3fyXeHRYMxRPqG7KaRXy0ps
n+hHWIh6BqhdnBxb81k+oBNESF9KNqbaFXrY2wOni4ef5It8q3RRUWxvjYEDK67a
zZLf2+NS2V9DbMrUTTZzee1lKMfBEJy3WVV93jNP9iKBh1t2RBsMKzIOwSTSmHIg
T1/GGAgjTdvIfKF9s/3TnrkR6vi6qMZUWGR2ItgBT7fRozM+Z/ouTVR+Hgwvis/P
SJKwsiP2qR+WfbKqUsTVTWLtvyYdvIE6C0ejWFB4zG79e4t0BGUPKlQCy0ObaH4a
3i9ovUTYj6T4ycEWEVHPUpAXAyEbw61ccLA0/V9nBQIcLAfv7Rl+N1RIOzeL3QJn
z0OCfJSQuJkPjS+BPbhOvTC1hBp4ZMS843S2e+pVpI0d5jw/GCz1cqkQuEEbUBpS
yZJMDcK+7dut8Ag4hJLNnNLX7/bOVemEeYCbvMQFrmHhLRYJ/mssRbMH6KKGl8/0
AZMTNDSn5YyKgSvluU1sVAHGetA/7b+Lqw6AO0jfbfWHFMD1xKEKYJ1b1mAAOKEU
hUfRotS7/VUqqu8e+ZjHU81IY1pEfH00vKDpIc9iEfncuWvBHZ33xqaGXb8uBROJ
bXPlQt9zr5oFsIczb8T4u/zEXTRcqUBJVlIrbwQnA7cIvRK+JJqVbekt5RvQ63/H
K9NX6HTNcTvK+0TR3E27jCXIgTm6kouQOMVpimFOWtcvkayhmJp+4h4e5ner4p0J
/4oIzA5UHUN1eWI3dvf9bavFYq5u4l78Jgnz+ftG0RDFPkhkD6fCVRxt3DYurmgR
D7ru10NSvRR9zCw6fHqq1Mc5v7YJykvl/mXH6UZVZzKr2MfD+5rapaa/pwwRF1+X
XPVOmJMeZPNyto/4m6MD6c+mHItR7G+lPIK8BMsUPgJk8NMpdUnq3vCe5HAVyDzo
juBoLJS4bwHBLfYyIWDB2CTkG6hij7OtnSrgT3tXIgqT+TIlDWVthyyVmqVS+HMV
rSYF9rlt18+DkQmjmnUgySNrjHZ+nn+MxeNFYdgS/LFQ0BwKhXPLvXWWLD1cvqJG
eOa/LPLjOQDN8UuqAWWCa+QRU7daAhRg6n0JEjdmr8VdFzrLRWcAOymyqk1/sk/9
TbWd0PAtLbtkJlTuI+Emg45OPZnvHQ125g2khcu0a9GPIaL3hh785yAN78hgzUZf
MYj3L180b8zn3UzNAQ+63t18YTff7/fjdTgDEVvqNmQ2SUhkwYkF659B6B4kd4V2
YNJ/WoRPXDUPfcbTfO3AG3asR55pdFvaxnVBxBA4IberA6UJ4/on9YYypyC5JYxo
SzarilCY3WI39RFj25iyOKzVEWnxJc9/CVBaC59edy8m3cTB+SrkW0fVtx8WOb2S
HEA5WwXpzAIDT9sthH90z88wXl/NlOS5Ljqh+FFLMW+YTqaYeAuhY5fnD3d3eBM4
bKoIXpHP5+sVnrgsksQMunhiQzLS0fWhUWw9/llRE85BBlj8tLuuodKNCwO6lxco
cG9hfIwo4yxk+LxhXIMgzWvFFnp+dimcjksS7atG1VEe8LpNO5kqinUiHDBSx4LG
wCDH3HbQFCEuvCCOEYaBLQR77uisbsOUZuznKRFjbbD/D8eYpqN37/qei8KEe8Px
XVB/T1zUe7LEKSVAJ8PFc7KMNMztS4ZzWFEJC/4fk/6tO62K+d528sO765zdnKD9
7maGSOVikL1xrAZMA9TmcbZLpRs+yfWzytehNR90Wg4gxeJT19/zeI5YfKgc85+J
tPmnUhRtOPTAdyJUCbdEYu4iUbOlcu1vR1BgLc/7fJ248z4/2aTJNBblIRa6pu8I
E7Gx6Ca6B0e88sqQ1LZLzeEOewYp1Euwt4419EJ0mhKtsohuoWBpzKnbucyAZd4/
Ud2j6/NE3pq8CUubTVTciN5sWedysu1fbtvPP/SR15i6T5Lyw6Ka4fEApFnf/EzL
ylTTU0mXJc2G7tYGtgglAwwBiaqTU3KsnHilHLuisNgdOAoweZuanjwjjFqSNdB8
SaIczYWSYXZAzbjfBRyNL42s1FrImuexYixfquFeatxapGKqBxcT2Fl7zVPkZztx
QegFXbasrJBFi6Zczi2gxXex9ZLMyj9Rr3xfxH3KN6JoExXoopVMBwBWKZl7mEje
acviYgLOzPHP3wozs/rL/0JLFQdjjAiGv4MFhAZoqfRDDqLJQFglFzFNr2t/CsHb
H7xL/cW/IytRXgpvlI0wt5gWCZmbsTM9CgNrjMfD/wd4jSaUVL6kxG6+S/W8X8Ba
q/SemNQMZFpIDUR21hiImDU26GKNzK8LYK0nt+J1ZESoHX2rLb/IGoY/93Rql4qE
zuAa5Kw/7QpY55T5HIUis04Kp8Wboc2GJDw0mRCbqbuTtkpE06832ncNOVB/torm
sZvRZtpRiSAkRheicSuByrL/WJTS2/sMdgf36HwN9cztw4wzOrEE4F+WSKoN06oE
PRkDK1WO/HKgpbapCwVQ+sDhjbMlBRLvjVHC0cHEsU+UCRG6eF4VFWcH5iXWTJoQ
BdMyRvc1iTvwGYMjoeS6WilP9782Sy5Z3RgR/wmC7A898pS0TCnegoh8KLpaIJTU
JhNnE3tj4r8PxG2qnT7gRpgkD05iWDivXxQbOGIssRWJiUNVgsO/uPMWskGzXXbs
vd6GI2tzPHEn47yRnBF7evfzk0gc6m99964piDwEBJp+gTqsDq29yy7edUcs11n6
M4+Cnd3k9viF84SqGU8BJDJbF/WufpXlCozVkThUEFlmdPTFWZ/udcGWmnxyMrWJ
AG/MUqhrlxHirRyPJcrNdIf+gE7Lc2S6hh6E4jLr+nRiHe0eNL/Fjxoe58a94v0E
QqPBnKzuqLM5lrX3Ipqdfd20P+5aMMJ/iwnpPWRf2ZMD991Tpz3HCd5c27yXafqL
vBz9v9bK7hQVIbewphKqE3uV89TqDOw+9pxZ0mB1xkUalTKDPYC0b8GOm/GWUSdG
/i86SOKpr3Del88GeDNc/xOjZtOeRYvBOHtOBS9fmhWpQG94b7gs0pER/jbQNP+/
olkIId0HK8w+2tNimqbA41zsHj/G1IJ36FTWzH1Q4fo6XXlfCzV4ovMIKE1ALo0A
2UG0YZvqJVkCkoZNgy8JvZqymoU9uGaCdmDt+UEGjIgdANZHa4NqyCgg/wbwxoEO
yEyhUy8ju7CNFxcUVeuX1F6C9IHpntOBn9ulHtFr3Ga7GZqNH9RzBN6qePXFAVsk
9u8wovmD24dIfSAgBaAP57h2/l2SfTTLGtUXq6MG1iF0HwiGpjwhJdMZ1IwFYGUK
xuonVAGkfT34Sckl/0eeL5ol9TDzy5I0jEgMxDvWOAowWoh0s8NjiIX0hCP1gNte
tzivFhSYskOBzamcHdDhSJFJ16OsookcWGCOEhP8kHRLhDIPkOsib5xVVUVRJBLX
9G5/7Bh825x8N8BJghpkedVzjrkE2EUbic0mwUhBQ1ui/xsA0HjIuY8fZ37k1so/
CdvB3YFdCEB7I+bEKE1ERLfkvrRPsMzJzYiw5H4UaoQhQizbUnXF171kxCf8+k1n
OEVj5GEfIr6ar/pnPvy5+UpzPJr6C6K7XuGC2yyYVYcCsnl2C1bBxPkfCrcjNz2M
TvncvLCYcjKYEeJT85HF5pVytx/LNWKbCKYlxnaQg4MiO+xDhJq0i/MpKsc9Tq91
RPc5AGpn1rIdgIZd+8uiIAcbEd3h3cZvUaj7kRlWrmWgYX7VdxErvhXtoimF+gE/
uaJ7bb8oD5dTPczAK0dBSluY33Efng1c3KMSfcXU+YTV51ujYCU+1GT+BuPoILqh
uHkcAWeOu53BcfRn+9W2nulggbr6Ze3THNOKupVNmttb2H8XCZjXVYfOKw+UInD0
ZLyU8vqfRFqzqb0zboKctWo0dz/RWVJjuJMMkq2TMUUQVg9Bg/ZyiRPLfC1YJMRP
cp+4cJCwDruv/AHPd9H5ejfAksMfotpcG+ArAPzi9/UcCzcnQ+sXu631fXmgZ6/8
KD13Mmf/UGSID/HrpcU8aoONIntwn8pnCBzeUprxcIHdJCc4oeEmicbOSRyoceXD
0RKnilUAUnvKm24huxsalRwQURxUP2JPpysg9kRrj68N6dWPapjXazp+oLW0Bsvq
c2/WsftHdVjIaitXQoUG2TuYZNuwEQ9oj5IDRFDihlfLp7CcXNE18sepEzxf9zQ/
z2xiceMtEeFexgXxJquyfEXa6mP8ytYp6IbdnwLghwToQT+U5PYqqRCUjIbhol1A
vheHsbVZceXuoWnZ+R1kzuR82cxX0+v6wLxELyweQ1kaT8XTMhOvwyxnRv+NmXII
356FxKzemJ25Fc2/rc+X1urdruSikxLTYLDe1xPriz2z+3gJaq3w1cMQ1Zd5y3XE
ELKrHjxGolQRVl60Nq5ccJArvVySd5IuG/ReMvyHPI3AvJTyiIPIavWgQg3Kk1sW
X6sz0zrvz85PcG84IxhGKgU9/LfOvV16+ku7MHyfndsOGWLzyJCfkzZcbfIAkval
Go/1AAZvDO8PuaZPlEcJrATpAQgqMR/RKXbop9NjtVDuzfsvpQ5F2OKlbqK0GpTB
1/etv4BDV+uHrY0dN6ySFGI/x0N7fQyMtEItF7/UNQsjRABNAjpQqE8934fgYC86
WjqtesVIfshCKEYSjMnfrQkVvoc0mWHYJsi4rtcevBQMBcpr3/3YzW0eyUSzT3Uf
iqJKiL2hZhABypW/035hCCa+yfS5UAH3oMh3bg4HCqjCr7PtReNDNflhKSpuKMYf
a7Yd4i8wRCOXb6ypIRD3TRlR/sQ6CcwGzryfc6Ri64EL22p/jmyXpH5JGbF6muON
/6mFL60qjtGYcSg+9JSV3fKey8V6vBhyqlryDd45qRT/tb5cD/LquRcM7HC4PD5u
qrQENA6gJU6p9g/Pcc4VI9Sk3q6UvcQbY6oAex3gf99XDd9nY5JmdTqS0BvS+Rs6
w6ySg75YbF+vRKzgUIgeWWx1ct4CmPVOIONpOJxSKrbVdOyZ4V8KWMoC89vJrpJF
ypEVFp9xcq1LM26JU6T2slqBRhjSdhfI6hEYWVFbOs+UxNG+5b3jHNulMaW8iWxe
24sggOenoORbttjFLTxkaNuEIKKxYHEtPRlRABkijZnxPscUnEFSy1jBE8kn4Cby
dlS4oUtx0PrwrJ7e+n5e6Ove9lfSIdtTCxPtkhriB4s1hkJR6disOxod1nxUb0+W
fWSkw5jgyF7p/Ef58KaVrJ0wvSQaOYkp1pn6pMVEromb3ppT9dYu5uhZpgNIvznI
cIH3d+Yr10PmGReIqAYuFT2LeZ7deBXrqRo2dF7u+Neb2FPQDAWNWUh7Wk37VpBK
v/OfQxSW3kGd5f9rhmTQ4D+6OHhWYdxkjDdsTK6MEI0IYDNoLJnkbqLnaiB3xM6v
YC9gdSr+Fcef1Sc3RkYFb3NL1i8YsMk/ZD1LlKhc7/2qCzG/31K2+ortE0hMOvoJ
qeJWBYaSyZLU75tU8Ku5afnNgGqWShhqwWpiks+0nYFdLu+G1qAmiUAeRup4dY5v
jwUIoJ6Qhd/aH9vzGBH0Xm60+JIBj33OQvlTac0sIngq6Rv2v/Cg2hd3h15oKvUO
j8g2wSzwyG3QbjX5gMvwrkOFFIw1NW8ZIQ2tFU7hKbepTmIoZr+7rUdzPL62QTZ5
F2XmWqMapKQYJWm8t/dtfk5XSR5P5QVCkB4pi2cbsPLhvNPH5Rjsx3E9sQhp4Ngi
Z/g0mC4Uff8V+9CzCyAr+z251y4nKI0GloTEk8H+UxWHoBqE7txON6sbJlHpAo9E
uZS/Da+iewnYSvMgiUmCcF1i2y/rpQfrWb/mf3ID1wBz9O8uOlKSwe7uML5A/V2Q
9b8/3LP4GLb8Q1dMdOOQjRJNuq2ZaZTn2LmqyL1/iAdrc6RN7ZWjrLZGhY9n4J4p
x+sYo9dPxs0plLOmJZbDTuOs96Z2E9GU676E1caAFgjkEyEas0ulTKhuwFSqlOSe
BQE2Swk3WMpZxx6O5b64luCNX3kmetqomrkh5COhjXNkT/F1uyRjYA5dm44CKTPL
qzgKH7qERcwzRKAxgKOVh8HZd/nM4sXCvVC8+gQXlDHdV98+tX9Rf9oIUqvH4M9z
rYLF4y10puXp+e8S4rYGtr2rTrLQ6Gv4NY7v/xwLdSIPBdhFuxC/6xT0D8onNxBh
LDG7c6VBd104ITbSI5j3dmscpiUiRrEyi6zAdd8vlNDGPoE+8jT3H0Qmv/zOUDPv
/532beWcN50wMhvg4s60hrDgbA52FRsp+kqBihkfK+pJ/MfrD/6hR4HWyRO9I7xC
DcPpSyV7E0y2b+57CQ3bbIakh9OePB53yR5I+V4olJZxSX2NkU+M2DuIbZg/9vGN
1omnkeL4b10cGoXAjH36RHAVp7suS+aKDsH32ev9dUvTxtz8y/s+DlpcaacAYzXa
id0HZiTMRlnI2cqRN5qmIMax4ZyT9TvVMkfxtmd3ExZzEycirFMnBEeVjttXl0iS
EWwvsvSvACaB8noX8BSBnAApKFrbC8uNo3RknHEE9DBdfKQs7aaFysnJZ96ADMD2
qxpVSI+JibOkxBcBvKtR4PUSa+g5MqB1IBg3n51nRmcGoEBJnhyVbC4BIK6L1R6d
wxNdhNgFY0zjrsth3Mk1dCp56tOh7GVfqXeBr59LC8u6/RaqXbHlHMndZ1GchkVh
cRG49vWyK7fKe2xqQx7vXXVTXT7OVzDHXlqFJis6oetKAjEjVEcY6nwz2l17aDwo
uTU9WuPlG4oMey74u1Nh5pyFESzS+hUmo4i1LRfvNIsbv595ZVXVPjxzH3ZpWuaj
1m6Ba1DSu+LRxq/9wzNV99bcTSTO6WQup7eZPhZO3ht18k9pQ9sXgEcO2U74KhgM
es1cbPkBH4+ZsU6kHxE28InnoOqIlrrHjMzY84yuis8knJ/wDQaQX4uwxaC0MB0/
kJi2jc0PNdViZhtb5sMK2g7M/0GtgJTX+93woSsyMDpOzoKFSJlHT3CTwy2oAdwM
0kswoDJq4QHNKAZ4Hfp1kAoz0iDnJwNhfQch8nBd65OPA95ew0VAwKn//FNTGFoF
A01bnO1pisk+dJ3eW/1qUK+7Mka1iwQh0pDqCgTMDALEFyX0X3Syb5UIwLG9HbMv
AeOn6uUOA1azZ4n8kWzASvpV21tM7Ttp5i/KyL8niuSsOs6yRLdNQ0JCYn7nRFzm
be37lZiew6uwkgV41A0QUup24f2lPuekQGLXkVSSKxx3RuCXNqwtVhScoN7W/ftf
rA3S/qwoWNP7K0t5WKbocJ/xrp6wM3wd5Mw+nyBECoCfEYz0EPOCHexuEDWTSJ/v
kzAMBHsHMU/awM9xPw3ZCvXxdahsHIl3zvYSr4ugZBEAAFcVR6qw+UWJivC1xpKs
d2ArfsHcLMJloNXtKfMhgj1pcVdNgLc2soMKo4Wgg6HgHI4RaxOjLpUkC57m+cVK
zQRheH2L1IKm0OAqFCs7FWtLIHoVKPiX5GzF55XROeujeFj16zH+B6lTpuN3OWmY
1PIOeNYA7mt2Lk7J/UF3njGysjzyWMPJQ6XZr8eDdtrMUzpMZa183mZO4Vab3RV5
71TKd8gUbHyXlfpEpmNhRBD7B+sRrEDFf/UVRpKfEZpuO2AoVF4pGOkHPiTWZoUC
ghKILvlzOWf5gzSGhxpZkx/IYzp2W1zSYXZMZKyqgyhjb2LHTemkwPRZwI3cV2ff
U4nqLVj/ya52Wo0wIB+h6h8sDp8t4+eqrnnkZMKH1lZcSirjyz2qECeBlgZGH1rF
SttGqU6z4eDdrqr7KqBimFqLRj73H+xKtcdjVB4vpS7kVO4cR43e6cyMiD0Drpxe
AOyhkJGQkIzDrDYjFAFv9Ll2xPaq4E0WeaF4pLHB99m2ZtufDN1kYembfBzmqsBe
mZ7ZyphwqsPHcl5KG5g9hi0Fxsnh2RFHwQkQCvzmD9QqNEVSCxp60a0kYw1afMby
DuMw+Oagavt5alDM7zbiSG3SArbbvC3PBeR6MRG0x4RonfMw6rUFucUcHnV2sleV
6hOp0fLxuWkAJ6Q5PlSUFlyYjmVEeJBMWjnZCg2HZxhwxbCLp2a34Zq7FqOWAHKw
EX/LTDp6uR+1bvYGKzoXFt/ho9ya9jbQgufimU8xFylwtEdS6y27sGwcUSeOLiOi
6Btq7O/gXC+0QnuFjF75LoFS7dlaVpeCDlHqNic+LrYQat8uEBe52Z1lzqXZUqHp
ETd2+vn2QFYug9h4zCnvUlqAcpt/5stWsgigWxZ9D4qbOKHZAtdz/cFlhT0BNlLb
B1lKbqLzTZHzkuziONiHcVD0d2xGo1aXkb5r5fkyhH7YkwMVwQVIcnLkNBlrfw4Z
iaIzMdwgvIAJQkF9T058hC1WVisa8nqypFHG7aY+4v9Epb+bSO83ZDwlcUXJ2fS5
GJpiLk90+bfA0HDA8jmoulPXk0tI3OGEjppghgNFtkghlUBupUSMCr26qVqpTpXk
DYGv8df04dPJmnXYnEcM/F9z61zbyWYTSoFgVAVQ8stOWuzNGQXVXSM/shHBvH6Y
CjG1sMI+7F+Sggsr6K8/rTGbNLYvo1whg/m9ZH7pLwLPFDa74c9EIB7Cf9mwSTrw
aH7+qDhPapE/yVCbxt7zJbX9upWoFQZS1gxl7PeGci/TLXlQ5Icb2E5Wxj+Q5z1u
nvW64o4EUaNyyslLMptb6NaWVG/4809rWUTokY6k0lLsP6BVUU039OkbDDg0sU+v
HC74bUDhwrL2x9umbgpN5T7Xs3ucI6y1ZJ2fqciOkr6rRkQiByWRxbsNrU5f3Mcv
w59UG0Btb2JsbGKN+ytRhmpauRrLEDhwy9V9UuaH8dKr5kfRT6OvA/fQjdYtWTN8
nXE/Yb3OG1YIa9ZKq/HE+ySykvKk653fFn0H6Gx/GhKrdWrz4ZEGqlcfQw+HElZI
XBRkluTyQBZ9RygNbWbVEzFNmVymqBv1osspRfEegl5sKx4rDri3kBXKYHNM8Kkx
5d9PAl0ZNIXLYEuffWN8bXUKSSwJgI7qCqfd688NoIW8ug1SVSQJf3IxLmUgLNXK
FBRa5nC9Xxe/D6sVJvkYTe7fBKFjHuekMQCh8cRaYithmkGx3eDqNPa3EDhubUis
R/RaXzYZVDSfpfZ9WJh1UrVAqC/I6lH7/2+56v+VIgHfuvG5bYnb/Ufdyi267Zgt
qzcrXNeklRszZl6llOqgVWmyFMcOo8qmeNEiqD/xxoaaxufNERUAyNZusEHgcZC9
eIEOpj+208SC0C6GUELcgbjiUttV2FuuetL1Lww4/5zLHRrd3GqhAvFmPELqvufa
FkGxm6V3QBjvAZU4FPMDNyXwp3tGow3y79oBoVct/3SMkBBoGegbzYn1R+VnqxaB
VqvK/aB6hkbgKCc9VxfIZJsSC4q3i8k8dHSoDEuoLKcqS/A02f3lk4wTIH+D/zk5
6x7QfrN63WDIOvarULdofUXCa77TAVrc878r1uXsB+62DXt9SyAJXXzEoGOUXXrf
XV1pO2eIjQ+1wgjsF3oIpAhiARBOgpdKShfnYNyhzWUuYU62zAUBHaSMM2HCBYM/
MSFlfHONPhM0HYCodygrslZeTZevyC2UbnBI2Kh926NCjmwbrr6JBiP1qDow5o3R
i0qhl3ieuaiEeTf4kbLKA1Ku/fyzTzYPTWQuP3w7GNBSfqnU14no8aMh2jMhCH4f
eSepduoION/KdCMQjmHhq8ExNSHu1BOAtmwbQ9D2sbJiYAb/Es/z/3hvuknGTqrZ
VxFIFArW3e4WdL0luA/A1/rj/MgmjyxOAU5rSR3iEsVQOs03ER0CiFExnPx3WnGE
NDrxc8DB4Dfe/6i6MsWqcfURvNvEZWLx9QH5NzkRFbhuQ3rn/WLY5KHJMxwy3tq2
RYKMm5fRF7T1XUw/XnL9s0pj8fzmhcXvDbZz43hrQXz0NJd1y9y7MKCVZZ61NeQ1
GH5B5sqNEiXBKUJu1YSJXUmiD92ZSwjiua/FzdzUJ4oYugBsX+uA8xh2/s95Jk9k
B9Cpviru+oh2y0ssGSqZQxklfk/kZcBNMxq/bmY4X7ZYvAMEgY78/qZ2Ap98s/fI
AIZ46NcgCJifPi+VJxwzYsJw/O8d1UUrcVOYlVa87eXZ3fCrxOpHUD/0lO4s7ogr
IpeW5pipERCS3E+bw4khA+6TpOQOQs65qsGAYzgwXVI3byv9un3qFZvCdiMYAKSQ
R5dAZzXaPFLOixwPVVkOZ3tQklSL94c4fktK7IWW6PPgWy3a/caFXXjNsbMsoOwN
RxNYO0e8U8OMmg58OaUa4or6Jcyx1GkNOjMGAwE1l66Lrndg4jZrv7PBqi1nmwfR
Th26VDuVFo/mpDZHsrEPnSb4kwzZZ0xv5DezOzkvicQJt1dcUMKnsgYvkouxPjd+
vLvLjuJe6zJdJfzgxdVRKjT3PqfN0EREcwASSx44tepgEswXXJJpOX0FjSnzedWY
KBEugGeAk+M6B6ZVviE2/7y9bg66/GFOfpSIZH2mSpdvjjCRjP99vEJJZ4hV7Dy1
iNBIOx0Ix4svOH4xT+PI6dIsRGPap6jDhNBMN/KwZmUy2Ryac9m2A5qItJC/5nII
6rlIjEK90B94fyVEwUJ9TsDkFTGzTgK9lG/GTb3ok7CRz9l7OSwmsHwfOInUhlWR
72ZNXvWTPU4KP+RdzVp+8UtmiTQ99q9zbjtSzVXxbkg2EWiWhZshrmdvbZ3Jb3Vg
7lmQLdYSUYyurvbDdGGqcSIo91jguuYA9M8sBFG6uf4WOTLv/HpnWxm7rUm1UW+2
/bNqJh3/s1i/BKgUCucsFXhZI2uKa2fQ6b1A1thYE4yd4H5u/QSUsMRMeTZcpFDT
V64eyT6zzzPGJq+/OykyQiyzJCK7Y7FBcqtgwOPuBPaXUkgl/B+1shDsGMWFUFty
ZhC2O0jFCFysTDSQ4YBLgymGwvazxqheDMDESjNNUrwH093KV+IEI3DbMjFECWho
rIhikGs4jOXobNNJgT1gNCktAGifn6v6mqhaVmtZmyCZYJVnawEml5HSaYBBiFsw
78fik173MuRCBprUPE1Y+o0kme2RhzSnKjk5qrmIb4kF9Ef/JFTtL9oziwrRywQb
5MLSLVeEaW1zcGl9I8bi+lb1zi3qe0kVBdPtLEKUaDZV9GDNlltxv6BHxAsdKYFy
ZOAyK/WAOn+3lMss0auXixuhraEUHRPfUK8vpWbHPCYa9iXjIy/46Y7vxdZDR/VX
n2dDk5wQZZgG4sz407tgBj6p+YC+SI/E5A7GBpiM8io1hEt8XbOvZEKyagGYIXV5
Z7TaVMU1KBna2L7WccXIJqulL0jVtFV2Y9wRqwDkvVJOxiE2yUO9PMb5IWNdywWC
w1YhOnvpjDNuLykELAmHHRqQsTAbGKax2RHoB1pfbEbfNI75GeLQVn+PSIrPulv3
Jc5nv+TDOGqqb4rfxL9FAowwU9eysDjc9GhhslCMcKEY27Z+m9SfQW7BYOVDA0p4
cglSZFTAeF+Y8PH5JDuBzwAhpcJfaPSopHkstBDcXPGQxGTrmMfn4OXxwMlbHo2y
CzHEpLEPPcfZw1sQIl8QnltCzpOWLSq5LL3fQ4TimZT46l3Rrv/aQFRsHKzX5F51
GWLVlKzIQs0NKMrhwHYk8FdUuwQZXaYsQkRbZKrMSY5EV/EDZgT5DbnrTBhzWx2W
8Qv83g2D/s+UZIK3nlaxTyN/n13PeAwFOT8hGfxQnNFC00qDiAoJhkcdHU7k4dfh
5RvTkVXXtfes2MwM6Exp6NPMFpuHu6oGNmlgEEgwawgOEmK+I2Ik0Bnc0pTbpzPx
5G+e5oRu0hiE8wTY80SepDgunN+5bMhdcKJGXXSCrqkwxbnNIfryHprllu6+pKNb
fMgjxFLPxyOP7yaXX4woVUOWTiLbHs9YU4h9w6hgTUGHDW7Ocgi3Lv5bi/RN/Th/
bUxG5PsMSZP67m8VcyT/fMvLcjOFa4WdCw0FFlrDFP68aklTadJuq/ZyCSK9Ld4t
eyBZU3hQE11YHeP96KfbIPK1lc+3qlvOQP9Hhr3ImADZN2OnHVVDoYs11GkbKcjU
8KN1PhN+iixY89Q1Y5OZgn8VVCTCPTugUxoFYQ825TKFPXIdSyzWaCW0mXx3LInF
1oY35YTe7bYc70PE3BalngMFwys5shqBQ0p4zIO7kFhoLJBlsgnL/9+2Zpf0B2cD
n2bGD6gzXeL53zdx2yfS676WXnBI2vADry14frS5qElze0sbN4+Dd1hvwfcMN9Sh
B3PEz6Wti/86ek9lTqUlTivb7S9UmrcMfTiiVZiIA4pRhc9fPLSPzYvST/s2Z5i2
ZBg+vpMBkeaTXCFiVASrwDaQogn21uycnnQBHo/JPpK4fhVeWriVBv2uvtgu+u8M
W7xy5b10YLlXfEa+cmXbxiqvEmBhCFHLkXFEAVTu2Dd3MwwXqnexUDxLj+EBzzmY
5/6VOGCBE/ISKTYrytWrenQuXKcVn2+hBy9b67stuYnjmzSJ5XKtXlCV+fyu2Aoa
k+iyGWr069osMBhgzkkMXCpvxSFvKbDwFF2GpwCzSN25X7PmNH7HtMdYZJ3xoqkG
FCrnrIkdB0FI7kgh4L05DoyCJFJSoM4mhijWvJMVeKaZGYNL84oKIy+ePqpKPXyO
03p3CABuBLMz6aq3jRKPgKhT/tFdqpSpMRH6K7HlV+lnuRAq1yALbjn7sAmTbiSQ
XrBRuTUisxBDzX+XOYrkw/XjlvVrKJFa1Pu2DHaHYgylDFc/QCVb/T1ged7Hcm8R
EtTOqy2YYcXoLIGWyQMWPpyAUCJWyD50bpoalzATSxyh2GNi7A95IPpNZbDg1s1u
LBAWSsv8nld24ny3oG9mVbzGOgUFFn4q7b+G4/f2CDrftXefcVqhZevkdXmnF2Zl
lg8xflcr1/tPEqVOQNYUUS1McC687AnOw4q09kVD5691ZW7TeMcgHsbTg5opnLgZ
O9zoWfhxSBO3S1t/JYRQnzmoDyk5g2R7cNA5Q99ayHU9DTJfygA8XHsKBQohn0qd
Dp23ZAcagRkVXzDb8LxqSw57J9Kwtc8JZPZdj94Dk2r22OBbKcv1EqsTrZp+xVqS
K38Qj/JvVttfgGWgVbwv8Z7C07AZy2YUXWoOOmwzZKKiL769Zye+DSdTVtFoTy0B
iIONLTha0a/RZ/LHHDqCEiA4vxYytY9aUBAaE0tLYnCd325DNyW2TonSd40VgQr7
e+xCktxl4oPEYTDcp6dAtzMi4/fuvds1zq4oWMlQppvSo37HMJLFrwY+E1u4nDyW
8uSAmqoeaerF02UjCugKPtr1QVTWrnAPD8qct1XyVaQiYFkBfiyI1OeLR//PPfMg
FHYcukGEeNpSMsQSuneOKsqvWHlhsg4LFGCp0iDihpq51gMH8wBcCopyO3Ukn5o2
AmdCIiLUJrlcEvziz72mLvx9hsIEO4p1CX1TCzBn4iR+CE7R21SOO0GPDkeU9oBM
md/U8+l2jVjWU2gV4P29Gs4Yx4QdcKjHyA1Unjf5UPhR0QVpmCAWfgmKivbMq1oj
p9pJ9IsNbOy/LWswVEOJCCvCGVhlaZvhoZFPcJd/dsMUNBqCg1sXOUEvVJn4/M7B
xdiVbw+kDb/H4ysT0Q3URN8pgpZRNJ6N8mROr1NIa2kYv0vRfIIhTTo4kTBsdwft
r9lJJshuwDDjnWiiNKKQFg0ytB/2VAwe3GGxz4oBU8AYACBrbVLPVCXPynfDwuEg
1DnUzLHNHZTzyj5WTuT5e+wqk6u9a/Z0INAKXhFHFnxPQsd0FJpXu2KEdHT/bLW+
LN/1wPkLt1hOPd7rs0v9USYK2Xx/oWUqkICwDAN/2DWgTEdn2+cQYZ5d21kCRWCL
9FawhQzs+284O9aOXfm3Dl2dOovdAEVy6pQlORDA2c60khIKBecwRjo+sLyrWHJ6
COSTshTFe8CKFCH8DFuL5rYZgpObEWO+K1xvf2BI9Cg+X32hZomnseBZzyMK4ydk
eBcJziFQtXPyxUytGINi5bhOoxm98kVs9Mv6P0FfojTtLiv78m+dtctgwoxEEqDX
GYB5nW6XwDmJSRdtzQUb/pZ4LodZM80SlAa+ElHvYx6CUugiWOymzfKuvpYCr7mI
RMaXPT/xKSUuPA8NkUNCeQhu6z2dfHvUBdIxePNBWLjCb/hXwFAj1EDc2KkpQ/fF
IFO2bYAacsAuQVy+VofPC4934eS5XfmCpJRSaINCui9RYb4a4AoJOZ1pOqJwu4n7
0yRdreW5DDLO4WyKTOytv4U/hCuZABfpdqsHW5G10RNDK2T2svhURsB4cX+dZsEo
P40jan4wbM72dLzEjH85THvelxWFSZRbmT03wwWxGRR4nlid5uF69CUOjc6Vb3vf
4YSsYOhjsHf337dGPACktygsAMyoSiv5tBl7At9Xh5mEICOgpyaXFIEv41605IL9
/W6ybCrYbTvNpU9fLExq2/a0pGAqEJYfHQ5I1LQ+XmRauDqy2MLXjlex6IPTnSKF
xpb3fYyrM2R4wS0SQU9HYRsFKQBuQIiius23wYVlX3gYLiyvXKCxgm830x/Iw3YC
C7QGwHuc32pueisrB7sqGs2JYNXvglj5G0HuKyWTadailw0dBuKUDkwMmFpeLLYr
PF4CMLaRRm5uvH2EeUBu0hxlvnCoS/s9dzhNjqAe+QPSE6TfreeZfgj9iFZY3P3n
7IhrEYWUbn/Nm9z/v4A8HM/7ixlHaUnx7aswrPJyX0n+q+1YjPwfOzcaT68SFrwI
I20SkeQ4bn0ufaEJmB+0YZ41s5h0+gu/gL/1CQ470Gt1MLhzP0e0Np1gjwp6P4eK
fvQ+2d6UT0OkKOEzNPVtJgytHfktj1yUlOLJ6vUM3kjSWAmV/8coW5pUn1yWxbRb
lvmSvOq7FW0IybNYGcR7sQdjxK9uSlOQqy9yhtJa2MauSw/GBCfEq3s3lN9bHhJ9
QjSGUlteZ+vlZjX8/omHg440aAC+I1dAOjvotW3aJXQidHL/JiSNENoOXNtUXhJG
xPJOEU3H5e9BJljqaKwWPr+BP9n9d1Mf/qIv45sAvI25c3ShcMXqMTXJMKL/kdDw
1dQciGv8GHDwm55NJpACpu+u2FIe1sDhfm1eCCsL3rgFJ9U9EoBLIX/PcWlBZSvP
JULfD60EEjJKpJgAx3K3VIlcwkVPFU6riVW6i6c078QcD9MF+xZVFnK820dxNGLE
bLadbdOSW/vFrhVZa+mU+INIpIRz7mIT35MLQ8Wvr9/a2iHMzupdPqlv4Q/MSH76
v4pothMYY2tC68jBVKJrTfjXMLAYtdsJF1/Hg4g3/qBEf09UR6uaKAPl5xwJukW4
81tBmb5SuWv/tjJ0pDWZoz+oFGr8NLj2Wz+b0CLFFyqlB4i3XqBLi5FI22AgWxzV
7MOJ438XL/bcD5pWxVCmDVmtcT3MofbkfZ4Jw7n7o4/ppYSEwquxDLs4OkA5xnNT
yh0NfSLu4u4zovRwd3mJRGUOx9bvKfFITZkZ/k5JnyhVqoLkXPKCE38KXeNYdJ1t
vs3+AOceAVZ4SRD+jGKMb1ImnuyiYTyvVTGjYxQEgyLfk9Kcv45VVkWdca+1i0eu
0DoBZa60jgzDia1Qikj4niiqv9ywMTXh5aqW1+pUB38onHFWnXJfdXMZCuO1WyNB
IJipMHWVnUX+XKtDr0AgTYXPHQVzJQRH/NZFkQD/bVFRukkz6ieEEKoxkY58TxK/
bLAooMdvuTvjwnAzAsKXo47+EqZEMeTLdug+W78sl2/ssPb/BcsgxMPXNxl7c9Bq
DQusLm6jpVQphTZ23Zt/S7tsqfSpqhtrGPu+f7GAy2qdq30GXXjBQ6RKyiUTUqZa
65xrCBKc/ihKzdIdRFefA3UNn+BtJgNEdPSsVompf8zrxCjbahpfx1EHB1MoeKq2
zlOzItnp4mYZbvF+vkdxwJhKBRNV8FDfZAGE6Ty7nLJWDS/md0mSRI5GblWMwMKW
DLK69g/q5478+Is4gnUP/KTdR4F0xBLJXm4XGslsu3oXYndvW1weEYCOrosWvjlz
Kc7XfBmk5Y/evsht+SGZywSDTmF/UtS9xYfeZ84F722VDzDnCPzUJJG0TbmC+YfV
kyhN85g0ZU39QtSJ6SIHpX9ptdYCFC3dHr/TrU0tAI9FvAGnAHNyvKq8xBFz4WX6
6Vcftf1HryJ3E3WuPCkpgVpe533+mGPRIKaJRRptEnuI+77AnPJCOJrw9gqFgYpZ
oydBVqBduintleIhOdaKIul0/JKcf5/JInwwtVqYx9Cs0jSSCRn+XMFVsY0uxf3+
BVictHh3iIvtCEn24xhJvI0muV/GEC8ONM3N1tDk29aYTI7J5fX+JyrNySUaLMU5
U2rJYT4PY41GwMsDBuI/L48DcLAhs55oxBb0kD1YcN2WjugwGUgq2eh6lp4A5/2L
TQeCLlcESNSCEH3LtdvJwi3yKq+3CWR7IbRBvNKCx7XK6XZk6Ll+SM3h/e5UaY5M
6UERLk8gpMi5DFrcEHGsX2mgdgEEHM27CqHHOPVpqj3RJ+XTR0qhlGs5SlaIJ+Ff
lJCns7KHjxoiZikAKKwmnnxGi2giQlo0pFMpA/+R3J1leY9JsExPWnvrToSAqW3E
T0ZDr8SdsmVApbRusm4mlTNVSTWEGBG/BvV4QOGrE67cMSCHy4nWt6V9/3ecowz1
+2fa41+/jGOVNjGCxTjexaMX9uf3q1o7z/EMHTBinKTMaYYlThqtBY+yx7CqfSt4
DJlUSBJOv3byki+KXOgs3OE6NDlthBm7f+c8uEP3P29Hs/rFdYmG2pG7aiI12Q9C
gvc96ZmCcqcoDjaaSwpljqUUtpaPfRxwg40QC1GsevjiepEMMDDJE0FuboCqeqNd
oIxsu3vJCkjKUGT3HSYjVhsvuZli9yKAbDjTor9kH5dMebtIB7cWTWjK7a38Ql7i
spkvOIEXOoVk3RF2Ya6BHuY7cvn75aKKteeDyLpTND5UTJoGnv8Neqjui5SvG62N
8ppoLVntuoArlHF5Z0PnZ2EtqNudblmx2jfKscSvLuS8Z0Pcj7q/gKDnVR61z4Y5
arv0hdPubQki6TTvG8DqeBmr2MUSydzxJYK2tEBdhnU1N/u3L5XmCqzMCPAz7mn8
02YZnnntT5uhtQFmREI+u4HOW+VirgbXysjzzzDgX7PzWCLWcUDfCFForbbip65V
rFLrLtEMyQYFZ4T1o2f0V/ZKdRiLi3+ahFUe1tB9BX0ddA1X5z0rRLVDIcLTM+Tj
d8UghJDeDAttIAfl3Kl/V3Yah0UsPLr27q5Fkei0m5VEOIRAow6GmhFW7jcQcVqq
64a6IA+oCPULl0fSxDAOVqoKzPZNAIH5nhChkAE3PWHdNwtRgwxXUtLop+ys8Lvg
QM4AQhcU9nVSY5CRXRX+/amOCffuV+hnZjV8IXBy/KkeKrRnU7ovtTo3/BZQOjoK
TrRQqL1P2aWCwIExWV8LKdCEXf/s5XjemvtJbJjLI7dlLn9XNnfsBJPuz19g8A+U
gQNuPv5hNtCXuZhM504yMYIa/MnuHJUsvu0h9XDsnT7M/k9QS9bNkrZVwKg1sBPK
lPdPEM3HIs7IhcbRcNkHg0FymYDIdvljEaveygSgSaMRB4fKIAQ3U2hgFtztgjK3
91ARS7qnxHZt/8hf7+SmG7K4QNpidJqN3hpUPr12UtX0ratqnUEAxi54j2f1TJPV
DNMuMumM/9b1UsD8vN3fT2BPjHYwfGAa75snrly0JALaiW7ku0XxdJ2ySuwk3Gyr
yzboAWQGyrdjxpUoE6A6W+GYwcwEQeKyRUgjgwgf16C55QI8wf97yJZdV1+KcPQp
HpNFfuAhGJSye/VZduJvFbbRJsHaxZO6nRMFMk3fhB7sfgGPiLHcuc/Aj+eui459
Ub4gxuSkH6odfH2qE/vnKo909Glw7avwYDXVbYZiOtb3QMOfaYS5CM3hdFR9+W13
9YRrA3UFoEmfZctyqQ7gNRhSsTAq8azBdNI6tYlnGvr7/rbgxWCQ7260jOl7QQBn
Ze3CfsVf2QylC+QTODjF9pDmr8Shkmdh0XMG7h2vHhmj2C4FsTPhXQeoe0PPtnB3
EdSyHip/7rejsYnnfc5u/EE2pdNFNG6j0AHyoJgN+9I/b6HnYy9uZEV2GAmCYWrx
OmQfpwdZ9j2JCzM92AcUf0e4oFVCoPBdZgmDzw8DjE/huPGYV5Lk13PNAarMi3og
NhqWwS+7/4KH+f+95+VYJt5kfw7JCs91sISzUDl9GdVBfN4dfRCIwtpic3MArvOo
McXjtyPApsjiVxglAytrJt/3FT+djVpgFLkr9guVKdQvqEJswQLDT3wP5e0NV5J2
flNe/08SLHMENv/7cyc7xab9t3L8nWtQjIVzM4Y2nkYtIIdl3jR/qV8TNIDmG9Ak
hq3dzY8ddFm4JqeHE1OaZMlADK6Jci/OVFPtNqlM9JaqMbCvOM33hLTF+5HhGRLS
Kxh5UXtikYa3cHH0w7RgtpPzEf0KmTlmwnwKRXGJpji4TjU8E6I4+X4vKFwbHKYR
DBt/uKtBrzTqd9wjQzN3VGHvCG7W3jgPMUYqpr7/9ExG8Y5shjHcupu/rvmoDWUK
TE1Bdla8MnOlbtvjmaA9cnDa7fIFVOeSsqIzMuWOzbk3u2O8PqRdGRadGKHfncnM
OgUq02ts68glJL0RSblsovq0KL4QqtwE25MwcTu8YuE3qR5B5SopHQ/hjqC4hnxM
17GR8VmCXzpNKwLhVlHuQN72LdBQrRAYwr8BDBj1jK0n2qjvS2aUGE6MN1wiacqq
x/y1elN0S1oWNVVgkADFqpI1zL6t7PDnlJJbxY5tXBWdhrkUyU968Jd3CkochZ7m
QquMiNUBtw87rcHOZEOuxIr6j1mkqz9BddowVD39vfUmylwjno1omrNGxU++eqXH
N8Bq1r5u/AjUd5Gg+XOkp1cgyTzXuXoXjPu5hx48kefmfXrEiW6TCwSdDF92GnGk
XhgdDyC6kJCYbv+77UBUb9qFzfcyxC7kjHv1vyVx9svGD3mwCMOed2ATwhT9SAQm
U9t8+XWmS9006gVYc2WkcrvYuZTTxSHF97+aWgUrdcr0C0R/bN5yZsqdSBVO/unW
rClTnkAEeyNpJV1eALYaJ9XWa63maZo62BEzUKVzg53fcK61w0nQgHNmX0sm664d
kXcIQohpH4DLuxY/dib1yfAL5YaSEjE/6+y06FgGkgqG2URP7mEUvk5Sjui3ZOKS
f1cUrnzS7QMd1XTxKNhShxnhdZbn47nDJBchNeZm8aTtHFMaaJnUozfDJX5+9aZa
YvpIkFICK/9R93OEmBDqRJRGvZ24XyIoX5njJeltJhFLvEN1f7zwlBvrRypd5aQ+
fNZXt83IUciTCpRNbYsP+fI0LOwW/rFCtGLlIx/rgYpjLrnf7rvNbC5V8sWEQMbE
G1uYYO+cnF/MsAs64nIgYvr500c1ah3YAbRGJMEv2Zu82N69aTeE4od+/4FhJhcS
jeyt7Kbf0L4S41tMVb3j4W6wmPizT3caNhWjA/Ro+PxOTBBZewUnqGUlLDpSrwsl
JDrc1mcf/alEsXXQ3qUyWpO+KFRds+1sTAY7j4DDSkyupnC5cI8NWStPcijT/eCB
hG8WATjnyrq87gzZHywdrkwuY1W+jisXe3g5mXMQRrnEZCc76voKMbGJBg/hcHhd
BNlo0f8e3+QtG5XC5hB9Huhv/KhgzjYx3sX/TBz3cgNAL4Rb3SAAc3S1SK8v4ZDu
FvGwxkFdg90hfINWBwkU7CdqLvaYjfOFElFkrxuosftTqO0oZJnBYK+ASOvzt/ZQ
KKtrCGOYEknNBQavE1ej4GbroBUi61e19GAEF/GG3yov0fL6148jI6tR5wddxCdE
Jz71OHbdxtq0CcU/AT7xKqNT3mlme5if7PZZiclf6tAhrYuBOwIpasq9qTKj98kY
Y4Ll66bd7K7bUQ5ytByYWNGrlfPnhDpBZMiQuLiEQXxCidEKxNeVWf7sETNEabVM
O4HGrsWrLThWsVPZN2LyHrmsGgzN1lyJ7eeI480FsvIIcJUiUhKU21rIAkyY8zE0
iV7ZrVRZlDHulyRml8JhwQiMa1jEAUXW9nyEfiGDrFSHh+MDt8XOmUQTAmDSZ9rY
vd785Syo/a8TPie+MydpHoJndARWtVovTmvgvrEZuErQILEbUe1Ytvv73SmELMw4
gUhaK7J9+UYBzwMknOCKs2sbeT4gpUI2gM5IgfvfH3FvRZ9yXHzWO/0zZtkLghwr
jCZDE6jDM/034iSrO7hAfsojQ2uVRAKg4U0a1a5Yb9rowR0YRMDBfJOOs+33TrBF
7f/FnSer/q5P5L8/5ZU1m+JT2EIOmI5A1HnzsbosD7O7ms1lkI2P2C3lUHfexTAf
VYc4Pz9575mYtxE6CxOwCVatfrYnxlFIJeW7aiv3hWlzZ8XuMWQ+X3M7sFs8vB09
XiGLKQt2o6hFQIpWxTcmgRC5xS90OgrdjNFpygx4hJBv8JFFufZ5so+WMdZjU2tW
1g2ymQLtu1etjxY0MdBcS1Me63uSDQpAjt6PmYduUBjheEBzFVC4ooUckFvNbFKU
0yxZDm3MtdV5UgLDhxL4ckkw1kTvHVF4GzZP3KOXhQtpu/P3fxoLQbRWp4pfYSek
a+mldaC0loIS76REvGUeChl3HPktt5boFvHfHy7zd0Utx6Ukap1mz4T2TV7bZsJc
4/viO1gwAF1mcF0HAfoM8ctSpVlrZwYu8Oi/4Y7E+gPKOr33d1kNW5J/J+dAQu+G
oAU4StBfNBFUCdz8Edqdluk5NwJ9Xrmvx63tI8Ail1K6O2sOaCMdRL7hqIs2eDze
b3mwov+x5A6Nh3z2QGlY6ocA4AivmnB0qykNa3JDgjmvhaKwDs6XIOekh+Y5EBVa
l1SsnJ/tyf84sIVOmVnkN/OjiSg+8eRMEIo/qbKo3VmVZkd5QfCaXjLnfrmaZLIg
IzH0aqRyjWjRWRv0H9ZKEpH5edU0qqcCzDgCe6bPXXh6lx2xJ8ZrnaHcJh9pxThR
qjJMbGx39D/NrvhDKSXgaCdeM/M1eR/nMGUUTQTe9FBpVl1iijOwrrHxUY+dMA08
utKk/buUM/EiVKKE/AOQpg/AX1mlNAlvNQDzn2CclUcL1EeGRSXXoeSdHHpXakf9
hA0Bh0cyaLnLh+p3C9PN8XxT5WAfwSgYcVgOGapQqY7Kt9bZ6wh4X1CzSPXfdf3H
Jkmy4HY7C/Z7njeH1sVpKA0psDHfCQr9ab4RTUGL1fL5VRqpWtmZ+BPnplLFD4GL
hnCh85HR+2IawbqYsvF5CgEtf9mxiU0jYXbCCRywaqML5b3pIxxPNa/e6ndEBynR
AOr9YWNwkVGpraWWZNybWpUiiZe8zJMgFQdOlB/u9hBC9bTK84rrlJOd/14mawxu
lbbx3YWmu7c0Xf2SGFWJ8TrZGUu3tte7z3+3IUnpUGUoKvemaaAE6i6FkgAF+6/h
tyAhDT9gMID0pc3e8hye/UeXHGKbAg9b30kmKR6UuZSuzrRZWwN9DiJUKvZ2fhvF
Voz+vjEakqL19OsQyKxjHEZElqIE9zMVPbs1BMRB5NgLnfvjcuuEhiKqr02tANxX
MKdlvEgRKMS8OOXUtCmsYc+PrqdWT4k1j9cCtSKoRh+t86uPB5OF87w8fbxBsW5n
crr+1cjRh44wC0iIqAdKeSRHc5b7wR/mMwLj1V6fjyDDInkhhye8jLSS3cPP8sio
zXTdjJ9umWf0nU0dIo+zQgCsVebQwbN2wmQJ55RV+yqvAd/m2c6NQc/dhRlTvi6w
1Jq0R9uUyDTb1P6dvcfcHIIntzV8/961KnbXNDkqU64KgNouWSlrMz2s2nN5Sx83
OqIfJh+rKa4hzb4ASSju14jKzMxSNBPOqIon8ItEN6WFNZrR8/PHcbhY1X/FxKov
9qzmtQBJSUe5SVdU/qPPxtiytcQ6qfZ7ttYQTSd6GR/20J/cTqZfWO2gQSWmJRvh
4Wp9JrIxR6ULG4HwJDNGibl38dponftOGKEYhmJUkuwq7vUqbHmZWM5GiBYog32x
Uwmuw4CKKCcJqnFq+fkSTvvy+lu4vxVHOiAmDrBi/ojDXw9UzjcG/LPH4JxSGx7z
VJPS3s8HLC9S0G5mS/HYy84P3P6ALaGUoGvsYUAXJMbr6B3768aOpUh8ZjW68I31
rORgszDUqotH9134Bj7LDtxgnDjoA6SMK+cOa7QncSxcMbh6wGoYKCFLHBwd0f3C
3+XMZE7Lsbum/0O0JBeYn4v1k88duknrIAeVM6+sM5UZv5I99LPC5ru9iiX5sOR9
5UirNnm6K3ZJzs9xI8YCgZpPhUemOmPFRTWUg1ke274Wz2i6JH0aewJYP5gPTuAl
kvozJCppQguNZU3s8EHgJURknA/Der9DpW/096aoxRtp5yaRzdS2FQfDbNiEScpJ
GQocfkzLO4ucL9Fwnb7UuC6UQ0+OgpNkRS732q+rE10E50F1Z7c7DW0cmoweF7dk
+bdT4X1KQqgQubKGQ2yL6wZUAfLp4M8CX9eY+D5hGRYiaiQg9CueaCxPPSbqjTEP
ZB4e0efEhpJHl5UVHS4W+zMD2jKaM1/H3qvqKMhmawC8HoWk90z/h4CMYTKlySeG
ZD3Ojd5SDw6XKWQJL/cRJ0AIrNIMPNBCNDfKPOoP7mOlSfcK9LVi9Vp6FSeQ4M0j
lunnQj71+NFp0+X2HyIH7Mfu+0sEefanxnVLzNwSncjgH2U8edDO6WdC2IoYrpWY
OER+4ud879LqInIngGsvcFZqJJW6lGEfs/pqWdXVKlr41LpMLUh9N0ATiZs10d/9
Z16HdvIQ8ylaMZ825J8VklYiMOyTqU8a5dFLNvoTEILRwRcoMLq6j2jhQd+GUfPP
euGOMhP8MafcT6jLAMsuzkgq0DjHUXY1GyELKRT5rPie5o+4HWRZT3Dox1IOCjhd
Bzw5vPvulp+XGwJk2vZjRmuf38qFFRj+uFlLe1HRwLJnFsA5nka6+OSBey4At0Nb
6/DwVtuPlaGpUp99hYqhnrYkRVdQzpji5d4vXVrBVJ8XOrcaLzLIyqetkVxKv7my
2TxwTwj50NU0uZRto/73bctBozKcp0BhTH6N9azNPgfAQbahVxkj+9l4txUnmeai
wk5RuQKvFMsYjbEe6VCyT7BpChKPeyWS2jEx5UUKXJ4e8Si/2ZB1i8hvhcB++lS2
Lms2tjy+dy0ngHnKf4JZ4EM74ZVDyUpMjc9D0lj59SpECZtnH99DN1EqvT39EvuA
QMdHUqm8bVFFTUlgEVluuFS27P82HuqMup26GyAqRytnvNF4hOR/VQodEmFhxRcB
YYW+lfY8PsEpk/PuuSVMLUwgkVQwXXDX1wG2oz1V9Ql5widwfAHTzEoUi+J9aATq
MemAAY53vqPBqH6nS00Xe3quJss/LePJDPDPPdkqXyuvmpE8eN/QICW7RipIltKf
T9iHWe4cCRsWlSiY5Wgdhcd5tV42BSBpmLCSdAZwXZXej7KHSWz+ziTOUHP39LNE
pCj1C76RgDyPhXRuctbomDWalxMVxohM/b6vVeSr6AzAsOEoCMwN/c8fPG1atuhE
1RF8U7VdT+EPSL1FuK182pbrJ5qYrN/spEstvw/Lv5TOnGfzd5iF2UG1nnX1tUV7
5/Li6NgNUh5ZHyyjwb4ovYEPwnxfgWAZEvELQhC8ssJHCHHTFHGDUN8BD7JEaIoN
ySDosiQ/gZLiIMFMUsZ/q9MQkT6f/ZhfCp2B22DK8ro/eJDSsIGcdRyPw01pSvhI
kcE2QN49hnj6HWd9G4UCSOUrLs/71D9Dozf0yc7I1shcCYjLzu39CrfD+1UzE/3R
FYAesWvg9SvzCxskUkZq190WqEZjtulhxk7lMoosFDjoVVxFblPaeY3Yv9xfX0GB
1VeK/7OSmOf9ozAbaqGpwkW2olq8PIeaeVj+frzmzn4sJ8Rn/z4OwlmB8gtliQLm
rJRKIaf1jssbUgWITfLr/yN3nSCwYCXLWrFOAcgPhFFWAX/SBk8hWj4WFRYII388
UXblrOhR8UdehWDbZJc3rFBhAyX0zbxRNq010VlIiAb3DMO0DMRRgSOfUeISeiyD
yAEhq4IvzvUqVN1qQk3t/4+MZWhehVJXwU0/pZNQXZNk/DqVFV6d6vke63cN6W7s
CIpjCQeDfXsYiDLpylUPv7j1M+aS2MpZxdpg/pKcIDV6VnEQanJ57lZrVLJCqjaw
sLructA9pPCwpZKJGJdsc2pMRMFbwXa9PiJNQLiugEhMn3Yhi5FLNDvp+WmFEFyQ
xuMoCyFN9R2LrUrjNGgw8lNKvi5K6bOZdQCOwu9PBSR+XfVXJa8UoIyhaPCrffai
X1oCkLzuonsZgI9U01PglaXQIg4XlBrrsYWZqrLPlBsFdF0FgxdF6kEFIv47N3+B
hLYgJzRaw4ulAl/euzTkrrB3KIUxx31nsFgCZ4naJ2v7jSRzk/C7rZ58wUVc2bbS
JqL4chF0gu63Ma59FvAjndaxmFvy4jYzN/ZenOFHAXw1eUtjvy4tMwuv/XDWb+sA
IKrsKIF7v1on0RGN7G9RctmWLBtZFrEitT1dXKvFyUOF/bYEAVrT89X+ErV2GA8o
J/Grl/5Xj14ZLuLDyY6nZmkCpDGhhM1L7kp7/XGBSggSP7CLud3QYUnv2b2j2acY
X1Cc4lWMTC0R/9h1zjBKiki4a72lZHrCYNyEfZUm64YoIILJhFEpLG1c3wIaLfI4
uC5TMBszpfq7SCU+n08Ss0bXrIQhhR8g0lWgl3RRlzLVbn1lsMhxSnCon5JmyuZa
LLCANajKVWOOs6QTZJ2DjDGIUX4XxhS5KhgXEoei+l4ZkDVf1CrGQGCZcV4y0gL2
mcmViaUg1wJFrt8toBop267kG0JzJxiHBlPN+47UhIIrMlAboCcP8xCne+ATMJ0J
9KVvjPSA1X75WBFnIiKC4Ta0mPDJf0UVBH2e6g7k+5K+MLd8PpjP28A1LkLvEJ4v
9DiIC82KJjVtdgdxCaRKnASeyFqayPQ3AC2Rt1b074cvuJVz7kmpC5+GvEqYTHvu
p169NMVIyYnuuOTNBbcEUG694ObQensR+DNjshVKn7wZ9MUf3RkvCsI/1ZDUBL3F
amgoenmw52gykvYxvO4GXezaNHgVTgt3xp1unw+BwJGJOdTkygf9ykJly2Iy4ua5
e0m1hK7pwkxEzM7tLBBZ8kPqmgvdOwsj/hzUD41evoT7DyUWiAdnLkQz7GhVx10j
VG7PBjhnicxgHZiSrP4gUQqdCRU2zo9FO2bpWiAiie0D6arNmuLD+/rEGseo2yuh
Y1BNrjFuz+ZTccSONDtk5WFpLFdcSjPiG2UHvOxskR+n6xRscRYEyDRYvxMDr6qU
pVtCJF210hCd4xqoNG4inSAaNM4iJPJNOyQp9gr2eSZUOtmdydim09shRB2Lt3AL
t52fiBAUcrVcLES+wd7kNtSdQUFFFO7qV1YsXA2UH6Kl3noVR3r7BZ23rN9fiVkd
TsgzvrZtCwy2WWw6XnzBkfLMt7GUDBulnCOrGLdoyEkVSwXEAHOxDQV8LIf9jAaE
0QY2viAIRjXcnicR7LNhtnY5/6bQUFMQZp9hfrsaTcXIDzBcjO9rACSzG2KwN2MZ
B8G9haNRgFhtcAVny3T8HUc8e+IW9xed+/cH5CwUfZvczGDhD+WRgMjw7PmrxQuj
GwJUDg1WFGvjBlCrUsGvIcENtlrwWC888gSG6tsou4PiT11LwXQQdymKDYEAvspw
whE7uVUNw8uyOYos1+AtYK677yG5VnfxPkCC5pADdFqDFi4w4DSOJacjyPgTD+Vr
8QAmVRTWGsvjOgpllFOPaCfgXTdB2gWQTIeTQzjVq/aDWA0zoYthwKiG2+75F2I6
lq9Ofeafk9Az/VP5XN1EhSH6aF946TktlTSTAh2wuVCvzKi1R7K/ha4kbjAQYsDx
uiHkbJMf7FbATk0tsQ3ZyB5w9jTT5qFwHslVuAJOjd+1/O1qzUx6g0MuPGvFZxmh
psillcHqFv9hfJVNq4ASZZRAjFjuCVXvU7Yoqs5MpFGZJgiCq8ok5HkWqgdn1jan
ldUAULl3sCGALXHFadxQotteWIyLovUbTLRJ30f+HHuZXNWFyUo5tXAAtM4J1bwN
nWa4ZFE24BiKj67I4vCLPbP6HpBdTQDHfMNgIo2nS3eHwaeEcYV5UbJv1KQMEmqU
xHIC2NE6R5jKwG+tNjJ4/2a8D4OUFWyUlcY7+R+f50ca2xNSl9Dd9UZHTd6oMbPQ
xoAbEOXwughZyU0TS5ZEi1ONEc7SHEydqhL7d3Oh5jfzTpb9LECkxlOH+mxQ00Vw
aFOGDrgq5nkOgXfsQc7f8DyF8Mitl+xXax3aa05hs4dd2zrsAUymqNOQou5eQALf
bo49pqcpgDxWFZh7Z1ek3KdXK3aepgidSIBHZpyEFnOPPnQMFciMEAg1hLge6FMd
YlhUcc4tb5tizbkbVQOZ55bIQu11O1Pq3d7Dz0JGp/dFaZ/uWSLJgcHlIWIHlXyX
WMfz6pRi0LuCg9RV01wSIcaQyEsWBKaq87xgAv48oTQKgVIi88m0yAXasXP1wTIa
cTQ4ca4fEoiFP9USWrSiE9aV4dsCHl82KQmTOA9f9127CPU2ljANCEHAWlzCRGU4
DNhxWOlvJYjTkRhp14Uc47ey7hMB4KXTCBe++dr8ZDV34jjZ0iVSKjBYBkAWZz6Q
GMkhz/c4cyWm8PZXPBAbaFHXL2brfTZnw2exT9wAlcYRcktTAid7a3y3BswXerg8
i73K5Tx2WppfvObsImDA+S2k6wDlSENnbao43a3yvdWcqRYS/ylrcIYD15LXkazx
eWMiCMDn8T1DP7veAB6iTkYxpM0HmZfPJgAA2VdWgQiv5uEPl7+R75LLWTbtdMsF
WPsghRvB2taDcwHUhjftlLj4OEn6pYNsG66j0JGSkqEOn8UyHVRnREal+Fw+6OIr
3amSipbvqYCfXY3aJGWvMQCD51i2KzEuoTLZbmtEZVKbAVSbPlbIqKzHgZjkZ/4r
XwlRzOpDOo59LnJ5JlPfgbGsb8r/dNjjwvwUTq0hmxpqPbhAHEDxGMSnBTNxX+Zg
DOeVjRHUK66cHvL3xmFjIfI8FYnvmQhVAzS13PLRnE1GKw4L1/xnvZwH9KrVat6e
jhnGHsdtM7K9Wwo210U3Sl+GukQ8rm8CeYBBYI4u6zYJVH+QGx1r4sagPjkinBlL
9BhptlFoSwmd5UZGAR9VUwfvaMQADUAs1J2ubsLYgUB7Up0iDY88fQDWOfEamvkz
M5Q2SHWa3Si4OT25CgP3ElRWU1JtwzUwsJGyca6qLek42iUhWRKFpY2TK8cRkGur
Kk8hwlOelwCA/Fl0B2T1ZnTLRVy+oSTlwrU5uaX3DLTVUpaVoUejYlgUsroaO25j
lgpS6+JuanAblWYgMeONmxkgNaLE2HF2/YP5+8RRimYIGz2P7pn3lpWQA7i/JQFP
lT6gQnQMUzNKf5wUL2MAsvR8iXBkrTDzIEUgVtWucTkBGK0/BwDo2MucKim2uINu
CM/Ng2bedTQT0Y7UntrVumB8gffABWBDc0RwsPqNBHX/3wLlOsftR6jYgTa72JRI
Czid13L7KaPCxDWAF3+HZCsgi9aXjWAMQ4J0mlObV0RYaPpqpeS+qnQLdQrgHlhe
4+eShmIw2LXWhENky4BWAqHTN1qy2q6iDSlKIlLVVrcjkVlIocZSLebfZoUWnopW
amMbFNWRT98LukTuXpxxS0xOxmCmMki1x0Rwxxp4/p6hYfP4WqVHnBjO3ebomGUU
sPqVgaDO+0OI028HsswH+3uSftQMC+wF4cYxY3OEUYVDCyAvH4xS7ejBp4DSikuX
PvoOLAa2LzV3L/XpaZ82j1IcZPFSwVBWNqU+OxWWFR2hHW1+npdI0cVd7TU5IuMw
HwU6Df0W4yA7w+pWsrbBG9Do/mkOU5j3Q4FKQeJXbN0eA9EbMnoMDL/1qPA0NIJ8
rMuALQOEfjevS4nmRZdaDjaYOYpg4z2hlGGhRS/3OmKXgd9++eryHASpmd1G6wnh
vFFklOtB2L3gD+N6S7vPCrCfwoMA4CEHXAk5j9cV66yjS/+GePNfSVQhTCULP1si
3Noe3/XU+5NxQOA06HkM7JXXzZr4+RmAXwa3DuGSLtIoogtHEnEm3A+wZW8xRSUZ
a0Hfa2V2zaiNpwdJjjaucU+eOHj/qbaPRrOoH+xIcndCz7t709wieHcchUPGLjmh
AM1WKC87U6FgppIIYVZ4oGW7Psmppkry+ExGfbQvWKIL8YLO6na1hpQH2Ip2VLzo
ag6LeutIuwPkFlVMbGB10QRJfSI0zxHXlmBmrJqFMIhbv8hoVZCVdJVGMK0RpjUm
fZ4GFzNSzqlcNr4Xc73xFHIDFzuaZDtW6UP0WjBVFl+YSJiBartoGIYWWvxVo6Sh
hzsGq6zEhF4zD6/EcjTVAB8Dknr91ZFv9TI4GRDvG2jh/GYzvV8Hmlf9Y//TKjkl
42Npr7tB3WET5Q+zka9QWlY2sbePvguGYWnbrpn5Bvkwsfje1j+bwirJpJOUfLzp
aN90k2ahAeN7CECgy8CAMNlBqsMcvUa7pDveQCTBt8lfvlQDQHotz9SbDgd87jbV
SC/gH9Yt0xGUMdnZRYcbLocRDNQ8PQIM+vJkf8NPL04KGbqj7rY0arqh0vONl0Xp
n/i2veFwmyqyuUxNujhChwhzYRIRaaEZ2VXzQlI3tHFmk73NfIjkS7JB1GdcyFt6
9kWn2LK3ttIi0HhZdd3NwyXoU3Lrdh4aCZQaAcYrreNE0Q3joHEit2o+EPcexecF
DIaamGaKXaADm4ZcLy2cdwV8gQq2zwYhMFbpmCykwLKqjdxWi4kmioZOWBmx1380
RoIFtNbZYuJDBPz//PVv9JMyoq7KNZZAz+c0fYMITM3WIHowqUPxslbpVYYSl0o8
CDq6uAb0w57I5mMYmyZJZqVG/5iN753G2x+zF39SzK/6Po88tccy4Zci5/4ALFlC
xtBSvcDU39tyM8bNehB4EqB8QNjKgrgSi1MaOFbpupdEfdBx3nZZPSJwPCyttXwD
3cdD06xDOr4nIwWXPbZ9tl2COgyWfZRraZkX3sRNSbWvuI2azSMBEfFXV9Zfak34
56FEJVs+x4zh//yfFLd3J3JXGPE3uqiG+KPqqPyoPfYbAfsxhEN5By0IIGgjryjs
ELYHYMzQgabxQKLhBG8vs43UYWHfDMzJ8FrLtiEsKGIL+29CdhS0mlWOfCsXUaJA
DuLVJlNCj/zNj6CnfOw5y6gHlJPbLgUtG2PAurBF6/EGMl11HQLXxo6ZDqETcyQD
86sczGua+UzRENqO3EABGdMg+wUE9DSvKhJLC/ee+LY+tIa6miY3EvbqsIXlRDc5
7/aS4eJ3kWnfMHkxgEixWBx+S4v7xypEcjA9CozJs6JrPY7ZJZuPNRIzlBLld6Ng
dnKxV2/CkDcZ/9c7RxGBvi4gqddj+PLHIWlAPv/etGvzRglNEftRw2CeV21amgol
bm9iczqr3KkJBLpzqFfAhdHSJhxJE4Rh7rBFzHUUiM9YrFTrGZ2tx2AB92BunA/I
q1RNIn8ZH/o1k27fKMrrRm8/JAlmMZQdGTZR3sysMV6Ppoxrfucl1MGqRTw/Fna3
kUTrzZESygLxSOC/7SqxaapJeTqxaCcnkxrhKqArTx15xyi3uvRXeAycu1MC+oLM
AczocCkc0lT+k0e/qtzt748UOVJOt00ZupTYmyBh1I1Bdl5JC19TxV/Rxz5nrmIE
7wLntn9dU+XIHByhFhkuioKKVEf71YghKMDWl6KwVRmioL3qqrSuMix8rh7ytHZX
y2c/tB1JqqAEyGfyymy/TLt8g3eGPOZgoWsVbE/YOBh05h1IhooFHMsEz1Sn3u4k
1b6tkIcXLQTtRhBG6K6+Ftz3+Wv/3f0TmA1MUgX3C8Yf60RUqh6Zzuaq+E4eUzOe
5ramL9o+TI5+Kud5lUyiIQVOYeGrpaWTa8gSzhjSsuutQ16kHkWXEsiLgUymXV0Z
a4WLGruRHxkvhmCt+4wTL66N5kB0/tynheqXyBO3jkzWOpmoD14bK7cou+l1gpMn
DWqPtXHVX8W31husOBi8V8DSPcw4Zn9LyY9vI+XIS7OVFUMd/t7UZxrWmv67E1SS
ILw4j8PjGKCYXj3dzF1UeY8F9nUnwnB+G8w8E4+2Tgkgf1hxGZiDDkF3MUFleQW8
RNZx2wqBayha2ZEzD1ifgIFzRsrn8TMHBrspuFlg1tBsxHzFusA9sBnOSaC6HE2I
ZhZr/ijW04270M0+MvbiAJMEPDjhzg+1BaPr1mXzrBuku+Ay39RY3ejSU4OekPcR
Ssf83JXKca7oDLTdhc9hSdlGymxY+/kwCgJN85wZW/cmQfPuyDMUkUxZpk7Fn7Nv
d/tdJ6Jatuj5GeDDpnEiIrJCVzCtpfDLYK44OrJacaZLcK9cQtD7L2izGf58SZ97
r+8FVKIx1KbDi1Ejb6KSlua3Mofy1UnvsDwWRaoKl5bLgN2Uw6LBAoIqBzMK2YSG
DTzy5dYFITbEbaJRE5F4gTYaeeyn1B13n+qlYFUrt5kQT3n1ZyBztJCz+ebkpvuR
p2mprgBw74uxJhx1dZSkFm9ICWLIfR5r4IPTkgYXQHLqtVtIZEoX5d3tc+8yr/8t
HBZnfdHhfRO9yvDkkNKBVD/iVyRrTItqNRw5ie2ragDhAqV9sOvCVlrLAq5br3NG
l3vEqRruTXR/ks1Ile5LJkqrXyzaE/GS7XDxsC1gFWQF8rYvW16Y6TYipCl0I0CR
QVkQADf4hGxF/LVhmcJEp7U04ErtXUKj8YZNiyxWhadSAHkiOBtPu5kl5VeQyyKp
kXubcgG7V7X+a3T1wsx32z6DzK3irxnMZ+w/ACUgZvdDAezEXZjqwhWwtynE9ail
XhuqvV90r7Xb7AnT6/ChvT89S63vVQkgai3XvzVNF5tOeyTlJcE2BQJaERU7PysL
Mh4TRZDZQMKSPpjo6FUtLm1bPSUD9tyUTFUH/tRxE6Pns1Nu8+RSjYU231Z9yLae
1mWNxIFB1x/63sjxumMTBA0pYFEjBNNEd0mPjNWps6kZ7bwAEF1Tc8i60NW+FSUj
4aSsUhWJbliT1Zxd3tMXSU7JSe5mpsYbVkBMT/oNW/glQYslq91hM3XGZMbywNv1
4rTlTb665yNlDF87cj1TqGucPZwbCs1Gu/azqQnd2d46i0NKHIhBzOQOGt/goe98
MSYLjZCrXmy+W6FxBz5mMjD2+4K+ZzHuTGwwtKw5lAN33S6xcl6ZagAeGWjZbAw6
HK6jS+XSuckw7WD7rtcv4YD8D8J0wWuo+/Ppesle/jYFH7gtQctQDGu2xzIveM+z
+Od6Betg+HqRr86I5SJX05RftCGfVYqg4h85N17pWrx6NBzPg7w8SYYibgxkwMR+
NJDKKQW0vWcAmswya58q948GJddjhbWMmVwyT7C1lM31lWE/Mygo1s80HhQCP+dR
w+7JL4kiUyHHHeVxiutRHhfiJoatlAk/Ao1vvqScvTjTWFLInXIE1seph1k0aC60
+5Dgz0n+xexZtALLTamnUVTreVDeQv213ZG9f+J2uBQPQE6xBIgrBCaw7o04zXkF
JIpd9Njw65vJ7UwceN8uopFYAIGjNZS+CazqmrXjEc23JYDjjYx95fA3nrQqZgGd
itAptvfVVECU/kwez5UBjFnCImuMCgCiShaRW17jGvkBmsvRvuQbqACU/iFqWZbk
YRpLiQpdUFq423yK6DlYYQyszFvAFW6yC2dMSkNoG2JrlQPIxm5g/p71s74GaS8H
oNQLv+DzYdrdE+1iEmDb1cNzxicDOA8lWXPPsmEkAME2kSCd/mfPPmQQ0b+hQ4Nw
M3CAp0t+SKw/eNMCF+xzQ0moUaGeb3yQOrPF00daceEB+8wHU9ejp1bpgQ7Sgiec
RoscYaoc2AOSwT5SIfJ57GinBwvmQ9GjgwlTcd5L8ZV+Su6PCQQp1Ppc/l3FWTO4
fYkcO9KI50zHGcN+/JlVkojyWg0Plhx2i/PxPY2R7kJRgAcBIVsBbm+rHcSO14lW
a8g2kPpVn9oNq4dxK6Iv14VPN+Xw1XWq5mZwx7WfeDyuIAoHqcXVvyMqmPuIlRZ8
UWvRNObl2B3gSxZIQ7MW2pvR3BhGG3n8gHfSKqe8y5zU56HYS8lIf8SekXSeAt5W
9LFKRqhikRmf6JFH7ebq3Mwz3JZlw69xAmEOGT2gklHz2VIEKmGvqsCCt0e6n00a
LeFg65OL/xTwgd6sctbsW060nJFSNc7ejAqupEmdRBqaU51WnUt5EcL7LBYxxmf4
73W38oi8m8d6B8BudABBq1V43udysqkZQw/PDGP+Q7PpUDveGlppsp8LhycXsDXL
DOHkbjNGmoKqmcfXxYrdeCyO0BPJZ4hBdgzeMdS2cfy3VNMX6tlhNd83qUZgdX+8
FHU9noXVdIZiCki7fF4RLngEbZGlzxbIER6TjQNdDIYQEBCFYnU6+XnyFk+QrXeC
FNJzXBlYOcpTOyeMhlAIgT1VHE4nWIn6Xy3LNRhk6UuUMF65XAnpXO9liQr/NFrj
tGzXyEakhk8EAX18h5hX0yplHS2ILc/HsR6CC6CY66FHavq/VUbdFeX7QgwXzlnN
SE1PYtmAgMtQwLOSK8A6z1kxHFh4mqsCyYYw+0HFPfzGrEe2euzTB9iu8easgvkv
fQ68F+ZJFv7IoG2nFecxE7jJmKeE6Pxnqorb3mXrqaAGhhWE9KR/YlNN2DZXupX2
j1sHka83io2QVj1q61k3/Ys4PRmszbNqEQtpoVyMq92zMM+x/dxrGYlxXrUzd6h0
E3HAshOeOE0nAcVluD7YAGehyqnyeJXSxVpNYQz5mTN/w6lTAfVwMedfkFuF9Cky
a2kEYhKEN6ObrUsO2PVetRH+46heAu7kjnU3I3u00wvuwF7FNEqwURmVhqP3/YND
nBJFcdyWbpVaHgE85UWCiJbjA5mA4B8RD1TFTgc3OCPzcSiZxqcl9ieN8guzS/ZE
FZbnpgqKWH9yf8guUTWKrXX/TCYUYyxRvEkq/q6tgRA00MmSc/2btdO4474/2ar2
UE3hXXkGvC+vHWK/6GkLvk5JghWDiHZCd7NrFNQ1NN1KDJ7nLHZPjEMIvO/6MP8v
6+AKHeRmzpH7e2E3Th0boeJfpwLxOTB2EhtBfnT3UktdcthdefbuzeENRlqVg2TO
1CQHUtywXLtE4I8/LjwTsVcmATUGCY3hEhvOjSlgNEWxQoqVWFDw502D9VTp/8FH
uOEdRcYFGs91ZXK03Xj6mNvlnCzKBNBdkXzJALp7xZu6lXC7jbTvij0aDxHlMSX7
tKnFoNkV3HH/zM9NC3n2napCek9/r0d1m9UNw9GZlS5y5BHu2hiRtzzM+h2sL4Oz
7NiK9Hj8S0ynkR8erM6g0RaRZiIHEPZWAHEKa0tHiiFCACcsEqnoiIBsV6o4Usdq
6OaNQEDe6uqRT+Pz6evJd8Y0HKo2om95ej3rskI3cWAFs1ra0vTFDSC78wvto+Ih
OCF7Oe1gWNA2Hg0RWRwtYmVzXgCmOruAx31/SC3pRMxPUe7sd1B2mkC08dhv7nAS
QNaqaOiuYBZecK/EVdd+6quostAqoHNf2NiAb1gcQAo3aH50mKu+VKbCw3ooro0b
lyBCf+Mdicm7yoNxpIrH5OfrGo2blslsJWrH5xGOgwNkZa/ewQWL15ExDs0/lQVe
OhFmHfDT6P1EziAst5tf8XbmUfTnITrJPBUXdQkot0erI3LK5QtqJUQ3OeSUwyqo
k/Dckh8fwWui0kxw66AH6OZRSl++Akbj/Op201/5Lj0BI9sjuDkYMRvcMC2/7op0
HURDE1svCaCfzl2NUMBMbdmjkOKMRmeYU9aUiIxj5ewz4pMJMqIUfSKEK/oSkAIC
LJ5ccMygd4LPoxwkVjPUWa7GVwqaOFT5R/bcLycpNNSa9lnvL/R4SBrJiHeviceY
9vpsLNu6ZBzH+O4yhb2q3D3IbkR4G/oeuRn/THw1BsjJ7pAGxWS5syu1vkbTg5Ro
OMxNLQYbZGsLLcohYESU3E/zJutgvnN0UDidgToZvixPv+NYkXGlzMy6cxQq8Zbn
+KbHzd/TjfX/esKqRLoBPiMHeLF2ps3Ta9Osj0uS1aG2W8xni0/lEC67XS5bBK2R
LOwAd2v/dragA4O2ulwP7TfG3ecybfFlXi7ZNeLR63aDlUH0+oXGQOYH73jdEeb/
8bJssbU2wQyvFFZsY7Xnqr7h4qnemL4xV/uOWLc+GUbrCI6z271RghTibPMmUl+r
ijK5lfnwHIgPJnTAxAA/OmMvJNQaOX18fPq0ehCqxc18FCIDXdDLT4BZs8RrfK9a
s0HewXUkYkzoYwLpG74d8OxW0rbIpf+Ej7LuUfOPSBeohQDekRgzBB4MWUMPD9mX
+lANHXMMiaO/PZ4xS2hVnNLmi1lQpIDyl/GpRYy5OqL3Ld6gAKwcOghTfgQsauHr
AkJxg69NxgVEbsYDyhTjWH1RshdDKcLlMu3k/G9ECVTvElm9n07SNf5eyQkYhNLZ
HKho5J0fFCwZw7ZQdNuknIiw0/62ojFhqtbu6MA4wourx8b/P3ZO+cZ9msod9tf8
2Uqb4ruf97sGfLMf0eQoGj/szsfEo+StRVFl4vi6q07PlzwNzrXf45n5YE3N9BEp
td2B17I6dIhGYQvoxhQtWdq5adAztSi3uxCjicJbmi6BhDlculE6fE+86/pGNs7w
P4VIsEK3iOnmyd5ot5aTznSoTXp8eT9nO6gvkcHG4FiMnRW+ysNvVdRLAyMtZGAr
AkJhfLs/z2kw6uURg0KGAjFZwCiGNBbS14mk2VDR37Sl7TcIy9H4wZ2FEamh0IXy
Z/vmLzI49nVIYCU+rsHY4JWxCVZPdvlGKE9VbFAWgP0AywiaRE0LUHxJ3SFtjlPB
wD9ZCZ2MUmHS3RXI8Xdg4vgcmw1wyRIvP3ql1kg/sYhJSKnzN577UIHw1sOf+GQY
0ZeoUN/jAGCfOzZUThcWtbwIuksUW0StcJ9dq5e7R2UpB4yksDBvcKfkAJsMLLc2
/i5treJ07pG/PwubR750cbmkM1BC/XZYNZCQ1X0NW33+bJv8EhVToYoqPMHLbvza
4w5g3R23gkzf+aEVv3BQYUmJAEVe89y9+T8qqjk0XslGsPqh7DD/b9PE9Fgl9ToC
CixDnZWgFbr5xsxyhVGaSNyAlPi+Tymc+R4HRqgbWvbwXgA4peXuXU57n4u3j208
Hi8Ytt/QZa4sYUbwDJRYt1+GaEQ+P7PyBB8/sfX3VntbMRxZTi2kEKTL2GDNXoBe
YyprfrGECQcSgl8vWLbqO110prs78eA9bbueeE2+YbcC3o9kO9k4qvQKC3Qucdeo
IVDkXCXc7QAjNMf72iAifrcv9+2uDCeEq2te7P1JWDHJiZs5Jb2BpnSz1D9mF71y
+MhQaH8kCDGURvkWW+NVw8gOKGuzNdJsugbt6lmNoBNnmnbi1W4mx3XITEuIn/HO
kXGWoh18mKUrU39L/zIWhR8em5c8qvtMxa1zlv5qToeS0rC6ueKdipeV6jUvc2W2
vAiJlGn3axOfL6H4ZcEzGTCtUIM+/HxSdi7uo1c0qALn1haD6h5RQevMZaxmW49U
99UpXWOaHa7JtteCRu4PdjuZFqs8Un8uzTtbkWfD8utTM8eSyaNE06pKT53S9KhN
l77/v+R+nq/vZs3xX0xmV/F7oBKI/aWaTI9pF8/XJfm8OG/Zv2iy8gWogHSgCoeS
7NUsQYVQHvv9cGBYpCkhySpiuYRDB8nBc2cFYpBF4wPV6v0NNcTLoUuXaeHnQG2x
mVmZdFRYkUh/xkTrFuU7mRTrPzCuhKdpCdEtIuIpEoSGmIT+AijoJZE6Jl7t/7uS
MUrTvdYIVSjAL100l87Gb42FvX14XlmZI/SvvJI81iaR0ffdOqHlaziysYF2ai1Z
Eczh6gfIrCPfBUJgCXgKtlmK4JcnR0SioDtjKui63vCkB1mo0hDa5Q0WWrWGaGql
GZDn54MFIQ6bn64i23nX/A5Mn8gNMjc3x3rTjTHi7nduGDKNStb4zvFRDmmSA/F5
W8tkzdvoeelqgVYAohW1fL/iiPOMWt0x6e6SgKd5yIRXD/12E26iqTk6bkhR7lJp
BklEe22nbkHeHrqsaMqW1+6VtyKAKL7/vctCO4YuSfb76iCvVY98sIFTSp6lAtcx
M0EAuEWq6uXfw9kgC4/Hkh3ilWQ2dPdm+NgJ/hlsuzdgP7awLcZpm32bdHNJDmsk
QPiDZ1wSA1564VN1Ilh09t4FevNPbIXaDOJ4O0It3erwcIoECLRnF06S60YXMQ5B
ttnPwDSmMievXoOJ2yx+OgnFWmOpixsQh9LhEWKX1HyjMbfMe6uaMhvd5P9U9oRA
Ejsuy0HxchNw1yorYTVGbfEoVS4JbjjMwWh7XE+2CeCIU+LICbdNLVXZDZ25elka
ziE0mI2xgwphH6/74oFdV77kYQbktlMTC2XgarU7HGkQ7cRwnNqRVsy7+E+6Hq8L
h7oYEk5zhzWd/LKCZEbHGWSH6EiPvpe3NR80cCZxF/umhndCVoAehxbBs4WJ8LZ6
DJu4F6ceJqNTuH2+cdRpfAahxPfkwcXoC6WSCN3hYps+EKqFWwrqEfnw8qgE93SO
r4cfIIlX/4R2+6ZMG5iOPNQj/v4q8ppVY3t0EqJ/lVEt9iBphejfl2m2aJi8BYW7
igTKO8winVcI/l+GsNs/Wxtwr8R/FjQUR5fC6VO5G9saUBakVPSaroV7gRAjk3GR
OFajPxMRBhyyUgnI+zubKLKS0Yjto7JYme+f+GrWOpiYySPcuumv2VpVsfgIe+tz
2s219ONVSdOCfehZBxvSt70+u8FrhZSgUtiCfy3VFa+rLu3/YG0gsgIpevxPYcPS
hH+rX2CfQJceYdT/uFEUu5sKdMJQS2qAseOCShc2NyIAVQy/fekqDqo0LdD8JpM4
tJZrvDSdIid7pWdyWb8EnYqiGiOQHpiVWYxR8zbgpTgZof5+wNL96imbfTA3qDtt
tqP8M1JCCEbWLj35po6LAofAZR21EXWzh6QowE3184wOU9ZV3Mnm7rdsw69iyxIF
vLiD7DgEIWhpcPn/urey0lOHosIBMgZuBTBAntkJaRbPV367IL67buPOz5u8eJqj
hytrr1WSGKpqblO45OTKjo7uw2A8dmLjMb9xX+/M/GHPgX6ZwqjybGJJu6ULF5fz
fdNL4CoPGqruXBmLDdpWDuaICO11/mMlWGU94PqH1VHsMnoUXhuHmmJ1ESj93X0V
A0231ywDMo1OBc/sJV8kOMbL4vjeY7TXXzkWCN634LXX+76R4pkVKT11m8cVo+is
UiDS4xesYs0u8dJB+LmYCD80Guyl3Gs+Mg9k+KLMwUNlv+NTlhlefgXgZWSG5mP8
iwiEg0KLTALhlFArtYVOCyTtb51NeeeSnZ4F4Af61TerOH3ENex2VLgcf88Z1b4a
xFOYpvKOzX7YttUOFN8cVOwrIdAbHyQeJFaMc5peZmRKujWKJU6Wz/yB4f8F5x3U
L4EF4rXrvuR2QDJbUnQ1ZPFX7vtue4cu3UkicEq7BFgoxtDzKSSGLGFtJxMkISiu
hfCPVedmhbAuJTdiTUS5esgq/ieY259RgRqfs5mOpUriRkNCVYaoyIlDcyDB9IgZ
3ymA0vn/7GQZ7tM3gf5pZMGraVBOd/ymLi/iMsfJeQ5vlgdnZo6OdMkWw4ZTshx7
AH7Wup1kjhS/9FFNghylt0vh4ANbugyuMp979j91Iy+NemjvbTG8tuFIpzpNnQVV
qOcmioQO/NF2IiqU2uIXm7aEJJoCzHMKJbIeh/4dhKHnfh/Ubi4g0N8dsAzAvY+p
KxzScs4LxTVhdPExZG1Ox9EBIAgH70/XIJzUGgi63xAZSdlBWE6G3FxhjphG/6M6
ib8Oy773LFoxoJTrQsi4UM6oWatiFcsRu6gM7QSlcfYSHP9ZU0PvwAEcLmTA3WsR
JIIXlm9wUVkIl4Pjl2zFJ//r84lUACosUdkRniJ9OwVyXKUNhMeXn9kiNqSMRhOh
cKByii1jKP8QKqz8PVvnhU3xOuil1331LU9m3QgRdP2XTaBYKHy+8pjVGEHoqobM
XKuzBACfEBObwAgBwdZqzDkbmlh4eBTjsPKP2pDPOTQKC5iQn8UYQHqqzri+uDaL
BUt4cIn6eTT+DH6l5K1gjmJWAkKLu2AwTkS7J8GtvXUlbCK+mulVHcernxx3BvGE
8MMsZeHglVaofNUKo7bEbxFcRXdc6xInJia2oHsjyVydJLRVh7qfj8NFG65pjm7m
mvnNR57/hJVJ21kTd3Tudg+J/jcUIepnq7moDNkqMKmMIzqWjWxJleuPXMSvAvQz
/AwcsXr+as497in/+83wKy2otyp4/Tj+1GdRA5m1AImgSdKR8ZGE7hvWZb5gczYE
1SV+ymFsTc1s+XRTTUW3W9SoZmNig7LypHQgzfv+Z9F/kFmplN7bYfgjS9fTuF55
kye3F8/nSNW9ODyw/KO48/JEFzt3d5BFgo0luQesLNHbyQ/6RmHHGtgDQZCb9jvD
6uSJd6P7pbfXKekZaQOkV10sRdy82GV44cY/IiD285kI/myE4V7kXPXEGb/f0zmj
H/B1/O1lW66UgiXpBhCOvOKyfmbrj3G/DYKIzXZk63YN4i2xb6Ar5DwZjgwf9fee
3humC1Jixci8XyvLgyfY6hzRNVGzZMjxvqsRquV61bsn27RPIbTzyn2BLtnNAYxA
SdE1wc4fjrxQFfiKzhD+nqve6DlhnJ4iEtSymAsZnkgbK/R5IM70ukjbB2wD9Rvq
i0MzL8XefKfTmNV2yEwI5pK9GzwrmSKJC2H8J50/PIP9GmK+O3rQhdSX28k67Q9j
Fa4mj6OVScA4RUS38wiButgtRL4O/zrNVgmOzvEphvhnQ0XwWyQaxTtKwXDxReMT
met2TTQdMkDgLwLMr67fuqbI2ugLhzfe0nLJs35TCv4kUl0QCSJb9DbJxNv5z1qm
IWG7ObRExngabLih7IhAfQL3FaqcEMP2yqP8Q5+Ii2VEQKcwDDu0fC/y5N84krZ9
PUk9c6cVTKAZrbR9TJzI1JiVyLtXK0P7x18cQBUuQqoi3LHFyKH01MJdcJil5F2m
wJRSBGSi9GUsQNAwjRvAz/DxpqMaSyPlgGYD8Nt8kx5kz9gNWK9tIkkrB9QPlnp+
Fy2H1idGL1htgctBnI+guqdJJAC9EiZ3wzhPRUzkTsfGM9G1Cjs2oKC5zTf5vlUQ
hyNKLcL/gaxhYlSiPqziKvoOZ9hVUIy4Nn660d9oKqVpWOi71Ma79xn3CJWS09Dd
z+AZeQ0IPAWLxHeafbuRoketBRzepdJtGTANJG0lSfiLiVtMMdFbOwhp2NhJr5Gz
VxHwz8oUM+nJvwgscFDB/aKRVm5KnOsStmBJVR0eMIye5KPT5Ml0NVoYUYuHRWYt
33OpNW26uYraYNM8CFpswrMMu5lt1xtw8RK7zWk3r1K8pPB6ZpQnsEtP8l7gDArr
2gHlV3bO5gRbseJdCN6buAv2ISbep/hWS1kpSI6hkm1ivzqy349c+TZuFX1WynK8
iYmbwn/cQHOtMvxopPNXqwj+GTkNNJTvr4qvNBGfztmxx7iUYCEO8Ghs9CVfMPOs
0J64MliUmrqSE2fqv2kzJmMbhUTBAJJM3AMGUcp2wQMlqIwXrxu+aZkLtv20Jisn
kcHhgdePggDMJz+pZaFjldB0xUySqOVYdYxQjXBcXbhZnALrfzykzJRmuc5TCevJ
d/ZhPHCIn4PIyW75bbPgYOdqyTfzCDWOh0mZ7wrlXagILLDK3X+X73abkB9TTjUx
E6hhZgn/YSxDsDamSNtBY0HxJFP0uGSb7IUo6X4Y+h99OSsonpD+z9W4o8HgoLOH
BxBiyTc98UwFrr/V4x0Gv5NYEOF+2tl9tJusJHh6BhfxQ1j7ywkO0csSOHxVWjEN
i3uHXnh3cMZSBWvKP0AD725bqh63JTWQlYqrSPjLs/WPlJ4oyT9tiNWi3tNVJ2wa
hgq7AIPc27hjvDnqvkV5l8+P5W5MgpK5C7ndFtDR9KmCT0jqHV3EslY6jfubHiAb
0EQFQTYaAGNIb1Oofp9iQi+vMIegdECCmk3/SA/Qdo/nIFHsC6f5X84X9e7p8lVr
IDhSwiYsmDE5PIiw9n044i8BltQv9Un6Q4vafIOn9SgmIdt2vdHH9aupcoYKoAwp
MsSxXKkHQ4mQsDVrcYrRvT06FppFg54rBHnCQwlVuDG5jJILncnH3UmCg7p/9ff6
c1s4AvdW3SsDWNh2QX7hD5F+y9ds30xtr++0PD2T1ybjiRv72ABpdrlc+6EeJ25s
VarQlwzxJ7CaLwaRSWV4WmOapTKNqaBD59wri19qqqQJjxuNGilG0wW2o7sV4hJC
hqHZbcToxRF+Har2Qo9VoZcSdlDWmkDodFBYdy2qHPTXUfmNC1/I/wMT8W0rLfYA
XfiNKqetKFGP2fEzxcJlkMfB/J5xHidjdP/NSH7PrLxlamO4bsjQ9x48dEEnJPEX
LoYSknoM5a5/1KQ5t7g7cyjPjadcTOJwJuCnyA9VOt1lMv+ZZXefg96q+WLx6tEs
/gwG7qC9JgMaqegF2jMJDI+rXrERJdkwIpdCEpgra7VQueiMz1bXtwBkif+X4yMu
tBuar/AkVlMEgY2Sre5BcRv9P0K7n7FhS1XMs21Px743g5a7su+uQawWReJ+kBIw
V80noZf8Vgd8QWqdX2BIiVtxhDXkNYVmcv+Uu1jtqjkNjMPfthFVGID5C3oyQ3k+
4HyH1nz/CrLqxzB2iXuMw58hGKDk2fC/9ooyDL14YnNdGqWRwhVHVezRvZDUa8TP
42YGYg8pu326TEEjC5sVIlBajRaRMDv1DjOI4OyyFkhkCu7trAom9yjStqOAPs0W
mt3RJ59GlLJwQfAR/lTbgwgXQRvP+ovmtYWb/v1FW/skpkv6e2s7NrwH7Fc0KvvJ
ekj3h1FWT7ke/xl/Mmoy0IwFBTcLtPXFbdHRbiAiQ7JfVzZQPdpNarUsRozYmwjd
Vpogjz8d5eQ8y+MRVcEwAjIzSzjFdZHKv6Wk7S3r4o48Wb4JVrtf/B5DXKLVfC9P
xU4uj3d8rwhoxR8y3AXC4frgz+6Re2UpkXK+x9JOyfMoaKw7E3GaKEyZOCnpv4Pd
98U8GIUvwaraKxeb+HJiC0aS0MyETJ8a//tIIFtr+1PzuMaaj6D4FxCMv0OhKAPe
qALD6rZB2v/1S2mbNDE7Mn2cFbswOKoYXRcqbvhwETRlnQHzL7GMLpxr1wbph05h
tz/NnE8vM5ymAEEHRCZ59wWIqixEWJtIqPJ4VcFhXfglct8wj416hELHUgcM7l9t
LJUJDhmHmK7qvduTwoynThv+8mNfs8pNh+vP4PSNlnK4rTKpnS4nN0t8JT4vuzFU
+hBy59ZHN4nxOwmtZ8Fefxxlx45ubYDn26ceUlLPbp4/4ZSHaKOvDNHVUqdZM6Ad
2OokDzlkYyZ+r6kqJ1HQaGeJ749T0IVy06kbAD4J+3kOTq8t4RfwYhESvR6qMbwV
nxeFX8bmEZkzQ32Ugyj9xfW2gFLDJBfrxGTK01Ti+8TS6qj1f67mlBxowCukNE3F
AxJxTMXxnum45SCduMaW1C94OYCP/9hWT9aCywGf9LoMBZ0S2SIyx3vKdNE9RuZ/
9InczTuEIDNNHK7Sb+fxWvANXkY2uKeeppjiBShtj0hqoDozeRQvqXjp9r8dbSIw
GIZVRubIKe/s6CQzUmj2bJZccGmQEZL6ZK8n5uKzBZqo0s0nqTctCDYoBBKfevOe
TCd/5qr8rDml4vC2K8/REVz9vTzk1QS16O0AyV3ZgrP3r2BC6zOP5QdXJrTONCz5
FiTgeL3b9xDMh0wjrs13iMOlq7a/3Qq9WzK4GeJ0olICtJ1P36RextcqlAS++f4C
gIx1PDcUjkXHDk7H12xyYsTX120KbnDcn3xegRXtT62pVBgmpUNfiDNExe0rpohV
WGqu8cTl4QdVadyYPDuj6ujy85YHiHF2PDNYgWebgyXDxfBHf0d7g+lCMzWE5Rd3
4k9nuxA9FMXBk9qt0nqAVsGfpsAOux76TgYTOcNE0fdn5zxcRspvJOFf2K2FUFG2
lcOizbqCEJmyCC4nhYVThOosVZltYIf+yw37u0IZpAZP3RWfGHy7sL8kHiHILLHf
9XkwF1oHALQpdNEoyP1eM+HNb+GVsPpyGkYPjvavt1kJFhmijGQDNfAkFE7EW8uR
7HkhXhUtHKFHxkxGahiYlEXXOgedmOvgNq/fi1zFIRJ41GfnCuS3Xw3Dpt2RHr7A
T9qovtm7WM6h4AVepm9kBJSo8+xF5dujlVXrp+AaYLIWARNWddjL31d3Iy5zT7lj
Tp4B7g5xll1rFfkGVPUFuwktXbwoAjtp0vfrLsv/omRJcxqGjY+tA3X4JmHJ+tkA
01//ZQHdhde527G119gdbJETYqm3lEpHunYk471BE3DQpZhWNNqq5LZLuzTQODbV
LsdWFteUzLK8eTvCjdYVcX8xMPh2bB026bx5/uHonOEIcOYEwJ9W6UaxbYpE8Akp
u0ckDA4uuyjjRpHlI9HlTaTaNRbWQj9ry/VqQZQuIVbBmfFZzxL4y2gMZqm+qAPN
EKOfL5ZIXelY1CACNP19GPtave3vIuLi7bEO63PuN49uXWfAirpecplLbFnLRVmp
u72IbhX8RvAvsqrBiI9Ztey0zEXv2+/hdcjyQ8DHjTzt2/RqvNzExavabwyB2XQn
EsEzyA+J/Qklf8rWgmChlUDwAEeYgvl9sOXbVazMc07Yj1ZxIPcPsvHDIWBJo1eT
nRZ6cblBT5uBT4ZX7hDvJt9B7K7NYr4YIp87wmp+0TmTMt1qBSxLklkFjGUEq826
d0HvZXRIwmitiILcGCFlD5xxAM4BmfIW4oWYspomuR1msMuYCIa7QXBgKqEYecR8
F/vuVfohuiNqNN3CDhYRh4mMycgkhEknavx2AxQ4r6L+av3mPfm6zN1zWxVl6VIL
RFc6OZaRqGQ/DsPNf/QrcqSDUYQnQRQnbuqokfLhNBZuG59B7NF/AulFBR8PVDsf
8+xz3NP8FBDdAMsLanjj0YsP/WtVQ0TTnl/vNazZNqHZjbiqFFreXavS/CFTAooz
ZfHNK0YMk18IMkdiSC/blJZUJSpau6o/sxZZUkB0MN7unD8VGlL6M71jVY+kbE2c
ZvfF+huKyWPGtehyO4xZ4Y89c5xN+WS4zZDiSIX7CobDPVMHVi/CUvcVtyBONKD1
adOzI55UN3AK9BEL5ptb1SU4HDTJ5obDOp2aObYf8i0LdxauY9SqfmoQHRN7ZwAh
0BNsiLwxFahI+2a3xKzxbAyIyu1wv9MiINJSGNIZsZ/OXdaWLeskrB2/nZtM7ufX
cQ121DOUwizSFfr0DPO39oL+rclvjsySBSoe9l6S2Qa1R1cYsM8T6e+/QoVqg7yB
PzOz2FHa0C+560O1FLsEUBOA7IFKlm+DlibHSdWSWinezkj8J3NekcgAutKYykUm
Tm+VDMqYoDPZozlVWPA//uabIxeSSk3Eh0fch2GYZ+cZWnx76Kl/vmB0ZWR5sBcv
pyP7YhomxasZnKJHW597tq1drf1vVRgZtKM8ywRncQU1r/WdiKnjLaniPIY/FylW
l3IE7IXVpWQSvieDxQm7zozUvKfrh9SMj3dFz1a9oH0l3h8gaspHPRSbahyM97sG
/aLOsQxlmE9JTdhRV989LCiAj78jt34Uj+7WmwpEaODDResDyKGIacP5VYawjt/l
iqz8WnefkmyVMFPhAL+V26OysihM0/FwWXsqUVc/IB9ZRfGgaP0++Q3vWKAbRcre
thkw8gD0rACHqwhxkrE4dag1PVokPA9Ieu4c/IjoaonVjaAlqkyfzA9acl602kHe
+FYJDpjp/D2bEv0XVBN8R8ZjaOgrlJO7fpbVZKJ1Ben/NdjWfc+CZfbN7kXhQc9h
5drrzFPXviPEVoCGcLqtE+bZMcgMZJqRNOK5dxZtWhoIQUX7vZ1UaaHjMnBYKspu
8/Dy5PJmqBUAppg2Lk5i+7HxlrNW9US82swDdLhU4wI3ti+h2/gXV5Mxm6l9YZKu
ax+Ddfm+mVIUqZteBS413JEu7EouDtY6hdOWSjvauGYVXexvihrNX8Toefhm5GIQ
hgI2Zh5ts3W0dxsbEhQC/bFnydF/9GiMy2nsAw3Mn44G0CWSpehqG8G57n7BZ19R
NgIU10zpReV5SBCVAwom5TQuYPdEtrxY8/vqntRE1+dEs02gdp95kL08YwpT0Qxs
I8BA3mpHmRzbEEVJWgdv+Eechlbg1c1njA6gHsFdJgQxuaSDIWrPXDJq/VYKAthx
ALbemWNiYQf52hcGepJ4mOPiKJYpXA8B3+8tgDW/gwKEkEDSsLKrXbS10iJISh/1
+zQcAPAUINsNXMiUiWqLuw/gggw8Qj3BEQy+CkGbcCGjafuP748cNuUDqr2WK/cZ
BBU7kiEGQ0RxqttdmTlnlpWNdgP0m2XfoUi+SqeHCKPguvZfdN7TAybj261uOADN
eX9kLMvNsE8XoqUaC/Q9PxCIG6NrPX8Zv4a0HQOHboGZI4L++hTgttVJaGal53FE
u1sAbHRwafDC3m9Ya/2wI9sL+ScDpSBxSnJidTbSpOrY/jJa3/FgM04kYL7TOtrp
ZDJysvZ16LeiosM5iAKJsHAtZiUuyVRplMy8jzDKu0/SBj7T5H2Fs3vm72HWq9op
DLYxfmbStZEk23Mbiwi5ET3y/QVT1q4OIUDFmvspaJboeH/ZfMjejVMYvJGBhQQT
NeAj7lcATJEeY2SAJY0RfKjLO+0jyosL546v7zWVHeduTkdZumc08jEWBNCTWNOE
3o70edskudjiZdoNf5V7bD/dHjXxrNiVTauD1FK0DOjgkQbNMG4voqa8S4loojYr
6XwB2X5Taf9f6hnNQWoWMAPROycO0HFs2CxBU0AGCWNvO8/95N79HBODW09q+czV
jPdECCiuhrSfiV5vlaLOvnd/bp60dUifh1l1sHGfFnXprq0WmhLYpeMIR/XlEYQq
xRMuOqN+y5W0216cu8DY6ZQaHPUbu1Opv8KKuLEi+dpOTadBsFfZyp+WZInwgqeO
10SASmtkAALfiwiHFb7p1kY6tWRLZ7nMnbD033N7J8lEmShQien83oUTxR1QJwlD
TG9NBfW1defXFlRj+JXVsu2i3yN09mQ9bM/Ob5bXep/VcTDkdDNB/Tvx6Wcoynkd
KVVd+swE7jllSiO8knDuBTiH0zvJq0KV3TJqpfTGA7msf+RPAHPGYyCToC897QZ/
aFHLRyBLZpyyh6y1RRFwvULFh1RqyOaHyj1ofM1PnXwRwtkQF1VIAzt/1VhKKmpl
XN4lnlVyE+SJVKwyMP6LUu9zpUy3lgW8tE+1lAFY54Zn/QxHnyJAsND1mXY5TJsf
JMhhP9hMZVxtQm3pA2DSgRm1ZU0xw3djsfTMmOCAGLAJm5qGflyX/OXJRw28MKQH
us1plN5An6c4X9c5ARtkL0vZJ5WJE9GfRAa5klSt8PkEPqUqQ89jzQ4oPGIlFU+j
rdlplqi7SQ/Ewzbx0A3qBVPxadOa/O/j3hku4/nOerQvUIVnIfyaG+iEGiPxd46Z
23YORrUwKqD1/mTNZOldJFql8k8qLFbWKznOeHKN0Uaudn18Kau5DqfHQwcmNy5R
2cufy8KvhLeyTTEjAtQYGYLB6x5bR7si23H4VJqNEq8D6ICaC29KO34MDV6MjRxP
5G2bsOuZDH6aAomQzRfQfVisN29jXct1Wpn3V4h7GjksllGQkJDEvQ0LJRqU3jgx
WH5v6JQVe5HfUgGhhGaA180feLvKhnwamgh5hEQNSwtk/VfPXpqJX2AS9eZmo/2J
J54feQKLr+zEJDWZIWd+Q9FYaGo3wvgdCeMqmFx9diHGNINSGlQM077iyBoEP09F
AvzqLNgxP6bBFGKBIZkrXj0V9/BBBNEPtUzaMUfwB5FiiBGPhKhHcD3YlCKZ0NkU
S232wBPLbEvRITtZ4oA4K7QIv3Sq7Sf8fky24iaiJwGMnfkS22GldwZseUVu2syh
kWwse0iCHAwjis72OqoQRaMIAmqI9ehBJsn3pbeMBnBEzkoUslfvZaYOZh7RtxNN
yJT8uDFy3S3PM6+y2e1j2E+53YVwn/NeDj5xkW4qYzNKq5pQyeNTZJq4M4zIqh24
WncT430t3eifmB4h6f9LSPrMK/bzv2bXV/Y7sxkSkTHiat+J3JeetsMzMJObGDEJ
9ZSlT+e4zQCmMSzyCblIqhzE0qqrRj5UzdfCmCrDCcWLjkW33JthRR1wFc6uF5e3
ZwSUq3ubmkVSK+hFVqWsqEAGn9JCtgAfwib01K1qIFHVRV+Oi0mmWb3nxJTG3Ddi
IxcVTF9eqrwv8O4n6cM6KWvKyEZjOEspVKlG5R93XJLE/80klMdJHGPEZVNkjwDY
8FdKpUR57yz2yz/8w8uINZcFhj97W+21pSzFWw8DlOE3IVNO1D6TU69WCW755UIM
CqJikvhubeA9oYPg02eAmKPz00s9eXyDuwJvETgmax5pWtbNRDW5U6wu7POHA3mA
XDdCpf/P3K4q08ta0Ao+GAUmc57eSKQoC4Ykx7F8PwKlGHgHSRy27vrSdpKSeFfa
upRyMYxZ+hlxGh0GbmJtt9yQ1PUP9uu8Guc62fOGwogqfis1t4FljTasxrvMQGQ/
NzeFxzDcox6EuukU39Obcbvz2dIMXbeyEfPbFGR1/74HUQCINTu5di2nk1yhymn8
ZHm2l7gG6Ndajk6GPOy7RmN7F6eZfmbxf+lfnJPvzKCTapcMzZOsxjuydidYCYVh
MT1JQ7+Wgdh0eqSpQmwZhnnamqSNOYuhja/7/svbb/xvAz5KG30Lt/P3alKAYbG0
TW+w0KRILBZXESghVwKo5KWaWSdkjbB1cO93dbm40NN+vLtw1KlOxguLgx4l5xAI
q7yw1BnTAQRuBmhQipzH5uM95L6QuElNkVv6swsdgLHz4nQBcby27ffNtKRXt6ij
4s5uz1ytcbu3D+WUFCxwoRhAkEyHJ4PhXX3HmAYE0Whw4fAoAicR+EgfYdz7u5xm
LO4cOgJ5XwRp8JUa8KJncIO1Fa/vBnLvYt2lrwr0VzEc6lNT6rF5VtSuvT5TZckb
sSLF5g4m7gSAot/L0xan1Q7JG5pbt/1/B1iNKFtHeaiP7M+Svqd3jgYCJzMOI0l/
4suvkLV+szdoT1Xzx7+ya5mBeP+JCkdvW8SwqePZqWpNqJwxcd+lAMQQRqrinUNI
mfmaORypVxy/IFvQrdBgAkAj9b5fipYVHyfUFDgrhL9y8jIFG9AXWP+xJwMun2mj
eQ9QLrPOPiJeZBBB4YIQ395pyBa6L0qH4kxXg0zoXZgL99Q58T5O6evSb1OCZb/b
v/EvE0+ILyEpqOJa2Ppd17Z5PxJGRGDBctTXPWkTegdp2TFCH+ySxE2Zw1XSzAq6
5wG2NHdUafiribVCjlFTDveEilamMmn5RGMJhK82xz04ULclRZDo9+qu/cQ4dbw8
q0XABX2Z7zNugA7C2dEv82VwrFMUnTwmcJ7XovaIVr1edwyhgXTCPV+1yxAhrQB/
dq2dvZbCBaQ3UHPLxL1+vjQ9WgizLU4sJ2Y/VuaxOkxYMAXn6URouua8gZgK3Qrs
FVm5yQPLx/CnXXzYzP3Tj2PGWdbKsS55HP+OlHGJxx6zvEt2C3gTbn8iI3kDJ6/B
TfeKd2mlNCxPX/oGt5qlJSyDLQ6+p0li1qh9RY+9TA1DotJWylkjOkSIYtLqJVz9
7djkeOxWK+xNka7hfmOEoBPesg5A54qrBGfZhIS8FS0yq85cxbtp9w+bI3kJMJ2q
LFZcY5S/GtJt2EyCu8AXdv2iG3zb0FRpnMTcRQiDPJZ8P57hjTpMWvgNoUGUHv3c
lUnDLjijX7oNUKByyYJAcfjtZYjzbBsJB55mkqpIk5pIiTnsY2wxGWt+m7mXWsEG
+gtVBCDm0aJkbPjIeYp/m+njed+t6y/DM8EM1F/YD/DWi5tverRW8E5QDbK3MGWh
VSlPz+yPvkhMmamrPWmEsgC6ZmEkdKdUcuS6buLi1QtxGolnGmthONRMEpVZ9y8F
7CpLVovE70EL3pEekvPYnJFEcqB7n65piSfzCfkVbWqSK/sM8CyuVU29zPR0c8sM
0lBsz6nLevLnotSZ5Xa2SUfpdPM0rxNxTd0p/wdaqRec66SQwscYXp3SdhvsLqoS
vvEW4p0YfunwzGIkaxPkmAd6XmbYed+qIEMGQJZAv6sOXXbrYYDJpHOUIaiPSUpK
r4rZ1w200FWAaobP8HITls0zNQHWfyXp7ZYn08S+GfutHWzPwH3u1t/UP5VIeKzK
uYGkGrB8jt7jsnBaV0E3eRlQFf92TkJXkEjScV9S06IPLSey1IenJhPfaBHPuQ2U
9NTAHY0uDeiSS23epatCfj508AF89IUl6rd145rjYtsAw05dt2lqaxS/qLMtAAkG
B49ZAoA8Sayo0BYgARlBOADCDBzcR7+selzEYIrHPn0wZb0Of1VdkuZXsI03SvaR
DkvIGBjY3B32xzIwWwaD5G6l1XXPskkL3XB4m1bnz66Mjw9rPrSA0ioYT9/6gg8C
lpd3H5yUZ1cQWTTgO+f/gFUZqXVa2DmSdcAivmyo32sQeQbVI+2qWvZ4UcxaKjZ2
gR/1II+IQcaZwWMqm9/shQeSAlq140ybnUl0mqghLumUmP9YQauhn4iAtoEpMfhq
T8TKaTCT0V7+x+ItgQWtSi6HYELsvGzeuwxCWwYyHJB1sc0cRz9RJzDLnc/lmnKv
eoA/I4VIOUFAVc48x2xVYKk2d1Vev3ppQF+P0PXsfNyXfxPlWhc/ylc9JK92UscD
A5ZzE0ZuSmf7CBc2uxdqYQpD4XVHIP/4DYlh97g+29zTlP7Y+APVJfncfdMhX0mU
5z3bTAG5U0aA2Rr7PCADMw2QB4HQLCfKhj0JkDugEiVDdtZEVlAqjV2IVx0RZUk/
Ri4nrY8sNxq9NiqhOGdXIODiqANlukCbAawFI30fh33EagypStoi/4X8l3dWxIBA
Ng1O5VGwsMktyL1iqb3OYWy+JqwkAYgwXgK2UxoDTEjnz1ZUuhbdIWxhaua+HWZq
2zYmzbSuGWscONUT4xwZAkS8FsAtZzRlvEhyKm2940Yv5RVqLVIRgBDg2lme+Z+L
xmO4fbTTWgd4efuyremSFAcwRzGojnLRvSpgbYM0FYx3ILcQ6LEzW3JV9btFVem0
hQNOjjESm/wE998Ta3yq9Bt+fpV2RXeiJbyM5Uc7EtAz6hEVl5wA7KTuk28mJ7oo
3lu3+85wXlyBM9F/WlUFzBC7cvYQJkfsXRJmiBzQoycy+rvMXLdw/LFOQi4O6rpi
a7P+auauRuiFxtFrNGH3JwLwNDr59G7RNqYILkTFePfcqikE/sNxAgyZ7KW3yFW/
hqL3b6jTsjwy+FKIrOuv2MoBJBP+HQAHVOKBn9HN7U1zKXsDG+aKl3ShlfU2z1xE
xYjFRasp9mVY9f08tr4sexbCaEYjuoy8oy9Eu1oEH8j4xbFLnNr6UbuTWa+EJTMf
JD+cmyRS9NJxwEbeSI5gswN0BctdVv8LpGna6Gekytgyo9y+QGspJuiYcpfpy/fi
9HGpA9K0NjiJOD9LeMiFFIC4/YT+QbnF+rd1PpRv8OBoeRMzkXoLkPUxgvoyocI5
TkHXarkXtwW8HsiyHFpIPbZN0jq/JVWX6nNxD2IXf/S+nFF4Prh2qPA3a0H1fm74
/RmOtDO80pW/AMT3Jjel3M4ywbIB7kZa/6HPvHSku7K3Jnr5LDZu4u4tc/uiXrRq
BKDsvX4S7SVMuWs3h7lc3rGCmVFLxKHqdQ1ln7xNzMaTSSY9seQYWv0LntqM8i0v
5PIE7S7dGkCnxhGzP999ntStd2Jnl9Rijfwc0aeKYM1KRsyZ1U6XvM9ZaHKNDqid
yHzrMi5JVJ82/aFS6tyGATVqI8R50MzyVQ4rRSWnp4fR1mNO2TXsrnaeJHrNbA0c
S4C0AqdAyI8Iaj4aIS+BLZcCtW+7sUj5bmzvtjNRMEZnDvW4SN7LrylqHECzbWJk
58QdzyPch/3q4vBpM/ulSu6Lzery7HhwDq4ZnMUpYokg5wCpH4NwZoFvWSCzxlBi
tgb+zHuigb3AEfttDYq17J8WBBOJ7CTvY80Ihl/JHULE1BHe5kO7RnexluErAbo7
ZodQKLpczqMwjSmt5VrSirRt2ykG8y/GoxCSZbkuV/z4P0h50pc2RtW7nzvBpjXn
qFyde/q7ZmNvtyQP//OxSMdZ897uUe1dxfjq7qeiBmNQM5gfcum2ID4Sv9M2PK0F
Sql55f9wGYEOXzqWV+jCwUm6EHn+ibMvKI6hSmBWJ/ZcyYllDNO1j8J+W4pHuuMs
WOyIMcbf5gTKHzbTPSVKhSPKg1wBww1OA8B+ezrYphlx7oJ0/cNQH3cvt29EPzDv
Um33eL4EscNX2hlmD5xc/ugGKVY1Qbkb3TBLufeppEoP4W9+5Z49H/5rrCKrkLGR
k2RjKKUti7H4kLwK6FY2zuykEHo1pLHVYawV5aeroVgYqWMm5yB8vqYkUT9OAvVz
Q89CLjFs1NCsFcmAu7zSQ55wD2AWPlRLnDMrtRtBK9F/SlYVA1UYCI0ORcghw9dg
sAa0QUJFf2scmNYTuo5QXrzU+5dgwP5aScko/eAL0TriuX75OuC5wLGNha/tXZiW
CdMa/Ek/ZXbb4x0YFcjrncOtXMA6LfIq2ASPA9JCXtJGNN9A0diFEM5sXe9PYOtp
QBuvRwZpWetI5PN83+aR/PWwKAXBUGgHE7X+UGEb+zTAciCLEyf56dNJqcu0GM+8
d+PApkKEEqgZ0KH/4xbG6aM4zPuKWQaMMald7C83UvJIl/2zTaJ3QPToI6xINxZC
norIshEjZDmYv4DTnbIRQbIl1fNo+PvjpBiNYjkTGgEUbOhiSlgXXAY+QD5hNFqw
3Eg/h8Vl7x2hlDDpmZt8ltQbP4XmtYIkhi59olZ4QQaQ2LXFKKGrjShVl0suitVs
aaYeMBU03kdex1Aiaiee8MOJ/ols8xW7zsfIrVpfuqoP+NfM7Xu/1ItR1C2t6iLn
Hw6Qq3lX4WvhNWUIl38CgHHxEhSu4hXTXJKMkG0z5Qhl3iebCBDNvkki6BlbfhFD
PWgyttjtXNaZmnrtF27/V3AIZj6t+q/DFa1PLUsUsDJGPyc7kH/BIZhXokvXn2SK
PKz6EoKcyg1mk/jvg7zphGkYGsWo7JEKmtz/THijZvx5x4bFneYAxbQvYBPEnNQ1
cwrdx0Lh5ilvuqrF1bzuvqYajZXRUpqkC6QyOVS+XwkkzhNAXTnu8QE+UmQRmvoU
jxVz6kShdPnxF1b0n8McyuI3Lvk+bL6eUzv6HyFEJvrwzpTm4gxEmvDG2IXt2pY0
lqRbidnehYaBwTAEdzd+eehr7QYC3K5cxXaO/hVwXg1KVmpf9g3xSe+CjneZJvVr
rSMyFVNEMH1RhLlYGN3YA5skObsHggMGLjAk8KJulndlGCA//1OEq+/Ks17h6gEe
UihQWp/hxgPK3nq0cMPUsRiDIZ4WIR3goI3tJba/X975Ztn5/IkQvEP2GmIWAuey
5HEGE81aJvzy/f+omJOM+NArs3DfsTdrE62ebfhWSgpHlWGqJsikK1RcqRIenuWJ
P9I67t5U8NfAf/wyqImaBd0fr1vpxQDJvRFBSjQPXU3JofWm4VHZkY6nkWAGznxp
mFxy1XgmAx+SYFbHNvQ5uTzTl7Ef1aoreUlQNBXWrUImV6EvMwQ5cPnEMu4WdPID
r6ueFYnPoCKLvPZXa71qT/eaHJtsuWvxwIFIWEYxZTT6cOdhDDVK7Fs5eikviKrK
xZtHGfpG0nhWqVpqK5KeaCs1f02nywyFBqMSgze7/DcfzDEP5S4DxBhrm81seSv4
I2t5lZBSSChRM5jNV8a6fCXRiC53/CnoTnTihydashxGQOKpx/fcCNRi+jHbA7Di
SreSmTy8tP+WhPjQKSntJb/2oqvhH3HpAJeKFhqnC+uR6w8HgnrsVKalrzL7jfsz
FUrO+bG73NnlE0LC2XkjWaVIvP+1m8dEuAt4fBV0JsY9/ku8aytvkqKdJ3Ar1otS
9nYJCM5Fzr2da9smosCYNlQ/z36sQDF/GmXkLcAdjTbJoeP5wVzfZa7+H5cW5ZZ+
1+XxnU3YXwjxmuZu5MHmtE2qOlw5Kpup59YyxozPe4weIo5oNLMnS3PPgQQRdyB8
1HifQXviJOmOZcLpS5vUon1g9fmrerNSnu43VEA8dUmEuqzAi0/fsamdajVj35ZQ
UkW6egANFBgFw1zaiq17e4erfHZ4MXYezlQ8lxPeghXkc/06yTHowuCYdUm9tbWM
236U94VzII+4dpVjtibPwrnqD122BIMaS0it6KhCT2n2pmKawx2uDzriCfJA0T/d
RK4b5cLGTPp/Q1oViPA7IoRrQDVAidPhciv+WXTbbaMzzszOLXnvgaaC9QlnFzOH
UC4yYEFHGufebtHdq6AlCDQ5QmpDKjAhUC3eA2yw9SuNCaITsIVfaX2QL8qguLpI
QdOovN7Lbcz/OdfIWWIpSZEelQT8igDRAIJmxmb4tG0ffT/rB15jNi7WQfHvGSkD
JXeXasTrGyC2nKNjvwY19vkQSAwBTCV+irzkXl0NtNdbeEy6jSeuXUFsm6Rj67nW
68tUm9YFQq0MEjgtyCcaZO3BXg+RvzyWFR0/S542PrmqHW++fuPnHxrtc8xUA4MM
zoDowhtb+9TD4LffFuL6UOb/QymavtsIQKID8dp0gQTsZDAifIpf/Cvv8dPCFa8x
GDdBw7JAILWZ9YMGPNFmk5wYUnKbzZ78d/xEz9WjOlM9+/5zesQ8K3C1S1xnYnbT
Ga6M9DUMrMRcgk3S2+SsvH3ZMWI5AJS4ZwmiWkzYAKbGpoeMp5TcUa1drAicMiVj
XKrxwcrsx62gXoyqBX13Tt8Vwwe7gNGPIespyf755/HeY+1q9SfzSKfaYee6odSd
Vw7VfS11ldnQSJUy1DobraHEi2+e9+sluhPFP62DHRXTgPDZypPeGfdqwq9HMp0r
XW4t1WjCl/ogIHd67xPQbViawcwlGfbZkMPwI5RXICIVObjqO33bRRNvG2/sTbWh
8LBOJje9z4iY2a3zxJ+2qw6hbC31zH9eMLlI4bqVYVttN4ui58XPrWZiHehwl1PC
RKr7agLVIjWgPPOG922OPsS1qPa1CyYXLGwqMobz/7nwSKb085TXLA/a/bf9RLjC
dujf8IhYi6OcE2/PIxlZbhJH+K1Vz0quhAKBRNLKMqA0+LJtGYOnmzlHcC5VyzgE
vr3BfLdBlOKo+YyS15SrOnbRD8mPQamyjbdJOEw/gWniLEHfTYfiBC/dtl4cUMqc
zWp4tfptBBTwQi/tC1N8Nv/TvK45nzmGGVhHGoKq/lhCKgZ12EhkUWViKyVgZ2U5
UxkHtjX8804EkW7PZ8Ovw90vktSl8B43AEc7i+bizFpE2mpj966/Myulu2qbMxco
7SyZSmCkbsU4yonXScVZH8jXx7IsCqrYas55yG4Z72G0egh0vb/77Wp1fcAHmkRX
P1R3ONT/G7l9d55st6BIhoHTvBvx2Ao3WiJhVMd12x+B1zNra1y8ejaB7rGt274Q
fWBxZZ+uXfGczdFdmMcwcw3TLNNITIvxS2Vk0wkqkkA+K7cJACpPQR20ZojeFN4n
12VrvLvQzl4OUavlgqEnKiZMDJQhctaX6lNd0RQT4dOal1SntdtW0I3JQnzTyqgQ
UXfy7+VjT9SXETJSvEKbI78Rclp8fwp8aQbdsdE1PU5SlRCgZ7+rETrE6eDdT+xM
twzp1tCGA/nsSbSgF3sb5YZA1MZjK7h/7egd+DCCMS1FzXKK3CuP0bn9e5txKsXj
L3m1PH25Y13ERaNoZnUBhzpacv+oE2OhweX7FhLmZWaCybxkhNYoxaczaHY469rv
CUUVoL1JXvY+Cgb9GPhU/APVWzN1Rdxf+1yndi7N9DuNLMvP9Ay+Sxj9i77Sh7Lk
My4Lifi2orH8Ck1eFNduVKBi0Q3F6wB4PmRMAeefweFOG4PNu3zJHvtGVP6vTv8P
lwOyyHNUnUGubOwtih3HFz32bLe1Ad/1ekmTUbtfeeyRr+b4FIvKGNWWZgYemQBU
lzdfCC2KlX07JqkhB6t3WHdv21741DeV0hOr0MKYFa9GZGckDRgQ++eO2UP2pZPf
aeWYkpZqdUxdtZoGo4DwoQK4FzMCncM6O/NrYVSvNpNad/8f/OdVnVKrJxmWfJiv
4O3401f/CqYx6rI2sPgtybbuSGx+qJOYlc+IMOK8VEepi3hhvTahx89Ll14/2JqI
Y1vJPmRHTaYyxoYebsrEkvhAq5VFAoLFh4WLf4KhpprRnN2Qbb2UDHZE6aiDFY6v
8Ex0vee2cx2yDwogTPRAN06EsSYUsjitaorIBpOSlNdfjpz7auq160M/7cqKQSa2
MuHsczj8+Kl92/Jxagodzjd6hyPe9zXHtfhVdKr7Lz9uRR8wVfLt38NZzizWrhVq
iT6kx7X/pmi/aYUloE++x7ha4B+boh+5dEWj/aPU5ty85prWkAKGlFdnEXFxDUUX
haHMOBGJUrI6z9b49pxZ5eMrbMt9GC4SUZAeYIW3dTo61Tof9gGvEL1fQL8b81XP
PuQy2Q5+WRz69rfB0PC0Uu4dBKAc+V5aym3K1D3+oKf7fuWQd1Y07WkrX1YgY7UE
fdgg1aMdUffxdp8D2gbJbYuGM46mSqg6gWj690+Uh8Xy8lflYabMhGUKGkO+4whD
ON46B0cOEbWemnwg8twdSlLpbGJMo8WoSIdUimqLvjTwIuDgXYRNTFXr+fJRjxJ8
e5c9J3i+LP4iGIVAdUlMyEE4O90Z6snnCkkIbueK+SPLnTV3bnE/xa2mLB0056iq
vVdpF+wSfDTx92CnFd1Ab/qtV649VRakIruHKa5/+Cs84+K5nZRtgqT2q/t0yIfp
ePX9i91fhSCwaig/Tlxlcxw4kUllwaTfKhGBVlNZTN0e4mFfWSAppD5fS4rW325m
CKOdavRx4iA17rbYrwrhpkBFF02v56H1FwmtVaQucteFxBR2offcBIO4MQRBkZDV
zHKCiQENqwjY0Ic0CR3jeUFYydfGoJkdtuTaLG3ti1scm2yYpgRzKIRe0oNK26wR
nF5xbN4zCKNdfDrwC1TYkTt2+cLrYV1XUoKHBOZyuwUSWL3qUoR8RAl3vuSQfhqR
UF8hJwAUiG9k+m73aSvwy4DjNXHXv2j4VjgCvOb5pBc/eX077CyEDhyl+NwBtan0
vYVpIsjdNwhpaSLLO4uIorFcticW6S/CYGENPx1fbZ6ck0+ataIKltfBFlq7QOs2
W3SBtWuG45hl4tEfGNxp50i3UJ7tZ6Voj2YaD6o5h2wSOhvFobxPCQkFdiGXZ9N2
xfKRUIyIR+faIyG8l3lpEQiM5b8OpHjGWziCKMwWcU2VJAlNaFwdetv+h2Z5Zwf4
CYm3pF5+A4hf34Rl05z7GLfi4AIQYphzoEQFMO58Zl6/2Q/+SBGznTGBBOImbokz
NPXq/Ex7/UcJiG2UmRKsiOYhnUa620RzRnGZgsJSzkyjQShxgzaTh8IzdGosNHLQ
tsXzxW5xuRdFbzz1jd981IxZYvYsYQOwtsP12SkeHYLKXnfN9pxT6V9R6ZrRJuN4
v3IalwRxpEV/LgiD7XdA9KsZc4hxFf1eURqPkH8GiI2FErMLzinL3CKUiy97DF8H
ERIVUv6YxNUWY4w5nJZP2fDaUxTs/GO167Afq/6DmmL4ctZqmqsWA4UEPy3ds2sW
gZOz75Qo8ICTrq21fOBQVyZccZ9IdFaQtEaZhqE1V3vAAUm7VwnTAxFOWXBlSrkS
3sfsUjBdCD71KM6ku/KLjicbnJrrpZ8r2IvIWp5ik5jcUaLxCiRGfwzu0qh/Ooe+
igrl87IucmlDynyTsZ5rY6RNxIiNMRsIUhkmrZauXTWheVRnC8CvaRe9nQWMDvO6
LHW1pdE5n/pkrnOBJJqmg+5YZPEZvTe1eVS51B0pcWsCCRAV+IeJgpsW22Xcj7nN
DOB/8bXzVAwotfW7wHV3L0x//zis4DL+I9gX8IpeW54uAjLd3kdNJ7XSWuWq7rta
CiXUUd2qA6SYHJuY0gtHS2oibX+eZcWmajJWUz3enQEJtr4Vb/HJHvBkvmWZUZgT
2pNkc6/MnbqYbLMwb7aBwPZlmVkpEqhliWXh/JnNVf6FmH4f2qoDKhcKJZp0gCZT
Lq2FsWqA+Vs0OzCz4zvZabABBIEbmY2UClTcLTNbqWbOu7J3mHhUQqlAf1FneT4i
Ddtot+FIg0kF02/nFsKo5gFS/TS9fGfEvQShIg53KOaVhM1XGS6DXopWACPkAmP7
iGSWd1fPq9GrgNPnOugDHFF4EK4S0Xo4LCQ4JFBrffPDQ8HUQeRc5hTSO72vL3xH
tHrLkD99Dg5Vm/05Cc6MHYrePg6ZsukB60Sbq35R0a+yIpMOoonjlGFsZQvhTFRg
d8Ik9OiJsbZRYNSx9L27XauruSStEY7VyC7AS+M6hghl8T/H/JG3aSJnQu1fPCfC
7uRCFgA2QMkSbm+jA8NNIkaBgBYhAxdFCqGKgTqNARs6A4r/00ptteNTKtSUGmDD
stxrlpemJybexGScUQIXZQ+KVKSoF/DHjB83TCEQ+Efecd1GRqwB9gHD2MYpMTl9
lPagu8zja6q2pH77Pmx7eu1C7saXR36dCudT4r2YtJ1JDGof5eU/WxWSfZhKdosZ
l4Y2L2ke2vMx9BLPG0pdY3cDx5AXE/XRbV23j2xT7wkJIRNqvYNSStAh4iHqJsmk
3Um9a3e9xxYM5Z+/xPrRIWSF7ZkX9NcX01TtcgmkmBiZvuiSq7G8bV99uay6NyEL
dba076zLL8kd2eNSAR5Dtg9bgZhwLtHL8EStzSKcK1tqNAsRl4OfvjKSh7vjvAvn
NG/wkCtbfQtfkslD8jnTbz7VygDz9fCrWr25s/pOeJ5rQMfoJuzoyzbLZoE2Ied4
bTt9mOzSE9lesRwDweYwf17AacQkrZ/fIYikJUNTRjXiaRrqHK/E3J22rLjprLR4
EAh6wWWfaDVQqeGe7i3DxOIBFZ7LVke0vVn+Gf53aW0hnbRShEDqI5cCwRSQxMXi
ch63VkhC5YcErk16fYY78UiUr5vex+GCOYRDvuNA53g5vtAoPehY2u8eSjPzxxGf
9ci1q/JchbfoOcXefiW5DoA1YTIbI5tcxba3cIal5lEz+LC/kaIH735UgrkRdq47
wjMVenJrUC3bs/PLOK/O3sJMHYPUK5Fwl2d9FHm8Gh2m098LVBplXi2+IjBs1yDR
eQcES1cJogtPmbLm3YIE1qpjAkulBKLzlu57Ec7Y86pmPOfCZkytjwNOOAybt910
aT9NsvD3nP0mDe4nR6Wb2FKzzra6Yk3Go05VTmTFJ/RpAmXYgpaX59A4ZMtnALdA
1334TRPEC1FBA8dKSLSDJBHWzDjcRYnpu2ZIqLzdiDGR96pUr0ArgUwpTdTY27zk
iKBNwwnXusJM4ZagJ475q8/h6OLo9onM2XRYGsB3z31r5j0SPqCNBu60cTKfQJUY
xUJuDj4gNBJSxaAyeFXc40QcILhF6/btWyQ6YLpdw9uzfL87L3UAi1oXWaSeFX6f
1bN5BtEs6v12OauacdvEgUxhBFn7JdO5bKVJEVXdmL7nJ53KNTz2ChBhBRkdoSZx
uXpzUAViPWkQE1AgsuJiIaISmi3kWGjNSdjW2sJkEKmxeuKX7asQeyXC+6kfyk6T
gknRuHZadBnq+RzH8/kNbFjIgo0xm103NigDTIn5Df22VIcgQ1AnxrrPOrRpsuZb
Ixbg998FiqHDh56EXJa/GtEvqmhCGADpyEu8waaqflBDTVC33s1A2ag3wB5eZdNk
VA+PmlJgYDEGTB5HYuT20TiqotFSwPxvR5gXxwVlKHsQot4Ayl6rAoErW049e6Yd
5xmaUFdCORBt9Y55q3FQR7fw8gQon3LkOeY+WDJop6AEfmUqp/oSe50ayR5onKk2
gS50twbFQzYe0Hk+Lj3C/dqboU3Hp7tOVrVQ1IJUhn0e6KQFcR69cdnpJejDxhEC
/+/yF5rN61FCNM1ufa4lI6hLziyqQa2KfFBRWmOyqyhC6Oe1sDJBY+74RVuiY7WP
ihR32uMpJmOE5xmXycacNDUrsOnRZ8MuRxCgv8ptOkIWbGv0AxD+bnpZdSbw5ufx
BMZvWDEB4fMRPZ7xsDAQPB55AW3x1WNKKm1ES03zZkPQSqwVdN2/3TsBJ++O3Z8W
A0C+CaHobDrp+WqcF242qNZ9MBQNiYZqjfBGc/931aqRo333x4P99/rsxm6ygowy
EXwxjXrktOESlbLak9Vb3W0+P/UmxLJnlJQDYIaqgx3R+w3Z6OxurQbfnBU7F24U
6d4n3MiiucgpG+fn++8gPbSt3yqAn2qar2ZGOUwFv3IToB23Y+zb4rrmv1PTKWkr
ETNa4DYY8G45s3cjwPbVWdBfGG/J970uKw8lwFoZzLCElqDsMBKb2dm3/vD77CGN
xTHx2fOh89ifJ/a7vZXpeT09UHXECvP3txsFwGtW6dwe3y5HRxxw2wd9iVkRx0Uk
WntREvnx+Zr0bu4V9wOyzXSOXsRoHdOTMTfFopcLth3SEa+aKgYuPs2/6zDevoU4
gvF2Kn120MjRkVueX1IT8z5N9tnn3vYa4c0NNzcuuyiu8UbhgUcYj6dr2Uix+cJm
Y2PH1azk7VbOoFIklJTQ0Rb6xMUXS17vccgsddUf9IIRQ7WHS4/I6tGFO3sv0YB1
mT2Fh5dWHPsErabzBH7o9fiHsa5Zfn/pqnYyPXvLBJmk4xdkFc2v8zPq5yAwfUgc
E7uOi7CxRvONTSryUioLqN9fQ4izf+YKqZD4xUQGQ6iocnSzvZIf00Rd09DckJr0
+MXpzMGlYaXAOhT5r/tHIXunx7B4re75m/Eqnxle7iX0X9Cf2drjSqZeSH/uwBNB
Vy0AQ3UBNtLRUwgVDPD1gR6HtApjssh29qRjsIZtgRZs+oa1w91gSl67DbXC3AOc
Tfsr8xzEvIbmarO6g8Zve/LmH86h+7T9gmMngjKP9TAiYNC6rJ+AQ1rBBa6OP23M
EYkJ7G7D9czYJB4j9oYPPUsv7TUZrS0BUiUoT0m7m5i4hmyDYx0ftni+3vTquCcs
oPePvSGT2SfTtZ4spg/AwbtE27K0rUyI8eDM0n7kF6MIMo60LY33mbJTZBigXfoh
v5pWjYKK3yUNNIvzj83QQLy2vGkStoJyRo+NSmQKPnc2m9lgbZ8KIoCYkM9xxLJV
HsX1cG4lVuBTAkAzhWHikKvWDk2tvSUnwGY0j3p4husJcjXFShVHEg9gv/+ZTl4I
9ese1YT1CDNRtbru/8rXwD7EKfIicJckNC+xVRWHHyoB6cE6/5BUOyCJ+tXeL3KR
/XDu929R0t5E/hMAL01I96vN/kDWaxsB/9AmIyVvpf9K5YjOB80dUBceMuCm2pra
JqT28aXaS3gV86eRR5LF73DDENkYKWbUsNFiAkjAJYszn8Bg8by3mhgpiBE3/p8r
MPPDd9wVMZQ/VFyZi1C0fC/jRyBm25nKX1UHUisDvTj03QClLxRkeoBrjbj79qFV
ioAN+m1AYx2SwcBhJpXpt651fSrWkgXu8raWiUof1mdY9bbikzaNUX81NLCDML7Z
6xeV4Vuem0zFEOaczoM5MjogKr20ncM/Rj+7sOMVJjT297yrTsSpBm1sbpTzUX8t
lxcAbg2qhW/AYemWa7l8Mx3olSs2ViEHtyhjWlBREhablhZjDJQF/YTh78eAI/Y2
Kpq+nKfw+KHcH5WA3OfM2ONs4M+I3VxDbo0pGgUHe6l8ET8koGaOzKF0CNbKXHli
Pn/jFP1jhM+g97q58AlCHjP5SWyflkMICQ+rr+p+JXqmeMt9JApSC9ReekrXR8O8
FcMTvb8Lnet1tbyM8OJ0N2NZxpbU+8R1FKxkkTHjjkjSfnQZDT2mwUZZgWixG9Lz
BL6tlFFqRWKO18EqkvBU+7OCsUabwvxoL2V2L/zmwsX+nbq53LMCgsFWt1wVPA02
WQKvgb6xwgl83Dh642zo+HWpuEe9WS3n1pkoPe+KP37Psorhxh/tAILJvQmbKFl5
ROXe1KxXA1sJehudWtCnQUjzqNqNI5/ZfdUkEGJnXyhH8NnvIrxQXcJYWjQXzYKY
r4PeIz4K++6UMwvAdZcRcUNoyd+h6fesgY5ItRh8lCsQyqnO5oltzAstF+WXkzo0
AkArDpBEQQ9YifZiWeSAE8gPbCWaSLAyiAvFj+t0oPW7YvUxTe6c0G7q/29I4PRY
nGFw6ZQKl2R/WAAuTDkzJaOdkqBjHX0r56hzQSY/Msh/XeLNv1jLblQh3yiM2VoL
VHz3DTqH7+o+u/uAMitH/5bE7iwsUoJrwIjuMF4z9XF0SCioEACAa46VKMCe5KDw
7reIbyA2ueDECRoYjdgPqBfz5w9mqbdycRlg7UPcfxuUhA2k52TkGc1ZTTRlw1+c
rrKe/eZ46He9cN7sPFnZO4LHxtrlfbGpSfpkcKz0ny1+3r8YLNyuzf5VSRUWobfp
X/KGWf1YdHdEhfn/09/GO4/pGbBt6UNe61yx3ywbnhrUM4lLok9N/sp4h/w5O/4h
aYbpN4WQydIBBO9gYWbUzF6tNGDfenEn8sKXt48BoZwyMBDBNm+NiUgVO9PDa2k5
Zf8O1orMjnNJJzazX8aSPvtaYIrygmEzD2Tw6yXEqKkZBQ2ImeSGbxywxhdMHo2g
O3e3Pq0NhCPt2YlfThBCTDg63ylfNL2at7Zhlv6u6eFn2pDiXk0KyR+u+5Qjv+bh
PYHHnjECt7pYG3fwYWD2rb/Er0/lTnlmH9sEIDpHK8o/iA2K7rJ1qQKz9yHIW145
V5aS1SQYbgjEiMpv1a8+hsn+Z8lPOo7+8+IXIKE0DJ7AHppzt+6cGfNtQZXfVV4S
ed/CuNH5NO8Tam5/GrGFBazNTl8pBaY8AUXJwXRla1GkiTpS3BnLDxwICviOQSO0
gx5bMYG0ihveafWRxy9IcaVItt5cXERbgTiwsyvDyUrP5axu53NMOe06XigNlmPG
GXyiU/qdcogV4zT/dY2ZjgL0IbEI6zfeXJ5GZmWjDipr2Rl32OVuqcrV0Et+6Sf4
OtOfg0d4DQ2Yn/7rB72tGRDs6uDgmvIWQWYvJeV/I2eOHQbinX1NysVF+fb+5GEr
T8rYN0W44rrv0lv3oBEMF8GnFH4kZLEQoXVZECYKQmhu8LtHZV6zVj0u4YY+Bpr+
aFldCV7rKqJj32sjn7tMcNYb9WXA7nKst6QCgZYqXAvjd0RFv0mqzcWYtDdSAo9E
+6Y/TXILvTBU4xzFC3d4qJJxxUpC7GuUndeFYRND8nWKu1InrDDw1zzjM0Z7bFVw
MavzXawCAnSWx8Fzlcd3HbrfhmS0rSJiLgylBaI8XDr3OvdBTPLVz5fSJVzDhwCF
jXYI+t2M+6f50WMCXfPUpIuFOLGXToWxLaTMVXwaH5NW3MCJim+G/56S9fyx/GKN
YTX0MI3bzk0ZVGGlphYONRzpCmicsKQccrXCiwn8mjf2jnztArhYd7WvJk9WpuNm
u8SJMjpkdbTPUmW9rzvZDv2hz7JaDapOBlb6Nc8qHUpTdYAZ2beTD543YlRAgEyf
nQfono8MgetXxXTktd1RVXgMvzXNrIyVmTntPE1HcsAnZPRPT9rltDYZa6lDnPh9
0zr3Fk1Fcv0oz1ZXOTy3zj61WC3dLCnMTT2J7UbvPVANVcQqszfgM5OO+6TYU+1r
Oat2SchpXVgaaO+l+HVP2YrC7J9tFdOip9/hku6Aivrkj1DA4VHlujISGQZ9mso3
JQoWk8Tau39p1liUTbMKJzRkAXOVZrclUFtfPnOtQBzzxo2OcFkAxX9ejyY+7q7i
IQWTmPD/2wSyFpCKuUqSc4m0TIxhtVaVCaFGgtzMFUWd0qnKZKKNH+qksrjkPEI6
SxHul/3TMdpv6p/AS3XsCh9uRxSjoKOif3+blXSEDO52q6zks/gVOEdiA6FIXj/p
GGez6asIf+76lYJ/5d+ggWSAJu0pUmfCB58PsYLBsdnXJi6HuviHiKJ9XN64vd9J
qG0LbA/P6h9RZMlLVJXoYEdj7MNORak+1JXBV6MQ8663XIicQ2HNbPX8NriDb/R5
18do+iuc56kgWG4j6rgnMyA26u7iv562XZCK9HzyNOsXxIIz7qEbF/j6wltJwZsU
psfdThgCw9DGaqqEMk2eeDxaQUVdrQmPey5S2JVLPSTxUuAtqQAx/Fj8DWJ1NTOf
lKWaBT+3759I4KrwVNFHD5VtJH2ISubRbzMMDL4nqNDo70P9vPa0usshgSDcuExE
QgyusrZ0z+72tNfVMfKa6xyR0ji1WB1awOQfDLqJ7u22ydBG2WaESuaT7SxZQaAY
gUGrzASss9P5mxwiTTjF6Q9DJqnB+lS4WIcr8I7+lGUT8U7y57QUa/4y5gSjUw2z
+dc0FfVTHce0BtrHgl8mQyke8Oxd09Ja6Qltimx4rH9xy31Iph5zMTXGcZkM13Nf
Z8TaR4GHUtL803MeUK7s3QjCi4bSZOSC5iSBGE3YI10Z+wPlvfGE8IuOd/p+yj6A
R9lYQMotLkL4BvupdxtQUFoIlv4Pl9rp8DMO6LyuoOGxnxftB0/9ueO/ovO+Jh1U
htDNlhpZgHeMqv41ABPka688hE3YjP8dIQpFuY7gjg436rYOw86RoCJVS+rADIR4
s9uU8RxOfch7M8bQpPECTBa8eBIk57NocPiYmEB1o77e5KZpMb2jd0gcGV4bK2I8
ujhq9KNzlO+S7P+2ZUKnSX7325/cM0Hq4Jgb6scdIRxSaIOJrTWgyeww+2at/i9V
9vPeVWaGGHSLEFsh/HK7ZMJVI795bdZrKLdaJaFZ14S+QI6FUp+R4+kCvuWQDmlU
wooAQdt9ExLTdOdiACsnBjDgu++yUhRakUaY1zxKm4Gflvv4RQwkne+KcwYl+5tV
2tuUWTF/dV9Qugatt1H2GSeVYU+B7FTKcgoo/rbx527paxPdL3gHXImms0pDSSF/
sToT6ZjjHko43/fq+ueMzpkcw1s2tw0mCQJLnp4+pw5sGdgJ2qtUJFqYc5KPwsUG
Dur32ILFUa7LKxkhFS0TTQ99H7TG8PUEYiEV9Y76RahH/iAif8U8t6jyq8eWlBHI
ppP4w5KHs3mNnu2gY7b7fC11XtqRKeRbnsdlzBLEXfgacDCFRJXv02PRo3myO5Ao
F0Vznd2ai5PgifcBKF1pmYdTh3/IbJ1/RjjFAJPTIVUJ7ihBMTX2WC+Ppq3PmeMx
T+1c04SoPG27oUeAGDQOzEEgGRyRCVhmrRhCoQaMgrduB6BvMhqatR87pvJs3SBB
JmTnK9YqufMizXcCkBDCP3gxJMurkZzoBGsI3fYXRvyvGz0sayaWDdR2DPmkxdXO
ofC6sfpcKCGFg88t9hKXUHLqu0lNBnBCaaoMAzkIEZrwPexqD0D6J6UYnR/1Dgi+
sLcm8oWUjMoKcoSPVJ1YlCqiW6Kczp+4pgIQrjOR86jV2LmlhgZvSDUO5WmlB7VL
ccAhTZkuj0zWksG0gEEwguux6rwH50pnnqO/bBom/e/7E/yOwoZowbiFbL1Lhr18
ZKSyy27K090tEnauDw7ZRPkVsn5EY4M7uTQMueKfy9fPIgqE8445L+3uSf9RH201
1hXBGcyvlqiICUht1I/iU7QEIRXcZ+gpmJPvYKEXS+F1WjfXAigDQHKDkW130xZY
+HnTGMqijd5oE1L6VvXXyCMj9OclWxB5NYQ4lK2hee+A5fM2bZqaThCNpURkXehu
i0/rVzyMPc5mxvNTHxRwRVE0KykAzPgJF+Wx9TeaEbyhi5gGi9Ky8f9h1/HQ/Gz1
D6bGh6duekoKAuqHOmZ8KR9Pv8HIDROnaLH6G/0+dzfrlcyFkX2OwjEqBAPrWytj
BaV/rzu4qFxaGqGDRR+f/et6XqyfIrXZ7J1eAcpboIl0BmGWGAXFrXOjUjmhurRt
IAZKipccY1dvwaCYU9iAzaNAhUslKT3kpc2xpwqzokZl9K7jC3dI9k8kWSNbPwwy
tIigkXkPyTmQeqNJ9DJvS4qrJkxKBTRKvA7jXKH9bXENg969OZUafPsOaHTHBLrc
wEAvPZnkZsO1xrwJ0XYvRq5rA3BJzBY7D8q5UNRBNztcyOG7EpyshePt3hkZQxk1
TyAY8NT0xbzidvuAjc1eBKO6Epk3uEqBtziB6hBHkbPPPh5O3Ko38iigd07zVhaX
mEh2taHRrKGj+mO0ejyGPzou3Lunsctov0QH2rnllysyZlvDs++R07H+b5GigyIM
ow5DM6wBIvlPnC/SRBxYbUqM4lQ2qfVSO4IZjvUAQAB3RVf83dN7l0Itd2/Eaib+
lQ8Q3kasvmaX4nNgCjo3gtLd31DlqmQ/bngII0hETrzH9fXc299XLhwQFTejwMZH
Q06m4/4W/F/W4o6CJOXAPsch9FMG1zCRkUuD0fzrvE/Pbj77m+u1mKtpKH8J9mO4
sEMgemyHxb6B+2V6SBAd+QZqpMFIM+zUx1hh9Jmx6iWbc8IYVRfEhiGPhHfQYKSm
vo+i3Zjhz1Eha96swod4YFxRvtwzNqknr5UAFvJu7UdYEH9yyePQrqRENoqMQAWt
clLc4OybmH473nA9T05JEKM/cxzZUbjUGVkoifwNFkJa+sldwIswEIFk3TWybrVh
0pnjSbOpw2YfHSWM1/MyR+NC6Bh3v0l00hg8DgrRTGEQ90/IEfiVdFUiArd9BISl
NiLB9lI5o57f3JogUwve/2yv9r0rSy7Ix9pDnF5QOlSHGcwJYngP+2563uclF0jb
aLU06zYs3xNUrDbMitcfeEfDkCG2Otj+uWtSSbGzLu5l18m4hrV5pFkRcqexSUGt
NGMbJKgjEOu5YD6PR5z/pvG2zCmZ6LXeIUhj7r8RAhfi7gBNoOF6B8TlPy4Kmqm5
JX9fJ8XImYi0y+BY3nvA2w8G4NUHlVayQjUvBqvo2nUOxFDzB7BYXf1krmTrZ78z
qkR9gYLiYxyX9DtuoEFud6jRWPV9MTqM51pOmI/8ruJnmXJZXo5u1biYsGq+DBG7
PsRF4SvIwgr3Iz/dx19r46c1z9FzadlxAHp5IlKJ6BP7KkF6cU3BC8IXdxjcuOQx
WeYorecIFdIYFdKKJJT7Iwu7IW762i6XQCZWloggTg9uLpMdW1K5JV3PEyfFp4Qk
8lsigtsK7804pp6MeBl7kdJfCClMR20TBzLym0r3CiPsHuPIMI4iubqQpxr0Peg7
ToVqTvjLx+4o92byL3r4b0oPe/Rl87ZDYvLsHJNpz1eXH9ipe6Y6SSLHKZvTxzIX
eqOUx8CvO/K9n1q5vaIFps3ELbKIvpcqXO4KeU9teiMdhBbPSp+xC4ARcqLIx3PK
T6/AQmZgP+BQKzBiQ1bdDbWeII3mIDOjFEvvqrrRvqJ+a9yCweIowIZ+bjQHYqYj
Hhtp5RdDx7EHkqcpQz4XISZmGspv8Xs9jFxcbPxkUVdMH07fXKguM90A8pDLRehD
XCgqU2mWXsUSf1v/9lPkkiAyxYINnSoKj8NKjB1fg7F0dnGMmkgF6rINi2SXHhKX
S+np5zd+VbTCQV+jFH+52kcyHIYRCFJUXOy3dK70uCPHr5yvt+5cH1VEYAvdwEsg
Y0zGmqoBngxQzjpPTNjT22732WvnecSlIdDLhSYaoVojmGoToWtFHenouvaCTmRa
o+yt8XBEZha+/t2Gm5OlE0D8+ZskTg/7eewtIw5iaqCVM/oevsuQJ8GkJ4eVs9s3
2IQo1ex/K/lP21d/VTtppBfYJA7PyaiS0P4bTuVqfwQhfju5Uc4HSxivWWtjtP2+
2LAEsZnzLXWOXfL7QHw5UxTpHyMw8Z011Ni9Y69eh4i1CrBAYD93HHd+wRlQPVkp
33Xd1iZfcdOK316CNUDJUyA/bzLFy5PwtRubf4/95nE5yP9S4yWd/sbshl0QEwJd
OyZuDhPw6xxBhFUypNhbXM1voURWhOI0MQvEflkxBv3c4NlulHaYo93po3HqF/Sz
Vn3WyfyUTO5NEi/x9xgewaJShIdmHscZuS6/08LlLqu/DOU3Iac8ZCFXc15+olzq
MVTW/yaH5FGCVHD+mMA5eb6Htmh/oOGQjUZg4Ba2uyUGQzVXFlCY5hLvTnW8kd1D
AbRx11OmkWg9Umu4mw/8eKGMVRPP26gY+xVcrRQTXPvAiuRUFpFry79wKZ8z03i6
4PJ510F1cZAEtDn/F60DvrX8H8qgDZpc6WgQe/v8zU1Zth4Givd49ZvobcE0nEk+
xP2dFmFdpQDe18X1AQimcYcg1nplY2qLQPmfZ0mxPsPFvzReu5fKhW9rEmdG2MBC
LymgQh1G2hrfn3nUmAORRYBoPFVQDqHlGlja28aXT+xC/Fbn2iPYu8URl9HGQvtd
FLKWhgmSeenFKIVVTklZNemJ/E0tCRIbdv+SV3PsP1V7pmaok6w95jq0plYV41te
Ani6AM5KXVBFDkouxL8scxrlROkWHo5Y5ecvTu1Hb+/WFwwKkyDAo4KxslLyBeNz
vLyd9gJhb6LnRu5tegjZUCuZq69JufobimF4yHPR+6sMFqhu0AIh5pzBCnm95KfX
yOUe3s23TJVeIzPo1smscWEUxvC8j3UAKhhSGgz8WUyHwnfgqBxOW5XeAS2m1O68
SDgiFgAWpWmUJw6iZ4QSvnvX+EOk1boW1XZ1na7j5VF8ByvLf3zEzgJnPQS2eWV+
xXUmEmd9Gd+Bw/hlYB4SbLrSlpDeLJz4+1bTS0SkHkT4EFPJNZsNWEzxxEkNZZLZ
Q7qof7toyTik9kR7Oivwjp0q8r1leRo8PPnpqivc21UfSVkv9Jz2DkCpmXknNk9t
juENBR1PdjE9kWNqavlhmCAoMMUITV7cELNKm2+dXM/ZMO6h3iGmmAbo3squI9JA
JHmCovMnF/OFz+dkY8G9+lnW8ipWCOnAC1TjBYIlsPgl3D2XLupufkNnAU4ntvBH
iyqrmjHldPO/3SoRpRNicadWqWMY7qvw8XwMVGZiOzFCwpfKPKHloRxSNgas5SAu
Cs5rrxaTMhXe0KGPs+IQ8Ze3viglEqhH+Bjh2d0k5W4qV2/EqmLG0orHxT/Ejal3
8OXvGbHR6itOmLjccMe9OB7/8j9df1BRk5F2lM2HJXWYwywSTXC5fWnDcMZ8TrJo
TZc+i4Rmx0yWzRadKVknlYdy8X0AZXTItmhk7Iq0yomMaTlWJRktaTmHIJA+Ukvh
mnDzKWJW7aytHr36uPr/n0iQJMsw9HjvwwP4tpGH8I4MfIiKqEw9q9jNvvOntEYh
NpakPmAN8MQ+DSvG/2CWzPNWyuQtQojn2Z/ZJ8wuXftPv7Us0EQSYebjMgyu+LAc
r4+hXQxNdy5/N+kpxwkmsapqz1ERoHnwJeWXw7JpZeazMqnunqqEF/5EWVT0cs0U
uNIblxPHvM/u/d0kyprutUhK+LETXC+w5HS2ItI14qVDaMIpKj/BP7/KancRVVc/
QqxZWgHJmbve++W9fhsyQUyAYJjUwyUcVsixjCV5MOP0G273uEukox+pWKwooYmk
gAadXgxY8ZOoyt6ks2r5NzyvkchRPLx/mtU99PZYjoO/k/pkKsRKOUbtMnB8lOgW
wvbLObiOqWk6r5SVl4xAIRMjkpXjqwu5KBf9IB1GbhJ2PzzK0ooxnBQl7/wKH4AA
UQem/9VyFSupeiQ9N4xY5suJPLN6Gk5z2IAH66vqNB7B6QvB+8EoUEVxuIlb1vPM
VnQU4c3G8Zz8lNAKibtqmSqIDv/4Y08lZlkQ+at4ok1NLrVT3GChpLZeXGUfsDjO
iBo3NKPyr1V0pRChWbfnYVRzbd/3UBLrSBaUa53uQ159OvvzDsmVfCjIvoc9epuD
x/933Rtz4qZcdrFfPX1JZ936QVHIVKI7/yRCGAbRsi2aI3oV8ldEqcVcywyOTcos
LVnactkgjehK4f9w2I094+TqrtWBvH60QvNtluWuwXfICgAktCoSu4U4XDcGYIrL
C/jQoe8xlTvcOM06PBAXn+vd08yWd06WTLhKjm0dFI4EZgsOcoHDaCZW4NaZdH2K
WFfJ/OBJXKtG1FEtj3ks21EK5raAgNyj21Ep/LX7cbQ/588zVXPhb+wHjzOtuYM9
06geB49Y+NmdgdWolzFYjvLBkqXsRQVocZ55foC3djWmmc+aeaxSGbHbVaNTJc/i
0T0NKle880MsWR2Th++YCjYNjpodaXCKVmEuFYQvY1dLUAIyv6r9PfEJ3rtI7ZY4
ZbMcHMgXK9j6ID+r9vwSCXHyn1isLzV11WrT+Bnb7HShgrhrBCegDqUJwsjuT65M
Nd5CSLl1wcAJlLO4k9RLgcSTSA/nuQ8k+H0ok8s/ioQ+bBsaB/YDnQouICGAo/Ng
lPd+1BqZDBnwZsLwP60Ta/FJoEiKg5uTHKmdS8ALHWD1Ilt4ROnqRESdSQSZPCJw
H1P/gETgsGZ0ob3eRrEl+wbWsShToiS/BqdCy8UKLV6Q2t559L1RefzlN3yOcdjO
UKFAS0pbT1sZmMCX7qF+7XgpVviVXzsBbRbV5gEgmvk0FoYPsTXjg3mlB6pmqA96
+sWq7Nk1KxF5kTeQ7b7ReBRuDEPZL5Flp5jIEyKq3rhzpSu7Hn2X35Iz8FpQiE7B
qL2dDVTvJu9/2NIlQl4lRxvZg7Cg2qTkC7xUynSclVZHgqXvPptfPm5lHwFYnun6
IXyHrUgpTX8ZngTic5wgFzqPIF1jpjURgcz6rRJFNrtfjNEvF4bQnefwsIpmNDYc
tk1Hx5FONerH3i7GCQn2c+LsW5BCFT+y+0kqTMmYeewUhWKyecqXIArD5J3yHPwW
TdaFNamPADMgbFW2okPCMavul8bq+xx2HZhXGVnq8Nk4Nv3Z2o/EsFh9ZUEr/NfK
2uJ05DFkExinAcN7GrKIlNqmwlNqeJRXO1orJh3nDv5hKA3Kl5bzQU983F+sosfv
nTgX+Tv9W56HeQlepnI0vjRcLzbyRU6U7zVAcymmzxzh2+Zw6pVXeZT5E3Aj0Y6J
CDiCzfjREvlElezMz+EOR3pb8kZXGU1ZaRERY++ACG047mTXDC+7s7SpJin3kqni
CetZmtXk+bY/eaedKgcKCMu+dFZkFTmFBxr7mA+8gDwQWPuWNTwB/hEH0gU0+3xb
F0jwFtpdOhOGCD3Y4thAUXoqPd8exLLaYPHn3qHO5CNk05NDxT8yitJuzb3edw9K
RocqhAEqckaHIGKoWRTJIDvFX6/r341IXctFUvkR84+jRONcNOkzFa3xF//6v5aj
/ICJWboa7UZj/+vGpL3ZA4UNx6ChSHT+EVH62tKs46mFvFyECTlZvtkM6a3Km2Bf
pokbCsHPjpoyEL5t9PcKCVomflsY9owyGhifw4PXQ8WvyIeyVi+FoP52qr9XE9DH
iTkqPmn2KG+gEfrJ0A9SdwKOvM0+PteQkU9L3YWxj2YamU901JV3MxiAa5uOfhtq
22cb4C52ashbDHw9rzJAFyZL6JHpVRxVOydgJG1HTcfHv6croWdFP7OQCqftibdh
DxzQtjOfUXLdsOgguWdtpCFiu6hazFvuhfC4g+jaeucPDlFphsECPw1iZcpV3/Lb
HrVrT8uv0jHWpIC+tVbL4LdNaw8VmLfq3HXnJpB096B5wOLbQ4wMxxtNm4rXJDND
Ccu6yNac4q5WfCWqYwVGzI0VumYmgJx6DXmtCG4TWSPqmCa2YMNg7oJtsFGnsmkS
p6HyOW+MPN9Z/9vwjK1v9WhLZ4LaGGD675kXWFw3lCHjNBVf6wJtVDr2XLjpBAjM
o32G8JGMJTlI/NzqV074vIohuq2pMGVe0/b1mGzvs5W5p3uesn1zzayLzdPYgljx
ppod+Q+5aFBeTpW+hvGbSrfV3BgyMQufyZ6b9nOHcCtdOK/gKDgzmavkNPj54OTz
3PVawC+GvD1e5xNgLqGp+HIcS7kgrn4eIPAPpv8NjZt5ey6QOuBg9ZCMmjvqPOxw
1bmSyA2BDzlzIC7LooIclGXlLFadSq+l0haiEX2vUG96X+onLFmbQSZ0bjP/k/UZ
jnJtnarPQlAWL+WelGVWO8PGunYXNj534RuriXm8lYjeUjg5kTDGhFwIZHRounBE
iQua4ISCX3OjktRNZxQnx6aBx9agInuQ+Nk8d6pcptqAE+8PGLJuPunD5u7bcsEl
iKALpvYQzRuwD7L6Ud6yzfxEfvym7TDFzpoPUCybjIBp1eOfNzxshD+9C+wkbl7U
O69UTbhtR2Fv+F6+Xk7bm4cfBbzjPWjXppOXoS6FflmjbWMQTdfvE2hR/ciy6abu
tgkwrYFT9jv1ccRr2MLbnSUsK99w3YaIRTBhwZL1S+P41ZH+xXZlKJyHCWhQRBNB
Zcr4lezW7sxMSUBE1v2KPSrj7TacaFCSn8r6ob1lbUEdc5GdIZf6SSmy0kAuoB7H
0WomJHZkHSwpYN4MEzVFXKz8BjctB9hyd7lPYwVBXasurA6ySOgi3hArFIK32Vuu
n/pP7naMfPIm3gpo7IehIV/vZQg6A66QCQ0WUqc4ZQPS6nm2KW4vvnf9aljHKm8M
JX4ma5M0ekLVdLZijhh4SWA6LYadpAHy8aj4RqDsRVGJM0Zv4aM8KL7b7naT+Zs/
LsiaXPeEZmIDlEfcdAt3QjlmVrh6mHHM7+32+7+2mkUTDob6PS01zSLfEMNAk2B1
+ySuRSwH1JkSKirCO7UBjeYNldRw4IilnqcFay+wrW5ErpXhDpL/SHRz2uWHsOKL
gF+OJdAfh8oOFje0uUryHn8qMCKPkqvopKyFGBi+bvJ8x/eDjq5GVBI4Jw9BgAxv
E3OGZTkgFc6r5vqA+CT62GGdqVW50R4AP/XUeNr5zHfEh8PWo+c3MftQAAw1IvEK
NPrdl7Zv5EEjrkzslb/rk3hrgJgBtmCc98tqLkT4czxJVqHbLec4HPkZpw/OEqv0
3p5gLuO/AM8d8Y4ixaiWBdQbbozsS1MMG/vaV1dSUm++5LLQffOHgSUN6wVnRi6d
OPFqtGUN8uUnypxCGGuGfzs1gHzD1TeEScscB1o/h0ojvb/7ERilHvjQSA3Z6WtT
0+k3yquXLjL52uWnPg8amVpW6ywbtO9On9q1oYK8UoSYQGVbctuIp0AK6mNYrH18
5aKiSZNviAsNhRlI3l9OJjHNBRAljpwCe8fYesKYe7GXjShZpqX0hFBDbH4tIe3m
JrPe807VnNQA5hqwo4cH8AKG5HQph95dEPTcM0grjiiJA9UpEX92agDAdFI1oh9v
jcTYeS3j1Lsks4ASYUelwGq2g94GWxS5gtZd2+REpvMCimqYWZHVWJn0mRSFKZyv
N3/HS+weB+Jcap6mdro8MPmTjHQRBwQB6+7VMq45LAoRygyekTx9PsWNfRFdKCx9
rjKnlc9w+ZAIBa17dsvubc5wm2otaeXs/pXH0V/MrSHYW+MM7/H91BlZxNtNFQAi
I72vsvxwnXgwKR0EHWnzSfYvYTIzdrmPGrm9aO0mml59GjYvz2+TnWO17o1lOmi8
5f3PMo6DeJh0ERM2IrpgeFASIOAZHklYYNR9LGeKxtjXfUkGCbChT88yy3ToVEPg
h2lQSsh/IvRwcsNBC32yxFinGWfp2gXX6tzGkCbWSZPfxBP8HAKq5uTf2NQzG4pt
VmhfXCS9m4QjWdrHLIGwE7lKnAfpg5G8zALaF5Uiyx8Py3G5Q/bg8Sn5OtFFbVlQ
7zT0T9/5vaoP25C9rj4JV9y8UctYAPioQUoZ8Z9g9Be1Vpxw8iL0QQP0+TA1jiuq
p1qkizbQV98InyOkpIsgfYXjMEXr4P/PJya7GId+s6a9s990Upoe6FOkr0JcHmrO
jYauwDH11OsyCamIsUSIFQwpHaKvEUs3nbX7kopxv4/CRrmjnupz/zn/HC7P/wuG
L5tshmK8pxbIAq2fcLqqrsgpYGXDeKdW7XdPu7+e899P5ZpOjtGVAE8wPy/b+L3/
htC2GW7yiOhn9MGIBA/hUCrjvaxIzm3Xxt6PCZG7tACrAiqudx7OwhoazRaOWruH
xqFp2t6tIMjEIi8SO6BVP5wGArr+WCp66EA465oi4Ig5BeosbUFfZyfbp5Seue14
TgJIDGMdTcOLUYQTY+IvZ/GarmH+lLTRkUBmwhuhtRCHHz0g8mN4zOEOO0KM+JmG
EloEOE56BpeSuadMb9/PXA9AnajNA6Az9F+zMJx7kVr/DxV1MH3kvC4iNgFwZyuY
4Q0ttu4/cKzjs/SPfZSrFpi7qDcBhpzfWSEDIS49Q0imWN1WflBZEpYIPVyhqtkQ
+AWRo0I3u3sRy4wE8xCeUmogbju9fVaC31RajPsOBI1kjAczkRiQfq4Tq5GkIdEJ
BABH7eCes0RN48s09ZVsTtC13gL2yqDWKyaD8MaCFvwATyGRdFQWUZWS5xpvGrDj
X4oAhx3+EFT9/EEx0tJkE1Bl80ehcIQJqSY2G0sJcvYqMsKgeR8E/bpZXtF9hgzL
Er1PJ7arm0lFEYiqJc7WUNugBS7Hy2P0QKJ9v8GJ872tmywacQYXLm8wsWxo9i9M
eRvOg9oPpLd2VaexVP8DHM6N40Hbx5Cjha700x5wCY98M+7LdOEVe/i9e05+aJvC
82MQEpMx657K+uesjQeI/cPnreaO1rZTi0rLc6wfbHKcj9Hkcr3g8b5aclmuLjWY
2f88oNiip1+gmXsJGIlPYm63zJpnVJaSPbgGZtPm2ZJzkxN2z74h2iGi+4j4ypWA
dMRXlThIHQXxZa7tdt5gWO6/7SQ8avYMhKGeadlI+NRxfToYtxbSfKHhLiXu2EQS
uDcZjrH2QCS/6W34Q3sSK5BIFfnLdhKb9T+BErbC3jfQx2fJpUnHJMiaw8Qv0hqM
QImiR8NMIt9NhzpzREreDkww3gi9gfFTzV6ip4uG3/PmzYV51TLJI2XNs+N+Irwa
1To//y8Fzq1XScZ4DwuavYlhSZHVFdvk4yGoYIzqXYw7dRoLQbdJwYVTtkrnGdm6
1XRsYO7znZpZxK1EhjElZV813Z4wkyRjJcXHbLUENe7t1gW8+KyN1InYBpLGAA/d
q2fOSb3u5gDORblUZ3hGq2jwnhForJDQSpJJaP4k+iOJOD5Egqqt5T5bQicou/Ay
71RBJlRzoSQDokcU+UYo6Js8S1UUIKjC03XaKZ8hd0ZXofw4t9+jxa/8OLgUuqnd
5t4P2YMqQZ8WpjcT2FCRSh/uuv57FZyBjMbrqTN0fNe8kE4QVDq2srvzgYthDK1G
SahHwEiMvaxw907VuFtyRUZZKHvqR6sYU0jStKTn3P7Be9LHywHtc/UEtrbNQnqk
QJGBbk2h9wVwNmzgESGvg5i+16apgqcCM+L4ZLZ7DDN+aazCbBfFA5hen0OBb4DF
Ru1eyTSaEmX5a4BoLVyEsVH8n1VZVBbs3DKy4nR1bjxBqNoCeuLWeNxisNZt9rkV
9tvRY3FNGE6ovaMS9bhIl51UaYgZFKkBtypGbFCmAwvf8jiS/cx4qLC/ZUXcAx0p
2HDS/HFJWWV2TR32y0/Hzi+pyDPJiIO6Fi2HBlZCcCzzDiHh8foxlzZD6xQNsv/2
vElg2qFboHuj+weMvbwvJEXdxoQHTRSTgOu81xqZJB/XEG9Ego3tpJoc3W2BehPV
xnhEvYBrASlIxlRLiLkJe4x24SQVf+lfRYVXTmv7wJl+luMqrGJRxL/7zMkS2bQX
mYnRMSwXjr0UxH4gYDDpLS5h5TUPHn6GYVOnx8nbI/A0x25xIS1Z+C1zp4n7YsEp
rDmFFrJI9tSORjZjLpA2mVGZruJuXIF+crCyZ49oQN3a+PKAi1iOORlVnmotRS98
zFeJ9AErdIdvPB0UwWWaeYBhP4ICV/uOHybvwc4LU/xKU0EpJMzBnpHtFJRfNWJf
KuFqm6o5KIkbwMgyc2NRCVj+++lzW0Y3I11HYAi4I2uUruzPuE/8sRBkpB7lhRAb
8aBwoVdyqGyQxwpQtZ3RDRXC4C5OSk6J6CYuiBcdvjfSbnXZYBiUyGtzpVDMfop9
BK7crsgp6AYuWWmB25kH4FiiLFTyIfJbbv+loze6YGTescNm/KvMraOWNml8IuR9
JczSowEU91Ny5A7BaqXwcyz/Yy3csVp906t12CRiVweT3+Ga5zSC0WArV7ZZC60A
Z2WMu9OwcM7mNn0/KfXVhzoNm9s3SmM9LkfMu1XsvFpQJYgHHdqSopk+ABc6JywQ
PivJ4yvbYelj6ZR3ohA5P5Cf78j7UsWOV0Q9WHUZuLLUFFlFtFZxk+aYG4tuv+zw
5FYBdr4Vnjn2ZP8oZlUM+4tnofsi8I4puJXl2Sl2rzL7/ZTDEUzh1yF8n7l7r84l
1R76ivZDQMh5DTWYVq9D9ph6eEMkbAbvZAxWEnn7FInGY23zbqAtdZQk52gbmmFj
JJ+phvosPE0xXY64yiLHcavKYlHTVg2nBLk0qy60fht+85I9dykaV5UWSN6xeuZ1
v8PAw3D4xO+Cge2i9QBcCC69JWhXwtZbY9B4sBTvW6kkRHEVPT6lmsWYdhdb1zlE
NJ882snlkJxV1dbF32yLtJJy5JiWiasqaf48UNEDqsYNL0tfe6xIi/JNn3qOAGLO
y+SV1QSSUIs62F9nfSZXVKnP1Fr+TAAX7yO2U1yLFL+vTgHnFLhGurd8LCsYJJ80
GsnyoMSSwb2fjscnzCw277kvAuRg1l1Af8d2ut1n3tdJuQKwOg98MWMAUlqj4PrX
frtO00HScFW6apA/QthtbBnezB2dwFjoGIn3dnM+6dnVE52u3Pk4EtipAz1wxS0M
6U9RXMXYzruT6XPMB9WzQRkgJ9zxMyKKxEqOrPNlQK5qiG5E1wnDcN0cifT3yuSa
f/O9ItMV+mayokSViq1dVXtURt90l8gbSamCwzJp5leh7BwEnV407yLE1thd8DwE
8orI3dFRGxzDP1BofwGP7SKRQdJVeOhXMTaWiIb3mT2lElrprbuqvrZmN++pqeAz
9ebFGyLpU78/84ipthI0CmCX3V5UgC1iHar7RRvO7hI7xHBQVQHAHfX07a4Xeq3p
vc8DRs89E5U71Q2j01uPsf6guyF4PSycE0ejIyJ9wrgeyXudy5TQzMgQWGUg0w9G
2GxGYgCC27Wlh/c/hfZxmL2sEIuSXuDKddnrjrvWCi09aSgyZEhDFGnzLLHMuSv5
Fbh2Ltfc+e+dhAEabQGq7btmbf39VAT0tFJXqWl5WCZP5iOBadq9ZBms9EjYJKkk
6v6KM0icqww+3zTNvkTviPm9W6VQ/px3eY+RH/TZNeKFTvtq4YquzaNtLIVeOC+k
EjlNqWHYJyNvUSp61fDrkECjWlqn5H62dYQXNNe1OmEmWSdiepillkhc5JVVzJQt
JPkdf4nRI3x1478uu0j71M7zL1dinUqVnCq+BOHVII+eL5tvLmxnNaFZIGadXF4z
31pptthOdVrPWaWo671b3SIhjXme9IdjWRK4qLD0coYXqSAsIKjiDVNHOd0kQ6KR
2rHwodDOWi/aFc1lSyYiq7pZg54tYcmduXGKSuH5UAc6jmd/YdXlUhlYMbau1xT1
881WtmeCFhphSHErD0VTaRMKJsFXSUMf4Tq8NEa3iy8wlfgq3fDlMZ27IsiUh/zu
poLIo82rvGb067sggqDhVK6kMnqzfcsQv8i6hIiQcd7er6X2xHV1qqSqv2xI7Zuf
dSa/d/mK7xMXRvTOVIn0pa+RneVTuxCqVvYModLyZgc6Jd3PQCW4N1hcg748TxMs
nk/CwsFJ/i68Pmy+D0R39oQf7zQvw4pGzZLQwonfHxWiAUFOg0yKdP+9MURvyWu9
8ZPGrzDDlQBiqW9CV2zI5Qe7f61sc3ONeAo4tpho50B5K7Rhw/Dpv5yNMN/nACg3
7T314TQRSxVLFpdu7JKlj2UX9SQI1+9vq/VhsKm7/XXt/kaoDBM7LbY0pLnvYhua
r13T8qu7z0sGDuiAoyQET6DYmBLsv+BDUxJoj9aFuyeHmSdoh1pVIN/WVZ0heWJR
oWqsigSiI7t28LClyjXF3akj6xeB4CIugP+6PB9m+fhJzrgzkokWv6HnnS1E3dQS
OEp9DKsPnobV/E/4qTmrGhn6Y8Vrs4NwXgU7abKHO2ERImb39Fu3TYidixVdVixZ
N9tBbFd5ioYXlzEXM66McyBesAFZfM79i/FgYgLDwwWns1bW4Uur1ekZ022kGYDD
wobqfmT5ujd1k/+BzKJrIxPjqKK7yio/0hClTi1hwbZJWnEVhgd/2+m2i/90cjdY
zbUPSlSmixRKEIDgOpR61eXRfwYwOPA4eMjyuWjioStLi1g6vKcX5XJYQw0sDE3N
Z0CegZxJLs616bOt5JgbVnPKKDk1AjjQWum2WUolTOWzmKDaiznAHWAfLSkwuCaF
7bvIglepxR8yNphiX0znG0UQqq4NBJBTC+omhmuiemZeR67JCUZJAmotDK/Ajsv3
C/50kq8GfeUecCY6VU/qhMlQG5nVkR6RgUKgqX3bGItfsWWxg+wF3+4ukRoWhBMU
eMzcz/HxivDblL4n0tGhbzSRBannxeOuVA3WjeKZZR519pEp2LyBY0+B7nIzpKEQ
fQ6+HinaswF63MVTKkYVTLMXxtFy68OkUQGF8N7+ZKhp6iGtamZSWW0vK4HDzvIH
DH/fX3tEtSdIGXb1JA16E5M5J8ahMxSIHZDel6ebd2JG+44/QR0PmTy6EX/DQUXu
veafn0SWI+bvqWMD48p4tfqj09hzU/l4ptC64zCDt9jIgjZmYS7GAC8FfjM15+to
zMJbAje6o2PbotDn7MFEwnJpY4FwXASh1qNtoCO1GSHKdpW1GjJ0siPqEFoeNJuB
KUKnLGL2qNRCIJ+vbYpQYDE6h9oY+jBw4+x3MK9J3Q0KEIcv0dfnUJpjXXf9XFuC
Zx5lhxbLaFd+IVNNDSThRVx/ohNQNoQp5B7lL93x7KFza2YFSM3OaM/JId684mzq
0cVWjYwOTtt+gatvYyXR9as16Hg0vzysf5JRiCBiX5Ac6/2P0tikKNfHDRUYnPBN
EGhcXWSA2ATwMONaT4zzGMR9JqYtS5o8iB2q54MBMir12mossRUHvns6OTKZ4JTf
xbjjBbcGVOyS/aS+clZsMq5mDl4AnC4S4h1QgI8YQKIe2eX/6EAKwSmtTSWOdtHB
9es7T5/VRP+bMxMYMFxqUdO35e4w07KOv9OhEhCqxc7XxR+DO9QP+qtrwAwUIRTJ
ZVQTqbUJ4R8SMvtq+zorlkjJtaHMOMo/yLTGsAoj3preN6MnJ77f/L8XjF/3T1Y1
nY7+dT12ei8zsD/+DfF9vWuI0yeYRo0YsMX05IEszjer9LVo+E7jTDYylpbeLfhq
wufnZQF77Tk+EE1UqGy1OHQs9h5x0xr7pB4CFskKJdMtJmEwtHEA4Xvkpn3G58qO
u18NnZfq2HCVSc8RmEJpkyGir6AW+ysuOQ5yAGwOJp7hOagpXyZvERALIBitFOXX
IhrKuh5OqLlvWIXYYL3sDOJVjbbk+GWbgedkC26s3wKwWGgof3/FGV6nAkUxSuWT
jomtCRVhyOVwWvpE93ll778tYGg+Le0bf6wN54eVHLEDo4MF6vsk4fmDZu+5zUD/
KQAfA04WUa+RLJVFHDabCrwaVe2Tc40H58HYXtog2iucTssLaMQibKkoWw86r9nz
ZR8fSXmVW8+toTqySDkFSEqDfYjNbExgwEl3lzcUWGkrwMnbQ/9EVfXMHtx7prMd
kGzlaO0HATtY7DlwgjmKpCGphwNQP8v2qpLhPLFpw3kz9gOHTcgzTQ45zd/ZmZNO
aulWbbAqDzT+ai/aZEzcvoPXP3A7QANPuJ42FRb2uoaCELY7F/DDT80H7dcAc5JP
TyIgc8qgXWXrvJa13ozYc+AOv2RjHJUVlCmuFoA1UDVLeB8rkuQtvA/m45HFxksM
F00TcmBHL0tlnAj9i49SM8R0xnQKg34qMsytpUFnfEcHyYWymSRyQuct6H3AWQBo
A1PG7jQt73z5trF6U6L4DyMacCITBLH27zBAPAXZh9UrMCQkanOK0yCZ0GasrF9e
0NCCKmdCeLYLxPIEQJvh+EWwv7M5UzXI/jGi62gkPdkiyqUxkOy5BcgKyVM/bOYx
xKtXshD/FZcRsptuTgHu0+RiK2xuMS3HlgPqYgPANBQEMHjPsqKsDFsWyqkR+BcX
DxDx8sQfxIk15twAUYxaZCs4h+J9gpWnNDkdJtEM4XVELpLMxLw2Pt2ZhCmwFaUP
AOhafuifaX9MPtTZ7qFHb9sIFsaepeKY7YcSrvF3f74p/PhFavQ8bruBkuAHaaMq
26cjCaByqjKNeNq2RLL3PIN0KfXNZIrbq2xUhIomao1S0w+QvWken+AQpL3PzERC
P9E1lr3xUdGhdj568wsGo8d3fpIrtPrDbzymXlEPrNdu1Z/rZ6JAwHuWxzSQWTAG
l0ipkvrOxu1tRSdpoVHwIZPHWXSU2NhcycK1ufdoZxCvXQXWA9T4jRL3zi2DJnC8
gEHMWlW6l5Wp3vJ3g74H4Be5XFZ5vtjuKkgdI9DwgWfbnkXlEh/NnjGIjPvZKywD
LDC4PaatwpctjGlah391ZbiLMCDCXZe8Yv6QqpLJ0+OV9ZAATGw4JERpk6LZC1zL
LO4RSt30bXGGnAF4JqWNxvRCwsooPtqMNOOU/X+/FjHJTdOGh/yeNFkLJCr3R5Zy
GNuCQ+TXge6us6Mf0D01HMEIGwIN7AiDIdccIVBNFfbZDkgeNbPHN2zu6paSWNHi
+tOJVvqs1n6uzAtakdXAkdaSIlKY7EBJw3DKcVjgfk/fflN74M2/r+eoLFdEcWM1
ddItBc/kVfeHoYI/50DjH2cWgTCLAfJehbB70CMlmgZ7L1zr3CRQpbzNr1RXb0AT
1XpIlM8wpUBvSdhpOlg89GcxTOlwul+C9pEUreld9TB2X3ClTtA32pq9J5qmi5Yp
c4Y9qSsif41SNC1XRgiTVO35mcD6DOkykhRgMiI4t4lZUdANwyDMSqnnNQ13C1Ff
O0rdqHZiuC8UX3htymPnzBtLKEMWJrmO+/3Cu8LfYcliISJ4lcfWDiszJD9XF6/Z
ohXwR0bIJ2rPyppkXq9Alc9GqOhS0MTe3h0rIK7Koc3NVKoGOdXpAp/Y7TJGfplk
wjLQjj4WeUnjyc36cD0sLpLZxeeiouwickW2y2Uot8LiWyHYz441/vxTjWwii4M0
BIBZsjuzw8EoXdf7z+Dul0K2XUYzuTAdmGZwRZCTwHgLDSEcWvZLoJQXkq1EoSUx
XXIbtAwUqEgZ0nTJ8RqUzTFZZeILV7ZlikoLRoXopFz1TKrF+zn4rM+GXqmhF6GI
h8qMFYk5L585skQnHkChzRth2ojK9jzFHivtnmkZKCJ7wYGkDpgpEbLH7TfudIrh
yjK0UQ7Eckncu6lBQzFGufjZQBt5cbHwAnvscQDyeBQHjk6f1qm9i/G76cuF/K1Z
PboWxB9YyMrL31J4j80JqzODymUv1ZTetBkQc1WESbg3Rly9NvTdBPp6E3kV6LLY
A7IfYgW0uq26TLWy6VTpby6kjBOkqiy+CIweVn3aKOMBJ168DvjmbgwAgnJEQW6G
DBjAX6QNpeeZ8TBHEr7xL6cy4kOSG0dABa5D9da6eHT3sq7HklZq2nOYpdC+j9ZB
e8jfLpHN7EGkcoyUCFVJUfAitW336gJleZxjy72V5wHdksLkToT/lDqsJejZrR8i
kyiO2HrpNWFL28HM9e2wqvmZeMimwK/vTlR5AxaX4i5n1GaskemIJFqalyLLJ4GR
IS4hHixGRoN+4lrOxblweVzNrCArcG34VL49pVTIWoQctnRZlh+kQHFkU7JLpLX+
1A8hnMz7KQb5Ixun4aRqvopfh/7Y6EL3t6iK8HCXAPNGAl9mhLhRJsNRZKSsqyy2
/PTZIXHnND2JUcVcw/x3Mrfm/7Etd8MfuPECHrpy1CoU8lbqhKdHf2EtHdV3ux4c
3DdRQ6GcXQAC5CdtEehxPcKMFFhea5Sb0+MIrYsbS13SxJo+ofvCtkuuZFKQx5SF
8KKWt/0vMZN/ZbNwCR9szp4Gfq93ZbBY+WeT19GLeDSAQctaS0+CUT4WrMWHKHL7
baEp67rwksrqpkuCnP2QmR0lf4KbsBUgurbCWb0Fujl9rHBjw5GY0iu90N9pr0Pr
sVfZUqbx0wF7aKUtg/gYE89K2sQcO+QUQc2+D/hQv6m577t4y1VjsekgnbK5VINS
4eYtJOJd/j2jdaC3iXG51fC/7p4S6sDoZxETSooSou2yY1p6MoQOAGTvmXhYIoca
HkYGhdLt2d9s79TD1KPZEV02F4OGqJTcSnUJRRgcYRKjaEDi+A/XXV0mZ1j89mq4
S5638XJEF1PEY1aJvoYBTpTrYL7U1+Za6Iu6uZgkE+x5OJuoHPzEEdILdvFCF2Rd
pEECqndKG0pGb9yCt61zkga4ANlVIVFl3JeXcSor48dj5KCtUWdB+tP2uO14z15z
/J7/xrj9ERf+1qCPJD0YmKTaJLI9O7pYPUHE59/qlWYaGP9sLV8UnMwOCGImNzkR
5J+QMPCc/hDZ5YHOV88M+W7fB7sHJIVuGn/E7yElHMptoe6xujVeTGtCcY0G5NS1
UkKRfgipdven2v/eLyc0WnhL6sj06ezlrdcP1OxlHk4KY1f9C6Wvv4y1nXKEx9S5
CMiyb0J2nLzFS2ljpdf1/yAvy62r9aRHI9D/8/O+WB5xVXG4O946OsMpXrxaaqRr
wyxe/JfBP7Z+oc9oouh6yJTlKjHvsHkii3J3rx4sOWmivBeir3IBvXEoVlhKBRmQ
FteDN19gt3Hoo8TqwN1fl9nO6qwh9hXAEa9FuYzUEJIcqn5hkonWIHrvjmnPCvRH
nB1Fz36Jrhxr/FiRAJpN7ah1vlOSkbNyfMGOfnjGS2N9sILTYwzFdnfIs1EBUGa9
g7jWyazIPU1P8UCaRWcFZku8Pu8GX3L1j6HLNrcFfK3Ab9SPWwO0N2FN8Oz9sq8O
xLkhHPFURcEvXVugWwiZ6cLGqB0DE32PA0vmBuoHPB/0Cmizn5nOkTC+oGuR1A26
JkOp/LITJMc09Tm4rtugWO4gg2AxWZY1OAb/hwu3zjtJRkhA/gpn2jUEw1SYtvYF
Za5YYyAipA+FNNsee+QK3MpsLlfJpj0R9WkUe7vmN8195r7ae5b0oeM6k8SKyEtD
zM1cKf+4rT52UYW2ztby8yCAe6IpDeUgDnRQrsdp5DVO9vCa3sWJvuLeBaucoVQC
C4PdNn8sAJnSuL07+yV+yaTI8T7tMT/kjEqVUdZ14GhhPXtIRtJrAyYMOc44XSKR
GdLXwupNspJwLzZsseqTDch/BUPG0CxVLlzlTZS5VJoylqvmVQqYw4E/hFpX+M6+
8aF2JKvdR/XWJ5hfQwIjWpjOiJQd2yJNXylANeCt9/dhP+lfv+v/JVk/F6m7v52J
7PWDHZlnQVG/wBZW6BTzrcOOuyhkrgFWPbkKyMdvd0CETnSEKqOUKbbJ62jxGspn
h2eWhx0zyy/u9H6MlNgOtj7R7x/BU8DZWwzc2YAF9cM6KxtENN2LG+Ky6bfVhVfU
uy+1XXWOyRU12GU2x3qdxIQjfc/rlA5hV9RPzU9sIcJbAeUUZFKLP2FDKLQ/3Ykm
poaNEUQVw1rqQvO9s/uoD0d6OJ8hl/tSXmnwrMH/PKAK+6tUJD74Yh4xchDtZzEp
+YjHSpfOh7u7cyLUSrNtcR17NIUJ04WPHU06WrKZS1fXI+uGxKHz8iY4syXuAkW/
Cc3H3/huyu9mYfGsQpvXJ+LBe8swI0uHJwV2O+SUMJUv7MfpwIXmcR6+dFhXxpR+
pn3atVEaaU8DcuKQfP5/wcMCHnPYywnUj+hLZVgoPwE+7lTehhdZBZVFvhhifFom
9C5MVCdGltcvVju1GIKY0TY01zNyPmtBranvG0EEyOvXonoK52c8gI2J3FsCAqW7
nt6peXKa/thhTSZJyp/KVoJYGGAaReAwaxeDuVny3BvydXfwWBJ41Ds97o7rco+7
rexbZNGi10+pxLrUPVjiBuZ+C6bT0zSKQshyJntfF2QfSG8/LzfJ3GLO8EN/tiX4
Aic9PsZpMBuvonIoIzpz5nZaKl9RywsJ2nPnrbrOdmmBDweg33prJ+e5yonnj2Ca
Ahn++VVkGwutfGJwRwJmsK89jU/TZxb6qTn1Ga65qvf+n8rCh25iyt/C7OZy1MJu
aBws7IK/xmB/Ug28ZJnmeCufz3XDO2O5Fb9kIm7YSdPzh4+M4QCQc3pAiFK/+H7p
uVES2MY9v1d9rMv61f7Zr5AICl9K8CFEz2gCLHlGI7akBWfjvcROJ9Yqg+n/FDaV
uU5ctRmHQbRm1v5mSAqeCoRUb6e4rHWrAtqM0BS6z6KYqCc4lDwwE1d91Q9YlCs8
vykl6HVG09T4LFG176Fprp/gI2zJrHcz/c/JQBJn21OvWSrdubIodgQhqFH4E8hn
crPZmZL2nziuMrI0AGMaxhu6gmSTIm5v2cWw2SgmmsjzRMVdjbqdeSyjDA7x7RMF
amI1+gqMvsxOksUKmggEDJFPPuR7EjqEQStan7ZgbxCK1Y+DQUd9I3X/vzuKom8e
ENTDTXZ5gy2MOqs70Qr/u/RMXAy/C8hkABTdd4OPwyx5RazEMw12pW/5GSS9otKk
qBcNPuUcAwPBTu7DG3IpSHBg8trkarEvYRksvEHAHwUQnd6uOsf1qsSzVh/If/YO
CP3wRE6nrmgjghaHR/nFxaDAnu915E0FabR2k0KQ46Q86WToKRBLJk0yRrPv0k2I
hKW7C4FgesqPAVOL/pMBvPkkXkEUdW9cr6ojLWLHp0Xm53EFpaBAFyFhznsNgkzs
0BnID7QX7H5sHAepaz9vFbJbIkLFAQj+TdYa8kI3rELFLMBiTf1I4hKcdN+HdOBg
iLEGKOStnqj1rStKVB8T1vaX23jAzqiXnzDCy2B4NV/t4ef2qVY1L/BVVNRf5WtO
sdwjpuSXQJdI4j5+kMNkFunkEMpDNpoiOPJJE8Lsa0KPrtHNYRLoo3qFnrwXJQNU
rO+pNoPOhvXQKECi9PUZYxn1a7v0j+eaA93AB4FDdYA0i85mclmgvoPDf7ZYQoIN
41XZ34oQWJ1Zfe95l5V8wffo8npv7JtdQDXDnbvmyUqGNmTSpNciX7I1bnSH0p0V
SMVsLe3WECkC3ObJm55JjhA1LBz2VfvcUugQlz3tLcZnokx57G5zb9ExwuwfNrk+
SzdjZaXcXfFbMmIWMjAaZp803kDKpcgLoNvPT4S/zA/ethpJpWn2SaxtOcZPaikm
HDyezLaoR2aWSdMBZSCkAuExDgYfPRLN7bBFMB3hcYZFrQErOm05x2TfOGpiEXKV
iAnke690ZgAR7KJdvm4jEaznRqK+VRYgWmNMDSakWJlql9grBU+aCv22n97ljqQ9
Q6LO8gWYzaYraiBhEiB/VL/9ZqkzBu/mtar+0SWL9hs0RQoKDj5kSJ0no2uOMoNj
IvCj+KHR32j4G4/DuJb7kG8nXEmBO4hoCk0haebtGrsxIxuS1nC8HO5kT8XcoG5e
5emPDLFKRwAA+EOcfp0b6e0sMfav1I00jNfjNY+dfr1BHTR+Bw2PIyNyuHCgwSKk
xGJM12pgzTrackmK7xVnsr4XbcY8vZy+Olb+Vxf4paMNvMKrRtwKPrwaLN7i+8af
Sz1LlHOMOTQLG6ug3+gYxLq06yNezZeiTry4QKzzTC635iyL+c4/vksjrXE55siN
rWxzicS8HEehC02HbQ/eZQqFIqpOykVZ2++JoB9EQ2iJefrfHKxV+jA8qRc9cwpw
V/hPiCbpEXOPXGUNfYNj7m0sCujc5qbnj9xAxpZGsrVSOUkygHWzCUGKEYp1TShN
p4SDmBvpSjKmi3WSH6aBTqb+3bZ5fOJnvahUmXy7dz5gGcQDNcKwKCwM0/p0YRBF
J9lvmCLA3Al/6DjRUs9Zn8QuwsXA/sh0/gAOgI11cPZU/aPO1eek79RzXojhOaGU
r35zyl0wXSjGOumc/LVNpzqf2wS3g8BauMz8J+JovP7dVZOFi69o1f+n+YeNcKWI
yxtQZxq3ObC7GitTrHMsKjVE2M5ARWle1tjAv9ZXV5qxVfKsnYvhPgLY2t6csBr0
snuU+SxOhTUdfnGRPgBmFVPDnl+UczyJd3u3SgpBr1jH+BJKqn/AqZ7YVWduEu2A
hepiy7ZaFhahLIPRR4K0Gs7JQ1Sw4VOrtWjvrvR56oL1kXLGt8bE/fd8NGqDhXJc
mGO2bLFTkifkNSSBfxEypC4t0fPnepEZY38tGq1PqCYP40KtiLJtq86Z4TmT6t7C
qKy4Or7Yv8Xqfv6Q6rg27S2D/FMbO4xYUQE7/ZyLtaIeLPUSkqy1xNMtDjlzbOep
1LmGg7WDnDf6nwhZbN9Ar98XOas4IgDKa8LJDXcXa0rUNptW5+ANmchOUnS8kSM8
Xerqru5gi9xi4+iYn016QoZ/s/YOaWzeAc+61bDozJ4h0VnfzMYxXZCfSXK3IZNl
kVNHPOzpXWaCMbDMiKAxhUaZPBN4cTi7FBuIdcLIZfitb39t7blDn2qP3c/wPnu2
UZR4zttLVr6Nn5rvFBQR9osK3azifPp4nYvo5TG9zjk73vLM8lmmArx4LYnTR+VK
JxuypNhlJzvTTgLYwKZuV9bHNvM6UtkijumS+z5QK0e0XVtH9TN7iuCUSxG9maJZ
pOjp5FDk/h9RdiTvIG89HRUl18WwccNckoL1wdJuWkjPTJHwNuaR64Z/xBpYGw0y
U60pjlmda4YwPrK/hZZ9oDgKRyctNTo+OFXra/yxOFxjPNttKo3jW29afh68NkGg
kIS3JmPTosJDl7s4Cy4a0/hB4YGlJoXWSc8X7ZWx9vfw50N358g67nZURczR9Q5b
wpfqxydKxLKN1IZ1VAMRCGJ9xTHO1A0mS8cQNLeUTX+SrGxU1mY8bSnz/9BD8W7k
8Q6w3MCzGRiGj8GN43Uv3+u5MeZ4n12+Sz4wkT44j3TbyxjwgW5L8iee0KGRVuBb
qV/Hrf2+ousoVfvH18IBpLKZB5WhKtqU1Ocactwon4jUvEge7P0Gv5bakselk5gN
VVSd4RacegV/0ii+dVU3IHhhSrytyiuGq2YuL86XEk7lfd4tb7dgIcDuk4h9rrRe
N8cu1tUqpHVXhIN8MN5hNr20/+Y1S5c1EWllw2Bg/nd7iKFkJqEiwNbVM6hhuxSs
+YGYayeTlqLiDfMIcvSmHmgz0LRpyXBeyvC7yuYJ7IIS8GVWyGk1Udh6Vu6Wxwmk
fKutIbp/eb9HI1sQP3yzWhA1C/Yb28YeqCc96h23LWlQE9sa2Puqu+q9O6VZWvYT
ktP40j7FmDX1VLPppHjjAt4hVB+5ETHSiooH2PC1zHtWAjif61oy/tFLH0JZxHXT
qslnlb+rCMEmrCtsMIwjLFBVjh7B9Rv/6TnU3rhFJn/EWzvkf+EUXBvB0fdvPDy1
i44EA4A0NN/98RiljcddN2c769QhU2PIxMTFg8mu0Sb3PAtJLJPmkmVFZw6HSl6A
fGuhVSiBAHUA+uKaimwMqWremmcTgiSuJcudtFFggs8ejce6Ax1yjwsNwC/Uc1EY
IUdPmDTKHQ1+lOfdOL6DYM6X0DqtEsVLoY+QAzJEl+QKFZH+8Thi3OHIa7WZvL8u
NYE6UNESkwL4UPa0wnr/QoykUdTdO2VKSMjtiTbcQjlFPiMQbF8nMgyuiAd2p08p
3BEaLvqID3O1lSxYRTJLN7cXAvjv7vkI2higdwexTZgXuWhOgMoaDotKt5EW+qX3
yfWMtw/PRE5AtwRYRyzSbZiVOJiiRnq34BSnS6kf2pKyDyIy75T93gvK7HMMF/Y8
YZc0sA0nzjxQ2mWdFduxSu5qwTx3m93rnLrceorHHCKEKNCcEnbladWu2ZeoUQK8
5snFPgbYlIBrxmsAF4Va7CPK2kvMIt23/qlzxDw919AdtZ9jL1jpDRVi6zXCz2A/
KV6rCzcylmO9PH9Rt7UbD/Yap1sF+oqhLAeBhP1vEhNs0Dtuygt80pSAtwIXPTTX
okYeM/9drXANrx2Vl+jFQkOA/10xGX/VuMe/oD0lJVFAEU6tM3pyWEvfmSPiqq4x
IbomVIPFrPktvn0idAXs7/qdkk7T5B/XLWRvrwFZDizUO8WvT5fB6qhIYgfNkvy2
q9T0bBcbjast0mjG9KZfIeyhs6CxPa+feymj84pntlv/ZDWZ0fgRlNlh/rZa5Khl
euuzgobaXjoCA83j+4GHL0LrI38qcNBh9mE7UikBa8PvnAeuAcgZ+lIsLdymJbB0
tqwScpSF5NWB7R+6jqm9puZPGShUwLZNnX+jzfhQOkCwMJQ1KIm7bBL2TWYA+OFD
PcFYfeijODg2/HNhcKLipOcsERCB3/S6JkqvedfGfVBFzUkSpJUa53FJH6v0rzfw
3GsvL17gbiLxZNsb0GbdBOlZ6Jb9EAepakzJX/JatXFB2yfUX2/638tFhYlakr6Z
Em49dtMcqwqQig0ZlTg78mXcZ5x9trdfRW+5/FosJsMmUqxc7yj/zoILnl4Jjcel
8qVP4W88ws1KXZ21sqattkZIovgkVvSXV45+sXY8xybX62jfDBPmnL/OZbnwp4mG
fM1WrvApZ0P119GXFhjjRCnLh+edLJTpG6uSdhChVAef4zQxh5tPTt/nFqoHg+su
nyGoR4SWuglzlw7/w9OeYUwJ/wye+M7VYJy0NCxXkO8nmhdm/Kn52CJzcoOHV8qW
r72KB3QdFkgN9ulifjncemNbgxdEMeJ0y8RM3XX49IrsCXaWqtxO7EEGJIHuPQQ/
H3EXgRrjRxNNX2jn7A9GpnPl0+Nvyak5vC03b2MtKC/gdQu6xKynQNYX9QPYjH5x
F+/RgKX5btbPRF0XnyhNNv9DZvGem8e2JgpiU/HEOAg29tRz1yhES6khbpR/V+Pd
Zj0aMdBe67Xpute7dcNE037E8Wb0vUmfOOFEgHWC+1pdh6n+RvgbumK9e3Toq9WS
+c2LnDAsP8RWTQKv/236kJlAyCYCUlqJdrjNjqsDMPwNjTN+23+TPjLlTnSp7KeR
v5gygstV+cRymcbWnTPbeSX7+Gv3sI6yb3vMZHLgZgbvv1qx78WtqnAq+JKojo47
gY6IGMP4TZAH/tAztvBmAXW8s1fic+NFSAIQAqp1Vj3QMUg35CgUvhGkSH+5YnYC
QQFy7wQkTpWk0niNydvSJecve+wtBRnNvh/LM1E9UTwmF4RNpYoclVY4+vjBfSdm
Wfam0a9f9g6EJL10adLTdkKfBhz10fvKHjJhG1NvEuJVxb2LuZyMeUHKKBJaJK8M
MQmCX9vmaNvU6I3fhUcm+cn+r+EzA6tj/Ap7VzWoOx3Y7PDLLsuQKEzNndiwOHCW
3aVPZuMlEIFqxYAVB0O5jboC+5e/kL2e2mDeoiLJmjgVCe9JnYWSAE+oqg1p/n6V
tUKy5ccTWpY5iZ89uUKracKgo7DZKeZlub6ntO3Pl2qx/BhBNdxR/3Fx7yqSyeqV
52pzp8CJbU7QG9yD8jmxKhtkT/bCS+Zjhz6qCa00VIfD5NH1F5W2zU0bzKhrZAWF
xbeRrEjDkTMil1OBzK6RP4BzjRfb7MLVwrAwKQd4FVk0e3aQOFyYnXf2gIpwPJ0W
ytdbUBlM6TIvw+Fyjazy3Q4xQjXIcyQk0o3RvIRFpG9d3xFisPCylGDzaoZW5zPk
MCI4HiCQpm8W2NRmvTxC3y6xLxV+v4jk80jTbIBv5jI9bMK9JHepXYT5OsIINGno
88u4d4+bxr3XOFjXCQjjQLyeY5lT715S9OzsUXu8YDS7JJ3I2wZTxTMe5P31GiFB
IAHhkkqh4X5V00UzE0hUbSTuR75sj1UB2QQ+TqH1pXJe+Cp3Qc+3PZyGtzq69Rlz
lobT7Z+tHNHpdse5RI5w/5L7XUdVPvQkgPNBKUCbk/1ek3pLig5OZEUNwdUTnWHs
ojFO6roby/uYgjt+9HQaGE4TeXRjAPw6uVMeuf/dPS/8roiLwpQsMNXqb9MmCdvE
3PLy7LoLfJLSrvHShTPBBoF284VnigLa25rQxqZIC3NIVmtgZDi48xxcLW73vpiA
8pfqBKg3cbqev06IKRrol0vzolvGOd3zjmWJpilgn12RUof+gzgQ3pHhTvxtCOfs
jUWIQv6hh+Audd1BcIi6Enq+16wEYyVy6EiGubLZ23rp/Uvhs9MOq/HIQj4XWone
2U6+oMG1PA2hT1AQMtgoPS5mY5zhg+XHLGKgI6N6g3Aa3UsHIyjbv+YcTzF8JhXx
DDJnMpS0rJsFK7s8AqW/0ODomX8pFuQjx/BlWFvgps31KKIl3KlM1gaoD9/gN+6F
FG3eYGKztR/xz9I2RVVmG2hrki4Gu1gxLc6XFM+DaDt9umcfgmUrvfgA9OXzN5HD
EEI2o7xeRLJYl4RicMhUrfvTH9CniR9qbicxsbcgq4BPhmBViXgPWWUpGzPuLLpN
bUtDIJPqBAzGrYgrxWeOWuhWIjgCsj1zpG7dm/tNoIP+YSyUSliYJSrSG6hNOhDs
VG1tdPfgcXDwHFxBflotl8t55zAFkDA2cTFdOFIw53NGl2Sz8EW7mLqcT5lKrGV+
+BpERGcWv4XA8O2mpgpeBR0Q2t1TwIAgKTEXf3tm7KyonmYM0EhlW9LcqH7Q+Jtm
hGpK5X/74AzNkie/Vd2RvIzDb98qFDeB2CyaH8Rh2YiTNz6LsmIjfFRTkPZLfqOO
spaOeqYqKs5LFnrLTl9QlDpllTvqKoRDZu9PrC1LRSQJXoC1Rm/tQThDm7xyoEYo
/WIeG4ZBJhtT5FQdu/FHd3Gx1JwRVjUVNM0+OKYL27doVEPmZNG0wiEywXs8O+E+
heI3Ukisj68vSXj16ofts8lcinrZ7UeE52VMqC6Gq7zn0tkxWNyy26YFp2+WFWzG
mZw9XZGm+LwnIvHaYIS520v4LU5l/E2wsP/DtNIxuy59l7714pTWogTkb2cMwLjl
GwY9b8EYDBkBHw+F3yheiWo7od1q9n0MW9XZYt/toJ1d6yGd7Ytcj6bHpn7r7plg
U0Sa53XdTZ88uIgk7acq3acmcMbouL4duk80gL7mbRMWV13sIJlMTA+wjnwKxJG1
gRWNc6MxvI2BPXaSSXd3NgSDria4cM1jYNM0Zny4AzvFi1sf5+VvAPOv8sei4ihA
lsV+12rQBGzvNs5wK+YM8GjsZg17Gg2XJEDcnD/eOeP4tfcjON7PKBk4cr/GpJBH
uI8kClam3mKhrfFgJ5T/0XasktgoU2rWK2qD3L8HBtQQJP8iZYzf2U4ScJx20wOL
CbT210xgomQfQGHEJIfe7wf7CvbMHEkDI553DQ/yQF7PAOLIz6JfUWOKQPjkpSJk
vSQTOM6dejdr6xuR1PPssUce5Ou96TwPM0hnT5SkYWZ7Qr+BIt7Xy4LEOcVK1Aig
mEX5x8dRdAktp8Hq6SCezMpdJwDCs4UGvXOd2XokQhQdgapWl/QPBnWdpaex9Mag
qIdEmySyzdOJbC8BRxaZ0U8aanOqO+AH3b/pTW0cGTNXV29irtkahfmIZW9TPp5m
47/k/oexurSnCz3sMvw4PW04z5hO64DGdoTy4KZKLCYGZfj4UCOVY7nzRLUIfOSi
Tq7eoITEguJqH4Y3s+fbvKxSuGwnhPRUj29IWjUZFQ9ialIa8lEU9uOiJ3oqlPtc
QXzq3CBFz6hjegxbSoZmkfFOt8SIP493gYUKfrXXQ0TdQzqSJw0N3Oz1XkVAXVrP
VYbNADQwRQG4Xktte+UI6C7fXITE/zAGpJpVR5Ty1+Flwug+IDSyj+2kbZPDez06
aRyESrd9+33l3zrz9bbX4NnmAcQudF7BWPMr3riwU0/Me787Co/U+wNVLhgpQubb
4KLAwVQI+d5wMdxELCTUHJQSqSfYR8tuEGlDkgA2BHbHfxWGbGa2p0rqUVFsFeCu
iLmrQvz3d1B/6sIkQj606YBWyr7bjF5CN/uhirsdm9sMNlgkvWGdU4IIODEUio1u
Wu+EiZdkh2k3ngYkGWe0H+/0/yZXsbnYkKTBsAg/oWWfSCfazz002poBP6q6z5va
l9oUH5ITwckEpg2Z7V5s3jWkKx0iFJnIqfdkcIVJWAFt/13zxLFaV67OE4/0aQlt
WZtO/JP+6QQSDhw/UXutn4866Y7mwYJGZxQ6g1YmkKpwJJzbbJbjtsKypP2LmS+c
QgiD1qD1r/E/rcrD78Eiumr7I/2jsNJjF3X699sv53SMzAQyI8qdMy6vulFrJcDC
bVGfHajgQQKIjvR7s4WGdmK+AmXWuNhW3+D+eTamJmN/qmT0A2hDfBxYzPzyHcVD
SmuPqPpKyaiYnEp5TZCMvOP1fOHp/lZWYCbLDy4cO9vhJS6gYw0yMYCOGm3T3ec3
ICUqK0KfMCQ+LdA3MaBaXAX8OnbB09fI28uhAbEUROClUU0FY1u4thiVdUTXiAcb
OhNu6HVsEJFl3yiFEDSMQxBdDI7xRbMjBqlO+qN/3TgUHRJo1Vd5BYhesRZBIE0f
BNrECKRncH0O5BrqumISUJO/xZWgbq3kW1uBXSKoGHfYtaS9LZMDaDGFY+5czgN3
Xov6cpUjGy5fOI/WeJ4Yw+W/j3uD+nsfruruWxFBTRy5dYrqJnWFpQb4mMaVNHXc
hi9NgltbF1SQkeLTdSPSXdKCFRkOTFxAOLKhENi4XRSxvWydm2+Vbg3LSXQLwx5G
eLL5x06+mLqULR/wTlO94Pdr4qAOC8ibvZSY/d6P0kUg9Q8rZgJPuaKpg+LTWU3R
NqjIQ69S1DuYhkOIyxPP/EhD66HuK7/Njp2Z+/ZSimxpNd8k9JExs4UBSnEFh8y/
k7ij6aFmfTIxD+SUyXuUI9F21DDnnlO/ounT1p1+UrxzKLOaCxAptKbgGs+NQFei
EKf1F/ktj/svKAyYIhcxt0jgnJq0B4GF+UA/it3hWOVTMrHxsv1uGAKYodBPBih6
mD1JfLZHQjfjeWpYkAvN6EfZecoMaw6WDT6rbakH5gRMAB6/DI/t2PbLM0AAkPJI
/MavriEUO1kDO57FpRXhmg0si71AW6a6cC+YI8ydDBMqzc1K7fp+lppm2yazB8I4
S6gEFsJmR2aqypCrjL28jlqH/ycnHeaTNmxoc9Fuwxh0Wos/hxAzZsN7sRxj3dz7
5EuM17h9KQzC/3RT2ipN67ythidWjzpHt1ZOuFjss/XCKz3p4iQbyaqTxoTdfUjZ
Sk5UvccGUBbSMqSZYmgUTlLS0tZOvrfRsPy36znIIak9PLJ6VZ/r4mEAqk9FFDNc
kR8s3X9NlrkIAcaRObtcoJK4nPjgGLGnsjNizIupdQRrOLIVmZ2RpTt4vy32AQjh
rmu4UfeSGMmKUyWmrSutQGxprBCFu94kzBnkeMXRW4WnkX2XhfYl6UJTjwG/bwxq
Y1Zaa18AbLWAKBRMYsM9XaAHQjYk/3G/pPnt327YOaDQHpWF9NXmwlrx48w7m51/
hUcbkr0durWV226oach1bEAywbTTQS5k8fAbvFFOMH5wnSgtYW3dn/ijy8ZLTqBu
GgcZ3LuACzblGZsanLwD5GRkvNeWbBWaNjLhzfD1BEgd/uu9t2PRCVCNIJrE+pGF
+N0NqDXt798WVWfQZcKqUz4VFun4eRA6Rt8Gro+gDu+ste1at6M5A9PHf093cE56
XGo1PMkWJJZ2rM4TP+kJgd59WcQ7fI5HODDdxPS9Z1sTQFWInCaYD/k+5JkvMRQt
EKhM3Ex9eTVXckwFbXo9r3/ByM/rtS3vSv3DOP+GJzoJAJhSTOkiu8MW3wNC7UgX
n39c1ew7ZeNUvLwPWmZS1tYLkiZUasNE2MBGXMvPO6Oyltw9vHgIb6WoJ3rNqnFI
w/nsIZDm84RZ5pZ2H8qzd6MzH22YtudNvRpQq7heQJx4z1akhfCdpISqPPNF2fHz
UZd2h1uwCeh5q8gXjeou5g6ihgawEGZe/Hkiv8wkN60WfZ1ENvkPwNxJqD2q5jBF
eIZLZcZ5z1IKSO+2jUUutTOeTVwbtES8a5t0V6owXqiFCraUC41kFm6iXWlFYbUV
TtauFBXWMOeZxVo1dRsv1D5hcDxL6VN8KKJTGGcta6x2vSRUXPNNbbW8YOxSsy0Q
Zleu0idEA9z8S3qHCIRL+4eL5hIqjGBmettIKoh//ekIPqL4krJLPl/4jmzVDYcA
WCOXFB+2tNtT55bFNY1DZ4RN2+bMxnYqeru2fvqBsIQaAso/ATBXUk4JKJyUXw8z
3Z+UjJsIG/9D5ze0f52MwdHLXmkZywH4/19dR4zSk2JlkZf5K8/eN9xWXLt3k7eR
rLnNS7guKPHhB3GHeApdvNoAW/A9G9/K1WoDiYHaOVDAbFkeocl9WJnYb/BBasdW
zDd5u24dTpAMaoLzjBBf7xBoMXdY5Tu/v2yz0aD1sRML+m0CFS7iByI6Yf9KRUte
YY08XqYKM7oVgl0YRlljvsoNdocVAkVNtXHChbzfF7vYIM7hDGH8Xu7/rauvdahb
TjTjir06ETz68NC+8XKz+YPdv+gGzBLZqiD5lFJ9jG0crGaYQMLUX0M3H64Zui9V
u28J3qgsdVrxjvpG1ekKk/SEmjBeTAPD9rjcwueLHG99aej3SXLYwaWTz/MtTXaH
dCN8K17Z8OrvVqIDYGzWRC+eKjUVKmLnTNLK+dI0N8zND17qdpqy5CaHwZwNw5rz
gTuM0x6mGGw+zYYOzqeGWyIWOmw0SRptuns9M/m7sV7/BB2NaEa0PLy4OYwbf8wS
GO+Ztv51Pg1h5tOcnUM7HOUcl7OXUAF+k8dET+gsd1jyEjRnl4nw9d8P6tb0L1om
JMDY1iF3PtVUdDlTemxE9tfXbDwXrB5xLz5WSt1/HY+fnOUQ+BruC2GctOgAvQ6J
c9CAse4FCfw25fn5ASZc1rHppVQ2mzUqj5tSB1k27Hpp0FH2ElfQb0OhS6Bgq1at
tSuvRS41UQQe4uegXIWJYXDQYaRHBJzHNtSeoNwdoUfGQ8OBYhRUSi8CWT+HjdAA
XlxmHEkpP2JP2Pl4WqwgFTDcSbKInoNoN1m+h2YfBo/y758w/B0fOs2LNd9I4p59
1Uq8PCNH5y1kUxyLen11BWDAOAmjM01dYjUuW4Euo84ODmoVEY5sbG8zyoSIv1FQ
AFaoCBlTAIK9eRCvakFvHGI2JbjkhgnMRCtQWGw1TIB2NX5UjCRi1qtfmLAbAyRH
CBnSF2c1wsL2BexNreuocTCUhRd5nyt5uLtcCjk+cmlK+aicSftCF2ZYYxEittjS
umadP4uM8yUZ0R2vZLOXAkBzSAil62tv25xfLYTVfS469iBPi+sev0p1vlNlsJ9X
E+uCWQ5O1bD4KVAU2M95QdPUhQKZhT2EE5rrq3iw+6t6luN+FftpSBl94/m/Rmbv
cO0JwRHzyG1/ArNkQq4ksxjbeeB2ZnVp4usPeIRPMK1aVHsR+U9sQWyGB8wCrUcv
sO8KFlTNm9rTvspDGiRJQMZx4NvivGcqsfc637oKXgMYTRuAUzw2U1gB6iO9GrDt
XmNQ+uqqi2J0FqSrK4quc4kWM9/JCtfgwp5+KYsZCxMtBU18ppzLRC24mk0DrRSF
Y2+W/0z5HF5BU9UcvL4eLXlaQgOJubcjwOe9NRjVMpYyqyrQexMLoUPBZOsbBCdW
mb1BeufDRtkKH8Wl/edITzTfBQcpZyQrFKmoM58nF1ekCfm0juELC4y96TMCarvS
R9PmNwnRov06C0hRCuCRUMgYh1X8PRM9LVrIGT06jxHRoMUU7isF8Q727U2Zx9xi
/NwUCVV2s5UdXaJ/jc04stLmq6AovVUl7FcVw+fsEsNSy+mHbi7XWgwP+J8PzanX
hsGB8o2Tm77kMOGpcqAg9xOVBKiEU8koh7xMB+fM8GQrS/NjvAWrggzvnXXJi7QU
W3tW94uZua5WzjRjVhSUn8dDd4HRly2wWrdKURhlUpC9Xif3obA0mf8gMcJqZSA0
PBU+ePNN7wQcNymgnweDrJmHA+ZI0zAHqwlaZiJvx+ZJmf9W9198CULqWGl8N2Pp
iOn+HeSk8kkWSncnoQF0/Zl7j2tq5ZLtihKa1awnTEJFXMTxN9z54W94IvXpZiEc
61YayG18GwXSwm80AE1lDVFhdI2E9Sxm2NXUxToh7L3PHMtiz1R3ZzGi2KSbYnSM
89lgrJ4nrm1r4UQAEj2EtRL6oYI6ZrpqKFA6dPgj2d17n+qzRMuHS7nCdkI1Mqh8
G2GWzK3RfTY+ix1emqhpBzjmwWk1nIpgg9lO1LICLlb6SfGGiIrDE8B92/Ifzinv
dWPwtKhNwhU4q5ucwvrowxQgBu7F/D9M6vBTyfU0yMGT3LiNfduXnk1NsYxws+3X
zrhwUURmhppXeMUF+KuRkWmtMCoRE9+en4w2dpDzAJ7d/JzkU+uc6XdBxKA2ltBD
p2l6bfyyyXteEx+2hqYdb5wA6kEke/PeiWp5DCqP5VcO+e/Q351T9DT39M51xeyq
aQOLGzU8rjures/zqWiQkejoX2PURNxT1NlnJX2oD5SP7rU2fVfrm2ScGRE+pCPA
M2xkpPY6SXG9KVb4l/hYqlokEQdEFmk0WSpg+/UaYU2EOHCqdIjMBFsDlx646wHa
Ihr5eg6juJUxUyfnPgql1u/a7k8PGH9i4BrTbvwRtufK4AjVVWLeJgbmKEDzEWLv
dsGLNh5gjV9dwOL3VrxWuL5rhakXUi/+cf/1J+gq9yW0Xxun4od0I562uV22sTZm
g9VYoWng0Amu2BpACtzNeOrt+pldVXKUi7t+xAZLWiGaT3p36vMKWNjipTvBeMm5
9RU/RUkqiZD3HHfj2AffOD0qLa4sAcqCL6ui/1zOOrYLu5pYBf85N7B0Jmqh9JAh
JqU1el2oFyJYRVjYoR0Kx8lNKukixpxoRyVaCh1V10uwXIknDcDpb3Pire2hGD1c
CAdtw+Fp4VPK5Tc/qfsMcI92Zhq26LMQ2q/I/rn6VqtC8/tl7wlRSzpXe6Obsdgt
nBjVxEMWdejJ89N/LYM8GZgV/XtLxbqpRq32WJYjnLZQ4333x4Cc89tXrt40Il0d
wyEohRUoCSq4nV5WLi4rYUTU8rEDvrp4fXD2Wj8x8V4RHIW/ayTOtflnDRwEeloG
b8wAzryFU4gBT4pW6PXfxxoW0CFvkpw/BwJDAQciYz7YFm0JDf3MoIJNyMhxuQOL
/pUVEEfc9EszOZMQRfBbw5u4OYlPfBAhHL3ECUlINJsuHpfDJrY6mjlhY9KbhSyj
S1Q7KJ534YSsBUXiPdjT7mGk9S9NydhGG3UmFzZ7zZiooij0Luq4Yjo7MKqWIgu7
RnIgU9FEJ945+EvaLHJ5afeGHikqGXGSi1w0J6vyA+7CoYfERwWZc3Oo3nXZ0y9C
ixywFpdU4hxTgTyJZxXLnPkUdLoB9ClG0WRGGAu0qEJf8WejVwdK+GnSXRriXbmA
V283p4801ezvb6GMzEltuWEqH3TxbTSGQ1Wj/RO0OImPSNUIOxlq4dOOsnwimInT
lakf1bvGZQt9rodZIfWmf1+57PidAo4UBqG9WMzfW54u6dEFn8/ZyiYX3Uas1saw
8uXH14T72EAY3EfHQq5NpQmeeJNFU01B4xw8pUZCcCj3Taj1QzJ5CSJx6p9A9VLP
Jjkb8ZJWtYlduWj2GB9yAGDISTzgn95eaHlUahjA1ESH2D8wAb/fnLwcvR1Dt/OT
K0k7X+HNJMBYq1r2TkWmtbakrGQ3ypf5R0oGiqDuraOPoBGkTHFVyJ/GZ0NySNAn
hIhe/4DYbOxMjyJY0T+Jf65yL28vK40I4ZS+IXJbdKYHU4Ajlur3IBGNF7L4hckR
Wv7AeMbld8UUXUZ3TFmCuHowLLpb7Fwbo5XDgdG64SgQxn+v0ReFC/fWIloTAoqP
opoSFU/wZm6FKr6WqtQFdpviklsgwiF/ak+h31cASiXbpUAsf7isxz32IvW3enru
ZPfTkibznYVq2tNhTMeLo/rcb+Ki242SP17PN5e3EknZYQANg0kivtU2SfQmNfHy
/tu+eECn7RKITBMPF1ru00zq1DzrgFHZntYU7cX+7svkHcxpqusldECEf8B6HdYa
qKliYhajqpjQXKrWEQtcy6/sTHof8J6vXJWvEylAlQ3/fuQmXEZmKjiCqJYb2DwI
hyCvk5prc0Xf7GV45bQuAD4Y2jqoAxTeuvIqe4KsXSpuWdzbNovfcQ28Elh+EU+k
l2Z4FSFwFN2JSHrU2PbMKxcAWgZmxkHOj/7mzApDNNKrInCo9cRZ7/hjnSsGrgkf
kloCh9YikhwPXfmLI42Ss9fC6rQXp9awKEBo5eOJ7XVAAJhG99+Afw75e7cGsm3j
FYD0maExYaGiDvFiUGdkpDIa1rDiu6P54/N300vEJX+DU510Pm7yrf2eYc4hJL4v
nVm4BJ0AQa2QJOygMUj3ZENTPvHQ0LtWZ7uQf42Jb68/EDcAdf+4+0CP/ZM2l7Eu
3W/o80oG+PVyHWEqlRz+IOyKLaNsUzQx7vk1r+TTpeWcjzloVg+vxS51avScjM7O
hu2WKN7tjxfa53epboZFfBTbhYQS8qrHHe18xWutso10j2FK3KlWIgNN2//VVyN/
dL3Ac4zngP18lYbfb8vVAo07eX7n9USsrJQig1AV1B0Cf84M6oe+2VZPfqik9r65
QmPMt5CFhAxFqh/CO4Nzwz4RYf7T1/7HmU7LSzsf6hvAuDPszqmY39idBBTdsifY
jiKEtgc7ZzOm/gOgsaUXN0a2LW//QPQ9KcLI1AnOTibYRPO1L8I3FaYIqn7VyY3l
xorxKmbLQO8+wHK3cBjjaGeQSj5M/Z5/eIiOipkvXaEcYwt6XdP59SnZ4EC1AEgL
PxXANF4rLIRJr7cfEaEdsYuQ/7vsKfVz/wLsUn0mQ5ZjQ7xQRtMkVNN48aIIpbza
xAWSJK6wUHY6Xf/OUFd3rv08yfMWekiAQpM9RqTa11y7vw5sAGObYPVvdlklqAtI
AielrNwcAjcj9+8ek8yMwGkolRCr/Ufwp3riDNIg5QYl8gJ4drL61J6NBjxIZ0/c
2gPZ/MtxqTlesNvw/fqQMhFvLKSH1IS9y4DQO9/iLquaCWIb9UcxcV478fCiiAJo
V/caorS7MdWSQiCS38i+JceQ594yCHIDco05gKL/rC3ENAVM12l7aHpllov3eChc
TT+m/gdVt1KMTTuXlAmmDuNwF63pqjIBKF/HfkVUmsFpacdlhbJNtR3iZx/kvkuS
fBmesfb6q6NMyu2PX+KTfd3fNx+J1/4QLU6xj9FqHnO5jl1dxpdBk/HNlHV00k5c
BWLRqKYL70kmRDRCrmLf+3HOpyYF7XeU4iKcCP6MvLE9jm/QqzGxhIDQHWpCzmq/
Wz9pwPN6PJiU/ns1v9rCxuexR6wu7TPCrD3UMcUSOyNaOI49A4iXSJX+f5I6g/lo
QQIkeDnX2c6SfNlus8wvf9w/6FfkG/v2J502G4hiyCp1YwYPJvbAyNT2yHvFsrpo
8pZJCFsPvj2aRf18dlzP7aHtCW65wPl64KRbjc94060ROrVAgx2gligDGqMTvksu
ctTNnHHgC6RszoSo65teeXb9hvPm5VU3u/ypu0/eUZXkmEwr+a7CM8lrQMQ3x1vo
Z54XuYtEBEg8oOXCLjqqUpKRfCh5ua8XjFjLV0hhZX3uJKmq1MphKaUUgb2kxwtj
juokb2+ZaGB+ysFdvYQDCWuSO+2ZRIZf3u73SASoz81TISQtJKhKoF0u21mmcSoB
KCCq2NV6GiaT0C50mWtmeUJUYm6k6AuwLYjZFb4PheZKxVLrVP61LG+cvV5f0SQU
tyLpMbkWLpu6GAbq9sncjLkwrg1b+LNkexD+LdVCVi5XWrY1jh0r3sRce2X2htXZ
3DwC//oLc8JNxpNSd8BfrTKz9+FXXTktQ7C9ZmBakLaMXRWwl2CkZa6NMFjEmacN
YE/TXuYUw+W1KVWfYZLehldUoGVKrOpSb60GcpmBP/N3L7JwgRBwJWVrfOqxzg/7
xMaC7Wg0Ju0eXf+CnTDzyH/354F71jZ04H6we0aojSvT4+QP8KbobQdFnVrNzRsk
xO+kUDGOsyqQC9kl/MvSK2NVDjep02hp2E+EWQfT9Zx5rUefWjr7r2GPFTR2V/E6
Plla0H10n0odW3cdANTuIcc+iIOQIxoKizLBbNnl4KEo7kCSLRoofcUXyaoNFwBu
ZcnviBaWrc6qaDaHQ79+XFeuGQkCef4BbjWHxZqji8LrLBZW3ve1hsBX/BVMTN/1
ad2SZBYyBzOXTW3bT/cLeQKOpqZC06fmbR0h8pfm/FvvCFgqnqf2wDdt/as5GiKc
rG3kcnVVNRfQTtdd4DPaYp4yxPo6OJqNmN88Osb5oMezrbRj8KTuYJOMytTmUgw0
ZZqNMWPWXpEh8rZ7o1rMRZHukjEZ16/U397uPekYVjLig4v9xc6FbmMaVfYGUUBt
gTLylMg32hdxGDaKhpCV0H4XIOW96cIxLhdLhHxoDpkEKBG+GxrM+bGnjtFWeOMv
ruAsyvVB31HrUlrXizKXy4KpmA9vv5oe8gTqA2DDICcnXeeMCeUtOua/hAKqF7Dc
I3Be3IQko73rDV3EYN3wHRHW8MiMrbonCS98EAJIGnNT1symOCOi9HMuUqEirgyr
efOTD4SexCoIVfwDLZ6yjheMV4npUPUQ0ybPLY1aGOIHzl7zMkyJs+0oBAg38pbj
rBsv3taQcc7Zm9uqao5dRCVO847qNYpfMf/qjdr5YeARE2c45gDB3J2f3pLorFPP
KK1QqrK/LS7Rdisx7c2QJBwdzK33Bc7gp87M8V9NCFsyDaiv26GaQ9NR9OJrFCez
1+ClJgu91CAm/wc/3Ft/6FSTLhwYx8uf6fS4cFdZ54capAK0ScV5LgcL2RkfxOPr
Wp9HOHKgF82BhV7lSDPcNSKGeqpdDE1f9/mqaJ2LHHZbvVqKZuAiAko1M257b+MM
OMA+AETPyeQ1wwFMEMACzIkSmMw4aTwGuEcwnhUb9vjdDPHPwx6yZeSu9JUunn1C
q3mWYZE1Suu4zkhjGe0ZrRi0vhiTR63DbMaOXZYaTHjIODhywHt8k5jicDjJI85y
xF0dcjB3y3Q7YVkSmYExhddkatEYTkD7ciyAUy+ynHTLysNxWECIEc/7yioo6fGV
qNNmFB6yDpahq+P3IysucAtsPoZNM3LzplceP3g1XDc22tkM76irE13MdLnYmhPS
EdONJ3xCW82EI5O4mS+GP+fQMb33iaMFD8mlsLnq+GqwcovFW/Hbk99ORirqBku+
7g9iPHskRNB3bO8LWAiIvUsjYRkGvDA58F0fJ+IS7ERIVPYTgDtsGWZ9v+VTXUA6
DOCmS/Am8MAyyg7slEWJQj4xtFdn2MLuvhLvtIFHcKxAOnfLcuuOr1Q2OyyI1a8T
fcroWjJ3Z9vFC8F+7u09fyMWXz+Ph1opJE6dhsgdmwhxTEgR6S9EESdclFmBdEVb
wJKkdUIYaB2SK3SqNjgqHDPHoj4dkpW95OSFZd3ng23DZxE0w94HmrYQ4DZ55BuJ
xwiJk8Ln1c7+gby8rrq0NuBVUMAqkaOIjCXHyyAdfWt/qXh4glnFYh7EK3uZP90/
8MTWKXLCe1z3jsMsoOCUwaaY0wYxdN27m6OAocdl0CMv4fp7dDZV/ILZnBocioWD
dOaAQqkfzeunmVPIgJPoqzPrkFsJLwf491OBGNjx21uhumtrEeEOj304fQT04VwB
aW2B3//4N+kl7fYiwO5vs0YjF5hWUJjdwjvMjgNDLo7G2fkT4Fjnaj9u0VpJ85L5
f9ldAsR5+bsnRCrl+3GM5ucvjmW7uUWI0ZO03jkKum9Cwd1GXPOgQ+L1XWAyUUur
0CW9ZwQzIttF24oHdgI2TSKbr0aG1W8Rg4Yl37Tg4MvrHiH4sDK03kWuUteLh+lG
NCixZ4qZLxHlt4nmvQISwJ6zdI0WZMrv4b24uIh6e0ezHvzd9Hpc9b39jI6+fsVq
E3qLHKryoEZ6Btx65aw9D4C6+80V8Kl5RlW7iUEXVaat1glU+JBQN54YDkjhOv+w
f8wtt+ECOh9PyVth97t1vJOnMHOjc4weyFDp8R8ZxlKz+FmiGe6t2iM3uME3fZhB
L36wY1OJ91vF+M13dnPD5vTogAwseS4aUVId+GX2l6wE6dZsUgh0L02dgs9ovQSW
tt2FWBsilfqzCm3Te9mVr0jCEsS1gfHCwIGkFysPT/EQp8U9RFsDozlDpENVkDY1
X2SGOE1JJyzYphYVwHQ9FkkjaurQ+IR7fk5fjGBhWc0Jb0tKiluy8HMMSZv6w2Oy
vF8xGuLAC53qkF1SEq4vFMCJ/BLc+EKoGrQBidZqMZdeBwG15/EsJ3AiLfHsKRqS
N70KalfY9vk8owOV3s57IPdxG6PO8IyN3DE89nCbHnkiLAScyIuUd4WQFbGXMzwQ
1T9LxW54bA2eGLtkfFZXWcEvKUOluIpFDjm5ERf6lns+iPlo2wQFzWswEuPPJOdr
SUN2vAs8XFpr9N6HN4Y80OvUR4eFYk6971OJaeXvzWiRVFMnI4RHUTmSJr0sHkSA
XVZrtSe8tupABuwW3sCl3kOytPi2AwzAXs18B6ACh6KfRj9b6DGDckwOc2Xti2Jn
icxMmSFsUgfWbRZiQxqN6ekc9t3qqJgh8oeD2p70lxQBSuMMpNGbCf+FxdsLweYh
q2+SQKf38GsRiOSDvjP6KF+lmtopg/D4sDUIPC28LeyFS+Dbq92IKm4Bh+id773B
g0BuxHkcWvJMiPmHwjux4zV7IVM5k8MNux+Z8/tIQvaTE/u0ZjvRZvnXPWoCKEu+
U791ZHU+gqn/jRXevoLb05/bKpMpNGIS4MReoZyE8r2534L3q70vvA3GUkgR3no0
wJfdHcwF3ekQ3ORmITegyrWUsdDmav0TE6U5AvsuU3XeoZ5fplK9NnCKOoTgxeO1
hClE+8CNyzgl4NfzXd1nrsy0/91F8ZA+4zLOqRBoOD/8zDy04iokKonQ2q6lARSJ
THUjoiAQniD5W5IAj9HDXo1bgw+Pnog6q0MZv2IdMrH1YhKBObfShcUd3ZeZuuSy
jg5AxhLjhyGnow4p7Usi1omgZSkcsqysxK7xBgugECX+M3T2EFV80vVmY1K95B84
tdv8xMLhTLMBx0u5lyv0ASEHFlY2A1ZNILNUWCogu058lPOiYL7gIhbtBwWinbSX
HN8Qjso5ta9frgyvT4A4+CuEk9vWa9FTHVRe9L9JQbIDrBXjMgrUNulgafYsn7JT
wQrrTp2JIjuY5xxxGQ1yTSeUc3j/OjSQycJlB80iP/ftQaEisAG2dYMU+8KOhFqU
IK15yBuC3PjN8mQdOCAYU4zLxmeYj4JBlj8EUi65da21KtsIm46PK7FSRY7l4Nl7
aTtJMz+gyrghTHVAnmednz+/VQF7pLyBWORO7VJrqWMoKN8wEFek0G+c06kcB08R
pZEBvfplkmfk7ftXm+BujQGPtlJ4iWxmD2oQNmToYgy5VEZFmeJs2s8BCEPjhahX
Aa585qYKbg24GZpKozgm97bMzKAFvdOQN1c7w71Kmi/2l8QJGGVRssBfcltKSBkI
UoVBrF5sSWVv6TqtCHDm82ogDXRlBQuQ7EWo8BLl4XfNVwoAIqfqFB61sITikVTF
xkuldV+eyv0L8VpbqpMdEm0lTGw8y7k+nb/ZPzFwbfkTGXSUWJvB+HMClPDi2MPD
FKqU7Eexn/qbRuyOVruaeW5FGk/n0AueiDh/E5suOAkD2mRbaUHdduU6oHXU86OJ
V68qVf/gI/bml5Q4DpXACj8x429DvRi5nvTBHdlS02JIVxXdjc68/KdM2VNQ2HJT
33SVOjVEQu2gO4uO+FN5/PxzBs37417Bw6DGv6jXUqTTL2g3k+QS9noZAtSa/qIj
DjxKDat6UeArjwkL/tiX7sWM2VZuhvmf/g0kn1WNYxRjxW/VSJKz9Cqtrb8WqtTD
FMvsociu76CIJKVLlPcw+NLKdpDQlL8dwbYPFWMhuMz6QfjslC2GBWLoCvcFZbJC
gUOSVQZNggU5lW6Y1hMVfgf0grN8GdmgJ9IL6WPcIR6J6uOSq4BOvePC9jzR91rF
CL3GTBfEdfqTR8g2AEWCeIALLt2qUJ+tf1fhigigLBxWJRGyYK4DHE1CnvcF001k
EkwFemtxIy4KePnXlw78ENmOetueDvQ1ERIFqhWv2VZ6/oO3FZaj5pEIrBxpPrFr
Jezz9jqOlatlKuwm743UwIZg8CkuIZHM+kJ6QV7HLGQueGi3fe3sDQNEUpcqcHkC
UPAxfelKJPSMCUSRCD7R6uTwnB1xNCgrx3YOhNeqruRkctOz5DnkFSH2q0jDOFMg
0i+6HKufJDaXQBYi9cBTKctKGmkgHMMZRAVd+Gz0DKsprmtFvk/+/CS7XHo3fIxf
Gcd6LzgjIuUJu3QMG+RwY4lnXoD9rpqqw5KdZB3a3imI6yg6foUme8MwhmN7L7yO
p8McV3I2O8mudP9jdCzSFz4xROr7MsQk/257cWSZZZHGn/gMLzSeIC2Ya9K1zWNP
sG/EcWrGkLDDH/VBjw5DbA6YS1KvCvcQOs0Gs3ogI9ij4sGA+j5RYqHIzEwCVJM5
uadYd8j5zm8Zz4tJ5AdWnThUEj5wmvlHox5GCXXa9CtbSKqAwl0A2NYhhBAyRDEX
mTryuhmih/j/XWNeFiYMSqPkT7rc3/dJKecmcw0fcrRkLHegf3tgWNj+6PPvp5Qh
S7o1cD+ITNnTUoZKeo2re47NUKfR3wEZSWsa11i3PZV9nQZC8vwsC9MwUwJRKWZ9
9OXjc2qyRczKUZ5WJGwoxfB8H9wvc5OrgLL78xuILr1e1eDlh8LDnQJCqCOD1Qtc
X/jxPsv+XULCqro6HZj7KKy6FUg5yeIG0mZDwdKnGThD14WT3gHgpZVKKxbwyLTv
Psco+CIeVAyISfDTDe03TdLNS6Oa0eS5otlnLrG5HPWFGwduI98wDnjThNd1Gwuf
7T5KmPRWu2D0loM6v6P1YLAMhtaGJcpxyQi7rnp4T9p8Teq2ABCYQpcdKN4oRKCr
9Kjayn7Gao6hQ+xq3C78cJbcV5ZvBXDNg0kLqbjAj69zSyjHkFh0YkGrFlcTi5h2
Ome/dgrcJRySRGnUrX93c+ZlCo5VX14kyIA+oNYqlmBuYTNp8jWur9S57bQ46LGW
VKpiVnSgKsPmQxWB3tf7LmjEjqyutg56CXfoVgDHd9rz2m/384T9yMP4nXODFBBh
wYqQBwM8UFqclQ4sB1xhcfk2lYOdavGHmjW0vGToBrSkMgMHhVihrrpKgJZTZZq5
uqHg6KOnGV9FfE35McixY6rnFigA8Z8bMIL5fcaTBdNeLyGzD7NX8DVqKG7qe78i
AuD4xL93qg2hAn6LCagEbU5YY+5oVhrwFhTbJfHWNz/k9i57oY8PhPlOibLKVlf/
AanOSdq0vEZVSdWzb3O0v1lY1w3FOFPYHbfvhJdYERjTcToEBmfUc6zAWF93QnCF
ZVoHTeJSKBuwRl0I0bKoyEQcHMyaWVxo/Ye8g09cgaBN7QvcN8q6u6EkRWmJVFys
faqR3QirNQeedNnK7Oy9OewAsYu2JvXEuqHUqKFiH7yI6/xoh+g59OjEZzquTEQY
0ITIQ4Qcsy+E0fDs/F2lZJIEey/sFPd5dLRsRu8ZFIwPo97yoiNBhyslfTrpJDKU
Y86EaQfLb9ytwrpv1qQaeKnebfBnPNKBzo8hhNfUbr0IkwtskM9yE0vjJd3oplB/
uSGDlc5EaIv2pK8eMQ+Vmt1FH4xKwybo5yMrFuVQKmX4/zDDh8e7nFi8TEyyNnm5
T1ZaH+vVM7REjcc2yns2LZYjXW+qo4TxdU9I3jFICmCxX4XN2UjAO1iDei5QlRE1
9FJXjDdX0TrS4POYV2kUgJPXN9Li9RRtNSy9/fblWOqjAtHgGtmK/G2qKZHO5Nne
MeG0qEUrp9rO5Z887RY+ImzejA0Lq59hDCgN6Ms0WVm1uS9IfP/unHsVJ6MNLzut
c5Mm7UXVryBL0ZUeBh/eUHa8XdFI643hwzuVm6JvC8D4eYmgP/KS88kpEXs69m3o
svfVkP67CdJWi3HLay6NmdcoiyqdP8QZJ99YL33MtDsbpi+8O33DEfKYOnwIhP59
imszqNTIOFz0/zAJzSXnjgMM2QNYEQX9XBLRW8LaDMXDz8lmeEwqzMDERpntoAm/
p/VLmaYaRElwlJbZwaAakb4MdC/jH+Uy+MXejgCJGFBXRljTu0172oM2zeRui1Kh
EYL3DGrEDLCfHF66fDxUsSNHoEnPEC7bq8YwHBmElUnmO7pRRN6EsEEBCpFxDsg3
E64ZsUf2uvAoUBYUdpYDxSvl+USujJkAFd4svI6RxYFpZQbmQAtq1qSmSCyfHXqV
iH1nM/PvR8KuyzlFiuEgQWlKxe0wV/r0g5SG8y7XmJJchv/Oye4B0CVO6qJDT+To
57yg/ux2dVp/L246+wLaVP88oTDmz9EvAePE7H1KSNwwweHKo4p9UU3u6lLQ51nD
Qq5FIWBZAY4hyFxfR4SmhPAhrAh9ZFu3lU9JFA35UPAfOJHfTqplkTbFXSlm4ZR2
ZWXsIMFKn6Yoh9GGIxn5RXSJWoW6Aie7X1W01t6ll4vI+IdYAphFqI/4eQdiVZAK
YNOSUOljzDalOkH13XlpJelzaScs1iEUehcvkIkBDyjdjFQeBSYDTkubYFrODRLt
8i6/lHqQZwxKptGc3exmoQS/AqlL30wo/ATbh2klandtPBYYP00QCp4O4M9tiZuv
2CGF+w9lgbGT8nNm0D6V4XAfr4FgBK0XfBZc7Ff4WWoJpDn5V3PUsK5eieh6bS+u
GdlvWKnziPg49xFAeqoU6vZiZUuJuRELvojrhLhs/sUqY31KslY+WhybOE+eFo17
fiFj8U3FdmPOTFWnsZweIxB55UudxcOLY65/S+RQJxwxgXDKShQ8EHIiRNsiCFyz
jRLJ8zMR6O1ZC6pLxsz/rpmKr73j3s1u3zbdCYAEwQMnajZpJXMLICvJ7bEiMM+q
QLY4ZF8Fii4lDJ1h1MkTaqBlsv0e1NPsi05z6foTNdnoQm+8iNSabj1XiI5Yj1aq
nKLamUQbKgMAd4QkZ4pJEYVN2S1K0DWjuYcvQl6StIpz+NGUQqA+i82q8VyhWRxF
YihjnnIuMkw22aA5In5n/M6DDNNounb5NVecqqNR7Jmpm8ksNl6d7WipxIUmHNsM
m2R09XFEeXKxxJ0TIkat0HZW4VnIrYC5nv7tcGlYrRoaK3U0UtX9eeowfdEfT60P
J2R5P1hYtxVUQhcs8M+PCLEy/kjYdz9K/3VDPjP6fRtXI9JfssL+HF711+0/7gTg
rA0Puxq6VRgf5huhX9HXRIC9fJ7l0T3zFhukjncnkabXvBjNyaahtDwk8C3SBWbH
Q7243gDYUpBBRzKMrBR4yvODy6nyujTNQovJN9p6Qoos01aYaeEAhEsnSMrMt2Tw
uPvwFBQUmMcStOvZU3FJuJXNfH21tHJkdUj9gZA2BrhrPHX5dG8AMBRcVc6qEjls
EoPnwP6884qs3Ur8RctLxq9Q4LWUjW5jcjR3lvNRt99R0XVcZJiYWFwbagcgwuaL
npWi4QuzkZMor19C/1muoS0HOdwECYLUgm9coi1i29RWMcqwG2Vy3qxCtOuypEis
J6pb0I5JhRlEJ7qesyBepPGuRMWFh9KHbco646C9SSOL2wuOgRqVEaUdR/bvRIli
Ly6XJ/VIcH98f/CxBYGVM2IoG+Av02gmg93i0gGZc+cl8cH0/72jfgjX0+QZXbTS
h7mRKcXhVF7Lc9XSCMjW1r4AJym52HzIxzR6XZ2ZA76RsXF4ISs2/vOK0W5L2/FA
8ZS1HZovh46E4r43c+3mCGRqNUG5IF7+VEJEgs4ual7kHT0zEDeBoW5EFjAaINgK
d2tkgxNhtmOqJYdUwbM542TvHeKBdNBa4XJUFI9GxjcXbZVMjanvHMqRZE+pLN7r
u6W397vdCX+FbHI4aTHUAEqU41t5ukoldJJNk0RMy6IGl9PIuO6baoriVlKU+Ddh
WttIU0orJwJLmd1eb/zEVQsMs7rb7AgjQYIyS/VkYwkgpDdIUsntOQ8S37BeQvl3
tELpmX2N+mSoTZMSQIv2l0z8UhTLWINViwsXkVHO3jdI5KmJkW6i9QEal2cpYiw/
YR4cEovZaDh35AER4mHDGExd30Jbl2ERNErHbypD8STVhaKvWXIX6oSnUhlkaGUn
MPaAvYxKqFaokfOM11IhXqQ6kGSFUoOtVu0WAUcHvKMHD0hXvFQYq1gt3frdUQt3
YuY7ZdWk/1XtJhtmE9iAooXQMTG+4/xTJ8vLI/GdLUg2PwMUWB54rl/S7MhRMI4S
mc0FjMWN3GXwGsWmjwJQdYWwpgP9TuR7IvsNGzHYxVG1CMoZ1DagJ1qQPooCnRop
VaMTFtHtS+QOGPoiqa7ZGmvRuXy3KAQuzmwirQIYPB7YjJkQtYS62+e41GlERb6M
SBZv2s3NsapR1xZbRL/xDaMjsgo/0109NU+QnxiHo2+JsxYr5XAB/C7G15+OW+Wy
/2jKv1CaikdOqqVBVDi4EZc23I0mjTR/pUfuvVZCx3ButOrQLppeEo0VhqxHLwEp
tS51Ri7rJFNrvRfw+UAi4IOWKx0+fV2bPoDkWFxwX6KyISJBHr4qu+8FhWfmS/Wu
POwAaobky2y9A8IqBpWKQgBt+JNqvzfP8Ce11nUgZ3QPxMWa928us2128ID07TND
1dWl1rib1g8JTynuAtSP5Oa75sEHqRGhDLx0hSY9U2W3oS84IDu47u0wA/VhGKxH
FqI4Z52N3qlLLI9b1OHL8lFda/2pfp7hP8UxMQPiIsyEKQsKlGQDzD5XDXsMzIBB
s0TlspwFvpM8/XrXgOAYLYuipNFCrUFVLrSs1vE9FJF7SYGeYLNMCmzVu4wREIWj
Nr8m+4eSTLiiugaJRJSduL5P7aQVYQJv+m39n0Th3j7jD7Zc9AoqZRu8wsHhv/fC
kbM8W3Cj45QAKEyDvXCTcKDBuMwMWag4DFl6FLOJRgfHtZVYNvMShj+OKgm1WMxS
oP+3Eji2zNxxKYY9hwKj48hYv8rriCmeAk5iPSa43rEjGkqUIjDfo50LHU9gWsiP
4RPbnSoAgBQpvUG52QpL4WJjPJlzQPae5R7941a70rWaas3Pgpp9EkK+5TDmRB1O
KIQUqKyByDKQb1RH8JKSHNZU2bka6bb54QIXdj8gwYAAhAQGN4dWvu0yHtwELiP5
L9qNzGJlbXpODCvgCag4652pnDCFiNfA6XWnrMkcZuYzz98mE6WA4AStTbeeFW4a
+TTIOs58JkUcB12bRF5CWclCyrK7dGI5I3g14b2t90rpCyg/jE8v8CPQlkPNj7CE
TbFuszNEGBC0AVBlvwRsGVlOuhOFTD6T26gAq3yHSoh8ipjiUSA3Sc+XfmvoDYT8
rMBPJXcs+B/t7tofWEEQchpSu3C5nf60cwfyMHAtOJGhgGey7WJLL7ILBwKzxfUP
k+nwZAFXIjvWfaTOYcmrsgFjORoPvIJMRTkf3ybN4zv47VieK0/VPtMA7UC3Y8Fc
6drX0KYY3/P6i0TN0hNx8Ima1yyIMLEPyk6T86R3taeGTrVFAIbkPLhwHnWQ/NEe
bJ7dX8dmb8ib0O4mxRJt0yN2pWAdGjs3RGH3OgpyNmL4YlcO0jdaFt7t+SGoNd3J
Jwc7wEuy3fSNKJbZKjXBUSch7KCpYazBtHDttCGaw4Z23FneobB3GWPODczpTryj
37R3v/3KIGwgR5kcSUU2inPRejrBETXVZRHLYpzIAUD+WHNsd6nRzQtTDtowDttH
4anqHbnzHllE2T/dyFUpOSyx+9ryY6+av+iUDGa6RuVKLBo2m2phAnRQytfhlJ+J
/ZA1Vn8PB5mvb5qMGkz1ejV9/E6qn4L25b9IaJiOyNHtx2GYQ8cc+L1+w3aujKG9
mD9rt8Igh6QLle/+OmcqfxWcJb80lIJUc3aLEu+4stOSQp4B98lf6iXTa0VsS5ZR
zV1tjLh+ATR29DRdwygV8Cnv8e8QzM/MdttzTlEDTy4e4QTNh630Pe0BhAmCGG8P
7ndGsTwspXe16m1t/8Aw4/8MQcWT+UexoZV8mtdVHp5rjob0s8bGsTaJj1EFJgXr
l6/qvvFYG14I0Nwge0zj09GguhH4xICk+oLpv9d6y92PaWZwhtalLP7zk2LVMJqW
+zox+U+kZvwib0UIKqcF3cCQ8kiwFBzXiOtumSAxy6IQeZ9zDpKeI9Il5J/LkZzc
xgCvMuB9Rf0JGMSM89yOVtjUhP1YPN4OjNLSJGrXwFzoEC5pNze4qBW5uyJAkkgk
ordBdyiQbu0//cLSX9zmGAJXZ/DavqK9JtS3xvGgCAUjss9GsnA9GVh0T+qTtTFn
UHCzEiM9V78gVijSuPRCxBfoIgA5HeoXxKawrp3mgZyvL/ob3JZCxqJMQd6Q/qw/
+n2YpIE54+BB+PRZsKRtxdsOlcDjJtvsE2cFdyL1LXZxgV8oIxD/U99Orh0FAjdi
P9Ga/xf7cCvGYnO7vHHnvNL+LysPzwUbE17RWBPr9SwxVznK4LwZlk/tA61yX7fT
GsNlwJmRP6qWXahTkLVI9MtWJC3idFWpvQWrtecdL2ER8dIkAWQMCl+IHrb7rE41
iP5m9mPo13dCkIGUx9Uegzsh4t4t96NBac2gMZU2reGpKbsRV+4EJs4M0ejG/6hJ
uVdBIg1FvtdQwEvN58WaI44Tuoc75gxrRx/U6jg5gisonk4Hyrm2ctoNkmIFdhRx
R4gXUI9bczJt0OmzubIZz+lsnjTAHhTNCNdjCCMn8xz4Gh19fm/N8KCANZpsLKFJ
RKDoDK1tZpOVUtNmxpvMO+D1/wiK/LQvTb8MXvsY1mtl757a70bvZburHy24Nj6l
OyucR48XevKxIoaxZaShg/Cd2F3OwfdJKIQ05iDETEtLLiPFGbaKMfQ+y7A58Qt6
5RmpSdfhg2p36N7n/r1bpsdBHNvnyaUuAvy2jqYOEeEa38q+3Cy3DZDMkqyA7Oo0
V4GmVao3Le0nKOaL53XhN2OfkSuUEtWJt3WWQKRvPjAm7DJKPBhFCcYnZr5QdXG7
TG7eyhIrSy/ITk6knqlETEthc2jwHkRyu7JgNStXEmo6qj20XaEaYJrHOI/TkmVB
Ek/zRLZFXf3hU6wHtgeRr0HQgiYsE5iv1skum7EbzPVVGkWbMqtTGu/LrByC2uP8
C3N9LuSu0APrPm6VmspAiSHpax5x1ChmdIwiRewukZddGFRLzpC3BKgdFChgO3so
IaRaXmkanYJAVzgsOnQUw1fq1fko+5tQ1tUg6lZcVtGaE33hkQagmCv/QzPPRMKu
5BkEJjKIsxSJuTtvVQAoJ9QzBrJ9bpBpSp1fOiDjh3CUfGs9q+QS1k2pJhEOyKEF
8NtSm8jwS/QXxUjFiHJkzwo1KxEEpC0XPe2dfXvn3Lu6/UjeLxHtjwcNpODwGpA5
zmq2xVQUlTvvuodC7h0Yu5DThGdUaUsoPruBE4AMsy4b9TxFk0eo28Ym4RuQnXTV
tFenqaJUab/B564jD4utQkArmqAUn6lLxOY610aoKm6n/X7jYXFvuoFVXXDd42TU
syP1nTcLiadj0pD2C46aCIcYYwWmb0ewuyAKk1MsmaK3VMi2BUlXQIUEIo99yv8O
J4LSGTyNWsc5n5L3cgf3pYxQfrrp89RQtpLtDNt1xN5Lb9Fjkrbe6fGg5kG7a8cB
qIqWTzcr7G7X/HuEEcTWqlMHAIIueU70EhJB9LvtSqmNoqpkRh7kcFSq8cY0YaZy
FG8E1ERhGyW5P+3GaQGe6Kk9T5MEeWzY87UATdZIeglzCZ94lcFeu3LzTaQ6J0Cn
bLrtJgr7Irhog54qSqAIs3ON42d2h8tpfRyzlQHFk70yiwmDP2s1n6efvEwYUgHX
pkdFVdNCjXUmlnZtESRV8Ja4LFMe5u9EkTWqpf2BBjZsVceI9UiliHt3/jN70ZHx
fK2km1o4FxtnYrG4J8m0q2uStSFKtDDc74eeDvM0AGzAXj1ZhVzQ4leKzn7vm3sb
idRMjIQs33jHB5+jOEdDKTHWQwK9tVk1oah4VbMt9XrFG1x+zIFahZF6906eDfXX
wDdeV9e5j2GvlDICffssg1pLZEEJ94aBSGz04V7qdYjCW67K+cLwPykyUTtE9Jwa
nFua+NcCFebFgfkvB7gxwoPKpxBO5MXKN4gLjR8CutnuT2ACV0OP33wvDfdv0BWd
DlMvGKFLfugCerQI/Pt3XkIu5yiafPu1a9W+yIYrykEUiveKZi9Qky5POOkqwezj
uCjktFE7ICpliIkvMmjcPqk3TigpZSUgkZn+2P6wM5+i90HvMHCRGgOIy/1Rqum0
/aL7kw+ipbXsoIZaGUQHNsI5XqgSrppP2Aq2OFbTIIunSPhUhfh4FCgGIXOYEaev
zY8x95Pn1d2iWH4UnfTXkjsdr5u7BWTK0f+wDQzAc7dxkLSIK59tLnl31Sxr4Njb
N3WX5/jX6eqzQkQrpM71y+Bzf0lqHQQxcTn59nYeu8fuCF9kbaLn5mqNC1X6OScf
HFnJ24OvtCq885z+Lc6xdpro9FC0UZaQ6Hiv9oeCSa3i+HJzlBTgSVSu0tDCNGMv
QCo4WTObyiI3iK8WzdE1hTZPrfm3KzLMN/UhPnJlGHLfujjW8aiorJzrYqr0mQ0Q
cTJcsb+xgrAlkZ2l/vDz+ezz2kncdxnZrGWuAtVngix38WyKozlSxJFQG/8+3afY
7z2s/53L2Jy4M9fruey7pYofBXToETSjopjzInQnQ8Ma+ulV1dxnp2XS2DMywx1o
h6evzDmWSYfPmv1k2FNlQqx9TLlRA941bK+5gyLwuJVxkAGtVY5mRmwiyedX6nFy
oy84sFw1b8ZX97eeBX7AlJxN2Fbw04RSnUgTPoHLClrMZ3vnt4QU6FAomu8hGfHC
b82U9FA0cJyZKTCmA3qois9g7gDZJFs66IfYapn5pDU2q6qxNYWMT8BJtl/a/b+e
6Tmviq6qrVx4HqcrL+fgr+ao3GF5g+1bUV5/sqJDEg98W/t1PNmDYL82MzuDWcX+
7f/B4vi7lL9yv9UTqD4Vyuds70fDo6v/PgcCmRRJ//e1HIHXA35rqW9J7hvSK7rn
MCOkfaOdfC/HNcHr6zpu5EExxbKa9wO5PN7UbMmEVqQPgQzoHBgXF5O8u40G++8W
Jqxi80GKLEOG9oj5CnCx7GpH0QxTz2V+E2I4Bhc/QteYfrwU2DBXWNzBqPu43cyA
XDHJ8ysQiUXsv/aSIQRe9DEaxUxxtzbKvZDRuUfDVz2u4kxcpfgEuoTlDaPJKVPS
p6zKee/VowG3rH/TAy/DDeie7zIMovPtTzVAwpabRuNu+brQJPmh3yEiU+oxWKMp
AnYqJGK7j1LTptXGIsegntrs2gcX+gSwypHbFB73rMWVRGWjTp5j5UTV7Loiw1/W
gRUSYPNO/uX1tRe3H4Wjouv+pI0I8FR768d3Z/vR7c/WZzHcCTKkkLbn3UkGfPYC
c18FVo7Gu7a5zokmmulEqMDj4cS1C3qCFwxesAYD4GYHiiis3jrnrLjiAFoyDSHH
wNmJoI9TqSPhzaWH+vSS/fy2+RozOvegnuqERgLK2Tf6Sx9ynbKkqvAvLrQjlo5T
Eaqm8EAeRMN6eJjGqo4s+ZhcYEoSZr+y+x5fTtB14JGYEHyGJ+6GjWgveKZSDDst
gRohM5aFApSnbto3bevU7VDbT/Ov2qHgE58CuVWu1bwacxuexlXj15gfRZJI1En1
pVeQ7kn6qxomzqrKkiZz2b/5PFfjh6XsQcst186obGUto8TL9AOfMchklXxKdx2l
8l7xHRHZFS8hg8MkFPNd6qJ5pa5IU9nXOzDq5D/ibv/wsDmTb3bXEgTXz/Ai9pIv
beCgsEhQ+fc/DTLYjcLOJhlQc88Rxhg9jYOv92jqQPH41Atlhv0/ZQKJOUgFVG8F
XytTMLXRSOskFY9O/l+7sVzcsPeIbanxAa7STzPzaXg65QgmMSnrC29VOaNLMtIt
tmYGJILGZ76fOuQHrAyjvz6LBGlfq5rRCagK267NttCshO9Ue0ICGD2iQu0oUGrT
+QUrT18a8kyHWFj/Ws9fu5ct11yQHcshce7YIjt2064gSqFBMcUTZe9uWjF6rx96
TInVtPiLih2zJtXRD59CXay0opli1MU3adoaOzS/pSYEVL1uC0BYfYf970uOwFoc
fenSdqepbdfrJMjgZ+faueREwY/ihtq2HPuej10V5hAs9I/5g8hEw/cRMYDjdRmI
QzQoqG1/lR6uWccUyujfzWeeq3khiB+/cMsv5f2OuHxCW3AclRWs5sCwHpc3/qfT
1FHTaT2OLH/rsgCqYHxIvp2rQCTgVPSQUOYgsiJTRPAJYcjAHQ5GOCjMQyqkBWkO
0C5TLFqZUsrzrNW14YAoO9nkcbhGGy/uKNMYvSqukenl/96NVrLD1DNl1FcWWeF7
Z8YiXH9RqyTbymF8llQxJ3hvxQgDPwYRDJWum/Hr0DQRSPmiKw4nCrsaVUCfi6ES
uInLh2QfKF2WzKeFYG6rbMKUx5+rih/9Lv3DbrSRO/e8KBqPjDmauRRHfkh3tzpo
Nvvp1YyK18KNACwTrkyeBQSeaA1ueAfZdckXxafjJpeBgQuJ7Z/0vAOcGq3AZsfm
vJH/hsb8vm3wbxg3dJhObAVvpnq3LyZ/LsBpyjYRB5UXiXqGg4NGW1l+TKcPxkhW
1qTaMsFc5/l0hAs9wXwUIky7tjHhv4qLa9vasI7Ip0vzi9O9kxqsUMXNA2wss8N2
pU3eXEPg1rxzJgGeEUqjx0MHkZp6flzxpm/8YLJjah3bAUUqOlzTuqxC3MeDLfNc
o7s28EO9ZH3O3bR+0kvUAnDtccZ3cjEGzxpDmOkpzt24g6Ki2l5rJ5de02TCZuBM
yF5HWlGznQ07KuBBt1GAPJjOo/4C0W9rqaVgam0ePMJvMLOdapAscE9yLFdGaYh9
8MZLPkDxxzlYcoxr1CkYAsMCVEHXLmayk0k/vLaRmKbIzUT708DDQC6aClpc3J2Z
lif17kYgcseOaXIMEVEsnd0T95RhY5CNiJboY/hRyztgNRFRZii0UCnNIOxI1hlA
ZPhSCePOTUIwWmLjLg7lvTLlslP9KItDFTaouaf8XaR11xPdprU8YALbVQBRmuNC
dqDEk5sdf8g0o57n716A/WM43YIyX9cQ00Z6GkosSsrSqhunGajV5HRfScPryW4m
oD4Ba4d6/4eh3NNbcCm5OETmbQTrqvgk4jVAFioyHvXGtVRWmSJKKFZwMYeZCDfG
SbYe7WMHJAX9l0yYdGPgTtfD3Vy0YZH0qSAV7ZRkDJtYUQBwPn0cVbMESNSRMCrt
WZ7n32HUstxiNSoGIstMd5M6uAFx/R0qvqrYAhhFzKfyK8N9gs1EMp26UAqgKDJH
CGIeDfvVxIAeCni5rqKV+4bwYqsJrsw/LoX0wxaXUtbfDAiH0hi+t89PyMadYpvr
UHb0pIQ5II0V1f7nWW6CjKhSH6mK0PvX9ohTaKtjfpgNZvczGFnQZBB/g08R2FCh
xAFD+VH44PT5dURJQ5VzW7+CSfKKUz1oFa0RupmciRcHjEf9y1zD19fFjcDk9EVa
veSubwMT8vHeT/J6Y2RHuhvTO1WSzlyhLSPPCBzd759K58gZI0ZQ49C4x92vhh7z
V0NaLtKtuTQyLQGVTlptOj5CUzE9HKNKQJZrXg7TovyAayXoiczEEvt9mAmwR07z
GRv2DyFARAsSzCmFxsn94UCg1I9MifuUGyM/roj3wwbmkbU03JVjcC7vwq+47AnS
+Ny+wCuwDhIH+rgzZnztRY50iBP1UO+1DqIl3WIPy/EzOm4/hgIZYp8gW/42wOUE
w/xHMds2m38rhjpY3CYMWJz+WsPAQY1Or47v6WmkErjoQ8Vr3q/1JAbVIudQ6ZBE
E335fo1rGzqmdWuyd/U+NmR9O78qD+gvUbWbH/jecjsMayBYlD/LdI/Y7fpcdM6Q
vrKwLz58Owbh8ccCDwHO15ul/f6iXWUwR8YT1SMcZnd1SeIRvZjc8CAmTc1La4xw
/P4MNPHtX8vFvZh5o1oVl0W4kEkWSquNLHEMqwbdzpP48AmbYA6sLpAM4pfNbj05
sACq2pKl8Vr6NZMVXuBDV76pn2QDWWhC6Sw5lcoqxk+5W5TDiAVEHKiZY84c8dyT
+DNQ2vIQqLPvlfZi/mfqsPptcGub2zpZrblJJBVpd0XzBIaUxM99e2qRfdLYOzbE
VVzdAHXacWVDWE/4qEcabgPvSOHaE7NtL/ddUmPWhLfMVQAgZDqMDjucKKk1B+B6
qqvxBAr3Vcy0sPJvygF1wDLCzNoYYqKihpK1zFd8mTcUS3k8T3zP2PJgVGkoV+lJ
SapGgADDaP0arru9MpsWUcJQ0L0ThrbxgmnxabFEHG53VorqU852Ka45qoM1rYVl
GrC/KyjoKykBZOQ26L+R9dRSlprCswIusbAIPzveLMwuxD57BFDSnzbTlEwanLR5
yN0xIKP72A0PGdZFou2vck7oRmOSX5+YS5olPMmknQ3qqDr6r4H3jUdKrJE9iNGf
YiLtlKR+eM5ZDAZMkKEmCEglVCEDmX6GI04NXMUVmS0C85PlOVrymXWvs1w+yjix
NKZe5GrNahJ+ywxTP61QV31e7MZcgGJQH035LH+0YEJHrtI0xM7LPdKw2mNfAIrW
xbbP9kS9r8E9VHHkgj/ffNnKmgGRPylZEnoCfEURdZjPsfkDx77kM0dXXHv2NME3
qh34mSc89HB2Ycw5h5QcZvrHWWAizST0XKD+i07Ew6Jn1ofv7ZbQ9LpfVIUeHSVH
h75zDMQPX6TmcyiOnj6wh5+R5GpuQxDK6Xo7yNAdV3sAd+JFqqi1v3jHMC+YFc5Y
KR+r779g/QNriBNl8JjZ460nagA30l/IlXjqXNbCZoDEXNq1wr6hmdu+Z+rAwCLc
aB2092OieWrtjMg/N8XIxrxWS69l/+pVq4FkUgYdq6Diez28tjJWpDt7fxsWiihA
+bkJgNJF4siBTWRMTiYkYWKb7abyO9wbt4WX+KXBcn6BVLxzYWhCYPd6jZlktVZG
Es25qlLw6eHxiY3Gv/QTl3wP0MvtprQ1wo8SQFxY/ipF9UcqVe0Etx5T+HkgC/wM
evZvvmNvsgiuINuol/mix907mACBejnHtg3coZgTaSG9mfMVbAWZ/+EElpNfpHV+
xMtjbyGWQ+1NqDrZ61CZdFal1e5+zADQMJpRjssGvjY14O8nuTW2hsNJKvesdUdU
4Ml7Y3vNoIEzjem59QJR+yS+F9zdlE34lhKK4Le7Yknf78CQfYkx3kjHEHyPvE3C
vMPFQr+71sy61qKG2IFP3O4I0eJWQFI2PIrJsS46m9MnCFVC/lW+3FASsdiQCdQq
rt36ijfaYeppA8YlcD2WQ/VJ01ulX0TcMDZFH16qsjOsMwG9Z1z9Rq+ybsytwmAN
hp1Op0eP24YgYYfl4uOW9Ow2BbQS4Al0uTiw3HfowMPK46aAlejUgSVXCxRR08hK
RO8+V20HKZYN6bjnNPTjcTuJbwYbKpYY0Dtr11a1ns+7kl09Rmwjl182hlYnuCK9
Kv0GemDRzDw6t+X8eeeW4YCWUOswwdFvKuz2fAROBSzUvkrx7DezC8nUJ2AnkFUk
w3vFbAntjFcCVMHUp99eUu41wL8OLeAXzy/bDPK+C+PMRFW49kGtYtul4SRuCOMT
8XtrklMVkZ0ypf8mPY+k+MJw7oWNE/Ls70XqmXgf0CyXXBZCaq5KR5lHT0RfcXus
/jy2gaxRMdUrO6gKB0B0DrnhQwP3oPYAa2RPGV7XZBfg1U9sIzOQ61S1oibsQ86Z
YhlfTBVXo9eqSLivON+p33jFC0haPIgFow4g9ft6oofaqjORUa9E867/6oBsM5au
n6kMyFnAlJ+ZoJFI/0XhH6Qzs5eqoGiruuE1HJlhFMbYv/CjdwOQlWxPAhA2rhsX
Wzfo4PcZViWTE4dDMWwtCinO8GfBdAHaClVOWkbUt+wm2oz03dn2WnsCl/dtioK4
rqZlfxZU0ryj/u6BYswDEhzI/2cB/eAkgnmnF6iigrZcB2quEEjtQI78MXfOZMcY
xXZm/dU43Nxld5yWZhJXI8KWvGir+DqV0QM9dlkCSZ2wtLH8S6okhaCSb0xRylco
HyBpKJZNVZn4tN8wXVnlyybLrzPRNS2+AREtYm7zD7J5MhS1CwDzWlIE0JJC12kx
1up1kDvrHFBOK4rYwLN+DTIFI2tXAqHNMGOavSA4RC8oxmoq6iv4FT7RYBq3UvRm
ehh6+6LcuY6L3l1FFY9/gzbHWH5XimVNl+28r5Ndhz90v3SRwGBP0jLkpcuJA72j
MDJlm9oW9n1NOCaAegN3JzU8YuIDt5F9/dDpeMSeycRUNGuXGjKrJjom8iaKi0gj
TUqlvmLZ14xtb5wxlWBJ0X9s0JeM+QicHuYkABacsClpc9Mq9bwBBYf+d5J8jZb6
5jVWyb5xBgdp7t1xQY151A0ZLzeUN7PjencL5j4B4bjTy4UwIYQD1hPDCgwpvm18
tRGGv7AWsUw8T2bIOyZcP5hn9fqIy+TwJ1cfoHSziuMSTpGg3IzNZ0gxPICPaSLo
bNWC7p038St5axiGscxCzOUQGswz5l/ZQ7lAVXJxwl4CvnWDdY2VtLkDWdCEbV1g
/vh/lL8QZF8yjqF8bKK4EF1IaCBU31FCoI9UxiMt/6jaalrXiI+rRPP3m9xqUTer
gCs7WZkDZQF4bWuhfI767oVn60c7Zk/klwtsKhPGhbesxyvkkYzdIYlBi3sN3pzw
5RSsJHEN4pPOgGfJ8vU2idaOn6Rgj82sjUR2b2ra9/5IIOgVohhNGkQSZGaUS2Rs
iroO2iyKjA1n0GmwZJffkaKqAOOX7eH/OJkGCc1JamKSXVArs3C40BQaXhG4uxdg
AMJwV4f2zfjSzmUXR9lR8j9pCmdT5INqo7BEHQWc/N4IALUEmdAxR7nSB3xS5/30
rrEXeqLLxlocX8LjrMFZQYCGzxca91oPJfHbDDqRkmgyTh7WqzIuEXQdwSAkkVai
A2y2YowChn9R9utAXJ1QmKaUtj7Z3CGrmM2I/bqxFgN800fY8lshHmKUBbu0Md8I
4B+LkpXAEbDDk/7n9pbRNWgF5FiE/ReaYDgVrlY4BHTE7DEgiijYWZ4JZm6D/2CH
6zfjRrHJwJTQwp7faw/uYGXh6h3fjkUIaw4V2VVtWcVlJlqijWbFLtbaKvlRbJGz
h8UIXiGvsFEolDAWegjeKR/eSkS3V0/i7fMB1OrY3bJZr0jzABpz4HD+gEacp8Qs
Dc0INav+kygEeEUXe6j28/uYgunVBZd0UV9lEi1YDBm1p3rKMPr51OGQgnjHyKGp
jKNinRoPTgVFv/K3fr8vb22llE52GlGUS115+atqesvPgkiyc18tQhcJ3uQNoOzU
g6G8/hhPVnnIdoeAaZzUxaOrTv1QthsBAdsXLPWgHVzzSO0K+bqx+UZNIYZYG7iD
49ML17Ej83EGZI5dDem0vM+oXGik4GcjyQthxjtOKjplQ7mbjMhBWOzrjkwjiy0m
I4r2r1knGnfZaF+x/syRIOvvI+1+XpoaWJicWw47N8QxsnJOCdN0HuANPI3oFuXv
5J/Dznxm+pGzlhmZM55GrMeQj9Ukff9XcqfGuIZRYw+vtLrPNVkd2nn4BYkQZBM+
CmDGGf70jaS3CJKLeHuR3wOfB4d3ha4AZgL6o1VfmbkXTBCHEeFpyZkK2F0s0u9D
9AAzkjupxqL0joHlJ5PU6gSduDyN7Io7AukU4sgPtZ6BH2Jog/OpdaKSf5TVKThF
X1QXCZsQhjrHzImf8OuQ46UfoY1EiOX0g6knCrG56qJG20tVWbsFKhMOHwiFV1iN
ImkXywhtZOgZ1CL8prnyZQM7uq4GC11UtDVo/KuKRvQaGLnf7Aq5nP1zKT8aJ+HV
96fSylAb729SP+zBdLKsdC6MMJ/u3BYtvhQY7+2FEF6SljFCD2ArFXDBNGXJn+G0
cj2SA1SC8bL0pLSNuJheINw0EoJp0GJYbozX8SXMaSADcJVu/t5qPnk400OwIHEn
x/LUSHsy7YaVkFDnOERWejiuAeqj9Ii64goFf099awQmn58B15/ujXdGN0LiYk1i
AHwiHJvyHYjDfNYZTrtmWfuBxF7ZQ0EzK2C88khN70wbrOfjrFwZXJLK4679hY28
hzO6eAdmwWtxyYA+axpMxnCy+hr6LHJVTa+KR3KGZPD2fRmAgRYNMBtIC2dz0S+q
vjnYIFeY2f/EEviDw3DoZSIQc2Acpp72b7AvL0+Iz1iqq6BWy8U76w23/9gRtgkJ
YrPI3p73l8yfDtYv16i+jBkn853PK9QCzqpp7Mgd/fZCWhs/bZPNKSu84NNhByS1
hnF1vEpihqr4T1I6jn82tzyolUbfws+3h72B6oVnbXK+t7bZpL0Nou3iji+FoZGN
sIJOJ6zdFBd+THfaeAfzJOwBaq1hd/+0MrEc9c7OOqrMtChYKlA32zs0GhbviB5z
k8wThDzE7WVcu97Iym/PJ65W1fj0EG32EYoNjK4xDXMHL1hMt9oJ0mikEt04pj5r
S5TglN8WXLNrLmTsID3aD9RIHmi2Jb2Qpvl1JxRI2WPa4KLuAzZ6ofOzMGhFpD4D
OP5YfmsUqKjnsdYjv7N710lGU7CECWR+8isOZRVbD2Q/Bi1x0YdhsNebIXth7Dl5
qF92iUXYO8CK7Odke/gxUPW5UTpPjk5KiXggRjL5ZvBeOwUDM4XJy4Vs/uGQDkMS
w+ZgQSzkxmgXRzxMoeFuNNQsLp6uDZKlFln1mh8VsXdrw7SVCkkjNHAZt7b4c+6W
wbIinJFUU5R4uuPKMyb0BOyULM9bjh+pE1CE1S2mDtuBiV341N4kBDCg3h90HIyU
Xh94TNs08ORV7zqZkgd4mEq68F7NN1QHjTeu2Vo6jO7CGpUL3Oq4QiuvYosYutpv
1oYcB4rASE7t1l+M/0BvIklsvqTmytkGL1PYfn465+C+U1nEuoGQllV9pY+pLPK7
Q4UpVbsq2BBZMIBFU9v5vXnmuKca7FbgDkoEAzMo8wSp1aWbCOhfucrpJYZTA5PJ
0JIeYm3P8yFJYsokwvKASgfbjMqmumkiztRCYzcBjJrKFSgdcfq4ybQh26VCgPoI
jrD+x/6npdlBq3DMTdo9frRr8AqYiYd/pf+sjAFaDu51uvXrucVjIU23mJ6PUjgM
ZQK7U/9eBQjw3lamC7lyxDbVeO4uM3NtA2MYultjeNRsk9lE+wACeCuKbKGSCmu4
niMhs45kyMrylBshGrPzxyI7SpniqC3ml7e7Mcn5rozKd6N4s6K9Y60BVuBALiG8
Wzqjkh0B3HBwUF9kuxxiFuyB01/gLfhBjtjwP0IVA22GlEGI7Vy7lkzgcmmon5vp
jHKAAvGMUR1OSA8+MQ7WLGyQoVl/mqKr5d/WZSb00M4L82H/RqkfqdbPEChkgPCt
zI4vn7P1XSkKw/rAqTTkAIif5+HcCjTmei+NPRCaV2FK6eoXIncievJV8h3ewVdx
FXlHpxaRpq42QsBCjoBoRSU2pUHNTCruzKCQ0YrdTZ5gixNb1nWB+U5Kp76/HTNP
GtIWnazMNkIImL6TVHVs2J0uMeQennqpDzTM0sdOqdXWUCkYvuYIJIFnNZQAAiDZ
gAsL6p1N/gh5Xe2Q70b6ZnFv/3Q7APftyRWExPgRdv/wA8uoFejk70zPVYd47Tgw
QmZoe/isweXfFCDvGk9tw2gYyJbl3Mb5bvc7rkZyzpU7FEeImtHrwM3ewl600tBM
unixT4jznZHBdPuwJAYEu7wWfIgs0XCocZTj5qD6zIlMm2VEKi8lwwfWTNVVuEJj
yRdGbtH29UECCKQtNhUBWrzvZHQvgkB4sJKMBjBefrCz5reutbrm4LJvUEYqrDAg
rZZB6jfOqtI8gtlfC4TjITLq6XCrI5uDNID3u4Jns4pE5HjiKW+GiBtD9BA86NfM
cYIWPs1ItebiA6tjkFXxgWwEeeFeRYsSjb5DC7KOQEv0IDTBU3FDdCnAYpSX0D2m
Kjr8r10+Se0zgkw2iFt+XMfaEdTzFWUDfLAtZA++Ib8TDPR8D2xB1kppSOlLCZb5
wNSwtpSAMeNfOsJRXIol6IlBs1QD4usKNXx08X8cazBicOOzKke+EYLS8np1Gslr
w5gzwrJthZmhJwrvqYBUoa9aO738/KXDhcIhfhAZJRiJVHf/0yARH2xJH13qOfFN
D9C3m13H+NMxFA4bU4LGEyVy9GNO+Wiy+ES8LzxhVhituJwPDQTRiI63/+K7oaWA
WUaG4wB3l2XzfI6+klnSOuWCojivFjHg2YhDoIOOwGSElBxhBBZ/7WZdg1TVm+7Q
07bGsnIuSSZJ5jF4l7Nn7T0eUmF2Osw/vWIzoBlsQMMdh7p37/VfK0d3JHiufS2/
p1JDSft2Q/0WoKhMrVcrQ22MixKmB+qOnMNEzuQEbYoT4SsNrgVa891Vbt1UjL6W
nDqayxE2xx1Sx9eNgT69chFAiTA62Nyg3C4TIUb0/2NvbI1+/Jix1aN5dV4vha85
mV6PWmUFTWlLoI+WRRCvhBONHPNfGyBTE1l57LUqi2OQdrMj0tSlZIn9PeGCEGNw
n3bAGCHEgxaoS4DX/AIkAwCZSiu4CctQnHRtEESEuNzgWZACpApBRcXjh+zPHq83
ZOeI83w0HZ5mPK27G87KTpkgImJlhP+LhOXBmjivoEK4Hdh7o6w38AnzJ6TYSuP/
oHjIrAh5zUtGzwtF512q53OhP6P+z48bqQ9Nzs1g1H3gFS/jaa89wa7XlL3ccz3c
QUUdLC14OK11sJ1NBrO15gj01x+VkTAvFq5/yz70LqcXSKWYnCJ/MowDWW2TR8ok
zzgzoXTUtQi2/lS+oMGrVpWBIdrl2IrgjYLgbv9JJmN+aNVLmRWNSlOtgGxSSJFO
wSyc8uCgVSQIAIm4C3oVoaG0xDbm1RDRXT6MBVJ2ohayY3ErRF3zsN3PWlxn968A
QeMCSMyYHy5GbvuGpHK2UvT1+PEWYXfVhc6RNoSVs40xqMMHhOgWQ9tvoM8aeutz
NVLnSjhK8gRmfhmKMjYS7upWrU6TkffXhuMNYXm0vaSUvIjVaqPECHxLMb1syZJ2
jnkCJ/CpUyAVIm6HE89SdCtj4/akbSLRsFyz/GLTYORiUk9CTJT34GwN6dOrEloI
j3+ekiX01B5zM9zIcvXWea4WMejxxGPPWICKCDEWslvnp+5cwfyrnJ4rfGsGeVcg
XKtzhpFHD+X7WE77IYq6NTMMnzWaaf/XJ3WrRWzZxs0Bw/uIJrTw8hlTqIU1ci6o
L6xw3NknUGxBEqwEpjI7XPYS8YMRMvKyAogrtHO2HTiqcBIp7CVR7h6c1UYM4NuD
ep+2koiNBO+XQUxqZ3qs08ZcFEPOzDbSbfRSvE0O9jlD4BZWKvIsvwDKqbdYwVA/
djce6lUtS38OtDJds/WL7Kc67P1LqOrFhmXlAiAWheW0XFgr+DQo2pJcy/3uS3m1
AiDWeIrMeey9MtCjv/Za9fAY7jZrb2IaL2xFZ/qYAB2uDnMiqBsJbnJCDyILxej1
y9MU+60qpQMAC4YGEjr9DR3QjYuMYzBFozGhZeT//Cba21wt71+v00J9YyULZ0K5
thNonIi99NpdenthXYxJWd9+nN8CJzb2wOWxr5D9EyjC0BxBSbtnF8WFByB6vDzH
R1wO4d5Swt4XRrcdRpahIuIb2lGtsdX7kggYH0pXv6qWXjQJL+MZAwkaWNLRxcPF
BPuBWWjpO8NSgnU2wVAJUhmNtcLhZUEmckwnh5o6iI8rImM92Q0KEsoSVx3h7eG2
hnpeGaAuxp9KOL2xF04OerpTjaq61W3Fph9pPZ5alESTNOouWkn1o0GlTybVT1QN
h+Wy02sZT4EB52mVybiigYxanNxQ+VALLYn13kn2Ly6oHr7w+VHDBs/zDWVj/RL1
VcgL6yy69c7HQ+g2WWn8yo4RoPZzqmgX53ArdsGtEpihV9Ns8ccb139KzlyE3xWD
LI/1Ba30JVe+cTt+Bf1wr5Ea7znbdM1GSIyo/OzzDhVOJXqgtGu+Tzj0mXqH9HFP
/H5k0Abcxkvi1BUhj1wGJb5+bnMk1TL9PmDU/+rIosDl9WpOflQ8iIuAKCdhH0XZ
MB2Tbnf5j/SS7zvK8bgDmHR2xjQGA67hv8T9N4cO0JtOEIeIyYjVc7vIN4wINPhp
dWPE8fIguGzMjF2EZMTMjmzkCLlxcwH6AwUht2ivrVJ6k9WQC+kJevHBzEg1tnpI
SLHLaaps4/ITnyyvbscsvTZrUEwjTVVd/rAAnLwtpIJRz5ZHKJZb9HXdyHhzlwMv
wOELm6D8xD5Sb0FtQRG5Ftmh+LGhOwSECHUrI1j4MV5vVozmFhmI9lzY67Ye5Ot0
aTFq+mz+cBtYP19/zV9QnwSdadBSMd+oIGtMVlqSFt+2HVSWsm4IbZ6NIl7cHH7l
DEPqzCsqHWzZhJVwgS9FjtozjLN58VXcnZYd6QuSmRfwPJmiaCBolYMOWuYT4Td0
9WPHjhj+xryOB9h96VUii1Jw7M0C1K2tCNR3Eww0IoCoJJaRG1nY6KRFB6eWFZs9
Bf8StMqLWhDEsSZWFgebpnZWQRCAYidR+kLmVn6t9q/Xn7qTWzaWIs66Jm5joL6D
ofY45fx22+YJz8SyIg4MMQQ4Jdc1Q5LZEcW+fEsZggA4xV5J20nahfsDUsFMAJy8
edRnsdO9+Yn5KDSIf7uyM8aoarGRgR1ZUXyiWB7DQQT5D3WEbHd/rbgJaViCEBrx
DihN8m35WJ8zyJf9ggHPltDUbZWjxLgEezMzXMqJ7Ab/Q68b0uNEQ0vM0aWWVSt9
wdBXzzqyEn06Yzo0giVMtFAx3xPrgTJjAXj+SyDbct1Rt5kQ4SaqSbZejhrLtM4T
DFifllLKdFx9ivAhotoJg69nIbkq1Dz+gbcuTrUbzp/FKkOyiTMkalFEJDWgTWCR
DK6NMDuuc6+Bsqvbx+Ew5oPlo/N052DsaEPuGZWq0q/dL3iJjruARZ9zyl9TSkKl
25BQ5duelVBPiLT7SVUQVepZaUE2ipH08ahyGgfc7UXp8wF8jui6+Um2GRJALiS9
UZ815nYquYA9BVkciman3QvtBpWA3I4LQbspd7HTT82LeqXNBrRwHYkIRf6x99aB
ShrVSIPIPOtSAdwTSZkElqjUWxc4kFfu0VQQp6ibLXGB3ZtjY16UgNRToq0whBJ+
nXvOm+8PzdCgCSWnQlOjLihHk33pcO5jsvOW0ZTjmyF+o8dAiCoKkFwZ9JBCDR67
iPOLvYG2SLxFRFSE2dF0aJoMOSbcyupGfNfrlM82ddFG1fXRtDJkiUVXlXNaqzX5
wSwIjIRR0OVuzXQHjFDFx3uWYDcM0HfN6u3boNo5wHk7Gy4smyeqMtBynWOVyea4
wmRmndV9r2C+o6lMxpbk1l7Kp561wsipQslhKHinxxuuGa+HFOYectCN3L/zx10j
yzudc9OkIFFJdPpIT2sHeCasukkTFoRExSCFTU742C9RN4PV2r/2jyYgHehmQ3o7
WLOaPMeZaUjX6Lsy53x1uWl2OWtIjRu4JTyaiXqX+l+bBiY1AZaF7ulel+/rqpuf
vi7MsAbtCM8EqVhR1p8KBNUHizptQO8WHVCJmxKZklgDDoCYXM99+Pl3l1ieYsQl
0rrZKK8eviOqFWOw9sPQINNszSw2VJzRCR3cGSJSiYfdb0ycVmkPzNxk4WD3F138
rBJjud1C45LthMwwbebF//2lKUY5eHaUuIUTr6dBIlNkoMHm5QMJJdnNvCy8f8su
wa9ilbMhBZsCBtPxrMt5xGwqAulaKo2XQHiTwsQQFZEIRS5TRC0+Z/bUVPayrCv/
+jf01NnYEmukXGoMAA92ELNGP834p1LqGTQkweyvEAbRNImRVKBnmo/1zhZNmEpJ
MBdXqMpq6NHlAyoscfZw5DPmuhg/AvRDuwDteHexja8okKJfY51okuc5nqvQI2Bd
MzwZ49Wp0MyejmjwNCP95H7bGJWCgbsHb9pTELPlM3UrHdn35g7vZvwIsYJz7ipV
Q75qvMTj5Jy0QxCqaKfHZ/Uu75BoaaEOEbfplFQBVOE7MeyxFLYWDLf5SE6KlbmR
rhXewe6++tMgObdT8wzErjrLHds/xlqPDHVaXISLxKAEavIn51mSOil/liLO30YI
NATN60koukwZ9yHVsWtXRPon1rd6NQnm14XCRiG02vgF9ha8nFwXViQnDUAn5yEu
AVGVZUyuljP2vFoI2Kw9c4WQLzZtcSAHlMyeCKEXWcRAtNXDeq7zvklVPq4QiFHD
VcGHohhGvdIeh0KjAVQW1Pua1Zna/e2fPOGx6zX9apn0dI2VfAA0f6Vv5tE+W8IN
C4qw9j9E9Y0A0xhPI/cteIvditgx/8Dfm5cGOKKC1jUZ52CftV5HASQmQSkiglE7
ufpv6mCKiJc/pqFmy1O11fpWLsY29fH/88LE133S8nx4gi4rBTYguTUreNdgG/uV
h6JREjfWUn6YMusU9nY32w82h69xlC61PLUmK+yqFVexSlbphbemc6H3JK6CPqPT
aVc+iS+8uHFSAPfxQFZilc6weHzA/AggSgH+Pd0O41yqikt5JMYjIK6j2lu3BFlQ
EKxPBoioLhgYq4AVPyyb1tGixj/9lo+t//KR3v3WW94QX9t/eFKEJ2M2qhKKKmPx
24jjYYhSuun0B9BHaUOObWs2C8XLmqDpPxC9KnSgTQvOCMIWlRJzd6ps5XylLq5N
jJ70Yp3kagkVSntcnY+hUjSU7GCaVoIvfqjxkKixtjJdj0/Gsc6z+OKKcuEbkcLs
P8EzKWqJdv/5XQqk/PniX1ZLcEOZsvBaY6Kwq6IqUNYCOzGhZYutAG25ON+hRoVw
rpeXcLYIv0FmT081T03eEO8Obgp6l8hIC9ABH8EHcl4k+Sk1o7xrPbnaqwAcsaVQ
FDBLJkZcou6aldKOsWuLW/AiLdB616PXHMeKxjYUxzAq4mBZRecwoEVsYQAexJvL
7xiCGZr8KunRT16i1WQOBD9uYo1l2OAHPs66Cnuq2yCBSKbi8j7IvCotFgLTp7Lv
Z289/u3XByaFFfusQ2+ubZfSZjR3wC42cmOEx1zOGsSCcFzB1BWv0cYWWtjiQaNj
JMUG5RtHsSvjkfB8o6jS7Qdh+WuKEyAIIvKRVU9W84l7sMnIB9TlD50g9Z1yNpsL
S8nVJLfQ0+fQk52Ly1cDsp0a5zk/POvpDNMgDW+VWqXj42LF6qLgoYsu6PrrkvnM
r7WyUONeZtR8hFAaLmoCy3QMSmtBJWVxg40iU4TOCd28QcW5KMuZJzfTiIof1dC6
bPyePzC9Ecx/tmUpoWFOFeFhdFja4Jnn9PPmn7ME5OvFmh9JtzrU5NJkZc8G+1NM
ZGk24XMkyljqgeBl8f7ajnNpuDdXN3/qOgT/cY942RzqPLteexITvcZUHMrXTyp0
ytvPNDuAyU/AZzT4dk864q4H0TIIiDG2vXAnsR2TzOG+wG1zfgg3xGxf/xX5Nu37
OoO2aUyu3vmVNfY1BbK90P3bY2aP0Ry3KimTn0l9xCmjHsSW+VQnf7W4/SzbpaCU
3kX6a/gkSleGVGqMJk6CRmMIN7texMw+10wP2a+UJoskwV2OYwAtbjLZXpN2NOk8
P5n9am1QhW+E+/NxWCPVg7+RrimY8W9+bPguWDnTpqTQuXAz/WCCPa4wF/qsHUyj
k3JbHQYZ7QM2l98QXzKuX3hOkO7mctKzqTuyzhRgAsAXUxpg9onxrezsswXTfqnn
y8ptBJYkcMGI2j0TagH3psP18lAu6BlGy//3Th1y3Mr4eA7oZehT8xNkZ9K6jNGO
5Aw7ArEES2yR6tSIIFEsKp38DPCWEk7ifng9aBsAwpWGmFDA03dM7kwCoyZCa058
ZtPbf0/AMkLP7M+Ojq+Z0V5d75YMZil8WvfWW6XiDwPt8M2DMTEgJxXgrNZRAfjj
Dr9O+kfm3eca5FtpT7dx+VP/oD4dpzz0GE9CZ70MAsUsWSB2dnT6Kcuns2DDKiK+
X8gsg4beJbiFxBZgnx1HSE37pvMRVjKWUEAguhcSRYl1bpgMskp2brzXA2hgPlHU
7ZEz8tklnmOVUXiOxZ1IqT6h4vu+W5elszPArLGW57x4ff/USEBgLDWuT3RhlAyE
uvFvIYK8mUSLRLf6tFWiQzLIkFR2nZmoiMPnO/RjsUGkvTTuTv+iQwq2VERAGpbM
Vh7FDg4Uh/zVoUy2YEg5s+U9dQQXLEGcle2Zgziec+DPdgUXmQndk86ObQ6QXxlv
T52sYxv5QKSyrJSI0h+NhiMi9QHlDfawUmQEVFXaaaEyd8g8GtJmp9RaUL/icnkN
JAU4guw0nM/sYiKaoGZxJEwLN+uzTyXNPA2FRM0ZAjYZIQ8LRZsWFqm8AH8Vy7Cj
99TyVle7J4Go96NlfZVD6cL0Ggo9JcuS+e5hsJfXOxkdkya9VQfC/nCGyxVnOV90
r7Ej6VgGNhebqJ1gapAXxYIR1uZvGXBis+81Xf+sL6LHQ9HFLW3qWXavdDApPK68
aZ9B2vkuJkkm0HiMrbwm2nKwB3IkXxJMUACboUm4YhDXZBBtmGHKBQsGYaHiTEPq
yRR6jITPRd9BI9YGXORkGGEgYZCXO4beJQJFrA5IXMbHO9jApoBMWUP7fYD6t/Wm
VNKmExQwdx6sm8FhjwOSawEnsOr4x0s1NbEEA9QJ77nesMH1QfEet9cSeOsLHM7V
j2EzCkvm9AgALRnvirhEBq6vnWQ6CCoRIcY+QAvPc5MCwQg5jC93YObJYyflfrUS
dmfmJ/qWYWDMGQ6H055j9iqUIJ35K7Vv5lv25cgHY8IT1osV1T6uLok5ixIlC0Rm
LWhf9QEk+L4THnzyWeMU8dzoBomkIa3lSwogmMif9iSw60cq7xetFi/U0zwThUsl
ueAJbo1Vpa96zxzxT22rrUNNjMf9a1qcJ1+6vvtF5zFErspnbOXbcn7bCba/V6ij
UPs9s6BPwwPkAagFPE/6XoiOrY6EPDOf0ixsWU1yzAdZ5WGGMIX/yWbBhlritcOl
guEpLSuFEPNp7DhNjDFTls4fMxmMCHQTwTksyea/EqRToAKlgQ6x0VXVyADgVJu2
PaRZ+aFNJJMU2g9ktnW7sq/qZq50HOm+djWf9aIYOQsuhs/HmR49xIznZP/m/WTL
f8sSnaTyMTFNUTUufvIZjMLv9nlj6y09TJYthotbA/uQVPcfwetNBgfTyjTfafUu
oLp8NTaAqjUolTHjR726skX73+P7LLRvVCN6ryV5sLQh7oOuGgWZbomQ6LBDnwBJ
6ws2eIo+mL9EHP98/fTqPSvZQYclOatV3vNgcmHLrR8Qu/IL7ZdvbIskgqsfTn6P
nEYRVemFd5Lrt59JBH0QX7VDCIbH0Tk/63PKluoJEBA4s+2RmHCmIG2lL6lSrwkz
7ON8g1/G8ynEtmkbUEAlbUe/ypWPDg4F8Oppaw58A7ipseIhTq34uS41580dM+QF
OTuvqXbOZ4IbsLhsSd0ByNRtQu0KPVnLAfhqNg1JNGC3CPEKsPYxhG+NEsQMEjHf
5R5DhUGbI6gV44FGh/+mC2I3qHRzCcFuoJbBsea+WR4u4nlMv/QRqqOyfuPW4wWy
5JNmAmRZVLyyaF4bPA4tKYXuZmN3T/OQEoBD5WALEyabW3UQ+DzGY5d2nO6/FHpu
Z6YQ8OLEIo58OpVdeNeaNRIlx/eOFFeeVEGV7kQ00WRzhClUf0wAUVdzmHrUoXzv
VzC5Gh6MW9OCjc0b5vFnOKbmN1u/wn+bag84XNGK7pDrLUakBlg57zt7i7RS/8eO
hUX8bPY+xeDm7vR9kIX7BdbNnlFcReGcVixDO865L5KNZ3BA4kR96Zzl8hvJR2Kd
swYztxnb4cF2LYITkFpl+kf/rsOR6hGjkQ2gpAPtEpE7yF8NtQ68xDD1jIZPsmGw
MBT/6z8uiKrmkcWbjKmRWFzEjhpA3lTBhbOx4ecRsbmipjD2vfTG0TlfafbKut2m
3HE1JceARMrwRXOYD4XG3gMnalq6Arzgs7y0hCVg1vN6NsbY53KOazzaMfiNmQQm
POXPxsl2rcW1a3fyubNZPIta3c8/VPeHfl8hIRd7sfz7hUBK6KWi1Am+fXXmw8jY
OJE7eneRPRbaLkbjQ5C7q5ffzNe3qwx/gn3XvKHHX6KMt9DE0tTX8D4jsnx83/z5
LQ6SBYQlXVjlJNteOhq9Lq4O3W7YOMcUrJNvYOjHQCUbsUVl0F/nIE1sb5PfHiGu
Jrd9NV2tNcJRsLNVqIX1mR2SJ8kqf4f6898vZlKM28E290aMCPcXNvmHvBXQ4LPn
tpnIBG0xPIy8mDxbSCK04KQAVNcYvImMjnoJ1kc8qrbzcZvlR8rLsytWqGTF+1sH
aebRYCoolSCX6PQ/6idH0b0YrMgF0WlBtJ7xxpcuQlw81oBrUjsnGMrtkuaXfB8+
ZhsF3Cm+8SIXK0Xde96/Hxv3Eh1T/lpbPJX5IkX+VMOiOSZOfwS0bGFO19k0szGN
u+5QXWSJa6hPq08NkYOk7IYMOk7GkbYgoXIWXwQ7rCBSGCI9u5zZJcUV+7/a/2Ph
39KB2uxn97wA9NSRoyhcozV/pDzK9c197m3b+VvGyQ1fs3UQ2h4Sc9NWHJkLkDgT
VL7wN625+jwXQdPh1qaQR2U8aN7ZrGBAmW6krIteIzYDy5O6l0GQhNSqEPOIVrbF
Qh3CUU3xDHiUN4AuSXR2O4sAjJqNFzYCCEx4YQagUmv9g85ifykchwIVQ753xE0M
sGBFTYFszFFWxIT2mHn5tW4fh7py/Azm9YoRWBHpfn8aSCBoLuttJMuHMKOrPbSK
qxiwkJTGm/abydSh8i9FY4KK2PNoKofaUtwQm3LApuOgaML0I/WjEVXnfHPJAyaz
JN744v5VM9LYrHppAoBVtyJk2IVK4sGxwDmUkha/8eCsU5UjybfcqDCS0p+DFPOl
DlYhc8zchx0f0csTCotLLFLVwKI4uBTKUBxm8DFS4dQfDkr8uPi0q57opIusB5wy
InX/OHl2x2MIcfTUhA3fv2l9wORG7xvwuWzwpDUrX34fMCB/O4z0yLuZ7pXR+EkB
OwhfxrWEYg/kxLVjnRcmdlQsM+fd0EKMXQNygPtookx2adZyUI/KxcxWcCdt+JCY
fEipcvr5UIs+h+yh26ACVNU5b7tgJcRHqXKAfyFSl0RVG+HYXBWNiQvQyjVjrXIu
o3B0EYY5VrqJgRAcDHHPyHM6izaYMcZrFc0D054sfnFCRm2oVCVEhUSyAw4KAhHV
NPIOB1oC0y4w2oe6T1Bk3pVDvTm33sYBt+b7brjzlT2PwI4gzkFoeS4A+k29TNM4
rHHCpVJCEkhN1sbbIUH7FBXfJVWCbUbzjZR/SVGZ/DgjatqWY/O00fIRsKkoutaX
cMajL2qrC+OWLNUmWHVUkrszJuX3m+QWXgjOiCZVSVxJ1kCo2mC3vpPxN3Mcp/6z
Zay3OaTPVv84Ak4T+AENVumC0/8haKZ88sBsVCLM4Kht4caZVO0YEhjJdiCqzSSx
M/qIpWt1iKryGi3NgKXfhQvqQyB91XJ/VYeGaDI7PJglya2QicLc27caQPgyOk+q
VPeF3NmoE8xGcst2QaO4/yzHwyzFWAEROeba/BVOMg5pIkj5V0hHpaTBigzZp9+L
fhhwwgZgP7gIbMPYQ+C1cvHonkonjgaWBviTd5dUAkmKxATl8co3rGn8WDEAPe3T
jKyLMxRNciqv3CyTgyQ3BdrT1Vk4A+ZNqmoZIUjfrpJ1+JZaK829DNEyHGo0yP2K
kSrurUq6MgIx71GdIHRztq6/VWBtAczTF5/RZRmDXKC8MM+ZHPqvXZhx407luWo0
fH7QvtBoCWZXhxHpWGSQnVfXe5ztsjatSUluO6pJyByBIET1g9AjZhD2E1z7tEn3
fwhB0MhLxf9xh/h9FAWJeen0dG9lvl8/vsoAH9ui6PpIboX3tva1iKOvnAbF7Ft6
Oej0UgyGCa8YMAcXkadSWXjaeQEQTSd1NT7ITsUppEMGcI42IO+wGk7qbb//Bvgp
1b8z+E6atA0sHsret73H94/iDTaP0E8GgQkRXGGOLzdXinkEtp+gVjPk05G08lnL
6PrTR+JHsi3ClVznJnTtzx3JzuFYzur6T6CbNjRuifB3SrBdVccs/NPyQo3RBdii
OYGf9rNep40zliIPtC9X7psZ7EbeZnCtCf5IpB3vMupNstDDL2jiU7oHWEc/xBRw
UBTOseb/X1TNPeuE5xM9gpHLvAPI02SyB/QkixZOjLqAODfA1CT+wT6CuNfy94AO
IWGWPUBuewH0c1ZTpytAj/qr/+Vo1PnPBWvrprc1ViOiJYySVuglUhPJ83IXLYvy
8aNRXz7bGfqf3nnQuPLlYIh9Inwkq0FGB83ub5pracxG4Zk0vi/GYwUe7MTagtV5
iROS2uvsrjDc25/jnDSJduVgK5OPzw9JPEdUoiwwnJzoniZgZKlknod8RkVhcsbM
zApsuf/aJuhYLd3Mf0Cx4gL9EW6hEM9uIYgK8+km/CVo0PEkQE7lDIST2HhkAMZG
M9eB3JzOF2C1QHd3g4yzJ5CqtGLmFf+S7PhqfCDb3cSI/BIRoz9xnzGCbYNlTbjC
TijSNAjmfUCE8tZnM0P4A6S4mQxXeToczSZTCr3QplWHB0n5wsCGJ1ub0o7HsDMp
XNq9DuoThonRbIR2aG9/XTSgYR0EDaq8uLObnO4M6IYi0Z7qGGd5UR/NKonXvkvG
NktgvV/H3fdQbdEH0z87wPbG/KuqgYvo+LndaEGB9XpDCqCHidajMnfuGeudE6eG
9AKw3mEh8utRS92TwQU+3iOx/xrIkZbHybxl5WT87jXpVnWibwuGiHpp7ql3DE3L
wblt30yDkz/YvapZ1FJoNyVvaQciT0UmG1fabLMw0esg+mrPcrFqDuxium7tGNvc
We3BBOGNaLb5RXC8hGX2nqCE3XCNF5DnKqcjK2Zm88I9FfPjNSDS30zRDhuNudZu
yv5bpiCOkDtZHlz+VMlCJLA7xgl7kf1pBhSd2LyiobzwEJssb6oQSs2wRx58MVAp
B/S1AW5gO4/nJcagZgg/H2o2brZzfbg0J0s5fiQmf6KurVoOuAK1Gxd23fQI2ZjW
BMt+9Xly+Yn7qxYDEBwy6XowKS2u+0MeIbbRiiIOVE51YglmE2tgFDBMy5pFtwJQ
cP/2E5TZLcaJBf6MCuJsTemWeNCooxXiGPrKdXQvgCjzRIS1dHyS+l6g3uU7wQ2+
GFFmxOt9fc9MduQlyU7xwpcQsGiL1fBbzin8dNlrRNXOONH+I+TGBlCZMFm7SG0J
6FOjqS0ccjNZRxOMyVgqfGMTtX5ecwtpY2NIigO76Avm1PXLuzECAKwFXKuTkZjs
2u9TzAzoDoW3F/HtaZXtW4vCS19I1WeTaOaLn7+P+QEkFtR9/zejBFQHEot/QX7x
0mQDMu2svsq1pOjBuDuxJymygf4LABe2PzDJWh4EqcgBqbMLrkFq+XNHghveq8RI
iYWhrT93wB1Qesbl0t3yU0K7NUXEYOqdN0MKdVGtHB9N9J7gMxWeRm9ZHS9lxGTG
G1FRPDDtb0sa0DxUO3WPzFgg3zsjgbO7lS5cQLctIke3pyEJb/Po3HmBndqcDfAS
yIYTUhJD3N5fEHFMakzLyaA0GN6M0oVWQvmHockVKlC5bwQJzW6vix9hyEUU2Ori
QIF/5FTRkzv+AC35yvDfgWMoRU1P62XvlG2aP0FzQwNe4KqwOkX9h+2yDNtP9Hvf
HxkyqMdkJBZyZ+ZiasMUi4Z2vFcp8GOs8euAeJm4F9aKXfkh/Y1tTvB1FSd7qEtG
Py3W8Pxoar4hY8vGqyOdB/YhDBYO/RUHrgPotfMpJcl931L3xrZTh0OVVM6lTCdz
HeUil7Ifj13AgCpRZKX/1UeWPF4wYO4Ll+V3FnPQL/kn6VsDWkyrjtVcVJi/PoCw
+IKnfyFFkGTK4dTqExLpIV4qhB54XocTXhx3QHYtZUg1PrymxlbeqGLD2xBEdEn1
L8nTP/zUIQatgKWUIikM/WuMvw5W1uh8Ncbu8bUB1qddQLogVoWPavk4HJAEn1jt
3isUZDPOyD9DddWwIfoZFx8cAtfibCkPgJ0cuBv1TAbOiUFvhMk6nIDif1oLULR1
O8m2poZ9eC5G5ltdORcfdqIBDZb/XFvJlsnNYZiWNnJntxT3iNgPYHuKrndl4/nq
HSerVd7YWBpRnyD+V1jKGBpTNz3LzGd7yCrRLJcDNMvRqhAOrivGhWl+RgJOaDdw
4P8AobwiSFMrvEK6bnjxirrSLEPzC5LBOr6nMPcj4DP3uO7ThOhMOMSLZhbftM7t
WLBAcwWUnoYb0muzOPSmFLq7El4O4aWrH8iW3KuKUfZqncj/ctfbxQ//n7RLUEXg
GkNAkA4tTSIFZcZBTSnm5jxZ4pw0T/NRC1nBPQtt+qe6+IDHrtchCkGtq0xP1/kv
TgOp2Em7dMaVrWklGTdDyQYWhS3ZbcWVQuPv1RbcftNCm7WrOEQVan2otXiyq6Go
ghx4uR+XYMs26IStHe9QcgXddEoVFCmP8QtYLsKeaHGisibcvgkN+lNZUA9BmTbm
ebpTTk3e32MliPq6Hkl15luUOg+RcPBrd9Zox3IqPJvUEmGpBzfNhw7e3p6e98RM
Dhttt2xvlETpCauGpER9pgmOFKYE7Cndl3MwUI40dTPgMe6/sfe7c2ghCVldyqx8
VEHUkrO6tLbqy1gqstcZP2MizR2ZN1wUb0qZJqKmgTs+VP3WJogzNZcVeOME80oU
o3t/Zrp+ZfRAe88GnVbJXzlREE3ev1iuf8y4b1i8ojQrAQNuvNMd40bnnem64XTO
XDELIXzIyhvpuD2zsUScoZJw4OSpTCTdanMtzYtj2gVjNb0jithhY0WRa9mtgT8A
pkPFD3G5bseVt9RoorbNiIjQb//4lBCYnKqbuYOCa+0/vnXGUPsIR1uSTm1oI3Q+
cX2iQzrdQh/sIW/Zyt4RK7QguZK9NcGPlUmFHWbcBT/ANjx2BZ3xFFn+F7qoZI4z
trLklN53hSY8NDCEuBXq7tLCxgT0cOPJv2B+jL70ya2jn3Qy2bG1RjCX/6PPE0IV
cEqKk1AV7uYJOQ21saDO3aD8xLPLeoqe3UE7Fknft3UI7sB+xosMGhK1VnnVRpKA
vKlRaNL9GscUgHrsIMl/OWf3XMTw70A2LxoCpx5pC7VnbyhxNP/Bz72ora5U50TC
ELY8f1TrKlDa2HzddwU4cQ45yZEtawXwFwjTIXJvSW3Co7kUICFlzz8Ti1j/wRv6
QF6kJc1n78zBBnBW+YQ0xa7fpKo2Ai4hJCXJFt4R8Y3TTw98QQTQT7g2yVYJN8AF
Z0m6Sj8axPBq4WAhtn7TMY9aDrpTOduhJ8oJ2gNz0H3JzgutlAZHzyuIXryW83Lz
a3lcjkY1TuOwZMkKuuW0InJd0TqEdcCmoMtdYoAyXQPQdheYC3Hn6/MjaH85zTem
WzDqmpnfgAwaJjyLDUovqzs/d01902Y5nsTbNnk4pPbJRReWkj0+1/1EBHrvBM6N
aX91x3yXHsQhP+/NvfOMJqcSg4ZaHG0iFu235kiKu8h/sWRGSRBEHVXTo36M7e18
UuS+vqhLtL2AwNSk1WZkA7LiRsV5DCr4OIgK3wul+hc8QDHVW/ixH/dLpS8vYWuB
6YWACUYF92gf18c6Z6/wzI9oDGAtQ7I2m1mXZERaGC+GipItsP3H00cZAh07ro0P
vaVOCFL5KimlbaIpv1cOejUqwdcCOQSgBOOULVhS1mcPIMJvqlfUzOC3BSYQ1wn/
LyXEZlfeKz7ddD0vfZhIZJkquBM2yE7IjZ9T5EUa8r6+MGo1AuI8OdNvw93FixD+
tFsxicLv3dAot97TA9JQUtyCndQwj9v8+pT4jzu4gXMI4ykRODKRzEl0GTPXofIh
Ochhgw6uJS5Qsz3dUDE4jQ48xOTmyj6ZJiAN3xFrMJJ50nMpBgjJMQzzEmpVnXvA
59yRyapyVqEgJpatLgW42OjuHuqRsKSWGkpWOEI9ZDAHx5Db6CmbYNRV7YCGu2Or
G//5GjIS3LjtGXVV+M886rMzQvUfOOwP8RnModjAW1M2KFb53rruWX9h+kbKS4NH
6QGmSL2jMbbhNOvcwkM/26pdjVQJLyDxOLP3WfkWJ7DgZNHHdEEomAeHRtofr4ei
/0aITH/ppL7jCLO1Qn8IE923Ou5jX+/C+fgcmZAC/BJajIPxu/68SzycIqanwtVI
Wx7j6Mj4kb78SINPqiyaveyyLy+VBzSLDNznvF+drn3qwG36S8XC52Sl902lW9Ou
UEQawMBa/WSbJ+zEIGPLT9g4qHWTZ/8ekXlekRGE6AScPoRg22jeklI5P9UE6FZS
K/YRddjy2skNq9PVVVEnH8EQFPaFGbx+LP9hjr9eIjxK2Ah77wWclRVvXJTTgPaI
5JJPU9wGNCotMfhCULBMgItsN0XbGfrMcc8YEptvPYV1urIr8JTMY3nLHg6BbWRC
pWOpBkJ7a85n8DKMjpFkdYx1T33NeErh1suPdZ135mFJ3xMDQ4uYbM1arzSmLn81
y66Cp/dby2XePly069CwxJH/EeLtIHNm3P5T1yVmhlTVnEIJUYktMWiEmNJGHXG0
s7aFHXZELKjjvHev3OQtVY8qjs8buRhEQn8EN7X9zqIIoa8mFtibeGDT7T4xAjyR
YlIjJ/asG6swa0U+XLHY6MQNiTy2gOmi85CI83eVD9+xfEKjO5jRQNbotBqy8K+L
uXocL9KNNzun2opEEDq5G91zhRrPx2QveLMnuikn8Zjd4OtNbps7yY239lId3bZu
2KKfZDbsKHsj2SvjX/UBNODuoOhxs2Ne5vs5bcpKfdUpsDnH19O1Uzr069Xwjfp2
ly2qDK8XqgJ1CM5iC+4ffP6ihnynK0eRDGymnCMOrBhWQnfk5uHOQ9oFWRhXie7d
B7FddovmwRC6lUSApFL2/zHmfm1QntdcwGYMqm2hfvvAiBfctCNIvyCOjMHJnKHf
JYZ7+4FQ2PSCHguptUTrC2ZMgIruZuCwD4lTUzwiX+W1FZZ5LrQ6NvJxfBrOU0Sy
hdSnO89J/jveOM2VzVSb1hltECc7+MmpWgHz/OON0/QhDjEpxZed1NdQkvEpfA5k
8p0WlYiqyxRcSTfyTOfGQoUs4QK/ZY9FlRCr2g1n7RBQsVrCS/PYdHbgWa1Cm1Mg
dQ13xmlMJYfiGHpl86WfJqLuWPO7nZZVfXfKutJSn+QCNzp/ISghxb31lXu3ZeiU
8ME2DZg5r6ixT/dV000bZoAPzgfq/dS9CAbskVdDV/xLJIPXPxqAOSGRVJEj1QLA
SR1EotkbmXvaz3r5fjzDnP7X/ATUxT0ievWmX+/R0I2sxaFQYggB+FZtCxyMaARC
2J5ljvDjz0adyQKoJsVdiy0rU+zA4hA60eroP7fRI3llUg4HS/EIEJ5BKCRta8as
+XTqdAvb0QCK6jPjxsEQ7cBaOVWgRBCJuuwU1HOC5Gm9J2BU+G7hCw26LtGmAx76
5ceesaZU+nHC/hREiofkB39KP0MLmgVyp215QHQJhAHfVcSXYhupVvahZBn3lmvn
kcoQqsWZ6IpvYd4iJB8y9Cbvvc/lqmgfmVwuIOP1cqo8tGSD6sXBWNstO/lpmqOp
AxCZdg7ZpBH3+Ncadk+zqpE6XQyhAzLwyIUdk1VfhMVONBzHDdyAkUTKwYPZARjG
d6uQP4i368TzQrRSN4TAyyjiXY9tHefvWdQI7ic2BgXt7Q4nBi67QAj/RJGjknzQ
7mnB2oT6iSxuycRH5IEtZVjyfoWALVO0UcVvrBXlyA8F2QAKlaSBoOmtM+Pj1q46
YmUPedm9SvVL/Q41MHTR0RepQSLKOg2uavFrzcJDqlw8ZqgfAYxQSpk5f3mAMAmj
TdPA8Bvp84QhNWoxaKPx0tDRKd3PMgGbuT0PZ4FA4UsFAro1di3gT/AnruD3HMFl
aoQ97TCY7uTwY2MecvaxIltBoDinzardr2GETmla0BSTgUm8D6YzACGfIJ5Wpsqe
Rdvqf9XANGmN+SeMcHRp2h26fsdI+1P4ofkQAjV3dzyetI3X4SsfRvH0VIjEtC7V
cge07JHeDH9YxH+6iNJRw6FNdDLuuZkgA5UkA8NRYpDHL3jpAAwf9ay9VYUYhIkh
VemPzRBl4K1KOqz2d5YKV/58AZYyzLpn8pLbVD51D/YvM3bDulJiS3GA3QjDl5OX
Qn1dNIuZ13YSCaElSxgnzmYTrqBjQ5LSpCb08PJqPsqGeBT5phLNMDR3X5+qMwTS
CuBb2wUqPMFkBtLWb0VpBPQco83ZwAjD+FHcph878FVY161NL+oKdXYL/tlwj6dF
fSNStIr2GXuBBj9DTqV3IDVfiNVsHZEgCWw+bhY22SvIxNqT77cgDuPLN4jGRz2S
maDl/uicTi0zWtavt+iwqoBh3vtK0U+qR9lrgm5XbLWbHKrRdytbc+MPJStBoS5w
yXeN7qUzE2BjQ/cmFpvFDfQN5HQplC6E2q8JrZAutcLxaGYvit4ifP+WrkfvpBOT
r47ez4/+PionKhPAdvhwRhBM4/hhoUqA9J0BX786L6M4PB3mfnZNCzYF2t1asqGQ
qiZwsyHxYkC8dlj1LrNcwFyHuXHPDcNQx77IwdBYmwkgdsHNreyySJGKjkC7EnLk
+72hgXHXxNJ9DFtq8fe0cO2k1G06MjepVWMZZuFFFzjKxKeWnN89ZC/W+XD+4RSH
KK8qVzO9LyWYaqFLAw9QIvah4IptC4/SMjWxcqOPomDcyUiNwyWaWVriwrUIR6TV
djBmQLezgNUxRgCWqabszwore4RGU8JjLCycFi1NHfN382wyam2q9uSzJtvDtUJO
3DGCbTEa8siFSB5GhDFDoGV3AesRmysm8JwA/QIpixD7nw+Dco8hPXHOGCWMCdd8
GusX1AnGi5CrWw29mmZZxVba/kI395FUBSx/DbEBQhET7J1gBCeSm0lovw3ybPmV
bskVrfOIM6hmcqmhBQJatB8K9y1uwB5TKPQFPE9hbZpZ8m/ZbZH7aKQOhyOyoQiJ
9/h8a3k6VEJy02Vu9+rPKnq2CZ+0JoLpE/Jok+kJW/lBE0ef9jyflvN5Btk09IVk
hEIR9ZcGc4S3GWv7GXPuJ3Ok7pOAYK6ntBGa7I91Ssz0YkAzLS1pLfIqGHqzNz8U
/B3SdA8Q8TA/RHhFhm2MKzVQQ4s3ZK37Sclo4co+QQGp8MdUDm7jVsq10HHmmyvy
kpR4S6U8b6f1X5PwKXWLmY66Df2pZtX6kMVQYZZf+oXbGsdpIHfWFpCQRtylEWhp
1f5iy6g9rtVirlyVQW4EK6y6B25ZpXwVwmWpc0DtKQZB9r1t4VX4IjP58IJ0wL6r
dDGN9ZlOLYd/Bu+ZgawkhmJEEZfiDL1hmOCfCI7kDQOyRCzZvpGXt17b0CIQbt+W
XJpqM7+tlppz0zfBs7YYXz7Cr9o1zH8d3s+0fv246D1vXXFx4ZU2c7IDDbEqUJ2w
XGm73kLPNFJ4G2atdpyco7IoH2Jdt1rZUYNktWQxFIoVhwPZJ372iNPXKasr/b7p
zT/3Vl1mSiiz2kw7x2y0MY7JssKUodRX7hiaDprhxrw6hbhiY9RqIRIeUUIBboFn
/ACFbszhkOkeasx1ZjK1dRdwhAnRIZuQnmd1Ycp6AmMUZvQlBq+5P+c9uVMkp4xy
PkCJE8PBOxA8ouTZTX+6qrQJzdL0HEPC51bGAirSZiaeRx6GZVsMpsRW9YPdLFIG
+1d51ngYF4eFCujZdUEybwzCBXD8/qr5f0A73HkSsHlFE+uiqMaNpvGnQZ/NqYy8
AM0j16oieBi75FVvTlhZ4Tjxwl1rLaiF7ltD3zbZg8mUEOeRyQ/b//8fVoKQu3HJ
90aA4k3lrLsJhCKtfInbX9PvyIS1pjLqOqeboBnhqp/x4DC+6Szzu0H3My1zmT1S
SI6F3nQq7YOjhwoz9TXvA6EijytJ3rWYtUkNMYlqMBFFUhT9UQcb0Ep4H5KJ5niB
dqZMvNg14HRpANrAO1uxhSyVUYAPvoF6EsojZ33fOv5Dx+n6xQ1mRmgpZ18bJKmU
pqNdAzVEeirnOsVFhyGx4lII+rLgdjh2f+5Kkj3Ogny7V3918Ew26pYWwRvD3by+
VwIoqTRYWntY5H6xMOqB6MDUYVaHXPmMpGQrqd+GQW987MeDPNYhT04Wf3IOP8Yx
MlM7NvLxvkT2Fx9fbXKyss8mfL+ig5HkixsTHKuSAp3SExlkoaNEhAExcW9QCm3W
MbzpB6sEBVGFBsgU6qmGDyetn2NYaBcMD9GPGuyyhmxUhHY+zfBRD82303il59f2
Jo8wdznqVOMyV9qBR6GJZQSu1Bbm5lkEucxxqusAUPbkcoj7aX8ssAVAmI387ut5
cTYuR08sY6uZ2zKj1JsRjTrQvIJZRBKH/jK+L30NBYPdzt4DcBdYK935J9flo6nE
LLBuQEvgbvtwajDgm8ySBjpn3HWdBvptf24AU4++C8v6LG6T1rXgaVDcZFr6jkLB
9WmswWN2Unw+GAFsyZA6hLzK/31UeSLO7YkLwXrLfS45tGX+xWZZO5crUs22ACcE
hH5ktM7/68XHIFVYT120hvSYd26Ksxg38cw9F9zUt67jdX5s5kaghox0Q3jET+Uj
E8alHp6bW+p58FwdhQOxyURqdeARoDrx+k0C6X0Ila2T2yYDP8E2Smor7HvsXSdu
0r35Jm3gpn9xAzj38ElF3beoF2ofRz8khSxQbvhyc1Qlrljutz/7DunLshVj8Yw5
aV7seP3rrDxQgSkSX4duGwj2uEVFAQ5klUvHzdl/a816Db9GKjGKUhOr3jPk9dSs
m+z+n9cdtb8Llohtro/aeV1awZifNJXsD/R+KGk1JioYgvdjrri9mU335l0gjXxS
lLUbSeAgh7Hezc7uA0VpIqKXDwDnyTZv+Ix93ZfF2Rec3qVBj7Ux0XKw2EBsSkVM
X4V4/+1tH0ldQ42iXKriAP2i/i3/cb4FR279Ph8eshkcnClUPLDmTPTRfiB5ys3o
OUsQ0gzh/IO6eE+rYtWtyC7//1TG6BrC0MYFMEefB605XjK8Ho0iaBjksQhtJfQq
ueIYdtxc/MSB+xppqVNgKeafFWfWDO8ERfU3p5z6qlQoQe/76kx6w/SJhm7Tr4r5
HRgZzUFKSRatLLp7t7ImlxnxkJ6ksrb2uoVBgidScFjftXb1Fkl6h+RaKhtzBQln
xjzIKyl2FgdCdViy66/3aCbsWdCC4q3tentUkuqWSceT4SK+lrrZP/J7HxZkyj5I
eeFhUqnM3I3/2aDr4iy089UNXp9imIJtnFaGHf62mFYIArPC9AEmeBvSxQwp1LsP
Ui0D3TjwLEK18PgTCLTKkYP3gia7kmTfcnoadJCk85QCDD+SshmvkcdDWnwYXixK
CG1l3sgpS1NiPjp44CLzv37pxf3BoTIvxLctqQ0NSIkAdDaFP2sTYsIaRBMOfSUe
umQCXPR9LgoyLMT71MNrdBW/HGIg51ozioXBnZjS9G83dcPMEZqbPjwVVHg03CN0
8WG7DFbFp6E1xiJbi8Mkq1Lt9TTnf02OI57y0oUTiYYSVQ052ps8IpuU6ngaBI/1
opbRuGaLi0h9vwqYchTaR+E999San/GzTidxz093bNAuuHTBiHHlU+IH0m3OOK/n
gzctgHheFcpfY8JWmlAXBmUUWb5zrWw3o5pfjDcWvSsbwXxGP0dx9zVR6d8JXvb2
2nuYuZ5U2y/dxS8eVZ96QOxMLvR+PD6JgVGUWprKYFZnmHhDO+LZQ2RC2jPZFOrD
EXWqSKJfYcT9bSHPDpWnXjlaNZCBnsztKxYheZbaIXTONdZNOtnVOW2N6TViDjQi
QNaOMSU88ruIWd7CBeCfvpuoBehHFUclg+9QU5NLuinwpb9q+3FUjLR7eQrrw+tv
2oZqOpKyQviPzRZ3bKcJl32SpnoEQ7+hPu6b4TpGfKtFF6tUZFuUEAhGJRaGRIsD
fVMCkc0njh6iw/X9t0AUrn7T1LE/DpMdjGt9gsXNMZuby+z2URTj0Pjd8/Kh5072
uoAibgvkurPyr3o8AiZ7Egn10Y4aBOOX6n8kWuyO4y+g88de7OHLa/BGSwxeysZ6
dtdQWy27xbih5kxwYjqbCtRaVPYYEhmNgu4BOfeOjgF2r616JlhTU+1OyqW2EZzw
NBk5m/y4gebjOoQo1vI+9DTyaiVsJBZspoxybpXlt6kEyX1+2WwVZSBzGPHS3EXL
0pYsCaD1+j5yIOwuRKqSsGKKjJXK+SMeWpQNLs2ob8vmUo3PUjq7qQ0Qe0u7CRJQ
qbJkVqNJiSFpsZNG4KyeoG34UdrKYS8h/WbLkfp4bs4Lkpmwl+OPCiFTRyA8IY5B
d0SmGYSHnkDKVT6lIQLbVAll+Biui5K4u3esHerRAiGchxDuilD35PBJTj4rEmsu
4UeazD+Rl+vBoQMniVqIMOP/8nrlCdvO5TAedhrt7Gg7BxmZ18GzeHhFi0cRnzDp
Ma+942nwQ9WcLi7UaeFbvBDxX2HEdVA9xM5w/D3J+2D4nlhjaQujjq/vLRCyvwza
plBJmJkFIloEyVplt/JvZ78ijowomCUefHCzioOPRkP7f7hWFyDJMMagXt6fnDbC
yrIUUX6OOlzuWfcFMmwsK/fhvrQhOcusvI3KjOlLV+HnS8VHYH5AWJnh0i4N3YSw
C4Lk42nLY+l7d875YeiyVhYT4b60+T91R4kcpWXuVPAO9qf1Q0OH8GeH4urYPrpi
HemQtiq+fvY8Rg3T4H4eoWfOSqDOPqWrlZ+pE6PHB9ABnulcXfq/6CEL0umC8+IK
xtIkbgqz97eUXP94LQdymL67sfTLbdzjU43Q+/fyHPcXl3STgi+IsAsAFd2JjQDD
U2Sj+tLetEg5UEE+OHzDi7Oi/4j/isDu+eTpD9lgGV8D83nznm6jRgIJ1spSofyo
537FerfnjhHVpvIdDL+domiIpftPbjv7X6NTlX1ETuSC72zG9KTEKyZZsyKpk8QA
Hyrt0wvyTSEmwT4YSJHzelfmq+8ZZUNpgAJI0gbiIPZ46FpNvUuEBgPNsRdx4M+C
NomiFXH+nfDvVwoG2RK15DN6k1x1ZjMyiteNTw2TekbooVY0F97ny3svHCaSiFWk
uxeEJY/45IebgGLL7fK7vKgOJUiX1sfRE0/VQoBdchStoK8GjGKbKFP/JcQJDqvQ
R9ooxtO25WHtDN7G3AOa/aTIb0MbKL313UptLOJR7nkgD4JsavMLxc+nMUNzu/Rc
7MErHXhlAALqUj1Tpbh24Mz7iY92lzCFXQXZ5nJJYZLzZfC7qz8smVyq0yvsxHmI
vbjKhhu6pDuElJzFF0tqAoewbXfaWta/3XSn0d01/qzO4Fwdp5DpsZcNbEh5Mst5
1E2Jhs+VFzAIPQoFUzmeERy/f3ORFDNckTPHrPSnQOQiePsCyLkmQ3GbPgBzOQoS
M/NymLNPjAvL80ea7VsT+wzSwGl4e8Xy7DOmRaWYHpwFWFOMeSfIQVA21BeO+BiF
OrRSX+hMlPwL0AQVrL7CXhm9O9nOlkX2fxEPvRm33sVyHk+0HB5jAXRgaw9YR+2m
uX2uEkYHILy9I5dqigo6kAEyCgRWYGV0s1htCGCuABMH5TrgWdz0bZm8VKpdZQI2
6eUpJirzQn1eZnEG+6xNkaln68EkmDnzInDcVCPiEfNPdWUq6zQp67iWz/GKo43l
+QExSQw+weThfd+x2rK1ZogUgs97ipB7xqwDFFJeVuTIuzcvUqto+4LEmH+Mh5Xj
329p6ZXDxVGdDv4S0SWRhJlqIfAKN87FAAGMl0PnbMmLzw9bNOGtZdFeans1H5/B
3FRe8QV6cpuamgo8wVPpGyVA/w105oDpAZEmZP8yUWPXfJdKEGn04bGIDdRj/wwc
i8r7TpFga1ZLj8rdOYHoVlwhsMyFXAPvyxyFU0FG0w4MeXWIoUoSv5pQewEloXCT
+XJALr31BErxC/Ei6JAlJsTMIApW5+BmVnn/qyuT91zFgA096QJp9skYlJMoY6i5
p9tvzQSuVpJ/7IgWM4QIuSNHbSIMqnvVpISLinojm42Jz/d298aCaIuVA5RSzYVv
+Z2diYSJB7mAMpZsnaDZdZ5IKYzQou7zODxHb58tWnwfdMFcbqs6F4c7fgUVSi7B
IGY95V2opDQ7JG6DKgqkc1QCmLM3Sy6HJ7ofo09xxtzTwIsTP7oDPNYcQzEPv269
JrDz2zOT7Pd1zXCBoq0ZNQgL2RQMuxs3zBDYXRuwSzKKo18+iBY+JY1W5G9uHThd
aVm/DHg3ZA0UpikHpTOU3AIHk/SpXUeFdWDHQ4UbX8dWfK9CGmaNVmVT23s/vSx4
U5JX41HyrgQd4MtupbkCXadE4w333NzDBDTDjb2bwCI0qoG5NITopRxzMvkArW+o
gjdKcvUfyLO+dYh6MGl9BcANhWA0FwGU01HPBHDgCUoJvB1PePFTjaUinXVg92fJ
5GL68kU1rvjIVuMRcC42FNCFrUBYsA9vVOsVIcjDsp+xlLqX7f8gjDMA5zjShRn4
ahXNozXtti8GNsJop+2iUqT15lVHMVDhzKIKgurYX/d3a7LY3LRPnLaFYdZaAhSt
iYMuFlTKJtVBHrzzrulxXyw7GeF96XagJauYBKE7bKVdUJRFDngj3kUL7y9fsVAq
S+XD8215Og/uY/k1TzdpUQB3M4Cjgk2Ti3IHWF/KdTpLvbH1OfbrJ4R7W/LaMeD5
4/HbEzhgTmTfDDsCMrn5EqUOdZduh4EWFsdqKfZsSi665YJxrFS1NndqMBx//oqH
wWTVUpuOuanGKFj93Vt0glD9qZmNvZIsc3dfieUxnND1XmrRpOCked9/f3fLChW+
/6i3br1NjR0AW/xua/qXaoc8kdZErz4Q+6sSoiKmrLI25SJs/zo78BMM0vWZ9Ucz
SafmNJ0WEb5z1F+45sRDgP/y3K/T0tuNVDOTLbuCxRSdHaAJjea70CZc6fgru+e1
wAxdBMJZHANh8T42BI8sFMkzZyO1n3iJ+9e1zss45+T00cxPtS3MzubfarsK/8Ck
emwpy2j3CwFf0XOpPQ0NtSN5RmVxN+Xh5lPX2b5ONqyPRH5KegQh8egnf9PgSEwK
CXhofOQOkAtB6fmw4VZhZF0i1vP/5/ZylmY+2sDGJV2MNRRSe5sB/SXkCym75A4a
auO9jOHJB37eUg299dZu67IYiVXSk/lzknYYzofUU/bQC2iQfpliFY1GynURUyIt
m8RKMsV5vBXVM7HGXFNh4XRfiYfojGaX6BeuqnXtcLa+tK3I4sn1rrOJGRZmSJ1B
v7irx46sDlVHOtOR+kJAxnXLDYjdHVMb//Aa7KF//A4KUxk6xznDARp+439GFn5r
8oLqe7Nhjpd/Us/I+1tZ2IN4h5j85jhmLFyWwh2iza583umtE03+pclSOVrxWIFu
ZQ6JEwHMq8NLoA+nCc7mRdjE3ZsPxrKcreo/y4eJtVhVWoWNcAoB59CYZRRQi2eU
PfHiSOznFbmtXqLXIGwkayo20PWdeNmXMv6Tg1BbmqeuB2VOOzz/S5Ug/PUgSiR/
Lx1QUmnQ3X2nK4B5YVAQrw/Q0J9lgAc693OoecEILU+irBegoJGoYuVghyMuwhac
OcZzyz4B2kYGtUL/9H5lTxFGm7/toPpFW2mpFh1QEUi4pqHeG3J5Gfglt556SFuy
A+lLW91jb2xfpaxrTtKe8z9i57KqOiAEPoT5ESGtcAO2VOB24cSpIFsciZn/Cn0H
7RfWFMhP8HRGoTTU5YvY+10CVZ0y3dsKt3TLGVEX6Nx/cebvHDTnxscEtP/hoWxn
53G5+d7ir4YBG3sjjG0mFtGFhIE1dRe4eukayX5GA0tLn3QsYFXSnSQmaU9uKGj8
eoI9E5qvezXQi/QWOPkVYgvnOwhYdRVQGXrAZJ++3aXnMr1uGMtjyzIsC7Q+8lZU
qXiRC6zpmIg4McQxMOywG7GDqzb/K7DBrfvA0ZE/ZVel6lQlC8Qk7JUm0uCQ4i5E
iqnofpCKCJj3+rNoM38V8WDQOgArTcs5kQZZUl9U6jr+WZFjHOmgzUq1Ppqy3aVP
24NV93D6GCLxwgdfGM0X/UDN0iVbAPgRR+J/Dov0yLI+7bBq1eKwviZjZdgOQ/12
vFPuDrwsT380KblqzkU5txUGeT5Oy8puigC/p6fm3MPwOWzXYOE1XvUBAm7cGaNN
Zy5XPdEWoZi5jHmfdOwTVY/i6xcW7Fj5iUzH/NRusrnfo9rSjVgaWqVDDpFF1G2E
ieF7r8BETy+6ca6BvxMWaP1D4esVbPbkt3OVi0TZ9+fiFHrqvDBEV0XtyWg3GWlF
qPxALv42V9GF/9pjTaKnvMmm/OkqqMT+USfGSA+cj5cLLiXEKa9Ew4iD6lJMKnWY
XuvSS53ggnOIAi4N+5if2D9FCnmD6zxIe+jgDbMsrY6AZASr6pEaiUOKto7OeQox
TcCEnYJHYuqfCL7hIi38OUhHWhZ6xOl0gnefPXUvYeuJW4iKgWUlJvcHD3yfz9jA
9hfQUQZxxMuLJZ/z9hoX/WgujPE0KYCi92KAS8AzazIOXyp5q6o6E3k4CsPi0x3l
Gg3OsiSLdrzkNm7QoQ1i9X/xIuMARH9n2znkU3JzQw5hT4s6gnL0eMlRJg0F4Vrf
RyZoz6rOZEg1bsHYHUrgziDEjjcTdRr+S80CwOyGZ8/JRuxYqUDxeCH41jn5c7eb
M8agfy0pcPeX9Qwki/f/iy7kKwq/s1Xk9ASo2QVUv3fQDHciVYVtYBsZiMj2Ub/w
ELV9aBT8INO1t5ppHL2UMQKBMHMWmWPyaIBQas/838toEJ7QpfRaJQE6hiW5YZEa
XppQ5OgohoGQqIQ0j0TGsOcq3CtvglmypLtZBtZ1Lr0bx/foo6d5SJfzA5frEwn+
5kRrgpFz5WY09j2fpXNF39+hZWjARB+2Diy3woiRLN1x0MJQtcK9BWP5MQExX2aR
EvnD+GvuFd9tSUgxCBKjNSJyP1n/Wi2xxzVA1Zw+Nd1/eZb96GrD+oe3tLPU3D7T
0V7efnD5uFaMVLxh++vmFeJOltgHDDXENfpLPex2Y0Y5o4HikiYOAiO3bvyJDUbE
BgZ9328pqNeCVNhqgIeqRC/VQ8VeTaGOCwu6vF+2r28VMZz4UkN+ifRHXokoN3Pr
QKyPR1O9j/8Nn2UBx9C5gVq8771I37B7oBWtRmk2UIXUsZ61eWujijCrLgHmcypQ
MqWv603ZUD86f6CgDEXCOq3DutZ3eu1dlMRJbVAlu8PJILWKad5nJ9QHvd3lF/7O
wxRC1wzLzIk0+jhBvnHcABjjZZLW12BBpehsrD0rwIdOzL5tY/ppkmhH6geZ9Y3C
8CuuD9z0tL5qDZz0MnLFCqrhzAB20JlS4zbv+T/uaH1tjdN46hrLwccLfzOkVORi
hSNVDL9pfIlCnVqcp5lGMn0t/zaxRCHQrd84+cp+ZSeQzuIwDJ+Men87hkQjZS6b
xbTfMMShwwgSmrqltpxErAPSFtiOVGmU/TzVhJUuHDGmosrDYWQl7xxvTDbh1Y26
ACUXMl61fvEtsGro694NfYRF3osw8scvcYr5d5DVM3N8Wta1t1JZJidQKe7jRXE2
j9eLdbvLXI4ETEj7kfY+Vl6uPo+gvxke9rtKeaTemXpOCFa0Ysc1gQJoKsWwP6JE
8b7UdIsEHzGde3AKC1pWDhBXpcL87eN544/P9g2l1yKyKENVA5x3W7cSd/sjjvTe
kf8ssEBhVpmEm4Vi1Eg5q8+DBNVBJ90+MZ4zP+gmdgp5vs4Oe+CTUDe/JOoyrCgT
x0GmFPvTuUqCS4vbbdOhb0n+CyiwgadctcdltDQpql+P7VhE2K99NEDKerptSIRD
XZTxdxTlJ/9pWxUcKxcMcMF+J1TAv7Jc7EOklSGJgfpIXomuVxXK5u+KqFMmFLOc
2WWZj3Z6+SsF10InrqNrEsD3iVTolFsJD5Qtj6baPgRiS371an8dLAs2ARYNzbtu
S8/ihzOUnRQIIS3qjTms8jqdk8ft3JU6TEO+0FNLoXyA2Bf3GrnPdaC3Nu0VTGBS
CH/QFDyIAW7QAjEVgQsDtymmYjbDdiqvNyytQSE/v8Gn3fBI1ZcQDkaJuhmGl5DS
nkH8my1aq0rrz1BGeNncQlsFDpApMb1fLevBvVH5IsvoUiFkFDT2akgUvsStnstn
I7BiaES6/eq6k9fLnR+uK6Yv26/j5pEvEMPcwoAi4lrDLnjZ8y5oRw1RjfU3UNB4
GoF+yXSnuyICruwAXADF0ScR46uTuSpAEuoAUxiOpZt0UpuRTk1PC2OAmnUrMe0W
RRRMd5xAu3f3l2wCN2DQUMkKc8amPKCkRtJimF74mvrv7JyClPkJ94cTVoiRI7dC
tahgrXgd1AyzdzPIY11ZiSURfO/Ph25B4uLwumQJqODo2UC3fs/Yy2dBJMJrhckn
dbRJDmkMtzNqkDbkRHZFC6tbLpaci87/9dHSn3qOKrMlAZNFvJB90NJti0k8Zjnw
DqVWsbKsXyPknqylM1zb35aXiq0yLPkR2OXJgMPgPCmTLokrfGQUDYYlP4SscWHx
ieasXY+2p5Z3xLWDB9dn8m24kq/Xtn8iZCmzkkTfBMEnWSKjwQOtiIBi0MliHjQh
BTz6BtebCrlOGdpxDYEhIiAiEUunMnM2a//PVv7MWMrPLNn9yy2idJtngOzziMC0
O+A+rGjjthwIKjTmSkZq/lzNKL/fwP/abbUXlAOlFyktTVzUL5h0qnXvefDoL08r
XPdZ3xaNVtCU1VYmC9US09TcRZWwc7prewpAsXXoYaq6booJ7V4/Pay1NJ9Uml3L
FpIBdhmaL/k7mlzOd64gJ70HMlx2cqb+dGAqDbzFvlbAV9QiP3vzDR0gPiya5k+b
HzVGNQEtuWadcJqiwa5SzW4sXc3u1oa4A7adWtDa8W9leyzucAf7lrkHM5PXCYbj
L7LOfJCgvFdYv5PGXS3uhSOt+xO3e9Ap+4TDyclLFLF+eu9fIfuAm9eBnKL4rfny
7674JMNDifU/7l+14JsTVX2/vZiDRwI4ioTGfTwlXGBywiYpE9ABglUrJowR3S6H
++cyxKEJS/CZS0RzR2PMQ5xNSbJdzaDrdJBXKXIfwXD2+FrjbTn62NU+UO7wxfIP
w/T4/w4cY4MU/SfUyhShQW84v9exzSunvdUSNgwHhudsbfhmQmSKHBO596sohULB
vmGUuqoMFwf7VpGDMhp375cvBzObf6TWlP1BREjTZPbYRyQNrIbQ9I8aem0AY8NL
/t6UMYhE5vzPczpMoFPSOyUQIIivqm2HzVP9oIJNIC5oyPvJrggpg2ldpep16fzq
HU2gNqi3CX0JQ236AuBVdMamf2hkHK+UW3RHnFM3yQ/uZuZQzZNztNvYYA25I66P
s3YkDTVu3iBuLmfQ6If6ESjoooNqrG2/LiMB2MU+UOyPXGYWCDdRpBggijroZILS
tRr1sMKhUC/147tb8dyfwwRxyVHePvp46XbLYpFlAmXFRQT4hugHk2rMY6mYEtLM
6HSGiADtfxVYlOhTc9wyV0k3hVpZhPsA1ALuFvihDNgKNI1w2WmySmVA8JWHR13b
yZ2ZOIqnFFoJxFXXFGqVru2eoVo4vWm6J6V1GSGQAIcLKAESSH7Ec1I7BCKeo5VX
Cf7Fu+9pb9A7LkhyBOrgHkRc8Ynl3sc/F81FmOJFi1R/XNDqkN6cuWYGRQBt1bTq
U/AZSFbUhJR/lP9JYwYd2svPU5Pgz3fxCEcFDryoQtK7XjwjW9McnHScl5zWhki9
29eJThcOA+e9npf4fZvSfpZKYMLtneUr+ecCBggBHwTGgFOHCTPrBk9p5pbnSGm2
hAsU1clYuKB3QhMkBya8NTw4eU/T5FoSnTr4jHS3SRQrhk/ivStw6vYGG5ePXFnB
hAoELDSyu1g6WVDgEwZT+8W72iaEwz16ovY++Hmj2i4ko3cjtR4pBp/rkEfDrkxF
22Np6E3gO00VQVisMG3iVQaarlzpWytizoCsKsrlKE9gCJblleIdMA9s5ZW6QHKF
y03oPhgwRCzgShLEY9fhzEcknPyzZy0LYuO6WvrRbjIKvS2lWNvQjXu2VLHaPXNH
EtDkrKjtMEqgXPsP0ZvL+bv2IyDYi9n+FjmDaDvpx4+i9YZEbBV9EeqiDQ8WRU79
TcenHBJ/teXq3iZi9l7M1VAUQCAiuisLX6fGabXq+2g1Evpp9veF8nbqGYrBsFQy
Pjz7b6XAz3GHy2V5dCGwY18tNY5p5TZ3k4/e7P6tymBRuqSzWpCqQQjJrOl5xGw1
DrZmajWNoL+tyLR32qTBfupZybAbm58X3DlIBAA3Y24Z9/jhVRh23oZPthtTxBMy
z4SSLg3eG01wiGklLpz+PwbaSohOpnvLz3T4N+uo+myZCV7xAoXPNjhGliSVP0VT
sOEnEzLp1hSVSIxMRN9sLcL8+9RDeA7/KLZdAi18aFDewHDzDFAWB/xmDH+CLgky
GDeslzg1+xb1HmCLlmiqeqnhg84Xga1nXeCQpb5FlNjDQdorJmu4lwM13Ew3Ag+l
HlhvoFS8D0hyqslPJ3fhmdXb7yEDqYxqVE/VNqODgRlSsL6Pjk+WnXjVlMfZm8p0
9x1O2KA+ntPjWfkZOg/lrBiWvHb6ethqcNUam/UtS7f74yso+pnBN+jvmvUEauMj
AdK4M+Q5ibqCOE5OtKbewq1WbkF65gfpcjG7YJ6TXvo8DAsjVx9BQ+jP6SlH7Koe
gsAoDbL2Jf838/ydiVOhTrgMN1bzVMevgi1tFuW+lxiE+A6JWbuNG2AcVxis3d1L
VRqjx8Xz922mBcanX3kmOlhUZZOxqfZIVzNGO+HzgpKo+BXZZwQC4GGUKw1aIIbL
7Ur9h5LTjomMJTkQD28HxD/wMvRZtVFjziW28hirR/SJzYBlBqgQdNSL6R4yI/Ax
oCDtufDBCSnLE5breRnGBrCInO2mks75j+ADK00riIJlS5Qsk5g0+JYS5YxtB4sd
W20LcrNEK5eMR1FTesmT/TJlTgvluf3/Mqz8J0BDMDL7yJ4xzt0JHmzcRy00+ukJ
DhHGjDtYO4Iwt7c9MxtJhxVK63HGSDRmOnN4IWLjVZOYvcSd2gFFsHaB3Qf0HaxY
BZnA3JvWmJtL+KLnViKuhqlQiYsVGuoV7ioJm5hehaPfwhia7oJjLFsSpxx0ji9r
ljHKBXEGfXSjfhchGADhSGooIMSqNryuJuEh11ACXKDhWvxIMy75ceAMl7l9eJHf
Dez01n7WX9DZM3oWpSsnO3fq/NUJg6RbA3PucqtdpOZjKXM2Y/cfZQk0itHb8Dgc
OWb1WaoeJ/uXRIfZz8/XGhJ+KZ6HZgDE4/Nt1pdz7l0pzvlphudsUJtsbYcWYMVt
VRXbYgtPa5cSSAg1jsa+wBL3LUlxxJZiN9+TajrR5jREmz8I5G9PXLy2t0mXNuWU
iyBF1/8ICaQB4ImNLoq6aDnKC6RT8rqO9rukwAJ6UdOOUMGDAB8YfHEFk+LVngtO
2o37IAbG4A9g3N1yuA2TUl/f89TxbbSXhl7hI7tpwg7kP0junRucQdXAebRpA3vN
J6BdjRCw4lvOCQvLXCutVwlRdIdOFko2UGhJcwn8nYbA6pcGR5OMS/wSw4Gmzz57
Jm3R5YptHGYIZZxI3i/kcRfCLFq15cquDrFs+lkesC5uIIsJ+O7vfrlgXid42u+5
4SwWoDocPpQIfeiL0AvWumHDrQy4vsvXH3BMnMlcWOmnR+8qbl87YfiL21JxLmEK
4VLNRR8WfLOkz2JBxAPIp/zXhNZVOdy2Bu3ssVmC+EJi5oAXEWldIcR1HAJaBkFa
i2jS4snFuTmtSlxJIW+GGAiIpfPy/GYLz5B/VtAXUa9VpFboXzoN40BdKbBnD7XJ
UkhRtW5WTt6YYahSqNsa7C7vNdnCbNcXJLjOfSdOmF+dbIY0Or6KE6say3FuiDPw
MqJlrNtHC3jswztDe+rqYNeE9ag2PHMtW8lde+cZbR9Et0pthx6/0fyDQaaqPgiQ
mp1Ar+2WWOGXPvSf/SlPJj0MtYkNAXHjExMjvAdrCcYcG7ZaC6OWYJHdtjGLd7OJ
VcB9yi8VtcZRLfR1erVKynffPiXIgCABTCBRN4eVlhpib3T2OW1TpehxfHW6Fyu6
+JnD/jAtHfM0mAq2LS2TUCTEmtt1zl5eBBJSGBxn1JRng0AobHOXStQIixoff8AA
aGtGZrSUYIaPYTXXhC4w6JLpZ1piZd68EfTp2xxrjT7dWVI8v3CIJcRGSbXBVPPT
7X55sCkZVJEF2O26JIxSqfGyb/BuAqbRLvmIWI66WIglnL+DTtmA3itbM6Kkz7ij
fzByG+B7FzxsdgmVKd99nKhHZgWyevDWdRHO6DJdhmgaeugFGXhXcMyiN2k/RjpS
6N6ZloCYXlSEFQveQPJt5Alh09IRVKA0TXxd1tc3W7n4TxfaJFGeyoR+XCU0YScZ
Snf3A16S9nxCRJajsPLYieOYBbuThyZKpjbYcVxaKKKK7E3Lp1Vc1QTKHPpMtPu/
ymRB+8eZKZX2p07OEW2r5gnzKyXXgIbrveDgRp2mi8FVnFNxhlIBljMuKp3ew5qZ
qRMC1vplSbB0BrgJkze5KkAHF/kWFNn7tdHmvLjFk6YFGMlyetIjb1KUpkhOR5+M
s9s4Rgn9LaV+AAObFDpKAz9gfS5ReqFVzeoVxhuGWBoIxxp8hmx2KdHCZ/roG7U9
OH6c/sAgJzSPM8EmFs/ctNbKHAfW26uHpc7B3G5CUrG0iTdkRzcuNCSqF5tYvmcz
KCg113LTcfUH9ZfYE66V+e49kWvX1JnjMMathGITpP7sBWYSCINYwn75WukfFdoR
DoDPURV3e39vPwg/Fk7hmOomNMyCx33fh9BEW3LXAgXu4aTQG2wRYBwK33i+/JCg
mzMNx81ryeH7zIGEmwFv80TgjSS19HpOwob5hSYODMH1/7CPoq3uwq1KDR26u6au
1Bkku9+9zZq5Xu+3wdTN3nBqaAFT7uvDfrCJ5OHltO5OKBmyxxWOMHM08u7Kzigg
3HATfEhrVbDAtF7OSMYnAbZ2WyqtXAjOcfMlN+v4MinQ2nP5SlplGkzxosnXvDOL
lvn7HlxssXey+H+4lF+GmWuCvF0v/7m6tBWN7UF85LrP5/D4UcsnAacfeLfmzjQt
/y3a2uZWw2Utfy+ukx299IuiEsBjC+mocyk61/iDETBSgmf1NnMrvIZ0vubnJKqo
xX2Rjzv1z+z4L1F573qklkSJEw66EfNbRp/AdWHX99pTpOB0Zy3nsLPZeHnn/Cxh
n7UhQ896GAx2OWGcz4ySVEvg4hq6aht2aDgdE/DOOBLg4jgcc41kJmfB/RpoWEVV
KFG/ru52btqoyybIzzzArwM1FfJ+SFXMfIG3MsZqUp8DxcFDbP4ZzaKjDYZwpEKh
nsu7HtpRdKWxtia2N+BwtOgzXjwIM24zSk7Qo9hpuM4VAQC6RbI2AtfcPx47qJm7
oC3nH7743/G0hBYRSjxj5a8XgDLWyhEKQ4efQQmQ58JzgaqRh/NU7UkrWPu6z6qD
LLmtOPtF9MsEDcnVcdquHEKEfHP5wm2UQsluLONqgLQCBbijrx0T3rHR4gCPpFeP
mR1U+LlE31c9EuAgG8UDrWj6i7v9/5vQXVGacIv66fl4Fg9PregQUCNQe6yx6DGF
DkFGFU+udhX5y9KFvElyImMvsgVHzt4ZLbX5VlmOumzwtC0lhGfCPuHG67Sj+l5m
P9f2PIUPHyPF3+WOGTEA8r7JsIQ5N0oe0b2TuNlqjmNPaKJ2+cZ7p29bB/wHZqi4
5alNJ2MxwtQGMS/kCCP1cRrsfCHwCfLDSZXASL8O2Y1rTe1TeOhV54qq1yHgtnSK
bNl86tyoXjfgYwT/7V7fecBe02qqm5ageN26fshDIqzwm8uNn6Vk6dR/9xI65x3c
q22koLh4lwizYljUMonGOJag1W+mrz/6QY9oapz1U4FhHZLwq4uvo/J82upZROb3
jkBbQFT2WZn6ExT3q4mZihTw2NuLcvwK0gVWUO62B1dTnLK+blQTCBz/sYgow5y9
gkNepQ5GBljKTiQKHWvb53AwNH6i5TdrgNaZREH2iwH7nb4bq5FtCUV+xPtc43un
v6ha8dCCFg9QZCMjR42O5Ins/xa7bDqCnaVPwmB+0XR9GXEFCB+04X/iXg5yzr3d
hWIxzwxSAjADL4E9WdSnrnNVPm7K8caXruHUjaMnTZe6vVlgPUsftIA/M5c8fAjf
bhVsyVulvvTM0bxNhhLQ3u9fUPml0CixFR6uhyUIomukkcfoYFsMIOx1rgCYPej7
n6oZHVLEhr+fOXaQeqXliyjFScCVWVIZ7U1kAiv4Z9HXAKzTgc3ppJQxxhH/cUpp
0I89a2eEE2gAFVtWKGlXMJ6nlJOykMfUJmI2ECcyxyx5AOE88CqqjQGBmy/gP0Vh
SrwLcfMZ5tI3gtupi8SPbyCa057jta4HZvWA2lEvk1ghtlNtIoWx2q4T8IAwyGhd
aB+pywfdG9FvAfaWuw9c9bFBLc15UmXS8F5eNviSl5f2jOOa9MYYoOQqBL4RSRWr
mDN8fPTqK5nfE7AatE9oEDxlSdUj0MbWQe8hmFlgdc+T285jDDEn+TANpxW7rZHP
htVqFyXWOemTX5EnG6b4qCjMRHmoYGHtai4sZUmz6j4gPDJWSBaydCHoSQag5ccD
9lru46dhQd8UBzj6cmFIcuOOPy4w1jFHV6xGXVhNwABHVpzCi491imH6UuzNwfPG
MPzR1WaqoCn2mDAugXrJ8B1VOP/LkWEhhcQkTFmcGbAudO1KmElGhu5zc0t/9Eaj
xdlupotUsUfYBu2B/Q4MGXz+BqnZbaGS5SHcGdIFDFoTIBR92tTBXN0WjpJYMCWv
DmVHL/JovdU+SwjHzhzULNKUO3vZOHBwqAIl1/cLZfqFzsPn5fYPatBsquEdZO1t
kzadAsIVYkvwKqnshTApPrVDyDf7CZam80cjIGrAUlLpAFL9h2gKRdRxy7P4tcMi
HkpHVUiCnURQCLKF4Cx8jMXS2yUiOWim5G5+ph7VMPWPN4BneR2MKZG9ZrFrlKtp
tqYhfktGeFLlNQHOdRX95EqGwKveV3gSXPujYPbc2UY8m4rARbJt3pfrPc3/ligB
ALwXx432sqm8jBM/sKGx5qEwU5gWQlQKlYu/I5xddAAJcPxTAGgIJgFyE6PfFKQt
dk2CY/MoQ4AYY375RXpNZZ6DgNBV4KqXRmYI0BZO8NFjMTJlEhDAsk3GFzSrwtyL
BA8xhOfzjFlq+836cD7F3u5c0zuMF+W4SYz51tAtz1qH26sMKQMtYf/esu2R0cJk
x9g9yWefz+zKdBKeDX2yJNbqXt/Z0wfjJqC046hXpZ52RWHzRxLO90SKbErUrQO5
Lg/joQi273uvg5L84S0pUxQYrF72hEQQn6YdiFSfl7pr46cZ1bDKjdtyDcBiwgRb
JUXudQiHRFGvgx8erHNfif/RCtybqXjItKwJqTRCuAlYtVB3EeuaFxuriW9rk4ti
PlORBUlrP3xJxNxn9kisi4SIiHyd1dqVz/jn9UCby8DGDMnj/LY5cOKgD0k/uFLq
UkHO6RhswYBrkoXLTsVjY4PBMetYeolnX4aTIG3z0+LlAC0FuJ6lMN87Hhq674Sp
cLtoB+INmD9kFJgAXMRea8iqfHhVkLD+fLmCivPD7NRQIuucuwcMorWfWJubo4rY
WptPSRw5oozXv3TLuZjW/hcgvnbDDDD8UMCe4W1Z/wkHHEeLS9XLnPzl3fyfs9S3
yWqzeOxwC+cU0OuxHdWY8MwukJEtWXWySwpMEQmgHGj/6kwecs7ZgjX6l+12fR7Y
dySdwJxV3uMcFBbmXMw0CUi1L0Fr4+YSMs6gx8cmuqwxxbcEBEG9EleY0/u19fUh
el64IkMtm/eY1E59QyufTyrXJMHFxfOSGEYC9Qfdt+1eEYzdgidK7GEBwKF+uhEy
NBCXquajfEnLagjMKTdpmf8LgALpkP3Mre5EscB4tdgS9H2ITi3utPmLiuXowZVq
+5m2HZ0XgTf4IiidLtkfczXf6f1y4WH03QLix0ENC1D29Aa8RKRhs5aXHWvvFrBs
Ap49jEpRTzanyJxkB5CiVhC1VR05m1dwRFh30dmKMUCguw1pRdSpcM+9K8+jsNwa
aoM2k6tzz8EbvJJaB4jWDBk9WbsF0N2E73aBXbX3Vq1Xo7DCYjUuuQ4uYayknuLH
Qh6MvyhZSuVrBoaZHGUvelwhVP0KU9+8mNqYLzl2VUJfB4Zilc53ySEX3wvVgJBn
itoN/b4MeRv93BNWQD6sI+UrdzSRSRk0b0Jp4nJPWZGAF1bgiFuuO8bIWpLY2ScD
RLYCj+w/IsNUoDSqFRFpJmuqARaGZMYAXvUoju5apzTKU6MNQXDyPyhoWZK/ILtj
8/tle0ojj/hmB+b+WYkekE8VKCIEg3vcqFYbp18BJPDTfOJGZmg1hpfDBNGBoqPN
u9tJOkfSnzNz1ScKJSb08PlzCJX4M35zwIX21awHht42Enx6P7pDQRRF4tsG0Pv1
iVOWoFPH7lqKOEfld0KoH+dXr/hUvItH4ET+m6OSUOQpj9GPG2ahqwtEyoJVss8Q
ovxOmE8sKNyv/Ful95rlV55Q+uwHAYaiJg/DJmz26ry2GsT6tUhaJs0uHuQi+c4Q
C9+qXJJGGjvmaLZVkaKA06VSouXe8RKNstivY3tYKIOKLGlaZjDr/TlQj4Ka+HeU
luH+Z6i1o9xw1aFdoYcGMfy3o1cqhPkC0ym3bG3GE+4im+p2txwhEy0yz431p1CV
drRO0/64oeUrURf7lX9j3htwkpNWMFJElxO4IF2KI22Jo2Fc7qxm3lNv2x3IQcQW
+XRkCCmU2+zD+t+tz5xYLj2PzPMYVMJZq9qE6GoIYPQbkJC/CpTCXY6W4sIc2Axo
x32mLzkV1W1Vy7q0toRvhNTx1g+pmcgSXinvEYPjNVYbGUP7K9Q+BhoNHSW2/nvi
R99qQTJQAsd5HagR8ucovDzir1hhGAFfosf7Gv3RU+DUJRIGtCkFYZUhn2N8KK2a
5JHySXEE1FfqVdwgzPrSr4UYbfcjjVfmsl0/v4XS8z3jREEMnrrCrbr+znW7sayi
2vn7IjZ64c8PbryQgbA+RiyzFwPloemhXqG8EqnJKuskCcZ0UgpDvqVX5Iq5zHVh
gTC+xcIArONnCLH8oGG35qkDIUD60vrSk5QPaWSrUBtcJwgLYoLHsq9aqoLbC+gt
XLgbIDlpchW9v6IqltaAs54SI01D49bUEinkUpBSpG3B3qriMjZRxbQICEvVjVrY
qNfaNcV5wE5NHZBAvbFWeaB6i4Lw53OSRdd2pgfgi1RYbu7BzfM6kRDBjccgPkxI
YLnYVuO2ZrFkXYy56bFA8B6JFh+Tu7jr4gSBVv+iiA0FSHTTBhJv1CcS0uO5EWqO
XsaPqDbPB9pKLDRFyaK3/YcR2EH71+6+eew0tcQ7fVlk1OAx9XbOAOZynyvb90WT
8bAyOsAI9eWvpzK7c0vkjwLtGQxE8QI/JcmCwdAlT0OZRsfkE2IEDxmvg/fVrBhS
6lox1c0n2Tit0z9pgUOfMvac8HHviIZxn/7167kP5NymHhHIWaSmnlZWMVuFiTKZ
7lGj0x9l9YjCox+6wp+ApwfCdIRw7JAtY6OpY0tquYR2mWm/1ZNgep8jX2QhRusp
hDi0PXV6vwmJH9UUgdidxzX/TNHH7Vh19wyZakXhkY0HpnsWVo/DUfc3obqe8JkO
ocA2OWTpS+X2fIVQxqgVEOI6HhAv5mIRGUDUqIFJjQqe6MxaQbsfQy9Kz7k1Zp01
dPp8Eg9pqJ8mgzDGFYguxwjkd3ccKgdNDX88E8zaIPwMoK4CKIhMdmpMRxGcoATj
NBF9PBNbuBV1+KmbrNC6LGJ1unRsNO4eALlA1rvzi9jtqF68FB1u+qsGvMYgkXkm
Y1XQBLFHLbIWCblFsxs/RxwF6RHXaoHsFCkVjpp2NLjX5tZhgbyIg1u7nRI7GiVI
LX1luf3sb2zxT6ylQOEF8ljO1LFrLLPuYJ65N9k4INk+e80WNyJs6lDVEieaXyky
IooU/lZGQo2R6k5/o9X/qGW686FC8OGNGlI10Los7l6qVsuNFSwUKt3FXcX3zQuI
cQifEbskej5Jy4NxKw9IyKixAa2xmPO1Tw9zBjOC4pxNalJE7Ze9DtfC9ZQgsZjp
0xcdsMzICVqJWuUbkg59vYpCBGgvv/75SIYSZTyIdVwp9wljdbyq30zaV6Mj7zEf
++ZeJ2kAisMZWXtMEkpKoslwNpXjjiPvaQzuDjf9cOBC3wAlYeUQIOKF4xz+bJK1
abvlq58uh/4opDSnV5wn8iuMFbypLsqjzp24YgWL8iajtDX593ZxtIjzNO8aPIJ1
CcEFt/oxNfRii+MNiVK4IWLX1RaOJt693ypHolfk+h2s2QMFDvsBLEr4A9pcXGA1
Pfm7n9pZg345hM3Mxdrq86+Vn9JN/tNHq0OY2u/rte4o8uUQy8oWkfQCp9rmba1V
y23iHJ8NT1/4sviJKUa11NNGGNFfsQDwgdWDmzyV3+DYYntZmmu4dWPrnSBnTgr0
+fKmEKwGyuc+QNJG8pztbHuLLs4dhJQJaQY958eosJCKcInWXyARnNke9nZzVCzV
Zwlj9lgkBz40glZcnrVN4c3FxfY2KtE4UCDsRqJWdAc+/IWo2spTTUF4KWGAoSav
vFHWTj9xeH/4JTUI9oPAEtazP877O5eCysvez5/IZqWM0Qn2WsivV9azlVGqPHmU
KxQTRYRFi0b9EXHJrcZP6eE8lcj97kUfj3a+oGqF4cDR3f5k6PFRT1delBrxYNLr
gD66eYe22zVq75T1JHtgAdn4KAd5fsXGBUX6BCUXd+BlZyEYhgW5bPvhQYgmUptF
k0uM9GQu+u/gfW3IszJRQZWbsIMztMBfqCzQMyhZPeMg/C8qh1tahYGN2nvU9u6F
LiOCyq6XmYbdMy6hrPXE+oYAkkdxS4on11qIwOx61LEj2kO6M9zBBuZoC+OxWR/K
M4QIuHGpFpN/dDLhy3+89yKEERkHj4MHb4n6u1iqsMWgAT2vnBC6QkJRgeRUS24X
k5oYMF6WaOvp6cf9S7o9oxAilyytLdMAWn7QZvyrsjImpxXYe/+/j1kj0eYe/U9k
LV187yBgv87/aWUtGb1rwKTVKifCjf9EUlgDbkRsBn0TB9OOVKITzeLQsm1Sm4r0
dV7BHbMq6Phh6jnP5NMd98QSuftyJ+tynM4t6mQOnv7P3aSpniMHG4/CIW1EciOO
rW0UsShxPe/fBEUAVqJbWhM1/Ap2hDuB3T6d3ZE56tOhBoq1bydb2zklMvf8Slfb
5FCEWfGVDwSh/d0HJUqSbQWu8/c1QdsXzp0Tq3wARo+RuLdrQFlYd+iKIj5kMPBf
3e8Ss/OYWJFKr8w6udcGYP34tj8X+OycTqgKX6hrnOBGia7o8Ln0y1EBQoIYKXkM
a3vN5kEp7ENIaF+XhU9jllGiu6H7gv4qDUZajPqdzL9gFcdI9mLyfFlLLFk6iGNu
G1pKBs2OG7mScbQU1gFN91rOWzTNTLqNXvB1BdxdlCKoMiORrLYxSj+KnVC+oPMm
LKlVwHhaQ7JnITrT9AM7LPx9BAe2dgKc0kpSHRR+amqlKZF8HRvpuEJviMuKoyVz
+4GXyHy7HQDmTQVylnMN3AmBEuOmip7gc8fk4Og0BKAN22EpBBU+hGnco3WqHVqh
kRPd91WuaxKwgoK/Gj68Sy7cGr8TRvvdOokh7M1YEoAVyRFolJ4+5HIyMVTgVpve
C9/gSw2ap0dBn2pZY31qlOkh6R3VqZom8NF4aBDF5UE1U4sFoYtyXlBmkf4k/Gfj
lFs8anz+YHcpAUA5SwLFm7PGA+N/Y+V8x4oKold8SO9dekoXu1bjJvJ7+aC/6G3Z
CboGbdOLly5i6xfHi3TN0eahokrrFWGm7z5Qg+D+I80qx5O+T8P1aSbH3QlLQexB
6WhBx3eJSda1bBqDGhX8zhmg/7MS39yxPuBHfmWokm7N2WQC2amdeXV5jbJAVasl
tm3G0GkEhf7GcqxYjb7/WYsr8FGwRJlGayrWSzWgBVfS9XWbMNdpcsQotSdnUGRn
HsbsSbGv6v4bL2H3PiL2i9qyUW3xtIznCzVKPSKNLDUjZrI6B+XcHWHwsbCvNqZ6
0jJO+6dmRcSvxOSees6HwEJ8czRTVQoR30EVtRiu5S+6VLHDmhmI5gMQguwx+s53
b1yCuIVqK25vaGxBOE+KZ80jzHLhGLCiuvN0GA9g4D/OdDLOEMJeq2v4/0w7Gzir
SsDIsP2WIlfNmkiqbBoOBw5g7ZMLjUIpZA7q7xIME2IzVUzUt58yQfhFMuq7JhYO
BjoHtQCQjstigz6ttojBnbk4EpGiS5U7ekZZCn70p5KcHxuKjmp6wcZEULvWGoWg
3oeXkIk2Wx/bDI8dSe9PgiP4zVE2K4fjOgVrQTgUnPSxpj9zqnjogZEblXB7Zohx
JqAeVPaLY8XhVESCL+7Tv0MehFaxo6kfnnYc8+WoOcR/hvMTm0spuoC37kF45XNF
/Ij7JuVqHXPg/8fTlJy6iOxfJR3jByVMrS8Pw5uDhpnWZ4lfrxVOmdYW+rs1wkqh
qrCtQ97bpZ1RPrzRAG6iDYrWZc6mU58GlI5uV3oKSz1enSQnpM4W7nAAOYmXO5rV
BFz8wMRcEpVKhDq+vjP/jrVYaZ8q+YY480ApBFFX7TxirFDUVFm62kqu07rq84eM
+yN9JWbGZRb7fGYmbjVPhjYxmmNSN23EvgoDyw/tumOQefTErTZt5Tld/PG30LX3
GEFf7w04kCAvXzmXJ1OHhKBO18I1sODSsNN2zKpUbgQ2XdiyqdLgllG20nr8+Fbz
6fDrSCt64uVCJGHBF2o9SWlW/kK1+a+0KbGxu3wr8o3ONE79BZ8Iugtieg8HgkSK
TeQdYzgRASzb7JPF7YybO1SJA3OkuT69lrr5NBw/gO3s1A+68TNikleuNb3KTNOB
3l19kwxv0e3TFHkSaM2rywmKKkr+HQ2yrhMm8VTk7ffevRfTOYQqF8XUhdmbaBoK
Hvq6Zl1UtSQPZTAcxd6eB4sK8uisqFzVQdnr1xkxB1n2H+ds5+2M6eYH4dzxTXVX
OGADxPff8rScqLW2ClGZTaS3OztRt/VnznIXDmou5moX55iiEdF9iyxXGQHjvKg/
SBoUrYkZCxaIOcdmHvSM1vBhAtaTGx4/zqGKDjHJKMQLdDE5eDIujrcBDrtXCB5d
vEmfVY3iffjvx0Yv2GYbutOKa50TSSrRQdINrnrUCuUTgytCM6e0DsppIVHaj+9I
ZLwfb8lbzn22R1Wr9vKwnb+5l/GK7cw5a6283555H+zvS7CVvjai6HbfvATww2sF
63g5aFTw5evAFbmy3z7bjtixe4XcOzog6SmThLmEZdE6SitPHn5A8cGKgKN8ejag
8QA3JdOnAKJUWByklbeVFqm/oTd2jW9XemBKxm3ymhWe9plM8PwdHd42ML4KQnsR
wCW5Pr+d4hMntwh/5VXBT2VwItZs5kNFXHF0hT2jVaTUwluA2Vl9yof3ooc/Lzjs
7oxuIqj2a50fezbPu3E0eCSdwnEi9MgxLgxdecXDwMC5ZOh5UITwlOEgLpFIBAsn
U1dAOIeEseReHIlQMX8Bs5st6tAg/j+r2DheIPiTPO3b9IgfvgnrZOKu+HcnDAby
ub0VjHNjhVnSuhvc3QXuQzsOi5Oh5v6dfEV6pTaFILH3TbRF6Lu23dSGi5fO/tgz
0CHOjWYRTdSzM8q/vnlh8Potj8zZhU9MRrihxI+ugBRjE6MY9Dzhddg13oI0Zo5W
vJCKErk6yf2GCHAXt9KrytzbEsvycu/EFkUTrIBl5Xg5lFrBYsLAwEqNVj1zzOCZ
ISIFI1wQArnDSEXwAVhBRGU0JDT95wwC50SqUyO8Gf7OfyI9EWl7gxXmteFllw4H
98KH5AfSva0VLqupqknDDgoghg0wA7CCEsR8ssWsQf5UKLrqPt+++1lGTngpcwyd
2ayjw2TCd3NJEyZcnZmO6fVZGcejN5U3PrSrpbIUHTdBOT/rHnZxaowJao+OEeBH
xtOFj+LAfCAqw5njEkk6YO/JXL/llJ3xBeiAzA97ao+0OPvweqRPf+KzLatWLySZ
M9KdYHC38LLH5s1Y/WRa5R+TuCalfQYmcv2+laXrdOq3n64IxLzm5JLtvMzApzBw
Io/iypjfukfhUWeRPUjuXT22DKKu8hbhBJgrVXTP20Tydw9pc0MStA+qzc7IrxfP
whWFmcBvm548GJ+3wqradWhDNnBjegd09aWR2+mAVmMDu+W9Mmz3dYiNIuTyTRNw
mVGM3jPzoK4y92BpNWr7R7db5YbP1229jKdvHVAl0EnuOj+4Do7b1/jxEN29qKwq
xE/QkatwC159AfGF6hXuJLsUYx/RnnupWVmHBFScTB5zIYedIOQS0Xbt2oawK9vB
qa2JiRB1xPgWmVlF7dRg8VAx450NhXpDYvpeacrOAR8/PdWaY0DLhlQXmY1cfZKV
2k6xWTBx63n6grotG5O/FMBcsMGcr28Z1qRal3FXVOwM91xZvFyThpstTJSIKBhT
m4eVtFC0ZUFYYSsuQh+c4yza4No0dgUcBEF8F9leDpexmYFdNWveTNaU3+e+z49t
mFwLWi7+6KjHYJllRn5A8d40YAyc+uqNNif54f5kxvXYPEHuKGA0VN9dBQmYl9XU
vAc2X0vnJJliR0irL/XKuJjj5RutKjf9Iqw441eoHZqMqhd6xMFtZXwV78hFcilX
vwfxCg0EUyyBbw52TMamPC2haB9C9RlMltQiP3qrLorUO4X9J8nMSTIFOJemgL7p
K+37ezaW1m+SFBwU4nEJRq4xmx18iXPOJ4OpfQSYdnZPYw8Ase9HN3qIG2518/JZ
FO6eai+5QJLS+aKI1UcyBRJUbH8ZPAOerF8SOIaHlCPoxAEcRa1AOHEC1RBp/UqV
Q3MpiEGuaNlNQOlLMt7LOwmZOmPxUB4AKtQYPh+XFljaiSghjC/14ihSZyPr9ZyS
RcYOQsc6xHrMG7gGmsYAN6NbQgsamXg7zGiAlvKFBPbebFmNSbmNWaiyaocOFfXl
a98vp6n+kam3dFYLk0Y69t8evhhL/xp2jqiLf2+He7Qnm9g2IHQDzN9JjJOcgim8
/I7X7Psyb0hMJhZa0J3BWz5MLAsBeZePy9bDCC3jKXQe6cw6bSLVz2lbx359ov31
3nLYnlt+53HAAVGbUNGlH1howrR3uz6dMYNJRFq78G4RGoHUb0KyffsZjJzOZEMm
GQWQvxar+9KC3e9ywxjVWhG1jB6jVVvgVC0ttwyAKW35/sJEaFHmf/dIk5aHB7ZP
vIZjCtxmAt9Or04SRlDISm2qsZZAigEHI5v//GBGhmBPjR/0Cc//9/fZrhXaSk1X
1x1WvV3JviBqIe6mfIPyrgbH2Mj+0+JWFHWF750aObQvT3EiEc254pwrHoAZowwR
RgNz7BP80eLODauCBQAfH5UniVutMr9csnZ4rwX6Pb4jNisFTdJfNpoxBqbLXkyh
zxDdFEMGFxjHAVYPdo6/3SKMA8IhsLzV8xZn7TwwwL5osfuwyXHu/pxn4MyIkFfk
ABuanWeFLxYTMfUgHqDdvY6B5aJWikT3uKdcXsB4MZ+gDYS7YSAx++KUHyL5C7Ay
8MOcih5xvXuI19Esb5i52QfKRyonx4DLXAZP7zwyaq0HRqg5OMGlOnj3fc08CVQ0
vGSjw9NhIUG+CmYbeiiVXCSvZtJw5DbvRWdTG1C4r0k0ZkiWBgfPPovTCaT5F8jW
fQD4nrzvnRtSml012B8XkdcdErmB0phKbEs5KNWG1b7jQaFYTwX2qH9ifOzpMSgk
K3dTrrLHzEp5NORk2TvRK4O2I4zFfwS7ydnkU7lUAqY8UNKi5jf8wH3npBdUkdUm
jTCbkVp+Jj3hufUs6ElxsIfBXvDyplqiB3S0/cQCy0CkwC3NpcqPJDHwDSgPAxBS
8juA+jK9GdDob4ReBYGELVK06JflrQ2iX1wbvbMD7w1Zj5N+zK48+WEjWd697kAs
rJxq12N6s02kLR1HKzw2AJ2pHIs0QMYX8yqsOboQ49t+Sf/R/cEm7z5bMIRUKMCf
Yn2heIX2TYgP5OSbDfQ2TQcR7ILJMy12kXMwbdR2906aANHLMCMRaYZAV3hQLbwa
RTgBs63LN2qJtVy7dRpG/rzamsimBG7XWI/u1g0FI9ZwhA3VamEM8YP3Q1WEyNWg
w6ViqBQcd+9wXYSWrCwN/Wa911uhIfRbVGdCdjlJ780+TmMlXcHczd0a3te6QpST
2U0PPvZUodxsoRKdWZV+//vKk8L1lFHb1xSwoO3w7HEj0YWC55bOT4FKtbBaj7nY
bRUOfdO4CC4aG5l5xM6UzdDPtmWpUpNpRDvWopWrp0joYSid1a6yyIUOULpzpCPq
Hxk9OEfCUAf/XfI3KZrqFVSRJA6DdMXZASnhIz6U9gPMCayER1W1cR9jUpqqPztt
Tj9CyuPmTx7+0l/eSIB1voa9uJzrufBSL+7L+/kG13r7MO87ANB02Sdy6rbqi55l
yoeSlHr7/fOPON9M9IQLPYLSTAry+vJjVf80Pt5tkqGsr2CzT8iP+1fXxc5SCRRv
HLvXCLtI55pMFElU5F3MX6U3PTHbqMiOJl8ZQi6OXhTPBC+sqCJVzqIe7edZ7b/y
9cmZr0SZ3LrcOSa9MioX7s5vJrZPYD1rqK3B5cMV85qRaFVukc9iFaFOLhReqvVF
oGrX8twCX1DgHNEwrLrDdpiIJ/Fy84nWdfiCv3NJ/ZXTtOgZ2FEXH8L/naKqLWHL
08DZO0cw1+HuknkgfBBfn6xUg+nhI5PJvv+lIWbsqbie4r98r6zzta+RKGcmM6NJ
kcydZkJz4IBbhNPn/UB8+6tjvq231oG+6I5H4LvhNTEToepGf+D8fGYBJDgYjgzp
U3IyiKfvP4Z6a32Ha2zkFg9Ej/jeEAx5OdvBuvYq5rqNnX0XmeIH7ma3PoRlquuF
NsD24/g8hXX6a/vgAyBJ8SfsQ3eHmSFDHKR7wdbcNg9bYeFlujuCmoVMAIbF1HLo
Ti1i+TOrXTsctmto537cnv44FlCD11JPGXKo3YOl/6ot5gqumFVmrwukEey7ln76
S6bTKi525eGfVTkDiOMuMvpy8PUKylHRq/3LjP+PeIoJA0wCjWoKOkZ+dSEvgwUT
MzritS4pa7Eq3qM6MZcUMec6pmIqG7BiFoan/j/ZDOLvkCoCYmE4IdiIt0BszWEl
pu1vdGTyomyVEdtPm0hz9ggeFkmUcDEYkI0hLN8RTsIj9PGA9hc8fyM7v9tQ9EBB
fa0+18wipKPt/ONse08o6AMZK6jpaNa8ZlMK9JoaDHveZbHbPTKHxAj+6Qt7aP6S
K6Dd551pylxkZp4G0Gsu6qxbGGYkfjV7d0Qryyp6MwcHGKOCNpHJyvOMqHbOdbZQ
cRqdjGJU+mVfTBs1qYB6OZIAsMkjimQbH6HPO7n1smYt2qBP7EPyYakrpg8R17t2
1wGTFbkeXoPvmz4uXPwWWVrEXG4lJr7QG6F6ppDviiQ3FFHvhJavyQ3OZpEt9H+H
m4fnL4ajqeartlYJx2J4hubnnX69XWmxuSrPZs0h0qbI9yTlialGZqDt+PQEHg3a
fo54TD9vSsaNjCNidBmIlgWGO+40Itx/+rbXEEJuZAHhHVRwYBLQPm4+L0aITP8w
xtWUXC6VP7iOnmxTMVAIGr9rT/kISoUaE1CZxdssUaOazZzcVl7ZTK2v/vvjHE64
eu9oeWjVQciOs9Pv//ZCAzU+0iksstGg+RmBgRWBJ5aWesEP99A+r8Nl2zIVjxmC
VhKOr0IuLuPVhvTo6Ck/YqEA8qMhNOohEZ3u2kzwTaskftPQ3Z8R1f1Dw7LAQ/qE
8swBkhA4wL7sX58mXJMUbrvX7zeWgaXteEULLPcJjVBsXVHVkmEaTofWp2bEksB2
eOEcbZo0c6he9xtqPRKGJBKXaaOHGO4rH3N7uJeKv9CUF+iELTbqUwqHXsNhDju+
ea5oB/1XuOvuYPATpGgxtIRxYFaezRXdCxMgOq3YDHLXk1gNWDiKdDbhN03fsDSA
bhOMVI0mQH6yB88G+pKJsT5AF0yjqPulCJttdNM6ltI4ol3Ec/2D3ZE+/IWSwpxs
5gkqGQIbn34y8R/Lj0Wsm+VKcGmCXNHlx553wSxQ05KdyeppHal1cVtwlNxoFmqQ
sJqx/yxN7Fz+/flqYSSKnmifPoREBJvpmUBJ+L2GnR46NmKBhX2AnHLZyaFmRQd1
mC8ouXHW+M4yfcgrA+kQNjevbSWVUhibgrnV0SE84CRSVPCeJb4rQ6GTiFeR/5D2
VqN95PNtfZ+fNMHEIQSgyBVqe+EppWUmNBpcY53pCiwr8DcKbymCiRWrGGmCIwVT
+GvLXheVo/xrr4ya4iDbYTA22vLzda9MweFmaCz6TuiBKdNRG8rsxHRW56Rv5JkH
I2cVEDMN6dnOjHv2ZkI3IEQHw3P9m1+1G7zQcg1rkbgyRspgCyCfMN2Hl9Psrfl2
pcdfACwQCS7N9+gJ1NcTcKAfnDprYuLRLO3GTSh3D9565rEhnTOpLZWYXWLTsuEe
+sX49wP/PxAki2DKNVcVS8sX17MtDzYEmysCrxSyIop0u7wwp1EhG5Axg4d3o72T
6SOYoGKoHY8R1hYEm6ERzfTM9641a7U8yd1prCwTqiA9sITsyiE+VUwKFeQDpsLb
oawhATVvX4+Sr425pVvvdTHTRWLI6wswj6HzonPDyepEWeEv19QapTRicM45hT4U
T/JfE8EBN3GXQF/QHx0qZCx260Nit01GiZY9EmswbgjzgetjbhG3+A2QCW68tEAe
wfXB4QJF3sZUxmDsAC01Z1BtHvr+Np5ym5ELtxuCxIL1t/f5iRZ+YP48UQLrvIof
Z8i2ufcaVB59VLrCuexfXg6tRLWf21gmuIBdB4VZzNRt0mUb/Ff7cv+4pmzPmQGH
hz4rQ4aaX0B7x0wN1pCixB0bv9hcYdokS2ME9889FRt62lwsH/EeAMF3CgkHylZ3
kySaw9SUOXqdWhPUuYIbDYEao6WW+4oSWOSnseXrxEum0UJng0GqSTtewVSi3R23
vqQs2l9LVPJBTdH29jnWQ86CIDOjFndduhxtnRs9aittM2wsaqiCPOde3cGTIp6k
IFcjDYL+7wKrpuuuXdUQvpJvgs4DdkKzaLje0yiapkXdoIWIRVpNFOjJlIo0JKOF
OSLo8ilYmCJT/xmM05LGgTqCEYdp0EANr+xMrnoCC0oxl0IFUXNE2tjC/TQyxDYH
y7Yeww+jGGRxXLet7OINUwjmEK8IPEnr8CBoUHrjzI542r9U3SI0IQUY8FfSzxAH
lJBHMSxGDbKuK0JdyAMfEGDWFaPzijipA8KZ+SMraPBgSUBsWHRFsb58OyHsQBXH
Fe+QgK3k8Io0Kn3wN6wLDGlydJGVfbVl4tpSoSGgJIHLv2yezwj+VwyR+tsYL5va
VbfSpNYUcGBr62z4vv+lU2o10j2c5WZnrbGez5/DuSpGzx2EMS1HXoX9kJbBXbnD
wvZh0ryPV9Bs3woupbHJWWuEfBs56qu3pcKBqTIcd1P+gtB2/NTdUDeLWj5c8WCT
ZKRQQyeFCAkGJ7BhplYlDIQWtIifWPT9nUBORAjBhHr7deAbCYm+VUrLcrfxK7gt
QitxMsXgYq6v9TjwDMT4xw65kwE/9MT1j/gnUWr2KhAZ/o5ilO7gutIwdIiRpsZd
f2o+nXREosLBhDBvNTvJrgvnYmYt2y6gCQIkwFmhw66pttjjcrZYX1xedtizyrg8
7wgwRcYxsgdNYqYyW3el1YKI3Ca8/00auR7OxrVEK3TC/OxWf95VpE94TeIpb517
Yxu25aEhnbtwoAc3RMsQjpUx/IDlj3xkf/AsmISI2EgNejhACFgput9YNwr12MUY
aryUwecUdYaZSavo38K3PHfRm8/enri9s7PZJ9W80mKnX94//ElhXWmU2pc2N3Tt
5P/qxnsaYeBrrYP2dqkPp1dpX1uj3xzOPG60R+OJ79w3JyZZDq6cFtvibLqRhZ00
M8owCtc47LfLGDUc1/Dba/RqJmqe3IH17L0QEE6NXznPP6SjA1gIZYMIYuj34DOU
eAVvIp4NCCIv1xuxflODZZS5K8CsEKmBd1+bnDri3dEKUgpQNxTbYn//JV+Vvi5C
YOlar6UmqxhQxkuq2lXl/USxBkh3uBAa9CGWYe9wIg6OUv0JZvOucwmTxx0u+Uhn
DyMymNHO2CmdiyQnPZiTS85FoC9i68Zl26BoI8Fw95Yo1GgXrWPS9H+KNkMKQDmF
/0k1mXRZkn0OUfWDjULQHC8Eog5vqYHQeMvm+0JaEvXveBmAy76nVLk3rYuo1g4a
hKmLtme7/l6zm5AKjooZC7KKaG+T2C9tOdwgTvL5RykXVJOAgL8nqbKD1pE16swo
/m3rIDrb+93YIFMLTtvmGsJsUqOK0hbrMMdM5BLIgzypBtCXZ20g5tbaoOWl4ir6
J7pbBO316HzHVfdnJoTXh8fV4q6nBUYKZ6hpFxwwKbVQFEXfwYyQpr0/aONxHmz0
Hv6Ih8lxs0U83TR/iNwHlEGEz6XOQ1Haj7h0aHDjFXViI9/rGStEoBJv529eRHjU
DcCnJFRsWiVdfzwFlArg1EEi8Nw2S6BwvBIwNeKAU55BvXRQEyW8R2qYjMSo9kK0
XxG1hU3oPrAbJesH9OanAm8YsiHLTlscSQKHyYyb4BdQY6uhX+nxznXup6iyS/ub
bE1+Ru8ZkyogqOKvIUFaSD8Wb4Ucf4fCm8rP5DVGMEDhmOiCwxpcSpgAmR+NIzty
iGW38AzpJuJyWjjGFhAQ9wf1Cu7GPaar6klViZ+nki7EhaDHqs/hFnOPQAZiZeQj
pvd6nxFnWu77FisVhDZPvmfRz1yM1lxW30pUJBE5gHzmhnN4WWfI9C0jxjg2larX
sr0Kk8TsN8sbkv8ZDTZI9EuPCYtjFyQOH+Mqsygnw7gx6fy5pHRa/+gKhSGZN61E
58cEj64sBOqF7/GGhtPx2qhv+XD/YayTJEikF65dd83INLtC9mfRxKzYzP474mKN
/j6UwtFtiPrZhwuQtsURjTe+iQReLCjVnEqWJ4qrFWRed/gkMGZKezSoOMyV55ZQ
axsvAqrq2Bca3b1dJCu/GZQfag1SBu3X5CZvTh0UUqlaDrl7RRXYpwXTWDfdvyYT
D/RJVLoLIeTUO101kl+q1zUDnl5INX1b+8AK97sJAU0O5lweVYod65btvm6zj84F
IDRwH1Qo/ANq7bOu8Smom8jaoNvvX8RVrYun+pMylZ7409mUlpIkjuviduxc1wsT
Fr5OyG5fujrbtogJaptj0L9W6cHWyVbovZUJ3pgyeZ9HcgabY2lJQEPCTQkkQJ9R
++2csNHQGFTFe89wOUfj1AZDkt6KHTH08S6Cy/QGK+H83FGozBuNhC6wScGdYs2q
R92WCEeSr2DjUwTqHBzTVzv2PJz6b2pm7Mdur+Zhz0bRRvayXCdGIPCfyh5c+b5r
ZjVlOgJzQ9S58cPlSyz4UIlYQ2goa0NP7HMzlAE0HySOPm4zWjttzzv331NOUTd9
nUIyx4BYSVir4lmefWsvT2oqJq+vj5HDzkADF33Xmk8ak3wZY0Xg6lpMbRZ3qcZA
HjYjXIZyj2w2aaG+J7aeUnfhORAx7As49B/r0trl54uBRqj1AqEC+OT06YP/OuRK
w4vTfG1ilzMa7zgx6RZTUzLERD0uIlyNwS0eTsiVU2GcNOAwkIM28wu3CHRjseI8
hCBfXSZqqIADlaIJfP6nlpHfI9BWcDez2Gq30i1P6DVZwbE8SyXGDYFkobedUsZG
cfTl2QksUU7gjqZRI5C/4hC6+jZJxO+JkFgfdGZ6OqW4YssDkw9MeWcP/hhWziev
tJ+PdhMnX+PqVdHCiclvq7Psuu3Lbj07KLyyRkkjO09DqQhf6SbeHl1n7qSIDI6F
EKr9Q3DDDshmGPPy/N9C7SwEtL/06tpzakC5hkPn7iBY2WbtpFyW5Ua2HbxX+Rqy
MAUUNZDas8s+xcquVrvzIpWVCwUdOo9snymcmSEs2U+ilHzb268x13akXRxkplw+
2XRPgJE647fxkHqyuAJNYhw11Xt9uyd+i0CAJFdwMyVLKETfudfHWkrSqzGbtpIz
iqtKxi5PCuy3JfMXhrwWhMzqQwRmSwt/zX9XQICdP0cidmQE0QDxJnMt/gcpKwy9
cGQ0bCsdHfb3Dk8xhty4QV7MC/MggkIO/NmMUCiAM3nNoWKfADjE6i4zMVeXF3Sf
St8580bC9qR7I6pvZt9C5ySeLCrP3EiGvl9jkzE0yTvvj5uB9dtCPxIwQ4RNudrn
cFynhlqFkiuYs+3xdht9Fp0T9gNNNxEAYi4+zooinfhiB/2oIQJ2cKAYY7dHLif9
ckNHqq8NISVswrEWICYdkkJLIdaFP2yGmiR4C9ubdUXZcoA7h9iRKYrYOTnqbsqi
hJc0Hk2quEBo4kOLlcQpIX8Ohz3KFRV6USHP1B0Vx0Z1Kc1ju2SqSE3Oe8MWasjF
byVahFV8QtjMEn1C4PECvB6haMINuwP3IuHalQjvWjMpxp1M7yw9U85yx92IVYzd
PLOrUBckURXP1yKoD3sZ7KU0ekRW7W2BrEawayEMd2vkPoPZvfcNx99MM9BVXHx9
bS07L/SdmKIb+HB4hDblnVSPi04APpd1cPaJ+ybAF7xmeMy4lkMi4B8+KEUU9Ufh
ajHMfNL6V+JcfWp7dE9nv58/YlR2994/EA5lJ4g3Qc4Ose7uFE+NQ54DVL2MGmZ/
I21oVGf0ziwXZLrowffaRZJ4RUcDYPF32slXsmZNpKOIQNG2QF/ymUuffP763tAt
qUk6GMUOg68wmBehQQ49aCSeEZpM+0T7Us1j2vh4J5yeklMH/J0RaydXs3dRRxCd
mrTwkQbWjX9wvHukv03Ca2aS972YQNpG3pnF4bBCmNrpeIQZE8DjYvRKjU7Gp/Sh
neFlGyP2MQ6Z8qcd0hVYGIk6lpjjLSpFq9QJqZx0oL2olPP0cWP4xQ0bfZiZosMM
5Js931pzGm3kEb9RhxqRbvsfP+ZbbXQeva6bILtiuqD18eCyLn2wtmIeaV5h8rd3
i31iMW5mHuFDVkg8s0UduVlPAWmngLHHwu2zM8be2AoEq3OiO/ehequZX7nht3sS
PIBQyYDMhrEDVdU04TlvGo95uoOnfKczWAWzXAcHrkWJF+1AcNGUFU84cAsXpZY5
f0O45+b0gDFLWrHE48MVAgvLYiWAUSS15hs1M2l1ilWm0v82Xystt/TOdYROVdM+
BisRu/Sr7n42Y8B9o93romQTyEn08zj779L4Bu8cIBftIgrqKCrRIskZeBFhp2dR
uuCyLY/HumcCFnbJ5BDk3yKar82SdZg90vSntKXh/rZpGOoPLg3eUsvSbHu4Kpzo
PK8CYusdOGZc/6T50CexAHY734W0pxZiZvLhQxEnMRIVIfn/z1ZAddKlqfwPWH40
R8dRTFfUg5x+LMwZwp4/lnaum+R72DUwKw5vTPMuSHxTJBmj521Slh72Rzmpa0AG
hwYoI1eHWhfBUcTvFwRnCriqFOPuFCdsgBfW2/CS/cH9r2sReHOXoAyO08R+2DsA
ARqJs83xJSJDU39AUzejPod7KxsaXqFyrSwHbZ+RR6tcRXj8yZE0mpSpkUaMkLXp
IQTPgkbNzkHPjzSAcXPKLUQJI6hZRpMtqVjaAsP/2tG/5dtIeL2g5/TxaAUbowp3
6a/+V6gLW+lSrEEw/bLbMcSOMbc1eyf5HjjKWyPlLx9EpNHoODdgWiiknrJQHbeA
FocRBbakrQxvKxf9nqDxcEUm7ytNAoHGljkZDPlofBcOs7rRj9Jq18dJ89glh5GU
rIR8Sy9QCwlcivXa80B8j2Htx/93fSVMyCXyY7Sm8QcTLIz3aVuY+YFjh3eZiaBv
uL49RZ4ju/0pqSN+Pn0NU+BHetBFpVNH8/maj7spDjPmHVNEELz2dHONVzH+itkF
Tj1zcfGBVrdwBWM13GNcPDz7EXUyErjnktYF4Zx6iMCkU9VQgwXqcWmS7b2KlpuE
Xd3oDLLUP33FqHodZR02yrFOD1+ybul+GPAepwX+jJarVuIgFDmPuCV4pdOh1z8Y
PB5iLfBzT8CXNi93B4G1r2hiHbB7D+WabQlU2g4miWW6LYMBB0zI83ip+1xcEPco
/XV/ptRoZCBnTmTPBK4turc8IVjFonc9tWV7Ts6ERfvMeINyzWtMUBAHJJRBhbl9
TEkIITOUbH0k61nwkxDO8goq03VdMipZD07ZQSIAKjtbA6cbgJi7o35R8c8U5X78
HCR7AfB5qcZGPLt6NjiyY5F0LO/KHFYr5SAFovxs4J+mdTPVe03LIg/D94r0XaZE
+9G/HTn5DPIPoAHbJuY3KwQItKfUNT8ZgCHtQxkv3q8xgr1wl7JLjpqIkmBKiJ/A
Z9Wy4fE8nwGIu1hfy1NaOBOFQEAmb/K0u+DWO5vQ0H53cRpV+FWpUBSngF9CYsX6
M9t76oQAfXpbIdkB/fisOWL2ktHhBcXHU/5/F6WiB61K6h03sChq3mt+u8h2/ayi
PQs/kpkb8RWIwVWF7VoadQyboKpSDNCq05e22n7PdRAqncFDut08VVR4oJ+XlVdR
GQHieiUjWCVIVuc8TjMOrLvu5lJnnyZYg5eWmxAx/03tQULe2bcpv401LOFWPLwg
WVnOFoTd8MdeTchqq5lbKgIajq3NlA/1p91FYMptnFYbXqrwSovI2gAt4VeDlX5j
+Ocw+QZNhLKH4cmrVZE/qZNzY99L4i6v8OF1DEpP7jj8aLuJV9ZYsCuo+kWDJG3E
kVGJ9pIYtmUUT4d9P7ifyuxLvnW6YlhSLIaMudJN2lgN5ry+46F6RyfQdwMuc2bI
FPR7zvT5xnoeyS0NP8tDE/fojAL5BCtx1SYlMva2WD25aFHQKTszPAnpnw7yAePR
uagtO4ooV6BBc1T/tLQritQ75ofrAyJilYSFgGmK/sIFx73WYlULAjcmjremsX9r
utUpEu9DZ4eU+OrR5BsBoDCB92uuFgQL/MIAHRDl20hjlVXgtllnNZwfLNFHLR2Z
iCPn6d3MA27ERIjUKeJx1sv6PgtX2nuPU0imPuglEQSuCa3Xmq1hPvXBJkMniQ4e
smH7dwvEcGME5GvlPJrclnpC2i5dPSaGUYsC0gB/n3FSCGF9mqwFzTvudlRBtPBv
XPv5eL3cjRuMVrfkhJU5vxJWAem+9/HtrzVb+pFT1iLw8BeAk7PR8cOkONQdwxdu
+DcpiR35jCQV0L3Hln9PrWKdIiszLFIOGDt9Anb+4gDwj06fKTFGO1OyhiZtRQB9
H5KD512cmWrccys4++AiAEBNLV5KBlOLdAEERmd4cvjmV/OXB73BrtRH/gLaOHwX
xRBnmXJJ4ZkRIQLhBP+wp1JraoRHzLpm2GchDMciil9msVjd+S5U5aLuvTRDVDBJ
qqufACdIJ/mF2xqVHLt4PtDzZggy4/gwFwS71MeNvxCXOFxX1cRBdCrnnnCZhLxF
1Uz8WaKBCaHzdLVBi0E5EbdvGEl6ovTiEKCLpoogJ/0LKC7VJ2l4THpcDc6Gg20E
0gxYFXsnzkSjeufMt1uNgZ8MDCJBzQBPQNPA79YwM2BpYLl03qO0fWrj8LxEFpr8
QRr/hRDRnBn4MJluOpTEY74O2B00EEZLKIFjz2loT8Po3CFKSaUGwzhT1PShpLpa
4+huzNgDEfe3atB/jg0iiUsXzozTidHv/CrfDsOjcpJtKToBiQqIjosuU1rk30Hr
prrYvqJXrOaBPHcmyqb9/a4VzdSvi61IEYGrgNx0wQIa9jsluXcDtGoe2BSQWfkY
R9/s0EKHs41zCpUVeQvTq39jdhYOFBuT305FzACWFuiFyTioJWk1IK+TMQY0NnOA
Ig6nHUyZtTknaVfsiCymHYfgpQcQqhJWISlZyXtUSbK9moZYDvCT9Sb4xNdkUrqb
JL6tcJy7xTlJvTfsuAheVsHuoJVa07VDmh9o/TZCnwS+fM2cjqD/1+8YpzT2WBHZ
/w+geXEPNIli5TG83KOZiYIt5TTw4uO+ktvVU/9iY7hAnhg4vip5orvJDEUOFVk+
c8tntkEWgTVxpA8ARyeTRvUMn/1HPzfjeWT8WZNaaMQqT83wJyD5oug8hvMzqNBn
ZCT+5buSSUpDPKq0KaRXVps+u/bF0yZigzAPNrKxQQinDhgf+SLyzLrLB26brsiK
QFgI83a5IFQMa3urnkcSdLt3dFQXxn4Dr49iFe1Hs7Hc5adWUQ2ZJbgWltFOzJyH
4bAtmV7R8DYVRr4eceCPhb6AKO4Yj4zbqa6E+zxxHHhaYNA80vdUW3/+zOryeaoZ
KxDs+88xGDhz3EFhfWB00BWz8bhIC9y9SXfov/RyiIZb3cKwtWPqEnxl8pDeI/eN
tswgNBmxoqLymM/peu/ATn1CJHQwgJ7I85sRJ5WNtTHing55gZiJoRh30ues8+zj
0k9jyj2D6vgHKIhDPEIZfEhKncpwgnzQEJwZkHgy9OrIM2iVma1Ozt8JeMooQy7D
nGfzERhu6lsYvsKETo4I2wJjtsHHA8eXbB0bHxYOBE6/siQeqPlAD+cvNbBZhl3W
JuLaEv0DjQgJeh84cXBXW9byGmaC0Z/7Jzzjg5BdJQkDOghL7tqR/LL74I6w6lpm
NvOBrqo9VbleLkziktVQEtsdBlRSghFIImlvTmZiz0cXl4af9NudATYe3ed2u7N5
PLc3+8T7QfhhybkblCTOX71L9h+F8dNSvDMUOIIa7ihVew9MQgOd9pmEF67Lqj0a
9hrkEllNGvnlIQyky7VIKTgx1r9WVUIM+N7LFyOux4Su0QUwxvxgvrF8AC2MHgBs
+6oHnWGzTkLRMdrXZWvz05W3VVtfcbc0QxYl0NHXPT/ncOzzMzB2W5EHkxBE4TSH
XEbUKuETl3ncQF+nnSdg0eXej8nqHT7hJElJLDoxtIVqi4ex+lkjX/zmKfSBd/i5
df8TEp4crVRdGR3Nm9khknp6SLmwe19bC/i355CWt2HuIY3WwnGVY56Jg2/NlZh0
blu49rjoZ3lCZm/3nDVrfFwTE/yFTBzlVdNmGpFRCLeXSQnhLK8KzbOat+HUun63
1Wsl5EO2PXiYTPgW7f/XlgfwujA37vVHU1z3JABIgGeyRnUBAUClgdVHDNAFIhZ+
kTeZx80jk3fTdXSBGX4tUI0enE9M++3+UwCjKHvRKI+spHwxiiQLokuhBPSTtZSp
I0vnpkrHcUfHU7FZsEA8es/tn4HHIlVbmNSPPY58XO9SQrsVhBBKqeXv626ZHuEb
+Q4P3CPsAu6kA/YtczIS+Ih5Q4a6NYaa79rSlTXfBlVz5NxajhUYKs5YFtIjiAPK
e1O4bijk5sgmhgP3aNDwxhubjDutRvzStgLSsoXDIro2CFfLwL1g8OmNEX/nRhky
upPfnCUq8sTtXKeAO2i1htzKtXVojfCiIMhdnH9OvOjyFf/pUD8g7piobCCwf/JB
coj/JEtxHcFUktdgjc70AMNhtJ1v9kSVvVfOawmBV4W+gtc0WrPPudLsJUeNyJF2
5DPb57R3VikB6IhjPTeEAj1uD3M6GY4ExaNbjao85P86umYOhoVTmWUN0ZzqFg3Y
m+GlFOr4laiO/3QMkXS7pP5szhmXS3TE3+ziLhDeECbVeQx09VbX40z6j7E8RBef
/5IIUtZVv6dcvg/KjZydLJcVxaOwyN89ijdtJsH0Jxc4O6JvDSLMIHiSZNBcFQAh
/exoaontVpwVSvnqt2P6pqFZ2VzkLjVd5ERUZG9sR2+6U3dugu35/hFNrVOG0OeM
H6myDmzKBoD2F+Mu/R6YNj6D4FgM4GUUhlt1va6TW7yAuvzeeU7TZ/my+i4DQWxX
GpGgDdAw+0dinRGeFiin87IVb0bii9u99wYehamNtB5J6rbYgmzUgh8z0h6A++0a
LX+ZO3G7BOj+l6C7wv19z37/xJ7AIi3wf6fDCdT4fBlfpukmBpwNJx3ZLzwpjKtb
iRyEKGXhe+/GHcgO5YJpI34hkyjLMLP/Gf9zpXf6IPX5cPXIugpJz7mUqbFHJ2ah
Hmk6GCWCRd7BtXSf1Zt5otSlcP8crzAR0vg7T/LCvF7/tvS5cFOgKcNpCGGnznw+
V7XcdRs1NmjCGiGmbe+zO6O01P+cqb5VSIJ8KmgLD6zae8JOlAYTPiIoE5NJspqb
K9BfaC7C2YsEQ5BAlBswgELFGvoXgyAgcB7VLAyuOeetIosGB+fOToBtp3RwwBoM
5j65Tpze6S1s37UIIOaY6jF2znyRZtgWhpZaqjSpLJGEdON4X79u6Rub81BhrFTr
dricB6N7xi0V+y73svkbbVJwuPAdJv8VTH3skTkKBqEf4sEGFiDN1t8UcvVoJt5U
+FqjIhFflfiP+/WF/Fxs4iYRw3hUb8qruAMvdzr7zdxZkTZRqeWvKd5qGr4vgSC3
uU4pglPqCLLINiaThWuhJE6NGcFpfMm0rO7887LWZxmfuU8F7Y60QGZoiCCwtRTj
5HfxVcRQUAeJsnluL1FajszALntrzq+6I5x69OSfxCFNjWIkWa/PjsThV0qQR85h
2DL9+6+eVYrIEEev+s3W/8cB1q50id/P2/fE/4OWNcMaD7pGypJU71kcblvwnyVF
5dkrgBpgdZ0NdGZAnuna67oqgE1JocOUDYe50PYLGy3YaW1oo9mFuqi9DShSh2CD
4WSYpfnnm2tdQfwYr9hHYgG2UyWv7eSoKpXc8tf0Rvbw5MpKagnwgwOI2VuA4Auf
gnr7EfO9B/hLqXc4Md3R0DgBnLADMvARMQpyOvZw8REtHUgRG3y7vu9OPgGP3ZCY
kPc4ZVlXFg9fFeIdsBjNS33DpzNg6XNWHWb4niF6E+Ra2Dsrm4YqBt4Wgu+3MFDq
tmLs01wgg72LpcpXpePLG9D6Q2cAKvT4vObxLdYxm3d44zKoyUVa8brEQCQ3G4j7
zHsQ9j7yQIchCyYAKPOc8GwU3M4Gc8vafrkntDud+II76q7xsO3+rY69knp9+I9F
D7dNHS9FCAEk12fZSRaacWT099YHfUQw5Yw1/eTvodEhOB1StKtsIHJuUHGYfU/g
YlgHt0In+qT8CVoQmLUGCs3oiHK2JYfGp3cUzhei+cvyG9vUEReFuLq5W+K2pPc4
satLdqLgKUICsGeshoIeWCdZI/ClqJJTIL9FMxEffJE3egVMjveVcN6bFD8lE8n0
h8zBGj4hpjm6Un7ZEn/kxuavB725KD8H5qkZDp9GLXr/ELIC++HAMSDax44bClRN
fIGDXR5HeZMXz1yWVCJOPo2IwoKGUh5AWDAL3VFmCHLTOvgXQznilykPnA64yPJK
9VPtDnytRLLVNq/F1WMaFv+x0f0ga21gEyX+itCEDLmsixYnwNlvWtj6xe9xbM+3
pZJZfX4heAZn6wzBRXRR/P3O8ACSmOv53bE/85jDMkDhi7DTUx9L9rbFgsr1CjX7
whac2iztAA12Kra6fLvdOE9gPxA9I+x0/QARhQRE9zzc53nDujtjjQrKu9EcUrds
Fh0y3S9H1SXK+nlE3b3ivI/wLynrCKfmrJQxci9sRTAtVO6XxcZgIyKm5mEfZRR0
WloCgY97Cft7wOvTZzciK9Ih/J+2VgJQCDboPLbYxmGf9iPXOAMRjGJPpNf8NvPH
EPV2O0zA1H4WYrDq9g42a8qS8kr2/otgw2Op5p8c6VVEvSrxGPHd/QFawQYQOOcc
pDAF+gQ9pP7QHpb+ix5Q9FcUMzMktqpYH1K/uLPQzsPydzPBcG4RZUtm2FQAcqLH
L2zRvsxVF1RMa7JEJcjUOtZ7HYcRhuZP4tXf7kl8aHcOGq2axJmHfIHeS27Tfo+3
RnoIyah7PmUrj0eJYCJDX+BZqAoJ1k2z/OfK82osOhF+tkSoSXZlH5QKZ22XR2Bw
COFq/Ur69Jj8wsGJpYVwXod17dsWMPCKjXLUJccjO7lvaZUuhOkaq7vB3MMQFngX
RJ+2fH5OUYUao49995xPn9222xbHOAbVEpdYRfQqFYMAgwxlwk3dX9QsCWfW9Ld/
R58i8pF8+KNmqRVATBCggclFN7qVNUxP+ylrdYbTrpBomc0BjWcaZIZc0YubdFCT
85daXoHOcXNAsoN5yxy5NMXfaH5cPIKctBH/uNTh5qL7Q7QJUGLm/+GCq/pfhyEw
LipgZRgyPQWmoVzbRlaylqqC/gAM5P7U5j48TeURCt/auXTJ369WNKjuMIuqmZoI
ASYTXSCzb0pUo5b5EiYBWghLoVbWBz3SAiavfhsG6kE8V2zBvRaX6nnW7xnfozMH
Z0L44sLjvbsoIJahZa9V7ssEs49I+Eh27VVG8aPE42PMGG/TbBuXOLSqVdwYJL4l
nKLktM9K+KEHGcp8Lwb/Rx1kfBeZyC6kBUWJ8fhbmH1ls+ubqjs4nKplu+2aITEt
FQONmjiTKs0a5zFB6jYOYwUcqp7TBWi19Zqkqjl6JHFpmkGMD78GXPn1QDZ8JfRw
Jqeorqu6QeNRZHSWQDwdTctFxORwqo/K/mV/8BuYI6dzonJbjshb1zW0v6wgA8j0
gTJ7hMZkeWXjjkXi9spoEFLDXXGuvM0NsO9IOoKwxffTGGg5VJrqhotPKabzWRwW
s7e85Lm2o5g4Yz6/lb2pufJN34QFWngHmhdl/7dJ7aLch3a9m85FRSYHcPWcLLNZ
pWa0CbHP/sR/Aqv7zn6p2Nqz0CJ13/OESeTBW9SIc5Oth2ztpSuZ8ZMuvEtlyzOb
seVZanooOUHT4gRHmYvWjX3kHH5tHEHYsK7z5K2PZc5AOvVZ9bNY/BhuqXOjqa81
FGBbYn4t9SfCieE+w6ehrfs2pwgmrc7hhKj/B4pyBQ5O5NO2TqIyd7JD+SYPwu3o
e3eexeqGveRGbA93uRZCv4HUbeckdGVsLjHLCm/PdukVeCL79WHvYxVWutSQmNY0
Yqp7csAdlogFq5PVxSPh9WCwA0bx66oN3g3BK47FezmTMCYlg/+fiFlAiOLAARwM
eE5s8Av8ZVxcNmoahFn+9zKMYZU/kq1cEbdJ9P1DPBuPOlA+QAhvOxUl2Y6Af5Uh
jgpCOKH8C7VrNGSySG29O+QpwI9PaIRlJZwazCw5X8ynLLDCdju+v+BN79eXVcOo
H2Oobw4EfxOMRPyJTX0cjfQmtRtseOutvnjFjisjeK1pAIjTaHia0d40m5zlBLvQ
fOBV0kgjpuqcf8YFBF2jymV6cO+38wbuV/sC+Z6uS5iErrZg7OTlWV0R0rI7sGX6
jAEiGBbPTqJsvevT4HoDzn7wbeaQ3CTSblJsL0oFqEN9G6O7GLLDSZ5Wl/dEsguo
3D0lnM2E8qF2gjqvFyogZsuCK98o/XdsYzzOOCBIiCdnW3ncVPy9YOlASQTU8cYb
Jc8OsJkcANZ68ubIM3Rs5VMidTYJ7IFrC7EPsQE78uxtpB2PpkOZKOnlckFzNPcE
FLkeeoyX1MzmuQJAk5Q7ZwfaTgPJtYO6UYE7kOQnQfjkYT3WPyJS5PxbkKXFqjrl
8xCFy7A6jXD2Em0YZKlytwQIYD96i61o2OgnIbKM5A0w3B/IiUmEurPC2Zqt+EbR
iBtR9Tn/zjy2n57apsbzTfLrAaOodthRyJArN58fvbQr5XZv7pXDyG0t6ULKan4M
LHS2irnj8fUUHBgFPRqgtnrMz2Vp+nSTVIDMe39nPBse350LHoiF2gQ8u6b03odY
sIzLDhEiOEzhEqdivfhFHvY8mMMlJiI++HHSRFaXGF3BWtrYWjv8Ok0EZyQNsFxR
DqLkcqX9jGBiftviWCx3jDdLm3C5TRbK/ME7ojQ1wmeLsEX4F9qRGf/kqiR3/pAk
JuuUBAJsc797/6klEv0nfRN25j1tJa4DpssBh8/RMCnWKiR+gTOhUsPVueVccc6B
R7p3LUj7oJTr4x+3NDc9bi0U3EMA4mD8MR1r+aFjm26ZZAdkQgYQ5/gXCoojKA4b
o+yLbzJS3kbmrhfAiK0PtfbkNIezFjXYFyKGrP6yjhLuyDQDfVLtaOZ4mfuZEDSq
0gRJSP/1FMw8ISR2UwpYmGeYp00Zy0o/lHK6d2vwx6opsqYENOLtJTlOkABNG7Ea
jr4ZmrlrAcF8DFvdnPYyrT1q+mCo5PSBPmCu6MSLNjB/odWxIyg+U57od/ct2xXH
TkgiPbStMzsPTeOmXfAo81Q6EzrJcaOYOO547pL5CcbDVtlOd5Xmimf4USKmA7p5
4GIdTYHT370LtPy6UvSMuUkeBV/EyceUY8BZtVatAerwKtbXdveaxrVVl9HKtFOL
qwg+W31jfqWMPyCCwOet8EVIcszeB6fo/z53hoZDMpd1gxkVdVvo/eHLq7FF9xL1
UG/KtExufHmvlmekOaEYPMwkyqoI9AJZNAeatvtQov2f1Te0K9gIpuFM24u4Bt3p
a+YyflCOnduk/gNfLA0lFRxBrvUv0hkxM9HCTRdDXhUwT3Y+QzyDCf4sTanyVkuW
POPYRLXB+VKWc/OZdeUcAcJuEhFbrBDkS8cDTZiTD6Gy8qtu+DNl2kOMCzCkPl5R
wOPaMen/JWD3VlfDmJ50+f0LuU0cFwNV3aVoYp5WFsv0JGAc+HfFEGv0fSa/01qf
KP+7VRgnKcI/nEmoObTJk3x+caYF2SoS5V23S9bAnwUDC+hIVvq8AkOtlRlC8zzE
2qwfyxUK2qLVN9wZSWH71AGt0P4lJh5twEAWnnpitKHKpG73vHeCKvgXUWx+zUwZ
rR82YP4MKC04jABkfcuSzsFupJM/EVYmQfV8SS0OKj14791Oj+Fg5KNXMTQOFmPi
kYiFnjeHoYJf4bY4eeyLTIoX0/zaieEIatyu9NwlIquhddw3dLD10qYkSw0Qsudk
ufdD6WnEbL2C93CbmY1zIl73cco2lOTmWhLGv60SKMgijSEzes16Zcy+ixPkSBou
xFUMAtH/RMaS3yqgWAYbSdUphaWPaNTwd78kuzhwSWtqrnXHm+0U3MpgUh6GErCA
mAlJemq4phiY/p92sZNBc89baeP8Mg7MAQrPgDx6tQ1I9M+scoi5lvXCEPlo1Hyq
2GLmjdfeTB+PAQdk/DCEctLbDDvIxX/hNiJwtEMqwLJoPTvvx27Yqaj7N4ooN+eU
8u8JrDnBNPYhbnfC8g3EEfeyXDb7s78ISH4PU0H7fLP0ZY/6GJFfdHi8ORaft7gI
GX9pk3ga33+FbIDUruuuMNDQ5SCTP0qNflrAyBbFBRaU3RS31G3osnpDz/wp1CYU
dToxJludsnw6+Wi+JWbONpoJCrIRW6Om0gpYktm4ExwBIkhUHyn04UyC68m8LHKr
hKn7wIa/X3tdfFIGaX/tC3Q/DhyvlMxnqsGaohBwMdhdjgxW5LPXBp1QoI8YFZBl
pqkSRuHFnjIOCY89azanbE6NMpK9mf3whjICrWBbK5YtphsBOaVnQz3Cq+rF+buC
S4xXgooYZFpOgJhdL1uR9GS/F4V7+5Bd76pTwdwZdUBTigD7ZeKXM7o6bqeERjLz
e7j/simuZwQg743uy3rgEwuNlBxpvP5RzGtDQ4M3RwmUZgxJj7rFXtkZp4q67r7d
rxtLAITtJ/zFGXh3vw2i8ZPMt41Ma5xmxGrg1TOn6yYEHCcBegnkVudjjAA1ragO
aUmDsPeYJ6ncy/bltu1KbCOGsPE+Za70B8EDY9T9Nor5bUAy7t1O0b/sDQ1kdqhO
FBQuGVD8ktkPWtVgECmIYJnxAFn6EROwDUAGjtOf+5LeyTFn22vkenS2JC/Ml5gx
aiFAd4rwpK3qu2Ov+B2mKlIVvYIzVnfFzWknlJFzM8wNXqFXqw9Lql73HdZRGEo3
HmPh2lLgb6BE1DeTiSRxwqj/gYkdGPNMnz4nq3GcingC31LXk+9wZp59bbsFx0Ti
MlajtraY9Glw6R22GH9B3CvQdw1GKqrdfqmklbo/WdC2nc4r77C2IKKXlStsE9ZW
O5BT86wHO9c/7S4bzC0b+4Qpat0GS7C7sa1NCJtpRFJ76HhiL3547q4wq8rKdj9g
rWk5cX+PhsR/MIXqeUZgDJZdaCRHthRC6knM5qDQETGSs6XRDZGixagoypFURaaM
G3CmTaGOd6p6eb3GQcDcMpQwzOJbe1YVidSzfb5WVKmA8fvj8LkpDzCpDcfq8Wbm
q9RDgzVitlXcIRAQNI+XT8Rg6NkU8tDMI/mZBHN5wDx5B6vkSq/1sXYTBi00sZrr
HHTv2TvamoJnBVri9H3keahMxhHBu8zKnEcqz9xL+iFQtbAnurZhhCWvEdRpQ92t
goS+ogoobN1DZ1JnNR/EKzulB4xc2yTcVPDS5YPER+9KbADMSao/CjL757hc3h69
y2XovgBRlF/HaCj5KnzaFy55eg8HSbiQhhY6rOilzx2+IPfAlg9HjGR1AmUjn0zo
QJdnokR21A6FS3vxga/UQrICH6870tw69Y9zACTrByAZN4UMD/D6mgnAG9UA/jOV
PSfhlyHnD/zQ3FWAKdyCMcspXqqBmUkmefuVGghOQMT2YJ0GW0+dmf5n3Yyt71LO
7GLCFpZWo04Nagr5/bP6Yn/QQn5vtrU+IXOe+tNY+ItJ7cziVeraSXuBAZTyiCNl
BTFBoIW44ofryLWM9V1U6z5TjzNN+u+BqRzU6U8hsJYGD9PDNPi7O+zZ31uxYVNt
L5U/+1yEy5gcPt99SPVfm/Kuv4o5ZH8uS9nu5ENfZGfiMWqyulMaWcVaAq5tZ4lr
Qj9ZAEF0DWnPi7lJXpsG7TiImZjsjFMrjfcb1F/XsU+7FjpwZUaSUmSszwYulzc4
1jxV4Z/6QLb+n9qMI3BR3wCCY66H4B3vzLzMJ/VRDPDq4m9/ynSq1aZL1FJuT8Du
5lKbwl15w+/XyWlh1c9xPgFv1kCUYyhjXCe4rf/bDgny7XPzErobrFwGum+d3ku5
EZiN29AkwoFTmuob8VaergJADps3m9DcFDVfOdDijVEYWJc9JWUsdYWmcAxc1pYf
pNiwx2MxiUAlRPdIr5NVr2UisVMxTIpmIoo5sJ3c81j5I+nWkRYiM7lJYURX9Mzl
J2Pd+v8MhRbOeXSwvPkWVCtDGHjKhM//zxXd22KHtVZj+64QuRr/7A0HstlRf5Wc
JRdm7YrisISiZXBPEKk3OvVfn6elZVNFwF+T1oySf/zDpA/xAh1nglX71Bp1rE61
YzlP7EbX1DJmuTmCGn8TEC7m/ilTZ6HjBMWA9YHN17QEdQ8WhOugjObaeGgprHtK
etlTEcj0ewsc2+FoXKMQgJnj+93ODgqFjWMw/cULocX08SADqmtXB/OslDP72EUN
cqCVR7n0VWvK76jy2FjIhOlk4PUfqLP0kYpZVwcuvUI1hm+8t9ANTlhO4kiz9qpr
1Uql4auohyTTYWIxkW7rW20XjEfWlfmM6uDkSfWE+yAY9iC3UDcxsX28d0d8qaHG
PUtC9LFMzcBGxoMOitGXCsUOnQ5iDblrMbqGv7MByC50t88TIEsw3gszYn/PAGLf
PjgDL9qIkxNOrWTjzd1ERA10Eb39dB/dyqc6gutu+ZrUpuPnMa3W8XcwHKasJn8/
xqeoYzMqu/GcS5OzjVuZGAkqA51u+TllYp3gIssdpVJL+kH8Xx3dc5iWMsJzfldr
6ekClhEmvRy0wwX2uSRBoR79a3cxAQw//o1YPCi149M8YoO6tQN7QjrX3nA/ZFwM
PYFus6EmssKbYZonMZUW2wMwF5IVKypoW+twoH55f47rr6IXlur4w1P514pDhEtk
NSQUU6arCM8hNKKT4M+mwdRN4/3Dfrbcn4yKSfK0Q3jbpPEjh6ep0o9I1ZO9mP7a
Q4vEoWJsDUjqkOqt3YSaUFsR76H6slAwFOLCmoZJe48hAWJGsrSrd9xetXBVM1Y4
4DZNcciuSLSzBW6Q0aLsPpy9EEYW7yaJHkhfOSxAfx4YCeJjDty088AqfcOpBK3p
oOEO2xWlaHnlbytTM29+3DT/jLmOnRGbTKsIPxJvqb9t6p5qo6CK230DPQBu5yn6
FAiMINicWgI/hnObNjOyKWwcr+RUh6wXRXTdNHOddSmchrsRDGTGCdP7V8jcwm3S
B0heCksMYcpqIQb/vMFrOKBGbt85c+vSnXNsBF2sx9lmMbBjyL3tTxmUgaYXetcV
C7vAahlprldh7cY6qrAlJihdyOplO0gw0IS5/ppxdXz7dZ//a5sYKMTLMegdJ1G6
QSdCW4U1vjMBm1xPKu1H5Koy7dHiqO6Sgiih9sytwOZCtQTezDlxzy0xOYuP+Pzu
SCJRVcgLIJKYBfGsuqGGTmH2gOXlorQ4EYmOwMZJLAJws3yCI7iigfPluVkFHY3B
jeDNxSTy5y40jv9lMdIs9U6lcP8TaIHZJt5AolGCIHdJ8qG2zAm5zHYN4GTNvqeR
cXVq7idlaEtvLnpbmzi3yWCEgHP35mc1VX57ZEr3qYLA0jTfSAVM9HeeVq61TTD3
b0CEzAAqqkQPY1LJisMpnKA25vf0xM+kEsEm1Wqml7FtjL26l+5K9AcCip3XVpT7
NmYUIi1bZTwMcoisRhFFlj5bHxAx4Dj4zMzg1MqWLVOqXBQT5eER5hCso11EOQpH
Uqyu3S5hRG4of8xAJnSnbWNbbCSRU8Q08If30mDQH29/hjt0aoXiDUC2oVxVYQAq
SEKciuPmpPCPfCcUWsUMP3j6gkTWd7ua3o/3HKB+hvbM3CT6pm2dtBNF6i+k3VPE
XK/coKdnRMGBvQLX0XncTgkfaF2OhzzLnJHCXsTSt83NbzaVYcZD+7PVkDRZ1Gc0
uUFZF+jmX1xZ5aqpdo4Z5RMJZYz4aqGTcX0bKUKZpxtNfqSTiI93uPqtRFl9O/wR
dYtNUaR7TFKQ5K5rs9Y7WTkea5cxDP2SrzFWoaONh5sWFRxhiJsz/iqYWZh/cxho
VPDo5oRntHagqaHVEFGhy11R0wdURhf3Xzb+s+/CLcouhLjympbIEauZGH+6qeox
EjzVs8/ittM0XknEvGqMMABsrjpJgNjT68Zv9n3k0JODIa+VZTLyosfVSzOKxjmD
SXLUCgTTrn/i6pa94LF98KGfaQcHY6wOONugYep0GPbeEDrWAHaQix7ksN9oBCY6
zryKJCfcShL/qywuiVupsswHnadaV0UfeeiMYMkimMd9BvsmlJX158Tng9tYxUty
Z2M0BrC9+DMkq23+X0VrAA5FoJ/xgbi/tPV4n6Z+Kcz09rzov5CjelT7qTG3lvPs
emp3kCpSJhr/ImEi8UmoRqqHul4zX1/pgp55/tJpsjtxmiImzL1YUZwCh+WxbCNc
Ivf7/NjgEQMmD8DH0+zoV8uCqE6+x0wPx1r43Zf2zKZ08a+OmRtefRnXNbXOHE9Q
wEFIsQoVVCP63pZ+mIeH/d6J1+L0VPUIOKvCv9njs8kyUvLIp1O+hB0J26AN3qJZ
7a45NPmoiNJDCnHljptAIaAYD+wEOZ9FJjrlWOn7onuUPcj9O6KrV0XZ+b13AIpV
GICW35LGAI3oKY0YogvmqDkwz5m63vJcyYa0km+nP+aYJ5cdK7Ny+FB8FDwBcao/
LU9XEui6/jc8H6iG/RF2rwYalzvFH0sYt/iKTx3I6d+cF8A9ejDXhQzoKrlaMAK2
tb11ILPi6hXI0ek3dBPXHIp+h40c/C58tbIBtCLXpNd+8mISw2X8n7KXFCxM7XdT
fDVnw2HnlJIgpFmux2u11JwD1yikHHnZtUyf4lJtPDuBG8gjbacGbS8QuKxnZ0Uo
k6J7k8+eP/uR6FfhIAsjdx4ThgQIEbQfv1Cp1uK/JxbkmSjA6Si7G7mqJxlpmcDl
wqnkX2m9aVxGxKRH5nvuxEJEqXs097vO1OX/XsGZOKvtF1uYqABkCzXEEm8oCPrZ
49ucXVB8Nhi/DElzzeV3VKUd7dGAAJGjYWgQ0yLkslIYRlL/Y7Go8nLDs2n77HBt
mT9OBUpiqR7Q71cCpncHIjDDnc2S5b1O3COjBTkIyuPoljGJ1sGTQqzVCcfeD8F2
EPRpnBTsqitIw5N+ChD3lHx14+d5pVS5X4kGEVyCDNVadfdEOvr96KxeQKTXMSX4
O8ocC5q3SC/TmhlFLep5caN6+6yxk3tlQ2l111kqDAS/fL+fvtcHDNLxo23Htg5p
Uqdi/5/h0HZ5E4UlEN0bq1KiUbrD4wsa71Oq7NSRBkz5iPtmEckn45iNpbqGXwTO
SNO8jLdCAP9le2cXAP1uBSc7Z8sMbe/okye5BsBx9gs53KkbRY7x6ROpGN/3LJ5X
B82aGZIT5fgELYnIqXRndWTtxQAoJU+ver49BvLtYcl0vFXnsZrLN2uZcpg9sHUi
EMV8VGTYh8JIPxahc7YT7a+wgirphSgUkVHASmEUBx177tOXzuRvjiUTNzHtSEjl
G+Ii5HkLGMJSOOZYeUfyyYB52cVOCZODt4/6SYwSEf41kVo3VDqDzN775NZ9sOgW
JT4+klLXMaWY1jXswTrKQ7/aHKoQhqIdTiYPdc7SQQ38AqP2tWylLI4CGx1GwyQp
392GB+y4ON0Zsrt2fumqFXbGXOoGiM0SeNvYQFcfHIYa0Flk7wrRYm9cyWK3wJU8
JoTXcq9LvA2UzkbvoQnRkRVt04G8SfBoA2+Lqf4zZ9jzcu7QlyuSAzYgXxFUOCSN
WXC+5c4oweGBv2OvNcpeh4d6fS+ObQIxEHrSksK3QnoVy9U488j/OHR43VeTNuq4
4smtJvdKqX9nA2hzi8Qk2c1fZ3n+ODT5FgWfyV1FjBF0qURqjfsrqf4Zb073GLNn
XYLbe95PRi4uTWlLLeJD4FhbtTPcSmweghVZnlAvuNoh/EhTH7+rsbjB1XOpAUd3
/uN4nbg+LjX1nSNXRHJwop/TAxEKMoNJGOH8z23FSo14PjiCeDBIFoHMQQEPIDKU
3Nr0C5Qhn3fa7oJkjnWmn/gKanxpgLn7+6C/g+qHPuCCdaI2zsHkNrc9sd9z8g2j
ZPmQYfXlHYevY4bm3RaTEPU6EJda1b+ANXuNuqZwnHoeG+hN5cdG49yz+thDZ5cj
56YOiDBnD8aTjOzfulR+Vozr/6Q2na/uujFu9iaNArEPdWLP5ySJw60zr+77f2es
2aLYwF4lHgd/LrJGgGXBb3bW8C+zvbnw21TE7nPZ1STYP4SQdRJX4/D0ijYoILdq
gSmgvxijLdOaomFEYmZ3sQvSUYATwF7XdtpDitNpMIa0P3VGiaoG91P6QdKJsZFA
xxlWNjOBDHBSw8AIdEfLnLkXEndQvdV0ts+y2YsMje56jDMTLBnTjMAmB/Fz9fR/
sEHs6XVWONxAp8bVzdMF0tD4WkJHd1o+WiIZZXP8TN0fodY6lnz+GF8G47lTMkKF
l6RjHKHGIVPNtocojWL8bcQzOAwAb8zkTs38y1EhuizGFzo2iy/EjrINbJVmdpzc
Ghkaa87/oUmwKMSRkYltnt24cbkEJbJMdPQwgN0wAL8SBHZViUgg7Znjr6azYPXi
cwrxuRhWfcLOr1D/R9iZKzuSMh1WggEGipj0FTSjQ6W1KIGCDHyk8zORGKVeBEsa
QCyGSzswyYlEXZq4u/e/caqh+EgJwuDCnGIhI02xRwWnuB8DBZWBaTRkNIiHLWrj
4/ubr2NQvZY3vAtvT7jf2npHnGXK3Z5WH1CH1vOCcmlG2RvCKwKxhUvgb/0e/FCt
s7gJCYNtjaVQz89h2ev/NTd2U0bDulfLosDRkw9v/0YMOknZoTACWTvInbFHXqni
BHj3vrF9J6jrC/KoA8NXEbEEYcZwpDmp2JSZ9nC99XgnEM/HWGVl8dnCsATL5Tgl
NnorAc3CFXtasR0jkOtWrJ7RkIFJ22vULjMFu90LR2Rcrw7O6OvyeV5Z2XduPpd3
ft1leVbOXQrWg1K6Jp9KouzNqzxOPmTEpCOSoHvFEEb7fDIleQCUHG22F9lvIRUF
oqWOQQ+v0F+f2c74aDoZE4XvKwzsrltZvrzYb4g/5/nSwJOmszxyb+RTFCeRqPSQ
059qUjxzxziwjA0YgETMeXTBAKpQlqV4LFrN0vnPDgSj7YQMYJkYWcBRbipg3jJI
6xfYRvoEWyXLErScOuaeyvj28pysm7zODnzOTxV7Mz+Bq8E0ZaPm8rEylZZjcZBS
Taw/229ENp+daPX8zyD5zgK3J85Cm9vpOxGo8xNSI8GyBkgy0BPDfnIeSyNuAH0m
IOX3MVkPgVEZHROJE7aB76N3JpsxVGSftU416pgoWuMUrRkm9/SCBtE74pnAkwh8
SgO6xpiI4BGx65uPtV5RPDiJ/2S6Nf6qcb5Jlsoa9SRE9+yB5lljiDeSC8QUThiH
HjutYu30aw3MYa0fMgf3G4SnjW9pxbMb2BZmGilZfbYWi/tKi7fxk9csLBwe9fqd
fEpNTD7rm7omH2sG3VILlkl+DzddV2SKuhzDSN2KrPfpnT6y0G0S2YQTGXfhXJNb
+rzjQ1Ywr0J+1yDW7nE5h5aXKBV00JJvewf+gZS91yuf8kO6E1Zge+iK+Ll5UbdX
uNFV0UOqDgSA7ac9eC34GQ4IZybmYHYiNBPrjXbiNBsFwgane6SJk9UcdipraPy7
2Gu+0MNQupCNMfkcMVffRXHJ3/tOoEOZmoQsbn2W0olQIVIPBmNLhQs5gXHhPZhV
0qHpDKqjCIXIElwxiwz1oiPuB8mq1rfL2gLgg8pDI+WXFahV83Uv4+1yV2Oe4W7V
pe/QwxTQ1oIz4Qmc71ecNx0qtJDX7ew+6Vf1RjUqlDcrkZsJKG0nMr1k6c34NHrb
U+Nz7SFC+N1pvyscfeZ8Lv/iyZapg9borxLNqEUKYryDyPN/4CzH9xVXNjlS0KYm
jsFBAyEmeo9YM9SUbF4f+7n6DLBAapSoXHkRdDlQgisox9pZVGbqOpOTK62SC5Sg
grkSfgybR2asbrd6TGvbPYkV4sPeHHlV5FsezIL0CyJ8PvXt9h7MSJewA7g2g2jH
dH27clNzgv3WxOqa3KoG6/HroRhF+ddz4Iy7TCk3bjWkGX3YFPE22OSW898P/Nnm
F4LUIgDeElgqTmt81kMxLRWoK5cTaJPe8P7sJay9B0S3I6Fo3f26zINmYsnc6x0k
ExCGDJijqv5wVOGRFiL/AHHzxxXYPlzqCh6H38wkT6tRuHLlOWA7I5es3imPywHd
i6FAhgMgsIbcmKYTvPJLaBqOXSgxrxTIh3wplLXQDSZ423wLNJ8nYcYLwCjgLg0v
DsPT/2PUJFVBT35d66nOf+YUWF7yXQrOolpWyAjnBYWIPcvoQA5E6J8H8fuBngsP
3nexCjLUGpmLg550kV/sSXVAEbcjXl9ovfByXCO+H1a+yVARpq1wlH/EkEf8muaq
ZqfG6nOCMkF2hB18htDZ4U5ThxMnqVr04qbLMjB8Z1abc1EhiWZG4XPdsDyUggVS
fd4zvInmz9bBCN7pJdZGudzX06YxB2U1FzTyDboPgo5sTk3rc+WYlzmZxDhW0/8T
CcO4LTeH/JPzz60pK00/p2PVdwq1P4LT8GIwY8E/wzvQIJzTLBbDIJIqlQCTkS5s
8eo3j78gbv0anr9GSEWc977QgLONqtiHA05pKLxyntjCVLCFmp1dKSrY2+I3Jkqg
xsLdL8knnz8941IHnTMOX+3TMsq32iYK0gUGNNTgXYHOmT2W0iHcvQ+sGcTchiwv
eoZ2+mAfpD5m8ZoRHz7+/Qtv7V/ApjianpAXF3KSk84ndokMibEvVxJsKZQgUhGp
YjQu1IBleMMJ9nHIkh4ZfbkSkGBbirlytSvpPaOLoM6daQXZdCF+zVn3Oi9a5nPI
PolatEjwOZ4zteC0r0TnA/GFQWNrDEj9mSdAV4KNkQVnZgP5TWm5jmJPVvCFTFAy
wvFyz/kMEW7LGzYSr4hsW2om4PHanqvKpPYPXKWeNZMLOOkXlVwrGp9+l3vmD+J6
vGpyVZaQLZuPT7X3DajPZNzrn4+ZvzNMqNxbdIWfk6ZMo+6TDlMcHwJRfNGduT+G
eC14e1wS2lEvTejtwDALElxZk8f4ujcO5bC6EGTF35sZG3bpK6Q9wSjl3hJxK1Bu
D8R1stkATmpWrrHRwCm4uvc0FXaNJhikd/YbzuCgoU+oEc+JooZh34XDOS6ey+zP
UZsdGUySLovMV18s6PxFpm4rPtZoOx/+/h/aI3quxSPuY2t5YuOlGE0VYGbG1gAv
E8grOurQQZMZ1XPPFayBk/U3834Dtw4bTdJ5QLYC6CkvSQWm9WyUt8f8406MwFxD
L2xnJL3o2QI5ed5SIlw1x0VoKvsJLesfqHNgRZOQmIuUiwaLWD1TpG/K0fGOi34v
37Pm3nzsioJRzh2rdkT/5petZspgDqCAyRs516VuniJ5JLG9QMfQaX6/TtbED78P
MZ2uhfnnJyp7DDf818/QbtAYHzedkS4JQSgknPoREWFK5/vx6pKXHIamPmRmLK3H
xDg8P+nzi9deMD2zeUmBqc6qLtUyZLjPaF+dSQjPhyY68cwZ5j8Ym1srNNyxjTnV
PlxaBOmjGJUNBjYvePEGLqK1AmUEz7uOb9mo00lok0yIWB4HSIt2d+ozH5JRr9Dj
KGOtbw87KrMwVVh04qhiyvvV0MkHd1J0pmjegC9VkObLlksBdekBTXkMUZK8Yrki
XT0Huh7rM4cF0iZREfHFWo+K5dRYsp5Swc+OSmHRujdAcogf8PJizpkGHVcaApgZ
3dleTBjCuQ/R0ZiktKJ4x8v9icPeueZvRRc61uU+uwd0T3yGyDBUjTw1AEs6LA3Y
r2V4goWLl4TZolq5/fmi4CoSXqlDMZUCIVXS1uj004LNPp45i+zY1ouF648L5lbW
nDbAG6LJRKNImqe7DyoJIq8k7bj3x9CioLFvIz99LvWNQdZUqKgr9xsf6JUrEM11
K+sTnIFl4uZaBAUCSp6CdNiwj7G8P25VFWFMAk6dktyg33mcyBhsdQGnlf+SBYnK
Jtm0nImkW+NmkK1RWK61W28y94Ua2sc45GBI7osZAoZAeZfJUMWqQE0NpkE5/JrZ
o+BbeQXv+p+BB+fy8MPGZWN3rt11pDLZttnMXOKYr2vVG/X4wdSjlo24S46X+bKN
HJK0PFxpKdR1/4/bMJX4+tTNIbsyRol3WBeRCL4fWnXezeCorzDfivPKWKv98rf3
sA9watVUKLLqz38FDWnpdXwbIz3Uq/oHAryrxzNbrIwFLryrLlGg6d+YeBBXgqqh
tPusT78FfBPODtDc9yBs5f5HygqYNGYK0cOhl/fRYbWwfaRFZ2BJu/vCgatEBLOD
oqz0TaX/+fTcfGul6wXzzCfvLX4p27KLD/XZG5FHPdH2/0DD6lOFZwjQ5kqp9y1r
9l7rVbRa3V/hRNN3ua4kBmZ/Lt9bjD4FX8dUhVpvgmaPPTSAqsuUDRrYgyY21/cH
pvrFEPOb0KDltBR+VvwTF4rzG3y/6DvTDL+2xfW60zak6XT4YdaSlHZO8k6uXUc0
mU+JtVucM++3GmnDOFnR6CH0MwdJxDNmzyCA4HjZTdBS7GK9YzklxFQCCTCguPZo
yNPrRSZrTVjUv4IotXPc6zmQeHJpoB2Hcys3PC6Oiv/u8inTjEY/SjtX8JJf7mnS
5Etye+mHXqxS2f31DUQ8JuNj/DQvzbpOYMlCYK0DvUrnV7+hkWyiwfEM9+YT5fCV
7hg7a8yfOKt78eUCMo2YS2zshzLsAu64oOA2OKIm3NzkFNCINVrv8RlGauXrZ+dy
72Sc9POlSIT/WlBk5ImYfGXcQuZxL/2DdwbW7vkJ449VoZG710ZE5+1BBghi8Y2h
zIH1mjl9zRGvK3wfBRxn57V++HbbkuxI6CNG2FCvaqlMYQuezfmzV7juKA05i0Oy
iDWVKMM4vvIgA90P9xv6nn7C4Zz+Ewaz79K3JoV3G9zonBQ+e3QuVVnl0DYSBLet
d/2j/QoUtNV3DRh3o21ZgypK0u6mvF/3s5HGp6BdI+4zpDpEnB4bzs/cBfksfj8/
1DoityK1eWVtNIW9cYB3ynidu1Yx/vfiyerRMJV06nJlD5xbD4g4HFzHd8otWB4b
Y8IuvvrmdgCHY41dHnjUylMk7UeOq9GUkPecsAL5JdoOBRGmBdLHdVykGJi8lqt2
2sqrUKMlQdOkRsdHjaYdmL6oupwom1DLZOIPPyLllyykgSiz9fze1WOGEh+D5NXG
vot9AlD5n7RTQbJH/Q/mKjzBPWRKvlQDiuDKLxXR6JGkrRhNBfL3ijsq47p6mgM1
/SmTuYCZMBG12HZX0jE0nZlb2R4M//KmGhr+bk1D6dlF39qnuLQwP/IUt0PBr6Gi
FhxeptvFj4wdzEe353pcE9ppZn6MwdPykHkutTslR1vd/DN72D8E3y7vUtXRphyf
Ij4wxPlQoYSOPERADBu7MPVx+SG8KpZ2tGj7ZgsW9X5YRfk1Gisr+PjJSOGKY1fx
FNg0PYTz2wS8XArQPVtUQRNkQObs2TUHazrGcDI3UZL0VVut4GpJZElMxZxpIYgo
3uABLR6/MbaXVTRgxXBRSIJ8A33l/gVsDlK5HO8F0Iv4+qTOef9UWvrhTB0kVbiS
UVrQ0Rr46dn4O0VNMPfRNdbgCjm/gvm/M0JNFDgdXZhaSAHgxwU/en6fnlQq5gwZ
gRguZalcau+3aLiXnrc0foSFdGVVo222JJ22KU+fSSwhv9vHMWYS7x7rqfAufClC
tIwEIw8HnkAPUu+iJRuLY7ppZEVejAIN1poK6PdHMUsRoczb4rZb1cLKFQdKWRIT
c9Ga78HVGo6C+iNwSm5T5Ey5u9rmgz1l1AqlFBrdHsx7QOwfwWdRf142UJdd750/
ZepS8Vji5/cScLxhw+LyudRDWME8wudGuWqmA2IBwXcSC/6CfhwI016+JxcW7yCm
HI7cC75QUuuX2wl/gbsSGpBa5VnhJ7bPN2dzZMoepZkpbf5WPlIljTIqlnvpmk2P
F6l/RRTgN/gHuUZbxLLz/b747y16nnuBiA+JpOi5CAPHt/vSY1riPHSuipzZEC9d
H7r0XM3jzp5L4PBjC3HIzOebGuW2mN4knu+dmTsTlk4zbeiFqLX9IwoVaUEWTFtH
m63m9HG/4VCWJOa2woCiXt1IS3okJHeTiPtdWyZ0SjF6r8PFvlLkOWXgLllo4D2y
ZCxa4MV9Kawgvw72FG+d6Jb6oGJAYyPBZJojPeHo8v9EnQTk5Z7x7LITw9PKPUz0
P6hoDAF3w3Q5K0Bg0apVlctoErgsfoa//ClAusSOm0ZYBVFHKQhX/59LAdScqTk0
rbXXNLUIW22Y0GafHnGmqSvplciU1918HM1tDjfBA8kcE8nHCNLdRdxKaTCI1y5G
NoNPVeEX+ST5Vnk1uIW2fck/3Th95qIJhGBqRp+6XW001BHAEZaJOe0VyJ97DXRl
6cmgYJOjKCskt+1Bm5t6yKPLGmfqPHMfzoLHXb0oxBLxtTDG2dW9wqpy7fU/svlq
0x/UcpItnb6WOL1MynO8/HQPFXv9sv7nBgxnvZe4kdUON+GTarmN4g4mVM3RTxbk
WMlQVLOQiNiOPcQHwE05YSiR/0pf2LhEoZfYYc0YYJVI5JI/j0uVQyeiOedNUXj2
4Q/e3nmIWCOdiS+PS9IbuC1kYl5sH33IRalszAtisXCimS++PFUwTTtmPzkaluBK
FfRaGG78589wUjEeqUw11wO5gqtsQbaATMMTd5qdysbv88zEB5YRIez+7IU793mR
Wx6i+N1/vdSmy652c20PlQywFd8QaX0kS+uFiQXl38BUc7xhrTQMYIyfjW+J9w0J
Kf+Rh8XAaVEmkpA2uBjsbVngjL2ysAICgSUlGhMxzSrz/L7I9VgSv4dpaOfyUOzz
3sUcHUX88MWkGkfEQXgz/4GBwYFN9lcN6fz4VbPCHsQkHBVZPtmr1TdKHJ0zd04g
BcmV3frHwspUXHeWWcBaTW05qj8o5JQQ2z/Hj2SE6JxPiV5jJTjJwSMp3iZWKRX9
5JYxofrtaVYr/62HAs3PXh8WgGAlZEocMfg2jiL83QTZzTqPYNGIdl5iUfEBWh6y
bVW6vDQXU9OTAy/DhWrB+SGLdrVOqyvzF4AJNzwEuGND09+RmghBQF8elhxcbPbD
TLOnPgBog35Y1ESPTf0ZEtEWE8irU8B8QFTYCL7cGamwd3Vk+9/miyABqSfYrxVO
gfmamx6WUAVafBXvDrgsbBtobp1pGbXzhwIGDcPWHXX+qPtItXYkVVLNTcWcFXZQ
A1tPN6BKX7JCDd3Sw+rzAeyFkZ+V5+8oSoP5SZx4WPlWtOzTUMzcsb5xmm/oT+E/
O4B37er6Ro5Sm30powid25T8dhJbhsGdEAC+CVyOcIyXo0D1fsMvNrHoZQGDlAlx
p74DJ4+BeqrRTYGKY4WeOUbVjB5puSC6acjzZZ5KIu7UGJl/aJIDINkP8+/APJxs
P3eUT3PnyD6tClL2oKM7bLnSe3+MhnzReoGgCM8yCffKLb5FaR+7lu/MuYQ2/iE0
Lgk6iCYSvPOuUDNi5I/TTK9unWFT7tDTEvpMTxfjK3G+M6FCJQJRkPk65yLUQWwm
GSM35wkr7OiT9RfpdMjErYJM9xE7pTDsT3/YA4K86zKIdcTbb1/ztSFvvA+CCLVR
Xs2DU/PenhT3qB9HKSSS92JYRNLYHA6kVzkigxC3kQgsGybvCwIpWR5RnsSIWBt4
dijiQgVdbdm1LfmVHSXcdQx5HvMBrr1gLkOqJjLerZ4jAslw4MZkjai423ePaL31
5v/kG2fE++UAIZRPrZS27V6ACY9H1rEDTYPnSW2iiPfnXD5XOXd9DXzhHNlX9+nr
wCYgfF2eup45KD39QbwuWDSDFZ/7IifJJE5i580dqMqs2ctZkcgNV8L7woTF6dkG
+4Rmu3tA+G8gIgXI9cHgAolD/z5h7nP2QI11PmUzO4v6LZVbqeRbh3uIJWwe+4eE
CdY7d8Ou2m4CZSSwSpCaXd3gGtlSTfzXc5PVLme0i4eOsozktp7apv4WOCF5a+E0
SHYPPi9n4tLAivnMIV43cjwjEAC/e5hlAboop6ULaocxsKoVuQES2Ap6HtaZXgYK
4hVfxXW1ww+a5DZvYHBGnGyjdjLJM3scfWxs+WUt5zUabkyHXUrjcrxQaeRv21We
htuU53wZn/cIAbCxtZMfalEZHIW8pFsIHxaHYAYuDUqCPchKhnnmjW0fopCSwhUL
NIHI407f2OKobt1pY53IHlRe52J9v0xbttYoo+4PY/oF9pPEOCU0/GVx0oFArtw+
X7lAOTDri9Ysx6OSJ2xuxhu7MKNHrVfSN3S2/4ylpF2InRizTSf3f+KFcMg9iy6z
B7yE4rxeX1H7+5XDoFbqQF3TQc3HPUtd0Kd9rVPHKMnLRiYG+rr//YNWRCBPbnea
vbIkdGnkHUNIjX6GUBeRqO+4mwWCztBHvYjbwHMEYqCr40wDY/Gyy0koSb1GxHWa
0DIU66cv3BHLFt8z8+30vnCoIQ3cHGs7ISQxsgH7/Kaw8KMFq2VtRE/hFwGhtvAy
vrQzNu9ERbIeZJpU90zBvhYA53jaI4szWNxiy1bJhjQPS7EN0G357e3B5cI27hQ/
MoF8fHTFbbweeKBbYoQytSswzEHQW6xgVTAoqxP8c9yXGCEU7J9X46uud2j+9QgJ
c+Za3tL4LRmg/cQv4FBXu78U8BikQdaL4//bqz7K2JERzewcO822hwHJfEMA0Xnz
ppa6sBqmXVkgyxSqAKEg0lBz7kXiwTZoA+SyZJjvy5sGsLax4AwpsHWdTUzWqZQ+
84sz+692ENHh1kS9T21rICWJ4CE52V7abISKVNIOYbhAXIMJ1rrl5u4JQJ/OOlgv
1lOzVd12lIfzRctfuplUUNYw51LBxPB4nSXUSpdVUJQQvpKRormzr/UjU2IqBuIT
j7fpv3qMUFcOXaSuDyUDDvPBBRgfn+ZD/Tx/9BNy61Dy/i4G2gpjFs+XQ6cw7bEV
Yr/IqyxVvDxyJjft2nVnk8fNwiHp4xAHJwznbmRWdCO+U3ByIEtVEP0VzHDzi3bM
dSbZRis/o486jvKCs6SxE6MOVqy5TWm4n7VvkhojVF7FItYh51S/auLVmgPvtFzI
23nIcXjvJEgxvX98XQc18HpkOsz54bGWQTBjVK0em0WLSoNhoVWRL1OD+shEpxTi
6tCeeZsv5Eae6MN/tOm5DynCVfyNfZw9J9limppiaglAdrbvjc5OgsghI/j15JzQ
IGLBpEpkV/BFuw1scl78XqY8U8avbEyUaT/h36/XzD+zQhruUjJpdOoyc+qHYgcN
ET+MZX2c0MdtF/UpOLw71r4C7dPbn+aRqJ6y4Gzoe2ZAnPCqUCX8f2Nx7bVfIodv
kmAZ3PTOgbb70VTKr73Lq0fS5ifGLx1dRFcBZPdCRASDzPdyNekthPvkPGsLwgOy
F35Ks2uMUScwxtZsofRfrcmL/IhNO8hQFysXQnOo5obtDGks7DH/gRiRrySQatVZ
SBmpSD8ogsGE3VtY24exHqiUDo2/SnyZM+APWQoP1L8ZyXay91t6jIQFcWylYXZd
+69hEhNYjpNGFoJCG09E0V+0slSb4moLt5shzyzQanrTYS+fCFaf5dw8PUs//fuh
BGgfKGcnamYXCeBK3WNd+CTFiLj0yCMjJNumoRVJi0xDURVlDausTzTqLjfXhAGK
q8E04Vq9A4+03D6hKC/PVlcF7rBmD25am+PnLIfywGV9uJ063XSIL9/s3u0sXhYo
PwAa2w39HtmBmOw2BGGBc3d9zO5qePdjEZ5SsQ7jATbGnriHcdEANLLN5cK2IVPx
LT8asgrGzmbuvEcWbc0tnKugY4dFVtGpR96NIxYE+kAY2Xhg5Mk4fExczLcjXcEw
JTqk1h9GA8eXwRX0a6gDYtOo/aaFgEgnKkAj8+pK/KgqBhC8OibTCB7optFvHtug
p15QeLOFYMUXjXEiMj6hpNReZB6PKrZ9UOU8eWklT1hItk4YZZYYMydZamDNdgpo
IUXx63jj5EH+3vNU5yfJ6zirjfO0g2Vvy44Ff6ofksrsT3bul0AnkdYlqvmeoyZF
Uihk9YHc38m1/wegQQ3Bqz8wmCHAfHTN1s5zydTEluxX/dFVLHgrlc3ZsIZjqFIf
31vwvMCaJx5jiFoDsvRkE5YWKmcH86rbcOrnNqW+hdLY5OTh8VhJE7D5ea5gMjL9
YCUJgUUWQ6mluI+adY4UaaVtcGae+2P029TqjrnH7kQNL3E0clFzBJTEJAvUzzBA
U2rda6szTQK4uOAYYAf2hkH1JAXY4+N/c27XIsIBWO9zhOIcfFj5ceorp5L57Ir2
H0NSIAP6E2nU3fKsG1q19pbBY7Bi/vrGZ+ctecpWf6/wvnn/EPyjZtp+Sq3/Nsmx
SiaFTb6EAJ0nnWmQyoLqfTiZmxGRbkTIB5WPXFFf+MpLUucOwxnp3flLwypY+BjM
A3jl6Hh6QFQlLW8sUAJhbVwhc7QbvVkmbkOmkypK274pzls/0uT4p6v6PCz2C+x0
H3sEPBVBaGWBKhxmba0edx5qc2h8qKSIh+jDGMKYa5dT1TbB2QmbetE2iOTaZlur
hWJiK7a54pXeIoJlVk6EYf/O6aRepg4QVzW8Vl/Kro8k9TSBDmvJAFvd6poRnMQ7
bfT/zx7dtRImNqjclDI8FNhh+juCTBO7IFQDfpIKbgsMcfMo3Xprk4eXr0z7OeNe
VmNuPKD5NyYzcfLeJlVs1eSuOGFaBkBvcTXzevaygcM/YPFc3s7rYI5vl0Xme6x9
pWIEwD52EF3E0nsxKg/qbxCJCIA0hmCKT7BMRJSnAMYgVrhxwH5qLRqbgaRITAou
vIve2YbdTNsgxBDphVCmpxK3u0sSifUdR00UqynYz5hAsD0mO6Ql+UHYwF+eqDbD
hLJPJJbF/PLa8QoIrXaiXy8v9tFa6UoTHyBwxC698/IdoCT92zK7uq2YgphsYktY
12FzeQCqkvZqhip6UUm0DsdNYm7I5AbQXdBZAnV8FnFR0LrrLoYKeV2Xk09scvTc
aH3+ONyaVedyINnsfjTylDBWAJCIuqpWJUr/P+UtNZLNGh9zw8OXd6B7HnUs2L/4
e7I0vuRn/J/Nn1tp1Ppgumgl1ToUjdY90bsKFHC/tNcDbLCYBreeNcqn7b0NPHVf
x9Dktn/AYVTjQEveJtog1H4v4xHmJpxgJTJHUQ/RtztP4+W+HoGJB0mbnP5Nun7B
OZJnMFozVQIro4eWjjE6CkvcfOFLELS0fH66w28wKhLUzKUIh8rphlhdwdWXIzen
RSRxguF474KPfZvXTu/kn6l5RilZ0P4lARwYgNZWd6QXGa8yZzvBA7JUdxlW/ELa
ZBJqXgmcxARqXV8QOjSLlyP6kkfQvgqs0mTlRF8vvayCmOflhdNokI71EsKEyAuU
TfhVt/orFXCUJ+7BHXQ/pEZO7tzn6rKeL5M65UZZw6UQdl+HF0qQBtAEZM8bz3G1
/CdNsFrxtF9SUuzHpMlaj+fWL1FhSzcesI6D2pBo5im9dTOykK5l3mpRfRIOq0zH
TToB6fOdV/QX6Y4ETcjxouvDVRUbbxDUescxJdwnpiYhiYqRY1zp+XKzhJAfrG7T
h+yyuWB1gZNzqvtfmzHTmGUSXUYl6HT9T+OZ47pzZbmIeYa8on1VKMRqH50SSJUX
GDRZdM3iwwmsj0+mY13QxRyFpEhubP/pr1Ow1Kz/wiAVjt35mbRs6H3bpNnTdnO9
kBBCsmrL/bRjNmaBs2NmcY/Xc7sdcLc/yZgGH1tncCi5EawlT3GGf/BVF0P+/IVR
JurDrk3T5K4mTp9PLq/LLeZSfYMHIdXBY8quSoclNZsh3BEr18u7iWI8NnmGL4Gd
+kJ/1S2SxxhH7c5MDoZGkzN2GVTA1RUklRiE079ZBmvK3J8gNwT9q0/N8ImvhhOl
gE+NC230plGSvt1eqWj+maaJhYKCzU5MDe4+tZ5Lfm8QwuOioDzo+qt5pdzkUg+s
iFY2u1vOobBjXLxNaHlrd8onNS7bHW42QMtHHGDY5x91o4sbjzivf3lOMa4nrG3E
QtaUeBFFykO8d5wIHpPkXBnz6j42KSHsKweso7YZZkjJ52Pflmf/v25Ips6aJz14
YOIsp/OzscaK+A2pwJdxIXtNez0zou7u4HB559AV4nh3ffYPW6Q5tstDmX56E+Yj
6O84cWuz6hAwQeIvCCW291+ghDCbP+VUgIJT6y3UmNTl7rGYFtDkvRJZHlHR8F1O
iN6Ndclj/4+JHW/fjH2rm6QTg+ktJM21TeFWqRGP3QwBxzgkVIk+208BoMwS+Xeq
VJq3R+2EJ9zemxoFmcxU5kMeMBPwO0j9yeMvGhJ4JYJo/aMvSYkts2fhwDnKy4Pu
IZerLTmvwiMznNdbK5HT9h1MV3SEp8mv/G3mCmQBnsAw3m9io19ZohJQaDUhrlmC
8R4d2MpS1MFkMOeFgti4YKuq3ql/hBVSD7oF23wSu8TWtXMHAEoKYc+5uujOSOn3
0Zk2rspKWtdE/2MHOblkqIggakPCoxwGSz8DBlBLIR/ksu8IOWG45/gSiAxyIjF+
EgqcGb6O6JVEaIw7pKdqP20EbCR7mm36+lIR73rAuVM/k1nDFQu6tTw0yU6l4RdA
/AemXWQon8aBgKbKV3VLUNhZxFqUjRgkALizv+R2EJh5rRRZroBWuxIgq1xd/hmr
gXjdieF1leQpFdDjct5Qx7uWYOjiDCkWVQIulVznFFPZi5TnUoa5Sl2IT3qPPIL6
sLeyhz1958NnveW8iFPjtrOl61/yoWzJjKT9Sy1sHxRrMv7n7lZP68WHu/I5CgvK
fWcCTLtMiNxsW2MGqhbzrIOrKrgKk76w8dafd0aQZc7EYnPKVuJ4lJpSu3lIeSSX
d19nLRR32eB7Fo4nwsj20X/OQ4nZHPE7RvKZ4W47MzAbzOF5B/L/FcpIzpHLTb5r
FbiXeRau0x4ez2XAleLURDWWzwAVQFSUpGPM+yTPUVZEaEKcGBi0J5R9OY4bAfM4
ZH9/TyRDdtqEgwCPwXH8Jq1xmYUfwfE/GJDqdeye2O1Fr0cRtnu1C1LKLHyJatfM
cyLhIxRstsCKZR2rcWMZLBAdBbfnK1LGjHnqJlZP8jOreaOAXXKf9tG1lf179GKi
wMniVLOdT9guX222VanR4JS7rI88pKK3uab6vrVzb00Zev3xpzy0XoX4+FHnuUyZ
qCiNDJuRJpaY3KWyOzLgw8vJt/pJMskG2nMcLG/E2OGp3izgfpRJaM6TLQsbPunF
NeLdt/yjnbCFbWlzefyfOQgNtJK+baYVzdsnQmnAj7GuONIJIyj0GeALdK4vGvDu
8pyDbW7C33HitQzA0w4yOrt3WCjlRzntD1nQbgrWg5AZRFnLnyN25M1I6s8XDI6N
CwcBN2TVI+fzFroiH/wyrjAKS6U4JQUMZB3ZmtUFedBRaHl/LrvoAO7jXvQz1qE7
Pi9AW4foBO+eAfyl5qarWrTSWbDYEMSovT8hvHH1nCMnq/f0FX3vcZfWtnZUWxQL
JChPB+MyI7GSKcxQDtmeVrkUhfgm2dryKzVH3syBTlAIb6VnJ4+kAbT8hA4LfaXf
OaR/t/XlYctdAQDZFZVnSZ1nwF+yfOSRGMuHw9cvy9yDnZs8LOQCk7vZmX3MBL+R
ClHiEUqRYyQBF8h584i+Ht0bwo4VVxFWklpYa5qh3Rh2GucwGBh4p7e13PZviygn
TKZOrHRFtKvZpWFA473Vjb7oQ/todbA9eGV481qXn/+m+cMrMHKgRuKfC+qs9ON2
pnGb41YaEXsIAruakbBZ3397koPWsZa12GNdGGost9dLbcYk7a9C/Cc3ZLZN60JZ
1n3yKFxQj7WLJ9yicr0pc/DDNjFyB0LynmLPczhXJS6trC14Lj9Mk9U1ggT7sYik
ZSLYtk7Frvsg57OV0V9ppIjHpXtlQ7vLmgsoyMJp3Ed1XLvRd8m9+y4xSO/zV1KQ
t21PFwfHDNhPmlwPYFYVcnpoV2YJ2ktYPoHYk/DZXqCf7rUFRzqdrMHRcdRnZI8t
ZVgem8wGMIYvV0C1MZEPty7fBtBgY+3Hl6WOqhf2nZ5RjhZ+pxH5/yMPLBuQjD14
lvkA7BORNsmUTq8+b2AQAEU5UcZ5H2ugfMOv2fJ0BwM5mMWL6qo+bHbejeEnbfrZ
Oh7lW1RUDQzGrpOQfInsrtAD/uw2VFr7A7q7Gp8m8+8zDAul5qvJAOcwYozMf6Uh
swmj76QGPKEiEt6JHaTpn8eL7JEsNnH5hfbzJOOjfit3Dl0CIWueVFftTTLwtWUJ
mRnSBPbj0Ymc0Dv++FCW4LIqIzrlH6F3dXMGzgqLzisqXBPBjcwde+637yspsDMR
wANrfxRt5x8zKgCSJe7nZuAMoaY52sqg6e+Qwc30VCpKWLjNPPNKrlxuW9k0tgFn
scErZ2/rx0fOZYmcyf0jJzIyqeg+lrkndFPcyD5DeHfIFsruS4y1f6M++A0/sU/c
nXF8tZmgcbQSFXM0Ysyea1e+LeBWCRkp08KsGI3VGnq8S7wZEFwTCd10cPB3XTrg
ut148gKyiQrnYC73DAWLoISFd7s3WfQYwowHTbrp4eumF0rn+BalAyWwBKKsVujL
MDXjSXhyBHUJBgwbKchEr2j1opdCpzHfU8YybnCoAejEB3bcII9Icawl5yXptod0
xuvI9EtA0UL9haSHmcyC4PK4iXYvwBOfDj5VX4lPC+9131be7XeLtSq4LwfIuV/x
D0wFZ4H5Ndl1Eolez5wROa/AEBq/VyFWo8yy3BvnNqg/8agSQmLbfp0+EMrtSJim
dqKhMQBznN2GY2gwADylI0wHsKFgC5inQW1hGJ8Z1ovK+4/+sVdHzt/SqZLfiZMu
ck5peeTwE1RljA8CZUQp0lT/a7Q/fMGmjgGOokFrmE/FGsLHUFWjYegKZd7v1xBy
4/f/ouF1soMJGmXyhkSlXYNBLu/q8JGUwNZJMQb6yh/gvHxIHdByrLgFLECMHej+
fW1Sp4ulUG44XZy4JKCwAMLmUVNFhO5oHFGLyslPkK5/pHbz89xGNCLuOqeT6RXd
lMMwHeXr/QcW1zov6Sv470ZbzXSb1uc3A0SMz91B24hcHTJpSuk0S1ZbCzllz0I5
JO6+MEiI/eixi6F0n8LSM8m1eRZeUADP5xSsJrO87+KxhVFGv/GSAt3Df2y+6CQ3
Sno+NJgigKDg4QFqSqm0QNkI6viV/niHLc/U6HmXMsC0BgvA2CQQ0DnHZcxQairl
Cq5uVFMLa+Zok60LC/5Do2VraCdgKN/R5O5FljlWDbSZ5H4wjFCEmOzJT2LBCt0X
d/qVwlwtLAr5toWd7qKxlfhcUS8rARPRmgV9OmVR5ec66fox9q+lVZB6eD7bSNCJ
hWXlBmYjtJbhH5ZVdCqwip7W3Op9EUJC/A1BgQGX1OHJ4feSZhYMOONYoKa/CmnU
IJibPp8lk/Ci3BBGMdkvfCgGEEzICgXAE47Fd8DUxVGmG/yXRK79U+EfwQKEToxz
Z1qBpOpGJxr3Dj6HgxD8qDbU0oqLGuU/tYE4aqq/ouXgtJWa1fKQeKunYtccxMh+
XaSfmImfPGxChrW+a1V6KXoYw2YJUeI8R3HyR2MvsHF6y2ptl6TZfPx/7qFoHqBR
a5VDu2dO4QgUv6XWdkQh/0da2gbS+ccleS+PcFwgVk8OqN/puMN0SJON2bemTCRp
rzoIG9adsYZxfdwIj/eGST168NqtTHtdD3hloQMyzOP9PXk5Iq+gOjGHlOwPangS
O14BirluYIHtYtdTb1udWuNK7003OAjykYi002buGxkcvrlno8XAVdhP9FQoRgWa
1CY3PhHC5Yytjg0NZdtjwGzPNCNS58z1Ns/B+dr7K8cEhCNOnatWcpLtffv39mNS
0MeOzZ5fcVlnG0olOJBgjT1L4/Y56hm/7OcgYEJB1mKhIy3EhXozbNqCfAz929wM
64Jcx+oMzTnF4/cQUc46X9krrvUf5Th32mJqIJZx9N5I19a9EUBJR80rJ6M9heVT
OEKRDcWMmyRoB0spdBptfqEPrdNMSfFyj2L70VHW11YemkSKO0tAcvi91gC32CrA
hTFK5c92WKHSDTuNx2m1uJ55CHUGydDQWtV/3ICi0U+ozbaVZVFimOgkJqOn/YpZ
HRsP2z1uL89EYGAnxaBz1k4r+HBZvNMagVA1TuH9IlmmjmKwWwOoALVKVmaOOXNb
5YV2cPzAMdz6NSLs38n+W33N97LGW754FnCN8DkLtBIWvCP+SnbMnr14Wveh6t19
oWFI+wlI6H6k3+cv0sjdnr0f7dTo4g0PCQ7ULakBKB1zMdJ9UTQSl3OXNvQCVH7e
wVvGcQeI2xVBD82saTy21Sb4jQVA/S6uiau08L5q6Fp2LMwNhQ1nEX4C1upbnAE0
1w4ww3mxrVKGuFXAAS7mHrCVxT+WSoqrO2r7jSzhoW1wQvoWMGT2OGU3UsJ4ufjK
8b3BGUyh97qVmJlZISWP9oWj9Bw+gfl/YzVhqsOu7RFRzcUZRw1GkQ5S66YhMCDR
ONpowh3Zyl3W7dLjcw07djtyEytAEH+ExSLlzTby0uDPppB6XjlT5JaEwwYvum2g
gDopnjsI1l3I2fcXIkULfXZIesnzaznUdwYsRb0kLpQPHsB/Q+wjokQe/mu2uVe/
ynFU21hDd+LUgilXX7MdrK21RjGV+Un57uK4Y7A5p8IQHu/gH1uX3UI4q99SeVu3
ppnQPt9zPuowTlSCcUNufcfNoOViWxtMxJkH6/RSN09AEyfwyc41QzmC2zngDXcI
ijjfEcfWcW25/tEsMxkjZg6+sJN7QWQpGtNAGZ5bjNr8ur3u+utrqh67l+X5QjD5
NM7XpvhSaApK+PHv2YRzuJUN9JcBY5Otgw4TDKNWBoFbEcDORd7bhGhh+fR5LbgQ
efXMajAWBi8V74wuQhgRrCqfFjQfoSpUY6bKroycjWV6wfy4ybTej0BVqS0T1Q30
oVGyloke9OPnQD1BfCXnFle0I1sK3Gqy+oX+2FqBBiFmLfny6nqZkgWxliOl1OXX
LLdzB751+vSL/vzab6uIPQtfVOqaeVZ/BRbQbyNeVC789w4vS/yz6ahOQggnN0qc
1jpIrJComG6J1vHhTaTdpYLmTLYvpyyQQPwxH2VBDogJnQZ2c+WhegMP0EUa5d5Q
l2Km6Bb29awEHflz6t1eWSLyMz9hh8b9r9EjbtuRjIxlchZr4RTLsrVcJRtnH4At
O79w+O4upijQTlBtKHkYdQZOoXkf6dhPaAj+yxfeb1dZSwgfSls6NqY3X2UCGcY1
Wt11X9dQz5qHfFvi2ydIAmh02wnOiqYDusY8KP/AEnE7sI+xkiTF7zVK3xL4nh9T
sZcIx3izVixmeQEKdqp+rMu0SON9XVs6H9VNPX4AW6VsZXCe/AmxwCaNUrhfykgp
oRPEBk7EnplyXoGe17daHT/8Qfj0uB+/FLKl+ZjOD0WX1YT3ggLlcfdUyQs5N8+h
gUrp8M9o1YHTnc2+xKqoefiEDb5NoniqHEYg0u7bbVBRViloc3gr/viCjepLdo97
52yiV4BPlRThnsRNPvU7uHBTxFk6CtOrY0uN/8To68dixmm5j6RH/UpfHyOka/8T
dRkicj8siIaNIucD0xT493+pHQko739g2xf2+ZLpytHfg0kMowDCu2l/mL8qP2kr
0HEwsruj86KlQNsf2ImghuqgPTA7Nufe2NMe8KapD6JYO9zOk1hTn0ylv1rYCoeG
r8mC8RBzy3I9fgstgFHriS48PmR0kUirkK4Cg3jztN+sAsAwiZtLcFegLlZQ7i3m
cImr+NWC2s8/YZeTL6mLUay0yEwSRoiLM7w/GVmE8mTYGPgEY3aG1KmcT+1x4jDc
DVGKv8sawwal3EfG6aezkdVOKAj+ofu6WKlt+L8Dscowzq8kqvC/evTQLzaEhBH+
fmSIklcTflnRda8i9dkJPZbslFl86+l/M0k4FqMdt1oIQYHC/cOHhAHzAiHlXDwi
7mBLEjtW/UlZNbthSHJ79noJyn5WYW75Q8w8ChWbRxiclKuE/xO00io3MGmtNU7u
MUpTHDzngLWLio6NcR1BRHthwU1Q/eqDAdXvrt8rj6U2quMfmphFtYbvbXOZSWaO
Iu0jVlqYggKR95ZUDZFGoidj5NW0Fz9CifEfOPlNcDE7BrwJv9dYGbYqSKV0SObE
wbf0Ui4FY+Znadgr3F1FvzmFoksOGqVwu1d18gYKudpag6UQKYOH3qjPtHCbf7cg
KnqzQR+2ZYp0D0N6FdfJeJcwKLx9xp8JjmuV0k0+QM/uOtLgw6WyNgm5uDIFYOVP
w7ZjzBdpB97gMggbs1X8qExK0MuIOzUSJdZQuMHpeC0+2qcE82tGIIW08aQNG2T3
I3P32KnZVt2+jgl0v+l+s6aZl9Vaw0ZqA9FEz3D3LTL6Ya8ex0y4qlF6qR1KiLk6
L3Ln3q7r4KyQyhLJkBnlnPN/c9cJ86f+pyvgq+psbC84w93iYjVBqAw/39Z5/KRB
7R68KGZ86kUiYVu6S4KA4bnGFY/IAR7U32yEYKgyR6uiJA0EHNxtOHpVDTd9t32R
kbi/0FcvfazTMYzvEZRxjXPPfb3M+NKGmALLcmi1A1886vJHIs0Yrg6NtP+CXgH9
d1JG9LuGD2hGgYqar9E5dvxH+3v+HnrDANfLl4AZnG/2/gtT+ZfWL97mcYPvFYzO
JIWwXCjaGnSAS723ihO4tO+pMaz1QG9231vH0kACOxLTvHBjC3VXiHlyxG+4DRen
NRJbMBhJ2M/oTOVJyK/gFK5g79UbSgoBQ58ijGAl+pSj5QmTaTiyNuFyorvoxYkk
o9wnTy0OcaQLA/RM/PGkF4nvcjxeUcdZHWdhlHxgVQefSN+oOxoilUFKE9fsBbLO
lpyT3UigtjGZUjv2BhNY8v/NF94rex8MzrcvkndVMiwQ7i6whleZSQdw7p9AiCoN
3+LLTcs+UVAvf29qq5cK1YxKLAx4CmFh8YVJTcucHl5+jNrs37bX73wxKPCecAch
D3R1jIM784ky/q7mUiNtkDPOoqoJ1WqldS65ItG9PpAKvuzhfQURTw5Q3AEaDT3n
6NTFQPWUROxi4fE+0Hx5ru4a2x9fMJ5OcXVsE7Us7LaRT72zDq3OmyMS5sAWxP0T
XZ7I46HMDzzq4Q4fUSmePrz1VLoDzCiqUn921LEH3xNnScMe5noklR2fOng2sktD
nFl0KIPXhZJwmxxR7PWRuUvJ0Ot6aPzGu94CQhxHo/jWHLoZbuESPWpjiX2GBh+j
elV3oJJqh5NM/vvxuJmcGGuCFdWYM6SUKoEU7mc8xEnLQu5uHOk/COU9vWrm+TKC
Ki7anqRQZE0YzGayt5V38U0JX8oBshnPonZQPA96BMInWie916r9hQBBolPXLyPW
G8hlWXtBTXlUH1jdcwO4lUEc4NECQx3SlC/NuB5uQceCbuMwbeY7Kw/2GSLgwTyF
Bblsc1i4O4Ehz4mNZaAxDULRtM8ZL2Zt5UiFB9NZ3zdaIrLb4sM5hN8LO7FXaozK
a27SJWTK5Db4ZqSdb7MucL3zPPfr/mZAymqd59HnpwbGdBTvWrOxV971A9NQMunO
E+gp0cc54c6++eFHcqripSnKzKSZZv4Jic8+lor/AMEInhEKg7foo1NvErOIVv40
Rakbct3PzKHm2YMigdwzi7EaqaD1ngo65aD0ABrL7qI/VaPbBEEVDkRW5fv08yYa
MYtoTtSwm2I0iUaPSMLfd/KhqiDs/i+PdAUTHGfC4OMDuu1BVQqzDKFMq9PFYqwk
WdK4KQULYcynsJgfV6COwB/Wsc7HnCsA47F/LR2v5ePBICZBkt17nQlUDki5fEZR
QU2zKb+MSfLB0NJnEPlsWrEAufbszfhOfQE9e9YnfFXnxlmIxV8l63CW9tCYUDZM
TwzS7QD5T4xZ38P6439qumgUYzT67yI2Tn0L8JS48GnR2a8Iguc9Mxm/v/4RYAPu
PQ1fBpiZGQUBUGjHtN77ysNgyR9fQi8cMF2NBwQJF0+InavR95Hfnu4mdlpIAF7b
/xH2Yej7JRkqNQBSeaHH+fZaGU1/+5rxOt1rdM+HjqQ8qICxsHht1q3eQi2yOK8o
gqUnYLGPXEoYKNc2raqMf0oyVR0/lYs7njePW/UwskZlSjbsFoQYepFl2Lsh4aPj
/4PHti4KygSmueppndsZXhue7HvuRvvA5w4sBIwUkWwTtSAhD8lFThY1rY/BPsDo
+JqWPaIthSfKXHZsfP1kBhiTqe3xVvkfUSqnHHfBbwlalUTF8ty6OkMlk5HxODxl
YmExNBEUusOo+/awlaEMFQwmzSGGw7CYqCbcX7Nh3d3Aq3HfCDwJ4TzXVUPsR3yS
U0jy3vLcZCG/wBFYkVBpqdHz7sRf8QxdGs+rwZA1kutf4ye0unfKOR0P0rDPTAur
5LjV8JqnJVPUkFL4Rf3c3yeGf9Ljjt+cL7oofni7nemIr4SySIN46K2dMWWu1w5b
5I0jiVmApinpZ1zzynan4O2IDYvmNAE2V2ptmYqoxl3G/K+Z+PR9Sfd691E+fNac
rv3qSzjbY0voXD184MCxTvwcJzRWoM4fbXv1axl3vf4H/0W5PMCqtEf+qDip34gC
KhAnUb+WoRuwotNMA3UjuOp3/zaaMaunT4Hb9sh1vt85en5+M4kqXNucUbDVGJFB
tYBBra39W3qUantmF3d2TdpreYcQmAHiEnoMaNHu0LZ4wiv2kUcPxoJxsA/diDPk
DjQPPxAGJWhe9Js+Bw3WWl5CieROQSpPtXUnzagCdhdiAP06qbNQSs4iWIaUUrZ1
EuPU9r9ltPGMnxUCWhO/uKew3pXYHa0R6yWsjYxE9X7g/e1KoSDC0LLsM1DLkUGC
mMVD36rsUJr0iwN768rLRjqiCU4WDQAd/3AAYp91JHqiySoufpGc02faMOOY6Exa
Rw7R5om6ZFXQt2fJu72ueJRiGIfS9utnNvqn3PVY8TASX3hcj9T78ppXVrUOj5+T
CZtkVaqo6RgWGLBgvABsJoJTr36L+8AdemSbQmp/MTtzr6IO0uhFUDeAg+gmR8Fz
EdBFGn0J7svPTUoiDVWu1FrI0vGqtmrUOaiScgLzyNj1ldavkEIMbG2MqkFM/mnz
v/K0xwWGuB5cDSU5zJRrowwAreZATqr+x+m50B1NuQcYafcRY4daqA1b7pwfC5Fv
ND3LAC646BZDEO2tjj4pXnXaQ2T4Cpi092p2vTKazBV6WVZKGC5aQXia6cc0psEH
PvOePNctQGmVDPaXz0gSIAquqfQeOkYlMiJf4dhdcLFQycpZxbDCfpm4ehhRfl6k
YuJSOJZbPs9Al4nYRKFItu8JWtcE7ChX6wdRlBnrvKsfifffMeiiv7KI3yy07bRm
WrmwN01T2evsgYOjHQsx3oai+QZ8rPSa0hGycujLxlE8SyiNqQCreLdrpnIwhhl6
+/TspNsXnk2/uwDRYXWr6e3Bn+YiC8xux6ulogApwDd5QR7d0tgiP1wgUkVAK1pt
V3sunVLP0vuuYytOzbHGjoPQ7bBZQ7YAyYAzY9rBwEhxelBMTe51H8F+p81bvuZE
wfqNTGBCLEnLOfOXljqECy8WQV9TcIT1ifqoWxgET3TWz5VxXqsi20tycna0Jpva
YM+kZBIkqFCu9XERIr7xQk2Hqt6/pM50bULVB14NTjjguCzkB4Nf6I0+WgKG2GVL
O6lwYtYLl4O6EmSA1bySHxwxSOoy6SmyZOnL+mTe2hbIWtn3xjO0u3EraH9EvlwQ
rz13aIm8BodqBgrLzLQF6EBo9s8Gx4UrfqdAavTXZQ/QDra7SESqQZfQgqrqRm4h
akISD8LIqaijmyiTDHADjS0/b45JppZxgWQyqrcF25BtunUg30SEWfQiWmVB5BT2
7Wi039c57pURWlcdLWU31+lcCcfIV7BcjSYzPblJhzZJq95BgMnlWSzJSYU1xe08
tTtQHQrbGbvrZ1fIvzJrxnfQdbYlCPZxTMhXs8dJw6HhDGUHEi0tT6rYonBdpr+l
ELIgzje9ReD+jnCyUv+KOjvHtZs87LRR3eqN4Zw5BGx3JC65Ts1OHtCUCqHrCMMj
ieAJVMjEA2Q7r2vbL/N3ie1Nw2Xv8zNnNJ9aVuKva3G3Yu5NTEiYukoAxvRkf302
WCS1P/+/OguevNT2UAWtWLMxChSIOvUJ0wP8sIhxweO80BozCF7TysL+H20fP6eG
HCeaJBQ7CC2Clpw35pzqLjcM2ZoVlH574b4CCVJn5J9KpHPCs9imE24oOg38esSz
6yl7zQWSX8WtNR9Yr3V9ygFbeVcVKUrgJLEC6xPuNgZAvJI/qikLSfYxZ+231Yee
b7aWlahatP4xPkRFh1MyG45J/7FW9LmjTDh+x/Qxi544vFTSmiBlaKWkukGC2k9R
DeAPk5X3uRmgbuvu84+MttsfZLgkBODonAGTDyCOSF9zafcwdbDSb4ZFK9AQ2+fP
bEAIhf6+yUxepbwNpaaZtT04avVxyW0l1C27n3u6K2oLyKKIwHl6BfPRv2P+orwb
p9lUWCzgDkabiELHqEVbbmyOTNcVMoFZBAneXgicavNQ1W0+TfcM3AtwZhJreHF1
ITqrNDELqU3suXNIxRn09s29thLTk1Gld5i9+atl6rk2L+52EP80toBNls9ZnFb2
YW8zHbtctnAGc8Z7R5AvDmB0x+EjYP61pq9S/pXYrtJnX7AnOTbL5IJ6845YLgVc
Gl92mopmlD7qHsIyKGVAUutFl0gBWZrTbGi/mmPHBvREuQvsEJXR5wx5wesUef80
a6osfwcRI8tM5iZOl+U3ODqa3dq8CSZ5zuDdiuzSNzBNUR8b0wg0Azn4ZCR0mBL8
/lhcfuC6edPdSIm5tklivP5CPmUwbLecIp54S+Dz2n72zeUnnS+TET3GyrYLQEUq
+3uZdpnmKeXNqYXRH6ZPtnwX85vu/LCmNcNqTvUirP8wJRqlPKdNQr0K7jQsCQiV
CR/713Hzy4CiZLwwbQ3hwyo4sqVvZnTxbBugOdlOpQL0M87PUTQ+EaNa5eI/4G8a
tLlxhVK+1mvAcct6SAGfBt2DYYoOK/1zfEQuKmHMbCtijkgxcS01EjP9F1D4E9pW
zMzrlkaeC4+R5ogwu26v96kL8Fj8VXWC1z6Lq+SgDs8HVc1LOuH/E5vFdYGKU/AB
bfnK1aToeNaLoyVWuqoWQ4sWjkDOTlQuqurEFKkblBHVzT/PXlo8HJ7A9rrh5Jv6
nbTnn6A8gsOlMBsgFE6zWekrcsKAjDPr0QHjVM5z2EjhYuPQyUA5N24+Hq//uJ+A
mFd0XTRdUPCHwB5++LlFC/HkAqiA5hBqaxorDdrRvGm0KlTo2q6p9zORrqoLFert
kXTN75ZCMCkeGh4iV/Y01VB4pOFyCpSq6oI+9vYnrA8cy2bKz6f/fsmyzQkYQvMA
hBkgkPcc0YqsDQLCUj0fxW13N+E5CzNZsuTZtlmZ05XvnNgXvXWQUiHyyLmKTyUV
wGcqD2SaIHIGBApkHkj1cG6nczqn/lxAeFuic8V72xjeRLNTwsKNKuqAFvL8/y7b
b9p5DU4XyfEyV29lGp70ynDmaH6fQPZWuwQAC56z1Gykmo/iNPlfJQqVRA/EZILJ
M7xMo6iUu8kYack9veRQQryXcWPEjl3KmgNF67WRLSgtSLMJuhCm5hmbLQVoMpBW
TPMfcP1UOh4e06oYifzaG2ZlP2Dh79mshgSTa5M7cxa+q7XqojlBV7bcnkdhNqQO
NISlddXKDM/hvrOGAQWwN0jT7zl3ucjSx3NpO3zSJHrYc7eTYccsi+boTWORgFBU
hYCldncjPnrg+hzIacjBQlbS8cA46DLpnz5Nb0LV/RImEdT5v9SmdVbAGTgATHTt
T3Dh96rKmN3lQmIqqsXo//imFQ2tlUf+K48iLnxQi8wOL5Wgg7qlk7buBwjFoDwe
IDjSl4jnjjfEAB0Q6rLotXIqIKj5dSGAfUqqqON8Um7v/40M7goo4vTV90qBMJ5U
vLrnCkD2mobGxCPehalqqemokkD2tdMPxhXTyGJAcuTRFUos5DM7X/2IXIsrWhzp
EO5zxu6nrZyqPZ/Wxh7xBwHvqnl8aJfLhbF+qHj9SBnSkn9C30dAdMZl8HK+P3IH
EjzQu41kx+YpKOejn/QzVdu06OIid6Xg6Fruithxat25R3Qq4wYfNh9qqDurnZgb
BWVD8TF4TrLwBGe0SA5LvNYjaFBhf2QPKZGUz3jd5o+pkeWMgLIo6/ClpsdfeFQC
Tb4UyTBLGyrGPddUdxYSPqjNuURiMpXG7vr5KFWRQT8npLNtR4SO77QwwOuJXtFQ
+Jr/YOv0AH4E0XaW5J7Ylis/KG7nulK0qqTMsMAyFesS/EeTMrrLJ1kXLU8zM6FK
2OD8K2GrXTC2HChGIzm5w2buMqxdLihgBZJ4IeKKNExzQmc721cMYY0JIRn24HI8
0nwFkYLluEccrvZ5FjcGDA57Nv7jCm9FBItxtVZjjlTD5JR5YDI/Nf5UjHmvG1de
G5/otuT1dZ88NRmJ4aLYOAcbum3XcgL1TY3VyWxFHzmYIpHR9uQ6vXKZB1uuSW2R
H3mg2j999jkiAZs52q28C7mAgjtt/frPNn9V84rmvIrBz+v/A6XLyhcuzXjgIfrs
MZUqUY8IFSVPGpuCjVoepYr4oyPtMtPvh9h+UOXRltqpv/4WZXyiOhslJ0lB852N
+RurYSqO+dsGv7pvi/UmVYrLJqDUmE1nwttXIMAC0kvojqx9OxRJ+Nn1WAHxKtXx
YilCt2NTqox9e0wz0+paiHkyuahJZY/Zu+YFbISTbgrMLZ4m8R0gHkmpg7bHRlMe
25o39pSyPgH6WSwvYSxggfj32N59MxZTTken7vYsvqgU3LFteTWehpCbO3Z4j8Xj
3FeBV5i2/Ii+NFzIkeF31WmGIxl2SMrVTOAF6ufcvXb6GpQpvvR09TScH5nf0qBw
ne15dNoty3XJzjkzx1yPC6WMopGAHnzfLDD6VIcCecoEUfrYGboA8xOvP6tWPHMQ
USWpLA805sQQGblAxFmtf17RRHXcNOyFSB86ziqWNbcgndxTUP8FhV8Gw/SCeBmd
l+N8rTL0ViZyskYp6njafyjaZE4aWvoHYHk15DkJPFMFdZbA6/71tZZzGRnK1FJf
4xCQtTKfFtMY+9umhKDKYZdVccXi9Dsl774Q+c249lUj8UxaF89zMX/Zt+H2YJ8R
i8mAkA9doHGdTy9igLZ+qoc5TYVbVqd3X1WWkdxhHubSWj/GlQtHDooZR/ObKozU
CTg1IKFOLdEqKN7SWI4P3A6OH3egHPrESl02Bsfz3NKEZJrNEsfZzVkYwJWl/bIf
gtm1ctu1ZjJm2wbMIA80N9J3bnJ4xJ7e5kxF0uUTXkjufPDgg4ZMzYB9lvrttOXJ
3uGhvHDu8yQAzZ4IDKKMVIxC3z5+Hx6NWvzNoyw2Tkeu8XoaOy/vqaAYN41fSC53
ve2QpcihG00abGTT1bMOzuN+MhhwoGl6fsYJKHTWr4Vv4gmMv4QXwX4TF9SDw3hX
de9IZm61joXNzjK2X80N9BuisdW017K4FPIP2qxuYu8tJSGV7qMKk7xjJAuybOmV
gvhK1UXxljBN9fuKXHcfcidmzEfLD1Vg+QCigjrE3EVquQ8uUi9M06N/ItowaJbM
BMNy2aAHTIXm5nSbrdKBjYmRcd4FkcXk+vpPE05iAIqcKt6/fpeZdBP3cX80RCrD
VDNCzFFtYHM3dlRON8lpHMAdQ/4lhqu6RQtKiPDkUQ3CRe1lhj2TNpNp2VyNGeQZ
tV3gPooVgjPRwrxQIeB7al4ip2ApXynyNvXW0Q6R8qN/sGOZnt1ej7UZLBgnZwZC
gNhu/tz69P9c70iErrewH/9o3Nzyr9hrcT9GF1mGZeQNz/+T99T76FkgDOJ6g5xf
MkdrR3Q603Bini8NspJGjlvsMPfExVSSsl6co7O6QxLb4Vw35u4Ryr4X4tpmsiiD
BUHGdMuwDVPoJaER6gMw57dqJgE2q5tx5h/GKXb0sDhJMF362+KjX2gTimcjhfNJ
9jqOJJ6vFI5a2uTaiiPwM5xjiumbreP5WfJgXv92T0J8Yja2trqjdGzdAcuyOsXd
aEeLk+/qSOwTotqXg/22ChS/Qcw90oS2mNlAtTyR2cmDWjTe61F/4ccp7bJMwD1+
0M4IbUaNB6EnZEteL/xfyvogoItDxOE+re5R3t6kY69tDCCWaMPlh7rJ5Aww0nx+
OVGmPPW5pFdZ+LLLE0rNyRWBJfMWGGRhVMh6JFDz4z0CFOFrhKt2ZGaJcCwau3VW
CNuJXfXgO/vTkVzKUKp+/wZ+r7A6k7pKXI+YAGrGK9izTYkHSxo0zfdBMe4LTLqB
MTDap20CpYJConOair2k5mcvfQSITWkSN4qKADgoXEeQQm7BkVBRPmXZrC8UsXWd
Blew0H5iN74lwJLJxzdPGxxSic2iIV5h29T7mXuOGITx9KgzNF+SdCu43srIVy3l
A+Fi5i9KTVict1qKIE3Vu5ygn13lpsyxe4eaOkAACsjIm9CgZoiJTfIKm6yNF8oX
elI5rm+OwrvVNHEzwVy04eFwopURBTdbBGkYwDbl8MaTWdifYkhayoIWLi6GOYrt
i2+iJ7AhVotA4GvNef8QRg1GlE06RQvvO6uCPqtwq+16o6Vyt7N95swW41fjKoYZ
jk2x3BaH8xOSAJGDPLcBRNPEkgYD2bv8nfMrtQpyzgR+R8cY/dM5+KCSvm88yX4I
RdMpMR8kJfai8dxoZTkFCV6v6C+PVF48C/EhxIse5sQdpyuru8l9VVHUQuyiCax5
dqAsOYC/WodipMvPH8eNDaEMEhtSdnWAHT40vzCEVaFTNGdYF47NWQfGHIIZOUaw
A7n7s1HZu6EtSe0Iq4K4sf+CGPYJHZfKz4Z+F5Hj1A5Xxmyp98r2j3ARu8wQUXi6
gjLGBh4hGAyCuo0y7YbSSjT1kOaFVBN/IVgmAT2Eu8eW2p5W7Z5LvttFiemleB4s
dFgX+Uf42eMVe+weOk9nIdMvW8iCzXQgwMVWSoyggmHT6MtSz6gG/Qj4GvbGuVaU
5tAzhwVrCveNtB/kUQhPzl3xa4ydFTVbBph0yfJNqXRJSJC46oMmP6xG+w6bhg/M
PzAHcjX390+GL8h/ObSToyyZ70PVUcVHauuyePk77tCwZt3rScXcUDttzte9eDrB
bgxMQHKW25xs65OAl+px33Nisfm9Ysxw8k05YnOO0q7x9o43cXLDNj5hRzdOFHIV
1ootKVYGfNqSVlbv7b8HzOlNOEAqkjGFh4NpZA3pfJ838e3DASnmIg0SkJ7woGGg
GfCQDM4KH3P3Eh2jRgcSisyPreBhi7vcqEvAMSj1vDFKY2U3HtLffqKQXJq2hLjA
ejy8/q6AwaVnFhLKx+rJrH7keTvWvYEGBJhM+HW1mnA81Wy/UmilDqh2at1LLOgS
Ic5S8tpr1/IlVa5yNsl+5idXL65cDbO8S92KNdnnEPHVts/8okI9tOfJwNT2n79s
nnYchVL4NSUSndiZHmZMYr0z2R9ffqT47B4j8mx1aFrQkrKUFq1ZQPpyHNbflQvY
NQh1Yu4LXE3aRSr6tCNY4m6kvjiXCYUkw6EysJbBiXznkgOy9gNq9lAzfD06VOk9
OXkI/ZyJxm6pmmnxttnfXWJoMdXpu6NQs4HwB+VXdQMhcwIi0hA5e6J2Arl8VUrO
D7o4rfGPyNiWW/+PMzYInJG6MECzxbdw8HtTiJNhWHgoMh71CGmy6nz0ORXCkiVB
bmF+ZuAov3TAtbwl2wryV0HWWqPzIwrOb9YGt3ZS25hkiFH36Ld9Cjy6wV0xtzFK
+qLhIMPm7YQKXirl1U3WFfZN+gAhovCPil3DgLeahVEHBTUfjkdnASGXfYZKpCNh
V8fuMScHhLHOEpps0ASSVSXARcUkotMTs8kzbllJaQRIGcnufr9SteLAUGOluuGL
ZDPL+g5C5/hNnfuHCUVvtrajYGWV0RlIq/9O8JfZSuJ4fEL+ury0AhM58w4v1IHn
6AzZfaekFN78J8d/631bpO02Wbabvbl8hYt7ur6KoEg5Rbu4J/GzL571iVi60C7b
LNh/nRUgCejlssk+X6NLeSbP+/0JHy/94c0YH/HUPO7rIkThtqu/ehwA+Gyds5r5
eads65Erg01oqyouVGJfe2K05Whj38lW5YcT14QM3orE1IPknpA9uOLkjst1crYI
zGuFHYahzZcO9ZXbKZiLK87n0yRWDoA9W8QPjLP4GjQ3m3xhniEp+/dNlW0NG+9j
n6to1rAObJOLByghNTMfz15awTA3AgS3SmMm1hwHLNXeeQrRhrrZp7rvZpflElYz
PB7/jgGSUQsMDZPovaEURwrMe+ZYr1FUMueF0wnn3j0m6ac6IrbutWgjo547EJmv
FgM1ySYWPzt1SoXYp2zgkiQlDYVl2Px0oPq1at6vtLtJoZf7ox3kCnSNPoPrFhc6
v9HKZiZlmFTp0ASNaliki/gxJJoq1x6hqQP0pM1rxSMQg7B9htTdnUDLby1c3JNt
C3+ujosMBWZpeD7K+AFSjDSlrIaXzoHKK5gkEY4pQat/ZicLs8UdV7n5E4wqjkI9
7qHlmIUlyRaqxMDxvM80ITkCVsnb6oK+Gw/U8psGiMDiXmHUKnsEFv8sscp4rRQC
rytY2NIJh/hzvekBakYXLniNmCLHm4OjxQk2yuGdA2OBJo5ILQzl/w8e5FfoFnr0
xmZixhVl2a7dC+Qhi7qp5lTvHGNoHLo2X5JKP+izXM9UEMOGZ77Fsdfstw4UN1/8
KsNF2MwS0XlstGVXm4vL8Bw8dpC3mUBShda5Xjq3lB/5sCQd3J2Xkxf1cv3W90Ts
JCnYrGEfA5VXKPVrHebfLUfP0e+HIKWO0+lz9RlCJGJcEOkHzr9Sdhp008KMvS5B
d3/zXoJoxNw9UJMT5uJkBBCUbQCTS63bVIvlemvP6QJmFGSraFKXGlkClRsts+V6
LBVmP8XwayyqXk3qDL9387eW3A5NlLq6xbSW5eE0RMOpPrdAHGBOUN+FQcFHCB8e
sPZUuLv1Om8QpQrVu/uaxq5FmrgetFqHwG6wsazYI2QjiBqCYzdTj5byNX9am6fh
YqiyQEJ2VZslxbwNulpGtQVwcEyfARSHVQN2u2UUGqFRCPIFhCpvJkj9xSj6Kr/P
6CXhuBdcsjRnTIww6YCFu7WfRKHxuE7lfyv3T1bvhZlTj1KOfDKaeONo3gE6f0lg
SFxIieq/vZNCiA1GN6q4pXnFEAoVx6PjQt0vQRfayk6zD58fD3t3CSv0aeyLbgxx
xdV/M87wzFNQ8IPRs/E/xAJVl+ZKcAfFVAxTlzgDfWz0IpVlkK73QrhPznT/p8BU
gh8ey745sNc/Up6duKgRIltv+ok5AppaTET2CQtHie1AD8SAqvsENAHooSFaNAJh
OVEQYMLFPMJkxgMz6KAhrexK+ut/MhXd3ajc+zKzzXYqY/29bilaWBLBP6oI85D+
uRzLpmS8C5MCwfPA4j+fFAiSK0pSfwUfOpIQuNcXufEkJjSduQJY92nY6cD/aEez
jIuZND8sLZnh7UxwEIR+HJxgUpEBPUvkX7jOQ2027GVOWPiASZ7HgETz99TT0pgP
DjtFsGcKMljdnUrbm/iejfl5Z0rE/Zi63aUh3DGch3o3DTmhrSHxbMTZ8ayzoUwH
F5c6vGiDLkud/7e2ZDr9Az5/ESatXflhpWna8U5Q76TqoGgqHyn6comLI2+Vm1so
mEx1zT1WoGOVAFmRZ3FZcWdgyEh8POek1W66r1PyUaGO+wI4wakxfc+tqv8lcqXW
ko4o/QwUJ8uqiRD+Ym8sZAV4Q/ZOlFe0A/DIc2a3GgQVKpf4RK2zB3V9V01t95bk
t6Hh9K79UPKnUJwcdEvbu0Zet37BN5Gv376WMhORCiC9v2SWmFnMbOgIsSjTuXtY
RNUJM8MHwFwbVw3yO9OA/0A9v0XtjWYnbJzT2lCzunqgVKUhD6c3UUhFzjVW7f0J
oCg2+vjNhvZL+Wxy0g+A3Ibl7Xlp9sRZT+ZhncRPctkXNec78ShxJGgUTj08UKVp
Az0qIeMVNl56fr61/HLF/0FiDP3zBRtLb+JDc8a/++QMw+3F0oJDSFV/1HKothKO
MZxOV9LK//0HckLdVsFfxLlwukopoFSAJEfSSVG8BQKV8kx8Bst4e//KI86D56Vr
aUFpc4r0rT6BKKLOJxDc3Xdh1k5kFumGF6ClRYM76ibOJjyxgFTEUfX8cMUzoppO
Sw9HQdtpfEMOqe0DOzN784bzSN0zIc0W11M3JkkwQ3PkWlC+hgObZUdPRnu7v8rY
B68S+pEBJhSAg4FIAxHbTGZKeY3oe2Z5WVxCRA04LwI+4RR7YY/Ez0bn8IbFW5kh
nysd0f7ius1peyF3/qCgAww0f+PPUELUhJafuY3+HUZxrpvZQjWGSXYSl2/Dou/c
JBRQIZ5mwox6qf7YIa+9ugkuy871jf7m+TdqwuA1XkK5JbkqDIPZHGzneSfbaBrp
zw/yyGgL1w8yRrdf2ZXy4pPKzqMhPB6UhlKeqGpoGSPmIf3G9CpKeR4n6ydHN++u
u/FiSB/dChoEP7lYSbFLKja54WqaZlyhKDtZhmKLDOEiw3X8DxnULfNGYylqCi4G
IgdL7K1CQHtNjsvGcezZgkD714JjHaMfPpNQFlI0GSw/KyVQSJC9awzCdzAMl5rJ
RsVoS6NBzAf4Ipf1hRa3+8GEbaxMiag2mdrThVYXeHk/fShfGBuacDVBODs36BNi
/gznn14gGGKBnign5xyNS4xN7rVrOV2YH1CHyK0qhpUuOltqJ4iW2bFuxYM5jtsn
eqmxJKU2OwSNGEdk0NlLaL4l2BEeqRr+sFvSbyaXwqmMkQpPkmrdheNbTk7A0d9v
oT4aMfyo3DlvQx/Nn+GKvpjQBbAHZcv9qeBFk7uTWyBYWexeHShF9ZGcDKcHtDHk
t2f+wv7LImldcchhTXR8FJVkwV7V1pnfeugwDQHijuRqHI8R9+JJOD7G9vTqATlo
9JIEJ1TBpmiyAZooGlyq6XL73H5DTNgStY8pb0lFgqHqgJCGhNeYtqyUK0PygaXm
YdvkHDkEkGKF49o0A6cvpmtPNf2GArHdmCLk+hvApECwp6fVdGtt1xhbLDLROHmL
wzLnQHKGz4jAxvJ1nsKZzMhc25sTYBIDpuY+l9ZTugcxrbJbiWEIKX+xcGLDdJOh
FKsw0sgFKqTzBJ/u3b6uLxewHI29b3OgoVuv6gWNHDI3z17tulzN/RiLG+uPt1nf
IpQax/ituIiZ9l8rX0NTpmc53PiwwqgFyu4Do0luK7fYk93v80s5x2PE84vWI5aM
inTl8sNBi++oxexGZD5oDn1/SBo2YC0YpPF3qLQ8AFEaokRG1YIgUEeL52C53Sjx
8Z0L/1xG11lRz+fVdgsctcHkOjc23RnVZpwMPDASQ+zCDWNXPeOW8dj2XEVTT+6f
iBXeD6Js4VtomGttFkkcShqlhPT/OeKBH5D85uQJ+FCWvzIGi3r5aki80ti8V2iz
UM/PcSCmPjX3btsoJt4pbCgicGJkpRChuDCvZJWnSmLYnNRkF/g5X7QwGyucFwhD
Sh3KgtVimiGLbl+oUQESkTfl9STlHH34yZxoX4dTchgQOkABvHUAJ484uj0fcr5d
5VZo8pjENM9YqIOyZh26KbBBkseyaZ94EHM8r22861xB44mTKtsUn+SfJmjEHOis
h01ZzpkrF5bT5W1ipuEjMXsGgKWW74Lpahinm4RN4oO/7kkUIzY+39SnfQITWsmM
Po7jGK0Ok/jQXCs4Fyd4hPosmDLmOmAdR7SWL1mvSXCUZlmRF0qP+zAmcqQm1v+e
ZxHXyruYP/6NGq0M4TUsJNeIuO6CDh1R+E/XAaahKq0ZLhY8zyGj2/77po8ba9ZS
DArWKbk64fkmflfznZk5RtysFa3CLKzXR5MxeN7KLnDZRzgZPsu5jSQ0rdVYlEo9
+i4jG3cN45hYzDogqIM73MHQnD5SJl0v4iZ1WdB3PMSO17oegMiHlTfAjuiXLxyo
fPaCTUq3kQcrgG2G1Gjlt4lN4h7KL8d3tjdAUq3XnAlvuvEa5VPa3vUKoFWd4/MQ
zZz2I/q5fi08EMXS/00fvmLulEJa7i2zG3/zeME5GGBJG3H+4ilXYpVI6LrTxmGM
nVB86zw1dJcXVc/bcrURPY/olL20/NNNUhrz8SM028SSb5Ksi4bmmKtLBx6mdKC+
R4hwUc4hMVSvEuINFyDJv2qMnFt12QuYVK0smcQAmvjrp0mEJDy036Ynfhbvu11q
iSneS2UvesSKxoIEI4Uogg6Yz1rwaitPXn5I50bWqB6hCXPWjWmI1vZgKg6Rsu2D
GDNoVATIRTLBnzgo6zvLHzx44Ev9HaKCCcUsYEuLZfdQryqKtPEQ+yIuj/HwbmhS
TP4fh8F061ofQzwYWPjWvGdI4Pp/xBS5foPHYX124PD/xsQg81vUVsN0hQZZQPUq
HFXIZmog7qp8QbIn6WWD4OzSI7TG+9+VeN5h8zdX8w76QNmSfheZw4GFAavvhR9Z
xqMVOXpYru4d6nkfYocZlzxvLrmmMnMsCXfhlm5IXAuIbtWMlxQ8uoaOdtIl4B+v
j4ZDTEd+TV5WR8Rur6hmi3XEslBD3FMbFTsTciMffqNA/MXQyz76KrXoEHkVNUF+
nII3vqjTkueuXWSKoq8F7gq14pFSCiTvWiOBXKal5gnFmsvq3v4yT+2VWkhMCGgV
25IsvegJKgsfxn5LrZGCQ9oAO0om3f5XbF/HRKs2GxkTBglg1dQMhRvzNr13SdV2
d7QPzAfSeKj0WvNSp8jwUkfgrSz0TlVs8CRyOjxdXzhDf14Lmh+lB+JsQVEEVh3w
mlj3yK988qArWgSoa/JRJjP2Q+35wVb1JdSD4yi+apw7ajcyNX2ohOpbwdq6N7cJ
q2wmlhBwpya5DmOw2ZcLnkSS6IlMtqEwVAaoNTGcPz7/ffpBhILdtPJI113wjQYw
Y1orQqXQbNhe05xWCG2V/gIKWLVBp9iMw8ttZdmaw9971nJmqVVZ40ZfSSiDg8+C
4BDgLLSJgehv2os9pIGYUPE5/Xbtj6cwhyKhPHG0M5shyHZkRKJX8KQzC1IryI2h
PU6zFMToUUsdkXY1LcN1IDoob720ZLUz1zbuDezVc7yMc2zpErOYRnhQe02TX8PV
DeJsFJcHca1Nd4Z/FusKKHiCyie6wV/VpC3RtQM0BTEqZPMJcwsP8AFC+C7lQ9Jf
WkDtVCAZw1MSoZ0LteGYhF932vKarsY+UhIKd1QCi0AoJvhqma8Qyh9KjZ7r9ixh
VyblWCBneds8FNKibRAUYQvXsaN4JhhruEHl0MK8xNEkctrulqj5ukCbq8Qt7OKY
as0I1uMfTOEsCoedHBL34T+lToDb1yfC58j3WtVDR7uPUYdQTwThWhIYk695p0gq
PTct7XHvWa2jNr+SXExulD8hsSiZQpV/Z6s37ZmMds7bwshXD+klOOrp/WqjqtLq
wnkI1ZqUBGKnorIFA0ZKGK5RaWujnrDIBRat8y3G6eiLK9dOkFJMxGrbMujJhmBl
5I3ovi9fo8g6HIvgtwCJyOMW66urCs0T9H7DF6lIQhfMSC3ydz5pH55WLG3Gb+LE
Dca6uY5LDhiXEJdQIcDTaqhAe3nCJ6gS++WbwhS/tGFk1f869hfa4Gz7HsfniHYz
wkc6w+jqePx4BKx2nepDNWT0nCVwzUFU1wYOGiVXk6wy0yoSLq9e/x7I1PRODBC/
Z5YAUObNwzY8W6j9L3e8KomkAH/Wcm5HFQ2J+i2J9aZPn224cYU+YZlv5TE4zlA6
e1RDrV3sGGh510R0/DwOrUeot1kX9npvS1E+/yzDWqTVtrg0lN5i+L1kUEGcC98t
bSXfuozSXWX8ZDZ2EQxb3hwyOfRL2tVsJGWvidDvLXQmgHdViB9Dzvxp1d9KUnOp
9OmxDIHCrHcwHdSeCPsoDSC+le6Exo5yCH9wDpsbT6mlI151OLArJrxitXy4ojWj
0egPU+TYS8pRUvFu2gPdS+KPYV8c/+hmnlD3I0XmxWJ3L0V4eSUz+mdkUN2frX5n
ZI1v2PhMGXCoyBAZwfR2HPOFW0yXDBNMGXIjXjJqfQot1nmpn3hbUBCEHTzkIVt+
PLCHpAs9qXxiVo5Ppj1PRrosBA0R14MC43VL6zBeFBAoQ2RjYOWx9fj1Wz+dcQJD
83l4f9Kih0P2UNV9f8bNXgr6qn45L8mwlaKiGdDxW+TZ8krZPQlcoYhb+AAejica
n3MAOXmOyQuyyugsdT3efwCt1WCaMP/GRl8bW5KerN+Xs4DDRUM3xPh82HMkOua5
jQmSNiwQvHT/MqDxNVGHGzHvINR2yD6T4su7eExigLfkeDgUKC+egR8zKex6vz6C
0CGyJSkcyRqq6m2NyE9Kz44o8w7OffkixF4b+RsTycVZNsp7f1qVcgQLvqZMiTUn
6C3x12KQ/7kDAa+rLRncUtxv9PnEMSkiRznZE4Jt3KQBew3j5HPIq1B5jJg7amTw
KsjuDrjGygCb15Bgo5VB3JwMRw0q5bX+6dtJ9aHle/IjQzDoLV9MXedJbWEQe+Z+
Lsf1EQyyyopQtxKBH+tuBUkkd0ZCtTpQQWA34CXa4K7afCYrJRocxz/VO/TvWqlZ
RMxg1HftKYHDRaQbdJEVL4LfqIbjZ4rcOoy7q91RW6vom6PAccMRIbfxMJRcLBJM
f9ZXp8ki/gWs/CHAqo5kaBOeUZGw92mVPppQGk/+tzXRVSIXL/VhypV+r4+r/vFH
aHgGiDziVCXMbdLrPlCedzIW6Qx96kITiH4mOYMntGwizSyg0NhTUpA35tDjnwLg
bX5/AoC/2/4NcA2OAPeOPSOFittpHVp0sAi+N4HO3kPUlrSAhlUZ80E00khSyr8o
C9e/UW3yaQdaYOJ3MLbid6kbTUy1VhLrll8JbvhaMbODnalJgGOohKOvZIjmEykR
LZuAsIw8wxh3nWrJ5ce5GJNaLDuV6UoWBhheONc5/yF/rjsQ9jmnLvRZ1YflfCE4
NCqTWrgjjgcQ8VPx5ZykD5/iAwnc+JBYH9QUmuleVB5NguXfLSCqWwAX97x6tT0w
UNA57jXS+UFvie5A+vWpDpG2fnVuUeKiFaX2VGO4s5jFE2rUnYWvwzgqMYVuH96F
wK5yMBj95IEumO7Drrd46zLRxNJgCHH9pg7cRPzcjTrvpYWIFUvagcFiHGPvs+9a
z1KwF5KwSdK6FzmMV5i7mq09P1yup3etZwJqbGKMsgOVO5NAC9l4mcTyyC0y262H
nmH92GWukxRWtC/nc7tDMaPyKChfHlDSa/3/9u+GxuC9+uTdWQA49vWb1uSD0+LS
0VEOfR+9OaTv2QqPOi6Zs2v10iD0VJngY4/P3KKkV1d9iroQVZ5Q8XJKivPrTvkG
xZUh6q3zNDcaY1gVnC8RdWFBmQSjMnAJU2xtn6ZHCKvL7z/Gl2CuMF5/aT79jfgQ
RSatBNLBfoJgA/LLLhYwbe/3JrSQao7mYxT07D3LxHd9/eCgRCLdTvrzPYB+nbX6
XvFJ32pp2VLXZXbdNW2b2qNoCX9XWgJKIbKIfHz3pxH4DzOnLoAXaQJbll25t/hG
8IIn9t56jD4GwTA8tSUQYQ+OqMAASWIFj1pNShHxouxtQYq1wZ/3rP/NsWQROGeb
o38VGin2aSdy1msa9BQj1GQTbn6llPOTu7/rDst9Obj7ZN6elWELI9OsL/ZAXUpf
1Ls8VGxcOigdCUQJnIUIvCfmphZru+WgGdBouuhG8z8UBsa36YGk0Pow2Fd/jJSp
WfajIPjIJysCcUrGeSDucsJ2RzcLbJgm3K2KUsA+tqKhAk46Vo7UW+WM8D+MW3Rh
IUa1iB88bwNFhVBq8LlrUzSNpvLFRv4oSoiD/S//EgJBQA2PW0XUsFTzX04+tQs4
fIaQjm21EoOc01t1a28YE5nMktOzez2wia2+HLR+uRDJW6o9Hap33A50P59vuTti
w/IEIijb89UUIJ7v+4OqnuxFjwqIiSLW5/SUqnxvxcj2zrapGNkZbIpXMVBrb8SY
EqIN1iLyW6IA2x5p6TMUOMMN/Y7Gc9JwVbYhMrHLhciV9qtC5CaHZQKn2d+Wnmq5
Ka6orSfGubmpGmyOWalPaJWjGoFK1PJVf3KKcFAFrPSv7FENwFfmRmDRexnm052e
nczFKzwm6Tb4YCBt7qwR5Phjm8NlBRAZJdyDOL8J3+n/AKRbziyuys0hKRowgDzy
hvbPmpUT1G3+Pp6/SS1k7qez6XZ7/Q/4HYAuoRzNDnt60Hm63HHUaKKk8qh5c81h
dZARhJjXcmYEb9ovl/fEPdZpL7X9/CiB1RfMVjZuBoWUyo5H5Yve997g4BKXkpjN
1vtxtILPYyzLyShaVSWjxjbc1cizv0kpu5mV5VUam5mLTBVpCg5n3Heh7DgGRXfS
cHUZYo2HRaZ1MK0mktUhXJp5IytDVvu72//DRO6PFK6tVlEtVtI7M7ue00SHHnyk
mqfPy7s7wnc4jaIlEssPOXNy0nsQAaU8ANQRdyhbrjqjut6JkntQ3iT4umTpvb0L
lB/5PfifhDqdjTN19N0OIbVLa4QTwi3trlemqRPComwaskaxWYm1Ai7VWu0NVjUq
+uGfl7N/01EU62EEhRgAcipI5g95wVv+mHkYCoDFsdpVo878CjX/8yMnIfvI3QOf
TgNf0mD/SQTsFxGGKOqAxc/D6YpRG/ihlOe18jFH2pljvKitTHOFDKTf61K5nYv7
4M27W9DppzeafkgynCERorzVgPX7vHI7OXdiBoc1KIdVwRWBE9RQnL/7OaBGCVAG
Y9m9eRYgD1JzU+PC3I1u5cUCr2oHXEIB3p0+AKQGsrhywLyygKiWExGEcZu1WUcv
C7RGXBufXOYZLdPSoHE5cb1qUVnWLRznR1wj9gcvbEAUH7U2/4gBWTBEGP7yFoe7
FD8BQSx7VVLtlw79gMAg5Ae6f4BTF1j52Xy0IF/7jCUj/MZZcrF9onNXgIQQC5lv
xAE3Zk7o62halegB/0HuMKgbxow4syJ8rBGMezLkt2+HGw/nYH1Uv1XuWjT3KSH4
UoIRaNLuWYt4SYp/+clOtlpQ+6k68r4FIie5l6WWI/XfXFITtIxYtd7m9qn2Uuk0
VzZM5oojSKsb71lngdgtSKj06W97t6CMI1pzuvsvVOi9tRa/7wvqKJHBIKrFvB/0
++9xBh1UZFZ6cJIt7sTG17wo3D/loia4bgKqLQTbZ7yHI0uCPZQ1zb8frXEWnJEl
doQRtbicn3ieAIC2sw+7zaKBL25NVTnwmt1IG2zhUo3ze22ZqwY/VCapgte22Wpo
F35MMFlwwqMdJphNmZkgieEDB2MmAVRgcYQ+wlrUSkISbiUx72+JiLKyqBqG8IBO
aL4JMKyhoU2YoqWUHKTBeh2y+W7A2JIIaEkK7tXoUKXWWY/Iz3gjLVuuROySj8dQ
BU+jM5qJWCS//C6bPZp6hmNLXYkWDoB7RzEvqsqNSc/nwgCJXD6TrQ76SUROkjwD
CuVIevMC8jqzbKogJerj1s2VvFbD0hJKE3u3lk/HCgSlpVziU2SaWxGCeKI88tcm
FQr+NWVIRkTjfcfe2Y4MLJddbSQQxTIwrD2R6z/CHo0Wn6MRhTo/SwF8/nEKHpx+
rRVcMoHsk+GQvX3BDpxsoFHPqK7f21UjMNsSJOZ3KoRqy1zhyyMmNNs8pajVxsI0
HuTEq30n2a37ahQvq2Ngxiaw+57NygDCK5eij1eBlFBmdy6BlULvqmhcfvVLJPGw
fXV9WIZstpIHK8Sgiwve2L/tbanTAE4Er4Jxg5M09OqLwvXQ/fz8PzAs4HGzxewB
fdGMqOSDR9v5DAsnP/ZNTMTTq4/JLk4s3pU3zmz85ttQYW3stJ0DCX4BH1GwMiWq
NedVh74OjsPZoRJtxwaHUi5eTpy/cjQyKRhDGuGZRlbQioDsOys00Qwx6YKkYwd6
KesRMdwjWRKToxmb6gWw5B3phtfLg5chdL5TF1AQt2ctIcaBV00LKDL5ENGDq4dR
TXzAGhncXJgRiW6y/jgcZned69cd2HVClrjBRYA1j4SALyKh6fAsuaytGeP7BQqs
fc/9hR1CPE8C8DPsHbXgYtceUZUGtbOlY1KPIlVUMLXHkTTck7JBmeuePrp3QhEp
3Y/pO7qPw8yo4sCcG2ZANWnpQ/V+uWQO6UiGEQjayUO20ZwF8RTkxqIFBbfHVcC4
kQDwx31eSbG1BQnXq0t62DKkmrsa9Xkr0Pcm8IXT26GJUc3RcP8XK5vNO3uiNNJl
i4tvP4cu+T98Mm+cl3/MEScBnj0mkcyKMmT6X7Rz3TLJPsuTuEnXaeL9H5z+Y0WC
WyGTzcGsShNfxMXJoSvx7Vm/erqqtmMWrt7q4btZHCenYM1VUJRJZ4+IEJVc0ysI
f8BXADPfCIcKzu1lxyFBIqu9MeCjdHY0FN+2YtfEiPTDYkY9xJM38gLKynK8qGgi
vhpNHgLBPaOH4rv+d6Xf3SLKO0JoLlqJwrWo5lwfexWSbKMddAnEQptkFCWrNmI5
bOkeihbp571qUS0zhyae3pdO6NSwMD1z5rNlkkpxdT9V5oAwaBtBsdQzgbL+W2JJ
UOj7u3+YoJ/ubILCt61kz7bTGrCaNnGUrh3Lrs2Rmkx/MvzLn3OpamxOiNl3jgzv
OVo6BU+ctdToIBVSUZB8qlcBT7ptdLRqJJ2fljgCYF4gZU/Vqcsrg4J2TDBq7qWy
S1k+SMZAXuNTgygtBkhPVTCL8LW7Z/ELfFIyZ+0UkcID4pMgPV8KQFTI+6JcB8Xa
GkrFDskoQl8WIyaCIaX3fVNWCqIjC17xeRVC+PfqC96Q9f9qD0PX3N4Necb9eFFT
b1rYmAQcDlJvUqPv0pPMr06k2ZWIAmWHcab7EMODpXUkolGwkXf8n6xhY4tUU/us
v0aXnnwqJ/2/ISX+s9EeHNKKoZtXJ60jXBEBDZY5KLEuAFXxkrktB5deCOuWAk8I
/9fpy2u+j87CaiRNA4SRHAbpXH8qQxXSWkr2pup7FfQn5BVwgYAq3NRbSSZ2YNKJ
pj2B/6vjHM4R0Rahf8tmgXa9p30zSwHd0bY1LyEJeDIWR/41Ypm6QF3nJfpM+0u7
Mdi/+bzGEK98RUkttIsL8qMv9ECzd+v+KK6H78DAv4q/4Iuwn5Uj0BfM8skr1QDd
kliBNeGb3sAB09CWP6wzmFLisZhe9Q45X+z/idt5LhzlyeGIGukXJHlAnVgf7vAE
25O+W8qmoJp/HLAmCmMiiIjQJV+R95TxdzbPFfVEqQoQOxOh+qP23BY0A+nruh/R
vMgr9S1ELZvGMAt71r3Ri1Lj2P1ZB7/Z8txH2g8G+xZaWNo/s4EiApXhEk687LhT
mAvy0W9SaXMJuuITN2vktGHBHGhhps1ikD+/JpaKG1epxszXSIUB0wpl+0GyhCLP
EeOeE9nzg6j3WfaII8loU8w1zGunglXQb1H1IhG3pcs1nysUl140Js8lt9vGsuM/
Idd++UyGQKdzI1Y6XWWw2hoHrI7nK1jE9LAvNGBLSwjvs8DX8DsikBAXtUJmH3a9
MWos8aYjlfMJ9CsoWgDbQEypHXMpLRb3ouwV1UzS1EJds9SiprFmuQiknZB1bBiz
xiLN5L68Da6r1N+WgPPQKNX9S3dpnoxKhMiowzoTAuJ6ixtCBxgB5PUkJrBNnmLf
ieo8Oc1HRfmoVTo/eUEzh0mWTt30I3YPh/MdmGLIUT7lHSpw57mvBfE8N7Aqv1Ky
Jcaw5pNer5nzyMvP1fqt9lxRstcPLCExpbitd9h084fiisPt1QPfSkwJitQnNHkW
uZoInhfg1j0z5nbNEksb8+ufBVgoauLtzvZAI5OrxJbVt9uGE/C7YQYDr2bTgb/8
vtiFZkWZwZfXHHHioZzKeDyrQpot/VWp5Tefn6nHRvHTp43qB2Scs9/vl+wzpA4y
M2JlwjBf0FBbLTq07zaVVFWL598xnkK7iJdy2Dhi9f+mXA+6lvsgGFttH+fA6pLg
xc/SAKDMsTP+K1yNyNhbdQnMi6krhyjLUlXgrTkKcaR4RkHpnAFR27QzA8ZofVGQ
xsgFMkMXxN73zsBEwdugM5xzIrlKb+ZOJfkKQ39mIwe5VtC957MJNDTVtS6XbJcR
KhbHoMxylcV19Lq65MRr4uPlyUsL9/gwrjV7s9Nw25YtOWaNpWZTjmFnkqj48VJg
NPx/uisoqtzTrnX5QNK6PDYlfqBGuKXtInxp55yy7bm0n2IZ5STeN7+74v3FloHE
B+EWNOksPQfzPeMDT0EjFp3yjWSaB2xdk+KLmO2Q61tVuWiE3kHNFwuEgPhPIBjZ
jxGfCs2HqcOg4dowI4O4CUTorKhvwbUhJ0dpDQxr2BV5wQUQ5kxbZyvDjVzDFkZH
BIpuH2RG+4J09b1B2R/zupAnfPTkny+4Ifg/6JsA/0LbNMN+2xhGpynbYbJZrF8G
VUgbRLrB78LLuGUvFlwNQa7OQMkrUXvnkpwYlia5iGTcnPgl0tgjmlBF7j+/1/7S
TfQ91sEzI7+Bc3KYkx8+oTV9S9PVMlNBy7xZFddsfq+iY0IHrDFEaNEo682uSW4D
LKUAs9tqATqHKe5fa5eUGm9nGhSoKFdl8gkIEAstvhtNyP0gaok9xQrCFiDcOZEi
h8s5hN6gUxDbA9APbaHTYn3hCzLN1jGPKrf8DY9ZbMAyLQtILI5t9fU8AOJlhKmx
tvtsJl8xVZHNX+Vdq2v9lSYzJ2hvyooQnFOs49aBjDXGNmxHiaQ9OblgIcZxHmcn
NopVKPhbJaiWpRUhOsRkjZIw6l/T3RCk23mawCoFzYmlINpyfpHcjpMLJ+lRQBHb
MKzvfQjsr3Uv01eX9DTwxGQtyB5SuIYhLIAMwQZ/ocQLRxXGVDjf/sHMZkPqytPM
BUpD8WFWCfz+qH5gpSlRXO7xFzwIpt//p/q0Bb+fxhnYod4wDo9nrNZGas5nLFpD
pXrWtZVmLjax5jwV/DNsNIQQF5RLvaIoIWiNjYOXqo1ppaBu3VTt3zl0j+l0u2Wk
hxzoumwgslST90C9bGGySmi4qoS8XS5/JA3AKPfiMdRc4csd7Q8TFopdQtgx5kjP
5l+Ns51SpBp3n5T22BxQylkJIBaT6wZ2l7tOVFflWEeQOEF4xsE8bA/TrpLRpEzU
Srntq5gtYBj06h93t4yWQEE6/zAaTa5SkI7GG22rmnammq0GNa3nv1iZKA+k39so
VI0tFrU4idJswd/xcv4nsUU101SCHj6wxHmHBtypiPsspOE3SAggyXgSrVgGepaR
0MwFXTXZYzZGkbi2q3eyHQlQJfJX03S5jeG+vumutsTTS1C5lV+Kb0f3fjtYKjCR
TtCfRqiR8xQlTYy1TRe43z93Ez0mnKbNYXN08LQ0cZWmdIOtu4biOdmE8AbDJM9n
TEtPMFKihjYx3bP7r7I4MpjQyvTBZ/Rz9lIu4P11DHvGJtpvKprDNqY2KOKMDzE/
Do9XNZfTFoKxSqVoXbAyc1VwSg1eLIN2LgptRIPKJutIR20U3/yc+DTiXoXD5Drc
NXA/SjJogs/D+5bKbLdD2qcuheHkxwM7NFRIbTPJmC8yPH6kuGfsRYNknrI7jWLa
Ah/vacOwbDBpPQp2UpC2I8sV3jiqYoj0UuQBjYuOP7cruWwGOcfWzle82hYGvKKu
F3zP3a79NeeSO0rH+NRzZCpI2w0L6D2Ze/kjecaDaoqB8uKCtVHd2P4EGC4yKtZU
O/GfV0dOkFxa3Md3y8148o6NV2lNtkucjY0C42sT+dy+cvFKc9VR1oV7GYJnQ1Vn
JxUsQhJIQuLq7E+qPXgJQgyX0cVtwrWnQI4i1mKiFzM3rvV3yqD5Q8NRazrxoARd
JZiGsxNIa2qbrhKoyias6PHyeEf0/VKE/sWr9TXDwUune7xxql8QRLPdnUz0nA0P
8nan7XcjuAVwVHbwNUf5hY6IHcnF2+geLG7RyB7bM0e8yPxDHI2XR9LIuWaTrC/O
pnlX1zCOKVFORcRI0x8zv5luVuXTR+jxtx+I9dcsPxZMolsojGvhKL6rf0pfDeUN
29Hs8M2jIWjQYctKDQWBcNbm/MANM/nPhSS3BBhR0mWeD8LrYK6pmLdV4V3KQQY1
pQVrqzH2OsjZ6y+v/UTGrTxikw10dlrRmr7vQLnU/reeX8SBhI16AD2BR/EV3pEt
C7Gm48OKc9vrysrJEg1e417eAy0sNUoEV5y7fYc9KunH2BJGhmstrGR0iTCI0VvN
o3S2373QlwkQYPvMbYNIM9JiGJ7JxoRz7NyHjxt1iMFAVUTThVp16rpkVx/K4R4c
wkSKnWFDV9FaaYqKnAiaZ9BxWO/o3P4bHsIlDWuit+/+igEy3N8eejwToUWA6D/8
tJum8dt4YW1X4deW3y0JPYEKb3FnFEt1puQx3nS9wss3hA139VktcGPFSp2eOzPN
Lmenp+6tyMsjxXyXcKrdPCdIqsp3K4D0DB/qVujLbP7HHQODRsc5opaFDjcBnckW
dw+zrDqWIiV4C70dqwzwknEEAaC8Z1A29HWHHF4/BTMw12nuB+MluE6ReTjQq9V8
+q1+upVKHKE6o/t38IYdsQfuphB8Ywi7DcsgO44jZhChYDzovLJ4tL2Lz9XrHxo6
dHI+3V5jumBnQ8mdcerDH2yNFNZl6tRklL9n8e/UOFRGnGD5acZiBnZ/FGAmTNJg
RPrmyncTj+oZXcOKue5UCAF2kBqO6b6eEdW6WDsgCx54iM4L/4OJBWG+LYN8XFX5
akFoUaXMpHmrKHjMJBgIWG93lR7/NIAf4+6MQgoWhl3J96O+OTnKEp3/vKytgxyA
39sHQqzNPJuYC5mGqZJQTzEILp3rIdsCWR9d2qXJ0dF9tpk0db5FCt0fo8L89c/d
S2rSXycv/VLK96AD4/V1q9rcn7wTfnlzQZS25SQhzyfh/a6jw0qTCoRNVmCA+6ax
jSPwgtWGvA9aH0WOVdmWYHzkwGzeEBiA1+H3uKewRNFaNFAwu5MKXTyk+7t0yid1
6M1N/8hQnD3g3U/NtMABCWm1vE+c0rwYEZONFtHI3GsI/LkUWVjZ6xb8rlcirCdV
vHabqGqCZjqZfwhJZGyBaMvH7DArf+qul/m67pIiOqCQbmjT+0C6unZwlWeMz8aE
m4hyVNEPiGuhMeIU6idk1wPb3r2SDBuAW9UjHvgMc9zUnbBf7tGHWCpvpY9wOcE5
Q30US0rNNlLRmouQTbsWOG19vkpyFLTyeCzxSmRmmGOrED/mNhHklgBjPl33n2Rf
MLpzAMu3Bs0WY+oDaR91lAdXifRb1fLc7sDylP8ArVA0fc2soF4CCxoOItfNA87k
x04VHu+fJBofd8eomc351wrkEFoj+cCC6UMINuUvpRpnuE9Mo2Qg57G0auPlTyV7
Bt5V3kQAWSOAxWtev9X+Ii8ygquiAOGDOv6oyu3PWFdrCNsbj9zdlDiMcOVHVeS+
hTpyesd6aA1fFdERMo9hmkN+BCJN3xQU6cSJTwkNiSU8Q8cKqyu/I6D4cfUYkWbQ
gRlVlvhNms+2Jw3DMxs6srzgA9g+rEveKqECegdzsNj1stE0AzwXV+v8eEeZgQ7c
l47n4Pn+aPYOyBgXv0WysM04x7t50jWjOR3jsTGtLly4f9FhDXqk8L/k06qOvXQQ
zkrsQwwgLb2SyEp33KyawcIOJsnzCzPbv+ep7jWoL++Yv1+ToeQqL/2ajmma1w/P
YYHJwGGVAwm+jZY3TYrNaWylFhKPiePubT1MWp58T9oi+rZO7UKVr2J8wN1L69nE
pjT0Ym4csCB9J4PZ6NwOzfn3UqM2ZSM6pAnC7kmIBHasflvlhYZjONg6gdIGLD58
Z30lh9shSFzYzm/7Uj7V7xyMJORfJlQxlTS1py/fdxGh/d9WH8+2zUelkkV40FVU
0rNwU4eXG81UKeCh85eEPaf6tpEblIFJA97xow3+iMdilp2FJLH+S2dxXp+8AUsw
3F20fI8V17uLXdxAPV0WXcbt18r3OAt+pyVjZTuekJgWGtBLV1L0p15a5G5rPwMo
Ovo+emCunr3daKsrZdPRDI6lto2Hrhx9TZGtg4dfu/QfkKjQfpwnGZewClFvqaSq
64lFZ7jQEM4sdp3NsFMwZxfayvEezfBNfWOGRdCFoucDBeeFqGSNjp0hon3oKsti
2CTFOmKSqvSlM6bwosvswFdhNT2dK2ZzBuMta20Z335P5s94Kmmc/BriL3NZpSNq
xTFl54qhEreFyJ+aZeDGGg2QvnngOXwvopZzTsdujVZa+uLe65PJimQDQZHCwxdg
oYn2hnnVXlopn+uEAErnFVMUPFaUi9vJ0Lmsq+Xczv7RQ5kvJGLkssyexr+vceU3
GLOhQj6NQcmVqnVdLWesaOBeiAH1Yw+ydaMdR7p3bgyFb4OpN131jDduookJOGeL
vFJHSN30SpOYV90T++ZBGSpsO+5CbBU+B2PvivaUXl3c0W7UV6icBPaQdLAwznMw
b0N9eu8LUkI7VwyJ7xPpTKyj8jm/E2zAm5oFYPMG0n9ytMOVZrZOJdiy3IsIh2oU
+zssrlJDdTfsnb8O6H5hLuxis98bYTe6ubztN2ENb7c8Ma6ZPtcyiJRpnD/4o/Lf
Qfqwo24Lvg8BiKPZeSV1658I8l7KtettYnlOukSGBJe29InswSkN2zBucWTbdbRr
xJAmboxSRYFYJPC62uAXnDW2FU5UdIaQ9WaynIZ0y0TWr20QWzUI1EikACWd6yko
u6i9GDUhdjrbWHIOBKTWtl13I/zZS7WpsgWuXvMaTHHeuoBdsbGcQRqBuGabZvUh
ao+9X4YPFWkk9he971SiRLlZaDEGJ75DRZ08ZQndCUCTj8wLXnnIXqGz3cF+FUJM
wAqJlpG+7ISIjQ8o4+2WhPi0TIlNggms/wZGliv7Vdt12hzdZZrO07b4qm4cvlMH
VV8mh2H5s2Fl45UyqqVf0CgRnB5QMIFojlDs9mbGpwjPKP1+1aFVfErAAPWz1kRz
5uRtU2rJ1V2idMo7CX8P93JdablmTiJ5Jlv1bU3IkKOqkdeRV4CeuptsUNQpW93m
EogkIlhbFX0HBEYTCgzG169mWIl2rkZ7klZSiJ2VD8rBKUFdg5igR5VEEs9HGU2A
YRznpFNt7kA5ObbhYnEb5DtHwyAJPGfndXJqJaxLui1rv2pnjFcfBPn3/gOCAG5a
/s3cHpAVB+EVfaHTb8Sq7xk/9rtrRShzW9ak5DLBVfziVVvSU2+1s5YaWi27GZYX
YIwEszQXPOjG4m/f0mSMTGsxNXqTz0MxDizK/v4UPMjjloNDZ3Qd8aXIXnJsd9Uh
T/6k5uSQbIQv3c9HOOWHbudyu4PbKiWoJuwemIVakn4fMUax1f8QIH9ZfrSgutcQ
ugpWs2AWwSlSOPvv69aWBjOc8CJveLjJXb7B5POI3xG0j+Wfy4yWAQVctwpb/pnk
E1Z0xTgxid4WlM9lXkMKEG+gq1du/5sOygJxOWIaqDynqMGlGTzyFa9EAnzoZ6cF
e2+XFPIKEy7iOQ000ODRq/6pQvIVP1Sa4ipu1WlNDm+seJYxJ5s+77DvbDxh+dDT
u9urJRkSek6tMIAht11M6ka+doMEZdtisffesiseeQ09jclD1hA2w7H0j3QCJDpG
17bOKWJlSCV915nLahyfe+p0R6URPRcV2qSnYsDcw7CYIDx1Z+iGROUyJjeU95HL
LL8ZFHdgZZ3fKTIpc9o6+dwSxNxKqC+Vue/1R5S4GpbSu3wy4jE/jGUwITm+pak2
UdstsLBRzM71x4T+thRPEna+Uj3f5hhGNNCrDVlboDJTQcsaRqVBE2YmrrCjGCNQ
WZHeXhaZG4SgpYqcwzGorsL2jve3hZ9W3UkZjbBh3BAAVvvuBWnpi/zs1BMwT4nS
e7TKk2yr/BhNIFP/ebEvw2uv2cALP9uWCO+JTVKwU69slAVfggC20Y8uSdaLKWLs
Lx+Kje161aCZvAy3yhdn33D0XR+gv8PRVu/qKA3TJ7c/UvO2mnCyhpFofGdNIe3D
T3/gcnDxWNWI61B5OR0Myv0JILX3JLyrj1YS+2yJ5q+KLz2CcWVgXS8fY/6/m/46
skb4+IVjEccooDTmj+SLSurZg8Av8EYDGdd1AdnzcQyw7sfeFqMnuyzR6i6mexir
JfAs6rxCTfQx5UhloTj/LtLsDJM4dqnJQ0i6PBRLL/rVrA+AGWDCC6psSCKf+/Rg
1tapHNMIU92ybOWL4vqxOzmJLXflvjawU6//UC8bIJ2baQZz028WuHRRJTPRcmGd
W3/+v67bn6pZEhh4E8Zyl27dPUvt0twYc87Nnqzw10uw7QfW2R786zvQXsMJLChk
0I+8RCT85CRpCeK2ClunIPYD1PK5Q+VUvMXKTpu/8pErdaLh4JGrTdrL+GZPa+K7
YvfMJz84VFV45OJsq4D0sJq/yYwS7BBn+mKB7eLidNDAB91Ob8LWmKsUR8hWLN08
i5BdeuGQNevbSTWhq4VDX2MCmntXmb4LHTqBs8osz1hciapDVBg7al9IyqmROW9z
hCoT45R+TA+PMR9uliF4NYISaHxZ0U6/c0gYkzMYaK3vGciqseJ2LvHRfuAOzHsX
HzfoxI7Weo3QdZuQzGQujbxK3bmmXlok/c9O/pS6Ee0iTNG3Kmn86NE+BihSj2zu
fxGvZtZuJ3UZIVQz1Ep4nYJhIIMlILCp3E8J2CyKM+q85V5ntMi8hJOWqAKixANM
N2rSNHfNpenUjoGJGzf1Pd5BAkRP5kCcvaDLk00dFVqkLnTQEDTdqbve1DZKqN+g
/89EBv6BAFoimhAaD067R9oPpP8X9bJX/t3B0Fz7iEk658UjmO+5I9Godg8qJNL7
dXsNHnkYog4kDOnl9yxS0ml3YdJt3lNrHtVmVyLzl7c6eloqBz2k6J1IMzTbQbls
PMjrMjhVOeqN8AozG/IDEbLfo/+Awuw0wrb20FyrfrN8Qw3ZV2mOn1ZZ+qUagj8B
SjT/cRrA+1fFswM8YsAjgekF19knwu2r5MPQTS+x2tH3rSNiM+WU22n9Xbwfq2X1
39UqMsNwzCste+Vs507piK0qDxaoWWHqu0UDT8fqeiEhed5ivC5ZXsnA06ZxwiyV
asGcdX1lJEUEYQ/O3mXrqDTeV9+rzmO9XYEcis9MCV8llYx36mRSAuT8LVZkDexm
FV+wQGGe1826mjadfF4wspr4G8PHWgNNvlrfORA+VOnYunNBK6m9L0BKiQkoMqAE
etI946JtCgLalVL89fuQz8K3cxxESV/ZIpTKJ8w7MKMQvouLovx8iJQYt3T93i87
/pccgCl7VVZcmlQ9DisQPzfJ+dMFQ/1j0r+gyrGNUzQB1FeGBcEqRi86WNtHFxt+
xKXHtvt06biSkRSFTCkgrP/eODV6yvKord4Ak3iRr0x2DkkFr2xl+h6/CbGCKlFP
WkEqHxUgXMEY4J0HRVIuIDFgELThiDAqgME6WXImcSi9mXQd5zZcmSjDaxOrZ5UM
Uk57+Xd+hV+VTMdFDnnsKZhaELNw50ZKNLBMOoY2q/ibkJ3NkJ7htgynqjFDZ6m3
IBrG4LeCsMqcyxSiSLY49jNJAWAiKty0M3FoRYaLktziwSTMk1vkrYvic34MvxgF
WxMUqVGEbfFQwBtVjIQgXn9uS1cgzlmXYBDq9yh55aN0pwN3xBHISVgMe4Frop6R
KEYM3xey99WHopeUd1mcm3jbmB1vCluYwNKEpG/YISxjNFcl+dfhYp8P3jchnzDX
kp8LBifKeJufBGubRDOfy6n3DAuDH2XXHnOp20vI0zF8AZRUioGX2wTXTiev7Bya
ac6JwlB3cwRcyXGC3iZzQBagbpa8afEw2yWWSaKnU9T2BwuykN7q509TJXYmyFMG
fmVOn7GVnaIGvj/f0jlaRbrR0EeTJ9yoaBJhJImEsCnP1q6HkRRQ9rYcT2FHy755
uLNZxQ09hh7HRxrDI0qUn0KNWNifzh+1kIoCaVjJsHyJNDmLVNqHAOSmmsMD+JGr
tBzPR3QDA6OsyxacoB2gCvtXAyNoR7iTSEPhZu8waXWEODvIeWyDa4LW5F+FZAIu
AwmQ6/r9R8kqidUOplQo8FS6pwSfwQlaaCpH5MWJEkRN4ncH5FhKKkrVr37XmzYn
FckLw99Q5m04280SXf5M+Ehs8PXnhvG305wpSKy9Ha5C9b8FImzGltSpHsqUHXMx
oAOAVdzUcLjttlgg3J1kxK1U78I5j2gevmLncBO+/JwWNSXkjbsxvr7UwPvyZN+c
dde4GeLh9L3K3eUOiIXqObsQv4ujqsyDibNoZ5H129L00O+Mx9kGR6IJqNhea7nY
l1hIJF0934jt85zydHaA4+7qNrqF+tIxoYRm/M6hP/4sFSoFuI+v7GgKaKwTjDd2
Uce0kTqQqvE23kuXJWRd5MJPpcR/gWAU8jRtzdpmvDp5iDH3R2MLliYRq8jif1Gm
J2EN2EuAgr3x6/eipyWFoUvlQWzu24H4abJHglEEQuTXYOFhFR9MhSUAI+G76kHn
x1RW8QJY8ndAmEiJj3zEL/1KSyLSeZvjIrk6f/CL0zIbX9DplVkJvlgTnDErEbkb
kF1Hdu8quA6feImwP2HcvJKFXrk3vc1V/3i76cgSFvl5mRHgpR7EzJ6/8BTYp8MS
WbePkbHqBFq7fAUnV9gBqGY+fp9lfrETdSe+8MY1TUfOo0aI+jDoKLhWoy3oPiX4
j9/cbPt74RgVrsGrGPKkVJX0tmuf0/5QudBF+q8+8bSCLybpkPkwk+Vl9VPSwvo7
aFz4J+CTxoNq1VgQ58PsdFXsZQEpKd8a/kZUCAsQv4oh4M+jEDLgCnZdZaAaACw1
wjUvtQ4fN8jwOTYZ1DQI4Rx4tXQocdou6tyhOGX+31ItlAA5zR2+ENkN6ifalA1+
8DVzLXWxUamSl+G8BBTZIyQD1gmcWfCiGIokuB4XaC7HaJsLfErvhGwv+juIWC9i
kC8jZi5jXi/udmpFgEzfnxrSHTs6jiXR3DV8e6EkY3bzr69/PjwPsrL1EaeqaH8C
BBGAWNF36cQmcbKxNi/Etq6N+pyZyp/uFk1RfJHuA2E5IbGrY0SeRujEus2dapqZ
7svAUxkBVB4KZzbCeQu/AXLFAQn6JoWC0shc5ARwWjWlVmGnzC4c3fNt1nguxiMO
cuqoNtD+dpRkHCazS698GFyDYquAVk3B4G6MH5BM+5sd6HicDEQJgN3ukBahX7qt
+BhavQ5zgLlTDqmpfmS5aZm1OrGlHrPd229AjARbhru52KOYzTUvthavtw2PmjpV
3unjzA1ZPilA+duO3Pd0cgsGSFbOGmKcj0ps4TU488jaAkjwKn4uKHbvkap7dNVO
j4ptlIrP8JsjYHsyVWWiSeIXOw9y//l5w5uEZ/yFrEBw0KHd4zZK+Nv/VksiLGvh
C/5/tXvjLUYVYJuazs/Dva9JA/3Rhcxz2nMAMr2RVIqXl6tS7xuPn4WzjarNs8+k
E9wmLzD06esh269TlTQmdyvoiswiPL7DSZDt3i64S+0HUCOcLQyht8mB/lyAbFK6
0dkzuSvB7A9K71SwXsRaqGQ8v+4zd6Di5hnu1/nyjcImiHJbBbcgQHxNQ6G6J2NB
aUfekvUPlJr2VdvXqmwxb13aSgdFMe8gnqI5o+nwoP/q8LojKIMQbcu0whY6LWP8
yWHZvJxRok7bu79KvUFSuwxm0q/dmGnpxdurectq0pd/Kc7UJY3mMho0f50Glnnw
2i4ZRjuw1JWxLPuiF6DTqqICZbyuV7J5qGoo1/7Ax2FiVnasRuia44ZFkfBBH4fM
u44yHfy0i/LRbk3ZDFiRQZAXHJI4AnfaQN/c6Mz6SOrPEJz112SFOYDVZ0ljaYfL
TL1OCwe/92WC5FCp2pY1WiwxusoO57HKQk4SqqKHFQVx/fTNGlMehpI8qTK04nR4
zBFmx6L8LxXeOD7CNQzBr6aYkyV9OF4ek5FVrNJmRKyupGgx0gRrZAziCIKU7nqR
8tLEXVUNrqzRRBb3KodqwO+CJN2JaCQz/rhUn6Kpe45lp3tMwB9Qm71fYcykB4J2
KhC36mzt3xKzVf5yncpPnPQuA/YlYUFv8YU2mankALLy7Cuhq0ZkARxkVyDNkbML
bLjmZP0yFcxe+z10xyFdHC1sc3MG1rID47Ej1ZRucIaRHkRHQPAL0YEAuOWsTXUS
D2ixfN4Nq1vneQgPLOqriwvv28rv+1sT77txNw6cGtzpa/HiksZoOCh7YiUMURfj
Clqs54qjXdCAysX+/d9LcFgRQMPgRHL3/5gEF8KJEGkppt0rfY7+3M/ryIczKNM/
jk2SaUVZVGBC/6BO6S/nJGNJixYRCPCpImdeSubz6AkvSCrvUWeSUQe1d00+mqR9
tS7avL8k0Q+sAvRkyzw7+BuojQa0Cigq1P26WOdD299l9g3beM316tq1dtkFJrGl
MYT8O/7wyVdeae7l9FBAcU/D0tPPTcqpGGtxpvpURME/s/xaxfR88DAH6ShiRe2o
cKfpQmUooNuuHvCfh9A/TUgXzRCvJSYlB8gHKPd1oLHD5/9SQKZtlrqj/gAKg8AR
W7R+oAdfIHvwCALyOVAM2Y/FUev0PvWHDFe3KKfY9eB03zYbFSY0hMP1vk4YLr/b
uJGDcd++e5WI6gH4mV+UZW+bsG50rC+f33BzA7+0vq/EiR4T7kfvtGDbEl0HZMgv
kOcPtSEcSvES14Zg0fBxnsYzV7mN79/tL69nFMDXwvge4TkJEa7x/nLXvFDMeBmD
cwa+haHdyNsFblAdIZLJeBuJrRGbZA+8uJCggEfAhFs3oPPRHS5/+/6GIgj1HWuT
Rib+Y1mGC4A0xyX2PzXgbmJI6Au1IKnYSuuM02VRHuPkXaqT+E/iBbt+PhqMnQhR
expx5/+JL8xMtz4kUjqel0k/IJPVS76zmklDD6dmM5Q9InHzxWJ+pIiPK/bFdZ4n
YQKuY991Qk8f0lLEqneSaeyb8Wp4IS7aGcoCXJbI4k6/LlOiBhLfaKeUH6vg1g48
ygMMTqdqe5c3j0IVilcFoPQJXFFCmPlRhKMEcarlT1/c5+pIzTqjWhWmCVaUGfJz
ThwhQ5jiBrLtX40zv4E8NLVqOlxYGfp6QFu5NpDuF8m0ihwdoN9v4xnlTlHi3gdH
DYtMdRG32WW/rs9m5CIFvO+FifcmbcoJXNvSn8uQbn2XEfuXMY8aMa8TkFU/onjf
lGhEvHtKRgutDSRsQQAuDIEIOXkTpOqP4EpeuoABGEjLa2+sZFSDXrsn8AZb2esk
xt3vx9C92MU1kYDz0scgSF7CCst0PpZKU9t13B3+T1g8JXHIGF7HF0ocHkI9iKd2
a4B5qP+SJnaxD932h7/wpV2GjNiyl6hkJaUDQrqB0C4Q58/FtAaaP/veRf//dG2M
iXKByNoekJzX/eemj959JsXEXJnqAbU3WAkyYUjW1RclrtRRWQbm3Homd8D1Uo07
/yCDK6Pm9zaHYNvC7XsqgMmQ/oId99I0935FcctoBN9R+p0sBqLzNJUfn0PLu2fF
S10FGFSZkLX7zR+TB2ZOZ3sC2931le3YIIzdeBMWbQmbbQOM9hBY9olqtM2Im6EY
HYOJLY1XrNhtFED0nirNIX3QgHuSggd5XHdXomlJO17kCLLzby+o3dw7DnAV/Gfz
3qI4c6mxdL7NsMQUhiYSumsdwtllcgrwCne/c8nQZYhT+zG6RWvMkXJMslSnUYB7
oE+X5b6mV/w2U6/lqdLZxqqqzuW4kSq9S3sGAFErKoYWP7y9vNJNg/Hi3SldL5kB
4MLWxdhd4I2LZByB3xXmzztnFUw22JFI7aI4v9sOoww6eo44GWCKs1GwRfIx8yiL
o+BHQqekNfzzfWQLJmGnTf7sOXdIQN6nEHJoW87oiIbK+kMNBw1uvXrqysKgVuRI
FD/L6ZHnhZD3nUMZlFLW2JhBeT1ljVaSrtm4ZzL/YcK1qsoTaY2gpje1EHffsZY8
ZgSd0S0U65mRrJlH3Wx0yj+6RIRHYBRVpgjenkGohAF+R6sm9Dl2HoxUpKrREFqg
RTRf9xQFX2d6kGahVy6E1jF/y7I67tkG4JmieTBHgYlOvJ3qC+PnLLkY0yY5iLTn
gFJMmi8TE/WWIk4y1lCnuvHi/E3RA6P69iDNXXVel/tp1mbH7xfV24dfl1djCrnC
Ub9BN/gGViTWkLDGbShGb6lcpMxptvkBZtPHLwuRIG0GmNlp9ASUb01v90YVEUZp
bmLNEVQmyIlBFK8nGdsh9DXPYm82/rw7mAxMNLjMES8MfO/BGQHNyGd2hHzUp/ks
QVdZMqA684PLy6syfnldeoSPM3/+Q7ycLtyI7eURMff9mGdcMDlYhVBmucUZkDcv
pY5FSd1ATZ/kAz7ka4W9Kgsvbf1L6PQPXUrtkJQiJLd8LEVLRHGI/NwfK/K3ussj
4I3hNpD5PxPGNL2pub9QUJ0M7fUGoGJ74TAZ6fEWnmrlmlf11JQwUWra53AUvzCQ
5pf9V8MFsfYpfkr/+x4QHkBWhskNb1PVaApg7dBR5JYISYJ1EMO7poFYzxGJv1dg
2qngUemLBrSS51r2F2fUXm3OWMTv2gxr/MRbi9ENFZYqIdJRGP3zhtz0O5U3kBB4
zaBKq+Yi95oPteflbh5OMVlNWsbLE+216geKyf+k3GQjkqHO9chQIycBRpGh/n0p
Ov0ffQ69B78jS4TwKpRnEqcQAGevw2omVa1UKDqSQ7bmCVTCpInwOu5aJeFtfaOO
63yAdckImoA+yjH10qyc7LIqguUyJkF6qlEdgXcebccNKOcrFQ+A90U3pw7bIb9d
p3ZK8OyThAcC9AgWkgBuyCS6A+HMbby83awn5BouK1Un6MY6/iaSgzdtfCg+msA4
H1lBxmk9QHERWRS4ZDjmyMxEJKHwhYbmzBGw9fD5qtAWX66NUybCWubuE/fKsi4c
t6DAl7mTieM7TSiJ5bs7jJdNwGqdvZsDrL1LTesFuPrP7FuVPPtCcYwJiqsOeW3+
1G/Tzsc24Xdk4Ls9Fv9FjTLSdEy5jpb5x2nmdTLRPHI+1QBretvqmgbuGBu6iJkx
hMa67q3KF3PEe7oLhU6ZyqqXNjHIKt5eILj1xImFHLngJaZHX1n/qOpKyHdyTurR
YAQ3/s4KltIVn3QHetZAUSzVlnp/jU+R67N1Dmzz02su1bkikcus2mH370bx8htu
UJ+HFRdo/zT793nWeHVTRKGQFL86HRRSnmTf8MQL+7yUzmZDbteUsjwqbXN46bFk
93jFYA3Y+0Dj9CPf2eMx32Z2c/1fPubFFN4Koqhl/p5IuvPDLIcXW4RERaYJuczd
8yqqoN/1xLLT9CHKjZsqtWc5+mglBrEhzGmGDjaYe8W1m/IN3KFxgb+RQ8Fsdr1h
kQKjlL8itG2e7lwMvjNJtnlJEDd54LZ2Gfd1HF5nvS+VzfVDKnFiJUT+R43W2pwC
cO5zkm6Ww/X0nqxJOpWN247A7OGCZe/8K2Xke6DH3jcISaevdCckFRCAScXa8+xa
6P6agY4dGHLFXxP9Wzr6agml1SYxHEffjifBenRmhORVSQKzRcmUcVUJk/XiGuE6
vKwuGqu9WVX9YARAEv8Ewo5bp1QZ9UzUTlxZyrS0GYE+HQWjXB8JcghfRaFArEsp
y47pYumeMx1k5SR+Fh6KFmEayzcNGIY+mZiYmJUvWZZSX6UbQSkQ9ANNr+nZvQcU
tsDBBrt3OZ/KaiQmO6A5SCieT+o8nW6XHu6sqpZufUNm0I0+hE3CJGcgyNm3uXDG
x4x8BQX2nSmM8qBNl2nxCfbfjyZ7xJ6DUEbioLg/kNIFMpYTuecBCowKf9Gz+jxV
juRfS4czz9rkbUy3Ej8jMPf7rBURKDbWsOIFphreGMLpdpJb3sP8KK3iMyxglIw0
kXb6cuZrNx9+8acYIPI1g3yRIu4FjRZkYcpw3dU7aUVSS2upkmtkxVym6PTjSVaV
98i0vx23KSOn/udIwqCii+dYZGSFWcsyr1YdsiSXON9UOIpIG5NlP/jtZ0lvmVLK
um65K1mxUMGyzWxY4FJlwOGIG7OJfWtx/SOOmUo4ZbqZd5Z61wfEloRKYHrttBss
m8gm29/kjwAr+tQvBYJywNzLPc02HuRj/j08rFUiK3No+BAlHtSvi8EEOwcwUACq
DvXT+7Qb5uMFnLBjeqwgze4sqjaue7rU32Q1U1bVaYVJcstNsRZlPot40tR6qgta
UNCS9UAQxMgGlDcbAO50StIvWa/YERajo8k1noWmuIYPD3X8LB2RknArycCNRqy/
S/Pb0ehHuybJtrDKBbg+WTXT9FGXs1ML05hfGAxiuqu/oNTl0JBG97TT35OxWDgk
cFdGBD+X6spU/M6JD3cveXPnLxfjXre8JujlAlbjfxT70VXyIxGduXpU8clAtrTw
W5DF5KQA+OhiO2AG5Rsv2iSb79Haq+C29jlhRg0OJeKtO/rDlLrOY8Njm/qRk3Do
YY/Mi8E/qFNlgb8iTCJp5JhEwwwgtheb7t3E4J6ScnjOx3FjZ5TRSYw+ZqUVoVVs
VJx7uE4mPnT4D/Ro+L9h+/I51yeTTFzewWnUM32ZBwyhp+RTjGKpJ0Iy4AwqxmOG
XBiRFKrYuJgaAeaIsOmDnBu/eliHPsaZyH3ifkjoYkuLiy175FS2xUcL3Gyb68U+
NvK9CBju+IaRo2hh+O7aJ6EqWtJU2Yxg1i6jKjYKv9eABTsstl9Uq0djCGd8Tx+S
KH7bcrh68RA50WYvU9BBnFpaXmbPGh9vzg6PuFrEYkNj7NRmx/G7hljZwJzNquSH
CXuOntKG/aoXQZY5r5+/wL3cLkCwztSm/7hQ0FQo5jCpHbVhfjOgx3H62/Nh18+7
MNHx03dl2Ti9tOyJIbFjvSsCKxkxqdcVKJmL82NOyUbhSgG56X3k9AKKbRwcCrEi
9SuVqIQaGJAUdmztq884YNF2a0SGw4OwmfBMQLM1Fjcq/mI2f2TqJp9dXlpJSgYd
IMIb2NFkbyq/7C0Dbesb9MzHqXWT3lb05GIP8I8zeNdh6aubOdMyoeW8HgbjMdz/
AbiCGouQdgqCgBec+9wR0hLNehJo+42PyhubcNiCCDxzD50q/KCeB0v+7ggiC1cg
ubtvHzcTvpsCIsH7NLM2/BmJmKQCYYnaGapZYfKsFGS6Q2GpcsYquAZ1TXplEGvI
K+xjl2bIGJoH93nd+FBrlav4nGjCRtT8gop4e7oivlZY8eAWKLdR+v3a2VqqJTa8
+OjD7Ge/ZZr35pN8EOgM85rMBMBPvYL8SBhHjeGH5WMg6cgXZmWYF6kbNs25s801
8/XfUpW5qWVMt/v5diy63i7J0KUeKdCt90q1RBEzX5AuHU1UMQ0Oigui2HXan3sg
s5ihd5V/dDEkcESB+qMK+gW+HLIbrW80cAIcz4RuaRGZ1ziICWmWKT8bzS6WPUbS
ancZ8Y3hMhRWxIknSeVeKfZqNcfSlqZJtOGk85Bbuw2JVKwOfHUabv/ZagwsIaXb
p9pXdF6x5s4nIMYwXlu3E0mHBkBEwhPOl8Cy4ccQuLwNmA7QT4xr8bdn0CbGzmG1
rjK0K+3FtMQGIFqvBXIq1Mqyk/mNOSv3Qj1Tr+oBVvPn2BWQ3ujEB4PqvU5ex8Xe
vL2oz+CgtTXPkaCJjVDRMScGDrq9rn7a6cpxixHOGHoSKLpmzLxoggjsf/0Xi+36
H6qkar4rh2pKvYfrTaYG6pglEgm1gkFK0ofcZyLCLKtrJhAFcB4BuDGMeylqtPYk
3/V14UweSwqrxDV3DRHS0whxCuQY69x/UTywrP4gLXEzrkSSah3i2Q2d6bL1GtWY
XRQQb5mIEOawq3ix0b8v0xT7QyvRu6c6JG4+LIiRK8mf6JxSabXdL4qTn3HWr7XN
lNgIN3Ae4520yBF0jMl193i2V2l2CebpViYY1bvrzsRUB7ampW93liO8vxU6zDdv
ZRemEr8CQWAJyZKScgoNU+/g61aFMKbt5B0SyBXWPMxMpzVJggo+UQBEnQeas7VR
b+jQCD4uyEKN7/p+5WOWBJnQNZSHgw/JrkxaQYPe4i7bpko5gPz2jt+LQM6n7gYy
PR+jd/JrtkIhDcitk+SWIo6JpEarTLpv27trl+vvHlf4ix/NZmmegYkRoppMJ+0e
JkrgHNPBqhekRhTjl2rcR7PYy7nwHBQ8lR+1zkHviT8hxno1U3xi375nUy92DVnm
veO/S/5mtmwgWaDy06AqV6mlrp07RFb3eE4ntk1lftI3OcpEuyfIhnU7ihU3ZycA
b/XGx9bSsGqvvRWJ5XYWgtXMAPQ7DWyyehpBw/ViPRbEsE0fEJPRwmUUXu237LdD
QaRqUMN2Fh4fkrKYG/r1Ys1kWk8p6aHraEwOVULvqROBhEksCeGbT0ixKhsVBT6Y
KRMPyleGFjKoAl9oX9V+HCi8BxbhSAi+4crfW65/j1Tq1a8/dHn8eYBlQK59CliH
x7GQpqCVa6t57QNnTZP66VzS/O7Ny0nzXu/lJS2c047xMwJjjDfJ9akySebp6X8C
XWwrkpOFPJkgY82P7JJC0kuLl8YpDmsw+1OoFcuXVgO4Ah4Zxl7KjSXNR/t995pQ
A4seLG7nF9PvnlByfxE+l7GErtkvtL/FVvwew1YOT/3PW9ic1YqKPRrZkB3jxpqG
LtwtY9LlAXd1wBolD2+cdsVbtodzFg9li2YXbvrMmLYdKwb0BRuX+P45yAYVoK35
2otKgBk9h1PsAOozhoHtLdpDd/P+AAolyGboMarSTRU8ygBRQn8icQ1l+SAmjnJ6
XVGz1occ4ilHTPhuC53V4vSe8G9dE79SGfAQ87d9I5NwBlYBb1DR/Q3IZYwl5Ya6
WFPHIZoRROnNS1kQg+u2GgkDrAWzsvNv0iuQ9ZdKnLvJ0LvfIQryNk+7c3cTuM8r
S84lNF9xArnY98xhpt/Wif3dRIV1OeGwUeJILMYUnAvcL5d/68LO+F2eWb7NezWh
fv4/wYvNz902+l/0jAOHunsoNp4zbLrto0PsH0jLSfcGM6zWaoHmZ1h7Wu5348wA
0CQje+pH5rQL5GxKHM/RlpWF8wnD3l4gqNTH6rGUL8f9PXl9n5ID2HB2jxkyjdpb
fIgXFZdLnKO/6Lz0RVKloHMuOkrtcAMlC6enZ+3piCJoA3TXN2jvkstpi9pY1r6y
Tknc3/tXfqMrWMRAO1mGvFin+1J5SrrcWMuzIDkzXPcaurdoIFCc0WnEVflljPbs
LwAXEa/JeM6dVUfm/an+auFu7cFhHaHGx4Cpjgw7dGBw/qm8xO0LsfrYTTAqInDF
OfvY9Ojvl4LRgoDqNV2WIat98rRZ1z4f1pGzyt0wTGrC3h+OjlaDz+wN9mfVLFrl
09lzXbA51wjNMlkRoudscYMPVZAdsWjO/QAKcUhtSoXGMsIRzh3Jzrmdu8btH9ML
7BUhiiqKRuWSWMR+KJ3c/MqZk1zynN/a2fk1Y/PXKHDedtjhc/BtWvx/wOaFU0yt
Rsr2gBqRtZdv47o0yd76R8jfvQ+D5N39QdUV6CpbQav7LhD4JkUNMpB3QRFPTRcJ
1OfYUlcqQA1QQqOKwiuJTXpSWkd4Ggv7B6KPRwEYnvYOS4fnrWPcqaot2B7JH7Y2
L6TT/CGWlqdFuXhKeuHyfq9KPCHUqZcLRsIFllvIPb+KHV3oQH5E3dOJV0WYM56K
yjqHHQzmcufDHBO4LxJ3VO1b63Zq63Q3zxbueH6HlK4y7Oc1CTtBCYFoj3D8gpZB
C1oUASVn4siewouSMyOgg1rq00WqB9hDDr4/QiPzxJmLAt5Eu1PbKkEvrGyeiHZQ
q3e4BfC1Ib3OUth3pkXsvW+a5UEe1qI6D8/+eIkzrsb0xodXm51fUoTYNQhUOzgo
HfHKzEGKhgfFzKdaUEdMsbxytbGJDrceLFFsoSDeQcnTHMQOA8SroMfj0cfC5Qls
VBhcPdM6/NNJw+x2CkRVh1BVuZndvTUJD//q/vjPdglzzWdLSDRwerW9eQZk5zMs
J08HGYPnjRAIaJnVXCTt+pG6g/YcgVU5NjPtsfWGIxM02e7BbfF2BGzZ6+kV92Yi
FDXt9jXn7kv8UA+D2PBxrypt6lBYN+2FalAWEKnxaJotIvTKjPhyjNr6S+aeHSxO
zW3rmh/AbAYpEDk6EkFpB+7FKcfRvjJ8YvfHSgojPU6a+CI+XhSxPD1wp0UXl2AC
ZHFZlCczhpD6JqBmIHXnj1ArHTqpDLER0XxRQicT2FWyguoBrIdCOHlAKUqpCl5Q
02BU/i0QKg/Qvk8hA5wWOcJ0gFmcrHqyfi2UY5PGnP52WKO6jlJ7Qv1lJwaY6Ndv
awITvMCb8JGpox5Mt2sEm4pUONHIKLdUtRHheQxu2cJewwyrAXislnlaE/eLPzq5
UfiDoJmeYyLG4Ct/Liwcg24gBmax7KaJS1Re7obdJCQaT2RVc68qQqVccWEuQKlD
zpGFAyag9xYWcNCvmPHN/YXXqS70uad3M2snttXsUPg24Vy4w/RZeyw7tTWbjk6Q
KzRw6MrmfLDLbwVGjudPETYj97poFlHIjPWXQbY0FcirxLQ5wWhfqQpOzN/Qubsj
n75J8tkV2ncsTsYduJXIH0IsHeQkm2g9fDZD3+vpMRfXO0PUDGN8HHuKy979F570
EuJrh+2jdnbm8mbAkqHqHrXSBzApu+NEfwYKxs84yoS/l+RopTYEH8mGVF4XHrEk
fnlY5Dt2ZlNyFc1NcrZ6da/FHpspwsUd5Ck3A2iNbWRhKGAUJpixMZCKmwP1y1QG
qb9JDtWRX/8lRRiAh0Jcytwnn1mYMyHGcZ10/udgFeDQ+DLcAJxKxS4XYYtbcha/
iAZ3o78Icg9iuaEQCreULaRj4j+ieZ73MaB+mN7R6ujeItFjTC/KDYhBxIi4ncfI
ONH4ckBB6Kws4Ry16CY2REKjmAGlQgaVEK6XZ/FWhmtu+ikbY2Yz9pxfSja+Nany
ba6m0Am9iIe1HNJIhNiY1DYWD4cY9g7+Xha7qANdnWCKo8V/jC/Yvte19IvwX8Tw
6SIAWx/uyZ6GkB4sk8aNNwEOe3dJ8z29eR3/oigh6RWp08CdxilBB6NO1yd6tMUo
C2JJr9TO8ppKrLSN4awVK7ewEOE35UwKoYJKM6dS4yd57sHWDDsEhTwuJoAif9FU
VrxDmjX9P6spYvSI83no28Ux3I04ttLBKYaIyf9zzshLdyhvsmE/4rvL8tspBVc0
EM/MSlYb08+CAcfapOgdOrqIdSHUwexO1EqP3KPGYAFlx5P9U7K/f7guzTxOaaRu
anW2LXOTt+IKhxZDu9B7KrXLe5WIkwJGGPZdLRI5zmnNtJfyz2YxMgj7PJv1De7d
HCq1v4sYz/SMoffqeXab3diZPgLV+PW1dmqtAxilz7qxsSGCvhHdne5wo919MZej
+wjp+6YqrPHxMDSaVGScNbvGs3XfrOrv/hu3ohVePaTcZGgAi6hXLOawMEATt7Vv
EUHK2uGnWcCIa072wu9nDriXP2kwLvIbFJjZQzl0K+wmAtMRjvB8WXVEqzgtKPnD
r2Ed5byo60sVQ0T37g5JHGM2PP3cpBqOiCQHCRRcYm4gKPe0jsOoGF8/Nt+5UEGw
lNO4qkTphRkZKBJ8hJnMlQeQj+GzDdUbUbEzl/9as80XcaRzJ/L3BBvYIAMtk3hh
crBtyeWRRuOnqvXr7yqzdhmb5T57LwAKrnhILXSImuiVaYpuFIfk40RNdKQFojmc
p7jGR3b2LbpmF7FShH6Z8JlkLQDAySj+hQQZUL1J1TEBB1Yb4MExC9Mr8+4HW/GU
6LbpKEzuyMXxY7BlR/bUtgcUAswMtwTzQq6W1oCvzLcq6sDkkYZTjV5oKe3b0bmf
n7i1Evq11GxFqwlFymyT8nP1EahoNe0wdiC8KpClhiN7VBpNSjBKbfuv5Ymdt4j/
FyVMRH4g10HOOtyBbaAqS3DL4XkWZecpI66EOB0A7IjtBsLBGrPcAoSt2RZ4/ebN
+pZJJDkJ/y7vZSBK/xujn0CJ5FCw82Hf098u2Dv2KsN2ApL/DNWsH7URHELeLyp8
E3n4prPmORq1B00v/ahZBh4x/sBCk/GKtYadz/tEe/RDYqAPyo88wkzf1x810s+m
COfmA88cT0X8PrqBDGT8pMxqKmVcpLLZGOMbv1CJQdyJjm4rmkyGRIX0n3drUSGn
4+PFYYngxpAr81IqoNW10mZ7kHiOd7Ks3rrFpqOYfZI5GAPsxTGGDkF/smv5yBYS
Z6xDCkFS8k/lrW+6N8uxhkHJBL4Oy+82kY1TfrzOQVIFBLea523ZCt6OT27OFANu
rRHcvVuS1vsl2Vx0AhzYGbXUny1pkQ305iA2O/WCQmDF7kXVgf0RQlo7bF/M/UR0
M2VIDBp6LASzvJR7I9WukWABDaJBiPZlFKaeBBwsUq8KoTQvyNPbLDdkqMyd9wNv
ATDYhouhiI8095A2Laj9Py/CguN+Nyapm3qadcPrY4a70dawN0bWkaakl5gFr/u4
GEOWPQGCGddLmg3VsWJSRQPNewtrJBphTahOyUpXTiH9C1keufbiy0zWH0UwEg/P
crvvIEv0etmhmf7qy+JykmaUJz8j8vV2hS2SjpD8Y0M5nPd3OkbbKFo8iG3K94dn
6N+p1MKuPjtEoJfg+sn+jp85EydQdiq84H1TWpmecOCPOAyjoaxuALX8waIjntAG
+RAA53w9MzOQzsNxLLbuFJzA0Ws+wlKvQtJY0A84fsAPTmOLLEkLbOPNh0xLpFyK
CgjlIea4AzqwcWBzmYLg1EwOuuHpYRqOUV5HrjHlzsMS4YxbjmbOEVje+tJQNaCc
dqbp0Sjp65XAhLmP3AkdlraO7rasW4Jz1RwDKiN5/VM2/U5p6sdo9uRuyrr2tNeQ
bjLpXbCTFQQrPt1tmPa2e5ds3byFKK1XbCOlCrPXogzqV+B9/JpCG35y0r24Sv2e
lLwqA8HlMWvW/Y/vk3ThlYuhnfcu8GvYAuTYE1i2ZiRTxaTOXBgP72lqpC2yZtlr
2wwMFv+x3eAQKZhOZD9i23CYGuIW40sJwihJuHFXvxEZvK4SXHHdjTvyE66CIUbX
nFGvRcGMfXFhFwHGLzTa6XUCJzgSo1QhuF95ByVc/jtZiBGazFmcxSwGlMM4FG6H
uEWeJhhY39C27eothB6Ft3Ku6VJhv7uGwa3/IGs425Uw1s2DZkoYrRAqJT3bokgD
lhgOg3h/Z6lAMld7WCXn/MAgpooVZ6G/gN315pmVzBniLDPD4SyBLJA6blWn83co
LQ3qVyklLmCLrEYPsYuxYQlCRFgEUl2JytN+WcYweKPfFu2a7sKI4Nccm4r330M1
aBCT8oqD8B+iNTg5vygV5klkhIz8VZubvxNtyQPuoaZAhCvFHx0b/5c1oAf0o3DD
kY+dR+Nfol1o7hOS5IPI2MJabdkfBXg6/OCCBg+O6Jsn1Eeqn1evAt0eRNCmqBlT
P41kalGwyL2RHUu54RULdmYA9WE4HuM7eBZheFGy8HKZx+2vSN188zrDRvTfxC5A
/lAZGpBAINPxdbyvOlIumEtziYwG0RWsdadE2p4MvzF7at1C5hM69raSKPb7T4eE
R3NKsyOKufqNwxLt950kwGiD0+VUZ8YDpdag5DqgTmU/2dz4DBe8OiKYTW/DZ3S3
RqO/8x3sPJZOTjrl29L/8gq2d0c+uV1TgOiTwmCd0MgS996W0p3DUPp2WuMucMcR
xGdLajU5V5FaE2go/kZB6Y0dXNl+i8QvTF3S/CH9Id67JQQuv7lVj6FOczdCexrX
y3zJC7ysYszvb3HsVZWctTgNQEASevvIZDQOE0pcclEnqMZblr/q3eJh7Bxp3M0x
MKHXiQy1ihJg8oLebiuGLNVQ2zTHDh+7qrCruLUblPNVWKfG88Uw/UIIfCTiYy5S
qWTrNJwFG/NzoasBzefNGia7addZ3cI2dTEIGD9KLsKWttB3rJoZxTkqUMvDCkRT
11a46ayLjCInp/P/F+xXBHN58fjjj6Yju12EyfOlaF2l+U1HscUtZkpt61qlpcYf
T1iz/KSE4/NYVFK4CSTQFqisWys+XDUtuyP3/bJzdzZw9eqaJ3eDAVwDNjIp5tEM
xfk1tr0EbjuFLUfTyBKjYFF9NC9c2AeKMtUfBN3nOAM4XFEcPxFebxJsMEctusFR
AWlCfRf5f1EdBoMvLvvm/VDwmMfo4GpZKSJRo6e8VVA/sLacG7AiRAWttkJ6wpv7
bcZmnlGk3+ybOjWGDvIL4FkNtmwX9yntGTWzpoueCeCDiLlYD91o12bC5vysU4jZ
gKN+MYlvFGdC7DAKIbvzqa3bKHiNSLwHGmu7LeTJ+59sIa3lAp+YqNkQtMfY9eYF
dLsioLQbYfIfAtMsSJ6xi7gkPxYLig23gjQJwUYHpALsa2lY2uIguBqKJb1kkefn
CnIWOUWO6QWLaWpYkANtskMBY+wa6t3/X7G0mwMG25ygEKDnLbx0CmitN7LsoZnU
lJurLBSYVDoxlxLsTowi5zEU1s8Ihts/Abj5QP9w2N7AqC9PD4+a4Or07Vq8YvHw
gZqNbc2Qc8NAF/d6gcGx32eqmU4dk26FaxDW6QBgsVHZiyKLr1oi2VsNOoeGad76
/8nhe6SNORegFUwMiHk/N6cE0OEKWofuiSS3vDfPW/JZnhbebPv2tw222E6Mv/nz
aEqFJ3EM/4IQFEPCGhJwgapWqb/64AVTU/UpTXPn2zCIbUpHiUHWwHNx4sKsVkmM
yQRUBcqQgK22ez5SKxsNIfvBsKR7oJ90Sqe8R7voUz29NDZX8UfFIF1yqoy8wpud
M2FD0QJnE8wQHCs4jozOIb+MeCu5S1Jv6HZRUBvzcrp3BC0w4MpnH7smoqspLSSo
UUJZq8TSGj2swfsKddkQTdRNira/9JFdKLlg4BctRTsXwgXEGY0xCLCc6XC8aG6E
uEMELTigWXX3gug7PPC8mVwrteKACmuNzB+jyccI1DhpDZeRUQKNksFwpUbokD77
f/b0xU8ywjLiDIV85LYcVq+V2FKIAOeg+Y1460gVIV7pOZzyg48tAadtocu0j2zv
ajkw1BSP5cUmXcoAcm+5aFSHgYFJjTksRqaNjbxV0ynW++0I07fshMyg3jwXkJAI
PpuyEG4Bm6Hq1ibAdDukqmpXjhy/vI60U/NbEk/t1fCNA2wH1WPlgbFXYGyRp5we
V5JgAQ2tsa7LHQhW2zwy+my7FuOphm48tYRJdK20dxHpo0gRljSJLmGs7MvPdS2h
eSCrI/O8+K0LGNY+j9HrCo2VFqDoHJrtVrVNYfIMKfQt+J0YmKG65WdznEXGEBC3
wAqMpSmR5AMiwZ5o8QYofAOvVKddD0XsJ6WsZFSzMUlvSagjDcHGl+HSWu1ut6ve
0csRDT8HjZCmZRfPD9yRgaewZti3t7mRfWyy/f9zcwXdhpicpdGBDxmYDPOGYI00
Lqg8dB4wxwhLa2eO41JUJOtyNKzOblj4UXa0agss/VAeoZ3M7zlyHRf9yIJUriBa
mjXoi5SH+t5ADidWZGKx5GtqAo5hZzWG7RThvzycSiSoZ1lJ1FES6hx+BQxXSXGd
icLJfDiHcgQfuNkHJuHPihj/BwW7t85mY0rIP9/dbORs28cjt1Cg89E4o1f7SeH8
uhGTuma8SEgLjPY2S/75nVbNZKIsNwSedWkH4Ym9N+JWxKWHSV+IZbz47oGtXHkB
dZUtYdTo3OIclZWxedx/kfv9rvZbO2R6q0gIMNZsihMb5bIr97pQZUso1G8aKeMT
qehwYvyWTTNQvi1DbWsg/9YFoSNdvdTVcADl2EVzbz0Q8cveNXAShxXiKOddaKHK
CpSvYli4SO7o2v2boLKr9bT9cyGXOWlPHhhzqAS/x6s7d9JJ77Ha6UlcW6x0Qxwj
YiRs0JbnXoXKe8k2tnzUgI/8XEH3NMlnjd+vqrPz/vNBsQJIFapfizvVHGDbI86f
vczMg+4gQlsYXrMosdLtEFv0DHUJlJF50SO2l46nxPGaelEdBlEMZ85gcmqZs9qT
xZ9yqgyCED2dQpw9NVAbXBdY/DERlPIlT0kgacUuN0vcd0cPAiWD0utlH+V17D7B
56Y6eb82FPwgJb9oKgYzUAmNphze8bzqCHra4VwlLO9afFjrkQ5FFe8RrTEpTnaq
EM1jlv5WDCsC1BKkJR2spM/ZohjZSvt7AswibUsp2oUDsNdgHoM0s+Gykz9/J3NL
kCJGifiA5+U9xaQv7msA5Z1u6GKUEwkGZGcDQ+c7zoroPUlyvQ9eQnudAjzx+FQw
4eKdeIURD5VzZWFQpjw+67EMtOwTZ/Hxh+y8UbPzFL4KrmiS41O/PJByfOfgKn55
SI+3bv/AoVug2qDjo6cToUnBJlzIiSMzfoxhuWDaFcd0gGRzidM6/X68xcRzIZ3P
hccen0QuuM7Co5aAeQaLOiqOZeL20C4ejC52s6kUw88m+Ot7LtelN0BGMJo9tpBv
r8EPBXF9h+W5tTLYwjagKjTum2QOd3Ei60qB0vLfxTZSjv8G1laa3VJpwUXoqF+8
4ceuIiuuQaZVCARP7Jv7tk08R6QVWnWjTif9oY+El7GUNKazH2Dy5ViJWC3wxsu/
5Vyz7JD4AP6U/D4U6NkRwrsRhSOqsMrhsY+/OWgZn62wz5CQpJzi8rRtOPIJGT5W
SARu6HkfsWKK2d7nP76rugTNQ6UMtcZIxRDHvoicrSMxGI/Rhg348kGE1AlOp90x
lpS0CMP92JgFDneGlI907XkbtW5Ng/nx7J3yz9ot4/IYdn7PcNV0kpH2dk1Cd6Vo
q9KGbAGHvHf+yATYvyMDMU45o10qSmZiKGjf9mYUGD975dk8qmDSMtfWkV1Q8B4m
0tupYjmpWXvpciNHP4JqYDt7+gqNh47kFRFEv3pUWHolatbbIPZFuIN/6bUZdn4k
cB4PMFeANWdDCTkrwgGmbw40f02SoDzBtlnliGRnAWXZS79P8RUWhtufKeiOiUOt
HdD4rp8n+z9EG3WgVs4muEIxiRcqOP04hTvudo+d/q6xBl0pe2rPISp6nRwn6NJ6
Rw59c0rA8gR80HNd3omXDOt3fQ8sIJaBSsy0cxDEg7RJXg3oWC7P2kPP2Ic5mqT0
O73WVtFINY7/ZqyhPQbA5VB6INnc9B5upgrvszBkWc5EkL+lo/YTUAFizl0vQ3lm
PeX904veXgyuSZTPNi6AJbbiH4Q7CsfFDRYbMe2jHedlEEVXs+wl+qjDuwh+l7FW
XbyeEEXveqW6DrI+8+9LKvuzOJC6AqkKc49dvj98CFMTuw7SKk2GbX0DCe8F4c+j
t8pingmKEjSomQTwxow/5M1N6wWlCJGti61XzT3jP2yN/aiokh228XWRcY093m3n
CJCfidwIgg9awGoIlt7TyciaRMEANxg+KHexrUugX04CfAgXgJtGtbxpID7GMtkh
WUaS3uFxVyBIXfYb4Uw4bi23VZ6kpLd3HtONhR+SvwesZCzPJqm558pEAoYasBbN
cesbhyJ3eFwZTjMlh56/HVZljnxiuf5ouuLk+pT6FeEgxmcXv2Bb1dWUVGGaprRw
Td5OkhQet7uu6zq+ZVYEaesclKVBToRsrMmxs7ex7cNQmyccuGoPSgA0qu3qBa6I
LiJZA5aQz5Jv+JCLqWUpU78xkiu6Lz/QOaKXAyVwgnQpDtb9X1IEJQfifwoC7BLE
mROKh1d5qBAHVMiVdKDAwH3OhZahsAcV4HrM/SLaDHtwRZ96IEvxlnr3BMARBY1i
33MZJN0fCdh8upDT6P/SwvVx/Njpl0/M0Q1Ym/iHBPoYiuEIxW3SEDqRGzvK8Vj9
1LBoQEE8qSSRjd7CK0/EOcoQL4bITrA0xSEmWf1RUZYHsswe8FD5arhEuT/NlgEB
zbrHdJRP6rnC0rMrms08euslDDcaQuWhKONE41pK0Fe+SeVlLQoTx8hCFYmtIXks
SRgcEAFB2JM26Hpzeecy8BDdcyNvQ2E6LvcEB2BoFfRaPIrL4oAoaUKPkqe2wyvc
Vqar0CJfNSZIorw5nq2qEONFTvFiO2k9BSSr69rbWaEaM/X99M1rCApoiLxYUkhT
olnDeIPhkJkFJCem5R1Pvo4ssy1/0kod/yzK4fSxOVPTFtkXhHAgqam2rTJYoGgS
nG78wKjNiRiQIXfPXMh8sy9/O+fUl/6LkmtrLZu4U1IQDnvd/aDT2D/JBp8LJWZp
7VN/NU9EyrJtQsRvuIVgC0E3qyQujRDtqFQQPGEm2wUcQUc3sOxWvuEXWWTbmwKL
W3tC1Pm/wvMOjgO16LgUa5+7Y3QXSetlMiu62RqCSiu583v4NrK4zYza0DRZ4bpx
F8XCL+qWhFu6rVknczM3Egly33sptXiIz5uEKSpM5XiG7jSupYVLpG8qJuZKRaBv
tPHTg9kStEZmDoKnKaFB0Uzi3LM0Mj/62fWxYCpTS848/0D5b1+5f4AeMBFx2vkM
uoxNGEvQInb3I9ho0c7qSgdws+OnPDuXdHtTQHotjcHJw4+ok5Chm+WjcREqMcdh
aw/r26p4BY4p1n5mPt1RzCm0LNVXHe1Fl6+fhcU32Ey3fM89c8vskAT6pbQQJ4AQ
1b2tLERJ7HRKysiT/4n9KupxP+gbXYZYE6AuicwQ5v7ZMS9qjNgHxcyoXvrZEVRx
fvJmu5fTN4B/kZHgs7I2jKiZN9f5Li61SnD2bgFYllBOJ240nLtrTY1zEsejOxEX
ModHOqEPz4fxGUrMtXUifgqHxvDeo655i1XSOSdyfO2vAY0RKdTIhXLp/Tp+01ft
ba9DprRlR9meHQ3NVefu5OTiAwbwLyBmZ/GH+q0mdHHliE6pjquAyBF8HBQbJmCo
j/s9Un+rIKKUh5nV+Vr6gLaTpa46gQWzUZ/M8jN83hcim1H+RZ1oJsHn8VUwIbjR
7PTsaMcEnFowVS27wWiLsMm5+q2JX0F6aINgncFhHxbFdQZWBYmdfUmOqk9t4e4C
hD59KervMqpVX/yFe2V+BgIsbaC8UEzhMZ+04Lk5jlo+HECjUPVZ6/awCwWwAsGV
6/toUpdQFijQPK8YCBdy4Ed+3JCz7knAgCfrlvO6TYQ0hSssWwUKfaixsEyYg2MP
HFaJOiNsoeMMYyAWFb4YEuUm6hGY/rpuzbEQLXsQsxZkg0lFKJAoiE7V+TH2NxiF
wN+LPKFQ8rm3P2PpynNuLH4nr/wkOg+MV3Vwb/1B0cEeCqUwxAaXL4g0+0JcaU8Z
8FU7UtDmu+7ECuPE0wre58tnGF5J3IhjKs0fEOFwbF39HgANLZtDTkpEN39loZuI
3WdDI/RryxsUGDy9Hr8hbq850YaHzhIF+JHqCR3iOqw4bTGYihrcs43DePHsO8Hk
sWO85uh0zNU5Zc2bgct/QFMqChwRV3E6D6LvOfwvP1eHO0CSYgsA8pFcc1C4bWm/
AZOOZkry9IWbLr4d1Z0bCYj5H06ByKsKx+UR7z0qmC+9n61kWL4uJ/2Q0EhD2NPA
fh1HyNvtlTC1PQnkt5g+2yly4Sbc1vi6DXauh4G6mKR/Xa0dHqlIu3k9zm1xLZf/
Cqvg70CReYJWJg/OWIRBk5+MgMaIFpuQ5xyK8WmoTYfuSriDxF8ZJa8Z/0dylA97
cI6A2OjGt/NpsXPKVJuqHvRD/+tY8jSilqUrUMXhw8BajvEPV/PZiTCIMxSsqrw9
KUd+lIKsQPhLTeMufIhK52LYHlrth2zOHyyH9VXUMMnQKz+4DF4RRKlfdyGJVcfd
DnMg6K4xaf4+Y2blK9y8aPJKWxCEb0YtmQkmi7wucszGK7cZWnfEFXQRpj82Rubf
6sPwFpzO2w2lxB3r06rSuflPayuJfuU1YcMEVqUrIqaWj+ErFGoR28s8KFX1XdUe
KQ5XHm5wnduywH82DiZM1u195Nq/XJuFm3VrZ95tHYaLcdLu1ZT+iN+SDAmZaH8O
tYw4qyoTBN60ATWGPbqWB+cELdmGjoNrSHDE0ZOkUy0zE1/8e0ySxnawloq9wUOM
k7XYb6oCFIcOuS2GXAMKIOwX5gIEKHTeXVf9LFWDpuwQ5vLycXrXqTjceJu+gIm5
oy3yraKdMkDYtfoO01gLRVfyuiUxU2mLVxYOLaVJFOPlP4dkEhqelYnpP4YptklB
mLpTycCu9tvD/LyH47OY3urUWWOP+YWnm5zh693iPicoLavtxdihml4lc/srHj06
VdSfJFII8bSsZ7tcAwwXT2X+i4RTrprECcZPWD6ZScdg6vrI2+1bLHV2ZbdnJ1dx
WPyertChz/+EAmJIy4u80kJAxiFpDvt46WCBrhgMpwf4cqBHs1TPixZKev9XADS+
c/rI8T1NeJ20240wCXMpyQb7rsUCweTEcQldnjzSUd26SYPprO0JgzU+GGt11UWJ
7PAzc6nx/DocODgPk5dwHjj4HGi4ne38QvUGb3ai+VzQ5p4sGGTSyasS3QfA9a3v
Bo7nCvwM7HqDRHqu04fCQ1QQc8De1ThxrbJnVzucrcWYOM+M5Las5RO4G0H4XQ8b
BUvUbOjNNUT/HTeOPSfXcBhbJpC1ACA1kzv+Ve/5fevNlRafybzmKADRbtedFlEk
vWLQl+qqQOzYjFMcsRCc7gUf9wSQg/6JHbIx4K6uzTcE+6Hp1+KkpZJnqTkx+7tv
4txrzDYrglcfb6bGYZcqP66Yrj8DT1y7b4691W4g9qfA2SMM1O9htanfwpPKGwir
LnevZd1G/+CFlePeaVeN+ngboNKt5P/ABms+XGPlbTIZjKYiCC/j7ZSitRLWK/EK
awIaoJFXnrZGUB/gZGLuDEol71cRK3BNlzP11iMVaLL/IICFZsIFY7370f93h9De
5n39luBNnqFtAJ/GhQdVDDckYcSsBxeX4uulZe13ZPJdPZv0xtn+N8ITFgnms7nC
WtKw+L2F/hEMihgp3JNDOj6lq5ctFUvQi+SRbbshKBm9nPYtezlGdSwfbrvrqXSE
GBaFmOePQjbB8Cku3ZkA/Y3+lz05rOZOASmOnUg7VMN0vUB5ot2kGuLkFKdJIztK
B7GbABxjgMcllaY4r0Fm3ZNj+3hVw7jhDR72TLY7aRrjK1mkIlDGobO/ZMBDPl7O
orSE98rvmXHyFDctPBG86WTTzWymj2/jGcWDiv/gNJMmgEHgukRW1eo4Noczg76S
AuYMCg33aoGWSWrHKhmyJn4KqGfYkexoRoMtlwEo9Or1c0zQInEls0CjyfYX+rbU
5hBzFDnB5umO/sh4F/MJG06v2rLXzL3/NHLG+wVVOGwtEJrOA8zENbROpWn0GIdy
V8eKf2eyzN7fQD5RdgeXO1bnnR98pzvAl6NmVJ84rJuodZqNIPy84VB6RxZbtabi
BpvHZqZ6BUgYaXRiqLBq4IDhNnQN0JrHz+P4GbufKvnmuJ+5Vzv2dxhDceRtSOpC
VcXzPQLWqd6nTGczoYH0WPf0wThkOg4Nju/kBO95zX/Eq9yfyzLiK0Ax9FZd6WZI
f7wldhTIjPakiofSwuv97n+3CV0bO3nvXVX9+yMHkWAHarvg5SwIA0cp3mJ7ATkl
q7bxDrqk7ZaeYM48SHRHJP2bPjR+RjQUSAhYoVqhwv7kaFJ76ty1iQBGFRnQPY61
xeECMxna7ukKbuPusB554I0kkmEC3CcQ0jMkrrzsPBO7g1PNLFxNjdgcKOntBQes
HJyqeSk7UD7Utf5ijhErwoClpdOL44W0M4Geh7Ktv7d+KFB+bJCEMNBp/xX92Ms5
17wmalbofXKoTjCLwwYi1Suu7trFRVZklV1BYeh41985LhPaJERocMCsNW+Sy7QF
4SfrQ8eCOYRwmI4o/MODbjyhkx9mo66G+2Ix0buCR48/lkodBufyDEhpYjnlT6FJ
J6LKfAhsRSPqeodqSbf+pM1XZsk9ct2jFD4V2YLm8qtdtgj6f0fS3kdPX+xcqJEp
UM3VWpZ9M2ZRWjZN+bOarKWJlz4rQwp3Sgl3BkrcIMtPOwnT8OhDwyVCVqzUc0r/
jzYEG+JrZaRYL0Gbf3DsD+MBwPYgFisHJrYbnQEKFLnz+FicasjFg+q/jeUGDEPQ
XO4CAKI7QVVI17lyZa2JaGaGY6Lk4bwRgVfCuM+gf7yoD27YSDE8rD/3AS8iyPsp
srdcE5tVX5MXgpBYivP4AFsiv7MqdnMg39GvoyvoZO1CGQJTM9LVAQNMYiSKhTXv
JXSt8lvBkaGRFNumkiWyR6dcGMXenZvDyUBwAnOUKHMokoetNmNjjO25vYtGJrH6
LXLvBnOChG5OaR3NpkTY/zGaxuQPLzwUvoIDaqQ4AZJ5G7M2Que2dc2chUmu7cvx
vP8vtFQpQWRDU9KRD1tvHNzXDBiPaEhRSoIi2ivmUbfHK3mNSEewzW01isqO+a6H
dvuvqYHO8LrjAQvZESig4tvkfJlMOMXDyq4Fv4F1TZ4BkZgLBhP+bEhvdXtmiW8E
kSWYB0ghGNhwQ2DO4p19IrmhK6OEUTZzX70VbJPFhg/GFdtF1tmFVqtRBAiJWWVh
Vs+2hvIh6W3gaDN4F0fJz9sNG6X++n3b86ypWX8+uSVoMxumv04pd14eabtmyfMv
P7WETBnk0kfAa6DBYCn4bV13PSkiBNrS+AStZ82ExJCgrAxuuM0fYtXpBK68Zb/3
ViFyJ2bdPL8go/z/l7AwAk8ChOm1AFu56gRW1aJA9bVTfpaliDhdIQuo1RpFRYIH
USIpJIXV3ZZFH/Ro3X+8NEpjwLocTxk47dDKit3pgcvI6JnLZLVj8ECIySegmwoL
qwv0VxDqbAKNtrr53oImZYWxwtoKcEd8nKneucIMsYZR3Qv0bYTEVAWIMJcH+xgM
mcHQKWDtCFjQrreFt9tbcs0mpOG0z04Gjabnr8KvlCzfqeHwiMWHq86zUSgs1fPd
HubEuR+mUqpKCZ49BdjKCZEThkHw83juU/DXzanwsF2yTyC0TrmRK358Xj2IAJYI
2CHqkt6CnhwlU4ET6AkrhJIT5RlfP/kS/gPWzCSGmfdlIPKVcm5X7THur5LOg+c9
xRdO9mgppPrC2CR13fvwQgxS+WzkEreWLWIpj8smDpuzWHDiu4cI1bsFi/dhNFY1
8uROAUU8Ydo3lAsrJGcRrDprEVw2h//c71SebUwmm86sCXVkEySME/bxSmedq1ov
+cC3Rzn+nYrFNLAewBV+SKk0eVX7YhOK6eY8Sm1x6pTXbUpoVxvsQ73ZkvBbGrmk
zVxnf0PkWr8v3zdsr6iLhIVouhAXYOtgk6Jsj1yjatlwyv2uA4P9DkWUTH3so3dZ
dQtUjJ8VATaZcV/mjV/6qmyL06rWUyTGcz3A1TfWjUpKqhoPZQm8TK8+q+wbpAj7
5eRtuXEtBoWb9N3qgikdXAFHOn2sA/V+YM6//1JcJntlaEIjCHrmP7So3zYFzmjC
c8lztXrtE7CVWeKNGsfpRfRSSDUgb5p34roN7npxy/z2yh5awZ/h1L40fD33rcb+
AwNM7ztTgSfRRxfX8DKX5zgaJa927FqpQXjzOOSSyU9/NeImvwu2Lm5iTT8lcSc3
T4VgUTaiKATmefcsD2JRkyITsVKwE9zUjT+sTJPBP9S8hGfEPFVrLBWm/fzTatcP
QSAso2X0XV9RCqND1i0YpSH6WCKDJRsXEGyXVMI39/HjkDwsC7aY8N1Y60UMSLYh
4OjipM5aNJpmYaqWD3QHaeYisbW2pdjfcD3elntq86jsBH4yzBdT3eV6MuGPaRAW
I9hH71OapFtH1jjw3PyTeAYhFd7ezUtO59ty8n18UIUSy86l9awZO+P+lCUaTbb8
xgQwDLrWg4GKP69umxJAPt4x+Qy8bqqiQQ8qDY0esmLzf7yWvNHHQj86/0dAK4gY
29nRFS467NwcVelIivN+V9eBDYqrUks+/HCQ5ZeX2o8yLjQNB2DOnsbf6s133umL
anNgtdJ9tLZw09U6d5YJVZ6RAuim8xPgWSMrmsOkUUIiAOxNhAod/pp+qNSolzbn
5jsRdS4Na8FFXY5hBE7/V2JmEeiiAnfz2XcTPscHcWkIGaSYhrukiOWKBFlVcEyh
cvaxR/B+2MvY2gTaCs3aRsxToxpRbuPddkh4Yb+KXOY4MrU1eEOxunIrPnFCWOqk
0E9dUYdm7MwgXYw2COGqm0P6Gj49IP8CdMkY4XZWEBGvmvB3XpDMKMpFzc05X7Vf
xQUo/xYiXwjAxg/kfK/Qr87smpnqrk6MDoV8nK5jlU0B+x63WYAWTOMMH95mQLPg
RfxPtv1qtimeknzPwIdDlrkb5POEBEMtkPWNvhau33y95HuZSiLvhCZYwHUkDDQF
2Hb2+gPxTP691EDXYHEwWZCnBFpAE+taiyNUbvvj7ST0I2R7G3gt2OIwxZrBvEvB
mXPHP6IPRyRFubxQFC2IINwakUtzeMAsN6vIUXo+agHXqJhbzpRF7bwek/SOkEnM
dSwzFN/o/Rlc9k/BG+dCZojlYVx2AuzaceM0GtVB23gxP3UH2gdNxc5BO6LbBglw
EwHeY/h1zVIalEMRQuL81AwLQgLUufVG+r6l5PcrwsQCpZOjqswJ0BL2n/Y6w70C
Tv4Ns7gMBKTAOPMlvUV4fmhd7DAA3mBQ1NLclXOIRIPHuAVNcqU6zGYsGyaYpLxN
AP+Z2nMUMDPYm6Z2BROcmT6dyxe+PdU+AxEZn/e3gw1M2i7Ur7GzHQf3nNrwCfoZ
aYULPgfLEj3X97//2bi9NimoXTLleUAS+t3mAeu8KLXroinKA+mp6d3mZjiE1sQ5
v5VCko3GB5P+08hr6zxsb3L+Hv6eP1MSbQLV+biweC8oPPkPVCKnOvUieHT6KDN8
Xrk/l9vboahs8q6/dl3oezGMjvZhWeqCNeE/uMxRvr/W2yu8uDk6g0rfffzZoGKd
EFFvrarmSLz4NSUMqeuY8C+GkfxR/wXxu8DxMc3Aw7Z5U2WHpiHFUs/rzqfQdxcb
c+GhE8R/4A71i20BOYy6CBK4dpBcj6K95Y7N8ivdYXTUfzCvz4piDImbxmMLyR/J
rp3ve/qHQyWA0TxvYrXRDc9pVWTIPhqT4uo8hlgKDxFjTQuXWEVjZtab6SIUi0Lz
VGk5edObJZM5PmwSGtPolxbxIcC1B31fNVaC2JJXqLh/HuRWlzRXKfCyWj64+uBV
raW2UYsl7qrBSNQtT+uujboNTs4Ugo5Bq6JnWn3w+/lB9F2m2Aax+uFN4uZghqqk
OPjIVzY27ZZDQ6Pdqu67nqkM6+yoyeQmitscuKnXuOJGjSXT8JhTbMj6/LWunqIK
kcM2y9o5Vb6mXJBc45D/JkBTi5nBZWCmCv3flllzy1Rr8hepzUee8f9VWBqmiwR9
iAmWiA83n9rXromw3CXCh2dKXDgi1LvsTyZJJ7J50q0v/e5n9tAA08Mn86F/tHwE
zQ7QMB6hSVkeRse7xwCiLPrUwJQeWW27YIOZnTBFuGVmHgJq15DREe4UK9HLQ2S3
rH6vSgGF+EaIGFakDFXyrzu9Y50toS8D8GHQcGidK65tq1WGC1ZEwN9b7oziqwkv
gRMp0opSI+gsDGKzBbcJOPFB9SBKO2D+y4uqGbXke2HfiHtftmrCH+7EeTeOhh/R
mYRcs7xxR/merzmM8iXTCLlwhvyCruarzpUXb8C9p7XJcJPyfBr69kL5jJfF7Zxw
c5g/25pr2WtFW60NYKmK2Jrl6+G1/i6A1A8N8+VmRyGnpfcyWUjoqLg0Nzc5h3JS
Nw2pBBQkS+P19KT1deaOujAXENgfhz3FzCDsagoGfIOIxI74FvrewI3+bov6NGQx
uJAkklxcWlTacbBO2Jol+wPO2Jar9LAVtcead+bdUA4/CPcCGEcod2NFGmsPwJM1
hGYU39qfwcwBywZV/N0RKT8JsdU31rBPC4SBpdbsLgSSr476Biif5LAnAnr0YEbh
JocsSC0CkNfAlwBf844VDrQYiJYNNWbBQ1m3BRWKiV5gU/4Nak1Wy9QLqDCUHOyk
t+Gld/3woRHwgnsBHIp1jH+J3KclblHR6bkpvxb6kELtX+9AFhpkilrR4/VloU0x
6T91sIA1d9tV3ArC2H1kk80EA/D/d9xQz8C+M7Jq4GPVHODSK4J4lGFXBOZ8mIGP
rKKzipnjVtaFpOGZRctqVUoeaAR41A7IdwySycZzWcS3+ChLtLFB497jxG0QRr5n
9VA2yEL/IPzd7JWvAME/hMrr/YQqWlbSAUW0SPfDL4+qnEkYjlqZxFP3u+/f8vxz
mJ2lSunvDZVC41JQmDcwuenRMp8uh0XM4z83PFwHocnw8AbAhJy2P10lg+/z5ctY
SCukGOU13RqtDCxsv4/e/62hJIDoUEHawH2SuQwMk/nBD1xxx5Dh/kXGiZyiL2kM
BFKU7heF6EYGqrcm4PFQDYEe/TOVViAg0Fu8lexu3MQuG3dToLJgbzctAXP2QugD
2her+iohaLftkrgI9esBg52pWUAR8qCS08r0iXJoptETpYWRbQb9AQOGzo3r6KTZ
ReIic5InNr01ktUd2BFbv4gSqZLuGWEFzJV1FI9GRAie4QCe20BjeVHepyhPJO+r
RrIRNuECxKh2OG4SsFpLlVLBnOaZ35EJxKCCkbF9p8MgrMz0JIMqN8HnopNLJF7a
ZjHEJ+ueKxqw7DCp3i7aGat8XLCmYtSN0KFbeMGeC3rNqvPtJg8b/Jc0CVku+idc
r1Mb9+Ukgb0TEdhTdze6G+5gmY1n+ahMo1RY6C4vjvc6GKuGOVZ5vsAkq0KShm8y
2QRBQv8Buutu7i4+0NCYde4B5uiSI4x7pNjKmbj3UX6LJwfxMvNglK4wEGPfBVhx
k8G8HNE4IOyp1IlTUW9ITkEWL/IRz/oQ+8+AETatSYz60sPlEl3lMu8g3nfh9X5x
5/67EImyxdc1CpwYyho//6h06EUEYr+BM+EfMByDlXcjear7sgcrCLNj7D79c9Eg
RpgqAbVfbUGF2jZ0HhizcFX+VsWsJOHiNZaypkCMhOnsjrBt6Wr+tg84ZBrQtyiD
su4CPQ7t49qz5YlXmNUFM8Wr7TIoxvfKmhjEbhAGdtziCTwj1HqUc9tPN5FKNzda
42BWJ9Q26KVO4RkU/bl4ef6zde2o4I7Q2WTVNVfoACHMwaTXrJDCpD8KbEJDMgtb
Ge0R06VFs64UvgNEV1BcM2KcMOrnSugGBgaHK33B//VyGx8jHfnb0zCbP8twj+wX
j2ou7bMF+f9IijGezM2ywgcE8itUdr+oDMaM6ydtQDhhFJ3v+8zDJLb1diq9l38M
SGUmJ2ntV4ucj37NIJXPdSmo6bl0bo5HBjen3wJxOe6FL6EbhXyed23SS9306Cp9
mhcubtuxtKXHquZScF3iXrVNfh6T4b3gw3RDWxeotM65pqbuA8ettxXtVDhRV9DM
4+wKKR0aPY2pjEcua/jXivnNi5wiAbAUR2EcAwzlTnjZftCy+Wcw4C80zziBePOE
T76ktWZXwOCWaeOmXnP6wL6wnrHUaZOy2LOasCfblg1QoyOo9xFWNabzZM17kmqy
T9F5MqYwe/ijqza3O6WsFaESMiIaQOkIcBMr2wmllsrs7bfWwBWMlKQIHuLYznyB
8pqB/WuXYTjChaSOAFYgWDROAgMKbnQqYOQkPAu3v/gqL0Xl+I+OogW3+UR27CIV
NDOm8X93BE9V/BLcegivU37cxV86tCEOycO/S5Nx0AdyoLBYPf+PqeCNaUuOPbX2
g8rfulkTZWV6lfoDrrlSZIAgEpI46N/S1M8B15hh91gujqChtUgF74gujvQ5iBvO
fPDUPg5qtKJfW/MMxuIlRF21O6s+aviJps7iWJQ6ZwR9oqra0NxKIeJ2iaFvb3Vn
ecCdAx38+iO962J/xbUseLmRcYCwU4hwBJo9kwxWz+nk1skErmBVN+/Mewv/uLv7
65St5D/nUC9FCQV9FNCkx2/vFd0pTAjrDPmrWZdr58+JXjMyNOcv5sycO0boaJOr
GXaFAfgMsxb6Hf3DJSlbxg1gBdZn7T+4Cd95fCcf/DSQYbcuEnCZADVnR6bhBZA9
U0gSe0BSnzsJiSEMo2eRV2D1Gn4wPELO19Bvp5KwwtgF5bWTmVj4kZ1OIR/y2DIX
D0FH9pjVbhHZHZV9wNKzUvNEKCEvvqBGea1djkJGIiObgJvSvir2cms+os34vJVE
zeFOw+xp2KTCWdi6SHi2Z2ObEBtFpXm4LatUv+5TOp37dioohmTBb9Bb+8wgZwqo
b2+JMG73fQObJo8ObUX8hHzFO6GQHaDHVY/cS+bP7FkowDNtNXp7mdg+6z4S7/An
d6lyGHbpctC8xkTZUYN1CnGyYZNg6mK+qGg7k6KHyGOBTG6/oLsXFWxlemXB9xQw
EdbdNEfWX8RRWDHThlS9hQCAtI6jyZLX8fS/Kyk7Df8aIoZz25dS71JHv6Mg7XsT
x9D63LOmfKNauZc+d8qD8jx9ynI7ndd7iM4hqqt+RPTEJ2ilEbFAIe+vLD9Qfun+
bUBGH6dK+K20A1KBTc3ZKm3VpNtEDUzGpdgnehvQkaGWwUnSB9YrJoAteZaEF5+s
h1DzaM9PBvx2DxdcdItQmr178EaKQtFIAc+8FIFy9Dtx+FS6f/gJZCNoPivlB0RQ
mG08HDgcro1VdZ2g5hb7XERmXO+mNqndDXXP4D3n500hEtzQ6kCWxxB6JvLyZTGV
CzKWVFeMu6fChpYAN7bgvA1b7tJGQ0DZl1199NDFFBePl5ZDz9ljP5XGxYAifItl
Gup3Cd23Zrmo4mo6hIFw1z8N7JTHKR7tcCWKffkYql6x0vUasaVbjAu5bqsWxjWI
ffrjdTSScQsUMLn/XMycI694FsThy6TfFt266y2tTvi7+B1fihmDYwpdNZCjEbqp
yNzJtHoSTEdzaR1RJ1XdpV4psmfi9EkXItcyjCsdHd+YwzIreff3OCOTTxVun7+t
ZGFLg5NYIFo/3aYoPF2soNOXjFfh+BShKys0w3wqr8dPrHpwO/I9V+qR8OKEs2UC
sIjhokIeQGJc//tRxh+lyCAY/VwCr8XureJSfUpiuZEM3HtpmPKPhHpk2lQ/mYy5
Y4vEIakj6bRzU8qxqU33Y2/uxeZjjsTQwLDynD7zb6CUDSSqpo/HMAfyYAKQxpb3
PrCzwjl7wgt20hE/BpHjJetZGTlT9VqdDoeX1ofEdJokBbX8FtJlQL5UiAkJXd1D
L44F4FxrW2twMMRWTR2XVse/PgQjz4xC6f0dt0StBBEJFdDwz9uV/Q32o7Q2mT+f
uf+96xzAKu738kJIRZ/TMym1frFb9S4BmmeCKGDX4jaWcs2CoDrBY1F8spqIAu9f
6gZD67Sq4K+YlSaxxkk4rTBNpjPjhmviC/PBbmn8QaC2NId5rpeOoMK3uYT06nOI
Pl7P/jNdtKffDPgSFYPk25mr1XBg7aFJ3erqcX4QVnQuzW8sTMC0nJuLDBA2lSrg
C6jMZOatd5cq/tkBShcfqLYFnQPh/nNZ1eMYiL46/gOJ1w0uVmm8DsVlv+lNrfw3
vI2diSobZAKxxGpOX8rQt2WbdKPFTl72AeVYS3yJ1m22Zz8K54gPoWwhPfdvoxYm
cjxpL+ZsI3O1RXpKlN6WR45o18+HBaO2oaDS2Z/dRoVjtkoarprQTd3dzeoUnFyk
jKWIoANWnLUTpRaasVkR6gEkP3yJTcWO/5nm6utXp8NFvmznjqZAq1HN6xJhZzzO
uY1b7vTnmgGhhcwnu5JfZB+KmL/oLV2rX6HYHuu/DY/A91sXVCOXE8RIDBE+xce+
KLcPataD79/Cg6XGh93/eoajvyjW0UtxBs/j7wLzM6d7y5Y7HyI116GCq0YM17NL
tXZKF3HitJ3lSQXoZBoRv1xWwZUgDLOmg/3cKYoicqqmm8htOrGDHftq/gbFUw5v
cWJNN621m7gusUAb607GX9bezxEsFt6bWjegHU+SiPoLh32xSgrvbPh6w8wZ1Tpk
+F5KpoHrrWPbKgdHZJF7BBPB7OnN9utpmzDNehn5qH/ZxUbMe6zCJsqt705JlhSP
mMGCa0cdIkutjqm2OSKeJfP7TcqnUb3+OHMwnEne7e1oF+vEAyHHMbfCZXlftVAd
utTE4MCqj2k//GfyOQduM6rXT62fqcgdQaZYZN0tEIjL0mjT8XXekDcaiowMPyJw
aU4dlqg3W8cYgqsbYDMjJQ/1q7aKJHivgQJkESSh3qFFSRr9rz0wpyM3mPQrSG9P
tOazlFp/okzFPK6mn9xYhKfZblpAdoM2ULvbY2CSDjSxgNW2V9gNb+aqvG03XL8u
Jqtr0PECUtPbyaf59Yyp7R+GBD4nxzmeYbTTQ40dTVoybMS9vKEfZc7Tm8Waum0S
yMpos1bUe/IBapTajoGc2fx+wg5Ax/7VkAynVYgPTBrXfvj31zinpab4HsSlsMwU
gAl/pDvvE0j15OSsiCbaVoIfKUE2USJhqkVSg7iiAgoshLbxtpmP3Vfzw12XXbR8
HLmo8AyQBWPRxoHs2bg2M2JHFveUlgwQDN6I4Gle1qbeagjecDk8yYrNzDntxZUG
Q7v7HC31bJryuTYBsqvRDC8P6HUvHdOhkbskfaV0jzLW9rkF97X4Y0WSMjJwd2cm
1PowTZoLeTnSfURKExYb2eTRRkDfSq9H/2fKSeQM3+ZLLHXzfe2QBnKih1+g3Et8
D7UsZZkjbQFqZbRmUg1V3MbwaDEOVXFxIvZMt13qY6STTYOw3yzonHpggjqp6Ng9
oeYClHMaEQ1gx/yjLREZv3dIHyooyVXS3RdnFS/1LGPjSaPTplFgNe3XAzmdFWCr
uL62odCXNviIJnoHejU7V43ybWz7kj356mevvkGYUBt35UipN7Pi91PfTTsK9x+S
kz2O2l/ptw8A9YSaadmlwmiGdsrFV5u1nwNo8/8oF2Mwnwgk/AL5QoM6DuQNF7Bk
9vMCFuNWUZDW3JjCUfUwAobq2jLo75QdD19yCTkclPIQKljNg95Dsi5YAfxayI39
AcAx6zPJKyW1Gy0ogBBiMB2eXTnjRZjpkFJy/LlCgf0isjDqa7opzB/0CixlrLAM
W5gNhKbRqIgD2M0L3UVXuqg9QMVY2q3VujkA0TNthhRt2jlmGCvbnsGpWm3dwuua
80MnU9UyMsrQrxBzvTm/t6oA+UFopLeogjeYMXzzLIj8oSnTrl2h/sOmG27fFDMr
DpluK+Sc5DQz2jM62pyOygFp6+oM+dVT0A43L3QbjoY5QnjbzlTmH9ckQUX8ynir
nnUz6pFK+/SZffn4RF8gtXPL2955DsRLLPeR7yRCyCN2T+t+OoFm9ouoTXd/O9sg
8LKYuqE0yhEr5BbW+O0pztfjRYOJyOjraxzcu0dgt3tU+L4rmz5ZDf0Z66Nqwokn
8+ORYK4STwPNVY/5BfxgXfkt9xc8oUnJyXynd45yYdfdARQhi3tTE/f80ev57Ku9
M2RabjDGHzQpLEA+gad3ZEIj6NehlC9jPQ72eTrLUiAj+hCj4t89EIKtkZe6IP0b
fDPI936fpJWiNgq/DK9lH9pi/wqSkUCpmFEeeIsAzpGaLvVZy6d8cvGcwKxTqB/I
JFlArNIDrO64SCtoAnVZW9xeEN32MSCOQEhyHspiy4OAYUXPRFIwU8vPm2TLD+DD
PAvqsxAlAzDmgyt+3+KGjwhF+f48yzcfmcVW8t6R/fzvJmr3B2vS1CHlXRIFr422
mNt2DtExSZP1Y8AskTUMHqRw5fwVff7bUhKZv8LqWoRSlXTaniDHkBDNcPpst5Cw
qsFoOKEH+aU4s/fUdQ1zEWzfaquYj4sfxERrC1LZHDgyRTiK8R3howH2MAnQhHT2
05Ww26Nfe473HDkAAdW9eSb0fIhWJbR+5eobD0zw7SvCWE+Zi2BSPpXDHVYDzUcP
iZIqH351BOWaXapQyfsVizwJa+1pEvI8bs8ibNHl5DQ/HMVf4D6gJ0fSDvvkZv5s
Stk6V7erRfnP/Y9WTNLZyWnWFZ2Wb7r/3GNUx/hKkE1x2hZIHBMHuDUY5MYkB6RC
A/iENsa7CodNxpeZwoVZV45/CV0KvzkxV52+GOM8utWkWSZkAL9CL8HIDFN7Nc1C
kGF0wPaxspJxx86AbvblXznmseTtoLUWqwFe//nv7oWKdG6jfoCaaicIRhI06ts+
YmVQy2CYscXn2IM3eTgVT0CLxuPKCUrvU1czADtTVHGFBOOqmpi5YJE0efi+hODO
WbkGi/O2vAOD7xCkhs/MZsQit6/U3TmSwRyyERu4L6vM2+xfy3d3fMCnRskQ78Sm
Oy2c014TlnmIzvNZ1hYMVWwnd5+SDQeMLDL0swyJ28IAFsdBZdJB5LFzR3g/5clC
yyhgCaR+77ZaO1K/09x0i309fe/BlelVf2EUtLFdhPYJf8P7EddzjFIRcdX9AdjI
I/KeBYiPCP4wHiBCBFrdcpU4uqg/yM785eF+M1dJKv0FBuuYTHoqoAu2TE30ZLwH
6THQ1mc/aR7iL3H9eYQRHzdqHbqpyCQ80VGFOHd/j7iPDufHyHLrxNqV5Oj/tXLa
fFpoObY63xNKE9SI89kO2q1vztUQPzNQVuzyadEkuSNfmwtVbaT6p8Rdg9VZ3ulC
H/pdx9H8H3lLZVm+WvfMD08jQ8U2lawv0xEuYOeYEqOKqGCxEAamLHe3cKVXMwHp
M3yGMksmcmtufQ/qMklL+ntBYtlXLTiSyCsIHNaZJt7l3rqfmAFoiMKhhiP02kV/
KhQ+X5gULCxJBN/K14CVStHCBXVt80Kf5MuzUK5kDG/qHyaGXQGCihwJA0tPHUh7
Dnowc5wkU1HX8QDiocM5wut53TABKaK7QhBFPTAuLidS/KH0vKZobaMEabl3nru6
qIDmF2WGCO6SifERM23sF6p+gro2AuZu7P2PW5MQxvS3JW7CvscfQO85z8a0hU9T
LjMMTt4ceeDXBTKgk+017+swLKK2q2WkgVGp3wT9/69MP3EzPg279Epcu0Lf9sTn
lzpKXwre+3pgqMc3CUBdt7IqPMmfCksMh+a8ZrSPb4PN7QeylPGqX/J3pBUIt8VG
/YWTEmtKW/JwUfoawA8fCu+jdaiPxp2CWn2ZJgc6qp0y8+33nfHvz9ZwP8ufsM7S
4VSW/UbXKhGPGUVA7YE4IwdFyL6Oq4Y7K+dilB/qNP7yBJG0XkhLqZe/UnHedtK9
K1Kywh49xjpkawpgyfdhM/sDgpFySB9EccpjBPyPRW4UCj+D6PV+RLOEosuhhdgG
BdheXt7p05yNJy3bwxaakW4S22kup6W95iAF9g/SivX8pD6bWmkD0gP0VnT2CmJ/
QGhPkuURwfe+SM+i3MXUvDh/ipTCOXSWq7k1Ir3KNFOqcjHcCg7pq4XhPgxvvU0y
0JDxeH+uuZX1DmTfdcgB74kbmz20RUHdHUsDQuGGSmxbR93Hu9zr45M24dqHN1LV
3E0PnLkieTWvHxJr3PjiqEPIsYArM0BQnRTeMdOnPAAo2XhsEXk5vyjRzrTrYwvN
iArzOSnEpZ5snSUdH3Us599fGa8U1YHwdyuG/3lHk2XBu1DRosKDPsWMLpAeaAeZ
nsY3NZhDZiTkOpUc4N6eCGdEjzmHR4n6bX3qzWF7/gz/g6vRjQYOuuRJWPtv2wK5
J5nkDFp7m0lkh3qxvqwx0w8H3R2iCuFaEtD/ph2N+tGygao/dRfU6rkpvCN9Eniv
rBeKa6sKRElmDepOwIkAAU6ECsWh5s8OXkKxDCeZR5k/S/YA5B4HqeLL+4+ibpA5
29fpYBpcEDJ/GpjqcH90nLCysk0XzPt63OI3uNG8wqCxOFqcYPvUC+x2tC21UjrP
NXSW1vAb8feLfeAhyla2drUEsC+qi0iQ04ZycsDLj2gN/pPQcaVRZATfwIZPYj+t
BYGcxj8DgH5s6Yf/qNEBOdpyKFZyoH92xGQDR93etNRoTenuM/TIk9SkCNkoBr+J
4leIAcjPMocqF7U/ld51Ao7aDcLC2SAnLac9IB4k+lvDv6iVMgxnTa8dd79GYqo2
wvPc3ANNXUJhHxnws4aFCUgOFqwvT+NZM/9MAxcY6NQQWIS1KrE37xZD+ff3yQpx
ePbgKEM1UngqMbyNhOc0c/AgUHL2X60qC4HuJ6jNXuwH2ooLWElpm01cJa0/6sQ5
/XtqD3yywGX4DC4Eq3WR4KeVEzm2VZ+kyrX1GQpwoBFEdbePiIwpKZlm0kFaWU2d
pRH7IaXODpMw+tYBXP4tD5pEOayljr5AxNBv2I74r9Abl8vnzJk3D1TQQLB1k6ch
35fi//AP0vq907ZVdk5Al8PAKB4AyjesOGlNuHhRxi/mk4k+YfeJ4Dscq0/V31j5
TA0UOVSa0jDWVK5ZQZ0d/qfJUCRKkes2EQnPUTCJFQk87mmXKMaNLhT5APWfBGCf
eJs8orU7s+Nc9diaHqieSHQa0XJ3HkX774QzgU4vGX1ZfRDYGcqR+ELvGaM1tA+U
nMuYzxY8Ax+on8Vp+vwFjyhGk3+hNWXfsMq9EIWkP+N96EE9S1uGSkKItKi8wC61
7F+Rq7wcSHcnxk/CKPqddSzeF8UCNJodd2mTHgNgGeRLFai0hbnvbtlkFfQ3JMol
30svi2vcHDV0bEOsY0qzY2wBBo5onbk12ivv2L2djPsQvnfAia/QehxIPI9LQjgb
+m+eb3ZTfX5V8p5ArOrZHlt+tYOKke6vfKDe293G246hyO+A/afCCDY29seLLq0d
0ZULxzQqq3Ar/1EYUvLAFrOQpJO6zNRV9go4Xp1hHJIw+hEDwbQFgt/jAeUY4+kp
4B51asHHMZLCMv3j/hmMdwsPmgR3vVfjzY7gwSCeuq7/55T2iVrU5RRfCGdeiH/R
ifkYED61cA8N4wEljskPTY6wOVQ6nRiHefyljkVsRw4R6YbzQDDhzt13GhBv1yTZ
K0r4NhYlfk7JjjMt4gFCI/vaHFAuUf7KCYl046pZd3VnfgpKRl2NPKh4l3KuzMjs
FoFlKWbcXUvnabjN3QSbeLi/dR071j0vNgPKwjYvT076wLAm4a5c1A13pkKuHbAx
rUFE4Smtgoz0PzcOzkXpbPr9gib2b3FSvD2t86xd/XCWBze4bzG7X3y3bWtYdDWQ
8ashfF2bC4DhRvPyFeknKljH7jpVCMfld0//uwHw7BJxEv0OimGd/AucmyJQbnjY
VwvEn+ZH6ouTXyXixP4D+WHFQki1iedN4qFsRKlGg1ie49z3aWFhVsJ4EX1sW5p0
i88sCqwsEjzp1v44PaTMYCjOBSsvemU7kY1ydo/FABIfOXlet1hehJ7TA6R6ImPB
MwT6yeWgTeL4+68aJ5lIheZ8GgW/6psUsZJvEQWWfdQ/n/wbys3PpwL45k0LsOWa
Zlc82VtI8hBQc6s3cpjpfqmRYc8ZvFnqm4X8i1IFXgaJyaBEDiF+xU8U6+dfZ1xQ
uFL9eNr3orKEDWuv5olf7erCOlcfIYWL1iOIMqcVJEnEKpPpYwc5l8wbBtY64KdU
E8qcmDOPdXt7B+wPEnh09lcOEEksvbBEBFLdUElP9opSQ3f3DR9Ox8HW2i5Oih+a
5zCeYOHcn95iq59QoVHWEsjUdGETWMNp0RtEcz4y5PlrYmAYUT/krIj/CcDag1HC
nOlpR/j8ACiH3Xkc4EXxoPX1RRF8rjqHlCaiONgDZr8UOkBy9k4SXxLcmlncPPEM
xqXU+ix5OEXABDJ4B+/RbaHVQ3h9xRRtXfuPMVi/b/J3R68sGAx6ei9S4ZhSWLqO
TtNMnFzR2Cxe6SiPU83v7ChC/7PUXsSS7ivJCSPTuILHCOc6SnxR6+Eh6XP0Kiqn
pQXCcUUKvMx+r7S3RKhtYg38cufgum9fs6n2N/yaM1J9wz0pEzX/jiU6dZBwdAcP
DpKGeIrUAeX6YGpwAqpNpMncj9aNqQ9AXJTVljGG7zF8ZtV4by98yOnvTdr3TIu5
3AMqI8cyfpaf+h07/mMnNbsvkrmG80N2PyBRuVGIBl4cTItOvDK0w/Nyy91v/4t5
eCpIOhPOrUri+shc7jJS19AzXpZ+Yce5x6Iojt2vw4P9DwA+ZFcqk9ayVspr/Bgz
YoNalOmmYuKJL8+OKkglo5h9ikjk3g1pPJw4T8odW8mU3IO1RldtmKKxwH0NRk5y
2OOOczPFS0eRrcc1u3caE7lb6Lh1wzcNLMwAhm1itLDIut3OjTutD7YNZIjrUrh0
IHVs834G0FsB958pifEBwJVXKijseEuDK99BkTeA5jJxFUDu71vH6rZc+uKd43jz
P72VbNbsU7neay/hbMEqNKt2ppdLK2ibMGJ5MrItHysxuuwi6k8+JFrQpR2tVPJY
PnlsSxoRonNWZWnLh6HbtEh47EuqI4YhDH3NuiYDg4E+dGbI002nJiHGKfthO9a+
/lVp7o4wEloSSu3ZzBIXeHwM5iZKCYpIObZA5e+RneALMnKjFBthErQ0XHkThaLZ
DNs5QiEiZ85W9JmV3g/y6dFwQm9hlIP08IiZefkQlHrpUYTEAKag+nS63zgEYyZN
PD490qCmvB/wKltXoLdoXXGq+lkSDi9a3gOaYZZDbu40LmqGLGctXOuRSoHrWylV
3sw1LqldnA66PPRZhLXNhzzeuq8YLNVHjywj6yDnZEiI636EnzNYJs+qpXpNKT+7
bmD00SJ3d+IfnFQ1fdDFJdPT9tsFJ32XrIoRHhdIEk4nOpDzQNddfhPnx4UVz28G
I7s2udNo8rkSyPdcXlmHe+tnGxOPosWDk9/tfTXsRgRN2DKaKvkyerQMznNWGTDs
WeqhhG8kBbMC37411m4Yrcxybj/restqOWh7Dhewzc85/VJGyGSILo5wF3fkZEZs
Ft9tFSf4II+RrO/QfkeESfV+aIymqPNNIXe39z6WYxHkPdkeb75E33r9Xu7PgdZX
DIqGHJv2vih3AqNypxHBfnaUspoMWwkZviND+hsIRqXnWXPEhSPkliF6MWmliq0G
RH7r/jtezLCojg4oCqR5+sFwAaI8N1cN/0V/A7y9lb1/BawkqCRCL5N4WnA1f3aO
ZxwC4Ov3WZuKKewN7vBy+RytDiKsflfgvIl+DFkD7f6g7GxiYpK5SUiLHPBBVhww
D2pLrRboaw+TkIB1Pv2loWiLUhnaGy6Fiu34ayphqxcByo+I8hm7LtoP3IW3eihE
c1ColtihLvm9dZTEDSlUfFAI+m+Bn636HtS/M0gIk5t0Pr914wHljZY4Cvsryh4U
nqbYuv/HV9W5mRFglJrEn8D5Q2nwUB6yJ/qRepRL1/DbiIe0ctx4CBU+0zP1M25l
8ItZdfCNQz/ds6zy6uVHhjt5VPS7ywDFimi2vQ3WMXVI1P/D8LRMLF8tSlTmf+rH
BuxOdh14R1D2eZ4C2AxbD61bVCRYjA3nYXkbop49TxVA2N/wDN7IbQJbz57SrZFQ
nOxiLUENyMXmBzHrTAMTGrpRM1p7/ZwM+1nIRmLnvdqIQ9VK6I+t3HeLYAkLlfhE
AUEJUhh/mpl/eHqw9C7glrrDw/8ixot80xOdlL1Cnngj0kcZCPANZGxVPEkxRQSq
OmyVBxh49vuyCjY9AkbyyfZm9E899kuI3F070kAmEpdYBOgPagFISE9PIMu9dlZC
mBv1USM/YnkC3jT0U24iWccmD9czm9nwQ8U80RJUGJNLYAV1vHM4JvaizQrm+jui
bJwhcGnU1MPoj/BZjp0c2bCVebFAJP3sxz11Tq29VjSZuJAQktEiJ6TIN9h+F2rk
vWq95XagK2i1OYI4ZgQOuDI6BNnE+G6Lx/tO+taIo5whlNnlamdIdJDdf9uUZG7d
uPZhWJtT/8N41ZQ/uYD3Mb3jWOSerofyuED3p236yOBHxBkW6dmqsQA4tReeQOHg
A+ckNO1RlL9KtlwLz0VjsvW2IpBj/RsB4v6C8FlB07+xtrbPJrchoq6belb1RMcX
lG9newdbLUcE3mxDB3jlvrUGvk2hIfY6BxuBkfFxDlYZ9ReDPtdhm1rjrZwS6DFS
aUyLrxvlxav6Okh5sDgxX6VxJSs5Dg6qzhnj0V54uIes4D54XjiSkFxcQyJ8RXeL
y0wx96CE8Vk1DDwRkAFdmkB/vQ5yeu7rWR0gDRqzU/GvZuZ/ZkxbwCCBfZXPbZRy
N+Jb4f7QDY9h3ScwcKyBBoYi+lRZAPHieCXSBxCCF62hP38Zm+c0YYCBrWh35hwP
FLfNIPGMM7AC+4cZ7BZyT72DK1yOcwOUYpOiFqWtRkWoEGj+QbZ+3JF0Kc/CWuHZ
JD0Ij6GzgZBKyfNrHO6Cr9ZF6EN5ChqqO6wDxzQaDMyXJxrff9mZ3JdfFasQagC+
c/wBgmSK5zR4ZRO7l7GEiS1o32J64HkuNxyjjn94IirPjf0oBbjR4EqAr7Mjrady
j5+y/DYhKhbrJG1vwg2Bzup/Ir4Y0VIP+CeX3nwGCy1of8Py6KaMLM6OhviKpoY0
BckoLRUIaVdZ7NyGmXiuZsjcR9rnof+2UiGExoVlYYlF8E8tKdQlGh9IstUaIsvx
t4y45hLOCLaoH7wUBd/4agXNX2mM0f1+El18PTkIL+kSFSJnEWlUJs3R+sEMiFgB
xXD5H9mbKA7PdzEXEBrfplqttshMVoltZjY7vcstPErUY7PiHKq/DPSmIOkA6wlP
yguy6qQoIKp9DrW7fosuqdamv9werRcRh0iwH2eKF+zak2uPjYlC0h9G/W1b3pcE
t66vhpbn/nXS+Z+nkpBF1t/xB5qpzsEHcTgEi0fryXA6C7jwqKIEn4AaWnmtBQKi
CbyYQVmEVN4FNwkpP9kvC2lQyu1mL0xklg1Gk1HdT2Ab/UWXiFdzaFNBMKXwcEX/
AaRXzEvDFg7AXBkD1Z+jPpB1+uEROEIsfBF/7G7EbBYureeijKHzYmt33qKaNEJs
m88QbzI5Oe/l9MkeOej7Ya2czhIJ5C41Wmyxqj06CjyMcSBdizKDoXyZX6/fZgXO
vAwpk/D0BK/50sdsziOc0tx+v5DIogQOHL4miinUq9+hh95D5VYi4QKHvmJ/YbBp
c/7eOeE1MrDWsppLoMw+O93FlxBxIc1Rgzz0+gRMDatLetr5ZEs+hjlXMFUxgOrL
zVKtcfQyt1YF9zQm5nezxtmVjWiF57Yy/vRSeN3iMmpT/BOFVNvZOjDw4O51h+Ys
ZujRaeNFNkb+QBuGU/r7JVmSXhDcIfrzoMpkp67CvRwCnzYFMlNrQHyN2ttxFaPH
X7g1AKg1aBT1UzCemfn88kvL/vR/N8wHhmD0bhANrKmquZl4ofzoJMQ1d8v9cxwl
UgCye6/9bWQ6iIZIaP3diwph2XrlOwVHJOTrXb9QRaEJ4a/PUgJk0D2KlRYit6jE
F3kUZH36aTfNJ9UpDzTqtLKCXok5UyzLsGV7SIGCXYr/UfFb8v7tjHrk2QzTvzNd
B3/0SXeDhGHI5A+UcbfvzCwGrdJGOwbWuyKjkLjoQXtpyqgq6IEXKhHR3AoIBgam
FADTQOFTpr1BT7cXZjsovYZOrb3eE2giJyGCEyaTueg17x/yG2dDkyYbttE2rBYL
vvpriyMrd3k97Dlg7g1KqzHKtIpyJfeTnCSY5x2mdOxXbw/MIeLL27ptQLHVZX/B
8ytkpD4NmGPznowW1oS5e2Bka9XGFr4/5Mcdq8eMNUpeOhfjLvLeP6XdfCLxPt2N
k0w8SvucfoQWyfAEXs6TD9dATVodM3GcKotLUHkps2UN8yPy6LesXoXdYLJ/1guD
WbEc3TtiIoOnTPKazgG3aC+03jwJOHZyxxW23XDopHbjnV0SWDfBqF7D4AVz5pBV
EalRkmAmopeOHk0J46x+a4NT7gM3BwUkCNyvFNsJUyI/Z4uy+vOQxVGShXnBUXFI
qusJbzQuhuA77EtoqsnTQm1rUqnemQcUzdzpLbPKTv1IezacCSOfucR8VrMrt8OX
2acG6JUspeyrWE7EeEmSzNSZvWpiEKyiLDc5mb54pC+Ib0xAtqsF0S+K12c3S4hP
fVB92v2Ezc4q9GDBXh1wY57ji9h2ao9qLxompDGMJsi5lSUjJl35udpf8lPhelcQ
RedpD6ccx7AfwkZD5sY2fmvhcyMNKbfe8on8nugLjP75ZgxWgLIgbWidqYnKCJ6y
jUBifYx746+T9jkXu++2DA5+5p0jlVGb4SYK1GTD39Md7SO5Mkg38IP93Z2KrZFo
rpfwDlTLKUEkG1oJuNsKR7Np0h8ITbKjnbKvxyz3KFM7IVhdASI9qYa+TyvPv9dX
BcGjqAvYRhoK3r8rCATciWb8c1qPu2Isxj3CSFfQ16yVtZFRLl+2aOmoBW4dj2Cq
Qw5vcXskxS5MERGlVg4Xy9iz+CIbUM1iUHp9fASjjg4cvlmLHixWu+BF20hWsi2U
vz+SUhysj51cwkychAX2MJn4AXUvlRSeVEt4C14gMeyfmC3iI3kzWHoVTdvRC+Cw
GcrNIRxFanhxUrrb1Wz3vUES+ZR9IIEE2wYyF8WKCXljOe9e+nBMsVpSsVfaP/4V
Yyc3wt/L4hpMl+3sVqeGLK5ejSRPrkvBqlJ+bjylv0mbPUC7HshkmUHDFBwwxUUy
7X53rdDf9X1SzgItJ7YMQcRo/RkLk9sk2V09Zy1/SYWjKAPdCa7et6DKwZtGxLO0
OXq3yBuBgNFEFQnzqZpnOwQ8p1LXpK3TbwNt4iKppL34+gmDMNjNuDgmpgHe45g7
Wj6m3Z3PvlPbw/fp1JrP0CKPxjNqD5oeb6Qrhw2e0f0dZmVyIfzxASLyy257MEKQ
TgVnPEbP+17uKGrfLt5e1o8tdPmwEOqvNQB33Vgn80K7KOv3rOL6fgIt+eAlWN1F
ff0N6xcyH6bZQ+iNAZ9g5+2XJpQMiXkx5s1Kfu7zQV8P519Epa5fxBCYkt2030VI
uCXmG4sbfZMGe7wLxmLSFkd/MSjFAll9MWKAuc9UHqEW+36WGGm5/a647h8EueI3
CqdIgYVDGlA4QL5xzKvulBUjP5fOm3XZKPxI4Eahvx2ITXgIkRp7v4V4xUlYjS6H
w8BkkOTWmDVbxHcx6Ew6xPP1NDIvzlgrnUGs6CyxL0mZCEWB32YHbCDfppHes42g
xq1m7AEY/9SwF16yp146dF7c8M/go80GikUvmDwIDSkBinIy5RQjYQfxVCXv+qjo
5P7///YNC2grr69gOee71VB3UltGlnU2dd6ISE8dI6ZmOhO5a0l77psDIR8PfRsW
Jcf1l0dUjV1CaTM7pnV3QASNPqFf1mkDePx8HYfpo4dQWySkf9+0J+et1tZCfz1N
DmHOmyFUWYel2l0xCe67D0G8tp/1TcqWEaryZE7YkdFAd4lfRYcz94wDb/UniUC8
7/pQ17Hc05prbwBt6qIntLPOKeCwBGOoVc14lT0jFNHmnljSl/cu6H0DuFdryBvZ
VUCdBUKtZtuim+WIa38QwvEGGkDVbqGo07UqKpMD8cSRB5vtEzKujrMZA56czb4f
MsOigerxsZde1zdE2aj3twPHT4Bf99lX0uI2Myr7K+6jvQDNUc+InTKsZJIiF5cr
haUWRj77e6I365pEJ3QsIDnQO/JskYjT+DeCveI/dGSxj4w5Ewja+DCi1p9ga3HD
vLID2gm9BT01Y+7NFIl1/9UtZ2UO9H+XUA3E06+RemV3jbDRQnGUyqhtdY0ZrrwS
DJ33zlr9x7Rh/B0Nna0OBtADwQxH1OMOJs7xeK7Cq7HQAHMzyGs6rmsN7N9AJ4Wa
Eg0s5wLg+Ua43DRyaP6kb1Y6Tr6ZwFwjD9uYKEXF+wRQDPL7uqefbJCJ4NwXW8+m
H38dP0WhlqyFstTf6efGeDN5NvXRFaRzxO+XuBzoJSGsUz2RZOcsSkJMA3+KerWa
c/vTxwMcmDEHvuY5ajBQfSul5o+Q0QaUp31BnGTH0teZLk/EjvXXDlCIpeKaGLt5
EtlNtoBXer66Kji7+jzJRoEhL+V6wydsfO5QE1CwewhDx/Nre88mJCQqYuIeLaf9
c4wt9xWayzBhFz9dt6IZFlZJRX+xSztYRWXB8l3IO0ZtOJ4rw/4S/qAvC4AQ06kM
ehhXx8yoCvxG5Xw+7Xpd6YJMT1KbYROtNNL4XAG35yV6S52nLHk6O2yUq6dsRmJn
9ojIQIzikTrLz0sCBSecbNoz8u/lqyYWgut/VvN+3hpS7EAjJME6+iy0NnsT+60a
QS4pYW0NSXn2+xRFVmqevIym4IsXMqyROXbBgiCmy811IzwoXvRPdRzr0q4Z5uB+
7oDr7TGTDKIAfokCHROENJaDLxZknX7iU9Y9Pn75BXb7rOKqo+RGnxcvExa9Iua3
Gfj0oy/UZhGuwrGfcbSVmUDMydQGWk9vLgFEH+G4spIT1c0Y11aURPLDocQq0GC9
Jq4k5PeA3/tg9fz7NNIbog/GfqAcmQA6Ho31ZifIPUXksS9KWCxPvYv9X2EFAKy7
ga3hwLlTQiJ4HAlPjFJg/F/4HryAMNpNoj+XCgN+qvZvD39dQJiD9/ouux7aPdpx
qnNyLS88gYR96E0TQp1y8GWIt9M0N6wtNapsoPJ035Ia21OGeIhQ0ZKok7x6/dif
w7FmJItCPrq1Un+9pXctUI5W1IDuF0az+bttm5gftM1+i1g3cA2oVBLs1ZNKea2j
AImPVvEh3nhJW34tKQeMzav+mN41jC3nlcW5H4EItTzc+0vYlpNYkWlrm0DNglqh
aAhekxH9VAnQUoSpm7g/Ml53wk82B/8vu/PpYR1Tvvtoc3c+sdNvQOVY20OIvywT
sYZdUITIrqbHTFq2zlkwUzY7d1fInyZNT+UmRwELNz/hUT9dUqgm5+vfQDgQhHP5
cV1CbZ4wAGWMpeR1nUpC597i/rYsVM44u1K66NyHM93ieim098CMSsW3sAqc2koN
kI69HbDTpvKDKVysueZYsyYXcWT03K8J05KUUdSdl+Is6Ww0N7Kp2RDIupnPpl/u
fmm2Zrwl2WxSkv7l+ZLMtdo7Z4ljQEBSK+lBKFxknQS3wNyrkDgMs8Q5p69jksVU
Y7LNP8P7C5srptRkUypVf7lE/zc+exKquzyAczee+f8dGdUbh5YuWgFGXi6OVqhx
7R3N5t8Z8mh1xjs+o9TrsduSeAH57LLQfki/8Bygl7qKPFhXfpdfMpiSmKD2flCv
9nCVzIxSD2X5wPCzbv2vTMmX3tvEKENTyNLwEXGyPJjrwSesm3aKhYEj/XDeEE9M
kkDsg620kyxO3X0lhwS9wnL2d2jX9aMdAUqN5a++URWfsRCPw+uouD/XHHgpE9jQ
Zlb3pJCCZHXYxuw52PazEM5EY+WSJKNk8RbVJjmxnFGHaIRHY86qr11CyQ95CHCu
mp7rFYtlb5Bkvq/fWq5FzwPUJn13FFYTdWBEwK7Pv1/Y2GYAAukqerD2Se/Sw72o
WpWcq9cwFWgn4UxJClg+t8wrtnz3PxySZSh+EIMyC8Ntx/3zsoZsqPcCwMD+5YpF
0/Cht6iBSXWi/1icFe7k4dTK/2YdiWGRmMJ1NXjmiaQdmITBByEJgcm0Vo/nusjT
G0WhD1bVSCw8gBx0KIZQfsCHA+eQ3rozSK/z++TDFE0H2t+S1/Ew00BsIUhyT0Fn
k2zIaEsHnehwpm/sgV80+DVe6ssOY7qF8p6Xi8p6jfRaAxSxGfWCzLZkT65Vi6jW
/JR4mzS8ga8c+yc1egRsubd+vODLi+H87Jusg7+Kljl/SNFsjFxKzYRD77EsyMfP
7LC7tiBWZVr2DT3w59nhJKaSoSPLlJueowLock14Yg8Ao4UVU7dOQImXJUBVhauX
ntYp8dPi3gBaOSrXs4dnIzLPtk4U6GB+uv6Fg8jkwS8CoavuwYRJctdiSM42tWNK
CUIYhsvXkR2ymqNrbgBFHvPWJzN3cq7jHlP9pnUAmglJF6xjSj0bL2gal/VHHRKT
y+v02voCBQuKhjJXOWVeNHSCaCtx2KxhDiY3gqGiJ/PO9EuBWt9NEAV1uAwdJUMJ
2dSsqX1oXU8wrERlSV+tPIeZPOELwGYVbEITeyHiEKA2wfcN8dM2H8b9cC2RiDbd
0vN4A8jU1xpT+a06+7s0wT9J7g388kohISeZ9zAes7DdeLt8V7I3ICuEJ8F2n0TW
1UXnzC/wI6gnxFcKggMT1+65mDDEv2Z4qttL7xGkPW/O0FY91mJz6cBC1cqcL3wu
zgoJCLaShN0MvdIP1RCV6EVl5nNHq8tPE4ZjcN4xWmzLy5fgcV2e2xLzyUEoaZ+F
kx41fnGpRTa+ml2QHImHuXOasNw7AD0MLN3c5n8VNzn60jkWbmLx2AJA26QugtiE
ni27ujpu/5yjhAG8W38+dzgoXyz1xlGw19lH0sKhVlpvp/orMmLx+c0BuY0QxRFh
Z1DqJYwaom4VuivSlgzUQNCkW5p3BQWCk+M46vvXphKE8Pwpwk+PDM7wfyOuXHGY
CDSI2Dlgcj8s1C9tSya8/oh8zLXAyb2GItdv2/g1l9Aii5GP9DqxewkbdJk4NoaY
yGaCHgPxyOiV2pVKgZGhrrvL3deLPNmFpnlr8EYa8QeVBqvZ/kF6v6wQm92W09t7
9GR9x3MTtZv/1o+Yp8K5or9Db+Kfu11haQLd4SvOrxE1pXO6v5ktBK3p98mJ4AhZ
7Cuj4T4IyrxB4byZIR0+ySfHxT3mhEVMZ1afRN3FAuqIGJ5WHVgNdxTp6i7sqJCc
vY1CEShcH9C8XEh9JoG0hA8ACcY1+rxLEYLogtznQe1zj86jSKnkExH4X/JcvfTx
PgVxxV+GVIr3+1+/Kr2DUxnknIHuvBIjWjaLvWuiNl9T1KhMnA/wZKW+m0zHCW/R
snNhhYcywtcKYcN/7RFSVVGuxalm3Uw5CN5QFFQDm1CFmKLpSliCvqL6zbsoN0Ax
nf+7Wo7oTAl3ztAxdYiAdJtJxQyW/0idMMWO/DJtl2Xp98i3E2tm8KwMh4qZMESh
4VWFYIF1dRKSNzBHteYaPaHOPOAMtjQVykuBiw04QThQt+P6Jf1PCExFPbVXOlI0
JKJSZdM0BpKkzd9u1ubIKidmG6hyMxPDhViC83RXO0WZZobjzPsXoyisxA/8zlwt
jdoU3kcuFWa6BUMfP8doDDOHy2UIetTZSlS5USmoxgDTlaxCcawGuNw0ab+wHkld
9ecMLQ9pdN2a6vXFtDiK0bfiWK7UCBALxJS0Ob4lf6QCgORmuG/+JQLo1xoM+QHG
XrjuyqxZmj9mzPlrLez62SsTuQVEnrHqWcrF/ZgChXD1MQ375YzBmD+bUMC0mys1
j17X/9vO9hMTddUj5N6yBSAgl+QS/2CpoatI3TvYf4MbIkAnxSA4dYXdY6DKN6ll
JjHjmHWWHQsaEOPplpa1mdW3970pwBBxbuHH/bSjcQEG8NjcjVnSwqliFXY8pWPe
5QbYdTdtOMcCryxA4uWe2n2zIvHFKk49T2y+2asfqN/OxJmByaLzluP3V5xL6Df2
6gGt7QKT3tOFvXNvuFzNXyPxhY7S4y7OAKHwobEeQ2G66VMstNnqH89kDfwoupnu
1m8weEdAFiCa0QI2K83LUdcDTH/ZJfdC7MzKyUoMh6SQL96O6E8+tiumb+UJi+rR
+4wKdKLhI33X3LaXJAJhDPzJWsWQ5gpXqwRtVDGEq/1SiBsvjkyNQwo+yhaXbCwh
NIlOHXWxVi0FkukbjsEf1alWFF2NEdAsLnFbUrkkI5Ko5HhVd75khv1Dg30lPB67
Z6mfz6paf8e/5bk9J1jKMmrH2bH9nSeCq/4SWeDhzqqUbIKGYCCAbj1iF8z1jjDH
eoO8KnPocxHcoXOc9wnuUUf7nRsYxLEE3VXp614Sl3HPWNSr7vU8kU1ZPTZeweKC
XHtOjaJBs3GzilQKcAtuLSgVbNGnYEjhV/hEgzCt3dtBNBOX+IQ5cIFnAgHpOzfa
sJ6DM7bj11wB5EsNl/Ov7iqi5yg79xlRv7b8DJU0H91NQL4hkTTdH6jNkAUe3t7y
m5OcJe2l9XPmS/nldCmfpiaVkeqZOAXj1sLsXf0YYryPr7zTILFwe+DAon7PwBjP
aeQkodjN8eyoOMW5k/R4eqkDFcXjZhPTLiabycQgS1jBZqRMZ50xr93MnHgkMvvM
8KENjld3uOT92U6Zhy0UYaEdd58BQxtb+QwKvumKY9QzzTE5UUiWcomzxghbSaRJ
SUJbcyGZDEnMWilFmNP+3So58CcIe8pAYyGLD/q8dq5q1pOWZg+QSs5Llv/vO+HZ
FrCIxyA6EbfxuirRPvfwphPqmBs3DP3QdIBLb20VRpSfWHBbZQ6TQqevyhfR6rXl
RBXjaUfWzrtXXXRp8TqsFoAD8/sE0i3BJ3thOghUxz4kFSmHziCnUTpp3ryqYZM0
JTvQarDLybZeHHfWd0Td7C3aaTDiwSU4f0XCMA1p439w+CJWdeYZ3ACFPgmNfZCG
Ozps3a6xohx0KkIuZA/lGQ0vVIXGqUtGkp+Sd1uX+10ZQQojoeBa0wX8IDgenshv
ghuhRLmMz/juGqfCyjhG6pS1Fx8CgKOQ5ZFf7CYMIrh2KgaLiahuxszws9LOXadN
Q/ldAQ487eLXWYVSeByvKhfb1xiXneFfMR3RWNq5bwWkH29AqbH2Uh5fplcHnNAP
SOw6gjDc9IE0fikzyzawxe5//Yw3BQQCaCfL5mh+GFc/moQ9hc1nCV4oEcLz+535
ImAeaURDrnKQWAI0Ui8LmJhWGubSronM8Ox727RHD9+Zc+r3fjH78DA3vhC9oW3t
cFghsZxyUCHUlCyrYR4A6fcGnfRC5NapZ8z/fN7BWe13sJDjiUKNboXO+6x56IHM
0viEpwUMMak1p88HVjm+qJ9Kl/yF2iDaoCJq+Y5MiMe/L94cBPJuXZK3/Y4SGGzF
xFaEryD/PnqvnE8WIFj1F1LoBsxYh2COaXzXktE39R26zuKXZkMJ4GXd6Cw1N7vA
/WRrLvywZi9gQv8krXfbROz9+bU1bC599ernrqOuvjweAbnqHUQRgZouieuERLuU
dn/GSXSTcT62Dvwu7pCAw+VtLmi+8XluVgSn5OXJS391JmMzPcIu84Id0p5JdRNJ
jdmgjS3FxhDNk3EtDDpNTPnEMJYvNRZFZ9oSVZH+hEjfV+aKxA9cEbEItwbS7MgE
6mxWJh9sbCVJzLlQnswiWKEabOQJicdonQmudXEG71F7ioMeRgPgv7+szNj2t2xm
DpWejfmElXzL7IO3xIj2WrpK3KqMrFmNPWA3Am3NHgpSSdHLtxQNSUJsi8gfi+YL
Bn9aiabaWnkAGOrZ2nLjh7IPkQh5Em+CaSiXMr1UsXx7vuGxG4RIyIbfBqg1XKhu
olCV/0kRuSMTkHRbzR5kw7VHFLm90u+49D3GKk7MdpdqcRcS0dDGk81Pw5XMCCLb
ddN0A8z7q+TCtnY28A63nQd5DQZIJPUPzj6h3EjR5M9KtochGMz3hC9FAiYsTtgx
poSgVqLcflZ09aTanseL4D8V/ijFmSAmfzpzJLYAiZ9sWCr99GdzgmSBMcMuJvNj
6UsiAQbUhurOxcO7Gk5B1lncCL1ct2SY6+WS/PGVtuGKMwaFHDETe945xUOw2tdz
ivUdxKWrEZmryMGmOYxVWDsMCQBtl3z9iWqtS2qt4imIOrDXEBzogHlDzsynA+W3
6r1V5JeQZrIlXXVHloCt3Uw+OXpJ7psNAeH4fnRL3LIN6+oeQZMcAWx309NzxQHT
d2WGxl1HNYb8yiaPjyAjw68j015mJY/kG7MwVw0u5dqeBMKV3P7lOieXCr48xnmT
4ZHOitv8B/OupEr1CY4vynGnRvuL17Vyvvs07Biexd3+khhlZGrpDxVxDUijbqCt
XeTS/2UvOaH4EXwvdFwwIp73nM7nuFynXtjzjjnuqsJuLngXVu/tJZc9SXFsEX+Q
sJhT6cvAsu1GSPqf4DLzO6+m0T59Oojf6VwazbIyTqTJkOmPIKbNzZPdSK/lf9mv
tMfczvfUcYWZxbIoQWzRdCk8krrnY2eBOp4JEmp6z3Y5BtEe3KpbAZx88LZVf2io
NvyPcAKi6pSyeoKQ+FS5BxbTeoE9gimZE+cBRcHK5LZTY0DTPnXZZYGRS7XxFSlV
Fo0R3t2gm2rOBaYQQ5hslPwg58cYlBmH0Qv02gCym3E85yIZUuZhClMc42br+U4O
++9sXYIRjKASOEOQgFaQwpOwl3KomwAWtDRaRsTIQYBuAi6l1KAylqoABlthVtcA
6oipKBpBPovUy/ryjUstfKvDoJrYxnFNjCcdhsArvoKm/4Z1DIuN5lhOE8Ya3I8s
ojZXPelV1YhldEVTXCH00ussglmvSxB6APLSlyjt5HZfUmPu3a77mnsBo3Hnhw9P
a5aA1Bwrb+myIbYWtacffJaRGtcRMr3keFsDCmcXJo1P4mPvL93YD3p6b6W+dyB+
pPgRNTMegaYyNywLa50zgoly5NgmIeHFCTbYvD1FQm8K6KovLeV+y1GjhSQAfvPC
GXjwz2Q5vWWI39a4sgWnJFfujftz2udENdm3eOZb2T01u/cD2m73z0rIrnsb8QR5
zcnbZGcRF2f5ivFf/EhCiD6FLTPYXLD/nLWfopF8rWYXtqjGwLMbfRRFxneFxqO8
uMqXStlMOw+B3oH/pkJkhS+aMZYUwlbS6lPBOjhyDzF9rLiu0PkYSxgrXLLSoeqq
/VuOMJ695zypIVTQ/yBr7cGRwZhlrQBj1m35X7ZpwKthJcyxEi+rnB714vG97bLl
EDIEFFfrtz+ivoGQi5dFQ3PGLnXy22WSKPn43oa5J0AwsXYqiOJXuWyDciGBDDVQ
/W1tb9PAb4KuCP8zTRnkfxIK9iQHVH+zCjm4kES80hTczFnegM8HaVmh7nsDrQeL
3hOHQIWEs1kSvc6wBk7PgZEzA45egEZ+yup1q3UjkxMcQRnAfXDZMp/FpV8KaWLo
ySg0d9lhqWcYsANRWt+pgwYgd/TeAvltYVPdJzU8zyhz5Q405cs+NbOKf8JytQv8
hgEIYJWGj/PIZwacu+AE3DyUzmp2vJrixRZWwMUkyQ2ULgszmLq1xHr2j4+swWxJ
G3ysqbcS2oLcxc2tMGkPGm16VDBcXy/OvyMxAy/AzzXJ7X6WhPwMzSMhZCAjVhBh
cv72e1gK0JjmKhwjLKnkjPfuA8/WEN7ibvutg1yl6wH5XZtwrbT0o/of3mfAfyV8
4wEZ6sr9Jg2N+qFKMauBHTvc6m6+OHDKNOV/RVRCVuaw03jq/LsakMH/yzEKReht
EbXfNdt99XrUa5j5NcsDta5IC63emGTK6zVhaXmdJ4YbdHDcXqQMdgDpJMhv1yom
1f61jR1xigRvSWRHPO7pseY+3x+7In19stIZr8KmMDz5yhGi4MZyTQvJ5YUVNBn7
+kz6EcB1ENsmt9MEDW0RG+L1VtEHbjiyVL677zJd4R40KfdgkKtgvT5G2Yf7docW
6w6h4aGG8ad2H7B2Gf/9Cvawpt5dp7SzP621D6DRzvTdpKlMyyGg+GibbUTRZCLZ
V2i1ydtnU0GYy3s+6CGVekkY+dwE6GJmknzWyPoe9do7w5wxyWMLGtF6j2ME1gpY
SGnseDAcZvJQCHNkqmxnoMqJiSd8wXVDmJvvyiLo280d4OEneH1NScLZYl5teBN3
yNrtjxL8MWFjJEyahu/OVgK3mybotycVBpAMZn6fov5HoF2lZQVmfRe9L83xoAXC
N0b2LosJiaC9RkDkUVs6uqYbVGqe1qYFGgQ/qQ/xAw62FYOGI79lSmLHVeFinjKA
ZNK/YNGA/I2QP1pw6GhiJCJStlGoqTpuJ6Qx2hdUNXI6b2W3eqAJjN9xNVOyOiBs
CP4tqM5YWfQsF207d2XnGD3PHcBGoyGejsvXe1owkfn7iABSxOaAhv42PFMn4Lc9
lZjX1Q0Bqv9m/d9XKM1ndLyi6KmpkT5ykBrMdhkGcvjtbMJdZhgFVefGfK/7ctS/
p77f0KpCoqpkNUpO1yVvsOBMrDcras+/CN6WpeOG3nc+KdRkPxgY/LxHhC/UxTXL
DnlVlrG7XyABkaFdZHxC5+xmKip3oAKeUHky2Q8xK2+pmkFvXRATHx3uTmeN3QWx
Qq6e+5twCTXjQATjxv8O7+LF3XLsBUOQPZ54UiaH5JyrnJV4LcNzze23PLB4CSoj
3P/6zznZAiFt/x5y6CmG9MAE3zuiTINw2oH6Vlq4G8z0dm39ob3Q8B9l1Ap6hq+p
qOUDF1xkDS6VoRyGURs/6f/2y4w2jsLfjdVxPs3g5/Gc4sjGB3csL6IjFftJCXQG
PTw7MFkmQIQ5XoaMEdJ55+s5uASAoeaO3WZ1ZmAANlb2lA2CmJLOobFb0OMf0jP3
Dp03aH0uOFqXcUvfY6j6+PWl2gVxeyLB8rGJJq1uZTjC4PDodAO88fpv8HmzlvmG
dKmuujt6aqwbOdbDOh9CKioUb9EuAJrqkCNV7FVKZylRBuOB9+PWqFBzoBpb6+4s
xiKKcQUk5OJ9tP6xf/SwY5J578lTOtop64+hpRRqbFZiz+WM8e7u2z9g0Q65hd6+
kRTOPPobyTQ8UTQbtA1gKpttES1Q7x+Lf/FGwUb4H6P8hP+X8+4ySrO7nxV1MImL
7uSAIstkVpmwpjM/ZiPk1wDnXZrq5O3CrSpX7ZHENu4PG+Jja8O65kNigIKzW1uH
pyz/srbx9D9WeuL2str8vvE0BLuD1H6XC+6A1+vLaO8CFNYTu+Bss8opXsO9HH9I
DtNZfmM+HV9tlEhOMFqybYVxDhiRcrLHD5tqHUjHxsCVsonZTlJVw9w/4s0gE0bE
d2WnZTSEMKgHwBfxDv5xW8xaBXfdb4JqAbbTzp4jMSGyVpHVPqIBreBQNHAjhD+F
cvR+dG1dE08YDq8/0KvjfznySVuoLgTWzeXXump27xaht4EmAOS+SoEnYr3FsU6N
m1M4cY4O+HIg9lmOZWjMLwd1IQacm0KEtKczHBBv93naLbyGllw59HnC/k41OVUB
MuM50PQIJgyZpdbEr6RgNMwb43/9uzrfMtEPl3bxsHEw8fcp8Te6BjZJEgcIB90L
PJl/GfKRmfWJtbt99pvyToAaujMKuI8hWB29fhCLZpQes326yhc1/t4CqtmELoV0
KuKG6OvKADTZSSLtbE0nkvGgaf9iD+cUhmS7in/g9Uc/jTWMd7lIR54W9Darv7Kl
fj27UK+SzDvmGCamIvq+S7Fh2NMwy6+hIGXwbOE+SF4+uyiQyGJQ7jNGjU4vNEZF
TjU34LAEOKiA6CeMaImx9pF81NoPQV9fQWaW/as+8U597w9foukwuZU17lcFHw6a
rK9Ep59rH9e2kpQJAD9BSqCT2imODBgWL8If8h5pM9n15FFA838b1byjg3wrLesm
q63HurP8EwMmcpx5ifl6GVaIB6gNpiKnJutz0jxXcI/c7VNl5RGd4pkqmtdO8txL
4pPZBt4erUtk7nLnDQIhjuY6CESUc2esc31O/O7CDayyNUEhS7z+yMEqq8WOma6k
Looy0YzqODgfw30aNNZEgCYhoSIoOyhLLycFVRNCOzGV+qZHvYFOn8gVvo4ULiAC
83E+sitpVtRZGBkJsQ+XM3T2nB1nWrcOph8XKFyBiuPc1/oPHYeztcjH440kBxW6
CCtSN/6vBf0iArsYZOLMhSpLlsAgLRs27cNBFoFRN12P9QjpfS236autbj9Jui5p
LOGnaXF6IwlPPJP5kRJJGOFK9Z/rr5QP4uCVHRrIm3PWckY9B5Rqcimxccb6RJOX
KO07cCoJ5HMbXdmZ9r63s/cWXfwWdjpb2XUSbUTwLsvVIkKDgF7oFdcpoeFK4f5k
DwYgWCzFSee5OKBAUIW0L4MTKTzpu/qKnD91yHpmV8V5c+p7WXAOqGDqdm5ikDP7
1lhauIYOtUrwgb0I0zmO6IXgpJ2lSGrZGaQ8iL9GMOmjLMUXW8zsjVitZnP6uHrX
JRPkl2Xhj2A5erHZh5hHuobComy/rmrrswTnclKyHbh+2DUWZl7rSbb4XrcGOopx
SQRLBPvY3ZdfRmFnAQg2bNBqSmK734Hg7HpuF9uS+vFGQXqXEe7SdRTz5Zpym7Q+
AmmxMEkHbL+hEQ7I5hfuLdX7DEvuHtxCD8WRZ8BkXeKZ1+Juqj4pGaJIkKSlWRFb
BJIffAG/f6iJ0BtPpHiFST38VHqnrqpo3Mr3aaiI3D7tvjQZqNXiXgttOeP1yZdL
P9eF5MGfa9KlKiA+KvaYq9oN1iQgvH+NyPbV97/GZVtSoCtu1bUjAtelNayvtKFd
9X5iOiFZXc8GL0jOV0arTWLnP1pPKHe7TJFs5AMLQ2IaGptsMBnA0FlAEcfXXXc8
BBWHP9fCVXKxp2gO3SBok4dEoHw/e/ISWyCq9Tu3ADJAAsqrPOFYrAbyyq+aZpQD
+/Nh8iUQlKAwvrMdZ6fs3sUnaPO/qoHU66RE9OjlqguViy7rIyWdrOVsdlvquwFK
DDwuwWpKAvMWxPiA5LHOxvlFxuOIcdVbjHcZ/6awAsv8nR2y8PUJm5v0J7/crl+r
lkDUdc0eKRl2o+uaC8799RrqnXPpO96RasH/gpyRag81BhcijT7899TZtqKE4ixe
70kG6MGZFVGj/uBhP+g5vBt07yFTeFK7+G8TZoMLX5wJ+mr3AjZuFVImCJ+XDl21
PhCKzbwyTxEPji9vys2kMeiBTqxsBAD7rs1Z885DorAQWFR/tFVUty3OFWoV/uwL
VPsO7WLPwR879NfjwHLOsvk3yeBCwXx+cYQTfSF5RIQi9oyn5ti9oAG5c7zkV5x2
CTrQfSDv4fLb0Tc8DJb0Oziz+Y6DYYAlTW34omVZItI9LONwEkvdx8BVfUxfXtqX
194U2TawJwgDuJEW5/RoGZnOtkvKnVmHgqOYwVEg1GVg2kgQ288OZpPpQtFJPMvs
UOFoT3VvjXM6tIpZhEjXpwRNdAw3GrI0xyzVjSYGB7qv2a/ClJ3KMgHAUHRIsDVd
QXIxHw3xrjoMa+lvag0lGrkrizqi5KR3TPEFgnK4me2LFijewLrPsmxanVr8aIUZ
Fo6J3dg+gV0hEI05VRpSU1ys/WbCRMEUc3MtGu3Oioi4P8viKNZYk2JFSdCqCmZ+
oZk25LoqWNqPLTjcdbD7KIWhG2cc3QZSSwferhCjqXcvQK8wNXsg+Ssnki6VQU8m
5+4BcWfAhb9QXxbdP2I2RlR9zGbDjeVrlETdj7zxsX0w9nz9aPbm7UpCD/VCBCxP
niWfWdprUc0CKwYJafjgLV2001d4em2vTFBAzyOSOtXEI7Wx6Hb4pcjeg8IMZxAL
KxayXib6a2J90qW/lIL9qjwmnSBT4DYCMUFFF/4tQiVrXtWqPRiw4ta1wSnd6BuA
EAfi6s6DCCGCk0b9Z+bJW9d0ACp4CHxS7X/0gjdlxsYYg5BgR4WFpTGRgxPX1jVR
TQJQHWxMOvvZ9x5Tsu73zIGIGftdo3NJfEE0woTfhL0jS+4zHYEkOo6X3cDYF53j
w+1+FUczuiict6mU0TyBF6eOBed0VrPY5JQ0H9cSKkdCEvjTsgpN+/ycrcXJ4jtI
9wjhFS1udJ8dhtcD9CltHz151ZwUExSGkethEjiz1LkG0PillWz+IviIjJrSELtY
c+9CE++8UW5Yv6xDYLJEoHUMar161jtnLbBTLNp/SCkfBqpih5wa/axADRVOLQtw
iDGA61QAmZobs4EXkJLzcCe1aAAmZGL8ibaP2rb/eAEcgso3f0OBTSdQjLYrm3CQ
oIOnRbqiYZ+t+rMAeEokQiikhVnMSgHlMlJr+PIelQMUQJRf2ClVZZPohBfSI3jg
Yzt5P3spuXkgYM9MfMAtnJxrbuaRBlko29BiHlh/lncLSjNlAup2CAwWTTTi/Hjb
Y3F8/H+Es3D3EfT/So01JUnDzEKmRymvBcUHGsLSjNavz8L3JUYGzYhAJW66KcK9
yG4GYu9U25ll6SIvBBDlvzHDOq57pNVz8agfYnUKm40z9CsWRXw8e5eFVlVMa9ve
48tXdw9mFZpkbQGidEkWyc5pM8KWk4cRf0PQP6JS8V7vgYtMXj6UQvrwT8MAc+k7
2Vu9U6JeAvr+yOTQXaLvhPHUxr/XRFWqLnnsutY4S/LRfxk2WWGIKQPwtmF7EvQI
9VcHG8CQMiTieUnZhAXEyWLlRc25kSIwzZ6UJO3ofoCXshj0PsCyYTlZNg0nazCx
/R/EEjX1nbweyk+W7mN2G4yp3W5tWFmrUTBJLKLf/67mABpI29rjF+Bs9F/e8993
FCgst/1m78YdrWEVCtUHTssQS5Pj5ZUN2mo097ul2X8ezLBX47KxHxH9tgtRH14M
pbCWLpBCSeQyx1Jn98WB9kf+/tj19+bhbrkmKl0jJ15uKBQadaghyMc5X74iYx/v
qp1F/CtuXRqFSSpieHTMIb+yLvmVnNcphX3qelxxadOniuSQ5sqcQTaQ9QnqsqoL
pzAoCLa/R5mSupDjNxngbeBsV8SRSs+nlib4kbtqNxCJWI5EgNVDsQrXevCcZ4W9
7uz1NzLXYn+tMDlg+/6rFbR9uHCM/0Xz5DeYAo7FXzjQ+qfoooGenVTZDty7YkPi
rewRLlvYu+OQFlnKeM97zvhXM/74kSfJGGynIL4YegMoj5c/BiTi4Z+pu6D/nhgH
ITNdkvfvJYDUr41JyyJ93ucEJ4y3MmuekQ09e+OU0eqS8/vUQ52FJYOAYXS4l2SC
6ON9DhjNoJlcXfsyGoA4SWK92v1xxXUujhHKrsAllWfibcm8Ax6qvohDWO23XLI/
Udg5bex9a8b0uaaCJxIM9e+02peBFWbha57YSRXjaY9wYl2qTJRftRDd4zrdzngb
A/QXacLD3YPvllqmMzcHwVUwyVy4qEj5X2qCJUmZXK14JXwJquh0pV/hqq2M7acX
/hXS4n6qj0JWIgeV+M/AL/byX29s/XDqwQJBZVeV31SnCTZK5hE3Zj6IYlA9i6aM
WzJd2F2RoQOzGfyLEmTkbKaLzs//iCmL7S9JXddYFGP+wMQA0botDchBtSpoEIBX
aKfWNvHi39W/+gRoZvUrfnMx5tx87VapLwdYYjRfDAcXNI06tgKzQOrIcdYlVoQW
m28VRyUJ8o/V5GsGG5BoAq1aRd7iP6oRr6BRE848VrMiiu5ebSZ2CokhVn7KRZIX
2a6Y1Ulw7sfmZPWuytdwLWZBDGKko17wZopKTZFTImph5x2XGIVW6ILEwmEpPZYX
ALt5ODrh+Hs++SYDivV2Z4mcnh8QL4yrwVtO47OXSa4/AKqgC91cJr1Idk8scYhR
MgyLM8U9qxviZkUAevEFpQdU1vSawJPmGo0r7WYUqgd8QKjyD4QyBzGXRElC+xTZ
SB5vxhJYOjeW/01cUiuIHEgBR7NVWtEnrwXWy+HoelNkjCIXkfqJas76Z5JlTmTS
zCpe6ErUNZkYSLrY2F6cjnKjcKXdDhU4eIe/APwD2VQ7yMk1SZtgwOCYbCsYJNZ5
X5q2oz7Ez0V2q0JCI93jCOwXI/rvfrv/2+PFzzIsdielPbWjFdDN47Uh3ZMX1zse
TMMOBmTWwL6pxVmjv6t52BobokvZ6FeG0nw28gc7EFvA8jGBuDIKpxUI0C05bNFY
A2yyr0d3wEdbq/0Q5AdIXyJvC9N0dFNzeH8sQ2Q0xAGJ6yVzc4pgEQO4gENZ7mwj
NJUMQoz8Chiqt0NXlrmARgRn24FKPP4TnH8pjRV4+kPlyo8NrQGLmFsXSZzH1+UQ
C5uuy7XeIkQY7hYFfs4paovmP4xK9SW1Wal9ZwYdqubZICYLwtKP9tfToyJrRPpq
4fMcsdzgAyeoI5u+haZg8/1mJctffzBrvktb83A86X5foMCZO48k05LiObuuje0p
cMBzFajH3bKsJNSLPg9qJHpHGCXlF4z1gF5gxI8vc7HTGq9zPdaDE53LkdY8u+Gx
/10/IEKCorXd3t12myUpSBYhk+87bIFicGKmevzyCpRivtorgZGnE6IArK0wCp2l
iBfyybudZ6rpC1gzORhbD2luLTzlkUezv9HUyuROI3bXmRAdZMmeX+YxwWJcc195
jl4La97V9f58TK0vux4EBiRwZ8w2mstPUoNWns+bLfoB2HyCEAoXVQnTeeoh1zBf
G8DDiqMV+tUg7ms2QJkRV1sriyEBoGLXf8jFO8GMl4ut6oRWqqPSVkQYHcgncg8G
3fXk77RVN6Fva2fF1BcCBIQz+CIDgk9ZGO98PKuZwvGSAz6rCglzrOD3ivCAk3mh
w/z5TLo+Xm9cuxFhFaW/xMyLAxytpbTvAeicH7nBBpZzm2olsFR94TWKT1OSdnME
aAUru7wBBSlVZ5TNSgCIKcQy1gaSG4Zk6N+R0Q8czwwX4alKv+tcCkFStgqYxeBg
BEZ5Amr/4t3WCwNpjZFwxQoZqGJdabg0JoSnQBmw1bew5CzQj+vkn9IqTXCsNniT
JaWljsVk4uic1iccbkrE7do5YvagEJZ4xyJOCBqKZb/fyMHKdOd+NR4aI9iUTJYY
ofyrmIQ1qEsmNFjd7NlikNcL0EkESbgPlT7TdHIl6b2Qmz9WfZsSBDqvfsHGbC11
TxyuMKe1TvnV3+Z56ojEeKvNZ/gAMnx97ntI+P8ysKtf6nOTcK0zxnjGO6nkmlMU
etqcUw9IDAF1X7Oyk4QIqTHSNK0owaUVY2zczaNtLwbX3uQGzGV5yEd2gbzCBOrH
vQu/QrKP0k+OsMKbDmKkhXKAg0Z6Sg6oqBBB6OAka2rtaTm5MYK8OcDDZgMkKqO1
frtD4bMYkrmTB/r3OhCfEdldfE/Sgt+oj9X56INMrrgECsBShYu5fgQdOra8Gl2T
4Qgofbz2tRV537hFwa1Db6PEuHSDDr83IlVC4J8Hn7vZvgVM1hpoGHNwLAkpIX9k
yHHT5KiRuLy41I1OZZZmaChSMpYyk1ZMvZAX2e4/V9+F2LQhpW20/SaKwBlQjyPv
x86/bJPrM1vbqJRABx1fyzxN0lihnIf2dFWes+bJTVSGchVRxm53NdaLkOkCjyQD
KODiqYVaAridcdQ8eNXolnwkvcqvRwsDriBmg5DnsILMTMys4JI7xyXgZfxXhV6T
88EUPlnVKU+9xDDI09UYAjGhsRaxE6NCf8Rry218R0vu9rda2QZNVVGAXxNoTVP+
W1+cyG0HhmogvAW3UG5qOsAOBRCym6jL2+7CPKZbQLhKcIEfVp37TSN64shiXQ/j
Jzigk96GcW6e6/y4lhbR3xnqGnU6x/koz0czKyUwwRxHBagl2GnLfQ7ZA7cpi95r
gO3kwH8YWippOcMOLGRP/u3580VB3U4bkxFvtV1OdLGvebiTRV8aZlLIX9wns8wU
lnwt+Y7v1KLhY5mlc1RLjHfPapNKYienVveKx7RkGhaj7xpDKeWNruyhFt1hsAxi
btTwVm1NuWRLESLJOzjOBkkrcIloojt6r0zs/53PnGaz+xjVYjwz/ebkgjK3DDIM
FZ7UBCDoA4b/WkXkziJKo7J7GjP5i9jooGkUF25pYTYuFn4mazvaToOy95sLJLYC
0mtNsi0XeZiVr8gZsYqfaNXS548NGkVx6b2Uj2zEBGuxmiZWuoMCTq4WSBzUvAwc
ezpOVBOiHTxwL5YjLxCpWEOTzwZWzam2W0w5sAzwRXmI7AujYpG63GVO8aaIA6ns
w2lUPyn2a++NrCve7wQbieRj+qBt3uX+jpnLYuH9GD1SRneVN730T5HpU/te5TRP
kq3dFY4JfrEDa70zTeO6gNf9+zsJo/5tudC6hW1El9oUIC7TT/LBGXKoPr7Amcam
aVj6ZIJk7Z+g/n2chda2UunVznzYA50pUVcctT1ovg3TYA47OyxhBfC/RvY8n2Lj
KipjTOITQIrod6PNANMo95XjpddWNT5df64/Bz8wsMYzqNxe5yE5IaDDZKrYq4m2
55ICF7ZMneg3pm2/JE7j03WQnEbqW28dGJ6GgDDaCa/MBjLL5c3mKkgduzT6L4nt
yhR+1SjRTo5tZCsbI5cFuS8WEZTOFCJguIPLoIuV0tRJjWlw1hYnbx8lyjUefgv7
NVTPW83VZu03xfJjc672FjBqnCmsIzFjPv7HVe7jgm38pGaWAKGU26I0IL6Zbeg+
et3q+M+6ab2dl50PdN+SKSyRgijeETB80ulLCwO/AsG9aPAQMaK7KIhIuHm2QlQA
WS9wbKVTUnVFelB85+mgAbLzzOz84vILt38+suC0uBnrjGysRZA6EBStQ6Y6VBjV
oZU+tiIvWfFmnDtQm5gE5iFW+4cYOYz/yFt3kAkfdl24FBtRYtSQzpM7fLHOJ4Av
6RiUbJ+iYHfR3CUoGDIvqRhTjrKdASTK3ZoxCRuxp1PAdeKUw+MN8Az0KeZ4V7fD
QT7dPOTQkmsYUBsX2TI6Apl+Pz9ElLCFlwBmURQmpUXBE38MlUaLruAcR9SabpsB
6MRRSM8hDgXCUg80UcbYyUot9hXz07uWYu7Z5srbancveoPB9L0K4piAPVIZlXXE
1Sr9cO5g3m64rUvsDoE+mHxBOts5S8hrf+0khqpJk0RWFMzf8Npun7ahku4jcL0z
IXQDUOMpTxEV5fQLtb+bBpuI1E+kDcfCb5C/MnScrV8HNDxAkNOfX6A2bIEFJX32
hmLygWSGwF1v3d6dKYe1X+GjxT0wBk9rjFu2S7kQg7JkJ1XrngG0Y3fbUADWCow4
PTddSxtskSPbktE6nwCYqUYEY1jmZDa9Zkrp2ppz9NzWY+epsinMRO0ggDNnCV1p
KzS19CNK2HMnVQx4CVCZDyvmZK4nBvCHACnw/SY/rmcMiDiHccZ1TS/pSDegJXB4
GuaLycJm/7k5TByiM9565htbtG2prAJvHN30qoelhHyot7BotLRDR1yyVBl8r1+L
V865W0+fddJCRYPXPB7NgrgZsoTvLivzGL6fZeH2I32zAUj3v5hVwQE+bG91vwnE
A/9MemjtimOZkJzo0+XVnh5070cF/eknOKdaWJjPjPFcBWZmZJnaPSJYTEbFkwy0
gHr7N0gIiz8PdlNmO5+uwdJkFnzTU4pt8G3hjToOx8jSUWQKyHUCyqzKV0aZfBmg
zEQeTD6J41kgQSPRHkXzrlPD51m5kpicgGdpYkVLVJfJLaGXb0bXoUvPIcAvrbLg
kLVHA1aCQaLNFvZefy8Ci/nXff7nifn1rn0xI0t1VrP4Hx1gHLpB0g1BsE0eWeYw
fkOVMETRDzP4HxPy1OkWAj6uYx7ujdzLq3VduPGZbX0UwsW5L9PalpjhtQH5zugi
wHqnfGpYothHS6+y/8L6p6UytoxyX2PDWAs+GKZtctg4KRGNycB24x1qtfnpi8A9
+R+0Hy4iHZDEbB9GGgZ7p8SX6xhyabID6Qf6rRJhluME8gxR8Dt1dPzUjXj0AMHM
wALSi7a/iizHJkILi7ixafoIj+XX2AotUOMQE8IyeMraOc/h2AhbBerQg6ydA5BU
+frot8M8+cZ2t46Iaol8YyUjHXbWctrkxZoqFCzfbq7pBi6wmJaRqf+9CeVKB3y7
flgARrV5sDMZ2YcYkNg0h+8pfJ4dqoUqkFvhTPReN8k6omfcqwJ1e5ywCdvyegzl
DrmSQPO0JmzIG+YgF3WKBTHvUtUNPpWtrzHTw2eR/RDC1cqqzvY9cOl3BvVRVjnz
+kpgtbcWcQ2jD6G5l5caMDQ+G19kkzLVrnI62Iyo+rOuFwrTeDutYiM+rnxgXNfU
8JJWxsma+3xEuMbGmmXyZAslvEmDm3Ko1xhQfopVqVgR/4nL8c/87O9AUE+4ns0t
FP/mjCK3XSIot71HlTb8u00MAllAVWdT9nWHio8Jc7glwAGKqUO0bFHl6T4lfPe2
NIKU7M2oKdejbsPnLWoG2SJXY9fOCqMxpUPdYDBa4lKCXk/FUUU9oMpdc+/n+mxy
mfc4WLJKvUA5Jr8j3GRkVrlADIRzFrB6vZKt2hyIggPf7WgnC6J6Cm9k62s0rtzB
6IalZuSIXtx7jxr+39Onsa1uAl7lgRNmwwN7EcjlJyxj+ns3GAulDT2483Oe8dYX
5E+a9sYEzayXM1KKnvh5v6qtZIlFmECBfl2Rbs4rCgQciCVdUbVZBzBjk4sPWyuN
OHZYgT5YDalFpwvAfkrzyxU05C7TyddlT0Hyx9oOmdpY4JiB34g7mPaWXpdxfMPM
rJzXnDa3nsw8sIonfBMcDz+6mC1cjaRc/4ddmPmffckEjoDqU+9iSVRbJrRfU1o7
JZzNFuPaHCcxyseSRzGUQmaG6wlAyomR+1ziFykJQPWTzlWEFz4q/QkcFkEbdniS
oiAWQHAmsigxf4wmctEJVs/Av82jyCS12T6cmf/atqpoysjCDasHpRXE9xkDVvwH
SGt0ufHead3vb+bKbDlr1r6I0P1Grtu7SCZtvzvZSR9tw52LJNNRIBrI8fXbDguB
U22nKSN38d9DBcRyQpdjPMLvrCtxfirQd3AIhatRvY5WDgZDKclI1IMOUJH8PIY7
GXnw+93nytiHLZpm1QRk4aUOv9gHWZrs9IRUGlkqJcMzHp7TOLLib1O2v4gG7arj
/4dO6usDraOv/XfAmcwqLaGbGdH0TIiSbxdWNufBoKhuuVnwBC/+ryJg/MsMuV8X
xjgbfM2ApRqnTt12kzyGIQDhjPGo0AKjODsW4qn6tduAry9b9M8htyEdhCIbAr4k
z7Tx+Ca2Em0+yLBZC6KDfA1YOsu5da7Gd9Ubsxg5EIe7yknM1/+Uq1bfXSyPVLQY
ZYo1wXjGhOz5i6LIrg5ib8D8Vd35nXSu/GsIRhuNWvdZgkEOZUcrjpZv5RO7jIA1
vn3FWRIiOGjmKhcNachfXZLQjanokgMjJtKPM+78/35NPWT42WJeUgxnyjl96X3J
C1UwWibXvENUiO+i+JaDYheTb2B3u9jJ4W17+GgR8emeX1vuJwJcpj1TunqPLob5
Y5TzAIrPCyxymL7DhPpFtXtKyykWUoM42tPyzHLoA7yA4P+HKK8AHWOFU9FlWefG
yk/Yd5cirawq6mdmr3RnS6KOBYip1OG+sZgNOc1Tqb+4ADJZdgy+st/bWIjfxLFR
SO7+wBI2r9zqSmGYTq3xgszregWqeirJyoa06/6RfOdVAlXEB0qigjGerxLO9ZvO
eQfE9GzHJPOWZtVFgNxIJGVgJRt5g90PcA8s1RHDRqnLqME3iG2skRiRH2zJ57E9
1WbyAPJbtw43CC1YlYM6boiZCf91kS6nMUoRz1Zp9e+Z73m56FwHAN7OQD9bu2XV
2NQWRERcUOLqKpUceVOftpcWE6nXsVtRU8FJN/Uywb3bTRGdlHbCnwFhnRNnCDRg
uQBUp94k34nOsjpJzFEXAxthWF/9HJ4Tw7UborvAMMsoKBl+vsnwZZXSAgy92TnP
gx0WmxuCoTihF3LNFHyZnIQv+bvk1y+/aE0DktXexISWtvXbfVEF/zbGMgi6+y/J
o70LvQXjlfYtMzeA8Y6xQMlXpcQB+4uEjdlR5aluCONOp199uz7MCzFZ+zXOUm+y
vjRhk97QrYdFMmSPjYtENw/nYlzEZNYPBU5yrboaRobAAVNBaOaqAVHpO8/SnWeq
ncS288qYgrU8rfRHrkFL6mZpQmocPNWFC9F3kmefwEDoqkQuzLsBfbhgn2iwFlLN
MA0aHBRZGKsiDsTJglwh16QV+oHtDGtoWTBrEevk4DovHb51R+OLenuAZAjWsj8b
ArQ5CKFtzQ6AwapXmcV1JZR+LlT6cEapP3AdB+4S6pMv7S5UilfC+Ew0GgSjEfiy
7VpaDADqTlnz9Z98eHYZ+fLC7us22AhygNdF4Z/qb8Z7buD8vxLapCBUDx6d37hD
5Lu2PAj11K7XAnQQqZqy/Dzj6gMMrJF0d1/DauM7/cFuR9uhaRbpFG3BKP1IzLyh
7kF+3JhL8wTsQaifJIG/23UlU6OQy5YDEDVY6q4LXyU4gaY1YmZNzG4adAcYF9QX
axwVcjyM3MPigsj9xa+5xUm9iD2X95f90GvUhHsOMvejuHLsdYn4JpQ9D/wk3Ieq
lqOhOZkTDThZCCqYOESKvTLkE4pcqOfk81l1lgxrbC3GksZjBoMKunNT6GMK61Pd
9Hvh1XVz3WhrvQHaBeHMLfPkQriw+HXn6hdsWYc2UgFFcU9Gehrdwd13cPcVb7jY
xHyHF1O/EzsDIkP2BBeTlT9MhQJ597trLcV966cYAY7qIcdmNHMYKdw9hgxbfZZj
BL3hnzxfFnrXmO3Ylg55IvG9kWjqFWitBWhicsH4hI8TbUFkCdAkVt0zriVcQWDO
WJTvraAmFQ7GFdnNMnVraDC0Zf2R1wRA9r9QXV1/XjeZsGWfjdPPOCento0S58pA
WByUdIykm7bBTc2LUFmBUjdyYmm0tPEz6Pao7EGov+Lvbatl1wyKLluBeVwFLV7X
NV5gjCdR/Kbv1naOHSz4aWc9Wj4ylKtzpwQ0pBRTT8xc8kO6cZ36VQyfahkpQv3S
Jl4Rsqo9VRPFoK2bJfJ3q2CQf7ia1GW9e/3G/J3xFjEmkk8ZwIq6w0yCRn27NaJ5
cK0zhHMJ2Xb5y8B0s/il70p1x6c0pFtuJ6PZQH3a8/sm/0tjoEiRuOjpg/Te7sry
NEvNYrfh5fVu9Z+JSgqynWkKYmQ1UBrT1qqjRQK0Xl6v7WxIlTi3V06a/eGAdBTT
jrrQHKtfPu6X8//QNHi6pGSpBMHMIFe+VOrKH+sZLIqObfmDI7Wm6DXbE9IypcxB
hLfeHHfHL2NSaQrOgpbWEfViz/RTNFF7s/qbfVRUzRP86VvjDfrSj1Z1hn69Lywg
cVhJjdARZFc+6kw1+mOcK5BYtthbrcTzZugn2W8mxuxC9FX1+O5V42EqOe7jQlri
58c8aj5nFO5aDQR5XHH2ysAnNNKl2BNiEJslflcDB4YNNNMseyitXbuU/pXEJ45G
croKraRVUy9v9SJL+mpaUI4zwWifa0HMmAenMw9QFTP+ViF+jPwOZbFFqtJAyxSo
5+n/HmXB2Ce9sdKIgD/MBA9r3K71x+qwr0CKMnR6/WUBWg2YV6YfrMnJ9pgpkR+2
piheyGtSYe2LhDcHfPzQ8FfSd6M/h0kp8vxnL8DXTQKb7PN1sp/iMnEPcK2clZDi
13Urq1+jRZ1PNQ2kCnmdYZ7bz7pwjUUM5km/BaCx3enKjbC0wQJm7TxnfNBsd1DG
oxRK0FtmPU5pbjNKlwr2qc1GyRB8jkHhMMJaL9Pcq7nPigu3C0R9361IBAFB2mG0
Qmc970lPgLGW61FVALW+7CToc9fiVjDXOXUwUNBGJ2v2uL45UqlPGQGJ0UL4wsHg
llIAHNZ/Oir/XGS9g+mJIU3DGGBfe2QwmvHgxbttWOIN30KTP6nNhZE4TbUdF+xr
tLieGikF5UCdFvmtyOJKuyDsT2hRGtJNw2yuqDMODk9p3duJpNP5dqBi7Fi4ao5w
MDSwlaTxvrM9Gelrf955FuBWQjmVEh0whClt1tQ0sjNkUpXKFEuDpBdj4AFM24da
Jkx3FVafnR6sVo8MFZtOlY4MedZHf/stZ0/9B+fc9icv7RaDMnVrN/Eu0ZpKRAAu
1VhuOAqKymuNGIf10OeHTASU/ZUtZuXBDExQOR/QjkhrdDKPGNf1UuP1UEF/KUZ7
LMINPW2oEOTYKqqy6gWy1BYdj0eIGFX+daJRjNEmzfO1lWzGnwR+fWbsTwHv3J38
C5Y98h+UTkVv519qrMVe+8mBWi95DSQs+c0rUlj5kFZf7lQ73MTxFSAvCO5TcwIO
HUusONXI/+ZdPu9x0FKT0uACg1LM2bE5Ui/Y7kYL5toDXg9zSbp/toD+L8ocLA/d
iSgZ69bYcmoGO12lkpDvhrA339ssvt8DP+XnUzAVjbZNVX2hSPK5NgEdFsB5pvBJ
NEhWZ9JpHWwErXOeP3r3JftVJliujnWAtMSnIJUbnLTAz9Ly3BSGUSoQ1KKNESHC
EcvI0JHlXG+E0+LZYGtBO/ooaZUts9YD+GXMHNJ95i2DssoFc2+qfMqzigDfdCAu
OwuJBw1NnCvygWpMcG5G3Pnh+v68BwS6Tv2n26sA1iH9C9COqGYrU2vikZF3K1zh
ZAM9NnH7XzGQUzIq3+ce7L4aXPduM484GgY8h1gOmAvXCiKJitKNtLSXAOrAUrHM
7s3RNSBrxHASY4lV1TCpITc67729qw8JBacFKS+wAY2TBl705ADbrxr27yv83JHT
9A6zsoLTswQ/GJ+HTFsNqqg7L9UBqde6RTFysin1vnxuk4UdS0nuO3GveAVv2097
BRyni++7TsZoQ1gdePxyHZzyzA7B7k/oMR9M59f1gig7Mf9IjZZCS5sK/+VSszG7
f0C1RfEiiSO7qCTTgviGPQ6CA5t9Ov3drlElJWX5CPEW4EaJSP8ss5ZPe8sWzL6h
LUVVIhYKnPw42mmx48aDQfeWaOiz1jb/TKhtzYbevN2FACOTWjVF6L0z/dNhgEmX
Gg8iayR0lspwbO7Jzq/gY+wy/jm9lacB0AqDIo0JPu/yIW8GsV086cwMEoaSFnsj
qAcOixqdlF4ffo/nAHz4CG3MK2E5fpLiACSYSuDs2iNQD/jjRlkrBZiLOj3wkIgO
CjmC+t4CR41c/6bOXaTQ/eOLOs9Ts868/SbGFQuKoP3yo3y1mKAxXEj6ZZIENYIF
IIdEdfUeig7aIwnOpPj9XvQpwf/OHo4uRAoR5chYHhIeS7p12MqnLgAY+eIPtfSE
KYRdUB1Y9b2a/tu9x3pF7pu02c8mBeUcJVw4wArkkN1VzmjEd4S1K9pnnpWICQ5q
Sd6r6d1yYGXDZ+84EXUozjcUP81qCZx0Xgod72VcIncuh/QZpPKD30h4ej6NF5Gw
NhBY49hOYQuEUGaB5WLVKJiqVvbb32YPnv6ETdcJH+Js2i9i+aUg4Y0xir+4b7XK
i9WqP+7QeHAQpT04jLS7ghrpe355sEi1ATSwK0uyVNiDFvmINmjKMQsXLeW+iN6w
X5n5adRhrLMOGLtv1ecEW3l8BH8337bwQp8cAZSQCGZB2gcz1JQgd7BhZNEcgoXJ
3ZzkiZI5T65fCravBaefKNMaj4fOouBga6+lLe5ufMb5AiXVnIJ2/Hfbu4QBOMRx
LOWVTCy5rlrImYLSlPzYYEAVUrBqc0SnOvR/OQMS8iSWCXEdhUCYLGxVJ2na36AP
5Q7vQft9bgJfsxxXcRmym12BPZ4Sc1poLITljh5KDAeVHvET8ROmBCmedx7M0+fZ
Ts3v0JzP2tFOnfm7EiaBo6PPwiZLrbspiK+XpMhTAXUKStSwIU+7rsJDQZpTn/04
YbQuw+VIBQlfelNuxF0bXgUL7D+0NlhGGTYj7GM3CHOYa8CM9R02hpfw0XMwLgpZ
LzQpROA78XpIMegzcZR7JVs/YinSGEHrqlH/Nmf2OVRF/ivAP3KObS2l9dWgtk/Y
IkezPf4faAMqR/XKzwRD3WiKhmOr2FRuWtKMwYnGW8RuWlGPx6lYzcaGaLBNyJ+b
7lTRkRvvCB44gNkSF4aqnb0ZFFmUW5gqWOaBq2mwgFUsruYzEBq35gIWumoZBqr4
aB4MH7N0XY3VKOi7dGQ5XeccJZOZMDV3pXZcyJpQf0jxRESvK3nzmnkc76n6wNtD
VuLrQWMSoR7L2n93maX37gNlwmjEGZDW3W40Gt9xxnINRcItLswVTz0s6oXwzMKt
SNJMFH5L6+oXskZBjOnUTwM6GAfJhZpPgxLjxqNmqZm6Uk8DOTK/L1ov5FNI4mlb
Es/RYX3OX//I4C6atQkL26lhLRcCkoBUUh+twjB+o6L3f9aDxZgA7TvZTOjU1a+o
DcDHCdKZPaATIn0tV0YrsIvdbTRhL6TfRnK2f75BtuFajxDHQ9RyO2DPDOXMyHyJ
rEj8FSBeCJxnEJacUalTQlrSesihBFWNWC43YcnPiYyBgahSJIfb8h3G7qy3UK8w
tjcPN20P4i6G3cpHVLYdAk/u/+5e51rEwKYrvFS0yqImftVDz+/R1e9BMoQSoUyQ
DRMpTrxgvgRST3GgIR9D7YW6DWRLNJkpzUKXGRtxRu16MYUyuDg0xSG3cmYcDiXG
hpDQuLUvNlNl1hQOfx6tDDoaAvgjWznjdNwKUAzA2Px6/9SSTdH37bvU7FmEbaE3
C9dTmcDSljyuS825ic/KOn2mlLcHPABL1kkY+9DBY/x1p9I0hlStDwmwQV05OhXp
sx05ZJz8UFkBGBpwypNVCuaY1g5jIxomk0nFF+/AHIc4xE+VpgprVwQlHM5S/82K
KDokJNAMyS0EPI+s17pX0/8AkWafYopv5XIC7J9ACc6k8GAlJz0lqs5uLrY28ovr
h8OpexwNFKJ/nWzqEIz8rXxg4kol9x5QYBXgRlkb+9Iniww2usjsDUtzU3F1Z9fs
gnbkwvgJVEXsWCs5A8k12Kl3L7VQaGJNftPDbScQGAP8IKyN2dkimKqbW8LHE9Ud
S5ZE4NYsCoitjEwqt25CbUqoB10jLCpfhlltvVbXy3WlM/c7u8M+Mpyuq2UAOAXn
ysJz7ZeTmLhLyl35CBjKZ/rhQEE8Gm2dRSe7Exuf6RU6MptWuTvQv32U2Fvq32Kg
XULxf4sup4gsOFsRlwZV7RhiRTNQ63vms49Yvq73cLFPJMeFYVXPRc3LQyQzOet3
HDwOQfVdMVc102aPsMbXkNIA3zqCHE5n4Dry0HaDX9mGlKz4MPnalP3hyNuoMf1z
U4hvjDr+j5xyEozA4fCh9l2Nff/87S6jxHgq6t5PGqyiwyKSEJNaouHnwiO0+KgR
SM9OFLIprJLzq1pAT4rMThudwoCuiQoRIFi5+OnvPuhS7zpA2wJ6mWm8CAeeT1LX
LzsYH5gesNEGe1Bx+hAhlchWRjVnwhpu6CwvftNtKpvg5hLg2TB3Fssec06w6k0p
jCFBZgQXPnIZJEE+Jgkwzxrh2Q7vX+yw33+HTHWxv8Sutm2tDD03Fj0T5TBz18Xt
O/XAjtSei5/d5MoLCRrxp4gXAaAiJ+3Bqs+X2k3LEqVYGXmr1O2FPSxQ37tLNKBN
oDWpeBNYHAdiPWY3Eu+DA2kuUJ+Nc3oH45Zp+Edb/j/kAyh1haNAYBRFYSEkMKb0
L015bI3/WipTDB8l/EpV0GPslOLpCj0hXVFP8FzMwkQl789SkvNaYu0kZrRAotz5
te/kDx6AzuOZA27wT7YzriM/4wt6R0kkHYrVmuC/5/iebqZDIRB2CcQhBek2X8mG
kA4dfWE9TLNh38Q4Naiipo0scdK3wf3XYki7047C6jgLY/s6+ljFVfKoRARC/5bx
vYWyupgCBTkV36sB4rMpyZPir8xyYy2Dg5n6zK/jesc+UitfEpuSDDPJ1HtOBP1I
ALDnwrossLb5rHTGP7ZKLW+PVVbjQ12H3W8MFNxjDIvjmHEHdrmmVd9/hVMNGa8g
W8uN352pLCiMzt4bb2yrdIW8FkLq3nfvzop0w/qQAksxebqqlLPgL6TNPaQe6Zcq
J6m2SDa30JXwadZoN8ma4cosxRR7XkQG3W3P0xfqCFDAWUZWwUBGxaahCTUZGbMX
hspFw4vwodpQPFbJh1BMT63YwT8NOrDvMA89hI4RbMbtejjq6sBVumI8mpmbO4ff
ix7AmSaGPpd6m4RwfK0FPwdZhJS9gGyIZTz3SfxCe3n6kg14Rv8qnJOcwvwGMlpt
Ca+3DGK/s7s9+IE5a72VnHFLTug01ScgExbbJ98FzANnt5Zx96z1I7wZpuoe3qwq
APbKHg1Y4EvOPQtRylknlV4nS6ur4rzqEC0s6WYpY6jhbCx6DQE+Scs7Q9pehE8e
yN8yo0JZpPJKyz2udP/ttL8qlVL4ofvm+MDHq8z8Zkg656F6uUc8Bgn0n0YKdc/R
rlqLWijOpWrKCcznYFmikG57zMkAMYw38fpeKPTgcOee1KZxn8NTgfJvnkX3o/Z2
/gIiOh1MfTLqDpM2VJ688uMvmVApuc79d4Q3uDJSj8Y1CM01XakPwzQdA4/XqwOu
6eyDgE89Lagly/qtM0sdkYBsGjaB9kqSbyhFU3LpGU9Lz8qh6nVcaYy/0LkOZFt0
9lejQEmGcjv9eXZvysQgK2jT1mmdlZz74nFlgxjG9Unxiv133LlEeoequz7tzshk
eQzKlkUlK98vO7OXx0xqcdi2hJOWmzP0wbwQ6J81Pdj3NsOIDGNS5jeastm36J/c
lcnwM8nl8+CkKbjH2Gq6vMURjexTSzlnXdR2/nRB5ADOXMU03aUgSpuDQHcqqy7C
0QUROZ+37fETSBj85bWmlc5d/oS0GMBn2TNk42F1E+sXuoVLIn6YxF5cwqh33kWR
w/P1H9bSl3wo6j9B0Rp/NpyZlCkt0j7dr93XcpmjTgldbcfqnfXqUCe/ILb1StEv
RQ0a/SkmmWTy9XQVTNaO1OjW94/J329ryIsjJ0uRTElRyW3CYFXyw61Z/mIKvQVS
jTcjghDw4Tymz03N6w6ViLJkD6DPYORRUE29yt6EfqwB89rAaOApuFTbh36wss2u
OhK9+w6x/eLOVGKXe13ze4VAvVOT4pSj+THmmhDmVjq9VqmCHZvYL7f8QxMZMPy0
j9aNTVPzqznk83UhSsRyBXVPIKICQyChmnNpiA9Tvg82Mae4bwIdS04kGMn3j537
uGW4fqnvVD7Ixk9jwxgsqxaZcabC+5JphC0ySjrintLPIRaIeC9OJk71lPDLOutf
LylY3d3S+zIhEmuAnKznXFIfZp1eVFQenjKjyWzb2YWIF2DlUwQ/nZECsXGAcuTP
wNqXOh4XaLih0XPZrqhF7ASY8y58b8ueIXfYvx2DGaoC4ru45zpveyYrLTHI2+e6
vWf4nLkc6Wai5yP4PzxPSMw2pyun0qKcsq9obPfZKaH+v+Fjca3SRVTQ+aZJgsvr
g6hxaf5i7x2Vx8sSuXqhzMwiQjvxlus6jiiknmp29j3c/ok81eU1ygu0A6dQ1xru
gcWFSllkcpVrTb07LvMqma4gLiFTYecuH6ujQRUkugAA/H+b5UZ+4U3s5C1im4S1
nEVZFu2a3YjF8BL2KGEe0tGpQyWPqYbU7/bXSgvnkl2pT1e87BxGV2iHRAzgnpj/
XFl4TYw7fO1M0BrF6HKp6TakE7ZT+0TxjvmjHAcDwmqVTn0nzF5TUp43P1HlwlaH
pxdjz95t2PkWVRbBTxVeyt8nzaFzZcY34KF20KnlMUBrzDyZfan2wOWTj/F4/hxx
sBlmTgfnAImQlqox+V4Eon8zaobGcmOUjFQo11B0jv43K5vW1R9udeMqQdvjt85S
E9wlVIKYouLfqEs18GkiQEsY/Iw18WNNwChh4H/P/3o1Vojf0KU4LpqBceTPKsDB
5XW944zysZPd9Zl7Z5ORP6YtaQ7z77b4ZKVHl5vF3oJUYMhFiCgNJMk7Yf2rjMOX
/z/Fn1xQl6EOOBClqAJqCrx9LeAwnuoj5c/qgGjH1IqlCoxx+3ZoDKo7+0eqtWml
MABJKrI5VonMfJmksr9C3iDARATOgg/nSZ6RfDi27TwLedgnyAzXFVfI0qcZDIR1
3UWtPcDvTJq1SD8F6QWxlLwG+ajhFdl+x10+LpLzAdR4+ytmyPVlD+ahAskbXrGZ
qZ8xQ2H0Oc507Zkxc4pmNu+KiHU+2qxZe/raHJEUZW1wKC9svVwdHkRu+U+BBuON
pdqB/zUUl3NzJ/37EuqQPOF6+l9CHpz8C6hrZY1tcVE/fZ3U3+RuBPe77RWzP20D
K413a6qSqspQ2aHm30IUB62anAfMhe612Jf94WD2tWu+TNNCSRpm+3RCP3iDAtRq
OMCb9TU4DU2VHpAhHp/b0X+XhMfbcZsvLghuzN1GXh/D1nrsWlnqQ/0dJOHsMkqg
X9ViMpCfYof64tQrMLh6v9nl4hQdm1BDN2zvJNV/3t3gMnX37qm3wetXSfodP4OZ
DUSirmiI9S8klOQ+RhMkNdTs5YDaj8ZWnp8Ni4FFb+3vXl/fyvQzI+HU+XVs5Yxn
PgreGZYJX4FCEFPBxMjicbDUTiYxzlVg5+TeIyP9B5U+lQ5FQ9Qch1OTC3n1F6dF
pZa/iuSTXof+upSJiRjziUC3hLdSxvp5NTJ7SqxNFrZWLymNT/EdR18IqA8NNefY
FJyY7tBtfznIK4IewJRXS/pMsZ9y4mN5qs/fZJZ5gJbjLgm381VTSs2af0Fy15QW
YPcwclwTROl0CVRunKSIku2QhlOgQdhk44dtpRfGRSZfShvEBqFgWcKkF9bJG3JU
mwIrAhL4ohKRRIghTmVTwUkz6IbcHscTDITmrkxvf11vDKJ7qjoCujVVmhu4FFo8
2zwbK1xtH7sDzJtpfAAjaR74iiKyWPPs1bfR8361qHNtt8HHSnL48LbMTrE2aQO7
UfORYSDLLiMC8smcNLcVtDPAp7lMSnwEMeX+y4lUYBKaVlUxj1ZAb5TSOCsFApM6
cRMW854KNXxiPfdzuVuvclDFkUDKPx5N5vOFqnIOjYrGBSwQdSBGlUrrB5l3wbXe
JgHy3llBbJrUgI9tPdzlvmqCdNmYh5N//XDx8W5Y8aALk3jJsyJIiIEYQziYV/XO
wLyYVUK45V13wywwp6rF28r8/2BK0WmhVVeSDpgqwIoOkaYkMoX3E+iwhEibDhKm
LoX3TZMyQF9Z1FrSotRTJS+p4WW/KbLe4Wx6L+xL5lDnXbZc+leLVGbgT2QbgCYS
9J/6uaHLfxnSrxU/2QOycv06As3Yvg7j4NImYf9HWvFW7L0wd+rGccGiuBmZuRNo
Jn7hWU8qBFQgI1e9CpSdN6LfH52n7x3Y+fvztdxJabAovUFu7TFK47/utA5YXY99
jWGPn67pJqWqHH/Xc20GQfGuUrMgs+UQPtfb0hMKJFDnfg0VGrkHzLFBwhRu557u
Hf7eG4DHNysqWRozEfgG1yVQVERwLbpUyLOM63sY4rYqAfzOLyIVy3E7ievQIEnY
8e/Tzj1Fys3zSL5BG6k2O0uo35hOY91DeZAlzku2ZujXa+AwdxyKa9UGrHFf33V6
r7gTU4Z04p/fWE9JKz8BATXRTffC4DlejjffrurSRNI3hVetp4agyBjSxUEzubZg
LDLGjqPjxv2VPqK30HGfgaO1waG5RvnHEVvu0dgow5FeMHrMW2QrksGKnoZhLJx+
/6+HdW0Wfx3SySyLy9bVF9QQwM1aT6J2mzoYrs/0H0g8AVE4mX14sPGtwC4uUiEL
gVyTxkhNVTiz5src1esKceoQ6Wg0L5fTgPf0ruSNE3iZN8BVyCnWT9v4Kn05QUQp
BmS22NwWy8ecoikYP/g+H0XjsiINVIY9NeouxwD6aPlk2eGrWidvZVdY/29DyeXe
S+5SpAG23SvRtH8IU8zynz1olYXJcC6Fvq+gNaxCOsjL0Ebbx1aojR41L6AAv6c7
GTwa5X4C7U5Q2PLn50+7IxoBbV3FTeakEy8/WCI1D3huWb9HqWnuKK7XLC4QfA4X
uHMRHiRjzlcpmT0ndMk9PcWdNbqI42whNu1gPcMua7qdyc95HsYcdGkGfUZaeKOt
4zRmIPInoSVBK4pRSmOI5IpSM7/AcYofy96Any4nOI3lDik4VtPxrg/N0MrWkbSS
tXxrKHbtTarKMMsxJ2yM0qoQ08PieDczoJv76i1B8MOCDj1xFUUL9zkre5paE2X3
t4F7EFP9AEFhgcn0NH11lGlxThWVAK+WZBlwS7RItOVSKf/9iioUACrCKtctDv4Z
mgMCC/ohLzcY7wWSDXcyy1Dc5ke1Qp0W4PFEAHoMWONVLZiu+KAoQpmYqs4BaY2i
lf/GMrybcYBn++cOJ7KuF0/Sn5fKS+D6n7sBQUZKUNEZ9z4Ye8bAbCPMBpVBGSQU
dC7AHVSDTygJIK63ErEI++J8PrzXpE/xcszTxnYImBX7x6QV0E3lnV/I97vbrw9i
bxqaOj2xuzmkUxc7BWa7BHWciCWuotXb8XcIMRJZmMWt8qenBe1VczGAwj/MKWUZ
UJ9XF3SffY1d6NeUAYkfMdcv3Q3PZhF8bJ+QGPhDd/hJ6OepSrNPF07Q3UCNOqsd
KzG4gbxm9whuO+M0/YKFq2gpaXcoLoJbP9hukGTgUFwzINJpnPSIZEhMiB0nof1I
vYbBgSSoiJBSFVyV1rqITssA46Cw9YTW05EQF1IrYSswaXsFXe2QnTXrh3Poz7Av
RyBZdQ4U783c6caSG6l4bvMkrlSk1hybnSu50Q2UY+28xRBQ8BaWTV0Sv2lSTyxC
SnijkGJI+/jOEjsFUbhNnMWrv+nY72/rxTkWSZt0b9o8odpy0g/MfYpoLAZB6bxJ
jDrezPBrfLSBgIRcHol9lon7pzMyoqHrutJE/sreXm6I5CqbKBcD+GROFUfZvGo8
UUZdFx+wquuaxYLIllSolVHXiNgDIjgVs04NFqodIMQoTi/gclr1CVwYXI4Lc790
NeWDbc+0ghckyC/QvvCChvGo0SAucbvowZne2Upi61kRrz/McrE9J3tyxWKs1eUa
MLjSRnYAAJRMXL5gCFyE1r69rV0/Sj+SNtg8BpdAQWT2+xRz+CesTyF8mMXwtSI0
tIjFKIV1aEWnpkjFFO/T2w4aoRPah5cYmsw92bWz9NUWAqACIk8YKBF8roSKpyjl
FSVp8owCFESfEBlQX7YJrfg/kolf9AKuMyjxlYCxOCIAKtVawFtEwvqXLg0A1qDQ
V9DACyN7FHJJ6fcJep6MkVvZzYGQ9x3lSqoeR6W7OI5RNXchFGvj2lTuAlYiRb+7
LgShg6iWxj/pCa+qw+RVebcDzTKevBR0AirSUARtF4iX9J4AW7Ylk0b80rCRftFT
SiHrbWYLfmsJC3NuAOL0bT+v7bmYxMWV3qHnZY7jvY8LTfI/intgvkAUA2N7Nge5
qaoTJlVybOLXnYFDH0jgM7+TUXuJU/YZC/uTQ9mvgt5XjasNayLkFsnCHV8vpOz4
4zykm3XL5XWil9GK1siMrKMQ9n70DVU0BNg3knR7X0KYqb0+gAI9VN7wc5RzlZrM
V+vYbeFKFFxWvxCv6Ch0l0OhySSjDKDq5LVLxBSCfXGhr1PtFrmrFEhlwLinbSLw
DS2Dmb2xermkiQklWSm4UDNUbPK5Wm7OeqGzTliNNSQdK7MjcpeeNXYhpeTr3LvX
CrLCPfwSmrxUAVBX5JberBNK9jVZotmibuq64Vai3sAlnkNyle0IzWZ1zGKmxFb9
9uyXJsw9eQcByLC9zBxgqvTpt7b3cFQgCPly5bNPrB86ubfg6A7ODMysnwnXPFp6
JJhHmd7YRtzya+laE7Rxt8c2sJHVnnLm+89WlHSYcVkGbxHDDPUHwBrumwOZuTRO
WfQOg5AOTrL2WAvrcUfwz80C0vb6l1DFWAxbMx4aQzlrpGdEYqSuSDCTIwH88kl7
FiBuHtsE8aTGUfqeZ0nvt5Tc8A7ST+Mdl7DbZci1LzQobhwQyIwmnlpt6TwAqQZP
RBYWNO1ssfA5snSYxk/rTreGRZLv/sy2WQHhMdu3hnCrNh5vGS3qs94E8N9B2v89
oJLzxuqNOphVg4JH4cW8J7mFMLhVzTgsMbOoK2cI+bqiQ6OS2yRkCWOaD3Q2EJZs
Z3WjKXsuhi4vaLTu7YjR880iFym3/GXHE7xaooD1ci/rGFElmmpVutkVKzUafwBq
b8PMcxj9p4yEPLVs411bbw+X/QGnbp2/QBi85U7VRXhtgQ9ZbvdH/4Y4864ohx7m
JDqMSQxTANTyPebd0p70Nb63zi3revWKN5vwvUu+5ajsLdpUU+SenBtFqNgZtzbc
2Yt2tJHL2gCBwsbq3uqOC7HajKk25pe/aoJ9CGnnIEs7wPf1zaOAsQNppANB0fMr
68ojFGorox1hGAD/jdqP4xFdmrYqW9uDgoJcBqtioeZAuwcMpJb3ROq1YcGOijkr
yAOi4BDMxgqNk3GCgv90zV8apyCrPULpYnH0OuMZWVvXqEbLUnOs/ZSpr92CL1Ug
TsD7h7VL2uRPegFolYTpFppVl5416wqMhXBfMKoamPQsUmUq+cZvatuq5fVd0Kz0
1y5jGjmErVPZSX9tVct/XcauB5EhFxRC5VFzq1W2jqu+MLkrYcIEthury932kkX2
nAyf8iecZnrqsdIq7IlLXMw1mL6h6l4jS68yMMvvXYMKyoh0/TAgzNaFqOcpgnBu
7yuiyIjdroarfTtY8gqfzoO7b3xFqQr1A4fKIW2nsIbhexY7wxHokwYUyjy/gVsD
2Kxv/EAFw72eN7HOsze8FNPTc8yzrL7n9LR4j87kbOF2Hmdi1WxAcMyyjy+8OWgx
XMJEiqC8ukQ4RlEOE28NHNMHLz/iYo5UxtseKsUnXX4UtSU1/YoJgCnCDe73Fb5r
ULuzxPCE0DpIQJnwqZ3x7Wqbqj0fO2JPc0svj5+Gd0eftw0U4prAMos/CVg5F0Rx
JJS93ppio9rYnZNgL/TGQXNzfKrZCCZC1m40YWminyxsgzWfs3fIlIXV8kHybIQa
6tza1RQ5hCJ0dQOsi09p6+Ye5i9qRhG7rev591feOVtsLx/gNQ4CXJig//Y15a59
fXetCyjvAg2vFw5cAji6QWm8Ttw1EaEZPCBAgFMEslV1P9CgxsMuYwnTKrJK8pU4
VG/59BznqqCtlOHbNOfZ1rdDpzwiQyS5oILpEDIunm3nIScivWThOL+a41iZ//0e
sAnJZen+E20jY2hmD6Kv4MnfBSr3Y3CLr6VqyTYIkWP480ywID6IP0cbgtuqv1D0
0bpOs5mGJOSC7zhxQt/ztp1vkGyBNvI37g3AmGT+9IWC9kt2kBL4tTH73SysIO/Y
a5+cfyl7BUH9CK7qYU7QZXa76gm90mSGMuzgBoMkLWVuYitOqBn7B4m8kYP2CLdG
ilbBEuX4uijO4MFLbg4JVPyvONbu+eBCRq2yyx0SKXaMBIsXo5mzIdDlui71YRrn
kQGXS+SZLXCEjlqgFSijVRkwM7DugI6XTY86Et/t3rFgTzGthsnmnpMZGui4v5J0
9x+Y3X19qHG7Ya1kIndfwZ6rmjVZORlceft99cXpRyMhqtIz4THI9KO6tQb3+UcO
v8mV0gMKc88P3tuHlb/jWFXMbkUlTpYlmGET/VgZxLeP1ar3QlOA//YDOBcjV3AL
MV4QZto6MTml1PjxSWOBe4AcNcjX77G9F+4WbZRlno0sc/R3Kwe14nfuPET8rhDc
skoG+xVKQ+N8j1mZKiz9QU5nYQJjhV+C4Y7lJ/GAc1ZUXrwBhntCdv0B5DRNebNK
bxKXR2H6EVs7YhhVIuZ0SiIxuzRTOHzzEmahPSjGM7tS1b+ipkXfRSKZ8v7w6Fzd
6PfVV2nZF3woDOcJ4F3uK9g76+pgfFbfCT+wpcD0UifNBXEnRDfIR29D0XYCscNM
RNmBD5L27aPLOTKGFMVMJpvagMjplKWnmjzJdU/FZ6TYQJns0/QE63XaBws2V9uS
sIw2TYaQlbOH3onnUXbi8Poc23PrJlvuw5Xyb8Lsd17WetNn1/S+GKSrEWEvpy5i
1793AQ0vQY78yIAMncCcaEAQJSYq6C4PIyOB+sY81cBtXrfwJuIakNiU7x1+r2fu
Pui+HXCa22Y3G91JtWRDbFF22b9ElqqjXSVTetCaXBnD6UGsDR34gPvMu3RGAvlu
fDVFzvxcjy6hlu1u3QhXJuPFZsxYDiPI30BrjR++DELc31ERQ2/niHPpCPGodwJN
dbeH0OIhe57Xm1L0VttJ6VL3ur4rqU4PjICEnit4makHs/ipqwlbTbRF10mwObJ+
JIRdfkjfHaTiq4VjogCTNHZW5ujpz8+67V7NBL1iSvuHMoX3hLSvEMT8oFXGkt9d
xc02n+WLdhe2P+Q7thF3huPL7wodt7EgdUq9zgNBM39mpVQ6sL9BQ9IGWXv+wwd5
Lu3IqxpUEZnNtLRZBOGKi/wV1Wwy9V+8UF5ZxAdlljOBEvthwIW/uXoZg4SYvRdz
csEUOgPYFmbnt5LepScrqrqPt7iTnKkK7DZdws0opUv3ZMa3SKB99vzeCmAottAk
ubpt6QtVVom90okGwy+H9iBKXBT1Zu+jRcTUabX7SJE5Hq63L+RLUohj1vUFDpAy
1bKJeOkZcEwz99V7tvjUJ1cp616qDFS8B5cAv1ApbJOUEubiEl3pWKJhnG6UZkh7
q1UyhDycDxV9RpD/buTwz5TuZ/2rkhpPjSNNjekeTFCjSVQfNxuebcM8LBej1CSn
CyXGwpe55iRLc0bqV4hWZjJR8qX79KxVP5QMTqizQAAIy89/22tKrshdNMt9XQKN
A32al9+WZswNYlXugkuR4urJrcZbZiAX0XbFjCCfxrCJbhkrTt6cydHw004fxZCG
wfryAhlim13b90o4TdoTqf8auH9WQ7+0JKtfBJ8ZrBECSDDfIF8UI/fO+SKmRX9f
h30Th05Xz1f9Vg5PrjZx/WmnnmsY9Oov/esGY99jdGXhmoHS6xDloZRrMUl9WhNj
IlOeelCtocoiM+WTty6Qk1QcxBjrB6Sl5D47gR4XsioY+c88AI7fH8jozJKiBBXj
ROcMbX8DOw0vB7pQKXvD1XpHvVGFS/+RDAdISODvpxh7O/5gMhEGy3qJFkgmhTp+
r8ZEIOLaG//XAZ2BelCItWrJljJL2eFmUi8YacXg1IgCqQu+ROWrYveUUW/ob0yH
RTtPeugClpsnCnSD1PKX0XwH1p93lgwJiHQ8WAmBtLuLIJ6nWixIA72fmAG48ltK
OHTtJA3TD+Racdb6Skv5TvAhf2shBpNa/d8jpdVTToLiFQvSUjBbBz47j2XoGQGl
dRSZLOMNSaqU3//8+jbRCF6wB/r8pX0bUEuMEvXGLuUocqbZS9zfVR7p5jwMTwAX
xaXbNr2/tkXkXK4JE8JA59H8YRwDPsNobkrZco9rumDTMZ4SsrbMBz+dg0g8OHw1
DzShU9R6vuciOqiUBNop93dY58Vuuf1JnRD18Qnt2+PMplEPLdzHWwYyUDEdYX/E
y5nlHEZR4a5ND0MEh0rY9BesFzZDvkIHkR0LNphYWs5WyafSPFwXxPXrDyagqoVd
aMHFHkpD2QCKQITS1kjj5+KjSs8sPTTTBMzYT4YqIAAlzi1sTXtwooo9oQ++AhJ9
NcvN/GI9o4Dnj3Ikmr2As5Y1KtITtgZZMLljqOxuvyjeftCo/pUNKWFzSjNI4whJ
IT89bLAuovhxKsRIPIViDkP7gmZYxFS2zBN+vAFB5lk9mYufJwdeevgwRnz/Gpz5
kUP5o4iOU040T4iFGNLOiWxgSOLCk+d3GaHSVMCA9iGdT7EFxtPrmly19dcspW1k
o+fyN+0keztwP6lrjiYwiEs37GG/SmpHicdHN47x9CK/4DNkqcLpLFSvHFBYKsF5
I2gxj+RNRUs48cvfMsf4Paj9j7NsoMiVQOF580vRmBb8+xa32Q//kYVNVBy6xkiy
BfsHiOGkIQT/9tHZCKauBg1ZU2i2+WRMfWRlUoAaRg8cNRfotOHhMmXbfulRbDry
pC15UFsnYWbgl/ZThEvGVVboOJg2RU5qxDpUgUbFZYGceRkxeqXZrEXzL/m2jz3p
qo659gCBHK4Nl5CgwlhPJ38YYuujQPqfWF2yNDVZfXJjWDvLdpC2kHScljDIC+T5
QmRuuPIOQxH2VcjNmZ0zOqc2U+q4YWddflpo8XFkZveT2ymkIZHW3BMo9HONnfHG
YICQ93If0NsAPWjeeqZrP3f22YGtg2566bMeQNPdP+muC8M1z7+VhaE9cbl5ycXL
bIl3GSr/2fovgCpr1NIxe9tsjI5cGSjRaDK5ZOJ8rIcJiVkIMtgyMPdYOi7Dp+4Z
f9YLeih32Mw6YK2pypv9Owoou5YN5iM6vBLRQEtEKUUIMGyTUq9TPVMBLWUjIzaH
+avuKiNhetJaYzW8F8nMJHF9D3si4pDTI6/KRNpHuo9x5bI0bbTKk+rPoI4fVkh5
b7uuvEZijzvo7tgXZC9WEB2SRCvKtFNoMDh06r5U/LwUu3crHt6tyBdu25qhFC7D
XdtbEzkW1Ee3Z722nOYA8H0z6xlMzmbzEPsCEnpIjYRNiRzW89Fiw+JDXK46prBv
R55JFnPRUPGwjF8BJE2WtyGfTC2uoHxIj+ASWYeuc6Uovg1GdLu4Et57HYxsB7oL
d4hIYY594hMcjJby+Fye5jXIaa/r25q4/UKe2RnWPre0hMoqLeE1TFNK9yQg7uTt
6AwPuzm0REARNbnUEoKg4gq2nKQ2/+kMRTrn0LPYZrhuZ+fzk2FGeovyA1zcng7/
EDFy6lBRXbyhDE25roPZwVTnwMfNHfdiWgYv8vOyNbwHt4uCrPwQpv40j+0JsQ9v
7Z8vatdDw6rwUTnkE51nq5/fwGL1JnFTXSZMCM+R1rw/w+NQFUekke5F9HmpbsHk
iWAoZNjeKwOmw9SrnLpPMMOM4h5TfP0vf0Ktw05YxXvH+Xhi5PpJmRRwOyFmsEee
fO21TjaN7rYEVn5UFT/hotkmMx0sPQf5dV7LfLX8bL8XBOqHemB7ZElCHEPYSc9v
x0diQpBt+T/FR/CXHuN3K/V3F2ejgqbnAa70q/f5dzmPtxYiyLbCedauZO4PZc2M
cuLxqFBchrYAOrXnmLMeGUOn2cyNsjEyyh3TPAI5bdRzh29P9yOyM84yOSuhc+TX
cxfUFv189py7D5K1iESgBXz9FxMoobe6CmovpGx9z9jEcJ65alg3XcGue4eKCjUQ
tlpWmbfdiUmjPYyDreBd9Q/CLdpyCapHO/qcvhwG2h8kOWXjWpNRZnebqyFgCwLM
v5WzYV7RyoMK7B1MCCigcXDUECx+y/hBrEcpzf3etXwLtFyhNOZRnSEtp8VUjpm1
GFvTD7aAEqZrnr8YRQ8jRyOzEcbvxdw26PlACqlKvvxIts3DTZaUQo/v4NnM/Im1
XaoKkWAqKfOPBAmLK4BtrIfcXAcMGrLZCGOQDhmHHu8f1oQNCrzfAalAAorN+TY8
9LUVNkt9vacA+JHIIx0Yey1v8wKuJkBcwj79zyQ0aGMJ7kW1n/JkxKoTKk4S8x9g
o/4LSP1caS/OTBoL+wBy5oRkev5PlicDSlcMgc8Y4SWg2Si2fg1bz/Mib/x/LWec
eKzuvXS6FgQueI5lu6LJ8rvpoRTNvkayuG333SX5p9zyo8vgpV5iJwP7/JqcI2OB
3nmY0qfNJp41O8XNz/vAiZ+exBAXf1wpX1sAw5fCZ/ZvgKJWyfwXUtyZ59M/EiEY
H2Ci8QaBISwBqe2N4DzgIJE9rLWtvMp2sAMOZcQn+lMs7M2R6+6udbOBbGjeFVwo
Z3dN34JvVndbvwbfL7P/zGXX5FeTfgOQHWTpYqOHyJl3PZK4n1uanKZFraE4JxUg
CekzdcxqTRSyH6Dje6KS+Fof5jEQxuqrYa4aaFlnc/HbR4IeFT4o5Xfq95m0i4v9
dCAwuUDXp+VxGmc6l6xpH6HQFl+DJVILMOUQjusYVapbPHlu5UpfK/AdVYNk9Pkx
HcmvSbFYlaVUB3T7zoEJn8xYqQaPufE5+zNhq1pogv2uN42hWLKjZJigULN7/WaD
pRgl3/YbRNjvyGa5vdgjDXJ8WGj7byrw72AFX7hvZ/U2+AWkd233auvlx4tE/dfm
JecVgpWs73SaIVQ32zdo7A+h8LHJrtSgtGm+DAvO0AiIl6VVQSprzHWpFxwz8+0b
i7ckbFSkpklbSRlz8iDw4woRAMOcQ4CvwVpNsF1tXc+1qtLGwLNxdHcHTsWUq4Vw
HVwxl6B20oyb2/KzGy7392psewZ8v8c39cYllICLUSV1f+eVWjvhVAu3GfvBQRfB
Kejja2wzMJUoSHJ4M5hQYNy+aAgX2gFs252hGFncyNABBDD9OYD/ZH5t7NcKV0gX
lfOAsMks5E9vSnMCUvZ2imkbA/G/m+pUEp84TNP1n+Z3KdaFXY7hpfN4Ljb3RS2t
fSWtYPxf2jEjOUshxa/YPrURBmNCQAIQH8SFIIBtj1Ss/bctpUrliM0Ewr2HeemI
Jle8C5MOk4xdM+IuuRx5oiCOkImUBYf2RhpUfq4VuaS/Q1KH1xv5WoufeAQDFdTX
Xp27h7BTI/Vv9Z8oEc25/wjxvS+EpH2elYb5ELpdYSU6NxUg35nfHdJoHckA35+4
9iOBdqeWU4xhK3x2+GSi8ZqRNDM0ODNHoUSHBMCHDzUb95daI3uPz0/q4EsFlJUL
QZlM7OeKlP+J+yNBh9g55MGtc+STfOkVnAJ0vfnP+3GAlBVuc2tf44kYSUnboGQB
DwCMOJbDzIvEVzOYhxFjl1/i10qeHc5QRukjgTXOFa0MpFwrWaAjfDgd91SbEH8I
6BcuezC5kQ3Fsq5LPNvMXARWpUGIo88PggvChaCXX/Co9gxFO31y/ihrT8UnHzHV
9PHh8pz8d+t/ja8gUo4H9TDfepGi0YpxmLVuEg23TfEvR2vYwRj/GmUl+zefFpLh
bsmECuJtgVIhmVQ0DdDywpUovb28p7YUgyd8vIQjYvHTgjh00npOI5BBSAlKlu+s
FajZ5ZjzrKzQldSrBna3Zwnd6+kyEgZ+CsNUP1iRQTwI4vyX+mm722GIXtrhsgTN
XHcPjpcZfqbsZDoFtempIfrlICj3I2JIQKtSBtXp0okzkEG2o4zo+aF7Cw3oiD/P
bFE+cm56b8ZFLze5ptXS5Tlm7qoa+he+G93PYtqJbuOo2Gq7Sr2f/M2L8zQtGegK
abKwo7pCLUK+ex9yJqwaJHqXV6qM/2sPgUHux3IOgsgwXUs17WokzidIWUBn2EKm
Zjy1lY4pCLYVux+7Li9NOsSk9KpmrCpK2vPdX/C/sOzHN2k97nbpfNE/OTsmo5LA
sriMNV8DZ3i2PrBqxthFY+0UzPnYuQG6R3hcG6GaccRbvflKzKaWDWRv27OF+AT2
ttsxp1g6b6GFToXIK+oRLmxaiuFfJVzgd0Y7Jcxok3nDx7X+ifQM7+FUH3LEtu9t
2ZfoAvVTa5DJdWxa/EhY/l1DdlJo2Tz1RqUvc1qJvPIanGJD6IYpSHSc2vKrjUR7
Fa7dhIsrZbierWNoj1HLQl//p32uK9iNQcoZgozhbnoYy9Wkgz+OXceW6mQXt4DW
SEq91JbowYm9QJkSZ3po5gKeWNaYxr1QvdcbaQZR/uTupkJKsAstHBpBBxhkRwAz
DaerEX/KS2t0uNOO7K5bvb5tf0Cedn9oc3WPMIV5TfyDy3STvE4w1gn8yJaOAFM4
H2MOqTat+9FMUhqJhmBbAp5R09HIHQ46emBrz3K56BDDbYNdxhJd7LG9jjbdqVv1
uxKTW8hIXXvedKu0zlMU+TwdLinGanMTQ8FoKk0CbVnmNjZjFKaWFcwWXTp+kAs5
ZtN7rdFdqtHLeczsJKxXiZMHGQBZGXgiX6uAGn0jQFREUEdA/h9G8lukvDPzaEe0
c4kouNUSAWQHFqGE6fdv9rBYJtodfTcIgaMF5RSLJAz7HTyHAxtr4h38AxRs2Fjs
u51sNJQ+2JMMYsV/W/kSBMhh4I+MAq/wTKzNTVKI1rfIKoo++W6yOcO5K5pqo/af
oL6V1MJ7csMMA7mEiufcXbJa0wlg/9ob3yfCAF3av43mzGn5K5eI5JbduJTK7f/N
HXFFLpzRWbG7lXk6QwwVX/qPWegGmOpyyjuCsKr7T8jAYST6AciqTbPBPaXckSmV
rFdNj51h2uBzn3ymnyyT7t4mMJVdfmfJUww2/ODNK34019EUZs/NNLCJXts43ZUl
teD9pLI30A7vIUR4o3iVzM92230C3AlW2ozOIZ0smrCRbzl2l7M6O70SMJj4tIsK
Nk9JGM2ESJkBb8O4IAjzgukcrvHWqLPvh8fQ7rv49bLIt8a9fTHyOK9m/ei/9E8N
zXidnIbgmbZQX/FgJ3ccGBwoucDffUlV6v427L2FFv7esVqbYptKVmHp0Z8KcJOW
FROky7MrPuutvxkt9QP602ARGSQ/hIIPw4ne5JKrHIX+FIXrUdalZTCfwCBAJ1Ke
3ojFTAVxf7P4zyP9taE33bTXU774439vS4s76YOZ1KIxs2q9C/YGBFKSn4arp00x
pJqcNAXLC1XmIm3fXsphoymNe0980U04EJJ78ojXO5+NUCSjleL1/t3u51CzhHx/
mU/iDVbup6h62HB+ddwQ+x1zyZKYts5JZDt+XE+xXk3xOQSKEZmZz5zL0fKhkSKH
ZEUSqix8XIj2GKSVfnxmBkar8eDu1A+E/6F5y2TwEl/sVRKKQWwqvOhCR6eGm6qD
k9OurY+dPLYa476AskHMMc5OlatYq0/H3Vyrm00Or1SwVNwACSsAf0V/5y8ql0el
3l0jM2T4rV/nmuneUNP/uiOPs/QrHdKoKRQPsLXx+7TdhISfFat9H6jVvB9+vwfF
lyidaEk7fyvxCXpYEv9lWD5pjebvH0TX5r89KDWHBRV97Xbk4e9S/qMIxmLVabmF
UdDF0pVxgWnGHmPkmB81yuQHl9A8krQbNqBP45lkTesnzxPYkBEMaPxfgQQm/7YA
ZCql+LKD1w8uLuXMsmFvF/PYtdjwmLNJDW0w1rVW/ZuU80OU0E1LmB2Q14j+dkfN
cAVhfDb3OwHZO6uDfeqoVUgBI6+Q4PfnaEGPGEGbk7Moh5DHkednofxNzHmKhKJ3
6I1w/h08tnxp9WS2h4Z3t/36RvY9YP0KjR9qtwWC2FOYIOmf7klMZJPk7Jtz2tId
wC7Jdr3zw1nHCzntUpUaRveSs/pDbT8eBEHBrmG3M+zQrhSFU2NyBASTpvJ01r3/
4FNTSAEIF7ekX8MqfMXUcLd0lm4aJBp/ZNc0GZ8GM+u+WfokvndcWcdV0EWu8we0
eIdZQluURe9aS+udShvpyyTmiUJ8t93UXnJ+1jGiW36/fH0+kOyywEmvOlTmAzf/
elO5vIoooiELSp/CHjsNliusY0T0txky3RleOUWObuFywZ4azP+RLwPAwdoBtsy0
nPVL4IVHSasm/vfz64EtUOav4lOx9TKWFun5qRQZTgdPPz28zMRF3gTdoNlnjykB
kzBEzW8qn87CYZ2bMLcVD/DfLJL2sD5CV4c6K7V+tSEIDj8Bc9peL4trB69Gqc9g
kaDa5DWmgleSwplFsgdZhviwIl0oO+5+/RO5/6ajOi75bZajT3UqiOAAFDLRWx3t
bd+5PYG6nmHI3+Tt8lFXmXFgJde+FcvfSZo492pDYbZtu5s2xveGsxCA4zA/Bc59
loMRFMU+MbxE8xdmeeD2LVKnci85ZQ717w3oaglQXhftmd6rd7kErRA7wiS33S/C
cEEwic5FYiERaCaa4hdb7gj9QqiFXhvibuVjOLnzhFJD9N/jNZ5j/LMZUE+qm2R6
tGdAC4Iu/+jmyFWASGWOcARwQtSdWXicdH3cc7PBGxa0vnzUGlROqfGB8EKyjLYO
BQezdcmCHsoP0ZlkU/kTsvL6Ez++sI/bYoli+yv5dABkxLb/BoyUTbBNbW9p5Wt/
G2Ic/sj0vWZvcVY+8j2i2z83fUCUP4WO3K7U548sahfCUnYKqGEI8JkyHHUPZQJM
JEQnDMDaT9O58nV4n4gpLG/2PCEi5JW68HRr7Ay2Mbw9RIDTsgsAwX3e1Ka5kldj
ISEh4RoANrQV19CsWfmWdQyCx20kOHGp/j9DPfn6+m2ygsSKM4KakbhlNKAH6RhP
bAPFKULP/AIe7kCKew8WbrNCAK1ziELkSFRrrvGFcBsgcxLaZK1LivC1aNvaSA6v
+kzYtm0QsyiqmxC+lhe1I6OWazDeOxTJYUKb6GlfriA1+g4mxlvdCcZXEX126YNe
52Wvt4qlFAcwuNx+5V3yRYSPUI4eP6LoVvLOSYw/V1oF4w4lho6rHN29iUGCn/Wi
QLRkarTyn0rzhPHmrc/CbgLzNQvWzmMmq/RAUUaCB8MwCbZxf+SvjLZ7e1CWOn29
mO4tLF3IKHmscwaIJRRN3qq5jEO0gOnyEujjBDZj6AvmiXdcYoZAvR5/kZfXxjQF
kMdP7P3T3k3AZF49DgLxWYdt8cBB/BfKs5fIIJQ712uZ+EBaweJCaAmxEUYEDqKp
2175a7xh+Tn1tmGLu5nw8uGt7tbrljlcJKYA667ESFQbL9f/TVAP3lSdrwz45z+r
N18g2sWuCLJ6lqZEC4PQn1cRWVtYaIGlRhzOENWJvDgpTAX0I2upiKFGkF2UHDH4
JmHBI2I6eSjaNV8ifWV0phDfbN84ARjaz/+Ufu1SsT6kgEpUSADHxi8Wxf8AY/03
IBaRckTzwcVGYafrcVv6VF6FRGYe0VOF92YSH9vOJvLhHbGxJ2XHrDi53VR2MUVP
jWtIsKnVMqoUwxo/e4zbZIJqT2JfS4mB8KYOWvkXz+zbq7HXt5SIlxcfGI2ccYoM
mhYiAZWBwLcEUzLzQSieqrJSF80QIxJdUbjyPimNKwYckAOmfzPOtahhO+o7Qyix
OJXW0Nst9P/aAuixuhG3Ofk5kmhRlWscNqyGSaMyTNkCS3cfgSpwHiTGLKTyXLPN
Hb0IVqHXQsUTyOWBP2qFqG+GSYZyczdBk1XyvRVL1teHUHq89ji5R1LHQr0yJQV7
FuIZF7sUAwZc6nTE2rJsL8DbGzMOEylW0uriIC7fveUclAaxc8NoBBFKveoJch1r
dpwM4bJUN7be8RXJwbpEiXQZwtwu5H4A97sMnxR/xew2zg0foX6YdE1e3uhCu8cB
RH+51bctTxLqr9Q5416Qxj6hGSuMFXDQEppVs7trfqilP6R80BnQKat4nGIRevWi
0pLNylIWjIRmNFWpOvLrfKhcidCIQ5A741xTVIqX53p9r2OIW45iN2cOFHvuxevD
gB0MlUTUYnMkweQPizvz7hSAIy5aCv+7fT/2Zs/1TAcpBOVeqlrfuMtcGBn3W8Or
7DqsayGyY2f2QP1GI4sfHRP54EcDrXfv2GfBWtcPZ6foeNgjLvtKQvaHcJlKkau0
pSjM2AvGOLUb7Nbxmr2A68EUqUR40bEMjscikumwRKQNtIbCqcz17eqe9YvSF/ss
W+4nNMODv00eIO5XmbMeSjY2R4ldC675DF75r9LrwS33d6HSN6LLw29ADdehCE5F
GVr/qKef8W8dKtyX1Hy2DPEA2ursQYpqDwHfh0n3gokKe1mUfd4oTeoT53Me8KZD
B4Qiaak+pIy1mrlrac2hKjL6PKMrneZPQJXan0ZFrxOE2ZTW/AdUPLbl+VD/9eDf
oR9fRKVsFBYTy0rbovBR6P23zyPQIRtb/5xS2q5XKf1oCXBQZ3WbtSzFtGigZYxZ
a2CsMjS1XJEeCtmUWGPSNgqZv/R3gXfpXcodfMkuFEyA2XOKGG0jykD7AxDPVfMF
MDAGevt38VpT1fcAyoZ6MY/bIXeJKN7+onWs5bxUIOhQf9hSTvhSywE25jFc6VVO
osYSV7YK8VQj8kaM02RXos3X3EEwJPFulkc7G3Zh+89sXCugWw/nXtprwR8b1SuR
fbe93ZygSwlR32sc6Lo/Vh321ygu0LvCRtxvv9w2+ODF2tKguS2VtzJlrq8kx+mk
Mre9625AJwZumZOOw+v+WNiRtcMqEo2RbIv7mnR5jBTTLbC68Oa8z1l3pQBCfjm0
fz1UA40gQtxRtcpBnzqaNxrCQpiipX7UnKus6Y2RE4iK5y76onjie6HhQKGIv8SM
GHoDhoN6XIga1+wlb09TeaKU55qPILwmNWpbLO198tsiV1gvH312lv5YwhLy8TBM
ODZSBuSm89PQ+HDojGJ9B0eYbB882hMa/DebJJ8CrKDf6ODd9Gq+7IwmgwKxw0rB
G9QYlmR04gt9jIaOKhoJBKBvMjETRBTJ+uZsD4ZWQPIHKcCAeaFvi0Q6+GUM8gzV
aQTq96b551Emtt1s/ldAXZ0sBUgmZeFd5BaK8qPjqGaAtA+2tXU+smOdwWj08U9Z
QhsPXQerqTQVPnOclX2yJIvipTCk9gpnPR89Qfbefj4RMPROTpAynoZdD95Zg4xR
IE/7bv8lrAQMKIEYL5LqCC6uY9BUgLwI2CwOfbPyxjngBGOTuK8ebgGgdJQnhmtj
GAvViYBCg/wZxdT+mOyNs2oLNcFMqCaxjyp96t0sJAbyRU86tGxWirZXtT/lsxbC
u/DLl2zB18yh+gLVHauVGrlpd6rmEjGPbWuz7aSX5MNiaueN0eFqF1Lw5rhfpOso
XWD7BK41NeNZLDFXy3lEZbc/mDX5ECkhdqCsZKA6PG5+b6rhz/88vDTyynBO+Mw8
Ijrg4vaENC/tSfa5NOk2uHxZ3XVSfnU8mh/sP2GF1HwVWfX/AlBGEO+ufLycvldC
pXlxZqssKS3wB4t0DKIvLtghubDA7ZNQuXIuvZVnmz8Z70yVJCVXPOirghz3g/eN
U5UD+iHk+goXv24y/Km8tp6miHeyKjvfdlJmkhz9sqWN6sVP1ELjxt8/H8/FbOxu
Ah7Dsarot70gT2JgHnO064yAoJBLois3lKY2cIJvLjGBqw8mH1L8m9Q5bENL880u
ICEhWLiNJTUJGnBmCnL8/mXvtz/I1qxZm+z78ltkLOvPCiTBOX/fEBBQUIReTpra
uWHeSj2YvvaZrXs0WvODRkC2B4zmeUJ7/fngXetjybf7XA+wTOyYUlFwqMs70uJs
BLhlMSn6P7oJIvswpIom9FVlxoyCho8WUYdU8ll6b3z3OLsHH0lxeEvq5WF2kp8n
9J3dl8jU9JMeIeWCdVzcIk72zrQv4Y7W98ZMC+TJgbeRb40LX5+eZjVSlM2Z8tAl
8YukwbQzs3ix8fYLlFti0UPxOXNusLkJe6qJRIXT6mqDLoX6mx/xCCnLA4socgxl
k9rzD61gZds1ttgL98xeIVY1jIUqFUcw4fiO1LkPwVQU7Cy0bLIEEI2vb+/2ydyX
v2I7IkD8vLrdh5Kud7IqQDZvGyfuEg9d/hun4fJztOWVTYQ0ZrHie4Mu6bEDb7Rp
fMdmJcCtC35wM3Tt6MKBXBh4nzGOJf9FL9JsbhFAONiAumzEgOBd2VdYPJbRdIkC
/WNqaavu32EgOugaeTWhZMKY1lmx6y66mz28P2X4R1l6+WAafVjlrquqUqQye4m+
I3m6/TR7UAac14bw0KQsLx3z6t3WzEJ6YTuqT65K7yD657HlsW3c5UvCCJxhKbs6
YtQdTOImsj9rUWdFu5MTOe8yb4QiGhv9s7rDH80fbJJV65xibYm1Yx1hx5MlBUHG
w7t1qZCa2cc+nSLl85oyw4mYPVz4cR+LtwW6ZN63EiqXT+nPy2CScZ5+TuO0/hmE
4inPDmouWA5XOPymSBN0nCNKO5wXDNBNiTMTtDDg6VTIcSCiVbFCF3PqcYolaw9j
8j56Y70dhEgXVCysD6/sSYKgLZaTf+GsgVgZuPSm/QxQ2sIaDWUZGMiYABeoxUnv
GYs1xXVQ4sE717DWAQ2grpga+evkC7v29ZuCH72dafSQ4GIPLrV0OU8Ox4Ivjdqb
cBs6LvlhFZU/6Fr6Chz8PsdgUILbKeZuHysu97Y+JTXx7GuB8cqJcOYUueYM8cf9
WgB2CXBNzQxEs4qQOBWSjXGOxpEd9f40p1f5MvgtXJ8by+yr41kh8o7VKn2d9YHJ
PKnnXnKAuN13QzzkmgUgBMSz7SWDmD/htOXuuxeyTEVT6i/kndzKD+WaPFsJ7mk8
A3eWV6nGlcU3o/TSCQdQb0MvzGDcsD7n9Jff4BsmRcEz9rlWxB07vZ3D5ijQv6+O
afEB6CPa+LjNNjGnanhoQAUvZExjpgVrK+M3MRkv+2j5ReUmgLUjPqJNpEUosHAy
XrX2HOfpC/VZ4MUfPhPtQZx8YcqR3CkaqbAWLtH4g5QD6aZdSnnlkzDetZlditmS
W6yx1WO6k4p5M73B66QMCPADdiZrUPocVegsGVWp/MO2osx3Gkth5Xzsp9h8Zk2M
X/XxTjBapwg0at6ojp3A7Z8/+tOAVOFDuU66lU7TxB155Hzvrsd0g5pgjAD2j9Bf
Ih+Fk/pwlkhYQF9OPnl9eafc9Kmg7jSfubHMVlGAXr5TvWKVgiroXdd6+GD7jyQo
D79FJb1ps6B2mLib30jb6SuVYumq9J5e9ItQBndTFutyEAWuPZTKymJnwdLznhNX
tuWr79zxhaps/iUAgmo8EBI69lZig9+CQu0dpxP1NGkKOt4HPyvMUEo4WJC6jvS1
3mxWM8687hvEfnHJqq03KUZR3Dmhst+J00p1mTAH2yR8QbCVPXS4wbxYAiMX6JJG
AUJTqC9mRH4FkjGrKZJXfkntNxcsKq2JbGNmYLUWK2v+VvOwHrjRJyTTE1lCGFP4
HXLEIrstLcA9OXyHLSV4L2q8+/62GxrcSDgKbzJ2QaIOYwFMjMEWN19LvcP4GfWO
Hg4GEkWB9XGAM2T7hoP3AozIlwlGto3PURQacO4rfAqzWpbH0SFdzyRQE437Skc7
NK/HXZ/bpfylZ2vOBWWX31IE/5K6+fqmkea0XwSoYCTHIu/Z35CxYx0kub9V5pd/
HJ4EJg0+hct7s/ClDUggSB7rk/Z+tm9xpMCzVHv2p5AFTjFEKcFBWWCGqjbCHw0I
0o8wx+QVnsOc5CNR+LE/VKFFb+IFJNMb39TMOmueWTY2wsMQVKflnLmva/GhU3AY
1jExehXb4xC0Oaq+G6T6zQzkzip2cIGYvMlJldk+ASNlHD1loop+dNnK3EcRdKS6
jhruMx+EN8XmYkOjTUkHEiaG7+qO7ppvNNjEOReTNjeUIZi1vMiiOY4aZBBPtpye
jN3aIwdLDBA1fteuibPKRBdQvO7F0+9MuN0nhgOHys8yPm85Nl6oW4Nk3ZD0iDae
JW+ebjNH3T9tMESeZ3VQGqvRY/QzyqyHFEhuCAjZWa3UWO9UzZQxsrlq50flqqlF
DwHTBn/0Lo2/bm6jK1rzr2J1LI63Xofztuhv8Qj+R2Naa5B1pEFzjrO8K9DknfUX
fweTfMwiCeJrZSCSkxUOFeGwaoyGLqBSTl2GNzNBGSaHZvebBULY8cmQPxnSU5tI
ManGx2p2oIZcdJ30eI2LjhSaySowZz0HBj9bxEB7DzESVCAD1VFrtoclf6N0E8CV
qy731frTyVosTa14DE0tNDuTqKLqB/ukk5bJ0Mwh5jwCHi/jwKpUqQUiKkbanuUq
J/PINbmTmCQPfbRSxaKgIVFBQMSmjC67+mb9A92JXFy+u/P3AUX7LJVVNUepcG9w
830N47fLHkFD/VRx4VxK9oD8IkrT2ScGro2XPpUMgdZhekYwo2xzdRH/t7d5QXeG
QdkMu0Tth4Iv78IgYAbCkGaFXx4YdwGt3BPvAcFEAf/i1cR/K7ZJfiESS3G4d0bl
/eM71crG+pSeTg0sgb7vt3PJtCe3EAYxtFCQotrAo5foELBZhefmJvQr07fczwi0
xxhCq7R9o1VXxIPor6+gGiF+fWY0ngOcUaf+v5T+64WxCHEgNMpU3Rd2iw42I5Pm
yJEt3mmSTgHYWpwyDCKsmX5J9P91Zsvvf+s8gGe3tjEuoq2fRVcXpWy9FyJpPdZa
mwRuiugTbjYd2YvkiksE27EXC7WQ6fD5wlHHS3/mNTB1tIjdVOIkbIydnqjgETJ3
01sGD8w9khwODY4ZzSQi+2a1iiaIgnOS/M+2HDZQBbagOGZI5X4d/A/d5lp44bAC
MIpEXt41dJNMiBUCFwr85tTkfTLbcOx9lEqrJsWo8SWAOrkqtGmqnJ916jcDIdDe
QGzeHe5FqNc/0mOXQG/0qKtZZamZg5IqatkR0MKCIikMPlB3XJlxo1kiylfqTNI9
/KN/ZEZ1wCCT+teHM1IBW6rGeAHSag5pl9QCkhMN2UXoJx0cXsM75hSyIOCdo3b3
pIRoa++5XG9SIZde976a+JCdITFady5CZG0mtTlGshX5M+FqrJ1GuXwoVPnl/9ff
buQhwyhdc8bKMfJA9VxvFqn5QDUklvoNAA1y5H+jdszw5eXFliYRlQwUAE1F1yGC
4mCtGh2nKo+48pE2WKydtzf+neuk67ACN4lkgghPVCUxZ5Mwx3u7Ri9vvv4o0WIz
IPWFBs+lZjcPZ4plj2aW/qjd7FpCfv2TqEIEkIpWiw0QLeL7x3NDaeMuGW314gMj
6SygiLYg0zxo66DYvTt3t+FaTzWVSg9UnqPujKyLRM/6eJETNfN+NcAXFKiyudVr
xd50LRz3i8WfoFhHdsLXCMZ24P7Hj4wBR4l9Q4lCgkpmoG66qXPFRjAgtpz3CfIG
qP1FAzVZb5Be1oO2V2sgHSrdTrKyV1TNFqNAk1ZwqD/Ig2+2QEj+Vh1eJy8BBCa1
pITCLOkPLmV41fDy1G4MkGu4zCukJebW4gcHsLyhYofcVwfyh9O0tV5zsLLxEgEC
7v+GdpWGg7BV1u33Uofag+t+Gv9jFNXrd5/ACnlgUl6tusK6y7+8gN72iGAdUvc+
Xy+rlAWw1zuMLcCLVAK+pdN5/Nf1g4cTxoq0ULQwX43ZK8AvBgxTrhvpQLEy3MhJ
bcHfX2U90Rh2poAV4B1NjuVhUJqOceyjar2kgtL/OgduZqMD3g9bptFngePrIpti
q1Mff9Y/g7OyY4KAJ4JaxZf45cSej/PN5mXkQAo8rEjfXVIY4VV4Lu/sd7DWdgaz
JNzIpPb5wGEzwgil+Fn7IZRbHBfJTjSTftzvr4mRIzYCbRcD5NKNlt0nhdwRDF6+
Fh1Qg3tVrttTsRhqPSCxr3N/983bwntZANqf720n2oXdNB7p5KaM+VEyDI/7yCVw
6K0iJdNotHGBPGEFyb5ASqm2lELz2Fgbw4Tb087ksco4mUo53MAz5HG1xujELf2p
ahu8DRCON+6oRJjmy+kiw452QIwywJL4K4D/SePp1wfRdoPnHw2m0a2f/Pi+djWH
orbDI8Ai1NbXxjVOerSlHXPb3XhvIzT48HjEMuR2QghXknIuwn4IAThVbSYlBdnl
bNATMwo/i6lfZF47NQVSDDJITfd8tgt6NCOu2u02Lqs/OcO7GistK1EKjzxrTxIj
LJ+Vbi2lR2jiwDN3rulCTd7ly5opgdpLqcSlnHjDL4utxhd4Dbinyf/49j+gWWxu
QqaWcvVignoPAS0OYGq3o+Ma8Xy/Edi+tXM6IVCj11qAkdkh/v/3kWUrTPYFJBH+
0kkOrPLv3EE9SUlfi/6507LTM8Yvnuz2dtlKJuRow6dqDGc/EzvxUoiwqVieJIpu
vx435y9EAA5q7J4s/jP+yjL2kM2Ypyv/MyAIuVfP1qBnhC97Qp6fxGdDvd77ajnA
j1c/oiQvQfTUJw+AW9Sfi4fwJkQlRZPEAbRfeHy1YAPYWBo6mZM2K7dC4MQCPRPV
QS4FGDMIpAqgLiaxJp4X7jDHbm+yjnqsq1XcOTXr5sl8/8owFN/4wrYaaOorystv
klMsp6utf+Z4FyJHjQ2QcDW3NGvFE/IxDlpmHJdj/rOEefCofvgkYKkuc7m0AJPx
EjvIwLVgMjojtN3mjJQVRQzJKZPneYvEXY0J21/CjLO56bMnqv6GL+KSURMxuWP6
KJD3qzBpkahDFUJum8TZQfRT2p0nRm8LZb0smuZPGalJVFUCW5BO5w3ZtfnIOs4D
Dg4tvuNfk21rUYG7wLoGi23qhWlSWO8p7afB6tfY07GIOCWN5x3e7F5RyCDj2RFp
Y/nmqT5dEapf4qS/4n3GSLxf9gxiyKabd76yHQKCGXU2wJrmTvmoii8Ja42UbAna
hOiuvaHPYAb8h37GOVBjL+xIAcylSk4tpGJsHz1ZEuh/nzbK7UzqRsIo/ytICPDV
Qw7eomNo6Ni7FlmjQWQuXcMdjoZNyWoFdiOBL+QJ/81L1LcUkMSG6FX0z5URPuXv
l4f00TheiSRzc9wjGoEql1E4F69oEdyK98YFjgtSrdJ3LQbsiF4DsFNvZjHR6eRr
gz60N6ANmRT9nDh9jE/ITnwbnTsk2b7at++oXL4To+V2a8Lb7IgESRysDW6vON9i
eKhvQwBe8oaTLbKaqIf1nNW7KURniwcrw4EunDiOZN1EjVeM3wHVdUcnZveT7k5b
RKOQpn2qoWTQ5t+XmGKEuFmckWZvwtfoe5Nd/5A7oQdv1QJvL1nprIwPMEw0dBNP
Rk5KcuDhNaeUedP/rwI5KrFUYHI6vgzkNPA664/Z5Xv8Ck6Ee8UVket1K2JKX9MZ
waYmI2jE3hI7MfwthPYZClBN5XSWStl3pw2tYKbuvX/fS0ZF/9GXxhfMa/CMv1F3
in6izc3b/Tt0M/WHAd8lVdZCqFDA618GrTWZtt/gAvPZ860NfqzCWNIpqAH2Pbfz
xCDZOEejUGENFSzwG5kJABiJNqHwJ+wdf5Wfoa/jDrnHb16+XCvSEF9/KUK4zB50
x8qoGfVgcHzq5ED3LFNfbvjWrP/LzrY8a6mtW2N21qVeDQ3X1PRidwXKdvj9hgP8
a6zcroLAk0JK9l9f2DGxsYuMSXvZFDVYYh8qMsESxaMmcZ1L3deGemTSh8XCEHQD
tEBJW4yFeDz3XEAQugO56ZvHNDdOSMMziouFLw0koLz8cUDl34tzvo24KnSxfvp5
YNcjwy2/NUjSaCSGobPV6zkG9Tj5CyzYWilh7LGb25KlezUEmYsKoyJLm51iDUPj
dkskAKUYHDujyYs8M85Kn7NsTLOONv14dB/TPxkkrdLXB5HWuIhJFF37Zk/CAVEx
4nq68TIQ27UV/9c6+geLNHd/ov4FluN5ffv2LZ6LuaiMa1xP55kY8513cHA/a5uE
R9HrxfwFLb1SGvPjN+9GR74F0N3OAqWt6Dgm0kFftMyLAnrlMcyk9EwTEV4wbo5s
jDorr8m23Xzvr8j0qp25/SZLMVP3wj15HldcRtY26jba7rl3o2vPzExslAN4MfrA
8NWY6AM/chlZBgHG2i2a5sLVyssuevZRwRChupGa7w/vZex01HQJFiLX1wpil7ab
/2jNADflybxkAbDTC/tvU7TbaGCof5TC6cDKMNLALIUO7Htqi4ix3frI0TzBegRD
uR7N2US9ivk5UnuL0gg6qKku8aj28bMz9DqgDidsh5eNLcEbcat8bFpwoJbTJlPr
TKighkaWbjtSNPuTyK2vyWV0en7t0ELiERQadqLw6tH7UyW+91o4dN4RBt5p9Grb
QY+zZJT42V+WCnP5Ke++eqP2Eah8wLi5i3vlIgnLcrKSSsod7Sy4BiE9M8JOQWQL
wgpRfv4s8xATQ70oq+a1nXxj+1ZS/k4N3KUkHojS0Paz7vaFh2cWocHz/uAchz7c
hj6zLTeHASCfUQiyM1memU+K7A6pvT0N04WrwkOeVXK2QhFppW9G0F0OFS29z50X
aFLHtdIZ2jxiz6s3JgjJPllnW7H/RxcLTgfAro8sbYxISTAfcyb6bDB2LrrjYFQm
gbUOkUUVyVieawEhIFg6XIEXQHUpOypRQaqU7J9W9fT5Kj9H+ypyng2M9XpI5ZwZ
9SZLULE1OCHhKUlF09Hu59ViFrHyBjGuHHI8OKbaYwRC4hKppT+gUOZyoN/81kRA
F+zaaNaDWq3CVmwK/rLXqnzfPrpIIJoVbWC8R0GggIhy+SfxIYtKmPsMCAZ01MRH
mxl+QY8X66yducJcSnfPf0nqzh+C9H5yfmeyR3Vpu55IVE+jvkwNLTTuq/FkjgBP
nU0jBVluKKiwMti10DDrwBpA64hCvnxl7Cba/amQHLaR74OGLoZpwn6qy1spLd1U
OqudUkNqoaS1nQsYKLfweAvF5kvPegPbruXBo/3iEytpl6lQl0fkxxUgTw8ZGctB
+VN7jilWzia0J57k4CMx0HgIvdq7dRrtvfAqCBZCEtkywLwjILO9vzF7QGERVJF9
ypbjmJMAROFeaxUf8jieS3q12kEZlBCpxxxjvSTJKJD64E66JVB/iRhwN3RnvlkR
fXJEpzUujAlnIr/mvEME9pDIM+ufRKAdQDRxGGSLWdo6lcm26qu6fgXBazjTyM3g
bDai2zbCHzvoE8bJGCv7X8Vh4p+FGg5Wf0LJ+6srH/vSmb8NnuzToCzVj9wDFTIp
wWjmYmYoQeX9XHPh2yOGGqoqe2d8mcDF8da6ym3aVFyqXp2OQ1tMb5lUHGOPsbLs
3c3hVNZpBZJHVaz/sYP0t2NKgrmyExOkyauMrCK0Ft84sDuhFO91UerETarROCgY
DEZeAJHzJ9eevdRnKs99X1H1dWva5vB3A0Gv/iUrN0BYeVsTxcZVLP4QuAU7KlaX
OCJkZlRqV5C11OlnOMz5YpcSZQ/b73RXB1f73Dh7EfPZsEnQF1UF7fe+rgljR78F
JdljpZmf5pgDW7TSR8kQUXLnndp4oE84CXhUJOz02aWg1j3+gfJSkdX+GOg9CpD9
h+WQbcEGH5dz0cCZ6I6MHEH0pVDQfT0qr0Dajpr1y/cjhn9pkTYG7EcDf2QGt6FD
MZGAv7A67/+dfZYJko0KE9cZDZc6MP8jWZVFG1Jj4tgvLF6jFN0jPPFSDLC0RV9V
rT1WAXuYM4HZ7eut9tWDHMBnrBS/Umpz6WSDLZPwG72b1f9qVRkXm7QMNXgRqkki
dO62t/LM5XFrE2xaeddXaeexGzHTt+J7QyFqkeUv3pGgj67GJ4VxUVBUl9k0qt8l
Hf2I42GZg+Rdpv6I8oM+wH+GPXEcwQcC6kotM2qRgu342UzIrFVgfkhNQQ7CCGnM
BQANmTokOq74FA0/emZdhoGH2z0HzH5woTpr1gHADhnHpg0eALzR+ZCvKRngWjpe
VIoTjTrI3wWOKESmV9W+ddAjc7nhwbhMrwAgS5J67YuQbNfbCKUntT2vckn2L7tB
1C9oW7x4Wq8dNQCLZryObkUjUU3oqotbf48JYnABZztDndxAMezdKBr2ZVxKSynP
A8S82XvL1tliXDZTtOLFr3vI1cxTPck9lKbYDj1zo1E6VedMl8LZ4ZNB97Uekx3D
YThnRpT7OK7rS8xCCpjt96GPvu7jpxzccP9OQEXnNBH1bzZka+q6OMaEEUv1yrVm
SyYZ8EAI5AB/RyL7blHKIxwymnnnkvWXxIYt7aAYPvXVVuPLxibhLLE7MlH6JXXr
wiLOCyFPzNqz09AGPRHPaBppnJOz++qBhKAuolzqRHjrn3NHwtaBbBqMUsKbSBkw
OzfEyGVniIOwHjYVaE/Imi/piEzVNmmITC5Yn92KUrNsOJVouNrc9sivtumkYoOF
mmuXzp2PX42GfWhhRTJRq/u6C5XuXvlEM0n6EGeSkU9NPcku1PEdl7E1pMVBuYVr
zC4Bdkr8F39iE/iGnvtjMUs3udLc22g2Va+PDGY8xKg0LwsVXMObdTCCg7ljtEAm
JsTYcNLlBsTBdfoNTfjkIWJqhNlgnOBflF2nEJydJDWC/MXrFaiTYhuMfSwppiE6
eLl/OvIeqlOVonhFejxryQdNMTj2GmcK8OhyDiRrjQASJHE+4IwdfrTrlCOkXYtE
zhpDdbqxpBcfzKcHna1NKEGGqA7HyfG5D50pl56mm9JT9NHDERBKR9PsieeD5hNX
w47Ex6SGEwXzz3NQ/O7zCmRkB+Cw733YpiO4vGDp2P6ophhaz61gL1ba0vbwz5pt
vhBWsGuyA857WVPccP/aqPulBQbuBbvvejcTJyEj6K6DNH2jzNoQaE9mvPoRWPp3
STQjNLKglZ95dwrLLLQ/6Xavvs+smrGGJHzCvc2UjT6X6sgiHFf0iqYOkLAw/OpP
PbevHfuu2a591no57o/Fs21vesy5NpIy5c5XqDq7yyjYtYcMCCdKyynLfL0BlgdR
4LXMCnkrHRzrzXOY/ItdilhApZ3zv2kpeYPL8vCLMHGRbNTY6IpQwT6cxEZ/jovq
kRynCyPu0o6QdHHd657itkjT7bvT9rDAHhLqms6LcvAyfCKFINkVZqRCYYWES2rw
eOvsimyrO4c86OjKFNAp628LZx/HtJ4cNyhaNvh5vGPkiDD+LmURHZQegS32XIvr
tS5C4YnxfW10gMox/CaK5Kt1YaRgSWwEkHAY6cgvmJXdUjHyzsPXUtLU2p32nRZY
k5MjQS4ATdMDlOOEn7oJHCNl3U74X+fz1l5aLD6FHL4Q+np0xQymn1MRttZ5iRCY
orgp/ioaYXxxJDQkNv8i91xVMm0ePIcNyhXL6FU+RXzED5tbVrn9U2k+6b+51w99
OVjopCzQ81pvaKB2D7DzmSnEhHAyHBunlgZ+bfPKW32dVlmkSK0Ni3e2pTh9tp2q
Uau3BPMTz3g3AayE2JKLVmZPKgs+GTYmJA9NSl4PZSJhDAAaJLge35f62DTu2/B6
RE2c37h6x0EiLsioa0gn/gW2AHEzxbn4C6JSk59asWGIfC35VW5HjsldCxsULKJp
HWADExIP9beuH+FMSXeW7TmQTEUaVFwZRzXT0QPOWNP/Pej35YPFXOj8TE0st88I
SRrXM6ihBTLDum2zYMpFtrDa8r7cus74JxmmX9r4ouoqbZsTi41Jn/biDpmQNk9H
cKfukyzIezSq/6eznOpkG6Zm73tmeQHBJSrY3EUhya5m83ArVJrvsKZz7jbilRCq
4nUW2hm6DvyB3+Wyz6nzVSn+hXtdfa7FKBhZ5fdWT7xKZMzpMrOtumQdsRDaMG0m
wlhAK17pBqIdZWLCKOQrVOFucPh8ZxI5rOKkK3qClS9n6U/uBakLC/w6nkXwkr79
Z/rKSP2yzuLFOd6RdNzuYF02SC/MePkaDRs0oDsHfEXRtLQ51iv/xveU5eWWcNPr
oYiz8ti8GqfXpvxugZ76firmXoR+8Ic0r2nJ8h+rmi459HnSHhGYhwaa5pIlXRQ1
FpfqZvJP9TLAWF3TZR8JnWYouLB5Iu7H8WwxajAy/L/R99DvYPyzPb2YhMLhHSu4
dHVqO1lzcaMbTP3oazvBu3YQDkQttcqsFb0P4X6h/bQkGO/95qjza1dV9Q44RZD8
jIoiahUnBT9EhmBv4xzhBxZ3tOxnKQGZ6/yJRZP2cUUCtXRirp6YKPVZBOJpsVqF
hb4yuIyw2rdZZb2JChPZ2xPqTJwbs5G9LhGGO6i0VEGFKGf2GXAnHxXx/ny4QBZE
sp9Fu0JRe/UOFVaaznFKttMgjdgDuW+N8UbLvy8YFdQoAP+gfY9V0eSe5MQW9hM8
1/iUk3w8WglbCEHgKt6PIFal+Uj8kQaIyoXUQ7a9nH2bB2vUitun/7tqYd3pFkvB
AqAFOZzl6dgFqgBVBS/9Py5TfsRlO+s7xnq1XeEuz6T/XVSUZaJQStey4a/nsb5h
zidlQW7dV38F1x93v2+hvT2tMmeKbQAciknDVPrz3+EWgm5XEy0zJvWjQThO4ldH
4RzRm8hHDtg//3PSZXC/j9t7cgNXLVFDBwY6p6XmCVdXAXcvF2WUke3s28tKEfMg
qT+LGhsGuh7ollBbZGk210R65MZ2dX1kxv1Pdk1hJxtgU+8bIRyQMlKo+9781Arj
6W3ox/UCD7P1aGHQwuY4n0wu4AQ8EA2039NbVC3xyNvB/NKNBZuJSA1u514cyRTi
Mxz6JOEisB7eBwjHc0MTG6h08a9SjPPmDN/yEh3hI//IF6Uc/bKp2FEayIqH/Jdv
MlvQnKphtTBdwKq3hzRShPYfKyWfPHbWMiKMWVtGbq1FnpPLz5iXU4wvX+bzW7B1
9yzlwDnoCtfBTfUOkllZWi9s0N1ivt926rWFGegFVTaSaHsWz7/uNZgnk03QPhw9
6IEKrO4ILj9XNDWcSEgJ+wuQ1+UtvCo5eWLWQhD2sQxUNHjXXHL3Z8AqWus+6SGI
xOkHX5EY5POdv05MoAqm5L0hAF9YxqkKOEcZlGOH2/3aIpKXrUOx7kfT+npjTk+e
eIBaXzn5iH77IcEBCMcNUhvsr61QnCY4pLHes5SuTsQxK579zfPctzuHm73HPl6W
wi86WVDsEPT0RqyhCX/MybR5xz6xrsJlEDgt3UDVov1S+vqbhsmDt+TfuJdOqTBp
vu/KVi5x5CHFRXhu4iwq2noMdcknY/hTLdUVVeIakFyPMLFvNGm7hnuCS5xuH8JI
CAC//CqHeOl6HalCK1lrrsE8AYsaklm6omLa147QA2favTvf5skL0a+Jufg1Y1Sk
RHvnnoLLBpfbJCVTDBznY7fb/fF5Axjeg3i2MOAjY5O7Cn70lH/T1WR/8hG9IhG4
hx2iJKjDzSePF3yXguK4C3gE19WrMIHn/isN9N+Jo96R0R8VlwQyw5IafEZ03z4O
Q9AZwVX4gTBWaKqpMQQ8D8iCXOt1vKnQ2+W4TCtCjQzOxj5zJQyEXz7ICxrsfC+5
xlnCL1r9NhBx56qhYC/f9R+wZKvp82XO5iN6WspScMEJM7vIecWMuFazWE5VF3rq
ON2HuWXzfdwSJq9RUrRYqIUUAnKs8TyqBhisiiXSHr/guC7x0h69ulOLgRES2yOQ
ZZ4JJZ4VpclpL69P/SXMw3IdeI3ClDOVhbt/aAmrHFjDmdAU01ftlLCtQg7QcBXr
3k0GLDEfL7B03TK6hBMZxfkdWUUxpOGVek5+m+u+Nz3SmoCMbIKj6Jyxi/NH3Yz7
ROa5NMfszd1rwF3fa/zz8ykMNVE1xNBqIbT6OjR3ZHgl0zP8ri2dHYg07yDl+5EU
8eyZnrPb37Knhax7heYij+4l8CnougFmL7zSAo+0m+71AyAhQb2USMnlutVoOnA/
6rV7I5M6U5+3fDawmm7LWHpq1lfgTRtYxRUCY9tDabsCZuRfg0ns1sGb/DX97ANk
KdpNNBUecFJ0rY34ujrLCG+xjTn/xXhibkL3jCBo6bt1abfWRcNAzEm1ZDxYStMS
lIz3r9WcaV+59QwR3tw6gpIz+NPCbNuC2UxDMHK8urVlwqtNVrDWZG+VSKH1fcWi
/mzDl2Q1iWSCn826VBR906Rg5Y4uJP0+KGzm0ghWn/ovF0sU4M2Fiu2JtKrufuOv
f4C0XI85v9qj9rZGr3yAiKqZbZKjs/wzG8SXngEO4JAh3kFXxO+et6HG0+mvtDiJ
1AGMjCvsebCJWKmHGXtPeO/oJK5tsI3j5eiRLzuovNS8ayiH8FyPjUs/La3Lh6mh
az7KRRUC6Fy8LaqJjCH0/kCjuP32SqLuHhosSQJsg9k60kbyCxmqR/dvjLnzj1IX
mKvmRzbufRICvvzUQf+21P3Zf8yb/LkAwodJGkcJXGqTZp0v6rj1rlmmGLj07Kwh
0BOoK5k/kBMQfGVoogviHDjVPhcFd6N/57q4F3YgoC8WJXxHN95KuDiu66LTbl/Q
qXq6HdR7i2S/Qu9ABPt+JgmzzsHOu7WMWf0HkdcXKPZ8XybcYs8T2NM5G51fq0E0
dm+Oo0PsqRpp0ql+M/ogYSsh0+rXL8mBel2USPf3RNDnNtHlgjFnwvPfH7WB8fw/
BNDHmQX4RGWgDNVy76TY9HhKw+5qOelycQpWSgTloMWJdpar7ouhf+0rOky0TGOX
M4zlaA7QfhjhJib8KDOpisqNxgcyQcIZeB2u98FFHmRTFScctCNYducCkAnv2TzG
7LNjwHIOF56wG/wrwOVyt2NYmGBd/Y+cyPmhEu2x62od6ra/6YkC9Msc3VnjH64d
QuVli6fTV9TOfoZ7S+TWO7QNnWo9uhTp0AgyWRvVDVn5bzQ7NXQ7BLTZ4IT46RWe
56fP7AuGO9A5YRxBZ2WSKNW7tao925QUvyUbjbmRMySz7q6i3n8dKaujRNE8V/sk
lH/KnWl82u8p71+Q4j2tjQQSliDV/Ei0/W4kHjOSYHRjRFI/N9ciHBvECzIfv8zi
WsTu5LABf0dXQ1G9mSzw/2oOMR5CF2d169BiLDtyvrSGRkxcuaGe4tsb6SQzQ79u
zbKfbcqalLWz2cBLgJqoXnFOg0AP5vRyaoWJs5m1o63dOFHdpTn67N3UK+TSA1gD
2CzgKPSLLXfp9p2IHURJ9VY+HnUYpQdcLcJs/m92+7jKxo2CjTnDpgPCjGKboCzQ
RoErXfrvZgto2B8PSUNtzeqjmP0ftzun4ZrH6xK07vQyg4viJ5lEvFQm7LvxAFhe
T+FKioLCGCFFFmFFyE6cCeu+2yujjP8BNrcQuJVqByC9MK3tM64jXJFws+E9ZU6/
JnGdmIIHIM0kr1uzsBIlsEfCjgLNhz4b2LysuYSvk40fDMzQQUn9+kVGKZ5R2B96
9IQYR1Gcj8AqiRpyzD2lHqXeTy2sTyBQXSE8JMkxipBmcfYgL6aGRU7QNMtqtyEa
SEP0+uQtjNvrtNExv62SYof7mp8y1TC/FrX+4jx6BH8XxdX7AkdiHFQoUu/CAtfj
+jCJF1IvrV1YgkP+s5Da+4x2lRj26Msfl8hRQg9vNYyBsmUkJU7WxQDP5porGdKY
wiCJbrfqgXmwtxiFIQJFdOX1bXLmYurMQBLNnxnu1QMytm4FSYursciNHbXFQQlR
teYhvN4jcRKUHkhd1C4hpf35Lw8WbtuaqbapUlYveZi2ciXRgP9uviqiP0vZCnZV
d3zMM0RGvrY5nwoB3/VtMwocFb6l/hhepkKfwnXzofoVvYAkQlde3mzeV49wHNiq
bJj6mQ2xIJvmH7CUpZwzy9RblP2Tv9js1V7tHntlXg0LSLM5cNAjaD7HcKhtKdL3
M3opddpM1k83/dgFMu9PjVZbOP6NoBhfdysP62Ne6lYXR76Fgr1IsQXNUPGRM3ug
BP9/jMP4sR8WBot1Rqo3BDo8H/udbBFmRHrEhPUXlHSDDl59vt9MUF5oSSskhOcJ
LLH859XZpj+PhdcbqLFmFHotnNaQyd4XR1CKbnlxYmUsjXC0KiF9A1oEw3T2SdOd
he+wdf5garkMmkNu/UDP87wUfocjCkDl1FtolLxDQtXjJ4+cyr5jq8QVIw/337if
QjRq6oNU27AKzNU5p5C0GCIW2B40Cn4BkVGpGIhpKYcwmJ4T9NUE6WzGrTg4O44z
Wjcf1Zw/ccADhP6nJTHkJxyM43FGKlnhtPzJjUompKIY1Fjr/5WZklaXDTB9mNyI
XP2G4BXi6zAGVTSzKp2i/Knn+4Vgaj0p3bIzvoKLdMuTd/N+GMKsLyAAItCFlQR1
yEQqkSAO5u2yN5vlnpP1Q1scWCdHKGtc8y48lXq8XfXPPY7/HKetPCaeAxYobeX5
jqu3gjCROXr0WdK9BPpAFk1aqrsmNYFQb3v+ZuBU0EadPqK2Dk4kIEqr2FfyuDOt
DOZZnNcjqmKrLBIYykDKROuIjSeUOt+bvJFa+s2y/4gHoJlevPh+a/SVTvCUBnmS
WwzvmuIBCm+dGRYzyMOBcN/5YGnm8lqoEOLwLw9ANhDnPpeeaFGsE+Wwf1Bu5z8V
JoZ6/gWf+9q0zmXEhYjHKhReWNTaP1zEG9R6rZEZkpdnB9JP31zvpqdqynIYpooT
ut7Zp0DWVjtPpjigl4wdnUqE9huTHyzlfqmULQzyhCHwkUhfc6KyCUlaI5il4m6D
EI2Zwb0A4OgXOO4HzBgOMU52enWuvXlsD7DIlC+SgOAz63u5P6mUS5lILZzxpzCJ
oLMsuJaPlPGWFsj07PVYYI7313CAt1p3F9gGAqZagsiEf8lv8cS5VU4z4AWlGtY2
/8lCZRYHeHnc0fKIMAX9B8v/5WFywwUrHS7ck4jOFr1blixabtDseeRRE5IVFDm2
wMruQ8nVRxGvvbb6nkhy9+KVM1R5RMLyvdEbUQznsVrjZ+QF8bAjXlvt50/XT+53
BkXPph/qAPnx2VpzjsKPJ7xSkkfQ4Qxg4OvwU5p+vzEXR34fJQUGC1rcbCVEz2kf
K+lOsiHO6BNl0956rxxrYh8il/vaONxtZ3rDOnStTzyghP8sCql+QBDriFKld7Ma
9bl29MNwstz8hwh8Fg31u0P0C6hz/5+Ypq2sUs+VXHFImrFkolpohNKLP0GCT4no
KwJCMz76Mv+kddT4QhiYZ0koJXgt+9bSI9z9ZJAmQtmqwBEtgJrfFZGLeT+hMaNf
DDB7IbeVGtVjAVo7hVqg8enpxEPPjR15YceqChXRxPEnFdZQ2BUmuhAX7pZz7hjT
ZP5sGHUWw/rLyclB/t/VIY7Oe3DHqOvqL/IcSBmGAVgZnSnfqtJodmrV7GIsH2vI
5AdYA5UuAhN51CzlEzAxG6D9D6W3tYbGzC0XY4X54spjEO1vGVoKnExV12l5FKwH
xI+jurvALq8fihUNEbVFXc1C7qElR/SWzpDobvRaBz0Jj3JbXBYEiCXVc9tBsWZ/
M3O64M/qbheU0dcvWw/HOdYNYxuInzYx5tMStDHfwx4m6tscMGL4/Us/zEnv17Ju
mp+Wpr7HaUIFGXCVh13P3CFI27aY2V5PkOK4fTKCobeeHyU0TZs1fJja2Fffalsx
zPIvYEkFM9U6NCZz4vHeaMcZz2HGga82+gkpK/lYW+ceA7r/cn9rZDVmYzpXLFcq
O44Uq/jfRKSN2Idib2LNC+Ui42+Sq2zyxxa3sBRXyizvecpD2VNvVwZSucqOJiZU
fqHIbFlvxf12a3fQVv6bk0ci4BnqdCGr2sdOJ6ESjm7e6JJU/Bmv4BOLLY09Z9ue
sxDDdbLDkZcjcVeu5p/W/LwHdFfhlXYnMgjJPIm+HcloUaCMN1h9nfb1wrHMd0Uh
60T6HN2rO3T+tFltHDHL/bNb4H++bBLIxcbtiV4oCyXLdBILfvtAkuDFcESPJwqM
5KnDf5ceQZjw13cXfE7+xGx6obGNjwbunHbqXpXBXHnqIKLIU0iV5L8wpU57955d
Ha+Lj1rNRfWBEq9aT328S2rGaHGXyV7c9Ni1K4QrirDTJSH8eSXACgVqPNhHKhyj
9SEfdKnyH1655UlMkdYqKZeGadBTZ0jDtxLZmeTzh+nOG3hrOUQWSjjZEIqHExOq
7Z/IUJ++MGxuIUCT6Mbq08wHSt/nZbkDcyy0gc7b0jOnIalkd1qYYq/4pgfWdIP5
dD8qKqTwhflgNq9zcB+BUiaZpea2NEbsrA32wNDwdTBNI/Dbnk7b49R3yfpnZfIn
AvlZnX2TGNylCzMAQ6p0vKHb2//QbPv6KzpDIq8b0zl7zJVEdsDoTc+vNJbTRRMp
c26d5PXDq8+XX0el8XJNnK1KL2xd2Kb+SptSsCbKaMnPovV2NvQK3h0Qxrpu8cOX
hDtizzyZCnxWqMKa+K2QTxSBDdekO4XsPFMAd+geCDjExsO2dcobDwHlKDzlqf27
TrKc4mkgHKkIl10zDOecn8ZwTD1KsNEVbtDzgfE+qPw6ZG4KtTYOT0Fbh5DG/+4H
vMT98mswSR4smZLrm+4KYi7kVsPspt6IJOHrTRNweWk7h3V3jNKn78H1N2sLmo9j
IGd/CFe/rQF2zSu/4+5S3WHhgzBo1sItj+WDMIkeGuDg9xIW3uUMhecENocdpAkT
sIe29w9+gJ2TIdw4vqRC7667tJEmP8B859ZPgGyF4MztflmXe/bhWKme3mv3u+gR
xxg3k92XNdzTJzavDgxK6JTF+cKsL3EWlSV56VoZ4up3sMZOEolLH9PZ6TKZWcEH
M2BhvMvFNRYM+6DkJU9a9GgXOSycKugmy67I23ofyNnbeswobFD1g/2JYJtsmvpw
rsneUe3d328oM3oYN1akcgDJsFUg1B4crFt0KRngvSeCBVH0M1fkAT+5NZDKikGE
LvPY9vlfwCEtTrD8L4Ftcq07wBDd6f29o9Zc4U81AhziG8oSlry73Ht9Kqlq6APd
wph4rJSuyoqNHsef7L2gBWT5DSs8HVfC8qN+fL+Ahhv/eNZpwB2SnJBPJ0Xt+mU2
dNu2oaO7VHPXOhcT8PUcc+/3ia+43KcSBWNQj23IwiV+AbCbpo485mRKIXPunFQi
UfO0fWWnncEZTUqZOo5UK0EMjIMKGdqn92V35i9MLrE6MV8VmM+tOkQmDHkqhaQx
ezEO+TMTbtCMYKrrtOdzhQYIYDZQUCERwK8a9yDHwugFC4YTvKJblaGUQ0dZpYEB
Ujs/VORJyeeLmHRJHaLoK1M+b7D0SIycZhh/1PatvwDpbY2zhCbL1PQRbU6eX/eo
HaNqG4zQL7H4EaNS9WOpzP0O1uBHr4RSnAmauh6UXI3Bi0YLwyVQZuQy4jIFp0AT
pzj6uv7j2+F0boN7p+Om+UtyLqPmpmVUhf02o7196kazgibkZ6xE1bREHaQ3fHN1
R483KDJj1eP+Ti5ENeBsJ3YXDoqCqHFx3R2inXO1fpjq1ECalp7jD1xmjuv1lsUL
DK4b7h724ElFE0jwe6mG1WTJAFXHZDyAv2jmDST+PZXQMrGkpuM5pQaMXoutciyI
f/N5iqVHFb23QprRYhxaFoYMC6UMkmKHnT+RtV4DhezFDlCkCehEPv6IRn8Fz4RM
mkRc7SrHgIaiWUsJ+GalJnlJAfGVovroO89X/e38ypEFEiemIMeCwO5vTDn/nv1h
imP98Oble77FoeKxU6x8AuGgoUK+KMpTh0eyooZhPVH76c6OuOxwYgIg3ntCvRuN
VpTmi+i+cGXhmMyJ7s+txQmlfSeyT8UuDCt0gfTHfRhf5qOG0w66phPVkLOyZjf8
sDpXBJnMzVXF7DV6zmfcX3mYGgU6t2sWEQ0WrzTugYHxKQqiyxV/pWMkYWFEu+ES
P3dyJ5ImBtsVjBH1+oJi2U+mV1CpLnf3TJ4o2GKOeZ5YWA7tYQSP+ipk1HecZ5pU
GMrPbWL0J3l7ZOPPuch18A2iytEqXySitE4v6adBADajkdSMNwgSOLOz47unt5NF
veujz3OYmGOpARWrFlH9xe5SEhdFdrkgL9Bb2xRZJG8x9kXFC0RRvq7Goet7AmV/
V8qQ4cl4rYy/dqf/+tmEveyOKa0TldRVoJ3M1t9XqXWmiz/lwFqtG5eYHtC/HaKJ
7Qa4HYjTYjdThHUuTNXY07HO9rfjVA7GztL0ip2lcpVRFPFxNr0cZOII3I6Z7Nw4
NnhgSfkhxG2XEBeK6lhNO26Wq1QC4GvdoMIVeFoMQL3x41Y9wAbqesmShCQVw/PY
1HVclU5NU+jEyHj1sKwyFGeMemoebr2zrm72l7r1PwYTaYCb/gO5J86NUiuZ/Iyv
HcSBHHLf7QuipM7WWoASxhpLw9eIxwU5c397tnfCyopa3EGzgQqnpk2ScOB6J2/6
q5g+FwcuQ96Ol8WMZDDs8KDI3TL8HNCViTpwLMBW1+R2lO8Fm21MmGCAXc8EvwJJ
srhdiCqKvXBlIA+0NQCZu2AoLStIpPA8yxJDDSk6wrSKMP+FiahgBDJ3PX3F2BHc
ArDtPEwKqO+wQesloYtkz6QTnN5lMtpT3nuKOXaE7nu1UAxsbumhVTfSb9LOsJ36
N5dnyn2SNUDJWX+YtXSZtgtTBzhDKKc7T2VoRjNTKi6LRxG5oXZqF6+bJkr0cITk
G/BENUDSzsEMXiQWrLnu35piqcb44ETwP/o8HJXHsr0ndZ8FR0NC2Mk7XUz3wMRM
8v5gfuMnYDRnpk4hnb+GKvBYEnQhmAj2/zOCmpIkVpl+bJaFMT2gO6gbJy48qAsr
/RH33IhtnT2aWdn/yv1iI28cVSPfcCMiUATF39zP11fWI1nhvcxT3p2u0CdaaA0S
hKvjoeTy9tkcZdJ6ftVg1HtdHEPK1HgAOmYSSkd6yPLXg2Uh616kFKNgP0he2jTy
7jvEdfkH9Mp4Y7Lg27PrVzdfrkadDwZbuEUFe5fhXzb+dNcNCEnoz1FPYp3ho4Ph
HG8Q35/c5NQsVx169ppyd1ARtN0aTzQWx9Vjhesl/K27xku4C6EOt+syG7zMBy6d
STRi+su/fj6t1SfFlooS2IwYjFtnlQ9nPlw5yypN7COBglCjUQo2ZHfuGlDo+Jcv
AEKGUjoDXpSCt2gPPLcF+k/PMSoyo25dRFiOu0tvzLSQoinYPMKpR8Vwmtjl75w9
S06yCzFTfTjjZiUWS4lW09WTbdsIH5gsvAu/GtmvU/6IbC4XWmgnaLbmcEOOYb3l
AJfZa0qQl0n1TGidc7s/RPngEjsL3PpaMUaatdWNZuQGLoE7sGAZ0eoyRn8/hBl7
BBi+6Bgx47Dd5MY59SujjZ6WgzXCCyeKeRDKB4ozpkQVjKuOmMFcIN9laDXldhHY
s7kvAZMwC8ryRdz5yCYYwc67EkXrGZ0ZWqmw6kMQCtBMAtae6ugCLDlHwbkupvCQ
q1WZeiLDriZTJXY32yj+rB43bBbsLeGZSsE/A5MLJAGVgQMpHHFIchCo1kCHi5C/
xqCfNNVzjXMM44qm//zcCavErnGz5wd2vbR3oA60HA77JUdfmST1ccL4yoE+o5Bz
dVfcocs4ba3KZvsEEy/ZZiZsDK9B6oOZBlX+3jwtrjG1ZH9Vbva5vayJes4q28pT
LikLtD2DdcX5vldMO30wz5cHZw0g0nY/EZLwSs/9H6tTShWtyglJuF9YmWoJoGHm
VtAsnE91Y1WONFsWPpHpBm/e8QPxvD2I+ejLbJCtswIc3R21HbRYn5qvTn6kTnni
R6u4hkj5wZ8DC+spCySBbJw+m6P8jjB63hewUj93psYDMBXbjv6H4Bxe3/mRBzkn
sWg+rg/01wxL/0ZOY9OklNEGoRTQ203A6D47zh9knpcNga/QgvlmT43CsjeI9EFO
oyMR6j8EWZsx+S4ejxynGmfND0JjatllcEnMblKBxqWAIdDAvcR+6chFtQiJD3m/
n1G9TQnn4dfYR+2KIDM8Pcbe+WyC0PldI8dRF7f2bTLZ5HN8xo8aZoOlatGoZctI
b9yXI+4a2BNKlj15e7r3A3fu89921GuwC9GRCbET/7NqaWTtbeYfxTx5UkpslU2h
GmbyHttejOEfbr2jNHsLCzjs/WSfaeUk2Rm1Fsp0wTIdbih+40TW+0wbkWl/BGgx
QSizGcx4rI5u5e4fUDu8C8Xhsz99H8fPZKOnBrq8fXEenmRPQt7hDQaA0vStRcSP
Cq643nCN1FT1HlTgwBSUUm6SahySrN+7hcq+TTJI7DR3ULL7bS+AStE+IPC0d294
rWWzjjuAHAOED0qoenX3EvwBmaDjIXIUFdVvRVMCNf+P/9DRGB2tHM4XTs+ZBcZw
yHx8ymC07ebJLIuzOV/7Zk16ic9PNtZV30PIgO9HXLwP/VpSrrS4ZGNh7Uz5j6cl
281FHaoZBNb39QJPnuEB3EE/ZR0JqN+LFXCscY4ga7Ohqt/z13OzBgILwC6O+WS6
i66TN8APA5XO+KMMaiCZnDCysTKwF/JJJY86wqkfPcH8wrpLvkXX4OYPTGI3L9pF
kignhr+RPtFr2OEbiZZdUh+8uG5TOmD7m6vNILmFmcthspGOMS9Mahmu9BX+uULP
gDHpeCQ0afmlk542x5xtzQu0sgzkgmzJKhqyEnQ3+SMKCkLzsPS9qeiZgYKcPp2g
tPqUob5TcTcJszelj3l2gTHTFtDGIOFGC+owhucWDpw2Ay/BfZ72EPvpO1bSdv/b
6mWVxktuMJaJ9ev7tc+XW8GgBhLhjnHVOguqo9BtmcP1qne5VnZLFbcJTFYON+1N
beDs9kP2d5qDqzpbZIkHIaE9hXvhSrAf3gsVG/Zp6jOJ904iRdt8QTgYeei7jFey
06z6/3nJeI0siGOQ3I0sZPq/J/auCTqIvlwbuD3Dkad02Unxmh9AoAeov8ldW6Po
lPxcBlnMa7UBpBPsmFKfCv1tWle71H+IvnpBU0JCYua1+h4Zr6ZGuWo+jujp1OD5
frchusBs19D2BirE25+zgLEfJbOAfBdCGHOibSYpqq/ILlTruoaeBZr/CSmoYpG5
eDGQlClNd/feKi6d06AZ90ZQBbFXfvGqfAPRqTsWGEQNAO3s5VLljue6BZkmcP1k
j1AOjkg2nLwCzivAKEvEJzFapYDKRPf8j/zotKDrcv3VfgULxdYKIr3YTxwK0piO
KqbmwQGYZRM52QQE0sLt1MZE9i6oQtlZlsT79BY7nJAWJzlQXf2uRWwc5uzRaeHY
OrqazYGpEIGRS+VBB6VGEyfxe7fxFXlMczvQEb3aV1YWo2I7aXW0nNl2ZGUnkZ3E
v89Vf4BvXCXreN+b1kOD0G9zdyeTIGXwyDbqWjkzBSkbfQB/4sDUk8cRgHA8nUz2
1LP6EbFKk2+qix8UnvWwgG8SgV2G9LHld4rLVI/YEOzplvQNWYgD6tPnx3zljKQ1
px/wRnkhyzeiFwYX87huuVK/1laUIDbEjjsRSipyHVhiIqHJFWmBglJKyd+RRlvk
9z4a3irPOd1VoRm6LQdPn2Il6mnve3LpvggPyva1/D1fs3WJluscO6hGkvu7uoob
1n+2WVmnzvatkLRDD9Y+xJ6viyvUhJu0tFi7IYJ0dMV7VtdZmUXi0ks+Dqn7w25m
zpVdUiR3lrznnMNg2NQBVFzZbclYCnoGeaEYtpgcqBjvlzNOA0llBsyBWmuFtYk5
MdD2aWesqxLLR6lnsoizEXlUEQ8lUci4YyqnFEJe4IqQGS6WufwqfCTBpElHHVpX
F6V8CA4NLOGVRkUds0cnVgf3RtQH3huYLnBRlfl12m72mBxdPoMH1peyyLSJytHM
NJIbO3t930Np9Zkxid9Wdu+4GZupSrIKcVVgRAfAFFDPQCy/215QG1/mJiTHGAYB
+4vAwGRtbbfa3CvZ4GwTEnBnQ501TlwlBedFoKNcKglrbrxJIxEHz8YFrL3C0QPx
+NMCmCRX9vLO6HuKir1qOZTmQWfwesZzeomlwAn/m5WL+SjQovKTc79FexJBr0Cs
7SGCiCyMqdIozZsG8QxY5NG//WJGt2FrLIDrVifvI8xAuot8L5MGL7dfQIh69tY3
jW7/c81mWr9JmpGiMhiiwETQorIRMOIO6jbX4eoW02dGuNHGspgnIWOVlCf10zdn
Q8QTCPpdQDbXMLJyDHMHyyBniMGZPJYkF1+/EveFiGbHMEGp9VkFOLWhD+U3IC2y
4HFmfTfuMB0Z7a6cza+uj9SsUCdoiyreS64wfhyKbpl98xLWiR1qj1Xu4PXadoc6
dtyhLmXFk4jHproh/PCqB3P9Vxh6t8kTd+8qvi2JTARNIfdbaZwJnmAbxXLr/hyt
9QYH/MdqgcJlyzcUrAedy/fwcMUyhL4oWsDszXyKt/e2pRF0CyLWtwnxvS9S2PHX
lnj9jeSiOfZymb6X9wGDIeZtzUhGdF1MmPDI6agahCIBQQbhSBnLPAjXGYxwHmyi
Rdrzg+vRPZuOBswwwTORFBdpDkLDkpw3jD4/taC/H52q3JSQpQQYHMxbA8nqxJ92
FY8CDk1+UQpSyRN8Cg7Y7eYQUdT712kcPJ1vcE7FYYlx0TtO6hKdQxL0ZWoSxb09
03KvO8RIQ5HTmpO1aukHKKgzmZHQteL0KdXtV6R3V7ZtUblB+efuy4uijJnnDsk5
aVTtaF8wXRSA2Kq+kV4RUAJCgLzEEf2yqwwQUCA11V5WsTVdlJKjMJlKzzoF9cnz
epW6KzzdQgyOZOsD3M8sRqEHZyfS7QZRh8UsSvSKSYoiXjn+gjIj553ukBgiNjz6
jrm5WjoYrnB3Z3bLB3W1vIWvpZvyFz01GSOM4bD97RZ+cAJncjGBObN5NKBGCLQy
vHsJbHXVyZSJBz/9cSad0scY74v093oYO/et17RiN1BW1PqOA5AFbAvXRhlFt+X/
rAPSgnubA3cotz+PL0/iWCY8/7nKK9RkphR/jbTNHWOXkVNBF81Xe4xX9lOeStuZ
btom8/ZarhhSjIZqwv46JUSkkSoEGnxxW83KgF1Mbc5nQ++b4IhWhF2Kn8UPcJTq
RY72QHjGKJcXWrgHlJfOpGEYEZNbjUuS0VHl251o/EvVppOqLqxg2XEZEI8/egSV
IICba7UroEA96yZvqQ/ekhBhhfNbFzDjPLYjM3q0gho4vTq4aWNheqUZRuif3Dbz
9J317mrikxFKYbtC6/SzsqB5nHbK8Ci6suoYGUHSjwyL8jvNyO7ieYFvEWei0ahy
XuOuq/aW705/3JLgrlCLYDIf/DUKWY9gF5KAzOZmtm6t3lm7z85GJDmVUnnoWz4W
t6paLkV+tm26Tene+qioHJXJcVYGRriwCK8vPPMBRpEOF15Lo+4lRZR5BAye9T3Y
EYEtgFyNVMq+dA0zNlusrwM7YZTLL8lkgJrNus/mVrid6devOx9MYiWqVS8oIGq3
WbZ7PAwCVTBWrWRnhJjregl8DpraQkZudj5L/Bbj38ZtY919/k+cByteuzjv3Qkl
ucUVVqid8FM/PKtjstZB3+hzUFLrb1tMOz+9H8HdFUNgWZe0+3YMT9h1BHY8YN8B
saKvgLobH1vQKix8zsawg9PzeQ6EPua23U33/OrDlkd0UPbbPQx8H6ScHE3ReH47
6yxibwUCmXt73i0S/nazqJLh8ZN3iAvc6cd4CO3XlwWwV7NdrSVF4RgrpOwbX0Ji
WyiLzGv4VvXxoW/ymIp5VsabbRmav3u1ME4FIjAdAM+0oLVM0aMjqlfatfsET79J
3AmxxN8PAO1f893oxQimpuy1TFuT9KxqUy4oBos188JQLgw5JJO1Iv0AYDjsMAfl
ih9InzkSeP/2aGn/po9WEotC/9o38jFAJFKVR8rTVbXujL5qKZYoGuLAhSbw9n61
f/HyHTXKu/YryLjAoB+MAQDLH8hnkqQ1//NgJo/IVFjmcKu7gjpjG+fuOcWj0+f+
FzsbfOrQGIjJUjqnkLSNwQwcZpIx7SHcPdE+B17ApOd1U9hzYiRKHSdzJ3eBdchg
A73X2X9LqimdTdn3YnJGrXeL/j1RtOUmr3m5U+vKP/ck4R44oD6dPitJ21mHR+8q
8SFo1R4iJ+6vKLyDx6lPc149K05uAuLVD75aooMKgPyHQT3qtowIad2RDkEmzRJE
jVkxC0qf/z1BKoSvXx6/EXRWHAI8XDnl44x9DS6WcEmcdf2zVCQTpsObFjXL6WJ/
Y7krMo0hhB+KXl1ZK7r+ZTU1ElUx6MNBTlMU477wi7SrjYNau3vyWZsP8AwWipqK
kXk+ZX6bLRBmYcWSPXVp9Ui4yI+IpnbQPNVGgYnHHP9Im8xzGOz1trj5U64CQ0ss
jFw4GvyqASiLGlRMVstI8B4c+NHcWxrrzpqzRZ8I4ruqs05Q4pXE817oazcYJw2G
aqS1R/6VZ4DzoSWiFfu3KAsY2DhZy3pfeeZeZ7kCUn7z6YgSGlymXC0YouCghX2t
tFiMi9bwQHgGT5NWN3ldGpd9L5+m/sDxQsoo9g5ix9KN8xIaxDu3hcmZfsQhIxhX
kW7XV064M7yTQRxKJ1yhgztszHdsVz6maHO4LevbFMPUTH1u4bduumJGXzW19o7R
MABukuU5wT7VzP4rKSzOEx5Vq0akoIYQ6mWZxJsDx/W4jEbp3IPE3zxY4RBaIcfM
BeN0/DT70rsISpL5QXLXQce8rJlTXptP0K6WtCymD4Yx6ldQU1rMHqxa/ATMYGrn
nUwdmsA7qOpxHev0rYNa+lJKZo5WwAJtgUSfks8hEBjDejD39emxJ4DSD88pWdaL
CoZPFNOG6Nicb5Sz7PghyvxkschXaht7DiPXuTqdngnwhUn8vBZydxVZavET0wQi
KfqDg3ZjS3cCPEhTtZ5ZqIuSQeaY5lZSj1TILCROIegs6AjjSJxSi5VoakxZJ4V8
Xxd0OV2t6jzTxC2PADpXAiNc2xTnvItZ7DH0QVLSckK5AeRhWG68OvK7UpTTt2S2
MIpKS6nOu+TsQmxAVdE4MpH1MGPm0HhRPVcf1W7dk+3lVzqNXvDru59H1xVLOTSA
PzKlUUlmxMC1Z+Tg8IZapjZCbzGAP9c/AKgB9CYt1FzmfDhNo5DEN8+EomgSEVaP
ChiszqTrKpautredYTL0Y/AJwdhLm0djjIDrtVVuRjDvRJ25sKWKiLB1//jAD2Be
/RIeqprk+Qew2evoZp9oZ4d5POa9/MH20hMeoLqr4fXVBN1HkDGZr/5Bo8QED3M2
ryPS1TK7s4ILwzZFQpVoB36Plvj4l7VUclM8xTfpoH1SERY4N8wmusOfF6mlIpAq
EUWgm5ikkMD0xgC1Xq2tazYPdKwK9Y65xBlARqre96wchNyP7iONHJsKuhMFf7b1
Fv7CENtNuoN8JPFD9YOnRTJwN3P7ZF2Qi4tPBFziQARIdIqnkW1FLxUD3tZOdMJx
im0vjcjJaC1SjnMu1whEk+ngUj4LOjt7Kxxmu4YgaoNvN/unOn7ehMnyFRducHwV
w6krqJ0BHu8wIGw1v/t54YhDXdkZzJBL/PrWiKQeNYnbZTBorhQjKEkYlbsWqc6k
paAw4LzDN9ZUIKISCNoWi29+FJiYXdrx5uJwcSttoDSz7iXgLFaOZ0fGRyBb1Rlx
qYIA4dwGwrw1VTJCeEKwmxdduFkleVVax3H7GT5ssmXfKWefnjhb95kaB8vftxT7
nH2vwxLZGxqksI/hP+8Da5g1qUiyIxm4REgRJPLRYfeUSr1xWdrFSKl/Ujfqo3sC
G4rgBSOOGHUWyQ78WrxH0SqlVgs+bqD34vYKFFQBNsYgUyYdcvI1bL71cZI14XtG
aDhPyIdzUM8gG88VKbwafvMu+EWP2P/e4RS3owUZ8nVW2FWqySELrDkfKWqWr2XR
t6O9GmfR8DDXML11JZtbeWKB/CnFA+NNbNS+W+s0hRGb3D/OV3Xwg/KCgkW12j5Q
XEbWb6wgt57B7vHQhu0rn/uHQSxGzgTgKUzRMVqM02PtYQLJTmUzUIM5/TJOGT2C
MCRg57VBxOy4cyXgZwXSYof7VR8ZEj1p3Wo0/V8+3kInz4HfANEpZNpQo39svaBt
CjRk5WWRObVFFOVzhgoF5/N21okgux0LYE7MWTzwyXZL/Y9IEF82CzM1ipzv2Xp9
ny1BzcnmRMTSLqLucXkNjKYcqaJu5+MsN4OLdZShjVpm5jlZMx57QY9HnN5fclea
KFyV1B+BXU1h3wLZK3ZD4U9ufPY3zRKd/8wyyxZEJwx3IEIfWt9e2l4zSe5NjoU1
Pcv9WgQ7jVna0WW+HUCB3nWWyIBli6XjHCKthEnGgPhVP0Y1J+Ou6bwAr3l/nAHf
itSOZzaW8GaJWUutSo6ruPcRhJk9MJl2SrKwjtwTXRLqnbkqI00bg9NyVmd45RnJ
/Fm6bRTy3IjjUOraAuo/qB2fWXXS7jMq3QxsMvRm/PJW8AkZZwDolrl3WYQFc9yn
B/8D17xDjd00YWXhdoyCd3y33cbgMmlys+uMuOpO8i4EYe0W6w/3Jio/cuYYAl8A
XDKkcevmTkiHHq0eTkiyNTJ+xSYBsshqFOL4HVEoctRqoAEvuOrDtuOE8as+AvYA
TCWipASzGBxB6ENPl/a3ki8IdICQphMMf3yNjtwhxJmEwx7mCXIc8DJbVxsPyf1x
ZehpHnRZKIqsvMRyhIBB7UscfA+l4BudCDMXisy1oVpp0Ukx8Xojs0c8OVxKkyn0
sVz5y04e6V5SoK98ZhWW8EoVg45O7IDZuS2ZcQsq0Qull7qupLFWQ3L+blTOyd68
nIdkLNVVVIAMaDesJBrUvDqGBuGkCoj4NMJgNMvwyAr6W0mXejYQHvDYCjl4/gud
bPZuQ4z1Yj3c1Ai2bTYlLDu5kTtZD7cD1J+hm1agbbTxHG2cJyb4jkIqA7eImdII
pIyYfCK7O6e5OgKq7UHrD2ToQCAucR7MUh7varnao0HFGvLlI0aIEUA6xOH8WmEx
/S2mwC+6vtkr2Zoi5FmF51xbblWBnhDdkWsqgPL0+pFywlJoSXqCbpYHAk4LSGOg
vm5T6I9MmOrglir3VA6Id5/2c459VF4TjtkhBzUS4gxSmRlrAJ4d7HlW+3+jjNC2
EJSpGo/UC7voeFOQQDzN6uIYZzdkPqWs3kXncsao1dp8WnoN/3KwaI+vzVJIpW4v
87jf34elP/R9vBy8MXoC5z8WByBvcIhdbcELCso9wDfw+2ACWqk5wNh+VKFv0EWD
9D8OvgPaLxAV0fVgvmvl6ARIxjdp5JK48FMGcwUqJBW4i5s6RS9r8ty3OyAh6j13
IypOyjSE2+O+trGAqiSGHXWh6NCFlZYwZQJ8gblSv7O7RF3bJHbWkL7wBxyddVkw
DiM4JbMGZom2LcoJuuZp1rRhVNMpgYV68KPGAqM95zyK/KiRfaN9KaqVbAPiHgjY
pDCCQmVEe2/o8C8nYDvKNwxRFTO6fsupogywpHuVdgF3XfpGnbriPMIxDGYqngqz
naKtwMxYiOhnBOzRBNxTgjTzWX+J7qk0fo+J6Db7EB0GH9rxjqE72+eSeG9ryrZM
Tv0WXYgsfS1wqDtrv1kELnrH6tVhuXewpB4wwACF4J7D/fmSb+4VG8nkcq0/OACW
5RfrNpnhm5WWJdSyhA/SnhPK8YIQlhj8VV7WrMOWZYXcVR0FOtJICWaP1s82GIAr
+Ocrx52AAID4JBqY3VPYy2Kb/NhLbpIB0P4iuOWVZLfR9/Ecz2vhdvtIHd/JCkqA
49KFJLc5QcmBZdZha6Jyt8VN/1jliKMjCSXopo59U2rBx5RMRudFp+cAhGk3s5Zd
7VSO4YA6n6Dbd7NJP2HjB/f1qaiL2lRp6nkVqMGDvBjJ38EcWtPLuwVZaVPmr61A
gGg05VS8Wo+/3fcNcwITKaOfqN/a+XhEr57kqyhJSAgErieQja1G12r/nrZKW3g7
cnD4Xr/x8sQ6OqKdKQqyV56PQt7JzlgKQVIJNrkEciKqdZjcDZ/uskTmtUa2tIg8
uC4Ko0SUPLYUMOW+6YPd8dAjYjwMAG3NzSTesaOP9XN3a/5blq5+QBMJgUysELdj
CNALTYPTfQIjbCv+Z9o/FBGki7tPCOuxHvodBUpCOKy1iSIFOMLdGRa6PUXR8Ch8
J2l8WTPdR8dH1z5Meo80qKuVr8fy0ai5FnmKaOs5pr0E6v7H9zz/ybptONMe/NNV
9ngDiujkV03ocSHfsNzCPdDfdQabZztPElSf/tgotjD9ZnepbY9RkN4i2s3ZiBSe
qRFwSX3/xsvGJhQq9EZYoaPu7exDDkSRB8BlDZ1czNE26ZC5HTvZLeIJutGviLGR
gkl8YARaPVFploDPFctjMcpIodpl/TTidQdx/CU3zBFfGPiBXhVZjZpSwnnABshy
0YeHqlFhhcfSV7SulebbP9NZnVxbxAhiNz49NlQ/X8HpjziTZQRSVgbhmwa1Eyrx
Q1VTwKkN3jc9XBY7MZk10rQk6hCi8goVE+BvIY1OUhvmNOCrSeEH5QW7+fkTZRiU
gqbgrD/UKyhsJsRJ2XVvp0Hnuoss8Pwvc/DyU1pjOT/rhbDJvZ5Xy+qOcwKeLXGD
pfswntdR9DQpdZ6e1VvBqHJtTp7NfXVBrH6I9qHNdfQNqr5u5ZRve3BliIatgN/t
VzXFeBtJLcinLFgeeg6Tuupj8GGz+l9cCQSvCa0h58FF7VE932peWRlWzLiNq1Us
pj42Vz8u/+A/VFyylMI/iGtpCFy5FBF3HusWpg9NP8eNQpYsM3/3BD+2L9dnVokz
of76xWD9espWKEFuRNAeCiUgXkGiAfgjMXJvF0cZ77mSjYHTu22vpFMhGR0H0RTS
bu1J04K0IH0jP4Gh2+40Q6b50wrgCWWVczKRku4gNo7cFppLEMklp4DkebM2hT32
A1sXklDPG0Y5Alap0bY49j3gLnWYyAYgO1PYYUSS+/piMaTfynFKHcKWIQ0DhljF
jn6m5j5JG+yUgVAjZvGaw15ii+/b8G7bmjr9Nc2QSnG8RSFRZdfj7fNYBMd4SGll
zQZQLRZ4YP5h376iMyiNQt4qTDvkXkxtNBX0RbuBPgHk+Q5UhyoWpk/bsUtrvkXZ
YvQtwQvvHsovq2IfHCGVMtTeWUjaxKGldtOUQ8Ejqi75DnPOShVCQ+4mYnlqlqI1
N+m1oTT2peCR/DncGx4oJQzxrvLxuYqlgZ64GEH+K2Dt0lekf2bljWE/ysty+9eC
89lAq54dpt84ZGQXMK8zHCrRpIXiU6FtjAZm/Q0AlLtQjQcLtGmCIbONgXduI4EY
4Y4niT27wsXsXPEuhxuNXqqkCiytHtrSD9OwBBkA6NpWksIIyxsHORjBpiyzNfTW
snJO3eYkqiVvOvzD2SoEKKedtF3XHf+ROCtViTYCs3bAMYrMpZS3G9SctDUKihe4
36wX/mtQ5ElFG6DQ9jdQMoUJIn9eAqcb7lD3hE50ntLiu+EdZWkoYSu40pkCVka3
l2sbDFHAP3WI+3nIa2ZU5la9Qmt8DGn6p6NEmGCOnEtkc0z3cpB+6wKVr5OLo7ld
VVs+xf3K3ZWtB4/FPYhSPMqLOdSaoI/Or5rk4KANQmD8fdtDTM2kUNlmJymfhS05
GwqFglhy2twQjnYCCggkHf9/j7JSiLds1FqGqBVm1UB0w/lgZULdp+muGo1Hx/6J
ttXfI9xfQrGGHde+DMA+chQuVKHraz0cSx0bptf7NSox2tRMuvsI5gPwjXzL3eFR
kRuSIIQ53lj64wJfrjJ7RSa6Mc/HTpNLRnya0XwaHAaED7KEf9ZTUCq0ZI+9p8if
M3wStMDB+YOR83Y4vDJq6lfmIxbLXbqPD0Qgq9BKJB349S3VMrsCqVsKQrZg4zB5
lEL0lPmZqqp/FojrdZh7ba5id7pY69oenHj2BbuDqsnj4+KCWUo68B+qQMiBvrys
xu3up1C5W+w7yhSeUUunjvoR80TEU7xPxxagNefd13cH9xHzhNxikVdOIrA9I7Aa
FtK2Eq2F9kG+o4x2jbtGIJJ0qe0aDn3p+9ERwRsJH6NOjYidk105S0Q/KVktU2e9
7Te5lpLsKpRlpaMT65D5zhUwHvkJ5clti5wsF4tRfm4Z/3BQ5baV+yfOLnHDWz1z
m04tpUBzmUjk8H2wzlUFLbx1nmwewfSMKFSVEGuwQQiYs/MekzvcrAFxDOF1R0VS
0ccoC8RhtnRuFRR4yzXtr1XijQa/l1wyBD47pTUu8l0DXsxjUbs4bPN94lUugwdP
3N9RSiFnrnsGABwAUNx9qINex8fg8kdnSlGWa8/CVRnvoUDPZw9mqLwRknPTFLQ6
opZsptN1FGAmVfG9BorWAHx7T8b+g00eve1yDqw/LppH1UxYSV/TB9cHyms2ZZxN
w7q5o3oklc1VAVvXlu4hX+XZDNjuPzMkfXtYG0iPa5bdmJeWR6IRbbMoagv8cEci
9dqcSf3va3detvWdD+poh1MO7NJtXE6bz9dqaeO/OARrCUWDKK65Q/g8aqyjlTnO
2PemGdPT3Zn9DNF/FfVIaehwTWnsL9sYkces1EzDSKwMdlX7QsvaObEiooC3x1Tc
LXp2XpmkpU/hqPPUd9sb288U81mVccItjWEMIwN1Qgq91aEGQpdtBiW2FLf/zqC9
p2WJC758AfS1wUgj/TdHs4aT8E6OlCYVn0tsOrFEayLcWCewq4ac0YfbKNHrUM4t
LDYmA1FEytEqu4fWA+K9yTHib6tJQcedxDoXZKRl9+pi6TfFoubczi0O8SCiYT5t
s+cHpX09T0NNsNF3VFEiRALW/exA8pKK77sY3UqwUbuGzhEd71dx0pEAirgTjfun
+rGw0V6Yzmbbj406URqoNE0m5lvhFlFy8BSQTxGXLZv+32R8tdo71Pd2A2Ls8Wxb
D6FtxlC+wAFGqSKqzFoBJNAF7kqYHevRhINTNBkpxKJRfWw0ZNS+YQdKZsFUFr0I
M4v4JYyxyc/b1Fmb8xk0G0K+nY+I2pFHkojnWpFpTh35+HFTjZsFxPH8Qh93v1Fb
5KfsCQiW+MHFihu4FAZhrcrETjBB8GdvppqHg7ORG2LNZbQ9EQ5uTpd790pxPx6Z
NwoAbqGbI9i/4hnTgOGplnhugay76kUv28qpx9hv3rQCUCLR7hsyTHG5KSMFlQJ5
zlDyETS6UgECSs3DVl3QbUg2azhXNLVAgQK91b+SGcyA4KrxPDkpehIbObxe5pkK
RMKo3KTaS2TpaYCeXqOsLhDQMk+LhgtH9NZaX0ESQHr4TvBDLsi/u6kglmXFaSEZ
3lyEceZW9QgI79JKh5x61RNfXz4rgsbQ82PoSsgN3AyFgR7QQ3MkbVeTmGkVjkOv
9+KEUvEVU9kZfOon9YVQ+1kNbksK9vm94JNwOgS26ySBKi2H9vsHedUUFcJ8xzvf
CtpRuF/rWz00lmvrc0HzueWN16CWqYALBInIPM0nSc4tzB+turtUtuThOFGldJ1c
CQ79LFu/xuFH4Mvk3+lGdrVP5r4UZUjeLh3j+H0jbJN24UJlHcbeztmTCwwItE7v
jn9LnWwSDfbdc1eOE/eXUdpsylIAeX53bo84Kp32/4BDJyxQ9ChWHWWfH6S2A0Qc
21idmZs2vwwDknWPTnkrccCKI+Xy0sGeJbgE6+0TfWers1bojWiE0m/hpybGmkgB
g1KFWDpVumofpG5qd2doLfpf05sBC58TU+03MPzb+/t1CC9VCH23vf9yHtAWPXWR
KGurvqRk4+VPI9a/GM1bIUkat9M26zuWiMNMcNfwg4AdUJPST9jc8Hw2ukoH7Ohn
g19G+w3qU3/siyprHjDq9uNlcz1p4YxzZlkgWIasKUVS57x7+OzqCPFxlDz70vwz
WqMJ3BcKhVGwk1ahWSdsd2UDzqTBr+pjtG+GiUX4UAqVbMddGbGXAjbJk3g0dGyc
Zj3EKuMiH2vQHMQYY24M8bUFSvSDuhpw1hKzg3+rejSfY5AIS7NvDa0eZlrTmXJH
a+aeh2f6XrxYSiOUNnQjZfDVOV1MT8/Jc4WM/CiFS9qbJPCCwPyB3U28QFgWHiaX
xnwluCzdxIchU9jt5LEw9nLf2HKmLY8/npM+YC29HLGCk/yE9pzDBczUAiElADjf
Y7AjGCm1qvdX7Iui8FWmvofrRoAea8xnkY0mbHoGZR+jyO7nYHvLlvA4rGo6n5mn
7y05gLflLIAwmnrKMN0O5qGY10PArQbUu0GuQiIeCkxrad1dZ/4mc/rhMNOEg517
kaLnPhNvny+GBb+1VIdWhTG8vwaE16+6s1XvtGxHx5Gp/kbp2Li6XHjSxHlm5bFZ
569bRSNiUkJX8kpNyz1J5OQu5SvtsHOt+kqgzpepCR+1F1x5UAOJSM07fa+kfuvb
SvRCnl6EEyMrO+qH39hsWPZ+xKEZK3cunaShFovGgJplzKPxtFIzpJtZQKcYxDTu
ubuvxopfr/TnY+TGr6a8kKqDDz4J4I2SrX1llsWJgvH14SCi9MqTD3EJ1RjYnb34
N9X9sVeAE9XdF4q/MBNeP27HQCPIXZA6rMT44iAVpThG9umNlgSFm+JD+tk93KmQ
fx/mF47ccO6A/TSULOSQJB8mST8G2CaNkYWmV34IIujk3RGDPbDopYgyYw1/sCp9
hAlthnON1LVv8EfUw5vWPK5xgOWO3YdxptGlxDrulQhvQ1kCgGyeXbtwliBkh30v
KzjXXqj+Q1GRfxNxh5pWdmX0IAzCoTpjsStq2x/4EkociqI4mA3AAMLBx0b8LPAx
Oa4B7W01kFBBqnSrY9L03WVL3Zfd184OcFRk0SAxMaAGgy1VAJKIZYkXzKBji7Y/
dkMCF5ETdEPW5KFZP3m+tw==
`pragma protect end_protected
