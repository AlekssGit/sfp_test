// send_cmd_pcie.v

// Generated using ACDS version 21.4 67

`timescale 1 ps / 1 ps
module send_cmd_pcie (
		input  wire        clk,                  //        clock.clk
		input  wire        rst_n,                //        reset.reset_n
		input  wire        avalon_mm_read,       // avalon_slave.read
		input  wire        avalon_mm_write,      //             .write
		input  wire [15:0] avalon_mm_addr,       //             .address
		input  wire [31:0] avalon_mm_write_data, //             .writedata
		output wire [31:0] avalon_mm_read_data,  //             .readdata
		output wire        avalon_mm_rd_valid,   //             .readdatavalid
		output wire [5:0]  start_ram_addr,       // send_control.start_ram_addr
		output wire        send_cmd              //             .signal
	);

	avalon_mm_slave send_cmd_pcie (
		.clk                  (clk),                  //   input,   width = 1,        clock.clk
		.rst_n                (rst_n),                //   input,   width = 1,        reset.reset_n
		.avalon_mm_read       (avalon_mm_read),       //   input,   width = 1, avalon_slave.read
		.avalon_mm_write      (avalon_mm_write),      //   input,   width = 1,             .write
		.avalon_mm_addr       (avalon_mm_addr),       //   input,  width = 16,             .address
		.avalon_mm_write_data (avalon_mm_write_data), //   input,  width = 32,             .writedata
		.avalon_mm_read_data  (avalon_mm_read_data),  //  output,  width = 32,             .readdata
		.avalon_mm_rd_valid   (avalon_mm_rd_valid),   //  output,   width = 1,             .readdatavalid
		.start_ram_addr       (start_ram_addr),       //  output,   width = 6, send_control.start_ram_addr
		.send_cmd             (send_cmd)              //  output,   width = 1,             .signal
	);

endmodule
