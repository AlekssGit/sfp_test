`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
pNifBhXtxGdLLmsOZGrHlnRuIRqe7hhQmz0ZpZDomHi/0Edmw67w+xyU3cwrZftg
HRfdfaW23o09FEw7XBeB3WRtw9o73CE5PwArFPOkMTmkZBRATM6yywgtorO5hLC2
QnCM8Sm2kWGd8XgG5NMeQI0xUEK0Pfo6BHfC0RJCBzA=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 31712), data_block
kVEwGak761BMbyZeBFDx+J1famk+pWUXKvwqIjxWAhPNMxTMIPZpaXqYS4YHtLvT
qkWQCYhd8iH9g/cCCkyz+HcE8PRZV1aQ3vWU6BaM3mdumUevlo2CMf6ixxzRRod0
jBsfFK87VRYHKAemoQaaBGA/zIlEbLp7VGhBlqbqOH8BlurR1jbqAf0qTh4gQV0v
NEZVJK70QI8kfA3dnvtbQ99W9GK8LMR4XxVraDUysqlQaUzGibqcjZ/lfWTO17cS
AFbXoqkI962yGWtWgqGAH/LiLALKdERuM7Mb3sOj1XkG/+KmwkGjrCpL3U/1ogm9
aY9lJQBDAVusldZXDkZMEOmud4Txd1gjgURnRWJEpJXL1TCMAkG271fq/019/CmO
WfyBBttoRaeCiXupcYRXLslwp5C1yLGuki9sT30cmoEVoC++cGiEsuLi9xQ/dx0f
eOlNgelyYyqvbfQeMHCX5bI2KHdgfAKUOAd+5LwzfgQW/nG1AUxINY9K9Xii/3TY
KWvunMspQJDreVrDEw6QdHH2+ypLoIrY181HjYmGnnq59GN9agIp7b3lhUyAxaRV
q1sJhfFdI1XyeDmEr7o8RenDyza6xP4PVxycYJs48PKkPq2LLxJImg/64dPYEomE
ROMXmEz8vs4qBB01KJ6kQB0gFKHALQsptgkSmoRWjJwaKjCpl4NIB83s2EhsSndl
pvOMXG6ftEzujlUSuRzMo6TpVifduiJxNI+aL00yh3IuhyE7vjZN5uCJJoJ3v52i
43Y+gimOPX78LoUrDyrg4nRln8Hslofm16kMJTMG6ghaIQZI/ZHWLugVeV3Gkcuc
n03vGMN+eAZt1r84wp73xJbcc7pCQsVjss2jAogYcT6lAjL3QJjI7I4aU7HKpBE2
EdE2RkaJTanQhGmfefW6ZzmiwceYrr/tgy7meH9cXs/TtZGRsiNHG40HJfW/IvaS
hw6BFDMuiAYPp9TxuskK1JMmjHLwRB919BD5v7szIyp7vxiVzJYyhFSuIPGPOsm8
zUXEchrCg8RzzeqUu5RWfIF2vfyJ3r+r9cxvRhqeKYWwVQU3w+DgQ6SeP7lyGPId
C7u1KQJpkdY9NsZWBhtUDdBmOA1q+M9ZX7Y9P2sjM0OmwU8Gqgqh0fL57n6/d9yq
e8mZ+K4WDeZbFSpKpKHnEKew6IS3chU1vWP1u+Xft5yJnKufZPiT1tsC7PT6t3H/
Sx1x85ooPIRBSsdHFfEuz7lartdqhGgShz+0XHRuI6+uG4rjQ7egh+1fiTDHRa/g
vu2rD4Td7CrDh9Zh4X9OEMnG67fX6RwXH1Rs6DcMGRvjlqurRi4kFEMtrix/h58f
MbWhitOYXgVp+bLddWOG0CUdpGC7HSRwyrYFwnENgj/TCpBcQjMBQcAweHJJWSS4
C1mhV3F1LGTjJmxLC9ECR0CMPy31xlp5jUuGfYzRwg80nbe3OwR06ARoxIgUHkwh
Y8EVfvBRjLbvFRWu4G4HuJhneTboN9/brzSpBramb6XHy3NO2XTaHMFSXWuaedS+
Au00iSPn3mDm2BgHaAeAAhvHoo2w1MsbKVIRVq0C6Owol5d+CJoDX0AsAmF85pLs
/VqxbK3CipLgR4orH4jzU7KpTkuOBLQmNfoeWi2rsKTowq+dsohidTR7fTu5kNzs
CVZ2SaWmRILf5xZBldVdp7NfIRQJzHhIr8fd1DO4lrhVxNKyfRu5CY+ogfgdN2Cv
2MiWO5JWdSaYpj4Z5m+uou5ui9009iIn6fuINETTyfzoyqaxDF64ulbQFKTXrBga
Tc5inf3LPAtYZe3d+4+GJGjR9bemILhktjiT8zlp900Si5w7Eed+kmoFX0HGhDwC
ET4vaAFPEGgqJg5z63sZ4KFcci45+rHvVdcI+HJT5zLI9ZUCLRbdw+kmR/az7xsv
GtN4sC75j64/Cp+oq708bvcv3dIwesiQ5bpiAEyhLu31L3YOYDOpsEozg+Y2BzM8
wf4CGlwKHfwZD9RYNiwHzVNjFwMFdTrmIoE5gldoI0x9oHNzbNlSZrzxNnWrvsO+
hMzj2u9EHaho1BjG6d1nVYkia4VjErh9fq0ZRS2azMdxgKt8dU/eBwc0mNIx1IGH
9UmM7uHf3UlUbP80hqfPexE4rhfaBXOq59wq2mB4iuK0KFiAxTc3Whr7/ismm05I
+qdmkRbRQEAoW8yfxzIJZohPPGG1HlMSO6CT6I+Ostb4xcgVdZyxJJlPSkf+HvXn
XV1Za5N5EaojI0fvoBWaDIyLoHD5CvMebSAhiGxWMuiCtCs7YTlvJjBLRaUVLCeR
mEe2BdYwwvwx00haAwNXViWuY8QXwdNibwT1VvrUn97fVf42JJXWXdWJcrYr7I5u
cjgbrL9VYhobXds/KzTSJP2hH4yw8JoSjzghhelB58rOREybDvP61hz4TxXHdWlB
17NiU8xkFHiiMNPA0W2R3bSKkBskLdE+O4liCFO91gWxtaeeVnPmiy0SMAi3cs8V
LFd8vJKwGLeOrfP0UV+aWeEa8UtDSu0OtvpV8suHUKzI+8p5bvnHBsBxHq/hof41
YS0L1wF6JBQ4+pYuXHPJRHHmdPSzSJbHXZ58unfQU0R8pcnOjml8ylabP9/aYxUB
rjA/4yOY6SkM9oFiQycWmJzCJGe3Zn8P7iNonLjT7YDYBq5ljMLYnOrrt2a3Eg6D
szbc7DnY77rRdKqn5PDlz/SPmxTFtaS8PApMnazplvXujYl+TbjDZXa5/rmNZj3A
jOSyQxKdF4jigz9oZWGVfrvNi3toCtxxhW0ik5MDGt+ZgILpOedcMnaHb6/w/D+I
/6gtQKnj3HMSxHEh6WuwkhS/M24jRWZ9BsXJKm0pMXPZNBhzC/XOwhOSIrk4HSda
RrI7sA3ke2spMv2rKsDgPce83P7YtwwEUILu7L1NgkTmiPafWqeqwHCOxEB8xfn9
hLjlsQmwcj01i4xhzsdcdlYfCuPhbjR5ZA2GZ0Msstuv7auQx/sd0w2T/9Pr2U9G
ZCJ8q0DwvX2FXg5s/Esyn0DbCCkUtW1mBHs5w5n3jyawZdvTMASi8lL32Z3Y4YuW
7Gmu3U+Z3YmJWUbJxpK8/Z6DtOCn/Ki3KuC1AXl2XKcyukhBZ4Ioj8Lf7QdyhjFO
2yRvg7TBmzCqtngbK0MidUAEujArEGySktA/YVD+F21pNInm6ooieTgDrXtxGTNV
BJTBdOEyJb3cHtP6BEZczah+ltuO0QNkKCwKNGkq1HLb8h0Xqd6SRkZhpef4Aw0D
/ePkTp/ZpqMHJfGOdJsb4L6ub+v0pjJr3chFamMld+Zt/r3drn1OECPK+Wu5D8Yz
dGgEEkxq4zWsHA2rhARxRWaPdBuhI+gLMhKC5yiHp/UoQqOyNZIDHk61ypmQr/4s
qWpDXoXH0RJrPQ55wYxZW3uJKOJ7lVmzwhMy964womuyhagaASA98gUjsuSDLzXB
HMRttMwBsacDR+7ZbQC+tdqSaBUiht5FQsSUOCH1kLz90Yqw4xe89Y9k7n+5nabl
zgXGObRiwKDwq4dOPJz91a+sE63IMTKT/WiTAHrxr6NvGqfnOx7fUkdWtpfxmS/D
aPXUFdJHB1YzecJDi5QU78bhsom4sukRXjPzPAd8kQeq0eMSKHjciOypRK5bEx5V
fyN4kIIDFsZvCqpfV2CA1Obl3RQBaEGX0hqoV4j7Cz/709x6/8qjo5VZVniq8/My
QDvlrOD+pO07mxLTBYfqtlFySoJ0g5RucRs2g6WuRMyAbcxlJQjO3L5SQr9mWZIu
H8tkGv7v+nDijpPwGcFaS1HtWdAjf0f/dlFh33bh/j/QDgLa0KHPwt9iQwcviZGB
DCCGLVWziCMzZLmN94VOWmOj6B9YvYfT/Rcok8Fl6lxjyptuEnY6lwTfd01+hRWB
7hMSO8y1Mxtcg2nHPaPVKUt53oQ01zMzC0lbtDSAdFA8LqlI+WGBP6F73IqcVxAr
LLzy6Ktt0JJpfn2Ed3v/HZLDfyxYKHubuCyvBPWjH+tLXSaB1qFSSCrfjpLeE3RR
p2tvX+TSN7v8KQ7a6xuqBF3szM2RkZqQvZdIm5P72gsk3qRJZUcXo1bo1tucsjNg
rq1eYfMQsadYDz+jPGrOPKmB3kcAl8hQ2RV1pGzcGM4iikrCvnjUlKgDdbx1D2Gn
lXYPdPU6X3VXtJVpKYLH0ZT0sdt5Z48VCTORIHBVbL3ZUuo+1/I31XfQSNej4srC
bHa+ANjIIHbmefiXADuppfZKpTKs6zdsbYU5wHAFqo3AqmVcHOjIycmi3sFUNFva
Bi+p5rLqPJUkFvOqcioTDf/lzJW2dmejlXao1Pgu7a3LfqVoK0w2oZ3cbYgibw19
xsNKRXlhDP/rn2Cc2w3YiAndc8I3B1M/orgbFz7tvsiCyFTVaJYmke6k7f1v9S9o
sIpOPde7AbM8dsZVb1eRlXTR9Z6XM3/ycoi+jS8PzSqxQ2ZNA0lNIsdNRO4h9//c
2phRv9s2Qz9vqVphwlnPHV1+6icOo0QdoGMOgRsSvvRFSSFO/w+VUg1aPQXENeKS
PX8Cn65o7x9flSddTxjzWfGSrrrPz21W5lPs4smwMNi7BNHxgnBxRVzH16r4mlGf
U/hAiIhogI/q+WnFO11cOvNN/m9UmwZoyS/R7KwPUL1nkbe31vYxw5gLosUqAHqr
xKolPX5Ci123bADEqpU3dsQcN6JhHQsbjtHqat0OI8c7iaAqROckWu4AGrqN1GV0
GpcLHmYeCS7dlofuqU63nMZVg6akGRRdlhmpOPdeDv6tvwluBX+4YwXco/IuSW1T
8u1a1kcoCJQwaRVmoCWr+qqPsTzQgdcOY+TuPBo0Z69QDJjZ6WcB7ul+PQPykIQt
Cuu51GSlPPKbe0uJocgnRUesnFyKM17e4Nqf0xVtoGZZt1D1QUgcVo0KGOU6EXun
CdH9K/60awASk87S8GBCj4EvQcxTtNJUQLSxkd3CekWFcjfnzU9VY9Glrsd/yujf
GYOF+SOvWJqvhA1NqT6ZHgv5jy6Wr7FLoXf7bsDXys5cHtNyd0FzBijJBJ8cjlSA
dHiIKvTgYnKzDw8ysYck4ZK+G5NO/enecmbHhJm2Hi/r/On2Mta4mIizddZRR8Wk
3+onSAtwCD9DNQbdn2g7Eh1jv3DbWelAP+hq1SmTZz8ZypyHc/XLvYh1k9YeNtn9
GtDyuqJf1wa9pUISvfZlJCdqdLKUMsiuHqGT9yqJyoj5nfODTX37xCSCMck0EGNx
2uV+uTWlLP8JawY7CygeaK3D95NY5XgDUAk2277ytQ2fqMzKjRgX8sSWuY8BViIr
anNITHiOI3H9TDhw8kd4Qnu60DHCh6Cml6UrmkKwG1TtxL2W+qZrxKBpIm3Lfnq/
y7VJCY1zzXgZ4JbM0ZnsqRgw/ZUQnzxCk85lIlj8zGhUen2twNtkAXD8xi6HdiaY
6TjOh7weZ0WUZYBKaUpCj8tnVjz+4ndNFaTKAKoRgA+1XR1p80AIvAu6OTlup1zR
0KMnvN1LbuWZE11tBVbzOzCFojS5LHDuXB6fyiZZAH8bh0YKQVm8uZNNlESjj9zt
PI7ObWe1VEoCrMx94H0ivyOo9vqz4i2/FhTqtnfQuyIy1yNBNAWVk38xpX7JDpD8
S1w8POG1FrcxaEuho7NdpszlQKMIhCyYKY7cq1a/5nct31vBb7SaSBK5bAq3yFq0
oQ5NRgFRHE1rdH6hvn8gtYrCIMa6LWBbxKE63r563ilGjr36UdhYpgYuVBOCbO1a
kqo/7XmAMTw+5Aw0l8Se6jb8cyQQpY1K1wmiX946qvOBupLz5f4Mgdtjog0Zqw97
eIibxvweovzp3ASw5YN061hN1gjHnzYo23ho1xSPt94zQwyr7q/uZAlMA4irvWqE
emi9hqsXuBTxW4mgXTu4LVyF90+UZRVKNEBxM/huLRykGY6jQeYzgAZ207aUtjnm
XtqNOKr4p4Nc256cB3Kj68EwFrYbCYb3iZx96tuUuI4ErWtLlhpHQnpkqhwe8fu6
UspKnbCJLM4l22flRz4wp+w+qamOUy0nQV2c+1ps4JRlkTkpfH0q/E13ulY3ntr9
HqMl6g4SUn1IxQH9wELfFKY/M7LRoEfcobgIJuivnyXTlyU8ZPOKatvFRleLo0ZS
wT7vAwk9heh38OKyAtBNhrUGGitoCdn1UTZxtwlkwdYN8+2/OFQmFbOwQskiTJA8
2tzBhYIkZ+MU2y8Lv3iH/DfE9FqB8p669FEDnR1OULag5mOzxzg1oG3Sqqcj7QUQ
GL3aHO8XDHJbkyzUgmcvSxaCmQ7pS58xwcIZTC8ahAKT8JdvFKwE1DgJflx+XhKG
tsXQJ/W7wO7Ilm2IqbREypILvteu0eyUIf4HZwNyREN5JwbflXVloKpZvSeqq2Zv
CpoSajOhDHCwXtwpn9bgxRx7RNVNANq2nzraZcLV0XIwufHP6WkNCtACIBtEN4HS
D1qs6WNMLzee3zg+FpjZqyg0N0E22n9KGwua3dfudMoa/bnIspry5kSrEhrPyiQZ
qgB+cU5jC7zArKdPP5rR+/bhYbWYtFIa0jPw3fSE8rXJesAYda1euHpQNs3D/YpE
1vULFiL2AzOHVraTzEbF7bExiy/TLzRCS/aaLqXaiKSpNnrPYNVobWM6K1UszxiT
QJHOpYBOUcrbzDAnNen1jHZ7ISQldEh5gjokEXFDgiJzW0qf1PDCkyULNPljnc/d
HlOl/SEYFsf108x1K/+sydN2X6AohwyxOKxCNegbcouHJPKUoBtsyK1IgTXTDaYb
tdgAnZNPlMmM391tVrfyHJeR54JFNpEK8tTEURLolAcaE3hwUqcyZ5aRWIzZM8+P
UfhrgwCbsDg6yuGKyPbNcAreh/xI58ybzVJKiyxoyYJm9Lc+nljqcKB+m0Zofu78
DVv3v9Z2/5rz18Ld62pAK0RHNqdMocKhjmDOu7OvELX/UZ+fpjMEd47xYE1ZBHIH
ViREx6s0/AeMXiavihLIH+9FtlNjDsO1UMNjoeB1zKptnbW/rkKWDcz9xTCa+UoZ
aRDGw9BQ5RrUoLKoy0H92GdntwC+r7WO8lSuhaOWfaageGoF/360dO3Ko5+DiiUs
AkCQFMVuKpHWXM37J0hu4XIqrlYsDjT9Gcl7Q3djYn3JkKiZsPDtPI6nYNf39CqJ
CX4uerMGuft4omIP3iOH6VEA435142UwF80LWWbtHbTixu07Iq/so8EHY2dptvNU
K1hTrdqP+7AvfPNoQp5qmnTy85vSRSKGmo/8TJ09LZMejY6szn5gWzWJvnYIP8jz
qflbM00npi2FSPwrtuhXyUo4FAnLDo94YFdoZ1ewy4flS1BVMOO4vVulf4rUlQgC
D8I3zu+zlKfpsgmiy7/tqhHc0oAD5zFvBdFeWIUZnuuZd/BOUbQ9ZLC2cZEAiX7X
SiHhpyd4QaC2Xy8qRrdT7YJ7VbYcb/oFH8HvJEX8Kk3S8zTd6wuwtDm3ygVBsDjg
n19ni87Rnbj0tjX7zvZz7k467DlrBnhg7MezKQxLMDx4aHTPrr7saFgjiU4dZTaa
Jskvrc44qSsVQu3QqGtOfZHtmMAep7zDM+rjYiSkpszR144W2r9+6QLBTMLlC8ra
kYPpJeH8h2Fc9TFrZAk4urXj9WDvoB94Q5mwv3jT5FReSKdwLZqakBRx1RnkG/fP
vhUESp72iZy92ot12gJcNJdyHsyIB0QMSqmoa52qYXPXq+xma9EQfdipZRp4JnpO
T1QnzeZzaNBMfQ/U0Tc98tLNNlLnYwQrB+j0OzOlUfZmsGcLzml6zfRDRk2wknOk
A8JoFmeM3+N3x8vQcKvrfb83JpZ+i4shNwPMOJhng0EsrEPv+0pwm2JFuI34b20o
9lEslrXda+L9zcguzEzGIlzHBCStE6F5qQE7On9Ar8Ueq6CqyQ81QOlLX6YF8VRs
EgYv9uz7dYgccxJzLEqoEYLBENIK/MYLyJREMShjOKTCF1oL/FA04vGRbU/WJY/w
abnts+146Fjh7kyaCfUtZmtsmSdKSKVOfHBDjPfdgKgcGV8PdzaptQmRI5FSNcmq
rtnrtXvlIHn8sQOcdMAo1A9O5qaGHeZ1Gxx83WTVyeceGjHqfwZY2nlon2OPGKX5
1MqtGBGzhfxG5eaJCKv0CwFOHCz8Xac1vVBqe63x9KnbFe7c10NKgXNY8NTQJmLn
iXk5Nq6uPk+Bb4dRzWok1KAQrQZmdsDaHbCaoPLOcFzLYAae48sfBfMwwvFZoFaX
9pjZ2hRY1ASNwzQInrmYQFK36LY1TUvMSWOmLwCn7o0cRN5tBXAioOT0cy4ZFaSS
TNY73Df7odz1xj/UtagKgnC5IkgRklCDdKzzEQDRekc5cbrw5QzTy6jr1CQeC6Uk
JnoJyOHV8mrJPvo/QiU7K1ToVuWf0YCJ7VjI5MMIU+wohmeSEdV1dhvbJuu04IUL
w9bFQutQjHv0+x+lhds2Ea6cjVE52XeD+nJi0kUaA4OqypaJCfxUabUlnt3cuith
xY8LVlMS8sTYKB51+arFR834BCM8uq3LEJ5u4/15M0tBAfvHBo3pMmk0ASoDpbny
Sh+MbzCnXde7QsNqhTpySZ9eLWJ42/DOEWRoY+YSSkEyAwuYZV28yghXvRF9uyn9
AWbT3rDqv1c0nyBv0PyusJLoUI7LK3yyIDOYxJKayn478wQH6FxhYJDpzAsYWV0R
ddTwqwNgRu2p/OUR7WQn23YUSPFey+pX0SHUXrGpacugliA2IMiVTcBjdDzM+Nab
hc/A6T2jcyYn6cNHW6ocQT2uV+82VjztD4wHZYuPgSvlrUTD3CxSthfe8/8vW4CJ
e9/wNR+SyXQwTxydJVJSir9QOXB7RgA+QSnMosboEpfaj96IaNyx7wDELfTYn+UN
U+RF5qRN4sauwsar32pegwy/AaIKh+ItlnVTvqoIZLvqj14KAmymONTwo+WqxML3
qHsDXtjBy8eOcCoTxnNTmr4roQOydjHyNBlelEHlpLOTzy+lnoGc/PEqm+ELy9MU
Q7vLbrRPIGIlkW0EKvgBCXmX9aiC1XxK0+rjqP6BUk7PG4w5RJfNzLfBxDzNB+sE
65+s6QmqOqcQNyTNFxPWaCDdtyqz9oSvDFeP3EUQCrXF7r/re4tdTtPr5lGhx9nI
J5LLDVq02UKeTFkxkWhxzPT4KcfLIAW00bQvLqZ3bj+LOHJKP5abB9WBFERBURI0
nls6n+fsHA9YSnGVLhxs8g0xuw/ANjdVaQOR9xjjG+0PuRp6AAAJr2JsnLQB+NUW
my9vZQ/5U/oVWRgcDwGoYhyczHi8o6vuPSHESB9Psa/+O+fJ3TU2kscXjWcGklR6
8lHd61v2WeoVUL7d+CxpHxBuokKBnSz/6dOcIjZiGx5aHTMxTK+2+z1cFir19kPU
Tf9o9Vs9Ew3b9mqo5Al2FxotpskrgLSttnaxJWWGFAfGZY9Ys/VRM/yPgyuqUTB6
Xd+7YB7cyIYcN7d2AqxFdp/oOBTAcaEg2HnHRsWjwcmRupb2A21WIkB8Z5NNwFvd
tBt/G30A561040UmOZf4qp0a68IiXin1StrE1Peqwt0mtHQQzLK7VWHMqBgit2Cm
UHtwq2Z7Y7jjGsEyRZr/H2a40QNYzVLGeHb9QKeEXw3WLiotg3wEv/pfwckC2tjH
3atCQP2unH2ynLv2Dfk5+q0lNEN7tJKu9hdnszhuGiwe9/nf5010Z1YotsJC5fhc
NnznnochvVetLgQHcSJ3uTKFUf7d099C+lzAIXvjj9KCxryUTlp0T2HMI8sXt8jA
jl9mr9bF8G6uMIt7ge3Or8RkGk9w4N+Xgu33RT74fJPpw8TsKE6P/xnIqmHI6vdS
Lh/gPo3wby1GzP00DpYrX3YdECOzDxBt5+o1A1YrGCjRAkBraXrDwk2CuXLgkytY
H1AqCebUNpS6hpuGYl65ssQtkFObunmt3x3YwiGuLBWZIV5sPLYF4VwEI44DnpxM
VikLscJGKjzoDIxRx8x9j2IwhvCuaydRtvlwETzzU3dq5inRaM7ZEJWZjCMsOQXR
isAVd2aoVMcrsk/LXRQIF5WKbn6fRf/xYwHE8237TEIhcj5CIXxSB3Ku3edswd3Z
wo0+091vpTBi791ZE3lv37IgUObqE1HE3UWJJQDSLVqXwDt7eqKb0sOrwoRhz0RN
oVOesV4Ib5HQT8aVzmsmmvuAS87Elensk+01iOYFSHYJGyMdbkLqLB2+VziJG5AL
Ku32XrNJ8PJPHCBHRbiVUsvjx3kXhWzzj7jyREV+wf8TpyOuOwVNX1LkFdQzRDZe
75VEXLhJG03t/+2pnr1q0Un0MRRj6/1NAa/p8pKqk6a+rC1TbGmxQHMBYO5X1uLq
PHS0lJ30EY5zjPHBnTO0r8/e2L6GCmmIV1zqajSni9RfP5il4EUpUgor8odOpL4w
Nfz+o1h8WqzMM9j9xka24h5c5azCBknk+wW3kIEQnq95fqRJNy6bEIqF4TRg56y2
JvnulkMfHNV9yXkdi11hTg7X0ba00ZKnwbm+jMrvqFPSq1TdlFMeQYl+lPWJvQo+
D44nfcz/jsUiNNSq0QTbVCuT/R7mLTN01vkrs7+X9n+bIzAvEMvN9UR9Ivqe6XQL
/Ic26xv3QKJ6W/0y5FWfeWuFdF/CG80yU2mbPNP8hnzLboiNSxS9NaFXZjFxo4Fw
xpemIHE9xgSAIgSvGSJQpDJ932O5vcobwPlmZdi2qSeZjL5gWroAAxq7Dvmxeuv8
dZAdZuUre3x8bWwB6gzkgCErFL559jEsvWb5OypDG7Of5Zd67MXggeIwuqzHg+cr
IKYKoRvUMXJ3SgkfXmlsilq9XdX0F/DukLEo2rumvEorWm2tZ5XmYixQQYTs+hi0
VPiC5TQ/aEh7pmMsZIseTVk4ZEgFJN1f7nTjhkXtok89+amH09ubKX1dywneyQoJ
zJkgaD96h5SV1rVsO7Qy10d2zOE4zZ5OzDaZZClrRAg9uTZq6pmKnxvofDiP/j0S
Rc1wEdnVWzzvc9aHSg+2FkDgwvQ1CH2qDd7ZbPM3LvVhnzio7T+XEb5+Pqi6m1ZQ
QKrGhtDJvPUM4jH8I0/KQq/z43Nu41eOerPZnFQvOkQ2IrX9Pd5tkWcty0QwUiQq
R6JfJXcGgbf+CKSh9nfCSC5AL2MgHUjBugLfZYzDraLHCUGFa/w/vAv5XfrR6K3Z
9IwxkyGtCpjHzBA0gNGR+wgQHwORDaaoPfXnFxsPLJ6iCfN3tlDuIRk+iQfP7sjL
G+BCXvFAl78AxnRZL75RnQ1pvCeIYj88313OYPRKbEHoGm/pBoTX6CIQFoUoftl+
d8JA9Tuzcrf6R4ha350gVgkrtQ+YTzKej5nlUsH+T4FCJjcbEJLdPh6U2MOnXE77
5jUCneWsBMf2Qw6Lml9vjHfkmPJ37aG+s5ItY+mA6H+I8xzhLGQ0hhdeCnC9EhMM
Lu2ZK5Hclow5qvk/02YQNToSy2Uw08vdUIUxASiIcEMyKmg9LS2bTx6iK9XMWc2n
pHCyOVzRopMHwOaFykHd2sdFfps3MDD293R9e0z+WgUJP4rZvGESXICTFvN7ERx/
n/ebGr/C5PaKGCE5WJ8SWZhGez8/pKTsE/XdrL+87DlsZIrir6yvdHGrWHy0//M0
zEx9y/yNlG37vo94D55VXa4gpZ0pVVQOwqt0aFzeZilElo42UVuLf3tDoGLS3nfQ
HK8/v4G3jNQmkk7N/bK3rHVYTS3xBbbmFa0HH4LQbJAVDmBdXJwMjCEUGf4k7i5j
IC6ZGaeuMrROQ++o3cXGypzMmQOKphtky/yWPD2F6V2lOgeSuRWRgzio8wKp6bvj
IqZrm0ZHqk9DL/741xBi3yhcimTXIQmVL+GfChA9Fkng3BVEwEjikK4uziR7nqxd
p+crOjO92wcZjOe36ked7S6Ij5HwT1RuhhIIFNhZPMiatVST8Ogi1L2HkgyulIMb
nb02PedGNAEGO3ADmlnanltFTtjSwW8Lo4XoQaez6oCluXCRNTWLy5auUq+l0Qny
dq1fXdT39/QGzknWps68Bp9comZQvppQIlVP2eQdcL713uScT/GoF5oXw/NwVBQ4
QJB31hyBwMOgijEyBfJhAbHsxuAJc940DSJOube9nxRKbloLP7LG7AF3X4y4Nw/M
pepXsmdFbphZxJ+B2vSHuCXnkzqPzP78iTlvCb843kPh2u9SK0DypJnPclhA1DQp
Li5cV6gHeaXiT3BmeYZa+TlovlpTDuReJLkkeskMocQ4r7SbV7ZHJeFhxcg29Yip
ZDBTaabt1Q0yASLYgJ3VvCps9C1lBkCCdLCajFAM64c0voKZ9k0iUAsHnkf6swMv
yyORmSp9xvXBnBbTRAsFOLnDNHqs04z7UgqH4fe8qw1TVXZ//N47dVNYkcIkCeqw
s3pFqxeq7YzGa77/joNHlEaOFF28o3+/JjW0vTcDlMBmAMWyotH0d8Gy+Ep43WAm
os6ncBIrRp11A2ABsEVxB+AnqE6ZD8A+stV7xHYWkDdtuLzOi2zA166lhDQgop+H
perwYVh94xP12J/EBJ+XPXo/AnC6dG4Jf8DpuyznWtiseRxY5IZLq5aYziUmUvmX
xV+SMQt+t/7iNydgrosLxe+7q60W65japo9047+Kr9apG4ss3W4IdKcBimRPZCx4
+KYjfQHE7sZX3D8/3q4fcvRYKeFque+AMpsJkuecpQ0OFqjwB/AZmZI0PXfZekNv
3afe86ppEZo0XN41uSrZBUUjoi129mORgl/rB0GcItQEBXLq5H7M1MXQH0TT9cNu
GBQb8rlwLDSTqPgKTxW5nP4EkV+V3Kfll0vVyEtEwxUwM5MiG+7oKG869U1PJWgm
vuqYXPRbmWF+kk9JFlLMWXwCBk35XC4/ToG33QTfFlXbIJFJU8Xu2bjmPN7oa1BD
9I1zItJkLeXZ/N4OL1M6X26HyStGj7pQXhww4iAvVMM8JwixWVIuG5ZCAgeSJ9Za
rQfLY9k7tLTVR13Uj2OLdYlrCUMZe3xK9eYdVsj0jHA10YxfQS8i3zqe2/mSdsVi
8CNxZL4+9K0JMSOYwLsTNWTLfnWyKNI7lXzvzlSEI4IWGY54hgoNVAciDDuypgHM
QeMsFAr+N+bitpOXquY8LPge7P99iKB3WtgdDaz26cFgZMAfwxIFpjpP7+/fCJ18
zZ7A116fS3ZAe813PuDwcWVWOQzr3gYUrl1+UBzsjepOprb4jUDoYK/Z0t++1o+O
ni8pN1mWHkjeT+qV3PbTn1BKkKEfz6nZn78VwyXYd4VFVAU6A9ckm3q10mJbKVP8
bVeBxQ4vOnFbcZR1vGJLIseZb576/Y8oqscU47h9+JXwutNtqnQaMtEKtCnVsRE4
My2eR9nrfHDv4b7mr/yF56UaZx6qy+pLebL1t1h1L2CjBmgHzM0yEUVg8pZOsPLU
STji5xrat2Q+A3frZF1WxE/UPKxD2SsNsxWbv1bc1t5SZuc+UHZ1QHyk0tmNMFOX
K6a6BfCfWIHphZTuhWBsKzgrmv8YA3IdCMBlOQKExuJHEvZAVYCJUKjOQs3d6Kee
CBxfV7/GuXfQ9DZePEFl9dcHY13uTpwGERsdDDvQKjJPgTq4APdC2nyUyymS/U6A
IUcTD/MlHV4oQYID38TAcxpQyNwR5fCUFxBekrKXsrY5GzBUNyqb4ydGzL1UiaBX
sY7TBVw7QIrIAoeeDnntKTm04qBDlGt+HRgRWZac0ZHuxBazfjHXncUsY7JbciCA
TwIAdmomgpGTfgRcxwucHheSjsH9Eo9vodtRm0HBf2HS2bEVUKmAgMimAsKDRTGn
iudVbTIuqaZfTk+Yh5iZ0bD9w+BX7CIwQCJAcIPxaybykg9UCw4kUint8YEMlvfR
4r9woN+yrGymVL4U2gJ3ZD0IIVz2mJEso9vHWzN5iR1y49G+CwUZcEQZp2BqT2pk
eduQkXqlJLYrhL7kWTQqH8pz39jUYXWuVLsSO7GeaRTM8fTqPc1/ki1gtt9500im
ni3937iYW6EGNOLScuUAQXu+YhPjujgBw619Wni7Ux4MVSna/tHA57oF62vnU69/
XlPMr8UR2EJ2GGvsDMAW938ef/p1rmQM9wepbO2MTCNwBnyLFcE+mKyQt9vb4Jnk
vFlM2jxaOJKK63+zdg2bvJBFcclQypAmY55fdspUN3SXtT/4xqtNwHZd/PBsdzzg
amR7ClQjH58bQFqf3g82p9ts9VFkcxIy3wZ6yFD2W5b2i0eeFzSaVmphv4dkecNj
JcHSGZQo+o01OTqvZjoHO3+1inOkwfXUNTJ0yquOCmOjZgWaqwwjQuHggw5+aZ5a
KlH0zAm01/xNADrboYEwpwzRkFJ4aredEZNiQ2d26LBuKLNn27iHcF92vl7CoYrd
cvkJhPtzpX8V0qv7rqSGj2fdi/90ct1UM0f+9bphqQx8RmtQm1cuIfJOZr5J9vjs
TTADtNM8g8S5gJPeb9Fe1KlBfblinENHl7I6iMnUvkJ2PVobUxJ/77SbOmrvw9bP
oZ+JE4Odn07zimplZn19FdQZTwMemdocVdDhtAMU/D0+yDd3drtc6NgW6f+QN3rM
rxjBh3AqfHDOkpjaLoLAcpv8eokK1iFBNaTdFeWFIKwKLuByv80UzvncoOwUuJrV
XO+sM4aPdhyGIt0ZS8Y6KdFrj1UowGGWBLKuhZ27dmLaNGMTYQzmimi4ulxzVxhG
N5Ki2u/ff1FHqupwP1gSz7iBbjj45ts7bNe4A7CWIEp0aF/ddsP5gQ+QuFZ614+m
azgENTzAgiBG2toPvMFlHnAdxEBYANH+hrbo85UzNamkh5M+v56B+57T9eTwb2M3
f6nhUyoPNQGfgpTeO8tTKWJKWcksh7mvpEWl14sRYWxQN34zkYFl9kSMlvnwnURj
M5v7bw+lcCo9+qb1VDIM60He77UXlOJ+iG4LnrZ1siCr0heif7GxERyV3NKOUxnq
5tIMPwFINIEkahE6neuGaOpy9Sz+SDQfts/keXjKzOSfYtMz4v5eUtwTRyZyy3EL
QJHYMhLzoqhGlenCBBCcA0QZ09PPTfujB593A4lA2RtQp4RD8KwNYThILJom3zct
I+vXXpqL9mXp+R9ieb7cHws+qM0vT9ICvaferW6wbzCxKhfbc04P07ilHzMq2gvS
/Ygy3dPsoOB1rPL4fZqurRvLPSjHBVdsOw0J5zmjlBMAl7QNbEUe8bhf0aGa1zMC
3Hx8mh0fonmpo/CFs1I8FGE5Bxesfn5sFlqlc8EiUruQdwMLsEY+NdQxNxvMWoUN
e2sGbUfLjwxwplUt4gBZ1/hALUlwN3mi5MEQ7VvSXpzriXrDziLoAJD+KpbMNMcm
lAhkGsyfGMJbJRa081nY+kS27lgZs2zkIIYleUY39wAxGMLO2CZKdQeQiaatWYd7
QKNTsckaG7cMNYGDrq33rbtodrr2+rnNWbjRO+PGexQXJZtwd6giicfLBD62556R
3lJuhriWTKhDl2yXALW+bT+KID7QnEbrPR67/4hcbDfbF3i2nASoH/5g25UquboI
fYwDzLcnRtlUSKb70xk5UdzgtKc/IJKgT1+/ynwdocvkunYTfU7UH/z4iLVkiIh5
Xad+fuJlDLd4EDhOFFO4vlrppHsmqNfbh/6yDBjcJLPrjSdo0u6AvNp8X4omJAsN
01IvMYDBKTSogYqzuA34Gr+2OEdvTpKRuOAkkmYpqiChuysrMJFBrO36aEIhb5hr
EvEpxjwFvql6uvIoVwrucBZKLzhUBdDcajmm0reyd1NGiVpYyiwZZ8EYWikVN5KZ
3xkWSq7Ysb543MXLyx1KKc8iPp95z7+8kJE7SDqWy+ORdbvYXRDdwMk1DZeY1DbB
GoQLABr55Musm34xwa3UTTxYnlkX5DKj/aHyOreZzv7xvSFmTGlb9zgUWEHDAMGn
JRRqB0HrBlU6+yse7/tW/64MhAKM73D+2YtGcCNUG+k8S7kqs6wRjvfRDVhXOmB8
amz/2ujGavzV/WneeaOh2iy6lewArVnzBoIN5oWUuAVa5+hHba3Soe8YiSdjD2uZ
F52Tzgp+vgXK5eVp4meL1F0hK4g4M3ToZf4yzXih7o4D0ZtO8+OsZI8vrgEOqllb
RIA3DKMvwkllF5MEMJ1RzNawOZbCqA5QHnkLK+RJK03lD6qUFyNuam53bxS8D8TK
hKoNKd1sTVDiXKntF8Ebhf/9xPhJVOd6aDOKEtT54EF+jLn1C+7SOflqW5s8A8Y1
QsrZoFzNXj1Qc2fs/96ODxvunMx0Nkr97Jygb1bUIeR6Vz1gSod69fPdKHnJgFrm
rKFeBYhp2wE+zkR3sljf3lydhEXLy9acavqibqFdnCQzoAHyCUg5fXVQslJUz/qk
Yi4kqo34wfELvTs0cOD44oWrc+NEgXl6jVkTeemIlwfqtPxVgG8IFSoCaSZAq8KP
szo82hWt49kJqixdxI1mxU6n5fQtbO058l7Mn8bfbwmxwAi84HaEflmM4UVft9IK
/lvJn8q3TAdzYFr/TBjLS+FffYFWrM8hJO8mLevw75qDbNmR0fdMBbGOd+XkohXx
redF9VcoaJgZYwauIulIngRMEp2m7UsYQsanGwG48x1uqBXPphISYBxF1IppHrga
kRYipC65SvV4cp7+tDtIjGr2+WI3v+jxNVb4VnOucpBPNkrsjtKZfkNTbGeKR5p3
jmZAs2YnmO+fdiaMcwaNVjw3qLld2LgUb+QsgYtHad18gASKWNZUo2zWaqtTMNno
YPwtdy0rulmrfjL9vrqnomA4WuGHbm6XqrigL99NXVqAKKrwbiDTe3n5Y1yhQk2X
GwjRCJhdH1o5Jl8wEwLyFx25y45Y9PUfPh3YsEk87to4xtFXvKb0De4ehEfF0pfD
2I2tnUlL/1U0ZigBUg4IyXasBrVaPPuUfTcvD24Bveum6tUBYXnKZTkIkz8XD+rJ
1wGoscFLg1wb91N/TVgEdb+7B3i7Nmt/NOyH83AG5Fn1scMBNUjdWjnXU1rmuNEW
2EFCInEqM+3IL7bcQ6AhicHBGjGZs+WTAiZTbmOy0z/dnjcyRaQk1ySikMfs83sV
J5IPQogBvcADSsZO//OvMw+0caxvWS1Li15czmK7EnAgpJMbuZJ+9q/pD3NJDwxm
MTCTG+GGpRY5rLCKQualVHcxDlRyqnPKS0Z5aguuXuOKlwLNf/70E5Khr+GJedgR
oOO3NqMH1CTqu+OfWEYIAEIV8kYZdKuWVBarI3HwTHLFAhh5tzpvHZQSMjP67hQi
5V5FiJqDAvbBkSJsA3yrIIau7SuY19fjzReyf02tcs41W08INotLgKzikp4jv3qL
d+ZFfjigNOkve2SUVs8W/xUCgAN4N6uF4LlWp4LRQc+UDvEjdNJfYq6+eEWy1FnR
lAdCi0lR4YvwhTAP9QZPMlkT58jE8NBCFkPYA1hGYUnSAY5Hl7HznuFgz1NWeGnw
nrOlaEkmSOOup2sOaHCSWwaX9h1729OtPCMZA7N8hCZIByVuaEUSmNKce+BcPBbU
fdQda8x/VGlXtWCbjFtxrfL+XNhSD6lEfjTsExupY4hHuQCfA2JwGv/sARW3TVTq
5eYTUyxslrT8Bi2k9H68HJTlvXpNvt2wnzBEW/1Np1mgEFemx6NEveNjUsaa/Uz/
Xn8FXI8AJf7+Ql4LAeQD1++qn4tXHpYCdGXmB+0BkoDOidlSF+FeJz8gTAxSmG0Q
/s016A1VVvI1Mz6WbJk5CcpUeL49wsp7paH81X+CkT6HW/M15vkD97QNPgX8RHc0
nTRvA11Qo59QJSNeTKtPl+RXJkDParLaYQUPdMU4eia4O2T+yti/SdFWOSdtFd0S
khL4x5hl1H1baHE1MXMSKBjv0VCF5XUD1ymefsRodqOCqCMDeqKDCoOGT113aKbm
0ggZhTS+cVDgqMbssevAV5kmXW4/6ERx6RlvInMNe0ZK/+dSZKlyGQy7PhMS7AaX
DKIGJsO51bXLHwD1mTuou2C++62cgkGYaD/joJQGiQfyX+walQX3nffY5roYBO+9
/OOcMgQJjqGDJM9qPa/KkJqcB+YTbuMJMAfxsSh5kTjYtkl8LiyqE3KwYxUjVXgW
B+v5Pomm6OD9YDX9cu3sslcahNmefTzNiGLC3LaA1ZHKCGy12Z/Wki8HNWoD7uL9
hrVAkOvGVtikgS+bpT5OJOw+XX3DJQkfwsCL/Vj8Uk6l80ohwHiZ3vnIU0iraDHB
cOLHV+Oa1dm5Um/empIr6HlZjvRJdbSLhmgd6sA0m89qffDEk7SzwxC05e5UIkeg
AyYYgrZINiE68I2MCRjx66/UFLLeUFzYqjcMRAQn7aa/HIXS6EekXfc9iqObapmC
QhvnFhmJmWRUnsrFlKl4JVObZG9GOoJ0EeHVfVeAVzeIw2zn4tGV2J5G7M3saVDe
QOwRsM7uHtYBqYfsWS3URZpjG2ryMi00DAG5KFc7NN6LoI3WTS4G3W3SgoI+kN0C
R+qP1JkXQBC7aLCJiXbLkYirV2lXiE2s99MLeF0U33gpmnAauwdaud212FC8J7DK
14VezTnjWSP6b48NzfjDYKQhWiTBdUm6AmFvYqXvuxEis98CiZr6LRHgnDUrf6m8
fJ9A3+GtIApDbycHaWdLcI4zzydD7eOSbMGucva7im3nuY3c7bGMNSWPUQ+wpn0K
z3+1Sib0YCUtcS0LQtzIoNqY9uHwyPfBH9j8YobBtt9fgvRJuluTgm5e96Kjvz0Z
pgmi8dZd0TW1rYx5rTKpEIten4jH/IFr2eOHtsC4hx6+1SNcyca+lOb4v82UlAD6
RtnnyIbSaPl0kPu/9UAOWVaoLdd31GgV3c6ZzISDZeARfgGxPc0aZGcrxkJmhBG5
iwWjzkk3fQm9GUYHnkPxGQkm4OmT2eSgdwVwIWCyNHye7g6TzUgp31OvY+5R4KdY
O+m7W5lVO9oW/lL0XpVwY6Ng3+Q4GUT1stJRqvlMfwwQT0a9LQ5IP+hJbbEh9q8z
uO0gNWPZZE86i3816mgLwzN7O6HAvST0k71pX1WZURpVLU1nCGosTFIUD9e+4JVk
ZOQKCypTqg6k4GuVOhzZYHrAIE9k5SmBMib6SC9Mx9ydPIk2V4yLmQaSBiSxLVRe
QT/mDc7LmNoYTM3Q0hqYAyxb/CXCBMOrCW/0KmTzIGvS2tkD1r4CNIdH6ET7PNza
s95sGXqCrTHhCbez7ZknFjMIm0micIef9xvSYZczrlHHfkOgASALViZ756vIn8+B
TCflbvbJeaUNwdW2hOF3zlbQqVqz4bpiV16w/WPEPn27L+PnMU9JSJezGQsfvaIO
eGg0bDzZSfr67GXjtpLDtIUfl62Kdq/d6K6p6TnHC8ICK8YUwv8zIpGgU367ievo
wzcXGappyabxiEcx6wv7uOWopEcZmRmSp5+hKMxJP8Fk2Tfaf5WPRXQv/RPmt5hh
oVWD4B18/1cl0fv7nPtvYg7L6kDvZjQHSIWTMm6H4sdk803rUVtr+9WyUik8gRgF
6q3LAUV57HW9ffjtBVtEvur5OUlaEhFpiYBJTf1iAK07a387RBx6mqprfU8zmhdR
VvKJiFO9h2wuGYjLarDxzUgXAwS1nHHNMlf/Zw9asEXMjhZT/TgkSyUQoKWs2EG3
tQLe0/QakwJpabu6CAOdg25a/gXA8rMA1ctue5ZzFDkWUdHDnVY7MWAxnZP3OZmF
EGMAL7Ow3Q/lh3ASgZcdnghtw1DObji9/CNS/cnRtZtk/RDy85AglSNCLZekMW3a
P6u+le9urZQ2j+unwmW3qST0XjoHKY9YqaYditpxkb57zbUDhrDpW9yuIH3VbarA
Ihc0sphRRb+sPqCEbdKpColEJq2TpG0z4yaxNysUeAFlcU4pbgTmw9wyQXFd1srh
HbCOJjH5HZwgNf4nH8/m/iH6S3+jJ7L/icgFMfeiuqGbWmlcSm76Qf1euMfCTX4F
1cmRlQBFKdJojolafWpKcX4T5KxbMxZt/UraFMp6lvI3kIowuDB0ZA59tB7i6inA
MVUdkQK7phcVuNrcSYwpQm/vvY8jv4nEEkUSKQNJWobFg02Xf2oEinm+N07YqlLR
zIlQx6BlgvnIRyNl8WsQhCrpSYlj1xHgyvA7FCloEbP2lkell0+ljzlPLvW6uWAJ
A+t0fhYyqf9yhWYGqi6O27chrDwZqCPggJiTonLHXL3tfNtR32MVVPmatgDbXry0
ExmQNyWlCazkG+lf+IrNKFtSQbja4V9ivR2oAYgE2zU/5AlJHsU6QsbjOjYJIN1a
L2cPTl4g+dBRpufeAfYCI1+QjToHI7EPSvNNUMCky41Gb4FgaDJuPHMkuKHHSKbp
A5lRjLgNHv5O2r5qvFgLhfltkV2zXFyll+IVPunOtJzHt/mvjB7hllsD8zoCFH0I
ylTgK8Zick5GJyRO8Rd9x7R/qnVNzK7laVkBtgFjXzAVj2j5Olr4YncVrTPU5CtY
18J/cPDziW4x+P79KO4U6lhUNIN8KnrmR1SL0Mxe8iizMYZSC668JDnQoQqqmit/
4u9nXg1k73aCwH/7RTUhsZIaMnAd6DXORg2sCmWEYIjZmOMPYpxMnglgdQbbHTxF
uB/BnHvDylb1opBSDJP8FwgDQnGZtlbZLKufG2wT0tOKoYuU8EsfwHzIGB+zhWgM
P6cd2zGXWN5H2lOkTwF4eSNv1p+1TNpbUy607ciXs1G0DAwB+idxIoHBjoe8Jql6
bXBPt4DpvpQHww8pNKLE0bRUYOIQZgxWeyU6ZjdlTmlBKdeYZPTk9AKkiAnbYskN
aG3s8GD/xFfhfdqe7EhR74BzGCBHpBh4NpVKp+tqDIEGtszIinymrxdIe+koMy/O
Xwxe/HBrKyYk9lLelBsFEguYKOb68w8FmDGVd+POf+vlGulMS7m3LYESF7xkXf5A
KFvME7f/KgFtzFQ5SM863ztoApDzScHizK2iSoNbe78WoExD22HhFcoqY76JBIrw
KR8/LD6JlsUlDzjY/wWHxGDwjd2xu4GPskR8lU6QsCpSMJ98UjGzG4QileywA0zE
ZSAbbFw7kSOcg++2eJ96041pLGajrUQb4u7LhJhS7apgt1kLOJ850koBAS9m4H2U
o6qR9Xxu3opbVWmtS1El+czxycya61ADRzlsWyXpwJPNuwNBUfiWhA5vEBts9+bf
eskvgpmuIVyoDfeQDtYZub8kRlodIDAGB6dadr/AWI8qV0u8QEMJG2KUdk8hQw8i
spao+syiaPfQ9bRI/y6XBoin0tXwiOPnLT9zhXMiqZF50O7tgl/kVlJXipU7Vu6o
/Zn9k5E2QEqV8pqXrfq6S6yzKPkXP0kWgJ2pNv/6QH2BF+zN5+7PHwWZMx7jjzpq
Qc+ruDXgoUjC4ZrjNxBYhnIJpE2CvsdmGeEWKte0QGiLpxCMzgtnSY2OU3MoLx6V
ow86J5G7/+Q0f0xbJk3uabSuu+deio3Fjl06/bvVbFvu5ob/hid3ZiDZAQrcMVMA
aWGXWwCLs0/dXOqvw4nXsd8oGavvN3TdmR1poehvkUe9vBBRfIndusY1l5GJ2bAW
g9tlfRbuaAGk4oRSeEK7mUUWNfHUMHBHy22HOODWplktdQXFy8spP70bCnpSMlxK
GEtNO0f+V37NottlT8cBRBxHSox4kD5/pCnrIg7/lMM5zlYN4ZgGEzhFHSJcwKbW
Khm/BFz9vrlVMxTyc2tdzW6DVigTKXWdOfW8JE0AX28z1b5KNqNC3P/sxy2BHjQE
+7PkFRWYwzPfnCoOJEUeKcb3Qcw5akDk8FjE2cA2mUN/cdz/fBq0uIN3wp4clsbB
bKAlJ38+XTTkpnOd7Z6Shq4uXC23fICE5N+75IgnFSebuw75wZnjUM3dBD/0nsFn
jpvonHeIdJsKJNwywsz7BSdM6fKBxDcSuo7k7yPP96htJvF52DVlTflSgBjabTt/
/6aOp8UG5E5WYfbRTsnbQAFkvd5IDklpqJMslDVnV0u0EwcPz/CXShSHHMZCueFb
PY/ma3Hc4FMqT/38dGUdcRZEl6/BCW/QRCuZTjNvTQcSm8xMzFiYRyLRWkUDXQiD
n+WOvioWV0mIYXCrmUq8jI2a8+p+R8XTJNiMAghvTP30JSe+Rp+0A45SE827EaQi
8OJ60nMdcV4C+59/o/v0IbDoa1soYPswD2D8BrBz1V63e0mV/MwGrccn1iCenU9p
y54ojxYuT3i2zc3b0+QCcyRSgifqmNOSuIHDKui3VMB+DpVf7Y5IiyJ525nbbya7
8G+4rO1OkfGFncDUq9afYpUVTpL0araYDWzSaI7DmVdePYrQ/2EOEUB+mUfIjSsf
i6ipMaxuucO6bt6bQh1xwAEmJE5H+JVXVrwhTg2tAFMrlhQdCasj7nL0cF0pE5xD
CwhfQ6EldKTNebHTrQqO2FSNqtQthnFRwa0TH3wDYo0BYOf9xUAqUBjQ6eqdFQUY
T+opnTtTrPfbK/yB4lA65aQg37H7m4dbSSV9GlgmdFpZ+z/2BMVL8V6rc4NZx7Es
Pwn+ZbnK0kmfyXC4lvIJ2irSYQ/OcrkDIc1DDC6PmXaexfZFoxGfMhr1T3U7SUQV
9LhHeSaeF9kiySvoTLyEn/LP8StP07Nh2MnlTkEeLhmMx5f9NHeO/pq3OWEuLw3I
6Mdz2RClmQiYN8696ntqoxUasESEU5QWCgI/kNBHELBj/ez1Mg3/C0UvAmt5DTIZ
YvYG7/Wh7iHiuNSnpaQpCAFJ9sGgOcRGCYgMahGtWnwyElIl4kTLdK+HmLtt3bsy
OQd6gqzoKCBlfFucNf6WpCxOtx3Iya8ZUl+UrLS3h+gJCVA7t5cyOZZdsk5D0HUu
JyZR4BXk833wzZmLVwFFVhFKTY8eXatacP7klxPFdcliUK3nQwLR9uO8iZFOrEoA
EK/kMkLy09rYlNUskJsp9bysGkyNtxObomVZTbUXowghdueAvgtYAmWORmZKLXNO
BgcvxKp/ui6CGdc/7mN/DnDmBzC8xJ1URlA/CTc6bRnMBIhJeX8uS4ZH7au2KTCX
n4hVPhdIbs29Ppw3cIhspEA4fJ/Ob0L5VdYYGQ0sJIEe/Xf6WOEhstdWiF6gO2yv
mKnVnhkXmx+sUc9VTK1uCsaY5t1jFlrzVDNCyYp3K2awp/vhTbEbI79vL7Ma/wPJ
0tTr5pIEFKcTTN99y16bU3U6KkR3rLEae8ov3G50GE83Wqn0n3QjuL86rexJ4tUY
t5ytBgjqJBY4/8UVCWj0mxRc6Uvf00u0F8CORgtd8PCP7Cvr66glNaJINnxSCIxf
glPXY6iV9ZCLYQoeJdpniRA79A1Xya4qTeVtPnI5mwcoYP40XjkuxAe18E37/rRf
LDpw+dXFV7Fr/jteXEYvZ0VHp1J+eQwfhZHOFZonyXHZSw6sWJjf6yFUaYVDdDZe
wEglspvSvZWU8cJ5dyciiwYhYeLda9/b9UTbujkhVVogkB+t0EmOBi472UO4cc4L
bcdgUN3GWKEsV0kR3HXmRz5FUnMFp0KDykCrBZApyHb7JPnH/TCw6cXhuQ9x0irc
nShvMsujCIp1yFLq6J4ZYBbcNujKJI5ziCseZV3o3taEak6k6bheINkLBSGp6pCj
sBKqwl5oYIQQ/4fCAN8BYp3QSk4emBPpECyPUErrERSx5YQCJOoDvF9b0aMEnjLj
CEvGm7dSIM2OLl3LByiaRllDiVtJ6p0B7Xg8BmFjkRkQF4TzFVz8fbohdAa5Ncar
pQPRvfvsWvyYOztYxgZdUjdexXjKkR4c1Kg2/B/bXPpZOxehLb0KBpp4gNUhBR96
fS5akHMRVJpQB67KKOjIJsGTyMyfVpgd9dhkuS9iPhZc5rw3ztJBrxwlB+sRU4ga
HfMpHy7bopj6lTTRcOXd2cBvbUrpYXKIRVQoL78ocew+BKSI9oS02cwedXFDXX9z
eACaOosm+8pvOpEwE69aEF15vLxSi2A1I7x1UQQghPQ8DxxlzLUvNxXG74ebZGhd
F2UnnAwIs7LFMJTckB0ZceAg2sZ5a98myYpzg1dE8WpW5KaT1UUJoD+egqYEsWf5
TxjnsxEe6NIGhew4+P7yxg8T+ews/e7jut3Rdc9jVmeIKM28u8Qmu+6l5hRxMAIQ
hIBMLZWS7CBP6b1qcmU2/VNybhzn97VpeBRzlA8NgfiSAS4IMvUCpFjfrVOEWy67
wTtwbCO2pX82HjQ/LbGklB9N/IvNDhW03WyNeEmg78kP3wV80QTjDoHBT2ynBpQ5
D6ylQskMGdQf/+H0Ql8QF8DGCyf8GgoW2Z+sNiRQGMqIk+6HkxOVyvRZXQo16YHy
YE7eOqlR4BEalgtIUq/GWJPQMZkKRPZxzzdMSdyuPBIT8Xk0DvtFXV3ES/I80cqu
5GFzeT5EjlnPNEkUujCGMSJZS66vJiTuPubKD/Fed/f21URbN4oDKuAR6ZhrmOBW
XNmalTM0mq4/ycqEClis7rYVfcwJGLy2cQPb/K28Pnn8JOKtgOjHZQn7bDiTiwK8
Vq/aXy/iBkaNGFjLxM12lA3oOj05j6llP853PGEPproeRJlIUCxPUBPe9/bzO0+D
jSXCqMIbLpzDxWGjagHKwjNsVc1As4SmPRiM+N6f6mQVSF9NPk+18VDmriCKuQqH
5z/Se6ebMIdU8+38+ReMNhvudJvBKFJArZKBAmoNGDtxwV08KPMtgxf8GpxcCWj+
7PPjlGgxtqaQBWh3N/QkkARO5EFsGgUFCLFg/gNftVmLU6uw6WpQmfA4Y/Qpr9T+
f8YudBfIl9Mc0HmPyqmXwpg962E5dL+bxjrttZRl1BbnbdXup9Aff+hYgbmJPxzE
7YamBO9GunFliu2ZDR5L103CJqb73ItsTO3bok1gvxHn1TeYLkMNnLoDTKc7eIWE
EEb1QicZM3ZcscZC1zeJ4sfsYndH4zGLVWJqXKnOQTCokOpA/drTvubP8XLghbFL
yjpZ5TN4tO5TqGV8PoqPhAz1TvvqlepDl+kLOBdB1xl7d/Xx8ZYKV7fGC+bmDMkt
BiGCzYhF3A4KZwoOACMtWuKUD/mOAr2G0w3Jljrv6u2wFsdNl7HX3dvk89XDJzU9
S2azcP1eWCv4uSIo/9ckC2zpqpjM9tRhaeGqDK5iCK2AIGq4TzjfS8TLMYzbxD9O
oHe/mhKm10aa83lKKj6+2XPlopPRYAxiQVE/oi08Kk4/wO40Ru8HqoezRwzlOV0i
bdcQ3eOijvY1xTJIBhtqil/uOvVskkUavohqYjvpIa7tabwYpGOo0vdt+c52Znhi
JMqNcYGLsWSLvYsohGk31abnIg83NFMxT4Pvl8pHhjsD4O8bwRUQdKzazoD8NXjz
sN89zI90aPPOvUMU3iptgWkH7rmW6iNoIsBTKDoC27hmj7XdbbLK8jIi4eQI4cFc
NoLgcmDdJJOkaLWOO+Q7jofvjsye0iIMjgGWthTBsG+2hecXG2DsPTYZ3kGySmyW
E1t50pUxSZ8TDbXzXkJZgOZ8xz9cSqV546JkQXDkEQAXMQKlUgbYp543NEjHDmrL
bGb06ijld5Sw24BnjM1OTHQZIJd67ULxOJBYIL056A7payG+cIxjR1Y4iRWKZzwU
GFuGcBCgFNt1i/t392iMDzaVS6BXq4+MPvPUFTl2X/iU6+4pfvn588AjUuy/BH8l
NzJGbGzCZ1SExBTB21JhDFxZ/X+dXQ0YzPOjOKLDjAeGGvdRxn1VFIGgtf07UVY8
Fm+jAchCiT3lgLrrU0HuKSVkXT1wQEawlOeclGGsJtZYQo+V/eSOduM8BQM5kT4K
bkUv9PC2DHTmYEDxGMOxlRkcxD10UgO9Mm3tH8237cH2psDuTArrNuDEolK0jK6m
xLNbFyjNZQMF18p7yGeQ62VaACXVbHQwINfXT32HXg8xQXv96BB6jiZKjMtvAkNK
T1mM3jwsnwtJ6y6hn+21+Xdp7seyzgDiW8qvIJacie7To1eBLQqgGZ1z/yBQMeI4
43v7KocLw0Mp1MuEyDXX2bPpYL5tbAdTSxV/qTkca4j1RYQ43yXl/Ur5U1C1Htgr
ocOu8KppmcqWsbxaXXIaWQDIORy8fsQtUge4vVHVXkvfXPmb4DM95y/m2qegv4w5
MPYmFnhzfVgZAbR0WaDiVnWdVk+RChRNzRPJRXBzl8fwOQEWg5rBDkKxEk4QIpwY
+x1MD544wkso3JRIJrTTMXUIWM3pjTniE9DLb325MgPnXPzhgrizqupwe/MdgDmU
QNcyLRRiPsD6Y83a1pPDaEGNCVxW2uOtqkE97kHaWLl4rpNPuXWcQwumCI3qen2a
o/u9COlBASyPN8KcWmVE9EjzCiSWbpsfx6h5acScWeLN7h+QL6tfCdYPiszEvv6X
oDTvEcy8bKYr+mVOZLoAY/4juKRZUw6bUwu905VIbt94N9xdRzK2Mkcwzhvge9ch
2jkYwR4x0bG4C05Wz+9RoeRsuVXnVtwqdLlk5NuN21CDrZ3S1Cpg9ooPMuCavjCn
7r2hMaJbJI9npltC6GK9pYbi2ST2u1k140DLjh0QIORoLUJZgIt9pMaJGD0fQGkP
ugYIklOYgVOo3X53SFYQjxs9RXCxIrLRdtOa5yqZAFh9RoVAZBda5h/sQV4no12t
kCgEd9BAE7KhuknS9nHrUQjofxi7d/VzzyBqd7CoSdMZv0HT58Bwp0C1RfzAeohi
BMcRGgKPLz4WegR8ga1DKbIsfaDtT1zN79KIh4sYH0QLJin/b2FOkYEjbQ9WpaYA
EQNftoU4blnvPdjRYXK/Yt13obZo5dz9LPo+dfxOXnq8Joi2jhGTffu3TA3f4gKW
YgOE7d4hYgCeE8So0VJoXQQVGN5SvXqtSqfREVu8dizd6oj63HDobwG3hIlFcUG0
Zb8uNC+YeWHYz9aIPsbIJIJ0RA8GX51XGooJP6zulqYjd2YQYLU8dDR8a/+NwDE+
Dm1iVDAjyH8UJEIW5h7ZFWbAukn1Kr3pNuxptiGQym/DuKoUIqFaiRw7h6qCozCx
FxLsj0T727U0w96BTbutKkef74GDCd3ccLLwr5SwwjIDxTP/smZdP1uctirNaaVk
BqG0p9tkQ97YQHnoDzutFmdzoH9fxUDOeAAj8Qkir4RI3xcV3zt2fTm2IR8aL6zU
w6uBdExqVknI4HO4cYRgLtKgYWiSselyMCNLZPNlrq4uwS+8uh1Gu1y57BBqiyOh
SbmEdIyu5xi0CY0N1cmKIBsYfwEJv8nhxNEgWUloQrpeD/myL/LC9K7VtX7wPQn3
+uN9ztBP5+ljuIVQhIOFqbJTuDZLWaQl+Dqka3v+MJpf7pq8QgCbsFH3g3pQ4DGf
9Rfd6hkbztXwSb8qBFA+RigpFXmsraKfQb46p80TjVKNzU3EdkiIJz0Fx71oLrF/
Ppzn80U/a+hOPWuFwoXF9Ij1mi6+kDfhsKK2gHfAkEqDdEvM6MV1W7Hr458bIgx+
ONOOMCfFQb2IpD45U+vttskmXaQiCKTR6P321GLTvzZc3uVpi/cMGv0JsHJguxM8
fh2QW/Amn7lJa2R7HGJQtFgkq35B/Qcr9CtiRzlOr2xUnYE3hApM+Qk428rSAKNV
OIATQV64KTsd7Zo81mHCWE1CE7ShXow7YIAZEuRW8niCiJPUIXXIOTrA/xAPxYFw
M6BTDxtiZDeTKmRzGmn8zxEPRfWHJGduSySHSSfWMjYVk7MgFH8WhzzzSxngnMi2
xgHL9P/SKdwNS4x+bTLzFH51E/yUr0TEbDdYWrLJxmPX145Q/SCbZDWEvfTlqmSc
PMAF5yfWDje1uLTQyA0QEXXQY6+ZcqGfq40B48IWJ4fnJ4hNnszYorhsnyVim1U/
PT05rwpCFIoota0P8ukJQ/vYQBn171H2kejjvUpSzfBG34+bftiDhxC+Xcen3ZjW
RwR/WeqtFBykTr/kwcI6q8soZVDdRBlpXBMBqaCPoJRQAJfQbyE25WSltirByvve
TJ4feOimtiuIy7xE4YrsXFQ7Xe1h5cxPp8OL7EgQ5zFpLqEif1IT+zL0AgLDfe9+
eLGkWJ8RK03Bg5mVQhbjB2JdeCreA3atFIFEfqSpMPKcT8bvH6+j8pc6x44pkc53
UOk5LjWArReAjHu0u5l0V/E0nN+5ZIKAUO8QAxROJofRP3xzSNesgA38hY+r5ciL
JkrDVcmFWkO9KCco1smIyXF6c61rBDt3rA4NnW0BOHfUTr7VjEz7AmWHvpXzB5Nk
bUvVmbhKAEumjNcLyZMeJps/PXaPTxxC9GPRo5qCg+R2sqbRlOBJrwhrRvmEbZeY
8TNvTxO7BqbDNifa6jLj/Dvfdb+IE/wwEatuZlFIlyMurJS+C+KimXaE3Nadd5eH
sAaxNVQODwIaUZxjBJ1ksV7VxsWMqnRKxtLARNdCGIyJKBIHbI52DymT1IoqkCkf
uAJWsWvIxkWbsRU6JF9PMG/9/ANRigonJBq3dRnxUZaKyevyiAm/LlhFVAt7pU3Z
hgGK/2JQFI65f6+U1Dw5M2ioZ58mXNQ7z6zVOzvrdRKqB/NBv0XcCPzNEGz+87nD
DFt+IXy3Gz81H2I00QX0IccxGhUcHx+xKZap7Ab3nfQWGZXXi2/5Tj/Un1MKoW+/
rFOIF/htzBL1o1CMnglRwdBmKOwiSHPoNagMMyT4hJHtqJWRtMBk+nFF452nFvyZ
PGKGFuPZZHKkuUEJ7Zn6uQOGmVrED/bxVacqSGSf2CSJClZqEko7l8BH1tYS/bsP
OVpr2q80KME5xWFOBjEw/x0pUPPtaiLbV3ULZQlzqIPRkLYkoy/eTeZudeeY5P35
Fe2G5oEwPP7pBuWlG6QYf6OLlP7IxrluwptRdl/j4oYO+BLngujKXbZwAyfutGZA
F1dB8boXobOvyEaY190e/BZQEnDMIpWEuRfs5pnSkRo16do2YQBK+JB3nxF2Orq+
Y2QBMsDL5mxo4NIaQcVqbypsGKVqXLPcM/dZrhmMIfADtebe0dAfemS05P0LnE/Q
yKfz/kYzwAdEai31D4pYwZ9Mq8ubD5N7fS6vlqUqa5yAYk9X2Hz1VJnon4GOCMDB
s354nwGHC4aBpJd2j1rYnk4an7uVrEFwq3TPNxk0HWWmRyPMurmSElOti9d88TFf
dKrR+3kJsZM0V4lOpaUKXCOapxDUsiUQ5e5e2Bjj859Zwuw/t7B4VoRBR8wcooCc
6Y0kYh4Y3lbqHWsuJ9qOXDhNzqEAFEk46fZooPn2jalkg+EPFA6wV+nVGUA2NiTG
gB9XaD+yi0AtiHxNTuWv6lamAhOqad8ED/O4BABhVxFN6nb0asdP5CPtoQMlS/+Y
sViY/lfvaHovYA/rquZXDWRWH6htPRYpC3HA5PqPXQChN2JcchOZcLfmEQvaa43h
FNd00IWyOugv/TS+nlcVSwsKdG7Jco12tet/O//eYXQhkE3iW1NwiyMX1aldprux
G7g2qcsTOxZLuxaGpDk9JiCNYsb+gjodpaCYe9K6d1vIPqGvu9+yrRyUeksYFP/M
RDDB6f2Tq52cjcRgizJh7+76Hg+qafG89AvDkB8cJyo+izjxUnrsT6OCmajFnx7Q
csC8/MyKFNE/7bY3Ym0um5yc4J9nebEZ/Ju1wlZ673gMZrrvHHy5UCkENHoipydM
A39oQ4IlyYgFsdyEFmnfvMb5n5ZqQy8f0lSyY7b8YT9SwIqu6g/8+FE38XNbaJ3d
Jwm4h/qjZwdEB7NlGPXCyW616Jw6G5Ubtjl9ud7HUuoLK8+lEGsLfu6+idi1yv93
q6/xBwXsgjboDplOCJI1/rfHoe2aJJxS/hdlXf2jD5rxYVs0XF5AV2u8D62YJiJV
WIzF7+iAXGfAxXBBajPxCNrt51XkCB2caGOZ9VqMsCEE6ii2J3XsfUsMbwhlfJyq
nTKUW2UUD3hHXv9C+D+VwrYKp0G1qmkZ4+6XpD2bJ/DTLEsO2MJ58G7SKF5SCWFt
WXZ++oAchDoFCb8au0PAy464fKnvocI3+V6d4w/otHcEqWIN7qJXkA63jNKmP9SE
uvMVrJcYWEYknLiQeJ4+aMmEmisa5hT1za4Goitw1+ufkmZP7TAvqHKwHyoClxcf
Jfcxknj2eY058LKILBdNdRH0P14kOIDRjHfY/x+/Hc0+eU1WjwEAIzcldhzQtmlP
U+Qwjv9rERAvbY3kckQO3PBOm/shjr1FQCrxWtCuriM2x2SjL6HXhPKjwB3DQaXL
MXZnLJZ6AyPSDn1gIUIgPASu5VYPM52hx/EDURf024Ne+Pcm2qThab+1v9cGgKu4
TvmxqslfZ0Mm512AhKe+9x3gN6+jFPj5EX0Xj8CMP03MdU/YkDDyZYk+5xSHaC5p
L8PCDBPHRn5swP0baFBbzBd8yNqSuuYb6OKHDUsDy2FmgVSiu2cugPQQUMyH0GCs
hI8hErF7EtKi7EXKNhRHAw6lHILD7XXSDkqDtoDDsx3L9IVLYIDPohtZK8xk/7xL
bg66o07qvR8GJ0cnC1eV0LjE0zAfOt2hQhP6bZL57/SH3pn40GG68oaXOMphyO4E
5OTWSAK6QUEG5o4zkQXlvOkkC27hZxYYtiSVNEhdP/PSXdOEq0JACNYU4jPMpFMP
3hUFeXnB8SfBbiEKyA0gyZxe6JBQOKzJMcSNkOH7GzI0CNmWQXJejbSYlRFFjP3m
vGik3emGVCikLYptYhag1BhxSN+Es5k2q3l98K5OEUQgk26/QDk767drFMUjXIO7
5WVe9FrMalUJa0GtF71zlasuadRZbkSNNYPkokdoDL0LghsdNYinA0bgulR5nK89
fYp2nflIIHuPib+g/Trn5UlOveYSgU0WwNwxLlXBWBQGGDY5nxkJRSDlG018dBhn
B2cyi8TUN2S2alvUohmasW+V3z+IoTA+CwqKUXddu/M4Yv1YNpzqW438A966aJhN
HQ9ouXnSnvgc8rqC/fufgEGyjxDyzofyKJDMuRh0FYMD8r0CcUtv0w/W6XYJABOv
YS3lOQYO/P1Yv0N3mL1umQyr9gTcX2onJXT+VkxXQBZMTYWfNgRa32wDHpO8yhyL
k10k4LzQs+dPTEV4fiJjgTFKk/ihuCDW6iN3HtNtBwrOBUFq0EWvUS3MsjSunaCj
QnxwgLDbFDJQOPVyGvSnmJW331Mqi8O4NZ0Kf175LwxYafcQY8fn03VON6OnskiR
+hIR92KMuABZKYxrUPOzmo71OpGmUkgLLftRacl9XlvZmSdThPK3pGCYEM6Yvc8s
JPLsB8lmi3dizgRQCWrq56eYr2k9vE2gUSL9+7ZctGyg26zNWPNRvLMSaehl1DNH
SoNEhpxrJVttqjg1G/xAKBu1VZc+92sk7jxoBGAS8EHJ/dtvY4cff+3VZWTzgXz3
qun01HuojjlREhLWGSoaD0YecWx6vm2AYm++v+XU6DHVa9b01riBQqXFRsbMqwyN
v4ZLC+rtq/vbU1LDSIrSLkLG6GxmC+h1s4uvg24h3LSD7B5If3rWgicq+jD6snK7
5AEl59PpPEsnF0l8erLelhzd9K2cmtgd5Q0RLkgwajNzMeChApxgVY8skralUc3a
C4SEW2me21NlVK3jm1J3mhX1KOlK/vHbYFlzBrGApnqcpMuLo5x4NErInjPb5+dy
PXDKohHsNHELIAu/QFTr8uT0TGmTMyqjXYbf+AI6ONeXPAmZXVD/XXc8LbkSvH5z
+9KPgo/UzebHkUC93t4tfMIQqz+cGMEbQRFkYTMcjkOa20INAsOnxN/yL0haOLp9
U5oHoXeXZ8gWe8W+ALA69imtUDdOON9HSYlQWk8Xdil2B/FAn53KKUepxUn/Bzrb
J+/i1jFyrTX4FJCB1TGIvCoPKzjuMLQ4ubd8tZ4sOmG0tn842IvVewz+cxWWJhcj
PTvMBGeNVOxQZt31xMi/7YZIgsOgScnpj9E8hqAhfwlgXPyjEXjKPgRiwfEL8/li
5KbnSWRHAEawLHXlEAWgk74NEXNFU4Y07kyIP6gw9g0/wJm6VJue0ZDEdVNU4ry8
7y0oyqN6OcnQPbJYjHw9TrCW1hdI8pJBj2nm1WIxyrKAT8YmXSsqJvmwfql1j1oG
G7HFtVQKrWtts2ZNpZsMRnZ4EwHXBnkM7FlqUBaBaRBuKxGKyiOmjIE17BNjsunn
4pLhGhl+Yy480He4zrC0gi8+tzmHEL+wbbNBfBH70IsUyFGLyxygD3O89rOtx5Gv
zoZiI9vLlahAV9ORmxwky8D0PG42vTMeyuib2gqbgz9bLq0rTQutJvOpD8SQofhf
7YW+Crm1Rwqd5IAPJG2huOitBsHOdwk0/ymGtTU29w9rQP0oGNBOCtWZqtww+M1W
jfzWymBaZKb7DZOp0J+Ebrr7Od4mJwbuZbXnDhulVpNpAEpl3f/h0AQyW2w8NDnW
XartHNJ6nlk8+QIeeNFLpvE9Xhz2xbsM6hzADLVZZoYLlNo9pttljm+JcBmLlYSF
prudbrAPCYNeMEjEq1C5fUArT+yEaDEVr2RUXpSt0RMHcSdAVJQFLXZdYV3xm8Yc
cwP24BCB+X2i8cDeynKspcdrXowJRt6rH9WaLWusACJPmRAKKLTPYN3XlkuC/M3V
HqTOGYi4cRHTrs1rb5rk7bkgwdUbmovoJTO2W+9untT5Kg+eYoAD3jz/NgSGb8zb
IvTNTXJQLllvBGrOB4T8vmmyF3nOD1c2wvEDv0z/AxwXSGCGYeLU1IfgEXXFefp+
1H/LHHdMvAGXwZUThk96CEe4hKqOVNC2sOe0bmIrrk1/2RjLDhpDZjvkdPvlbULm
1uhuhXrLrz2V5oSbei8XMLP+tL5y6G+DaG5fSj4kwdQoLWCW3GzhvFPQtjZ6s+az
WRpSHL3d83xID9kJ87pOdTteQ0Kw29dWVtwC31oWxE94rX/5jakxxj6jnj2mcnBj
8CDf8cWhsbcV8iulncwaBcGPl68OXr+6LW2mSb2DQIgzapQF+2oFVLWcxhGTLEkB
qAOLZ+x43zX1o5S586KJpYOxRPdL7xPcKpvGidD+X8wzzG1gJV15698bgcIQ3aJz
c5/SJKxdLazQzk5iuOFuI7GLKJwWMUl9qROmzsTbtCeZAzVc1lETRpCVcr9hYO6C
I8KNyWzKXSKMHPDD2PnME8jVeSSmL40oiazqS+d7VGEFCGWlaE1TFrDAWzt35L0Z
rDAd6SiS9xZNQZbrS58G4UsULBicQdJlCTpxug5kx1nuFTpS+Bommmzo/HwCfOo0
kYzaG8AykyIYGFeduh77QSTHMBPec+YPsOYi/KpdvIm8Yo7ZS/X5ZAPLqThkENgv
ElUk5lScl/FAjb0jGPfsafJpiozKJgUJ5OO5XCsRPw/h1lYKd+ximesReklo6qCF
vthGx7eI8qe3SScCH2dHD1bHQahpJY+G4hJkLhXaqo/P94GyirsAieauLT4gHdhN
ZnDNYC97EMin1CGzzTHaokbTPk+i/WUeH3AlmHJNnrH8lXbXy3Ea3UGuNJuv8KA1
xmFxoi4uSOS/rY4ZtfWvANtTfueh8/DXTglhJkEpZ+sOLHuZKrDgfDNl87OxtRni
1PDq1AcoKHvOabPu6j5TaCYLHMxoaK8xzH1Jh/aWRABxy6/NMaaAb45smQ7n8fAW
76XYgGoAWKjtEyxC02ToWeJMALhczTIoigRz5QyGvvQO+KgwC41MxzDW3Fx6YNpd
pHj6n8gZXBV/TQ9fwqI774Ups+Hdr2x/uYL6JlwNvao/irzq6LzRHVSTxBubClnP
Daz2QDULv84z6u6xLG+uZs8lYEfrOimI18SR0HTWjVxGR5I+t60FKetlaACcZipl
caJcAEIL1o52WKk/XMNVWAY+qjVr2eB/EF5AOSgFCaeHcARAqdVYmDH70FW72NIm
JWTXp5/CuOy6xiIuyoVdZEa8P9RFmF4MVSeGN5oX2pQ/sZXgk3tx836UP21PBwl4
T96jNQun/fMJHTnsfZP5jiIWEWcf/a5ohY+iMlRQjUrvbXqjagG5JGMfw4BObfI1
mNOJudiwX8/BhPhwHmUY5zGuYNp45pYM4ouMfuxG55xcYxJKJV7RalKXp/hs+I3H
vdPLCIjumFB62L+JnBuU5wsFt1R81QKaMsXerK4AEL6YyJa6AC2/+EVOcMhJwCR4
cZqdkHCcs/bI/D2Pkc1FgPMDLldune7NsXk88FyWd8X2HyhU+6OGuF5T5HPmDie9
f9cSo8nVnEvHuDwimD0Uykk++TFalie85hPkCrZA2tGtBLysXt9r/kscTyuiVA2Q
cJuR20n+GKxuSKF0GfiRqFkJN5QmrLmEVhDnJesggXM+GjC9YAdxbG4Ui+VpL2O1
dg1Nl3cgf4plAV020GrcxbyH9hnmp8G0Hobg/pJQdY1rWVmOBTsyaTaQ/k/G3YJL
zahLDlIrsNWPIBIkSNRsfqdU4KROaMkr05kBxYdBl4W1amquEJEwtdJDobVdbVRB
TX7VbszuOq5w6XfzX/rJfebUQ6Cg1sr0BEs0JOcE6ejP+QSnrfraFC+Fw33KRwQe
exgmOc9pzwELM3fFYG8mPHp7oH0bGeTMtzf3PdZcA2Nkn0HfakMKl4WVvoWtHlGw
qIcuVILQQf0HsXo4OICasp8Hf1xkPstIGa4UxY93L10Ye605QBUGpxJkPaUyNaBD
00Wz3vrKlkJFqE3uGFhkEsTd2VzR0VGXHxcboiP5xjxBtbci/uwnNEGsqDF3DB2C
U1/xaaFFuXW7xKo523f8KGffCiG/SK22aoC9+IuRB4/s4IgtMoh5sN54n2+8SJSb
8vb73CBdWAUzCL7j24jmA2CRqgB34GBGV3l/Q2cm24zeLw3hF53pT3UnRguddJPR
agV+otSYAqxiCOQ+P2RDo8hFJwRsoGJAgDhh/WK+22uHKC6+3riQRlkFKyFypueG
wk/k/Izm797LogiW1LD38skdyS95HTJ4ezw+IeJX3dO5NM5+HKqmuikBBMhwtX1e
ErGlIc1Alm2ADyrfwDVmUziGAu+wVif3ywKrFghGi1BAoEhNURmg/qeXvupgS1Ei
Z5xDgkfLP8RBK0AeoPk+QHlloXKT32pZ04Zg+SnFOFmbZ/fr74CT0NsyEs0nWbK7
9HF91R8J3tyZyPnoVBCZlGTT9CJ0zefm0CrktzXh4r/O7V0vrF9sO5jbxtW168E/
wuLhozdvwjVkl8muPELaNTGYOPEi5tfH/17K3CCKiUjqnDDZA9/vJ/0wBc3MQWOC
z5At+mUmrhXhkwT2Ii5JGj3OLxG9KKaLzbs1FCWIe2nNS1ZqSxrOsv4mPW37PFvK
gfvpmjVP4xl6jjJC9ub6z5O5NmMeqlREPo9vKK7N5Tx8G4wTooQT/nbwF4R5uDqG
WM7Rw5xPyqyUoWmivcAE++zhIumk0EVMDI2nqO0x1JTPr6VtT9s+mlroA8wIq3WV
9C3nuuHUuP9TSEDHIOll6f2JRaiQAu79d+LZFzFlr2EY42lDqtGyXvSRBQPvh2XU
J6GJCF1pvvVX9O5JJloZuGp+Rb3VgKd+IbedsfcqnhusM1Qukmh8lGRJHg9Rhw7z
o6ZWJGnOAT0jbmY1ZxkQJKqDP6x4qV7xTR78TDqdBpG4XF5k2vnC5vIZtl8+CrBg
6wOs35XT3CgeQURKNcjts+nYC4Ejt4VKheUdfivLJrsAX6FaMtC4Pf6+lQAq9+nf
S6ruZKTOQy2ugp8FtL21vJM5JwB5djiAIK7SUEPWqycAFdw7Cmrx7K9OTZprOhNU
eSdzxtmlOWysz/GW/EC5SlNB6r9AoFdnavR8ynppeayL+h/Y7F/9WrhzFGegZU3r
6CV34Wid6E1JZ2Awms5lPGu+cQeiPOL50i+QYEWrMagnPNH6GrcfmXPFvEiDd6vD
tURpNQgQmPEXqGEWwbAtVYPNXmlfenboN23mbytuk+qfW5Fd8V8B1YH3E+lHS0De
UZARBvnvcuB8PyGfCLIeA9xmAnbvPyk/5X6oMCT047JSX0UNszaXpbzIMdJPPeSp
TYfd0ZSlIs6vJMPmjMCVDy57Abw600Fseepi8WLiVKIBrOsFwvmrIvnHyLb0GGEf
zEA4zMwsA3IynOexs9cvNdgYaVSlEWx/cvmQGaITnzxtakZQ9emsCxUXSJzc1o0U
rHCwWo+IbNcysr90heroH2K0eY/oRbuZd3wULpHOQz3wyQF/bLDkhMSm/Yhhwpuy
NGfJSCEQMt7cPLDoXJYzm3Lk6idJrfscrAMev19iFzA41/LSHVVXPft5fLv2Rj4p
nhsFscUOCivYMwD1ugXowDc+jegIUzopfFi7L0EClWd2sI2SqTibdK+eUtpepCMf
/oIMY7U6RBfJsW9W/c/pLArJV6gGUUd1ZufDQ11v8qQEJv+NNF2g2OuhKUwxDrAP
QhZO2ETSl952Y72gF0EiONkoY+juaV0rj7P0u2GYhzdQqMHNZF8vDHB93aNWdwVD
0o7qmxOxl84XMpnROf6XAg7GhdUCHykzdi9C8PMfjmF7rn+Hvnhj/76LKTk/sy42
Crx3QjkRvOD7nyLMCu3Abdj0CMoy76abs5LOcy/5mmw5BfMUesgwUnESkEepFl+Z
GERJEpgnT4RvnuGE8a50LSsY9QbwvmlFN29aFPWnEmbMkqYbIR9+1yUjTUFxLqUc
PHEaxXjE+bvtHW6es2t3F9O+SXk2MQrr2sjPS6E19cfTpqj1B6YCgJVM9QqyQodS
T6fdNPukOC+Ze0cFNsEiIE8W7SUpcat7duSTvoLP1vTTtM7h7q5p1LYzKfWL2bjl
HtJPTuQNX6D4XBZr8oqfyhNYvj9Nlb892LzubT4kuiJLzM5/KnmBWuXltsfBIy1y
Lp3goadfPDEhqwQRwe8j6IKaiZzO9Qi3nG0+I3qKN3LRRiEzTjtVarBbZl1+kF/g
07vsXG3l1L8Yr4YEbOhEVvJ41l1hw+ThWXgon0z0rEa9Gfmq8+On4G5u6u1eKjW/
fr7UtTQQc4dJREuL6F6B6zquSHK4YzKSh9gzguo1KDbTb3Bzohc2aCF3Jry+Aq+g
IOE6ppFVPDYN4f4ZEyN95xnru3A/D72Ko2TjqsUtgXm7BSORNRbh9Oqa2gZKO58Z
rJSCy1cIQvaOEMoUANFZQ8CtBH3yAgdj81G9BlvgEouJGuwtKjSbRFJabVOMM7Us
tvgdTg38vFWFLlMMJFyN6Q5Xn0rd1eqQaUZ5a+Y2qqK3u8FGW0i3t8e8ANj6zNim
9o/KsZCipMvpH/EZ1VscfDKRRd62achr6PVMSPf27WGTvCvvwl12V72yh11ft8kr
i4lTez5JTFYFs5mtkzust5o9SaEjryWtFMhgeLbkfNfrsKNS/7mp7qIeckeg2Wr2
9/6ThTy2bRNCPj3HDmX3Ri1+b4QOQDb2VJFC2GfcXw6oMbCUtCpWSWKUkElFdrMn
kNZtgXG4NQSMGhj/45WBbXklAkaHvipANs4R2iMjslGo11kxmd8Fpcxo0XsCz0/+
Nag6BHBXX1BnPpJCf777NKhzFD/JhOs5+G6mMl1aQN2swGr8QkrIKdk/u7cltugb
YJnZHNnY7CChPSn/JwbUamg09v92uV6fvJ8sUCx1SAWh89RHFo8LVlS6kjUoD+zM
0Xhmw9V/EmnrMF6oyikPcXqx+KKFJ2tMvdTX/PZvZyg49lHby94a4zsObMWtXYcl
DAq5otBdBxU3EJPZDHBQNHrG3gR0dCvGHBwjM1Rm4gnRJGkzhqI/LWkJwZWuWhXe
EYtXowVkmD/4kn+K7x1xSOAnp8KptSthJ0dS4VvJpe+GO+Tcs9mqJBgEU0onB1iZ
dTSr06s7Lonvjt8Vo8bPS8K4nF0CO6tJTE6PPZsatTZ3wllWvm4dmAlif6mW3B9c
8hDlDGPQB5V5tH7Ew95w4jXcyhGIbrKkp6ZDS2+WnHlILsF3wlvFkhjJjAXN2pU7
5GE1x68/RCt3gNhlq4g7ZzN5TXfKWHosTTRrARnV4rpVYY6hRIxYpmskIOW7qB8h
AJnPk+0D2N1ByxfGtesRDOYzhsiN+DBWt24YPrjq1RoL0eikADNs0v3D+3fabTLL
CPp27nKiA5F//K+kmR7gbBa8+A3471c2kz3+DwesHyk39EuG/m9IYn/KgORKX64N
jJyWRsodT+QEEQ9QFcdmGRfDHm1sEnqXQgE6AYOdnQI0QUiZ/7pLzoWImu/ia7De
yswSWAhrIPeY7pNyv253CyP+hJY0z1ZEXWGNFCPaUyAPHpWlJCXKUmsVKrjnWbpJ
aqDmCntdUJnWLwC/590qOpn+ab8DfW/8hGSxg8Gn0fJaczWcGUyhODhWfgtU8B7u
hL8ltfsZ4ZGzTG8Cjz312qZDHk3cX+n5NJ6cbHGKxlJs6V3YXEP4WoQAfHkqjhD+
eMeiRdtKny3oyuznhl7Pu54SQ3kXIekntqFcdyZRI9U/rR1mY3c2zVu1+gRumOMh
Kq/okpMHSVTEynu0ki+Td9fGNRo8Uu54xn4FDbN0m1ALd+EfMm4KAvM2yiHVnH8D
p+AafG8U/sMhrq1chQeye36fBtQQL6+l6j9QCdFeHQooJkirVyju/A+3Hul/EBdr
dVHcXPxjcT3xlRdOQlPugM+UmAfio2L9LKA9A1nkol9+E+JCpGyB0lqKLTAFMU6j
2NTTbQMnh/XQyb+naaHqTZjW7w4Na9dGOjMbDvcBz+mclr8MIgzWPk7OyHOXSqFe
U5A6+PZ9TRyw4k/aXhtu4y3gMyXHo/SniyKcXez7BvPSkikp2eqMD6LNsdlEU0MY
JgRklABlbrbYUc/wovGNymCOFnIZkuI4irqko4W3Q3ZGg8VPcK5hoEc0qhOFhDvq
dU42JqvvoTx46qr4OZ7LXJUKBiO1hVB46FAZog6hPsMZnrUzyIlSK+CAxxaOXAMu
hMUkg65vHDIcC0M1Y17UHYspx9wIswI4a3XkkcF+ku9e+BNc6MbfFRwZivn5BkeV
qEZMpQ1Mc96zw69ZsFuPIY75/v/UnOoANXX0VCaG0g9ZN1bHT+ukpXiVxD4uKPjJ
nrUKK0A7xMwDiFLq0ylItO31Z61o7NE9zdbTokho49TxezzWlww6JNFUSpnifWq+
2iiUqFtCNlYTm7H5mLsWVadTS9ILbfNZXUDAWFeoJ2RFR86CbL3bUU3w/kQ+zgWF
inPCAOmvoA1tShHUy6d3tXY55I6jkzeYYhu7M831YW03Tq6LyN/9xLuGrZit8oCC
NkOFuaPJUdbq10F5F2nmbKWavxxJI2m8c8jEMw10dG9hCnQ2woR7S/ngcEtoiX8R
UdMjZMWBgi5ZIQN6zk86S0rvia2A9CN+oUIfITwjIxzRmfo3f/S5EpdNe2m/7+hc
pM0iMXi0vgHmthT6Jc7d4m9AZ7x5CI5QLfndLBE3MVXkpilpMzpeuaQFZ0DTn98y
QntknRodEPN11lafexyFXNt7+Mg9M7NW00KDS/Y7scqzdZCz5QV10ly8iSYAstVX
H6jYLM+agvxhzHsDU3MR0/lbLrvRkLy5fFeBQqSgE2VArE99FhRQ9hnBQrRXBYSe
Z/vtwJm7KSTqvOzhPTK8UhAXKg0HxwY1k0IVIcBZuV+3xmvhqWuYLPYmvn9BBv5d
JUTFkhNc87Ly9zxeoUzarmZgQrqxLTo8QKjNwcGlDZCHZj3btm5VXBsqLsmTJ3h+
Gj/o3Uz9WGfPFGW67LOdwTiSP1UB/P198sHPvV3lECNdsPQMZWHbUZArNo0HUWGJ
kpYxaoEy9bxDSTMTBD02qhlHRwLp2+rIJEQDrt/oVkG1ugKzSqe583BfQR173Djs
6aGoex03aSJeHUUO2KSuiolmOgpyztbbVjl4adXQStXFp/DvzxuKGry7centp/K/
R7e6TAI2PHVMRrzjKBLd+T23QF5KsPuKjFYIk2SSDY1+lS6DfYbt9ujTKv4Qdr4s
JHKsYaJYQXqzSTSgF2gBfQRrNbId12zV7SlKoNvnVrZewwpdF/nUzs+8OJX8xmoN
aeJTHchgVMpitr7YQ/Sx5GGaJjP36TlP8O5fwgLE1jRVuf0DrVkB78I3iJfEMdJF
MXz9viinZeHtaiKWAG+CEodLWjdAhGKie/13XWiQKQ396yyYxdnPceulzhTDWmuU
JTs0gDQASOgpFCzBIDgiURzwiYsowJX2vUlRvxoQkbDGghe3HqYnpf1TrskTuwFD
KERvqpQix28n8CaAe4zCVT37tM5fg70hr53fIi5MTYQUOA2qNmlEGIHPw88rutXr
8ore63qz6tMCEMGNRCXMNw4L1NxuQje2XIddcLkGtTgxQir3Z7ssYT52oGFIRGgP
Gxt3EMx2RP7ll3I3qZUjJzqoU2y04oP9CXvJ5PMasr2RH/T90Yb03PVxHVU2ch6V
8JTePsY4yAa+dGMcQCdRS/VDnd+ZV41CpSZPF299dXyxH1LSV0ZaKLX+srg116ci
tcVh4+ftov+edy3FxtJzqA2Q3bmPZCOV600UreKvKwoSgCEKpkyvGv9FFJ/g9Ksw
FMmxSjA0gkTSzBs/N4wXThfIoo9QV+iapACpAJhe17MTp73RmgYlVd9j1Ca85V7d
tJ37E0v5Tf+1SwtXY/0rwxxUJFO0tPpyBSi8Bd8GcG3a363AUByeXJZcwt0g7ijR
rIfjHeRYeH0O4rB3tLjba/5fIOo2a31vix5+kOUPp7Fh6quxLI4AYCi8dA6qkhfi
SartaZcLoJFaa6mXnmfZ3J1NuE74DHKSZ8avHquGXV3bMB6BrD2JTyXy3cJ/9wva
Wrbner0SBuozIkDmvyjb2b1Bzy0JVv87US1aqL8gRbCWC6se3fTd+OrNeSofaRdA
alv1C87A4IwOvdUDpD9z5VKuGR6QXjtNVOmHc0a8iTS9ArZ5c2txBAYyzmGUzYV9
sL7ePCWlqNNRTsI68OgxX/MEGM93Fks95dvEnllv4lBVEdE7P6AbVoE/18e1b2Hw
FAX0pAjY5C6cu30NlZnn7jgotlNwRCJC9AeIUalV+PqcSElkwJbQcgsGTzLhdaJ5
bATCIOZknGHJhxtLVKKMvVRShbMO8MFIxiXLUUkwksv2a/0fsO+qPvdVB2aKOeLO
7p/Wk7FoMrRodP8wOIvCgPRyngv1IJArfgfICXGjDN+Nwp3kr27OooLm+M1HxhY0
qnpGfS+I2Ilobu7mKSbVvYzUF3NOBhioPrIYXRLYx9QNPV+CR33OallFtK31Y+TI
NYnyjpEB1toSgwLDl3TuC68lA8iD8zRsDX4zxo7Dtj1NR8pWiRF/q4TXbQif/e6s
2EJQz/eU+3UnqE/Om44xewr4m8rrNbHgyJkK0Key5MccLVn+L9xj2esJoBd1zT6d
mGxuzvf/dK6ttKoU7ELyaaeoWy92qDXFUxSRhgxvsea+eisETnGQZcuiepTIKHB4
VsC+pNSdT3dXB9Q7flGpbMpJVqGQvBflZPCbteLxcIBc++DcE/BYMqb1lP8qCh2v
vlitViwtq7uPxeT9dtAzXsXO1ifMV66eE5aHHf9Dxu8Ht3HsT4p0V24jssGdXbBE
b7Mmo/ICGz6ARf9hFnGH78e4wh0bouzkQTufcQuqyVUvMO1YI2P7dtkk+Y2ofQhe
JdbdVOB8qb+GVCpjkQRkZ5AoSzFZvCcrF1QlPTKwyk0mz+m0skZitsSUt5RaFyVv
rDouPYt8MjIErWe+2io+UJFo4dbSerdRDSCQGmb2CCB5HIdHxZXfwKHPzRG2b4Hz
MtmxCrCpgFceawBeKwZI7UGBr7/rP+z5CtZXXLPHrFXIobMlg1BkSwH5EnoGSijd
iLUyAyZQjxyPY3HPcx6aCtkUx7LaB/u7iAea98cxO2382gu946GAOZoab46PQV5F
Fc2epwgmnxiYMIpME8O8Iom5B58fS48EuYUny4mOOcedQ8PI9uZRmx+Cy3wYWDvH
489RgSfLY5MCKi8brIA9Iy6CNkgKKfZXp6E7tZRwy+c9fnYrzOcny/ulhtJyV4xw
ZjbhS3b3f0vjrHdTVC/uht6YL1gzIVm/uAmtyNpup+g4slmuoGx7WFSJJP7ZcXaM
H/6TjzLO8PEbPuRPiU+t99Wy/d6BUBM1912u+NtA7lFJWtnAp8Bg/7Z+YGDajRLb
Fi1b8Kw2JBZXLIqMGVd1rljerwCwd3HIzLkJbug1pQxuh3Y9E1GWG9f20kTTD0Sy
tsremuDm9jvWxaJztd8YiFgbXrMFjGYAswHXJTg/FcMmYb8gs0x1o6+rEI5slWF3
Nk38dy8b3j3uXIK3eWAce1ihdUURIvbhUof5io7hL5xy8lP8hAZzsWOlRfNl6bMO
weeemrI/htoCxlOpbQE7jwf2ZdZT2fh7RMVI+kQ0ZNQ=
`pragma protect end_protected
