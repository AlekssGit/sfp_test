`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
QiXtQpmaq44kTrHx5nS1lS19Pf/kFBVM1NoEcFagDJtev6wz8gVWPYL3jSfI1Dmb
KW2HGVd1u33Y/tfHV4lnpiYbx4RP9swyH+ljbR4PFYwyuk06hqCkPyaw9lGBQ+2G
fjiSt1uvg2QLvXlS6DZtp1x7jjkduB3pXUXFOlJ/FDI=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10528), data_block
3kz6dhfQtR78VzQDuIAxFXSXgBSOG7ON8LCcb4ZIDlbt7IWcOKVNnEDdHV4dz8r+
Lnkshj4/4PDJBSORZDs3uU6sVVvIsMZEvnbz4/35qvkU623iUSAfBd+UoIysBDj9
uJdNoLIMQDr5Z+A9oBN3o5JwQzrkQHAafH0TJfSwpPhCVWuKhBsMmzSHzpxsj4kl
Nrl5uN0WXSFc9bf0CY5UZssDb+UUYQ+x5npC3MvXur0hkWR5WIqRI/G+vA3bU5mC
LzyFViLYZfyRo+LF3IEr8U58LUXqqRqMvyPiuZR6AKBMCwRMhwQmDA45I9PUZ2pD
Sjl5ucHR7xe46MzPklM3Gx+7T6jr20gSA6anFyXewbyykd4Y1MPXbwcEsmL+kzMT
tmXObaQlu/N6m0KJHHcE/c4FYey2ahieDLePpnkJi889HkeryJgwdn7dN7Ppoq64
66CLGqKNsJidDjRUkio+5VGX8a5t4/a+PRMGFeI1/LOUrV5n5vI6fx3L5JmOnKAl
IbKhq/3mi7K51/0IVE+8haljH+42RJTu7rQylCKxY7IiPJNsEButkpeBLIKdYvE7
A8CA759+qfwOA1/rSwrauo7tyQFBdDPlJgejRBBJI59CSJgzExfYoKe0OV1QumpX
q/o6YviBL47M4B2FlKMPwulup5pLmL7aSHfaIdfVaG7e1HPLBZcszowhexNlHXiZ
hn0ZEwmXJpBIo1Z5jKbSrQlBa6i3Ulo+2ZOmgnbiSvZHMHOlryA3Y02NaXxELCJE
+yT0Nc4FqauVtPoFaUnxeeDL0wdZI8N4Xbs1ly2dtSE+raBDCL7taO6YbH6N0yPS
bgAvJWN0YwnIuPKAB/ltvmoJECMqkzLjRl7Cc1U+LAQeBZuh6yosdrpf0wMbTXkx
9PxAZvcUtPxc4WBlq+kPvTn0hiB8RF1azfS3WIsjEPe8iJuKxl0JLB/AwpPapqg5
WIWD0f2IkbK08On8S/j2hNmnSpMWkpfnnx5vx/Fpa6/NacGFCocMgWU2221ql2Bi
Ex6jgz+AnO+A11SuvMxers9f5RWAxPWtXLm82Do3z5W3aIdlQJ3EHL2AeDpZ6Xl/
d0rkCdNuoF0z1Iuu/D3vG2o/viz37lXF8U/JnpXuCcnX8l55OfXqOxHfL5UdWusU
ACloYqfEkJ1TaVh0x8XqxJWgPLRxnleK08D0cONwoAlf76rEpllTlj+DJ8zQ4Yrg
9ndPWkqM6voXdvd2k9yW1S3My2mIEe0eWmsuRp7k93bJaFsmbHolx5t8o3U1q9AF
f71nWxWDEJaFbcxYmwtIrYABNb9mSE8RZBw2wOfW1ogT8t9Gs3ntJbG9PtdgivfD
6fG5BHKwzZzG3j80PD4KHzlCOZM7hnsKzaZONR2pwaUDTzx5bsKbcnX+36whUABT
/0SQAlzX6E903vQOMKehXnWt6wNXYsOLaENBJwGz2N1VI/CcrJu1F88YKiW4Rlct
M0d7IjIAkODb4EAuAu9nM0qqWtpcn1yq4JbPtsUrEhIxT5LKYCdf/h8FBXk7kgJO
FxyO22SSlinI5RvZGRfK6MLKzyOQSgTds9WzIAQ+jQgc1Q3VAU56V/15oPLPQ+mo
vdCrPzqxSMBGvbOBGhHeK8NBBdawmgLBaD2nK8uv3SyX2lcomCJ/KVGXxphv1H+E
a+NKq0fPYxuMGex8w5YQcQQkJjf4YVvLS/SGc/nXBeWHecEjkkLcXxNGPAT3Ez1d
jizWIphVClnqR+Wk5/Rk4MTgVcsPAUrKZ9OFTSCMgaq9dNxLdaYiRSF2eG1MwmAv
cv8H8062MuVZO327FvwdRfgCD7HCDGXHroNorxXM0vwfNcq3jGF8twpR9Bpenhei
nJ7Dv8LFEEbt+P2P6GT7WpxPtmcdKXbGz/g/fxvdSWCxJTv1yDwBKbcyxYJLzO30
JczurLg+3E5jkqz+rcf64A7rH161LCyidh2Ufxo/TrSZ70SoRWZfmY/CR4Ky6RzS
Dasn+wyqvuupw4/srUrH98uvOMBbL37EyPHqk0Z/GcajOliEjbQb8lo7kKbRsYTq
5s+6+uolL/EiTxApyVxaAuAI1luxYcLJ3IeUpKnA32QSa9+23ediU7BLfjlEO3CE
XgDfyWw9cyxBF1P6Vnzu9gKsTVhY9aLqiY0ilTuNxaJADZ909bGAEedLMoysErKO
gmIaaa+8hB1AAOeXFjfEqDM/hmw3Hvo9wxAaY3pJI+90aB+lCsDHFthPgaIOfVVh
sInFOab5u6Sny6jMnsItGsz+KJGVDqxhojjJqNuzyVyLN3lSn0nobosS5OwYp15J
pFhRyvyWKSLy8DuB9/+J8oEUUs7md5NrGj4Y2mkB+GUV2jdoGRuhmVF0hwqdMQtH
URUZj6qsK9Fi4H2FDFQA7Q/Hu7mAVkMcXyxnDHt2yIGEEwpoaND4lI+E+oUkutZR
Ky2mmcJz66lLMCAGHTN5PaIv0MryGmpnlqvA13Rrs/QcO5StFWZUmUXkFAFpKjv7
yU1ACPKNqxsAsxUUi6OK5EC+d1ozOUPaKFUIpL0bb2kwCNJvyBgAolWmeQXsYZHm
hcQ0kfdl73c/GqJxVn6Ma3cEglSMz4eBK0qUvBeucQkxH4a808T/7gQ1REQmEqRv
I5+SSXUbQEf4wcQuVtXTxvO751tKAXbvlzgDiOGpMUou3RSujXYyRb1PRyGpEXRP
SjNyk+wnOH5wK8DExIB7SaE+vCOjphwpwuj3F48bVU3AqXniDWBjBi2OHOAh0+3f
aw15w9Imxy8s2iKKnmWP3cXqRq7zUFLuZQ6htBJGso+z2MHt3w6M31LOSaH2noEG
qak/n74J2h8FBa8Zj8IoTAIYChqGhVjsVc0U8qAcBxZ/ymwF5G3G0W+g/Gu07aPJ
MjUrtCqTGpZb3mi+ffPHWFUTgUESPmdsfIUWrb24qMFZMAOobAdOrgK7yiJa1AnD
qXc2h+CGCsl6g/8dpODLbKL1KAg1bvvec8Y1ydPvbI4Uwax8eLzypHf8NvUpukuD
JOqSNWf8e1WG1C28YaLmv2wv36IuBHzxyAN/C1G3qwBZLDXKf52+15ZJiknVe4r/
j0RCegDioziQDtsUow+yzuPbFQssH0tJZZzznXLOiM/VO16O+0hzPCnpg9PawLHE
VyQIBDuCUYi6mOqojmll4K+D9+573iOgFMl3dlDcfRLzHrHFdufNITIgahY4cVL0
VAE/8hur57wtbgkQexZkeQ6cH8j6Q0eIXHyZ80E0G1J0A70YKQwiQcScQflEXKQZ
uR1AXYC3FMEql2MWu1XJD3vgZwVzK0cr9mSr0lnVdrw3uBVfsLgcPyg0d/bRpXTo
ZjVvteevH20PkUzALRzeLhOA89+j7z++mZbbYPXnZhzPp7s8uW+5SZckWWRM5ROb
RVwmBHg2RtHS1hImzpob+mMdVkMrsLpMirav+YpXLVMU1pKgZjldigWeEj+esNAd
bseVQMkYnCoJ/8Q8Dnx2upIYuPuy7rmi6hfqkpMXMp1J+7mIYaCJvF6gUoKXMyiE
gnr88v21aVX3V/Na11TeQjJu3x5cTgoqmcT5q6qwaOXcwUGeKjALO61lCLNqngAd
/fRYkEQMG93FG4uBgzBW8LdsNAbxdV3Qi+yDtzJ/MAo2Jy8h0vNpIX/oGM4dQmId
KO49HDZDKAAK4xSc1iqkZikYcVdc88GpiqXIjQ9Q5UFNe3lU6p4opTdDkcOCHZpX
CX3EagIw9G/V6UPSXTvHE1HFvJC5LCZH+9Qg/XDlna4BJvMrgQu9MZkhEOv3S1Dy
KGH/DuWAXS4mgVBvx0yNOLnVZ8E9+p6Od7BhZqx7z9GN/rPGVq5ODLyGr+e2GLZe
OFT3s1xp6sXDOFp1LMwak+YM3nXGMzhC2yIlvuRUxVsBoElbWNUn6SCwQLMGJHTc
iUdefs9zQzGssux0WnKyGBVv6DhlBKBvaioSCWLX/pSs2eh4whmge+gdiK9/bLMW
fvGHB5iZ4Q5u8Tef1rX2gOsd6TzwU3Q9966TltYpI+6Exj2Qz++jY3pnEI4rcRjy
15hn5TJCihRx8YeteeDeUoSnzRv5lLZ/QrcGU9ifnAXEsVpe/4rhovMszJOkO7QQ
a9WaKoKPy0qIOtqI6YerfXB0abT+fPYBOxNY8PbhA8Hi5xO0S3iHfGnd3oINFj++
/xi1iqwxfAtruE/XpXdtptxZtlAfyCbriR+9F7pSgA+7j8rnJ87GdXsSQRPMB+xx
SembZw7sMUjTSjcK1PGc3tAbTjefSU514At7azUMuqlwrfnaOCn3KCfW41Rwj1Vl
g/s8cIp94gLVOsIDcgU0mkB19i1Ognbs28nBgPs1Wno05zNJOhO5u86sm1670lsd
zAQdGxNzG4CBkEXKG0yVgr4FE3J3PG6i0OSa+fvaiNZSoDQNAQBYdSrNS9riF5mR
LI2ZG56NPMrh5Xdn7dGgP6+qPgEU3UsZFEA82+OENGMbxN7ZZfg0+3rD/N/We9m4
iaL7qJSH2Jk7mkwyITC7js59kFsJsIVPZ3IsV66ByRLKLQrPQJzj6lS3vUk58obW
WaZL3bzKYqvokVG+ziy4VEGTkdLhFXoIvIjx6eab5L/kzqxHejW1D8aVpXlITXNU
JYI1IDemx5FwbK0V+z8NpTRlYDfC3eZK5LChkvoxHj2oRO+cjiDGohfAxj38EBEn
n8VMQRV2CrdVzj6Z84vCVOrviIoYl/WUlS7E+dPN74CuWoI6DOgMCwXGuRLGDE1A
SqdgDXbVUsnLZLYzdgGuFvUf2NXf9v+jdfny7csW5JcKhOZFGHi6a7O6nEyP55YO
9ydbdsuTneL49Hsw30VzqavME97/avPorsLdqz1/8Pq1mbS04ce14SsEsJp/EhAF
PewqDepm+N5I/8A7DNWw3UKwpzCiDjNn7+oGNbzk+gHUkSurpwoRYb0cTfHpALyf
kMMLnpI7gvpylB+wVGJrhc5Wy9idaBgG+c6Y5NJ7sdIPOhqC/dzDBCOznJ6NBdta
QDPe6YvCfb/PadyTTd5tJsjuYqQu6rZifOP1YCruR1NP917jKiOZJjNT9PSfYw4J
NOBx5ZU4GwpKOY7y1GgA/ZNjuKlKAEAZz37i6aCc5vE0tAY7J1hRdb8tqRR1cKuG
NEHxgB1V1kAbqr2aHADRmLsUiGNpHR7UTlMbLY2TPKn4xenI1YNs2KqDCYmW9/eo
rtfvKbDu63hX1fBDD9CkUjMCVwQkaf+xGBkURBh8w6ZhAv+Q4f21lOFkNYofGkBz
VVBLX3j++NNmwpKHpFwUm0UOYDAKIAjTEiudxjZ6GAU7ED7CjLdmNr0XOOQO2mom
5egrYjo2JycPTa5buWx3tARZZEIe7VW47BCZ4ftMCryyji9+JCoELqdFfJJN00SR
kpT0q36cozyeXyGzRVECJvL6z/55SozI5D9SbsxULg2DPCe6MGgDtfM5UtgoU1N9
22qjuVAoOhWN5Iany8r/lX6i38rKu20eOiHBcvTfcmIff9um4jyZtArw71qMKV2L
5OpLO/fTzYq6pR0WB48VKwsKcVP/sjBkU+Iyi39VhhUZjuWb7x71n5eZKCamZuyD
e0QecEnNqKvYsEAe6DqpanfnVT63yrytIN9zGzflRiYFqpzx32tvABHJkvy5I9wG
5fDOiElzHC7oWW35M9gSy7JjZgU6jq/ORBu4hmbTXio8KFFVa7pvkagGS2otkZ7e
G0CEiHTLIKHY5pzsoy8RXjBce+bU6SbFWDCv2yfXc40j4OQvSUTjxXE03AvO7fsF
JL8oYYBtPeUq4mQNwEk7BsWGLlz6HXoQxY7pKG2Vd/SeFEAWYrnkPPMSIbFTsD8/
yBGw35lYar9WTP58dXK2mM21MRwcJgQp7JJaRo8kRgl6JjjRLuEjmwMlICpWzphD
cwKcCY0H7wtA4+miBELG8kzXsXSyObeBwJHYcYMU7fEzysXkE8w6z6TL8HEMPrER
OS9vVvjuEmnivjmWnnWYNbdx5jT5ZOLXr8oFZsV+YTj93WSyDi8elPO8ExhIsHEG
m1Q6ZroOvO1UzCyqPblk+70EX1ASQf6CH3ZXwZbPJZSBCcq6cBYIw6XbmW2An3Qw
Sdh94vHFQtoLAG4njUsw828GtmZcCQGDb7TUnwPJJT67ZTmPknQkBvwGEVIXhRSa
YwC0e9R9l9M+GKfmarSOoKijZkbhoSXazoGhuiDBDKnMphZHDJlB4jHxb9JYb2Og
t0ozQyWIYM0cRvvc36CdAGrA59MjPQiy7yZ4y3aN7DLxlM0okXhaytzIi0hoe/Ap
NVKfmwwOmtk5syTjzlDIkzCcbeAygoJOwFV0O0N3Y3Yl5UT4l2IkBx5LMOKc/KoU
mBhtPkxidYntVtm0oy0uTnP0qUwbh8O3dBCojLO3YpakN2jhfCXyjP5oQ1shK8vV
oEpR319jtJEHYDI4FWFWEdcWTnsYzu+Dyz32X3IbrGgoPDvW06o2MeW51YsYix0w
zNnv7MzmlQriIGnIrRLyNHf3xvGYcSUQRHsJ30VxfX2EKRs9phsd1p8wqxTA0WYL
wusfBD5KsZQiTIu/ZfzVRMZKgKrsdlPmz2oWUet0UTTD8I2hiKNCT5i80jwuKDK5
UlFyHwP7TA7O/2vdvTozzMTosfCrxZ/uQWc5VUwPsiqQ7EKONYxDp7YsT3qojnJa
q+ZmpJF5N7sdlu0XQ2z1+1WwsKmftpDhRLJrSWwTavtK6yksfn3y/zAPVsrLj3G1
cK5fjFMGO/oMMM7mw33KcGSeBY/g392JcYkCHx2Wo8CJCgpygJeLm83Oy2TN5Etq
pRAa3ZFqCiyaSXrKtzYqx/td745jTJbjtNtfDnxhC1omIx8SHpb44zj1VDiKWxnH
5r5+LDF+ZCF/02UnON+Anpk449Zs5DWJipY8Ij9KSwioqRFC4ms+gakGYBxKUA1n
t0NqzvNm61uhW8hRAut6qsmrCRFA1V4iRywxDvgQggMzoT3pleUzV5SKBxLdxKyK
WxmfRXR8ygK9TnN8iZOmPQRxJgwiViw3/0q+lW78vYlmfdw10zJbY98eN17wT26I
b/BorWrALjUSSThdqQmHlLo8qBrrbk+enatFHE16tTQ52LpFAuseWfb2neMxCWfK
op62RtNQNw5cHGmGyS23C6CpAmMGHZX0/uGMEHqfgiLIrR9YTEn+MPGTbx6Ef+Qk
+hnddXs137/LFFZ4sW3G9Vkj2B4pIs0hiiHPw+UBSdTqKwMhYdDPvs/tJlxuxoxf
FGp+VzdwpPFE6zYTneiqidP7tYEpf3xTOtjMirz2XZ+7QEC9tajV+UA3xmAMia6i
/g9sV5i4yv9rxx2Zvs2XEa3FvuYkjkaL0inCTOx9dvWFc8RbOJu93Lco9IRXQNTI
66VNQ7EQATZf7bbJcZRSk3KsvN9VZprVbVDOOteoySI8V774AvY6R3Ub8HICe6AC
oaUXelfp1LMq6QrK98vnPOo/tSzBnEvD9HDXF+jykh0S1Rk057bXcLauE58Yoj/z
yPRsLYEmxpsO6g5hFe7wOFYQ82lPiyjyYXJnDVyL6C2DtpQM/ymMlnDR4VTTS6aI
BubieZ+tCIwC7xslieRAi36j3kyCoJdbNaAm/7ktpoWgIDHCi33/DDjMPe04xfNx
4PYl/LjOpstStcHgJlzJxURY/G9ADwAD6uFLimlEiPjE6w8yk2o+QskiA8ExS2CT
On8Xt0ee70Qg58oKhaNpWJ9y5XD9Wv0VM4BhcigzqXpb+CCmWruWUpGN2BG8zYK6
xHXW4DLA0ZGaA1ZP1k0lC00JGhA7WnfaH0SaQ6c9XA1RjXDjwht4fYR7N2rJfQeE
iDpHUETNr4SGI6qiT83CokjMbtTKdvgBpp14ImDgc9thfMScJFe7v9HcSYsbnfPh
flqtK3ZSzjSfBpqcbuL1mNBFwDmWJ/l+zfFQ6vfogyB6vqH7UHxtw2rOxVGnKfMn
fxHQR/XcRjY6Gy+yZIARoZRuc4KCYs2dVgebNRuaBWKKjW0pzPU42V0QuEuq7ifJ
vtx6s/+KphYfJG544Vf0TFtWxT2DOpDAfvA+J1a4LZ+9z8K35o1IyeJ5hXzJgkGq
co0/8JVTW9MCigDV6mJM7LEy88EIXn70FiOAn/U47BAD2TkBRrCSZWzJfsphx9Tv
+mfn4m4P9ZlTR5NYAk+UrVX61/HLQVZDNZmgeVVuKNyTZg/aA/yTcmOTw4dPJUFJ
da2xg59vPpehfkCnT+LBskFA/1KSPr+HBMhrWYVZAJCFFuRJe6YIuM+vMrA1S9tm
mRDhAfN3LLjLMp6fuTFk9KxrxRMnccf6W01hePQX08otYOuWCwgozDHLh4RaTsTS
NfEVmwadATrDP4pGomtIpQmA0R3cwCzV5XF8ASY/u0CxcjCPsTNuF94bMC8Pa2sq
w3mdYH+SN4wI4BD/FQSAAUaIB6RxJ2r2F6JeL8UN0VX/MTnSL8VDKJoJTf9adjdW
VXI97wf3ztVXg3LDVukGBLoIgcSP+SiAiXHw+KiO7x6O1PJlhMM5SC8r3G1bpIhS
E0ST64nusqg2EJ1Q2QwFQIDSyC5J0WS19aTPf+zNZ5J0LAs0Ee9oUFDJC6Z82ZUG
RfoigWJf+Z3Y7AJsXuoZn1aStM3kCOmzL64ewR7OBiBa6cBaqfuNgAuIOueem0u2
4vWyOsA+aEDoG3Bp/H8NGJW5UTFkJhhYmKsCsYGBFcy5gUqQ3aeAeLuMr/agUjg4
pQfoEiWIqTD9Cx76mCBilQrFPaCAO7ZyCd5hNBj1FqLdN4GK/wF2DRI7V2abiKU1
k9lpqeZCMEIwOtUxEg1wJv6tgRTjj8HumXJnZfBZlVpVlIuScMnELq8w0/jKJ15s
6kfYsdzIhmlosWZfhZCr9PTJ2GpEVBY2XoKpZXw9cn9nJesEgQGcap0hRjl7Pwzo
24vjZUStYWrDJMvXdb3XeBjaGgTEompWOPNbTlBt7tYL/W+QpPXINW/oKcvFzPJU
C3iohGjv+ndH3An5Y0t8OA2FWZe32p+5MzZ2uoroF9Sb9OGo38RI+ElF7npYct9D
MA//9apvhalGAfzGU/JyEVIuvt8mPtDpbeg8LXHR4A9/BqKTFF0BqBtrgsbN0vPw
PThDEAcmrLbtRT1oh6Mb6KZldOwTK07PfnGOqnPXHHXF3PQ254gPyDE/5OUSqGbY
ApZFvxb2N5Cae9kNrucCBdi817Q0Vtqda8Pvx/fHAZ0+6e9sizWoZZ/Ge2gLpJqN
sodGDTxFDr2BIkZvdMExFdjx/QlyamRidskNydv5bW7aAikPcihun6Fs1GK/TR1U
aNjgyTFZp+4sxvtmq3d0dMaPeNIvjcD8kPD8x2RWazu7dm14ETRG3ruRkxQQbm8w
6xnGLLOJJDYMUBDKP55AlRvfJC6Vl4yYTpdgu4MOfrWAyac3RwYIoCTtXOVxlFJV
6HBVn/dWAY+nRhrsNITX4KeD6r/CJA16gESMuNRxgw6FSBFQcQE4YNcSU9BMScaX
kxPgKarHYErNwEORjg5+OEXjUaao1v/ZChUGGK9e1rwPcEGKziD+hZJPwTvpzZlp
xxBmeRhCLg7mM+5TLw0NpPaoTUt8UV1WDOHKLQQZoPqJ4x87UFL497IeovTAIyfE
nFjf1MGNV5ayMt8akhWIDLmufqcfzo2+YuG+6MIRQ0LMbXU48NKMcjM0qnz9Unmy
UThEWwJC9y0fLHI/k886G9gZt/m462qTfz5kyelq5y9yG3N3Yp41GIWFhqmTeYhn
9eEojXsdIAXmZSYqRUizk1pDUvUMExG3a/XqHGmotzUC1dHTj6hEiF6lS5WcWK8f
UuVxvGqcHnZocTG8HsT7gtLw8o2FTx0VKXStOxvL7IGWMyEQZ830bGF6b4BBtDJ9
PkQ6nHKttMZl96ez8Z8jOiFtgqa9KXJ90KVjIaWxwX3M4jAYjbgBOYqyWY8IubEs
x76EsdWNLorSrns7BVVyuvnkPpz0QOCGsth/KFOATLKZLmLY4Zyxd6E/cK7l9DiL
BWmxd5GBtanC5UhozNyFLAoS1VX+/XO/7r1o13q2w6oP9DtUYB/f+I5kT6vsARmA
0aSAPlu0PVkBcWDHLuM0isCurGTaZEsQqGkKB96RRNGarmaFMh3ze6P3F1UV3Suq
dds2B7khNG0QNkSauiZI3qeWk/W/717KcFsce04OcZHOemdIFrtzw8VztXcxUmcM
gieWtxFVvTCDeqGm5DDBHNVkgO15xh84FymLIJPHXDg0grM+74QgacAArK6FG73T
ADmyypqL44o04+smkb6CGeLNHSRA18TxQ91tcFWf/nbmTO6liF1rBJiWimMH9Xp7
WQJ36EZmFjqjugp7i/Mh2ZG0QuzofNhDEkpr5iyxOLM1WHXjH9u2dJxMAOSgscUg
LFdoJX4c/uhdE73IkC2uKYqMm1RAE+9tCHk0XWLsMQ5pxXxGOiiS1JCiWKKhvmA/
+haaSTh7eb4D7HJDHDfUNBOAiPmNDoddKO+5ill5wkaj8kpMKz0m6cq/6PfauDTt
Co9Or59NMbqzBcpgj5QtO2DYPvDWwRLWhrc7IsnUu6HRKoIPXThQUDh5PZSaoSQd
n5sNzhTan3sKkcLSMBLrm0RwTx/pRg36IsqnXfZqFds6zH9/cyTsel4eytjWSp6o
4Lld+ke9JJAf8SHRTFojEyGNsT3PDaQE6bjXnLEiz837PeP27GxuRvJQw88Iiv5x
vH/QQV6gqbvsYGqiC4aS0+fTz3AmC+h20GYeVVnZ8QorOdRAWJyLZP7ZL+8Nsury
VSa7/tUYp9W/4YERxNHALFavJ/0lEFp03BWlBMGzzhtl86vg8hTjKKhli68rpblL
RsiMfeuZMgYHJRcg76NbCfOfksE/YHQn+jp6Wi+GCwxHkNWWlMWr6LgFcRajee2K
VjXEVQWZHniQujfN06QamR61w79/l/yCKU+z1FnFf1sqZUinU6L/Ond2T2NKhy+e
YWgAyEbyjf5Bypys+4jfmOYedOwHrHua/ogGf2PNlwkxLjJJKltVRAMo/djYzHhL
e0LHYcPl/YSg1eveNCcfpkbGiD4DF44pj/71MelZLrjuctrZTkV2+moB1VBhLORT
Cn8TqpWFSqHk11wacgr133ThCFmgE+BjLBxmOFcYyW4KS5UT3bZkjiREgs9rABur
Nc1ll6d/q2S6JVY3PkDdBB/xIJnWPWS7RvdTm/BuRszL9bPZx/Czs7LjKF1FA4bp
/z81bwnh/VAwY9eQuB6xr24nYfdY+3XP4mG5SVrKzuXnIE4KA8Zwxht02jv0Nx8d
C0ljaZEGx/h/g/2D4HuOd1Ad8A0YKneFFrWFUlm4j1EkFeHw8MHLDu6dj3aldhBj
3QGLHdpov+qqtLxsGs4jZLzrehST3+NL49qQEETKr1T3p6Xjkit/g8OCPsvHiKwd
CtI5sJQjG4BrswuR493yZE9SIq+Po0ZMCVe1mE04rDNfXQkud8l1IzAEKNuxpgt/
CJrKM01qrLCrrsoxRQS4AS32r3MN3GyisFU2EmDoH4ZL6g47Vn2hovWZDkZj2LF1
Q2aTK6AbnL7BFeJ4pMfyG+GSp6StS1kiZbf9AlogBL1tJDO8BEIFuGkfbCrcOc9q
cPLi2ThjK6dXr5mTkUBBGsPgRy5DxyDIuniDb7c+urY/dUaD6jwyt0v7SyWIemN/
x7m0krzYNHs3whflJTSDLFcbGMn9M4vHmupo8orJnvBoVoCkcpzceV8LsofBK9fq
g9XFexuMaIki4+Hp0ZKjOJDqYxN2gB+kgf9LYUaZRSSz3hA04aut9qAfH2+gIuW9
2ivnyDnoxEQUQbNNpjYsTZbyUY2g1M4IJumnMEVpgazdi5IigfvYG11MN1O8vptk
tHVm6nrIyg/h6mWrW6kTDHLxZjOgIHZpwxE5VZrbdrCfM5EnEGOpllgupNmda+QI
ATin9g2Qmr3QWYwfa5jfcT6GroGdovZUbP9i3jPx6/Z6WnWPOda/Nw6trmwbwL+a
S6O9LOgSSmJMwKId/LST28LcDRY7MuvP3/9ves8gk3RU3jppWzfo2t42cXJ1mIFV
ovCL5YcN1s40yJcwL/4UZncOzWgQo+D3lKDixmj8tocu4fPCS2cFiJ0zD8LLFhWv
vNJHuWehMaH/cNcKWEVK4ZANH0LjN9/MXvyH/VkOWPYmetC9O9x/SegkEJ1b5ga6
tnnDPuhKCnZg2i+59a0PBakwrx5c0Qp+N1CmXSVSzzbGJI9BOL3WQs1QI9JXPTrI
qGNVLVoN/rPuSShDOXNxSkSMl/dxp+OQ/vTkom+Z5FdhOX7KZ9ymEnoUg5laPElX
DtSs1usRQzdj1J9iPSTjxNZe5qWiO2sDAOGQi7UJbWmfUsHC0WBrVq6XGNqhj73c
ufIGz56mdnlkwadlS+O55l3VgyEjC/EHsj3kPvYVl9WqSXCrf9VZ6h37QMfPhj3X
B8GR0wNSBiImYtSB1gKjgzOSBk852vMI0tm/6HRwVzPhm3hnglIL0UoKNt0I7YyO
YNaPF7De9xNzypJAilE/ZESgS0/+u7Mb2DUCs+Txsld2etcGiRLeGfz/2GPAbNLL
HE+rnnyHCGPIc+K5oDzpc+go+vSGkZVo91r/qKnAgcICo5UvWtJUctv8l3AD9yNk
9TDM6IdxUeDqHJSdLgB5v5MBsFHkIAQDNOAgKkA3HwelcsV4SIOXVfJtglgVExep
koBO+62pD5pN9hAjDemNXLO7gFfN1B89JJ0UNi0Og/B6kUHfGlSgMvqxPfUZUtF5
u4RoRATlwFXpQdbNgPNykQyfvS4N7kiiuAnGxWZlxiRJ/l1gaVqlUwRo3jdkFsmG
aJ95ZT/QOJcjEoIg9UERZcSHHQd9xv7yfDomOoSt8/raJrlfx2JHeQzqpyxxez1y
LYzXQ90YVU0POsjUYpa328aBGjYtKLJNaKUmuYh8u6kRNpHRmy3caMY4zHQbkcHW
t7U9v92N3SwzPwuhtttoA3pDuMk7k7xnvLd1J/xL+cJ784ifgVh5TCFFVa5QP9Ac
+3UiQs4/zSMKU2jixiyhwGIdmcdVjNFGMJEuHktuwEncalD8CQd0/xS2O8cz6pXU
3EVVVXo7Nf3JlMn+QoOHhafP9WJ8HrLjTZVnSqeYgeci1WdT8VvuT78xkFUptu+2
bwv6PSp6Z50WRIqfpK7ux+8PDyak7V7LuPCUeQ6eOxy3bRlmEPfYH4uiz9eL7kzZ
2gQw8HJ0HqDTQHey4P8ZtNfsNGItsLErMBkDt/B+NmPi+HqCA7rQ72AmGwAEHkBE
N9sX1yJGV0IKKhTMvQnJzBAJIGPRqVD0ltSAzsBzfUyUIZWByD15m1kEnjvdMw6g
kiL8E1BBDkfdrK2rptdh4/YAUv26zzYAEQOZEA39R1RkJ+gsoX3QbvJ11Ao8U8XS
y7ZOwiySABvP5F54D8RnkLdSoLbIaM3+/a+Ja1ipwlmN2LEpf0xDsmMxbk8BJOIu
AipLutH7hvwV941PQudMlEjkHl3LWsEE4veynEWZoKzuzgoioTNsu0F/0IrPPdkH
ly2KpTkMiFSNz93WnJ8FhZ1OxTL7LuuJqHU4vUj8Ex0QZPWbDTLcy7LbC3A6d0Sd
moq19NtQT9pZSl/25RUyfWKoc8KbP6mqb5g7a4zxssNJsUcDmirXsyPp8d/wGruz
QCThtstuHOb0vnjjpkygwodRdMjOax1U/zUGfX69Z7VQvIdsZsiDOLIHY+a7hsog
9tXvS4bBaihCqlodqkWMcHLDGPSF8e4w1UUeG7yzMx4F9m/6Ntq99+YfqMI1SxFx
sGr4HCvMUNDMPVy5aDQCFv1ku8gQg+n7OWLH+BgsR6SNuZc+a8zcblkvewvRQNuU
q5JkoD9NMFN45x9E7M+RIIaCuvfHU4t8hEJRK643sgDl2oxQipm4Gx+89tvWeDbM
CikMaatQ5Inbut+55H1Gh9E8BgVKfUCLFGEVGBfFHU/0TB1+UpWn+mw1vcjWAFrQ
P2fSYfIOpYPiITHHjBv/AzhpDNiKAde5qGCpCgqxVoc1ZWu4TC1qahj5V08pq2Zg
arI4/tyxZrl7Iy2vz1tTwg==
`pragma protect end_protected
