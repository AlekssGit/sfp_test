module clock_50_out (
		input  wire  in_clk,  //  in_clk.clk
		output wire  out_clk  // out_clk.clk
	);
endmodule

