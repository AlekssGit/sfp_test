// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
kDj9J57cTILAdlcvAASmEkdYSgY5m5WNwN8naAsg2cjjf1TAoiit/wwvM8Rl5GnhEtDhLKG+4R9u
OO20NPm0yoDXrAraNrnQDVNgoBSUj5nJHTh5O/CipY36K88Nweu5/XxW++rRCg3zswBRQxUJ5fJF
V/Tp8XkK9PzrBbrcvOHbSDXVd+ukSlVthvABVETJLjULP8g4fWCf4wyJo4dx1GeIonE3iECAqrAm
UcuyVAKzP7JI6m7fL2jgbnCqwEQn6Josx0bvHyBQL2Ux87luHuu7WElmf8e4/FaJwn3+c5I/PAgR
2PXLdDqp5m6rTRR9CGCljzz51zuCTh954Cl/0A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9248)
j/ulbnn/R6CRLVkkplktxwDrrUEiY4hQoGXkUoyYvyzOS5lMv8+O/9gKI6V+BqTvJ5hMo3fhzsdZ
Bb4aPF3TuTGHIL66Hcdhv/wx/bDt4fdKzsdnYVkUQLEL5VO8aGfJJtN32nwWT2u2E7b+im7QCG0U
jsvpbfjgl7K5w2yxMqDhLm08Qdn2j+ly9Rucry+A7e2tW96UIbSCcyDQg+b20Osu/4R75XzGlKKZ
afK96KKEZ0TfqMcS3NRjvJoJDW9z45KgsOSFeAj1hL0NrSTJnr49feL3iLua5M9IJUt2m3bBRxt3
Q8e3hd3S1hRWxKQD0Sbz1mAzL1OrjrW6f550VqISmxcEQG5U0ERFo+hUFtaHp0qdSP8YdPQNwPGE
dhDYkmag5wNZ22P3wudOd0xJTRrq6OTmJkdiG6NYSe4ahQfLmMeOsocNq7K6GUh6qB8FWI7SMpSg
uUrreCBWvRW0v8j+EE4bwBQv+ZQjB1qB/J4qdyXHGnus303sc+P/6fNCPKR4fgLhLAsO/jsiftZ+
XP13RhJQGlpErdutpxBURA36uCRw9OlsoMGymJdUK/DvKxW4ASdNannPLCgjtPsnzsD3igUO+TEP
sma3WqEHVp8ECXMUumOEUVTrburxHxGgd2Zq4fkngctjGWQnRy2FCwV95l3qje7y34Kl+2S9ZkdI
WjWXt6s9oOW3PE+WT99obxWRiqtr4byv8W+btIaTQWgfDxsm0li3fyMzTpa7IqgA/CiiPvBhi0c/
fsFTX4xdeQfIK7p+oU0lLoWpTfPP+JBDpR56I+lKFp+8DJU7kt+jUFLSln8yRQhqMIUSINel+yAE
waOPr9ltr23LgIYlDg2mD2ii1GA13hdYrorwXcKn85d77iRoe4H22xyGE9rRvkAM8yufSNaAuGmt
fIizTreKZAVfNWLTFvx46jU3fGV+Oh3M+xEYQ0OvJ8WR3lBuktLPW3cRbZTdvr0sf1QCXPiXxGHI
c8ebbd9cZOmPcMj6lui0xA87pD0amCNG+sJiX745Cg6dRYyVhrm61LNLFHLNJFpUPpFccsFdWDnY
s09vbU3J/yTaunt/n10N8ZgDeU62YMTjJqx9UFXRQhpVLfYZyhANud+XKb8ayv7Vz/VJTmW+Vb+W
4kjv0nLqaw0J4iaq5hWXMSvLLzSb/OkJ7VJDHitAEM7kvx4CwbQNQa97nP5Boko9/Z2LAThpwo8t
jV0+CWEH1yYx6g1YMHIT6/TWVMfXNmgrnRW6XatfHp/qotlmVNoCQrQdlCaZ0LiWq0EUAQSVSW5t
bntKsKQV2AAa9tlRUl3bLR/uq+GjDFYXJpFY1OP9NzIL/6subge3sRIRG5jFFuX5jjx+tJYj/yt+
nD0WVGOi0U7DyTYEkMo20+kwXv2YCGAhyAYmzE6t2pZ9GnJzUbQ/j+8F+vf8canY/+RX6geKKedS
f8SVntyzRSdckA/t4R9N/L0EvcdF2Zt54hQYrs0z+/3vlChWYYp0I2NczgLdYTM6K2qJqaFkqEoE
PTFDCbZW3f9ZxC8Bn022dknMdlILv51t3Au/EcQiQPLZEwd49RG1j/YYcc8pL4aT4Nyvkm7jTJn7
+l+8wSGBg97GEv2QLSWK3SJ9CBKmG6MXutiTvWGIBOkzZJkePvi3sLsERoYSPiLREs5BCqPcl3zm
3EDtUp74Dyxx3qmM7bt+Ii4iPNP2d8vrAYWrndewT4B/Qk0us68Lee0X6fHC7+zDzN2Uoe6ph/Of
pkNwo/j4W/fVIuG/Lm5N76lwhYDvflpMBrymThQc3NDKCQHGKFl1Uox7V4l+hCvLXeB4rpjDmFUq
js6DKbrzR9wTSyv5mKec6n0g2NEO8LzHz5499bAYG3SLeLTTvdb2pfPe0LRmmNVzdCYN2SVVpEkq
ouGq7RJCHsmpQBr1WxWUJyAnBNTvmdiPXNVzBNqakTUUz/+SsQqsyxrbFZ7Tv3+dLYoItulqf9z0
HsFBSA8mY2XkfPXouUuvRwY2SGoHlHVW40AbhEaYNGkHBCQ4XTGF5B/SD7HAaL96idvZDFG4JVxu
des0Z9cHLzO5x9ov+KKMdZPElkUBL3pGohs+UhQqbZ1j+N8z3fC6T+/wwMFJdMHiIQbvtICs1IYn
TSg93Gh2thW5KFqlLh3cDMAJJUB0JwKIw00OssAkoSAsBDM3MhlMDTs8u9xb3UfAgh4MmcMunQA+
UrwqVjeZ8x73/KiUWiEcRCZWL0jxMRhg0cwn6KfQT1+M/LHD4hX2jW7cCyXWyO5ikLsgfXrpKLQF
v37lJrPbQY/azTjyDMn+3kDHI9YV5gYHPNXj1tIZqq54dFQUdlC9cgF0cmk/PyYMZqHr0EWvsYCE
OcFxNWGBjFBv2KojGyKvJbxLPr4dzqf8OY6aGbMHGU/MRv0+Y5+UUXJWxZb4bOYEYjyjgFvOohY9
9zF5x+21kViGrHP5Hadxxl+9Lqg0QiWVvA/vhebpyxhIP9atiK2WaYC88r+aNJo5GjyotOTKAP6r
P/E121OyfLktzPiO6bt6ff2J1APrKIaj7jD6Q6hrl3ormCPiQDFCAnOE+c8HG2s/RBVTQwivWaVw
WKxXe1Rihg/mGgfnRb0Y/CEQnPAHhc5tntjF3cVGycGMJHdGHqI2uJv9I+z4fbgdq1Qw3NKQjSDx
0eFSOQaV6A0nO+LCe8P9W8VpB3fJAzulAK+eQqC3cN3ec7cuAhYTkFvZUSOi0QPv1fmfvEjLdavH
Is4bgp8qJKwLI/ABEJ1JhVdZT+znLMeuYnsGgcrT12B70gffLKhfdz3BreHuNLVBheJU9MX77+Ag
Ck1Dwbw3IbfN7pCjAY00ITvf5UWx9CznAbUZqxYumMeA/fGB5eOf08kcStI1iUqJ83uWVr8Zaqa8
qDxm8GU0HeE82zZuo8FAcz9mGV1jK3a+/duuPOw7bMSQ7YxJuVtuRAyDerZSuKZa4CxQQkDjEh66
4IPLwcpDPkSTavDNCA3uwuoRmvBVhee51KKzwmeeD0fpest+pXvfxTGkpes8cPjo3vBWAEz8eoBB
CQmiuWg+CKOQZzYYgJR6FgJakEsQjWxEmjnx0teJx1VjuuQKraY1IUk4mwISedFH7SViDLnaffly
Vk1tXWUrWjLf3P71nouGTrW0zSxd+GVd+4MGUWn7ZkxJQTmZuoYyyQtCbdiYDGbJlqvspfvxNnFk
ATXhavTuvfYC3++6R2VZsZ6BxiQieWOHVlUkVGWgoH/xyNXmTk/PSc4LYJyDDYtD/cYPbJcozmB7
pzIHbxakiBUndJYaxlPrqtPf73O+eP9mSxLhKs2qvuvkZiaZN+x4+OBdFqPI5G1aVduwh6cgjRzY
2CJnq2ZQO5LSP7mzYEE0XYiIbw4P51fQE2gGZKSGYGvJy83NuM5OM1Gs7ESzsCMLqLNevJa/jqsY
9BaoCHHXopExKR1AKNev0n0AtkoKQ6xi/AnMNCFgYxXbUJJZao6mIWOqlYmuEAgdjzK2uWscIYMk
DJQiVPJf1YepnNoXJ8OE8l9187VLugVrdvtDhKOXfZJjJBSTdHG5CcSOiIpu8/P4NUde8IqUP+Lk
W5noUEF8OqWsZ0N7ulouieUS8n4JQVPHIgfre9WAnnAYBDJAIzu6btWIPKe0E7OymIPa5QOXOsQE
YeDAK/mKk/r9xrGlDxCJxXX9mmgE1MOvf9I5SQS9pFdL8KjmQD0aMTvczsuAMEsjrSgjE1AR/M9C
sGviPvjbR8xYtRrCKdje4Rt1X97T+OozcsRDlS9TNt5PGfVfEKEiRjVZtyGgukh+z42ePPPS2DED
DGmSuAsLXJWo0WNOmLBwDH3KdmwX7idR0AGybARXRKluZ+mCqh1GR4e/RwKHKzPui4/Flco5SrWv
oFHOBA88nIL2+j3Ygk8fLXiAZ72uQZMt/jKeqzISc6DOP8IFocoAR6OZoI8Brvmb7Ayl88Y9+ubd
hmNnfpXnZSSTaUOsEetv+w4ihne9eQtiv67uH/Ty0jtw/BP45QKq4gdJOmYKtuJQJzHwXmy4EwVJ
kjkasDlHWowzqfZ4QGJD2OJtYmGVL7H86HC682OPS0vyafUhUnfyMwO0JVbt9VYddVq32yNDCKtN
flG4syY7MiMVAnU5eTarX+Kka24sXdZ4TNLcaHX1KLe2//LMV6xF8S/u305xsF6nKZv9lTcEr7LW
1C4qHdXDXTtTJ7tU75ULiqaqXQYRZ71I3qeNT1ttTqwhD2s8E7i/Po+W8QveCQElTfs6ZwRLY9uV
T4vLpR23oCKX/0c5EKcbIbSz/fUOdakpDeJEUcVuOxDY9gx1t/w2bchMXM1IPM+88N2/F4ofo+g7
dXyB/Ov+M81TKuyAsfPno/t1YfF/1DjU4roo8TuJdx4UpgqDnXoEjlgfMx5yYnSnDcatwpF0FJTR
K7McowDxzvxZqw8BeQjLXs0yP7YM5sJcq0FeBZmkfJNm29QfFPbsH2EoKk2N2bm47cXDGlTtZhpO
//HULhPd8vOY/vnRQF189KcpuCtGlSspfUP9THk3tKN05kYj/pT93WPyfeWVsoT4sdF+EtxplIQm
QZLd3wTWsY+K3l4pT7+BFIsKUxRW+SKP7kBpHAlTOfTmx9M5IfuEAy8srRUiFu8jsWDhL1tP3uHX
sjgBSMrTW6eOnNF+mVmI7GdJJigsY1RDtF4+OpXODufYUqKj5j6Z1qyCGRXXZ2crOoHEIiaI5/Xz
n8qB5pcxEn1F8dG7EzA8nd9OsHuom8OGjTu3OO4YRbhEzRk/m9rjqJlfwmiYU8wAgANWq2WGGx+V
wOA1zDXenr+ykIwd6YENRN6P+j5XKw8isgzROHemvpzmCZ45O/0M5PatFV4KpxBYkYGyXhSvaX1S
QH7i1Am4adapB2LCdlCHc0JY5F5N4CdirpXJ94U2ZRw/tDnw6NdtGIxlM+OmYQMgXf24l5rArj4P
S7TG+zIwwL/R9HzsekC0/VWqSxAwwjle7Xr00iJa5Ex/h3xPTuJLFm/CjNn5sdHn8ruJ1leQkQIU
YHsWCPq9XBGuND/rfS/9rz3mBwrJITG77lgQJU41WnGdBuvmX7RabnDt740ZW4CmLT9Fnpr7rpzH
0A3YuDNgGYJbA+AXmnwSenc02knV4cMC9Xsj6aD+WKCLDZ9SDLltXEJ7AVLyjNWKuhXvxu1zJKWI
y3XBEj5+bF0psHb7naeOW1q4dFS6Z+/PrZP4c0uUfocv//T+T2kcZaqLuSqyH16gpPvDPUJJlC/F
JWYGLZSvPoivlArONjVU6rfTu4nNdfK1dC8ygcLHrOCdtgQCn8EeQgIQWCpvQzVTTa84SBnojTzl
Wq6bxWCF2fzdkJBNbD4VTdbR5raVUqijgwOSN2obmdqgked6l6qRLku6sgZiQRRbepHQLfE68qFu
HhLv20/Yt/eYZhoZD25yWUwFoYzAitvjOBcGuHaAjpFT/qDlC3tGhUpz1I0BTZJAMCsd/dRrONh5
tGJX8pWjLWmEuRfEVXLoX29mDRHZXGwKkw3vz0qv2JGdb+wIn6jWkLAkeccgR9UehSGIf6n64kNQ
3BfTVnXAcpjw2hvhou+ULxNxC4af2L3us/YEdBom7eSXIyypf2Ve68+yqtl89GRsy83kUnha27Od
gXfoe2XVFfDxHBP358HD7B6puYQ1zqPIJltR9n5MR6quOrFBlPVALYHPO3aUc2Es1McBccyrhLO3
R8zHGiuHcZVMdhRwetAKyxz43ygiBuifuBQAWYP7i2/1AISXQFTY1Jy/m6AaZna5JIUsOwowzMMI
NmsqMO98Xus3V5a72M9XWMIkAbyKUxkn4Kes0+ZAuwSx0AwcGDO6ms27XLw+cdbUqltASvX+xN5d
Rf5pu20sCqjzq9bWQ/t+vAQf/9dX8cp4r5D1n6pP2riOjpu0/cFvemK4gdMew1iySvzP1B4DU62d
/TChr/PMkSAdUiE75D8CoTCtjoWWQbDZ5lRAfDfLlXVkqTbKyO9XOVRLFAKz26bRHAxm6pUiIbn8
Ybb2QxqvTTW3Sfp/NcgjFRWZWUfhYSFPu6uWRQnWF+uFzMJDIpT+aii6eOvSfcvd7e4+G2FfNHkF
mYJvTC20TBsOSZkAkQlATFiIl4xDuqYEONl4cpzI7emfZk4Tlc0H5mDnyUV7eH5bOnCeYGD8VDwN
BAXVaIvLjkySBCtHsD4+N+EnKztqqJjz0g6i7ZWG3Vhc9XtogYdPcR35nvddDjHqx3KiGXsCDaXK
ntJRHgDA7knNJwwMqKmJN7CpRUyfhlMyZcsNe4M/LHH0M2/2raBgZT81qqnc1pLPvMWm//XqxP3B
cmxTyb4W6VyJ+SJeMa109QivtcWuBF2HYh0boq/lY3Tvrcf43A30DowhD1+Qy+GELpzq3mavRxUn
4dqVwxyEJMuxS5ODF3laZspu9U19nEMhhAevgxJ0o1nQzp9imOg0ntu+JM6TY7r51dpk4EXUbNBs
hTkfvXjODHvBntLdUnBZbP2pz/Bm2L1dJCu+i0oY60ELmAYhn9Y6+q7eh8oJ+JTVyTUfeIrVWR94
/GOIaLx+yIcu1+dyvKAjeO8mUEKvO3SOLTXEJcRSSaiGq/VvGwWKJLP7oxCXUCdewlCB7xjTKyxJ
eC/O/rJzPfxqaQBoNibVWUyuWSQoTl3RAKyq5a2C1qK4Eu9GVdfnyyRpezGSpqaCB24hfjEqlhxK
6Fg+hxUzML1jCpKYG6Ikd892Ru88Nu4YM4swwPQteG3YjPvSPFRR84xJzd/HbnQdiVM5/9jOecZL
Yx+14eqUjbvkh3dmadUo4ZbCJuIs+RL+MNsVCRjjN9SgxaxKqcvrcD3iC5B+JKgS4nfkFtxcQkga
jHEdxg4TXj8qDqL83fLz9BYeR/yWrMWUKaTELMunJ2eU+NBfw/iDbkBUCRrlgMNAxgADypF9mB3k
NPrdUtNgF4qsfbfVXfhZZtBML2b+kgWe+wN+C6rK3lnt27z+fSubc1v3RvhzAaWXYE0zuoH+y2OB
OpZUuWYW2JxXkNqyuuXTvOU+XKBxzNizPmltlqZw/Hl0cEKCi9lFCyB7UXAJV84pKZHK5NF2t+BK
vASPjg0m7e4W61ISpR/RkJjmpHp3wADZ03Nwh0ulohh391i4bsGtP6hMBgiIAegQMWcKseQKO3QE
Hap38XqEBTQ/Wc1i7EBT592LPh4/IBqVmhBQnoqLvbLC+TRPg0P/Sa+9vTSxLqLM3fKerOBQPnLT
eTArZp2Qbrj/cAYJzpGzc2ikL8392F1B0RIhE71uxMocm96AO3XWrreDh0Rt64513x/FmYlTmkw+
YXqGZsUJCOlOSH0CHj44VGqom7gQCfaszsnRxFAO0WCFtiPgPGGB4EucUL3BIzxL9MWsUP/YcJu9
u01swLlYGBd4501b4VqBs9TOA4t+AF3/XlqzGfPZ01dmfo2m3bUeTDwZMhnlCx2GTc1tId/qyWNO
8ewxuiWK+NNhxYTph5OyeEx1OwF/8BMfMARLDCLKEpuTGniElpvj4Xj3r7TqYPVQn5JSG/oHGZjL
iGTllKn+m92fo1Rec2r4rw9DBM7maM1wZsM+Wv6uccEvbB8w0uKWTxOx1C871JvoYYKMPi3y2nS+
EVFKkAY9Y2w4/0N3BFA7df40640/7or4g3pdLkKFtBDAnqHyy706wcQN5rI347nJlB1sFuvhL1Dv
jZsBO28rjR0jAaUq5TG5/exPZ8vArnkskxnA3KY8RNnsgdnhkfpUsaA8mWslz0p+wmi0qXWkQInh
+uftzQUtPaM4Iuqkh4D8pxLJeddMNpa3hfFGV0wynSJTipFh/zdk26nyAvXUEArAV5vzlPhozGpA
VxM0ZX3a02Elj6fXSh/VbR/Xh/+Z6IfF10Sq+AU9ZpJcbUtZLUrroucdlLJQ1coueKy0alPXwg44
NfW4SnMxTA5YeDQzXpDLFFdO4/VGfnVKoXVE62N7BHyRvik8MRQ9iwYXIusmsvu27E1xmr7Y6NN4
NDlZDk9dHM/cWJCbbKzwz96rinnZXO/Cd1h5nVEyuFhvJzdAtnY7MCwR2HiW/3V85ju1YfxwhCp5
nibzbCW9DYyRCDl/v/i0FYYQiFtOq6kpACEDVkEyb7IULMz5rt3fGYLUcJWIHpJITi6xx/PhbR7V
j1EHtiXBwtpIB+I7cZmac8oPcNH1AnFTO7kP+pNyi1Q+Qlqxx/hdmD7Dy+mXuH2+EDMwIhuCYsyl
xL+t+YlK/Ro6HswuQJ/p+n5KsTg2FU7FPt0D1EYHrOqKWb3O7OMnl/nHOoYb1jkgozB1ruwrPwNH
IE+8C2OSR5UMIqvEGakehq+ya3XGfdLOaz5jt2zo1tfg+jJdRP1uEjpM8xcqh5WM30/l+1izDUvR
kD9N/pDIYGoa877++tJ6FXsYdCJlKxC6Jcb8emOQOu58KfJZiQx0CoUoXKUfaS7ozjc3qMiHBJZW
RprAn+1KJ0+a7qaYMCeEw/TelSViuKOPpytyNz/b99e564A3YgM+XnT2fMPmFfUGhJe20OxG/NJD
44N9aD39izwsAg4KrhSRDA8Q5ThSxhFkwQpHlqrGCJ/p0i7PPSUcL1vg4rWoOEVOy97MZV/68vPQ
h5ZfsmsPTO8AVkTgFK8ou1iQgnORyRWMmi32WT6V2e826y4vwmIF6Blu1lyT4qqmNEb1kPQYXIyW
8YfLSTJLm+fQBS9nuGvVoVLsxN3Tur5TZWUvdlZ/4rWQ0hWTwBI4d07ZyvmY6HV8uGT6uv7x1pGv
sugNepDFrdjGE4bIDGc1XeU0VsRn721MIpt87BMNkOjm3YXz2z7rYcRAIc7pqYIzMfSByViRCOVl
wFrEIq0yPxicodx+9gC7JdjQQ/XWtdRy6O5qQ/4hzt6keUlkzrjGP4AYbT2szwEFKagHNn/rmqvD
OYkAaMwaukKLSRRThtmfjvHsURVbUluITmmLf73BiE8s+OVSAhvIGemhAhjDW1832fykZ6rZvtxq
RTqFoS6pq15t2ZRe8/orFJPx2+ZxF6hEEV1ijSpWK7fbMjpcHulGpbLq5FxJnUzAe1TVC1Pwwpa7
SUXkLLs7o/0dKO/z3+k2jI1RinJ7uu2keihPNX+yv7RZ+tfEOMUmkI6G73Omok0hJ2ktvY7lSrT2
sz3pkDINbaNMFBUK8Ii1kPnNPq1YwLqADAakYWlKp3g7MidL2AdoZ2TlmOtx9PFBtf/slg/NMYF5
edsEwX0eH8WD4suEz5jxgh5GPgeWXx9fU2/Zwt7hsEv2BLaru1T7YKlD2DuMYEGMo0N2e0quk7yJ
t2rPVXRf1lros3IxDAcivnRJTSdAlUJIRjFGW9AtqiTU+0iCbgXVLa2S2D6RjTRDH5q/xfBI4ftu
0MwVYgRlrJfGjm8/s7ZkrAQfPNx0lqRVpOskm8pjgqzzfDur1T/DBVH/SFQN5/9YfifXNe4pg2Do
cJRc+rud85o6oSRjdFa7h9c5BKsCk/NZtPx/109q/AVX5VZx365kww7I+2UCRfIY4vn42CgLbjBI
iN5TDZZeph0OVhXIzIZHVdKKXeq2F7aDvIgOVHxcw4p4YtTe9rFQ06+TLNKet4UELjuATnRx5TfN
Y7dHDOUXg4UikLq/k3OOWAymbGKKG+0+9boOcPGbz5i0cjh5zbA7aQN0ZmABuXKnqfowTtX2fvB3
KDVKLu8oX3z/3CYhRbQ4cuy+qPQRpkvq17aI38MQ5M8kvEQdNXBr+mJyT8z0jWnpgsPa9zYkm7eA
K8wVEJEtOmDhcws8T+5hjoCb3FjOcTmVFMcKz1+C8XA6BHsoX4wF5kBpY4nU3WhZsocc/RFgAfRH
yYed3Zpu8N14Sv9+TGI0hoOZekVTNWqbToPkbwTsythALfqwrWIEBLdUjpbYmBEj+kQQ2eeMVTUy
ievflWBOs3rLSEoT+xW5LCbEV1SdUqRGiaF2vRdtEVTBWjN4OstoUdi24DZSu1YAPh/9VfYKnQu1
zds3T3D0EYry90hSVCDyq3Ka4DP9CxuTGtViMioyEAlz0rE3znqt921RD4wrqB1+10tILaAe8egA
MaieYULTtGISDkZ0Rbm4ZuIGnPD4KHZubDlorKYaxOri+dvZTYP7wZ+q/NU0QbR4jGs6sF6ZWoP7
Mj3rAN+V3RgjSgjO8IJltoUTPeBIvmrCDetkHZ+aSk+symcuiF9r087zLhjLAasG3EzIHf0r7nh4
c00seA+ByCtc+JUGSbGSRumpePh9WXBrao1RjlhUx7azkG/KYrRfwVTae0waO46LgePV83TUllGy
aM+AtjGsNuIiWkZQFEKNw2uSvGziUEfYw4zabpqOq8FEy384/b4M5heaaQdNraUU2bnjzOnzLeCv
QElGCD4Lz7JKElstTXJCmyvi4j+raSW3vxZAwTXRg7KGTO/q2CH3pLsHjyJgBeujz69eWSy+eaZs
P0mmYi8oCyo452rueeH8yCEGL3Do5QVNBr1GaHsLabInAzvgvGx5Bbqs4Wlw838/8EP9Q/I0yven
Pv/TNKtMiBTZZQnXfTNBsyaeA/GHGV8MyTQWc84DlgchqB96teuXqNp+0sS4BChg4mdCzOFXS5SC
2Uj3I4m96hxuBtqNEbxPUy8fxNYC/Pe4SvKIrzjnBgyDJQwKzAYz3RhQvYw9KeYQ2r1L7OcY6KpI
KW5BpD6AfVJ7NONyD/VlgM0Yo7dY42Yuvri/PvWVRU0OvFWgl/k6ybymYBLpplYUOXAs/SL/O1gI
/YkrlmdI8NkodcnhCScs8SGhGv/KUeOhwqy1eD+Xrx5LHwkdMfUm6mS4bOiia9SnaKax/OdoRbaF
Fm9JsKRE7wLWGG+k4yRVNdL8StytL8kdA/YtCwv0sI1wmBhJyNfvKOKJAJqsaOVhQfkKWYSvMIdY
yW5yMDmod51WKjy2lIPwJGzQGue7cl6mpIsgEKvLVySYvvFeYMAqiM/rwUX6T3rIAj/GqBzvZTtZ
oPV/4wjeahGY4rqIWNODFIypiuZGOI1k/gJMlg+N0PrScAanv002i0g+Kqyhh92Y2vPnbMBAhvjB
4X33bYfyEcf9Ej2l2kaGKNLX9rSw4HJKb/5J6pwfzvaKLI+AwcQZqAGWzpNjhIz3FZPCt77tZpyf
jmyNGmVo7vy8jEteAL+ChsdBSpFrPkA1tc2dhVyejLBrt6/ydR3LqIPzhdbWJdKdo4wdSwMtH7d2
Tcg6TmCNUEMAXi+qN811sU4c4wQheEHzt4SEolmfqKBgcgC5D3IqO0xfcVUVtX62benC5acGPuFA
ubow6mxTc61WWPuhpCIbjU3Y8qD6U/+b+7/JA1XffIDbq7L2P+hwEuwQQ9tZen3e4WnXgq5aCE2I
b4O4Ibym+WVXRZEopD29lt0p56VLm7fwx7qlT0mB8DHcFhGGhgtNPmlta50ubw+xtLXLFFCUABfI
HyOge7+sH2+d+EyMu10QRCJ83agXHBy0JCnpuchSed9/iqNXQfiNLeODzRMlYXXoKnzDUl5LU3+6
GTo84H5TvDzYXpPUBp7LSPj+r7yd2HrGl74ToYELiglhGNZ8O3/yB82quimzT8fs8q6p32Pt5R4I
SJzQaHagIBABQ4sELJ97P9g5n5NFwoo0+kot9XutAHeeuray+5En3RGd05HXyj+H6AXz7pZvHciH
vDok/cPnv3F4Ftd2qK5xPnaRzLJa/8gpsgnucuZwL899N8Si1ABoFksYxPM0L02J7mUyRyETyqHn
hyQdWFLTpDOgHvfNASrqV55QeGpiSa+ZFQGnmCcmh8W+4VoPATGBFL0U/4SJnwIpHhGCAtsguZMW
r36hzoqxAQCN7OCz1qVRvZvuSCAlZt0GfnlERlQDmIaVOgQ1tYFUo4HnN9REwSSHuaVFuA55iwF1
//nRj1qiO+W156J5ad/qVRuiTq98T1F3H/A6kVglvXEBaICxfGJo+zvtxQ3FaRRFea3x+0rNQg87
TKJABO9X1LW8V1e1Q07TkOVwE+dve+fStv2KebfV07dYK7GrtlO6e7b3snsMMqjzCekZWboQqjOX
Dq1ocmMCN/aT5LkX6e+FOkXkS/HEPBrZPJdCM8HbcdSCtFaHC8JaDBjJEjITC5d8LFkseRtbFpKg
K53I3xFjAN1Tf3ydRV4CoqpUPQ1zmPUVjM7VQ73WwP68YVWnzhXn3D9d50SKDqdO29KecMzuDW2B
3n+JwF6PBADDoZ0fEjmVUI1uU+wzvkEWRnRBXjha1z+nzF/hsRa+uQKL68DVe+gi4o1RSdvwyWyR
Ug3whgavKeBjjqksWC8JsZ3am4CnkoFjcB6p5Y/xrWIa1sZcngWLyOnGZbK4pu8QzHUoH442VR+x
nVvaunLln03cKYv3l8Q=
`pragma protect end_protected
