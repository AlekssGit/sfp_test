// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Yzaj+JNmgaDAGmomHpklRrLNtxUnKH3aD4fZc3f7Hsbobdl+t4ulH+l1/z3Iu+ztgm8w6z8sCyKG
IPhM44o9fvzvBMX2yNFcnH8xtJJg8ejTTtG8eP6VJmm0gBpeF7t8fmcZ4FeYPioOs7m7YF9yuNrq
K09AskW9tPiq7/nmliSqBZprszAiCoBR/mtbDSlmVQhMqn7Zxg0NR6uAaLYAS4bhOsJ/X02lwS0I
j9i+LluqzIPnebpHUAh3abFhXVope9cfTj20vUoa97p7EG7BUTndL8L/bzK0ZkOB27G7y4hM9oz2
ai1zQVvgajYYXgsYJxEN0IG1snoT3aqYcuw29g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10672)
/Jy35jcOs9kCsUefZ/oTAPb2USPDm4Bm2LfJafqzKcTfRPoN1PC/u39QvZHOaShrfeAAoWFyf9av
EV78/u2qWsiVJE2nHdP8iaB0pT0LNkFqweOCDlMs8D9izi/pmpbtHdsKJmcpuZJNtw0Ua09C8XTX
5epw9gEEVdgUJsX+BxW9gapA+HsDFcwXqOte51zqC7E5+WF53FX0/aVgHrXyMEW+H7Es+AZMy4w0
5fsSCK9ZgL4gIIyvpU1OcYnYOHSq0tvzc+coIsH4xuf5tdwYTAjMaOz5Ve2TVs7Hh6V067QanrwY
zri5FlLHNf3EmXE08wUpubK811oCvs5XIgvMGJJeJGAirX1LFq4uqw5TPhWwdOY+TLsj1H73NHUL
bWT3tjtdHhlMp57eRPfNsbnaSgEleF1I9lnZVoDN0ozMUZDZiO17zh/XjnjnIe9tPKPT09Rj1Av/
bKzHSIQdxDEq2tDt8Z1/1d6B2bkjPmBzW5H0IVf61VepJNi/oMjRnMe2Pum17AHdzpBM/tvJMqnr
TCC8/Axc01H73YBLbq64qXK/KuNN2sc7paScr0UWX3THUyRkDCIcUEfYGfCuN/z1ZsOrRNbAM5c2
TdBppX0ZKcsjWvpbFwCxOGSlWleHVs0UJoi0hWaFn4HxbQHsK6M9CfSBHq+ulrbbyWWk0bde6hmo
B/Dn8VIBYOAXXYrx5PYKOj7zNx3osciv89zp6wqBTZVlfrU1VJdzxxd1qF6sGv8qdheFKxDUc+hh
qZsgtMZBqZJeWYWTcMewB3ZwiynEODzkkqqUUmNtJKA+tzGW2JsJ55eOb2rEUDN/Iaf/Mkt/IDzM
GJlLelJTF3nHc6nUH+0F+zruZMUq0uUoRw/FwPBcw6Nyhf81068rY/TnM6IMQ/amJ1+evVO8fHp2
tjDPam8tio+iQAw9BM2/gvK4TzY4KHkVAUjqQ3DI1AqpnRRLQylEvuo5io/WxdUepF/QK0pzgelt
sfc7+QCAVQrExnotz4A3hJLU67N74j0x1Qwgl3PGymFmorJHEsIGw3JVWL102qVf5TNaorpJQ9wF
xoqTPEJRdJAdCqqdsAy2JPjgzRt9lL+ilzgErZVQ5cEZmv7/5nGssdAUvi9g76aDIUpNOrJnVriC
nVLq4FUh8pbohNXnhoxQoTG1Z+EdZNZxq8qJZjCLJrp9TIhbPZUvTp/RMCD2gmLInC/jzXXOGRpA
jBoZB+La91eJeS4oHL3i7bFYeELZIvZLahag0f4C8s4jXvZrnBRIIrPgX0q211qVesh8A73UoWSJ
wFN3/Ko6EmGPb9AHvUOlfgexW0+YEYWiEcoTo7jFlhC/uMp3qO0qA78CsrLj18IMsUSo94lrdu/X
KRsCydikwWMFlSEOkh843cVaRolSrSwqXnyO9M5kXZLIRGGa/25uOtCRMN+kv818apFojKPdSfrv
6x9yw2/RucgIQTwGf/s/lH/7iDfTsTIvoFCuP/lQnla40NgcZCuy1nmlv8Lo2i9F89wsQht2XIYf
GkGn+Ofd7/x7Ul4tLIAf514quhJX689sk0yc040oC8naiFmRKaYrxQ8UDOi9E0YuTzuHsGZXRwa0
W4wdMjCp6MbBo8ANeUggvGhEZO+1G/Cl2gfqMXPudJwmwFzNSPvKJHe1r4cPkI6BPYxOi8WB8QOs
M+vDS8yudqRG5bDJkadtxAcni3PFjAD4PksBU9rLx+h+74+RQIXlk8vRyOULsVsXGS5vnf9gV6+l
lVSwJN6LOkV8+AIimUCuHFlb4KviNH7NIktydDqY6Rc8VyMyzdr9UGpEZaP+4RX/RidjuAKkYc0J
gktVqaSiwI3bEhmwKTOxx8tCsW+rq/PeKczwdZ0paKOBhdxB4kwh0VpFBPZ+FrGh2SgAaAFv+E7h
GEslkvs3d/17t9PEOsieatfYMsDclPAl2jJoX+SO3csgLgHKrRtcOYeLQP7CYBI30155RiZ1eZHS
t/XCsyX3qNW1wik8K3tC1rTedXJ4jcaRo3w7tFnqInl3sSVlTDFcrU9Aya+kplQ42cUprfFSHGrL
xjnoAhix9JGsfu6PXN7wHqcvP1I1++DITM6m2tv/1xDvR0wzI6BnySoXPyntSaxHf1vU13BYnuC6
kFiDO5ovYyZ11Cn3PFJ0Z4YegRZ2sbNa2ttmBFBBoYiTkRzRoNm31QdTCJfOkKqV82gzo2w10j4I
v2jOOU5QaacT1332/Nze/vHSa/zhYniC/N45iMWdENqK7duamrqqQCtF2LDmakmW8Wev3oqVm4PW
IyATjrtIFUn093hZTUVgMj387kHPF8UqNylPTGoeFt5ML5gvvBfdi4wozXcubRQZgXMjhRM+3b6P
mm1kypc2ZTtKwU0BHzQWtBxEqppqNCNqdhsvIb7VXhRoInSzaYRUjl8SrqNxk0WbNGtpAFNy5CAD
xfTtUZCt7ElkyO5AdS3R5ZRB0tsiAKzoNKjEmigevFbC1Z8ptrX+JzpgTtKkVkwTr6aDaTtYpipR
eTNvC0zHxAsvUUexlJ7QirDY/HKzBcSch4DZv0h0yQO3L1ynLlJnfT0PkGu8Gi/1o7Sf6DW03B6X
jSwWHV6QvhpvdgMMrs9qFuBHaQBuf2hul+SmN+hNrel9IG6gh3jLhv2AQ7UvlSW90SbAMwOx+nEk
VjhoM/ZAHEo5M804fn941cQ7neL3nDqqltLbrpmzvVMszC2xYxAb2n3l3v3UeVDtoQmpOar4QNbh
+BAWXYoFQND/Ws7vUjeyj4heQlZ3tC/o+Dvbvsp7yK3qrgodQmeuL3nKUIh8SAaZL41Psh9FRkna
5nUL60hsIW8ZRphz3OXX6rbyyu9kE04VsKFvrsUB2xzbCq5tEnSHtYgX+SkmhtPimAB4/niGMOGd
MC0/Frj9csusrr8bv4LW6TFTHz29WMS40x3FxFiEkQZu+qM1FxqbzPRPnulYmG6f19tKxgaxwDG0
/sGZQpijCeCRxguKS/VwV6U1Lh1mScORWYPZgwxUnandMg3i1QBNFMXJjX+0pXNRFbtEK7Vw9+GU
k2pym4L26xVuIYpIx0GnXv67yQrgaAL0oYLCjKl45ndxdPp+J5QrD9vuMzWYLyPffikm7FJtKQkD
CKJqcHIClIQHxj3VlVQ0fTKqzTsPBNBCd5bmYDynXpyvVdw+QX0MB86kh2JM6ZNFe9xzMfxbOOmH
J950AIJZLp7B8NmsnWWz3rPoByG+IdgtkiJxuZGg6BlKFVE8uhrySp3O0JQHYjH31v8ZvKuh2m2i
bXjjOUT1e8MKkLLiFc9hqdlaCzqQ6Eo5MNbx+j/Fxu39Yrm4csj4/qqbE3DlrXfuIoQoIDgFeDt8
ZtyQI6rJQRGJJUnC7KcjrJPNZUZ1yWiaFxfHivBx2hs/HvVatR3MhjTzWWpEmyrhsXrwY7vzLWrq
zb/pGLcRxH9n8YgV6TM3SBxOTW0flcCS7mdIRsgtJWm4GZ/pTACEKqP/fsPzwEbA4ccQIgnhh5M7
jzEKi5b+TyxEq0m+FoKZL3wXHqgyFgFS8d4N7qi1PRCmkyeGDQr/ZgTQpNekKNgJlKp5Ahq5/hUQ
G4GuYUZeZrT99zhCNpIEmu3mE6Px7bHmDa3+bfTqJaFflvaBRnVZ8NsXwrRIdpNMy6EZzSODP5W4
FQGxgBtoKS5btSkrioX/edKPPlWWYZE9p4vXbYK+mtQvODzbgO73vZI2ZNGvnmKdVVXwE5+8u7Jf
9f75oTKWFNLMl7iJzWh4rvAuIqIRY/s65jScKhfFTNmeXmMp75YPjX40C55MG4HZqMZ0IAAq/GeX
naJdwITZPI0+qI990sIni6N0ocJawVTribsOr6/mZPmFH4TySRmnABMzcpn9o6w8XBsZKVojuXzM
PAmc/HtOFcDDslA1wCo7uDeqHOrog4YjkrKrUz9JyBO/awYMftIeu2MbbKdkjabx9kYM9mrxcuRz
HfZp7nWzpvp+Rps5jHb6pkHZJVSz/gb1yEZvGwcl6fIHMinvp8KYhALEqw9ggXZYB3bL+SEymd76
3Mz50v6wLaYJufWPRv0ts953MTNBQRefw89XN3yyRvImfEQ9CXAZmTCTDf7sa3Pw4NL7psoLiN6W
X/bZ3ScuT4AeaNI+SggSfdj3l3xFaUmfZI8fNTPUMrDZhNqmRl/1rEBZWHQNTOUj0dkjMdtjXi+Z
zmojvgd92Urg85SXhWXDBFu+KF0FRn2x7QHkXBxn/lF9oQBep/T+QM8y1EB/nE8mr+kVgy8YbQgj
D81rxGfn4sL1sYAJkTIhXIpCNKfV8uGmqMeQC8JYHvndKGilELTzKxAOb17B28ubUNVCB7btgHs1
aTLTxml+6mW1m+/IhFGz2MMvim/E/ZPewKEgjEsYyaNbk+DWoNSzbGecYtLL374knPnuZkmG8yIJ
L0/yU2xsjVoW1BVbKSEp2GNSlg+Gx1/Hy51Z0QK4q/dVaqL3CU8BcpbC0f2r6IK1q7wjJ5iokYKJ
X/5FBuP+hNU2dv2txcHwjxJzteHuuhN/i1cRwYbuezdWfXeSAJpFtEJGAubd3g9MELiKQvhbZ412
uAaP4ES0wWD12MFpHzCnLjcmxs5z6tX4dAhVNoGl1zN+s+bX4HbEgjnYL2HMgRXuHFFA21AgNl8+
9u8BJ3SmmkFwF3L2u2YU2+PR6gsWT8DtjiOgEOJ14kxqgz4LwykUoxZbyj7bKeem5Y227mhwisgj
Z/2hhCrpOtjhh2OrV36p+edq7gImLu3iCF0xVgmYdOHlCtmLUIXc9lcpLdjIlIenxaHKx2kjB2up
SDGo2CW+U+ylyUYEZyyH/vAZMUcwExtsmjubl70gfsuD0HPLBP9QfNIIh5CFqj2raUaWzyB/NjPE
CSdpqI/GbVLSS8zE95Sh2UUFRbQoZd2xtu5mj0pyPQJ/Yn+pMtxBp3IfUVk/Gq5l3KXqY5nt7+ls
JzWp8V4XGMh4MGaR+T23tCCi7tbaOYrz7tvDYrwiqkuBhUV7LzuRvZ93+o2MquQlLJZwmpKZ092w
S/3gU4lgFFTF1LSTsi3KKZigCTG61kRB3aMAMSsumq2JORo2R6IrVCq5aXj6BHGwMq+jKbvSX7wL
DkS3x+dq0ZCpxb99/ofbVNAbN5zPSWubnIPGkImoBhdcmkX7OuG6ld+v48GuIKH+Bqi3WUUsi7vO
6jLz38eGuWsd4IKztAbmDMzUUuQu4Zt2reFbR0uHuGo2rOVkB6NIn+J3p5MbzJDP+CT9NMfSr/XI
Vzd0BJMv4E+Qfh5n848M31GOHCwmihaNbi+IPwEeTZMoh/2SjW6erILrepij5pYxnglxrsWTnaem
1zRrbhqGYzBVSNvh0AT5pgsuYd/iGInzmW+z2kNZIW/mCXxpy3vkmqczPOh3wQdHZTIWSLu0UiOl
4WOrA20TO0u174Pd2GSWN92X/RliU47jUjRj0IvEo0wJHRbHsENtwbdSnRvwSrIVLhhu0Cc0UCv9
D4/37e4I4SOBp24Ybhouf2KPpdseeJpHo4NIa+lyaU1PzdtHcKQMBMnTI7Ik0qb+7vmRVSzil/nL
IautkavCbemf6ciTG4iCfMBYyO1DZpcBgceAHFTQJnUd6xyTJB4X9KLatmP8w/voZK+4EmQ/sJuN
9w79WUovs1LrbQNCLTn7pqRQ1ZJm09VLBiY/k4yc3z3MxmtFF/BzvvZY5KOZwp6GAwWQ2WY7nsS/
Id1YzKebXV/q3a054LwoTBGGh1f5qN4XIS/zxsUud5RrVauxQNp97JaB0p0KKibh7zSeOPl52QD1
3vcH8IbgpTYrqEjjXg47fknrXRykNQTXdQuUZTTzKtx7mOyuWni5eir6UFDcKMyYc+KgachKXUI0
RsW+e90oV1K4Phmi/nQhPsPwcOqQ4XvK+u8WtAQqTguf+R9TEYWCxfZrwZgHcTXasfD1CYVjaSxV
0+h2+RHpxvySDSv5bJwThsHtePW38tFaxJFpD6aHMZzxBeiqYYkF7W3AEntVgVKMn3f7AiO9lEXK
sgsMt5ZBKXN/wtDfRky3zhw2pr8TozNAKHYmM01p2235fHT0BJtkIdESIuRKugv6MCCfI/MyLmLy
vWSGiw7o++0LSR9MjUp2cyyLZejJoF4yRfAGCqN7fLi50otmOavDzFcJpQc1cuVaEfgzgY/4SpCE
HeUG/W2+9Ur+voqSVpMUD+dDxTL1McwtXiL3RZgKlhsYaAr8LSCZNF6jmL1DDg4kvtAmLgreedUp
eeAqT2h3VtQQlllkqpw8vmKShPFjEzGGkKZZLBJ025Kg20G8gmMWKGcUgV7l7RMuI1QmUo0gqRKA
eeE2jrn0EuY5pnCaTTQm6rh1EmvrHL4u/QMfduZuSdqLGOWl1iv3fHnb7q2R8s+zGOKsqTEEEXjD
8cb8OcKkk9hj3YuDCWhfcSdKInHHAMiob5HpFsNfWf2szdyRZw7+gH8OW+CqACq1RCoaa4PypBjG
92f+p5gqxxCRJ/LJJjp4xSvaFM4LM6oh4VYJJI+Yi+yuowZuYVy1OaBv6JqcBT9ZzJZAnx/siDiy
iqSbviP/J6WcLiceeEOnis1JLj3JMT4zSCnH8j4fy1/pWZw5W+3c9CVM4KFdJV/lFFPrtuf/17fP
k1gmQ3O6n8uJoOXfB3s564kcOJ0A4Tcb2edGmZ/1q3DMfRMlLtUuydyvcXvh4JqmkQR7jrPym/Gj
FSO3zNR3h03rKWBF+W2iBTiKm0oJwIBa+Bb7NqXq0iETZK1GmgyZLUGyqUf+Lk/gns7vNfaNMGja
3gQuliOW3PDOgnShTu9NaNM8ZWuB40cY41/ZQp/LWEgK/YNR4idDuqcvxY8b4IGKtuOkp2ely6Ek
6IFSGRieuZprZLuRMgF+m3odDebNZrdgeNL4r7OkA8VV20dytCdGvqFCpWm0e9Q3qmaGTGJDNAV2
mrCUcUJc6OUD1zROjd6DSS8/VwHXRpuxd7k208lb8xAhzdBpe5O5EsKsJjp+XUzc3lSNgfmAUff0
TT33mP1Dd/kfXwuJjOy5BtaY+LKpx2G72wESzWYCMmfROrjHmuh2Qg/xbnFh0jN5sjhgqPhLCcbp
T/T4w744WXPNFKhYrd/g2+QXszpGmb3gh8i2kH/ecbrl2wiCFRA54DcvWlrRQSS5Cbk7E/R5x14N
OJiCzjGZgRKOdDmiDQfGM/15yx23iazV1+tZjE6/dfvD2q40ypMA8KsySwYMZAoasbpPjSi8u/uF
fa7ZZJtGOGC2Ft9hLRUaYR3s1h7YQQH7GSCYFLTIAUCUQE2dpNr4j5PVhmoxTLoFkJAf5HNy4uST
/f+UNh9ScD5Ny/Hz3CLxkk0CEpNVa8G5HMJSBH3XSoRATCZz7iGDeLOfjhFliItLh1rWsEvjGOwl
C8Su2lDKhqTB5PPN8UfCTRA7JtdHc5s3o4A2G68ScihQxqiC75AV/bJ5M+sB+BwiTBL9kPzqYEu/
uk0BKDOgUc3iHCvjHylRcoJdhwwIxY1xdza/aIo6hHOWzj97bpdjdFIm5+jN5I9YexmT1q1wXYu2
nJWpacCya7vpcSO0lN13EUhpt0HSztQax0+aYvV7Er2NrGfETJalh9UDcR5YV3zgk2cnTJLkIVaZ
zZCYYW4vdJRGPG7vnt/CokAN3NNy/HVaXbz3b6NV0qS1NTPUdskrrZv/1DFKd2po+nzYPYngsASR
mnAb3B5p/HXwMah+ZhCxjyWfpeZmtHRjPUO8CDgYP/SbdEM7U3zUIirtLsdnoUf8N1h/vG1eO+jN
kJNbZxkEdhFIYBE+m2n4iF6Uc9mF0aKGN1hew4nQTCrTwi8CzjS9uVUM4STk9dr5Fz0tJ7E+3oh2
9ZPV5OcZTgdIuSrSbrSdQ3p66zfqj3fKJOt3KFOohbAFOcrKjmHtTh7LEx7GCamuclCI4wPpg1kP
iS6FYnOsHRnxrIHX8jQ7SwcBTC0INFQxpO05UBQInZ4DCHTqCFJW4QeN+jnYrnuJMRSw5cyDzOgA
N3rzkygYQnl7svGVDD7ZRnWcBbpQu8mor5+eKuuF1w5po6ajWcbiZMhR+8k5WRoag6qZRMhrhliv
eoK4YWbHAjDeKvymGd+ZPjp7Ud9jBbie/KDk7nlUiMXQ1BBlUaSsTvSfnf+TGuifNTdzxUqLrQ31
zdVVC+zY3nnbIB/V5FkyB6b6erEOI7kETdHzeOoR+EO2q/ZOowCKP95aHfelBGcnT4fkPbUEh+eD
rRnZB/HLxQ2tjH4e3D4sFIwpeIHrx86H/sLv7oz3ArfyMn6QfoEdf2OHhFRMvp8yAwEeXHIj9TOZ
wAPeYLvBhsgdJIityx+qIrLxaoDQK/V5j/gH/41rehgTVTwUXlDpWJEz61uh0NZmh8EE8YltaBxn
6F8Jb4x4k8zDPkags0WbgWRcjg5kA7Ef9dyJwXFn1sx9SLx9OjyvKfxxZt84LoKP/1KZl1sex0DA
zZfrCVT0nH/pZrvFV0Sy3tRa0TQPzPhoj+eC8qL2kDumHnBVZW+fKaxtxbRRcu1AOD9IZdlxK+6Z
RCXW4WzJc4SdpsaIhExO1RoPMDlC5CNXEGvFBETZ2wv1Yto4osEq+O+zQ9PeDQXC1J2i++mHR0NV
VQ4UHBsCMD6ZxK7VdXogGmFwpkvk9DHsCFzklXMTEL1ULYEip/TLquAxa+BsviUZeKuxI6X0khfR
G7ytIQ6zIm8tLa23gBOfqntz8LLrkyUryJFpQUsTfmZ8VGE4UDcCnxL7qbrUKFf7DHyvhVX/f65Q
A9H7n54QCgtKnM3SGnzcMNv5VcCSMsBO3WZcsZ++EYDm2FjWVaayrqODSHDQkExz8ofQJMp+/rlw
29uMj0WBGVLV10jTc2CUbUXdiwp/VZHFK4uWMhNviSt9kHAd9Ab3mW7hj+5MBur5sRD5bTPmpQjT
WTurokLsKn/Yv1o3txr2l0ZmDh2A55ZylPldmN0H0unQOCZSnaziwSKAn+S71eCLUIW438UvuffN
jlPDIglg1p0UhxJKTNNFVO4E1DJK5Ew/W1yzNbartD3mOlrYm4zfyH/g+k5VJj6ar/iC2zjQxgLd
MPV/PSKIuuJKFan6huK36zRVwe1RJnAU1Alzmq2JaUx89pvmSSjx2Yv08AYjaAl4WTWzCOwORXMN
jzftuwqJFAxuXSINhPuTt/1TN7cX1pa4YHo2FwR7nfOqWjyYVd3dB7TlqYMN3a43NoYs+wH4QqPC
4WuXYZMv/Rj3a4rX/N7mazSrqsIQvnzIKTeccF3txANHa+X8ozAsZpRoCe9Hm/S/tQ9wRj/ryjDR
XmGHS8crbnZDYyGUlKvHKLYPtlY1JNIjh7r3vKd1EfT8aH4qZLhB7ynq8SH/0VINktZGtjDYXs6D
WuEA3evqmnfDDZx5eCTetxXHoB8+1UXpMpTGtRZs9iBF8P5qBE9eV5IePRo9c2x3iCOjtag0JDGv
nHTIHrwgKpaKO8ko3V+QdK57MRpZFlSHF5rf8BXgZBgtbTEYxeJ8hgO5GbBu9dBvdS8DI0e8S1yS
2bFQO6y1Mlw53zhKmhO5aRrAoLPO0w7RT7O9CT2K85u4pi13RWToihUmQbQmXL18ft6cx+j5s8D4
mjtdXEQ7wmaK5QcFLHXeqnXNn+Z9LMXqghkS5jz+rNrgSs6UpcyMgU7Pmxz8HbqEfVZyVJqv1cg+
SwmfXpplTcTxxdjRepXxHCswp0juuHtD28b/FyfSaGu04c9okIp2RKEaMD7YHiXU2HfEi0Hg1D4j
3SFDy+vMcLhptfHjjFj39ohCjWurKLLLlK76sVfypbuJzPijYm6byEbyWLh9sf0HDvdPWZ+LoMDB
PahS1Jo6BqgPHxa5/LFVAd9GBpcibAO8N0GyOria1Yn/OYKOCtkE/9DwoYgD/XH5NVJzPRbal/sx
hNjfatQCmh3M65gTtMswrcoFfb20bguxCUNgxl04o58jrNxiWjb2tNZRWMlaeIDpktfBy1GgZTYn
a6s50bDqpm4Xbq247L9+QuSKNOc+Od6JqyffZJ9gBmSiEuXu8yTKkTRYa31F6pPnssHXSsPXu/mi
zsVs4Qj/oCxyDhSJ3Ak7ZlLtnHqhPwv6fHugMZw6Ej1giC46WVZVsX5jyqlkuIQCYVUM3QBW9Rlo
kdymTjKFEnOqr/VjtlP0ash0XEKqfRMuxJE9JyWkyraV0SQR0WbB1u03hctLBEOTdgsGeVNcK3F9
Twe0kmoHX9TfgQVVDLRpuMJAeydEgf24zQBLidxHQMt9nyutvVzwI3IUqaS8k+DYz2T6AD7JZcwO
4R/G4kZGp+DvzQsXv9mnxKIKtxZGp7z0vqdZprvSSN6FQU5BvnwKU4lWkkKLugIAoI/bJW/+GsZR
pvmJ+lstOVBjARdXnrwDyydNCwb/Foz2MQw2iJSealc/kRQh9WXYl0SXYG+S5tcTK/91yU/1ejL3
nTFZoVrPY3v/Hv56+lDaduWPiE0SUK0QXye20iasQ/IV6qpAoO4I0Lo2jAa3CS2pBMckAI1QHIhT
chFnJiP++91tufGNOSlF7tIPEMEe8JADfvsS4H+H2IckTVmGSSSLUahKELA91J54YcUcI/xYrzFS
Z4Y26X/P0A7GCcxslSjff83P3FS4hGrNumdYV67g2zrtsLcQVP1Ll+L7EVUcx3VnpwAIU6VOkj/t
VYQkxQj82onknJ5YFmQ0IKaD08ExgU1+VzT9yRcJwtKhJRBAMjc0TmLgprqxeJ6oBRhmJ4pnY/b5
+FZyJHWDL9YAZiKhUw0p0tkC2NqBHB+Hij954moYg5ynEIistQOpylszdrX+VnENSP9Y3a63s4di
Fe2HKLHza9U2tDN5OhEvToMGs4gh61mqLb1+XyHfK8A56iImqwe4aRyFCvTTb92ZUBraAulJl70j
XeieA7du8h73bGazyCHtQRgI3dCYodF4p85EWvvP6uw6LSV+vWb0a53njnocO997J9pj2NYrFEOi
18RWLeSSVUcvPi68inOxcTmWOyNXBE+9eA/fe7/HPgrWA/YW60Pp0dIRSH2IhQ3mbMp+LSvswz0O
NSiP9u1/FVqoBAXZr6V3RBrXziIx7Etvc7wiMiWf2ZJqYzyB0PT5G3K2c+E6Unv1xoS9GoxBAshs
hzzqTIUGe4wtBgN81ONtein5xmcSIxJflrI964XlJf1NdETkCaNCVHLtiM5iYnRSvOMsrYVa/4v/
SYZ1J5l62isviTxhZbE+z8Cs7zwKTYPsZ1Ve2mJNEiFeDXdgxFD0SvrpiYp9lybwnpT3UIz5FQZZ
SC+3WX9GOQwQVHdT7VIl9koe9HDeY9/NfKus+uYQeXOGvtgP/85GPpln7ZZZ4m0pfev1ij5WB2BE
uCu0PuLVF5GUuMJO7TAp8nyNcEgt68tDqT8j3+YHnrPVlNcE7QvqZ/U+KEedUCxaZlkMM8qhxmFb
+CMKhLOerQ5qM66bBlCV/oKsmLTp8bKx4CZxa+ggx+8w22oOihRL80qtdXsMKQs2/TaMDCKiz44N
6swLJI8CYCGy/6OiaTfeiqT1B2txl5uMsJ45JIOAo+4bM9XuM22s0qB1tgrUb8nnXMdI8RZ4PLLq
p2SZqYOFjAsZ/U8j51W+S44Zxc9xDyovBVuDSpe/Cv277ArVusfVugdnRHi0mbw67z25MaVPV2/Z
v5Sxl2UJarqWN5kPayqWNZVs8GwY/yZhl8FpU/ycqEEQAnAvWYGWBEgHxdQOdzg1/lD32+C4SvlD
8H6ve35v68NuUMSr0kMF3/EmX+HSxEmr65UOILbp/ovZ2o9mowut9wyUh0EwW2TfQOnL273M+2My
Nv2oghebeEl88LkWdv8kNireFsndVMQmfWQXpqVtOqzLRpTW588wHrAEvH8w8rHhrCATmh8mEnUg
7+hZ5cpEpBcx1P4yByrk3BusjVZE1OgnpOR2cSBSJcHd3vmU3m1evTMyMrwC+3raGG4LUofpOtmy
o/rcbN4J4pDmDw/nbjRm9+0ffDVE//GxrCJp34uwY8seNvqgc71X49OOuxh7TZGP9/oUEFymJP2g
J7nQ6BBM8xlZPxsggArzPxDw8vt9BkLh462j6BknO7TjF4aGhMxWwp10/cJVzNNJt8J+gbMgdV56
PIFusrjANKf5sobBRW0vgIJxf4bAt1ggDe3sCYIL+wAR+AtFEXaafvr5UrOBd2zcXT84FSmoXzfB
U3HWu29R8+FBtsP9G4PCXoyKqT2Rie4RwLdCS8YrbUeJn6vYRNMRI6+FdBG2IOQWhADO4yJHuC2C
p8WEHaO2F6Pa1eSfBaiyfNoyEC9k7GDn7cn02Mi4fyo/t5/aW66a5ggbLSNC0ba6X0j1UPOcboQL
QoHPTNsNLKI6ZDkqkso12FkcqwStgroNFmw8A/RnG1c41k2pwXUEizgCl6DTrzERXa+cf02O7VhI
uPm1gkid7E7z7fmZWmA/qAN9EKDWW8Stojbv0t1bQUiDDMrUfDHRNRqLuy6jKdtGXyA9km/rQLnD
dLJkKChyJxu8OS1/lDOdJRjMDR69EUOqpu1uOVS9qN5WZHt/FdDTLa8bsBPb0wHtrWBgPCiczq8P
jfihZMTLIQ5LwzjVtpstlo0lUOIGJh08k0CrJwFMgGVSQS4YA0YwyBFFRHA48fe7kFwCR6L0clMu
WIY0ocIERNN/mQbUoelEAaItkqCqqtj6HUWh5P+MPC8lg7pfXPLMIma8bZuSemn+jEnAQyoIule8
7/SJUO/FnQnEHh72V/Vg8HPWaf7QReQfMaKBb393hscxZcHR8YOGZcT8Js8sD8CEiratH017uPgJ
ZShY5NbV4UoxGgO6wQj9l7s11sqTC6iWd/KTeLf+DCTcDHD/J+pr/+73nxE78KAeTZD3rbhgrlqf
pgMxUCx2BG53G6ZVOMU79I4vz+QW8hEhejHeLXCOYJAV5oFHTKTWvh+l8QzcdXqiRgCcbt2V//Fv
MHMRvFLVbBNCowQMU44BDlQjIEdBxj97XPMStnEkyhG/ekecD3HOWj5sZ+KIZwWF/B+H9ph6rkRO
qRViJ06I6dAMfq/lpb/ZNkYzFshQFnJkO2/OY7Vkzztuj8sh+k1imsVeRkbtfS35/W0xTphjlPR3
luBtWbI+b0GvZ7BCd8f5IfilFahB1AizIMdev8FoKzNuhPU8C23bI7C0781Rz/dSGfTeLox8Tb/r
lcM4CayOvkXwLYbc5MgV2yzKiEhbEnIlyHTI0IsP+R8FPJxU51YnTx2mD3Cxt+NhnzCU10j4ZNQQ
bPPqNawpX1jk9fv98zBLh/XvuU6OMWo8KCAEAKt7UzCVYj/BkKJDeCy7NYl35shoBAvJO4HgJrWk
kRYUgEY00SGLJaUi6iAk1CITs9GrfSyEGtFEH1BMS5kWSVaw3TfHx4seFlHEcq6O0LEaibNZXigb
wCfTr3ubDKISxqtwUXG2n28MEPRHQCM5inE5Q/NdxrZVXh5+0wzJr3Y9QFZUZKSwDn92+j6AXmBY
IBdrA06TbHb4Xw4S9ZbfwHjyp2S7sulHtR0SgHfHs3kvshtKS6Flv+IaANNakmsOjlRaTF+6Z5b8
iSFyNNcQo4CKCe26+k3vdKqi4l7OGDAkBLwQbPwQbk5kbe7RbC8fNZTprg7cmiPxV/prREshrywf
zfGJNcpskjnPRqi3WFx9Ik9k5xW2em00j7dED8FPR7lEfGyYy7npKOO7TLYwBvdxN2zY+0wWexPU
FSJy8HFEdGl6pFsh+WiSOKjidwzdY5LBut3OdUnIjrcNmG5oTKchKWZ1kTGn/ZXoIXZgRkJqNV3C
uWk02kU8ZbpRAcF8Z9TsrzADr8BvXZWZdPSho1BNNIrfx+k+houA66/Hv/uVE6qONASfOvSwQr1o
vwgAgvDyEIXYrCbZEhlzCWQLYoLAaxgi6ciZgR5DSmnR0tMA+vmlaPYXF+qcvH3VWBjjx8QZJgga
8RJQ3/NMa3mpldRACoxOJUQM4BcpxP95HtxuEaK0tgtKXx613UC2Aot2pCMVB1O7bcKZw3oIrRGH
l5vRLEYIWoR/2PPsbbbqSRZtb76hEIUDutG+D0/PUOASx3jLDOFA1N8fPh3vmF2lAHyb6DRoZ8Ms
JUNPiU9GxceAGUxu/krPmGcGbkiU61Skpf2qFKnGZ133+qGQflf2thQ30f1bzUY7wjw1PHZ8rQa+
Cd6Ixyp+GyAHunrKAk0de2+tfUfyVzQfkVqMjIPEDwR1FSomeWrEH8efrn205VatWfj91h5NrwAJ
BK8+CFsvOYBDcaVjgw==
`pragma protect end_protected
