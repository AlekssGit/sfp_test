// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
msj7MA0tVpGhW6h419o3Jmo6+FUjFUaHUewIYpVRoK5X8/Ynp299nc2sGF+9tUfS
AhCSFAF9eBQHg8IysoXzlJh6i6BTdGUm9cWcOOAfvOfMx/nSELPABsBMYGdBy4Pb
6zsJBVZUOONEB0OcYQOkVUK3dtnqwFTsFmT9otcrI9W8Bn3EzzAAaw==
//pragma protect end_key_block
//pragma protect digest_block
c4xM64CSSuohVhbhLOVlm/vj+Bo=
//pragma protect end_digest_block
//pragma protect data_block
H5jKOEIiajCF11RwzAc/AwnKufZ0dK/dd95z66YWD0r+tI3do45C60rwX9bBx1rb
/nBGbEdg8b1tF3AqBaHZNUH7my0ZSsKJncbTKeBS4PnkZIjQLGo5EiRKxeoUnxOY
kw83hb54svRPhS8C8O7hntmJ1t6HKqDJ3srqzjFYIIgdW2u5qA2SbZSGwmfHFKWH
yrLQYHeUZ4raZc8gRya+YcDst+K/2zuKXzsI2HcRT2MwaW74rTGp6u1ALtDaou8Q
k+w1ndZJ0Gdvj8Xozm5rsk0MrNutebpN1kJPdK0qCcjPcTVPplEU8u71wMZ395ZY
w2gkWWzxvvoWq5rAttvlc0DuOwRa3w+40o2KR96xULxEF8sTdB2w/6A3QJ5tMtac
bmgGn6yhyrdGZSzmojS3ejpmH7Vx0cf4BKbmHogz99VBccmxt8QznamvOrJ1ARA3
7Y1M1BuTWGzgu7ktMBirn2uq4Q6A4XsVMnTQ/O6u5gfUx3Ryz+a7gdEeYNbIQJqh
3nFe9JD4m+9uirEV4wqSRwzfZtL/rRGz19xCT5yk7iTDWSiNgd4pVRFp7lCfxHMH
+hsh29hXJzZXKmxs1+jhXrmhpxUnfakVN75P350LbDB3dIhiQ+SwEcheT4EC8kY8
hOq3M+z4UZQHIw4MkkJ1Ktp3R29TlupSZNFeTzHPSKtjnpW0w1n5ut+JH97ZWLRL
GsBLwlSc3xzqv4jG9WFO53k0c9yvZ92V5mJGrfXj/9TQRcKNH9rCPoKKctHd2B3m
cTMLlLCn/RobpHDEfm3+sYbno7mPYYmSqgDA4qWTgABgpAXduNnZF7QJ4G12id4V
joCgto4+1aUCsPmy0O5A1bXvukerfRbOiM892MomU+LjHyfAh0bZrY/PB350gJD6
iG2oFlm23Kkkh7RwBqSHS1/imO/+Px1cakisy6kxipnWb0CBrv12GqBUZoaWKGVc
xsDcu/JxqkpMahGl68LSh8RBN3r3DlHlZQnLL56j1R4MNLQcbwHx0EY6sL9CeG4z
LLoIdMfq1U8mlBij/OXqrUV2AvHfh/BnQXzyueNoSaMyiNKRQYmLd/e1Le62vbK5
f/LnvXKDRyTYPMmvDfoxThH4Ct1emOTctyhKtktbjFsohrsfGDo1kfj4NaZWEcK5
oDy2uxAPBnSKIPkWavJyopbWcD3nxY4QtKpiJAu5ZDjVHfkGIvDRiXCulA+GhVJw
3ygD4zxodTQbs9XiChJxwOg5tPj57yROPmYPSNvRnsRF6wA3uPI825oXd0XVUeMy
hnogEn1v/vh+7OBvRZVwrAHsjCpfLODKnhG/rw8d4ivIwyVSjynSNU2K6XongcA/
6x2ZZl4Kby9rbRVDgSmR+mO2CbSECb2ai/mkhfBgwiU5DkMMQnusNMzugcRWrRup
1OK8ZDBVVVd+gJ8DNVMJKoqyRpXeyrs0k0wa2GK33xDVpxb7D+URciVu8XRBZ3m+
MatMB6o3xiS5LDfI78MLLuHd/p86fKaPDd0nTPi5BMO4rOv0GJafNbT+RIqb20rt
LGUYGPjK0CJZc1ZbckhfnxsvAxKsyLp6c1nnQT5eY1v8JWfRpynE638apVTeZ8m6
MpnDphQ2oHfH1tHj9ig1f8q8PjwVA4qtB+C6K6DPmNv1RLSLm8xrZci/Mmt+veH7
3DjnO0ImSz7Aw7E1YqiXUxpC8cTB1aGKwNPHeM7eMPb7HPTWSu45YcqObgvFh8It
c+8p7E2fb4phaAFKoVOZu7T0rIAeZKo6WAAl95NeemvcqOuAv8qdwO6wHssyulR/
LrM+HeObJUMmHr/lc8tMShKYTIRDTgRi/L+YHaHbMYLXK6rzSxfQgk/byDCApOxZ
rXvaccXgowhBTWmcVEGBlnYiBed0J47U19ehylM4M7qldwxLlZjAp52FQyieWtY2
VrlB92lPFwLk61a3fBvrwP9ojIjptv+Et1SfT/OLaVeygSfbPMweX5prox7U/637
9ZSeO9j6Szdq4yRUR13lqM6zUycfpWVwt899QKuWAdLJlUquqLzWHWmFJYrqpE2b
e4pxnIaAUuRU0yUHEjgtD8abQZ7KGoC9risPFgoCCusyKmsAUhXv9EcUFQY/nx12
lHqJiJNMJJJVxztAqeqG/YFEd+pIQLHZXzTrXyYggpNaByewD/Nrdq3trRq5KPXU
zqw0t+YvvJqGlcARtxIXgw4pjHqPoxXp3xZsISKN/AqMvbi8EEGJsI789Fo4AzwV
2jvuuxYiwb+2vQsaOR4Zm7aFpgrjlcgqYNx5aVhSo5z/MuVFe8ntfMZ/3aIakyp+
/ruRiCo5/K9SmsgD6fQkbHVH607MuA0QCGwbRuVxVtVSmCf/HJjUMHq2gN3eTkGs
lyqi5aBR+MntjUDjvWJWyFLGnoME3myL2fC+U4yYiU64eouH7wz5tSWdUl83ReZc
7A3gze4OdKl+tJKtIX68+MqikGfTGdEUnDtvu1OwoQZF3Z0J0hNkjhRrjNNa8xS1
8rCAgQ6yq2mUO7ANvWnCsF12KDp3jWMphTrCM/b7x8H/ZZSo+LQdKhJjEYrjJInT
Izojt1BDVw0aCBupGs4XRax1CwU+eMyXTYBfpmxeILai5an1WqT4tXBi1vqlAytr
fQ1PRQES/JyuJ13eRk7DwiZ2EdC7TrYpsGAU/kOjtb5CATrmj3gcM080k/qf4eBE
9dntfuAAOGCjY57QTBqm/wnEHtQLW6gAD5gO+HRWOU2o8ieoTqftn4GelvWxFwwI
HYi/oh3/cGz2D1608ENnze5KCHy0kqTOAFw1HF5xZZeMoUXB+2VcdDuKzenvH4Ta
zDNoBKtP4haryAN3kYEn7eiYng72Nbc7DLuJ5PiGoYDvSUcKo3ZMr75xo9i2IX0C
O5+OeFQVsqoYopt8gAZ0gKAgDt1NXDfrVrgNFjzCAPwikZy5dB9mUJ0dH+DZQIyP
bO7lR9p9pcfsYCjeILH1Aw/cPWCIoaSssdrtKT+dcJnZ9A5BGeEiLMoehgwSOuLL
yhsWvr6JzsMKGilXT1H7Epxf2K7EV/rVsvSlv/p3Eg9H1kLj4ZpDrJF5J+ntRNwP
sP9YJKvSp8JGZ7NQOK/4whOrIInqxHBATWTVXjvnstLntOXFcEFxdbBww2Y97QeS
uxbG0qGqUav1lZFvhKykh+5bDAdS4bVsZUcM3XB5TXK4b66rGLeA5jYTLTTbJX9T
n9+UPwDO+l6l8rnxv3OSAbwo3JZ21OhIIglScYpv67SEu1/n6/ukcjhdWDSblHia
QGJ19fQJeSLe980VSRRvctf3IpXLwvw2GlMimJ562yGVQzpckr/cr5fkRBMpfCzH
u02uIwD17uCpVJ7rjreudBatJfP5yJlfXfOni4XDJU9BV01bdGpzXB/OKeaywYk1
DLEkxw8e0aX5QhiQ5SMqq6RIAZDC+CC+cj2HgsXbI4pTNRArw/Gf4D9GigMIQVvc
xUMmY88JE/BtVwlFLOYho+Bblyt70mszq82SEt3eVeHyq3SpRGAzg42mEqO1bTSI
OcgedFcSGhIWxSMGVtFERDede/7ZzLno43UzLPzrBeqOLGZ1wUk0Aq15YVsmol4Z
2Z/H9RDIG8unxYANLvk4eMWAYbjCaFlVoMc47oKhav450YGp8OVXw74P9cyX/uHs
6mFOojYMOv/s07Las98QEJ18AdMgtOjyWLEuiXZQbGJ9VdtMRT0PQRhsC6+ICjp6
dXziNqCeEhzeVYoWG7g/7kqMHJn7pmjS+QDgla2RpuBwseX81rRSWZ2br17YZojh
c5rV6UPJev67w1+s85WY2dGA04kvYjVMg24FQyBBC4nGwEBGWKXAGa30NbWjXsK6
0XTwVDt7uLKIpiAw7Mvy+v0kY26JDPTJn0jPMZS5g/tilIsI3aeKMqSo04i9bF3J
uQkuSVk/8aLicfp2gk3QsGLudPpzGw1gMfsRblJPY1ww7VN1DMSrtDl8Dqxf6pEV
JbzYY35cKWTgxj/AmK+GGOua8LpNu2RL76YORLU61JojMctJ9joSGbdXDjr292LI
HyWTyAi976H40SXF796rtrzBzUDTlIQxd40cv+NbHpslDbDHMMm2uUheGbHH/JxV
6875bq96eTRuZykQGFNKASzZ7xnsSOiR2b937v8EJ/6PkioIH747iGQ0kfjiAtlP
cQ2G8svEezmP2+MiMBjQ0Pf88vtes9ItisFENaatNQ92vLoJP3UiU9liyep23aBN
rNnUUCRvdNlfWUZ89l/bgUDsCT8tFCIcPa+33rGZ//jd2cKtt7YEB4LDZDzaUO6m
Z4hfJVUN720/7/JXAydmGvsm4Tqyop5TGV7/hZFUtV0H8UMZ2o803orHkk46Q2kp
27Rb87/0ISmsoUCRH4Cp4w6ccJS+GK2xJGVMl6fNK5Ei+AsMpjBpji9YYqK4K9FK
Yq5VOaEDbpeTq88Iu0cGpH3R8PFB7yjhNo46r+xcF0aDJaDbjPJTZQMBl+oYUgfl
IDPtqR88qg5h5qTfNGQIId2ty8rq40H/1hUNMtqS62yf128uitfs0NwXpwWTnjDb
7dYaw+KiK9LWcINTta+AwMQ9pd2+Jjr56O3Qc9tbO/j69xY47Vdf+xGpszR1zNjL
AuaJm01yY0I36Jv8Yp+zXrCuEODBmgNqHaS88a+5hn2+GT8t/FQnlk3N/rARJEC0
VdD0VzflpNyxNzNuVcLKq0r7DIUXFbvf4aZA6tWecbOIjLPeaNdXy4fmHGPEUr/p
E8cLqv3H94lKlsI56ZA5JOxKSxghXhZy2atShymeOeUSNoZmpjdfQ5GxcUVdhbzi
JqHhO5davkiQRcukbjpEAoZkKIUGXvoFSx8AfwjVwPHXRVWJgWEuFHbdL8L90O2Q
5La/HtUo6k9fF5MowTInvc5HHOh/lxo2ZFvmHtb1QMtOXfHgUZLcMxieN3sedTrE
CCce+UVQ57pXqx60uEpZoMVlBAt+lXraJi7OaARkR+KZiLYLjgwvfw97Rr2HvmM/
UX31165od2qHuDMC/f7Gtm7X9OCH9h8tF6afRb0JZ2jF4JVGYsITessiC+LhLHwf
PpTWribS0Hei1XcMCwFST1wvDV0naNtRnXOg7YfVQdcxnm1mHr+lel9DuSpw4o2R
400vcVgMwb1YexlRT+jU5JFDkPjRp3eg8Ux0YMUdxNuE+xjpJuaqixjp6MEBxq4C
/As6pX9bWbeAWXrda6ohWb7ZKSJ8BwDVWvNbMP0YmljFtDxK7dh8CKQ7hKnBkbcV
Ll6ff9XaTnHnrpCe1D5xtdwVQehZ5wDPFdwy0SewsXEjDSv755ctEDnwApe8pcnk
5mPRbzene4wlMG7BqzcSQf0bGuP6RjHBujAfx1pG5emxIGFhz7N3tStXaQuuocxV
lenExYdsT3GB7T1IJge9o/Db2p13zt0tyyixJpa2cXTodkf3erh7dJ5ohWx/JZ+i
WnSOsbmkLHhGCkuGUwM9Db7Vs40qTlIH/GVlhA8F6/r1yFI0pcAjt95ivQKF9TJ8
dJUOnrsvbs8kClx7mjYOWPdSCEpoihESDc5t/HTJLYfCy7Gx14o0zwhP4MR6l/sv
DCGJ/6UEAnExd7+kmPkgP1CLOxKiKg/rJ+N2leC8bzfoKdJwXV/5Sb5INuDRjwqE
VE0TICAQgGCFgLEqn9U+nZaoA4wv/TK+QTDZPMY4sxekBrKKfe6M+JscvQeGm5Wh
aiqcEIeGAYdNrJMNMeetwH2W62glUd7D1EK930gKvSY+heCya4tF5oEbM2m5TB/2
XOfArQm6XYbPzBvBQ8ph/1NBio5uiknm1NeJEcXS0Qe1pyopfiXGyxWeywTCx4i5
mBbTy8c4FEqD/XFhmE3o2Ds1EPdtj5s7hW0aqThK0wzJ5umf1mu9qwXaF1JbgI6a
b36F/vxzL/VYkzb1/35lA8eumU5XRpsr2H1rBEPdYpxjKNeZvogDUwh561dBFEV1
dL60PgvBJGdWgileh2oFwcw1z3ulB1GyXvQmjg63JcYCefkSvoMJgdVublPexlYA
in8z2dzBaQVOuxz4EdX2AeMGuEAB+YUx0R7K+HDbb43+TFFZmENrF7NVgHq0n4I3
aqiIucPCxOy3vWZiVspGTK7vn7Zr8/4taIArzaYil349umHibH55LJtCnA4VvPxf
a+sQoIQryJ/8zWOweBRqj6uW446WZs3w9kKAwDPXGTzQeJZNDBFFoFXVheBeusty
sglg+MTC9i+sWhHck/ormW444yJyTiLJMaJYwKnrirOIj3H3FeXAdiWhwoHs6OEa
ivfeIJoxpuZ4M/TKOoGCKcecw4wC/Orp6QWb6SQ7sb0MkFIz8FotG7ESW9nfxmNr
6ODXjTC1YlbJCck2VkwKL/SFTTe4Tp72X3mPTMXIFXg377TNf3ssF8N/6HG8oPjw
ddvyo+WqvvdNgnfjv8sNmuwPmgUfP4MOhn7CQAqZUbRoCvYMZ9AME8+QGeyQN0yb
iUch2GLapU7oVsJm0biOtsnbfOJy8S6JoMxi3wMEYABdJS5Hk/W56THwYTxAW6wa
x/vxfURbB29pxnjJiWEPHNt3f+PSiWG7ZBS5QAUPC1QzWk+qs5Y5oA6usgwtkxwN
P5cXmntq5qpR3bz61Sn8f27jE9NedJC4y8fpfLfEOKJ/v4uEIg6t+g3QdliP875G
fr2b6eJ7wfwWPWvt0l1jz1/gCjxaIcTFaF4W9ARC2XrLf3hLoBa3mFTeR/7WHLvK
OibxfHs65GeoIHhr3upmEmUJDlWGQG7fLG5JxzQhu/32EbpXZyEUmiIRHMae0tN4
DXQB7Ljv1rDZsse9IaVDn76akT2hHGPIwFgb9I0vs/DfaJePGd7en0+dDpLAbrvU
2B13ojarSj4RF08EWHU2dPTJGpfQtEAI2U76VxXfUyAExHXSU5rfxm/4j6GTtCeJ
eDu0Hq8euRBvHHP9JfzXmaPQsomSLuuFDmPXQJxhMfC0cuxrjXIjAHEssFSyCq23
b30M0SvRDxvGcs6RVNy6W0P5a2qQf17+UQYjhoD935q9RkN3G9d0zMjPW9dZ6zQO
J6CF0/FO07oivrZJRRFBbUEqJ4sgaRvLEH9zc5pjInoNHdrnwjt8uWKYhJpiDl2l
XaRq8LbHWqZ1HtRxb4aMwOc9q42IBbBb+m4Qj/ZAWuUjx8yQOTJwxcXjjnQyLkqo
CnEhr7Cs6OcRT9ygQSOw7U7ZDS+pvgC1UKjXm2JHm5ZlbbUegUNUZlUYSlfS1x5+
YfULz9IVG8jJVYObxiVFL8RnoZtP8CKMEAQUxoS1DTJ1kKNr8xBxNSLrvojAafUQ
QK6g67mn1DFqqAOe7j0C1ZHzumJsQTrSTgKRxVZWBq7Re8XsXcU1WTC2psDP2qjb
UadspauyzoUP8fK3OumFa4y9fWyaCXzbVFk1LjDD6KStBmntRMAXf3AsoRIQe/dU
m5LKpxhYAe8/Rs+D/iZE/09H+Va+T3e3km2betIAmquSk5tbacd256r7RD8n+j7k
LGvwmrTNTMn9aSXjo8wGYZwnm+rj9aVNQMbfZsUpB2YAsnLDowvNaFhNGRSQoWej
hJ9jdTqoXqCj7y0UkPYD+/BSrE2VJ6Gb75g8iNm4f1YXX0qrhYv5IDGjI0BxfoX5
lZC5zNkCJGBiRh6OyXyBpTDRIEQ86F7IJyDOZkWztSsqfDU9ZQcBBdkK9DeqrM3K
8bKIXLfaSLsU30Psrq7lShUt6qOri8dr7/r3fOtMlfxQqklwriRdmMqRu0BDiO1R
UrWwz3FwNbe8bb820aONvA==
//pragma protect end_data_block
//pragma protect digest_block
80kk6B486sGgNo3nAwYm5vDpAT4=
//pragma protect end_digest_block
//pragma protect end_protected
