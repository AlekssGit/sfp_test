`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
TOxIx3XDx2Bjj4t/fFPLsoxk2gNejN63EDEPDAMufIV5oPoKnB4yX1kTc6E6f/I8
f6DvPL00xst5cvqkfpRuw1X63mMPl46zi0d/aVIDUGJidYdbXE0Ijgle5jDDhfdB
adXiET7BGwaMC98qMR+R8xmJchkf954y607q2UxKHHU=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 468768), data_block
0KbtGjdPOAc2qh08Da/9T6BgynqwIcER5cDf9Apsn4QYzELdCXwTkLWn8xH+m8aP
x7RTLQ5T3JwpRITOy7yJS/FHQI+joWNI8XW2tHnpqJlFtOul1yVKYhO9k7+iAQTs
J+oRvINUzqJSnT65Fz0SY7tOXS4wmZ6VWbvMkiE8AUOjFHYZrOmmbraaGefjjgw8
LKJNZV1LREOmN8PkVgoyK285KIfzYaiMpMev9mxAgNqjKWrTKOApAn31ImXSfEWh
lLyDzou/fgMQluL0+45L0Lgb/oOWlaSPJgFQZQ+vvPr9oze/ccdSNBinSK5Ou2R8
9Kpyub0GRQJtptqrgKOGfAyweG8nciN3o9Mr0JqdDFbOngWN9T5ZCMpBzzjrMMQO
7tfv5xcpeVm8mWymlpI1/Q5AktbtAE5Lej0CnbfftWRM9ubbkQSUbu2fDfwT1h3K
QUCESZvgRj6JGwJBXlgjrlUJH0vWILbwhi6EEzGHuzt3pj/w8nFhKs+wCggiOJvU
/4eUNCzQZ9y677/R3BarSlDnENICpegcTZ8VBvKVZ0OAm+vmegknWlCam/uScOTK
TJE3rLKBnrQGa80sYrQxr885ROHIiittsrpnYYg+/ua6NGWVtGwh1IRmBtaGkJoK
FgBiXaGDGHV9QyN+IgCrORVg6PlVa3ca2uvvmO5KvCSgTAOfcVp92LSCfbcfpw/4
gsd4OYSSHxXdW799YrY8xpyjKctV0ByuVqEzGwmSqQ3AxbfVU2Ab69fWBQsP5oa6
bCcjySQwg+OZ1a3HBHAYy2KAVSO2ITpal/jXRMFQfz5T24xwnBk+wMFQbM/zDmXG
kkPiEhN3A0sfFxmZxLKWoTkkJpjiN5bIhTButd4r7xE2cxYb/3otfkW7KpnAHcSc
/ObA1fpaI9IePb8WopHCyVuruMKq2YJ/be0Trr9Fp/sesaa3ke9NzWZXon4MFjvy
7sus0uHd1N9b/xFgdia6MaVVFm+m6xLR1lRGlFBEgwqolzNphBdaxc0loYUBt2xe
38DvlYdqx47NZNMSjf1LUmktHk//W8aAO2Fd/q2I5xi/Ljmm3z3f40WW24pJ8aIX
dmRTAVcrGRY+yIeLEidKzpnPEUxbkv0AR/7eEShy1xGD2CQvUe/SNdydt6E5X47M
FR/20a8aw81VoezYQKb75FPAiShOWU12PygBmj4IQ/Q9c4TyDTIzSI11CJ7HL9UQ
Yor4BBsHizCeIz8ULx6A9/yGEyxUtcprx8dyZ2CfgB5IVcFf9QhaMHlIHgoz69Ya
iR6nSmpKkZK8zESbA70vCFq5qIUJ1DmkpdrCAcy8agn0Z+3shuRVMdMJzu572jUL
NTHWoJ/NVTkMnmISRb5D08BLp6X68rGiRhrVq8jnWdaus6KbwAo47P2Zflp0cwic
XWxa+HCtPyp9QhTTK6CnNEuGu9rpP3KY6oMarXe7RGMj60h/9U+9tgwc6QmAM1cy
F4DQ7032LScbsWVW2E7rZK+ptX0ETyC/NVkSixNPKV4O7ZbtgOHlbludABT7luO2
pn8O6VLdc+EtaGcfIz0eupMBibN8wdpObl2m1raG2aEmtCaRiZwcAQ6vC3q2siaj
QVeDXPf+5FuWy1T/2crXEnyt4Kmt69/JQhlGZN9LM0U6CBmG8KtplMRN2UDiC0Rk
CwsDbWhbOfhCy0vhCDgPnEiXaulU0oXKc8JTsY8ticQ4szyzz0MJz9GloEGiOav4
U+gQ8EOdMyFt2fv54pW7pIV/ocFcRoErj21a11ZXtoqw7vz8e7oN/UnuiesnWKs1
sSHMVq+KLwMNJnIzNy6PBJ22VDLodEvpTM1SG4QngrC7hIP9MBMUeTKWBwquvMXE
L9QvzoqZP/DvFFsGWcFbkhaJPQ2b/EV6hZfIB6LeK04FN+a2RtPD6qor2mHfIVI7
Txo858kyQJp+T5TjLpBg4eiZaGOq7gXVakExbnfG/Be9xvQ7hQ0iAIEqxaw5Wlzw
/EkGGP8+ehDFF1RV4db/2J0g4K0fQKDob0TB2UfJsCHj2ocSzUbAVQ5kSf09TTgz
5N0lfNue7Vg5hqxCOnVxI2WAaipJL4pRwXWuOhddPXt7J6Gjfh6fvXI4HnoOujYW
UkAlx5n+DGmkKbA12KS4itgImjqLbPpsiE8Re+wYfBuKtF+ANqvnJoqZatJsyWVn
owVqtFAsAGebg9xiIbjqtmkC/BzpNcSMPV2ssmn/QEuc30eVsARqxVI07qG7aXut
eqRHEQoeB96X51q5lCa0yLPIm0PMjNS+FmZU9DRnGMw+azlFl751yTr9AWnJ2vtN
HJN4RCia3KXd+ZtoGNisbh2sjlEi25a8E/FjjJ2UBaTGsn9Wr154h81H9tZMbBIc
ulBqdTbdNQjuGtEXnpsafaDIK8z6eBAbAcubMzGFAwae6bLC8XQC3WLQcENn6SA/
K+6NbkxZI7Pct1wtGP5bPx6qXCKO1LBRAfN5Aq1UYhZ4tdVBu7OdEUTQNrhjo+qx
q9xFBsJkoMnxLia5i9dMEi9To8nj5nVsustvgbie8najO0JHwKgevgcJDGbW/SIH
66p0b564pYM23QSl3osCFW4fNwRu4UhvEINZSDMnbeg9CXd8LfamFeKScG8PBvEJ
8Gvw7hygiO1WOV9zTCImT3iCctobjqaRt6h6L4kDG6BYJZ0bPiW05lrK+vrl7ntO
P9MfK3xQuF408H99Oygznj3gOeeIjJq7vMP+QMEPR8JJpH+QKRrB8LHqgEh6aPqE
41uVx+vnlenVzowzXZUucPaYYXVZ6buBoYndR6KU/BruTUWgV7ETx77uM6eV6gPa
KD34ML3fHnQX9yrChbC8jJtD8I45CJ5NvzPL4Kvtr095As/AwD6jHkyisGY2d6O/
EqIf4fjLjJxERQ2aOipECRVZ5QL0prhhBFBTz17KrhbuJ3VQ1Hk+lEPIXly2UaXP
oXz1sTBDIVzOcYkY87p1P++5HfbmU0pUgfhZnlcVvb8Sq4A/R8pXSHpnxAMnGMqb
Avhh9cBuLzbUudDPEkskrZbJeADgnIWtMvNMm35XITu3kDFZSm5op0WO89K6yQKn
28i0U+3+yfl8570/Z0i3TA9F7VJ+JeudL0eolqoJblvBMigangCpr1e4Sz89cXze
Rkp6De6YFHEhg62Me2tbzLjjzKbjn/Lj1za0niiUpcM3/5rCKZovdPBuEki0N4UG
vKhfI5l+GL7XE39SrMJHErwzT+vhv6LDFhOGlS2kuiNbU5PDJ/HknPdycGaGU+bn
ac62iCZPs9V7TImPemF9Ss99kd8K/ycC7rxcYuPO8TOPxs70kgVVPwkHcbbYNMF7
ZNYCbZw5V54GlvV8bNdTMbWFfE93deTLermD9VIN+nVOesRaqSpco18dyV/UXKuw
3DZDmPpeThrAwo/41V3YydiNr3aeDLBWVGq0z+H4k7YCv69ZezN8+fzzU5p6zDCp
w0J3feBC+TJuGXKZm6s9CLSTXAgRtS7lJTvQaghopxH5lG/5uD8kDeye/1y3Dg5p
H5j6jkEZdAUU2BvX4G9I0ctRHySF1cGcS9OTehIRl1Kxs0SEE1br/8GI4UJ/+fk4
1p7TrBh/8QbXHHlHo2M+rku5263JVflasPT6Y3UtKpPbeX8bAYQYWljQa9xIlGfg
piJj1vHQxZJD6Vch3VUuriAvbWxo14LPIBo4XeeFELGIYnH8WmZuDEJUdvEZynjK
s5tlHMX0xR/vNFGOg5MMGdNBZNT8ygIUTmEoxuWTwJ3t8fSdnXiu5kGayBPQrwmi
S+Y0l9e/gvpJIkbdqF5L5IRiPrieYTll7cGyjLq2eAcxvvHRGoUebvnchZRUNxfk
WH2BLZRSvvVZsuSkuJKdM/4pq9hnQsMXGETvlnchyFM3Goi4t0/btQS3agjFGsDy
vYukGZEbL2pY1uH6mcjgaaCwr6ZPeevBIaVBaLqTcH4HxFLsUJmGrXw8vrcHHfTJ
CQWQjNHpTVez5f3vz/q2TdQsyKaq/qXVdSIvhwjI93aDyG/63kp0e6c5NExHgDOi
UqCrT4cscli2/NMSGpxKGBTm5J+Ty8fCDVZc7/hfhS14yF4hkIBZeHK6bP3Tf2fY
nSb2GCa+E0RpICqNVePa5T7resRX7OHHEpoSUXH+jU7IOuDyotehIKBKhvYmD39r
GYJpoHRTnwFIzsnidQRGBC+1UJiCF8Wpk6n1m9ZrqYzyaLDBxzjdgQaR8T9CGRRr
AfVQEuewdnPrYRPEzB+GXpNtX9c/515Pj59WNSqb411zkxu2ou9XYyqblBDwrjQr
1odXIxQx1K3uy9oF/I/uz2KSCe7U36cDCVWhozr4E0q8Jvz6uYBcLnax1H/nOgfY
PzIDhJWZ+MWc/cOJQGeYtl5G9IbJaJAOnz87rKoEl/0yDA4KnLQUrNAJvAIiu6g0
DR7AFgBA+kNeA7uvy0KmZaYJ6VScQHMM3KuqlpLUzvzbqjmKEMW5HBxrHuDiQOeF
DfJiBEubmlH387ExvaDAACIAw+EoV+q+fMKLnNA1eOJ9FDnbso92SvlS6KYATIY+
WCi19MBDJbbdseCrvdNlVEqfVfWpNwdPUmbPw9lVseXTFvvp7hTu+PiMr+EpLASF
M2jbcLgNACnI7IwEKyCUYr68ijyxcvcNMgNETSAmEdsUD+bqcZZMnZb1pKPWsqXN
7kAxkajZDmTfSkPtlMQj+elWXpQHl44Wa6/259/bhv4OIICsGgFHnHsQXBbqBG87
DWU7c4hTKUkw6zPS/cEWxpevqxLX7qV91cVw1DBOduO98IFFRJhV1xOTSO9afhH0
hjpkalG5IB11hJ3K91w82vuDM6P5xw8VKnx7rU5RPkft+VskjsB2sGqVUPwGY8Ny
oqFHMW5fQHPRBDdQCeS/kwE1h7xxdE1Wt4GXzqufhJdaLHCGgvwCTsBLVL1nZcr6
lD6GjnYZkEKq4N927eTYyjEMQ8rBQwWX5o2p0g79aMPuZYLmcktYg8dRool7YM/T
jDuA2trDmI+Xa+mktf1WL1A7hG0OaNfDPFfmhQeg8vZL8ILjdu9WHe3xdLDWtf1V
RdgV0kKZuAk9oaxWMnJDA5agEL2qaMzprYxfWDaMItlwjcgOPgkKIXetWrJYcJLh
Ay3007E4bJVO+SNjsf9akPhS93wK3iX6tIs7IfhF8BT734xiwIs0lzyEUZULwt/b
BnLapPwMewemMkeT8hpuRzmkooHWqBKI1H6CnpuWpCcLrv9xWAi+kJQ3T1QlfvHX
huXXOM64VsjEycPo4sOIhV6dSc12QTd7gGIRvYYhYdF/daHKZqmxw9dCMc28N563
4A2zvNSczNkHX5pYWcnRTajs8amZ2A1LbiBHN8h7cmnEO79sql8fuJDZo7zlLYk/
f03N3cDoo2DDkpQPIHpUPl4hNxZt38m70hQ3I31KzdJ3MVT45Wf+xd275zlHkVFY
PnPortnws4MkpQh2IbGSPBxFNJEe61qm/enPkkYcQJtjiG7pKrCAh2Y/CjU6NCmN
yOV4f8NoNyH4itWytwiw2ng1U+b+bCRqg/s6xW9F7pGX8ck8JQNd0xGojVkkELKI
tuVuHiqQUaexMwiSHG3nbCzoZmdaMzmrbR3jkskJFmK6/UXitemN3BK4BspIiG4+
7uZgDpO2IREPfV/Wk7TL6sb0OETSND4ff1tczFgZxKl6sFjERyLaAQnIee7LD+jL
5eh5U1pjMp+QcgZo9f2tL/vkRLW9sLTK6FhIXHkg1ki+8sTwDutac5ZEj74OIcEQ
2o0jOO+aHHf5DMUKg5ZFk4+R0mnC/AF6NQ8RFvBRU8zoMoCUIYC2Hx/lsMkKFnfO
EHaTHZuKNnPgluzeNUOCvH97kGU+wU8pr7sDnFTHGvPIpm09pI6y6j4yfNPi06go
2BuQN8d8+OO0lRZkum5l70WnWj9R2yqzFOoLtJNQ66CnLwgh5lMGmTOTghyu1EON
VEVH91+4MuSBayyWzbA+zHc3xg7qjU0ikZgOCxoyzsNL2VZrmXCNKTOQBhPCwOpO
NUxd39Mg1tyNgVSD7BGPGYDs8ClrYCvUz9/7O6tMfdfl0pI2B7RFbPtL1a7QOgvx
tYgBcu3HexDTiC4VuMZzHEvV4BRihFapCgC4y+h51848eLL7LuTk7kgFqWLSzHFP
MdjFUx3bsJTWrJEScVvneOsEInxC/fBJMB5wWAr0/1OvJQ9Qg/s1tG2G29OcPScF
1lXoZFQ6TXuy5kX/GDSCJf68Z53YvM9Ji8S9RU2Uy+mRNwky64j+4prLUXXh9ouA
od7EHrwstSsQ83q4grse3WKsCQF6tMkkvcDFoRhcxVXpDGxQakoITI//9IILu/fr
/ZxHB/K1HZF3plDjyTvW78VIhP8p5tUymM3MH9anUzfHM/wggJPmBLqu3OlzeNbq
CRBcP0ZYS+pv8OuNQTHRZLbqirjJP3gu8AxBPpSjPp2UyqewdCkfqufwb/n1xqCV
2iC0tNN3wYta/Oq8yAvijKJox4S2oZ2KctvleTTdyo38IrAzI/lpw5N06ziKxYHo
wel5Egnf0E0TaxDM7owP0V0TkoVQyZjL+/dscEykpTGP/zEROZpdlNO1rPS6dM8C
wdo0lP/QuRpSuI3bA+KRnmu/hupHGcKA5Okk0uE7NkY9Mbmd5T+ZjRJXAbGdycg8
/DOm5S/pIkpu73rAyXXZ2lejt6E7JGMALl3iWUNOAKpQM/E0dL/fmF5VGoOvpuCE
s2W+pFj4MZl4pRSWQAAkekLQ8ANCbZ4IOTq0OZs/i6pGyDiLsInLro9nhrgXvY4A
MsO6kxJDqAW8G7KvrmKIEI7dPzsNLFcdzl/I2RF2nAASjAk1At66Qv6yDBEOGe6G
KWZ4UhA9/A7kpOHcSseCd0xRTNKrzDaKrM9RTovVytGB1ZKFfeLesMk6B3Ftp2gg
g6/4+cANc+Ii98BdmcMOZL5SbKuk0nU8W7kJ0l5LO2Q9ak/nIjDhKnbBeeAk5u2w
ZO1+T8HzLtHwPNCgitSuKAx+KeeknvGDmlVVy+oYkUx+b5tirNBLgdosABWNqtEs
ARJXR9d3EtApbUVziABirPqhISDejv4ycE05wdCNVfyp6bD1TyrSYkR025AnKwCv
dM8LeHQeP4Q/fnzVHnQSiCazCpx+wcjeSjbUnNn+RP3sRlvqp6sFX5Tl6gPhGL+M
FG1HOGKym3FFZEn4gvSHXtJvQyCxQlQspjFAYx927MJzdsBe2lBFHLvm3IuAoDQQ
/+hqsFp3ITmHEawuF3nOT1xPn4tD8+fnCa0g8DMYfkM65K+Pak5K3Bpz7JEHFgET
0hzUJ5XTcOrmVNsyoYDA9SaJ27uzzcQoNR9ru5PkZH135WCjIm2DzOH8PU78X8WJ
eXuCi8OlUKNISSUCmYSp9makHdBM504rAsWE7eC2xvI1YmXLMjQGh5JXXbs32U+2
Xtgiyu4kO43LwyWOlgw3MJ1l20YDPnXb6rpovfUMw7vox6gB9Bn6K9nT6hChJZqd
n7ZlyJYrrC9Q9W93TiS3r5tyww24dF9quEFrqdPTyCp0YamEfWvB/RW4PPRPQ1fN
AStwo7TCeBY2+x8pt6IipiCr3OfPDgARGPauYpd6H7Hrhz33MpiL2mU8WrJOsSPt
/c4k2Yup6Ob/BQNs1wNLD1WKWnzDtGUVsq5wtD/ZWXFgzXwyUIHeJ7nSXUIIg/WK
dpOUGb5+3Sz10L3FlRPOTY3Dn3xq4yvKAKy9jpjBNORWMOCTSHfuKdcm3YZ16qI3
28NkQ9Y16Fb7mkzuTzqqdjtv/gXML+Yc9QK2O6Xw3yBoFnE+xlRW17hYiemyeA4f
omVAg6Cw+ZjyMOcb+DgQWZ5AZ+9xYTOv0To8V4T+DolHMQ0JdakSBuPqLXoxHjIW
ssDOJozypDsqYtTeadyHQnhvKS2BDH227YDJSnj9V+ojKkB7ljYQZqpWsgINm8mv
lqIPWFGlc7nYh3BnoNpNkwQLFtaDB0bcf/GHBPrrcKjbeSi/XIZ6tJiCgAv8f3Gq
a7wWtxx91kIfy7WHMa4uzrgHLr98XN8WcdS7EsTsaMZx6li6ZazoLyaLwuexydFQ
7VZXozQrqMJWzJIYQNYjWMdgYH5y7e/e+/R1+jC4XCvHymolropOQ/4p5IK8z4LH
V13YVSCRnygPrgFsnLR/R5RH5BwJNHHpfEySVTwcHseHsMp4bYOacpmdNtt0gEs+
3I2kTetS9VxfB/3syyLIRxzJ4UzdPuKQkIT//eoolpu+AH8a6pdp1GUK3Z1Tlulg
gtrVuDmIggfpxQDkRLLuqKAMEIWUkjGDvLS0AUvEqSxhH4XN8LuLZMonv+DLc+pu
zuiLDrVyU4W04LKHDnVrkcSzNd9H4h840R8uMXEeFxlXPflqlTQ5J9JJdiXEOPCW
3/pZ/xlYewkfhetmaWUN+VllX3dKC6A2tJhP5id2LaPYLtSIt4xrg5UcuF3ns0R3
aBpZq0I+uJ2qHJ8CXlj9Ul1neumYSuSgH4V6Kqxmcw/6w3Wa5CoCXbxR0jb4Elka
PMXJTU56eUJeYbRBEqXuSdin0IFSNwq7P/opnhwNA8FFlai9hKjO8/om6F84OdiX
0CAz3grk2qtppryCJI9vZFcEtzDUwXOKHinxSOJhwbC6RFjFxoN9k+4DIcL80/LS
Hj51IZUi/20zM4KxO/3aC5sxyBOctqi4qC8unxlBDlmEF4PeWhxVYh67E4FghlKX
XBnhigKQ2VmvP//7HQrzIJxXZ8pULXw3R/BYMdqSH/KlAlECVe0S4tWADnIeh6IO
EnLvAunpIf3MO4qrWe7BeVIcMJVadXRo/YdtujV6qUKwVNnlO2lQu2uIEuVM1TAj
+F5gvboYFJCsF5wHq215GKIKRVdgtN7+lSkA+dpDE6+vz4xr0V7tMJBpS84LRQiQ
wWUJjxjAH4nTWbu0wYtcrj6ByVi/8GtLJM+1FI59K94dCUf0DQpR1hwrsDw0nbGz
uj50yoHkGF6g+XJ/+cSqck5Gf69+DLtdEuobZGibaGIvB44qRJ6yTFohIN8qw4i/
2nGWv9TownzEJurPYKQnQhUksmca/CrARPbQiwhVLFqjERb6RUMgeXl2bGshfwkU
9s2jGbV7iH7er6ORSe38ENQTmFoLEq0+2qnUoGNxa5m9vnRVcFX2cU0oSw0Z9rBp
+WFUHQwymnGCjtO5Fkd9Yuk9rmy9nD1Ebv+yl9HoI8s+BU543jiURj20BiMnKdp9
b2bPyZAp92q9U2t/76T55FEInYdshrQujGUxiEeWxA6MrJA+tV1fcED9iaMhaJM2
J9l5aCGmEbA1DMIuTTkU7wr/eFsL4/a927OOKLQGUlGbj5jDFLqysVKY9L3TkDwV
EkdzZnMUWWkXpk4X250mrM5zAZdZ0lKAmeIKDFLXioqHtao4RITLXsmg2LYQ/+Va
WC3m+N0DfmZtCl2DrbaKmhV8NqNIrVQFZcL9/NivkszOhaC2KIS1lhSn8YcGjvzi
ZcRGuODgKt4/FwYHXznz3wDO9Zkj0WqDbYhBBBxeWOnO+a1kx4nym6YIGKq5m0Oy
cZEiSIMiNHkaGqXXaD6YkDvPTRKKq82uSeeMYm9uNsUxjUS4XsfupPaUJ0lAH2ea
nar+mSvQEi9F62OmXaEfbzaVRhzAy8XrwT7oN4+gtKVftO5AotLcjClZz+EW6xCO
JFI6mWJnle/IDIHnXnTTBl8AG6u8OFX0GAmz+3QCFwZXAc7F2OGK5k/+ldQgD4C1
YIuS4kJ34M2tMKyMppWjRzBqMBJa94R4xeY7aOkStPIBK53PAnDyD7SpDg79D7iI
pAcQR4/L+FS0wo1aUN5J99W1NU+hK0Fa0pp43QjNelS2BHB03Xp8Ene25vxqLEbc
WYvy6ELUw9mqM++H84I1ck6IJfiUU2u9Xty/wktAgpijsQP+DPmPombh1XAbszBr
OWuD7iqYZLZ2j+bPHKo1ndUsLAZoWHHPyqrha6KXfqnWeHOVz2OxVTaOJGhxpzrl
oIS8axHL0zFl90Q2ogdIAahLLzCs7UKFgdvoMlJo0U2RLh80SvJTwXUPlrAmFFKF
VdHC6LLJH+lPTGz8My295K78T6NFPZ2Zcy6Cb/KFmhMdApZM96WzNgs6ZBhgmS//
LiwaytQGdQiatW0SE7gPRdpJql4M3wv8FoXkrzyCNZZmBnR703pBAupw4zq5zpC8
VVWn/xI5a+rDlWxX7LIIyUU7ViubxQsUFv2kombLx3s4Q6SvlBCfPXcrIarN8nC4
Fz61rIyiJ+DD6oQQ4uFFeA875hjHDBPMFJUQ2kQ8OxmFdLoQj/93lK6ztydTZcBm
AJdnKThD+s0BGdwWYUFdooPzre4l0/WULYsR1V2bjp7tHulq6V0zWG+bSkxYad0g
AfT1k1uGyeSLtZ9briLW6mTqAkb/ayaMvOhSoAXjG2Jfsz2fc+gbUXZBDy66i6OF
+aQphAGcnqiAk3xiNVh90zKWzrfF3+AFNFrtZF6RDh2pT63+qAO9s6iz3wZs+1Ma
iSVhCDDcwUaU0svvGQBEyDT68WnGrDVwqDFRadVFijsQvWhHKlEDoU7zZdzBh8G4
v+ifcb/U/azRvmGl93xXBN4F7TDO49WF9xSHV9HlaTmXejTWLS3TdUfipc3N1dl2
IdU1wvLAm+mWYurze+gNm6n9EzMZLKx0gIEHB7dgSfjKiGPcXlFQxHU/Id+qx6lV
1TP/hdIyZAL2tbNvOlWBeUuhLkxL8ziy9IniG60/KhN+vH6a1+HiuAyngWqeh+7x
Gxur8WdRUYliL0bakaFHsgyjqruh0nCLh79vrlaHdTKQlJfsR++ft6KZOX/7YJNj
N4F79h18gq0+EDwN7ZWruMEPKCrkLb0Jx+UFFMdQoJB9hGpkBbGrOBM9X47YBV17
rCcc8dTfjLiD4mn3LjcvLJTm8i4ADMGo4yi3I2aROTlUSntoWfnNIhutljiDAvlH
BtbYqipeNN4PO1re/3Ow1Sjiq65rXHj9dDnB3g52XkpOjVpNonLs1CxmzREo18sS
qLEP37+pZ0J31n07/MMebLiHA0yVSUcOchz6ArW7rA1TJSpxs7PEsD+l6stF4AIa
UCgYk3cv11ud3knttZiJ44nUfdByUSnHPGZ3vsxV6RalDQm1AA3zl4nqfnvsqW9y
vNC73oZEcuIjwplRzN4ROOKzgJAtmcDcQCKNRAqM8el0vmVwaR6KYKbIYq7sp+MW
agNCLtyh/xGjrCjbmAXOLZ0dfESo12OELtSJaXFMA/InHJYoIoem4qK8kGYPelqf
bINHA1r0LCvjRbJO/EW1dnwf3syP3Ef1xSoWUKKvlP8tKm5qrkmm17AiXlOOTZTu
YFuJt7MTDzaWRYITyK/DTUyfHv6q0ROxRQC9Dc35XetkEYNbk9PxPp4yIkAE/QGi
TrXOAweBlAAecSuap4WPbfsAj3KZBJ0E9IZ65X8KFHCI0H9Vh+wJFF4xUakJ7OhZ
PXUvllHIjXFLbHV0lWhPf4n+wamK0w9b4CYqFEokQ7jUeW8V7HJJnz5ebr4n1FA3
ku09FHrcHElwzCfTb+Clj5yjpBAAc0rSM/kiQxMzu3ILDqUykdEhoXlDgCoxa2fO
OfOfd1rAutsGdizQkAEaDXiDZbLKUF12majP+tx6cyzFHHDZqaiBY/pbAsAJpFiB
ggpV4yOyfHCpGPL/Yj4m/bVdroT49YCnHDuYSaffKUtMIIXvTatUBxcD63tV30J1
B5qDEPEzExI1tSnjqvDxZ+EzJhRkIbbHnkzbdEuuQcYzAFH72tSV6ArDVxgPP7UP
N2cf86bUica3TP6qFmkLJ61KY+CKT3QlyWVaLvYuKtRCKXbWCcy0xUYcPNfB+QbB
so+KQKMFVbyKnHHJ/NhkpwSevu45cAdq95IAesd6q0mZQaJf/1ApAVMnGuF5WOLJ
xGqZSRT5f5tyfgAot9uiP1oSyM053KBSvogZByaQs6U6RhslVaLuBAGvqu4gL80Q
ImKhc/tlSsHl6Iqo0W65mu7Ss13uf1VNgTb6jXZVggIfsx47ej1flN6T0V8aUr88
WQ7mCBXmpI5+nNty9mR80r3LsECibK3YANztRExHV7tA4I4Q0vLZBtUtUyctA2Fw
yXyP4MBZZd7N7zg7kCwKffjYMrmyDFh7T6PbbWPNtRXLcoIcYJy/n7Uv+5PLQODD
5grOTtEjKxqlzsAjttLywd2hwjIosFrG32HuqxgnDvm1wsbvJxfDUG8wrgZu9GBJ
3PZ4lDm0IhKa4XUuuX7gEOKfgPYIniEnZVnfltr0u7i6j0B4YOBDmqFhT8U1/05g
yFlcjLUN/85eEmU06oWQ1XNloRwimEaT8BwB8OizR29eJY2Mit0ueK5t4NrTAkto
CBzBOnMcFfDCHWwDWb3jhwJxoV+wvibilsS3eu1OKD7BPDBm1s2YuqNmzpMPDUQ1
MfhIwU+5Ndies3EH9o6HMEn1qJvTkE8JySAiCRd7H1Afasz74+wtV+2FHOYAVKWg
ZADJT8tqE7WZI1szCRAE+t33vUvbrCGaaLhk61KWJBZa/h6BpTBo8uYu9n6/zonH
i0eAzQQ/a+JZ5R/n3LrlZ2DJM3IaNpXiXQWzXP9n2SRneMsCGL7MHCgDHO7IvIKB
2ibUoUX39f+e9+XB+xX0GxUNUJNzrHRZ3bImbIWEdIEzWOVDbKNAiAxakysnRZch
mhl+l+lGrbEKDHmNriaD7hUaTZhfnXa9fWo0vPeMoc/58KfoEt22+PgTobvBNCwP
N55j0KB7n9GJqZ5osMuDSopMDORBmTb1D+UM9cjOMYYsweC/6N27Y4C6tthgN4uF
SUpR6wCYsudMPpywW8MChyq3QVxDmJ8KC8x4OdMelmEBYoJHm03teK85kH4zWQ9f
gW33yS1tS0styx46NTWGUP986PwV3pC2EcM4/Xfjy9uBsBuXqAX6m/tTugOzJoAS
l/Q43xyOORPHeddyw6KAkAC0YPmU+odKZF35q4HqoP2aYzBfCsQjPcb2X0d7TkW5
liu/oS4wu9EayaM5D0w6eusjeB+MjazFfoYJ78uiFDUoo5BVcSo8j6QCF9KueTn1
Zi+JtIpRRgsC5aLqF4ntbOYJy0tdFGW+Z5y2QpNyvW4Ua/zuQhpX+Ox82NJz+k0j
5Av0fDT4lZerVv/gUvj/pzrfGqfrAn3Arp7lNuYkDTr3xAByPgV6wWtTq+NsmWSS
V6dHp1/tLNd+GMclckgLsmX53UuE20/cZujGDvrIkoeQAXFXeGgcAGis6AzUM657
qhEe+glmNWu9L/WKNohmP6eW+NvkDelr/dspex/OIfc3eXwxvwK3RbvhHLlja6wx
BF28fm2blBHJUyNkPSL+YqfFeS1jlt3sJ1EYfGveIDOlgvXahZVUAsVCmfR51Xdf
eYHy0y9c0MZkFp5O568YX33S7jyv/KaSTfGaCUgm95sFuj6poyJjHweBuky+KzBv
TcWgXFOc5QXL9nmr5NHDH11OQtSyPsuchYZf0pdIxUXayWPyEdL13ZOs1bLigItd
m8TrFBMu2WfrE/fLSodnXHQylyjVMg3VTCQ13AF2Y456FUr4zPf/X5eKpQ1iJpYI
ENB2TFg/jHquYcHpM6AlrZIP39b+9saIAUFdNTWFmmT95Mj/yHZKvVxOYiYqprTM
yPr5UaP0QBKJlws1snhjWPMAl5F2TIHApWfsvg0nnye3khJeAf6TQH595360mp2o
WXhkShoZLOP/f9KvP1yWvJsd5XiZOu4CjkcSElZJNWL8x/u5iA7ww9zOJPcsdnQA
eAgkQrpuR6O+8pCFf9VzoAhjxbheXrcdv6UEy9XyvCeuewXAdCOnB/ajXSyxRTEZ
41iIk4HZeEVO+E8DVWH+YwUcYKOR0VcUwzx1FXx8Hglw7PP14ZpR42tI+fSvW7OU
aWZB2w4CN61VdjsGlfwqpUyXRrj9Coa7zvYJOQ1kfju2Y+JMAaxsICjecyLbONXE
JNcsOxHpW69dJDUDHPUl8lvtMrXU9ZsHcYQ5ckPdHd2IueiVE8D+ChqiTCb+qCri
re9bAr+ZdgaDmZfRbOmhl6mWg85UxvcRW9V01ZNFr0nwREX0gR0+upcSi9d1xnor
k3qlLw1t38vw7u8p6umvGBN2ZNdytBmx/LDfHJjSSzf3Z1CB7kTzX/Wz/3SH357v
7dVnlj7zwIbabOTT2jG91gwnBvi5RRRyL0KXvDjafF6S3QzBE46WHTEW+85Gyhhw
KzelZKc57mhVFknLOqe+7uuasFuuqeC2FsTd2hWnqyjMizEiL97JJkjAr0AtPmo2
olR+GLRTdaUaJ36NJZjrIhnZzHeTKr1+qBYbZevRalMAOcByx3dWMKcbrzpdL6vH
ojvIDdkxDgX2sbpQfkaV/vStJSBsAbUuu0KCxyps7uAGTMZ/mIoQLhAIsyf/Uc5W
MQ5Xk7Q5J7jQzTlsg+yzxV9AvJ9ecPn3pFBeDfce46nHg4U8ff118qMuMyMd4rbV
PQhLfn2HmdtXAF7EqNbP8QGJ+78sFDjIlUPmEAzE3/LgBNoEILQFJ4j5KpaferFv
9s8It2FySDXeEXmdBng8L88eF1u6TuMpxaUHb4yE7/psjK2VeZuHhIoeMxWHmvtH
XtCG4vklC1ifBCdusurBmmNLxZcJJTmnI6sS8ynYdvtpNcdZGNkzXZUzHzQRrVTr
6gdgTnwUTD7HmwoN8CjSTlKiKUnRSWRLE28Vcdx406x16hyHbOwItaWXXo9tpkVP
7RIlQvSPSEd0iaaSHA1Vta6qmwfkeDuVorTukl2A+9oBD8dMWsKgjf8HebNi8mYr
DFeJyBPT6wAgeZ7iP41odZyzRxiPKQXQFMJicRAlFZZmkVthLfDJCtadjPQ35J4n
1XVknWliuO60d/dlukOuGOPnClR2GF/sScNSNgaRVyYZM47/D8dA9osa0mKTLKZI
Vc9uS0+UF4rXTdIrw2gARkRZz4aCarQ1l3phKjaONqv+FcIjpjlq6CMq/VAfynu9
rBZrJTome3mLc5bXIxTiH4YOb27okh4t5Q3ikGOt2hql8jA9f4xeIJdbMzGQQJnw
AmC2dvZjak/KykC75pzC9V3C9cKmAPIfC0UfaXer1AWU3Dqtw6XOMwajdgzxIwHa
GR68soPwLe+McrGCX2MTc/VcdIYb9nLugZJT6xRAXozNJSGj9p6Lv5zkYh8tRC/R
e9FH54GiQk6zt2vQEVUADTf0BCq2GvaVquaFFr8l/KvvZ+M/GcJyIoTUovja/kSH
ykO3c9cVq+wmzl6dYVYvYrz+3H/uyDTwY/O5CwK0DDUomyAf2VsORKuV40u9x/eJ
zTFmSNtbbaTaGQ+IQ32RHBrQUe0zggmHB+Ynen8VJQkmTBZibwGhgVN7m5L6blBu
QF2+0/cx4rMgfSxLMySRIM31xDZ/lu4t9JDzOUVLzFzereCczPKgLVnyoFS/2uJE
H5QH6EvfgnKZxwsfSWm5VwJzLwAyk7X9b7sFVjRYUjv46ho4H2Nojjrp1ffVrffB
5Uh1kjSGg3CMkdGwcBKkG+a9W/OClet6DpJPRpiseBTsEkb/D1P0aYUWKElxYR0u
rZFAuAcJ4mecfjc9s2+I3UstIK6SbAaU9ksUjueX+NiTfKHJbKzecXejClLV7glr
QdKw5ZSqDI+vZ6lYxGf+kzGywAMLokYJ65gTg7leZiEpALL/EIi7K574Z+MhRrXa
qCBsqVpDp7iSueDK0QCMrKVjwAZGybAd4RYC1OYrMUCBlrK2lpW33JWqx8om3ijz
IfxHYSDdtnXqgYjbIiUCfg4UYEMh9Se8gxa8mBdjmy9jFiaoELThuH3ONID1ybSJ
6w3bV03qFSwgyKQV+WE/scBbKJL/E7voz85MeKuTj28MNQPx8I6TSx+ZsxcRzyDF
mDZ1ItZTUAOJbObf+MSH4w+tr6dt1a3RJ6cifi45LwRFPIOZ4pHj3cqUEfMAWTum
by/nS4rVSM9j1G2P/J9WbmLYo+nKhCN75mEbMZT5oCpj/DWCWKmeo1GQqk68fpmq
pGLnIfLTkQ2h0gKkHwOLIIltTVjBIt0Csfs1H5Blm6KJQX7wMPyeG9tR0ZHl3Lzr
lQie5NgbZbfis1eKYoD2GY+DqpjuYhBqtooV5h7Ypyo2rOztQ2IV6nHObfqMiu4p
ZNm9T5f4NjOnnXcjV6PTPUXkKdLy8XdyofnQPZggJX0kyh5rWz9fzKzjKQm+YtI+
TTmxaQNhi+gNNygd4Za1xfergBvky6Wlf9UOarrBzYiKMYLJ1ZQUWTMMThwAsO0C
BISBo/PPIUvweahm4wk+XQdu3qVCOVG7wuvFf7FjUpJK0Mf4+dzOxxTMOO29T0Mp
mu6iAn3Tp6qtiZMCjpd0q5Iku3zTaBECyxujvxFa5O9tV9AZiuG8/I9nlA9Whs3q
QSJpr1Lb5b2qrgtyJcSbXlc5ZVnuMX7femaF2pMQHhvPBMGPCRYeSDci+zo6ZfbH
5r9ebAs9AIznj63N5P10KgB9K25pe1NOm63IPI/no148iMc00x0Ef48DTiBo0bzv
f4mIqkR+NcigZUawUyWbP0q9MMMMpg+ypBasRpaUHW/lauEquwFhC4Pms5WPYQ0v
WMlRGA0/UyQzYWsMq/zdzdKzviuz48I8cf9A8vBIdIhQn1p8O+aRngqVl/40IfxH
egQHen61m+Uq1ayli677lRqc9Vi3anmg74g5AW7EYwoXaP1LAzqLFHD9UVMcIYfO
goVcjrAAyiZSWutUaiG9ntibWuLuc9SRj71s76k8b8nVObZivt3KgF4uGOd73IeY
esp1KWh8WoCsIZyAHhlZzwSyu7RBO6CN0+FCWXV4npb8oL8pA8uKkMkwobdTZSDh
5BApN+7cez9Xg8IdSQN2Yu+97+ukZNAbrVkafLxB8w7v/3czgNonvkpStnYsFHRM
pF7qgRuc3j31yM8elDiUkvU0q0nBhn8HFNq/urjpQYELOWKVd5hYXw8UNFRbXQ3x
lFNsUV9Spm4woXjnuFUZ+vu00zOAnwIOqdanjyxvBUWTLcarEtdSPgOBUlVCOUqn
baN0Q6seBeR7A+U/2Ajj+Tx/qxxoEdW8zIkJd6j3HE1Q9BlazvNo8GI9EqKa9cOC
MMK7DqzDKWXqg3a/SNudgAvjlBVSzUFP6E58mE0lnJ77Qb59nbYzKE1CrrJVeBbu
acDrXpUQJM/LT4AYrRYUcfsXIdqKzg1jlMbFrYpq2+X2BYs21niQlgW0zz6z8hUl
aH4VpNmEIS+pIX6rJ26nF9nQY738vLao5RzUhS2Itu3WK+4PJgc+8LT/jiD5vQQv
0FL43uMTMKsihvNrYLKV0BMrjaMW0H+QeR9GV6JSFtyaztCWp6JCYarcfO7/iWyk
Brynz0mZn+q3OS5m3I1bwkJyu7qpNTje2mOB6ZpWqj+Q0DeCTQ6VIstG7m7GBvce
sNFbqH5Pk9k4fwnDPPr+P6Sxe0uo5LqeJ04j+sJPQwGxpAuzlEyjmsxqK3pCE6gr
UtzXvYR0xDzEc0RW4hipKj+h/3rahcPNjIZorv3iy3+Jhk/PU97dsgZ6shq0UUEe
9pV4K6LTbpGr4AORRUHHUNky+uwM2cOPuKn5JaKJhd4+Fvqp1NOugunyekqjis69
bHVPdrZ2jP2/MbuBjKZnPv3IIaf1eNSxqKGvaSCQe7krHqtBWzRgez20D5X3+BGN
1w0nqq/oO55D1aVSHrJLvor2FWAw1zRLQAAYMq6QcS0rXTg0NKu8Ltdr2jC+ZHyR
i1kCCHkG38PMaF5Bva8dGMwlqIj2qU0RavYSMtCowLfmof6CwVg3VK+NU1E5kHOt
Zt0TBA0Qwihj+2QW2z0fAHX0WD6oYhwheMVaNos+jWKrGrPBnijD0rV08uKYPpbc
UuGo67IRi2qS4EOSasY3XXF/h0FmYishNwq6IyUgdgCKPMZsHSwoqavmOW3auiNM
IXxCZwlEl+ZasP+HA7wup+0tJd7paL4uCZKJz1kS5/WJ7eBXPFWQeI5cvhZyR4dy
jf9ZymhZ26EQcO9giygGXw1TLxnQcxbH4Dsm7yfKPlDWrbHyabM3vRxP6T6vTPxQ
io8RUZ523e11W36tM7jKd/+M9Cq8EkqHc5VMGzuFxxYGpDx3dzDekQufFkOi61+D
bBTma709i/C8j6JM14jwB2WtZU3MA5uTZ5P8dOlyawjao7WBSqGaRAk+TUx/WajR
R7pQiNIe3QCX+NDdKSo0wLrNyljVDGFu88EIyR5A7PNekcPY9vofVtr+LucPHNZF
EAMT3pKNW7OGTqPQ1ziF/1Unyu0qMs/ZUoN+gnWOKkjPoQEGrA0X8CE19FhYpF04
eGI5fuUkAJZLyGFVRY54L5JAedV8Vu+5kEZ3S7ozcoCIEZxgb/cfI6c0O+Jo1Shf
Jd5L1jehCSLzQCRNaXtZB/Dv1IsMDzd1fR/7SHFEa4e7+CHmhVdpIwnPean8vNsz
sX2Fycq9/2J3r0SsaKx2c9h+GgHsN+CnKJVMz6Gl7Dl4qIivL5dvresk7AZ2ghaH
/akmHP+/Z/xwLyjv7tqBJ0kZ1DUFTQ9C2gTnvuyZhslj4Zg8LxvXqrvHyusBADKT
ie0fGtTBTKfF6+Y7GwFa3lnyxzMoqcagyvFMZUigNUiZrDWMl4+9b8C6tV4HnUiY
vAE/PS7o2aT+gLaFAKWulTxppouqQ7SCcncijeoxkKuP9ltbWbRcpQ9ou09oX7ao
qJnW6Ko53VHsUqOU6obE3YwuE/qrIPbfU1sYd2WcVbphy858WHcxq/cGQAy6Uu8e
qc4zEz0XZCUaDCHOCTnS4k6giv8PmnqoZ0KdAUup0RXcKuoZj1Z6KjivzcrfNGZG
hnx2T/U/WHBRQdFd0mDKejOa8zG4tVhdLJEcJoEYbR52ZVAL+kJXOlZYTzf9VyVF
itA0idzrYIYEJlseGTHTa8Rmma0IEEqP4+CHS/EC20OSZwZyUObCc9rqt9EMDGmg
rJu2xmOhIrpT35Q9rWIbRpiihl3sEa1OwPdydu3J/EZm9w/Bs1XraH9gvpgh2o1z
t9+FThIX31S86AfPOWhWWLAEWXn/iZa9qnOlP5ritlmm5stLd2JXY29WWQcPSNYl
deV1CH5+G/1fVOrfnxxZtWTofbeq7EuHKt66Fs5M3N4xTpMX40bxOGE0t9eStjXT
WSp00FsFG3EZ5Ei9chKHqha5NqV2jr2aKM3JpEQ+TXWD8lae+j1b2W4Aj+2AmrAi
CdsiHv5v2ob29EBfZaFF36im3Ni3S88kKlbGNgjxA3TZ+6RFM4OWG1IfKL0Er4fg
oRTjY/7Wd4FsmE7Im9Y7FDAO95jF1pDhwmifhOoipWlhlOldV0tMvQhWWRIOHzRd
bUiuxC2rY9QaCSL7SH4SNhItZzn8sMjg0ZQOX3tmfY8IrAgWGPvE9vv7d4ja0ep1
cbLrF542pj6XqiHg5r+ckn9MolavtBDFiNRQCl0dYbmOwyBt2EcXLmW/E1qIEuIe
VqYlfc1fLeojpQMLL0/1vfU2cq9JDwE+goe3mEpnFWnNMZq3rom1yN7RyarFhfus
m31vNuPP+NSXWt70iV0fnFfs3CGeDRkCSqw0xj0lAjA0R1mOWRys/3VjuFBFWqrO
bzvefqwpJ+QLCkw1g/I0tTAwsaion/SNiQqKqqcfuon/+COVQO6HMI7Uq7e4isks
x95MNWxGPQCjKQ890DjLQYpRynmGUZ/5yBjlzCn+n8LCOMT/Owbu5NbyTnZL8uPF
J/7P8VdpQllIgigYedVeguVt/kjwYFWToKcw3U5ue/4wozBFXMSK8QMo/QlJDnoU
8GgKuNPD+glCCzf7HBNo6Ms9MhH6m05evuBhBywmb5zLQx81sopma1/YBAoSsL9W
oEjVwvQBXqp686+q/POFyyCDW9ySOvuekTco/ztpExA/C1/9Dn5d7UBrA20M7H7u
WZ7Vx7UUpTXPx/bp8wLHZ4QOyRCJ3W8370+hxAQto2noJWlifyObKAUFPtFgcUAf
8kAyMllJ/N9/Js1AwnQmiBVGDsf3k+1K5FP1QV0c04cEK0DkTn7iQa14oevo398s
KbEBiuhD8GWupxKqvg9tirGGzYtdMAYWcG9TZyHkliBx/jmh/hVJSVc9ArZnBLmU
c8mb6lTJWH2tCWjc1hJHlGk5KIygxNSNBXFmWM3eI7phKaM1T2B6odwMxqieP/X1
VTDPtOXmsP3FeFDdQ4VpLvPkvfGbaVfI21M19DWD/7EGwhilBfsNAcZrykJVF1I7
c26uOId8jlzwrRBmGYjbhxixieFu5QjjSiXVG83ArkVnF+W145Sj46DkiJKsnT7h
X46PzCdMjGKd9gPDIzBCcSNcg0swxEzZTGjuYlVw2TUqR8/fYvJm1sYqq+epWVV3
ievYbARB1zjYRD7rC99tTiFqkkg1ElopTbXzLutHMl+se1sSecdQZwoNBIwPuyjM
zPcuxIjEugtMepa9BSQyLLsE0Gl3e5o6neemeHFoDNauID6G17REWJsZNSydDfuE
ApNfbYYT/R/71RrHv6k9Db3T+W+4g02j+cyTOcEWJO194HLFwkxR8Be/zTGYt09t
08mNb81aVL8Bfl+2SzWyuDgjayqA6I98Qrrjr7fApAVt9TW5BYjqf50lIiAmcBoP
OLchMU1vVubQaXizSW5VhC0/pusxaxDeuQeCTNXY4wGMQD3bH8g72Fzmnl//memd
7NKobuzj1NoAkeySlcEVR6ox/nXeKLYhZdP4oKyjrqU5avc7SXEEdgMYPnIy59KG
dOeH6nuBf7GCgvtgeYYTk0/B0NTU3DB/xOLpJOyhtx8roM5YWYM+DEDxswcfwHP2
VSdsqxKkpkh2V/qyVfOrB8ywsN80M0GdOwAO3fDlsTWPqMqnZPd9R/pHx4j+Qla4
RgJclSU1u4L9RKvPSCJrxGdd+fedbuSV8pOiGn6LiCKz733bAq7ZpYgc5m5f73KS
ubFESQOVSuvaIwdbbhbczR2NeF9I9JjtC9yd32EvjJXjsVbdVXs0iGm/FFavpLpl
yYjIcIkyernr9Y0Fe2l3DY3wt3k8gd35jutYycCeD9dILNXfjWbQ+0uayhs1DX1D
1dtVY0ZMVSwxyCmd7sFQVtFsitWYOSp8BWYS7NL2lzx1g0ZXweY4E+xOecbyhNx2
y9+jBRP9cOl84WXPJhxTvlyJHCcMjLmt7zniBiIwjtmGEGn5jh5AaGiEpd5uWVfS
o6COrwKwldpx3vvDT4t8EL9I0CHzEjqhljIo6h+QWWclYGEfs/dyJWD0dXnda69o
byPKmcWmpQySOD+Mxd5voSbM/V0jPDx1TdIPGe2MIB/TfvBVHIZ4inFDWQNrOn/Z
Epfn5V/GBO1/B1mUszh21+DG/RsFpAYyQlpz5fVroMD/nkKVEvwWVPjfJdCjf58D
JqhwlsYo0tDw/njgFRBeLS58vg4dQaMqr/eZ1sz5wpFEOIa0SSdSaLg+dUqtGwjm
DMLAgkrOOn1SNgXxVd1m2EPLoV2OvLLG1akVXmwDttSJ+AgbTNhVjhfVqm7qNsgq
I/SCNI5rTjNqzsPscGxqUrei5OdDyfqZmTpa1VM4PobKV0mZK1btQzH6E6VprH24
6tpriyhPOIjBA2FyDtFdn2VqaPDl9hHwVO7sht9CBpEWYaaKxpmWLXWq8xDHeNd2
tb2LfxiiULwzr13FK5vBqh6DL3qyIGPApQMZyiKag+phQR2DWwqFg1dwMZnIuu6s
/SBAnw2zQy+xyNt1SJj8IoWWHtRQHqfiOpARU4eQp6PWlVk1oDb9B0kzEwFYSqLS
6vMw72bAE+GmuhDoiC2WempPoORYSfkD+k6PR718T/3suDF9t9c9ofwLcCrpWDp6
kouYOKwPmVjuO+H0NL64A04WpYWocErB0PtTbxlUcXsnMG1/9xjwgwHMV+h68kHY
rVANoWBQa3oR7CcMt5RHNcNRLv1thLIjMv5ic1cz6RL639tgW4OVz1fDt34GDrRi
sKvdnwjSqeOy7l6SB1/do2ISmrcp2sLNTLkApFi/u7alAESfkfBPVqmbfdIZf/qd
a3uXTzZi7eK4orE9W716q67x0xkcoZ/wNHD7sK7Mvk5CjsRP8qO8pZ2rbD18ZwMt
3wsgDXWvNv0BHZ42vKaFEudmOfOFuTIFRXfUjb8/FCIFmaBgopfaJhuhQDHYoNYa
SwJNnsp9MjEoWS0c26w/BEmIBlU8WbCeXU4GCb+4ehNBp524Qov383xcfQPERwoF
QdcJrJ5LICK5PfPWzLNdjVsV0d7k7Z+lMnZqaoCP5ZMmLHOAghyrTYNfEDqDVqxz
PkBR0zFm1EtyRlsvIFKQFYi5jgv1z/xHAhpytxAH46wo0TGZmoo3S8wHTJL2rBRU
+f6VuFtFZEEurmRVAIiK6mG/yXh9Ns8PR+YIMWX+D9utTCfjNV8cag167V3B+hcS
E7EkQELW6HQTtQg4fmdVNHXF4/o4JJHRDhkbsufyIZ7lJtmwrltlHE1X4TmIruEZ
2VyGNkE3QsSdgRZ3GxgxDzK4JkMGpHvPY6irZbYOLLckMnfkTDb0kag0ZRYJMQ9d
VD1DCv/ZES3/1bot2PqNYQHEWNWCg81992ecAT7Os6+ubA8XmFuCMTtccQd0iGCp
ohJwJXU8aUp9oxNyaAGs0GcQeRF4YT3NFJJDRlaNuDMy5RJwInohKHe0hiCvJSvz
o9KZo+TgsCdABlxEyb7hSyOMsxANjbFJRMEZuyR2n08AUvmTJRUR9SxaYpNfMw0v
jBP+fvo8aj+CXY4r34ZtBSqEl9tNBdlo0F1yvYbSWKZ8NXH2KNSSxx18B9K/ubSD
n2GuQpAesK1aB5DV6G1FZK4t6wfrYptd3J/1RN4jlePOcA9W5iUbToMTSdpVJvaK
mFGH793lFveYtBiREuJ0QMz8yBJEOzSwqxGzfyGAqGz5X26ylXQKTlcTENPF1ZEV
itFDQxZDSHN8KbxkIrz3rc3p4TOBhEhiyFHDeoDRsr4kgynkdYpq5x/Pl+Z/xM4k
o8NSffu0TY6YymTboxFoCrlG+UzBKJev/4ul0WoKQ6BAkcpwxQ2j0XuKhobdOxIa
kml4/QSyu6Pgw/0Sy1Pw2m3gTON1i4f4HMCeLH628LQ2qk+/N3s9QuOR8VIunM27
vLo3qKfqLsCTzTxlsAhxnBFYzilWs7xS9YvGxo1slmhlzTp6QF+XTbwb0A/5O/Qg
Icw1kFA8Sp7vkbrhyrFdFDh/H7WHylrY8cG0jwLpS711w6MKseX/fiZ2f5C37RCI
qTcEoqXG71/1u76+aABNrrhQje4eUIsmSXuWU3tE+Rh9H1YaK2uitX/LlpLCgBjo
nTQlV2Fw9Sb8v8uDZx/kq7HoPzL4JUrN9E25JUIFcYMdocHkjKfl0uYRXu4n6st4
hmnPZHQwSZrNjsDTCbwu6ducgssNV3nN6oYDA1AYyioNoeIM+WexphwAqIM7725k
kjYpD+cFE46+WW9s0ZJr9wAA6P1xnB7fjzVVlvjQa2d/7XDy/MvELO711RIgsSZ/
1Y+loHfLbXrWnLnLBqPj4jL3KPhunsXB3uzYIqdL0aQcIYvZWiA4DPXOS2Fmgf4Q
3Ul3XBGwEK3RpUvEk9c+x5llrNrVzSMC1v2H+30ipjVgX55iuAPkeQZKHe33BBFj
XAaysk3OAbGYx1bum4bz8u6djj5HS/FuJ0a52oVlJ/dvJAt9G4C75UtFFbfbqSq9
jhbnmoW7gu+Di83YHHIvUSOkNl1SU/s9enzNLw6o6W+Wfz0OCy0sOGkstNylrXLm
1O/SKaBYkcm5ttC43wpdcWDEedDh4m7zLwDmbwRCWFJatkgM5VU1u9lTr0oS+WGd
c931UUAhQVr47kbqas+2a5PzieIMlDdifAVhvDxWtqVq/Yblp7Z0oX+SO15uj1v8
YE5sa7xEnepNdGcFEZYAOJAJVGxx3CN9cHdLKBO+Vi4iwuwT5NgGNdzm54PF2YzQ
VGP82QilQBDbE6rR06UZO/XHZk4xKzv4hxnR0a3Gggbd9929xv9ntJRpsRPZdLYZ
6E9K8DyIf77BV/2ez9E7586PCvlgiF6PBxevWzhhRb1psS0O4vmZ0wwEyNYdKuH3
S0JPm3WnODzjGZ1zWg5C7PdW6aond+oEXzJ5ZwjwrwA6FX+c+jA4q3sLCjGlgH3Y
Ff2HQtStWPnAspyluEM3o5SjvBuO9xj81z4HiR3hPLQvr31/qHxWOLXF5r4lV7Hp
2efWiQTWIre9jxGMeWCuoMj4roFSgKAxyoYEw72NyNwN8zXfYwQAduBMNv51By1U
LoAr3ytCi6n2fzrVjkTUzpPQnZrgUCG0DaGl8YHJ7oc3FPam01o98XUNJk8SN3kX
DQT/0or3AgaWGFxshH8imzA79cOAdKOAUciQzqS4k0gM09LOc50l43FW4k4EADX+
i5XJIQeG1rn5qLdRfuYOpkTS3Lv3cQjWk1QYdEo5IzSNx6uEOszspdhXvYKlx5lt
GGY0ZwiTeFoJwiJwiol3ctSTdBIpQERG1ovBcz8qOtp/RPoL3L1gli9x1AZAq06w
uag/uNJEF7zAVdrlb3vh5lMvyn8KDrUPT47siQ/6ts9Y3svrF4AotVCgZ7ftVFi0
lhvyJHcjvTe+899kBmV5ppXYh2CIeXilc+wAS779u+VZ1du+JhaiFT9es4QFeEuv
Dnj31TKPeqUQ1v8Cf6PrA3uqPYvCWyCgCngY7wxRMRTqqC5O5bBGBEyLQVKaSs+T
IsGOLMOxdR+xwrBYrKnOuJcXMlyKlKJ6+0F/TfDQ1OPgOwp9Plr0aMoVgi3pA4/P
Z4XfW902utJvvGfEPmZlqDPTC1liz17wS6q3+x8TWsuFElAcdFe5HwmFlWdOtTIr
Rk5kAuRCFzXgCua++oRHzIHVZUrmPJWikux9Tj9V+mtDvcc2dAKGiA4DGhic+uUD
eokcfxX9doV8Zu0RxLm/h4PhKCaEfBZabLcaMeYrHaT4dqW1+RyjMHNIkTbaEltB
Hz3/gX+9OiTC5Y3dqhX/jNl/xQumxKqV3XnXdRI5I6/rh5XwXMjs0PKZ6sKKe2dm
9VNoskiQsm/nOSsCj+jFfyLNrWfhg+WowylUTs654jG17/LBcmlm/KZg5EyHTUc7
g55+p/d2CDVfh9BoTF0mQidcN0192cnv1gY1zAotN6dArDLZ6EyQFG8EyVFuuehU
aJ/JRp9uE35f5k/wubRszCT1CIQTRBKMXhfz9guPkvDbRIFbAQYCpHxg/W2Wzx2S
Y3BJ4jz2qjyPBbRDJbGMXAZTlhky8w6cqFDzh98PtEUs3c767pPwfbJjHgeOjb/Y
ZEI0qAvSD36jOdsrj5rqozjmOhjQIAyZDTkz4RQEa+19sCVxaxy4ixy4rfKmGjnB
d0sI/4R7BfuMC2eOKFltpobrzOsxZsBCggM4gpum99kM6xQPprXMbaNBTAzQm/w8
zfs0Pc9gOd43ENH8ML/XXo6oR8UgvUz96mLeemJfrSdC4N+fYit+BGhzkVbXSsSn
G63Laqj1jzjUU5qjgsbY0q47gIvDtRanAEzHYVTQ1798zNzrUqp0vwMZz0Rlr4x0
nlYwlV42jwsMo2msEJieKAVvlcOBk5ZvtIn0aT4md5ObsHA/Pqk0m0qR2ACpGGVf
7DOTXud6Np9akwIGzgiCI25D3j4Yd/c6GogpNga5uagQnT4d49t2bSIPJiUuOdYM
wWs4qmiDAOumnfTfWgBGaLQr0G93e1Bc28hf5J+I5xl9HDldeT8/bcFMyUKxP5O9
BVz8b6y0XIGq+MWLS7km/qoUiV7cBe8NIxb6afrR6aLeR56FOKo+bpWLw0ACrthR
avwyZH6Wq7AWUimCmNgO/YKh82Z7PH5bKwiWSiH+sTiy1CkILc+G1QWkIMmXislz
WUH7E6Lg7P1QhXEk4QLo9PuTjFCYRfoJazHPAngmJJBJL82WRT/6F41su5mw48Vp
BYb+5iQ7vAnpR+h1Q+WpYKnYDl33ETt7MQrCz9my22RTt6gA/RjFvLXCT0Nvces2
z+uk7muoakcumsEGtNhaKgM2IUAK28e/kU/hvji/eBsKDKL9T3YnBTtMSCpGrSvY
tQmEnaOOrsejoKo206rp3en3odXXlhgy2yqY7v25D92+lknz8pbfMlgKVv40hHSv
Gt9hZ5EW6pB52fO25V9VHnem0XcGmID4+iRbqHE85LshdTDrTc3zoiQvWmu80tL+
yJCzeIDUX3FL7h6/E1VZqoEadKPBNZYqNVGD9AFNHc73BIbAVKCdiU0J+8owWj6i
XxD91fHSBSZw4DEFyPE195Vg8/2Xoz7SLHGk7n7EFZjWdj/MwKXvhBAnCEc9gAGc
voFqdg7JoLcqFZ4YL+2KRQ01IMwI5QsS7GZM0rZ2ht3OoqUo4JXE0pxQzl5AZjHo
Sw2734i1D58Ov1qFuSNEoEs6k6WNKD/mCCi4F86xApzOH9D4b2uFbyvFvAXJFlMM
c5mjnfQVrw0of9EHM87Bq62yIHs8Kkov0KJOPFqJQGihXx5OKR8l7XCPM9s7c2cA
emtqv/9DqqJohw6kbdDqX2tbtGC82VNnDxbLaIVSZSkEQ6W9Sw1S1TUx+uuepCVy
511Ub+lrQAp5oSKIp7SxOzkClvm2ohd7b/kAdXeFZkvDEYp95AKbR6a6FQydNJmm
OImu295uIydDNhcjucZXiNGcMwFGTlGYaQjl3/U5L+WvmGkoe0i5MJBIhtc3sj/D
n1FasXHmy5oC3mXDPNBEz24rZQqiLvolmWx0IiXlWh+J8mlEaQjmOOU3D3D6/8yi
R/tsVg/8bHOVGHv2Cpv7UGfIC9hmsE4XJtg/ZqEHMsRGQNe8Plo/OLBsW/xvezB/
YK72uHCquOj+UaDVSGDLfnd3IehEK1mjPv90LrbhieSYpNcqnNhYBH+0pu0ZMxy5
8+OgaCxKSZOOq3P/w2a8D3hzTBaIlu3NSu0ejJCWdZlJSDdVXch9wiokjGUxDlNT
+StnwgfURc6d9paTsrP2yZS2m3igrc8ZYzR3CXsReusSHyVedbDSHhtMz9HxkrMs
8JlWMt3JKDBT/kH2cw9XDv15XGtQGlRLyy9nHm0jUMyHzaLbIpyV+qTne+JYCmep
rhATnhDGs+PkPOUOv45po0Ywf9pGdpq+EOnobHzMnD7P5C1asqjipT1uykIY6Gx7
hS2kNitMNscJRsdFvaQCZ/c0NtoequKxMUsOL4AD9Jt61yP+tUMYocOP5VdeR3Qu
RLp73O8xha9FVytEaMuN9ycHXupvtWvg8SzyToziz2dsho0xZF8kc9FGgYMdSyfF
KLpOBLmWIKUQ5YDcg1rGaiL1NnSo/FNm1aRrXWj6fGgvQxFU139tx3kje1NWc8L5
O0VWbILQvBKWhQYkNDaLwJDAul1V/lq8P19eYjMWVxex9hIY0fO5smILcArDptWZ
i1SXm/2rBtkxkTG/NWmRO0r0PHmvKAJKVq9d+mCpV976MST4j0llF4NBKMgTIUJP
eVCvU/9vupFKIiuLwd1cCJlh+HCVun3Az4iBDGcLdjln3J97c5pJ68NL9XnRcwce
egcAAlVGjWte8dUwZ/zG4Xc81AkF1eJdykVKEv8APABflNSHL9Ho+vlq6jv4NG2M
dHT47ypwMr+pzju+bBHtSkKhkL1naS3jNuBr/oFzgZKxe9uTW0BY2+u7BbKU1kVc
H5P71XdRTL5gwpX/gAfQ6HosBU1fWZ/82+5mV9RY04RZd1rTm8qMTPpUiiIPZ8B0
ZVwyeNyENkq6YAgLqAdobGuHGu/AOKzHgKOW0oToamwsMBfxQzqZDcCPXG6tpHrP
zvtv9GTOizpekQAfwz88dEkk/N9k6hD8quoRqMQFyAAKlRo5dUzhiMCfH/HnwzFC
ZDJ1JhmAQUF3rKsQgyDPSmBDaQVVBm1c9rL5w4j1GvNCRcRFM0EAPcsKYkb9K+U+
uv2/yLKSrGHMUnfNpbN7jOD5JjK4sL2eGFeRTFKZ93sPyNrFRu+QV0ZW/1k+29bu
O5UntnmyOo8rVITXLQnQzUuXQZncIKhIjj6+FMBwlv5eNymqN7fLq/sKrNqr7gST
31dZl2K15JkgTs36LZF4wREygGgvWpwFjlf/8WeKzYBi9sY3O3j78K6XA5aXvnu5
zvybILjri7lF61HEV1AZmB5WghtUnpz6r4JghRpGKE3hMxT4bpD5yOnEPdN0Q5jQ
yzzM/H4mt15LMXXrQ/iF7l5WcP1hXdKmdM4Ov2KNTb6S1xihaaRHalVRa0iwWuF2
KCjnik0zQ6Bza4Qv4k+Xi/Ayuc8W6xY4WQSmMAS0u7WzPv/pwzR6c1XN6C4KAKWs
Bt8dn9+CAepnLrBv/XxLU65Ou4mIj1Xw/7nKEW0kbiGS7lBXY5UWQXNio52oymbQ
BTnvIXXzjww366+AUGG2Ggwj0p0bhoGJJjHc52W7HvGoG47Voo535buproHROy9a
mpJNmgvo/67xrRYpVjLSXUDF/Pyps2542nh75OxwC7BhBG+G3osDNtQK6t13i/0e
RCPSpBAbGhWGikfncC5RhlSBCdVGOACKi9EENCwmt0yY6k11IOTtedGKhSp5FUzb
WobZXg028WoHrc3XzQlV9c7jcnIPC7bM+lY7EHrbgsswzJ0q4NY0xpp5GMGJvgFz
tY15DWMDCzzJXhdjVqko8FF+zH0A68CZ1anpPcECJouUWG4jSVkBTUe2gk9b+DzP
FY6soG0+Va6dD8ucaZ0mbLSFbcW5t1K1F4yuv5/FxuELDNmIE/5O0Kze60gH3wp1
mqSmlzZN//kbvANMdPV/h68osWntXFz1+ZmIqgCO0CGuQrL7GHsZMKfw6ABIL7d/
B9XDAkvEinZ178ihpjh5XeYrvKe5wvG/zWQ5NDKEy0R6V4BlyEVmNSs4sZH4dRX0
ez1UsUlTNw8RnY2Adzu0OUc3A05nCNY3lmbT7g+viaqLMALzgOLwD+CGDC6TGvCs
xZ40zP4Wzm0jqDoGgNnVNkygyYtdmA5u1cBkz+6mlSND/68bOrKcRmtDiychN8IK
Af7T2qQ/AKUunaMWidYbgwC0os7vLH6p028jAMbQU+aCNVbAawUnZgByi188EZny
weYfx7r+xRCr3cUi2FPgI9bmF+fQFyvXy9x77dm7vj58dJhgXqT6/69ZMI3KhGMT
w5yYRQBWPhnpKffO2Pzrt5VKUG94bixuWpOcUPHOaip6tICnb/IzAvUsl35pxle1
rSFW3zRXwz1CEx84zbC7G8tcnCGjjL1ufjVmi49q8zx2rpJfNqrkUH3LJZu7Gp9/
mUyfuFDMHfW2Yfb2f6JznPJcUlh7LLaSLuLxKFk3kf9m38KumJqTPAvaeP/upPNo
j0FuTEhGPRckw/UrVNB2j5V0iwhegiHHtxllDetGWXszmcEGKFHORGx/+DepyEFw
W4+OWJd8ZKYNwiMvoUoo6niX8EQy3098FUMLsb0syK5Jgilk3SpakqDKQgqSZ3sl
3mckXgY8xTBfUihViH1+06od6m85gBxp1SBrTq5I33/m8VYNHR20ZOQB7/bbSYYF
6Yn/Nq1Gjq7sDg2ue13x23FzSkcGgSNBT6+t2Bb5nVqHSYFL6l5YesI6L5Lz/fzo
0e27bv4I3EDkMkFhI5kuceG453Usu+TfEKXCkXjxRhOgdxqHohOlvcife3fmGyBC
sN4YYfcWJWKzs3n4ikc+PTtbmnYmadMsJAHonEQtuoABmP6rTVoHbrUf3EfqlW4+
HvYP6AD2x0fgGvVm0PoM0fGVB8PUNztPHfPlpC6wF7vK8EdIsUTPOkR9lVWfc8Se
HJs8xMr5v1v9+G8SR980Ps+eVK+EhEaqilFyuhMXX2IeIMmdBGREKYA2gX2Yrgnm
4GRTrmW0cQOY9ikJffe0JnGnawq/giecjNPvgFOOaZyfzSqE1VoXG4KMfIcRsHmL
dJPvOCO7IIa7BYR+nWRVih9nK6HY3bWT2L2C7aDjB3CcdIf+hGESzFdgfJdzRaOX
8N4VHA8+RbhIzU7hCAUs9m3YQnmZ27rGThp2asiCnUbppVCDLBHExBa6cYHNmODk
NqPDY52GnlF8pULgOXj1YAME0CNY4B0461jjCixRzw+gV2hiliUR93mnNqV6T2GG
EiGYLUqReDis0NYsvtTi9iNy2ZNxFfH0DNKGsRmRUre1k0z77NtwQM7FfWeJANt8
tGcL+uoXC1nYHW9MyVU/MfotseNwA81q0aQu0XlZ4oLvTYxXk67sAtHJVrSHUxK3
XhrO4G12oJWEnLZsZTOPGtvMPb7XwZmaSJePgnya9y4Lg0GmAsj5q4pf9Eg/TPwH
te6fU+RgcxoZDPhPiaoHEQB2rSz8DsitZbvcBw5+CIsKAsfDOZeSYAUNtKqigj6J
uLnumTHi/5CdT1EHYNZEdVsfcCdx1gveV+qbQaQRfx/5RsovPpb7PRYZ+VAJok7r
7ehb66nZaiXKOvcu5diaeBqx6A32t6L4sHy5W0ujTrKrRgAo1Cs/j2/H83/Anh56
JcyLQ3cq1hm2QxUkUhq3fARPjPCLw5p1yj8o8wVT9Ta+PpH3hpFgp185L5zalvGz
bc6G4Ov1M8g+DBL0Ai6RszyWyWTYQXVHeaGCx+C5cZz3gX4sNfoGrQSbeKljOm+4
MXYNbB2swzZy74xBZ/i3q0H98XpdLfHfNCU+XwsZvu0lH+7pjOUHGDiuscEeYeiK
qJ/vn8+zCL3LOCokLWLY9FkiWldhOX9pH5Be1pRqgFavf57NfXZrRLgZhtu10NKR
Zv2p0VvWl1aHcfj2ToEWYJ41Zkbisrbj2S0XHiotYeqvvARSeFP0dm6vsn2rn/o5
PG8qMTQ/gXhgeqpAIKFUUNxe9OaK8VugKkdWJChy26ow28T9O0HLih3nSQWfHsIG
g0ScMuY+Zmu3sLTU+FqR2Qb/h4Kil6NulL2GRhzDL4ROHepNWAjhuv7iupystUbw
sd3T6LWNwNXovwIQF9zXy7640GfOL06vNO00Pks3B5uZ4uuWqYrG7AzcrE8BIMDx
oOLLJgezqKVmM59lvmA/yI4uz1/T1Rc7AGu9bk0yDxaooZHofDdieZF6FmG8qoqz
UNIwgNIf68CGgHeAsFQGLG4690flfrAiHjhl/rgBCKkoY1c+RWZQ+sNZ22nrCsp1
rxubOwOQdjdwSdzvyNMlZLkAiPKtbCAfGTH7W9lhpFf789opKO3Wg+aLeP8lxulZ
fLb+e/5Y22C5GUG6bfkxzLtJt2O5xwKarvh676IhqVRAKKQI6LRc2QRej3SFS/pV
m7tIziy+sOt6w5TQmX0c1pd9vVekO5DDiWLJT015pcXExzI5+3Vv/VZPwlDf3PDF
NYO02MIyDOAhpntmpi6NFl2d28uvMLgJOPL63b1IxqNKCgkyvlaUa9IfM69+EJve
tR2bZlJ/2qM9/WzJQADE4n1O5BN9miNAQPwg7R6ID3kux5/t4qBIFnMdnLmfCO8Z
6GlZnPyd4U2FVXv/31wceJuVOZOxgmx4D90YVDUEbDQuZMMWWtzdqzedN6DtYpEb
cBa2yJe5orAEtL5GaF6jZdWCTRmyWaHmbgHMGn7XZzmn4qZCas9OYcZuTCZBWAbq
HvkYHBQ4oLN5+Kz4PS2PkdDBR/mcHPuDUujyG1WxEj32loU72TZSBIR13NZGLs6a
ANjUbMMiyGNHYxJaZw04shFxYfP/MlOPgHTqO/+NNNcjic/CQAlKiHLJMqhm8zv1
WvkBm13Gl01VpzeWxkGK9wnQfQITbhsB7JgUaVSD+TQLDpr4+GQFgdrxGUEix8+B
vhoAfqOpENBftQCq1fIZRspf5sQYlibKxD/fFWKk/xXL3h+KqTWw2tpkTwcoo7oS
15+D5dxIhomVuh91Be+2Gctt9FZKKksL2MKK8Ghauu42DYXvwqGxzcRYQlvCiYg5
DaqoWRT3S2MnKRa39nLBJewkHkNkFdmIN0z8Vwlix9GCTiMyb1NTrqhVzgyaRAEB
vKVfUq8al5gKGjcvOmYUtOWANeTnkBE3bKQRhoajwV3KzRuhD8p/fdIZby+q9i0L
V3d90ljpUKE/3ZHNVvMHF2Gcv+eaaMgGU7u66zxpoThiO/xcZA8tSXPY399GgWY5
WA7bFRU6ov92SnFVH6XPIHUGbua3SSJSCUjGIwhRQ3HbtCKdXqfHvfrbHFZJWzgg
LbOT6PcDe9aJskwWnBacH3filK0/qyZuFAgiZmK5Jcei0/I8lOFpiXrHgFrJTsA0
L1SVIZs6tLzh5+YPywjqR90Ti6DJLZhHCR431s5uv+OZzUhjJASDaDXlA06SKKWa
kUUYbDbGVoTDIlDY/iury5E/FSeg7updq2PLCwCmQzRXzGEKEQROvNJSgkQ9ubrl
mXn8txstsSeqH2cuTc6hGJLXSRGBfLRJitxpGo+M/QqXaomepF8ToS6Xuk5239n5
MfHuSl7sC5y47rIXVbhiDcviYIsmrQQRPj4vF2ftZF+iX1t4MNJgLVTB8Hs7qPKK
+dsUbe3RiM1OlLQgHh1GSz5B8bF52pWzNNbOHRHt2VCTUWR73WpZJVCGL0lP8Qf2
T8tXmLU7arH4kutuoLI3dJZ8IS2hPJveAj7oLvBGJGvjAxt2aYpWM3+uW8uDOvX9
kWcxc0V8EwL311L2bGZbXi+p7MMvsAasGJGLraTCnRP0iErYWiQxDArbD152czBZ
DrAFavAj1tt2ODDIExJjV9I0Y+syIw1TNn0/u2DvH3hGSSZf0E1rnE+GLvjekuEk
ey6zd1tL7gmslWjZks0Zty8ATwmD9U85ZgXYFI9RBiH2InbnhYJcfWiXOoaH8XIN
7+B9HHEI8f9jWHnjobymM+WAMgf+B1L9h/fiFm/UmzCHFc9ZbKKSEne8JXiRg92T
+ES7FHTnitoeJM8ecF0h5LZrrLquDz2e/8MdGQF3Ldj3rWM+xy/Uo8zuVvRE1qcV
xReL+4Q4//WPd82nt55nnvqb5GFRDqH6KNQWHAIIgQiVQGcrXvoIpSUZ0xywLt9Z
yZftBdIpOPIrkj7uo7oUfkXwX3fnVPVhiDM2dd8YSCfb5VF6V1drswlmFrHP63KB
pZW/zp9AEvj2IOrG2MU4IbWTIG85xLN+s1JHdRlzGVxTopJNIzeV9IOHDKuKzuS7
8axN4s6TXST4eoJ730ypClDuQYzcYd0RziU1SG6lQuGsWMh8iqD4uo7p3Mvv9L+0
CFyCDCurBISBzGqWxG3hJKN0v6mInx/Dt8hVVuGto+4J0CTO1Ooul3+QwVJeVXEt
GXo9s56wT3uyBSGcVhDbeV+xDiAb6cjjCuU8v+25BOhojNNgeJ2lbnnCczkHrZJQ
psI+8EOdEjUYl+nx1BxCQ+XWnf49LGk1fNVEtcSdZOf1o0xrolE1Z6c8/DDk1TSO
sqw77dEsRb9QET1vKJeIG4LQDxph258eL9F5AjpuPgurNrbosZvRJRpddlORIwcy
IuyUzKPyho6ry4In379qQbV0xvIYj6rsMygxxHFByqUcw2Sv/Bq1ilGlhBCLqscB
jeobMfj3yqAcyFA26L1qzAFdeacmvTYgIaiYMpsipOgUANNc51c7ijb56qSCAQec
WCtznfPF7Bikq4QgPBkqlUXQSwyOD3V92TSugkOhKTBzNwOFwezXv8CRakOgIAAW
rvCeAPSAelw/pmWpqJ978Hc5JzdSGxgT7xYGjeMe2nCGrbzAddkyg32ollt6tdUI
IiVLU0SEEoRkx/R6JykwFPLzUdq0qGGF9erhBQQ7VPhRpQQ0DK/S0nDWIG89vS2Q
XuKBslxWeUkmGkAsqT/L9gvXukrXWynh90Z5qgtAXYEcsG8d+SNXltWjT87JUeAP
oDDDtURZA5QV0U9/kG+Xh2ftGtNxld5vWAwxIfoNvOMShy+D833YL1/wFM42pydO
xzhdGHfdifspQ7UEUUfVjb8U10raYklA4VcIrHN/sGZpbMu2GVV2xmazwNWEadA1
tMZceclqaoeiiG8O8s1gUc/WReZGbf5IYoUofDolcBrpKVAfzFTt1Q33fTVLt2Nl
gIydUzCRJm5gRf1RJsLn77JwUGVDIg1f3LpKu4P9S/u7LPrKtrwOekfWr3OwE8pF
d8a1ApBcB83mRFV5wEuMliGkUdFn2gmNwoLafPYdEHiXp9EYqkW7yneDveGN5W1A
H2JYkUDgXP1rDsLFIpSiL0H/8g2l6Y0Vi9INXeUeXR6a22EjTf3MJrycITEJOmZZ
ZVOBbZENgg1hvzZVj8WBQnw0mNIFaAJSFdv9KAcuJ2H3MkvI2duA865bmCtEoOhX
mV7eSlIxhtVHi2LtqlT5mZBcmvbd/veGuIBfYtL++Duv5m9WiOvCy6dUnsopwiqP
dkQzDjhFeGAMHVt/o04gb75VydW6uu7oLXDlEl87IKuG1WMhnxuweENAlso4AEus
iX7boViOkxBtuj0fBbMLrPGmVI7/zV88xV5vo69YHLAek/FkvIloOlKTZ0po3kgO
ugv1rzzEudJ7GAjdv15UP7YVtDMd8gu4BEXSRVei9MQW1q6ZrUZ3sBySo5BEI78F
ZMl/9povUQ+KZ2ka4T5Iku2Eqi3TP6X+dOIXWuAIaaxJxLz1QT/bfFDVMc09oRKN
Q8sF+QnXm+wdvazOpEpjMNTrmjwLvAZwf1Ge0v5gKZZ4ymc00Nl0eFI39QQgMGJO
1gaBP3WCSGubczFPm03WQQo1Mvud7LMYNwhW/NBC8u2WlzlO8eIMB3gn3Wud9Cxs
Z33bHMbIpmcoJF8I6BHbA/0OuZIiaRRl1e2olIk/uPCAdw1NSO6T4ottC+tVTK+w
qjKjZBsXEVIb8un0iBL/GuWautCTgYPpAl/kbIAPg12YV+O4PQW0v94+F5jJ4IcL
ScH4BGYUX4s2egzcBpcntNpIqyMuaEwnu8oEPTYIbEX0Y+65di160xdmVoqyX+/V
MvuHZuV172Z6CrL2u7H/SSygPOh3IxbBBJWP7N55znRG8VyeYSuFrQa10cHqDhIu
VD6VUxkfEZJzpP07QYgqSMGnBo1TwiHgKkYbj432Ze2iVAyJgQXs/v8h2ei7xoSu
6pZ/9CoZvJOBGas31drH6ICR1sqGbdFkAUbuMPHICLD2MQaOcSa7+5iV2YM7eAiJ
+FpqHegAooVT3awnSgsiK9cF+yLjzhy3sRNHd5lLsn6SMRrTNQy2m9TBG16zPtGy
qZdqo9+axCntu/JIYgvxt5qCZFX0wfUQA8WeKh5VTT1pWObLQkGbYQQu+MkxvTEK
WyPzk4eyYNLM34t+HiN0xk5LI0F2y3iEDUQuxLON8zAXYKLscp+9cO6hF1Bggywd
jmkDBv/biVYAKkGjVYFAZYJYRBXfmP5y4Ad2uvneKwm6p//mbneaaOyxYbBRp4u7
vYaJYXIGoaBNmaD00bp/HSsUb06pC+W+OHjCjTT5P7gTlgxi53xTFJ7WgFP8zRlm
EeP8UsPXCOguQJOXZc8owk43bA+DJuu0NXqXVlpCmUYlnRk1hD4Cl5X2V7mlcISl
Sjkt4z6IFS3CpkLl/fPXydVHGMBg8vxgaE6ZlfpUDONw07vvd5sxRi02+gjgDn8B
LuG672yydBi6Lba/wZYC9jPwb/ENSY29Q/K8YVlD6v/9BWPbN8dpKDLvLpRTJXiK
onwzAOprUw9UHYoOdDmTXuDUjH6KSNCwQCr3hbo6Zb5RnZt5tbHCHdBrL1vTFEZ+
BigNMrt6sE/Q/3hwtw0EkAGmT8QWqWbihrMnMJ+lflf60qJxzlEWjF5eSzlpBIs7
MbyepSj2oE8GyDlekb+YsIIxLp1g+nu1+qaGoqkaGjSsMO0mcOgQxJ/sAiXUDGb9
w+cFxxF7EJnpJwP8b5he73OJRG328cpBg0uqcBD42kqQgtJgdFdd+9vkzrJZsqvN
QZO6wNN4TFCKE/93miDNpFwe7gByZ5Oe5seOdkTByPg0yjsMtEyviKK1u7lt+AEh
Bt5Ud8VwtaR/t0FflSlxBYdeO/YGb2fgk80NrNaqU3bBNTMdd74gazmpHJu4iJwt
nG2FxG6F2mRMHtRyX3jH3gStd5pK+tQ28AFvmvlPmsDEY9gGEFp0Au/2Hg4MjrM/
c3feWEyEigsB2p76l/SP+4T+Z3I8irkY4Nd5a9KqEazvXhnZzkkOCARD86OoHzxa
DUli0d+MkhFUt+vZHJTiVkIqm1MnUO6LkbJzanaQM+SmX8bslQRALtbmV6BcAwFb
Xr5OmPf3N8f0r3divCzKnN2tKyUBDMCuJ3uCsIEydeyPDnIZvk5TXSma53Q8fWSw
vVqFs5YbpH96fa8cRBnMKmCJP26vFGJxRH4CF9t/jn4IkPLvOqVHy91LujvBoZg6
XxCdTUC1DXn5+CSNUvSvXssAjrDyBF0AmPLp4EDae1sMKV5ufq1ig/7f/M204N90
QFZ+W7okKs+T/dCSYNWkPTzd3dLqDLzbidSQ10ZQp6ie3lAGrXo7/hEU5Wr2zbY0
1wEidNlABrQD9HGhVImo7Mlsbjl5KJdNX4E13J2ex5gS3axN8LuabhwQ3Ju9Pf6u
4P+kz5Mw3+pcjkmJXQuKDC2RQi2rktW2/0493XEQsjD9VDMEL8ysrOqKrprdk4hJ
9jTmvedvDIHahyd/0KFj3nsSiUTV6OVQ5aMo57QTW0tAqUDyItVtMCZhLIKsPyWq
byB6eB6evJ3eYmoZiMQyjxRiUkyTgAJ1MGd2eXJ+TvrRXI6UUlOKVpMtLrX243PJ
NMaEBMRYzCtDM4naJKW20orWO5FSSkBniAHBOkHrrySlRR8P8400jyyyJ24leTaj
8LCIznou/FHJK5Bp+QgD8H92aNRZgHFKeWxkKRDwH4KxL3vdSpVhnKDTalxMGPFk
Gv7/N82R9X/WoLRyK4Enya6a9DgiCl/FkU/iNiS1Qydm32DMcAFXBW2ZOw2Y8WX2
thRrKjwVSH1GJnHgKCUbiUBbcOSF0UiXIR2F8ZHaMZ5ICwoWiTP0+a3RLL+GKPor
cbBT4Vk7khD58SM5eIZd2gfo2gvXvPJDbb6bZuxGRvhA6xdKw2eG/8QngLGdaWFR
mHsT2JZKmPequYMPDC/ZkBDfN6yjVCWsun+K8M0aw6TKq5xXBHhMm2hdftse9BVz
e0UIrjHN3s9loogA0rnLynyMXcVc4h0IQ6fQsfD86qDkukXJe/F74XulOF35Mloe
mgkLfdzJRrozbLEbEAbtOWARSoognJw5HtKSt9e/EBVLbrB626HOziGCcxjpLsMv
cjPH8oshfHYuPrJ0ED4cCgMxnPNexe+iW6EyDSt0fe/aVpDqu/yHwdI5cqQBbTwE
dMFpgrXaE990gqdN4rvU956iwDZ+sdgE90jexx5iRFEc6QaYhU2zjK41aYtYdQbH
a0ab/HpVjd7ZYePemkxylWv3KrBPWEX5N7XPgYsRB3ge7B28J1TawdJh7wkJUil8
va9XE7+GM9eoTKM3pBIcwIQOh4Nl6Gv5RRQmFzgblsN5S3mxChIx4FguEnDqd51U
jT+YVwS9+2Uvi2OAHYohCWiyyTLi1/kFet3anwUf/TfsfchRFqAz92lQ29xpSHLm
4RAKPPuUVVYDgXuMM1sBN+MqEksMi4iUL8Qz0loCY9CvZEiKld5yUpS4xEjzoj/J
IoIGr9SoPiXn1gD89jJ4Y1THjh8kBMhs+7jSxaRxScqlgmJKVwCs8/4VbhFlEwOX
871/UtcEbfxVrwKswBa56Y+cyLay60quudI3ff6XAWD9/HocZtEC4jpnsSPjL3Vm
VW1PVy/a/Gjp8gohZWE9IYt4zodJYJVcI04/LDgydtEWi/WyPWpl7M4qD1cz30DI
LMh5odDEvc/S1ofDxTyTiLBT8crakMXA1MfljZr+o4A6zBQAKp4kVskcgm8tWYHb
ED6Y5joj/yzMScCzSUixiYsfOXI+b9JvfjM9I6wB0re3ObIn/rHdi6qIXXR0ZD8+
XhV7k9wr/Pp5C738Q//bVvR3OcJpxTzJSASRexiqtZ50GSq0LwG7yrcbe4PRFA1j
/BFJydy361egVzPcOVoNtq3aFjHvuyZbXq1yx0GSToyvMiHxcMNT6HE50yNzV3UM
EzrapvBEuiwHacFrhFJniAerOdTO1Aw2Pm90R/YURNP80iv7FztDwR1VeikIykH0
xDeUKAdEbTWRTDqJlcoUK2Ex3cLUIvlsaPI970grQ9lJn/rO+rMRj1lZA4MxuWop
ChxWjH10tEDlVKcPLLskIl/JR9gGvAqcMb6tMPzSiy36HIVtUigVpHp31SstjEZP
nTNPedO4nhxeJUKIQhQS8/SNliLI+ZpcwV090vhqZU5Cav5YFl3vHKX5wvdWwbBX
NY5ILhqMty9z+d+oTTnnrq8ZwMiNMnUbhT1jqBwuZhFHSysQqq0woeQ3HEA+Ezs5
YCKDqRMPfQHVoNDizd3ub5d2r3+InGNdPl6+A4GyBG+dCBd/feLlP3AdXU8dOlBR
k+PV0GotyDLOeByhni5bB1Hzcs6IzFbJ4KNaTiHKoHFXFsINnn4L/i1bLpYLSkgL
UROVzjzMna1IRT/Ttfo7PSHNcM9pke4fDuHgZG/Uxh6zSYDiwEafnmDKtEao4njt
MVuSlA0xp0uhQ/HmHHkpT3+DT3eVYyvcKJSBH/WqACtVHbddSLXp/l8sxppKPfe9
527srTW9pDVWyPGqCtPvAETneRolv7CxbsQKbuUEs0r4CnR4Tk6SYgOZuydxLRwu
E6GiU1yRzyyiyBWbrZec/bsA3yghtlHtaFcP+pePBzGkY0wr6mlM1dMaReJe7S3i
5yCdilDtdV33iy8ujHFJOWYhqpQfuAGs6vrB83Y1hliKOsAKNAR8KRzxWC75G9cD
bu1Ut1rbkv1pdXBTuIfujJAy2kdpRLUVKy8wfzCQyCnMVQjuaIHc5Sf1QR6i9sko
8LISBvzV6rHFBOqPFeAtnqc4YQjnsYYOs36ts78SykNov2/42z9AanAp5ES0fRR4
NX2cJqbuQn/fXULgWI8Aiq5nbD3gR3/Z2MhXjlieqCn8gHjOkBKLvliluuPhwQ8o
ozCSHOXTzfyoU3HoHnzyLNPBxV3hu6V2M1Jmp0PIQZxYDAqAG0w/wIdU0/I9XVzn
u/NF0oYvSM2/8ZYkwHFox23g+6dMkBYCSWcmZ0mUsMuz7cbbhZ8xAMXq7a5GYyQ4
iIxw0zGnFzYqd2LouEQZVo5ol7sVMSI2oK9BK+QMtZz+d/EAoUKaOnP81Z+Vvoad
yNvkDk+1d8UOlRzHiUVan2VAO46SilOUgUv5wlZg5FWjAT8rLmkBlCiOoBCr1AwN
uvCDdXxOASx6UjBQ9H4C7VdHrWtNjCpAkFrSaBbKAYeKPeQgm+zKkSCwH8gZs6Bt
4SodOZiEyNDFh15ByJFrDfC/r/RGsAO6tYETbbjpCkpg9uXRGytg+mCXGsZuhwXk
zMT4rQpxpiJH/5DaJeMbrPYOxfx9G/jlbm9Gkj0vmegmHMnC7l3ojl8ICU7lCdYw
EcTderJeMcI4xtZ+KQ+eI9kYAggBvz55x2NCYnIhEGTv16jEs3ONnnygVBEfs7/C
e/7ru2aIS6y+CQ3d/lJtJoNlb2PkfzzaLbAcjVcc2GkzmvEEsMWe2exKCKoUuPVv
kJ3LkrPUOl8oiFlQCNTD2gRhQ4aPXmXgL8cMwGacVeIbnnCXn3zL2pLLy/swi2XW
rzNS4r0qc7I2shp6L7LXS+P+JAMFnTEQRpxvcG8hJj61+IpyBg9eLLydI8u/MQjG
906FFyIheoZAyFGQLvoVK0pZSKGWMLGPqGKywrfETidB0BDe9npQmPfV3Y5v0rm2
OCFfUFs0urE6DabkCKjKgMkNzmJwjOiNQFs7TadY5/Kqfv3tz0c/8fYU0Qn139yI
ihUa5KvjmIJbsfxultckgmze4mE8RDXqoPB47VJ/InZDGFUDkmcn+a/arH7997fY
XyqtCWTQrC730L0JfLaO2JY4iFs2BP/6jTjiRSSwALROOTNIJlm8ueZMYYzxpc/D
yKLigjJ1ABFmJCTW6RP10FMukipNo/clA3yWtNxphsz5p3fWMlWh41J0KuOaJlvS
aWUl+JTbJScoPvUCsXCGblqPIJ6mTTAYcMo6MXll7JRN6S3jfKoTTFpN5IEPZI9k
PAYnKdUkvALQqwfcJudR7FuVciJ+mk9z9aKU+H6sMRyVLKqoa7H+mWgQhiuLZJ1U
icX6QIT01dA7jbrYKxA5lJHU6Y9Sn/6X+CsDwEkL4UD8SsKt1z9MKNHMbIOPaTHr
10JgKFZ9Ux9c3ZrFbeFyV+/VWrD8O1kAuUw9az3rnAzO78A4N7HSG+nFBqajWyvo
OAXVLIlQE8cfVMvsHreR4x6GCTQqfl8Ci9JN++GJqx1PYd2ePNdTNAfaNqRHJeaC
OPaLEyQ1U7dDVLDf+/WjdZ1VRqIdElZhksCvBnrgMyjkQvtrfVPkQd3T+yEa8rXK
s9tLNt1ix9AyzRIXxRoL1QEkDaeGlY0rE4LZCJLdFO7CA2iaKprHOzQPNYL+vuME
oOXl9FZ/wJEwmLlHAXOC5UW0h2yfht+wTAJtfCzk0SVw3VrNDH1Nv9KknOmX4VrD
kCxYM8VDpxUJL0N+CoXVHX0Ul0uCKOjy+UFga87WHeOmvFwYuxTVOFsHwQize3Ac
zSiAwLibGAS7cu5j7/ASQuKLBBa22BF4Q5pB97bVB4TT+lEjC5QPizjE9ye36xzr
ulJZYcFvbPEIjDss4U+h5xSvHWPkDfDwBu3dF57c9h3jbQy6xvSfsao8g7YR9LYH
xy1qPevrIxx9jCxm6L9ZX+KoPrIaJx0UrOBxSemWD7GM3HPgnaiqLR2HPL/m79a2
I9sXBVb7m0pH/C3fWrabsBGiSAGoJ9C41I6ebc4n/gx7FRS7Uva9cPVz++4x5biw
GHtvdpZ1VbqH52DTjX+eYgZpgIBrbUgGRWia41Uhh5QvpobquTbBvfqrStJLRe/t
iF7s35mg643s5jXkE+1w4MxwGCr5aNJXMhcyMvmXyK/+fCd6lJKyiHqwzryOKR7B
Y47d7ByVJF49F5MHTIq17dSRRoHyq1g6E/QTrjnes33ZJC7kignfnW32dw8lkhZS
PVAdMVzNDZo6gjTHDFAoAMV2AHvIG4B0L/Pu3I9t+uuaKoFRGKWMLl9+5Fj1t9Xu
S9nbBjCGnoYdpADW8RqwrYOvhDeWxJxhAlfgIe+GYBW8tRnhjcv8qJOS6j5eRomT
iaHhPBiAQ1gS5RnEqyeHGnpV9GC1PQa+zAQ0wIBNrmyRWqjWDPmgLvtvnFAF8iuM
dGXcuV6zEhCB8aEKjJPHS/lQFDjUvEySotLpEwVO/lQyR2WumMKlkKoUNCmWkStn
imtx48ZHsFGjm2/OsK5LNXP4zdIg4Edl4NvUGYGCSqdelitMIqXvbf1k5ne9eFip
ub+flBD11IkU8Gluh4w/CMr+5yIy8vjhtd35N3qT+4A+8kjG17m2KPbDrkV1snP4
FvK5Th4mY6bPEgCuLmzXQwQO+xPtC8qAo0zkG3jFiEgW/aR7ZaWUqxMyAASMeum5
2fBYjQVYyzQN6JwI+H54PKifk/Q7mDCusymuHVAEauNW8x9yGYOikCyCbHsxe/MN
cl0VmSY+W7Q2pqWRAAzuzSixBqn3H9rng9rConZ0bt5DcD+yTNBrA8S0ZXSCeisx
yxOodPKByJ8RZ7wqezPWn0zoCNkXgGaAedlF/jfooebScJ2XWyak8a17OTK7SFnz
hcTNsMGGt2nnPXEkjImw0NpmQClD7idx7YnTzwkWCvpyMgvx2zbk/pdY8dBLmPxP
FLaNdJe+uwYAMPv1UzcwrcSVRz6xdNBVPZiJT/MFOr4xltZWvqHXT8CJQeeSLTIu
HUn1XahnCDMZURdOCKfHo6RJkAE4bPSj2W7p5xJU4g1WiJBJ4Q5oyfW7NsIOxQpS
uLbat4ZQTO62H0BgnYaWhk53Pyma50NWbc1JG3IYXEC+L231jHImQLyP2NNif0dr
4kpDR7yynodiL1EGQo5IJiWRm23ZxtXDkAINO3tcD8za3VCYDY3d89OrSvRVxpbn
Ze3wSMV68iN5b+3xUyepwpZ1yMrQmSBetOWGCdNZLSVvhonpJos+bZiLkIA3H4U4
kzhBnoakosRjxHUDgJG91RHSY3utqmxHojncggxHVvkWPgRd08xuRgvOi2CetWn3
e1q3iI4S4Qbvx52NCwe6GdQFmZO+voAaoNs+l4KTFUthITAW3p0oxVSaX6IRqLXr
4t0klRRygVWoHDjvze3hRceT+1f0OSsOWFcwBeDCLjHuyZFc5Q2zECUzHK4/+tPZ
AX042FzIQBLEuQOq2F5fH9fdxBv5olZ8DT8M7/leARtnGOSLvF4hKRqynZps6QJ2
IaDfBJo6LrHUnV8NqxYXUiyraKtkEQZOnsUbovgnY4v6P8P1Ogr2f9s6Hx8zIL1G
dEltAraWv7uzWybOobG88WFDCAhoCjAL22Adjk8h4d/WaKQ5ZhbIe9n1GDmddFNT
+aINDsARHqwdRPiuwNJvdq3rqo9bribBk1GAepvqdUfzTpl5iwBpJcQyY54WGD7j
MOBRMbDEPby12hR8Ms4e26VTx+u5UdcNGX3R1tXMKdKjQX1wMC7tLnByals3CrL8
mTpgM0q3p4zGCES5gr8o9hBZRbaSTXBWaxsRio08qyc79DmXWBBqb2i0i50/qqzE
x9G9oF7WziH/OY+gtTIN7jz2UGgCA7F31C1FXsWy+Mdho7gMPsQpOZLmXg5lk/Hw
1AG4Kxde2yB609RFrxvbeky272uBK6+FMvfe1LwVNQgN8DfM8jqfhKYuwU7p5Ngc
GFWCbkYnEn2rTsRebwdCYkNG/h4t2Ul4gz3uHmheFFfug/A6wm9WQVOE9hwlWPgv
y5Q/8B1jtAsJDj+v2tWd+yNJZ4sN676Zh6WWSU1PIyMIFXks1hDpkpHDax3DdWss
H2AxzsCp9m1SSASO8xH3DH914pokSHkGwq3t8aqboxisGgyR3TFvOAwzA8WQZRHA
HR7zjamMlPZhlHavVfv0lX2FblKvzsIK/d9+w6CsShBgK6uiKhmu5pffmtUe6H+y
vi57V1pYpchBUYjFa3pO3b/Yz94MwnQ2sqhz27Q2jVy1vswhxOpiG1jdjIkH9Qvb
1H0jSJSuKRKc7ukDDK+oqwiiC4EAVwrrVLE4CIjmkvP8dGyHsa1Gte3OD9XHM0Wp
8VK4Muf8lYQZduS34eL0PWm3WkBQmVhMEvFTBeAakGKGcgEXPEl0gtcMATQt2KPT
zErM/6AY2L+B9HEc8RheiZXO2BSgvrRgub2WikNa/7tCNVfG8GADXRN7x7B38qn3
1xgvL+kSzTCL266uEuQ4lIcRYe8onpdBn6oGfz0yYegY67cJ7vNsBXFAeuImQ4zM
uJSXm61qHoxJrwOvmV1HFzFW/E0JenEclwi49jvjgUvHz/sMAflzSE4Vm0AqNOLl
UoTwfESxj9v/zoUw865YNTb4MUB9yCqHbAUoyj1mPtQLeOK5wS/w1KVzx2pzkzpF
zawzmfLAM6EiorgqVbRIBGJwuNSOL+V4dgCn06D+4yigygHH9HHLQsJ2nj6fXm+G
sPHnBx5bjhAdPsexQW0lBVR4z7n9NZnjbA40gYrbO6M0RH36tFfreyVCb1skZaRU
i3yKzwmWMd4MlhRYkSg8o9oc+HlHaYgrDOJTdsChZVTkCQ7aQYx8uGYPQ99Tej+M
3FOAsj0CtY1UfV5KUCJJGRFlwHlyRzLGbO+RomZmynr14LvVKfrzVFiz9QBBlgxI
mCbXQxuKTfnH5VkeNkmZrATOdj9xPEBKIBocJfttwmWdo6t8QDWxim8A4DysNK5c
zsKxgT581VSCW00v1rSPgYoN3QARh86pTObTHUq0eONd59sg7UiEOV2WZVSt/Nuw
dK0HBx4qbgZAYTIYsHZz/Rc+Yi2yx9QowFp8lELhiTpOr9xjQ2AAlhroeO3lG6dc
NnYU6C3VCabVB6M8AKuhVzom2lwypmkIYUrIITNa2w9GMqZsLNqb5XDlt5YRCC73
unsf+Rj2XCTd23QlENM8NnV2/usfwnmg4Vut/GF+3D64xMigox5tXBI7OaqaJYhZ
P6yYp39ed3JIA5fidbWXADuI+2loc5PADmtRliJrw+bWkCrcpZWFj154VAqZzYsV
VvZRKagqjmTjxYCR0Lm57YpVFHynAomefQEUq+nmN3k5kM0ySkbxamGM9Mmr4EDP
0iS4YUkjGrYzgYR1QXqTqtj7peeB16x6Mg9Jv2JnusKZ+nG2cvwpflJPkeWlv5d4
2Jc4xGTcGym9anIzK9ZthGmo7qeMyJkMEao0IBKfJGWA9y+krQrFCfeNkjwc/h2m
MwLrERhqlLeeqcQDP2/jEVJAVRSTcbou6nONWx4jn5kucMnGldHtWixvyXOJVlzz
UDPxIQigbix+ZMnTKr9NoZjXZekqRcXVlpSCvjuSkDTsQjWyNZpIikohZlmmXEfa
z/qhCgiwDvfbfglryzlPFEumtW1mB4tbdzsJCIRjYZoA+qx8weiVjs3s/hmqt4q4
yBydHCymuIeNBflFE/NmfzpLwEJjEPEFGTgBbEV9DhaCzd3m3zQ8CCWRXRIdibau
D64Upg4nI7WItTPHmpQhserxc0PJMSP0lIMw2JfbOOxfkHKkdeFgKk/ModguvAA2
L+YjhvsWrBcaZdwTrA0G7g48hkhf2UDtWJ012lSe8GgkUaHQ3Mv4N60VlsPNBuqE
oYFZS1kJJssQQAjjPdDNyUClCcrDWPVwKqPwRbz32PncfPzrFWbO5sAm99m6EYHE
EkBk6BSpn4VQbFSEUfLqAo0osfJALXlh4Ez7y+M+f5KI9N1gZe3EgeR8q128M1nM
zRxYvaH+49lzw3XbXGX1AZqvLIMeP0luL1XtezooFXiGzReINKjBA45UZoI7u2Aq
19HLm+wVj4tG5tw6SE9NUfWpZ9ldh273CWLUM76/3RB563tFBOBE1+egvpXf0FX8
RAv2un+5vrKjHwIbVdoPFDZQ07DHMsnCXUgMYGzra1cQ6k2BWvftyYObcShj3YmG
EVdxh2mLELFmjYhvnwcWA8UGq8UD0J7MIiHe+XR5G7QKq7aEOSyZ4sxN7yFQDC3C
WacvdmYFiBeFURh3LK7F/aZvr0xEyQIMDaWJ1mHu2ckIGmLahtAm6edbE5GgdLa9
MEXZRa088IPbg3xGOFfQWS1mLawKJuQTYpagBrz8CCNa7WjgnK2HYt0kChZiF4ai
ZHNoemPg7N9ET/5uqGirGdDsqmFdFVNQG/rUtmUtDz1LK47MWvvPyO8BvvrG5gqM
8DNKIUuQMBeONvRcxxlVvBG4nj0WwiDwuV1QHLFIRX0iwWDsgtm1sQ3ypRqzIUY9
feuuIad5YYfPIjNphzTWU9VJZpaprlgSVU7/GDUV5kM43UBCE+aa1prfLcmumjeZ
W53L3Fj3Hbt564DKxp9BBAlviow6L+fDaSbvUDsnpYwKEaMZrluSTLk/CArBCgWz
KcWvK3TEQiJRidX4s5ltz8fCNKJ2qr4IgdCJJAIQKY5jYtQvkXsJTlgHZIR9hdvf
bUJBXf14wpNMDIA/Tvs2iTOBnxDd6fnbHGxhAWUdBxQpCfrkt0qrhONdRP+GLBcY
BbzUDO4VDoArYrtBqFLuEurL3YLFSL7M2js4zIjSuuu6YHoK+u2uqdpszfPMxoyi
vRbid8/DSUbF3AHXr1EGRBbb7UwyEC2e4uuxKbU+B3NhEO+oLrgA87axq3ejjOmT
Zz3VR2cls8WgIXP5R6ag7WYZPzPdCPz4ghXe6VqL5/h+1zAQFfGzyM++W8af5swi
BJIsP7tOi4MzPDvuTVCrlFpxoRefGv0NTG+ctsdchrRMRsXyy+M2Gf42seT4XMYi
V7GEkcrbg+1hdMRqOTsR+yxje6IyCl/M5se2PfiGHKYHsbdBuGRmwKKFLhcQPxha
JYrzLMd4Prvf5xH4eTZ/e/eq0PGKKe5RBxcCKMtWYTCJIYxNdwrgIFQZfvUkL4DJ
u4I+NidvtguYjeY1L3BqQigQKRwb5+IDfOnqia5LVQUzLEzCv43RTAzQmHoFYd1K
VjKlXUSXsU4NzfF8r6BqfALA3XAvAHgRHrSYbjRXKsXCWdsnUBeaanNDQUiEcpVo
WcnWO3Xt6OvXeseN+G2SV6/McJ3r9XNWYeRH4R0ZNwKLnJrk9vQ9/NXaHpFu9v20
HDgpZoDlgjapCauRhjIgXn4e0HsW0KkiUComn5cL1LJ4i+io+fG0dbYtOI0+rBRe
twmIgpEQq8GypUbED4XBXKxYbJ4BtX5a+D4Jb45HIbYFl403PZW9xwvYNM/UaoIm
XefJrVKRLFAgL7ZWHa9KmCqZ1JccVq/QQvDPI8gFGrU5XSNetNLlwv8GMaW4NpnU
9sbENruTVsRfrh2kI4sJKPNp+ClYPQrzNKQPq8wLn2U217XqS+krSCqEuPoDDwwn
G7GSACzAp67Ow83tjzCQLRTRmNj38wvVVWCieiU4g4QofWNV1lDwWt7FozXPONLr
dWZ3wki3o2AkUI7TvYgHEYXw/mEcPP7p+TuxEMxsTl3LD3G7cFJ+wrcFHNINMVFX
BeaYsI5IplFiuEGaXdk20JU+72yP0lhPS2tv8VpB0lhbZ6ctlTvTFLqtCnNWTjda
l2VdmUnMEfNebEfpHH/Ku3L/cxChvbzo6Ag0ooiqi7HhVsvG9HmyB/crDgBLm6Cu
u4O30Bc057K75mhYrK2vTbErbm5LdJA1HPOJVsJggthNsmX+9bep/2SJVwpn4dCi
moygKsxOiMG/g23c3f8+OoxpbkpN3ymRBhK5nFN5RjH9mignUKsA6APBAzFj3iia
qbY5MyG4udB+bWMljbGBI1sMSohYFzgUHcsJgx5j2RZTUlUyJzm2n+w4s87cQWqw
sKbORlP5LOXmhW+IQOELITM5j4qfGb7TdKaTeQw6ZfBJjlFFUzG1VinKjidhMQHz
lMjw0ZKkEHu/qrQvC3SXaTrEmNqM+lU5dPZtEwjAokqtGnxHGHg8uaJg94a4VMlL
EJxLkFFtxynmop9JKNQMfC8AwWVh7E7NjEWrtIwENOKXXnfPMMOFGQfmdArG3uAt
8oCTEQLnnXKaYE0heuBqYJ3oLZFoUmms29WMEzLsFOJ0RT6sTJKy4bn0fGaZzpnt
50NetDObmlSdC0HfaP1EQtpt6/cpp+/OUuTyp9YSAw5Ak8ZzE9lTkV4KIJhMBAMS
u0RjgJiN6D3Z/P1kIsbBwGw3AjQ884EKGedVKf787DK2UO6cs42cPJ9dYBZlq2v4
Er/0tDNUVIoWh/CqRGKEqUh/6Y9JHv4Z7SqKY3L1bSxQacHTtqJ6+8g+4n+ZVqhi
FTScDvCvFNS5+A7j8mg9A0m7W/oRuDvWlUbEtoKa3pheaIue+a7+cH9JGLToc8v2
N526Of+4OL3OmkA4Ls5FARgGIfcknLnpvzMW9W8t8mz8IqDsKg0OSUcNbYmHqRi7
QKRsIe/9axDVTRhKHz/dxNaQL3SpzGqFyf/pUN96vDeh7WHtN8ml8A5ejfZMp6va
tGXCcuAunPJVOfWIpoPuqYJVL2BxFsXJIjKt4bd+vkEpXnYvyz8faSPf6rtHbXGU
hNvYA3YeZnK7YJrKtHfUzAuNDPlNW0hYGdRBQJ533SVr1OSpmyKLHnmOQmR/QUSM
Nu992ry7ueqVPscOJPWXTi3PISZ8xaU259pRSmrnByDb9/i4FXUs20bx605amEUu
mND182+YsFkZS+AiWi6QbGPg2wxSjA5HpY/wdVt+WBwgJ2I+c7TWw/mkxRvBJSRx
Jpx6m2H2aR9CLb8erL9aRX2GjJVHAnDlNHxwUzX6q0Tb0ZiNev83zb7AeQSu/j8J
irbmrTlQh+zmYYI0wBfPqGKj86SbZ7v1Rs8jqrUkUAocTCA3RxvcJ+Dc+khk1pTI
vXHvtqoE8JVvZooFwlRPPtU+WFgPDuBKduAR1zUYmO+mgLI/OMaHAv4RXTfcrG0u
30w30qRVk9RwrkS+MyhKdn324ztTkXkIzuxT1LH8hvT8LobOlhn9i+e9po4TwYhk
LSPwA1f8LneMbw0hG+J7TwXXX2cagogDzoxncbSUNrTUBHuG2/DmLTEg6wPLy8pO
2jdcwZ3p+9oiw2gQmifm+mdCh50aLs/bOggNfZaH4IbDR6c5aQsHUN1KFHywAcB3
V4BGvnD9qgufUkRciiCGGN3HWzwUUIFfB8T1d7QTi6xLJm0oCBwcufUwz5CSojwd
I63T2/PjGWZ5noMMBRXYfIkQTRo8KrAtGjcQrC/4IlEh8KLOyP+SEC2NJkCGqjdv
bDEKbSFCgBWNWh1XXXSk254SSBSN1DMLCTjMFn8tcEBc4vpniL7ZzK4F0PjDQ2xs
Pi0L7Dm90JgZoRFTLJ8dyXLZPhg2UcwYknWbigBAsHzi7P+Sv8FWIXmIv0W83JHs
Bc/Dpfe24dO0H4BdBN1MThJnh5Ijb2cw2X6QkoiYyS9eVDeztGhvCODEVTbgMpro
H21q1LC8/bUqjWN7fgS/a3K7bxU2INKetNa+TGgWAmGGqNpavUiCLtET0jl796+B
l4+rQzSRpcCo9ffzeo/J6uvbikmcHmNGZFgFmx81K6QREMQygh+iXrjyAkmzTgqb
amxzFQ1+7NsW6MxQwNaK1Tk9+1vx8wGIGXnCi7GJfaC7xekJbWnCPduuG+5qGxAE
A6VsciCCGmAVTIcfZFvVXq1dRw4vJKZwcxvVYnXsAEf6cm40jJUbdAFoh4l5yjOo
FsSwHSyBvfuJf3HNWLz5sh/i708pSJ/aQr1YgHxZMYJl9463EGIdiEtmMxkTfH8A
SXHWzaNf1r3OCS0Yq4TT74852GYuJ5paWaDHgaKvPOdpVwYD4pC/bGcR9WsJ0/MJ
Chg5JICCowdveIVcXi/T5sWY1+B58vut/DSN5OrRGuW1tpleXwv+e37Xy91h/kHC
Duh4ikWzGygok5rs062KI9ii+GSj/Uni7VnhHP+Z17o4q99gHTa8J6HKNpOG/6If
CKNySvoEukqWknXcOjLb4LIVz4fWbL84Yjyu9dZBY/PMnXN0rAKjTnkwyyTcVArN
OaYx3HgTaVhPeaMMF+5bStnfyLAcm5fTgCTgictr7tCxPdIMHPzqXdrykd+couTy
qitb9HMbzf2DRkD0lySYvRRQ5KHWkBT0dH+bPg+MRckYFfi8y3Xn8yAnPgal21rh
t6ScqP35nTDXP046GQ0auWOWarCQFSnwVDbL63lq9annkJdfFH3wU7FgI+sGN2kf
qrDHCu+RHCb5Xna6uHnv1aUFjVK3+LRCl2ZmJb2ZYoezQI/fTz425usc8o6XuWCr
spLb5fQRPq3JhBZrawNJvCzsYRiK+79zGKXQoVP/17Z+vJ+TNhf/Uo/n4KPS6bfo
1MCJ8oo/a7cSNg3705ovThqrHQsEf70XK3+wIxlKNJVUDONQYpdJ60Ig3hyczyYj
z/WDk8K+Gl85tgRxKykyND7b7/nIYVe/yAaD15D2VrcnOpd3iPksVFKl78g8jVvW
WoGYtgSq2zHfeQPIvYRuEQaxHEIOXArplXNe1c7gjwhjSoRf4LAFkoQISsVXpUyD
tkwjOm2EPriKHLNApN2Nha1xrLxwY7GQnjUmkQBCgZH1fUIkvv5bpTYcED7ulXhU
mQCy8r41lYqyc2lVGafC9TumSJ8iiS3KQX8y+8ti1or2PVcXfTrrqefRKMdNC5V6
U8G920IPOy29KHq2YCwmsHX1moq13gCk4JcRlBtn4qkVSeGwQwQ+LkJmHpwjvfN8
M8xoz19N4Vnhlehp+PLbDfrD/lSStWp4t9ToO9J3RdankgYwkp//6k3iN4HBeL0L
6Sdffvy01j5LFCK2eBhfvb9fU6aIShy27ewcUKPSpFeI3bcbh3iRTRJbinqlD+az
ALxoHiGuWUAxtIa73f4u8H1PLzD1PqTr8EbgpNllkBFjsjKwZGeXAKUxMgKRXCYN
J535EOTF1q8/jPI1fiV9dwkyWTG5IoaaJmNcenVhXR/WEy+mxd49ihZ/Oha8GG5I
G2kFskRhc3AuFqrJRkFD5rz6McjxZNkP1nuGIP+dy0/ke29Ll5y/ja+jfijgh+2b
chiG9UvtZtPb2edx//woX3iUFSPSr6SJQU4B9lUfvTGT3skO07ID0VV07z4oBxWU
UI9La8OKNB5OrX39jV6mCKZkodqBXBxz22iII3c+wzXH5p1/rH9UTGH84s2PCnM6
mbFpPtAw49KhlfdUw4KHvf9TpTdP09Ltopz3DVlX1PSVqg4X4cNwwYgMwFRwWWI7
SSDWg8tdMOmX2dcyWjZ5zEnx86zpzSOorQqYmhOa2029V1E7PeItSFcPR6YlQyMx
e2gF31WZuxM1qXVUC3Sl0dpZXe0CbHMYNaArv2ezap2u4jBlLB97eCZ9aWuYW7ht
xN5zeqVw34W4xK41XWkscIMbVM5krHlO1BoUut0JlzmHSRBSgCSL6VfaLWkUrJta
lyqsK9NoUIFdV+XrPKYKOwYHSpj+E/eBWWExfUP/vCP2UHnhPguf01I4t34G5x6Q
n91jj6rmtVXpAMCImHagauBz8FU+0z8rqnekPDbG4M+G1MIMN6av+YbcxCkKGgI4
8LclnVyxmWnHpulipBLgDvCEoHj0PZqIo4P6muPY1wyXKGNvZg0lV2f0bVVAwhOd
SvAH5MVkf4DZQWW5cGs0Rh3YbWTi2Qr2TJdFh81IiSNbNsswS367QrLtsa5hoVC9
8tYycrqOpFNylEJtOEt3SKGsvBhJAWsqKcsd51yGCCEdZa+BnsTHBMmDjKnxNBSL
0duG637ivP4UdTn2uO8XhemcsvLCicG677+LyLCT61ms4s1h8khtm0GsolQTRbZH
02fTKc2OWiYJWZIVEU+hDLihX74T4GIZvZghkK7kW9+3596VPOWDtFBsyea1epPE
fIl8FWwROOEA0GzWGoTR08p/eC/w2EYeLDKjuj/1jI2i+q/bPuDD2eukRHSAzkW6
UQAFTMaYd/Zzqm6OyX8nlkbfdtN18Tz9C4BIMgnAkonANGDVqAW0NbuQJ+g8KryE
wj4QBhRxhKMB//Gsql0U0Hheso85KjaxilO6rEplxIf79Rd058NPHAM0jb4DIjrm
1Gc9s4a0zhDYz/qWchGZv4Jz/1hqmRIjEFIP05CtAVdB031Pl0sVHbdRRfpT+T7F
ySNkH7gEEKusuFSJzFRqueVTtYFUS9HGc0duaFgCXYx4kfEJp5GNa75MUHEGvtau
CGIGLeDgQGkBZvjl3+Rf20smvK0L4Ty2TqkUhiisxd9nyeXaPhL7qG3WI3Kz3frz
e4FhYWmcTqKXtx08tOIw60rNXQDhvxdvfWw0uU/OYwp0484apYYygx4nPh75QBk2
xOoL9NzIftEBEF9RaawGFnuau2Gpjt4MYjtUAG6g9hYPRPKMalpxau+3/h9XDb9r
Psm1STBkIceuoDpQOh1Y1nrUlRyE7ngCYiqJ215ZQ4HypnzL6a7nru4Wv55LXtwO
LOlmH4SE3oCAvTL1cvhq3Wp1fxaJeRsA35VmmT1O24A2/ivqcYc6KrGwoEdD46Bt
71y5tbFkXKVfqso9OkVOLcbNAwuOVtAilaZYvHCCFWd7zb/E6E2BSzIa7ZXPLQC1
bBhZ4L2qR7os3E9DsW5YE88PzIPF7xtJ+El9yi75hEjQYIzg4ZAo4iC7Ef6rcIt9
dMHNxp+VQAfUBmw/mb3lb7DxigQK1r/9QzlPAvOmOwKMVELzoBgc+UcXIdWgoKZI
c57d5e6WKCYm9IM6R7aDCXM2heQB60YS4JkYdoIEFlSUplLpWG2ejT+EX12POYtB
9iW8ecEB0UXD1P9xYl41AzmOTBxsm2L4bf0bTm/H6lvyXAw6K7/FJNlMW3SiSo0Z
DilDEVh4FaIMn1lQCkdSFPxae1lW3FJ/AFo/9/Vk/H+Vb09GspJHonar2e6mwg9y
gKNd96SRBkvUqQZJNUsLuUOp1/sk+9dLBFLssLwWxA22qwPBEGnwsX3ELm5XVa1y
ga/4VtL8gyg9qw70yzTy3DOFkuoYFPZ5J3ZncrqQhcSqFhwXaMnuReUW5pGPFo7B
3S0JOwKFp17H4JEpjtTmgNszSTEXlH+i9ss8ZQa2F923Wd2iZD6EUGyl5woM+Vls
p6gVdjCo3o2xgEbDQOlzFsmXKa7e/ndTeO7+602LSa/hBvB/YS41ifjCqApxFOv+
jHD8VTz+tvlkGrrw6L8yHF78H+x60O7PzHLy8HUqXSegLx3/PUfeznO+NnzclUrX
pXbzT5YzgtWO0gwbgJ+O5Nj45PrJcuZTc41l599sL8Ei/bAFa3x5h4ycvT3nEClA
1fJgkGUbR6JIz3wj9bZLt+v3Zlu3VFeKQSstuBBld1rqsTdebhexHueNvS/v5fP8
v0k70VH9pwt0KL4GQQAVKdJWrA6VpuXMhcyKdeCUc/C9jrDxXS60zKRPN5pyq8iU
AhFkq2LoHVGNs4Qg6y+5KyQY5t/HBwkF0kKo1b1w+T0w6Xjan+DPV60l/q7+pVKE
nJ/wqyopMxSAKADnaL+csfTgcKcFWEa1DUlVklC/cPXd4pigKL9Oq7pvMXqZbz8o
QBz5HlQQE58bFT2MhcHWqPIT2vF8oiBHqenQ9jn5UosJlfYo//eGjCdQNug7SksR
oRmh+jEehXGNLV/PR3Uo3XUL+rNvEZAtEtPTxXLIkGwpS60lAnRzOy417GDs3VXR
2kGuxda6KFZrFbOktXCcBDIGU/ht6Dy2OX38+VJj1Ph9lg5Y1SIEsF0DEQ95B77P
fkQoJt73vsyUVyx3Ly4x/E7Yql3qzRX99dmimBZErWOhuL+McZ9heJwAqu5iLA8a
zO5eDi3JzgOfcmYHeb+ftkGg6DA7TTghTdVG6KCuns/QITZRG/ifnZTPNy9sVl1s
mJJdKWU37CrrniweMF50DWg4YpiAZuXpRyza+0eR9Q98jT0RRb2dfYIZF0ZlPGYY
0VzZ/ZI3+aqQUSMTHO1aHwi4KlqROYjHQVQhCwunqgCYx7xb09tUnxRxFzMVx8V9
seS9awsubS7WMf8guQhHZQGLKQ/gahbE2mfDUaFB/hZy2W1SZRR94hhU1+CI2Fw2
ePpuqHephiPSXO3bqA+aeegWGL7MNPpFX8/EqP5xNJwODsPD8g1sM+DQn7nZ6s6F
8Izz6c5Y9G7SUBLsfu8kX1TwwbtQxU7q4SV4Yd1X5D6vt7mm4OwimtZliHfdu6hP
NjEZo2CRRaCeAp6ImfzLGUkBgJ0gtIrrVIm7Y3axlbWdsFAwlNPTLs0PKNxciFeM
FLT9/p2FKC9fvhgUok+ktO92qQKkOE7oI6IxF3RVCir1rPY0UHKNYkQvOngApKmf
g+fzVuZAZHfcwZNkYLWXPzwNVUjFBSDEMnNId2Xg5HNeL+boKIOzlw+eJiokFAI3
bg7FGlXlBjZlyNQP98q2+MMpVKkzPdx/j2zmcPpwMsmWms28PjdAic7me5I4zxQc
CpcObPzzqMrGlkS+fNqp7UN+dN/Ih9HoVivObiHFPxvCCeWJW/GSISINZpH93T1n
fGdi18fAkkjPHUnV771RxTuHzPjhhl30zcC4SC22O0m4qFuXOWX/6DfQBiOGBoyh
fOO90q3zHcsVzS3sEHbdqEX+XrlX6tVeJvgNybYy1B08AFZIO4/6FbN5Ll7N2uKP
TnI6oCKvGJwIQm7b1yPPMD+n3Zf73QxBLMllAKUPCUB7m0hkkMxdCBWfG1mr2Its
LwxtmYdd8GBog02rPybNhyYAmIkJiWW43cGOC5ANtBDXcFsHikhz3QwKhXUWkbDi
YqRrD1m2BVpEGN/uIr3qcdaKwa3uIYH8yDPFegxlP9pwcT/CUkzwUbFyRfc3gEEr
2X0AZqBeFrN2pkqZm/LNOIATal9sFIYidfMpdbt8Qj95z4nih1ZEOZK2YfreElio
ELW2e0QwYx76epPA2Y1Vp6QO7KmKNdQ718KVrYQfpiaLK5Kv+10JHl1SsbAGU24P
0jPmlpTdXklxcTfonK62xUfZ/Nd9cwNnYVQBjQ/T0pgq8c1ljjBYMnsIEsyUgtQO
wOBrWWh4huUb5tyKgdSLEPULAodsks8nN8crzuAMXI3ntRUCycYY7jkIUQuzYNIa
GriVXnCGRuInEt8XXqvS3pcxNJ05e0N90NPVsHyu3X+kcTgzGMQf7hHTxlXEhrBK
dmkvW5sqVtfAnV8AHByL1Ju9rYMG08YdZbNy9NxUpDBlQ21xekCCf17CX0cwQCaN
YTiDSYFaw+hCRpHhXyMpGlGntwHzce/bgmAKIVb/0sIleg8Hr53yT3n0SjahiwW4
EuEZkkqix1QT+yh8dVWK/ara34emjP7P8rXdpjBh+UnK2LmcFIeSbP4wn9hcWENi
PENCmy56QLeYNfk0lnAhCIiNLK6FA+BHMhTNW74Ict3okeCwhnFHIWSXKnAWLMCC
sNtRe7XErqgOL5KDVQU5ZreZ57MGW4d3l0uXHOpr5Bu1mWtTGkzM8xX14QnPNVML
rQqLhu+/+PbCV+oZae9hh8dLV/Eu6GQTDeOaenWd6ToLfaMSq96IEMTnuEvI9S2K
uUoEmAo372QO6zIYHTDX35ObMWE4PrHfkmZmG3zKiye7R1CclsCTKk/lzs2KFB+t
+7shR0ZAfvSVz8HMKQTDrjQmJJ1cBDHOKfYtGqwqZiaW3AUZYTibLUFbooPILq7E
8MS5Duc0d9USGBqMXsxOZ5FGSZ7V3mPgFcATu9CqXdzNF3E8f75i7EFAthO0o3G0
uiw80Fhl18OLCVSYAmcPYNgTSEYHL9unkig49lKuji0zt/0e6NmPIi/U0XcO/CQe
YuJSSQt1YzRMT+u+5Lo7KkKTvfyJ7414Sholzt7qIMPjsLFXB+AkXvkKemOump6y
1I+CazTw106zLnu80n3uBrncRUZnzYc62/EYoBN4hUHz2yqZywtHfFpEUXcTk1AP
4/rY++lyImElKc7edst80QPe9JveuEeiN6DndRxgjt5Ks4KfN+M5cgTSHJGpHd7e
AAc2pE3tS/b9RckH9TGRJT4wJpe8f5mZTHt3j2Ihh+p3XCzHVswjexRTaRcdrKAd
Ggxd04InEG9W0WZ9dmg9Pw7X8L9UMETuWSbo3xMtYBAfHFaamXp3zX/TgxbKCaGu
lzqnxEOgWdAwSIzUfJkTKh+tQJLYicL3U085O1I7EPMIk0lxR/Warwd9iDmFDU+l
kghkipGcMGIalTvvEe9Rgp1CtAIMl6afIckk6AdFvIVeVMDn5QrvRC9jPiziEEne
U811wTSkopKEzb8VIZxWh3JQ4YEFp20WyJAEwZolmgDYKXEv0dVQwuWGT7mNonX7
VCloMRm/vScsOj2LLsg5g6T79l3+db9wA1uVSC8rS5A9ObxlXCyOGW378bg7a1S1
ytWOIZmadk9us3SR6ZKjVdDheNFLIl0qur+hYxBCes6joXvVPpeR52EaoRt9T89D
d00jnNku8Wkh6/NAtJ/uVu6JO51+qVaWygYtoBbxYIYs7rr+Pd04TqeajBC0503Y
wTaqPldh6pG39RR2LB85syKyzFXtYTivWwsoHP4LB2d9LX9GbZgr4AxTXvUMo7K3
10rvuSSFg/4SvFltusreNcck17TAG+dEQNL301H1OrGGoQWQmsjPUPN+HzRrTvFK
Aq69Avi7MAQpIU8MsIva0Ql9UM0H5fpfFx0PXAj5J0rP+0GvVasKA64h9caLYEzm
EODHeTEx3iWagxp1R4xful2Sjj52UcjgZhlRrknk2Mu2ACwp3wzYRim1Qp8FPAO4
oeRyomJQcDGkQsgdRNw/ufg8s74QOfdWt6rsmOrR3obm4+ciI9pYEWnY7NL0hTed
5f6Cg4bNEWpXnBB9Lp+q8GwiFJtQm6OU2dWAPZmavFW8l5JqLwiixzX/CB9fC0Ef
AOyNxUywpqiRUXVmxLl6PS0Cn4LKaRuw1xOQAmaKKZ4y4iqjizQ1DzSW1vyAMAUJ
MbjcEIPWn/ZkZkobL5/++4aYOj0WyrLsY+fHr1gfL5wP6LzgXLD340CX8OPcHbVa
E1shhAy+qsDruTnJCxH2bRi/QVeRJXfrk8TOKdbp89c5yk05k9XISa3MFMCK0Dzk
tI0M1tqKQv6RnM7w+NzQuApHqHyLsfQk2uSblOeS5sxZvLkSmEL73viUi91LQtC2
OhiNiJn/foN/FAc06L5ht51JTIp1qkobjBbhyWm7GHj6NfZm/HRHbBEyKGlq1Knc
aDUpPFuia1Ofz5UYI9UOlbcZbtJLIm42Hkrj9Bwmrx2VFJt2nUBk6Su8t+9qXxq+
DTPE/N0FcfixrhjMBn+iSryYWNHa8+z3AkK3a3eS+X9ebeMlFPU/TF6AV1pNbX8+
c7kO1Tx5I/KVQ4MPAc+bT1jCZDs1ztkYbghJGKqcN0YsVvXsCFkXuVKFfVDeoWnJ
X6GhtNvMpibCEOokNPllde6WyVE7mb+W2UNQcAJk/6ABMy5Sie5TXD4xoXuf4kQH
EYO6KyRuLrJd6OZk9cunbnq8OCbjiOx5CdzvqfdY7smjk8MaoVlsS/y5FpWtjVjD
6B1OtwSGD+0sdK15JHZPOEfkzt4zTYHz16uwkB8VSQOwmcT3DHlBDdDuIN9QpXHR
3AVVFv8DRWjkc7N06VT4Bb+lB6iJ9d4Xcx1rHkMx+4JnsYmJmvfqKnGJsX0AFbrS
APMMAfEJ0vTAymBkz0wi8ytyq8x2mJiGDgPKzFPKLq54yj7JGpBt3Lh0jE5MSJ+U
Z9Ba8Jh5Ma7SMWAd8Y7pv6fBsziY3gkUHyqLnAlF2JeIw4inFLRyek5EkI0OEX0S
h7LYCKPxvdo4Wt6hKunLLQx0m9A8Dc4MftHEVOIoKg46W7n8p2T+XvYhgMNBC5+T
Upn8VEZoW/lUxfH4EFtTF+ychWxGFjmsw9O9yona9uAqlf98q9GIX2Uct3nojFww
PnRe2HFFj+YHdP7EU/yyDQy7oKEWbZqjqY0dxRr3vY7acc67HJJzPHztzlJYFje9
8hStsEzGZ4PM7QcAMNtv70jHddEvP6LOo1MRhBN7Bh8ZMqoLr2tf0sxlLh2cIfnN
31Z73Qh81zNAStgZ6WKcWxvo+TZm17QZ/m3Ydgy30ogUbnID2ynm9QWB3PFvApx5
iE27HbbRYwx5X/peFeA6shmsXesgHMOVeEwe3kJHphCoJNHKxycNajKSJ4mdYXIC
kE9BImE3Mepe4b2vSB/3OBL0/eoN7tYx2jigmrtLA3UX7eJHpLwvElkVpCfOOaBq
LBNRNh9/nNS7RqHUuVhtg6wDOQMsAfgy/f7ODjdRJ8ivoSzKXB7IkjfRBSR5i6cK
M8Xay+oOMB4ynaW6fiOzG5U7zseDmFXndYoWfOEDOC956gRH1Z6/DOfajVoZpynt
5k25ggc51p1cMfxvKhdpGVHe5Dnx1xqxseR97YLOBEzjSlStGqWKYEroXYWOMayV
clAXrcfpcdwQsKQDsjkpgL9Rja2OHUCbxKVdr9HynwRdEnn/AInjar5rv8SuUfys
1G8fUTdaRoYLP/jxTRQ21xizUife4oQzLmsg7qn4ByCA4sr+OTfgYEcuPh1JlXZQ
vqppl5YuOvx4wL3vbOBZDt2F/4g6WXlDpPuB7jH/kuXLrlT6wQIpI3JRisbCjEWi
DuPBTASBsm/ZqAhRIUKCp9f8L5QMuZNMk4ZIY6rLiPFGbvcOcn0y85jVc8Ywgi3+
LuI1ktGVAcz5ifDxAyqvPImkq6pQ3ebgm2p4scHDEa/lirvPZof3AkTyvXr6tsUW
n4DgPBeUsByBcyguIMeJNZ4EOoaU/pIsKugMUHP4dVC3y3HYGaBqFfqJu5jIelU5
4Mym3rj6xtPg0h0pJwilkRDN9kRtQE8NSNGDltTyg8bQ/D7wTAg8O1XReVoYIFzy
pZ4sgtW0Zi43DMXq0lDsDAvNjkKolI542av6yiIBA3qw8E3GGcJr3qCk+2WvZkrZ
LC04RFNAYEeNWbQ8bRn0rWiDnbN7trF0vernM/DiZs4gxeJ3ZTV2faCZBWSXN8YY
FvkvXc9GqOq/oMJ9phQMMsNYyd9G6MoYQmlk0Bxj+nD/s51XERJHsxphbO1pV1/N
TBB7F7+vYK+neP/nhtAb7DAkPYujUX9mmui80tFr6zFHS14lYKynhFAcV1rZZekv
yBHmJooQ1XLj0mBgnnx9GJSjWzKpZ50Rz3XnPBXyk/nKCVguZ6A6p+8NNl1PaAqx
6Rd9WJRQGWsh+eGz8lK0EZQ8+8mifn2oB6VnA/jeEyI1KXtYbURxMkJ2cN84KF44
A6rtr6AmLlaOZF0qm4TTVrlBMbMyYa3A9uIfBxMfzJGM6BRJ6S+GYRp50RO9oeS/
uNVTKGgsUymD6rVsuAfwlZ8pGKCZxZWjrJzkDMYq8arMAmkd+Hpm5VZBaA9PKKd7
yJoCSu+J9p92eevs2fqKLHvqqecenQGFxLFRrYD+egJM7MnlC9cndXJJVNMMTJzq
5HUdQYMGmDmt4KW7BRS+WVdHv+T35925IIFaB3tPJ553u2b/2ogy5ed7XJJut5MA
PeY8OyZ3DbpbnHvIgiY5o6BbwuNoJ7Rt7xAbvcluxj77iYEAf7hzmU5bNRTyjivP
WHUEcwCuGXo7nyMmRlIX8dxxvxkTamMb0mOAxH/MQzHdvtVnIv1oLC5i1/lnoFSb
qlAbWFdNMUDLXAiZCOAs/J1OaZUG2du68QUQ9WHt+PSCV49opnx9ltc33y+Zt2q9
tSa11r6tK2e0B93SzA66dO/uMgIRcr3Ge7kNKPBQC5BsbTEaroQ1mgeV9jdy3h1l
epZAqdIe18xzKAKiHzoe7jgQOvAJ/mMNogdu/+szh921CzsMqNQ/DYC4wYctY7ur
HY++zKgxvWLyyhuofBPAqBwfLOaAsuH8uKLCl0YZmknnAyiL3/mLRQZVDJVZunUC
YyOBeElroCSP+F0jZt5VfBu+0WmuIkiQpqe1qEr+oh5u6zTsow3e5bdjZYO4OtIC
hdbXeg8/8qP+NW/I90e1ARAitKDNAh6d7ks6d9+OBbl3P5i+b5UycYaWPX+ekqGe
P6yP4uR1SwTBhlG1ZnPVqSktAHKJrLKl/s1hzPJxea9CfdmXIqmHS3YHzhDHxCnB
/aO3TQPJ3vnuMGEXlNm9Ix7oqSZ7XhNxd9fuFVjXUS0ulrqMJR/rAotKH1+wJmxX
53m0/K9GDVSGADSjNWFcwXGaBkImKfmWqk43TA9s50lWodCyUGlqWzMj7VJrEQmx
rbQOXLIzUyXfKQJxypNxcz9KHHeD30Zf+CtvkA7/q4iOGgjAR+cYZeiNYkmiWclQ
0ZMXJBA2PXxxkRD6GhXYe1+nB8Q7Q2ew1SYtyrPnEexrijKuSSO03HsNNmNqA21X
SAteBJ5K6fzOh66AG0VDkgpN8pq55EYctGO/f8VuMEopDPCil/1MqkiBJ9GbG5Kj
SKXZIa04ofAMAuf7PmylG6DCUVvIHCKMOHmglhi2b3nutyvho6PpQgBrLrjAgN2O
mmh6GUHmPO7ib7xU8kcuHHRcQ+BJcYR56Gzt1di3Gi41avNS1WjHesO7qjzbzk7G
atyXu9IILM6cAMksQzjf+mOJPyKOepvq/hXT/Jv6jIGMpZ8WCu4zuSQcICbtHj9o
lhuuJBmIFY2UMzVXkGIPERxLPUUFumW7I59dmEsXi7qj3BDvqjCV7r0wj2r/FsVA
eWh2pFS0/i56okYiJcU7uAWh4XAT/MH1Hw3lAJjSUIR/slQiaXxf7sQ1AVYCSogP
0FNrL0aTWZ+fjiP0aKBQvfnfD/X84lzrJt3Wvts1ycIRQ4LGEoJMK4737zG5a+Wa
VkOrpF86l8FIOhBTje0dC/SFtRMx0TnHbCoqwid9RuoVweVUXu1RC/GAaY+K6msH
xTio9/UBJcn+8dcsdeecgFZ1U3CU7/Spe6ICE7z5b2kZNuVi75pM8HPiTvxNZA2p
no0X//r5jryRxBjBDnrbXp//jZGROQ8kZTJO/X8e+aFABZeEI6W6vJ5hyauS4POy
Cd74+Hx5N0EgsIcVsu3SJH4c936pL20O1+I+y26JPhFNfKD+QzdL6XJhy/7dTN+y
xtanE61K2s/sMKzmz7X0QqJfNsaXtMRZ+KU/LRbT0KfDOW7sRHC9ljChoGNp2ZOf
rOvfHZYZbiquNs3hb/wolMSSSeB5hOAu/aT6oGIsYOYDSXC34rAX50RdkoNIzjfm
K1irGzWPGjdjjjivy3qABxrrJPy1WxIzKWSfK5cRV/tJ/ljsFTPJyKJxJBNf8emi
9FoYAE5dijE3TAWHc/j43VTqG5Y62V9AcIIFldzosgYIWHRALnZvJxfwgIRKU4HE
01c2orFqv4qNvXyu/SYUxmrjLTmjtI6EEOew3FJGS/c8zzlec6snyv1ouqsjnZ5V
g8oxTEI4Z6mTPhunS7HxK3AIJjgQXueQyXakgsffE87fp+HTdx4z7ouIivCNLhkb
qDk4nq2gy+GZ5+StnPMFOrszGCQLExLl/SGN0utId2XxDfWYTPgXYwgAF427JgO5
GeZAYqESDX4p3SOPphi+eSIlOEBJUcPFsQvw6rF+naKL8I7KsJU11m6DTvbbw/11
7xQ/q9zmv0QYo2HO+RYdo4vtGKyQN0iVWh5GcAzhdOJ6K44BEQh6EhLKvTgPoxeW
o8W1oFoAqxR+Nu8unseteDfTf8RmdrvrOqNvFDS/Q2zwvPsyukUGdv7VTvc/twOq
3GvmUA+036Ovh5zf8FEhQllSWThEl5kjONuIa6oePu9YOg64tKHlc+Gj6WGO54/g
MhJkj9idvxdHvCbBdePzWS9qwZgWJS1O5UrHtDIH3GEoCVV+BT9vr4WxMhmPR2hq
VvPp6Eo9feC07sZ947w0CsPRsiqX6iq9FKcF0W4aXs/7RdgcFYbx6n3K5KgnUuBh
RKvHGwHzdDTY63KwWBfUDjq141zJVU/is6q+ozmoIVelBoqDM7mFFXnWs6btxonA
caqxrxTw6UxJqHGEiyVcCm6KtYFQP6ZVFqoRVV0aj1pbYKjCe3wdgLevb7ECq2Nm
Elei5FQYXgvXsD6+dc5V+DmpoDQ49742iCjOLQ5ZaF835UF1WiSdLw9tbOfN6q5v
93Yzh1R0s37GdLj5xGAj816I7Quiilu7rS+IZRsHdlHyDb+s1N4koQa7BGiqe4zw
WzmfcBlzUqK0wfbxcrVRXT6oVWz5YtmyhFLASb/leGCtVA0a0J4cQN/EAbJanBvf
MlghI8tOwBUDXYh7grpfoZm+7sbQ+hMUZx+BIV+LoXZBRadj4cJS1n0c+kt3x1tx
W7lctc7amfJHHJ2Kb3vJ5fRPnP6JVZKtT6aRKn6ZJLI04+rp1Np/nPIUYl1Do+sH
pgGC+/mK6fuOKgox5sQwgE6sUgyNoFQrnaJ5Ipek3ErGX4zYEg/uFjYa/EN1CZLB
Y+jf2grUzIHiXNzniYtA9260NrFtnExjUUSIbMZlU3xu8LuDEQpsq9QK40o28y9H
bDieIo5p+vDNcbJ2UgwmQZzhLPl+9Lcqke4DqKm/O2vcUoEwHMi3RWOJkbe9iEnY
6LutsCXb6AgTlwRfOwnjoKxXsjYKj5VZAGUO8PWagM+61646mjtGgFOTrB7Ob8ew
/i7aBNkSKszHbliCoFWiyiuPHGtZPIut90yAyvR1fHddpDWf/jY22Ag9PaD/aTq3
+zwlSr9FSZM4PvaS1AyaJc5Uubx0LKi55iSyrGDtCeL6ftuwGx/brhqt+6ncruEE
Ouq03DdabBdAztqqWCCX+PHruJI0kd0f99cEHR6RvHs+FqGUXCkveJ+EwQkcKRlX
/PIwVCuo1GlOfJ0RFViCYz0i0kdt2JYaE3R4FeoXU77Uty6a1p7wi+DcV1QkePNc
Xqy5LtiXBH8o3FkQyT9qojQvjS5SD5fYS1ybOUDohxq32HUNedWGf/gmqDnlf5+5
OlwCxDRoACEgv46J8gNQuaQ5KGxr092dFBoUXCnfp/HRfMBhTsCldHA0giqfF9uZ
1AhuyY+yyA7Jo+c43qf/C6+tVac5tG7EM5GDDFljwibkL6kkWVaJNn19jIK0cgof
DcAVJ0zMMHIWIi0IMUGMH9YODrG40R6DNdO65WoWMj1NVZ3qxhZRZZqOO2pGGrMI
N/lTesLmhvtiC89nQQmOAyCsw4rla6NYdYZu82qSKqGsGN9rthMjR6WT0kf2Uo1B
YlESKEuHu8ZXsUoHdiUkBvsZoobsjGBfgupVYAsHsTqe1UYtL+N/jA1V7dDpgwB6
+t44tM4a2JYjjdJCnoC/vL00e7Ite8L+dKVum3AErPkEHCneJ/s3JErZQW1+gOPT
u1CgN69A0vYVZHfG2sCR83DrUwlZp13RajHSpkna2egTKiC1UjOdlvKjtt7pVg8h
wG4Ll0ULpcH1CZiZz0Z4ahbOJupJvrdncmiyQbWo4ChkuijUOt2U4gvUgwgBnuVx
DS9D5AtNm0yKyhIa/hJf+6LSTm03cu0c/uHrQG1o7SQQWrshigN4v/Uz1c0dmOWQ
lptjaQSB6iTTbddvCr4u7FO560xPMhOs52TBJXIhLy7hcRWfMs5ehjZHMXAadHqR
pCAVG+7s9SW9DIMhXi/zjeUk/y8WkJ+9wntO4Xit49m0qQEfC8PhhzjjlR24cFOn
tNvyfbDCgj4zf0GroUcVXuImaew1P/AIcWVoIKz8iNyjDGft4YluwjDqQ7rCD0TJ
4cOg/KEJM372hJcsK5+R+lSWeXrqApFo7AVyKlPfRV1bdwiIXNRrpAvtbEG4j37g
p6bfb165xOrBbfpQ+OJtGU7upRFBChazUqiENJZBHKWN0Lty94IfseOL94H05GQ1
7Ek/hUu56DIv+mhZm+wFT3cP4Zi5i53cfmcpHAbCHnXx2AOvshGoHxr05G1E9tDr
VFjqwbjLHr1g+c38SHKTQ11oHstcQ0uUbQHfzQfNlqpTKVZQPLaMtjJHqHJhDNWJ
VXkiLzDz5rapXlPv/2tSdnKR4ps6Q/fCtXQ3Q/lN0Q7bQ2sQeWOFKgvzJfm98kI/
prH99fk5s2fMq3TKnk0FXCd1srVkPF9jvWSd2NmISGvDKme8s/awwL4iHoAfuQi+
cBVgGLQcqh0QaHd0lxj3j6gvNXv15maqdIuckwTS3fZ0LHJ5YHJoKlD/rBKUYgzE
QtytmEWetWyk9eVtY4PYEknSPvLD3A/U29HNx35TUVWuikr0GEQfy6Aj0RECM4we
9ZU4g+xKFaMxny6iaAx0ajhsXfRWFGdlNWlu+Hd9z/C7gc87rd5AVLXb79NvfhG5
s+rGn50VsXigtwatKyuZz+dlMoIy7FDyklhtHJdtFQLfLLq+Ongfd4yHw9fq8ioQ
84tVlJUqq1/lViffj/GY8tB1m6LoCB+sRwwOyGI05R8YpPU71U2yx3LYLdwyzce5
nOnU2n4/XZVaXffnRs0QC/cdLZjH3N5hO6bdmMJb0qtyIi7iX3WcsCii+TLzedIy
f1mD1O9TrMnNCeuUuKd2YC2clxOLYzgRvmqlxouAnPhfdYTw9skb5OXhF1ptY5SF
UlKXL7Zyg3I43MmfO/WNIYstWVvbHkWw9TcrHgXoaBzmmNuN2B2jKcmUHVpzSxyw
JWJHvS3XnLxTp7J/gl56mlXi2iL0AiYWSS42e2NLNpSH+zKOEhz7+ELFJLnl1lF6
twaoz8ChcIgfTmrUATj2q8KWhUMMscY45rHWzDeJPpHQpA2+xhhtEVqvDZNV5GWZ
BIeFBkx4KUVFeroojR9w2iblQyyNRVxs+JHkwGHqQLohFy9hU+eUc5dnw4qc3fSb
MQ/WbAFaSBrNzVjMH/KIykE2wzGmlz7tbYGhYL89tfiatHzqw4WA6mpPSwQHhwsy
D1x68bJ5XjmosoHcN81sZ7+EGlbLREPeYRcVXEDD6CrjS6ae7H/tpgAcJ+UcOvve
ibh8KOjNwd5B1/4pDkcHporYtVcIiE8xhrXXPN3xu5v7Pui+dqLSbYGn4afDxd4k
4TPTvaOffXHLSVX0foP80eZYvrFEN/I3H1/YaMaecc9iO7vqFdlCgPx4WoezkW0X
ZRwEPB6h6eztXJX88JLph3ETuTDxbK8zEjESRsSag1wXHhjkVMkrtT8KehVqcBb1
uTMPLgfHdyrQbPvyJ18dIF5VwcRUtHqv7qa9S0wDrRp+mHJLp3Cs5A5YX6NaBi/u
jCgwDmt2O6rpLkj0nnQYVlU2uK8//ljqMhrgfQBSwqHuNFEWenZxz0PDFWMCoUaD
JCPycVQHYBVcukBx6gJ6JfvoaKGcSbPVHOmWyuKGUHuvi9FCE+d1CFqYFIo1Lk1b
GWYZd4a93fDEmNWGsg3yWMcmwT9T1aJfjeYfUWnxCZylOSlovFUMF02MBFQjgxb4
0tSE6uemTSHbJ+7z2CWqbW6xJ/7mtZVUuGJBfw1WT7I/slsGlbUxA7WBrmkvVKtq
rr+hwgLnqDHwgOpjz/zK3HQpeOhuovNS+pGjFPAjmPiS8rZ0+qs460dNryPY/STR
l8qgqokUaiidID3q7kbm27LiHkNWDsFZ9UMaE1nKGVDLVzPaBAU9+gh7vl3yjY4N
2zN0NcJa8zY3fAkl92CVTovJKkApINPm4GqDAU/26JNNrz0AFbtt7j7poyXqfmq2
XSRq8g3jX/20y3AaynuHZruvHB4XM5rVvfpGVm+6PVG6gUiFB4HdUOvgplzVqyVT
VyD18kbm26OYG8Y37PoY20HlJH0fqy80VQ7QNNhha+1He1nBf/i5aMxuyTQNkye1
EU5bVaG3cEq0+o9/a/sR42q/yw8wPbD6pr8cN371D8mHlzm4j3ZDIm++3fyaeu51
amQPL1k2qEfVF3/RQmIvfwht9xU0JzfJsbqLFPGw1dDf8TrseP4aqTb5gnlbLgoU
VIvcIfTy7AYYg/H5iYrwgrKynBOs/lEhSuuou0HkJR1ySFdTc+bvOFICYb9cdP0B
//gLglqBDzlsFkSE9PBGZVOcOJbqtN2puM8wfit6SsXPP3E77fJ61Q6l/VJvoIhI
h+nPQi72SHqZT+cR1iFlQvdhw039OenrNbAZayyQ+xDcKqjQDRGYPrnL3uwFvIGs
WA2YkPmutBOQ9rVBJfbcIRQXdlD2Aw6CHRlYUgt/wlLbwb+6DtnlL4RHt2MZdTOl
BqaopxFXbQ1YqQsUKqVxZED3rFkMG3cxiANI4xFnHDclgONKPBLsdSh1DH8lSR8B
9pP/wcIk85UGuzRoRrTps30BR5b+zoqMsYTFzuBkO2Zbd2qlH6wczXGcngWf+1nu
VmIT5TRk74SODeFaccO8gwp+4z7U5hI0cdRVgzsg8CXuZl3nOwzDVEzfx9svdkcP
8dqF356ZCly+cRFMzWSmZW3xEZRp6cY40F/G1zoRyc/i3BQ3/kLiGAGUTMrVIsGx
nq4qFG+GQFj4v3wBmCVp7ngx2DaPG2vXyWwVq9P6OQyv1M9rpiwYoYw2I/uPyLHy
AKmsZhh1IMp9mk2DnFV1BUk/+zRGU1mOjqVsW/WM2wDSNuUfXRne1D0CS+yuL1Bt
jJhjVFqAKse+/ErWINJahI7FHcu1TSzRlLKxBvmPvLQb+0TMwhAQaYfHEz59OtUn
aC0ElTcltpRl4DaSMz9j+qE+dLWerxaZPx08Bhczr7LwzvoWv7R+R3XgOGfDHKCt
AqyXQDHWJu4j2KdBPJ4992T3zsNiFe4forvAZlHMaqiUcYFKSl92Ph79aV1tks/C
WY9U8JSikchldhfl1k5H4swTHS2iRLmZ+XcFf9KmMClEIw7DnECGdE1eiqIVa/Pl
nBOF2EtQo+7gDRLQ8dTIvDDLVOXGihFEys8qGq6OZHqS2qUpdM9AQXjgRszlLjQL
/ssq++ChHNyQ1Tx5xc6yNbqXXgoCzJhXl0QZ7A97retrK8VWz/hzjPm5BOwvODIx
2rKP/9kMlnSsUU47QRSBDXAktjvrL+FWaphH77Atn4zD+vNaWQFo1QKC2W6kNzWv
jw4rYSt7Fo0s6Uy1mNihqxGuHhprTMFxPB7kV4gYHRin1eKH6O0r6b5+xYezt9Qa
46Cog4oAU6MKPPoYoLhHHI51jC/ZL2QkueULmBU5IIolVbH17Y0c4eCq1jo30YD0
+pVwfoVcK12zfmmCE4Cbq27f9CJkXR8gHO9TmsuA7OEOjfCilDwyu3Qt7QjQGdGK
/0pP3YW2ov8ilSDeMsdonp7TJSX1GRTNZe/850/d6dsGh+4m641VvE6IZrJnYx+k
jt9+hEufSaokECZipvIWOB/oB/s1+7EbHhPWc/NtGj86aN5KhtJJCuNivdUQ46xH
NnpGAZdmcV84sFFv2bFj1/lq/QIt/nY90+G7bYx+O4wNzzumNbX212dQ0fMueSNw
rKGldjduOydO0ALrqGfzVoLOs5BzzLGv7ZMMMJdRtpWGkeHIBjuUDBlb9YKbyig5
LQRbJwCGSv6PMBghVgcwq5RAOGMEgrpXo050wq8Yy7BOymSJBemZo8aRvffIKtjQ
MPmGBdtC9onCfWa/IBJwe6tqFzv/PyqIhj2YNYkAWiVDBfiCwUAcex0yIrJj5NTw
dU9WuL9CI8kkpSyLmhmrYC1ULPdkC4UlNm2kS4JAeE2H0RvTA7u40Mr7ZcPuPNtS
3GMrwTZxFFwv24ZmHeGwwUsY6R1EvF8E0Nbm/U57YRTcNHWE/MqmKGLT7Lp2MHG1
SDaTj3F5jVTamonPWqOmdnfMBy6sqnmPGJCOb5fVA+7vNplLS12hOQ1Zc2ibd0Rw
UOeeH2cKeH6xCv5s0PecYNf375t5F7Php4GOux4AJ1Vjp9Xkj3ZRNpnjSW0cGe3H
m7gLgnqvB6K9CJbJU5nwMJGLRe093JEjgSwIC5zGJclH7sfK21IbFqDwB6xe3EpD
m118EV0Lj1WAR9oLPizHMci1O82W4o4oGgLJNni3mEwhEYeBWlHiL2XUXC25WUWf
F58MaRIRCV9OQBXFEGWErLrMJwERapFS7eIpN0pvrHF9hw24k+XHNakKrT5+gZ9v
j/Yh5AsT+0k8Df5WUFpz1Mry8esUOlPwdm70gIcuE4ct0nn47BvUNzckMW0eHTqr
5xpa+jppDBSpmTQ3SR3wgsTqz1sGqpda59eCgJKH5iDccTxX3K8ji3ddXo2wozaz
bDUQy4QuBwDTCYkt5HGJ487+GHIB8Obz7lSOQ0P3mZZG/LoUbw07uiElAHRK3D7W
L/Rjh92b8AGbRyVeW9Mex9JLAa165W6RTBaAnu1gCq/efuNSY3bYF3OpKrVT/Nr6
qzhk514y1BMNwwDDElMdPIIxNhbZpL0OJ3xM3D8//uIXBJO2mx4QAKh6n45X62/2
8ik/TP8eYTHKPom3YN2xs4xwJyJq/xqAWT4tQA72/ob5QNVP5ltBf+nxGIKKR2Xr
TSv+U8SpKViStPfHyHNJo2dbiPaNFOu3Eq2zxvGIRpDjcPoJNXmkU5uaqKJWnYeo
AvcP6jDKZL6nIoP88jHMEH473zhoFrIvKDvKpKq07lRd3byBLAbbXQFBRNhLisB7
Kg5dv12zz6278zuTvHL9XRY567kEqFd/rrIBGDe9g1GeOTO5TWVVwY8zdno5rNJv
Q85yel/qioihNO8WjmFYCAf3YeKKCGfksAdDludepZQS2LuGc4jIeyeJT8Sdudwo
CoF6+THIZwWP2goq5WqsSAnwIye8RS6eL0FPcsnzivJm1eJky1SJN9Bo98BGtapF
83H7HN1ebu9A9xsNV2SpMJ+r63KCpnJANsJtl8C2wc78ui4RQINyX7WgXVuB6zAx
1EVf3bij0h9EkQXOEFp1DteFA50YfoPDZ+I8DmbDIabw4LXdppfaZSKQP24YR1l4
shyxNXK0Ayc+KM0PSkqvYT5u3DmSdt4KGaOAgzsa4gQCi7dDFJG3ErNcjnSuvZfg
zhdJ35xng301iCerQGUw9oNNiYWr2uqkbi5vroqS2R41aKsdraPaTH0RaIlvzcND
T58EGjxdjZoiBRoCbARUD0vmG5HhGrbvV1tzrbU6diKc2qsDECWDhefV2/NifcA3
UVnjKrJ8Rl+cxuHSM5R59vGAi5RTbzoKCjTNVQOg9cS1Jc8ZJviuPSqUJEf+AJe7
Li1XAjdNsrtkP6JNQOa7OcTS+ie9C1GTYEjR4MxYgMwaT+XrNo7JA5rjfKrrCc68
bfGHYq7hFRVioPAsxVC6zPdJZKven8E8xeScxFYhI/3MbOr/0PTYYu4/fyy7n6Ha
h2dHWJpxAEM1ZeSXS8BxYlF6t5mJp1Sj8+NKvPn/s3PROBADfaedIqXDJG07pian
O0AVVUiNxzI/quhgv6OP9X2QwuL0Jg+dKhZbebC20Wq9uSVi3bjrcd0S6ii5Iz7P
szXWnkt0y+q17El3qgXCzkx0VltIgJTxjp1iDV1dUTNx7nY5/SeTyylhjlwCSh1S
fzYPGlP/Ct/5ADYSFImNcuMn+D/yqUE9N8NI23rDyGUIcKjwLzzpDxAK4OopzQgE
2eKurxMEeGauNmasCaGTpRUhGUjmofBIJW3fwmu5yIGsqJFOAW8q0yUYNJjfXryb
xL+8cZVISTPRrgj0X7RvIO/74g+dsAe+jpA/q0QcaB0D3Zzg8uBlK/4M16kOTzYl
pe4UT9qYpQJVqTVJnAoN+yUj59eR3JjY9NOosEFS/VJTI/03bAEPCNaBXIqxKd7k
9iAiZIB9VHGkCGSUWsWvgyLfwGDHpqHiBurUXj7iuYISY9wnYudlilzdA9yWOY9A
XJmKWD11nt1Dx8UNYO4uVILDfFgevUf9AQPLseZEptH9SC6gxGIGHtM29qVcHNl2
Hz2y43FFqrNEayTuxAOO03awGUHBfF+USu69gh7LVe8+EXQ/mtVizLNIvwcNbkKL
sNGMa3qQ5AGR6VW2Axxe2ETzHm5mKV6pp3cMiPTlnqPPDn9+p2HRXGhkiZmcd7IG
B7MwXHmHaxpq0a4HEMCAA6E6scKo2yi87MN1VwTPR/v84K87AlNDPSKDLvaf2+Za
JltZuQLT7U5ehrklpj7mR58+Amqp0zviIV03x3DW3v0StUmcfid1G+y7b4SK/eUp
R8ZxaToYH3MIOuG/1a5GLTS/+bHXXtLCMcIUO752pTysVbcVT7EIf9gkTsT/RnZR
4ICr5HJzqEsPEx7GjlO0OQNfFV+Omol3pR4D+nN1CwHUANg+EXcwu21MoymPLMmD
cF5xNLmtdlMcZD9F9iFx/Erj2JkbfwOloWcbXde//LfcGsqdAjc2WljHJ9O1r6gR
Oc07py0dLlsswh2QowezmQYp0YNVqycbXazdz3k5MESp9mIMVXTcYEjVDH0qCH0f
yceTMu7Yo9sJLX5+9RpHO8or1V3m9tubQcNjy1L0m2yH1oF5nsILTFBkb1VP2se/
WBkL8XlexDThoTFqhTsURx/cAuzPSR2s1f+zXWAlgaBlV0p8b1wiN3y3aRk0rU/n
y9yG07dXisJFwUwvYBgHDDWJvrOEyCHn5HRNT/tvrbwdFybz/VHJL5+5tZHoQNYC
sMx011EHaOGHff6yXnO8V5Ba8sWIY2I1qPXXDcNUKvScFWlJrYiBpt1VJMz6hZ1o
sNWOpm47QMGa0r4EoL64FM3qjX7jGQkMzWq/xiU6jRgA0gFlKVQXRyF1podBpwtN
F0SA4Ii8RfvfQrI9LJT28azNg+86jXuW+i+sn6ark2WcSTOMHhMX4dsuBKruHgfQ
XtcKTrbPoFGcsJK5eBeIwfYqole/rn7KqWJO8lOVhHWSsOqz2AkAWexXNR1ijO/H
7PuqyCKj9P/L+uzxitZLubUinJdfXinwjzHX5CYZO1e8gyRSrlFaY8s0F8Yg2Hv+
MC4WmV9UNJkuSmDoKsfXAuE7D+JN3MJUqqG3oUiO9ERLnCa3hLdjOp4mrRxcNkbm
Vcx6WYmdxK+IVpkAwQh2VKYABw5q0qEWSMhgDzF9EqGC6gobFLLlWKGSq6TcJuVK
RzRulA4qtGFos9GbojtH8oNGJ7OqRxPR/g0rhavkVR/MqoKztHdSvZxXjkMZUVh1
1H0vLj3inCDdai34gWY3/pZ6JyvuqlScCpHoxRurtS+RwhxIOjt2bEcQKLyXAfwf
1cZRR0Si1HKL95oYNu9Tv6dx+zMh3RDtipaLhYM+tqFtiV7EPS9ZwtBjip6ao7dT
/OkiSJWlif68ShSdcTLMGa03QmDwX+sND0FqImftbFn0VIpMYVOprf92H2gofWgq
OOJ4C6krxzTurpOET7BRx6kycHJ30Cmgitiq5Pq01GBE3O6anQEfbHF4t7YeCEMw
d0gCTbs8zUMimXaQHvlrDLZi1Q0AwNdSSMhg0WYUM1uy19qYh1pyTSqwDx8VrTgi
cFsBN7GoSMwjbs6MhIUPhtUPDFYZMsFxLbetnghw0LQbG4ifxezTJ0QOIfme0mgS
TKO2XDjwJbCV7B3L8y2Wcj5IkC2tLiBUMkNcAnbGVpO6MLoAESambbu7a43KsHO9
IUKQxeLfWwQVUqyBuEU99pdtYJ/AkxheViRPqXC6XOw0oyTdAUhnhYCqWTF5x8oY
64OWmRZWKqmvc2iecydl7DfwAvXYv7hMHgZVsyOwcM7koZDIAxz6QRh7grGf6FRh
G+peFe5MwIEeUBrUVJN/MmQY/8U0ySCuGn2MMGPo/irexsQVqs9kcpCIx//n5NXy
+KFD1GYDgQiKGMHqZeusBh3bk/5sZUfEEcMFYxvJ7OKHSbu/plDPCcT7GRKmt0NM
yvee3Yh70eMSMO28TUdIb/VPyPTIePM7XchVymFZnPrXH4hLtJSquHpCazryzFvc
rVc7WxmamAKRous6L5P3Y7qrUOCw21iPwX3PpxCMGTkcCJo+7Eb6G7mS1p97oRc0
IzRLkbUUvjYIF6qcWjTyd38gndrWhocnSh0VHhnqSdsT7JrNBsxbBarTJMA4oQ+5
SFFW5ZlMh9Hag/84xhFB5JTu5Tay0Fg8QPOZvCGCLaVrPDxOXIogvM3O8x+sQvyl
oNiEqB2r6r1qbzmxqsxjeIRq0KaQqIx3ZJTAUoozjvb/UkmgOC1K41381IwscYjH
HirCWbrynAF41U1Zay1MxVn4FFRdJgl1tSFYBiT8TwA3BPec5/kCJktt2W5Ip8M9
+c6OD5rfpLoRCsipDo/cq9QUaYhE5GhPAMo95VtNclnFwoMFBMqAZ6XPA8hdpLe9
mvr76ci3lYt2zNzkc9orlAutUc6mNPE1AthgVO/TwBsceQBaspkfw/S79JMbYprH
vsr31tYE+R9XvqHvlS40X2Qz8oXVglrDmuv1iz0RQSqKkk5i7ZNY7u2lDUW+Bum1
TitLZuSMe+zDR0ACgDznpu+Umzl2e8X6My2UnLKgP3VGf5GIzaBk3HUt0Ks/MoJK
l06lL1RVCHbV+yxahZPdrqJ4pisa9FVSx81WFjQeNgBRAe0tjjL9nPa9T19DdPJf
jV/30WIi9WJ4HkO5pBuJRPL38RI2jrAsMO9ZwDvZU1R99N7+h/e+p9hn1ECRHxIN
Csp8hY5/fnrej37m0Vb5kjoL0WJDJOvvFfUiXNPUcvO5KSU6tsz1MM4QeURYIC78
ENlitMOYb0B/stTymT5B/oVxyFu/gX5DWNKai5xnAPaVRNV2eoRqbFxtyuoBHRSa
mNJveBWVksjKXFiRq8ib6mn6d41ZZwtc8+jEZFYq9fdv154UAwrcxwpFBlm6p46R
cEh8n/PY/9wN2XBUdVflp+9Y7PlzGE7IW4uDXGN2w29Og0fW0AfjaWQAB9lVhasO
N+Him1O4QGGnSpkG21HiLy71gMjcg5J4vRgdHnFDwerlXSJ7LvS/5sZk/EeRuKn1
Z+H0KnHDhEybKx4p9UQioP4VCB4os/EQaKgxD7XlQwLr3Be3CKXES6pwoBiAVPgO
t8Rg0dALlcZFPvUsWq6zgbZY1HbUfwKBDkioCzmVV3c57P4Z0M3Yt+pE+aVZ82xP
QEbT4z4O4RC5Uh0o/dJ/PZvYr1LsNFHGh4FfO5BJePkRP2qkpblEB0eQqo1KgQi9
oGZRSqMpfjRj8m1s2K/ai+VD25d2Yp+z1eHliImC/GmIfNeTlSMlgaiCZONaS3Fc
ijR6zo5T7i2o4KsJgfyMmQMt+B/Nh2gjLPacrWpz4tJpY2qYaOouoC2nTEKbsfGF
7lqpKafTF53CRNpt4KUYBpIb2KNiDooxBTXyqYCqZhOw5+GdxbWaneKN6EKoQdKA
xprkP5AStWK/xsvjyLJ13lgRL3fmblh0zLpBrM3mGRzJL2ge+qwYDqmZ/cZY3vL0
67GrcchKEDg87QasDxIOE5o79zrSr2pmwWJfX4wAXCSN/v6JwVUoFuglQwsmUs+v
UxDzn7FD4DXLBtm1kQ3qHKJu0miFkZEmyhM8BCf0qjSOEge0/KWZfV+FR8rEW4uB
zg0HI5r1PSfVfXcvIW9a6Wbh18bdiJdS8uxh6LcbLIZOnnf8gsXU7znr+M64UncQ
Fqhfz4+QGO4d2IieXO72GviHxpFwV2NQnyVAiOQcxRmEac5rT4U20pPM7Tb8ENdV
zFu3qLM+dewp8mTFP1wE7gq3vCPGqLz4ak2wdGYY9BUlIBOhg1TgJf7eY104SD6Z
+G8a9qIvpX+0jm+daj/t9vx0QgeA/hQ91QFItZcZ9Tj3rdts46ECTh1wFZCIUNkB
bow3NkqPnWBraBZG7d854XYUd2hOJ02OjevSCPdf/nINuUQHPlE/2Yn1mFjfJFZx
bD2X2mMPJUmek8Uh594CK4YthnClgyrdQA4D2jMp7c5BwLvfJ0Y4Y0oKnc/wFNbZ
g/sH2FGRfEZZB3yA08HXHjmIu8m9VZx5bdcDy0e9jfyjvyrK6iT5Lstt/NofcyEk
DwC7xHfhthfrIoig9p3mDjD2HKQ50PW/d1gz4C3txyq3ZyULpjTStY3u9kQ9sFXH
868ICTinKyAH9kj1ecmzN8e6Zy1u78ngSfHU2eFq+RNPO8EwPK9nLNoqGuNKlP/x
SYgDps+IQqrpuHaNvSgAsfdSnyYPN5BNp5EQiVJrWECdJwJnXEe4vu8Hfc4QK3Uc
CUi/RgpAQ66XzNOXDXROcwjledaCBTkOZTmUoVOYbhEfm1dH2pDp/8G8gk+XoT8b
bCt0igVEErO8E2Qf651IiXrvANxnVx0SwuZit3tjxIWuwzL53G3jdtp3xtDFmWse
TbMYADx1HU//2FyHOVUb49WN8Z9P9yvtRJZ30RjMzbh78bBg/mV6LCVH+z6SdLk1
+F4a7GZR+/D5ThqHg2FMzJmlMgvk7nkQwNbBTF8gvRRuI3FHZ3c8lq2ut1LDKYeQ
Enk4AjqlJ3WufnDpWdy1JGxartXy1ssX+lx9geEDU/HDPLSWPi6TvsRvu/2jBg5V
xM+06aTXNoa1GfpcGI7SUVHDTM8iDmyDSgyq+lsUVGD+8LwNxmaY4dmKZYZCV/My
XuR/3QWp3gc7NL5LyS028z90S7zODf61p2rRAJKKqM0guisRAwNii0CLYytOUXZ8
AhxtHmjmCnyJHFqMiOdIXuwFvUZwDgBKy3B8WkzEaFJN2OfIww+GNDLor2mlZd+f
hEFmo+seLA5IDYu1epy7+KvOa9uJ/7JiY2feK05bMxXUhHDkiarK+GJKukK1TeR7
6DGwvXouiDRM38wFkxBLhqatkbPcp1Y1pygfyd+Fc+fklswSw8D1dONyXjkLfWJ8
waIVmkp0I6CKEH5zhF5uZgIH0NDBs29t3LNxAlky4Sp+YM2/ih2Pzu9lyHbnXT0B
drDZOaGxv1QuG3Fk8n4M2pUlyaE5ZNuwnRgKID5zL8QKT8apqh4W7nMv5ReSQmAi
sXScmlfwE6bxzQTwPsTGZHfq3Yq8n1eSt21rl30P5UZmNA1O80/UjMcYBrkGf+Jk
jGIDUTX5Cs2H4TK2YEdfi65PfvScVAH3O+dizt9xFLnMvMQY/EehQSUAQRgIyW68
2iYkAQke5aTHNyJHDYC0CoF2EvGDmeHsgorvKEPYTIF/3r55AfhMjeA+7yx0y1rT
Iu2tTRxauELwa6EwE3fZ0dV4Tmkk0C4rdL+ty+OWSuxli3Wgdjja7FuSleyxSCu0
KKkZepssyrw/I26bNML5F7cJkq2ofgzcf7jJ6Gp3cUp/hxr7a7FPDqvGdvHq7Hu1
aT1ZsPbG2nqxuySeT9oD3NAAbUzHhI6fgr7cedHFZ9FBf7Wh0xd1pjetKj11usg1
kXiug7hHIAdI4VfTYNCtuPSqpgnyWkyww7w3qMCJxvYYdv3mlKlh3sGUjeKdeH+G
nadC89EayjY63XO+ethF9CwzJqpW5Uup1jKtGWIqZ8xa9sQB5mOSbbMXX26y7cfz
xXkcxIHa/Z946r5M9+8YbO+s3OwRCDvXAQVihw3tnY9Dt5y8gv3TOktyVLDCym2N
bIMk5TLL4Llbbg8rqYZFALEl9kADIwXyVhenD/KAA2aeYBvO1AA8BZ+0VKQ+fXE2
dE2GXkqlhywIJOpMc2cN2hF2FvJx3p1+tpMZniyKB+2j0S62tqMSQp1+j/k08GS1
fbfTXSzQ7KAgY3TLD3uJCsEHHmtZ++k29qCbCh5Mx6BEgExDPs6OuElJrhbea0kX
+lAqexPdjC1WJdEQUFg/Eb9kQmxeTIrWgKA5GoLnoe8Jf5Nq1+CsRF/xRkLEnqG6
346idtWZ6DfBU5qpre3LhuefZOa8ga+TIPrgVVSDIP0DtO5Rz48cU0aMnvDMpbYQ
+22ECmnjpHYlwuKc6YQsps+xPUGSfqIf+aSQL2Hc9WOlpUla/tV7iNJKDa31L8a3
/RUy1Yo6rzZwyhaElVodux3FHY90qNwjinD5Om6CdTeRtWensxse/61GRekG2ea9
99Gfra87SaCxJWd0IRutuKs9SGCnf6QLeX/I4leoecUIfWrnOp5vehkru0D7Tabx
QzYuHpRStvmHPRUWnbwjpE+4nHA1NEY8SEyKAXO6KPumWc+R4hSAK9lZTuM7gbig
VdoeaDvrcbuBJt82X5x81jRdhhglLl7AD8RkbG/YHHeM7WdOjpsgMCXJ0BeUdE6s
mRmYOE1LrQQru9vSBU5rn5Onz311vA2wanMzaxh5IWMe/EGYDVsqw3UQtyiQ01I6
uHFt9JeAU4xr/5qYdHyvkb/Q+DvsNEhA0FHbY0TmDcJR8BaAQr314Bgc0Ao7W7XM
0IXyvIWPk8QHpv+h0guYg8PJ5roYgBePDHVm6xt9gk0pGLy0yUTi5GY7gbBD/Lfu
nVD8TQ/uWItrVg7U843yHv6Z2rYrOPUYR9V/Rlf64oJkt1Zu7S/SMwaq17yqREKZ
5SCRrfS/k9kzLWFq0OZvkIW9Nb0MLfVIFhgP8ZBXjqwcfV0NtTBS4wBVQWIzjPIg
AfNdWM+hh0VVrjjmUudq4jUFLbHgc1e13Nu2TDQiS44nDUo7/P3ufaWZTnSGhT0M
fQHV8GJzmElVYOh+WLYVxHd3S6qkYFr+Wg/vPUKBDTopIqczveRMre670ZpYeWSo
hXbdRSWRbPOj0cPWqD4GWZ9hZEtFpGCiobWxdNAX5z9sNhuLmToGWnBd4xJVcROT
w+y0siuxPFjhYbK/qfdb1W6Vu0h1a79xC/UgGDsoyU5b7eH3+v/mxqtaa54wd8k+
qpKXPxqurKzH8pUHxbnjKBERi8hPCPL+eMdwijqZHZIE/r57fqj1mbnpdDuCDLYs
QPB6gPk3kON1/2GEZ9DWz6LcaMWc6q1VGRrVhD7PyVGIKnGJgBFIpCEk6+UdE1D3
Yq4fr2yGDN8x3xvgerC/FzhrxVSa0iGZyP6tq7rxUD00q79ARviMxUUG6PDb7TB0
S0MADNY0HRrApb3+Nbccsa/pC0/K4IslBOyK4fcZb+5rcCBMVUKD/2c1BH4BMAIk
5iLoAFNxZJ023vnr6FIm1D2IUps6mhV22Oyxt2b9Jhauoz6b3pyR2lqgVzMr0pv8
MQ0c/xK6n0ThYH91auvG6r1bqLK4pVbi+r5xITRtyzEqoA0aIMoQMaRiYRBDTzOi
+yXtXhTbGESki+Z1xbPVh8A2D/zoOwPGxm5rs2Bj9hCsU6/86RdQxcLkYN60F7hD
mJP0042Sqa5WBvk2UlSUXeNdOWc8VKpD8Yff5S6iC69GrSK2/HuOH7fjYaovlJs9
PLT19/eFje62bfp9Xwi4qocGk9NulZp7sECamxOKojRRBdk6cMhR9PL4/YpERuhM
/I4LmiyEt5zj5qmUIfUwL7v6JSEqZotDgxFtSJM075bMhh0shEbk7XMjuswQoR5p
iJQU6SQMxVDx4ALBCgoEv0zBvcxq6NuG7zsKL8/yy4lpHnV8gzMYRgMyzHfi8OYw
UbYNFCt8O8xwOwDj1C7Ts203ikQfzZeyh8YUU4qCcOUB+ooONWP9XgkS9KgEre/z
CY+5OQcqBBKKupSQA9hjLP/x+ZbYNaS6Lpzpw+1DTZSDyqdBuU+VMC4x3hvgwBdK
0m1gmJ0UAs1SC/Twfkg8GA7VDKpXdxHsGhqd/liG5G7EPpxczvNBqipxP3tcrheX
M8US3nPKV+s1QPNnu95dANTq2IV14C8NlPQYFQD6GCBuicBadcTYx5KYrw0S/LUq
cr/X+nOihYB77wPFXgq307dyuDXKChtgfbIPoQhAUFOCoQypXwXNBo6jX9beWpBB
F4C/es/yRmFbI6I71rASyOKq3YEm+OKpp0j0LlJ3RxG6hN9SDeOzvG5RKeaHS+fb
NGs7Itn+nMFbPl6X0OTzAIqMISH+7FY1WYTqitNjcDL0sgCA4jW8e5C2GE9s0SNC
rst4n4JVdRlFKwT0Hxrooe/CjxJBbMpPiEPiG1GWWezQey94W5FGdUxOailmhhYk
27p4qlQ+eyCuwGzQcXxALxoSin23/3sd/lpfcPImgT6bdaQXrHt+BffzMd4wSgzP
0PBe1iZDakgwJTGJTMiEIi0Wfn434Ye7fdQb+sPtt6UBBqo2DhkL2hIJUGI3Al12
6Uhrhgiz1QvE+1u+EZ7tFeZBtNu1M7WUjD6jXzrJnOwuM/pGTWzOZAe4V44rjjPX
RXGIU5yguHi3YnvaES1rAKYfpXkaDTRHjWgqhmJ7spnraaDMT+l8mROB2Bm8OZfz
ud0fZd27rWUJrbW+d758XlyGkNwtXC8cAgWUt9sPmI04+ZugFvvAoNkZ9VImUUO2
QzE3Ldkmbjzv14lEcNeDkscVdYzBIXL7xNCKFAWokEP1Cany/27n3m5NEd201w8J
9zqLXbB8/2jQh8NEQcCBQoT5jfii+8kDuGzrWRoUYL7OA97B6/b538ZnRsECnoIf
4aQHJSBblPgkD5OYLJ83nT85Lp7HX3CLUrNWy0L0Uu2vDZcxC3kIaFBDLaDChiAU
xB+4dZIo2GCLGH3zVWlpnPksVYza19+TDsmtt+WVmOzcX1EWuNinlVMa42UL3+V3
QpJQWKJAoXDQvilIt9PKcfVFjKKuyx3FwvwDiv2vi2eh2/5cZiarSV6QKQi1NrMf
bAH2ToUMEj2cabfc8Iao2/7OrXQEwMMzmhEB6O2FlxuZk3xVBp21xdNbSlXecWC+
ZjgMwa0GQkVsmHBd1f3dgl0gpDx+cNzrkM5Dtrjb7sM7eu/7WBGJqjIFKKdhtb4p
RamJME5R51X43U7BJFAnazkvhdaLxdhXN3B2DsmlPDY5fYzWMf4xsXpNevx30xTc
Jq/YHOzNaU6oNMX6nozozZ6P8MjXwoZW6bZS04kyA0lvf4zkf0YJvsCt05Z3oF9Y
K6fTyDgFoSvagNvyV03PPEo2DyK9b+voMLrkz/pdMDtpdo4Dva5MRYuzzkkQUyJx
Lh/OVFJV7WwwgNSqgQxI1DczDAinrBOKH4+yVTBExNX7ssKte+cmjSJTdogAxzzX
U89OOJAw6EW/13AyIq0Nw4hq/QuFcOZQal8AcQjvGbYw/sVZpn/JRehPI28R749u
pve02IBwljvOHGrVowTty5LYEJlfX/CeSFVmaDKSHk7fYV/l2JDaZLVVfFJTipvq
kFAG/hmSke2dRt+U4nrU0fPyX7LN5KQVPmnT/saokuY+LbTSmvQo2A8lz6DdEvXQ
U9V1mtHRE4aWHAjwTDXXE2IP/hbfTal8y8fldKTedklGx176kJMy92AI+N5S47af
o6flQeHG19ltasqpN1r2k+JNNOIx6kTEbhgeWnvKiEMhQ9r05xR2aqOlqUFSo2V9
T3fAIKRzy/3BiMYAd4zVz1SFFx0l8+iZDAiipPK/hUvMfMC8kb8M8MLx0b4cQVuk
hoa6LX0dQwP4q2ze12143IFq1rfE0QenP4WcE+c/X3awqcFh5dMYlbg7W8RpI/k8
4p/4LIQKq9CWOxtIDeh3m3DD21mUl/rZqfqkYwjdYNG4u7cpxLeGZcvnGx7MM3Wr
7P/2Md+gYwKSj37Xs+/NumqL7k7N3aREuhKTlGrwX0vzuF9Iq4oN+nSCte9S/3+n
5kgoJAN/d3GR8cfuyZywxmOkQZM/+waUTgR97Z4qYgpRmz6qr9xNeDvTUE6MlgQG
irN/d0wl+5gMu1KPpuWEXM94I/gGIwcwelha+6AwuE9vY6/YnMvQam8KRih3/gDt
4UyUFIOBMiVKM7Wh+qY3Hidjg8dZqtiCA1nzjiTueRyBHg72wYXOkG6Aw8lGCZP4
ZXCYss5bgO8dhlAxMfy7rHlIQuxTBP/Vg32k7p/d9jBpEp7HTZRuRKrax8R32wY8
SNP8RMy2Dqwo6zymxwjUksjfZE/5zhS65SzJ8KSsjpMbTNUJ9Ouq7ImszuDQ/Wom
d9AcQXOWQ3fc3DAs3LOH9lHAo4iPve5A+Wn4EGgwwQVSsMrw1yPSdHlqLkI/Pvyg
sE6zSz5i5yJ6W2aHn0fDrKXtxcILel6EtcZPPyeqTRXt+dbf+DP4xN2dGU6sGRtF
oO4PNxq0Ptff+BA/MJh/ICcgzi2uw2V4jmwVWkhm6aDs6kh/cro79bvp6vZR/QJr
skaj5gWF1c3WjMiH77as+qz323wU9Uo8eihOCbivnmIwFCAroDxDKEOlIu7VbSO3
f/rbfQyDdapae6WaNTH5F+A04vU5LoHjUYP3xuDyxZszX9IYzk8iEYu3cwMz3jMx
vOdKl7f6YcHJ0cDX1jfjlh/8aIFneJPv1MoK4XucT9R8pdhq3aaEGDnORgzwuSlQ
yFOpBHyJGky/Vt2VF8XyZ8nCNqzDONJn4oSpwBWF1Tfkv8SG+WK1Y8aL7vhjWzM0
dtIcocxTTDhnL0NLElYwJgO82NYOpYVaxiBVGJuRlGKMTBO4NYbYV+JY6p42Ai0c
A9CQjHIj/oTT+bCnJr+UAbtiHeQqnhBIret1m75ecN9Nu2hlYw+I5EgWgxNM7D10
ZYrZOm1TTKETMZnGTHyY1HjgEVOh+zBRk9XERUPDGZJ3+W+yT3UAvyXLbIgzVQQe
uSbsS4aDUD6eMS3RYNjwFcJ24I55DLwo7MUne4BddZGFJhq8KPaJYaV09DxPv/9o
rhQpYOvu29XdwhkUpuPhI47sXVDaLmFBmswbvjs3PS7ycq6J2eFldVDR1umkh4wv
G9HyzRKnHdRd+OB81waCXgyOi/CVJJu7C4sP3cgCDAZ/20hbUlH/aMzCJzJ/lvrI
fsj4OVsXLcx5Iz+yyKpDEeS9p0AldGSmOs3xgWbT+rtuUwzmmBcFTkz0XTu3rs0f
/4Gdxr89I/tGYX8SlEFT3TJJONdt4N0S6VjV0b8UGqr+R+C09oXkhj3BRyVwPERS
sQbqOsKfqmFMNFY0biJWpdgvKKDCvXjA8bo2/fTrPFsood5UkYf+SXx//RiLHJVe
lgu3K2O4yGFXZzOMgFIQNMjDRQoOG8ON26LkrvOqClipLnqJdCDVmP+ZDCawgB0W
cw1IsMRUjJQWvtLac2NKU1c3b47q6tQgWyyJyRZxtSgHC+XLvMTIqjN1Vj86xwRM
zbxPx3KBaAa3J9EoxN10JceOB2DXNLX8psBNRXLFzJerp0zc+JZNivua6dvAENmW
zdyyUIQrlX+bJZAzPU9hNpXZmdJ+nJ3u2RJF3eQL+cD3YOggemZUCcohFYWNgIck
pfytYJrtU9wzlBb5q0AFRxO8su0BvbdhpwRzagGOR0uFj90ieqw0ApERw3IV7ado
6p9SNQKvFDyV9ZYr/2Sh7koaTgX3yWwtDwCAvdyM0bZ6CUK9MScjauXznWCHVTlQ
ISHhUu3E5cUI+xsxb22+6JpxYaYd/bumHKmjLlARrd+iRW6Tld8+9KxZ00ssOran
rl48Q1DXSbbvMy6ZTq4JNxXrkHLsq4Tqoyww7y+g5OVXRMSV9UIBSTVvblX0GEFy
Xo5DqkvXr5w0QnDsKmeso6V0kay8ww/MfXoIzcEaG67VLChvyZwoZuEidL0CisJO
czWjggU0SMhcSxamt4D6MX4QGkP4WgA0WbvYOkP1JJ4/7m7kMBzUEGcWJsgKXPJ2
7RiifZGyBl4XavLFXLPJIcVLcfcYogBQVicNKU7mrDghdbC902ffmN+kiWBxVEUO
k4BqU5pjfjSMnwNPiLKRKUXhXMgeyLJ8BbtMrQCzTU9D7JLm5/ywO/ejqIwTVYrV
VT0KdioapuexmQIXLz/XtKCOaClw/EpUDZlNF85qnXjs82g7FMYzt1Zofc/v6Ub1
Urfp5cmq+7B8eg3QYonar3H2WJExDrNH9l2HOyxQNr5EgWNoLOhpqY/R7+GNeEBl
DpOebDXMBAArxoKw0XDW7Gn6P7sQw16HHN992O5ZJsBdquvi3ZSpLzFI49sGol9S
RxSI3RbhcBjhzfWDxGNh1kokriF4Adjf5cKsYAskj8ap4S63l259GV27Cg750TfA
84eUeSQsPZTCcf/ID/EQ2Xy36EB5Crx1S0hU8HknOCG6wSYiZ4atWOdS/lfiqTSf
QWHZCR7G+jEM1JVAnac6oyxnOXuqbyd1kOhoPizX3xeMsnFEXkFHJBBsoxUmsFCy
ZZS6mgu1G82hMiAEShSC5Qcxaeq1HRPYDvgzzvWp1S6Boeaj9ISu3y+xmysQnddb
oZRow/yQ6gjzFe9QqVjealswDQqwmaaKp2N8Rx2FKELo9qWCWwVIRt+0kwLbwy05
oYSexi1C3AZ5A9lsMzPXxd3bSGSXwyCsIdOfHftwC7gtNjS9Zslggon3UZNVxOh6
yKY366P4pZW+makfPrOiW9y3JLd00HYty0Ej4x5v7qTQ7zUjSKtIeceUgypXMGWa
SahQToNmkRmWSNo6qDcNWOagwHKv6v+Xt3pxtpIbCjrjAS2dT6wlWYGI9CHit6Vy
HojTZBWvU+Nl8phsIPpslYdgn1ZUSB2DqroKzs20d6XCFt0gt8XWSBYToc7znnLB
IaG1knuUWbhyFMmzpfRkyqLuGSVJaRmG3Z74dkJzu27PF6Gw1LW/MDYFN1cUzvlx
k/o+mOSZbfo1ZVR893XObmx0/fD+UNKqVeALSrRosyhfTlLx0sWe4tJ8wByYbUwi
7cQRNV7IlZJSXI4WX+kW1E+/SvXVaPXlJvG+Uuu3sSm7QNyOZuKKvOjiQHdWEa7l
1rNMT9gI//AeXKpqWFG4RZouykhdek7Onz9F/UhD8h98eA3PgaLZXeZxNesHNtGF
VUS0g7qRQXUlf1K7Yev2silXOrZ/o/pLtKnGW5AX4xIsixFYnspDedWua9e7NLIq
yiGxJjd5S4zn0+It0UPHLys5KsFWvDCYizkdngZKWpTBZqQHFdiEDpXNXsdNjzhD
EN7q1dlZBrZPoTp0Grf/Qy1B7SuKiBArUH02tkZMsRoQ4bYaNgu95aTWlvgufNP4
86Eopx/FGPRlbV+ZxzeJy+J8wnrzYc0KYJ4x41n28+qL/vcqf4rX3gCJSHcw25gA
IriFTnDthf/E2h9x5U12ILp9QPl7R47BC11RHGSSQ8xHO+WgMWBwXYFkNZod9ieb
9/8+juCKgnw7tZyxsO0LYHfgrR4IYHPtm8jgt+pcS8i4SywWbv2OXo0Ym1MnFOVs
8ZcokA0eF4eGsVUWgplaBR/9VEzmjtS7lChni4oc0USDmIV3GCfutlo2YDYi3ZDQ
nengAnr32ztwiIUSqod0yHMSfj0qvYna8ouNoVQC0L6ug9Gm0BnQgvZqOdVErzyh
lZD1fo02Nvwooy9swQICm9HRGj4GGj58U/gDgAerxS/ZwA1rO6VPxFNqmeex6yj7
xJGqluX/sSW9pwYI0AbGJt7QlMyGSMgDXCE/5Ux4v/tTzEW23Ylt6a2fV56XVW1W
XjsXOEXjHkJMGhY8FHkFiOATQ7r6a43l2Kxr0uHfLhkOgIPEjvSM9pa2geIAFL2l
x7bIkkipsgEQNkfJySijsKql+KJmLW/Kr0IQkVG3P2lHh+LMtiUb1RwD+YS5bOXH
B3wzs/jdMxcNypRJxwtjJFvw1GQuxv0D7cfEKgZtBm5QR1CtEkhi6oUQRU+1+iMk
yGfim9hLZS3WTE5+Ovy4RYDNcwWSdGic8vOeC5SLzyHQ0KKK0tiltCBtMuAIjE/B
9e6lKSUVc/UGZ+pikjL6vE9UeHtxooI1Gk45420xVTl5Gn2F70/V+VLAm3amhkQT
PBU94Nz5FcdLB4Ie9BM2FM3fq1S5Dj1qAO1kcpYAseLXZhFMaNYoRrNeUFNEKVjo
V5cGAVvlcI5v1coZQSTKPC+kzG2xQepiVNZrfe6FNBkXTXT8DkVRQVOpwCJlaZUd
Ec2IRRx7rSuhzbmAyh5v5ywsl8kvm5kdCotzR+mKWAOGSEn1OOoA2oSb4J4XB0R3
QwrXfFAkAJtCeW1AaRo/1Dk+yhKkKcSahdPXoEgvfAyjNRoFpeL6ZtRsi1337bCg
9hJmHdzwCreZL5vRYGnG93CWaURKlEszeWC581uA6e2ARI0EoMgZTC96BMe9UmNE
L+Khm0rzEPBF8uSWbmA+woMTp0ZmC5p6/+m25yLpaAJmhHuuR8X7gpdzV2nf99yy
YmA+XW33t4b3mGA7n53JYPoegEv3ytunL4I3Amul0dS2CEbSIHqWwjPuC2JCIXl+
wcy9QHpqleROXVNhaIbB99n43ip5gcftVYoKCDfLCBtQQkWareQBu9nk05yXBmO/
KUd+9+0BMz+c6y6SJ1lMN7CYc/NFc3zSUSKj7PZzBItoMGXdjC4v++wSd/BUTvUg
0rWX5sMKw9TY2ykYVTwoL5q5u70ta/0dcaSbSzZlKlsh+5X2GKlVNUX4+1zSEW1Y
dhwUhHbKVUa1satpK3p0ogP4rJJn5ThAln9yDivM8l9EC6j8EBJ0vzXQ5HqGsW9Z
WQ4g7TbnfN2zrEezQuQX0yACss4wv3z3LtSvvlG1sxF4Z85u56YWzJW/l18OjbqB
umickzZoWlYpkOecwatseB9dBVX+TGagzoO3dQpcCrv+eQqTwcbxwBJPJlLHFITv
6WTty1gV3m6uDin4A0EhM+Yl+g+g6SscDh/661RAV7gAqu8hl7fSN7czoMdjNxcz
GLEdJVeM6cmSne05yRKpzL0lGhBXBlG2LkaDXnoExPzkpZav7oVt3/vw5z47LU6b
Y54I+1kFqzFv930lIaCaWrKDZkAyCfNei38HgXOCDeXcfx5lS5zn0BsSiPxRWBBe
Cp+vscCxgLbhsPeN//04hYXKMY3fIkYPH9QDRzh/oK0E3oapDKJsQ/Au2GUfZ91s
HiKQKshf510iQ4FjWttHjizEZC01/1q/XbUsSaDNcKwg9MQfmoF6aizf74P6zKZh
D1scIawAE2YyRAnqApizFy+VO7smxM2qXYbTI6yTFqRWnUkBNqzmAKeS7M6yvEsu
YwFJifcanMqwjNFksvdrdGTdFhqHZBnHyB5GHmYEspzdVgyiJic/epzLP+yNofJM
vmk7js9zjAw+cCnGYwswk7+9wbMOE3qH2KMPd+IfAqOD69IrAsDYmlapxrMlcs1m
j7pwzTubDocmNtKQOYFpI06GNNflWsDr/eypeLuDP1JJdFdoS3tIrVED0shHWVgb
o7kT5yQbGVgh1HAAPyyKl8YnlJ+16kbhHCLTKJkZbbC3OnJVgTRJpiRUkPsK3EKn
B10yipCdPYY3t9Hp+y5VLhYFVom1GMOJ+P79FfWwe8A5/rdpT1moQS4IV+4Ikv4W
6A9YAGHHoEI65EMvaamNAfN/wRIfgAyhY5XHWo0UeT2UYO5h7CWgjhoE1/3PCOgT
akiNgTsQ1/7xopLr0FdYDCHUG1cDb1neqJTTdFTHlNwexyZc7fVU10iDcy9sreKm
6cmqe5+THjcEnKDzY2RqTk5VLCMgH7ABzzFOEhbup2Cs1LdRogisvC7gQqmSNX/Q
IYj7I9tPbZi1ULwZAFsI9ZjAS19UOugVEpNWVptCnQCWEUKyd0U36Y57WiM6ipDY
4BmA7v2Ue4ek4u84xTetxOenhRVFE+Yni80V0UZj9epPd0bJP6xcp+2hMIaI1fmx
lei76Gqwar/6sIXM/V4aHBZ9LXsLeY7aJiSSYUZhcxBHUbrxpJ8Yl534ozNZrJDc
0swYLn1C0WVZXI4632lponFSU6LCNYuD0efDxvQzPrMizBxxGA0mk4uttqXFeEhb
fHXJ5/KxxHYNNwywMztWs86WOmxDTB6xS0OWvz3NHXA5YEOyZh/PhzJHx/e0hUcf
2OHt3ceCMnw2BIVaCTg9Wj658FDfnBR4VmPWBFIEcC7Qh033wWUvyn5IRd/7KX/H
lgAP4DhADWGlY1V0kcZGpnYB7Tq4ie6XSHD3i/Kpb1LWo/h2aYzR2/XQbIpu1QUi
KwJE9AVBBpdSOSK8kQ8Zsuika2HHRAfc7hD0g1Zn4XJ6ZG0SVDVhxP7/oE+JEU9J
H4bxvGFsbsfeBeTmaI8N++sTBmvF9eHC6vkmzCNfSfrUAPsHl/L5FNllZ8zphBzN
3w3VyTMOH99c3F0WRwQQvK+bJgqbZHRikHVFIJL9XGnbh+o0OX9+eCn0EibPnESk
o5oqE7Xj1leGaKcvX7OI/KU/T4yzUp50z01cqDQj0XovB+YqubvyiICwxyEvqloU
/SS2l37OEgmMyIQvNo64apmaLyitKtixi+//+0uQ08VLXJdmM6NLKcCjxZAlwQ5V
W3OzGQNruXzNdXGJrCsrq0ZwsqQXfHUmuFVzb/pfMT144ExnjVjmHtADxvGIZEg+
vfv62FekexhbjT37fv/u3DxUdyXszOt64rXf7Xtb3pA098EZ5T5+buAD0MwZElgZ
x79DJ95UsCaxeuFWh6t68OtLO4d41e+SSgdEsZ2G1+fcKtOPhw2Z0X2ziIkQq7VR
4681cGdwCsoU4S7PijTPrOaLPoF1h7Z/6fCtHtuVtkNcqQMq8pny5H4COfr1HXx/
5/F9LSTyrsU3IvfxuA2xUmWlg+n3eDsrY9fj2qwL/sAPB/U/GxaiYuFrPdU9QDt9
xXrZdYUYRpkYYWY5V65DQpZ7bCwGOl8yi1LvZ45K9E65XZXuhRPPLal0X8JbVnT8
igL895vIV7ysNtXIGPaDsh1tA7JYs/TFabh1UG7RCCTdTeIEXkEmDGPCo2eEKmKi
f5ce8l/nqmrceHZOhUXje2XMLj5qi3jbJ4p/8cKdIF4HqEi501EImLpi5uVsRoJQ
FSOjY+2gPfZTURhVNANuapgR7EegzUmyTIR+8EMAr8c3hL9uR+mtF9H5HElxBSxb
B8NRK6YjR6eaXU7QJxglVZRmHFMn+Qq2uFMdnSiU72vV5laLDhEUvxWuP2fhsRre
f+TmBo2tv3GsPHyv3QV4nbVrBDpM84DsqW0qQuvztwdH5g0OWwPCRlHwG8qtniEd
e0Yt4kdV9plC2IAXvh9Xb8cukRMU/n59SpKoClet/NiwaG+Mc8wgoMIDnT4TUm2r
rMc6EgKOl0XgsPNBHudiBlHSXmMTa3s6vHMpdzBCt/4norGBNb+3XJMGDRYjXNlQ
pxeT/e2HTWnqhvLRODu2L5sqK7glYKDn9GVZ8mvQIFHFEqitjcI7CnTVFwPV9zNH
yw5cz7vRF0j0cSWhz3HpqA2+FLKEQPPvIZKF6uWm36xSEPtkcTazfiznwkhnmtE/
QFKGAbKR0T2iKTj6vCho7FRRZMMEAOLHfKtjIHSVr8awtUxvtPNn3odmmji6Hhz3
nTClgIUIAqZYjiRmaB/oZKZyGeB9FgcJioFPjT6APNeLOswBExQvL/aVCcER0yMC
M7/POhrrLbta+NHpdWce+AEFN4LiS+BE0Vrb2of3bq2BepuLp/PytXA6NBEFfZ9v
dXk8wxwZ7nBbVW9APAprM/YITuHyspIqpAp7tpEH7cRPqT3ZaYIII72JV6yCBRb4
Elg9TK08mB8eZ+WB2s7cvY2/gNTy3m3Xd4MxOzlwJ97hxRp6C5/NXDhUak/aAQLl
mJkxad6gTHWZB2YzEyu+AUCywrcBE8c1aF6IPX0CFO7QW7o/Fa4leI11kBK7EBFV
7JzQ+m/vRV6f7BDcSdMSQtK/nAGF/L2PzJG2+WH7q/rDe8GWvfT1AYhzQjtKOlDS
ItJyZ+zaPyeWD15pBHeTjlDlSV6La+G8bw6J/x2BWIPyBQPVIe2i/K4DJ9ch8dgz
Q3/Jdgn5MXR3SCB8IadFND4lxI0xbG1a5BYBsbPxSh7XVf6xnMs2Ba1qTI6zAUKO
apl5GRD8iM2zd6pOT7Q7qWtxHa4xDxFUXipj2zf1v8g0oyPyBlrVZ/Z8jOfcDC1d
O5bCYP8/rWxJ5xlCm5fPAeCaEuiny9Vk+gdD3OPnQ0v8sCWnBY/PkgqQkRqsKAo2
P2M1l+XkPOQdfCNE8JChqXLNXbSqPGEK6IWh8immEzGWvzj+/RhJo6AsPgaiKStK
yE8Bf3rZXFB0wc29NhZQLrbWXFEvGA9APzJBYPJ+ovE2aEoJoFDdT7gzM5zCJ2yQ
unqFPPpPoqPsG1kuT0EyRQ2uk/EGGkLX5HezJOQY2bskTQSmospiNkz0h5NIzp6k
rfEUaClFU7ypvwzc4Ft5kKKNyeVC3W51KezasptEHTVTFu0JESVWFrSUyiy6pOTv
TNJXeLWRozTFRQzxa3snwsQ5P6nkEDsluQ4GtUpZmydgINjWjcMAhEQUAhlB+YK7
Mbxu+nefR790quhX35bJgEknOp6iyovvKud6PECbpjS3XzgjJ4YwG9RzGenB71Qa
O8lNIPoeCjtJhYlA4lXqgc09hpGRpWwICTlfRtH8YJ5RagepKmmCjGsYahrlY7F/
NhsG1dnxuF34E9kSWp6aRr/ds56Tk2bFpfrAHO140HNwGEspQSPIGJIzyRZJ2Fc3
1RteDo/k3gWF8PYQKgGQjjgLTY/+0K3vbDPI3Pa8DUcrp6QoDjOUZ4E6bBZ9OpRl
hUIJ4OJ6oPx2/a6btEI0LFfTbO3yPh0XwQRaxxsoXCCi1LvcoZHiDASaoIx0BdbX
/SgT/gWhwdN/+p3xvPGTomyCT3aVx9HwLpNBr6rWgaJRVoVJhCtMrJCHqYd888FI
hvHTu5oX14X31YwanlHCRj0v6S0FFmbYsJ+MfpZCsE6LupQzelKN/9xdljfG0wCS
baLYWtnLceQ5LI5GFiiRv3DqZLg0oXEel79XaEzHJ1TQQdsoe6AFcIpavqsmapcH
LfwP8Y+yq9fbPdlTm/Ivur0F5KPpoLFLU/5w5hylwTPU2jEowcqpNwZ6VIuV3vhR
bPvjMlA4o/m/JVjuaWb4xJ+ZmWuSQ31vlqm81LyYVr91joGCNzuiyaiR9ztaObux
ge3HKSOHnoWEAK2EbxidmhBK0NxQSRSiDFATPrJcnLvF7l6uMa4qWvcYq8EGCFrQ
62YJbISl/uJUIRY/M6Cafj0VRlijizI1Lwurdbhn6oPBJB7nbA1J888N5NmcPYVL
4e/+lPohagqfNMsrttL0kmpiKXTgL6zGSjW8GPoqbGDm14xrSsO+KUX5X96B3Ntj
8liV+QRBs2xDFSZmaRb9LZluzZeZXrWAf3FMjaDuPCqztrUzjxIzyhEn0Qchmo51
BDFAt0ZMYOMn3Jmz0CwECmjNLJ4hptHUY3uHaUErHXCuYfkE2PBO5GsG5S8j2ndp
bQcEEYRl1bfk0cuK03D4pakg39F2V8aC9j07DTgM6zFHooI0hsTEyGlfoqF2TV/k
pldAFcJjT8q+j2k/BiqMSoTOpzYar8Y3knQfvumSY0FpHUHZpsGX0gjG5SMFp/sh
Bd5uhPNIFQYeYbpou5YOnOQKD7mUib5+h18nsWuDAs9jSYz34XaSeswHQ1DX/VoT
0UEH2Ni1anQJSrdPotrLN1L21HRTNMa+bfAsbmvgyTqN7p8BKZRCGqcB526fe4uv
fAsWaTSckYdxHVveq+JZcVa1GOu5RaGQwbutBbgFCw2or9u4x8pBFpRoTVMAXGNf
TB2YD5CPrLcJwzJEOUD6I0QynIgiHBgSeB4/X5u4IkWrz5jOsS+o+uMZ78bmU+ou
FPOi5NhB316F6B39CerKPq1Nernvgdqsrx4F5gbGOEFfQzJHlQC5+p9rWxQHJpDu
kzeXUowMJP0+2Ar2iFY5nryQgz3/od5xqTDfKEBJlq6fFwHdLP5vfSRmsU5gPOKz
u8VnQgpDkR3L1QOskxbh4k+CK+X+wnavSYI0sXQd3X53oaZbW+6nEmIiOV3GW/hr
rweyFU8ssNRhDw5lqoONT8Vypsk88OJWSrxlcExMDxsfovIgIWHccQJyZPUyHNuY
MOrUOjbp6HHZK3x8mI+M3leAmLAdj9LGTSBrLT3nAWG6ly46nujAf1xvyC07HRip
7fH+sAeyysScbtc8/rWH1IDg7MJfbWko8BQlXRfjyObC7iBeT/jp1ommwTGw64/A
LfvCNop0Pod9EXnndy2mj9eLDh+gEMB8vmt0nDqKX9Nystf+rrjVcYc/nKU1CqFo
/I7/Fz274m2tQXJSkAH3U5h/OE7ZO73Sp+DBzUa4aDVofn5e8Tt7OAwEqkNDGV7t
YTOVS6x9lDs+dnUk/9AscLTLmKk+MPWLKYYCZmxZoTVXZLf2P/XKWK8Kl6RKc49t
Eiy6TAc0wl1E/iFTb+21OQpOHne1+g7f+GqiClMNGnePfRueDiGLffEsYW6rttvJ
vJQGm2vKELy5rzxeU77vIlre8+xxxiKKmcgpxNumN1eetsr7PNZqgQtjvxQjaJ07
GCR86CDnl1sJ+q8y0lJgyNtdF/NkkhUTvM3qPED3xxOObqT57xuJ/FBSpxq/v0Sr
d5sh8Db8M82eX0Dxg5QLv5d8be63ep9D3LxpBlKuEd7v/MloAYjY2MZmG7E7JlRB
Qm4QsGha19sDQ3L0HyGL52NMCRCi5IrGHhGvb7qIDAe7pgx2AJ1IvjQSyIjyIwtP
6Ifz2WD//nJf9+k5035FhpML2QCwNHCqJ0y+o+u/ObZYkWXjvVCigOnlOKGIW5rG
pWHoQP2pWtSkL00uWu04fklIY3ziLOQvYwBjY5e1zWhaZCfGwAXzAAaacRCVAToU
392Lcw6NRxTRUcDAmNz0/Z/L4OUe11EwLkHCyq0WvuSVd7K+M78dgBjfmMkBwOtw
qPm3FXBkEkHj6gaK4HAV7reMdJ8xCnAXjbJ8K6N8pdWIrdpBgeD9Ey2TuZj5RXO0
QJuIWEyWpEKC/2JNiHJOgMb3V2mHmsormsSePU1jXfHlkEbg6EMni2NComxnu6qA
EeHIcr9OlAUdDSmAn9rMCmA8WYWCKOpdKPtwHIuLbelYm5Lxg2jp2thFRTGLeQSx
DwSv6RtkFDWDPg1czw70cVmuL7ewEBXTqGUg7XiLYrFwRdI+/9TLtJ9Bk4/D+LgF
JYmGGtbsuP19D9U7fjG9f7E6+wznlj8Z30QSYLh43+QMIZ2Irr0PuGof+bJw3110
T3x2f75w7vJcyHJKzmiSju9M3wPBU63AqyuJucYWw0BPje9X0aKZ1fxw0oWBPnmo
QWJY1EjUALq343lJxdUwkPCp6OngdSqmEFAd2FhC40tBAMqrlIsqVXxDJkPNKPFR
G9Jy+Xptcig6SIDcVQJdhRq8OHNZK5fRoXMnYCbzRTHcvjL7RtoQKh6naKdsDfbi
hwHLn1OVb3Px4eJefRScvHiFvucl2Q1wFusKFwDOkLtMxMQIhi5N4fe1ZtjtAuBw
r9JTqc3GshKWRlEhQAxHoju/Q+0kVz2+LtFC6tAB3+sb63VeqUSTjIuXNR6E1367
lIvlCBHkzIVvGOaI7IGARGOfLOyJlQWFPKDb/Y6/nXJt3jZ/zJ4tRCeHu+DREVta
9aG4Dy+mmTaLo39b0G4zHJ70F2gDPEOLEiot7fPXlgWYf3fojkeQYWue4SWn/341
4gdUt7LdO6e4Tiji7kQv5Bb+XPhPWxwSmIKtS6cKTCABnD+FMW2QKZ8Qv2o5yO/v
f6K467JYpJNvj6oXhv5b9tawauQpAzvQzG0KiHlbKRbkiwcBoMWSlQBwR8E6k9Zn
441q1A3eM8qDystr0g+Mj2yN2VSu3A4FyvWYdi4ctjvD52NOrmfcGoJqgtMHZ9Cp
phkxlfltSATNDMdmDINpmTjHd33oYONV5Duy1MJBh6jYLmmiUX7S6EZ7NmYC0JXa
9AGJULwW4oLwEW+AHbiAFge3BrP9M4M1meMKS/JWXL59wVKbie2K9hBz+lVVjXF3
B2PbTOTSfxmH99YfHIo7NT1YJfERWcjYTANmJtreqQfAF6lkM8QrZBcsT3AywpDn
YGZJ+FCQOuPUvO9YyZ9Jvg2xsxoqGjJwHvl9zbKe1ysbreitgN8BvimuKt5Rwfb5
VmBKQ0mrjGVklPDw7NvOcJDyY66MpHgVo8+VkXUHuHwU4VGm3au4gO2V68a6iYA+
B3oGa2WZ6lSpQoW8QwV43cuUOoQ7iTq/E/KKYpJq3ub4DZ4z6wlNRNtNYaC+oisw
zIqcf9cJBcILR9x0k+UtB83v1WSKHb4YGi3x8BxdhlS90LRzeU+73tH5cYP5N8IM
tp+xO/XFr+WpHoj9rR7x6IH51d+dy/+g/LauTUJ3sb4AXXGYDn5e2pB+7JF477/F
F47VLf694RQ1CXWI5Hk7llqxXk0bEa5kZ3wUI1ZJHgRv+p/9L8QPBKq1tREOAOBL
+/x609BOuf1ycy7MZPNUyol6mZPMR5jH91XFoqxcWVxtLFa686f+mwgjwwn2Tht+
kBgXQ4/XMmoHLNCOvoeB9DF/NG9F2qIYp6zRJiFKcd4ndibxValVxKBnQMJ9UBvo
U8YoPZ60ueGB8cWIeqRqmAc/u9w1ElOhurfITtXjZaDVHWhumYEHYJZmw1v34XDh
hiP+EvQuYY8+r+FxDnuqJ8oMK+jZG6UX3jWzkJhNMdcHrFyLTbkLL7ErBlNJSkaW
mwLd3JwHf/gdtuGZLO2uaM3eQr3oe8+w34KcF/9UKVNqkAJOX80LVt5g7nkAKARH
wn5edluKwtVGv8lnso6GDWDNnGY+ciOaw2rvdq9NCGcwYjWb43UyQ0CtbrtSImnS
fWbG/Si4bdHfZzyDEDDt8nQQ85oLf0mfg+Igxrny1CKdwuKVGEORxx9L8VX+pz+V
6erwX8rrE2y7pN8IMzqzezm0Z4k3RrupX/ceg9kWJrZsiDHfho1nR8NEL/s2x2vq
dqzKdNFJ9j5YDp3l6KtAQzlI/HXUCUK66WEQgb8vq0VFFGAhlpX20E4EL8Nn2jlO
4m94MRG5yp0wA6DqVzG9k14ewFiR9zGcXuGux1SUIcXSIsy3h2WjYbYd02q29ci3
uDrxYQsiUR2+XfBsnYMEvsUK5egV/KkmDoELKpn878qrQvSzbI2Dg7ixyBEK8O8a
N1XFmb6kRuT+UTlRUh0UdJGtQ48A/GdnzGq5o33cCBYNVr9yJO0Rgs6WOvguQDsX
rePk7WknQ7UJcNR4PhlhLMVkXDRsoHtcL16uYWfE+9JrnDXN/1LH/XG5A7VqudaJ
x67HWt9uTOSItkOl2oIbzTvlypWaIIrLG52DrsdDZO+BudHgZM+FQaixoFzT2CT9
ZsD0HV4FYspVukdI7WiqMWTYCc9h+9FxDaSY6zhZx582ChanrlV5+kGFxg1HOrBx
1wtpbUUlArrXAOdxNslFrMOoSonNd+ESyghyJROIocCMsu7s2L5Xj8KxUk5veMY7
uLZFFqWyXRjfFOfJtnNarPucwnJhvEAznlJ/ahzlL+zVIXBHWauI2wz5msCNwvQU
AyBiRuogwRQ3FkmJq2AQRNmVSyOWagLiWeNRprG4KYH4IahQlzQ5f398k5TEtCih
ZxFJN4MVx3jCuMu+w2+v5oebJd9EzmNGvCOgO6yn9KM4O8G+WmFUvtC1oen6QKc5
MAKz5PBKXpYotlmYA7K99tpYMqLi/eEgpfPKhybvJZ4zvZQbIBpYaGeMIAgeyZvk
ldAjsLAIwMo7v3iRUcMPVNMmEaQcy3ukBsokmGP/5DBLlLZGX5KyEo1sbWTsHeHp
BqiI/jVnJUnU8I9quyet4FZLW3rdoeRGTeIyshqsl2UU/GpsXkY1ByoB4gqBylas
BaonXCo/XiSin/WGL0D30GDd4Rhf+4o5kKckzOZtKnMRuJ1k1J+yMR8RUG2Xit63
0rFCg1CSI6EDQ0pIbQdO9PDcEcHGzXKug/5igUep3rEk1UaGEEZxBXqxvygThfry
LUhk6sXPkIarqJf8PhYqsYXg+OFwWrT5A14C9v4NThfYCTEV9L+19loF/ILe6PL8
OOBiEOZCkIaWLFnj01b5pgDBX4NBbzJuBk1OprmZDcIkPeS/dk23EItaXEnBJtdf
R1NcrNBBCQZteiep8tEPO+mW71nTSRVv6jQPy4j50dopfy1SIMLTP7hH1CCD8Me5
h1QywAjx3pyceMHLSPcMdBYBDzXvB7Lg1H6g+4/9UGgaNbcnm7OeDOv4RKuAXLA0
VwhVtLM/KnHYpnJhmyvnOW6b1lFUraQiuk7P32LH8aMHiQXUUFYUEpHgkavdPQgS
fj16/gF4pXbVRmLQT5dVtL9v7FZ4VlBp7v1gB0NDYeb6rlfzrvp1kgzsvKMePBPT
mjPB1UXS47LlDUyfUfqdIoq2VYrBd7q3WdLQMsThU8Xv4Ws0K/3Olr0TLHfivE+Y
0aJs6UgJvNTNbw6RJ7kBRwYTlT/UIcBYDXGv9qxbvzhe7pVmQrX2VjAh9VwYR1lu
J1uTfhzjhPImPIw4Z8pxJ7yBNWswqN0Y1AlUrIyzvUb2b7e1LReHt9FY2v1kvjhz
aYJ+G/UGeN9HhFrEvfpZbdkK/HiAFHq2lGhb3IcAHZvuNU5S9WyxV/E6SmsBWPPc
uzt40h98jM7hCEXaePGhSFsGBT3W/OHRNvrPJD2AP4/Fr3S5suW4uQmKemSQCrIa
7c1OXLsgEgOXBNxJYecUcurm0fX05RHrd/VJLreNQ947UY0VRVcZ7pGJkBxLQcDA
eWuobjzanBuouXgKliJQHR2kJmYwoF2d7tHgLDEJiajs6Zz1ANWbd7gKtKWqP4/V
aQ8PSyfKqKttDiezo/7LdLT9lAqbVdH2AIDUrq7qFYa68KyswpvisK+Rwjva84uw
ufcg8xOFWvW/yjO3KIDvdHqfh2Ok+XLRIj6fSaVZRrMizu9eLBXfLttobD2kIr/M
6pnPy9Kf4CUxlHdNTAdrkU5nqP1PqrF6BzJv2NN6QbOe05JsCMsBBdkcSDNiDwoO
Cnn8cjDn4C8HOXxu5IuI68FANKbUQI6HgYF0mnqAPZ+zWsrIUr8yEvuXv4xSDyeN
wPzDiwmZDBDQFMSTwIEQhaql3VFunrTotMimFrg4iDyUbb/k2o0R0NDgbA7/0bsu
MC6pFBzlLWC00+mwPxyndQkWDtsfn9B/06h6gA3VNsUlEaV2u9qxKPjfVJhaAg8X
ZFzLMFk3EiVCJQ07dr0NrGgZN2GMkqzB6ZBCVzmhacbtefMqmR/NZ+/+5Bsu54q1
GZIoV+fcRwepFiTzHEoQ2Zm7D/B+xa5Z2RaZ/YgfUrPNMsHj5NQzhhbxOVpvma4F
GnaHRHQrsCQaX3o4Ygk1pUOvihWKxedR0ceHCOOJHVR6fn1yesp89QGjt6Prq4Rf
wZhy4rVifDTFYPNduw+geya3t84KKv1V2XvrnRjTSGW9L47aKIAu2IhAN85ZMg0O
CKhNWxjfcj/0mavGwhn/bIIvFnaNKR2gOLWgwiVfNdvM35kJMMfUW0uKLPaiLUza
E0dK2rfKX6lSPeGPWd2//8Y8npYHx/05JW9k3ljBFZ+UMFGNx2VOc0f8BPZ1vAmf
CnkfLVz1LzoClpG/Fx57dmp/w8yjn2x7pmBUgq0W/8rI3/TojRlgDJXxkkC/hM4b
65Q2AOf0DhXLxkZCdsDnykecEngv/IQ/0E74TFuW2AvyLRw6YtbFk+PZ3QUB4Vp0
puEalv5QrkQbestFJkdHAEnx2GExxiztVWLA62f+PyIseOpxtVqB28rm7aWH83qw
FO9OGUvA1qNNiIV84bOF+TYeqYEqyha4I/pA0N8MKMoHz7edQ3WLpsRlUHbpTReU
pENdx2/4MUOYCNGuzxDDfbPtd44RTJjQyh2dtL84Vz8ybjm06Vr2MIaI32QbjDWm
yz+V0faeuFWoyTck57XwhPnad14cB26a7JHucMBo4k6aMBnuTtAVRBzl4Q0L4w39
TR125Q0KW1pXRcmcMqasPTqrZNK/pMxHyHq5wNg+2aQbyyWkFL263HJPK1hCx7P8
9q/f1+YLCKOprp217YifD1YJSuGTbNEG6xLA5aV0PksCS/uhTfhfn0PB/0z1DuXW
t3F58uvNSVf9IXe84S3st6v2Gdy/PkgJyKaoMdErFwlIc7t70MaAznMrQswaI++a
GHL2ZvC+Sf8a40E3jZ1IOjUeLsSfGvR1TTlcuDRSMS+ZIknbIook59OxV96KvQIX
Ojoto4N1e+CSlcb0wCNEzEMtsm4FWwSY16iy6ART6h43B5iLg9K0tUZ4eWQFo0qp
R1aUFHTKA1cXa3PJ5rhD+N24MD9zlQm2gFx2ipjxxcW194pvue/K2JQeoq74rqh5
FFG9Dz9h0/hpYeAPTmStuOQowNsW3BCCAhb5ir8IIqt4bpoaSHXgjTtAOdSYr0GV
1Oc/smL0c6zzo4jUdEF1iVpN5ovICrzr3aNYAUf2SFUoSl5pvuklpTRfyoN5WsDP
t0Ncy6GfQEgwolWexI+eDh5gl4Wlr0SPfzuJCMFK3xhCWuwX8eWEqK32vf+BrY8o
xt6qU1tOlUw0ajVJU3u+M3+uNI70bWlQI3h4y6JYwM8rBsbAoLEgzmjSOJgYwe8Z
MunCOBSlQ62cbVu9FV+H72j9PMuQ9g6W6KR8GNiheynv13qx5tm/cSAeu7JchoYu
AqRwmcfvL1yJoPv3kPGJ/+TxbJPttlEh/mdIEHMozgaSSSKUkCT0OTD98jYHI/am
hjlcV3qpSK0tAbkYsMgXUpHjZfOUjJOxUwSww/6Xcl/MR3f5p07kmUYa87O02OWa
Cu78UdmrS1dl6ODVIM6bSa9WI5bPxTVmhGEVS8Wq6p5VU9uWI2Itky+Sg+T2mfyo
GSnhIvZqrzqXzt2QI2MBiyg2LI6qA/KBs8MMxzEHkEid1HSNCx9sDpEiAlZRitKx
sPQbtlFSaLjCLWaZkcIz3SWjtdGoD5s177UA/SXFWYPaFt36PloGK3DW6GpRPMHw
1vnZ9Nra4BwysHGdQB4HYnWdiQvffj/yksE/PGVZf2F492I3BzanebZdOoxibkkC
LRB1EISOyt0ED6tz56If8tfxJoe4TgIgzQbi5xsQvIFFDleWtL4Tf14Q2YmPc74j
Un/Z+CXBLVJAo+Os8GXzbxN6EgpRYnu2/AMEXXE2e8dR9emPL4DGPhV0rW0YOnyV
rpPczNCycQiwg5Q7ZoLUeHdLwcWSQjzdZ0z5GnuvXlAVx6ZIFMVfgJPaalPZqviR
Ub08loxnL2MQtt8e8A6aBCiNear9BFQTpC+dsFpT81N5q+DQN61k2GJlgnum4roy
R4lZUqGrdKAt0DLXnSiQ/Rkp6JXotLCZMxS1alsMQCc2YJpjXW24JSkIpqplMWF0
yyIthXDkVcSl58N5nWwvRF9RgSbLdxhvs2UnnsWJPTF9rnsCQ6p1wy9Z0Xbx/bzL
w+YpV2E7mld0ulklX/TgVFEuMkeoleHJmkSiw+Tb6IdjlmcXjp+iKnm+Hho7NCYh
NAgyX2Z5a/8MM4aNeb+3Dfn58QivcIcpUbR45lyEorfLxm+S9gE0MnlMbnPR9A5x
u9BrEsEOpHG5XbQPpdWECDIEVUdaUryHseUa5hapOFlRmNqJ+QZ+A6QKM/tnfwDR
DtAt5nSGkOtBTz8M4AMeDjBUNKSzWU4vRC2DBEzu/kjIE/NSYoV4gzg7ycfFsyjb
vycSfzE4BR+9A+q2bJSj6jSO96gFqQKDBbEhxyl7v5DleeQQrAFOJiTgv0EB8PGh
Whq8TYmjbgKBO4Tgm0gcLpdF8sUNUPP1HNr+3xI3zHMFew2/PAStuyrDvYrkoD7z
SshXCYJ5VvZwmhSHpu1gzg2AjGRHXfNRipG8mMxcv+ekvQmEBhj3c3R0zu8sS8JH
yUAd+4iJpn9TWn6z9kYcKFGx/2OPieSK3EfuOsZ+apACuz4hXsEirpNF/nCr+cIw
7kkybjjP8nfRvcr01Zj4vXBJoTCgSChHlaQ95OXc7plIKOcW+8TAeW/3ty/HVtDL
yvXehYmoz5GAUdSNj5WeJmzGiAfjNNUkw10Bty7Roc1lackGKXS5U/4NbOpGrrk8
yAXi9ejQS98gXSIlcHapNUHah0xWKs4VRNeoR0Tibt+YUYfbGKjhL/aE73jXOHK+
55bvBk4H5O1qnv//NTduVRCzOsRVuJSGdh9Fsw5+IEF43K/djONYl93zJzYINnPO
8bqWBFfEmjyCG5zmtZ4ZBnTAzKwbHb5zq6/Jl9B86pRtiZDqQcAgKJmX2jegltfr
bzi5ZqH3lkkvf7ah6nZ2odi4IJpp3XY0uUs1VMTTRZQw/jWsVPbQnBjw/WD0okkI
fPUsy2KfTfUb+S3SfDBXfQzX72uKDTXvTHCes+HOzYIe4188X1O7s+2p1WA0Dwop
28HTvLsScnqtePsKo3QQwvSopnL+b7aUXh0PCxDTIUVVxq3wZrBAWvMqjPOkwUah
OPuF/GWQXv/5bi0DYxR742PcrrfK+rCYfOvvE8IUiGb0A7LlIHgN+u2ACdlUHck0
dvIKOCIJTKTVKimi4mKmBQ2qyBzqUU40xoIF8tROSNuw6I+S0RMo9XSBah2GkWUf
4Mw7Db3jMflayGTeP5QiR9l+9itIA40BOvkbsMcIH/pM3DVIHBAoHIHw1vnjApKC
ubk3HLdouUIyggoaoJD66gLVO5XrYi2X9HtZYHCuNd8PtBhLIqtmtZZn3eGrIHIf
RrBRQ4h4jmz/Th+4Ns5pduHBAfPB155cWVAyVzRZUHDZUWgztRr83Ls5IOKhfKaW
N6oV+Sy7GtWRGOJ0cwai7MhWsypc1it8BYbFsoIIuBKGodvVFjw7GOT24KNywLQw
sF+BrolQjletIiaBdO6szLiwpsmUI6RGc61c8gBAL9udpaVNWsuW1ckSU4JQ3GAL
+/7hOwQbpha78rnFN9DjSsl9UhmG8+6DLvqZt++lWyP0oOHsKaG1WGE8smtpXxnL
pr3YyumzjcQdgd5kzumGc/YqI4mgjVMI5WaW2npI705/VyCYYGwfeYqtHo5QrF7d
T9sAL/2bqgLZwfra2ozYMcZmRkfHHPSlgTNb5r2Cp3UOI7cGfKvKlQJ2Nn9e4uKl
Q3AdMztsKM0+UOW8zWGPmFKkJQRVDDOz0Hn4B5bFmBz3pyv7byUa4xL+Hwza01lU
+5oCC6CoeurGdgaOm/X2qIHHBQUhBwDwDKOghsey3Nk1gIPfS0rO2v/JUTaYYu2/
TsxFN35odKrh4SFwhelM11ORUy1N77ESfyHViT9Eqczy5IyvqZjCCy/3MQPc0K65
crw/X6wPU8mGD9Dwua0Qnf/pJp1v8ePQIldV3PtRDOT0WM/H3D6gPLp2/WpPFspj
oUs2D3CLHK9hAjUR/9TqOP4PKDK7RU6ADZA1Fzf2FYMrdeMhbn/IZvSUa+tvRP8G
PbvTE7PCG/dTQUxKSi1Tbh0D+sJJMOAprAYeijgpdmm52diKJi0WNEB7B2Q+wgal
1fasEG7Htl9N2X5qXOOFlGV05G+EZr9B6JxHWwqx6qyaguVbEoiTcwIcWtZNkQae
KSCNwIWHZHw8QA9Ipg5Z5EvOMUr0NSQH5pV7RC4PDzZV8o18Pp42aufZDffPkyaF
E03UI+zbaB4GojaxtnOq4LfsuuKsnB29a1h/VW2utMyiwOoxJIAJGIUXK68SYhj1
5yzXfINonI7XybhMPeNUR4o9Pqi2Hl4Ibbq590BaD1LAhFpMwOnaE6eMOhAZmKLb
PTriwH1uuJ/ROMzx3kgwqGj6flLX3NQgLGYpn618WGu4gVJjBsh+X8ZD8n0VSW9W
91q7OngysSXa6PaaSyZ+xUHdYvoPNHjI2r0Ix98X+WKnGVoHMyswrrGabjeAKmwp
drjk5dJrTHBLkLUdsiAPVgiDcM6O2QslDH6sJpSYQzPtSYKMbm3xZF70QL6WmqBh
4DSU6siSgUUJPR/XxxkkWJwAngSivPs9l5x415LSgI/QBD0cltDEc0RJIpk7keqZ
rTxxAJk375VrsrSXzGsbxT1AO7t7cy9wN2wrnchaqa7ac3fYGgwRvcJxeO5fPw9H
GQImZ2E7EkRmyDryjq6n7nud1ZO4FSzkJyuMPiL6JcCNvkAd/tF+w8AO0iYr2P8M
D3gTpKW8iZow0pU7AjJh2iV48qoRpUBbaSzv1YFCswN6nzV0qnDoOMQtVNdEQVP9
NVe80UXeIW2jHqYlthoxjxVKvnnnQe+jqqsc7FbAQDdVVKOZC8siHUYixp51crU+
hRff/wvZdchRBVFfDwS9ch2MdQTrUAuT242AmSwC6goZXugdTVZrH0VGINn/c2zu
BPbaoxDuOe8lXFQQj59TNqv4EYELEZ0ceqT32GGKcOBhkmVfpv4pNFLzsJsoPafO
2RXB9Dp7cqvZTaH7vKtzINC5MGIO2WNpAC0B35WFB9iKmULlaBaaSI9Hgb7w0s+R
xcpvZ9/o35r6Bc2p/ixNtzIbgyi7Zb0h3KtNFKzSDLQJ+B4QbMkRLBxW3mxrROfh
Hb5XwuoJUhxjco6mi9GhbN4t1tIIyyp2aALVcZGRmJ2RRqmphnunP1LC1rQDHvx3
HjxIioD4xktUhs7S1vTQgE75KeMimxZTALlaUAwK2eRsU+4ZcIvXlbY9TOMEcmBC
WW3mkhrSxhNxloUFJq/wRK14EvytVr/EP3jQhbqF5QrCHOYsm/ssV2GGAjzJ7/H5
Tceb+KwXqbSjM87xYCHuH5Hl8slw5j4gJuYhwa1XRFnZUL54ZzopFLkbPMEILVNU
364u6DHQa82lhV+WQJMG36XSQS9DpXeAysg9NBBYFi2RzamZVL/CnoKDSSPlQhy+
M9rM4W2cHApUJMZ4xkTjYHhvJHzzmi1ZI5tCLXGDksdQ0pNHvPu8Msx4noHS1Mce
GGkyHdqeohA/atQiv2s56ybJEmGMQDaGn5Ugx0/jyB0F3cT63FYe11O8x/cnFcT9
bWhTqVBbxrekLKkI60iUt7uzMq0A+cyMAsbodobPYEsctLNTChWX8SYhrwuVdf2q
MWWeCdmUBj89Z1HM5tPxMAGd0hiZ/g26ZbYYv3P0n7jQpX9yH7XTQbfic7QN4+DF
cfrfUTUssnh+0HFvQ6JFaUv/8/WmHDXGmO2sIWl439dWVIIxYFi1Bt7h7DnGBTu7
0qL0Q1E8EHq1CsAYZgsX2AjDf6cozRcgxmJQopz+GpgTKZDy2dTrtSues2iJHL/h
CiuljU1Tj00vYjXEsAT3ysFz41/kovXLBcdlOvXdSVXSPz5k50aY1WCeEscR2juX
IWVDiIXiMrpB91ZVXh1NDaZjLOUp/XOCGC16pRxuVN3NGiilSbmTDYcdAgO/AlOs
ItAOZkTixvU9vIdvIYF86iarf1mYxCiBTVNRk6G4DqSKnGmtJZeO3ZFgvJvtYaPs
MJK9+/r9IPeumhEpvJJ6h+i/gWXSA67pZ0DX1gCwRge8Hq/UdbG4oowPwvdil36g
7GTEVvcXx5lykLqoez9fwEOeGmruB16j14ezr15SnHERtTewfLgYovaAexAlIA2D
gtoau7pf88SDzDDRhboph00i1FvtXLml3PjiGqKQ2TMNcZYGgBg/wZtt1y0zFjv8
heYlsbU0F84doH6I4WPt2+5ntfFrk5Mwn7Tsyzq1jD0Z8tuUma6dfx/M/9mF66UM
f3r/zMkDKNJ+ZRHWJDjYkWXew5n2CMcsU1eKVTue2bNgnjUYl4o/UiKAHjrqeCMf
q2VAw/MF4Eo0e4UP+Tf5xdNQSHtepl/MVia4Pa2gWH80HEI0stcnCkjbzWLHBbAw
Lsu7ngxLYYumb2mz5b86v/ktUMZO/zO+apKZvVNN1GCIvtmrACGEy9FFm3Y6dduZ
4NiXOtyEs7SvtLxRBJrMeaclCMmhqKr65HfmAYxKvTAb2e7enEtyCQJpPPhLz/NI
lOBEnxzHKJK9P8uKsIgXtjzWioibiri49iBWqc+v/68GLThiX+PBz2jPfi0b+JNi
y0tYQvV2W/3ogTPfE8ux+5YVfH4G3w7Lb1tERjP4IziYf00wXBSLIgSm9YECEWS8
c5u3Oo44d83k+PNaoCSWwVxqBuJHftGYMHKeY4sDUK9ELYV+gOOr+HttRjC4vn9R
zbClzwpXIRvAwRTYthOCSHFb9caqyQFAK12KxphXFMG6q6xA68VTw8ahxHzO02Cm
gb4xeL9+s1nTa19rwTiNfBMO87FPD7s9vrCD7eq6yKjghjkwd01JABn4Nkw/SCf1
k7Zg6tNKSY4wxo4W5gPZLkT8/KqFwSdTaxhYM5y811xYb1soUUG1X52UQCKvlPIq
KGF6h4mAEXH/y7FUdjonSZAbD335j9vL7PJzW1GTKTu5VXsNaeX/wTwaeSDxMUkp
Zo7JzMemn7iSKPb5LMDw615A0jolXpDcyntGQIZQkvOCxLGKTglVG/Q1M7RfkymE
pK8jHLqxsI2+/lGC7NqtdWqvE5QW+ILZ+iRpfCuqAND4sf35Lwf71OgZA8H4XTTK
t0QdfIlkjNFnvqknHCcbfq9Yr4AeIjFQlYjT8D4RsuUbyeec2yy0ZKZRRNp7CSLZ
zhHeNsX7ERxk1539cjoMsfQCrFEcaPI25QjLRic0dRaf1yv9lO2SF1jnX4Ixqtoo
DXAUUexN3vaqax9jHNLBvRoUmAs3JIYoUgWOgLPYhuEcI8exhK6tttcuo8UeCrQc
+3J9dUIaOWUrnIrZ2sID2eLXNorUuEYT4o0Ukzapo1EfZeZoDXoZ+R8IQBVyYT72
TBo66JddduV98JmIodUAjCfI0sK13vcZ1YECvTKlYhlYjKNGpdRDc/0xV7ncmSaV
ue0hj++u4WJ5J9O6wOCpw7YUdhwTbh1b47soq3iouHK0HCUuqEFY/hUwpCAsSGMU
1VPUl0VXmSpvTrY8pUS1/fim+6nQvdUbkDs8SYwfOFJERaJNcandDiNu4gOZZFGV
n0HHlcHy7yZl5uewQ8Nyc8FgccSq1lHkBR5HEjkbxib5bUNDz/HDLouXcGILbDhL
iKoeJn0+WWGXtmgtT3bIvrkbVmg9pU+NNGOcfREI8j0K+d7maMilIHhbv6cZp3mh
K4Zcwab2wqB3OujKZRRJBnG7b5YSqYecVi8pV+GQah4KFjop2afxC1FsC2kfQYwI
nq5ZjNiDSzpzZI6r8UJ6gE5oXIMU3deQGj2YKB3BXNKE8FXpsSKuTW0jQ5a0F5rP
QW9Hn/zO3w46kmHOg5dnbp+ODpqyE9Yp54NNmNBW8Lwm+bs/Y+6dy8+yU5SGN3IC
q3aoG+i5tbpScnHtXkvLf7NTGUuDHYBrHIYjLQr0dArAC4TXBmLH6kzDx0LZNpXB
ECzbNllPLDzKnSutcwIkWqrIUl8AILFAZGVB7lYz9VOkwsh4v0p6dnP4X9LicHoN
/oCHtP/2Cjs5CifXcmDbO1Fp7ZCmmzVOBpyYD3+goTlxlBFDzawbVWNlAkKp6ujc
NP8QqP6E8GU0wZK7L7rtQpEtPiiUjGnJ++wcaZMSYnILybwHMGXhVRBbz8QE8cB9
uerd7f4LEhbsb8Sr/gjd/Fkob/Kni07gLiOxNIYF9GlhyuH2NGQes2Bu4ws4IN0Y
EUl//j03js38zjF8Ndkpu0yXpqqIFWB1izpSmbwfSUQrhGnGkqQ+DJST2GVpgpX2
mN3+rgUiZsxLos8QnQb53HELD5vwDwlygG4zLyZ3gQhBl9s+ENPU7yBGg6exhmFk
uYoKwsSEWYiw4vUHIFHHkV6gXHxqdti6sqoARQ6WStAzn07nfNlB3P9teNGuS9ap
ljtWOTma33AMG5vrAd7ofLFT07zoOOoif/ui9TfXwNNE6lrMQGRhhr4FpHpLHicc
bpZa7qg4IM3zcv2aY+JlVtuNTFcYaHQlt/FzxunWESveZ2yzYe8FP6mpJHZG7dz6
XGng7s88+/la1Px/DDK6B9G8pUSS3Hzb1Y7q2mjniHrUfmKlZjRHSNh78y+u8Qk0
RA6mHFF/XwjiVs2qvMkA1fB32vP+NoeQPNL8QrSYPw4ZEXEkTsTMIiWZFLMyj8zW
YNrv0k26kH0hL/oXJgO1yaVvRVm7yfwEN/h1fk+ZlVbQ8wfREZhzW3OIrr27J06j
T3ZmNB3igs+WxKBHOrtsT1t9f8G9jBxNhScqT2YH4p21dXe7Q9HSNqvExJR6NlOz
XmHtrgMknuE4I/vQDTWnUXqRHZsq8U4v2Uht9WhxCNfiCy7BOYohO/iWwKFhKyV2
2X/9rKdpsnYghKvElOr+uW3iWWaRnbv7HTs/0YJ4ytH5K/6e5r7TPAYsYQXxSMQQ
Le1hlz3HZ/r+M3cz/ShIMy7QOsPQ/AVD1/5voUPGrCy75DB9IJnSTS+bnlc7JhvO
D2fXWE1mZEzYxS+6JvWMPWOCCNVFADa3fqSJ/BJOivZ76NRmqiJU0R02Akj4kvPr
fg2hWqmlMuG4SfE8JeTPu/FafRoKlDS8OQ6iQCQ6DTlSlY1UpKGN6lZVbsCnfYcI
EJ/sgulIJx2hP/Ll9egL4wYFf/rm4+AkPRAgX+vdp3c/QIoah0VQycDGfv09skvE
5K70gonLaJE/4iZc/0wysqE28SjeYoqXTviRzQaArCGHslnE0df/KUyXDc17lM/N
4cyizduDldtYeC3y5zeIkQydTz7rExJOXluAtcETvDfFk+rjuziVkQtKeKm5pgGS
k1nIa2X7lBtupENH+dQ210BSfPoHyqW1s0fI6xxS5SnodaBic8HNRg/1GzU5HwkE
X8oATOI9N3XxRkoGsaNiCsVkGxTOwJj/YkyW1a8XQAxnxG4m/nOBSDXS91Rbf8cJ
yabnENprJw1vZv5KZqVyjbcJe/sYO69JZCBQ/iWfelbmovtuBuOVaj6kKEfI9psU
VA/mr2Tf2OfawARm4GbEXmdlct0NQEd1mKl+rDarf6BJK/3F70LE83vco0fAu4hv
b9Ow2sghsvovx8odHPdvwhFbw4YDhL6uQJDDvcvExfv5lAr66m6r/kOMNlUUk2Mj
K7rkdRk+XkCfR4OmpnjB8mmh4RdpR6CnQ1KsXa+u4ib3bC00FE3/N+BezxEhnfqX
XM7r5c18vcvQilPrrJXXfRbBFmQq+SjWweC9yabGhLO9FNhzmHougwcqQUf8Uvsc
jUJjb4K2Gv9hEnjEm4eemOGSPD2pz6KeMLojoYQrOxDWrAazoMGVwjnzl8tUrNG9
iZRGQ9zpw6nkPaeM7KsL66Dw8zVwnLmlk7CKTP/ZGZKi5VoocGpZ9toQaBrsmbMz
q1Z5Y0j3RMeFwcvcmrFC8nDMKFgltEjFzcCw0yaylf4VwuCBBq+a5uOHK7hwd7ki
edqVZtmzjQs7B2EpFPV6uc9X6nr7vyovidj4uTKYbdQ+paSPHyGS7HwY9fNs0RGi
9rBgxhhSbDZhalJZ6XX7qfKjwhoP/K5ONugxurC20zsgmHWgg1bfmYX/fCo5wxoI
v6AImSUvUpk0kbsMz+3BKNWbqyrbTwNiYwHOwTAiLK8qcTQENyGLU8hnlRt65k86
nWl46UQsFKa76WAHQyYk9Rvt5Q7a1fen+v+tc0uWLUcwiyzYdDfuWMRF8Y4h6cCq
wnUigcMneaK49hFS/gAXWbrwcvXHzq/hg3dPTXPJphEjty2Gwcg1/5GMvJzqL8lr
A1bRXyHHpGCpAAfWzJCvzNdBOzfl65R7Lxg0diOTwl6c3xnKjSNSJiI6YSRdB/kg
3TDkzX8OQMnrCK78Rs6DZRsxvhNoxzuMp6rCkn/D/w1btDHJAjFDPCinukxIXssd
pZ/CWJfe/t3LJVf3vDNnlEcyav0xVGGxYCw1TBTvX3EwK2TtfKqKs820sYGUDJ2S
iK2HIQOHgg3NUTBIaeDRDkCluijZB7TWxzZIR2W5t5QaQcXi20SL/SsKIVp5gbi8
i9rFhF6gp9DjP26bsOEMbyikrCSd0+pwd0VZnzyiuPPvx4PW76xfyLEsSFVfPQkw
2RKBFRaPTjfe5DD01/XMvm3iOmuwjO8xlYbEWgyZMvbEwtE6OpjFGKgResA5U3Od
aL9K4gFPTkNaPq566rrD4+vT1M/zd78XlqzDz8vbyMTTq0tbjSwk9CHMxSE+RHfu
is5vfcceJSfBZ95Wu3SJVLyADblkHKa+ddZZk5nIpPv/6QG1fuIyfJuL9L0s1dH1
9vVbJ+G2J8PGFUzHy23ytWAsZn3bXf5DhrSYKT4PpcO2bBD96vbf5CmmaKH2ZItM
T+gzPztqtMM1KhpZdCDe+NBy94BFiOPyye8blRoQ2vIi+wedF+wbDQrHYY8pSBRf
B+97TmFy+qyXkP9FnTbctTrc8GKNlOTnIH3oNyU0ANd0VOt+iMrUbzhh9y834NZt
dqG/BsfCnreoK0TJKaRFYW5Ydm8CLppet80LWPwh5UDMfsGvkAWts6NJs5kcfOF4
EWOGJ50av9OKOhE7+KZq1UJ6ghQm2JdPLNPEhZK+f7fK/829KR01+eY8xfNhXghi
ECXYnU/KgV1gIrCCrs02e5I83SixMqP8+sjejSqJHOAmxSgV85qhOqmEsmhlQPBT
PjN3LC+3OLZQ4ZxviueDrsWN1cvUv5zBoOcP579RzgxkVjmCbfM2J8SxLqImtTnR
2Uvdbf9gcMXf7p5bDURoTmkkOaZbOpHlHcsEJ5VaBctPDge1MSDSI/AZQ6jgb1fI
ydf3NKXf54t1g9bjb6gaboaWI7jlfZmqhEkM1gP26RiDtGjHxdD8QeKcc7fv9Fnd
9NzWjGFU2ba1n+sSTt3CrD4+bjvmf48KrjumD14pustt9vf5NFW0qRt92stdC/zs
DrqE7HmNqET3908Fm3QeiuM1g5U6j0ORB51GU2HApaLa0l8VwVSnceoDSYMpzfzD
02CCkI0X+lwPoKzJgs7+mh3VTHMrmpdCJVafKcTTYuGCJKRItxo50e7aPhVSfShD
94q12gLAIyCl4mqgnUKS3Ee9ka4cTi/9FWlNjlANOyxb/XkbC3nM1pnSe1h8NO6Z
1AElLT1FWAT728nUsvnen52aiIt/IJcaquJ2AeOhzLlV/KA9XzBDsegWLLr+ysfn
kAJpEoP+6tWH1rrtmpI+nwSjDwkFR1nnTZYg2QtweLayX6CbTVkPS+KVKv2ot2Me
CCHrvbSYCZOgrPH5h9OcdLgcC8jjMFw684M0IM76NHT+yVYucPztSW/mk3BXh3br
xdfiffr0zDLQA6rQfVtqczWeTR/BWUsDIv0uZvDYrls98/TN1IYrn9ELtqbziruU
YuoVQM4GUeUqvS2eZSHDTTiFZuigmgRuW7E5if5/+P7pCzWSCZBQiY41xWdpcAoI
gSOFqrcpd1rKDB9QLyBply/bDDh0BX59dOV4IpcorR6SZNBqjQUWorlf8hwpOVgC
qhBE/RTkoPutGOYRoh+bpuTu5K9UNh0UmqGORTDk8WwgZMnVJUvdvz8tj5EMJEIB
+W0cyyWA8+6WxyCErmexgtDy4t7CPWfYJ9/Dg1ZJXcrPztQxt7uLywxQ1VU2UzWe
TeFzwpROi8fHZLkpRDlfgyZsJMqu87GpjCbQNb0QpDKS2MpN4mFIP5ijXPv718VA
UkSZBSJXNn89sAa6Dd/lgCVYm2sMdJ/Z0uOORz8LJdYgmd8QUwXQrsHpJ/KmpwAU
tXNrwwH/pHJDNo7yW3WLGYmqTCrkpkwBKpw2kPbCvyBiQM+hBMOMud/t/xtTbFpm
bXWfBsmjHLAlO8zMLeUY9O5i/um78774wbaef9nypIlq6p47LlOsydV2Q3pOEwIG
x+MMBaDpXhIApzKv3gDs5dkmKfgFEEFoTvh5BMgg36S1gB6aJl4IJ6KzKzzFyuVG
xc9kTgghw5ELkHLvDw8JbtNzQM8eQzR/puhd2FTIVrrbi14ky5eIehRljtgTVE4s
8PGMe0THwJLzfPcOgjn0ahOsIlvCsSp11NiV1dn5FebZPqmmy21w8zUsGdIj8KRm
Ug2AG5N2j8SHKWViVc/VPNYtStzY/eX7oNMA8Iy9uIUDo/lDshSwIoIy0Lpv11Ad
Yw2N+sYNihMY9Rubz1WyZhtBP5SuAdh8RJvzeb46tr1SEocikDxPuzzeo+RPPXG6
V7WWSLrNppR2KveBKCGFRbnJ2hN+G8UaVD5gDjw4cxf0+rlR0Ya1t4bwkFjioAgd
Ha7NtEwr/uDAEb1qRvPiStUFzaCJTwK11uNd+hucthJRIHdwaMIqgg6pb7ITfrJe
o0RxJThVeHEGY3bw3lrBoYjIW/MI7f/yum2FdttMqu8RRfUj04Jrkk/LyVMh+lpk
mQ7AZfH3W5l69ShzyuoATJV+p2e5LkpklwFXua7FhRIoq4P7/dzaTZv8R2TaZSTC
jJp0ihIEMsAzvaLl653JoHde2bL5sGH3JGD6N5XCeXs4BzVvyP0yVm5GvvEpyjnQ
cjpvy/mct2oGUM9JigqpR5ZpMXHBDE9lnD8GcxdqK65HPF+tuNzseDmlWodqmxhW
SuH6PMo6bNngICiegvYsnBPXDHQiycpF9d+EzRFoAonMGDscP1+CpCui8xnd0ZpD
yqWsTr58bwebtvZKO7F2c034Pu6rotNmoyHNzbBkT2855PxgqMCjBpLmK/LxEyjF
MyUs7gKHnkUZ5BvpEzhFFV8mw0M82oKv9kZeKStwgN4Q+m5KdlhuE6A8sbOvQ1Op
IzPLRe5uvUuW67CyUHIN88c9Kl9Qh1Z40dhm9SK22QdJyXuuFh++LKzuBWRAvizH
O3gPVbfmz2Vz5DyWuZxTvvlSr5UnGTlntpg5enJoEN97ObGgyQrzo3XHwYFNBiJ9
iM8FVou44UXK8oOujOLdlIoQz+Ig9NNo16s9ACk3/NCFRGUyJqN0lnd+FAhc9vnI
i4a/0dG4eu2N0NigFNn9tdXWCYNRfiOlIVA71bQwYtzWBM51TLCAUUxTrPC0xqUy
rovd7csRZ3YliEd0O51f9FzsMTvphc9kheto8rncqDYcs8mH2sJJe21QUaAMpACi
qB1L8fAjFjRf4ErD9gwa2annmT86qg+qo0NsCL+ZdGcPPhWiiOMY9msV30t54INc
e/g5ZZt5EV6wNIL/+zfZCaPBpzVeHNKslJmaN2bcHK10QrTtB5PFp7RenExXb6ja
9d4CeuKOrtWY72mYEkfpxw3HSR/cBQGGHA7RXyXtT3pkycerE7iOMPwJ7ZVSnega
Oqvq1cYLKuKcPIvvyqUkix3xvZQyL1/NF+An7HbzHs4QznLSLdpnOXlpUP+0Df8/
WXpgJkBf7YtwM0q37zhDPCfYxgrPUK09fm7tQWYYk6WG71VW672lQ3qy4+YWBAl8
3NRQzMXClnS0rFZ+suCRtMFJPC39Jts5g4027e1yfQVkXEKXj8u2BTm+avYSx6Nj
TKfNGQHwWfXZ+jSiiGudoyuR3Pq7eyPtOZT1NnNAtk0enmP5hDs4+fA14zH47/2J
WwTCSAGqp5Ljv2l3+JYS4bhapEgT0b1+gODvHzBuet4soajMUYhZZBQcXMitbucx
GI1vWSQDYuH2E2S24/g83XpwdZYjt5udzvS9F1dPFsiYYcaM5btTUtJ1Ui6f63cb
UT9Jpme5NVRVVhR+QEzu1mDzEh8n3FosqeedCMJ8f94k9MFIGDhPJZtZisWLGrNV
LyECfHAylY6NpXuH0vGUEtLIjc2PJhBzERR7JCX90iozgkJkSGr7arwEXIqKulSF
m5oz/lz5NGAQJ5TvXa/b5XfJi/3JR2BJJS6lGTgibFOjCmSnoLiw2QrkFZNnK97J
3Khat8ZfBT6ql2P6awjD0c2mRBfqqdqU+TW/qfo5ABlxsPFE13NsG7d1XC+h2a0x
vTeprm2PW4WgETZFgtMDHiOoQ6+fB0HZm2E65s5ud9AESY+SG9A0D8JQ3A/abSb5
9R/wuHNkNDzPdqmdE54cgCJaFEsr/NURDdPAwCwAsvbXAwc5eA1x+gDqLqM84i/F
n0XqNA5yk5+DXYL6sjR5rVS69Uhf8HNfgnkO4g8HZhkuuQmirvodPqvTFBxwnzh5
cuwTFfmJRiLyX7Jsl4vfSwFACvwJ9QvUGgseo4lhl8BHias3t56x7gtdC9OM5uuL
3tr2v27jhc37n+0vb6XySD4p326J7GfVgiYTxSSIBDLcJgSaDBLJpwu0fm5GTai8
D/Ec0iPqK4sgDfOgGNmnQebSvGDbFwLfi5fFw8EXdgxAXEr6Ebx+tC7O3DJSJdqh
n0M84JsbPh2LK77hZvv/BNqmUqpheiuiKO4gr3GHTCyPV+B2uEk2CyZ3uzTlV75C
Ar3nbf0B2WQFsPdH12Ydxq7DjYrM1dNt6NDtSEiRKar64z0d4r3cLzv8JbqsNK7Z
fK1LYrQn56JJt95y8Cbw+UBjImFUWzrKtb+mreMlkiM6mXzNWpO5wbuPCbxRpDCG
OxuB0GtK/57SrvqYcEW8oI/QM/Uh2V4sp9k/doVm3VlgsQnxCBd0I40gv29zFzly
ZGAq/J4i2q4gXYvXxslIWvt8/8eMnv8Dj3CZu8gr587xcyUw39OXH7WxSY7KDaPb
N+x5Rugb8Kg4v6jDGdfHqDlid8MUZuADc6GhQNA0JkMLK9jCTRPH4/lYraY3ASY7
GN2vvtP8UVStk8kVRg7i3Ifxs/HRUDLkPIgLldrfX3hbGomDSn68a3OxhaEyvLvg
NNRzpOhyBkcShApNdoqVA3hOz3naOsHToTPKMuDM88k1UUwEQrW+RprHLBJhAd8D
VaungBRPRvdNZvaDJjFCZvPHy5cBu5SJABWxb/jsAJ//3Z4WRaNh+n/BTHM8V4B2
g4E8uEgjqHWy4fI9W0ixmn1Y0/+hCHXLeuMRr1C1/QnUCNW14oia1Vw8xVlofX1S
WNZ9nOdoB1mh1NGqDwZf+pbe2zZBFGqUdZ0y4krBpKH25bu8uKfzgFsLiqlCW55O
tXN7AOhIdxyXztVHGLx5RVm+OrY8EYQKOzlMJyfDeGyBqNUKytlg7IQ6vH8LjHG5
znoN+EJ8fBngRdZBR9xyXXHp7yXjcKR1s0z/IyWLbib82daKsmdgAiNHg9sAAEUM
RhyYrbqG31WyYoDAmT4f45PZtzV/qkoc+c+/mvbB8RDvnm9gIRYYi3Gqu6nUfqUd
+EtX6xUMc+2zbJDtbRPfygwdAIWzhHuLdiZybzv/PPstKqxzaj9fcYPrBzcbT4Yq
UxIB2B3fq/msUYxYiT/sVzRE0JlLPPqSUAXY+18eWaLhsKD/1N03g7CUXTUGsxmO
Zfw8PNCatQcGLffg/2leoCTe9jmpOfti3Hpxiyp4eJnS4GfNhvP3e1yb3u6xYzC7
WIJyk6pXVydciW9sSw9vH7hhCO5Hnr6dfRe/L9M/HG9zQ9KQnnahsaJmdX0mJnOw
NBq+IEax2QljfNhthZ3XtVvA3YWRZXaRFk4jcs0hlj2GUsGAQDROn/6usM4XGBkY
NohwS/YC7dIFOqG7Jn7vhnay5YlilhyF0oROgTFepT7V17rCrRCury29EDwolho7
OjmTuj/1KM/gGnYFDcEuJO9I2Cxx2Ha+fk1ezBnplT+i3TD/yZ1Sse8GK7FEImzo
AMc4aVgSGlOLihwDiGu+I4c0eWJ8DWgupSF50hpIgZz1VILeH4ttv70b92hKb6vJ
LX/iEPg5RlQgp7nl2F9Fb7M7mjA8op3ixYjJHTz+GXkarazm83EDULXw74qoSK04
SSDosgx2tKntqZSe81UnNHBY5vda4pzd3Fm/UlV+VhMokpcG4JpGXOclNwv4Eg14
e3SB60ucZxylDsloXeILkxg1buO5ktXHMeogLNPZ8F4rKV/JcBu3VyJCD4C5aY+c
PTqzhdqID9pMDGZByEk9D8XrU6Hc2qiJw7YlLLGHw1bCMLa0XR2Ur2fmiuNtrQbn
PfEDCno8fA2T6ASw1VhgJHhryIZVTTz0D0Fk+RMk3Uv453m7CE6GpPFF5Ls1RFXB
vtU3JHpKkK9YIvrdGow0HV4kAyCnPJl0XgMJLyv1+0scgRpEnkFa5U8Rhc8iOcC9
5cs7ojQqqrtkCl1xQUEeQUoHrJKua+4sjXBQEHrNmP7DE6UCika3T4hJMR8HTYbt
5EhifSVKQJ6lW9TI3xK4nRK2ONys2EXyNHC+r96fzOvfFeA5oFXXIUD2fNgmBhCf
lDqIQJzxalnhtvHluL1HTInit4nr4OcYmwXX2gSjcI/4Sp+5eIDM1Z74GFs97w4G
+qfD9kQoAhSgCyPJm3ZbSAE/Yo1uOOwOwIVWbj7YsbQQEbM4pQU0CUU8ASu3WViT
fCz0euKvqZNrFOiInZGS+s4o1b8/zx0oWI3QVMT/U8G/zdTNIHcgMWhWJPG4snsn
R7jzZ6XcYimHCmtIO7ZOj/BAxO7zLjChNiE/5hQ/hKvEZ2xQ2vr8FPu0uPjhJgqY
cb5zbPefJsCQ5lFa+DMFY4LHekBE9xxjlsg+BDsVmdpwzt5SReooYM6Vx/Er4Q1A
PzZTDMJQIypudX7oJ4QOK5LtGjgtjRhOMZESfywF/3+BmPEPbVBt6pnk8Lpuutib
jkkvygw+En5VzZKkTvqhYEhardngKorsstE/UltBhw/uejSyFzTPKEb+FnQ6b/6m
WARgUhIndi6a6coRsT6yAuOlvvw0mG2+xHOCfzCdpz6vLvYTu9n5LjfNxYqsk8bf
Dg7O72UgUf3a0cdTcKSB4lGbBOnB/U9oVvBXzhumC5JqVD86HyNxjjGcAhuBPzVP
bgQ606VVGvluayE/E3w+lGR6YObIRY+jnQG5oUTjNBYSefA0HOOrzbaGrzF73bb7
j2oyXwwQZh1km3UFK8FxJKKWYcy2xmUsadbKxU7e/Q6/H2k1GrRJtfJbc2bct4HA
5k0gsFn/1/N0xg73FEam29wa5WhEp+wZwuM01idBvPtiys6UoDEd3ZFE/572R+tj
mkOFx8xmWGc9ReaVJCxR6GIekXLWvdpT6AZaguIoRdqUFv8k5YqnCpSMUGil8Iug
1RviTqSr73xd2j8iP31nzHqLWe2yvENouvguoKb2ytuAOk0zdSwjHHRfF23sQ/Hk
jzWFQuEaFYFrJAV5PKxFdS5pygivBu6PkbwMG5o7fVcOeQSshmW7bb4agUTLiFw5
0qRg/l1wNIVzLRPigvd4aVpemjKT9hlb1Qdudr4tpiYXK4LhMhVVq/EeQv84gr6m
5vnniUctGWXqjw2WTqWSviaU4kcl/BZvku9WOQzFqfq+t6OqLJofTM1F8MsW0KV+
CnvYEtTIEUvt3KHSzi/6zRJyDs+1FXvFsxJWOEWJMx1OQyFyd1BhZw2m73SgVMjk
jgOKX1vppuICzstKnn1bqNKdbP7AFEVgLr01cRLDyscaC3VGh/IpG1ToDrdf0KjA
GM8eneiC9btCgRpM4Gl0EMd9V83MuSI14C8WM6j1WuJfCkJDp/k2gg02423Erpel
ihCpmPScNHAS1QUOFxIctVv5R2+bzUFDpJhpsNLZANGhxcYFweE0ONtnnO2QDefV
+BJQcn3hJNhI/TJWKkitpaeo7sfjXkHbfgHUsTWa/WNVJt9jDesdcqwj5estRc63
BkbPjo7eYeAG3AMge/6hREt/ZXOVTFvR2j9Ca87ibLokro4SM44Jko78bvSW68il
j3s43x+qTKaIY4BrPUZpm88DmPfeLywfpyrBI+SIxOiXDaY7p0rPVYPcMWlcWCA4
5ZXrIs/3QxBQ4UDLXG455eEGC9iW1ZHiOoBHvrBMm1XZvq93OHLpvjB+UQtgIO8F
4KKdjBXPq47D+YfGcSwrNzJMRbiDRLEPNNZCZ0JIE1AJJ4y7pFRKG+3j8q5NhyOH
EVHp5tNxGVzpAne4Zrzd10oi8v1iFHi8juSj+CyMpmeDbeCyLDUQ2lJVqXKegdFG
bobHU8p1i1cuCIfSHFwivUoPyMa4ZHY3JdShI2OtOyI/ONt92FOZLXAh4iyVE22i
KSBU08Ub7qk3C2nQ4YLfKNW+EVc2rgfunMG4RY2avSB8V0oqgN2hMPjJawNyBcl8
yN3Dt+PRFDDoP2/go+n4XhpfZmkA8gYzk23SHUQ6QwgYiBTA01qIkK363u5pxw45
wIhpgYFJJVUjtqwhTFLneTWICFkIPtfG46oS/bTsgd+jGZgJVyZRlqhDMDV2ROmZ
Kj4ehqX3Gz5n1iiwgKnn0j/8/hdSpAdB6yEuPWSx33pI44itCUkTxJ/FKaVU3qi9
a3SLSm9hYhhLrob8oGu0Nb4oKvFg25oT7acW3FmTJnlHaJU5BaD8KWapw/0CB4iX
tejZs4Gqmiw6EwiVvHec4uNUH8KrVktV82Dd+5TGo7TDD0l1r4kpH4OYlHNfqDy2
XODwpU0VXTxOquV2uEvj97SzwwYLcbKUM3++uVcwEUec8e4qAwXHq4dxrsEBN9YA
LEWVe6p2rRBz30k00Ys0OFNSWfJPi0z9kdLSDacKSYYzBB6WausiceAsdrnuVWc7
QlAfQIWUatwuA4cbTV12Hb0/4recDQAE/HfLnjpvuCwTvzQ8Rwzy9WaCN2iMcMFU
DRPCTunhXWen7l4ctkzCjnQjKQNhkmG41tvmKtoCEaOVs0hcMmU5tqJdo6WDEH00
8t7QfUer/M+5U2GcpS5+Eb4orktvlLOqSwXFbYyVBdsH1UHMaPzWd8ogXgYHehti
BkX+LVDZjEFX5BRHDphJyU+vNa2qv2gsM2f9TABc9Is/2umNNHGT3Sr6qylTfCZc
Ee4LCPXaHtkGCl8q2kKcu6t27oDxr+htdyGTpxIkGkfoGaDo45P5X1Lw36BgCOxw
oThxXLpwUd2yzNYOCsD/SiDiJ34f/IiH0n+E4KiSPmRDS0lj4Ea7GvBPM/V1giBv
FQS7KtXSOsOS1ca86NY7kUBlAgERKczulzZsWidI2fKeq37soz4jMRAQ9B44ZTrZ
JY9eN59tx0FSOZ3fgGPVsKjVrrivSYeA9/chpeeT+lN0Unq1/oavGugh3diFE4Sy
jlcRIuOl3dUN+0RaEstJfynqu9NNVbVIOoldUWlkoEwLVcAEHeIj1MGN2Pyh87qs
inirxFop7AdJgKRvEAIytRWvbnXUq4E7GUcEmmm9lhTBi0spG1aDmg7qHcFkPZMP
nZ7SS4X7FgZBd227NWW+iUzH3hpGJl9u4Qm5D7wHdV3tnytU/T4cRyricAyEhGZP
TmOVogAt/wqwLt+7nX8UEhIEAjD/TPNUjou1mfs/chCFSLuYAJ2iOQ2zBR3qZqt+
z/UI7JLFJdYMgts6Xj3yJTPn8B4iKIuETiJLu3NaJVuoJuKTxQbL74Ho+OrBmHDx
9J6ftoHA6JJGIxTCQygMHqqHcRSX9hxcwVTVA1JiTTcpY9qs5P5zyF1QW+KoGafP
AHFJ6ZYyxOntg5ZM/UOcBdOMRrL2GwZe4oHnndLR4arCI/qGa3Mx+cRO9tRcXXJx
Fcn6R/awvBOXI56Ir8KCqFrDFQG12P/Tduf6XtHjQlqu1b63wnAF7p+wIDM6rXCV
tfVLFB3ctAdZZ9o91jRFpyub8TeAV1ZWLOLcy4Vejd7D0/FIqNDFdnZUOYwHjB89
13yIg5HrqJNMu0Rto5NrukttZBoinLly8SIYIN2HP3EV2e9Dxli3nDTQAUn1m6jK
Gg1+NjeZfrNfPDTfMjLW8lg5C12FZnUz0abcfg/RRz/aJht1NgwQaFaBewOkzyZd
Vk+NxrLNSaGcMlY9TuDWGgoudYPKmPrt7rfuh6yC499huPFs2kWqIxUxXPSMsFFD
x97h42rvnsKYpSCtvCjUWPI+5Vjwol/IPCUVfUiEag1XctBvxEDuUkA5dG/TXXNF
a/nPc9c1ECabN4cP2VaNIPH4fKIzhDX2CQyaqzfsqbMhKDq0FVGy3+Ab9Ckt0fi+
eMlelR224h04yNSKUf3uLrIiTUgeWgcW8w8EjCvuItXBNjxYnOSymL8cSUiGV6Cj
JlllPXv5zUx9TffQ8bPdnSlDn6FPHTKGLGlnvroqq4PRjNcZ1Gw4RzO+nCsD+JR7
bTogjJJMWgeqp2vOxKuLnV0Niuz8y9mjihw8+LicZ9JvzRHJBpSBMfinZjM2g/h0
CXpJzU9TOuXZ5bFgfsXwtUM7bBEy+frImWc0SlsIZ1E2hyEvMrFMPPUW2tjUk/M8
/LgVjpNJ+3uDhuR49gZQz0lM3lxIxP2VVUkrAIOHTB0NXpI/0F+WSM1mXs5w7vFR
c03CpqLLTA/YVxxnEU9YN4dw938cPD2nur8TfXJwhjuJ7dUjuNW5oI9uEc4HaNxz
ypFqW0/cejR5iPnWlvBrVXMWWf71WhBXElFPxXREbAgx704HZqxjOYi6TSUGAB2Z
ehRcxYOy3+cfiiI6x8xAFeE/oFX0Bnfhnd1eaXH7ZelQayEn0WjUjPmDysDCKQk3
+0lbHSAsbgKYcXCAa6+brBaE/ATeATiVwke3vqIzZKoEz0xNxIkJK4714Aw33lFj
sX+nd1DdFM+ZWFAQW47IQOJW15H1kS3VVtjdbMS3Ki9/oIwPJXMI4w7u97tY05Br
XXPlHSa9MmMg0arEjQXyU844bYPJxMq8QLQTkE3zZKg3vR3ZFNmuMBoFIJlFKnOq
YqMhTRbRsFXfBZ3w8ec0AgK4EV7sK0K6VR/yu2dU35ZjgKbSqDaxsXpDC4tDrhq2
+j7gs1+grZmgIgr0iflHo/XUJ072p3su3xn+sSvZiN1vSctSOcybFU9X2UxICFde
8vUS+pQddOvdPOKLg69uwH8AU63AXexehBt32BF+4TFVwWy94xAjnOBEtSKCF2WX
/pz7RmZEcaTflw05e8y3WJxkzMfUz7rs8t+ZnKtkCzR8ZWT0tnBAXh5dwJPJwmDr
pac9uEBef5DhAi/rjFZmaH5dxOBp/CTSYMms8j4vFwsY5MWRBcmXC5dmlgkTlldD
gOqfrZ7uAZMJiAmeiABpDVxOaP8O9n9+EO3psSGH+np0QXe7LLzYd3powX39cO59
1ahS0BrewNaUPFMDphe8wVAh3BAuuENyn0KbrLTbwQOl/In2rawK9i6tegDXkYqG
cJNkcirsiF+02rb0qPVzC2br2gtCYU2xHpXjEQoTTxCFziikSbfvvJqdEcpyShCI
KUGZs+/RhABnd0OxKOLXknHGy4K3WrRTwh9Gx8+6l1kkG93vv7zuMhLATHkSrSa1
7ympG5A2BycWt6EqikYeDZUViFRJwBgJgcrf8eqi5uvSF2Z8ssR5mtAe3W/Rn6nR
ixJBcKll5PSzyt9j/XbJ63BAbzBJmbDRu3OzKG/U4jRo5G3tATrKIjnPL9TbtKC3
JYd1G+h2vCI6gP0jUPYvlefuS1HEcuifx4OGkEw3KtXNQ8fX4//455LRdELPZLMV
agUHV/neIjEsfxkRqoQNki40ZwxZUz4qHEdVf+3OihHgI0sp8S7rmTrB3oPXnLMV
avGKM+UorbkZo7/rCAiq+EYz6NFPrAUEGqOTWihJOPwzwKXgHK4RTINVLfZCembf
oPtpsBaITRsT4xgYTWKaiEzY8WD2evcKX8vYnDy/J6TXpfM8AXaL9knB1BGHN5BM
nLlVJhHHFoH9nbB8FHSHuKzlROuthPAhaDB2VMi91weYzP2+ODNySEIbfruG86gm
kG5bYGBZ8k9i54pLpClFRplTY2pAD0Amq2IzAFDu83SL6zOSexNTQK+g/MAFzaoh
Q+kiC++WwoT5K7rVtmJqsdBzXVBtX6wCI2s3tjv/1vmryN4J38j/bxmj1O0QdFYy
vZaGD8eyYyPtI6g5ubNlzPiXrY9M1A9EmbGPWkD5QncUQCq1CB6sLcfVwsdbG620
BXlNmEaWUph1MoX49UtcKJR70FIlFlgbcKtYHqJeZjdNffICTrTD1l9wqboT5IyE
0iY+pQjDGzZ1C9j2Hfn732FLCBPqlHvGRctMIRMIGOObk2FjGGrqEaa7jbpmZFHk
G57hpwjLLRt3RxACBlZ6R70fG/RSoCFGXOAX0uHsbLpde1SHCSJ2Aro+P3ers1dg
ZLlEs355DRAxAE+HmixQ+C5ICU2XmVwrFubvO0hKObNV+QXEoB6RPoRQvhk3hhxs
eJEs/3R9i6Ll6PTvF3Z0IB/Qlz/HS9PQSakWYV/ekXxoncjK7BFkNZYH1/sARf3V
UIbCWdzFg39Wi70OsE3ekVy6ycV9NX5hcLxBswvtPTIYXPV1uO/1rMip8H1mT2FM
188pC/N+8939/kFwtEjVxI/p7+mch7WUyQIvZQXDH1iOl341/FkgIiIyxf8Z4Zbk
jloLuqX26yRWZXXbkcw3hUBx7lMj+4ocWieClm8AS+K7q1K3gjDodfZr3gzMFbC/
csQSs74Y8x6F39nsFs5Fm/ydxTB53l6f+q9GxYThB4XzeHDd7it8shL2DT/8lNwn
gHcdPYoGmoY2U358IdNEHdk4I+XjUBCHTEprZ5CvqnLIbVKyaeAZM0ssoETiNUUb
StSI/LpoqoQjOQrpq1B5JuDHH5A/a45AyxCqh/EdHKAYIasY6m35NO2Nmuxl+N9E
moR/0TyPNcr2THXk1FXP7DHtzKkv/A3RawyOx+87xozMRyOYacBoAS+PXX7l88Mr
KZi9NY0RYn/wTVWRQhJf6X9Igp3rFZKmWhjrBCvNi19TMuTezCLr3qJVJTqP78UV
AS7L2mBw5U9eJ8p2DoA70yvwt+9UcxdYdIQl2akJAxM6De/4xi2ckmOjEPd4pA1k
SQznyagmvED1agfSrHDoQWh2lhhpcgu/jxgSytt9DWIq3zNeyY90JtTumvS3qBp1
RlqgdcX1RNnRUwRoamlImTFYvUO8yzlM0C9JiM9EoEx2utvs9lp7Z4I4aE+5pAub
0sxpLQexsjS+Rsfv/wTjODximFX+5iOUJmdZOShrVGac9bL1/SIC1xZRocY5+XAj
oyXbGAKQRx2GSp1XdpcQGsaKk1tfzGEeoFeEXbIQZhz4r/K5aT5vyOSkf/VP8gwa
Zf58j/0HPuSSZ+cc0K9IBzBqRRbEGfxdQgI+/kC3VxLFgwdNo66j8ydHmpcQCuQL
rddpNdS5ngOPl8yOOsxabS+7zpwAq7k2H6XJS/aVeeTCT7AE9D8Cmk3+sz32Q1+s
BfwfuNSU0vTdyYhNwwOl1nad7IlcgezpiO+EG0ClHULHZKFpe+G5jJoqd4ybRiC1
ac1/nnsw8LyhL2U2AlKPn0gxLRCaOKF0OPeucjT23ekMMJ7aoglVmdBnD/FzaELY
KeFeC1jq4wOHNReuaVkiM55e3r7zgg2bjQpYYoXfiZXEMcckXVp2TurV0arTViD0
YrAa8C+NNisHgVb5sTee23B4wzttC67YPZBg3P3BO6MJylC/ciZ42kFZ5X0plFhD
VF2bZExdUKQvh6EfDg3fFUlzcMty1O7bYI8IwAPC22eXnXh2lBbo5G9HaxhHgstv
SNCxSzA61GuvhRSq7jEYJJEy/2gZhKoXopPMh2rf/AdViL4ARWSd24NlcHfdRnm8
+G23jB/Ewhvm5qA0YEODK717h1mNaKC0YC4s0GC/bAd62CN0L3fhjbv7VitDVupl
ROxrBzwxgIrNIZ3ZeotWJRuDz02Qhw1TPQmTUcO0nVnThuvshgWR7giMyKlBKny8
WZ1oG8LbDbheTzwOyeyK5RmMa+XJ/P275RYGnY54jyS4Nsv+WqfBFRab9YU10QTr
IyfEwRaF1+rJjUxqM1qXyQB6VKLu2Nf1KueIUO7pl7buinr9RttHpPLOjHv5hmEJ
LyhjAElfx7KuTQ5GUFjjJYdvHo+8KVTSk2WDk2f0r/hKRiCDEnUnEbIPlSdXN9WD
kJz7m2Yk6LoVlSOQLGuSLMkWK9uIcNR1NeJts2gESf9hcOraAM44rPy295FGfHju
FFD6nwwY9OHds4olKN4251SYhnDAiGjC9owxzvyPQNAcWyQxSn9kBohBVoPv2aDX
IJPUrfEVe9J524fYNUmeSisaJBaNroWV/IvZbR1zKTRdkUw1cH3j7DPKeyNfSvCt
6jO9nka+lKDv5rfnk471lyiT+zkWxZjCpeM4c8KKoacMS5gDt3IAT8AE9fzhaDMe
oszFhn/GS3rtsBFLwvxd13WrSIg87nAWbds1Y1+ienApt96lE/JLgomfRJX5XQC3
YNgqkr57QNYzrdkh7E2PpI7qdupRJVgYgk+lqmRYXdoylNeTn0BSFDeNCa+qbPIa
PoutG77uZiLDvSPwmZ+FGtd40XANp4OAi3U1StAjTA4h586HKJElMu7DwI3hfoxb
A7jFIcmKcxD2+6L6lu/9TSks7Y7o2utFfTwGfbVOK4qs6Cyt6BbK6o1VgUukw3/8
880esIwwQch9r+jta1rEgV7k8IdysIC1tRKOQCgF+dr0fjSKn4wIG0jlEPXrbRFy
N8zvSuD3lk5WGno8Zm7Fdlw+gibK9s+seMGmvd+181STECfNnzVqWcI2mFG12qSC
sKnEom8HMTWuH1HAcUE2+Lj7mn8lqbIn0g+Bd4HkrfCMMLDiwWU3Kh3MWJf2ASJG
VulFKxG2xqugCH1UdICb0qchEwPA9v24npMDf9EoRPiMrEa7wZkwUxPleue2UhhB
n0iDkwhl24Aoz+ZsFZx/e2pzYceGYEQnVHT061oYcT9GIeEq4Qr/n6dBisl13s2P
5wQdXKmiOrbhItjITFdx6noXyMqULa2M6HXB1JPjZ7O1z6oQSg4C71HdF6yX+Lfy
QU/SQ/TW7d1HD7nse6yMCVGUVl4HvauLPJklTZisH1vowYG7Ti1coPYS4jIHP9i3
cHOtJZjOOIYWwmIdZmB2icaEmXbw1xQbGVTfTW1D5D3rTSew5ZBiF+A0DonNky5h
2374N4Tr4Jugp8KlM9/yi1CIdyPNaTbaun3/J7gTRN7ybgU5+nUFElUB85SX1IPb
dPNhRP3ZD+5Lw5LUyGZhoZi2MSZn+1mYY7kpEsJCuIOJIEfJy9ZbfnFIrIRDmduu
1V8OUTHXPssoX7beHM/R9xbZpGzJ0dWYskoIFujfBRAfI5BLhTO5GGylto6bd4UI
LyJPMEc7Weu1uCqxPmgzjOKbqxeQ79OpJUd6EDvPBAblJKDRc5xtqlqqlqAfkCjq
DqiGEIfrOEJie2Ol75BndbJnoYiakMD6vSSWClwAUXznAxY862H1NsOiI/GgerOe
a603A0nw4RgZQT7f19cfbf8sYCXwg3eFCbL5spnnJ8ts1bz/c80FTNi/S4E5hSAZ
nWuuQHYHWlOP+jizc0nniKSImEHoHsO2xDWfBoe4uS1FYHsV6z/1y6sfE/d/JWn/
GBWe7fUA93uvu5Rbp269sEJEHBifSbh0b/95vxHjQpkFPhl8wRzqIP14Glkkruxf
Mj6JGK5qd/czw+dkNp8mwEgACfltt4Kslsmb7akgBOtR0NZ7M6PqbdAsSteXFWNM
54ZfTpujyaTCsChPql8PQbwddBMr8npiAlkfD+L5Gu+8y44dsb8CCfx2AQ0eRDjk
YB0Wo4kSP5pLyePGYYHnOBLPB8/vuLW/PeKdLBcF7JSzCCkpr8c5POUI7KNThy5J
zMsFAXjTT4wUV9fnQ7rYVPc3jj17uEhOFPuVPjQs9oiHY8J+kAJpHgywdxbK88Bs
ioiEqY8E0Ye7gkcQmk71VmkqAoOLy/fTDm+HkpJ8TIDYVFR/vCapYoXKO5vFmzAF
lijj+PuUN3BOpcItwBPMh+WZaB8lyWyDDolbKb2i6txX5xAXkmFRquVVzvAWgA9A
dnHx2kjuTnhL5FVcZnYDmVIYgBiGjB8q57ExGdis62w/sCpeoceBqkE/Qclce0Kj
yYhP/+FIVR7BLz1sJiDRJn3O7X8j6USwjXKBKybtGgXdqJ3Z1gofoHXrI1zIpFwM
/vXT9NKwZbutog6UCfsgiGWCVF5Xyyr3o6iklN/NSzeDcFd8yd2yYXply5JCZk7K
NpqCTeh7770DuJ1msgq+ukBLD4iZdfCbLW4JKjtUeQQHpu5n0ALByWIwDOhdOVbj
9XJ4wgYNcaUt+2B5eoGP8VR1NaU65705si+FDT0Br6eOzpa7aCBZvega2eIHHeL2
Z6jx4zyFXdR0cBzV3xvo9HMo6giG9J+HXfNMVUjsxsvxo3dNvsWt5cudAO1obMWj
mGfy8VChWghIFGXp5Sy2AevbsyQ1nNRAYBrH00z1tDM+dH38tYiwdO3E0V5cIqAx
jNHlNgyKIjxe5Q8JwpoxwcbEtIG7uu2mXcl6f0r6OFBWDdSS3uQheqVS0UuApKZ5
jp7PoojMpY1zsiQytEnKUEvKlHzSvPg//DIEFniJ3obcbTJc6WSgSKlI7ehqzFzt
ApLwsamqAH2zcDJxcnkMkuYVeiSDceXq8iFOwklVFDKnYqeRfoxBe+bz2RlH1iuR
qWFVYOQJMMxP+DIWq+ASUVhCCgRSQipwWVDgaLtqRBt+1iQFIg5azII633MqagxJ
IjbFs7fedcgsqSU1RIJnUc/PvN2JhpJ1kkOEMclJL2MBjI+9yg2bZz1oR57Oq24Y
Xp4veCaCg7U8m1GEeXHS1hvFBY9CYSh6+8dbUPYerHlun1eTXSC7THKSL8Jj0aiZ
59Ld768Jj6b3ujdK2/ke11Cf3z3c9Zb/+05xdJpDbVUh/F/lGhSvqzTlnDZS9kkh
8i28SgvE9KDWdWa5Kc3dCFcTzyYbRQD/hulJsPBqadALt6XkzC5PusGpXTNDUFPe
xmg+f7LFU4QZoMuUygeSvI+zfv6QwJpkf7jpUM+d8IRdXU0A+qFOnZ0r0p3yJ3PV
hbTsEX/+9b0UQI0ENS/d13sbD4oF14EKrzz5ChETL7xrGBZujgQCPKFRMEmi4U7v
QxE/+1edM3mhg/H/QCyS1t3sk1Y6V8TSFvAqnbflmzXpHqStvfljZx6z8K+g4S80
YNeHgm9+CkJLWAhg0wvR2fwR2HSi0K7o4X0g3KUxpj244wUbdichhsrlQtHvgbcf
zNRPHpW/QjnX8sgmIr1YBMRTW9/BYddkyYHTn++G4jfNKNgxDCS18TmhR7rb8z/d
i9gkuoFokBSLc7s07VPBalT55+8OOD6T8jB/TOJIYhNqjYo6EF/+nbrdcBQooG0e
Q6Rfp5AGmdXWBX0CVkg/zSOjEkg3//eZJF8bBrMxiGQW1pCcDd91OgVX8RC3O/BV
2BGnHXRL6+wM+X0NHAvTBoWI013Wb4kyJAhzyU9WTRCms3fOLlAD9BxIh1whJnMx
o3DXPoiHMAgC1udwhKxD7Ox8hI8KUTYCm41KiCaEj3kk123TRQC6pa6Dm6p0AMQj
uHsDr9K7hPQGEhxLoLsM4Qhaad5w6oPHYzZ3ySQJmLZkL+/aXqRAc24MJIKj0WYu
7rkj/fnkY2wsfLKYP0H9Beaim1ZfiSu8e5UUX1ODTeKj4zdTwctpaPjMJ1ewFGDB
KHCoZEsqiE4REI5rGki38QkYmdl+T4oh2Trby7u7r4CEcH1E0fjG+ssUKMUY3JzG
vaowwS/sbQAaFYRWXaLXPN+On/mouGY8ZrOIU2Z1nqEaQBjyWmZnuKP1i4jvbzaY
v6XNEG/W+Gg/Piqg8U31lOe1nGThsk5xEV2r9hv9Ihjvhl02PjN4iTg2g8kfi3o/
WlS9BPa3M5rI4BETc4pgZ7TxPCLIqqmHbVJlCEvyn9VObKYv3aksFSAEqN+fNRpj
dkqgejYM/bnkpaY9nJ1NAl23Y7gb4Zl8jZjsuFR7U2qCSoe2Zyj9nLc1/SXlmKaP
WFlSfKZtzcrRLOOY21+JgXRP81fwa2SkgTKimLW4M6IMnp3N5QMNLBPjI4u2AcQa
opx1J7ujmdHEmw6ICLmE/PRj49kRtQqSW/7u1/N6kriHhWhSCWTb7TsTL92sxCG+
hhh+1il9DUMHjELSM5RHmAeGWwdk9pcRBDKRJesam5g1CKXXxkP3ftXyxVNOltVe
A6kRTWltQSACLKDV6ht4gXhtSzgO6WyniSIhFmz1A5w/7iQpKaNTTEZmf3UrzaW9
gAYS7ggwcu14JaIYEm12BNiopW8xSLFJYnE9Lx/bf40qWFE3HLJH2KapYEs98X0i
7mfxg77OJmYBHhwq3/K8wwV85/MlEqpZn3v5Vm71/Ok2ogLGa8oRF4Fr0DQALgtm
5mtzNu0nCIbOBQL9zedpkUtVb42c/WQoV4ZsqeY1tUufAtAEa8HrKXkV5EDvJmjF
iZzd2PljMYEsIf0jHxvjW3KHgiznMfM3uUYxWmRtchH9oypNFdcbxA88zx+T5iLP
aQRxE9wbiOdlb0tDBaojNtgPuTCIbBIOXVyZFy0PYllcBBvHIRpbmVpc+8nWiUHp
mbqL2YPTPdzpRgiWwZ1Yq8q5MV7FYTj9IxrTT2VlIfUqH5Ysqu1TZW08rZw2kSIx
lVozkWEIc/rDcOwSWvIfKnAIyby8AXqMF7FHPFFwcN+cCnkB4KuSSd0+lArLoc7c
M6FXuRBiTVrSBZ7OrWu0FlGeMil8XOQlVMvI/9BzrTy6Ovl7QOurWon8aZVhGhQ2
B3r9soOfLROU6PusdwP3HQS/XeW1hzlWAyS5ys3ongJofPWNhaI9UG5vN6rtIU9W
XOTjDwwRmiroGOWPJrkJTdUiByfTUI5CtyjWD8bUG5j+K2ljX+aRlso52DQYx+wl
DRlUcNV9d2h/YrJt97zRy4SBm/pYlXSBFDABZEJieEs2wKMdT/AO7DopcY3bhqfc
jfhGP66MB7qCRb/n7pZ1SqMUajdGl8ZV2lLmnw/h686yWqb+qRsrdY87j3tN7B/r
pnuaqT11JU/S0UE2gMtIXUEt+bRwRHbaUsvc73hsYPSA2nZ7JLlcFT5W+5iHiZeR
hFGNCbKM4fwbWLP0kmuSlWwy4Zo8b008hqdrP/hVitePuk2KmDHe+mh/Bmj2mRKn
jr6W8X+p6tTdi7Ob219Lj/I7noB1CMDwwyDcBLhzAl5uaCc/s8wL17/wGgr6MCaj
G1MR6FOpmBDilFS6v95FGzYruCNbzh4PLvO97Orys0xDkgcI1FTevj/vJ5xymWF5
yem/h/ez3KB3I+R6wM7QnCnDQyd1Sye6W88B5OjzG20eS8nvEuVChXYMPj/pL6u8
3nCeZCH0s1NaoqdT7ooKgnOrMBlUTFEFr7LBJ9s3lAOkjKpv+nBnH9MIDvcgAPEX
l95jl7OqeiMNFvK3S1zbC53fWDgxiXxJfpgMVmtI1EcOIIkBu7YktFUpyGSgyvY9
/V8HrI4dtyKphbhCzrG3o6d5TLNIC1PCdQ2C0c3xj5zg5UNLwx7w1QNX/k3TUgDp
KswF+BuVUvmkABoyAkvWvDgT9fjolS28lHnfH8wX/NCUIMatkQh6k9fbAKnzRzpx
0pfb79w8bPe9E1i/9ikCfuzcYw43cYii4mqMe8/ZDr8+SVLV31m1vZZoAWVF1Zm6
Ny0VRo5sm/+mZnndDwBDOOEokwZmUb5VAv3wtMEAeVkSW7TpKC/aQMMBGPGiK+So
1+FYzqOnKQYv4lR2QUtuzZ23THNy6NnWpwzHKyCokPU444bZMsTXg4aSyKfvtgMR
Vo8jd21wrTegCHBtx8zSGH51YFR1MF8D4zKzknMIJkPTc3bPSev+ujjcIpr7R+yO
9unL3kul1ZLmfOsQRIZSdmtaQd+6F/lTVRVIRS3+Kk4gwzyjzGRSWjscRjHRPe8G
xCB2PwuOel08oC7rPb9+r+bu0dIX2dz3CbIADbRcsdRtYYFg4LnBcK0tGvS8bDEC
CU+mOjtwF+JdAPltxEuvFSl51YC0/3+tLjDR79KbkAMckEdmPXSDZr2fi1JWfzSK
HLr4/MTTd9Qf9uVBRbCyu09s+uGGfZuwRnBTxifYsDb6woXK50he8v7TGu/pO0Ku
w+XmhScmLBzVgXq/XqCkpiW+V7kWCiaTLjTAe2c7khZ70UJRpwXO3EmH0KsqM7oh
LGoIOVECbBwUh5TvLZ9ov0EsDTXuJT3JMS0v3JDI9+nHkTWIPC33sydCargJXkne
0Fz7vSehNk63d1SOCGTgKdR3wu2Yv1GtKSeUjGnrD9zpAT+Tyger/WCwjO70+Ssf
lYKAVCwzskCaD3lSkdWpOQ4SM+glMnbYN3wZVwOboB9UpV5r7meAacek5ln5Eqyl
YCqU6iK87OlhoJmM4bPDoIJRsifpmaSshd87ZBffDrp4EueuiqAsfXB2zFnFX3K3
ZprJ6VJeg3DOAJjWAu6QMyabCroGXuUazk7ojSJoHXwZrWnmwDlOXceLFydYeNUd
0vYLeTVC15DfbdkwfJ5puIlYJo8yNvBUhm/bDBRzmSFsAQDD857vaMqMh1I9yDoE
eAPH1PQxpdhC7fk2nPlxyQj2Gj1KaXLwLBCaskQqP0l6Rt1GoqVyEZ+xC9vZ7DNF
SQky6iK8RUYbOjvU1G9B3C3mektPrLowHOZ0Sr1j4juKRbHtlYSp1CZUd4SqTwiD
ZyOGgrNCmEv0LVlbr/u29KfqWXYAwFLdGXQ/XVFhL6+2W50tbNRzwV5/gAq81rUi
lG8aWxRhXW7HJ42fjSie4NV0VwWdY4aYZjBuBZt2ag+pwi43Lxj9QeTg1Gm0jPOR
jCsa9/Or9/wdOFv1pTvI+8etiJlF5Cy/K6v1B7DhymkvT49wE3m91brG9Fcknp5m
FiqoW+rQItkqgmUsjX9bAmUhOT7ikMEPDuEYFBpi9Ta0co3dtnsT//5KiwLimR6C
HNSlzND8jCxRcrcB7aBEa7tQMkcahLIJaaFNZtHQgX/5Shm6QHd0w0GobP03VsSb
Q+qfT/oQOT8kgQTdgW13w1W4v8R8pXLi92lwSlOXJ0mFZAWmzvNN8kNplH23soFo
op4A5L5l6nf8YwS2xXXOYxoZYXV2tZss+Tdu4V5fAzsiUkqi/EEtdXeLMEQa0RbL
YdrwLDwuX+gJ7/N+QlEL894nRtgoWCLe1Izyly7jQaBbHkNbbMwpOXWzpOHqq19U
LZA7mJCaYcWPndnebxER0KiHcbR5MxMgZnBe6qZIG5I5Z++ehrMod9BANrmb654s
VjfxIW16fpoh57Vsi4y5Azuf0uOO+L/rcoXlWd/U6dBSBpGn29vfCNOAndhI25tT
9mGef2xg+AXLqYUSzQrdIIp7a1meI3Vr8swGxYvZO/fZVSt8sI/Ogk6Bg8AVjcjF
uJMDmHjwX25db0nmo7nfzy5yoa7wCpe52hYOq3B89AiSd8a5LFwxMdaX3gPjYGpz
KPETuRz9KsWzQ6FnjsqEWJLgdENJekHLb8giO38Zd3/EY4SI6Y5lJft1xhgirgvc
kindFr1xCQk9YYOYm2s3scX4hFqeDiVfXB5lXJFTtpAqkGwou9jN13Nad0uzx1Eh
r1K5+S/JFhGZaLxZql4thqB2AAPP9feIG1VDmx/KIeM2q9OLYa15SDjJ+ZYJYSLE
bm6HP/WQxuAeR8l5yrYgw/1z+Vk8bUOREqx28N0Za6JoJVDLKxhLsuReyo7s/Wjb
FYTv2vJ2nU+XNFkelg8PXtBkYSDm13Zqf8DnhasyBbyyOFLD23FRyvj/7eSlIr6w
/AL6t0d2qcsOAwMHt9gxB7uvulc/AteTYgDJZ15zfELMbUftv5p7/aBVaA4Rpmb8
RQpt5SqsuFe0t3F4YzTU7uaH6NaAm+E/s49C5fv0ZZ+fuCJa1oDDwcg8UDw9GYNf
1EyebL5DQbfEye4hxMqv0Q/N9aHjJpowiEDlh428SKIOGcuS7wRiwkDOhTr5Ae/V
AjB789jZnN1py8FFVFrxvWO28IbAQDoXESE49JmqyLdd9iGkdWT3mjvA/Gt2kiMG
EealvvGRyCXigzyziRdWyDYR6P5N8x29nEr2i3y0IMe1QsChrp69b7HZmkV/fqiY
mk5zo6skbreC4cDu9jVZZbU9Gtni5OgxT6OWwL8SxpR58bAQomt9B4Cm+0zuFtPm
PjYJCFGWb+HqA/mYrU5rqFsfERa0YbBeMr6ITLdNpcnx3j4nx58nW4pmReXvk2P2
6Ppw8NKDeb4xUb6WZRDEB4++XMqVmMzR5G28NfNN2QwZ6Dtou2uaG0aP5RiXQXrn
Ow68eMDDwqgXIurlJW0j3GqiN2WwVclZzKzdV5EB1y0PmOag561+8VBmgMSlDROb
SHvyiKk5Dob9ok1R/tk06FmG/bR9ckjjXua6yZ/PI23UDRDXbnqyURofXGmUvGaF
BaY8rVcNQ90Lo6Lm9+3TEGoCu0d7uSLtpS2thVdpq4+j+HwyN8iKavdOoYg8gFqx
G8IAwlhE89nMAdPgAfWxAuTowjc4QFlUzNxFyBJjD8jiuOUweKqPSz07Vrrx9ghm
FylSNwextrS5DMdz3fdqSEsIlUmPYbXNGALN2B+cDBBXzryHOMlc3LLZ6g1sI4wq
gFri3h/VNr/YD02q7hJYUv4HZJmkj03AvXWC0nqf7nEKkrG2KRpqc2d78S9Q5BN6
wbhbKiWwpoZ2Zkr9901EICHptlVjCQUFKX9gfPjAtQEkAbcJaNesMB2Isql+h6hp
FeDGeBZp4yd4WE8kzOAz1AAlRV4TJ03CzIZh3lx7fvrYMhoNTy1SoTV/HIJk8A4O
dOQ5nhQBUe91SPqLtz55GUqiqnRORieXXS8WDgHoiOLrPaJn91W1rgFBW2M1D9jC
o6Dg7k1Rakl6o3qHnPT6ILWNWWtrMR8JAR80MVmoiK8u2kUOvLA9KN6je/vb9RJt
Y0G15Uyo8pLVTiYlqkYmzAoLP0w3JUa5q9l2+9182mZqs3JfJJbJkTkA2ZUV2r/j
GbicV0Ekpwg0GMPAfidmDyecDIPFaXJD58MJdDQATm5PwigjUb4vI6+rO6fz27ZO
P9trHVsN+GyfVgtNEvRTR+0PPZJi+F785wJRvZZp+485byVNfNnZqXiVp5GjQ0Jo
9e3PF/PA/4lUVTfoDWP5jQcJgBM7WFmLBsa3Wn5RFhwxYK7cwm+BMZDJY6b+M/ki
iBn9ReM4CNNuNEDhDqMI9RVmrz3auLSMY/ZXXUD8ixWKbEL3oRaO5AAkptOKRcOJ
HIiExgTRAntsjH/GnWbKiQXCmgAD2uLrglSRYabwut2Hy1eAzg+1J7pT/sp2hK8Q
bAyFlDCr865exyKFWw6F8XYyRDIMy1yENiDWc02k4uJT/ULsGDB7eUbKuG+OgeZd
niCG16SjAneIW2fx5vrJUzRRLFuuOSqIcNyIpxsxeTdzbty8tuE9/+netP4HiGXR
/zpgN+WlCOz9D/xjpyBj4LZY2BgCMWh2i18zzcHPd5kMTETGvQ4aFtameEzC4xcZ
j0aqbIYmSKSIQepc88Qeddv1HCODy+cKP625YS+khop4iDk56P08WYIGmOGjn+Hn
SkdtqGFiQJc7+Jm+a6Y89jRsToRwD+jsoh3P8PlFM4MQ37+ZcQzBY0RoDjv2fcv5
z8R/BHLf3F2MKF17jOKCyjxf2UHgUb+Abqje8qXxfvX3kMVnSAC5RAJZy3vt/Ttn
QTSEtEVcEkS9fhSTO7CXZeLQX0vy0oyKG8jkAloA2TH1fwSvKs5axB7z4CpmNLSr
Uct+zxKqQ6bwTuIUia1yiVccL14urqGrEgV2d/pDIFGBomde9cAk7tNhY5tcCjUG
INfpVs30XfCyOGLm/ffWcNxWJJU56ARGZWahrVhA6Eay3F8bN+agEzTDdUTbgUuS
cKolrm0J3jwnIWv43p2Il3jTtevbZTX9/oDyS30fYWx2jsZk3ipkRQ/W9Pkzl6l6
X9bXSvobKgSFs937/046fNBGMMBGiOS+qVkMDZqlYEciR7yUSWil2MCy0rPDs/pc
1KGVZyF0ZIn6K4NNo+LQ4twZRlrBXFl18nMJLhINshWB7Mirk3JqRv4rnb2Zf7V2
tplsZAw+LpFy7Igd0EJFz9CtT+njoK+2Svl+qMM9Hi0Ef9Z4p2KWla7MpwyCdzaN
W3l+tQbNU6M+H+Nu/tua46gfIg1Px3mSAub8bLX8TK49ihuBoXdTYxk3ben2dCXM
MTxSeSrrVxn1d2Iz9zVldu+jPL0E30gqYjjeIdTDjt+HNFTrSXm5mUA5Y19FXvu5
OPmxPI2ScIHMHwP54qNIJ62T9BQlJo4Fg4IlY+OOMHysr8Rd1wrT0caAXCVnqqhy
Mqvx2HUlrjvP4J8k4qpJjBto0N8Cn0xY47WI5R7yUWOYQlVuZ489vYjBQYrQDsXk
8aJDlSqHpBWvE22pgOXjyxrX+GHQiE7n0BDP2QTDGPIHkUgK5IytELm+53Gl1Efu
57LXWR3Bi+zXaV8UywL38F6zFJ6yWbwf7dHZRRHx0zYSUJUzAkmy4FtgDqtDN1jr
aqZIayIWtYMp8fY5TJucsKconIoCYYKxv0l8vOo4Q9nTrUhaVCGYoBF7+7p0GjuM
Gh/Esm9KpLv5ND4sYTLJ5XAs7i12LTKB6Ue+1muwq1kLW5IoYuMFKdE2mGFNssFS
hFFrTjNxgKPdBt1yPzKwAULpa6LV4bE8fBh8KkYu1BpQ35Pf5LQbjPIhFwG4nVAU
DJdgACTpFICzNaIxbSvjyg1ctkaL4uKlvtrXAIzyD8zjgi8LauT5Z60OTD/aJzsH
99AdD0yEuJJjrY+xQgIicx5mmasBFIgGRViD2fsXXv6BAPBvBhN36dR0sNBPeem/
02/F6TPK1xrz392eB1eDZKfOIc1pPt2Wpf6d2e9h7BJcweyBn6MDvRkCZJDP7nSS
4nxNjbfQa57uWiGXdEjz/9CuzvKbZD84j8dpwX7jZMqdmvZzDIrHwkgDFz6S+QM5
YvG+sb3MK2l3/QZug4alpCMVCI11LOo4TDfFokzJtdTNhqRDCkf1rHN1nNc8C3Hg
OXa4maC8jRTBhbSut02Jr/18HDUPFLfL/wyvqa6lq+Lhab7ruKgaaXEfvBk4jWVF
LaArkufGVF6c6214c2fU4gDKbSr5qWgynTTsL0JGb/T6o1dt7FlqX53WCVZyJpJq
AuJgFrxdMpHQsQSvizQZ0mh+zPu6v47354cNjHdDCVSYzCrinO4DM8o4UapwK5S2
GLmnelbM7J+UHof09XQkCvcTdUzteW8OVI33faBgAtj6/8lND6xhImbXAS5t3Dn6
mDWuLGo83nxybcOmsgAXVWBAH0dnqsld3ecOe3iWTjI0B3fCrT9r1smMdQqnZSB3
hDBX8FW5Az1soDiVQlQs+eUKRwtt81I2MBzQ1A2xapXWsC1q5O9J/bzHjkNWnrvw
cHmJaFUpGYPwonThw52nEWCbnZoIQ+VKzysoVmh04PsRoFar/EP+j+ahSzHpRegV
Rg2maP9QnTP1B7sZ3CWIu67eOiLDis3pkCZHvvLQvVXarQrq+OhIAjHguXgSpPMv
XIhEaS1C78qoCVuLa7fpKWC6red7K5KqQZiEgoQn8qypKbvrCefl8Gg/7TtCJo9d
kXMgqeis2LCB6MwIKxIxoIogtLjOWs+dSop6hgqTjwsKTvrISf+uEl80y8HTZeMv
mof0xumyXYOJ4SnV01Fou7Vhn1xZOuVIYIGfGgcRNn8bz7QTZts38VLF6t4P/lP/
1s2D9YsehP9R+F/HDnvF2tdmUOa14lgBwdlSToHmaLbG27CpeaOjM/NzdslSh+Oy
TrXaTnr696jZXFYv7kdOiLOJb9cBwRW1EXvuVbBgn0rRccRayfIQvbecc2Zo5EQM
7Q9NoMylxSPLXApZ0GtJTS3AzgLvoLtzbJM5fQ+MfJtRRf9csnViEeMOABS5Kthw
vcm30dhARwqPtsiEXfeT96P76B1XDyfAsoj3jz6BgzI1bIZbpr1AUOb8gvILZRdg
DmoK3kuXlbcJ6EWs4eVeiiXNuNWIYc00CIHRDjeVqA7K++N/ZCG3YwjXCkgvnPV2
uDusr+FHbFqyUNp4CdjAeFfPw9aTLWs5UdoAX+lpyhYDSDtu4ZOHUg7zKT0yGAjh
AXlu9dAYF4ucNgZmoaPqmhGyawMmc9RrLfcuC+rRWak1aaN5nU/ZZb4a8r7bFZTS
FRVVLdiRdculm+kx53dn/f+UReUgP6NfHOp1CyL2WBrcHTDQyKEMaKHUiI58IEOE
KH8XFKEbBIOdquQab2xFmcLihJO7k3LxZkSY1ewCvFOBRBqeNTwTbeMXZ1orBPi2
likh1/0VSwJVxlxJQOqumIEkKGoTC5SCLoD951FwxPhs/2kr4PhBGJHLOY5TdPAa
11Kdsw6sqCe5gMDfhsYf6ljeenTNnGMl+pwGKYrqIYLQnm7tAw4HiQGxy5X5jglB
fLcfc0n9m1XeB5VTBHhZh0m+X6izkro4+HUi6zDFkxAK16Msz10Dr1RWF78AEYjX
ZISndcIkJMeZQ/bbJeHb/r3ZQ8xH+rt0ltEg0vu/l3n6EayByz/hYZbOzA4vYIQ5
xBiAZZW+PCJWv/0+tM8fxy0RD9Xu2ajBoMeyd+CRItJC0W/NUAGkOjskOnDVzSpp
MJBK+Lvov8vydiB3fIOr0QoZuu33gxrkDmyMRUucmK7abcvwDWGv9zUZGLsbxZZG
C5BcCe1qdPzx+4rpkVPh35508u1x+b9tnIRZjdXZApIpKCm7q95nEa904hBVCA0w
heiOFshPOHzaLAN3UIPqOGoZFXVOZLmsjRddSgzmIcnZb02g+ijY5Xohw//arxni
Zi1tzKRdoXlnATHQASbmOKaWe0YWnlqcHhXHh01pouq3RVZY8E1o8KNVqH5dfG2c
LRkAeQuucySNEZ84W1SKr7rX5oj+fvlA2Plv4cRkBwLmlaWIW1orsIpEsQbI0QlG
h/drSD1D/XWWfZny9qE1kpqGjSi+myMWK0ZUCoztZ8te2DmqEMNyTegsHKkuhNHm
ekHcDnMFztn6aaAm81P1d4iilGVoMarfc0VdfxkErhh7cey5ELWrqFyz0/Tjzpn+
uaEbKKmlduYUd2SKyfFFdW4UsB7JbiaUABFotD39DGpM2tZYtX2cSemCT7jdrCuk
P0VHyfd7txEmFxb6Czbo1z3KjFdhC/40N6HtIpaRH9Fhq4UBDPztQIv6ab3GW4K/
nlUx3oXh3m6asrWxSTbg1cKVXfXmTtwsOsqNsEsir90s+qhabq7YyyhrXxp26N+J
4NSftk4GbCkA/AH5mWXhR99d8Ag3cxwZTAxdd2l5MxSOqUKKk6K/LUg/VSPxbn+E
m/zfu1Cp3j0LwMDBz8y10bReNUy+fdbjaCOiXijelxZOIuYzf9GyY/BmQi2qMX7V
Opornf9pUlFFt0U7GwOlsCAXR+FOYXYY3pJb/KZj1pkxu72Wy0OHR+xb6LjxzkF5
tZfzFph4oCneBr6usTLeYQmuq0euUtN7I1GWXZqq29+HLbKRYz7mWa9p7cWGgXt2
UHkd+7ulKYlEE+Bp5KmirsNb53uPxXXPC2rbBMTK1YvuWxndPRKz/IXKnLL9xIH5
IV/0IsBsQtxFd95qZM7UDFJevH7iiGCCaW2SMoHArYNrgcQXp6wnakOf/U3bl29b
Tk9UphXJ0Xub+7FzkVpxkd4h0cCCjNW8GQ3CtYjDJzYVNS3YLhx2fTowpvqurme4
l0Mhp5qG97EazH/Sy4Y5xSTkrAuBO6n92fPPPjTyAFNxmOKzFIkhtBuhziI27pZV
9mc7t114OWL2p0UM1g4Nfalk7meKko9uyQ6p4vxs9uUGjsCaxuJXDiARHvX5zmjA
xsbTt+jhQcoMOCQFFJoFrFGPmG9r4uvNOo95CnWyGKbTpRULrmLDfHM8nYeFNrh8
qxxNGJm1mfe6Za0C7BiKy+IdlnsMTpUpigzAYonKlv03jd4MwbYZuJP5m2pQSv7I
JAhxpszHqr1qBDFqZG5tZTH0JfWfBPQyEgiYFor/SRxLGS4+veIwIB5jXc6UK+dO
oNuIiRyh7IhW2Zu+bnXCSp2eDM3gTSgQfUCJnGSS7x5Vzh44HtNqNwOoTkQTWJ+N
EijPPcKmsOJTyt60M9FYHmjQrRuklKCTw7RzD1rM8VRYC3nHYR1TwmbHbfHMeWgp
KXa57XV4d1eowFe64iJ8vGQxNZNlDzM2LfNeGzmvz+nbJxvdIhhYDnFVhJZNoprM
r148O9Mfw6IFbwkl+ndESPjOezQZaZGZcOBhBITU2bjdrPUpDuRpUbFkQ6o6DJ+Y
FvfF7n4UndE7UvqP6VA+bwjMy697r1pkHBca1TU9AaWSsWqcp1eUAclWgU0mCrT5
CvRHLv9h9mBOT8O+y9g6JygcjagAzGkyoO6jc2PrOP1UW7WhMhT1G7aUW6IMenW6
tMCqTy6FgH2xGnf9C+SPMEcrCSMo2fhaE9jluhyfdAVho9n5t7LoGGVoT+LROxJk
rPjxIGmm2+iVS2dbNMewm3TvDYm1IrwdIsr5hqqZH86GZtwCWQdxIxX1UHLzZfy3
Gp9ESxyiNWODYUs/8KMIanOOW4VgZYDz6/fbEj1ZaaObh+q31PNRE3ZHJVhvfiD3
NISCAhSPAei+PrFu3vyBLvVv+TaPD9pnEg3Fegnh4xxlY+7fYEoijvvY53VMPVrS
waLKHM9ojC8h+BOTLxfwCYoxotxJJdNKWURYIvzWwVUezqyaAcnCJDlJYOB51S4o
VdQnV/kos9LR6rbo1qQZUvlVaI+/sEvze8uXWikD1ae0WHbQ6wCrSrMH2xb0RuWW
gjb/F0unWzD1eSVpfF90tSUllzfPb93G2cAUQDWrNipyqrW/dXZEj2cwQ7U8HBQQ
r7ESDix3suuqxoHoiwcoHKqBsyK3HXK434pS+XaAJSr7Bx2YnTL4Z2Oq4DU0Lx4q
ScVPRjAv1mzLsbO/fzTO6uRRZHA1fKvaW3Z9pUdS6H2i0NgNwe0Zhsaqahrmwoci
ry7xx79SwXXDqdhtjiBJkDsvmt4pEjUN/VKA62lHNssH3UE57P1Ptay7aMg0RhqK
aFDsLyYpYDYE+zRrUDnaNoDLmIMs7V/Zyb7ubd28IzVTFiR8rWqDYxLMhI+6uIw6
/EZ+Xv2Psg9Ne6SKr4jI2D1MENNV2t0gyiZAxxCATAb3ma9MCrLzS0v8VW0BFlnU
Zs+f8FDX5cIvw1u5uKuDm3D9JTpW2s+ZTGPAeejUTomDFdCSzqeIWZEuzA+kDIbq
pgKxXY8tkJtqWrTjNUiZwavGwyLMTFWi81en0HRTurQo6U3UAJBBXSCxXV168aAj
tagvS+wgpKi6gAgrSmNXA26Cr46bg2/jh66wUYdGNvI5pl4JW73l/0bF5+riCQO6
E9LYEoGJzEYcfq76iFmXzNl+sCJpc85DVvWFP7McTxm2hF92sMWaFSGvQATzv6w2
7Uo2XXAAKgCcJcy0lN2JDCcp37zfB6L2DO32m2CkhTjnWgExHonMFBagdV8oN0y7
WzD/BZ6CTfSC8eg8qdgdyy5VQProajzXrbWP7WwFLw1c1yFpA4VDfwwZ70FGmct8
VYbw+BSIZcOKZ/NAUC5UOjVpCk+vG+s9OZx6frmd+dU+jOz/OXZiQSNSixKuWL98
k2vgtcFogU7mPh/48GdYDqfhjeRpWq241dqKBhiACSeAdLnAVMnO+EoOqVV/0LjO
ZZVDGTUUl23Vmc/FtJFEw6cKHziW0xAUuQE0DeRm13dMyVQw5dD25Pb4igrGvBn+
GP2MHZwjJeIS0UpKmQg8jDRUqiUY5BOwDLaHZH4Y5zakLU7BnCcy2JvaknBd0Y+g
J3vUJlW9/OW47My+fBt39rtzKylswNnqCF7Y0ArFXGVXYUHmcyhf7pEy3cg8Jegl
bL6Rzftwq6k/x+Xb9dJ66USgy8ZaBlV3wG3dhB+rYwag7R8r0cPpZxuGEOi+JT4w
IKt/D4fmOqjite81sX05NGyAer15q0FazoEAEDsJnlSVctwW2Raa/CQ93iGoYXF6
aPI15lfTkvRM3i39k9BiLUTyX4dmplCybuwjRnPBYFWpPnjgSEfBwoelqhZrreVk
3onmKpMgDdJMeuc8rkpqADSyNMBaVtvxDH0F1dLJTkuYrOkkV1kYcYCF3xbOFUTm
XLFsn7nBPH38mI/knbSKBE9kwG+lYPlDzVKAmlBUFKD5kCvyI/WB4ipAJ2kn3v9Q
0sAtLlud8/meLPMIid2RNex/FNXYA54pIJjkSMSu+kRS1TcpP7kPoowJDkS4i8IE
8HCJYawI86+YZSZCVSW2QNuwBogXiHeZCMLCCJl/iGdEKJi6U6LoC78aTVbb1/On
ulNSDiVo4FWGLy8N+U9aX9eWyKgQtU5wCQL3lwId9U9lGEvl+lPQcRW8rBuzeK11
A32dmeOxujALrdU6L2rHc5sl/xarrB4xy4uzpgIr/y/vtXZi113DZHvetP77aNIz
cc4I8AgemoUM6XMR34jaCgwVmmbewmfspQfFd6yyLXfg3qsCXLd3ifjTAm7aVuM2
bcuXc6ECnQBIPP0BsPOJGjUasl1VW21WFQddffdTKsUmV7qMPDiv+ncUy8tndyUP
J1EJatyNrsEpOVMauDSkAPLBHyKLXlN8b6tC8ePktDpb8wIxdYOSNXZDGxEI7E4q
cHGQZ/pItucxbR5CmQJAe12bGOKMERN9G/XWqC15bnQobj8i/lfjCfa96E+qxX7f
zFfZoz253aNRRE5kNseBCXF3M96AuZfrthy3/cl8NCn6Jem5pXyEb2x1x5yDW++4
4u0C07rWXNbtaWXVQzEbTMdiQc6wFCpSIL4aGZOsB66CDjUnZQsqhkdHUxJ+rqpN
cg2/lrX/WCUMWwrnBf89Igj1GI6nf/YoYLdPh9bqX2iLBRowX5+CfYS2hIziB4YC
hbYNP1TbGM3/LdYRGSlTcqpMC63TCPSmsb40U1Dd37SEd1f0ffFf55UFm2BdHjry
cfaeCZJ20XdD35UFSxDZeTchtP5UwlvV1OzR7YNJs6zsRujFKPkq5zMZxHV+Va3j
NVnX6JSs9g5zSRxBB1F3z4slrJ2+SvpAQQvkMsFIf5t8MzRnoC1gO3qaHmOg3h8k
Fdw0ILyEd3iRZTZynafIXlmAWj65LJYiBaSm3qEN4zh4iVeBZt19TavKxrXhjdCo
9fHotMhuaLOpxoPgmgvCvfdY7Gu2q7nnSNGZNCTrdsrVXl0zwU6mHDe+Qyk35cfH
8TRkFk4y7ojSExx8+IAIDJdqUihouuvhOBCUj0yxqMI7lML6BXHWXrUN9YxfvvWS
FRsWhbrii9MGbiD2HAXMIfteOdfPo9EnixTLuSRk3RiBxBKah8evzd8uLQ+Liq4Y
bdJxLpmJ9HbIEzGi3dVwKJ+HDCi6NHyIyYsKZ4l6ckHQu9tr5cc4z7tQOn/BSTgQ
hohVmlY2njR4m0cblNSG84OQlj71Svy8LB6/eDVUOn/WY+zBl94OMKxG68fmlrsm
sCElDGR9vAeDrilwubKM1Z7qB6rnm5BCARnatyGw1tMCpaOITAvbZkUtxTkahqt9
xYirbkNeA26JUj8Z9mWcPaO1b5YFm4+Fy4ERie6c9em1pXW3RQZBlJfrNZJTGni6
c0i8n4lShQH6ZDbCxXa/Gu8QGC53ZeWJnVCSBmk3PGBOmXnF3Xd0O0QyhR6IqGnh
koPraPa2pKGmyyo8Z6X6OSIR6BRz7JOwhW+UcPsZ5lvRjjaUyZoDtk7C3PvyglpY
Ies77YoYkvfKhOhOr1rJtgLmGPbVqfa+G6ljebEYvvmQjVaOoXRiItw6HAM1qj28
ZULt1HUW0o+t4mc+a6u5nQTV/iUJBKaxVfx9RxKTcaUf+c+nwx2/ezHAaN25wBoG
czKiqEkDJWV2bPJYYbFBbYPWbRKrVme17TRfaLzpAV9VjZm6QW3vffCx2EXpT3O1
XLV5QWYyczeNm7/G/GSd8tktBTh//v8p6rsjV1jtJJMa3cG4E+SxJFwrz7sZo/Pj
UPGyYlmyRpl6Hf1Q6HgfqjAWkxCLMYVe2LWM+G4a4xSZKYekazUhkWBDBNzIMaCC
UWdKg5tBPiIid8lD+SlhwcBxCea/hpt1ZL3LN2/KxnIlgjBQfjMybOQRJw1YfD1h
SGfQfXkQEM08/qjI0h/MNCkG5M3Z7KVPQV7httPZ5CE/Wm6+iee7PtiHeWVqpV5s
/HoCgXD+KqgEhDftaDY2ftA4JpjhPyc3vHSH9J288BrZYWeXlEOE+UXj3m8ydPmu
H/b5A+HEf2z5c4gSx31Ypir1kolfIriXXJ4Iaw5GLWv7IR4Kyp6HaKC1ZM08Hl6j
6ncPU236H1xVbYRMLU+OBv3Yz4Ws54Mo1ECwXoJ/uXqbBEu6RtXZKiA2PbBX3HXO
CAX4RBm1ZsOjkiAzIn+3zcXUCX+6bcGdnDdUm+QaM4ejtZy+738HE1+xdIDbH+uc
IzM2O3eJg3Pxdp/lspGVhFtxM4HZV2CoTNzSLnNxCFypq97GOWxm8gQ9EE9lUJq5
yuPm66/f4+dSeg4MPIbT1g2rE+cpG0BXhKpUd3hg58Deo6ePHU1SBo8S1H/S5SO+
1KpH3u4bAznnO5zZUS19nnQHKKWJWyqlm3IAABSuCnOXs0pxD8iU8vrOMb4BHMSM
4hG7+glaBE74eR+YPTMn4AnyAKYnAzIBFIoVelLjACqHUDxrleLg8Vbx0f+gffpU
om4zXKZtVmBJXh66Cwmu4+TmovJr3tKmdQFViOqS0xvbts+H0cWGi8CKG8SWf4rV
UI5WGk71W1agUU+DOjbWIrOCRbWeOXxLRktD9uz/zEv39s8PNohKXt1Pktyl0OE7
TWgp+tz0PLZ7uteZ+7I5zcBFb4f7/bFIo9uEqTUUdd5tU5y0ndkc4IPscg9c5cIE
jWiZX0YcHfJuHPdip1VUinBq9AAqJAS1me/5Yl+yIvMkVgsZQhD/PCBf8zoP9TD2
Xm/aVExtBt+OWN+/ZqG8V24UrFzXYVGKH/JOIy+4uc2qnAkm2Xq4yVIXG8jaa6rY
EqEBXd5+kuwYNEd51+xGjhfvQYznSwDVf/wwlxD5wt8aNWKPCV99GtIp0sO/Wj7W
6yN7ptdIpxF0CojT6dfmNyvhK1b/Ccwy4nmtXBIJ4O6cOQjYerg3hntQlyOfVnZa
lZ9G/NYw4g8HOY+/Y3eHp3aPjzbGCmnJj1pnXrJukNWKZi5HB9q8soZID4dYsMX4
dgZWV48gwJM0ku4UIzg55UrNEA7Yz+Y9j/JaSow6zAl3D5S+cEO9luVEqXfK+j9D
NedVszyOC/Mlcw8hR/zwb7n3BzIJfVwmYWbCOJhMtvKLUCUgHNrxvRKcwQZr6xwX
qzYBsA7o/7eYpoDTvFqzpRx3E8LkyKCTN9timPwhjZGhp5jU1YDbIhKI6uuvj4n2
HMX45aY6kX1S2THUIf5jncXSsLgP/DWUta8RbyncrWrgGIbzzGuZ8xfaAvXEL8g4
CLLsJupd6cCTwNiLtpX4p8LTchmtsSXJeaiEik6eVtEUKoJZWwuU8goGaNWw/fER
x27cS+Tv+tGbLZp3nBtuzAmemVp6BqCj+G+cwnYrtx9xQ7JXcbN0w4mCH+07JJnq
JbVEMob2ncZaT1PBcNhO96O5UHbjTjH08FmZhLspTJsm8GXus4/LAJzX0As2ZA7V
mEB6WsSpTyYI6hyB2kmaHLjgP7n28CNJe4TWbmhe3PCvQyKaOeC8nIPi2Rg3jsvO
0asEQHhZVOrqHh83+u6b+lL7DdOsyEzs0c9j03elY7mBi8KGoG2yhgBQY4ISJp3C
+3Dj6/d9G3xF262bvhKEF/4H1st4W5OBGWpWrbQQOPJXmXwENl5srfIKsRqipc1t
PPZJEDfJA/lDdupW+Ax6hl+Os0oQC3kVwYGpmh20bSk/sOm96MAUQIPGi4VF9xmT
jbx2dbSxF7OUvRa/W0hAzgsOXD6VLX0k5P4xHDt0qyiavssQLOoC5+vGroBBChBu
2myheZ2x8OPuK2U55VggR1s/fadccOf2a0j1ImPyYlTAJgtUlCQXp1zpsjKCS+MH
4fnpFFW3fnr0zeMDNc24mKevLXQQlcSGWva5NSW4WAkoq2owIpUqdys2TvCmjJ1F
ukrN4bFYLlRrU851IG7U0+1aDj/vxs9V9F1nyvFxQi3Cov5ibAnlgJ+fmnk62Rb4
co0LVdTVJnjeZIVRMTmqUewKnq3B9VN2rEcG1H6vKXkhjrqmE4cTVDLdLeMpFrTR
Klg/Ml2vacMu30v5hxd0U240q5ptEf+MAkYNWSevraJb9GKXD4jnWv6Mfqf4jB4a
Znc5BEmmAPymzN+T0/iVsAIzeDcxuhRmdwztdvIHfV8XqAfNEa/drVKKDBto3aKA
BHn5FKlfp1SFREI2JOkxI+J682jdgXrOX8HCyhs6Fa0rXXIY70bIZph9PQPgG4rP
ARvDAVd43eYwe1Zff1OV0+dz7V79t9BUv3hnGh4/w/z2Mrb8UlJcvlqv4J0+Aonj
lgACeXQbktf7hzJ5B2x4GXC15qJX2MDKoFJYpa9ko07PDoTvQ6fqs/CxQEVJ5tVq
KlmPWKhIfNTaJmOfFgoTp7/6GGbLAQA+qLMIfAv9yPqLGAbpJ/spALoS4xQgGeRR
EkfHcutGh7bRYgbA8vTTeBXjDuuU2tyneaMgMjFspFRwOOnjwnFxyzWl0pWBYSJg
bqlw7L7/to3+QpCF27WEZ8moWB7i6NEHLXX/cOQGXvg35RThzelHmWSDeD3MFGou
9VOdpe3SfL9JnL2WK2dyiCtuL1b+Aqc6K1iuxB4H25sC9d2FJZMf1XhLxzyJFJFu
G14hNnluUh6GChpEdnMDmYww/M9FC6vpRs1hFzVeTV3+AKt7v4twoF14CChzGRxq
jlET6FkgMkCSHJC0lV5LGnJ4DxCt0fwHGNtvYS4A2avyJ/9DAF/QGX2YGSQLhu/9
fy6bgP0EWJ/spkR7NTxyeipKr3ETcgzXCoMGrK/3jLLrPRTR62G940NuwKoJ7n5p
cvh3CWwafGlr3t/32NgoQ51+4HkU+cGcX9ywPWohWPweC1VyzMz4SwpaKszmFsmx
aTrv6EAjp0tm/70lWoF6HSi/oDUrsE82oqhM21J7oFcuhxEFu3Xp4J/y2yHecoO7
kQJqR06fwO84VZlu4ZrA4+EuGLhJwPlCspbRKQRCYUr6cIIRNTankBrqWyHus7al
0sokqE6iojvtKQ/5MfD/wUKxS9qqXkCTqfvODideBfjRMY/PZ0lAl7QlNNUuVgRG
mXwxKT7N9/VcO1u86bsfWVIwgGA6aYipihiTjRNmGWEtmRSD1xKIJB3QAgHR/dYV
mcd9OWXAtFuJhLdcINTt3AFAaPzyHERmE7OVnyH+/Q4ZuEMn6VjYcT/kd4u1ZmBN
J3OT9rui0h4GkRwQUpDjfnPbEJLa7PP+nIpNvZlewS3eLub2HSYscZhl1KxmgNnn
Jp1R9tiuu6yq8fzVzOc7mxBSx/32VM2qxpWR5lVZkUjQxDQAEtKDxRa2kq6v1f23
kZOf+5KIE6BJaqVc/YYlcWynfAPbjTnvhCYUkHw3Az5DVxtx6tBEAUQ8KOakagKb
CDUQcbj0IUz+BE37jlEQczySqd8KAUxPftS2S0b9f5csoKc1qiRK5EL8NTkcUgC5
AX9vdp+cJDhzD44F+c3l7iYPFeUlW4rXBdSnkbGIDaGCXJy8Obg0bXY/C5DY2/ah
LgrfzU9M4Y8EgLoMofjRdVQnPUTl1n41irUfvFpownGrbfwAkC+Ms5t5z7Ww/8oV
hxzArXNJ/0gbxowS3igtewrUCuuCuCFww1jvXXidGcLekAMnTkG+oC7P3oEZqbtW
iYcUrZHV3HKUNcGhJsFrZOekmdvIR1sm21vC3U03CaWgjV03C3ZOMQNw/N/61APK
OfmjTfn2gXseneOzSXzLGDkh+d+zj9cft8wDD8TAEezaA4W5zSZrLxXZnJCqiiRz
VVthQnqUywCSNoKYe8rg0yEHcyquNUhcnKaC6yUHqn9Ud8rBwX2cL/dKg1Z4BN2A
EX2ticQgLwGahZvtrcZ/5i9wt+A7gUtGB28URZi7hNTs0Z8DngXICrjsznBPpr6z
RIjPagwgkoP/Qvc4QrxX5N1eHymoHXswVp+M0DS4Y/5h4Bj1gMLQkgIXI/Y3HxMa
EbL1Li/UTjtyTdsNxWUyhEsgIbeupjLVMtsJmY5XXV/ZXigSwxndYLWn2bF2Fkdd
dzKStflTK1q2l23jSdSyYP4se1FYybRPTqXlQzGcV3HTvsN+5wvtBFXdfJatTXQG
s3n4bLynmWmQACsldRYRJo/xc5pZjyo2Gn2FPRjRY7HkbhoG14bFshVJpYAj59S4
3O9iJ4GIAU/YlobsIoUJFdh5vC/W0O8hreDEreh98X91OnLBnNSNBs6ugAmB615o
to6VwJ/W3rNozKt9GPI9wpIt/XCH5P9e8vilX0LzZpU1wEhP0AQGKAyDkn7dkH32
eMPRsE9I9JHrKBeYLOnb5HOGcZxJ0ZRHvoRq5aPvhWXt5bz70LVBEIivNlWmboPD
JT0Rrf0fRQpxbgZXBfDy7wHY5sqN3r/1grH7wfK+7xQWuyJ8yMz+tHL6r3vo3ffs
DP3trM7fcIzmbUNgYTvycIQ8YCU6nnuO/jtbQhf/aDJPc/mPhGj8KhyLimVSGd4t
+FXfVOKA+jayBPgd9QsIMwdZA+XiIB7XNaF730wBlyc/QeA/V4lBYC6WQ2XbRwCD
G6UrQjpz8RgRmErPZgZ6wV6DS+hvjUV37usKSD1Mvogug8i06x5ALOWd0BhHBPOr
T2aESENZ70wVMTcsp9I/4jpfoQ7itzj62LSYuM8mqpQCkB41eECY3LOmxItVWvkN
IjGYR8NJORWvnOOtu0lsqYjjIveIoWIaYaDdWTw8twYMH0J1KspfujGwrukb4Zdv
vkIVsLpRZCKDMApSXHhLofzruL9lJle/vHpQBWdwR28EnnjRW9XNubtlybOdYsrJ
QplKrGmAxraLcXtEpG/MKB9l0SxbDLP3y2oAGQn3pADMvu3+pMzmoTqF+HKe7wvK
Rc//qXcjKdtO5LkciApFsohB8JHZBbTi69j+dWEC8z86C/MkHQs9QrQcmandQZuu
Q+VjJauyXb5IOrcqFuo4F7OgY/wZrLoU9e9F531m/T9f4noZEvbN8x6kKviFZkyR
ChKTyZAoVElHJfZ6gtmd75wBhNfBXsIHxgoj1H4540ISamp9TEaITgdLNs69c9w7
7cQslvF0Ph3GdY+h0Onc2l78F+GV3Q9Mv/H6ijDYhwi8O0g0qdhKSdDPVBPsemTQ
HqXBzsg4yApnJgFa1qyOzdYe5hUv+ylcALdH3ZYh7eK59vmozxmuGJa3iwKTSq/z
6zPe5R/iSF+dgiIJItlw7OoamQhaB/lhLccobhY+R2FUO/YiKAUraYOTzntgUUnr
26CXqRCKMNiQ6ZJ90psFR/6jgr39LGrXNyb6CS99Zp0mVo5sginvv9y/5neb5gTp
T/63isyDRjDcP0tw1MDFn5tecZzeFIxTcRVNRl6//Xp+oSmZMm5s7Byvj/3a2HOr
/lundyqEQ5f2pSp30noiZ7z2+9NDoHtmARntFjnd1ttzTphUUL1Xhbjv+lCIpRfC
bDlLXndXar0tz4jd++EQlp3n1Nwuv+0kbtrjPPnokegsczYOrpd91N49CP6ZrOKw
XYQ8mq1YExXVpXLBYWVKJhVZs64a4hXas+DshGKdWqaK+N05XVugcj36RrfrohTA
ThSQZ9EpsBzBrHgB7ApKXua+QmQfMBRvF6mb3KJXoMHmaJ4E3irrHFI5fhhdt1Wi
DpbGH/r1Am/Ka7hz/UQaQ1RG+KNwIJUDuSfBSNj+mwO8Kxep6F52ff4td9RwmLh1
J0z0OT/fQQZU24IaAk70S6vNzr41bBb8NWHwQHeNR3tlDxkz39AaaubLBJc64+Vc
XFQ5kh9pRehNCufsPmm5oiIy45zljSL2JtGg1psUhAyfkRXZrCFCtWLlU3aaau6O
8BLwLmprA58kawinwxoLh6binowKq104nHCOvu2Aup3vWypRKISAlovC/JzY8a+g
N9C2rc8GXVfEAhONYHUB4r7Q8qSAil+Vhzy2BmSgwNhTRe9yEOVeNAwU6EO5zDky
AImUqA9vVElmAOiEGfw9SWWuKzphsNgM6Kl6Cv+QtbF0SH06UYYKvZrPbzQMWyzK
ilwHzFmleJOCQUkS8AAzobmiGbiCrr9pOwY0QvDkGxPUUoN63BZ0V532bLmqBTIO
ZQodwAhsH0tGNcPAriqAs6lTPDXuiaVLkB2c4yBCeFDx8aQpMRniX4c1LEZQduwI
K0UW9YGUD4B21AOyNPqhIKcgXo3Ty9R8ZPG9WQWBZ9b8bGcFNEDM7Tv9fFuNDjZY
bt7mqX8L/UiaaLCcm8yuT0lMkFjtkNCvCsjyvlzZ4LsD7gqhaDidNiMYokNj4DG3
6G+hbCCH21BoE/wicolSAa6agEaoZ6z0x+m0MJdxHaLbIOV3suBSi8pch3PC0+Pm
n8DmLn9kJNdW7FN3X+YNeIFH/t8gnj5N1F/snsc1VX4H11cAZbrpB5Zxr2Dhg9v3
TV5LIB3DTpB3mreZC+jf0oPMsyB36ASNWaFj9SVqNPDVJSb6pEfuG48tRKqUy/05
AEEzN34WvuEPknRGaVcqVZFzAothSHrg3mo4i0zuv0eJVj/HIza04CLF4+NFYHlj
SFdk8fCDsqXcRWVgsOfl1JqPs5ZqOo5Nd+Rg3a103h0H4oYRMau/QotGN/5S/Wxf
Iy4MzgDyA48dXOEnQup2WzynqANimEeout1QHVZZSfXXtm0GV2FGRZj54L9Va1dw
lUGlsrO134T4BluWvI6dF7MXN3bBYe6kbIOnBEYIO+KiBBjRtmxtAHbdYdIHZOJ9
sN2yIuKMy4BJZUaO44b8g1iJh2KEuG/ylE3s8d7zZu5dV1rr4G/gHM/LrZVQq7h6
XzCxLSOZNHweR0TpT8GWlzDpvs0uIlhDfyZ8CAv7mxJuJyyqmECQdSZC9TJd5wFy
DMhvBYJKyqFn0Ylnji87QvyJYQvIeCyxPxQOKQqEaUH048e0qt5nmqztf9U36zdR
DB8YSlurMFFOOQAbfC44YuYr4u94wOiEGYizSVmMsZka6DAOsPcvrlFMMm2rzPz5
JZi6ntjupjsZ1csgcaS3Kw0Ovws5/i3J/NCRELCw5Ig22jI3kRGJ6stRAA9tF749
htJber8TCXEOIFhF0OtcJ1ZbwvH5zU6rj60cfndds7CZNWg7pM2Ub4ajfK3Jdq4c
1Fhl9BVm/6XwwawhZU7uatQxAywHTbaP+gmiv2el0MV8oGyqtM20v64bqCoIMLEJ
qe06uwVtNdTmiBmlV3BMuq2Ri3cIEWPIrM4eIZcxNlO5PANN1oQzZM0l+77vhRrm
5cdNoPIrVvBYOey9a53v2t0oON2GOjAqP1twpiqkqK8CrxIq0+lN2mI7lzmZ53Mi
NR4NJFfjwHTqnoSEu1t1ocN5A3cIzhjrIIONnFafV70AuaEOTqxfIo43SNChY4Xn
3K8VcebYXhO/1DGuiiLmwBFNfeuvVhcQyHKj63K1w61lnbUo40nRJiUGcvjxzfIe
q1f8lHyqnOeJ+S+R+jnMg16RzVPFvYGElwDMYDx/IIg3mTfgf+m3NeS+Ya7oFZ8C
gZGgaefoLAK8+Kk+1h4KXQhLXmqwinFjaXbJhRxh9fOWf7pJDSZ+oChkoaYIRayS
2+oy1yDo26FzQY1+hcHFB5pN3qlDwP1cp7f1GR0mrYeeIIGdH/woML6jnRglqdEz
2/NLv1TRqa79fu6FGKfqeCYVUQ7AfZVGmxpG4SOpVYLYBluXsaiGWltwtx4GJnbe
FQnnEYvDoGp8b7AzPoJpeyPsaWdWT7pjtoAK1bEJF549q2fn4jcPcAbU67WY9BGP
wcvoHhF4/pvsZylc4Y0loptrziYFc6EpRiY0M8pdHqCtBjsySGpEFrMIZJ8Fhntx
q/PExHNzXgL0srIFROPPXHiSJRhHnigoF4O2OmrjMsDrTM8drxMUumgLR+APotNE
B6zGCTsxeOQEe8vonzi4L+A/py/3XPl5BkZb0FyJpYB3NeDedeoiApAptOEuADxj
7T6xuMMGqWSbBxFfEQ5koGukHgwebzevdDpb9L9mJiviF3KPNJtIqgSFTwNs8LdJ
382eD1Lydxt8IUxNlc4AjtDc/xLrLcLnCQlQc3ojnthoW5DgwFa1cxdNe+jU8xY6
nh/QsvEgMkunUp8wA7Lep2GApIeiA/re5dO5rd8PLxb9W/pCa5viOXb6TosoT1Jt
JFh7u1IHFbhfQznrliIRdq9XLKpATxMjT7mibc4whOfDV90iNi5XOMiruPI5nYlF
WDaVmtU1yEbhIqJGnG/hIJrh9g/mf94zjTEyFr44VNTu+ABVrYRXWv8Su3l3TUHn
DGxgifE7q8ar1krZFUzCgb2yIds0mlxdz5MDY/ccA2RGjAp3ueECW+WAIXJ+882Z
7QMaZHrcwfyglX+f3GvZd5mkU61RK8zM9bLK4g1JeKxVQqdKk6QwjILyUzk4IhCz
ZRyBUWSyO3tky1j4kakehpTirRWrHZKwP20qyvIFJD6/TaGsOOdgtMPV+n9BQRwW
sBTq/PX4Uvwcfz8V7X8EziKXS/6dQjcN9EZceJ+o7x96asjGYlPjxzHparOegUF2
qEA9wVRoqSO+gJ/9x7MoxsunGPvXiN4ANP3VrGTnz2MLHhrTGQXuRMeGQH29OFgm
pLEXj1xw9lq6BCPaqodOoL1/Fy8oQ64C4X3XCopQDel0nMOFPjJF5czeiBLinVHv
xjFpiE5OPc5l3IJ6yb9hw/fadz/3Izt5sggNMOCyZcMS2zLYN7etaHzH6xdHKzF9
p+Ol7a123J/2tm9kySGpZL/0j6YrWV5UXyGgFZcBc6OE7qdtbGAItImwIR1XxsLw
QmYIzVefWGNYQOiyIk0arRZiULU7aCsb6nvHxirvU2nx+b2GIkGVcxdBlaGYDhjA
f4vJF51DZD+LrqP9n4G19lpOJIwNKo234fSxHxlU5ULqN1Oz1VIv6IdH4TsjCmzd
lvjkoSh1Y8j+ucY8V96GPQlBIZW5QG/PBuTvjUjP0WE8LIPCYwX5kd6g8+NbqaOX
ojsEt69UH5S5HnuMLMt9DxXW5OpLEa8FQ5QKvZEvSqjxF4aXB6B952Nts6RSpExc
lsDZgEOt/rsgsZ0lPcJC2ccnyl7L4gDeV2wHhbkX+SHBPwHvBw/aDwt6AodEMZZ3
weD+AuVVkozkBqC3loiUR7ZsgHiQL3iFvfWBFI3xYTL33a8jY7ky5RBsMHFUuOOG
MXqQKfALVwKoDka3rENJyVLWiWsolbgel2MOLHxAkpG7nEF2tBtfS5cEewLmQShk
IvKNPvnyGc0pm63+EOxtxlaQuB4q73MMZSXDwN47tAYH1pEfLGOOyqwt8TxNSjSV
X/p3eyV+JDHov/H81OMvAua5Oxm9PHnbGNjle/vr192Zrx4fFHKdNM0vt5JVJw10
bpNnqQP3m9x3HSNa4rTtaanwfKhS+hA/aEKu1ZZiGojoklLy1hU2207sIVpI52PY
aaW0+Yu2601lQkIlfvv0EG649YCM5P3qYxESXYnVTrNuz9bmeWR7QnQ9lwZXBr0x
qyti/e7myNDcvrVJwlnP1g0ovRhmjgx9UZbdGIQucMGq/0pCu3Hp5mky7gvi8Y5D
4IHFKW1hOxVskRCxnOmS/WTf/qFSO9b2PjA1sJkS9hE3IaoExR638uyABQZrXYiv
vq1JzXNdgxv+U1ZdcKE4aRgEK8n1/MhIGJcdFwJPllbUfwdSmXFG991mMyqvQFB0
XLAfSdjnTLNUkshE5ffaxTpM3/crrvmwyIqrlHbBKNMw05yb7jYNYYWT7YJyZynY
+BJL4prQFFGb2Pr5a7bTK6bTcbxvIu9hdjYA15RDBayS8HMSC6Wxk2v1CFbw2Mx5
RE91m/Kcz63GOG/KhvJyd1FOt6KmymZJCckMOtUH2xl+PDdDi+09vDiKxrvV0mjI
8YBqUpyoHPk9E+fupodHuAuwoVvVfc2xL7B/l+j7PyE7poXWEPPuXhoserwOO2K0
5VbfI1PXidh350F1LWfYqL1XPL+y41Zdf9xkgVjAVcR9QLCS/Chf248thb2o12Lc
mt6oOi20gv7fRNLNnlAwniTk94lj9cVtIrVEVmjWHwfFs5dVN0kHVMysivfBA0ui
nbmrxJScZ4wA2qyA4274bGXkQ9WirhUO+6SqSsXk1aSkPzFWD7zl0+MegGvh8HUo
KGjcocbUQNWiAMiyHAi8QA9Kt74xO1NNGnSsRiIHaO/vIf/M1109V3ewO7rfq4gB
UIfRUug2/s4p23+vaVwx+oOJ7WaKw8gDMtZh0ryPVvYAkSydMNiFKTgRi3RE/M0P
OlEmyUh5p0v2Jgol3yjWklgMCZ/dwG8PbHY2qrh9KqDD2hD14fq8QBcn89IZCNVK
5kTZj6I5+nrc65rHzu75ujkZSsRFXDRxfKiAiicPF/2FjJiu12ueYII2YHRRUwvi
deFKGc+pQLmO72NvbnguG7Vp6JXY4Id4PJAouTHXIvqbgrqibF1SRE1WjCOFshdY
SyoPdqvB9h9JBJRauPR6CUu0c4uQEGxVoCrDVJw9NtpCH3VkB1YJTcmml7NUOPPq
n56/ytAClFzNOkEcAKqldfhP7rR/XL3gfW572yY+dtNVVGk8Z495AwyJMcaYVeyw
2b3/XwfpgdHHJiyZCtpEBzPEJdhx2OZ+lhYLhVFhXHMesim9zoSxgQnCOY+OCasj
JwQryx0ezBBezZ9vRfXQROwFs5JoJDnLX62uGN+pcyvMfu3tLOWhLDVBJfwQaIcg
HUD4E9TgtJriIhJRLtDzN+2yKlSGSRHdiC4uIyBa5BczZ+UkcoewJa12kYoP4inD
VhVUEu2JQpqBFympGRVmUNPTx82Jscj5pcb5lXOvmTEelh31fNxFosQ+hLXTfNAG
dz+tjPsYbi77cOKol8jwjIXjLKwnCBWtYMwUjtP/X9YYQfFLF6mJ80KHD7Scu6xd
1jXQMxzEz7VZObJ4vGY8AvO2NFk+L07X7WNoCCwb0F+wCvT59+BmzpNJjI/CB6hg
CvYt4/3XJDdloCCg9We+NNtlYgTcsEw4abFWWhRgGmMSNLBbGjAd7R06s5viICTq
0YDG7zhckTbbiQYjdGW/k5WZlle3OEKf0vtDmOlXuHm/xHRiGxS1I3pwoQKmao8l
OgWQuxt5nISregbJ+LYMRbHZuqksQNv6CZDvcgMBVWv3HkaSUhh7TWtH57nptHf7
sqIZCjus+Xbw3UbMgQVCMsFXRawQw8iHgpA230+xHoKudL4SqLFjn5rJtKmXHV3P
bf3SEQ2sL5FxAiHxdr1V61YkYIoryjGme2eZxNefYMrivy5MHBgdTNeA3h9Wy1Si
rCnntT/51+d+7llFEOTtEbEzDLJVpyTKgdMetCv+jWJXTJT9jx4y9zy5IRsYAQJ1
gjRCBPCR/y8kNMIzLus5bfyX+bDo2ipQgDz3KOHAGClwp7gYJGuiQfLB4bRpyJlE
dHzi6cgpuhrVxyuYUNkssbihpnXYmUjVLdPNXQniioMbzupPtszIb1EHV1JqMT7a
uSQof4Wl60qEVquxjbqqHt8f96jM3CelanK79S8RiYoB9C7qFd2VTUTcsbyJDSr1
oQCAS7YWGTaHqZ233wCbLRrihjTEVou5WBCarFTk6PbAqv4GHnLFy6gL8H5kOwpD
xSsV3nYKE0i5C1dp5uc89dNC8FMu1PsJs5fSncSpxjWeBjayUwyQ8GLTIAU2H48k
+gpo0vaHBfYI91xpVs6LWiMQSKLpHjCvA80yByGHHfbElCjlxrDByLMeSCDd/Moz
ZpvInrJk/H4EnghK+5GLmx4U/W80MRB8K6QpDj32Gv5VAvCYl+io0bhwWF8hPPlu
Saf4uKLon5OCqoW3BzFc7bsNV54GM5A6H93Cnng1k1EmQMDju8HRuLnPBjQrAx+V
GEHyNFVsGr1M+0P3zQgF/iUqyjQYFh+Ev4xcLksw6D7kvNnljFL3W3+ynQC2pF7F
dcSVekokxSAZN63YKBnZK3aX8zJQ54JCHNxKUFSJMB0IkLkSrryIeviudY9b9IdL
Bg1x0OOGNcLPZzZcTYrPp+mY6UlY8Y0aGpRpLl2vUHFXs2gYVmmyLS37LiLI1pOH
kZXvRwAInNOA8UK6xLl7tjKplkKpo7GpnNxrgMj5Ei/bkjguJzMoAC/p8/ow3fZ0
EkM2MQVOOCrCGEGbb0GQWnovXZ7q1rxpiZeI2Mmx/p9iyhnsbyhtBONxKgt8hMqJ
gZlst3qkWuGZT3UzoGQi2JFTNH6H+gneGrXCabsc6ghNFrbJsSlCFWcRj0VNeKM7
9lW1mUDuwGzDFI6ISbMWAdijm+GEZsJz3cM04GgGHKFkZTfrpx/ZlzYlELLIEkRH
FK/VSo+TntUpSBnJ8XAwd18lJK9crkgTkXAM9nDwXiO/lilRA+KS6KVGcUpPXq/k
CdSguPzmQMat4ahrq4fnCJBMb8alUmzeZKCYqRQsSkCnq+bJ9yxAkwZ5cY4FPTLk
t6NJx9h2IzTPU6FPzOrd+g9jEXBK6FG/6PsUSYTBSS17PRe3A7aIFwfz7sfdYWzP
RrWnGFZYNhDt1CianEUNBbSJRdmkBfd/I7FU/BL7ypnCwoV9j1ks2WMCnanFOZ+V
IkcMU2mMIZvEVe3zSiwQ5/9n/bnJ2Crls/Y09Ai2m8l0a1Rt8o1lxKvTDwskGSou
7Fv53hACSTelmZ/VhSc/qWNYnmD74T7CuepCEGcJ8zAtiFrq5Jg/ynL1UB3Sg1aD
lmNdRJAHP/Gbf7o8sDsU6BmPaXTnhi/UNtWd149ZCcwzSeDH2ewPuMz7e8YKL/E+
/2cNERE4Zfq7/yF4lGqcuziSCMUHbNgyuM8+mZPbfQCRQYLfNF7PQpOKdSmgw8xO
jnd0iIfC3dIUmVVTgZKLB+9tOpky7HyvbG4YY51y6zFgFam3ojqqiLfpkMpQQFrd
vA3PDwz6SqJGioUdgoOZwy0oyhPoajGokWC1mccJImsh/eWyVEtNzjiog/YCyVzl
WTWPzxLyis7C2H3OQkXsbwcieEdlADB6EDKixUqikA6Di3nJT4EEN12FFY1SAJWb
FmFed+2jeSs1s3MWQ9f2dZWUJheZFhxC6nGtfgtN7OHmCKLIIx7j8h43UqrJoyr5
2DlZ2awqKzwCJQg20NVyCXWtZi9dVHO4Sq4oOz8ivpXnOaD+W0RHP0MAwzeWFJBJ
/PYMHa7XKcZeo7+40xdzmMeiUY6SME8M2gEQoIqq8HsDBTbO87bJrZPObFu6v7MN
U9kA8kNfONfbX1aV/1vDuVu4w8W99fQDi0rNhsZ5PukegRsD6m0rkzydNn8z0cbx
L+zv5HCLX2hMUgRdxBPeLRPn7cz/2zgWMQZb5hpvv6weqPTvhb4GfbPomk/6Bxps
QaVeHzYgbjmKZMOdYiHszFJXM8HG12FedW5PWSe8ylk9Mh0HrPvfHxMs36K66BGx
Ha88bmBAb1Rt+Yist6h7WbxdYckf8Ua85T8LyadmNGAXnvDgnU3OvBhVD+JouIKm
jdvwT4sOvLg0ZQEiBrZTgRXme3WXE+egNuJE2qB2j0ihI7A5V8DPO6Dy66hJBfXE
e6xDHNlu43UKVZcP3TqlMxwNCluzHDv9xaJuqPC/YfHgxTlO8weXj9LTGmbjITId
hMdXa6LsjtNOyOKEwnThQZ+r2L0yDsDvaHTkDZUv0vRW84QNKdKrI23dGnQNXO7M
KyzG1Y7Jz72hKEYS+txwMlEBU/oLuH6jqoFSLptm+HPOoJS1KhT5ZvHOix2XZ9Xr
OB8sGr7g4dkzNINZYDe68MHS/0U1kKpEwyZ0wUfwFCQ+f2mlACApUicSGj9mpTwr
wQK4eknyBNe8JWJM6EbEj3c9OLSEdrvMZMFPkEtjNNBIIH2dmDI/k5UlQAmqnaC5
OMn3YMGXPh5muQsInLjUAoNgIT8jZbeTWLoxSvyJIG1vJoIZ8SsEbtD+Q0aGBgOv
O6tpF7YGlFfo+yJhL5V6bai8kZf1cwfkKr6i/R7tS+8jp/e7rlsyjE1ScdW9pWCX
pXch6WWBleQLJfvRfB8wB1sBQrZ7VbGBYX6cRjrTY6Wk9zY0bjaWoD6SYNNKM7lf
xZyvqYZvOX4ere3X/dlkAyT2XGm5XqO5GgfX5NnCHWlpou1AXjN5E3glhiWUVdfx
89PeDCUNhJxKbPLYSg7tjn7sqsvt5DY9tyBTtbTEVwD3zphY28I2wORb9IDN5Q+O
4+FsazQvH4Wb0qnekaQA6Ju2upgOLHMN8h38wI4mDPu0wUCOz07FUni/yxlz4dn5
u+ne2vJW99tpQ9waXug5sCltS1/1iY8yqmqw4xhaRN8Ja1yrSh6tYoSdtHvsbRU3
Z6j3BREDrbT/xMhBtM5B7Ch0DPuq7r+eefEEIsh6YUgWEFAYaxmTr/TlwPPahmTy
HKSmx2AmP8C9Hl+0FFTWy+h47L4J29EvPCEDeWtwoCfKYf9QiTSd9Tbg+sDh7Ygn
vWqgwLO3eirvDdcJTWYq0UfmmmlBMtUmlCC26DOeltGO5nM+Y2GjZ9HnQ8Va8DJC
ANrIUvfcaXuX3uEjlqNZJJQQno7lgWES5fB3lrNNn41IAsgbbsaBx8uccKQtNd4W
V86z8M752Xlhn+CIlYytBlBO6aYawdxJQcOcJOpKe4oCaaR0U6p9/TsI5P5nGI8e
/W7GjApxAqEKnDZQGjFsjCgxGogkjgqkBf5xlkq15dAkmLr8ws3hCBLuFZImVqre
2V099M2l5v363tlW+Uxy0uLWWMu/bvDxEGNLxPpUy6TZKBHp4IY23Hs4onyI7Jwz
p/sQns1y+Zjvobvt0P0Iqs05kDAey674kW1e/sFKToxjydj23LPly4ftz29d1G22
ztbK/LFG7a0I+oZUVfIkagAGDdESqyeOVnDGzEO3ADO9gqhgjYaH2ytmChayOVE0
XmkQMsZyvzyUwgq0SFCK1pTaRE0eEnT1q1TByxlwfvRhIzwZ//C7YRoTBR76gTcL
pEBeNJQ6rc7w8/OdYNplIwsinXyC64BurOjlUMF1X/fXFirfvGKm9AZ3YDXunEoH
sMhqexkrc2Ga5FQAcvMi46YjlKIFE5ubn9g3KcgYYopZ6zYf3sgrg37sKGw6qDeD
ser0wpUHGNvNfWw0oJwWg7+oS8gLuqN5I+zqgYfxjKW1MmeUUkpuwhDXc3Qs8fWQ
Bj26rE6meU3IDBlrcCj1nS3MsXGKtf6AhgCQQwSOclEeIxzvVrCqRv1ez5j3DI3N
+t6iHzoHoW08otRTm6ySfCTA5mg8P69hf9whPtqvVEKjHxCbddOHcTeoFO7X0Xca
/9BWgorn+cIRv95CEC0WL9ggJRqympRAATuiEsht68MHOeVY/KOHBuEzZxyVybFr
ui7ezG/g9BzqL0/c17idxz+c4k85xncx9FP9MRfVnkPEwWflW9ptT2Vkn87pMuHp
M54JRwRx2NH/TkaiwrNoqnpSnpv3RfUiAewy9hPdDiIzzfGSOFa2NmG3wzpVnLrK
dtNLR18DW0b15A64QwSAJpP0D6jSnsi4ykblGB5bWXao85R1VKqBgOrIDRrVB3zl
8Rk40ICpykDnEojqCxDwU5PAY1yh5kYIhG87u/bjomalE+5ccx/JOMBg8cU2F1LL
t4qiz8L28EV+fIWLn1eY7wmBk2a737ODLr8En2u6F0/VqvEEnfx+YHPZ5Psic3JZ
cFjeBW92SLp1LoT4NtAhBfSQFZMP2T2CkNOCxsIZTKfHpAH+lmgTt9VSltlKz547
uGdznbU+SKKts0FTRoykUl1l7oJordZFHL375v6ISIAQZ7KwBOaPda8AYBJc5+8N
CYJk65BJH3Iu3ipLYRcoHrR+BOpHu8Wsgs6XuDmSei54gQU671Ccc8rLXZ6SDgze
ckcW+tWhf666hG3BODJgWxXSnY4uubmfPmi2ywCPsxi4MphTTodsrXUy2oa0m6cl
VKFoE0Kei53b7s1S0slSVXs6UuBSl6UfLz6DGcTgLLTDsdlM0lNoI8GdU92OAJpb
CH+cry2GlsU9Cs4LVMOLwCrtknVoXdNXhXeXUmjipwFWdAKN4tCzAzgYxnzjHDS3
U3l/NUsi6ZLVNAvbaVTKB4imE0ENxknbRPSIMaNKVpzeX4nXVAB/z+gyYEliAeGf
zk4nbipK/qwg3Fm1z1VB3kMbK+WRPd4K6O5vzLKsjy1X4omxPNrm4QRDB9d4qvuU
rzJSTxqYjSGS9dGKLFdDAiR131dp48/Vge9gzx6Gu7lsIszYJRIc3XvzUhvAiK+i
L/GeBKNDjZ6fKvsb9zdUcVWE2KWInCLMzJkClnp6LDAI0E1GnNxx5tkcH9RkM8k0
t6nPUKh20ET5v5corX2tDmmBw1p2Zs8VBIX3W8bF2p9V9wCeUHW2oQBpQ6vki+DI
o+bSOF7PVoQaZs9KQYXfw+tvwZr+1cs6k+DQZatQpOBwBGVSuZCCqz5thtHsAbKS
z8gm3i766Jg9C3Xo5xALec3/EoZOQStcdlI+7Y3UNqNrvd/wc4Qfw3vHSW7gFvFH
lTozb8C6977uwxrOFUnSV27Fcke6q6rVhosuIlk9QIq72wXGGU0UIxEtXq9ZhA1F
qn/VNJhK8bhAU2E6h1YOYCk4DbcxGOMM9pUHzAruRIEE2tvHGmsUMMaU7ueUk50Z
g/pbCgjDHa7Y3vCrW4wNiPk+TM+nIByxNKVCEjiIbtEWvOJhczDwejxcrQWO/ZJO
kHe+JoDRNk5xIkC9WkPT2q7atSZQd+MTvqzEU3CbbGX0FZn6nqqfJkbS4nJjpESX
GF9R10I74x52OLWe8D8Sw+bLZG2dYsNIeIdrV7v4FW/xZ/gt0POm0lB6IgvKCj1F
MRAfHK3BmxoIyVcxqgjkyx8U9numKcnQRVI2k8urfAzRnn1pBervKw7E9ynS1jgw
xVCZgkk4/XRCPpBeJ6k77SAIjY6RxbH4X5M0kVf/125kF8yWzPhCllHDBGxM1z+F
vHZHSgB6V/+5kG0llvQLdKCz8AzlONjug/IKT0pXUgXwsRkQC2PKO/2xQgfHrltQ
DMj8AkmvULYcLNwLKDGAt86aARILXDrDLREAyl/djKi8kTn5y0TeXvRUc34m4FGO
OAYJ3e6XtXxGsx4SWUNIMxhmn7L90pzTJVjcBY6BpZkwYtxcqwkTAPvhl/WUBMEt
/hTPBoRr2vNAJCTPVpWrnE3JQD3kQvcs0dEBs+Ycx0MwVrFvuO+q8NqKrm1/byN5
Nu1k/i5Q8AQFKfNqfg5yAL3Rr+8969q4YFqCQsysjviQcI18TKy9QRBEG0zLRr7g
+bmeNNBODxyjoRlOjuukuHEo//g9FVBgu6XZNUovK7BrBqSaMBUQD9Hjt8Ay+wNV
wST2oKGoO5cu+Pf/n1j5nurqSyItbMkzWB1PMQxoMKuXMgo89H5zC9fvkts8eRCm
djGvIl5527CkBkJphS663eVv0aUEh1FUDwYyZZ9pwbwk2weQB72KoVNiQGGYX++c
sXHdyQUUw2o5aVH/qfkb7lmqN6oNycFSTlurVxbAMXljHCYNQvHOyrxxCcvUFI7v
f43NpxiP1/0BMHCY4AtxMppsdI24cSUT9IshgRfb7Njtsa/YAdisQ0f3y7ZAaM0f
eNedmsUagE9TJt1xPXc4g+Dh3qJZSKDaMFMBUEItodCZznP+BoKxTwKJ6VmbSgOY
W2zOcGOnXB8t75kX0TRvH5FNsazsbYrHM6EtJfOt8JDcohpO4UsGIfY+aqi1eyBg
cusjL3zvRS9/9PnYk1t089G3x49W0b32cyoC5ASLb8aPTj91onOkmLabJ254L3pe
xpZy5hmQqLlThCgMNx+S1+7uRdErd4IX+U2aWeKgTY9PD/sTUHjjZVWDKvPuE2Dj
shbp1U2M4NuFy+zMn1jI3FJhdgzaUyDq0rLIQjqbPbh3s0dIrxuaMv2cbehIkkkE
xA/gfZtgeNSxeXuDBVVG8j7ncFkd9ULrgOD6lJUAcEjBhA9nPnGYtXdzE+MKruHm
OgmAVFYlaoCkaxFaOfiI/Pxpr4kIsZeJQx5J3ZnQDMao3zP1JzzpF2TUp9BgIvva
xK+ZMb0wNQDnBKfToxmNIytuhGpdjDP+K3NlJB689jZFw+fdhZjcx3J+kTfMZJE5
4WSZppTk8OeNRhGy50swIHZGvSh73QGX54BA1la8fhm3p4aMz7G1TdHKl9pPzD/L
V9IFrLlJNbMkgGvNLB68fhGjlvRIpuRElkotuiAx1R1O4BYLJZff92lMK5AtwwQh
W7bGdbNaCcxcJjOhhOmQPG39Vpd3BCfWiLg/Nc+AQZCxX4vPQ9dkN+Z331rQTV7q
xdKCdafNfxa1QZDjv4JyOty6MqNus8G6qmghA7pEw0B87WmEokN3cJAejg6P/Qk2
eQ5+AE9cm2DWiMKBUoIIQLu9DJYnU+s2BUdraOHJgjveHtVyQIm5iz2lcVYjKP1C
ckx6MLWi5v7wmFY7PtcCn7tBaXgliWIVWh3Wa+dUaLBCGfQ7XHhDsOK8StQQOkkA
QPrDZgxxoRqcsAdSv/aCmrq3JmM42xnieksIHHbSb/7AzvhiWfx/UIEvGRIAW4XW
edkgktFdsqBolfMtlp8uWWaD56kodEoUbKBpTyXloAhoiiHci7NjvjY6vNq6Bc4f
fYPPED0G60bWiwViVjFh16gE9ZCOOvs/QcoYRvf8qCouTGewZdRzbHO/oesC1/Ck
6U3u0g2In+yn7J3TOIDmFSW+e5j2mT+2sIHKeqBEF2RXIcUqMcj3cdmaV4pAzgg5
7tgN/lwkzMbaCrtSmrK7OytoXskuWJBVsl/ZVDGf9obxJeYqeijyU/ipWFTWxhTt
9/aLn9TpFWwwylxQ4rjRQiHFzkW+F1hHBH3N/4LTtjxQYHg2UVYME6Q6XAD9ZVvm
syfJrtvedMioKg8yp9sNnNiboAC1AHziDmVH0kXk2oBGllWCvDnhd4pBnkvv2dqd
0jw75VSnzhTG3gnMR9BR9FLZPmP01ubygXlggqwMk9BC+2ex/sACPzIaFrcQvg9Q
9up/Kd00qpsh8LA6UOOZ9gHTBfYVD1iWb1qNpV/k4Qqr4TuC5jGn5c0xDrEPTjdK
j23YHJGZASe1aUHmkpD/eghOnQ7i+OIEQAjjzGadAvt98aHgryBX6X8d9OQVptqj
iAqz4c/HgILGxJmH8/dG3gn6/wPKtH39TmOULRiH89lUCaJL8D0zZHgF7Q/TpnjZ
mEzEvg6yf70USRW/Nhy/+KnZWQolFc/RRxnbALqA3dDQdyBajtTKU+sLi0T/NWJQ
2vcWCZI/XrZ/Lk6xL+itzaHa5xR11bliqzg7aLMgMD3FxQKTetQIv0lhl17LvNbq
/JVEozgodY8hMns3NHSV7r1anB3ulhyrIpQ1sOlbfhAArwZmUDtTzJ4vdP/xNR+5
jhkXZAg9s8KmyeuYXHy6TstDNkb8ssM7au6/r6sGE9LMOGO8QCXK8gtZhgwV2tLC
I7999RHqQoZp+uQj5AWY1ynerTQLiRbxsv0qixdG0j3g7i30tGsIR2itJioSRmjn
9JzBhPsLdw6xpGJeQ5Z5arSLxMye/s+rPQk4dvsDRoTcUQQ7nBQvKwx/CyILBiWR
NlvKCTZ2uLWutXNGKIa5USTdX8Sq8/fz5Fj2vN19Fr0kHpuRtiv6Z/ncIUnKU+RT
gYhtSEbb6JiEH1mvwDaOw/x37xIMUqkwQ94XSmgNfnUdQC/YWI0jOFXUWQs32ENY
kuga/PXmxl5jwmvVgawrg3xVs6pY/Romn5KsHaaIi5JWdaYECSnmVZd0yQUFlivz
u21f1VVDo9AMEr29/CUUDwjLuiTv3Xu11VYO8ey/XHJMrTFf8cLppSTpkJOteEvK
VukfbOE15dEI/GG1wLlOGXAoNpWIULJa4aBZeABxTtR7CjQyX6l01TF14ojX14OG
7XidZA4nJU3FKJjoPgz5QkcF0MwQNrgpVNaMNatOmsE27CRqYeGTvODJjggDQfkr
qxXfv5eUnfEUyfjuOPDuzHsPQkmPnbMr0nba6Wlng9MXVO6nxvkUcqAa9bGWNdB6
OP2kXWIK8wQi0x7NLq5b+s51dL78oE3Rh8on1ttjW+wqt+xKh4wV3yQCp3FWlFRb
JCZKV+i2t8usFbE2+P44/8kA2bZT2BLvxWpRTu4D2ApnjiBL0+V48sODjX8i4xEw
wbfNA7YnKjQCOTT0IUZUtZ4Oi/L9pogwe3OS0MmH78tG8pMUPlah/pVao+RfXGC6
zP7LbaiE8sZCR+QP8R6RkYQ2i7fCGP8VlnSQ0166WrLX02MuyvrzpXuxsJl+Oz42
/J/ttVZFTp4mPifuu4fYcnSfu5nxnxBf1uVquJjv9A3wVCIGygr0YTPdsKpx3/vh
siESumIBeP9XOqL8BKApLECSIM88sq57ok98a2O6jCATZ5m8/n6zz/aMOih0OREG
kyvja82dBq29t4WhzTPMJ/wnONyh/IRGwJZz04uJPUyIdsnST40vYjJhJtJE8D3Q
rb8ejXP6R2T05cwDV0mAtaXVclZNjhCTJT7Aj/L5ol6CEUqOV/RM23sVBh8MWcJY
JVUZ4bwueIeVksIApwfcSyi7CGXJb81j+OceQize4KDVAFie/k2kUK4x+v5neB45
8TbHxRWBo/ltkJIafEwtrfPeXTX9OJAgWqqHhCUgUIgsn803WOCsOOXaJuScy2u0
Cauc3q9wxvzOTBBjAmB0PSHxpbkfuvSf0LFWMwI1TusLLsU7Mw5vIU6FlZQtzhVT
HhJCZ+w7wsE+YLj4GCryXh92s+CQg8mIo+vClYMviCZirQiV+gBsJJp6N2pQyowi
YJCN1RBTnCaOtuEulx2Z7oYFfFHYdDpVAkHRTuFh8FMA5OKX6JF76pUdgfgfhwNW
Syer1jJ6CMRqnvW8RdajpE4651yChbksY4E0GO6O7oCEsXqLTdTDpeZI8BMjNeEF
lBoAxXA9ejmj0wLtCBFymArGsAodfz5OITt3e7/xV2Z7or1+sIWeyGv755ydeAtz
ZxBIawP3g7Xn6r3dURmrEZmmGi7p4mACdPajccudyjU28cwPfEu+66xTWVGmuhk2
Ry5G5liC2tRtw3KYQ8bjbM05MGHADbL9vZ4PS8w6Uqp23humMmBY/22DgevLmo/q
Gp+B1F7oMIsb9fXh+hYFVjzBRrIBY1CwVTPxK4aSKRhCmfhMMqqSLrEp6QnMuiIy
9eq53vSIF6RM0PU19YH5WfOO6ZYfEfwu2jT5qqchIsW6kWc7DBANbHN7smAAOaSP
pnIgS7l1fIV8n1y7QZGz8OgJNgY4HzDDpRBjkX0J6bXOlIbsdxGbh2ImDqsZqYby
9HDEFYVX3goIIorirI5H52t04z8672rIB4cLZZZc+BnPpSwQXWtWgGNxIqM5nZ4O
QRjboc+0Std8y2ZmiGyKS0LphlWh99vr6sgP51w/fIxKkwKh6I9G+8hkYSrHH9bE
kjJGO5cUf3Tdm0tL+AyghPRhZ26mTeG6pehudrkPS54xxvqnBUDRJ37py1D6Xkll
EArkDdlYOL6B5lLo9aFVwGkAD8z1iLXN/13BwZ9roMtNCRghJg/hM5TbXOjLl1F3
26DVIZMyJwBnZTaF3k3fkpgfnFt+xrkqtIq0DgjT6bUT0xYdK+mAzFKtf+es6dfh
cTdJzR9pnU/XAfu61ZCzNyk6dBBASeHQCGM0kjvM6VVMCfrEAOZLFxnzrRoKrgQV
mvv5EOLSAv5CyDYZ7sMhvtqVnr8qZ50AQHYxD3MnYUb6k5AquVbqUJUKSDhRZpI7
dPbVTv9DRpdxUOPFrN1WXEkoLIMXcIv2wiTPPWlrjqSYkGIpuva+nKh1ZNGTR4xo
AgUB15uO4Rw7w0xvZmX55Y3irPUMzQUonCKQ2H+7KZ4oJc4nBD/HmjaWMflhCh2t
mPk8liSccy0B6vj3CuzZBfuHF1llge4P1ZmHk6QWPPwGXfzaqfIbv7h/1amSrRKk
iTLjquTFWfEYUUMxGkInJeZON9jphrkFsG3xzgpKqm/Q1ymtxEpsuXloP8mBv42g
sCRD5qTEJ6Z7n+oTknsT08Up3L6W8gDFduyisAu+Zx9TtCZsyAfj+v/Rc2X0bx51
rAKTStUAwpHE1oVsdw+pYiz7pn1ThIFOjwKys4qQTuuBSrG5wAhyorte+0tCdeMR
GEhjtUDzsQOBvLreA+T/vWbu9x6d3gOsZcBylxv0PMxwluwAu8HA4Q0PjbPM88At
3SL6wplLLDpno7ZkVksD8ixzVoAWImCf712OwaRfSh7NpGTG1WK4jhdCBZTOwrNh
mnCvzfCjXFZQdpPrfsrxJwpi2uBfOm3VM8RjMEGhcUYeleV+rjVs7pHgVDv0FoWh
uFFGTg0VajLgbfQjYWMG2kGQ6my9SLl7qvcg/zkTRQCDwSgP9V8SQzYf1Rxz9ejD
+D+B+6mUjStrDVeVei1daiK0qSLkhW9zxeYkX1SNt4DE1rhRqXJA5wsL/0H122n3
fjacy/Y14qd2+1qedU0g//B4bH2JTWZkWPWcVW6K1lyJG9RjK2lRZQKetlGTGYQ4
MjW5iWwjuxuCL32YnwVXTZDBH4Anm76NHJ0hZa4ek6FL7TXsiLOKpV87itVsKKBK
PxKh2kB14I8PGyI1zw2wq0t1ezXSRQsx0I2LWyBFLt9s/GQcZKjmy06+W3SHp50G
MBU6x48fknXJ3zCLbVrsSwdY8N6q7X24B+8ET2wB89FHnrfyOPC0suldGy/kR84n
YHvZqbqp5c79+8gkOxyzDYKMLIrdtzCk0vwjU6L4AN51oWNjLePPSTvLoIMk2UFj
oC6qdidJNcohnPqUOCESsNQALpKiBYSH5uPb6IfkgDhCj0RPzwm8rzk8HaQAS19O
CDSm7G3aVgCP58Coa/8iGbM0l2DSs+FF4rqJBdJK0nuI37cmyHcCwIOGPArebJ67
/bnQ5zVZKuo68qMunfhMVljMJ6vcikQtiTrTYHQpcBL9oWPmAgLDoKTdJ7mDx4JG
OUaYyCZ34IS80IykOgja184TmgLWI7NGwFZfQ9uOywpLKK7iqd005g6gyvXb810y
tneg1tqLlOlgFEL3pFyg0tUwviYZaxfZY6s/XxGsIPHV1/CjL4QlhLkDXciSgLDe
XTxuLZYpSA8fOMEepN/R0X/wrAzOpywrT2iZshDKb9FY79eVi/3mY+0i9Zgu+MkF
1ZmaVDjz/RF+KG+gSoovM9mFFZSS7rV3iTaVVW+evyZIhpdLR1CLo6GW4SUkJCzX
1VlwiAGaCSmzus/GGzVY8yoATvkzVzVJHMVa9+LadsIK+TuDeVuBTMhNjJZyx+7Z
FDgEFjZyhuKvVbyDQ1RW7rhFzYuu165eZIUBKQnI+XtpiQdS+exX9ZMZM63MxJOM
9k9BbcxBFSYpigo3MzprvCuDE2dOKo2MHSqqBCT6zAht6Oiv80aro7NAbJKxAh+c
QRHbDd36ynXm3DYULV3uG9E5dzwf9ZEzasjh6g8KB65fwXX7vGnnHHjpS+h/xgK3
2wIETk63/kiYSaaDqcRswCtRCiBlPu9/uUU+1WC99sEVv9RvXN1YIQZnxstY8/dE
7Ay83zcAzvATl1tXtaLR85nPjXu0ulxtg3CSiNVdYmA87Ao3HV09tfjodUtvH6ps
dv7BaooizyWPiNzvgBaD5rVnjdd/7T0J+xtsABM5ig0sOa6MV7X2vcLR8mqigYzL
xqILeCnqzp9apW9MAOAlOlcITOezTy29iJjdX12vunLraU14PTxiiBHvDOmr7GzU
v4PppXMzJ5+7gILSfRouG5v7QuJ2ON3XjkzBk4124qTblfs5t9TbK9kRU/TnvFtc
M1+vlKUK2zzXbSesSE4UajLknF5jS9M2dS+rohplnAYvIYZU10xXSlpX6svElXYD
ewGU27nSJhGvjpc4+Z1Nd8WdNqxhuMgUvfMbAc/s78L/eMr0wvrmCabKWJ9CipMC
c9vFIf4eB9UICOJMsEymRDEP0+qgn8RhFPp06vXotSjpA/ysjmUuAgVkwnePZ9Yn
capCMs4nN/tfOXC1ZSCMvfOnWTQr1Cp6ina7SHYDLjW7qogRvjBiUYoawfiW0PyI
5ntQ7Bt5lEm+Q/sW594oTDGYw3P4PxNAXBV501CarIU86hHdftE85HUszDHxtadJ
poMoZGkykiSeg4ekssA8ukW0A0l/3zW22CxftKcc43mfQ5JTmf638nO9Vw80wmU2
VBMEMIz3g7WZ+AlRRBoj4UxYzYsRgecHsYd35+bce4uZqAFZDbGiPIN/asS6lAHQ
UYHCm4eZzBe+FqsRrie2AwhI0wRlXSlr8fzJAxhDqn5qIELPNeVhUPDuC2NJaQa0
FnjL3HnXdpZ4UKukZqhF7PE+g5SxfRHPnutKhOIwjbMDxuE2LlhWkYbgPGuOT1AH
wyFTy6HxHpB5a9rSz5iGvuele2Z50P8wab7xpdKeGkOD8/Aq5493rTcCJCLEoa/Y
RqcLAUsoCu25PeTKMes02SmQGDocPBoX3YmKEfF83fASNzpFYzSE/QsrfndmHCT1
6Jfr0Ve+cYHQr9Rpn5nbJVxwrlVCWVOUuCDs4vNqX+J/1FN4AakGYNnKbxoO0R1+
XPOIAZmtUcXQN++H7VPLg6dA60+emHABUL7eSZMawiGUhGFxxD+Wu5vAOVkcs8te
3tdNNvDYPuyRIGsTxT9kuwPGmOK8xywd6hbMcdh7b32s2gzl6EjBmstC0LJnigKY
4KUCGVhPmNrZtvTBsSUBPdLtFQksRmFX9Wqa6WJs4gO54ib/Wx8xTAFSTUa0czce
mPSQSM8zuGAFmE1XfzBNOf4CMtpyDOXZ/83cSOJnCRELYxZMWr4C6aPZkXonlnO5
AUUjqYDbjSRPH7xKIfQ5xXAp5hCzXEVqVOTHLzEq2FTpkDTFsAo/c/nzxvf5L4ba
QgPXTLwzASB0n/WgP7FrEnayKBaUVUqFFEqJT7vgXO7ki8/b69cobs8JnmNIDROA
gDj+V9/zvAzTy8vKGdSYjGDlS5sS9BRqtncfHiNoDzQFvuOD37uOr1dDx/L2CRee
H7N0mI/s9dnrON+gnHaekiZMS3NatByhlSN4o4TMa8/OcOFlo/h5g4cUOBFSmDl7
+xmD9pXHOMSTlEFESVajclK0cwKsnKFPkggdAwg+yRAhFfCbMDIZzWgk58vXc/hA
yIfbkpiaPB0jlgOaK7Jb4uziiE3BJVeLNN2MQb0DMu74ta7UmkS0Zk2suKZwcoYM
6VM6f7XlPR/EAG1kb841pzTN79HSubGfWJ+eauDVMSj+dXT2h/vjDVx6Xjkx/qqV
EwCnLfNeA4uYjf7sQQlsTlcKp6VoOlJe3r/l2jUIWxeCYGbbKKSG5l2HWce23J5l
pdb1K+2h2xdvgxGAnJWuFZAGW46rb7ietaw8qiWBa/Eks89M7NyU8S75FXmT7t1S
nlFuzIi0WyI64IVzPqgekjRD6C3sqxOXZkH3NIVRdINOWm6Kj9wiejwlVIORJ6M8
s72EX22gqhE3Lvz/m10XqtLqBfx9MVzmBbbNBeLyILzgvaQLhyrG2ioQ7WgNq5YF
++X5Q0+vQ286EwLLLzLEWqA3sYfxq6t21gps76EZVezsDEcNm5znyGjUO1FV9XyY
oB0DWSBdUH7QB6QaK0B/rw3HL8ybRtFcH6DE4OSZ09gBAAkUeAiMYQpku0naz010
t2JF4nqZ1B0m/G8fBFiF7ey3gDQ6s7yGl2eKKnnYEu8Y9kUERgNTWwXhCCL2xJks
Aqx6u55iFY5TTuc+u4sGKQ9pAKSsK80zHBsF3wq18VkmArLAh7Z0KBUGtpzJz4f3
jiBOQ8xkAlkDVs20HD0x3cOaQwr3DLOgFLjFGZLzQfL89NXBf/OtrHNwnD8uT7lw
4kV/SItPhkJEwGGXRWEmcCD81cDc2I9fSqQuNltS4Mm48H9xK00bU2mBOOXD0jqk
BmpONcvTn3LpV4nzc89fPP5fglwHYCOH+9Kt4gtYzU5zwlAEmBffnu5PhRIA3Im3
XE0QFd7hDcIvwmpfcK5bGyjSQ6nf8qZ2HgOhyG6cBF2IjNmtkovkuQxdG6lFQEvS
AG1cOP2QcdxTW/c7Zdj72aa1ESQ67ojnJhIv4PDvY2XylC/3+IArzPEhhiFgWFHw
NkWrk8i6JVWJqOgk04M0O7lLQWHMnts3aCP9Gd22dRYQHrOJNalcqyuhGqtwPjDu
MVf6uBFhON1e7vr+g4oAbzuxF1fR/GLHGxXWsNqbwMfv8PdFNf0O+VG/b2ojZK2v
7ivpQYepyL9bK7/UzZbL1GhCTgZ6XkrbGKhSSTxosZwvBc5GP6P4iBs8++KO43u6
dkcF6t62pADXuwoi4UjiitCyASTAI8uLlqGxA12JeWzmlB5JVdXLJjBbgARQ1PKS
nWkATNudYBLk55Fgl6DcVSH2S3wdp2Ma7jx5YgRw8gzv0KoR4hio8vA0LPnJ2uvV
GWveeaSdHAgvdeMiHAUBPJ1eiXnPKXoRvTPQPhD5UpKaEDPSf/PLs+7JDL+FC9zh
q9qCSj/DrjoiTPyxPTxfd4iT1QwWzlDAfEAKp0ZIY8Bzb8ObKLQ2mfsRnD58yI55
/eHxgOeXv72gULxjT7or3lxaxOCX9/VmNTNM47gYp8BZZELnNFchjjOclJJSHy/z
lzAE+on2L1SAIemM4FmK7pnue8I19mRhAEbHKZmTgPbRhQwQFoBr/ScZatWsIenk
AnaQxuLkEIho9S0j1xeYQAdZxoKeHK3do4jH+oPReYkTQx/26fMJKaLeDudXtDWx
PYAkVgk85tu8h0YxCx1jg/VLv4KFtUyBq97v3o7GoKwcrhOn+s+hVxc2Q/myL9Zh
+XAWe75VNNxgBH0bA/b/1RsXlx+vp1Rd9UI20d05dlHzP6hQ6HkBuM4pPP/+9HIJ
BjaU0JpMKiBxIe4AW0sw7NL+krdogKSrG5Hr9sVx82UdLwv6kmIvawpVgHuqajBy
jBDIe7g6lF2oqJ4+ynjB6hO0ZYBT5JTvxxKAmX4fIex5g9Dx9SQlCpExGV5UG25U
9NpbBYWFZCh1iajUr/R6yxUbmaNo94dsNOcywzVE9wK2Zmu0+FLzvNOhA8s5uQCo
ZS4cV6oTi1/paO7KJu9bdvQGmU6ywMqXXkvr3oZ510qKsKqsbuyAvWqEccQGq1Wo
N7kVdr7PtUHvieGRtogz6b8rntHNomHFVNO6JK+Kd5+ow3laplHBMcy6GuhY+Ekm
kLgqVEOlqKwY1qLEGZwfmQ1ZB8ursAdNZa5At3rB90eTSRgjbUoOyu8F0o4MqOwy
GimWSh9zmWnhf/jYapEw+nkRIFcvQx8Sr9KJDM1P0L67+iifFcfsjEaz+TktuBrB
SkSPU7sXApxZ3eWykOpuOnTehRhXPyGxBcpdXWxCYMLTMsVaYUgVaT6WWJ32Wzqn
Us2pYC5X2J69T5q1qBNBhJSE+HJve2LiHDWDYrPnxOqwg+IrmXN/FB1yjCtxTxMg
c+VsiViryOsBp3Z6tGoQRVg2sCmCyO0nizYHwJeqqd0I9GNYzf91zuwL2n7OoUPz
2ZzZ7UxH6JqzsGMviidmAfp7y4OHDCbQGG2yu2ab8G4ikKsuT+xAepe4EbD07WWZ
19kyR2+qeK/ftqJ/ajamB4bUIcVL5pm0Ygx6h977D7JMO6+9SRbDEz1HOelCJBYC
QvKeM1uEnWLx9qFDaeM+1JKcx0kjolcUKvkIa1Ut9AJiaPCH7GJk4Q02dhhCVNXO
M3NT+cC5SJTs34GFIIZxIktemS8uKTJHCw8g10QCaetHFppTiTngmrt1kPMkTogI
uMNNvWWIKmxc2n5l9QHBZZfxxUf/1dSup3QbtdiN3B9XkqidrRcjZvLbdH6b8dIu
uyuM9Jg4kGv/7w5wzRN5EeSg88NXOPabmDtvwPE3b4nX4wyntqtidZEQKCNSCLn+
E+3IZ0xnzth10CVGLb/9nTiPTNUQHT9iqCfkcMx5238ZFeJn5C9T1zVD/p7BpfPf
e4l7auvtGIuSds5VAsUAmlrbwvQab8QBUAkrJfSHAVLY1+gSrlLtyzaQekRhImhX
SBUksng7k/u6xO/nq3mZdxQFUm+lqcqJtknN4ZLknA8jW/l+9a8v88xETlU0r5To
cv91CC7Y7K7Mf8T/o7wmTMNnXoVI1s0Z+YTvLv0n+GmB1vD5iJvSHKR6gBKHfNq3
kDk/TjxBV/LVCFu072/PRQ/2muJwI05ZeI0MoiyX+jain8LXHQt73/uSQgdd5dvF
CWanQb9RH6IPUpN0o/DOx70Crf8RoKpPqSsnoXTo2Hpvgsuh8Fsb5o635GBy25H8
7s9wFmzOiaCU5DddDG5Vxlp8vGZIZV/YiBfOlDvTm7Nf+4lCeOjAPjBwOW2UuCQO
QO2ZrWYVFkzIcWYklFJ0G58tGL0crz0wZ4cNhGrCU4IQ84Cwl/LySfYFzJWIFdhn
wLsDu5l2az43v0I5m6YaIrQYhtNWVR7PS2RySdEthF0Tnhd/3btLrSMbsh+E/O39
HD2xbA/Ak5c6cpFoVo312J6nz2FsV5aPnU9jdWVD+hUBfjZxTJY4MJJBhfCEQGSB
MrMf/nFntcW3j1e0PT5wqMx1O4ehXBoYt33Rzz6eWsb+WFpiamEYKPesLOsJAuNQ
eyibDp0OTBcHGBRyR3OiSsXg3rb45YAOf7v7MC0vYClrc4LoyTeX5SEgKQu33voN
SrL76GR6CCYukRDytGP95TzxYL+ZB84enAUIngbMs2aJK6OzjAOPdzoYGSfA0QdO
HKuUW2V0OZQsV4yqZxzcTwnaJrNmlVmw7GHnZ1CpJC3UxzdelVt4e7+C39eeaVKW
Pik6UP5R3TQf0OcamuLe15n3cvx7rqVRvcS+hUA9KICAlfNkaeGPklqktpaFgRcV
OKRDbS7VsmzUzuDetgupsfxtgkcsm7OUF92+h+B7k4yytPYet4zl+YQ8VokqY9/9
Hrs0eat1tTto3wgp03H1YyeCfviQMo4K8eLNT9sWsO5PrUT+L7N1iRYIHZzL73Q7
pHTPh6uVN45COdO26Khn3W5IoJ/7MmQMsHorvBpSJP2mrzSZ8AUE5hhGUxbx1Xu6
Ru059uKlmUyaORrB9Dz4KNMPX2JjzCEMmVrCG5+X1SCCIcM9f2MJRRtT+0j8CUPK
pmENoGvY0KZRNqqbWlQpg98SHA4g+eplBrod58UyDGtGXQ2SeFvE42ud3r3rc7Dr
6wpQjKZlsBFhQ44FpJ5/WKevxPF3ouVBSI4tdd5iGxLTWmD21Y9MGBEGtaZ1NUvB
OOj9ag8H5p5EX4/h10KmZryAFTqqzcOxTpWh8z1KjhJCN3ahbUuOk5VGGKwPUjnx
WUI3s6a4BgN4EQBlR/wyYr12zHNHXXE1rSKZgx1d+yEc6SFpNDhUZoj/DiNTQquB
Zr+FDUDKK2JdkZTPTlQCcbTz6IfV1uRf5XNzC6HjqrR+A20HuGe6T9+mk5QS0GM7
puz3+ubz42dpvzHKzXBW5D8peIt7gC58uZprsSLYChml/oVEs8CbrZcuC009jtQx
ZYrL0emdEWxzG0i2v5x9gG+AXLTMoLFN+KvhkGtNxrgRRjgia6ERbCG6ntd061MQ
uK9f2rlDOrVGIkitZI0LdC4oNCtbpIrZbqIocUAWsEfMZvPs2Fzig9Vi/pyaQLYl
9TPzTFrd0rwgecsiMqvzrCusfWQcClqHAA+A8MnmqYmIf/pt2kyllDZJOVZRo2De
DUD0I9BbgFPAM03JNrUI0MZ+WL1u3wsyELLlAWprqoAvbADDlYx51Ogfph879qmq
1rEAz1+VNRjlLtORsTtSJOWrRglNYe7tgXUnIOP7r60JX27Ad7Bk49C6VLgyCDQ6
fSanlHkSotz1gY5H/yP/vSlhpJSyV9GEN+lALbQ9XAs/s8oGjlJGv7wn72bXlTXk
lV/bAFIPShiz58v6KKGCcaXUt5ekO3mh2DyUanJsvXejPa/5xR6mYhE1Y8uDtzmo
Wk7e/j6FwqlTP54GfI2+HKdFSyKO0FlamUv5zxVegdE32jG1rk34dJkMZA6mluxi
xWa7xzlAlweJ+W8JqHUvh/ZPw4FCASJ1/PrQ9OOOYCfEP+2O+D8RQ1NbSOLVshrV
JjJarPISCUhm3h8oOqNUGcD1C1phiBqhbLbh5uvjDfIM1wraVwcT72S0fOA2Z2Ob
hu4WUBh3emLvJiToSmeL8KXgfQj0FUrq+V+uJFqrNunOYqfikxF4SOl+hC43cwsS
86QffOPS2AaraXgXP5dc3z3LZnSgAu5W8D/jnx4c+JZufg2HYuP3Y7BM3J5YdgsK
hg2lcHCJS4KbJB2/s8nydHjiiN60uYM7ovtf2gBZHRQF4R9GGXnbgLtrYQQVK3P3
aGSaWowNkmj7xFneTf23QQbSgwj7Phe0i80E2uDbdAx5vxBmIcMI35nEmPbyk4uq
/hzcK0KtXdw8Cg5tUSzNKCDJy2tg7bbN2tHYTwn2Rd2E/cKVoRwnDJs5NjWp20/m
FE05EUff2TRddllo7mX2OoKyUwP8SlRDA/cZjBdphXEeme8wNjQ9Pu+K3zqB4EPC
u/dVwD87REidjSZbUUvzenXGnM6ecHxGvL5ItVu011gMVvDMPtZTFpaM4h7BtGOL
rkyTwKAK43T7XSsNkjKczcmvE6Zi0ISk/YmvSHOB7xp3Nbb6k1vJaPKUxqUgsjYq
FuAiEz8B3gpToJZTma+8ec50aG9kXgKA3p/jVVbeIBLzREeZeFlKdmdwmntJDGce
y/gZvLi1UU+WbfU75OcN7wS/Fr5y/er4dO6CWQQDdNAmyC3CuT07yu4eeeTMzp4R
zxpNsYsRaT2eKRSzaAOTNv6+nqqrB6BQpr54/N78J2Gj6Kf+GAfIGaZXv8bzo5dl
KWraRK+X7ccb3j7jdLNEPAGGuxufRc6eyBaUGo5Pn9f27G9Qpaw9UlJSSMTvyS8m
lBV+K1ajvrKcCwVv9HTSVG53AvHvsQ5B1AqNfoV0jIXZLHD99HCEysxy2IbSxLlK
660AaLU3iMFuUPl8NowYqBy+Mpl8CtUDfjLrwPaV1lsdowQAMP7ZNJr9t2Brq8og
0t8XBlTOo1ljBPwKnSAmHM8uLbmdML3pzblGKz1XqIQsPhTRsyE3hdX2/5TlsjZf
fsC37n64rrBPDfwu+1s2TLhfThMsfCICd+fSXjN6FXXeAkzghDKX1VfD8EkxuqLH
xIWiHL6FXAN1DbJanMQer1vYULB8GkgNsqOcDdo0sZb+vlpDhG3XRqsp7zeibPOt
zX38HspDqktO98fkLDHG9IWGrPAByPJwFsyaRDhtUvHNGXUoQqpJjuTeEgpb5JhR
bdt4WkyKEmqLW6NFvEZR+QgpG7PHupTLYGbGLUA13qt8YeMARayZOgd5DxMntVum
o30+QiF7s0KOaROg18WWtkF6kDPe3BT2rEaD1q2o0yJSZDNBH4z5Ou76TviOaxiz
bdo22EptYS5wKNM8y+D9GOXQJNQXL+IfaUs3TL+zBu6N49czXz5mJAVxzJKuFqns
yA+g0N6Ha9rmlCw018Se3N2N+xpyHUE87DpQYICc7lEa2x3wByCbBtXx68JRCd5Q
bXiwrB1l1pKPVPRhxWgxuzmXI915GLedUeIRYk/a5G6c3AhRJvaGEYnQxbk2cN6M
LTeRWOn5xphoHK4Nzt9smjlJuM1z9xrC5f5n5fJ3GJCI7B+JlE2hZbunpDeGUZyh
jUuwIR+o22IB/64T6YiaDcejd0a3w8s9JBm/gqXtGTT3igtyye4jzRtZuXx0JSNu
M4w2xMfP7smgOOhJBzV9/NvmqQWr80djdewYu7KO5Qb6jmEh+hDlTWkfU9FgZcD5
US6Dxbqz5av2uAGZwD/8jlDOKYxpSlQpZOcHCnP0GzyFybMqT2g7PCQnGOB87N2X
WUae1r3hDmWo8xNFgMY0RuC9T049u1YuDuu0IzWwHaCY91GcnCMyioUHSGndPwm9
GlfDgdXOzX6go18/iCmJgWsYIdCX3jZeEFzXztEmL6hxIYz6rXhrJ7+5qKrY7Yj3
m2xI9S9/23LPdHu8Omc6uynNq3UtECCs160PddHKY5iGsKeg4cyXDPD0p1+68DHE
XGZmr/j/r7yL0UF3dS1XfzxTwcejghH/k4Q1kynbvfSXeeUXg3Gb+v6QtQTtaEDy
A+NJ7b8Ha0DFI2ubUp7U+fN44UdaDHETcC92mvxHDKuS9zd/qdtlRLytS+hi3zg6
zj7W7HsU7hAkjeiq3CzsyK3CWTic/JL+7wNKyhLtPNW8t26dIA9ySmtVlV3afzHL
2hvnrYpsmHmkr5bmjMYf/kYN0Wmt2kYC9yEC044eYfT8t17XAz4/y5HDwf0JcHbW
CWIAWg++dy7JaBxn7KMkJdda076PzUU/3Htagfh7v5sHKBVn9Jn75dwFhx1R6/5+
NGHG6TeUyugtic2HIrRJSe+X9U1qNMa7pWKKha84IzRARTUM3gEqJwdZWStRIJnn
K6TJQRCbppT7NXvyMOCnnSSfeyWZBO9eWf39MVh6GDC1kbhPYAOqiPf9bF2a10aa
IKSmc0XPhDVYfkcR6QzJUrASDDTyD6xr4U3kAU1WXOfAtl0XNueFcA4SmkpAJUhH
T+TcM7txJhqANreMb1h2/PcHfaKzgRfsmvpV8r8dkiw/3U073meCYd+ClIlMs3Hj
JSouEnmJNqw+r9Ucf9ktnQ4JFMdFNrWgQMWdXgwSaOPsU+N52qG5TKW7wnMuR52C
zVK9F7cZr/GMy1lOVZmGV7E7pzmv4WFl+lyIw6kppt32YWLwxlFY0pknE4Fd1W7D
RvhpWyUtR+i4i3SMhuw76jZPkHGmyJFu+JEjOaedSVw0edTSn4AD0WuFah94cpUQ
IcuWqaInBFczf+sIX1Bl/Y5S1KJOKnWHBjenI9cGkoQgOyGjY6aUILWlP6CQiQCi
EYdXtI++UgZADpvptTfTDfBO2qMz8EZPu5b7lCBBJRYsXj1msM+8u7qUrDjI3rMi
h1KrgpwC79Lrld8lj3NtHyB9ASdIhpLvRCqcLChLzBh43NGaNvMSBZEBnZQ6I95L
8tW3r86AR+KHVnmiOCnGlR8yrMpasVBt6sQfMD3iuCWFyDzsDGX6JNT3hoUyW/jO
C56VSfMQoNQhBAzGNUl6sWkTGbDZDoDqJK2FQQVPoeIE1DnJov96ll2VFHjSzh0I
sfw4UU1o02vWdGWAPG9Kydl7JhqdU4m2VIApKRoTa9H3WkM+LZ3icwdkmSrG3CEo
ZtRREVxVY9GS1Wpigj9gYm/IwxXcFVoi4M0DN6cA7Sj4l+Vykv+BP4GyCT3r2Irs
i5tetz3iH63sM7sqyf2pXicGEJvQz+v02PpOyMM8+nphUckDiry4fkbxnJf10AFN
PnUrocMmPAAJAgawiy6KxhuEc0tn5CtmbBKkb9YfJbIAewdDSu363NREeTxwFYHV
k4PJu9Bkm0317CJTw0VNkbfA2wyy09Jecg6XlqUaqkK05g0CUU9cZUrcVGdC+CIm
v3imGaDoLAgy5qsfnChlgkZ52TDS+WZ9ZrXd7bTZ4f6J32RLG9ef6sQUSRzCjfDN
UdJpdvjm9hhpCIVC30hl+HSorJFHXko9tNStys+THOBH0ddDu6scdxYAF3TkoEwF
yOUUpbWyNNfbfNwF3b5YmU+PGJg+dv+JQpw5IGl53yC7g8LSkgY6sk/aqX9nADte
0zFUxYgVQ5ac9zEfuevzpPoR3/ykiC5DUhEikADqH0czS/KInjxZ/CkSM2AuqWEs
VRgYxmlSxNk6pS/nG+CgHkUjnkhdZAd+IkGnLG2NxCj3SAgEcWBsEVjUmT7cz0r1
R2ZJPbxEiHgFOSXtMEnoc+IYlAOScGgsZONbXNd7NDT0JRrJzdYK/Q5lMJUp0K5Y
Id+BSF9KImkFu9V+B60+uKY+GQ51xk1quaH1z1BbQvO3ab8Nj8vfek5bLqX2r9VR
d5EmGlViZFmBkJzk7V+uwJBID+tPvR3CXnOq7GH+fE774LqMPUre1HOrtMDDlT6z
RSeE9G5JapM3VmWeDSz/wjOw00wDJtUwBJspxaSVWh8/LXtzUHSGQvdMzR+nJ1LF
NC5xX1Up1bBuEI4JZdu/6RusxSc8WraHMoYX7DzbDARX0bQ8GnucEZg5sxUnyCLk
2021peHd/TR/njy4cWMTeeo6yD1C/PUYJNZLEwzYkF4mhF+Rio92dpYbgG9+Qp02
1tXN5cnlJpd7VYPoaTT7h8wRD/uRBhT9wLooeL56o86WSMSuM87vDIs4J7G9U+4M
bA3ESbe/5x1nkGPer+ruwpBxtOgne20VWjqwHQSl4CTzdcKNIZ3WRObHvp6ht4md
xZSyjyIjk1GTkxNRX0DTNujHwhLit/6Rl4aDhDEt3gFMrc35xbldsRQNHeoRV/WV
nzhs74OO3GsgEp/4VMeFbII5M0Q6SZcarJL1ebJXndl4T0WHW/AhKiZWDSOsFz9T
o1XwismDanBYk0uL+m1XLePvGSfeYxLCm+wu2RJxVh1FCj6VFGwm/jS9KkFSIYZs
fT0GC20nL28Px3pZR2xe0RzfwBcfgj5eEidsqaj0W0zSnvQI1WvGQFmRATXZyKb8
PwWADR5fvWCe0mUZeLor8iczpUnX61Jlj7soToR2r+V4Xe9onlXmNK349BYUJFDm
lxjumkQ2L7IfkMGbE90P+72jFVngiqtxJTjPAQjp0bfYhX7I8wtV6v08UhVFvLBw
5odKJNhx4PchLKjU9270RK9KKpPf2S0bLD+5zprjljkgGOt0W1cSPicLlCcpIvbM
R5JOUQJvqHoW2REexuFqb4Zc74vy1YlY5i57ikdEmtv29BnRgSpEqkkfcpx2HrJI
8h3/fsWnHe92c0BRamxl7B8pXSbzvfGyHh8g3iyB6Sx8IrJiGpgDpkSCXqTggHfj
Dzj3/Yn2yA3//XJPOy6pEbl3FfS4Rb/qtEpxjvTCIMEpqSqOgzN8I4oIb8B0BDpB
9+cPU7XSEr764lR7lWcycUpsnhPt0WDI/pExJJMHzcAIeu4yu92vPrA3/K9afa1L
0VgZt1Pd7qYPS4FWwQa4gtcRCOGtHCESFKmXLPnyUiqsK8k4wiezC/uQEn8tyYUZ
xTl/VKnwFP5ur7igAPEMABdYoTRR/T0LyN+AaPdcyOa9CsHk8/oaaq3/emQ1osAg
lJflQakFfDsNwFnTj2lGnJwVWICl8b9H5+FcHz37exxAuAmFh2x6wPPECp/XQR6U
lAuGa6vOQe6t1Ao/VW0ICF8ThsM4A3gq8WfuDYsfF3QkKrBcMbS7YwNOy8VoUVH7
f8yxMLFNBMQlKdBGAB9mjK60mbCf31dtjAjA40mLFz1w8vvRNljTA4JZUpuFEJHM
z7fFk4pj1EE0zYotB03sV9Hhi0/avTPVHuVKU6gGLdtGyTu6cuAG+6ffU3GloVPJ
R30gGW5+vHkYix6bj7Yjg2MZT4U+MhW9LeCRWueaSIMA8/8YYBWti9+dcTjv4gZW
KzHa8Vrhm1g9oWWgvke4JASneCU7N6geyNscL93/bHqk4XRd25TLhzDyatNeIh0P
xC1SIxdYkAAfHPDcISYZPWRWvpNLH8TXFqZEM9V9uICg/VZETr4LO17rI4KaNrAl
T5o3OL6S7178+r3mDhOE+U2QoVopSUAbgw8c3KMsA8bCcWM0Tt9w3mrUAbwaW6OK
p6kIjyGQUcFcNxikoOKzpSIz66gCpuI8I5fTMChjyi7xiN+Jt71aKNW/rtXzSHKU
dPWRIfkmxZ8iE07S244P1k9w43ivYtrVWO1XqSzHoQjKJmwskl+ygXgkdp1VWl8x
wKYcKRGHc008cfA/5t5KaZgT7/s0V0ZsbXeUyVtJKTWZXAus5OB++1ylKxySYrv9
NP5ndVXaxaVgc/P7WF9ho/s7Q4L5yzo5MVW54tGhsdfbcDCiqk70dPRuH4M2/y0k
axoDEQzhfYIajr0Fxk90+L3c4cERBuYOBmpdgCgXm6QheUMYEoNvfAPrPB1fVPQV
JFCYYf/kSY4Glty+8MKbDhviu38mZbdxDZOt8Iw4mVEfGY7LSQMdZASMW1RCd1nl
yMDZX0j29+VQwu82nPY7s4Is1oJkOKN2vXVYnF3ZQ1XPrfV1MZz7T136UWJ9qf3E
ayed0y/WmftS88kkeCDhF3JVvL2/Rjl3yuy5OZXpJG/TwdE4QVd0YOJZ8anQSUJp
+h5RlnD6pqCK6b1Z01lbzynp5JyMmHJgYm6THRCxGMO9nQBsCG/rfGn4n+Q8fLrU
4qut15iANqoFhvbep7p2LeVlUtrlhi/Aom1gQp5ttZ4FqigDiOxQomtWuE6W3Ndt
d1tTaWCmFMtIpiGMmRLV3N0hFOo/L3ILkXghGeSAd6hDDUf36jU/sJnj6sdlndmE
Ko19WU1S1NywRzUPw3Ok+CYs5bjv/HU3lAM9alRwWohGW4wJtTfiSK1posSzT5sK
WlHweqRFWBuNQfmmkifmqauV5CuM+z8KQWQ3SaCB0/FHOD4pi3HcLo4lpEvQYiew
ayfSBRfb8UpaeV8E0Bnc+dPhsPpwXz5n2wk/ES0pxT73N68t11LhV8G6MENpuYob
M/Z6a76uwfsb024cIGf5GUwEfeTJRtyBmL+I2AwexppiSK2SV2+LOKd05LGqf8IJ
RQeR+/Ngag/FrAbSA22gTIxDRl1YsNqxmhBZQ+SALOIq9zD7D20JLovV7mMX/C8O
Yd/ZpTmCRb2L5ARzGvk3HoAZhmjsEUY0ims1AhdQl62FdJNK5XM+CY1HunU9TpGq
sp6T1AWAY+r9tfi3AXU571rX4vM6mRlGYPag3xGkF0ECOetE543GW1BMbaZm/vFG
OtRApGljXAgU39O8iq+T4XciBzfeJuhuxWC3k96mr4YjkCVjSKhvX0YDiDwEaSR1
1E381m6/VQrM58atW7ibSuEM6pLqJS+VSFy1hPJw3IHjkSSMSeijZ/ZU5Df18oVd
iTefvI/4FlNg889OoDH/rfWWgiYJsoIfwn6dktE24VTlofD9m2taJWU0/vnNLUc5
v4Htt5zN7sOp6CECvZTjQsEM/8fVeQywCCBZ/N+Ja4uAWNNmsZJHFP9WtZ5K/1DO
dbOwL4DYne+NvUndvNH5GX1WdufXYnIVNn4iqIYthH+EHbuvShowOiY2/aiZTKiy
lZ/XM5QMPhXte7E9k1sjZewixu9b6K0X1jb8W1aa1uo67vRKZt5qxYjk4txokUJI
5x9+pd/SuX5GwpaXJGV+xwWJyatt2Km1GDrLgOhFzbcRemYTTx7RVwzj7FWxcgbm
tgVXk384fsCFghM8w/cWbhgZc3cCZG/lw42w+AwBjw7DZMbSBt33wjs6n8HveV4P
ybucrhRVPpdgInJqW7sN12dFux+TfgvbuYVa+aL2GZm1Py9Kp5CSX76+G3R3e29r
XzX2n718DQj/eGyNGyjrXcF/bAcBBGFY4Ar19BVxnH/ot1sQKBs6LOJGq4P64ruq
TQdg/tnYlQ8XDKW1tYy12gJU6HZogWMoOmneS/06I/UgAbWSn6r4BO/ULXUl1x0r
tVpHUNM6aL3SVxQOxaE7ja//NV8KnvQU8J8QKTkXFbB6llrrC0shwCYkbmcLRiHC
HPuOOjoLxWsQ08qeRG+FsN+uetSvnhmCXYqbHa75Zm+ykQBIo8prjNXArfIDmKbR
bQD8erzJybJT9Dh0J0NTGFEwyxG4beoof0dwSPdL2LOTcVmdpnMny2Hlc0qxHA35
w+oGSH+Cw2B3p4sJCFE4jwDXY8FS5qyWIE440bMhaDpMi1YRqYSeFbIsjzzQPCaN
PqbgFAPhCKvXj/OFiRPGU7e3PsPEN6nqmrATe2QN3nfeviwnls80R7Ofy9FrMlKb
hxERxev9+vNL9F2lDPNQ/IKCOwL8jnWMkVHYH5JyopRs+EtRHGZdykrRBSecvocH
twgq9gCEVQI6fHzvyWC//j+rdQWKuo0hxR3EsL5W/paaIVJ6g+eYMU2qqondhmuh
+WTYvQUaPrzEYgwAeoPM9b+rmBJX/TDRa1gJga9yV3PK5AUbXE3Vhd4gI+R/nlVG
yaLwQZ1p0VPDvjz1fUGtGmleZxLPRabNb//tg+9cKqasLGi/w4EdsmyUKc9hLeNc
09uYbwvjCn0q28BvSVUzYH0WE6Nbd4wCAlcsvaVi313HJXek+VT3pbu38OS/7sTq
DSWvOGbIlSwqfFcUiUY5xatnJfwVX0UPx5R8IyjNeBtvREjbtguZ/wrJJMJvi3t7
DhLeMQJY/BwHetUwL1uafuPZu21V0Zd59Lxvg4Dy89b4kwUP3KK9euhVW5Rj+aeE
tLGosYg+zv30+jnG68RVnM7RmGcoEVWf+wNwqDujRRm/W2xEmOlZnD87BFCUP2Uz
rsxY/7gGlk4YeDOjlZjLUUqDUpTCeHVtTzsQScEKA7RcdGXc4JtE4+u+KEd74B/r
Vdm7Q03dpdCoqJjDnmCyiQvyYDWoxf/kryjzegsSfnX7QfRCjxru/oGffTwuLjxv
V8g3J4HDXl8x33fY5A4k2cixGtKjh+XtbxTmUS2DTiUaDUgAEzAqF+l1AFbBJscs
4fseS4Y2aRdOe5ULPMrSpsQIpI8BEwu1y61M6IPemMER75umKA1jxpWVPLaqvtu0
HWf2aX6sbfIbwMY/9MDEYWktuSKtbTwLM9OI6V8jFA8Bm/m38FxHZVq4v9iriQZv
VuOOcVLiCPgKyEPVhYgr73FzKrqmeml9z+tf96oeRCNda4zyOn5/mtWGGqV8vnpa
uIcob00+qfXVEU5o5qQwJuZbIOh/jpN/UyeM3+VIxAdOgK2IQs+zPy/Tt8wXaHcf
yN6IHbscwkp16suuCkDBO1jrMJC4iwIM2HPWPhyyfO5fIJZ6qb8s1ZrtDN4xUiBd
InTqG/et62l4Lzb5welAqEN5w8pwRUR3bxSy3rK/KSKAg6T0sKyJ3Ij9DQb7QZt2
xq3K3s2xgNA+oIxCVZNj1bc8Ie5JWI3Vbv2Ex35Xj8EmfWNxVuBcQFELTKXo/0wH
VXXdjpDzx48SLXUkoL6iuM7HujAIK+vdy/q4np+HDfOckyTtlF6ILkk7QzaQlN6G
D/ufXZ/nEwpS5QaefpUQn9H442Mu46vfdfhHBSVCGPvIHSfnA/X9t+SsXEbvocnW
jpZ3XbDwiwlKNfsFo2C8+FoDvudSfTqNXGKH1jbhXBXNTeZhspUBZYoGr1R0HrN5
34AXN9IfzkUstMGglEbBPdyPbK5GIME6byvovu4+MRPYv343nQZFs45FUjxXOZjZ
b7rSaFUifLGKB2QirAEVi2AJPSlts6FMlAtkP++iHV8zyqgLWwy7Z2ugbTw6d34U
Ukh1ONsxxGGHig6igL76DorA/kdi5dgWtvffvS8B0D+fF1Kzg6fKP5T8VoxQV+/0
Gkou/Ipos2ekT9AuMaASAA/iLvmoo9wP2R+VD+I8hBjg16w6usBBuvTs/oADVuxe
lUMoSDKSDLxuBgJyns5TQc0gGAvZTYE3m0cla8UR6LEbO6w+TcavFS+jHqu3mIge
jsIVEFFSX4MvwNM477EexkjykYz0lrKfOpLbw/nuGGIa4UlautuL3e8GHjEfE2dJ
nAPWjnWXY3tE3B4Mp8UUEVt0gG2K3tNNLbuQUjVfYVgtSN4TGliMv01nv8zBq1U/
yExnfN+rvfrl/gGu5Aq60PtHZpPHhiHR/gQnWLKrEY9RqL7JVNOqvKQJ29Tiy2Tt
4KHWh4uB34wW+UjGEGZ9Gi1ZItgK3Gs+Yp1t0lP/g3jxKgvtG4V/HdnkrR2lqsEc
MdQIhN3sNPlEtYALybMYHOCg3xYFCxZ1w15vW4+8XTQWDwkkC+58bmUzR3uvEWnA
4JVTcDNvrDmz09mp9A/rNv822ZlMAFavOkFFtCZvjMqKXdyOx+Z4BbsDtNUp7v5Q
Yc/vQffxDj4XDXA8k9xi5uDw4y0jEmz3gVzXgORgMxyBJLOHMUJVrbBOVvxV9MqK
SzwgDNSn2uFO4r0LJFDc8Y4soZRTY+mc7P7K7azfZtww8P2TaoXucIRgbjcI/6XB
iCH/Lf5Wt73S7bzC4LVf/qL7Ih3jp9NXD4s7leIuaPoU48RwieF83WUXPburzHgP
rPAkpP6WKioCw869RYWMcQWfvgnn6maeiRexUx6Mo0b43nD8EtDHDoJsZpk0cvjZ
grGT6+A+sD2ThljnEg7CKPbi15oHdnm0obNDvdBqRRHyponYYTh/SX5fQ4ZV/FUd
mHwluIfFpRCmqd2/bJsnKIfo0a5kxCbvdaiWATxBR5TAPI4TlxOPjyWiCBtV3gie
OfQDfB9hoWJnpWHjJ+Um1z6n0JmfSaQH4M/Un7tJM7PKBex4tzKUmE14wPDCjIRB
9Q9+sYPQepzewGAM0L5OTtshuR/ZsHjKksE7j31tsr6LEDcxCIFm8R6lFzS4TLUv
JZqQZjJ7V8yrI4z1E2DV8IuJ9i+efJr4+ys77qUyQUgcagS2PSRrnEdMHDpKjPkB
I1FNwMoTGIvmRrHBkY1x+zGahub/iQOcixk5hnW0hMFFLscNM0X84+NPKc1O+eKH
HiaBcr7yidYBSxzLlkj+e/47Ijl5syIvIzhc4qDBOCW2gAXffvIRaWkrN82a8Xy0
17InJg3ISmAxLMYZvZXPcnqm2cZH6s2JMnfmdoRk47hZs7FxTy5vi0vzf2FHDfZs
Ehu7Dv8Vf4+kpGF3wZrn+CpbnnOAOi/9zy54/JN26uGWAXlQEb5EYxZQ7jr0jcrQ
EVFh5ylR9GumzGsV86tZM7HDcxtjio7/9zK6WJCJ2D4Cj+MRh1z7E2MP0yK1F8Xe
oWMppeawbNqNXLjttM9ijteS89aHVNcQ7vm7hrd+jbCMehMKH/cpyU0HvbKXE71l
GqvAazGcAwFKyRUb4w33dTzb5ovXkI2afXDgqeTnv2SSN78gd8L3WP1S+wI0dZ3S
rC3B+bliGI4bkv+2zDetDdVH8VlRD2BvJ7f4aZ8LoLoPpXYeheTbWhu/12PIW+jd
KbcxUV3Wk6xWGyqB1dylFn3Vt61/Y68jMDfNuqjAShqP6uUY9xfjMksBVsHNFxtd
3UQq0oARuc81LRjwIHnNfkJbpF2yvdpd0nliZ9tntidCNbiuk7rQmBcjMMoS5BUv
oYG63vMvydQEd2I4HejwwBplPqhEhvDgo2ZDyfLEozxs3sX+ZSa243IswLfZ5X9k
ztZVmFZZIVkwd6wAjqXRLrquTXugM78OsyPEP/IzffYkQN/fv5bbhIyRjgPOPT7Q
ITByVG+Tqi/L7opiX9ejnEEWTzPyZ01asdYC1/3HD372cZp5ko3LlS3l78KMn98x
pSkfMmPYfZ9SAJIHxFHxVaClQEIWOF73rh0WdoyE2RwwIZOqUN+0hi84W+sL3HBh
DO5tkboQh/Hi7aRj0C9BWWWX1totHoTpgQ1NBIFdWwroEjP0okmj4AMQcIkMlxtV
k2q487pGpbp9b+CTbcx/t+TkTauT+HWk4hPFPPE7669ReJMHNU0hgNbRfxtxKpBl
Uf9SWEn29A2RrEuCJuapVexzKxiAtPtZUbZZNHOGf8ACRFvln6z0yRjSRmtaydMm
nATczCO9DWJ8GYXTFIdXuJC+ZKR/Hvxw3tPs1ypIugdkhZn5Wb8UUzTMTVZEJ9Gf
MfTdOcJUh7UnNnsEf2h5DVlntv3kpNoZ0ss0/QGpSJWIWMyGa4RvcBhSFwaVOeqy
kMVhGK0OePpGVYkZ601oXpLHIEFO45oIefibh+kO6nOlZnUf39/jLIVOEblrlsoi
n9QUnub0GpgUrSSKTD+Dat7ThGSG9jiTKeBfxxryq93Ds2501aYj2JLexo9lGUx6
NwORvQpsVqiWQTvXTerjvzMgCHb2Qowiemtz76/rohrlECkYxGMai6OqzTb4Ko/E
UOzsoDB/cnPSoco1ESlBsP73Gk61XiiOV780QKy0RrosL7hIKBouo1VDqLxITvib
D34E5RY0e3lcY9KPjnOuZiUdEwhDk9OBMXEZoKtgKaTYq3tPdIBgvlvBTnlfIgs9
sTIRwxUpFOOhHpSFM0YcrqsGacwzxpaGCizn2e4BOTYo2BFu1NNYBCm7xKm9Jp6I
nn28ah2ROS+Fzk1hlYIgmQTmjUzvDMJu+v4ox4Twk1214T1x1XOk8VMzxGGXT9tp
qzrySrbFfqTQzuYNclLsvJjhlGRNrJhJ0Z/x2dLl+pXRIOxOrWX0lpGgovHLcirh
zTtYDdUsDbWTpd4PQuv3rZWKePSlNQk/IbdibYb34dYCQGkmA8VkmZFRxN+NZtlN
aNBgIPS7ic6OPMOP0CtDCy++RyVT1tSWjsY0TVF1rYhx8xF9PVtKiVpbTLBVLVXD
M5D19SjMqNpSMLhc2QU6r+gxRW/aPsqvDnPjZOaC5vg7Rup8Z9gENi0pqEsBtdKg
6lKS7QMRswSIBCeb6IejnFwl6lyw82BpEhtBcRqREiG5Auvu+ID9xktBE7R4gIb6
XgacYnAcEyyMISzIJjBMA3lhoyRxUTdydWkIIR0xveiMhBWEPSnlFQUUiHe+ad1a
xHvw2wCrh5E+wRCRNAvmr9ZtG+VT6XrXOZa6276OfEQdcThu2QFdDuDUjlLQXKJH
RGbEWeaICLCGfxlp/X9NZvW2XBS+kyf6wl5LqPWM32MULdvPZjNRDVOSiKuIpaVY
cAxi+RKY2Mz5o+KYi/GhfOkrBD18LlRYh4ltwcJbTNpfaWyREFtOJ4lRQWNBIdmh
9qPCFvZ/2Ak6jxqTz+FzXQmLFuajVp6wKFOam+2MIg7UCIj5YMOE2iGeF5BJbN8Z
HWsU3EjV5EQwG6ZyG/V4HqkJWLD9PNgvQ8fk9Xqp2DaRxsBgmjo5sCu4Y2z7Vw/6
PAnvdXuEMR83s3vjVW4W4YhOTHlRaKvYqHFbm+DJbiALVm1AXmlFxqPKDp2AnRX+
n/ayjcVY4u7tZjAOcO1tDmxFqk2bSkDBGQ584HS7ZqZ7oEutt4O16wCSweOAGR57
ezhnyfSCkcEshUp0cg1OJ5nOY8RwX2vqZnK4THiLkyFX1u5zW+1a84QOIF02fLWN
FbswSG5BxFihRns4j8G6vCLX8dOGA8ndqlx2FiFOXYn5/eVB9bNlrLWBqbPClm2W
tw31qIIi0FGfCAJ5bYJ9C5oqxxbhSdVYNsvgBsIVbYmPtJioeMJwE7/noD32ATXT
4KbNaM2nEdbmPd5Mu3TxOl5lWgtNMUVGnXjQ9CNE7lv+0C94Cn5F0jxa2zz0abXJ
dtK/P2pwa3cjd02rrN13dx31KmQ8FHkd/YPrhmfpwN4NGYirXL9TC9OioMDhTJ3k
/OcYa4cULhWQ9iL+yiYFKu3Rlec/yJLyn3MnU06cj0y9fUpA7FMnP5QU2v5tIqCL
8b8rEdzDjNPkc1WMtt4O8xYQjdjiPI7D/m7RTmusqnyQq8/z2bDyz2nBbHb4CwAj
ZyvKN2nMqE9g+QGUj5JDBC7A5zX0dQG3M3SecWK1s80m6Q/6Ey9oBezFM0tDPgyU
Q/zw/VBxkWIpDW3FrTnYTmraeKEQNH421dHTuu3Fil4jhTD9JxJKnJ41Pqa7hmiz
rwTX5WMMPqPG+wC+ynqz2oU1pNHk2ZlNH5HO3O+XcxZ9KfI9o/HD5RgmPK6uWSeo
7tTt8BuyCVwbEpRvxoRMdZcZSI3CBDGbvC7m2o9MBVT+aUKqM0/LfJ6Izm9z64sF
r1Rehi7miv3rMSSl7HFo2pFYvjWFrHAC7Ycmd62ngaa2JfSyIG75YeofEJ43oE9f
4L0qkmZPErb4pNGoiJBZDgwVZ4GDwE9RILJ9wQMFy/gkpe093yCH9jsAs9P3jkZG
ADeKRSeacNBB80rRVpRonZHopAyyRH53qE0NiYBDVuDLckwwr5t3qswjdmE5bqhQ
QEyDv1fA0iGqgfoFHqxRuwBL1X9THP9v3sN1mlgX7QefIRzOrsLv+tAOw8EHwTD+
e0ij51KzyLhJrHDMed6kxHEdKQb7GgdGxugWu677G7FDsPNhLXW2NhXAkbe4QJZB
D6lkaNRxypPzrdwFFB1IJIKKAZBSPHmn2Q3iRZZAFCVdEaU7WovT6yk0qTeRiTiX
/tkJcQUzB5bnGDnirYL71dMpxGJnvEY3PV/yeqDr9b9L9htbT8hvdSQ93h2n0rsY
H3d1W0iGjFO+ZFkM5u1Dt2iUIWqD6gGiuHnm36mZTV9uyv3KkE3j89L4Zr1FTUAJ
uu9RFdVW3APcceKiCszt73CpHTGFqDD6XU3Loi2UOeE6Ge2r/u/Jyg0EwLRM1V2O
w+jYwr2FVTps/rs06uyEir3bjN5QZxVITB1udFOujAzLi7xiweFcplh8Tg7iVDGN
m4xJnP4wBz8mtws4nEPaCnu2wHj9oH/OMQGCvrrEpoi7V8DrvpJxLFE8FAskEypQ
QJmMgkXgWRHRmEkSrpbY9zoXbhu9s71+BN6cTAvrNZ8VioyEnMcgWHxFBAbNpUTV
pn6RkPA4lAvgtuLGYSDeTdy+QLc4vF6y2NbJBUkwF9JTAUs07MGFBB4g8LNhG6FK
92kDl0vm0qKFmcCdz2DDxGS7x4qzOjWbdu1ZxgUCe5kSGcpy8FM7vEeDsgfMLiHm
g48w1FLSh57My2LaglXtSqkRy/+40acrU3dsRb0HnOfoBZakVoxX9fMZrv8MT8Gx
2A59JejYEjJ99ZYwT62KPnDhb6c9o5By/PxLuSnkX2N8FTTAFEXbUvKvlpLJftLH
X2p18O3gmDuASAt/y6/TZfkLxHHPVoNRUodV5aIF+LM5UJuGvMYvF7SA0mlSCfv3
mRGrveXRb/aRkGQWgDq8UeV9DnZnZZyHZqHfkXqPfsJcdbpcM74ca57x6WrZSiQf
aB+bgD5jiQCObuuQB9ZPU92uNb6cSJBjfyhMUgDcnC+TV6xluYIzXWq609o4uHHp
WcbRpQQ5PK4br7d9tMSXOfDkSYdo52wdaUxOOlI94rFGtmPZBgAUBgxIUWut8yud
qY+hDBMsNEA8lu5pmP5Nn/IZ+yGZaQTpawI7i3BWIES21s7ZBZUFm3J8jUr1IVK8
xpf4kW74kS9z4wc26Ys79nzNjmEAtl1SA49yilB+1wGcnP6qlXhpWLrsosJlk5d9
c/mR7q+gOl8yOfnOWhGcaZvXDyET0fppV12QIcPwHZf+tByb/MJnOVisOQUOGRzK
+hE7AqJ6GcKPwMp6XViluQ7NJ3jZcEpoXVyAEc9uQTlIhkY4NxNMba8GyiJZK7rI
JWnBwFHjjbbrNbRZFvd83xdMGOJEucxcjL2GOTBMcrKJZ/0+UWKZXrhpRg+51tLw
lirqm9doqZ4JrUVWT8NksLeNQTvqxf5ZZWnOtHhxNxhcOAIguWIOj0BOdECjM1WR
si9wfVZqtaHFqq/0gLZDRbjwEk4n+ziWgtXn1U9E14nIdxwePD2HlUes6dPDtoCF
Sgm6/GJ9P2Hit4R98rMaWWdlVWtpwqYuVyGNM7JH3ccjuGosRObeBmkoNatin4pm
LMxsbQgyXhZK616/crGrtpbDoJmp8fwTNtUw6zGjBZRykyHf+12QooIxr8hQBDlK
cPib00DbVCW9LqF0UobMpXwCt/sQo7y0kP3fQgm1qRNyghppKz6e25y8ZGOIex9J
3eb3hZTfpf+6aFwBKZ6tDghGaF2szzoX5pXFvIuyaQt7uFvXZYwFk+EnmMqj8FGE
T2Wf7nPsIy8O7DRIujljTE02Nk0+M4tJ5uQHI4VxbibwSTocqF0hvXILlqF+8w+p
W6Hj/M4jQPuEmCvpkDcJ4HQDPQuiZrqB08k6Q38UZpaGYy0lb46lc8L7bJu7GwZL
WGa/HpLMmYRKKMFPOoSFZGm0RyFOsg/tAK2/TDXI6b87NhnUTdVQQVxA2fhUPWIN
kM2TeCQMqWbnz7Nh/2HKbKBcrr0h32s8dURvuZVB48c0Yj1keAbLumweW4jDAuXW
KQc97uOKhVPUUHHan7kJlOmPtmeNybglRIkmu47ZbZi05Lv47k8dGqSM37LhKoOy
XdScXqwHmBlyRt4FKu048xmihR9SZhC1f+l6MEQQlaHeNvRdCPNxH44PqhHvMkdu
MOaxGaZij/DpAJ48KqjR3XJjSQuBo98RoVjC48XOF9QJkxx8AbsaxdQQWJrPp79H
NwPXDadS0hIL2PDuVy61QMNsVj12uZEWFUrPjKk5axUgJhLGoN7JklOk/vxOCitv
ydynT9fphbIDxWv+7Sc7aRGa4FN74Q9o6ThuIFtAr65AGbhofvBzROchmLjv5Gew
rxYyPZaSnisKnUqOuLUM30wwZ3GFIeG1vAgEQ2mmse8hjy5GTf7Sc3vaU94TrOjo
poOX5HUxCWvPTn6/qbsi9/+Jm0S0cs9X4wl8lU+E5tAm9vzc2IAWuZFaEJujk1ua
Y6c1kUClj/OnJzcYOjfXqx4evt6m/Mxl66Pomu7EOzHt5/h75elj3jEKg1Hl/+DQ
GPI+NsCvf9S6uZ7pguL3SB8e74f62lSLMq0bN3QuWhpypw2PcVfNFw+0qcYgmF6h
ZaP+Khq9ePp1ikEbtjzkyLoxcCuNokrUIiZGV8cJ2qiuBqUC1jFQrRkgVoTYk5as
Mk4VqWvI+aJancnVd4VBL80VC1NAJYXU3bLu0/3qwXKUSx2wmw6r2ba12GNsdOwZ
S1zkEV1y7+hgHoL5kWUWO76M8XLjqj6qwvRtXKb4aXMJ4f3Y3ysTcJJfWOlbqfGc
MQpqSSTyMbfUMX13qlNYgChRLjI84AXVdIUZq0YXesEYN+WCiyIu9IaKqtmM8Ybx
y6WrYDeFOxUBFHCq40jPXGlq2WW2d1F3DylhAMaFiiYWOlTWbKbNGO5Xls2sC83I
u71ohd0xLg3WSc2A8AcnsavNSXZfHQk0QdRdUZTpvFdLRhZAFWiUJk4kNH8105cy
94nvs8o/YepscwRksd9m53DDLFqDueeNjnmbssDwJOO4R4SJyA6I0CkVe7Umxf6W
XRFP4fVwT+Zw3ObABOGm1MKhboPFYTosqONi/Eqtq0ksXzNsCmkVwS4d6+0DPX09
pnm8nOnafLS7KX7Jk6fGWRY+MeyccUFRq+Ft7QwrDjXRLVz+DJjGdw42dekEJGOp
cwlVimRck94WqdyPjbC79rfj8jgsWkhVd4SW2VrQouQa6e71sp0KeTIWKJQLFgnh
9/ZLDfdm3a1lIKH6JyOK22US6J6+WyDDk+kV1m7SEIwH5eJ/TJX8l32Pnw4H+jia
9/XqRsB59LVpa/VsV1gZWekfAlQ+rSzM+RdvcRXmG+8Y5qg/+3rNky3LaEFbYCMa
V9/uy1TRiZH/RgMD9UdKl4kiCJ6PRtZHdL0pPUUZ7Dtgc9yGCmp0NQ5+KfJC31cL
YCXFumzgLiR7wjzvA0VGQFNSxyJGOvChDhMMwUWkwbAK6cofKLisu30Pp6VFuSpY
rTgP9ru/CLkjnw99nxiU+z/xyfDs9/HehCLtipPTrviGdW3TK2IuUXpz9XlJAakx
36bEJkrl8XevTzoAsCQG1LpvtQRn3AAjBPhmirZdIE7lQfcT6gXjJ7e6/gEEzT/x
vTDgMPEfrfwvdIau3oiGKcaU4MC4Gh4lFkIolw2uUxv5dYbFnX0w115lr92jajvQ
f5wIQuxxffcDSEGEwDLJk2qchrtYgrILc2IYU18chun3vRpXoqzsqPHy2VRntN95
ZwLvsufwGJji/RDGLVpCLuC4Io9DNFotYLw/LDdSIvL4jE8PpEIbEpIZHm1F0yDc
6KccDTJTHpU5+/OTk3aMLLQ4z4r7jNpMbXOush5eOlddmudztNchG0tKbEdSuSlL
u7EZ3U4pF/hwKG9qEWkVQSnJMllN3CT6Z2m8HP5nTo/lj2qMS3fgXshscEXkweX5
MA8avJlgnooP1zEHBEpXj7zheIXlej2Eq8hQS0oVsL0nM4Ohu4WEFz+MnfyP5fBv
RHaf5JsLLkEpITkIzaoGF2YgtXjOJWsyXyxFyI1q9/YYhbD58sWbFMLYqqb5J41o
RuQzYdJwn5toy/sxG/rCfFsfsAV8ld5ZOnB7e9uZa4eIviqVU9rwFfx/r/PtYQU1
8rHXkqOfTpmQf85JXf6QG5okQrfi5LQtx0cYdAWLiUTHRTBOWpiYTmDEeuM21dtE
QOZvPCzKWn//JPjzUstx0tPQkz3UTjrflwRyU5In73WFYOu0x0edtzB7eQpJ3Yh6
AbHfgELydNYIgRpTUjwH4GKe66+KkfKjWHfOPZ1uAcXOCdTb/F3zVYIdGF5kzrZS
dselNhZNvSUNnWu/HuPx6OUq/yM5cG+ABwLY3Xv9U9qtOZ0gkYI+LKIYyj3DHiDe
V0fgAfiYEViVPZ3kCNRNZlUZU8Nd/P/tFUIH1SMzpPEavIWajkCoIev4k93rnUv5
KMWjav9k8+ItHF+zu8SOAUqpnbCxzbUYQhA9yM7EJpF8DpuNoogDdOt4261b7U7u
TH49U5MVzhny8kSg930rQGLABDWMALXrQ0COsede4uRfbP11lwu7ImBUxgx/Qfc3
AsknWWjW+LEmFKlLZQxS7qXUNme8P0f/QrOwWkOsjJ9D+NKNBqcAKDXtk1lgtOzJ
VLLCej0dYpj5Kwi69YstJGtGhxUNbDDCo4HptayBLQh/LHsisB0/L1o5TzTNuKC3
MnqWGwnygchVwwOf0Kr9PyBsuL4uvL9JssGs8yTJV3hD1Rpps/P2UG9Kk+7TZHc4
dh+LdpgxJK0/RI7ux02Zu6n7gMuWIiSmOJk/AEFT8C9Ju2K4c8dX1sUb3tkuwoND
MShFOIVHITkoQetxRbGlAy+qiEgME1QVlK9uLwyJIqfG2Ah3Yqx6KpXMLMrWjJYp
5lej3O9O+FvogmZ6uROuhS4uutc+ekRZ8u5uBYgDxLcex2oHY94YWe2wuI2+LNkc
m1V3v645ibCjODwdtrweQxuPYWOYFQOaOYg2UPwb6E2xpz4IOj6sJrB0GVEKjld1
qwdN8/S+aL/n+GmaV63CSY4xboJRDtjeAFgq3K72Dg/ZTf/lpfGZB5h2u5jKUiAh
lkJPGNGyEDd2gegdPria6pAM9gIL4qlZpNsgcg5kr1iLjiVHsBlw+tTzIUo65Vw/
E7RRxOv0EOY/IcOhF7SZ0qzacVUmI8E/OqpGS8vChUsvmJJ72og19S4dIC6jcDzl
AvUZGLxNj5pTWaLPci2gdcvbtpQh2BtLOjQVQfnnWL4VBO8KH/Zf9WEJR2G0Ra29
O4G1MXU2qtLlIPE1TXT1serqFXMl/mDFIfw7bTI38WsrCPRDnWFl1N/JsMIw13rI
IVfyldC00msX1+V8vNcJgd3590ABPArkKO9CtP1SXcnrt1EX91BugpX9AGeGd9/X
bsDZb7SfKtaojcI1AstOs7qnYKyKRe4Fx1MggnWXoyHT9Y6FW50SyZlhiwUOAFTR
tNAoVXuo+s4qAPwhzCwpsnQzAiB1y4jJc/l7lye2+R3ahVefZfCIucHGdKwwQ25H
XzfN8SCACx/kiPqt2FjsXvCM00XDeP3BIZxSTNHf0XW4Bl6KOzpWOoStbnDUN69y
bO1Mecs2fiPYRtXpfYRBby51IOY6xSv/PkcraFG0Y8vqqXquxf0ZnYnnG6nqniqy
1EJBeGEWxvtv0ysTYrg9Cm0vx1QLUXnA6l/tvFRN9oi4E5V+WW85jGM/1PUJJKnA
2Bh7XoLlfGmfr3AWL70jkbV5BV8PBeZsDVsDwEtSAz6jRYPad6lQGPJPMjz/p8Tk
JeKKLc4zN4hcJj9XDWb5byDNywqnA9xCSwIMgn3SwXZD8uoVvg9ou53PrQHpmXJG
WiGQnILFlLhI6zGRWGYuPdanRv719+CvGg84dmmL1cKko2g+2a2F418yjXiLSnGy
yHZtfMBzJIVBSGCASKdGQotinMeUf1Ui/K+0sQYOsgPzXv4TAOqHTW5RWeSJOcfT
/B/WdPaiO5VKcjvfqinbkA3tRLa0fSWMvZX6ch0WFGB+ZDmILmuanwPxevDMTXWr
2B4Ziz/EWet/E7DcKeKnGiPG9bg9mGs0AOTNNiUAf9jI0/+j4TJ0A4PUF37S1MSK
jU1H/oG0C6V1RosVcBOvrCUcpOYuvZJwHXlPoGveolBVQf1X9W00ZntdoHGk+yKZ
SoTHNI6Rswc1JUn3q2zf3F/nRnUar1S+2J3Z3P4wuyARc0xMGFM11gK9ib5OkwkF
RM/NFMM+XvD85+ta8jkOFEtLhB8lzcctNKpdKDsPADmoxU2OAp3Fsj9oN8VD6iux
NZcwZi8s5m+rYtQnQkFtm8hiDpybeTtcwXYz34dqgieNFtzYiwF500p011sk2tII
nrXvHoGcQkGMQLzToUHW3j8HDzbXuP2muNoMIXrDon96rTZHlH2kTXO/RbZzPuep
XRGnOBuKdKNxsj56BqsBVfzNwHGhwaut7AqO157KRJLeyS1J94IQTk9H3V4cSuIe
bpy33ERKSZWR1dnmzRhzD7a4x1Ex48zG5yIOdLjouoyPY9WHl6jXhtfhGqsR4K9z
peJ/rW+1gGqo1PCqQ1vWkPE9FHeKqdLISW+8/0u3FaSOuYbl9zYA8O1giy7y2lik
2+VJizwflysLD7RNU/ccRdrFk3s0N1Jv4Y6U4bsqwfwctt3W5UnDYSr2vfSHKf68
zBR3IDjA3mKafEs8F37L5KuEs8VjuII1Sg9PFCCgCTBL1aH5LDfck6+JyP0SwVXC
nzhcsHM6LfeqUauRZXj1OxGtXZx0upQfjKidSWNNOot4J4von18y8zxE489QyGDk
Iq2JnJ6RV9Sf13AC5MIFaIoWVMpMqUgtyKB4xJDWIZ0PpSd2g/FqgGHQ6DiTIvCY
OPYd8a0mZjQuKDWAYzH3TC25BnGbmThYE4kkG81gZ4VpstFfeNd/1n2/4DicF3fY
i1MCJiCFmO8UUNTRo20nqih/9NS/QldP6BFLp0ZPWfjfbc8lGx3vNY/v8U9IkP4V
Cods6zSLsv1eEA1CosqWUOZL8qLAUiHil9en4ONK9vzOVHFcw3TDJb7uXLUxf3X3
PytJZeTV4SlAvXNb2ZDYuZlX8nEhqmjAnXIp8R+MwnbzIuJbxna+t54a9T6v57VR
LQ7fFnjem94K3gfUN62cOQyD6hOO+yAtOQctIzwqOCLhG2y9cDWKQUhVyxyz16DS
Rn2GJwUTplql0BFWMA4ZCoN7lepS9Z+Oca7voRMcUWbDn5Ap0auHAmU/lg4Rhbta
EjshLixF8zga2eoFH/LE/GXqjr7O+VIsF/wIrf1WEpQA10okr3Jt2dUvyxJHELV0
7Yg2Vq+OJUC3gQFggdD7i5m8Um5LePC6ghizbCryoqJz84tC5P5f5IDfpddhg656
ufMOzykJUN8ozSRttIEkWz9KY1GuLmuYEAPi6GrkU3aVjlp3yokX+4UhQUpItDxL
LtCQJH8LayX7RZv/0TVrhVrcJhVthsgym4m13xeHy+9vmIFV9RwzJH48uVKBvVlc
s9jrjdcTVBwhF+REjBkJP7upw76SVtWQqzCQSQixDtBLPO8rC+Teyq0FfYaliF0O
OaOE4jtFOKlkvfUjtpElicoZokdYGorKaEaqO+lOMEXElgYVtMuJgjBaVV0D2mfl
mX7U0BKpkQplmSJScBDCdf1Rez+9XzHPs7bjI7oJAEcXzzKlGUh7GWiq09kB6aia
58Ati5zpSBZ052Hq8qi+DVuY9BRGMUDRLgZr3QMeie07yTpJaBQ1CorEJEsoHeOi
duyz19HaOcBarnMUmxh9djh/XKu8465zHIQFIQYRErZ4dZseifs85BuUlEFCJ8Kr
vNdp0imu5/hLzDiYhSbz9+9oFd/EPbT+vZn+ATcRuFR51u3V3MPpIusY71BItLEV
IA/W7EhBu/s2jjUQi8TzSCtOBobSkcDAUK1gkWUQlbTDLDC+g3IOvF3B+8t/SIAS
hXoBl0QUuph4ySzwAwY0+mBjNX+ZRQyyMKzx/iYwdalah3rQPveg4SoZ3rEAc5Y0
iYcJuB7NQwqM9f5HdGT67RN0JDBg6I2sjCelfT7W+fESuwDcbDNXhXXnFb/h8kz2
/rcrQ37d/vc573POb+gIhrxevmvLQpyL3MyIcah72xR/+UHKV3PtOI4i7LXuYF77
5ahUXA+jpE9zDSaFlqvQqk2fqc+8dUi1AXJiunEpGLlSPKVgNoMHwOXBFh9TFDJ2
lk2J6FGMFrKoyXOau95Yphr/y//C4SFIcXYwyhRgZqaytkw+to7c/6+cXLKYBKaP
6D+oPLWX22N22bPYiV6iBK8boo6A75jVV10gi2rLIYlN9m9PkWyYyCxgZFIBXVvO
JBlEX1tntMcWhawKliCYVcX9FxPCftyDqFATON0AC0yMPuHEmmMwOlh4LDD0OW6o
NHJo5HU3AJW8rkI436tlD8jr7QZah0pSnLC0vf3lwGK7dqQapRt14qvOosjOVhFS
7tEXJHbFryhcr5/R6lc0mVLIspTM8jGKc/RbrmwXSACgAEaOgP07CigkrYyPY5OE
2kOwmgYAzOdrCFULewr+dIhSJpeqhl9b9VEuGNhWU7Jg4ZYNUoZncCXMkObUvAzT
1ovw/rv/4IwR1/8V0kVA44d+0Ge4wzZ9i0g1nnyE95IzJqBfo396EgomxzfxSSDD
Dv/dqtZIoa9Nm9dgNZlGwiAOuoFF9lR5jFgjSmi+1Ywi8V0LktsHxseggirnGRGH
p7xBBHqNDl858mXSYlMubj/NZ61dgVAkRF8lYykcYefwyuQCRb2FM5/sQTROWdqt
5sE94P5V0ea91mcIwypAagKeryEC9YGLaZ6aN5Suukq2QApBMNqqdRdxUwDrKUux
zGbS5dLsyamm8cnr4KmvwpwGiMU2xm2O3qV0Fqgzn/9vLuGjaZBov3xrmT6hUAYZ
/Ff15Zpqz8+Zs5R5CfApph+VBt7Fk9dVYodHNBcAA9raT9byfShW2oqqPIXiWnFd
bCPf/uBI0kgdJIxm8WLgnTzdD4ALY8fcXoOrKO0ZDONtHMl75tivMC8p7Y4JDrQT
JRg5Y2zY7wIuvO3Pk4KKEIIu/aPDWR4622Oxk5f/jsWf2jdHM+u8/UR3aRxSK411
RXdYaRUHMlFdlfi4AwQGIumdzssVR0qV4cpdeD6gIClBAihGIb/5gLplGnrcjV8Y
Rns/pvLNj1avyctRHI0T8NH94Fcwj9s6bCV4EucQBZjGGbdRwkSsHlnEPWOkzIuR
+qUPb7xI9vK2idhsfZCY6BsLvo1bxFWANr0UKhxk/LE9PqvBN3XOcrwWXmcZkQLR
mr59MJTyqg5QQC7EaLLe0Rnfgf7BQzcp4ohU3lqMO4W3+dUyCiHzt0U0Fd8Rq5WV
ras+J2eIQ7P4yiVGKoKoLH3aos8khlymheVYNQ3ufYrN6zo7X3hWFVttu8LyvwTL
HhIDc5rf97N8b4TmB9tcVUYSQsxCILMbMHHuNggV/dEtQYeJf5hTzpxEJZtH3NmK
BWX/Lgf8sT+hXTowf+asI+BzT6XLFcSBYf0zXRSPRNOz3Kj+ir6toTJcWR3VOHGx
KRUgP5D6g4lwTVan5hiuolcrKfpn9ZK5JbwdD0hK0oEiMRVMeFCRXIa19uMCr4BF
AUD14ShIT5UtHMWfqrnZndyJWdRz1e7VSaFWIJHAW8ABlRFQ3ScLNEJUqlIH+OSQ
9igcSCylkwfQAkgONPCLTZzSIIojFUnaPM1MY/vYFiqro/Th1mQTRhmLVsgkX3Bz
zCVmPI3pQ6IeSf5alR9Y1zzv7qeHtBen1C0r1QbqAQdoyjf9JS+AOFMth01lmi2u
orQ2YPLSnADTQjQ3LjK+7l21oGBRihat0rfBFoQKq5iVukioBMOnNxFD6kMXA2Fy
ZvpiKpw7dDKIHQ2tClrSPfNBn0getAAhYalXjrSr1BSON/u7UT85UTWRAbZdeECe
QTlUBrhiY3ji4rh1u+HraEurUIbjmj0DlPJ06fOu/+OHyuTvn6uqt5/nJW34ONfj
2BBpDSb8/nJXYglm694J2/8zGg77VrABUMBjaqwaFpTUf9qyCXb9Eg+iGExjwWyB
M/qqdazXh7WmNi0PD57hOpeYj4GaCgy7ukS2br9JL/EwfRXJ7oeUFtCQ9mnSdvRa
e5o6T5jnhkl6aMZgq1Q50poMpP7SPF6eFuhCG8AfESfaZfyMy4HyI4WbWKxlTRrY
cR/oYiaesneRGN3xrmbNaM5KE76mkw1eEMhlpk8z3v3kp63t9Dqi1hzCz3lzEvJ+
gnfRr7fxOBPd75X+0WWpLRu746OE1BCnG1uB8LUOyJCR7EJEzHoxDquPVgsS9H4w
QhzMh6wLvZj20DwodqnmJvIA9DwkbuYWyQNMhPgXsVjb+W3J03uws1ecplw56+go
sNyUDYv9BpjQTaq5M6c4Kkxy8SWiyloivaJdhyS/DZRrWRoM34SkibHxQiTDssX7
9ThPtY+WIQKsxxLMtd7gYpqsnma9PuJeefwYH3v1pU4boLBFssOoT7S4R3yTuEzz
zcYicU8Jnk8NGt9FENX22EDXcx/O4dWyFjW+2uV2rIFX5265cu5gEmkJLahORj1f
g7xBMepbxYsO1jMfxOwlMTX4rujVP//iS/jlrbvihXMC7UDKBr/Qq0gS7kZRKGJ1
wx4qptKgZqScQrS8TxZsHblpkVztGRu2RaYtnMmRljM+Ut9rQgWLmGwHZKYzA752
aQdY9lvPol+MOyPUNq6MvZbPYugKkzeY1ZuwaVnsBsqTveibG2nZ9/4hj10GCjJ0
8AFrGSmiMrn2KQdQv8ekBDREYiBDUSDVUGWtC4X/yT3E4crdAabeOjWhnpwpYX1v
JDiHjV0ypuSeyGV2qxvx+3S05JlrhGVLF/IunedmiOBT4vpAdYOANCHaucnFX8f4
WoUKxp2kW2WP7juCREOWTXlzvy+IMFTeLzn1O9U8yB3a6zksDQmTMFSiueRhuS7T
NnMN/kvO4hUPfxG3D5Uv8Ll62nE+fHzOTSmX3pjnjqjImYbswCD/dFy/8Qg18/xP
UL7OqLJAVQ0weznaO7gEOZL1mk0mnqTsB34JE37jC5WUY/DfJRXzGnQBmk+p9n9U
0KIDH9lvrltUigQAy4/GCuikjQtr0f16PttGvBnCg6PQEqDNVHKA8IbqydVhUxY3
1AXbOop+wCj6WoFmnjbFQqkJySqe9PjRSlGB+q1YaF8QwY8h97EpoWmrWPRxYRCe
PDVgv6GNfKBc61qyj6kJoW/U9epFrJ0LGxU9tBzlW2R72t5FOkWt4JB1E/5Vx9X8
V/PYFB7R1gq6PN1832gxthXoewZq49/T/2rSWX3j3e7tUCuHtIWULqF69AQVu+/y
mOq1OxEzFxNQ++wyEiGniUSrGarwMIKfZblojtaIUMtF5Xkk47nh96lrT7gLZ8aN
E04vAFA1o5ZVoNwHOFaUUKatWHGm9Fyj0+gy2xtRT1dA63RjsqAE2Fk6GyeLmzTJ
7B8T684sdCo5r5TOeknEKQfP1zFEYwAy/ZpPNv/wpg05UP3OXAKH/n03nEhWn0Fa
OOoBijuWnhXregAm5LiuwKO6GCaXCy407dGx7ozjB2vSL1niyVyQOTSlzyV41tef
e9n8qV+Y4Jk9uWRYT2lSeXdE7K0VZGhTf5W/t/jNYcVtHK3tYGMqeG+LipSPil0x
jqJpwkpzY1mLoXLZPn0pw/igkbbRWYDj344aJI/oVJvWvnOsvgO6imfHdoQF9pTp
2k13IPHc4vjENkx38rqmd21+cJOPGfTdIGN4shgtMirNXpeAuZzzttJZlZI1BKR1
q3ADYSPL4rCraJSKrZqpYstt16i+hZjb3NHNVjCp4qylBEi6N64AODxDaImuTS8a
Kma/dbuOnAMSmh7T7EYmBuzlzVvOEWbd3CYqJ4mJaV1jH5Mo8RIc180GW1n3GHUC
czhsMfFTW/DOP6IAR4xa0g7olsrtJ7RFPGAbk43xmaIGJHKspWTT82hiIlpM75d7
GyQJHDJ/n4ejzOX09FV9xMBIxIWu7wZNQlDtwPz3IwjMOUWCIQG7SbA4UZxmSZhy
W6iPAdyBeKM35rRTJYKPs/4w9YXxGxvus8uP9se1JWwopont6ivw53Ay22vGW+HD
qHCo6ejIXVIgdcsJPMwBqdZogbXDxDgXGFktdtkg0V4/uy51FM+8L20V0+tPvlNe
8I4tXmjeNmpAWJEbJ559oggCjYN/Sr9Z6XEv/Ng8qLQWayHWEZl1wsj3Y2AImOT+
ZSdFFqPggZy4Qj203DLDz4hGLE2zOLBuVVXf+tQMdVpYG4EZ0kVLBFaCwT8MOyq0
GpIZIWmgDWjQCup8SYbQtcbrJIMl+NOIBRejkNm4v5Q6MjHj0fgqT33EDhSVmhZm
ajXtb9qql3QiRhEpleKTpRTkdv7MeVkAEyPtdJpPP5zi/cVtxWk2iOpUzzsbkBhN
rBrqtoPelqKgGddSIu7VrP3DDy6NyrajZscumVKXP2vdztugiwqg5j+QGfbqAPLv
58hxzbKApA9hEZO5rPNj2HCTxsjsipIWBXvt8Y7AxPhAqCaYOtg/l6N+xZPnT5MO
5BKFDMqDZB9Dn7W+Io+cVuBdYw1Lxnf6O7SjkXTgWQznVYQK9OxuNRHVb7YIqukN
FUVP9qV69IpcdJ6eSUhXhG/KAEADgMxggWbQZBl2eKvy0H0NF5816X3z9mQQghAU
I8cr5ZcDabc8V+r+DBYtgCd9PYBI4k2EJpkG29oKzNG9la9JfOZ7jlHu6rcbrHUN
O+eAdM5hZnUozgtJmKtD75IfUklRrX/GW/JQCXNpnHL6tSKWHEIT5KcOEsCShivW
0gppXoXfZJruSYt8+nbdfT4IIZmy6E3f+UHCO8KjnnCDEeGpsyYBpqRviqx+E+JU
UsZ3ELlN4PxBhuNP82UNVxvNo29Ilmqzn1z/TOk0MAOiWbbCDPghl/D9/Wo+Tdt1
2GPd1K2YKoLFwTCNfIVz63dMteLj+SzB5jLnl4xD9/pbHr0mV2GF5ZFfOR6k5SZ7
EQdjzV2bDf+rIeuSW6zrYSQQJZBDyFSFxpbMfMORoywgnwfvgiVGqpAxV4u2g5Lc
YrkVr+2kMPdeoOSIM6MVFEibp8IGeeg2higT8gnpIO84G+v6WeOnKxJEIB1VOgpx
bntAQAfMpTYD7ay5oQFrSH78KhNfy7OBKAd4rB9pJAvOn0rbiq75PAdbFaRaRLJ4
fxUp6ytiJ9qh43qrrlxSv0/NFD02d6/Gipe87FIvHSbCp97S4uQ+s+En+kQITuwG
LWwYJ7pMdb7A/rEUnGsFSq9O7jx0LeA58alBAbotwok2lPMu2EyOVh+KiT3C5qk5
HWJU2IL5QAAxBHEO0mwUfdVPGiqFCH+NyodWkEl8NNUOjJA6rHpmrrG2AzN5fRbX
bSOv1cC5uaL1pNoWNnUB/UkxIUvrwgQgMdyhitsQYErfQmJybMQUvmJEgDDZdfe5
1HkFzZc8GkhRv5f6ehTicNbfh9GCASXyF2EUSZz3Y/S0Q3PsS2wxHee5iavXBSoq
Endj7+xrj0PnC7HgFkN5ljMpgznTPg01VTOWXfPUIfGIerjcP24GKwNiDWV8ApK0
fA8V53uDWjkCFdkmmD+EA1FlZQcoprZbRVBclP5i/s9DF6NAurbrK9uizDrcctg6
7gh9PI3vh93BpeKoMoQSiher8RtBfhi+VxJ74tyOPI797ltJYtx6dY2aZKsKvQ/r
fDupBHghPkKNMs54UMr3iy1BAkbUGKMTvWIUkNmdqnnUjlYJZp1sedUNLa//an/S
FA4LPoLd+7T15unvG/KBYRDUTe0cKIfsdR9m28M5OtUKaHMTt3ERAV6JjBexbmyY
aO7Lz/HPkpxfAjEm0EQmNz++lqoJQgxNJSSDfyjtWZdAqN3zOEPHkCez2f0vz2JM
R2xMsUSu9A1s/U33E/JwWB/Qg56QkB2Sc0jRzPlTAaur3jZJwO8wjFTO9tmyYUTt
lXKhLCZyR8KYTwt71rYwVMtw5uSV2GcxU+k5rcRf8d7R0JvaYSQevBvRlRDKH8oo
8sfxKgoQ/vzxHcWYa/AHNBR6BjQVDTpsnsvoLMkc3kboEXjhC6pnzOdWwsubJ1NJ
nxrPQ+nDSf23owlJDk0XSYJ1NIlICOYfOwd5T1cxA1Fx9HPpp1jWRVDirtzNfkfH
gsLpPTKNeeCmwD/mUjIYCg/XynxjgRQHV9sGFHKy/BRurLRRcLykWTKliPvSy62u
EKXCDGihrgNTDZrdbzWkOSuHgzyt1MPAuc1lT+TW1fTb0lG4ntmFe3qNDQuhCEuf
184ksVA1OYW1ZdiEZjslHva0uIN468YbaY/89hXxiEugqBPYYPSl+6hJcGzxTAD0
baPG0xYxDsG5osBHGK3xjFbFd0+BmWyfMTq9OW8shRU4ldySH225P+JpC8k1q+tp
DmHFU/RTi5CsmNUnJwolw5A1m/eB5nLywrNWvSa1Spd2s/sXq3czXrp0sdD/ZeDl
V55e1lQBtugizXYfXjM3xymwBSq/hmlUcEKgaFRdBX43l54c27cAAB4uCphFmis4
tymqAHcUnQ3H/OZ1YfIEjCjAgvcUSFvMyqthBoFSW4DfUu3oJuoVUdE6gq3i9XmX
xjpPuLUB8zechXKP1PUZdxU4sK1XIsaGyYVwP9rGzanwwCMNaGh5txpJJe++Erpn
cMOuW1u6OATAmm24vwpp0m8BUtwbmSsYO76MSv58/vI4vGnn2C3A7CnPa+7rEVRO
qMTZjFHu6tVYEwpXJhbuHo7wWthRLnYQwSPo9ufuZu8pSEg9rwarOCP2qTbQjrba
WPGGeGKJRYq0mHZIUKRL/ZfkY7PM7/bLhBUL9EgaZmSuz6gTfZXwOfY2S2x4itdi
ilxSOajNJtrYR5Kx1HqrxHiSLRocJXMNVUk5iVwGwgASw95+jCYi+Q3XX1Sen0GP
a3sfoWAoR2pX/tOs79ax0ioL5oO78PQfIQwd0lX/NQR1RvmzGeGxRAA4slKeSUOI
QSVxgAxYG23wEKV4rBRrWgHTj0rXa1PLKVQ1ArmaJTsXYElWRRROVbswRkE+1zj9
z9rVEZODCZKUpD+7NQmGpcS675ySVe2DcCDDdeJGjdCqRfsHb8s9WcCKlx9B1bs1
GDs1ScgV/hEEXowgj08MVhl1dYwbm3g/ea3gavZUYCt8YssFmcT3W0G9grUpM2El
arq4KxrRxNPz6R0pwEChUt8+OozSyBZh7cRemxs49waauNzdxWQTHA1Jeetq+Xw1
783AYX8zZj0mjFktysPtJCfd++gZeLLty7Wuz9CVO9EqDn2nlDHKVFwIkn/Xzu2E
uNmJDqH3GztwHL94Rkw0KjK8O9YXoUWKmjLAmM5OmlBDGUfqcj2WHp9J2XRT6HLA
yt2Y9NqxCYuuF0pgYju3jWFswnwUTNV7aXwXu7Yk05LR/2WxN6d6uB6oGflHSXcL
GeLsodbZqZNuM8vIziID88OVxmTr/SH8SNRAeCXImylUE+fzliiCzl0UR1zpCsHm
LSLPyjlNUeRnsUhc3vXMwAd7ggZT4vezRUPle9jR0tnDnZ1I5K3J5I5ZeGevoFvP
dxIVY3YuKveGqpfDYWtj5MJbJgv871m2r3tmeOFBMyvhsvMimxkpkprCGVu/KqY9
elWRg0ZC+i3ZW9Pp8GItY0ZghbNfviPrVehquCTELxH0pVs6l8e14REyDh5nB7Ha
Cijv3W9kfWkdRVphPvslwMQVOAQUPSZPJupji0xWqBRs0/HYBGfOHHXFzsGt/DQY
zK7uuCBL89iUDk3/jT4UnoGo61oOn9nMsaxC2VxBYO2BlGtzSBYvxiGFuAhd6v3P
Pyt1W75cqVWeqvKNIGoaraGZXvC+NZ6IwhHOBKeFFA8inaiG/UAc+gV/5N1LrWNy
TnYVZb1rmaGQ/YzMd12EWX+clSpznGWp9bshJ2btbokmpTqVNP2M9W2HwiLCxC31
mdDI+yRKG4fi1q9g+dgNlpDGeLJdZo2mnUSCzVQadPp+N2vcuBnz5oNKk+cAlin3
KVq/pEsv6gZzHbcDzcpl+3uO43+yhiKgCdEG2nIWsqgATEu7w/EoXfbKmBO16O6R
e43atXzeLlXsPVmXbrGntStkY/bN6HKSI6j2SwHNlALQa+7pdEySyQDrVAnUgg+0
SEhU6/kZYzjRsv7pV68e1+nu2mw6mUnqfaHjYM6LWW1ux/ogecv5YSFOUa563Iy+
pRmx5NRiJDeaETShTXr0Ekyyg6DiILYc4M84JxhgSU/xmoZIWu03mduSR0etHyKr
Plp5TTzKX4ta70E2GNpKY9gNPthAQlaYHI08dkh+tVmMyUUUxefSw0wHeKsjk22X
oYsoO50c+NFfVyOkwUyJqlLDGxC9xioQVXY+eFvhWZ9imzm9dJVzlgxIflhs8HrH
HZSsz0KS5Yc3q9uKDi4Qb3re7Wphq0H2PA+mkA5qC0EJxabfRaO+I9yhEpU2VbGA
TolgWg6qkqdW2abTzTYGdEwa7x3X0VGyY4usrmIwmNPdSytJ5yvk/EdMs04LHqXj
B9mFz+TRm6E1OFf80ZxTi8vT2lD6qbQeQ4bupe65gaoQ0MT6dj3t2xCKcSn43/tk
9UUKdpUhCR23dpQKwjiqdKFDLmQx3MllX3sfXJwfHYOWMJt+ETcLgDYkOpM9fWci
L6aaS/frWPYKQ0zq+iz6kiatgj4i1XwAg7iiUjIxd30DauN6DSONGzUo+fC9R4+J
cvyW+3RbSpwVi3vQxutrVhqVLMTGQHb6WjG6TJxJLRcsowIcrjZMvyLMDOqXeQ3q
Ynn9nf4kJZI52thYILLv0gOu6fh+hfFJAaLiFCVBXZxdFVtjNwBTpF64nnkgWQt2
VlGKxe7eTqSg0XsiB41dgm91l3A6NeDFNW41U1vpinFAnxnRdlfT8zfm/adCxHRm
b6KJiyjm3V/83OUDNdJ1diZY77ThoHaoIqWgHu4zEx/hnZ1Ag2Rn/mCakuDFqRd/
0mY3mcVqNhmyIUtT7WucR/aJQl2tG9TwBbf0f0JIuZ4cWnCytGhGItrQ1raj4eT3
8q7bwFDwBFeG4onCkR/p2l7gdZQwyDL9RgVV6uCkeFQG/S/8J/VVMTcSRgqAUfrN
NmvcVR7XQvH57/4dKWZRUf9tVUQCBKjwBS/oYgx9oto+mwUBh9ylEvlCmlI+32uO
5EE6P6Tq3aRUsDTFidekEBzfNIGVRcx57TJGRFtZBirtst8BCKvNPOxvZEdStZ/C
zVUlK7ZR99qaixNJ8IyDIqc1uQ78IPN/STnwYYbnyczmXyIVYfq9q9YoximgMW47
3VF5OoJA8n4t8PkMfWRkw55TBS6PBUkCNF0HD1O2aztOotmXZIgz/gGg6aAC5q7g
8tb9IyZQSomY+efQzy3ZrxF19rK3OMKfbcYQj/zaTW+V2plJ887IYKZ3ZGuRBaEs
QvBboe/HW8rCmE13YuWed505LR0+EwGLzReyRbNj9OOOv+oK+MetlsjMDSAqKfTM
i9P4ln3mUW2FXipcZWfzl9Lr3X9s6f9Q3JcOiUp9mKhGMdFoYCnxtnDQXLu8YXHn
VmRCqS/xSkziQ4VN8IRbpZsfXTt5YiNNfZIvrMpsyP5v/LIwVtlNpNueR7kfui5Q
dXZCL07kzJx8BKFsyuVmSwbrMwU7H4v+aCnUCLzJiUwsSmtfXDQA2Fac4OV9XyQR
eZTynano/Mk7b6DcfGhFXtI6WorpOSYkArF7+xvgHIcU+80HqsVahAzGwpwscihC
o3wvjX29C/9Y1Y6U8KECYbJ4ugYBgytnV6vX87rzy4uuSGopzGLf6fLAQsKQ36oY
Paxelz5IqZZKEWlY3w4aGExvvNogCAAq1floRbPPueJ3qqTzI9NFw7CsUaRHbmJd
CJCm1SmxYJAHSsGt7KzPwI+7dU7/MbLg7dAlEH7Nh9ISzSqyVzsauXjQjsKPgPNc
XJ24/PiWw3L/UGMZNNWz2db5l7wW+0p6sYTD+E2uwl1MwfcTDMODRklcc6tHu+FI
+QtNB/B8k2GvW3eFnuUeM3qFdKUgYa7lx5kOvEqJlHYMxoalps6cEoBZjjpaeilS
SumRUCwA6JUBog+L2bAR1DL4Frk1nsi9MgMm+nwkmFPJ1raRlKQVkNqLRSPH4Nl1
zXKLsH1vbXs+1Pq8RUQDUmlQQtbNxw5gYp+7mFAWAmviR1WAyFBJqkDetyIdZDbG
MNROda7Yb70WQw+C9+gC5PT2pPPjWtG8RWJrPePbZsHSPVmjvzjGpY1mfF0O2Uno
epHgck+cmQo8zoXB+n6gXqQ1snJKmfN+qM23Drj5HzBZOkk5kLU71deV2PnnECzP
weYUOjbV5TyJiKNGONZd2tGbmJn16ORCmn+JE9tK/MS1GAvAxVtcdnQvFlx3WvUP
ViYQQ4Qx5R3KxKSzsMmKvc34th6ITwPcHY5UlUwquHG13F7LG+ojMAtvVaZJvNl0
Ipq/kwd19opdDK7yZNkUuC4vp5WJ3hxdfAYWsct2G0SrDLa+ZVWeSbwwBgAWihtI
ATD+LWLP6ruSe1ro/8xzmaRYnvLlwx3ZEdnSmZN9Bz/hzpzJ/3hLIbiXNIUaKuAZ
t8hINyos7KFF78StJOclJZsJ+Yjm4xnCoXd4RUU9AiYicfydsQQJB9KGACUtGckW
aBVs99SJlPB2eMOaxGm21Y7xhz7K+3K/HhdwzI0PghC83lePm3ocwvVsiObBe+Yh
uXV11aN38anMh73/EC5NMXO9qdxPRhGid9VnAnaiNxQSgEa9mAjMCiYGYsZZBhpL
ob4x+YbMXlxNLy96yEPqxvpE52+1l3pww5TNXx0Wudq9jPXYbmeY6zRcmTSxS5Fx
V/OF/pyAjg6FyYFBv2Q01Mlwf+7PdSYndVVfvv7ePwaxEoxrVotkcSavG7DH/AfX
ogDT4a8TPNNcWI12c5h8T8IBY6p6dNyWjVGoTfBM5lAtnyULinodIacXxblA/0rI
zxyLO4oiR+2mGVRtrCXyxzyrszy+pQhh3dXTaBH2ErXoFV6vxJor+HoKHIUkZht0
Qvu0a79FtDswnbXEmMglsa45kqFDAxcxaDasX+bO8hol7BCzvj0DDwOskm3AGuIN
2lMDxiIPDLHPAEXUCjRd65Z6UidssL4Ep+LQebxf4wOt2JJxz5bD7Ce5+N+Ej1Ha
WjRUtN2tukbaNBAu2VYwUGcfN2ZAiiCjGxrq0v2lWN8U6o4n7FUzt9nIKCeop8AO
4RhKVlEmPLOU0Eq9AKdkSVdNCyB9eJ3egMvI5mzVQIqT4qD1HGq0RJr7kb6YoPVe
HhTIR5CjEbmO1B06b1ZhETRXBpEXe0f33oyWu2Vq4AoFdECc+r0iugOqFGEq7jVi
CrY4tJuv48iCW/UpRpy72Zi6xFFGC0yIiFl29GyXw2glHEyMW+vtAZqqFwlJ117y
Qx6vLv9tT6Y6TVzlK3TRoFf6auS3duXOG/NeDQ3bKhgA5JMmOJYuVN4i9MBtYsQ6
N6LkmKJZVcpHO1gNEJxMwK77JddEPcPPN4dIw2XntdVsl5Gtz0t97JMJWsAs6VEK
LKjgM0iIgCa8vYoKNFBBj1OarEeHKL3P9J0iIjc1+UyO7xAgTQgycRIvPX0hE+6N
zFNuOLh0cMzoumoQmzDHnLzM5OYmcbXnOaL3nmtlxjLC/r7fiiiS3WR68bdJkKmW
QriZQlD8PDHr0c0EFIXcJdL2qgnAmPY+1e1l2wYEMJmTis2N3l+118G5ydMtg2Hv
ReGLS9CLbuwRn23JlGYjZrtVb5TgU4lYJ19Oieq4/V4Ppzv/fsvzYgqxcwNJKkTZ
rqYmCAZ2QaTmU2odjtQYDC4Vw2S8Mbyh1y2J1miXkJczkq/luAl875Fu3sBW4aph
F8MqMuVxXW+yW5TW6g6c/PC1ur6nXvyclBwRcNJ5ShZIGgt9eRVZ4Z9tZlXaX+F9
AKsiWocj8sFvAcFxahrko/Hwu/Qtyb/lEtR6FZXoAqjrhXax/F5LwguVDuoqlH+W
Wc8GpWtjx4mYOT0cb/Hq9LldkbaxkUuZikkBw/LU1eD3zqwvKowEy4sqZrz1zMPl
jgoqDiFIBz5HYp6T4n0+bIpDDhBdUlKdk/9UDE2d4h7E4ejE6sqjKfNYEjSZG0E1
x+pIJXWkmVfslkmin2amh+iJxv5+oSJzxS2H7d2bqz9ctmy8ZlVqmvtdb2OyKDPa
DibmS/dPZ932yRikJ0gQJzkbR7Cdw0El+roZYFedrX5bIwxl9JfWXgAdYrRkr6jH
P/PbSX5CjzP6l0CKHnfYHQ4pb7W5XuqH50U1oEu1gIPPqkQ8o8+8YBpxfu62N9T3
Cv0M57/llaWhdRcwieGHZUXz6eSqdDObTPl/7UF/LkEdsbZBI2ybU1v/c0zbFstX
rjBdV9A8Iuzf7XtFqB4ie7zYs97JVYbkDsqsROOoywNufbGtbTILlxghgI10JApK
49N7Bby+Ei9LcCsGEFs0ZB74ObqMv6gDEOjlkG/b/zO1Y91MiNX/UUKkSl1yB7lr
OKVm++28V7lAZ96jNJNFuEXOJ/D3QagK6pnRPNSD+W/vCvIt2YgO7HZFMuunTc8y
tkJnShPmb9Ajfin58QtIltZC7tvmfnyyg5jDghbzep5jK0IE0zoVn3nc/Ecoms6n
5llEtwzfpkQkjAaTp8AqL3nIYx4UvnjVyi2ppl+JMkQw7tAcbCT1c5RDZ7TPo3jC
bWniy1hgsWUGVKPbTSSCacqO3R/vfKiv38YwfcOQvUUyKx5PodvoV81A5Ehv07pQ
qR7zMt1pb5uGYW5j8cilmHk0VHjOSZYInWAGeaXC0zA0Bfq7T4TgHh6Hesdze+aZ
ZNzpjassYvvIuI3/3NudAgGCus0BBVcdYNltlsfbB54PJ+xFhghz7iZ7Qo2N9gVy
sq9pPHBzCY1WipVNBWFfWPWoLoeeUTFU2NsVVna1tTYuchnctLseqqdtWO2YVnZ3
ZrPwxB1zVVI44hqx280V5Jjl9kfnXYPRt4zh5PciGQhS63CvaTBxItx+FUvBQWCz
GkpR+Pwt3IbZ+9p0F6poOw2H59Ge85XtWwx3AH1djdcA/9GWxKUsmlOopmEkiVQC
G5CVXBh8oKTLnnpai3CfIEv2dw94qT5JpJg6rwTlEZMs7THdlAYLEHjiJmssDpt9
n6kjwS1Z9L0qPxlummhKZHtriFYqoXiiRMb27vvIX2s8RivnldMvtbaBk01QUXi9
Qwxhp1trtMgqGDAaFApzwH1slKwvTMzGVpeJGPtadMKPQDLkxbb7AYs45KRjNyHy
LPRTa34Wyq7BocmW8VTwRDo2QYVVw5UatISDGLeXshoLBExHufdBuGbqzd6DS3xl
C7wW6VvPgWbLyKnoLvqWVAr0kGrad9fTqig2pdk8JUzCi2Wo5UsMFzkXKMQ5rkp5
BvLcNe1/rGtSOK135RBprKg6BfmSP01JjHYAei26gwjCbN9IVe6Dd4XUfn5GCrM4
fFpQCCMtaz4/4t1JRH+XMoUdIFRXH0CdYb5x4wc+MVCPWZt04emuG4YJYVHfZZ2r
NQ1AIImYfZU3JEcg4xgZNElo4jOWSmzdwLLOFXG7mANQKH85aCUPknlWpB3sC9PM
K6tJbkNAvpq/imo41N5ki92oLESVdSfZ3hY1tZkM/2Z03dmnKNw+pZ4GSYT9CtDG
R6sJhkxjNZotwZVfXJJ5twZaQ6QpgTFqjF4JHckcMvjZBp612NdZQwAXFkskxw8B
MDtwOE9gXgYgWHC5qwcCWsxHCUXT/rygpc0zHkSllutkVq5BZJNehbUxnbU3j2jt
FpwCpT8FfqDKJJpHWpDJNH1UHWkoTIGOoMm2M5aEJSL/WmiKpztwF+9gj6WRpdgF
pKoNErTsNJwjbdCq2ZQ3Mn5I6GVXBfVEXukKBt80x7qhwRmaBL658zr2xSajDl70
5uypk6MVuFZxAIo2FQcZM6/dOkdrtz0aKN61/TxD6ppXKir/JlzMJ89/3tMC33/H
Zg+kSfRHzCJPQkdk45QX440HxDvtDdyGy2eeCb2Q72UbibRIbGiXcGQPsJrnI3dE
gVwrfaY9TCbsd54QPEVTei7VkFwLdxMm7EkA9cW/UuD03tSOzokOIx8NKB++rHno
ZaErsG3EscLqBeHDJJeCYQ3A5uz9K0erNEm4X7iU9zSF+EXaVXBfQYfAVU1yChtD
28GE/P3J3nzbh4NmeecPrRvLyqAZ/ApxmWGJnlfBCCE0Rsm9yWGseigQjBWyQfnn
EIdonXjY1e3vISQhKoieIZH5mtedtoUFxd9wu3UWIsqR86BjDyE05MSOzzgTMIr+
KIgMIB/tdlRT15gbvThGoRB9oKGuqoaBlfO02Hhw/1MLphk04WCUsM4YExdzoApa
WgOHycE/vbtiQ1i7UTxs71gVGndfjbH74THm+0NiM32TVbtWzn4lL1UxWn6ypZUN
csuJ/4FPvhzlskTTK9COjZV9mruMoB8VVEHz9c9Rozmqzsl2VDVAhqhOeRx0OAPt
MMi9wb/RnjK8zAq3GkDmRXd9xEPBQjnrbju90PMlyVt2sRFriHmAJpzQ2zN84vFs
btSJHkFxK1zhosfCSObRtwE4KVjXN1ofT9/YYWNiTJpj5eA0FLYkgjyLbJbeKetX
MRA4Ucx1x5MCSYBz75pPgM/BXQwr9LsGXkIcb+f43XdE1hP1/Mxeg4dV8dVr7qdM
ZY1IuxTcEyoarOIFRgnrkHkpgE34qR9pdAETRC5DZak3gp1II4p93Qv7LIRfc5NL
PMaVtX+1dlzqlgNbP+LwBuHKc2xY1OZ3kM4HAg2DEhn3uZem1lb8c4FJ7nSvtg66
yOBssNOdkNZ35J7H6DEXxFjIbRBvp4TP6Qz2wW8JQ6xYuW6CBKXVreYuyEUSOznv
UmRMS/NYVryu5J6f/WXEUeV9W55rbdSIjgPJTdxT1O2jVL1GLMtAX4qK5a1rOBKR
I0ExSeadJyRxaDHtWZaK0k7+r/Ty9hQRJXh9fA2Ve8TJKzDEkvFWqWf5Rw6YQ12p
TDb+78e/b6yW88a9sAoTH0D5dFDiK/PFOSmQ9Q50AfNRl1W8UViB8BJr1CXeO8Wr
c8aJbiUwdweYpRArP0imqiy1VYHXwYSmTCcX6Q6llk7gqnZZT4z5Q+/cfLlN1/Yd
UlWnZdsmaIKw/MPaV5x+whzaKhP+jJW9SPP6lbzAq4vHpwafz8pSv67k6FLzgyPS
FCu3Adl/RAX+8TWVYOWYTVJmWIOkpNsDRlJ46TFGYyHUWiTN46NNX8exXTVwZWOO
mxE3t2tABYQuPd4DCLgErE1IXaDE50hW66hu0/wgx1doiOU31+wIyMo9LKvZVtpc
OnhXkZGxOiZXTwmaugk/jslJBWkM1NIVSnHwUQ0x3oKUoo8psBwlTVZlyvdtFobR
FfN89o8Ao50YpyeX6eXFznBBH4zoiSHpt3hoDdhTd/CcMzTWAMSl7GInY0rNQIza
+oa4WCs3wOB4JgDyDuuy33wluib7dN+S9fulmmVmgKNJa+D8DHbdCWVav44JDT6F
CqqCEkRigCaoX5mhcKe1BVMFiN13ZDOzFsoXRHvVoz8g7PFyU2TAfwQ9Bl7Lo1yx
WLwE7sQkvWoT3QzLpexPXrzXZ+nEOmC7k1fhRq/MPUIHJ1QvgF7LttHODZBEl3zf
dEWTyznuL2kaFPpewXDcR2tBw1jw4CyaTbhzdP/r2JSL4l9L6wXd5JRnrVFSacLz
CzAUp/f5JTpU5hYHe1kF03FaBSHHx1X+azYeAJXotWQEvbghEdgbDIRAULuU/Avs
F6vEwBjJ7vpzvay8lvLLLHo2Q6iHvGMJY2BDv5cbDr5zfnhPi/qpMq3S8E/DVP2q
0EVVSC0Mznupt53L3mCoX5SfnSuqb9kfDa72ueIpLTUCPynDj+5Vt+vqLnTuOULs
402erUa+/M1XxAsnhatlM3qrzwic8l1E1HgI08uFfHG51fH6NzFY3fU1+f+CkLyG
c6mZfac7tM9iN49AAwAh6urpolh7JMQErjJWJugkAVNy43C2lBxN0Yn1ZfGAVRix
MQc4WeK1t0WWhq8lhd5H/6P/BiQjPsXRijA19O7EtaItuhnDOOzq2fEDd1A7Ywb5
FDNFehC3VzOj+p68sJoLjAyFF8jyCc2YyECqdA5pM/pFi0VrB1ctxp+LeL73CYzF
wW5s6rkD822mjG1U7Ebqm8+GIOROIzyD/P/M8r/I/PS83xKguD+Rh7jTNUdzvvJN
pP3q4bNDtim8X2stlHwRvHc1Sef696/63q8phtQ0RuPQCUbcWfDRiNTW5zmPpBHH
NJU1vw4mndr9SSwQs5zQFSyxo9AwiT42eYl2mKBnJtbO91SalNZrqh5Ti4HS2zFu
6tgYHQanzCcs08LjTz7eQ8VsGyjVgAuTjKKnpHEFo6ZcB2xKrHrF/l7feBiaXWI4
VDVe6/Eef7f1V2BaRPY9xePjJIVzcBx5AEkxKMVGTwtOiqBbym/B4rOkTJBmV9jA
It3QR1Pik/0Rhx6kuK++3zOIzfeEiWa28fCYDRvcF9ChejRHrogUQLhMA10mjHAo
X6XIf/ExOxxFBnzNSNv5L/kA9esS5IUh2tN99kfquCdTRNBRZNO1/r0MoNUakuEX
imTIj9A0EuzqUTYeZ7fKDRTLbg/Qer282ZGcziFUdTjJy+o3yUWoPIaOho55NK2Q
xm2VM4RmVGKSaL2cTF426AWUhcT0V0fCVuBYWahkJWEC1W9TfsHT6JyHYSGdKL2d
23681pIPaQB/G3wivV/tPsf4+VqdvySiJ7xVHAfWs1TDHTY76qpBNvq/E0nBUJUw
4EwfaQWYLxWegY6bMSG152ZNfFx2OgTNln1yJ5HkxUqKgf9ARk5VCmOxga7+Q23t
DQzE/NSQ/DmysuM1gRQYCFOrGkyp4thRY06fkzghgN/WgaKU2jsg1BJqwwi72csI
wGAVMk3/RJCsimJuUpdWBEvrJj6qjr3ztza1XxbDSumWRb7d0Kv2ipPW2/L2b0tL
Ylq9+Uwvxq0ce610abApRYRBCMZpsbH9NSYgn8gSOO+RyjPYBv4x3c6t9VF7xS7/
gxI28ZsdbF1O9O7X+LIdYd0jrrpAlFOOvdqcyBVOh8amCI3st1LcipP8SlYTxGBi
sjIUDowxb21ZuIk0gTt4tCdgkj2tPvvOvGdrAaekSIL2HhU1Ysvb3EnKggPWol6h
AHJF2j7h6cmFLK91U1UbtswUPO+WQ1Yo0c4P7VvGXHSrXzXgyBEQoG6JLcIl14an
KUNRhFP0uiwTxLCgpf9RjvuOxpBjF6Z4PVYz6JMMKpvYBrC2MvDQKULw3O6mAOqr
GPTa+tRqUL1brvoedC9iixkxYySlpnRzAhcZM8xIuQc6Jkdk8eOLL8+zYAa/nX9d
RDOUEe0WXkZUChIPnF+XIrsfC/c8wAvyBU0nQBpK0TXe9mFN2m7Itd2RMmoQzQ/Q
/EryXfJvPvDpISaOSDtlPZ26OCK6Ay3o5FGtp0UCkKM8siCs8LTAUiJ/Xr/adbOR
joUgafW55x1GJWuMi4e7WPzgf0QRbVlVmr5OOGRPUghnzvV9tMzsXFFzJxQNz33m
AoHUHLewGs4tCvlaJnOIVrR2I0OwxYU9Wt+TUk7nVPOUXbXUI8KMOkY/yC/gsy6G
EtpdHgaddpZ4jFVJnW+qFxYQr2WhLRt1Ud6/bBRVjjSG0cXSM+uBa1Zm2pGDaZwi
M6jkkTWHLY2UDbZ4qy4eiC2kgJj/tYDGEsbkGKMGOWvxRtqltxQrgaJwnSar8ACx
urZeFvnIoz3qCLsLefQUjckgVpbHOmPI8WGruluJEgAyVSEKw4nYy47cEKp1N3Kd
h7CWy8+B3CplIMFjEizBjk2bsgFgGbsrpYqKo7oW7KaqJS8yePRmy8xLeSxFgsk7
NCxTnSqrurA0+StpRucgMQIasmaNE7wHymLFJ+ODk5/F0islJAfLo8HdhR24frzc
ReDAIWdippVn4FTihNGv1gdXBGdl+j4XFhDLo8uTlhKQQvdKysVDOJAcFPNZzcUy
1bYJKKrQE0NX8DnmAaxGrxSBqARkGNIk3etJ982PpgsynlMJOYFaJGvPBSEPi/Ya
aVDEnCr/UavMZoz9ANydEyDPpcpbaynqjVTf6HcgL8YqzE62os7viWvFof6zKktj
b2a9EfVKzbrK5EPtBN2gfiZbzXuU0ve9U1fdPfy+mQIqRLrXu2H/n0KI9W6wr1Sn
7yLxQTsTS+IT94B4XgRYgOzS5WgY4+U1VPgjNzmmRPbZrSSUas0Y24I8gbSm8n6f
3GhZayBVM/qd6Ep/IQA46zEKxvF/+gs4bG3/M3HNW+FO8ze9yn9mg4/99MLQLNWd
ymaMl9Bdb49zNGZPLjxorwODidg3VBOUZHcLdlXtT49j9WcxOV8nzMPnUum/9CCR
cUsW313kSfQDYqc/OcLjiX4ycvgdOE1Srp8tRLj7Gz7bLLZMhROvBxvvM2rxk2xP
voGag8WPfwO0ZTSGLPsYvZE2jzbABjkF5PNqvCUU7MlAgZ9Mvs3d5wA2do8M4nny
VLsVU4PiX+VbJgMUEf2PhzTDzezmCkbXJtd8+1fdk+R0okruz7CZVK6q6aj4TdT9
I3o6Dsg5cprOh0XyhvziLyj2euBILSOt8bGippZ4BVT3J/yulTZHXC+q/r/naGXT
YKqU2UT5I9TKtiyvA2cn352lj7JlAJFRCWKzgZGX+7qSmR6TooTaR57WDSXEcQpJ
MFOP38TWrhafj6i/z7t0QSc5vx1IMxyMqJMpHvLiTq0+F8wIgyvD+yZJLYTmQZpd
R3F9HDa+Ob1zG17lOquHPHvAmF98xOuGuJNQ/e4mOVYOqsFdyk1shcvVt8vAssem
BC5OeW8W/ydUomnQS+cBOPRl/mWbfhPJfDq383rxQ/2vyQkSC4OLLyUaqLv9UFKb
VCessbAABclf1gncPgoBKbTNoQMJXZVksLbtew4AKc4coZarP4pgSZA7WkRccB5b
IyxJJIM1U0Y15ZS+9khQkcJ1WocRu2mN4PmEFN6tXoL/YiphtQmh/nypFAAR7QYh
fnNHy1boTiiFx2Z9jz0RlCFUxkNLM1+Pr8rfZS5MIYAXFXsho4pztz6/KcQ67u2j
kKhCmw1iHHJy2bavvhjGhBEGcUUXloFWbpFkNiEC/DTe325BHOPb6dmKrjabER2/
6E6T18kZogHo1ZPwdmLFGtpUVkyDniNwv+EwEF7D02fQSn5H4xtzxOSpPYP3klKi
AozdjjibBdGeVeUfCrkeocl1l4F7Rix35DkSak6S69NItDxgu1LjNxzoB32D9NN9
mf+mpu9vSQGBfPns8UVMn7LoVA3ZTmHZjKL1zMzjlCV7k84NoCHSzizwE3efag3q
LcVhhJSmXVGuXUlKh5ikeZfRWDS3XLI56qcktgyIoHGjUWO1KrDOyHeiC2fPOzxf
f7OACB3ZfX9LKmq+knuyggKlrXjH0fA0+y3kJ3doITsYG19bbpbKjPC7oUXnxCAh
9Bewfi3w/uhh1mog99BJKcpPCLicrtKJIUh1iLbmLOXeZHoclVOr/PX0R6Fm9qig
AbiEHIrG+X2hcAXXOwKfQ4R+m3Q/BaZpI6tyZj0r/Eu8y+TOSg5bUqxuXrPUoADh
zB02V9zsqoO/eYg2ExldSs5sWWNLBFCRnx4tdhbGuANjYU+8/EMNP2M6Dp4dcRxm
0lhj11TpCmD99sO6R7WevzY4B811HEJJjOJZbk3wu+NU3nS8DktRVbsWW28h5ENr
AIm6x+e8n64sHYpO4NFJp799rFGGIhMg38MmZdQs3BxdQW9d6SxfQyLjOiF4zYmR
ZJH4XeY+gE5ZQ9yWRa/OlmakPR2xvKIRWw0tCFsQER20aE/aehFQ5Wr+Zn6vKy8E
tq+HOLy5nx+RBWyWuRRiaybzp/bVQyRlVMIZ6TYtpLXfALusfHyzxrcWj4MdVM7D
kAwmXqZUKHJgV3PfvuO2Sy1EC8t5LjAHLqXXBU+HKpITNZZnp9ZO03SXqVX0VkK/
QnfIbKzEAm4s5ey9QpOKaCXkn8D9ZKgJMjsKoMrDluLZyK7Oua+8tKPopur0Wk8P
CkAB0IRyfZuNPnTpb749HG9RhZScH0GgcoGkyR3T6HBOqBkvvMH+7PftO7VWNSeZ
I27R6A5FDMIig8Edo0bs07xh6t4lirfygeR6LmNwoLw9LG8bny9mTj6cij7oVUc4
T5/kWhpnra10LkqEZQ5ugQGE3ZqGY+t8yd1hYh2TRrlVhOn9LTVCLcns//rtNQsO
3grPxdMXcy0qq9lefJFlrUqB8YbMjVhqeeGS3nfBZSDwyGMR4B91oA9bkDfAo1iS
MV7VF7CLLdoMX97ea0HCT2ARbgqwu038tXY0AKx18NuAtR/4ZFWCpq7ZhSbDDb1p
Z8zu3xDQthm3Otai5vFAOfPtg9KLbcpvbxzY1cD7Nq3UdpwBdJudPx2hPZPtElbu
ljIbPvj+paXwtApp3KG+xopxt7lozC2yuLH9FdRsgH3fEG/qJotD1VzjjhkfjlNe
96BeEPxzrv80TZK9mh68UWemG6u5yGkSPlaFsinWc+KMwMHDSw3dFMmYtzjk9XxJ
TVAqvOzC27Ldk6oOj2VQciJEIAs6pqiz78/479gSDNJEQzQTrM7RNLtYrW3Z8x8F
UFfOJife2YrlYPgCgq+oCk6THLdcJbCZus36k59mAUsrwOk9OexBbsWOMkxIeI+o
K3r6fHqtZUbE8H3tCiCHTdR4xaTA1GZj7E9Ozj8lauyCLt+HxQ9vW48vPIb/XsiZ
6XOAaJzZKXwGVDZS4eWbEz7O2Y77B08b9fdBQPkbYVb9qbM8y+Q4N7f+2456MCvf
ch3XWpOdJKHzTOGlmUKaO02jYe68mAYOSKhlV22dEfNCfBT623Ysu5Jc1WlrOIM9
j1rnBMpMF2xvpGe27+vnUyvvXSFncNYP2hhGXODQVbL7Qo1ORGNBPg5Zh5xIbdU2
Ki2ZaHVj59A2WAL7Jp+z+Kc9c59W+3xfVkTOUIzFP6f1Z0CNuhPHaF5txDjXyTjT
osA+FWD9kaDjN6S3rea4BoRq3qB8+bhkwFD+KnMU1mCYfyBNkH4AnArNtUsviKJF
8ITKNFlEBwSzENHNXSOe9dUngFIb+1MVnBFdgeRvA+BxvDvexsV7qFPHJekpcqLH
6VeGAxwxEoNQb6KmevGfPsqOUKOkUWJ2EIGStqKzf+CfdsHrAsw/+Ubkeh4QGniD
0s2FFuns23eUDBXBdus78nQjN04HmyQrVAvowbD0DLmes4E78cPOrGEjjbGtCcJy
0iiNCidfAudszLe4aY6gJ0AD/RVSc7siNwqZe5mTw6zfGBFCZP79XSCkoTcMYJOY
eUHqZXZ5INPhFKCsl44wtYJKvBTSjkK/K9tFgL3HYhc0YEwwSHy6OvQ2jtfLRfoT
dQL+iKc9XucTk1qjPRtqxQj3yXA8Be5oiHVvhfBxNn+zuFKACX2kDR1v8go4sI5d
PqmwMxmYMrgeGyfndYSYLWu+PE1E0Km/A9CAEvDG3dzDkXJby9E1gqpW9xR4Gr0O
DeRPxsSFHY8/fuB188oBMqfcxbZo833UGkAHzTI0iB034ro5UbPNZ3F/fXmESpdz
RXYmWuS7VmiMH9Zo9L8f6yy+ZsEU2ztDoXzI72/RqYueohS/ZLNDfwppP9SR7QnD
H7bE7BZEGt8U3YcuDfQNKIbPds0IRE0dPyJLcHfMzcXqImI9YtIk9xK9Oly4Fg+r
CRxEturVoPO9erXZ44uBoDzZzzcv/BDacLhU01SiRmjJd5sfvKWqtgpc4whJ8ZTk
3JUInZtpuXYRDP/pH8eJho1xMRVEssjKuL3BDnOoDMsiJxwuo+thirZl38BEhWue
fAIJu7CCXpxLfBEVHzl4qSs+hfPEHsuNVZf+14GLvK3pnZ3BCtwYU5ZnQZ/k2yTm
lyMFKIUWEhAx4Ms5zvMhl7Z4lYl8HKe6ovyQqhRQHGzBuELpQ/96P6M4B5U4Oqm5
y6hYsO5spY8GU1nPTQ7imKr+R25+ucRiP6jpHan4IdyTHY3wLSfTeVnwvgBHIuqw
XyAx2YEve+6jwv5H/j1oMNXzfTBkaaWrkDALnWoT7yl4iNSQjOFqaCYORhjJ7BZo
ucs3RiaYQuGprvWZ7mOb6vYneTMO/8FQ7h/RIl/Nz1+2p1eCvZbNFchJzuKsR4dP
cNWAZbTkCSXsH2wyb7I8EXDJE6E12ICwUh7r0qFczJSgGHKNANmDTZ/o7JiLvSMp
9xP3+IwYjoDk4Aat4jY/DJTvZ81zZUI1dpxN0BWX2wLOvocTESYlmd/QVv1nPEx7
YavEFC8OJ2b41hTXneL+4ZcOVoRWCroMVLVHpQAN9BP0L68nWoye2E+tr1AOCP3R
PiRNG9V6KmwP416IDlC6xvIiW+aO1j10JkFXbnSW2A4XfKg6ZomVJ5uOVHE3tzck
lXO7ZXDd85PIQplwfdfBDsv2H9WYW+x7ZHjsDM8LcPaIVmxHc+M0F9ZJOoJK7koI
E6DmmIqm/GWuoRBCD+RzWwan6P6ldYRzX2RznvIpuPORUbm2KWl4GWNf1wcqzu8e
wrNddL0WlW/q6n1fcHsouDscwbh7JmaalqrM3KBBOSeDluPZEgKUkT3Nro63E1RG
7roLodfk2IQKejyw0El0s1NfMOeZsQ2oVVPbOHFNhNd2kWAKyTFFrEuvI7wcKyv0
zdXeJs+3JCMWLvVdXtc9wUrdXHZiPFpdhElROUQLilJheMfiRPKmCGl1kis9p6AO
aWu1h3RbVVh+w2fw0MUN+08VPoFmR7NC+cgA3INlsIjn9fnQNRpepUVhm8adZ97W
BkNYFz+kwGX5Suqtld+LuCxpsFIuMAy22DjMyOVZ1pc2ByWT0hV/GHAkxkqB3TK3
jVwZv+KpqBRKqhWqAy8la+0WROH+NAdQBFv2TDBxhvibNzFBxDmed+SkLqqaxwQv
SjfmZAr8oxTgdChkNAKZzXqKZYFHzEZjROmaSDRDuo5O8DDD3KyphMtlvQVb666S
2ZSEDGFEyiNc0jHMRNBuu4pLhpQHzKmaKCl+swDuwnAw1it2SWntMaCTllydlWhS
L6gS/Us61oK3cd0art8J/YZy+L3q4v/VK5zJSzebPPJYhrlX/Nhxh3THayeBe/3H
hApAuxkodBNWeNQ74o8rHxq6t6RwMp2u+dQS2MNLfeahfuagSoYYVczrE76H7f9M
rYKsjg8UwuoiRQo2BuE1D1NV/cDorhPEOVkr0aFxVvlvtmtxlUEfpskSxMtWb6iK
eW7L3qwxIIVepkwEmDs/G/jl7tgHVdfhahzxOr9StAXanA9DSRtzgm+fnzmhFe6r
L5WhTGyYS37lAtEry5LoAbFt0C5naJy8JX+epR2K4pCF0PnlEdWqQfywf60WwzXC
ryQ1vkvxAMg9Q625UBnXiv3fcI7ItWholOfv12kL5Ej3xG8lYA3hmynH37JtxXOz
xGXxhKfb2dvIF38ru8Lakgn8GSH50SNntkV/CxExnF0rI4rMRRqXOr7RcpJsPn0X
uPs2jjESIJDe9zHUpfwd0rFMBxhoT79zH6l2flL/taF0pUx2pATPeXYvNF48VLo1
mLHhmTEDPn9l9OgpQ2iqr8p9wR+E6Ij2jryW/l2DoEbNTgPymU1lzH432nqYa5Lg
nl6Q3h3jVnGy0Z8RU0nVAtAN5Kua1IQVvUi5kw5ijf1VLYrRtjvlBBatP32zFuK1
40CJHBMsDT+DWoZXlEQBvamPEuYGIDB+zt2XZ3XUKw8+tY7sObyKB1Sz3iNr+5/k
teTh37T3CiiwUHV9DsBMCMb8P6kzVdSgo19/OBeraIVlCIxZ3AvjChyGTgN5NwZW
mSmZCL+HuwrByXTdQ9p8FkhHytHhZrAbXE6FEZ4d3+Jlpz/PKk69hIhwXRe34hJb
Xbw4Ap0M/kMbFOww8buWCZODXX11u3yVNiMxJ03sb8EwpCMKi80OPK+sZDC3pDDD
iBQuDetYC8dBToirGjjDeOozp151qdfrCrIVCnrPFPE7mtGafxTmYTv4ZwhHGzaV
Y37TBoRzMzCepvc7NlB8aWGms4xDv/IkjzNSsG8k0GnKpnS7FBBX0Zl3VzYHistM
5ZNXfQY0AH3mezFAIvapl0dFQCKiLmKZMeGw6RbIMVI/VyJccXndQtDFXk9optt8
Bn6HYv/OxznG34JlCZ7aVlOgkWMkdw5sQ1HWIHLAlPhL6ulU7yzD4lHKAKzdDnLg
9xyZ4JzYflMPyfz9VnfImMdpVkPryJoGiTUcrU7lD8YFnLvAuRUxJhk+tc+uB7Pv
Da7n+Wmm25Y/kJD2mGjseVUvRbFtez7SAXZeBKcvOKZ5s4wNL/4UxYshkuHvuH7v
S0ihf2trB9GJu3aT3je18wUu8NkkP8TZ6W+36wyHoEW79wajWWXTPOR4Q2m+u6AN
A+zSG1TU9axfONXeUUM1EjR+uNifCHyY3mdth/uLngFy3fa9fX3lTVnicibtV+Wq
MGNqCJl0vOKI7EOr3bE4e+V9pXNV6aTS37WYTASHCQ1GUjvfafxgrRti2JZ7VkKq
Pmc1fvG0Xb4tAMoaLidw+k10QgWs+a10ho37HFMZie5z0Pv+5vFrjtN0kmufC+8c
B+bqqEje99dth9ie6hDSzKNM0jF57GA2cFhk4Qr2q94EEeJna8fyaKbh8JIwUn46
U3biXCj2YMIR+4mvv7YDyqUpGzweJP5RygwMe9iU0tBX/3heln48LM39WV41g17C
GVJ/354g8R1qtz7A13b0u/Qi4koVIz8ZVCTW6/foz8Eo5Ngpo6XtjZbGlHyBzRe8
nLPHxG7oOSj7j0AI3hAgV1DsSEhez7uVi4Oqdv0t68mTGPTAP+aXyNv7Pv+33vVY
SXVzn6LUHquxHbifB8q02q/9+vpACf3N8dPMhdEQBSCaL4mkGeZACgDDfC9Nyr/q
81CfAJNraariQdIx57dInefcYjmmhtGwb2WncOlf5BwDCuWpLYyzu9vJeuNy2by1
Ss7vYBqyk/g+T4lCl1g6pG4W5Ml3FUzi8VhHRXXOMmmboTQ8LMxxj4nI9a896o8+
EtNOrv7meq6FgLlWpQlbpFpR/Wj3SEREfQqADdgBAOE1CvgOAK36CfgKrQC0brPD
ZR0yefBMVG2qckSYEBNG/2e2UYourQBV7/NurqdK4Z0MK/Ru2VqSWCc1o11aYbWH
XudGOXboacMJzNawyBlnqJPSog1jNSMKz1OTGXrIOvXLD2J5CR6bSZrnEdQDQ3NZ
rGlpwwxnu2AZigajQjSe67sXXZT9tI8dAbvY/4NtGFNKpBSRkRmA8uEM6jMxdp3z
9nnODhgeX3JcrYocfSDr5aebSbHmPAXDm6s9H7e+9ehcTf1wsGfE6ymfqqS/4JvT
qkRUKDlAiLF0nCcabcCQXFxn86EEXBgKUirblrMet0gArRQbALtVgq+JQiBLt7jR
8JW4tc/D/GU37l18xtve8HDUQ3LG0chptaTfLwZkm4ZWqYAAL1axsV47te7rUEKA
F+u9YhGnewhWzSwHvMgWXXjUZkLX9c0RV4vF1mRgqt/Mbdu+GrXD5tZ6mfW+q+9n
K0TkwwmJN0pgMifsHGsTZT+Jz1vqvEz1uL05pIhHjJhb8kNWTuIkfMlN01+lttjI
hndZ5gbA1vwJQnQ9XBIilqD47uGCufl2RvQIX7ZqrQWMbTIyBhx2GYUm5CBLJYVq
HkeVme2j6LTjb9eKQwZl+gHl6NMLF89R08R7veoiQ9LPuS959/2pSI6me35weXg9
t38/JddBr7EfJ+MMws53F9hdN/5gXFcq46jxfcOIn//LHliTsWXFpekeHAEniS2Q
cOR4G5VHgEEHXZJZgWmFoXgUCf5dXtrVNcYrxT+wN0LuqQU6u/6O6brgDKSdV6Nj
lwEpco/fgJjKIqOrDTLYP03S50dGcHCv9+R2dFLI15FGILBnlq1IeYirACpLISrf
MhhuDsHKvg8cdDA6rjJfaoTsyC2kYgPw4+UJG0sQU97l1vctG0qRTEBoAiUFLS/a
NfL3KXxGHt3wtX6EOUHRajVpJvi7URdh5ZXYhPmBnMbQxQUR42Vaol4+xpUJ+ziV
ATVi8kBRCvbCuxVBW8l3tT2enUQiQEx4C4sDGA4nJICzEVwNKP4az/OXpIhiyIWK
vzdlRZbgas5LdfmxahXN58eMqCEK6M7IhFN7wO6w8uTrhl1r94LtKhuY5xhpmM91
kD3GtgSVUMX4Xuuu3yVsMpQPZ8EF4qdCuXsu8eRSiC9/VrRcmbk26RKGKU2ImLth
EMie3ofzU4TgRbWupm/KVckQ/uijEMRA4IIpocdpg9d8Qv0RgmF+21kA4UJjGo3c
E+Id+cxIxJkw/HkSJbhANhsWbA/mDoMmAohosAKKhC1XmjbF6lsWz6jX6eQwmfpi
4q17zT9n4rj8wRDP3hcbwA/1k1DthSvf674CeJGBhaheTH8AesHBHRsWbeXBvgfo
OveW8ivdV8YCZIp5tyCgpsIbeYKxwT4fWJVY0f4u7HVW6yScxwTQkgkTEcCZkejQ
p1QNuHuGnZYL451luTfLbBQ8Ewxn32JKvMbg4weOOLhEMSm998Atj80FFfGi4Blz
I3OQut4xSn1VBOi4qPnNd51MV5Td6PKdtq5xO6YN3ok9STeSM5Gv0rNO3zMumjOx
5UKp/Br+k7zi9LKb64541yQMhmiBAAeYl82yUQUQlw8auny32g8LTqz//9KZzdId
4voCfHPGyM0GK54m2IbRNENnC5jyxoJj+UJmIGjElb+r0rBJNhcpnzHF4XMgriz1
HRzekoypiMdLfF0ccWMDhCt+YXqaPZ7NIfecQJDJKyZDFDFXAMilIAWgpMZYUs9V
j08PeDxlwhVLUQb5GElPwp2/bsQyMoaht24zs64NlhE27gcaFDtWQ/X5lNiVbiXj
G+i+DUlhNtCsKOgNltSX/9BnQIwCC318x2G9RN/H8DxE8bcAg4sxRbR9PxG8yMa4
UULOjwMOOex8HY9BihhaZt3hMUF8sIcastkCEhgcYp5GB4rqbgiTRJ/SMan7NMK/
Ice1cSUlIRcH6LmWm+M5yyy+Yi0DHgsk+65I23wS179jNiGX+vE1NUfpkWY+7Za6
dtpHWy36KBXmxMo9hkhTXHlb5dgBMG3/tL7Us494cT2blr7QUxcgHEWC1gN3gp+r
LntRQmUrkITygmXeR9OhlPPCtPlaGs8JA9NwbpNb6XbxyLnzoi0v9Neh/z7biX7K
I4+EQ6BYGmKPYIQRFRyOB8VipK3zn2htOV85jQv04EnEdaBxx+LC4jLZKX8t+g59
OjwU+O8PGfzwj90/CNkRHeHhxaIxLYCK33fa4nkPWPQI5slKR4l7pySPgpDh/s+S
pC9x5YHz0R5DH6Sv5Sbvm70r1SJeq4R9xOJpbnK85CwO5d22aoU6l5hsLDeeYT8C
2FzvyKqlD9V0a+q3dmWLlgLxFeVietaFxbxZesW3MSQcDeAiwGtI6bQmupnRifnG
piDJoOw5RPwtPub7Fl7xKugwWfgYzJYJdKMUZj0Kwl9VwlmB462kjamE0OcIqqDz
sWt5En1cIKAk6NGIffQj+B7jXG90etL7D1S/HlaDoIqBv+gfPAVnT1nEsTZUEyfP
FpZN2G/EwKvDpp6qkyRYbJ8aB730wDo0WGBYz1e/lOFxEiJc0KKosjaWYYOMFlNT
kbLiIsblZuoAzdQ+cgW9yh67cRMlpW9aOW3t8i5KaqgQIcOI//YwjvgbdaJQmbGQ
DAe76WduxHOzAdufI+5MnRZ+IbFAAxSAhiJtOsBxmzmkekM0rpyn4dMhA+bblT80
fskfz7jv5i71Vk31UR0qCos+ECvOg51Ou3ZEIQSrHK+kvYE4U8MCXkxfnNErhHY4
Q3oJV52dlVuvl+SM2L7YPs1fnugSfBYp+mM1nmAUMUnjCMeO5E1HKtQmgTW1KIjf
2+Gfiy4suaVzCDM8P+eFqRrnp8nYGj2l5YxEe9Y+vBD0GDkQGU0rdeCO3V62BV6o
GdLTQcOqw2YLu9SUFrxPdFgDOCr+hdzTjyVdcJJ7cwN9XFyQtwhtNdz/bEHDoyn+
wHVPvM0waZZZo740fiNvVN2YgGxGCdl9LqGEkoMg8RBKIonNoLdDdtXLFf9N7ZPN
a+0h72Gc++QYtOkJJb0WK6Mg712AeRtcTFzTbUmI5+WzznFvw9q97MVCmVfPv9+U
dXRC2+UHl+YDbXjX0kZ8aLobKLYl2eYEH1FuE8o0ZNf1XmNPmpZQ9E/J+rX8Isjx
K9kmcMe4yPBAl/48kKkhOdy03gNG6Ea8tztPDk6oFxY4HB0v32J61qln8qRvPSxw
ED9esrYC3B3u7RJ5VRxUhguPOJ6OlJjsjRd/8BRtZiiTNcyqUyLBGdStjRTps1ke
cspYRmXd1qGC4YnLTcoEICCPm+G0/GD2oNrw5Ie4lZ2agSdMFA1vn6peIp3CBYBL
YHroEckrHX5aeajuofBHJdgfmy0/ZQ6+PEKUZMoBwc+R0/JuMd11H/3cCwD8yvUn
kwIXqmwGLfrMd15N4Vwf30FodpM00SUOD0MHKbvwfskAsLguvOFlpSgvzInSHPNa
jEO+e1LV1i/Qxl2idPe4B5VIWcGpLfq1rvBcakgGlMBECpDI094oSi30VnCefFsI
8wjExLwnzdR6Isl5DHXs13Epiqy8TitXFKhBZOqrWlwAD+Y8q/NW04VfRBqg9nP0
bJh1IFZnxTPzModK0Z0kxBsJ5c7EC5Mo3uzrGDC8IzleS/O69ak+M9o2R7iAyExU
T6n+4yFH70QaY5VKQd7LpHGxyXArvrOTP8L8xAJjfmiDtrGrrgQXL0kR5SoI/I6p
H47H293EkiAJlBnv9BO6Bar3921tKatNqFhQKaR9BgN1NlJ0i2eSNBym+cpMJTeG
zMMohe3RExFG2OGVVt1A5/JdgdWfl3h1Tj7WAGa67cSKjWwberOwTfq81q1czRYD
YtNuEIX09ps63EIZLwwtAIdQTnZBnbi/WgVcVRUZIXPG1NgzV6gCC8HWun1lC1uI
N8zHnCzrVZirWaKcCKO8ZzUF4Ev88ijQo1WWazps6UMAoOEyEu8NEligt2caT1X2
bWSy/+1CKSyBNftUvMhSB69QviqEmw1KkBKubPa80EUgPMd1Z6S5FRKmAWxui0Ph
mk7R+mNbFSu2FZrnglob+NyPU8iSWTBmVBhtR8eaGizFebSMqFCin5dXR/S6Bg7B
1Wer2y20ZvA4dZgWI+CfL3Bc2//1WQOjmfQ0NqdVDV6K/U8ByFzdgo8ERW3xi/98
Ea4oN5nO1fOQhc0/HLYxZ1Nv+ISP2TEv7ZcosvLn6pvyf39M82BF29IfbraK4zNP
ZodTK5+nPSE9fmhF4MnWP5exko8HCcIv6kYTVv72V74NpP4HBnfKzI2QCM4JHNEW
cdep2cIcF3FQB/zxgT3rv8zs0FuAULXl9qoTCyWb6hPCDJZ1t26h9zNalXdlI+wz
zJvUhZonbeo/wDsYZQE9GFbZ6BeP7/k05djlpGsRU7Ur88IzbO+6yep24D7iv7qL
oWlAVxtBcYho/3yyfqj+612w58CLfn4in7/3c3y7YNGdBvTf//GraMSu1sKGmR7+
3XQUcW66zgjlXNEDxvzabto2t7AMRCZmBy6dU7cHWwWOeFzU4UZ07tfCzHr9qPcr
PMstVPu+lLP6qRAi8MbwTknmQaVXNQfXA24e74CZOkLdFOhr3alI9N8yT2HPgFDF
lYukS9y+T/XuMe+Uy0t9P+OgOQq1W9B6nOc0wTYPmhMkaqstdcO87yFgL4sJof6l
hB50HZZ0IJuzOvZ00rju/D4ZhpXHwDekAHLz5ade25XryptuPGaGu/ekbSOMCeRv
oEvMfkbQZCOffvwVsT30QFqtPIWwmLGM3LahC4gNPHVBvx24YpnJM3Od2DZi5LtV
7BHEwXkvERAS23iRdkNJnjbPxd9EtvhPYEEspWArw61riwrpqUmbfCux7r9YDpTB
u5n5q4tD8fYZkW73LLzMWYbLBx0Pfr8RIqy+5gkmcJcrPnCaGK88wHfcsM1HnwI2
QwL1JxJZG5mrCmP2EIj/hRxMZUj6vE/e0bu5WK8KmkXehiok3Mo5lcCHbeVnWmaH
ibkiLENvzpsm6RAS4J5rwtxgi9Az57WtCH03QjkwebuzOxWh9PgOOw03ZCmqYx4z
GUfwNDRnKDSg+8gwg/LUVFO9jDqU33k6S6h+hhlT9zURlk5iXR2JXO50OgFqA+WZ
ApqzszZFm61mDGkiOrlBYpJYpS+boDNExptuj3vZhYM0PbLV3gvIpRwT6dma7gRH
kYU3WgF+cj4GzvDW7m6SKQdb7m4NR/1p4mR6OYdhIeLqmRnighB/PyWZXbxdjcYd
/9/yETsXLPM51tv11MM8zt+F7tTUzfKavB19H5r7916en7Pnhvq+CJQkpnZb53ZT
pUun3ZSo2bNfG0WLTk+IzjJTIQeSj0LaKRAIt5E0U3vDnRh7hWHEa7sepP7bzwxD
wqFkjSzoHrVE6f6rRRMIsXyPzh+8gY0lPb2TOsdCCWbKazJU1LAo50iqLeMZ4XTe
cCFTKvOOvA0BvbZfe/vohH2/d5b4bXVvMRjqISaoDiUyIrm3O2mJNS2IHjTfwVi6
E8+XHOW5om3jefa7/MpYyF2E55Ffv8DfvJG1tQQYDLCFMNNAB+tUJG0trk9VdPyY
ImdnnJv0I8MAMJS+n1Qbnm3UtlgN5tSSigzBM8GzAlE0Xfiv5KPQ96yNhYL58eOU
zqhuIgl/9aOFs1QoY1uS6UpmC1//qdO3oOdrDfdqE+xdUxvO1vSXKS6kV20RIDhG
xkqVaCYsm0AU9+GiFFYDDZukpcuqzNAfIPHA0thC9BDUP5kV+4ZQyIOHftif6bBV
o855CbITOi1H59JbNVLN3VS2qNNuB+BsTTe5oPqwFTvXNsZMjZYg3Ihw779DviEZ
rnFgb5Xpyii8trJA5eAjqnWgN1WEgBw8hK4sHria7YOql4AFH6GblTePWCC21jPM
c3+jwWuk8cDWovXyXirPHYbfVA3W9vv6zcoHePHhr5SCQ8RZw9QT4k0a0UYnHjRY
ONt+gSqadyv0wSPf8SIKwQ116HEL38hlJhlC7VXyGCTjIUnWZIs5gDVWFkvbTu9Z
pMS3yt72qOXHSeI9fqkPYBkEzMF7oUICA2y1G+SfhbyCQDWgmTc+bvos6pfbzGhN
j0TfDRfzft2WrXQFYZzWnLjZeRRtxw12h7ug4kk5L2xvrmLyMlCwkcU3B4oYuiDp
PWQrSyx324mOLQ0FstndJhckU4iURLfkQujk14zALnDcT3q/zsS9iHOFAokroQwz
PxQdRaywJ/d7P0Du/RQ/obH+LDfMbk3Yprh28koKBSr7C+h2Jrv+tgHQ7jfMWJHz
S0i37lLXf2BPmd7mZeuoWeYMJu+//MoEX8oDuhjVS8IRczApSLuqqOL5O1k3US04
MlnFeK8OFyq7iceUXnS3+64/YZQ7fhMqBkuj58gzKOmBYbNctGQ0lOzVG6XyVXxZ
+Pkp5mUGTq/dvgdWpOldDQ5enhdUWAcvgz/kC1IxUmw9oiHMGz4Elyu+nAdjsMpC
gmZf1SFp+BXuJ1UhUFTBYmCyrXTJj7SfN+ok6/z97cLYMd/xMQHodxb4wbCzmnok
kKC6hPhwcRIlF1FzD5tNGDVadDXumNx6DJtetKPbm2gBcPzJjzbwgk7KHgnvdCHR
nXHmDs7F18IZ4HAEvNR3FppO5MQL0z14jb44yb/soEFqpwoorla0KBPAMhOZXNqC
0BK1UKISvZ53/7dRPw5vYqIt0X77L07jsYfUaqCfLZKlgbJ5yxpwPSZqFCVqUTno
pIV5AMSibeJynBX+KzPxUgZoBF1Mt9ooWZnhPSWlx0OG82TkBHoJNoM0BvjmN18k
0gqSxxIGFZ4oBvIrvuMK+awULzwZY4B7zlFHxVFwk0a2kcTEh2c6J7cOxEmwPdv6
/DfZqgHKpt3460D3WvfPIQwdaD48sKfyNjbegZEJ+jRblfZn4wkIHFoHsOR1IyvF
0B3ORVtcHi8owQH2KRfnJeewuehSwci6DDxur6JfMGYuCr98434szPjEUl7zMwuY
Aska1pEJnZXniwThBU+WxX2rvOW+PG9+jDDWKAPduTv7nqwdODXo4Sq8cBSPMLdO
5soScfI67lkvBI7AICps9vJ7O3en1dpRiaoZxLkcAxY9dqovSKqSbC/J/yyAj8Tv
UIefd+Hp3JkWbUd6a/n9ZvYa7oXyBs2ikPt7kbBOmduYYz9d+ajeQBwPJtIzB8rJ
+QLf7J1+8a7ip5i8eoyGaAxTPW45ooi7XUhelDJclRArGiVPuZJqjA73AvEiPV+8
vELaO/29AxwcH4cqVLDUcrUiFbx6/5AmnROisg/WIkUOopfiqI7KEeDgKju4x0lL
BcFiWmCzyk92DqSQ737KCp3GKRuIA+W0tYRviSB9ClsoJfctQs0lYskCzGLIgS07
KIejFPcu7kA0mxrlCOhiOH3U5yjV5ORuC+/YizDGk3tHU6P+vTCIPd687LY+22vm
WsreEYUeIovPK3JpcOh1yz8bUXNBWoYI86nb4Yjl52vOplxsoJY3GKx+iCauHnji
41gp/S6JA010iGX28H2eHFO1+dYNnr9Gw1O76ESiOH7Y7Qfv+jxsDDu1OEa8o+NT
mMw+mOM2DfMk8Kpb/BRPFy/Uwm5XdyisK4ILwPcHaOC2+BE5OC1GfUhUF5Vhzke9
nEPnqD2rzEfnNrPhnSflp8J2M+Z5rPGOTOcTs3Oiq0GwnMUF3BMh/T544wq/IcnQ
RncC4kL93UgmlVCr+GPYu2oKcHQCk9DpAHFpQzTG8y1M+ag/9L594LvwEJ9fv4B2
G3E+UPwFPeETUgB7MQs8n89FGhJx/tQ7QZpBrx2IBqByl/rKzDPY7DF4EFXJXcDD
jQjhJKUrtsv1CT1CuED+sXc3yY9RVaX8tnYQwxVNUAT6GSmIOYfTIbIAhSK7t/Wp
KiR+e3g+/snPnaUILWvJd3Px4mrAlDBe28q3aoA/UrE1hZVwMPmXCnEVM/egJb1k
Lw/SEFwEWATW1ttsTNwzp13VO4Z/JjwCBAHiaSb6ut6cGYs7dMOck66Do4FqtHC3
vO9vg5nDG8KObUo8wUAYf5pnWRkBU0sKPPohChzANp/GKOrqQTXKUyb6p4tEYFTF
dIrk7wb/hzMfPoOsVRz322FqhDVurqvr42VysCH/j7qsGfcCtO0lKTXL5QtjnfEs
RVghSwjz1idpmYdMV9tkeH84fhkKKdde8dZvFt2unBy4EIl/1AnYxGa3RODV3Za2
NVDRQuMtAOY8lS1JTUfZQXkLudQIqx0nqoPZpg4rNJeZ+d6wmatfbMNKhsWysJqX
sDN99ZvYFB1Y7QK7covwzygj7JfFOee0GmsuRamkJNpsO3jrj3s7TEyI/pJKI9wt
uWXN+D3Oip+6lTl3lDC6BMAZiyBJUGJijpmRBOmmb1VoyPq1G650GeR+9WcWDnWV
QH2bnvi0X4ENvcezgou4Bbrj2zZ5lRIUnrEDCQXJ5QkUZ6GNyCa0sF3+tMslmuwD
HUwVpelh3Iqn9J0iypL1LApUJn1HRcPmg8btkGGs8iJhm4XxZu/uusovzp7T9CY8
iI8YFx6uY3GHuaCERM9TpbpFC4dQO3pl2v1qd35b10MlY/87kY/PrQeSAhoVrYMJ
esp2/IxWubk8Fzf1x6NK44vO3v7sSWEIBxgbL3lrUQgeUqC5JddeLW+SxkrFv4fm
fJqY7FwKWGIGCQ4VUPWCckF1BzF9vSU5AD11Qh1178patmVaGbcZsPSY1Y1VqiXk
xh+cBi2otNsb2keyXcf0Agn7/olXb+2roUJkcTLczYtzgepLpdjZJeXz+xTYlO5r
iY85A2hdFIa+r1fhF6pcPZUNjS9actFaTxrTtyndZfZK0dUvXB4xi6+PM/0cFyjC
P+aHkY9ZkpmwTtRpI4+jbzSiYSFd9H5fIBpeMzgQeR5ja/S8lALqQGtHDghS6Njh
eBJ6kJ7mqROko3J0jN/t/xQTmdXeMqiTZSfuiHEr72SHh1QNJ9ZVicHA0Qo/JHA5
p3H8fySn397w6Tnp2CnBJqznMDi808dPwHgZ9r6LgWsO3jhuCIoiVUMrnOAcTWA6
ph68DJENzgxliNg1RVQCg9z4puu1EmnYwLsQGuf7+gTb2OEIiQ3vX8NOA49kkI7u
NzzmsUhH0lQW4M+PfmRS/YNLCkPhQGWwjd4W0hI45s4oKtIjUde4asTHOlqYyeXq
Au6EWmx4bQkY8qzvuaL6Ntbng1BGNMmMIQgLcJnugoPlEsOEsOCLgLxr6Q1gPNzQ
OHGHlPaf6jocyIKHqal3fdJZOXT1Ha3riixRmASjlTPjRH2j4xAKpISSfwoXdIQo
WtHrbeclana0fdGGdSywwZBBUhh/MnSkvnvjTMlQz9WU4XASw5RuPO9vd/ZY6PC2
IZF/09BtEM1UKE4f7kQ2S23CrZ+5z3g+CkW/xJ6iRl2Nk3owWvCSJySgrjs0Cmhc
Vq62PkDdiuKAXy3J5m7sMRf6ok21n2kzqR8qjJVoXIobw00yHe7SxO0llrPuJf5W
oO5KMTL9hz/v2G3uuQ9qSg3SgzAYXWfHW+6UNIeaGdA777UX7D65faOtxb8mgpGZ
h13/e3X/EkVwWWCkBsEpDnxgZW7RuyzRR6TQPaeLJpzAzil2+easOl713A+5g9lI
/m+I4wVBTzCWgt3qZ1U09Ea+W4An1Gjw4vId/uf1g5vYJRDiyUxv+kxA+SAopetK
1M2m6NLS4s/iGGCcphPrm9FaivB1Y2dEtVsmXWnP9K3Q5ML/G0oKVQDDBqRRbPkR
P9c7hNGPRFaDpv1RLbowa2MhAHaZGI6Demgwc1s50cXJEeUX9g2VjopQ8RsGmIij
kdgxENGV8gDHhWYS6m3QG+K1c3pKwNCtxWo+ZRBXcATo7IWO7IY84b+Hpo5pR/6q
hqapFMvA4k4fQlTO3VUw9IwTCHcFDlg+dab5/4M5TvhINgBwCg3Giy8rGZPHiyvR
/KHDm0VbiMoiUXu4qDrXnfOOhTK5+4PdrKk0Rkw4wsaXuV2rtSo2avBPxwDWHJea
dC4azvXhZL776CyLU+XXzxgErlkrKHGxKgHfPE6mtSaNoZMcAgYhMiLclSqjcZaj
Hks6OnO2K3TmDpV6GZ5JipulFBPZZI8zvUvEcOBcpmKLIMro59PkOUE0FrwbfBQv
ZpH6nk5fKowHysXcdoLTGGqVccRxn2dEvt5b8aqi/QdjNMnDQgg5Cj3I0Qdwbqeq
JBtLGpIDMuo5Jq1er0kPKespaX3auOUUYfzp5mo1Nj0glbMEii3p6M8g8RHU9FiS
nDKoFjzlzBlws5XBft3pzly00RP8M+Q97W2V2G0tIG0LzEKEy2Uz6a9xSuJwXib5
6bO27BzFAoWCcUaEBvtZAJXwnbkLFTEkw3Rg0ABuet+Wf2bZ3zf4m4Gznn/wlsOT
OJMFBCGILn8Nvq1/fRNbQRr+Yw8It7pkoLN014pvdS70Y/Rl3qP+5HXH2ycgoEjO
TtCxb1lL/UpKskThe4TmjpQzHEnZDAtIEbwj+cEf5xaGtg/O/pkLd0109IgjLAzj
rkZx3jfMYtAEeREw099n/RzSocYp7MgMxd4nIWXl8eGQbInuwRyWmpoEw+KFK224
p66g+AaTB4d60hTGecQ9bmUBLeNoLX2BAboXy25mA4rakxKSfQKgKFbge7ovOvIb
hqjaY2oprbd6BNjcdv1O21ZX4EUx3bDDLeRs8aT1+wD1lsraX4SJxf6NVFZ22YYV
s8e1xxbgYnbr9RR2d6XyQUk6MTdy973UtZ/rAjPQsUs/ZbzWEvWWABTCDnhUnSUo
Li3NQ44FE9RfFZ7z32lAUhaUzi6brTnwpIJ9aK7P75qlsCMTaTLU8OLWdHDbZR/R
WpP5218c1cUYR2oDgGdxhRdQ8ewxo03qvcRrXFZMnF2x/vq4doPf8UFj5ASiMnmY
UeJK+WEdZi2RRnSxtTHi4WRLWQePGHu2aDgOPyQg4pkU59IMsb+Q4X0OZNinxdPm
XdmptfgLJbRhKogkuBDAUcnv13Ux6J1DDmiWlbKXX8QQDCh/ZfXm43eAkG6XTaXW
Ua5xIhIOu8TbXPwsr8bcTY5bkLa+IVkn1NVM2GzNP9wLA2H0fmsn49+GNNrPI1Ng
yB5OomzMcTPhqY5WWXQ0p2l/nSjg+R3J1l3T9edl48sXSK1arUVvrhQZ4kKZBl8v
poRM7cXquRrDB37A3InoUMzc4ju/PmX3OEX9MNI9fDqefadgLedmoNxJ2I/kph+G
8JL4bNYd0+SIqu1pCf7C4XLlCIvwd0GwOzRl1IeVK9LdgQ5oD18jg0rFeXyyZWtU
KV+fdoRcaxGPu7x9sCcvUuFYW4DyCSsjvNACKUDIWa5s1/EmCv8cE5Y0SsXUlHWa
X2P/DAsYesrt/e9W2w/7evhbtvsCUXva/kV8j2E2JirjC2pqU4rKZUV1IW3c+80Y
bHIdBUnSCGEoolnhgI8y2mNuZxV7sf4ubfPRPFTWO3qLv3oxuycoM8EJFI03Qf2/
PCYgG7vN3GT0fp9gOfzpD0lI9G+EbxTYJoNkpuu1FhdlbbYuZc+iPODQaF3rqW0/
NPk3pbfLUz7OnDwmTXLwsX5w+oM2MB+i61oubXv2Dt7irgUOnJUml0/wC/UxJGIP
nNoCCt0oY1B6Ol+hR/SzljFp+nxQMXu2fKGfFY5I9Zea0C2dKpQ7ZWcsfsgptDHz
vijKHAV9M6oJRWR3gEq+Dsx5P0M5qxFsnd4g056pFXaRT/gboJHf8+0gQvJydEe4
1sWu3YBKev7iLACk1v2BLWEnSPAaPatJJCQWtApxL8ecn4GoxItD6Am1ZySR9S5r
VfZeUaQNfnV+cPzTVIGt5z0V3MqoPLmx+AaGtkk/C2BKahn2+G+Gwe4EIdlxh0my
2vyNMLYoqzl1VCnkVlmfZAXANo+arK+NysLrSVNG0nLweBVkX5hrAgwfKCAVThJ6
fr1MejNju1+MLHO8p36z5M/1rdnqNCo2Zj8LNr0og0jPoPTMJBRj1rxImCy1azoc
vBUqL+q1Pd1xLNJXz0zUd5HeYSJ3fasVlIUCAJRzisIBRh3LKXjqzC5OL89V9Ic2
Ucvs1xiGElxpzq3B2ETMruVEa3DxWatMkSFnG6ggI8+DaTkyLm32MReKMWzy5gNI
igCB1bH+K8YSguqHgIqFtkPE8z8anc+TrtLUoP/xCE0Gy85T2er6kFmGCUt6KYSQ
NwyKSR0VLhdPi9vEO1AWLUB932poYqOs+NA6TFhThwgpMWpPzRPI7Nax//jTNUkR
J1DpGU3zt6QSd7oCBjXNktr5Dhcs7O/eIiRg7m+XGIAone7MqORjihT7KdHeYEZi
wHKYBXVFG75noGIMa73rKYOT1hR2y/QBzBytg8Q41jDadR8mEZniEyHai1h6+lh4
GeVaEPZOUpTTnyHzI0EiaS3B9DbNHybGlU7f7y7XU2QJUsrsXdzhFfap4NB/4Pbh
jTxaNxOeHrhLFi1toWymq1qsobUeDm+a8Vd7r/9RX7A1Z06qIQZE3u7UL/xzs6lL
kdYnyiZPDB1AYW1Mw5cPX1G6eo14qB8aLSGmaK3d5C/VmnSxd8WXU4iQnyaKuicU
1pnTZO7YIrq0djUGNie9Zj4NsyIM1u/3lC/q9b7ZWlrRzHVDbTJt2B/6CPSTV0Wr
keYPq9h6ZY8QXbmOy55lks/NTyrlKJIefJK5pcqzWRHAkEB+2EC4sSeDTKndPKu1
qWjmYGFll4vTwWqCTBXtzf3QVsSvxMKBBzx8r3xwjJoGW9WnYpfimWOpGdr0c8S7
BO2Hz4yPuXmBE6XtPVq1cQvkQr3Xmb5eBwDUqtbNVdiEpNcJ7PczPvP4jFaAua/e
DR950ixwpx9iMi601ESAR+3eRUid874UFp+o1R6U/rlyAslGigiYHRrOIndFFchO
LDaBIYjhftyheaEEzmtovTRTxma8HuabC7CkRkOiDNUvFaAv50WtwtKkWKXJX72d
3iVMdmdQ+rY4f0qk5dWhLU5M0sQrS3IpCYgDpLsoVaZiYy0Cc8J6RVwpqJjOrjZV
LTYqDUvQeoRpfaWBk8ylmdjyV9CZIjkQDp+FzzT0du6sAsc7NMhlK4K2pXsPtMIc
4eG8wyzQDz6vTFsrFdNEaZEOPKUDmkM+/75IgsOuxUMuySGGGbX23IoW2JLcDz+P
BSvD9MHYtQ+Kye8RdF3mYDMcbcK6d8Yg7J3PZE5WIR9ah5kvqRaZl2yRkf+r2BIe
ran9aSic3eJ/pYS/Lj7PVcdeeg62Yg47ZsWeIteOLHA6fD3XWS7UGjIAogd+rqvy
M0KPnV7yCgxkVmVKLfrOhZYIFD5qLbPMiizPXd+veCcUKMqgSEo5J7K/If7gJVLV
5YC+aTTkuu21iSbYdCGPMuLTrOgMC/zPHpYy+ECAOGV/T8RUH1pNLUTfGI44HxzM
jRwf7WJDTCmktKAainSt9DvvULMaM06wO5YuXbgIjmZLaVs4ZGRnVlaa3BZFC/Ru
FQGbYJvzSeesRvx+5F09KsNm779iFKOzOvO03DdDHBrBm+t23hlcpMBexU19TjKh
ec4a71zi45joE3rPdP/J39SXjDO2jq3697/JV8LuqkqEQEG9WV/05s2n3zrSqBC4
DkoyWp7bS5XitMfH8QubXuQ3/Kxk1KP1vqCUZYLlScA+xl3jE3QTRDoPbhZwpv4V
Du9Mi9ZVxVa3ZGx1L7xHyFfS1Pj/XU2ond2IMHzpQbbm32QmIdQEGMlanSDXNm4Y
feHMSYr1OKeVZtuijaVp2cYprACiN0qZCA0nE/BXZ58M1XmS/9vvSK6kl0KKbF+j
c8puIaQ4zmkM6LjqH/w8h029Svwc6xC8Kt6N0Qvyrk9F24jV6MK7gc9f39qbZe4d
5kCK05QAwdOpw+vYKoug+vyzWz2gmzTw/i5PxOvGWoC6YQ8w+2JGrvXXl5zsQZPm
pZwPtJuR1bdZfoqTcDEqeGXILYQ6k4Jb/vkmnoAUbXEXnXWlTvgrmvK8hlHWfjo6
+RalIlgZfAcHufUsqVVyxfd2Hg9lWN4hEZoCRPXycDIE/yxD4mUGjRyMMpKxQg7b
xMMJ5+5Xg873eL3cUx5EcgAnX5OGa0ckuSvhCUuwnmXdH4jl/iWz90nZJzHcjrg1
Qal7xtTLLfWmQlYPuXBuw8SzpI5W1Ilh3RZcbuWnmDz0RNS4BGX4X+p0TueNzdi6
gaarvLu8Hdnjx/Bm+ChCCj2dG8BiBGHKFUbrmuMQkrvKwNfVPzw6gcvbxMCKpD05
lS+B2wwvRdB9UFDSRWRx42C3ucZ1FslNkwPLIgnXv8VH+OsiiGLc8023vNr6EAKR
plabAEgnscrB9k8G4w1CyoVs4SA6ArxU62+k2hzv66E37KoL4omYL8bKQabVND0b
3ve6AESsrN2a2iwnqCyPQLo6CYlqwFR9fISQQ4GpCFKYI80MN56zAD0Y/jMh/scY
Qi1B8gAZfxsRcRrYxCrgIWtAvaNzrTL7xFJH0q2QqA9AYTBxwoUsslbIznYgd6Al
R37E8n0hQFuMBo+mXkLtbIGS0rEhDH/wOG+EkjxdCbibMOtWLlk817ke/4EQ3lsn
s6HYfuL++8d49W9kPdWYwfvK8tWTbQ98iMwwpXmW1FwDB3UiziuteouGQAd814/E
kPVlcqZElUtO41NCALGQrSKBen4E9ltEmhYksGttJTxL6pLrk0xgIxKQsh18He6t
8J+c6KpS1ibvSRG2dI+kMPwDJGKe56vyJhL6PkvribNwUda+A/6A0YGLegN7Equu
f6uKFfw/+yKNWWG8lV//CGtQL1xhYzTO1rBEDo/rYlOJHPcY/lE4tCihPPkfc8ft
iRoFqsi/UkBijCEiREXhT3BG1m7e/66Y4V2BbpKEbavhj/XUrnFyW0qLbjL5/unI
lbKRhTf2EfYtuMjgqpCvao0nFqT9BlToo3Qpco9zs3+wWYhtQZf+xVDnc2DGzdO0
o8HSLUXcQqajAWoQyMUwAcjeKLY4BHgcfHCM1vPNy5pQIhRkfa4S6fQuKCHoYm9k
5LJIOq2N2nCS/c+5+0XAun5bmaS9cSff0ZFDyiBBlTYcTMtaxzg6AiOKoALbm+oI
wqQLCzz/WuoIRg+6Ek+9WyAwxOP77UPbFY1+Z0GXc3WSd0d67SDSxvcxKM0VSV7t
yaOS3FOdYqBKBjXcQJeafHsDD9b8JKwEdZqMFLW2IKdSKxp4HyLBqaYD/Tk8SqfR
mLQeElBaJwr9+Gcr0L9q3UzZa1U9cy3vsWQuum/PYnrvYmPk9xxpdYlkxNY9MLUL
tpL+rWfErYg7n2n50wKprjv9bBYo8G0AcBjZfLaMl/6vuK8a9pNu0GIe6wtwWXhu
b4rcdFeh4HXsr9SnRwwES7dbUBZO5kd19UWhx2KdLeWmlhgcHvOea2z6JtrHexPf
biUYcFK8EolaBF5oZwRv6Fsr/EholVONSIMtkAHhDoWhLvrrOnPKze55FP7Ye50E
bTg415CbGBqf9BfhFZe2mL/h5eMl2dc7gpBNeP1i4+s7D4NPRjrzgM+MaXmH+2UJ
rLaXo1KEubbDcVcUZlzvCb1hXRZFJqxvqrIN63R1AIXIjQJbNeXz4B9ev5ilIYT2
irmAOQ0mNpxuKsokZxf+wTxklh965N5WA517J5zfK0AO7Nou5VXo3TljY5cYsxRo
GLwDZPOyVdexEoAV6gyf3/T9s5UvOIk4cz2dDkNs3gEAMf2oXiMRsa1ggL19Hc9P
g8TRlJ+e82i1EBZkJq1hI5I8gD0DWzGo6uR0QfBjIzccrMmEe1OBnFfjBgeIyoHz
noRVM84W2c0um1sAGZbvjvUjFcWYDv2qcTZzm6kOvXcFmgazXKtMzeOqO0q2YEA7
3AybP4quLYGA9TTSbwzKybvY1BhQ+wzsZYRZyO+Iw+Pkvr6s8+al5EsETgz9iCvz
Y5FpLL2LzzqguAPPiM0zXh2MliU0Lmhx7zDDZZGd+KTOyr17LcE8q3HGjTqr2tnC
aZOHxJxwOrwDALyXP70EMFuN5BOXJsPKRzXZ6kznR2H9oCV9/dQpYK9Yimn5WO5P
Hue4BTGYmA3UPPCF8nFHdyB0A1VCgTEJ4tV9VQ2LjJHY7xO27pq1NUbCXPqLKQ0X
JVVuGYmLXNJaLQNgVX4gyXLd16d+FCgt+nlL3deMwdgE4nyYGjOfYmz48iCC1JbH
5UqoEnviRra+xs5L6nF38shVQHlyaVuM594cPu+mn7mIND+yFtHCCN18amuqUWRi
+6CnZ+KeeC/9lgH1bO1Laf8JqNBYLmR83EoiWc5FU5uoqx2pRnt3W71qzqv90xyH
pehn3G9XSqnqXqAznGeA99ia3SFcbJavCr2QRdRUpepymH6zfvs7djQn2RLN2Yv1
w14H1yBdkajJ57BND0v87315d2AxpcEw5kuBoDFRnrNjUqZd9woGTsZlyi30Yale
f3tbq2vimquDySHMKMtMMy6zMmYpiPWPvV59Frh1Wysl+DVRQl0eueRI7sYk0Y3K
wCUJ28ajGIHdOqFzDucQ0cmOMlmurf7sFFpXDjX8QLW/I5JhxSMu1wCj2+dgdend
/WFYXCsXgGnTSO/cbkVPbhqMK/oKYx2Iq1/zrGc4eTiHq3VI5cspwpml71U6uggj
+xfPOtpixIH8Xc6dQFsARyonIBfpVaRsXzZ51ml7OSsDMHKjcqkJjQn0cH4BrXPA
RyFoty8nesDHCAb3ANNZrZPnxw6pLaDfbwaQwmkNEGTwtJNNkR4j4f0eiMnOR0i3
3G1zeb6f6bWB7qFyL6wrI8J9H1d0ozZ+DT2nFAjyf/TCEiGc7Hi5ZslKjrPYzkDM
oIDmMOUcTYUQ/2/2Z74p0Y4yU6gMUEyQE1JzaoiGeHu88kNs1fVk7NJ6hr3kWSXl
4E9dasdQpcJdbD0nwa+yYVsut2YDlEB2btP2TQ3wN/T/AY1r9j//x7PSRWnHiwm7
xrpg5Vy8TgdVGdgnJYdR5+o+lY+nIhGkFirTjSb+TQkZc0O2IC7Q6TBGe/UIQSZe
yWj50qkCFz3We4wy63fla8mZdOJecE1V8HzmOOotRqLlKxCal3Ux2FUFYoMpLfhT
fipaj2KABI+kcvLXnMtVrFUirkC7dOGJF54l4yVuYA6bBnsagm0rzsSJOAN7HTWE
TLrvRehQbiWD5ZTmw8lYF+3VALplbLOeOwJXC+atSPK04Zn1G9udi9lSo3GY0slW
JaDp7jKIuBl+0nqOZh0RQyopBzPCEC8Qq2ulbBJQdwOJM/u28+RCDRzZ7d6/7asj
3fBJNu5Xg2+sSE13yuZVRN38Z0Tlpac9iipCUaNvsNCFEOj5DEYV2+leW+CFhAAz
1txVnBVXhXcw1r7Z6NXKZca0qZnpL0JKXZawFdrL1kUJQWZWI1Q7ImDH1v3fVg3S
5zkQ1N9zbH2Fhvix+Ui6Ap1GNhV3jOOAdvLK2U6yKKGkKVifak4/otKa9IxAcydR
JzLPgGW4jn5Ym1bBnipf1olSrz0pPazfD+6ZAKMqLZFEmtPb9ghWPxOtVfBIqaGX
spdEXM6kI6ObX9dBYDNqrJ9ZqtB248Trtiq1yTZ2S9t/kwl1skPlIqxP+tZNQ6Gf
SVDeKmBH/zVpHMgqCNZxnkRanBqNoZlOprBuVpw1cULUJiOoiIqBIeFbjkvAvGXh
3PqWBcI8Y1zZmw8/IR8Al6m852r0FUXsZbIWl7NeA6h9tyyzaq6/4FjGZsU9iRiw
bu/vVTbmwumakvoV76D0iQY6I9A7WqHiE66+e35QwFGI1zmBuVjZIglioo7to+Tc
bZ9TXAscrl5M3gf2T32oV+/LAprkltDWoI6ysqIheiI0EsG6Nb3eWwuxmpdH8et4
f2mDVgTTDIKfdrsaHvgE5u7Cm/7KURWB0DYtB+DhIAvR+Dju0FDuxP7wz4TRLn6Z
J/EUQiilYHRO3a6qqQwLvr6Id4oNBLgS/v3zgybHdakUJWroN1OsqTBjQ6snQ0T7
LaKT346Upiivg/79+8Zc4R5q101k8GQa/5u0vElnA54loysMoSrSjybSRBnW/HlI
lpONaOoausBCVwerqc6/wulh1h3w6OKKYmuwlIyLbJCdFjj56s9dSPLmH19ZnjNg
Y1pMIiEYIH33ja2wf3waAR0FGZ0hBjLcoJKak1vLYPa3NmAEoA9Q+SV2VO9C8ehA
r0ljtl3l7+PWriuZbpbLRMfdj/NwLg75P1QmjTYTbyuxc/nZH6p96o0+QjSy8x99
4g7VaA70RtJABSmXUzQaPc3dYLWzK1/Dr+iQVbmWUcKR4cJMedX4IW9RPu9q7uW2
jOYgLPEvroludMCDF103RTrW192/6Bj04l7AmCNu2FL3dGcZH+v72aN7OVbyC9f9
AOPYuimX6AHdYy7WTsLzZDQfrx1Sn98TQwXc5/rg8gccPklIctZgJDr5zgR6HO5h
UOdzkKB5Plf+V/zCShJzg0HooppeXmA7MNf6zf8cCb6Jn2f0Iyud3qzdVCQ9BEG5
6+v/LS7z9W0eifa6NhOPDEpViz5ARIWaeJdFB5WtaHcsjzJKB7RLf89OQHO9+ehV
lLQk2l8H/ovX/8l/j57sqe5s54N5ZbRn8upeRPmqbxCaSaeBWxqbcw7/5WAPOPhF
y7oh6JG5qlBpIrf6+YjI+keiknwHM/DevGBCQ6pwg7vi6DTXPR3nIVdZqtxOqN7g
7awOo6j/sNyeo7rUer3X2MwzeJe98C4d2kE/LJwjWACBeVJzyaq5gHnS5uTzr+Yd
pBtoTltYVUz4aK+MqYyz9LGu6MsmvCIr1TGYoXE6oKI3jFLojEIZCI9Cm1q+obpI
98Wz2+Lou6jYCtz0myWo/dbXeuTUOotAZRasNBhLXK+0b/kHjQ5pAGKtjj8oEfbG
wt2F89dBD20xm9i72KKy3y+bT6M1AsQGiVcAj26RksJQFl5SX7P3LqCQ1fzgSttB
WUD9Gcux5yBsqxvUVLHxnOzC9E/awc2QZwSdPWpHsCUo+O3RZi0gAcAY1qhQU5f1
xzho3e4hGme1xo3E/GS5cmoogv665h02r/Hi3h/qPmD3M9oDQJjf5tgdLasfQTdm
IZxXnIgk2cfGBkAjTrW5vXufNwVUvAhW5ye/cqVfUpX5NvDnEDLMlQlsqep0u52B
bk7hbHT9EsMDKj5083/MUz3rFAaMfRiQzPeuOdO7byNuglX1M+nuYcTJ357XfB+A
mImc5FmyHLU+jaq0iiu4ssBTREnfn+xyVm+c+0zstK0HfvGmocVrQueRyEb3zvDU
rxjxRHaLLHms7wDr4xEvy+CA/6OHlBFXlcV5E1TbbcKGdMw2+Q0QHMmWTm9fEcbo
RAXP75zuhFS2WfloPCjl5dOJMvnbilL0UF930SMhFcEVNOD3ENcA6vn2CF0TGC+J
MhEiZNaxAYV2igeU7H+RPZqAFxRUk8aRh5HoIDWJKIRNW3yttgikSdIAqE7I4hZV
bvQI2Cz1uh8jw2oRdU5dYNQK3zT8goPF+8WXx8xCoIVQrWS59u5lq4Z4lInLpQ3q
k1rsippGUW7XKiJ63nw8a6BOOiE2CzY0XRZUV82OIj76X63RtNAL2qxwSHx+8j1c
t40UGWv79lBlqQ2h+rV6JoNv7i4WG8VSBnPw30m7SVPXiT36EdMUX3QpqqaXJuln
pIR9SgUDFwpGxKFhVWGtA5th1m0//G4u3fMHN+GjjN3m/4vh08alp/BBi5HY7qEm
9jlHuFdw6ZUiM7+y+266z+cfKQmVyWY4lUHeIcaEjiqZWqoG3A70+PqaCium1l7G
AIV7p5a2cNrzEB+SOIjmsIlDAkrUYB1vtzXZEYx0f6qPRQh/zJTsT3G1DDTCL8+Z
Is3eOGNIBv7Ly905KN4JxHD6e+tN9CA40+pfXiU7sT2rDRfP9dGYqDA3a9CCClNw
NKH7anbMGVEiIC7fQYhEH8QhdNG7AHU6EjrxFetzhDDJ6sH/qaW/+U1cOmQYavs/
2WFJ/Y3DdIsANrDI6ZUjzurOkf/BLqsJSsrMSqu7N5ojenWBa4/368OnqzSVGNYj
vUEdTGIeYhMUPl55Q4pv3rjN4LEsN/1WN7rjxR/k+emjOOBO/gksqrKTAT3N4FDp
mdGWEyVHmzFwxBGY0yToiwnlIqNrJwQ/DwrCsFekeKTW0bTqI+etJiX1AvZT0PM8
0UmSv+OmXGWGrtQ8nmq92T+m37CmGPOJYF6yMfqPPgCUzcRDTs7fuFDwEPJV3Pwq
bMkX7QjvvtNl2Jp/AgnGD6TStRKNQm2V9qI5kVwfayRuIBsxnTHR04gR42MwMxwi
wC7JMrT0GOeVtbpt1FfVtyFlUzDWu+RyZ2crNbt3qyFmoO1DrKSQkadfBKuSQF1K
QEFA5/ZhdaX99H0YcEz497ubcZB/XRDDrNGZQ7vjMEUQ3985+Q9ZwanFfQYdtqh3
nIru4T7yKGpRFUsHnUjR0L3McqMdZpWiDkmPaHm00ZjfqYnOdL6JIxdCgd8gSYgk
mjYzVibfz7UHW/n6vO9H5STQsbZ12AeyRgy4YXpaRR+/HDi0gt02R8iTooqJf9Tp
ym2gZzdv9T8NLx1r8NpRuYEpgwGZbryVWESpM3eThd4ALJZdTh4EcBcXthWYFGZN
Wpp+8JjXWgjlbEucCM69EWZrFkoEP+OXKo5i5x9LTdVZ4sucG1ML+/QbIc8FaNw/
RicHLUaiPlg1T4F65rFbnChHwBaxq+ryOyTToQlmdtgK7e0Za5FKHz+bSnR6QsbT
YOGy/6IIWiaqLI+hYVsuUGrtbFOU7v442JNYtS6pAeoIqFdLUWVPFsCAVDvqYDWu
GsPZlFum9A8VXdFxoKVVHzSv775xbYQyk0Mmd5uyCY8FArQcKjJw3eO2oMeFAR0w
o6hAK+04mv6pfrnqpTofA0nJ91F8b7dODgwEsgEZMTucO9g1kTBfvIPQXkV85D9c
Zs1PP7JubvJ9UWqoE4AECqWav/y4h6TvUn/8CPu6ekn1We0JInf1zioWHDuzq++j
SDrq4Th3PPIDNSGUOgun+rOt6LmSj/IoUIVVoYh+jggqNkjcT1lQ8j5qbpzCgofO
Sb52TK9AQ+IY4I4yeGtGdP0cBG0KZRPD+sxW86LNWY+HThAIO9K2/FmcRQ3bmyxX
bVsUoNxDlHqDp6AXP0HrkAbwZin+JwvzdcaHm6a//6MuTmqTlEgsKJ4jgMaA6EA3
sz61s4aCa/xvQOY1sT/bXVWkBxBwcZXo/Xjpy5KiGFh+YDWYumcYUsYnlHe7PXof
iX0/XFFGICyXBMo/ZODYqr+7qrl3QH4ntiRpR11unF99QE8w+TkI92oLRq561GEe
6IQUrGz3TBKbwp8uR0Q/L5xBPu6u5zo7U6OFILUoZuY3vGQ5D3H1K2TQYUdm89Nw
LV5C42hLMp27NjwxoxA2rghQMwzV/Ev+Jph5N/FFDkjn83PHYB1LDv8fq1s9tNcy
xP38E2kzvmWA1FgLmQIvX/9tNjf6fLhzBnPrBioTEv/ogAmArcmy44K8fd9WThkW
xcvnnOs32aeC0YzF732a2YnQ8UzCriNTM9u4vONlAJiTye0hXN+4zkBoShNjW5Vn
lCGkJakn420vGXIVU46VI+spQ8WQI7vhH7qOG28YlUhHxyv1T1wRRcYFWVeBPNbC
MV0CroypfCWYQT34AfREiw6Oav9rOesXdhO8CcPs4Jxf7aa6LMo3LZ/2wTRaNn/8
25vaEA8PcsoscH3WZtkf7Jbld+yKej0H7XZmqWA6PqSInkB0p6hNwihqYBRDwdwO
DWYWDE1U9gfFLZRAjmWYGbljhZUE9Alfod2ZXhIYK9XZVAEjJ9ncb86gBVHpLQTx
s/a/qB5KVI9CbAv1aV/glOd8RZ9tC81ST7Nb7qniunJOL7jEyS5i496hqC+I9/aV
23Ltda6iu8mRzEigQeqIT0P9PEmwrQMERnoFuORfW+ncMGRe01NVrj+hMK9KdkIf
BIFPRvh9dIQfDENGkXKcP5xDobml3n8qukg2Ja2Bna64QkFikWrOWEs0M3N2DY2O
6U4KChaXX+c26MAX8qEphAt73N6kXzl1cmlxIw3DZuRGSbvaTtJwQZ9C7yH1HpQ0
ALd294WbMespg9jJ5Y4e9QEuHX4NWmVtuOFlsUMkt+XkIYyd5AdMarGIvxdk3IN3
Gs5pmnQixefQ4Cq7TAgGlHW2sN0EcYnCPJ9L5afKDlW3A4Mjle6KaiXhwvi/U+uQ
OBwO5yFlBbIZJBRbADegN+TPzOZ2hAdyKDB3+6A2eUmXBx2GCc82g/M4OhvIWANG
7K4PaPjVhiEK2+vi017sDtXuVHlucZf2OD4PcErg4o3gL6slZJcU6CFxgD930jdF
Cqv6eb3mAGCsZRJYxc3tO6lLvbig/1GlB2sblUVDQw9rn0087ExOOJKTMgTHz81e
5oVjTH+BYe/0KRM0dZKkcGXFNI+7jhcwldLWf4hpeUYIL4PG1e0xr88fmi7UKdCy
PH8TtPML93WjEoxog35MiFeJf4+fA8kb80+Qqb4jvSuSpQRhHV4RExDCL6RFU7Lm
jrb8VunlW0ysZt7/t6+uiVAGd1bUd69EzNlkrUgWaEFBJtYBQPLnrhZi779+6SvA
oXPtTwMAKzajhwbg9KdWEDoo0ASkVFzqrqaLQhC2G/NG1M8jYlLtrlZ7v8lMS18W
E/snHcov/+Kv11J/eiMilXcgbNiml69DrTihBlFaQUKLweMWxHfsgZOevyhraukM
B6Xyv6zF3LXfJ2MkstgOLE3bNuQFSg2/dnNWIie9p+gh56uGvJNdPo3l2bLE5Poq
d6v+WOutHlHm7xCIeKAixXMy7V3+4iG8k5q2umSMj7W2obRTAiI1bytoPqWAC2Mx
OtUy8uxebIXX/sTcM/ZF/vyNmFM8UQcUuijyT7x00PRBQHOMqxNqYaAFttoZzqK/
opFIPciWqmxGA3dExkxeE9s8L6LqM4T2moDklKhrFQDEFXQPWwSItek0EDMIE1fH
eg8nJnQvPJUYLULiZV/UQn4mMH6JOCPwFOAxv4MaRDMtE81Itr1qrvKg+m+gDY45
g+NwznANcxyxZXTgwlm2wMA39H8VlSwiOGQHH5nITGWIjnAO665ZUXXjPX2JK1cd
MxoKzloCIGWF/dnbx2LH1rKuZaUfQXOfrkSLMrUGjxiIzRH6eDNtPsz0ufpxWdpY
ZP4W42STP+OmFLdr8ycSwZ6SzIA9lLiKT1xaWvYThL4mxTd0UJ1loHv7kekpeZvx
B8UK+fXBPbwcj77qmwqcwU3c7qXHtMNU5GUHXNyFmQhT6h3lwNxhxMpdvqyc+oKI
2F/U2Cp22pNtGJznKA3Rmau1s+xg4PBxVFTDhEF2auBWpbxzKCuOhTsG8wMG7ioV
EIOqO7+atAY/V7nbqSJZNUpWRbG2Dr7R3GxjK+oDviQxNwMT+LX095UM7bPEFMXf
r7aGkzahvAoY0UnObKjLp8XE6/xJUI6isBXEI5ict/geHe34mLPnPeDm2ExyZ3Nd
eZbNlByG0jvN6wJFVLTB9kNFdfWWiFKOGGFXseKUCNS0RxwRGRrblk/+u6xyv/Tq
ylVTQfsTCtYydr+vOIoN5y3JMUkb9YxaGMvE7owXgVTTG+ot9DUw1QI84VdWK4rm
Yg3dyI/V0bGTYxG0rIQ9T3jKH/ay5qzDa4/JkGbrMCP6vxE1Q7FB8dOeXIP5Gwlq
PCPNhFSigheFtOAO0pez3wbTHq4w44eqgIjbRoY1Fv467YMZS9SB3KdEhwNWBWiV
jGHxPzP8JOFaw10i5CaD9cpqCtfLcAHCUL09HT/YBGTiOevBnpOvjlYYtXRS8Np1
mRbPRvCS5ng1q3WttnX3hJngkRP90f4zHlOCPsTD1tRUPuwQgWVePjzE+NGYYCZA
YK1XuAJTRIcixL5qMtNHpb/1OoqvcA1mZkH101VuqzqY9ZpqGWZYyhEgSzmSUU2E
zLbA+4FtQw9lBZja675X0ksFWd6z0v228m4Q9gNr2C37JlQst+ZMPSky8SOLIikC
FJZlJ/L/ya0m14fp/VhLFizrKf4O2ypCAqyq0LpaiPmrgzmKLE+Cm74YTDEM3v3r
5jxIMfRa4H3W9sxng+r0ORHV21WPMhRaFmxjkUlPZDxTLGSpE3arXSH6gM1YanOr
+j8SsPpQOy5N4gUUWjY3MvmfiaOslkaEKG3IRJUuNMB00kFxM2GcTAIfJ6sXxlUJ
U2Hb9ZNp+y2m8Bwloy9bokI61Knbyv2gIXm7d6UaQwzPGXQlk8b42kyneuHIDYDY
1yxi3a/gEzIL1Xm6cXTSskgwY/TuIXGAWgADTMjT2ZQwOOdwvrNnzj7x11yQ3LJl
YUkZzdqB/lsEM0Xqvp3qFBwzcWnsn77Bemy4ebSJi8Bfq0xOdwiCdKgP4NrQZTdB
YDsI29eak+I02yK3SKJsQYgcgacJ0NhC1iZZwC67HtPmnOijIYI0knzcmZYzcJ+o
YKSvGsb89ajr/iLL8wN6Ye2Bgw+zi62rymZ4sIanBuycjhx468GAtF6SNgJ2gIrG
UrXAU442pBjrf9gj8DEPTtJlpkgsf5X5mgbwKQzb5NOLkG5WBdjMgmmIcoQfNekN
os9PIES9fGvAJbB81Qa19W0jIGNlCmXOXXW/dFY05xRfpbwdNWiWtErLebnL7iH+
Sw8vNIWndGP3gxOfa9bdbm2DGml62CdvvqcnlFyxkiJ4BsjB/wNv6atl5LuB5J5p
NKFoJANqiLBg15pDPlqBgNCsA1G7dYuf9LF3sLOzBnyxqrJWQ0KabVOGc+H1b+z0
0sDWulkzNMvkk67arbX/4W87USG8hODWYsmUD2sXzzrYuaiCEDmPODVKXgi9UuUk
9fa90ki7XdPHW+zTQpRtURr4JCweDuFddJ3ukeO26mAYOlEcQGMp91jIncR4nLC5
0TQad1TtmmCGd44Qu5bfwvZZpbbWAWZg/35Ksusdud+kTUPgb/hLH08N/I9AJM6g
LCIcCgk9yY4i6pCTWfaYccylIma8Dbd6PyiFuqEaunhnTD3INr85Ms7ucnxP9SBz
qwd/7+J92M2Qh2MmL1wvJOJbMfFhPFGXz0nPcuSDje7ylbPI+T9BYLaPjWpmPJUF
/c+v+6FojDeHf36CDA87rclO9XJSO3+nwyhCCVsmsKyZn4mxRy4L7SUAobqoHW0G
QkTl2kAYKcosDZNFw0uzi7tYnECwUJS2O5dyIfNLbZrsoufrcxZSzhaodg+IP8xk
720rh25bY7UzxX91rin0j16ZkPZVNAM+briVLQxhXc/3UyGPvALm6MpeuWtp3O6V
H8TsfmdLt3LRRygcmnaO55SbUq6XeSPZb/7J/DvAjE7c1PqbXphdConmU6LTUL6z
Fl++VgjdBHupeAn5NA+sG6dK/HYzAaQbrW7YZVFWugpLX13YqTyGqUUyZfUl0Dkv
TLPx0n2UqCF2VPsY5OUyVvSRu3pqmc3QPTE71abYDdv0Go5h/vKb8NFGNMUGm7SW
djrlpNL1/6LbV4PJ+bTDE9oRZ8jxnUM51b6g+qG1g167OYM1n16zeFkro8uw9kqL
E10I1Ju+AKlpnxPoLt2HG3NZ+r2OwjMnI3ZeFF8U0YDeAe1VfdAio+Y65VdjH1RS
gFqzN19krnW012DPfcfVmWaFa27IirPvpYmRkAMnY87x+EnSMKwJ2rX568K95mHY
cGZpc7MDdYmTCHyfP+Owl1fGW4wKdTX0gXPy/HlAmIB7nvP8F8dptjlLbzLkhZC6
wtXEWAywl1BlIPo7oQP93gcAPvxqe5SHQSXFLlFJ6HA6gULRIdXzbhxNOe8yKml6
qDnBi1FFB5tN153icr/enx1FXXvQCQKL7EHD2VChuIsZDXilyXJnIPOQ0ciigwY5
U5DrcJiSVkfYaWLRm50Bic7EEgM/t3sFnRR3fPLhXPuCGrDJN8+DQmfVdjK0ziBs
dVzicpKkp5OrfvwGbEHmLiVXgUYSIXe06LA2TuXCzmNkkWUOG/wTLiGCA5abIxV5
HoU0UnBe/2AFbajp9Y/qE6a/+rQ2DHhCieLSZbgCyZxLZOGUTPDM7Jr7YhMBRfVx
jQm7aI8BWopfnrbvd0bd0qRrAtW45Q/1O5CL5bDbBEZt1zCvHm39bs+K8zZpuO0x
yi50PjvOeUeN/gtUPZ/o7jXIOCWubWKeqGhNnHdWI8VWQHfDuTlbLx3Njh+fnRKj
oSpnUMa2iy1jMGY1O9/DFFHZIXkPxNR7AtVsglSYqx+j8pOoDIVooXfrNGQHQvEC
23ZU+7pKwLW1AHhO9qY7ytzBH9iMM4U5zRG953xjQA9g7vbT/EL3otlseTyu81aF
EA3UI82TieU0TItkvItnhQ/Vr5qtvWH0fntIr3uYfoCY6PI86bJtfhNk9I/nkYHU
7UyB+5qlDHv9qXi5LWeH+1GqyUA6e/s2wibqskqu7P6nXkH8vP4cnL6q6cbILXBu
JBBV4oc+LLR4zu3bvqsnKdWCzRLKjfqwuGDBjOqXRDd8ZMDo0PPdKNsqhFsZppO1
pvdMOmazNgw9YkF4kqWg3NDitzwtPDFeV/MKynZ5EkDc2NT5WKDgPSTpkFBqVr4P
QyKPHRlsjxCKr4ohH4L5CLgCiX7Hl0aNNHOhn/99EMoPe/vh+ytQc87MmqoB1vCj
SK6OvExC+onB/Wvoj2OdRZtVJVQV2GNN9BkAgMpWiWFBL/5GJwc8AAu6LnerhGNI
Fgl01jiapuch8AyM3be2xjqyxwgXpr1tgqwHEMGBqPkxslU53w9cy4EB8XOywR0+
1SRH68ZpIcTqxxmbB7QbDur2IMSF+nRQBJGUigEWRUkXvB9bkC/QdKqeCXvHL+XK
3SxbfaoZxciIBH3tmyCSwigVryJoSTz4zcHl10TLK49OyNB+FyRNDPu4cagnxpKn
iByKUWVzabvGlrgSzAZVLWoajytP+rwFchFDT6wlXi01zWD6ItdFL2fje965BxJn
2ZZ7rUhH2Vyp7KKWaiwKXeyKSgF2mkIgm5Fwn/gKBMGbnZ1sqUVxhDS74xDQBbJZ
j64V4Z43VF59hZTI7f6KTXt8jkHfC6QkWShN6VjWkrl2osVmMZgQINL+bafuE/tt
nctrE99W+DBbEB3W6BANvSNwFCMcS3+CM8nhM5QqBFoUeI+bialKKEf9NsZmwVHQ
0jmku2r+KKjL/uuuyJu65gLpRjoCzSBwKXl9PMyb0xw8WydGN5lXN76FfAJoPkcb
0cwWkZnah2KW79OGga3Xj5AapGbVcvjC2E1qR0Xr2Fe93XiHBfDKkjTQliQr3D32
cChbRd0Na4w8rgDNoRI+rD3yJ4q2yHpEXDIJHbGDdnqycjrvAr7tcc6ehNwZRBbr
qwGv9ExEScB4bX4D6JJ6nNPH0brk4gQqvLk5uZ0lNEPu1ZvZ+82lgVHAZnYiDSxg
suXPyi4QmudN5aDm6CTpGbXto/ln4NwT6Wi5DBDzO+pjkDezbnbXcdNSybCvNbAB
hqepthZ8sREuY8qAtzS/NevUCKYC3zr7w+vZbm34ILD00qIOYju/+VbkofEdNpM4
Qht3ZI7F821t7esote7ZDe0XgqpShV9DPastbisenNUAbycZvPnmNGOummPOn8Aa
3rY+s9YunmV7+bbnFZTsMQ4BXwBmZCsOQJisBWNRAlygDo40YfzlD2Eh3eKowxAj
MaQR5V0W4U9JN4F7OwiPpEr9X87KC9UC0Ra9NlXwkpQ9zUIZ4dIFXh+OaJUlWTd2
Iu6ex4B3JNeZz6zQaViArp6PnM29b9Lfn5EXPwZokjrldMvmeoRosKDLYPdfLLlX
/cGipnQseKSGUmqYHX9myfa+RlkXsL/0TRZeX/R6qtm9lPAkGCxmjhSZ0zSmLSlZ
9K6Pu+ymcnhYrjQy1vnNsaDVFHQSMikaGAF7JWU9FpM+p1XRnItIvNCR+q7/wNS8
M9S0XaHS4/TuuVTdqFagdUuVpemkGh/NzycqIqcCkOraK1SAkvfGWxsJmeD1Wyqw
xhXVxzPIwmNX1FpfZZ8dC/8QiF3YOH5EqS/0NwmtwrW5VJLdR81j9jDef4nRJc5p
tJROgrildzIgddR35J64uS1qG32pjesMaHCyfzCforUYQxLY/03cIDmRWZeq52zV
CkZZ2ufC5mSLI5EDsHV5YlMZ+/CBpreMStTT6/m0u7gsSJ+ta9nWeM2ujqGHRw+1
sw73lIr0hkSq1KZQBQ+Agryuh/SGBrd8/CnOi6Dfnf7gZPsu07SC6fqSQVzIrbzV
tphC6ZDz4WLSeaYluAhq726xnHJJPMAujDZ+6GEEwUS6NwNkGDd6m6yL+MY5/duw
1eOmL/2qi/5pj7PT3NZiv6uuacKPTQSTFj2nfeDr5ZNmRXD4APWdcPp9+P0aE9Iz
QSULVeXnkZFPklu5qE7KwcYyiqZgnccD+nGg0xU+YGsLgpOPCNXn3wwixNOS/mJU
qAMOVmaHtHgDrm1oQbNtJ06l4ECNWncr7/nJ6mPxrkE/B5spAfnHpBWpsnrFwIVm
/15blIkRBc80EKwgl9lK0EaA2pMaH16mt5WlGvcJL3ZKJC9h21liyTakDdheDHNs
yK+9nJJ+EM+Uyyx4Kd6g/WYZPdRWwWVS7unEEYDQxIJ9JGORgbimlNlCFHXi8cjV
40BbWSFGguMC2LeNo+bWha1Xu9BELAsNWpODdOb1LsG3oV/CyDXNQ7e8BU3FrCp1
8QQlRscm3DKMJnVTb86Js8zm/K+pVIjgReYSu1bde4wVhqQ/TulDCl+UNOqwIkuL
Z9oQnQ2Q9mUAT261n187F1vxXiyUGF7jZfypy+74PSZL4mra/ome4cI33H1aHeV0
tOFGQZJaOOvdpkT4pwAaF7HkEaMjWndh6g/cO4dacuNlCrQVzcPKmD+WBcjHNDVL
XrD3mzI5yhIqOauzRjS1qqfw68q9ZqdUf3bs3vjh3UvRcUU8Frbpk0j6FFTZ3uO7
tIfgwSP1uJb2nEdi5EMkAL24sqgPLuMlXWMIPhgdaThIEaTWHHDArxuDHg/Kceo6
Q8NOyjQpyLTGGJTmXbwG/hheqnFn4F9dSU418oSFz7E15+rlfQW9xUCA9rA0gAWI
62zNTvZG1+NBv94VvRqNSW/FnL2bcpIwd2i9LEqYxHSHkp2fmlxlGqBD7rv1gZD+
iF28pdQrd9KM6FqE6B5bBdTSY5Kp5NxCaOvOW7uVB+OzXh7S2RL62S+CzCR9xLeW
ewOp2xhv82xIiqJg7aFEyvTJyQi9FKRWOTmwhg+pNA+IUFmRDc3XKflrifT/k+M9
Ce/W3/yugRv/fFdu/Odj2y/2BfukYQzQyl/C+7z7HlpozOhqCsxn66kR1+36hz+/
XvN4oBjO2g9h3Hs+VPkHNcF+dXZSitOMKQEbAIldvwFt3TBZHHtIUWa5+Sjr9hvg
A6wSWS6Z54eSWVyzuEYjaSVFXD/X3EJlq93Ec2ke1pKA8KhaINo/jsMTEuJnqJwM
X73Fx2I6NOMlrjzlXBDgMoW8y3NIdtxhrrqHMb8U3pKD9ary6VpeeDS+WtFV5tyZ
sUfwoU+qMKSRhdUhmnHNi8cZHt5lQNTzKsO+XatcFLwZp9IRtqeJTP8skX6aYoDP
qvLpbJBKxvAw29Yvji6wz+h/rkITZ93+fM//Dv38l9SyuduuWvoU3TpPcRfzTJ8p
dJx/nCJu2897ufh2yl5NfJPqNIHaq6PN1z0Kn7UPk+4g1L0esQttSWhoBQ7eJ9WR
XnfPgt6VhnuNKqGAV00x2WxCpqejl1NuYtMPGstF29E+ooTABu13K8zzYSz7Qc+6
oFshlASUoow4zffmnkvYtiOip02bwfmzcvVZTKv15DD1XqOTPR9Zz3jJOaYUSTm6
yltsB3NKUvsKMSkyfKXrj3epmmZgUj7R82OkHN4+PY878dzLHf1j0jYZ5H0EkdQb
eahhdNy6bacxQ/G0a0Y3yGYQo3Wj8J4P9jF/TVu60DiqL+FpP4wwlXt9IVFGA527
p6UlMnvurCYcAdO20Ywoi2QkxhvrEKdZTXH7EdNJraqqShXwHsXAub/GpWQ6Dun+
6/UGUI8APEKY/siZiKrvxOJLoNo3JDKXRbCCN+/YGmVySovdOPD33gXw+wxndHba
7m60TZV09VSejHKcytHNQFV2txQKt8/7+u7Fayb/548K82Wdzfe0PqiAdOuKdNbQ
lPF5XXegb/dncjz9nefugeVxiHNCj4N5KcKHvxp0NBgI3frFTQLP50s4bLP7lfTp
5Zl5PJEGYpAQfZWT6b1BndX8LfrytqMgW5yR2DN3AGFRDJOQaStrFypEIuxdqmZJ
i4LAWq6LS27/gCs1jdx6cbaSaCwD9PjK5JjooZtEHcJLtkvcoOoB8fqzNSI9jUWE
8y35HLqxxTZYrqKhg6Wg+NQGfr/nImux72vOCLcDlzKDKgG56vUoZYuhxekHbI+G
xJmHwdpD8Ih3mTmArx2hXzoFdv/dEUu3GaMel781o4APIb+vmH6g28DFn6rZTeMw
LPUJFkU4S7ns2pDnF0ddacDTICjz3otllqfZPapyZbgTNqTWJGpu+cuSXwQX7N3w
SEClqR20zss3QhBNID42/qFC/SkbPiyiHUhHNRbuHiQDpuqKQNkxZikXPXmqjaTi
bglOpG0Ss/NIoiHUwbo5BQRzX/rYs4cCiFc4BHQzQlxK17c1UoOxfl0h+fnS5uDw
TjutZ4u72qw+URdeV3NtznIIXSQHNxsF2kOZpkN+DJjoRinv537e/+tQnpmjez7G
18Sp8qg9W9EZW4KtGQ+VEOAQqh8GAwPMbZlAUw2TamNlvzmTJX4r8rVuvumpsYd4
xourbZWmMcaoa6muC4TimVRo1+8CWGkvqQKsGl275bxFQULImm+/SXD2QwBPS7oV
QwLdAxZ/QmXds/iaGu96atJBUkdObRYHHAisi6RTAtuqii0if//ygcyZ3T4Jf8ul
a31hLrLxA0PGc5EzgKrGWTXnDokC2zInKGd7MSrl/bOBZUNA6prh5A/uj7WKFbJ5
XMaZ59FiysZASbGIvFMag5Fzv+T87FySPOeQwoP4tUKmLrDydGcPp5kWolWSyo38
W7tFl8Y5RfLQzhZj/XcB545tENcrmzL98Si4MKkCe/Bo+BVYUrWLahBRpvspT3oF
iq3V7MY/WnP9LOaZSymM+8aCKnpisDcO7csESWJRQXoKLPaswsy8ybxwMv0nzpa3
PTQ1zNaYdd+aj6UoESX154L0yvGBKxXM8bkTbKEPqOY9/SMy5MIIO3h8hNjdsYf2
Wt9rdofG/aKpwljp70PeDO6LwSK/n7833B2Tt2eNsBS3tbwpy8q4PYBvBPn2/7il
Ruw/xZ+2WEoryTmSc4pedyx+mjg7OZQzYqG9WKvY+cV04F02/OeMiKGo4NioAjpG
8ARv+q1etCBfxTo3Yph4cbm1k9cTa2JsRVnz90Ki+bAGeLq6F4vx5sIDxPlXvlKF
kjC0oqLFCRC7ym9+O4cO2HEkdH217C/DRdKHNjcQZ+vK7UMAztdBnKwhr+Vio9l6
OVhFUm9skqIGC74fYSO0DBQuLD57CaGAwiN4tiTEWpS1hjLyvTcXjtWqO4m7p9+0
BXKEhHc37ng2Sn0quX03P0ytq/a7DZJLi00RpwJ/Z1CCKq606ObHSNymFkToG2Uc
XxxwDUWyLpQnv170/wI8WGiHgUfMzENS4JtojU9Pfe+NX0oVNQK/5ZqCMQamTkEz
SS06jsQN2Dz9YdgDg/gGFm2GYZvl9aIuXFtNi5YKRYNhaaJnwLCdY858jtxxWZ3E
tOo8LM7ToRhUxDK6k+8zy1pLcOx54LDRT6qLMT6VIu0gcFKMWEkukhTx8k1a3saB
86ie+GVnPxsqZXewzgubS03n0BtNIhGkIcPMO+7AkUSaAY+p/armvg3Dd+I6UVNP
PsX+wx8Pe+iyS3Q9wfWz72ajk5xHGx8k7/1bpfNbkcD0Nt8NGNaUTfa+W92Q2LEK
gerNF4UYll62Z7jGCg/NuJtMpkUIoSTeg3ByJzMRK0Dpfg7YV5PsNNjojQkJ/saN
De7MzZCAoEtBdLHUcN8+/MLeTHtS3aU/qTQaebpCxK8PFKEZdUJ0rL7dmReHu38M
CD+6PLdNsp7X0dzZV1QHlePQN9r9suSrxkCkLk+av9mkyPHJAnZVQNaxfpnl0SWp
x5tH7AhhyI55RAqdhBrLUXf928dj4jiVgG+ACCr/laKrs+JEEJYE7b7cXy1OqGIN
kMBVH40D4vMZ7pkAZFTlO7uzq0ms/Cic/+YMiriHtW6q5SPI1+kadRPi3QFR5KiP
oVcjAFrFSxMsVo5bPAqyKpXlrtikEK/rKV/bZhQjCYoUqnkjouek5eLryxxez8U8
Dy+cGfOkb2igsr+o1o+H3asTtELoyX5zxS+bTfGwJ0B8ApTYUP8WB2Z47OQEudez
w0tRZez38SASvNiRGhtNuqplRZwPCsOi6sq8sVoTN9wT5rXGaO2cwJywIsavtXav
pmKBxXyI4Sf6iXWNkmbfF7bze1D3ijbCx2BzrpsIfjtmXRZCi+7QaydqnSRDbyxs
v6L5RsYWU7biqfwR058yfSQHtfYZ4l9gDxBK9RDiRLqEnXD3aC4DPzwoAdIoTBgU
o9IuxJMnIDYL/xZ/vlOQUb+pVfnqOqflCQ65D8KXnCS4E/+CsLbNn5LkLAzEF/bP
/4x//L2Bojq6Aiek7NIYEw35Mmza8anHu3C7YY5/npUHqJXTcUmupRgfYdS2dLrU
fPehkwQF7vLY0ZTNaiMXg7B3aCPrUwxgFcNN9kKMpuOkwyeqep2bebsaWA9G6sHL
a9V/qG/bMHzqIXSco5w76OsdXvBhTkfRNR70JLV/w4CAhoJv7HCfE/XkgYQyThvt
2/Dh1RsLu/gK6f4dMNSGjHby7qq34t01jKslNcDh9mE6QCwAyS5GMEQgh83IDLdg
QhAq6couheploIY5yuahIZSNU9MIaB/ObKj1uFFzER8kQNdyiTQdPnlQo1cjFige
Ts9w8KZOV6HEbBsl0CAxggoaCRGiSdB0/nDvOvLlGlQT5dQMzUnpBWwklvMIWI/h
PbOkK1yO9LCKYJi8vx9GehQK3R6VGbbNhDPq2Z/FRY9MemRfuIvMIlpXLXcDnjMC
9gpAjylWkRy92tIMyKZ4G/Dy3tWmE57uw9XeJNN//RALo/UEjjW/pgcCPH5tumQW
qqkiK1bMZoZvS0G9EODl1lLkCM1TGwLbZaA7NdBmsFZxQkv443IhOaSjKQ3nqEZk
MGTDWLt8C9O5G92Noth4PXBH7yyMkDI1V0CJZqv410n2Y1zla21Lc+8IE0ipReaG
j5XvCpsvCl0bT85a6DMZFkOb/rLCxWg4kjJuwUx4wpr2LFZsxWyMZ/DeL2oI8m65
mfLaL5phWnpI4cYjZAEikr/31YCeK1vPZAFXOjTmuHLhN8fHQD5a8VGjLSlHUQ9o
QiRUwK9dNNYz87NSfi17nLA9uxH8pcmDdcGTHrQLpGIXfvWqYCkEaODJ0l0BGORG
s3mg4v/VFcp2Dljwq6mfHCYmHrfD/JpWyFhqzi64MM1AyKM/BctEwRQYxAmUtx6L
pnvxSCvnsm765/bQjywVZe7WnVxyW3eSJTEQ/HOjl/JU6a6g53MGnn+LRYGR3p5f
yQzPsoNuUG6QzbuIqvPnDXd3/QRw23Jtysa2hhbeKQOm6eTWHOQuqitlzdEcYrQ0
I44JK3yRNI8PI495dxwzEiHwUxe65g2dkIhaDSNoCymVDtPcwqFtkwt3R5Bdp8Bp
RDsTnkNCVpB2sRDorwaH/PydgFlusjylzYrZ22mL+xK7UAyZRh5F82tGlnXEFOy7
xLaQyXPQqO+pUGujJJLX5Qm0quUTOaTOd8EgQzfdnnEAG1sZAw4PaA5THnq0cyWX
wxg/YsymEOG6Sl1cluVim9j8/enCPEaTK4HIrfL3rGyhHv+VpgF/T4cTGvjGOI/7
RdqHRXOlAi9gNRbXNjeY/dcVpSY/58+2r2LE1JFb423N23fOxX+jrhdN3MFd+XCR
CSevPNR6ddWNLV1QAnmiBhLmKxDif+P7RgMzE4UTx4+90ieGqveHRNTx9HuCQyQ3
W/Am+a9xqicgrsBFROrmVAU6dsG1Kx3iDpSrO7Pd2jXUm86+n9rcQyaZSBEKp+iO
eZotJiHMGE3TT6+gUTHNGqRBB72hOKEJiVAUPtQJrH/CI6V/iecWhfxTJaAasrn8
QdS4mrq0/DC7AMxp762xl96eGm/ILGIFuQkoh6GhWASpdl6Qp0MPFQ36NmCgogcn
zWbkRJeFctof+wdM6zqqkNeaiMslNk30Qg/sDs4UGlAjvDkx/XTu7k+Bo1suD7ag
IiRNxeRvO7I+/jfcP2OrHbwzTnYLCpoAo1QGdq3FwKCtzKh9IspFN78oxMjWbL+b
q9SQ8BH7l86tMF/rqNBb+urvP0S45zgEr0InkmA9ajzGFGmAJxkZBlMJhfNYLKDO
XCDAv/0ltFMyIm92WkxTKzdv1JhEXemntbEj0WQT7Hz1UIwq7ikMyDHtPlGq9KZb
2ctlXxaMUUM3XJcYEBhq+ZjWLezsJsQt8QE4/DsFp/qJUTyz6KUhgqcGCtGYTeQ+
vB3sjqsupgFsEqPnuGkfgXVPG+N0bSpwELJzLtafUfeARShQi/a3qa2fK0GOqAqh
uNyUasubzF9bwXMNMPGoQO+J/bFQxYhGSA7+v/t3/NJyalAtpJW60G7QVUwB7+Ih
JeEB9QSubOoCq9W1g1lsumqKJ4eHA/xnPZbbaseF2IA/KkcT3M3tcVnKB2j/JskU
3qV/HbIzP5zrmJBucPECH5bXYhRmSkczVbowoWthdYR6KL+xyeFNlIiv9Jzfz9Z7
jnoZwuTKFseBV1cjTxJYAMgMFdmq2KPzzYX4dKcoU9CsEpvS7JjBnhn7GUFxC8qC
Ohk8JIYMcWtjoq3ANxNOBeEwcwdUzI1Flck8RIZiJ15awG68Ur/jEPgjqLAlGg8g
2XqmQovyrA08UWsSMiriTEa3eSsuzW+CG63rUQDCOrWFxszrbaipIE4XGjle86uO
c0CFT+gN8leOuK1lIMzVewI8dhPL0ty9ostgpNPE5qpyboKFEEu6+9p+BeS4NmeW
NnoWvJ09Xsm/uwgDn4/eSOuKLFHpDeyqRNji5CM26YIbZB5+GbS2Eeg23GNj/SBf
tBujqk5GA3wERW/b1E6EDIizfU8hQuSTaQpUTqlqJu2pOO+F74UX8EtjnNwP+IK+
l4KnQfOPoobjQIj2bOMvJzaj58yYjZqsEEivHeSs4WEMyEz+yGfE1L1Q/Sgdo7gQ
GOVqmCQ2MG7Vlo0KVzp9tMVAEFE6MCcagJzGFijh+K7aPockLiOrpgVJiZrygdfB
f9RMlKkEID3wb0n7UQSwX+jd4Rbf4DEV4TXO2T/90hSqL14gNs62WOyIm6NRckea
lZtxKvlR/UoD1IBxGPIClug8P1JCDKsyrwkw1MVniWowzLOKGqCRg7hBieYO02Zw
n+2kvvkESmCcwufA9aYgC6ip6yi+qAATXni+Z0VWqaxSlzvGe1/YzMjvGWn36XpK
tKSOo9+y2g7j7q0Ai8gl/rUOWsCLLT9c6mLPCQeb+xlRiFzUdgJDtQUhE1zm5OB4
yXWex6fS1rfcI/mS2W5n2bzEmeLklEkJYPUKezYmgIDIpnTXMB7iZtDZ5OMachc7
O+NhDN1eMHELOZ5La1wGWhpFMWih4PO3M2qvRW63Btkg07xOu20ZRiCNP5tCiqpj
UOQ8+A4pZpVnYeTtnC37JWiFjF1Lp3uEly9ykukIOoXhW0HlorTHiXbgHpLihBUd
yXPV7Rq765Pk/8Y4p8VeXjtwPe9mEyWskm2CpvmYKAeLJ6dxfW6+1uOXz/SEuZso
GB/notH8gzl7ow4RLi1CR1ECYC0VJvyMuDwuiBVGIsgssHOfxaEYxAjvb5A16hpo
Nlpe069cjlfUCgjkdMfC+ZtUw+oSARdbkb6JcYSEBVqdVz/07v1lk0Vq0gNze7t4
e9aRNiV0Se95Y07awOT7VbUHAVEeqdGG8IbuLlvgZ3Z1shOypLDYyyBbvoC5SL9Q
YNzwYhX+RmXZvk3m7Cw+9Mu6M21kGHKP7IwOH/JItAW/UCt/RM9bXRCT8C8aKDRY
ekCjSgcz5BnWDIOgRD+KKOF+3S5JBrAb4v8lWTP7k8tjVA+xH4L6Tr0Qz/I45tni
9thwdC/txwTz6OyA48lPXwvrRrZ/2cxG4l598szMT79j1N93y/HEoYSPPMxmdrqq
oqsHHkjieu35HHSTANpikS5gA5M3mpe+U1or6Wrtfw8hbM5LmYCK27LaZa8R9cRH
P76Z5n5aE8f5Y2Rb8XxyQNvJ2n/LCtnj0qSFR167qtknf3gjtgbRZtiEC+Qz7VyY
b0EN8sGGrDbHaLWFLZFolhf3pDpU5BiScWbMCQyuG0cwmjPKILtPFy4/Wdg8gCP/
g3R4hyNucyCz3ee5FmmCmJCBYoWlAglVy9ez96/cRuG2phx/uctHH0LOpieoDDnG
H3eYmUc3axeK18dVLLhzTK4318EQ1AE5f8w9gaLZ5D185noWE4/uwg2yKDJLDDCz
unG9WoybeBJrScoyC3BuWXrlYc05m4gMStf9PzM/xO+2yVhmEqlH+7x2OhJ3Z0bU
9GP8c3AptlFRMMnRIEcfmbqNghrSO8Dzy/MFY2gLlqW3XBzYGHNAme8iqzePd28f
lP2xFXmzwzbatjdBqkCUwkDl/w6kGA0AY7aUToA/y1LxTIp4vM+yFs0E3+JT3kZc
BRUTDOeNrDhklRFUf+ZqrdRede+snXgD03s3FSnAniizQUEQ55zOZ29PW5WS7c25
in0Di8huQQpR94DuoecDJTZU/rZsRpTWjgReMjdPwzlNg/qhuBSadjyrzWIEfCgy
8sED6qrd3ibfpIHVSZNSuMxkAyRrnOmi87ShU7+GpUDFxS/V0+SbjvRHQfDhaSy8
kZq3E/alNX0IdIv2HNnNHeI4uIe2kfE9zJNAyEUvIpowNMha2lxifqK8F9QU4s0l
r4+GRs7YUM2s10tkLKkkPAVKYbktIgddb6scSVOWoNAR+3pjcesz6X78vfm/mON1
pDnUz2P0XnNj4yu1TQMHfue4RqLPCWwIos9JDRAZQ/i//RAwxYlRyHof53bwKbqH
CBHYWPcta+4T+Wt7PS65pCQJT0ZviPFI2olOmEvWs54Vgy45HVzY7Y45fqC0S3+d
agC9x0wREehnAnh2Yg5RYQh18G8cdmL9M3CKbOfcWsq9bt9d/UW3I0I/63k11Owe
/hbqBdfDHnmfySZMTNsAGUKFntPH59iVAWkcODEu4K3UvC6/cmVgCFNLEaA/Qs3c
Swp4sDTst48sLZ/Q05LTE73p6IiMKACS7hG7ia9fJHm5VrgCb2bybUKY21EpmjUN
rxhOfbqaIT0EoaRUD07B7vnTFGFbYq/KhUo7QGp/+vNh5fzDalCsRih90le/dzPw
11jY+KFDSG1OjXfAqSKTs0Zf6A1xfcBWrTkMs8u08j+980ryWA5zgHz2sXbxUoir
atInDsTU/QLz3WezWP2ABDk6xnScIqXDfbLho0yXaPznSFtPdTOlE/XQ3T/Ca1JM
NItI5jjZv8bO0G0T0hoWW6xYqYtVHk45CnE5B6OQYDmq4FHClOyw4bNanGh2lAAa
EEGZRlzRgvgMxYziKk3EErOEC7Loue3FnOm6INmlk3WrxNGxxoN2nJBUESiqf7fE
JUNo5zy1YLVkybyl3HybmaznU3Mf2lkkPb6Ia2qtutXx0tgZupYoIlBzE2x+XAWK
2kpWG2/ksNnao01Yhg5Jn8NiodpsOpptvKTlQjJJtFZf55E821S08+E3te1JRHFe
04N7pfURVZfMv4aOiuEU7wb3JNbSzwMjkXnjKdeVAqSgKtDJwzoeDJVk9Zz4Zir/
sGJK5EQejSLhlZ98UvpEAE49MPD3ms6dh59EmpW43LHvoM1HxfvdgDiHk7ET2mEK
kDY7thcgNqaoKGvKI7X+jwPb7AatjrzfWmx6G0uDvSeo3+j94ZBE3hXo8+1/srJQ
UtaVl24zM5MLKitEQx60UDm0FYkJ+JPTUxkKLhG0IZZ/mK+gUmnr9FVrXJgkpBcL
7ztU2FdyODUMnDQ+OlNSP2W3VQlT+E/lT4dHDD28LVPzgsGxFW2kUG6TMfmsyXdf
RT3qhczrx5YXeTxCG1CiHyzzKDfkzkYuLMLpB4JkcNoEII9WiKlRTOuEOfZAzY5k
tXOxKJi0mioe/AW8sfYb+lVGKrjfeVPgQKOzTWS5Ji9ter8dcEsXgZ4SXeqdtmHc
6Ed9e6qtk4EC8IYOrOOtIu21fQFK27aCkDQbYCAABAExuKTXyHhbXW7faUwTgua5
Vj2N1A87/vn7z1oJeVC05sRz+ro3zROuwSW4BcDvlWVMx0J+Kaj8wrpFxWvyPwdC
dd/cSJJ3WjNxTQkxG/wKAQEwSkZd7UyIHm28Byp1cpi0Pb82yUypBTD88291xyL6
FgdHfOVK+sc/NMqZLRdlUfzN1QxaqVveCiBU2lEqC7kyV2iG7hrzr+h51kBWDE/E
jSIq0Z1vKBoJtY1vSwkrpKi+Pew+AuVqCZKzADRh0wYe96zfH0cCOZ1qxDJI7Fgv
SlxLrdSBS81tgk6bat19wPjpheb5LFrFXMlyO5SMOz834ROoXvELype0z1iw71eZ
RzxXaZGCQFO+bKPtQJp14OG9vw0K1DFHomc4F+yVQLrWCacR2/eC//7pEIsyx8nv
n7FZ+GuO0kFCQrsiT+yJLTNfHgzxG0kdtwni3lNzBKUafzzJwJuVF2+MCK76IFDu
EPVMpOatUoTsrhqjnyL6EdKbeHd/k+85WLMKtqTqC2FPy6+PepDsO9PCx/Kt4TYC
FwwsF19DWNNoWcsDwMNK6ig0dHEB3rgBc5H2P8fAQZa0X+vlFlBh5byFxO5xqVYr
gVNNrhoFcyprDMom5ccHlRI2JRqHMea3giU0cemfder/u3J7w8HcMWsig4+dPb5h
pzz63JEAaBq40/e7e6I0aug++27IECRxmAhn0MY8mpFez5Mzcoa5HwYdbnODyi7i
JmIwkBHVjSUFXxMYaAbrLomwdXP2hqOI7HZRatf1tSvVIPtUjbiv9pNjjDR8zkpX
63MZQdO9sOtCl3FuLSwTbtn+l7QNBQx+AzXVCilnv0E33ZdLgZxgFIhSpuQqwnOf
FX8JNDkEWcjlS4W7B+y88DR7FdrVLyjdXyshqsPUMK/1AMVx7jDb8zB05tlyUAEw
ii4xXHXi5LDXbJDqVO0HrP02hZYqYnjf57Q7ghozAbVtnzC/75K/WVLRLY5Zdya4
8V0WI3f7OYG+OAiGaf7F2LEi619tF5ZBRg+1xVO9Iqiwjem2Ltna2kfIBBwH7aAY
4dXtnKRt89wfGKszDHLouJrq+VyMomxpKnuEf+d3Tk3I95M7VrO1Lo+zyqZQFGfu
t71mEnILxfR5RLNjdu+gYRHLvAoAfnlZ4SPJSCGOTjH1YfN3Sqo8Bnjj00g1W5pD
QWPRZMKQURMcpDnrGL8VnFY3EQwD4z5CLWo61pZZ1Md0oHxT8+TQK/Va+4/nsPE6
g6wAQ5IwiCOHmTSPrw5UO0oVad/lYIpIpEWGG76hunDYCI73rdGyYRS0LZ6pP3qY
PKgym7EcA7QLirynl4gccf6SJu1yQERJ+L6ueMSDWlZsq4BnOqgwYFWyvCOqLHrx
ti/2QtDk0wAbUf+Tzd88m5zMAJrxhA4sWNNp0bhuJ667jjb8Kb0+RDGZniVmwBps
cdeX4dWnPCbRQneRTGEAWyT3gOyY17qH7+seEt0d/7dB9T2uJZwMO6LO9l+STYrg
Wi5VYBbiLbxWMagw0PaHvX2u9tdMlnBWquN5JORE/khiHJbR1gJy3PK4I5X+HDca
xQcIlQFYAE4Az4m3ygHCD4Lfz2Xbiy/79SECjN8L0511pcX4Elc1FLfAj3a4+oAT
ut5tZpeTL7HNW4AEUBf8cm1mqyiVFOkUFwgkpHO01jcwsiBD0ovxHuot8QzaWixt
mG7BB8i8uM+QY29p5jkVaCo72NUXmpa0UD/XhDmUkIFOs1iUhpA2pEDqGkA5p+Ug
JnlgFO0+jxUOhBHWTJ1c3t9GGt3tPRZ/Dn04/vx5BOui0HIRd/9IcyAFzF82FdTL
m+8B8gCoJX6Bd4hDOOrYiOWBoBZnR+EhI6OhXz+cMCAdhcpzbT0YoPpFkaQYjBWp
X0o/RkWwPJHcBkmyfnrI50pIYotTVN6lNjR1JkOMGFgIPz1ArhUZHGadJEXoF3K1
BeQx569H7jy4c/0X/y8I+l9/VWAmIoEU7BCcljseyrSBQ4qYKqzGMltrZQIvcXD7
jiqk0MZy62di7XmLMZRYU0GVCsT7hsw4PU97LymF9Jf43ZrJ2pe4f1YVMq4sLpLl
NK8Quunld2f58nXjJcdn/y+UIXYZrslGN7zG1mHqou4zJlv1JfsUJojzd2f3yrML
YS4Ce3H4yfHBhs4AnaG9w+13IXAzDrYAWVyw65P9KqeqXbTPBJW0BEGtQMiqqNss
LvdataadmXAa5xVEwja29orX5OA2g2pmjb+HTf8FgEFChRvQ1cSuyqzuEprt7msz
XLOp8Tb1Y0bxOATQei+Z3dhmYmTYsRkA/73HaDUBWfcWxRVTuYX/HZPFS2yoSF+V
ajWNa5m9osEZXa9PKjb6PkKxmDQVbXAJV6PusaDMR3aanJhg3Fti3jnnZy6wVtGZ
6KqdeffLCjKc1KwK6yMLWCLcA/MJeUtThJwsHuIHYwWe+77+XSH3Mb+8fuc3qHUB
zIo6tklFT7H5uECdnbN56CyioU9ypdNJHJWLAZYNHcKEIeX8BXVPdGfRYCobhGTb
bqbSVygVU9rkPx9A7FgqbhJSlod1mA+p1yVvux5NEcZRHjgCzTJ33/Vt0e17ldsd
O9B8YIwuoKaPvyjSDIwBAIx8INrymZ/vzl3d7DwVIHdHUlfdVYrSuhlvcWdSpG+A
k/eKUbUMjPFWA2iyq14KQDtmOPIxUgaos5T4ovNhLIbjO1dSPaYgmhfbsOUEucgk
FTvE92n2rTG/Emuw/BJY294U1W2Xg7o9ZM9JqmYQRcR4K+33FSlm7kk8ASOwOlxV
3IiloUM3hN4cQ4ROCTzjltnixGdBTwhyvddqgzX/UVclUX/dRII4ET/Ws2C+XYgg
bopoguvAXKNq9aMITLwgn0bA3TPLS+rw6W5cIhjw8lj8O3IQSfNWugoHIML/e4bD
4ofgRvh3rZPbOVpuF85PD9e747WF7rKrZiExT7/wADlFV4uErV0I+yE/aWs2drdx
Gx9FF1qJPU/HzJ+6pqygBIfaIpHLwQOHZguNQmaXCT8XpXgooRTybAHaaPlQaoUq
7bJHVGzLfZzvJZWgD2qgij3TxQPoj8GctlyanWWLDqkkWkKgdoFBCBN4IrRQtmCQ
IY7KVCObJPg7mFhfLPUZLuWnElWa5uiz5VR7bavXDziQ9fjisWQuCLDvop+H3E8t
WykCBCWWTx6a53HT8h9kqr+XgFGMtS3CTpCw7RgVylRhsvk6LDLOtWHg28rhwOZD
pOnAa/NQ7gAmHKQPdOkNefEXvajDln+G9cwuazw41d6ZKn1hN8zk1CLWRSm5Itha
tbb3rOTZG/3UH7zMqReni3A1hkt91LbBTT0G8VWwCYvHmzrNc6VMF2pIZVDqjyu2
M3PYH0/qDWBlwnvAIoqI3gdEe/HQy5NewCYajRpxLbPNz7s00UqsBfHAKcwb5buL
bLsfYX9DJdCtetNOzCZmRU+2sJm9CQFezNWRtbkBJkZaicikq7xSzeHQdump3N0W
eRml2jXUoT04IalM0wLq1sPwEf4yfVWD4OYMN66LX0wUoahNG86kC4TcqcyGaUa4
rPfzXapOhIoxFrdrEej9y9I7Jz1hDOtxQLg75nim9zBSuprSVl+SDKob88rowfG5
RnnO0Af3g7QdOniMMOZXJ1XEsC306QS5e8G46osZSsef0h+QL4aZHQI3CIpZHdzh
sHHoafZjFQZKCD/vtK/2FQwEMYKOEyF9vtlAlWvA57meHamroaVzyjNsnqBAStMq
67DK6BJJpdnYUBOfHcIljHDpEfMQxFqOmcVrRtXYjYqvAh7YyAu3bM24mBCu3B3H
Q2c0jEaZt49WhPffuA5EXc48f8WbL8Hbyq0mlud3x3rWBKPK9RSbJj+BBZf4asfy
X4BRz2mV+ZcdVIuqnZ3EE44u6/UDghUeHFelH3WiDHrYDoP/2VsQB+KtfEFPKJQw
l0n7Kz8rlxp7Lb+EqS3svDg9pRG/RCSnTNVT3bLvJFuwJfNAW7gLZKRgQR4bnunU
S1Fz1hZF/oJSc7vhN7i01IovQVeMTqn6YsrA2q2mTKYaRjDS93A3KwxKtUfHyq6k
UAOSyOSYPNfgTwKCdvuXlpkEsxznUMiVFl7xtXf1kzuQBMiyFacfuYFBCt8MCvUc
t9d4OQhfBXUH0tQqjgbVPr4u+eXT73A+Y9QwbaC/gbDcJ68LqEQpCoPIJERF4hk/
q5TwJiko67V/D5r8iP5BtWQbvFGqqEGf0GjPVAsNcV+pkfd6GDnPyUpuBpFXOT5F
QU4gcRRTfQnniYzFojQDO2/SP8JBzydpDEef5eJ1P7rjg+DFdpCiAI9J2N+5RO02
4OoeNpBzqrrvIUSw0Ml2SHlAVmllcBGE9YmmyIQ16NMp4qjyp3kflw+EBdUUg8fV
7HBNfwcgyV9ooVVXyfK83HkV/HPf64A6gZc0a1es+mymvqw9n6K1AQ/Bxt/u8VE+
f5mfzqo4q2GL2j6phEURkQnnSkrnJhA+SLaetQJ/FmCzYJTq0anRFczs2uRpG3Rs
+vxL5dYOb2UwDATyPWVNdJXXj1f0SSUnCW4sleRO9Gmv2CPr3X9qSWeAY/Jdgl6n
z88EzXpS2L4q4iB9WciU6UkQq5n3JhBIf5qk1x8VoSEGHFy1YXpg+gBpY0at0KRu
bO9cv+bcJDR8sawdddXmPYKowgbLU4Mtur9fqfU/pcatuMEpZtTzWwcX5XwRBc6F
8PQ8CyIyrbJPG7FA2m0gkm4Wx05gbAjFEXgBgoz1uhblMYhLnBCWMkCJPC5rqU9/
SZz322+D4eEhdLKzRi2DFIOYLMb32LwJPlaYT2hL6lFb3HWhXhl4rMzqm32Tz4OM
TZWVM+wqMHwEu4rHQ2tAkxfxHVDPf7FjpnR54Q3nBg5ddjUE0OaJYbdRI6IXFtMs
teyOnw8zC3lS/9GPjCfUgMDDWXMnbbn2nkTs6++akOx3zuJFSjEPmCOmDa/D+R4B
EZbNDztJyfBmrCMTOHv2u2mg6jVxf0GD0vPzSY1qFYiVK0GTHPzx1gsy5CNu2vxy
/HHsAajsGSEMDgV4pAlp8ROv7/tA1hNSU2mh48tlyyWCdcH04umcsFcAsT/hUKUn
k5pm8wzlWfoavaWSM7todNPgaQD9d4u5KSJEYbp5XZA/I3klC/4FjjT+egk0eV3k
IZ0F/lL1G2Dc4f9W0of7vEwrmtdQeBhqmotTrt7iI4Cue+b2gr5hbYaoHQCfI0Y/
5jQcr+NbHWVwfV4LtzJWkB0n+b8zv1CC+QvYday1ok5l0+5GkZnn+ngh3nnQqVgM
lgAfOrUpg3aFV1BRdqyyURmf/mmayADEy7T7NEaVJs5PGC7A294H2iFe/cIO1kTc
DZnFn/E/OSmm/YqRyRX2MTIZlncbX/V2be7dn6fcM00VpfnAt9n+Vty420dUDmev
H5iRxX3isOWJq0Sm/Ix9TukP7cQ5UKIVm6fIzsPYzvyGbZU2AqACip6slXX+8+06
6Pk7pNZT0UE//49ET+gn7Z/0oRD/D7MgPlvipofCDx3G0KqksjaTy+k6l17wrQUR
x85/v2gWShb2+n+lZzrGXisLs7OnhfErxdNvRO6TONRJRtsgxWC0sYCZeyo05f0W
6g5FRoLu2PWLKjn9PoP4Ts/+FJkxkU8fffrVnudTgQsyCCRdTh0BXjFIzQY1UB5X
5m5r2ZJu99afxKnj+mxFaxS1YsHaWw46HDpvDMf5OrUX1NLLoVRY/jIl6dZMnGtf
LLsAD05fBGo0Zb2hF647zoo+Z+UhFGH9WtdKaZ9kMZr6MVAezTYTstD2b5HQXyuB
PC6iHaJMIWSSUmuipGNO9iELLI05ChzJlHiygaHvb5RLI3sTQcekEj55MXTq+xvO
ykDbCbF7jhA+AMxM9b9TiRL40ud5vyCVBr630EtTYuSr2vGLMY7Q/WpnBHlzidoB
YHBbA0Yc8SY5zpFtRzBgznpfXWxX1tkXEx/3VUkq3uEf37okXBuIgyN0+hz3VTtx
d/pc4Ph/r/4MOmytz5T/1MzifFVsbMYhrM1b0ehkR5WmrFhNZnDiQuQRsFxFVhEz
+wxNiKHEZx2qYsvtm5mvr1QTHQ+mtSRkBHTWfhh14fpM6B6jOMpwZD3Z6M8beNgy
xfWjTwqqpFFbvrB5k0nv6pkQOtnTu1jJNVSP3dXl/pSwYD0DQ6gkq8eSG+nkxV2n
14EjydJx6GTIt//PqRAQxZfpeDD/LujU7hI6TR3qYyMrr1Og4HswC0Ybsb8/cKhi
WwwRpPTht1VOJY3QE7KR9LVmF6xO4zgwrhXqBkSmo1FH+t8Pt+Lg4Y8FWCq7n/ii
/9+PW+dg0sruM8mJ7ssybrEgo0bHPCAoL8zRmUyGGBqx9Zn9hY1tplzf3qoY5Z/G
mqgwoOVbQP5wOIB5DdY/I3gP3XGrNGU+++P2lc1A7DSDk8dJyBl6geICd3qTerm7
xNzzCevjuyGVvM9D6hSI6OpCMIC1Kb1uVZPOGmZnCCPo1hOgBAHU/GtfNPi6lwH8
H8n/ScFJxR1iB2og374M4FC0b5VUWURXaW879kduW1NSe6xxnd0A43Afo9Nxbb2A
lV+oRpEKimlpftYLrMYoa4vBA4rpiwURzDCi9BPgeeHCs/F33q3Dv2iTdPf8uBZD
Hu91nXgnSQf4/cYzklG9Qqcj/A/D2M/MuLPGiiyPoF9EkfZdMzuF0qMhsnnHtbfB
5PH96cKBcQ3ylSK4u81S1Nv8FFFm0JgeJQTb8PT4nHLIwJKOPUQoU45pP3JD7S0D
PP41277qDdqhu8WMhNRAneKjvSDdVjxuyKWkJl0rcwltOoVKlxhnAFRHVYEBVUnV
+gLJCRoVOmKg+6lI9Uwllmqi9s/sFkLgSxvKENET2IKlD4tkhx3xjnr0R8NF3O6F
bN5RmGHciJcI0kR0pEZ+qcAzVCN5plcwBvY28YF+puZv/nk3xaRTE92DhjpYAWtz
sey7W32WZ+UmpXf2iA5gZKVNULuLFa0RPRb2eaOGJnnpjFTZ1GLcAKdPFG+ZrPZ9
gUTwELSt9KVqwuaxfEUtG91fbRTzkzjrAmTM9Ud64qDbvUJj2ZhVYFVujyj/poG6
P02eQ3RC0crS6A4uT+qOZdRYDqeuG8xqxDAgZKa34zhih6VU45tMQ6Cn4LzEAIt3
4XOzVmyycr6/1OQSuIrvNGIzdFmkvYKzWBOGcmORGcr/UhFjqrn38odGen3utj0Y
ZgyN+nYxMJDht/133qKpKFytuNqh/AaxVhlG0FxBtKkV173/ccOfft39caKTtV84
CNyRpiti1jNzP/bom5WhfWGLJzlOyZ1v3UmAMNBeu0dzm/OrwFR9LNFOO2+A5CZX
QkiWYIhppe6RAUYJuQSSP5HquHuWiRZiTby9oLfXcp8d+j7yNRsSWq0cvdhme2bP
DxmypSrq0ZsiT8aQSN8W39RKrM+lNi9kzz6XO5S4yCkhnVjdbx99PYYZG5NzqXzo
pr2bZveBBKK1pOkKhqS3XxpqbTlBtvWVxBx5IRSbWhFckesJtwjq2uVurtk9a5fi
+TaizkY/WxShNxldm8EiU0/KYzLfHpydVsxJOPXOYDsIsjCV58bu9p4nvZ7Atq+L
S51sz8a4K2kZmoT7ye2T1lxF/F0AkD6fBgN5Xi+uzV47/7yVR5dusY4atRJDkQpC
D86yjEiCpToPxEJbXezocT6wd4NBw3urGzgT7rc1kchcaOxyMJyQD8JstY+vXbO8
A6HtsOXn57F5eWddnky6dOb1Bg+Tur/o3yvuC2mFpfKZmltvDC7RsS7grI7JBDnR
ZcL/wh6dbLTo4aZ2uOqz3zplMbfRx7FtNX07VlX7TXhjewPLkWfYGMdqcxu5jWw4
WipbQrsoXEZgU7stLQPG8tRKXDgiwaFYEQIt5fRipoUm2NAFyPLtGoRaQUVRfRRF
Fd24mN5kg70YlIN93auACl9UuSoFWxD/BCyU50WQvOFTjPvMHUk+WAW/bwckUfds
LCyc7nWPcsuG2UswkPwfpFbgL/jbiEESBoojqNC94GjZqmPo94IZvx3Z5bl7Uiwg
6TKqvll3D6Th+/ToDgBmr3eqETUQmK0mJIXrkPwKEHS9em8uttc8iI1kg5FYE/DS
BT01xFPTIhEInwSpQqku2wwKp3NsE7FDo46bIavcowBhJiQ7ZwOCiu5W4nFiuHlQ
VYE5pnuXLZj6HY9IwoMbqAPWchs+tnXNCbRmToMG18VDnufcUO70yxl9gg6pa5h2
H3ZJX6dIDFnUXxJ+IwCI9mSvhps9eEHohBuTfePI91+quiTHbJRxSk6VfwFLr9hg
ojVIvTeoLBpTbWWdG0KvuayU6RxEIaINHgD/W4McrMVTo1aCJBxiLw4paxD2HqEm
8QKAv5Ps6LR/6VQeSZy8v9r+4E5F7VH9kG7pHcyAP3umOb3b4FlLNgM/NHA7qrbH
K9VsaBFYUVad9BMiWP1UfTq3ymo/BC34fVGyqskW0SGzlgZyy1F3IdN2e8MsC3c8
qHV6q95WaIisgcjkzldC4E5ntT6+XP2VC7CwNnxgeTP2NBvdXCN4Sw+x6+EwTvHv
Mac5mNDRhsILFDxUKjV8C1O4r7R6DYVKvTis6EVNFTtmNJbMXNwP8tx5UMiXiCvp
Ork4ZusJzGiFkHM/ydH+Lg/rvqFOVP3erSwqfRbOvk4cxT321pZHhRBJkq8+WB8C
I5SN+BmoVwqfwDxwPqMwjecuyLxBE1o6f588vaIygV25wjv4l82FdtsuJFVVPO17
lTdC7zsTsTgvJm/HHWT1io4LCRgovH75NB9tdbqCMk+7cblrVtiZLWmjtjsGo1Z+
4vVsiI/fLmb2iV9QmBpYCCVVkIFIXeI85iwn4D72IZs7Lfi9120Dhhzojvyt+Zua
q5Ac1yqMFuzU+8YPgPHmuiBhajqhJhmQ9JLsuePJxa5IcDWIkUhAu0ekeD6PkRu0
aFQzwsK/FKYYniBucluuhvSpXmLnmWYKO8AvetnIU/Q7Rc6Y/FvFIMVKak7ed8Zv
ib6TSCHVYRIdSamqOA8DJUTRs4bIFGtO32TIsstFVCBbMQg3Y9vR4XRCrD7qbmdF
DMRFCE0XqhITXADMLGUqA+iBI+D1PJbh5TR9TATcRgDQ1f2NHKOVWLFSeFflPfqC
AqwXnFIRMYDtGhLRq8XK8NUaVO6BnJ8Fl/jYDeWIpMllZHbNsLvEWPe4nJeXlai9
tL90hT6TRw8P9Psn6Lt+lu5ZxBkuQZrTdZWo2Kw3LC0jOU8ZkCCogWsBv4bLKV/+
e+EIjBVRw7kENeMj+8KG55jDn6owb9w61k3UnlEOgiJxRWZGzKIJlIGPb5Tflevk
eFP8f2FOu+KcGe4a83jPd6C0qEE+J7kgGBVjxhN4XcbRzZR10bkRt84eZj6kpxwW
bUpVREHB+aCR98ZXTkUnOc6O/Kx5r2ZTZOX/Nw06yYce9Rd6D1QB/ihS0SkKa/M0
SVAL0Ba9PwdWZegMeTpeeFUKhxDPcbRykO6UaFSckg+8srADZB/wXyRCPATQPy9k
EZHt1WgGEfumSMQhnwby62yCHddx5oK7kDbZPXxsiVIpEyOz2dVV7ZL5OCrNDGOq
8AiHZMVcarNhP9IgwfMMT+DGh3MTpZSh/Vqjttd/TEXr7l7k+8eBgrDJ2mMKFOV3
37d2o5GOU/rQ0ZhtEWkvzGDqxzHHqq4W85NbL+3uBJHHyxG0yGm7u7uJ9PcSUVBN
OqS9ByApxscDFfzR9EudQ80SxGCM38z4aIjrPl3Rz4B9fMsoiyKQQ0eKTGhO6ubR
DVl8fA2OCNgJaOMO0LP97Qb8DF9+VIxKRdDMJhCQCx5RmIUfSvWb1Q4po67W/Cj1
ggs9lyMLXQY2qssWXOSuwYwQFcX5+/F+5Rd2JeXMWgrXcY42sPYjEBBxjotbX7xf
S5fFk4rmYuWDdMIoRRqihtB1McZC97PfDjgsKwB0IkzmTQbz8f7xdTMR3QY1Oyck
rgrDiKhcw358V9kUnIrlzgN9fahK5zcTb2YoUSB/j/BXhKc2iBs+kswi4B9uB1Ew
vZpF/m+o7Pf6Sc3A4IYmiERPe15SpPFnpxPuggfWyZVnck5fquVIcYhL1GlFB9Lc
o5lFqKCO9iYXdqEK12trhrarGbFYCzVbcI0rXIDWl+ic9r0V6kkMqte0D18UZ68b
aejQOKd1ujcymGfqCtt44GngLxfWv/87mNDYLegEahaAal4S5k1jV7HPPNSXgCgq
9YFD33rG0ODkcNa2O/NxbCdtTZldLw1/3MANortn3TZDZL+1NL3clRUMC+fz9S5h
gjT1LouAqJghwy1ZbD0Y8yXcE7Hbrh7EmUy7IFLlPzfNzOCQmgHYWeC2GwB5+3dQ
F8l40jZxHdaOslp8FCx81Y+R209LlVyvwPIrFjMhHkF1ZHm4tGv7ANis5nuc6Pnv
9gKT4/dqWu+nNI2WrKAwonQZ3MohOT6QmVMW0nDiRwN8+U2Dm9aIBjoI79rE+xTD
aQ0r9w7BZp5/MSFwNqoEWM0gJIj1HrlR/JgxmDdRomg3Z2U/YrM5Aa8nTgkgbUeU
ckYsNMe3T79AM+viYtQvHaxBE6H8TzyJqYqC5e96agCgIfmzHAD0fvJJ+7AsNVep
hMT1syh4jPi2MFqgVE3R0xNPI2Y7Xgl137o9euh0zr6/s8hEo2siA9kZ6/u3g95x
Afc1jDXjX3jxea6nkHF8YOe39DWicK6oBHNk25G+UnP2ONCoafm2ZbuL5HtpqLxP
cGuXbiI/KACc+0vj7LKK7+KIW9rUXBCkibcBTgQI1An6Fr4pOXwk3+JfoX0hJfHL
ZPkiS9wqbF7zbp8DRoq0QW8QXV0d//OZ1hlw22Ou94a6iCUtSfLS+PjREyTiUyXe
aMHtFztMgv4s7eEbMgUrUYgQv9Tg498dbVVR3lg/u0iPsIhIlVPrQmuzi+nEkxjd
RSabkHA29TSR4YFNulGi4RA5fjvUdLgyNpWl1NVgsOBgNNA0Jtui9zUvHCXZeLw9
s9QmHvXDQxplieFb5dcnb59ugEHXHAyiui5NCtnG1feDpqvyAkKbTEcs8D5zhPYN
ZuG3wUxhy9p9pN1QOyrf5Erlt2DCO27jvcuq3yeif2YitCo1+IN1vW6+ALfotyJi
qCQ9M3qMkGn2CNJDns/Txw/Er06yPCZmdbHBwMBompvhAUzX3NGm7Mnj8BlkyAzd
B0Srs4WA/iws98TT6GOZ7PEAHDjdTQR9X/kE3S2wVwETrQVivFVpu8VcUDdetb8x
z1acRKzN552DXonQ83LCT8N/LTGlAHApyLzWteR1o7TQdaxGjVMrvYZ9evPPJS/p
Zocv/wSudYut3QY40jI3ed0DYvxdnfJbFy0qmzGAZB313WPATC9wznO+1+4Wa2gJ
scituoAP8urdHIXSOVyuhXiEE6cjFkyLwcl4kKVM7GBPdp1Pojpne2utlq9qhPRT
tZe4tkM8GNnkrPDIXbpMI6QLZKqn4zJoUlJfTfqagqFYn3uaOWrAW+zyQbu7fYJd
WtF8MyBHAU25Iv+kud7tYJZbqvAWJRwdjWa19N+xUVPTMfcTB/QbivgjgZUSU3Jt
bui4ho6AYJi5VHK+RMkak+c+tuBFkAyiq/wSPorOPmLDhiWOgBLrrJbMSMs2T5PW
ZCXoA+/IWgb06bwLc/wQP4MTXHZA/GXyPFZTKOovxPOPZKy3rRey/avx79rIML+d
M8crYyV+p9CwqJ6iiHwHP1+JmwFgd+lbSsejgKVQi+SyJzQhoqFwdG/4PQbgX2eV
fCLKbO/CpdDygJa4KiSXu5rt+AosGngnjXZ0Kdk/w4O8QE5qXmqm9IVS44HOaITG
BAL9Afut3Qj1EfjFUoX+zo1RpfHarllSB73pXKlMaJcLbIXehpdEWmH/P/gCq4Hy
VPZhfU8zoUYA7cRPDezOhmkmQ2KK1xdUya468ZLCR2MBI2rOsb5Ws8N/pmiD9ZXl
xboXCdRrSGBmdwSDs0f54vGfKX+HyVhbgy++qP7SB0bKkd93m+IzmNJyPGv8yYx/
j0LEIJ7haMYaywoqJfc7bTPU4zamd9CQNL+6mC3HgadG89iYrdcQbyWhv9sYxFSP
YNDITYfnWM0fk6CRG2LQtQHOvv2CsF/X+7dL9ufSZHm/BuWDqe95VbigrMAnfSa6
a6Jf1sEc/xlbF68052lZzHVaIX6h2qNK+0HC5D+1JmSQafEcr1OkR/Mk9tFhj4oX
YkwXfs4V76ZfVK0/xk+7C6BrAp2JVHzi6JKel3WN7M0g07Re2hmLpdfSFTTfnERN
61sFU3wFIDnOgT/iyLi1zNJeFATYUTXC/qCMq2NDCsFhcW28/O60phBYy0FdR6pA
8irfNpxIKC5XjdNjZ9D3tWBUbwaZTrMfHklIGg9Qr1vX/tJ3+QEubFFWbkNcBU08
OupPUB79xlg7jV6g/FBsvJEz/vh1ZnWmoQRNG6plBRVEaiAaCb7ltSLYLLjf0+Q7
YYXkrShGYsmAGKxbSqpfuculcDwsi1GJM58ce/ff4TChbT1WOKLPGsJcZhGVoS0Y
aRfpX646O9kLmc/+7Onj02U++FTjxSlp/S/fRvZQoSb8ApExRIpYeJLhnxdUEOch
Awl6uGy5HaDMDwCdtFftZUyxAxnCfycsvI3/YHcamrWds0LOAEAaLStMTpZTDORu
dnPsEvNbQgtf+mX9IVcI60UnJQODHyKyjqXULoroEbi63QmeA1GjOcrvhNQfplIc
JoScHvJu+mJeHIG3m2HpInSpKZUuC1xYc2ykpkCWdYsQu7ozFG/ZfX/c4WBlv+v+
RA6EOtcR7yVFUmhZ70QriDNqomm4Ob2uSnOrx/xt+HLL5PFAlHs/IkQPM3lMbW7B
m65BHyd/BdxTfaxIwAaWmAbwsEbE6w3j//bAJBG8PU910Yyne1HT5MQJjbly1mPh
fT44shPAPoqKUuQXTpZojq8W/s2X9wzWsm//Qv0fTlpVuzouETpsoo0CnPTwce5b
PPuJbcCCdGVjUgW5bPe1ITdABiaBiSEaLJGBZjTD7xrkMQ8QGdufzFxaRhelDsBP
QDaxTmctVPQK4O8AZl6/PH8XPNxhRC+lIxqPXsmb1LLfocPjqFSvaIb3UcCjmMxF
82BHNbvObn43DoRUqT21ZMmIRHp2vBBeJK+6t0RtR2di+MdJt+uno1F/gIsh3G/X
zwlIKY12QJrHZqOo74B4nPYbeadH5MIK0BJq9F4AB8awDngAjN5lgXDFMQ6h9NPX
GpktFCqhe8ePZJbXiNSAx6lYmfG0LKZgU0tYidLCI+edEcspgOAFzq8f6fYHrVS7
Qiwt6ZY6i4FQnmji+7n81+k6GEz0zOq6t7FXTT8wdwU4WMwy0uhUDTp6ULyb+FQP
G0UUqYM/KdA0l4Fd6CuCpJVKUyr+9Gp1uvXzh4XUSvuJDoY3DfrZR0UnLWnj744W
rk/dMO2gb445LYTJ/mmsSwBu4gggjqS41DPTOJ1j76xpXhgFDE8p4QMSqB1J37KO
NYRZLJsQHFWIdN4MXJkr37g8/+dft6ZzzoQhf4762dBORsqI9Ehyd3+FrVixpwW0
HD6Ey1HBFTKx+vMTE5xr6jeQWAJOgtg0NyoadX+JA30Dc350GG6BOOOqXduAGac9
x9n5uwELbAk9fKwfjrOn+BMytPjc7rj2xG1l/qOpXnnbxp9WZOzSNFcUmRznBCIR
+EqT4d9VVZRMMyOeK2D6DV8LSdjoYRuCK8qFBzVbBazOoxq5Kq+LAfzd/mVa6moP
N/Ycm9o537p26AlnkntX34XbV+283QSMvPWsmde9Grri+kxCMxQg4JA9clFEvAiI
lWO1ZfoLqhk/4o23s6U5sHi1MknvnaW155L1nQqjVR0RKA4N8ykKeL/S3KNVxdi3
szLUhta+wACv4XfuRa18zuiZpXnd3SXzMJtI7YavmTqKIv6j8mevRFZUFt3VW8BA
7ssOmm0FgVOCDFdz/9omTJxBLD0gTtPQEeuVupGIXWqLJhAapQiKnhe9pGSXrXhX
HigYGgzn7E9MvhEkSiyQvYctBgObXA92j/FCrYNLo2yXG2q4u+wZ8fkibJxX3jEI
6ILWGWs7YQs+gitRoAcErPwKfxPxLAkG9Rafx1JkDIED/Cbf+zlr+hA950xlh5ZP
F7XT9MrwWXcaxVAuH6LUjhAgPljZlTozuT0mI4gvdi63lUhcOCsT2/F8b/wImdf5
ejVMWuH4Yns9ePeBzG9EoUcLYoHEj8tVPUDatLZtJSeD2BFLLpS750Ohrv7SfhQa
Fi2dPXAfu9J1zezITLuVTIgw4LdjUO2pGEwHyLVtAzLiLMV8ZcEpnOjG17BELyXq
Xod12d/EuAT8V5QvqHix/DKDiGmrKufVCNHxx2PZhPIZKlG2NLv9ZMHZy1tQfk0n
vhI0tYEFzPvkQqsXqSCUt4lNwdbxYA2vbtiw872DU85NdKc8OpS5jPtuSgASOldw
OLc5cRVQsMhGXm81BMMsK1hRhYsTenAn0/KLpMwiIZNWUkCkbwUE5xuZ1yLw36BP
ppoe7+V37abCDY6ouTdLEy0xYturBIgZaxJzP2adQB4eaw29O0YrcJIxHLAlID7n
4fFL5fijRFwo7hPWmxqRvslcKICMvi0rJRYHazammlTtqwP6EhTLC0TV3b8AlF2l
lf2HYsQAJY/4lgxMs5hkhyttzzzFLqZ0AnrfCsB5KZo31k62WlAI1OP4fbA8Ar6b
POs8AxWos5i0XGVlU9smjPNI4wY/WEXZnh8KfoTOHaOH9K94GJjOOaCv3vguEP0V
D4SwcGtaRA+XIg129dOsvRt7c5boqMTfUaVIm3l992bh0Thr8XSwkcVdH4zEsz74
i/BjtvZtnlZAMAwHpGjBzRtKowz8ybmL8mEfYh7dVornWIJwZv7kt79+0r4ELgCb
U43+ST3or9cvrc3SB7I3QZi+HE55SXOogdZhP4QTtPLlf8yi7IGE+jOsnp070dnk
dxNadZnGJwX6ZRYeg54kaeIbEIDYUQWVxH8xvJRFwhgg/PsQTRQNPL/Fm2hGpO0/
18Dbw52TuXm6FuQTCyWz8vzzLV+JGJwgJmY34NZ1bGZPJVdok2aR30g5/jCileWB
0ZB/EpeT0QaaaIasNind/JRDAZXUj8Npq6btJ5nmlAYqVytBjKG1Dm+b0mvSAqbi
wLCydlBq0r3Sryre+ipfE+5CPTVzaxfXTaH0JRrvjzeERL3ZRJrjMhB2yqbzmZB6
slnSr/UiV4B4qjV1ai8oH76oh53Aefm5ZAVJseD2NDfGUrsbFMvTChg/3B35WcMU
WVsStIdCApHhYDbL/tcMxKRAG6k+3itU1t5j8ABOy0kE9J5YJ1e/knDMf28U8ojL
SDfL+m9L67H+JTqxDHIXwcfiQhTASMD4pacMZgq20y9k4eMX6sq9siojDhYeec/o
vcCrJmCwpwJ1fW1IWeyTIiw4cmuOKbrH+Z6V2ssTZRFpe60VBiPXgQYdUUM7Ax26
hP8gIWP+3vaC8FtNio4OSU1AbmHhHoFBMo4f3KDHuW+fGiK7uM1+sNZ1MW5PmvCC
H0qrgnnP7VV8Nz9EzW+peUW2r5AV/7RGazxtrcAqIay3eEAJTRyiRJMKz+bmkS3R
f8Fee9v4kU+dTuOJLFgJZrR/4xUWCGxGbPCDl+t6mzRlc/0ueneMLc2SDxbCy3IC
bvLOutUfdcUTTyQ6y3B5G2lMJ1KBDkwV40o4ECFVls8BVxvyOe8WZq+39ATx78RD
RFKMCbnVQCcnizsdi1UTKDcuMySzO0xaJStgMGCN60QDRvtpDY7EIBmXaG7zm/0B
I8AsjFthJ/G5GX4owj051pAre0wBBLO+2pollfcGhQI+itlQ06fGmAJJHYrRG5qR
JbaT33nAnjXV7vTGMq7wQeLNOuDEKFnp8OvRJaagZjsj2EnZ9jy+9ywAfhl/xkoI
zh+vp8ZFSqMrGIQ3QPSzRJZSKX591SAhyewxca+X6VLSO10Rzvy8EoUanwM1zFeZ
RFfHKgHOoatal3JM9H6DF2APYWW1fNu9CQTJhi4k2aAPYvBQC9t3+8nZtdItblzZ
K1kr/L2qsI3jXNOconUtZnW9S4GI2jBfo23bZbD2B7Cbf6RWDmlRZKTEkdiVxkpk
O1fYBLQjN8XN1H1OM2xLrfqiDdy5FByt4yJWYg+OBhCfzkZgdd4ozXLpu79qglRW
5bcuIt4UekZdd2G+IAAiPDo0e0eiqKUGFxpY5bU8xVRreBplPqnDh1KrtGOh17Yi
S4pgIYJGsM7k0zEK2MAtKiiL1bGhjSR7d7QjjtwHhiwzSku9nqHREqPrVEuaWArI
h6QG+5q7d7SuPJrzyn1aRV20RmPKiwrVIfl6gSkClkdeh5TmYRYDHpfv4qW6NkyG
EEZGXlUkNsQ97FoTDA6LKgV3h0DjP4GSypMWNhw6l7XOKG3dB8reR3Sd6G9Al0lC
pXnrIcAQRH8CDQqy5Z35TbC/27WooIfTCHvsB8Fu/tMNwLbhadfRv+6fh5+ZoJs4
iguvPqO3nK+fpq1+ROuPNoLeMADmvk7lhNXLm8I68VNi9dUtg3HNKkae7GaPiusP
y73svnCInpM1vsaCfP2iLV6ofrd+dZr8fbwun8OPtaXlxr2g4WwBkUxBvsYsCZXs
1GvZpTy5dJmXd3Zr46WGrZ/0sTjnEjGELV8NQeWpx2ZQWKP0a3jkb+HgdFOC5iSB
gFtNmdzGxD4jPNokA+BbHK9NqVA8QbXbUASOvYWXPPEFSuRyr7szG5ezLNHPKFRf
7WvCmrp+cKy0sSD4c6Ah9XxkUiK6UDF3YiICr+ZSfN7XsR4h/pV9z10dTXWoCEQH
n2fMihFyt6MpEHcXBYaWCgL4q0M0hcl3ZfmAre8gaE5sLdrUsriHee+V0BTCBqpW
EZX066HZbc7Xh7nrPTZJnC1ARZ/9KB+xin0BOMqnYBu5VruoC/mVrYTrXMfcizs8
WdDHlEAbUkVrT1dpakp7b9R7i2tMzLUjPHiWoSoVSixzxPfzFrKEKCrPCyzvMTbg
mCJ8EWY5/EYkeQaMjzcH7MpxPamxMD5PgItDbgcd5y+rGYMTKiUZolvwR0xj/ejx
WZUWQhLOOO9yGLeELVGyx9SGaq+Lc1TVPlzWG+pKlo5fNWZ5xEfmRxyb5Oj13er7
YDyXBTUWwWxgrTb2MUtWxC6owUoMeGs2KP85jSUoJ6FADSqMZoJYIH24Q0sv4t1p
tzH6kbPCqmCkN22tmni+RrXifqa0xWyfb4lYzgusrm1NjP9FouXH3u5w7vMJXF2M
j7ZSlTx7YamNAOGyOZsW4hBw8gmBp2Otnznq2dGxfD2lNYfCSRLm7RsjYqaTSMQq
VRuEcZQA+4Wc3f0x8MJ1b8FOG+lYZ9Zce+L6JOsyh0wP6UZ1ej2Jb+eTqnByNrRz
50xeJrQxWmG0E7kpSWil0xG1YqpPLXg0WSby2j/SdC35TdUUFDbkXxUhtCd8cJ1G
2gsrPlOwbdLJ6SiS4AX8FDIhv9BpsU3xxPjP8a9tcGzM3eRXwR/av/01Y3F8qk9Q
IN5Sql/KYPWbRFn0Pa/kXeia2AxtmuPpDX7S7Y3+RygCtAFvQtXGwi8blzgBt5QF
qtevZBheW+hw893sQ8DJzU0+eG8FHRi7lsnVs7C80zZO2bU2UJYKFX7j4ArpUbws
IefLZANlZzg8qGSK/wYO668a7cYsE/ocu2crq+vcJwSePENOR8yV/0Xkdx3rdZ/D
Q4rG87YaIAgVhPo2giBNDeOtvo55Yi9rfS+O2TX+6aCrFe2wLakyX/YCU0yiZlom
BggKBu7RAvVb0QicCtSdrT2n5KCdxzvyQscfJ0h7ymlx3HCcjOSkosxiURcFVvOx
CDHyEw8PpXehjoksOq+OP3aprHLdRlMxfqd7eF8B045Tj6rN9SnF0noqKN3wJmxW
ruAyCcdwTX26+MZ1AeJxUV+5Jy3VFGAszSbMtWI6qcAdOBdUpTu7dkKVf4O1698u
elGziSBjOvRCRVfZHFYMk45YzQPXy9UDvcuKBPcKvrDs0yqf17mv2zqc3YfMCgqQ
/J57K0fQ6xvsieq+TReqnNBl8zPVTpBNAojQOnXRvfjUFYsa7Qy2v3wW3UePNA36
S+jOaUqguqo05msSRRQydOHgxlsUbXZj6gsBdV2Hq1VF3vFNa84vYfyxwJFCOX24
KDIMeM9CQ0yEX2nXwaKJx+yivK2u24RrgF1jZDsC4yvcTAemhSw24XAxN3fKYgXz
XBdeewtYqtncb5os3iGPj9X5xrsSeA1WNWp6RqaQwzTcNgoSGCmDPyaaNez9lJ3v
RJ11817cRglCGJIfJwC7bWkFxElgezuFhlr0k+lPeZM/6uRRrLPMFckVAtUHaQ/g
4eQtwuuuy7x9zJmGXmrw1Akhk9pXnhsZnCMc9G//5Uw9l5CJzVMZiS+L5IQR/clE
8S0j7J5/5m7TBk/cIvlTUV85WeqJwK82PEzEKgScrnA5Ld0dWf4NpQcwUpFXAHah
3Lp3UGRqEyFVg2lF2RqrDMJppWrMbGDydIdb3/T1Er2sf+lXzS8ExGkOCtH7HChY
mhq9x2eleW/eRRqthLmwXr2k5D9lRNByiGbJg7KLU4GE43Hoy0PZaro/HquSsPLv
GLw2WWnESfUx4nF+SNkPbVY8wmpSYfEMRgefJ1PCiCBR4sZtQ26Rbpsi1sAMK7Ws
F2gClwgLR7jY4Ev2U8k6epBvDf7J36oZNT/NtpWHwL0fFymmsQZA99PeemNLD2YN
U7NDc0H8zoifRHn433gRv6FG5nTXzmsdmkrhxN8KzR2OXBnAVyGkwRXg1rT05HSD
I6TohKbk0/BWjtqPrxnaG6mftoa1FshWnLaySo3dMLQGFet9FTbgPRzDk6BLxc/f
yieAgkYKh9mmc32OCvKDU4jKfbbQVVLhPbB3McRRt3lf4DTU8oGEjyjTeJUk5vks
xNQbO87RFTsXzcFXNGF3cvfFujb3dkduOPFnYVAUqRxvtnQpjmx5ggIilVV1lavs
+ZJhOeKLj+Che7zW77uOfoqLvEYNAKcQjiwsmhkUFwmsJIOY3+/CjDTr1gyLPIXP
f6AyBManXNvLyph+R0CBniJvHxlra4fRcOkvNznpsE2k5u63rxMab25sp8dR8Yeo
wZiox9HzInMxRrajFTv01NKc2jXgTkQiSifjqKFsbWqPFmr9wUzva8Y88lbHPplY
Oy35RIZyHcGv18WpwEycch4rrEfMVm6JwFJTa/+eRtV6k1tBJ52jwdyU2t6OgyEQ
ardwa/9D9y01kAr1E+Co0UWwGnbKbA5xShKdTi9nORUNjfELvjE6FHQ6jhZQuVo1
6AMiaT/5rqD7xzvzse/84cSiPuwsk25+QbIZthb83gqg37YRGHUvdgb2BlNoN+Pl
Z625jQXunxUBgo/4WfERrQNUXYFoIXczX4+UqWzC2s+UtYbczsb4asi4BWX7VrHH
PZDvlcC4UtJNLgq9d90kjjBntZUv9xQhVgDSirfF1AOnVmXC+PqLJa3/54L5vAoi
bmJ9eBSD2FSqJ1vsHu3Gpl7FTNcfgBVs3SrfLPW7SwWQMLSSaVGSYY0lbaIEtzbI
KVY7NjNiyYKEnUDZTJfJF0AGx3SAFO1IhN4c7Yw+UysymKFM4Um1jzuUnBzuSHD/
HsbnRRSzGV0oGKH0np0lwAkXYdodkcCrkbUkxvveoE2uqIuq+TELFhnWqIBMDU9v
l9oS9jDoP26416e2NQAb3thTgvEvqgTh1m+esPRd4M7xYrKx0sAT4BmnzxK//faw
u02rCf3TFdzjTQDtwodZWw4GSkl0wF2iBEHb5iQOiETtvqGkrAZGnoYyAH2kAh7p
Ux4uVmTSoxXH/dhS0Ii/h33MDubTK2SpqO+aU/la4kdU2vF0lGc6mERJxaqrdCkK
HMhxpzOXCcvtFnIvzefDEkcX2iRiSPlcfP9/vIUDjNItZs8GtR5wUzUEzWqeZWea
x8bPwviGlopA2lPs1EqT2E0U8vuhUXyhgt6cjOaUJM6f0idrGsxOZdzsww1XeCQJ
1tk4i6VhDbV9mC1SwLfyRuNIYaT/fO6UPprRRDw6RLOXkVUbM2FD3hOZT+3/Ti+a
xE6pIzrToj3ldL3JAba1f3JdV5fv2T1+9kfX0KRfEfe39shrhTjGtbasKp9VU6BY
lEKk3A0NDg4FLyDVbiKPk5IKxqXRCyYkPkgHBJqrte/4Nfu20qsZh5/e9827y05f
5e4XESiBnHb4mSJIAn4FDd1Lm8lpiKIEHa1dUaJmwppfCksHDxZkeeJ8zoO25G2g
wlWeheQzlY06gfTKYQsnsmYxwQe2wOOk1Oar3xwCQe+BeS1tbadSrtpMOsKtgxnC
FwoyQh0Nl8ayYYeWMhz349jlz0DHfWjpD8mfjUFZ0IrNxSM6b9b0/llKz4BKKNM1
iV3xpa7V5IVl9QxxeThu1BYSyBQtvNsCM0594tFRPmm2CkeqyjIVoGHuIUK4jNds
N1Jmiz4ihnNWXNd5IwQG2LVNGb2zjMF027qWmwX3Sjs9DV/ZAe9TW3vwX8ewVgeQ
2MNLyZYJKw6eY2fS8Hk8hohDbvwH1yNwruFHHF0SCZBOKCaE7arg6sh3Tp/v54TC
KoZFxurVLn2rwDGDcx/nWUwDFbxC36OGWLi1kdkFuwTrqFJg+W4V3n+KWZuvaoT5
UKAnJV9VzxwrwT72d/nVLTpF5x3/Fl9pnW8zfzOGJA2u54p3mAnos6I5ogmS3kHX
XMVa+XuVzH35hgLlclc4ZvphSzXTsFZjP/sHErzG6aatMpTkIKp8vjgFKV5bsQPk
u165CHQYcSrbX9aYpIFNVSzDKs2ZXU9vEkEb7cORCqLyUhB9keO0IxSw/c7VapVv
/v5lNQjlADXtmnz9E7pJasssFHW3zGvPdW8P7tsNa0STgu3aPBjihGupusj+7/8q
0mJsCwmeWC7nJcBikfY+Qy4PLWoX8XJWxFp0sm1H+PuqIC9mJilNPU2D8bckfA7+
+/w7lXko8twjqv9AaB0hglkPDr0t1EOS5EJsrG687aL1eLzg+dR6EJjFd6mYizLw
K8mCXgH84unk3x8qMO6BR4+ZIHqdPcItdV5N0E7E7uS3juMnj3veFMtKy10G2u2G
OLLzKX4CWj4e+HMpWDxmolQSU38zx4Lt0k4GMf3K1DX7ctaMdEyRwO5fsOVIrYW9
WW+rGfIDNhiihocOP1RU5FhjZzIIXcQ6J0aZucpm8fZRIs6lxxR6IqFNtUzwCksq
LVRSHTN9kmtXrOoY6ROuJuKwPjmx5Ra+eVeMVqr9ZHQ/k//ujv5ZcQO0Zxh6/7zL
PwQ+Xk0xjP1Z8Ua0qpG9xXRCTCELLk1/8UegCMp+VHzNh9D3TgmiWnWQld1dexFw
i5rtLSXlLbjxOYhUkmySBmfIfZKh6LEqspNgIwuEpELS5qg8KPkvw50OgstSuPuh
LpAa2njBMeH7ahWfzzHOftjHKM1W35hH5EVhr2Uf2AD8o85fhHSivtW/Rh25SnlK
qIuzhrxDaT+ZNoPTs81REjJrFQBLi+b5R5NC1OaX0Qv8O6xKqnknEwj1JSzP4xno
gwTZrohIUXBnSjZp7BLbZhucgtO2vEN3Iy75mkP+osJA8xVFlFkXazSdHLHgY2+5
StFIZv8nAytI7RHnix46EeMvNzfB+MDjZ45lI6JQxuQ0Cjh6HpG1sy2B5KSlPJhj
pgkFHkc5SYVCFn8r6+6dLxZdBGA2tO2f+2pStBYjpLcoAYb4OPsA+LWVBvHor9Fk
V0/6Apt93EB2/WD4xzK02PKZvh2xNvyP84qM/286jKxjB7HcswLFut3OKaVN3/ZE
CU6PefFsHen+2sXEwJWEStZzeDZLULzYifv/WFI6+czrMxYUmWuCaJwDV+ockWzF
RmGQekdSvsd9563KVqCApfoaRsil6FRMBEncJoKGieHH2Hz1fXgY7USGHPkGHU/s
BqkFLsqZFPCqs1zAjje6a1VvMHf8PtpuBonDd8Vu4kg4AWMRTnTSnB2bPjizdX6g
byqJ/sHTeG+Bi1RT1ykZL8WZ+EHekUAtVy+iNcNeDZi3iaNy52U2uue/tSRU0D5Z
QJxn7PiIFchQBT8M4blo/g2qCsP8+Nr131pu9Zgwv0GLjVJvwvxHCstusK1jgzBW
kImpgZzfZSHU8U1GOb0Y3hyik0fOf+p4KwfO79SQy0Se5A/77rjxLT03pMCZj3ve
AAICcPOdJCWdcH3KBZCKeLzlhU+kX/mMGku/sELBGdSwXX5bKYH6ql0tE5Xc4z4X
J04hw7o8Z1a4/elJ5F7TOYxdIoAqFFK5wcS+Px7Yx8q9zpe1DcXeh2GG1NM4dIcw
cR5Zgxmc5LK7CE5Udhegti/LsMK5g1ZRsjvHn+H+0XLQinzpIfF3QWJNpW+LFTWu
q/GAf5jJ11lLFDH1OATq+JBMhWL8QKktVSQdtm64nFzd5V8P1jxDnsztnaJDNbp3
GnspL/jVbSLB/a+6hU7PttuMiDf08krq4MX7JcXuWThklVoWyBelJzrmio55TwfJ
VPmX0ZYpENSLcoskJkhYg1fZhy/W42nxi+pAFmuN9fVnc8XQr+GUJn6aRXmk2sha
2/grwj6aifhql5Rf+NhjLKSdWeibXL5GXUsQOIVUpPA+FKvpnZoARFGCs2VqFI/d
10amTnML7psSC2EdW4v51uUFerAdia84bTEHb7svQJyd2LOZmRZ20/8QV5PHiL5p
Qu30wUY3H2RbjElpcUz7T8KLcUWloAjEuuxKd+UzVY8RMR+y9ddqzK55+Lbzggsb
89huPo/4LHYnaNMV4B72ah3c87hVBRUWWnKfGgUplEHA4QoPUVdNRLKC5YZHu9tM
u59BF3ZV8p8O59VwJ3sT3smOFH/14sz8hx14ZqtGNNu+MWmH9hh//hbjxfy8BIG3
jNfIaP9MZev/VF3FQiqMCWpgiT45rtJ8aW6FvMq2i+w/MRwNibKbDGQ81mC8UVZA
Hph1+TyZ3tz9DO46ItsWEEZxN7pluUiFIb1PELNEwsZeozG1gqNBoWTT3MCIuPIR
Uuj8r1EUW4QxaO2W+CgL+EA+p/UXUaiAtc0hLhUYkFBLQ2NbOBFBbghqWbGpFBoK
wGG+J+PNjq0UwOGtdilNChuYjy4uULwGhAI8eenKn7ixEtHpszT1EaKL3k2Wj6V2
Eco2+zUUlZFFW4/eCKgZdRobx3oP14iAzeGOkKH9/pEycLyElF5VZBv46xB9zYXX
Txbh34vieDK6rBOGbexgTU+4bKWOIsZzvltsH5xdOToYl29t8yopcyetQK3+VcmN
FEpE9PrOv9+hTxZNUE7cFweIqrPvS8iotcup0vlZN+Z6WL239nhjAGMTGDoEB9Yy
1DMfgE+AlMCkbSp2NDuJWoz3EmKqg6jnjRY0c+w7HQBAvrPhNwCtRFbKto3hMdXx
4BNZiH/WMITrnj4NSAmucJM9N83ry/BY4CYyF5kLm+fvSYYWw58GqlDwmgmILZdL
dhpQmjsszcwx1yM0v/SX8X83DoYfZOlae53w0RGrxvtLIQYRgjvzQNn705YjE471
TmtS+OLR1zFW8FeDDsmM4Un0kySvjst93sijK40MJBBw1xajECb+KVbVRtLdRZZK
JA6mVDoUfiqbYgy1tJ4uOKgD69eckdchYYzBZ67IZLajgtbcX6uoJPciuz9+E/Zy
DO14z1/Tf2g4wxN+sIg/Mi76r4CPNECbuZQkzhH3Lf5anDJl9vbfTdS5nFtcIHVb
69FjSaYOtRKgPl+8rYUNsqoCF1BCQMThOpyboqtNgiqKjJ06Pp8BysmJjfdb/U+q
67o0QjUrnbCQt3KnOJzyETNhh8zy3hcYdAWdjMJMKsJ9NbPTCUsglhV8wIRi2w/2
hjKppFzGdwQIXnilHvLmAI3AAUt2zEHISAsuh8Mrv0pJ7majpfhUVgHmVDtn2sFc
S+IwHL4mUXy2DoKsMVcdnA4NcGrbLTu6k0dckLSwErSWz72rPI6N7AeLtkbN+eyI
NVyz63cyQd+RUIXySyhdBAXrf29DxdjZ80/jilHsAYJz0PLJ1Uff9FfLXb8NDVH8
0JFH8OKdQ9dnPoZ/Ead+iVT3zXJ226dLLn70r9fRn9Cp1E8+agEBvspLvdo8AuMD
rI2wCm49g/NDiM3/BktJSxotfi3tc6b5VFqTDOfo2aWv7MKQhgY3ktlopeVbKRaB
S5Cnm/OW3wNbZ1XENIRTitGpGWwxWyU9DUnXKcZVq3pyZaU6zvS29LQT/s9/YyWC
r8pdUjzr0LN06FakbkeUkmRSk3sgAFHW0jOdX999pyXbXG+MLvJox37gMbXQ0Wz0
uIIi8niDMYH0E17an2RohthGBqTrkT4kwcHqJiuMzucrNemPsUcwJBa58LY34bku
9MNFyYXb6GvoNAPsawWQSI5I0RL85SlN44x+zNuABeah4VXKU+hxxaLM7yrisoFo
/f3lEIHq5w4iv/LwlUviO42Lb5ypPMc61Mk146+KMsfFnjsbCTupW5SbWLoAI+ra
s65XYbIxVolas1jzQ0JKUU/xwHWcAywmZ1+Hqg0lgKTjaJ4Q4cdKdJYKQvHLoRiK
/RoWtbDhuARa7juRgZVPFuZB5TaqzdLRbpmNaJbaGtAQ8//L0Nxbico+yr/adaRP
kE4ASTtnOOgnvFqFCL3IThz456YgypEoq7gwTNTexLqXfNtw3p56kB+JXU45U0Ow
QT+9EFjU2Oz5Yigan0lKVDhfxESPBrNGj33zongl0v8EJjPbolrIG26VFTXSaeJN
k8YbyzCOHUiPknV8vL7q7RLtoopJgI9r9861c7S+kyzWsheT/8VOuBwFR/2I4tn3
KHY4fytRzGZ1nJl29f5soKbp0Tie+0MHnWKx61M0lwYvJ/LlxK6umR4rlPDX6im+
dRK7oli5RyXbyDtBmQD81IyFKgtkXPywfIIlfRxVjvOk5O6neQPQ81o4ClbmKY8a
bgRN4PjnSdblCUKKcyrWNiRbnTVCwWLdFNd1QeBEeqtncei0vHbFQYIqNmneAd/q
MZHPHdCvwpt8y8KlUWuek2weiCueJxsybVl+g5xHq+pmZF3BKaXXwJuu5WA7zj9x
yU/G1UwZH9Im9x47HD3YF880DNmQj4KlmMHliM/yet5PjYLNKHCj5piihi8pyKGK
mP33Iv2HVWpgXTJu+6P0Zx/wOXkxpWEgKQExrw2/ni1+AtVbegATcfQ05Jpxg+zQ
JeIz38KRZCvR98EFwyhWbxvSTIlP1V4bjGfYhA04NwHKODZX4sRrgek38JbROv2x
TN2aOOjeCD3E5WJFDd2KzC/uRs1zhq2HUA7zTR4uwQT3rOvei2KXpxiLOAWObWZQ
1OfwwHALLMqkOiVWZN8AZkM8nHNh25XW8R/Xy8QunxXSjCAvdgO34h7sR7NafdG2
pD/OZv08JvHVWqxn1ipwhVHR/X/fBRilI8Yqup5C5SSbICjgZ5L1e2FyUFCTv93M
eZJkGnrsjsQJF08I9nwrcSrwNodMwv74Dg0R1WAAJ6GFZ3LNzBZEFsCp9kZwV1b7
/38LC3fEyntlm4kaJdDyibNFl3kdJI9DE4k94i+mlTfFl8Rh/O6ChPl+StIas2nm
7+HxISzMSbWnEfgA99vFkDk+lpgEbRecdHpUFhY5wEJYOzjjVgPEzkC1A7mg76iR
xCl1UskRtK/tDXZky7Hn+FfFhr3A2AsvcqmZvRs9ZFQbj8FLEtofR3Oy8NtJlCn0
9dRH5UY2Tw7cTG2IPlLXMBMCLEyBOVKigBvV2WeUi2scrr+O9xXk8/nxQN257tHC
/3juo+uMKGzrasTiDTYWNmmN95ZHSyweZeoESFR80oPavXVAa2F1P28s98F2sK9t
0EhmJqZZ6az8UglyEQWbHyhvJikW+JvkTNmxmOT7937TH1eawHSHGURCkXqfrBbw
SOhiVbroztKYyiw4LgR36aX0xmLmlQ1aHs8EY2bH353TZFIIZ9useETzDEJ+ltan
OiKJ6VsbzGbdjGGSvemf3hf0oWJmRvpcyZ7TUe+Ld40tCxvvstVGTuL7o8iWsTTw
OaJC30XtGdb6qGdFTxqe8knOqDw/YfyffRiQEr1tcGVShCPfs7SaOnrG7qK2Umlk
CzBKUpCDllLxzUkvYGsc/TjjM187YB7/y4JAtl9AVh+rWdRins/bu8LPZ/Y3hsFx
cH73hb9avW1Xxb2d2nPjnfWyZOac+oqx3BI9rkcOVz7VQU3HrZmq8vC0myISvVwY
qH1f9rTTSrY7y5WF+DZNjAphbFNqmMf5THRx8NDolhHTDW313nH7GdNGlNXzDw8L
DbQHalOK1MgRmkN46ZCRaf91L8Evp/VsA6+o2v5faUtVp7hcPmS6vObjiRyMI7t5
dtuVWivDFGOMX/Z6I93qz/2KKRypwq6vt9gGvBR6sbkijh5oeZUHObSdNtCQuB4E
Mc5hr9+iMrjnK849fiu3iwGuUbVyR3AGr+is15oO0a/sHegqrpTfQvpeIKae71sf
gAfLz93mupKbN71xRoGuPslr7TN4DY2TSFourBpKdjcXk9nIizZe8+GXbilZsLhE
FtMr9sHLWoryUxtQ3Na1eFxy3cmoWRDMQ1bwpggiQPvDpafjc5IrPgD1hyQYMHWd
RAQ6SezcDoIx1iwXWmdvh9uSIOvjrQGwUdlQiFy7+6WD1/UMlnLc4fmpWTm8RhRk
GakIeiVKmdZsqxBCrobOsNNRgixcLDoopLkDqe/guRr96XjMhetAyVNEB/+Y8/nN
VQh7Ou3ZDWz+fW305JnNFJ9oIztSfAuqO5cq5pcn+xluQ20oknUJN4O8Dp6AzCRe
maqz3koXtljPt0HRStPYiinUTW66zclMoM0YVDD8BUcy8PeILQWYC2OQFh6G5Bs6
9FJVlE725TLLfFEtCFeIUrX6qIiDYDCm2waKv8twUoTiJnYPSUxLGGT3pcsCOAj7
zAQdwPBYwxCk7wIC187j7uuNjQGe+Eh7RMAGFk3l0i36AU2xTcWEHHtvYGnkR0Kb
Nw7O8is5UXSdG1enLkeckcm91rb56vilosmnzQtUI9bfg01GBquBrw5RMVFtK6EW
qj16Srqk4ZFqfBfjlSZcCsJRWW/+QjKKgb7QMCDwSz2+6H23stJuhjbE+2iU3sET
5GNsAlFwZVgwU0roVKRuk+Lsx6kGLeS3kiJpr8WS7ZseQyV1jt1LZ2iTtjfRIYz6
nmn5GvqLPwZX7Z4vkP+5KAVBFC7XCY9Nf+jlw4gTd6XfHSrdhl31plZPCWq7Oy33
hVzQ0cEuHW+hA7i2l9QTTOlYSNF7N0og9wCA48sc6N65oGHox9foP0L+SzqW/L/C
5FVJcYvapC3rAaj2F2BQ3Ll1hshTqZOsciCey41+t1Wlidt0rscGfCOMki+bTxS+
Oa6XQyQ+pzJv5kv4CUfwEY66WLNAsxOrB5PCtAhyy4Ppe9D6T5KCAHIzMAi+Kzam
8+H99HxB8RI2akjvFMdYLBcZORvKnDq3gb8iFHWgZSzIUp5VVu16ZF9UwHZny605
Zj5nwn+035vP6nj44EN4JBRJjcbC9KiDFXQ5LCrE4v1+KaAGvThVgV1aJ6BdgZYy
gtVEBDlkkfDka8FkN77CDeHuehPIRjDwkpvU8IDZdZQlQqzJGRe3XeCmjs0a0twn
ttTfQKAg/Xior2Iv6FkPO05XNZi21FyrHVMOcK+hZejqYSaEL/fTIKnsTAb7VPHk
BzuAvXsXFVPKGaqpE/ah+aAf3EU2F69NJ9mlCzqU2qkuyME4m/fXXYhUhIryK4kb
FHW7xoaJR1p2rlusb+TnrCBdnxPQeU1kXaQsOyjY9vA+8SMyB+Iac7XixabAIrMJ
PaOwrSNpJYyg2K25cbn465QEDxqTaIWYl92U7RQtB8QhnAJGO4Ug+f/RSZFbTXug
qjbtIsfU2S3KV3AF35vx7uNBYorTGox53bwf1Z8rMvmBph4qOmCISt/PW3gyxQpm
teH6MaEYpAP8MFpoO5n77gCSxTGKClXchgvE1p/+c1CzvIQ0VUzOMfgF/UZ1qVoZ
zA4hJdr0KiozcgfMpnqymaE9/K4DRsuo7iYXVwmF5sn/cFf6swSrH2LNKkB8qo6I
CM4Y82/A+y4pl0jvjVNxHrkSuEYqf7HU4m1hFs/HM7MCEfb4DdBe+Op0t115jMOu
K2IHUX7R+EgnirC3XMuD4gbC+OBDIYVl9upkjDkypWgjtfHn0/LH0bl5xI9AVYfv
VoYY1f0un+gpEW6EpR4hx3spGILWVelCNPXr4y3lWQ22F0nvcFrJnATkuFwnDUt4
JEDzbNWuvxLlH9z20zaOuMjI622b/B/H4X9iL8b08ZhkNtWs09HycEhe5i8fMm7R
GRmvQtR5ahqFAza9gevhku1Rto9p6A8JL2PBNywycboB76CLgM3/aj1UW467ZiEP
8mRLyWQo2A/CqGg4l1A5oYO6kNa0HVp8K4alJwbkjNmeCIivMUEMeFFlbAIsrIY9
ApB/M8SEnhmo9B3CeERRERTG7cvgI7x4u7K7zexK1V3VAlmp7Iw8vHJC3FMSWWl1
kGVINl7ZMcUaXlUcBR7aYlW7IrAoxalaBs7udVoDJ9neaf8rokp4LnWldy2X6hl5
1oMZIR7o//2VMZqfa5220EH2F6B8C+ZJL1p9uAycsK/hcA6joFc8Z2gyK1QKmy5q
oCev1R1B+KKnrfwxFIjTsck6jUZIQ+FqvCrME/IH+RT9+XeUt1pV+P6Lz+U/lWgk
A25r/gMZlalXSdcfrP3uV2dpNdgjU8dZbGJ6JWC9c/zscqVlLQ3HyNQEcJ7UiOY6
sGRnu1HAM0AicoKoCDCYjaaD2FClUn872uVeRAmQScDESuVnOl4x+A9QjYThWdEm
Ax2gJQprLoLfULdjjXhnzGpjiut7lFUhwEpgtVwoIKow5Ft4TtVUqB+M9GdD2RwS
MfKMur/7J6w30GAYOT1hdF69owpLsg64WV3PcBGJWziuxmoj22fS3Qwp5vyGYRz8
wvtfsR43eJf6dxsP7ERghPyiLRTHWwUtne8m6Qlgs9D186/2AgUgP+LIc/xEfdSM
kn39E9z8xnmy00MfvPAX8dB1yoER/cmTrhKkUk36GHLygGXg6bz/4/YCsCqdRCBA
DfxGGbak8Rm9xlgYlXG+zSUHrH0zuo3ALQ4CaEO7vphMdtibhG3eeTpKvZf990jn
t0hXiMnyfa5M5BbH2ct9sWMGAaQmT4ek1yohkEC9RoR4ECS7Xhu9WNREQ7d38ysh
h6cFJnwyvTa1hSpdZbsZhHi+og1emZWzHxMkec0ugjsGV79XXoiOXqar/e6S7zOh
9JYmnrP5hCQ8rd8ZFhup96hE3RqlwkQUEgbsvcnSe/d1WPJLtIteBhg3ij1T96F3
bzqzf+tg4caR6Zftf0Ji0joMjzHxC1u1/lMHhzF//zqCu8Te/0Aevbek+3AFCeol
cQMy+8SvPw9BEjaw7YmhlmYQg7rXKNB9lbeqGaAJi/zLFMnTK2n8qBMvPBU8zYKR
SIqn5i1W+k+rdcEiYuzAyDgjV4kTY/w0X/NQuQFmn5QX64uLuFmMASPeHuxyIRfZ
0V2j/1OP7NyfKvMq9UuQMHqC2GNSTP9ICtziWlhysyz5ahcFrR0O6nY/Fy0MxNuL
QqhHySisHBgO1gqFCXIOH0B0GNhtHZxBcLzki0x8yFKqTnP1PGTKxS+YG3FBxtOA
IsS0OovQfG0wy0M0l3s8O0KO2QVYbDipXZORit5vPsd81/Sf4s3DB7EvrewxgIOr
G8nT3vVH4QPf/YK0iy5kzUO44iNCSEn2WLxWJW3iUEWy3Jc/igbPcD9Wt0/KfhqK
PKkpJYQFLJkGTZL6JP1WvMMNgALcmAKYbQW/Qd5eaHpNtpvmGioODogATsf8wcHS
PKPvJfiXikq+oMCSWrHQgSS+iEqcdb/ankdgC1j85RMx1jULJTtSFi25ku72gUO7
bcsezva0JCFRf1JdatRy7la34t7w1riW2HFd6kdsIn0HS4IeRisz3nF5wWbhIb+D
zW0VWwcCp3hA/dV1V4suwyqkSyi5AcwT7bU71DyzbXbR9rvNYYH9A9QJ7GH44hD9
urg3f6o4vYnqXQqY4QmPrRL9NjhUZ9+D6yVTpgVVXk8n3Lrz82X1wPfNKEyPCAJn
dYMB2555wlxdolXf8hiBmnNnO8Vgx1cD+jkT8YfCv+Nxk0toZiMYFPN90MX2K/fO
Hg4DRbS9w1z5Vk5vZS69ubGvslJ9qboBzWW8Lc6KcxJTf4SfTInHAANO5MoC/Cb0
UXnzp6QAYVbE2EMni84oMXHq6u4pO17t87OShvju+H8bSEFVNGIk7de0tBiupdVL
HkmAmmfeJJDXxQG20ctQdQUOy2Z1mmAH3On6Bx9gRUwbW3pdxXhKqVIuzqhpjIO0
NWnffM7zwFOqeg7srrXhAws2BsHdv8MnR59OrkjJHFsGDW31OJeFlKa7DcphOVR9
XtiR1xZAxLzutMy8Og3BgHbI5KdmnCYp/xbG0PuTYph3KFG8vFumZ9zw+EziDowD
4Hh4DSyfrFhPAZXk+ponEoHYk+aip0VE2Mo5lXqNuhpy/RLZKAaAu8DYgfNLxw+4
2rgTkNfNHY46cF8s0+W+CS5h0FaKL484ul1ECein7zRBHVu7slTid28EHPQZNm3k
aipixQq3wh4S8J61ZuXvZGobf0LhE3fB8PbqPpG7D9qm+mRIQQv/cL1sQi+abW91
kDxygADnij2zBAdpfSMp+6o+dmrMshX6kv6OHPredtpgp8F9cM0hN+iZbWH5bUBR
lC7IV0M+zm9YItj/yLizluiXzVpXiUSXMpW6nbQvJ8Ve/9nWPsz7R010J561Ak43
MpC3srPBbrvuvN+tFSb3+V7Fqy6XYB00mW97VzCSFB+GcOJjuz9D/g1K+sh7cBnS
ETgYcLvJcyuA67Mw4h2tkI/5QMbtkR6Z8p0I+cMWyGMZzetRV2kURfwomx0prqRF
qbt3i9S0UwPg4wH1V2l2O/uLLaNkcJNAvPOMeCbfueNI6tIPjuTDbFbkhGDXC4jN
cQayV/RF+PEDeGg1pYExO+pUIA/UTM0X6GBmlqA8s48eLrnqXE/8/u5HgnRMFFS1
7Gdl+D9w874iBs+7xLKCno39AyYU/6CHZ0owl35qWiaXoIbNoXnVaMn9fM0I6tdz
r6dGdch0HpCs1FDkUBsYWKGoqq/oyOCBxXC7pHGeGTKabtp/ChsfGSX1f7awHNrU
+Oyo49Bjg6JhWELS6eMJqOVJyNLTdgKS9CULyo3ZmVvIfxnsDnSbKOuF2GA25sp8
CpVGcazfmxZ0p8b4H76cQR+Ld7HFsUSo7cBSizuqYLNNOpp08WnbbxNJuq1U/jG/
7N74zxuvEsx0L3WZW1r9hya4JJQebBHRSdvnpRbiGIhpfHYVpDZdbxpuTwxAtexi
/fNpDbgZmgo4OKafAqJenUgvIli+MOaKw95iQ5QmKjHXVWSlEIA7cWnF91NGtkt2
aeVy0UmCdu3ORo9z1slXU+ZBwto7Hao3MvIQ3PqWDIyOMiyGL94mrWqoVk+FlCfL
O1nPHk/66wE+axuqmzfE9Q08e+XfF68nmsKkF3GAdJUx6GiNTISp+AP0S7v2e0Pe
rVyd5lMd9xL3zFg0v8/py8zZ4sPSu5/OSrNuN2SlqvJvue5Hn+aR/dvovyqob8aK
CcyJh5w2/t3jzY+GA7FCGiejhxQXG4uKptv90R2wKJ/HDKekKxsmQsYMkkUIKa1q
6hD7qQTd2D9ytICk+CqQMi5DOO5SF9A3J+bsRAKoVmB2BdT9Gnfa9KqJakT8XEEN
TQ4jwslNBvpe1npoEIpR/nAYa1bqRfKAoVejmp9AF764sOMf448v91+ItdPbLA2U
CPhaG3DgI0+3XgFQgJ95fZkTDijjRfNMbpCtD1ZavYyg8N3xIZZE6tE8GVgyiH6u
+CSDtI6d6qavZR2+Pv9isb6EB5EPqkLDPN2XviiSRJLvHRaNmZE4aXwEZRQ40JE/
FkzdU5cKIr5ZP0mup5W52XPor8Pp6CrUonQvsc1c6DCB8L3shszYyMuRe+S5YKk2
cCML5XaYhh8nQ8mb+turn38523vKoQFssatVdZf1zbSY/DP+9B0F4C686xgc7rLs
S9zV7SAWTEUMkIMrH/oUL/rv0KnQdmFwmf/shRhq/vZXrSuaHRI+nXnRL0YqKIe7
DdK2/XPFQhBwJNg0eWOSIkp3qOwKVwyU4QPw1/BxITik/+vfG8uuNCq7ZFT8hzJW
c4kFROKpzozRb9haolZu88Gch1yjuHLlxMC0rrwnm+vjpB7HR3DJEBgBbxrXEfu7
uXA0J0x33HGWX64m2wVKVXyMyfxuNLnZq3Hj8sFaM/azgsIdFNL6sMQ0vKPNyNVj
6jPXYy/xtduo08cMLdsYLx8+r/tBNRj00VbsTX5fRQiGAOatmcRqCPi7C7jpTM7D
CkNZi3GI7Mv7RScb309kkesZIo5qdsqETIQYHYZGQaah6OIM/szkDocR26EM6A4V
KWabzEnGMqLTXYUn9hHh1pwjvQHZBEkiGbZ23gB6s2uLAS3oaArF5UHQLSPOjE71
z23AU4XwNL403FDw1P3Xk8sO+4C7qpRx8nEC6zw/EsOnXfZFgIoB8FLDELIeiums
V2kvA3LLaFapxPk+c8fjv1Nrl7iLZ1DnfptJCies46q4qQyG0f/hi+HwuCpQCh2H
1qxJAaRAiFpZ6LvcXWbNhJYOCP2FNKcNCLjQTEzxfnk7EfUZsfAgARYn2xyy6VgV
2Wp+p2+ApEEpMtlyxmkC2PI1AqB5E3RK4FDU2oB3dhOEBD6CeZCpNPWPwbiEtdJl
cTYcmLBUeyKA3Rajt2JE8MgbI2MP1SAtZiu6xot0reQjUQBvhuG1Xd/SgpgkRSYG
G5ZvsOroC2MoY5zVxjOfsIVf0gN9ybZPg3Hdgb92NJHO5suO7nDglsrm5Ivr1/9z
juf4S+hHMwjiFZt08XioDTNsZyfnOSV/r5f+sH4OnhtcWqKV2uMO4P04yJDT8L0J
Vl9/gut/Dv9FP81pbayHKq0ZWJs339Ef6Mb10H3Pk54ORTd919jy3bXe8V+12wlK
dcFRAnYSoDjCp2NZgWYrZC95M+I5eldC9x8oih1cTdV+LwqtzjCf6qukiZNf9bd1
os9TWrMs5Ql70ONz0+dyYeyg1yXPwEdXyHo8ale7lJIWLjbTevdsJHXBFMsIMBZp
Hpf6o/yBqw9EtulG7gykZNLJ2fDSm+oq00eFedb2nvhccI+yWkUK8+6vajE0SGSd
F8kgZicdmwsGqCpThzGPnJgIkdVTzG/FZwyKyGHjg/qBTBATR5Bl2XCN4aVBNkqy
RAec3LVapi8JOcjQ16baNFySkMY6eXBZm0gYB1L0UFYYkZHrYrtLsul3DyS9FYR1
7MEapzJTMZ1970uMdY1OFMbiJ5Mlu4tQDfMxjM3skGRJCytnt9osKAGVgLoIObbB
R4ud249OijRe4HJLA5SpIDIDJtcBZKxKnla17CUPBMq4asKumHpCmvhKnBDrk+sv
izDeWJ3CqK7PVJOMM15xmfEvzhdS9Ql8YgUXKqk+80evNiruz8L/hR8pgTZSVVN/
l88rSiGNZthPJgyKmVlfdDN/9eLunq8nOFAgtNPcgHhlANeBaboIOM7QJI1Q4o7o
L2WGJWJ+rVW5O8RzIkzByvc0v85AwfG8yfUeL3FbEaRcVxrx7M4oAord0pSRrp8y
2xIkY7cmltzBBNTZgSM0DWi7Hc4CNKXb0tyraKhL6Z8mGYD4FWc5XrjuxVr5Pw+C
7D8+eRW69eTH1DtMOs1uHATvf6pVIcPzP9MRXlK8Q5LkVFVwJRrER7PUmhVxgjLz
qHs0p9x0VKb6fKG8Yg+MoghaXz0t22gAM6UNZjRH1kd4jvh4JRwgLmJ5/UUA6sX9
GnhT/pP+jCV9ir7rqiT6RvI/OnFhGBj/tKhXTX3B1xtN0TU7OpBr5CyWHKcT8pnB
tu5I+Pn8ziGP13n9/+CqQtmXhBkzDIj4Zxs9G1OMkG5tARLiRurTzmBv6RsuTjIS
LBX2dIr51IwmGq2bqSXQkQXp6yiA8qGEpt/pm/kfOZCVoNW5xxgdgEvHs3TOLz57
wFjKeEI+BuSAaco5W9Y62B3mbseGgWMTAfAO1YO069N0y0H8QLroVW+V7bmoTYlN
yc353u9W8CopQc0J7azu5Qhvvr8lLtZ1kVRPW15ZkEoBOWhFyo+I7sg/AfFCXsIb
KHf3yfm3yAhRm95reWfVog8k2KUsBJQbUmTKphr7V2EnH7kL+/mtlHMIP/rp7Gdr
DmSOI/k3+ayEiI71xMTiqz+z92ELxj7uRYCDzlxKOY1KmJz5fnAuBfJgNXF6pBLb
VpRJKczYaI1vaKH7ltHMQ2/C1ZB8OTKibz5sdhcuh5aBAEpc/PuFeTsqPEsBjKRD
OuN9yJWRGqGbP2K3Iz9HG2sQwhTjdq1EZSsbGAR13mCm4AXrF2fWYqen5Cr6T2sI
LKRdfJjPiAKEJBYALdIJluPKy4lLFjRQokGsnrnUbMeeGt+UTNFy8H4wx4M36wHX
KUgFqWSs0uC9cRCUWfBppgVQbfUqSXxUp4sqgyKz1G8GtRN83MwdEJ66abQdeguc
En7hPe5rqwFB6zOHZZGTbpT25/4vfzhUK4maewt5m9xN3V620EbnkL2EHdhKew8P
C5YFcQKvnCfB+i/Wc80T82jOpsc0hXQ8W7ErERNDqzqVK4hXYeLERm0yPrBN4ZZT
fu0c9Y/IC67K/KqKN5WkU+J6ia4BZj9WkmRXKc7Tb+p3FRhzYfjMpnPkvt6fyCuu
rcCUy4WSriYAFNSEoZ2i4qEu3PdW9GbGYs28Wn0STtGYZ1pf58pvjSw+wi7rZO/1
0d3k6qHXbS2YuO4lTB1T0RWwb/zqmqlfIxaV0qxgqEhCakda9bCcNvDMqgBgGAOa
QBy+KrYr2DXsgazAU9iY6FKvVXYbJl1lhJVmOzA9fC8iLVPgQ51Ze4DDG4W1601G
5U5IsgwwN1wVODDZKkYPNtww7l5di2bfEowxorJw5r9tR8erEEt75ku3ozdcpf5u
O70QHpwJ4lbeVsoo6Vas/aWk6fx46rnQQtzix7YPH/I4a2nL3pElMnd63pnYMQTP
QH3Iqv+VBdBN5pCd207IhF70rVfhCJQUPoZiJnPrOQAjpH+NDZ4/uHmIdSV7qtME
JE9u4gnZeAonLi12livZpDp1jgKW7oy5pRnxfhEP1b1Wbqxqo6FspNEDp4qhRlVo
wz57NX9ZaKHhDAy0X2SXMcJPgh5EQFJbZlWAk6XeOv0eVf5c+E5vvffu+HaN4r4Z
tJWG11FUJDhiokjjc/a6TDD7PKyCvT6v1Zk0YeX2xIZQFkaVcvcBGrx+suO3vsgd
wHhImvd3N5Y3pbK7XvE6siY4VUsSOQD/clF4onFN2skvRQ3YyEp7w1W8BM3CjkyY
EI/ea/mhpC7NjW7YyOs2Yi4UqJR06ULsdqCl7WlRfiq4w9Sg202oyOGx8Y1GBk27
KRzYoyCvgLWY9A/rd+TJ597YtON/yGpw6X2DNK/vtQJ7h99jWskrlF17dPfKtHim
nlUTgGQu5VlQ0U02rOY8YXf6pLZ3UjxU39nb7u5oXA/SfaKV3LUhabWbSUmMonnK
101Rvv1PcPyNuubbOLdMYLY49FWCsjDkbKWQ+23Ky+BKLBR8x54eLaX9BrvabnaU
pxESi2m8/Fggl5Xa/cK7dyv8OobB1+nQ+sLXwWqMTFZnpjLueoNkqy/vRdZPm9ZW
yXApbTVwpR7tEGPaF8peQtXs7cXAVV8swuCEEjY8KcWKwA3gs/IAN+NRdPjcz4bE
iD3OAuhisCGPKgmgsWsJJFLO08CqosSLUsP4ICg2FVDk55IWiEmON/Sa5sZXnrY/
Z5IZO2qSu53B9YvjgYZ90SjJpZ+TRZ64OTbr8u9OfRw8ULG1huoUGtnY+vez10Sr
6JgUB0D81iFLOlGnqmSBitb+RI9OVvYfvOsuUqT/P4hK3Um+9JQG+yX/dRcf18xs
PCw6Pj7ZU7EsVBs1nFwjBqaav1Zw3x+/Jj5bScBZLPf5/Sc8r3+bJ7xIgeqd8GXc
uUt1Z6swgwvswQ1reK8oSgacLxlT9KMIlAROxlnJoAjlYs4JMY4uB9KdYx8WJyyS
YDW+9Mi1s63M2B5qoxKHmSEGl8aNNnPLHLLQ0dJ4QcPeO/ef/mwinWZV52d4QwBw
FneOejZ8vZEIGLIuQCBCIZlO538XoeDafgFYco7L7IGadTQx6qjvB7+jBE+CvUC9
lrnSALPB6c+RSi+dgzzfWbVJnzooq6AT5Cy1nBjZaSGzSbIHCSszfsDaztd5E6b+
eK/jwrSsfh1b+AmHShHOeFcW2Q+81cLt6lkUEuBD71a4/q7pv8K5b5ALDZopG8UT
QGLDwMfNcFZuH1JjU/L6bqNAid0nVT5NNFsSb3lQFv31k1DOR1m9k1yQBKBJxnf5
Id+gaMtKrzlmkPP7PsmpKrUhpjXkl0Huv5Fp4WSzPhO2fB2bdjb9RH2RAQoaqT9u
AVQjFoEztTdspJnB+wl4tATwzymYfm/DKc5RWLEKxZ7UdIXNckbscgr2J3sB3wrJ
UN1sCrfVP29UTrTYFcZDoDTJXXHyCyPNkz5imfo9psLWC7dNFf9gPSFc/JUf4xUf
H3OJDXhtqOKIuegEt4PU3Yd+Xfs3brh8+ccu19G1aw5pGkMif+gcTlE0YAXirSQS
NUh+/+TBPmwtrv4HAUg4bvpohdAsat5c/tbWxTdMKEMcyk55cPKCTGHO2VdIJSpA
xfDddqBaucanww36xxRKLnLIgPw1wXws3l1uy8AmVyAD6YvKDMIAuhBCXRZPlKTA
FnQr/TLN6Q3Y4cSu2vyvZ9eTjg03NifYNeyB+OdaJ/d2RgRn7lyeBOnqV7nDyZkA
nbz1HsG5GN6GGw64YI9s2JZlhM//n0nIyp1k8KTpsKdUrPjWF+fB9LHGIjUqCnac
RGW9ZKF8B+RnhvNAJJDXVT1r6+ykNmEO0KdU9jYCu3H6Hm5caTK6wPfNDH4BoABZ
/xPRyfV/Pr8v8qUw2jIrdn4ST3CQc1PB77SrIfIvs1gPUNN9LuBcJUpiI3mlODU5
1ZWxkMxjW23vWdw4LN9EGB3TvXuNnGplQXGxXm7fNPjLVtz+8FdEHuEObDI/9Cpc
OKNWNjprzZ3RJo4TpulaSRrrhiaDg4F+Jz2H45kmv6+SH9Mx6cn8sLL1VAWqHJvR
bNaMVNcTMTWbZ5IMwFT3TKkEl7yG0VNt3ZDUhDyPnP07njIvxLTjPM0V9Yw96SuI
eUqYnFq2g4hfKkcGVPplTxWYlgRWxg57zJD7nXOJW7lomo0XaQYkoL/517+UeN0w
FbRau0wsr3fMGj1QHKeqfsqzce7Jo99/T1xP5Qa5y8tL5ih3qUNnxysrfBk0oqAL
8fiP2XhD0FHAb4naYI2Jiqo2q9t0u6m7r5cM3VpBmBX7+u1dYjK2HGKGCVslgh/i
mg5V82DAMs6W9OsteHHtRSmc03cTA4u/hSSSLLUsnh8bi53xMZMq6O7900lLKwNK
6G0XLiHTL5Yweii7/db4sRkbQG21VSQoDmq4y0hnMESyvNmSUYLl98ukgQe9TsZj
d6GHBeerXcFBgb9dpZwkszlbwyMv25lHfNh713mSp9M5YBD6+M4uSovuKY1s4t85
nLTetUdOR4zJfGlD2NZx6EE7I0cIfw8FYQUw6R4Z75i1L2W/iFWRlWBxpLnpZzo7
QqflCHnM488E3LRl1Zj9nsZGRLCt7o4Zt41o4EShFPOQBe/cwpmerCPV3frbc3oQ
GX8Q0Mpy4wdvZ5IDmJyddGLYEI5sIgGuu/gLzy2JIjEz0mbZkbATJePwwX8stvu0
1TPB1O/3s60gTML4a6JQX48bDtlTqnGv1nA8+/oP00N7HUX09tq0TgEsVDwZeNUa
lnMlXeVkO2P/zw4C+NE5g2XwG9/AhfZNpTdf+jxCsoAVXoGV1DFeYBLy4yfBONye
fz8Dn+sls1G14bWZPe1DX18a/xWdYyX76y2btdeFBs6hi9sjv4AzbanXHYDP0GF9
gp6oe59id/EYYW+RAq+8XR11xsBeu4UUgz+2eVoVA0Blb4VCVspUfabaplobZoBb
nfgIrRegMNv9b1Al1jN9JTvkzs6XgyKvEX8CaFzbLOkcqJ3WPnPf8qtzNP9bkSFh
+rBKxYpcINxhN3K5Fh5QSkgIxIPXkgxXxRhYhCQDCHDfGsvv5LpNqwOzr61Eupce
1QgGtseord0M8nias5QC3JrlyDmBreNhXd3GXl+o+KJ+FsLS0I0UX27n2THRzVzv
b9mztDzwLHxRm65ZaWSGAwAPlKgIYNp2i3eElk4cVzHrEnjxwHkKmPzupdhOQo4n
XjsGv2p5k5n/5iy8NnjoXFoHVOpK3X1i0XzJhVdrqfCsnOcUYfguFcOYLa98hRAA
M+n/0o7OS6ZN+ximYcqp73KXUAazVBez1RWYcArNL5TUlUctebziJolNPkuxI4Mz
3qmDRTf4my1p9ZbfLnT97RHxpJybX+7+JWdZOAyKw+u9jIGoWkVcsNOXplDSL0yI
8cQ/b1NAfXqIZ2g8VYZ4ai71TivKxw9mUE99nPuTXS+j3wBnimNe4zAtUB1For/o
g8ju8ads34pgfGuRrNlKPY8CdgBK3AbE6SkSZxDocFoHxHVO18plYlzBaw9ExW6E
mP9QmYWGOL3hQ2Mq+17FcL5LnG8LC42SaVEpdfxNFBZ55z+0GT2Q2alnny08tDiJ
alixgsWyWKZj6O3OqH4UVnqSf1zJnJXk27/9wBFKNAuZpwdmxt2QwhIXuxsS7Wzf
tlNNBq2EdsLU55vWLKLxuj7HXjj6ywJuLW0eeviTGmogo1eep/xh2svnCWnY+FIa
uEefqQdkSZuBt8ErfwTUpznfz8mUfbyY/uOFjop9v3T0G11am4EfIAore3zePh23
gs+/O1aHB9tLaSrB4dLm1fzau2Hny3I8csGpCowaY0vBxnic4szkcpAgzRDzwXMO
A7UQtFt36iCp+ePcf5pUEK4HSmpV4c5Kq/5CwNvNoQGOXw9LpNwa3gmfHo/rg3CG
bZTKEergObP8sVz8O24k7Z9C8FNnTsBt09g/dxedN/IlnSiRjihnRsOnHntT78hT
dqYnvuBSzujZh34de/BmmecurBkQmAbbXbQPApA36jE8v1CBmLiPXEvBEF5l+X/H
BXAPS4xSaVU7oURTCHobgS1oWa5ANNY4pk0xKvgq/gDJX4jUz1Im4NVTLqRP/c3n
PIr9S9WqTQBPoEOq0f34d5NjJNjwZw9gAOy0G0D/bdZqScmtilldaigh2z3sSj03
RMsw/svo+Y2T1cB70h7s6wWAoUO6oL+6UHs3dDNu087oiPoRDYzjIV19KghAGq9T
F+Xky+rNnFGvqiwTcG1ubN+4W7+55BsAAtCmJyzOOTqV+0FxGoRU/xruZofbucCh
W5FS9fHRXw82slmbb86SgqvFuPX52fiOAQ2adqBQLCFW6SbVlUYYFe+4SNJ17adC
WyHckYoFyvM++oud7GH3v40TApgRzqh9AOmXXGzS5IhUTii9kRUjRYiT2gAhe0ho
g/WQCVunWMp07OiKo28OPn86a9WdAtfzzHPUh5bb3D5qMjKG7IaLQeciIxcvRJaO
qo3QGrVndTgCyhwbjhTFY0AuiWNEUXMnbXq949z6tKktNG3Lr3tZHlgMZncjzXZ4
edlnGWACh9tdk8YdcjpH2b5DzVjMMi8OnbsYDvVMriii1fkImyRHH5AsOKfEZ6Ix
LloE8YbYSwXAazV61QKwtC7njrTEI9WRIg6AYGohnqkYre/9wDRgnGUQSuFie+r5
SMhH4Xpatgb6+3i7RvwaLjk5fyJuDjdPLGmwbFZkwx3iOaQ1nR8oyTq1FRVOAHqa
O7IOxs644RMyNdAiFLsSdMoLmW43XZ476MOMdKqToHhivH3BQr93kwBD604vToOm
JdKX0cXytV0B56l0Im7nSXC+4hE/X+tE/lPxsHqam2ud3LJlzxEZXOrR2U18lfGa
SmZUu2w2ODLulVkXpyCCYnovPCqEQ18bljsLWFsVNzw0HNt11PFqoV3mX6YnitOJ
Jr9D83OCeHzsY/6qlTePe4++CFOUzoc+Y9KcwmtZEYX0PWKu3ZiiaKCbnfJKcweM
tpsiI9YK3hJN8pVystmhNB2zTKsLY3RKGCfXUh/AWN0lYIOKKqboxxgoDPbbaLeR
hLV/I1bV/8bY0GjeBM2nQIXdV/JSwW13LZHuo9nM5x/xcbk692VuZNIaehgNF26/
jW/ZayjsvZCAsYJwY0uGTmQ6S/d8rlqeIOercfXYskVGrZSdPIKB6gXwRqf7gNEo
gGgpYkOzrsSOY9iJyy658C5MOj4SdMiJ7+4FK2H8AseBpZJHxtc3U8KS0h16rcC/
QfeyiaZlrMeRltJO5X/dhXIwMvB7rGF2N9T4Nnuq+oSunp6fiyYbSfUyrhTxmoLT
23X6pfOCfgA+2I09ovE3bCJ1jbET4mRP/s5LtZfegnwPSGW4Ao1o2p4A9O3Gd53R
zCOAgk3fCKgBP5aO7YFaNBqcgNAEXqXSXk9F4zineGmzkj5UP5bSi/ULRe24kvW0
pbOqm7sQvrMPmuIePj1pF4cw6qM1mLVNrmy0rX2CA3QgOul5SdJSQFuENW+dvRZ6
1IYtCDlDWuLe4TKi0DoTGV6miWi4aJR9LrOJuYa0cyP7Y0F/+cwDxReWdnYIG9WP
BR1oSW5e8cgpRdVIYPVLJ8RL7c1nDb6utobb7cA2UFH+qiAvtc1jq53kK4cFpwFX
quXTCOUnjpCIkOJG/2JVCCuoLaU+CTPW9fvaFIIHCApLoFDfeQQgW1uAMsHw9pS5
Kf/WD0jpYZHT5StE+rh1iWZ5el5hrzTIY0EBKkQpIlLeuZ16lowyRTrwvBwBF8xY
YsSDJYrO+Zwj6V+2QBBzYnZpnOk4CXZOnqw58OK67sYf2lMYCN2fRAvMjhiGJP01
ctohSnq0IBV06rnIBWjNTPbVLJO8YeeygInl3vwZf/pCs1/5GzDo3wHCzvT2D478
XWtow2FRXbkfjfGqdmg+0xN3biBpTQzvW6UuSGqVEeXjogR0owcbIFf4qZ/0iWRa
W5uOe8rJrsLmYyT8WT1384PBnNYLu+2Pe29ke88MCN9DV2BovbWFHnH6fB1iUKYo
DOpJvIjmQ/On3z0Bvz0wO/keKQ4ttW8r/hmlye4vkEsXXTAmutSUzJKu7YtRDbuW
qgwOAEy2OB9GAexLu8Vg02GNUODiaOmWCDfcT5eFkW3botTbKGnzrPlaLJgDPW5m
H0pSqTywej9vsvPee9B7eifh4nXRyXpdlEOC3ExHM++zKIxy8jyESvMHlE/CFC0R
Tc9RJH66yNfh4SYJvWBdrzWwy6PBzy5bNwWw2ghsAU4A2PwD0OUox2fpIPZFnxZU
yK4bK6XCtYbiQx7W621oClGS+ElGVkIDBQBZK756QiOGcpiOrP/C96/JbebB0VRk
mP5e5KQMbkFIoXzYMbtZYEvmuKYm7I2R6EqboSG2eI1AL0+736vGW/J05gUloXya
z0+DhrwX+NHsvird4Sq3Q4SqXV9WJUMKJk4wXsJ9U7vRlRMN2Yf2soYmV8stCZt2
8PY8wgSrHPFnpAfwOR2QdIZzN9NlNbvfSLRuh07j28IVMUpNiO6kDkoLZHC1SxZI
MaZZk0RweoHQWw7ahx3dzMzH+MkfTBDTmK/rKa46KnGHsYcTev+ugnw9l7r+HXBs
OKAboLJS12kui3qkEGuO1NxWIzxviMDioAdymkckm17jdGPWFfuq98bzQr7zS36Z
+u3yoJUJKYaQwXYyyNkZywDAtu7OQKKhXR2Ke9p7q+MG5vntDg3WHUd9Fzs2L5Gj
1GrMfTS2MZuPQDhZ2MEhoPhe2DU5nsuyqnla+k13rIzEIUL4mA2nTrRluNA7yqoo
iSeOSpQ8NZ7alhR6xZBcAGEq9qZdGpCX77sHSH55InuyUp/Kg90i4pq4c1dtNAGd
wPYXh9XyHkgWQWossUq4syLq0ps9OmwGbuJhgBW3noAcWoa+UNA8s6PDNlVeG9jW
Up7VP+o4wgN/Frl52/jI1e8WDEWfsEOLsfeLXJDE3eR7TsyKaIIf0+g1w6vUABQf
dKHgbr2z9fCVSEdrvBgl0smjnKCf3Zur41C4kVdga43Ym5t5WsIgN2KzSRSP5Asb
xBi81aV/Sx66d3fv6HaaI1J1HLcRBOGrlzNMzVuoW1lmfzzA2OaHbansn4c8Pgy0
WW8OUXrB7+XNuMdNqp8dFrO/7mAiY/UIAGpB7WWifVjDH0RdLDzjoZT/teReJAs/
GO1lQrzVwI8oOQV6obHM8bbXEK/rLGOk39bXa5GcaBQmNDXx6dealY4EpUjsSPds
arPq5z7TjBngiMEk6yhWHmfD68k+HqHynshP37M5WP9gNfLem+gCmz7lYsZUHvil
Mrk8G41uwywygQucTj4jS4EF58du/RwFkIBU48CXikgvq3nc3rSo7H+1OGFI8ZhB
y4BZzd83oy6wsDlqnAbfGrdaER7RpycC+o8zSTvh7T361Fc51iq8xwtEnOAdhwbp
vewpKlyak0WcNURvHJFuIYdb7WZwumUeCe5nkYiPipinaq0KKnjvdwWLxKJVA2A/
ce758q/RuGC388dDKSJDRWalA+O1JzY/uYQp8S0bimqoHEWOvp5d1KmOS3nx3uxL
1m1bvTFHB2vAfp4SVRBUdgBW5YFDU2fpd2ZJI/LrjjBa8CExZWQmpOWt0nwH6AXO
/+meYZM8fOVu5J5OCyAi+BnEXGsXgs7b/XNY+G2LZotYYehboBxQDvz80v2Ms6/q
V3u01Y08ZwoqWzfRrBgaRepTCNSX6FH+znbHHb2IklcKFGfrpnUjI1Iv9/Wvsw72
9EXLUWL9KmCMg5XzC8Ac3z0IEAwnZRI+Ey10JQ0Y0id5FK6Z9ZtNyxNtMqxRfSUi
/5T9CEVgujgoN47MaNEAhCvMn//fClfenX8wAy52AOXm6nLGjJ8JcAcUoFu0obPt
dM/jFev9o3A7YKCuG5A02X7Q/45pHSTrlCscNd801GuvBcKHP6sBcXMRhWNKX+Pt
USnk/TSk0RWZb/17rLSCvsqFX3jaObAtBwcnBSmsLIB3nDX/seipR+aOuNBuajZo
WhUgeQ34dt9XKxSPo0TA/vo81gnIcO82c2pH7Lwtl6uL7f/+oZzKAzFuHYWcjzLJ
ggqfIRu+n7IcsoD4FRmUOiEQomeTgYtQih7jdPtxe29qWoNXUh5JST8ez3Czbfas
RnAEy0f9s9rx1MPEM5diZbwjr4loiiBgQGgFgPwts0Z0FqhpxLhvAfIlM+cFkM40
OMndhTFYU4Z/2UFJ8mRStZNMyEwXfiZn33hdzETS6sV3tNLAl7hRON57rdEYymPT
CR/jma18pGM/PxZuJo+zhGB1Uukv9Hf3TXU/iS+lKvZRvOaS/iFrWCQc+c0CrgHK
99NVLnw9luR+9A8hzDp5q5sJB70SBpPAL3wWSxz9HK3KkwjjIOJbjA+P5zK1spC4
7LBX3TqK0DHm5qayBPJdMLAGOYzAZdvHYfIRIIAUT6p8FLxGZ0hWe5qL2fckfK8P
jzLcVW4mKTD+jzezghTCbleHfhFWaTIhYGDJqUYJ9W779TI9q+ARZF0XsWMyJXDS
pQ0pg6CgVQFkjecThw5zhWp9uNoiSLqExesBr+bSPtQi7FtJqy8OkxN9E8YJsuFG
0bcfziWZL4FwPJE7s7gJdIg2ak0v0+rAzt1b4QbYpfb+FvNSXv0F7rROzVFWBv5Y
BuV86Om3VoVsoOLuvt1lhqguwe1AQnwPXLrhjGGDOJksnZV3ZgzIKhtNEtT7GbMh
lgbiIAVUU4/LJuT1rVtXDK0cYvWQmY9R+G4gXaIEfspP2YKDXqIr3YUWbvQKuSRP
a3QBpnNNKJxkc0/sPkrQGHX/o6ThxgP3sg+8U5RTw2vEz7UIY6qK2WYYChWq5x/T
7qbaOmEBCZwkV2/xgMLBtk00brmXt7s5vMpJZuWwGJgAoacWHNSPyYJ9aZFbZ9WT
ps8sEhVVbO6QhyRbca/OHqAbsFZbY9agkrIF5v6WckqW4CzcsLg2KImqlFNVyF/8
NqwxtNkrOnDtJonXkjdqU0WA7D/lr/8vLaTcLgJ/JpEebtB1YsfxpDjs93RQTqU5
XnKXwnn2b2+cyILnA81V6vJprZNMfz2N5qdSlUBjZRqxxPUdU63/waY1fsuS+YpM
GOU96n+HtzAq6JQylis9iCxwMtg+CHI9nx1DO35eBdFAm/Wm05xHbguOpCTTL5AT
h5dHPUbH0WGcyNMEPKcrLq+T1uSLmKTQ2hgTXZnTFSeV2ItjTAZ8vtF+YklxwX+q
pYjgVrR9SAk5VCjo+pSaWkjwD/EmDjqgPU3LWYZv26Om/en0QaFtv4xQLGTSuEsT
cJ5Bs2m2RJzQlITAm+O3MJFXVW4zPCwxfjNzCGSB6PwhwyEjGzj4Tf/5ZAJimacM
HeHUlxWfvVpTOGkotG79Pm11VgrAj74zyJ5LTVlaY/ekNZP8NCIt6GbKNH18M+Cp
EC+VpgmRJsiXPJD1Wi4G34DtW9q9s8TIKnjNi5p6HzwIedmSNarqycU6fwVz9zwE
8OZya2Gh6L+daOmRGm5G0uhZ/NAuCUG1PuoKywUCVYijbtROP4bqj40/DYXMItM4
rKxmvqw6yfANuaTWHhjrjXUNu5uz6h9rglmyGOIE3me2M0lmPndXRWep3q7VYONA
2EnOGIYMTDM61yEoF+SXzhp9IA3XgW9lAPP0Y8w2Aze4ZX3ZwQ1Xod+j7r1ZmOSo
YOhKBoToVk2yYWxV4ES9ibdhRpcG+sD3Dcc+PqQh9BWxBJqAhdToMv5lnKSmdhql
EsTAOeJhQWzWq9WekRSueVxEvuuxwaJDGJy5TXHjBm2B1bj6iyNyUtYHVOg5bEMs
aA8WSkvH3VfLbHqoxLlIuoPLl3ujb7/A0051k4isFjRy2G0dFalRcL4ENm6Oc4KG
vU/owlwrO0nystM7m/ei014Kze+tvx5JIEqB5SwyQeowU36+KU1womZHlgnGX72X
sjdUZdFzFHxtt14G4aXn8oMv/N1HkMeHwJ2rtayBTyIvxHXO6hk22LaPSdQyuB8v
DfC02iyCXIEX2m97PFEnjsY2Wajqzl8H12jXLX3J3zuJsquTfiBezaWV2DYLsM0t
9WU8+Yig0XUGFJPELUAAUwRRT1t1SnZBUIVSHtPIjNScYWUgbT8417OrlFMqJ2vZ
PVGH94j2XE+FahfVJAmulv86Kl9fOfrjBLp9/kP84REbZmpemCwpQZOaybI6OZju
XSAN4MPu9QBc8/kGWV9kceOWfydQf1XYWji0Mexj639ZsIaZATpRondL/EmHOzos
0dmRcCUK0aYiYF7yo2/pe5HQXEAk7XCW/p++tmv9BQ1et++XboUvHR7YKrTFybUc
Dl5MA47XoGgQdnLj0a7HQ9XBTvjJJhy4XOsASogwFeOJY2yR3aLMAbGfFGAq6qLp
U6HGH1hf+mSTJvFMB5jaB7QBroOKMJSEtRS/aWYM/+bljeqwg5OzZlUMvepk2lBD
WNSn1oOMbt0jelxJJCpwWvolBswCdHKSQ9RgwVC5haMAKpnjAh5JETVK8Yn/yIyI
9Nxv3WOWXvMaOzbI51g19ZPcN741/8xmW8HDeERj9vINwF3gt4MkqzbSgz9XHoHR
wjEfyRn9WDzH5+7cJS6kxm15NJIMsLpwVRDRoOCAiR6A1K2Ip488KzQ1qKsmarq0
M75I0RQ0GBvZ4TeynMzzyceRU32Yyxq2p30r4Aq2L0dPZNtX4fOkmUAb9HluNC3+
SgtG/V0SFPgPOiS3KiMhVwRveGYw8fidEqJy/FVFdS6U7N+7vTaya5cYOVC2m8eJ
fBGgLgizJ9IV8rEGNs0xzxhNNdNZBJqfyDSrBjM8nrY6jzkqR914JbFxDefjX5F0
FwdvF96Kn5/pSNAYk5l97q/mDjxkpOonEyVLbybW8vuFA0CLg4wwAK3VHTEEP9nH
eh1CJfuzRv6pbnswWMwmWX73g6ryPFgwXqdy130FBBm/gs1hhzQ69c0w6XW2RFHp
QvGRyPasj71LGmB91YmZ/8X2Yt9MN26qOrg3XRCNMsSvFtE7WVGjedVBg2hdYnU8
6srS+hKstsJjTufdVn5KKs6d0iLLSch/kkDb6T86o+kt/WRjqPVS+bDs7Bwkt0CY
rWXZcEp0WX1nidTQ95STU21Pwyd29F1qwTosZ1icRkjEjPBdEVKmMotDLKUMhFag
3aRIohyhszxq0Ni0o516I79hfZ2+UwmGiW1MzblxfXJFh8+usKlRA0p/ItG7jMdE
0ayIwYQJPEPeB8uk5eczcL2w7pILzWXiAaUJ54y2+7CvwUa0F3pHDeUq20JS4RDA
rMKWb5d+X9rsmuUSowb6hqWzPfYkllJFb83uKgKrNTcn7StjSYN85mTi3Qv7yTB7
Nq9QYEEo6704o4xLwKlfMJPuK4OpZ8fNC3HaI61rFZAzWuIIFUiHNWR1mYa6rQWZ
qgt0Pe0S2/QQUNlHT1VVpgxJuelFeJINtWA/4ONzgXjyP7oyA7AG0Qg+4Dn83s0z
ZMMJzyfFZ0lOzzLHNSqI+IQ5I2poUcx1QpR7R7Dbd2EsE4fDByNnx7T8M8HvIdjA
N5DVljdvChJoBb0DLILwi4qmdBSJ1OuhMVYoTSUsLaPS1+RxV2p4+OLoO/dknWjc
LECpIGX93Mfto2+YMq4Fc2EP02rXAZqdVH852yhqtxpV2mTqfFajF7+3SYb34Lmz
/dFM2rbVtjaXUgnPPjp0H15k+JXDgE1BBAfHbzK7uTS1ecfnwiqrVAeqc5fxoTZv
k6aG1arUQnwWJpmgf/PySe3jNy8V/xUYA07bshpBgP5v4tSWMHFQaI3oq5rKr9Nx
yoei/pQyEnn3nPlnLg0b8V5V0ibuRq4lFrZWZ5bxRlDcVdNoaDDH5v8/DKAiEObw
4pG9j086NDG/KlcFEOKylKKYs0E4V19kM8ugRjwKX8a+WkTIVWf5baS/Si9KFLPs
7qbpi1gH1F4rpxhVPV1hFCFMIstCe9IfTzsKJnv81kO2zZxjp87Jzy5v3RJgTFcZ
4t0RYqQx2SAA1Nhw5LKByV6v9MaavhukbVMzg4bY9gfiFSAO8WqrRuu1DKYARbG3
StG6uVQjFtarr47p543iReV0oQ6ah4CtbmE1b7Ng0+TbgalT5TWkSCp/Xth6FC4j
n38ISOXiMEDu567bWfXpPlyb8HAjXoIAefxh+LzJdPRXQZYepw9Wqj3PGKWKDltw
pNEe5NoS7+0rLrNmcICMjY1Km2hvKKYDzwHiSfVjuXQlix28hYkybr9rDivuiYTq
KCsTdezDmkr/rXD69dg5bPmq1nVI9vG0Uq0jW76DDVPpYC6Q5Hgl1bOjmZZZ+Dqp
Y6UDK9u99/tUTQ1Ut7eifAIHxB1W7rZRJgdYllG2vZDPvEFS/K1pQZPG1aGVLk+Y
wtxDETPlOqTcsGtQNuLknSQSxyUx0n0saBhIjIi9lm/co48qUXnipVWc75RF6NqF
+4ZvWPuktBG58//rrl3F/YeA23zs/RpFRmUba84wGuKSCBWmypYhs3J4lTF3wItW
uQ4BCPiUGHN/esOIYYJPHYSFF3jxXMcmL2G4mT8b9bLcNNsTFMdR69+V1sZvO2v1
uT14ESA8G+2gjhimF+A3xgsMCJPkIfakD17EI6bBVXvlj1mDJ7atquGPnWJ+myq0
+quNeWIiGtkjK5JTAz8MVJB2AGhcx/rm4fyMG3GURjlfy/g7WyEzoNIhjzQ/bXJP
diHzRmiDNPEhjklan658XRpQ9Cexi7xil3F3eVpTKZCjaf05nhRSVCuKVdtRc+xU
hLoy/WVt0hfG6CF4SYmwTMKaNb9g1CScSbedYRosROayQ3u0EArgQ4UEl+tOm4gn
0RwozaK4sgzkkUp9FFr1/aoGZvWn+kPgAqJMWlkbepa0ouI8wXIw8T+AuCr/lmdP
XzeMRcYqS105i6UJAVOyabd9hN4pE76CkXTjkcdd7mkHfcwU23Ur92QPTMDf9gxg
P2P1bRCEPTg4n+nMqYSDMaK3yGcRepbjgu2gW5dDqMF0ZFYq/C0jGHqI8svxssSp
h+in6VRtCmJ8E7PUwA1NKtRCy02bS1sxARQP3PAaKWWCf3uCWvOqRgczIGzbMGE6
ozm9CIG5LbdnMOCOVM+bSQaLRCnznAugHu7ndZJyHjNARbkZG389Coi9wiuGhgK/
O8hD9/rg468Yyx4FCKhwPXEsHZ0qiYlDTQTyOID04gSa2YlkpewsExc5lNRrgdlS
+PJjrV44aY6DDjBMDPfrhmvF0jIxNGdRxJMhEF02EQAPVL1pU4zi2uOoiJTDE1l2
MxZMXMbRBbcR+1n9AcyvQgsKGKgBmATB/JbUFLwMsgbWSDP0d34UAN42oUXM4zhQ
MwjgZdedrP54DJcFfqRN8cHKh6oyHi/jh6XyC/NUnbhxT2TC4epA/P9rExd55qN+
X3Jyrikc9rH/wPqEYI73XusIm6V6JEIuH3l87EADyQHng6zX+cjhDa51j7NUx79M
7c+geBjTvb02enToSD45j7Z5l3sZYb909DlUKrqcPz7YqjlvHRNcGm4RNn+13Jvv
8x201vPT95/xSSTtc8BGh0Wbt1irkUOS1MXLnGSUfqah37f5gNzgy76gocTYsSyY
iV9TC8bc3WQzVpkJeY71QnepAKOuNPJ0d19BP1Y6BWTI5uoiFMqdPUUuYrvjpAxI
V19Voe26htiG0JnmWtFwIhBIRupx6WN2LHWiU3tR5eV2xyx9mBFDLhg79q+B7eB/
LbQZRQ/8ORgtdOPLevDoBgDfSNwrG8f8mYgdVBdTXhgPYcS5k8WLR5YC5v05RFkT
7HIjqMKUU5jDlcAfBWvvG2nGciFdLn/1+fOS1FreBhQN1UylSKGchziEMuYpxgId
Qs9MSpmtEwalunPGfaKqwTWA9kdKLnhsY9IhK2j7sL2SOPcR7SU4aUbFleNPKnkK
ECZWE3fRN4Awc4MK5LUW9IGr1NPOQt7jMrQMQ54zwemw2xzuD4rHWUbWgDMGOED9
BW7lFcERpQzcvFu3xSnTuJEu+BEo48kIRDC5I6tbuuRGezCuuO6YhBFYjIB/uyYI
UJijHWcuMmYh1naCRb+uCZfljXUPl3ALCKJMj1yOJG2+cMSXvjz5B+KRfQyWZSev
6PL3frvbUxAI3Y0sxxiF6/a5feJxEFpyd3OnoHM1Zb/BHMkjye5OX6VyMRanQXub
p+XjOSi46eyjIy4iIlj/KCGulfVUfO+KeB5kDJ0Cwx2GO813HoM4HiZAnYWoEJO9
Cjvrpi/87HCJnJpKMv3Dha5slYpWbrMWtOt1VofmrNexTM7aRsQC8gASmZmFZtmA
CLSZAvwiXQfinWCYBNRGA5Jz4sstqGJ+Uk7TTGwwtDogWjwpntriFt4HcYxJ5TYp
DeN9kB+X9s1O/q9AOEB9ygMLbRDOyEs+Mw9K5SbG8JYYaUxDqXfsxoGBDTomJAWs
aDkupHpkdfrIgkSmFyoP5Kn4+t4vj0dp+BhT3hjFSOSIfdpWw8o5iqrF3/FsoTdB
NLd5RaytmkRYyLCg/BHpQPRGkFYtYJ0lW73BH3kDMi7oiwnBUlBhkmxRaDf7XybF
BXg2g6FWf5il8A4TOumvLZVEbmP0HPHKv6aFjHyN487d+6TPiJIvPzIN5FDQ+bii
aZgYvFnzFWl4/0RggFvb8YER8ri+RSBWAv/t6zfD3Wf63c1/9HNBEr1luIEqaEFp
S45qmDZNiSdeL1ArCdSoPWMvT106knN5zh+VWvXFxV6RgWnkth/DKz3Gw+U/9s4d
wtm8aPP2G09XvbCkYVRF8/awa9Zp4td4geVRtIfSzxb8oF9bc1jvDuhVjsWzBbfa
NBwin+lAdqaZDYH8mGTR3iPX2AoyyqDS+LT+RsOLmHICQFdY7vBwyXq/wgHJ1k6y
mD44o5fCMWjX6k+LTOrLLvQqXpUk8WE1s5PXEb9YteJnDf61wcpPRlb5X89v7nuH
97YUwoRU6qYy8B+8Iu9AJZDmxhL1yr3Er3ENlHXrzV4zW4kIFG1IjiZoAfd+9e7Q
aQ8cylKR5H4BVeeNHZospZTiDqiyq0L/JdJ/gqyrvKQ1rF+ARqpjOTGcDKBcjud4
hsVSAkTVWRPqI/7udDsdsknqNNMgHB/NYuykYRyFyEWz4gAG4yXm/5UMOjlZhtZN
FVzhUMpGZOvltkpoJCHYhN2ppMtKCXmFFjNKP++aMI40/00Wgolw/0e0n7aFxFjh
aSGNdICZDHk0VLOfFbj0qLJlxmcBuXQbzBH4qpY+3XiALTlyCgoa39kyFvmCCFhN
ewZxphDWTZChE4Hzmuv2m7fcdekSzbisO516cgYCcIFGqKu0uxUZ8p2JjyV2JFYF
4EGji6K9hvikYtQjAr+AJv1EzO5eLjV+0f+ImhIhZngGAaf2gwLsaodCvpkhroTM
sL9uw46njv86vOedKO+HypzzIrGlHSRTO8kBS1N2Yfhe+Mk3v3weupVFgGBfKBtg
DF6NDmHm/7rstDQkFIzUu56OQnjaVruio2UNOoXm2mep701CtoZRMq4MQWbffbNn
7yY2P899aox6OtvWzQMTMo0y3UUFwlQ/m8CcgN4u5CPiJIFoP51H8d7CwtXZg04N
0UeMoulYAGgHJngFnweyNgye9d2/wPIKZO+85KVS/APBvfP3vh7jLOsXUjFo6NEu
VhJlUNRxR2vhTVVehbXVcR9cMVkNtnLGthsJsGD9f53AG6c6kOj+SX7hJbbASk93
0NQRdejfNJ9Gf6LyyVaOMSMEopwjNnPefOepFUxWsOjySK67xn0jsDOTDRdKuQXK
ISgGNBlI+RVU/tMQMgeFZW0o9CY3ZC7FUK4+CZ9FWNGrnXlhQjCvXKo3Y5FRv4Jp
syZgNuMVn+vF+e73a4tktXuou0WxMP06H5zXAJdudW0S5xX/0Pfh0SFPQLrQpAB1
+ZgcrxhjZJR4KR+f1ew1nYUADQGA4ykutEgQa0Kb3mSV7Mn+AAA2GbPNij4bqvI2
CE6xZ9W58oXnNO4PTXMd7G00rpfAubH6CnSeZ23OsE/sFy8RVhJ0tawZeP/5YsTp
eMaCoCeLznujQVt3ZFR/XfWqhy/Dk8q8r4m9pPhyftqz2zTTcA2+wwNHmYO6j/dk
7yTaWF7Go7s6KV/hWoAr0fjmeI9ZrYbbWruczXsxPjo+WIIQu8TZQjpruhd4wGFR
8yrKFJiSmyQ8437SkvZLUZOLOMkIn2EF7yBzooOD3vpEx7BxtXeXPWwqkm40KNOU
epRjqwvhq65pQ4RjSxYXbrd+d+i3EreQzjAt5tVskNBbZL7cbbpRP/BhtKVVgvJq
UY9DnPv83fE/8naot4Hj0KI+aAXoiZI2oYZ8IjOClXZ7Aa0auvRZoMPgkR3XOVRh
UZ0bOLvM7I9hEmBBvfiP+1KjZQxdMWEzgRWOtvvzlZRlDetgk/mpjn2gQ6peCoGX
9FxVa/jnQETiIDFSH+oiCavNvtwyHEL8CBzVG60tXjwNsFO1x5P1F63GSwb3gqYt
uJ/EmXCwmeSlyMRaeWYGCECNjunk0+7MhVV+CUvH5E6MwgcFI35XWP48RawfjtX3
IETwWSKpVvRVXA4KUGQrPPpMZckSdP48KJ1fcWjh0CjugzCmUVxS0rQ5lW+KtYqH
kMnz2AceYFxqCHPTRLjxWbee9TGsqTypImUXfcHXjidIybXP71S23gtiC4HcqUAP
3rWyMj3Lx7318QqTEwMcZh0PHXp/HWvChtflAkolM/9KMc7C2TwKtF6mMS1PMHh5
91ZYfoRkWjm3jy9Y1TTPnwL3jgFRcfB7/jOA50HoiPHQ3taJZ7nABjvjkCDGCMNx
/Jc8YZKiBIipat123eUQaUQSbI6Eosl2kcy32r4XZVEkgK30zx+slQdU9rDv4y9u
/rZiIcApjW9QKCJToQ2WKJMFmhIcAA1m4adkjvU0lUyxT2NhGU/EQNmMncYeD2xz
6QKdaA4zenMnbdFBwOKE3Ys83F+y9P7bOSyuyrxwWXApS3C8v5Ydm5GWZ8+X7aT6
/FQ/caI3gYzFbpX1bcn9FSdEGA7WIWyYMi3AwfV3v5DVmZL9uD1NzCtQPXNA+jj3
1pbRfxs3xKZ3CJeWiUGuu/uHFF9KlsUIJC77YRhwIiAoWQxggPZkjvzoZZaAzIAi
yAtlhRcIVafeJDTMuW6W0pVX9A16XYAKUgzYiCyAZ9pl8bkpLrU6MlkYSBrS7UlW
pKeluFQkmipshvjn313A+1LSixSY48EyfiTffmKM8jzleuXNaiYZ0T1HZScu06D1
X+O333kfmB/pCc0wrg8iBoRMlJFWGN9FCOVNY++IWWm81P/Eju44cRHosdI/z+i8
GGnRW+kN0LxMUtk9uZB59MQdzLZW9VtTyWIdfptgz4cLizHCjNRwFqfVpzb/H7OG
Ivj7KNU7EBpbmDmHbGdASmkwctHWGbmEyyUP2j0T0uAeCrZSlaeG5iTZeUB382r3
nFzgo3fZ8ojxNuZNyKb0JI1632NBb61ha+TBcORjBOTsnHzQ3c1bvFJ8RKxxFGGw
hEKycNx6K4OU5jB9yOe6tcust88IFBq/DGnQG2z6dFbrMObByx/p2i0EOCxLWLUz
m53AZUXQ1ALN2s8HKoK2evAUqiwj/FUAthgh+OQIa/qxU8nQK6spwtuHAW8wz1EF
gwsCnF+OVUWh8M8hXOhPKrE+vN18tEw7OtTgUpJ76bPMFkKngFZRT9LzlW2ctLvw
ur8Y4HRuhMD0pW8EYmKCnkZifGj3DV1R248H5xOZ99EDiZVgWUhPiGjmRIqvvDNl
SliPHePNebWctiW3y8SDUsQUoNK6alB5YQeqqEnXkLe6GiSe5Zz+cuRgzNkCj0vD
vF8ehoAlWvm3iCMcVjmoaeSoOGCu2uv6DSPH6Ij8+oG4Er3VaYennK2DDR8drkDo
3GXiHf/+AZMxOfav2C7vgNt47hIuHLSGnEyYJ8hnwrGxmTrGX6mFa0uv29u971M5
t3SZmVO3YTwEpho8q6nS1sUfthdKBM9p+ZT5HBLaS/SGAcqBhRoMj12CU//EMKxp
mMEpcytRKp6HyA/ucijQc3Tgc+fMVDqk/FN+8+/yQaS4AhqEyH4fKQ9UJRaGlWBW
g0Ovhc0q3V7k9uKUNkOg9WwJ6PgPm1UF91qATbBOJyDOA75tqgvxBFczDUhc5QRJ
y4RxuACmym5v/J4ENpgy9GnK4TtfWSzKlOFVkE8nvEwcM4mrHGbsGZQ/Ymp9PE9F
JHBNXuzHflb8NZ/eSXtZDPA0b9blVzmIRp1l61ke7mAyBlvDHaHwM2rmRv1l7JG+
eh6eg6aU/lGom/hHcbZ9//2hJQoPDwTsJU/NHBD7HAZzUKpo2kN8QkhTOOoU67IS
eHWchGGhY5jV0AhnPvrRJVB5oW9VwMeT/4mYmP8uzyIObsTA1m5UIzhqilLcmzbl
MQ5H03hO6Z2T3bFSQ3j9MlGkrddrldteQyfeYLSlJU7opaDclqJEOwbqj4GocfHu
tMy39ZU6k8GPY4A99ZTHnrO8T0FO+Mb6WUTR5vG4EEQznVO2Mr59v3v3LzfjPDLO
EkF3Vprc2s+gLE7JOEXdIEQAd2jAKWW3QckZxQSvihdV7pf0GttROK6ZwWjVe1x+
ooIpJZ9gWrEsVM4EGAnSuMg9EutdkTXa/0JaIycyOy/D8Jk8uCTBarBxOS0g5yMv
0uYfWGU62YI/81ZaV5E9Eop1mpW80iWYy9zIDLiaX6VDaEOUUOTmyesDEzteNigd
Nb+iBpl4AagNsoe7iSBKhioOZUfRrZfqK8renY46BaEuGhS+fDH9tD0Dgv/T4lXg
Tf4d1VsiW6fWQbnOD1LE/S2PHxhCNqBFKlosA7uYp2oqfYxrPAfhtUFDUjNPrJom
sNGlCII7pmO4b1yQe3IEoL8IfZlWSjkcW2AbDhBDQ0gtIqmp89TwB6YdFIOMmAwo
mpteaBL4QGxZqm7DmYdbJU4LZz42V0pgQyoyvQ4esxmf7BtLDHArSTZyvU48Y95G
1VSqR9DFe/40of5CBcUemKjd7uXj5N4Kod2pWd7RgK3IW33WWpNALXzbHm+lEVlK
FemCdX7pkDi0L/ORmDGamIEcJ/F6R5OWSN2awQ7zhlmnKGvAGIjSbo/BVOR32ik6
JcaXwvm2+3N0B2RpA9UE4CpbioR0bjiAJttVKVxj3V5I911ikXzpDBiF4oZ+wc2B
75ZhvQclkTeviPgfmw7dExvB51IrPYEJB/PB9NR/PNBAyDEDe7v+KJtdhyE2IsJU
RzemjWxwY/FWRPTMhBCV9UZwt/NPLbRQzE0GpIzOAXLOy/5amQGFAiCbXucokXhe
shLq9sGtIkTWvuU4OgzjzEof3SlGl+AoGTnP0s7d1hR+EcEWWJS25vGYvd8aAeVR
VEX/6Q0i1IbWOHyJB+kklfscbuAFa8wBbNZRQPh16P3XIe/97Ate/hxBcutcHc80
uzPdKaacn3L8Wu6i+v2T/xOkUHfCMl/G9c7c248s6W91KMeMwgqZbaoEg1bFI5+S
YGe8wP7FFHTURmkPS3F0G812gvEnTKHNkf3MtDOSq7akovK/UZxhcxwK9T0ZS9ds
xXePiWzhvhQnIG4TxLeE6nOcE8ACLBQXMO/mDCW39o7MW6B8VuEe3jlKdbEzf+ps
f2MesDFCsvI+xXzEI1BYrzckNekJYSBhD4YjAk8s0jk5Tm7lDFPSHJ1dWN9XpaU2
a4pe9Nlbi6Z053lOTAohVQ7BJR1Czs/1UDi2I3/ZzlQRRqnLWxtFquxAExxGVsEO
uF0FUAK2u887jSO85DLWNYgtib+oc8ElQOS7KUib64PNb2un71YroOtfkmbaEkYS
Gg+WE+xukHOsygsb2vdJhUHhSq5kbe6F9SLHJDLvCbdgN2PB+9CmkQXhxkyfnaot
i28Tfu2W0x9m7cNDjrCtkg2NI1gSnTPRz3vHJecQ53cEbHNsFjaHLiqYI9DDX+ix
9gavvrk5JaBJJsCJOBjONeX/HgnjrcsgLRcGlVm0vwAieJW6Bto6OpDJtv6fEfKR
IoBGGiwRu6D22GCnbCDCWH7HSHSRm6TV0NXk9bndLNwiObOfoW4t6aLiqIQ3/o/m
E1fgcC9OFXZxOjrqPB3IAlDRQ78+lWR6sAE5DXCEBBGMUMgxwyqdBiodzTCyAndJ
YjE7zyvMnm80ZELb7oZIRRrcyhtfmPEZdIDMRVNFkUen5tIj+ujS7v9RTlrNLii3
npN3QN2KQf/qTfX9N1eT+bQ7lZKWjYN057Q8lc8T5qqq0i6i6y6GR6gYm2MrlEVt
zOO+iHQzekAKRvU95XLHQy/IPR7XwZhKo+u3AKINKbXj12lFOZRuugb8X9ayaJAb
++z0Jb2+R3Ue5WVMVRLST/spBcATl/SKJkGcipvdugdumk7X9WqXY96U6B3ESql8
Z+Cc70dvm+cpkVqDJWOGpSI71VPNbg8KegDUsaRL949f6e1sRfU7zfDLOvke8hgq
flbSzb3MFPwrfmmU7tnfu7REwow8VRcy4Fqo8nUuDvOG8YImUDhg9RrDBqZowXaS
PcJ7wMS/aNLEEQI6/6bFmcn+HVRWrgBQvxdw2/dB2Sv2vqhyLf3WZpsulWx8/mNC
hss4fnRMFgZrpBloSVSoUsx3pe+XZ7eNqRLOhj9YCWEAxYBJzxhqXgllQJc6ZARK
E0LM11yjd/bkGYfKprGgfRxtVc+OObTFRuhWi9UDdZMejCAAQ/6yO6VWAeBNQ9qi
wk8DRHw1c67Y5IjLpTx9jIPgnuaqxPdaklzFlLdACvk+D23wtc9Cfa3gccOoYOlj
ZC5a64GXx/0l0KPIEFyXkDJdipYciUcKRRbLbv1RSgbYzpm5Ija7I/tMh9avNvQT
MSCF/M2qWYhuxvNP06OFvM/Q52U0fLW3igslu0amStVH2Fw68fgJKouqR9Pe70lk
vYaPjdzhRnlN2685O9zABOFLu2muONLG6cXmMdEgCnJw3CGbE3qO54InC9agAyjx
3hEnxG+DnFrNh0XOptRxoz1JzqD/Kpzk2FO8CKMB4qowtgV3GnLwuuYNPGdMA5FM
yQkxioC0dxVb4NiTOpo0MOLjOnWM90Ul7qN7TZ9KX4r6tW2nvKfcjtX+U1v38tjc
P5Wk2r05Mb/1ei7vpCEgMUBRM8He6ct+h6AJa5PAtA5aRbwotLhX+OtSidLIRH3v
eR+me1t3yo7XEizmhmz57ld9ELys8b/ezninse95E9LRZKEG6Lj9kJRW6dWUL5pW
3YcW+2985E+nYAs+RQhayoiqy+ZOsDxg01UJT7vfcMyG6/+SIUQlj0tMYHW06e4W
FVwVDz1Llx65CqSuvon8rq+FD20zJi+/9FeBsR3qJHqcHOpMXT5F3GI0xfK/KpsM
STCgJO8pHvBwaFTSfWvMDliE/YMcJQwLB7OTGberdNy2YhScG4SkkrgVUma/PEQf
sjO4QwDEqUSbC7PY8kSexk7cCg8c8E3lt+el3BCGMd6WDYvOluiFBImYhRzm/g0d
K5YV6EI42Qdc0yuoO8brt7nIECPqlcSYNlA5bPDgG/Um4rmDzqbGaEQ8/+J4pCZZ
bzC0pbhPMIQesC4h2HrayUfx8x5iy9Aoz+EqkOk2GGdJAueLSnn+HNExNaOCHT6H
p6lLqCRlB6MgPb77Xnd92smJt/VNpEV8haPwOawX6cEax157+oZatK2RgivYHjOR
6iiz5NxyVXBbwKm6vvy57hLewmQ09KbliBo3VIy85sms03bdsquxaqFVk1YWTAqD
so0vA2h2IyjY6R01wH0+0mWXntY9QULCP5F76DI2D4njXhcLeSmZ4wLto3k1FLMB
udY1Xe8zWfcRsrdMNr8ccoCSN1aDyTmNam1ZOKfjGPRj1hYJcRpmPPi19I+TRQte
+X7tpBNqcYGSkFF2y6ZRKTdQTkgxBZOTSXkA5/vELEvN0RtDz5wNoqXrqLhCzgAh
T1c9uLsVGYJfH93sEfpS+wGqHXGv/N4Zh58R04D2xAA5KNLQ5is7kyqZdxq+yJRz
jMmsNY+tcoECJAd8KFWiKQwNfube3Ud6r62n/UQOPHaWoS2gAFPXzoYYjWSL2spU
PHO+K/Wdc5PLCaalzAKyAj7htQjTDc/ywNGHCO5Zki23bPPa2nH+tVAv99ShKLhT
/LphDvzZ6NDs56TiA9ebj0JDZmlF0DvI2dlXLHgIQ7wgeUtw7+8JlVMHZOMHh1AS
OylE+IFPD9ge/2V/66xHp7UK4agKDQv78vsLH5+VzEenoO/hIsq36mk6zSf/n0C8
3WPN2aRq6k4JOpGZGzXQzq09wfLVNFPaiUdAPh2/x9atTeRHpF745p4phWR9Zi99
L8jq3569iKKcuSOfjyJ3iBwYKgYbe8M1zhjnebODP2dWBeG5y8Z2nUPWbcO/JyOm
GY5FsllQp4uwFziI3ZbyGa+oT2n1CEzmhgfM1/ZFEgt78SBXv0rz0pQaS2G9oFHB
rOzyk75ySaH++Aavp8qp1jf0gN3cL8RFKvnE7wel2FP+fB4ExdqL8hVcZw/ouc9x
+Tv/xpUKQdm7RsZJVXhbf4w7EykVnw+9PSFYPFiPMj2JTh+5md83XKIjPhR39sCE
k6jiCO8Uv66K9NiFyxafyuGpEAgzLbzrqTsPNY+sBE7h2ODKmrl46gLSpaSp8SQ6
9EwHbnAU14HAFY0fOK6/5LgnKcNl7b7roq9R7F5/2sUclHxu0o6SXx5RyEOSbMfi
5dIBDneDKfK9dp6A7yoevaotQqj3/pb07l0rgLfNqscIOmm6um/DlCihUv/yBXQt
Cx91GVEch6duVnWO/WnY/hyCWNZG1ODdwsYv4qNTZotE+LdgtpafKtmpM+O+UUiv
izu9IIj7jDX7LMAA1Q+7WvHjHZhnegomOpUbm0M/kAoUGRA3mdy3CVnsmaLTveao
CPnBF0oZSj2gJ33FYSHJ9jDvpHYCTh2D90EeCLwStSK7JjK27gEWbbd8iamWY5QA
ESUPs4F6QgTzi5TFsVvBCuXzTBUa4MYP7D6Nsp7RXWpZjiKV3qwEMqQP+gXUMoV7
X6iYdNzqpRradqbn9TtXYfmT+RO8Js0/UWd3F9/4tBNYa1MAvCCvQfPqnNGEQgGu
3DqxHd7Vi8rg1hNqeaOyy8Jccs6mrP+LaOPSQrmwPSG5m0uSmq/dgBgzz0qsk81b
ixRGz6UloyE8I5nKF4RS4Is+qRTk9ljVnY3+AVYbYvR/HjV3h6qudYmPwgDLq76z
tEsgDdX+kLLnvxI2syJpVkrY7UZZ0N9TOWj95Ivq7gMKSg4cHAQFsAK5Y5JJktFL
JuHaHfTRj/BkHD9y+Z3bsB0USHFtmpZjKSLbnq769eK7SYFLiwARM4nYBqoDuHpa
8s4RLJa4Gl4GwYFEs1P2MaRMQlGgep6K46K4pkBh2N6Am6tFDikGTuMQJGmTpPPj
xZr3FIFtmThOQEKmjPNHdUhHAYXwKWOqnTSy31Vmu15FY7mQ/iemgGJuL6nGJNmm
pnK2fvjnM2LQIOm8r9uX6oWZsu+9ZihqsoBJHxUXXwhKZEbx1fRjHigcie0sD4N2
JdPcG8LQel8zUO8pODCUo6/Y7lXt2f1ZAy0aLDGzfiqcge/xcnps0aj0WKRntzdI
SPBOqZ4hYl8X6J6fvDfXDXusK4DN6lWKlj2n+anCJ4dATehBcbMmedBfrgjgSHak
7IpZOrvmtIXzmO5S5hvlBBWrMi5wZa/2vTPMTuOTf16ya8eCt/phs2h4VZoj4uyu
vSTJ+9HlOosqPiC6kJsTKUChvRoj/dU4FYXTXX1cuO5ZiumspU7UqFwY6SFaCVRB
tqlRBc7eH3gsqqwXpc1dnMERSjBCeXMKi/yLv8IQOMw5h4vWgLV3LnsskcAZf6gq
G570vR2digCULJ80CdQDMNTSVEX2b/2OFPt6TAczTZ1hVkk72doW874h1nvmD+X+
YJwchskc+vjICRQeY+O20qB2dVcvVL9hilr7gnqmGIP+jwuAUuNle7LQR285kgfT
5eETe36N0IsrMyxdPUjwcv6y6Iwj8EVAp890Aq9K/1nlLdu8nxjVNRxFKmqobAfT
9pTtxFQXC318AEG/jw0Hf7AkT1TbNfrDKVOLML6ca+xwYN0TqnOZYlHVUEDctX14
3v6nMquPeGb59u+awhjs1ALGTXUA9pfrMUQ4VZqraiAmFqjxbix4V+gxzPWDpZAw
Xu9R37cLgqY+nudVRKC+7/ar/XcuQhzEOv9HampDfazH1eNzvLoMgwSY5EYa5uEi
aoa6MFSjt2ByC8ajB1BV8VapE4s/M5k5EUZvZYuFQKUYFqZrmj6oxBUZGpcdg0/F
AtpzAquLDGOKdyf+gDwRcpHG3doRVBxw2PjI8/qc+V2Mi5My+3z+cCRYPuCDgtC8
B1MVSwJiHRRQFULSYmx+lv98T/ItGN5T2Vs9BmiYB3D/80KRHKeXJ6cqdODWhf87
7IxNj8d7BNASAbmfHj5aaQO/ZFYTaKRHaW5+wJL9VrzYuhO1if+ooWqFeBRHz4RP
nieJxvLzfbfgHXwPxKs1bL4Et96WI606rwDajsfvHgpghJ+0zpq0TQSfeG1pQdoq
VBaCluI0V1k/6WNRphmVDLeZWImB4D4mXZ48UTnBGQOod0ladBQlTydnKVW1u2zn
8azEX4IhybgNDv6NTl7UiQKsybW4MLi9h5eHXq1XpMLS92IYEfFzGdP2C+gQYw6P
X8s2pyLqGdHFMrpb/+3MSNcO4GF3vd0pYTa+3K+Sjce3nhOu41fgo7ajGZ2jIQaQ
MDLNV3c8OCRx8CRbOAuMzOzjfEMGP2XZOQpT8PhvlCbVmB4LMCOfVi3zfMN7c2/L
90/R6X3wIv9RfSk7DeWXngfVn79yQloCHQv5LesKFywJxy/MfO5K0HHUyhkRRK6Q
eqXbgGKB2ZI9do1Ewmv82QzgMTUt/hRs4G38SQQw4h19o/YiA0I5bY/nblq+I4dZ
7cdh09KrdXRfFrpcyAzZJF/RJHwtjSQXLWX8pvclrQE5eoSQrd4OEKHo1t8rijK8
m/Tejr7AcDPuX+3oOC614G2sb12NWLO90DB8lMs2huRNl0KcHPVjlO+IN9sOswyq
wTCBSWrIf9XOejzch72D6tK+mQX7k0M3oVDnS4InwWGgX8BiZTYJRyv+rVTaOWM0
7n1dbkkgjhVT+MVpxkV3d+6ayC5+dZ8/RvN4cHKOz5MWAY6eFL0CS9LJTyX6t6l1
N7pcX0gBmMaAlRCS2eN2+82Vb+Mungm3zb3VhUIgT/SekiaxXa/Eedh0JNxsRl1i
5VC8TH95mjtFzQ5Zvj6Bh06fa5dasU7GN0vKObX2l2QvSMpRJ7smaF2YNHg+1K9I
ep3kdMYZ9MF9KLtkU1wVijrsQRwnxSUnODxOP7chgStUVT/WkRPWXFCzcHiU6ZjH
wTgcssQg4nIH1gyQDu0MEvEvrHbaNjSPgKwmSdzl+NdGLH8lG5g7nhT9daxwOn95
WFT3RR8ASK2LToUUj6t+ZwaYgHv+4LiAIWu78AeaKKmZ3Tl8tK1CC+EPfB6uFIGw
rXnFdwG44eWmsyLsb7c8M7nwGsLszqXEnFu36y1A9MOkxHutG4+tySSlPflU7qiw
+Lz8vouykQFd/jnq2dp2YsJZhB0r+5IESFvRQGkzmCATg9pPDwoGo+KF4F9JggUs
EXaX0FvYFoIme2AmFrGLVJkLSkVOKurAxc883MyenpcuZVioPRnorllYbV3EaFO6
ARONmki2SO+9caY2WwOgFuYPvVoIXLHF6SAPZC8vRqCpjN0cA/hCZmMJaxCCYOor
9Hha2DYg1YPf3b3tAmRQxzzbWy4IpnGqETkTPWqJk6XNOI+l6QxLZEd6uWn0Lu7R
CZzx5Zx9e6NxyLWaW3vibqlytlFXR3j57yJcu4NTCkzAxHk+IdQElCKdzRkOSXoz
sWsLSRVmWHWJYFDvoe4nDvv5lYMW0zem7jt9I6s+bhhh276rPOY2T50zG6BfHuEa
kIUcbZZ+fVdgg90HN5R24I5MU5AQg4LqJm4LeQNesMirLncLNtUnZxOyzHeUWX0p
Ika4eYKL3Vd0/SjzNghYckZrOZXQDD1Izetu1wOkzZ5r7tOVYvrpNoseZ7ZHwDhj
rERKznYDQOE/lHstEKMQX7IvKNqayAcdINiLcJex85JZWCBE1t5jDrtWwIDENaCX
WLhS80UxrQEKK5tQj7w+IWm78WwkJlzjuWipDOwLhVopG+C2hWGuR4efv8Gi5Jqn
JivTskyTDEG78G2U3lP6N8YQKkfVhTl3yDtONw9NsMNHJSt4EXvfWbpGaYNwO/IY
FVjQB6y0/diItqhc7abV4zI/p2Iy8TqHgoSUxjy0kNImLRuNhjskrM2F9tQ7BLC9
+HZnBQs+3XDl2o7uMo7rJ7rrn0+bTRLIE+vFZgSdijwSmHSnPUzH0CUZyanQbU1n
xjHNbwmyCWr48zFKuHre3OsUzqfHvdDLXbfc4jLTG9NOqK64/5d35NZibZtOlnVi
YzjVgDsDvjoS1NFEYOkS63IS+dC7TucTnwkKLabFkc864xz96bfJHm/pVCoZgVta
Abj3VrLeHYlGMJyxC6rubLMzgDOHnW1OeG563bxQ8MDmaK7PITOlV3mhU3t3CjZg
mNGTvjhGvzyPQI0P9UcTukOOaMFfy+5flwDMZNl5N8zG+XgKcJ/im0FkBoxgS8v5
psgA1GH/vgCiW2GsG0+/PDzJsDIMohSWfSfjfHUf9oko0angLu93XiIvIMP7hSJY
BFrLQO2d1dl/REvRpZYKR7EgwnT7ss4cmnF3Td1Z9i79558+Cfr9i8cAyRAagz2t
lkBKi7M8EgL2y0HmhxRuh1L4o0pwYkn7IqghRCDA2tSF1xXnvX7KPQjxQJ4tMHZX
/7LicHEQqAuxMqxbMHT/MsqTbu95gGtYigBqna/8snSPTraHvzHIQA0GhNEMklgO
j6aZ8vXMLBYR4z4E/fEdBbyQ9psWsK38/4tI0AA3bee8nESLSf9WWujOYNFnnRBx
WcAO91Sc/fwI4v0j4S5Deez7UCXh2sY5g2hP1CqbLdJ3dp4VZNZjQ6sXeGFcGSrB
GGVs2nO7XQZuF1eNaFxBMzEuDRBduk3QLqhfq6LY4MM29qiw9kcUAnPLdSuY1D12
uIZCKe+p0NFB8DES9EfeExnYxN11Y2BYeEN4CJcjfE3Pq2cFqdYiat74adkdB2WH
nt1nAu+WdYQH6jY1L0e5GDQgr6yvQCtVnT2V3knLwmqjluqqSwPPnaypgRK+0XZx
vlYYA2SQiX0W488nfhAFG6XQUdeNdQ6dWSc47OAwRE1yOrcICwWvgGEf4nk0dFyl
VrAZ1fZ2nQOSLwxYGC78bsgzKx1IdYuqR8VQWDSeuYIAA/4Zf7JIU2lSVKh5tR8y
kaMX9M/ElzgNhFjSqqpiugJDDydpzz6s7vu1oK2oWXNeibeehgnhO8/5VywSnptm
ASEMoz2TUaEObQ5ZKCt0I6VGMuaMPx0kgjp6l1lV7Hc/APZKzpPV/j+Ij6buyaKK
cA/vgZsszaJqYSpd0r+0WrRutSJNN0i6iYqlBHq8H20XZs9GDdkn0tsGuegbHVmT
CAtSacpGsP8Jhek/g+awXfzKSPKWQFFnmWxg+Q/uVet/9i4kZZlXPNeZ3Fi6pWeF
cAj+fAMjPkde9J2a2Ne8jJjt6q9Z3BQrb6UKVgmgwT/a3JFMb2QGHkJAd6EppQcK
1sWpb55IdJTVtaqXvhbrFee8DWzHbFbOg5818zUQetQbPCHVhmAjS2TaGcuRgekL
OEtdeyWHRwn1xSsBSsJG/I4T2TvCxnD9//DHzJS/0bmiTwE1tJdluUJiKZaeLPhF
OFP5LU5GQJ2hsxMn6cLLIE29srvqR/dQBf+Txkx0yZ8e4LYNQxC6lHcMaxM+CBsK
yiD+3iOBl9Xr4TFmM3fyJC1jWvgkcoWnowxnmDOc6EK6I5N98rTzEngazrDWOvhY
lRHdgaBCkqRyVxeV+fAufp3e/fQjQKvKvfXNpwRaWG4XHD/zCVilXtpv8WSfgiHT
ILyJKxWxffmfpgyJ9AGwNCcFtOanrd3IyDeszEL5TwBpBelFUPycbl1KIbYK3OYp
o4EARqAkUXUicFnY5zIZ72rCbPGNQHoj9KwUqOAM3RY573GH/W9QCcGUr3zJGwCl
2PqIoZApbWCxRlPqrviVQpp4xVHnJYo2IFPoSgamtmRulXPSnyRCoSw/YtdKtdAN
BBBz01YK7m/RkGiD6zsjcATpLuvJAEbO4rUQEoeJXNRcgXVg8Xi2NMdMH6hzmhYW
hUCZGcGRGnwDrdqqTY0rOmHJGZk82lQGcWHPJPHtaKvEBLZAItJ1kL972vrPBhOl
kDlaq6O95cE2UGsbas9OrRjXDAav3FQOys+bpbuJhHNyeLA025Uo/8AxGK5H1deb
eOyi/munhWPyGJsFk1tz4seepwkYeEY1XAz1+L+n6mq+MP+Y4xo3yzjiZK93ccpy
YpRlLxVIfwUFytIDjkr53v2tQ7MQOrmS9Rnicp4WnQ/JY/b2lQZWiyLdMANYvYDR
4RXitKtmBZ7XXF9dvqA6DyZG/9WhHmEpXvWvjqoct19CyqvwqsQTL3drR4Ea5RQf
UVs+LgOEzW6+TF5pZetvODzHw8wUHe5UNZpXnrZxdIB3o1n5pn+ayiVQglKvgiZR
X9nplm6P+QjOa3nQexEPswQ4ANS239Rr1ajbn6CrPa7S4nOSQ2AQIp0RH+v7EN5t
+9Equs3QTpH0D5W/x8IpV4EXXy+ZJVWGwk2aZrWd6msQGYlMZnZHPKl9KL+T/xCM
y+4BawSydk8yt6JIFE3HhqnzNGH6n7DymLR2YhTOxtuFavM7FTmgNUckg15pcWb/
T6j9J14yP9+Bf0RZmJ8Pfq51GYOZ843R0PY811he6KR+f98u2QXmucGVLFB1E1n1
QA6bOGOVlUONrZFyb+RKwkrGPCpX203/Uki39H7U6G9PCRW1RQ3djxKYl0CDIaab
qdSY1tFe1SNr+zKuB2QO1VjMpv6ToE5TMK9TyDqwoXMiZrDy69x20+etrgnBMxee
V0LwgSzcjukbvxiBS2f/vJGxy0sNt4fCdYKRiHKTYt8aFOpJFpKO7B4T49EbWrQP
7CjJEDyAHXzcsskt626CvPZA3/qAiyauwFjITn5JJlNkwDhmzIEtfycitngyPBa3
NsT1tvBz8JXnCez4brZ1qArOhu+NfMhUnfbf+byfOqLBku7yaX7xlDOjRg4SXg9N
FbbifQiQDYmo83iZt9a+vkoqUGJwLt9ohB/AWGdhPYy1kYJEgMgBnNPsGV9zEAVJ
MtVPIcNfwUAnOkvHowVh4nXoyNeryDVfblMhP17yg5Fi3JxzMxTkSVjyy7RYOHSD
S5ql+5zdecXxxVsl1uMWdjwhJB5LznxswLxUllCLLngS1n1F6xmcX0v1Fynmh9N/
8GoxCRY9bdxvOOYVm6f5/rSj1yyu5D2kZWhTgvapr/Mz+pobMQqfEt/mzkwkuEGY
uhX57rAUxf0dToRa/iTm7OH77GxXxntbCNrhVjJvaDAf3mwm/MJ5nYaVYAkmgiqM
pJlybqCEVkhrcFCCyWOdylQ5LrTZsJQgl+jww2JNXkVAkCV9FLh5qdT4vCDFDqRb
YLfjavx7H6+vmAjq/34PXWfUDnsw/biBwsy0caLa3/ADUABZgx3BsHU2llY0ZTq9
viKZSq7nRBD82wA/CXwpRyct/cXQjPBVf6qZTOQcIg+udVq/YBYnIAqZ3s2jgQ1o
5+N2+KMkmF9JZXoem7qT/0Gq3P66xUi5wgXKY18RyVnFbWvGtjvpZ1ybNkYsofNv
uPLLne78BOE3FI0MrinjX77jMVA7TSr5e+OyjOwVMiU9xAnrLC87Z2kV2KLpFPn0
lgolX9lNxqBKwjZcWLh1sB+5gmlUEVyBBRyPpO6ZVxDsHfM7wRwFtSGc2ZEGDQwh
mRZxX0btrB6414CszaHuzhW0dX/z3cAF8uoIC469xe6QVRLKvN6+zbpMtD/Gm5Dd
Jhn8fxnE3GJVEtpxdGAR+4KSX0rBSuUzEzmEhdMDvHDB3uVhBwjQ8JNHIgZTFZ8/
NNj6JKqrNQwhOCSXFJ5pW2nDsNVRCVX6xuecMALmEcVXStPZMElRdVHxw0PsrBN5
zkPblNvAgfdid6Ly2IjeyIrcZbTheBYhBTYdBgFR0H70be1VcSkNmWZZFY/6F/eR
Ep4DvU0CYf3R7J2zhsOo+xIWwkQTsX0y4j2K+PvQ8vMY/TGAW6k6S/oH6gHFf8/u
rtlY9fPX5Ge/OXUSQHrViWpbkKNUlUkdGNaFW/PDMK5zqQ6tQC0aFTiE4n0kfSJc
gpm9dwamoypvs5x52/QsnJGPajifCROJKM2qLA+hfhiL7iewTINTWNYi2ckPJfRp
u2ac8vgGpNR9nlXkAYUk7QHHjzY1yx1FxgatNi1wDUmLQXYaPmLkFwbhOLob/uOW
fvmu8/EamSCLzDrxLd5tndFdYBY0Jx4SXOPvwZop8opja02cSJnC5tRqth6yw8kb
KilGvRLY35RRbKahk7HNKhURd9b74m279uU0OTAUFcKK9aXnOZTCQpKhCWP0KT/2
bd5F53grF+f8OR/Q1gPiAbWF+8uOhAw5dlwKYz9h2WTQ7eR5Mc3f9VjLcnqcsSvA
iwB2Wl/O483jLaNJnNgKvFZ9PgW5SDnTercl2cxgwuD35fGTAOk9EP1upAVTK0jk
blJgMxZYuEZCQIqB60E1/Oxv7fUqL6yFtqY/t4uBxeb2l125UF6oYuf1KrPhP6/+
r8pFpYAyKxbdU5tH0eT/23ReHj6Gn0PTBl3Mpw5S2jgfoc46Y5hux4RZtfpgU9sa
yFP56mzTlB4VqbH4+4Ah7WLnWQ8y7jiolINEUynGbAklPGptKxp2WGYJVJHqMuqX
03OAyovNU4N8AS7TEqZvlT752zvf+1MP+P+iRbY6TF+oiykQtlJORTHg8bKHuwAJ
KiA6n0qqtztaJew6pbcLnAXy+RahEJC6Xn4BLaN28x69vIRcyEwL5TE0iJEnCQZN
ghOp5YdwHFFiNNpgvv5AOPCXS8eaX9x0gEgEcmdmsq9Qf0nCTiq/+8H+WeuwdIzj
rGCN0bmuPWj5Oqze0OCe1X1Nj09rqgiFrdc86Ln7vM7gZfikwh8SZdrcxp0KdbtC
I4SlC1tfLyLjjL1M0ErtREtRgozgzp7WO2uy5YDyetlzCeaDARCqR9/IVYgWqOrl
i/XrfttINPVe5f8b8rLoZ6xQVkbBIEv/gx0segWvjbsKN1VXMnNmOjZXPZ+T1I40
NuzuFuk+qd6Joq4DZdtx9N40qYh1hrHQGuD3CaT0CbVn9armv9OlN32WmG3vS/SS
/3bWUiuGB/GGmSgFgKhm1yhx3PDSl0M0jmuizSMvW4sGBuuYsnLSfjLi+3wW5ZYR
ms62eQdukVR6YdNNLSNY1P04YKjd2rzTDNnQ/iwi0BJ2Ld/ua3e7WmHkJA4pII05
X39a7K4KtbXRdLYW6x/esylluOxoshB06WWCdL1TURLk1TnwT1nsCHjh4koh6b8c
nEkVHuca21jspG3TLmClaLWGStwHU5rH4AFSlyDF5jSryvYjQ1Ko5UUEMUXho6K6
5fVF/wxitGZW1rFbJTu4wVNc16TWF4TSW0IQVtJm1/0vPdwsLud5YRkPuBKpVsot
adYe43AyyZ6ygMhW1vDMqdxbE2ioDOHbqeYO9T4/CYtaRJhdCn6lPASLQsISSdp5
SN759DlPAObyhTHzU1ar4aohtQ9BtKR8GOx4yB0FMIQdvjoiqdwgVAiBuRXRRZfB
/LXh22CyCk+JbSYpwrBKd/kXbFH7jB9ufX5uuZCZIrqcWsB5g0781q7T9GI9fXNw
Td5n72YvBagCK92VD8rME4ECgqzt35P0JcU7O3bA/2TwK7I9nGuy7KmQJgx0rpMW
yrqk3kod/ytY1JgAEDaimLtnoztjH215G+B5JB5LlQq70HT46ywwP8dRuBH9l6od
nTi0uuKM0rAvOZEglbjUBntqXfg802uyr0iH8yJ80Q3+dqaDZkCQZrMzhMxNJpEk
dQw35bpS1Kg7URFgi5rqNyjilzgaO8jdHHLw2AKnY+9R6xLILqN3OYu7/Iaqed5c
o+JsDgfojRp7EVwa8oT65qYkrg2NN9AHl66Xsa0viB3aRhhar68wMxupkPZeuBME
5pea9rm1xgMez5xSuqWHEfdVrfJqJs0etwi1GbqnQmUkvxrchNq9CK35/jUkoppO
32pu6DI5TdAvpQUXXIu+e3u6UCbAiP/EqH7nEiSnDHyBlFglHZrMVXBwruI4Yc0d
1/TKncNRSU0cpxVKvDmQtvAjUA8AsDWgLNpCYbDnNp39zCoImFKepJh4b6cSYPp5
erYzl8NgJSSnDnqAFidYbG+6CtOp/qyGJBReP02HMFrnmXf5mrlRrWumLXaPLoS7
8dOd8m6vTxequvQ1Tu1ISxMS/gpqOQJfiwNBZOj0SqMbmFBk9eQm/bbDgAvqXSVi
eLO2rfo4dOkfOUUUkMf5PTRMHWlzYj/torQ+F0krCcN0fwjcKL4hAeHvilc+ukyD
Xq/2Z0GE7diIVsqsKC1jIR/kq2smsgW5uf2tKgKUNw8PbImSPkefMLb6KnZDwMRa
CXi4yjnzCOGPV26aQeJXZHUh//yjpf6ibBf1ApUvmIuwhqdV1ehIHKZwekSkPlNm
ul+kAMOfswL6tzAPsuetdLS4FcssDKADYwGxtru/rgEDR1wETBxSS7q+aen4EEhF
SNwJJOTSr+toaY0MVySgRKOJCj+I0daDOFe04qSJgMQrAFA3swEqMTFRxlYMAZdZ
szslLMN+D9h9Uj0ZcnYlRqEXkt2fHLPK7hAmzDUTvGZ8n/UJXUSI7971qQz9w+CQ
gPg73Vk1ra6q/La9E62bBEsZq6ryjAHp7eJv1tVmh9c58xsF8WCCBKOKUMyg0Iwp
xLSQpeHwT2znRyKUE9AbSw7nl1LiB9fK/qD5gLMxQLJxuE5Vyt6xAw15Onp3x+Va
nXcP4ULFRv+elBidwihV76jtqkzqcGuwtbbyKbfedJEiisjSW6+w0sCf9qqMcdTZ
ozkx1gogoR7hLAYwD6dmvNh6QFsfwlP/JD4uiBzCLHXhAkecR1uTRUiE1Cz3gyay
NL+UB5vhAaEuWBB7qx1tLyxWPgyMPrIKP2/lfORHDWp5iko0Odj/pr3Wr9fWEtHZ
EKUMrR68YtUrLUPZc7lNsMz0/hpxFGr71cNRNU9APM6RaZud5+WYoKjXOXnMG/Ry
FjhItkn1l9ED9T9I+6MxszfFKD+UP3Ux5jt/ptvZY3lelxcVHPlVZcrTe4yNoPnJ
uAVyUnER78W0OitN4N5Jzuwl3t2hL9qzYwBxG46ITvrwipzH/9juS0hYyoIqiyqX
2JKcjG+XkB772Q0eoZqHRsNoy+uJKdcsXR2fTbxSOO7qwxqrM2XsKvBkGe0L/mub
Qbqfuk5Banz04XZSv6Ehu9EqdF47Qkr0KtwsY3GyB2gvWufR5jUa86ecG2hX4GwS
W/XJRymc+5XLGL9L3i0MhjMxW4stkKX/9YIb1ZK7GJ6s+yJ++929Z6QdnX1p15Nb
YfaB/ULGh4V27eJHcrwOgv7ECRJXzq1AqtyCatT2lS2VP29JsK/iwmjYpzKPBV5N
kQmoKQqFhTfRoaw/xPuiYHzI21CgtNdgQQkRHV6sBQAgAeBotZc2Tv7Wk4byg5q7
KwS1Nf+Rxnmb0T6pSRL8MJs19iaWOC/wd1pUaq8PvBtit78Yr6CE33S6BSdM2NBb
zZ6rOQaAwGWWPHXn89pKcXoO68uGqFm2GWuSs6YF3GmIxQncup0lNEXK1JY/z/4W
ceMS9QxonLxeYoXa9AGGlQ32dmFIWdyrV/9ASDiHILOTC1vPLVJRDhNKEuZc0KVz
JX+1TydFUsAW1PuYVtpEog3hMVCfcMNGrXp0MMiZ4UI7tNQT8V/21V2638tUgTCG
1dSkhN62uygFhcT7GIYB6w8JIg6/FgqR86SODQKVwR8JmHPXGQAIHnhKRu7ScWzY
EQGa6yHCMBXvx09X0keKuT0geHEogyfMzJIyWHLjooxWzH0fY5TIqA2UArlsgzWm
KWvwoqzAyQpPHmr6fcWMqD0PH18Q0TOE/86h21v7qlWyb5+46kqMIzL/L5HfQMOj
XRTV5C8X6zUq+wce7MCmoFWzY58WOHxX7phFhyUGrbLtHeoVO3z6tx9xHqHQvUY4
K3+68EP+GTm/PFHx2k3Gb/4HznfOWLJ8EKK9jZ/LwnUuKeG9cjIQdXpUtOItsMqj
iZh3ehEaJ3hA8hIhxxS+YCZ0AzaqMDzIpgJrIbzUEvqq7s7NBM9F+G+y/nGPq+HG
gcsKkZA8ppGzcvZKD62hfOceC+iXtBVnSzokpfvhl2MR2tbs6FPIrOPiRsv5AYOO
O9A9cyGRP6ljl7Xrru1lHoKxZnCe9+bv3Xl4Xoc80U8lyEatRDhznzMvHkpKa3Op
wExRBZIBdtxEfsW290+dWWYfvfHiyhbYPjRJR6D6yNAJtnQ0gxq1U01IkSonyTcS
YuJfW6e6WOWcKEeEBaznPq5ag12avGiCN+HsVsr81RpprLKqAxkVrzOpYRupdF9o
dUYHcdhGggRix5KgcKN8jf1o5yb+DquqZpGzYLkNbfw+y058MsmQc4JMgTCXxNT0
MBzkoEXikfF/5ku2fRQplR3MLrY4eff/ubQSm6bdvjmX1MrJwcR5oKXxEmouSQOk
jKVXY/iKhVk8WcQzHq7sNCBZ2rvbnv7OnjYDqv3HaEmrCFL2J6kdN2soe0fLAOJx
hZLkM6mqKf7h2bY56tBAQrBfIINPcTyIBLoKfUa193lgMEWO7EqqG1eo8bIMCCAn
8sullIzmHwHEtiBdoxyEj3q8vpQ8DgN0bbhfpAq6DB60W5owu9m8AyOSWAlIUQ6P
G6zPdITSUWoxLRPh55/seb3cyBXOiOBoAHJwiEN3xRXjuDF1txYpM/zBreKTi5jO
LCkztz7tpObQPawd5sKjOpomQ9wHIMaiodAAkjIFB3Vk2L66xPvhqLghIzZ6CqL4
KHvbySyTx7Ega2oEiAID4yeMk/IRwfngAJIHpYt/AwruvnBetUpj8kZRPBJQwZkU
4l2+pvFuZDXe8Bq1voyK4IcWoLTRNPlsoGsGbMGcWJwsPTlrV6qDCC/w8RYeDvGT
WzJHrm30TiGAlPaAH5rVYQZtNJOW/pJzLIdbu7MnPsO/vIYlLqVytZvLQO6+aWF9
8+P6X4Uv+GVcYNisZFRdrtbXmULgmYC0sWWSsHcsLcIZ5BhZBzL2j/bt9biyrXF4
gbsldqVDbs3mZs/7zI8sLSh4GLGxNtMLq4sx9xf93ZN/KQ748WUI9g9zAptGhjft
ITESMo1Q6IQusl+nqziUH4YyRx73XMVM2BbKjF8Jn5oBRiRsSqjEtpHXQM0IZSiU
490P3O2EIJbCC8Z28NUh0ADT8U5DMN+PvLooVyYdVjbNjmhe07f2JqCaFIRit1yU
cAdlNzZE5+kK0JJIoQyBtkYL6IPwI06Cc+6s7OQs4QylG86FxyCEbMtjY7snWDQy
XWGS6uoTjKfxRLXN8nQfxRTce7AfUvXT2muxvlFlkycz9Jo8KdJpxB7SiuJEHL2h
i9Tx5HD1UgNngGTR4ljxWKH9pT0AG4UJPkV1o2YEQRraDL9dINfJuf9k4DHnZeGn
yNYBSmiqL90r3SwNpxUbjSbmvNbNHvQkboW18DsEecBE60Q+Fi37q5UBJWO3Ap1h
2WWi8+zp9QiXLHe26U83hOI1lTfoGW9t/A9RJfmIiVliJFK2dniB4Wn5sYI3QbLU
3nw/7V2HFIlVe+D8Qf7Y8qopcmiOIUZzO3MpXoHGRS28bUE1o6G89DSrRuN3OjrU
+WPG+hHXDYV16MUA0w0utJWuuearJ10Otwa+3wpbxfETpcWnwG9KG86AL6Y4+W+s
IAxCQXTPxqlKVI/62yhG1eVSDjZY9Xd0+iyAAvJiJe8xmw0jRvx+RxXrthk5zXyL
oyDLaeWKs259O2IOZjnyXX+6mAkE0QoKmsMml+tarHfk4FTFjEIPyjGgVdrXMazn
J7NnIoZHkZ90EAVnzSMFidTzQ5Vfloq/GwD0SJyT31iTP906IXt1b1WplWyfuAXB
dtAahzFJUbjq1ClZPID7B6K4km+MwMTUnwLkZBSfmGHwxWio2jlovM9z+AxMSB/F
E6HCv9+oWDUSqToULKJqfQEJeSTztWWxVNNb1qdSQI+8X2/t4WXQGH7yXbNpuVEb
k66D1fc+KfEASl9Epa90ocI+EeP101G2VB+tvzqMqDTIAkIcZXdtxSSS7tB1BMUx
7qcD+U+QdycEHDPhwbVbVltEslDqjkcHWeOE+5oJ64s2tbtZIie5byYRbDwLkrMW
iFewY3rZA49qqOJfDxUIHRNx4ctYc0FE5QC7Qn4rfy3V/OLQLQL0FhvcvhaU+F2Y
6k0tLdcdEuxbLx9t8jMliDOSH98+0oNVeSHPlMCMWFijFiwNBA9Wq4O/HCZtW0wv
txt27BteQkLQ+V6tZ5oGsuvCED3IqFZdSj+aZIqtnJf67Zz7yHwXSC+19RYIMiMC
O9uyhaW8U2p2mI0EgyYSWbNQ9tH4sVgx2Ua/lk07UIYYUS5wGQZC81tsyFTPikTc
3nrsl92IW0gBlaNcq4IYgJCCxOqGsPJr5/qfkApeSdqltV1RR2TmQCiP7/oTYykU
v/j4yrBIu2ZrgxPlRELxBZ04yCugrv06Swu6DuK4/B4vnR9JCWLrRa8+L9UWT57n
eJIzuFzBY26IIxPlEToldI7gzoe+w/rbntxU5W4ZnN6AtAT5FoahzqBYnmHBblvO
D5vt2sInSCyEK6fslDwfFuD9jJZmQeMmarc8jYIT6BLQD3SqzKhTdjbwWteY/HF1
1MOjqBL3GmPazpTkSVhePEvr8UoCW+At68aJDwKb8VR9xj1tGDuZ+MgzsFe8DS5I
YKY9u/5C78VWNRwsFyql1hiiuPonKIFPocFzVvlS63RJMoxs1Q0FRjtXIRARBeuD
HfTURVahmHkgCx/xts2LZ2T4oNUUv45s478CWbRaiWXBWM5kZ792U+2py6Z7fOhi
N2YiobYN2F1pk9tkdk6c3dEeKct/G4hMZ+ytRnPsMzFuOMaTXV1qAmtYg3eX7Naq
IUvvYbzZ0TlIN1p4psMt42wzFXCqu7GpwRCMznfORZX63y7WhIqYR93yXcLsZpzb
YeUBBwj7v+UmYVRepiIFKbDP46mBNzskkCWR/lYo8qWJh7Zd+uZB13URXeUZY0uE
DVCHcpOd7C6b/mn272f0qxLmwIykU/7/PRqWyi3DVM3Q9psHtHRULOcYIKe7QeLR
GX9OW1GNc2aZyWjwkowAlj5YNfB2AcDIDYxhkjlr6hjDVfwtdaGW3UBNmM+4lawU
LcdFdrHi3XTgdf39cB5EuoJDIM+HyCH5mFds72fcNdZqL2papQ+/8h/wXX4IQViM
5n4zYZ+BR4+ioTt88YAHWKz2lvesmlcJwwZyreDgLnoYoSSfJ3p/+stp88Ae7Kec
o04Ii2qr9wLRabz8M1/LWqAIJdSBdtkmi9cENO/lGdscF1R5qeMNvLqgYnoE1KxB
ujsKNuiizP3OrpWMG2c5Ry1DpSi7u3Z+npfjQsQ3yTFC50oEfUVXYWNXddn/KY6x
+AKDg9B5bVveGIWxXL1GRzQHeSKm0mNFFy1RHra5RcfNIgA9BJUKy0cgCuQEapIi
n46OS8dIw4/VquRa5u7pXDWOhJXM+BKesC3RmGvZGU6mdf8FTdfaM5NyY9KXJ6jL
2JnN50adyAxoo/vvF3WygDa+uMVjGJ+nLxC7wQh/TLR4X0NXRoA8QGhALpdE2z8H
uXnjHH/vHYcQ3w7/cMOf2i6SiOTnYUXB3l5gGu/bDZ3ne78UoJLZy390lVO/HbKZ
AaZ/8rttOPlSr/6VVgMEd4GvCZGVVX3u5QdoqrBXWC7r6aBnUfIQ9yI5ziH2nNhl
2pjZ9JTq10UeUsdgB/jmuxBljz9MrO1BOe8lhPwRpfdNpW1wRhcp3njO1XFURhiP
yOjoQuBGPmB8BgT+WSvsMsnvS1Gs9rzn23dL+ifsJrYAe2fKBtxpbNbxfPHIssjl
BUaoOKPOGuZxgZh1LAeUxVinHgyV1RQ3cCy8iiW0RNoOiomyj/9WT2kq4LD3KdMc
pdWaua6bmbdQRA7m/+lkF1rjPNlBAQhFTwDdPiRjuk3/nhBDYTXMC+YOhMSSo26v
HKsV0RQVAXP6inuPpL1PdZ76md42SBxh0fQKRaS0jwtE8uKkV6wyeNKpIq8Wk0EW
wM+82IlnGPZlnRg4p0CS7/TADT75zt80N4GMYqggpz2lAUUIqJWY94QOQE8Ux15t
dgXttdRb/npY5Cj0ygKtce8gTaDu0bh4JgrUzIyUK+DfSr/QH9tbf2Sw5Maoy+/E
N8OjlR5PQQUIvrDFnA2nJYH6/VfUCSz/hdx/Xa5s5LTtIqwG0R30Zqfhqa2roZ3D
r99wYfj+MGw784V1n72EcTVb3QiYV/0PIP42UaoDOyuurjpkJcSI47DGJAKlsPXw
2zFoyUb0pgMJFDCrdxCGJFbF2YkHs/Z9+En6mkvvu9VB7nlbXNdrQtGwgj29qQqz
wLZGPMSxeb1TrouZZb9CaAdrvWHRp02hABXmdHsyJSieHTPuB6DcqxyUcx0dIuKu
9sy5K0Bgkt7RvZPx88d7JXKRrSpIMHgV1RNhTgUN+F0bVKkiFIIRoVA2iZf2E5u1
Fc43XMgU33JK1z9sUOIK3klD6WFRFq28mGFfkkPrAHZcPGmBrt7o3Rr1Bt/8ub5X
zlC2kjOxcWCQeTfrb1mwXnKX9Sv4NzE0/49LEWUrHMqobT4mltFHw6/GX0EMWDAq
UI+CeHHBE2IfGvm/EkDy0QHgpZPJqqQHuQBckYCZQGRTXSvYYX0SvXsuX4kO5AWh
fZmzNf3XkSySbCIR/s66OwtKi5YbOWGNk//bHJ7Rfgp7pdVyjFwapp2qpW3X+GtA
4oJkgHcXQqQ+fsad4Su4sMDRTfqlpfaE6GUxQ+5iA9sVvnaerCRIWpydA1GDa5NJ
XgDOFwrCNOVknLPk0smOWx1o6qaDB1zerZ2jiNjSZNsMf4JPhAGh9xq8ssJCae/9
fHZVbnP7AbPioeDeeUEyiiSVKYyExmnq3WGXKLWgw8VXT6w74m+/FIQtqKHmFSjY
ImXcNhIsA8QUiKocFF3insIoxc7HI2cus9mks4si8//upiGIz6zHEF2mhOdVXXm9
QBYVV47v/PCYhukDRDQjLc3viOW4ZYRwXQYa8gW4OKQLyIH22ko7eLExFR6bhPxp
6vj7Aj+Q3WY5WpsYcUgoU2gIBE8s+sQ/wYoiLVhEp7Xr+fJ5NOh6fUkCES8sWXMA
+TCF73qGc4GGPdUxDhAztB499rprw91s+Gy9cyySyF4qxGz+YRxAMMupcllOBo/5
SYHGttFmH79PZsGxGkdpAovEhRDkRKrfleD5EfPtTc8BRMAcA7YgCKAukTbZOnZe
+2YX/MVvyKMwOrRd8CrswSJgglZPEZuBbsK+uwdSTvmyjmHY7xtdLxZ3PkaFqP+K
B7X3q8yyJUV0SU6MyEJicBZpsGjJf5yb4KQysxxILUrMpHPgRBp7q6y4rdxkKOYo
dMnYGvKjaxMAqImkQI3drboPqoKNOS2c3pxzs2Cw3SMu8n2q5DtJfn9TUbAxBCtL
9xTyTbhwBwaZiWowjfMTbGWzki7rtq+i4f3APqlEYSUIbIgXCzucMjlFJbh9+wMe
DimqwSa5hgrG4fATR+8DZFWl8rPFOGbnD7eIHehHe1KICEcq5pbR/g81d4BOx8iv
rkkgCBe69Yzr9eucjRxyMCwypI4vAKCdL0cOIuT3AVl7QPpO3bL8Ry+tdIuiApMv
EUTpCYmjydLBJoyY9klkfXu09vNmToLs9xl1OMUJaCsFN4YSRMP1kwf1QaRTtVss
/lWvPkBxGYc7A08ChZ/54SeLRMXm5shiGoPhKFCPrGi1rggcVlEnZziTITiIzPu1
/xUPlD0dCtP8MVKF2IosiN03uo2cjunPkm4mS2CFHR02bM2Svv1llrhonJapdV1W
GhVxJNt4IOx+mnTNOAsx2EgPQg6higFiHpBgneoegpRRWnu/hQO9FJDgWyxRsLdq
hk8hNM1PXrZRAJo3/v0UAOngSC6fCSNRCxST57GQGF7nY94qMinLtflC2YK2Z4K0
YIoNBMp7Y0yN4+lIsnKcYIm/I7xTykpPSxLJRVpXvyelJJrNN+XJqzv/kxGHfWPv
GE4rJAe56cAhOU756lz5e2KBJQ+vII5n62GqkGa4aRW8m1ffVpfi8X2K0Rgp0Iz6
+eN10zO4cYctqp+jJfgLCTk0nr7vAbnjW+oc4K1gLD3X7S6RLPrmQGz9Ysjb/gGp
kVygVz/Cq3Ek+ygPGVH+AlUGsZt2SKKlw6e0B8OqGnfdPlLOwZazbLxLUjem9ZqO
T88gQPF+fUcHfG8fhiin2NPDQ+En4SiV6RdwXNnEcX+JYpJqbrhacYxhT9I8Es12
pL1FzAsB5tDT119dK7yAIqMVFVLj/5DVFf58YJBTIHHPywg9sYDTn6VrIFGJSiP4
PLWluyA0hTsiUDs2w5tF304Seddp/4lSdIHVXC3qaW7aydNYzHWoLPzXE40AolLn
rdwAnuykhvyhsIW+9cGstIgjV4KJmS9NdBGI5DLBQWcxkCL1uw/yvQzApXmCO8VB
hKOJ6866hdvVkVfwVgyI58wb4vj4+uSehOi6j8i6wpwufVYncSCIkLUHsX2Kqozb
oG+SuzQ2a5gBIC8r/bidyQzvCGBdOWbQ4e6bbiQ8SVqiuHILiHzXjnD8KMszuzQ2
ayhPFkF9V30m31gnjOWRJ1PcqM1KwlV7+Dzm/k13qPrMdfFEslx7ZCJCOmvDxGuX
1NZDyg4TkYdgxrIm/5kkuVVqcRFS+e4ngdWBQ2Y8MGaCl541AesQXLrTv3qVGGXi
jpMAYqP+N/9CXrCGJtMVIVRy0+ZwaqgMQQEmq+u+cpYpSiVWkwtTvSk7Z1cjumHv
Z9XcV839P8VApjmY+0Iboleqp+c+Satykuvxq5WJWDokJY9ifOsU/166WnLq3Xlm
hxj0Lfr665L/ePz8SpnMZr8iiOUILAKtIDLFYekvD7N9hO6enRfJkBZFrBugzVj6
xUB9O2yJmHqSmoBdc8xQJBQCYPiy/VnDOKn27Sg2LamtATJDPXcvAnimWbyY1gjV
wkwqY9gNQ0Lz7GLcVWvRdW2GFUTz8sxSTOF1g+loMAFOeBdbfAL1/wqSbBE8NDMk
beM2I/o2OaYLHZ3YT+oOjECO43UQvYNuJXkdoF/I2G7o1/ff8EzbWsazKQKj6gOl
4TgJBvdtco5Hj24V8Ai9z5wKknYZ07U2r5LpebjUVzzkOHGiI5yJqzfZqf9LQLY7
KpyIYPObGhl6YhXe9BnJNFzDY4POmAZ3JB2yufnii6Okr/xJJFQEAG7NPm8GniYV
2ZTZeHQ5BeuF8rKiY/kmfeM266BuSUPIINOwpzsWMq1a447S8M6tUNqp4fyCYYgr
jxgruiMCmq6+TyKh0kDNzfBceCZyFe80gr3ujzB4hoLer+LfYpXDQAYm/cmXrSGR
brSUhw1Kh0GgqZmjh66fj6WlZaaQ3mbPA9C5v59AGRKoFZjoIjzOQ4VMSwtF9IbM
nvBRucgsAQX7BAAXh6A6PLjeT216BsMwsXLzJ9ivDvYYfvwswY3kh8W9JmpJM57Y
g9L57xKwjLWN+jUK5bdUQ0IsGn87pHtXq1eQ4U8SOXJwVRQNCyJ+4nDuAaT2GKP3
ysjZ06sONu3KYuLHi1Idu+UTvjV7F6fPmZe+xillSHq5XLINH65yWQB3TsCJGjQq
blevlFNjgQ0XU1SXjvYqQUtbu1Gvfn4T6KuwTs5yIfe2MXlEx+Rudt0SjbjBmrsK
TP9szaUDsft+uICpepcPW5RSDTr3Z4Cggvg5Sjsq7t486divLe7HEok03WC3mFOi
h71gOT8ZJNqNpQwrKP/NbNhrwZKv78D2x1Vw3uOdka2un1y7br9t1qElqm8Y4Pl4
odSx/emD4qd8m1q5vdtODVoMuidm/Vf0KaRB5y8Qj5gEKf6QSGzcfmr/qzcVvM+Q
KVGD7C7iI9lAwG26mbTGvtfZp0r2tYYoNG4XVGX9myahetfGFhkCpjD4oAm6doeq
nDuJInNRm4hp4wT6+vVZzV2oZifrxQxqO9ohvl3e+i8bogfwVU+X8egWHgbV0zG2
Sp1KcaslMrIdEqTPcSDp3mSz/vrQJP45qDaG5QX61gU+ihW0/ZpMuZ//tA8BqpiN
Kqwg3V/knLEXJU3hqBauVdXBuN7zUk3TV/63qObOkHREylsByUdZhlUHW0PIr8jK
gpYpJ52MLToyybnpl29w1eqbsOcBPh+PYfIy+NvBwv3eza7BnSbJdUJJg+333MAC
4fmd4AAfCnkkgNSLPMq4BMPe58Pev5OJH5EjksgZMHhlA/ZUL7oNBgkmKYkeQvGi
EBvHyA+KrE1AlfxRdb3q7i4O1+2KlKa5lePgPzWhmKLaB7IYd+PHu3Vc2towmFUC
WNlhDphUgOgaaHVKx0cqPknf2y3rv2sIYz7FmZiFvtJqJH81aUz3gnvoLQ7vY/oQ
ZjyOQFsfvAEYT2kaQ/cXhIWnTEbc9vxcT8iRhSi7+4q2Lv1HHTs2UREZu8F1lk39
tBXYQ/AcWX0zn0FRL6BXCVgFxQiFzWzEYiMdQ2lFQYiO2ijUw3Bl+Z9a2/ZjdKWa
BwwazdnzBKFnrnF1C3iECVTrPxh2Keb7R60yf5kuw3X2xW4wSzK0+HzqWrmZKFyG
USEj502HPp2bIvEeiy38aIY0H07cBsJVK+98SyeDG9fsuwBljEhETINCWShBZjqq
/vVuo1kgxDV3rv6hQQRWjvqNedqJYouWgS3HiVNRhjMdYEserQkJiwJNk46Y5o5x
v2I1rlOz/1oaSq14ZSl534L8DKPxQj5Lkm+wIJ8pvXr/3WPdkvszCC4RUS2ebWgU
JxYbOx7KHZ6NvA3xMSVTUuJ/Mw2knt+nT9Rp/zcAlY0P5sdHJ+b1yBtlm0mSp/bZ
kmH9t3ZLXrM0S+7vl9Z5RKvW/MUyu/TwQkLNL4vmEBlIK4Mf5qcKfNlgndiHnO39
TFyPLyTom8q6FpXUhgzFDySib+ux8+vHwPLpKm2r46j/vSTbeUGifBaWqKZg8+Y/
mHGYkN5RmCnpXUzjarl7dj/qwLyENp8AOuE6MG5CaC9e55HZ+A6tiDeBLTswndrN
zAN5uP6lvZqJJ3zsFg2huQ4fWvOfc76d/fHKibpxnDz5VOGnIfkZJEBJC/dxbkX0
lEmNwuE3I+S/bR24K9gheuDwE3xhtvPB/8Av9w3yRwsBnXEVIxxbK+/cu+Yekice
NTBbyzBMgvIvGYTn2H76LGRhXIxDG7xeaFtbo7A02iUoH/t+cUNfH+6bLbh6Ozsg
b6yhejcCpT2BM4g7/QVVLI0/K3LUv2xhb1v3vjMrWDAjva/vHPqWnPEwK1ZzCdxs
gcSB7JYVEI3mxsnJiOIOpgAoaMtaR7IUVqZRToycLNVKqoTrisK/sWWZnliMbsuj
6o/kdQb6iBt0ZZahRYKK6KZDLAk6cLGRRlf1otdK/ULFK7uqsflgQaTojrS4sKdv
5ns6ZWnTNm8mZhBzUgwK8nnmdTL0o9n1rJxG0/WtUYFJt53g8X7kKmfjrdsR9Kmv
ViwDlscPa/BslT9TMTR9tKyCGWjhCO4c6auA/R0R9BccPQkD4KoxvEjHeUrKF/z9
1hzD5f0rRj8iXug79p+QoLpjn4XE6/RYVHuNDBWn9sHOOZfo7ScsZWrR4Rx8OgYX
x9QkjajQzJzrfN0yUzY6ENUDTedQXdtqko6jEn4dJSuA4q7Rd/9UfE33xM+e94eL
W+ixcQyLcHqXLi/SrOb2EfvOOU2TmkBpokETcPVaiF8YMcq0lEZMtjRDTbo2cC9f
NqE06R+QCmH21uhUqxNgZOe2Fb/PBQ0pr6is+Z+I5t5+yoMPZsdFrmW9msoKe2dH
AlCwMyAfaY3TC4wJLoJlKJmoAEwR1SozEgnCetaPN+9O9u1oRhR2t7TDyl/YHRiP
QI+tXNa5jG5Yu5J6bJsgDUqX4++CkV7oky8zHvW2MrBn3/gzHqTGCza9B3rViGZA
/E22ECgvsGTDcCK6BVaHXqM1x5pxYc+henIfNh1XH0qrG2EZJxOxK7XE46uGkUMz
//otea+qpDyDbUCMN21AjkYEKDhWTBb1ZKFlVHHTQ2zuBZdMSRe1OtihE4VbCF8k
sueFSyPbJAc7yswBenpyWzn81yWbTO4n9XWwx3KD7jGo63l5D70BfrQbGGA0L5Jk
+ZR0C112lwkbIKu3U0RIC4jh55zSyroQ9j9gvIUjUFJS5pachwxDNOA6BIHZnLGq
3JVDlR/r/BRJpnJV7J4ftta9XdIXFQv6OrQrBAWFQneiPiNZufjz2uejonw3mrle
4yKvYWl88nzUBZa+Dk6h2yqfIiHG6Dq2ZDmg19SyP/a9wRrkGydHugSSq7JZMhlm
Ynu/nclqP73PogUWMYXk5/6P4px2RsntGrm4h3E2WfVKAlh4XzAskzIBiRvOC5l2
6MEreTOLCWF77HkiUTu7xkV7DJwyhEsUeqWrvzzWtab6hPmeSv0AJYB7Ot8/wvcq
NOb9EIQ58dWBCMXbGRGFT+eF/ERFtPu8TwT/MNhyBP8nPaWembO2NJ4V+fjvHiN/
jUDOZfUhhRxeVTI0WpwNIuMFuw2cIQegnww1k7M0oBd26cV0pRvO8Q1xsS0wevJz
/KelRj1KGyIbOkn24VxDFs/CjMXE3jlJPjz4s4AX/kYVXgF+biwmuS8QyDOkIeGL
iQjnNgb35HpowPnwjA4BNYEL9GGYq+ZHk4s5szSni/H/j45d7qT3NT2hdeeWou9X
thgzg3bxQBc66yStgkSouZrOd7H8HUhPSFtDH/tVnXEaw9iJtxkhUz9n9MNnqcBU
CNjPS3nGngE7IqffYmfw2n4vJWV9lLXFJ0qMk1/gO2dLrXtDEo3BHZtKuscLHMNv
IvN3Rj8slr4LpUm1qUPWegGGhm9XCL7VivKoBDrfZEB/+dFCwi6BjG2o8aRzKjv1
zH4tUskVRq2gcPqK9kQsY3W46qO3p+Tl281cxNYPojaAStMGc0ULd9gGgzeQXl20
SYnNCfSpcuwv/bzXqK3+2XHnc5aT5kkQapyw082WI1Kw8gHAqBn4zpGyNN7+CMpp
XUjSzaxBJqmH50xt8GC67SbkBOrAKGGBCu0MDstEgjobZxX0K84YdaJecu3q2Z+t
VycdjTJqR6V9zy7IY+bENNmXcOfBgLULlB6XccWxPppldKxJWVejBLC0eHC6xSM4
kwP3nnRdbqot11mUDYU7UJrwQMYwelZjfxbvLG2MWjBBGSZRYGGFkVkRNL8SMIjt
I4uw/FqZQZ6kl+cxgLUh4QwWn31zckTh/KZ9FoE3tgz6jAuApT905SX4J3pZk3zH
5mREkTQNAASlpl8Kb/bzSK9+dvgqpX2J1dyhMYWICg+iSN8te9MP3PH8L/eDmjuj
0o1AMN2x1Ui5cNM4DHVqAyp1euzSejy7/e/CqeyWzLkwKGZJV/j0Ve1BbfYisdWC
mB26C/qvAZps9rV1Oy9idvHLTCgzzqcE3EyaodN8nyNHvfz96yGLxH21cnMgz4wD
hW3VPCo+N2e/a1FQRnZOy1QPHgooSyxPQIHpX2c9Var987dELoVdDeHEjBFWd+Dx
S39NM1XSrwEoFFvk8EqxNyFL6nqxoBPV/LjEXTH3PYLZyw+bz9Y2QHZdOyktkSMT
5X/18myquW3liju9SfPksKek6Ib4b84jgC+0XO4V+3IFrFM2H9jql+st8ajTglCa
isSuy58EkS6AUB3mUJx0kbid2uRMQWsZ7JIPLGziVqzcziniLtG3gpLpsge41so/
b1AwnCPucOiqzdCG0SohhM7FtPSEx+IAYy9NbirEqRpWU+XeASGKdAWKhVcpZw8V
B3L1X1tCqTA9CYhyIqhLKofHDdSIaxT4VY+02TOdFAgVKpBnoSRkVF7+0t07S1yg
g4hzDTSq6u9wI3Md52TDddMqZRUcCv8LcBkhqWiaiTCoJC7ySuhBBUPWYqsRjzno
YPW5qCqQ9k8PrU9KZZdAWChS6HtVUPZSlGJ7yC6w1b1pDeruym5jwAQfWmsEpv8V
zcrHDgnNildKMMGvK/I2DeTzc+D3c6HYqzDvF44A9z1pFTqJjgqcHGZHQLNsXJ+V
8BegVtEOPVxAL2U7tzpRWsfhF76bBqnIG6sUY/mbAUgauf38Zw2a4zRZ4iAhD+dG
jptaTDVsHkOGlkE5oPtbl+dOdsWcCSuJLq/jxcQIC3hRAMX3lpW/Cl/lM1oyflbL
tkEwdO+GWV/K4mlFcXpcb4Kit6BDZMqjrKIR7l4sSUSN9t7q0pUcavK6oBTiHDP3
szJYTEeRvyfReKEcSaoKdwL5vrOGv4/JzZV+/6sx/zEoGD68++WHahqzTwqkQp36
ZbQ+z/FSkj+Tlg+9sABSmhpLU0b8yOoP9J0jxDblx06+hNFmWYNNh6VTgOKTm4RN
Jp3ck2N00YC42xpIh5bIqlQvg4y5bMb711m+8uf07CAcAhHVxKNKeCmgcxEUtz0C
jsxhNkG3p6JfHcB6QXTekmmtTbY1J/sWwefHKlDV+Qzz8gVz5wEqszKcn5ilegy7
Mm4FSdm5DC+y4DPao28drSYA0vOqbsU40or8vyYUOsrMQ2oJJRlOEYgC3Xpa9nf6
tQCeRL2jTKs6WY9NbnkBxAfJQ/SWAR+Jm5MmdfaqTi9oMtwAOC2SHeA7+635Um1E
Hi6hqnwZCY3o/GxBD3DI+wNuuRL6cQ2z4HuGZyCeLKaazjf3zM2ckhBE8BeZNb2c
IxyeB33hoZXDRaVlzXRWjpqAl3PFgiBTfdXNIbQjreppSWhy9OisSSbgZo3auWe9
FJfkj3/FyHZcb2LrIJpU8/v1BWbrAt4yeRU9rk9sgBhkRx2pwIo9ub9CKSAq2t0l
FpiteVM1o7fVaaOx/79HXQEle6CJGk5MO2I1Wf7XgF5c1CMXdib7AZZjRmvkE/Rt
Gy6T4y2hPUwxyMx0IIwKbLscPM5xSU2EUKoXHaGD+Q/6dMwi323nj5oTOm5mOq4X
VDN/EJuyC5Wek/F2oWesK2RnN9m65ju9sWPBRLHHolhJ7+aijCo2zpLWQCgwXoul
PGBR2jNBwvrcSGmODaUztY7JXgmfzAoL66+QGZrHz4Q7LDY+ziZEWCGrnOTF5F8M
W6shSeSjfDAAwcMc/x29tkFwbL741gtBdoZ8SdwJfJEEWLfH4osgg8V+MrGski/D
NqJhW9U9JEheDuoDkY52oZLqm/O2Oe4HIJXJpir4RGoUGeH36jcwieQi3zqSq5iU
/9FdWmvMTSiZrHFEjWy4thlSm8o56WnRy2Jom7jYK0STPb9v8NCSFkJQam407+Wd
wxdQAdA51hxc271R53vRy8uIz1/480Q7GTRV/135PXCGAYGHC/RslC7ce60nC88H
TdbHISXQ5S6yRjbqx7ivDLszpqPf6CYVimfGNz6LdKmQh5UDsP8nkWQkudlEXrdq
cHNgCeiR6F5afuhTr0gi/GnRfyWFvISqPROr19baFK7CS5/uA1cUBPkGB5PJ84bX
XF1tMeHHQ2LVHcIKrM/+ltvHyRWwoSIQHOXXhipbtezSaEXlf37HJHx03AToFch5
BFjipxkNiY7CdYNpBzLm18zpn2sa0ZQ3Pa3xp/8wKYi/pgQyHo2HcbwzfkWzlhAR
R+A7vFJchY53qeQWscI1U731z2kSzLnRhjOCMuAB8lbnEww1W5lUVoBX8pJvcdEa
zSQxPN7KjP9+bl8dr0orseHM3Eo8HTCTFGXSxdrY6MPZ8lU6wfTP7Z7dzjkwWKfg
vIyX/1m7UvtmTUn+oEuAQKkHEunrpOOnQaUCOtYSYlh1lKjB066yvHaa/Z8pV0qR
zYkj2qcAqnG09u+Wjucl8Ic/xsrJmu88b2XNnNT7PoUT4wivTrlveXw9n0/dDOI8
CK/iYqgwFSEmOIN7QK4u8RSFw0BzbLLvnpujdgxiamocLLnAcwLTvg3Vi3ILvO4Z
eR0bY2GuWwVWOjw7MNeb+ZzSUiNcso+LCosPwYi7UnZSyKH1q/4RLQ89fXKtp7E2
8U4wviUVn4SxuZFGVlDku9ooLUSy6UDeqrVxmGq4Nc4Bv9WHqSmE50cRSr2eKR/8
enZN9ZN4Vjs9J/51xF4tZd9D6RIlnK/PdIxUSXAFls3SHSPtxSWcRANwccEj3PMk
qWM347ypvEFg6/1JQez1ERiHZzOB3zACOyptp99YRd573DrZnBiORyxFJHT1FZVv
Ra1Jc+0/mLf2VxpdN5yQYzRCR1h7A9AFUYsEJNFS2H0j1+vAqDy6rZAxkea6umW3
3hUkN7d6CqaLNVWQIOO4hrhcG94jaS4fyBGLxeFIArWZx8BWRqyl7bD9H9wy3+Q1
Pxj6GbGMO1ItGr+lblaH99GsYiSBUyHWTPF6gDpUQQPYtc16B37Nx0cVkrIlOYCU
k04DWuDAb6kYQ6JGUQPKtBUuuU1RZK/Zvwzgs+vwCNsQ58tt3TCn/SCWtxPGnu4H
1sF2+jlIUOIThjSUmtlKZaU3/LLjg5ZAgMLxDbPxcrroDll/w5fj7z86A3MQ0e7p
ff9ZmJJqSFDwOhauqOEKAchCn53yAdzq+CWsgm5HntwT4sjTbVNrGbyaGLnHX47C
CPnJB+M0fzBo589Buyvp73Sgb/37km5lmNzaroucOqHvn+JhkLWxc0g8ubQe72Vr
ua+JOvLBXvJR+dOPgTFLPb8fI8cvz7mXXYmxmwK5k+49tdMQxZOwOAKAf9oCNAJG
teK0lK8k1mtwIwI2nTssZdEnnwFzzDPRmbtAK1J84EgrcJyUINA0S+SP14y7mhwH
HWrAy2Iifw9tFwdTmQQv68NKS90cva4LkFlgMGiY/iXMkMrQzFs8VHvaUqAbyIA2
XWzc290v13vhvL7reCHR5hIkjLkpMkFgIbY+El+oZYthUjCM6RYsSp5wm1RMrIrl
Q8WUJFO+IbBApNkZMPfRrb/YE+BfKluQXpR4KYyTSf+OUtMT9x14L3sOiPIciumo
rlKSk6hfMgrXFL8S/TjswQwV+hWCpqo3VvXe5kl2geSQlvWuoJrLM/ErYV/uLAEL
h4cwygonZGQt8fA+khJF2u11A0lyusb+tw5/t+cA61CLdXeYMVno0Pul5M/GnRT9
+5wLO7F9rRBXTPIkfgafuxFOXrH2+np3zpZcqrz6/eoWldlmEtXBg67bB6wCq0MY
Wkym2yQRP47tFaSp54eyvuUgot8LtrG4lzEswjA/8mVO8vyTwFqI8b+bpUHiEncP
1llEWpWQBsWxg4iT7m/NGnQGHR/vVBMZ5B5UaWcfb8ryCR0GfG+lmLn+qm+E28e5
mC4xM1tDOR0pnHuZOtmYm3lkmFlch3L4Bo7TOqreeqzQmrw7wlfSp2uzGsfV+UHV
CeSox9ASAkIG5vuUlh2P+2BtCCQ256e3N7a71kpUy5cfRZqgbXgEWtA/lCVyAQZC
VsoyFWLY6AvuRzY7YwBjyml5xog0dCSbjTvQwFlxsRqwXZ37WGAQJ9KB1mozAZ04
Yu2lyByVE9COFI94vcAsMjrcPsHEWkFgq0mjXZ2r3Fp4VmuH66WPv96fF4pcxZh7
+azvVrIdt3newkYVxO/ZNzhMZqIj+DKO0UiwGzxj7+kHiefUDecSpO2Tv/GcqoLO
nv1SqWSIMLAMUEkcVRVBJepbsST2vm62gdMOZrgUsaN52/5RPeKq3MZgvmDVr6WW
nT+nDcjbDwrEq8agAqjTNIMfbrHkF33d+dFhMjMVP4xKTtrU5dMDoYRxF2fH7NnR
XICi970Y4m7ctIuwD0eGjZg+u+D1Wqo4aIXtSGWb4OTJihn/uRCMM2owZWCle97D
vNWvgbBtIotJ7B5lG4sSQo6TXpgp/2fvhWUn2dvm90QGrYfJbfbiinPB9zqyhRz3
1PGVBHAz06svKiStWnDILFCacLOOlPDimXTionQqxfMG2SokbgxK0mf0bwlk78/G
DjBacSoDqTsk49SqXx72W7360Br24khnXFX272f9u2hRN0apfJik9Nhd8OQfVZ5W
cRnPxxIdENkAoiweytKkICcTy4kQ/qkKFdd7xS19VIwRmMScfV0VCUcYM6VKx0uS
qlDJPE6Mvj9++giJUVU7En7E51DU11xh5MzZJUwNphyy7NqanBHxI6kjBvxOQgx9
gbWCaAExKO8wLa4TMcv/+bqGPEwnfzDPoxPWtSP6phMMC1aEoLdoIXoxrummltKT
HkJVZRnYKkxNJC+hY9iaQYjYQBhx0ZevdER6EOJkUjn3NLaka/YGGV9c8KgAgZ1V
1z18fktl0Mv4TqxB4DcDZkEyTVpKffEAttFJdoI+nQwS1c5lbz4S6Sy0dh17EYWV
BM/cfnqYBAfFOCwA8QJ0P+he6qqWmt4ALMjFREmW1hq7wFMbMbboaJQZrfaZ1JN1
1AmDsdLePzzer1ZeXM2j+ezCWvEQRJuugWsGDT/TkgFXDl0/C5cDT5xGe21MnmJ7
4fYfSVVjgX3etR9yNAxZZcnnLXkzyIowHjV9xu4nnzn68HVcDkxG1X8cr/J/M8w8
T5m9zApMcPKGnVzco9JWrCm91oEzaEJMoAo1UE7KzrCX8vmBvjklq/DpXRvTs3lL
ypjUS1e5V4bfrAYtQwUv24ymDWsnw4oT5AF3wnXuSde4kGT5RAAx0mqUaFPUPARe
tBOahEg4p3bfaA6uQZgrRsel0BT76GgL6mtPLZAvmEgvJNUvuF7nhN16j9CpLWgS
IuGPdzDYECe2zAU2AdieyeUQv5Vo/6N8ZVFuOGkZa3F2tfOGL3XpGAamAej28mDQ
aScddhTgCdFquTsENvFK2p0h+5R/LRltxnsg4qITE5n+GSw+Hpx35eg8m3pP7VnZ
kVc1utGGZOPIYbez0dDhwOum8L5Q4OLU1Ub7tl+E09dkQaGvB3A4DLHKw0jCyccE
3Rca3PRYFbUV5xYuTzsl6e53pGFK/0zV7A+tSi0FcLsbZSkkL88vnL9MzxhlDJKN
5JSg2l1hIXbDd4Mkyme5Z/tLlkaeendLPG3MZi/7Rgb57CiZN/1k/74OH+fzo3aW
Rd3/qCSYyhQeX8sz2oBSNmbJ8x4xdhqkyWP75aNXHUYTpNRRvF6vCaDuGnpl78ye
lZyXvIL2GHYXE5LG6tu1BEX2DImMa3C1aEIvQrRTulf5a8AcYlUISJwKnl7sjA1J
at5TBmiBZ27oYWrNFNsO0u04R38wMHkN1IfdZGQqfccCeWs8uJmgKxf3WSAxdHqB
37izbaxUFIzVn3MID7NWv7LhKzfpAfJs6u/CMVKazPpIcryYpWDBurq12PtmqtIt
JehiNWqHRB6347gZxl8OKIu1iohOFt5wTTSXkhtXLyivFEHk/ZO1b4iJ1w4C5NYS
wyXnsq+Tos/IdUP5zRqZ0ymSRyFTkIh1PrVP8pTRzgDkiWi1TCdSv+SmC0nX4Y7r
7CvY1eBM0GyuC5kaa3l/xxA0MPnZvtJWevMQwl96mwMmmw+UkCYGeEzYohBdUcNO
Z+756UvEwVqd2EgMIF9S2OBCIVglYqh63x3UQEVGpYy9lDgiOw1P4K2IYf895cNg
Dd5wzPtJE2kcUvF4bmzhh8GsXrQKT2KEgBeC44DghrEibe4rRG6sGk/oqQd3DaOE
fDtoVF5zJvU9yhEur/3xVOciR8QZlEFgKvIYNRFCBypClV+sLwQcgWkuMmwF7mwY
PqQiFCyhUe1TzOIBZ2CbeI9/cfkQVE64b9ofzsW0LQeB3FCjNEjLcP9H8mcxMByg
gkfVM3tVMx4S2LBoUEBI3TcdT9QnD4LQFerj1O9/5d364hcVYp/EOOSdZDxaCUsU
i64fVN5YdYfCzWyYj1J1FBn7dsuEzN3Sc3UXqoJBmn3qvzk6dc9bEM/DLvTgqnQU
3+ydmEy6upxzXSbq+cNqs8PDb1a/tHCbOtx+jyf5M3wTtKJrhFXHbOl5NRChgZua
rtm6uL/JiiE5cbZEprbKDJJqa+npRyEKrhXXacbe3GBvx7Qnfnme5MF22Ye2wchv
A2wJHabVagv5cgEHoUrrNlgxGQBU9SE88wPcP+exdKAmaTVMmPyFrj8wmuZ/2EG8
j+MwfkthV6B7kGA9ViECtJQDI5++JNjEaa3FH5N6egm0CVOn+l5e5NGWCCKJiEuZ
aqn11NyVCyhs2YZllrBmNcWM5CWFpxK0jWpZlkZ8h0o38SquPLyM6OHv9PgswCFX
xfZVycLsw/UfK2IUwmTtHQlJNW7gY5lYNlxB5IbRcM/NeMetvbYdBHocgFVOeuro
Jg8SxT8KNmDBMJsdwbVI8K3QKfVMFXqyuGjihwy3ynsvYs5uDJmmEKyuZlkipmJ2
zdrQp3D7N7hl5yXnPjThoyufiFA0WAelE+XyvstFFhe+179RAvgqGAzOMNTovSlu
QvTp38G3eGsH1hH+IoZ/fpi88eLXwTD5ErFbBD8vEUCOwUA6uQqpd/TjvhyxLmUN
76nP/a6fIJUOv3ver/W2KBTutYy/4iiZj/mu4AV7pt0+AFcaN/ckpoMbmLWA/Kfw
8y025LOInKalnq/W9uP8aavApj7J1XGTpXzRh0sUwCh/Mjt2/QZ/DZwa5PjlWPc7
2gAOz1ryQhB7X1sFKAgE0UQpVdJG1FFgAS35bSVFKD8oJ1lrKpQc3J46nsx9MgM2
iMFn8pt3rUXwCogY6jsDcyBv2WIbxmNGsa02objH9R2uXElyi3QK5e4ngxMAlgHK
OpRcaADe0dh2iQ9vy69NC7KFmCVQb6Ydw6RegcT5j+2DAVc0jcTIUy/8m48rHGSZ
orJRU4mfGU0TBx6QQOfk02An5gHsUci7oWDu2Oo/eL34aZ0imBRPeaUZkz/Y8Umc
uE/do6RQWtchkAigL8tZ4zWGKrAc2VfJknyfNJVWYwYSfP8ezapctfj5taOqjowk
gQytqawq3hg0pDK2kM9dth08I8HdYTFYMwaMPV3EZmGpd6PGUcXkJnPvTdimaUcH
x4oSoJ+OCTDDqbDkBPWn2y7fObTn4vZc+vXE4Cuqdp09Hmwd2JcIr4Zsxy3B71xI
ajPY78vHO17CbP8ywh/fCvgHEB8PRdp2E/2+vGJCfHOjmIHkK7YFJ0Al3U+3XFdV
+ld0Hb0+z4qWsdWXtElJukb8t2JOzMyO2NTdbj5v+Er6BYST+MBKI5hhM5bsOBhM
yphpIpzuJ6WIMD12dIcxofV17/RUaxR6ip5Z4W+uLcAskufgcTXN1GqKKEYcvFGe
M9G1jNxUUp+ffw2DzHLLSxWOUpfCELreOzJrusoRZYeePcP9uzZy3yixdLw2Ii4i
D2o35WTkVu5CjONbneTzgo/W3NLPEMYlmZkUAWXY070JtkELAZzfCDergCGGazwX
oJPHMe8x3EZ/FyHriF47DPpeBSFLIapSmDiOnYhkqBCeT4FbGylJbMPsBhF8E4is
8WSFY2Sg/LSZWZf6T7w8F0PII6tDwYjQySs5mtevElU1eRaMloOTENROKdwpHW74
ebTzYCb4SuKjciV5qFUqmbSe+MA8os/Rbvl9XUsummtH0f2ZC2+Kth3dWh1NiGUu
PnCMxPKTl/ofLJFAhHNnuGeF2J3OG5EQvDytFOk8I3mI8Oxpf7hn4Uhx18CFILL0
rIKDvf3x0SZCqNTl6wYMEHrj0R3OVtT3LuESftGfpKFAACCfPQZu0jpKBA9OrRsn
0Vv9FBd+7wpHwVJ0qMfrbuS4vdP+S+EarL6+TfizB7IM6KRvO/oxD5HVSyG1Vtw2
VYL2v/W7t2fIWlNoEV/K+0zmxfDxOB9bKiUnQ30fjyisjsH0i/GBvGdYrF4BJpda
vPhJ/lZ6N4VxcwZpTKuWYqYkvFh5h1CmPL1dLDusgfCu6ZwUq+xgzPwsY8F7iPhQ
f8uYqcBXWVX5iZ8wPmPqrbRYUXNSTwuW4oSmmEuDxcKLCt3AxRnZ7yj/yMdwTdZr
I8L5WONZCgHinrcxIcqFUssLufs6b8u1gRPApB5Uke2beuYPgji0MgdfIftM4hFP
AlVs7Nfxac4n+pqlTr19KvIWb/Vg8igNfOoNIffurdS/uIZOLY63UA/atdGBCJG4
XrH62dT8rk90LStQPvpwhLUSYGsp1n6GPcWuonVnFnJVSBnI1CsaXee0nS6NrrND
uafGLuh+fhzHfn8bwdfsO2gDFF3JfNaiH1Yr3NlhknlHwwJSeUWsHpHh3uoaAJop
JmDJxNKFaktEfqQ2GvjxITHEMIoDItr8H77pKpL6GWQ5hl+CmYlPqJCDylPvNuWZ
e1sRl41pduZVJZO+UjqMQy4HSYvXW9FtU4qVXSPcR163BLBqVrdddP9oRTaO8Pf5
piLG8n8tyOyLY839N4NsKNOllkGNgF5tbl8xoJbtfGwhUdjq7xTUVSKk0lrr2EHQ
oneEkpy2HE7EciEpNdWwMbOJkn2GyjozZlsbeSm0mOg64P/FOH5XVwjNL0TNLsk2
r0+XZp1rBMHgyD+zXMNoXEpDmsgdJ5Vys3Np64HsZyywc9h67GDWqpdUiz4slbyj
nx94PApKMdul8Dsr9iss2elMTh/DyQazMtWu6FXzpv79/lulyX1BibciVPZh0rVz
V4HbX17paKQbTePiWFKzt5/lCIShOE9Z3oixHQ1BXWcFoFmOlYixaQU5e+IisGgZ
pWY7atSHvuvlny2bO76/DKtPUIq3UYSr+zIEUDH+RRWkviHs69g5VD4NK3qpwJTI
wyeCJN+c3GQbIL8BOS+3PVLyflS22E/PePHJ9O5e9FVLx92CEJ7w7FFUh6pFZSzG
5hNsupHgGqaRRepfhzCZ6ftU5kkdi/aKnB7VbQ8DKcLkMFYChXs1oor3fIXhYZlt
mYv7Ku9rHNoczNHdCgzEZ12uBrkBZk+1aTXyIqzhG+1VZ2VZBBEGQDntp1vB732f
Dd9HWeJSJ1e3045EjE2UWeVPLc8umpy3mLduSkH2J2pllsBDjr296u+k4oPVXT2t
KIEP87CzqsN+UZNSL2V8m03CJGWW3kJ4fpYz+kLKdV2XoQ7PvhcT4kp0pxH1bgIP
BSIjNo7tU7v11/IZIdwhiRlseouhqXTKvxyXas9+K7zBtFMSNCCcgT3kIOeDT3Uz
ppyLzPnQBlcZ3N8RrgHDuWAZXeCqakKFEJNCfxfGSLcEL5RgnMyXLDoJhH9ow+n0
r3Raz+uCQZgIP2hJavLlEUEDso6fFgx/gVWnfyN687HiIoQaOYSc2aFgiC/EyI1Y
mif5i24QZ3Ir6QHymGP5Hnqv1hrl4mpF9vH5nN2bhJtmMrxgT091LpcVKGAKGgJB
1UPY/kOz9vH6FYXdcHiR7SOgiGq2fUdVd67geM0N0ioeRnqB0lGcg9sjcdOexOe8
V1dWFM49aCWhOIAPVZUy5DlIa29IXuCy3XhJxK0XDDJuCO4xxKZQ9qiBBEnVpB6Y
bepUOhKIb2DK/HI66dUaLdF5GVU5Rslh2HXSEBrW5MPGYNkk+pJJ/qpwxS2y4Ybc
evUNi0U8nk8aa7TPXzWePOjnFZc+E7AXYXk5Wjm1fE01d8AD5L0mQ/1j3AHKZiHE
8mBGtYo/R0lXRIYgRA4izXT0dAIQx7PggHv9FAcc+/H94EY4rbDQMHANL6/twEQx
PjFZntMNLih8Z77kVlctX6lywalYnEmSLkP2ORb4Sk4BFM1QMHI/dB5qQThHimbs
CtWLoktV+iaDBf2iq1ioKuosZYHOrwxEGZh7QXjyHGRNLeQYLoW1OGXxhzBk+uOj
Fq2h4lS2oHJVr9JP7B9F+ag9mm6zl8kVdkSo3RiYpKqvsdy4gfF2bcU0FoZoNBd1
OPupbXfEmxaF2Zs+11w2KUaUerb/TdrIqro87Zx70uSpJWNgP3i6sLWHmsdIsNLp
hFUrDwrz3Sy0i9IdRSdYH0hqFUPsd2ODG2nSYNIuFhJGAkuIfJMF3wYUf1OGnGC2
qBFhEsClikriGzy1zXVAvsVeR12F+yXs3dLv8mgLxQ2E5tZcay8CCbCY8ER/f3M1
LV+E2ie5OOAHfyaf5k4HATLcA0ic0oaP49QVNfLN8eXW3KyMxixzi8x4PjduH/Wb
WweWfSlPy5Svy1uRNTRHOX3imv/9MvVpnkJ1wH0gHJwOz8HIPJb0p1wODlsNnZ5c
TPSzHXBHOd8JZfzMRSg4pBgufOI5/3DfJQIi5VpIrFiwq6ltw0uGHliPbNT6Fe0C
lFMeDlJYJQimKDQZ8S/RdGkqjaQfr3uy+4iWvr8WMOI4utqrgD1As8Uj9rU8/fy1
Q67mKVj2e/tkYiqViMILPcNpSrDvvdeOeb//6ZiOfGg/vMoEaqh0pQpAdFKxJ9z6
UBABDmJp06FoQuLRApVIN0EbIA79R6PwDJgmFBpB4h1PIwCrdRkTwkvxL+R3Pp4O
lperPeSWBV/rzTQRH3sGDuOyCLfarUFUavLLnRZLqk2vbV8zOxipi9LOE62x8WDN
UWQR78Jg9jh7mrkNO2Ca6Jd2rCP+ga+/QcEQyKmJsqmx+WAeYIl62XdIxW3Kee9m
YBCleDs30Fs+uJsCt9MJxGteHtZpb58vQgLrH4EV6ZOHnnRJKmxtvVuDBFZFTxNp
gFqYlxGN47KRzyHCuMFQIkngpxYS1/2p+G/moARgKgL/KcVmGA8daF6cknk3FriG
ghc570a0IbM7aO+kFvo/3wfEfufOD8jxCIcEO1R12kz39fXhFDyXYzqJQiYmrC5L
AltzY7X/I4hlAhtuM1QoMWbUUxYRfC9MYWZdH+GIqWEyV2v0Yu0VDMpWlcGdV64W
Q2h/ghxprjhoIIXLq7JdKijewtwGvPC4KPxjYxNtHE9bMCg8cJJ2ROFX77GSmN3m
WzXDOdT7qKUKeqQm2DlaM42c7A9oetWRTk98PK0Fua4MPH3naIURKYFfNxubVDtG
JyhHY3Rjy05dVMagxVYr8Aq3JZf/bubd+Cd5QVMrSweNHOeUtMU02Sbj5QfSekhX
Z4agZuo7kqZa0IdD43ztuFr7zwq5Cd819hMnLC8akYmkJN6yE1sAjurxihL+CDSr
bCZTe35KqpRohIZFgr1Qe+TG4NX+8hsP1Dd00W3H1CsdOZxBp/4SFnyd/xMse97C
CrKQj6ZOzUsnUQw3pz8pZ2nQSbbV5jFpYySm5RyI4fyDICRHL2ce6qUX7oWtPJbf
wj9cD82B+Zy+PQRFHez88PAg+qLSH1H4bpbfk62vNplfA3+QaxqiBuQ97IaAdS+O
y7zTOtecGETkDOhPxqsnv2e63WOosIxe8It3nwm8bdwTDICZ5MxqQyynJnRIPDl6
1FQwCP9kkcXeE8gkT40P3pYLqcoVDKL6OR6uzIiNP7ULabgBcX6q++vt9m1uyel+
HMwjedMTRq2ectU+kSDWMp9M/qU8AhsFHuSXQ3wQmPy0CMohHuL4U7E0tGxryBGk
z13nij0yIsD39dA+awHNZL0eqeFGfS/+W5yhTZSNXabzb2pO/VUIg0JTsM/jOCDD
UyW73AsmNPU4shXBUVgJgdKombyO2HDrHu+B+dbO8ZwlVQWmquhbSxpwVqtvopQh
3uF5/mGkc9n7fh9mRGMFWCPBSX3j17nmkNfh9Y2j3xdG3dBXlVCpIA7Em2u5EbO3
vvZy/2HuWYHddPuAnYoGec/tGR0k8PH5abgqMHJxV94w573dOOBnfQse6rEMxVYn
q0FFKSJ/OMsIEvAwCSuUW0Ky2NZUmWIdncPEXDjl3DNTBHTbx5Q9pvYs87Oz9v2+
N/WCf7li4p5p9YozmwSoZ3MeALmHZ5YkHO9XrwOez4yxJCkcUE6DPKtIEzPz+hmA
/5j8JO7nfIvo/CdjDcJFb+Q69mWLRG6l/TtPG85onOkq+oXdztfPWBDiiS8Z1H4n
Jws9vlhRQeBhmrOm4aPaswq5Campyoy5bv/I30A72S4D3vUv/CfSfnz0POAfjTrw
yyUSm+DLJFKHLcyplaIurQDW4ch/S6vcSktGL0QLO3zEtiwC63V3G3k9whKsIMJY
PzzGZ4Z474C3jkYM6alilOaTv+KRsTvPY7BZG5eYdEuoktpA+pDxOPnokZ1CxTtD
5ZWrZATA4SGowF8aOdbi24SUjEyYeFWsIsDGDk7m0+Kte9Ym29mqG+J//D23OyGU
taW5HKFAkEtYeaRwaSZ8n88maXhXLUamDjU1LeZDMZpVdIYt0117dG/aoD6fzJO+
f6h9Yk4dGSSOg0XCCxeKfpXacFi1MDYViyEJq/uFc3w/WJoIOgmL/WYl8g7UV58U
9mP+3BmyS9qDJvuP+rV83vsm8sh07ylFSWYDXmJps1T4AhY/RmiQ9Yrh46v7U6AY
cXAjRJbS3Pow3PZ2d7kJslsyavjpCxv8S0igwUdsbD+RDVSpvXr83HdsKvCFYEEZ
eoHUjlU38H6L/yXpcmPMROUt1CKsTFP8AN8qUdfO7146wx7Vopf8HjemjTF6cyTw
Ml/Szl8DpbBnXND79aqA0yKMJUQOv1CUdOvSBhZLqL7GIaMn9XpbmUAxZ7dKVkIq
gumLBny/mjiaHopIejINVU28wX+7HBYXPznSBUt4GB4yhK55q8pwj7h4Ot4LclEq
+X7VpK+10rFWy03VhjtXwS7rbs8AaodspyNX9GmCauMIT+AYlTM/v8g3xwXZ6/fV
vKELUFH3ihfCprSOvma7GYopGtzzsORtx0v0KxLa2LqHcoyFfxYUrGOdUk8s9aUn
/3rKMEUhImwWIXWFICAaUWkNdTOxXUDO7EJOVILnrRf2tol+LdTuznn0toLTpmvm
YkJ8NPkQneZDBjtOWJPbR8iJYwh+RZvrQxQCzfoKIpJfPbCEt7eAanYK82c0xzAo
3KHHW1qH6lPefozd4wab6Uyk1jUjoGOXMn1vnrNdRkKAU5Z4Op1VXVjZCc9sAToJ
F6fouArZ6ID7tqoBpMLVT2jubSf9DaDMpr7fsmahNpJboOkHEU08s8O3KIAg5GQn
CwEc1Pp38cvJEmyuMfTF8zYhhYkc/eY4bA2n0ruocZdXAHt/6oe3FsJv7d6ouL3w
rmSZRzBsltZwAzpVX6gjbwPbE9CtycELm7oEwmWLumPJar9MFtoiVcRTf56+372i
bhUHGcd9fqoRXQB7wxy2T3SoL6Lru/snIl4khN8NbDhEkQmNM58n94hMS3uIMfmk
rPmT9Yd3RZDngcEbg0bAvyurQMZch9zcSUWIWIUGYv8Sg8ToAG1X5V+Nqb4nmlJ5
vYVJPt2znvlZUmRlPM6qxHIPEYz6GZzmW77liEVGUk/U6dif/fWH2fiRSykVffBg
jNdP43V3nwdHbQ3tcFDyVFwHj9z06flNOdeQdF14Qf36xfsVlaEKp+iL1uIcnb0Q
R9Pb7zOs/rO2E5/QtiaAYIeosCs202+NFpwx6Vng8oaTuWEnwW89Ig/JzG3h9v5I
zj7HS5J9MTQdle02REbiLF4D4hyrAvroqGMTMKG3PWkFJuW9/8CjZVIXAfs96aW4
g2mWsq6Tj8uM5okaeSj4B2Xl9CFGCxa2gjpLspzBgHm+s9UxP7UuekPnh2okT9R+
PZngcqMavugOckZRfKxmyR1evYu9Oj7D0g/ao1bZExTG3Hou//viAfqf3B7/pu+t
kZuhVbdj+hjpnKE5+TvoE3pQOEh/h28aQ8rOyUeHYf2I9OAi6+YaeA5U4Vqb6JYU
zeVI6qmwDRhNUQsrSmjEYQufDFoguYMr7B4pNl0/eN2wm1pjt0H8ytFHdS/WRLYI
EP7JCwERKQfNz4MxYgek9ZpG2qDNL9mlBJcBcK6jEYU0tByTEUYx7zNRPJ5oSXig
aIlU62FlM8cMctpfM4qIfMEgPNDu3Zeh6okyhMk6jT3E47CDqc4i0dABEgSKbBZp
rW6135WG6aqQIlM444JKDRPUIWLqwV7FpKPBQ69RI7ghfcIbT08hbg5/DnEnJUcU
EUdNsXfU12P74Ncfe6wlQ9xxWZxSDAP+iLtaA698JkrbuqGV/5vFcNoCKDEXmsNj
gpus4zOVzXnZHJmajMUWXZTIGFvzJ67qX1lgRrvmoBF+vs42/dQhIlQwxuEEuSE2
dvuf78cA9cgiW/aSIp5GtViYPVcKMoEDrOV+gF30Yq8/QUtXjT1nvbv8bloF+syL
EJakB2xFCVAh7dr8+4DVkHY6Slrdu2kO3NqnvOD7t9105mfL8cNwVJHaM/aWlPp3
skJJ0EQgYiN0HJFDZHd4TWqWykyEiwZjkjS4F0kq8pJzInlYcAPzeS6YWKQcHHth
0GOsHE9HJYls7TSPjgL0lwO/LYkRNC/4k5IfKNvoZjSHIBlDZbiu/mayG57+FA1g
gb54BA9rVA1jwg8rjdGAkX5eJjD9uFi6HCA6d6/JUq5ChpFgPBy2R9oSd2TvRctA
tf0eUgq4VcofM5DX2CKlXwmIgPBbHmmZUo/MiNfkvP4APIgGH4zZzS1AaxvfieKD
I5QCryN8RWD/wRjtMsUmUpB+gvOniUOcaR/Ajjx2nH3vsqulZZ5hNX3JNTEME130
36Z5rjomr8LQZj5UpW6dEhuB0dnuV6IIT9vnJX0WKX2NI0ERHm3U5EE8N3eHyqsP
WlcmG7B7IOEC3kSKol1Kq3bG/TaQP2HUijW6qXToDxdHPby1HJ4OE/eguuWi/Wya
GUP0hyy3T+TR9dtGqKCWrzbW0QZDJ/H1IITfNmdBQQeVhhhbNHl/5DOI68bLUYvJ
TTPx8Dr4ix0KhdR2GE+D9YiSu6p7z7zN4m/wYGUhr2obX2ZkQBqZBuhnaD2f/VDA
2WhjpEObdlip8gszuu5Ct/gQg0GINNBGzuWEjb79GbURuY+TlNXQzh3LkcEHwRY8
SB6nrA5/1jGSYuDOifK4P6rria3Tdp7vX9oQfCJqT2Dlo1LHeof/H+Pni25X3ICJ
Saq2nR/rYTXH8nOqJzZIzNVvG35lquwgfeZleBSjrFS1hjZnABiN6v9l0Nfa+Ef6
tvxiJgfZB7R1jzBW71Um+Ay1ILKxbPYDrqkGkK9BcN54l8PeNtobBL0bmEwxFrOh
/SPzuelZ/UHZxFBHjcxH1+OAQQVkqLX9TpzBuDHLdtpZ8MJEy94y1BN1Y3SyAmTX
Q9wKrR4p/3uc+S0QxTgCK0ZB8W6V23NRzjsE4LGJpWFJGqHKPxePkKzbQP7DI2yw
xS4J+WsrGAQlTttckbEHP7eYK2sHKLctym/0oLaJPyrQ2EA3BfGpNGai2ETaxx9V
3hbY8m4pq2Ycjd1epLPlnc9+T6ALsQJqPnSukOCV2HCWTuSTmSSUKISSEKKiLgOz
xAv1A0y4aKbxf+GPpAZvO9ncfmr+eBS5af8B2A76GY+eg0R4Q4QWWt2P/HqBhzps
xlzZm4rcXV9jaSZj5trxx+nTJO50BO6FXU2N9F9ESgviuvFUk8yaViYG26A49G4U
+QJ5+NoUCoUgYYns69zzamOP2p7nMRYVCpDP5J3w0Z/C+lwzculCEBca/onK2Krd
Uvc5LNt7ZkGxxbTK1SUam4PIsmT9OvflNtcOA3eMA9z/peNo9f6dytQ+vQ4sYSCr
MMoeef+zHMHNQY0A+ZT/fqXUgp2/mfCQ9o8vah85RQ6a2j27zGxmH3rMIJjwrf4a
tOSk6O89NI4HQWy+hzKme2fvN0Qfc/BGFrhBlzeAy2fZX8IdiLwcPSmhpmyVL6Av
YEMhZ+wHkR9RTD0HkhqkuFQTBkewm7Al41n9MyZ9M9ULNHaEWeLsqA4bB83Cr5AA
adlpxaIv7c9A2aYDw+rXqEabnW9rksZ2XcSQ3sBTJIuF5ng/7vNHdViDUzMGnwqB
WKT4X5oB/lgFQbfG6ZMalkkJCzK5ASb2WcDGOahA+K9HI5AH8RSmaiWeLDI1BNOH
pZR8zAA7tz8zUkBy5uAmd5PAWFQ5UzlqXY8jo+Vf+mpiDNMh1Mlnin3vRRjXBEVP
OPupiutkyjbe0Kk7rdOGV6a5bi6MWtqEtKKyliDbSrzRPRCIRKqOhBLM6JN4ydl5
9hjG13hnOzXgdnTnn+T4ZnSPgwir3Adml4/nXfpOZx9YM5VxeijFMEgjiF7SqGat
Ve+0HHxWDx03QGMpk71HqCWcQTvexsgZOq9Gs6aV2XKd5fInKwnK9PKDu+01qaXR
bMfcqwb70nYyaUwZnzCTAkDwjs7UA2qcyzGc+4257H85TePgpzz03yyMP5LrWswB
oNTcHak/I+EL5VKTugl0WBleo8JcVwh0xMyb3H3a023xvvrZvhpCmpQsyN/Hp9wL
pKNA6wB1vdaTTeOhjajON7k2Amm75wyRqjE27FJOurvl4gZ0wjqwoiRc6yUciI1E
tdkRJFfROwUh+WyIBQopZHIIixO8NSHXDSvV2CBiEcvmAmFtRGFG6vaD4BRtkUC2
v1zeS89voeA3ObE/BsSYrCAHM6hKxX4dlm49XKqvjLil8qZUSEU1GkUz9ts7NdY8
lMW3ATHU5ppbo7sxct6QPy3HkuSvk1cIwk6qLPs4LsOYoHhliUMALVNvFB8+II5n
zIZ01qoxJsERH+yhzdb0m3KIPZLE4YpWX0dgLA6erKIObFducdqWDVvmqn8omZSV
ryyL4DwAhJdm5KJ72kd6nu/rhgRBvAROvYHNlCqlWUX38X7xhM/TRjEjYDgxw93b
CEtPtFtR2LFdjmRkd3l3+j729pr6INqSTII98R0A/5M+TUeC1HxfsejBdA+pJdkT
jKnhV+EIzFITogVWOX3BfNj7mi6I4VXt+hKfREp1j1TlVu4EWZilf8lwKNLm0b8h
S3a3H9Cz+WxwdPanckuiVZTV785iCsL9ZldTwSm/kdLLlV9AtgVlVxWDOIJZ9Luy
H+FChaJGRJSbVa+suPnR0U94m72c/ifpl9vgGwogSiqZWXBpBhGJTJ0cBqU3lquz
iYWkPqO9aKVr5OeIVxy5WtF9b3cHA8qsSFXFbwnwOZcgiOA/PX4vmzgtCog/Tg0O
hRYYmA96GWN7RlF3CCj+ArsQUpSKYYYral9NhufjBXK8VinPLOixNYpC9MYO3N3q
rn4sRGODquFFsd9Xy0VlgnvL4Bm5cWFRyoPKECi6F3pKY9jJHjVGNfTpC7+6M/TM
q5VGROKxLP0ZpccZXyvkUk6rO+c6m7faCeS7kOIZno6Ya1/5aq2OeVBGFFXqKeGz
y6tJ9VTF+u/kQSaacYbbEfVGS+lUntIjyWEsFapjD42DLTuxfcTO+mxKC1G+d2zy
CIKda/rjMwFi1bl/ZslRuyJ/axdi+/Mtn2qpFkeP5ZvlpEEhrlZeE5akkIxBh2+t
BJvbtRL0JQ5mTdw0CNxd4YKBzbnWgZW8uJRSkk31ZE10zLzRWhduGvO3YzHxD/L2
CkzijJA2iGpi5p1/aXEdHIMLJQ6xLU3Ahn+Cige7eeaNgrcxs9iaV3QpBJxwQh8D
tdINcL2pPuu0fC0cL0kDIElrbjfC4LA7yVjOnaslGXVh8Yf/vHVSks2cTZ0FrI7X
Hp+ZKlt2Wri4kzW2UVdWvEVyptmSlFH1OjXtlN8CBFVL8hr+//o35roFQ/vdjiCo
MAxze7wn09KXpAdVdTCJsvF1W0pPbPEVnm938q9MZYB6ykX7gyRdTXBDl3cGJ/d9
/2anG/QjhNokCJrAZ6lQnpj59L/GZpCPgoXf+Zsp9EQwSx7T9Xepo424tv+eGBYv
x2G1nbIPLX9lz/LmyOXrQsKHAIr48u6HY6DnNiATCTVZvLXTn8q9KGqTMLsBuQtf
Vlk35jr8lEUmfVJj9ATXeyvqtG3jizP0vOB8vhDdzinDVvDjKgTveObMXbDKxroE
W6fWbsEBcCp8hN/kqK1yUareMyvvWntjlkCEd75DGezH7Lld8iphjnSOqOogTuCS
QQV9XdfI/Omg9Rep/bNgaaBd7oXFRcKXR2AxYXx15HOS/1wdqf6tfim55ue/Dt3h
JAbQXcErKJyszCgj6njmgL+fZ7XtSEPotrMDrIcHo1i0WTXY6LfH7GdFPV6pmPAL
FxzpRfEGbvxk+JESZWNeDoeuBMjf7a5h8KWunJKwv7UCCUkNBBuRIFTotSppo3Bq
wwue/B/Gj2L+J4lydNRtm8m9ptcCzOPp2p2pn045Mfvu+FPRZPyyIEFEFSsaikkA
h/PFCoh8V2XldXxGQpksxkhzCuE1VqMKN2L0jbuC3HU3TrRW/G9jU6P4NI4e4xLI
3qF7pP7nUmA8J403ceF90nuUJSjKeupZuWTCeYAGCiQleVYrgHexwUDTpTUGXLCL
uDAzcqhmA1srMW0CICfnc+v/VDO5y3qjjy/bTOCwmWvkNQro8ERmI505FM869SKP
Cz9NeaKYuSTTkxAhKh+3KprX3ZQxwVeGPCA5Pv3qqWLabIA5aUZLwrFatN5TftA+
AhL5QychT11BfW1QSIbUxTr6RW8zYjB17W7oOf+UoOazIt0af/hmGD9dgHZRpE+p
pPJEDmlwCwzmzmbYwDC8kSDzG3h6lHD7/R0r4qkTwW3SzJRxdwWA+hC+vVjc8Cgj
HRvdCpvFMAKwS1BoGOuJUQf+BbDkl7ROPJ5v4mJgKQiZ/B2Uar6gZnEVmoON/+DW
RNj2V3/m7rNKwCNCWjI8k2g3vQD75mb3xh4q0jdaLd6a2LQfe+0e12fQPgfUC5YO
mHVRhQiy0e4INfnG/xkVeYr6KHj7KGv5TfQpn76Ak5gp8xRfUUnb34QMIl0dd1wT
Vw8Lvgtv0TyhEII2+KwGYdgw1N6KhpSBranOjkT1L3PGPeNuWxEN5gLgXdQqJRG6
+GudbdrYvMagtq946zJB4N/jPvR9pXcuEGqse+6YYzWqPOTWUMHNitqUIADIBFJz
Gn7enim9Hqv4vlhZX1Pnrb8MtAPmiCUisoFRLROBP+KBfaumz4Yt2kP9tevIOQND
lmcsX9eG+3xLsCoB+RR1LeaLe5q122XRVR3XAt7DW0mTw8e4MgXtT/LSg0j+s1IW
EfsTmoFlvqNpc7aeprPR5JfNMIpYq0IR9YAiw2ugGsncNfvsPE/zvcyD/XM+vKeV
SDhJgpZO2G3hfM3pXg6EbtJshqmSlti/8xLwr+QoQqmoQ/B5gcMTlODU/1Qg4OiS
V2L9GBJx3/+HpYehvxMDMBBBqiwwZf8bSlcEn0APzCQ0wj4DDrUtdJL7HOUAwPys
vxVVsQs3kdxiaKHvDVLPGBbZuy2enWVH1Il+czR3nk6h+9rALqc8qtoxx4Qj7QC+
HgSW6rrTpQ39mT+2ahwI12SUWoXdYvvcjEYIhMf6Jtf6WGEJ2p49sujChjBGVLsS
VX9XlCIRp6GG73KojRGIgOI3kofhGUWKqmCLReCyquFiZ6sp+FcRQ3ud+24PU6EE
eLv9rgKR5gHGV6uebWL4o1UKtGuwtqto3FBvTcBJZ3qp9bVipx2s0qWO2ki5kaVN
Pzim39fAyvyvxrAKJ/hZP/+zdcF67WgCXY18lvjcV6q3hFi4uJqfCtyC6494C8hm
ZicAR8MJfu7O4f9yGB4/fhElUjqUnKA9zCfwnyKlXeK17XmOtbxZl5nD+SzzQEBb
lhaGotrti+5E+oyOP+6IX1Si3boQakKKWEX3gkh2plt3+kO0Zmq5h7ItLsLSiBnR
0WX/fH7qHK8nOCgMQdY0vza5/LiAh/UmupOwEqP7e4g4z58nRgcI1uwO7nF2gq7Y
ra0z8USqWrQ7o+o/+3K5FsX+AVbEDZL1DcZIUVk9w4HIvmrPvVQN6qaPLHgvh8cb
woQculjvVlRnPHxHr23cPQNS/5LlAOJ6nk1ns1GXnaOfoWfRArK1fRJDrv4uncI3
uTSWZEdkm7ZKDM7NTVjjCVXUDuAwikDMWxZIwCvKtlazCkL7bHDKXlgSfnT4vDu8
FRMT7iPYp1OjfAsSwwHMMad0oLQyxLArRw6FjI+r8CMPEoe5bZPLFnyipUURYZ5j
4fKSA7XjeJUG0GzeRH8DJfWUkmwyEPfDhjx18gOrqYFymDWh/Lc6lai3qmOOEFts
RpVVD5gVLFBAl6XffUO//KgmkXG4xMc7c61npH4FGxh/vEsdC6KyJF2LHpr1HnBC
G45aPT+Bz/qE5UeVZTA0minYsEKW6PBQN2oAeyQhgasyXbSY8w6xJF1XMyZ9TmP/
dHmr8lshjCCnt3XpfOLeGzAa/aqs4IKC4Ks0OtpIULjdslPpHkGnNRDpeUpOjwST
0UtL20rFL5e7NoEvPCrY+URHNMA9ZEMddOAC1TYBvxtHt5qawJYQz+NwJSX0jKJo
HZPntz/3B3prEdMh0o/GThLvfY+a3W+18dAv1GDLwIbOwp2+QKkV9Z04S7z6DptR
K0uLtS2qo2cZJlK2tons491BuSylfeYwN6pvwAy4zY4e/NfF+BJS2HJGHVvR9kOA
4h8lc2Z7a2ARem1zN8tWhf4b35m523f59YgItkOh3OoJK3t4bes+xqxbNHZVSl4O
9wxdi50apOll65HkRVBW2ccw0WHwiaT2tOAQPPUzRUAvHddX2iWEaYGQ4atFz66m
QRe1fMsoFn42o4drY+T/KK1qo+DcCo4EdZqrPTiv1b/tKo5Unh9ldZEwPBadcTpE
nVDtCGyU4LtbE8Z5TTDU0LQsussCUvhxR9c5BxRMZS29vsToRITKEyWPtMuAQ6vv
6LyxFq76KMiXzM0tqQkDEulIXpiHyhdaJDp7/NgelIRMU05wX5LmNz/m72cu4Ep4
MoXassncgF8ZrdSmFJkpfvhOuN0c/IqEFkFui1j443efSREdN4mRymyGfhqJ/0By
H8IG4SiCmm0L08O6aoho9JcVY8lbVHdU0cEeGUbxYNX9Vrs1Bby7z8KznHsm5pS/
Zv22ouNYrCfXDGdUT3A3pLvZNqhoO4/LsNyhCWmWl3/lblhCjgMTK+RQ5iU7BLbz
7nK48mwQkqge+CPh6pGQ5/64ypVBETGkCBZFc3PKjX2w3ua5hlQZKPktCMqPfyvZ
5ZBCYDMuXKOf+NckJ//BF1uO5laoy9nTi4u30TcMvFWma7NEQVH0fK7Mo1OhaxKr
ybVi5g4+kW7BtNQsQCyScCNcTewMcA9hOjBFyzfY3SKzRlqOmJw8MDa4k9JL2yVb
0klqsl1pETuwDTLFa4Tom0r4EGDsMgLgygbyDBUXudasmzFTN8UhhElwTThSHW8B
UctlXS2Vfeqb6qpKHgv1qz0ql60DM+1dZ5C8oeUaCH+hEJ68NzWbIhgIFkhfAd6X
/KcLWHqv5k2wLohCb7lXTT+i0+3pPgheWxNUvmnh4oii9D573Mzf6hpebMoSV/AI
d9okPbjiwLLn41gMdqi/0wsKQMWaOoP3XL79ixiE/3bsv6XA6YzBL6hiBrfccmbH
blH2hALqpGHJwFExHc73inQoIBtfq7Tjp3LecXYdQYBUaCeHqZ6t/7Ebh4M31pwG
cAgaZDnnYhEV42Af51NPLlsUgdY4AH/cfUvQlDsLZBaW3HdwlgmaMGXy4dxuSjJ8
nH75ZECxGPCCh4w8ZN/T2k5kScVdL8jCV6M9updvPFMHNVUF9Tw1L+UsOnY8a2Po
QYo6MjkSubWu89H32tyw3PIUClbLRPEyJ7YgcMOItAyCWs6uvqiKzBlYVPzrKaWz
XuQ8jc7wL1xqF7vkgf/PEbfr3l12vm/nTTc/cWALSYNVTbWr02sfxT6g0BF2IOi0
4vjPsvMp+uZo159p/eQboV+Kz5ldd/mWP62u4N6U95HSfuasrnaZCo2nA6rrlbbA
0vWWcgvdUPRMiMUabdJ7Q0O9Eo0gYV2WEpdEYIkDow5/HG2Gl20Ao9X1TlxR645s
RVmcA/DiwD87ky4zLQEj3jhBmUJL2zSbbRFlpT1DZwO4yO2mL51tCvFFUGisCVhb
pixYaGklT6CinnWzX5jMLMTNKrAy+0iCwSBVxIzMsShWcbB62AWyjzsfydVc6sHU
YpDkWgjZLeYKbqLqmCU27BwscpIlFxnY7RWPFsPSsQHy/+2JUB4WiVWs+5Glpl9F
Sb8gMUBgh7HqLiBRiEKm4x3m5UqaD5BIQLqoHlcyhuQV2E+kkiZ4sEwjnHcGvSCf
O5VH0j4FCgK10WM58o0UWFYRTYDxX6Qsp9g4I5OEXK2FAdwCLBmMncKpoWD+DoLq
u3EaBN3msbaFEJQfUCi5k4RZXmzgfhSQ/EQ77aAMVbirGLex8NdIEK0/AIAbXIgS
Ej1vAP21wELGBehBwPw1Eouhc+KDTJCovLej1JutuDXPDiBjlegA5bVOYH0s4g6d
Y57zCtbf1wIX/OGxFsRjV6I7/liRSCxCYbNcW0a2noAXhhzIaSVc8HB6PcQ8IBtq
sdcsAuxAQewMMUW45G7DXaGM46tSxBl4cLuwmFD+iomtClDkzELBkfHTJyjCUp4q
jDzyKBoMzLtG3wPRg2AcbvtaYlmWqz3gJ5bGQB2NBdPyX9kgWCihQ94QqROhWuWR
842howIgvY+CKHg37rFE0h35IdJafA3kIDOZQHUsYWrheAVN4ykTns5oitLg82VX
AmBRvOJc8dN6N1TFWivNNTvzRrWMxSB1vqpc0aKdmjnoZPNy+lZckaBC8By0Ro3b
usfg2KUz5jk7imu/vRqeLlupNTzTLNh9XkmFAIKXBbmivN15HC/aD1x4w83Z5DVD
gtTMYgGCTa5ucJifLYSykKqyUANtjoosUtHZxpIzx33B67iO6mejdopn8JfDT1Ws
cWOiBetaYNbnlAh4LikbmYnP+qv9WCic1OZm9fnG19QzE2GZSAYH7tWj7tkiSibQ
YD0usUODdjiGgLxcjC2tTko/e/V1wnOTzjvpJV72Bm0NmD13+EdcHVu9TomuSLm+
iSIM4qmGKcQBUy/nJLNqYMEtAhvUlYeCCKhxf9Cksald8pPCfRWwPmky/VHurVcH
VEIapr0T1bCLWrcHrZH0039Y28vLZXqz54LUPeQ4e4629Ov3UAsv9YUO1C/NzD3k
Q26IwlOZy4yXkn2heJPEoZ+dUVCnfnEiYXGbyRNEs5FXSLZk1wmdY3LrHHH6xkXx
ezHndqjzljrH/mx/n4oE4UrzwHYaXc4+2dQv72HfrOW4PZPa1n3IUcpFszVT9Sps
2GSmBB8b5pN4mKl6RFwFFL2oOgoAg5CjK3X1HmwGml1CH2RYSIX5xxcJdDcKpXHq
9Zx0ft++ATu+nfKVy8ARYEqH0XrDVrD4ae8nb6pyRbOP47Lvc5xQ6mUAzm2Qg0PV
dUJR6x/Z2lLBKb6Rja77YctNSSLUzVj5Whonfhe24cTfEUZquXa+3MranaxDFfna
00H/Kvnxywkz3/diKDoRhvtaK9/fNiqMb/FpdLvQ/6eE9eyH/U1+GkyHmvZzZ4ui
ac7oD8moK0g6bqmCRJcR8Vv/941v7fFv9Fi67Qh3Af5ZVxlynYUqaJKNW1FSfJFN
wHTh9rTd8uhjssLrQn8N0drswXQ5Q5RNj/7oUjaTaSHuesL6JOVcd/PGj4MYbSdt
oZGDoGC6w0K1n1mS98sD5XpOvm+9c8rPqf5hCYKqr/cF3UV1Qsc+Qg11v1VeRUgq
W/KG1PEPdaB04YqfLPwxagVJGjtoiEhuF2t7LcRflBj+oJYs7eu9n7xxE/isbWQd
9bL1Abj47DgZuhHOqwpXgNhoyXTI2LPwYkpAH2Fg0MJwx7LfgCq/4jWQTiY/gcMh
iPIi9hhHtY3yKVywqiyjx45q9lhr4S81dan3yow5p/ytRXxtByEO1dImx72c+23e
IKIa/lKqaaLLFlncNHSKxBaWTGd86dq5IRm0LcbwaQ/hwR2kVnmWaBMSM/Nsfv8K
4SODaaERM81gnUMJCxyRhW0fhLaZZqDok1o0ap4VK50XD5kH18hCXj7u6aq+tpTS
qAZTYLHDYw6LvZTcSa0kfZwYtnphfsE3JvVn5BAV3NVpTeM3f8vV6FvBlfGdti3E
Pe1tAp/EwUduGPdVB4mHJS2xIZ/NFCzIbIZWVWPmL7NAlEOHaHzjAMbICsQi8c9n
itmN8b+tQnzGvN2LH7j+SnSfMjgU8H6L8bkVnZqx55VzGbwU3RgILc/sIczEwYiN
hL0pN5hhWLlVE9nqE69NY79NoFGjWNZzTFxn6II4IjAN2VFCbxfBOr120Ivfp1Fs
0+nwnDl0rVyvsJplvQB11A7uQ9dytFgce7LTg4MHVFsSzN290EgZ2N7t+QDMQFM/
FfqaH03L/W+HNFmObeVIesC6+M0P42r9UB0s/0fhZ34DqQksEDAh7Q0Np7z4pdug
5AnQdoLebxvdjfhaUPl5zieXp0o+5g2xt6UJLcMH2lkz/FakyMjeZ4nG+Y2D7v2H
h5U6nnTGhjowlDab1qn/+Di5xyXEXJIHe+NDUgLCeBaZn+TCMwc+6qBEKNUMO11k
cfV8i+O5I6rgLKgCrNo2BRtx79dGp9EAhuSf/4ULaejkSa0TlLOVnibt9Yr13w1Z
o2KgQL2mZVvUj0gCgYbMX7jqf8nxPHiSebdNGWhj3mwyzcimBtMJY0+75Nz8egTa
GQyzQc2D+MfzSytjQ1aiSS0IvCGayTQs/CxhrnynCE58Jh80Js5Vb6QDN+mG/RI6
eIBR3uhje7HZZElDKiH8xVe1m6SylGJkOWXo7NdJVzhQmC+YXHxPLNJDr38mxOq7
UW5xy4WzHkvXXWUKdUsJSn0qOjPULD7b2uicFIdeajkDgBUINebZMB3drF4Z1/0j
BD59t023chFWO0KLn6OvXlY2/QDAqlp8IZvXNqU+n4XeuXUoYnqvzUfUgUycXMPa
U7kl/93qYoVfR6crjDcTWQyNVJhB+Mj9npqtOgT7PzuNmW+xotlZxb5AIsNY3+PM
/As46wjurC4dy3M/bI0bzU1SLJJQnz8TqZzm2tLm7njo28KS4b745HXijWuNJ+BF
6vgbaF3AV2WBog2c8HQJZlt+XRr8XTMiN95toYcS6j5J9wQRtdAPMRNzCwvIb1sI
9aIFhfevrW6oTZR7Avii5c0QDSWpAU0u1gu3RLja+He1HLJYUhv7Jaw77F69DN0I
/VCG6wZag48rubnj6i2na7akYH9Gx1AWl8FAmKEP3os0s67TJ3faO1h/lHoS66UC
kJdOCmwKak8rlVxvzwB7DbnGG4Gd03xF9jJ9anMt0KhwCpBMJmIOIhAkbVIknHEB
tYPj6wI6eZu4/83GWPdui8hDlGLTQEgupzcP/Nqrr8RR2Rqw8SGAHKwNJGI8bE2P
hiJxKvj2D+xEhuqxkRu/ZG7f4rg7mWO4IAxpyMX0ytsm1J8t3JO6LsKfNg6EZ6v7
Mr39x8SZ4p9vMjPXS+1f3JINsGZAXoJiHvCjCoJee3gBy9rfKx4/YrDdoFu0t06z
YKGzHwUVrUdktOB8FDEeeT23G2sPn2QLr6t64TT6hvRgrxzloo4bCUk2epzm4sLN
DTVpRI/RXFa3f8CLVXagOhS7v5od0IrNI/5LJHhT5PT/vj3n4Trn/5pR/HdF/zAI
ovTGWvAcX/20sUpzS0qo+Ia+UevKmU9uwXmbBX/ee2qu/A2n+N96c7woSPHXUWQE
p7Yl6XZwCaE/NMpJGjkFMn4w0K4sd22iAjZALfl0xCUtyhaEcuOmdUCYl89J6PIs
c2axThYmfd+o03DuK1CuTRuStF38cPp9hUQiAxWcbjHPfPwYK3eEkx2xzcmLRg5j
xVHVSCzBir1u470azev2yrygtYbgH6M7m5RhgKjKmzpXLjkVpFjjcByPupcXsGAf
RJRdet/GwkwYLzAsMkT0NFZDO61ZBmtbiZI/BzYQbZ7Zi4/LQNMlUHf4l5hzR/do
rc86+HQpWGRKevM72B7FvwXk+zLF/imJRnlxpkGX4UKsmNa8kY02LcLJlUJbVxL6
HZV4ZZ+VtEiuJ1FXO8JK3oJc1jaoPJSdp2wJn2efAMvXWSMjvTYuXq49qVscHIWe
bmh+iMUmgPwUoFccqzfIpSVK02GUs9m2ErEYvFZehn2I2BkzKjhwMHlcEPaE9+cd
nbaoIWh8pcmfNIerbTZUCUqv9nyVOnFAbSi/6oI8ysfl8vHwAUZVxV0JmNPMtuN6
aucK1hm6joL8ANRRnerAPr+hIYRVjTJzsWIevJ+WdXLO2nM8ozxzhH5ZvhQr72aH
A5jh3YsoOxiZI/km/2qxm3QxNPoCqzfwhqhGf/E2pCSZR+YiA1SquZlhl7eKSYc1
1bTr5/Qxuyg3qEdSNZz25HO4t0o2eFSldd0AOKKHwVNwb9GUTVw8Z973mEfFQP5r
OI7M13XwUoeY3YCqGSfVwwdmp7nETndp01m0YPVLd8JM+V+LS08H7U0sp+MBBdTO
MDjkD+cx7L1naVII5SNpZ6qZWyGH3bt1fijeEdMLdOf2rPe9luBI8DNPtuoXivEN
kJYnuRKmSDNhG6tQ8VtgxNQLBZrWuYV977OCOPVCm23dnZA0TfpSJUihg8WVpJ64
9Kagh6YVIylC7h7gP7LkXsLMBtpTbIPgkA3ILRgCq0dM+njN6dQhxt8fb2kXPlob
EquaRuTdW/uMKm9HesziJc2nSC+XCos0RuaCsdX/WifJUIz5lwgiroaNF4XrGrz5
QVTJHLE7guEmC+rCX8FEjsYhc55ylUVx5IqtEuc3yt8xWIVbDXlzJd/vqGmX2ccc
D3FlnoVghxEZVGQnWpSpgNpI90R4/8OR7lJGS3QRPY/IWMdgg0gjbrCYPuf/i3Ag
P/RsQXO44jKBxTbZ9eGyllJ5/jTYgW8dVcgdm6C2CuEgyCPb0uwijsso/JPDt66n
fVzmP2ydv83kp3W3dx8a1CiZT71BxQcPxvTvcSrJeX2ZCVd2SMAdO0uH7rS/ww8Z
Z/b5bT4TBVZys3VjOxEThTascOzP4rFlDtezvKeoaJ+1RljY50hIbnTKtyjA6hey
5QsMMOx3hyApCxIi9s5sIKS/eEnL56YDXmgvX7UvlJeNQa8ZnglMMFXpPltDlDZE
PEsZmkYMD8wZPA3QFXllKUE/6vkHBvmW15V2kL04kHB/71W706jJLZu9PVFwrm3q
msPfs8uoN/HSyEKIDF85Ig27L95Diek/LcmJCZEBXamixgvtl5IlLSH8OCshtQs9
EIfVSTkBddL6x+mqphh7ntruJmbDB4Ks/4F8b9+kWzyaGNEJkDaoRszEf4FUzrxo
oigJBN5qwP71gbhVprz1Nevl8lJSissXaGGwg0BZ4Rze6Fr3zvpWdQs6NYJB6zqj
1MZbQ0Ies+ahrmk0+QCi/XpGymcoCEpyH7S2r+KAd2OobITcjL91x3mwcCu+lQ6C
b8qSijb9X5unBKuL8eH2ELdOC8+id+pZkZvCUkY+u4Wvd8xXumdwvJBsKmjUrmOo
XwVXYjYfTnLVXFssRyMvP0iZ3Yv5U9nmjpjecvRbS5fsL/3ux5ZFqECGCq2VKoxF
CujimevrkGeI87LwAkOsNodNeQeMW/iknk2nMnCt9O8kvY9BERxd4YQySQPIAFvG
O5JKZOhcm0BvBnbdKgZe7r1lj+0qI2GfDmwAcrBuz5h9GfL+tZmNBXPp8coPUxEJ
1rjMdwLUievCGr+n7i75GrGPBvNBHcMvkVGOz739Q8BCgXKla3sGBk21VBBIIPR5
YXiUstAx326VBrJbcKSQt/KyR2nD0eMmznFfjz2EApha8Yem0DxZLxqn9NvW/XzY
AyLzOnCLQOMhey2yliIinlxqXGGmXbiYqr3QSuJTH50UVtHwax1vk9saImz2mPfT
ygDXaXaFfXdcf5icWoteS/M0KvyyN4WY61LffuSMAydFzoYcvIVXqCCNbRWFDeuz
QLOvW3kYep19oBWu1B52nos04ZATwCrGHhxkbSDDcnGufQgyhrffLh2vq9MLXNAS
fiOH3AgVwEns0NwlTpSFRAT1kWSeRQFYh8/BuELChXbJH8zrfhEJVKeEhsxp2Sj2
fxZlfIfL8/iZrCtwse9165KRrhN+ZsHcDg8mXaIRgcOqp9CT4tW88nKpNxtQqJIN
lFQOwwBiKJ5Y/lZyirLS2FmXk95g4DmFNWz6p4ZHjXrohq0bmuiSAxppSZHXyCQc
HuxUOorqOsZ1u6H5jQZ00SoORjR66NXfQLIFkX2KbuAIGhGkJ9HVfN/daGrlPm2C
hHOIICwF/ylBDU0CJArSIdbVlRYRotTUmiHNATY/OyxwYksRgKjqROcjA+w2r9jD
pJ/AjNgknCTep3766JWDB/xmcfzQtbknhcKjeJdnUIbiQwv7KwwCe8gwN0Bu5RSi
/Cc2fd/Jrgsqqn6E99Hf+BPG3WmThkerBS/W5PuE2hzGCTP+ijTX+oT0br2aNuge
LnCbj7kd6PXEv4MtH9vk9MjWNd8qqI62zprDMbeB69wFooIiIxbTxaNG4JBLUFUN
NqfRuN0hQ6WXWDPXNWP9vyC2wdIRoNm0iJjItZJ96Sk3PJgIWu5J+evUO1Xh0uVn
A7SjqQ8kKXrreegUIQteIFpjXrWGGtA3jh4YO15gZAn4P4DdglCB6+07b8QS8Hh5
N79vquIiqUzAzPwECq1P2wrHC5TBs7YrPGpKegsdLG8JbOqOX41oA0Y0d+sxv6CK
S/iedhWlb2+Tuwgc8vmGPj011GpVqbGpT5V6I/qgm/X1kWe1Kdwx+wZ++/ijzDmL
4+Bu0aEzATBRoynF1GW15DX7etwBvfUSJmAO+tr4T7wxvipBjf7Z1Kd3LHZnB/ss
2UB4OQ/Q4K9JUU7zNJGdHy9ZlonO746V49Vg3VSy/J2YKlTOiH0QptQ1KUrPxOni
y908ssNlm3rb5KoL2gvLdSjAyhsI8B7YHD0hW6ppj4aFuFVDdW/O8IPllQ+s+BKh
VjMR61jmDBSmJLlz9zIiJ7Chyt5qCdnc/8ELa0eIe+62SR3i0okEoickuGW2Be48
XBbD4cFjQOdbeZVZqHuYSzsfD0eFHaUDpr9XTO0JB5BZVx41SOY2SdcaVoHRvVFF
HPOKw5d8qyYugqkzrZB+bAQlhjSpRPHUDwz5u/PV3dZccMQwgY2UdmZHuaXLsnt2
lbR1n2maWfnIL2CvOXi69Pse7kP7nYiPQsiA58KmkzgXyrV6SUboBXeyAdJp6Bv+
EpVVmlNrzMH45/qwlulzKzqipENCeekOBTAFQKswLWhb9UTWI4uor24oQgR03YKm
gLaDaTamYZoJeunY+smrC4RHKXbCCFtUy4O31bXYm7Ct/zRMDxS+yteRcAYNgCj4
Vd9VJwsd4CXmHleAQb3j7l2WGQctp2BnJdlsRO4a4Oh6KxOGF23PE9iFOtMZNaIj
siJIIeSOPxOurRQ3V5YwU04lTfD9WlKHUz6YTnInf5w4bbJO9nKpjAbECsHSzlOS
7IbwEbq+JJJUJ/5JDJlsrceP28Zv5lXD8so2tvYVJvn4RPgLPrxZdXypodorY9pn
fJ9vIABPEUD4s+Vlbe+lOhVE0mBLea5uuQScJym5MKosv+F1DLmkrQz7NtESinNh
JRothYf/HllJTg6TXPC7Y4BdxxRFsNzVfvEkRLUDjG6sZdorfuFrHUtLEEvw3a+Y
e6k0Tte6Ml+z1DDATZnlJeXGqb8WzdSUMo/Z8+ks/IVFAlQLWcf5JAoeXEZv5k/x
vExdzsns+jyGsRu3b69HYl8xLZZ8i0wPodx8d0DiLyid3uOgJ1p/QZzgpbDj7y1z
MxpYjDESRkMuWrHoehjJe0hrQFgqEkaHDqBdlB19W0xwaj8ceS8W2JAp38PvSkf2
QDR2Qy4DBUMbOyCg3HqqACvvsYyDW5ihrewNgov4qt9l+ff/O09dGBoMz6+k/7y4
DLIu7vuB/+MA74R/VGho8CPBCDm5+Xl884d5gjrc5WujqPYECpYD7wB5FxS6r5M1
vYFYCrsL03rIDJVaO9na8AMzFI0lnlgrannqE6sBF2KAyOEonM8NpBld3Agqkt2D
2gi25P9Xk4QFip7Du8HnbfRvlCSDzzrVbVGf5e88Mcudm9Z2twZHJB9GZwrY0559
6N7mx73Xqtc3mQlevGCB7/kwcTKMFWgo8/ZQtBtjjK9EK+QyKjKaLCP3pqOptVHI
nDctoDUhdiB1Rdt/hevP38GnLeCkFBjH9OfSUcJ+clwx300x3S6otUZHb+wtXpVo
4imkVy9noUrVDrRbGZMePbOo+EUcU30HBMnBHSoyifZQbj1PZpEohkfCQUaH00Ih
28xx46lz30gZHAt+PkM7aaUlrd6TXwWUMwLlTKc9zz9NA7bk9zG+tPny5TaXBRP0
6NCCNwPSXSvXW9iMq/Q0qZRFIU3zfMBOY0O6o0zle2jWCPpRLfuBg3c8lLtlnOYl
LlC1BaVq9RO3JZ4l7Q/g7zyYAA8x1f47M52ruN9QLX+Htm0PeL/0PQO7U1ZB01Nw
JlAlpzX+N8Tk8lhMGntbqEJb0AOA5kqRYmi+F7rru8xSR66PJEjbTBNpRTS1Jr4/
XDUp4eRj+0W0AdYffo1PwcGrilht5sI2AXdYFDpoKH7NIjL1cwfgyTxiyk2fqsJu
t5W80p0J+loM7EUsRZpQtEu7AXGKlWCmQ6WIBKwyyMGnYsEicKHOhYZHsvtQH20f
VfgWDmoTDO8+s9Uj5x+pm8e6/45ZPNG1iCKdeolPucynV64cbiCfwkqAxuqMhVnI
erM5kylLt+XAKjDKXfkHlb6HGteHc7rwhvJULDaoI+/3ATI9uEMSO57HYso/9Cha
LedsNwG/VhsCadxV78VKHfOWUXPWeMmFZz5AxOKAWK06hQUHlSGTtNScmcKWCw/n
PG9aPkQTGDu3l7ysh/3zFBpBIr9moo4q8hdcL9hJ+4INT2Eojyw3hkHIEV4Dn0w5
1mLGfCwqaync6aEgf92vLWjL4iwsiBaPzuAaQ+9T2xz8bUaHWqLns9FAsi0Hzf9l
wPCkTrr4Bp6ESV7N1Yr39iCQMHzndGxjfrhs/Z6YlCPhwJPIv8b99n3xdJDRZj4N
AC6AnPPJdzK1GssTOSUztrbaFq+KobGiCMUDKXQVw+hbmRdc6cn87uiaDwHzkVdV
bIwH6iFnl4okv9THhUbClXdz7ELwM0eBKJzWOacu4p4E5opSp8YyK0YTCTwCMmdp
EX9DpB5rvLv4IzMYiREiqq5qnNebK7QqszVdE5fZhJf9TFhS8mKVM3ZcVvmz9w5Q
8UCWYprKyWMtZBKZ7xTMxCzgM4SGvd3/EUrjTP2RirJkDJh7w5ACBL4YMBC057wu
GQpMRDNAlW/YayL501kYiZtqgczmwDUOhLGzt4OpkcV8ooaAL2inla3pn++N22Iw
k5qFFxfLLPaNOvyXhFoNetemUCAZf4lS5vyKkIIbgZLjaOYyIC9PYMGZLdnG9tcb
NIki3RKgjBCvgcyS8pychSTz1Z0JRe+87RG0IWQzUJJ9PBhnKUAXDpRhXFsrMjCD
Rupa/554dkGXBeCmgdz/M9S+DfaJklilH0+G49IyCU0YrpSy9O3stwKth27Gw0FY
Qzdchpy/0CJQg7OHwVMdyH4Bj9LP1RXKFooOsKNyITFRrH7/QDkYL/qrA3moJpHP
W1uXcGXW1w10Bs01d3oU6hJWWDAan5v0wjDnopO5rKpZBXgdnLPW1+5GMpBcWch+
00sbw1L81kbf0mK6i5XEwXcMa5HloKWEmgkFoAuRmGrmIuexP1zNQEurYpQYvNGj
+fovXR9J3swFnJXZms1xNfhQDpoOaq5lhioOpJevzAtlmMxsIrMfAOiLelu+kSFX
NuUyejYKMKf9+CADtobov9maq/gjicPE+yPXgOVebhWmquiQXn4lZbwJ9sZ9w4Zd
afGVWKxZvBDsC8wrWQ82DNH9/sergglEQYJzMYuSGxyTVmD31w0iQ+x4pOIOpXgG
F1qBu7hYfXepzvdpwi519L1q4z0+LXJ2nzgrHPzgesBtrRO/TPjx2YAmO3zOe88G
b0hLaKnK4QoL62sKfqGENlg+FbAFE5+nd7dzSHjZGCSiEJbNWsGLwCMrYD3C7TbO
HTfkcl7DXSefN2rr3WV5BPO0ftSVKWQzjCxZsRiImK2cOP6zx0LrbjOcYVt2n5dg
c/wI2JMDn/dbVsbOIoOsJQtx+/lV/gzPo0b3KV8tEAJco9vg6xQNI4MOwlg8tE0h
RonOHIJrf2Bm/gONc8Qb8abm2FShIsYy8/7rNkUE4inMGOVETTPNcHDzKo49k4Ae
QkWjlii4TrAd87baC7LO08t/6YVEGX3Ka3mzs82Hh74YJc2iXkO5JZAZu34GpGFB
72CrBzNs1HZlI4O6ecSoD7FlP75KyatJKJPTOGpdPD8YpifpmVcTE66aGxUozn+f
TMxP12fcji6vQkBUtd+9Q9uWHTkDg/EfENnSKZIrmTJGpkduhjgKqs597V3Svn8g
fcQ7xP2JMQtJg3lSSyHF+TH/CcaxEtZt5+criD6EqOimA7v6oZ8z/WcXWA+ZTFVw
Q1Z7NIW4qDHgK0oSTG2FuI2lNHZcc5ZgCZTUoHmphS4DjhnIaQG7lJH7AGg5yORf
jjaGAYry+CLtrr/XfiCJn7sSMO9tTnDMrxzu2nogYWWXF202h9Rv4hOwbIMmMBkx
LCQaWsRDF1iJpuJPVK8SHpzoaTb8sCVDe8ItkKQArHvwlcudnaAqEHpaVHBaCdVI
n/l8zOo5mHPRwbgosOs++0mdMPw+hbtNdjBBNk4dwDzkrtvTRlXyzxpqyz/RxwT/
ylnFMS7/rhsR7Sfoc8Sj9Gl2daYKN5z59BVa6JypWtv5zRJVqAfKV70WdtBGSWej
kkoQfF3NlbMdW8fZvTtL7yC7mBW/nFspUK/4hqJIf5MbXj9XYJRyB6+GLT2i/Nst
MzbzDiQQ4VwaMgnQstC+sOo009seSYzEsuf2rtnkY6E2mfUWbJlRefE/gptQou08
tDUbNkFtlqB4CO784mA/amBvqdJoFsdCP1wyxy4JCimK1lKx99ydeYqECZv31/0J
tyi824AjCBn+SdUefr3QXpz/rGVjORcIbYzILCk0Rtz8dL08eyytWZW5Cf/Y97t6
aHXiasu5hpHLjMIEPK01OlJbCL6P02qVWiwXfFekZecXHPAVoaIPCeGB7yGvozQP
EQ/dTlb7QZgOFZJkXSxcFfApa80/GR8g7Q1HdBrs1a8peUodPp3K+QFlUrScKJtc
b/tFCMzar6kIVV+it7+Yaq+XbSEb/QXx8WR1Rz1ouCiA1d3+GSBOy0AbEc1HFMnY
o6zW4zi/KSHU4pD6cNjpMJ7WAyIWpAn0+xAc2TjxO4uBlDYTC8p0HyVq825tCRow
YVXUs+sJSnoumtqgfqj1oRycg0CycDYc8qV4WD31HVV/G1EUSZ8G8di4ihYz0X6g
A1jwAklo3rOhksONYQXV5m9WrtzASZ176DaMLrPN4UY6e5Vxyg8YeMN3z9olCgID
Y8NW8YvzEYKW1R6/RNgLDDBKAqgyW4HbAi2Tniy2/MZDwUTF06HihpVQyTq82TNv
dqjRwfQV7PAsKA79CVkDj4YtrAsgIYd71HRRSgax7iwMH3CGJS/eluTzffEJMAtt
OU4n5hzMrZ9Bq6y0YP2z4OU82adf6V30jC3aJC0AnfVcIMpKlS7qxRwvPxIdZdLD
dZz8S2jSHZWzhCNG2ChatgIEjC1MzGtFiSGx9G+QKkftqTGWzBViulkPQ94llfh/
/67a0u17S/FBkkus9rI3C67e4pfxu77bc+GhZ2uCMGpwxJqjLINHOjzIdLB5u2CZ
vhp9rPy5ZsgQnz23Rx0Yoi91/TqdVZwQPryEW2LKlFcOHUZPlZkWZIzYXM72I1Du
stl5jdV02Fku5dYJLEgM9LIyVxYnr022DowVGA4vTgivbVOmksa6FH+YkHmslapp
4YGLnY59AnII6OMy4QfAmAWKFbguAesCLYAg5zJwRZBP3UuDjWncAb1cT/vl7dMN
5rlLAzz+t6FSSKcbd9WOZrjcsxaLfnFMhMlacIaKCKf9wyHJ1jDrGlgE7ir/f7sR
+RRTk0O8gjBiuZvrbAyF2y2SAXPnldQCo4fq2sG96AeVg6XSojFoVl6uB0wk+BFG
dvZAJWiWLEsgQ8pesclkrFU/HkGP5MmA4gsNAxJ3szpP1D3kVmxEPoaBxcg0J57d
s82Cjd02AbPa4kvpLGukYLd2kMYNelDw3zqOxuQspDNgpKc1xXfR2BaIUsffg/cy
qJkBVep0IMwZpgU1iRcRw90Tc1zglyj/WjLGRYQnaW+Luy4jg9fQSZuGZhcX0rco
sOWAZs/mV/DiCOtSVjo1dR5k6tTd23Nt+hgVVgm7hlZMfXiFJT8qYlYECsHAkZh+
2f+d1Hj3XNaNdKMEUZOimhktGpN7CmdNthRddnFov4df7rjFH/VY+gaMgcA5mWsK
xY0jzdj0sHxKQUZ+49+qA/oxpRqJyD+rSet91NJKbzazuJ9AhOYZ1TPNtvkKd+TE
JRjECNYDdOxHTH4YhxSG+g+exGIOaQG4EifzuXYLdj5DJbwQe7CBwSl3/mrg/juI
NL+LHBtZ2YJZ9U31z2rhuBjXETO9TOHelaIjjLN5rFT+eecZKErve/8hzfF//ka+
VVzELE0piQ6oRPs4B46gQFvcvOq6glYxkyNKKgRgMElZ1jpCBLp+/RvfWIjxFBcJ
hyUuJ1lq1AV22dKGeK0000IoYlt2nHlqo2hIkHRa7rgQp7KzFR+GCnaIZRPnAqwV
IrL4QGNq9RxkF7zLuDI4Vigw9GFVkP1xL44/fmEal5tW8O9KcWICK/0o0Ih1fCQ0
/K+FzbawYdp0PAdmj1RDGcT77NhpB6Sq+wEz177kik8sEG2nMK63eXGD5KEJVoya
hNe5U4yRc/6y2RCgZkuMoJXUswmHbnTzDO/JuTQ2KEZE8xsb7q/qPzb40wOIubHs
aO18bYicPVv1HdnwYbJwdipkTuqha8hT6qVoCeQr70FbpAvcbkDrSAcMQEUEvNIp
h/a6V9VDxCWz8hnGnw0IpjwTIrvEMO9DT/3TfHJbjK4Yigtt0UMOfnYTgBrqp/LN
s8GLhqL650x2zWsNmoEFXCx32jp5FbmHrxm06JzwVCjKVvWuwhjXcm3aYlxVUExZ
XXrubVvs3oYdmdANzqTD3a77e+UYOTmufegFqYZLfTA+yUoV5dPA4NSHud1n89DK
nrQfqKa7ZX3VCzJEcsGuzGJfZjEVPyt1uWaeDC5o29Yh1Jsx3qGiF/N0YWAIMDas
B/5PBFm550Prb1sZjsYYqnu+5L3UUoUKF8E6+72zGHxmA9Doa+xaPSA42+GVybCg
16ituHPorw4OriiV5d0K9guV/fFegT5axEuhRZwpr0RJl8raALYvfiI3ZYDbtbtR
+u1i2YKftN2seztsvC/Ane52om5CHA0y061O+7zUtJboweOkeAP8c0xr729yhW64
KEqSrGD9ucN1DtwmJgMnmIkVS2VjULOAGggITUScg9vIeUK4iRe9V0fmC59kbWgj
Zgrdzl+U2GKwtIgZuJBoP34fLnLnjjRZeN+ChyjQ5zjUrl+6RrQqoM5DxD8tDTiv
gKjcRIsNz4nmAM0ZizLtXpZS4WFIdppmuWDV77FqFZAhvpHMKd0Ru3ZHAKqOiX4l
kPxiBKxVfhaYlfYZvhmz/bkEsFsPcYWii7BIeVQbRpLU+JLkXbEKUoCdFDewfcYT
SRHovL301Disi9/jI5th3PkkSadJjK+i/AZiKK/rBntAGWyMyPPxWlIlobIkMRYO
UVvhwz+X4Z309FL8Zx4TBYvDRcb648XGmJjeAtMkR28f//y9cAtlI8QDshJKO0dE
5w6YYNbdMsg9f/BEUz+exIKXqA5susxdFIudC8ug6mk1jn9W4xmJhJot6hZr+PPZ
eVzFRzeeLBkNZX7yfsI36+C4rDpASEC9qujsmKYjCn/Qjaxk9YWzqTeVVZJt+BSd
6PpdhZeHYDKAl8YvdKjVirkABUppKs/PIdUteZMcBEPx3M7NTjbiYc1hOuocLb+O
9tHB4UEU/Tjk1mqPI17pPKSxRzMni8ucZ+SEF1AiuZ41PytaN71nq4rE5Y6NpHMB
XowlEtdXeztGOnpgmYLyJJBzlVvKZ2lznQHYBhFXXacdsAUfG2ZulbUtreQfx0Kb
nfXbqZpfgDnXdAUxgc4cf79fWaO+qDgKRWgzqV1iur/gRfUIzJyoI8ijdYZkRe6B
Mf18m0MTpd1fFGgny8/dRGRUdAzgwkgQj8gkX8Sd+tuyR2RwmifwcFkK5G/2jSxF
qQ2Ik99WXK7tsC/ylFnZM++18OFOm7Z3Wb4fNRowjA4tgKADGFjsKn1H5ww74lfz
GU+0YD/lhS2hwKsGfQ77ZyW7p3h2sHw93V0THx3nAOlRjXgnN8ybi5Te9RsH4vEi
6ggm4jeMtOUCvHwtFLYvRZ+XD3hRKvRdUxm/22PeozgcYAzWNh5N8zfcUlYRdgpx
NL5lxXl1DWHkvxpl9xiL9r78XROCRogGeK8+ygVM+TNpMWmEH75+ajtDQN/x4KdM
Xpbau7qWFlyg6FccfPZQRx4ITq4Oax+GjOKdmSqEmIMdxpXl6Gm9mFxxTHzk7NsX
jCPleIDV2Yy0OUqHc5bH6E+utILg5w/zdwDW8IniVRZHAYVjal1ZTXabCVTvzb9D
iUosJF4d/LhEsnr3xd+V9b4B1qfyb/ZYR84fd6FTllT5KNgWh2UhlM7WhgioeJzv
uA1rSzY0a/DE5wy/scib8voYdOK9kxifgC+0PfmodX2GbwPo/7+VQiI6dBg1Aj7a
SWrHsBJ8pU9Uu826g6IkZ4zEtgHv19bgj3UfnOpQm9LoctbVO2inx2GRZ3mSWdjf
35dP/7YRBJTsazFunE+fe3zC1y6icYouBGW6cmSCuWySgymenuNppmXv07OSEs/j
HN8zHVKfzyP+IOop7KMTCGgjMB8KCNd4umhneEwF01dsrkhR1Hnb80Z4Pskt+hiF
pe86pdcuoN/R5TXe/n6kbVQBC2NiiJLxXcpaHW4yCD7rLuHyvIrJnWIWc6FrnQST
tk6yJQm9PgETZn+uKG+7i5mUHMYplPtRwLbMQ2xNbiZfYOUm18YtLiC7ZCIpalky
+g99yVKdSWAsSsmAtwBzfyoA9fTSCoFPYFMCs4nhYbOFr3CAq4qREj03OAcHp+E9
hj7n8bNgoveuokafkg0a1sYy4xWwcv66Yq0uyGQhBjEeF3Iv7cq1NeYdG1M3C8eY
YRxS+xrtH5ugIwU2lvYpLCdYuh33WeU9aPs5Kcn6+fJV/RamFDzIvhDOZg79LTtn
zOjfOcmm2uTExUaGAr68e0o3xbwKxswpnO8hrbrjFIPS36i+14R6bK0tK/1K/Xx5
bgQj2vaNcs86cLfPQ/enXZpkYh309bfTC0N/3SDlgY6SPgPGuiwSVAcfoVThARq4
J2q8CKjr8eJOGdTxn7UeeJ4XwDgc7wVX9VMq2wfmQ2GEG/eFMldPd3qWtgjE2XAZ
lW5n12tbhwpXURx0eRYnJuht8Ls4Y0yfF+v9fgK7KsNMuj1j+7XLL1iPQVm4R3FT
PFJK4edd33Do8oB8TeuEdr5VqQtqC2JVRfcoNZ+a5/FbahVCNrjj4NEnM9bVq0Ii
Aq8DlHZz/IignvMe3Tb66Op6HxUimQlOGE8tM0XFS8afKKEdvegSlLRBWoypD545
SgwsSwCBrLvFSlT4+rfB8XR/oHQYJR5/xL882Mxffy6W5FC5q7sV0sQnuaPjMqtU
J9+SUug7jeHYblJ6VGdkLbAn9diqmjDVW2vDX2VqhwNw74iycgtgbYYtDzZDZuT9
A6MZUI6WQWg2PzaunT9NcLLZfggVMNdiuICqoLLLoi2WfmDq83QGa7nufC4i+hZH
UQ1qj3OdI1c2ihoCSy+/YHFwqHa8NUYV+0cWafvUVaewkO0/cF0bYLiYyZWfOfrV
jFurNsRGbU5xdqBiFNp5zcJz955YniRh3aYwEtgVvWgQpo1ejqe4uLQbPfEHedu+
WV2VLfHCKJK6uRabU4WIGhBEsx/LHJZ9usoFtpT7PZwZKHycUZ0o/2lTig2egFUc
SFQ3XTQleF3fSBQ6a5dgRrR8MePa2jYuXSxXcWPfvyFWlv/bBcNwhLJ45rP3cu6g
XpQlycx3XwNB1hK7oC3uSODLhWFq6shvU1nBKUKniRDpBNAl9584ih1DIIDAcaOQ
DxXYvfEgoB+NoJ8K2Vc9qh1VGh8IRMgIGiCiVw/PLW6zUiaOUWDnbKQwiPIRUpN7
R5Xmm5gejJlpXD5KYrq5yH1ek5fRTPOCalEE917Uug3dXBMM0z/H/z+sweqITF3k
ftTit5QWAxEZsSfZgqHR3cGU4gsL5ZEdD3kNPUIGAgEBkDdSlsn1atIbz1Ukhpss
wRbg3q1ehBhvmdtq+4ujQlynaCKiF4o6fM/6YlndDO39gU9D0KFoziKFkjfesNR2
c+X5/m5YPCLuZc+hGRJiWWzHKMVj+BLz0YwHvy8FiKMcznQpMVh+jrqHzSuy6m7I
XYXGo7Xc+4qf2Exnvc+DAeTbsjbAt0SSAvX+I7aTue4WjwWdSA/ru1mKIrhOvMbK
Lm1K08cu//ydPKVxYhNbNRmqKPZjYXNfHc7bVuMVj48bjxubFhxtQwXSMVgyYL9q
oawWrNib66qf1cEbXUTx76+Pr74l2xVVmgBlm9F+ZkbbGMxGPHEqDnmM952FCzTg
r7OiRZgkYcIRn6CiOjfavpIbnl8Q9tAI54UYF3cnWCbFaBpJDdCkRQJlyGhiZ93Z
Ijx8QkJnF1rJvdj/umeXYbxNqCPnjHx3K83HzqB9yK0xnhAh8YV285tVJ4qvbHBY
SOAYKpAu81fSo3xR+PyLXtIEAYCijjgKs0K+GHNPIunafqmhL19ghYsFtyPgH/Kk
/6enlrROaJuywGmfm2JgygHNsgNBPka9eTpriEdXWZvEMHLgAGAN3LsbhIg7kYRa
cBO8oXjfqcgUcne5eSirmbXTRm6BNfhsYEAR98n0JnBRcGcygykks+a+tg6HNIyH
WFn+aEOj5W1M+mAp9EVxnQLcxQm/RbK1Bzinio/KSjLeMxSPjXq4aZtgXPDX0Ik8
VQJKUONsSguOeMJsA8PJ15UX5FvjNX6JYaokE05nYkEPhUE7V/NrB0rZoatTXGYP
sAru5ymaJ1LRkR9QowEO9cJ0xUoSGcT+mLz3OkifIBQdmrd4LB+l0ftI1NSFcEN+
W0eRszUs5UWZcBC/iM5CdUkpDPpVUtt2JdsM9WMx7Xlg3cWNe4eGCpI1130g5RSY
IQpFj17jTZSBRfG1kJi7JJOmIE8n49A3P0v8AlHr+out4b4TM9DLOV5uHu37n2R4
/UIJcKTsWJUUu4qlVQrOuSJ7Ki5qwdJ7JbUl55Hd7si+fDM/UuEyjd3EtOy5Zb/B
Usn20or8ilHJthaGATxJ3ulM/HqP77yL79n0NXpH8LGCkYePiv9akkCBpYZYuHoJ
DqSQ1A+L7OUD2Sd9z4HB7ZdfD4lcXhpyAZBOL58WfP4O3WwZ4qU8rQu7Rw+6K7dK
3gXrAgVNnSJN0Df/fi+ChAouJQ07y5nyLYjFIrcuR+nUI57HoPie8smNgIUgMY+C
AX8VQGXjMG0+HXs6RxtYUHxQjbbjjmObzi72KM3lor/CyurNO9+EbGPOw4HfENh1
TQSDfUb6H2uFQT7n9wrorGcSjlniQCsY+f+bvmYVDb0ITYKTG558xygrmDwL/55i
+Odxo1GhyjORMzKnfCQe2Zi1dbt/w7bvsxBZmW8IWkjEFX+u+1kaHhOP7op5CdaX
6SKAMQFVvlMMlpUoX7R694OSAJKcPu3HeJqOB1Yv40LNO7NAn9OAdcs7JhB72Rbc
gzg5LHlg8EvLitg3LDVVUgHTemgnSyreCX6nSK6bONKjZ7zKTbTMf5kLwTVtOkDf
rCiYgU09BMwPPwArccp1alSqg/Njcace7Al74Ml+HgQ3en6NLfm9obwkV70AoPg8
PRLMpvudi6+BeuvXpBf1tjMcffuTg3Z2Mkaq9Np2rlymYbb5lA47AXWs3tZ0Uxxd
mtpF5NJShOY+GmD3urvgVFiSbjY5AwSiDnCqfAp7V0RJ/B0Cu59CJMj/+fds2Gdr
fSbRPO6mg9wPBXL8PfoDjzuQ4tx0mroNU1e+MJFB1FMeu0sdI9pMIcdJoVI/eSp/
c6Yw3eqxi1Gx4VHoFXrr/t+8e8zmQl9VvnVxNFGUoB3wibBvsYPSfLCGNGmrJU+q
GgyyNhnNm4xrdf1PN0p/LewSf0+9VbA6f2WFRlbO5XPhegCD/grr5NtJY/86jCnu
AcKXjycyT7vpxeA7Rsc7RS2szQT50Qx2BD2s3rfi2DxBZ2hwAtAqGAXaYsdX/Yeq
SUh+LOQGyd6JLDUJZW3tMrZQptiY2u/8n3SriEipF6rtC8S8NaYn1P3UAKtUWH0n
B2mRXpHLLPgGUOIdP4lc+GMyVn7g/9XCTvSZhhWTk1lQABQ84JWoh+Z25Y0WGE27
KNix/WR6G7EKbIp8jlTCtGToIc4pUeYWVuk/eCE0TaAG9IdY7VRyF8esaDICwy0z
cNLdQhFtL917qvA/3fyOe7sqWbtCw4O3/fujupu52NTmQdb69TDSXCBwyJd1a7a7
LoFwQqZEe2MNgawtT9dEcmKrtFgGRoYaGeKj8z0ehtb4HRrfrRoaizcZdiETs2Ye
GGn6exTa5L3abs/Pcm7Yb3z20g2JxSN2wmsn2dc34HcLJTwipHHn46qCAOrmPwPU
uL76o+Wc1trjciKAN4FahcWtUYxvZOfQQ7pIFGnSTsvnMqTUmzShoRw6g4Jy5cLo
smCIlzY580UsI3ygpCY3rx8jKtafccSruM6x0IYeAUaBCplBuWb+y6ZXepRgb2nI
3scD/BDyPjjylxrYVBBDQvvImUyApjuNPspcm+W/td34d9g5WpVjRLF1ESSv5HdN
mWyk8g48DKW3IibY9uNvHOGjYSHx4IDSPo20eXBgSPzDbPbPbCH6O1nd0YDyuuTn
3EuFuO2mKjD5UkQYYxT6ZsL6cbNYmvxa+VzkfpzxFjmCqCk3AAM+H+c/1lgWlxQI
J9wJWXzlF2fyE+8XnhUpKSoSg8y6JKvpOuKyP+LAQRBB/xYUMzqhriG/OUtS07Im
JKsKhn/uk2lHh+VyJ4Vr2uBol+9NxnqjLUT0FiGZ379zjx4J6kFTk2IUIz6+sW+Z
3IwkHmicuwLaoClUjiUMqnBXdPJZ7uUR9YFbDFCWwzKyQ55vRT6ZaRwSqirV9yC7
+9tft79du+xR+ebCY6Hpgj/Q6zluT+sI1+aO7xtCM9rm59LwS8gb5B6IOF1ldCA9
iGs5oTVKMUbPxnPmx0/MhlxGJ1Wzmc+zgAZpE0Zkw8vT+pYE9eF2XAbJ4b5DX6wA
SBMzvsy6gyok2EHdk203PPX4Fv0bDSLHKA+uBiMJYnIMCX34m95+3YOgpxk75b9p
dAdbq5nk6ebvCFepDE3jqpSS5vFEdBUyseNHXAlMPnOYyjpumMNbI2l1I2z5ozsB
0casqX+N5KeJ7rck30MZVBRboqTBHXX0SeURYGG2fl5VkiTVafjtSmcDhh0rvXp6
uXw/SAMtEStOjKBnK5hyEkc3a7Wbv5GndMdWSTSujMrr7Lqrl02XyBpBqDMuIXF2
y3w/2VXJJGY3m8NDO1PndDp5wMlv/uVlRrVEtphKqdZ6U0gGmAI/2zv1tXS6oVp4
iRrcYsQeQM2G6qOoRsBfqevVImzme4BLzu1+UdqtVnmVh8L+WweSIakCBRYPGks9
nOmSCgmRXZf+rp5MtDpXpeYHNY7ZztqRva93QZQTENbHFxwfixzKiUZafcrUl7fX
dzlVcgrTKUGfh1C1fVnOWwsYqcAfANjVJX4rKOqO3WHAvTz9dLC3CM8SVn/mxGbN
DTZfsSccCak9KWt5DhgdfdDnbs58I6cucor7QKrZwtdZ65H2aAtBkAkFRWHEy0wS
NI2uPHItT87m+M+nMRdPqDcWqq48URmFYS/De6Xn6ahge0J2NAy6Btkc6OdPz/94
ZO7cKpPKaB0K0j1De0YcjErreMwsTFGq/C3vvzzZSwqAJDmDKvdGMsMs7JS+D6gX
60B/QB41D52lED+/fx3/da+KOq/y/B7nEmqedUrrq8DgUnq5Y6EusvXAKwgLfrj+
g9siuwDVKuiQn5o5xIrcUDeeYnk46OkTG8s7XhVDmyLQ10cmkSoTmCbL1+bIpFps
KJCF5yy2ePnLWfzkSdQ+KRGQegpwhe69RWhItoHJTHqO3E2lwfUYB2cbfNQPrNuS
kOz0mjZ2S+vpomszUupJkHeRpxk65ADd2HLmHAtu5D7VHPmWtYnWUV2gDJ4viyxd
hnX4Xxqsch37U8b3xF0c+/5XKn0WbV5weNW4cW5mbP/EfpgD50Go1jXw2rM8drSd
XAU+FdDYkwKFx8vK4kqrCQalWsiCGnXgohDBtHuh8j/gXe/5c/2ePzDW+boofcV8
4rrofHCSZ2CFHKO/vE0MPOhKFOX2Pu7E7wrqDPLy8eksF5xuRI1VdkQqbdK1/SM+
/y74PUnB1CZGL0URIPF28GCUh4+jUx/ps4MCrlukwxRWsaheJlqvAwiOu29UhS2x
KgZxJwrmcmhcLMwnUY3nmM/UsBPRXGmGVI77qm7HY7N03kDVLpJW4I9D92Zh9+Rc
D+lh1jPkQEp97HI2jM6of+Zfn22mKWvM2Or0ufD0dz7k9vuQljRBPaRA48ptDOFU
N9iQWMZEbVp0WL8Y2cBXmJefaHRhj6ieM1LvoenkKaoI65+bJbmk4oxDq1hZRg+0
MdfwHwpzwGfJDGCjf1ieTLKr8bGkdL99hNx/x9Ex3mjLV3O/LTvJ0kbJmM2+9Aah
AS4EK+02tfRILh1ErGh+/UOq+EYvGesRpa/vx4gJzBpy/cx8JYWtHmFDuNGgqqFJ
li1upsvPkPZAHb1pTsAAO3LLHP/l2Xz4/oXYKjxrQe/l6qQ0fw8Bj7aw5k3HvllU
uC/x2Cq8gNxRvixXS5K5/r9Yo2OMBcJB12jYy7bxisJ3E0VVjU+jbh7uFmIE3+Fs
BKbk/RBjTA+jRHbeGkI3iXaHWNYMR73mrElruNJ7hsEuvj0GO9/sj23KBjW5xXvY
KsHs0gbVj/JxgFvBhOSzpyrDpFfhqls9jnvFl6fvOld7C1wqp8nbqig+JP1YCfG6
/EQqLAsSHNouzFH7wrAoOjCgQeD6h1nqzlvnFfR9B354/u3UIhz2XLJTfr8F80di
SSZY2a4R5uEerH2q+3QfFFoxfbSJ5NiiuaTQjNfJGOvlevLQ6DELOgdbWi+01qwm
jxkqOj2Qw0OZPLGyez8hnAPbblr4dIiMGF9qVdMokiSv/UX/m3nPiH/ChESp5Rd9
U+b4LKLBgtirydFFI6CPGFynJKxr/tD3NDFPw++LtTKscV5kRlZqLiYcftEhawcO
kXDTmwx8FmJfx7tLFmaJd8lB4IJCTUaSltBUPlC9HLcy3N8eQrwo68xvkSYNLKed
2QQXGh6W2VOnbCh8DVsCuUXaXYs8IBNlsV/NqiZQzChCap/3uRj6YWqGEqXenKf4
gzOxS+CtOV3IfLd/wSZ8ZPcKTPHBKeTYGx4HtCGd9t/eADgSTG/xUDYdFhw+8Bgl
c1P7y3jywejn0SCXdaZbbyYqdF9p7hxhiu3rAeMDbAXLUtMUnaQKHvQ2CAst/VAJ
4zqivr4eO9KpvxkEfJtuqYGuiwYzfJRoyiCwpM0qr7mgQXfESrAnnP7WPdFC2pdS
6wdUpTWucwQpXTsXUy/6D+bcRcVSezx36wOktu34ZsPD+cKwrAHSXjQV/Bw7/Wn9
4Cg8IOaNwssg6/HieC+FHRCNgYzJeBNMd9t2gk0bmRvuMg56AhdQ4NS6ONBF3TK+
RKy5Va8HVXq9yAJ3m16P4ePkoRvRopkNZ8/+JENz7vVlJ0BQmXnH9EtKppoNdshW
DC6GE7P8rqHCrEsTVMgAWs7VfBNLj16lPfNngNBYLt7ASziWAkAeVu7H2Kuy+nIv
ugA5RlAdPTL+CtrFctLZBHVBACQClWCscPdsQ0AdqGU80WQkDQlJ7mS3No5jfnvX
JQp/gynkNDvD/txYo6DM/A+nCv2svley4Rb9+aCP3vrF52UUKmROxHI4Tj5YiQ+N
dype1BZUTNBcaUf2SteriwSR+KYEMyXF/RUwR6wKR+8toTTa+xHekMNSIaWCe80L
xl48EbfiW2n4pxUxx7eQsjvxHfsjApCUr9vkNHVKuD/1hG15D1SbT+GEwY2L8P0B
l9rJKLm7oOFvUiVsmFXAq/cbBvP3XlJ0Ksh0/cgX5a6Q/Ki5Ih/qehgrgGQMNuPV
eweD2SAFrgkQshzAb6/WBiL/Z4f1qlDZ1/x8ayZU28bOgFcDo0f6dsZc2hp82hzx
KfsuNsM5a3r2R4+r2H134geyn6y9e1XBwyLJQFOpkrHgfIBoofmJJRUfqbKDBcrh
cRM4xAGX1Dt0GAODZSVRTY1zFpnEeOA24qlCdu3GniGLeUOOMmnyu79K8jtU8FAD
s57gtnkHrTCV+zL2E0mRvkudoSys4KhyocXKZ3RYFQpG+lcZlIexLKiqtf/1mYXy
/OvXVFuw4qizgcUkcjb/mkXUlpPEp82ZbYdAbuF9Hhf6ThkgzU7B+yeIyNrDS4Qr
IMkAeVRXkk/JfZEPTh0YPIE1Syqr2x/WT+2+Evd1RARdClKeLGfuvfKh6UT3p/ru
DBGIRjJ602Jvt1B9IHtoi66FY2ray+GKCI0lmkR39LUd5sGWciT+MJwszJLF9NqO
QXNClPdXSe+8uz6cioVMaVFH7eTB47amjNe8m0vnkPEod0oaqtzQp+Dl8Ue/ReJS
4rDLpwV4VLttzIQ0t/8ArGlDEVFYcuIx70eMVNSuLsFEYPbkQ7HEr3+oFdGHupmS
naDG+/I2pVF5/qO1L0bYnhs2XRK0BLbNetey3uHO5qIn6MGHYPDsqF3JBc1CPCKI
zs/DfXJeBIsIYDzWQdPClfSFg8gtFE+uskbGPjljGs0B3ZMeL9NFge97mnfR3Odi
9AI9JtI3SwkGKrgL2Djx8X2UM24wxyEEkYeiBT8iYYXPjg/5QZ3EKBtYjNKPpKLp
CrOFcnopQKZ1Dut6Pm+sF0ccxRbFY2a+19IlPO9C1HSJOFBn3cH08mB6PPilJW1D
tjXfTUTEtClhoSczUNTJUu4dPQysR9kbIivCgJNfPPlYp+MKxj7PJ6MYgA8SsOle
QFIiog4yqJ5igB9NA6ASfX5kI5eeurbeT1k83d1GaPzE3Sm07f4VRsQJvt6lokXf
SWrglpfvJkZERRKfa39QQxFwe4zsTWXAfyLLz/pKEbhZaP/jRUl5DeXMIoWsUHVk
py+87cy1HgP56SS5q6ZmL+5D/pdNhAe0hlPLJeBUBIO7movNlag6ycT1O8C3V3Q+
WJj/JF7n++rx1RUXtM3w8hwezKOBG3mFmfwoKF86yK0QEUiosCV1YdbeT6wxsn4N
gKEUEyghQNCaW6Pp0+2WJrm8P4ECauVaquC/OdCcsyNlCdL20JKbiQArUrupIcKo
dac4vsDL6QpUhTzbNzmdn8XVDhVaqXB9vwaLpuh7Os3j2ghBaYYjy1uteNJCHLv4
9vhfua+Ynne6Q7cbb2qYGKv8yqZA2Blf61K7WC2gRSrUbhVaV+VLzJltQWpuL20n
VhXchbhZkCZ+Eh0g+HEWW+iBYbgQ1g0GgZDVd+HD1q+djSei4XjAoOlRvpYlBs8e
2C4nt9MvpyA0d8LV7XbalgRfYvSVTQVdrTAKcPmqHoD4yqm+2dm1+5CJBPuoQEr1
WenG5auc7oF2VWWKZjecYQDoyQFffvUW6N0O/BjXN6NAN9v7iX+1W6P4AGC5j9BA
8DNzRrnz2Z1yOr1B59jl6GNH5cuukwyJe5TzOxdUX/+ZsXVU92pwqaOjYK62Clow
LAAbuooppi/OVx2pwtWI3gXPXgwqBXDQAdSKMukOxIcNPbZMvEyd8h7//gpnCGNA
M0likQ+fbHXngFdBCtxOUIYR3FlSyISo5WAhb4I4dwdkfleSYIpvo7+1KduB3KZB
RWCQq7s6N1DKNoZw2Y7CtE1haib9/t8zheTN5LC9A87pN7+dduEQ72tQwtYjzax5
FGUpdrTqysKD3+Q5ts/OkIk3ROw2tWLp7fMpjbAEl2xneLLePBL6D6EuCAGyPGY0
WIhdvyZl+y/symYSch3aVlDvP5Qt7ici2nE6DiTKgkV2vIgeJ+B9FE/Pf7cxyFex
ZI+NwY5RUFCVvHj+Z4xogcbyLJGxgJGbrrMi3XjZVXYyv0gRwjtUPa/A3RPbL0Jo
FwlxoFaTL6r4B98+raSjdrJLJ3c+ZwVEUHQX/pPJimA79yn+Ceeqc2NdB8G1vFJw
fFKbT7xiCeb5Zcim9v55bQEQoy7vZpMOjsTAzRyOs9Ty488v2WmYYa9JRja8w64Q
Dvc9gBGCy9LKnnsvGuDiaGTLXBdlHxrqOUa8EmJXmQ66ETX3yb9p8I8RDb6FpLg2
3dzVNbGRNLLk/J5VmDTNA8PnqTBZGGYabznag78XmosWaVOBwmcornpYmKgYAAk9
dTPPvBbcK4f8tDonVzkDm4cOJ/LqCgldwAjBvme//es6UMF5hCQOq+6uqrsz4aw/
pwRqav7RwuRcJHyByHaCiM4MNslvTe39bh9ybphHa3SrmMKAZPOi8/G3lcpOYcCT
8Z4oZP8Fs5t8RV+Fso6Y5QcEIF5VcePRuhToUJvCMiED9rrkxJ6ZHm98kjXw0N1L
BYBPSQbSPIo6BYzUJiJ/YK+FfG92jSENkFAX61Lraxr7HVCPVHgudknZ6Jl+fzMm
mWh1ej+8CHw3b/wzxmFL7oqjbT/kaFqk8KgpAsb1B3pLn0UJUasd3nbIp/0rmGey
sSFCX0h8+f9s+oPzXpXmIr+gIxj2B6vR8DLe/JpnkWnkhhOV7IyG0cj58LTm7xeY
rfuWUyw2SyLKJ1kwa9jyqwDU+poUwnis6MHA5DpRzRhdZK+KwycNgQvKIswez+JI
SvLLkuBz4623L1r9LlKdLk6pGBKIvt+ekvtlF8yu1N2poyB+pnOy6oiSqHVWnscD
qmXrMZya18ivkKVmZEvNxeTF0WwQvOHQ6pdPm1BmbilghNdB803V/K4uCOFJupRI
pGeuIs1lvvMjycfVrOeZT579NLcSB7Dd2DhndWfIIphTrPynSOEoO8B5/t/kj9Fl
2nSDxsjy6VANG0+rERbCgj3MZ5JoGXOQ2BnbD6X47cu4Ks1ynJDq9IwAhlotXGdd
YF0h/jwNvGDJ674+vJOSWmDLZ8Lz+as0bWa0Wlt0SWKuyIjV+utYa0EBbW3rnEQ4
Bky6vXwR5P5l9Tw907hjdQqqvgo3ndUbWCSSdHhqeBZ3oqm6DgP14dBOv5C8YU6j
gbGi1kPJzgr7mAjmR/Mkibc00Aq+6V2ZKDoBLUX4EMxaDnip8wpFTZtUc7stYxE8
LNX97zGm40FMAgFOMnnVfP3pR0lSvapDb6Z07cQXoySskQ97FEPF1dX4NA4RACcg
keDG3nS+Ow7SRCFIToVMPEjkd45+2MJKe0vie25XzEMSkqyFAo7UI87bpqGMpmiQ
SsaFtmB7eS7WhAX0liZt5QJgPZqaFLjeWXn/FFC85Gncn4CymqcgX6KmsG9h7ABn
LpvhbvaYszo5wXVhvHAo7HdAgdUhWECJ2XKL3A3sxdU82Rx4rTW6mTU77l6UAQ75
T8OXlkbKhEyDRLhHuc9fV1Md/7daUTqv5vsA5r3ySpyfeOQOnnYYGNAKSwLQh32V
5VVxyHlrvgZWRLr6XwrC1qio3Vu7BkSppC0K1X75RsZ/TRuX4VnLL/REQoEumEP6
8yMwHfXsJVI4av/aWByb2LytBEJ+zGLQ4whsxfjyWiuYuHw7dKBI0UnzHPBrbdJb
eoUfkp/C/A2Q1qd7xtx2UHffmmoiEiu6flOJh4JjkNOJkS8F3qw5J6fcT3NtWvbt
+wIwaGXXFT+Dc3kP1TQgxyQlnTDaKaomB9nFqsZKPZVfogHut9df0SlYl2Bry9Ot
xSypPaptbXqckkCOMZR40WjkN2uIBLtWTbS6XUKVrwvKkebfEcYbwBNuGQDyIN1u
qmLa6xt/wqKp4BA9Xctqf/39xyRDGJWxxCns2asvThkpEsnDBzAgWqa+FNspsuAy
nJEHI7cFWBCUU6cxr7WO/9tE9wht0I0LFtq9VMSp+PxBn3gE0uhYeI7Rx6k0ziEp
LkODOvgEu7nJXXNVzOkoR5E6CLj2mPZiL+r6IePsrNgLLBBkIwe2vP/1PBIYEeOP
RYNhDI9+7AA5ifIJTqLOpDxWDdDEJ5ksz+GVYiveK+xhYIz7eQDJdil179LbNdj4
ZqTEPTPAiJmb9tMGy2ivos6Y+cEPwr8F9saSmx3b8lfridPW6sqxxyWa4fQpk3rZ
AeuYozR7Ok4Rj+dQhgfYPZSXEm4sy0mwnZENgKGBRUYEHeLyrJqVrO5Rjjp/rSZo
mS4bSLPVlUyIzaUwq1/nSQONUUWOOQrVIj3D0aKnX1wrBlSBbxLFGMnrT93ikIWX
jHu3AuRhpxe5fc8ahkagirbnmgIUrBPfZ9rCt0qtkJYUnL5qqXnPFwYMVazG/g5i
ZWJES8FLSZOZOo0+nujZw5hU6VOh9rX/Xq6mqtnUm1ASRdybHg8/pA8cpOPYxKgO
5PhYV2h4mLDJCfLOv9HKi5H0hPFwxeMZCKmZUORV2dpDJm9/1oKu5AERv9qgcj4d
Zs0S+Fs/RUnffnlz++5TIEID1QkIC1xMKEAUEF+m8ePYTXU6IG2lDkzU2Wu8jyzP
MNSqtgOvYtlDo9isyWzkUt8xwrSIB6XvfEnfPhTs3nMduaUOCIvD04rrhmHij49/
b5Ia3jZzVFXWRS3g8YA7PaQYuUb6mg6lDvMFHUgXVCuzoZRIuFhVtST5wHn/qIWg
uTHOydV5OevTkP1JLHhArzS7H4fyTO9xR7V5oz4Qr2EmHn3mm5yJa658yW5yk++7
MkjHDhuOBYYWQzsYXJQb37s2E9GVn3UcOOXy2550qiEbed6RcnGrUJY6ygHhu36b
tbo3xEVqiQeusOWY6n2CLqoc8Lwt0P615jl+7Z464M3Tnq/So6KbRqJWlGp6fSN9
QNLRCeLus3CWRTNlp9W+N8OqpMlQOVhqWYx0fvUoLBj/FZRDzGirraidM5PsfLkD
YXKdNjdHBwbI5KOjEqOJax/fXFPXYkhgTq342cKI97JRI69ED7W1Rx6Maa0rPe1P
KzndqLC71bUDwrpP9IFs+NUSGjHQYjCQPVjkrA6lUZN8a8olGU3/v7m2ccp/xgxJ
bfRBIzmAoE56NDNLC/IixKG+mX+b87ZhUF+DCf0Tk73wxFhNTuq+n2XI302cLn93
IHdox90LD0b2XnsT9AwxLkYU5fIpOPcCaoWeqgRhdmrMGi8FWK8Nge065DeBMHmz
rbnswfjWxleou5cc8M190cHBqwTJtEKqfBf7kuAwUoNcrjrBJmjhPDxFgLcfHQgq
C/PeBFVNwA0PymXnBDYuCywwllrZHn3YOsk9GbkZT6TD9Uz6aFxGtWJmEI4IHmd5
nFDOr8XovLNmi3tPa/dkqyT9ry1bhG7kUyBxM7z4Uqsv0ulNZAhUZpwG2sEFiF0d
Fa/i/ftb4WhMVNxuatrcWuCJ4nXcwaNjitaCyfyEaitzu6LskZJQxVPpuVrfihV2
jSC0Ko/CyqMyEY9Ri1cIdGvjSyodqc/EsmFiTYvyCrXNtixLbo1be4ggnypsYQER
rPlBvs3Bi0bIeqVom6hfF8RajCcwQL9N//eTpMEaMtK7EXIPM5N6Hai2Manq06Dg
KhCPjWWoQ2zx8zCqt2LTRotTQmKlHnewcHPj+6prAlX5YHI5VIFeYchgIqAfkcKK
s8QcsbyJddgkffskWARvVTDX5pen6Wey6ZMP1uKbjwkbhtzGWSkBVl3GOjqA1Ife
46P/dDfnCeJQsEfHC4w4kTwmjLHlZszaYoL4DvWmH3UVJ4TO0tHQdOs3N31w+XFx
pMW/JQkrRO/axEqrfUIK1JErgAqUg+sKEj9ZoM56IPXBcy8wyl2x1ufrKvTBEw3w
6q4L4IL/zSGKLcteB5ncsZGe9GR90Uh87igpVoqufNWIA2MztumRDrlFXxlmTvgC
s05/YaMlMfAbHyDmhfjIyrQx5bNeTHIzSG1EoFLG4Ms5H4O1Rz/5W2BuLqnJ4dkx
AG373uHa2GoJwFb5EasyoKbz6vbyWD3OeOL7uOLWMLCafcX9nbDQ9inEaw1ROEIl
y8eaJ1lVSsBsTjNLkcUND6z8Nn/9DwuphpqMvgBj+Sv3nFeFHUckd5IofB021I70
AzEebtVfMjXLDXU7m4B3RGnMVdI3VQR5x/ItPnhyxbiq/Q8X7Os6EsAg7r+fKPPd
PAp//0nXUyFqPzxuxvKQflPDZcDauT7LenTYGjHWkBJpsd/SLOYjCuDf8HdGMmYz
VCzxCqB7VCHiYMCtWzf7ffPk0u4NsnKs4g3pmpWTg9hTuVZtzzFsLds7eb5YmV0y
W3Dt0XKgKkPBCReYcONwJagx/OaObScqn+R4bmggkehRfTG4RaBWG+ABC21wJgr2
NilNzSykoY5O/GGrznHgCyqiybWhBU/F3/l5JZ620eVIK6iz5mgja25ZJIC63aXD
LMCVAm78mx4J5qFy+09QhYGjjO6zyd9wSbt1xTcMhosJEuR8ExnarilfTsj/fNgh
4ZDNULZiCrAbleZUB7mkW6Otu4S5LEM8aXmeRdb251t2eAu2m56SOlY5Sp2YZ375
JNPHFhA6JD4pqAJpv+P7XRbG5cyRRVuzNaba2S+JTNM/tA5YqbuVEozIwVIcEsOF
kvsZbfpfbXd2uZw+4mwZBmKSaJ7DQckr50rH/krdsWdVvdGYxr9ZCz+lFEY+iVQC
HCptC0El3rYs7p6uEs9dx7Pfakih2yPMYPX8BeaX1IOGVz/I18xviYJhTLNrVp96
htuN0DYFhg3wYXOKny74xflr9O8ftz6EAVVO2DGwfN1iWlzL+MArt66e87O5opdM
l0ZqO1H+Vb8lhE4SJ+M0i7OV3LuMHkEJ1SkQ6vH7VuWLW2iyiIBVqtZhdOwJAFlP
AADJApKsrv+n2vV4v5shxJ2Z496QRA6LferlonyT+BsCzUI9jtUjG/knSxqO6EuV
8MAJJIjDsqSOPfWZcl80oi02dCCgovmdZ+GnyhY8ERQ/GK+aNgf36cRFCEBJN5l2
vwl/k2rU7gJUeaDB46i7sZ0jNeX1VWCAOM02n2xFoUSK6r/Sz72ZGLpH3NkXXCVq
ogF7GZJ4SSUvfd/NnYXQPDmAYIxuvglhTo3dHEcvxeeYBkKbY68ZMcanM+RRvrX9
j+WssTDHyyAghUUavAThN2FqNlqqn8xjQ+2RHYToMDMoJp8gdnY3UnK/EckT7N7B
/OJtjCByBrfoO9D0vr3PGXysST7cpc1qZUnXMn/4qq0H9U6siWZmdkkTL4YgU5yr
6Rd6jO1L/6BOzGZVHMf6rT1zZ+rKTZo5pzBycIFgKQSfavT+HS70ivBUe6D4/oBx
iYH/OEXiPuUDB4DXBcwXyMryAPrSGK5r/BtiMC1GC692uaadUpdbhfglT1a74KTv
ZAfo08fnaQC9Lnz/7GeLUB8bZ8C3L+E4IYNHERx4g+pWEfuMZzXVu7HCoJLulECi
aJxIBJiDOsF95mW1Aic2Qqszufe+E0DmtBeGhfnhMF9+zp3ZPynY5TPLUVU8Un1s
q8Q1V/jgqu8uJjZABL5cXYzGcgYfJnM4juMyYbHoEVCDFCKlQVBTS/QJagHy9VCH
RvMT8x9Rig9ZBKP37J1UmnBnHjwkN2l0hK7ovPRl0GPyAqJl/+ZFGWCnirjY65OS
9KAqb/oqJZF0qpcnkjCTM0c7sDq7A/c5CDlYFRFgjqKHYTGLrlFSpF8NHqJocS10
PGWdY3jcOlhM0O5nsWYlAv8QDkdsmFRbA3V1+zSGFiIcVoKv0VHfqMJ8mdFxPM7k
w1BO41yMTCKrhU3qJWYP2rYHJEgTkNozsaXGyXJM+jcWdJOrPs3GEz+WJz6Q7xDO
T7sVTdHZA00MqjAyzuz4cUPrIGpnJnHxFNKfRXhiQ52JLTlMEhfJD4CCMycNE76A
2ykmi/bov3FzYbr/EEbstHkjKj6tGsqpdTcHpaIRXRweSRmSjJ9ix1OGzJ0Ypy7F
TvC6vkmyj1dmCPrstdyQ3pkecG4INDSbKgDY9dxPe1/S9rWmXrtiZK6G5KiLS+PZ
+jOhANBs7yS0Tj78Y2oLldBhuJBV3dqIN+z1rQ+HOhePEsHhCBwcI4EQZeCT15tq
MdbghgZ+OfbjmeHe+zHzG2jSZozde1m6HgcTHM4RLZIGhqVHQFllnOB4ls7ZOiNl
7lxL58K2CaUK3W+kAaQ6ciWKurWvlj1LnLDlESU6ocqyQAOKto2PlhSP3VINKBT1
N2jdLe2JPHxYHQUlHRhJuQFU5BPvUF3U9r3fKaVhUlHZGkKc+dYp70BGfsZtSUl0
OMOmcYNyS4u/VBVoD3RAaCHoCbg7n20KJDmZJgSQK0I5Ts5BuUnpOEmAWG25qiMH
gybbuUa+oErry1cj8Zoo4ZVOwEN+o+PROJgsRMaCZfYFt6dhBEHm2nT0h6fW8M53
nMos2pkuDk6GwV+XRcOCiri9OjoAQn0pKyJg5lKaulAuPvulPf6zcurmGWHt+Hu1
eyU4t+CvNRCjR5d9qRlYuZ7UtRErd4czAYyr2hbUK9GFxxBWNd4aEpaBaeLvtqZt
lDJgnmB2oB/TsTp8pXRPvS0olUm7T+bQt1KNSBitSHzGQrdZYzNixryOxAjNLulJ
y04fwWT8onYcSTsDok+Tb3jBfgiHrmH7o0my/hmcHuT0nptkwQRvGp6tp8oQ4SGr
YzBAf+JrqZg+pVVsb85ohb20dNLuAEV08WA/B8Z7+KazkpkUnyjoegIvZ3/iGci4
3ltt/LCsUzPusri274FM2rUuNQh7jEPkWGuaHE4r0G2h7atlglBJxdJMkZcIEBDZ
jiOyIeSy6L2f3NiT46WDBU5N8cR7w7fyxAHPYumig2ZQXSV5cUwLLHS8aWtUaOjy
Du54GqHzO7wDNFlhNDqq2we6DlhfokellbMRGOXoXup0nMsE+8A9BcNen5TNxQqD
Dxh14/yvDgaelHb9ct1Hz0HZpup5kcx3XqaDbG1Maqz8VLJvKktEfC+4jw5NJp9h
DOYzjcWyd+vjcKqWgx42gFzjknr7nbSnbtIOCwzhPgJJA4QrlqpyIlHCXEA66+kU
U+Zr3zOMpRGNYyBybKnbmM2t+4Sh7rYuJ7NS+znGhTFYLweRwVmocFrxvVDoGcdk
HR4bxxqrw1N5bSN5eZLZxKvRpwbRRH8Xt1GCR5ECwdKkwMuks9DmMRuKJRKiJat4
i++B91qmoDaAWQQPzw7h29WOQnvpjIDKw2icn/uhfL/Z8E1VI4O0vmqAZRzJL2pQ
XrTmB1s77vnWYcViB7vc8r4+Gqs26ekf1tllSdQ6tONWkt4IrHO7F1/ho7sWh7Bv
oa215tmtRSMdwADJUXzQL8oUMY0GW3qKgcZNAnczsxU7LwZOlTUHnb1oA0PaGMEW
982Wvj11fHtPNnegKVNBfwSw7mvGhaILJVhfrWk6vzJqpxmjS9AGAe9z4+e3oMJ3
nwRNrWhByvaIdqm/FjEZsudy56wkxCDu9Sx24eaZfdYcSBv9SkbSjQh8nnTnjGyq
+qfiXF5YsAMelcS/ce/TIIqHszYt0NQ2IM4vs7HCpIwqiSP1MEVqw5yO/kSKxVgJ
T87EeIq6Tyc5z/8heTh/6kmekvt4B15htUClAIazpB6gZ3GbmHU98mk0z5sMTcsE
WSusmu3AjgWYY/j1cFxFsX6ZY8+gymYPrACiNXuv/WJymtrtJXeErDxIJ3mhtDRA
X2T6739LLl2OpnhjdO4bxFBM79abnyHCX4uTn2ur+eJrCDgv+iHQSjbwloX2Gkq2
ycrgOoa74cIMNfClrQ7MRNHy7Zi6+h5DB3NEavkozmES32QibLFXBdVPGSzRuq7x
vtZYVE/RJTow/x4a1kNkf4biCjnk4YvwgM27N42EYv++KbyA/vo1VJ60t88D/aDT
FnZ+WtUDO4rMyTC1l3d++q14OeecgkBWLzJrWEtOTngD8aDBlPleFjCTkry5iYEj
JiKgaKNVU3ciXgyDxSmvxuMBL2KkbEZ9EW9TYur4NPtScVMFVeoD9OiynL3bDUUA
Onj3CcuMeW3BAHNaIQFgI/L5uFMASRNiRK7tiURl0XhdnFBX3Yla/7BM0RYQ/tec
cechpbauhyqsCI4wpANoWOuJDfEN2vm1R4s39HUJlXXUmvSxxQzWUobKbYIOMgSG
Zmj30vUbDf9km/o9UPrwnm1HpowrC5gn3yRzsxPX5Bvoditg+4kQzP12/cRFluPK
opYWHDZoI9VJzhoY1+h5rZbVTD/CfSXH7XOvHZ/FOvNy6NnJm2dXlVHJF/0zyiUv
g13HW3aE5aVo8SVo2iS1SN2a12Azj3wKUmORKqCkeGCiqirQm9/MAduORlARcWzE
iE/bWw7XWmTx9EY8XLm0NWX3j/LTj1hhwtm5NP9tkdPpbXxgQpHZhteVmzjTcC0l
jT4DycSZU2H8AJBASyiYk3LJbww8Nd/oV1MQYK8QKw/kgHrUxuC+QIFx9dscT/p5
sd0wlGQJxcKsBeCwsX+GPf6HVzlmhzU/gWnI6eZfY6/5SjUfmRVSh4oG2JIuWrlk
vLj1BDufJibcdoqEffsNPyXEUnDJzOQtjYFcOObyCmbfdsSX2n5vF08fswB5s09F
MEXSzg88iomnQTNU7hFo9z7vS0QC27re0mTuC0hSHIgbrksdj778iExZ1qxzLZ28
oureTw7VclzBg84IIRZRnZVE9gE6OY28znPVweWa/VyXhm28eQsqyWtPFyYkCbV2
17vwhCNw6zhh/hesHd274xhtbpqsU4BWB1KHUmf3tnCywKru3rN1wZR+iHs5rBCC
MGawjjryvkN2EEhWXxDJiPxyFxWBqkfnVDukMQBeEW6DWjnWF+FVk53N4UfVw9zX
kmei9+85zBauKwNgzGsMKA90RVFaRB9aZulEj2sSUIcYF9gEkrbr2j665eyxdMvZ
hN6KhQG48k8n2aRksT+S3Ku5V3PURCl1ITOkTh37MsGef8/dNaK9VyzUffofAG79
AFHYYLBOSPNCzWuQL5E5KH2t1FlNM2dB3nHnB646k+5K0mHx184udZAWRRoeymTw
6sIN6IeQpvRhyVtZw/goLgy/kl1THUX2E3EACcRY/pCpCDL+IIEjVPDrNHFpU/3x
Kh8kFIx18Zo14Fa9ev1z697QO/NYxbyfCV/IMR6Hw77eJlhqiVerXW45CrRBnDj2
X9LKteiNTx1Kh4wzj3TJyg7kgXMI+tD9jcHcK7XH8QwzomQFjnOfiG+Q/OrPd43H
Y7OhPxFdzfeeKLAsQN2TD1rN/04JJXg/iOxtxJ0SQBnkgeXwYRgfAqBOOf6vy2pU
9cAIofktgzkuNmH8h24sqasf710Jw6VWpKEyiua4T12AFIjXAz75J6w7ZxKrppY5
S+cESPPu/R/vRvPZrOM8oQ/QIotz0XbNUKeSAET+tIbiY2k0IY4/RU1MCQomyetO
TAMXZuMty9nGpRqaiwLb7U0ZDTQsakjwUty+a6+h8rduqg/7XRGWeEjfXgUccjvg
BnqhDTyZtb4cl9LEAU6UKaX+27cpjZj8R3F5+1k1CKY2HZwSkpE+EZNFrJEc6VfJ
NQ3VantBl/jWht88WsapyQL4iVkQ8OHjlh+SsIAHpnDCHbn43ezc0f6BumcRo4op
H5vN94AvAz3npL5SaWBh+HfQiKXynVRevgTBCEl/OUtzK/ITfsKgJfkwEkVmCv0L
pugjiR7/9RcciQxWHTulnUASRBDBeS09mTx3HZw4/kaug8UmRyYEQCnlSUHrExJr
kYBPTosnlXC2C4BM03lc0kiBALJ/f2NaCTMirea/BQ9P55GIF/M8Be6S9viknw01
sKqiNAbI8hBSdHOEtKREy/GM9w8YvRJOId1slCbpGodkYPOJ7i/8Spuogo/GNJld
DOzZdBBq/eEW5QoCvRw41p21iH7t+bQHW2eZYcJTQeD63yu/065KkL3rKy+Els/+
/dS/PBZPeXqxBNZvjgEFGf9Sd/lTRw6sY6mXB5CWVFoJPtel+06r7FIqyu2tupY5
9GgZd1iSprEHe0H0WqnytLp5uXEG0fzwGH1CUO5AjrvQp1sawo1qH8pemSn/qSoM
ZNZY07VYrRWPY9zwiaIHaqUgkbx1UWuMF06aW8reHbMdwaHMUjYT3WoTZgO1j0H1
LlhUTdn6iC7DFJf6XNOkZNEdSCwZNwJ0KP42xPhkGccYZmpr/3C8Ybhq3dHyAJQ+
Ok0JXKFUcWSMzA8kdfOWjSvWb3uq6SbY+RStSlIpCVxekIRKQYkogPZZt8As4oky
uPiCiLSxjjGj8A7z0/yIk1kLd4Mf17g7QM5zfW8IBAhyhTvyGCu0202Qz4LviijX
TUq78bb3UYRG3LXr+eh8PS/oJQ1/U1W4GNjylOwV2tM0X8M+uYaCY//Ty4ULhYpX
s8Vfs6+Q2kZND01kuqUSvXfB8kJcIXM+a5m1FB7eOHCMSvoqc8FlcWG/XiMVdVAZ
zHrh44GewYw/lEhHiurz+B/VcZCtfNNyrM4JK/IYHDOFDjejUNYPQbeMAs6B7vQQ
FPVbnmxCl6ZohGrVUf2k5Ef2Rq9QMkkrtSX4IU8r4J2M695DQBp9qPVHyIEbyih3
WPqRWcWa281jQR/FH0skntN0PHIPMmCsbruBF3T5RSL1nK7Wyz8Nrgcm/HBrEyH0
/ntnB6xr3gW4aPQ9Bw5qYu4wwqwgIksTUze8ds6n2xhL/mZMLYnsOV8aUw4I8YQR
tGwP4CfghsmU/73eLhh2+B5we1JEdDazJ4C+u6fSUEEkAAYylFjY7DdVEwWtkjl9
YWkAyuIIYjIV7d6gqlVQ49jNjMWzdUnXNYteFoQbzt5tQsumR5V/1KSdgw4wwmB3
3zbwipTwzQUB2xnNu6NQ6muzH6qVpEy88rY9TCJSCz8Wuhyy4uE5+PdOjKT7XaQ0
Nb5pRDzVpeekFErtBPkinpBwLv5ZvUYwOjlWbOfBFiwGM4gnGFFGk2ts4i9lvVmR
S+WF5NPJeJitFpsTEnlNf5/S52pHfg1yHjbXtCD5O/OT/KE6UwpjZnamr7S2/0z0
j2Z1Q9UikybO8XmbGwidBREu23ftD0Rz71swcJYKURJDCuvaZNapqN0NJ//9DWs4
UD5xOd3wJxI67VG4zLcBZu2Ma2YLWkK+088wkRwkZco2+9i33/jE/F/Y6yIlawKn
koQoV20mY7qT58dXeG4FD02hGW50O4zExLZg2DdO0Z13box7hqsrlRgmR39aRi+Q
WyuAGzskgOTIIRwbtUbq03oOi2PKrHQAFqxcPgCTRt2BKCS186V4XUEyV8dBDH5e
XlgDxyNy5cXaVFa4QRsbL7+RJGdDoWZdo1FYvJdVDTrVxyBhMFZigMvtffvBzS1r
c7z60yqQmfaHB5IX+jpJ2M2kgUxOmtb0E06XJYghxLKRtPTFfThk5WoaBkZrgDUQ
TTw/qV1KgeAt29jvBiMC07elKbYM4oKtkQNlnYu0e6sC9WkJ3MjrHN2lgD6M0Y5p
r+ODudnuu+0ZdxvITAp5DgLDbeVzNNimtaZmbmdXU5pAdljnDT1nXJG3jwQ+uC9E
fK0t1bDUvJ8jszR5WTWBRfS2GycUf//FDvl+uVGPUPnMvt/1jO06E4yU09GgKHzk
rR4hwxRvsXNZbmyIKP5hC6wBy6q6VWM8FXZUdYqEVZvgW6ytFRha3R7JQzuyhbKL
/HKXs8LG4kNsNSjyKMz54cGWpIjAWQTV78SeCum08JhPK+7vFbDFAC2Bhk9aJiXv
IJxFLkyEIINRWQuSbT2S77oNGb9QTOJM+y2l1AX/2TJCpJ9xZ256DvC4WFogeEQU
ImXNAxfy3nXn3MBOUSsp0tZKD36pzHl/2sqKhGixsH6OIcbBBO4GyRC2KeY0oAsK
GEGF47Fn7YFTr+rppkLlacC2UkxNORE9352r+PCya1JNlcgnA1bDgJmJwseViduE
ROViTdSG1P/iUw9faG/dQ5f51cum6fmJNKezh35Bo1kLXKLdk+P3Njr7K24bhbX7
Yl33RV9j9vamCejBmuKTuRfEBdvAG7QlulbUO6u0/D+lT1LJMEmS7tOtNmsEw+tj
SnFsCfP+BXSP1aVyEaUYRR9AyUY30AOdWvfEgL2LmZMbnUtc+qtAl1CJJJLGZwSA
0B2LDnhjoPyXDjVfY+ZqM5chpi2JeTvfXW1uKsF4nYuRFIF1AKr2xBpPLXrBaxYF
ruKwkDBelZ2md2AZpnHO1wrauWHaOpkJlsznTDVXtrYiEnVREzuN495NOBmiTxNK
ctSVE6pMEi5EqN5TtOOyo5Ch1BwbRsAW15fLdxOxfKWRJ57mn5wr3V7JrbFcZG/P
oh+3bLS2o2ylQG44d8IR9lmrmVpzBdRjfE4CtqNms8fsvd3JG3DW60DGte0A9h9q
z355tqBjS8KBRqOHQnPxb3utzqTfa3czEqlXS9evkc7DNo+VTajq7j28w8w8Axk4
mCyzmQ45dANvfdpNQztX2orup3K5hYfuG5NQUVZlM2UbVESf9lKA59nLHAV+IeQq
DlJIrdehm7Tdr4aWM495RPn9uIhF9RUYg5PBrTEaZmGvLei6SOS1IWkNO0q3ghin
BaMaOnfsp9eRagvTAgr1TuttzEkXrW0gUyniKg9ra9p4qDVoxwodjutaZRLzgVUo
E0XnyovA+fTqUXuttCEscQh10mvOIvEQhfg7EhunbGfyIbQEFxKoYQ+BThNeI5ID
DqTd4MxhUrHHZ9i6Jp6umlVyrhaoc4HWncdfSinOj1Eg75BC5gGFE6Lv6psDAQD+
X3e+WjyDzCCuwgLIV/hdEFYGyw1Qqhcp4jtP7feND7J/fUoe2h0c4N90P1n6e8zp
iUAfbSrBqZUhuqf3q4NbWIWYBYyxXR5LSfRUGqCdynSv/WXFh8nXZM18D/VLbkGv
phL1QlyASTSFj6eiVfD8bFiCSjmBXFSF0S1dFXBKm2zWSmjajVdglYdd0DZYg92B
NiIbqsHCNqwOzRRtHC8agokDVdAdDB5qnaiJfHa0yeTBrvnjCYQ5IPMWg4B8xVPM
Ff5EbWGSY3A7aoN9WRmiO1S6MpvA3ZmlS7scl9E/YsGKAT2TVTZYORhbO+TzQSEy
rPB2DWw1wyGUqDnRLDJq+nm4FDH/Dl7gRp1m+/iwkJz3f26wy3i72ymI6YNnUmpF
i3VzFpvUoyECgh+4gmHyDjLBCKA6PnXeChPlt3z9DSSJPJkXz+iwTIULlgD+PLTZ
Kx8FN3tpmjUl+6mB1r9X/dRd6OHkNbvJCi+8zqf3OukcP8YI3xFioBrnWqW6wlHm
o9O1mkxIcqua979swfv4sdDSRCgFmC6vP9K1ZWIf+v7EV+pUTg/mz85abqnPdEY6
WBuWQoda8EMRsLv8ZD/xXsy/8kbHwHCYvuFuQiCcs06zaBuUGPvtXUVFaJAVWTI8
DhIFeogRIpy+FuWpN81OHbb0o/dZty00TJoR1OyButqbCHA2UOtLCsQPKUHDttpc
TetJxjFnohVB78zzbzzDh96arpIDKBTJBr8wSEZGBigUKnN5o0W+cZiW+bYc7TLY
1vouy7S4tT1b9CfQtKhoWMtxUDoVnoofgQU5G2VemoJnMCvVET+aKjQm609/+CmP
6qtAxyHv8CKWSllMJ2VCvP876W24kGgrh5bnwnAS/qq9AMCdnGQUJ9xGVwHqqdMg
E+qJVI1Txi+0iNflo3V7qa1CJiozvPlPX781aNs7XZRLFU8fjOXTadBL5oBqUXSX
WVE/F7becQkpeG2/WVX8q1HEsVOM2CPSSNRRxJw+oXRfbNo2vd3Lj/f415Y2Uheb
6c4SbqKWt8SMSmx4cIScGCnvnF3MAC/SFNE0Hd43xlZnsO6bIEf1oSOpxmMpWP44
MxIo7XfDjIel2BcnKebIEqBxgOC90MXQPukFc8b0Y6O5FBYAfE7CuB9CbRZ7c1dF
MTRqqjMFEM0iu6A+wPHIW7aYK1C5qnDHZ8n4XN9iYi9hCSZmD0FIqngUNRpuIF/U
ZhT6p5fIrEyLW8whvf5r+V6oGhB1Y8YzDmP9Ep3LiCTIhOqni0JUCGojHXCuW1bk
uqRW0yFpJF7sx5/hHQdy0xkJuCd++qGczgHiOkBlFKdJ6WwcqM77hPzeBLHu+zEn
mAI+uCKnOENwMdpxy/8xTANtYSGXB5yWpVFxCrmLMc2eR11puLGRRjK9JXZIsweV
QDQJ1XzllBggNfpc0HsXuQ41NaTsfUnLIUJbf2aO9YNhwotn11ODuoMEQi7OWsfc
3J81LHuUwXSL2jnlW3DRqOUT5mw75HU1LLdodMVvC7ykudhTEG2RJST8ztWsR2wU
WRZ5TGKl5dlehnuV+SXav6Z6Z2NBQspTbl+/9XL23r82Zt7GYCMUXrXW8zLRwFIs
fjtmoWNd3+WmYX+lrtEdG2P3mHQw8uMKTc7dQG3TK/KMAoSRR+m3cm4fwFpRSDlB
M6/bD4a9A0zO1VYzwZK0Jz6qaSLDdcdsSlr4UFIBGSKS6a1WNNTP5MpB709LeC8y
BLjrjzxg2NbPq21VwFcohazVaSgOnNY3CIp8FBWzQUWi4xW048w0SPBzjJ5pmVE+
0o0RO9TxXEWGOrUzeIgV1NMEoKnA1Rq3IFoDPihuA+kq73mypPLPOckKEUjLM3bL
XJafme6gX2qA8eGD94e/HiIDtmVyFgi2SPvj0lUCFyXPqHwYivfXPIcQ4Eov9e0m
hKVhrmTJfvClNpn1n21FQ6wkvxtSTUD1IpIxhX3PeZX1mteWC0hDb79zkwflcBki
IQWWxdGgaOzEmEFiZp46XwWyKvhZL1PN1elVcbQoLzpEkbGkRF3IDRtfsyn1LY19
v2hrF58wjcAynKBSm+hIkWQ9k7lsKHrclJdNhxA1VXJAeXm82Uw8GEKD2LMFQxjy
vAfgRpjSePSMrPFdM2sGa7NCIUZu47pZ0AjWuLO4WCDlGn+t+Prz+dJtRyVhs3Db
pNpbk+U5BP/E/ogHwgdC01TNiH2Bm0zDbKYG+7vUhNGh3DZgak56chuHtdKUL9N5
yNRp6unhd0WkYfNt7MUhgbyMwjXY2Mrq+8wRbE1Eyh27LbvjV6vCQXMvPcPcuGbu
CNLlh8LAL9rOJ4nxQ+oogUpguEqU8DGaTjsitZ3BxNTUSHeY6oS4mPWCf8nsSBdA
zeripXXTFYQ9jY0Ena8NKdu5IoJAVK3I2xraRqnZWpy7Nt7cPWmGoAjyVDJVSmni
PYp1//AmdjM0dkurNzq9DGiPNbfGp/x6c4SD8wuSPprQcHUcxpZtAfyR/wI7HWWy
yOKJZ22eKplN3c+LY1KH7Mi+fTy51/L7pibSkw05Jk161PpNaS8BpycFL9Z1vs1v
3BUTvXibIX3+nyE3JUi04cUYxULxuybKs5pFtpHA62l50sIPa0qYkGjP7jaPyNOj
L4NdxIp39tVcT6xu8zGNEUsGS2lgn+fWhhKL8v4VYonSXmKK5XRrEpBGA37AQSdo
ROhILIQRn3SR3wwAMg89k8ubFnzLHiJ5dz8GSpW4ol2buI69AiOs+zdq1XvXzAGJ
6L4s8CqDtOU3RxrJIn5s/91/LlTyAxMGXvVaPIBm4q33uzTlqRnecBasFwEeTi7U
ckMK9GUJBwID7CzYtvwglhXeVI5ouHnnVKaf9rn9+jUSVx4HlsRgnraQFVdgHqDr
ge8y+/2FlEtUK4eyXCLcf5YD93OqfMBaJU/2F8rxKePpK2qWhx/s1EKYMnZL1qrO
SgkSSfY+YLwS1ZnvWajx8Fl5m7iv5L3jJEP6pMlxPfF5RBAqJqlvDPhxs5UTHvGW
PUMndCfnsLM6F7S+pekJMuAR38tG7YoQ7gZzEEkl34x3egrQUHqIJ+90l+mZy5eQ
ooDO8YyoHMWgJPnBVNoayWHoIoywW22hQ6Uf8fF9E3Jqze4VTzC+8ac6XDQiwGqv
AE3Puaem8TqNTPpyezkie+ky8+CLvRZz+bZh0I93w0yVXbsMCLRJfI3+6Di1Qqrl
KeMKdZ4F4xZ/8gT8ahAo4TBvYty65BKwNI18bn4A5tBZim5ky+WYLr/Tzrz/Dexx
4KXoLVmlgj80BS0jdEY8IVilYZuZC53iUx3lHWSfBR2YN4s0eA3yZhcrZFKFNFvU
RBYBhe3oM/rKwb22sIkzHcI+mGVYboJzBA/KpoUNbNC6z+JEW3aOShvc6Ubi8pzg
ffjLhueVzL1BrVlwIpAFMzeaavG/yWYKTnGehVJ9MXYJ0UkB8hpwTSwVW9NygO09
SWpjq+ZqTjNcAArtltrNNFhVUENlmxncnn8hbRw559V0fJcKW0K9euLnjUP9Isfd
HGN9GrsKAzrL+g8LDWn0ymGUAPs8O5AYVbq8Q6/QiM12EujWoOBYICbguiQRNpsc
Jv4/GeD+DiLYbZYYPMA9FKy9PfOzyCdxZpKJ0w+vDWJ/mND1RfmXLY8f5Nqb8F6T
cpOT94agfd7yeCKeShDizZrKtAmFC+idAcsxNAhS8KzapPe5mDatt0vUR0hWdLfO
GQKGmCbvSNFWNEGL4y/QUEvXBl2eniWBGDcK671AYnsvHOGsxE5mRGz6AV5psK8m
JQI8+/OKd5duYiVgfjJeHQ4HDbVXcTlnEf/29DYP5+32qXDz8dFG66GkdnsDxqku
Rlh7ZQA2zIKpJ0tAcfnwxZmttGIigAY0ABqJQmXsE5z7kzJKALZqyKgz4DN/I4Gy
sRXULMaLKIGFAyUVCbQQecZz/NFtDcT1g6WqSsgaV7kODvzHyd13eq5KEE7sc2PT
Y7xEcuG7SsDKeAt1j+gBfwNISyMnzHyb3QGsbipJzIKoOZvPj47p4o8cFik1IBgn
E6SALqQoFLcPSvFtKf1XsPiwWQAMFSl1w02/kiaUMjffIsAFWYpirzhjukdnORmr
+nuAz9DxXxutHIkEHvt2iW3ELf8lj4qGA0nN/L3ShQRTu27Yg5SZEVxZWefYhjJ9
ccRmuQ7eLRQWl+kZAdNgtCKGM6eJ4MLdQ2tdAiPMOlPoG4wCexz9+bK55wA+coWs
JAUMz+DFsL4OHEUdfvcZQk2+VR6jlgS4aW/Pa8Yvchz7U6rbWKz1z0XCR4iNhNGW
ZvDj+phtfnmZJcQCrPM2p4RhnQD8FCIx/lEVHh/55utesvg+PqqLF36aO1Q2mAEu
8kij5TgI7BgtKQfHjw8wgxaznMioGLG56hT5i3E/YvJYIMf21n3zg2Oq/kmTbAYa
iK0eFhEhAD54DaQl7QPIRr6aSflQAtCbnAV63RP6AYTWxOXQ7+bVqXh+EqvdqHUD
3c9tu2YrrTSlFoKkDiHmf64o7aHR52+eculfIACgyl3xI3WKB7v6sKeuuRFj9kxp
Tx1lDCgPJolA2n//OYA9hAc/uc2ieedJqzVX98BDWkaNZ5SdWX2qKujLhgsqC0xg
2TCDYCsCg3luD/DCawSQZqAsxcT1a6wTR3lapOddjTA6QRQlhCFZD8Q3uGd9aGfm
gUmqwFmavNvG0/lL/9j0uNhKuBuY//NmVmqY7+em8eg3bGqh5skjBQpjc8dr84Pl
PcUVIcW8LhQJpq+TfqP61RHMRjfcN1uka+IWtpRdKJr1Cn0o33ilXiuKWjVIOw2u
K+MDzmLqNVdS1FHwe24f1OMkyFqzFEyRYrlD5nlI8eTdnCyleJE6fXiNcf7SUd8W
iPoFQsyCf64TWs1/un+CAyAv0PIEr/N03j2DUzIKKl4REUxsZ9HpsQrwkPM5dkyX
V7UCcTo/qagUW3T7iaQGnD7XNRXmMeDO40tSF8YTEjguLdxwugtzEdnl7YzejcIW
aTMkrujXGAb8jF5nZPH2zdEMn7Y6uK1NhI/9kwkc3DUy1F1IcDFBux0WGK7UjEIs
byZPvvEqxU2nWNBXQAWc9vcl64XYojuqLiBn6I4euEF8AvSuxW8uqN7+kb1Achfs
0djOJfNUx5Gs1fhjcUHAjjIJ1mDccjJDerao/536wcWiFAmBwzalGiTBuCTET0PN
w+Dmu6Fp1a153ewFs6Gf4Jeu871k/dS4zAqjQmcXh9XRIrU+0XnGERThylxHTuHI
4B68hZKassPkoFxrchafCv2qqfHpiKFEsCdSbRQsUaUHt1/vtP0i1aVzFpi7h0ba
TlwmyFfFiPG3t6H4I1NKZ7XktTMhc7vOYWWOfCd0TfwqMDaJXhLxL54OWwqiKXxV
5LL8/limZMkYV6zC9o3Q8Ug0Hlvetm42DADPIoWhRhuL4c4OINhgVss+GokW8TJR
a0dejos54aj60uoKPomfymYvs6T5J7119wvBQdOrku12QIjOsWQx/EjCHUsK1KKv
ep3aDxTwcoS2WkfouufzCxF+V9HwRPXcejcDxY8eH/WM0XDW1tngz/uWz7zKPLKr
EJL0uqAWaK1auyGtHNIrOXTBLQUujdki4RLVlouKC/V/5Qcv9OE1xgxNgIYSYkDj
2IvGHwax9K9q1NhnVwTiYR8nyK7d+6JmfhuF2w7udUypBGaSE1/z1Bbz7Xc0Gh6X
421YqNP6EIyPr6UA2lOnJyjM5PMRBcsoz/Z3ofBb8JDJjXiRfoZtUOyhC1TapuGm
4AkVaVvngBtDt63nnYoEt/brXbe0WlsUMPz4KJ9dXTXn4jUgPMt5cpd5PeakfKXx
4jp8uwhYrmi+g3wWdiKf5c4JRaOnbNYnuGGXkEjGOzetVT999U1g71Aw5BGuHC1J
vrRABodnjtyBgoLD99ELmvVm+pBFV4QYbGiKJYV/ERg3XCPk+h8IuLYbcHt9tgbu
tE19M47ITDG3iEDcljLT8gYDpQ6ypSsaeNCnLBBedN186VHMUXdDMaq+w0j8vGO+
+IEt/sWWY4M5lN0h2CafaoLHJhWKX3Tt+xl/pFLuV58YXGMjUtiG9Sfruu7pKcwO
9UeuVEpfRwOZsfCBwytwLBNji3dHJnb7fktv+jdZbXoV/852uQhdK6BrPfAkgWXK
A/rhEG5DQ5wE2QjRNRUvTLQ0ww62Oh7XLP+UKEdZyASsEOc6kQtkA1IewhYt2z+6
4vF1iqlgHDLBjLHvn+KeaTTqV2P/57IaZxt5IgG6bNtYSIXEelI8mhn2tzlWnMlJ
Xn6f83+f5rI02YhYt86epj2S40RXkFjcETg99Ig89vQypcFkPGWBdTNg1ligb8a0
ESp/8FbU0rvgorLvdNt1L+h9Ki1cTw2hlYst3r7/OmFUkekLItBER5nxU6GE9NJE
0JDM7z7/Uef2WzvGCoyXchOqQ5Q8/wup8Iboxf0qydVxPpqdJSz8/Ba6w3zzylTO
QSJh48t1vZ8W0F6i9TMZdklH6C7rIHaritlGKB2PyUdLuOAXRcgZ0HDYsCGmtAq3
BpGVVLnfhT6878w1Cmvg0XruNDbVu8PFnEt0tqrsScnFEkZp44n//FZeqga6O25j
Ag52FIsYuvxwH9b8bL2NJTUnLvXuiNWTSEmivTGDlg0N+3riAemOaTfGyf+bT+Er
XhMwVVsxFsFmSI19pC06bvJ24Ui0zqv9Be7hmNXywI85Bv1l9L6REkaCIuRtEQXO
XWJDNkbc9Tg7SEfLClMxpn9VYiGoOhrxPYj504JcTS+l7aIQ4Rjx8h7ZGuXcLR9a
BR9tfmzHhoj2n3Pqt4cKu5NPlPUbC4vmUKtykNagCXzV9w0twQdiqEXKMurERw8m
otNQRzIAQCpgMubge7NfNdfh0e4ou30hjYQ7g/kp+NSoXrtfg2ya8BbApTRXEeZR
85NLEY4vVwThNJ47Cs8vokDTeK2GzkwS2kffLLH3snMbkpl5AMxs9OgDBriAJ92O
jZi67pt1FyAbuQBrykcnLnHkjjpR4YAi/472Nu2r7WIdpB8h63XFObQTTFXeWmHN
hM4jZ2plxVmUvBqJhLSbna/04k5Q9CkElmYDK9R6V1CKGRyYnm3SaTruRRtGZFUI
IpADYXyLuGxmXtU6qfqdTJ0di1Ox03fM0/b4FgYaG0jczd8JA44u3ChqUbZ3Iyc6
nIc1o4Dw0tAh0CPICGme7zQDc7sXju7cDK+AuCNFuNW3xe/h9H77gsJnin5CVvRG
SIkobntA0uso63il75D90j4Nr1KUvfoOKvNzPMx+e8LUbHgYxdl1yMEDtZorWAXH
DKcIguQMWqIp5pRpS3dT+kP8EcgoaJDBQzFWK4lgsLhahZayjcXEA01YKSiKxSPF
CW2gKFQpw2w4BO7ZwfxHg/5Y/T+Qe96YLCtXeBO3AMNakYT50bzMQupZ3w/aB9SL
2rEbF7R1qVOzkv81GPrCfxYPmvi6CjIjV9qvC3KlW/pjqB2pL3/JR8C1D5pJksef
OdzAKX4fq59Xn3WyE85pkHNQU66kmGJKN6nDsERKcVrFBbX9d70wU3INQpZnQ0LP
LLNt9Za9AysE4fldwU82FnIoX6za7MuqhDSjF0mkfCNgOGwhl/lBtydClY74hxUm
5oropWZDUXOGBhu6Yea+Xd3U2phRIGKOIBbFhKH3ms0JINrCZ39k+zBjxSqTSPNl
YYi6UaEA7XUoeoLvYQo49BLcXj5Pz3wCXqCbOrB/Z0wNs8Duatn5Q9/swk6NBaNE
dgLcKfsDQQSdyHiptNo5vll6kWmk6MCCzW8PFKROkr05SDOs1PGmbL0oWRJ0wrJx
p2A5bCSRBCi4gC15X76zzvvQz+j3Vt9lNinSXEv0UiNWFzZPPdfZrDgEPDY+hKO9
Ox1vDy6wxpiR+hwjbE9WZkrMEK/wD+F65nfQhUJS3T2XYTKa7wK/1RexYL113p/T
j+GIQ9zp0cwo9US2peBMBnachK7/7GenefW/PMmLh1wxaLGaG4uNO0rp7ZqR9iFy
wjnpa1qUm+0+gBEeGbzmpkEPP/vfuLXsu8nUzDbBQdC32SlCfeS5qTCDU40p8cvh
lb+FwnqFghceUqq+lO1A1FpZmg/ZD4LZXBp2wLZY7a3zizuHxSsf2gzhkI54m57u
RH3dFq8sJD2WlqxS0PCQt0oupjsXdrYNngYhO542YUAR2Xv4yKHu1CDn+ccP/5B6
HYtcof2LpbMs6Ro85pmd0OcQQ8KsxL/EE2e5Kmmn4KYD8B9uggCUSBKKWwb6w/vZ
h2woMZshgzXOOHLCVO6F3QzNTvjCHSV3mHifp/3Ks7PF/VhRbqul7UOT5PPnilLf
Jb2Qzy9o2WR4bbufCBUMljRAGocilMpA35+yCtPI9Mrs5lDumGCQvl/Eq7t09AHx
9PvLGJpfue1GlkI+phOW96DnxvtqsvMfAuV724z+l6NJLfE92ijzDFGth+CojViD
S8kfQytqlgjq7Z1mawPfgI1zJo1SuDWG4/pHKnjtbrTZ/BKIz8kG9beNGGiERoNB
6gGSQdMdW2nhMhpxqPDpEjE2Q0gYrjHPmP8IDor3K8o9XIbYjh4D3MqHaqWuqawu
Onxs3pP6es1IXglg8B2Ua5MynKXHMSvMTylhBvK7tkG+MwezX5cykuCg5Ep0eneb
fN60xE0xtZgkh0u4DMo47J9tbKKQ3eretfQyaa/DR04CxLhOm0tsO06j49IGl41q
bCuAgppHBmBZL/+6rUSN8x4qv7JVGnqQOfQnYLo2DDbnyOnWdMZ4ApjuQR/tYQsX
Pt9bz4KTyYANKqCc+dL4xqt4N2UuygH40ErqDGcaVhJgHFTq653TnS1gDytlnx2A
Jd6XvqS/tYjeu45Zx82UAbP/Afn/QBmyfbf/fb0W6D5FKqawHSj+EnuqSts6XZ0f
ddY0gGPK/nqeAOAifh8taeRAT0Ap0DAYa2WrWnuhYaCtVMEtFHVoyCktqDN2vV6+
KcHuaTNWPUIqKIo4tOcIXP5HWe6ZLN/Jj46yLrJeRviQDCwkBsrJILQrZMydBRzw
ptW9dul87JGWppnfh4L7BY7hI5+zTGdJx8SvGj4OzFP/bjZxIm4yCxjBpUZM6hP1
UYQogB91aGofQs86ln29/xApIgOsNtm8DE6rYWRYO3aRMwit+p8ggp/IhkTfF6kj
zokvnZvovdaUPJcnNFht5+SANSDBbP0rrGDMdIP+24cksYinJTP60FR6GULVWKlJ
PV2KSLHvU9mYxZvHF9MAsk4OyyHDxijxipRNygX9thJ2FwDA5sJ+bmydHQDumw5R
nNC9Ts8PiU38wTPH7VU7FBbA+d21NUhlVjHPUo1hxvo1kpo/FfcsSGgqRwHwGjVw
sxWMZRFnVQJZVjC60KWG8x+8rl70dySx8x+M0SlCUUEksHTJ93uZblD8KF2uhp3g
ySGMS6rJeSu7sWUZ/AszNumytL9zPBRV4Ol1D2WysOiGTgkrae6dNURT4DaDfK/0
0jp8ntN/MlYBL+f/GnQIDHqmgK2M5oTBR3+EIAY2DqDTPVUQwou/xmmWG0RBSWbl
MNm07DRLXpzBZL6FtbelB7CqgqxuVW493pt/xa54NGIWVnZpXZgnuBxxF8Kwf2jZ
y/2XFLjot6KpnZC0359X2c8TWKKiffhC0dgnGWXttETsKPSgVKx8E5qOmY4aryzf
ekF+qYLgP+Jm0gFCaee+/M+H3r73wou311+YGFtWRPZTk/yd38sLi/G9r5YSwaou
G5OjvtMbe0OmmJs41xl4spTx7bQ08W9jNwZLMPujDULlVVBg6OS09PXvy21uBzO1
LMSrJpXkBpaFMsTvSdwTZWgQ2kiwLimG6s2uXKLlK4flFB+bT/ttTT/toBKRftoc
V/jHYi8o1pBasqvhgdX9cFtnDUgnNMxAde3/eKSkkuTOvTJW20aUAUTVKDmuFc2j
A0J8/qmriQgbJc5XRytcKyO/3cFAsHnEH0h0g92w+8CvXb675GZVXKjIxhyYA5bc
68zmchsikGUE2i9e2TSbJoCoxpdk+f/Que5gIbavUQAv5rznDOWnCMTXQySmcgwy
POj5/ctxlmBfd9n8Xl02tD3Ypv3OHpDGecwkvzaxR0IM4WfCbsYiJNqECRlg/lTs
Tf3Q4ND7hIDREDRF7p3HcsxbRSEe+DKrvONhJwWSqi/VlHs8g7rRw7O6FX1/75JC
jbMScWUa/uohQEyPywwJ2k8MRUCcLolnxlLd7/N9BJx/koNXqkqDjzKEwQkz2u3/
S4+a6+iS1bo2EIE85ROT0/y57v6Ia6WhY7B1OUKcv1Fq6mTatYRRlWGFqpJ577mu
ugZpGezhndVjlNFQv1tQ/yrDKXKe0KdrUdo8woNU+XjpKXg1Rhdwy0Clf+RXlonH
gpztMlpz8qnRAF8hAxTccHBdRDeoU5fftHdSpIqMEKOM89iXVko2oWH93A7CkW81
GEGyIDddcXSAsaaGzJnVE2PjOpaJULHLgrPhQunqKBUUhXGAku5auGKRAqi6fOTw
8A4JjEqo76A0xgBB4HSCwkzj0UiCgbRCzv7rImsdKoYJJ9P+5Cw615P0C9yE69sW
VNJpF+8Ep6q73C/PqB23mxWaeCCHWQ6MX0O3wmJ+jQaFnr9AVOEcnsrlmwEnS8Kb
ozvRPy+uEVBPq8gKWBv+/Bf6cKCZsEcZBwctYFMz/Xi+gYwyuFayD7ktwMt8dtrc
TH3ZzSBEBtkunE+hc2630lxDgBUdRS9tsqVN8GfCVuDHw1Z8wk+/D+mj4vcpasmv
H9BWvCfel96Rof6rbZdbOcYcXB9rfmlogb6s9E+wpT6fKqsOpCtn5SoY2Vp6/YGo
FemT1sC7zutfo6/hBCFucK58k7y/6Hea9AiWgy/hUSu9MqzvTAhow1J6STGFMVFn
A7a4QXIiMWMAchsLYnTOWhNZePWYtWmrjOCXlWoSGqDMUG5LLgL2/RN4DOEMo110
EJs9qPi8XCR9+0DXWRrr6fArBY/fGo0ed+WXDIVLt+8HdQ9V7kCGK6uYaBAhhzf1
tzVrIfR8Q8yCl9O+xaFcDWbkSyQox3I5INvt34BXUCj+G4RyQj/WWYyHrSBdUMKr
NdK8ef2satOpGm6dmTDASh80Lw93rFFSAvVk9GdAMYCDXLrwsopRlp1kECbzLwGN
tQWoWdWzwX1B5OX/8803kiH+nhXavb9hYUjWkqQyxhMvf9Wi50tQxWJ0Kzmr8f+D
gJg1hbjjsDTpSqF2HtMrDGv9NieN3kPZj6NXDCisyzdcGIxshHFG+KB0Ehyo7oGm
Y0X8a16lgNDzQqoFsZgf/b/fEOEuQnr8L1yQB5K9imk2Vl6jP9XnTpOdMvB+ko/F
gcPGVocnyr3yKgJDbpRgoQR5sY8UOJZ7YUWVdHClzGv+44BmpGeesVW8WUNBrRnc
2FqtttFVIrCIkowIRQClKbTRdjt6X08ylbMIITHjY1gLm8EwBOV6eMHxYsF1VQY2
fgnCtXiUIvuPkN5msfVXMe84RJFxvxvnmG3/wyeT6wXIIQa4wCkmz23IFkjyBeXy
voHRspLVL0MFgKsU47/2ykWJZaeSrxVL2Qz+U/pM7fd9+sz8cS3yU4v4CIZKQxJ6
5q1C1Gqh2otLGpgh2q3yJ1cRCGxgQmGWXd0F+VBLzidBCLNQM3Zi+ZXO5lkuJ+1Q
HN/J4GaHpg+eA+A+p6aMqNQm9s1dRHJYlBXg1OMFagbByY9gXfiaMVgtnd/pxB5S
IxLrPoN2bjiKVf7wtKFF+yOjgx1dTTQJExpVna5R4GaWGCUK+zsXySVmxKP9RYVx
EJGOIwJ3i+NN/q3ueoOzaDRKAo4qvdAlWWEGY0kRDHMOct0yls2lfr4+yDgQ9+m1
DCV9ozs/+ARlTQd7JgQTaI7vHmPG2QGaNOKFOv1N4Tooi7GHEdEmiDCpgLO4z5gX
23XZ59czj23tc1hiySdC3xAgocFk2wmtLSxrbCApifhQqQK1HUlgxfFeJpwJf4z4
oPpd0VXhsqQcY6ahZj3H84CmjHTAbVIJZ1DsX0fcHO249xfY4lkxpQjMtsPcpwCd
GMAMTPkFh/CRD4fICR25VAAsXs02NDHJ0fMtRyTpTGEOEzIcClvaWgY67K38/Lam
5BUleRD/c7kOMbNVWb5HtRTe2IrzsF63xsv61vERi22i+snsm8KKiIj59h9iJTTB
XFbXin6o91Qe1fZprb6QObtSBSVKPTdvo3ED7xbxEy2SIgOO58d81Ar+YB+H4Ega
JmxIDHjqdWlaotcOSTmdOHlcNaxkxLJK8IwCyuK//FIJL4Rf3nyvq61jtrbVMNE5
e2oFNlaNgh5xaoOs5WgjIRdZo+G8hC6aQroJd4PTGHpgkOma8/MWVucmJN7HO7Ws
ceId2Vbvqvb+7w5Xnlh/QxAy/bPaXVVoWEg1YpVnY/NmVthG7igAILlZExOGMGlh
DDFCbC3eeKddQvNSIWoWc8DCc14tVdTDhq0bcRtg6DckRKG5a0cTaa/HGC81rYxi
HrCW/NvH6AfAX6s4MMIBhj6AdOGB6O0Jp/CB17lpc9qIzstateVPun7SVECrSV8m
PXjUIdeg7E1KSaCtfmw0dzV+pshbxgvd8hszVgeI8TzFkDo2/i+0MCJBZyR1I912
zEzhS9vZjcSzyCs4vXbrlutJB6NGUInZFESioBp1Xo87/iTHSIZJ0lA1NABRoG49
SyxHQS+sCNNjdTUln0f5tQmoyv6jqc0yC9JqpRYAYrJ+kS7uFduT+80usUnzEuym
FSTbwJX8Jacy947cvV0dv0Tp0Jcco3S025rEqdsjpyOWax9LYTuqKBO3tP+U6IL1
JMdpxFz57Pwux1RjumOG6UnHTS6n4Zao62YkOnRHYnosPGP/eZx6QvAhCcD0OGtL
3YJWUFYNxrCfmaJI3pMDs2U/xQbRWhnNn3sdPiFIyeZyht2lfCOyZpmU5L3PoISe
rAtY2vQLNrP5MaeFN+N+czYIQInnipGvasfE5/XnqVxCVx4p0RM0iffHnto1XfiU
iIgJ8NENscjFB+kzttv5z0w8D7Spen8wg4yo5V2TGMwSHLs32xOJkJv4aDom/EbW
GCewkcMboIUSegIUfauf8EcPNqyll8l5TF2p5jKL4qeCgN6r8aJvUNfAk7OHHkNn
DZ22u/PDe1zX2JsNFiMxl4VDIa++/LWU1uiAVy4IqHLdvzeH/Vz0adJyhfOKiBZq
R8hcdpTWzVd5o2x6DkCp5bY8j2cKxPSjL0ULxg6+9z30X4kZNaDFrja6b1X8DS7Q
ovR6GMDNbJ2gbXt1Yd6BPQm0cEnbvDTDfxztmDr6/4fBR92NVbWMK1GKgWdGSpdP
ehxf3QwmQDX+Po3nwCTAcFHBjxqhl3tbTr/gpDzcg8KQoy39SfPpo+jlswXsoujN
HPI/v3eGzCJ4fMODMtiNhhGsUslM4QPpylV90dbKeICqH34NVrs35N1Vd8Z0kr1L
xh1O1PDOma6SdkHpwvIJ6cN+O6bgzcuQs6NXp6iCq1BDVv/LF9j8m+MpJ5KYLChP
ecHC8UsgrEXHVu31liLUgwSSHVNmKG4twvGijCTaiCLD5iSeqTcFej3X5KD1ZCHk
B5e6lp0smRu06rh0SYOjbM+QPC3PXKIMejFzt/VuAzcD6i5hK1h7X9QQCWlHWGM4
VnG/egyQhWjnw/LNfiUax7nUdAVnhA7WpioY2CPlK08h8tbk5fcKPV/ssPTOCjAh
9xp8vrfhMZqmkDMYVkVH5RKCsNs4Gmu56dgiWP1pTDUl36qE2zrO4OB4Yzyd+mLE
r+8eettHV47wjzdzJb+CBpyTYdmru7OJNrgb/WSEemrNCiEa3gSbu3A/JUn2cdPu
AQ3N8APnAKXN1TL8LxKw8XyKzFrz0YH0oz2r8zbQ5++gOMjyOuJKA1AF0zI35qTC
SkiyFDMQsAVwhNROUOI6sQ46uZDwko0pmeg0SaEN6Nxxa6PX2mZ/zt51tyKAq1x2
/Ewu80LcolAsARAvge7o9SuUwkTmx1jZvl2UbgqBfLgd8c0r3AwyXnZ5C9lf9e+B
1GyRWw7EK8XoVSuzQTFnBD8aL2QkSZeVKujnmhFI335YIyvE8uzalzQsm/8v8gbZ
rXHDalN7JH7pw+0Z2e1GU0mmSCs6EzT9Sac/+Zx+rlCN2nlFSaSZcqfS9zIBhol5
TJ1DIwmo0egC7z86fUSy4eVMsm3pYSUYP27ew2YIvMbNGKL4cmG/EAX9lQ/N9v6l
cqsOKPUJjIUV/j4XwwOFH405K0jfb5aQ84rLpEMG3xy09pO7j9Id0rufWXIPKLlx
qRxPgbx0XdSTlVxhBpYvt636WIqiNwFMnKLnoyvxgMJcnfdk76VHN5i7nEHYsZJs
g8CZCT9+jANJijUqgrjY2CZNjjf3a1Hz/iHcLHWQdRVKcE1E9KNv0Ytd/egMuKXL
CZaZliLA08VLHDAprXewOac2quc3aSsaGZL103oui73sJMNvVKtyNIFQ1ROIKfLv
kt68fzwY+LJkTxZAyPmlCr1gwpZyZ+60J6es5tzJh5crUeah+4dv0akMiG9DRlp+
kuIE7y0wyNpuUq1jw5q3WxlIkAARnUOSGhMZ0+uRuQ4yAhq86P8cDSniirQdxLdt
+7RD4dooKNrV89asYcCY1unbK/2ggXfWrL54IkWcpAV8ktFfgOwexH38lFXaL/l1
pWo9QNPceemQ8iMuL3zqxC6NVSEqKhJzdw4AndA9ag29YjVQ1S5L/8xDd7FWS0Dz
zZuPDe4rURnPJuptdEuqxghVHEJ8jUjBgdpiPmksqV+88H+ND9PwAn19cAjE9jcQ
De6/TejSnUE4lynpDzm2ZsfHR9ExB5Jef9Aa44PDlUgSmSP9cWgzGla48SXOf5Xt
zCQgaG/znHbKTe+yaaEeLs0kG6DZ5GxmMsKh7tuYcr8C5QhdRPpkoTmNotP8Zf6T
YRCKrWZPDtayL8X1Pz2OrTJya1axsbChyfPsuNW95eFpeBleYTv11jXFAhe1XnaI
lY05FI/fAckHLBOerNajsXUhztEZQGn9S1UeahLB5L6PN4ftDU7VXLYaT5odNmay
Klf51GRQaMNXJj5htKJlPaTCeWaUZbMkRVLm8ZWlxHJCkJexS38wgqYL+A9AgoFo
36K1iuxeVglHybSJMipTZ/TB9pLtwLJOn7ojsPO26UvAVSOBwqQjVAT+zqPkBlNN
dvSU8+qdMog6FrdohaTHnH3Y6gV306oRVkpm+AspQM0WE49tWLMOZi7UQg1JpvQd
7b/KjpsY4JIFtQwirHh00P97yWNNlwh+ZlA2YMNvYXRo6QWIZpTXfjpsxInIdW0e
4KEZTGet+yO/cK34mV8L4LBLPRO3+awnFK1oseIWZoQ8josLR7Mo2myT0tazZxGK
xtbT84JvQuXxodl4MPqBo3HXxAsLeA5g3HrY2mGSaQeOC4H3VXamkzN02BlNH5PL
9OFr8S44piQThj+rU1iOkEzZUPp5MEw73TdcgnETgWG3t1Og1RiLFqQHN0FQehvl
cyIeHZ7GHI5/WhS5jUrk9eMZJvXeUVzXsWL6qXxMTaEFx05SwyhBXwY7eQRYcrdh
O/Z4PJlUjbbKTlwQbMvXjNk1wwXFPo+mc9nBgn2oBFvQmqT5telXG99yc9MXH7yO
3aKcROKQDbRYYNX2PzTgkdrQzDenCqZI4ApEujYuubJh0XQJ/Bmwto1FYkmR0mHe
+GuaYnpeAX2lGqTsRZ3R6qTJkZIdstlgqhIjNTiVcrrYs8kqvL28o5NG9NNMghwE
ZlWSTsppVcG1tgxVJbza1TqHD4Wv0gd1mV9pqMOURX+VgenNxZQmBh8252XbxcF4
PjWO/s3xmui26Jshgul9VZWk6hipJCSmsxLrEE9d0GYUCZlJC2JNr8jxyVfEOR+r
hX9eMyPG7zXOZQLKOhMzdjqolU7KiqDoeya5EDikX8LsWMo/f749MWrbOVAUNjAG
ChJV6ljoKbhJn3Cjlu6fxzKVFfrBVOYa0gCagm5vJndW0whnkhB0T1dVa5m43rbj
ZE+Ld98poF4xS7dpAcz3Y40jvnSXnHvif804NXv38Ot2vCxEBm0YUa5eH6GGh0/g
DIwGEnHEAPBxXzVxpL2uqXz0W4UGRXWbnjoBA8wCTlFOe1XtTwdVekkK2jJwaHNG
oTTYcNeJz0iQMQR/ygFrVXtfs0Oa8//W+lfqyZWK2a099S9MObXuRUpih3QSmMxg
d2PkI+wG6+0pWyGdlqANFugmN5l6rnf2iWhPA8G/mCMsefGPeyhpgt2HArIRFIB2
bmssL9C5ZAWxgwmIKb+9sygj1qp88bf31LUUww26U9pvROSw1UqO4tp+O3+5FWIY
5YO01HFRDVKKBQtSqoYwGw7VHiJJAzbbaStnkcJHQgXPAG+rpiEnahffus0Ov1WO
Zn1U4PUszgkeBz+shM8q1PiYxv1YnBSpak6d59QIJyGmpqpB9G8US9d96xwLEg6i
PxTuooMpqjLNU0DZgw4TEEG0KszNRBLuYjTwJBRTii1E5JZ21lu6Le1U4G0ORYEr
u6YL/THwFFPS6QKKGKRhj/DnOs4tnZcrVGRY89Icqjz8wlmrf7M3Gmcn+IbY4IQH
oVMAxmagu0clztk3MQVaSfik9PNh5Avf5GYqyZ69jugPJlMg3zxfwfgALhNcJES6
RqyWRWwD2wuSFTS45Dhx5E0kckfJCICPKg+RnNwDd42SzbcJG3aF1J/006FdlIbX
360o/JTPA9zv6nlhvhefpwWx2D7egkQRWue6TwrfyUAnAJ3Vjz7mq+tYBb28CsDP
JoHCdV5NOmkpu62tRXRAoYSAcehBjZJrkRopPdkeWajo5thcPeEPirQFHwojB3q0
SpnYs0z+sOGOOPZN+WA241hyzuCmpXz3nS2OmZM1svy0oG3+XaEwC8qscyhE2pBS
sRW2zbvWqxW7xtXarG7050P7mueK8OOs3httSf1CWj7T+Dxqyx3ivBvnu/XtdPT3
woqc5LEMxYoW132tvM/NvMvrbqBEcGKhk69yhCzwVP0kk0HCOI6RpvJF7ZLaNavF
cW4ixFsSZVbJmC9ipWofO4ECSQIp//gXQ7ZdNb4rHLBFHgocPImIUHTNO9I1Eisb
j7Vj119ou6THoNUPGB2daf5jbSFFojZsIL1hNGtrEyE2HhhbTmrEW9H6NwF8ovoA
XAsnp93rUB0Zloq1jUIeEp1oImNLBg3j7K/WkfxuVPP1IVaBjb56p6CstWiKuN0K
jZZC2ZgDBEGL/6NV4l8AKkAvoeK6Fl4DCkKJuPyJYO+3KScrR90REaF11iTHfHwJ
Re6MI4NHJ6mz1RHL/tW3gn/YotRe2UH0go0QHj3bRy2iR5PzqcZChwUedX94fdVM
CmMaSXNyntpTffX54PKbJPvwyMZaLoMQIZh/qdzyt/KHVYfiQwsowIsQrsZUuKAj
mMFwaOw55BFCcwEolQiDh1ibkOusnIMyt+L+3gnjmWTE+LFmyeRCH8kanXS3nO/3
v+z9FsFsnWFbtSnpB+lQ5Rlv3zm7+JsD0gHVP/VhUZRVEGrIhIk6i491A7kC5A6Z
L/rogExSokz4tgAb47B9EWF+LqNSJT8nCoHz8tjFuEcSIa2zOdcqSQcLHxGHF8SA
QxK8Hav26QOy1dyLlj9QYqge6xnfF3Fq2cX1CXcy8YOHJ0yvr3JUserKloBgx/6S
8mPn7ZEyJoleFAEciD+lb4ZJ+46SIzZdUsEMCZGRBUZtpo9ofpr3P+5odE3loATs
4T9IrT2y77KP/SM5aM1fza1Hj4lDIZ4UNwOagmyaj8Bg2ky4m5NQLOldIQfWbbJq
Znr3rF0u+VMXJxaU/RcKYTxGfNATjExWVfqgi+9gCtYvjH4jWVnxPKx2UUT6Chj+
v/1wSk0Tz1EdZpHe2BXEUIUQh6FtcKDW4smtZ59QTYaM9oXizzKooMxCIxQ4yPma
PgM8hzgAz5I9c2NphtsPRc8cYW0jXy456oHTKDxtgHdoJyT3VtKng7/xu3SBqZzm
jb0y3/+ywGy3Yi7sONrPW2fq8K1i4lygazMUQTvQtrpH8Ojl0zQWcVT6QR9k8GDZ
D4IDQBev07CEeWtQ+aMJN3vcnSiPBgnkPOk9JNTqETZ6iQHrI0ZyfV2wUpJPuCvN
3o5Ns4gi2oCXfsHUbUXGpI3VHpxsQqTf68TdSfvYZ9FWSiuxFXdgYdXttwnMOyML
RVtU3yXZ5dbCvEE8wNgKLbuQ0NPInuGMGcwitCaQ3r9ug64GKt16QSe4/mdLlB02
qhlhXaYNx97Caa130zPZAS5crbX9M+9OrI552atoYocYYE5I1cQ7qmiB7mMCa1yw
szI4HlgUmWw6QeqjSFaL6FtCZ0LxWpcO2V1p/1pnziedURkC7k7QxvPtjIft8Dvc
cMk0qr1kTdJaAvUFUgsnPSzJ5dTjxf53bzDysf14Cm0V8l34YH4HfxXzWRyyFDV7
lFNmDKc9fsmOT92Xyx3yjACpc2ztURRri/OGqk1KgnO/KErh8HLlNYCEunel7EgG
20FF2jSrAMUk8Z74uxj5ZCGxU5wp3N23MfpSUizHh4aUAiJLMin754VlhTJoE01z
KxML8C2DZQC8s+EAbrokUr1/n4ilDXXXMENEi5o+5USwn1WVDokSURH9gSsIkuVc
vMJXc3jkQJiGbI5tCR31CveLxC3jvp/d74T1AI8AWhWeoE9rDo9PtKAnloosJwNN
kg/Kn2OamDDj/nmsN3nNJTL7I1UBCMlG6aIrNRDKqwvzfGesvbe4qy4eaQI1BQHt
wHnZK83W0BhXmC7tZsRu8K0TXpDfD11ojUj0XIqJSpd4Zv0tEoXr8FQPODt6fgkI
Oi2j9C/iyEKoZHfPB/zwzTP3c2JFoZPVTPItwiv7zU+hjFLDd/pfQKHPkdzkj3TB
/6vAz+K8+cCZgLDsz3flMwxc4M1aN/w2mdWMfbEfiiT+xABTWmqjQ2EI90gQe9aH
dQyNIS3tfdP27GsR6WsH1CFg4tieDuofL6jPYapEoYcUZsHkeRzGcvv+Eve/JKAI
XBAJydfhW40YAsb0fJbzqavNBFWZbfBlC68Ew29gV5mTeVmc2yroZ5ftPz6SUDIY
Lk1UWLQjz/CHIBXrKB+DSU9IyJ4g0jAxjtCnZeWnN/vxHBtYrKvAGu9fJ0kHE1qX
hwqY7mqMR08BoEYQvzTuMjmqKvqaS5M+QVncjIJ/YysdNDnIYaWlSrp9h+Nqp17B
JWSXOlZcw28DmfU66rM0GCteRjJa6DZDu9kXD4jCeBHzORZvLm61fGyD4F77xJri
9GOM+q1Dx/9UYOvbCzF6n3RfEjoja9arDN6oxZxHMRVjHxicsE3dGwL4XgB4ETHE
jaT7eXp7A1YXwKcFSnPDX8xB7Ur+58sdjqRyr/shH7n45rTnbpedyoNn3aPu6Vr4
Xr5RqZP3ICjLms9rYVubWRzkwbw+LFdZT+3iqF00jqnjzLapK3L+On5kst3zZvsu
xD3Ug7Dml/akpnbj0hxzchETk4fyy1RWGknhM03Giku/bSRRNnjEus4cXNPH13VZ
j/28XPBML0dV2ShjNNLCRWXGWrjR8TfbOLQU3ltZ92MVdcDGir6DMiD1KNvZ0zTX
O1tqg+3Gzn8bUi2M3PIiXiROvfTQXoJ0hCXNosvE4HGShoROJFIHOeUAMF8akpXR
Or2zFLLZwwh9LlM40k0LIS7jKAWa6JA7MPD71FfUOzOObyP/ZMYBndkO7BG8topA
ABgYqVV4Qwse9xwNw47GYfOQZ0Qe+mYSw+QTeU4u/z94PDaArvA5lmZCe5KLhHVW
u0h0G+7GguFaMhdRWo9karkw+26sGhqNlLkagfPasaaH97f34zAj+WBCcVYCMa6W
ftRpNBWpI/ItwJTo8PzjJpJSOeWXsUzFp6lPYy+x5jBiJIftMhmr/7c+QUVm3Yca
+UrdpaThhBVQOFIQFaN0379dNiYDw8WiApGDVZxXqWeariO1x6lNe/2RlbSsH8if
JGa4VhUP5hajrJJt58GiOKE8TuQ36/dj4Hrs4jistj7K7rv9EdSMpHHh+YIYv2HR
wlm8H7L3aPiXQa2bX8untHVmmPlc+KRYUXM/ew9UHr5xE7HYJOs8Qt8Cjj/+2NEO
TPg7o6Q7qfdYEVmpNxGTcYi8t/M0uhm1O1F7DeBv2q9J10QM42YQTfMBlkX0FJ0T
ihTH4YNAmjczwZkasP4l7l3WhelbsmJtXk1RiRQ9VWSEHETS9fr7pf28tLP0N6VP
Y6GAU9OLnaOW3GZ7A+zUETf0zoypfAffvAxy+mGLt2o7YtK1P75I/FnWdkl0AvlZ
eSi1vVjlg6UTHLJic4bwC4utZsO7zONnNDS5qWzs+0f0VQUWU0F3Ht27xqSOKip9
m+c42lRFL1mnzxDwP6fSrKlA0bABg0A9TgS2FKGHQX0jAQjZ3Il+5GY82zUi8zrY
HURQJIfqQ6Donfp2lkOiKAKP0eOF1Mg3Ni5gg9UL0m+Tfh11RfG5h8euPa8cXZtS
Ie06SaNxr5X1I1sCNoQP11QR+2AwLORlPuGdNb3WXLvIh+UDQMNfL1zvSKf1BEiU
0rlDkxoLT66RUtqxRcVM41KFwggzLaqcHgtk5mJ+2jzDWX/HFVVqZLwfLMkJiKEF
CCzIHHbpc9g98wRcCPKvROKYR12zg8T1KtYDaapalsMVh3pcoaUw2NpsfoROF+UZ
iP9cz2r8H6TgS6cQfMav2e3tyM3a4dMyO9GBDljlKwxkVqC+IZAGCQHfIOwcWhzP
kb/g+qcF0kGh1/KJa0StDkf3cwseHNLLFfb790UuSFsrJ5HX9vT837mvUdXXG6gX
2FksHqFPvnH9pcZWbV3WMrOcvS++/haA8vCFq+6gpzrmcC5+pSB8kJXK0dMuKnNI
2iOOOLmACprhcdBt83dm0RszM003K3Hh4l/XeJXUzMpxnZelIz3pq7zSUebSD7Hb
ooriAi7hY9IUL97M16MzmkMyl/RIsAoLjj1TAsSw70OpD3i30TOopvAQToyn2u3M
/cg92RG/8xatFwtTwY9NpY3lqdX8BDyaVoHGr8tEom23BjU1DdJRgywQshLpSrhs
8G4zQeNVVK/v9TqDhyEq2N+xlJD8jHRoynbb6dTojZoZlQCGXtGixb7QlxwpccFg
iQnUFccvPREWGR2Tkki2/F40LqchY1t9nTpNhOj6t7NGw6GDTeG9W8vY8W/YZT4/
fKQF7rvqCJzGDuTWGe5Y1f+tIFxhR92WBfNpblclIqKSzBI8KNYbQtOEjeQI8Aeb
n0/OLo0BYrwuXfh8/lq1bbks8zvcXt/0b34O14QsIzTyoreas8hFDn8bS2BEA4rh
HOOpe2S5X2NLAGVO26xHJR9vEfBY24HMHMjoh7LwwowzHA6EcV3l1Um4U5qIH9h+
GnHMwJlSozLoyFBXKpoZMlcBDI8oyOknKlg/hPiOleVbqLQ8dVKJdz8HGp/OMZvQ
s33fYvwdJWoG4d1ZrbpszSH7okHyjxo6JSYTdklKQlz0nfs5VDzjbKr/gH4RtmCQ
OriF2tR0qA7GGwK57YcuWGdAWx9MAfjgs3gMoGkiSn3z6IlwD245z7f6cRUid7Cm
0wON1Ay5ebi/1Xtylh8BlmRxPLweUThIUBmXtvaiCxywJXvf5XZBmYEGCk6G2GWK
kLbx+ZAOdTd3KnJc7ftsWhPczNwYTj1V1f6RU2tQGiSL8rLGTGoMY+ele1ow97gv
rkJuoGCCTPg+HkZogD6yZ3VLzE1UMjpYUIhR0y/IGqFd465Vv2lnqgtPmT8h8Z8A
nnAM2XtLghHGGPjiqaxeB7iB+GhVckUBLG79y1RlElMPocPwMZpkXGt98Mkd/ymL
zH5jVUAMBbfSdtALp3ffPZY4K87LuDEGqejrxT6HZXy23ETLHr6nuW3Px1aX2yEE
GVuR+zh6h9Lga/XbnyVT/Kr4uSkSehTkfDQbJRQX49VsgbqAoDvp7BmxmNaMyJJO
lE+TZDz5u4SmlrXz+8ujD0kkNY08pdS/7hWXi7rjPfl40gEtltHcXuCPfxLXzygk
crmse01RCEb5L57E/l4uchT/iR6ChYdQpTJ20Dpb5S83musruuYDjxu9ww1fyevt
QwDojqPkFNmxlhYa/UsUI/JbY9ied0cRUuAcgEvGBvrpYDjGVbXAndw5zXsDfw+A
0sU5K3BOq66vGF576w17r4/lyj1HHgVwIKtls6mggsJUJd2g6XHgEOLK++nDtQy2
2gjHvMiwdDODiktekawz8e+uJQlYssW+o3td76BXn/lOxzS9frhyo/XmsSPPArhW
oi5ITNAPIuUe/6GS5DhnT5Uq1l9E9yEPssj5cLCTTwjVnaz0F0ZHYwQMeJHAnVJc
yVDd+sDLJR5iGpy0tvBiaUwhZytGkqJWERGNjGSsDHn1H5RASCbqmiO+RJex1Qhu
vYbgBwzBARMcaEkkdKGU/4eC2Lgy/TsgnH6RL41dMiDh9cgrTBtMHGolnExUvEBB
5/GW+ETum2Gg/xZl9SX/7yb548B4FI1SBOF9UEdAnnaqUFFkdUdQc3MuDLssYTjn
Eibm5yQVl7ERCkpqKL7DyIOAYcw8Bo3hdIMfeYhlrGKgy0NLRbhx3czmZ8DDa25x
lC4wTCKJYGHUyXHsPhZ5TZCwSDiLYeiXRUjAcn9hWUlTFOoeuOJQuVG5SH9gmYcs
l2tz75CZ2ii2QSXHWpW3vLQeAhsLMntMDP+q3lSW3NFSq8uTjDOqNrl+uSDg5lnw
ltwWqrX9CR90E73NTP4L21xJvwa8RgBKQ81MP95O62HqV37W0d+Tp8TwfPjMJAVn
+aSek6haWKp7TW8TAsyvWOJXEszdBojrVMu2oSdQqZStCfwoY1ZGLFQ4LrIkBBJC
FFhrF3GZttoY8dDiTMHQIszrsOBZEbx1t2RDXi+P6XbUjJM78a1/HLC0GlfFtB+q
m43bhmSsuYFYGRD7tVBPjkw9d1e7MZzE2b3juwr46/k+VQmLMMWv2IFJs5lcMdOp
Hy5IWN6cHc3OPfdr5QreOVgw48C9PxTv8KOH3PTCmwqyziCoSUkbaapzcE66cDzG
kQV5rxSSeG9LYDHHpN5TGBprQS/meNNB2VDhBSDHRdNwdgVUDH1r3Qq3d+xkB7sW
bd4CpqZjoMNUteK26Vwd1fipF3KdXK5K++75SPgeJVSggT7hUBtyH9p/YOV//h4d
762yO9qvqvBH0memByct2h2d4MjVJH+Hc5qNAy2ZBHvsrRwAIZ5NPF7yKRKZUBdw
8NCCnmw4AHj4oXQSoEWG2citkA9y50kDB2N38sk6AwpkYQ+C7rxtixSoJ12VtlnD
jsawLh+fC7rup+NppaFBpjMu8BB/aFEjQ9lSS+oj+lY5tno69M7iaNzJ3kRCvCPK
GlADOi2V1KVl+Tr0li0K0XOLky/aTo5Gmma+4uNVhgwql/RZ//0ATQGcUs91EvQy
yUVsRAeF7flWSWtyyN5zKAz4D0CmkREGxC9j3q1z68xbCfDLLBZyhUABm8zp+pEf
jk7szfBl6uTkfc/dmp0IhM63hmK5TgkTWnZ0VKGa6nWGcqnxe7+w8rZ/ZwCMndtG
VuJWIerCGJ1s5rTTfSNY61IfeJrzvJn3t4dPNR6Govyj9/407t2FE+1bojZTe9wM
0dgAHL1uYP3oNCXfFa/NI7DnARxzm+V9a+PHKAWBRCdyjfQHJUEJKrYeiAPm1Y7Q
BbaduBDSQojk9tsD6x0AImoqLcJ5k2zFxSXAwHC1fAUKX/A/C9NB3T6Ugo8nqvIm
AXouHdxTpBiuDcgwuZXRZcGVRGVOlrogDzQHAYEE14svkBcHNeg3PRxoR632oKNG
9wRMNt6qmwn/GrUob4WgN6HVk3RfKrwmTbFq9rP9/kRxvoU8a3v4Pc0JVsmhqMuX
kgFqhL1vkCwN8PXo/gxQTMIQG+lL/tlIeKCJXvdlVX11dXEFDfUaNNWkKnpcPvMO
g7LG9rhpYG2p6m1ovfQRaXSHmfH2HNfHbH5c3ZU7M2EPBhn1xSbP5xxbdOpgmUlC
SmWkRifmTztO8HFEsvs8SIRvMCx8JxWHJhnqdPpGZwj3Kv5zS9atYhe49wB25AQO
4tLJY1tshe1rgfVlS7crR8fIQp5bF1mLyn0YrPRafy3Zcl64QKmJPB6NQKMwcphW
sueysCDF7bJKpltxqfLeLbyYgGjssXS+FTtB8ftg4p0Uz7AlGtFtnWgutF7gmtq3
upkJ8EgCuivGEHaos+9oO6h/Ee6aREJddrOVfKEDtdhR2nzfj5AGunNL9dsM/4Cb
AGpMvi8J0LnNeSDYALcOPNlPwikieHHGWtL1BTM4/SwnwP7cx/qxbDoqphNoL1wp
m1Q7RDnWrtImx4B0HWMLyL6L0BLYc5iDkor0AOpkKOjCus+HxmjvwHAW2y+1mScH
/sB+UC+a2u3UKaj3AGawWDACmgmJolc8NW7FXbZmMShSAWlzmRBaJADbt+si7cf/
affWD8yQLErDtwhmZDfOuB99ad/YCJMxKn+XK0zuQsIsZefVaLQl1dqTqywHGaZL
xp2vyO1ZvmbaccWm/JIkRODJroVG6n6FN9e9fYde+mRoOlCehhRkHVQUkj1JYIqI
qRN5Mx2eU7sIwWZ3d+6TwYKrcdWURbEF9ZtkcjbMxQPGRa6eRdWVl05Ylmh5DB0U
vJGRBwzFpyOdyCO5sjTxWtaXNWv53ys+EMPwdpF8c2hibZ7R0Bc4yiqcvrdqYzFv
gVNKhSvEhTiO/y2aD8+AhQQT5p/3LXEpch6MSxllBBMcWGwhqT5yqjuw6Q5WY8/j
Z5bhTtaPcfpUemOAbwM0Yvqzlmfq4LyuoKH02pgZTc1b8yoF8JyOkQM6XO46Jwur
tWQXaN7CMENBwjc/3N4TOMhely4HviB3KCAVWsQ+/z+jFw11+21B03r3+p+1kEHu
yhp+sj7PSNQ7dsQjK1IhPUuh4Bl8Kbu14ncs+zvt6wxoFFu7yHUnqMqdhfD/YZI4
pHigD/BGUPGzogT/c/6leCLw9u2mBcWTrX5pZfcFtNnfd3EdvJH0iTdpxIQAcVij
mIrDbDNoQ2A2iPYyMvSQ1D2W1AP5+3VpFQtKs6Wsq8GMKYufvoSOZq5PRVlSg3YS
+F8UoQuCDAzSXJI7IvIM7ygpC5z2Jb7uv+/e4EK8rrDSgqJS2bVmoYtpu7ea/D+C
M4wzoUSReYhhwqwmwhE5sQLUECHOvLjKsuoELb2KELMnm7C/7qCx41FE9jpXs3MN
w6FtccYiSlIvdqMgv2JybI43u/Mfnk05Yyvw/IVeNaJwzZoNLLFgFCGmle8JuuiC
daL2R/AOJbPIcHu0tl3yhlpoyu0qI5Vcn+4BbFagAl2S7d5pEjqBDs1QDD6w1IIr
3+LlidVUuMVtNmlMH1Hw8UXsc+2lm6HmoO4c8/lM3TrQtecFPV8puoXQuecZKYHw
yVuSA2VhcAqA+kXsCI7OzIioZxdMDF7/nw9k8hJAvHTSWuI486N2gECQlp+9Mmys
59H9tBK3SemWZZBNDvOZuQqBZLnoOU8MsfmNNLY63afBc9Nsd8XlgKM3ILfNKwia
KIZNGD1lwx13TiaALTPvk55XX7JhdLdfmJbqkpZXuihcqXCw7Ff0xAQxR0tUBlFg
+r7D7jy30pEzwwgUO62FcQyTGQAZA33gFvoCmmchs5Uk2V1XW/eM0lwxUxgI+3IB
oMrdnp+nHiauDo5R0/7yFsdVJmPTfEJrJ4LmN/cu5cenahg4xd2God7V1nSnAGTK
e0FU7uy1dh5ZJv+BFcRr1DvW2MPGL1awAt5dmK2cWYfq1Zx+fcihRaTFfQmsjLca
aBsEcIpssP0KmlTKkeVdHZB4mtLdvwanr8Tf2JLey4pdB4oC2hqmfafkfWXoaSAe
F9q5ZwTSYLaWDqYZov27EoXN3dPbCmon4NZWWGlctoFD7ZSYDqYdMLE+LbnQhZh9
xfaUuaokukQsEaWkw2QjjPXZbcyBq3+Umr4y4k31u1W2cKSOF+qlkSwFDkPVMGmJ
HsE56s1vbj2U1XzY897w0nor3CT67wHSnX5JDHPttkCJuLgXp4JhFO87dqwNmCAU
HfC6JgJLoX36tJJfK0QBvtdkibyAcygBzHIiDUOrearor8H/nAO6usnKb/Dqk/sr
A0KIHLZw4l4y1Cwf5q2zWJWlTsc+kPK8yfg8tqi8nq4razT/dDNXlkePy+f+PYcM
1ZW0Z7+ir0O/OOfsijdm5J0oqYdBCU/GPEhdV9/tQ5J4+MUOZ0mKvcnb3lhe2V3j
Iy3TCoIMjwmMhzI2omEpOEQubv1PpNBxe6GvSOmr7xELj6AR8yV2+rRbE4hWIbkR
T2wRim6SDP7B+5T8MMPPYBI6bnaj6Q60551MCWEsZlEcIhSpuU0mBnrLqnYMqv/m
yrNysmXQt/AKPzhU/pNfjU1KcUM8lJNsRd7xghHBFzVubN1Xa03NMHwpsxdevC3r
s78i5K1gVQ+6FVAE9jh+7z5CuzZP4YZG26gGo7gRXFfhpbfCSC8c3fhALXe7HIH6
hAqhfnMKpeLV6bvUU5m3FiZFNB2e7gQMssYxLcXX9+niibfDexP+L2DDD8/c53X8
irWhmGVCMOlMeh8giqFp4D24X6GvWxyt5wOT+I/GU+fzr5e6aklxBmHiBIcupEuN
ImN6629aBOq67lLJvRJ09TUFuEIhZri9x7IYzjb3j1mE9XNnyYstve/PWBcwLAkT
/2x21cHCgkOqrOuzHXU13zKJlhxBwCCUMYzq3PxwcVJVqGB+3fvpRkfDiFRhBr1t
ei6oUQUkIOGcDFkBRDnKZDVT1gQeiA5nOYF2SBQCOINm6ABKPyANCgaoobAduTr5
BJOQh0Z+EudbIkdcCcfKa6yoMobi5qET1w9oL9UxmxepZqnObNXpzs6Iw+E0zd+r
4GC7pTG3Nw6gl3EpRTrxXM6jEqouR0UPBDvsC+hCtqvvqL5XALzXl5rxocBEegVh
wOcqe12kuTuFQX8RwY18BgtQz075ORDlwtS9LjJDPSkd7SJ2mfLyLh3x34KrtL0m
bZCczjX2JgF32hD/Db5nzGiZxTiOdrJFwwDod3cxzV4eaF304ShDC10vNoN49nz6
otFxqhCayraRpJncjeuK5uL9jYyDe9Et4gjrGCG70JnsI79yNuJwMr2p3x0G0/yw
s7KoUP4L/u3K05wcjYuHTDQXuH6Y7yHz1+3LffJXmir8d9l0OlHfe+uQksfJ+PzT
tJ72HpQEExc1bse/Ndq95O1hzCzbS3cygrM2v69pvcbNNgoPQG4Mfzopaq0aGOVH
2eg8DUnD712ZLgrWDw+srIB3CTDtERrXl6liilOeoBTW+h7pKlmVM+GYcgGtHflt
SFMp1uNRMP2Kx2+GtehsNHMQcU/BdJQhYp901roRl/yNJtfpbjfYLfaT78P1JpLm
25DKLJQ+fvbvBruA+Q6ri1xbW6wgkUJPLyEsUUsATp51ADNHJmzxgaOUTy6KVwCW
dth8whC60dFPfuaTXrLocDZWTbNlKdSreL4kuKCzCyKi1rPda9k4e8VwQq5UCvYR
nfRJgEHWqjOwVCWXwNJQtnZOYM9MpbYnSsAFSfIpdb2qY60PNtX4ZUh3D3OJIyKl
xnUQeZtsQlAbzGVf3llHE+7SvZDNsHkrzRvwvHcd1RQgu85YxWHCrrT3moSdbU8z
jZ+XurVtqqHf6W6kJ0JveUod7K3917eWeYv25rML3uJA1eLUIhfT6RXjJ9u5vyUc
REvtC4+p9V3v1iPQANd4GCe2ujmalPTblXbsp3tv5RUfsoRgvUMimslDBe2J4+9r
vq0KiyNUTCjK507RvB0wxcyYBP8eSg+x3wxp/Rw9BhC8llewvAPFYilBAdjKvdb8
VgOZoTbtAEV3oKaGA/1wFoRrXDspBj+jFCDnPhx6/3IuBuziffws8QFmERWuWi6U
P42zcGQkRrcFah5i4jY5U2l/UbMJKf1dn8UjOXvyKfjc3dKoyiGQkHiwQtoECjnl
Tn1Df+FjpqpVoDtjig4vk15JIJSO5yys7lt3sKryp3GcT/9ehmy1O//sMEu3ktM1
PJVcBUO/FBcAaTsbSTrsreyoxhDSgOgFbjAuJBSYSFH3q0MaenweW9yRU9EAFHLP
TbEfTqOREIYmqgINMexwHYU41TmgVzztaAYr+3UeBIaggX89twMsHgAXGBGEqJFy
7JNdgYl0YpVhOIpiqntV5VnrufXlAs2a26tbJ6VOsbVmKzqFZ+eaT2/nG+z/9EJ1
ryQ6Nvq6v63OpF+aTJkLokAkwqW8pYmh1be+ZJEaPNbxBhJgZw1CnayinJwFN6Ii
J3ESbq8XdVuZ30iz/LO+wx3XTYB8iWZIRaC4WDomqJsGEbllPl80aTQLYGF/9uAK
IN43kYkK4Uhea5xkT9uKQDgt+km8iMqYGt91X3Hti0wv7BiOoC7Fq9iD52pblevc
W8SUFhK0E5tvKF4FmYlkpKZVpB4RenVehFSJ3kRZeqzmrp+Wn+yqWwUKq9h+aLAz
uKy/UxizcV8BJX+viXQeezO7L0ICtWcYVMNNqUuLx0Z2/mNbf1LWcnuxCpCJsQb2
5R+uHZrmCUX07iMGxkx7/Zfu/31/n7JO1WpYw+1SWnQQEN9OEGC8MuN3hiQuRwpr
xQirAExPuJ+p1BlfnN472Rwsc7kONLD1KFp8yqIAzbKYAyJxNTQTyMnyBPvKMfa/
C15zVtTqv9KAITxXLtQcHcarnjuPZSlDrIxwfKx6KGQzxmHLfFvUa2AbKl/bgQSL
1nTDoLFbtD+MAK5vODEa1msYY6M19ED3aR9UO1J/wW8vzGWuFQjpOS/9YVZ04+h5
l9MgFL4cUhGl+Sr2yob+LrtWE+0pAhhkfgRll6V9f4jNq8zRKJohzJX9ZJIm28v/
VSaqQlj5F5Bh3sO3gJJvSHui4nFLAlK+p76+xonJN9AVqNoiX/8PX2U+DkOm1SIp
GI0OeRjvUcaE8twqBGMsiNFD6wmT5DBsV5D9FUNhVmQq59FchWsjsta2so8f81dF
JjnWLfv6alAAIOGDvOPwDyN423tot56WZmCHigP9WC/3RwCqEJtpeVhCWSPc0rjO
QCTQdla+MMvXX8YDphJmVap8Jl7GTIh1FlcmuKQ2Sy4KQ9QGnEDCks/NtgrBOfqK
r7BXb9sGdl4l/tMyUBwEw2W1KW3SiX1pZ+1aNercCIGHnPHNSj2k4nb9+W+1r9ll
rnlZhcvxaxeo2MU7pTKoqwF97Vvq+jLy25Gty7Ipdsk5kXQ/sdcnwTKwOwdf3HHU
xZnq5crXEg9Ycf9wz89PRA+R+o/EdklQ44/TfvPh+lK5VcquroHuFnU+FSXDrcQN
KBizBynkBAd3jF09J0bT0OjulST6mL5/aepu3a8PDAI3pgEXKOn7n4rQPQgP3VRC
le+GmsOVr/reXQxJqOcOvfqpEKqrNzKAMSMZgPHsorE7cQVSNQ69b70YYJh7uyWG
SCFVA2Bq047iWpVhvvCUcouMexJklPJN6idne+aCWpDeWKcg7LYGoe3BTmk74RGT
Cx3q6j5eFvT/onqg2+GN64wmTGEcO+LUofNeFu1TO5UFVfs7XmqfZNpue9s07YCx
3pz2luYlVBF0naeRq9rJIXlrjViSxQo90LrrkLNjM7WAvJOwWCIx+UUdbwpM1B8o
dDnhX8+4kNNtzB1iQ3O+fJvP5E/heOabqoGpIA4iehlfrfE1G9NVrUZ6VjcmtZ8C
r/6CuG9r4w37gORgttxPxwuZH2I6K92kn29gc6YwRzrGLlDLj79Pr/KkaJZPi7Ks
Luv/2uPXfmF3fRPHveaHxu8a4XPCBDlGcQUh+J9NfRwncIXF+kaIEj60VGHsukv+
+dTmg5tChQsnj/0r0W8mYFpP4WhUaD9nuSkfv/uuJuUlidvr63lDpI8J1tPZ5nUh
s5TPnimPzFR4Uk2gV8VtHzj94Nl0XRgqpYlxW19IDM5rQb0iQAb4fe+UpmePTct/
jxu13DWaUGgPBYa4QeIvJbyLwPPFExz+G7hQ1ZyvRPTFt3FRDZ7OKRU6dETcqADY
CUQDd2gfnuH/a/t7o/48DdR8a7LriZdZ3HWYjzYy4BIe+wHIHA0LLCMY7s4j1AWS
VYXN5EanethrzARFJ+ys17Wg0QQJ4BFdaeGZp8nkk3Zw7MLMRBLAHTiCLyF3KNwD
mVmS7ApcQaJQc6YFt63PnfNMh3fJ3/Y6Ezn9BWp057l2oCVP4T+UhhS0YldFBgyJ
Ni1e5GMoi/RD7Fdo0TFuW/l+bQ91s8t+JlYKny7gW8gvDBCiwnTkvRSo5FjV3VJ0
KO4ujRB0toJBkun5prs48eCgv8nV2tWFjiYVAc1AjqflxBFkOSYwjv+nx3pX58Ae
Kn/AJxSPWwyrm3KpRTpE4+9D5uxdfkJvDizCbDrY98mX/cwXeSqVi0F333ozQndF
XM21F+Zwfu1+jZWNJZkyvddoJ7jKNbg/SBhU6TuBCq4zFj5G2KZ+qLziSibgcOi+
jYOs6WBeGAlup3/3tBtsWIm0ZM2cGg/xsY/6dbSTmNtBxWAKrsO7lfTSh/c4HKjG
27tfiO/BMUF2mPiaxc2svGFzZEAUKEjhG4KBsJ1aCOyn7iP5qixSjzDEpqxJDt7Z
2RwS8+MC0Vf6RHYYSdK0kYyz7vUl80ubo/mbXi9xf7ElCATpucR5guiVQIZ+OMWq
1f88fZju1ldF4Am4z/kSd7VMXqMoh4+DWbgI4MKXc2wDzEaqlgl0tTk8qK7pT458
HhC6iZIgJlZqQf6C1E4FcmockFOufd4gylnxevtJ09Wgv4urDBTBok48kKtz872c
ygXMmuYfNNb2dUqvWwfuc4f8bNDumj9dvJTNoFZmo6XVh/mqM2GljksB8Oc6MDX3
+fdS0tI7CYv80Cal9zhKM5V3lddZELAnpwr2UBdb3yGf68zW1NjDFDIB3jkixhtB
v8qUOCAmqQeD1XT2hiD7e3G5Xaq9oal7R5cQgDVW02SK9SEgt1thPC7exaTFSK68
g94VQ0dUX175/BDW3FXYBtGBDiKSZLx5fwQB45yRfuNgYyF5iZvQJXsIhvz1IyTF
0xNK8jBtHtS4GfOa6shWd1KZpjQBuCIEsxtz9aTnXxwF9qUk84HqnhUnMIIdyz7c
L+Zs2Yq4ZLj/za9Ku0wFG2MSagEGLms7lesuOcA00MnvNdjGWmFCoys1V5VFYsr/
sMJp16V/UhekoJvit3b4poXHdbReLxLZ6hSZaj86L7YrvAujRXPWK943D6CjSaVY
PHKHop2PVU4K0id5HfQPNOfww5+L0UfRf+/DVDbGm8fJalzTMIrP7qYvOUM5PM8V
5RTUPI6dyeefOL2QjBsyDH5YIC4zj+coUj2580xImIWpVslVfvxMJdiq1KM6kKya
zoSPgQugbJXcBJjp4F+tMLv21qzf0VBi6SmsqAJfTW98NGvb4qJ4KoAx8X79s3Ug
ofZ1zoS7BQAaxcY0PcKL6/fjgzsG/ZSVkO7UbfY1JNzlpUq1gcSgp2llc3NRgg2+
QNK8XMBdw2d95UgU7ptI8T8vCk8vwPrTCqtu9Atiyprmy2KkvL/fSReeOPc8EDw8
TJtokqte5QTVT3TW5O6igcr2LUAVrdAGRF1MtO0nkzaiXziGQCIXeulr0ao0+ICM
G9OtXZuGVywwr9E/SouWBqNNHXs3SbZllmqHokEaqdNWm/FKPTyJnZ95SCfJkfN9
1+IPWgzMAtseMPKsZX0rUFxj931c1Z+F7HSGJmGeFw4oRNXStldtbadeoZ/p8KLu
IJs3EOL3rpIpXgZyGTpG3GfNFlNPlriALm7bu/RVBWRQvJ0ZfB+Deua+LdMyt+Jd
k/BiuAfnXwVSjcmj3F8Mn7MMDdP3HWv6PQt26h0LBPj+uZmsMKjr1FQvgvrBZW2V
sBohypGquWTVqTcSnzLQ4TiK6DLeBs60DSccvXMmflO5Nt6QSoI46Au/ujME0/pJ
3kwhyyfp0lyLfKav882PgAvMT1wEEhUsJeMUQEOm/CagEQmDddvoEMzsaLUVla1p
SGCcjU2aHrNsKCdHtygereCiGngmJYtJUVizaUB2PJjfLBWZq4qYnH3HHu7FoWAu
HXNw5cTZiFE2NWwthsvHyhatO+Ocu2Hrn/iM+CCyrqUy+f+pFdxX9O7J+pjjodU5
4FA+SjC8XPwdHNXmyLQ/Cg2Or1cXFfOw0qtBDBTlsQVMYx4W39K2JqkLQr9mlF20
K+KCZ5A7xXE6cCnAXXSoFQOnzX+KQW+yAgVaogz+MUZlpihRAC5LIPd32nlqicuw
VaHR6LwYFcE7SwchiNz/NWVHtkqTjZcy/X9sGnfAZk36yI6Azf6znZWIREiXLElD
nPARtC4a+J61llODYUoj05AeXeSfXFmXcT36w8DJog+bP9CAVQyrwzK2UKKvLhdb
tuOFeLfH5mVRr/PEpUwmGhye1ghu85CGxoQjnRGtCPFlG8BDpslSKzMnMBD6EaiI
S0xdzFoSuOoDGBIo5+RSACOoHO7A3cW7SHqe+sge7l9XDWPE0VVLVZfJbRALinj0
vhOxHzHzL2QbivqWhi9zR+vAaofuXH1LG0fOox1NCz1wahIhJTdt3lFUS2g7iD+n
zoVzCJFsHCvOsYMazgmjZ0SB5UBQJSJNSb/h1oNBuhkWwR5PFWgO6XYUpl10ppjs
k1PHpS8O2N1cVxyAi+Lns8hH/WkCwvLgDnTeLKXYGPoDe46GGhxx031NBfll9ZDf
aoTrOLjzWOPLZBygNvSztr3A9gi+0vU8jP3ae4voikLO8cYPOH58Tc+X/XKf48nK
Q658X2NWz/3hikQPTj5rCOvmsS5JPonYpWFLQ9uBI9lM/m0Q4uyNdMtZzHnsHHFM
jFShZ3NzCE7ui0SycwK/o4BgDCHgXSgbDI8VUXoE0GUnrF1K57XMdQ1ZZCS1+H2K
7/Z5sMdu35+B4FROKyBbANoREeCKlMB4VL+iqaS4BR98/Lmn29/FGE1exCF7PW3f
I8Uv7FZ9FjWCMJ9uUH9tzLTg+UDKAw4fJZbJ3ZGRwLa8JKmUM+p/UBsvrS1RqU8j
ewdX9HNyefTghCqiFXT2EuKIMs5xui6qy4BEUq90Mh3wNWbjZF8FYYKbWxZZbdMP
WxSwCt/a2izqJ0RrL2RPKK0JgbrTaNuJcWFKL/9UbH7+w+b6H9NL7dS+uHWhhAvv
Pp5/0nhronQTFlYS6IzWHdQlzb4dpawtGs6fN591l983kOOaW+adHphS3H2Cr29/
XLbGDENyEl14cZBZmJFT49ed0svJPiXxE6gkZUNHp4i912XS4p8tBwamfsh++ZL+
Y7pU+U81EYSnIFI1bpuBmp+o8IuPgP7TQvZ5emHfg1yvDpp1HLZh/B5MFgxiXpYl
ZVs7EKDLfCkQlYmAnRw7sRSJO6k7/2gMn4OTp282LVi+LAc+vGIL1aqDdR5j+Dg/
ivn2ui946S6DkW0WGMgWLZK9Ixc6M2gjzr/NSCoZdgKo/Q48v6DWjzT7IGZ8HM+H
dOHqDzZvpmlNElBspnje3+yDgdrraz8Ozhf/F2ENzXo237+b2CZhZ3ue7oXTyGn/
zeBtP2zF7UMRjVA80YLrHLn+KEiH2KZQ4m/0K4bkVQ+xMAKlT7PpYxEgBXpMauHO
jTNBBfz30dz5kI6iJq3ZLniWIrW0Gq9GT5qrhcKskthr9ReE0BYBcIB7gUR5GlC3
PPAnMsDPaHXdbH9kCpFYbrHEexH4lUKjWSkfrPfbplLBueh5RMl2i0WHf3Ps0vaN
pm1d6k5FZGfoS9xowudMi7pgPVdpTbGx5LVMV5ZrfOovnRjYMJcFLgQBmVpyLYsm
kXeRcn6Cl/tQtlrqd/rq56LWgxP7sgWMgR42rsV2GvI1xTqiSToHqBsSqG7tr6bN
IuiGdlPELkLWldoQd4N9wWo0gXkGsuFT9WwMqMWEOSfqJ+aPdaSG7Rr2tR5cc4zr
D0g0JTj0bQ3swN1nrpESm7KxJrMwpu8ZuwVtkCeOc9kzqRJlPicTKZUU6fg0cqUa
FDyDR/vCJheQGyg8N7ZJ+q4QrjEdf8M4caNcLh+tZpfg3Ha/vVuDcRGZ7Tke08DA
j5pT89BefORu16jinlwuPi6Qnhys0PxhKPevgNNOitgZBAiQY2MNeNTdPQwYnRiT
m7ubMyIsw5SIf7S6kFZ215skZlcgVNC/P/xMS/jP0FPS9RUM/SJQmjUTrMKR62QZ
ZNFrfCuuawxUx3Zrl59xDxDbPVKz9ibsRsmo7HERh2oFyeTEmTbvTnXffpr/znG/
ijlbznxtcfj3Sr4gW50qule5xDsZ0g1HnTWNHMNvr4IOFkt1oZLX/lpuppN5LMhr
qZlDNLlRpnSjrUsdOoS8/0GOIO95QLm0N1I40Qf+v/TINOJjygR3NPtpApf6/X2R
MZ7u0G0MBOSep+Cv1LrmlXDdSdX+tvIWTORVJvq+ZdMJsAXPPVu4Z+0uQlWwdXOf
lz9Yki9keoj3hi4QDLBnsRsbbe/Vh8EMRAwJSuBog78HDQkDpw3/VljX/KG6lZLj
FDJaKCRBNU4XmrvPK/CQmyVJjgzYl0F7GmvHRAKj5SSc7ToWxAaIUj65+QDZvk76
aUmgR2p42Z01ZveppvOeZNqh/MqMU3NaDCHzdVXDh0U/YHxkFm/u5cAxOuG2+xfb
n46Dw9Z+eSXyYucGSpSAUsW6DHQcqkdeakOnET3g4AjmAYPmQ7p8jr/GMmMzHmkm
4j+Fx+GmmKDGnJ2kWZrU+01swYluzwM85vBtLV5sMqxaMNDbeoFPoGR72jx24MwD
3yzFVI+r9oDqNexagVDlb8UVhW7B0mxFY/7IU5VEUmvlbaXCyeKxvnsSnIuPj1vq
bXZJZ0hIWG+UnI7e0aF1H9EpzleFYwkphtdl39ViLhGTgsCpyKfwAHZxkTO6cuaw
U4WjXw5u0H6IqEhMTQAdRJy7XsObTDX3aVVVUYszP3+upSgiBe3USGr3ph9q4mhr
wdrxpK67/i64MucGsVjMlET08ZsOj2XZR8Ssp3bx1x3wQkR8upH5Vn2DDvec9DQV
/5yWjCuitygauU8DQXi2sucmToBOyUsSWwtbbSGIBT7G+iDVoGdC858eMlJkFb22
SXbcpPXrmJ+GTqaEhdSfZXzu9EuAR4NdX0eNgH9qSWTyifZfm1kQ5VyXBe2elJzG
bzGBZjKfqnTAnMtkBgtbVKtLf/GFSd9tyuwSSStvwAdimtDEpJtj6BJNVde1FGJb
esx0MV60gAC/zFK0R+y9qvMT/TwPJnXbEUgYHHZhPqQaA+SYRdLlHA7Keu4LSN94
d3jS+eHL3NsN6GYI+MK/yOaGV0A7EuM1rAW18Qpn2rfbsxfzht9hIRTaghDLbB1U
IAmLgKY9b8qmnsjh325LCB0yMtOmxYK3CD6ZeqrD/0tT/z7id88yhpYTgwIZEOny
5yLEDhO0FdAkPMM7mAh6jSzj3zmdoRBHQuCktsJ+sGBHx06mdjaByJt+B9JwkF+5
vBWUxxEcmXWnQsItEAr/KSuZznMqssfRr2C4kcQB2YyfMSwhgGpaRf9qo4BvCXBi
QQDihyjfIEgKup5KvK2kg/iMoDU1HCTWkFG1obAcaXopjt88RvvDY4/UIqOIEsOI
Ls5azgRIBYsUl3P7YkUH559YDz3Tnfkvd6MF+/ASOS8fz5wGtLxR1Ov27pGrTjYV
am4JBnjXdLbdJWgCWf4ETtwVpD6BeP2fCwhCcniZ6fYepKpx/SjTKdJQsguUcbqf
uEU5K/ST3chmcfrKLOZSb37V5uJpwlxyIlSMvt1VCGjHAJzeYhnstB66ZpWgXccZ
XyPrq8j1jW5//8zM543rmkBtmzr7yU8gCNQ/eGXhMak2dDtu9A0hvAXGNWMTZEzo
Wftg9ZxhTWEb/yrV9o3rGV8QqcInNFE8pRU4IqD3DWM/7WXW07ifEcux/U+MzysO
MwbZMnwfPu8NCUipODLTvjAAjhuUdBqVdn1Rst+nVN8Y+FnTue6izASsx2LiRLzk
/iO7/0lP0YCthFillrFboEnMeFs8FkmxWLYWXbd/NBNPu8Zk3vuCgA5l9PDMh+R2
FvTMzkNmbUoEhdyO3sZBNZ65Q3PJzRkL1gGvRHvfUxtR6bY3LpgXT0/DL2m7sEnr
C8eukXKCE3V7nCgxclAtG2bPZBzpdpNXURMUBkAWKHXiK7w3jSLOh+ERoM6YF27D
xrA3/vZymG9UwcLnz+Api67TJmVUwGsZTTeUMmrtq7EOzhYOxsJwhZbTmj4jlGgg
qM8wn+bGLi5JmKfqkEIsKJgctWcTrVUlxBYuRuJxdf7xk3ADnmCJtm8UjUVd4djC
/94T3pQybqu3Epeuc7R+KpTqekEus+JAUPDf7QvJAeOdL6KqHoS+VBKN2W947X91
yJbBUhOGF4+bHSINacuYSOSg3Qn6fA/PuUmCfdvzhEF8gYhYqvmGbe8q8M5afSsf
9iyDIChK63UMJMgGK9/0QlD9N2kgjQ8eZVar8FIdTdMtDUQd7NI4RH9M8B8ba1wS
42GV1kdP7K/vaKAMeeIb2I3fy5pT14ES32s3C/evTiBU2Rufsqnq2QTMTBKQ4ZZr
6PRHwAI3jXUMiIkWt89jzRcWsS3Sr04aK0McUZE7fbmUJkS54JgkljNW88hU9EFN
Z5XQptdbReTt0KgIdpVT5NSgx8TxotF8SlENYdXVuOFdT1GkB/YEw5IeVzTn2gH4
VI0wufKrWnxb8dYrle5kt/DizXZ3WgTP7yrN3DarnLVEayy7YZIFfIc0HwJKMgaB
bOyM8hcTrje1ZcEMxlPYkU5R3AA2YnWkeR8tiMeuxtyx2Eu9F9oQudeu0+wQE435
xGq8S7pDH+2G6j9GhZ7btDQHq1Xf3jO6pgvDQCOe48pX6G2x7xbktPqhHaUEleqc
398O42zaeSkegh+Bn7nch+cqAaZMdwZ5LE80JQPs75g3aOOC+SwF/CMtXK5mGHvn
UxLVfeVyXQBKq8HMjyhn1yVofCZaG7TTo+/W20jPdonUGoHWAeDKw1P2FKORtzDC
NHP5Yrmw5QCaUQifgVEr9sL2JV0CtJYLF7Yu3OF4WEoUsIJtZeJk8Pn571UyXHG8
gw3zzP61LfUXL8tRbds4/eQbMis88xACXr0NHDpHLBfd/dL+5JswtQyySnW8m/jl
zRdAwemc20an00c28akgVJxiIHX4ZibSPwWugPrsUnBmKEZG9EKtRiiGMCC/o4bx
uvUmEBfYUOYW87jUWNh84ea0VUasHLbfyE9jteWq8fXm1fTH+KMpeeksyKanApiR
0Ux7cdMVCJPHyc9bqLiKEqe9WVmX0mAxK/YEhTxm3PBU7pG057d2SQW4j7pyRNcM
uvVwIQuWwqOquOtOa/vE8Dky2SOq9eaptqRCIysXiBRk60n7ZDS9vhkVkfgXpBTS
pZKVViizqJQKbBJ2JYh9vaM18HNAmC6+zH20lA8m8PmJJnr4h1fBFN71OB5B/8rR
eyZ6Ec6Ps7uG6OF2fnopRX941QFerJ8L58QPTrlhAMcKDlYZHIMil3ImcBrUIgtl
NZ+Rng6P6Nd1j8CHegmGqvO+SkGKEOQkfwSgHiHi8V1jVd6DvZNZmxG7kzng1+pw
jSDed827Tm1ArLeg6evzItsJ98Bm9ejuH1tgSB1Ix2+DIOy9dj/A0jArYLNd3xAC
JdDqVXyhS3SOYZH72r/XldJUUED8czotYR4Ieqc8jGiVKpCBPJWGB4kK3AxlloW3
fbpjbXPYIArDVLCxIXDs+ssiAuKil79mCz3THpUDOGqH/A4LmrpC3NNdrx6gPOXJ
14wlHm13X0hFXygPWwTahrFaYxaPoDh3zRKsIt/MupSvxhNm3kSHSKfddYm2kSbW
IPeEH2hRcH7eRnfRn5OH6iUEPZAnkEzh1Kle29lUMYDXFxrRBoycfMhlErwvqFiV
DgdELtNVqhn//FfXggjNwGL2Zb5UW35/6OALC2YsWK2A92sNQot8pq3o+l8IU9j6
4cRE6YT2WIzuXufm+l2It/5gTxSHaBo+aSN8Hbeye2Fzpj532Otwd/keLGjsJeFQ
Qi/cY/HPjOLBSxLB517OvPeroRL3FWBExqL3bp6S7aAeciDB54y+9ZsK3o/2SH2f
DP+GVg9vfj33JYpi4By+IkoXgdpz8bhfcUs2jEu1Ms4wPJrBjnMx7rhonFWltgVw
YL+4D/d31JCbkZwhWUoqDfMV06nvSKpRuBk6rTxWp8BlE8uTW+FlpAdb7iZpCKFO
e+RqrdpxIGabOKA0Uc/IM2wN2ZBslkeznZ5A3s7+AuK5Z0Ht+OlxuXwmLivxeQca
FJ0sFulD3SBHIyk3/92GrkV3Ufw47SpHweNAoCo28xkC+dSN1SNu54ZkBxm+TEg7
J6kt4SSXlQF/QokrY+5MK+MJVlq/5d3ey9EL2KrfZ0ddes9epej33BInI3ovXXJo
T9k4TXKNEn0s9Ng9fY8tvWrU/fa0L+gU6x4AcjwE4bfECri+PM2UxRUb3ukfC63a
c0g5SD3jN9Ic/cE0zckc4azOjz2W9RnUQGoE8QwbH8fEcnlEkmH29ZDIHunRj0HX
jNs0EAbm4yR+E6RpCk8lkFBuolXJgF+XIf+JFZ7ZQhf0g9/2oSIvL/52EmJq8TRM
HfGoqu9JjAazRkvgkJC+3mS6ck33Blf1JsymC4vxVhjrOHbZNJhC7PIIWLni57Yw
9rHEZugKGSxB9xTPgjdN+X4OoYz7oFm0umJRbuHq6nnOVq9g+YU3eTqI0saGjD3M
e+gyfo2++Y9osQqz4qrx5y7g8Pci1F1VxJEajKQtik+nciKIM9gArX/XcF3gf35L
v1qo+66hyb8R04kSqtyU+spGZSMvn3p+EB31P4k9+49s5CDSEk+bT/DySrbHEC5G
zAM7lys22BrX29QANo1nfmLTArt7SNCqLXs/FImXCcnDZwkhzZdZY6SYricyKcfM
Q2kTSyboKlaP+9FMg0rFv9NStGviVhS0FHfdwl/D7LzzJWG0ow8sPUZVbeaO6RUd
EmCA8Fc7pmzyjcdrCevohisE4OEHYD6xBl2hzUApjrUfbuUbaJ3pFcvK2f54vEQY
/9trZJZ4/LwZq8tC20MORwwOLAZYXmda4zYTZ352/dl/Q7SGfuvwIeTj4vY4X6/1
yPzC6q3BAfPfrUKkRBi0zUqOtPcOnnc70U4n0eFGhN/8XpIaWJUR7FQPS89UuH1m
EU7PC3rgeXYpq5pBB0Pg2pf6/Bpo7JGS0tJdSrUUHvaH49kMBt5PENjEPqmXgl9X
GV3gejhNGWv6K4g6lv0mpUixwOrKW+Z6196ekhSBv3d8ILlDEJLItfHhtSb02rfx
r1fTrrXQubaZOSA8nE99/tRwYBbM9X8WfepI43HCr3Qv+H2C38X3KbystTW/32wC
jTlkn/8d6ff4pKo/eaue5j1FxQqQY7xMcr5qbu3J70PR19GSLYFDRYHxFDwqvc6L
g6eAc+PZdKPIfVUl1GCZWg2cnPH27dC4peJ4HCEENcHVig3pGC8a2S5Z+9GX0rwh
NlV2BRfnh1+xAj16+3gj8lufFY/hRPhqBG5OtAee2CCG5w9fLqUxT9C02FnOlpcs
GNVHRjRtIDUyVp12otozbcx0QW0UYVbb9GExr+TlYmvy1PI04eBwIUG0g07UdKIS
mAnFqgAEu9XBFnP9i4XNufmQq7sbayzQetkISSGZNEbchUb86UE0jnjIPZSmMJMa
pD8p2JzADxf7RRtI9kwbZOMP7zRA8sFSXyPuKdmdSDeb7tf5N1/IUBAT3vlH89gM
n3hgGR0d+33g5jLXhLf1iqEMCTC10vl/DXfMYiQ1QMqWKhu+FrWpDyKLyFD+IBm4
PG6dYde2EI5q4a/ixZ4m8IyGNDbmheJdru/6Gg3h5zEL8iUTeIVxWA0ROU3oe5ZM
s8heTyCXV/KqsPmw5hG10YA/crsd6tV7opPIlxjWp8oIJRjB6sKtHlOxkefmGnUl
jHpZeHksXIrNUhbXBO+gnTMt5+ZmY2/y+EVr5YI6nOPE8NgDU++JRD4OgKMOcSjs
tMRUul7VK8SPUMVhLhF0caa/0fueaQi1r7euabY4cJlqm/zN+oh/eg3Sq2LTpmJg
n1rElFPIjUtM8huZ0nZYyPapx25hX1pcU5A0Wnsdwp/AgvfhOR7Wu1wkc3qJgDTc
8FUBCB7ijOgoOuubkW2rZWpk73gic7iQkF4cdTapxH9UHUOxvygWYGcuWA9Orxmo
AUYcKQvg/jhBFo3+wDloD0hcThyXWqYpcOO06Zrpm7pvBNTztoHVc32ThPimxxjQ
zZiVNlr3pmLeJn9SzeZ0ijnNfCgesl/kJvTy0Fx/ReW0dli0vqK6uz7PkyClLbwD
DKgzrVU8IVoNnV6/gEiPqRydrt1AIvuG/AKPmov4959zdhllmNTUdR7OvSd7XZv4
vhWb/4MKoZOKLnToCJhfO25XdafvksqoQvhJts0+phrAbrkwL8A1sQM84Y2vHcl3
jhMLIr+8AZew8x3/OucCrNDQ3xlgeh5nEWXKcQWJ7bhoFxiJW12KMU2vMV6vmR5w
hsKvx9roE/VHgPh4+rLralVie1vwqf0222rxrFXfgIVdlE2aualFcewEEAPAfmMV
XxZ+EHYa/9e/jA4EE2e48yY1dtMoVzv7Kg/SQdYGgm89dZnDavR91zP0kfCLvjT+
j4Pnxcd6lZEEU4j33uaF1g66Deq1WwgvqiTMNHnU4QUpsrpU4CLjx7LWDIMzAbay
ozBj7zZ3PBVLrSZLirKFoYYnyqd+r7+eVXu4l4zPhQvXxaw4VGjLXzf+30FtLYjN
RjfCCH9Iyd/owDTfs53LtN3xKIH1DtJa6SVdz0yQSmPzgGYyYNOyostUDNdROy0c
XfEriibzkbCFucA01h4RuXrrIVvP4d8MgryuSMv8zYlgnAkvCesn/LY287Ma1e/6
+nnaPhcaRxlbV0Isr5tbnUxrAN1pXpjVSoOjujQmoxz9DWpyVT7OzYAvqQxk+YrK
KbC1HRMCQM4bdRisyGZ3gjzPAaTOud40X3V4zxklleo4OwazvCF6Vg4c4/AGEAGI
VoD7m6ta2liQxHNZjOUr7wyZ0ebpoyVSMUzf7wPZmGyTRcXM9bsbyJ9fUFEcJW0+
t1i3mdZYIqZZ64h7aYFn1d7unX9a32f2TkSUOSze3FjmSJSWp9oIWKUfAqApD4Fk
dKb77qefhO9LU9tO8I6TFla/R/xBtKBa6IKDsz3nJUdvA8hTOSRkMT2q1mEM0pxX
DCdEXlAzimPDovxMG/hQotILmFAMnjB3LG/cOpbn3e2q5f47prr1bjDiHiqV3AOV
ZvLf/I1GOpVmOhNky4c2rmw3UPlIshqNknNJ2KcAYt7qBgzrxWf0qGj5dDXy29vt
xORXhSeVxhv+h17/Rq72Nkr4NfCr/MHzgsWS7MWB7tgtZLK3FA5Iy38vWfFC1YnT
n4+N373MBBuYDkuHWM1NPwqrPZbVsoGAL/C6NSTMfBRjQq0w4WsDJjzI+6p4+1HE
tX+bf7DIwYSVGch3bKK4QjqbjJosVgobwRuwRiVj2iw5grXR9BWs6cW1evQLPuHk
kV/xhutnLZbDiUccur+B3V9Tmq74+z9KrxKq6cwrmoPi/hzAf8z8knI+sdtmvL54
3SdBw/oSVVSZcjsCoG9BHEA08pS9Upzw2rQIBrT8JbpMHuaPf04om/skMUJt+O6e
bqlu9ESVnrbyzPNjCdXLlDz/ooeEH2f2gzF0VFkfqOzhSlgzDMlqOtAa/VRGEutQ
MI9AaaiZKQrBG+czHkAbSYYI0jIOBc0p1Y+1SSAZ/GNgGw3AhWZ35hf7x6KUzhpZ
v4KZbTsigZjRJh8KAxO6hoTYo4JkpZFrtXC7a8IIv/fUgngx9ITexouXiwT8UqVj
4/xGsFb8gdWQoy7l4KNnTeP73l6bHPUwiaq9/PdVx3bprJ1r1EJj+UsPKVqCidDA
FgrkMNoO5Sx/jFOl4Unem7B2pMs8IkcCIKgcxNu6R/nupIM4w4M+Doq8gmwUDVto
4C76P82JKMTWYwLi8ttwRk2kpQFdpbV3KmCFy3e0XuYZu9M5wKQp7LCWzSwLTQyJ
Psju9CnsXpLK9QNJerAsdJ7RDT88UuLeXIvhxSNA1h2xAn4vY3Q8zc3a+MryhtRg
SQ55Da0aDfx4IEGMpVdKAspmsYK9WrjrqP/JeAC/2oBVQa5DEsEJCxD/OwqqtSxU
ic4C3uUHGeTI641uWqPgD2pzOW5kcJHD4INpBWswyDAPzXM4xB69wlEucZDkJKgM
z8r0eggFaCoDLuU4Etan17m7S2I3HWmsYyQ2fGTyTkjFgZvGCOjXB8XP9b8H/Ih1
zbGdwmSGPhW6Rnh6ZA2EHFs9Kanjf4kM78Ff8Om6CbPRtcKTDKfi4KQlFWjoLOPQ
qr0vOg5JretrzDB2x6q2HM9YlMmXKonHSDWAAfQ3pYzESwId+XiujGfzloHlp+co
YBGiKnWyOJex7mnCsoMWcP2phc/95y+6rCrMw3e/3tarJdqlAG8VUzbrFnxginoM
P6+HBcGRNAgCzGmTI4z/9PBSOet/UDUVQXwKKyjvpN/6VeTlEcVHTlkfKEuZ6X/k
tHeDi+q8R3wVDAtsyfEkKWB8DV5si/waS5XGyRgcuMq1y8A3GRDW2OUCpVsCnDK3
Pri6UL8fFdGL/K5zpH3CkuEvFggxcugrBwkKRZa2oi37DA78j+18QgtEgCR5yWpQ
AIhFOHV7vd4gUMm1sJ9BBAX8Uv3zQJYzK34d1F2Z65nPV2HYL/sYXrdbiI3RwCUE
3FwUYVlX/R3SonZS6AE143ra/YOQkCgkyMOe0oFMF3vr4Nmqyqp2FJJtEiSzfP7c
NHQxEHx/idm6BgIWQtQq/EA2PYrwiWc+S97U38X9STn3XYLPYdkj13rZDehZZBKo
e+1dEnuS0jZJgNC4ngpsA3hWvMhuTL3k4hRfxL4XTzTrPIycELwcPAG1kdo3OD3y
aBJU5D9THLcyLE3J87yYgV4vXq6z4fBap6fAOxFdztxFsN3BAyHwMDW9RENRI4IO
OmBumUOE3lG38SiLMf24JNT49dueHpXp89ayWSO9oTQXZhghWnmrBGqUBmISc0NY
UC/m+KafcYIdGkb5mmTVioHjzvGBMhUFJWQtyi2aemLqvokDANXQ/xxgU7MZFroo
47nd5A2I+XjvbRoQPEkUupc1AYACrgV6KjvFUjTOaDmKS39fXTpNcYgQNW//eOwr
/isSf6arpzu9hXV30lCino7pSRUQCrzpDng6G6bOUhi9XD9Uri5cNPVbkxPW+2c6
G33szRRg8lFxBULRkpUoeW/SLTCvU4IQgflEsyYi0nrpXdoIRqgcB5BHpjjcjYeq
sgxg8DDI4UBghDEV3TnVgYIZw0KtZwIzdTG/Kp1rhqdOqH6v5zQ2uUz+ZYyK/NJ0
rcmuzG49lh+xk3yezINF+PcUHpchcu9a21tt/Nv+/54kaILKA666FYALUNODMah1
wgldVwyygMQKGAk6ssY5/lZUZUvcmVS1cnHR/5G5EG9+hHw9viVMV4Dkaj3hGANa
OJuvqCPvdx41OTPWhuRZh7odAiYTB09DANIvj/v4/FwJZg+TxxRM3s9QFVYMzf3I
ehoLM3Pt7uGPEnc5j072Mg8b8tlkkuw0f8eNMGcVQCusmtbVtH8q1u/xbNnnSDvG
ovkh9WJQ8g3U11Vc46KSRTWwvriMCbTw2xn1F95XRDu8ghQUzKkSa1Eb+YzFfRH4
3nH2FH/vD9j42WgCVG+G8Qz8Wtqfq3N08LHqRpeZWvFvfxgHZGAwvQPy3Gy8xeW0
SdeyxcTHxR23Db3Dh2zdNr+dTjj/kcoAYqo74CTqRsKV60jnihspDh33Im0ReYvC
3oyzThoUUdrnEsszwgGmxN7PpgNdDkfNNc+2LyYKMhmm+MbZj3PgamOhRueCb6QR
/dywUaULPXIzozgmGDcw0IMnUwIg9Z6InIIK6X/llKDfBs0n4+LaK3gTxscgs013
TDRrVV45TKTuoeS6/Eyn7x50e4JQ6eR2djd6djeZS4KsdJ322nHylTBLCIUQP4Jd
gpDgYuBfxY5cdSvpkDRp4FpNEsWXdvVyCsdHib2+dehuypXVnywfSOYsnFhuMnZR
bDNvIcPjWl9GrZFXM8APx3KdQ7j5cxOiIhCmxH3xwa65lZCH5C3lmCjLOpX3Ah7V
/2Wi8xc/Vhbr8Rj919bEzcZ2hcrFeplpanbIQoPNo2BmNb6rwEEuKOT9SZ27sxTO
GuqOgZvvrlKyYbDCihRn5LAoJAolKZritnxYObq7IuI10CCpJxDC3XvY5qj1sboP
uJrJFy3/x53vX11irTDOVWccpeCJRxtC43V7BmRDrJkTGo+2N/VU4G3BxwpbpNLJ
TwUxFnT+omjbMrbTwZX+YZ62pV4bcNmkONakxuwyzg1G2J1YqIU36b1crqNhobbI
REi8/hzXDzJtfIDhZsv4RMwY+WLwFG9EapYgOA1nVVGTSb7T3cxxh7uUh5i/QKkG
yr53+CWNLvsUAY+CvsPBjUyHKfsSG546NdoICXVnYm/DLO8AyzgIrrMxKeU5m1Gy
tNFMNV4TlbBrFxQ4x97KQx7HU9jlYvkhphGWjL3vTpup57v5YEFt6HcM1D/yILJu
utBmf4IlFr71GUhBPdk94lwDpNVfUu9A+myidaKsvAuHeoiv/LNoVvIdW2w7Yngc
pgdaZTbvAb16uFSbrnR7cA3GSxRwJmuYZpW2JAyyieR6wwHvxjmQsEq/hfHPMtcp
rLAz0VJ3Sj4Wb42rGapjKgN0vuwx4WEYfR5oE6ZNLIZx9G+ixMwjS2mtiPXPwbYb
bL26MIM16tUUQDyia8oz7j+81bkzSRrRxs4tn9I0s+yF/t4OaRVt/+UKwrq72O2G
J0qiJFxKj3hdjkJ6+fWbfzAnm32qw8UvCo1BFcJ1jvznSWon4BJyuMqHmJ87R65j
lA3iV+sgfhTNLMiZS1JUwk0yA3WbxMg1WnmuIr1gkqav0y2vos0rYzIs2OHIYPZX
9bge0moAfFR9AnyNqG28Eec0e8FLKyosqajXrBEje6yMNfKK12aejowznWMkEUD7
A7gcujXSRs3TZdpO5D1tI/rM3T98kD3Up7CeuXUzNt2Vh6kYu6bKdTDKoU36F+If
JFpMI4aAkH5tni/UzbGsLTzOMSnfVn5e6RO96uCLZRj4B3LS9S9Gq0bhu63RHuWd
3crhJQSG4kVovPk9SiF7XPQxygY6QcL2oC617UmngR+gmEH4sQ3E0NG4mTPqWDnY
dqxHX8i9uqorBl8x8XHs+Y73iJeY+cHOUW6ThwFNJP8+6HXMbR/+XJ8t8PPB8XDT
SK1nqlxyDlwBoPfMMrzNuc77omI+h5dhLXsUjdeplzDzPkXeyT9Lj+qxxIJxCW1P
UN3meUMC8JKkqbJCMEGyhW22QREeLBbBQKi+u8LIDLghujvD5KgogkADlBOSIJ+u
Al+ItwrQVDOV2K/CSpSJSa0b4e31IDSRdHkcXvkk9TyHbr3A2FRqhjTsbRjiguz8
T95jhqW+114nBsK8FX2O6RXBdj2cPuV5jiRdPa0SvAaz791wASvKnb4mgd8UqtE3
31lBkrwZBNvSWeTLugc+E719cO2aVQCwYNrvIydV1DE2N2q4s/5342Y55nkHLx3W
0JUQr6vP7/NfktvbAxPLgmng50sMjj6tf+TsUhWooVlY51b7ik7T+aBbVZSD5ZKx
hH8CJpNn1I5x9/lKlqu/VKawFxK+I7ZP7wsQkjBS79wV+nWULKz8+62VqL0jXZEu
Ndo74qxTAHDjauNj6UcCAeAPGFmitEY9vMJzmOY3Qg2ue2194rKNql7cDiFjfTYz
jHZ2+d7GOSZ2aRwL9wjifuaxWjphJgF3J3ZkQ3/JSDQQmDThAIX5qjWCv6NtqMXH
hDt/Ud9EZstBcoYfbM56Q5Viv7OCB8bD/HethbKvsT+JPu9V9J65ZsZULL/+NZsu
BDrpQ6PaT+naEUJ/OOQzi+Ly1z71U9KiMD/uGmIjAZFkcrr4TQPVbhuygavOouNf
K4OWWWMZLQd4lPLXiNuQpzK+ho9IRYx86FSe+E5Vh+Ebm0S4B6llRxhHCJsTb6R9
w6IBS2qlzLVr+dg49trFAF5VZwi4EsjEmWcKgkDiyTL8SY777Wp2Dt800QbRu0I4
m5Tej0/Dd+b0qCtK74H4P/3CLWLOPgENWmjebK7d9GRGh/WnCxOVqmEHWlp3Kg1g
rfOUrDz2t1t1aaMmvpbYp0KBQRFKcSTxvSviSFI7g0TobpvDlS1DJFbvDZy3CYxT
iqGQiEi/YIB/lYn0Wn1sxw0id50EM2dZzdLCjDQgbOnDwx361Fv3oG8W9VjTBeLW
DgZFrt3D/148fO8p2IGDhmKMaeKhj7xcLD+Cc6EnkIbmFfRdraHEI//PHLYupAz8
rbEaJr6ykPs9WMG+C4U6l4b2EVnbdxq1nD4+nFH2CMR1+iwQTtzK+ttFB9gU6b0K
/kwkKmGWSoSsl5U5dLbRC1fDJXcgx75VMzVUHicF1/VpZbybY0vVJyjRBWJAiWkA
vzoz20tcvjxrq/sbGUYAU4h+FnyuAQUjSyOO4qBNuZIfgneWJdpv82LKlmEbBEWU
a6i0C6IyW1cVwf6NnzvlTp3u20sIkUkkwXDU5RweCs2RcqCmU3VzuDtWWuwaOAiw
ygwyTFXOszdqOqTWjrjwdRDqmPJaM9v60BP6eUpPR1ETI6UgEw7SvWbRM+Vj6Tuf
Ro6S/eMyioPfNodTEswqngp8utQPfuQZ5ZGwPijPOwFHOvDs+Bk5lNU2lVQQT+YP
5mN7M3BEgGmX9UUQXIS8TGHVYWLo83VhITFIx7namqSlQImIYM3tqvkCN/Siyu8k
QP7oimXxuEo2A1K5iFBvyCLQcumYQ6hB2Rm538rxXwnmUSetznnZz0ZD0akoxWqS
QxTUh7TvwRl40/xBwhSRbbWaljEVhlDZxfDQejwG7LuUh5tosfJOhodAsZZ7aDE6
2jxnHUCO3rq9slVRi1QQikFIG1PVVOqqVcuM5eX5LZUu3u/sOgynYlJeG0dLRTs1
zVKj1AJpJfzYOxuO42WX4BEOTC0nICHIPR32RFiYB33tL72QCv++h531MAsRbMer
6Fx7uqeR0R6CO55NsLpnBXQHdP1NUjAkvfKLTDSs4JbZXSccjmj1QqFmsTs79lrx
eIzcyjym1hwRF7l/e4Jr8jRNppE5KRjMKzptKZgx4R3m+TOJLyzMe+zBmKr2NfoH
9B+WZi/3GVl/ce2xpa6NEJMFCl2ppcK2dPXHKASuOV6mVi1k5nm0Z+jhsTHZJG4s
bKBe6ghgW2WoOVe8BgdjxIIdm1vgBp/kknRUH0jVIZF3PhWB60NrbcloCg6GZb8U
v/y8+YFnOnEF0q3YlSTLhdt1YgXkwYeOkYYIvficCe7+x2i8kJpGhWqDZYVNX+jp
cDk+mhiC0cHIPOEeonlJFw0fDgTTGDSCESMJynWF9ZncM7wNN3Ehzvsi2g7sVtRN
HTvP2sHC4wZ5rnv71k42nYEFfLzaLjdJATFBT/9LjPsQRWn3SGxsFgr5Tw53rMW7
42CQswAmlHfvVAQYaOI0vGmSa0Z9zaZzUQZxABklYccH4u8mXowZQf1IrRgtItHH
KSMNAzWJNdbYqU3P2Blt4ma8u2a2/FDnX22lvCU09Ni22JZ3QZc5bIcnR92Xao94
Fv/CjCwSp/4dsTkCdg0v7CJiZo1AdSa92NFSw0C9iORdu2PVIEV9Stos1Z1FvtGd
nRiiDhICok/Z5kPB//qcbFvLayd10uZ4yqYheR5WcEFJXsAlhL0Ls/SIH3Y8DZlT
VzWQTEy8j9BZwJUQZGPkGL+5wGTZRaETO5dzZEGKYfQk0QxjCVTLkelk8No7P9mF
o5SmknTKpJfy+qjlRWNcTf5N7O82B8sZlvZTcq/X0H/0VeMNNhteSYOdvSNTv4HF
Bb1Ba5Ok8W+34v2SKBGVSgb2AsZOMbIlioiNwXH2lc1bqUFceeBnWHsVaaS8vp1R
KeZmu8AihrrvIjQGbX5sFdTXd9Bec5QJxzwCZsfoMCt2Jwlknm/BugOWyzyqG6Yc
mRTWWeJLTnnOa5JvAN2+QQ3/GwAwR0AntBrrAhc7OV6f5FVQq8p7kiASragdUBP2
2TqKGKgbQMNp+wOroryb8SY/BGLbYy7vj8fnnPYWd2AZlvEzdOKlK63AoEe1qaqp
cZq3pylH8mXi/or+xTUB6jm31O9GMtbCCcvCfXtZEYIjOI1HtxZ4dI9PhSBrOse1
jiK2xvuUPOILFyZP7292VPXTCh+2uris55DCob2mxon+TnmStt3RJ398GfKAWG7q
JfvDePdhnCOSupKeNe6SVNy8R3fdb0/0XqQSkveOEuCmi7yrHjxM74oe977wIYdd
hpLRzu1QsE26ujPz1Rn/HbJIC6Eh9UB7mzeVL+RzHwjt/TCCtUAes25dMi1WlDvD
nKNlWjsIWzBwL480KfTCC3boZMN9wt8fj73TsHV8jqrQ8WsI/TdfEt1Q+xvAt4Lb
mANlD5YFcQXE9COF5LpsB8D1orf18qyisvSdEfeWGEH10rYjzfr8H3sNkr8PBXd1
1fsvFupoVL9Zu5c53o58hIdseJh5FQ86koL889pfBqhpM5nIljwy5ocHEhAgNKCv
BXKkUn6cJNx/I/fvA4zHU9IxfnthQkbeT5Qu7iP9p7C/8MrrncTPRBisDTuA5cvm
od52KcOje7nZFLekBH053AqlzrlJ4Monz3mOYD+TwbhUCuNbsh2naJZq5XM5X4NP
ncD+qjr2zPiVsE1QnnXhc+sp4yIZ35l/7aob1qUlS37PRZxn31uazQdAqLe5tSf2
J5kJg0EMTq+d3M3Ki4pyodJhKlb6oMP8/FaAMGGJSBk2YubwS7YrLXktySfbytVK
x8JyIYuDvQPvG74TnilRmVKiO6zNqHUe8w+/uVoMPX+T6gXeJIAzI/zM6NSQuzrK
9AjHRvlniwPVcE/aPr6YfTi37hMIVVwL7UWFkEaybSDjZje3llZ7jVFTZFzw9bfr
GDButdbKtpvOU/sl7f9vC2LD1r9EefMluP6Aeh1oWTwGZne9qYtzravOVecSFLnS
Tr10LClhxh1wUvlexCj0xl8sXtJIW6j1McvgVM3UaiDZQGqyLghTnseO/j/MM55y
/u2gpvj4P9kO79PhvM6qdJgXGltkMHhpaprNNaimXk2fO757fyz5Vz/fB2qdJHpO
dfeb558UV7Xpu0PsF0rZvfjhskGjpJWiglKdXq/TLBg8NdjdS7PW1dRwmVf5EMDw
K1srfJY2PDxxQPZeJXR0oFakwponlLgxiqHJLvw+FajWaLXbFOcD4w1Q1QGMqHtI
byEwwfFfHSapG++CLIarLImZtXtNnV3lcHQ6QO3SSrPDPacqeoy1o2msdDqRIU8+
Br6URpZmU+NYsQXWxXBK3f0RwXo/ScCTRs4L84RR0M/e9C2jg8RR2HVHmbzVi2Do
2JXisFEl0UM5y5SN7Sf7TN8EoZ5G38Q9ZkJDwZF3Mfp//qQgR9mwfqm/OyPCvKgV
uyVfQYn6w4tMiX3yzh+cPIbW66SwnxegOxOgQm8BwlsZccd4KC7VMiATImRrICqH
RvJg6/4oxAFVDPubhwAeDAZjp7VnhA0OlkcXhM3L+VRnzqb2FgIRbQZqNlfwg0jU
ZUNrHGKjLE27XyBbZgSMr/FSyJjw2THsoRW/WJOSuIEaGikTrhyk7XlCKijTxKch
+7wB95wXma71GmrrOlX6czhJrWXncHAS9+FnDfGcgKr8cofOdLVzJpIuvUaEy8G9
xLq0jIRHoU2VT5h5mHK9bKcaYRnWz3NEy8pKtyzehL95SN88i5Kih4IJY7DqJZXh
NmTeARkrQHN+JZeRt6fzda3SSJzqyE7QQbL2NVXGqOdAuNn/fpqhWsr62zENoMYp
IdFYVEDdFdsjqen2FmW3XGSqb+cSNoV/WAcK/eA1Mzl03ENqN8fysJijNWfaDvLa
xoyYPuTLjwn8n/mukf83ohXflyB/I/e5pncZyWjhh9mZ4GQtq8RlTZo2qQEfiHjG
HFjvZmqt1LDagAdml/qJrTMBsO5UzsKNhZlUmXc8fZJvcbfve2fci+q+E35L1Oqt
wbCtoGINA0ab5LROc7vLKXUqk1OgJzw8qq8zhz3pNeW14/Rg0LEA21jtbqEZKgrR
4SDHoKpbBWGM11N8xdVTINHbS+dzWvD6Txy+/GdRqgSoqL9usBNMVOxByy69Rwir
wM/pMcrv1N5jAajKVIsZxtGvLno5RZ7wIYhdNlqwG8IYWc71Ayp5UNFrBNB6y0v/
d8saTkxM4T57BzoTM/Rnilhw7nFQcOJMmMJspAtSthez5oUsOyWqQiFPENONUWQe
0XWpLOiRDm3yqwzooDswRSVlqSqtuTa+8aZL6FzrmMIeYFxt9OxG9xaaSX60/9sG
sIBzeiNIeL7LghGRBQxaO1ONZoRyIEoM33VTw2kJg83sN6PVfWnNOwqwX9qwanZL
RbY64UJCNntaGAS/aCefXUUaqgLYfaABEOBMMeTRhlkxC/CTtfok3+wncD8f/sV7
qx+egc537pmLi9CzHMVkmj7fFsekj/8W43wYSIr66Y6UKGVO+2NuMiLXeyqDGc4Z
4Ob0MTxotkdxuVyYBIUtLrutYpxvCetCXNEk2klAkngr3IajhEVxQpMUTeMNP/if
NGBgVQ5iV5RWTrfJuhH5EGzLo3zNXOfw2dTImT8ozVlTVRfx1xoi09eEv4jSRAgI
aUOBltD5YOTAHgZNhKrfaT1ZBGCrVE9R4k9cJ+aHh6zC20Tbd4pcV+NMvjtbJyPI
A2dNBz8J6JzEpliDKbkfMFL7XfTSe/o3jgn+xCrDXEpHfF+RebEhy4Ugbb5SWo41
fW5w4qqNtKkmPQx6XdffR9da+TxZr1L+l1vQpn2HMElnin3BdK4+wMKedh/vP/cy
w+RT9mJdyCjOySCji9H5B0MUXsL/K7Hn5UnqhdrktBpbNToN/Mc5YjXFIYbGUcj0
SmZN1raJlIaV1FBUxZEYyd1X9X519gDFRGSbU5hna83rj7yjEHF44zIT/gslMWj9
9Z8wZmj//lgNcKlMGLS6dEowLQUU2dXQgy+QUYu7FKd0ruDCa2O0El9dxA8Z5BUd
JOxEyIUWol5vd+egwCuAZyOy5PrfZq2EiKMZThMiT+88vf2wSvkA7hF4cOFK/cCD
bAJQEc/da1iSjC1aDrG/Z2h0b/JPz4pWWGccb23F0QGfrasfeYhK+wP95wNmJc1k
AE49AJq4ualIz9wPXwsS202nXu+IEthMq08idczxS1F5aCaX4/ZWFkPq8OM++lA0
KF59GzUrv4HbtevMBp7djHBGzPiixsGUUPuCCoxK1Y0i+HMKoLpA2IGCgHezMzNZ
K9fbrNgji4n3aoqhTyPdoR+lXCt0FowuhVq2JJCy84jvUNKrnjksy7UQfA7hc95V
peWA/efgzRI3L+jpnpZsp5fVHE1xmspqZj6KzqMlSTdvygJSBw7HG9jfCn7cOH71
uoyXF3G8TSrcGeoTcgC+77kwl4+02BplY2/+KR4WgCm7yMjOPQmws3SuxeE7NfMv
vEl51WGyDVlNf7qDlgKhkByOakQDmArkAtrsT/fk2DmCKWuyJkfWRZHQQUdN/xaW
dM4ZV8zYbnzPewmGBPdRphFv716NCPDDbXg0woaVWfwLCsDLuPA67wh+u5GMdfP0
l80fbnbfWtqycRMqyYaZ1KdLHvYf37cCAluLmO+F0vSQDMFlZpeP7ncNNxbLozin
A86wup+5uTmf9c/PuSJu524QJco5PeQz1/s5CHZsFls3HEkG9I+csfY8DIQATFdH
4Tz+PVLaYqgpvM5P/q3WeUDgKsRTp0y4Zp0WQusPFHY2F5jwTd6w8x78IzjXqjU2
VtjleYgHJESta3iKSUHPirwmKrtM80VqT1hkjCl9fXL8eLp99lkC/s3eav+up1pz
O/Tmou+ClW0vwJV/aiJ3uht2Yrm4bHOo6YAWkPYZH5OL67AFhkY+b67XbCUZJgjD
2Sy8T4Dae8tS2I4s9vx8QFPpOHter1BB0hqgWOgw3T6zXmWdsM2g6LY9H/YE4z/w
um96471ThNmxce+N1HL969BPNe3ygCRMVie/fN8tSnjdehDsYgD7SvGSAm5IPp5o
xtS3Zrq/UOsar6qne4aIDCcQ8s/Ih7KBnxt08rtP8IbkmpkydsuMtkLWF1iL9BWt
NheKf6lIrrjRueJw/U25Alx7zXOhLW+3XKH2xicuvf0Vib7AP7fyxW5VakDcDXiP
ldLBtTRZF5Y1YhRvS6yM5nJux1sQJDZv80wB+xYgXVofWfKDr+qpnlFQh1UO0/EP
0V2uHrwbQy/h/bUO2gptuaK7HsctG/wqRwZ27sbiaMyrB/ZpGHRYM1GnIb0NErGy
hw2rYf4jVoIcSnH4oCW3W+fcbBiYzGUFjeEC8XBHeGM1EhnT91dYoxsvV56cjvGW
3bHZn004btU+G3KGh8WTesIBqOq+1cvUQh/pzxxeFtTgaE/NTjprbSb/pV36fLaQ
NXQYB9V4G4xfVAfur6KPI/Rs8ySJdJCAifa/+7T62JPnMreJyMjg+7ArqlJyMvqz
Jv4QVhhgUT8w4lvOT69E/CD5oeHJGHHeuIPpGd+VtKn7J36unr9MtXo+56X8WHfN
NtsKu0SKFq4vw+aT7KE6mGg5W6uEMOwDzd87kymhCF4WqmhmDv94aimA+ofjZwRu
NbP0ANt0Nd9htlTfSsUhqh26M+QlgZey+pCLPdTnBTNeGpADOGTWwW/g4c3SXIi2
/+zicljgXwTJuzXcWDiIYuzgoShWvVveHPUjvcxnLC+JwYVR2btM0U5t4EDAsbML
Om42j+MuNVwnkF86tMO/c3IfGe9L74MAqFGg7peOoqtqdZFzCiH95H3kKEilagWs
IxRxY1ZpUq6dlZ55Z+ACAfpTdLsK/Ryo0qA0Ypa46SgoX6NUZl9dZgBc05PxhoO/
yLfGvAQpwIgiUJuEeCACWMkkQCdu9JdC2ysLMGSXT5DBFu/KU2KVKbR8uB9Etwf9
UfBzimmhcsx/mqLZnbSya0L492Dj/DNThEbE6Tu877EF+iAnWDZtew+2NGKr1BIP
9kgxSe8s9D/YqFjHVhdi7HFtP4KKosyzCm4e849blyXozeAEZ8OyEmJ7cq6Yw3W6
NfFZyTAkqg6WH3aVgP8Tvvk3nns5OfBY2K+20DxomfL/331YmRu7XUEISBYJMmJK
JVm6+vEtpfE1qfrSTUWbYDO75HuzYTk0suy1Gy09Qkc9PLQ7A8cMSeNnYrtbWagk
Wm9xLW5dNWqjwHPeSqrHIH5w7H4HHUasjYwsWwFs03VztD+Dc4Aa9S7lioAaLvrW
j+TcyY39C1Kq9NzOFBVKcYQ+iBXP9PUOIezHsze9gARr8lb1U72rt4ZVZDKeHpCV
z1fVotyqxwj87xl1lZ4AcY6bIO9YTwWKpcATyibPS2tYWkTx4GHjKBxAV5yU1lzm
/t5dvkEK/kEy+ghfx3UbLy7xqOgYS/jZC4ouI6MqP2wZdVl9CNT9Om4NicP8FRfl
G2eIYWbL2V+s4eDsBTe7fjz8FbuOTqeKJphyYGw78XoWV+RIpvrz1agvMm0kogNX
CsYt5kUryT40p1BpvWWRFYhMjjVTKxDs0Jp1M6/t6RU7U/f67sYV0tyvgBEmBzZA
acAR5GapwIJD5x3z44uJ9pakN37mWUAEkFM9Y2UJ6Mw3r/r5MKo4jl7PIor7tfZq
Cm6wnrhZSCvhTTVUf3pTN4B+NfAcGWWrMHSYBEkoILxMwxVBE0QjMTPYgw4A6wZZ
bk5NB83DkT4TM6g0qBpqU7hlHDevZkhUsLUmrxkutl/GBOqjeGUtjDO3j1FuGe4m
ZlVIZbuwtgd65sx8qWAWYQ7viHZ49k7cNY7fw9IvfW7D7o+Y4ALIZMsgWB1i6Cth
98ZSFiCWAsI+rXUavvXuEnwoBKia1a1eSOERU2DYu6HvSqozEdSmiqZyjn3st6B9
xj78U7P4pS4hWaB2ZPDFgQ6GhDSs1z47DXqJ/qAqi6egEy6CWges7GT744Rgskw1
wBwQ//RzymFrsztf900oebUdsSNzVyOlZQq8yZlrjL0O/xqViRKKWD792q6J7W37
yMZy6MrdJ0mQW7bieGzKkyyHtXwuFIBU+qGdf5oj1MXqCRTWlYRTn6ionNz7Bl76
cCyUOvSibtTvSmhvHbohMOABtHYl1OMpJEzHFuSobn9zCSMfPEsABGPKfyzKipk1
bVEfNuycANZP/6X2sSNqQckOcqi+A5/T9oudHqldgRoBct2/W2wxJFiZlg/ulqpg
dhutloz7d+cTXgwWXpnasAsEebNcVOAYKAWzo6yaUHhJWjY6L0QbGtj9krgLSWp9
/Al1on1/iIh9too7RPWwuS22sQNaVvrwlGevrfDLOsn7QfDBLOOqm/s0YtEyXieq
lUM+gCSBVcgT2MrqIgICfqZyUv+PCZmuj3iJMgkaXb1Djj9oDDoNs5CnnWQRLNPS
34rTVUU/7yQh6NmPRxyF6u+kLxGNd7Ebp+GYlJWL3JYwzkG6A+YEg3i8ng27DhGD
VPF2RiB7FvmbJ1QtStqQ9RfFiVTHMkphknW94zt4ZK2YBt9FB13s+kjP2iIV/k+v
AWLl5l8oZeqRa7kNsJ2JVIlMCOLkXrhNd+CpOxZSw+oVG/M2kL3ZxvvbYn3MQ4SX
Vu2sFavk6dcF/xpEEkzoQgO01VbWUAJNcrWllOD6s/ncgVa3PrCs51dcNqCwUBxv
9rj84REdLtNEVY2a3JUFiWBkB97GdNchUEYtVbg5uduSKu1t0ZpqQaIO+Iy5ooSD
W4CaJPS+sLwvQI83oGUM28w7neZBF8Vl9pYx/8dW2Ch7zsBUfatZqLe1yEd02ueD
pTupGtS4yCp8os8+bVQLLCkQKA1dOMFKPrZMF/uYdJ6ELEoPbaAdhkgYrvKpmigb
BRTkoJ6iZ9Z8Shl53VLPXKiXWCn2Epkew91eaTmCqgtQxsn6mpBgUc3iwpfNe6h8
ub3wDzvUyC47DM+k8gWncOeZEhQ5T44UuakJWt7zKo70EW4NvBHvHADfMFlkDrrO
DfdkJ9dKupU3LX7TQN7hTZaB1/lpDWDkwbVMZ070dBG+KMKL7YxLnSEeC3+MOKbO
i7ux9tpDfauRh6z8jT77EuxML9fRGak0g4D8grNQnqo5QZ5onKsDomAAFIqZyrv0
ugEa8QNhemGsismpxIkFVb8ezlUHYGMdKGLXdS/JTyKcjz+jUayGkoPgGjteCxEZ
j11Auj13s7V2JNZTQnt0rQAjoSTJ/YAQqEysHiRYNYBRptAiOCoTnkjprP2M+Gee
u738pcTMxWL0nWSKfUi05cfMeWGSiZjwCE0LRZYAzthFki973YYcyX0yNtI5IFjd
AmyirDUCXUmT0CSyD42zZ7MmytuFBWHFEPIj6A2Tgkxepl5MRSKINVshn79Js31v
7fbfxmXKwPqlu4gxwwwmj5uZaM0QJ9MmnYP8xymIGJ9DbbZozf+n5nrR7iOrVS30
gE1VUs4VF14zSnAgj1CWXGmp8ij/pMqaSit2CEYNj9AhXkXCGVSrRKYw6nFaliDQ
VhCkPOdXezwn0TOgd8nHBqYDUd1XkIr+PBpKoaBW6fnZnIIhA4uH1ct9y8WCgPb3
4vulMd1SWeZYZoloEU76b2CGPszzMz422p2FfkzGleUR8VqeJOdBhC0FDjnERzyK
C0pbQ1U8HOy/uaDny69nJ+fWoKQqK8+7UiDvz5e9pm+bU/cHEksWO4NRqGRAuSMR
yWuheQf61fobpExIIxoFxgkKJJCcnHEo/EOM3rh3URsdwt44yRpAry+IaDTRkNIs
inIYFj7yYQmPFXXYVTlOjMjukuotlc2rl7LK/ed6M8CrW0aqBrJzU84+7Gp4tzpp
tI4JsjdNemVZO5s+pYe5JjvI3YMnGmqfmAKu8GpVRxHFykPlRIWBCpwqOEGio99E
zhWT72S+cA36VdCtAgGB1cN/PhfBmWKueMtBOZVSK6CTJ6eXQfKPVa3qBL+iKZIq
mYWupEC2iQBR6zKv/S/DFgvdFdI2uKSjQIAvbrZwyx1ynOfUEyCwRS1ckYycWIZ/
dbYcPg/9reNlWwv5yOLqP3brBWae9IxZCQHh2GI4EVvCRNUX5yGW55lRd7xSO1Sq
xbVlMhdPe6qa+YOo0xEFHQRPeBPdU7hi70GUBFGaI8diNIN+FuQ3nblLFeXzQQGK
nok4JvdBVmL4RhIt6XfC155T8W3rYn2gkVihdTW+5adZ3FcM6QoyUmIUQT9D3Yn6
H4ODfrl9UoKn7e/zl6HLFxv2oqxPzK1zUozKz1cQbJ9HTjhbfu7wmmARqacaHtxu
rDJs2TOmvX6kOwOtabPV2fL+aei4hfSWr4AegmzUhtQ7lobvWk1bIhIcFQ0PMidq
mr8vBMpNxnZMzEklouiSzx29JUrkrCvMm3yguG/qTl/zMbG+5VnQH8Fd8hlWCUWJ
aRKLtZ/a34WVxdSM+oc1jQbZH9WbzZiT0LG5XWLHjYLs946frZazI/wqYTcXYL3b
GAt1P6VKLq4xhZwOgWDXHeTzitXwCTwOYtr2dTeYTfiPjmolygpGQKoFp7lu3kqf
O4aWHzYNM1bmISIeO9jrAqr9kyHMUZJVdSlHbmBgXVgHDAGw3lpVzA0n9UmZ/a/u
kcxDyd8qzS8SncmmiwkThWgn/REKBzy5AnTQEqEbHaNZcpizEqXrqyvCZQbfc9zZ
5AuXP/Nut/N2U49nuCcbXEVXaiwhCgk9FJoG3lIl3/lCJ7ShfcmzQu1WTDj1QnZ1
OWJSzbL2TF2sYtqqV7e/XLNvYJqhh2l8sAeIahJnoKKFWOadCe746eHuqahyUcPe
lM/cJsh0KSJ8tvzGQwyDG+5Avi4OckQghgeJjKFYBaJlf8vSxyoSPjSjQQSWAsqS
U9wxs7xmbAI1eaGqb7vXQl3ZjBDpBG68LXkE0w7YkA+E8EawLpwk+GetfifCk01M
m4atlkSi58FJVLwu+O9FdX9XxpfRsXnCnrfTeIZdL0NK3ME1SaSx/4XFBgUlrUe4
qE0aVw1I+hAaZ+mEEXoxDpypAwSMXSns/AEpExrPT4ytZa3s+R9Q2l5IlZCyx84e
m+MMwcU+pWYJ27xTOUQS0fXuL2AjMOub39ei2aU07tG8Rj9FZ2HxPQ1xXYZ0y8cC
2R6Cx3fT0403yoEvMHoxh38lU2xi3c/13EjnCmJoP7cDZnugSKC2JXutzIXiJIvf
Z/gfu4mwbcb3oZ4/MqCVi7U/I7LZcuwuqRswBKSa1WsVifQgisVa5grJe52Q9Eqf
ARMBJvNi3EjFLZJwVvQSrPlYZZB67xbxgUsBHc6qEEphaYGV7bdOjVvVmF1TeIO5
px5SPkSEMOolq5eUd2lVmEhkESu4zcYUo9AEZIPctVqCoaKh3D997BOIhHCezskN
i4MxEjsR/ZtBkmR7ER97+f8Adr3JovPhwmgvmyEgKbw0kGfwm3nijsDyaCxI34zw
6Utw4LuQ2l866BcgHlE8tC9D5hfOtmvSijaKrPKbuybJ815stjk5HqB37EEiZpKB
Z5+HbZii76SjWFUTFVV1VyvMqGZo1BjiAfFwm2BmxSgTZNo5Ak64kaQWK6gQy3H6
AoSqmEIBDJCqeRi0tWwnzQxx4alRDepauKwNawvOnVEsUc9yxSxGA7SVeOyX7kos
+QUI7nBntavaDeYjeohLFzmzHI5kYmdOl307bVcO0Ta1ccagwe5rePg8dAIuL0vP
sB2N6ZSwxqcY5BJIG96T6S5Lp9OVIoAj2OrTyFy7dJxC/ajQKgTJAeNeOPgQaSqn
0nDPR3WZLCAFA2QnVuePe6IjX7mAW8py3VIIkq/5RwJssg7Lav8SD2hqQq+i8l5p
E8EkcEeEO7oHdFwRVZR9wjKJD2UOWeFohy5Egxm0Y51/JRDIf159YLNnRETJgKDi
H9Seu4FzvOhUP37dZay4pWMmVgkS9QUbIF5WCp2uaW2K0WAqHg0w4rnNlQ11jo7v
tNgVP4HA88tl5dYlg9hMnt7kMvs/zzd/RvCDybRc3CanKCVL2qBLH9YG/bX/uOos
Eu4wqJhckUYQHTp41r/4WRuSxlO0KK2XtHPpLXERYItTNqnnRF3Pj5e06VkzQmlI
aA4909UXyqk0HrSh8aPZa2EIDdhZP8CE7/GhdSvI5fAkbXilj89WkmkXxsQvqVvH
P9YDabv49CSa7Hh86E8UPsp3ZPlLVzyqfnhwF4tS6odDB3QBFK4k2kz5Q113qbis
56N94/JV9Gl3MTa3nLwL7huYMh5uKQQrU2QOk1RniPyCWZZion5oOSdwHDSOjV6q
h6iU0huKrUmDfFrekXbk8cp6oGCf4EQzva2bt1wMp34tcltuoCesEnmthvCsq74k
RNlO6Fqga+4J6lptK2kYWF0LX7RGdnIqYYK6dYZpa4+etwTBJmoybnCwaY46XRYr
JqrxPTsjsD/Usv6eVnQmKeTCKrN1KfkAYU6luf0LlU7MnJ3bPDchTS5sNHsG6Jck
xOBH+EMGq7XxfD7I9iQWjWn78O9bbH67R5O0zafyGScTz65d0EHvvukarR2qr5LA
6VXSS7u5L5pamwsBvqem+VKFNyEX74zoW9gijp232IFeb9TEICpkWqptO0YqcKan
B4CAF3iQnNycr31ovmjmTCzYTIqJp1DFcrWAUPnFAJZMY9xb+fY5IBvdrahhefFq
Yf6+LTxYhtzfMmR3Bod3xYFySzPYF0G8AVrgOLxRUG6vIecV7+0OtAoiBC483Q8A
lDd2bxdFKUeVJkJObn7LnWYNtnXgXapH6k7dTV/EVkOWAunn2Snuzy+4St0kmrLA
jIqvIN7ixqQaKoYiIA8rvR2IBCEdLYX7mqAgF+IKa5i7PgpLWCYfntz2XK5CX9OP
YnaSqKx71yk2lgZpbiZbYSjd4vfKRq+jcL6eaalmcZll2B6LocGuwugZXgBxhTdE
RdgYshec2EBHi5JrOesCqLnjwy0rw81I12Nxn5p54/qXaJQqhS0OCGKAO+qehoIQ
yPvGrF6sFDYR3G4WUsJRn2fWdM0gcy/P+jl2WwxAKNKERO842Ki6wH8zRv4fN57X
lpuxMIo4O+HiahWXubzXeSdXgf7STdi+4YAsJbp646a2e1+WjXIqvonAF5taxvGa
k9knykONNMO9gccz3p9NvTzf3q+92WwWy6uaaBZEPM0/6ZZQkPObJ/sDDQNyq1vI
MUzHjaD05zbgO3vFt16+S33F7B9hYfQ1lcDUKgU4GIrs/Jj5she6rxX9wFtvleh2
E8uiALrY/8CdsK4Lm0b9ZICdMpkU5zSp3YwezZjvEAZRWZ7Wm9BxqNpNh6EzevwA
O6Rz2c7fFlHB9VNAWUOKcAGj1CLHxV3+gGzC0ef5imf+ChxteN4HCALxx/vC47oD
6qigA+kOmjezuBCxNwB6hKQgdVKn+Q61Z9vKOe9dNbEQ7r1scf3aP9i3L2V52lRX
jbTG8t9fVCFQ+VsEOnoIbf3JU6CutoEXGPLY/4ptq48HNwJJnkXCkDY8jDH6yxg1
GctTd2J5zjyKxkfLJ/eX46BT4eGHYtQyQRrmUtASZm9gUeILzJ1GOoVAUyBElZBY
5vE+qr/CyIebLXN6Hd7WkvIY2W7/Uic7wrjJ1l/6p5w87KrQMyuNh9yO2tBSf4Vr
pLc+VoZxcTrn66Soo+USUewDH6Wq0trtUgvj8LCTCAOQoSMSw/lKWcM0YCdbbHek
VFZ5lsMEuxijswblRQPeJN5VB324zySeB+WEVkmmCb65TdCegteWDG/LGrA4lA6x
LmadqVUd/P47oFiSsSpOgT4Sxx9F67qRuboMcQQ1lhPinZibG/ST1r+tsJBQhXnq
jUB3FVTXKnp9j+Ppa9PP/+lA4N7a6wEFl4E6JDN2GsuzKgY+e9jcWgMKj0Mh7Ty3
9VXgXXhsk7RGu+25TQ/loyVukZwIzuhzzH/PS9an7jP8elRcmsu260JVohEtTPlh
+Dtdgkrcp9/sOoKZAg17AajycDfDyK9ldLaMMnG9T1A1LkObqJKAY7U0JSyTuAnS
/aTFNJwy4n1WdjEaXMxdbVKoAf/BAWdZyIAVIt22okBaSwc9x+9GoljZwXC4QCn6
Z7u099sECqcDFOje4/hkPTibQCxFb0jWixBw58VasFzNY0lP6L8hYIQN2G39+Z3o
aEkbazGhuxF7LWzpVrAn8lLJtN5KoMjyUB5IY5vxTvJt2UP/+VKcFSwBvpAgQtUY
b+cY5fPyQy2X4ClTmQ2YSfc5gjkHvXFvQRdsxSo/Oqt8GS5dyoV3mNJQgHhPk9jm
WymoJn2QtmfzqC9Q8nAh5jqoxGFXMG9an8RwRQsUJwt+bTScWlMoZvk/Njl2CaLN
N/C0SDBh6VN6O8gjQkaHZYGDCwAjlXNbnzwp/+xkDGyftOXnix14rbBHItUBqUrS
roXQGfma9Wiw9RlXG5mxZL++Zd0IyeGS5MSGKjZ45Bcf5fwhqM2bJAHXkGD7+Cd0
QElUI8wd1O87QYcWutxiluPwxGaDvdsFAwu+S/KnxdtYX4bmtUm63g8PH6JafTB7
z5r05bEWU1b3F2sI3xpWmBnRMGKJhvnHlleISStmbiN3XNRCR0Jie7MmkEUWhb8R
8jhU15k8Ai+zLfg3TTiEI25R4o3ctC6i0m7ZtPHnypfyuwbRvTMSDOgcyP1wdkmX
8sTEcDM2olNwVt9+43927ib8XTYbPM7M+p0kbv5EBHhdIMnt4TLytffWbT2AW3Il
0H7AP8/wVXXdI8rm8JdWKsv/svjGcbZJlhoCXo+guR2T8TaDhMtSTA73nkhSDjRx
FSddvrN66wx+PUui1cJ9HMpV58VrftkyLjfmMpT0knpYJkl6meehw5xyq3ilZ8Xf
UdBnl6ym3TET0kIWtMABeuzOXupVQC1BKAFoa/VqtDwcPmjXw/tPGAb+sTaF+WND
a/4Q8rKbAUkMmjwMKg7O5yRFZquiD/TKwrXDlGlQrZB3sO1SXg7+f5zyTpkijOi2
uKjyxWk8CdF3Ud1lJgHdAhun+6JWDhNWwJf6LC8d7SInkPy433DLiKfV+nBmOO6a
55kMpBuzNKEHQMLiwco8wrsA8Ii9QPe3V0hkuWSrbfxZB1zy2KbcY+puSjApirAk
Vwi+PhRJNYG/caP7iwdyZuHXPDKIi8oIMHgN3WNDuJod+2LZ+JYK2EzAo8w7hHKu
9hxDVHhjIrI8H5HYVTh/RQyhIA9n4c2HqbsvPvKCxLNrSBT7DFRtYuPlN1AsL25w
Ey+++I4Q2+kOs2KLA+uKlfGo49qt47b56IIVLpJVw4W2kDL5alFnj5Fy9QO/RX5Y
8RQn6gNzKjDMqtMvkSmZa3h+mWe4X2riYziYltk8cLl3gSytweWQSB+fmycUSyQh
Y4MTVaXm2EZdUq26+3YT8kE8bZWjvlEkfFbNYS/YpOpCAwQtzQmtEJX5kZah6Jz7
mIp/tJGMvk85zy7pQd6wRA1+U+DViPKTVHt3UfoQdWwy85HCS9iLXnaUsG02uXwQ
J9Hhf3qIItjVE3FCdefq8Lhb0NGnJ5sleyaZ0EQhxCydwNcn3g3mxePcbcHnlG8v
LXN7FpNZY065Lb60co77Gkqi2NMpTrAG0P30Fh6GDN+IoMZ6EBov7T+ymRfZXMek
aO0mfUUXsSxPcuBHcoZ8CrvcaZYLSe8PoibEATM7TItSoysudmX7Z0ZsRKgH7/hS
xO58H0tchTtMcTpx57xF7fLitYjk+CU+FNVjTJcbMdofAW6mskOPok2Y7mKRGpC4
gkhRia3gByTbf5Y9PxRlB928Rg12B0nMsqnDKMjbL10nDuoIFJO72U9Uf+czXtzD
ykgYZUJAPzmVkjOz3bbAsyJrnPObB/Zn1/bXzDKBDwx17o065NEwxS7AGsR7EesM
FAIlZY7BmZ7DwGg91VR1D0Url2xqhPQ1yr+pV+VjV48NMQd/87m3wDacuo2CXkHX
UghrRX44iofT/p5lmVGCHiLKc2y9UPRdr0RD7HdShX6yOKwm+h2Bu5eM0HIP3GBT
wxHm4LUQh39zhVY/yYRaIq3s8w7082ZlA5S/W3CoJQ6eAyAan78hyoSLTUJbq2vk
bmVJze20trP9Gp93YKBUOnT5fMoOO+IcX5aOcpDcNLf23dlMBn8XYSANfu+Q57gC
r7zKmcF0mlzuUYVKmspH7Lkqy8YY+AiEwAnHqJegylynomy2GuUQhTrJypbgSyaO
hIt4febnnD96HHqSUcoEMvRFnxxhwvZj3Fc4f2+IdM8EV9ZXxd4ZYIdk6nx0ycAK
5XpZ9ThjMsXMr1VLCrJygteQV4NjeiD9w1Eqm/sZ+WycQC2VVjnEvzooxSU71A1T
uj6wLg/+Gay2pGbXce5j5daUEtVfhWr5c3OWZUtoWVNq/7G4UMLjAA1JN6WfGm+Y
xOREJ+0YydFlin8l+7garepp74ABkxKr1hPHFXntFsWrXPsjG84mAUWPYt5txGuD
thEDhdJU8NsjSHvzxjL/pwbMWzp2gvxG2IGhRSYYrAlR7DlexQRFAZj/HRQB4n5r
CdslzqGBun3ps0D7AJr23lNniLFY1VicUIQIWriRp84hzeBL21jZVtfX8veqiV4S
8PwIaJ65JiZ1YNiZ3Cnaifl0Sloi26TxaiN6eQpZMNIfiut0mWhdgfonAG40DgJY
kv9MkUJbA1S2Wugbo40lKFRHZUtsWiMwDuoTUd04A8QCq4O7ucm68eCKez1ySGHz
TRKJFNLRVzKdnjat+RuiAi0pXgqeNBTAXdcUX1LV9acdaujL6zELPo5TBL2ZITUL
tDtNDbRXU17fAyPVBhibavY/KTMMvk5/oFEQVYdJiMl7XArxBJ247f748AUNdrso
ftnbygq8Ul/L/QrXkgJRuUVprqjq0GLvkTmq6mWwG+VLz9j/qNdKD4dZeNTiWisw
EWNGuvQY5UO+FHQJiqcP0h172HWTT8oyHe6z0dPR+Psy1joMTpgAuQ3alOWaRnsA
nKgReNAE6HTstu5aywD4on2gHhpVl/aW2urJ5T/0KO7tqe+ERx98PSkowXvOgDHN
4HIDGGvjQj1UqBXGTqZDI7P6N00KI5A3BEJAYqbm7HklYdQfIyUPnpxU85QUmqlV
RRC6LNkLGz/eXaF7PvE7kxq4QFruCZVFrfIyC8eejEef3x4igtJnatuKQ+unIBIM
LIrOHssjcD9S7xYfjX4HZXmGxVA6BKvHoQL8DLyb0h3fXO+UKCbfAyaaCiSQ8bgt
hSG7wsXgPqZNwyPI/KhGAP5QjwvD9YSDXc+ULXQ2woS6IQh3DWrNlrZz10JGkPqS
4IKDDr/qVwxGrnK9oCJHMyy032iKCrJ0hgl22O85QVyQHabfoI4VBYLLrPI7AKh4
jsvyeO2p75B0tvhHfsLaSE85EPyZTXMaau+0regpdy0RU2+A0aZZtO+9gjM8Erwk
Z8BMk7GMGRS9TI+KOpAi94LT7x3x45tJyyT58ksHGrPS3ufup6sbinK64B5soqys
oJsJnw070on75Qvxc/UHFUa6pQZVA0OijJX7lJw6jAWt5QXZvu9aROu60KvL5JkC
ISGuoUIMxYb9Lp8gWy9x6uIfRVxSHqRDqj77EGHtIPvUttle1UUadBQHsSnrF/g6
zAketDtLIRJOYKuTeu6ciOPsp+OdIJAL71qpcol6wfnfMezDjBZLTNsZA92RN2/z
suDExvmUNN7ilpxrObTj+HOveMIoqSyqYqzyJjhphwUfwScmbOPiyfgdSQI9BJ+J
SYvjNQBpAj9xRGWxWlOE7tQbQNZrFqs9mQNrDZjTE3JXf6KVq8QoaPvRE+Qnff26
NVCsnQOlWXdSxqpywWzf0VHUSocMryuigOk4VJFNgJ4DoTBJ+JfIeTr1FbLBaD0h
Kew37UxTArLlnL33mFjTF2oSvqmi61JOOsPFxkNLEOr4ACGjBIJOITxNtn/h85ZC
lX1gif3qIaFvGZhrBiBW5nO+jqivHgvSSZtapQzx7PabbZwCJLWvwe8uDPQp1PU1
tZ0y5mcwaHJM1QKmFC6OeblOlPr0GLBhmi1PIk1RVTYfqQtQ0G79OpJMj/3Grtd1
CpA03wqahS7SrW0c9orDJSmTxsflW1quhpGYJN2MQO6kp+2LlGaL/0S1afsF2qJF
lpgUMG8OZzBinF20HhIrDCykbY22FGVH+YFc5gdvBydUf8Njv8c+kokjLHQp7iCa
0uWRjhiRrHInpCrIT0BiVPBvEsaoyxa6CCXERjUkpzXUb1ACa7hC7hEz1yLKIJ1J
jXsNBOdOsB2u3FKXs1MOhhaMG6wI0ScJqKk51oIV06QMo1xq5HHYEWgWURIWJ4fR
rwYRpvr0vnKP+tvRF+v4zeavgMtfIPjTLyuIp1qdnRm9n2+9o75/UmUXFl51vZkb
I0ZjMGh7GP5vyFDJWxdANwQm6J8C4+2c7s8LJe8KJjzNin6Lq3KWiaqzX9+Bko4d
HmMcwQqkvK8sP/2hOt34K4Yn0Wkr0bXrETIpdPI/6/rWtAgHkoSXOTjQW55Gnwhy
7G345EJHsEsLEl3mHokPlxiOluKqIooEl6+I/eRkkoOqWb8jceiTa/YPPfZsjAzJ
BpjRWH0WmNEBDz0G8QO8uRDJwmXk4+8zwvaDGymBpNbLHoIzlmdJx9KJWcCTzBiw
BwAI8sKOhOmEtpn1Cvel+pPbg3VjmizutDPGv4MmgUT2ECPOZaA3w6tX0OOqF1iy
zexfJ4rVE5S/TRurrfFRwmygKnzjJbEs+Gp2DGKrJfZ/8xDGIFUWn8kpdoRtiS6J
9o9JamjlAvR7INQj59KfnbKqftwMBshqcYuRQw1QMt/mEsF3A78xahBlN3I9VtGg
SGfmFMPu0/QD/vUMOpb0tEqfCioMKgBIov+7/Ir/kSfaYOZxOCL57dRN7HI92GzC
JOQb+prL/3lQG9gAQQJKPF2g/BKyJDQ5fSOD/Wjzuo5wtsc5h056ccp6rPmb60wr
jvIrfyWdAHL55Vs0oIKzJZVEwAhqIyEMTSDGGy/lzayyAToWt08aDNpIVCJmm4TY
siUxo8t7V/lBYyNsv78VCEwN8q+i1LMTgDBZd4E6Yc1O9fGD5G43Pvrc5PxLT6F3
qqPZU5zADTe+rlR59w6iDjkrzann6LXpA7enwswCWRfzj8WMepTGQbqqwkAeoOG1
EnEUlKhlQKNIMH8qfDZAxxBdcaRVXrkrMlEJZRsimtnIUNVE9hbLpzmFXexV3eiX
Z9YjBrFWpxvl6VCwp4R31gNCXAiItBXttNIHZtBH+0IwS21MS+vs8A9hqXDmhXNq
LCkGg8+78nwK59UTEwg8IBjBi8Hct25QA1tfmKfUBQejtAzEXpS6xq7Vvwb4qnZE
pjm5d4YbLyIhZVyqFA9upzuiA4qzVA9juuY7c2cjSfGCepFdpDbyWvrr/LoyvLso
4IXZJWVZwR+vcgyUeDDsSjMgS39v324suf2JTdIgI6dlEuka711uBTkC258dT3XG
xIK2usFROMjf1e0lBVrG5w9MSurTG62OKRU4DY9ZBthnsuDJSq6PoNmHlzgvvlji
qGYMhiQIC5KxpvM26+0+N5hPNtMYZpe6Fdm9/KvElhRM/By3vs+1vLscYBUzIHX7
CoNb9/Q1N1OrwJsaxovN7hsQ5pM6dI5qZ+CpXoM0O6U6Bn/H+L4FdR5heo8or8Si
3Dy9px5Sbb6QtlG1EuFteCKp8mD2r7BdOMiIi4j7Eu+N4HOP9r55RiFdqiMJSjNx
sVLb8cqGu6DUNhmHkQp2IyTXOUTa3fZ3qmIaPqt0Nt54XJGD8kCd/mRZ8yrh7PlN
NabcC3+x6k34rTOnCNeLQ6C9LLMkUScWqVbMLGdDc2V7A37M9sTrznHJfjvURqBr
qrbEjoVVhYiqkYRjMP9btiW8Z4HUhV+9OrRi2WMSLd/jYKRP0m3PtReSLMqhjzzt
32tjfwsrTjJpkZaEYT0dyS688q39fKkCXOc9ygp6WPX+5SpYmgsE/BG9rvN4Vu6H
JkzLgToDo+or6gIxY45dOT3u5WXcstDM/C1IgYFpHvRiTC12oZEGspSL52+0qJDT
CHeJtui6apwgfzujtVZPqSDye4PWgQ9opRc8Gb0gpCLmioyovxiERefpkV7vaAuJ
NXzjDdAWZLqnlVVT0sSgz6orZfF5g0uQRJoeNs+VSW97NUSzfV/T8QFguTliga6o
Q2X7/jHiAFTRB2QQoxQARwRouDQEwMABRpB/ZTKed8ZEvywHFipdwKq2fhOOdqKj
1aXftI8PCo3ELoTJChPaH9LxnRAWcjYsZlVncMNNqcbhecMvwaeMmbS8x1YIrLRC
u5z5p6hOIGCCs2B5Poqn/gitO60/us/zAKx36hjBl453OxL06VkubxYq7B8ckCQk
VPXrD2430ppiwgMsuTOo5riGxvmjYEZqAV8y8ofj/bbXW+9GN5g0BDQk3tC6qe9F
AU23GFIxNjGCC61UEdWVMoPmH7ubRpUog8zwsjvU9KV4rk0gX60E+dR+i73UxVrX
DLtHF3w4XVOpDaf6lXhAF5CkMBM1whVyPlwLGfnTCaXnRNF2kMXXFYcuoHeYKx6J
n/un4vPQzVmZRYazQ1FSj8kaqosqWhD6iZlMdqqX0oBHwlSb1o6Ivxx/ChU7uih0
dmG7NVRXMjGBiE7xEZZmfOpXpldjRL10AK4vvjsMI3aG14/Rd9UuRlWzTDIowApp
wkBIT0Xpkek7Y/5irV3qzLvjKxXRdF96OsaDeUVSU4t4UJlxbUbMktqEOFkTAwqB
cHCoIBSsfzl90yQsXRJhPBYipOTwzXfUgZWM1aPV0aVjc9QRh6IP4FyY5a8RC2GD
SGy8Tc90WvKbKdK3AiWOkpPHJpLIEXM1P6LUL4BSzqd/UfXGuMMKl0Am339aqXj4
sOAigdP0nBuA+fkQiwLNDUEqVuwtPNXryyc6WVq1M/9a6OiJQ0iFA2UW5dFSQI5Y
d68sougZLysMnVGyg87uLglRh+aYFoRTVQbZksxtWwYszOGUUZ+CI+a1DC/xzmQJ
wHUtuIw1WT+Y9q9WjRNkozgkc3Jq4IWDEdkghhOfTl4X8CSM5HNmXAlnUgXvZ5Mg
myEXHWzAIpNm0tDArsie62wFXv/YnDVkTDiNs5UqWW4mMQh1vXzzteEmzl1qiJid
+N6e4ID9f+3bBVKK2GmegxgL4yHu2CHlWBC/R89VDiYXtGDBo8d9guhTCXa3LhXM
W9iqbXTnC8MHkAiCIZQ8pH7oy2iWymrQK1udaZSD7UwKhfnApq6VB9VNVgXMpXHl
bA73HCrP3tDqTcXB7HqciwgVFBj8XOeMiYq/5Ift7InkOYMDMb7xC6zG8KokxMBP
HrCo7zR2MXxbXX1Dbs0E+PsU50nqdW0Mp8I1oDXEYVEfp9qaxwUaiwP+QquBanAB
p9dDdL5zLSG46FfFftILDWmgnDz1/gfpAAK9hBRJRVL8I3qhVdO8xnygpHDhj7e+
D5ka5/aWnaTDP4ZF6rcrzrPBcOklll71ITAw8m9Dm1PY9EK3WCqNA1ijvBRvHgRB
VnSwA0bWTgjB5skl91JGkZEXgOVTAOknVSJfTMDUYpRQfbWv8Yw1pCsrA2VVx/yY
zJoeEYJ1MMxdEuVDIbybotmyYIzxXe+2Lawc+rYlY3lCkW1k/Y2YjWRvMBWEDWc5
VRdrSRLe9vBuvDeRGSLNbhxcibivbVf4y4/BhOl1stUky2lGmLe7vvrUjG0I++ax
/bgoTdYsAFwcqCeNYCLuVoR2n+MKeFHNuTfj0C4wi6BX3BiU5ypr9hi6BUrmfKHa
UmrcwRbr2Xc3Hhchfzu/OeCQdvQGn9FMbwg2K8+EMfBqsupSyucwVYfSn8N2H1yQ
VX8pbIWtB0Z72gFAgdfpRGd8vx4584rkxfs/Bb4SKhtxoSgjEGKwqRD1u8fWvwt1
4uSQh4+fEqQ7Av9WOnJgiQeSKngQQbveWs+IDLqAP6Kzu3ksWrX4qBMt6badwoQj
clUjiwRzJEj/fSJcDyU/PBH8iWLi7QF3SFOpO6lNECmEZWznyuRpU6wht6DRjCsn
Apx6c8gDq5kMRrhAJGvlUAvPUcNfWCDXoTi7KOyx8y6bgyOdySEV/6EFaTXtLlm0
rrxMKR/6C5Nx0MF7djyevSYRp4aXjvG1RXysYIf5VEgsvuDQqw6RYWsu1JGy0lkR
/Yw7bLIjmBkBDo3VjwYYOuLHd/ZAmHslXqgsDtZmYH60sAVl0ejzpGNwQ3AKZdxs
ptaLKpc6/k0FcL+ynbVaUlqoFTvVSZ+pBpDgxF4NKuLM4Kn1StgiUl0RWEupMqHH
sYMRWGbsCKEF+Qvy3PsAKX4A93tlMCcRSJMaNIXj1/egRjjK4hFHiRjbT87GBj4W
Gwte/l3g9zWb+swih8bwYuYTvYel1D4vlCVKfTcDNbv+CWLLscIsLPYQVBJ+rbNP
6NoZ49pE/603qkSRGhHXv/63iaxKp6Y2U053BDGfGFrl0RtPPYxMVrgjxfgdONT2
sq/lDLaYzjT39Fw7CZoqNcAZWl3/ZBt0Vyfhv4NOcc2BWsNHE5ESrAUgF0rZR2Bj
sYPLd3Pvxs2H5EPeQnJXdod3k916OAytDTNaKx+h2Ef+Cn0QW3Cz1gldEm+sQ0dY
xYDBZwIZIBNICSO6syu1WiVN35gbi5gEUCTnlsqlvrc6JjG9ZR06Dsq46iVk2YUH
Ftp1rwKPPdzu8YypZNHNcbEi0idIiWsRCUKklqaUtvv9F321kWHgIrOAHfpyQFXg
y+zcogGFm8B/RbGElJmFS4LuSbWicwsbqh6jd3UGVg/fByShzytxyKBKQYCzasc1
vXIzhQaKs+eo2qoQgO/W3K07wWSQ8s46Ejxc8ypVrWBVMZRoHvtdTd0k6s6WAbV4
ffl/MzXkjJ4X8bbiBUhUMg6I0G3rv0plvJhgcuXsXA7XPRxfE2R3htLJYWU/KeuS
OOIdxkF0LdrY6ffb/UeDJqfnAQhISXL1NQsdIBaGdQ+eG4madeA/tYHIrf31+ego
O5ELDHi/N6IRk43r8LzXvxskOGD1JnWaoYmJU2XpuaX5a5MS3tHSAEZAcDuRhkuM
NBJSTo2SZRmypTz+9ZpUogadGJdY1m/RaJxh0JtCOwLxytyRZ+mTfzYtZvGZZsfE
WOdm8X5iRaYPemnWieE96g/7FHoblrAfUQRjKjsNK5Ci3rOkUES4y9q6jAd/M/EI
FUitemJ4acWg7mwh9rdDoMbF8VukGnHgc03Y5gVq5WGFcAhfmtJpl9IPn7cuZJ6s
ghVqZ2sCImJXQTjDKLEDAETyW5haS3oZOhb8DcNRkm/IMiqDl0HnLWTAwCkwSc1w
EIwLMFKmATpRvOe+FLh+ktESKDDVuXa/qCuZxlDSNtTafZ98xwtp/R1HNIQv4Qc+
4Nf2lOJATSI1msRwcz0nvqDd3s2NlQEiQjDUfcSDA1e+yLPu8LWr4JYU2TiF0dvm
gxUDoZCFMTszCHSSsrWpc1QvC/kJljcntBHgbg7bRT1kMlAXhmYIwU1rjfn1Ahel
2dMIKwLr8w/BqFmIJaDc/foFejP/U17MENU6gB7YCYf6SYl+PSYxriqiRxRhAPIR
5B8/zLtzAGPIxlF8QBapNWATjN/aAP2LFjsC+4G7lFCqz/ZplH3c6Pxn/IMBYqV8
uzS/hqhSEdx97EnPhvWMV/i6tV6UQPZlO4Yy8VzB9vVjsppQq/BVW9q2dn2NB96L
q/8mxRt5cnoQuZZS/wsS9fB0cX92MUKYsuLe1zDzeacsXaa1J8jKjLaljYhGRqx1
BTeWmW7pMfKamF9R1iln5OZ5lcLTEVQljQk2z5hhkR0b5oEwlZAlBH/Ic5fTx5lr
T//chCE3RxxOeQ6lD6au5TaaNMboDxXmkW6wda/fho+9Q5MPG7DK+5I8MlrA3975
j3mViA6xUqHbmBRXeBziqz84XLwNXWoicCs4BzgzBpIYCKz5L2aocksLuyoBS+tM
1eC7gElBvYHbSWuYf4w64OB3u+qt+di13akzv0d5g9NKS2qYkyhYX6LGu3dcxDor
s6HIM7jFIxR/b5i35/UY3SCgj8O5jPOscgJa087+vUZJ7oXyCnFkaHPjXcJM04VP
rUenPOFEvnNI0obBUuNnufjXj+fa/SL4Vqs/yuSFGpzYoar7LdFuDw2dik1FSN/3
0BNMMvwYgHv3tUP6N2OOFXCiHiVnc65Nau2KXJB6xUwgQHuNwozzNAYJZxl9Acq+
LmLTzCqntXhgzG56D9qjil3ZhTlDebB7gi47d9nUqFLM6QeDhgxVQSrhVrZMPTGy
G7ZhfIfxgyge71FkGXeQXYa/chuLVKDEf8DBYduAz2d988taSmeAG+5DAy9I97Wl
qiRZt4mnNBeilt4AmZfU0cJoEw+yIPq289Y+SIxcjr0NtwzqmqshT0IAziFO8Z9k
ZOoH22P30MsgBkOMTKy2S41oKuHwdpBKJvoeZEYfX40XcWQBB7gthqYHsXiTtbv1
zWlOBedUx1MDYRGjphgP0m0h4T5ReRgH3SRwbdjrfelX3V69/2FjyuLbMtLV5FSO
4rf6b/x1F3rlUtdJs+KCqedgZkB7pxAOjxYag5WKU/JFDoczzbQv77+xIA0WgMb/
stvwK4fpEdqFt8qyU8ZezECiiYhZuKKYUAtrJg/+eRxTZkI0ljGjrFbFAcBGvN38
0/5xmCfLk0ncm4IFA9Gtkwy1XFjjDme2Mkr1Rfxe2zEzGQohRch9pDx0VItVXClj
hsbFTp+31pN0euFN/9Glvwacuc/hmeM8CJmQ7N18L7XI4kW5PjZejKTXiW/11Haq
lhfXGsW4MVTcJ88oNPy/KZwE+MCKsFMuBUZruoMepeso3HVe+Viagpcn9aaHLmp2
queNmYTMC8ttjRus9pMJgoodDigv7YiLvZZJ23mn6AhNfyGw6WuhTu5jvwccRuQT
ZLexjOBMTi1IYc3CpsCEB6hzwnXJ7aAWLwVbqfSbLdQRItLd+GbabqFCuAP2KTOV
BaB/6a8h4exr0HCg70iw7uNxiReM28aV1lcWDI6QthQS+zgsCg2LcoGcC2Dhfm8y
n1fXGdq66qrMFMkOhcW3vy37NP1rTu8BCdNFL9mr4BsQGEsOWo494UyfRch4cnSX
HTRyj59NR6e2T548qTi1bWNdOFLcCGi1V+/kgpLB/FRoGYxQhUFwg55Mh6EZI9gN
aZYSB0LzMJdGUR9+tLkziAmrucJhYI4B30N1Ti5fjLeC1JwtalibbCYmpnYHxKeM
zmQnCUHQTJB509HO3DviFBiP6Tf51NyIOP+g7jSVhaAOeh97mtjNZ6Hb/Hn5eA+w
miYRhIZ0W1ckHho0t5+5JOhy9ZiIKlDaAnxCNpH6an2vpjqVA5CkQOO8WjkHikVt
Sk8hZUSgyCEXGjFows+0clvVz2gG6iihjeqflyv8uIA5JVt4B3qR5fhAraAWUfyF
GibNU9pKJWgh9G6bLofnE86Anh7/ra/P0RzEVwEUN0NFqj97j8i5eCchypW8QhYg
nwJ2gCkMjD4RgN3O6WU1hzFKbro37+SQb3RT74bZ1uSqfnNSeeLIjJGhes35tGG8
+h5Yq5tglU49boFuCzEY13LUKgho0Gx7ige74rF9KUBPhdF/HFTST7hX0/8e6qlJ
niJ7vAPGvNOWHJmFlNMgZCbfjki2lZDr+TXNyo74JDif60xI9Wef0ZqSh0t+ktIQ
pITbEwN/p6VSuEqHUD3kKD+dQNVySXihFlYT2rWj5UFBvx2PznWPskURx6dcFOBX
Uv8OyGt6S5wO9eyriAEc5RbzXsKidt31kWTWxLb182r7DkzGhX88dJcqwrap2R2C
7IIKppBMhLlxto5K3EBT2qMBjsyY29n1U+S5BlJdpFgr4JI3fcFnqJQL6ZsL+LlD
dUH0u9vxG186DFivgLloAWzpG1nXq1e87Cduq15l5iK8vqxAh2G0x6BWH18cBmjO
MEZOe5PxxtiYL14CW/FVARTt0yRfgDmbuuuL78R7VVbwnELRnHc+C8fm3lB1Wcrs
PiwXILFEOTLNuF6YrIjQTaQRoOMHcBxKRCYDPc2oQsOoRh7sI6P96GhyOCObjou3
3bYiKqnGsMRHmPiUzlWGlGI7vwyarJiqIfmJy7FfxTzAkodCiiMOgCy60oCfR/qi
7k95p/H00Y+V39ZcsC5noNWUF+SKUkzEJsvIXURC9C/zmt7RtulgmtcgMGPS05cH
BQevX+qZsEcdBRuHe7kKPcfE7V+7Y83FnQDTBZkrd4dYl8yOdUiC+nPLUm6nyGah
H8Mtn80QxYLumWdz2ctNQMUrSg4oTjzGZ5Gav6Yv2j4oeRqO/t+IpI1NKQaYKFXj
SN0TPWkfEVTaKbCulIbsnIW9u77+hoPl5Q+Cigc0NE5X6JRjU2EZ+3Bk3W/i66eu
bfXcdCIuh1T4qvQi7XlBEHTmrceiAMjygXPQRkfxFLeFlnfyutCwcNNBSnTf0agz
Gco5SYWvq+14GkhsaxJqJeiGu3jonCHTCijPGlsG/lCprUvzc+VeBfuuCEIQKSGf
1oTWT+bOaJoEfhay1vpaaWjqw7BkftTxcqWKx4lMxlU6970zGfCQ6ECQDraqXdUb
2vxfrdHHIaNVACbZ++gqcCye21vJz2o9mRdEs2aygpUwnhIZ7M8sz6NIWyv9RnWs
wpnKp+ShwkSbHZzNy+hbfXnRMIJTxaZSmZZviX/bQr6TkNbDN9MYT8g8/NhPDuQO
dnVQUU1+5n5KVOEb8+ji69JXoOk/z/t2Pt63gwVvxCPbqtggZmF7AzMT8nMOJE9H
tLDhkKQhaMpdwTHdVaVhwISIgWJvsBaztCwAWH14jUJ3200Up2xgA/0JXimBedEb
H72Flhlim6l60oyXbys3u3KdqYUzs4ENPRSNbtdCGG3GP0afcKHB+PfoXADXSafZ
zg8PlpSB9hiizl9ENAr0tXaEI+xTxa0w+RVhl6P4OrR6wbJGq2JHwyka5DAlGMgG
dx7WjTxpT1RqhmhlrIirhx+91E8c1/SYlGoGMNG2wQZiIUoA+uV1I513n5FeDuU+
m7LYnS/gz003otvWlMSO3EPEMDlt4ARV2L5iyK62PpoE9ffGtOe9eVjFsORAfM33
ioqJl1vQVSHtZ7AxOI91dSoxWw5+hKM9NPNJQ/PG0xaYKNHeFgrWMEJoCUbVWAJj
n24/kl06Ka02bDRZrq5+/10DeJrc9EGqk6aNIL1yvfK5kn8d4YUewKqq8no4YwOt
GQeZC4VSlZZ0Tp2XK3a5Ec85pO/Y2/cDBGAKal/fYorBmtxsrInCRJpcGRmQycPp
w8nVSrScU/zp0vaJ98SsHj2f4b/7kiYERtFAYV4pM1Nt58f/ZX7KwEjaEyvmaPk9
rCh0uBY8cWr5f5d3HYKcTYELVOrW1A9DFJNedtP6WfRRSLffIqrHsCNiJQL2SaJv
qHLsZygD+yKikY6i0VbznMaeHR8Q2DfEBEMlQX47p3wn8JWQNHfgQi+tXM49KxeV
km6wHx9ORUaIn6HgtzJpXcq+ijvENBWa0/V8MprFkLx9Vb7tly5uV2Om8j1q0Ajq
MZ4EtDL/c7GTs0YqOcD0oQZB8YAL3U5rZBBbObNMuqJzlgkoCxKhr0L7lkcmqo5a
NW+Qn+yMb0XsmeEdYuik2eXU98q86l9FD7H+OpvdJINnRPdAewM0S+LYfqtiBxvC
dEVa1KVYEXL8jJxLpFZyE8coDTwdvUVpzlkxaa05ExX3aEprzw5i7QH3MceGIPAG
sd8D8CHykTdEMXljFS3ZgMdRKlL3h/et3zAJPKSQ/x4yLKupioQGYb8lCy6vTFRx
nEk7Yn+hTOSADcRwGSPLbSdYch74HWpEF+wHuSrQ10xwz8eY+i2fMAjkI1zglQPj
J5gXwuXCiS0UETnDfQWkDM1vKOITmkVHPFpvFlRwkT8xgAnFFe8IDwM5LU3N7Shs
EfNGjonSXkoMPVTQDZK8WiAWmxexqgf8F9137BDVKs5EtXxWqt5GuNqrUOvnxyYy
FBtB8rMcbk+M7g9okgWNS2NjqMpB2ZrH7y378aD1vagke+QLVaGrF1xu4u1UvKBS
uN+2R9w0b/pWlLFbXxg/mb604MeqtP/xcc+8XIhr6IF9h3hwHCnjC32fShvJJDrk
W01lTgCksk/+mviaV0SZykwRYTaU+yhh9zH/tejexkara5e6w+UpsJxuQXgPHBxo
obdrcI9IVNa+IpG7EmxUU/9yIAnq9o1ewQgbIn5xZnvU/KXKGMYPz32vJ6rpwqYq
bD7B0IUouWe+Qy6czsgzw4jBksPwD+l30wH+Ki8aQKFZUGeuIpOAuYLM6XiNs4t9
x5YO4ZbyE9gljARyoNbDOkrQhEBs4pQeuOr2NcXwsb8H7vJQrPcphj/lT6BpYAFC
EAvF+FlWb7thkV7oHJ3hME1WpizwXnI03BFUQIc694DojKJtNZN1cV7EqQ6w2u5k
SOEY/rZCxBOkcQvzA+01WFdv/dOE2E+fg3ipsaAkXpkRW9cxD79JKzRLvxRi8cql
FN0ihQVVN4w0VXmeiwhnNotx8IWzmB+zHDoh+LfKV5KVXG8ZrsIzk2zu9VO2kgfW
jUrPlsL/OzRix3OUU/RyYmiQTGX3jKu4K6Co9mnM+PMBJgG6Acwo2GPPTZoPryDt
uTs4SSMXY+TqmySttN5Sc4rIOo9opATcavPtihDEUvBmia7LEKzQT7tTQIxIBp2M
oMFKosBLPyPCCStQWYRYIke/zx1+i0Jbs50lnXgJBBDp4/onf2OtfiI3yAwNuC9N
yUzHPOUnOTcEjmOdC1J5Z7H5wGVcTADawaRpjeTcYhvfyPItO8IRLW5uJYPEXpsp
/d8avC6Ri396XmJsOh8x3AZOnyvIW4f6DTpYApvDn4k/2bgBI2D2aa7aCRPSiyTJ
EKUFhSJOY//BTXIiVGUZUFv1UGxL6M2/0utCzRGf5wSGqRBZCIpVMeBKI/sBocuR
bnAzn9h4kNtJTTUNTiI80McfwT19AIfOIkSu8o89mae8/cxtM5GDzURKF5SkWAP/
+JXNYX21vWHDhJ8E56VaI4/nxSXxqp+nP30H/IfFJoWvMQsFjYZ2q7zk4A7CzcJ3
GaY9T931H/pIjHuzzDqo5HpnT8ARWvol8vKjrTrcAJ6k94n8Gp3zOxEqUJuOsfyT
tRgaQQr1EgxgRFClUUIbKihK22puxMQAscB5CpRIj77CVb30Vg1KckTvLV3MaXLl
BkpUMCG2dpesO5OcVz3cPc6c6TPs3a2IErztXswYCcTA1iudP68m7O3Ym+8r4lAx
B77s4YIT8tTxACb34vcwH7lgsmTzd+yFQ3Xp7nitqkCCYwl7KHyzpkRqdfcGe0gy
xaBzvskV1i6kJusO0P7r0W18NCe1hn9JqbDHzzS456bd/BNmfWzf2i5QdAU0fQm+
g94M7I2BwA7RN2I5xlqM9WemoDaRAON56m/exYeesEWiWLGQhuDWtQtDnPqGH8jq
Oe1M0OmwE63ChpGCbhcJpFt7Y80LMvEixoMKcEDezO9JTYwKNqtNjlVBT34rXWu6
nHgz6u1fOb4vuNTzJ4QbkcAPXYqF81PPr/SL+M/pl4IhGPmuDOnhnfZvguxb0kDY
QwmCy9NKiRl4ZyTCbJ9HB69x7L504hu9xO0OCYSh+pcZjDRyZ+D/nB6g3DLU9jsF
oUS2wnBHD+HfpgLz5crxyDlw1YWG06JAwN15d0fbi6cBMK7ErHr6Yi4+meucPkGn
YE0PV0cQcFrc2k+pWmbaG2AVJpqjNnQnDZGr7XBg2hy214KB/H3VTjEO1/K/ZMST
Xqa+aUrALloDRvzI+v24uBVPtR8HgJWRNaX4rWJItQQS+88AR0sfefR9H8BewE+/
SlcmkVDpqzs3w8dbZa6rB89n2Wlb4JM4n+5oHU8Ib3JEulOktAFZfzQzUPkAZ8F5
vcTFOJMvDAP0M3QA+VuzZ+OecCmfaXi6xfeBU5ULUkKhp/YHwNmWmz8tHFB/Umml
LDQ8JAs5dpnax0A3QCwQUNoKHep2ebKYe5wf+GpHZhZjZQpvFTi0vK4xAVhcePJQ
QqSn0TwePzYmaak1lsASI8MVuGqn7NkI3+GL2BujhFSD683CaaYMc598AhdkEbOk
gl4Bvjd2LIo7Do0KtTbQ0Hry/mvBMDbzC3nml9RdzDeWw7JwStMRSO10njR5CySS
8gJ+7myrzDiGTYJKupdYBSHiCxnEGAD95fMbX2QMnqYgov5eKe5jk9rSoqnTPCqp
AloDa+tstOfUXIORrZr0xnTtZiByUDpZi5yq2l8drVD2QpL0L5U9jDr6U7Liizhx
nuktOtW0o84OiUy2W40XxDBr/mymRNLq1VPrA0tDon+wiNWT4xVN9HAe1CzCGwOu
CthKM57pgkMOIlLB0t3jd3gc/8kqevoNQlcL3CRRJvBkhJmAL3SJ2iPfzuei3w4K
jGohHhzvqWkV6WJ/Z0WMhOR/xWjSUMzeqDs3MSeTw79KBMUIZIWLgjs2evZl1rbh
YSR7BMoenjAeIrvbizZE2nUK7bbc8K58eWDhpXPuSiPMuRS5ePaFBpeRBIpoLwxg
cbLgYRFp637aKVTr7TM2W+qbIeT9Q8XThtwSo9OkEvQ959d/81t2YMdBut/dAdzd
GadlRkwiOONYkN+me72WT92P2rXyXZZdn6dHyCbKFINkl7E4S4Je8t07w5NbRUw6
h5fxHFzIa/n9Mis1O5HymD++DkTte7elczZbt0V8IH4QDxJMjoOWVNIq+NpqidLR
ymy70p9o/lQG8HpOkrhyHzUvYRlaydGnde6n8PqAMwDznlO9Egb2hRwptzOoE+ba
rb+o9eI1RG16z0tQiIbjftMRxpW+gnLD+8/6LbCEbdQKXKpEF7XwETj+tOkFWDhd
xkpnMge4wbgBkMGMClv5TVc5KAhfZFeKzQ1k8FvBMGTR3Uvpw2wfw0U2kI9uG2Pu
AUPQY00WdanteOOE/AOZCW+vZv7aoUAuqQDNICVEdeMDqOSxB72LZwWahWdJ23dx
thjEDs9rMlZ6hEOkWFDS7hqA7/1hVyiGJVOBJ2TpxxOW7kXkXP4pavB2OVCO4Fg2
429eYEUvhoiKswxUxC622ojhtXFsAqzbIz87u2Dm6yv5obNspkE4tRgaDMO21UiJ
g8zkD9fwpXbV+uIMLiVxf5XFBuPmEVBIpGNB1rqsyQjBJy+d5EHu5CRlvqcK5RI6
ewneI/dNnNkBe0KXnVHqX8JZ/vPhOwZlEcIxa+USwQQwfkQIrvgMMdz2VKQ5ee85
aj0Ni391oIlsDH/FJxM/Wi3Er8PUT2NBVFEnMy99GhwLJOwhcagi/aGejpKVJP4x
m2Ftc6pFuILNVqybeKYBPLVyPu38Qyrbm7UKxIwiTjFTQBrTp/QyJLj6iFUN5+Le
3nCNhfSMIn6fBEH5afZ6OuCuMZ0lqx/BMZy2ZQz56AuIaMbsF0bbBowjtF5a2s76
oFErmmgUoDIFsuP7f2u1YdAJVRnycbI4M4n3p06+mMqbcVJ5B+2tMf0QXUQulX2C
O74+KWdo7oAqOzTjYUiaKxDEmn5A0GOrJjJ/mqZt+yDnT9yf+4iK3eyP5LeMfeA2
a7V2vtjnu+ot08auqwA6jQ5Y0pnWvK0vKXAE5x9JdndjPb4J3gFE8IiBPpegUIlm
y6haTrWhJKS7pJBjQcKnJPGwueoyVZSiqGFqSC03PQbwOx84qJWzc+9kxgiofLW/
sHmNr4AsKVzJSmwvkWi6nsLRqD+nfwnS3BAJCYdhreFLbtkWXHch0IWcj6iyekbN
nATR9dXqFPMZJUi4A+nMht+CbfMOpVytlI/Kvpa8p+popHOgyGRk6oTGIamu6/Kk
U9Mc+R5yzAFUjZkC8mwfuW/sqNVCmUb4XTxjjfsUBuOg/ZjHDWpnTkuxCPO6SvnB
zR70YuxjcNPaTEjXa2qJlTTgd2PVORbchMzzeOa/VeUrcLonQsN94qag6Qe6jXzb
mdW0h29rX98HItMzaeG/6j/z4ucb3jBRa0cJERtQx0DbQ7qt8wGKq07XYcEzbo8C
DCid8XreM93wRNvJ1ItkwrrXmi4nZGk4/ZZXc7zHicLIf21U2wjQ/agsHh/7110Q
o+aZeNq2/18+uJolC99BzP7GIsdC7AMl/J8RNKTemOoxI576Up8TrZ8eC7NFlNwV
zXD7xb3wSsVUs3Zht+ZmUV9vfW7wIYbNEie0RC3cEf4sG0+kpy+rkIxZHcwYq4oK
1ipVfKETth0+FWk/vOkd8vlA1BdB3Z9bKhpFUfmcS7VTxWTt932kH+GEcZEDoRUn
xmDnh6lYGeEPxWkhV5REPh1KcilVPTQDrEynUwe/zoxG4YOBZC2VnV/FJFMk5UOB
ZWwTo+eFxGCkqDA68Gs9hPnMT6J7gs3J1GM3o0TU24An37kF62q23gyf4dEMCdAW
4nT3IdOrUnhv8BV1xBEFyKwuhZefjvAyDqJ+UDNS6LhDIDmyexz6wOlHq9UsUFE9
v3XgzBMhXzlARanPJUIdVElRNG4ti+xZdr542R2T0bIH9QjmKSTogMSglRAt665T
bbh4NcXm5slCaUoKPAWGNdAsCI9Ch6DayQkNkZBrqRtbOdRLtFyx67/Lc/x97mqj
kM5m2FieSdlfY+jGm5nLXl/x90WgfFq/MFM4wAzEw6B742HlBRNyhGWIonxMTCRX
qhb0bMVJ0dwr59QWRwWDPV1j1oRpvAZCNXq8ONjIn2x7Cbpi0E0X07CWJNlhzKSO
Sd/nUFXMhIQwWTKDXQBOZn9NP0fFfltKQgpgYdQCTf5eYHVe5Ny3Y2GEttGQ1ebd
h4GWa54UzXAiDYwhFEhJaHU4dvhk1OIUBpBT0BiItiIvnSGfz46BLUC3nOD/Ulbv
+qYvq7eOMw4KFkxsb9Rvzq4Smk6MkFP+kyszdx1YverC35voyGktBy3QgOD8b15F
w9eqzfq8zt5KAJKwTeJOB664bh4jSC+vurzS0ZUc82u6gPCQHBTonLCEFbexSHh3
JCwfADb9mfzv/A/TEAawjsEw9Po3LnQNgnG7DCmPIoukwOdYDixhQ0MSgfov0KuP
sL+OA97IiNokKOms1RjlBKi1PdRjmWhiE/rhjq+XGVDAidfv8ZqDVG0uFKDnsJ2R
vgXRNXy1H+cusAJhnecuxwueSUUbska+2vSMiP9il4qkWa1PWCPfSrkcP+vgIg4r
f9kQZyUUyND57s4Sx8Sj+xLZLfHItaz/2LEm27oa/AdFWURWN5Y3OCRrQvVrkyND
SJiWJMm1QmLyjiFdc7bWRrcDRzKQZj2QPl1/w3et3aymvyvI/LNMvnLZlpLHDMXJ
uyZvtmnzEctNMFO3hk20/LhnVSsV+ByscY/EFSRo0/Cccs9y5qDlzS2glqbVND2Q
o01rMR3pEj8Wg791PAqQGr4q0pVH9qCHshc5W6kTF66DCgItV7NDj9o+6p8QGIlz
PUuAoi3T8Sk80z8/M0x0GRr3SArJ1y/3R1WTeiPUB1QvmRVFhHnpRczmn0dYGy9y
SMELhjOH77cVroXVT8xFlGD9pgqqhGUEF1dZEqJS4hVN1/wpuX4YUQS04mzEkpSo
G/xjE2BoWmmo2fTN6j8ILtU5akg8ygXJ4EPGScCPUCngaD0rNKGSTNcS9AoWIz5b
1QjikDCh/b2/cCwbRo1fEWRSnos21LmgkehThzW9J4GsylzxrpnjUx+QrHDy1QUU
d2K9Yju0hgIUJMbZG1z0OC9krsk8NdQQj/OAxuRihpjbD1q4jLy7+y8sg7z7uOAN
SfMkWnNMDKRhPt+mZ3dfEPd1Db9ThKW2e+WFtEX/PiL+zqtGokPMoNpdn9Ge9r9d
FfDoitcFf+19GWoPQbqpPeCj3GPFZKeV97gSgK6jnDIBTR+UpZi7m1hdUhmfOvWR
zb4I/3qP4qDt/bMzsazuGHMEYbtqZz34Zya4m6JT632E8/04BJ8jUjJLhd8NdN1z
YoXRxQHOnU8QCU7+rETKXFsybQmpnaEw5TqsAVLpFg3ethc1H4hnleZcqY3JcouS
MHIBa3Y40IhNRhFDMuYTuvgjWL82A6ByDy3reWyZhcmMUbFyPW8X0jMt0EPXN2jp
RIZIUlYjRl+CZqBBPTLJsW9dM503IGvlI+tZoeC5imERnoZoHxJvVNd50Pda+fGn
TSd4ykCi0S1wzrdWCLcQFPOt1Ao/s+nJszl7yqfSKQxPSe3GFg8HPj7sZGutTvzS
CJOxAWE6JKDUQ0zrfx0Bo08ONDCS6XK36d1HE2e5inhVRFF5pJSK75NwxvgSpZor
bynkDOLkahGcxH5mjJrm4Nptv7q1tycBIR/cG2vT20OSqIEUNhgOHikGsa8V2dr/
wu97c8jMQnB6XsjfmDKPPB42eFQJ5AK/oSNp9WZ6rDdAr1Krnj8JBHORbfmsBKLl
nOUnZfJZeqw1hiMnNzKMQ/yBAVtF+ZXlpIRNkHSECcNnIIovSQW4M681FOEiEHV6
4kK4lqXx4jNZVjIpjb8cnGYRl3is3xkjVfKMFNWWobg5vMbG59M4js8db5Fi8lDu
CFXV0HtD4WEENt6IuPgJyG66HGSNZObRt/R40NHU09p8oDtYjJGQdWbIJS5awkp5
xkfBiRtdf4rYkF+wAGitBFcc79Hy6B7mUXZWgHgS+ECIrTMvPXdxEkuuc/O33OV+
dcbA7+A+4RBUW0ONDiV3k9SCRglYraYF+c3DaKQFWWVWhVefDP4whGozDTJQyDSW
poq1f4DHh+n921iatu8WM86DR1cw3Mm3IEEt4jbr/81BY9IVc3aGgYPFn52IMaNM
rtCFQTdjjxyp7jy0IFKTveXFivSfxn6EkfhuN/4+gBIeoI0pzT6vTJyGLUW1lhtt
x1k/ZUyl2T8I85WhJUhFDTanygk6ww+ntY1YMmwXI6Qbds/ibGLe6f+jYTthWVIx
S+xBo0sk3qmLAQ5FuJvilVZdxqJsKXJh+lVVKJwRSNZn31EqhJUIsmuKw5ph04wG
wuxysGvsRgaZQmqzm+AY6YNs4WoNs60IQh1vPT7iz5/UdQBnp9j6yuVKGg2XvLuH
qbKZkxv+gFEumvM2RNJ02o/durgOn3bU6wlJwd5iWrT5LmSKc/e/ZVpOovFQSltX
v5CiQco6pWoC0v9O3gUGLhgeqePxacERKm//mqOV7WeE0/5ATLj0hklFQaft+3Zj
/dWC0x/5ryrTqNjJefwOFgQ/1Z0RzClmleY9NmY5CigKovIE895Plv4hbEOkI2ro
2RSzZlUTM4BKZbMnLmqJiWt1myck8v8w4irEZ5UPVtiwKcJenTdhmAaWaw5xsW9y
k7mGtASH19ftDWJaozJJuh2BELJZZSoDNloisAaxCW+eJmrrYyJb5mLPJZ83nEx/
0pNERgWFFfJBSpLmIWgCNU7H2b8dPGMI94vjmSL+Evrhaw5Y4uf7TncwM9uDjQcR
zt1a/0ut7TBMetpPNfQw6YnZQLOsr5iJ4VkhwZ3B1025qrorrtC9gYBXHiVuG8rU
MGHc3ZhR1830dk32c02ceJeR9ImqSAYPns2utcY2gdEVGhDO82OTd5pnuFYy8Uxb
988W4d3hxKFyU9mO/T02zI1hDNH5JeFz8SUjnRc5hKv/cxn5+nnI6/uyTzl6Cxm0
CSqCXWLGAh1fu4vKedkVoiweO2bnJc3liLNHAvXMnhsj4LOsdq+JktLTYNm2YBij
vzIlhD3CLvIP8JIqmc/gTJ3wKejqu57XfRIPDTASIebJ9HTL3oQyFavQG0v+glUd
aEtTXr1xRxGUsTOtOhoUu1Sx7NoieiHiFUyFig/9MI697fpxZWiREC0syGyB+VJJ
OUoc9aBP8Ugrgpep4zFQSEU02x19vYqZHY6MH3XFqkdM6W3CCrQwmjPQlTXdlf1E
BvwUDbKCOEqKu7T13sjioO8JM7vGQMv710HPXX5zKxffloRBEs4p5IscwoN8uYxv
/GDlykAVLMha4UaK1ryjNBMM7S+x5m8mlzi45WC2i/g/rOCiQ23x72TKM4sLErpx
WwJxT4hEjXU07Xf8QJLQGItNJ9Va4VqSgPxqNGj/bJ62CHqIVWVWjdTrYgtazRmB
4lgS9cukNCe/tn6vHykateD+LBXFXxGn5TSE6jiY3uuc+02rSgg2y9B23pk0qogK
1n0bU/P2NhuPiGrPUGK82G91smVjDf8XCFY8Fd/SCCQHOtS9f4NnyTyU2QNx3Ph7
4VYc0ZY4bd4bi0Inxn6h4zGm5sVaZ1bcBvDcQNDcJ7bC6OeAfhOOED9lNDRJ4XoV
ZuGOrPhFwmnPomHCmf58G9qtrpsIDHsh3uQ9fkZEqKKKECdomHpf4TeBlp7YNXbn
vnJOFo5XJXbMnjTjVVk8gYmn6fIaAydiy7TaG48g+1IKybvikfD8VNLjF6LlsbPP
rm9fT9bv7noYLlo7iN5JDOgZ4uETMUtJD2+R/VH3cIt/zGS4puJ6KWTp8dWB8YcY
Ek/pyE9SLqICFx5gwqJ0WpTGHgHf2ODzegpZ5D5TzxYVdFN3uk3ExNYtg+ZUjG+R
eehMELVZnXjtZNmsP9e8rjH8L2qT+DEVTBqsCiMpEppGnhrYfzymuWJMJG2BbXGI
w7ZScPpPwhzIvX0CTK2AbkWkmzqVnbxcZ2llYM8a8K/nsbzJ/WQEP6Khkcb54DPp
atmVQN+x/UG+kmQMkOUXqqEHUngmmHg+cBxnGayBmdfm0IDCSfcUWVXwyaxgQgGN
ac2tx3gNGpPs873pSm9H61k1qCvGbuKfLRa8NFLIcBIcn7ObI82rKg6zBOxmqRe9
6Wut/m+eV8SBXQ6HazIQ+kv+geLIiLhZxlzhf92JjPXu3yDJ9UMLOX9vPlGMp8Sp
DPUrXRXGWAdZRSrSM0lEDnd737BgP094EAH2VEEFhnEvMLlazjl9tUlNXoFa84J6
B1ApHjvTlLenGeWsyL+uG/qzdcHAl77mJnS7K1OdWgCExCp2eiqQjNFK5nyS4kGH
T6FONz1bn4BoIHJdAdlTmGHUIheZ8RBwDi5Q+vSSGEvUgRVuTA5LCFLzGT+sxXeo
i2NHTlp/dWFDkxx1ZRkvIdobV7NIU/mn7vv/6fBeqjJer3GkgVrG50YkwyrBemfe
2Rg2QcwZsPI+Xe/5dDzGXWPtaD260L7gXbJvU36WI/IbmqUfu1r1Kaha591HQ2mK
JE51n/KmNA7UsSq7uY0wMqrdan7b9RB33+2x+mbaKTwzDTztqXJbNUG00+6d6Rgs
w+XOUsPSOhKdTNdlk4SVgyIGgsDPZmlC+RsA4jJCkpqMv938KOJd0+kdxTNKzD4f
DGFC7oMaoAIWwj0Jte/k9sk3ZISUh5/m9koXkzMtBmDL9afaD00gjoNYOeuGLsgp
C9BmQE8YiMqyQxqu95W0yTQ3MReX56OyWBkA0In2PdwucEBS263R0cBBzO/bG4AE
1W6m14SC4qyIUIMU8CEk4qO3/7llQdqi5VkK9N5xXcts+LhsUX+e0nilZAMW5lZw
9Pb71SWfEATYD1hDowCQ/lFtwea89uF+WHgPzFWz84t6LCj+cHiaXc1eTQbMCisZ
GgFH061kloBOTFUhy1jUlWhknSJgaPC0h856wEF8aH7LAq9twuxY9VR4joIe1839
omjca7Cf6RI5GrfIxOtRXyoxAoEVGYfenUr2LRLHWXnfRs5LZScPirI/R6iM7+uD
unfeHDMAAWLVvWCT0yt2xmf8YuwhQdgP/7P65mHxBoGG5Ddb+hQr4aRG435Vvrwi
NzZa05/cAz5LlRMUGL4LcnAzbyhW6lDF8oRGmp58UTm9+8vf88adfuZDK+dxQmDJ
CMZWSwBJ01tamQhkxB1zVoIqIqGdeLA56LJS9OtQI/ylxN3TkuWxA7fbEe/f8elC
tWmgYBPmmvrsXL9YatDuHa0sA1AmGtF5Sy3gX2upiw4J6xH5dM1HCt+ez/Rv2q3i
nzgWkshlbEODAgyhU9ym9sXLHbZhmFqWL1q0K4SagyD9fCaYbSu88aM3m+zp763/
VYRE2z37zbDYx/a6sZ2+ahkA2O/jBAzmeVdPlk8wDACOo44TTueBEnJBsBZbBk9b
PeqSlOZWS3IVIkPlw6q2+ueSzkVJRTvOilIdLnECDHH9r0XSKVfMGft2MjaPWQ+d
wws58KFrTOemBzFNPGkCjikvcza3yoPaVzgFmBQDHkiJchpl+vZn6UuarWqLmRtm
H6bCTZy6vm3LKXhG110bL6sWPl1wx+mSSB+N72rs7J1HYRdtQlKicVZA5OExdQxV
zFck4GWqBT6Sv0UQ5FcSgWVtE1PU9ntdRdYQ9/PJ687gRNxlc9vz8SsGssKSx8M+
JEvhaQGxjM7bg/zA9axrDjiHxxfYnaB+k2FyHLhuW4EdxeNh8S/S92zk2DE8si8C
qNEBqa7wgAsZbd+qJ2YVNvar9M9ddXhrxA4pjigIwYfLQjM2mBm73Ii2fMtb7QwL
2v/ZGHC1rKG/lN70frsBPW64z7yDXOTEFSkrVhFFJpVGK0Vd3xoQqGqbmhQRnX4J
w2X/+XNfSgLc8rRiJgr3QMT83z4PpPvK8KatMBjFIPflGMeyX16obBMpspvBS30r
NzGllAdiaA4ew92sFNzqfNf4kF5zv6G2g/zzY5b75B7fRHf3A9svSzcWFS+N/Ye+
ZzFOzl6rY1+XDbL44E3V9SUha7s/vUJYEktsdyFhB+ffg24SAGwv2WpE1MpSohbO
tdLz9J+ASzcF4TsaIOqlptoT883sCSL6byiaQUeDwC9BQ35QwZ7ERpAuULSLQoIW
n117UAO1MNq8Wt/42+LUwDVXNFLf7Lix5L9ce1m9Wutc0Pght2LYIQTZUz1pn8V5
ikJpc+FdfAPaJrdTWNV/h/9ro3picFCgrCcoWE2T46ON0BEraa/Ltcgq/MHcVpKa
AsQD+tKrWWbxW+74k3B8CcLj6eXernB0rW8XGYx7mnoispLdEIqG5rvraP7Igaq3
0e9kWB0EKxCmkMW2anhurGIblkIioH1LChsyosoIWBzRxXJGwPQ+pjAe2PqpgA3N
6I1OqWxXmGr16gRv6VOOq9A1UFNbKUEquLug5TlOHc8i17lsmybvwVyEySkNv3HW
NWiCx0W+vRfMKn/h43C3yQVc9lbOhPlbFDKAcCGl5UBK68AwUuLd3zT45XSamKEV
9V8i3j5GvG6gywN5NkBI+tin3VqfMQH4kt2wykMWZgpD9tYWKQM/9RYBzgVAC6WC
lB1SWLNwsqwplZqPH0hAPoaK09jsOfRn3s7tyZ+iEDgYb8L8/l5+cJxFPoAz+Ldm
86PcLIVTnY1YCJAay9QXthE4jNUYnZ3jePT1GlG0f9X5t3qY6+VGgF6QWSktgNrr
o83drzRdCWGT8M1xokk5A/255S+tJTJZ07j6xUllOuheKG88M8WkIW4m6tC2Dnof
R5I97X70VNthA6SLgIAAELkaxcLMlhhqfu1LrM1Bn6JFi8SqNIbWgq1QYDJ/1g1c
kWqOWRGLOAEDdySTn3qXqj/BtUPqePalmr3eXBrudQuFIOSfylpGpo+8gNMrYmpr
1B/hMVC/pMOp/rQxJOf4NPSoySE8L2380Gc61rWTs003+8i2LRGxLy27FkLy/NWe
IE69znmIlmdtHYL6FDYWMQSjY3T53qSVo3g/9aM7efHa6MjlLuDFy6bU2z67bX68
BHq6Bgh+KCYgpfXSntMSK09ASklwK+ML78BQCtskBoaHyuSRRZweIhhbLPXT+0bw
XGNHyXjP84XbujqqflkGllHx/RDebbRJSlUJGPEsbZurFGy7vzeC1EN9MDz1CYcy
iTCeTtpG+0aqAigoKzJqE6AV/20P+ZoIs3+WT9Aypze61f64gLraW+yAgHCOzUzK
fKYxxpH0gIGHKmq4y3iSIJFsJpTe/r8RiitDAgeawjmt9hx24o76onnfShDMVslV
fLCrc9mptrJlLMM0ykzWm22j8vT1puy5Qvhb32+753SC4NuqOUsotYoogJLuiYDH
7X8RaNNbaaUTc/NngY5rGkBX4MZQn3NSoBIUDF0K7hwekRMdzwxoKwtit+aJhj1s
TWFfdXodFI03HdK8Kqz3wFRjYct/bJ/UWvSHucuYXYbNRSZEn0Rube0fJuhtvJCu
X+XA5tR3DtgF1DOq9f97dJnSgp+hdZasSjJgDV/fbVVT4bYBTcrRy9EXN6P5rXCQ
TxTFV6WLKl8M+WHzcGfosmv5pkImWqS2KnnfnUdvFt4Y/+SL7DuogJ0iym1ygf+M
/iF7oLj+bDgDFlM7je1aqMmI3GGgrVOwrY1d6173L+pig45npxoaDL/HSjf34QVt
CerXHIM9UYtE14jy42aRIOn+VUAJB71Qsu7Xd7wCTlXD8sMac6IepxuQyJGzarzS
i8u7oEj4ov+cu4hq3WtDLsrCuiPm2E4g/5LOBycJfQSE+2aD/nrwWjT5H9keWjLR
UOToXHNiTASHh+pi3giSw133Y2wPoTCaM+ZVG5IjVkNAbgceCeAbRx2oRah6JuAf
oGTTZ/ejcZx4XHZ18uIa4vNsLlFT4kxAOQ7JPiKO/CP684fkLtkzVYg0jbOqHlpM
h1kfCfzMw/5QUt59O3R33X3Wm+kbI2YYQ0DCWzm+ICZWsDwNTKys1kGmsEdNbaZ8
wLXjhoBYG8M7E/ZrIbtCtsqAiUAe4frzAGOsw2RmHUtirHyWRBgK5ttQCkKU/0i9
PRqf+9ypYpe1pFhLDbYfGhbZr98caKCCAO58j5pNgkZqQ1nnvj9Bz+j7uh7R4xvR
fqsT5gZUfiEugz6Re3sByeLo0hyzuvZ7nEymGBhcYQ8/B1RezVBtbwonfLJrmJRj
1wYIVln+qGCuE2c0HNAkcQlRnaFLrgVCBdQVLCbIxcL+xmE6ejUNUQ8xiqS4YU+F
WO1S8MArHXjTrYP0t8bIz58hFaDbBvKTyJpkZT9n2X2MPmsSEkFP2UjgQ/PyM6uF
pCTxC4OechHcgr5AMtP7PRpjBpAyMplorMKu9BBKZEX69u/Y9ft8Yvkj7m2Tb27V
30xXGHwnx01wTw68MwNEX5jPA5ADgXG8fyT01YNdQLYj0ASroamBycAqbTMbsz82
6EzxgDiHGZpiVTX7hu8cAZzkDc1p+TFyrdq6AG0vp1hDK3rCuFOKFo4/XG+jW3KW
iuWq/FuFEldPUm1WF62sfJhzMFK2cz7vSyn+uT139yFUZsAbFfQy14VQHaoA0jYW
rSwJ+kBo7m2AadJ3u1xBlh6dcfffvHSNmTy323yQJBW0/W+vwbKYWwyJdFU/L+3y
1mUdUv1mPuDxncLaDq9l77UkXzCue0WbuNSPX1x/QclorJ3pyn8ezcu1JVN1QTQn
jImcI0RIaWUQZsL4+F2HSSCGkDpiY0lvDMpLmnhzDBvLgVzJngfr3mtBpRZB8BnN
ZBGWhHpr0xPC3V/utgAY+W/9kjPDv+64TvRC5zrKLYYBJ8hvB3DY6Cc06UZnykWm
HyxfN9Dev3TxtnWbyoVp9QRFIesmR4EG6zue8fB9sMos9E4mSEuNEz0tHwpfUa89
BjAjuBARCY+sm6DzBuWdeoXBdhcifz6LBq9Wrny2A779IvYACwF1YC4LX0X/KvoS
X7W85+E5ngQSMyHsN+EUr08FRrGAqkV9WxerUt+oPiAKpZyzEPO46Qfdasmatmpq
IRFJtoX2Qw+FjcyqLiRNqFIDEeUDowzbVWRrojTyDb2Wdw4TVHCIqloWr2uncLhY
VGlmHg7nVlSyXJSz4pnrsPFgSalCKwqX/0LtRJGXC/VzOdDM/Z3ZqTSkOQRnGfxS
FX8OuzfEuv97RPqHGPOPqLZSfb4P9goWOmrCN8D035mf7euNl7sPn1rcCHTdz7yq
qm6u2LwYwza3zWpSxGI3COjWdGyED8z7LY09/sTJbnJlhRpfR1Xh3MRsOqAk06et
38j8U8mqemRDEmTybdzuWw0/jMzyg7pBaZke6/NxFoIK4zj36gj7mC+dzjwkGG7s
sTMmXalXGHutggxt5dFhDV7KRlx92eKYrFWOfTSrPdsNpZQYVjOB4/Vd8pEe++Se
nOAst4rq6in4I6VgNM2DeDMh6+yftmFW5EIs2AgVFrFmJP1jq8wgOmYHJpc5CYy1
pWU5v5/sW7bzrzsDqpxQkJxmZVwjUjjYxnJ9NTLTc/AK2uAk1pwlKcHrdaxkeIWk
Dal//S+oc9HYeys0KzLGFoGKvlFvWf0u9L/uubZfcD0zxL5rde1mjr1+qmm5K3Cf
gklpXy+Tnu1aMkBr9VAGu/sSYzP7AEPAAvWqA+kJX1zPR+P6jYaQap2oVH8bHzuG
DlxvX/aV/Ilg59E3iDLFVB1f3DJ0TgIOarguwfmAiyc5X5PlTpkS/mp6sR6Jmesw
63BLit1WkS/yyZGa+k2swQzgL30rfQjWaXgMgMidmUFAoVlqkmDmJSGNf6r+5ha2
4uf6iFYMIWAo0deIuB1u7WYgT8nmUbn71AtCOV9eQikJAnmiAd7otR0CFzb/vUvJ
bL1ECyBeY07DCtLHUGPNNsQHY+zg35dH9+Z96KI0DlBTLo9oYrN25La/aGMxQCah
uBLDCLfbAHery+JI3cYsMVkkRBoHzLAn+T8xvtP5j/2FtRZzMFCFr/WI+wTnBHOl
Abfm+IFMJy+unPMwyOkVqIpOyhhUjfjN5pcj44195jNz39c9g2AeWIvmnd2l5XsG
LoL/r11olkauWrGy2dw9pXNfKgLpg4Q7/eeerEllhEe0Ep+JnebB1f4Ryys/nTsN
BohepbpeKK0KrmXuSnC/RriyIAFBeLzpV1D/IEGb/kUoppHdJPUlX7d97fzOjuZl
HfW6r2b/UjBln0fL0inLiYOOryICN9NjX14m+/ttZGGAeHKFak7ouhr8lhALNc1n
PsUnKBY6laz019EvMwr+uu4eH9L8lTEZ1Iwb58nVhITtPjevMwe/U07Bs/3mKQN6
vKmj/Y+Doq8wbNu5lLkaA6wP4HLLoKONFzZCmf8rOZ5/BhmHfizKOr7gcxy1ErB1
ViP/MCiHTxESmCoW9bjSq1GbFAZvaKZS/HyAQCjM6Px4UbQ8pIOLSXOfw/SDNlSp
UvF34AtmUPMGiILYMUk9G0TtZKqqiGOC2KHwn8uIhNiyDkh1uKGNvxjQKbUa8oAs
YOMJa3FxI7JKKPWcC8gHClcjQ+B4zelUApJpm0iRpR5caMo08sen4h8/7RT9x+Xz
PdhdT8qjo+qFZOGJ4+36/GKDLTnETqIgN5tDEa9fKBPy0JI5hgDqELaFQAFKRmk5
Y6yYVMsVVVxV9/zSeOPeLoCc13906NgYr5SHk/Swx7FIRb42wJfFVKovocEWpLb3
+hem1g0Mf0ryItwnTYDXFdxEWdpIWcxcdK2MO3iW6uosy+OF8pk7q1BfXUnAQMM9
WEJLCNkfvVVh7XxhM1JMPEgCr5IoSfBTXmk+hte1KekKbyLkj63d/QarCVwqCGA4
nfaOnKg0RnHeJDo8W2+j/ffm2eot13B9c+U/r0/v/GtjA+QpAGGQ3vyvAxcXII1f
jUf6+3tELEyIVkZTrBlCJVrq8neL06/2/zvmCPjEsdgC8vgT4ETCJKm6QmHPKkqh
c3VEVQFEzYFXLJxrFfVK/xM7D33ReTkUVd8W1qHXfNnwG7JzBTQe+h5I6l9T8rQQ
TmjRkV1Ccv7qFsn3rZy9wBiTF9L+kKzgvzNVVCbZfw2wHDIKG/+HZXogY5GhtMI5
m0QB08GysmnRMjPdAk2v5UJiQLpldejaPJg1qvK+Ynn/cuJsX+Wxbp3wJvyEjWzD
ZYw4UOY4r7Vio7n8VrnWWL2V0Yx0UN2SnlCCOUaxYR03v8BtsijUVUMrlDQlM54p
R8tJ5jh+kxYGUVDldDmfzP7y0blG7Wd997EgK1DCuofXnGfuWo/99R/BFvObked/
y5cvAU3X/3qzQ4DmXsswlCdhxeYX2l014J29mhLwFvXI2Z/LWSy1jQefzfnLCKDY
5SM3NWsPzYR/rSrqtztNC6O9pfI2DgN8mu4i+7x9A6779QN/8NjJkoq7UugV/tHh
+yXKjdpkY2zqImWbUQwc7kZjMAbEre2VRgK59dGqzD6oKS3wJFbu2GO/O6BHTTAm
Mawuco8mpw9BehDaNhNO1oYEZ/7uNa/UZ36yEcyUvrn5k2dnnskAYHPQqHLG56LK
bS4D1KRccTyO4372j/Qn8Ksd9/0S8XgU0ukH3/bhLJAPRi3bmLafmAu1Su83NS2S
2TAPrG7OvEEM0uchmYqoF83RbMA88EWPV1KGl9GHOLrXsAP8gjDGUeMQhmnQ4mJ5
nlOYYt+Iap3LsfJklSC8H4qnU+WSLHPEdonCk1x1VTVkc65QXTc8GdNkuY+xCAgh
PD+vpDXC3mZDyd9g2VvHEzLYL46ckYk0ab63IqKT/oh6Xnq0mVOy86O8Bo6jB4e0
75rZSYugta1UCU/LcxSu69aHDVBX3F5xIiD28D1P7VZdr1UpIw3laM9s26AoahLr
Ask5yDhsBHBN2EvlFUD/oZcPRktf+q/saGN1w2jYx8cYBXTH284mrvN17Ga6U/Ot
TtkDWr1u6U1k6hysSu4rbdwYabLyQQMiySzc5OXIXfI79WR1Qr7+eCSeJ1KEho44
pVr1Y9VC/lb4DDDblLXZ/fg4b2oLzcD3qHOxF3gJA2IOvli23J8bf2eP5Qb/66Qk
VhUMa2kVxX+W2xFRvG+C4Jei+WWWCnYv+WA9JdLVqPsX5l8qOfNWqFPOKdWojtLQ
1jytK+bYANXs0/HW7x5B5HeIsHF5GbUCBXdfnZkivW01is5MozOFgU6OEq317bBz
u+ev8TjEiFpRIqiWYIRxlT9Hs8ydHgC17CjFldxZBDgaNIxSIA1a8NA/aA7j7Dlu
gmd1QJdSlJGuodqAqDuvvTOTivv7stDOY8f7GictYFeJj4J88Yh1OuxSynl1NWMp
vdyugnhWOHxZMQiKaHBZIa81ehc4MqUpr0xiV+nPYHbIrKhUckK6KCbZr9hNh0RX
hlfRqrVvHZevUfbADc3toWAURP5rvux/9DxjXKxweO+vfSGlPy/24msu2Uo7x48f
3G9bLAfZ/Lgo+HPoEJ2p2x5TJfUxjC/qRy2VAP7y8ky10d2mD/b7XNn0JyldNqf7
KDcxh2Wedq2iyhz89rbj4WPopUf+F9Oz6Je+EjSbM3Kw/PvdEL2HyW2B6CCY6mOf
s7/wsRlDQz9GICSpYweX1W/o1Fv+E6s+Vn68gACCe5Sn+RMiQupAVcxx2fF3s3OW
Tn821wlOYs54L9ITaoY5hT8RWKWW1Zacx/yUPx24SlC6vaxWWltqM1fmE9W+HdDw
tVzw2WsK7FnRX4L5ZT3Av6dibYbv1lxoy0lPdwDMTzri+DG9v2mLpaWgig3o/koy
3EshW9U0FZMzTfV2CmojOBcpxrCjpwHgdigt4P643p1AgvsugzmRcBQJx2e9HFp0
NueW9FC0KyR/tqvxBIKZ54xu3kmUoCfVJoB2AXTqATMN1GU7/orWXkbdZmCkNGNX
44yoxwzpvgFOZSTBgQpCG+6XtBiM+HHmLv7zIuYtL3CbD201QQ7BtNnqMYIiTGps
v4iZ9v6vzUSecB1XEEOOrtMPrXyhLSUOQnZlH+MK9Ev/43cDOD9eHimPDmmG5fUP
NbQlTXjD/GtsJvR4CbEgdVG6qB/e00TuQjkoUPa8K7CH5gJ+oWH80Nx2WYiTWGkR
Pn4XeTRbf2Os+iMng6wRGHuJ+8v6Q6lfGoIL6zHFqfa3mXHk8mRHHn/Z1X2xDTZ3
eQTywB5yYLtwjeqCt2bhvNmW7vaRVk2UoxSvOPRu0wYGrwZXpTc7GiY/V3CNDaCu
VO73ubmT2dwBgxUfmai0LPWfsLAmmwHm8DQu8kTF6SHWxtIb5zqt7zReu771wqMZ
jn8UtHOHBFzzPbXUQkmn53RbH/NQgimpE2XbR0gdROWg9mMqYxAlex5vBL3fJCGy
kRjpWjuTodJyugAE5PmlU7rfr8BJ41MAlDqDTay+vqWbepST2NWwlLicl1GhJZqt
LMIr0ybaQXpKQF7H3nFSf0UkMnSsBXw3Ur7PFGqIWokrGjzO8XgLcXwhjLx+Zw9+
idCILrABbJaxo5Hr0AFfO6ob39wzFbWT6obqbycZrpdVXQwZFQKGZXtijfNPc04i
MljSCpzC5bWJut8yBHouvj0Hf6IADyV3BHAgq4FABsFrIgK5jM9i2ivKrTYjJXWI
cMz1CV4qmfxerY38BKHBIlrTqSsY09raVIwuctr2pVdOuA0hZ+RnQTnRoR78SVTV
a3i0sB8VK6I6ZSpNXyNee0+noAvRCFPloUXzguqgNYX/85vPgkTURkaLF9IrYdAp
C7Xi+/GP32GAXn/aYMsgDk2VptDCxlg5MAH9f0hM20ZIVBeB5zDapCNMUy9HI14p
zNGQBYIKKRtSCg3PTtG3m7iZmhy16eXVWNPSAkE1b+nRUtDS13PwPwfXy30lRHyW
n49hAHENGHaEJXcvh7qelwSdBR8lUQa270Jzt8ZGecLBTqoxSK1XAJln1ATxPnxN
Y+Neo7tu9zqM+avKJlec1wC+dg9yEn0k2ruZarYx0iW6AUhXypnWBqlbTM7MyEX2
L9vviGUBfxZ3nvzJ9MLYVTHWmTQ7RMveD4/TS7uUYTiW8M7bq/S4vyrt8FK7EpjA
t9B49u9jxygv4kPQHjQa+L5WNo0KbMGF35pvwwljJsExVJI/vVhSdYDJ8BiOn0Gs
eTzfTEmM8EqOTQj1q9hWpZtgGQEsOMo3b6q969ev7yCM5NwsckD2Z8Wj/xObhRCo
O32jyiWrXttYIgWHseYhQql3jb9MwLviB8FHcbMv9nMVgSz2ou9s36fMYez44yYh
mOtWy5G1iDoYKb0LWI+P7Ayx3XMgKnjlDLf2Y8qDLr6e9s7yYQUcy9t4gcjRO0jr
85NTpdheyNgZfK7PIxhXtPjcPmhnXYtYmSzZbCfF8s8jo1POCwfcIoODXSN5etb6
YKxoKMSvTRf2e1wGEi62YjCLbEBo+hD+Nb/Ya9HiDWVKYrWn39zSRkYseCRQM+He
9Vx3xOMddCiyFPEh3GuTaPWSeNntVuEBzgCOWBKPrb53qxFTxjp1s479bpnq8VvO
oQB1rhseuNV0PXtB+ngGhRXpIjc46RfdAKDe8QQP+qhJ0QuMpOXm9lQDA9D8GavL
H0UN3/1kHjg/wWHfsGJ8payhkd3Gz/p5It/lseJB4nwPrdvAX1KjzmHUI4rgQsYL
/BqoQ665qLMTF4VsmZuauPwAhM2rUXPI9RtM0aLw0iJ2itsxbNl8lnW4XGUIBO4M
423spSwfcI568ajTcSo3drhCp02L+IOx+FHZXv7f8K4fchvcOXuGw3hqoXgKEnyF
5Ixb10/yC9TvEyVQCCBDJBSY8e2UeUPQwHiPXuu/oOvFbvYtCIVjGOI0wF2RQXFM
c61vv2uxeEhGaM1lRvpz9XmfhnMgXGhjEEEYfg+7B058Ksqgs4tPMvi4Rd4gW5tt
GXLSLwnEvqAlN0EroHFw/dVlYtpU+pcEakFZbqL2D1e+pTeeCZdr4n00Y8e/IzKP
h+wbmsO9Nx2/AVph8OUo6aBn4iZjgyZxdutrccEMN7nKzzWuHnNJJDP35+ePT5nP
OMKEG48niDP+5udR777G3HiDPFQVffb5HWONTXbk1ZgDQUp+VtLq3vcnknTOVfL8
m8wxETj6WZYsaP0CkvAsO/tRTaz/EgjRraYAu+U5/dcFFgeJmeXnbaxmwF1uJ1Q0
n+1ZHGBiMqFIny2sqm5y8vR2TFSS5czQmVPBdBXQQRPVv50P2XYNPNELXmkEkGp1
sDwyvRm++LQdDlw/YLNj0LhrQGQKHXjyLdzzaTkMzp5zxFKnGA+tdEXNPVbC9zqO
Y8GR4dA5HOirVvLjMRRHwYzWoKhdTO2XNLVYWi6zQPra1ARaQcGwQ5HMBR+kXR5L
G3rPB3P3yORzlJHSfYcxM3TYB6H/hXqqWhMidhf8IRjOb8/uJ8jM5/CcTfVPI9Wg
J9+RfUs+8zORppfSoKYoreOevyQ3+1apmYEODLAQnQQ+8s5KVTJcB5EeOADG3kIM
KvGDzrBUhyZe2CBmUZEjYQ0zm3LBG+JhvxU1ek26gnLpPxIMzYSVdy+5ToEHryt6
YSYnFPmAYd/ns0UVYIOCV8tVIjKixJtgcbfdea8/l/HBAH9mGN0/chkrYVnrlRdT
aUyZ/4LLuTPF9V8q/79Yxpbwe5wOgENcdTAwmdhpDu+iRhLee1cu2BSIf05yrORT
pdefNmjbdqMeXCZpgpQXAIEoaE0Coe82B3+0SsG499myDTpZszRKq+jEdBNUTQ45
q4M5wdmFTe6Ze5GBt2hPnezhP8H4S5CQqSvn6LLKF/Q+vdpwvJF/v0jgDrMMgIMI
o7Lycxr3sl0DpJI6IW0wPQORCcR2wKMLehQ19MyTxvfQhTm+i4nTLymOnwxrA5Xt
i6DJ7DvUgw57IZzmhpsXSgvmeN1qHDYFK9hVLF6iV6fpuYwCWmSD64A0eJYJFGmS
7f3KAGvUAF37wj6fQ2AM7BjyRO7tUzMpCNDQvtd0mBPz+/9Dw7e9CQc+l+8ZdKv/
jSvAHamh5vgXb24BjtfBh3lQBHQOuCJDeZvhgjI59mrsWiLwz1uER75MiuuVvfyD
cHoxxNCyGYkLFSTRYE81xRuBpSvYjIsI0kNCRyc3a2t2Bsb4f15rJc3YWE4Feomk
YiK5YBCzVgt7rDzeyYClCsQ1O5fhHd5qlqoMjlegNjBim5PkJe7uREb8n5TBltnf
fV6DtPinmLBD6BBFNGHMqYpuc8zPbqpI9kLjGeh27Lkn+wkWVpGtX3Kfw8WWxxWZ
IZ9WTshqSWCZm0dhf0vGR6pClcXFV/Gjnqod0uI7z7iPbc09Pwng8JEx4YjFYc87
ibjYbfN9CcuyI5Nxg85m7a1NCYdnVnht4WDBspu4Xwyinke9M3UsbCXGycFZ5/Cu
0gk1Q5aH5IGtHZyBOjT5J79YereEBB4HAIAXBzyFE+IiZ07AmMzm/0jE2oo04tsA
A37OlqWg5CxlHu9zN8nZi3azaAisZfCklUosohh4RtrtYL9R6iANtpmm8vtMr3sv
8xQ/21qBUy82/UG4EzQC846Mt+SZ1RoW8lhxuyWEhbLPgtiuj0tsR/Ck0pY/Gv7i
VSLDZ3f/csNhRkIJd83U8bY/G2L+eGmssxDF32S7JQRd4Ky1IAd6M52ivn5ASTEL
BJhf+V3fb35b0KrjsGemTeGrP8gY2hXvn3p+NgWQOXAcXVZQO6XoI9vgC5FkMaTf
rBZzIGNDiHgO2o9yd/o76iS0ligKl8uKK3Je3kKUk3K1P9R8nAJFT+R4a3v0smBN
YSf19eK+0VwWVCtkoP+j6D8H2GjpEB+BkrZAJCsHfKR4p99Paon6TyWvRqfi33to
t0vVtiJri5tUKP1rPD56fIiPGv0QBdw4QOGNknAVK4waj/rlPS5xQRnG+bMaUKaM
u3nLHUgaqUiRyFejGWYiZc/qNcvv0ZZ1qxGVgRi/WnEw4RKcXYnOum+8+9zOivvn
V0cf0JSRU8zTKffmow7uG1tzhQt5DKs0kAJjQQCybQMvfjcM6sfNc8VFYTngpw1i
9FgdN3PLa3VFHvCv3kM/liBLpT6QDwYY2wsgE+L/kII1PSXzcfQtf5N20BHHaknO
s2bYEUTBDi007VnDJTLz+bT25iJhqd9QSnG+bQxySVon8cU34FLvUlpU+1tH5MoE
PQUOlf0Xsow+nNaqc86xuBjRiPtW6CRYUa+07K854JQtD0sRW16BmrRG42pabbRJ
cz5g550R9Il45DHUQo8pc4bhTJbT8jr7zWvmLo+7H/K6+ypggguvitMmIcc2mQf2
zHc3NnNH+dwlwV4K30/MuEWskV5I5rxqM0dfamqST+9cuOyBd8bR+GdiAVn6tbVN
XBxFKcRRjGLYiJFAKmmFlJGAfG8MkJXvZE8Lyovi5PhVKWILVtCVEWFipeQBWiKu
QbYa4PnqOaiQYsdPU+6F3fuHUqYV+17qs0mmyt8HqtFLlHlnIPUDwUAdXz+upEb7
AVsJd9tsvjIs7Iup7IZZNjBXz+EUZUNztoCEBQPXSINSSzBJqHg0OcAcVXwmnFm+
x7dX9chn3E5L4z0Za3OvlP6/GrTjcdRMr8p/A63M5krZrRx4+PnLeoaKLv0wylyU
Jl5HzQiAl4eiyQ5/myXlWCc47XFiGpjngjKzPAXFaNI7l7fZ6wm/iyZXBiEPStBD
SbaXjQbuTFZhdP3eT06NH7wF5448ffXp2Ack9R0hCNuq6MKsuUSsdNQY7B/haEnb
Tk1QVjtarNmYTxWHA9wpjgeCiDUdFWyTPbfHIAWoab2fGkKOnlhvN4ufXgAV/PZZ
IvO6tf231oxlU+NU3rriwXAhDOK2eJX19SOLhWBctVBgEA8m1vCjOIy7VQFOSkBn
/tmTqucrZPkK2SuCZny94EM3Igf1Sf2FwOrZqNf2s/LaiExOqlqe6S6svOuxm2Nu
CcJL8cjGqHpyzmSb7qKyF6Snn2ijPATrLKlrxV4wByWH64rUhTz3xfIC7buFyH5T
IZ5QtkFLs6uUQtlzzvkEK/19gc8pjPPAHDKFQxt2KssuRZtKc0cegGNl5HW1I7v6
c09viM//L7jVIi5Li7gj0nY4kv4p8FDCjgAskjzfl0M8uB/EN1FynUzKQU47EakC
57rhNZT4s1qMSFcZxrM556JmCPsGPkRL96OOy2IZUUQBj/jQK8St2sJYUHjQLS+K
KzfcXgbNdbNk4yH5OEpnnIkACWjNEpig47UFKrHuEoNQ6A3gL4n6u+mXPMAfq1v9
ZOhzAj4XhL6oMyTcAPxhb4g6BOEbnIBgZsHFvJ1ue7cJiLiPyj/8tANVMY0b6utX
uwKJThXGXeXRG4ix/RRckPhrlvJavCzkfTut6OoxwYBMzfRb+cu164rV2X5XlBl1
/SkBE7QWTylcT+ioMoxPLrjwehy4STx5U7M+UeixtrRRbC/WojWsF/eRqG2XVrRC
xj3QPDXQBLIGGeV4oGzGWDGfhtcyhAxu6KlIrskXKqw3KhuO+QM0cPxwzOWCG4En
dtSCunp2Fu3drO7ZXtuERSizEqLhDP1rfhxKB/GVgPSIa0gm7wCdYmrOZBMn31mt
brcIUqpW0nNMnGVEu63Ql5di3bxu+bfPLZ/OWdBDkx4XMlS1YY2Px3qmvOw0xQul
50GjDmZ//5A4baLOXVD2fFAmHLbRvjCZW59/M88mr0baR+JmaJCKZUjXbvPM/gCe
54S5/1a8flsLKu3mEw3qEu6FrwcNF2Xbl13txX68+BYsejkZD4rkwr0yxUIsrKfQ
Pb96+ZLSDsUNjORCAHuWF2K3OWsBvnp0nuTntJJcCxG33rZLn1JpK0TBzXeIiBfX
J0fTQu3h+go64c0B7hpiew688GXhHDMFxKmyGGnEcwgv838asFTbf5YA1ogYVmh1
95mtu73SJ0pkh4USuMZcZMA32ECuUbIe1vZbqEUTmE6dGj92s392crZPKrkLGJzP
P1B/SQx/MU1bLRkAb8gnl6PHFMb2vdPmLV3WRMVZ2hLdfT5VGyx+BYdLhNhrFKBc
X9g+bDNhCnOzglKNcjc2Rs9ow9Xqtco3NLT5PqTUlHcFQDoUmr2yggrC7MvmLF9j
ilUta1LphqXiJ1I8Vg2I3fHev/M+7ZuDdAJ7OEUFLgq3b9t8T5fJNfrZMLHJi4YF
K2POQoaCjEj9Dg2hjRQNAlboVMbGexiLXCP8wnEic/0Z39e5nm1kWsL27zYocRVQ
l6s6F1FbfZyzf54gJ/G/LID7kSpsdemX/kNEDaaXB00o1DGt+TtmKvU26RPPkyV2
V/CewsLsN/BVCf/cEBgp1zc3SoKJrI+JyzSoo7RkO836RVJspl9wreMX+in92wdP
keHMPxfiXGx+Rl99l+rhPkZFcHLdan4tRR834+rYbaQJgZUlbF8ymrntiWKEENc3
pL9ScxN5JTsnoZMAr7tHBXkg3gxyAQXctb5PDxWRdcuWLgSuNccU19O+Ok4wU3iz
951dCSBCzbYyGdmBwS/aFoZZS9qD+cL0xhYTwGsKE32a8KRT1EW0eu00Z+UZYMbA
Tf52Zpt8MnbvdyOq2fmzEWMcSpzfmoWd2PwYFH+MfCaXmYBu/JMJbV3QajAUL9eE
8qGEeeo9TqSxsafj0E/Akp6u95TCnSnE1WnAt0mwkp+Zqmn8TPiRUrUlR4eeHnZp
PHSCJ+8wK+Z/q5lfkFD+hwkxIVEKYiOaIoGnZRQ5wMmnvPafbSfLEvRreb7i2VsL
eATyUwuTQTX/5jQ/aHUnRokSLg5hv3gWex8pab2iZJsf5RrDCsxgC/Oi8ER7sLq1
k5Pz7B9m7F4Emr6UMgpfQpxPT8JJv+Tcsd7vcYBnsfiwYY+w1DMFJETMLEz39vri
ML2duUD5gTwovl/3xkT8e5yb6KanqUoqgNU2B/L/iT069BUGZ5HP1tT/xrRkHWUN
2NljRMVMxSIwj5mDIPTdfosSi3GGJnvfsFo1BKL4XpOoe2vUlZ/opNSMrtORQQjI
9zTqZlVqaLeKGXF2/pfLiUpu/Jv7JLXqxNO1448YFZTMDQbRYh1p/k881dxndWyK
l/KKYSOgGrYKtcK7wa0wL75XJRv7qd7XQJ/aDuCwQEDSkuuPhTnWFW7oINF1l9o4
Mzu9V4COtjewxwy54hX2tD9WOsO+3+wE5jQjPREuyozKEF300jCjmeDeaJfff7Yl
Yx75VWdOzW0svSxMyt63oHF4fLeP+plSn6uUGFEmFNlrsqWeEbrFm6Wkh4hhzfKU
0odjcvjSOkOU5Y8rJyAO60nCHTCcsXJv7lwDeGQRJ6Zygr1Jh7hS0LIsEec1dHl3
KqB6nBsyfr8aX60LugzSwwpqL15z9Fq4OE2/pUeSJ5KWsMmQdnjnJMtNzc2s/FrR
WsWu0Zt9w744gDXxp6K5bJfOYZHdrToupsVL8RLeB/T2lj9my+WeOHATyun0BIsd
ZFbzJVtjyQpHNAFZ9zpkJo2XxFBKplIrAFns+uOHfdSJh2P1AniKNSm15vRf6cre
kYJlsMqMEAfm20ZXeVvD0SlaOBVbPvVjWe0Se5dBmM+qDBt81fXX+wY22rKzx7h2
LmdaexwPGoAId9kjP6K9/iIRqhi0TaTF2/zwu5iEYV5qEtKyNhi3Z2Z1uApxQi3n
Oze003qwD15mx3kCqfz/S8V7n0zQ2uIP7O2Sbzx3OicR99D9nVo3zuzqML5e3ncR
hXNK+lHKTgtwQf7PEVHy5kxphw7XEj1HrQUIics+AnYe4221o9sasNVe/acITMpr
M6YuheZct7zEs6KrOn4IoEyuSlJ+KlhOUN/7HpEpF8taFSqhKMviOHtl1pgkVEO3
cxHSyqYZQqRM9shUjhO9JyG6W6mpMOqgPjKy4Yprdh27SmsnU2pfWw6tNPnD2jDb
/08ykySZE56YbeNJhYQmLDVRI8aG+TNcUlmXhWe1UwRfsd9lvtRrqC7fAH38r6vQ
HDm2atPCruihr6pLm2n6c8Kf7R/SHfmRaWfHHOFaoGoBKzLQaJMN8qk3x9O21s+m
7tj0DKlRiQFODUMZpxRN6v73EuIJhdNLCYOLPcka5sc+Ob9382o+9P+B6eS6zNl4
HIOzIW/mB2MpDw8cDn9TxlvrgMaZ8e6LIoP2k68wYLR4QJbHe3rjMT8P2rvfh2Eb
+ALFKoqXUhssBMnsdaZkuVDeCqbMB6KE6r2NBxw69hfziVj712u+EwF60yT4dyO7
kebmTXhvSU6dESsoLTi6D/Nw2IGvMys0OTCztWUb3H/qI/mnXndk8Kz+NLV58Rh0
eOuoyWZ9OupuSkhuABb0Kk2ESVJdSXRj3wgLaZgk9FK+93sY981gwOnmxAUfL1Iu
dTc6Tts6STu/bebeIfKMcuYmE/TEhUsalhrZrmJtq6chtTLtj7XVNM8PvawWotbi
xEvvdqfk+9VbA/x6+KItWMyuF8TOWcxGLS8ZwFYQRLHCG+ZWrcwoK6mxDV8AYox/
w60LuMeBCPnurSfhsC0N/V8qbHLzYKnU3TvqJbNMv+IveGXRw849KKMeUAu44/5r
m0Z3KWT9wqF6oLvPtQMG1us3U+QhSps62vXTa6Dk/ngBK5rnkcF/vkHDsnsdNv/v
7/ZXB12gAH3V0N43hMI4HbNlJSVMA9mTaIju+bbRDyPyfPuauVxC/9RxW9VO0jvC
sz71Imqp9uyLkqYYY5HgCXN42Lcib82a/ps6RaE7fcu0ScNZ4+R1/h4GbwackHh0
WXZ885bBTCyJAGqqrSSCZkglnRBRIWzD/oQ2zVfrDavb0k6RtWRr/cUPAJvMSSsk
CjbQcM9P9YDkaCyoJ7ERwyXSPgqFYjFaJFwYLmqLvt2bkA2MKAynA7pHR1u9605H
qk5Gx5yvpVwoN5dbu9ct4msMVdZ9jh6mZBUlESbpIA+H1piAixD+MYf0jvcNbCk/
1MYVp8jOYPhfQqPplxqpFEHMqn8qxakjjpKYffsSYBEy4/M3cQl+f300kYvNgMGN
brjfouKm45Q+jijJ0jOAzpSXbK7yH62+/nUXLLT/Np3NQot5jL7YgClJMxa5Xlk4
ayaIaBhjfhGHUUCswb+fIdBqhKWiJDuJDgUtJMKCTwmcbsduYRj4cmj/V43hBW7h
/GJwfyvOIrzBgrtsOV5n8SJGqFu0D1Nveh8CIb1IWRk1KKa6soGLnJDGO79L8qKw
oChtRGApHzLF3m7LT1lXQqnK9IX0gPvzBrjeYIOdzLF+S9xvZ7d2EYawCbWbbmNh
udiYZdYfrv6iN0/6IdKepZCVrhlswWWHCZY8z84uKX7QPZ+/dyKUZp01ZB9uJ3A3
80Ep2oCpBR6Px6adyxcPJaHSCJ4JlcXI4B/ICeEkJBKwbj9BnoLqNx23Tly45Qfk
pbTXRiAkzTjc7xYTTj+iIZecfEQn+x0zQOya7AkB8u6EnX6ldkkdqLLC+63PInnt
ingIL/7ZoXTQnf9G+Y1jv2c0Ui9HPbJNiFnSWgP7AqNES51qn7ZXaYt+04WpuYvP
oR9mAGNB5s6qLh3o1iAiLbY6awdPOodqoSpeCFcEnrXK3nq2O6eKD8125ydPKxEB
seiOQlzr70z3B8Migd3ilWwO+tT52IxtzgGwfVJ+InWK7Rs6PPut7Dra3xTKUOUz
I7kLS+6N4MocH8vc3eXprAZVKx9jOm7wdinl38jy0k82wQzh5hLyPCFAen5MzMlt
V3eni5il/pjchKxXcz2ifhMq5qk59SiRj22eWQ4BBN6YgvqD6sZtyxwzN9zBbpWr
uogNHUdPqoj/SJsaPhAZfweZkFvlVrfSL49iUqoYm52jAEkEt0o8g1AnPlfd0ddD
3ZmR7RfJSEzRo4h9umYZwN/j4+Ewh+tpR+ddXBGOuOP3S9L+xiu7k5xHAyGDhHn9
nrJ5zU1XqE40cqctWedzTBRUHMTr2AuusVNModZstfVjCN5HcJlt6lvE+aCf+i3C
uPOlDlthFF1m0NqDgc+fGTpNOstOAauIEaB9a90v3zgsjwqAcJ370v2mEB9nNB4q
nzzEq5qiOJZnnZnHFqU0hLWdZt1wYbViSjrTLNDl3ts+EMw+fSjOrqMMyrBXce5x
HDCBTKn3uZiumsZBZVyD/VoAjXshjsKvqMsX64et3W14WKPKbRJSMMBuZWGYECsM
TS8pU5yvgZxkxzJ819SdZNIYqg69So8yqQgx7ohpKiZQDGul+yZ4HG5wBjiq/Vix
efm05Bj0vPRBLKiFUexQUSHwZm+CtrNjk7Wwa107hsEB+CWrkXmKzm9vVMsEa0vy
hCjV+qpvWy5Ijs0XtZ0qfVDJbsVYccUtBZV9o+vUApSflDF1s2wjOQKK+1QMt1cN
2XQnyadjoA7rMnzADOzoBhIV6u7gQVBLqmHaIAettlNMb2tqmZlA3EumFycqI5v5
SkS/lxJhoXrLdjEC9+Cq1ZIEbMWuKIQljOp8CZbw/GV2p5FpFTo21R+VdfqA3yWz
iqNIUvqN1NNfdD36kFK5xT22rdeJ0viFqAU0kD3o2adVJ4XPJTAawj9rKQwDCMhj
4L5k8tcdgQBNgnJ2niFbkRv1lMXSUv25sA1kcPmAatdPYvyRDz0+m1fbFITU7MqC
XTvrUDsNrfDbRyqC3ISEBWB7kMCRYDwmof2mz+TDS0cbh1FimmPHWaQXbXibXEW4
eGSMKCkb8xbTsY3bCmGL88A1HZl8vde/gFb9yeR9XKtUriLxIle8nm8WbC85rfbd
fTXXMaTCG8+G4ILozBbluyd1WwVVx8yuxGZedSDhFDy9fANksHCQiNptTaX5shGe
JTCZawn6Gj4DuCzuTihonijdOg7tyvvOnwo9RqjQ6cb5GFGw6zjUhCvMo44GtVgm
zAOo0FyTPYDSR4nYe5ph2G69tfEKtpennVzEaZAJ/ZQFikO/vnfx4kselMmoSSp6
iERU2q2NpFXxQQ0zfGExqKpaUcUHZYKd7H0j4ZXWkDB/OmhlnDUWVIEbNWCk33Gr
tFU4gXDWGQneGQsfm7w9ensT7BmlMu1xeHVvduGvVMXvFnjZ0UpbAoooarIDhvyZ
dmlihMoFn4UqjplYnToJ7qlVD6nwL30e5swimpuXQdIYnc1mpUpT/WSAj4FNSaMD
1Cpg7BA8KdoPBQj/UfE0/0tJVNDYlOvsrqpVZul8I6/2DdcmOeQso0ZKqS0/Fb8+
YfiqA2v/IgPhwlfuEkUNMoIDWJceA5E8i2nwSVioX3B1U27IFVvRNMzpFZ2IpSc1
fYgOh7qc/zJ2q82eOb+1RHT/ceyNQwv7ODuzrYV3Y6RoYL8R0KOgPPc6FB95eFyN
falxjreu39RF3kJ9wvlnxc5dO3wmeJR0fai+8kPPRDywl5DRySJM0Q/ub8sYeh84
7FA3SSrmOcyLOlqcPQmJjBroLf+HFXLM41tB7lNyEFamhNwVfexdpCM1mezX/E/E
VbDWPKwf1mO6KnQoXmkQzcIejppfHgpM8QX72q1VYhTYQmwb2JBPbfpK1tm5MC8M
E5T4NTHakQNI/ihtqJMsfHNQOMtcZG9B+keT/o1biFw0yRqImajqN0hRDnnAM5Y/
vp9gd6u6LDYI+NXinTX8aRR1kgZlJNdnR8azDo57w1KJLwkHL9nxO70Ll96N3V6T
Kjz/uQrtWYSXvKNSl28L3Bmn53IELCb6mp+6rhrWpWf9AsQKxTIPKx8Gri7ECP+P
mYbFHgGD2hS5WRppWCCD/bgWyPKnr5ORlX0Bjjf5keboDqPNkrSVx7EpN5jsdvAK
STyp7K9kpHpVUq+DJRKMrm/AnqeJa8rRNKFA7kmZPul7Y5EktqCSvoJcFVeSwah+
nl9fFF61a7eaZ+qBrkGMoT45qT3RRL6InaF0lKrryU4b61HzNfIWWjehF07QyWUB
2Ks1DJZ+b22hm2OCYc0sOCv9lcAJCdmSPMCSO9d4pbwlfm6tPmY1BJOrMTx0Amyu
+uMcJ2AwblRzOi7JiREt5Use8WXYuhVq5fm1rnl17oACkrR6dYO/ORse2MJbqNyy
kl6Nz/kVy3kgViEfskM/GWe5QGugGeLEew68APOPkNl0wkQ/5/Ir4mBo/pw2NPP6
onZR7hir/8q/PSh6Jez3Cb+EGFWLEq/HouIjbfiqa/NRrUs0KvKV0n8LU7i63J7n
/QnkgVD4Dr+GF6ZHArmy4dbWqF4XAGQXeMGRN2HdSqd2P2A7oaaBth43BUmNL83i
ImjvS4VApbJr2NqgNeOsD+91cFQvr9TlibJmR2ofw2DbS1ss8KlU1B0UDwxyTRd1
W+pMvMtBu4BQcFLZkJgEEbL7E3pgJdgjCiSlF39L/xmCqE7nUfwQMti336r4+cso
fDf8V4b5F32qdsKQJCrfDyGZpOnfHixzSqDjfFGkXTwXtionQQA1S7d7M4UQ0O7v
kwaVMfkeTf+w89rdBDtsq5LRVfaYTmQjBTu784ib6nbYkNb0p7BEPMDtzvUQmePU
iwk4uGkFi9bRqVztgRQDeYT1Qb4A+6IkDapxCdRQxX9sGvD+ZYdOdDc/qNkGNkRi
BLMF0xUz/RpcEsmFH0/rjXdZHV2SwMGJRZxqKtcwSVbUfcRRmJeAo66Mxc/XncZ6
61puPIvDz1EL5SCv/za9R7sUWB8379T4vcIhXGcaj+oLSPADPDwYCK3BQdS7JYQE
ml/0hS2AOy6ojR9Gsc4U1ukgkBf+GSMBSSRcoJBHXDgkl1yvXcFdj33qrAKMqCgJ
mLvfhXzkhLivcgdMWXBOoGjoNo7W1s5Fv4dUWkGRH+jQQwLCSiTOGgP9Qj6pXBsa
4sXG1GxgYfxTkCjK9wJPPyQmO8z8ivQJArHU3Nxa57pSmhTnMVvON/FAJ+KG2DPd
3trxioJq9J2ri/z2UzXbjY1vD1tFQCg/xwKENxkSEePMX5+jC7l4FqyJbJOgTb4R
GMRqtxOhpJa367yBKeFwikMSXMLRuSkCkCQzci5xDe26kOxEIfs/Z8bB+2k3qdZL
exji9dr3fbF4i/TytZHNf1lcNKO2///XnC+A+zZ8wOkNFoSExPJFBxhFFMUwGRLQ
hmkbVmWj/y6qUTw5Kk16W4O6tTi2NTxqqNFu3OnZ+9q3MJAVS6yKgUeO44ZT3fSG
5+tUO8DuwxF9ZM49oB+1aUzAbmGOGNrdWAXeT6XZzAe/309BEtfUmncYcSoqMkGb
hZ/9D2P8QyvPQmBk+8TW7wtylyb8qyy52i3go/gqi0MczfSkDoQ0gsFjiIJf2UGj
M4rRXxxwDltLWNIiQ0QbB80PJ87IMtXZQLh689tcwl+JXWBtI8PsNdYM58Mjl1BU
Io4+ZpZNNIB3RbkBbDhvCpaC1re9rs3yq6scMcQ8R3lfUmskvlbJS5LSPDzYxd+J
9zx6G4O5mpX8xx/tl+LMQ6F1i18EdjVbQ3DeXf8fv4RRq80TLsZxfUxwsPPxu/qK
gjRIkuiZHEsBJzb+M/KiRf5tWKG7o1v293EoewkYKcbJlLXJDhvoBJy6VoTMfFfF
hKy4d9nJSzGlZYt5Ya7qlevY5MLRPr5tst8nixAQKGTbneI5hL0DuJx+zVf+lgYn
8wAZR4zn61vg9uXwJgmWtYgLLWfpKvr8IG7DKFR9Qq2uItdZ4Pb+UZMtGau7Aix0
nN9AkDuUw4rhDG3Xqd+5om2mUnvhHgbKD8UbYOerxUCb9kPUj0T9HRVlYVPpE7jy
LUsM8HK60XQSeatfOte3/yMoHRGNOraI0UhPaKrJGsBWuqvZ9XWPKkNQDMJ21PVB
I1hwJfYjrYGwRiU1fy4JXB/ovHH8EJM8uCq5aFQsJywGbQI1ihKoxf7pSgt6IPxe
6Wvns9/fQVD4h0PbGV0tsiV+Vk0Ye8ZCIwpI0KXpj7AQxzmSmVsduV+jtdLHiSc9
n9SOVYOA34mQbBK5ikeVh6+v/u6THqb5pXjsHv+GTvaLEnVa41XUISaG2hrDUovX
3/angO/a2LJUy/96TmfniaggtnRbrbG1VcZ+G/hrCYn8NV3AJvB32GV1HxwBz12E
Vb8oCfanCrdHtE7UazuVHzA7KU1GBGJEjU/lcBLHPs07mmie5Ko1rIRTLpkikDtu
HuMdqmnUBVpKwpMlks9yTAUlUeDTyX486G6AfWGgwQHwWXOhZVFAjiHJYk1yu85q
LWpfCauFxSDrKVobsN/u+NoC/gzbw3F/ji4X4lSj9QzyRkmbuuaHYM/D3fW7DcLb
1oKQmNRFetDQDBI1E1Skh/ERpXJf7fliF4symg+3B4GFwq4KJr/A46R7nWYtN3O5
YZq14lC7bgRySxS+5EXmjA9qYaSTQOC0J6MucatKO1E9KsitbViHKdndrOD5yZjx
VwUp/+Nd5JrVm7sxCmBBtWp1bkKPy3NwzMmLl73UtQ2FWPUTXlyJ33xJQ11kr1T0
bYISm5VRD4UN8slelLpAETq+uKM8NF9lzP49myE7Nvrn9hHXTE+BrxuKnf0zkWon
31FhmH1MrXIwZr3dPGsNyvbdKrWtGeqg48nrGkqPleIKZt7DfW3pS6fPZ81/aytl
8ae81OT9A0Q4ErvHahqke8jsNFNBDAV+ntwUrbPqLXI7Z51tFC3mFAZZNKxFuZpP
tB/zBxk/ez5Q6xT+OKzaKEDpY1meUpxCgbS+/wyum9Ndkykcdyyohvaf0/GMjqcU
ubmyR8w2eh22txtIEsNYGPIUEgujZxy6XpSBruG6XrP5G6f5Avg6+RLNDms6srh+
mSAbMdAFNO57pxb+ZoWwivvxQnZE6nD+WFpSDr2XSbivyK/3/iNLuulubmdTtLZj
5reJIz+qIHpESeOMlsCLjevyVnBOpzr50hHdAtyQRkWrHzcd38tCCY6vwHzmkq8I
9vGRBTfNGivukgRXGOVPPTArRaWNfVCy/FhNVHy0VsG5rJbLgCBmW5AEc5oYSYQS
pGVAUlCVFSLfZyFusyuo0/ICQYOTKoBfxd423JaugYZRuF44nKTvWPf1jIADbxTj
CPahvYC0YVcx/zoPwX7fF0teV3RJGM4M/MXrHF6LyGiTifSUxyDiRw31Wd0CtNxr
/uiw1zFafSpv4O83TxYugYUTiXPefvwxJfW7X29c2NhwvpkcAde1OdTacszfXPRc
85k22KLHxoFOPOUTBNWa9M9XU2rYCzaiulYiYQhuXLQDoZfPVh7LbRr6TooTICpi
NSKweztAAv70AkryJ4rVer6a5ZBoTgu0s8C2G/vsjnmhF5+5sk42uQvbUmfzl0IP
ap9JnUAi3boWybg7EF4rOuBeXjhQjMU2o668ovxdkzEEroMSfKUFfuuG7rKws5SP
zI/wG0dwhkmAfy4DPljzr/yuedbEj93daty9mkAWOGwDEO80o+BUDf1MJUkXg3s0
ADGKE0vfDAXI6gQTPkh/5KWjeWo7KgDHPB3FdVjhLlTmvgZaZCiF7uRfIKBmwDPO
mYAFR/ET/iZQSpGUCVOFb+I5H5hgLdN8DkwAu5qWJRAb2X0IoDU2XT1o8z/77CMZ
8EEr/JtrKqo0bkIH1hwtYeNYMFDKKDnepQd51CxcZVeNBQgcp+xhoTRRGn7QV2jM
Hp4qkfEgaeUQFZUuVyLSq+UifyP6ow/PSt/Thor7mYGwjJvU+AzDNHFsoAyZAuCA
rpo5gB/ibUXPpTjEI60sWKSVH5LDjfXbwt4nfPCv5aJAt91szDqyKT22lfe4Cbtt
LeJoImLxhHu0Dy52R3ghzeqcq7TG+KkPjO3ZJ+Nm+bTgdItcj650WPjQtDTcGZsJ
KVscw9W4of3q776PWGbNe0CIOqHO0iCPg/nFbNYJ2WfPjKPqcU7bVS5xPcj5E8M7
Yo8ISG2KDKBZhqqhocEMx5KLIsAa4ZiY6lYvxDKk+qK9kKCD/QsK8EXxX1rMPBBa
SDc2NszJTUxz4al491TYiRZRhEqoqZl3ngP2PPWwh8I4NPo4+YC8uvtNG4jHXniM
COTka8UImb1at5JYIm9z5Su3S8W0H4Kc/LS1V/SODTMmOtAmeUpwjP8sIzsYd0Id
wRXF5NLOdIu4M5abKZzYR3eaYuuBJ6qF305Dui/8w22SKd6xn5/1OEbnAFURApJE
rKEDB0xPgheXpKgdNZIdjWrTPrD7d5RcS26+hjEHdU6vzMcBIwX3w4saJLYS067J
UYoZrvkPo7K3+0Ds8QJLk+8ODA4AXMqbmeTlPfi18XDtwA85mAwFFwT6flDF4djN
6tDEKsBfyWg81sXKZ58hyc8zIvJm66E1Awr46DMX6SpZL/W7+MRpP/SjztCUC9Dp
P++jumzfEy6q6RydzYZuCL4y0XRcUuZ3zE1jHmcKfS07YYpMGF2t9dRl7BI8RxsU
BREU5psYeXaxZhdLE8Ttp7EmHpsXMQrJmjaPfaHnNJ6nEJEwP95ioNi+QjGMU7J4
gvbSRKaeXby+CcOJ58JpPYlkUK3GlpZiRI9FRkWsmyWIjKL7YI8INO/pLtDTaUES
unE++3t3Yq4j8FRIinPsVJkZxxYT5ki7Z0tpSRuQ8zyVNHD8GW4TaFDahRwgFnwS
4q4H6A6swAN2mV9+i8Fi9WYUdmWRGzxlDE+nZ1WQeTIgerzfTKBwDCygcGfGJ83y
vM85AS1BgyDxMlQiBiKBKGzdLjFZcYuOILKWcDtlRRWOQuJG1F1VzdqV5BTAqXAb
cxCzDacGcIPwICLrDAizGXTUF+E2vl7ttGXoEf9bnst2m2RSkVr73B8VRL5cz9w2
Nz6bBywAh0wslvtGrsDAZkr5WMX794IE1BoSiTaraTO4nn8/NWi1Vm43+sCGmzC2
kHjlyxvlYbcnEk+Osc/SU2o7Bq+qpTNBrF2hqVuyqPQzr00039cgkVUgT015JLHv
1zPd0t48sT0lABjTn/Om/oJEnRc1sxagoEN/JlW087DB5aTeceie5WfTzS8vFd0Q
btApXusKCWQ9Ja9LyX9Xoeu1t4RMfWozV2CxGE7LkbjTvKteR+hOXCzFCivuRT06
AJGiQ1ScvVq1RqXL25JGGiGIzdD2GzuYteN92wBPdGDcfpNchK0r9oYAde+QjESi
DwVk9+zzkDrrUdrgXnVRXm3y2GX7ZrBmw7ffcSmNtt9Oe7EA8a46yNS0oTzo/Pc9
nun309J2Uzw7pMWWAeTg6Rl+vjAdz4F1ltDNKPYcXf1i1Qd5u/9JW4bU2C5th/0j
6+COwsJ/C27LMaxy03VI5hJIbbb4ce/KeymnVlsbPqYvQFx71D56HUor2qCkwgme
P3XzsyRhkTyHj+vC6W4hvyLyCTXhmDHz9bGqxNubs6lmjRjJMihpOKPH8pES1x5h
llA/EAFjx4+u81FwQd3wE2KnF6PdM+g2Vb/LY9RqDS8Te568oxSNTOovekvJOoLa
fZwHqhg6S7jaZBTAb+QpTwAxXWctOC3j46Vd/fUx5PvZ37K9FqfxSEUOZbfcfwJp
Go1tUxoPPuhtqS+4kCrk8zygx+5oN/uBIaro3odZq87ymdZ2zzQHJBfnQVGCjMst
Fh4gK7Tap7anrk/BQUOnbCvZ2jxJids2MR8klEVa5wavkP7vgM9pyZV3HRHXWtrD
ZgVFUxDuf2Wv1Bj+JzajB8z92vD2fNPoH+qERHFaSuJHIsYynPz9/cDF/EngRrR1
B7xAdv18tBH06ar66HjfazkMnrLaazP4mTEg7T77I0gIQ+SEAL3xiAvCcW80Dj/f
Ejy60oixthhlYgAlLbuRPyoExw81VNxfrlV+/b/j2u/+q1/UXaNnHZhTNBrGuFob
jP0fvWOgfgpQ65yQwayHMxEybwATTmrQ9vxerSaNyoG43vMA+saFvo5ZFAne8kUD
4yZbpjx/Xha8CsBP4OG5IGbarHxy86WAcwyqsw9Y2DuEj3dURiYHrpCJWgv7gRuz
DRUGYVl8lSvfgH7TXQy8scK2yrOUl5o/h2UxL5HeaxcFmiHo7aYEtepkxBAkwwbM
+GHwPB9SSYxGmSbCuiz4htDJz9yMrZ2tA6HEouthR171QSElnKiHHWH6Doz0uY53
nW5tE8htqjygtd+1UNzxnNhLbRX9U7qum5xZpXVjd3oUcoRcksoRgRW9fzb4+cTe
luy5nfsHr9g+FSyh+i36miGk/7QW4zm1OOABCuQuGWlauB9z97zs/Wadmx94dlon
thpKkDdx8iL64D9sEwUsOYGb0RA9pV5/TRzdFCSWPIWKHW9NxNSIuZ6i/TPNoXD5
7D7ZWEHnugBvLDpbqtv7ekjlTMOvQIYpifL0HOyFd8xqJ6a6K/6MNoJL829Yzb9F
v4j0Dx64ZyHynVQuRV7sMitWrptZQqoL6AwLSc6MXXu/Ce1VVAjDwyXEZMJLv0XH
RU+dETCgfVjfDpsrTciqL+FoRZjlI2x02SnGJUm7Qdu+qTVoZ01tVZVgN+6uRqZQ
fm3xEQMOaoaX2mogXswKCh20UQ57WGyRUNnZZUGNu8Yg72qm+ImFl6mQD/C4aeQT
Q90UC1DYPE0UFxd86USQKy7hdsAtUTt2yK9i4J9F3XoZH128u83X0AaF+Jk60cZq
VcM0BbCkBe/STOfMFpIE/kk4DbkuvioxF2blHCv4tFz9jVqh2VZWlT2bUqDwiheL
i6pKvrU/2Ec1Uexr66WTnjTvB3iuKEwr2F0LdMJssrB8IslX6omeu7VjvgAPaFjN
m9mHiIcPOMATbIF/0a6zbduG7lh3QOmZwM7xKCTnhoGHgfxY2QKBsjcai14dPEzf
F69Ly692NxGVL2n1Q3o1jra/YzLWU7uIxJhSH8uyiv5pIc/GYuTqUEMt3M/wAcGV
sfC2AF7s0XJuqjeVbqvyPo+ZAtWiMcTK1UDBLFU9/++XUtsJxn817txtraW1VADU
kH97ip/FiYbDp2PRDPdF52SnOnuo2oKm+HjPXYIxpT7u9c2e05jGsIxNCPTqbInm
mJXIqUtRlTyn4Gm1Yj25kUU+qGsrQfhF8IqtvnX6T2pYeJ6KJryiYO1vv2wcLogg
s68WeM92QaMqmE93wuvFEnBA6fTugMBew3khA0h/c84EPITL0st+fN2lB5Q7Ndv8
t4eft761liqgbF6NvGdIZT1jO0L/sfEMImB2rfKPHHZkxyNLz7VOWwcopxjO4D21
ZvH4En5/IkY29MBWmq3pWEiyyrc26Luni3eSFtmHcUIdHUaY0mF/3n7rxYRJFToY
ug7/8VsKMgbKfBbmaQIS5/HITojquyzMMM7yLLA4MXLQqBo7GuNDos9MMewS4Tys
Nx5unKZSL5lJqL5Yjw+44R7kGWSw/yknIje/NYRwz1vzoQOAH3FIHP21r1sSpwsA
ZNr+sFe2U6i7l07TEqCQWX1a0T50G6XBmwRcT61wFuRMAGOlIrD7ID1sZ5VA4i8j
r0yy1QMnOmLAIjjOtnIk65rf9KEvwCXyc8v3LNoF0R5ZiL5YXF1KCwLu9+lFd3UM
YOyPAhwna6qH9C2Ov1U2yVdLZ+uKDlzaJ+F7PZDD4wwge+ZEW/TvwZ7QMjDZAVxV
A9Uyv4VX940iZKoOlEuCiBS8pBaxvcQ/+dCw2+USUwXkPUsqr99EqXL2+BnlatC1
LtKJW3YYbASO0IlfbDUD+ZNrgbSR0QDKMaUB7e11Z7X5JQbT1ahT2sflN+B0kOYH
eKKLNWAb3DXKjtqdH3OjrYqtxJoS91ODkbqt2OiRSL7JX/ZzNAoxzpM7vV690GFh
FYvDwdWFJvL+ILYpdcVXuFtFu3JXJUn+NPw/az81hna0ygIbNpT57S8dsdw+jg1O
T3amEW+vmxDdhR/PVjykcH2Zaey4tv2YxWypsmaaX6CrsaqpM/U3pI5iFrm+RQ2R
YjFDRTvVMA3gpeaNRS6oJo9SHEOVEx8zKzTc/uaJriuTkVpmJExgr/u1/KOV53YF
PIrqXFkLBvHRfGsJac3hfKRhYW+NYBCVOl84d1oZXl5yrniAScdGjdNQNLOv2KqL
pbPavFcm0NDCLR4QJ3KHZwRAURQIQQLT6LfPJkXSmefzhs6QzMaP6Nc1TWokpdvi
JCP19oar1kh2ivLXha1jeXz+xz27PcOwFsFdtrj89DU0jj3NXkzj5o46+9aB0B/e
XIopI/fFFhHgFCVKMWuEIOISQ0WidZFrnLxSLTpRINtG9xqreddC156Z2+Nf5dlN
IxQiWC2PQCTqtKFXApKdkKcaUe+uAvtl0beoFHCMCh68nB7T/5numjUIYs5WxRSe
eAe9j+0bd73aIpBVidqLodhya+QkWTNTgCKC9MWVMQpkIkBOyUqrKcpZqvCEzpVH
FNdLwcPT6qQz72UyImCNKUdx/5nB/GsUh5ZejEDghC4Tc1dUuvlPcg2v0hfT6Xaa
UKoFzM70h7Z/Ost3HmVr8etnomgqumTs/eb/lPgwHA6SsH+9X5st9k570VTf+ZMx
a9cUCvoCvx3fp2ODGy3dCjuMKy22V4ahteZAPLiagKVfCI30x1fZgl+8PSOW5IiK
rRVuW9ZVTeCWVXZfSemsMMDj/uoxGHDQI0Cooy2ElqfvKBbqLBaTY4BpZe45OQ37
+rx+tJK+tFbWAZbqlXVT3f/aAP3Yf1yWx2+tGWH4GBFvooe6lgJNJCnl8jf4Fm/d
sBj2WmHwmwWrWIFV8zhAy2M8MSWWaTTuBwBMCALkTytfBC9ytbdmvbGad/4xuEYG
z9LE643hxFtnw6mtxEA/B9j5v1svHKlF4OkHbOT6cZAPbUkt6judRuvOwucMSh81
+LVJEF94qiey+3KmwglpEdqvBLwg1wurQapUKTrb4mLSXs5o58dnZsNfwR9itAwR
2753eGT3RX1UZmbb6Yz04Vlzut84TL4Hx3HIDDD7kOuomTMO7t1+/jwuprOpFBSX
dFtacwckMgKNMRsKTn/YlN/ubmk5Z8Xxb2pH/p1p1+3mDzXPH+sXZ9004DOedUCh
+xrcwmHWfDBuSTzGY+KbzTQT6IlUw+DXhJg44gKmHv51N1Gg0ThooAvOJg3s0of7
i7HQibFoVJkRdC2hVZieery9bCOOVVT9ldHLGccr+HVKDssXVhLaNZvwQ7NX1xOM
7ExBn9W63EpLHIHVXleo1M1Dx+S9nehQwRifHOhc74bJvMo7zwIwQmzsTWkRU4zQ
C+zpuhW75zOgJyqfWWpsRp7HPNCaWCOUKRbd4rgT7KnFOIChOT9xEM6/9cp+EWNN
iUWO9GJbOY/ytjq8+cQFB9nHuFBvgcEj4Y0i54ExOqjOkUmgvJusI2kTDyWxSOR5
ovu2Vf9R2sM/K6A4OJdLHikpdgRIJ7yDxowB5ak/QoIpbj7Tt6v2vgAgjekpbgKh
9PHenJ3GF3Y3qvKeRAgJNaKDkO7fBq4bRBbl9X3l6dw6/MxX4XqqeKr2Y/ugInKK
XNXN80v9w04NBVMzJ5csKUypBbv+vlhs/okieT8Wa+JOYlJ5Z2oyrqVzfQ5p9YHm
C9G+GNQSvmlpS5uCkxb/OSLFcuxZY7i5FcW9u++C/UqVubcpji0hmidF+wrhglSm
mUSoQ2CE88kjYvvjtcO7c7nI7uekDImnlSqvV4H4ZKatPzc7tgOVxVT2PSczqhlC
/IFYlei8u6TymlFuKuC2o/UsymK3XTpv2gBJCLKUP8olHAZcmyvCqfQRT5XSK88B
9oDhzke0BnhYKcT3WShawbQrH2/Xz/xP3s/64j7hC30qZC66s3E3CKd/HU6TgzPu
Yl1WTjgw9jJbbyabgyl80G7JqWmplrsy7NM3coUURgNihcRZLADG0UUyQkjUAk4L
BHzRGjp/MVFeF7hY5wsrpkCExMADbGL17TST7UiFoeF/aNFpD8Y7d3zZG3rd14mt
9s71wKCHuqyThyHajY4gruGeaB4kncsVB4q9701qoOR0asIFhDyGCs9h8EHt57nf
PtAXAiwwgf//x2bNU0yzjQCEOQU9sPG79nLqxBZr5t7GAQvZe8r2sjJput8vDxGk
ZRtj49y2XHz03QPDZqVXOeuOo/S3Xkdbvf2GmQjzrtACL8+hY+uBB3c6ZnTgXvO4
8yNqPbBrF485JMRhseX/T9bt/lML2c7jcED6PpVGCz3vM9tyYqJV2QzBUUuMk8gD
Pdci42SmG+kHauXfO/jPARcWXtG8CZb2weHA1K7lai51VLNXgyHziwA4vjFV4689
36YvzEE2DzUJ51yqWlEbU6E61iPOqP16UDN8yS3BwsuDmq5Kea+aWEeU03xHfGyR
FA+O3HtsrGvK4xJCg2oVn8KNSD2wRvxykmyLYRKp/YS25Wc5w/1RRn78pKqr0zKP
RiFg4orRG4j5xSQekJcIqYhkGDOaxkw+3lF4NZvQSBdVr2Q7OYZqB5r3y4GZWgnO
JQo8tALRW9w5Zm1aWgk6m3R0JrXDPrM9oR0OvbmMsUj+hwTcOEfvG5cAEmcgqNsW
5R4AIOIQhXcTKBnwsAd9NW/oWSWAkC0IHkuEDyDmIMz3R/NwWoK/yD4zJUuo4oj0
1fvgL+Okct6np9Cr/ujerQOmgNbBuPYUWeRul9SEr5XVipGEs36qKzFkFBHwhSsr
gofrrmQJlbCTJbAO+YOmBAiW7DTidXLfHVpB8g1bp3rUb4YS2CadEI8YWVotzC9B
hJ0v3GVg6LQDdI0YEos+ajHOopLPPlYZQL4yNUIPgjSGM5hd99kUjH3M8aYNQsVi
wNr3SHFZ13nSltZc8Cb+eS3CQDLbAe+K5+8rthbgDx0ewdP1Opmqi9zyggKTwY/q
lXFPkOk4080rMhExEjlJqohhV05WfKcO/wsTTHLYPpX37tZ45FDVkf4FINPsDm/u
NYf+x+ukDN38iIFcFrmDZkJ+r8LMwUti6YfxqokikaYkaDw+BH4P1hzd9GI50SUq
my4TnzXCJZzOgj0O/YRbN7yQ4u9FhahuH5FefJe52DNqxaluTpInDDZlLDW42sBn
OpcLWoSEyX95o13XWKnlqTaIHDm2p3s3my/d5MyRrqV6lqthG5PKKC3tJnUJZ7wI
/nEMd9RHeV2wN4rcklJEPEq20FWjUUVPClCrNajK1y5GoaAInPwfNMmmro3W7eio
Ydu+1AydRw6bXj11EtVBQzaBhQkCyV+tEPIAa/CBWzGoA95R9ED+1dIeYoHY7XaZ
tvDaa+KHeZX9b5CYhz+OZPdMEspOrT+XGJFH7xKqBQEvMpv2pOwL5bDQJhTTVD63
AH3OBAOj0eqyt2toot6N/5mkByGj8vzboQl25z37VJoaocJHpDLiIcyPqDCQX6J/
dRZGokdR0SqkCUr//Byqom/iZeX10mSqnXYf9i3tErYFES/IGu3qNYy9hICKOxe7
0TL3ARghDIssmwl9u0P15K7Hg2+1QrjU+OmiGJOV9RnKDL+bOWW6tTYod2Zq9syj
fGze+yqYXg3OoArptXD4wySmPfxGEG2wfB9hFKAEb0Y0GIVoOuL85RK/Grq6ChUg
AvAXWS+G7ryZ0w/sI5S0g+asG/P4x/jv3AXnuHgwlXHZjwKG4xxrx4EkE+K4dVr4
saSTSA2MpbaDhNRrNeFj1o6Wgozus+Iw/APbJn/v+cdJJPHAfuZoFQw5osRWHWlp
3DkmQiLhgVoJubulGrOLeFRuwD2DbA/pzW2W7N2SV+HKpvOeabnUavQqx8s4UbtT
ixOQDFUY7iGZcc1IwXCDYIdn7EMnoYm1xVH1ddzcXXqJ+1Kpd9zmzcfB/sO9Ea14
5Wj32ptysazV18CY6mCpr6d1xQ08CJBZ7bPPuBXF0c4xjjvAf/7RhTbdckPxzrZc
/EES55IQJRqlvs9uSRbXnU/Rt0qGybq7VMEO497tRn4rg/C/FH4KaYBckICwNzI+
a6LHFEyVZbu7LHrksF6efOPzLS/IwgQ86Of+oZZkGiAOeaDugQJ+z2R2u1XH93qf
PUO6vJHRltpFwbs1dSBC9QHRbCJn4gtmarSD5I+XhQEohSFFNuNbEwonAF/vDO8d
ZsP1Zt8xSNTHhYhSgj/4+oMi5+5Lexvfx+20L4pEmDfI+EIAwVpdIuodb1+S4Llv
JVGHHV8dEj0npYhoJJIj4VyHj2yJXF6ZAOg9S3RQMSlxGby6jxBtrvSmuLdk1M9G
BMQsZcDdMPOJjeDWyAaczAzgMqodv+fkqJXfBFzm4vJJJblACJmHI7YBK/otTrfL
sBskHJR/XHAQz9YhCaFS3U/GwRfPZbu9IXiEBkvfz18HSc0EQ6VA4rg6ArjTN/vK
MFRUkWtIedUFgFZes25QYfHaOEdXBgMc0+0mN5k7TQeanItMbmCwxNXe7nuLAIn9
wzqy/7pQnrvB1aky0H7krxembuRJXF+KyZWIb2/JdL6OWlt6UvR6oXSlNUagoA1Q
qEWFVr1YLFFMYIT0B2vpKbkIOZKLyzz10a19+neBpb+dIvd8d5InP/LFsO3zcwPC
UIcnrqAApphvY+r3Rb7DqIvUX5TWBxfprdn4UqH3Yht4WAdM5wB1HIO+b/qOVSDw
IZK3dO5dTWm9es0vY0YLP8CuzcOz0H0P5jWPUZO7UxZib7cudi6ogEbZRa83kKXZ
MQOrtdGOHJ5+c/toW+4f9MI3/TmbAhVajG7VqA693IYF+ohxbzHU6z7tFLVFqhGa
dQFLDdc5tYPui808qv1e42B2Yr9kRt5NIoxva0oMCxDVGwpx2os6+y9cE6k5dC5a
pZllKCrXcc7Px5hUS4TI2VykGwu17ZfKiEvoku1Sa9ElSVuGpy9geOWpM73pTeqN
UesAGpcc7b1SQbCj1vYEg0XqgkYgFELJ41qz61ETo3vTzvUN1uaa/npNy+l14rwP
fwqtk4o3gHCnkAvi8Yzt+zL1PQhPvxcCpVeXQlCgvdeLdr7tsVj2gRkLYw5zLHxX
l8QtzDTY4xgIjEsjY7wIKGfXJu15wu9YZ4HQ+0FIJK1raY5pfPuJzGzxsERZ013O
Z+Qj1fT3mC2ezMPALCXOz6TYikY4U28dWwRDC9Y+a+Tygwnop6njf4X3yF/CPyaZ
8psn3KwSU9YOSOrkUrPB98EOlpFZcuKyaKy7RyVpfMyLyCuDe5ts5RAGDaY7rZCk
WDWunyj6FX9BhTDzpDwQnuw68gNVm+/qAEfYZOsD8Q+nUVuZGTPgNa5ensZt/vI3
0RyUfvyeVehNGeWR01r1IKQSjYghbDJPTe6n6ebLpm4xC8pzJC3wzt748qaciia4
rGU554yW48nurT4w/dNv2wO9wnnE7aEKHR5GX9EdwKKnREu6AZpxVLfqp7//jDWO
rlX1iSwGgQOQuvG9EXX1Lfgd9VpafYotBvrrxLcgc1tGWFFlu4sJUDxRyRjIK9Yp
3ZrW22ZzqAGOO23dBRYHGQCS2Reo6bgOPy3BMIQLaB8xVjqsW8jqxVrMhc7sPVtd
RgrXN0gt3sxMEcNnt4T1Xv0F2Qb3TOn1HcfMGhpi94WXSWrjN+kNKVnQ7dzzBuLN
HenuVO466QGJtkh3AfNMK7Lgk+uDjxgfqHJWKfvVrjHFin3RRpYntLeJV+OGP9H1
8wH+I6E1Ntnd7UamF99Ine7GSa8qYhxjCM/jd8iEGd9BIAy6m1aVTT5GmBPCg5PY
1oLStZmXC5pF0iO66lJE2/4AyCXZNOjR7Jnk+1t5jXtJi+1xMqEnswiz730Num46
cr0luhWih2cAKPijNudizz5S7m+xYsNeTahuySISqlyRD5dhZUhDmRhHU47u3XyC
xdc9GsK/3qevUYICFtxuBt9nrQ4R5T4n7buAHo0ms3RGp0xFtgB5az8oNtw6d6aB
+pXHbaXfdBjG2OQXUQZIA3oBuWaIhYIU2Es9ATNII/wZ7eMFvw8VPUXTUWDibkK+
BhCvyixhn5ZhiGIuPY02UvDBDHvfUFI+SkTsd2ehjytprX11nzTkhgOgSWP/uin+
q8Pei7fDHlrbeerEyI0SyhkPT1qdH+MKoBaaeHgMnc+wQhq4QaeQp91x4GEyDHI+
uaWyuXdLNFxF5nR1+3UZrZQxut5cDs3RTOzxl/amIiZud8dnTqrEVbUREDLy5qYM
HeqMytqVK+Y3JsvrfDWze8+qNVpUFjGsb0L6knwN3H3YYQbhVCjEUJQejq/rdnEm
i4WKc/DqBWjsnnvm+3a1wD1JfDrez3d1CGjNIlL4c21JuFPfqWM7c/J4KldmgCNw
WEAaRAudVKR5VjBXz8VGtbg/Tu5eRsHaHpCM/lVvcXguttWDpGMISeL7HGV3zAkZ
GnhcIT1jjFGTogzXm4ziSGUHKt1uiPETCStT4lvzi32mzu4SLqeywmJgUsQObOjC
yG63g8U2co1cQZJ2JedEqehhMnQ99r3Cp8ayda/TyM0burcZJ3n1nn2apZonAnSS
R02r1gw51CWHPfR0PCZD3XOZ/wc2F/0O0Zh24yDQBnMh9iyaJXncFozwEgr3KbgF
qtBX8lkt3f0oz5/o6J6yTyFbw0x1JzwnSuzJ9+L1iGSuDHPZ9sQHiEnwzWyNpzV0
+5T8scqR10bFU26tFe19+OdUTH1VgGqm1++cq7Zi29TiyOhObB62eHt89+UnKTQM
Thf2WIF8oDWXkbXfLv5Y/Ek6wFD+0czXFrBmZvRxhcZDVSjOf6xZ+NjuT+C9q+ku
SVFFgOygTvAma/FdI/KjM8a4kv1UvOe5WNyDIatUTcYrVbF/D/qFT13yhtnWTZ7E
s509m/zKizfraA6P2q/aug1F7RD/ghVkiWYk8W8HDoHQCf+y6PL9U427mxPuMGAd
5OljwWP8Hq5yM8HEN9zae9RAXeUhroKYLTQBUVI0J0bMhXoaqWkSPlZ/vQKjzdBu
hdtVplAY8SjcF7hs3YdEykZYuxOJKbAH0zjGfyGeyM4CEj3G57tNnyzaVFuefHLf
vZb81R/PSeqARFrt9q7yJFEaMHxbABnAZa07ah0suFVrMQ4A9uaa6fFmTz0sWgfS
RUMfnZceb4/8gGv7ubvMrsedt/0NsW8MpIFfv5t2lhrgiVBwHXJeTtexXFOcv8Zi
q8g91sIJAMN98BMUTyy2FR1KYLzNXzHoeE2yeZhkX5bWyWm8jUwO5Y1vlIFss/jN
Qac3fkOx34H4iPm7wUIQ3t5syLhJBAtzAkYEaQjbtiGKLJku68+lEVvBAL0nfdxP
vFgvsFium69x0Tp4EZL/bB/gE/1PrXli/azbT++Aa9gOO74eUVvcJp7BxE+XUnHr
VALaSdVJL0VAYUJRk19gzcE0CykanKcCKbvz8MVhFlVVDsOXZuPVOTMRPSVCeGRy
Tvt0bVKcL1ADl2mEGRe+SSmVI/bxAI1040ztTpOtE/zXzp3E/BhLT5sqD0qJvPsm
Eq6KbTheWCplCU+d004ZV7rDfocDrZjdJZLsFfbw9eYgXieHntiX2EMQ094CG9G3
QcNiSiNZ8yoHaCYb/kj7ovRhgKk2TZfHpbh6K3qDHUIswcpl7M0n8nFb7Q92mY6u
asbdi/2puRcd9ditH0cyWhYTRip5m16ZNUqqhsk70LqAvjStxv7rDqeeIGsV2eYZ
CnVoKnxY4rCKXj4jNR5A2p48KM/3JV0fKrb9WbWR3plFJBaRqOXwBqBdUkbCV6U7
UViZ3qBOP2gXWVEQOq8xo4nU8sSOZlPK8EM/sLWBbbu0q7ayvL2wxf+G/OwqOXBQ
xKCiUy7scDX9Cb3JmwSrJNquNFrTSbCvF9ro7RpIIQwzGzvfP6Pl67JCUBiXRyDy
iQunHJdwO5w6LUTw/oXlI4oI7vmP1fTWndiGbhi4RUciyAxNQIuAG2+FjCAMY1jM
gz6ljxj8ciZe6hCEtD+2uetKtxlQ7UmPV9RUrqU6bsweXXtjMgIhFoCOa/mOFpUQ
oUFRtLrtu8lAR5N/UAr/xPaQ+eqMZErrUbBO0yHK2Md7YVD/7N58Hmi7czLW9Nai
mdbjMCm973CtqCgTB9j66m8bIwY+1KRed2x39/iAtza2YY9I5HLZCZSdx6CuTIMh
uS4XFQNx7/VqgwQhq3tRFKNEzcBWMjaR9D6kuqyZiT/4pz62C1tlBG9EMb3StS6q
72gH2fWJNDTRyGVzPfZtdTw/OXHcme9Sl6Up5nZYa2uUmMwHj4AQX7M8sWHkVw9f
fcg48uDEd3jlmoJJAArmFAnCq8I03uxtPWsDPvR9mdffoyw5PfJgekQlpSXtzHVT
33Rq1yl6vYb/p68oRBPWWnlHLbW4Rnl0xBGlnWHsT/6sTdzfJt3ToCTWzps8Sshw
9wVRD4ieXsCCwKY2Zkl7rGZkByMRzAGfk99w6BretCLofy1MNmrpXytCmBFJMBae
JgJIo+TNEc2jHzIu4q0cZqrwiHIlIx9SfHJPK7J4r/B7SGtxSpZ7m6b6BRxSKro6
5qei9ioFcl/U3EFEwL0TL+ShWmE+uk8zMrs6HBknrAVCOD/0ncBCs+8DSTTCddLD
S9ARRTwJnOzA659dc6+BqvTessE+dmap7x3DrOqYpHPUfUE8F+h9ZNv6bjPOhJ2w
DwkqmQxjhQfD2kIDoki6loduaFgYvPAajtvhrQ156QoK9wJGo7oGSJSx6lZL1FGd
PoYVSOAngLnsnZo1uVNTlHNjdH8TFPluzPzO+0RFkEex8ZRrTrEkZunC3OQZk9d+
oCq8sOVB4WVYoJUeSwKyYN247RRHxiYPo3ooWFncnHGeYsomj9XPgESJgUX8d9oJ
kFHShMYKtY9NbTN6gF4+2DYju+1+59RpRtcg+JNNjA4z4ti/nwqYmgfPjq9op92l
0eWMbPEWNWigqdt5rR+PB6NlqeDP0nVf7aX/SpEMr9GDJjfTYADMcOX9pMJjSrYD
W/5JdsojPlS/qlduM/sGYTVL8QF6i9J+u1t6HCGUONuuOIRxM7TDFfRnYCa1o0MJ
OPlv7MLYJewGEYsAQ6VGJHW+9v4z7DI7/HdWsIX4SoEQ+lQ59dBJe8Dp9wfMKT5d
XRDMvznbTKPTK6+/qlQEygYSr4CQ23lTLFsbmyawqKIm9djv7ApcQu/qDSHTlVL/
cIMmA7stCaDCbUC+k56Ujb41ATYhlubdRdcbv+c9oCYZsJXFAnCfHvHdGpcH5rrU
1qpPpJMI8bb2NKxqnLpOaH7athIKhBW8CE+HqQsHsUNrKmygnn1oJUqbmhdzaQSu
zKIvwzcPxEo2io/1ZXANnl3A0xCr+7sLCDBji5FZs24dz9i9rPpZHKOenW7Ryn4R
+br0wZx4jkitcTuvaPEci6LK8rrwHsDlAlorKXPJ50i8inFO4HVF2BXSxKwIbHeD
GEEeaZuMajHL6tnO3+8EcRydGWNQ+b+/y5ZSrGeRyB/daVGv9fEdxyb6ZLg5V+CW
Xm/5FrH3Tprvk0pAPm+hT8hrz8kFpQa8izjiZ03MMUm47Tvf+C5+aiI+QWK79vcI
R7jqwxU7CDVFXUj5MPBz/4X/T3m/lk5WqXhuYkVi6T5tM+a0QFRhmxFcmH9GhnqG
VxnUkP4DQ11IPDCXYSpSqAEq9yNx4Hf1OEO09I4tKvnZmFir0HoomipOd89UtNAX
pqwLCP/lhSunb95V6oSlcFH2CtdeCOHpR/t2BzWjDuBkUHEtBFsMTIO6+YZ5WQgL
r3lpJZETiGmbtG8tM060TjLt8P6REPuEE3h6S7JHGgXBpZDxvvK1VP773mdhsU9T
lGCObMQ+E8DeRvneKTfTighYrsJNqVG5l7a4zuhERclYWOkbiJmszzr+UYka04Vn
C3dGqD20ZQJlxb6pRq098xOoACT8trLz/oYoRPVsWtnqCnLgn3vXpEBAfsvUinRF
AaVWqCGLM0EKTXXHefdJR6W4CtJo35IImhe75SgIEZbbjFjS5KGZikSeMpZPeUle
sm1PWbapoxullg+3O0/kVhfUYbctki+OytuCTee44kPDbxim7N0837AJuUphflz2
rWKVH8Gb+N9XzURWQvBwmnSRT2u1J8nmVjorENczab2EtLwim+qjYA7OeN2fVIXC
D7Nmd35qybs/5ysSXO+R6Z84UtEqdFcsz/qdiTZu/Fok4jEoNjjGn49SYjjI1fb3
cqXARye+vdQ9+x9BDkkG5c8HzaOMKYuX148aZgGpgsHx8JqRI2LWTayqm2zKaa2q
gfsNtm6LWmIlS0mxBNNP6/rvmZen8pJMzY9MaYculx6Diu/GVBn1ybG29LiDvhmR
RseWkbfTX/zNg0qqPEUFvSbVxO4Pl/378P+N5kmppV/RVgY1EYSkRUDbD9+GjUin
LtPPTAQzd6bLOQJWqxc8ctS1S4fa+85obMcj7rRCiYiiuIYj30KbqtZGvqGV2K6h
PbB0WTEA0miFAhazBuLjgbLNJkxOZ8gOq2lq46q8JTPkZ6oyJKRogX2cbaosD720
iRDqqMHc0JeWndEmecMwI3CBqsH3CE4qlFGdyV2427Q3cuNU0A2CiT4mCpQVbLaC
GqlTZrovfEc0E3JAlUHQpqMfvOerV8fF6LzTkS2xUfGUGAfE6susxdyjPKgg8FJr
NEh83hXpDfubFeyu+CtKJdPgf/zFhUl03HJXK0du5Gnfu5aDqiiBAtfmZnX9VlpH
0Br+Ds91p/yW5OxOPVfJhW2q7mPGJrQGtI0jUeB8VnkxbHv3dzp1sHc/mpM9Xrkx
5x0geW/d1Sk/xd4WaFE9WGcrEKovJM3ie9FA5fVHxiC5KAqwLQ4pETKk+hvdj0Nc
sqDqlunu6cOGRBY6kaL07M7QorCq0L5iqeAt6e+VdrdUdKC3E8U8DRjead884lTR
Jo6XbaMZKSRRDCJbY2Ax27+qeoe/MJBLYgog2uOloXlkckQ/Old2J5UPCDrJngmR
C6stVwI+6sOfy/jrjvBHSEYimS054NaLARJqNEjES2cc8dX5sV2rPtGDZ3OaIeQy
TJHrnhnQ0ep5xUCzXmUGLtLK6hFdWvPfNvAlpeuwnzkaly/P1YLpXU8Zws/gdyZq
B7vji21xfGgWx7Sev17V7Vl3dJiGfHEXCMzHy0I0vJTX5Bz7BUiIOsWmssS1syWK
Bvr100NiKRMQ4shXYSHdEENu/no+7kX9mm8wa1iagu7QecS/8V8zQbplJGAnU1Aq
c4AHcsHdITFIGCbJ/YXax44iAfx7Pz7EkhFuSK5wCh/p62SYkb7WVv4Kyp+Gwg3N
4iryrvv4sy0qXHogx9+g0OjfYXOHp5R4UZaa9liqWgxRd+EzPANAwZuJtna5tiVh
4UGoI/fNc7KSmZpTQbpMJx2xxRutuX60Q6979xPntRpnfJEa3VLaYLOtkZIP9VHU
dhAp0JUva99mqUXs2rzpcwALWpv7JML67JwjyqByJo6iOPdVpIB426CLVLTxvjvz
FtIc5X0I3WNlzUkpZIKAxShm5lN5mabMnezKmraTT1aedtYRDzPJZT808O5trTCc
Ob47/JRZg+CAzCZVHgeF/xttdkr6iU/Jqanq2muG+E28VUduxeqpdx1i1TWTZ8jl
pLzUx4NGsRLdlyWLEp2h7j5nzUE3coCZzPW2kBvMo+RpcRL6qbJHjC7yR+HPZpIa
fFCzoAHx3mt+k63uuph+ctua8CiVHPn7dG7aa63DmTvL4DaXyGZG32sUjM+NUh+U
h8Dx7zYj+NVqIaffNl8nISl3TvH7QosB5/LM1l84x5tvhAH5NgkT9m19421v/ooJ
olBjUcjTdWpLkkwELG8kFvNuGkxRUEZaMDOymXe1VluwcfAbigci4BRkuvkx4iFJ
VfBktQtfYrNNe46UBINoq9BCxEQtChseRzAMezw7A/3va9mPrITP+6xXu6RSr/n3
teLsR1xayvt02nKCXVJIew/FLwLA28h5xSUbOH6i2h5d3Wf9mr+rK9RKDNKWNzpl
sy/NV1QSR3lKf1ITjkUP9mT7Mz3otun8IrSlA/X3RRa4n4NjmN1zuAKzPBaVrSrI
HedH+0GnDUoptJLPnlBp5VFiLukxUL/HSb3HNF8kkrTDoGDLQgVW14ElSRol+G/K
zY/Iqv0erZ/o9NuqtuabUswnXeHdVG2b4V+MJs+33XSaQ1dFRQD6DjOm9AFkzTtd
JhS5FZmctjCIaZWWOpFd3WTBx6vard1Q6rRiU7c3k7zoFPEJnYURV5Oi/XiuWsLH
HQizqrWgHOqJPWFMrnHMhQCXQKpl+NKICTkyXYKV494UquwMSHBZEpGarcVMs8ep
c3rET960S7d7SjA7Jfgln/89MXziA912pSsbC1ulKE9ltl2yjo3Oh7OQa1eN8a9e
aLkyTcBugp5qqnxOYQ0plIOVnyv59tAKjxS4W98n188dHgqhYRX45fOG4qMUJToA
3H5vNHebV9eZMnSvdT4h8Sh/Su43Cpxus1s6nNBmFyF472HZzADhYTzLzRIH1AJM
TPh2hLvAqsN6ahUPFnrasmtQCORBsPg6D0G7d/8K2Bjnr/mJA6AafvBfRqc3qsGu
8+d4rvvK5lxRUoV0CCZOaishHzsn8Es//tndv6m0VgIaLEeC6loTC2v2FMZTEMp6
wJw5KR4AxBVxksrCRV4/bmv7V4yaynrEW7brU7r+FQOfAibGrgcaJDW38dyRbhRG
dKJQY0m5S/LXXpkTqO6M0RTpam5CRU/yvm3QAAp3I3uDDxZedSUBgabOok/UhImj
VIXUGIj3X0tmnObz/fEUF9rhIkBYgXwyYEmACzOEnbKIhtFc/nmuKGyliCZQdoVe
7o2l2X6WaajNbYe8IeTbABewHqY2x6vHqEO3ZtM7gaFVhT3UvfqagKc/AxuZHvDS
sU3hj5v0UPK8T7bCHygZKQnkDlLlc9+c7K4qf9xZOk+9DgsTLHtYiBtzKc8NEl/E
09cxXuDFRJ54Rqqz+EAma4laEGShb4StbGyN5HCCawBYLtD92BGVDzHJTp08R6+Y
sjGspYo8YaECVFE5ebFSYAa+pxWGzcYOqGKnfeYUU2/QJJYOrFEQaki94X2N85Uh
njruSwhS3KG+y1+1QpjKfgXTSKOYzWEjBjb/Ed+65eEaB2S8/z8fqs2G+Tbrj379
VZFENBLsxvvR1XFMeKEdxKHZz9rNjvnCDmKEPQ/8Rqtm8p+In7Kf05jLepPocviV
VBKSBBVIXFUWLmfomAu/WdLSB8xC0i/VQ7y0XisGaMDgEcXHTeBOoRPbL4x0E3N5
VbDonnrVp/gGNArx07sr7FKmjzo8nNwbl7sOGjWwiKtYn8EviNa6grDPlCUg14Ub
WK0Y/5m2bSKNJMhxuXaiBVTx1c3WD3+XSTyoLYyQaOV641psrR58+VTFln+CVKJ0
mE1DvX1m8HLynghmd34152rS/g9l2c2e24KUkyt1vRsGODeGc5DbaptjLBVBwz8j
WIkSCs3q/jDhDuzyj6pAR5duVtGDk8shp0NRpeXXEjGI6jGGpgePRiZ0pApUDdZN
52ZjHASfPD/eK0mWSufuL3Vq1KF+aIOAiOnov37oEIWPuTf23BvRkplKXswXBCKw
Zyddk9epR2ZttNJZfv24nk3jb8cd1uPumKSbeQduXQrF0jEotriMyhWR+sDzQT3/
cVIxicYf8te035l8POoiChKZjn1qGGb+QL3RERgy81ZaOF8hWtILmrFyceJsC5LL
XGhJgfUc0ImLJyRgGAW4OjeQ7xlKvdv1BXd2+JcAOajX7jq6KZDChLfucmIasSnY
IeqgWJK/TJ6s398KpXbkNR4YeE2Zo+sfBKYNKPSJuyy54E74mjM2wzp6lcUubWRv
brmrf3/gQ8hLeMMUmqavXexqHh0ovrN3+i/APLdHTfSzg03fhwgHGRhxOaBK43tM
nZhf3tMN3hAeBxfudCOQ8096mNKZreSMQlx9SEYOgcPVlGgXuh+3nGgsOhkxqo+Z
wrwYAHGxlLcdVZSVEiD+9aroWckFRpKzZZgejCUo8PoiA7Pz2T5Q3EJ5isJokhSL
WrG2+zi/Yh22PNEsTqy/lkP22+SCul7kU4HanTiY4QKBkqlXdNCtgAGuEDgdBNr/
zQ9ctCvP+EN7xVs4Utr9RLfE34lXCQkkQkadOKRFR8UXKkqkFppT46AHB5EFzmjh
LnlL8k/Fwq4tP8/9SsPYxyWHbE3kKvUH1qOe8lUTOBhqcMkyitbKH4+NTMNKXnFa
pQ2zTnE8x6FMxxmGLtpr7P9gafjKvE5vB0PrnUlER3v6xHPCKEiIISKDiB+9mfVx
53yZvbh3RSn4Ibx7Lr3wBK414Fs/19eWFNzls06dvosEjPB5dYWfzcB3h+oJyjGa
iddtgZPTePjexyoRSFtrrDoKSpXB5Elx9N4yJyDwGWvINa7IZzxUBZpFtUPAWiLi
lkd/QHrJQaz4X0Kb8SjqrH1DgiE1/X0WUB2SDazJYMyWEP703lQ/Yz7xbCB450hx
exXJdEH3sPxLznmIVTfvgb26p+eZFi6+t+KlWmuSrKNrd4A+UGYCdHRwA2InNsYR
J6/S3PPFscd5G6UPMwqbTGLfbkSo3hTYt834XT9XdFByjUg5wjW1syWnhfVQKeb9
0DYifhAN1eyeBmPKfFidj5jrgnbGoqulXC7TBsMS2GZIaQxtKWXxpRKyIs3fYps5
HGKm/RaM4xVoTwPzPB1Yt23whbqigcjokxVBe3woNrlvEvbc0debk6mfE1ymexNO
YmwNBcjzNjWiuFnAa5PgDNlrQprbAOYMyy7g5pJ7PVTYjYocwwYXmlKDWu6PG9Tg
9olnly45HJCLqp15EeV1kEtsXmXxAXHnn17Gr92IeERh0J3XBbKHQseRlrO+UoY0
CCxJzRl5yWThoIeUDCa0apOZ9ofTJbUlTf1/b7J1MyFL064QpbXWBr16WO5DkWt+
iyQbpzxNWvccuHBmL6d09KJsAuv0S9ekHffEipVL3JsG0FH6uNiHy8Iqzreep4CC
TcvyHcRHQhr51s3ZUNrx39dEzTlRIXGsNcRgDpcATwDmhpUr5d/wuEGdHnRoWubP
PvI6/vIDKWHSWO3Nez/862T5EPW7RVnuYa5+l2Wt7OYDaU2Q3odeV9NN66FEN40u
l5y+PoFOuF3MXHq54xPsbp1UCCxYh2bDGOgLBQqAcmqfG2uo7Oin0Ew7QLv0FKZW
sw1z4ZUuSGY5qi44CQiu0xt26BU1Tidur9lL1kDtrXg4DMPW+BMKsb91YfIaD+br
lW3cPHc439yJXa50kf/syWwxIMIob/QVEbwE5aW73VIBH9OKzsfeKzojo5IjEDmb
//PktqZ4itmRVuT/vsP2Y7fthq2dKmdMSz9tYINQov0Chd7naPjKHYBkJDgeRylJ
DoTGAjDfHtidh5xGWeRaXM1iv/2vh97WJeiwMt73C0YutTbOggAuBWE1qZYIDZBo
SuOJXU6M9+IpT/6yP/Iek1RMO3ZN0XJ6OQgM0LP6LpWb+Cj4S+bocf8TErnbQifQ
dvxlNXmRsRVHgQGiUkIyVM2cLX3J/K+qHAc/sXJm+NXZisiwJOsLxyjDxJPtZPds
T4YI0QGwKcGN+/UcG0v6NmHq8PZtX0Z05xFJUngoc6anXuRrl6lpVK7rXO8jPCCx
9UQfkpXeaJ5Cn4KahUyifeYRL1/2CViBZmgpZLc/0b3ds8/D+0A6hEDdQKB3I6ej
b2YvvaFn2+n4N+3GbBkApI43yR41oTAEu9wG7swgxm3Y/u/cbpk/XX40/iBDvm5J
Nb+FHW8ZCR/hJF+M8kWcscK6AsNPB5AvOIPJLaRMxhAf4/eilaGtsanXu8uMti5T
CO3tSUiHZirX4cXXGOOAoqDNBrFKxmqIpB/i+oEOL9uZ8IJtBg6WqMHy3BOTFHeI
2bnDKxJjftjb27TkO+c+5LZAq1h7pF0mYfKorq0+voDzyS2fzi6Fmhn6ATIvaNy5
wa66br4PAntGQAxvTFb+3NYvPrReITR8j1fb/tVh9Hp9JBd4h+NpF3p8ANeAj9pY
hiRKFfPT4sidzY3N229PTvDtT1mD/z78zh5dfvjesx/t8p9nQn//iBo4qwhevHR1
U+l/dQTfUrpHLLMkav0DcO7P5NmN5/1AREpGRiku78y/5oGwzbY0nLSGOFN2Fv+Q
pNOGH4Y/5dbdxmGLCNP6l0U573dvPIlEu4p4iEQjf1PMxtUc+0AxPCa0c2N735o7
GTQPehc3MYyoWKP+NGodm0XFIuUIWoOmuqeNq3Dbog+nbTJtY3N6Lqu+FXSJPTxS
mvSp0M3kPF/v5wzzVe47e/oPzP+r+gH8J/S5maAHVOUbJLBezYrlzQ+ekjyKmhDu
IkiiaczU3q5Au+t9qBa76euDQ4xMuIJmm7cas/Cz+MazU8gdAhmOAvIKjAE2o052
bdBZq917MPNtA7L7lj5jbI+jnn8YL+XIdbw6SeFrhnUkbUC3lo8QeNTdRgM9NXGw
aNac4U3fTjlKb2ZS6CwRZoT0jJ7peD0vKaWg2IwtynBYY/MJJT5F9yYMY8XXQzlZ
DfoUvDXCm5JhCegJr6/WH+hdUcR7MRiOGd6ijfmLR/yWQMYnjkK7K0YolOuRqGIK
iEzPL5ICXm/wXs/xhDOJXncqcV+JVK3yHFEdP3LmFanerxd/1MHOvSOV5KixxWzL
Al/6sHE+DH6pr0BDksteFWEO0z8r/u/XxX188kwyTmHPPS1Ypz9nsf3XIE+VX3Oz
Dh5PinrJ26JcHzD21a65bIA8Vh3YeIxItWeA/3BOqsk+I+mksRRUoFoiFh9ihGvZ
RNJaPLU0tj8f1Zg8zgx/k1BMKfjMmwSJDZPpjnvZq4b4yMPEdN83muB4/JgN0jkt
GApNjhhjmMOqvgqmtckuGgNgAybwaAFyZkIHriQcYhDrCsm1ILCciLfvzN9ZZKLl
+/jrCcBdefwWh4QxGurfe+NLfNbbBGp8OOSd0pRgk8B1ahgxWxXIzEAqVK5RspdB
bxlpJozAEOE+hUMtCQ96Zl9JmOs2fWTfBOM4+1bFfowRxmw5Vno3tOkj3OLxHaMB
258qUL+dk490f0Pkb4xq7spv+JtS8ojdp1fgOuTp07GD2Ilfy5vGNDwBd3CcOIlg
cyzAE1oIo6ehZKz79+fxMpR5bEYCtQcsqk4I7RJDGO+Y4nE6bCjEhMQAX3JURAwB
LWt1Ly8I6/fU7ie/zMEYpz7XEqnk9tyh5mW+++cbXFGGc2GNY0zBPck9i7OfydaQ
IOJQ0IOWjTE5Zvnw3c7ADbPZym1HA9i1CblqizwpOz5mjUjezU79yBR2kvLT2vhH
WqPPhb86GRkxahz9n++iw8o7OjeI9r63Bl5wEugHJSaOzheHRT09iAOtK1Z+kT6p
jvyqtP20LYxwGHSvWghBzhWb7KcD4mOg5dLYUheHtxyae0DlboZbpylf73WYmKK3
xH8f9rVzclcWnqmZj3E9FHHZI3KmUetWTz40MbL5uHKsEcymcuYZvAemuHNaUTpw
lIgsujZfJbJIpWpzvAXGwg98YcOQntR5yUJQX+zu5v0yEWmi9fxbF2LRMV/HSzed
x9+AZeTjrcpxJ6I1WCeG5qAd4zpCUmoAEiwpTX0JdPUazmC3ZVQhTA4uknFjB628
hC3W3MyZqPPHSkVTkppP4rLEfVsbE7rq8o5c6HmolWZbwDepf6um57KFEDfYZy49
LRFrt7kd/8cvQvXTyd3GFMCLEXokxAkt+gwKzr2sUmD7ZFcvgKSt1S8hfzcW0FV8
7Ev/QptqqYBCisSv28D9OfG38RrIBS43bkVZC0wWxFITZyAWkezBM/5b2kjtz8cG
8RfA+Ec36NJIMaHpWzvSNNnajZJHzdq+WnV3NKvzzz9sVQFBmlXm2eNuVMWxP2op
LbnNP8ktbh4hw0ttKnoVO6/tZ/TxmTqIU/z+kYmSR1ZSTJWblPr4HXDmHeUxI3lY
26R5f9Mb2lq/go+5Ij7gv3FcGHoi2DfgcA03RV6omnoE1h02YtPHPVsIiZB4JuHH
gv+7cWi07g1W+5GeMU6WiuTKzzMBKP/LjI0dKBLYq+owFjp4rYivpSTCTHDziysK
rjoHQz/OVxvg5cpu1fyxU6uFpTuuM1O6hYtNKeoSRiMEi14YSUz+3eB/pmN4sUPm
QJL+IHTNQ0hUGvADhoW1cYs1O1hIl7AkewqhbRt9gGeBOQKuA8cMWIPKEkWnR/av
90q0FRBzmEW/R4rsBgh4m//Wm+MoSvs6XV84SXi3+70hjLEm0RO6ZtlFanJsWC2y
4cwPZYYKA02S58/d96I8bgk+7qPNBqLEJM/nPsZJAHzaspnp4r/qelF2YeG6Rnhm
XNBxH18vvgG1NGyKwUG6XpF5lAHZvL9LMOXIuc8qdaYeAAAoJ/RwoCvxuIBeMpDy
OWE8JVbBdfymA+PeI3b24Zit1bQXS04dUsMhgLT0QUMM5Trsc0POCmeXFcOzR/P2
RKnK/q+wEaoyRodyfqfKTiP3UqGM5rJwLHpim7ziwmJKTuGKxfauLAiMjci56pLb
L9DwL03SDwHoB71Q9Il2nScTiOoqZYsuzgvJT2Sbr1Hsbb3VG/9AG0Uqj/l2jFS2
JpVgrgJ54gA5xAiJQ08goS1PadkRSdF2//w5Aa70p7fr46Oae15yvzzODijDHSiX
Z6jdeiliTU9xpvQqh/Iiab0oO02wCGhc7KtHBM4RERUMHgdL7u2xaUSU2LcPll7Y
/OIBOP5KfKwIESxpm9F2YYPciNsGO5KlRdYP3vp5SSiTmy26jU1qIZrslSOG4TMF
KM4gc5yj1anBhp2Ufx4PGbKRP+CNHaVMCXJLmDDkJKS2lU7PW+8PHG/JmC5qbnPc
GK+pEQe6NAb1GkgHTYHrPJT1gKW3Xh/AN3qMDhfhoob5ltvWxhGPITYvpqgVhi+5
GZh3AgnBGvr6wTV3hmQbtrbx7FhDWUTZgyaNb6CFDiI1CjbBHPRfCcCYjIlBcduO
LYFgNN3aqm4P9rRwRHwFjUQP3mU7gdyiYQG5iCdS5n36FM9Wg9D/1xV3kfcNwY+H
TuWNlI46bVo1L/GKoLBzcDQmnYjQb6XjBQ8yN9jAw5GMEXaGiwA6aYKxmIgu8KcC
sgvKkb/ePwosYwxwBZ0RZUpE7IIMakpfg8weQ0YYN99UiqNUsuJoIXjT2kByVBml
wzmm6Tk39sIkvX3kEVEj8Cl01F+oCE6Vs5YQuX63ZbUglByMtuM1yVPhuXE/ag5m
05752D95wVlgtOMcv2AidDhGDK0t0O0IahY1IDf/dO7fFITjMYqL1++DkfDPiCKm
xemtoQaMIZmMdMOwnGqQj17BD/KY8XMHZUeC9r43G6vc0/IaSNJCVppwqfKJhNTD
UR+baVZi596nmtRiT99UNFi0Nt5VYAdkA2/jchiv6Fpo2po3berQyUWoyEc1rIBa
izVkEEjLBloN1v7/a/r8p/s/hqGCH3v+9CvNvVFxdDza5FIHgaeXLdlBCgBk5WhC
5wBx+6yri3rIOmfMaAD7Ew5q3GW46KGlWNKWhFbqdj+imPYj4F8BYD+ldRHWu4BH
5eW/GLGYkXKui9SF/zJhjcOB1zH1DKSX0gD/AG3SLyjQpgfXUMuNYT7TvifjCreg
hJvbpCpMQ82JFj07oOC1At1VYoqWHYT9f+eAJYiX3UtQFXdwBcG+mdB92UPXOMXg
+nr2k+d0fE8An7pyuBIG7ftcZ+y0mE5OCCvfoObnNE2/Qpu7JFR0VLqWPyvVAT2p
D4YyFok5dWwAHszf6K+3ZnHJiCjvKB1rrWJ4zWQwinwnUUUGyo+ZkSdzO1LV2ovp
WjVw6T7vm99PA0hnZpy6cftsScvZKcwjSr6MKGmoiBQj+fihGhzNXDgrntuNjhQK
KYwCnny2YJXYNxqoDZzFUiKbqSQtH9IoD9f63PuOquJ/hSUy+upQzHzUYtWy3qMB
9DtWzbnNjbHRa5TSQ0IGjEXhtamtkW4xVlw6aUh7BqahWYXhkXUEuiKaSYa0HuTN
DwZKy/W/3IVm1X/6Cbyy5Jki5AYJVZ+S/iWUG72un6ww4a5vGYAvj3s8gFpJr/rj
2hzn+3Es2X6Yc7Z5MsFXme9UdZDbRhfIeMk2y+Urilgt1kf9RgZrba2kvzyCN+uh
cHu76QS0qhz2Xdymie/y7/jP/ZKY67sMbiBPjMvYaO1D1fERNFNVZYR2Z42V75Tn
9yEx8e9HIsfTTL4NbdUZzhDLyd3652KC9KlPg/+Zy4NNE4ryYYCkKQ+5LITn/WgC
sjmeqsrORL3YFnNbGSVT5uxfyAJBy5dnPko5nOh+mV8+bCKzruCTOpqkDb05ZKv+
UO+BWzh9PDRUaDyfZXb7lm41NHBE9XdXt8uObPACHovDW8bfaaxE+AodXQ5uyCAe
iBdEMnN2RZRsxzlSQ1KzeRF1O6EyNVvb3MYWDy1j5fC5/Q5E3XupAAhyByQG47j8
a8JcJy0gd2hOqQlwIaYiD6PuSYGBRLkgyxtnDHeN6RKk2hg/BNo+c/2/ah2/4haP
4ipzRqKaBGkjrPE0BabcInEChuBcCry9HswDYPCZgqIrjZDXqiNYWXWdhJoPuZDR
WuufNy+cdYJOqzpHjytIq+jeO/WvtokaY9diRrd80U7NtJA4GjgAbd7wTtEXIO1X
A2faHa+12QypTzHw2TyQavyUv/DDNp+M4UzDWvTyCxT+SUkTO8smeYziQ8aKPBuK
Acw789F2TJowAiYdwDzCsMtLYx0qmE6LB9MQzSRkR/cdgECKl2J9IpW1Boy5cTl5
lKrdw3FEBbu3QnIfTso0j9JFydYObepjtELGTxd6Y4uwTISuehyrhIYSP0PoP+R8
MHyEBdpp1/RuLOYA/1Rol2a1TdJ61BV0HwYouqHoblkERF2JNq/DMXm6hlbPBqPQ
g3/3/DYoFmKAsdaDrlJIGDZHQxHVHzl3of2s13l6VAVBcxPJfozi7hIGZuvdoPGa
VYYrI+gXdXkMI8ye4yQmkZpHQomGRNGsktayPfnbqRHEOR+0LqFZRe3GdplB2S9/
DgurlMlEsoFQPABq4wkIs9Dtzr5YDm5Vo+rfWqGjoj54vbw2ZseB6qgWUgpGlgcz
q9rnEcqTkO9XX9qezFORhlRBK4XnyNgBGatmSkzlyDlhTZTU6cnoKnuHhh2G38Ji
6hHAIyMWWGsy/BgBuFoDCK273UkCrsTlcq9rMA9cjtMFHJ+m+6hRVNQydKYp5G98
ULV+9j/vK/zpMkHJlinM2fiAcKRNAZf0m2o0N3boE7V5+WVMNLLiEcYfDYpnn/as
O0V3OuQVUMk1JbEJ/bZlCgyOla9IxMt75jlh+nyjC0BrmoqG2mbjYs24Jr44JEFv
QS/Ppc07gmD9XToKUUYku+lYSVKN9rLT7+uaw4HPDO/8eUHMgNP8GDdU/736qHcU
xtRVuVJHK/eYC/NNC1IT0a6CmxkTAxXspBH4Pp2YkMG53hpFVQikETwuhdNWxtz/
FqerDJlERYxtiCBaMgxLHftL2ZampC6WPGV2Jf3uEB+pnU4//6kR+n3K9FhlSxTu
5HBV3Weq9bWcrbYHOXUau3DNU9J0joFVwkP09RStOES6spoIDaWylUouDYYfzL2A
5nH1LsHW/+yE3/E/3h1ALoF5boy1Eki3TnH1ES5azuJ6wYCDMOkQW36thR+agqK0
oUy/xZ6bw790veeMS5/c7tSKpthpKjLn9zz64N6KxPnu220Smh8kCxc9H36u9ev8
3ZSZ3OA67L8wMTg9WvKfz4OQyG8nlWrAx9Twc5z78NeXGd/QJi/W42ImQQUeuTPn
dJko0LYZOQYpTQofmNmk8RTFYWASB0xo/N7i8721MT6u0k9S21sJdJQxccMvSNnL
zqNIdUy4016JOT9pH7Qu/MFcOyRp0mBqCm2qx7VnNy+ot0+pCSobPhECeW10GcLL
TROncF9hEfmENLC8KeuEwuqx/DathdNqe+o7DG2N4aDbc31xTQtUfZO/S4eL8frP
Pv/LolqiJhMssWDbsca2oWHCSkAdEIiJKXS4NFB8HhGGIwTYAQyoGcF8QYRlPjcX
OikhdM0QwV8n2TIfXyyh2qzCS2yr+8OmdumWQhI799zi3NMvns4FERxaNXX/67Jf
iaUwroBzcmyLHEMWePKYG61wflxWJonxH9vouQtHz7zx9UtDNj8r0YmzCf/3RD/t
pcbtE7jlNhbuqPdbVbIARhWNdrkuQXaxrfxIo4FLO4UnTiTvUmBoqnPaIBP3dmZL
YDEwuG0xtv9Iik78H+0Jhl+uXFpgMexPEeYuYziqFN78qE2wjUx5IhRIJzeA/Dqo
O1KTiSyfiekGPVb2JCJIe90g0ot6owEqQqJUbhJzgMZgFAZykf+BrSxQ+zYVt7BO
USPN2V/wH2UvC7Pioo6ZxmCEdHEeVbG07tfx79p8fbZ36kEFAGaBUxntsDG/CZsX
fuPwy5C8uJ7ZOFrQdN56joWU4pPr+u5lFFNOFPZGWpXoVNVerZV9VPSrhWQnDG0m
DUBTxuQHrQShqZEH0LJpjXUjGdN4ijN/M5T27KLMtD4hIhoLWVYnPyPxVhNOwZxX
pdhi3d/v0w/9mCJFiiiU0YxxNn8yqfEnmVTjS6UOlnWmI1Lo5wTbpq9mQFHrLmmN
MvFi+eH4q3AKTuTo2kLhR5tYd0r/YwP+pqAY2r54bejcDlhqIvvLeyAxlaFFG6Pr
PdhLtyWl46/s8Hi6wHTMD/yYGADEdWxeyMUizDF520hJXSBhkZ018VJ/7Ts/24b4
pnu8Jx1yaD+1V0dM2txLUskWu1kk2nfIkeDVGDRZBfVCB/5jcRAg27NCAL9Y+JDI
rjroh1BEcZdxTwhB+HDbAjS2Nwyv9uCa4roB5f8s8qVYX2g1SmYte3gRNMd18xgx
YWv9W5YIDB7YV5JVGDoQvZuHuGaWh+ZYraubejdR4jtP7u3j0wc06IsEow0txmzz
3SwEnsGHYebHeyu6DTb+BwDxCaCGzfcw15XV5YV0/uHail6qQVqEfopOaM5Nt1nM
Jqa461Z3bAaYr1hyZWEaWKY0KfA70VpN/nsjbJve4tNuY77lJRh0qiifpOJH5Hx7
7Po/jk470zv6x9854HYS4Ubc8BiMgaAtLtLX+Txlr6Zg6F3O1Qf59D61bL0PLpGR
MmgY/pSuF0WkYMMQOpOvfzJzBnlcuZOJnllyTjTACaSrL1ofT1GTBa2UEIb6zwmo
kDjI4emCFt7+NYNSTmzfNQwTi/Zvm/rNdDDDNW4h1pJSQMVXTmWzq7X5ouISltPo
kDyGVT3nyt80LWYgktMYg/BVCbljMmGWrhixqi0oDOdT/PiskPb7RUh1vaubQvKH
5W/Mjvi3FtRRaLIwRCqTuE+6XyCWb7z1Eh5YXziBRU8gvLLwW4uXRsM6+Rp0RsIa
Kh1Vzzapfs1eoG9A3nsvzu9Scza5vsW289kfU8CV0DRGiCM7Vl8VAGJIz0MGAB8n
l71I95GoJQUPnsLLqWGu5l8VzVnKcNaNaTPzHPdrAox5Pyqk7LcMN+8CLh+MQ2jE
7tpIpBFURVs06JHwvWLQEkP2RnGwIGgWjKmKPt7OM7zagLEhI+226h9qJRR202MB
V7m9lmz9RrTTWh7kEzZvejVO3BLcAajHGsZGPakcIvjSALBUo2PEpjQIOYvc+eCM
aXr3xNV4U3ZtolgOhR1HsX6SuWX6+NyhToin8WjoAsmeVAPZUzj3/yBJ6IR+8d/Z
vcwotJexJf+EIt/PadV/Sg474OArZKxfeJ4Fw0QM3/1N+OZY4z7MfAdN6c5rm43Z
dLd5DmSeycPiWz1ea98pUgp+cYkwdBWxIe3Avyw+mzFT8U7e4RKKpSTo/hjja8yZ
Fr/dnA3Al2bH5quUqsSB8ShMdBETI+c75CWWq76Vj+Yid0LL5Fc7evPrYlHblFIH
1rOgX9qWryxmS+6Gc2YMb3V9a9jaeDXcD6kZLSEK8J5m8tevDCbWE7c0itqG3+v1
vRGKCqikhDSlOu+IDzG8+iN+Zz0dJ5uTSPkfLNmzXMCYkMY3fVPYVdgnUMgTD7KJ
UoCLeNZYYYs1LK1zPJgiIoV6ZMlnfoIvGVVwPeMPz4mZFD9Bc3i9L8CugW6h8KIj
ftTCy4TWBB9EIFrsf3fYu24HxyeDA3suomfSi4sBYmPjS/Jynipeynr5HQW1XjY7
KRn1Y2dak47Fkk4kQZGTHplrSBtsCo4WKzzXkPebdtFEew+M8JAawOgE9GxoekB9
D2Sa457tRqzWOjIpbDuIqQE0bQMj7+lbILrikEaihxte9QIPUMIwN50iAM/H86AV
HU52ej3F0IHMXfBkse3zyx/+z4QUCSvkw0H94wMsfdVeDCPiF0Jm3TsIObP7z8ml
OhUBScKhP/EGy1J0Cz6Cb7d35XgZgAD6fwrX4FR2FnbI2DFQf72TM2VSGlo0oF9o
sCiNVeAkRzR+8BnK9xNIJL9LhVFnZdFnvXnVrT7UNvigBHBAJskYCG9o3CloNd6Z
AunRzhSSqn45Kmbp80nStKtyd6WSviuPVqx/kUHrmV50QG1ZNqT/vI3Orf/9jFyB
5PvKr95J8cMdtpgF8E8MkqOxFmgGUsj2L/v+iKScddXf+Iieci+mbB7DaYP40YtB
QWouN1kwNm7K+T+2e5+TmxpK1Nr+K++uUPtoxmhSor4K3PdjGoJX4pf9Z86GwpiA
2MpQkCC51MKO2RfCFWGcriUybUCh3LWafbm2d+CRhUsVuikW4w6+MY6D0UFis18S
sYcvUn2rUtx6WXxJGQFx6qgYPk7296TKL7iMvJ3XJ2c0VsfzUehGfREB8h+pPXC2
n/cFoLzCSHnisDTnJIxn+5skNDGiwSVis0L3bBaPmgckGiwhOhZjtgXzrFD2w9OG
MU4N6uekTw5XewKw/FZwmmhIBbKNZhRi8343tgFPCxJ6FHTLLaJYTxh4bHIN8kvY
6WbG5RmJ+AwXoc+4bki8cg/+ATJgUKVakRxF5D+Is82zDbgld6JvCImFjDaIuq83
iqxuyqSDTa37GBE4ri+nm39nxCNJIVQ+7Q72My/qtvM5KvO6t4w8WrZJs8oL+uWN
uEwmgj5CxIDpGcv7hpcGzVCliBLsDyChG46IefEiQhe0lRIs1KvUU9T/fLDfzRO0
wcbHYUJ/uw74XsfgQGg/3mguajpyH3jnl4k2plIgKgpEe4Bg3DjWsDPSN1Js/ORz
+YX42tkm4R5thhCkIJzEi21TFJW64R80A8v1Hk3KesHZCbMm2sBg5+NlzODsqOC8
Ee1wSjSWvVqT53D8AKa+otwkbainf/oAIygtnlCHXPRJhL+MG7kaceBpysfwddmd
ThFS+CstDdfa+sHKYnl8J7DPidTdvi6est2ZQ6WSM2hJ4P0wgILBo/s4V37948zn
9Ust0dXEXsTjgGvgPxwtqSQJa6jk1FKEbsX25vK35NzahKDgQBtp65qGVz5BTKuC
9rxgisyehV3KVO4V9IA02DhG08Gb9oGlM8GmfFZs0Q8BRyzdckhHUfoabg9S+Nt5
sUs6gJ3fxBFvfsHeptJel38L+YJt/k56kUpzRFJHHho2kdEIR5du88ZmQROnVnn7
M0FOFlGMN2EEXMKcx2bpSr+BiTf5DvnEdZ7s53l5JiPIx7MMjwLH8fLKAhuyYQYl
kP7r+cv5WotXXUPyISm7aPZwi9PbVnogYgv85UyCHCn8nvzu1rKOonrt0tJoA1U9
neyTia0LLqF8R3Tg3AXAYax2Rwq+NhYoamF733L3XaP9o4b7jVGRA1vnDk9lNJMn
hdu5CdvckTuMOciGT5FiM2D1sMLgXCi33vh6DZwHmNjhoKCU/468SgxXM06ggZ28
b3mTXx9SGuarVYMaGSplSvIyk7GxQs0iPaiu6VAWXwR2nSJuVIDl0uw4s6R6GRIP
6pti812iijGJPsbG0PRIEVdhhiF6y7US5U0JPGQUVjLsRnnTfhlW+hNPCB997PJC
b8h60ml1bnmfFTIfyeHTD1iyPfgDEFq0LgurMkwbNDvmAfO1d77TUoIAcIgvthw2
oYbU+03N/Hoa8Vk/geF62bHhDIVWn4D9E7RmketpxjO4QJsF/B4xlyQUz4PsGRSK
49+cYMDCnZx9w3wV8TXi9pFJxRsfxXsduRNkP/VlgYtTljjWAqPvVMeeTFqBnhf5
7Tskqnc/rsMKUInbCLd0BKvzS8kZZ+igvfAvPUvUAvUiCUbPm7C1uwY4kT8FzJh/
FVYiqebuFGIEdk0NUAnTOCkvChtITfv/wcIPRMXUf2NiWPFzYY70SIHnkty4KIBr
3DOFOLyMda7htW5NDiteU2BVjP3spbikZp+d4SMZNGfw3vUDdXZ/S1Q6oQxCCpK4
G5/G96fbwKbVwEkrKnK3MYiwsxKSkAjfLYMkSaUpkR+VRAf4bXCh6632dZLMI3CZ
04CD8M3e59O0CZGmPbFiE8/sS/i1JiLWgW01wiAcvSYXiDwLRzyQQd7PCDGdpWLw
zmv573X7viDs0JktF44KpgtfDn0gIrp91BQwNNs2WP7qB5LR8WF8Qk8Z9WylVypD
q9S1aQdjMka1qRJtT8rAdSIHKpTvk4/sfGjeq+xETdEAvUvx0QkbfB+uVy3AG3GK
E3KDJmLhQcw75rPrthFrIFYHmoo2CH6SN++wn507Fc7vANL61qqkYrJ0q4Z1OLoj
SJaS3oZdTuOnGzwTr83PEm9ZEqLgMl2Uq99WAeNe5+T8IPB8hEK3q8GJfpnGqeFN
0gIhpeYMZhd6DmdGJLrdoYyzO2GeFzGHS3l4T4juerJRhLMcpr8EgVir3byQGHGG
UUqTCfMkDTbZ2NPD6wb7hpUA2zEV+t722F7gWVbgirNfPkvYDxHJFzNdkigkg2SK
9vuxtTCxlnTbl66wzxGyfDhUBE63BTKyISf1/HJAwgw5OSmRduY+6uksf6BEV0eI
TzRwMB18KHNTjuOwr+BcRjxwiVxy7Bd3Ye6Vw8aCU9NAOAyyr2HD37jDsHsHWj0s
YTkt9PoFAMlB3zJUM+ZHXyFCi2tuHKWu0n6qssmHrAqjTkjsZ+P6wm5x5t+BgN9H
8CDtizCRlGAnG1Hr40xgZRMaGqsAzMk9crVLsnuOD5jbflwuzk1d1Mnvx64cjRiF
m+hz9LoK4bYHgH1sTEeK4DbycxmG0v6UkvOQNUUkaOQSRlkBzSSaiYgob8A4mpMr
7NS+gQYwnWg3O6+1xDtvEkBCzdMCUGlVwqdxr1xYB2SZPmmio2pdal9ByWN3lvN3
8p7XgclGAD6jX0mPwj3bqjFNlxK13568dULLdekGH8x//FNPd3mjvk5Nb6Ka4XAW
ghW76m75eMwMLRxulL3Z15clP6VQeUuPvfKOKmv7E4mcaojO3XMTFb1CzIlM5mQc
ZaiJNHd4/3jrOxJBQtPuVQ6Rj3TW1n5zqS5o97DNnj6xWuQlZFd30Fw4CtQ3keoS
bNRsAlnRhXBWF0NngV5Guy6Si+5RdkzRVRnZZxUK/WMGEy1i5F0rKgXZXlIUyEyd
uuJPnabhYiB5V3mTj/CKw+cnHg+SONLiBkIskd2MIyn2GjVxZx800f4hgVdy/Vfs
KbfsA5GfwLCJXlWINpWM7erilWUz49k57Ix470m5c4OgEqCnMRiHMSglXGhOTmTv
Magoi8V+jpMPN384k164aotAztwk3JrhkxO3QSa6G0/DYxJrJokl1RhUTd46YgbI
OtaS7OPl5Wn2LNOjNgCWTfXtGSnsZim2rw9we4Trr7oC6YEtCvzzyTCKDeqViVJN
tr2tYxfT7WBc8vtumTUFediSS/pHc9FxQzYojMQ3h8s2tCLkmC0WaX92Au5a7/xR
bu5LjpYjm6uij+KvV6eX+QaW2H5pSaebmWiZ9QaC+F2jeNvxH0Ge7pZfV0qFm4m8
rnIoHu0hVhld6lAFFkPovRYZ5vEf3CDUBARTZ/A4/3YOs0R5zfv9+y9KEIbdY3kG
tNhomVLjogCXvCTfNIPQEiF1+x//Ksd6WcGb+Y+BLRMM+p+gegGb9sVBrnTRKuOc
ML0FA7uw/tIcdCoECAaeEQ/QTfEwczYSjk7odTFTejcb8wnMRaMDl6NypNyVRM4w
q74O2xH/YtPSo1ei4anktPWA14Q+ldc68n5qQaQYXaUuKY9wD9ZUftExdwqQuSfq
B/mmx7A2K3MHxeCbarwXw9szQOFcSiziJd7tkmdSqua7zUHxsH86m5mOIh3I3BpZ
BR3MoO01+vVSzofOIIDcJzKsg+es39tISDm5gvGONR8eLwfgF/eTB2YbRgRbiEoG
QX+iUKqhJfndyDEETBht7m6T35UslE54CJ+YKGTEk5r/xCW4Hsh5JKd6xAWxdJou
Ml0wDy1ts2w5B0JJCy2rjqSiOqxBOL/1F5cO3KIz6+TxuJY0d0dDGLF/zSaAVaLM
ADedIyqsQXNFSpZPrKygIqEGGKBfO8obBOLJXPL8zsKrpF8YSgSFZqaJuTQRXq/P
3wQDNvvAyaQJGB1DBisPo2TN2Doet0lmtxEqaixuuAzrfnVNPZwCDKb3s09IMb/H
7xGhJ/Zdr4Ix3/72P4Kz0FVm4kH1W12Q0SkORUERo/DdaQpzpySSmKTIOB8Mx4Bl
ZXzezgvAozrqqua9O1RlQiFZMVKLDgx0xRwjAMCDgMQWrbLXdppbQOJlPd3b6b4Y
grsMzw29YtRtaVjBmfKKVWBwy8xoDWFrYPBGh1i/dIKCKCYeWrIeOmjSI830Ye2S
gkHs6ecirg8klUTZ8Feq/C1D08t1s0tZR2YZsX6vISdT6cF9dYBsMOr023C0I8HO
04iU7ESmPWijM8AMheCaD8YZIy8kOZ0zmr2xa7TYrnWR0ro8uCyew9Vo1Q6pGJek
b7uhwGoBOzol+1exBApeIazbVyuBijvp0qEFLp1L7L05gsGqhp4Wjc6EYQlD3Xog
bu3/zqbOYd77O3ABCTh2Cd9ac4ef/d3E2TM2i18ZM+TEEZhqUkoKdT+gN+vydg7N
+ujAxq9AoB4OejjMH3Fxu18LtRfqm/5Pg6rl2oXh9rFJENgLhz+HUChsaeg3qZeI
OJWfX+VOaRoK09zE5J4QJy5FEz1IThaolDdBRDur8MdT0udHIuHrJ5rDM4zFdVR6
nDmXiBiseN/fygzk6qnsF/453A96nQJ0bqODLK4Dp4D3/7WHHDZ853AaTW/yRAGE
/eaU1JI2aRnuvJ6NYx3JNWFO3rpKLumbN0OllusmB51bFbEKx5tFwPrclNBa4ZE9
bnI85oFXpv/WafCjV3+p4lpIVQe1T8t40eQ/NbyLwIs9ym19HtTaRijE98XK4lIz
OnksMeUGN13RawYm1UASoBLyWmW3CKRMMOFQLpMkGwlYGgIpI17lTJXEnK1iphmg
H3CTKknBjZsJEkHLIm42hzM7+gFowClW/G279SBGT7MeoBEImuytAM22MKVaoY1v
/Iq+227cozKQzhOmrp2nFCGo/j7519/S15O82S9aSSRPqlzqF37yHbsW+UqfvPGU
fxwZpLmia3wVUpCgPyIkHaZvQkG1H51dPIWCPI2ZF2+bU2w4rMRQIykxg5+zyIpm
Re3R9e4alQn61G1sLxnaN7ivY9uDEc+lv9lAl0vEk+KcMxGggpKDLflXqTlSeu+R
HDqnhRTHupsdDzq1HmI9EWZzBtMga/rWcDrKTfhsX87lb7EN2avttJ5++2zZMpBQ
Znd7cMnpdtlCxmYlTaRMvNQnyBS+BTcvoXzQQLoFbO6C2gOrYIgzKAXR+4rso9tE
57IdJI75J4k1oMGP8WL/7mEPnumB/HzUc43DGYfDApzFa1R4Cd+Ox12PpeLszCq/
jyJTrq7FfLcrfJ/b2/Z5nsDQ+TqB9GE/afHFnJWxSpQYuSD9rUvFZzInyLSW+SIY
Z0nhaZT1vKVHRAhJrYhgP0xI4p1U80t0Zzd5vgbgR/TT7t/EKzhQdEVbhNE6r5z7
RCFY5I4o5lturQ59qHMDX2NGmOI2nYqWRt+y1wE0Qo/8CtIOFAXGaoNVJDKfoXDK
1SDgoO7exeYqExjzPFIa3mRYalu2cAFboVlOMNj6FzqEo0/R+2robnVH3vD/icBS
+y61t96LFvThVcViN9W6rcf+blet4jk82/sk2ruH/EyFanTUIreFzHE538cQ/8Wu
C3ul590gk8XB4hNo0aFGGx8gQUarWvhB66A85kKUvgErR9XzGMt39ddfg6U3kfQz
xUwX95zYPTAHct+bqNWsI5Oad2URS8ZMCB5S5HOmU1AGgEbgKfIXN8d8YxOkJ4/H
S6+Xdhy0kq3bHrWSX1LIVfSG8+uK6ZXyZm2fMtugm5XGhkUfIC0njjW7bKHS23EF
83Tdm1xsrOo1sJNuvCKFcOs5K2YzmyRfBlHd/5qDg7RYpBYSIbt34hLwAaaf2t3W
w9T+NAjEzHjKH+kgHD5Z3tDVdvOXV6PJ7JepI/A4dzG1z/QvHMvzOmSF/OQnLmRi
kvZg9gYHrTc4yBQsvplqp6p+HYwrKKwrd1DpC6IDGGTBM2xJvG0HeGAe7rKd6TQa
hauYf4C/jdPEFnLsIxdjWbKGShTVCu7BA/hvSm517uVwcpNdFjenpeY0gYuSEaWN
iPGabdWBZIGC/HeS3Xckny4uVMf8VYRenoAU81v8jd7GCCNw26r5xR5Tkh5ibYE3
P3B0EtZuWyjF3h+273WScW5l+/AoiQwQIU1UxSnkQSK0WvpQtFlRSax2E0sOJTYv
Z6xCZ777l1LwJT81DLItAId0VrVm8NUmmg5zIcWO5vJLvdnPqChEJLqCJ3vK4/md
aO8kFPsB1kc3ONWJwt+9LoYveLFcnEq0eF21ZUEsrD5B3F6EXVUh9cWRhi/BTze1
PFq7PYRUPwlEBTmmafB1KsGK807j6L33acb9NRMICUALAm2tz58mjhR4FSrnv7Q1
MEtL6g3TBFR7hN+R+kzvnyjAi51Uu/s4DZsMit7vUUaKASqtAeuISU01KYxLVLVa
/+NK/OKRktesjZpBKuKuBPgTlV0sHw2Yo1wtIr/6HqgypEMQJL+8l7G9ssYKLLQ+
LV+2wMWzH9uJf4PrXu4/pvSAgj+H4eWHasDMK/xV1kDe6aQ35o8Rv69EXYvSFfxf
zRhQVXmhV5fkCAye2VfypKBiWZm912dP8cFoWVYVBWbqpooUqpmpC8lgAI7AljsE
OkGJw7vbRKcyMYHBrLJpfIygt6vTSdBYVdewwS5Ca29F8aS+XKpgPH1iMn3Njbfb
Dqgh81SmUKraDkI/f/m/kmfy9x2uZ2rWwTwbAmMZndJZ0JqVKV1Pn61ilr9rk6FY
fpB89vWic/lDYLEAve6kpwPi397eAo4bVpdZ8MSXD9BMngkz6W53pwjqd8G6uYBr
ki5mMY1EOlokGMchJG2k2eZLZVOnYcpCkXX+MkC9ijPwzF6eMmznl1B9t76LOBHp
sPPZ0bHcheO2DjVac11XB1N++ZFCQ5a0cWygfsertAZTZ8edQNWxWzJDL32Z/F14
5zPKHYul1rSZkkAWqq2YDsEk1T6sCeNZSLshiQKLx1N9c/iIruO+vn91gUQr2HL2
LpPMqcL5AVbz8GLJ3q5fB9NA59gzgMlIr56tsdJ5EhMp9Z/H9kSl165VZLBI9QQ8
cG2X9as+s0qY6IQ6r2IN3zbMD9OeIY2iJkn8I5SYFbWDIzhuf9/ZlJMC/UWWXQjt
Lqfl+J1xeb5g7HS1YskjmKpIaKHtaKadApHD1stAOR5z0uTqfd5e4CvLl3ot1vgS
xU8Sn69HZYsJOplSGsB9qMjck4tPpOMuRcrDGX86GR4f+RrhizrxD06/CFUEx8Vo
p0bKHT+6r0TEpCIFtv8uUBTxWgq2PIj9+1xQsh6SJQlWb7wojg5REGS00OI/papu
oTNYx5AIe36p75IfbqjUiO+KUtvlzmT/DMp517TVAxsh6kxlGhSlXdZ0NNER9o6+
+0HVjkStyT6q7HmBpiZ5a/ZmU3qNcliSoeiCrLokWSZ4RskqDfow4BqT1bpbcjQY
GM/uscgbt7K2eZAWPvnCq6OnPuz1dQoOWjwiUrwyOKJ6+CvfIxG0sYHfyGvcMHVj
tCxP5HXvLmbDdtQ5++Jp5y7fGtNQGDhW2RAgTnPGfj0AQkNDLncgXmiJI92bZDQN
9QB9Fi49gBoCZVOyRXfMi1Rkc0WUUlOf1T8FY9k4hgKkCzbMWKAZFMwaLxZ+t6FY
YbGtlpOTsLA//T9B+qBdZoHYEqQ6dwWv1VOlm+w9v/a4DASoxQC4UPNW1FTJmC0e
WNrplo4PBoPnPjT/1ThuVFt3t12M0Hi3u7U0GmwX6QQ8WAmKCc98AlFA59hGSvYN
7T+5sx9vgEvQ18nuGw1apN40q5VoNf3GCs8hiZpmYpmXOIYYLLRxS5IkOC3z1NkY
of4INR7i9SsQz3uXWVaRYSx5r8fXhswCLaIdjhdhiXQ1/jG+PbKn8clfCTsMc/ov
m/OcwbJcp0/VyF4qY2cjqJUD1KyhcGRjRYqsydBGBope5Ckl6Zpb7nK6ZrNLP43M
wZdF9n1BjTE8sVeq/f6jAJVrStRPE5k6MkAN98aed24iZguWq6z+7WWG2P59PUIZ
5cMu/P7Fzt9ZITX8KqNEZBItkKGQnnP8H/NqebnJHBO5NfRrnL6eikm6kduJEYGB
+pQq4R5ueRyvvve7zS7T3kFuW5HJ5Au2lHf+uflnMAay4D9HuZDp4VLSuzhSAOvq
clx1JluzJlICitpwGBI4VNHI5Bp3WcAjeRcxhRQS4rPLd1jDeOHIj5c8HZaDkghb
+Fz0SV4cCiC4al3euoY+JVpVjVlP222xEj7dvoDnqIv3YTrmSXRDQW9tmQD7nlmu
uMI9ukqKRF79KfFwWyggEDLUmkI+aeVr0Rv2jtjNl+h0qe+JvCZsGQzXBudLcKMG
a5Pvvsj0UAr5NT0iMSNwbT6MOkPNd5aA8VUveSnDfHH4SkxpT7m0TBNlq4awDBij
/aJ8Oba/zv7GxN6jAZCYfL77dHKUS3d+a7R1+Q9BvWvly31U/xYnfzLzZIYDlm6t
CnyhYH/aPQD4aLsWcWIZbPaNm837M/ZKVnOy/0znUXFww/y1w4a7gNTn6xmmG5GM
2+bYhpwjlOtJosbyYwbFZEuu/+xXAALlK7p/4RVTB01VLUiN+7ieVyMLzu6gIaP7
8MEqUGZIphfNS+wSKlw6K9beRY9ZIzwtcnROeW04WzczK5L1NYCGg2337rOCL26L
EvZveALe4sv14Bccx4ghXReboamnOSqYvQ/Ii8Q3+MXwXb7ytaemle3IXQoLnI7z
bt/k2a5tediDCAyY5j6o/aDJnqXLrZJrEDqG1ab1f8+ptbYmQ6BGK4qXcv8M5nyG
BsTgGDBg+S224krhPqEBfdqtK2+h4bcaqS0PNn+pAFzjFbIYg5wxtAY8fI5AVhPz
rDaY4UF154wmlYUf4oAyRqFYTgqTavZCzTfZrmN3x091fiQrAfAL5UsZrIsf15aE
oKyc1Psg9TeSGOhlTZB+dSxWPQYhkvc38MraCkMmn2AKGQ5q9Fl5YqIG/OzkACsn
cDP/XKHkyMCVSqxSzYjCuJ4zKsOItjP0/6Lk6n04VvfFG72+0xGARtizeDTn2K1R
PM53ufD4TrZ4QL1KUapVDqwyo7BZLQ+Llv6y2b9gfvdKCQEjo3gwCR9+mb0Bur/4
Pvy6C2rmMj9+qySolqXgxIbAw6OF1j3qLV5Xak/NmoOKI6Ug5cp7Eji4oOT6VgP8
8ey01yNMkh6PD0BTd4m+O7IpgaVnP+3E/RSmynjOfwh4n6wP+lbc/72GM3zjGSPD
faXRu0GRupNoiUm4s4rPHLrte1VZiKCijfJp++MXQbT4v3/Dg2DWACnXxZhxDcy/
pVTKKjYbeL+3zcs7zS+Rvj3m3yGdw+G13euvINh8LYx/hoVdmbAe5U7vqEPLXCWS
dhlL8A3DhxkLcM+E02VpefBKHYt4EqaEk7baqI9D+V3p3aZtF8MTbg7BUJwgDftg
oZ1wJdtY+CnJqJ+Yy5nD5hthAmKD5XEEVTH6xSAj5iyP+odRb5lYF3F21swEftOc
Btorm6GNkeCCpL45vMQs2whI65s9t1bhG/+loUdU3w5DuaJFk9z2cp7915K8Tumw
/vEJdRzqr02ivydP9XdxxAEekHYiAEUan3GK/NMJA4eL0v/ndZnRbq04D1OJkGcP
o7vtxAWK+IEPO/8ZsXxkDZMXPN3domOd37rhNS3Y/S6wI5/g5+H3oDIxwQ3PJu4O
5lfM4gkHaQ3s9x87l2sqKN1mK+rVyb/atcY56P0mwqhcmZYoSaOQsw7OShiXO8gz
7EtWnlprgIk67rPRn5J4+qq118FTSeztu4VTpN6IwBU1R7QeU/exgtEdp7/Rb6U4
NpqmvKFBLK31GCZPlz0MzzDx7Ji29sY7G+3EdHPLVXhpim/Gc/JclL+HOAuxd+vu
jH6zILw6OmwAb2Wl/e8/rx8cjsIJ0KBTIBbaEUHpOo8PUBf+yoVhYk7BJ/xYMWEM
csw/wpE/PlPqKIFNe7Hj/mBbnEN5A4dY/q+la8sDM9PMaHIFbVhAcPU3AfC+yZ4+
PhseeRLNufh3AnBce4K9lZDyk5tq76X5Awl0vBIKs3fyrqVbazF3/Wdjtx7IV80f
z9AF64qW5N9DWJFeglm3KSu2oDgdvjdStfBjq0HGv/4IBCmV6OljkzOT2aP0Mtcp
3YArqi+6BrdoDD9Em0tsXD7501d0titVts70Cxmh1gMrl4X4mdrNj0iWbiU06/E8
/hA/xzRmzgp7+iUSUSzzMDFkqZGAqQz4XfXk2vX3/teiuDvGok03mmKYZ9uzddG2
dBNRaUV7yUS8Zn7O/OapPDDiEmTR/B2aTYZJJbbRBIqUWuuUWBdiCO57+LYYQTZ7
pxEb572VDZ8m1SMFKLHT/NWwsAQtE/47JzS1krZXA5d0VIUekuibAfxDidcadZg2
67Vh8ohS5kJq6QZ+oioFUxw/jQAIrUfc4U5KIKYi8WixnAo91hC+PMrnrfFJyuLp
ZVCSB9oM14DFBwNsR2i4rTmbZj0fgb5FQVEV3JODOYzL3ZtWR17cDlwBcHqge17t
ckPNcnr/h4CyDYfkJIeaXup4qOQruDC0R7CNcGU3cIc8pl7DZ+3/f2+tatIh4q5n
PzZK4HoXycdXpyoWadwc/PYFfT9ciAaLYb3p4/Cu1KrVIjwbquHl5FCzuPmGEayb
b8414z8GTBaYr6mK/tPNavXwkqossELAq4mwmSrqk3wZ/++xGu65d7mHnhCg5Cjp
++KN03WizWmYq4fqWO5dpl4j6BIRSQmNEwwduzyQcyYS3oRTsJrEZlefMsN877Ek
NMzmpPaDAqPEoZYlSbtZNXO+u/kqufVjGOBb1+cOFxMQ3RYkXSm7mtkChmfLleUP
pyI1fMkjd58gDszbR9JPqw78PBfXwZORTbdsQ/DNhsoacgJ/T6p/e9TJ4TLDQzRm
oH39gsyeHg0GyOVtgdbeNVT3hIGBxTE90kiHRrNcd9uVrxhZWQ0ui4UfI5ZlFWdt
OBnpq1ZgGyIWOu26w96tFKIZ4TMboC6xI9Lus5hfEZgB2wAdGMAOAb4rOKCO7rY6
ftBjvkyo41K2shWWrR0YzkEsYvo1I9U7p4EaViZ4OHwatquyL9X7UtZqBqwKySvz
6r5D6kbFmVOTNU7QqfANqKPslcSfABgxmF+wR9bNJyb47nPkwB9N63YF7dBpJvK1
ttjIdmYAN6UXENAejN6joz7jC1Tt6zXlEevIXAlB4YOYO0Abp1KiRtd7dVw3SXdi
ZkJ0hKK29kHPiMlrPN1GXf8KF911e7/1ZhPZku749KQEQ00o5q47W1akphmuyIcn
wNVFRdBoZ+jCPxqRc8ub3IVlyi8gsNSPpoxAzLUh/10tkB3CV+D3aBpg0uMDx9Fa
RXezhkGTqL0P5n/6Ay1MJ5lgXaNT+7ww7dfLkk4GoOeIMYIha4LKxZumwmGTEIMt
jlRRBHRosxFZTGKE/xmEE+g7OPCisInUCTzR6qxm5mNKbX12TQaIMlYLS7AePYjD
GoYsk/ISSYn8GgEGNRhUoqS8AdmGGMbU+lE5GWskbs1FSge+nrHWGH7C46ESdfVq
oJiAhrdibgZBSHWBo8bMpcX+KXc/kFV3Tt3tu659fzMLK+BxB6golsgVqdgzG2cu
00isH0WR6yNCh01EPLTZ23COm5mYp6Dm/mlLqxeNVZRpD9gqH/t9j5AYy62Ecmjq
wFODnrPKkLc05OaN8BrqziblO/wvFbPOyxK5qalEWiLjRoX/tyY6VaJC0QNueNcd
z2rzCc9ZhdjcnPGqIEuC2JNqEkRP4jlle7ekpXny6avSc0Dh1aZte5IkQlzh+3Qr
3QYkZBw57FdXgh3aoveuD5Xroxpr9y2jiFlNtr3idAx8Fba4JV/smbguA4Ogmmjs
ttPcHMsvLB0ETahOR5WgMYcjZKqSjCM3YDapTRcyoS49bYWOqH5oQMKHCMvtcalu
TtykwfsTisOFo97/5OHur+lo1ueGXtZ14ShcYT48Nhb83/AFdM0oZXlfFHGWXGM9
3h+9i7DEx8tF6yXsn5bGsE/BKY6DftSJvMzZJxgoLLZt/1cpX5WjUSsetRBUndCQ
Haigmx1eSWhytSiMecBZ6q8+vbb64+k0nbggndMX8GC4DLv0nxFrAZOwvq2SnJT1
mDFhZPwIL18kyfPn5XwTpXAiurys/hcnIylXLlL2nJh1Pkh9soFdb+t2NLW4PNTd
oknaHXMcX1L/WhQHq1VZe2ty5YlYriwnmbAURFd5Yld+Oek8IEvOUSqsHEG0HPi5
MxwxpQ7V+ahMrl1G0gK+eBv2hYFTBQNX+RVEAHnm5rqG18/FlZyCSYoFJBlVVB4p
P9VtnsfdTHzBQ6ZCY6b3ZRSMkKJnZQzQDcl9TL4s8INa5rusibbOz7hmqCk7D7GC
Vunob2XnyaL2NAherp06cX1i042+q7YJKG/wgLtVcxg0aEvlo/L9L2jm2pyesS6l
9IK4cOKyfap+f3jmckjgy7SfRe853IpvNCAeIT+V9vMTG7rtVMgShGvOx09o+SZ5
Y2qGS5/yHlaGk/CrN2P++Yo8U0gsBLVC6p1858kMBo2O5Wc8fDhyA6J4GJ19aH2T
vPi/IiYJyhHfLocqgkf9NGUUFdV7KURgC0kktC4z+ExMUMYp7IPoa3XMSoVIfjxM
yNYJXVwsgCGmqpjULBNjR7oTMhj7BlkOTTSl2gCLDg5MPSTuyU91oH9HPKYha7dx
+I4GoD1z/qGhHakXEuxZjWo81hpefypF2yzF+31qJg4Fgy66qD/PBMwCtuNPchie
spJo5BGTI55dS1tX3y2HHMjqTjNYpPs37OkphpdPlSjdiES4CL8mVisUvy7yCJtV
U3zjPd58uRhD/3CN4Xcklagr3GhBLAYf4EbBuRc/SewVOk+1NFIxCYXqvAJ3DyRJ
ab5IkI9w6TP4EjHDa8sl2DBU/toBKajzKOdP4o9Gcz5fTpHD4cefyCu9zR24j8S9
rvuD47jWnNSX4Goz6kwGz+KtwExGl3nI1HSHHBeY1Fif0us50ONZwUvxKP9ZZhZD
fB/LqJrmixwfHDFj/+bXslFAU7uiQAC7gmDse0QnSCAExlhjWsG5NA6q38E3r4pM
TBzquEQcQKVCDUQnhlLm/eQ97UsivCv/43sudLirkkdtSc4GPSBEcn4kpknuP/jG
f0kOVTIXnp41ooSrH7i6b9lUfj0yXfYHhWBXE0wo9xZ6tAInhE9zybw0/VNyFFqv
AjAWNSddNCniSlrqOSatjzRUkvphMtgrzdf0G4z4FxfsrEx6qPFGqbJzaahwK5mn
bpos/8YASqIteRute0hhYMIEGr5zr9RrwaCCA6P7tVFwcx6klda5nT5+E+Ch5gty
TAdF1fRw7/r7fBSEQfdOrpV+NP1VKrruLZ7bu76MYbuS82TcIu1ZnDOscphptDaV
3z6+FQCPhyI7G2pMuf9A+Lm6/TPdgeGUrCAIGV9+U1oy94gdtgt+2su3p9OmKQWR
jAJYLu4mHds7he2VN69/PzyqAaFl8h61wKzWLMEWRbmdfGyPE1niu7erPT2+w/cB
E/TEUe71GrH5GXCvpakJoO4zVcZTjqgJ8MwlaxiI7YfrDYk0SeQklpVgm4CAt0lr
dhs2VHfuBsKJmkBf/TvO9YijBeAFswzFvgS47Q5dW2kxjsaagWnILrQwRQ0u6nnL
hWXf4KychKyAtHutXW/36ax5Iw/ARVF/3vEvRbmQ37ZzrZo7j2Yw7jXeJjiS4M/u
mz81KvwASckz70idU+KHFtsoRCELOTS8n1bBXaltnMxb9ItUJxwgEf5VBspzSQgL
eIq0RSGQ2SkfzENk5wcl6VGjs1U2HhIoR6Avo6s2pA0rd4V+kqZUhU9Z0eHM+TGJ
dLgUjOkatDNnIXw82Kglywx3yV3GM40IRclsqDW3jqBQ+Iww6JwzDgbEmwXz8dxI
swqKIGsI5w+TLB3H5UXHybxj76TnjIb1lhwcOWY2B6cJ5RRx1avbuflbth/tkbAs
AwnXY1PRmkchCC+hqQwmZ10FckdUBBOayBgBSkXjx4kHeSdgrI1S/u5U1m74z/30
2mmUvtuD35qPtkPkGeF6g10kTivngfB+nmw4Xc0Q17Mj8o2I4rm9ygaZZJbvkl4D
Tpmz0AC8ykIrL1xZ422LxNq5MMknK60+1N23DiJ3JdcHY29LwgwakuF6O/W6mZ4m
HZbyS8vxOS0l8oJWIXZZ2NpTGSX/77/++c72m9FWJIU+FXDnEXOxOlmIceMcwyzk
R7WTRZtbrVflhvplAzVwyah7eK12eklJ1IOiR0vr5K11kciLy5+Ysf/G2oWZK+R4
vhf4WOTBeT0MciABfsiteWYGT/sAAIN/weDa73Uf2QLFq/+ipT9mXNX6FTYFWmM0
O/1WcM3UJqVVft9SAKPxL4DfdyM4kkpTv2vYGRr/VgibHkrZIyZ3KHwjX5DZzMMV
mNPtaIyXLk2lRmmRusg54XNGEOwlYImBNPMrSE5D7ceg125PbsxAR2tKOx4XRgag
Iq49PPM6CD7koth+xQ7JicLr62tZ0hauaBDJ05ri2cDdGZBcQhp5Mx54zyjF76md
BN92xFaIlLrUifjCUG4ZFyHQn/SjLnHkmIFt/PuTYEVuTNJtb75mnI8HIdAtVYYo
Ta2jhIU9jCg/AL1aK7AnVySXI9g4PiOK4b6gxawoiYDUT8QKK5etoDQdTespiyg5
MExPQ4PImddDG8gqQoI2f336Zw8grFgcQVHtpEhCC/gyjHN+4EcTn/vrGofU5LhI
tyuVINBxoM0fyLhec/+FE9yh/wkvC322pudVUKnpBmmM5dFQr9t/z/tx0Pze0pUp
Rugl3Ipvn+97aoqaiJuY8HjJUHOAsFY/TjGlEh2RbTgBejniXOrkbF91G7bPz9+f
4oAlkCY/WX/jGXrWEsMfrOpThI2LAJozzB3t3s3ohyUEPRGHDSnbslqKJV5WTANY
EToZaeJCO0UMIOGhVzhB0gqjW9pnRnQxi5jfucF/OaMBpSKmiImLhY0Gb1cVb2kU
u/fvaN35cJZceg1kz3/pYBQJW5Gw6aGRR2oK79NwYn0pogjH/8xH/aAqV4hcXRRU
hDdq7hUVkGJaSEDZ4Y7N6rkEw/l+U6mlHj2FjT6Tn7hFt7rdrpqCks6VHTos21QQ
ZFyPed5338YnTKQucp4eaYMIjJU67K9qiVrJ0EAUfCArHWtLDrJX/8BrS4yFrXtv
VyLxYCJZ3/W75e2IveYlaiTQym8pqpDxD3QUROptuRMZwBa/ebAxYGgFIbqMs1cd
wOdDZsugntpTxx1yJ+mQtXQ6dMJIBlFgbD4dvPp5wFpWwxRNxH00w1vNS7bvQQSI
U2PvkqXC07e6Age7OQ5LhTqyIYE1T6Yf25mWCV0zy6Zf+DJeYNvgXWI93LWS4kpF
0HsjIF4R5M/9apdB7bakHMJ75KcmbABFY6X/dtNBKhfcwamh4QQIbnl4TdeabXAI
Qop3JmC96vUnPQt9/1n9/5xfZG5ShvhfcLySHFJMsNXPtR2XYIOTlzC1efCA2vUb
asZY2WJFYSn1AfGL0RyELedT7x58hH1fLBdWfO4pm1VFPGhV2iCEPvveMTuJhXS4
T1t6GiO/9KAhYXYn0oznWypk3XleymX8wF8SNPOt378GsTs61ghYGiF/wrIeEx2k
mUVIDat2RlXN4tRZzdlMgcL6UTNsT45UkBO9WglQWDW1aK7+0FdLt/7YQzYuSV2g
f9WID2jX+IPOYeGwYuhfzYzH+8Yq7z5Iyhxo5LZdSO9wPZecWkcdJFWqZRU1CJMH
rJoQrYXvpv+zRnyBFdiZTmzs18fLJ4lWDMPe23UAoSzQlnYUY8BdXT4f62ZoL8Sg
1h8SgzJB4DPO27+vpnq66bsC3T6olB41qUmL3TYvs0NUvUdA361QHI+4S2umMbt/
Gbu/NzxxPDnpYHJPeBKllimg9elsVZMQIUyaRQKDPUxO4v1VRodkvc9cWIO1hYrB
ZiUxSzlyV/jdIvvbX8wBYLTF+0a5ITYFm58e5opIep2iiry+OnDeAcK+D1OuCSYG
YgPkQJGMN8DCeyq9ZkHvlcHHcY6+QFDyCVeeMOE4PXomJzKpP/0uDmk2ojb0fJBg
CKIABYOvBHFzFYdqSsBmZi6t0P4HibYZzaCWrkV2evjHr/6sVKJuaZTwUDjdr89z
6q9jeKn9ixqGWbCLWTM0yM/9prnnx/cNkevRCcbuWprWcYDF8MeeWoh1oZRoHWCd
UNU5HZF1Grrq7kKzN0IgCfqn9KKj3m2G0ATJ4WKnKEFEcARo1eSsj9tmvycpO0X9
pOURy5Ju/ggzXEKouZWt+XYc7nhrONuwk5An1iz8EDDNngWPpwcDdSy2opJb+Atd
XoZwZkXn3NS4w//8AxBa2vLAa44DzVZCh0KgoIIw3y/W8YJxFaFpurQThxOnuWYU
VjGaiAB3X8qiG4AEY9mAuvbFagJRoF8vjxhpYooJnMMlaBi8ciMvkYd8axyWzneE
+b3/RxmsGV4mMXLaji1otE2Fpt1S/gJk6ptjNy7FDKI3dbToWqbYlhI8mcJTC1ju
i0oyNHHOOhH2C7sW7Hsh8UpkAXi97Sk0DiA/BYW8ibSBG4G41sUXV12K7a6jxRMi
lO3UiRNF07mkignNH5oFHpPuediFgoGjm07Ov1WiwhfEofO7qCKIjxilRbubNHwW
zdSe85NzBjHt8RMi3GKaLgZByU7FQ4Yugm8lOChBMkZR6Fx4URVNi7IKt51Mn+PD
WMbkjpZihP7yVEE7fhWFox4iffHzJGMRHcHoJHw05/O6WGtbWR5CYiPLFESZqPcL
v+vvWYiF357o2o9IJqZj9fU5kpsTRhO305mCzjghkOF1TDId6d2bi13AjKRRJ7Ua
JiE3E0FxkJmdFJDuQTqv73Q3C+xw70xOIwFOscACMuug7dovOeB1KXMluU1OwhPx
KlsxcZjdcX5Mv55S3I8E92B2qFV7zI8sTnWaBCpTBqGtKiXzqJMbqLJ7aPUs/Oot
iK6motgu1XdiP8H1pt4p+pUjAIdKk76IkCeCAwuK8sqqv5OjR3u4m0mV9g/byDc1
icL4PG8WJYEzU6pOFzFFIhmiScFWJpIAr/nhz7AO9B1mvNMsT11KD3osX0joNVDz
OLkNUsG4FEcQnnwfUlUSqU6H+W0V3GHBDMD5xAf9S4i8igKIQGRyrnCw4bFAlzxw
8nOLMgccE8nbL1DuO8ZQU4CgjGw16awwZYmNQw/mlXhvCORWQqbVN7xWZKaTRSMk
Uspw7Jq9Iy5F46QtveI/4p2W/+zSB97inIUqxeXKFJqvwDEY0ZLvqTzYwbOLpRJD
I/onKq55b0HW2+rpOLa3UzD6mSnLFD9to05UqiCv//SK2NTWZZGYMxosD6bzspWb
G/avlC4HBvvajS53D25tp3KNGTN/X1wdhf5iKSoXtl9oI1K94ZmqkIQ1FxfruOPj
/ZLBcbMYMB6G8hThxqV3Xk1bhGMt4G/IDlg8F3gkwpkx/NE0MPtilhttByGuNxeM
epEU80tDlYpf3YEn8+NH1P1H+1M9Y68SRSpOfw454VGV1GqXt4bITFJdF1G3Lfuf
5O+0t1+bIe1j6xz6uM7OMHxK9mL2aZ6/LHzuvjJiLS+uOBBjttJrAQWYbR4IC4QH
r1Lu+1U/v6m546GGB8VLhaLpZ3KUfI7mX+i4F2eyET0m4G3B/UYJ6ArNwn24uc5y
JfTx1AQzbIiJYzehfRAPCArHUVOWcVwWczoh4L8yRjsK1GNhZ6tE6Rn8Gab+KJ69
PSWDPrhWe8pCNQOglhyBqMjBIMRL8RPKqwUH/LYlKg8iKvfBAU2Of36VSKxJ2n5M
O0ftNvt4PPD4h5hhgbvBhbHl+SNw5yQnWxv+C1ZYb50fFcWuwvmQY75NGZQOu1ei
FfHuw2m9YZFjQHEP0R8CJ8wZjko2u/fFUkBn3bUI3U1zjpZ4v5++Jr/rHpl/7G+b
buNL6O3gQg7Z1lJHUzQ8uOwt5E09ATij7av15lbb/K1sQz++dPSeFBrXmGtha0Kd
xMmpc3jAbfgymVKOVggPjwjnwLX9UqO0kAKZRSDQxWRwsl51iFbL+cNsnstZVxv4
hC+//g3fcnpBv5T3Vd8tPd4H1VhzBhKIaYzVziw3Vyv8uJzdGwvNuTVCp8tK/DC9
ORv5ykVB5jcIl/lFf//ivFFtETsn+H3c77SOjBicKyjE9BVccRcKZZ4eB9vb1sXp
tsPAPjtlrM5ClwAXUcNK1jD9hWDGMv/8I1upTQ9esS52UkJPIllGxoyuHYWUkiGZ
ylYj6Ul6OjXv7YOtud32a/ASaJe/MfLYMc40xkZ6xhkm2XCysCtdQNKnMCV5OEFa
hf0DXBj3dIaJj2hPkYPR8J3ah+gvGRqn7DWC/eDmpeaiTqmdhyrZ1ThcIgTTIwq9
EBGStQsSOeBChwpUhQ254GHcnvWtRY0HcgkZctYqTOK7c5VNBfpu1MMY/51niFRq
owdn7cZgYvsyVUhHv8Q8HB7SwJZ3IyWYiLl6V6Mt/ZrXWBMmxAqrjJhtizbt8i81
Ql2wGhbr+oDTlkUru7Ea/0SctKBUxDL0QoU8xW83k8S/RFrvr7SliLWAidtIkH/T
GQFBATWljEohHS8HbJHC/08epX9Ka8F8XAHSpjhcVhsBWPw9JtMsJVvwVC2Z0g4k
pf9w/LtmTjXtxfvEmnFXIWJ9jJxGjll3OexCYvRLRwDMcvw8oKVrwzw4rRydybca
ewVBvjTLKhrKF+IeVO4ebgxJUGUWTI9Vk7iLtvXtma5y1UivssiEKVEUOIQLC0Ve
1EsmN1OzuUi9bT2LmFhmW+jRxItdcTWLobZni2/tql4NVs95UPQ66X6EvMPTdf9S
wqKM32i0Hk8QBhSdrc+KAp4X8kEVfZF4MZRd1pLQOt/EbIxmfR0VDZVJqI0Jb9ma
bH+9/OPdqdm3e/ShPMNu5KEtnKHz/Z/sr2YdXdlpCj0Akq/zpvztpiFn+stBSv5P
IyoEsUruzUMNu6YoJZLZUqPXLlBcdbGn2myihJR2TsVE7Rxgw+jKMyQt0oj5fEVf
IYbJaOqfjzhCk2WZ4RyLuDO+SLDjlqEgWb0M6Uvq4y4un/UtEamVxgOfU+yyDogI
LTAHj3YKhS+t6ABgX/z0/0M6jH1iKTTDw3b67rukPDA9po3u1OhXGMssSK+Tho7n
L2wpEatDw4OAc+qFDiA1F0HnSrB+5HDAP2pfYu7WkIGR4WOCu45Ko+kozH4SEYAq
DjaBFWERfSaNagARAQCnLDjmDPzXlJJpEiB8zCcldrbClCF1B2vkud7xtm3y7Jh0
Q3PBrbw7+RZqktWpaU5AxOf96rjlR1eQ1BQi9rf8nSlyW7If0ugK0D23v5U6aVtI
aEktnk4C08fSlDDCprLZjY1VgvqA/xypWtC3Gko+sMMttYKlMB5DnP7R69goi3Mv
oNwj4dWvOAL4Wlaw2wNLnKgxDXQYoHkaePeYEfKhsp7k3jdXo0s8bUu8QocGgPg/
Mk9WTmoTX7fYg5T6kiMBvPZ48XK4Wi/VlL3+UrXp5nhzxXkFgC95vjkJe376kggi
qe//07lK8xQq0TRF6whp2qmwCb3TM8l9EJwH+mPEVd1TcpOGZT9QimFG0v13vk0q
hFkqjMpN0uEXL6aBvdHwLtKVcYuPrXp4IoCuRYrGDdy5CC7FguadNzAp1PVr6D+5
KY1PswyRwUgGMExVAfVi+kuGbjxXKoODlft1DZOPLTejfAMnzjIAdeUCQ1EJoeyY
F3IYXcZPfy7PPYM5SnT2BzbS+ycr3wU4PfYSnmK9y82W8fv7l7vssTsVLtGhvs8S
uwF1G66xxYfYWCTtp43kK5hYemoscWlHv9ut+96RdCAgp7WiMn/BSR6pgTk+hk4Y
aipTg4DlUthJnkk0FqhmNCPqhSon6XnGBhuQmZ9XhoUpVLMibIhZ5TF+cFkE6QJK
dqdfv1/IIPX70u1OJ0MElda4lMbh5eli6q9Kubsn9Oq6CdK0WhHyVzY0m5dhRfn4
navxnDLm07UqIaLKR+9u1U0tTfVyqerNBRAYYSwkmrRJIPGrzs5kzd/avuAJ01yM
iw0q6jahDO2yH9+uAaKwJspUBvHpksY10eymzxaICRtcQroN61KhTP+l/PHhMD8b
s4irPcjyjFWvwvwJcQLfOQN+fx4HO9m+yhREv2aLQu5y56NIA/s1/zIHbFS9kZRS
GWB2FEZu+eXv2PLlUsah+d25yUyJ9CMJhJFelPUKIfOXDs1TID1ZiZjGyOoYZoyb
9pVv4tZ3IQhmnWOT2Gq0k8Ac8+aRodM500208/4ERT2OwxDLiMTvfmyfkyMPcx3w
R9Mmg2we04NljcYmGiQ2cwX9HGhzEJie0Ctzjxky0Ekf3hc7ljA4MMQ2f4TfhI5Q
oTsw5ZdTl/vUPiyGm2vxWtkHDDq2M1/DQZlfcPHRtVJA0hN6kJrOz6uGNDDOtLjw
x770WSZZlVdBvG/oWTDumc03yPkuZyelEyUVkw9LxYPzEziqRRb62LIJdb4zQcOG
xJhXdDcOpzZgplmKVvBkkK5C1iHbc5TycpdDvImDZJwE7Y9WyoP2bJ/uH6ouMcWt
1hCCPzOD2IKNaG0pBaKGv8pcWTbHGvokZj07TVJXVOovXQF9vNvxwoyWQGrWutjz
AXgiR017CINOrxKLtrqpI7/tzCdj9C+du08UGMljzLOfB0ttgx53cANMX5UZRBCW
6d0e5qYWZmdh9NSDqSwBWkTFBrCSwWHcE308D2J2TEBAoV2X41f7QeOxlFYCKAZi
5QKOICWk/QIrSMlfzRZxLlWqL5+JaA+C2nyiT9KsClwFT4t7kugxuAUFuAk7gohs
Ggf/83kYsqzOmIZoEU0M5Dr566uDSdMvKm2OOvtF+GCwt5LbPaEiH3uEFH58UjvV
Q0eH1AujI2KLJYv9wcnpUuj4JI9gDUfLzoNCchxUhDtwf/d963V/UXS3olzwwDzj
hMOiw5lLP1k/vve77eUAfABspI3WUtNfmnFTJ9czpT/UN9QBmpXVCm/PiC54gGZc
phstrYrOqWmI2j7LSaKK+P8+CWokYs4pqeBozsUgYff7T6H+E0g8aslULs/Q2l46
7AxnVPUyItzcmjLSUT6tKLukI6ULNih7uR4RBJXP2wsebyLDrHwUN8+7K5Q4R0o3
38VtHY0qSKEAHPSDjh4rAYSjZApjZSe5wvQAKg524Sy5t5GvBLoPUUXlA1D/wZzi
ps58z4fAh98WbXoT0u+DZESlE/NvHqomdHjSnASPU+8SeGEGVX+cgPBhiHwq4csD
c0KnAF5L1nkCunXJrrk/iQxudvF4uxaZ7qGeVswnY3v6DQm754fgKme5T+KX6h9l
9q6l8IHq9OxbvvGySPcZvvkwQy51NTVflvXAbDfoGqj0PsUkNIGOpPCdu1Q15Eso
2ORaWJkSe7JrXa9JYfPizYvPuyEutrWVsc5JrKgg/5nb7Bt7FPO8yDKl0bgelJWo
m6n2tgtGUEtPfGENxtXNbsgdj3teuafarKflCxcRpnao47oEpR4RlWT1uy8DJu2i
DRi1nwpYFntdPPp9DNGMYmyW1WjUU1vp1hmKwLeDk9JBfPqYGfxXSYxPNNboOPqm
gk3r0pQs3C1sdFr+iJuEENLm5f7YdAQDUsePZziaueQfZ/7UAgkKyQMJoyx6poE0
gkFGt6WdY7latAe5DKAhDAJtTFcblKHkN4KWEJpmaD9u3fHr4T5RBQlPeVtfWj9K
rgIYAKBSslLtped8o1/Q+FhGLoe4+PsenKTOPiGuZyysXQwXODeJI/dPyqLqNp3r
7GQ/yjBA0Igkk0CPvqc+rsR5r9CVr6pwQNTODr6R4v6iAXsWTtVM+m1y6OvkINlb
kzXSUgE4rKMBgd5RTNE4e8kiau34Nsd6ZkQr7CBB65rmWzyu5Mqk/v1WB7SS9iwd
7rrM+HJw4CcOICvke8mTTF1DigPkPwfDjvGtQHr7WyrKhB+z+xnOvQtrRfR2T4xP
kz6tlEdR3gKXgbRDaNBwt9ckPTKCWZQwroGfhCidY2PCrn9p3wnGVom+CA8OYDpA
2/DGv6Ajn54nah/zIHjlAQ9uDKMdxQxl3OmNi+u+AQkMP8Wfj5JTk+Oc31rCkWHp
zicUk2zUyep30NnLzwJ89F42bmUiwVD66Lfn+FKRkiTtE0DpbJPNpiOSPwXHWbdY
4Tf0mZX2sMBc5p14SIQK74M11tSGqSAEndsXASYacrVpY9XaN4UxTOUoAXWTak0O
7Sc4LRjuy3o20yrawD171bnmJt3pBTdHscv5nuvZ0ltZnBfoboE/9DYToInb+INp
Ro8XUbNAbi/10ajZxMk+1Sskc2TOJ1tP3G1dJOWtYf+XHRWwIcn0cKrvcV3yQF1u
ZnPrB8VIrBGcNrRZDxAojR6qNOGSEw6mbEO/hlU4PCKesYRy70PJ5sz3sAxpzyxF
rIfPMnBbmXOfeWHR80iC9QmBZb4mcCTyiliALJmpxVY5muH7y8fi/pzLQecFuLWN
5cSmqqveRKjXUvYr3tMJn3pq4x+j8R84mdOlqcL4peN9MWqRttcfc1hXvLqsBLX6
UB9tBW8t8C+Zds5mhaWKMXQbfI91QXE/ABXA3CTjxrnWdkGBtf7NnSbbFe3BOcyr
Q9WQKIVwE0rDM/bY0LUwpzVq6zQTcx3yBhq7f2fEVg10QEiOVhOxp6sYvsfp5UqU
t9f4dVw6lk6jjyEwO1/vQrGh0JXm8tHt755q6Z1RwSt+k63CpC6d2jl3uuAayxaQ
Q8fLRfPjsGDsO3f8oNwTJ+cj+/GMnZ1mXFNGv72SNwW8BdriZIK+IIBpQHUYIRW5
73aArrTDLVTuzg4EJtIM/JC2zFR21YkxEkfcfK0+uVNS5YT9l3xFgIXZ+CUPc4Qr
CRGAImvX5ycUyKKvNuTKvGOYWIvg812m7F1SB3uGshnN1MUM37CTIVKo4vedPPl6
yEqBqp3XoZ00sLHgoKf6qEgTRTnYa0yRUY7//B2E1gbuublUavLdUxJk54x3Pn8r
4hwyjoU5+pfyooYqEgvfi4orCNZMNIFiQvaHHLxZl1/r51ok80qQPmh2PuZgp9gX
geye/qzB2Au67wWFL7pHrkwDgBoaKE0FrrHmnc1nCpThBz9bMkvsegxlzSWHnHG0
Fa10jnq+3KumBgn8i1wbmGGcGAMJj6f3dP6Be7/7FP4IOeQBSNgmZtPpFBD6Di+7
+GjH2nc6F7Cje5WbKRBXf9VrLXLfAfmlRYwsTu8/AJkqr/RMqEqSzcMBRTNbBZu2
gPjNj8K2lthH1bEgrHDDsK/MEv8FMuuIqMW/asJFWZ4u7uXKlMUBaazqCx1HA2N4
cNHTFM0EI3E2ULyjVA2vfUoaiHbHIz0vuMirIvVVCb42KEa4s3P12CFP21mSRk+o
gUwnKVI2bsGiqPmIEU2Js0GhNFLbCaRZ+J4Z7ypwRaBZtfUDy1Db/RSu18Bd8gYq
4UvMsmgde3BImJJhssIRH2pCyaQQoAhxTXm8kszK8wJKS7o0wKhpSK7SuxjJq76b
qestyYdod0d/vU0PyTrVGbTyeOIBoJNavPiNH9xbGVxuqZaysw5yT/LZt0z9GQZD
r3IrvntWe+ondVEoAeY4xxw62YF6le3k3SuGqMVPeLRLGD+se/iSpEyzRQmvxLhN
9oBA53Gy2cvVlOJJNq5/v/lJ9qnRcXDWPyycZv9Xhuc5nq4Xt4EvyEx1pYnuC6r5
PovuU3OHEEFT9AdQPcxTdryw3t5CwVP+um0IBl0m9JE0+0DI5zA+pG17w4sjRScM
8ley1bYhn7EJ2WaatYsIMYKpRLyloIgPfhO6zEFrXPuOPRfrG7bEqZzWCACOQ0bA
EUArgFBUT903D1Hr+L35NEfwsMVXOChuvHZ7Mp3aMOljpqKIqy2n12hAvgmagh8y
fV5eGhzILn3l+Ybhqc6TaUPBH9kGb5IcOTWmItNEavvkBTpplNPUtp2nKD/qUXr1
m2DWiGVRLjRTvIXoXryDmORQBGl+EX3xkNl4nySpIQWAYBlDfj2sF5e3JGBskX7y
hs6/8OU4DpmlCip2u3naTnBgvhvuQKtRdljcnadVHFvOFetKeHnBa6UyLDq+wDay
QZVRzufCkAZFPYci17w/gPVzvyBV0N7Us0q78RTUqFeoOGt6P2NWPEMEYs7m4FfA
JdgbNaZdsG6jBaficGBxQqeh+Qw8AKA9PYpThtCI2kRQ942AxFD7AVuV1YtmjdYU
pv3jhbebuo/JMbwbnfwb6zldUYiOXZ/wqsiS7s57jZOfFQ2YWpKsQ3gYf3IAuSxj
uURGEd8MTMOTqyFe+f/xIja9m8bqZmexYmc+271F4nIR9xPqaYidDY+Zfrc01yf8
9TZDhezRZnPlh8VfbysNgbxzjdOEnhyCDJWGS5M87Ci+eP1qeOuA1YFdPbMxLZbs
25CoZAK11IBLnZ5hG6U+RCn9/nrqlDrlhUSPz5yAuK1CP/8O1fQYT6wKIhoCcN/Q
9lI5xY81LwDHem2UgKlCVaNDaxvZ8r+jt8Er/Eg9SyYEjrv4yDJDMGeKX/D49qM8
F6h6IVhQZkivxQr6t9I17z+YJJWFrdf5Ox3S+5rMry7Aby3+9qjlAHo4oPa1FEQH
gybtUa8qTJMlr7hB/tvduA/H8rQbNoO6AtL7CYD7PyJx10X+KApXrbamBl/D05tm
RnJ1MTej4H6k4z/wUxb+wv0ueppgaLPmIapZ0rkMgxBpHp4CBw8MapZWNmPti3wk
Op+BTRyN6f8R+XSmpVq3z3u/lcQM9bnk9WR0QN+xDe2wnvX+RDuVM6Iqsl2TecLw
IJAJlV2ES+sVScu4eSgFTo4N2HylkwyCCN2o75F5/H80F2arXbDNDGuYgJhnF/lt
ZwTsz88ypCUyXQ05PtxAHlPx976Z+thyWCffBzfYpI51nDkn9ptNXKybTedZR0vc
L6YwdE7lCd0TIZpOd6zYqD6i3OkxOYWi4GSOuTQOduh0FEou4Aa8c4+azXJ+Nbv1
LfAHX/XfrSvNNZsXFzzrpFTxzN0UzLyCFmIglK0Ed43k/P9xu0Q2VLQgBeoEl4Hb
Hut2Y0GNrFcPs6q9TlNjii2kZiqzZxK/OAHAMvtOqepp1AHq24pFfVbaxA6PLajT
Vuvy6x71OG3AVkJ4qazFpC8X5oxCu+ZHEdHKigNIL9GtJFYEALn7PuVK/3J/MiCC
SjjfHMrUdf2xnK8WWVU6j7EnI3PAyKF+ZYo92Ay5nQGltbG1QnzS3BGgJ1kY8V+z
57KNG6G6pfkd/8Dj9Kfw+3CdmF1FjtbginKj4xlTQRZk7oLTDfcE7VMPF0YVWnLg
6eWcihuLWHq3mEokhzB8cBRjqR16mWNdEFQUuyFKlkCvrNLIjLigVcedpgS2lt/m
7tU3REjJN8geLbkXr+ynqnAZye3SM+xnZK9vCHWaHS75qm6MIlvpfzXxeZ60Mp26
uiyGsCC+svJqt2UBYPEQLxPBKe2Wg1ydeXYxBSj7QdaDNJPT2DUqBNEuIDqbkK/9
+w6HVsP9AAmT0phpLTwmdX63dSdsVctEZkMkxuO5WZSal8rEavni4qKpj88pJurD
vtL0e36dhkhE9/DMCVqAj84CrZpP7z0KJU/3TfYsC0mHB6+qJ6NMooldEST/hTVJ
tf2WWGKst/1vZ4z5Lo9bZDDO1T97NfONmYC6c1FtW201kdNUEWTh484cpXDIRbPQ
8U3CaUXxG6YhOELcSPKQYHYL3P3U39nTigGzfiBfd52jdhkxLNqv216IVO9dMkf7
hRlQ0k1BN1WkzuRPImEn1g0mzCSmx/aRLJvEvWg68sEjiUy7M5dD8nTYM9Nvxhk7
CNPmoCpXRsFUMM5dtXN4u0PumHQn/N/apRGmAkwBvwKC6suM3wytXzvXx1IjC1F1
7nPYWZET3VgHY1xMLf1BRNZgElr+sNsxw2eno3ihk9fXT4V5s0LSJWEX/2hnedqM
og9LspAPAuvyUYrXkf3TRmrhOXOp9QfVCT29uhE+4bdxTkdZP3YLJ6QrNhpnbyk9
RTODvLXrttR9sqFHjo2nOObviJTJdGKj9bhubyilCYqh18rfR+5ZhXP9FLWUZHlC
9fw77qSQlLS+zKAKIcK4AFKi25wl08anGhX+nXNaktfyBpHEtUg8FV1owabCTXPm
7SwuPYNcpYy+vTAGngi/py3jo7024YXwSQ9YCDpumNzWs71OzRCBL+lgEZQRPaap
IPuhe8LDFSZysHYZT/CFdwGHQJOkjVI+2tH9CfBHBqehC+tC2GqSmxYW1h/0DEdW
sqJYoXGk8CeBl1r11CMe7nmRYnOLR7PAxHl0HyUHdNb7nmgNM1RizYW/1Eu5c6fA
zUOiGIX8NLuC1I6aXsGBwbd/7zAJXm+sR2DqOf9FS2Y4fdiW8VdUjdqxnTtOYZ1t
qlK4SBKfztydrF15E65/r8BCA+xVIZYSE6EtES7oYv5mwWUL66bvRNJ/YRvh4WSu
3/3nYr2YXiVP9+8VIHMKDhvmyS2+liSwYDDWQ+tfj54dj+/BS8+PVYJaCG5v6MwJ
rFCMBrvH6iosRH9jHsGR2Qc9UBcYHFomU70aB31KliZa/4DFJxchn+jezejs95E1
B2apfopHEiX1zhDBunqCaVA1NN5LhWfjHfxO/8vLcjzljEVN1KfVp/HZ7F+V+pd+
eodJ8yMTmkBUHDlaZls/0qT+QUvynEHsKOYUDXpY7Za7H4D3RSFDHakOMBl4RVv2
qBkXyzN8y7v/2STg9xsi3Sfd01hdz+welTdT8yFYVQayyMVEEj4d7d/xiNH05MP1
5SxpEqMy5ymZRdcZGv1crangjFalyRu/mCe8+5MsmcKLCH3T264dOAArjZZxTvAI
Y6yzF62gRCu9kAks0S1dQA0PPiUi/Lh91kKFT63QN+Na3T7it/2M2FlLMMvAEWVm
ONCEzw+ZT5/hbLBFijYJgczKM1ky/1EdigIKA1DEy1SfcNfoe3nCSNihTM8xiOQ7
DDwgdAa7d7wL8Gtq6HDjvXD0eDWEZLX/KoQ3IUZKbV59tzItblSqWzOp8UE5weIw
WmYwBCMQmgM1lzT2YyGUSlK2c0nz1foAm4lQ+tr3mCjQsF2KJXk0im/BcsxNmn7/
dh765BAtaesFCbTYTC/Mxf6WcmcieH4kzgFU6ObmG0g4ShWEacSNXjTYzGqB8JN5
JpLWxrWqHoNKrJqWTetjsvCm49xgbg1ztYzrFO11YypC3OMlOAna5qoLt5OC+eis
Q3hB/Y2EpSvA6MWD7lq2roykSWeUtMM6Mig3A42RpdbC37XXH7rNWWbEHfnt8SFQ
nrZAIyFcodXm4508c/aNhlKGSqK4BDH/p7RcyTY36Gc7Dzm4IrBFMJsGuHDsBQ/V
t4Z+GLhUMle09qpV9JBYNkIjt8XzUuJJ6Jp75JLzA/7CPoYKHSZ+uwUOyQC4uO2u
UeFSMV3E7R550E26Jrhym7c1saaG3ixVTX4QGqp4K9N8p2MFe05/WocHRWUKuBk+
X3ZkKFUiZTRoXUp1mTVPEmIKUaa+xRkXhYsFdXPDbObRCIOUgo3qH1Wqxqfg5aNE
HbqhhHsiO7exZautxP/PMysHsOn+MEjiC5Kfh9xwxHWkdL5fLN9isz+iWBWGrpig
sbihcQQGfzFLs1XMkgvLBb3+TdeRkB+ZiOln8/OJbLj3eYY0NOPpkYz6AgS1Byyk
vrkzafJbkKbGVHPtW69otEngAPx34Jw9iVTB5j2heK78kk9tk/l2QHww76FrwB2T
7zOiwRhJVXXEG5YQDxyMniIbRpHosqGckQBuzJjQKtQkcdZXWQPTNUuyprMea25J
jGZ3CX8vLxhfrynYwHfiRjY/vqTxQZS6aw6Cu+OOJQx1W+1ePzQRfXjM6pNYVDDL
DsliEdsH0cCGoSNEZicBJBi2RJIQrKhuRceNboDwiVZTAtVugRYjuttHcpruXA5X
Qu7PalhsbDQRy8bmtujRSHdH4bABNBSBbkSas9WklF3GxgpHDPqRl3UK0TSNc1an
dCw6DoRlR9wouefuPjCKKegM+7HWK/dRy3r9TqW2Ip7aAlPZqRCxcXZsll8rg5cC
oOZKf9qDUX1qBBohb5F0KvcragRrpPWEfRCrsSQEf41VqAt1klbBGX1aBjfeJHe5
9aTxbzI0I6lGsZhBVSV4kU+kOtPdvuhKj7NYxAEKG7KoSjTVHYpYTOuhpS207QjD
YfC2BBEeFZof/cyMBMsSMMAWr2Bc/XGEUoLJJT1hIvcOw6MjHKDKJ4VUmYG6ACvk
zWanx869gh4lzG5GdwbSw/upEM6UF2ChXdv0Rdq1duZeC+c9InFAQAuorJGaPiqP
GaKC5mPG5dyv2Ti2GRFLfud18M1tgds/0cfnuKxwbtZHZr8LCvRRffAqUO2E9hY5
nhq55tIylWTzXCLKkghEKOKQ/q6UOrNAZB7whQmVGI4hKuuabbWMAfIsDEJoME+X
qygG+Vy9qDe4mGRdAVmTRJ71FYeZFk3ar+E0Qk8iQV1AqQQjK+2ojDBcvhuNiDc6
zWD6jFdX2AUrQ2cFPMVvLMepowjBb9LtLbLTEIKVIlI5S5ByfH1TSoBNLkUAFiKz
n6jgzCK9Yt1n/GD1XYrZeDf3G8wZ2rLexu8ZuZqkLqOKD8YNCfFv30zIE0VUOPKR
MV9+Ye+Q6m2XSJ3GQVA8yYNPT7+iBj5P9AQYTdVb0h80qhXv1FhGybG4ApnfpfKt
2tfTG28mA3hPliKy3EpLqxPFHGQR3zIoLKM+HCypPWYN+OWr3AC8ZrAiFEXldTI5
euTjrbDSbQ3MVLykBOErIF/M3LXn47P0NHXkCMNRx89Fsokt4HiaAqJ5lfza5jeN
XW5ijMifyzb3O2jYcRzIcTK506UWoZ+P3VIxw9jqwcdQ7LsxqXfq2HSQezSDD2gr
Je/mX4TYVqg8Gv/gh2notTs7wh7gmIIv9JdPOOnAW5i3ENySn+/pt+9/4alHH+G+
sTa2ttVhVWXxEKFdo1prhxPwuuRB3qifnPhNZO9FVTJ9JGIuq39BpKI44xaodmC/
Lgv5Ve7D1peGT5cJQlozNyGkBhwvkUyFWLgqvbJ7YFPd0saQePqzkG2UpHJtD05f
SUgEnKKJ/xokYLII5rROvFpF8nC/31Qr7ML6i8a87xCTNzlntOlZYEYHWDnlPrnV
FN49LdNbntTBFNEEyL0LjNed2Boh9I6wO2BAMGWeKkE3lILyrf2N00oElRdmbcGI
XgBaCRfq4g/HQsAaGXefaOiW3yPDK5kwqOJ5rDONhSi9d91btT7GjFP7Iw/AqjuD
eWxl8xWjn2k+wXmCPHVZ/91/o064/heGPgo8qnvVmxgKTTZDgrvn+6MLNTYyq/kV
qrOhUn3HhJ9W0I5P9z9pa+2eyku6BGMFhcJZFAaDOavC3jYjnnxDbuQ2qLsxZ01G
a9crcKgK6IL/rOA4N9KvgGfWA/RXOQUmXWAn+A0bYbFFcsO4nSc4LMP4BR+XnzJo
P8yQS5Rb6KNjM5Nx3CRA8DzHewuT/uZXKDgQK7CAHgJiHi0wO44yw+2EFe23nzYT
vNhliguTtp3+NdDwbRWnIhAP/wT55DS2JvHJf/aNT0PWt2rjERWkJbxBazZBdGz2
unEmYaGp1ilpDeDN6ZLQAknMjRl5Z96aLrYNj0UIMhRpZnZy3LidP4l0k3RveVd9
JgwyBCadWr9jO3noHqg6KDIPH1LpHvhoCxzeMRjLv4xKjMFwnQYWweV8AFs+222i
Eu8JTYqBlO5OBDOzP+lVj8rF4i/QIlQ8kSoWT7XeiafNZoD0kmQz9Idx735afFmP
jevKc/rqYblGTYyufC44FGFniEZeYwYLdAT2TieQDpPBCvLJsruXjScOnWCqTWss
b//BiAwYGN9U4KK7PMIGXDxmQTeYpEqGSLb7vLSqN0/ehixka6o/TOGcqkKVuJW+
/HC+v2Jjp8m4aa4aI0ofjcdKY9hIPmGMA49k8u94cKXfRlovJip4I9ZxZic1BulC
56y5DyDfQeOeyZhgNabodI7smPgWpbo/PJAYo0oCn77zAg1PEqnbdj8774SSwOf1
cYLntDMmHj5w2c1wQq/zXv9RGWnSmI0hUv5tv9nmG8OBzBNNVKg41jWafgooyg9W
nUi1h2RMQNVUGVPhoHT4dCdJtCngS08IXBWUx91ydNXhraGuFxGu1abXkKupS71U
DBiZU8lyNBOmAnXkMvsBN8jnOUWGFA8ZtYEVnN3xFcazIffopEu83dDY+poyMjME
tbJ+vsq8wuyZdJl4Hz90yGv2qqvQPaXI2vIwrXfQtnL720Us3HmenEwty/Pmqu1I
y9MioGGXlSBH3J1dag8HWPKLia7Yz8w7qsYcBHAN8P7OXqzNzHVRxOfXfTaJ1fNq
tJqbbTTtjY2R0RHw8Qg49/2cGtaNSNWAc44iCILdx15731mF4jMD/qANflcb3zcx
7utI0q76y+v2ObrcuZwXFlfW9YShK64gojWs8aUNWB6SSE+zqmeYVfEFCnlbjp3Y
diM0mLN5Ch/r02fSMLvRGBL3lGw26uOk2KQTAkUbIU51kXhoWCady3TnIypV8Ndg
QoMsmiOBTqRvP4dasUi9U9ooyNqddL+RhECJCd8KkAxS17IRqZjhaOxZU9rFQai5
Oopkdy5l23ogH99EyKXxNUwTS++8iDCB0GH7CUTM8YeoZfXdEnPlrQfbuWfpWklr
AS7ARBmf/JTJJVFAdH+aTfbacmgBcQPd4JL69x3la0rRnoTHMS6cvUiUJDT7Dw2c
/4J54cPuTTBP5Ur1GfYpmInWBkAqr4qjKxbBRWlNfW449rP8jOtINhco590HUB8Y
L6hj0wcDmEIWxBbS1xlISvXGDV5WOwZNp/jtzRqeWlKKZPHWTzfC1c8/p5ycpN1e
ybyZXt5aK2rUs8iT/XYRuam6JptrKaDk010STi77ja6/w7v4vctYun02eZM9yz0+
IJTFZpb6GbSK4mJChFfgwAUFBYjK1d/if7FqtkcVOJEREk8Qlc6lvQ6dOJOGXD8s
WcRJqBItDzT5XZZ6lqNjYDJYVVEo+vL9MdVNsduSTrVh3V529v2nLmCKhxmkaKD9
S56s9HT7u513d9uXJMFsqjKBKiUIcYom5n7TrbgxgLDLu4JH5Ah2xOpuZw7Psv4M
x+xM19byEUyD2sxrkR5jK5K7HR+B+FlWRCgPDBQouOi4ER8Q9FUgWSthT63xV4mh
TEI7Cf7L78p+CJ6b253HPqYTiijuoz+VU9kJh87a/PIPBth4tBFxvjY0MhCXh4+B
/O4axHEpHebYmovfL++2WL1kQFIW2tr0UY8k08ZiCy0n2pJ6+6+12vR7KhiV8v6u
I+N2Ms1ucmkZogl8d1Kn3uzT4aA1JBVojB9k1GN/jG7fDgi8wLemAYvreitoUICH
NaxGEobvYF9cHGDwe6qrl4G0nMR2z8wGE2trQi04bcuPwF5bejFY4b9xDQXf7xrm
Rd9AhpgV++wtBRPrqUSUgscdqABvpSTnoFY5hJ2QyF7bdHvza/yUBW1pvfw1A0L0
ywYaQmWSb7/1gGS7AUCSkusN9Jtl+wx5JLFnCZlTeOhGJV2coktSVBhSYt9YnoDI
8TmIPGrL3fmj6KOV61mCPofS6nSe6Q5Ey0SSvxXgM7f4SiYFHaHqppoSEdK6xjq1
t5o1yDVysEEKtEbS8CMHB6NBJUIs7zTfBA8PhDJBHkftouBtDIZ/sPmd+OIP1W/R
pLnPRLzMPKnLEXiBeVj9f7Lp6uhrRPPRz91no6FuL96RRpB4L8HHikwfMVUcGnmK
l13NQTa8bGgfMYTnsXps6DeUD/Dh5MRV2E9XNWBjvDg59dRqUM9xNu/CTtgbGRQJ
fCFBe7jOeifVLpT5u9YaM5oNR79oAtAzEgtYpyFC6gNd19USLmpKAP2ExM9oUIwm
zOxSdO3S7FpPoKhTyNrAnq6xW/3iZnnXls6JUehxXQAhsrINX2Ivb/L6u1d4wWoa
GshTwXam2hhObAK6KEIZA6q8kViQHeethZD/+8R3uoMLGuRe69xXImQQDr5yCbsC
yKYRd84+ItMHGla16kgM4UC0tc7srY51OvEc95Bal9UIR4YDbloFPzd2+XPqZ5s+
XGgUslP/BEwJ4bv8bvAogcBm/qQ5flQ9k44egokRs3I31UwUP7dD6qo4lN6lU8FW
BN0/P6EQSU+FUj5nWY9hiw3YEl4D+ouHYGbCPp0SxB8fL1m2AX5vlZGDRbxG9dVf
e+FnFWklNngqfO7XV7rAWdZHy4xeSRrvMsmdPNmo3XHAesJ4OhzA77ens2TAK/jv
GtsAyV23ik3K7iZlwCJmGfPoGa5OCD1O1VdUspgvxZz60/rD3W7w1IkCS3xmlhMd
FiMvhxz5734smjMIOjb3UXuyiaeS3USKHeLD2V0wnRNp8I6fyT5E+KCIC+MHj/zf
xlrubunFULZVQL0SNzB6WnFwG0YkbA9ITORLqa8u8tl16gO6JubYfqM3qIQj1wDS
5A6MYzIT/ux0rsA+IZJbWl8mNHGq7cF9Jxpir6xabsF7v5+z/E1Oh8PQ+GDFmJZR
uwddWqO5uChFO+BmOncOdQ7FBLRfPLOGta7Zoi64KOugnQrT/rZiQHTik01cGu0z
UTIUssIRW9Y1ZfwrKEHKcbbj3WtKkGuEhRdDl2YLN5bwXy4EHw/a5fYdRSu2nF/K
GqMh0wotWmLj+AEP5blBPZhfiu1fDp+BZRHgntnN7eiqF/66lR1/Ujm+NwrfZrWo
C90shb61CGrTQHh8cU5Bw8kpQrWYUaON+nZ34PgTVElx8hYOTImBSf4PIbJeIM9J
u8X7r6Yq/B9QC2T8ZZHx/vMpe0ly11DwxQsLFVFGHKZ7GfavWvr5CZPa6UZDPipr
UPH7Fu/gC3lOLo4sbvlFYXNIJGyqioCsD9n1bYp07K3dDMw0Txh5jwTLAX2NVvem
GEoim/5k9gFznKYJDE+sr/sFkaQn51B470aczkab/qgD/u8cY7ghceXetJk42DO3
Mb1r8/ADzXOOejAJhfYp9Ao31gt3RBoou9NyQQfEK5u2DHVfMmQ/IltHzuuMZu8A
djhMKqDVomlEj4gDSn1lljnw/r7lznbN9m2OQ9VZtYMLmEpFO8q08vHTW14PKcpP
x382z0aN/Bc/oofYJsNw4ax7v8DY64VN7XR1xhcz2C9wSjq9G2+8Oble+sgxv6Bu
VUO9MHOIbAek4uBeAo7WKILt6jkrz6MnY0QlqIhkgAecOfm6VY2h1LDdY1WVAwxt
dySvcONP5g9Qw7goa+pYCp+fnIuh6HQr6cqg+grPj1e9AunPWpRw5TkkWpimdKja
BE/SkeOPsiBxVPC8H1nJhO5P8qB/x5lm7ex48Z7otwFPVoaLhfsRZWxSwjJ+nYtZ
flA/jRKWJZ3T1wougjTybY8kIKHvn9z7US01D7n/3CYte7Ns8in9zupikaTlOnw5
MsaNil2KkAs+xOhqEVFdehdCf03Cex0Ewg6yiYBnWgo0mIFf+z2UjOtPGMwdXYmk
x2OOEG+HU1kUTyEFj8qyTa1ImigV4i4VnUgZStRcPNak7s/WVQSDrsKV2dSMQlks
v9U3eRAvrfKZgYYWkSbkF6HrfujyUtQO5PAxy5/tfJ2aikpZsrm8EJ1huW82ozTL
tfVlqN/RHt8TnFauhsewMBY7aQSbvBRFTaluf33Q+CvwFnIIgqft5VkFNrSkigNH
xVa2kmQ3TnEySpsLX6ODF2vWz2JGqazSN7H0ouuBUZPOk6vOUvQ8Bl52LoT6ko70
L8MItATmJDFnaLWVWKuIDJGwqz6xPjsi1yvkomr/qH+dc1RaTxHcng3ESP/HGIsF
4FccshFz3fpD/AGzrWomoFEekA3/kCsX6JCqwoRHtfF5AuJ7mRMcjet/Lw+S1MMb
OCwTa0PT/+OYf126fGJVIwNQmXuUjgS39qbc2qg97XCQmPLumriNGhRTl4VlR2vd
1QdpvVNh2pXQbr+WXAjHftbKPXuQ4KqhGiMeapsZ4miju5p3F1vp2jLtzR5WV9n1
mT2I2WS6rMZ5eRLPny2UdBTpmFeyiwWkw1MDHWjXaF3klkozh4qQ34ee72YMlMIZ
jOwIXi8jl0G/hvHxt50AvPC6Cq0nFf0VOLKpHWsxjilmjRGWN3n6SunaOwgJRRVZ
iZnWymQY8GgxxQsJIbj5/aGSABhLA5nxTZP2KoEOEa7DSsvHx3hK6+kholLk3R+G
pzIBmmgjp/cezaKyRkNumMnnuFVkHr0eRkX4ZnEYuv1dq5q1vgy9KGHUs3M+/y69
joE7BzFw9s+e37ISkxfcE07+Ap1D8GSRki86xfWjXbfUW3vSD0PegXDPDmaxOBsK
0aGAdSL7Mci0D2cupQOOOE4XNV/atPnwuNFsfn4TLyS82Kf3OOr4wu5a4wILQ2Mc
eonJdt8JrZRBUowAknrrNHCHkTzK4ePrfh5E1utTphSa3EgoShLX8JJ19o72TnLl
n3ilQfYqnenDFVRxvgRhYJxngP4igHCiwCzoWLM+8gP8WvP/K9rUelxNzw4PVr9g
n9GGL/7MlSpbQMugpNKJyCxhA+cKG3ebOtCeUfU5mRRrLInClE/rBDAuaMTeD7il
DlNHNjWE9K7WaSJ8y/FDuRNdjmQ1qoMO4P+jFRbvFhdYaZscsnSTYo/Knr7PuJXM
qzlEPSEd0S77Yw3eQE8b8YMQidSO6+7IwNaJtLOeTSLv3mMJVdtJ+IU1WjDgrdwC
WXdvIuqV7rZHjJ9VUtzZgNjDVEAYQqNq9r/cNe9sBNcIX1Lg/tfBCU+VQ7cZQfMF
lL4jyagaMy/lSg61fdr0PQrIw8FPzOpXAd2bUSJxSl1msGnkKbGw0rVPY41zqd69
QmwDULOUxtZft6uPRJXq6vlvMG9U0ROvssrvve0BGgxsZCNaBVBGD3NOqbtCbJGo
V11D0PoibCy6soRsQ8Eo+2mpTh0Mm1mzwO3hHv8T76TmtZ5ivwpejoiaaJI/mALW
XOY2j+9DcMGq/C9JSbKB3n459sIpzS/E2j0ueR1HC5d5JfVkVBpr8n5yxQt5TmOm
QWqeYfUWaueRDeWv5f3sAlwvBu3jt2jGnkVRLOu/+j+6Sv8D6f4u30Qt724tO0jF
dvr5qqhcEtFQDXDnE8+f8GmCeofY2nxGgKB4Fpi+q4Z/QIGTvtrkm69wRcJ7WhHe
BWSwfO7GLCI3f+PCKDHtUP98Vaojz9N1uLexVSeWRHg6uLw8PVfyPY9GYZKShKkN
ZHmXKwThzSsnAFV7IE3akcm5eIcFmcSvswoRE5nAd2Tq7X/AZMYgjMg0EjgKba86
34427MkR6BAsJcYg0HwWA46kNUKtTAFiBg6a7z60h7jp5s6FunbaAy6P7cGR61DS
Q4FM3+geHu0zayPoViqGYtu1GkOMruXDGRMgM+Xd5CWpn+32k/fd9rwgFiN6FY2W
4GKCnaiZ4JSp7VtnNVtFbwXCZag6eV7jwetgucNM0cd7vMqWTyAsiM4F8ahA/vno
iENPlXZO3pizxBTk4vOu7X6k3uDQNlyOiAO1gnBmf9eTxNu5ME4MbWGt77gtwnS6
UHgVwNPVnR3OMjkuf94di+mV3dPp1MS1VR3j/0ZqzNpNZxgp1Q+0bUZn8H8L+0sS
5e+1W08h8QtTPtbwstWNZnw1792Oh5w/a7LtEamQHgfbNEV8Zk2xpx5/TaR8VWKf
6PLHguRy7I8fzEuWCjmVvAbjLs/i2Gsu5eCNOq9sZHretiJp//FHVyPUu41RnFmu
jkuDG7utfIIZ3i+OGD3Q6NC9fi3Xfod1gUdN6W7ZDz3L5+W4U9HSF/o3v9vR/PpK
NSKEDaJDaYpckRRjkt/lXq1/CxDgBmJnpYj7N8gRYnNnAk3HP5lxPKY4iyQIU7aE
hugNUp7b9PspBFi98OEKGVRomPehp4et38CVGkzzbSAvqfwEOt69qu/F9fFBs/Cd
acGsYANveM6KoLc93vaRxTmQN50Gn3/KGRma1vYQrDF2WbrHxRXrT+rsTijv1nAf
xlNQEcfjmGAvYLDu5kjLKWVH6p7psiLHjC7dXFOsf/Ry55ANKI02sWARUlhWTPEw
LQUu2vStfTrvaH8jeYH/iHOSUxSLfyHbuzKDyXs0OmUDsVrLPZqaiX3vrQjtFez9
wk74g0cKUzRnNZ+sLZUPGzR9mStxrFxzAOPGNYK40LPRLG3MgkCTYyPqEZyRDklJ
8bmFwZGRYYn/5I3wbzKTLbwHnNAy6bMraKGp87w55e+G9uFyWQlw7eq3QaZJQDKp
YkeKkauUYaxZ0jOutskQ4a9+YK2Yb2MfTRx05UhidPboglQyL48XFgnO+ElykjUy
PTsXWEnfObjf9Sr/UHQE54dG2z66KrA/ly0KE1gO6u4KJKL2QmVrMfZ8tbDvB++6
fvM2qpMQ2sQyKoRH8Bd2OhQ57D1vczAM9hz3YwZCcR9Soz8fxF5ChoH51joetyfw
mbbQyg9YQM1TIS1tYlvwM1NWHLoPnrhbqWc9OsU+wx15yf68HnwTns6jDEUpoy+c
H6vgExhdsrWCPenV1xwQI2zpLpPvSvlGpRjeRayjDJqdwQxRUnT6CwdQBHHuF+Fk
mLggg4kn70OF9w4VMoMyQBU6YIlW7VvcAwnJY3CoSWZP7dTYr0QKyf+x19UaXhFa
MQ0rODSyVfSi4tZR2rBUXHJ8VPUMwVHkM5/3kg5YbpQ6K5RjIoAEHBeblTHlwG5s
19ehhasmsG69lmTT+SxZaKThK8XFADml/B5UhVMGrJI87tu97t+1/4+Wl5t3yqq6
2buQKfUsMS/R74Vrci7LibiYarCHhwYkWLSZKL435esV+ApeiKIo29UgdxLzFthE
3TdEvYEvSMFqVIRpUJi3oBSRJSDgB9altSYgkvHUHZ5w7fNDIOdiydHRa2xjbS17
Q4o+tWReJipPq5v1InyUtzHlEOHCG8iqPvE193jj7WtPYC7h8o13bQEx4T9in/jN
EPC9cRZtjBiC0C68phbCV5OMpl4TfLt4OFC2HfxVUlpDIqN6k7qcFuolB0I5tpZv
jHyfzheamr1MJnrjnaSRcCSo4grWuKjhkb7TManTyPBDofUgh1ToY/D7HPT7zhRC
2rZLk6C3jjw8opOcIipxL7AY1fYBly/BC6vOTNudTGWANZnsXwscTIkrg+LW4x2L
1dK3gDEb71bfUlVX3yb7o8GiXnuizdGWCSi8e58AAhZgNokeB4x/l8w7NoeuBiCD
EPGxYjnxSUbDJNOkKecJ2lhtJipsmGDBpIpy8t+e4uMEG4+IZHQW1obY9atNCDN0
+yfb0otB63eaNrNdWLRPHosOchLnBVfyqGhi6ejxMixP9jWzcxHGyZhd4L+WnG0b
QpK1/mcw5+F5tuAq0mnfYeS4QuWhe/vFF6CUtfu0+w6UvxFqvvt22f/yrQZkJvTQ
U5jlrECqEnh6EXgHzAAgwyejFSDNBB+gwRtcHDLCAR682OcO+g+CLjeeTkimnCNi
k15T4sy0Fom3i3MGSS6qbnpoHGNXLYc+HzzIOd4iWiJSEVYlDp0C5xeZ3lkiZs74
9IsRq0hoaAMUfz2rVVmw0hj24Q9weSB0raJNbaoXozwhbBHQBuhk0spa82jcjqm0
YteY0UxkrA7iRnu6uUNevQgV383mg3Nwy51DgH1RSXAxESFW25RQ8iYvfw6pub1d
PnzcnevhDMeskTa2c7kYhUzclmxYk3z9L22+DiHRuypxS2Pyb/1nLA9o6vCbMHYb
BhZIlqCDxKFossZqvMRuTeN5iobG9lyKgTgR/+Jemm/TXe75hfQKcIZttNZpEQBR
qYRLjtHQyyySTkV/udYKMPREXOnHoDqZplooGx9W0NO+QklzrPwC2zt8N8eMZc3J
0ZTrcHx97zhDTCG0hrbMYrTPNUqCQYvnGORbv8ODMBOHy40XfJ4XEJiyEP1Qo/+i
QvCM2oYf/6JBzpdNMEW3UbQgFwiwwuqjvYiUoYGJbQzuhu5SmQkKADpXEWj00GA8
wbHqngIl3RmOtE75d9OHIb5wn3Ucez9d/k1vbM1xWGIY64WjUb0Cbhb6PUEcLvEl
6wVPFJYYYCG31lPL7R79UE4XmEdCDqn1j27C1oRaJRYW/DNjCDWTrj+e8nyP7URF
LCIDBK0Qjg8vkxIXdxnvkubDO+ts2R5/xTw4y0nfriy6Azgby8Wpx24ODuGYHOUP
LRWPuAEsGXiRV3BrVV5FTNoc2aWtqMj0vtT+5BddJ3KAEFCdxyNmotb9teLVFy2O
tOLmmkEO7jEugPws5WFkv2QXaY3ZYmE9Ll7ZcwzlqL4HU1h7nD/lC8ygPhmLiGB5
quKDhiNErG3D9SrlE+sZgG1qz9aicEB3RT4tPuwI3hgqvJ7fM/AwMdhOvmo8I01W
jxSw/HgUmHU4uWHIdmwHl6E1dz8QB3zFn90pip0c1/GECbjZ/hjPZnh5qOI5f2NL
x6dF2FymL1YG4gRs37dO6yeXrijPXrLkJY42SdVrcNjLY16UEjSJpIsk0vaa46WJ
6hrKERYvGCc/drwv12FoA0xCZlA58Rg3Q5YvoyUQbZGsRo2g9HJu40Gdk4tQMWrD
ntvAiiUNHwARbAT8gSP0nWie9MArpk3TbXosBXRZAEe72yVRwETneQotQyAjjv0l
JfMLMA4M3+95wdrPva4MHEZODMlCSABrNonIDyM8o+k4GFIgFuWIEQ4xFG5ksaXH
dg4Fd4Ef3/JgmgUkRwFqdXn3LddyK/LrMJrI8Ldu3dd09vHT1L91Xo/cgbsR6LNZ
w1/vx8LZZbD6c/9UDx+vVlUtuQl8pzYlf0T9+FaRSFtTUh27I4zWh0OJaNXRSs51
90dV3dLWdnIiP6SNi3RN6mdl8z7GVco0jKOo+uZjpxaRrQ+sKXBvLkvdjoqSzW+R
l4lBk505lLXfpOwm0GmlIsZCFtr3GkQ7+1VWmIn07ZMrHEjrL0XKDNZXCuA201q3
NyxioJKYCv4aG8XHqbhLbSKbWP1GPZYSS3eOrzzYyIFBHuvDFT0wEjqzDxQepzXD
d8EFouagTtEwYDREy0W3OP3eExKdJ6JXk+tNLHvglfRpcgrEbClcfBt1T05r3tSt
gZk9swRk8QjQ5Bamn2tONPsB1dVSLW6X/wqLJU8EJ9Sz3zXEmeHvhDjc3ETi09q4
gO8eNcycMIzwB9L1K+WTf44o104W2dFDcGK1Kk8qHW4xF9SZ6vBwAKI3Dae8Ju6r
ZAf27z5ZG75wdg75m1237OaNaFXRJyOySenxUEE8nngS8xB6JHzi/xh0FpYc6qhw
FPp1U/HhAOxtopJO3DCZn9n01E1YW3ugJ40bE1sISbZP16W42aYhINnAPdIEOzst
dxuc8PkObxCxztlf8uObQBt+FA3YcGDpYSSNBNoOMmzLKqKBa86oPPEq0/5OlgEj
tcs9o2PeEDm/R6pHQezmLlyJ7VeoueIvRQ5eO60FoUebaABt/cumE8EQNltg6GsF
EsdnpE4HZq1ihd0BkJYnGeeI8cdMuOIU4+G2YGotmJpQ9dFe9CA3gya5s3RtNcwz
EY3xhr576WZUilvF/TnWBleoCDo9y8OLsUa+zt15033GivhLl8lkN8HclR54Wmk4
7WyzuxjFQl3j92nQAgoUFL9JWK4K7VI4fgwUXQwT67v/yLpjpuogNwr7Bue11HyT
+/QUcG2ToRzM3rM8nkQRgaZe8rcBU7TYnzbZxpFjqmQL+28O4aIYnv2dLTJkD+bt
BmLzd8/t8N//NCvG40030JV1pfg4BeT0+Udrg4APWb5eZN/UV6pt4fVPuC0/uLKf
2Kvod7/ZY1AB+dmYNcbt6dqKrtgQS+3QxWoBXgG0g4EWMxhBY3KwBoNyBA38Vtoq
b50RomjbwxpPAul3ytSMm7NHMe50mld4OU7xs60Zzgmi94GamhBKOzU2QhzoFPJI
RqJYAPhTIfzrnZ4QBVEEbxIm02DA8Ookhz7LumBgsVyrZdfbQ8HDdbWgIMveLPDA
NgGShOr/BHtCJl647GQIygElgJ6IeWbTnxcIqg3B8LsmWHwg11qL/+xGHsMBD3Dn
QEIHpGPgU5FDpRF8m71C3KHuZyNa/3h96iuxT1F7T+TTTiyzp+TjUS9HpeS66qfd
0Ud0DY9Tf6lnI86CtDRZyF1PGt8eOcWPQYp5GRBrxZ6Gp6cZT4XLuSc+WJhLvF5O
Dz8WRiX2qtlQ2kJ4CuuuPiTf5WKbCAPU0OWFA/h0LI6Dk3MPh0bJG8OZvJdCTjQV
b5c/MVAWHhg/r7gJFWzw4RddaFI2bK408FrU+q0KhSzEfNhC6PG/7nsr0O7RseBe
vRJXJWrALwBx5AhmAjC3fexyW+Sy7Khs0j0KNg7K/W2+Yh3vZF1/nOd8MMrD+M/G
LnvjuJsyJM61ZnSBoLehWY0t4ist6uKYbT7EOXOlPgjLkJ3Ab2b1OKcxxNvUltLC
1QKTEMyTpCkTmP7oRyJCz4OoFj8lVkJCEggCnfjmRVpp90OZVATmuZoVRRf/hIP8
0BA/b6XFFGMCMRkj7nyxZveo2ohLHtGXmw47w3zk2H7KiOUB1vPmqDyIiiKbgTfz
KlcYX9LOhg3AO8eA41kN8+NMAcrZl1lWUcnQdByumQmXfniKpDAyM/+tVzgmXzD2
DeyEnrsGNjiHIP0GH/22KPPFxwSo2uRWsSskuA+l2WmvhDvyfh1lx+MMp7rNpCcl
XITL545QonBLM18Opw/3+2TeGiyXzO67fxZKjz9u173hGNh3IcGIwHk3N2tIvkgR
w4JrwpbJfsNPtRsnxOUq3wOt1YTiG3LLldXLT2kxsHL9+Qna7Bi++GKYX2kqgU7K
joGUNxVjA2QBQfK8KJR5kZ5O3dPGFMnF5gEFrQX3tKI9o5pCNzJFViLZHnFxVAef
wrfZ0iFOnKCXZ1AAo7fWBatC9/aQqw2ndoJeBNdGHP5iOtuM4CZorgzBmLvW6JK6
+E+BnXtQyYiXEsG/LSC6+dpZs+0VLIcorqKJZEX4vE43fY72+BY1NOA/a91TF+eH
FHJxXnxBUvPVIKj5jyPH+KfLHVcGjJ0Y3YAX/jv2j8D3RpHZFgZLih+CCd02N11Y
lch8BX2bqFtK98xFqf345eYxBhCVlS5YVI5YN5dqSwl4EP/P0flbtp3yvE1ZWHTh
K3iw2LXyIyGOUPzrVrXGPby/MIdGZPQd1VdZUxry66XUYZMG8zK7R8sO7EFZcHoT
h9sgn22UuNy3ZzzgYvXvX36Ytnp0incVhmA9B522IMAATCHBUfTD+5DCsNEkx2E1
TMB5L2engFAjfhXXOW5N8H1ECND3ynjnlkiuWTuyOdI7pqeLDlM7VIHlZ+1zT4b0
ZWGoaqtobch7x1vEcuolmXSPqXLpm4eYJadSH7oPEWOVccPy3+5i9ACGM7oXUc+v
iymaZ2QhzYMUOYiv0SgB/FackGjCx4/3NVJcqLTPAFf8L5uiFQs/r+UIDvAZH2Gz
mLF5DUACnLkZ3byDnhjrI+RAvbV482ij9wJliYypHcPNBu60wsp1Ezz8xD+36ght
jW4A/zhk4BOQxnMBUPprOIyhdDSRtGKuWd4u7SiZmm7vgTBy9HR6SwddrruSyorR
OoW0MaEJWXn4ViBY3i25JlmHTsOIUh9BzbTV/Mp8DDtZnASgrvQUMLpl7mw0tk3k
sZb4g7ep5aYHd8VQd/9uwFlGV7PJHKd8FOlyuusMZsg2d+SuW1MiSotvwaf1H9Yf
NF8GzTnvZhTOdDaJ/B6sN6sTMVyI5NBIsY+vVumUy2awqBkxpfWb7lna0AzBQsHn
6+vzcIydN3Iti+ICjJnxSSdTetWmtgzv7lhiNZtG9XJnFiWC5HaL/GsQsRLcxnlF
5HNJ7iLeZNYdaFYDt25Sr9qED2qyAvVQvDhjMgUdSKtOoBzTTyTzkD/HHXbh/Hkh
IqzUXwcb9axW9DpwsqDEIQtj0wWUixFzK2OiAXa9bktlVaBERHDSB+rXTLT6Pas+
qSeFFBIGimKGDWZEpsUy7LxCJBhskdzmR6XMthdDqcRcNGQPd+ZJySRm1hIhaDhp
izynn4HWeap5ZQezNXzh1x5a1xi/Q7832ZCIsq+YwQIyGHSaIyGC9zI3i9CRf/2z
AaypLJr+Wo1V9u5eHEq/gqLReEh0cUDaAxRZg4lut/sWy6lRH0dveEXOd+MDzYDg
A8gITRRpTkwaZzze39sHJHzFFT0mpw76XSoiWAwy79ZYUB6mULo/ZPfnN2ucD3Xo
QHprvpI8M/8gJ7r9aLRiCo0YdE/5khBzSYqsooUpdDpMIMRjBch6w7hDk02fE9DC
IzotOIK1xET0v+62kXHFsYgIfPLj4XLudfp3C6Yox+ep27DLOS4LQDMxNYU73HrE
jcpVLKIdr+08OX0n2aRtAcQpvwNMo3BRVGqrMb9pUa7iV5RNX5PnF//9hzJlQARq
Ci3odAY6RM1+Zv7ZaCvAwE+QiVDVAsWHA+8nJ2XK/yoSneSskrRyotS+HKPBoXyt
xkg9yhzMRXyV5lTO0Ny9x/SlYweGLo3gpTWRwKKolcbpWcaWp9BnSSMfENDic3Gk
myN+Unv5Ecb1J9kTACdsJtvfYU+zSbFaY/4SgVyCYb3L+oE8aNkRQcbhpYDXqjUP
fxlwo1RPVKRDbsExlFFPFxSxoc+J/SJ+HBSGJeejJdUwLLyNC0q9vW5wrc7DheqK
xbeEcn6BzbRfwXo/l4sE+FUwT2V/Dqf/h4ztWl2Ld6jzYZYr1ciFDqU1KckMyVhq
na4cZfNAOtP1ipoNG64Fpsh1vNdwcVaX/O9GLOM/wlfgcS+CMqK7UTDF6poQ5qmj
Wlerw+muZGiODBWOVGTovxCuKM4sYX58uGiCyteVq+AeegA4J4HYxcqg/nc6s3Ly
7SaWwQPvgPjKd2QN9DKFTwlrwmHt/+llHKPdLoII0uCeCnpLIEr16o2smcRMFspg
98Amq/39mF3P+U3k0NYFiXqVgiWnVxwWkxYWSIZlEkSb+ncAP4SHKms62kukSgXT
dT4ehMx+3kIfD++c88X1ZOLBFREbKZhBdxkSs6mNRSN5CXWEFbYu3eyrU6uY5Rw8
kpI/WSJRd/HZZXAhQ6Bi21rdr1Pt7eAY/K2tj36Usx0xgvdYukU4cCWVrkJPSM6a
Jasinu/84PZ7W8ame2EkuUP+1dygj2iH4HnAO6SIk0Nq9klrdc4rabNSByk5b/vr
bzOuSJMcGz3rj1AbkW3TK9CV+qm7o78NBGxcB6j4YoWle5qtCvKNf1iv2VgvQ0SC
ArM+GPKh7RvMsopwoCcXiI3/cqidFGqnwZVkIz4Lu6/w/tXdSMPO8YgzA9DL711/
604eQqoVtfVx0GQLmsz/Cnkjk6808U7p+xOASXTMzBhk4KSWaw5unru8U6TwjnDh
MCO9/ZZ6699OFia4n/loDoxOS/vdL2ePc0NCFZdwckOG+QpYPv9bq4W2Oh5x1gwS
o2o0fn5+gsToOcfwVlbEazgv1KnCrq/EAHbkrNRwUGj6+musSM7wznLii+rYEOf2
Rn2a2GFbWhp+SZ6YURyX9iqFhKTGWlPSXC2SOmTmz6L65fRkQURnD8WWFa+21AIu
qutLchYzVJNdqLFgENL2Xer9stKf79nAwhJnRNWPiYqh4+mSA3T965Kr2v0zVvYt
0pol1znpryJ4XjLr+qaRPiHOH8TqltYaI8N2jW6mrDKUcPwcyC9AyWy820UsomAQ
eMZpHat2jso23bqngNDFoOuLqV7zHCCNiYZJAl3sYwhCZO9hiCwk8DUM+Ureotnu
w4iDHEzKQzzoPYV59bWeMIqD7ZQAFhR6kxeCsX6HxQPiFjRFCIR+HrX5WjGEW0Ut
8HM908pQLry47bTjFRmdevFKSlUCl8w6AXUnHZS5voCvaoVlo3TujW9OcPunIZiJ
92yIMqbKlZpimeHqD6efAB47uZB5xXqXw9drQqFYesAuzfi9sM6zrZ8lE2UWPphv
sSnmDa5Y7YGOEWi7/HKIjVY6cqYB6TpRuchhmF+OLSI5i8VUUpg6dpBWIdkE8t3Q
Otv9C6CFnawdzz2vhl6+XJdrM+rnbWQj4VF3PHppn8PGvWIDTjnS/jpaUbD4ujjq
el7fMq1PmDEST6pkdxiPZzN2JJ8JnO7IWtY4pgBHLy/HVpKnfOvTvXNYr2XEUWQv
tgQGR5pv60tr1qhlwtsVr69JLEmqNNW3atf0JJUfw8GcHao4GJrfQT6kV2TyBDrw
YS2jVx6lTKqVqh876ARDbVSrex+qY8jUSQAQ8zr/EnJ0Hgm/m7EX3J9du+lGy/Vf
oaxiud4umMj6xbJAGZafB+8cB8++Vrk+1+tD4xQVX59wtudlPsThDd+VJSI7azwZ
7Wj+me4+gB1fj4kMBQ2prDnNV2ZMz/lYzRIcHlcdt2QZjH7dYd5g2c9bFnSQZtZq
Iz7tFTWYWBGxp5LVIqvJeCOEeOfs2ylOmGjiv7eJjpfll2LqdPbNS6S+cIJBczb/
4sRwr5OctWPyl2rz7yK4h+ybIeWPFZ5qiOYCwciNhjwc26MAu527edsdTycGxBjX
Ldh/3oHPrShz1oLGefCayVpPbt27PEJL1oyjJKh1Q35L61WXK7lUHiQZlAsH9PQw
itHWG/aiHjPWkL1GCtU1GGWsRJcRVki2mNuBhjF5V9SX570mwHuEoo53ReTZ+y+N
RXruDx/w+j9Btn7ag+wn4A3qe8hrfgkcXKD4GjSmvXnVXglAOEDKYohmCNjofAQm
6vrsmrqwDSJwBFZJI2t09FmcO1WGoQbp7+v/mRWTXif4dqDUQ2pLchs0xkojCTvr
IpuSleT9IfXWHJAzGD9maOd/wo1Mi+haD3P9WBul1XB+m4XhtA1PhobPpd6f+2Or
GCFa7zhYDGboJALIvk/p71tKQxk9YM9UJIIXgkPlnwWl34P2PxaoKgORJBS+M04g
TU/WbWzM7eFBaak5RnAEbZWXsUP2/l9QSLUYLHpr+JfdryXp+8Luz6wwaVrOlAgO
cGA0htM99pZBisTjPEwd7OMdD28MxTjQ9Uo5o18EZYLiFu5kz9ldENF+Uxl2Dnu2
Cn6k01oFmi19QnaQiThOHvOpjUgMGVypkLxCA1N5kRtXbJiZWsvZUDWOSuYsdrZJ
hRiXFqWeXPwLM7X6yygWwsm3yzkD5/WbWks2zZLhmvMjPHC9FaEBapHlzwfVjeix
e2saEogdayq44PEL6O8wGAS8vgi6DtFEfQTUPA7vDYUpnEKwYeBtEkXfsQSCFhXh
2TFCBdneRpd7uvhQEhyeYT+PnXQgpBstgqnSvXoxZxWVxG2nF911dVSDtENhoqF+
urG1P32Gd3UOWcirSuac6MD8I4uoE9WK+II8psl+Y5yP1qyMmEHD/OiU54RQuZnV
4KAU9bBo4RyZs1VM1TX6s1xWrWy7CmJ23ftznhi8e02VKX3bQWbsqea6n6W/RJTE
8DuOY8Oti98LSAzLrhMZa3NpGw1iWP0M89TgjMwPvj1gHBs78wBEvWaFeH5x1OVw
8VLRrFn/OStu9+JXd0M9WBMrtCNNPJaBG3vTUUMtRcUBLHbj60j468amR8VXYfp8
PYAHn1vMMTZk7Ca9mxYIM2ZIIKxpO1sk0MJCmRsRgBfEsujQUqjSZGtM6BA6GVgJ
+bzFUhcyL5P8nKltMkU9fpn3vKe+2LMCriTPnd9Zyh2TgC3TS54zRADlxJGnezgT
SNUCXPzP0n2NKpswuvodNJwIKeuqCIPx+jvMdxCWRhErawTxS9kvElReDIfforAv
J0pcmGdg/zvVqCgFCsoCGTPSmLHIuxDMxv0jP4vgTHeYgv6mCpcYkQWCbXLGYRSK
76gBdhep07Nj3PLhMKurJvXNwY9tkNdkRkxR5ZEkiyrrId/5/f/Fun/sPyQxkAuM
A9Y0S3qvFeZpeQEjUkFLusiGAVbJEHLUPRrHQgHSY9cdZ8sZ7/bo2VjWXfWNRwzt
U7QMtIaijK1ewJ3+z9QF2F07EfkU9sEPy9D3Wuf5A2Q7w3+fDP7Ob3VlnugymhRz
7Ac3eSr1qE8DFUZeVzaG+7HiWjlv01G3G0OBtY6GKW/CRePaRwhqiE4UCnKBGAcD
n7ZezxFORlxaGqMCg92p5wGsPiayWGH/J3T0zZlXYVFMRK9uZdijJtMbZpOT2lJy
lAyqQwef+8EwOnZN04zAR49/j9tihWFeMOdscHB3qkP49cup9hYllnMg5b4XOKM4
smjpwzok3tnjitTcCsR8/h0jtDu67xgSGYN1j9pMilGhfPkmMhxDWErwzQCrAUsq
QtkHolpVQwRjChppe8KbFk5t12imsb9VGejFJUoir2fBIOHx3fzxVNYlLmbTFaTs
jjrNH06HEMWSaIA49sexDEKI1UJxZWy43is0mASOLEHw2ayaOfG2y9yUoOO9Wvr2
29FKDv7XJctBWX6UBAxOuTZINGOdhvufBYEkdhl2Uz5aS4xp6WuKeF12xvih6PXC
gT626NoT7HadTaMhe/frGrpgnLzkzQtpdfprHI2Eu/FKoHaYFI7AvqM1UuWKUqNo
mdZTlmgI22e+GqXaoJNpyx+z6wXLf1Ctu9aqn6j8rXghyZLisqnRmwOjp4NuM9L+
d60wHAcul1F/g07FuUc0J0GdyYVXXIOD5DC5h2m/UYxCEEc2E1vAUyfGjNl+I4GI
o0uu3D0OLKyWx8NhrbC+SgPgz2c0TsXDAY6Dy8ASkYjwY7T6gvdpghz/X4qRkJ+N
d8ozdRg5g5R+TxGynOYlgYxMypVPyJELiNtb3EZ2S3TtVnEX14UTHeyqbQxZbiZm
g+knuJ+ajOYkSRZCESboYPJTC4XWW4b8u0P+06vBeyXtRv0hNLfj9coLVBjsGg3y
Ig1WIrStBjn1HGRndIwWo3sYPwkrDmYyG/qs7TsbUK2yzXOSNYem2M6evFhuHbwn
h57rJFwAIfs3fqZ/TRHUZRRZBTZ+L0a2CueDn5TBTE5O0AqweHn7RdOAXNgzLJ5i
3M2mb4BhxdzjhbXXNo4XVj8v16PfxZ9Bgm7tpJDVZjqV0PK//yJRzq/2AR+S8oTO
7eHc1QgpH08l3EVfZ8y5wj/Hz0O3uhlVtyVDFm875JEykuYQVQqe8Rr+yWWca74a
0lJtPmW8/5sEsGj8AnxgfXrr2v7jiZZut/cjpL6P7ifoFIwdVCo+n5K3tdKpMm5A
MX4b3mD2cxxDEbnaRDYF9qjUBJmAmJMcZaa2u2nplXz799zSblRaTk2Y8wjbzTSS
Gl71sHAGJeNXb2zL2Eataq83jP8Zc8r0ia1mgm05vS+nVgbI+wYUSSHyYuLBB3SC
TpwoCv6rb2GDEOURFDmpcqCdJ299tCbgOsXHTuD+lI+xtQ++MtZPGbDFuAXaUdpS
2Sp4sYh7E16xSxXJTTXBorvT5FPzC+5qst3O/O2WtmpBrb4eSS5XuNkcZQKEW2ZM
J0Ir3gUHO4YarDxgE5v5vsHVTWsr9TVykge9KVG7ddF7bdMUZHIlrB0HXtvJA9OB
yl6LXLleYP8SC5Vsdcn1UzZA3jhv+8HYhAW6atHw4eEbqs94jwU9RBb+dT8q8f+Y
bpSEskhLHi+UOqqm/OwQQSm8pD0YpD1XxQf7CuOBl36GF4oaea1we9OJ1VJZ5X/l
fsjeQk6cVBlrGhGoobeNr5eeuspWbwcdqPPEnmIrXFEzDaJsqY37ChCifQR/D/Fz
bRYptB+RjErZD/+Xe8zFgQEnVTiy6JGarD6pi2UcCSfBLgjcyt4Zh8XHJec0Yus3
QsXHoOGkxxZDFPArBaWRdHthgnfIyqtXRxGb6St5bb8NpVqhOIVZ0EAlEaH92hT2
h1TaJ7IXS4QsBnXkBtGAExGrS+PrSXH8k9BVrtaEj1d0f4Yky2pufR1MwkSnL+ja
/W9zKjeU8llg9xDWhGfHi3hGBL4za/EYNUmHPw/5wQOWkv4970TQu1rWs6LB9C2J
sXQujP1rjZ0qWHigRTDs/SLxbdZxXliWk+iTQKCHSo2qWhb6P1zVuSuyMhOYHJjh
YbE3gkc7lFOcqCx/Q2oGcsCMkn8Sd8ED2IuAcmBtKaEtm7V5z9RvWYA8d2Q6dIWl
7C26cWMtHX9IhvkloPbiR2ydxloS8NrHz+7aYyBnhj6SDFJJlcg+Dw032ycy+tkD
AdixG5SoXIYXluuPyciDhlnP1b7xCAnDx1J0iQq+e5TV4KcY8W86BeuHbRREWk0S
0ZsQDzcEtA7Q7EjiptCJxDxL4D5uqqA+yt0f30pizy+xO6JtkZKCQj7js2owCifl
cNjDnNKlTv/vf1HrzZj/U5DLASaYR0BenfsAl+3D6z/dFaFU61zQLi5r4O9gXMb/
9ayHb2/khjqwkcTo1oDjVMvIo5WhFwOotpJLa/3vkD8Z4nA5nFIOATNdyUFI12j0
3SbKYkOkNapcn7OZwnKTeRxlPcx53T5jjgcHcHmSTN7YKYHMSnu7fzmNbnPkATmZ
hmMhewd9GKfb9ed1SueF6L7sH88OPa9l8CktkdZLx0nl2MylD1xx7UJf0C+bIq2h
yEypleiHyDO3iQllOagxHkiBsUwl2YVx6k1jtQkWUc9Fzw1RonGo3Wd5ylJDl4eX
RJ4SR25e6ZA5TV1WxnRzs3Ti0jeu1e7jD9XeYN2+LclfokQMn++SjGBURxUQBQsQ
Pv4ZFvIuOw/3NKAzNaWXYAnhvfvgwCNiBpLyJBIvkT4DrUFIqLAZnm/xLvYSn0l4
G9FSn6d8LNNNTAmZ7oRsUktwFP3fXgE/9CeZjzarsAjJrKg6gWJl/xDJK67Ejaat
scy1anrDixQie+GWB7ZgWRmW3FyRMUuQe9K4N0x5GQm3+8O7kcFfa+heZrlL3V3v
liVodkJrQRFthd7JA631em5UWmYi4WA0ikaCgTdk09vrA9NfYYclOYyGu2fQhsgd
lAPrN+aHzYsxHBfFZ9kvPf5F8hZnjWgQLHkiTsJtXrAhYXhu1z1reKwHlI1FiF+a
3iYNjHqsHfBL4s0dejP8Itjs9/O4UovVZ9YQCq8xDFTQvFPrIPgwiPmsL8py6bP9
yx6z74ys5lns/s0BI1Mh+wI4JzP4wCxZGbkiZ50YUVKBdVKmg5Np7A8coHDctYCQ
vaRce3UWWsAF63MwPSsz+utR+iabIwcbmXiO/Exc71DFlzsdylj6UA6Vb7I3L9cU
JyhmCg+KnEAUg0dG6+CBLlRRo1kRmzeJh4x7yvosIkgLeTaGUMNH0uskR1ViSG9N
sWY9BhQ74Qs39VyEQKMtcw4doN3mKc7+TXasL3lTdLdUM90X6y+wW5byu9WYPpZO
ShrEsgsXQCWL4i9pL+t+uaNcWaP5H83aV6rrewA0lSBNV8+6ezW2PdnZ0RxxtFrE
2EZ6mnVF9+0A4/nLg5m0EIFtpr7/psM3gmmQ3JvSQ0N1zQXXcPsezgI39wDlM7sw
HxHYxZF/YKpEnOTBAu1Pd6WUhWouhz6VEuUdRSL14G29abXIgmYQuKWHTrOHuUtF
U0LO4HCcdPlGtIfooSF17WBc+WslhtKKkxByidH5VGZhpIM78l55jtb94o5kNjTN
mv3ybSbnTkRtJHUUqEO8Pk+K+n2/FjSbKASFeUQbJ4wdHJ+v5mRJHoNEeHIqZIzg
VnEjZOPRw6PvJGujKA9m7glvREItLLM6qKr2Lymhf1tfz+iNEKvNZVW3OqWWiGsq
df2zpMXfq7wiW0xXvNNr8+5MPp16ZekNMGdP/HFU8Kr5Ls+SlVvmKFfRidSDGbvC
mm1LX3bO7eAfC0OL0NSu6iVWvoN8Qzlf3z9joSIxWNZojQO0BwNHPSMUFQLc5ZSu
oCTA68hjsrJMlBwfPc+Z84d082Sybd5vJs+DRIgUGqUWoDw4JtbFzxojIRicqJw3
dKO228gePm5j+4Te9eqJGEfapmrQt7WVgLX+AJQ0/OVr5mGTK0FVuGbJH1sz83qX
jiqebRZ4g1ev4YrCZhS4hMQoUyjoW7shWGj9cjq1yrQwsIiEXaUrGdpavvfLvgMT
3mIA+ZnhtGXtZ/9WWoeulCHajN2yDhqifmbBNKFhkkrXkQvfTERKRobAb+3vbI/s
v2+ZbTwWCjFxvytEwcXON6Se+cEG36gVD/8Txoru+J535Pb0cjisbbmZZ7fFu96n
v5vRRhV/hdCoOI8cO36DtrWHbvL8mg9q9ycbw7I2sToxE5+HaKsiS7DiQ7sEJa5k
6kFufHVBUCE5A41z9s8kQfBt8hChcqLmDaYwUqkPdzBWINHUUh7rOtiz281VobPW
gHymRj1v/76OO9QnJZi5qFw3VVMZE3cT2PPmGyo0HKTbOj8fCwh59M+UK+StlBqZ
pz9eNbAaOHpFJHBmD2DS0HL+r7nZeS8m+1uTdZOVjzxjqWbcqSzqORmgbUY7noUH
NzJOZ82/GQxtFXuNlskwsn36NCwgcgkrKfXbqpjoUnml/MzUlwOcqhLbJ2n/MFr9
O8TBjZk7l1kAEojN6gXEIN6++vliptcqW2Ts99j7+rsMiRhA6UF5ysg7j6KJ4Lqs
H3SuCBsW6Up/oVXPWO/J91kxxQIc47iLMye1im8hyBbtoliqYyOe1yd12CdQuZ0r
FXaXHdFNZKc/UorLHUgHUpmYBBxinoNxy8QGzfkS2IO0cOul2phUqbN1ACoqVaMs
dgig51P47PQstywczj4hlT/ltbnRgpuOZ713aqLnkF9Ku1YxXEK2SXIIvxbZGac8
avOxgv5O9c89QWxSjIcAKAFcWQpN08ra+/ENhFxtGNn2PQfNMKaMqMn4qjmvqJu/
YiqTDR2+aHziM0e5Y0Blr+fBrtuWzfB7R1tfQeQ6iBatB4V7uRYnb/Q4cCfojNRX
IqvHblyhA1v37f1+6tp5ZsoWubCWzceKBFtOyu/Hkji0oakDib3Bs3cYMTUZ6krv
tAzvtEGro2DnlKdy1+6itIOuszvRMvHf8WBZ1Shtq06VsFEx9DyYDXSMT+J4F5XF
cDYn8xwTvuvkdC8gK+EWzHFI2pRB882B9oDK2QfTHRqKLzxtJgt0s8+UNZO46Hw5
oH2QbjKs+D9OJ/rjGoMuBm6kFs6DYbRKh3vGTgr3Ed2TQofh+dVDl7S7kCApi3Xi
KFaDhdcSpdB7BG2ZPpuulLCXAT1ae0d2QLmzzSNchA6o0IMyH0gstMMXbna7cmqO
2yCf+WakNiPU4/s0zNsYK5V4+qxdkFd4/pYHfhmbd82XkuJ3w2ivQCJTc16BClQn
W4/RV9Bvr5bGhKyPg7E0rOKCmXtOG3jdFGsWNnHsdDQ95OtQj218zp2QwQC7Dsx5
ltTVAIeHlkQBAo253TvxQ41xnkzjuv+eh8NMivrvneRi4Q7deJUGmGXzCcxxweAP
veXFhJmm3+K5wxicwKelIfOo849f9r3CuIy39rZ8FZl/tM8zEFc56EkC8qhe6h+Y
clXLfP2+cFmsB00iO2e3YWxLNrjUdif/Xiu76m9/jWQnZz861gymtWWD0u6OhOL/
tRM4gxWW6Ylvwlxmf9EKG2YuYdV4xb7QWUnJ6pNojvZpixruc7V2++gDocE9r5Dz
pHxAuxj5K2IBrDY07geWeYk/SQ7t3ZscQq/aT5k7A0+n/sViucHiVmLg175WFYaG
sducXpPox3zCEQJq47UZCfkk9TSK3hsHz1uJvx1VmsV252/dwUKSJ5DaWmr/3SlP
3hg/ffjV+q5ffK03lovEV/rlcN4xsYOP94kCgmp65FjwFY2NmPls0amiqfvZavdt
BGbaH1IZdHvhGMrBnWeTuwbrTFcxPV8LblguKY8s+DKZ/9D8t/HCzt3/d4NKiRHc
+Y2UMHxF0KlS34ZWlNWrbvNgiIODHcb9KuSjtTaMmBuTQwP5Ta2FJ0XNX/o1QFkn
8deciI+HKHj3go32mvLNYRAgy34y9P8rR/+LmH3EG5938k6AOFoY54kdg9BdIPlV
70lEPk99mlf70rnjcT9qmN16CEbWlh+BU77FDHJctd2VFI8GV/fsCOtpsg6CHIpL
yv4dMYfd/wlrgZYcrYNZ/IQLUdfvFWNjhEFNYzo7r54nsELmiE1855UpfCEpb1CZ
XQpfz4/pOlwoy9ZjXl8ZO4VG+bSL92qpkyLIss1idexWrgL0znvRerMMW1k201XF
ea30KEXI2gUtKAo9uQvNHzOFCWhhK4F9KVLLYAF91c1HHrMsOUuGI2PzQsep4Br8
isu/AveGvcfcgFL3FCfhZ8c2GYWlA1owmCinSpK3yTw8vvTKh0D8ZhJuo2IunFC7
v0WRe33Sfr8GY6c829OLvtiaasaxPc2g/fllPRPrjoDF6oaILuIefZ9lQZS6JDZq
IrqFwV1scheJ5K+w/bUxb26wsP7zM+bxfgl3lR1rNtaNC3zyjXTRfEI2ju1NvH1T
qpVk/Ug11Rt/px6zJhJyObyTIJZXvXIWs0AgTt671W73CR997gPemflfRy5jK0YJ
S7yGbLhdlMylIrf6+1A+zG7kriaTarZb55UwYLp1WwlFTjBlDKmxsgO4Jc2q7tYv
c7y8UYiWPLQY5Br14TBUxp4GLJw7Vbt/EFh72re5M4HsQRU7PNFTApE34zo66AL6
8Nxvz2BDSRDdOVUWlPialdd563fJTMhPimBQroAUtGD48lX5THRN+DjjiDhJRJxu
SKqHgzCAhcVDB6d4LZZz5/2esdLDG19l+da/Y/oc7pZIuPh/H5PFtA5zDL4MyVTv
+cVcD8X+hHE5PZhCeDY+CdQYnPrva0/V+IcOphs2HmVyFQxRi6qo63qaZiCGD6Zl
eIgVbQGeutYKcQ3VvvuEUeGFIYLMPMsbmnqtlLFxAUBtQOtrJ2Zsy4OZC3bDJR/a
iKudl426htm9O/T2mYreW2IfmFHf36bh9I6MThjq0rBXLIvT8yCBcmchIWBN+Bu7
lscmNJjliIvHB8npVFsuGG8jgQzKBPgcfI8pyOJfxcYTFl4A30pz6QljZ8SWpdsB
strrSYPYOz+SK8xJxcds2ESu8JpToe+VQDE0pu/ycy3K/KmcAXyv7UN5DIIAy+7f
a1730vqCJDQj97gBRGzQ4DL6WIKsH6wtyG8xeKOPPhY+UgWlIPa0r0bkumU2WvO/
46w7Lc6dmvydk7rAcXRutw3HvyqL1hz+gAJlNHoGCOjP6YKbpl1lX11S/mdG8CcJ
PR4+MonLhcBONR5wQzrx1A2aMl13D55tcQxj9SyOE65cvlkyARMqPwuwcbtKYu9b
85gEu4JS0pRma2aYuATTK3pDadNpeQPmET3p92Q4zXf+814dOtZsz4P1tBy8qqCb
yYQfPBQlxBpbSzP2SWOb5ht3sDgebyDLofWpczu5VUMTG6u2UIdt5+ABID9k+oEb
kqbFrXBvuRk+EAlUtIWfJbRuDzapo4+uK3rZup+hSQiZTVpsWErOFEIJ1GF8+OZn
5KRklawyWv7XJOxGzVvSrXFKQ9JXM27piM3KSc0eFt+Nn8i2QmXuepLOBFJDoYXV
i4Nq2deRuCJVG5TsaSoaHdDC/Ds/O3Cha7E/m6ByuB/bK1htPrxwu9ZskbLJajtC
Xkpgqa2zBv81ioDllPXONKnuOP9QLo7TCHfd/n1jXnTlhx5gZO3MeGKRe9HeUD1J
BUFTmnh2nj+5V1IY5Mt7+51CMKeHbL1xFenKw7NB/GC4GLXlGxSa09St2KI5eL5z
Ljct41z9Vq8TneeLbRHSZqMGnLcZcWgal1Ye7tpbG2WE2dzqpbAGoI0FzJsE58bG
J0fS2XAc5DTnNtrptTXpgd3/aW7OvT9l5IboKLiticVNkYC7Oq4TFVwnowP/s5lK
mwD0SWHVl4zC6pHT4wNSlSnNWAQy+7pDJNe2kWBAj3M9AukRcyDCXgVvj99C3InB
m9AvFh/LTkANcBmnwQzKCx8IbGXv3ieBx6RLo/b6dLxBI+P1DM5O4/uYu4IQCgZf
MjjkNtu4sgT7YRTz3Q4kbtk1L2hr5vWBINhnYHLRVnk8SBZN6SdQBBiYfUuFTDux
Fdw3NKhFGG98XF/fNHb+36/a929eVTleotbgV9FlEMlNrie5nhztYQ5FxPt6hChO
sRYidwHS3KwS1yEVDteNPAp0F+7wcZuYPFWzdnfufujvkNgzFxoIAWfDPTJT/nqt
BlDLvlwlwwMxAzetkapJuOZg07SqTn0yWZY4KD0SzhCKCMn/tDGs+JxIFKgsN/Mg
8ULEvGHwGMvAbVueiH8wbZ+c8JPEpAO50ryGzibAaGLo6mCgElWxBPUf2z9Y8vHf
JWmIekU/TLAyWW8VcLbm973GZKsUkQ688hEjjjwfZoosAKMrVx2uStvZKNLeTOyH
LfUdnH9HoUactA+5itOsSAvJ3Pr3Kal7apv2ZlebnVxZDwL2ZdAhaLDtZ11WzZcZ
wdY2zZjN+lvSBnYcbwK22ubXqyfoPCuWiG5AYpi23C+ksttqt6y64/myhMRmN1h3
bXZw/EPAMDTGYvIZ+LSAA8CnYfdVxu3fgVpubs1f9/XKKCMV+ztKAvPCp/YqwVgR
CHgsXAIB49N50LnXKnm0J3HelDd6CBhStCaLuQwpjuqbVRGPcybYGTSWS+sALtyl
PbUqbYwEMlW1/zp06qKvPMf2NB+kCgFQZPPjohT0iJ3gtvxAvD/agLwAwcStNCoK
d+3WHRNt4JT5cW4CRbdZ5VLNxGeStgPuuI9D6IVyzEBxc1DUShNfxX01VO1OgzEF
kQBkeL6NHCICJRJOb4pOVrm9xoek7UiTMk78u1svWT0/AryGmeuJQdxCUzsGdTja
7Rffdpuek7AsVzWyhmQ1klVIxwKN8YTEfSUamnUoa8X2ONxUEEwZVkBBR7GOaNBG
MScKybnofV4+IqORggpix21ouDAP5Jb3a6DK77HPGcSDlWC+bdzW4AcccvLeGc6d
uV+kpeHlWBB7pQOnxqroZM+6YPGAvMIFZxPrhwuof2+2ZRr/8tFaQVfG49CvElQB
jlN0bMp/ZxmbAJ5oKNbKdEUwrXTFniCA/1kRxSrNLptywqf7rudXxff1lcQ6A1Ss
n+i3/0OD3WnRflaVWZZ2f6L+0UW49O1Z1eRG4R7Wny1hyhnYnmqDnYNsa/fiwzsy
OXMYaVyralYyLji5BApuEvcKyCYHsZuszdxk27BU5WbpJCTSeHjufIaqFEdNajRu
muWcX8kUnPk4yKU+dtOAaqJS4xtxkCjNOZphQWx27iatumnZLIztK74CyYZuB1IL
th/65MN0XbUNAYTovBseGXwMG3E46MAXJfTg7UqYfbsVJu2N8xIrpYcujZICA1Rq
V3B++55tADYWen3ADlva4TqqmnGR4PCSfvg2uAKu9E3MjrRehnbnDKkBAqnnVTlq
R498EnYIHlL66xh/xJi6I1wFpl26Vv59yAtaaTrMQZbtB3m3AFsYb2ftVZJgRazM
5TcpO4M3bL8MRBtH8Ac978dbFs70dRuBbuVcEbF+NXFMzBQOqicbIErJmxPDQHbA
T79JZ6v9ZUplfD+HnZHzwpBMl18bVnPVgfTGvCnj1TxgnY5FhYtlD8v6/C9CwWm/
57QBoQEwaW7D0NYp8z5gqWA0JvB0LtMdcWADibSoaAvVpRpzxeQpy++d6mRYzC9k
t/vc9mRUdtcrPOq723/VwyhrxU3Z6YDEBt88n4XWdkamarAPoOwwWHgE4REVvFcd
z8o3/4mlqaCMgwWKryWnev01BXK3B0peU1NDRFtACwia7u76LTkmAk3qkLCBuKVM
3kKZ8DV3ZA5IPK2VdxE0Er5ec1RbmIf1ytsB8MGkPtmQXmzGfXEVtX/Nv0+YDV5G
bY6zcki55bWruopG9tIDHgdiOVhhKmb+GMRHSYL/h5rfrnSs9Z3r512uhzkDmHFZ
I0cAGoyVkPN7uOjdavkTbZ4Xx65VzP298p3Ejr0beIJWTPKIoErdc6LyzNMkYH5y
KTJoHm0gUr4cAKUS51v3jC5ghQvi/hrsc9O2jBlc1fPh1dUNQqL3iqR7v9jzV6/j
bepCxUOcOy669kRyvFz4DXzCio5PeEXsdfHNwLWl1YfcON4W2xhC5dQibWyzUHa7
qoCOKflaqbyP3sK4PVGw+ePKtCohcyy95tBEyyXUMDIUIicZEpnwMQ1N0AUkFzFj
uF2hgCCOUwYlJYfNVq6AJlMRuNF8iZAWUVyHzRHkP7TmY3GxFcCvueF67+coJs2g
aNSV5obmcqtrp4VQ8gDDCpbIv2RBe6IUC9yyRltwVCTrf7tzKB/LSTxW63xujwrS
ekpBxkO9sxplnuQ+CVEaqc4p7Wm4hnamDqq5nFUabFjkKH36cuOR3YvSR1IGVlEi
Smjxp6H6ituFTb9Yw/JoreBbewbE56kh5VScb8kN938OMuWSWrnL822Q2440JEXV
wma1ZTQn0mULarRlMUWb6hPCFqqZUpsaJ5WV4FeVvrl+Eou4b3De2G26tHzXhs1V
hqpHa7ykX1Lmo2cNnwslTXC1V4apqmTNAu75ALRHiZNQbnmbwnI+eeBnr4YT9T7W
0XEvGlOYcHbp+TK2PFdoOo1nt5ZznDa4aLxLocwhz8uJ24A9P+LictJoGzdeoM29
fJPZLdL1iHUxjjXDTpJyN6pPryZQzMKKxvzx9tKsAreNc0quUPS95G6UqnLl4yfI
RNRLWU1eCWjthRbuYNwZuxqhu3LwhamVWbSf5zyfTL3g7OqcgdL3JnfEa6v8KCoA
spR3pdM9MEuZ7pGYWXKQlfhdStTFadUHKEekbEfWyo8K01xPDPz13kcj0p0i4qcC
6RDw5OwsYEoOWIPnU2tS51/xP0m70KyJ2rLxqhUi6aNDNSGV7aY9C/UlAyX+mqpV
Ew/gp7wnDAB/SBFs0w97TJ5ovfLtJp+qsygGAMzeTIDfMBLZGftvURQqXcNV6qe4
LvcktaJyZR6veqC0vMJESbZMACPdkMhgtSrUZ6R/1sNs5LPEYTKo0UK0SIGD4mfZ
skOfH0Tcd3Q5bWLFVN+GRS9+qEZgYKYg+r9K1V7QDb7qfn7G0tzbLKBiVuZxLQF+
WFDunzlRyzMrXat0eK6OXpxPWJ96nex809j0ertpZnDOkkbxwOpcIIA6K+vEwGF5
123By/uT/BoE1bdZYSRQ2wF9BPTHAHlmZWhj30spyoE4DWmahqKZCjd+SnOB5/lT
l7xeghQwwHGLwX0qyj3cooxSwL/dRgWWloLq00tk9cD9RtEfznAFvPyGVlfBb8Un
6KxM0LDcrx7lqWGvERtS9tQfMURFEwT2WfYFmMQVZacXIZO1GSXm6v1SqVCh+Eml
rhm34S/EOxXlibxprx34OM6TBzzsl2OsFgPJag6VkBMcsZDjElFqjGnYkt3I4GTv
ijvkbv79VNbci/fBkwqsMAiuqLIVdyXVw5F/OITYPTn9iTQFS4psenjwXiYRf3mF
5JJ4564W7YRc24Lr0CJVfw4TrxiNRmmdBjm6BxS01Gcnpc8KsvkSMWxX/a3vk+4W
6nWCU2rLdM2ABQOFl5MfkUKRYVVEG/zmah6MWyAEDi3tXOuyhVC1AEf8yvGN18lO
jjq/b8qozQKEOP9KjznfwwdkGD5mIgWrZe1ywdzlaB6bMWeVC8zUHPNovJQ8w6xt
jTHxtUGa3jYmNQu4KllTyLND/Fgog8rmBHHBTYGK31i+096JhBGCau4IdIvec1Y0
Mb/eW1zs046VeYltx3Nb8ycxibxnN2b8EzEwhnOUvNmv6w8XDGsctsfbCuWIGESs
FZUDS5iCxqP7GflGeifipHfHHIc3RRm71vsuOPWBOQsQw/RzZn7j52Mc/N/cww+2
ePAY7zuy8ZqXKQWmEI6LbjJNRxSx7aFHnn4KXnRJVSy8yvAs+p74ZG5kTmxvT/+Z
hBPVd42klUbORM1bxpSATcGBY3V3tplo0UqGAhOxGEIHNIlf9puILys2y0zXaHO2
enmqcJ5bZIw2BVpU5SMqmZimRG0pJaXE2d7zfI8REyKWlJlwSKz9yXJoxdgdLb7f
lT0EQuRxk/0fsp5GkfHSCjpla+DsnCIEZ7ZhG+eGuoGm1/bHEfT58syJG9NKDFH4
zrglSZTAt8v4gOdabtfwUeaGR/yWuNdd1Ov1xKinNqra1R+qSeP/ZSO2ZLJ1euwg
RY9J67M2Jj1JbfwaEj25i5/l8uw9K0UCVBmDlmC5UR8D7KZ2tFmSnrAqYy8gkuqy
N6K1YcbXV71OSKY+9gfEtV3B4Ac9uuJwWt+jy1LN3Ggbk/4UMCyTI7e/ffgUPLwe
VegINWj3uh5pKNldOVBmKuwU6uVywbnPJbimYQxHbfZOCDzKOeXSaUFvYvF97t1W
kGgcbwXCvJjJnH+yoaJEJnzuSH3muOKTsUsVDdE46OCRbB3e88Yksb3dwDc+pOj4
8mOb/FryVJBDlrcttKoa7id4tEhCV3VgXiKkO2vqYPFQJlLWUYpM8WTpGTMmHp8S
F5Nn4hZL+PwEzeD36kI7hTcsjm5bW4U07ihKPzy+ifPF9qqW4x96BNcITCMpfpsg
MjdabM3NPUq+J5aeEohFK89Zc1XjhMQZP89yfBtbWV2j5anntCXmv2L3z9jVFpFr
8s9ivWxdwcQgc/j95xe7obt6cxh2Nb72VaprVzUibOhtcRUwXPB/NjmHNtpQXEQD
PqdlrOkYpoQKPfmRngKXfGYZgbVotHQF6kPoX7NEcxeP8oVrhtDDSl3g4RC2b//e
FZQVqqOLExxLvx4hAeeyJLzu9nsIkQzAZV2iUFxJtiuwlsP5AuRHDk52bw0jjRfj
vY1NpS73dqiJyGhqNSyw9AJapCpFE9AOh71C8gOWjsVAl73jbrZFLYCEorDcFPIl
zJOqfsM32RzA3ReaTzL09ymj60TNwS5nXe0ytTEMcJJ3BLpEAJ35QZxcml/qtQXu
bqCBcGKuADPk9ibsKPKUCoDJyVKH1DhIIPgOCPLzOD9x5WPEP0npxI+SIfjVv0zl
qxjwGo53jl4KmHsAhliORe3Ueq204hGvx9uwBxeuLMY0J9BCCq0NE5gFSf8wl4My
edjvcjPzSXqiUSz8uwURDo5c+nHaCpXeXsym3wE8xfYSmb0S5kjlSpIYgJnBPDDV
/VaeDMropmu3olaf521KowRZN+fBbFBEUq0Rt+nCW7ir8bA+ruVw/YndVwWvPt3T
4RQDHFI2LbWAWod5ERzlRz3bW3whRgW3Ezbh7MF09/IaoZQ4lK8eWyTDfmVrQsWq
L1w7zA+OtsOf11booDH2dXFMBJKqoksiUBs1P7I9CaoaOwplz1pHebdm2OB4NPMZ
klhAVON1W0FimoCsTyUps1ONtxkIhk/j1UoUodugpHbk5GtUEeWLAgPO/nw0QKC8
7ZLpTyllZwGQPyeS8hU1NjKxdl4QF2OoXl7Mpcy+h6Gt8ssco2/Djszxu3r/Ui4q
nPDAhY4apCxVV4hvS5gRi3gU+11YZnFWg5bT9tCyGs2qsOJWaLQaFhGHnlY4V5tI
eKS60lNS5foaTrreMKBlnbaLngs+0o5slNYX+3Vj24aUFaB7OIaIRY+BxxChTN2/
Ow7A3s0Q2MSoRGeY7p2ijO3KL/uzsFid/nTGZowWHtd2wPieqXxh7mmAd+A9Yy1t
Wsk3qoFU8fO4whM85L8wxwZJkvaRdlmMpWCrjtk8X59psm+lO+i8Dz95wd8NghWA
pqk/R6zGI3hGbjUKxVvTJOILvIYGBH65HsAerGDC4aDHGN2UBfuZxcUH1iV6mqyC
Q1Hb12H3YcL89iSoMvdFDG3f+Tz5NWiupoXx9KkoYo/iRLJWmc183Bc2qm+KcjTM
7G8IipqYhvPeFlcMhg2ttpH74Sm+bE/lGsgdaqpvjEdccxTk3PUx+fUZMH0gOG2f
FO8QykJIae4Kk41i2Jx3U6NDNU2gEIVjzVyqApOP/Q0uDXIP0OBVIdUNPXwUsTmM
qM8gm/XrfhD0Wo35FDdbLz51P8IWPWjbA9oFPY6IEwrw0yPogEDZsRO2qNRtvhsB
VJQb2Ay7tXdE+5WlLx9BtHESW49RUgeQs76bikPh6qyPiylhH48YwczWCazOsG4+
tNswIHVuvyI6vZzGloqh1cFORgZFiKfbO1zWRPriicQEvD8WoOIaRyb6IGUtzHaX
BMzXFVgL0ctCRNIsXAeLHuiqf6eVWssDhfbrGJYLOVQEYlG301UuX/PfJVVYM1We
nKvhqyQDqjmN7GR1nBXyLGA8GV2MLGnJTHrAVjJWFN66VOLJKredg9vLNc2Znm04
wU+EJ2E5Ra1TpgBXQwcnB7DYyBMzxYNT6T0bXOx3mFMmhm5AcMEZCpjwcr9hgchv
8Z+yy40uxeqVtxiv6BqKxsWtmSZ7+jOUKnzjhbSXHh5/I2bWJGRsEhFaUvVEfck4
5epQBmtbWzVkQXtryxrgp8ksPaYN9RHy4YRlHFAqOBMN6qifhjVqaDIWW0jpvMZp
a02hgHdWzEIokw0f8Zadhbl2d5tKxstGUkq0/QyOlzDbcrPHNvzJRg0Z0VsvL5Ot
Na/qSpvxZk/bs6UbWZIEjM4Lo/hPYJQMQLVpESv9M462ZX9h/Muk8Cbm7uKh2Ler
gYh2bwauKc9zq/EdEOGJj8YBHkgnRdCJFv9h2jFSSiIhf+x7tuphqjnFn9MsffuH
bYJpoSMejkECBnQGA8iRyIBqfJfvvvPnAZvETljZ4CxunHS07ODn8ddZnYwjs0gM
L/WWVzjcnWsmfYz/AFKvLantV3dUguMccRv/RaKwnkm+w4za6bZB1DW/k9n6jhMX
s62yOExHY+p1cMeh4FbOSrLVt9JWlrUO8UByloCM3Y7eUaUI7aSXPngUlSNMMnFR
1hsyKRp2o+zq24iLIplvPBrPPdE2reRKIic9ucMHEjSPdjjd6KZePIbv4njecjH6
2G2z40dgRypn1WqMtgtaUGolrsvsen5L6NSZHavSbTGUEg1VXXpIu62drneq7AhZ
PiNwZ4LeQmuPPBnj9K4RzIQk7Dm2LUVCP9Sa6vWXoyQMVxPD/9eTCvz5C3Bbv2Po
LwYkIlSDQBmw+824lTRIZ74uQk6l9eIVM42oLc0OT+aHMFirgmlf1XCZ0bb1b/cD
UAM5Q1eesI8uKKSee3EgI1LDUc24lcMVuNmRCkxhmRwqPsw2ISzp0OSWRr2Ynl/T
28l87T2kRJ+vi9KK3uu17cU+BRltiPF/62PdkK5cSQnioSOH4+3FbCNYBWla/hbt
PDd0cVsLUyT5eqjIopkm+auPGsV6zJ4N2iedEa4ejKY48tpZstqHSEcRQ1yjKGmE
K6qlTAIDBbtZEzMI3lg+LFJkU506upn2ChWU4RzWKNLoMyBabZBhQrlXhrnIMwXC
/7Qzyy+nqb1MhcYDIGk3A3RqNt8KPadhn0MHy77DkaMEACw/XS0imTfoN2KmV4uv
NSL4PRAbGLCzwG+MyGILpuMY6vaCD/wmzChKbKa/I88qSStZeQbFpFQxTTGx/HVF
SWBQx50UAb9KiruT/Vd4rbdNnq0PodYJ7Fo6SmOWA/l7zOVIEm9G6BzAQxTQ35iF
T3uCARdrkHIJd87YN19p8P4kZowibExY8j51JFYXo+grZroL4RaHs9z5IGXusfID
+rafZlyCRSpFdaJJ3xYBaD7woaFiYgFPfRvdjGyiXCgY3e2oAo4haRplXosw+mQE
59Np8u6PqX3qHluKv/B0D02Sk7jZ2VEB2f9Kq8cDuOYyfy6aigpuCgXWWT9Hu8qO
7lVRkecguSNBs8m4vpBFFtV//hxpLPVYQ1BZXAgwSDw+L3u3+SjeH0U4aVvlLeGS
VBs1DxZzRgivd7WdskIw/OLv9YWSBhxW/TJGupoE68VZuohODHuDLNZ4D4FlMIt9
Kazc5scMpij5PM2/gPZLjxmqQ3zBqUVT+XOpAClzbqGP5hdhL0qnBcukRz0p3jgk
8BxfCPe3vfYhywikrfX4J2n+yDMMM4QZYFFZTXOLWi+Bc3xg6o6yTcIUyqeyWfUz
jMNeKOyUYNMWJ39wUz/YZS80MUuE7CwUmU4NojpIIdjHxqDL1YGbQoXZqOuJKW4g
Cgvwd70lRylvGNFM3laXCoVRPOyvlsAz79TVHfmRSLSQzU8Y3r22jc5xVF2BRdmB
ap0+bF4eq9XR+cSvLr1pGntbyv3ZFU4ZPzz6rQ0wo57nUxmSCRrjpJ/V/CJY+d3w
cww28tHIZ+00ciNfVfqvvTUFnhBUMSgX/Xf3RKsNAX9t6Up5dadPV8EtUorws0DW
AmwqxLPRPUcQENFTRbb3oWJJLeECarO91Ds5bQ1ecIFmNZic2P4ND0WAe4AMH3MD
r3SI0wU5QhiTbMLlydAHpqSGzaiA/YoUPdl7b/dEZMf5lqUsQV/Dza/ToDmFDyIn
lbMCPSkV3EJJ0DlIlsRgLAiAeT2DBeOZPGkLbqGN4QR5mI/A8vW2hAL3oJChpsl6
EGEVQkA8IaddfSaVfaDm5XfyO53uKxzbwI9KkcsYnI8zLfBonnZKzOaCHOYf5Glk
XEdYjHSmumDakg7pGQI4PIewXsrrmcfwWKrmWOKRb/bmw8c+b6d8luZNPZogQ1rL
RJOm3NiySpxl8rmefMAEczkGjR9LaZEPBHdeM8rGmFHGJVh/TsPxgbWmwGW3zpWD
GAdjqevliHojh3A4WDvmT8vqbs8oYkSSw/KzO7VLjICA9KnODQ+Kl/lVmTpNobOb
0yDolsL5MZRtR1m0ItPnCziMJbVWElV95KMBSsfdhssVuvRSEiqgupPcvK3aGpYX
dHVotY9hF68pDrLnJjuY/8LMYctMT7ekMY0ArxcSOVdJ9e6uPiqsG3BGd7orsKPQ
kF7Y79w4nNnS1kfqm8gL9T0i5G7glrWuX4eM4wKvXXfQLYdUpZAFI0kMFLIakQiE
Nsij4/3/bSD7qcpO9tCnkkiuGe+7AM1Sr8YKhIqTY13I+ZW4rIAMbmdTbwA1qV2o
jdUo18EQpFpW5yoxcH0P8/VbWqApovz4qv+ffc3Sa9eq8JZJ/aMJqSwF58QWYeHE
nRwjK9xETQ/v2xpYXxtdRKFAiXEDt64em7iul6q6Gt/5XPFrj5OrnOER/HE7+rXx
jfffRzcBbZQ+b78sjrLa4w1Y3IQSciI700cBvhPNh81AQqs//9ljPaLRCQ7oxglm
8lQmZtVRk1SHOH52UteQqpmrrujRruM7uWDtrwOHsVIuha5hq6vmkrb7uPSRhwSo
tfj/a6QRcpbJYq7DuoD8m+vbMkv2OTE9UypWk4PgPnr+h3fhgw0AbJhDkm6MfdpC
stzwDW8qNKI+Zmnuzcgp1PD6A6UuCTlKmJYEge4u9ZpQTwspyxVtrspsEj8LBjaA
3YULAXME7PwCyDrNolW/j362fO2owxZLrmBCapIKjXrPfKAvjkbmmKYp3ZOsF6IT
HzJeqV/Qcq53xgHiSApzW7I/gFh9s9gjXWwwa9RC87E6rtXG/zeP/sUj0dJD8bgO
6g3I5DfbVmjbILqM0XB6hkzzIcOR+5LKAU164GW9YeT2KVAUIh1fUfYfY9L5HWOb
PbczItID2Soq5bUIesuYlOJafg0PhmDNvjeod1I6waJvMIKNnJxqZWceXOS6ulkb
glC7scrxJl7nUGlOGtzxTtghUmiPwZdQf0mt7Uuu80ZgOSAiXqnQBxDuUejE52x/
cvlvr6v22HLC2XqWXzp0hbFHlYfecbeYZ9TMF9Dd4zpaGG22O9707aLaOg+j1M4L
WBmxOHvjWW1FIUSJbKaLnaJKcgfdoFsb0+iC54AJue7IKtnxBympmaJB46NtKqSd
y/rQBbipePlbFDOH3rd9BeH9jGBgIzUDFf0HfVZtJpfobGHsQYl64nrrwqC9Sh56
Eq/hBDK0o2KuJlylbWyCpkgjKogIYR9jN6S5pQpX/0ypLblIpJpHziF8tXqO0NhD
ZVV7pdJOZZ1WdiZYmvq38rLjqXh20Lz+ErKIVjKAgr4QiK67yq5MYPonRrJFr5hd
mQ16zYMZmGrlOiNke7sXUk5u6ZVP6TNkWW4tUVoHCqDGyeVqdq5Xwbv2+nV7736E
Vcid73pgAMcxH6nHEKog0u9O0+kQ19wL3Ra4tyvvww8f+x2yeJTbyMnh9kEzDH1C
MJDEPbN7cyk1p0E7fP0KskTf8uONfJZF/b3YGFNJfg5sq/4xNr/gnTQAppc5dkVm
BbFRzbIxv1DX22tcmA0I3q6lFabitEfNHEPJMXy9tWswmUHq+B66vEwAufqlcado
Tkz+wdeI3NLdPUddTbmnTecSxP//ONQRQ+/mz//fxXEikqIfTqVQOeQeZjoelC0+
eKWOeo0U8F9+ebTskG2jSggiTlIjuNW7X4UQFb+6wjYsOCCX3I7zfo2qBcSh710X
gornJtRrBOZfXMM8TTKazS1sLfBxkCRwbuqL0FXjge1HvfqoapbABatOCVHOiNab
BIuJUpN5pV/IIfnu3o/ubvIAGJsQyaMl4KvtKI/ytK+ZkCH5GIAFhITt97YMBdQY
gLIV2cPaLHuSaBWgqZHYPTNE+fHVaF5biyIbSCfj5otlBxZzeAtq7c8d8hhTnW6+
LiVbR40HWvTuw2Hl5ZUTav8xbVS0VE/oZuvwpkb5XTadSt1ZER1Zhfaoei4w7wcV
3QqIe9qfPd0jW5/yM7mcucHeVP/ExBExw0CfR0w3iHqkRhjdJtsVHXs7hgiVPEAN
rYdTYGAcqin5TH48cYHFEfZyi05KVJA8+ZHciwZ4e5W5w3mAWjDQ7/kc5chZwkMg
N0DbLAxGdv1SqqdA+nrf6ionODJVL+6a7/zHOOrw102eigjHkpXHQdWIiOxNALMh
A1LrF5IIa22nb+Y/nFAn2VuXoyTHZ/l80QHeH+aFZXKb//20SHjxHYGe3QwHOQEa
Tq/f/8iN3ymKu9ns8SDogzZxGHRNyQZfLWNIzwl3p4kAXRX3G0rQ+gdN/RULOhfl
k2eUVXDC1fozcA/So/29ZhG8XpkbHTftPR02ra61Z40W+x9SApPjBz4JA/aHq0Gb
x5PuSpy0fl8M2OjPldj1NOtnFiMwXt9N24IceQiM5gCqccMXDT+yl074EIivN5TY
BjkJwZYnwfdlm4BnCpsfJhNwvvbRrY/8wl9YGSqIBODn+SWQQt3DeR74Ec84Tw7N
CHXtuebEQc/5oeOvVShweY1uVYskg4CO8XSo9DX90Kn6jpaQNYo6WukkqXXEh+Jf
L5Xh6S2J9ShCPCK2SX09PrP7c/jWirFzbEL88GjIbJkg5J7VJoCYKcLoezfDnL+o
ysixvGg4l8w2mj6G64yzhx63lJ1iufgmKWYZ4Y58/urGpsfOGgDp2Cm0RXnh0Q4m
JUJZvaTzwQ6gFU326eE0h6/WTfdIviR5yt7GSHg5FMJJqYbixntjsYGrssgKYFQC
WXf4rbIp2GvtQ61O0/a2OIfPnfF3ssI9AGzI4AjabYbiPRMhwIyAxrJNCMyDv7Lr
snb1yTxElo++cna92rdcspik6IBZA+l5mQVvlgo1zZ04mWJjQB/3K/lI1sIgnLMj
EcmcQK4d7hqWWGLA9Yu9P8ZQL1+M2kFS3HsfrBlXy6lSYQzKd6VLZLuybCdUU62q
ovr5dB9cS+PXRbHe5mpLt2i+OAO9NdtWWLJklnlvSr4zuM+9VQk3+700MyXu+5lQ
HiPy1zJNLofydGYdX2J3spwC0+Z0c7eICfUMooSn8YHHkY0+Pw0eTBxJbLeXk4EJ
qBzfHEK0qT3f57t9y45/wTWYjZvhJegWyMNt7KIwO9Tez7LK/ZGZ1aooarOKR+lX
8uSQGHgQ6uQb5H5WyVKTZeuQmdFNPnGsKdZA21m8Zd9TzzdZXmjqTsXKpGLI3DEd
U0gMRu/skzDMAXEQKUE3sJtiQUDa25jzAdEpoD5z+lyxDAa3vG+o9wP/IZmisqWd
swGUwALhvjM3AMkD+IQdPpuPZcaIDnCI7uGveO84Cj8RUxfFyjBDJ66+4hjHQfsJ
1Q3NJrUSeuswMVJ4v8AZo4pQoRfqTB5EoxoH2+Hfzaz8dAcn1qT2OQYak56b5PQU
DeUvWlho6WJVUA8iho9QdVkiRm49nYNSRod1GXzqX2HMaeg5NI/3hduYcrub7WAA
3rI1f6GyIopfBR7AyaO7FY1L7xNUWUrKQBpF60rFPrB4s4LwHJ8wyeoS1A3SUqM/
25+fe77baa5Ghg2yW5wcPTFqvqf5dIko5w9LJ2rOQ3EC+b+HnWM+ayfQ74XZ8IiL
yKbqlQATQPMBlTDDUXF9RjvKbgvDXJuX7EOGHZUgwqJ6tEK096mSj4eIxSORXbRW
SfPfZ9YtytTGfvRzKECi0Qm13slNrS4VOKaG5F4RZg0Nkr7zOBQ+tpkmSCYqM76P
NkW0lZgo+yzVH267g0w77uk+o7jxEyzVHaOxT8/u6nPXvbgQSUH6lAXU68ipwR7l
wGFx1QlCobwtQ6XvkE89ANrs0SDxs2muuLd5xx6eEXxoinqYj7+myLTCxQsDRPX2
kekiwl87NpqwMBRVWKH/5KQJHRaSshXwfKD0AQFAdudOcmJ/SVEcJIAvNaAxxQP6
0CgMPSKwNepDK7FufPBluOabyqoL/RBV4mdxBM8x6zAPmcHUzg2/3ZB/2uvqxWu0
FN4qwkUElxFIo5r4jwN1Axm4GBvBtwIZh2cW+UhIkr5q5c8ZUu6/Em2fQ7lbDCuR
mjrDdHS+zHNIuH6nQ+yzxXxJmOeW2iDI+z6MbhYMS6BR9p/ViMX6Cr6GaRNytJwQ
UxRfg4P9y9ZYmBJN4+DrlDIqhmDHdzqaoXC9qgfXFweGwRPCBJJcnerr3rFaUrEF
z1x30QueNeAwnaVBHkTMz+muNHTjQ18/u9ov1D5mvUvzexlppkMVqrJcOC5HfvdK
NY1AeqJi+hagjuHQgvIu+kdprJE55Z9yCYWiFm52jy9YbWDy/7v36Mq3ZHnB6zFd
cHiQ0RJwy/OaKOwX2ECKkGEq3jSdp4m+yprqtUltvlizA9p5BQ9g1C+S0A6JHRMz
MtDG4zFImTH3fmtP69Xn261y8TABpeFevuTfRS4fRFu8wTMCJMnGUZXDp5bpF7QX
WYstjlmG7lUiTkV/2vA3VbOFe3agTcbfM7FOJFS0wq/HJ7OpkBB8DgH+9C9j6YIK
C3xCZjAviqUmaPvchkWSa5ImD/vpjfcEL7D+QybcqlbShJJQbeyapobBvMi/diXH
ZdTA2nQmvX/iTDK62TzIc+dKtiqqAyA1M7icBGpfPpeS8gvRU3DcWh+hmkTQwjKd
4Ym77Gk0foyhTwoCjW/HH1wE+qOUfE87UE3SA95zCfR02Ozj8aiqDXJlujKb44wo
gBc79fRNfBJbNFXxM/3fDY1IwZ3bTNP7QOlHOy5jEdDif6mDAO4R9U8L94mHhTwo
jnlSLjPJSkXLLtn+ARk7Dk7zusUDqX+kymjr8X6t3ECzHpTNPeARRKkv4OExdBRq
WppDrgHtHTiMcfRiWz3nZX5OSylYJ7tMucwESqaObQvuIkqN0vu64l8EOg1MjbgT
cip3wi9658VMyl4C408+BizfTl9qFxKiRhwdNkHVf/zuSkuTdqX/QEpOJaGR4maN
j6rinVXHC2gZtERW3lD11AeJGF4P3AUKYDAd5jwfaEBoEQo/Tk+rMMmCnfl+sdOx
5PkQ7HBsoh0Rjp+hsyGcSB2K6frg+cQQqkccP5M1AZaC4CYoXJsT1RFnsekruWv9
b8CJ674jneWDn603za7C7fXrpe4XAMH7FMHGUqy8v6fB3gL5pmaqgojNoUIpwEU+
75x/EBj56M73CS7ZunGNdb2AvdgaMcl7/6Tw+ZHle4Jami1fS7AXLTfnEyVYSafR
kg4rp1wl+Gkm+XEkycmDsYKbCz8kjTldOVNEBSzAiiDKq0PwodbTCs1IWVYjtlge
3fFYFmvAy0Y0SirKAAA8z6pJds0bv+2t3YiKE5epWOpBknfJyQ8RZ8ZoCFg3yDL+
gVSprqqgGh5ABDv7ABDXOhu+xj9lSh6Y6QuyuhazvfZZBo8sgYiKqWFcL1acRkri
XQc5/7YlsmY0IrG0ibQx0apKIM9HUfcSAH3g257S5u7PIFe0hl+ImFR5GYBv0mk8
z7Oj+mNFSbRIe48wKiOXXskoa0gq5cqX3jPBMzZ9OdHdcTkQnWkMCQO3kebEFlBq
3CFG1dvhld7PsCIHO3an5c7gzFKiG/vqZ+IBkKK7VUl0EAb9JHDcMEs2EZfhetWI
1U2vH8HZ17Sv3WvJJeiROSaTsJ//OiyUxGQxRl9ZdbwxCIQK/h/Jt1a3E+eIUCV6
/HjRkJSEqV4ZQdoBtWE1ycO9nHjPBh/7m8pjCa5dy87yjLfBrFcuLWkrWCWmuuy0
uqAe+tEEOB4Dnj1OSvdA8ooizuKHnphYO2AJCURpcEBcLP5bcmS2tt+RqzWv1y0z
CR4bXPWdTHtl/4eBej2ZoFpLfLLLxmbIWiX/hy7LBN08K9iOMeVFc6/kkKZMr7vm
Rir43rjZqHjGsfE8k+6q0eLv5Q1To8lcYprldrdA/ML4tYVDdJgyclCchfS96Hv/
/KsWg3JoX384rvtYRkRPLHooVSp6zTzbz/q/Y8E7jyARg22Jw00gRnenUz2x17Yg
Ki69xsIKjkgy4b4/9xrIasQkOEdJvVPqoncTA9wZFF/OfyZQQMSgph0TW7DS+yL6
57i+tnz4fmbf+6CXIc2+MTLLkIAsbTVRVxcRvUttrJ1Vq2MLvntqQ5G1uEMWM7ES
p0Wvjp7l8Qn3XwNwwaDTe2n6rMVhNqwTua7xxpbv7+9y3js0O5mFB5QChFESIgHN
L7hA0qYa8kY3UxLBQ7wPNMkZb6DHbHe6HIfphMZ9giAP3kULGa2i3/bk9SrTtevf
pm7ha/DcXzcCrTStJQ3SROYTbuta9SzNquuIrHvS8u8lQHfdjTqYRiH9i/weFTQ3
CXuWPtmeRqK/54blF69WXYa7frbkmpl++0Qqwe9QpwI4Lo/FTcO9SNMaZTOxEfLE
1yzzigzldsV6SgF3Y50RPXLoMppQCR2zBAw3mBJ2S0BF7MJelcjS1RSpKY+3wzGQ
kJrY/E5y7koY98S6zSKDobPRw/psKGCSVlGEmbF60My9DRIA5oPf2YaLEdk7R5tk
flW+oLeNBoikqfe26tHXmGsf9l6i4pJ+uvwhORFURXUySBsdTdk9X0vS6VXiYEm4
LOevsBMRaLbx7IOuXExLWaQg0ZqLDEa9tnNXWDGnD0fvbB7xBbeBkKkoGy8Ra8ZE
vuVXaCi60mRfwoSYi60Hu8tbaF5ix4ipwtPkQkBf/OHGbx3nYhmaftbX2CtwB68L
QO+4PUkAZp3e+ZZkWkwFks9qmvdV4Kzo0xbm7H9LldWMXR1jNuj3hCVnl77urtHn
dagQ/j58P82IpRE6ZfFdUWmSLGUm2LafFBQA8A0YmgzyjLxo8Y7SXeVVWQT0kGDW
Fy9+gLDYw4lvAnFSK+V0zK1jSGRpNahpzUOszvyE7DzyQzZdiGjlUYFf8Pt4T7nt
QhxNUUAVaRamUUzV1rp8Wbn4EGqILezaTz0bUqgh61RNxXaiH0ayeAgMV32plrP1
4u7YEDDWT+tx2CLLqqnvbleJouCJ6VrXutQRSpQ6EoTWTW6qxu8g2fls6CiO/jnX
GqCu8OMWSITunBXCpdIb+U6ZO9OytVFnoSZ4GIExUcRYKZltFFR/rEf34n7l7/7s
nIfbWi+X6lCAn7I3ioyiyPzUfgaV9vaI51sq3bnfiJbheLeT9nYqCTF3dIgdvMwj
9cBWP4zyWJ0PZ75v/j/vLtMzw/3/JwiuKs6XzQrbkMHfSpE/WLSsvWBu13+awU/p
ZI8PGd1YWIFlQG57vrHPcMc24z6vd/R767McPoFw9etaZb+AEDmFxeA/KjnikBSi
5+bMvUjrNm3wdS45zyJpxymCljtPPhmJTds2aCj+O28b0UDr2K1E8qQ2vdZsceFK
pVSTYyfwmLYg9YMh/odA6O2V4On7npxRIo3VZRVcmMbz9UsDgtNR83Iz09K7YVmE
4WaeR1ZId51bbu/jwUf4M8Tb1qKRO8o078oBqq3bWXUUN/rPl4oFI4Pi/iXFw9G3
jzI6tXftC8/ktIFw7IESIhPqxECx2/yNqv8T3gNUMKwwlFeoHpXec/0HhVQ2jaGV
ujb+8Brv4nLYddrx5reUp2kj3gkUqxZK1VE229StCshoeLGAu50NjJzkFWhGCGFJ
lZWi/thgyxYeEVN9ZMlJHsVpMRp8Hc2JipSQnh5LVzK2BOjwHVnTo6l2OZPw2Dny
l4w8XP0nm59ch8nc0h5/bLKHfjy7k1zHjTLKnq0Gem+d8XLaNQj+XkCsaP6OFKJY
Gol4L5QJ8RJYy8dcA05aR6zaViPfoygoeOXsZJMTIb4d3YIca/g3cezqrJ7il/Zn
AHw7DTlRU0pX70BcPfdU65Cndwy2Ugl3QCMAkOfgLsBoQoZf/FCoW8Y5tIlGHplE
c7VOLUhGeSmuVq/NQKng88S9l3dH5OoaGeW6SXS0Vr9ajf4wUAfbUajLNCrfqTdV
1HIi+3KXb2BkjrF6PnibyepFZgNa2bfLkZkK9ifOTqeW7Rh2YEoghpxEikiCkhZL
Ey5T1HmCzuSZh39Db2JH5DwJqMdt9A8YAmpAK6sbBqf8igY7GReFXyHDj0iOCd8v
my5ZwzF1i0gP/bMrBcI/mdhmCLuyTSqe857OQHFVgDGKhVDbEFOgQLAHicNc2XOQ
6Qw0bpA57Yfnn3yfk8RBHspvcw3FaWgZodnUI41LLETtZjqj4iE5lwOMjHnnw2hO
cGopGu4jFYMh7xBCvlwDxnf3EA7708ByYpUnlIui3quaE/G5LGpQV1sbx73j13xy
cC7uc7/giPFAGdKiwWdtTDv4rgEj98gMKcNbxxWuiyId3ljmEcRtPhMzlWMSsScd
FIPv1yUcebONBFOtb0wyeBLwLOTXUYpi1ep0n2J0Xa9s/VQON+W/EVugf2wH7yrO
4U5fmoRwY1oeRz3+7l+C9it7X3al3ZZw0S38rQ/XBdgY8V8QWWKqWv7UGwJx+oDi
N+hWOULSScM4EB+jji3PWXO/NqVnP1IpOqXVDYReTAc/J3H3LGRflqyUgFSzxiga
Ftt2zlQRylo0cxLrAY6aw5LMMe0TzqKJTeeQoziXV72MyMJ32p8sGZoFpyvhjuID
6uWw1oVB/j2NXQnP9232N1QOpQrPNQUgYlGleb0nEtP9r/HVI9W+Y2CXo7iKSJVA
AKjZxy1xEn0BvE8WoQwnvQFb18ipMhWWDQswga1JYrSaTzfXScUyJi4m6Eazg5eq
vDaKjB+alKR4kQEu/j8cGh+/JbOQLqrB9ko+kDVe6JZpwM4PRorXalXar5dNKJWP
XSm5O/PA+95F6GPXcZCer0QnOLMB9QfYxPztDhgNa9hEQbLfSPt3rBnIqKDK42lR
m7OhNhJ3hO6NbPi6SWYjaE0spDjLkkF0ZfMl9m1L+tQL+lC2BAPkRaOwDJQN8e4q
8SVo+NG06/bwzGwiSDKyZue36j6BZM4PFKBek5RmnCDHHdVhCyyn4TVfAao4G6XE
am19u7WrZCe/WJ7b6/CbNVAbHUaeTn1OO5+RHLp+lNM02zcQHYAq9N8/0OQJti34
sGC9OMqjnMQNclW2kUPvJHEYannIcAzora5+dlIJsij6C2nRCF6FY3mWsQyqs6wB
vg8wdBUIrRAO/vLyJFt6gfPi8So8rkEByfMTy1G9tx8+oXd4W130OC1tB9G8OXoR
7wuqNaGoe+gcmGGs3h0PWL8BomoVDSAZpvGl1+8zv8DaZFdQBlUInuRwsMpwXv6G
XBQxvO389xLcpUgyY1HR+L9BVXwoHxFreYuJtCKtLUb9f3vBngUCI7Mjs+UmZmnN
xmbvf38DXcugrl0DdOqn/K8YqFTr5aXe1JL8JDn2rfbcGekjTcfFms+pyJjNQQSv
qgLEHqwsSNbdwynnZPzrOdXvXp0rxpME1cgkkLIyuMZEU+yYRQ/p76555wwKJ5OK
UbIuXnoHB8A+LZYnVWov02frr/kR/jFfXcZ7D72Q0LqaqzI3O7shPMB0yt0z6JmH
2772F5s3UnIpCgKpqAMPES2a8Gdy4Qcm4hhM7+eH3xAOR21rnTBapP2hN4FzzE+s
DHZG4Tkoye10rPz7iR3wh3oVIunpQcScLG8O+lbpdA6efIpUC7GjbQKgwpC5BXqc
B+47n6EYwQYRsBtSWyfn+6w8rPu3Qo/l38jiFNudRqGj1PCWwK1HUPKsxSFNcGuF
VbUaUmw7cPCPfnUQybltYsIOyBR6rkdBiCgiyALZ/dY7iPa/cupJCTd1NoZWlAWJ
aHPEdQXEuBt6x6qiqMZp+JlApJ2+8GsGMTVj9r/ayLKdC4wCaUKCt5GRr9w2eMjC
iMo6EKxSFIdqdF5t2DRMMJWpqNm1B4z7U98X0wEjCoZlWWUz1Ij00NCeNswkp8mW
E5r1TFZV0kIsNcYmU/xCNOSD0jebGaTU1GaI615IIW+rxpIw1os+P9BJUKPdu4wd
Vuxi3oYVQLutMqtK84f+kBRtONH/HNSgBnKq8FEK0nqxv3oq6K1xGYuhRm53HJ0o
mrI2M6+qS3vA79wK3QRlEuylMlptBClfd+bVRFdniIGZs6xnNLgGXeICQw2SWVgE
G+1QTZjhfroG5e7cdKGOyN/s70yBB9BXw77hExw+M5GiVp6lDaM0FZXGMKc001vB
iPBAKMLyFKrRYkoQrxyLVFWbCxekGE3LYkBHqAF8YvYoPZyjyjxAro51261iVxCI
FJRCUq7mCQbmGGcfC+qIfWUCSQ6Q9OkzUwigvxac2zWv1NLLIXXaGrSIqVB9CmEW
kUZKu01bl/0kFEOPXYs1Aie6+4UhtFCFfevIKdxa6ve7pO67fhajskx8YYUp5moC
bPpeZ3Z23BHayUTYFWWsmS/kS7t4Rg+B8cQXTJDWol0zlzwEgfyN8O6bRyVf5V7G
wNtFkMPvh0Spv56kgWZ9J+q5uLLO2inbOhf7FTdS/SAQSkXv0MV3M6RgbtF/Dhcn
QLMmoY0GMBCvdbZMfklgDAcF98mq/9foV0iQ8xMC2o/4GlLsDRqlP5xcQPeeK4bh
AOKw3Q07wXEHQjcwmqe4S7AYS9A5dZ81U5l5K7dBM3m8nvpOlPTYjPwlYwknyyFI
I2Fbwsz7KpAyf5SZ02t+lt7v0bDaFinRUrkMSnBJehmnFynB0pxQJEu+SRKsaz37
sR5uhcNuPGuw6kT0jSYUqbVk8dwv2TLxbgjKGXN0j6Vfbw7hyu1SQntK+OQS6yTs
O7ltkTdFzezRpgifPQHJx9VoABjwhpBfUI9DnmTLn15oj7b78u8gGsZ9ZHQu9sYI
N+RqxQpZSGZguPqssPp/5q1YMSOBVyNrN8KyTjgXk3lbMNyq/zM8OMNp86mkezET
n89MCHC+C2t/jvnXYtIt+oscyB6cBrNAzCsUAUCo9KxgBiQ1UMtMYp0g/QwV7fST
bbnLzKRVLSmJyTlE2+I8V3vco6AuPclg4LiBfKxRE4BylvdmFoOk1AqTEFiJlWap
q0sfbiQT0u86XWS8tK2V6IKkVSfL8N5ApFz5RkjfiLrkGd0tJRHYzz0Toc3kPs/s
sjZvXaBgAIIE34wQPZcD778PhkGkXNQj2ktIi+r9Ez64G3bzUBKpsGf0oif/OEcx
5ImbBuMGXr2s93zWZItXr0LOldgqf7J0B7KIEpVlZJ5/xGIWs5LomvyLysJMYy4w
oplTRuWlbYx1KuPd733rmQU6pHTpKrCr9NMH7uQIxPBDE/Z6I+ftX356XsXSz8ok
XvrHWvZAUlEiUU3AsprgNPW9H4MJ2zoJP/i9003ghEbkCV/iPqz5iWTbXa6LoSpC
31Ctk7gnvDexp+rGDMiUicubKSkX+qG/cTdXuuQneoNTCnO4y4zRzTcfnqdb2Fv6
CeuyyvCTlEHp9Xpck6fgE04AkzzigTCgTLl/9ZVQEH+B2uSVuYw/F+PqK8ZAE4LR
u0mTGOYjtzj87SVOAP/lnsBvUwAjcTzhv4BTbsA+wePrRzsSEb/oYwooZbxaG/ik
B/Xzyofwwd29NsnKOjBc3rTAO2rcLHFnOvy1WKNyIqkCIR4VWWnHKqxjI76L7NMh
oVRuU9qLbArhKnSyejBZZoPSNDILpfvlELsifhL839z0+gsm4TV8TRD3qSCpMzwj
qjVL3pfOQxSbWRrIJ9M56OZd6E3nHY0XpnhQmS42LvdJFKdQEq1RkVAymGvOJwB5
wpGTZ709NlYcfhsbTVIXmlBMMGr5AsR/Vf4NGWDgulUlKGNJPAsl5OmLT7OMYTrX
NB95KiQ2oq35hMeJqN3NfER6eMSDd6v3BYiisS+PIpRel4TUhRVDLAlycyCTi7mM
2DRoE4RQtMaQ8MkEIj5jb6bcdjcE0eJfy3DrJeQMXQaQAC6DxFh2EbdApHwMhcf4
TvfpWjDuzquWeYnvZb45cyIrwrNcjnL0rkoxQ34hJHjflH5H87j5Sd283Sj9IAfc
wj7Cu765a/rgkT0PMxdr/HFnOCGpy5SvTAFM9pa+yz3u4uxiCzhOEhsCjuMgvZDB
7JVlmzcWQhbo/dbTtCw/6yIXhYhrncwz34f40rZz0EHBGXCpL6zDD7lAeFasMAV0
cUNdn5dZurC6a5dcaM4WQFZlQ3WPEp7teRRnDwsziYBzjdVhb9Yeg7Ommhv1DJa+
OR+d8g/7p8CwPgMx7jjON60N630g4hVr2R5y8F6XiNemFBOP3WG2xvYXNM3aDFvj
BqmB9x9p/Q+RsVa58cG3Hdm13B4/0aQF4rynl9ZA1LQdbZ+y3BlOmwsj7hpds2fb
sIPEr1SAa1cOs9mTCWzKeIMpZ6xy8iA5Njp13LnSL/Aaa5jZUPLt+KuxzMHLR824
8itaPfGkO9MlO37x4hvCIEdKZmDkNnjHAaB8W/9ZyDleNAoZUM7Vr9Sf/B6A5S+V
7T5iHf9Gthg4WeTQCXqU7hxXBWWWHum3G8d54xpsL22EdRU8iSq6msjsY4RUEJa1
vNP+OtLvSkucmXA8DmODNbQg9MwnWAE9NS5RYEXGGCcb4n0FfWphoIto0IP1oyYt
wgrwzNStLaWfZoUlSPgrbGKKLVqGQNEPuXHp99zONUHts/cWOXDbQBPiwo1xIw49
GCjwkuIu9igq63IKm6lPLCZkXqQnK29+FNRw2dS4ZXvWbujtAidk2XYOpzo7cifx
JNlRbf96gfu5tXnAgCS16hA+wDSng61AH6l/79KudhJ03NNUJuJDDLe7l1rRiqrP
j/MPgghuR5H46Fmtz6OmF2YTsR/La9mjz4vyTu4PiUdxeS8VPF4cXTvE1D+r37wa
h99o/mz97jEKMqG8+2uz6ixM5L/HtpoWFF+41a80RHEXsGyhOPOPa9nEUFzILgM8
Hnx2qnq6ujuhVJuHnrhEC23UHFBVNtsEVRntsUUw+dTDZIR8PjVc8HEQk8XCJ4ZL
iH4Hbm6bo7o04m0MiHcsR4gSSgkk/T2JMu98/AND84DuUY04hnTpJroyHspJMZrD
9ojKYULsCzFaLiE/WN5fqUADmkwtq0s9LK6LT23FmFYM+VaPsWQLadVZwoFZC4tP
Bw744McgOtBofI+NSfQ9rYQyxFXIgYigLqxNc1mRBgys5RJWEJ4AKgcmqXNrkDd6
PBOvYX3KJKE1SoGBhk6Iuo1eQBzvnc775NiwM804cbRFupwBrK9wPJvjbPqEEPGt
G7UJhtQORCfhEew4no1PQyjqP6+Lq8fB4c61byWDp0G8ERZWFAJSBLWNEyvDNImy
+S3S9AX9DDgYSrUDtUrPZtXflWLoJhedi9SD/tD8YIf3fV+VOxdFHDzRjo9f1mrV
qeaAWY2hPAYHzWiQLFZNzRrXPFjeL9TMiFSf1Ek8PaI5weHgVpQHo4jNEFFEGe82
3VASJLfJaAf3UfdhmPxNJ3B+rlagnenjxUd0VtBb3rm23kFsJFcVWyekOF/Cr6nX
2avPsWEXd6XOEWAxyKd2XVaXLulhPBvPbdh85O/fFAo51tDLbtHvlqSSsh0wOkIL
8nof9rubbsH0xqGHOx2uA+ROAQQ9VNSxfaHl6HcxC1YxRojejaxL4MZwNcFsfyz5
e4xLOR06j4qD0EK5GhE4W348ORyupPvJ91TCYE3QqHv4G12zYQISnl/vBEKCNvqy
BTKidiZIOqsZPBgbIKWa5IE20nOj6TP3dUpNGoA4Rq2SWMcx78yRWT+TUQz0tBMr
uTcOkDqhMDIIKLVkRvpPkEs3eYPOTrvmaW8HKZtp9GWNZPXDIQR+jouhq+veOey8
UaYFp6vZpWlx4q9eNZz52riApqCsYKn7tA3t5+mkUGyrzJ6ACRmXKmVe0jzvDeDP
iyBfB3x+4tssqJB2yz5I5qMLHg+p3nIBuQLmeWTuynqtU/1kBhbS2Us6aD1idZWW
h6HrlLB2jpn5MytLwTRXRpt99zG6WLKUEl5xOazQ8ldOVZfvOjWDX67fEgUwBfok
sw1V4LRmvJuOHpxM46hGYVDIKNgbHx1YKNWcNbjB7Qw2mPEmSa08tqraKtxxhYjP
Hyq1KkqDIAmOTEHPoGS/C+1QVhEzlGKuQPFoVWMzjcHjfRhOzr6YceBkcyMuNG25
7sGbfPdDCn3+6d6Tmv3H7BjGUd6NdXfBByG+E7StvM08YVmi3ELOR3cznad7tlzH
5LaXpI99CMIRtISXEsS6nJsBXQGDJdT30rgbs4/bDrimuTjXMtUcwiaa9YMLGD8I
njeWk3frlFqdVNGsnpNVELkqegRK+pVd/Zwbk6SdTDVE3OMfxzoXGu+DaNvwo6gp
TZEMgopUhRoHkbOcBCiublv1WZa1Lt4PltoqjCJQOY8bSPppVRsoCADoD5WEysft
ohRnuQ8f3O6usjp5kXt8C6eDS0rjwAQGZJwqLYd5BjMuJJey76nGqnAPpov0RAym
olEVz0tsZpFyAM1uXtHdjhyKRNP+QHTcqQl0j0nEMhCHZvMLpMF/PZV1ZF8PTksZ
h0jJuhIHLXt5nM3q1gZROKpymCp6rP/uLtMzm9m+HxIOTGrbsZ/p3B7WUmYsZ3ig
VVrAZuUgri0b6jodp9n7L0ZDpGlbXEO0TBfnKaMjwqEIxSJS+eioGn9ZUOaR6XT8
XpZ6z9oJIxh+rpcZGiaAFiKD0tig1ZfIZAzsBF2NmQ0c8Mjh9Sz7wjglvYT3mGYB
NHv1JeYqqIRgqhR7vd1wpj83NYSp6xQBGYsYOa+lBvnzEbHXnI6+jACxzaArENE3
En9h8COIGSp9pIrFey+7pv/uCvcJFbV8pP1wqQidiQwtIFRQANxAMK8xBtPZbASh
ta+IA3YZwBt3Q08sc6gUaQ9pZ4h3ON4XKN78+e0F1U9blM7eF9L+1CLdR/oboLa2
sZAL1Irxgfr6lvZcPAb7FSi4RWGaX39O5PKgr7d7UVksNGwhB+ynEGw9tnZ3s0gf
2OsxEZxCf3P4v/trsZeZysBN96OBr8lFV2v7gZzAG076BwkkNrowDqVkdMQ/JeOM
uWBoL5SU5/DPnU07QE+If+L186UPWGUWoLwyaNJT9tB48xbXtnSM+2/gk5D6Xzp9
uohVrINX+AnauLXO9b7yYHylHUJ7lZyV136qbcBD48y0o/55zS4PcPBUFtDa8S6w
5HmI53uRdbZ7XfzedrISBSSPkxC9E9+7bANapaueK4BjwVU4VuPQ+NvlETI0VSRG
n951gWcRcpPky+2NfgJKgIZT+7V9Kjf/fAq4XZYB6BI6WkQW+TqlUufkQ4I0zUpN
6ikM6TNcJpLcTIBMowJ2OcY5Bw2pdyH4o2AFMvEE6e9M7DP8xH41+/IZsTvK5tcy
10dYgyLRLxyDV4yebN8odGONjz3h/vh8VyocTpLTiajwr0gijrPQ8TTqKvVXZJqT
3qdNm0mb+O9lqyvNWYHw9yH+J11eHbRD69dh8LbwgA6YHrN4g8uGVA4t/mkC3wu2
LyIC3qEb4pHTgS7+7Lb3HQ+02yJwJdWyPmnAlFqZrRAuBEfg9ykR4xCUmZM8aZvN
TKFTfLSycA5Ohu+pQlWVhPH/Yj1bDiKhxZpvCIkYqdULc3XswmsoJSThMGKIojR4
bj25pSO3R2r6FkgaTSyXQW0hXgrQmcKZAKagmB/IhKhLdy2Y4e+g/krMdY90lVCE
rHr+b7SRQA0WhJteDQeyUmAR7nyE5V/qlF1KkQ5gCPY6OVbXkxarwUbw9AUgZc5x
t/w24N9uJnyVv0lLWRk7Bkyil2EnKiWClZr5TKTeHPvlS7B8WgWbhcc3aNFciFos
wk6OjUAWQekvufFfnhACAltMnG2vIGsLFbizgNLxCZlOGB97+nR/MreOrkhLY/ti
njl/4AM4Wn0wcxtuqyiSR3Zp3Jr/aUM1EkacaU7rlS7jSMARuRhu4IuBQDAz243e
iK0iOzRwtxNLyjc/4Kc9y7umunHczU5H5Gks02aXP2k4QgsLiGSKjjAHrHjfFwAg
E+gfoKxS7sUBMoGDZRydn08Ur7QgMQSwyKqjpkLigV3q5IZJnRsU1J+g4NVsBYFp
4AFsPSD4cKEQSyID6siZarF8cP/2lRpbvj8kCVCtn6QEDK7qhDiLJ1fGb5PNDr5K
1xQeK1Ph9dSuSBDXeWuzMfie1GdspZLnfj2nT4mowzAO59iAJUtTxqiAUvwDCHp7
d0BbuMY050MLJsNjdn1Tntf9G7QkmYwy7mRUShptuXZib1ncJ5OJnCs90Dd6XGZT
Ki0S3cG+AlJY3PP+5pquIHMY6C6NIGZvFKtwWEFiS/ncp8tvdzSpkKmerqi+SId6
mMw7HKVgCYHCoZo9HP4DAoJrVt2NeOw/hgm2HkRviUBYF8SifPthf8ilAmbJQIzt
g5v3gXxhbvxUrhrwOE0cLA4yOT2FXHKj5b3vdg8SI6eRfjx/i2hcESuvQU85tJJh
EfXXlJuT5W1gQooEZujXg4Am40sxB0NvZzPDdHmWhzfSBiIuRWMcUOMc9aLPorjg
cBoIsxGeWXbF9eZxUeVRP76Qdq9kuotT5hahKk7CJVQpUJzDCkjPLLPdOZc5sMcM
LWJxBvCMp8AbiDlG77LbuE+WGhys8M/i5YMAgE6Ybg4HtMAe+c9FcFyL4jTX2kbC
JeTMB0cSZUPW1XNWm5ddecHyHo5RVpXlMi0UBc6q/p7MZMkBU/F1PS46uX2/cljJ
poU4boDHwM/vG1/kM4uclFlMAHkHqSA/Qqqf+hIx7fYU8Nu3psOJqhAdfrljGWQo
JscA8QbIMvIWkm+8fQDCuyYk7vfLAyyvn5+qz0P9ByFM+ogyXS7QnB7zXrzoWbYA
OgHNI5YP3rec3BhnX1GU4YSE1qmXlSr2QVujHfpbgJu5vfy3P/n82LxNTFU+S0Me
Wibf51dZIum1Zs4S0ElR/smJMmH48uQCeGGlcGuG65pJuwgfwkuVCynmzrNPw05I
NmdC5j3S3kRgI5xYjD6YVVYWaefW6aVN01bISvnXvn5oWcGCqJV2yRIbnGpcRxub
ecpk2uNfT8pTNWm9vXah0KYqPhapPZ4w+0BkVTa4UZOEUXdONx0rPYnH3QZEhJ8m
VBILm1L6DcFDGKm3HWNr/1SVbT2w9qrsDnXr0iUoR+PuHAaPnqwhyUggm8ror6xD
evhUoNL0P8jyHAPGEDKWHcOZ4RJe95QW1m4umXDv1vHqMT1wEK5dnKKqJ817ul7y
3c6r8IVG2OhEzKpIWaE8sJiOEO6eVpXwDV7Ywqd+W04RwXlpd6WLsqc6KbgWEhon
4edGeE42NkvDkeo8B+mP1bPJcBFtfr3YVvnO73gYLWCmaqQP4lH5lVEDrWKi4WSW
JVSXrZ83fZhNiZ+5IUgB5UXNv5FBcfCdXVGf2lntNAFj3N+c3hcFRQ+5XzxEKbN4
blG5sERtX8KCXhkCRV3judgQbrO0ASXvDJjlOAKSJK6Hx9cJAz1jNMmSb87FEcAu
u25MOXya2Zp8IJnW6WZpEqBsUQZXrUk/+5OQ/M0m5j3ah/uoptjkYBXbqkLP+dwK
mVuR7LB2m+D89k6gZpcbfsMLIPqHOUuRk6pCX2eZAbnEya5Rtv8ZsdPAej6AAWZD
E6ww5y7tM1ctxdv1XRvxeG6XoRkBGpL4bpgumsXAf3zacwsUImsoVV8iP2GaOcP+
t8NSLJe8k2kjDZWfhO+qHhf0hdTRJuteicNcg9gNK2/7s/Yd+Ttl0q/v7aK7rSBz
m2wl0l8EZ4VhaKMLFYDD8BNsN6HyYHm4TNuBOQAJ8Z8tiIlpPAhLE9I2aVuG1qaE
Ugw1gblmBYtf4nm92DKRXpu+2rbw1dE0Sjn77Vu3aZdNe0ZYbpXUsQfIZDE0Bc8M
n6g+CMLisuqw9HxB5kE8lmSafNqDExFPPj7BSjKuUHGg4TxGrfSqTwXdBXSq++nx
+vOTHbBo7TkKVMeqqYLYOI7xXvcYL6+ocLLeSckmB8HtCTfJNhJWe6bXM+6y8scF
AajYlzWU1Ig5hQFjkwFGIbjkm+P1InWCGBwPi3mKZnHNZa89RztLHxToHeFFiNWT
xXgIm4NZhq1VKopuvaIdIzAycdBOZ3kpoc2cIepgOSi0WFllHD1PsYgaI6MPRfRv
PY45kdEvFL4zpiRzZSPZrcFO/WKo/HzaUHhvFTv7V7/owo3HGDyOIar6Y04Gn50V
uSpFur0zX6O0O7BfIyYa4WkDo39nAO+X8zHKo23SLWCaVOKgiPzmDFMpIQVYz3WY
F2eT7jqodQF/Hk2NEb42Bab3EVfBP7zUnMeHKyT/TCJT2h1Drg6FJq0VdmR3BebK
wRWp1vXf2Dr7suR7SD4EOqi9ls++qss4fbO+5Lu0jdUxu3gXAG734WhrAuGZkJBw
c1eHteoiAQullbJIOlVQeV1A/5tHM+jyow1Drjz084GUE4RBK1JStnhGXLI2L+M+
YAa9KHoSWD6WXZcVHh3yE3SoNg4DGBC/N3N1YrVpVDLISXKHvEVJphJxCR8dQVXN
ks2frXcf6ECQm0yLukwfQML88iWwMI6FjJKruZLplc6Lv+RmoV6kUeWetPus40pA
9L4uI+D7Db/7xtVDCimgxpMtqv6Dvk+aYXKvvwCNI3ez1+FFC7m9rmaWs1SsaZ7c
t4vopn78/VPkwxiuM4F8NKpxwNWRRTtPdAPwBGGO6swPH9F0RKH2f2gmqN3Xv5Fy
JzWl1S7HGQcrXYp/GZMjGk+IDolihnLm0jdSCTsLauuJazk1rsk+n1SG9IY2tgkx
ZOea2lAOYEJ3PW2Q8Pu8fYXY4TfeF17tSqKvhyvcbT6ZYfVF0fX0+5jLMLv8Y+P9
b+742LlMkNJugSSQMA1EyXfQz9avVL9UGbbNuGFxOKJjnBYvA7RkwUfd9+SEvX/Y
sJrvB6VBhJx628lYC+H74Np9AT5E22DE5SRy8fF5SLEXbpjbw8fl8U5k3HTC0HrU
S4BCvTLMbiGXI+f3UuoxsEXxK5bpyrDVudCNT519hFlPeCV7y14ocAIEmhg4SGSd
q1Whszy96Mq3WABnVaSxaYqf9RIWjxg9STGhhN4y0g/gFerFRnddqHqT4pEWw2hm
47mv/WveAaJgFd7Xe+yDrlCNljosfTjLS4jXDbnM7JiE2jIjLtEEym8kcBDcREXr
2aMcErOXUGA1YT6xlbW3R3O8pxgcZTmKtfLRZUKlTuo24JyA9/Aaj75p2hJD3bnd
SE0cyINhIvkN7WsS8IbH0y4fVl6fRnZ4kB+HXZZ0Oq0uAGQ+dp78gBGH5Q8v+XEc
X8nYQ+RfKXosu+t+q5X6l8IRc5fpCOMiCtW6bZq3m1KBwuDzm/JXgTJFqzsIOdi3
+By4rq0QCv3KHHmgqxR+Y31faXOmbgYhQNfCcYQBmN1Gx3DKx4JaQ3Lhvq8+xhtq
wa0eoAvUUFP31y+xzy3Uoo/nPXrf2VnadlXDbm1oPEgLS4sXjeX2hswjwozNFCpV
sySFHWBC0c++O/5Q7W8aWA3xRPteizSljSr1hbfFulTxVo8f3AJHLy6zLf5BVsy7
DWVmvbLlc9Jh/pIp3TQAqxmf3x8aLPGIqGXQmmArXsNmDmWlaA9AHQWP/ze9TIPe
O+zlotFy4XdpcKtSYl3Xp5+0iBLJ1EAtXEmYH9UNtS6FKFngTUGXXmFR/VFPgg5a
84GWNtuiIJr/7Hzo7WGy0sNFMxVVB29okD/FhE2jCjE2LpRiC5x6aI1qcLJoBiFX
q+rgkFVXJqEGCxjdxbncCXZ0+8/jQv67YgvRpd3iK2PcjA5uKfKqOjtr/yw1OGDY
LCD2fjZkvBoRoZgSIXfJ6oJhqWE/7iDaig2FpkmtfJGJ/cbNsVyFZ9SB4PJOOGyw
MMJGgFO/GEbiD1DC5l266uLDJbQWvOw5Hp5jeXAxII0tWGDMVF0wk7480lukNMRo
xrRBdYyO2QfS28jTYlcQWjs4lPcLQwIg9CCsWmvIhsI13xk+W1Wv0EiCKG0mhzix
IQQ+4HgtfLPV0RUniqn7XXZUl0kIaurOnFti3V4ex5soCvJ+jCl7BzmHJYvGWtKJ
vWBbMcX/HHwRNs8pUODyVjQSwzzQZq4LXxhIM/VhJ0kFKBUuK7H3K1T+k5M2QAhj
QxWFhg5xp8gQClvY0oNbI+RE5/J1UCQ9FYtZBxQfDofpkBHRUvBnsENIjMg+VX7i
Gmbo47HebKXcjO1N0e0IkAkveGgzqhtBdrCdNp6jGgQRrxTxqARAEPkkd54WKZhe
HP/+/OAQw3azqgIj/NCuSBDVOM5fyirTafcLNBeI3ZLOjB2v71Zz0M2kR7k551EB
B1wLm5LZoEthuUiNTlKLvuZiQgMjKmsjaWPBF3rCBQhCzoSsPMq2qkcWOAksFkmI
kMqRBssBRT7Yyh9vDav0V3tB3SKu/kjmhbpM5DkRzsprBlThvlO4VeVqKAD9zU5g
9HTtfIk54aqJ2+TIfyILZdZ8gciJ/7eh13FwaQCao1NVJ06EwpZXTMS1z5eTzjPc
uZcAb9qHAtXhs3TVPNQtEJ88aoH0Xxbkl2pz2qwJiuoqGtthdDBPwvkNUReTLWmD
sVk6NNZeVEQrznzjGSB0B+G+Ykwv5a4v9qsvyNvb2p+ZqgoSMi2u4kMAC5oik4yE
ZjiMtsZJ9WDFjL2I9ZPEwlS3I68zYghX4wVb5g1ak4vjDxgcFQbwBR9Doxc+7/8A
UIm9G6FIhEgWFEYh+6URTERgyYTigmWw6//sc36URvfOYcZiJz87pDJtj5M8D/aC
N8kgCRG2iXK2If09SdpTaN++RA/HZ2RIRBO9nAqMKBtee0MIHx4uFrA6v/1e2RG2
16/yy55j3rAL2FsgyBToiO7SnawO2ydacipZRV/uEOik5v/n8rUOyAHIPIehE9s3
2LNH35AZC3+8aROEzpXsMra3flqTpGliMzHRRUCpEWFXBfz1P8sBP0S7OL8Newo3
nwhpXwpCnTEs+oTXVzr+debCKJuCrj6tFF65/9tqfKPMlSPHMXs+y95EYauHxPlX
/38D66I1rQx7Wts33Oh5rASFQNb14gveZq77rH3zCKR36HoGhAVjCR9YNcIHXXGH
VyFxROsUDtCc3fNxl2gdoaKdprOvnN0Wh6UNymBpPTDZL7fXSXgY8EvGbMo3SYrw
51pLNaX0AwK2nYKgS6gdVO1ye5WGXG4O+ljPSutpZiDZcdLjyILSL7vUUXtfuCpf
3MogEc4hnIXE7DB4WdwMNqSfyI76DEW7VLwCN7LdyjHjFZPQV/6hMRXaUBwbwX4e
IoorYdWPx1IV+Ap90rQinvCH6/SC82EDsuRhhCQrAipyu6nq3sjKbNUQpQ2N37BX
oVrHsiEWWrq+p0BXL8P/lkE0WtsWJ6y9comWmmcgimwzFIg4vuOoRyfhLzEqIgD4
URjYX7KB6jRiGDwAs0CNILt6Ol9lRNNIexabgILve0122ik0P3byZcKy7KUeVLf9
vpahkW12/C3H4g87z+NIS7pJLdlnQ5OUAvZw6jHv2LqixvaeqLls5HbBaekGH3XI
ihtYGM8+V18A7UQtso9eqKasC7hPfnJW7U08cLFI0yeqZTq2bCG/qpwxKNmnHMvS
g4CW85KZ/AtUyZ+U1CvAiknG67yUPnV6PRlmeW+3YmcqusitGCkcJTBjiEZTLO6m
cjLIfHa9zuGkSWGmYH3k054fygHU/pi1frhr5m9DxNmy0jy64ogTXYzlVGymPYpB
DcufhiHfYgYNYhZOHKmiMu8NNPEVFguSYsH4KKAU+jvhlIqf1yvGPCptYMGh69Qi
4kp89e1eMgz0Hy9G9OQAQKo3pfCrigN1nicWWjdvDDTh7w3QumCKN5JJev1jspOp
yhz/9jRNdns8Mvfim7X+KnPRZAt4/VYKpVSUI+FFKpNGUD1kmUPf5tAmrYq5wzH9
ILPZg2Sl7zmx5nqEPACoA7odD9ZucOHjmFK9ylSk69FMQxSifi7Db9p/R9/sXNF/
Zu+sVONs4DehF6VnLY1UkDB+3IrS7HHa4HKVCqn0DLff3uEbrb0JaRCgWCKOyDHo
wNizwCBoLwFOY8ToRgmjiWxddVO3NYBy6IKaL5905VSBOE3/S/nH/f75id5Fnuk0
qMghnE8DsI9PuLGxuaqlA4j6TMCk9yPidWh6wsfONpfHdxCKw7gttCTwfLheJGRT
HY3oWhhDhb/+qgZ1Z042iYQ9Sulb6KyPCYW/gkLVrEIHOLy7GR9K7Fw3wS3oM9Uo
yBlT0+NPJUmivbplBajn7o9uA1d+5a5NBA+f010HT67GPnYqpK3KxYcRen33/zJl
WrfPwLt3Ak5U8re90GM40VBagG7pH1ojGa9LujND/4HLgtCoENqR1Qw+W3n9T6JL
hMbamnLsdEwENVYAcMUcHJ1+rYYwaR3qcCuU3eNrKaV3oOp8UgdbCZTU5MUAOE5E
CKF8l+kk/xUZYlc7RjSu+QmhxHRPbO7Id8tK3M11yAxKu65EZxhWcsKxvZQlbNsf
xbAmaZcxu72Uk9ZKeKPoUGvzvOZSw9gfXXytkJqDJwo8Li+fCQ2i7m+/AFz5d5td
F3nPTk0aAPcL5FHnnEoTnCZ805fvCcLMKplNBV6eiYJUyGPraM+6J5Nlfi/Cycyf
DP155KJfsBojKHL/o4Ruvt+9fqXkuIcgJBCxwICqy7i6cwHLBB8CJMRU3j+ITaBL
WbiYGpH1t2YtHoqjv1RHzuYldtL1YnTyMVRcVKv2GtfHWCahwFXqhuJCy+E+854q
Ep5utsl1tksvbgJZQ6DwtYKMiIGr3zXnZ5fUprEW4Hb6xanwfwJWN450t3BxfX8q
WAuvN2qO++KkG/ro/GuaAyezgraFhTrzx7BhB+7Bm2ctWY+1aaaL+SkWg1w9KT2j
+EEr2dbJ9wpzxyYVMUR1MAGvPH4ewxMcdgSonQtGNmKtQNw2KosTzMmECt5cPkm7
2tr4mUHtHpIw0UthxSGEC6ZQW/tXrFvY8UWfPASGrWO7mP+tgDKNzAD76vn9E5dn
JqLqAAsxxkCH0iT1yZoAmonluOLaeqOCU/EO8KsffpesCe/zw63cj/Rv1N/xvsaK
UnTeF1JCHfFaeVzel9/4tf3DX3K3VgO67TX2pDYiF5BAXqz/dT9ZPhsc0EIILKuG
bqafvxcKluUGanOW9xemyDjiO8SmZsYJh1t3fDEJKlnTI/w251yKJJJMPPMth+Lu
Hn7iPKlyzSGgcPAQY3kfU1PYCxh76O6ocW7QnvexZDbBSQbU89BOEblQeMKvVUTD
g+ToMYqoB+xFlP0wEcQlYE6h2hurvnrAAG1C5D3gJZ6Z2YThZmQECqQDrr/v9iZ0
1nr+c8k74RkFFcd4FSnErsHbAaEGxyE1l47FOhSbPYSmBzdvZ2kl8mjOyBcwoph3
OqAyx23EbTglkMH1YSxalf2FXVBn/JmYPgPDLQFhvnrX2wIlc77kobs1gr8JHxXt
iXtNXIcMxECOKI5Swto77Xcvt3+p3embfxu0BcT0SS3e5NgLRH0D9Ay/veFRRXcL
FvRZvEpmRLvf7e2UtNwS/bOz89l22ZTCLwNFMVio+jOUrbob38gg1HyYVUYUCzM+
ioH6px/vjjVKdMOF2iJXBh1x2r/amACw2srP3bTDRdAWkcXn7MuofDc8BOt9KeaQ
XbUxheWqugQpq3w6tXhzCAi9DoTIDS4eVyDq8MiOS24Talj9HEJhyFm+JmNK6k6b
b9Lr6YmBZHdqvU0YeU4NcuCCWB58MXdMJ0xx1DGrL9gtINP/ty1zOsEFbgeffi8b
ccLLmw4hORTRdrPPIxdN4OvUApwdyrfqya8PHaj8JQTINeqS/A1HWOQUYgTiQHPW
N9WEoy2Gq2V9XFPCiW1TbRlVEOGnZxkx8RoC17fvb4Pbppaco09lThZJs30nNCiL
PgsB7M23xXUDGlQS3XUlOUZyF+A9jaD32+ttH/Xe9uVifSPGtkrW+b1edEE3IL/x
CK5zveC4Pb2KO1yfx6r+d5Nxhech+IcUnAwqck8qpUrapbVHksVyW0ZL2fRd4v3a
Cmoo3PHoniFXnn2xs4pDs9cbEdXnTdDvwICIj7Hz/tDahHlYTybnsQtetQe+NQ8C
U1l1mT96lmt5TXvlG2suPQW6N8Pm3ywzHbapMjX5azgX6WxmF4ifn61RuVISSm9e
d2k+DnTMWe+rmtzRUlVYMaU26bUsl8zkL45DqViB2LHDQcbKgjBjwKVJDn+Sthxc
wRPjaCJsaEMRU/xu4AYkifVEgqd3D+yJ5yYswh5WRKzsq1CwwjTG9GKh4AHzjUqY
g9CP7srlFMrXoHwgSno0ge+Gdjb3PyIEcoHQ9mAyCMHIb/kJvRXvIGPm15SGN0bG
QVZYVXG4RgsrzPov+tdLvXhXeaPQMS11thi07G+iAYY5VpmVjc89puUNNe3Ms6bG
3I0L1w9ujqYn1RRB3V6ifinm33KDdUQNqj0AHofMujkmf+7Rm5Iumym7940pQv2S
327PUS4LMBEFaHCYNl3HECXZg94mJ6id9Ar9b9nlBzBHEDO/NFl18HfpXQml1RUw
lCCjiPQSQ3JoEH3zwjYm4djeKHwps1Ur9BQ9JW929E/tfPrclAYjj2i4yMKZuP/J
vMWnfKb6RqDDlsaquaqaKekEIgPcZJ7rzzHqpneVL/czC2oeqLL5oE+6RWZaK9be
8gjsHEfgsgvWCSOuz7bYhlT95zwcVrrlw0e8md2VtFPkmVKqPSKBL0f6XfWVYi9F
QofBcGC7GJZaNDDRXs2yTQ/8uK7i6p4sdJE/1q4IrkWKx60iVHQdlprdsaeODLnG
RQ0s6PmxCOWHcu8KTc0Q/opuj3W+3aXFL168nLQHIHOcbSbIYCt2pWMZJ65//B0z
xKdCNQmf1sukB7DeqDVpa2rqiEVaNvi1/ZBtcMcRWUZV7Vs38nnQLMy+xNC5jkjS
8aq5/dTAZ33vDDnlSApoB9dN41S8TmyjbP4TTQ1NJm9NnN/+714GzZ4hTZZZyqvV
ud6h8npbsprHyPAYubISikuJFVZIg+fqFobtZsqntp27HGM/6MeZnniH9XGHjvix
uWlNNAWUtZ/SscHNgo5klPD3pk9LJ7dJxJQapJiupPEyxOsK4Cy6Lv3xI8teYm7W
EewQHkLi/NOfKA2WO/zMhNkU1S+Z7yK/SrOV5mx9h7efr3stnrDp2XWQn4du8K0N
eFthQ5YGON3zF4vek9uiq9IqXCIpSG9y+8c5l0PzV1ssmebmMVQhij+CRFzWKP/a
KZRJUKVzvX56D7VBbUnYvGNZy3b/imOl2202X8SKJ6R9Lwz/GBMLeDqhvN4MBCQd
LCJ/E2LOTQ/+AVE6VxNDKO+3rvsNvRi6/izyMdBxAJfZzr3LvkAY+zfY9qLy1Ytm
wu0bJTDm61ybQvYFitpyAybUBMrdd7qtiz7oGINmmwxuzSNYdGe9b9Q7xwqi5eSR
744+C+7L5mA+rClZNNwtuIB2cKUKp/KfFtojrnDs28jzkXA4bYFaso4dMV596srC
ghN2UKBiL5GHrcrq+Nz+nAFmO0w2+OYofq8oM2qodidE/2tbXKkVSjYV+CtWgk/K
nM8dor71AEs13sEfzVg82bgONn+399xjbwA6Rsy01YCFWXJfqy5V3n6ZJznhpuG8
o1uvy4L8o/70FEVfo7rhy+7X0sI2pldicU4sWp8urwxLq/kpLw1NVR8t8KboYIXe
WDYFhgZ/2V6uU6iKNnBg5SQ5PQFZ/lZgwN/reYpo8D0aExSMBhuYmjbsYXXc8vKf
OHYVRko9YaAT6K8sXBFs/dSb/siOJ66MvEcl5R0OEli2oGFffvnO/0GRHlxoooUZ
WwsKhaKxFoEMNSn9bvh2aczwhEI3xxRTGTQtNCJM5nfUyichZHK4nLDfXAjsCMCo
rhj//hzQkDCN8L6ydVdTn+ESTNoM3IvY9Plqi7Na622Vej1UFscc/aAfSZS5n4ak
px0aDC3NxsOSyIFs2nxkHplUPAeBZ708eUXlmNEAqcvmalknRHNu9RdJxw4r93QC
mhL5EGiluhzXTwCfmxnd/Cv9aMMSMPnLi5stG6Mz8sFGRcRc95oy8RIBJyyu5/of
VaDLVY1XNstNZbsR+WV47O/UlfqQZdm9D2hnggg7hxzTEk9imTOm6xcmE95gdtX3
328R4eOhl0Vny5eRbsyzpEE4cX6ziDfkJy4X61Wp3yICd6r0g+nfgyl7BrBPV+pW
6LPgEXfHquTMDomD1Fz+3tocRtIUWiASUCpjBQe6SWNZxQJyb9i2eIqoqrSPo3pa
D/P3USd3y2vbHkHoBWn+Ai5AQr/Gd+3LmRv4NfbVUkLxmk0SrRrWPnRz9tJBgYeq
GaUMoBEuW32weM/4lQLHT2MJ5o3rcEI5gx3PNIK/h3KbtyOlTiI1KbYnE0Sjpuxd
TF4tVKjerRaxBQLAjc1WeThQdfrsYoeD19wxmUsUV+xspJf8Nx2Y9GG6TTADS4o+
CDDo+7xN+bQyj/iNslblOsVwvTS1X85pJoIASNy2bSr2UgRyTi0gUjSDiaZSGFou
ph3/mdeXMM5hObPjXuYXgZD6KfQNWz2IoRufCtjNlCUsZbdurpdM1bi8OLcsfBPU
vMFbnnT9ARuPq6iHvLYI8WJRGkeRvMCWrR5a/nPvHbXvGIuOOV3NCn30vHOODe/g
8/FS9lJa0zFiblEtr40b6X6h7qO28EjnB3mN5ribzFMq+iHSS3QAJ7lwW36ho9Ik
oIBtCM1rYjTX2TrUKtxR0RhpmOMenVgT/qlm7sToelZ11DbPfNYD7yS7b1PMnX54
umL383xidPGXbjhmv5yLeIkF9hauxJ9i+5uhsDcC/NrWvvzOBqr25jQMPqHfCsOx
Yt2tXDLTuPhltbnT3NJxpJ8t520qrhD2w6AhLY0Cyu+HUbsPQ8HLKIlpZ6GUSoOy
5WEaPd8i0akal3vrJNV8B/Dn6PIBj2uANlSN1p4hLh2eg4rfBHVUgpFkjkPlfamg
CV2HgKPAOlPN9QIgk/cK7w5eyy21YmWMrqMTfhZDI2nNYPj5rcO9jJCQBTepgyq4
geOy8aRndQR//et/RcmbEBOqWDIf/MuWLKHNrFbFL1dU1fCAQBqJZCHhjNzgkiVv
dT2OEYPbLBXhob8+Nz2Xjd0IrEFe3IrRSLQZlquaNCGTPBXTBsJmj6jHae9TxN9c
Pv+SQF5uZqpqbzkM1VItsrOXp/6czXcVaXFKT0SHErUt/3Zkv57YUD7nROx6KRCu
f/3DpksCbTeGwi9Vj/Ms+F9H0k0+/KCbk07CR4yX5rPH2vIX8kNoFDVY7GIPlX0/
Nkcw+ROp62gNPmTFYNdqlWuKRy86fYZL6tvZS/UHtjsIMGZBTzAWgce0bj+vLkMn
+oo30Tw/EeUSrLGjLs4IHLloNPaPLDxc97QyCuk0bgeRIulesbvgDE1MDvrr7cXR
P1BS2yxEHBmV0tXMSqh7MJGq7HBzFgh9mM7gL29AevIFeyN4XQ67rLrW4qYq0Z/V
SKIpn36CxraR67Kh/omSwmdMYzEqlWcOmge6vNyGZZ/FEEDnq3c2gCRe3O7X12Hk
JsXs9SePuYnSLotRb+SghAURu/zzGJFqmdnTgP3YMyqs5Y9t8NUSxIJe8acSEChS
xHnqEb3dCbkcdFirsgmFKSGzsMRwSG3AHKoSjRHmuJupgLsCiBS7/bkZx2k0Qr5R
Fx2pFPSnuabIMAUN2qTi53kyUW7aUsky4hqtOMcMXf2GNiGnBRv5KtYu2D5nl+2z
MiTVWDhU89hVQoEgdlJOEVcIwLHFb/Ij25cnWRlmC0uknY+6PLPPaVJWhnwxzUXZ
NfZYd2PfXZQRrsb/m574RhXpX7bk1EqKV6V/Rm21k2XT/WcAIF9jsBWe9GBVa4Ss
yHKcEH8KXwcSQ/shbI2WLBY+itUuxnr9N4ENJnNyylymj9FjPU6ErNCxZz68aVIz
MlL3vdLOrr/cTeyH0Y4iMrEysekVM7trfgrnp/nKJ5Q/osYuKFimzSRnvFlFyG9H
hHiSyCeF5fMAydc1bKLsY9OKNQT/chxgnUjpJhYc9tqeuCTQlSleVp9ZM9IDnk3I
tdOxtie/i9lmTugiWQWW75FSqkPRDlWkuc7pmSx2E/DHoK8Mhwwu+oMxOBUMDqHt
0twbcxu/1DZT0sgmM5/dx+8YgsUy3gtj5ljHsB13w0fOnVGNLdZQZ9Hzp2qP5XnT
fH2Xz2qiLljazkFLXRrIHj/F4aEC9OyRU41smr9PyjiZpvFPbfo1oMTp71d3JE6c
wHl+LSavN8bFcowC04N4ZF8H9i7wtNSUq8dIhVTVYd7R0PAPdXtCbh/DAbdxlzMp
JRN+yi0RUwWhkvqI/kgQcp1+tMCg5t2bk5y+OupLizgiRHCkDG25QBmsEIm6oEsM
wb9cet00RJEv8acVAP2V+TmbO0whDsUPJ8+hoe2i4k1R/optzCzFOCD6hLPq7mNV
O0QbZq+jiOK3WQ2nc7LCfjBzgUHqUBtH8artV+LMshmUGUmy3GCMnPV8nSK50V73
mS5xemWgp4fS8dRabR8RlglKFE56Ba0zFOgGkzD6IAYhFWtG51xTh/pzmU/uZE5l
QTa2sLP/KVOJKlLQugfXbRMUf5aMzUDtfly+KPswsVNjEbsx1C2d+3hvAJnWSKwx
HwAZr6KIZwhKslKy6N9jArHUVuW4SthnKjVZdVxOs6EytPq1DcAlEtIAwZfH33vI
MgeohZ/IONixZNXtW0+Ho+qTgXTkCwuWdTjvu4O1rkDUPihDiF6gUFaUwSnOmIrL
D9utQLjwNpNwzqQ0Jv4SGHS+f63OTGvE9CvSgWLp+dgDByDSXCxkRDXVCRC3qe/z
1i2crsDZVRzUcqdVVlxS7E9So5uQu+OKQyJ2+DZcKogX7OIWaFsYNB2nUm8kYyHz
hkzxAL/qAjG28BnuhDb4BnXhl9jrs3x21+tAi/LdVNgE4GeUaqveYVvGUB63GWBV
oeGoCQfoc7f4wWslf4lwVwuDM8JuYdjKeTeZ6p5z2CP77UcjRlYsqApggqaAesio
182fZKks1oxvpo99J6040pVjUjV5CFdf5uitvRSNDTY/U88MKiKObbK98Qa8MAPT
OMC9SEO3PQOHJBpxEVBmVMhk0fBmxmUjWiPGQPvBZf+JUgWgKF0fJRW8YWhulkIr
gpvXU3hKKyI0y9g86ODAvADc+kk/nnxNsnYtsVtn0tCaLptc5baUmQ9pt1j+YJMp
4HzBJ4h8i0epPoO2y8SzzGbSb/btOE6pP6p22qsakXfMAw4H3kNqmg8/LGwBA9ta
Rxh9rKv1kTRnPta1GCb/7XzXj3oryn3wZ5NH4q7EXY6CvZUIppXatiibYu5pm521
17mBJBYneXNHPT/vkmJZRmC3LjYV2yHnHxr5aM3PNWDKm978X4KOf6bl8cGRYWUp
V0r2hsMBoNKfAQ/CpsugeXYn3NoMQY5p+vNpe/pKD8JKuFP5U4FugkogQVZX3Vmz
NFQMwdrepMEQTXoZHHYpjTH5VlEBmp0+qrXwGkQk3+q0KYseNzk0xegB6mWUvGfv
I/Sx+Eg88b1OyyjfgoKz3rwK8HgqFZ/Mkke9OE+RTYhQSGy1zlTh6L3V/k8FveDn
9Z1RUB8KHu35OFTtLHn80+39Ou05QFy4uOTDMmL6EIdbeCULGzN1Btx07f/pJYbg
YPeriG172QLnRslzMBQ4FZDrcFTFRGInf9DBtzDjLyI/tU2u+x0YEjwZ8zDyKtnC
s7dODL90IMu12kmEonYTeDHR2Oq0msif0L9SC5B1uOBtsVFBksZjJf3CSEAlv4DP
YbFfzQXKbDEW/4G3WkrYj3CnbDUVlh41qDvhqrI57bv9Vl7PMFG0y/5gp0OPESxB
+1CCeBKqOVsRU7VomdHTDwlXnB2fikVFiMta55s0rWO2RE6+omA7esVweRsCBtj3
Va8HSNoYbcrPW4LfoPyFGDIQBV+J6Xg1SCa8PtgLfizZ6yLeZGWrKcz0s2mjU3ra
HuvBt08VuVcUJjQUHV7UMMR6rhyvyikN6E6ZA1wti7aH0t/9CEXfwmxagAfzuzk2
OtGaL98jJw54Th57GyT52BRhWgbwQPxNSucRS3nTuSb/s9SFSWC0ney0cnHWqBId
CLXNk1oCEkrknsiNJhV+NFlll+I+QFz6klzCosYG+JMcno8++/fXb107zwnQnaV2
upclAz2P6jQjiv0UGStQjmhRCp+3WXnwyfxiT0kfECzn/KklKm4+alJ9pjB43Zuu
zE3ExFrOBEyhBhrxZ1C/U8dlR59n5Mcq8XZvK7jeQ2H44u4Y/+QBQ+kRqzuDDnes
CfKlQ/TsBbTHu5Bbn5ysxk6q3kqLDI/uK6Yc9B7js84+mwL9MUzID1L1HYUj/kfZ
usTjExnophRWzicdRSqeTWPy6iWEnl0iMkJNzzgScrNki75f5w/eyNVIP3Wm91Jv
4B8JXz49U58Q2yJclEWUsvLoc2jeWKqvSvzPU8qCEIqt6a4MCKSQdOu2wTHSPrGR
nhzykQ3GEZrnzU3EW7cptEYcPwXhz+vojSmcnK+CnyzurIJktCtIAesKOLhoNCOJ
MsrauN4VDGi13d51XAvHjKYopWiUKS2iX9Mu/HQvvTK5kMDG9dd5UTzekbfPPKAV
ZRebhOQygc68uwlgo9hS40qz3jvyJOyyyU0stMplLD1ON1oLqPJKwxFspISMKl5R
ydpisnC5VL2Z3gPC9jloKGDrIgiS8pTupHUBNrhb/p8rz1PS6wPcj5gxsWphoVwe
boz+Y4/XLrr0g31CmvgSNvYQ9c+WDOxYB6vRI83N6WP4rv2Z6wrHw2IW/9b97GVq
dhQoPi2NeuBoCgGQ/QhM3jhYj5vsi0l54wPATeORg12hhIum9S45JIPKapXtfSB0
e3c/WWsqi2RXHmURWS7GsiHvmNmmwTnBnS/eRmXx4Yf+koJfu4kC7nTZx3jw+1a+
Y2VAMRVRhRD8MfalCS+hi1jNMOp6sR9M1fNtKpeR5hbQwQYfBRYLVKCsWIJaJxET
4vVqnAvus9ZALOFPxJRaly+I1vSXeHsk6GrN9QXopMPx10T4H4BP7JCBdhtBPdBv
YLiuS9nkQWv1ecXrqy+n7RydCkb112o8QMXNbD1LbxJSw+Npbz5DncezK/VjACzh
eXvyOJkfFYMcEvzqXD6ZtuDAGlGX341M1LIiecUFgJnG8DObrSP2y+oW935AWYLv
5b1bJ00KIqf9p2RHBiBaArsB1F5FZ/gQAidpUiYBNUbPUkSfBDdL2vh+RYHfDS6r
RxXgQwpPbfPf1mrJQ2baTsBnL+wpKz88iA/wtkSZhxmkJA0jiV5U/+UlbMSVue8V
VkwyWTLwgdNdP1F+NNtcczwz/ahQWG+Um4J6tGG5HLt9PMxyYeHNeWcKKyZv+6zk
duBVAMK2WCfCsdAps5sF7bVanMDv00B5q2eV3EjUcuuqxxwq54eXXVmzCOnsRCls
Hdzdtk54Z+oXGDZ38joPYwIaLkey4bB4ZzYo//N1oJoeO5/DIy/gFaezCaD7hdGn
GtCHYATVQypCLkmjQfQlqz55jMm4YKBCoGnNoTEKiKdE+eXh7zfIXpZ/GCHCqh14
ptUoZOoNVMYZ1onMpejUZVkxR+FDy064Wr2LLalIUdlkMpvXcWUEPUwR8gPpDQZM
wETwSFcvXUZ8QNiznVBN+J7DVRdO1E9xfgxoR0u7f8knTnzbttC3EYR5jtdRBjTQ
neAvC+/93Ha5ykmum2qXJPPfjWls3KIa0/eUw75TvRG7eGOfzIrDJ7C4QwPgqR5X
QRN3G9wl9Hs/V6fkpmZ8q+wfPysemdLOC4L4VrABTQHQl9CakXB+bOYqdFrWEPy/
kOvwnk+yr2LWd922s757SHThehoNyQ21N4RUFsGrWQaIbMh9ShIw63lHMpuZEhvB
KIrKtPC2nJb+zgeTfRCalCZNF8yXnAUd2m+oWJwsdtNuYeyGAPM2GCh+UT6oAx0G
vu2HvI2f0ozEX4GXs9EHdLyRpwGoiqVLhvyXWAW0PRza/5pImf++x75YgP28rRpy
Mk1N2t9jjIpgfwLJL1HxwPF6jRZlinDM5YtMbUQZNoTAxSuJjInkygx3GwBbRO0D
da5JcBzupcAr525BD35dawRC1J4Jr0lWVOeM2b6StZWp3JLx+X9Nl9D6/IUsejA4
Pbx1MArTf2g2WFMuJ7MLafFzwFdLxHCARgluy3GsEFqN4WIqJY8qdRclQYUEWhdX
XsgGRiPPgfBxPb2wzjxeh8eBYWepOv8fmaJEhU4qi//+mqyrANOmLyQjPNTdEnCQ
Wyy1A5rHQrMkyiPCbhzljvSyrC+XGrIaR0HHvrQDAELAEjk/qGrMhBJCt3JwZFVj
kBwfKLkvbrb2nkXIWQ52TtEG0rQ7m2WHJfAjEueW3FdQwwqP2y/d+DrIx39RUGVZ
DE/uihN28fBQDBlDoZeG9rvjEikby3r6WtcBa7GTnEnw8O7r5o964AVSb1qtwyDS
shXsmmNF6TDW9ogvIZhyCkpePXjZunLlNuy1ztTSiLLhXjxoISoxVLXjgoiDtBjk
clqbWOLv8XeZu+2AG4eXP7mmrOmuzPHU4zOeSqhHhsSqsnbetJwMhiUBGmek0+8S
aq37G7nfqmijbQJhl0UsxCMEhDD4o6eAA5xTOW9PpbYl388YCqB+7B7Yme/L+w3f
Ibvnsazvhs4Zk390ruzI/AndHif2WvP44YBlkcxIRLchSI0UEHRnBxRgL5URFd+C
5lCqUv7SXCI2yWEeZWzKYb/AKR33hmt839ou4Ks4hPKHbbATCnjpjdHppPAtstRj
XI6BgE94M6Y/WwMac/Zc+Y0XjVVGB+xC7FKMLdU9omjY0Sf94iPUnbnoMaWHvhb6
KwR/vvungkFtJWsUSRtxVWgIT+F/NhEBHzuH11iyo2MgTWUNyvgIW2g3RGtz1SyA
L9MSLM77KgVKcLXOoZTSC1VA1MHiCCRcuft+sQsRl2SnOMXCZRALboGjA9EirWXl
whQU8lLGaM614QtzIh+ZtcVv6Nk8yEQInPv92aIV5/ok9Be/BGhVHs6EPUEZkXqn
ygXMfl8siiaHyhP+ntw2ESsOxKiqnPHdoqO56J8IUm8fFcD3nynroB/74RLbL9QH
jy6sld0WkE2p/MJ9naA68NAlSGKvyBMHyHUQs0lcxKOxakTsjvSxlsO2HkQXBM/6
W6YbP/SSXM0Yo4RN421M7Na4Fq838AywPm7a4nbB7vUzAW88rN0lQa+qqzVrM6B5
xiq3ykTknfKB4j4UxpLfppx/PC5M858bk2UwygBq5tq5Iu/Sd1rWOQUxLdpzKpqP
+XP6+o9I5Uz5kcSKjR/HbgbaIMi6SZHGLdRBKNv9kcz54ayyzxLUdbsHwr/bP/IL
FWzsxY9IEvaeCqlDZ61gg+QEt2oXZ5xdwbue1W2K7JUdP+jET7pWGlsCG/X90Szp
jCFsU+aIMX7XyUkOpJSt4uNszv8dHIq4C3nmB2ndoyjEIlUMMHdv6lNbP6USradN
EAGoJfopegj/dfFy9UaeYUZnjgfc3rlSw+njiHNzsyzsW0E4mtZ/D3ogX9i5BYsS
XNu4sKUbPyw3m3+nXAHY49rooOhv69RUDEcamtHWg0CDQfxhp3NXfIdyVLkmdbyS
DWDT24O5qBOeRtHqfWOWMFORFsm+Fv4pXwLll9gqOwyYCgHS2sfupiNZfvbDzV6L
CVa6axP4ISS6OK4o3sWDg268RA0HgOsyQnBQP3nqLTq5dWDAc2Gl79QeWhFHNBpE
qinPnFc/mhK62JFRx54K4/MdAax0zu3CZeRJCUSBI/lQGHQIsePyv7Ibw9inxtKY
Y3MgoVTEHP/PRir8LoooSD/OQEA1wv7tIFPO/xP/YVciaDAHJ24VwrCeruZSaIBG
4cC0UAYVSJgpp2eDVjRQdRkdfYozf+7uPkpjCud/Ayyd8pvobkcjNJ/gSXeyLEuc
SnXoE7zWebxNIyUZExVYapSrqlMGEp31zDlpLG4byMfWlM0/Lc0i0QGJQstX/Via
FHV4rGK+U4ikp4bpwHy3d7vQHCFIN+0CDXgjubU1qBCqTfjPmgjQ9OFJKpqODgfv
F28rRughJqEaqkS2M4oT1+c0VqIl9+UkXrN5KFMgsBc4RksCVhOMBhlavSfhVjB4
LFphJ/Pty+2pFPjCasYrRiFwKrKDDTAjEC9hgwSs41TjdQhMXQ59DyaUUYRAYRPq
nU3daUUsw7n20rgbniwowrBS0cN52bU6bVh1wMUQwNRgB1/fdjVJOYMozbLZp38c
3H8S+gt1LekXGz/CBpSVmW9x888V39xjv4yR85MHIp+c0oKnjZHQR/WtXebVsvvD
mrIMrZ5tI9PVO2wU8TDDicZzQrJbCf641oYRCF3gmI+LQkD2tgoVnvGN8ZCRIxuh
nTqNcfAjQnU090FDehvRnFXAmHtelGZaIvHFHJ4nHjj2SlxjPC8+BHlOBQfteirP
eXx0zM1eUpKVZRV1KN7THRIe6XA2bwjnj+ZuGqGrj4M05O+yoUA5M2FPDjGgwuUH
QEDyKJ3/aQv03wOTATN3K5xxFnQpUr0MQm3j+Uyx1D8zIeAFewQUBVgZc07VrKLk
Q7FinXMds7mm9UP5aVxeSN6SSvcfPwNjZ/8fDkcydGuGZOHvwDCvrFvvNwdnEhsL
U4PbAnIFMv462+i9FhoWP+0Ii8cp5+Vv/jMLaeTtWjKdUEiDVJHmvdLgEbPw/MFk
byGPH8JtgJh2qsWjWGAI7Ilk/mhFHrn/P1lK1e2ae/9N2BguQJV6ALMZGROk+7i5
nA3Ku7RGIRFKIccbQHFAF/EoG2UcGZs8NwytdDIl5MDuoZyievUJF8Ldnsbkf6TZ
nF5pqMz5KtNRA7buULjiFMb1vLyuZ4rrBpWpQzoezfnQzUHURLpQm0prW76zJl5C
azFWbKQdLCAXaY0PNuMjxXXLCzGyzwOJTtD9U4MUDBHFF6UeflCJGHMeQOk/e/di
P04CY2lbpkAbPtRF1/0KB0tJJN1MlHF8bH31FYG7ywWv1+yOiOB95VPCxTk9z9T+
B5NN96a2zSTOxhrFScWUQ3SBFY5bDSywRR2sDghQqnnsEA9G3M3dw5F9jDmFjGll
AtPV0QUnEm+TGL7Ye7nj47jFZCQrkewI3alwDIKQyFiBhFRhRljKNB+gX/CT+f9y
AXXMVWThaIDrPUSMCUCTo2EPTJxJtx1N/T8KdWgq7veiT0+1Mh+6qvkJrANbgZyn
BCeHW9w0CPzUgVgsEeRJuwXa5jLlVuM313fwbEJ5PwCHKNAtJzpYUJwvXR/UsSid
LvRnndxPLBEA9NGB9Jxndvb2R1D2PIPt/K6jxRvQaoxshu9wh5N3wFXkDH911uAH
hDNkPYS/ivZvyL/zCOUdHSL3hrhlxkqdurPDZWSmjYq39CMVIBodoAngelbCyipq
8vvtZ0v330eBEvsEPeZIQW2+CAYkdJalqDWlbofw12ClOzRd6I7T0yqvl8T6TKZO
XtkiwvUFTUX3GVAqj3A9rPjYlpF/OKyELhgj2XhUKLaaFbDHyyV1YJCx70OygPCQ
`pragma protect end_protected
