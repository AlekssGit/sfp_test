`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
erWNKsjV0rKN/p1Vj623rARDpqyVB+6jCb0w+MoSd49FXT6qjGwFYsQIYbw3S6Um
Ri5p4dAGF0YllWOqDz2cN7ZukuQq5odnqN9l870+GjRicFzq17pC+8ttIpVUsTS+
VinrOUT5RuRfZJU5lzSzM+kiwK4TdcdnhJDl7Ydhk18=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 5680), data_block
E3VUeUFkO7scf8Yd7YykF+BHvyRAQzcDEhbUcBjelV8GzfEf58WaZLQWUA2BejH6
W9TfewVwEERJ+g1PTyoinh1Sz2LEbx79oN/Hy+IunNDQk+fasXYFWaESJ4XRM1BY
ZcNwdjTq9uW45dgDC4KqfBb/0U6BKa9hQPMqY5//TiWDJ3eJzn9ZDOM3JOUHvfIm
wsSjdERhLaSdfUgQQtDWqnQsZL51kooFPMaEkyx+MYnlLOemFw8B44YBMaJMgTjl
oJ3HWfgxIac3DDGKEidJTdVoInGS1csIhnttp96EPzYapPLSouiUsXprwle5D785
Qe+iwgLn53wpoyk9DJOTy92IEE4IctwKLoTilg+zT5ZrHrF6WleU5SbcMYRyezGM
xGwbxNV37WG33fWPKG2tTrqQzU1Vkj1ocil+VaZg2SGkC9qdlu5wGVce9Oka5tKG
hMzrv8BuL40TMXVWCpTC0FhV8PnhjVUxX+cawMx5MeyxS17AuermqvGBJgyhFm8T
Ahfa3b4WzPKP/kSWSSMN6FXf6S65URrxTfmdlormAKvfdXLWed6I7l1q68FcezKL
1uIn9xkIHbISggPZ+NZoOufWOw9WveyZXJHVMrbIw+9dFNgBpz1LK83Nk1LX3L9N
wnNeSnOoKf3VEQL/QFrO3XQKnBGxHVeu3ld0L1K8Yp624auUpW1rSlM8p0uJhssC
R9tJjOkeol7LlXXaZ4FRY7+4sEGO/fforeYgBfqICl8VZJA0vBx9qbuERVE3dYQI
BM9x7z7nznllCScfmrShRU+jwnqvsGPWA0pqwnVV0+y2YmdBUWf5R8putHSsdI5h
8z6Ms0UeLLm0M5eTH17T7TixGOChynXc6xKIPkOFQue+wN5COWPxAwMfBkoazT89
reVz4150lsPBzFbcbq3ogrsQ2VchkxgHds+ntRuOnAO/I9RoDMr4HgWt4PUCRazT
ErpFYggoKzmGJTL9RUZPBPWiV5FwM+vK5Nb44aPsorQI7BVdoxvA+6CZ6SQyP56C
GV7/vC9t42xmHIJoTEb0DOyIHxBBZGfrveh+WJ9sdwATVUmjdufwY1u0G3J/FKSu
N7oBNMnvPtCAO6XmfCtLh3JmVR345HYsQvGurSg+MCnzOMj+fHFQ9/jPFFNxmwYO
fZZuR3OPh2Kd4HV5qfrCmJZ2LnMsJINLRcjnOrErNkxZDvgUBN9lxKNjxliIMOMG
bMjGYxr1SZNq64oJgZtnn+zrQ1VILQIWX5f3YXu2qb9lqqwtIJDv7Xe9Vmpq24Me
5JkAsEwNvz9OavfDAICp9o8ku2aqOkSn8YxLB5IM4JpUx87RxJ6ErJI9G+J1mAEZ
FoMfdwh8q5RDsFmQvqZDLyK+yyx44YM1cQRBJT5R1kCZOcNCoG45vjSrFrxMJCDi
hQWZQh9nt41MJuMOnFyAXVnYAWCUF4bWPtaVyuZnYgL1rJ4ssg7Y8lir8e5kWi3c
Ie5HyO8pwvJuWAwa90P88/Mhx0B0hkFHXFg8q5qE3fx3SBEgAOQ/0dYo8QCzlBYC
LhXevtXfMWz0LIKcIThxSIYsOa+kkBfgSlWFNDYdwBW7y4TBoe7VN2KNx5iAVZ47
n6K0eFAFrlUeLFG61C2tnjHXpy9Us6tuF6Yf88KSl6IzvXf0Bs3UfgI5us8kGAWF
XHme8C3l/aMuZiDoRvJKm0Y3GCANmQUP8b4shTJ4P8NE7mAKQ6LqI4MyhLrhNQAp
RUJPXKpehx0UUevXpyGowdLZZ+vJf52K+qhW5ux3M6iLe5HyWR6ZF/0sOaaEuzsu
z3u23J7Z3wGBoh8DLC+nLUV7L//Yj488iMYNgy5bkz6aZi0sxj1n3h5sJMadVJQ+
mTOZBEOS9V5MMyrCv/mQzrW/OjPPYisA/bOWe61z+tVNfeFUUV7Em4YrY0xbZIg+
9jZ03FCClASw9GuYbTXJMRobhJLbp1gu0kyjfp/VAz28rfDo3vvw1Mxk7xOPfzeH
L7ywSBy8MsMtW2o6uWJoMaNaBVxiadVEO9nMwhhr7V4YY1HsWnjaaHyZjd3YDzDd
diSJ0Nno7+c9YTrT5syM7o7fyARITNi1GfPICAi10Wg0kSyukFQr8zmYonqV1l6I
pH82BHaYMOu6oPtPjjMs9Z3VK8xjfckg1oudKSUBZpJTMKW4PCJdXka3T3FsBeXu
PUuPLytrtwp6VLTLEMXcmWBQYY0wfFmtFrDn4Eum72ctEgi886bG78L6jPOdAObO
z2CrbQDFLBfklS9x9LV+R0Azx2s9HhuCcd55j7dJDe+7hWVI7dRnDeLLNNxUxT2f
Hk4OeKWxJSeo+aeQrJmBQz7siSboHuC8gvD+ilA/3hMrjDDgGsqUulkxr/40OhNX
LL7VdeYWcqx3gFnRv64erqPRgdZiYRgUvJG4lS5h1TUqMB6mOgPWaujaBV29crRE
nJ6zMEauWI0vEVv3tY3cmnuVgki5SCq05Q6BM+IrzaWzUJfiXmko0155J7QqFGGi
nFHlbFe8yWgfVXHM4Uukek0WAaf1lP2Fn90JUurniP21ktLcroypfZP2P3hhG7B9
xIyG8i4baCjdVxxX9uySSrw5PKsd65HnLUg4iA3Zv4YLpttvKCpSmgypQhn9oi97
sQGhkx8asfdZlUEuHVXAzbY6ANaE/qM2s30Si/nP5MZzlxpWDlHpc3su0cAZfbnz
DuZqNfjrJnhAhetM3KoY6BWVJ2xDBqxQUg890lJlkKrlbcZUPyPiph4bA2Iq4vwv
yLbq6RqSY2i1yHr0pppbVYdIkWg4N8E4j+pMVdDTftP4FMrlS72+wTG/1J2cDiZG
+77YMnOrI1jSRk5Y9rkI/OquQm8nm4mtGUM/YUxxGs22g3XYV0PVJCqFgmG7XPj7
ies1OMlNb0Uj17BXgFrc5DjqFWKl0UwYd7rdLnTsTRsYBVkNHsUpzh8D9HESx1ib
680aJVw/hNDLCAOhmgkhBWrpdqWUgdsDh6EwiN8ublTgJQyJ/6hf2RZfhzeJMApg
F9VicDdNFhjIQMLsdGwOzZulgnbFtoq046tNDc7yoieEjHs9vNDRde/BfhbJEeo7
UxGEBy1AVK+YQE7y8urA/QzHgamclklKvRo6X9RYRguChfdXFqsbXnPAD8EvUCTi
lYe3cUAB4GR0i7nSBLYm55XTG3R5SIp9yNPoTUuvuLDzpxxNgSvxiXghwFmiz+LS
JTzdINsY/wDM2CFOaMeKFNtDL3pJJWtsAf8n/dxzGFNSbl7mTTmM6eA6mrAZiXO0
A9pUruHaWEfKuVheAZKKKLZsYhzla8aqq+1sdouYUGZBL7cA7QxiuWw3ZZoWOzYM
z9f/dBGRmMIzLBkxowgesgBeis/4eTLE3bCGFjC54ENnPPRhe8+CTqPE9GIlVA6/
KjgM7jJkDGBqUbWyPOLCYF9C+MfGmlDGzvqMf4DJDGpgD3DP0EAMNss+I/8YfqCO
mQim8r7iDwZXUCVQRh+crKJvAnGhBWoUUnqT67aAEN7x+kznuHHYNDTioMvQbwFH
ajyMFMk3vl5Jj16HGJIf8x/gLPw0ocC+JnBV2N2gm9J2YlFgNKiU7OMm2T7ETbch
q2BOZeITxsCI7GzeO459YADx7zIhEQjF10BjKQ7Af9mtNJE/19+tikZ521QC41hG
sWkXtgdNXpR/h1ivPqmCsTpwXDLemCILaJOKDzh1aJZoY22e6jmrwtzscaaLUU6W
leYaV8RDleFLpplLTnJp1dShpRmFT0iA00udTSo1AwbtkjY41g6nR8U2ADbCyf6I
IPBYvgq/xgiKxX7QBdO9ziTx35tEY1oF3kB45NyXeEm2SbHwftxtu9yPh2yLiUao
6Dg2/nSdK1zbfxM5zZpvoASkHdFlVMcqPYgm9q3eRcsxgPu6ydhqjvsRbgUX9e1n
lgutNBpg6SnL+5Zs+dT1GQET1PonvNCavkdfrlFdbVehfRxZS9M99BJnfNUsRyfF
E1q3g+Pcf08P8tLXcgU+0KXCD+GfzrTjDvvwYKQ2rG0DH0A8Ap0ql1N1sN8U1tx4
+AgWPxR5ANdWToW2Dhn68oNnF7heXbu6RKuN5BYS9NG1q+ep0oAY9Q0ZO0y0ZNbe
uXwWAKp6b0BANV/Mw22eYRj1T68A/tRI9ld8Kv3jk9yaw/wI+u4QZV8h/9zh0O5/
wvRkQXWirzJUkcER/pvLGvlILs+tJXLPhHBv+9iRdjOtYDjbbNcc01zoH7pp+NYH
O0uh42mol6MbNCJcBakuTW2EgmewIyTDe66JK1W/8XvJQHQiHmg6/IgzzVANLwl9
QL2vtVkDHKgYa561nsVNdXO1J/+TecXiYZqunkmIcunOWx8eDkto6UZc8H9Ny+v4
PaCFm7LW8C4hkMzFYmGONYSimd/vtukDjhY1LDkuWy7TLnmyqXTYdrj9o6C+gmTT
yn5+r8oyPuX5ZFIwQ1HbhAGv42UrE6NavAIYxUZQCufmG8SVkxnz2FRVFe0zgL0r
n4nrinIlTNN3mTUW4pGZXC60at+RT812Q7FqdtsNiISJsGgQp6RGjnP5UtIm0fEt
Y7gEM5sw+rAZ/e2UDHwQMiq2cmIHHPEOfjkH5rvfcBcjdTPdkTyKeL89jNjwepAY
mA2fRiEj5UPiEiayPyY9MwLrwscb5I99laQ+x4WsMVlHWe5tfl77MAzzyKezFMYS
f4FivudU+xfSUWGsHsUgmuXoP6ZLuDYpOT9YFD923g4aQsbDm+4YAHcKs8Fy1l9r
8ueCIraUdRoh/PG5wVsYSxVy59evw2OEnNFJPQKZa4BxnDzoc/cIM3d1aeINGOpu
Bp01XXBB7GVBJGfGugwE7qYu6SeG93TXXkFBykWshmCYHmwS/ZASG3JeN2A4UlJ/
1I/1N11QqtfGGAMd9kbYBxnS9mi6lM6ES65gjWsG8e7SjyuOhTCpkqfcPXwNIam4
gsditE0OJDetEKjZ5dlm+/SMPBExyZnDFE0n8QU+3inVbDLg9K+6k5BwGpMamXbe
X7Vrwd5PtCYJ/Ao1c2iZ2QftfP+dzBpTMY7By1DHDP0SwRTagpcGcXPMqKUCCzSE
/lvlwZ0cXPFzmyFcawQ8JXL14t2sOJPmG6XSNVJKAHekNR1X9hVb6tCtzD1UvYho
ZKAnSIuz88t/rL/EyZLhDkc0njuCjQlv1Cas7C30PjsAZYF/Tg9VVponGMutKs31
CuGJQcy1gexcbf5I7caORKVp0h+bdRQKruBjBuXIS7X88WI2c3zQRJVTHEjgH4jb
Cypz+VzDUlimPy5jVIt/nNiY/hJb3e6XrTTB2X4x4OSFGI/X7KJZTL8tFueY29y3
ra5qj/q7+qM519NAZjxm9H4RoxQHNleUjpLpZn7XbrWrdZ6VXjVaEKEQH+oMhj9R
/1Vh+BCCvlznoBKlnbr020h8zPifeOF6LOYbqqjCJqLIx6CH+Pn3XrQDYqTMowc/
9dUBNrxu5ypP258VvTf4xuwM/F5EVuhmVvPJ0XoTOBRgEklHXJ70c2a4ijcMHahg
LCCqEPA39Na7/OEPncRl+GveoS3BWTtKsinNnEyXW+6x+gR+rG/Zy/dg3o1tBmJM
Bc7XTVwNhISvEsA1ZEhVzKud0KNZ46KioUFuATlgrxw7jM3mz56pZV5LM59ahXCr
9dbSAvrEEmgYrOHVhK7HzTeISnV7jvkJOpyKcqmz9vmXfNyOmuOeKIzFy5vfoDbq
n+L3l67Fnt+Eu796Hgt/QdtKuLVGu5YoGhTSDyjwgVnAEblTSvd8zQz6l27wV92+
J9N5p7IycSvgaXgS0hug5L8U3p0t64L5KaM4juW8msLPtjKDvcgPNBP6bvJEy/L1
MX/bzJmzTTvv0QuFmEoFYvNl7Vq/3mRPHgWO4xltN2/mC8ZQ1/t0kQrykCHXD1+N
oeQLPvqPRwqT69I4PEDc0plV39rMJwX3nJa7rgfSsMLpSsoGijdJ2Xm2enZ6xcSk
HjkmPPBE1rzMzQuS8NuCNc5YlfHb+mY7Uz3YraBR3DGkBVd9TkUAUL7Us37Gvj02
JtEqUBvyb6kWXdB+XJCBIpL1J5JiXRRd64f1oD2ucjiZUYzky4wZigw89t5v+EpU
IngkcsXAVPPxVAyQwk6ulpR9WW6urv41T+1hrzbujTO+1FBtPg87nVh0QPAJfCQi
eSSqRpfEuQH9p1uoGYNnLd1cNiLSP8lUUH+2dGdNYl+jRjw0v+uxtIZP864YqaeW
+bN1CJSE9Xqvzeq/z+H4//txfUMhUlDgjw8L53nEC+zVlrMGdSBTVmYo7EzyyhFC
IWMu/V1tJh3hN2Vb/C3YNIPnDo7xGyd4MwiJOfRJ3I3UaZnSo4bsrMocXUHUG83w
oOcyz5X/fC7owjqvpxLNVvag2RQXN9yXOSwTL/Pa95Vy4AlC8/X4d7Ti3L4GfxQQ
35Ou3ruLOj/tK/mvfeMoTbewgNGc73PunNuczmu7h/0btasxLpp8F+3iqf5owhfR
fqZDV4PpXeyl21VUjXCTre9eGx3jdjB17RA3qhyXB221Md6pCLAczPRivv68ZHfE
+ImrYvJBmu4sixOKPtAVx8ZOOIFv2DoNuUpiTrPBng9dsHdc6QD+9zPYYvmuMEub
ip8IJwjImgWKLILjSvH9DzkoEFpD9YxsIxeSyAW0W4vQHexbj2djSjIobEha/vk8
MRPB/k0Tf371VEXpRwjtJWzo4wfnJ//H/m0uZ7Q0tp5fpvHcXAxNr4JR8VCxL7Nu
EkheAnR0OziYhmP6l9WGcF2cq0Tzm9wNbrLdT1WpnhR36rzyYd6+pSuMRQBVOSL/
2XKBLUc6FEhmRv90tKAnPgK8Awv2s9WHgIOX83FYDB5/FpmThnIzZRnNLGkXXu/i
eyXO3J23F3wc9jJRRPWCYz2O/KdhBIRs5gPrA9yAZqfs5ywPQjuHpaBz+g9e4fXK
CiGUUOL9WleLSA37hBcWJ7B6E+Kd52oetKMcNXhS5m7Eil7TeKK5PDImHsXrQZVv
PUZ5LAfSMIPG3YBjfmJCvrsBq1f66WvaviRmhhERRg8H8p31sfHcgdLJB4C+QkWD
UU8vbEBlYvuWrCuhH4D+r8spKUnxNnDQQbYmTFpf/S9Z1T6g9XINTc/pBSRjIs21
KghDaX/6FNUgQlkc8ow2WCkaoxoerwDSA7y5EXn3AE3KsabU9/nJKUDpwoZ/0aCj
WTWUmtuXEInTO8wV26dt1A4q0Ml/DvyYVgj7uPp05XIiQivGnlO667Eyzcc8dKFs
wPLUzr7plyTHo+h+N136aJF3uSmi9MI4Re0a9AKC0vcSH8jLCXulR9lc8jRwMf2I
njk5IYHcKW2N4qmtzjCJacVtdfQrp1a5LQwmWtn6nku7IGdW2cHJ0VeFYp2+sCbw
B0PkA1k9/GMJzuAmwNjqLGUkGwsnZiKrz1xA+ztUtcKLWrKCXkFpa4BaKasF6QZy
Xveb7Ya0PS18SLJT2ir0hQLnA6PTPPabp79NRNT+QXBuvbWPpI8xE749jiL6SwrJ
KX+tHioXXLS9SLPiqQAJ3q0XhrmvKYRK0v/X2Sa0EweveNe4fnqrL9yFbuUyuGgp
I8cBL/YNRfyV6qRPg2tCsw==
`pragma protect end_protected
