// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
3H961NIMvuwvj/oZLnXS7LkRCJmhm4Bf+hPDHC711FHTUEvS0c0h4ycvS4W/pVMs
7/lQ7lZm5lUUc79kdHbyENhRbG091k7hiAsERpNIkfyUrn2D5PCscnf5CmYEDisv
0jaRKEA5oA5g7S1I8GqstrpuzFNcVbNgzNTQXHXLEEc=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 4480 )
`pragma protect data_block
1BWrrT51VdfMZ9bWSGRnNI0hh8hIOwhrK99Krjup8Co5KCQsL+QW2P4rZBlP6Hyw
1ZXZLwkdKKxb6xTk9rKYAsV2FdSPMWy34KCdiIiA/lJHyRnZFvYN8Yr+qYLKJQIi
/+TYsnOz9ATSHJrPsryTUE1f3om407aie10bAD74ZcPswEu+iVXL1W/tsxfXqT0z
XdEjSrF4HwEt7jKz8/iBl23h27K2tVoo62493v4/rjvYjo5mV4K8Lv0LhszE+4GC
m5MxoIXpNxjZF4F1HXdzIKlt5bgP5Z7GBxi20avFIznas39RtOkwlv7ZQUWHVksY
PuBeNE4+KKC+ufr3VC6AGBUDBtE/oz97OKD6vJh1LANBYlGKveuFuVrarpop5kg/
v/lZrOZ2nmwq7R3H+MUta9vdTQkn31+fHTlCo8y8AIdNyuUTPSBEj1rbMHheMrgb
b4D27JVv7KVWd0G62gfqdRFIYSoJxhMyuX5ECYPetBR6s2yIZWm2/z4vqTafvREe
8tUSYwUdA85HGvYgcODNSACJ65xCKDL1IsA+XYCsr32g+UOAghfHKnToSjvPTFg0
JsROz6tt0lfqr8MQeYj3E3+6N99sU32KwWoqMtFmtAbqSRLBrmoidQGCtozG1z3H
AQ/+ghoSOXedo3h32Au4ZzUVbncTBFyYilfGV/TTNtMNyuzCwOqHC1y0BVnkC6tA
RZwSJGToMN2nGD5mbOQBrBFZC1xnvVxeB7w9Me99QY1mSGXXK8x+AGN5gbqpnMY/
yX3nTbXCex3LptxBMawhd3JtaTj5tZkDgYRqeC+/4FVihSzFpUay4+uyBeLe5CNF
+iZc9//7x0gODKjJ4dBEdSUW4G6cXVHjXSLFrcNknzAV2ZWSo59LWqfY96sNP03w
qoWl1jFu6V46CKjDFHFZjgqOwh3DTIjiYz1GW7opj1Bcx4YT73KBt09v3WR3NYxY
3CKnWZo9YHl19tBkshR41fEjZCDsSrsZ09yAz+swuTo/CAy/Xr80u4VJlZbT3bul
mOL1YAIRPbDRJ7sxvOxm4bPz5DdGAsJNS81vLTRJJmpRA21qW3iia/Bqao9HyAc5
f7iJVaxBi49VweY+ESZxMOfJKcQPRfThForLmhXPG1NxMo2HrPp4HDKKd8NFmwbq
UFRXHmkd9JEln8Vb05KwX2H+9D6DGJ8cLb5jLP0QrwwQlWdVQVsToeAyZRxDpyMl
p8qEbZTuDgV0IcO3tSDSyyNhC4ypvS1jzMTpTZAHTz4Kg9euKKpzaQeqAwbaLUNd
dpGP7ljpHLVuGrBzfQrkIFsnS/HIAw+89A2FoMpEYXRvrMjDzQShEbpPWrR3ktuA
4peGiudeNYAjnib14s8IE6if93h/qfdhKKUEoYjDPAcuIG+NUpNPvuJSICAlbepR
GMjJ0zsyJ1ETpjvnNn/gJn0H/hBRxLj0suVqkedUX22Wyg22vAyoMrMna/Gi3INS
iIQBes5FbX30mS9J1qaMwGpLkuBeROnUdzzpKAn7IRv1An1PGrn2KJv1Q+NhhtXk
8RHZ49+c8N8jx/ftIjsXAv/Z1mNOKmEomWx4Rwkgq5dWlDJOhSr1pFPSBt0pAscH
O/amZd1p28ka+7EeyeIr0//p/8HBSzTv17AMA8GL7lMc7nXOx1RGZNFU366dNzDM
nm5kOJtlX+3xeMS/RPVTlzXrSqv2DbmtOXZ9lkO+oMd05jP5TcjM350vTfcPLCt0
Z/98uVyezKcuh2tRTaCExSHfi9Xrrh6Z4nz6n1kzjwPzPn4nnLll9XEei0tfquU7
XpkNHPX1qHTEtfV5S/Xe+nlAWBxS9SlKDxLJT2Vn41RXPDQAXWJy+zMG3TtHH52n
N0pbKpRn8q/36jt6YRoS1KqS16vmWgfSuzYQtcetSc7PIYKWwR+3TEIW9BUVODWD
tpphQbAEnEbyG2hwoWq10nTl0OwXtPEfCws38akdUGvmv8HN8KIraFLGlPFeMdgu
j83dl+XnLrfKvijeguMBDaZ8VtRADHb+l9j5z000fDn1daCHx31zzN4zCx4F/ViB
o5xqeyEUzfcl27dit3jI5LzdPVuflCXNvJq41cNhCQw+JHQO1J5BoCyp2+38D0de
FdR1Ov3BGbv8AkWFc/tgVY0i4l7N95/1dxC2EGcN/EOpOM0t5gxW74r/SrgV006L
NYTftzDa6yf3NeI7F/CLAHH0P1P4uAr9P4ycAuk+4nZf3a0rprwithKSvlW8Jr9L
hr0/v3OnGCCeVGzB84bC77OKz3MpxTQaThcr1GQdKOsPHv4NUIlceFQHCfKBketL
DjixAUsojVRTrZNxhE8cVpmxB4KnJRmi81NR9DhQGnZNM0PC8AJ8AMegTwe/1ZTo
W5UAUwlltHSOIwqNk59NmxiiDuuGZNIqdF5fZAyseFFDaVfV6hQM4aZZK+STcKpZ
7I25e4azwDRO/m4ZaKi+4vpOIpJoV3EzGxb2W4FCZ4qbwLW4bpqOKycAiPG4CKCj
TiS9KytOQibbRc1/Ma+ZRak/9oHaQrgwkN+d30f8I8IbvvfuEey8qJ4uWtJu1ZFD
0/l18IWIKvEmNh5oC+RblYT51hk9ftQLns79RltX8Htm9g6FLmIZtzdExr6Xfi+2
kFa+nhk7nw4W3Ml4rgFMNxnmxuxyr/X8xPPvxLL4Lm8PbGwujmuUr8/t3zm9prCy
W/K2op84A14/vM5VzjD5+Boi+6fzPrCfnqBtAbUt1+SHzSvIlHXFJm14YvWwjVJL
j4zU1TfdVsSMH+W5lypzGtZdmD7umYxLSKIX7icnSBj9uy0VIvP2cEAojUZ703DR
hFO736cf5B25aQvPTlABggM6BrOXZ63pg5afHvo5PScz3IqG+yD2voTkcZkZoY74
HwfXivlC7ameXAxcnD88XrINx1LAWEzKCbIy+O0pshFRLhQ4DcYKXc9Q4RhXoQE3
b3fRmoVd1Dr/Gm77RuF1IXSRDjjJDAfwF4dabg+0fFSD4OF5Iivl62cp5vtAfoCC
mA09LIJgEQ6+plW4bGF5wxfhrRvoizpB6YVGtASS0grLCgSZFpG2uDr/dVZtlFSh
A9P/rvZQ8y2lP04CrqRPu02iNdzTC50HBdYqE047QpywLDapfBvbnpWXaNHSiGC3
lU1uyx/g+JkmEqEqc5WShYpOPS9hZUC4EDCJ8ofs7bA83jLqURbNh1sTpTJFIRCU
D52lCFBtaW/EFQXNazyug7P62mK7H6P3Np7D+NmSrj21WtoQpZBybaTfg9y3eRU4
x7/SWJMsNtaVMPJM6mQBoOFJzLAgaSAb3+j1Ez58YPhy/QAQImZ9g6YogDsXXf8O
X+xI4PNwo3sJVuHbhuSiNGxa9Exq0j/U6DSz01N6A08UDcPvRn532lM/paAz7xAJ
rC2NT3ylWE3YI0ghv+CRoTUzh7nAFvBo3IggegZNYcaiy4FeS+R3UFQ/YDWoM/rm
OVYuh0rCGGNEH85m2AdDr/otiH21XsRS1HNkjM19+TGffN9Jhhk+m6PNzTh5UYXq
0VYHPtqOXwymLaFafwxnxNtJ00dQiJdaRpEDnc5dbJSteR6yQO+LLXoX5Z+XNfcJ
sM6/B2pEo6EdEM5sZddk4d8/S1OnpozWUc4e9gReB426R28HA1SrDHw4XKhDI7oc
+LveFwJ7gxv0K571ia3KOIp6aPvataLkU5s9OZcKQL3INap3q31TzXOyg5duV48D
R6qYZsbCHLJqs9SvstOTx2diweej2bHJCLEvKnIwPnnSl8WSeEFs64/0VYG7lEHz
8bz/PHotY5zxWuLelZbc3MAk1CyCjo6yHKLWUpGzfIevEJLpqlj/DGfhyixMB7jl
TYeDJ928HfqUbqLYvzdw9zsZ8sAHK5nnYSBf6ApfGlwe1hj4cxkQ6L/Xs5Y8irf8
paQfTomTEaSaVdwH1qt6D6DJHOvWRJISyeKd6rPm3ZX55vxuabWYyDHHL8bvsxfo
JXsQ8CDtTGslrkL+DG6tDDECkRNDQa1RySBaakG0gTjbEb2sye4S5ewHOXlFLNB5
E+0TQZb0tU/awV7q0/JvPPowhmctWPf2QcSG3FsoLcggoNcy5y3URygoq0439t0K
CQEEiVtY77CizJIqNJ5qTAlqmxRqd53kzkmovPuuBV0P/QRE12S3AJc6qbAoXjWJ
OeIF9oE0G7MyhtiF2zKoOmoyBOPRvT7gapAWU7Cs7AGBF1C6z+Repn3Ilg0Vph2o
uqwVa2jw7F9ZBcXm3RPh4E1IhMR9wcEaB+4cN8NTuNP13GMuxqi9UvPSuF0tPz4g
RtnaQTlrQZjA3+DO6zZxacnEn8/ij5pSu2bUF/kV5M46YNpqFQrICldWNGWeYaio
22ykKShJ1xLrCpvqJEFrjlcovE08aRF4plGLFr5WqxuHDBOfRDkq1/1SzGz6C5Tr
FNhWeThFrc6A7dE1zCp4Tr8POckUiYsDa2Yvd36Hwzqxx8jpTDBR4WjMHQgSAUIp
gkpDulGpVmhoST0ZchyEVr0a7EggltnI9udk+zi6NDCRQmRn4TCaKlW0xdiljiaA
7LCIoralYyxAiH0GqVr0TmxTd8Loo55jtq2ZdgPIi4bi69j6WQeQSSc3nw5zwskc
U0brR7P5HHqCz1t2+kWuvIkhLs4PGDX9qQOrn4+T+6L9av30TRkupCQsOFA2rFBn
S1EiLwUhYBFNEZ0U8ZEs9aQbepfJEnJDOGoaegtSFuZFxj3uNcj2+NCmlgnLEsSi
VBtcl2YCIg+Pdi/Cn6FvvIhh9Zn6VRvvlct1xXsqZpEbVXBEHeFBl60Xq/dueofZ
Ry1tl02l/SSZ9161Zg1/kOyVcFO8CY8JaMVWre7Quj+bOpj3g47JBvw6K/wj92Z7
paC1LJwMdT4LuHWW1MgSW79dl9z+GT2Vcioxc0Vu1Lx2P292YS2I6QsTPEF/Xz97
GdNF2bmFaXtFKoM2rgGlsN54+kz911bcG/l78vs3R2pRPTWiB6zWI/CT+TcSF9H2
LTDmr/g3CDm8zyKMK6esP57ZIV3v3LOXbmLoVfJptbXsLvTXrywLj8h/uMWsC/dh
ywr9KmyBixBtfrCoUjM23pC3G2PC9QUS0+zaqOiQJLPHsqoh4oPvI6zEza1lsAgS
ADJNFxVLA1PFc+AsjlvTe4YS+G5UFs7URPXiSsOMUlHB57qxhBifb97CWQAVPYLa
VyCMoa0SYr4sEV9Qj5U/+WGj5lG9oS03LqauZcK2IQWDFgArUYy6SaJ1idY/U9lg
BpNJsnPCwNxAiX7yUMJzjpIzCdghM1w1A6SrIIFPmkESv6QXFkL+l4Q2wHLolvYI
JkT87wanBp4x9C6/YPsEFBAZ1SjYqEZKzykw1MCPflPY/9e7eyeSQzCPdiUcx4Zs
lbdd1N9JWwUL+6K98XTV5HX4zVjMsE1b5zDrT4vohSFIhGDMDbXq6bzl6v5M0og4
MJGoc4GxdCjfQdBb/rC7vkm1VhaGKqw+SHmmJ9Pr/+BALL9jmvcMlnpGW417Su2x
4K5esD7t/u1nS2HEoTTiAy5dYVF+gPLntWSdbaH44XDxxdDHhLTXIFw1bmgxhPSc
GfAEW7Bg50jKbd6jT7xJFOgZsTO49KTVc+uu9zvX3VZbkiQeCPmlru1vn6lCW5aH
TaxIBCp20+tWdyVlQ7vrhPZFju/Za6OKx+gisi6mh6QANhc+vnCCrRN6ngTXLSB1
8mqnzeHyYWJzWlyWCGPaAh7DFCQqXOT6HwlZTB3ITmKPZhBn/U7NGfGnHRcyj3Uj
vM8f9T43YVZNAOUhpYqINlpyezo8R6yfGIYTDeE3XWOywmSKuAuIvC+jEtdD8Un/
GoeSammTO9s3xdiEzHUi0Lo23651bq1XOw8idCQbhng4r6R7E660zWSc/u24lYbS
co6Wobg+WrqzG1HjwjUp/R8umSFG8stYQom+S0gR+lfYnkZPHB4u5KxwCWEE0fdg
5FVuSkg1ax1xoZ104q6wPQ==

`pragma protect end_protected
