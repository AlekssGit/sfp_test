// pcie.v

// Generated using ACDS version 21.4 67

`timescale 1 ps / 1 ps
module pcie (
		output wire         coreclkout_hip,           //    coreclkout_hip.clk
		input  wire         refclk,                   //            refclk.clk
		input  wire         npor,                     //              npor.npor
		input  wire         pin_perst,                //                  .pin_perst
		output wire         app_nreset_status,        // app_nreset_status.reset_n
		input  wire [31:0]  test_in,                  //          hip_ctrl.test_in
		input  wire         simu_mode_pipe,           //                  .simu_mode_pipe
		input  wire         sim_pipe_pclk_in,         //          hip_pipe.sim_pipe_pclk_in
		output wire [1:0]   sim_pipe_rate,            //                  .sim_pipe_rate
		output wire [4:0]   sim_ltssmstate,           //                  .sim_ltssmstate
		output wire [2:0]   eidleinfersel0,           //                  .eidleinfersel0
		output wire [2:0]   eidleinfersel1,           //                  .eidleinfersel1
		output wire [2:0]   eidleinfersel2,           //                  .eidleinfersel2
		output wire [2:0]   eidleinfersel3,           //                  .eidleinfersel3
		output wire [1:0]   powerdown0,               //                  .powerdown0
		output wire [1:0]   powerdown1,               //                  .powerdown1
		output wire [1:0]   powerdown2,               //                  .powerdown2
		output wire [1:0]   powerdown3,               //                  .powerdown3
		output wire         rxpolarity0,              //                  .rxpolarity0
		output wire         rxpolarity1,              //                  .rxpolarity1
		output wire         rxpolarity2,              //                  .rxpolarity2
		output wire         rxpolarity3,              //                  .rxpolarity3
		output wire         txcompl0,                 //                  .txcompl0
		output wire         txcompl1,                 //                  .txcompl1
		output wire         txcompl2,                 //                  .txcompl2
		output wire         txcompl3,                 //                  .txcompl3
		output wire [31:0]  txdata0,                  //                  .txdata0
		output wire [31:0]  txdata1,                  //                  .txdata1
		output wire [31:0]  txdata2,                  //                  .txdata2
		output wire [31:0]  txdata3,                  //                  .txdata3
		output wire [3:0]   txdatak0,                 //                  .txdatak0
		output wire [3:0]   txdatak1,                 //                  .txdatak1
		output wire [3:0]   txdatak2,                 //                  .txdatak2
		output wire [3:0]   txdatak3,                 //                  .txdatak3
		output wire         txdetectrx0,              //                  .txdetectrx0
		output wire         txdetectrx1,              //                  .txdetectrx1
		output wire         txdetectrx2,              //                  .txdetectrx2
		output wire         txdetectrx3,              //                  .txdetectrx3
		output wire         txelecidle0,              //                  .txelecidle0
		output wire         txelecidle1,              //                  .txelecidle1
		output wire         txelecidle2,              //                  .txelecidle2
		output wire         txelecidle3,              //                  .txelecidle3
		output wire         txdeemph0,                //                  .txdeemph0
		output wire         txdeemph1,                //                  .txdeemph1
		output wire         txdeemph2,                //                  .txdeemph2
		output wire         txdeemph3,                //                  .txdeemph3
		output wire [2:0]   txmargin0,                //                  .txmargin0
		output wire [2:0]   txmargin1,                //                  .txmargin1
		output wire [2:0]   txmargin2,                //                  .txmargin2
		output wire [2:0]   txmargin3,                //                  .txmargin3
		output wire         txswing0,                 //                  .txswing0
		output wire         txswing1,                 //                  .txswing1
		output wire         txswing2,                 //                  .txswing2
		output wire         txswing3,                 //                  .txswing3
		input  wire         phystatus0,               //                  .phystatus0
		input  wire         phystatus1,               //                  .phystatus1
		input  wire         phystatus2,               //                  .phystatus2
		input  wire         phystatus3,               //                  .phystatus3
		input  wire [31:0]  rxdata0,                  //                  .rxdata0
		input  wire [31:0]  rxdata1,                  //                  .rxdata1
		input  wire [31:0]  rxdata2,                  //                  .rxdata2
		input  wire [31:0]  rxdata3,                  //                  .rxdata3
		input  wire [3:0]   rxdatak0,                 //                  .rxdatak0
		input  wire [3:0]   rxdatak1,                 //                  .rxdatak1
		input  wire [3:0]   rxdatak2,                 //                  .rxdatak2
		input  wire [3:0]   rxdatak3,                 //                  .rxdatak3
		input  wire         rxelecidle0,              //                  .rxelecidle0
		input  wire         rxelecidle1,              //                  .rxelecidle1
		input  wire         rxelecidle2,              //                  .rxelecidle2
		input  wire         rxelecidle3,              //                  .rxelecidle3
		input  wire [2:0]   rxstatus0,                //                  .rxstatus0
		input  wire [2:0]   rxstatus1,                //                  .rxstatus1
		input  wire [2:0]   rxstatus2,                //                  .rxstatus2
		input  wire [2:0]   rxstatus3,                //                  .rxstatus3
		input  wire         rxvalid0,                 //                  .rxvalid0
		input  wire         rxvalid1,                 //                  .rxvalid1
		input  wire         rxvalid2,                 //                  .rxvalid2
		input  wire         rxvalid3,                 //                  .rxvalid3
		input  wire         rxdataskip0,              //                  .rxdataskip0
		input  wire         rxdataskip1,              //                  .rxdataskip1
		input  wire         rxdataskip2,              //                  .rxdataskip2
		input  wire         rxdataskip3,              //                  .rxdataskip3
		input  wire         rxblkst0,                 //                  .rxblkst0
		input  wire         rxblkst1,                 //                  .rxblkst1
		input  wire         rxblkst2,                 //                  .rxblkst2
		input  wire         rxblkst3,                 //                  .rxblkst3
		input  wire [1:0]   rxsynchd0,                //                  .rxsynchd0
		input  wire [1:0]   rxsynchd1,                //                  .rxsynchd1
		input  wire [1:0]   rxsynchd2,                //                  .rxsynchd2
		input  wire [1:0]   rxsynchd3,                //                  .rxsynchd3
		output wire [17:0]  currentcoeff0,            //                  .currentcoeff0
		output wire [17:0]  currentcoeff1,            //                  .currentcoeff1
		output wire [17:0]  currentcoeff2,            //                  .currentcoeff2
		output wire [17:0]  currentcoeff3,            //                  .currentcoeff3
		output wire [2:0]   currentrxpreset0,         //                  .currentrxpreset0
		output wire [2:0]   currentrxpreset1,         //                  .currentrxpreset1
		output wire [2:0]   currentrxpreset2,         //                  .currentrxpreset2
		output wire [2:0]   currentrxpreset3,         //                  .currentrxpreset3
		output wire [1:0]   txsynchd0,                //                  .txsynchd0
		output wire [1:0]   txsynchd1,                //                  .txsynchd1
		output wire [1:0]   txsynchd2,                //                  .txsynchd2
		output wire [1:0]   txsynchd3,                //                  .txsynchd3
		output wire         txblkst0,                 //                  .txblkst0
		output wire         txblkst1,                 //                  .txblkst1
		output wire         txblkst2,                 //                  .txblkst2
		output wire         txblkst3,                 //                  .txblkst3
		output wire         txdataskip0,              //                  .txdataskip0
		output wire         txdataskip1,              //                  .txdataskip1
		output wire         txdataskip2,              //                  .txdataskip2
		output wire         txdataskip3,              //                  .txdataskip3
		output wire [1:0]   rate0,                    //                  .rate0
		output wire [1:0]   rate1,                    //                  .rate1
		output wire [1:0]   rate2,                    //                  .rate2
		output wire [1:0]   rate3,                    //                  .rate3
		input  wire         rx_in0,                   //        hip_serial.rx_in0
		input  wire         rx_in1,                   //                  .rx_in1
		input  wire         rx_in2,                   //                  .rx_in2
		input  wire         rx_in3,                   //                  .rx_in3
		output wire         tx_out0,                  //                  .tx_out0
		output wire         tx_out1,                  //                  .tx_out1
		output wire         tx_out2,                  //                  .tx_out2
		output wire         tx_out3,                  //                  .tx_out3
		output wire [81:0]  msi_intfc_o,              //         msi_intfc.msi_intfc
		output wire [15:0]  msi_control_o,            //       msi_control.msi_control
		output wire [15:0]  msix_intfc_o,             //        msix_intfc.msix_intfc
		input  wire         intx_req_i,               //        intx_intfc.intx_req
		output wire         intx_ack_o,               //                  .intx_ack
		input  wire [63:0]  txs_address_i,            //               txs.address
		input  wire         txs_chipselect_i,         //                  .chipselect
		input  wire [15:0]  txs_byteenable_i,         //                  .byteenable
		output wire [127:0] txs_readdata_o,           //                  .readdata
		input  wire [127:0] txs_writedata_i,          //                  .writedata
		input  wire         txs_read_i,               //                  .read
		input  wire         txs_write_i,              //                  .write
		input  wire [5:0]   txs_burstcount_i,         //                  .burstcount
		output wire         txs_readdatavalid_o,      //                  .readdatavalid
		output wire         txs_waitrequest_o,        //                  .waitrequest
		input  wire         cra_chipselect_i,         //               cra.chipselect
		input  wire [13:0]  cra_address_i,            //                  .address
		input  wire [3:0]   cra_byteenable_i,         //                  .byteenable
		input  wire         cra_read_i,               //                  .read
		output wire [31:0]  cra_readdata_o,           //                  .readdata
		input  wire         cra_write_i,              //                  .write
		input  wire [31:0]  cra_writedata_i,          //                  .writedata
		output wire         cra_waitrequest_o,        //                  .waitrequest
		output wire         cra_irq_o,                //           cra_irq.irq
		output wire [63:0]  rxm_bar0_address_o,       //          rxm_bar0.address
		output wire [15:0]  rxm_bar0_byteenable_o,    //                  .byteenable
		input  wire [127:0] rxm_bar0_readdata_i,      //                  .readdata
		output wire [127:0] rxm_bar0_writedata_o,     //                  .writedata
		output wire         rxm_bar0_read_o,          //                  .read
		output wire         rxm_bar0_write_o,         //                  .write
		output wire [5:0]   rxm_bar0_burstcount_o,    //                  .burstcount
		input  wire         rxm_bar0_readdatavalid_i, //                  .readdatavalid
		input  wire         rxm_bar0_waitrequest_i,   //                  .waitrequest
		output wire [63:0]  rxm_bar2_address_o,       //          rxm_bar2.address
		output wire [15:0]  rxm_bar2_byteenable_o,    //                  .byteenable
		input  wire [127:0] rxm_bar2_readdata_i,      //                  .readdata
		output wire [127:0] rxm_bar2_writedata_o,     //                  .writedata
		output wire         rxm_bar2_read_o,          //                  .read
		output wire         rxm_bar2_write_o,         //                  .write
		output wire [5:0]   rxm_bar2_burstcount_o,    //                  .burstcount
		input  wire         rxm_bar2_readdatavalid_i, //                  .readdatavalid
		input  wire         rxm_bar2_waitrequest_i,   //                  .waitrequest
		input  wire [15:0]  rxm_irq_i                 //           rxm_irq.irq
	);

	pcie_altera_pcie_a10_hip_2011_ub5pqua #(
		.force_tag_checking_on_hwtcl                          (0),
		.bar0_address_width_mux_hwtcl                         (16),
		.bar1_address_width_mux_hwtcl                         (0),
		.bar2_address_width_mux_hwtcl                         (30),
		.bar3_address_width_mux_hwtcl                         (0),
		.bar4_address_width_mux_hwtcl                         (0),
		.bar5_address_width_mux_hwtcl                         (0),
		.data_width_integer_hwtcl                             (128),
		.data_width_integer_rxm_txs_hwtcl                     (128),
		.data_width_integer_txs_hwtcl                         (128),
		.data_byte_width_integer_hwtcl                        (16),
		.reconfig_address_width_integer_hwtcl                 (12),
		.burst_count_integer_hwtcl                            (6),
		.empty_integer_hwtcl                                  (1),
		.include_dma_hwtcl                                    (0),
		.txs_addr_width_integer_hwtcl                         (64),
		.interface_type_integer_hwtcl                         (1),
		.dma_width_hwtcl                                      (128),
		.dma_be_width_hwtcl                                   (16),
		.dma_brst_cnt_w_hwtcl                                 (6),
		.avmm_addr_width_hwtcl                                (64),
		.cb_pcie_mode_hwtcl                                   (0),
		.cb_pcie_rx_lite_hwtcl                                (0),
		.cg_impl_cra_av_slave_port_hwtcl                      (1),
		.cg_enable_advanced_interrupt_hwtcl                   (1),
		.cg_enable_a2p_interrupt_hwtcl                        (1),
		.internal_controller_hwtcl                            (1),
		.enable_rxm_burst_hwtcl                               (0),
		.extended_tag_support_hwtcl                           (0),
		.cg_a2p_addr_map_num_entries_hwtcl                    (2),
		.cg_a2p_addr_map_pass_thru_bits_hwtcl                 (12),
		.lane_rate_hwtcl                                      ("Gen2 (5.0 Gbps)"),
		.enable_avst_reset_hwtcl                              (1),
		.multiple_packets_per_cycle_hwtcl                     (0),
		.use_tx_cons_cred_sel_hwtcl                           (0),
		.cseb_autonomous_hwtcl                                (0),
		.speed_change_hwtcl                                   (0),
		.hip_reconfig_hwtcl                                   (0),
		.xcvr_reconfig_hwtcl                                  (0),
		.export_phy_input_to_top_level_hwtcl                  (0),
		.adme_enable_hwtcl                                    (0),
		.enable_devkit_conduit_hwtcl                          (0),
		.enable_skp_det                                       (0),
		.DEBUG_WIDTH                                          (16),
		.enable_g3_bypass_equlz_rp_sim_hwtcl                  (0),
		.expansion_base_address_register_hwtcl                (0),
		.pf0_vf_device_id_hwtcl                               (0),
		.pf0_subclass_code_hwtcl                              (0),
		.pf0_pci_prog_intfc_byte_hwtcl                        (0),
		.enable_completion_timeout_disable_hwtcl              (1),
		.slot_clock_cfg_hwtcl                                 (1),
		.msix_table_offset_hwtcl                              (0),
		.msix_pba_offset_hwtcl                                (0),
		.reserved_debug_hwtcl                                 (0),
		.include_sriov_hwtcl                                  (0),
		.app_msi_req_fn_hwtcl                                 (8),
		.cfg_num_vf_width_hwtcl                               (8),
		.flr_completed_vf_width_hwtcl                         (4),
		.sriov2_en                                            (1),
		.enable_custom_features_hwtcl                         (0),
		.pf0_extra_bar_present_hwtcl                          (0),
		.pf0_extra_bar_size_hwtcl                             (12),
		.devhide_support_hwtcl                                (0),
		.device_embedded_ep_support_hwtcl                     (0),
		.total_pf_count_hwtcl                                 (1),
		.pf0_vf_count_hwtcl                                   (0),
		.pf1_vf_count_hwtcl                                   (0),
		.pf2_vf_count_hwtcl                                   (0),
		.pf3_vf_count_hwtcl                                   (0),
		.total_vf_count_hwtcl                                 (4),
		.total_pf_count_width_hwtcl                           (1),
		.total_vf_count_width_hwtcl                           (1),
		.system_page_sizes_supported_hwtcl                    (1363),
		.sr_iov_support_hwtcl                                 (0),
		.enable_alternate_link_list_hwtcl                     (0),
		.ari_support_hwtcl                                    (0),
		.flr_capability_hwtcl                                 (0),
		.pf0_virtio_capability_present_hwtcl                  (0),
		.pf0_virtio_device_specific_cap_present_hwtcl         (0),
		.pf0_virtio_cmn_config_bar_indicator_hwtcl            (0),
		.pf0_virtio_cmn_config_bar_offset_hwtcl               (0),
		.pf0_virtio_cmn_config_structure_length_hwtcl         (0),
		.pf0_virtio_notification_bar_indicator_hwtcl          (0),
		.pf0_virtio_notification_bar_offset_hwtcl             (0),
		.pf0_virtio_notification_structure_length_hwtcl       (0),
		.pf0_virtio_notify_off_multiplier_hwtcl               (0),
		.pf0_virtio_isrstatus_bar_indicator_hwtcl             (0),
		.pf0_virtio_isrstatus_bar_offset_hwtcl                (0),
		.pf0_virtio_isrstatus_structure_length_hwtcl          (0),
		.pf0_virtio_devspecific_bar_indicator_hwtcl           (0),
		.pf0_virtio_devspecific_bar_offset_hwtcl              (0),
		.pf0_virtio_devspecific_structure_length_hwtcl        (0),
		.pf0_virtio_pciconfig_access_bar_indicator_hwtcl      (0),
		.pf0_virtio_pciconfig_access_bar_offset_hwtcl         (0),
		.pf0_virtio_pciconfig_access_structure_length_hwtcl   (0),
		.pf1_virtio_capability_present_hwtcl                  (0),
		.pf1_virtio_device_specific_cap_present_hwtcl         (0),
		.pf1_virtio_cmn_config_bar_indicator_hwtcl            (0),
		.pf1_virtio_cmn_config_bar_offset_hwtcl               (0),
		.pf1_virtio_cmn_config_structure_length_hwtcl         (0),
		.pf1_virtio_notification_bar_indicator_hwtcl          (0),
		.pf1_virtio_notification_bar_offset_hwtcl             (0),
		.pf1_virtio_notification_structure_length_hwtcl       (0),
		.pf1_virtio_notify_off_multiplier_hwtcl               (0),
		.pf1_virtio_isrstatus_bar_indicator_hwtcl             (0),
		.pf1_virtio_isrstatus_bar_offset_hwtcl                (0),
		.pf1_virtio_isrstatus_structure_length_hwtcl          (0),
		.pf1_virtio_devspecific_bar_indicator_hwtcl           (0),
		.pf1_virtio_devspecific_bar_offset_hwtcl              (0),
		.pf1_virtio_devspecific_structure_length_hwtcl        (0),
		.pf1_virtio_pciconfig_access_bar_indicator_hwtcl      (0),
		.pf1_virtio_pciconfig_access_bar_offset_hwtcl         (0),
		.pf1_virtio_pciconfig_access_structure_length_hwtcl   (0),
		.pf2_virtio_capability_present_hwtcl                  (0),
		.pf2_virtio_device_specific_cap_present_hwtcl         (0),
		.pf2_virtio_cmn_config_bar_indicator_hwtcl            (0),
		.pf2_virtio_cmn_config_bar_offset_hwtcl               (0),
		.pf2_virtio_cmn_config_structure_length_hwtcl         (0),
		.pf2_virtio_notification_bar_indicator_hwtcl          (0),
		.pf2_virtio_notification_bar_offset_hwtcl             (0),
		.pf2_virtio_notification_structure_length_hwtcl       (0),
		.pf2_virtio_notify_off_multiplier_hwtcl               (0),
		.pf2_virtio_isrstatus_bar_indicator_hwtcl             (0),
		.pf2_virtio_isrstatus_bar_offset_hwtcl                (0),
		.pf2_virtio_isrstatus_structure_length_hwtcl          (0),
		.pf2_virtio_devspecific_bar_indicator_hwtcl           (0),
		.pf2_virtio_devspecific_bar_offset_hwtcl              (0),
		.pf2_virtio_devspecific_structure_length_hwtcl        (0),
		.pf2_virtio_pciconfig_access_bar_indicator_hwtcl      (0),
		.pf2_virtio_pciconfig_access_bar_offset_hwtcl         (0),
		.pf2_virtio_pciconfig_access_structure_length_hwtcl   (0),
		.pf3_virtio_capability_present_hwtcl                  (0),
		.pf3_virtio_device_specific_cap_present_hwtcl         (0),
		.pf3_virtio_cmn_config_bar_indicator_hwtcl            (0),
		.pf3_virtio_cmn_config_bar_offset_hwtcl               (0),
		.pf3_virtio_cmn_config_structure_length_hwtcl         (0),
		.pf3_virtio_notification_bar_indicator_hwtcl          (0),
		.pf3_virtio_notification_bar_offset_hwtcl             (0),
		.pf3_virtio_notification_structure_length_hwtcl       (0),
		.pf3_virtio_notify_off_multiplier_hwtcl               (0),
		.pf3_virtio_isrstatus_bar_indicator_hwtcl             (0),
		.pf3_virtio_isrstatus_bar_offset_hwtcl                (0),
		.pf3_virtio_isrstatus_structure_length_hwtcl          (0),
		.pf3_virtio_devspecific_bar_indicator_hwtcl           (0),
		.pf3_virtio_devspecific_bar_offset_hwtcl              (0),
		.pf3_virtio_devspecific_structure_length_hwtcl        (0),
		.pf3_virtio_pciconfig_access_bar_indicator_hwtcl      (0),
		.pf3_virtio_pciconfig_access_bar_offset_hwtcl         (0),
		.pf3_virtio_pciconfig_access_structure_length_hwtcl   (0),
		.pf4_virtio_capability_present_hwtcl                  (0),
		.pf4_virtio_device_specific_cap_present_hwtcl         (0),
		.pf4_virtio_cmn_config_bar_indicator_hwtcl            (0),
		.pf4_virtio_cmn_config_bar_offset_hwtcl               (0),
		.pf4_virtio_cmn_config_structure_length_hwtcl         (0),
		.pf4_virtio_notification_bar_indicator_hwtcl          (0),
		.pf4_virtio_notification_bar_offset_hwtcl             (0),
		.pf4_virtio_notification_structure_length_hwtcl       (0),
		.pf4_virtio_notify_off_multiplier_hwtcl               (0),
		.pf4_virtio_isrstatus_bar_indicator_hwtcl             (0),
		.pf4_virtio_isrstatus_bar_offset_hwtcl                (0),
		.pf4_virtio_isrstatus_structure_length_hwtcl          (0),
		.pf4_virtio_devspecific_bar_indicator_hwtcl           (0),
		.pf4_virtio_devspecific_bar_offset_hwtcl              (0),
		.pf4_virtio_devspecific_structure_length_hwtcl        (0),
		.pf4_virtio_pciconfig_access_bar_indicator_hwtcl      (0),
		.pf4_virtio_pciconfig_access_bar_offset_hwtcl         (0),
		.pf4_virtio_pciconfig_access_structure_length_hwtcl   (0),
		.pf5_virtio_capability_present_hwtcl                  (0),
		.pf5_virtio_device_specific_cap_present_hwtcl         (0),
		.pf5_virtio_cmn_config_bar_indicator_hwtcl            (0),
		.pf5_virtio_cmn_config_bar_offset_hwtcl               (0),
		.pf5_virtio_cmn_config_structure_length_hwtcl         (0),
		.pf5_virtio_notification_bar_indicator_hwtcl          (0),
		.pf5_virtio_notification_bar_offset_hwtcl             (0),
		.pf5_virtio_notification_structure_length_hwtcl       (0),
		.pf5_virtio_notify_off_multiplier_hwtcl               (0),
		.pf5_virtio_isrstatus_bar_indicator_hwtcl             (0),
		.pf5_virtio_isrstatus_bar_offset_hwtcl                (0),
		.pf5_virtio_isrstatus_structure_length_hwtcl          (0),
		.pf5_virtio_devspecific_bar_indicator_hwtcl           (0),
		.pf5_virtio_devspecific_bar_offset_hwtcl              (0),
		.pf5_virtio_devspecific_structure_length_hwtcl        (0),
		.pf5_virtio_pciconfig_access_bar_indicator_hwtcl      (0),
		.pf5_virtio_pciconfig_access_bar_offset_hwtcl         (0),
		.pf5_virtio_pciconfig_access_structure_length_hwtcl   (0),
		.pf6_virtio_capability_present_hwtcl                  (0),
		.pf6_virtio_device_specific_cap_present_hwtcl         (0),
		.pf6_virtio_cmn_config_bar_indicator_hwtcl            (0),
		.pf6_virtio_cmn_config_bar_offset_hwtcl               (0),
		.pf6_virtio_cmn_config_structure_length_hwtcl         (0),
		.pf6_virtio_notification_bar_indicator_hwtcl          (0),
		.pf6_virtio_notification_bar_offset_hwtcl             (0),
		.pf6_virtio_notification_structure_length_hwtcl       (0),
		.pf6_virtio_notify_off_multiplier_hwtcl               (0),
		.pf6_virtio_isrstatus_bar_indicator_hwtcl             (0),
		.pf6_virtio_isrstatus_bar_offset_hwtcl                (0),
		.pf6_virtio_isrstatus_structure_length_hwtcl          (0),
		.pf6_virtio_devspecific_bar_indicator_hwtcl           (0),
		.pf6_virtio_devspecific_bar_offset_hwtcl              (0),
		.pf6_virtio_devspecific_structure_length_hwtcl        (0),
		.pf6_virtio_pciconfig_access_bar_indicator_hwtcl      (0),
		.pf6_virtio_pciconfig_access_bar_offset_hwtcl         (0),
		.pf6_virtio_pciconfig_access_structure_length_hwtcl   (0),
		.pf7_virtio_capability_present_hwtcl                  (0),
		.pf7_virtio_device_specific_cap_present_hwtcl         (0),
		.pf7_virtio_cmn_config_bar_indicator_hwtcl            (0),
		.pf7_virtio_cmn_config_bar_offset_hwtcl               (0),
		.pf7_virtio_cmn_config_structure_length_hwtcl         (0),
		.pf7_virtio_notification_bar_indicator_hwtcl          (0),
		.pf7_virtio_notification_bar_offset_hwtcl             (0),
		.pf7_virtio_notification_structure_length_hwtcl       (0),
		.pf7_virtio_notify_off_multiplier_hwtcl               (0),
		.pf7_virtio_isrstatus_bar_indicator_hwtcl             (0),
		.pf7_virtio_isrstatus_bar_offset_hwtcl                (0),
		.pf7_virtio_isrstatus_structure_length_hwtcl          (0),
		.pf7_virtio_devspecific_bar_indicator_hwtcl           (0),
		.pf7_virtio_devspecific_bar_offset_hwtcl              (0),
		.pf7_virtio_devspecific_structure_length_hwtcl        (0),
		.pf7_virtio_pciconfig_access_bar_indicator_hwtcl      (0),
		.pf7_virtio_pciconfig_access_bar_offset_hwtcl         (0),
		.pf7_virtio_pciconfig_access_structure_length_hwtcl   (0),
		.pf0vf_virtio_capability_present_hwtcl                (0),
		.pf0vf_virtio_device_specific_cap_present_hwtcl       (0),
		.pf0vf_virtio_cmn_config_bar_indicator_hwtcl          (0),
		.pf0vf_virtio_cmn_config_bar_offset_hwtcl             (0),
		.pf0vf_virtio_cmn_config_structure_length_hwtcl       (0),
		.pf0vf_virtio_notification_bar_indicator_hwtcl        (0),
		.pf0vf_virtio_notification_bar_offset_hwtcl           (0),
		.pf0vf_virtio_notification_structure_length_hwtcl     (0),
		.pf0vf_virtio_notify_off_multiplier_hwtcl             (0),
		.pf0vf_virtio_isrstatus_bar_indicator_hwtcl           (0),
		.pf0vf_virtio_isrstatus_bar_offset_hwtcl              (0),
		.pf0vf_virtio_isrstatus_structure_length_hwtcl        (0),
		.pf0vf_virtio_devspecific_bar_indicator_hwtcl         (0),
		.pf0vf_virtio_devspecific_bar_offset_hwtcl            (0),
		.pf0vf_virtio_devspecific_structure_length_hwtcl      (0),
		.pf0vf_virtio_pciconfig_access_bar_indicator_hwtcl    (0),
		.pf0vf_virtio_pciconfig_access_bar_offset_hwtcl       (0),
		.pf0vf_virtio_pciconfig_access_structure_length_hwtcl (0),
		.pf1vf_virtio_capability_present_hwtcl                (0),
		.pf1vf_virtio_device_specific_cap_present_hwtcl       (0),
		.pf1vf_virtio_cmn_config_bar_indicator_hwtcl          (0),
		.pf1vf_virtio_cmn_config_bar_offset_hwtcl             (0),
		.pf1vf_virtio_cmn_config_structure_length_hwtcl       (0),
		.pf1vf_virtio_notification_bar_indicator_hwtcl        (0),
		.pf1vf_virtio_notification_bar_offset_hwtcl           (0),
		.pf1vf_virtio_notification_structure_length_hwtcl     (0),
		.pf1vf_virtio_notify_off_multiplier_hwtcl             (0),
		.pf1vf_virtio_isrstatus_bar_indicator_hwtcl           (0),
		.pf1vf_virtio_isrstatus_bar_offset_hwtcl              (0),
		.pf1vf_virtio_isrstatus_structure_length_hwtcl        (0),
		.pf1vf_virtio_devspecific_bar_indicator_hwtcl         (0),
		.pf1vf_virtio_devspecific_bar_offset_hwtcl            (0),
		.pf1vf_virtio_devspecific_structure_length_hwtcl      (0),
		.pf1vf_virtio_pciconfig_access_bar_indicator_hwtcl    (0),
		.pf1vf_virtio_pciconfig_access_bar_offset_hwtcl       (0),
		.pf1vf_virtio_pciconfig_access_structure_length_hwtcl (0),
		.pf2vf_virtio_capability_present_hwtcl                (0),
		.pf2vf_virtio_device_specific_cap_present_hwtcl       (0),
		.pf2vf_virtio_cmn_config_bar_indicator_hwtcl          (0),
		.pf2vf_virtio_cmn_config_bar_offset_hwtcl             (0),
		.pf2vf_virtio_cmn_config_structure_length_hwtcl       (0),
		.pf2vf_virtio_notification_bar_indicator_hwtcl        (0),
		.pf2vf_virtio_notification_bar_offset_hwtcl           (0),
		.pf2vf_virtio_notification_structure_length_hwtcl     (0),
		.pf2vf_virtio_notify_off_multiplier_hwtcl             (0),
		.pf2vf_virtio_isrstatus_bar_indicator_hwtcl           (0),
		.pf2vf_virtio_isrstatus_bar_offset_hwtcl              (0),
		.pf2vf_virtio_isrstatus_structure_length_hwtcl        (0),
		.pf2vf_virtio_devspecific_bar_indicator_hwtcl         (0),
		.pf2vf_virtio_devspecific_bar_offset_hwtcl            (0),
		.pf2vf_virtio_devspecific_structure_length_hwtcl      (0),
		.pf2vf_virtio_pciconfig_access_bar_indicator_hwtcl    (0),
		.pf2vf_virtio_pciconfig_access_bar_offset_hwtcl       (0),
		.pf2vf_virtio_pciconfig_access_structure_length_hwtcl (0),
		.pf3vf_virtio_capability_present_hwtcl                (0),
		.pf3vf_virtio_device_specific_cap_present_hwtcl       (0),
		.pf3vf_virtio_cmn_config_bar_indicator_hwtcl          (0),
		.pf3vf_virtio_cmn_config_bar_offset_hwtcl             (0),
		.pf3vf_virtio_cmn_config_structure_length_hwtcl       (0),
		.pf3vf_virtio_notification_bar_indicator_hwtcl        (0),
		.pf3vf_virtio_notification_bar_offset_hwtcl           (0),
		.pf3vf_virtio_notification_structure_length_hwtcl     (0),
		.pf3vf_virtio_notify_off_multiplier_hwtcl             (0),
		.pf3vf_virtio_isrstatus_bar_indicator_hwtcl           (0),
		.pf3vf_virtio_isrstatus_bar_offset_hwtcl              (0),
		.pf3vf_virtio_isrstatus_structure_length_hwtcl        (0),
		.pf3vf_virtio_devspecific_bar_indicator_hwtcl         (0),
		.pf3vf_virtio_devspecific_bar_offset_hwtcl            (0),
		.pf3vf_virtio_devspecific_structure_length_hwtcl      (0),
		.pf3vf_virtio_pciconfig_access_bar_indicator_hwtcl    (0),
		.pf3vf_virtio_pciconfig_access_bar_offset_hwtcl       (0),
		.pf3vf_virtio_pciconfig_access_structure_length_hwtcl (0),
		.pf_tph_support_hwtcl                                 (0),
		.pf0_tph_int_mode_support_hwtcl                       (0),
		.pf0_tph_dev_specific_mode_support_hwtcl              (0),
		.pf0_tph_st_table_location_hwtcl                      (0),
		.pf0_tph_st_table_size_hwtcl                          (63),
		.pf1_tph_int_mode_support_hwtcl                       (0),
		.pf1_tph_dev_specific_mode_support_hwtcl              (0),
		.pf1_tph_st_table_location_hwtcl                      (0),
		.pf1_tph_st_table_size_hwtcl                          (63),
		.pf2_tph_int_mode_support_hwtcl                       (0),
		.pf2_tph_dev_specific_mode_support_hwtcl              (0),
		.pf2_tph_st_table_location_hwtcl                      (0),
		.pf2_tph_st_table_size_hwtcl                          (63),
		.pf3_tph_int_mode_support_hwtcl                       (0),
		.pf3_tph_dev_specific_mode_support_hwtcl              (0),
		.pf3_tph_st_table_location_hwtcl                      (0),
		.pf3_tph_st_table_size_hwtcl                          (63),
		.vf_tph_support_hwtcl                                 (0),
		.pf0_vf_tph_int_mode_support_hwtcl                    (0),
		.pf0_vf_tph_dev_specific_mode_support_hwtcl           (0),
		.pf0_vf_tph_st_table_location_hwtcl                   (0),
		.pf0_vf_tph_st_table_size_hwtcl                       (63),
		.pf1_vf_tph_int_mode_support_hwtcl                    (0),
		.pf1_vf_tph_dev_specific_mode_support_hwtcl           (0),
		.pf1_vf_tph_st_table_location_hwtcl                   (0),
		.pf1_vf_tph_st_table_size_hwtcl                       (63),
		.pf2_vf_tph_int_mode_support_hwtcl                    (0),
		.pf2_vf_tph_dev_specific_mode_support_hwtcl           (0),
		.pf2_vf_tph_st_table_location_hwtcl                   (0),
		.pf2_vf_tph_st_table_size_hwtcl                       (63),
		.pf3_vf_tph_int_mode_support_hwtcl                    (0),
		.pf3_vf_tph_dev_specific_mode_support_hwtcl           (0),
		.pf3_vf_tph_st_table_location_hwtcl                   (0),
		.pf3_vf_tph_st_table_size_hwtcl                       (63),
		.pf_ats_support_hwtcl                                 (0),
		.pf0_ats_invalidate_queue_depth_hwtcl                 (0),
		.pf1_ats_invalidate_queue_depth_hwtcl                 (0),
		.pf2_ats_invalidate_queue_depth_hwtcl                 (0),
		.pf3_ats_invalidate_queue_depth_hwtcl                 (0),
		.vf_ats_support_hwtcl                                 (0),
		.pf0_bar0_present_hwtcl                               (1),
		.pf0_bar1_present_hwtcl                               (0),
		.pf0_bar2_present_hwtcl                               (0),
		.pf0_bar3_present_hwtcl                               (0),
		.pf0_bar4_present_hwtcl                               (0),
		.pf0_bar5_present_hwtcl                               (0),
		.pf0_exprom_bar_present_hwtcl                         (0),
		.pf0_bar0_type_hwtcl                                  (1),
		.pf0_bar2_type_hwtcl                                  (1),
		.pf0_bar4_type_hwtcl                                  (1),
		.pf0_bar0_prefetchable_hwtcl                          (1),
		.pf0_bar1_prefetchable_hwtcl                          (1),
		.pf0_bar2_prefetchable_hwtcl                          (1),
		.pf0_bar3_prefetchable_hwtcl                          (1),
		.pf0_bar4_prefetchable_hwtcl                          (1),
		.pf0_bar5_prefetchable_hwtcl                          (1),
		.pf0_bar0_size_hwtcl                                  (12),
		.pf0_bar1_size_hwtcl                                  (12),
		.pf0_bar2_size_hwtcl                                  (12),
		.pf0_bar3_size_hwtcl                                  (12),
		.pf0_bar4_size_hwtcl                                  (12),
		.pf0_bar5_size_hwtcl                                  (12),
		.pf0_exprom_bar_size_hwtcl                            (12),
		.pf0_vf_bar0_present_hwtcl                            (0),
		.pf0_vf_bar1_present_hwtcl                            (0),
		.pf0_vf_bar2_present_hwtcl                            (0),
		.pf0_vf_bar3_present_hwtcl                            (0),
		.pf0_vf_bar4_present_hwtcl                            (0),
		.pf0_vf_bar5_present_hwtcl                            (0),
		.pf0_vf_bar0_type_hwtcl                               (1),
		.pf0_vf_bar2_type_hwtcl                               (1),
		.pf0_vf_bar4_type_hwtcl                               (1),
		.pf0_vf_bar0_prefetchable_hwtcl                       (1),
		.pf0_vf_bar1_prefetchable_hwtcl                       (1),
		.pf0_vf_bar2_prefetchable_hwtcl                       (1),
		.pf0_vf_bar3_prefetchable_hwtcl                       (1),
		.pf0_vf_bar4_prefetchable_hwtcl                       (1),
		.pf0_vf_bar5_prefetchable_hwtcl                       (1),
		.pf0_vf_bar0_size_hwtcl                               (12),
		.pf0_vf_bar1_size_hwtcl                               (12),
		.pf0_vf_bar2_size_hwtcl                               (12),
		.pf0_vf_bar3_size_hwtcl                               (12),
		.pf0_vf_bar4_size_hwtcl                               (12),
		.pf0_vf_bar5_size_hwtcl                               (12),
		.pf1_bar0_present_hwtcl                               (0),
		.pf1_bar1_present_hwtcl                               (0),
		.pf1_bar2_present_hwtcl                               (0),
		.pf1_bar3_present_hwtcl                               (0),
		.pf1_bar4_present_hwtcl                               (0),
		.pf1_bar5_present_hwtcl                               (0),
		.pf1_exprom_bar_present_hwtcl                         (0),
		.pf1_bar0_type_hwtcl                                  (1),
		.pf1_bar2_type_hwtcl                                  (1),
		.pf1_bar4_type_hwtcl                                  (1),
		.pf1_bar0_prefetchable_hwtcl                          (1),
		.pf1_bar1_prefetchable_hwtcl                          (1),
		.pf1_bar2_prefetchable_hwtcl                          (1),
		.pf1_bar3_prefetchable_hwtcl                          (1),
		.pf1_bar4_prefetchable_hwtcl                          (1),
		.pf1_bar5_prefetchable_hwtcl                          (1),
		.pf1_bar0_size_hwtcl                                  (12),
		.pf1_bar1_size_hwtcl                                  (12),
		.pf1_bar2_size_hwtcl                                  (12),
		.pf1_bar3_size_hwtcl                                  (12),
		.pf1_bar4_size_hwtcl                                  (12),
		.pf1_bar5_size_hwtcl                                  (12),
		.pf1_exprom_bar_size_hwtcl                            (12),
		.pf1_vf_bar0_present_hwtcl                            (0),
		.pf1_vf_bar1_present_hwtcl                            (0),
		.pf1_vf_bar2_present_hwtcl                            (0),
		.pf1_vf_bar3_present_hwtcl                            (0),
		.pf1_vf_bar4_present_hwtcl                            (0),
		.pf1_vf_bar5_present_hwtcl                            (0),
		.pf1_vf_bar0_type_hwtcl                               (1),
		.pf1_vf_bar2_type_hwtcl                               (1),
		.pf1_vf_bar4_type_hwtcl                               (1),
		.pf1_vf_bar0_prefetchable_hwtcl                       (1),
		.pf1_vf_bar1_prefetchable_hwtcl                       (1),
		.pf1_vf_bar2_prefetchable_hwtcl                       (1),
		.pf1_vf_bar3_prefetchable_hwtcl                       (1),
		.pf1_vf_bar4_prefetchable_hwtcl                       (1),
		.pf1_vf_bar5_prefetchable_hwtcl                       (1),
		.pf1_vf_bar0_size_hwtcl                               (12),
		.pf1_vf_bar1_size_hwtcl                               (12),
		.pf1_vf_bar2_size_hwtcl                               (12),
		.pf1_vf_bar3_size_hwtcl                               (12),
		.pf1_vf_bar4_size_hwtcl                               (12),
		.pf1_vf_bar5_size_hwtcl                               (12),
		.pf2_bar0_present_hwtcl                               (0),
		.pf2_bar1_present_hwtcl                               (0),
		.pf2_bar2_present_hwtcl                               (0),
		.pf2_bar3_present_hwtcl                               (0),
		.pf2_bar4_present_hwtcl                               (0),
		.pf2_bar5_present_hwtcl                               (0),
		.pf2_exprom_bar_present_hwtcl                         (0),
		.pf2_bar0_type_hwtcl                                  (1),
		.pf2_bar2_type_hwtcl                                  (1),
		.pf2_bar4_type_hwtcl                                  (1),
		.pf2_bar0_prefetchable_hwtcl                          (1),
		.pf2_bar1_prefetchable_hwtcl                          (1),
		.pf2_bar2_prefetchable_hwtcl                          (1),
		.pf2_bar3_prefetchable_hwtcl                          (1),
		.pf2_bar4_prefetchable_hwtcl                          (1),
		.pf2_bar5_prefetchable_hwtcl                          (1),
		.pf2_bar0_size_hwtcl                                  (12),
		.pf2_bar1_size_hwtcl                                  (12),
		.pf2_bar2_size_hwtcl                                  (12),
		.pf2_bar3_size_hwtcl                                  (12),
		.pf2_bar4_size_hwtcl                                  (12),
		.pf2_bar5_size_hwtcl                                  (12),
		.pf2_exprom_bar_size_hwtcl                            (12),
		.pf2_vf_bar0_present_hwtcl                            (0),
		.pf2_vf_bar1_present_hwtcl                            (0),
		.pf2_vf_bar2_present_hwtcl                            (0),
		.pf2_vf_bar3_present_hwtcl                            (0),
		.pf2_vf_bar4_present_hwtcl                            (0),
		.pf2_vf_bar5_present_hwtcl                            (0),
		.pf2_vf_bar0_type_hwtcl                               (1),
		.pf2_vf_bar2_type_hwtcl                               (1),
		.pf2_vf_bar4_type_hwtcl                               (1),
		.pf2_vf_bar0_prefetchable_hwtcl                       (1),
		.pf2_vf_bar1_prefetchable_hwtcl                       (1),
		.pf2_vf_bar2_prefetchable_hwtcl                       (1),
		.pf2_vf_bar3_prefetchable_hwtcl                       (1),
		.pf2_vf_bar4_prefetchable_hwtcl                       (1),
		.pf2_vf_bar5_prefetchable_hwtcl                       (1),
		.pf2_vf_bar0_size_hwtcl                               (12),
		.pf2_vf_bar1_size_hwtcl                               (12),
		.pf2_vf_bar2_size_hwtcl                               (12),
		.pf2_vf_bar3_size_hwtcl                               (12),
		.pf2_vf_bar4_size_hwtcl                               (12),
		.pf2_vf_bar5_size_hwtcl                               (12),
		.pf3_bar0_present_hwtcl                               (0),
		.pf3_bar1_present_hwtcl                               (0),
		.pf3_bar2_present_hwtcl                               (0),
		.pf3_bar3_present_hwtcl                               (0),
		.pf3_bar4_present_hwtcl                               (0),
		.pf3_bar5_present_hwtcl                               (0),
		.pf3_exprom_bar_present_hwtcl                         (0),
		.pf3_bar0_type_hwtcl                                  (1),
		.pf3_bar2_type_hwtcl                                  (1),
		.pf3_bar4_type_hwtcl                                  (1),
		.pf3_bar0_prefetchable_hwtcl                          (1),
		.pf3_bar1_prefetchable_hwtcl                          (1),
		.pf3_bar2_prefetchable_hwtcl                          (1),
		.pf3_bar3_prefetchable_hwtcl                          (1),
		.pf3_bar4_prefetchable_hwtcl                          (1),
		.pf3_bar5_prefetchable_hwtcl                          (1),
		.pf3_bar0_size_hwtcl                                  (12),
		.pf3_bar1_size_hwtcl                                  (12),
		.pf3_bar2_size_hwtcl                                  (12),
		.pf3_bar3_size_hwtcl                                  (12),
		.pf3_bar4_size_hwtcl                                  (12),
		.pf3_bar5_size_hwtcl                                  (12),
		.pf3_exprom_bar_size_hwtcl                            (12),
		.pf3_vf_bar0_present_hwtcl                            (0),
		.pf3_vf_bar1_present_hwtcl                            (0),
		.pf3_vf_bar2_present_hwtcl                            (0),
		.pf3_vf_bar3_present_hwtcl                            (0),
		.pf3_vf_bar4_present_hwtcl                            (0),
		.pf3_vf_bar5_present_hwtcl                            (0),
		.pf3_vf_bar0_type_hwtcl                               (1),
		.pf3_vf_bar2_type_hwtcl                               (1),
		.pf3_vf_bar4_type_hwtcl                               (1),
		.pf3_vf_bar0_prefetchable_hwtcl                       (1),
		.pf3_vf_bar1_prefetchable_hwtcl                       (1),
		.pf3_vf_bar2_prefetchable_hwtcl                       (1),
		.pf3_vf_bar3_prefetchable_hwtcl                       (1),
		.pf3_vf_bar4_prefetchable_hwtcl                       (1),
		.pf3_vf_bar5_prefetchable_hwtcl                       (1),
		.pf3_vf_bar0_size_hwtcl                               (12),
		.pf3_vf_bar1_size_hwtcl                               (12),
		.pf3_vf_bar2_size_hwtcl                               (12),
		.pf3_vf_bar3_size_hwtcl                               (12),
		.pf3_vf_bar4_size_hwtcl                               (12),
		.pf3_vf_bar5_size_hwtcl                               (12),
		.pf4_bar0_present_hwtcl                               (0),
		.pf4_bar1_present_hwtcl                               (0),
		.pf4_bar2_present_hwtcl                               (0),
		.pf4_bar3_present_hwtcl                               (0),
		.pf4_bar4_present_hwtcl                               (0),
		.pf4_bar5_present_hwtcl                               (0),
		.pf4_exprom_bar_present_hwtcl                         (0),
		.pf4_bar0_type_hwtcl                                  (1),
		.pf4_bar2_type_hwtcl                                  (1),
		.pf4_bar4_type_hwtcl                                  (1),
		.pf4_bar0_prefetchable_hwtcl                          (1),
		.pf4_bar1_prefetchable_hwtcl                          (1),
		.pf4_bar2_prefetchable_hwtcl                          (1),
		.pf4_bar3_prefetchable_hwtcl                          (1),
		.pf4_bar4_prefetchable_hwtcl                          (1),
		.pf4_bar5_prefetchable_hwtcl                          (1),
		.pf4_bar0_size_hwtcl                                  (12),
		.pf4_bar1_size_hwtcl                                  (12),
		.pf4_bar2_size_hwtcl                                  (12),
		.pf4_bar3_size_hwtcl                                  (12),
		.pf4_bar4_size_hwtcl                                  (12),
		.pf4_bar5_size_hwtcl                                  (12),
		.pf4_exprom_bar_size_hwtcl                            (12),
		.pf5_bar0_present_hwtcl                               (0),
		.pf5_bar1_present_hwtcl                               (0),
		.pf5_bar2_present_hwtcl                               (0),
		.pf5_bar3_present_hwtcl                               (0),
		.pf5_bar4_present_hwtcl                               (0),
		.pf5_bar5_present_hwtcl                               (0),
		.pf5_exprom_bar_present_hwtcl                         (0),
		.pf5_bar0_type_hwtcl                                  (1),
		.pf5_bar2_type_hwtcl                                  (1),
		.pf5_bar4_type_hwtcl                                  (1),
		.pf5_bar0_prefetchable_hwtcl                          (1),
		.pf5_bar1_prefetchable_hwtcl                          (1),
		.pf5_bar2_prefetchable_hwtcl                          (1),
		.pf5_bar3_prefetchable_hwtcl                          (1),
		.pf5_bar4_prefetchable_hwtcl                          (1),
		.pf5_bar5_prefetchable_hwtcl                          (1),
		.pf5_bar0_size_hwtcl                                  (12),
		.pf5_bar1_size_hwtcl                                  (12),
		.pf5_bar2_size_hwtcl                                  (12),
		.pf5_bar3_size_hwtcl                                  (12),
		.pf5_bar4_size_hwtcl                                  (12),
		.pf5_bar5_size_hwtcl                                  (12),
		.pf5_exprom_bar_size_hwtcl                            (12),
		.pf6_bar0_present_hwtcl                               (0),
		.pf6_bar1_present_hwtcl                               (0),
		.pf6_bar2_present_hwtcl                               (0),
		.pf6_bar3_present_hwtcl                               (0),
		.pf6_bar4_present_hwtcl                               (0),
		.pf6_bar5_present_hwtcl                               (0),
		.pf6_exprom_bar_present_hwtcl                         (0),
		.pf6_bar0_type_hwtcl                                  (1),
		.pf6_bar2_type_hwtcl                                  (1),
		.pf6_bar4_type_hwtcl                                  (1),
		.pf6_bar0_prefetchable_hwtcl                          (1),
		.pf6_bar1_prefetchable_hwtcl                          (1),
		.pf6_bar2_prefetchable_hwtcl                          (1),
		.pf6_bar3_prefetchable_hwtcl                          (1),
		.pf6_bar4_prefetchable_hwtcl                          (1),
		.pf6_bar5_prefetchable_hwtcl                          (1),
		.pf6_bar0_size_hwtcl                                  (12),
		.pf6_bar1_size_hwtcl                                  (12),
		.pf6_bar2_size_hwtcl                                  (12),
		.pf6_bar3_size_hwtcl                                  (12),
		.pf6_bar4_size_hwtcl                                  (12),
		.pf6_bar5_size_hwtcl                                  (12),
		.pf6_exprom_bar_size_hwtcl                            (12),
		.pf7_bar0_present_hwtcl                               (0),
		.pf7_bar1_present_hwtcl                               (0),
		.pf7_bar2_present_hwtcl                               (0),
		.pf7_bar3_present_hwtcl                               (0),
		.pf7_bar4_present_hwtcl                               (0),
		.pf7_bar5_present_hwtcl                               (0),
		.pf7_exprom_bar_present_hwtcl                         (0),
		.pf7_bar0_type_hwtcl                                  (1),
		.pf7_bar2_type_hwtcl                                  (1),
		.pf7_bar4_type_hwtcl                                  (1),
		.pf7_bar0_prefetchable_hwtcl                          (1),
		.pf7_bar1_prefetchable_hwtcl                          (1),
		.pf7_bar2_prefetchable_hwtcl                          (1),
		.pf7_bar3_prefetchable_hwtcl                          (1),
		.pf7_bar4_prefetchable_hwtcl                          (1),
		.pf7_bar5_prefetchable_hwtcl                          (1),
		.pf7_bar0_size_hwtcl                                  (12),
		.pf7_bar1_size_hwtcl                                  (12),
		.pf7_bar2_size_hwtcl                                  (12),
		.pf7_bar3_size_hwtcl                                  (12),
		.pf7_bar4_size_hwtcl                                  (12),
		.pf7_bar5_size_hwtcl                                  (12),
		.pf7_exprom_bar_size_hwtcl                            (12),
		.pf1_vendor_id_hwtcl                                  (0),
		.pf1_device_id_hwtcl                                  (0),
		.pf1_vf_device_id_hwtcl                               (0),
		.pf1_revision_id_hwtcl                                (0),
		.pf1_class_code_hwtcl                                 (0),
		.pf1_subclass_code_hwtcl                              (0),
		.pf1_pci_prog_intfc_byte_hwtcl                        (0),
		.pf1_subsystem_vendor_id_hwtcl                        (0),
		.pf1_subsystem_device_id_hwtcl                        (0),
		.pf1_vf_subsystem_device_id_hwtcl                     (0),
		.pf2_vendor_id_hwtcl                                  (0),
		.pf2_device_id_hwtcl                                  (0),
		.pf2_vf_device_id_hwtcl                               (0),
		.pf2_revision_id_hwtcl                                (0),
		.pf2_class_code_hwtcl                                 (0),
		.pf2_subclass_code_hwtcl                              (0),
		.pf2_pci_prog_intfc_byte_hwtcl                        (0),
		.pf2_subsystem_vendor_id_hwtcl                        (0),
		.pf2_subsystem_device_id_hwtcl                        (0),
		.pf2_vf_subsystem_device_id_hwtcl                     (0),
		.pf3_vendor_id_hwtcl                                  (0),
		.pf3_device_id_hwtcl                                  (0),
		.pf3_vf_device_id_hwtcl                               (0),
		.pf3_revision_id_hwtcl                                (0),
		.pf3_class_code_hwtcl                                 (0),
		.pf3_subclass_code_hwtcl                              (0),
		.pf3_pci_prog_intfc_byte_hwtcl                        (0),
		.pf3_subsystem_vendor_id_hwtcl                        (0),
		.pf3_subsystem_device_id_hwtcl                        (0),
		.pf3_vf_subsystem_device_id_hwtcl                     (0),
		.pf4_vendor_id_hwtcl                                  (0),
		.pf4_device_id_hwtcl                                  (0),
		.pf4_vf_device_id_hwtcl                               (0),
		.pf4_revision_id_hwtcl                                (0),
		.pf4_class_code_hwtcl                                 (0),
		.pf4_subclass_code_hwtcl                              (0),
		.pf4_pci_prog_intfc_byte_hwtcl                        (0),
		.pf4_subsystem_vendor_id_hwtcl                        (0),
		.pf4_subsystem_device_id_hwtcl                        (0),
		.pf4_vf_subsystem_device_id_hwtcl                     (0),
		.pf5_vendor_id_hwtcl                                  (0),
		.pf5_device_id_hwtcl                                  (0),
		.pf5_vf_device_id_hwtcl                               (0),
		.pf5_revision_id_hwtcl                                (0),
		.pf5_class_code_hwtcl                                 (0),
		.pf5_subclass_code_hwtcl                              (0),
		.pf5_pci_prog_intfc_byte_hwtcl                        (0),
		.pf5_subsystem_vendor_id_hwtcl                        (0),
		.pf5_subsystem_device_id_hwtcl                        (0),
		.pf5_vf_subsystem_device_id_hwtcl                     (0),
		.pf6_vendor_id_hwtcl                                  (0),
		.pf6_device_id_hwtcl                                  (0),
		.pf6_vf_device_id_hwtcl                               (0),
		.pf6_revision_id_hwtcl                                (0),
		.pf6_class_code_hwtcl                                 (0),
		.pf6_subclass_code_hwtcl                              (0),
		.pf6_pci_prog_intfc_byte_hwtcl                        (0),
		.pf6_subsystem_vendor_id_hwtcl                        (0),
		.pf6_subsystem_device_id_hwtcl                        (0),
		.pf6_vf_subsystem_device_id_hwtcl                     (0),
		.pf7_vendor_id_hwtcl                                  (0),
		.pf7_device_id_hwtcl                                  (0),
		.pf7_vf_device_id_hwtcl                               (0),
		.pf7_revision_id_hwtcl                                (0),
		.pf7_class_code_hwtcl                                 (0),
		.pf7_subclass_code_hwtcl                              (0),
		.pf7_pci_prog_intfc_byte_hwtcl                        (0),
		.pf7_subsystem_vendor_id_hwtcl                        (0),
		.pf7_subsystem_device_id_hwtcl                        (0),
		.pf7_vf_subsystem_device_id_hwtcl                     (0),
		.pf_msi_support_hwtcl                                 (0),
		.pf0_msi_multi_message_capable_hwtcl                  (4),
		.pf1_msi_multi_message_capable_hwtcl                  (4),
		.pf2_msi_multi_message_capable_hwtcl                  (4),
		.pf3_msi_multi_message_capable_hwtcl                  (4),
		.pf4_msi_multi_message_capable_hwtcl                  (4),
		.pf5_msi_multi_message_capable_hwtcl                  (4),
		.pf6_msi_multi_message_capable_hwtcl                  (4),
		.pf7_msi_multi_message_capable_hwtcl                  (4),
		.pf_enable_function_msix_support_hwtcl                (0),
		.vf_msix_cap_present_hwtcl                            (0),
		.pf0_msix_table_size_hwtcl                            (0),
		.pf0_msix_table_offset_hwtcl                          (0),
		.pf0_msix_table_bir_hwtcl                             (0),
		.pf0_msix_pba_offset_hwtcl                            (0),
		.pf0_msix_pba_bir_hwtcl                               (0),
		.pf1_msix_table_size_hwtcl                            (0),
		.pf1_msix_table_offset_hwtcl                          (0),
		.pf1_msix_table_bir_hwtcl                             (0),
		.pf1_msix_pba_offset_hwtcl                            (0),
		.pf1_msix_pba_bir_hwtcl                               (0),
		.pf2_msix_table_size_hwtcl                            (0),
		.pf2_msix_table_offset_hwtcl                          (0),
		.pf2_msix_table_bir_hwtcl                             (0),
		.pf2_msix_pba_offset_hwtcl                            (0),
		.pf2_msix_pba_bir_hwtcl                               (0),
		.pf3_msix_table_size_hwtcl                            (0),
		.pf3_msix_table_offset_hwtcl                          (0),
		.pf3_msix_table_bir_hwtcl                             (0),
		.pf3_msix_pba_offset_hwtcl                            (0),
		.pf3_msix_pba_bir_hwtcl                               (0),
		.pf4_msix_table_size_hwtcl                            (0),
		.pf4_msix_table_offset_hwtcl                          (0),
		.pf4_msix_table_bir_hwtcl                             (0),
		.pf4_msix_pba_offset_hwtcl                            (0),
		.pf4_msix_pba_bir_hwtcl                               (0),
		.pf5_msix_table_size_hwtcl                            (0),
		.pf5_msix_table_offset_hwtcl                          (0),
		.pf5_msix_table_bir_hwtcl                             (0),
		.pf5_msix_pba_offset_hwtcl                            (0),
		.pf5_msix_pba_bir_hwtcl                               (0),
		.pf6_msix_table_size_hwtcl                            (0),
		.pf6_msix_table_offset_hwtcl                          (0),
		.pf6_msix_table_bir_hwtcl                             (0),
		.pf6_msix_pba_offset_hwtcl                            (0),
		.pf6_msix_pba_bir_hwtcl                               (0),
		.pf7_msix_table_size_hwtcl                            (0),
		.pf7_msix_table_offset_hwtcl                          (0),
		.pf7_msix_table_bir_hwtcl                             (0),
		.pf7_msix_pba_offset_hwtcl                            (0),
		.pf7_msix_pba_bir_hwtcl                               (0),
		.pf0_vf_msix_tbl_size_hwtcl                           (0),
		.pf0_vf_msix_tbl_offset_hwtcl                         (0),
		.pf0_vf_msix_tbl_bir_hwtcl                            (0),
		.pf0_vf_msix_pba_offset_hwtcl                         (0),
		.pf0_vf_msix_pba_bir_hwtcl                            (0),
		.pf1_vf_msix_tbl_size_hwtcl                           (0),
		.pf1_vf_msix_tbl_offset_hwtcl                         (0),
		.pf1_vf_msix_tbl_bir_hwtcl                            (0),
		.pf1_vf_msix_pba_offset_hwtcl                         (0),
		.pf1_vf_msix_pba_bir_hwtcl                            (0),
		.pf2_vf_msix_tbl_size_hwtcl                           (0),
		.pf2_vf_msix_tbl_offset_hwtcl                         (0),
		.pf2_vf_msix_tbl_bir_hwtcl                            (0),
		.pf2_vf_msix_pba_offset_hwtcl                         (0),
		.pf2_vf_msix_pba_bir_hwtcl                            (0),
		.pf3_vf_msix_tbl_size_hwtcl                           (0),
		.pf3_vf_msix_tbl_offset_hwtcl                         (0),
		.pf3_vf_msix_tbl_bir_hwtcl                            (0),
		.pf3_vf_msix_pba_offset_hwtcl                         (0),
		.pf3_vf_msix_pba_bir_hwtcl                            (0),
		.pf0_interrupt_pin_hwtcl                              ("inta"),
		.pf1_interrupt_pin_hwtcl                              ("inta"),
		.pf2_interrupt_pin_hwtcl                              ("inta"),
		.pf3_interrupt_pin_hwtcl                              ("inta"),
		.pf4_interrupt_pin_hwtcl                              ("inta"),
		.pf5_interrupt_pin_hwtcl                              ("inta"),
		.pf6_interrupt_pin_hwtcl                              ("inta"),
		.pf7_interrupt_pin_hwtcl                              ("inta"),
		.pf0_intr_line_hwtcl                                  (0),
		.pf1_intr_line_hwtcl                                  (0),
		.pf2_intr_line_hwtcl                                  (0),
		.pf3_intr_line_hwtcl                                  (0),
		.pf4_intr_line_hwtcl                                  (0),
		.pf5_intr_line_hwtcl                                  (0),
		.pf6_intr_line_hwtcl                                  (0),
		.pf7_intr_line_hwtcl                                  (0),
		.link2csr_width_hwtcl                                 (16),
		.lmi_width_hwtcl                                      (8),
		.rx_polinv_soft_logic_enable                          (0),
		.enable_soft_dfe                                      (0),
		.ceb_enable_hwtcl                                     (0),
		.ceb_pf_std_cap_last_ptr                              (0),
		.ceb_pf_ext_cap_last_ptr                              (0),
		.ceb_vf_std_cap_last_ptr                              (0),
		.ceb_vf_ext_cap_last_ptr                              (0),
		.ceb_ack_latency_hwtcl                                (1),
		.tlp_inspector_hwtcl                                  (0),
		.tlp_inspector_use_signal_probe_hwtcl                 (0),
		.tlp_inspector_use_thin_rx_master                     (0),
		.tlp_insp_trg_dw0_hwtcl                               (2049),
		.tlp_insp_trg_dw1_hwtcl                               (0),
		.tlp_insp_trg_dw2_hwtcl                               (0),
		.enable_ast_trs_hwtcl                                 (0),
		.ast_trs_num_desc_hwtcl                               (16),
		.ast_trs_txdata_width_hwtcl                           (256),
		.ast_trs_txdesc_width_hwtcl                           (256),
		.ast_trs_txstatus_width_hwtcl                         (256),
		.ast_trs_rxdata_width_hwtcl                           (256),
		.ast_trs_rxdesc_width_hwtcl                           (256),
		.ast_trs_txmty_width_hwtcl                            (32),
		.ast_trs_rxmty_width_hwtcl                            (32),
		.dma_use_scfifo_ext_hwtcl                             (0),
		.silicon_rev                                          ("20nm5es"),
		.hip_ac_pwr_clk_freq_in_hz                            (125000000),
		.ko_compl_data                                        (440),
		.ko_compl_header                                      (112),
		.acknack_base                                         (0),
		.acknack_set                                          ("false"),
		.advance_error_reporting                              ("disable"),
		.app_interface_width                                  ("avst_128bit"),
		.arb_upfc_30us_counter                                (0),
		.arb_upfc_30us_en                                     ("enable"),
		.aspm_config_management                               ("true"),
		.aspm_patch_disable                                   ("enable_both"),
		.ast_width_rx                                         ("rx_128"),
		.ast_width_tx                                         ("tx_128"),
		.atomic_malformed                                     ("false"),
		.atomic_op_completer_32bit                            ("false"),
		.atomic_op_completer_64bit                            ("false"),
		.atomic_op_routing                                    ("false"),
		.auto_msg_drop_enable                                 ("false"),
		.bar0_type                                            ("bar0_64bit_prefetch_mem"),
		.bar1_type                                            ("bar1_disable"),
		.bar2_type                                            ("bar2_64bit_prefetch_mem"),
		.bar3_type                                            ("bar3_disable"),
		.bar4_type                                            ("bar4_disable"),
		.bar5_type                                            ("bar5_disable"),
		.base_counter_sel                                     ("count_clk_62p5"),
		.bist_memory_settings                                 ("2417851639246850506078208"),
		.bridge_port_ssid_support                             ("false"),
		.bridge_port_vga_enable                               ("false"),
		.bypass_cdc                                           ("false"),
		.bypass_clk_switch                                    ("false"),
		.bypass_tl                                            ("false"),
		.cas_completer_128bit                                 ("false"),
		.cdc_clk_relation                                     ("plesiochronous"),
		.cdc_dummy_insert_limit                               (11),
		.cfg_parchk_ena                                       ("disable"),
		.cfgbp_req_recov_disable                              ("false"),
		.class_code                                           (16711680),
		.clock_pwr_management                                 ("false"),
		.completion_timeout                                   ("none_compl_timeout"),
		.core_clk_divider                                     ("div_2"),
		.core_clk_freq_mhz                                    ("core_clk_125mhz"),
		.core_clk_out_sel                                     ("core_clk_out_div_2"),
		.core_clk_sel                                         ("pld_clk"),
		.core_clk_source                                      ("pll_fixed_clk"),
		.cseb_bar_match_checking                              ("enable"),
		.cseb_config_bypass                                   ("disable"),
		.cseb_cpl_status_during_cvp                           ("config_retry_status"),
		.cseb_cpl_tag_checking                                ("enable"),
		.cseb_disable_auto_crs                                ("false"),
		.cseb_extend_pci                                      ("false"),
		.cseb_extend_pcie                                     ("false"),
		.cseb_min_error_checking                              ("false"),
		.cseb_route_to_avl_rx_st                              ("cseb"),
		.cseb_temp_busy_crs                                   ("completer_abort_tmp_busy"),
		.cvp_clk_reset                                        ("false"),
		.cvp_data_compressed                                  ("false"),
		.cvp_data_encrypted                                   ("false"),
		.cvp_enable                                           ("cvp_dis"),
		.cvp_mode_reset                                       ("false"),
		.cvp_rate_sel                                         ("full_rate"),
		.d0_pme                                               ("false"),
		.d1_pme                                               ("false"),
		.d1_support                                           ("false"),
		.d2_pme                                               ("false"),
		.d2_support                                           ("false"),
		.d3_cold_pme                                          ("false"),
		.d3_hot_pme                                           ("false"),
		.data_pack_rx                                         ("disable"),
		.deemphasis_enable                                    ("false"),
		.deskew_comma                                         ("skp_eieos_deskw"),
		.device_id                                            (0),
		.device_number                                        (0),
		.device_specific_init                                 ("false"),
		.dft_clock_obsrv_en                                   ("disable"),
		.dft_clock_obsrv_sel                                  ("dft_pclk"),
		.diffclock_nfts_count                                 (128),
		.dis_cplovf                                           ("disable"),
		.dis_paritychk                                        ("disable"),
		.disable_link_x2_support                              ("false"),
		.disable_snoop_packet                                 ("false"),
		.dl_tx_check_parity_edb                               ("disable"),
		.dll_active_report_support                            ("false"),
		.early_dl_up                                          ("false"),
		.ecrc_check_capable                                   ("false"),
		.ecrc_gen_capable                                     ("false"),
		.egress_block_err_report_ena                          ("false"),
		.ei_delay_powerdown_count                             (10),
		.eie_before_nfts_count                                (4),
		.electromech_interlock                                ("false"),
		.en_ieiupdatefc                                       ("false"),
		.en_lane_errchk                                       ("false"),
		.en_phystatus_dly                                     ("false"),
		.ena_ido_cpl                                          ("false"),
		.ena_ido_req                                          ("false"),
		.enable_adapter_half_rate_mode                        ("false"),
		.enable_ch0_pclk_out                                  ("pclk_central"),
		.enable_ch01_pclk_out                                 ("pclk_ch0"),
		.enable_completion_timeout_disable                    ("true"),
		.enable_directed_spd_chng                             ("false"),
		.enable_function_msix_support                         ("false"),
		.enable_l0s_aspm                                      ("false"),
		.enable_l1_aspm                                       ("false"),
		.enable_rx_buffer_checking                            ("false"),
		.enable_rx_reordering                                 ("true"),
		.enable_slot_register                                 ("false"),
		.endpoint_l0_latency                                  (0),
		.endpoint_l1_latency                                  (0),
		.eql_rq_int_en_number                                 (0),
		.errmgt_fcpe_patch_dis                                ("enable"),
		.errmgt_fep_patch_dis                                 ("enable"),
		.extend_tag_field                                     ("false"),
		.extended_format_field                                ("true"),
		.extended_tag_reset                                   ("false"),
		.fc_init_timer                                        (1024),
		.flow_control_timeout_count                           (200),
		.flow_control_update_count                            (30),
		.flr_capability                                       ("false"),
		.force_dis_to_det                                     ("false"),
		.force_gen1_dis                                       ("false"),
		.force_tx_coeff_preset_lpbk                           ("false"),
		.frame_err_patch_dis                                  ("enable"),
		.func_mode                                            ("enable"),
		.g3_bypass_equlz                                      ("false"),
		.g3_coeff_done_tmout                                  ("enable"),
		.g3_deskew_char                                       ("default_sdsos"),
		.g3_dis_be_frm_err                                    ("false"),
		.g3_dn_rx_hint_eqlz_0                                 (0),
		.g3_dn_rx_hint_eqlz_1                                 (0),
		.g3_dn_rx_hint_eqlz_2                                 (0),
		.g3_dn_rx_hint_eqlz_3                                 (0),
		.g3_dn_rx_hint_eqlz_4                                 (0),
		.g3_dn_rx_hint_eqlz_5                                 (0),
		.g3_dn_rx_hint_eqlz_6                                 (0),
		.g3_dn_rx_hint_eqlz_7                                 (0),
		.g3_dn_tx_preset_eqlz_0                               (0),
		.g3_dn_tx_preset_eqlz_1                               (0),
		.g3_dn_tx_preset_eqlz_2                               (0),
		.g3_dn_tx_preset_eqlz_3                               (0),
		.g3_dn_tx_preset_eqlz_4                               (0),
		.g3_dn_tx_preset_eqlz_5                               (0),
		.g3_dn_tx_preset_eqlz_6                               (0),
		.g3_dn_tx_preset_eqlz_7                               (0),
		.g3_force_ber_max                                     ("false"),
		.g3_force_ber_min                                     ("true"),
		.g3_lnk_trn_rx_ts                                     ("false"),
		.g3_ltssm_eq_dbg                                      ("false"),
		.g3_ltssm_rec_dbg                                     ("true"),
		.g3_pause_ltssm_rec_en                                ("disable"),
		.g3_quiesce_guarant                                   ("false"),
		.g3_redo_equlz_dis                                    ("false"),
		.g3_redo_equlz_en                                     ("false"),
		.g3_up_rx_hint_eqlz_0                                 (0),
		.g3_up_rx_hint_eqlz_1                                 (0),
		.g3_up_rx_hint_eqlz_2                                 (0),
		.g3_up_rx_hint_eqlz_3                                 (0),
		.g3_up_rx_hint_eqlz_4                                 (0),
		.g3_up_rx_hint_eqlz_5                                 (0),
		.g3_up_rx_hint_eqlz_6                                 (0),
		.g3_up_rx_hint_eqlz_7                                 (0),
		.g3_up_tx_preset_eqlz_0                               (0),
		.g3_up_tx_preset_eqlz_1                               (0),
		.g3_up_tx_preset_eqlz_2                               (0),
		.g3_up_tx_preset_eqlz_3                               (0),
		.g3_up_tx_preset_eqlz_4                               (0),
		.g3_up_tx_preset_eqlz_5                               (0),
		.g3_up_tx_preset_eqlz_6                               (0),
		.g3_up_tx_preset_eqlz_7                               (0),
		.gen123_lane_rate_mode                                ("gen1_gen2"),
		.gen2_diffclock_nfts_count                            (255),
		.gen2_pma_pll_usage                                   ("use_ffpll"),
		.gen2_sameclock_nfts_count                            (255),
		.gen3_coeff_1                                         (8),
		.gen3_coeff_1_ber_meas                                (4),
		.gen3_coeff_1_nxtber_less                             (1),
		.gen3_coeff_1_nxtber_more                             (1),
		.gen3_coeff_1_preset_hint                             (0),
		.gen3_coeff_1_reqber                                  (0),
		.gen3_coeff_1_sel                                     ("preset_1"),
		.gen3_coeff_10                                        (0),
		.gen3_coeff_10_ber_meas                               (0),
		.gen3_coeff_10_nxtber_less                            (0),
		.gen3_coeff_10_nxtber_more                            (0),
		.gen3_coeff_10_preset_hint                            (0),
		.gen3_coeff_10_reqber                                 (0),
		.gen3_coeff_10_sel                                    ("preset_10"),
		.gen3_coeff_11                                        (0),
		.gen3_coeff_11_ber_meas                               (0),
		.gen3_coeff_11_nxtber_less                            (0),
		.gen3_coeff_11_nxtber_more                            (0),
		.gen3_coeff_11_preset_hint                            (0),
		.gen3_coeff_11_reqber                                 (0),
		.gen3_coeff_11_sel                                    ("preset_11"),
		.gen3_coeff_12                                        (0),
		.gen3_coeff_12_ber_meas                               (0),
		.gen3_coeff_12_nxtber_less                            (0),
		.gen3_coeff_12_nxtber_more                            (0),
		.gen3_coeff_12_preset_hint                            (0),
		.gen3_coeff_12_reqber                                 (0),
		.gen3_coeff_12_sel                                    ("preset_12"),
		.gen3_coeff_13                                        (0),
		.gen3_coeff_13_ber_meas                               (0),
		.gen3_coeff_13_nxtber_less                            (0),
		.gen3_coeff_13_nxtber_more                            (0),
		.gen3_coeff_13_preset_hint                            (0),
		.gen3_coeff_13_reqber                                 (0),
		.gen3_coeff_13_sel                                    ("preset_13"),
		.gen3_coeff_14                                        (0),
		.gen3_coeff_14_ber_meas                               (0),
		.gen3_coeff_14_nxtber_less                            (0),
		.gen3_coeff_14_nxtber_more                            (0),
		.gen3_coeff_14_preset_hint                            (0),
		.gen3_coeff_14_reqber                                 (0),
		.gen3_coeff_14_sel                                    ("preset_14"),
		.gen3_coeff_15                                        (0),
		.gen3_coeff_15_ber_meas                               (0),
		.gen3_coeff_15_nxtber_less                            (0),
		.gen3_coeff_15_nxtber_more                            (0),
		.gen3_coeff_15_preset_hint                            (0),
		.gen3_coeff_15_reqber                                 (0),
		.gen3_coeff_15_sel                                    ("preset_15"),
		.gen3_coeff_16                                        (0),
		.gen3_coeff_16_ber_meas                               (0),
		.gen3_coeff_16_nxtber_less                            (0),
		.gen3_coeff_16_nxtber_more                            (0),
		.gen3_coeff_16_preset_hint                            (0),
		.gen3_coeff_16_reqber                                 (0),
		.gen3_coeff_16_sel                                    ("preset_16"),
		.gen3_coeff_17                                        (196608),
		.gen3_coeff_17_ber_meas                               (0),
		.gen3_coeff_17_nxtber_less                            (0),
		.gen3_coeff_17_nxtber_more                            (0),
		.gen3_coeff_17_preset_hint                            (0),
		.gen3_coeff_17_reqber                                 (0),
		.gen3_coeff_17_sel                                    ("preset_17"),
		.gen3_coeff_18                                        (196609),
		.gen3_coeff_18_ber_meas                               (0),
		.gen3_coeff_18_nxtber_less                            (0),
		.gen3_coeff_18_nxtber_more                            (0),
		.gen3_coeff_18_preset_hint                            (0),
		.gen3_coeff_18_reqber                                 (0),
		.gen3_coeff_18_sel                                    ("preset_18"),
		.gen3_coeff_19                                        (196609),
		.gen3_coeff_19_ber_meas                               (0),
		.gen3_coeff_19_nxtber_less                            (0),
		.gen3_coeff_19_nxtber_more                            (0),
		.gen3_coeff_19_preset_hint                            (0),
		.gen3_coeff_19_reqber                                 (0),
		.gen3_coeff_19_sel                                    ("preset_19"),
		.gen3_coeff_2                                         (8),
		.gen3_coeff_2_ber_meas                                (4),
		.gen3_coeff_2_nxtber_less                             (2),
		.gen3_coeff_2_nxtber_more                             (2),
		.gen3_coeff_2_preset_hint                             (7),
		.gen3_coeff_2_reqber                                  (0),
		.gen3_coeff_2_sel                                     ("preset_2"),
		.gen3_coeff_20                                        (196609),
		.gen3_coeff_20_ber_meas                               (0),
		.gen3_coeff_20_nxtber_less                            (0),
		.gen3_coeff_20_nxtber_more                            (0),
		.gen3_coeff_20_preset_hint                            (0),
		.gen3_coeff_20_reqber                                 (0),
		.gen3_coeff_20_sel                                    ("preset_20"),
		.gen3_coeff_21                                        (196609),
		.gen3_coeff_21_ber_meas                               (0),
		.gen3_coeff_21_nxtber_less                            (0),
		.gen3_coeff_21_nxtber_more                            (0),
		.gen3_coeff_21_preset_hint                            (0),
		.gen3_coeff_21_reqber                                 (0),
		.gen3_coeff_21_sel                                    ("preset_21"),
		.gen3_coeff_22                                        (196609),
		.gen3_coeff_22_ber_meas                               (0),
		.gen3_coeff_22_nxtber_less                            (7),
		.gen3_coeff_22_nxtber_more                            (0),
		.gen3_coeff_22_preset_hint                            (0),
		.gen3_coeff_22_reqber                                 (0),
		.gen3_coeff_22_sel                                    ("preset_22"),
		.gen3_coeff_23                                        (196609),
		.gen3_coeff_23_ber_meas                               (0),
		.gen3_coeff_23_nxtber_less                            (0),
		.gen3_coeff_23_nxtber_more                            (0),
		.gen3_coeff_23_preset_hint                            (0),
		.gen3_coeff_23_reqber                                 (0),
		.gen3_coeff_23_sel                                    ("preset_23"),
		.gen3_coeff_24                                        (196609),
		.gen3_coeff_24_ber_meas                               (0),
		.gen3_coeff_24_nxtber_less                            (0),
		.gen3_coeff_24_nxtber_more                            (0),
		.gen3_coeff_24_preset_hint                            (7),
		.gen3_coeff_24_reqber                                 (0),
		.gen3_coeff_24_sel                                    ("preset_24"),
		.gen3_coeff_3                                         (8),
		.gen3_coeff_3_ber_meas                                (16),
		.gen3_coeff_3_nxtber_less                             (4),
		.gen3_coeff_3_nxtber_more                             (4),
		.gen3_coeff_3_preset_hint                             (7),
		.gen3_coeff_3_reqber                                  (31),
		.gen3_coeff_3_sel                                     ("preset_3"),
		.gen3_coeff_4                                         (8),
		.gen3_coeff_4_ber_meas                                (4),
		.gen3_coeff_4_nxtber_less                             (4),
		.gen3_coeff_4_nxtber_more                             (4),
		.gen3_coeff_4_preset_hint                             (7),
		.gen3_coeff_4_reqber                                  (31),
		.gen3_coeff_4_sel                                     ("preset_4"),
		.gen3_coeff_5                                         (0),
		.gen3_coeff_5_ber_meas                                (0),
		.gen3_coeff_5_nxtber_less                             (0),
		.gen3_coeff_5_nxtber_more                             (0),
		.gen3_coeff_5_preset_hint                             (7),
		.gen3_coeff_5_reqber                                  (0),
		.gen3_coeff_5_sel                                     ("preset_5"),
		.gen3_coeff_6                                         (0),
		.gen3_coeff_6_ber_meas                                (0),
		.gen3_coeff_6_nxtber_less                             (0),
		.gen3_coeff_6_nxtber_more                             (0),
		.gen3_coeff_6_preset_hint                             (0),
		.gen3_coeff_6_reqber                                  (0),
		.gen3_coeff_6_sel                                     ("preset_6"),
		.gen3_coeff_7                                         (0),
		.gen3_coeff_7_ber_meas                                (0),
		.gen3_coeff_7_nxtber_less                             (0),
		.gen3_coeff_7_nxtber_more                             (0),
		.gen3_coeff_7_preset_hint                             (0),
		.gen3_coeff_7_reqber                                  (0),
		.gen3_coeff_7_sel                                     ("preset_7"),
		.gen3_coeff_8                                         (0),
		.gen3_coeff_8_ber_meas                                (0),
		.gen3_coeff_8_nxtber_less                             (0),
		.gen3_coeff_8_nxtber_more                             (0),
		.gen3_coeff_8_preset_hint                             (0),
		.gen3_coeff_8_reqber                                  (0),
		.gen3_coeff_8_sel                                     ("preset_8"),
		.gen3_coeff_9                                         (0),
		.gen3_coeff_9_ber_meas                                (0),
		.gen3_coeff_9_nxtber_less                             (0),
		.gen3_coeff_9_nxtber_more                             (0),
		.gen3_coeff_9_preset_hint                             (0),
		.gen3_coeff_9_reqber                                  (0),
		.gen3_coeff_9_sel                                     ("preset_9"),
		.gen3_coeff_delay_count                               (125),
		.gen3_coeff_errchk                                    ("disable"),
		.gen3_dcbal_en                                        ("true"),
		.gen3_diffclock_nfts_count                            (128),
		.gen3_force_local_coeff                               ("false"),
		.gen3_full_swing                                      (60),
		.gen3_half_swing                                      ("false"),
		.gen3_low_freq                                        (20),
		.gen3_paritychk                                       ("disable"),
		.gen3_pl_framing_err_dis                              ("enable"),
		.gen3_preset_coeff_1                                  (64320),
		.gen3_preset_coeff_10                                 (3210),
		.gen3_preset_coeff_11                                 (84480),
		.gen3_preset_coeff_2                                  (44160),
		.gen3_preset_coeff_3                                  (52224),
		.gen3_preset_coeff_4                                  (36096),
		.gen3_preset_coeff_5                                  (3840),
		.gen3_preset_coeff_6                                  (3462),
		.gen3_preset_coeff_7                                  (3336),
		.gen3_preset_coeff_8                                  (51846),
		.gen3_preset_coeff_9                                  (35592),
		.gen3_reset_eieos_cnt_bit                             ("false"),
		.gen3_rxfreqlock_counter                              (0),
		.gen3_sameclock_nfts_count                            (128),
		.gen3_scrdscr_bypass                                  ("true"),
		.gen3_skip_ph2_ph3                                    ("false"),
		.hard_reset_bypass                                    ("false"),
		.hard_rst_sig_chnl_en                                 ("enable_hrc_sig_x4"),
		.hard_rst_tx_pll_rst_chnl_en                          ("enable_hrc_txpll_rst_ch4"),
		.hip_base_address                                     (0),
		.hip_clock_dis                                        ("enable_hip_clk"),
		.hip_hard_reset                                       ("enable"),
		.hip_pcs_sig_chnl_en                                  ("enable_hip_pcs_sig_x4"),
		.hot_plug_support                                     (0),
		.hrc_chnl_txpll_master_cgb_rst_select                 ("ch3_master_cgb_sel"),
		.hrdrstctrl_en                                        ("hrdrstctrl_en"),
		.iei_enable_settings                                  ("gen3_infei_infsd_gen2_infsd_gen1_infsd_sd"),
		.indicator                                            (0),
		.intel_id_access                                      ("false"),
		.interrupt_pin                                        ("inta"),
		.io_window_addr_width                                 ("none"),
		.jtag_id                                              ("0"),
		.l0_exit_latency_diffclock                            (6),
		.l0_exit_latency_sameclock                            (6),
		.l01_entry_latency                                    (31),
		.l0s_adj_rply_timer_dis                               ("enable"),
		.l1_exit_latency_diffclock                            (0),
		.l1_exit_latency_sameclock                            (0),
		.l2_async_logic                                       ("disable"),
		.lane_mask                                            ("ln_mask_x4"),
		.lane_rate                                            ("gen2"),
		.link_width                                           ("x4"),
		.low_priority_vc                                      ("single_vc_low_pr"),
		.ltr_mechanism                                        ("false"),
		.ltssm_1ms_timeout                                    ("disable"),
		.ltssm_freqlocked_check                               ("disable"),
		.malformed_tlp_truncate_en                            ("disable"),
		.max_link_width                                       ("x4_link_width"),
		.max_payload_size                                     ("payload_128"),
		.maximum_current                                      (0),
		.millisecond_cycle_count                              (124248),
		.msi_64bit_addressing_capable                         ("true"),
		.msi_masking_capable                                  ("false"),
		.msi_multi_message_capable                            ("count_4"),
		.msi_support                                          ("true"),
		.msix_pba_bir                                         (0),
		.msix_table_bir                                       (0),
		.msix_table_size                                      (0),
		.national_inst_thru_enhance                           ("false"),
		.no_command_completed                                 ("false"),
		.no_soft_reset                                        ("false"),
		.pcie_base_spec                                       ("pcie_3p0"),
		.pcie_mode                                            ("ep_native"),
		.pcie_spec_1p0_compliance                             ("spec_1p1"),
		.pcie_spec_version                                    ("v3"),
		.pclk_out_sel                                         ("pclk"),
		.pld_in_use_reg                                       ("false"),
		.pm_latency_patch_dis                                 ("enable"),
		.pm_txdl_patch_dis                                    ("enable"),
		.pme_clock                                            ("false"),
		.port_link_number                                     (1),
		.port_type                                            ("native_ep"),
		.powerdown_mode                                       ("powerup"),
		.prefetchable_mem_window_addr_width                   ("prefetch_0"),
		.r2c_mask_easy                                        ("false"),
		.r2c_mask_enable                                      ("false"),
		.rec_frqlk_mon_en                                     ("disable"),
		.register_pipe_signals                                ("true"),
		.retry_buffer_last_active_address                     (1023),
		.retry_buffer_memory_settings                         ("12885005388"),
		.retry_ecc_corr_mask_dis                              ("enable"),
		.revision_id                                          (0),
		.role_based_error_reporting                           ("true"),
		.rp_bug_fix_pri_sec_stat_reg                          (127),
		.rpltim_base                                          (16),
		.rpltim_set                                           ("true"),
		.rstctl_ltssm_dis                                     ("false"),
		.rstctrl_1ms_count_fref_clk                           (100000),
		.rstctrl_1us_count_fref_clk                           (100),
		.rstctrl_altpe3_crst_n_inv                            ("false"),
		.rstctrl_altpe3_rst_n_inv                             ("false"),
		.rstctrl_altpe3_srst_n_inv                            ("false"),
		.rstctrl_chnl_cal_done_select                         ("ch0123_out_chnl_cal_done"),
		.rstctrl_debug_en                                     ("false"),
		.rstctrl_force_inactive_rst                           ("false"),
		.rstctrl_fref_clk_select                              ("ch0_sel"),
		.rstctrl_hard_block_enable                            ("hard_rst_ctl"),
		.rstctrl_hip_ep                                       ("hip_ep"),
		.rstctrl_mask_tx_pll_lock_select                      ("ch3_sel_mask_tx_pll_lock"),
		.rstctrl_perst_enable                                 ("level"),
		.rstctrl_perstn_select                                ("perstn_pin"),
		.rstctrl_pld_clr                                      ("true"),
		.rstctrl_pll_cal_done_select                          ("ch4_sel_pll_cal_done"),
		.rstctrl_rx_pcs_rst_n_inv                             ("false"),
		.rstctrl_rx_pcs_rst_n_select                          ("ch0123_out_rx_pcs_rst"),
		.rstctrl_rx_pll_freq_lock_select                      ("not_active_rx_pll_f_lock"),
		.rstctrl_rx_pll_lock_select                           ("ch0123_sel_rx_pll_lock"),
		.rstctrl_rx_pma_rstb_inv                              ("false"),
		.rstctrl_rx_pma_rstb_select                           ("ch0123_out_rx_pma_rstb"),
		.rstctrl_timer_a                                      (10),
		.rstctrl_timer_a_type                                 ("a_timer_fref_cycles"),
		.rstctrl_timer_b                                      (10),
		.rstctrl_timer_b_type                                 ("b_timer_fref_cycles"),
		.rstctrl_timer_c                                      (10),
		.rstctrl_timer_c_type                                 ("c_timer_fref_cycles"),
		.rstctrl_timer_d                                      (20),
		.rstctrl_timer_d_type                                 ("d_timer_fref_cycles"),
		.rstctrl_timer_e                                      (1),
		.rstctrl_timer_e_type                                 ("e_timer_fref_cycles"),
		.rstctrl_timer_f                                      (10),
		.rstctrl_timer_f_type                                 ("f_timer_fref_cycles"),
		.rstctrl_timer_g                                      (10),
		.rstctrl_timer_g_type                                 ("g_timer_fref_cycles"),
		.rstctrl_timer_h                                      (4),
		.rstctrl_timer_h_type                                 ("h_timer_micro_secs"),
		.rstctrl_timer_i                                      (20),
		.rstctrl_timer_i_type                                 ("i_timer_fref_cycles"),
		.rstctrl_timer_j                                      (20),
		.rstctrl_timer_j_type                                 ("j_timer_fref_cycles"),
		.rstctrl_tx_lcff_pll_lock_select                      ("ch4_sel_lcff_pll_lock"),
		.rstctrl_tx_lcff_pll_rstb_select                      ("ch4_out_lcff_pll_rstb"),
		.rstctrl_tx_pcs_rst_n_inv                             ("false"),
		.rstctrl_tx_pcs_rst_n_select                          ("ch0123_out_tx_pcs_rst"),
		.rstctrl_tx_pma_rstb_inv                              ("false"),
		.rstctrl_tx_pma_syncp_inv                             ("false"),
		.rstctrl_tx_pma_syncp_select                          ("ch3_out_tx_pma_syncp"),
		.rx_ast_parity                                        ("disable"),
		.rx_buffer_credit_alloc                               ("balance"),
		.rx_buffer_fc_protect                                 (68),
		.rx_buffer_protect                                    (68),
		.rx_cdc_almost_empty                                  (3),
		.rx_cdc_almost_full                                   (12),
		.rx_cred_ctl_param                                    ("disable"),
		.rx_ei_l0s                                            ("disable"),
		.rx_l0s_count_idl                                     (0),
		.rx_ptr0_nonposted_dpram_max                          (2047),
		.rx_ptr0_nonposted_dpram_min                          (1928),
		.rx_ptr0_posted_dpram_max                             (1927),
		.rx_ptr0_posted_dpram_min                             (0),
		.rx_runt_patch_dis                                    ("enable"),
		.rx_sop_ctrl                                          ("rx_sop_boundary_128"),
		.rx_trunc_patch_dis                                   ("enable"),
		.rx_use_prst                                          ("true"),
		.rx_use_prst_ep                                       ("true"),
		.rxbuf_ecc_corr_mask_dis                              ("enable"),
		.sameclock_nfts_count                                 (128),
		.sel_enable_pcs_rx_fifo_err                           ("disable_sel"),
		.sim_mode                                             ("disable"),
		.simple_ro_fifo_control_en                            ("disable"),
		.single_rx_detect                                     ("detect_lane0_3"),
		.skp_os_gen3_count                                    (0),
		.skp_os_schedule_count                                (0),
		.slot_number                                          (0),
		.slot_power_limit                                     (0),
		.slot_power_scale                                     (0),
		.slotclk_cfg                                          ("static_slotclkcfgon"),
		.ssid                                                 (0),
		.ssvid                                                (0),
		.subsystem_device_id                                  (0),
		.subsystem_vendor_id                                  (0),
		.sup_mode                                             ("user_mode"),
		.surprise_down_error_support                          ("false"),
		.tl_cfg_div                                           ("cfg_clk_div_7"),
		.tl_tx_check_parity_msg                               ("disable"),
		.tph_completer                                        ("false"),
		.tx_ast_parity                                        ("disable"),
		.tx_cdc_almost_empty                                  (5),
		.tx_cdc_almost_full                                   (11),
		.tx_sop_ctrl                                          ("boundary_128"),
		.tx_swing                                             (0),
		.txdl_fair_arbiter_counter                            (0),
		.txdl_fair_arbiter_en                                 ("enable"),
		.txrate_adv                                           ("capability"),
		.uc_calibration_en                                    ("uc_calibration_en"),
		.use_aer                                              ("false"),
		.use_crc_forwarding                                   ("false"),
		.user_id                                              (0),
		.vc_arbitration                                       ("single_vc_arb"),
		.vc_enable                                            ("single_vc"),
		.vc0_clk_enable                                       ("true"),
		.vc0_rx_buffer_memory_settings                        ("12885005388"),
		.vc0_rx_flow_ctrl_compl_data                          (0),
		.vc0_rx_flow_ctrl_compl_header                        (0),
		.vc0_rx_flow_ctrl_nonposted_data                      (0),
		.vc0_rx_flow_ctrl_nonposted_header                    (56),
		.vc0_rx_flow_ctrl_posted_data                         (358),
		.vc0_rx_flow_ctrl_posted_header                       (50),
		.vc1_clk_enable                                       ("false"),
		.vendor_id                                            (4466),
		.vsec_cap                                             (0),
		.vsec_id                                              (4466),
		.wrong_device_id                                      ("disable"),
		.not_use_k_gbl_bits                                   ("not_used_k_gbl"),
		.avmm_force_inter_sel_csr_ctrl                        ("disable"),
		.operating_voltage                                    ("standard"),
		.rxdl_bad_tlp_patch_dis                               ("rxdlbug2_enable_both"),
		.avmm_dprio_broadcast_en_csr_ctrl                     ("disable"),
		.hip_ac_pwr_uw_per_mhz                                (1120),
		.rxdl_bad_sop_eop_filter_dis                          ("rxdlbug1_enable_both"),
		.rxdl_lcrc_patch_dis                                  ("rxdlbug3_enable_both"),
		.capab_rate_rxcfg_en                                  ("disable"),
		.avmm_cvp_inter_sel_csr_ctrl                          ("disable"),
		.lmi_hold_off_cfg_timer_en                            ("disable"),
		.avmm_power_iso_en_csr_ctrl                           ("disable"),
		.eco_fb332688_dis                                     ("false")
	) pcie (
		.coreclkout_hip                 (coreclkout_hip),                                                                                                                                                                                                                                                        //  output,    width = 1,    coreclkout_hip.clk
		.refclk                         (refclk),                                                                                                                                                                                                                                                                //   input,    width = 1,            refclk.clk
		.npor                           (npor),                                                                                                                                                                                                                                                                  //   input,    width = 1,              npor.npor
		.pin_perst                      (pin_perst),                                                                                                                                                                                                                                                             //   input,    width = 1,                  .pin_perst
		.app_nreset_status              (app_nreset_status),                                                                                                                                                                                                                                                     //  output,    width = 1, app_nreset_status.reset_n
		.test_in                        (test_in),                                                                                                                                                                                                                                                               //   input,   width = 32,          hip_ctrl.test_in
		.simu_mode_pipe                 (simu_mode_pipe),                                                                                                                                                                                                                                                        //   input,    width = 1,                  .simu_mode_pipe
		.sim_pipe_pclk_in               (sim_pipe_pclk_in),                                                                                                                                                                                                                                                      //   input,    width = 1,          hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate                  (sim_pipe_rate),                                                                                                                                                                                                                                                         //  output,    width = 2,                  .sim_pipe_rate
		.sim_ltssmstate                 (sim_ltssmstate),                                                                                                                                                                                                                                                        //  output,    width = 5,                  .sim_ltssmstate
		.eidleinfersel0                 (eidleinfersel0),                                                                                                                                                                                                                                                        //  output,    width = 3,                  .eidleinfersel0
		.eidleinfersel1                 (eidleinfersel1),                                                                                                                                                                                                                                                        //  output,    width = 3,                  .eidleinfersel1
		.eidleinfersel2                 (eidleinfersel2),                                                                                                                                                                                                                                                        //  output,    width = 3,                  .eidleinfersel2
		.eidleinfersel3                 (eidleinfersel3),                                                                                                                                                                                                                                                        //  output,    width = 3,                  .eidleinfersel3
		.powerdown0                     (powerdown0),                                                                                                                                                                                                                                                            //  output,    width = 2,                  .powerdown0
		.powerdown1                     (powerdown1),                                                                                                                                                                                                                                                            //  output,    width = 2,                  .powerdown1
		.powerdown2                     (powerdown2),                                                                                                                                                                                                                                                            //  output,    width = 2,                  .powerdown2
		.powerdown3                     (powerdown3),                                                                                                                                                                                                                                                            //  output,    width = 2,                  .powerdown3
		.rxpolarity0                    (rxpolarity0),                                                                                                                                                                                                                                                           //  output,    width = 1,                  .rxpolarity0
		.rxpolarity1                    (rxpolarity1),                                                                                                                                                                                                                                                           //  output,    width = 1,                  .rxpolarity1
		.rxpolarity2                    (rxpolarity2),                                                                                                                                                                                                                                                           //  output,    width = 1,                  .rxpolarity2
		.rxpolarity3                    (rxpolarity3),                                                                                                                                                                                                                                                           //  output,    width = 1,                  .rxpolarity3
		.txcompl0                       (txcompl0),                                                                                                                                                                                                                                                              //  output,    width = 1,                  .txcompl0
		.txcompl1                       (txcompl1),                                                                                                                                                                                                                                                              //  output,    width = 1,                  .txcompl1
		.txcompl2                       (txcompl2),                                                                                                                                                                                                                                                              //  output,    width = 1,                  .txcompl2
		.txcompl3                       (txcompl3),                                                                                                                                                                                                                                                              //  output,    width = 1,                  .txcompl3
		.txdata0                        (txdata0),                                                                                                                                                                                                                                                               //  output,   width = 32,                  .txdata0
		.txdata1                        (txdata1),                                                                                                                                                                                                                                                               //  output,   width = 32,                  .txdata1
		.txdata2                        (txdata2),                                                                                                                                                                                                                                                               //  output,   width = 32,                  .txdata2
		.txdata3                        (txdata3),                                                                                                                                                                                                                                                               //  output,   width = 32,                  .txdata3
		.txdatak0                       (txdatak0),                                                                                                                                                                                                                                                              //  output,    width = 4,                  .txdatak0
		.txdatak1                       (txdatak1),                                                                                                                                                                                                                                                              //  output,    width = 4,                  .txdatak1
		.txdatak2                       (txdatak2),                                                                                                                                                                                                                                                              //  output,    width = 4,                  .txdatak2
		.txdatak3                       (txdatak3),                                                                                                                                                                                                                                                              //  output,    width = 4,                  .txdatak3
		.txdetectrx0                    (txdetectrx0),                                                                                                                                                                                                                                                           //  output,    width = 1,                  .txdetectrx0
		.txdetectrx1                    (txdetectrx1),                                                                                                                                                                                                                                                           //  output,    width = 1,                  .txdetectrx1
		.txdetectrx2                    (txdetectrx2),                                                                                                                                                                                                                                                           //  output,    width = 1,                  .txdetectrx2
		.txdetectrx3                    (txdetectrx3),                                                                                                                                                                                                                                                           //  output,    width = 1,                  .txdetectrx3
		.txelecidle0                    (txelecidle0),                                                                                                                                                                                                                                                           //  output,    width = 1,                  .txelecidle0
		.txelecidle1                    (txelecidle1),                                                                                                                                                                                                                                                           //  output,    width = 1,                  .txelecidle1
		.txelecidle2                    (txelecidle2),                                                                                                                                                                                                                                                           //  output,    width = 1,                  .txelecidle2
		.txelecidle3                    (txelecidle3),                                                                                                                                                                                                                                                           //  output,    width = 1,                  .txelecidle3
		.txdeemph0                      (txdeemph0),                                                                                                                                                                                                                                                             //  output,    width = 1,                  .txdeemph0
		.txdeemph1                      (txdeemph1),                                                                                                                                                                                                                                                             //  output,    width = 1,                  .txdeemph1
		.txdeemph2                      (txdeemph2),                                                                                                                                                                                                                                                             //  output,    width = 1,                  .txdeemph2
		.txdeemph3                      (txdeemph3),                                                                                                                                                                                                                                                             //  output,    width = 1,                  .txdeemph3
		.txmargin0                      (txmargin0),                                                                                                                                                                                                                                                             //  output,    width = 3,                  .txmargin0
		.txmargin1                      (txmargin1),                                                                                                                                                                                                                                                             //  output,    width = 3,                  .txmargin1
		.txmargin2                      (txmargin2),                                                                                                                                                                                                                                                             //  output,    width = 3,                  .txmargin2
		.txmargin3                      (txmargin3),                                                                                                                                                                                                                                                             //  output,    width = 3,                  .txmargin3
		.txswing0                       (txswing0),                                                                                                                                                                                                                                                              //  output,    width = 1,                  .txswing0
		.txswing1                       (txswing1),                                                                                                                                                                                                                                                              //  output,    width = 1,                  .txswing1
		.txswing2                       (txswing2),                                                                                                                                                                                                                                                              //  output,    width = 1,                  .txswing2
		.txswing3                       (txswing3),                                                                                                                                                                                                                                                              //  output,    width = 1,                  .txswing3
		.phystatus0                     (phystatus0),                                                                                                                                                                                                                                                            //   input,    width = 1,                  .phystatus0
		.phystatus1                     (phystatus1),                                                                                                                                                                                                                                                            //   input,    width = 1,                  .phystatus1
		.phystatus2                     (phystatus2),                                                                                                                                                                                                                                                            //   input,    width = 1,                  .phystatus2
		.phystatus3                     (phystatus3),                                                                                                                                                                                                                                                            //   input,    width = 1,                  .phystatus3
		.rxdata0                        (rxdata0),                                                                                                                                                                                                                                                               //   input,   width = 32,                  .rxdata0
		.rxdata1                        (rxdata1),                                                                                                                                                                                                                                                               //   input,   width = 32,                  .rxdata1
		.rxdata2                        (rxdata2),                                                                                                                                                                                                                                                               //   input,   width = 32,                  .rxdata2
		.rxdata3                        (rxdata3),                                                                                                                                                                                                                                                               //   input,   width = 32,                  .rxdata3
		.rxdatak0                       (rxdatak0),                                                                                                                                                                                                                                                              //   input,    width = 4,                  .rxdatak0
		.rxdatak1                       (rxdatak1),                                                                                                                                                                                                                                                              //   input,    width = 4,                  .rxdatak1
		.rxdatak2                       (rxdatak2),                                                                                                                                                                                                                                                              //   input,    width = 4,                  .rxdatak2
		.rxdatak3                       (rxdatak3),                                                                                                                                                                                                                                                              //   input,    width = 4,                  .rxdatak3
		.rxelecidle0                    (rxelecidle0),                                                                                                                                                                                                                                                           //   input,    width = 1,                  .rxelecidle0
		.rxelecidle1                    (rxelecidle1),                                                                                                                                                                                                                                                           //   input,    width = 1,                  .rxelecidle1
		.rxelecidle2                    (rxelecidle2),                                                                                                                                                                                                                                                           //   input,    width = 1,                  .rxelecidle2
		.rxelecidle3                    (rxelecidle3),                                                                                                                                                                                                                                                           //   input,    width = 1,                  .rxelecidle3
		.rxstatus0                      (rxstatus0),                                                                                                                                                                                                                                                             //   input,    width = 3,                  .rxstatus0
		.rxstatus1                      (rxstatus1),                                                                                                                                                                                                                                                             //   input,    width = 3,                  .rxstatus1
		.rxstatus2                      (rxstatus2),                                                                                                                                                                                                                                                             //   input,    width = 3,                  .rxstatus2
		.rxstatus3                      (rxstatus3),                                                                                                                                                                                                                                                             //   input,    width = 3,                  .rxstatus3
		.rxvalid0                       (rxvalid0),                                                                                                                                                                                                                                                              //   input,    width = 1,                  .rxvalid0
		.rxvalid1                       (rxvalid1),                                                                                                                                                                                                                                                              //   input,    width = 1,                  .rxvalid1
		.rxvalid2                       (rxvalid2),                                                                                                                                                                                                                                                              //   input,    width = 1,                  .rxvalid2
		.rxvalid3                       (rxvalid3),                                                                                                                                                                                                                                                              //   input,    width = 1,                  .rxvalid3
		.rxdataskip0                    (rxdataskip0),                                                                                                                                                                                                                                                           //   input,    width = 1,                  .rxdataskip0
		.rxdataskip1                    (rxdataskip1),                                                                                                                                                                                                                                                           //   input,    width = 1,                  .rxdataskip1
		.rxdataskip2                    (rxdataskip2),                                                                                                                                                                                                                                                           //   input,    width = 1,                  .rxdataskip2
		.rxdataskip3                    (rxdataskip3),                                                                                                                                                                                                                                                           //   input,    width = 1,                  .rxdataskip3
		.rxblkst0                       (rxblkst0),                                                                                                                                                                                                                                                              //   input,    width = 1,                  .rxblkst0
		.rxblkst1                       (rxblkst1),                                                                                                                                                                                                                                                              //   input,    width = 1,                  .rxblkst1
		.rxblkst2                       (rxblkst2),                                                                                                                                                                                                                                                              //   input,    width = 1,                  .rxblkst2
		.rxblkst3                       (rxblkst3),                                                                                                                                                                                                                                                              //   input,    width = 1,                  .rxblkst3
		.rxsynchd0                      (rxsynchd0),                                                                                                                                                                                                                                                             //   input,    width = 2,                  .rxsynchd0
		.rxsynchd1                      (rxsynchd1),                                                                                                                                                                                                                                                             //   input,    width = 2,                  .rxsynchd1
		.rxsynchd2                      (rxsynchd2),                                                                                                                                                                                                                                                             //   input,    width = 2,                  .rxsynchd2
		.rxsynchd3                      (rxsynchd3),                                                                                                                                                                                                                                                             //   input,    width = 2,                  .rxsynchd3
		.currentcoeff0                  (currentcoeff0),                                                                                                                                                                                                                                                         //  output,   width = 18,                  .currentcoeff0
		.currentcoeff1                  (currentcoeff1),                                                                                                                                                                                                                                                         //  output,   width = 18,                  .currentcoeff1
		.currentcoeff2                  (currentcoeff2),                                                                                                                                                                                                                                                         //  output,   width = 18,                  .currentcoeff2
		.currentcoeff3                  (currentcoeff3),                                                                                                                                                                                                                                                         //  output,   width = 18,                  .currentcoeff3
		.currentrxpreset0               (currentrxpreset0),                                                                                                                                                                                                                                                      //  output,    width = 3,                  .currentrxpreset0
		.currentrxpreset1               (currentrxpreset1),                                                                                                                                                                                                                                                      //  output,    width = 3,                  .currentrxpreset1
		.currentrxpreset2               (currentrxpreset2),                                                                                                                                                                                                                                                      //  output,    width = 3,                  .currentrxpreset2
		.currentrxpreset3               (currentrxpreset3),                                                                                                                                                                                                                                                      //  output,    width = 3,                  .currentrxpreset3
		.txsynchd0                      (txsynchd0),                                                                                                                                                                                                                                                             //  output,    width = 2,                  .txsynchd0
		.txsynchd1                      (txsynchd1),                                                                                                                                                                                                                                                             //  output,    width = 2,                  .txsynchd1
		.txsynchd2                      (txsynchd2),                                                                                                                                                                                                                                                             //  output,    width = 2,                  .txsynchd2
		.txsynchd3                      (txsynchd3),                                                                                                                                                                                                                                                             //  output,    width = 2,                  .txsynchd3
		.txblkst0                       (txblkst0),                                                                                                                                                                                                                                                              //  output,    width = 1,                  .txblkst0
		.txblkst1                       (txblkst1),                                                                                                                                                                                                                                                              //  output,    width = 1,                  .txblkst1
		.txblkst2                       (txblkst2),                                                                                                                                                                                                                                                              //  output,    width = 1,                  .txblkst2
		.txblkst3                       (txblkst3),                                                                                                                                                                                                                                                              //  output,    width = 1,                  .txblkst3
		.txdataskip0                    (txdataskip0),                                                                                                                                                                                                                                                           //  output,    width = 1,                  .txdataskip0
		.txdataskip1                    (txdataskip1),                                                                                                                                                                                                                                                           //  output,    width = 1,                  .txdataskip1
		.txdataskip2                    (txdataskip2),                                                                                                                                                                                                                                                           //  output,    width = 1,                  .txdataskip2
		.txdataskip3                    (txdataskip3),                                                                                                                                                                                                                                                           //  output,    width = 1,                  .txdataskip3
		.rate0                          (rate0),                                                                                                                                                                                                                                                                 //  output,    width = 2,                  .rate0
		.rate1                          (rate1),                                                                                                                                                                                                                                                                 //  output,    width = 2,                  .rate1
		.rate2                          (rate2),                                                                                                                                                                                                                                                                 //  output,    width = 2,                  .rate2
		.rate3                          (rate3),                                                                                                                                                                                                                                                                 //  output,    width = 2,                  .rate3
		.rx_in0                         (rx_in0),                                                                                                                                                                                                                                                                //   input,    width = 1,        hip_serial.rx_in0
		.rx_in1                         (rx_in1),                                                                                                                                                                                                                                                                //   input,    width = 1,                  .rx_in1
		.rx_in2                         (rx_in2),                                                                                                                                                                                                                                                                //   input,    width = 1,                  .rx_in2
		.rx_in3                         (rx_in3),                                                                                                                                                                                                                                                                //   input,    width = 1,                  .rx_in3
		.tx_out0                        (tx_out0),                                                                                                                                                                                                                                                               //  output,    width = 1,                  .tx_out0
		.tx_out1                        (tx_out1),                                                                                                                                                                                                                                                               //  output,    width = 1,                  .tx_out1
		.tx_out2                        (tx_out2),                                                                                                                                                                                                                                                               //  output,    width = 1,                  .tx_out2
		.tx_out3                        (tx_out3),                                                                                                                                                                                                                                                               //  output,    width = 1,                  .tx_out3
		.msi_intfc_o                    (msi_intfc_o),                                                                                                                                                                                                                                                           //  output,   width = 82,         msi_intfc.msi_intfc
		.msi_control_o                  (msi_control_o),                                                                                                                                                                                                                                                         //  output,   width = 16,       msi_control.msi_control
		.msix_intfc_o                   (msix_intfc_o),                                                                                                                                                                                                                                                          //  output,   width = 16,        msix_intfc.msix_intfc
		.intx_req_i                     (intx_req_i),                                                                                                                                                                                                                                                            //   input,    width = 1,        intx_intfc.intx_req
		.intx_ack_o                     (intx_ack_o),                                                                                                                                                                                                                                                            //  output,    width = 1,                  .intx_ack
		.txs_address_i                  (txs_address_i),                                                                                                                                                                                                                                                         //   input,   width = 64,               txs.address
		.txs_chipselect_i               (txs_chipselect_i),                                                                                                                                                                                                                                                      //   input,    width = 1,                  .chipselect
		.txs_byteenable_i               (txs_byteenable_i),                                                                                                                                                                                                                                                      //   input,   width = 16,                  .byteenable
		.txs_readdata_o                 (txs_readdata_o),                                                                                                                                                                                                                                                        //  output,  width = 128,                  .readdata
		.txs_writedata_i                (txs_writedata_i),                                                                                                                                                                                                                                                       //   input,  width = 128,                  .writedata
		.txs_read_i                     (txs_read_i),                                                                                                                                                                                                                                                            //   input,    width = 1,                  .read
		.txs_write_i                    (txs_write_i),                                                                                                                                                                                                                                                           //   input,    width = 1,                  .write
		.txs_burstcount_i               (txs_burstcount_i),                                                                                                                                                                                                                                                      //   input,    width = 6,                  .burstcount
		.txs_readdatavalid_o            (txs_readdatavalid_o),                                                                                                                                                                                                                                                   //  output,    width = 1,                  .readdatavalid
		.txs_waitrequest_o              (txs_waitrequest_o),                                                                                                                                                                                                                                                     //  output,    width = 1,                  .waitrequest
		.cra_chipselect_i               (cra_chipselect_i),                                                                                                                                                                                                                                                      //   input,    width = 1,               cra.chipselect
		.cra_address_i                  (cra_address_i),                                                                                                                                                                                                                                                         //   input,   width = 14,                  .address
		.cra_byteenable_i               (cra_byteenable_i),                                                                                                                                                                                                                                                      //   input,    width = 4,                  .byteenable
		.cra_read_i                     (cra_read_i),                                                                                                                                                                                                                                                            //   input,    width = 1,                  .read
		.cra_readdata_o                 (cra_readdata_o),                                                                                                                                                                                                                                                        //  output,   width = 32,                  .readdata
		.cra_write_i                    (cra_write_i),                                                                                                                                                                                                                                                           //   input,    width = 1,                  .write
		.cra_writedata_i                (cra_writedata_i),                                                                                                                                                                                                                                                       //   input,   width = 32,                  .writedata
		.cra_waitrequest_o              (cra_waitrequest_o),                                                                                                                                                                                                                                                     //  output,    width = 1,                  .waitrequest
		.cra_irq_o                      (cra_irq_o),                                                                                                                                                                                                                                                             //  output,    width = 1,           cra_irq.irq
		.rxm_bar0_address_o             (rxm_bar0_address_o),                                                                                                                                                                                                                                                    //  output,   width = 64,          rxm_bar0.address
		.rxm_bar0_byteenable_o          (rxm_bar0_byteenable_o),                                                                                                                                                                                                                                                 //  output,   width = 16,                  .byteenable
		.rxm_bar0_readdata_i            (rxm_bar0_readdata_i),                                                                                                                                                                                                                                                   //   input,  width = 128,                  .readdata
		.rxm_bar0_writedata_o           (rxm_bar0_writedata_o),                                                                                                                                                                                                                                                  //  output,  width = 128,                  .writedata
		.rxm_bar0_read_o                (rxm_bar0_read_o),                                                                                                                                                                                                                                                       //  output,    width = 1,                  .read
		.rxm_bar0_write_o               (rxm_bar0_write_o),                                                                                                                                                                                                                                                      //  output,    width = 1,                  .write
		.rxm_bar0_burstcount_o          (rxm_bar0_burstcount_o),                                                                                                                                                                                                                                                 //  output,    width = 6,                  .burstcount
		.rxm_bar0_readdatavalid_i       (rxm_bar0_readdatavalid_i),                                                                                                                                                                                                                                              //   input,    width = 1,                  .readdatavalid
		.rxm_bar0_waitrequest_i         (rxm_bar0_waitrequest_i),                                                                                                                                                                                                                                                //   input,    width = 1,                  .waitrequest
		.rxm_bar2_address_o             (rxm_bar2_address_o),                                                                                                                                                                                                                                                    //  output,   width = 64,          rxm_bar2.address
		.rxm_bar2_byteenable_o          (rxm_bar2_byteenable_o),                                                                                                                                                                                                                                                 //  output,   width = 16,                  .byteenable
		.rxm_bar2_readdata_i            (rxm_bar2_readdata_i),                                                                                                                                                                                                                                                   //   input,  width = 128,                  .readdata
		.rxm_bar2_writedata_o           (rxm_bar2_writedata_o),                                                                                                                                                                                                                                                  //  output,  width = 128,                  .writedata
		.rxm_bar2_read_o                (rxm_bar2_read_o),                                                                                                                                                                                                                                                       //  output,    width = 1,                  .read
		.rxm_bar2_write_o               (rxm_bar2_write_o),                                                                                                                                                                                                                                                      //  output,    width = 1,                  .write
		.rxm_bar2_burstcount_o          (rxm_bar2_burstcount_o),                                                                                                                                                                                                                                                 //  output,    width = 6,                  .burstcount
		.rxm_bar2_readdatavalid_i       (rxm_bar2_readdatavalid_i),                                                                                                                                                                                                                                              //   input,    width = 1,                  .readdatavalid
		.rxm_bar2_waitrequest_i         (rxm_bar2_waitrequest_i),                                                                                                                                                                                                                                                //   input,    width = 1,                  .waitrequest
		.rxm_irq_i                      (rxm_irq_i),                                                                                                                                                                                                                                                             //   input,   width = 16,           rxm_irq.irq
		.pld_clk                        (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.TxData_rdy_o                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.TxData_val_i                   (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.TxData_sop_i                   (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.TxData_eop_i                   (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.TxData_err_i                   (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.TxData_dat_i                   (256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), // (terminated),                                 
		.TxData_sty_i                   (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.TxData_mty_i                   (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.TxData_dsc_i                   (256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), // (terminated),                                 
		.TxStatus_val_o                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.TxStatus_dat_o                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.RxData_rdy_i                   (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.RxData_val_o                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.RxData_sop_o                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.RxData_eop_o                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.RxData_err_o                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.RxData_dat_o                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.RxData_sty_o                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.RxData_mty_o                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.RxData_dsc_o                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.pld_core_ready                 (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.pld_clk_inuse                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.serdes_pll_locked              (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.reset_status                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.testin_zero                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.sim_pipe_pclk_out              (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.devkit_status                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.devkit_ctrl                    (256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), // (terminated),                                 
		.rx_cred_ctl                    (16'b0000000000000000),                                                                                                                                                                                                                                                  // (terminated),                                 
		.rx_cred_status                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.derr_cor_ext_rcv               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.derr_cor_ext_rpl               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.derr_rpl                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.dlup                           (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.dlup_exit                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ev128ns                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ev1us                          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.hotrst_exit                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.int_status                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.l2_exit                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.lane_act                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ltssmstate                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rx_par_err                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.tx_par_err                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfg_par_err                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ko_cpl_spc_header              (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ko_cpl_spc_data                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxfc_cplbuf_ovf                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.currentspeed                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.tx_st_sop                      (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.tx_st_eop                      (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.tx_st_err                      (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.tx_st_valid                    (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.tx_st_ready                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.tx_st_data                     (128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                 // (terminated),                                 
		.tx_st_empty                    (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.tx_st_parity                   (16'b0000000000000000),                                                                                                                                                                                                                                                  // (terminated),                                 
		.rx_st_sop                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rx_st_eop                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rx_st_err                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rx_st_valid                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rx_st_ready                    (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rx_st_data                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rx_st_empty                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rx_st_parity                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.clr_st                         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rx_st_bar_range                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rx_st_pf_num                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rx_st_vf_num                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rx_st_vf_active                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.tx_st_pf_num                   (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.tx_st_vf_num                   (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.tx_st_vf_active                (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.extraBAR_lock                  (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.extraBAR_hit                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.devhide_pf                     (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.device_rciep                   (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rx_st_bar                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rx_st_bar_hit_tlp0             (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rx_st_bar_hit_fn_tlp0          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rx_st_bar_hit_tlp1             (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rx_st_bar_hit_fn_tlp1          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rx_st_mask                     (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.tx_cred_data_fc                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.tx_cred_fc_hip_cons            (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.tx_cred_fc_infinite            (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.tx_cred_hdr_fc                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.tx_cred_fc_sel                 (2'b00),                                                                                                                                                                                                                                                                 // (terminated),                                 
		.tx_cred_cons_select            (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.eidleinfersel4                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.eidleinfersel5                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.eidleinfersel6                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.eidleinfersel7                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.powerdown4                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.powerdown5                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.powerdown6                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.powerdown7                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxpolarity4                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxpolarity5                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxpolarity6                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxpolarity7                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txcompl4                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txcompl5                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txcompl6                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txcompl7                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdata4                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdata5                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdata6                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdata7                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdatak4                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdatak5                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdatak6                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdatak7                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdetectrx4                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdetectrx5                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdetectrx6                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdetectrx7                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txelecidle4                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txelecidle5                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txelecidle6                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txelecidle7                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdeemph4                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdeemph5                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdeemph6                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdeemph7                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txmargin4                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txmargin5                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txmargin6                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txmargin7                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txswing4                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txswing5                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txswing6                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txswing7                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.phystatus4                     (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.phystatus5                     (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.phystatus6                     (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.phystatus7                     (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxdata4                        (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.rxdata5                        (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.rxdata6                        (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.rxdata7                        (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.rxdatak4                       (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.rxdatak5                       (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.rxdatak6                       (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.rxdatak7                       (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.rxelecidle4                    (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxelecidle5                    (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxelecidle6                    (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxelecidle7                    (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxstatus4                      (3'b000),                                                                                                                                                                                                                                                                // (terminated),                                 
		.rxstatus5                      (3'b000),                                                                                                                                                                                                                                                                // (terminated),                                 
		.rxstatus6                      (3'b000),                                                                                                                                                                                                                                                                // (terminated),                                 
		.rxstatus7                      (3'b000),                                                                                                                                                                                                                                                                // (terminated),                                 
		.rxvalid4                       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxvalid5                       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxvalid6                       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxvalid7                       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxdataskip4                    (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxdataskip5                    (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxdataskip6                    (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxdataskip7                    (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxblkst4                       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxblkst5                       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxblkst6                       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxblkst7                       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxsynchd4                      (2'b00),                                                                                                                                                                                                                                                                 // (terminated),                                 
		.rxsynchd5                      (2'b00),                                                                                                                                                                                                                                                                 // (terminated),                                 
		.rxsynchd6                      (2'b00),                                                                                                                                                                                                                                                                 // (terminated),                                 
		.rxsynchd7                      (2'b00),                                                                                                                                                                                                                                                                 // (terminated),                                 
		.currentcoeff4                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.currentcoeff5                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.currentcoeff6                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.currentcoeff7                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.currentrxpreset4               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.currentrxpreset5               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.currentrxpreset6               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.currentrxpreset7               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txsynchd4                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txsynchd5                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txsynchd6                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txsynchd7                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txblkst4                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txblkst5                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txblkst6                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txblkst7                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdataskip4                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdataskip5                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdataskip6                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.txdataskip7                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rate4                          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rate5                          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rate6                          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rate7                          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rx_in4                         (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rx_in5                         (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rx_in6                         (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rx_in7                         (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.tx_out4                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.tx_out5                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.tx_out6                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.tx_out7                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.app_int_sts                    (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.app_int_pf_sts                 (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.app_int_sts_a                  (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.app_int_sts_b                  (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.app_int_sts_c                  (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.app_int_sts_d                  (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.app_int_sts_fn                 (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.app_int_pend_status            (2'b00),                                                                                                                                                                                                                                                                 // (terminated),                                 
		.app_int_ack                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.app_intx_disable               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.app_msi_num                    (5'b00000),                                                                                                                                                                                                                                                              // (terminated),                                 
		.app_msi_req                    (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.app_msi_tc                     (3'b000),                                                                                                                                                                                                                                                                // (terminated),                                 
		.app_msi_ack                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.app_msi_status                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.app_msi_req_fn                 (8'b00000000),                                                                                                                                                                                                                                                           // (terminated),                                 
		.app_msi_pending_bit_write_en   (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.app_msi_pending_bit_write_data (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.app_msix_req                   (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.app_msix_tc                    (3'b000),                                                                                                                                                                                                                                                                // (terminated),                                 
		.app_msix_ack                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.app_msix_err                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.app_msix_addr                  (64'b0000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                                                                                  // (terminated),                                 
		.app_msix_data                  (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.app_msix_pf_num                (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.app_msix_vf_num                (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.app_msix_vf_active             (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.app_msi_addr_pf                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.app_msi_data_pf                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.app_msi_mask_pf                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.app_msi_pending_pf             (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.app_msi_enable_pf              (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.app_msi_multi_msg_enable_pf    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.app_msix_en_pf                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.app_msix_fn_mask_pf            (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.app_msix_en_vf                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.app_msix_fn_mask_vf            (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.serr_out                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.aer_msi_num                    (5'b00000),                                                                                                                                                                                                                                                              // (terminated),                                 
		.pex_msi_num                    (5'b00000),                                                                                                                                                                                                                                                              // (terminated),                                 
		.lmi_addr                       (12'b000000000000),                                                                                                                                                                                                                                                      // (terminated),                                 
		.lmi_din                        (8'b00000000),                                                                                                                                                                                                                                                           // (terminated),                                 
		.lmi_rden                       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.lmi_wren                       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.lmi_func                       (9'b000000000),                                                                                                                                                                                                                                                          // (terminated),                                 
		.lmi_ack                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.lmi_dout                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.lmi_pf_num_app                 (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.lmi_vf_num_app                 (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.lmi_vf_active_app              (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.pm_auxpwr                      (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.pm_data                        (10'b0000000000),                                                                                                                                                                                                                                                        // (terminated),                                 
		.pme_to_cr                      (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.pm_event                       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.pme_to_sr                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_link2csr                 (16'b0000000000000000),                                                                                                                                                                                                                                                  // (terminated),                                 
		.cfgbp_comclk_reg               (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.cfgbp_extsy_reg                (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.cfgbp_max_pload                (3'b000),                                                                                                                                                                                                                                                                // (terminated),                                 
		.cfgbp_tx_ecrcgen               (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.cfgbp_rx_ecrchk                (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.cfgbp_secbus                   (8'b00000000),                                                                                                                                                                                                                                                           // (terminated),                                 
		.cfgbp_linkcsr_bit0             (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.cfgbp_tx_req_pm                (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.cfgbp_tx_typ_pm                (3'b000),                                                                                                                                                                                                                                                                // (terminated),                                 
		.cfgbp_req_phypm                (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.cfgbp_req_phycfg               (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.cfgbp_vc0_tcmap_pld            (7'b0000000),                                                                                                                                                                                                                                                            // (terminated),                                 
		.cfgbp_inh_dllp                 (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.cfgbp_inh_tx_tlp               (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.cfgbp_req_wake                 (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.cfgbp_link3_ctl                (2'b00),                                                                                                                                                                                                                                                                 // (terminated),                                 
		.cfgbp_lane_err                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_link_equlz_req           (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_equiz_complete           (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_phase_3_successful       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_phase_2_successful       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_phase_1_successful       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_current_deemph           (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_current_speed            (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_link_up                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_link_train               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_10state                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_10sstate                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_rx_val_pm                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_rx_typ_pm                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_tx_ack_pm                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_ack_phypm                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_vc_status                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_rxfc_max                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_txfc_max                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_txbuf_emp                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_cfgbuf_emp               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_rpbuf_emp                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_dll_req                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_link_auto_bdw_status     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_link_bdw_mng_status      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_rst_tx_margin_field      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_rst_enter_comp_bit       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_rx_st_ecrcerr            (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_err_uncorr_internal      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_rx_corr_internal         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_err_tlrcvovf             (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_txfc_err                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_err_tlmalf               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_err_surpdwn_dll          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_err_dllrev               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_err_dll_repnum           (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_err_dllreptim            (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_err_dllp_baddllp         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_err_dll_badtlp           (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_err_phy_tng              (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_err_phy_rcv              (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_root_err_reg_sts         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_corr_err_reg_sts         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cfgbp_unc_err_reg_sts          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cseb_rddata                    (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.cseb_rdresponse                (5'b00000),                                                                                                                                                                                                                                                              // (terminated),                                 
		.cseb_waitrequest               (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.cseb_wrresponse                (5'b00000),                                                                                                                                                                                                                                                              // (terminated),                                 
		.cseb_wrresp_valid              (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.cseb_addr                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cseb_be                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cseb_rden                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cseb_wrdata                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cseb_wren                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cseb_is_shadow                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cseb_wrresp_req                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cseb_rddata_parity             (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.cseb_addr_parity               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cseb_wrdata_parity             (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.hip_reconfig_clk               (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.hip_reconfig_rst_n             (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.hip_reconfig_address           (10'b0000000000),                                                                                                                                                                                                                                                        // (terminated),                                 
		.hip_reconfig_read              (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.hip_reconfig_readdata          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.hip_reconfig_write             (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.hip_reconfig_writedata         (16'b0000000000000000),                                                                                                                                                                                                                                                  // (terminated),                                 
		.hip_reconfig_byte_en           (2'b00),                                                                                                                                                                                                                                                                 // (terminated),                                 
		.ser_shift_load                 (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.interface_sel                  (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.xcvr_reconfig_clk              (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.xcvr_reconfig_reset            (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.xcvr_reconfig_address          (12'b000000000000),                                                                                                                                                                                                                                                      // (terminated),                                 
		.xcvr_reconfig_read             (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.xcvr_reconfig_readdata         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.xcvr_reconfig_write            (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.xcvr_reconfig_writedata        (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.xcvr_reconfig_waitrequest      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.reconfig_pll0_clk              (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.reconfig_pll0_reset            (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.reconfig_pll0_address          (10'b0000000000),                                                                                                                                                                                                                                                        // (terminated),                                 
		.reconfig_pll0_read             (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.reconfig_pll0_readdata         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.reconfig_pll0_write            (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.reconfig_pll0_writedata        (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.reconfig_pll0_waitrequest      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.reconfig_pll1_clk              (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.reconfig_pll1_reset            (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.reconfig_pll1_address          (10'b0000000000),                                                                                                                                                                                                                                                        // (terminated),                                 
		.reconfig_pll1_read             (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.reconfig_pll1_readdata         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.reconfig_pll1_write            (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.reconfig_pll1_writedata        (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.reconfig_pll1_waitrequest      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.pipe_hclk_in                   (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.pll_pcie_clk                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.hpg_ctrler                     (5'b00000),                                                                                                                                                                                                                                                              // (terminated),                                 
		.tl_cfg_add                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.tl_cfg_ctl                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.tl_cfg_sts                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.cpl_err                        (7'b0000000),                                                                                                                                                                                                                                                            // (terminated),                                 
		.cpl_pending                    (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.cpl_err_fn                     (8'b00000000),                                                                                                                                                                                                                                                           // (terminated),                                 
		.cpl_pending_pf                 (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.cpl_pending_vf                 (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.log_hdr                        (128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                 // (terminated),                                 
		.cpl_err_pf_num                 (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.cpl_err_vf_num                 (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.cpl_err_vf_active              (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.vf_compl_status_update         (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.vf_compl_status                (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.vf_compl_status_pf_num         (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.vf_compl_status_vf_num         (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.vf_compl_status_update_ack     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.flr_active_pf                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.flr_active_vf                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.flr_completed_pf               (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.flr_completed_vf               (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.flr_rcvd_vf                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.flr_rcvd_pf_num                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.flr_rcvd_vf_num                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.flr_completed_pf_num           (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.flr_completed_vf_num           (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.bus_num_f0                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.bus_num_f1                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.device_num_f0                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.device_num_f1                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.mem_space_en_pf                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.bus_master_en_pf               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.mem_space_en_vf                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.exprom_en_pf                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.bus_master_en_vf               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.pf0_num_vfs                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.pf1_num_vfs                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.pf_max_payload_size            (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.pf_rd_req_size                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.bus_num_f2                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.bus_num_f3                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.device_num_f2                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.device_num_f3                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.bus_num_f4                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.bus_num_f5                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.device_num_f4                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.device_num_f5                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.bus_num_f6                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.bus_num_f7                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.device_num_f6                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.device_num_f7                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.pf2_num_vfs                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.pf3_num_vfs                    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.extended_tag_en_pf             (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.compl_timeout_disable_pf       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.atomic_op_requester_en_pf      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.tph_st_mode_pf                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.tph_requester_en_pf            (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ats_stu_pf                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ats_en_pf                      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ctl_shdw_update                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ctl_shdw_pf_num                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ctl_shdw_vf_num                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ctl_shdw_vf_active             (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ctl_shdw_cfg                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ctl_shdw_req_all               (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.f0_virtio_pcicfg_bar_o         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f0_virtio_pcicfg_length_o      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f0_virtio_pcicfg_baroffset_o   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f0_virtio_pcicfg_cfgdata_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f0_virtio_pcicfg_cfgwr_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f0_virtio_pcicfg_cfgrd_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f0_virtio_pcicfg_rdack_i       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.f0_virtio_pcicfg_rdbe_i        (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.f0_virtio_pcicfg_data_i        (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.f1_virtio_pcicfg_bar_o         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f1_virtio_pcicfg_length_o      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f1_virtio_pcicfg_baroffset_o   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f1_virtio_pcicfg_cfgdata_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f1_virtio_pcicfg_cfgwr_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f1_virtio_pcicfg_cfgrd_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f1_virtio_pcicfg_rdack_i       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.f1_virtio_pcicfg_rdbe_i        (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.f1_virtio_pcicfg_data_i        (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.f2_virtio_pcicfg_bar_o         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f2_virtio_pcicfg_length_o      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f2_virtio_pcicfg_baroffset_o   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f2_virtio_pcicfg_cfgdata_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f2_virtio_pcicfg_cfgwr_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f2_virtio_pcicfg_cfgrd_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f2_virtio_pcicfg_rdack_i       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.f2_virtio_pcicfg_rdbe_i        (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.f2_virtio_pcicfg_data_i        (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.f3_virtio_pcicfg_bar_o         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f3_virtio_pcicfg_length_o      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f3_virtio_pcicfg_baroffset_o   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f3_virtio_pcicfg_cfgdata_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f3_virtio_pcicfg_cfgwr_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f3_virtio_pcicfg_cfgrd_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f3_virtio_pcicfg_rdack_i       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.f3_virtio_pcicfg_rdbe_i        (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.f3_virtio_pcicfg_data_i        (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.f4_virtio_pcicfg_bar_o         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f4_virtio_pcicfg_length_o      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f4_virtio_pcicfg_baroffset_o   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f4_virtio_pcicfg_cfgdata_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f4_virtio_pcicfg_cfgwr_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f4_virtio_pcicfg_cfgrd_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f4_virtio_pcicfg_rdack_i       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.f4_virtio_pcicfg_rdbe_i        (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.f4_virtio_pcicfg_data_i        (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.f5_virtio_pcicfg_bar_o         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f5_virtio_pcicfg_length_o      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f5_virtio_pcicfg_baroffset_o   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f5_virtio_pcicfg_cfgdata_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f5_virtio_pcicfg_cfgwr_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f5_virtio_pcicfg_cfgrd_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f5_virtio_pcicfg_rdack_i       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.f5_virtio_pcicfg_rdbe_i        (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.f5_virtio_pcicfg_data_i        (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.f6_virtio_pcicfg_bar_o         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f6_virtio_pcicfg_length_o      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f6_virtio_pcicfg_baroffset_o   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f6_virtio_pcicfg_cfgdata_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f6_virtio_pcicfg_cfgwr_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f6_virtio_pcicfg_cfgrd_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f6_virtio_pcicfg_rdack_i       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.f6_virtio_pcicfg_rdbe_i        (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.f6_virtio_pcicfg_data_i        (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.f7_virtio_pcicfg_bar_o         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f7_virtio_pcicfg_length_o      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f7_virtio_pcicfg_baroffset_o   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f7_virtio_pcicfg_cfgdata_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f7_virtio_pcicfg_cfgwr_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f7_virtio_pcicfg_cfgrd_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f7_virtio_pcicfg_rdack_i       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.f7_virtio_pcicfg_rdbe_i        (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.f7_virtio_pcicfg_data_i        (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.f0vf_virtio_pcicfg_bar_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f0vf_virtio_pcicfg_length_o    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f0vf_virtio_pcicfg_baroffset_o (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f0vf_virtio_pcicfg_cfgdata_o   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f0vf_virtio_pcicfg_cfgwr_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f0vf_virtio_pcicfg_cfgrd_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f0vf_virtio_pcicfg_vfnum_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f0vf_virtio_pcicfg_rdack_i     (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.f0vf_virtio_pcicfg_rdbe_i      (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.f0vf_virtio_pcicfg_data_i      (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.f0vf_virtio_pcicfg_appvfnum_i  (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.f1vf_virtio_pcicfg_bar_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f1vf_virtio_pcicfg_length_o    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f1vf_virtio_pcicfg_baroffset_o (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f1vf_virtio_pcicfg_cfgdata_o   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f1vf_virtio_pcicfg_cfgwr_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f1vf_virtio_pcicfg_cfgrd_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f1vf_virtio_pcicfg_vfnum_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f1vf_virtio_pcicfg_rdack_i     (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.f1vf_virtio_pcicfg_rdbe_i      (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.f1vf_virtio_pcicfg_data_i      (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.f1vf_virtio_pcicfg_appvfnum_i  (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.f2vf_virtio_pcicfg_bar_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f2vf_virtio_pcicfg_length_o    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f2vf_virtio_pcicfg_baroffset_o (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f2vf_virtio_pcicfg_cfgdata_o   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f2vf_virtio_pcicfg_cfgwr_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f2vf_virtio_pcicfg_cfgrd_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f2vf_virtio_pcicfg_vfnum_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f2vf_virtio_pcicfg_rdack_i     (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.f2vf_virtio_pcicfg_rdbe_i      (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.f2vf_virtio_pcicfg_data_i      (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.f2vf_virtio_pcicfg_appvfnum_i  (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.f3vf_virtio_pcicfg_bar_o       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f3vf_virtio_pcicfg_length_o    (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f3vf_virtio_pcicfg_baroffset_o (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f3vf_virtio_pcicfg_cfgdata_o   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f3vf_virtio_pcicfg_cfgwr_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f3vf_virtio_pcicfg_cfgrd_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f3vf_virtio_pcicfg_vfnum_o     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.f3vf_virtio_pcicfg_rdack_i     (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.f3vf_virtio_pcicfg_rdbe_i      (4'b0000),                                                                                                                                                                                                                                                               // (terminated),                                 
		.f3vf_virtio_pcicfg_data_i      (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.f3vf_virtio_pcicfg_appvfnum_i  (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.avmm_thinmaster_reset          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.avmm_thinmaster_address        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.avmm_thinmaster_byteenable     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.avmm_thinmaster_readdata       (16'b0000000000000000),                                                                                                                                                                                                                                                  // (terminated),                                 
		.avmm_thinmaster_writedata      (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.avmm_thinmaster_read           (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.avmm_thinmaster_write          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.avmm_thinmaster_readdatavalid  (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.avmm_thinmaster_waitrequest    (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxm_bar1_address_o             (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar1_byteenable_o          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar1_readdata_i            (128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                 // (terminated),                                 
		.rxm_bar1_writedata_o           (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar1_read_o                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar1_write_o               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar1_burstcount_o          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar1_readdatavalid_i       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxm_bar1_waitrequest_i         (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxm_bar3_address_o             (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar3_byteenable_o          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar3_readdata_i            (128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                 // (terminated),                                 
		.rxm_bar3_writedata_o           (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar3_read_o                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar3_write_o               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar3_burstcount_o          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar3_readdatavalid_i       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxm_bar3_waitrequest_i         (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxm_bar4_address_o             (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar4_byteenable_o          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar4_readdata_i            (128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                 // (terminated),                                 
		.rxm_bar4_writedata_o           (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar4_read_o                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar4_write_o               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar4_burstcount_o          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar4_readdatavalid_i       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxm_bar4_waitrequest_i         (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxm_bar5_address_o             (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar5_byteenable_o          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar5_readdata_i            (128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                 // (terminated),                                 
		.rxm_bar5_writedata_o           (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar5_read_o                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar5_write_o               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar5_burstcount_o          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rxm_bar5_readdatavalid_i       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rxm_bar5_waitrequest_i         (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.hprxm_address_o                (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.hprxm_byteenable_o             (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.hprxm_readdata_i               (128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                 // (terminated),                                 
		.hprxm_writedata_o              (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.hprxm_read_o                   (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.hprxm_write_o                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.hprxm_burstcount_o             (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.hprxm_readdatavalid_i          (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.hprxm_waitrequest_i            (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rd_ast_rx_valid_i              (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rd_ast_rx_data_i               (160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                 // (terminated),                                 
		.rd_ast_rx_ready_o              (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rd_ast_tx_valid_o              (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rd_ast_tx_data_o               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.wr_ast_rx_valid_i              (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.wr_ast_rx_data_i               (160'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                 // (terminated),                                 
		.wr_ast_rx_ready_o              (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.wr_ast_tx_valid_o              (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.wr_ast_tx_data_o               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rd_dma_address_o               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rd_dma_write_o                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rd_dma_write_data_o            (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rd_dma_wait_request_i          (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rd_dma_burst_count_o           (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rd_dma_byte_enable_o           (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.wr_dma_address_o               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.wr_dma_read_o                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.wr_dma_read_data_i             (128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000),                                                                                                                                 // (terminated),                                 
		.wr_dma_wait_request_i          (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.wr_dma_burst_count_o           (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.wr_dma_read_data_valid_i       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rd_dts_chip_select_i           (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rd_dts_write_i                 (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rd_dts_burst_count_i           (5'b00000),                                                                                                                                                                                                                                                              // (terminated),                                 
		.rd_dts_address_i               (8'b00000000),                                                                                                                                                                                                                                                           // (terminated),                                 
		.rd_dts_write_data_i            (256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), // (terminated),                                 
		.rd_dts_wait_request_o          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.wr_dts_chip_select_i           (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.wr_dts_write_i                 (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.wr_dts_burst_count_i           (5'b00000),                                                                                                                                                                                                                                                              // (terminated),                                 
		.wr_dts_address_i               (8'b00000000),                                                                                                                                                                                                                                                           // (terminated),                                 
		.wr_dts_write_data_i            (256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), // (terminated),                                 
		.wr_dts_wait_request_o          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rd_dcm_address_o               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rd_dcm_write_o                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rd_dcm_writedata_o             (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rd_dcm_read_o                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rd_dcm_byte_enable_o           (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.rd_dcm_wait_request_i          (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.rd_dcm_read_data_i             (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.rd_dcm_read_data_valid_i       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.wr_dcm_address_o               (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.wr_dcm_write_o                 (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.wr_dcm_writedata_o             (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.wr_dcm_read_o                  (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.wr_dcm_byte_enable_o           (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.wr_dcm_wait_request_i          (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.wr_dcm_read_data_i             (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.wr_dcm_read_data_valid_i       (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.skp_os                         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.debug                          (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ceb_ack                        (1'b0),                                                                                                                                                                                                                                                                  // (terminated),                                 
		.ceb_din                        (32'b00000000000000000000000000000000),                                                                                                                                                                                                                                  // (terminated),                                 
		.ceb_addr                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ceb_req                        (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ceb_dout                       (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ceb_wr                         (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ceb_pf_num                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ceb_vf_num                     (),                                                                                                                                                                                                                                                                      // (terminated),                                 
		.ceb_vf_active                  ()                                                                                                                                                                                                                                                                       // (terminated),                                 
	);

endmodule
