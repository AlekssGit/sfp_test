// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ZZp666AHvJvwNhYs981I9poqfYxHIu3/BRVxJkOsLj4B+lJUSHIJgRDVXfvnnTmjmBGw5RoHyVZ6
7Xe83AYwpfYyl5JLKqANblvfYw0VlEB76PJpj8MPksFXRNGYYm2NdERYPgilx2Ya3lUPoJIdKW2u
EDHXkKfcbMOjRYFW1VVYPp7LcIF7bT82W05uSUpmIvdmMqvyeeBoKisdhWyRs3sUFgiK935J4IuW
wWuW1HJEBM56Jv6R/9E1k0FDUUv03Az40H9lCgsS23vgt2/tXT77PuZB/9etV/bKaWbR3fbDU3+w
jQQRQzjAj9Nc8hkpLlBgvdBqEWdVxpfHjy3x2g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5600)
TzyQWmHe00eizAdFvuSyTgmOEyPD7QrBWU4AzXKrJXOdq6YfdzrLZ0D77OJLoxIgDlbegQSZtrbH
ks8H0vinXkc2oJ3O3cX1/PwAQ0viBSyTxvpQ3TT+ciDt5V10eqmPbb8eKrBIa/RGsayydZUbBcVh
xvSH1lfp1htrHcApB4avPP5keoxMoqnWyhlTvCxLW3iNEySflN4LY9oNmcqnRynFscf9kIwviqdu
ojXCvBTMLwe58hRmZE07eqp+Vb03rrlRk/flSJnNGG2iNf84vnuHFea8SOh8OiWkNunPt5g0AH7Z
VAn732TfMV9FLGaWsCamZ/pswJSteEEU3vns+IRHRdEBDj/kFb2JWU4PqABHlXjRdNMyDmQTg/Dd
2xrz9uGvBlf2eqXTurC/45weEqARk4LPDSTjpvf/g7b8SQX8eNO018aoQtH341vueBH5e3U6eDzx
5S1QCK46mQ0ReDUkR+PaADB+/lMDM9FZBFQHnNy9KzFlpga1zcJn6g52fcsOPHkVEQe7qdWLQs5S
iCb8YFarEfQUWmbdcwoDaBk2rb/WG8CWvIpry/OsFxRyZTWM/ps9xBoruzPXrsIu37JkDuE5XnOZ
uX+Z+zmG6oV6wGu7V2G28qD98fzsbiDPJGJW4nQrB8/B8YX4XSKRCxtcmsUkkRqrEzojBimKNJ2s
dQFGH6K3cZV60jSMxyiGVolAGMtYnTpvawfqlOk7RD6hW1Ua9GU0E/cmCrfXkyU9EhO33LnX7qNb
tdje+rO1FQrBEEjRInUqFjBJNmoHp4K7g1j1iA+OwR0bP4R1w+XeSIpD9Vt6kfc2p9EJDZQBvDFJ
6+njmwP1so4z+/Tn0Miafdvd/3ahIe55aUDP2oZb1Wkx1dnw2mzebE1c2wAS/si3UnxKNyGibrvU
Uadw+hS6ysm6AVGQIvj6A0EvmPJTth1XO8IBKk9//dHi100FQV6x9y1XAMzPkLkllPX6ylqpFkVU
doJg0SYICnEtR6MMNRXcOaefxTm38Xc6Eq3Qp2h+osKDXURJ9k5eeon7I0i+8UwbiQfntFIgWqyW
FNLYkG2kkzfnT6wzGd9zLvrrKkVdl2xdktLWfQ+d4BGuIl7yw4wbHfsyRUdG8KF8tTBRuBU/e+ca
4MPKYUn18rFeM440ZVDFphw9xEgAkylamKsYeCZ+OVtenRU0UI/olN+bTUpE5gHuXZvKOJD/1lCw
Y+LxwAJHU8NskJRxPLqzUGF2Ga4kbkVMhhl0tntvCQFc8KwsxLvEaYM9kg3pF6FKpjBHDl16dx3/
8QtZl37y2Llt9DCS+hgVkyRVtA5TtmbvPJjaU1h9XjXinm+735oG213TZ/3E3fYmoTFb0itU+Dqi
bo5OXr+yaBk1KW6IpJAAwz9KgOMCEb6kmca/0fgGD7Go+Z+s5G2dDiCuNvb93KFWswV3dZ5y/iZu
JeyKKueaJ0Wcd6MEbSvdCczyNb3pXbXtUPGyXwCutOwMMm1+bmCbRfJAoqOkW/3q37IW4713M/YQ
i82vGEAS5KvMWuPFyOV73sD0Sgd66Ee6LQqXTxvB/EcqCs2d1iiVgf3OY6FJMt+BW0PM3C6OXL3V
DTg/FvjQBBgCxFKxcQo3VJWF3097RxtZ48gjbHEcNXFfL2RA4ohGGjSFDm8ZBdaZVSmrlgCJde9x
W/3xtYuKrm0YEee3SB3/PJAHmdbdQIlOtn8C6OJRuyLqWs/ztE0nUsYC/+qSCTOOj04d9yxUz8Qe
pqSUNfVoVrl+1+mAO899HKagEjzaBrBzyDjYOXG/9ZZ/l+oTU35/tZrCQjxUAW9Cus4WswF8kqBw
UrehKsxHHs3Wz42i740JAnYUuKz4OZiF+pVnL3xTj26tAE6IrWmEmGG+ma9lzLwfX4CDd4OsQyLj
vnHS6XAap7XARZrWlkK0q3dSBjsu+VUW6d72YkUW9y68XA37MT98wlWA8n1LDkscWCsRMlaS7IOV
RVSZSU6x1IvdZTRW86rYso+64oKyyT15PjVZbxjjqop5kGtOOIV1tLGZg8twh9oiMgkTxd9AIToO
/0rPWAjVneXdK06+KoritaUJ7c97NECcsQcDJljFR//9cMrlNXkgBixg/hJMgyxCZvG/picbrhgG
rbPafH1szTeO7KjUpnp417A+xgWNZ1i2jWX+5J2tdRINuLCqFwJs1VhS7u7g67kEPnQtk01JFxXD
MicKEwjeyN0K+VqL4GNisPXOMDbB5JeJjsg1bpzYEq2jpyR5l9ue0ibgMfuXxuNbT6XlD1JUlBlE
k7kXiuH9KuUg95kD3GqfbrOZeFTp2HB3boQLlcKnu8EgeGzRVcQPHnlr7AZpQej+G2B5yJn72GDz
XOLmpT+jR9/0MwQqNwZPFMcTJes5jhqf41moS7hkGBxQ9Fo3Bpz//DeHSX6kuJKGq59oYVSMoaOK
fHpM1IjslFMq6AoZ++TDLdntPtxn6WsDb9abWS92M+yh57U1y2L1No5ErdSe1iyAJ7NsPXnnH1SA
GyuKk+imcGC2LVA9Ae6z8fakkNJk50YUWuh6RpraXrTdn4wD14LRP0EVFYrtUdgQp1XwTvjntDTm
yeaieYudWu839jZ1lVzBYag8Hd8EOyr7K8PGdq0l0Bt/5uBZce5qGBWMURMTFAUpx5FGS2FUDy76
IT/w3ah+5GHikpsrVsBlKzqdTnBO/CLUsKz89mfDdoE30vOX7yoXkPLtlVJm+8FwUKzHu0J1pO9k
oMWkCkeiAE4GBdgslkISOeu7sBH5rqE+ns5B3sVq4Po/Gfkjkna33C4TZMRtv3jpYJQr159z77Hf
cOyfEqkEDfEkc1R1LDAOGgS2pgzkHdmpbRaDXSCb/fZ5sqxvQdxOg47RcFIMXHpyfWhow39BVfYN
fEfP1W1SLm6uaIMjnqjZxh/1j8dm8O0h6ZELhoONycV+f8dY7qipOorEFJ/f9ZwYSf951vmpIPHm
uZU/Si7a4Go8h2aaxYsESjp5ic6LAUqBv3p+tNnRr3P6oxlXyF0RoCvnOsKy61Eb+hOxE9lZGp39
DrhckoBmrCU48/HTK63QXrJ8iTuU4/akHQgY5ofRVfVKCthmTVOuqhMINt+MLbzyCGO5+qw78eOP
5lP3rQdYVAveMCWr4G3Uk6zGfBpwqshLc65f5abweQoC7Bfw3l0m+u5TjtK51jAuRQd+qGr0ckUW
w3zIO4AU/iPeo5wwWtkBAaVqt3ryFIfwgAayQn2G7nZE1LeJu57kHGfmOcsuQxCauTa72f2SMet+
XIxkY0YpundFVnrZIDPFH6jVke2LmCtNQ2BdvfVNJkblXyL7yR7zokbXcAAfBd+fjKiSdSu4zbF/
CGWf37zs7ird5TwVjui7yMpR+YMx5cbbHM55/zBu5S7AG0IBr5bo31WkHCN5/z6W5mT6yesHnUn8
Q2NpxXYOg/gRRJAcfOTPHu1xNpyWOmUwnOWT+YYTPqC8ZZ1x030FFUd9qRDuVrgtBGT/x9i0gTbh
QLGVRV0ouoC0HLyYVDZRBXMahHfiDG7SLZ6baLySCH8Es9PONp4ajZj/qcxxG0V18Roo4f+ixO+g
YxQkLuYyl7phiyiWfRSnP15+W2PvvWay7jyJDpOe+pFdsi8eZ/AsJLorrVtxZKO84u2Rb4PpUrY4
43UfQxHOvUlzXZnABauy9H9IjoYQcBVSevcMhkr6J7IMMHyd20uOgFaCBCGjaCGyY0wDKnzMbGWb
NxrGqJg/e3Y6NxG5eitDdJGHFlpAwaj+iMeb+3g5kGexjqfngHay10zvUs4HV4nu4KdNEcqPLn2k
ekcUHut5zZ1/pAHqv0Q+R/OflW6T4i8vBAho6vVd/rVMQnBUa9VlfTVdni6SbyXJp8HnDL9YrRft
Oy6ATvuErabjC4FU68Yk98U0vjVPjf3r58V394nSBRpQEIYdEm572zs5WRt84+Vfegs/yqEs2rmU
wPApuCr9E/16ZRYv4jkU3/ICBvDvEtvjq9qQ7eoRshfpwo7sAb8ZZAQ1JUUNX8OxpgoONS+TenvQ
3Y8aW9AZk4zEppWFOiEKl1dseG8d4d8in0jKYW4oU5j2/iRtBr6LjfRvICP678Z5YpPjkstp0CmQ
C15qpBALnOTGLQofY+177ul7MMkLH9NIGWOFAh/fL2kr8XhEYaoeVed+u1azZxXogBRo0MsvHCza
BNjlgRqOq805xJAWHKjLkWMs6ZNxi9deZU2O0YE4YXroBMxcaGQQXiuSZmKFXGnrHIST+Hg5yCai
Izv6RoZD+7vD36NNkWJzK26Eoo6MK7ZkbUyLLBdbKKiZKkpJ30/csA6Gmz3YKlkAt8JMWc/YR0t7
UZ4yQe+pj5gknykn/VBbU45gQibIE3G1PLUdtlNVOUgLUAGyy5tR8tbOgWC7FxSbjwU0H3q/s0VU
Za+9O7StCxSQAzR/jt1g3QiJHq3kRZjbgZrEJ4lL7RJr9UxgkgSrNFG0VqLqZ7bbSn4xYxwn2XZx
v4Bl4azsivEggiV0Z+4T3WMp7CrTdnSf60vC7k8LTvOpTuy11oTSxFPmKGAVvPCRVAkfQrmK2zt7
qe9pd5AePE0kN8N+2nNxKj1HaY+vIqBskbjvl4bDXN//HYOgVXx+jf14Fa7lpTG9+i/I7fzz9Ybj
Azg8sZMkSqrrj+P8r9kNrVfQkqIYj4EMG5pLEXKbEF2CUCWR6Ysfa9ctXo4VrcajcgfuCarQF6Nf
znuskpVWO2cCPGWqOljRSNhm75JPYlNFQma4NfR3G4LBDXpldQQvmEz+DUVcduWTXAIE61m6ur1Y
vCGr8rBzcu4il1YHUiaQRSlGO061UrCU9OO6/J25wWgkvyc/XC8YiWwTRy9NQxKnZJnpbaPfKcBi
q8idtUHX4QRt9TfXCVpAq98d5sdIdBZbukBMA3AdaiwvwKMSO4HwsbCvLCgFgyowI4R9gKNJwpF8
dCCbWaypUWAhAUKRTsWpP2B7xnKjzkrSKQVZbLFg6MVp/tR6M2ieJ7chHJdzMdfOhaVL0MVJpDWo
qhoj08vv5MzxSlUtVvzOYM17A1Fh+IxTSMAMmiD/VuHbfvlvvBzILdWlyh9uR2Dhl9hST4Vu8k6r
mggtrmsWe92R6+yZLW8duHHRdSwqy1kQcNKYYMQt9Vob/+aCZj4qgf9riVsr2zmps7+MqqtqSEHY
GHBA8uUaFDLljmbpLJFQ/qb8uNN49pqjAJ3/D0vbrETJzqYMGudRBiQ/cb/uHhOXpEAkfKhDFpPc
0L6FvSBzl08E+JYxc9uXfa/RMiZK3tz1RGb12dyn8JUFKIMhrkRWxbW4Q8MCG4X/7ss5BGV6ezb0
DnF5owPxHBwfRAD8Fh91vH7499FUWbu8iq+Zxjb2fV7GVlKbEajaZQ6vrR8DH8YV3TPF1TH/vsoT
6UFw51TjsWLcWinJa3TgfUw4dsEri2Cmp7em+/SOimTO3h2VjdAFaMnWzJ5/YVGP9Pn91relWFck
6nb9vgsmCgxBVoXVrWW3WoOJrDbizAd6Nybo0TzFk9osJzcIVHvA2iisEjmzxzpmnDpLhBl7IGg2
tigDat2PN6MeVL0fEVHSAHwk7xWmfm6wLGO4DSS8K7obUtdxqW3LxNgfppWLKKyHBMXYT0HwSyz8
FgWV6iDvkE4RIlOoYPUKJwskjzevflYgD51oX6UI/OnpImfR1tPZFnSzOfqE2dQ17QzhGzJBICSl
ifSoR/hTt3CWiLUnUoGL29OSulimSYb9Dy2sSke1lWYJwCstZO4yWxpwb4stzeBRJ1a1PU4Ung1U
H/5o4f3pBNVxfxHIbj3rwyuoi9rZBchzDUZ1a4rColz+KX8KMLwqLHo2hCE+CLJ4xo/RMQZW9VPK
EYtrrL7DK2AN6M1dnYfP0xQM/s5uFz1HZshTA6taHy2VWnWONwMmdAdlDOSxt80C8qydefvyF3BA
B+8S6YQocS1qdFTSYLZ8CcDuJqQaoLBIjxh90jBMpfFGHrm9hr6Vx85F9bNcbaDvllwvIONJaxPc
nl6upPpB7rCYMB7vauN54FjGPKqaFTSenhyjCA4CgBPtm7/WJI1zKISuLH0EMcJ6iV0jteKUO0y6
sUnK8fOIzN8QvNU/1j7fjylpai7LqaaHa76tESC+aByl6b5avxvE0KGI9/h31NS2JOHQs2W8MIcp
suF5DZbksxCH4TLH9aLVMxoxSHOc94G0Z2wLXdf8+fjkLBEiC7H1sSqFVeKvoaeeV54K3UsVjnEG
N2hMCZP0l/4SlbUsjrvqeeE+6VVFQgxvPsRG3fu2RhI52cmK7jk1jYthMj7l+nPa6+OxO1AU2KlI
BR92XYlCg3/sWPXfJQ6ekEAxd0ZrXeyKJGNCs99Kfwbt2wFceGD8zdsLW+FVIyjtNpt62qdOEFv2
ooQzLUC0lNz92z+lxKph/oEWOqX51NPTD4VhayEvgg9oFZ+ITC+2dd7S8NVly80kGzn0IERneOl6
wQJjG8IQI97IQCCeMIAUrR2sPQpOMiSRbuHJKO1LlazboQTNcJZpTYd2bphVZaN50t1m3AdelrRM
k7/RU8esdq9f5p2pYAwOEFLf+L4iVZQSc6YLe2L5vOawoxPn5I8h6Qxz7DWsMZ0tWElid9iflkRJ
PpNMI4OH8sRYHHdUgOGUbI3yZGKdsPczFR7nPmBpoP+13WJkUSRggUxunVRGyGqzVLjuPWrqB401
uk5qH1OfjVenJYMxMGzo3HwMYJ9Ap4UOeuoeYZM9DPKKDoArVVG9h9yz5vkAV6U4XzJ4SQvBAftN
rYrNfMhrzjI52aFVrPMAVovHzC6NKix6rcGx+k+xUgb81iVC9fz4Gm4RDZ1ifXzNyVJmwnmSo3km
YgukTuBOrqxRxXfmyQ4ACxB5ih/Lr72FPD5JVtfrUhZ8jmtgp7oj1sJZVuCH+wFlzqdIqFpzCa7r
M7qrnXXMmkB6bTfRKtWnTsa4K5MB3rJ+yeJ1zlPPvZqFq7Ckslwb/RQ7Xics9trSJuOftv7faWX/
KEMjK4mV0C+tZEJTue4mHvHTztx6uhg4vwHYCbc96llRCYdobntooM1i5da95+tBJiAbXNQyFPj7
f09fVst9wBBd/iWZPZd7uXJCAz5jB7M9ov20bxRTKZJRB2+EdBfl8x9iD0LKYn8AhYa942nSU8ko
7eYtOnQmpgFDDF7jS/YJgn4c5D77WjIXCy3PDe8j0DDA7qVWojLicAOITbz4Fw26u+oEbEh7OCta
/rZE549doF6h9SrdeqTPgUbsqUO+LC47bfqIwJq79sd7gKq0jv1Oi6yr1EL45u9YzrsQF3bfl5Ze
pQk98PHbS3np0uy4dzPpxYmbdmS3A86/NsQR9KdFTQ8BTIU9lO73dVSAvYUBLtXXu6HN3N6cyzk2
yCsOhmCY46CEWVHruPBCTyDGsemnKiD2+0BnoSIZEEDimYjbkSIW+QyCZTy/yfcShSscmGzsJ9Fd
UKB3NSzTWGHoX9ZRiJg=
`pragma protect end_protected
