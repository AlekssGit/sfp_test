`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
jS9cINBdLq6HHutjvhJQVpyJXQeGKkeaSJLDU/U9vxHegSqsARgdVqkqGEFPLwiZ
LSomyxaznBviIHqIHUopIvNvYuJWdYLywWUtYjMKjpeJ0FmB0zN2Lj+kiE09U1Oh
sWg3Zcvd0EWWPoCvAKKeH0pVyBnAgRAY1YwemlaG7KY=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2452544), data_block
SNBgIZMRb8p9g03I3AMftaxq3f/b4vkCACkAT70OC0T2zMQbEulztoTIljDkYz/9
GsFl6WY4yEo1r5LNE5cMDAf4zEHsuXdVKxQk2gls7Kkwbp6XxhTikdiUNCn8uPq6
cx7fP+cNJfDnTfjapxw7e/Dllc4tJRZzxMS4U4GkloZa3OnyEZx05zRr/SEz/UJI
nR8Kr6QS92g8ahiTwtnKEVDHIPyTGc8UNm8n0wA/TbcXKt9mP7mp1J+Pm85hnz7O
QFjS+OLKk1maJ13WgcisBFMFXTx+SJee5g14bylEnL/y4MkaJzoGFeJ6/rbFnBSv
plbnpv0QRXhQZtcyudchfdyYLNOuzYzxJK/RUXE/W2hPGp7kIOyOohby0byDY4B9
gZaddzywZsdf+04wWVsFQzxqpOTADXIqfQjtXVsvr0QAzP3Frisnuxz2l63Cqrcf
yJ7G7Cs+p3UPNXg1suphadCuwRmzsnBv/eGYH6lXWIBdKe5NZEK3PHF9r277cmv7
yV7jrOwzCscFQwHVZkmA9pYgJ4+GFU1RXM2npmhLT9qFG6iZRqZ/Ni5NsQeKcUEj
bHAb5gRZ1irjNy1IOxhKg6s2+Cw8ISuyu0uTlsfsOD4+mlD6qnWTGgDp/6fGKYSK
ByZWNyupReuv055tpq6Y0orEeE4HZWsy0omz0QTkpL670UdnUlymP70lM2vri/6C
dW4UItHso9QbzrFY+WGdtQfHAu6WxZngF65q1psKKy4/k/ll+y4ebl/HeAzdANNp
77NDxrsGHkCi3WxCNB4oT+tTzR+c2/DmivQ6yGfH/tRc1uaGCmp29PV1UKf9xRif
fBkrlaH5veTqacTagJ3GJy3B7zGK8Pn5bq1paXY5kmrCLiTk278GaGfenO0yFWvW
fgJJAdN5jvRkPR3HeGvObSkp/VIXdr44SKhF/Doj1ItKXsriQz4/Q7ZxZzK86Ouh
uSkm5EZBNXmZSGSxMF6DTfo9mFPrp5OxNcnw5Fat5FxTP/WeMlKD1vgsM4R30ITx
j8qs885kyOBr8sJitDV1nULnIGgbWaiRbKXPQTVMN1cffQEaY9GPHd5ZXeq7P5br
2FjYLnEzHscv51zO5IyhmBbuD/jkgRt2q0AplJdFlxvR6VR/0LQHvz4NXwdi/FQz
kdOz2Yqp2KlVuS8v0aLE7lQR62lb2lxIr6pzhrhSfQzsYlwKDjNDPmS8qYutQZ4D
nGkcDsaNxeywIk+qz/aSDfcvUx7EICKc02K4m73yrp3Kg/kUuP3s+aWgFsw0JaK0
lZQ+JuCvMcKM/LL3LAylkmPVGyqnu9YlwdBNzLcnttcpVtX9cJgBXhgl/xGuY5h0
vtEPj46aMPXcwqTX/W7NyYwpgZ/UCuX6aXf0BmmlYnLLPfajoH3Q4q3AIIseO1R5
nFWBVBlbpfmurNB3RxIqnsl2Uu2zp3s+djrNBInx4C7JoO+Fn9tYFRutviTynD/T
Y1j10XP/27O1SYUnDCkjfMUAdkeXiMD0y+m97zIPR/h3PtVGp5Zxg0XW/g31cIXF
is9VLftn7fwrgGrbb4W4QkhPABzF2WqaVT+hK6ug569DiD5FgYyS4q8EwMBs/rxj
H2h103miKA02qln7MV5eWTtFDSo13AGZd9+4TwAwliXEfzdc+LkhCXaENDaMA0/3
e7ats5FavvULbn01vc73Gar2Xy31IDMRfHchnQmhLPhVPZS6H45G+Jp7nTevrD1d
k/saEQhC8y/AD25APIOej64W+pJEdsJVsJ+Z3xJKj5aaXjT1TCZWeOrRuCPe+C4d
NhffowJbi2ZnhqeZVOzPPzA43Da0h0mImpYS537TtscIJJZqe3tvjaWY2RVls2pa
v96BLy81fh7vO1YODS1eFRrVMyHn9ugRcMrbM2ZLb5Jks35R595cJUYfCflN7jiJ
BGnkq5aSmuIT8nQSMPuW7eW4iIiacp0BAaUvQhc/qGf5he02pmMmy4TmohVBBsy4
fiwblT21k6FYKNJFH3JsErxG2hv0dAcQvArjsYXqcwby7FY6nkPLsSQb7ohWnfKq
djXEGpR5EAzXPz2p3dU1fchcn+79oElcT3VChUwgW3u1MM+tsrGOJTQGGTagVJuT
c8/8wNze2UDIiSDtAbgOGTW9LoB1HLbnhOFWTukET00GG9NijA0NdvH8a5aoewL7
Q8FdqQvTeRrTXZX5qiSJZdBSOtdOepQJs/TtXrCaSfMkWpbs3Upd0pAE+ezWVoU0
+jnwMpW+ro6m3exA5jDDvsMZ/qBIbHM0JXNTspRCjF13q9hPlWsgeju6JoesTYh3
Mk/O/7khsQuFeaNPsXBo7foCD4BLvOSJFJhbixAAGaupyO0V0E9Qf2wd1lGg0bTz
raPPH/61pULYZfRZY1W1h7rt6x3phzteXsGPuqy/MwOKkeuldJGzF/P4WRaFlcD3
sl/Dr0PVcUOGZygMGtm1Snn0cJjm5cW61L/pLTg+QPmkE2X6pf6F0Ve6xYp1lWkK
+/myEGujizzmUKIfVKcxYp7Sk8/6LFYXK9xSU8UqpPEPNX/v6mWV/XWq1kjMKqm6
fjH5noGrquNzveCeg6xzv1CiKl6f4mfuMGxc+H8r6iCPQltA0bmKh19dZX6Wp7ju
ICvloECtrShv/NDiZZHEe7TPjuMGsa0DQI7dOXHdZ3PMWUKM3z0r3hyrrQdKlqm+
IFKEPf0ipe5/VSlqrMHwT9b/nyLWMX0BIUctuQiLSyTfMFdiL+4wq+kLUJgCHaiw
GjbQlAPO34F5RaKfJFXhf6hfevvoI4wa5Wr2BNtJA0owguE5GFWYiGKFxdIVMykD
P251EbrnmTd8d9xFjuCsMC2oRflYhXmpZ+gPCKhy0T1QXcr4C7l7qxcjJh3hHUH+
K/6G83LxnBMAYaLC3B1NpuDdMonXfYBHFPkV5d8hNlq88IZ8e52oqgNHpNddkjRz
B2OwQW7pMFla3vFjGfxfqhu3hVLfjLTF5eyzQuTcVmgwmuHRlpg3apTrwefcsu+t
lKxeKEKtPiqkikULU9TUqqSZ3iL3e/h59q2OaN971ZteRPZNvw8hB1ib9foUy92t
+X/eMc69i4+UNOZaDuQcjmY9meW7QE++uAgTGkqu6LfVnlxrzT6bmBLariYMYEde
Qa7Rwuh932gAEl2x9XFZFxgjQ6RVm6pp6O+aobeFVmQImEKKFEf6s00Gt9hLwLKI
LvMfQTGsv15fi/r/bJsFFy5yqwk1446/pYIN2wnoaaqQ8kYpMIk32SdrHDZd/0JZ
SO/g9J/2js0rCwXjDwQzsV4rnBrv6tUbKSsGqOlsZUMvlzJxq3ovYw2YB8COWg8W
LRskhr16I2xRxLjzWDRJQx59IOC+NEHuTnxbbF5k7Eg2gT7N5p3oGx1+1IQMV+ce
TwiM9vjkJOTynXNBXpiXrJ6CoX2b+GBRLWFDyekz9Z3Scp2F/HJDHtOT3s3YTrfd
2UXEf55pBtJSAtqSmJBbRhcBXu7AF9UAQypBfhqu0e6SvcwGYAAkFpuysJzeiz21
hVf/cYtOcdUxIKlXnPh7Tk4DwceXMExFCkg795Zi7Yt3KYXeIAky/ERXZrCfYLCF
m00TcGufT7tZT0JcRPW5bJrtqEWFWsf8SBhUv3es50C3m9hkXlyG7EI8CzOlSikw
1ZsvT7YpoL0NoljuzitAWNfc+9+xPThPjgZyxCFEDUXJ4y+9K6TNmyjgJVEbWepT
+yEdNopmLofG5pQgRNgbhHO1LFyMCR3TlVer+c1V9BiYL+3c5YOuyM0ja/esQEg0
L35CKQSFzBbfKT1egBWuNfBl4CtcSShU++UQ8zZfTL/I+Bjhl6nsZ7HvdsHm+no5
fLc8n9aC1C498SIBS6pAparemS2FICE5K2gqGn+J25KMK5OOqEhzMk/I7ffnOkV4
3ahF6Nc5I5fvn5AOKghxmXBNMJYaw3wOcaCOl4tdli2CcDGDDpShr9YmJzOnqosK
KkGxMFtCq+rOAa150YjPPgM7VZfU95N/TwJzkstPwHjHt71GUWQLdR0NQicmR8QU
WCaogkB52PoUQ3AbBJh2DlklWpOe1v9YKHiDrVJBoNTJnBW/83wPSyvjso7r1j3Q
o7wixLjVO+s65e4sErE9+j5ivlI7rb3likf4XClmbSMBJSBKwihGJyeJUzg7wYFZ
hpZdnHoT1izuccpq2CGQrrJC2fnL0ubj1xm4wM/K9Od1Lxd5SbJwtlsPol4B+ZPf
RYqi8Aesap0wbQJMoE5qcP6J7C9dL5MLWNpPWkXn9dOMIKoZPYhJzHnrkzaZMOzA
BKASfjgYHaJAhITWn5UxDLycBpS7rJ8/M+9kHZU8Oy35zLdLXK7phEMttHdz3uZi
SvK724+eaLT4eNkQVdqo9Hpp7cqLX0vxKVp3baX0zIbeCjvUxkoC3QRNplX5TtwX
ULPoizqQX8l5eHtQOr9odg2OYXgeMNj885QXvxabK7aMMT7DbOgTavdDlz5BWOaX
/ESmZdRONjQFH54NGiJ4m+yG28yeW8sPbcFDYtw3SMYE0tjBU2PgFEd8gyvSs+k+
pXjOSVOLyBNEnv9DtsVfZZcTFCdBhRpGP5oCISIR26fM3j6q0I19h+V3lrJY1RW1
Cvc9uc3I95pXg39lgfI9zaHpxQxPBerS+uXSmfhVEKKF7vA0OKQwcJsfK4xXeLZN
Ndm6zlZGtkpfuz3Hbc47oZd7A0ILO8Ke7exvHLF6XaTXxghRV+tgbbj/EqEMC6SS
Jzj41VlzzZchM3pidm9rcEtcgeuvuFTcbfJUc6Z7JAOTOzCJH/SlrBAlUwmdBxDq
SuXvmoanX8FUyC8C7D60em1R3MdcyZu6n8m0MgNQj5AiNnP7X0KYu3TfDhVD/mla
QImUTu9SqP6KXRcKULaZI327WUmkjM6B4P45LibIc3bnr10pYgInpOrKQaNFsfM0
tOO8GrOfafdFkFTVA6GZZBhTW867Nj3BTR82U2/gap6t6KVhox9OwWPmq+xL689f
N060dslmZbwh45rTexD9zBt1GuvrKIyw7CfdZCD+AzDQR9ww64YOyQG4yih0FBpc
0+gic2/1KRnYyfS+eJPisD2ARyPMFPE5B6PYg4LAjaZRr1H7dIQquUxPb0ySHyO7
x2oJql21xwKKx3NOT6dPeJbuACbyuLYu650rmmIjal/8AMDP7nfUOVIdH0hPnhf0
PhLajGE1+Npeffhi5eYUwMKJn7jX1CiGdsAeeeKRA43/U6JR2BaFE8ZXt/KcTYJL
I7G592EMCC8JOP7/VGzK01C9b1vS5ABax/mbrbFFezyaJOREJQSw2t4JIOhU5rvq
xvo/QEN5H49qBlHdUmM/6kR0+ApEle/nPNNe2TzAcrvMasdLjkkQ9qBi571mcqyT
K5Jylj/G3xSdJ/QCSI0f2OZFHmqiuokdMifJ0lrGxSvOX5+QdeTHXPfNpLhT3KOT
3FMpLIBd6RpW/qAUBTa8lUMr76vRw6FPvGfOuPGCbWgZXdSJ+xBkGwFCtiCm5XcV
Ak5kB9TZ/NENSrGeOK0UjxmyVtnUJzqBJTf5/lLoBJkY2X5n1o5macMHzKoiFGc3
V1qvQs9TBo1MoHpVqq4QB1yLrLo+pEzFuTJ9G9JcudE/NLpsAD8oBI4BvVbIYtAR
qjuymI++7d/8Xji6fHqD5SbHnWTii5tsn1SLomgTP9WE15J49bCNatD9K4qQFu1Q
wOC/2sXHdSIfdRiEvjL+K5fW0RCFShF4ZvBgcqwCBA4so2Z3vWptHz9+rvC60HGA
19xuOAcsHoaT9LyFpAys2HBBb3MLg3DWJVMCE0DihGvmlyaUfdapd6g9dAGgtxgw
oRjv1Wfsj9jP50YR1DN6wFe6/v7qZdqPv5KdK4OQmroxKGP8behoiqYKrZZxSKNg
98z1kecnM5+N0Os1CQIWRDM6vBRIuw8s+uexiSx5O5MUwosHD3QG7if0Gg9/25C8
tvHgt2l0VkByTkM/auk1KI6nNQ0Z3wezKVfHFssc+AHx7H4e9VHKUhEqHUoC+hPm
CE2R9c+0rrSeGQihzWTGJF2jppFfS/WIM4p8YpAtOu6jDeDTSmRlvT1qk0rSg7du
/Fi6Zj1xEq5ehdWfawFaYNwBCnkMncueAcmwRFPYEUMv0wpQ3/leORLti9QNV3KV
ZjknyWJ3Oq5/SDgkTBYUYpfyNycfgCKxb6qq3xhAVTFyodXoDEzGlGlvDjyw6gsb
JkOKMAoB2CP5QB5knf7j5lPSl4AMe0fLopK6/+WICqmawaG7ljSMaV+ueEAYOUFI
kKU//nqT86IQ/mdGkY7ZAgau75YQBmjfEa1unPXVU6w6h0iMsgKH7iX0gDaYi6o8
S/bu5TgpSGiE0pa+Zcl/75ZrU5XjOKe2iKeHTS6hygi8ZqSN3zddI4Fg7z356NP7
uZefz/jYIcQ7rSANF2AgZGuDt46sYacQ1K1IYYUuYvFWs/TSZoJzoqOUwxLxLbPq
b74Fs1u+g+DB3s1IdBMQbgcUeC8RpPf10fiJuePDJThey3ekRmX+M6DAo2bUEqLG
Cr6/dIqK7KJSVkGPAMMXS1RIByB7pMFodFEA2UniTKQ7Dam4EuNuqJss7NHqHzYG
9GbVY9Pxqm/oOFcDDDbcVI9+j018pAG+Btlgwm7R96GAjh+88wagV29BTg0OCjdn
4n/L88ryh9bR4SU58q5qTcXa0rPlttrlexvV9EwUcsaWELTJiGT0kSky1Bbmv7+B
vwSl3AKT4FrRdDXdd5gxB/zhjkUnRMqFWD2qe/1yXTNnVVginBGq11yYSdxDduRz
FeOEW3Zrg1LOIu1ysF/fI4J025NpaivedCkJHu93EflQ1Uj79xi2YgEin2wiGlk/
DyIKWjhHxbG2REND29O8JpXR1nQIB1HxEx4P5oePJNmt+9H2569Q4TYp9xQvZXk5
LTuv33+tEGGMIniliDOWnl6zJY83D+Drq+jVgG+/o1vvgnuMc1M4tfSoacBKn51O
Ytpv7r6OZeGYRjHdKvKOEq6cNzGxI1vRO6NfEBfb3UsZ+vZrm630zC6Jc7IunHyT
/Lg1L+VbbW3oI8uuaWXcxC9+2RW+hN8N9/xxmNYtsApD9cv6Yvim5P7bZb+ypdJ5
G5jsnpzBe2gbJHf+mH5CCukBaik3xrLZX63iKaWTgZjDV+NoizaYUtEzxmhZhsXH
5qFkcCuM/9sqj4/DuZgBDH1sVCztYt1K1o2C6ZhFDXGySLQLof1ZvNHiw4le5Jhz
zrRJnP9gEihcfpvH3GtcCdXBrCDF0P3wz3567Z20dr1xVXYijkVW81Hr4Sml9TuT
8Ptznadig7wMYpdCbhrEb9nJRYuvwt2O7+uVheJTddqd1i24C8vKeHl3EqmFoRZW
Cs5eqhSMg9AmfnJj1sWdoGJIICBlkyDv6mupaCAyRAIcNI0NrnNrQHxXWQPfe2Rf
Zps93xP8lWE7UlKK8B/yqmqYcAiz/mhZPdG86vM9mlRaRXNwit0SUKGGEJ3EAoQK
ya0xcWK+Mvr1vIpMZ9QtN/nxZQibNioJiV1mePWQaTpT/XETzVSt2+vgRVHV8pai
TUI7G9E0I74wSqf65LHmFLt91SNfJEmK77YlpY1t/fJKGL7rdr02uIYJa8LPrH98
RHoMJS0NWXzjbc/IH6yoCTxrZQO47yBhLPSkAZWBeF0vTqYaEUwyhp7yhd4HgJUo
DgW3ArmyGDDgPriPAhTPiPuvhNCyJbND6rWz9rwgignbiTcERJ2+OQA491VYOru7
NHcW9kVULEGifoPQAiXyP/jiWEemg/gkXf7W7wLQi4Xl5ma+iHyj6dTtNNGMEnIq
5Hq48eA9MN0LOY2LmQqTQSdde1VlTqNZNzh6XMpjLjAOMBx0Qxc+pZ4e2WHJ+MCA
+c6gK2ZEzntyHYijBvFJxFfwkJ6TWGTWJYnyOV3I+DwtHBfElWwKOGMrxTr8OhWy
PM8kenQlrpiVVTUmZV/2nIu3Dk+n1nYnnBAzsEUuCJxLD+hY4Xm5/QAl+qXZcGy4
0Zj/7ZLuTRXcdLyO3cC9gnwSg7FVZfzyIulH8i5FlA56OYtHJsqPQ+ctZapHHi6d
SMJZAWCKh+LIgmxdW809LtC0bvnxcCnmci6pKd70LSLx9Cq6UTPEbCtcirA4CkKd
BeQ7rz1yy0y3jpJXzWUUzXnqwEfqVPLDObWiTxrSdc4UMstw4n3zXQCG/EqoLrdO
qSjqbjZ363TZ3+kyXQ5P0QC10uK47wtLGeRvI375GCXTi1p4PKIZSHXrdzmhBYe4
7NXUif7oW6qvC1BYiMQlH25orVWBc5K24GgEj6wSpwyJmai0tUcbqEWoAr+4iBFT
xcB1JvagC91A8y5siu9WUhHr8mwCPhbGU8MlfUPoOJ7Qja8JPaoVfjLIqfXY7hvi
NhQDnj5F7TbBsJFpZj31vAf63lUuWS78BnYpRTY75rT6l71WIHInhkI6aEWkS1x/
iIOybYC639PEXksTKy78M+EXL43ZmZoK8IAVxaiT7kHB3MlLNLU9NvftDoGXTg2b
Vl9Vg2S+UtLDXFYE5myv6gfuqHgh8rBn+5K7bDaz2fMEliJSRIa/aE5C6wKHi4tr
TDtjA+k8sKI/QwKAN8wTlR8zGSpOgc4ahkEL/Ldq0U84vp/LcRZKQmAMqjnXZoVL
a43A2c0zJmQVIr1OX55XHpR0HBPFmfLZM9WEp57nHcSP3+hljjcCLdlL/HQjO5tK
1M53qJWzKBnrFc3o5T1yEpH936ZSKo/rEwyEYkWG7+m/xumpnP/Zn3RvcIDNZo4g
haZTiETIk4zMaAINKPrarammO9DYgcmyZIlZ/3qYwcH33fDno4EEh468kF1zW/j7
3bfilknUbWWnhfusW0MJ+APK7UtMeMTTgyeXJ2EE+rgMEek/gjov7Yi+iTXO5Ydi
vLqLTs71JbOfltPsEz+vB1QEpMxK/JTgklU3vuxl1m8IPOCiyBTljFLLBIHcSVWS
pdFRfZsMv5vgHooyNgdCBTQZiISvIsr5fcUJvA6rmmWzB2Tts3qJhcmM9eV/ivFo
j2fIDXDacRGLNKs6o1XdLYBX88qyJTF9KICzi6jIiKMrLIvLJAMu578p28j4vKe0
oHo0NsyzZhAwscfFG0MqnNekVWV1Jfx2udFkIMR8zX8ohakqQPQzygXOtxqty9ja
hkyEd4vldeZ/78PiA+NYEsFElXItZKHmnUwUZ4i96NVHva1ZzpKM+Qy8qWgg7uyJ
SU4MQUfdY8QvHkTEZ5ilMLIiWF0Gl//zt9F/pSjFes76on+qTAMDTg8OSPbNgtTE
MWHlGPO7JpIP5J0VFLcnXoJ6wnaUR3cPhR/f+HOVibtlHDzO1DTH/JfPl663we4y
RnZKig69hwJF9vRpco5eYpJ6JXK/s0Mq1KQbA0GaN/nvogG+jUi01k6Wk08F3bYh
fXp5LlOxYWIz4c1rt4kFW+lZlVZaOu/4039SkAuT35uESPm4XMfCJ0SbNG1N46JR
skgzFjqTOEG/5TM2GrJbUDYNPl1AFkqfAXIhnKYqVlnSfnWb3s9DFej8S2dr5d9J
6xDctX37G2zX5gvhAvlxoiMeT/pAx1g6PZhXkiQMQysHhUcy09JLy3GQJ2GorfqJ
fmAwyL6CG3yRDhGbeFVcIwi2aDSG/gtCr+Gw0jcP++V7rToSU9swV55WIPuxkDur
X7tZ/BZEHlNiZpc6Rz1hGOwF/8ARfB381q+iOj37ulpogg8uzD28F697hkPnk0qj
LzM2dFQ0Ol5m65t2KELtpPmyF6m7MWYgK4rwfJvhi+NQu2EZHtP2H+vNjlVePgKP
lXLnlSZFYcUj/E/ZgG+4oq2S5rI+mmwwANzFlgwFonS2+1AOJ+GNaKS+jfHMFfJ7
0kVXyCJVmAAUrVo+FKE9yFxNX2xEK3+aSUMf9ujy4mZ1HtC19LBoLWgTBTB+xoiY
V5XeqAhIImU6+vLSdjGsgG8DUA1DVFGqSf7E5zwlpCWLLAN+WphDnKlFygZmSv1f
1KKNUQRZpO8D4iCN4NbPuzsDgA3XxKaoewRHlPxDtw28W3Q3EUPVtwf9K6fDmqQY
QzmtNlYXNCtbbhxkDmoYcUkrVRTVdmlgfRMDG6MMmJVQYcvTGp8Poqjz3qsiZ0ZX
0AibgaEfcEXOQ3BvBsUaJuvypv39Qy0yBLdb5kEQGNvlhRb/UPZKDoikVB09dSIF
GecCloK5Vr/bFvh63g36qP8vAG0xtZ67szveH5G+bXaBAe9P7+SGLMWDNUuClgwC
uDI1eCMuTk/EPR2MiSmXknDKtHYw32smWxo/L6qN6ded00CkmAWRsMUejVgXTotK
hCSQVnPb45UdCE+0JFzsmb/xKl9nazqRoJhzcURg8TBOiBFXIBgUwZM7oMgbAFvz
PKgZpF1w1yFuUoZ3mulgTF7GHrV7IOU2M3zULe+AwP1grLCXtqG0jV2hY/M3+iFA
tSc/S0PS8O/4/T9vweck9B+vqSJyWVfPydRTod/uw9kQBDLmUEFRqTnxm4rO4o5U
udF2jv+tOOUb7QPr0Yf/J7ocVwt6qEy6gL0nvajLz6H6hxZbpPWS2wDbS9mWCBAe
ub+hJbbNu37Wc7uXgLet0nRl2+G886gYFPwS98+ssRtOGmgyRrLJhDtQMd9qPv8x
W2vtRT2B2gd/Bnu4WrB3rbLc4ZXsK0Vor3bYhZ1+b8cPKaK6eBri1ubXa+bHujvS
ltzwn7llquPhH3t5hOgAMhEcURV9WZhLrpRMRJq9SlEXJyb3GTh9ltDlDc6tnv+U
KfUfdvGClNTZq/9NTVVicho0ZwxgmjTHr/vE88PpAux+Atwf+bj3fyXDA19b3+Hi
m5yI7nrm+zt0LXiHtLufJnRjcQBdBa09+jLjH5xGn1vaYdXAvcxBfsjp136O4ymh
qF/H2Ik6RGYItbQMA6nB8ECyiFl9k9klVJljiV3orSZGJU5jA5aFtZlOCCQN5p8a
/Ykg7vfef0KGYgbP0+rdoWZ/b98YHlF3c+oOyivIuesSey00I0aon/ykD25keMyr
4yTtBUBSPeazPg6rYADBLmdS2a5r/5LpLahSpl5e/SP5nn8SXxuzACx0jBHAtDjY
/tXjJM8Lgv4FzAoPVmlDTTAEFgetfip6nMdsUFWnhfkgQ4nuxlMtYoSnF8t0HT7Z
EHWTSKgmEwndNwBvbWZEyK00ndRsp6wrvQcMEFjOp9tBD14aYyXxE26zb0CD6QM4
uGUnu52Cs2CpNSoC76es1jede6gXj8VW9iGdvPJTRJzHmtLvyc9IkNIpE3O8VVMS
NxE+qjPYkfOdj7HqOgt/L0TE432llO/xRDWXuXgxU0eshfjSXcmxOtgmaPe0Cob5
U1Uz/zrzsJYXJkw+z68F4R+ErCaEKMq+o9tqcXzTrhNEG+toLlckK0ipTwa2hkAi
WEMrDPhMiVkYYoEtNPn8Kueaw0mf1vJczsP05+4sOEuh3MF474Cms8d9axVMCsdW
lanoJkiOLHnSyNKrG9c1iIXzkuqYy/a7BdQDcWsl/1h/9hPcaQME550tSfA+nkjv
NDMA1bOPITw7T2tJSvbmRCQe7UKBft3UgAfb3lWgVwSnkKixvV5hQv0VnCBWQsGE
yl5pyU2dzQKtOp/T+tWCNDgbDiFk3kz/NkC+jzHm42Mq7MofM7MpdESz1dcQW7kY
u73S+fqi7aMllu/t1td+VWQEj4EhkRBrqDV82LPPSlPZSPnnED2gBS6iARQo8RRZ
KjRXDOezbD2VVgJV2gdmxmTbedu5LCKlSY4L2VNi2521yNc9srF3K/jPMaA2Ucv+
XpkHggzh6XM1zxeJrdYnEHkXpMrQEAyTnUQ9uTi8DVZm8hjcapaKaHnoOJauJCty
nCrHLwAf3bI7AaZIbbzgnC6n7NAVitVw699qgDk6fIbVa5gZQJoG1um5ibCkjdBs
54B/fjzQgzRv27yAKMSCtyNTJwkzS9uN6UcNVFtAEYNVnkNDUH7P5P1993R/zLqJ
t2BF8T7CFQzhrLyesXP8TjRN4naRmxc8DUtT0VOdmx9/gU81QfZOdUHQwHzt3hbW
Y1X+QkRHXlqomLU6S6E8pss/XhsDvgzUoZ2gNvQVLrQkVf7Gtzx1yI2evvKITsC4
O/88SackzNStfif5QNQ2Egbn02FnKsBYIaHdqOnpB6hKSkVtV7KKV8fX/DiQ17jb
51So+gGvLnGepT9Rl1W4/7HdywLYxonRDlr6pPd3nFYefHVFfxv7RzMUxpfxMu3D
L4zE2CE8I6VpI9QFzYHbtX0krbMw/xK3iuQ2bPnTgwyFJqfXHxfhFl0S2AVTns0U
lpE4W8fZcXQFkVd47mk6YF18wAp0lNMmqAh3zXOPJRYL6DNf6iDJyAP1o2qn/aPx
g2Kw4TGHAYJog0z8WE/9zaDdG6t91kNbN1D/8cYvX/Y/OORPFDLSm4b6i6EPxX+6
YzrcX6qkpbpSS53x0h+PAG0HRhtCcu355gSoVZlSZdYNlbbQ4/MVsb/VaOEcjQlv
o7QdSG+rOElwRd97k7zjCPC2gXC7Eek+1FUkdX51IGoY4TXyLzA4Ft+J7oi7ndfz
XIzwlCuYwGNzDFAhC+roT+zxIx4z5vYo9XaJUzgWqd+jtkPaEM1GoFb9r16PIjm4
9PwgPHetURe6doYcpAb5bHzFexTB6YwFYvIa+cj3daGV118Pth7bx9zSgAXTxqFR
0qpaR3KMspdhlLJ/isRbG0+dm7buJmp2KWXqYmKsopTU9s06idDZHXtWpaBzPI71
Q11iRPCAJzlzNE8hso7f5pcmNMPP0jGyrUxZWweX1iFGyZCNmumAUNmZfMWkFtVr
uUrb4o4sN5igyhdEiCTaF6i8+1hUJptzi6sjZEfnlFj9UlSlzb3FTVnT25Qc4XBi
onehigDeAwkScRaolMd/DpkiVQlgiostMZcoEtO1+0z8PEdcS7+5hkj1R5PRY5Ao
hl40dRa4ftVDdGBl0bBcZuOPYcB/gbSgW0OvTmTNzWq3xLgmg0v4GapGeRN+VKN2
XBU1aO1oVau7k1xyLE9IeSwKPSANd/rT+L8EUT2lIM+KmNMFOc72R+0NATlI3KA6
azGNO8t8wfubTxl6LnUapL/xC08cAMl1ydFUE2ru9ElQXB+RSVE39GL6Mdy/s1Ho
cBm/UVH+X+2H50bJiBzhTnTB9boGV92wHjcr8dov5wTTFYLPZtyIlu6Yh7A6xWLh
rBV+MShFWVBCU/uy39Pvv8DvNfba43/H+jjFM6EDJFjB2FPg1j8WghvtpF3w1l+T
559iL3B7Tw6nmt2FMjBGvHU7OQ1EuUu6oUka4M95f63zWfTM9XzLhSR/oURYpogY
Klm1VVOGxpkLJ1hInScEygRRsitP1swkUsYVcVcfdmKhCEaJBhICmbaekbdiw+wy
q3IUrZrnLf8WNHLwBt1gjCObLS2WKoMxNLGCCRdG8y+YVDeMy9BTeRhMFoRNw/z6
igFYqL1aUk8JlfFXmbNto6V8gTalsnwLgSCU3Bxt/w50otyNYtVdMNhJ91y4Hjut
V726a5s7SVCkzn3/fDE2rt0pNxUk2Z/GLKRuYRsO0YKC4jBVRL1QxYg50rTU5+f+
FFRXJUbjnFPjAK0d9RDAQq05Uqv1Z4/bKka5ODS81vf2IeQjG/40NQgJi14oUAl2
jIyTgbyY8/30QgiIHLnAx9bo6BOmhoBUM+nGj4Y9onTnt+VSGh/FkPXXtq6o7t0E
sGVXioYwrKIk8/1qvM1Vwu6Hj5BclW4DZS2K5vlbC3clYzFuElYNg8R2tC5S+m8O
0NNrSHzwr5T/P1scXc2Mzbv57XjAlDML0MF9qo1QUIDnANEnbeqVxLIKgl9pR8iu
BRd9vnDCyeZ941z7qh9tBToY4FuMkUtXvSQsU/8y9EV90xTXMnmXWd9//6//yf/9
SRReYrgKjOsr9oFHw8lhN6cl9VooN4xTUb9/UVhdYF4BQqCkINDlrhHQlJXvPdYQ
u5mmGiLx4NwomSW/ITjDgNEKbwdF2lqrN6d4U2dcBrqvCMBVVKt4q3W5nD0T8xnH
mleQhHsztHgKqJ06aC/N/51gTnrju/GMRZOkE4aQqwd5znuuDfstad0WOtxHr7br
f1yZxCDbmy9fVzrW0f++4NMuFprmSIu7kwRoj0L9Jwo8tc/1F/BDF7aZZUCh4iUg
PyhUIg0EyfJ4laXVG72+xrzaXyBJv8TZAqiijEqP+Q3Cet2wEiDRm5/VH0eyyrya
t+e/8Pb26BLqd4c1Vql0JP4SJ3ozWeuFSWugmUMJN8bi3TwPxumi9xj+A+Z2wzIQ
gCzyz6sJn8zTQcBbSHZbFcRJ3uEtB2tELLEdIoXZXoY6SfsupjLETIAWANVW9o4O
1OJYmxVQBeHycjOYA/Z3QQvHr1d5CGQ5J0YJKvwg74CvhekytPeOAIqluFVuE6yX
RABZI790kvu1UyG/mJOd449KTpO5rnxmyuIQZd5J+zuK7lzSZJv7bkui9SZ1PK4w
udxvdIEdgsc/tPowzEYNsyidWSoHU9JNYphH/VoAqxHX5ZwCgVrymJ1DoK63aLlq
NsOLhWb6VkiH0/ZPStsfwRFyuIX/Ladwota7tQOoh4nvyHCFtj7eMVooB0hdW1fn
xeki4FDiH6ao1RRq6zxJgtb6s+1I1qjSTXRa+vEirxCYCo39QU1L03JmdpRSiEQY
/XyI2jcJWOoMkUxgxdH74O8DQaQ5T7s8WxMr0KZfleUQkz0fcCh3Pxhzo3AoGmtD
cOgj0IDzLr5tboLtLkOd/PCoAPUTbs+/HDxzCxDfz8NvjRV4om1JSKBu10c/LRR0
x3H0U40ugaddCoUGEhiYyhpqPAZKDF5Y36mBjrBQPkhW/mcL5h13IPbOHD11BS7l
j3dXesA+Ceku9fbsDdYWP3dJ+9iCOIpLKem8c5m1ep3NVmILWmAcRqcfH9QFt/82
q+d06KLQO+oAaToG5aUiMwFkcPdKTLHTgPHI4/0MJYtb8QCKyuCt/5dkpV/gb5Ds
g8TByzrH9RAWX/OhPfH3HeRHx21UpTwGHbe741CmGE4q8gfXDtYVBgBNjCwMsrVD
zjQco9MRhb5dFDYm+PpsA9b1Qpcc2UE9HUQwfSxqKTEwxAX7adNDqH/ZcpKalZYZ
fIxbDAnPoqZQh/7IlJFGvxCRVM2+L95OR3Una1u3BhhGqdEcHI+bykQHRDR1zHrW
COm3y/id+u+CYe1ALfZSLKUEQ7rrcBJq/difZvRTv3pD3E3EupBFBjKwnzIx9eQE
kPeFraSE2PYK/1MC/HlNAPwkcpnmIw+961A3hAGamjUyPzMOmBCAX9hn0LxptEEs
KYoEdmcn8R/Q19jjPwrSfsqJCPsHkQ6txYs/pWwhPvq4jRnmZyCF5zdmx2RRFV93
Oh9UZo8oaMam6m/ANoLSERcuHo83oOR6spX7cpArFgGnIzfQMfJ8y2ONrnT5B/S8
dfQvWyK5+9Ep518Pxoy+Op+wT1LckCtdIndyZZzQafV4tJdVCf0KOnDTe/26Peiv
Cv0s7R8SewTWpgBt0D19T3mcOnqK2vLpIWpuqam/beOFyYvEYFDPJ4az5bAXzR8V
PyAcTQffLFdYa10gdgzNUj6buvKjbwni24diJLTg4TH+FS+wxDksRxNQLR2zZjRs
OcgcAmtkeFOnqEbUyTlRjkvuA/SK1C9V8qwmBZ8l/U2Z9fh+mLonMM/s5yldpJDM
R6mnTI1rjDId2ob8fnUoKr8yaBsg5aw4/RcUIOODfVSz9m/jV5o4VBERGkWvSakg
guonTR0Fj6diK415Lw4TP+O70oUKooEfAaSGUf+yK9XmyWzSLQCVWAvr7RoPZI/j
jY67JHB8y7kVA0R9O5tTeUV3YFmqKQR3jBb4LbE6S86AFzgpU5lPRF25qrcom8Ht
OI4la5i6kAMs+MHa+zZvoDG1c4cOK0m61aE2J1TiicSNX2Bid5TFecZHUP//eRVM
7AjdoI2kshkXHq0LkYJOLIPSo1fD0vN+UGrJ2h2/m/VWg7CwuWgkAubPYeLlXpP7
+KP6eiy8JvDTJoUTr/m5AKHf7N2BeHtHw9Hh6ibA++OYEcQmWNrbhxpW+tQUkmHw
j1hpy/ykbXJJnH8LOX3lvTdd168cZUAjwi5Gpv06kAF7Ll+AXoQlRkMjLpxUWepT
aItqfGcFY2nYy8tFQzNzrCLYaNdnfDUCYwo/Tn4C3dInGQOnHY5Cq6Zkw0bWM6Ut
VUaWVt+/WS2gbnhnM3wFw+opI0HcGhiP0w8gi8Olbd4UAXmJwplUc7Vsphu0nFdS
WU0IOFOfg1UYG4GO4N/RaVJ3LpWjftNjGaBkQAlSJGLyIymUJ6LDpOPzphdzF31b
14f48vP30kIyxaqiX2/1QRBr4uf68JTWShyBP/9DdqAout13ErZdVuxHN6PhaCVl
yndZkYWDIF4WJ392Vc0Qy5K3uwbvireVYcVYbeVz9Lf87hJfOtp7+eYDUVpoqUNF
f8MxEqRqUVUa9nXd8lGtVAc5hRI3DXGAFbAy1TBJXoTGZt7bZVtNqbwTjvHgUlhg
592s+FstWxy0nZVhnBAFvl7C61Rlmdao0xfDfTNIcar2olBxx5SGJykGQqFu0R19
NlMuYLf5CjbLSvRY2iXvGJ92DgXQq/NWetJc2cTqE8Koqfe4l58TKD9rj6ib+7mV
duT+M07SaUxqg9p7FD5dZobp6+qYf/ZlLZr32wUSfqOe09Ft+PKFUN5VjWjDl/vN
KLAWEHnpLwfzjTDTSApz4xLeA5D6rIfViZGjJGUJY5iyAXqK9PzVdxHfR1Gr4mi2
HuHOmqKUmejcvMv82q/6AucgO8Zt8ZoA05oWY6Rb6rEzFXrmtJfA1KT3AdcILfNd
irOlqrmbLYbs8Y7HHISELgHto5fjfITL44lteM/yyFcSo0eDOTWGEW5QScuMNwRE
f4+Jqj19UBi4oOkprhGCM9fR7iW1sWbLfbjSoqITUQUh3tVXx/SdRhr8m1lOLRZh
zJoYV4kOLgChezUh/5BN0FjRqk0iW7hvAS6O3B8265XlKDnmRNIME3cz0AgCSpln
IQd6cQJXN4odFAltEm8p+oT5T88HoJ+kIclSiLOmiqn1/HuAG2BE9c5QxbSeTqua
6gsodlfOGkA78WD6ZAmzogOxZ2gk+H+RApc3lF/j2yzfK0ZgyG0nN5hMJDCV6bVt
PXVdfoarWXkHQO0Vlruh+4HRNckOGvQNf31MjAYxlMJFFiTMu8ljYoMZvzaWcaa2
68qwZxoJoevqCDr2EOx+B1r8zb4U8nO8YBF+wo7yU4T+zSeW7fNe99FeisacDF3c
08AMk9DO6SXPdws1uO5qP2A1nXP+XZ21KUlT/5iUK0D4b7B1qCaCGcJQWiHXNfMd
JflTJrDwy9xXiyW+8Wj+f4sTOAIYM+OHBRfGCQ+PbwmPiDm4A713rjHipbxi3U7W
TQb8bMjsHjlYnsa4ME20Yi1KBrPqMcPw/9xV8wPS0dZpjZ8Isy5UQHgVgsgccma1
WLMzSXr2yejP8iuhDnUOG2NKbzf3R2QjUPC1ZHzwabHFOz2uCMecA/zy1Dlo737J
m/C9A9/wYjy2WbTqMg46UZwPQ9ZKO52s5dMZqYf0ZQiYRU5l2LhH3zB8D6DOZKDo
NSiNytGTEby7xakmOi9rcxY3+KU/plGUUecUdnUMHew8ZEX1A3UPhgRTsCpjVkB7
VGMxqVKZlt5jt/47JxcOZNHuXx4Mc+rnScwC2rQTabWgW1wW1z2+HsIDKOcWhXvu
r1wQC7S3G06PQib9ff3ppSV58wB3ea+b1gLuG6Rd21Uk/wTbL+CvpDTlTWrEriGJ
RAJ4BGAYqachHHg8Crd+LM7GgGeH0yxlWxDfW7pZuEiuJP56zAjV9jjRO3Ak4Edi
FNXgPj5EwWk2pWilgHMPA7NWYnhuXOqKeJMgkVn09isqTriEnAM6OGCfggNP279i
yv7fApkxmY86q/0Wf4I4OG6+Vn0EdaSb+FunwuqL6Wq2uX2yg52Bz0NdEu/nfPKm
rIh0qngsYaOzaUHEf/lZNx70w5TDPx7WKZmjX6UAFrka+rDuCYwtQGELfS1gfD6q
ix7T6GB90AAI5ljIETS6DewPZr8SpkVLPKId9OmEkVRFMsGSmJcxzyKGQjDcIuzg
dA30ayNdNFJs0+J+bmqUdpPPTUo4rYNHmwDFdYFxK6bJB15LGvThkBHvdVGOcsCI
++2u6b0rG6A7EC0pSukv6ST5uQ8fRpFht17OFawobJfNhlioJqsc5MIUGUURp0AC
e2zNYw/ava+PDnATLg0VSwJfX1BokwSksa0xjrF/qfYC79Qq/5uwcD7SsKoYafXw
BakM7qaz6sIDH+Cdz68T1G8gAyrELG//l6wYtz1GLGCkCWRxJt57krNGV+M28/OQ
XhLMZeG0NhlSLJOKgojC1X57vbqv4w2wgZ0zC43mmmmc9lFFkS5QFMwm59VmwEe8
dHDBL72j8M9FVjfrmAbkrjLjMW7aJwseIq8+f+9BESmcFoOE5dQJdYx2lbK2Evbg
5fAaTPJc+GMr9MIYNl152hG49E14pD1Q+f3eaLubqfH+45N0m5OpanEYP/D5TvlN
Psi6LhMODb7589AxKLas699/xCBFxNIsusoAh5obVqB2XYrxXKBsLJbcK0OTBYYu
ICfKTOBdDFG+0bhxEAniiFxGUliE0Z/UayQKiNHrlPJAYbsHGCLafTXmcGFplnQn
RFRILbhgmF0wLKTD5ukjcCdOS4A5QAg2cr1J1litGTQksfaD05nAUm4w7in9HQc6
nm4YTkZpYWBGDgKQEkbh9PVv1zW/jX0ZGTvTkZ2/P+32jU0t39ne7LKZxwF82mqj
WvWhvFj6N7id4P7RwRZjlb8eDnqfscDLMYMs/8DJ57V1hgnUhFSsCHeSdx333ckM
W11Kw6JNlm/rI34Gyn3/ZrvsxYeqg4mHpA+h/TZJVghSGOHw2rbH986ZR+bYWLZX
inhOMYrSz7U/2WBhZlcoVTj0cNKjznFIDgn7Aojha3HBVSCZeq941xK2dKyGpGV0
lErLS2n5gmog9EKvjS2S0tqARGl/NmMtxwcqJ2e+wfTwijDk7uIoTBfBNtJOF5Bo
cMDMHHGFOdCYls1iYy3veqjy2sem9XtN9iRTMtUIGyu0uKZmB5cdywzQcg4mjH+4
V2mxjk9NruabSIUDFqgI1luyHgrbWY8Qnh/7Ma12swNbvPb+vWlE5BGNF+9PFeeW
SfugzrovAZRaJliCtNVY7x7i0q21gMip8plsxmOT2gTcdemGJQqZ83u1iritmsv6
xP01zdAqMW7sdLrvl5mivcmgOLzhqNgg5OBkTg4ebNjJN1iztxxS4ULUNir83bCP
lbIObXZL3jiiZR6YzpXnXsWcAUrZwKovmAztex2UqHYpX7a7mMgHMFIjZHP/HXfa
pd6xZlaGljhbIdvQE+WihtxzeW80SzQ5q5GlYZoLhKI79/N8Jvw9VuaGEuGYCEt0
InPDF607O35jh25str7P9dLFVh0Jj1KELb5xCMQfkbSGHmYq8wnrvBvDYTDXhYGq
rro7yfjzRFPDq7otlYbtpQ3YKmm1+RtnHtfLb6cYR95W0Jk99vT36qQFI47a3E0A
RM7k0TYjVWx7R4H+MqNyVvGdPVc/MW1z8lQdi2xLEGXhKpB56/r4WDSVHGv5ePRD
jUE066lVzUd9PPK5+z69bxLbDadUdBVannmbFaOhpLHE5db2yE/t6E13AO5KAX0M
+w2c6rbIWmhpbx9jPkuGb3dlH/HWSjj44q+O84P+AwWDtvaK6hb8KkRQpFhQzzg7
+5NA6+1xEJb2ruy3ijmFCk1aGNk1CthHfn69/BhAhZwob2h9NdVl+O9ITrInK8s2
8kFhfaUuDRgM5oKXgzzxDE9q162L87wfMA49VNOOY/1GUsnU7BWQN7ep+gVHhwZI
PJJAxX+I/gBAbF4UfiJCTLKyWUay4YEpQ21IrhV6OfYDdkhK9YZIc5pwUpFy2nwG
2He+A3tBN1m4QPRhiFAeNjPQz0NUDkgS6nSyCxl19wPCS8paKJZ4WHaU92FrREk7
3N5V1J+iBdtiApNGs1KSfnImtxIu0sHNOVYMsckZLu0YTTO+S9deNwGRVA/XXqI2
JhnSfcLoWFjay2Irl/KyEMsPAkL0cCqnbaGXy+AFWnRvcWg4pdyCsvTL271p5vmB
gfZ8oCJjJ7zk6gZuN4hFDWi89HDb7BNflJeo4pH9tMSodYkAonHoOEXMvDYNdFj5
Ahw7vMuD0jMWy9F49IDg6NhxOwf+4b3K6TMfTPu0mrT6hxbhU50Qmc3qI7UiiwVN
qZVPH/9bJWdDuITKxRdacpOO7uqmVh59wjjTGZHBqos/IfpDM4VRn0FICZgvav0k
pRpj+nb/jkzWCPwYfWKLq0GrcbT+zcj3vihhm6U7vfxUbssmnayCD5V9e6ptnYwu
QVRYcez5sffrDkxrgj1G5QchTy2+taP2fs10dJfp+G7CX0CsdBY+qD+ejOiFgDcd
AoxYZveusjCWlw+NcEl3xM2faDEoJB3TeUpPi0f+Z/hhHA8Rvd5FGCDmLP89OmT6
Oic7xcjzip17xscDgYmbTguwX70ezo5281mIakHLqnB3RrCbaoCx5qSTTu89igZp
6Ty3uXyrolxC2rY3XThXON2VErtBrQQU8tD2LMDybF5vE0k9x8EuNx9oaVIqbkQc
aNCpIgr8UIB9NUa8qFPlE5HxAnB+fif0loLfPLKXpivumy68Pw45I1g5Om7HmOZz
sbGYtL3rJMrKQKTck/i0rrCmz4vSf41Yjq/YQIcd3FGQdGhbQtiFxJicId6QSOTV
rynj7wgdHcmmd5A+L86L5i0hIaq6194VkFBcbExM1DqAGaFsIymEswqLSxFYni+b
UWz6QmkX/9/SFyoj77jKQjdXhtTZb5Szq9J3WyN+FsK0owba6E9HiVOnHN0BE8vB
ym+Nk0uJ+/ffzpC/PVy8xE6+3Wf3XPrKF3Tu0hkCm4iXdU1uxvxcOZtlvi5hPdMT
e9Int1EoVbuvLoImbfj9ALMqYumso+TjV5bi3C/wFQWePOnA2eJC/0Qe//CNOlnJ
MOTMGxKkfYRfrcjkByJdcbqzQ0l9jBb/Jogv30xQdf8D7f9mn50uPf+Naq1huPbI
TjgeWzVUawsp2lvU7BZPsDYe7Tew7Q42+q3GtETEbRerqT7EGQLB8tQfbNblQ2Bp
rhXHqUZlShTcgUSanu15JuWCcvao0ZpA1Aq5M6qZxpFQ58LDhr8428zh8QEcXsqV
to0nhsbsoKiXlyb00ZShnROwlKWILJyAkIi6byMkHzMzPEorMCFGhzeEbjTnJyPQ
RbLKn1H7KLV0rqqQs307+wXjQvd0YTlyFEw/X4Ql9mQQAhIYvPhYgwBdcQ5qg/eH
E8GKE78ELpkVBNB5mNGW8mo/YpdiAnBjSb2pY5x5yqMEx41QuZxRBV9JVbxtAti0
waNssAoo3Q7X+xHeASZI24MY18Dbg2O6JxKnGJSz04CfN+xwVwQgpWMhLJf3e6LA
HwC3Z6dZwMnvvpQoM6hV8yjU2g8ldMmgpoApfqfLzX2VAf/sbSZZaVt848LdRmda
3obR6rnLI9UmBiEdju29PYiQA1DV2zsR+0sw9NChCkdJ6w8EhdytlgdeOuXV7U3G
nVBPu6skb2MQ4lKo+6DCWMnDEYDjc0O6QBshzV6KnX8W7JCU/stSkxNArraFB4MK
VCRYf4NVluMPmRaJFTteE0AzwThEa6297YZBowTJEMP8PWX8GSXdewOASJrY/zeA
0ebK2ukYX6MnZweB8MSmovmaEvDuMLf8vJzaNPDdnZEbntOkoQiIgVePk6zOCBSD
7VUc0EPhGEwTsi2kbiwSDKsrtO2ZMMByrknjaHkdukGuk+QFhk4n7wWXT2yxKnBZ
m9KK3+QOW1r/XrU6ZK6gZL46E+AjB9Y88h/Nr6TGblOKtUWrtHaUTITtrKNPYODb
9pzpuREZkEvDSJmuD0R43M6MTAcl4z94x1LHTuenv1tLV3ySKLnzGTx3KajEk3wY
jLLpunz/+nQT/8x+cHDhO6hKoCqhFGAPL+t5x7aHSIzeAE5upcU0T8uX8Szuto3A
gUpMXGlpl5cyv0TUsvh6m9W/wvMA/e91o7vtgg8oYJ1NdZL00rve1ovFSaS+XatS
4kUXUXKEbudTBUzYOBBThtuAFGHrFGuJf4LHbXZMm4w0DPMustkCrEi1UY3UIwFe
bjfbg+BTjSK9nV+kjAVmKUF9Z2eq4xn7sWqekjQt/RopcLClOhlbQIgfAbotE6Jq
SEX/7bCi+AJWfhKWT074H0hvlcSx9AnNOayPz9bg3ln6bnY5Z3cWYLDCSpSRBb1H
ctuDL3kX8qD60m+fX+cB5SVgTygmEeQ3W+h8OIhiHxBm2ezGjXgJF33mGmYp0X4F
o6DCEDxeLl/tRq4xrDDCar5ZFW1oHdIViOL/s8xHtvOwkRkvhWIeLo0myX7KYVXi
F00mUXrpULUa90XSquzPLydPmzzrwymrgc6OkjpMCo55g52oJKg06SqR5uolI5wJ
CS3yVMNIkuVvdgwrZKZ4/cdPEHBgLTWAKeSlgLoXtIVtaPv1p0gQOVnCGOtlNPBq
WGnLLu5cuA5dwjpKeeKXVSSbQ0C8qNLCPNxNAdA0cp9NbQO5XwvwD5DGL19BGU6X
7K8AN39yUh6sqzOCtL4Qg4Gpbzr0OeB2nNgvPfAltmXKUaygMNyITv1yMY/8ZlVN
1XkK8j411Y9qJA6vI50wzlJBQTvIHSC+9qaFkY9EKKpti4rG5N1j3ljDkn/eL0FV
vu0z4J/vntT2okRBTWqcjxVp2Dg3m0HFdfXRJ+1LJG3FcmRfDIaY0Y4FQd+ma3dg
Zx4AD4U0pjpcNWcgLOoP6zUDAhA+0XB4V/CV0Z3EY/jTbVxz9CxLSGPviCUKeG3d
vDc0zFX1s/kpP8qlyU5iKoKbHJQJ78ThfayDzks/cG9pU20lhhDn9f4bvHh4gQTq
kh5H4nAEoM+Z0QfnYMYz38f4qG45irg9id5xw4K2Bz/IHlNawYroC8fznmGToCrD
HZnfAUhXDF6sWRj7Y9Gqb3J1r+UlXcnpWntTpm5sLjrGdvLnE5LqECwANvB3g0E0
7i3hsHqO3OvoUy9Wgzb4cGJejWGDoN/0QIhK04OQGMFD1Q6wyH9w5J09MZ9I9Nah
fh5aW++0kBG5tED0ZeOX6N4z+S2eglvw0hBa5OxgqfNx7/q3OHRHhMSo5priZAbm
XSBZBHG/KC0lZ554g8qDioTovKCkY+F0BZaXLj4Kat6YVKejXeXb+dOPU/mLz5E9
/fae9l1S/cS+1p+8UtfcXAGJENVZ67/TtQa19vRK+FalGYMwakVfD/Qlugfs9AgR
EcWOpd+57skFw21qWte0zrgEg/IVLRS3xWwcxNYX6dKf4r+tgMZQkHou2Eq30Xjv
2NWufDWfCshgOotQJvtZoBmlOdBAy1MrGfMNRUHv9GpJXLn1Qgh4NiJvbDyD0WSZ
iutnh4Aw/UXKuy9G9uSadW00lPyejtrwCvd0qZ3WN1/XrQkntaEYmdiBBkSWPrnc
iI92jcvNotRwp94mvauwMLr0gA05bQHjCZ+ExCBsog0jCXhgqqARN3+Zn+MI9cdF
C4YbDzxc4bpgh9x1rjZ3OY0crXSL2VV4HIu9/yv9PmDkDjQk9tiE8DUyVlG7G2St
k80HaGGljFmU7i5sNauF780WEYPBjS7HUpJ99O4YABT+ATyGnN/zAvBd/pSYHoS/
lMHaHPU6CDjz1xYupmYVglbJFDmUw+wkYl+deHS7DnMUdTXAQitwBPsVHdw6G5CC
QDqlNAnE14dSYAuWJn8fCT7FeIvlD9TspIlAuBJkMsAMJNsFr9ZPUSCj6SgymRcb
x6859ea3A62/ELt4aJHDIWsJBcWj2P7M2pNMg4rKxLBZo3MageR6C5U0ivJa/3pS
hmIY/35mcMcT0AzaP/wkWT8GT3QXEWZ0zZBW4LaxkC1x6hWd9ITbjvin1CgXhA2w
TiRxSlCloFfIHZzbC5ZW+vixEjkutZIagRZZJ3kteG+1O+qbecV1hO8K0zJFVz5E
Mup32EySWIYH59hMaHp4AqRtBGS0FPal+jS+vjAO2Pyt14I64Vy7Y5fOPLYxSiVZ
y74s4KCBfALNwJubFLcpfxVkvQvbvdZ1jDqWaMcfDhJ7SsXH9X6q8+fd5TOARa+W
Z41XpOXIefOUV3I2xHuPBMtIVybTzvP9P641uuwp+bdTm7fniqiF8p/AotC6QvXm
qjIG7BC3sNGW83fQgt0sZGqwTztrUcdpHfMNR22B7jJHxkwh7UUYAyKvIHRYIofD
PzHY1GFcK/eeS5QYq8CZnfnRZV5KYCHtFuK2luPjAIF9y3PPtqp5VC9A0OtcmgNW
KfiTceZ/Mxz3LsjgL3TkR/QpBzed4vkE4bUKIuH6GF1b/qBDh75aXBnb7Kgpgd4D
aXJj7IJSJENV60VNM0za79CeaK4Vqqru4RZQ4ktLZTPuWk104UM3RNVxyAcO1NOO
3db4IG0lWBe96sgjK3dTegojYjPnTWVCxDH0cEtzxRzEOzW+5l5vfY7BnyILRL2H
e7JqG1dx0uNEm8oNGtgc9qpIBybF5894Ivhr7wrxjnD8dqO8SZ2QknWnzBKa7ucX
6eQUjQOzzoNH0hJX3ZwU5tiYtm+MSwOYqFLuMapE6bKXh3BfPbUkaoUxPiRSHN6W
Y+29YAapdFb9JrtBBh5uIvzcZC9eT09JTvxUI1btKKg5BEJp8b3+sbvo7Ljad2I7
xx1fODo5wePVjVSkka0+2nNvbq5/usGp7o0IHiFjjavI8rkMZziohtGqMxdBlJLL
Xn7Hjok2DnvqPBgJxwhfoZEzf2jL/5AKwV2UsSti9YBH6h3ZOkR68JX0p/EJHB7v
w/ubpFiolbEGAY36p/j3tzSET7iB3T16tH3qdoYxVGATW+3pKJ7C8fGMQ5CJg0aR
UHwMHE/AhuTniRibGZiC0Y/HdFq+EIU7aOe1RIMzgh98yMBDSdPmrqYHIZXgUuqy
ZnBPPvjUqKbkr/cr2fraVRHeMlIlrnZ56HqowXKFCV/sosxo7Qenb/ZF2yxHz3du
3m9+hcBddOmppYahGGjb7dhJm81EBvulSejBN285kGZJ0w5vRisAYWJA19vr/Bqc
ahFTzfUrIQeUg6TKg14eyWimgtG39aPk+mCAeCd5mIX3VxrWwDlW4YdgZRQTZHxq
HUw0Y9tD+RDRfK2LD5CoOdiG2bn6pfNlBl5Sbou5Cvyc+A0WPGULQm4BydnXsFCK
3sYx16i/BZTgxwlul5AcJTzNcRLx4fgKZ125tmDpEWiq5656bqH8MzZ/9qgtmsdT
nEMbxOVWPS186d93SCQdRK87OWkDRaSf3gLdN9950wmUiXs8jNgy3kJ3YOhVZU5d
tNoXElUBMFv15ugUwFEUmN2+fK3LrlumrZxWRPxVdOjK+9LREcDsbbnTKpmpO+1s
3u/6fCarEUNLjMkY0MQpMMpB9hmUBtx1G1oTO600hWe+/hLIxJns36W0QDTzofWh
+E3dsl66b62mAETdx9K158fW/kZ4y6wIxVfHebs1jyy2XsweI8YmYAXRUPoU65F5
Z/bL7Le9xtJ+t9/2x5IkR55Ws7paAj+BoXLeXuoE3463/EI0ypT2dNtxDhMT+VXu
jfCzstXjkS67DhUeIwTsiK7goSUSqlFFx3tq7X5zwTrf2fPM1LVDZmeaRIr8hVSI
JBrCmErTr4c8nDHXqG5e0xU5DryQMZTMnKeAHK5kJK4s38GcQLxIcSlq9qWP8X/x
cAZjqTXBKhJMs4BOqon8i2/KvTpN+aOMTGTDHNDMNl+uC0MmBtFg0IrhoNkSSruW
jz7aXzPXH7qxvFGZ5ssEZOPq9rlT0w9QJKfGEbbcyj4fsP1mQgp+ctwZ95gr+XHl
llQg1cfVITNXbeC3sKxBHflI5sHRiBiyoulIJg6oBJg+/S2GiUHXXsIv/yySUhw3
b/QbxwrI4Ptn+dVwI0u9sZ3Rs/+YJ2tMN4xACPaFGImy2nwsF1wW+K2NyuyNsmYe
o/jfAK22C3FAdrSLjxHmh/9OkMEBeWTz3MyHXu9kHxkAwxhe32QzjTkQO0kB1l6X
3GSpNKLuLjJOPxM9nSiuNY2OTtoy1BToQnglRvilzv9f4+CkbAclM88/DaiENZWr
GGI549tBXyZyj116jbL8S5Lf0IrA7rKk+Ab+JPefabBnWElM7YJhL4iuJ90yDtkQ
twHZ4qoGbpXjFaPNZ7eYyQHKnknQGW/zaAFJSg0MLaSMAdF6+IbEImNwpMcgumYN
3/RzJHrP9VxK7+VTwfa/aD3/WNZj7xAQw7bb3IQRNwmNBCAMy+4RJm2HPkydx3h8
LvnYO3Uj2mduP3J9PM1SFe9wHA6FzyRq1HO7uKIrfEEwAtxdxTBOPpi5uQKCs1Sv
CILML1JBWUTsUcRIXOLt/kRtKra8g6rg+ZrR1Zp/Cf2OI0IjDp57F/Qm+u9uAZiG
QiWcK0en4O+GV+OwjuCvMr5oZAPxy2s5Ckkt2JWEBknErwmH2tGZMVEGNNnhDuL8
6WrrEZzYSdwa6UGtutFv95bkwhRmNLcCVbvnPSsZNMSYN68fwrZIYD+4ONTTSdsa
7HHynkdLpN2Vq/3TI3FJ/05KQ3dwt7o8+vH26jpl/owRQYm2elOhaxlVbavGpzjU
h619oKAhC74iIfX9pq/2ggIZ2Qr3/m7XShb5pUxdJScNoLCFEqZ5X+MNg/yuGm9Q
aIVelD+dMewiESeN0kYQapwjKV5wF1ZBzWTuPmm+Gr+tLhkTyvi3khu0q36Tee7j
Aohl1lDaHKdrSJ5ksNBmf1Mp5LjENKTutvvUgkhJYRaltuQJ2mjy9zgeqCWokh/l
sMMxA+RlBw0EcQ/TTNZ3NyK1K2Z9UdhJ207+zBeT34eePUemxObJljU6mDBhee1Q
VXZPtg3VB14MMezpPerBSMIivOknL9gVTSWelhL6lBe83tsGOHfzL4oW4yZ6S5qI
US81QKtgwfD01uQ4ap32c7GI21yGkuGI8UKCIHTez5X8kTQH0Hsz7LDRrFD42g9K
+38JRb5pI/zK4Xk8SSd25oTH07ikTFczx+brHSws9ciVK4mENN5IvOFVlr2Spo2y
tXy27ui4R+Ax8RfdfrvORzAV7Aomi/Pf4ZRMuQf/m+DHR59G8+aigAaJGHuxq97N
tt3MYqDM7FvpUZ3qhYYbVX+aMAoVy070vrROWauj4qM6/TfwCQD3fVgnI6tUIFkT
DxHRtDc6jrHxIX57N8en3FFnXnu6nzOEk/fLS9A9/NGAw7dBZGXGkXRXYRDh9M0m
0fFW7Zwocd0+mwhaz+zkJCoZ3UIUNOXIP7/kH77EwiKM3rN2/eDjoh31isAjP9WF
TBd4mkFi7xnbGpG9LjJ9Gzd6N6/2ehIRV+9uEbaGn4YHZaFJzzbHhnKaikyX1LYT
wGN3mEJnV48TEnJW9dnDxWP+LzbmV/BGtR4W18UCin8QVhIGfzYU/g/wFgmE4J/S
0imRBBDXsDBK/PlijVfjB9cwioOR1FEJFWQ2r84e5ORJrBfo0QiJ6yMuqTJ/ql6T
MeNpl00gXzyuUlCbtOn/n4nTtasi+M45rzVYHQ76a+XPSSSLe8h4T+B9lr5Pny2s
p4p3LzHIDuU8T8UiuPD2yajBRq+Z2jm2VwIgUBA2b56bu54EVprG56sVGdhuDCEh
VH9artwaCiSxIYJPkh3zGNiPiDyG3W9XFCa4FH6WplAWZ/O/gKBF67XsGmlkSBrr
31OmIIsbWrNgQooa2qmxo9pGaQ25RjhoUMGISfeKbkXVBCUCeM4hsl4CCN1E/JPU
S9s4WXnjvDrYy1wgNCX4tGmKPVa/SFqds+8nOMEn+Vkj840LFtUsxZa1pGCcYNje
awZ7TSHvUUI4web+jsM7La4cGqQQgCW9r43GektFPzyeMXHIS5l9Cl0uWGcP8v0E
iouSQCR7tVMh/Ul3pIEHq4HZz0UVTrH7KAqRxIdQXhuCRKq/UjXhFHFjocb5lU3u
WR2hmk7ZI2lphvEcfoJi9CF0xcCzhOotPC/g11QkXjR9pS8Vl9nxhreilb1e0NNr
7PFW9mbUA2WXs7VpE5qd1GlivSBRgf4FClTOtU/jzZCv/N9Tqp3JR3/qNKDOBUtU
nJdYPDlkPtHKDPd1eitgRn9TrmHGUejP4Y2KuB0I43kKtH/1PdeDRzDngxl+NOPc
dwdY2qPs7fvFOnaiJjcwPSJzwRM15xZKGBpVwE820Rn3Lnw0bscv126lzQu3KHKW
H2/Xj3oomb1AX7fiLvti80f3irdH+4q9PkUIAWarY/4t7Ca1MdTfua+ZvaHudJLD
Urff7MaWUeD7sfKJJ80FyyxJeFWkI+RS7VFLzzNybcEMkWjyC/jO6PgCyp52k3CA
QRSdR1pgbFZVWKJ0yO5UE+8PGFLkV0NXEyQIRdju7CjJPxrGm5rzXZf1dNSI9xFO
UD2kfvCg4D06YedvJZdKjHlHuFYQkHQ7qaO6Jp8ImE8MY53lGpVTY3IOK1WGzmkp
S/dcvQMfHFPzE2tuI5JRQyHONtpFl2nDtwpq3dTZEIWhRnhzth6K340cz2ZD5arE
MmNCjH8zRX9Sz7OTKwYC/GVHt2yQGa02mczMo8jCB0tgAuRDqp5G0OLbphhLPYxa
RbLbKFnZSlhTqXGVaSXgXeNcqqw3pph2rmdezGGSdEh3NSXfpZ6bcojJPaI0lMW3
bm3Obaah5vSKM5VkIjRB+znAmLq0m1pN8tQBdZGEw4Fp1Uac9QlBOc2K3nocEmOp
w9imaWwEoRqnEKQ07gRhYvmrmpNCoTpinbe0mOSODJC043OO2VAhxsFj6Zp2xBvZ
u18bIYAFm7WUksuGOB0riS+14c+x/u7zh5oB226vUR5p2wXAIjCMVps06xjtrCoM
987vVg2akqvj6vPeIyD9LipBmGO6P0QTjQOaG9qRKmi+70tIyeTvzIlMKEJemQ17
GWxIPWcL7JCvWQckzsgL9rj0SPx8hNXHc2Yt3wTn3wU3Kk2Fcli6arbh0PENuSYr
MYcz4KRmDvMYrSmTfApLC0CpVq/4ZJ1hTVIno9QVjuHt+jRDbKbZ825fQhguTwVo
Y0efcZNZWC6L4IeO80uye5rqc1MuMZdz4JFHvg/jqcwnQid4POdbvLN/0l5nhs7f
xW42ZIX+ZyCng1FdXkaHgD4poTy5k/O0iBTh5EB58KvMJgG2sNnMM/Ahvz5tODhy
zmKHpGe+n6gh262IpcDHCTcg48tsQSpSEBSATbq6fcblmTbut1AN0sJfaggMnat1
ikdNoIJbeLLmoaWCjIpmO2YX+zGmm7zuKVJ85SFupYwe3q2fSt7Y/ez5kyvrRqxY
IwpnxalPzabxP13Avp12NlG9LPNi/biMNCJEQiAxO8SRGvojMR14fWobSrdLZU+8
vPnmFyv6b0T0XAPbEH5dwn2z2BVKlNmqJbzBi7IndhAr3kTPlS/a9bDFNz61ynm8
+VQXv0So56+Mm7uevuWptEbgnjxJwVH2Qad+/ABhzd3AYacQ/HhgwQ7A+mUqTPGa
D73WRbnc9AdxVqh0duqqVCERfFhNV/KIILbz54C3UVaQLE53+ckPshiZpWlbBq9C
7sMharnbL9KdYlP1YV4omxwyiNyZWvhbxKkdUv7j8tp2k7EWQtFfGZ0WUiiqPuy+
EHOBT0C1dmUb37qp4EhnNFx5Ei2gfKMPHCuU9cjwbNuZfDrZQ2/XYpPKvKIOL/1D
W0axMwZuMXEUEUBGyguWIT/4YvhdWqYQ87AqlW9tDdzkF9bbVqW15v5w/EqOxZt9
rmjsrk/bdPWgbW65erED4BzKU7RIrH0IF8eAODrsbOn7H+dVS/QtyepghYQaQwnZ
kW0zolTn1DfNIUXyxisKJOnF8xJyVA6TO2ZtCNp2DqJY9PX0MlCNwCvazGr9yOB/
46PS79hcqTK0SFK2L7aiRW4kRGUbCyIO6GAA76B4pwKVa6GDGH6X1VruPD74ieOc
pxpwIdKbrphsI/4REkkZ+jt1v1CBpnOpCrghcz1WgJL8Vpj//fYqLApJrMEdyu7C
91fHq3/YJxCYSXzLhjl2xRLFIPby1rTLEzNMCu0o2gRa+XRFENVL6IdDiP74Fc0h
kGP9rPFDA9qxaAdN+k1Lv0Vjk6YXzBtauSdQg4Nj/EjQa9xQscXBRg2f2Yb3P+US
5usEvYKhqSedPRNx6ABq6u/vfH3cJflVV7fHWmjtEhCTMuI/dxNq8Ta1kSSenH6o
83FJd+Df/4B1KDyrC1BZIG0pA3uyJWfF/5v1SrhUQViun6PJ13HLqlg1KbffmpRe
TNX6EmSGtFC2kZHPR7hW+jYDTLnfJBaaKkDiR0wRfnBePgPMugYMzchfEco+rEOo
BkdpW8reNiYkcWMxVA6OFmk0QTmpf/VULrUBZuuOmhss4YorErKyuVV2rr9S0bQC
FXoZDg+PF/A7xHV0aBnF1JIjr6tUs4Lai0BvuqAOVDvRfkQj5KPwd1CRRXHfBERA
B1qGh5D/y7jqSeYjGC2ugVUeg1CuCmuXcu6BxViL1cvEtwYe1MtAh4qfB9U82Sqe
O/X0FxLIfVd5etT0Zq8VR0TMV/hIlrLSf7pSRM+yPGSDmnq1YtD85fTtOTXUiIw9
02WvVSUi6WuCIxk8VAFVZABt0X01ixuANxV5N0nx0RT/4pYxIRGxccCg1i31UUN5
/DqBYuv6dYVuLPBzY+mH7lAT4H+zRDo9D3THrz8TzXWn1dvkhm5l81x9GEqSHeIh
VGVs9bCNjwvHH8URE3/wvCAEHxlG8NWn8y+e3vVanoD3Uoli6Py1xBDsbZTzELBD
R1BHAI9t4sOJCVrKQaDrAtUda+N3iLO7DzbUG2HFxAtfPjCWrw1n70Wa0IzZ/HZK
5lVC6oEraCbhecn095twk5QMXfg6HGDRkeDTZPAj7hD7KHJjlkZTrlY+4SqIKoqo
JRNQ+bkWNMv8lytlp0XkdrsHZF4IfHyUEY/q1vONtR8IpUv2wmxYh++cX3/zT5aX
NNDls7zWUrZXR4c/6n/zbfItIfEAALd3IJ9kGSokKHOMJ7M/FwGvP6BLbpcxJERW
0WSQuoboON5gvwfdt2YLkLj8UQZ2WM6/dkw3j6AxQ86Id2K1xTUNrQbY1GlV/ha7
YtW5+YLjCy8GJElcpnWLlv5sqBuXi1QhiSRlO1ykO5P5Xjx3i3FbqzoVBVmIXvBy
2AiHHpxvmh7pTUf1JskSO1WQ6JuUfWj0ysYvx3X2lAJZbyBE+B4H00w6eZixJAHy
8N3lA1AgJVzSjwvM2Gnx4/rPlqpt+dvFxfxuZfFXxYDVfj8sWB2CQeZtoluwl19o
iVlAVIsxmF9ZMBFUp2cBZDDeCIdVkCYyV1Uw1EPnIjN/IQwP7vxCnvIXC/tGgpvC
r/uDdawAmlvk4Qg3P4wrwYQhBmtiKhy7kxac302079dxoVkfEWTEbLQAs5IEoeUo
YGIE8wDhoUHyZmyX0vETSj5SeJKW57G4Edll1f2hXFOz/L34OGZKAMGuTSI510ZR
+qADtnmSGldInvV4j5zUin3MSKuvGfM6+gbPpUTw7HF0JUwS1YTitd/VBoAl47yf
wY68z4zAHxhh9AZNkdI9pQIaxJFaYC5ucP8kLXqYRZqX3NZwPPsH51I1YnMKSy8d
EHOUrYwyOq4y30Px9eD4VpLCl8u9mpzQbAS0wbSKjBhHJElHZoIQl7SudzSldgQe
njnQKVL4sz2EAOwd5HqqEm9Y/Tx9R32b63ng33V8AaCH4QR5lzzKqs99gbj8nnpc
XgR/lm2hVqvcWnZh4+fUrCHzDw3NwsEXYM3aSO3gMDuE4csD6ZDCgDufaCo0N5+B
zH0Inp9TD+5OjdeLDkDs+u2KR4bRRYgCyKkWBkk/jDz+aYE4i9Fmj48D9RV0eHCl
ZRJmDf7S8PEmYiT0YuyQj0iMylwWkdHZriqNm0YVzu2ZsfzeKIMjEgmrCrWi/CfD
W9tSkei9+LlI6UuKSIeSzeM9d8Bg6nUAeONgkk0GQUk8EBzp7Gr93NgYcHrkfJli
jrUkk5HHS3DzguQ0fzNAzA3pfgbCzmDifjLyR4q2qjt6j9BI1MQi7iWsm4GAbFZM
PuNzy0QBH/o5Pe6cx1W7Ovxw/+dHvp382NJG2/hlkXPO4+lkJ2YGPI04XO51sgXV
aQ1HAdUr9KPw+1EOrnmYjZge7/UrNPMxxNW7006HYb+wRNPiDuImt12VbAT/IKzO
05rdCOEo8ThEg7YtT6RymGPIlStkutyPCYthjsxU2sD/oRy5NSIMdSJuv+d9RAji
Ocv1HiLKc4NkckaoUtLq+tfhBbp6YNoF+V7Du6vSiso212RFnTwioWRVwrcLLkVj
sLqj65XI2rcEGaSgg3G8AV6E1jvMT663/wNdsmGek/HSRPLCNRgN7I0jiLsOV1ml
+dXsg0iOCM/tMXzJqWsoPh9R5KlBycqLayZuN64IIU0goPQWAq/b9KRxuCjONTZ5
6x4qYlfCym5T4VooGZPjXhAaryQuOqv2C6SDOYE79LFYbQOj1u2JDaPYrKuPaLP5
6a9xxnhzh28F5lxViRQN9o2Trh4GRTbhBuALclAFz4B/pjgozMHo3jHmUF+SMeyx
doL1cx/K6Uv6X+g9Mamu5L3hcaZYmL6Ria8Z1X++68AQYfAz5ubbT0N1UrAlxUJG
npEo8lFYg5m/ZOoxRJXXvU6dK+uxzdh9oyo6wEpl5Xhua2sRJH/fK9mUEI33Xxel
PeOjx9v0OHbtCrsxvyj/lpNuYElkr9ZWc6MmuV7ZI7eBTgAWrz0iG6E2FRIhu8Rx
NJ8aDNAu0AvaUcYLqpSAVXsc/fyHet2Kvwqrhi4LMB+Rv31p4VZ4oU5gAlC3leHV
DiPO5NnrzCc2me2juNUiA+mhMGXEHdd8YE+KtkaMggXCbtS0Igx6T7kRIaNgrq5z
STKy0hVWX5dlChdi1NYqjtsx0hYqWZr0ofmjsde4TyahFHUYYd72mwTq59Zj4aE7
3Q2d9P8wx60SY5tIrlewdGl3pW7h69IbxUkgVfKdDoF17GE3XxY1FnTfTxAcK7Eg
iBrPW6G+AzmOY8Zelnm0NA51obZSkkpZjdvQ/lItB/NdjNEo6V0i5+rbAfHDDrOu
LKC3ioKiFWlsZkmooDgxDCexEJqADim9jh3RWRbBseF1m5eecHZPL4Mdn/6+4YBC
M9xSlnBE7yxLknw0NwbQbdqy+obv56jbA2ymCvhf1cHmEbAEYF8Oq9Agfq3ao700
vkrenWcyWlJbm1ds/62rz84VY+sfTZNbTIX69SdG0FnWMk7TZuGXtFbMPTxKbhWi
T2wvxYCjXiW6HTWYithvia1w70vaX2/j3OgldFGPX4moWfXkQg6UEDGmE1flbdey
1uvvcSuQ7zOmRI9VDzeJkYIyZup72qif63Q0BA2ptxwOhTGtWKUsbZx4kpQ/fL6+
OjrOO8yrvpxHcD1w3lnHj/zIy/urOGOC2H2F2UbtUcHNonnzBQni8eh7/nv7PG3W
f5sRlV+/cOILA6wLcBDtpfYyB1G9jPIzLjtaqUqqVYLKE+7HSWXZcOEF3lYtj5Bs
57bMGmYq1+ZKqg4t/EK3XWBuRDb35S4bmhQV/Nx3zNdsvchYSupRm0DqL+NpHvkD
z6MwD0bw16kAPM5L/mqspObIPBbJaZaP6K1Bdht48GtKmWnL7UApUVqPM51pIRmA
rGj2nvy9jGTaXmGjuFrbv91M3MgUHyzoqLXgDPyQFizhMfS3UtR/8Ay7rvgBXgqE
XBBlx5l1ayfjnQzsEbba5BIufeJ93UCjUvVt2LGkUYxHRFJwZQswUa6fAFv8MM7Q
r9zMw1hx1jq9epEx9zpAVRW6RZixzrRjfMUSR5pKqbPOuNWcY5S53ujUsQsNO/9L
bOYTbEHZ6Igwzq7wLuR+GvsxqnYQc8nYSmFIxlzwIsCSEvV3JYdJEf0qJXPGHbAd
qIXexKKfAUeR8Ocx5wy+BKFj2tt5OhTqQ1WEInz2gwqYlKTjBBAFeGVi4EARRXBX
7GxLA8Y0Ewa9TPPdea17vfZSS2lohtOn8AIzKQXeEhAgPM30grcsgoz6YXPpTASX
8LhEIp1tgeEvVuloKFO9g0NdaLPT3B/7TawzOlQ8VLyfbzQwE3xsBnzg7IBeLCpW
FMgxE3ASh1phkCQ7lPaaCn339VoEhMLhEpYDh1RGcbHz+nF69+t2BFgfgwSbDgRz
A92tseAQFwWH3Z+ms8X+BPiAKPRg11w5mOQVA+e/EsIgGqzSzBBaGM7g1yQo2SJi
JMmreibsISQS+BtAfcNQoQ2j9CIah5Yjbhz1hjDbrmyTcSj4AK9/q1mMshzvNPzm
soj1fffHXjA8NFw5oBVY4sVy5JaVi5U7/PFSNASGehPxvISAuwqsxxzo3H0MwJy4
iMizQUUzzkpJ+LjbXMmtZw0PJ10vHIBA+fv5IO0iJPro7DaYIWpeYAc+j6QHqQQo
9PaQX1JgnpYIhiSj2HkWMyJKiSW12IZwxl9X6yflz1ddWTlHyS+a7LhMkfkFHnd3
N643lF9gHvxHH13EiWRWA0o5SpeJC4wict7mN04gA3Akwvtf/GCwmOxWaRnSXI+G
F90Yli6PgP2WK2XEGl2MNLODodrpfDlBIkMvl0uplYMFnWLNfzBNkasMbhwA++O8
2mHhJ+YGOkdWRWR+6FvfH18HkwYIKHt2+p4mQMYFvhO0thTDRgkwxnz2DUcuYRq8
FL9XFSZUkNWKipl8DXNfukzS0Ry8ej3ohDDlDo4urbj6PxaTVGjXktmi1rjewLJj
cLJZvltaDwKzBv0nW6Ed3xYrL8gOD6AvX5BQ5oac8BV9cF6yqtg7CiC36lypZKZT
rauBrja++jnTNxx6MScvPJh06M228hxhK7f6chaf/sxqSnDEvOJCjp9hDoutqXlr
FxWSUimDLZk4IooC0p0jxjZpkrwSpbOaarzCped3nvCn9uC+1P/H1RoKQbJ1JQsB
jaJi4hbTTcrU06hpFXlicAJlsO4fmXPy/OBEKr8J81+rVIlfVDqOpEaZtPqJ87qM
gWvRrXwIwS0NgL5WPgm9eXH3F4ZtYHrUddeuVBEmzSD+sbtu+A1QBEWFOwRdnU3W
9uol6EyQ0atqAsGcw07K7G+lpM8vOf/XDfTkojM1VspdakxmIrGVTitZ2uEpSpTl
cdYD7ot6UPCJq0WW9muyaNTQVL+efKIjeznSP1dLSkprFvpChpHx0F3ZFF4tJjRb
Io9rAmD2ttUkmtmqexfw7y/nRbi9ECNtC3PwK2N18mmfYdEtLIuiiRr+tT4TrYle
tBrYtp0hFlpaJaNhF7TFabTYEHAqCuTJTWE1e5Oo2S4ua0ONfeFQEEFzUOvXwl7+
KMIaT0jEmu8h7MouZ694oLTsJ7Wd9i6vPgAhunEPQhUH5kXtwiit+/8wL5faFS7t
Kgmu6gzQrDpEqAkx0DS+O2rZ1YZR1U/v48SGyc/1iJ17hMZipyYjNs7FKCrLj5G+
bMmMU6ytggiG3t27tRyM1jgcAxMF8EIFQp13IBVcXYVf5IWkxlIbUVtvb/S+nQyG
jTxMdwtHNx3kLZkFzMVARwzMTx5ITxUl+v0atoSJ7KEdZcdyXSex+pT1Wo5DIt6z
z2jIGr6jRTjShsvNPUkWl8CxCftADkRPmLRICLx2SvkguhkoXTvzCMdmzLEU6k2k
UIp1MI7j72OvYO3HF7y4EYIyFbT2/SpXYySKq8vgzXJ40yOpepHL35u9GUWjitO0
erkArVUQLvz2CKjqaDSLtz+lbmzg25ELIR6b+lUj/Ub8GYMYVQbSiHe+7XaWHPPA
Yhyh6kfBkmKRngsCQDasGoBhsuBe+2O/WZJF7H/ACZvPWTtWlEu43yK3tcBiYrsF
ZJ4BuuR7nzq/JWOBvRAlvVPcTXXq3s+Xzl1Ctlt5CL4M0e/0iwU8ebAVfcNGU+pQ
TUA6BfcX5dXlOCiiDB3kLQHvDTDBy58eisjQPIqZhGoGM7iRrAU5G8KBBEy02M8f
bLuNbE3yCe+DycPyjsfluNjUgkZYn+K2fXo3YVfAIwUaJg3qrgNg7rj5JgcvZ6xz
AQ6+RxvR7S+r5W3EbOPboR/WjbjQIs/AW9UvKnJaeIyqWVRqtLiJE0NMYBxzBFtp
OdTk0kkw5gVYvDgQq+QWEo8KVnePqYqAOZ3BkxfMdza6VCq4rwcKPHFg+xcQxMAN
FRALipJldqGSOk28GCmxp5mGOh+hm2ldSWCuH/3hMnASuM9t/rI2OyU9nCxy1Wiz
FLuA3pUTkyFNPr64NEc2b8A6fzKvyyoGnQhUlRubQ9Jzy0JKs0zuGb7PGmuQcu3f
28XCxiTqdCK802tR+tfmQng/m9mKPwQRWJvro5L9scN85GJVbeZFkHIKFml7reUE
Ql9FSwzCkxRWkD/UlKWXWgsBk1CvdpttfEft6apKCQ7cqXbekv+qVf4w/hJf1/4C
3NWuDxWXZLkuNQvvQkKPPppbL81Lsn9QG2FiTpVhw3MnCUhNLgr8g7McSfyWf1uA
XaPwoloEWdPX3DbvcrZHz2J5Sx45zM5fGcpaVk/yGvxEFvVfArl+wNvVedIlzAvL
L1T4QM4WLHpwVLDVOr6U1LWzto1DDcXwtI46q3U4LafYhBXarodlTGOelEjrqXoO
KKXUfP5ee0LXL0CvsTo3KJVGs8rr2VTd6jocZ0FPI0GGUjBaZLcuBxoz8xBGJQJh
7LeEaWKXBKu+GjSKevHovP087jeTQjJpBvtGY8eWLuEu6nm5tr4rGgVTY+UIH1of
aSb5md3JlNFl0usCnednctUbLr1WKRHrhW7LelR00TwATOm9hiicaZRZK1bHaQHI
jc4xe0ygZAyORl+L1Nke97moY7RqaEuXq0kw7EURkflYFnvFWh2qtL8mAeX82J+T
6ww4sPeKKT2oCoAS704dNskgCsz2iS77reWcx59MvL5+CTUPbS0Q+0KA6kukGRyi
/vWpfRsn/sl1gMP1eV9Lxdpc9TAkd4THbRkAj8SCLOdn91vmBm4dBb2QhKBQ3YLQ
sdCXgZDtX3rCWp0D5Is6GX/hW3kW7KPV4ZgugqGBbgNA8jXwWkJkKAgoxgbYvx7P
FFicssLgvFajgHGFhBg150nZUGnHEPeRaLVPlonyir92I4D9t+8RLR7wFpdX9L7v
lEFXLys0u7eTxFBjhaMkPrA76JkoM4X02muzN5CkYBoREuqjsOh2aSKq+OTeCRNb
ObyvnHsZ/iLXyKv8/A2WdAHlSkGnBQzSaU5jSk4iW3TRmMIfF6rIl3VsPBWs2es7
PNwd40KWmghuwGZtvTzw//SnINIrPVIKActIW/mdons1fYU3PgffspUrsWe57+K6
OQ1gqxBikOkwx7acgkkYaFo0gwnwc6AYUHSAkcl/5gPHwTsKMVAT0VUQosDG79ml
ULNekrIHcgZRprblwhzqEIFPEazq9MZeAO+Ni31ieHK3CCtH0HAuABCUyjkyICEE
VPAlywbCX9YZWu/1h/1Xa4DlZq+0UN0UGCrmoWkStqAowyP6D+AA6YjTrON6ATqO
A1fyg7Z4rD5GAGmHI66FceATwT0jlrWyZMxh5nIc8eUaXvZ4sobMwOPsQ5A1JhqU
5twZgn+1YBY/UvIsVVHI0e+7OiPykRqQdWGm/xl2aSjvbVLxgUZGtViMfFRxcLaw
ALypxLHDAgRPYlKUcfXksqUbz9cq7rHaLMk5jMqtp6Lj2x23vnLIxVsG+HZj5adg
BDfjXmtwcAngKfT5iWhyGlaJ3+iRntNKUN0pTtIyjiutu2l2jjWWz/Cvmlvmw88L
7si5wEw9XNpeLF3YNKdpHl2TvSOT87fHsKvD6wCLwjzMFxlgpHIxIjkz+3+z1puj
Z/sVmTgRdjaTZfPptXjfqpCRKHhoi80ojznnnNWNyC+NV3YAzoCkEteC6gg8IDpf
buDkeReyFXLhCatmhNV0GaH6XknImat6wDCaPuMwe7XAcaXuwU48S1hK23EkJH1m
pCiAGbX3eD1maZXOOeabdD+V8jzvauC0Nl3sH+VjlXz6EZKc6/vk0GEUiyO+goaN
QdDgdcxJ5RJLwn3Vj6/Fut4UQqVIZb/GiADuhQB5JxUrW4jHNcWGYuGji5ntf5gF
wyfeQb/HGiQv1wobw/wXSptCheF3Y9GlzDgGuAc8LJSHvFVJnFIgbfdzm3wH5z8A
2aJOkqhn4cV1C0a+WJNgv5G5IuGX1CQXAAnbFWfMZ3mbPXYhye8avWuPiU448gZj
Cj27g8p5TY+v/uB6ge6Zbx9h7zy0zGAbr3fhqOWaUlWVL97e1lewczU1H74rtlSm
r/OpmP0ffM9mIr59e8l3abLbLhJ2KKEgDIUd3OYUWLbLrUCL8BFBfvs0yp2J4Vhy
4XmkOKn28yzcSP9UNehHzb/whUyhBGJORHvV5vZ80b1IlusKCVR5PybgQMdtbQIh
3EZ502SYBVvCp9owKuPukC95P4NAXjeWgVPWpPuHp+7gLBPxTrC9oYOVc1iMEX28
nFr4hcf5AHYKxRk9X+Bmpua+iYmpgdN8ar3cFrhdtj58Uwb/zrLYWC3QjT9K3Xht
dwYVoLPeR2vSjKf2/r83HXQVuUXXhLnY6fybqOCPLhLRahMRZBfvHyzLxqi2V2hm
/aNd7FLzkQuYPIsX7gTgXjk01fV4AQ5vKxkqehKOjwjfqpGfYo/zdDNfhyw1PX2W
1TiCnTx/JsrbwtFM4SmmrmYiDMayi7GyD+ZR8zW929Yj6tc/Cs+m2InxprPVdAPF
nbr61Nuy6jTG9IN4ynUU4zXe7Q5zh/R+nuGbEuzHkxrnWGslPkzYhVrxZhuLJ/Q8
3Nf2Dcdg4yyMHc46vdM89DFYYsm9/ZEbzTVZHD1SgE8G8SjduDdPeQhKkQrwTy1x
5jk2LS9JMy8o8qJn3K0JuEz64iHNFdp4+cpqMaANHrWsrhTDz9Gjzrs07w8LIPqT
kpFABdWtdn0+AXXe+qjjE/MaaHHz2cWBFRHw/nsR0owe+K3LEjmp4qT499kmadyT
a8KnWU5lPH7k2lwKLbsUWMowtF8SXz1faiOc3Y2Qnub/uPzrGrDFtuBetm8p0e+V
RzaoPwXmaHIxr0k3KjtW/3Vc9KidkWuDAEt5v4+sdATzpwEJZcejHzu9X0/T0wgY
jCV3LUD3nQv6XMQHXdLNrTYPtgi2XXP43fqWG+LcEiTMMreWeX4gercowNXYQ2Ft
2+uAcNTb5fMjsFHz3jIscOx4aeGZi/bqotPzD/MjAM228qVkGCVQJpSKZCsj3GDk
6kER4dHu7wS3LcrPND5ZSrRIgjk4xIfuVamEBUsRrsBjYSOamQHJMWgpmjMjGZlM
19QGkITjHz3bKaBZFU0DRKbu/wk0rPfq7A5JP29LihyeG6GX0TgSKqNHYYeyWesK
hrI5zrCpKBaEil65ZVQzgbuyDhJdRgame0y7hyVnSb0ZhfI03TmMdSdDvD379f+n
RKTM4vIgglIyU/8nDY3nfqatJrdziSJMBBUaOH0oqN4TYGtVkoDrru4CmXnrSOSg
ivtac/mJ6JVDvyW5ZT7Brha5GxUqabk/M6wCct5ls2pm3Ht6zWPEr9QDRyIoD155
YDyrtUN56OzUM2HI+Aql4GUFsxzu2zdLeyXDZosfbUvpoNhypnDlFKvNTd96qGdG
wSmAW77KtObm4tvoGW6YIHqgLbRtbHZ2rCBQdEiaMglHCpLsaMeB0Ddgs0o4OYTu
9WwCDSNsFZfEaM7zIpTKhVAdnMoqHnJ7PF44GR9qg+gFdpf+ju8zcUIg5GgYFooO
eXhwKUTNdGd0/xVRSvuePeGBxSEotObdeF3W3X8y+fBqtimCFXhleNP675SAdcv1
855HYxqZSTtNBBSim195ejqewRv0BlxjJPW2703bygrYNyOierhEpZyApaMl6dyn
Yg7VWd78DAE305o6TtrSD7mwZtglElRikYeprF5a0cXEGEWCVVqaejW4PhTAKgXW
ebZNnz10zGb5auxZPO/uWKXbP/KwlVfmTdsKNheiInmQcwgjaH/UO0+nph5et+FZ
yaCYmxCC1PinVmCFI/nFTw8PWrvCAF1lJpClW4+9xTOPvIcBA/hjTEXsV0ldBTtc
dk2DH6/7OubhmkDeO7VEmgNk7u5cBzT+ATVy44hUK5f+IeKhnbnbl6UO8T2dL+T8
WlO6nMYAZaldRqekiz15o7Lt/eQcxsPcMUSWXwjn+GvtklfH0FfOe7xh0zMvNKq8
U4O1X5rsGcBeZZOoBuaMAwUSLIg2xvI/1KMH9HewOTacn23RAW/WhSJkQk7Jy8bj
qRcIOqe8ZB4O01bSBmNPYbGVKQxzL/oyeN4uJl7Xo74HyLA5nqpCl9fdeRJU3sh5
nstcHJ2lSTghrtNhYp1T5caa9ZqL1ah7nLO7yPO0CkySnVqcqb/rgiUWGFVqOhjn
k91l/NbTLVTihX5CsYDW91GzJSGHyhzNBgLybqum0t3/CnKFleC3ucrzcYY2V5wY
xqjzGmHU3Asm6G89+y33BRR7FamN7tzDSq+U/z/xUIZ0kOB2hV3o2JnYiH3DLxIP
mOXv5ixIJSSIoitBQPMYaervcVEXrnfG7ujH/hEPrEQU4orclsgfJENBQQI3+P4+
hwA9oGuF19BJZThQrzLHg/YDtlGU4xsSHGd0NThauBe5vacDaK2ScEaEa6ZdQA9E
ZiAJp8EhHkByVUaVstjDq6/9xMcxCOXeA4Wq4WA/4kDMXVf+CiLyp2OMgO6on2mf
Kaoc40OLQeact/HgmCIMjSpvRCdfb5UuQvbDQIYv2Tuu2oT41ZjrYFxFHKpFsoui
sc/hf3McnO6Roljo+2y6+2XUbIrfk1X2LO3GzLK06rPQuSlZj8bT60n8oVIRqfe1
stI975eIKjCpeN8jC3+HLjxMQGfBgy6AzhxxA0J/bVf0jvxyAWrgfrYG2TPYgr0V
QRAU/pizyhLysx4oWcVHT9oMfIdCo9/8lXrB8DxZjCrFzGB+7BPvGjvys85LPWZ9
+P4SCX2Xmy5GGHV/hPn50kuiitKnbQINE+c1DBcZsBvQJ7Ql2jfeAM9uvogoihMD
7NIbnqPbaNiTyqoXHLrxHQe18GrI/1HpdpJd+y79PTDphCaB0xTGdlMipA2WQLs9
jIlsnOS2tP9ZcN10pC111DYMtMId/m0cOP8wua8omjMKu0GJlrd1WAoiDb2j6mHd
AFfpke6Xm8C9HiEO1GIfoEFSBUyh/GDPnAFZ4uZZ3ncpITgdmMT3OGNka2JxqnTy
rW+LIBXQ+Gq+N/w4VyJemJXXUXKMCZbLkLHrSeR5m7zGtk0NnVCJLb7IrY6iglcf
KZoybCFCW6Td2si+06UJFaQ5tA83TZussAuRBCOD1ozDuZEDdKJjv8xIjrXrl0Zz
6hh62B5Grbp4jlB0fsw9z0IGOvK3hQywL83M11RknTH9sXh5PjpsjhcpSM3v2Uk4
DwtPdFZdLJWDxZoihHYX5xSIAQEuC9aHwJd09gQkXI15Q3kszW8kiiRgv7XrnHZh
fP60UqCEpiUkBGGoW4+RCoC92iFi7CIg3n85IyrgM69jyqDxK12JH1WZEYx5kELe
53PcJrvbMasdxS1Sh5XoNkgbDeYQ+DnfMou1xuuX3wimH9LKYT6SNWC6oQVR+vnH
KIBOUeLieorznlsZ6TOHQ9GJvJy9SijYqUsK7Y5mkZqml66fV87aqPK/m+QcSSbZ
mFlf5g8OlmBOLEeXlfEAYdZ0ba92pYBwCvECGohY2I1fMKm6YcZ75dK2lO0Df5hp
1mOMF0sEWfKZntXnLL7ibnt/pv4Zq15I6Q/99NbseOjLc6o6yudpMstTb4LfA1ft
aV5nMg90beH4X6L/I/0ofNA+RWh8jMCGCel0PoNkiYb/ylClxFspWzrSnwmcNngM
e9up1/TIuht6IhbyMegODY+Q1yX8VQc7pln86ghHMvVt9zgXcWAa39azwC3v78kr
rBgRoRt2jtQwWB/WX030wmSzOR9bMBrMBfbqvtGcwJswh18QoIAWfDmDHqZi2jwX
GcpN2eCOytQY4QmLS0qr5XK06ooD4+60eq7oj9wln8Ncb3bBD/yvnLgNmWajJPcF
hLlgZTFOFdv2ZCOUtRuzz3OixnwbL9WQYmkmhBe71wAvQDucwCKkZ57mEeh6uZ0l
EibPTHPP3qzRRR5fGEKIoW1NBgT/lDhrkp4UQipk9fra7zj7YB4IGq0X6tSLDcs6
Nau5fSTJIR95uhXf+lvlFon+oDi5hfto8qXBukM9UwG/fZRprH44i9xmjhmolQLW
QrjliVi29xAlvsld2GcOlKUlHM4xF3wHbrn68QgjXsVgf1U6Iz0Ke9t3KamKDJSS
Tw21AfAFxBw5h5Hk3RqyASpFiNlgs9GOYsCxmq6WfeaVAeHT/I5OSE4z1kdXApSa
QfljFEv3/hEmAooOcyex6joigZqlFQvy1GGH83GZE83MZLxLlvSUQIS1HpIlSK+V
AywvArunN8NECki6VBEbOg5Gj771Ya6AcoPUnve4z3deMoVm7J/B/ffCyDAx+qhl
IFCqxBUAfzzxP32N9i0cPlJSEiY2Fl+ALNFGkn85oqsD7SuxDNJOICtwsErXHLdY
j4c8yy3QRA6/ZDjNbcchLJBhEtot0d2bUKyihcMsBEGe6cYoAE+wOpstB54k7KcY
nXEdjpZ5kXB8HqpBqIlOXjJzZiCk4Gmg5LL/jGqjUlo6f2TF2UVxSCYq7US+FIBf
PLPFcxM8urmkGn5ULhL9hnWZfiD4mRvJOPoQthr61z56TsilABMo4rWbH/o//oq0
sk68y/2P7CEixnhp0njd291uU0bjk4a29NJd+ay98WxAo8nbX4yMVTfUwKFBE9Wv
OYBOgxyfnRQqqrEHvJ8YKv45DmhiPHwV7EfyMVePx95j9nbkNhEgbWDfIOj0A3uw
ueUiV6tuMWMN0s6AcWIMZX2s8RxbdB2H3+aOcHZ4HaIK2jcAAfJz30zEKrmuFPmq
7V4TYaIekQpDt5YU3KbDqqqy0f3CB3d1IRTE0A9g+8NsIb0O53aBB0T/7/8uzSZy
a5ek/IcNVyATRBNxW7Tuwxec1Es8mBjUM9X3fFxwOgI+tQ5ffmlPo/l+QrnvOAFV
25YKWCCxknnexIMp+e632nrqEeT5IJxJOnz56iyuh9IAOGPh2XaKSq7WuoWHEa4S
O1LkDywRtEWYZalF7OGJShygnPq+fDZcsex3plCU0VUYtmugIe7n5/Ls1C8ddiRh
h5a0ujB+CpGBPe6o6GwZvmlzDa49wqPxv9UQO296UECILk0pkaTh7ZQXiQbv+olY
FzC9CUVcMrmQBp/D0E0WSS/bYUCqsPC7ZPcyebCXLJ36Gca3S8f5i8AZhlwjnweX
qPMeVAPINLOctKB86asIEqP26GjzdpY7BNZtlSbKUDpk6yxvD3mP5XT1slMfB4Ju
En4SUmhwnxmqGkkNeIeUuB0F2VTDN3XAaRjvBES1ovk9Ton93sTwim/bUIH7qkVb
N3Olr7HnIfbTpfwUhGkphFCY16aqYKMnpcossgVofGkbtqXTraVZFWcN8AZn+a1X
hftRdS3JB3tS6OSJEy+GYXxQFm9nVk8zuYlZmNK3fsJS31cX0MIBAxUxZAs4XK8a
T2O3hF81wVVEx4jqfrCxrTvhdFdvHWB4lUAAmmu5y4Ci7QrF//bcrDHY8QL05gmb
id6EhUyd8A7277Tor5ma2CKv+MjtodBeNf9U44VH7j5C4XV/B4JAmOCaS1hjq3on
daIjw4XLkEfWJQ3P8WaJoMkjPYgGh7l5tuBLA2OM0H35EmmFBjb4xyJhbD46va7C
cVb8TxKUk63qXJE2IdYfqJB9DMK3WSIPMhWoK7DEwnW+HbwXub8qRLaNbF2q8Sp6
MSWkvNgzNViTDVd+TJuzZ/mwO8lWFkZTHRqO2WqQWQwaMXPLHz+Ty7d88szEdzSn
pcxiwcoSSA8J6o+CQzdz2m+ADcQWRfofawqjHLfClHXrOu5W9cwz7kG1OyNK0baM
xmhqDQZUw8k60jE0LFLjJVz36BTbnX16phO9RJ+A4RRAW9avQ1VtLhNuPBEnxTsY
o+nARVoIIxXhd6OSyRPkhXhaUAi+p9dvAFLJRahZFAAk1Om75w/eLTBcADba0Ted
Gx1rz+K3ZWweBDlvjvUBV/s8TCy6D1SGJ7HxhfYGnFAiVZ2DyCUoaRWUDUOmU/0Q
UT9BF5diVo8LKBsVhIszG4KyM2A1NvRSB+kZb0J9VAFvf/3fqDvY8oEjh7v7yZY6
L8bbwmhsyB9mEBYhhyEx9KBBdf5jwZ1Y30pz6QFHNdyg74gxMz/bABos/sZUjMAP
fh9wwZkMa9T/YpuQFIBPd0bH9HLecxVXpNqsLwOt+6gJacxkwf5Wrvput4vFOmQm
2CdIoduIhMeGdnKIf8yErBJCEYX1bXyM0zIisg7DthsRvtxlALA4GRZIFSCWdLn7
4pjQTy+W9AJ6nsRDbOkpTJ8bEsV2K7hG5UvO3eyVITv/RsV5oVp+ylj1TmnoQddu
q5e2xkCI35DBxGxjC3OyusolMCg7kb9Am3SEEL4CIbyKb+xqW370Jb2t6qUszQtf
rZDqddShPWLB5PD+LU1CcJumjphkof1KYUX1Tn3IVZchimuNHfDI6utzPS/2ohK+
9vHNpmb3aIV5nGg3yy6TrDBlY7C/mhQY/Cr/33+OX9Xohwbo3x8Zj66XCgqmUNTx
5HIkgvSzQh3rjrKWHrq9/2fqgQIEY6OZxLnQSMafI6xPpLMFfEJJIgcKUf0jsgvN
xKKa+HiEDeJX7RH+kMyWHAMfrUlOllOHP/HMU7VBGaZi09HNWdgyff8E9Z6NM9ff
4Wnfwzy2ld6V3tTFbEFqdj4TFMATRWPVVdU2YK+ionXnnZxhBtb6XkNb2gu+r7Ya
uecvkFR93D92s2HmkcgwuRhjKl13hlHXSZxw2o5FbhSzIRx6RVaV1bjyxnpHoiC3
TBTX/bOrRjxCjGB7pVPCNrCO8ZoeAKlj2jJ51FKQNoKq3zQLGSzNel9QIqPobsrg
5MFu4S7N+bKywB+vrYSD1wOkDw5LNySF+Lzyk9SO9mA67E2rl/bga5XjjL/VCTky
EmE3HhwyBA7OAdsWEPlqHTQ0QhVkRaGGSvhA12x3QXuhwXRPHNeHibnSh2MzQQBW
544kx+SWiVToHd+t9jDInAAwr9mEiL3yFmYB/nl4I62p09vdu4gvfWGigSPsVQrv
hp/OGWksJqqWELI2jHsWZ407P610fHKAJRKqZy+1Ln+MaWwj21mvowgv05NRLKL/
etKRZIK8sHR6WELaAKLea1AH5tQUhbP6THshsHK1B6HtHTcBXKst5B/xrGu0oWUo
LYxireWu9lvS5faJMgEFWLrbfpy187kIwGWa2+8as2b526NgEX5dL7VsUN290q5H
jhQfw3zlTxwjpt5gd3YXetJCI63D3VEqXg6gGJ7+CLKHZXg41m+e7e1icngAFLv6
YQVAKFJjxw2apauLbpMZCe8oa0MvCTOaP+nXWIiS7SehTaEBI3OXKL+WRiMzTEAQ
0Uti0idULF5BjOOITUtPZ5S6rwx174kTLgbmS8M04gXt9cMpQW7yD2to8ZJOERBU
MIF0iu4gpVFdELTOFPmTK78+N0l8sVNmeV5a2cM7JB6HOOGW08YQBHT995oynfN5
1N/kQ0R/ktIFEN8087NLdbUhp4SXyFpIjDkP4L1c1H55iekWqk9d2/pMKO4Er7Cr
Rz+w7dnI+0iFuzCN5GcrTGYaORqSruXHGgkDvxvgEFoNKIEFzCvpyIcWwboxxvGs
qgdpItKQOmVDG5b9CAqkm/iSnWCpC3zeVY5k32hqstvLrcdFZrm0kQ/x89mjKVRe
Ptl47PMrlRmTaSl2nQaquQtkQny2cOrHvUDImr+wzzTbUnVoc1jOoSUcwXD/1EwC
NF0vI+saCQ2NGq8FGlABixfrWePFD0agG4TxeJOXyb+e7ScVicjzpuzsvTqm1T4n
1L5hbtOaHnLsj2vU/BYcYTDh8mTkbkjuzY9ZqF+SeEwHg9bkmT2XFAw+Tile/n2Q
eEB1DbfjKovSaahiAOgrQPiyndWZKqULPOxVuBnlsgnHB3msTBGXG1Dc6ORJU9uv
t0ellGBLX2D784NTTl43CEg4zvOuBz4v9kUD2Hw2drAGuev1O79CtRZk8z2De9iv
mBzdBodYC5c4Im2z2HluPRgY30obSo5et3/D4JiIPJ96VUyh4z6gWKQpy1O+A3FE
WUdfR7WR4BwnnFIkT4MzBkKG06dWAXozmd9YlzwYJb7sknSNt+MK7i5jdLVoaD3t
TtIZg7fbS+olmZ345VeRMhRyRHDzenOKqM2BC6JQdOGTjokTt+QsXh8U66KmJepx
DzMsyUSbLww9mmFCibEuHr0jEMMV+gM5yIqZn1s6+Yod4veQaoktRAGKyp7GcVyT
+tlceLy1vUcvT9ZCI5TVGxW4rHW8xL/axg/t30/gOdgSu837/02hjW0hS6hnORjp
BEZWbZZy9MdKXJSdE0CzzvkBAKxIokNJ2D7vN7EuKMaii7btB5MEZzWBoyk8F4oM
M1fJG5VzwRqbgF3l4GNPd7SiWIxiDZKfHkcKBRMqyHhOvlffH/prS/oqmxxNvGgx
I6aDKD6T8xjmGufuhmICiYeaOSFhTFFVTxDjLEDYsolfJWWXVOEHSgegeA/t4ePM
8t3Wzlt7GZCVfG/gv+PDf5UxHRYUny53zG/Dm3KhxHW90RY5dOLaSygTPa2uMRv9
iMXItgOUDXA1B6KDFhulHHEYGf0qTRx7fle3iRdhpG2ZdZ/dcPvfb0FkXacR+J5V
DC3o0GEbtWO/cmMwP7pTFgDwwpfPCMAn3fHuqkqVKsnH+gV5XMJ7R+ekiOktuaGO
At9T381EvWxKD3jciut0KAWTv7HNuEuNmNO/HrXuLUM8qhb5bd6mzdpzbRALW4fp
OXbF02WhUDcbdD4HqeVD5b4iD3aB46HVsJnZqkRH6MmDhbl8FYdSomPYVWMrNe3N
1Af+EWNgj7YZgMMRM5Scyu22tHaOYdNvoqwXDWvjNkuLuefLcXgeASRidksIMV2J
esBZv2zMm4nbWIij5OCVN32P0HIqjTCtc2EoI43LSfb1e5GNiTzdXw2Sn3nQvq2x
XzSEwsWSZQeABpZSZuQ6X2bnMI67Oov7U2mYsN4L3QZk22Pdz6TIuV+D9APLVtgY
tQ6au8nvM8lBxzXirshWU8gXmq7rsZkqucAJuFaxgvignX8SpliWaE0peOFlKmDA
FK28plMbkZPokWb0VTRPedTXXUL6RsS4C30FfdFSoznSeL1d6gNx8XMlsacpUJTD
tjujNK0OGLtezIHM4QofKWpSZt9LLyhb7ixvOWnwQHBUKOEbDSrV0E7GbBcXw3am
dnN9h1ojW2dXodRi+PEvUYiz+WDJb8c16GUjla773V3Dko3Z/2Ng1m8uD4ScYQ1B
TYG2gHz1bLsAq5T/+99AiEbuaWJ8/QTRHCrFFqiEgJ4YzosWv6tIiB0TbvGWsXXR
UEQXAnzSoUjHCPs13gGfI4T3ZtyufGkOZJBPx5J1SeAfINfA/EFc8uH/LV5WC2vb
dx0xm5Kv/AETn7Gh6ynnWZ5F0kuRqHDlSkhCx5fUIZDTjy8m8+THLzn5owWzgqu+
nLe9zHv1p3V2oOXhxg8zgVzMJRAhbJC54ms9tNSgfkThygdIZABHZQ0sarFZL9Ez
LkIdrMxRqb8YC1V6gjwkgVT9LPRWlhuOE/ErMb1UuVtt1Lts7+0QugnegPKrRbZZ
rGN+sKVJjaBNS0ysT8+kPI5EERayYxDpVL5nhnr1pwKB3hmoEkTrV9LHU60BVety
rUskQYqwhiD7qzDbU37r41BKsQpnmP7BShkb6OdMybq8qezJp5n/9KUAGQodL/ic
sac+sH4FmVLAwxxTFxi9owo+esc7LoJQM/CKLxf3ZDUseUE39Mf2ZQ0YnQxGuvkb
dFE71XBsRDtg253TKw/RCHjGYViBVhafTXNjBmMpLpmEFuD6kRgKPj5B2Pky0yLq
Aw2FiOimsF/wiikqhmnMT02m6l5y2l2SgRRe0zhKBHh9OhdBz+AGEBoJiEPdABA8
3+lf/Pz+XZVRvjSpIjNwk5HMLotuBEUMzkFxLK/YpgAo0NLv6tYfbrirQj8HzXna
JyDqul6pCI5cK0Tj/vSEbImSR0pSD2eCMy9aC6FOWF5lsflB3Y5Qf6cphsVw9aLx
zJYuu9EttdmJLJ90TyXUxTYVpAA1mRBnl31sEwwiwKH9W5Bg0LNYrQpLUm31BDb7
pVU/r8xN/dBRg5AJso5x+INZgGRQg9aJw/vWdunNzQsfr7Lg9l52qHhEcXPsCdqd
xHPIBKryqJMtrjdRlCTJWqjJUI9O19OOXR/o61xT4zIKQ+hQw8syYPw/R/Ssj7N7
llDQCbkjPt8ifFH4YUpy1ER7h9W1GzxF8D65+rOmfkl01tgrsqon8/0rTicyEqKZ
u7BiWQlqIO1dxfUrZkAK8WqKwQ25Vb4NKHUWZ0xk5y73IJ9sGygQD8wrzR8as4C3
Le9VI2wLqYFW/gs/btKvP2xjGYf+q+iOr84v4Vwq9SYcB9SseErZxlVIHiVAcHL0
ldEbxxMptQfLiJQtl91yRcRahwsfw69LMvWqZWqyO+w1sJQXHkcgG1m7HoAX/ouN
GQTjgoULVpSZ0ShAJSY4SQpQG0eK2rzy0e2P9gI5KgFT7y/MJoTWwvvN9PuWt/ch
lVxnOEpg8RYufveRd2CLUmawirvnYY2dYLbwMYPtuCI+B7Bc3PmjTdP/ncO+XeuG
nn2OaqfC/xxS77VD0+JKJW4a5L7aROKEA+wMolbWO1cuxQiEPXkEW8KHRav2SGdC
NkAkIzmF6kHX9cfN59V+ZW3mSFEbuHMiYZu/6+Pcs3dqiO/ZZY8ibW2nwk7OU3f+
UktPbVe37iqFLY62oG7E69Aqde716wCsNvfNv7M7b8e2CLqC9/Ry7ihPvX3EVNgc
QGB2WPBlYhNmP5b9QduWDyR897D8nC0xPJV4/sEGae9RbM00z6oV+W/sJD3d8zAV
QA+5/BY227QGgj178/kGa128UsRnC6MeneBdz32VKSZ6lwgTXaDd+3odKjkVzRN/
4VmC26cQvQ2ynCahnH6YilEXLrgAJd2QwQAGEvXH8Fr3BFuVgRMdrv4X6KPgm5Xx
V4rdjCxJGxPLC8RqIsySq53s3GqIZk+MWB9k/B/3oV2Ajo03DSdQq9BQiY96ADjU
Ex4zIEFlHCoStd5vg5b5WoR2BcVU0nQvsrDRvNZlkvqAKE5RAUwHzWL+eqJtKFe0
p/dM6djYq/1FPxoBvfU9t1S8psK+ni1XoUUgdHT2iSYnrwDVdMMKqTbabBCCeZV2
XP78/a0M0pok8cWbB7TF+2B6Qk5NW5bs6gtmaSwx04xqF9q8wrkcAgWU7htnnxGX
QJe3WHl4PoNv+TRxxMuW0MsUrYGErSQcVzNQqJ5Ox9oi8PEkvlgEYGeRH0+ivsa3
L0bWG8aCg75OP7hCQy+G5klLBTnMto9kTojyJ5whH4OCCiDY5ttOBBQ8J7vnx4eW
cQBlVh14Aas836+qcsE0mADp4G0saan65VFD0PzuXgLo0JWGM4r37Wxud8Vs+B5c
Sz230r33Zm1SSBu5MKOwFwmq2ewSzJhAn0tzZuHXNi9ZYrDZpjez75me2GKDMTTh
fXulKRIGnK2LT4ixazdl8ulAs3ShH/PCFanAUrvNns/t2ghL13m6Z9bYmgSvhzsb
6kT4mkqAqMKICyIqfl7w6PTx9+zdpL290DC6lrg7jWCp++OWsnQXZ2RTMfPZEtIs
Jz0nmuXedQ3xSNn6/FELjTScJGTvJRA/3vE4+TGFfvn7eerX7l4QlpTCMSHRIdNd
Hd++wGhWgei66fSZ4eOOMRG71IFbE32hnYnXY9MU+RNn9+f8RIOY/jVv4f/7Jw13
JlbcwdzTu0dG+xC1b22IA90cXdsyenIEj2vFKhsJambcw/3ssZTSxraDKKw++C49
Csru1UTEbgIOg4qdiN47nYfrXvUmhqRFJjm93Y4n1xYVyAQaKO+ovsfsC8y0Het2
zfqkWE0Xs63rCrWJpqWo6DX3X/Jbk33tLOGckWhkM4tQ2d+R6J48GTfGfrZu3eDk
Whj0XTdSZwJ9OdWpXAchL12vauKsxr/vaIIZczWTJTQriX8KmkWfwJnNUOYQsRAU
gX3YsJvUe2Htb+bJOzhI0Va19OCZMUb0tv5NrbjOqTpxzjCUUgkTnKR497QUs6Tu
IludIKSqaw2xhP6xDvrMNDYyYuDOhu/ITwEJSr+ywPo+fZevh1VKuJphKJhssJ8g
npqvjACHk7bVJeCHRj7VfDyveDiwnGIPUlSXEc6WTd8S0ZO9HNJgxzk7UKjSnbON
CU6MeTkhTm7tnNrLnvdqJC+olSSQlUVTeQXWxFE1kh/s0ravT7kuH80WVRXHHRTz
rNUiA2l4yQdVvA4sVMwceRvTjCsyW86Zkgu2KMPiU9t4QC1Pyk1X6llNoviIDJ0L
BtldXJ51GJhHsvxV8U6Y1/GQtV1DCpQ9kS/V00JGXNFXqkzusv88dW9ZCVY08ZdV
8cLoPKcVG2wDpbnOqn0ezDp13DuZLFnCopSmKlfIyj6yTf/P0VcyI9NJx3llFbIX
Ea5JGY47V1CMBhIIY6E8H83Gpyy4Mgze9vpUutVcNbybFzfD7Pgxwxkq0YeoUilx
d3lkZpgivarjkyacD6r3xB3c4fpEkm+IBt5eNyaAwzSrtH9tUj143hOu1IZNtYPN
XIKBVBoL30n1ta7nqcan2EBa2S+P2/Y34K7jVGmyLu1jSgAtP85wF+CTDm0+STRM
Yq8zUcTJFl+k5di/Gon7VlSteP+8IPrDbrsmemZ3mEKVma0BHNALlTyAK20PGdcF
StxFSTUxq13D5P50aYwbuSJol6GcN3Sgdx9pY4CzRnG+6o0isrnUfJtZJVVzfyXU
BKYrSjlDCeENgsJyaokdPFyLrpz35KAGQot+ST+awno5p/rEOctlRXtGHMyd0HUi
xdZ+AhI5QJNt5je+y+6Ko10csPPglNp8Ng4ft+A7EQN48aKee+mufJUyRwu1qdRw
oG5WCY2n55UxaF0PW6k9pKNf/gO0Q7F9hdFGSfmp5Lzi+TLJX6jbgbcI15MKr8jd
nyvZJNS2ALAOk8B6Ij7ahqhSMA3N7meFem/9Y3o+maZv1aYIMamfmlWWD4je3Tz0
Phhp+72PscfdXGacHEkzov7ro+E8VMwi2y01e8kIrrFQAalbA+9/pWlbnxip0c1w
QgVqFU9gaBJTPQxad16aNVO34nBrHU20Q+SV/EEZyyZdUVQ1HbxYmCpE5EoKWqmb
wqUOvdhpL3zp5xuJJzBmkYsmyjUu4HqBytHi1p+x93YozilAKV+b9jZWwxqiHzTF
UoUmnxqic887EEo1GCrNfmZF7qQH664ZtjRLDU/nCVP2thpn2rqaww6FI0+7jsey
DoF07jvMU8GPWz/nRgMpXRzsOHhee1GI+DjaDEH9xnwt4wE4kLS1Du4Pnk8GdaMr
GJcNnjkwNLTIxjW9Hr/wF3r9dsojxE46lrIRF26Os1nm1FZBQ08YVgXurXYHcVXL
5CJJH34772tePGreKzXqOobBE9TS56IsxllXyCk537QyESeGFLzNWj+O2wk+Bkmf
zLXzABqs+O8VRJCmPozop3N+7zw4FOwD9JLKf7z7UtphMhVGQ5OVvUZnFhmBRPx7
wDLRbcWg4rOQbeb88sy1eXOiH+Zbdh3Hb4sRkg07bROOPUKsnoJIqA3dTm0nwR4W
LzS+7IX1fTMSDe1JLUYecrhvMdFuSAWkzexHkKQYG3ubpVj4NJdNUNNjg6EfF3Tx
5duUopIl1/DyPY0N/6a7AFbODwhzYTG/3CslVur66QlzBWoRJxbEHvVrQkHxjEXn
OYshUsCfV+ojOlwwj6N4LcnnJ5z4U0eIjGoIV94WtVWx5d5CQeal4J8Dq2WOMXG0
AM3Qh6CEKAmj+D08BGUGMj0O/Agc3YlRNnwHI7py69pYdBH4fF6EIMxcxKzAasvf
qGqy4nJPEKp2mUblnrs1TbdFaoeWld5/uH6U3D+tePXhOgeLinr2YlFBKfjO1/ia
JvNn5z7QbRYM7p3S4NcWvqIhgxI4drJCQiCJanCFykRxadNqF4jYfNAzQU7cwybM
7r7k88wt/4amrpOISrIAqgv9sSfqe59QaZfjflBsaaLPOgKwVMUHB8YKWD2b54bq
JfRJzNweCt93XG5OkM9S7Kj4FDBvWWX2E75luko8lmBQuXKrbDlNwUCcbaDHfLz6
NB+M0aALuT4ySD7iLOwWP0RsV/PmO07KaDck3FkdG52VoIPYP1lWmp6qldwaAzuS
xxNb2Hs2SLfsdkUYzRWHEbAeRkMRZ2cbBu3YTKC1PAZ5hk/V6sMELLg0hnfCymjA
78A27XcprNlXR+G2t123vKp2p+ofN9k/IfozPTLc9V3EUUzIosHb0PvUVVTyo5RC
Pz1J6TiCpJWypiMY2PWiJxoGcLs27ZueaAGTapwhwCLbhC7GnhmcgzqeqRVRNHNr
zRh06K6jFYF9P5FVTek178wgggTEUlElaVO87c3rutn3/VrU7RTSFctYZnkUKlW7
zqdhh9PB9lUeYR1S6vJ3uSceZkFPne3eKAtd/BdSq0D1AM1rEOJ1rnmUybiRgIWd
F3R8Bq67KLhEOB2q2L8nHX3oHEDtjde42Jo0r3ArXf1tdMlDCteeLEas/y3lbzOG
VYP4dM0JJtIhBXYJFFd/IGzHij20vcUalGRUxiGs6dgfw8s4rOJ8TftLhNj80sik
d7gU2Cek+mh//sMshJkcyDjDfhPLzZdKwIVBFHB/3BQCMdxX3jzM5bJxklaER/Hp
vhT9b1xcw5yG5xGXEbKs/9N/BpY7Fog30vM3I+9LGrt4KIiQrJgt9aDxv6fRAGMb
EOHhyb1TvVxR6IO9on5t0xlVURKWMHjQLTHh9XWm9tYNR9a5f55plWoPnVs+PUWI
QQcKdeP8er/HUDehdKoPiZNhBhk8Rja7FndaKzCvhp6SuftidfSlsOYIupbwQGsP
6Q0BT4wDpvoT7G85ybmuaCswBlX8MpwyxprHAW0btRL/IgJJf3syZj1zvKbYUCDo
qcx3ELxLmNlblU4n+eq7oolm3oajCMYcXulkCxLpRVfBkMP0ZLu2BLw+8pUGK/zZ
GU2f73gucsbsbhnkG3SZhs5UndQXoap6U4flmRbUoXzrwggomXzi9ZcIaFYoclv4
q24mR2fMJUFHGfmhFS0IM88OGPEClYG7Mz/Jc3LH8ksfv43jtg9AvVncR7T1OLSq
rllnoaEASjbPHJAi1Q+7XhgSfD6JABT4LTmTsdGB6mgt8np2jIGWAdTv792yHsgl
UAMS9Tj+EjlP7DAqXKIEUA/k/0BlCVlUE3fzCdsLGHsv5EFarIhfAa+cdAtRN3Zp
+nyaltw5FqSO8LJxXo8D6gsOkjgHPoAVC/HCVICntfuDZDUbN2uOm4fRqbZwmasx
tnXLhbkMfoiAovTzSPuTPllXV+Z6zRQcDGAAYNHHZpeNSzbaa0utK08zfQfKP/rW
WveDwU/r00XsKig4viNq0zYP46Ds1k9/cDfQsCgQtfp4VRhDCw9yevhoi0oFhoPt
0KJHD6jIhIB0jfuw7WfZvhYlhQxT9xIhVWGWTz7B1Kis0ADdHWPYneg+ySGMgDdR
GG5HrAVtmXVesKazgbkVnDmwKwWGCrMqMTLjQ3GNLZN5mXBooWJNGbWOeFZF9bx7
ezMEVmD5N7Qy7T+COFW2iq9NZmELpHlS84Btr0SQPEZHc9d9YgYrdunYrIi0xNsR
6USq+rFghs3pBvvaEUbfXurlaTAfPwW2vGWPNXL/l5N0OD/KMGofWzYLICULMWk+
VQghgqqFGTz7B8cZjWicQWYcu7H1JmMPvSHTFPbU3UGj9ZOmOcqjkM6l4Se/Qj7C
J+Q7AHcCh4gv72ZHaA3pb/+8HHVQ2+JxTnGKsuZMThaK+x3Z4n1giS8BsHDgr/yj
vFp5OPleuP3XW+WPD20+UHkpFb3isWJ+zZj756K9pvhxwEbrHdBcExEVLik0eQ9S
luJG6mkgZMpndSJIq0BOr25vWKi5kubXgufUYKbGa1X/8QtMKdDz7AJUU62/zMDm
77ANMW8dgbPUQZj9fQQzSmqMcWBjgxITeB7GbBvcBhTCwfk/AHUGliZWU3OZ7dED
GnkZWHvrEfm8yvEGHloAJuK4JGG+T8G7y6l1F4ZALuhI0PD2nUK/A6vWkXP4oLaE
FOnTFOnNx11pndbTRCfprV20clBaKjK0MFwQOXxe37og4bqb2R2SBwYiqQqSNyu2
40l6vhIVYp0/uYbeolcrR8Z+LXJGynPXDiMmomwxpRUVgNUtDXn9KiYKO93F7snB
Cj9npZYHUUG6COdCRCOCdvHfGEiz06JCHkenX5CgdsPkYsbB0WTxPkem9gLbfAXt
q4LKKIM8PBXC/cj9uLi773j8F47QL6t4I3+3dsDMWhLdwo3ry6UDuEKqeq/j9kGY
+mYIZ0jHAOIYZ4DcJsSmvBzM6Wjn1OExJ/FNlYtkXEmpy/L69Fe0U2t8RDJIromS
g6ch+v1IKGdHO8jSs2qCahLYxGaG4PIjsr8uTayChxhQfscCCPJ7HBiJVAJqSmRj
7NpWcmUZavUOr89Zh/G2utTZZL6bIqzx8dtNLgoNkpD5iPi1QhPR8WpNzv1kzz1m
bP7X4DSNrYFDGwGVbGvZ3pcSQU3s5n2cjZnx1LYgd4bNhXpOqhClfYaj8LAjBJfL
MRA0mm+qG4OfdPbMMugMQu4hyQq8B7Rwm4rfr2+pj9LnbIHrm7fdgKvSiD2EDb3D
f28W6YoOwkVECJ21mBafs4y3RK/MoFKkCsoeJ5Psk1qwQK5blre5XDI4TurwbwIY
vvdXLYA198RgRVWtWU1qDoMeIk9NMcvN8U1NZqFlPtqmkTwrCyvA8XgtdiI/9r3I
GN5UYdIPej6arwnqoEuFttfjoV63Af0X5bsj/aS8HQQPK21V5LmZddXN9MwgPGxL
HcMY1Y70hzfu2l30JWj7kyVwKDSWYD0OqxHrk3Q2XeMl8Gq6+5km+YVG71aCcSnY
aPUlasoeAVgFCoBrPZ8Ob7xMGP2zfCv2Tbp7CQuUlI1NooSMftVGv26fs8mhcOqf
LH+dukOmElQdftZiotBB/USTWE8ukbY3avp2KDf0dt57N/Re0AN9nburQPV8bAI2
gc4ORYOrIoKbGQHaUjbbfanj54rUU+QXAUusgg48Xc5kzeO4VQfOyqsSeJ1HJ+es
/sdrKjEPu+jW79SLg8wzurAVtZmjwICikM+UlXVKQ3TBsvumeTZGy/2nEjNlbRLb
YdcVXPY3BFb3KBadd6qzz/0nGwOGPw6GuEDzHo3rEC5hhfhKGjVQNOHUWOFWREZ4
zjhA8n2X1Vik9ucdKYWd6C3iq6zaKMgPMgyo9NWUwVGpH4ggygyX+Db1VkLTfCkH
/XLkGsv7UKW8oYmzSGaR/GfPp1gMdvc+Zca32K+Ch3CRJV3mIa1P0KaboCal/dtb
S8F253RKTPXv28LCrwWOVmYp/23b2mOh26OnC9JrOZbz+r1K1Qiv2sNRlNaQuPS9
U4PlFg7eksrTtX2CPtbjdR9o9OUMpDxfzdzFDjbSLK+eT356eNnS7rMyltAZn+hh
5X0ddpRDNk7eGdVrUMGVSd9fmFN09JWARGq491u1zg3Ys9Tr2a1n+HzZ30XCAygL
5M0hJBEMatA+dyPysTFLRr2M+f7LQjWrzCQIIeJGUclVYZ+ynf3FWOpkXpeXib13
0Yqyw1aeUulKunG1nw/5JUM5xK8iIQIztjpK026MWAZaIEsiD6MeP1tKSe4UH2r9
BsdwDq2rWsMv7SreuBzDM0uZQ22fBFWR5RhroQGoeQzL/Dyeno1+AEgJkQnyUH9j
QIqtT2AZ6UJakdoEsmFsrzYX14F5Xyd9l/nvUNQdFT7LIutgndzJKiH6JmPo9ilp
vCAZxdBUdJfeWsgpebgo/aujbgfclyfUtYD/jbjx7ZvzM+A1rSq/PBGM/XN6WuWc
YNKMbczejqYye47kqp0hULXKODsJk+6AggP/AxkkxIteiA89UMv4ljSFuHZrvW2f
kyDisGrJzmcwqMOJS2NvMsAJL36GiCtrPIP3ROgh1oda45sl6Zdf7K+tak6GgGDm
NME2FLN0gf4m/kHhtK4UOO0UVMiyntAd/PvHxBSOUO/KZWFjoZUXbQ0fwJCiJZmJ
Ap3WBeK2uK/sSsPgwolVxE+jGY4BVdZkEF871pcIu3E2ArEY3rsc444OYCXqHCsL
ggyxagbKdQ2ryUMaJwIPcswADXbvW1FGYxVBCxLUNNr81dJYjryJ5hON7nDoU91P
OYw6i71EykNVe65Z3xgOBLXl+8u99/NkfIp/fVKLoXqX3a4vLCLcml4SmgY1MYn0
VJ3kyeTCjpmCAlZHJQfFF5kqOqm0Fvf3VWiAXK7cNvmdv5RcyT3Ha4Ou4mO6CMHe
KrKo7WO6/XLrzBIu2qeQaCMxstaOUIzQ/UAGPQ8H3fq+CEH1sc1vYnwEFNnFkP2x
f2+k+MjTRZej56syJBXnOwee3Q3IyFFG8vf6u/iT0SFbIaW+xyKZ7WpiNUsCiSwS
v/vf64+tPzm3XKEFXXHrD6u7vh+v2I2Azs6FNxYfOytXiAM+nCIOO+7lN9rKuEeA
1n0meSd4afqYefHHXO0PqllJ+TOHpPQTS8VKDfvLRx4Ml72YUn5hIo648OoYvWuq
5oy3xQMEdaD/YKGZxwZRfxlGI7AGytv3U5GPqCb1BEl6uIJX1neZqlNe1rdofP3+
tS1CiUyzXZHpReW/Qj1fgvZrXBvCWsS8XcfFY72j0py04xSXGbfsrIBNlXSqDM29
4BomEt2uZzkoq38b2AejlFhqYqnXWv1rGdK8DpmhDVo7Vq4Y0lLjXomfGWfWzcOu
Uj4hbnDBbgs63JBqqUunG/xLkbumTTTTMVJgta05jMcNuNZKyY1drbIB1Mzi2Y5s
HmlZf4Pwh/DdZeNIPDCOMV2kplqA6/ckcPueuvTIEVaw3am4i+/Ol3aHi7bp9J4R
5zExk4e5KyiX5/ZmZ/7gTNUINE2Bt41gBo3OjWRYP5UkH5fYhlP6l7HZ8kHPA/LW
DHLuNuImjq/POhxaVmk5svIAj98HKL1/W689GaIWqUmr296rH+P+ov6hvfvwv8gv
CVWd8vgLoOjLSn+KskjkBAxfbY45zxUp64cyFwefLrMDmaanJ9fUISQLzechy4ic
508xruutiJEUNRfAgOrbd9w6sSBUZfPag2CqLJgVvIjNSF8jz6HhUIvLKRckhpfT
a/vG00H/aLOAzAPhdyvskt0dnlm84w62hOCfuGjEptgZzyKUAPyiP3atrnCggt3x
E7Cd3IlK+L+gIOPSpi5wOC5QC9p4xW3G+D2NJy2rApy744RokHQN/ki5I6wgiRCl
KsMR0mE9YUeDR7R+mDH7O5FPIKEulQJcwSd2dQMZFfK2GEr5jPnxpRNJ6dX3LTAQ
xeJLZwU4X0BQ2EvUx9b+F68rlC0ZmOcZWZSLpyZRgEeH6/UTL7Br9TfHRjNMZrRb
YCVKglBL5dGfEfejgMn3YsXW0eX82wKrOjuuT+bnfYkpnQ4024BeQaMFarGMZE34
5ZN8qhX0oxGvJjCsu5jtnw/gTw9bqlQxK0DqFAuTeN3KFGS2f/rePghf4Y0C1I5l
0Ygx52WZxX2OSBqME1Rf4DZg2oS9DdnDJUCzZUEu805+5gq6bihLDdPPTOFWch1V
BidESs09f0K8JH1j8PZpVKSREclPe/8T+ZpMJw3jNWPSZHKWZOuIBX7bQP5FsJrE
MmaHOSwJi+4wylnBwvqJYD+tg8G29HEg4b2O7/cLPMBmspXIKKHDWwGE/79fqxv/
KrNqhTfzMQVIlck8z1uXfOs49Pc06gcLbeG1DaDgFg9afJOCXLfuGdJibomZ1kFm
Pfbikk792Qh8b2wwu2zHn/7JgNukd5ObnIXUFB6avZLMh9CGwkR7UnScTSYZRnYs
VVsNZV3c28wGhGxsL5arSH8UrKUKkO5gGdzVJvUbHg2joCaJFn/JBWvxrKaA/XWA
AA7an6FoRNL7xb9IfLYl10wUkRTwdJeO5+cWwm60A3nsogcYGgtukQ05m1tmI6bW
O96MVorKtBXX3CB6mxukp0FPY9b8cYKHQvXtj5cfmSxCKgTKWsP6cUGtAz8NheHE
a/ThE5wlYOw8kXfVQ5U9mzdikOChFF/TNfBCf9hUPtLolZiELbgr9nqVeJoU0Gi8
CLXSdTQxckcpX7KujjxwEfebEMZSgPvLWtn+pmktgQdJG4rU1C1U18LkPByX2UeW
/571rDLvkewz+X/YfrZvecnVD7kYwJlaFlvRVAMtA+5KmsGLlK/ooMgRbN687mmn
EucUf/AHmND+4jxziWg+Rarz7d0EZviYwoXjaAZ0astENbL6rXp9ZABVEw1lHTIv
nYChSbuc8TGZY/xWjSfhNDLLPFhIOmS7KTEZ0Bvg0LKkfo/vB4zSJB3IAbY6FwYa
YrdCXBmozwNm+BV1T86Ac8dWU1RKA2aIlLwIz2tx0UPdtqZ0P8U+VNqA0rhi9koU
9/rfpBp38qPxpCeXMV19q9AbEs5k74GUYqZjvQ5VhLBdgWuF1iY91DoB8zg/MY8G
G6N60UqDFVmN431SV4FRMQi3D0XfJYpPyJZi2DQjB/z8m9tVhOg4yBEFez5qt0MV
UjWqWOLRSKD1HpK5KtGJFTGFYQf4r9MeCRhAExrpZQtt3jLGLIkUbSEs2GQSsfha
7ANsv2BpfeGQngTb1cZtgsDKoOuwdr7Ia41gNTr5wmamSC8Tm4Uh6u8Xvot6MIqZ
B68IcxAuY5eVRPneTQC8uB0rRcxNAa6NYpG8Z9Cr+Y0MUxq7Kl5Hvb8mzbwlL6Gf
JYDhKWbGEDUJXmIMzTlagjxBk9tiIyqstZv0NvjBxeftHdt67AVpcqyDxlyxQrys
FggyJnRqBZcfnutvqzw18urOswkprLqiIj01FkdwNwbycE0jCNdWFjEHbApkMdRq
tmv0XySTCOb3ae8NcVQ4s/YRmgtxzIi40OyfOBdo72TQMJb+s8bVgT6tGyLUzVFv
B7XQrnifi4HTpWeQ7WvrTKOyPcam1CeumeUpKSJWkliMJI0/iE+0aGHVRomh+qdu
9cMw8pBgCAFecsFLVXEw2Fip6+O5O7F+VM/gKUMN5koB+mMy7mvCFiDh9Qjz0sq5
+C9gMIE/vC5kIlL2qgnVYNVp3letAGmr+iFiy8wBXuRGzYZaH4UXYtrDLTPYxeV/
8h+HzntyFooFAFXnrZ7KGXzDMT2iT0dM3H8ZNG4LTJP0sVeSNcFr47PJsGYTPmjg
3BC6uMl6nCSxBcPJtL53Az9iqxDWll+dzlCQZShI/xf0r6S+obDFs3AWXcsegr1e
WTNO6Wdpq2ILRUGCcJdPTTcgeo13CEdQQokWw+HQ1kzmC8Sop+RJe32cZsOTOCnO
g8zMUstR2tCU3Gxh5FLpCV0OyLnHtLm4vux55yvYkRrKowYBxoJJylZSJ9g8jWM1
lJ0vEJlE6AUMHJ/bjPTE8XMQMZNEBAgcdMQ4CqTtvP5/uXYAyZ0Hju7hKb9Md3J/
Saiz5BB33BLoXw3m8aWNohONM8BsF+c1ypxzWtyr+KZdW05agBA4TZ4tNe7AVXGX
JyOCGzDXbJmMTz6stITWfXaTCNEvo80vk+fnmE6nnRvDVapa+O6OnDHSHq2AYcdx
jG3KN6cQuB7qg85SY7TPWbP22oons8NOIN2xahNO/DIjtMT9UvFQLogZsHjICi45
kY2ZtZcVwDX+V4NpVtox4PCaBU12zrhP1ohlb0sofWh1fkMD4AJHNhuqParsTHlk
e6M0YGt3gBe/c94v3T8AxM3nMUpJBVDfOfV+p2C3u0a75rDVW7TQhhK+49QfIame
gvpe2XsUmqnaKbrJ9u0vH1D9DZHV3IsGwaIbPauQI/ajzqjKuFavO9/mtELVC7Ne
zFa1UyfkKnJwWmoqc5L7D5w+Br5iDI7ayjGQp2KVUsO6A02kDp0c+TmpYmIY7R34
/keKmNfl9qmM2Y04WlZgZjIlb6MyUxQeDCW2J/JeOqke/OE8lshjJRHl9XdvvBwp
uLB+uylIiHSamnhGM9xtzrzm8CwVGWboz1CufjJWL08LEaVN8CTAp2OfuB5zYE8B
KwA99FjcPM1H6TkZ0HdteoA8IBU5AYYixCqpCsPaWstmd+qrlZWdh8Ty2a8cEzl+
cxpNyjmgwC0MbDRfdZq8BE8hEPsneLRZn7/a0k0E8mM2DeKgd8VyQPGoaqyS0VUa
R4FE1BUxQ5qivMuRSJRpRL2GHEOhZKf72+WXAKhSyAjtCDxiXT29v/09csNFfEd3
5f0yeVn6qZsMOBwRTVLIz8d9RbEe6CBbPiN5dyOxUl277/xdhsWGCCmwsTbDegE5
PacMT9J9g3Gw869YJ9nNkbIbqm3EzrYKcJ9EVqvGPnt1n5kR6iR3IqcbwWpyxuCq
tFhcgCLfUzw1LIop18w9upqoPdzhalNRWPNsn8FpLrsFPeSWwSC4CCRjh/1PPjy+
CFyN8XeZffGuTW7GNZtA3PJtgZv5GFRjj6CzYYBGScSOKihC5P3MeosBrqCckN+m
/PzSgC8sHsERgVq6XGZXt3iPGjwVvPTJ3p4r0mQLsAWHoNsHPXAhsQVLYr7UJnLG
j7n9702Szu5IZ4BlQCfDZ5//7foHPSwpCO335fAqQ4iljsotSmfTJZuvIGleXUw3
kUPUsivFjsQc+HAXEFD8GR7uBDK4s15Z86VDapMEvs5TudrKdlq4SdS5sDOBlVbz
imRKnrONmGb4Pl+5QxsSzY2OgvkPlk8yhFkOTuHCa+3d6iBDqguuXINVZ/Du3TKT
WSG8KhnPocHdFFIccoFWSIAifrLT9sGO+VPiqjxzrpqOUEQV7qupqfaLwTDuFtvr
NVZ0cZUcP7PlkYhHxzV8NM/fixf+WPpezJnjAaw3yb1vgsX2INBIlIt0HePqPM9e
Dj0pdGuiemyvjD4QrmvQvr8Jf6apvhbohxNonLsfohQAusoCNcchV1IyOJCGyioW
m+h5d1md0MT7WOcDLO1l0fHChCp+4Oslu2VAVXjRNKmnhE6S1iJvUF3mmqIANRBw
e37T3zJ44tOKbK4FQPcFYBIpvc+bcrhzOFqEB6m3C3pQoYShKNtaBJYkJ16ggC4M
cYcaozn2bivovxM1xYkb86znjlYjT/ObMQaBvdMRgGRzHDTabIDEP7lsC8zaGVLx
ngrdPPxacxScBCpKc07TFIqXNllDbd409LQ9hDIjs5zNEcwmy/W6a/DcVXyu1llA
KPeWAB2kkLIEmIi/0/XwKFrf6kW10WzIcQMjr4Fvfn/QEeA1Mj1hV52txAkZ2l1J
YhCxNicTzBZN5XQH8shB38dT4IQiYo9uP3EZ6E+3en3q7lXskMbh2M3BaXq3Mi2H
Hsx03wMypk8hcNn0CQ5dVa3/WAt0io68DvUcruHE9Ch+hsO6LZFVppa2pdR5z5B1
bc8YhHDOzrxdDoUP//tMvn9pHjBB27elp5ugWSCerASDHL/yQ0AV3id8ZvjYRoHS
QGdhJ74Ycx9XNcIgfpD5UVyrvub3q/hfEHjorFxboE/Xx9nxg0Co6jquxhMFzhVB
7cijKNm+k0mz6UQ9DbOeXZj+KJVzEa0x7321sJ1ohlNsV6a0J5UvBlAb0xAjUtGy
H1klI3eO0HABrIjzUB+foHjK4XZkzRGfZ3938e6pNiSVqBrAY0QgoXg2eNNQPKPQ
Gt2cDI/zXQn1TDbzZG6rCDgDOstV3kYql0DpKQ43HDRctskYQNIMY/FUjgSFyK7m
3q8dUpHjWQznPVoBjijXHZwLN/a8XfFctj3RTDFT3p0Y2pLUCLH31z4uEixWAGI7
urhP1O8S8hd+OkNCGTpXoPp3pS5+SAxN8ZdDRS/j6oJhEECJWJedTx7snoWLRxiW
E7yoJZdoqkSwBr/sYaF9hM7zgrZ7g1NsZ1O/8s8yGa+s3EJqSmguzn0aD/06AfPY
OqvaIM7hQXiaYw00RI9NAOjL/sKgNFGWpxX/K3IFpiZCt9z0S42K2AoS8+C4okKS
B4OU/9ha+AJX9NCD5PJC0p6EpNzzr7PVae4sC1Cx6MX94ia22vDExMOrEZmC+3gs
XEzJtIyEm3uY43y8YSIFMgp8xLWGZAcv9dH2QRaXnGibx0yBxl/+LGHngVt4I11y
PZx48NSxS3iMX/qfiAeeIRUtZGgYN80rzCw361FxIFm4S/tSrsFmOL9t7BVEHt3N
a+s28gniP5Wr8PEc4murUtxMfFdO+ZFRDs0oa99TlyODFGl3hZ8IlW8YVQBLH8zi
TZ6k04MZVY4PsVdES+cQOqxzf2u4Ixfak9cuwzqfMFYX6RQaFL9SvEyU+6Ah9dCw
3XyD3brSSZr6RK71vsB1p+jrDOWOnD0BdjUI/gRtUNQ7XqI9+Zt+Z/QG8/q2Vv7s
M9zykdlbXDl8QhRJhpKxl9Xt94/7+YXuRqwagXRC8F8+1icw8KnHl19+CL8R2xxM
WN0/tSoJKJ4XK20dxbXGtDy/64izcI/lrg9sVUHZvB+XQRWTINNm8g9iNn/xUpkk
CEG1OBeUIwby3ek5m99t70u2SKiHF8pBD20Tjm63ub4C5E8R2KnHu6bzGemuW7Ml
9Jn5SsPaFKPnpMPKcD0V7Qe4YLVKknUj0UN0qhoI7T73aZhVgiXeAMfcYi6uMpsA
Zi7MLMjXSMpgZHJWkVRjvMtncC+PFFewRYuhFgWjWPBz3ogK5T4XHQjfRWN7UTnE
JLlqAja6U81JYEj8usN8LFJaDYR29BYiqTQFKup9Jq6xrL0DZa8ViWX3NjBYqdGT
adQdC7qwiM9xm6OBLHXTWDWrz3HaOFH6TFe8oqRTdQHpFRDNTds7c1Rn7smcqIjz
dsNpo5qjel2/dGdjR0nQxeUjxYjBbPXb8wD14D+nIolcbdXLi4sxvxCjMDGZYPnj
Vfy/bDS3hfzL4HbmCbR5hmiupsuyioH61COLpeUGK9SeDhRjNYBDIQJDqacash9v
9mWu+3Fed02zHMAT6RhRKVmua10dLgcEiIW+ELUGh+6C8OnNcXK/DMHLqNuZO744
EP3EC2CS85yWuCH1QkFUK0b4Q3/1JogJyFqHdDGbP2fd37JB+H3aBlU//+YDD6Kl
zsfhA9T4Tg39zqtuJjBCae12JStkQYGrRiz+Qo9IbpkbMfAAQgV9rqNkQgHpqAsy
Zl06XYhoiVM/WxLFPncHgri/jR/FkoheodrWJyYYZqDvRPkR4W/V8KqmxGU0un9W
13Zlolicq2W2mXxdVU4WkDIEMpq2fU4iiLCC3psqkNZN4FWK7XhT+EbTEtSnyN87
8dQxbki188AVjoDksCbAj73HrFLn1qx6w47dX10dxTAa2jKOIU9EwBFBbyg28Iga
hRETXc+LnUNuYhcDda8fABAgmaC1LkmjebbiBbAz1mFTZ6BeX5QRj0RP2yVSR1SY
qI70N+3Ofos5MOHlEMkuQxz045YzQE09VwqGFxd4OXfidXrXNiACEIvC+RYURujx
5FoMATZuuj/fgs8u7JjgBtRjALz9uKNrRZ6tCbFkEvPd9jpDiHQFIgxil1m+AHAm
scF5Ostj6v20UfdrRt0AbdhZXM/2RECN8pcdslGnCjhs20yz2f32XKEnvaVbSBrI
HZLD3RDY6QxZ+oFv0GDmXaQyTB6GsjlFAVG38cWJDboLIoZHBpecdZq+kgKAlwk1
yAo1vfHVLvjTkXX5D/nyimun1NAf8w4VrWanESPD0YA5rGlrVZ0oeV1r/UWA28Im
7Ll0DUU9MdAp4gVy25EmTcCzGrMeVUoGL/pllp7iYLyaIPabhYpDKUhwljCzI0ta
n/VOPuzmS2pE2cEXCIOp/VjEdJswdJTZU8gPFt5DfV3+8+aYijzprX54HbaMcKXt
sBUMkaOomEWsUz3xzNpUZzx/6FvyC2Ezpf4+H/8UTgtWfJn8iLWHreT0e1DjAl8E
8hScIdERSLw3q8Y91Mw9rBEkax8dbe6Yfnsl3+8P/KuQUf09gpam/xLqOnXi4LrV
16DEDqlOmlIPSarYm34jNk8fcOnJD7kT+ZkcFnasM3rnZkrqUgI+jILUGVQiaIhd
/2ToFiGmYJPgSgVfXKJE/A0FE7IC97TgXXAO2nqmkzg1ZBRbek77X/v0/RTsP5c7
59La76brdZMRyW0KD1rMKel0ehS04BPAqn+UBg0pEYGrLS0uEYPsIGUx0XohLaRc
TYJ/s4X5mUCz92b2AsgWVu+I736qefCsifN4mXj+iIwFQb5pQO21H4PnZyF+XIQK
gR3kPUuLQsa+jBRweI3b5eksBQNkaziVMKVhmeFOX0s9Sh5Zoze4h+RbWT2QxLxd
sZhpY0ciHMvItUzHdEiRraM4Gszt3aEXpwI7hZtsxBpFH5YohOM9XXsLvKtpTPK+
HaXLzjDLXhChq/iH+yt44VtNxUi2jTbOWhOPlPJ1MIKOLDWZbMGATMAaG1NdFRkb
y6mzft4FPXqenZWnW/uJM7UhP6ooZXE6isY400H3VDGFfiJ+dmMYHae7WdIZJt3I
RyLk8O9rz/7XzAskqsFG1WOA9wsMBjbFG9APRcC/l/u5uDyuoxTLx29jJRdA1bFC
WM7jdI3QB7FkTFG5KbtaZ9/4TtHwVvytCr/UlvntBh0lgME69XP1oOBVlBDyL+ts
RWtSdpF0TQLiNFjCtq5MjLxFuGp2t+vHvIBtqr1xP1+rAgN/FW0tT2yKVcGDRN1P
eKnVxoGe+H0cA+/WbGzAVJhJTU9cVCV7lv4CZfTcKPOAV28BCMNJguEMSMbz1FtF
Zx1ZQy12IpedmaBaujUUvL7mkk/z2sJ8q0kod5yz4Go8otx/CZqz5G0G9yIYly2S
SHgM3ubIBh5jPXrhQcQ7VztdtpwD8gB5/6krzXwt/QTQS8DaTZosgTBGSLYCow2F
ImMnio4ZkWwz0Chkg+CeQWxKYCgOVO1vUFCfkWTrOO3foxQV3fXoMSZSBKDFksGf
DKf46SwxewFCYe6LStH+ZfA3+bjHT6y8A0NK0v6geFUyTyBiDpY4cg5AZ0Zxf7YW
E6wgjyveS2UEmfWuhzHmBF0Na6fa95EbCCEICM42TpWWIqGxA3tIU27QmKtlXCN7
j4kilS09+7DkIqzXXoFDJ6ZW6mMANlYKrIZ7PtcDaG0z0e0Z1xvBLLKQr1oZp3DD
Cj+R2NLkgClCsluBulYByaB46mTgX+wcvxtu3O8hkrJ/QmlXuOcWFA6EaBlAZxMe
rh7XYI+s3B+Q+rFujhk4R5b6WYHm05f4HzJh+LWhXhbvd2wrw6gb3sL0ZMxGg3FJ
1QZHlW+uz0PwImcQVYlQ/pYWvi1RXo24OfqOOgQbQgx61mk2YJ6vpQ748l7oJvp5
bAZURHFWMQ9vqinT5D6snlCLUkgu6+Dfp5HPF0oPzWBnWfuxpqv1QOO7Omom1zT8
hxfuNfAKlrYUbpY2xWFJkArTnq4JcrQ3ZLi3wtEdD5ZwVRUjpdxcXc4b4EPASuXN
KqPJK6CF9ulPQIsak4ZNwFxMgJojYXjAYzHCdNno4d3fFAmZ+ecNIR2eNcD9rSzx
/rDNecYXVfjrXSREhLknX+V4ikWL57vdeHo66YDyKG+fatLkP+o3Z5jrMDbz1DJe
iU9/iIsE6dmHOJbiOmgIB2kB3OV4JZcI+oSsdrPwpS5T4AQnnRy6iXAsZwWttFF5
XOJ7lZziszWrO33lnvgK8mTbDgSCxZd8mbheqZLuxyUgE6lPGgZg8ufIcHVAjMlg
OwU3K66nAJM1+fEQ0nDYDDRmjhnK77ScvsMkKaXK5E2P5pgIqx490w952JGr7m8/
YYNnIEH5MxCzeCDoCTS/xCVjCGWBSNbWb2vXuJkCOMRp4M2/dLsvpynV1fSaKLFR
y8yAQSftB434VdeOGFUsIxNAUVw9gp7KOxlcF1NAllU/hlc06X8S7u2j6+DwoRnW
Z2Lz8wUnSQnXvVaFydvLm/iz8Tt5S6QtSmUa/Sfat391AjLJrrRu3kVtW+E+hvS3
r/1PI4pAVqYPjQLmU2dXAdhHU0s0qd3SzHi6dVsvVgGz5EQWNawJWKaI8NU+Ef7Q
wqKkbPbzFworLHkBIHm1yUdhcMokFbrmzOOpzCFI9U4Rzmu1Vi/Um6+u9E9UfCtG
qk26DxiQz+SYopwxDY2no7CbpZCfbuGGdw6bM7SFtHbvwodWR4jxuMzdicuqhLcQ
Tkt81jL32l8Stbsp/2XqmgRmHz7gc65S2RsBCGjISV5qjKh2HyPe1EOLEUttG6W2
rpLQ7SDQLtfU+j0sFJJOEzwMy6VUAFM8Y3XmY4OuXNeBC9Zj+mx8Tpffm8w+d0wE
QCTRYMjAcnrr8cWQWCadifDZbaDTVPjeFWJfFyoOms8wmysMMJABEBa0Dc31JpWA
HvDXAEHYXGzJdTh7iNLDKBD5At8dBh8Hgois6bNvhmsDmdPXnYem/WfCdPsbjYVK
xUU3tvkAwGHs7o9n8MAbwAxiZ/We810BIErV6U2FixnMdNR/o9k3NfD7iEdtLaTw
ErlbBtJR1goFTUITuf6nWE+TRlWYLsfrRWELFCYaibwywHAaYoGynslB8wx7u/4I
XoU9wFa5COEFPMxFa/f7wED5UVTsRjfiac9ZzF8GbhyMnxJmRXvYt4IXKDkwdmeI
Zbdit21I4JSRRvj/IDBYlIUKIWEjowfB+J8G0f+s8S+ol9ziKBLxPOEtcAuomP1u
MK+kxPJU1uHt/L6j5ez3qkm6eoCyZ6lTsp5oJiBUULFkOv0nsFAIlsMKbsSCs9Ki
Hv0K+J1hcRmPW8bLhBIac/1m1gtzOquWWX5D/tcIMICKVlEfKU/elUObXekWfKOo
22p3iaRgBsDm7aG8xVRlp16O29etNtZ9JqDbYxto5AHJMyfG+ReoK+OEHrZlLWlF
XUPUeao0IyZIEQwvQKYdNd6IJduv37meFy9wrvZnm5pr5xqGRqqt/Zds/19Z9lcx
wplA0JvZVy18FaJ81a28Mu4OO6K9mmSGmNEoL068ESR9S9+w33sVnZPHR/GZU8cY
IuusNW4RkOQr1riHJ4ljBdbkxhn6pavRlwy+vu75PgNr5dLLK+Y0Xm7tl6dPi/kN
qIdCAl+MFX0EeUtKwquzuqO68GvyVTLVtmnFvmXTsbbPaQlkslJ/Id9KnE6QlWFQ
QG+OXnVXDkH7hPbJi2ZpdJpc5pYMO2PYa+xh4hITnu2z9enQOHbz1IGt7V5qhQ7T
7tzuZ4xg0VKemZHtvwuFaHtw4jGh2hWXpXhv3837At6/TuS58bwPsewPFJLFqvy9
LB7GBe5plSCFLQvf0NGcSV3n8gFl2wnRAAvHU+8ElW8kYHRiHl2yS8fpnAdnRDtY
uOYpt/m4l7fXQ0wZrp4IlmKe4EQ8nYuggBcIBoFU1WeP0F2xlcXj+g96vP7XJppe
FVIVst4kol5YQzCjrHrTiuSkKYraXxjhUFZNlpKz38UTLqGJu0IBZWY47F3TwBEf
bSf+bSfSyNZJ/HgIFObFnkqie0jgmOUk81Oj/BGaGpGZtjvJMsZaUuAXIkqH9qeY
mN6pWjBlpQUvO2oc9IxkP5hZELrM/lMW/uk8P0f0MbD0VuAyagjoBh6Bzj8t1fdf
8kDmk1NtJIFZl7EMwAwxihrG3qGblPq5MHu/TdU7+a304P+lgHg/7B+AxS8JXILT
CLxv97T0/pAF3OuJ3eucq+u+e9JsZWbwYMRyBk1khTxhk27YfQjBDwTZkeehu3f4
qqhjPaTAfGtKtQLjI/kS45nVrCp11xt22PtVbY9Iu8xl7l2miPhyc1uMRnjNKMDR
D6yqJ9LwMIQhU+QnEgB0uapfJtMRZCvHEaL4M4DAgegly6PZx9HiDXme62tPjR2E
Ai2KO/gFJxXxh1AQGpXV0uapsTAxKimiLH4Wr+8BEkM7a5zK/4+jL5oqcAN7iTwG
DGHrLjRkNWTGKMYqz0eyQEXbZVoIcJHK/7PZQ7tuVbh2YBgiirdGTL4CHUA8nPfn
0u8PqqrFz24Ug3jF/jUR3G6NXTxgUEhoatf7oqF/Khtc/55jsdiJci6jc6seX+Kr
Diz8ND0pi6wcLffe1FASygctdkdqzY6QEJPXL2QQuPnQGwI3c+2eAMHvjX7tVIq4
Hz20oM5W7dAoLIl8vvlxLijKdI+vBuCcf5pzoQhmZVGYoudPmtOmxsaDzhFTEMQz
sIUKahpz6+E8QZ875z6jHbBiVHllQGw85WMXa7H5pEhHp44kgSGM515IMaXI0pI2
LqpvGE9oXxmq5r4eXEawsuMeV7oDWdxqrjXMQRLIqd5Mv6Xt+PuhAP5nVxljyuAW
aZdukhC7JG3uWHqm0n4AUwHCjvnt5Hnlh1cIRsPJsMgPkSrg1PM20Ow9Qp8sM/RD
XVx9FOpEdJuL8tAnOl6tLVIqiwAQspMN2+EF7mJJ6x/3jDL+OUs0EwmO4i22O1bf
29MthcLUMThsrbvf4fCeLa1cIXnPYQbTWdm3lQKs8V79nqCkvRtTF4ie4BBRcT43
qABoLp7bP/29+ifYyVPvogbA/YlYhWhAeGjXQLxcKSqwzxcXaoLvH8q17K3oa32k
r6+1r/qoAIswiq+sgYKo01tvur8ha35LhxJz3aQUzlVIueoO+dIlLhIJG5Z7/+no
aEiY1sXQH8pIVcOD0mNA6NSJSrVsUxBq1GdShtFN+njPyAdBad9zkQMru/JdT/S9
VBDbOX5tIYe2du4ixxWYBE3+QZyQubn3ZXXwljAIvgq6wArIX4ou4ExP5EBegM7+
WecJdvPq+S48Jj7J9vCuwMkLIpmoUfDBWCFBLXalmAqzn7h8XI8U0uW2lBjQmujV
18kaLFEJEDSALoPLciPwk2OQFxgTaFx7Y0yKF6H3WLwVxWWkpc4Xo6Ia6IrD84VH
T66CglRN6Lh/HqC6JSKKJRygBWfbt3leZpqxhC28Kgpt0YhfqWIgBtd8vFX52xvf
KJlDDTMO8yGUdGTu8hGaYeEkSAgxz7204DvKSRwjxYtdh9D0j+ajreHzkTxjiicD
pfaFVhwTyk+E/vMT//VhllGqePvtrUTHqtkTU87ttMgLc9+6kFwLLBrNfrqNXn2K
lomYYGhZ6/ij+fHedsRo4O+9ysiyJaGQpbYSFssXkQj/qCKp4yP8QtiH25A8N1Is
yR20sE9SPoW3fwAVqukt1W/i+jANEBlUvLj3q7L1e1gegy6oeEyjylNf/7XKjAaY
SS4J4R6PqsNtKggKYdvxDCQxuI/BTnz+pMbgDTSUHS6rLTTWvP5bd1m4MuFbHcXG
HvOWrwkL0NFXu8bKQn0IvJ0p9JokbIMc+ASPXNlbJRxdSB8HzfKRHtX+fMHsjtT7
KsFgEP1GCsEjUgMYYa8C8fUOzRYtZsabgok9G0EQUgF1rs511+4DeGTB5xQp+ZjL
CDAH+arMxTYa5q3IGHBQogRCTyab6Aogd2ClUwj32TPPd2w/Eg56A66hNJ/QqeaG
QQT5NO8bsTaQvZElDucWWsjRn/vrPnJ0ySjkl6/jfJacJOfM0wutKhanAFGOg9ww
tlkuf9kZ3PtElHBUozzgIZ/X2Uru02/8tP6bswAIdt7ld43WbrQqXJPxUT8J5my4
6/nNvXZDMbqVM3Fzwd8m1Q0CAVxjpSc0krSf0rOqoWbPzPMECHjy7ITL5rQ4qE4R
WILbVtx0X6TprZ8/FV0Gn5jnFJMqKU3XZuGvrM0/AJvwI7zOL8rGV7O0KKjetwsF
Vxm6a4jmBQ0BAPsqIQajxRJCS/JdS0qtRC3k10lTnCMpNBjwGyObajBGMKXa83PG
RywC9mglURtDR+EcxoHi5EBOwbAk64bzFszJBR3NinT5BeutDyjBs/fA3SCmpIlz
2Ed9kgU5UenNhxFOQDFeePNwLqREapS02nJOLh3eswRY9cn+UNrXiGzlEX7ARnOd
ee4DueyJUFwbK1ss3Bf5/jVCI51YhUarCakUot3Vh14fTMvrjPqXxRg/9ANcGCGS
7z4t6GBuNUA2HKJmXde91t++RH2snKCIPXmwbc2U83Mbt/s+3iosyKl//EzMBMnp
tb3w+ypWEBxjydVRYOhzuj87yVk+A3x3KqpVE2QA9VmpFYOfltgjTP7P8YfsEdyJ
30Fnr2db9li0JfssbLub4P7s8+E3y8pq96TrqdteWycbdeAhH6DS0Z12y3TUVCBo
rZFze//Mf8meZ4mAsKi7lIMX2gyoSFY+JZC/K9T6NzrRHzNJ2iG8E2UTVEtFxUFI
9kDuLPuSBgSfsLdOY+y40GfABZaSQjLXpP3R121ZnX4a7bhC77htPllDGbsm7fKq
TzQHWK2nCDtRo+iAbzYF+Z3UAAkIwVsU4G14B/3q44s+t5CSx3FgbAR6Ysp2gnDh
xYQTdm7t1pLz8PbdnYTpUqipo0kNsdyywYrU+XKSTwomlW6tseT/E20wBMR6rrqz
aa/pj4rRY61rs8Gp+afWbFOtI5SgrlVY65Iymoc+6AelIAIZ09j8kL6efQim85Wv
+zB4euew87CuyPw+To5ZQIU9hLoxYE9JtPGAeqbw5pZ2J5fGecML+VuVkTdOYa0a
HrVBvKQW9Q04Abw7IY9dhCs1Lvs9569YhJkMteiYsTPOwrHH+2slE2VuK6M4XH3L
icl8KZmvs319ldFs5foUzQcxzwtMC3lXHty57rtFwdKpDUvTGOaOJyUGiEPqAQw4
dmYN74Lnqz8/Bo4ZWx7koV8+p2pbFi8xueTMVORZ0EOjhkfqHpdudDyPyMQF3Yvx
DFt84ATBTjfNUWxQsbHRN8pmZgT9bMIj33vTi9aIelHsh+D76m+peFlwBrr1POqx
tXN2iX1ARXa5XX7CzrWHFte4Hvtsze2NcMd1fPkrCLYCRLhoJhPn5n4POxhTKiq1
fgqWGXnmaNc4k4Cba3R4ZMSt+j03oEDJfkZPCI8I5epC+SNLTggZOdMspU5/5Ez3
w0bSX0bbXJ6QvvT1Acw2i4vNnNt0JRKekoTOEKf8DW9OjamyeIdooDuFQav4ZRlw
8ZuQ8Snmc+a63RMlqCcyskmG6uz+qHAxJfwpXoY5Mlme+3/xgy2GLducpxTy5Bgc
HZaWQSVf2S3dZyWhPZt7SYsL7kvIE98H4Zs5BweotFNdSEXaVN3JMDsGfmAWCeNZ
xS/r3XIaTLOjxIAADml+Yvd7PbMSMfaR2xDXo7cjJKYtC2PdqNYYPmu5yP6+G736
FEkm7qfgchTngSH63zehOlsdJZc4FR0CtKpJ+wFRRD+HRidRamC1hepnYH1mfea9
Ks/2wxLwbCbN6cgUhDhzQN75b8Sgul976I+ri8eLlNMIyr0gzZdtSAPPSlwUc9mG
KU8AkRCq+OCoNRciXWrIibfUFsZFPRQ/wBlRE7YUORbfC71PQJYW9cHDUgwkndc6
VJymvuZPCk2mErgtjKjwB52FJuaogSpvh569QZDqRacxfn1U3egG3DyE4SvAaeIU
5p/tc5dYUSsvTj8aWdEOt8TthPwJhcZidzKo7qXylesmCFh59cc6PxxBu/JzEnXB
SYM5naIEAAbt8xcqeyo7dYKdLyWqXtPB2eHeCwUwMqdWSzlESv38qJNEDToHs4/q
8SkvhCh4wRG/Xb4f2u/pSO0woXSjA0KXAKS8qpRBgmqox2YTHkWvs+fhmN1OCBTe
gian/6HHZ3/Z17PXCdUUlVFv8gmke679vbAz8XnkB2E2QJ8DqV4zi9SozurT2F/S
9NYhLAJPXVXeTjwSKvkqDhU4jHgY7C5HMSjookGuCEVqFE2//mNGYYosCe9QXmFQ
pOy+hh1xeO0XRUuJhh94LpSSTSJLutpydZm9pT7gPHVAeLcYZ4JaVYuhEPzHCHBs
5LTxHdIFNkC3TrwA99kUxT9G9n/2mCGU5xValjBvpl2+/KSUVLH9/TMAVDTqDTk+
lh3A61mvRaUEeUSJ8YDbG1pOthWmE4/3A/xh5gSowbfR6SAUfXV2fYILUhedmAjR
LFfzAcAwzoJQf82PnOfOH+M215aATju140B9b7gtFHpY4rcU6J2W0f8etu3vA+dE
sSQ7Dy18wEyiH1ItJKrrIU2zkN3XSdTczHSCWcXjaxHiqqs1bZ6ShhQ0H2Hv2Ii7
dfRaCP45Ebe2Q9ioL0rcnz13nEFlRfwMg4gq5z0fM1MzHN4giwH44WTpIl0Dkh5Q
N34uLiVy6NGLVWFmE45l+S+WvOle71fzmLP8R8F2ct0QtsiKr8ZJjbz5qHTptsgB
QgWdBwGwc41hY+gKKHGo+LXlDaACyS0iWIiF3VzJip1XgWxdGgK39wRxqWWiDHxN
kw5wudlzmusf4VbbujXguhDg6d2iR1LRYbzH+H1yAsqjHdrcLLBpry+hcl8+2WJL
T+UNRr+mOk+gbFI/5LnfIhTHlydbRWVVKszT7QeizBp79dDguf2Acu0fr5UELSNc
T6aKszoO9ZGobuC9PrrbstFNkpQuZc9Lf/yuNvKQJNujvuRt9tCDzr9WBAwrdfX/
Z1sLWNzrbFIZR102pCYbvQT8Vbt92FWOpIs134jlsCYw5eZUJCBfHEn0b24vUUbd
IyjAKvJweo+HIgxnbO4ZiRKn2fM8j+U4u43XCrsBw/Kn8cVTZOnyOu1Dx6AaCowM
MWKXg0zckfvbJnd8Y4xqKdORKOiTNfDWKoADIqOoeaRtgbzg36hOgUKeqZrmhuYJ
Rinc2HhXtl5CnBodqZs82On9gVx8kx55f8Rb0/Vv7PUupWXYOlbJzH+fJC5kDIiZ
gfQwaCDD1O7BbRmJnwNtdBf5eiZBKV61o+fJuN+oq/WC1XvRmzmV17melb8S+qvL
uuZYKXwZUZynJ4jLDug/vn5OVvuRNPY6CbLEwDqn9tdrFHRi1d1ltZy3WYeSH58g
jMhRJIds7HEeR4GSKKNVrS1NU1B0y8b8cKaeqJvnk7jXOqV6FzI5P0FvBEoWh5Qn
/e96b0P3GogKY5ZSfBYhbKWr5uorDsRpIUsUP8XDQyX6nrrN+Cs+rZ51TfZtKGqF
AJG2G3hl3qR8tum12XvtITvjXhhriuuyCz6FLWKhA+UI63sGHt8pygLP219Oxim+
yvs4oOdaKAWh7J2WFAPOrm8ZUc3qdAIVbfCNo4AHqCRACKrrwaXJMEO1UgFs/vpV
LA6oOtLhf6bPyJkG8N8DHLKVYpr92gde2JKA43MxN6qVpVqC5+cL3wWe0sf8lV5M
0kIL3Xdlf2lWy0hlhbG9Y27joifR7rlH0toSTY+SG0ChO/EbZkRH4eT6ylMno8+P
0/NEVj/NVnpkukCGMD/Mh7psErzGIsAiBSQtEKWnLpDbTwQ9p8EeAJOON43xRBxs
Ob1Vn4ELL86B1nUWKu6jeY8qWjP5V9Zx3cKekTq8+ZTNwg7lCrhoph5VnjcsG2D6
XEXWVRmLwUtkFFU3ukmfYlZVyKiq7yX6zuGUxtcFvUZ8Mr62xcE7I9aJ1Kf7O5Uo
jd5Ux7TNrVDznZVo5ddVZ/DQlwjDFB5l4CFHHKZbNLfZweZj1f1Kv2eVJ0EWYRM7
5HNyjxuw8OWjbRmkvjCYM+0oLtvh4y5ebRDReewgUHOGZfr2zB+MlpKfdZNb7J1e
0AfZeRgbjrOlEX/bKnsZ5nqyEBM4CJueaJvZCEjFIyggbGG3xQDBJb9HizS4vg/S
kG5qmPGT8XDBnnOjwzySi9yKBA3kL1EBbBG5zRGuPe5/4VRJHf6mIa0rhfnliHuq
dVgTskp8M7EMy4NE5osnQ4gCFO36nGxAeno+TzRvV/idjtl/0iq5CFkDEz1pXRBN
0bF30BrUkMAG3OuMEys3htec+tByWJUXE8X8rke3kCmjngvdiA89QMcT97Bw+1Bj
6UnOMrX+/JV19ZcieNyeVLnlO+aptH1LM1ivGpgpnlDg+/HFpf5KupXEWB6B/6PF
quWZ2H7VOxluFTneYZ85pxtcTN0NBfthvrlWbZwnBfBvZvPObTpefHKcgE8dFepz
xPFqIPjRjH68/vfN++qASQHXylJvojUJRcpNDtiyWc9YLxB91VUhteriyP+XzWxZ
51oDOoGCvtGw77PHPRNB7xc/57ZuIsmKhbc04R3IUSLfhf2gDG+lnaoWfb/aoGp9
braONUAHhKurMemTXXZpS5akdmptLkkRJ/upRVVjtOjAt8YqRdMzdgzIsNwoqNkS
ZHhAxgGGt/8S9g1crbDC9XrDhasi0Uwl/PG3s16ykY5bDoTTsbQCPcJykkJvCl4m
bAAFnun0DOznI0Qjv+HNc/uzUp0douIwGQ5RBBfAIebxYy67/1GeRW8bTBdP7ueU
WMTR5s0OVeS0D6Waz4711Gylk+bPf+lEHXdeU9q8SxL/ZaCzskxpUa5qXDF/uwkF
y11ftdHmq6aDBCizDIUWz1ztG6PoP/+5lR5aozFFoRP7JDh68nw+/SO4oedV5o3M
+ccUiPIgbUtIFnIkUwAcxEOieauTbAei0a1LEDLNGmxEDhaNNxL8rOG2znEIlZNZ
ON4D8UJxyXAVvWToipeavok++1wpeexqL26V03CLnqCGTznE6v981hHZfsjg1LKC
nGYhTDBTIzPwVlEYcaYj3jNWhyI6IYWM+qlM+JmjeFHMxrSaIz/l7VbPvIydmUro
HUpRn3vUehWn+u6F+e+oj+HCmAiQbAJpGKcbC43G6EHjBhXtLgk0FkY8fQCK9pmK
HXfhn8q+CJyy8WqaiR1jGJ8PCJ3XO2EVrBMSrj8STBFiLMImfy0eplLA8O2CJfa1
hwMJvGj7XV2+xRZhsqDw5rQloaj2YFSmDGmCP6ReaJB+BXkQKhxx4b5DicXAbPi8
oQTr9PxKLOcyzdrvfzgnNvLx+200GOUMzp2aVhnF73d9kTvWEQAf+Yr7KmHtLGby
vBIjo7r5haTlZOxnMO+w5Gqjn+U3Z8f3Ek2GIJAYfegQVVj9n6HUKE8sIBWjIp6i
UEcb22Ws76CjeDVsO3bI/OwX+ThlSEg2gJbKjHuJxFSSKjmTVF/rydzaeoF7DyU7
/VDUY3CPthdLy0cigvLhAdhj1jDwg1FmJ+qkIn/aqXXpF49IZ7dQrocfrMiLXmzQ
jWhpNY7VvICCY2RyH4ROzc4bPK96/MiDcgWOrOVbJXAdQIPSqeT8sU+tdTS4Rtl7
1aRxD47qNODnAW977yzsHtvXZoWyPPpBQEjq7T/MBguc670POeor9tvqH3iXWGIc
PuUaOsMbz+svJGRI2EJ/sYCWcIHNkWe3c5mwV5zncne8nuB9PhxT8OgNWTLLMSdy
/DA04r7SNhSTwUJxgNfqJS4bDjG87ki9odyBQBolzs2Cy2jYtO4XPQzYzMb/bB8G
DCNAHbM6xW/G8l3asmxNMKAE4mWHCa6X1JbAaXaSR2BAGGPm5cMUJVhpgm34Q5cH
x5bVtCuI/wnjzVospGF3npZqnbkJejOzc8hYTVG3K0fr+5rYNbwXH9tviDjx+MHk
nvU0/LgIBTRSoAheb8TRtFRC7s116j3HbNnjbkyNUIxc8FSIuDYLSW54V1yr2/e2
TAbG3DoJIBPnZNv7KIDddnnxKIDexrA9x7JQS9fnMG8orAKMit5lxOaMdPbUE1On
w2lri8fUuGUL2nKyYIOSVYl+2OtnxrKaDYCHXEFxLHDRyuU9E5nunIge5sgZd7wj
HTg4y8peJGSw2oFnKBLL2gAEQ1iFo/d/2N160GUhWA5z2pNaPfuvKt36HSvNq5OV
wxOFBdZguf5tzeOVc/PUx8zraKxN6jESBbJXya4MzCBVdS6hCaLHEUurPDRHPstV
qUWhPom0PRoDFOnwFgOTgiJSIJuHj9uy1b8YMaoORfFXzQfN7qP/0CDBEJJ6RArx
urYmIHIU7VMDswUdQUwQcEn4UNJ013vQY52FKelm9LAQGyrRs1clhWX7UuGKZHyj
EqkjAOSdrMSL5MYtxlapUeeZBQ21xEsVGM/qgyhTyRNU3bjv/UcuKL10Qx9AYw1O
gSFBPSSChOTL/2Wip2LWOU7nStda7xws2U5yabdzlN0kmu03k6WDCc0yxLVlImbc
8q6hBjEG3VZe5NI1GrIPyOxyfsbCe/i00+FSwqLP2/JL44z9ENnJmRZTuo6jI3jN
EJVBQnO1k+VukHZsJ/uyc0i/HUQaLZJLODFIpQZEakCq9BOzc7GEkUI7LE7XrszI
Y+PjKIAc+2m1MnMjOqr1zG8drHe/abrEIcQVsAxV8GISxMyl9uSbsWfYAYGzBKlo
HRFOp5S+vX34Z12NhI/yYpueEhWGRijuwL5TaJJMtjSSs7WE2Cf6QX5DtaT5N21t
VILxsVp5oNOhC8wgD7gmmyR22CiZazJtals3WA/vq562by1cQfKrQ8thGHdYLo7M
I1FTIo1jWhkzioKecBA1hqHTkYIkShCfu0iQF6kCHlUY6Gv7hVTO4ZABQxwIFHCd
HTWIRrfJ2r38PG1B1ychTpzIcV/sITzPEYMGrzgYjKllYXDYn8CI2NfuqPuIPDvF
hPX7uEg2nYW9OUGQ9UXL7qv45xjgZhTH8gzHBJQzQ9x5G0HldmpguCIHN0F8RMDo
lD8N3/bBzAEAS6CHDFHtwL+gL8EOwVtHBYn/bGN5clRV2AS8d/Ei9v/weIF6tQmY
h71VtPr0lRKIy2GzCs8kGjvkHbmIahYvWwrBKtYRRLwPh3zhBYFD3HzCQn97AKCq
5QChw7hwO7W4OC65g/vr2SlSzLAjug7pzEV69Atc7U1cYxJKGZiQRYSuZ1SnhVaM
NjG4PlEDWtWtjXu5a5bIMNWh7m2saS2t1tTzeqCzOE+l0cuqHFmbOFaxlGHYEy4k
fBgxXPN4zO+gYHDk3lXBZJy7QP3lFxjkVi4J05t8WE4r06lPRHmtBPod5yXC7nMu
hboLz6RTlvMjou1ubp4+PbvEhmUUVPgqRqvt7I1pnMu7i/y0b/AOG0wlpdejahNJ
2dbyHXdx/VzS3tmHLjCC2vV90uqzLC4wf+Mcdt+3iZtR2/4HreyzvD/BjwUxCo5M
20dfhm8Fx0boEXWDvwe+oiWh4frs2+L5ed/DbVXk0XG8kqQqwU483GstPwG0aoFa
1SFs8BZA73oNMcumHLIPWWIzoDQZShBeKCZwwNsbWB9rQ5uqr4PZXHDeT48DdUz9
dvAyfPg8jU8ST8QE8JWl8ZxxGgcQyRWHl6WgFEiaQWjKjyG+fMHwc1bXRrcSAvzv
kYgeb8CsMVu13VhifWkWSrB/2X3qaMLh4sH8pQtHd05U85rDJmL0wVwg4ArV8+cn
bSguztoy4OzVYEGMZ2i+lrNghrroMWokG/63RamwLjiOvOWk46b41+A5l7OqXILO
PbX9u+2h/MO9bb34tXw3ZUGGptqPwsBO6e7CZiZCLFssFKGfNNntIjBPifScz8kw
pvbKXetn3mqPsEICtb+QFobhr7wWwBa55gpfhaemFuVVXsrbwyHVENePWHRB42jw
wSAU/yTXzqUW/CH0ZtDc9mhzpiQ3R4BRBmwS1yyb7QPyaK2urLO4IliJXe5Dg1+Y
4X1/FTQ9USO39tnTJFWd7YzoAT5iBi14Icev6A5mq9ix3uTJRCNmaMx24fwjpzB+
WaqbtKex/SRHbHSB4yB40FHRopdT3t3y5TyHuN20HvzGuWa5v2XHkaId/h/5tYrg
zT1dCPIPnFN/h3VhxhX81ARaWV29uphDOGtNEOeBfCQzwS2/gfGOKOGxZW4RaFjm
UvyNUz5sE3Wkw9jeY+oQCDhr43V6Rd3XIfyI573a65rQwdwu+/HbukyZ9WRl6mjR
PC1Z8voD3PdFJVnCjozA+ue//QPdMo6YD+qXOC7JKNI/TzNJLaADojSZVb2e1M/E
f8PiNn6QtMwU3kx1uFnNQBRjIlfWlZQtlU7v+C1dReGgQT496L2RoK6SmTNDuu/z
KOAeYqusdsTLc/S8esZoPultdGMi8PJynxp3//oJeFgkcBcEs0eqsf9I48q/hqda
4HqkQ4SRvtUu1PHpP80JUi3Qxg1HwDQhy08pyYtCU/72MbpBtTiNTAvhcc6cHbQq
ToZBpo4S51rq5c0IYROshe9K41EhFnr/ov20nsnXdtgj2PTCwHiZcLtiroyUKUtE
VbrO9I9JUDwtqATUZJKcjjWHnvy5psYKe7tcNCphpthH23sV89MZ5GslWvS/2yoM
Cgg2oaqwo4PQ+BWYgg1n53H7SCiqCy1jUnfGSOPA4x7jRg+wCv1oF3AO6cjXrPAA
G+yTgbuFX4OMGBiCDYYS15Tjp/NmmiwkluXB/4w7Lcj/iTWOtgIhFsN+7d9Xnx5R
xcv76KT8bmPVhJY55XGayhHEB1GyzuBs5sm9WVVMDYGj2xxNJmHdcfuIOyFKzAry
ANyPO1EmfHuDHQeFNjz3NxXCqawptSTDjqSp6+ouyjF23BCgT7WJsvzacWcZoofa
HCbpnIJhBgDpjjH/QPzfRCKVVJpbvpZz5rXariHLgmg1u1/xrsKu3j4GSEkWxNaZ
Gxv3/iePHMph2UoXJmBHq1l8pD//z1SMbfjaTIzLkSX1k8ll/n3OMI4If1PfjQSJ
7GUkFUZNXlDYwtlOa9soLrD+BlpACw2chy3gCwPLtdq+zy2WdaETxuT+PVCDKuKE
DvE7nmI75PhtIHnebErlwXm4OcJ3S/7mqvFU97/mLUQJfocHPgs2UPXUsiua/7Cz
6C5rC6LYdLhAo/+uRkfLYXjx3gmiZCleIR8XIfQ9sFP863AspPnd2gH5Aogeb39o
lsDRyyF0SrxsCCAShum8J1PZcDNFuxL6FbQJiLAnf4ricU87e1cA1GXpJgox/66c
i3zps2IGVhouFqSL/JwGIguTC1XcfyhHlOTnXCu2voFxPpm7VPb0CSPwrU/77A8/
g9utPc8t5ppPtYABNE8gT9eH8k75ESlmVfS/Zt/rjWXIQdfHbixFUFaHxPjmOdYO
Hb/IjEZWblNsSuLGRH3sqgETvRMjN/iR/i6Weg8uLDIeUHQxrZdH5ki0XVBE8qd+
hkkS9PFCoZdcaKDJnHUYDFboZOn4129tVbC9Cs2fMh/dpvNMQGTG3Fs+96i4QIHU
z7ud6ltqxzRwtGr8OQhHAJmB2BoTrm5IdoFmCd41SX1y6LLsDoBcuH8bQMXVWLa3
HxnWxY+mkSZqJNapjB3JFWOyGhSy+GLhiHrDHmGoDbxX008rTIr4IaMkEhcnLlWP
2t5+DRiSjpqN/pRXSeHiza2IrmaSTdFlcJyacoN3yNv0BaLwp23XMiOai91e6ohF
eG0t1Hd7RzXYmD4n9iOq5etgoHYfr6AWXaYf+nC6EX4O+EGJRz/nEBxUUXQh0dJC
cKfKj4DVRh/ZS/tR9iKH5IW9Fet0dI8w8qClq2yCLEZ4Hm56zRXpVnNR/S02dAs8
0coiK3r+DrPA+2M27xvNrf3oiCxCKbgcsaShryjGBgXe/5pof3+HCpp5sXEFc3k0
c+ieRHpq+G9qNSFfXiwwnG6Whwlm8Ju7Kkrc+oaLZLr4KQuOiQAWBTTH34Tn0yaj
GIgzGowa7/bs0JjPKyZh1RuEklFhnYNEA59gitd0uXx+mSJpBDdeE5RgPR6Mhm9i
GhJJ4KRBc+XUCNLUDMEX1O0tkTuwPho/lKWuqYaOl+7j7RIvyAB4uSWgzWg+an3e
tYLtPLBUCIqqaaNFPUDkKp03wS1RQDh8MHn7O1WM4kpVSPW+ASNVMUKKbWAqAckv
WVm+7GgzNsvuqK4hJ8oswPyHS4GGL4dey+yisvZOJZSZSNnZPEBntV7AsBwM2cvS
/FbcayV3RGA2lEPoYt9S/D4pL77c7o470cmG2RbDq8LQCnTRLjgvfA6qkI/rsVXC
NWGUID1s9IHyu7XlWLIrhAzsxofKZ7zDGtJv+QWQQYE+8nWxBhZ/s/Jurvp2/u0M
lLWPBQDHO2gNyYN378RgBBqRxePkD0ebJtw/omL4dib0tHW7EPmcrssp0qJT+Lna
xAqntET7uWcz2HQdt+M3NP1YxNE9acThKTYftG6hibqvkXWiavzxyAYRLm9K6M5w
LZwKYbqz7yrFr6LTJunUgjNUsxtn5Ea3facxMEsGbVrdQOQBYDK4J5JU+ssmJJEc
I67An46xK7oKOyXI01p2RKoduhHUuvMzzx26AmWbhpt8pVyt9hzKif6sXMyPxfxe
6EDlTKA4NrmHb+e1GZ0qqhFz7zRp59uuawm4kO4Ae45mn6CJf/v1OdNxMXrDmoM3
1KzE7SzZ+qvXx5K2KnC0sAJjFKrhT4D7etQoposuN1GTqINodm9IOcYLlk5EJ8x1
t9j5nY0NzWirtbFxXCp+gqCG4m3Cz7baP2xMzcK5ZhfjlEeo/7VmWRqXFz9Mgx3a
oPfjqMnj6X15Krb3QpUnyuRPrO4Qo4l/tlEkT7dlV1PW3QGjH4lG27MZqdkDjbpq
LX+gukFFhW+rakiXqXiW9l7xRDy56d9aaXSKLGwwib3i/N0Zzc3nY41Z96xxKdYU
qioTrz1wxOU4f4Hlk/8nYa2DE48Xmvc7ke64REJZKBpiMmV9PFnAsnYgu3ydEkwL
rKKYNkY5FPYh1W1yqjyTjoYxAZ+jXKirxwCvTf3NCV/GNq/LlPfFvzcRR9KqgnbA
wPNBJF8AtmLsSQdUnhaBVcirqpZ6nir3K/OVZ0bxwYUpx7AnZZmi92nIYJC0PvVz
u9w7+sex/Xa3N/tE3IlB64RCy1xggiQG0t35BTNuYvhAfDpjr7HFS79lL2ZNWFXO
SXFuEHKWbGHPR4g22Z92mV1Q9F8RJUPi6gv3jMvbPO8kPjDfkJY9/MIIKJI/9DG+
45GkaHnBxqf8IiOxDMgCSpRUoBDxbOyKr3QlXsz/g1DDxUVBOwkt9bUFldfFa7le
95ioKsO+wQn95qkNKzBV1Hm3huRL5ZdeHFiwPn/Udm6Y7qUH7Q1WUjDlKWYXOLsw
oAyTp8ZVFX+8SBIYTXLzxEhxf/ELrlD3BwqlI+gyclr+hpEWK4q3ueMnGndppI3N
XcFbe8sqoW+E0CPmOauXx6TkyeOpkwzLeYyXyPmTg1c9yYC5LSpZYNGyv348RFGN
OowKZyf8vI1ACSohMmKFUItc+99/lotEvQkm2FEfclml+7y5p9ybVBpvwc6p55gG
Y/lnRpKhlMMLTuaHotBb2Ggoapqr9VxyJAr8piAAD1ZQfaRb9y8kZ01VWt8dsSSm
OJ+8+Kj4kNv+zXeViseMvC7Oh5aGhB3jLgV3pSr2ydiNrlXgEd1WiVeBLfzoZEIb
R+V9xVDT89clspnWJlDqvQffc+0ITTV53ukwFP5uIfuS2hy9UdFa6lx53Fh2EB4W
B+oE+Pg0o0HZ9Wh+ofc046f2unDA+SJ1XfJOVxWQNkTmGx7mkvStuo/H+XZCR+uP
buvHIJmINJcfr4X9KJywKcrubmo2E6jnpggY3rWtPK9vPjXsQkQgmm3TL0Brkd4X
a2pARJBP4RRuyJ0O5gQ99m4OzDr/+meCXp9ccL5GN6gifYxelAsJcbAtj6PX6efA
ca8Kjasrc+onFacsxOOST63g5wI7MZSVy7EQQV+yu/C08uyLiP0Ml3bChto28fNZ
+vs9vY5foO+vKCgSZpBZKjSJXv5j34gFbLvEa8J3vrkeuroZePndfzE7TWh1vURX
jBdrWUZBJZ27OfOEmQ5XJGIcq5R4364C0kqH30AI6ParuTRUF7c+8I/yCf8biO9b
0yQfteWJiP7mqz6J28uTq1XAjws5DtE3g3YMjzvnduZTrQK4/QKwAlqBXg4zexbA
Sz6wo+FQAoEedsTt2AYd/+kJdAXXVxVDA5dFXpc5jjiQGX/Y3lezY/QDA+zqigku
ngQ1ud12xsfKQzXmHwudv6lr4W0akGoYf83i46NmxtH9MVd+E3oeHP/CyCJE6TNc
sGY3701lq/67mXB3KlFLt762ZT1q4Wi6/k6hOuQlEAqIrjo4YC+KO1jnHAvZixTG
sr/T/TnAMzDAZOolnOftzK+BhvRU05rZLupYn+pmCvUqmBZ+y58jU28xZbdMtarb
DHxVZQq0FdrtEVcScKmdJl9dQa9CMhs55laVjJe+8e2pYtHLeP8RChUadI6n3ohQ
pLRvh7jKzKqgolMBxSAmBNZ4LmvcSNxwLXm6sRGJkW+tgAPaxE8wOQVvDcf9x8o6
XBIeONBulQ/ntAOvDbrmSAnQHZUNe3DakQOupy8nin6mwVbJwz7AvP2wD1xx0et+
k4EAZ3xZxDm/g11aDTXX2T9f+k90QgLgGxsx+9hxeLobIioMdRSEudI8MkkbKMkz
IEeqD/XOqN9RhZSiFPddANhVN/AVP/bTlSohPaewWZSHVHqy8Z13PEN7YThbgprN
5yNH156HmAFtgYUIyyiTNJbYd2xi9FZA4AJ1l2x7A+FaWC8yfg0U9Ousxm/8gV3v
kd3qECTZrW2FAk7bhqBVhM74vwqekzt9rrIak/utQHgkC1/+LJPXJ2xwwVKo6mMt
7Lom5se56rN+fqkVm+fj5d4EhRd/RCwKWNwe2is1BaN+gUSm2jpk5Dm4FVVwkCxs
Ezz2j5QYBT2MrMZK6pYDgz+5e0myC36o1nnszdByYoFyvjMVt/rylEJz4xr/2rWs
X6T9ruTfJNoexd6pNy36TmJoVq/XD15QdamNc/PtNnsRWqjWC8h88P6D0uIxRjP7
whB7hUEzyIzGqx/pSUQp5+Uam6LwBY4nyiC+/bpygClt7wFV1O5dhX8R6sNAKreS
lE/Iz9nROfd0DlfrPbUE6XT1lLXPRazMWtmAsKZy9LPwt8CHXw08dYraEGUjiOEt
JAPsXEtfbIU5963n/plPm/tVkyK+zhKz9S7bLl6SPK1SdkrRuyQY5C6+jGc/9T+x
Yy5U9N3Kyaj7i0M6j+IqWwwYlt5WzPTjwzmLRFVn0MLjBk/ALVi5W2nfmetEj7H2
T5egKkKcETYPAVPsoLNmMf95nqE41CKQxvQycbVtfisaRqjEKS4Ub+Ky5+0FGJer
By0FKtq56gPnoFhBdwHIdx59osukR0O1cjTWozkMLxaFL9UqUQz0Favk4dwLZEN5
8PUM1K1DeCdssH78SrY/DUX9JQBdieHK72H0xMTMwziwxgNaq9tHT74hAJ1sxfea
c3VRMwEkvhJNoYklvRSHinf9p5cZ0BwBuMAFCYAAtwTDYzoOfUoKPT+GpLgEWBL3
iyZb9Q0TeU8U/JCTm3NqyOA05QhYH++f6owml/oMb7fl3kY3nKfthIlDpSJUOhxS
6EsvinsFfMKb79t70bnohUJ8w0F7vAT7MJxwBnkQphR09RLRR3XplhodAjEkDmDL
RUJv/wqNIidT0L8zYTtSb94fkYpQ5IKavaAKpyOsiwkJ6NGRuODHo0MbTUBUYDWY
Mr/Mcd6+NQGC/UZrSlSw8HwyMZhLQq256VX0XsCcKZJ+YTB6034PRPSb1IsZfO/X
KiODLldUsoRafSjSU3JbDdH4dRabkv+lr1vSeI8TYaxLg10gaIw3Io+LeSWgGSTA
Da59BUtQq1NlblZc5lQ9+0HGyneSByecEYusjtNVxJpcodB7CtVg1jLqiZQj52JL
RZo0izFw2nV4WaMjxe5SFe3LINc3bgbArSMJyWDxnC+1YF8BHtmrsggLFw7Epem0
A3N7ZA08yv5bQCe4RntVmuH9s1nEk2KiEvxV1alUpnVRPfvu1RXPZt05ZSaogKaF
HOoiS6197Tk7sCNi66XrR0EeuMua91YHeyP3qlYrMMDGqcHUaSwEf1AuQNF6FxR/
qf08vHzgf80HGscbFgUbe0vFbvge130sozxFb9Sj6VADkaI7GaaJfbWsS+zaVu7o
ZVcWheLEeVcliSV31qYIAXx9AWF7kbrdJ15Y5bXChNLOQPyKMSesYKrKVSDUTj9X
B24V+0VCvm4ugUoaeLAM+Uv7q2wIdTkiuHX+owob0AS3Mimycl/KlB5re3ZzcCJY
aoYBXpnq4spf+DMK5D3mdZdqD5UsvZsrAGf+xPuhVn6Y8JrfPjbPc6RWwDS/PG1w
ai8JZ8lWeNNCekNB5Jkv3fRUFbCH5xDWpV3CM3f+/3BTXvkxg46NjojFVmnaFhxU
HkNFQQ2LI//74m+jmNABc79duDcvNH15QY3eYR3G9f9umc0ZtwXnLo4dujkK60/J
bOsIVjJiRpmC/6ejizj3FhgIQU/NGgzCYIRRlEWEPMRfEgnKJgBeXxfLQqJWWT3+
rtHchrH2sgEBIuIEvm+AOq6f4dc5mCs6Fbe+mTfTuyprI/SbTT5HTi0sWiDm4i5N
9CoyJCobaf7JRkYn5hReQn9b45ixOEay2lGocBIrnsYsrvo+rNiVyQTXoAL954V/
7j8xxOR+KbogMB08ksSOj7s4dYI8zQ1RQsRntMdgeNeDQHg1VDg145FQsKQcDXrx
Xnu2Qi6IFhAo46qmw0YxBeMmNSAjn730nDY15ts9lenDDxbjP6xqXlBY/WsR4IO1
fR3ru8zFijrJeCwqbJA1N4Hd1OGhGR2b4zjrBlSl1d4YpZxXk3LsKyV0EKGofAef
SNAGZQQN3XZQxgsLvbIQvRerQzHyt9JmxLIag93dfao6o7a8PKhbJ4FQYpJBitXC
pQ+3Dy6aLXrT9vtFYGk6RpX0UX8RTWupee7/JU/VmQLouOcKeu78CDA4FdrPBC1B
BFOFtp+ezEsFi8OjXGeGfLWRI+9sD12h9+RMjwqQLXgzAtdAvSk+RQnCdbFQnbwF
Rgn7NHjBeGHw33HQBdzK/H424oRy18wxSZdlFVUwbXTi3rhIT8ezlLCcozRxevuy
H+UBOdVIMo6PLgYmjlmct7CzuC0R4Jj/91ZpL9hG6AZk6wpBvWNMAMyV33eEMU5Y
n3j/1ZUn/tMjoCKPiBlQXJrIVRz3EB7aZkzwHX1+o2+O7UeiVkqW3Kp2cNhJfahY
OWr9fewouDULEJkwjCcHtgZgU4McLscBD+YM+O4Fau0Ont4hXyrk3pNOxphiMfrX
a+qmp7rvw7abNdu0e1EYce1gW29f/2TRRsQyP7nAFHBQRPXtkcklD4Iq6TWR9bQe
EbEnlJdKUQBYA6JptDRXuG2qHRExLBwPJv28Zm7dZX+5cscAsAdWqcEbGTvNUbBG
drhQ9PFPHzYkcamVwx4nRvAwKbm2MnJEk2qfzJi7rQHX+xxTGM0s1g/meFmFyJe2
/PswlrteYNAXi/P3r6y/TU2fYbjEeGMAz1bE90QewYG7eURtgbXxsKtZgfTHg60I
aEElDL0fXScB2dK5pX/GjlAP7pjC4slhsMH2G0toFlZRRS89sNAdo5PwS5cUz0NC
KQwP+IG2PYJxhK2bu/8zTS74G0VBktvnlcmNuWma7jWh1ELoCwmxczT4Nlmkcjtk
a+RJLNR/J1oDte8JgmqvAPoc3kkKR35ZncRnEH++byOGeFk/g6IKcl/vJm0WE2mD
4l2/5mIw0klPjyZ5sMLQuTrDUG8AtUmJtcvGNt1UMeBMBLL+wMf68RThD6PaUgZi
jfSJgiU+6b7aKnqWQTMnWOLzmqPlarMKFzUrFnnaysGGSA4NuNn4Ro1FslFbdP1F
y2jF+oKPB7ovY8JPwse8nkcxRvSwMPQ+o2dNvgwBMKcCATaDnpfc0qXZqE8cZHMz
RCBK6m6NtOiZwHm+EfGjnCTTSJHHq6HodxnLgB/M4b4tpHGey4aAU8OcgEaEQ6Rx
QiTIN/AZ8xkxeWuB/PLsl79eoOdRs7EmMU+ki1nlhwFZtIuCQ6nVggEbiJTvaHSA
luSinpDRAnQsPghu5NDrO5mxCCJWXyfZQ35CkwDdIUzoIXvCEZXuICYxun9xDwid
o0v4AorvTIEx4eeBDUjcGMRA76rFMPyzb4fc+JUDntnv5binRsSsLcBEhL2kPe+0
72bU8Bb/NFoG4dOLzRDT9Gge+Fpcq8UryCYllo9V0MuHRcgokzJbjxFYq4p29csp
FFfcrz+ws/QjQW7p5dI7oX8gBoKf0ghAIO17qZpKJclKZmkfwm9ZeqhZbUCjeAL2
dz0mET44ZeFhSnTzXCDckJG5yzypGk8HRL8GX4KA+7aCPKPexGn7HwPlqpnJpzG2
3ccLc2X1XQQlelqg1NcgUtYcwGanyAs0P5BJb/63e9sN3b4WPdS0SUmQEYW638HP
bhZs9asKrWfhT4FFhTvcyeAyHA2AnyHl+UjcKLkpTp4tHAElaRAE36RnUEj1PsTm
xwF22gylUJLZcD7ejR+zvxFrvNiuqZRxfnVeKagL1VtMs4pB6lqXGmZyOToo9V98
ShX6OQ3Bcf/UaVTsB6hnpiCpfiFUQtR3mDcli2F3/uSHq+Itk5RB6VoaRdklifOo
OmkPsKdZQWc6Lvyx44aB5RBRc39MKcEmN+OmRAx8CslMkLaACnVsDCn+2nGXRB6N
gSfcA+srm9RhXJXURS+ouvP3wuxB0KHnbBpJfHn7+JI+DFdBz1A7uimOAh4hu2aR
Sn1XpAlhjZ0rvriw1jEJEQ/WUwkgp5Kr0mxXDla1SY0r0fl3OaBVOr5xCd5DrPYW
/kMkUSX21O9h40collw2zgAOeF/gllUbSnPfiq4xIt6rgnjpXPCnqcVBqmdFq4c0
xWdSz8ZQ1FB/YIcbw1OH+KFUzd7OWG0+T6vkO5rGOMcABQs/1s9nI1XqJTLauwdW
uE8EAXG9ZOzR7aQMNfYvjx+iS6ttHM22M+MjJQgaovdDyPNU3gwdx2HtExhOezsR
2XTEhvCCvcbKN9lKtBJJ2o2J62F746IPYKaeROgFcdbX/9c8Sk1EeJNyKW7UyqEX
PmHe/u6sF7QheHD3R8uasCplKkJ9RmCJXbm2K2XM505MF8ScigymzwP7tXCb/Ngy
ohbPqju7YyW/tx/IH5UIUu5NEp8s2hRBq9TwURkkT+ldd4jjpp4hS8WOhv4FrBPl
uGy1PpjNiw/9ZLZZwi8smaSJp5O5kdcwFtCGlo+qLnIFapjA6mLrTjgGGJUxm1j5
wGixe7jJhskFCVszi/oXpxnlmCEmAXlUJ1QJ8QG4qzjUiVqUoQm7/E6Mfx5h0VrC
y4xvX/aJWYu8Z83JrnKyS8AOJWaxSLQA3oRSVlitD1FxBMpuR2ItdxRCm+wGy57H
KAqlrAMG7JBwsjXod7gzvQAUvB4EBJ3S71grqy0UIJMHVzSuGMJai86wpU9yxjee
1PbL87lLaxtCVOncae1VDY+kDV+iNuGJWWt2ED989nrOshbV41sKeC9Vr6abUnbk
Ty1wWeGqiZxQuSqyhoNLl/xPTtebg99jFlL18H2S/YG8uNiWuzPHbTTs+ZETBN7I
WbqN/sP9MBEGQZeNR21rBe8YEAc4Z1BVlhHZKY2q6DADC2t5usaJ+MCzRPyE11Qs
WbzbgcyYLuY3yI/85AX98l4yDU8lvPy3LRQZwEFCM0VTLSzZWIO4Fc1kgGFknHp3
de9Oh48bNBXCy9Z7WmBtmAEtH0XK7mwuKEU8v3ZlxqkSf9rA4w5fO9+lMiTnH3YY
N80+EeC9b6nW+qgNTtJQ9Ktb8eS4A/hR1Y2TlcOARaflEC2rQv2GJ5QTodYbjARF
Apl0OJU87Texf4GL3663sKQOBR55vXmMgWCPVYtYV9Xn9aWRlqqLhorF3i5YdKTm
/DCpylYDUswx8mdBsmPVGSiL3HjviB9Ag5frkUJ1RHnVchWm9SW1hM438f9FTHPC
DRazzClelJ8E5pNWiFW6mYKePUn3aCq9WBBdiXFvZVaace42n7EY7BE5XDeYcCv1
ERgksGXBwd4zLTi8spShB3TGxERoSueQbxV9SrTVXaqwlAXy0t4o+KKmtBgWF22j
MhOudnPLGlMG3Vz59ibFh4GfgCJqO7Kwy4bEtKst6SWYLUO7lavmwwO6ici/0qaI
mjR3BCUdgJ+LTuhNJsgVD2+5uI07eFasM0uJPVyt4DG02OprAE+VEFp1Tu2a2/1x
eu5H8V23RYkl2QtNS1x/LqEAHA7UYoX91GJabRPMS4o9ZzDbuR3pDyReTv1yBO6C
z5tKzbRaYBKshQ68UTzUZvhq+0Uzs1AUV4ttGTerZ0ZV6ln3KnlCpCr/hBnmFxOe
T0YW49wAOe8Qzg0BH2wmwMCCuMQk35OCdB7Z9hVbh6+6FUqZ03QkUJEqZCUcMjgk
IWINpI0mXK7/byML4fmzQ3xeLPRAyHjGY+P7PJK9q/NgSw345BL/91rIXmeRDb0b
6dt39001EhPdVLAAddY/h7/mhJRXhCP2rh74Ti6x5gHphjfVXdMiGoXCCM5o8kWs
cVYzjzuU40jBt2VLsAMNJ5arc4zEv6hedgLo+n4a1W2EYpok0O6Crkh8WzJxaLj5
wmKqx5Erp7E18VDCAD1KLuC+7NQ8UFc1ffkL8a2WLftFw0iuZDvHrMDE+OhCOLAI
3lU2kKa++lUFhUJi+yO8WBwsLlEDAJDf7+cyVG3DHH61voyP6mGK7/1l5bJ5saTW
6coPTx03E9Qc1XipZA1JJRR6TW17jKMqlh2D9L9KX3OaBhHUxY7i93kjYQYTGWs3
DoKzQRVzD6cGaRghIpApcA8nQF7rKgp80EtED6CTmLZSUqM5567ce8kQBSzyzb75
J6eOS9GToV3t1F/IJ5vWuzdRRqfZCQI8q+5CzTJnsZxT2uHxT18cL/4LMibXOKx9
5bi0pEek/BFqpax3PMa00iTmx9e1AG9zuZhvbsILwdU7WLelqqh2m1h/uexSEhG0
tkQ4lTko9xMavgcRUvN/4NjaPTALGTAaPVNuvEclaoErJueRUc203iAQl/kb2t9V
LJq2+38syne5FimFRGd/bnT9PMvJ6+HuZ6Q2iAHUzvSK+23cWeOG7/jW2TjeSFN+
C3CJNJnKzARC47RHzbefTDX8YXnCwY1L/ns4A0y+7/gjg0gFH6tvWZuiAO50lnSE
mTk5QsoIKD0jFfX6Wtwj+42gTHcrDzwva1I5J1gTATTOqbmp6wsssPGTiXpgWI6m
kPUpieEeuFS26HlxP5HClkIKhWE8GKZkJL9CSVLtnmktBgKxqljFZPsi022ZLBR5
R388J0e83Q3O9E/oi1bMT0mMdrFijMCyqo2vJ/DnS2uH/H7ze/MbBVL1O2qmDEVy
Tjf73CorYT7W7bP4KFVxAm2VplYLSHnzMPeWCy1Ta13BQ+OiRhXr10ulMdWLL9MM
u+O/t4jbY68OiyQnDT9JoPmWHoHSyxwPyiY38obajpFmogUUSeWVO6ovQ8RoClfj
7LBxHVMQC8wm4tda8F3vTPTuwj8f9dY6bcXiiRqX784fUQ/TDZri7YZLpf5n0+qq
LUjyPTtPBujvK8fdi8YWVlgtsJao8BUlfBCuha4bs1+b7OIf0BvMuqMhGPt+qmNj
I7S24VPQcK3Be2ifcP2llFQ4w0YC6/SQvplJN223YaSV8TOyiSgLrpgbs97qfyH4
+FFZWroJslUzuh3oD/fNrOI4tGD3KcK81BMAC+b0ELypDTM7Z23YDe3xobJTIddP
ccnOSABJCgX0WWXS6G0pRSH/7aD1VQ8kxdS1b6GTbdHNf/AsB7743e6/uRlURTuB
SByKu3296U5bwRlg/sQzMfH2bBoVHn26afrG1oQA20jOu3aFa4IY7UwmiUV+Z+Kj
GZcBbrINUgh2UV3Ls3UeAaNuIKvInbwj9Nr+bY7e60sQkSGOl5O+ORpw+uX84VFa
oLFOq0CRubTDHr2pTHx9Xz+hvGlOW7j/qO4bFgIqugfmdwAq6w939oqOUK1hEUFd
4ZTNhqWn0/F7CxSq0SvzwUfP+/CZtd4b0uExuuGSVLb8DcIBlflK6Oc+Jkx0LnAe
sWTZG+VCRdvgbX+RYxQ7DAT/2EhQh8ZX5zUXJC8AZd8A7+vLp6e3gFUNq2tKamh6
cT13TiMyZM0ymZB4xQlOx3JmxIJ19MHhIao39vifcp4crZiOBZgpbRTywRWTKGwH
gAtzG97pBzakATSmG7XY5PtPBBOSCjPvrrftfePpFaR5peAubbRNGmyHlsKbaPwj
UGkLqrlBlME0nIEgV58VX2kQGASHphZFe1pCNagossivE1CGRXWyFs+4WTqR4fdi
oVzRvS+F2hzdS5XisN5/3GV3BmIeAoiG4qgmhnGpM6AWE6z2S40q436sh8dUkiJn
r8WpNUa3X6vGepV9yxjQ4DJbi/rR5+7p3e5Xxu0m8zpqaHPsJu2XyJ03P0MtmeLL
YAVsogMwXFsCvZv3tsKJveMxTk8AvfSrOHksQV5/kCHurldq2nVadWaODFxc2WLn
WAgR7nLMRnBlU2zuOsrDqkqkgBLRy2UiAgSwOCwwlzdD8du7ZiUmaeBc+f6BY6Tn
cwRaGfzM7LtB6W3PusE/ZeaWwf++3ana50sNpEjyzQJcsObq2XmokCxtEHA1yK9v
edG5lAMbuK8V24R8YNqidNqftfmqTgWoxhMx7pzo2Mre8cTSIiUJvMRn8U/BizEx
PNv9rECc6uYFJPiLBuJAm+oY3/+SPpdQDscB7PSVm62GbVgfjpe2WKk2npw/xUpZ
/sBZ8B0qFma+DgvBKOCwyilVPeHC55juH/lFvUxG2M1GuDAWr9RJnDTx+EcGtkTM
xEtzThixv6VUgivHB8DLJ8EnAmOQP+2cSOVf8UWC38XjItwH8gdiCZLNLIHA/kGk
wCMhoGFbbWefJhnqOyPNGERAQUQAnlKTPFXhkNgg6hThW2P3KH9rKBEbCWhqeEMY
7NEINFQiUC6sa97XkIrk59i7+CKRL09DbuEfVq0tHGcXhbAQoXkdRQgZrblZUYts
fbBbaRQKbi8s8TDiYFmzqVPy4Au6Ya/OE8WFDuYDNqAUe0Gc6XjBDPpXHbDiBdyO
BRoyLQe/ZsUdAOXrlFNZoCL6t8WlWLBqHiYLlr7XM8Tb4j+5U8SMcLcUZkYX2MjG
wLTy7Q0OWg/o8FzZtn/5Df/+hVs6F62G9fa1v+12ISBJApxzgnV7Uk2tYzRnPUtL
pQPp9za+NHmZUBnfPZHsfAKMknLoGcUzspyjOPfbGH4PJMP3IaBBKEQ/8czfxuSL
1pf+hf1XGUdYI0JII5LQ2dYvFhFgk1xGDNJOmStRlL9XVfnZLW1wRyRBgmHHMgNi
sKW5ufMBq0zsdYr3gJEE2AdGk41D1cI37KBTHnDP8nDz42oScI0mqvc+1SREgrOb
eEFBwPzgYyU9cB9ObLolrdRLbSdskKeTgUCyxTS2UuxXFMEBu3EtLDT8KOi/26QC
oY/AnMf5/lLoBRUQKO0xXEigdwcvvW25/DYYYrfl/093e0toiG/6JaNVY6ZZtg6v
pTIGymRhzVDIv5QeZZmqCjn//uBY5Q4etj8v6lmkIH3xGmLnWNI3u30Uxno4fCub
yEoCjj1XXn8DFFVzb8bTb40hPjc1ACz4Zo3sY1KomNTBgEiFhpQDIVvBu3/pAHQV
VOPRT7+t8q5GVIUMnCVTTy/rqZ+cDmkztp9CgjxOVsOv2HLYDgPEgVznBwjFsAcn
cUzTaqpg185AaQKCmHcv4YjYtczcv55dXzByCIYGfdMwTxMeM+mIsw9HXfkC8oba
Gu02jriN3eIdWY08A9f/B/u9OQvQj3bINHFHBoZkySHzEqQ44xmsMP55OZU8uMKj
qPrjdjyU3WYac2NFXHvjB6i7LEHbYgcVrgXLdGzOXgPemEcjIdZPGPzAqTW2Rc+X
i0YvDD2uXimt67Vz7HM1/wVSr0FLhjWgNS58xChvGX2Osh0PLaKeuls0Um1lkn0f
OJqIYtLMWWZHeuYrKyCqQgtvR99wov2K6NPAHeQTUaSxbz5+X/ZccS0IOdEGX5Tf
imkVZb+W/yN9seFANr2kcmqbVkIgiFOxOq/4Ql81yVzAtKsJUoqJka4RwVWuDMWq
yPtODBu3ZymW6Vzpw3jnAe3J1IqInTPy1cN37maYAT9AR7w3nzKFgTKgLwC+oULd
EcaxRd371J5S9pYFG928LDqI3+YFfFrHZoYQfTD8S+GP8+o10jvJFYjjZCDeoB2+
g5RcMmmT+I5PY/e2Su7gq7nf5/+NW5iuVMqDHILM+gqqLKNFHB4c0f9dlocCVaHu
Z0+cPFfdfVj3sejT7dqSlo+gYkeizoLbnKjqHpQcWDan3hZo7xAojm0y9HjBPjCN
dq4E2BDZngDviQucX5WHewcXuIIXY23kl2QiHPkz93vWi88OEB7U4S273PJfU29O
SMuxlEJfpyE8xDvhDjt1HBAsgnMTcWV/CGiSMDcuXGqF8cHxDahTvxOZluKCXDtr
mF6pLPk6e6bWfskRUtsh84OXiBLYJ2Y9pj80wPmxMRfX73Lr/GpMjDJ4S6WCE+Il
2klAvlFd7Cci/HQPx/qWM884JRDYJdXxuI/+d720gRr3PwXpHGTQH2jttTsAHP89
+BwY6C7/fTwlJOCPtEeL68tQCDcOaUJ/+AY39R4+tBzV6ZpQWKruuL/mFkWSqaZK
pm2yPz11VYK2warjblUsY41GaPNONmeLGmP78u3OZpZLVLLugoCVnLdK3Js00puA
x1a8zrvYtlzUdAKhL3rAbH/KLzkrGUwvf8OTc/eJFReBTnJKilxo6ELFnf1Mt5/5
BxhPwbIaTHU+IwJU4PZ60DEOVCcJK8E0WW4Td2UYnQM/TtxaIoC4LCYP6t4QtYF/
754zTqxanSMUJRMig/tGHTJW0beCPlUHLeWZbicjpoam8uMkQ5bxndCVrWsXBCOU
PSjiEm1lmzUuh/nODr/sTu/JmZoepA07wGcXrqeXm0K9F2LHDTdjjKbud4N1EODG
dhZIx/XOYpvJ8hDeMrZUA+4TrP2YbJaAhnrjeEmxv+TMNQfoLTk5kqaIchXVIZrJ
52VSvQp6p9m6OdyvFx1RaS7b0+hkGN1eQaDbgm536IzEf8g/y9R33jtAuHGz+URk
QRIylaEMzWHoqxIX+ve8XKUbzBsaj3bdxwAb9WhXILr87wWZsGgN59IZ7Ot0J3rF
y0VtamGKyXY+1lPZO1leTb48KDPCjEkoNZQQajhojrxacCuzKS1s+8MK2KKPArJD
ADlY58ykUzIa7F9dC63HY6PohDPrQ4hCfw4IL1i309hivAz6vNt+kUNjfiQzDsi2
2StFyv0VaklYcu2XU3lxPiQf4uv/m0Bjx2nUH2HD2OeUHJA1j0u+og9bXyy5rSm8
2LbX9OCzICGCI9cqLwjYfqNnaXPgyqxKcclvkef2CQkfVzIma38KUmQZRGXbZ1lg
gwTL/eZlAMvo6xgFH96bgP3QP62ISHISCnbQ/fefhLgAMyIeihshvoqdKOudKxNW
kfpjWElIqvt9KETzSK9TwXqN5uCQmiWIj+0GP7znUW4EZs7fy1Zl/Q0oMxge9S0T
L6CbGY4/XFtDcqGM84k0XqyNmtI1jCwsyTKcAUeZZuDsAIrgGwqaHEf/9x6iDwyA
Nskq4Np8pgbt+ZdZrf/cmSeicfy2cicQIfpR7bZBkb/5jyEzK2l0yr2XDYOqdJbH
4wIZ6e9uZz92QqQ7hU47dvjYWTxbBWf/mKpOiyx702BpyyesDuE+fArohvDEpkCH
Ps6IL3bxkYSeJDjXHyfa/UV9PqbYHw4FuZ7O67Y76wu5a7sNIXcUDHLEjpOZPEl0
fpngZRP25jd6mz77Q5yUMRMePvfh2Yyr1KG2eUtwGZlSCNb4/KnmpCdVo1dNC2AD
EIVyQuqiekcSPA7InuiOL4sBDqYQ6rU3/2a56qriY8HqPlCw9FQnEd+AfhMTs7d/
PuH9vusUzOn6QrRsEQwZ73wHo4CvpJCh/4rwQFQqvtWuSH2Ub+uw4vbdLdbF2Rbb
0nqDkPabLZuC0GjJ4mEYTjHkcp+FRWt486w9lz+koQBvS7nipozBGau+8679NM0U
ZvyuUs33RrnFs8+IHIqKeh1bhavDFMZd0Se1DgIDwPVTBC4Ccb+Yr8XNi1B3LGRk
lMp3cstyKqTFLOO5+1xaSJG3rdXSXBLfawUyglKpMixaTBKrzZO5GOP9s9w8yY4s
yuvKJ7Qau1xm1vWVnbo4oD2guXA4t+WVUzWSGB1aSszJh3Ka76oMUUoOK3Io40xx
zzGciMytuIvz47B25e+nrgPUraB+sLxNWPflq444X2gNRlBSXffmQTRs9mFqWbJH
BfPPmkpeRjGr3LgaQabj0G9jbniGxUawQWgID4aBfsTGtx0wqeXQ76005NiaVSuv
3wHprpYd7oNXcB9ee42lLpvpILTM/oRCfYL6jUybgr88yu1qBtRbYAh4ISEu+6SG
KNmhDqc6h0fxW4J7sNcfAh6MrVKm6DjJ/6nWrWDL9qnRV0jKh8ydDbzUznfVIEGG
RenZKnvikVDMW1z2ufTqHQ7PhyaZxSqg0TebGe3oi0Qp6KlFtkGZNWFJZ+UHJqG0
QV455cjeWgvvFPlys3RFUZudoIYYaLFsFPhcxkS3OUzhuj0fUL2dQ7pQpqf06NY1
a+uIUeTCEIRIL0vpQ64HrHdVbhiNX04LvjKeP3TvGZVsx1Z5kZllgrbdgTq0lMZ+
Wtz1pG83AYLJ8nyMtDUcLqlET92e+gMACGAyAWV4GbPQlRm5rdQ/Gj3Xni4jqsV1
83m/AecZDfDWAZ//Kb1w9X5sIazIZqk26r6iOHoQVHZKrap6amcKzFV9IUjsHr+X
Ip2BMVPpJlYHxmVmwLAUmOuAiBc3IqW7ZuCxWFot5E/3O7b0YERsmaowysZ6vgrN
zCZOPe+nnOktoq48PV3Zxz06woXFvEsNdy4RuM9ruK/X0aXpiPXAq/T+MkNxwVAI
Smmpc9uOvALzUn4Cpf/4+5vURLqC970K79RyUdjCjA8Z+UFz4E7dQxXJC3/owzIW
InMmrmWXkht4QPHXeE9FjE+dZgWA18lX7EKqzYI5AHfLunOcA8jkayVUYzysF/mr
qJrdZQ6FECAVkZ6Sjixkcgla2IFCOKNHsygHISsMcuAA/W9g1wQWYFC1YmCe+XIz
VH8k1kGQUMDoRT+AR1oerwcoNff1yP6RGqbSj5OPxfuy2XS3easIhZbWTsUV9qyD
oHYz2opHiNTx43zlxBL7IuQ8R/G4qpiDmZmRr9wUYzKVvPMTszLRPoX/7lelWM26
EVI45TU714Y3z7JJfvZUJryQ6x2RQm6U7ZCwmxyz93AkUz5I66kAPez7T/nOeU/D
nRlbNAPUKKS88ZU3/86YhRFwwLUHMJC9n6QduFLbq72TsU6lDZsNLkE/xUE6RgNZ
xqXlD4BJwyL3nx4d3FPBmCPe9iil1iM7aGt8hP1oYfdJsopY960CjaV81yuopdHw
4fI1xXf29JZm1GNbcp4fghy3BrwcsyEEzhBZufovf0F5LftvtWWJJVQ/HanDAFcV
Vrg3Lyz7Wn4FplrgIwoOrFdTErNxbp16SKkiFpTJYgj2nYNpUUBPwJGfruwBG8xN
kUwj9fbD0ovpU1DrLuealsnoQ+UukmC/46GEthp9s/aynbqojUii1acKvcWPreo4
KJPyu0dd+IP9HEVcqZoVEulxfSufQv4l+AmuSTNpw05goxHHOh3JYB/IiU/1vy+t
RoXDvSkmPKbn5jwH/zyKYF4OmoJM5q96CJfW/WnHNu1jpi5tvTXtTBjgqyKwuNwN
8p2FdynZjv/mICskAgAnDNXEWVYuP+/Qbm9sFZKjqTPLS/IA8OQoBNlxLJEfWCLE
RX34f6b3semIQZqlnsVw7Cn9OD41ci+Zyit6BCvO9Ga5oXB62LYLw8T/4IuVHUV4
20ikFPlw6I55zG682Z8sWqoJV6w+l3zneTjKwkFBNOAfyMiCUElJ95L2cj31R0LS
PaJPE9Cp7JpFsIPx2vv5+BxZTh6rQYWx+gGhgIErZtKDblq+/nIlK5FvCox2OLIl
V700gnVxMm3mMNWzPcNlCQPosGsvP17EvVko5luP1bl9OBCcs//EYiA1S70kQx+y
RkjF6KYSz/uABQxwgMWkNqGsWIkMrEL58woduspi+bIIqY0XjL9RUY/WozSzphxt
X3drLHR4wfXjaAdnVT3ugT22q5kAcZEL9OTh39CHd3xa2kWW+kWbZvcn/gATOgpC
H8L1Hx6Rd9YzQL/IJFWX5sQ7vZ9xQnStljSkprPjl49u12A3FlB+mTqn1Ir68O0w
tbbr2KitPJYgtCM10M/eiYRswr0l+DbHUZsyMXsLFxXWzoGrzKNUh5RsldD92fZu
7L/Zo5PEQ/iVNBeh0CcVFXpNo15+SQr2jSF72d748M+AL8/5Kf8VFtVDlme/0HRJ
4dZQ7U0r3fvdcnWeECyTaFQzW+AAAl4MPzte5EmmU1BKfqQl03/jtKN4zD6s7off
ciHkna65VvtfRMIjatOGmzeWq5jpKsO1vvLkcSlggoRGojOGP15XI9x/AIspQYMD
tKgnZLCTeAzjVDdme8k6H+7n7oqi6iFZnxNibxzgO+tenyDoyv/fAbvNJBz1baHe
qvdzvq2R91PqyRCVNVjtzStsNUJcmSgtOLSXgD9bDi273dZoqyFYFhUj/c4xOyzc
Uq8fdEo/yuUe4FYKp1uzQ34VAHjceShv1y67D5/Yg/Townev62jwPgKlSbiq5TfT
qKZ2S8Me1inzJNmkMnGMhMSqoOMLELApSvM4fjrZT2gae3FgFgqSFtDIS6/gs6zE
t98361L+6ZXDrGs5+FKrfaR1Sn1dWVLNsjL+/0ZgVd29lajw1FrD/YJFi8yTii48
f4R+MoioB4PO3qcL5i6a0mwVWV0r4+MToKLqj4rhAqjUH0j0KSt2oHWfRH5YcodU
l5L+n94dDw7TKiyPoVn39bViM2F9fp6A1D+pKI8qqf6VySJAz+nRCsykW0dXKvC/
Qv57btahK7mQlQZImRhEGWGqRws2wVH2KEOwRXgh2EWv6rYEVK/McWGkhVVvwzVM
mnkrILH9ETBQHCGka5HR0B4xLjNfgibEjC4Dl/cpzbCTbQlVK8jeQZsjiedxoJKu
H/4WBYMNKw1tZ+G82EXhzia+YlT8GDKDHjN4QA5dHtyY/n56OIOoUl8yckkGxbId
oDNpDfkFA+ZtRnF7QXuOPwj3cpDVs/pfYNr38nmkshgRchw0ZrmLr4OsnMe30jaY
VdEh716zCvGNRNY1qEyo02bKjPN3F/YjyvqTlY/Q6unyIx/e8FKcvDbqOEv9zczh
ppOlotMI+4l+MjWvoNOvu/Ql4k2i1wm9d99mNoLMmbK2KttHdt3UgVGNvhOB6PAK
c1fmu4vckcouJ14Uzc59kJb6DHE1bk3NP3fOgqKrgtszD/eX9rtzBkI2HT/fPPSc
JtmX2zNw+xFja0jukULskFcadqf5SV90ElzuJYkMH7pblpkF6/WAySPF+CWRwHyE
2zM2YH2bseNL8jYzVqX3+XmIt0bjfqhc2yoxDTRUkxeAxXCIJ5muHTnWGTM1+gIA
RanbQYNYhbCktsV1MNLhXUEXfQJ7SSbneXs/9uBsfNkM4KzMxim10TaOAtaY6n/M
dKTh5NYUGQSo3KpDK2uoIH1VWZ2iHFN/TGbcXOy8NFmeJrUNtNCWZx1A1JVRmQnX
g9JiKD4U2xOz3WAqSGAvXWrEBWjPc/xSLRmHShmHqxRU5nBojcErevyHvz5ggg1l
NgTjazCYV4I3buntDg1M9ppKLh/e9T4cvm6S5bHjgRbrnDJdLSaWdHuQvzk+UsVY
bbALB7Gfk5lYkcNJ8+qaxmFJX987ectK28ybnTZ/AdYtkHAdwFqYR3uv4Kr3yJze
aOBncmvO3D140AZCsTIvN+t/uC9jz9A1nTIOQjWm+dqIYHZRA6WWT8AzQ9lsfTau
p+tDjO4Z8TjYISmtCw8LCbSPPI9iRPU74dtHU64lG9Y2whWkUSKURj9niWEKpwxQ
wi/3AZb64tX8Ly962giv+ikEwt+o4RSMEU8x7as2AaPi749URV5BtWBQccZI12UZ
9PoHXjhLA6eOYdxYMloRlCeBlocpFnY9KVbiLA2HlwwqObJocf30BmYdboB0izru
fX+9eq+nUu3+YLDNtLA8zCo4LEvgVUzARNMQvoTCi2SMY6WX6oZ0x53xuMzFxGf0
Ow+jAVSj1K2/6datuCsKIU4xd276kyFrwZYnvpArgvg6hUgXrp1rcXTVh6HleKi9
eKgUoi0FyJF0ArqKnqBPp/B/sblFYXEOmCLEBEYIez5aFQukYuKOd/ERypdeUdAe
GxyfKMwn00gzoPWfdExr/CQKoYHiVkiy0SRc8dQQK1mvAY6gjRIPWxJaJepFVATH
K7h45++S8T+tpT8yfkUgTpOY+fW+XoJmWA7AtsZx9StM6kIiuaIcpqBs3/Z/mxFz
rDiW8gIj0Wb4RJVFW6laCVPAomqDRYLo0440erhxzSC0cE0j6Y6vbRW5q7hdUVEN
IkjEVdmnBV2OlSbMlXZlIxybR9Vq29YC3d5Ta8cUS38nIsmg1OnGfWo5ShMcfZCT
zjibrYG/AreE0QoWkJEsddPmdfvUBMTxskx7/5AadcJj2dp8L6AdoL5YQvYBmRw/
bQf1wWDndMmuypGwh3TcvhdEJEWY5LmmLX2biiTwK2Zquz6Aapc6BM7X8gVjOnVN
MgXIh0NlVJIrjC5f1Oa8rpHnPVvvSEfw+ejU04N/XG3P0MAOBjnFyTHeamXrcxVE
Maqk/1eihDqbotMzjAx4OOVs0vxWkxl9AgVOtXcpLuc5yELGFmyLGZZU5h6zLb8v
d5+DCd+6YgGH9/DdKJEM5TGGYHPgcKi97Tt60ouIrsMEMRr33xB7V4vW5WH8tPN4
vGEN9Rlbo4xrlPpfQ3u4hsk+uu0pWHq0L7s1mdx1yhVdr8JbM9nAl9x3eMDBBjNm
bzIIy3Q8JRpfuW/S9kBEAbZt65Rnz4HauDcnT47zR347s4znrpZGfkoXcsFshfLg
vCjaQxwlDFWLYsnDfAJ9dcCs3QNEtftE8lSjoYDFJaGh6cLh9PudBYkFExgSZ0Ak
girjCKLXCxx3MAJarcfUMl4rqtUa3ydu48vaJCXe8GxQ7RQeaGL7/L8t4S1v5uCu
ZJR5/EuMczn7D+fji/1SJni3Vf+P77VJwopINFGfBWqtRaF0/Ih3sJFEWZWFuAxw
F2Jobibz3iZHcR6n9xTnB2ZP7i8C04lK7LZgYyugYnQcHkDff40t2JrSqykcfuNp
UafwDFJNwogJIzJkczf6jecbLCDGewzGvmG1FamFrPSG+Dd5bwf9Xjir8NFUy57K
1V5grp44Mbbs7gOmMQL8zGKy17MMcYHzrImtIvcU/O4FULROGeRXA9xyS9dPOlk2
woMcgfBk1XT3JZ2WX+cBkBO7mINmYXIfpdDhqJng0X4YIjJNNKAhElsfJH4TxS/Z
QNUAs8gs4nMtMwUOi2V9cnmWpDlwMjg4F8VRdQpOuN41O11XhnpIxprGWDpUVhQA
8DnPYufLi8VGoUMhyql4tdrEzyvympp+Ph7KMZaxn8A6QBYuGij/H6+/xv5CLc51
jvmRghScE02xDgBl4WNGRr0obFrlp5vNIqSCybrTSibjXaYOjJAKUs0bwkBqBuwF
lyDlmeqVrTj3kTAvcU7QSfG++iixtlvODkWmqYim5CdpRrKxHYocxAMWFW5zNbmH
ScYd/vff0yruYm88QThWugIn52rw/m9xEIOF98Nf6funZvjbxWJb7o1+UUAu+3O9
yjEvQwy4wGOgwFYY5DWo/q4ETU38YM7pVqgUJ/37fGMnYArFxgEWTbedtD9fuMyU
dc6/SvRrIo2U/d7pedit64oA1+RaURD8VHEfuSNRmL8FrwQThCGhbYoX80Joyg8V
QaSL6W9t35fgrevuQ2N31s+7mGrOwJKUPyiwnX5i7YFBPoEHcGVyYrnAHK/wSk0W
4BpKgaHcOgHXunn5x54B3IYUcGjWyBzb9L75lBP7+JFuac8EDhnv4lMthLXmnAB9
xoEGgc1Kp2zogzNDZTotYIQ+YiJTgm+C5+dim13PmO837UOIBgpTuBhd6VfsnSMD
mwddlDWRqrwtjd5QRhGPhrQTmadS4IOHCCzPtC2QTgBCz5ZEe034kuCedmPur8U+
n8PXd6N/gkDPWvstmd9Ms36CYP7tirXjnJYcEWP1hrakRFnDTSc5RocoyCwDei/T
Bb4Uhe07aN5EUb5ZALkvfcJs2r6Cb6TlNsFx1j4IGwKpz85p7h+2H8HOa6m9qD9g
UTIlxgC1L/IBeUSA5zuigV1eZqY6CwAyPlUdaGPbIYUKu2+U7OWMWXjlsSgK5uhw
FPRUCXgICekbXUmHpgZRYaSMRTngtB6ptM710LfI96xD7ZE/ZiH5MY6+0LfLseGQ
4dX1xJPYeQgk36d4TUK0XTlzqoftFRDR28cU4Yw1GwhHOqYy0JMc01PjJDpYSUNI
qCF08/QazSYdPQrCUNoBoo+GN/N1Z01jbqDAVgidSpu9Rv2ZnJgvpGseLjTwhfhx
RyV+XDHMB5unxMxWiawPzSYcg0yxSHwOnRq2MkfqfD51I8G8uPewsi3jgz0WnOgF
F9kdjjKnkiUkuwm46IZr8YffuczXGeJi5RngaaFO0earpu28AM20lnB7yCWESwnF
aSuxugU/MkncQwDp9mjN8FXeQBXo2E8d+yFuk5TRI+zav+7HJiPnPbyTFYxjflK3
t3UQg/i5rVXGI9sSoqrlpPBPJf3RlY94wDA8khuarinP7hEd4Nou2HahCf8pFSha
YFXqVWBigEStYyzm4D5cxXhrWbHPGMXuCyFN5r+pLAS1ZO3X9CjO8ZUymFDnqnhi
F3JIGNx7Q7jI1vjSALryi7X1KnrbqG+J3FFjPIRjwvjO2489GVNpkXmR80oRUr7d
OeG3XamAuwhhUHEQGfpYP+XAe6uDrJAgi0kp832dwOtTbb05grjg6UQQsfLhFj1+
6Ve+cWVSDETHZguuSP1ia4eUBeRM74Lm9plySeusyYy9LYfDfSCCOXEDk+O8QEgn
yxlKLpBNrc274YgDzWpTwhuDD/VzQNs69ev0uAoIabP7uzEa0Y0nb22Zy5zLji32
1BnSf7KzWOoFzohFc3E3gkcocrkHFKvsmXjacjrTA8rfTeONHXHnZkpiuYJE+syL
D8sIo5Hpbl0r9S7eju0bCxyCbHd/i2Sm/AWOhQ4QKoyskpYSFN/8BrqS+TmO/6D+
mtHJ5dibLJV3K2uIUez9lCA0pqSrsKydngOkedZjOGgxTGytQS40V91x/36qA4sl
R0yVwzbN6p6oeJv1TLjppZ9r+xYYEVIRC8ZMIBfG+T36uUK1VQm+QHZgcrPU+Rr1
CG5o8AUllsOb67JH+XVCUNpADZRLQVO7Ly98hTthBtXaXQJpLel8l7Wv0XRUKNi9
eyXTtIDS15BSo8k6514050saVyiOeTsSIwL94VlNWO40tPuFFKp78SmbIVelLnc/
6MAps4Wd+9Zjlc9P3/MiW0geUxZqOiFCd1lN2+h1EW/mMFuRtBhoG9s4+cjZaY9U
GfaUuTDPRUefi3bJ1TcfMI87nfhmBuP76HhxnEjH8+Irbq9G44UX6kd8GRqThrTF
PvE8/nNZEnAIEDEhd50eHS0xTwIEYXe7Ysbw5ZNBwuJe9f2fcDbRwAoPr6lJH607
N3zF8OqNzETnjWZ3cOy32CXGmHGfGmbAx+hjgD4y8n4+l20kQUicCSymcFS3Dzy6
16kYNKXqKw4UNRqN567r523zswZ0scX129deg3+tI2/GH3HfziTP3XojzgCvBApF
hzng2FbNdwJYSIYxfymEWEsisd3Q+buSQpBqO88pvviD8v+yscurfc1r4g8HcDrl
pIJ0xvWIY28En3FIgfYJS9c7waJjOPeSdoE/is91me3fwNThDz0XaHHAANpcLIHu
UwCWjs9loNLvpEXA0R8OIWWWhaeD0yIeChH0UhtqHYkD5OLsJOoIDmnP+C58RWOy
17kBjqTOm1xn2/l1Y/VyK7DJhGylYFdu4eq8+eEYLsAhIpJfHC2FWHLt87Zm6Ovr
cMJUOOyJaKspb1ZpHubCMtA7vQw5zvMdj3UC6hULICy2z+fHH7JBqJQSdNbA7eCv
27BJSj/lFvItan99zAXkMIKnDfgkDUHZGBdT/VaFvXk9kMLPSwYq4JEKytXRWKFi
AKss2vqqfEm6b7/RWxRexi4O9npLWMj1t/vPr+SV6XziDVCDhkjLK04kUKW0yPR8
Tu2N//rSk0zUtuoZO7eTodZKidHoNoXJQmrpIxiNajL4zzStperuJXVRypcpGof7
HZymhAdVWuEW1IriTYv4zeJvK8CuxqaYCt6V2nAwLv3BJJQ9Bvw7/mvdJukjyPxh
Hj/cVtO7/WMtW01CxJcYUXGx8d6Ey2rEnxHVmmJD6oOmUROI5Dt/zjw0lwT3x8YE
PNm9pLGutvsmbdGlFjRMnMw5WJuNoqAsfrJEmSgQI0Y7ckkHhBwXpotRe+eSnUGW
8G/yFXFjDsTB9kWX79PLY/DXD2uhzSXMYbRjKRbJpMfRfvwmfYu8X79vLRWQWV5h
1S6mpvccYYmsxy/kdwnuFaazJV7lJLQkZlSOjycylknTPZPCDMUF0+ZcEvRXFPxx
D5qkyH5gXfABEFuIbWFkw+x6zBavLeo+mB79cXZ4H3D6YbBJyycyvGLCJYTHFOJR
Hm/tv/fOnlILFOkGnHk+ag7Ab3Ux1vO3mFPGJrGPWZzpOYopUAcrqd3aAP5TSjfT
KjdJmgRSCk0OE9hmeYttt1WODx7G6w0QjG4F9ldwQGGE8DPLJvfVhuIMEotCq+FB
tTJOqjnnAwzkg2sgours54KSMIHhNnKz0rdUCtj3WrME1HjneQMHH1qZooM1tDmP
0zbJcS/R6iertyYeb6n5XKAdCTve7k+Q5IY++H/+Uw68u6O4JoqHYXEt50u3zcsf
8Slwq8RE5p1sTzBw8zz+rWkAtGc6UzChE3HKZ2Lvm9FEbxm5OoOgzxNCo7yxOkXU
zlnzRUyNRvOJc69/wy8ehgwbdRhWGC8EeStoLsDBb4LIAHQsxjojucpg8IMpM0Fw
ZEhDsrUuKXFgs2VDiVp9RaTykEEjW26OaueBcm9F0Hc6l8K7+FlIZqAjcev66XEM
xgV6IQuwmu0+Ah4u7i7emS2dXAHKjKmMaiEyXyvxVWJMO3dlQUmZPYnfJKWX9fYG
2uuUwN7Zp5Drg7qzxDDTZT+6oTngBuTU1cvUiK+LhHNoEmE4RN5X2Bu8SfpHQh9t
rOWVG3dF1hGDMB/4dhTkWhcBkCtWku7k5OiwH7JDKK76aTkDtlpBwrwRKV6T1Sbx
RqMpOKeq0f9RjEa2b+fEE8uzudcOctt65X53HNZjpZg+7+uLO5NeRtFSYQ8sCSsi
Cyeqon51VvP0cpE1E57MM5zCyBWMgU7D241cRJJuJ50/5kV121i5D4SnfKp+Po/f
HSK2O1hO4SSvm73B8y4e22y42uXAuBjBElAh8Kxg57HsJ3t2OpSmIJ1B6CMhTPdp
hq5RBVxNfyGVWG1yIibrV+fYQxLwST/DanQaKvUkc8Hbm5kyf671ze6WdzlDKbGT
VuPKrjngGAELZEq/333UlfSMUfVNMo2u7fIWwH4S6rTzC+av1gayhrKx4IxowHaZ
CsHTseap6MsiRKtGSfLLs1iBZkVuiRUj3ikKK1+5P07q2nOval+9J9jXWM73F8Ih
inT3nD0yqOdBwWCJ+0IhI9friYJD4IZm3C+8ye5Ow4Dy+Qllc63eWjDvUmvYPBZA
6UDX2ZC3EqY/0gPj0YoHqtZfZl/w7wbB0QopUK7C0+4U8Dk4m1GtxlAU9911/7U/
SYqZw6PM+jWrdtfXI7Srf+hnuNOFNvmhZt8gBcZroaVXDx7xhuzeDTAc4pu7gJAd
3XS8FEobZ1gixQshPyGCIYMwOImSATkJdBLixlEb5D+xXkPbH5iFCiXxbYFRo45r
FLe27XoWrSYKNw1f+Pl13ml+nPun4VHUaEbPePY5gAFI3FiMOzB7hdDIeEZOco/9
u+V0EgIFQc/A2qBgo87HjjcWkDiOKVUbl2a3WlU3ceKnfpj/n15Hc3wO74t8Aijq
q+LQUMJEv+lbRuN3fajyTCoiPUlxI0EMuh7L8noBWuKFdEAs93nhcQ9odkHts52S
XdWP2HeC7Ln2GqcnerO35UHn8+ek+YZzvRt6xCwbAOt2cj/DJa4mBMnuvatiunrm
Eih5UPo3p+RN7binSZlYP7qnQkdFhSReEw5HGjgISTPZTyXkXBXO7yJohSXU6YN+
XQCabapDA5ArTyHk5S/dg4/DTDDE6U/AdVRfltg/jLDYs+OLXe777mOyTxPHydkv
RCGylCrCblQIBEMICUQStBDC2EUJ4Au3RkEfWcyCUYHiakFl2KGQfVg19oh3fdBn
XXHS62Vt8B5O0FmM2tKnZKQe1vLSiljTNfQUvZ2QxHbwa8U4G0q7fbPMaosBseMI
VJH+NZRJRaOc6qDZSWMZfuYzjV5ahM1i6iDQqK+4r4BR9yyN9h8BGTv3h94ITR1s
VDtZBsJla6HSR17dPoTK98D+Ba/eCQTdzjeM7T7K78nV1JjJ/cmgzmSZcep51lyt
YAfJwWFqdhsjktvU5GfZLuo4rPxfZLeWPUaCEGlzmVbyJ6+dPHqWW1jNeKZ1NoDn
M36gwLRQBcAVF75yQefjZLcLZ3tCT9wisEWcgZpyqrwwzlabmA4ARdnxdvpaHWSn
boblvGwr0tk2/lvda8/cvQpN7WkQfKx1CMEBMWQ3+OSazdNqDl3YXVssi7+LIXt3
i86M5zqiQHzvWdDy/W5PgWplJ7oSAdRG9nLiNrQTpce82rj92NUZ7rGDlSNVqKOy
4pof+Cm20FNOrDxaEA1VXxaodb55n3Wf+lpXZMslV8WaUOQ5nB+K5Y8+jr0kqYay
Wl350f7ZmiYTik5MNVd7cBlN6nRvPUPgn0Y4EU5Os1/9uYaJ+6Pvy1mfcR0ofeoc
ROgr5hHzFfP7nOglnJAICR2ipaQRxbVOXsqnJRNPKKPI7P5uCSxLPgtOpYdokEkn
z58Egm1GLWhC3/Wf/g1WU/HERqJE69snF1YKgwz+6Lzuz7cQn9cZY7CKAHcmrrbF
sa9h+vEE+4ZNObhN5y0iChfeF8auRZ8Cais3aoxiR5wWpcT+F6uZmvgn59TGpraI
jv2sD/UEGwtITtjvZVkncxkJXYendNDu2nPwdwLwlRq8gvKjdVu4BOZTe2gjOT4E
0JHceMHRhR+AIbJL9ebjIICAvmWChpQIO6OeWGlbHiD6ZsLdVJBVFeg6CkBqoYFl
ZReOtzQOHNaC5FKvvY3nYASt6jPu260AQu1obrn0IuiySSreULHGETKucF5l85r6
CU/vuLy0diBXf43w/6Yjqanv6uXIF4AMTgwk68lbbRzb2StRmYmusOYY7jFWPgOM
GDLA5Hr1NwuReALhSAzSYDU+St3CxEhgg2Y9oVHY81JE7uTRX3Nsb+ITjxHA11v4
TO+86D1Mn3wNkiLmatlBqjUPaE9+djZuO3clO9yvyfVcjWm9oQMu5w0cCOzXgUXF
HKZAlDzt7HufI/X9GiulA3SaCq239sT3TD1b1ZVRJP5sdfFXO9qS0DLtIe9Zdi/3
QsYvUc45j0t+b1JMA6/ULvgzBRWEmfzA2W3sgQvWHEDnTLdF022f0n82kaosAOY0
orkbI/2mh4kKvuKGX7rsEeAywJaYRdqtkz8FuvLEaNJ3yRCqQq2jVwrC4zJZV/ZG
dsAA6syRzYxZ2t9JM3ZQGm0zsMrAYXqQa89iPSFVCsW19fUuWAfNB+ckL03DyONx
p/iuCB2OJHEtcOuEe5VDPTzty7mqGT71H9FGWvwDuJgFhlV0wpi0OPShokC0CwbH
ZvWGKx+QFzhimPJedTa/M95Hw1wENlCpOyL+PWV13uK0OvTgF1RnMraSOwVNtFW5
5edz4Cn1qf/6xLmOoVXEToAZScA6H4fsPuKiLjLB/4BKcDwtcFBbPOh+tQ06Lo7M
tI3UgnD5nrVn2vkCOoRDlzd4jC+M7rZgDoMb+AIYdie1VO979zLGJb0ugjoZvfig
cYgdVpt/faXo6sfFm3FBUJPnDYbvmsPEVL1mS7zUhvgrvbFsnQGuOGGqLuP7SaIO
WuSuqViwI5lCrWrcg9FY+ZvOQ5cwYiTpmoLqVWXYA5lpZkj5KtkmP7xlP8gppQOP
UfB1qR8ZPoGCq8WVWzm4NwBsrqH4LFAnqXziYgXiEF5C/Lcnztz0F6vLIadj0KM+
T4/l+/aKdEMVjiKVxV8pVZaWNFlVh76wgMF2qF6ejI6QgIULhGkHh+sPrTegtZHu
h/1JJwVHuCXEI6W8lRxWr73foVf2SNJYRrRsMBGASFznVF9p6oa/Z8kRCYNSGRNq
AnkHlmtEld1q87lFo/bA0xByFBbd57cSvbMzLdsfRr1KgaePymkub3Rj0MLgz9sc
xa8iadhQmV9FoVpL+YLux+yq6ofxDyIOLag8uAvND6Ad94wVx0MwDjg4rvz86MXN
O3nbQbhdDu9Vl8N0UBag3xjN8KANy3z5jTd9KNgBtz554vSFSooHrGxF3OlpO32x
ZuiXBgSTIlQbqnorS1xGMokO743Q6bBQ+eunDjAArNAg9cF1PE6w9rlbIcrPYIJQ
6E3QUUiiuHepoB4m4uK7/hEDfL/6xuc5/ooZtG45pb4S+m72HLzWpbmRzGc8SZeC
/OSM/bsl6eq2oHbHpNyEQhRU30XRBS090tyBmwhJyGxFD6CRQHYdyEhiHFjgIdPt
uT7Q1c/qbLyD9dyJ9l7W11y1xB0cFcbgPsG/uAoEwfGngvRwp2J02wFeAtO50EpX
MRbxwgL7+g+9+X2esndj9DhuwfVGX8a3tM77IezDcZdXxtn2oI9dhTMtb7Odcd99
VLbfcjoBS1AxFp7ThmTZq6REG4WEM9AhJ0738JGouxIQdHGmYUjpu9i3e+Afdk04
AY87QRM63ox/MEFoj5r6wfaWGGcla3a9+ozu/IJ/1iMpcvI/wXTAwLMPShEBWbOF
gUkCfqjJsEwmF/12akmIbQpJ+GBrSZYhsmzLPs+qRGNcVK1LUQ1G+rfLoCx5sRI4
j/TZokDre6QgSp4ps9kO3bP7fxXBAHPqfcix6TM+IInqeCZ34dUR96eFHL+jprsJ
CTET8cA8omkenqHvn2qP8wOVmKtSEoDc2PA4C/iOuwdtqs2sv+OYCFwrivDBYUcz
AKgEmxFwWLoaWhp0qmJO14TUV/FcSWc3FwTP+VCA0jm2EZShF33NO+Xp3qGmtzgR
YZFgfeTZL8w0qIvHy0ikvesJZQbng5pncfdnLEWDxZxutTsULiEvxwavnZx+AiOn
hiP3MyK56jmiAQS2XgscjmZPA+QQP9iY3sAKZ8pjL6Hh6bYE1L9t6Gt33Lqz/8WD
ElxjP1epmQyg+hXhc/061o/QhSmrQ2HiEuFFiL3dxDp75f3W0Khm5N6GtQU0+TJa
E3zvY30ng5FKo0HtR6ofFgEwN2N3YjspWlwtW0DkFuCd58WQbouMwbZHQp+2kVxk
7bwOu1LoOP8whLmkNcUgjfwrYn1KCFmXpczBeX+hhr/QDyuzvOhcJ3cZ7RkzDdPs
1ta9ad47gCeL8KR9JOBtHK33vIkxoxSJ+ANwGNbO7nNoT+/ouCvSn9q1Nk1oyBVV
7ypOMZV+K6Aoh0+YLlGc9P27AmhktqF4oP4KPzslP7y1nxJ1mP1pm/CaBTfFlnxT
w2SdlU6ZHzaCPLlPgoQYQQ+wYPjIOncpdxWBcwv8zK32gSP6ogL+3xhro3MFtvZt
Py+2np5Rj5gf1x/75KBx7DADCq09FK9Y9lrKBKuWFBTe/4E4SOaGLDi8zgzNFYkS
4OTZx4OYksC+t5UdR99CsG+8NGR89gsvqw6KAshBejJp/gLywRjPzGMr9PLgwIcZ
D2enElD/LaHSWNoF5xpVJz2QEmFPbPXafdUG7o8rCmZCb3zq1x2m3UYLwtu9Zb6d
cfqwuCmeSN9QruOeOmwIjAqv5ZzuK54HozarUKef+eHHFQqDzGmP8QzvcdXVZ9IP
2z5N1KJTC9LvtOs6sncjR2KRzKIs8rl+IWTttcS9zacn/cEWysTY95fM5LjSrlpu
Y+dgAI5Lo27G1pW76q6xFTz3UTAA5zc8b6DvTm7lPvbdsFrE1LBt+RXrnL9j2JSu
FNsEx1n/PxPq3CFjG2w+H+bRcKbolV6nVOqiMEV5hjg+/xgV3GL5iaw8lAq5FXC2
JN0nLj5+4NGcPOUwKtow2A6t4XIa6UtupMUH+hqnfe/PVc3JkvIcYMQ0+iER/WP4
XUxaBQJr0/UguZInyr3it9Bv+1w4jXc9dVdpEJ7+FwGRVV3FjdlwEhi9yw+WD2QO
5RrLKMm3PglngQdKEC+0BtZkhdaZ3NMJoFpiUPE2DwS6YXmZRmtA40GdHZ1kVjxG
eybDwL1hmiaG5VkCTDfm+y64Jsuqj0JIlBVOkqVHX5p1k/v+HJojzFIN7U4o/svG
8P/7Z0uxY83MuyF3+cpDcZORa+BwaIGLWcu8dYvMLvSlqxqI7GiuVRigxfwHOmp7
uuVb3p7WZzZz222ga82WshfOpNsB9lyGA7T2Lqij3Nlbx1t36/Sv926ticBWyAtM
btTYN9iaolseYw80eXTG++hS8siGylGoJ8X3svUijXS1ODSqPQ9M0m183Kdv6lQK
OULMb4VYMiJD2mpe1+wq0CU6dltBBdAxz9X5wOxiFALlLjTvAs0f0ILU821wWshP
3GZqdv+n5lh4D+uTgzHQp1tfKqL/tqdqdXC1OVwsffUb+bdOEM4oxLeAAfhgXC+2
gkK2+s0sHmOVMUL3LVZ2jHvQFStNDt3txzhOOkbHEBuDN0oMfMVQK3OeeYw6GOH5
8HtUpZeOeOcFWoBaBi71HNJD1ZU5/rNNKqqwfmz+h0GPipOM1ic+t+6FfXCpO5ev
ctBITWh5dYHXPLwnZxS0JwUuuJqYOpt4UeA9voK1Vox+R44dMzpaLi+YU/F0CreR
9ePOLYTzyYKEhlMtTP86ZT9CUf8o6Ka3ixI/OmPwJ/P9wk/mz8SYHQnY4lkGiSmU
WkNxEGn0bnYwqOgv7tKHQX3mWRe9xjrvZDixW5ki3IQ2R5S5/3zXhdldu7ZXvxm7
tusz2AbdbCrBFvAzuNaA1jNFTZFpyhQjA7dcQhP/5JrYm7YK4Af58kthSsWLro+E
ATIjhEQgP25XOsZH+giixTiGWJ4lzx3GKt8/p/iW60epr7fmW/XDzSLulb1SrDA1
um2Mpe+MxS+lNBhyptkuoA303s5fmINzZ2TY/Ahq0YClnlVxlsDEkWHinnVWNIoN
9nBwAoA5cH9sF9FcTfeGinvxBDuIaKvVrMOhJgEN53MQ12jt7r42PH2rOILC49z3
loFFCofjnBLQI9IKTv8kIBfyWRBc4E+1MxIqxkKspj8foheQFlRO9eaiSWGr9HEn
iQth4JHUHO7wwciJP6bBVugffPuc7+wSCueNJzBikY9hezzWxpHW0Tp7o4NnmX5T
ahHhNqU47dzillIoeuvNZrF2XId4gXtinyLQqLYUoDpBfCGkyyHNaMn70kBtFfU9
SaXa3Y/Temnnadb9t/PlUdH23fqZUOrHNU3iLE4jCBYeSo+ceDR5tyfQZvqINOAA
ngXNH1xWg50Xz1iQ4FSyc/U6xKZVDqzQVmjqF1FusJZYKWa+lDP8IkhfsKal/rgk
8rSAXEeyKtfi+7/cpq4FmJh3mEjlQ6lPsYjhW00Px7mV00YQuinwIqBmWoSP9Ncu
iI8/w5t4qx3DfliecZiHEDTAXLqcWDreJ52ANdl7SNRMTredlt4KsP0hS9EJN6Bi
vCDXEI38MJtBd7kfi7XBkdQi9BzVgnd1kAuXOpiPxkZ+Ae1HOqHSBMXaDU8/CAug
o0+kohp+Oabo+P5/CANAuw2YXzJKwrdJQCaypmRkSFjTLh5ZgPIA9BgHaX1KTFwj
5UPvNAbIPnfvYn1cBs+WesxnCEzLLVeMJlaEW6a6VLci7KLhF4+GaC8piVj/5vzc
7lAxKn82Fiia6x9SQdj6N2uZcK5qmSKncfKx7ZVTkoI6jv7KhKpAnmLDzKAMJMKx
Fy3yx+7tCmPSlnCO8G8p8lsWJJ3msKmAy6yqyN63pCh9q6uMrY+TEGdN5uoauRhh
+Yu2c+zHqskaJIIFeZl5cXD8oVpiEjZ1KhKJet6SYCwhZaoDmgBtBUiWfCrrp9OT
vuUtRYvBkoKTGCZvS+qTjyIAa/0Uu18qm76ChzNtdmBXltiDJUmiGV5Vfv5T2at2
wn2/hze8Cm4qCvsYxzpo8693Wy34OHeZ1Br9Tt+soRwToR3XSJx0u3GrsGEwi92t
Ypr3sNZhgfHghTxfLlKNX/AfbMtb0cEi3bMehvYEXbwZjmCxR1ots/NyulzOPztQ
HP2nCcAViz7BRe456YEB1F8rBthfc+wwFCOy5HWbPYk92LPTZYGhleLHODL4Pa0B
SXdNJwfVN3Zg/Z71llKsq89ewuCAWjuMgNE8QdQePZ+BVxaUvKuN53fEErWv8QJz
u3++Rt+k6LqObZAhmX0/DUkA8o9FgyDMQpR9YA35zzNE/w+6TGtTFLcX/04ruJwk
7U5hVUDoY1bl6O9LHtJK+VryMKwYKsRnFDvX354Sh0thACEiamu6qI++TmESml8c
xbBGoIRoR0PJC9hT0KnfL4wiK/7Xe42IvJoT2GEcu9KgqB2mjToBkLBKHO6/hxqA
cj7JcU1X2Q/8TPp4PXLoI0YP8hkugcU85n5EM3ap2yIv4krjTi1s5V16RaUOIc8Y
j4cPc8P49Jc2T5po3kqUC9NIu+4uG+C83rZiu8JN6EOXUQP6ZI8pJml2h00iQhkt
5E8T00cwLicBh9EUmiNhPvcHR+1ZAgwWaeGYslY2EFtM/GtwDUFgT9gWy0LSVQ7u
OacUDnlTDQ8rHT/CFlupJDQWatQbkRGcEcbYNFlqwrjY92DpcytjAdEP5F7cRIla
BP9Zu77CRioz+gR0/Sq3DABckV7Tk9vpTWerXB7SjqYiIDbXtiU7MOky7TneVW/F
vkI+7dX5WoYg5tDJQdMqsfy9+3LMZh+n6X0e5wvvrxrmxh5nuDo9lw5yQoxzzt8s
QCLJaXkI0HSRPoTM7fe3oZb15w4efDYsX+cJUuj0fxGaT9+LEk29JBsq3u+vv/3f
ctmx6QtHL0U5rTOCbkpYiEN1CJd4LGJNUyk/0veQv5eDyhoIbnV+y4Ug3xxzSB46
KOqaakC+B2Y5Uow4bDzgJVl1giUUG68pIiWLmk8kAbR2nI/rNRs3fAen6b1ibG94
h0KUEtEWPp3U9i/ivd7k/UE7rYDr5CUryZEHyAMK+wkflbCwtPBSq5cQ44AW04W2
vBLi3G7y7k75B/RdpBR4Nwqdhh7D7wyuiGCJhNAqFf7Or1g5yihF1/17f5fAEQCf
RSFkodoI3kIBfNECUCO0nAXDCc8gVtA6oYy1C96d2EVclwZ+fIvACa0YC8mBg2ss
lTu75GDhx/HbMXBL7VHTw4/oFQYYCkETOWZ1xN+CsPCmhFXyUbCz0JF03pfS93ty
et/vNRi6rH0o3iTh6dsqIGwvEDsITa5s1RO0sXUzDZUVSrfVHH06/2eFAK2u+FQj
FeJl0RFe4U8Z8IzijpX62bVXJ2LZzWFF2fiI/MxhHYipOU3LIMtXrjRC5ikddhge
FnCV22Y1eLHWInQcev+S6RZlKMU6crpeVlAQkvG0y8y3+ZiEa60KQ/czjcxXVsgT
K8pnrI6pqyH2HdU8lwXevZkkojrYGbuFE930Ahqx/Ca225e1eJtJvzPKPdhALESk
Vmh0M9ZYa1D3mckqZ9sEugWd4Bl61titcEubO/O66eMDnz5AQeMbVMC+WO0ai5NJ
u4inRapI15Ydqt8yZoKFsLZbSf4pb9F82oJviORZFCCuSbuKPeqMxX8VZfq8uOe1
FWHJwZyfy42Hb24sO2ujZgl0hqY/y+N8UbAW5qOFyB1lMFB1CKjEGD54DkxsliW6
QpFGBzEjw0aA7rjcgqYWruOdp9etlUEegLgUCaIBemSLw1+nPE9ED+d/GFQKyGp3
6MAZIKVKd4bAVL01SxeCgCHn2hbeLsKYc+93Qi/+LN1TCdhPghEwr/HVaq5QXukt
CdlEPQnZE0qqQRNriSO79H95Laezw7ElTxAEtMXiB/G2WL4/kTFqZerETxPsnadp
Hxc5LQtbaxt3JesEh/OggBqPYOHKRUHZ7yzZyjZ7dCljbV3Z9iH0xs2sO+o9jD0q
CRrgFoeE/nyXSeohh5M+l3+nmZcQT42WtX2gZkX7NGQe78YZ3+ksaLqjox5btEpR
gRQKq+vAaoItDKY7vO7fu6XDzSmdYUAzZv1jc92EA05m8le/W1wPV0ihdGu6ejlj
qmXM6IgKcTnoB0WSwc5+l/yWiPAmedp959kjPaj7UMMn4PS5E2n4m1Rhv7fj+xQY
np25Cz/bu14eOlloVpFg+VAFbt3WjYkgxy+a/CgEm8Y7cRRUO4RoqLCkRjatd+Mn
dpezyGqPKBFAoylCDzl0i19++VSoFcc+zyioeArwFPBfWwmfnYefFwmLRcEslhIa
pu7cRvm7jZ3TgzlbUAOIcGDzPmNwTi/ksACXxt5KRDguCj8LHYy9ElEICTBTHU0t
5OmsEpR58v9ROEIW0uUHni81S0OiJMqL+Dmcz2SBg0urNU733a0CqZAZoX3pC9BA
6xa0HYe696Tx9GGBnQQ1qJlQCRVQrLZhqqGgfU82LisPI+lMnbafCcdav6/PICcD
bTwfJ5ToxkFEom9hINt/heI4a2GqMGXoHRKkZvk8oROdAQHsADTbp2cG55trbr3W
bBBq3DqhNrKtUTDS/+igy8OMK7IV4Ruc2io/releBysu9KMicBHO49I5WkcKjlLj
bB6bqL7KoFmoBVasj3V3LsGYx15uVUi0UYWbF5ev5doESy1c7L1EUHvLKE1e7on0
+ZF0gKy3tZwRf88GBPdldAlgnZplu2oJqDFGMiRJv8+zug4xlzlsV6FeSr7+R/cD
9RTL4Umc1q8KKKw0dq87ax/hG3cRFNcpna6Cj89CXetM/d1q8QempA4XIlL0Mum0
Th+ANPzCr9rwoFjyNIAMrY/+8DDmTFgAhocm3izGd2RGsO5dDkbAnZSRp9zVDdp4
pksXMxcnXPVKWBge7MagvQrfTHtzuLtt/Qy7OKmPwo1kVrbXEVTHzV9WmyFG7dGd
5DzBT3dXMZpQiVbKsMYA0pQPe8sR7M+yEv5ahqwV7u9x4NDgo0Gxa69jRzjmCZwv
VLxtlmTnhhKlmxqN2K2YPi+a2yJ1AbS7IUqaipkvu2B6Fng20l2jfQFcCszrjGjf
tYf17IScfHrdWRiNx/OmXHyjuUuwUFVvjGCm4R1QQ5MOxflK3FSyUbgoiWzjlN91
FoKrB5O9yHoqxNjaDdn/4aMUU6En5x/RtV/80+EErLQxL/gSWU1ojysohLmggcvM
B+/h4R2PzbEfHkBtwruCOmo5yFsIVj7x4j8AmlZ4Q7tZ5PgmuJw+G1ML9d4ypBHF
0JZwDjgmfmGkYfftTwVgQDJSzRnt9Bwyq76+gcrG0wEdYToGRAQbwvZxWJaR6dky
Y6bIU2SrdHcGDmzr9SiFI6/PlOTDZ9V20VT4NJRJiUSzSR4BymaJMn0cXgd3pxdE
mlhJS+xBWTD8u89RxKvRo21k9ETj1/8veB50wOgg9YyuVfeeiUG8p1whaVrCZrVc
OZ4s8ApH2Wp3kSuXEY7tbVYm8Duf71AKMzZaQ4x3VHiEDIYupmxcH9Ob1N0QluNx
T7Z7b96/Vgm64mWp8OMmr+jiJdWHAnuEcKMK3sBsBzaqFdGPHwV2x9HZ1bg3kysp
4KxZPXGuhU7YcqW98pqInZlq7/o7leSq8eM49M2OGE/OCGIHlRdl9BDilduHH95e
Kr2rbZ6tMqeOjuc9AD1RsM6N8GW+Op+QDqiUbvMNiZDUPwD2UPvXFhsvw3dJDbON
ywtG4Y19aaGhwrQQb6Rc/gjJPI+elumKXtIUkngReVh07lVzNKecNyD+f3devBcb
3vyb/PIFOHkpueN76X85/0JQE8KD/zUQ5M3QIwaZu/h/t8TLKsxJXy5AXJVN4mZY
bA1Z5KK+S2Z5kqAvF7tQnS2lOhbwDg2gnqa5vG3W4JN+QEHtG5ppDcTFFtcRIGa5
RXqzv4Gfrs4vLkCLmvOK5vsSlhcTCxUqnL2W3OgwH7NdE49psWfIUv5XL9Yd35Jq
Hd22TC3c9mwdDqQD/tM0/tDXmOG/v0CWd94GXcFW7b4o+XTrWfRTFeA4aY0DQPkD
etrdAxtkWH5QSToUXHlfFnLMwTj4v2kpiq+cQISvSquz1SjGlVwJBg0ckVWBJ4lL
gGK9f7GA1aQcZKbWmbxVkI6A+NIuyOg1MarHuvjmUaE8tln1NCmY8lqXpRW/W4Hg
YTjkEu+BEat4TFhLaLnKiDImBVXsW9NNJWQVNcaebolFLTcSvXYTFJ1khwOL+jTu
o+tSX+mq49AhE47QzU/b2hWt0JIOnhcvfV0Xf+fxlUnxGewdeHdbpsq6kmRhEB1y
Wze43mYaYOq0JzxN7ukFqNlvwSQ/fKGABiQPFg9rShZbh1TLctBVXyhtfK/RZc89
q79qEpCnp25+R99qo2oPrqvk//EbcdpQG++BkqQZCGgJPR5dV4wGGgKKrIOLFmrh
Fj7VMLAE1WEUZW64jG6bMXY5WXAehssaUwDGe5bY7rLDub4HjfiOwmYyTVdYd8xe
U6K3A8TzJUO+iOYw4YED4Xa1bxQ3sEdritnWMqvlH8CwB0O5QtS1uKz4YaJnZMvL
rLX3Pp7/nUe4Zp1LlCJ3+H2naLjgd0UrK3jIdZGUoMFZ8BOR7Et6psZEpzthGBZc
HLZxE8hS2x4vEsV/YpKKLiXKqG8ZlBZEMq6hO1e80LhKayewgxzlHPQEunld82fQ
Rh4a7BE5Z6fq3A7WYPh/vA+b78Nad+h+tM1SDkENrxiit8+YXkoy4fSBkUmvdI2u
0g9/CdknzL2hMo8NzmgnO0Powc9UmSFtve7C9owrWmKE+YHlb7VRoSzkTzz5Qa1E
KI5yGUbE+ukWfydCfgsn4OCf+Y12MpB1K+PgoQ9MpS/DG6/0VT+LqQ7bYpbofrg7
ziZvp2z7ePdcMvS73PU0Wqeuq9Zyy4quHDjilPBpdj1CjjNNCBH8Q9cMe9lVNQXp
Y9wOpBKAbSeQP+D7HpI7BoOZeCMfoKiN2m2xFv6dDonrqnw1F5A8ratGISWtYFDc
HRSehzkovKUNgSZ8vdA8fLskZstvL36YAC6zOGW/f6kLIuRi1viUvSdhCBu2Usa0
g+ijfdTuZ2v7g5RToX2W0PEBOL0Zej6R5FT+a+VoDXzpPgggs4KmIAbiXqxv7bs7
52tPmlAcU3EmZWzrl8ZySrlRAA5624aeQGGDylOfIc/o7mEv9NNQGcES9UQCohp9
v6ZGQp6YP5/niVgGuVqi+trNCYcKuHTU6azlBlYoN3DUiNNooPDw3KJs395UZFfX
O9uGhuvCdbGm5wki4T3M7GOYt9EsO8Y+ornvNnQHz/Nh+X+uzUEt5VLGReXjSlJb
B7/SB+Z7GMv9gmxS4zFtLV8m1e1j8nVzLh1100NIaClvFQvQl7bMdZdxYJlkI5ms
sHIR+PO3MiIYyKrikNidLRr3baD+wQc4Rx4jDqoiYgTbtx8y6Vo683lv1i+9YQ7E
iBRJLaYmn5RzOyXDh/U5xuS331s3xLQHx46QuXuLsJS8inox0znsUoXtPXhGqgBd
pyED3djbdNd7E6s2yDRO/EUxa7r7ka9jsjhVDUPr+nc/YBR9stAg2kSSdpJohiW3
kSGAgQiGvkQw/5vCrc22P/p/RW9FJExey6CkOmOzczq0vRUgAEdXXV/KG179h/G0
w7487TkYNCiVTuYAkzklIwPz3CdmXlMpf6eGMZIiCM29RNYp/BrBfPpynH6Q38Tf
KQIxtto5ZdZocImSxs7AzrDl/CIzOP0ePM29eg+Ib8NK4qInBPi7DWs+a12CPm6N
H5G7StUw4ShL8719YKYStGUHu6/R0b5HUy7+aN8+WKdJOiBYsQ9sIOQBx5CzV/WS
73N14F1zyMfqh1Ybe6MAIdWtDpP0tBS3FXojfbjF6qN3GwBTmMWDPDBgZeI4Uan9
7f2nL56NC3gKcaZuVS8yBP8xERLVaJwcl3zIYEaSYpcXrxa4Qi5C2V9iIDeVc+5H
m5Q6wkQuM+eqJ6HMDxr6qY0R6fQscEewJvobuUVIgnmTO5Ym26TgG13BNkIP+CXy
lNFHQAIbEnoaqL06YJsCIcGG+v/F+JdRLuItmsSQ25zOkfIaYxVgTae6A61ZFA+l
9xUlNXZZF2EVhth1FIl//rIRlwmkIHC8iB1nVbQs7rphaQnhWwXYzeuY/UYTHMa/
3muV09x2jXTXW8IFEW3tZMrwzs934LcQIVtMpCCScYxPEjyTsR6zyQjwQsgWU628
uDGv86hfjR83598j7/cXw77z2Cee/Iz4lMvOn5seuWIpsBPNsMrK5Hi+aizqA3HA
b4AVjvfD0I60LdGqys8jPYGJeHXWu0j/oBj96ADRdQXOB1kkLn7DfPX5wLjV2Z8D
YWeH28zJ/jWcpAHnsU9zSwAAreD0NVtvsfOvkisN4ExWL/2eqOLa0sQ5bOg+WKeJ
3eQp9M+oOvX/cgPt9Ehylg5QGhWzpviJP5m8oGLTBlt5/Vig4o+V5f5vrKDztyxn
uVRx0mSu82JeKeUXaPBpq2Q6Jc+BkOzfzvxs7K9RCmGVgQqzkIaYahmxSFoHKqY3
aQnYCgqDi4mKM9KrBXq+jEhe+wjH6FbVg0vuVTJqURU+zI9uS+JQvJhL+eES0y1c
PbrvLmZhOcm25MQAwNIBlppc7vCnsftOpWKBhQFhUYdeb6MSNIfmXSVPKRBhNzb0
sKA/zA5TG/YuFeNzvCXHvwMHIonysZXxyP6kZuiwAPxpCx4/dRIIzvHupPpCR78E
5iN6b2vCaJ/5MObP23faO7+owolwmZGD1KJFxvPa7MXnrNAV7zzrmCHpH8UF4ppG
BR+jzs8xG+U3XuOtbjAHiS4VR2/h/lPTbRew0DVPNQU+IhBt/mJV22/Ul9wItbjP
FWCoPyNuGAG5fCCtxjOeFHoRh/GnSBoo0G6L3Ey7A+ZXGGdfyJW/aLLBiHLFKS4V
3V0HqVrx24+VME/cbzB/gH6yoWij8BoRMPeER6DGj9GNehurDzVkXtxIpnLYE+LH
G5Vzc8CcNWGbNI/FLoVaqyzhZaomGxO4VzGntxyDuXHtI8CZuk/6CnKRSmleVY+1
xnKZeeWLcxEfODYQlWlXqmLPil4KB+oeoBpFflYcd1uLwixhuRljWCPwUaEvIOpt
asr7VNJdmnGkEOO0gd7SctyahocrRkiDEDmhWBg59atS10ORWVBXiF/4V/S9zZnk
ngSCBLItUtOx5tHZtyuOm20Z7UDwkv6sD2+OjY2uK5jxs6OI7HzqosXwXrtg1WzY
c/AyOTDbBWvH9N6Gt51wfdZhmBxOyoZdLJygNyVOfOYoyW+eHngxcggf9SULFguP
mBMtlWqUeHjb846jClizP9R61EBnEoChAOCE+o92jN/D13Olc73eNHhK8+BSTl5Q
IIZepRx/rmhoLyfzIh84MByUInwtWocZwazchvdAoUOkR+adOz6SydDZBW/dS4sS
w0IuJi2c5FZ6VsLGuqUSPfVao9gODpxhyHpEFvmlMl2dIE2G+K7WqeNkDFxCbFvI
DQUD9MjIjlEbeQTZBsSk5XbHivWolGGIrc7WvNy51QBiRHP7vL3A+uyG66+DGThF
gtBb407WCXeLCCQqqVmD/i5tUpnL719YDQP3uud8lbrhZ32UXjptx6K4M+96rdDc
HYfUlkvrqa9Nnq2sBE6uRBKXjwU6NMN31yRYU9DEhWUGJiApaBJ81brJN/G7eWTm
Q8M/VR3/+ZYzAsvS/dq4ZsDmYME/BxSmsR9QhYuIrf3X9bKqEwPf0NQLsPnGpDfy
fII13aMRKDRDI3fupJ5uw0JQklKSgnUIdf6U8LCDs6XpFXIn1jfINj3zrMHA5Knz
evem0+xvH70MJp9EdRQRQDLVrjFzslRXmv8hlVqZysDKgOY+E4kdcD3vaaoyVQc9
57ku394/QUpmXz29BHDx7n/oWOSKAafl3yoNA2fQyyP3rLZjvxFRkVUwinzwZ9TI
xF+P0ZEhM15e0wB+kU9lq9hsDEME7gvarTRNPHgyzm9ojgH4a+a2Ez4/EAVkAjEI
5stxYt3XBJvFf57PvaoDykZfwl2F8/LY7OltuBAVDl/RPxHDQ6CPwEToeyJdeNkz
gTYoHi+DaOVtIDpvorqcu/6Hh4El3cAnfX2MJS3CA9tmBO60o2nfQ8URMbJzavif
4OZyks/v13vhqRgTpc0BTXYQ66Tm8jiSWWcVwcDLIYy0LxB/e6yBonlXHRPLkvSb
yos585fg+iVwNVh34hfCRhxfWDADRmqSKl6BOrMMxIt31ylCqE5XKkQfoiAN/ysL
KeTjkb+tzad74OhW/EKDAuCkGeFQ8c88ObBNZZlYzI1jw9714XlCLGyhsx3KlmZy
CmmWgf0ZPUC053PFn0DmNlc6eZ/zYCn8GQcRJp9zNRhEZPIc7LJIG/xG8SBGkqZc
UO5nlsE4OnOjT9x1eLiEeqxpJ1G8j2QPMwJKUjR3LBOnGMakgWG5kbi/R8c5SsPu
hQPFOdQGyMbmLZ95G56+d1FaAgKv0IO2hsH3Ygrmx2Php4KiykelAAWqNe4MLjIw
pWOsa3kZkh6PihqjA+/DcMz9fG+/ALOzVcnOYXsIQaeTtiXOoDvmYVnwjXsEtq4D
Tp/aErGedpUPX9UzytjJlFwBMlPKuq+KJsEfvhXblxlwD7g6+dzPMtlSJ79CB0Yb
kKrAf4Xj9zSrhyoE6MEwbNA7P9udWoKWjDeSuxEDDSvtsLN4OO+Auhtn2iRZr0Qz
ojJHGANZd0GjFykW5/CK9N4XH3GeBY63yCY/85F0KfeZG+VTzjg9nFBI5PB8mr/Z
hIggKm76/a/K97JWdw/bnEE5gf1Bc81JjUKXw87ZBxCPm+yJ6hTiycWSHb8Ymati
N0wSzr922wcBUit7IMBC/zQb+ZtCsSJzmbEJzTccV+5b8/Ytv+OEVb1+sPJN3ClL
RuFtWBBExDV3I1ex5tbWDkR1AJZSFRLZedKoquDrO2/HLslaTw36SAMzxs6mX9nf
Fi/HBamOi0Q6/FU9hQg5eXSTa08+0Dm0bWFpRYdRvY6YOKr+v/w3kl6LdDJRgKYk
u4+YhCp+QBBPqiKijz9nzkaFKEIDm4TRuitLmKuTPVOISM5nKJNIUc69iiltXo9R
8v9BfXMpRIo86gvW2l/YBoIAZHJy0QSEfQQk9BS/ElTs9aJm2M9Ekpa8GNtWzIqK
rFyacildSmZgI2UBJm9kBMqmavKmgxFqd6+l+hyBDYrTUYkrG1QsmD0Jl7LdvffN
sFU77qaN/MuA4c6uwN0JxFEAsYjlAqd94GDBNbU+NOYAb6/PcHTLXOXLICIzWUMe
J9Usdd/VWTHVrc9hdJ2R3v1dgZnRztIkLvtCdaimOKH3aln+4ygcI6VnaRbr5yaz
Kye8ca2Ut9qbE+PgCN1fUj6l2DxWiGkA3/3WQql7No6q3vQah4RIvjLQx6rWy7T1
0biMNcTP7dojiE/uo9U2MJs+hECabJjhqY9TPWdmgajWjfOmIYydLsl1KtU1FEs3
Z2wfU/puPwHdZN0U5kfDPtVcXatkF8a0ZIH6x3F4bTVChFQiCuDNoTqojdD4dttb
SSfWhsc7zoFPabZdSg7N+fXxzZLRKc2nGs+OZu1F/gPRdxwf56wJX4FiECSElv1C
f1fnC2idz0rgqZm8LA9KLHfpijA1QYZttLXpngsYPpZUso+B5OMwkA6ND3aQiwUP
o2ctFE4ZMKbYvTRuOkL16lcOcJhjl0KkoR8sfdY1Rcm/IP1XcYadUNxoBdxXL9Z2
x+bUFoklbGhzleAzmhN+ebryIgz2UT5MVUrlRDzaEd+UZZWL0rHHn4rLRbRhn/B4
QXlBV2HJZd2tFcIfAlTTz9CZydJDvYmsdFkBPf+RX0RD0rNY54yRnRr28YR6Cw4J
Xtlpi0dx/G7vH3PCkLJRt9UnwCpf6FZmPvQaMVQJErVx+dREyr6oxt8LO6XNn1Zb
gh6PZUMsC5PRDKGByg0nytwRzzVyB8c5Vm3BS+QK1Z0T0HiCZLfwpVshYc7Sipgq
x0L+aNA1fxQsIWuX2g2D9cJTxJQKQqZ/ugSb1xEJX/17bF187KlQ5T34c+cHPWuC
V+IOXmwhd1nzg+7V/J4NFbGDXrAhLb+v2NxXFFPVYZZ1oNt99QzTsXC2fM0Bdg0K
qINRKs44mqLoDdvF41U10OoejUmawhby8G0GQt61yhi3AIS9kntCa8bORCh5NwuR
KrV1G150zVMQ+KluFUtTQUNrUc8CCNq/00Hy1UTV3rmmeTRvor+S/a4et68AhH1G
WGjONfdP9GWSMBZvxQytBT8OqePxRFEWEO0hDApkifV0O2RpZ/6AvCYR1AWeGEYF
GzFOFHZOBeh1822lolR3YFnggBGTuFQA7IFUk8o02zCr76Cvl3yEiPgb3L2V7faI
PduSJsbg4B2V7kZPIwHN0uN5OIuNz/5anJlPRTj0s9wIvboKsDeS/WleeC75mDr5
LCXjAPKmkPRbKu4k6Ovbv6CQNN4/JDeKD+4p6O+2g5+UxgpUF3tJ3GLR7/Cw82dO
RXVD4pgsy584KDf1veamSf9oqfVy4HI54HOafllIGEwHR23yeH80ST9XK8jMhSIT
rYS893mEHhrhHJUW3MQ/vbhAMo2UVxbIasQFcbK02Bo+45YHahcnGa+ctu1SUzTn
lQRYod3k13+fBh0a7QdUe1T2ISAOSomKcHmMHs39Q1kwiGbL18SONCOjFew7rWh+
ExnuZT8RzQmtt5cpA/EQjUPQ+QZHvSKU0Qjv70ygmT8SPZSP5Hxthr/0wlSjVi08
JZrU4+ex9JaCG0f8qpdjlB1tpxBWO38xjjLc9aja+CvdcRgRqNxE/ZXC3tgxoSYW
IQsgjbjqnDPJCn0VOFjaChSFUNmK7X9iF98RktUc8IJUaDGecJJHn8OWOze+ZyZi
Q2xPKQy2GGQQuhtcbQUQ1+czjE4Phsv2NW7FgEpLc4ervFwy3yXlYkIlt+d5rRw6
jEvfPrBuMdar/fyD2ROYmGGyMumaxY1zcr/ulmx+5HBVjeVwKY0TalUJIDpCXb2m
iJPIe64JOcNAhB6b1nA1bIEOJ/q72zszicKaXmsile3P6P9dxduxcUJBTg3rQ6SD
hPRsuhO07TRdVLTTp0HjKnFwF2IIad4UY4LWC08bxfHQZlgsgv+HVfZsG83U3xQS
/Ua1JsA/n7FSqhSxp4LosZlVn19cC+DJvOoY8LFv7w+ZGPTIeZSs22Uk7lncd4qP
eyLXdjuLXE7GSXD4dD+USobVz93dHz02lABg1ez51RzE2/muYkS+jGD6ShkM5X3v
Ep/XFJJquJalbVUhEVxGZMF3iIG4/xlCrGmo9fNzwaxy/6V1KaiZsieTOYPiGWLR
GX12oboBKJ1ItxX7dXPZZadwLN4z9P5BqlufXOciVFuCwQF3/kOEV2hk5shELOXH
qNsaipxXJosTcqwCYS82AFDYsm9V0k7BHOYUdVEZ4sCL447QGatixpYdXk3bU3+u
fO2PvREY4oNY29bCL+nuHGTS+4S52NDGd88iftd+xx2D+QguBVLT35Y+HVtvlEQD
6E3A4S0oba2+NtZE6KTdwAJ41T4HsHtCFc6bKcQDlrBNiTPeicmBYyUTWmVL+Vfb
/b4aqsns7pe150cvSOk5L7AIvgMVcb8Mn4W2vcMGWALdIgwJEONy2YE3W4NaYy31
iDTt+e3cr3Buyrj5Z6VABfvMGFSOcA9qwYT/TqHEoeHL94hNo48vJ10uOonbRTss
QyvgNSjylsAgxCCslOJBpIXl8uS2aDMEN+s0mogiREuYAA3AU7gF1pC/5yGlyq9Y
8KMPu7mxaqNULO1xJgCu0FIbYJ76ef5c6tviU+JVN9IoBn5CxKaHYT5s8NBEw4Dj
3JdW7Rrgeg8quUe+Is5Zt0E13nA3j6DvbWaFein6j9/IpzjD7Li4+0Uwe9BNmPur
iNKRfKrOwR6W+doeQJ3FTHgJKaKrO0HrQTTcA90O5zaVnqhd37eMqeKsA3BNOrEN
XZgbUEMPLUILik9jdEChxKBi6/CgPGCgt1zyjxBn5ZHOt5BzLgwIYuOR85d25VjT
CjxkBKMALqBoXWryb1H4S1JqUAlIQEClK0YpjJhU86V86y4LoX+qfBmRiLGMAELx
lLz8g6yVyqWXCIT+wuT+X9wTBOZxEhEEyneWlF2PBa5xdmVVxHZ85wYZDzMqqwpC
iXbo6PQ7wz/4tdOwxLimpFialj/c5jcGTWAdkLnEyNGm+3Jxxp+AFvSA7uyStegd
OEGyNKRrTiFJOmD8wkSjNa9gLIQ7kTKAU6fSg536pdVkSknWuzPmTetly5834UJd
Fl3CJepjXv+VRJW/j8uItDXbgTbmSZzj36PCxTSZNjcz/vRPe/V25LROUFzbfk5z
5pqOykoejeRkqYGKHEcJlTB5jvHtZ0v+FQ+UJ8jCvhaTanEzKYp0poijjvdIVBKt
brYjTmUJEykj5VpMPDDFlRYMBS6oL0/gyn8OFnY5K8cFzOLhFi5L5Udwl+nB1Jb9
FhHxHyT3eJgRaT34DdA3lDponc/vCj7y1eA4qfiOIGxJQOUEySG6WWrMmImpadTW
4HJVeWGvwwDdleOOtW7vCv3nzajMzkM5OrQGzt9MZzQvRgBCJKwAjox00ggb5wWy
RHOzoNkUfO+NqD3lj0UM7/Qd+NEBY2jLCX2tUhd51s5jts9zFMiypVeDI9Beq5od
rAZxvzjIhiEDZTCVAlB9xCLzMnsFhBllhGyLqD67IwGziV4GXia2VHJ+wAj+wu2/
4tu+hh+QESs/3fwgxPktSw9AVAsPnId251/eoGQdWOJhvblehL95r9bcwDoZzlyE
zM2a8DZ623Lbdj2Bdlyh29xqI27GfeY8aZogC/BjIgPkehrxQyDYYRLAHvOXSzyI
8MeQJk7LZc5PGzvM7cA+3mCaNvBwt82EXFNQ3L22s1lAqlcg9Hg5o0BbmvdgEuva
XNQlLCcrO0d8jFqsrj4BhxM/cDjZN+mrD21TVTnpazFrFgmlr7Gl+UiQ2FfgBXSY
Xuf7vtE8VvBzdE0S0NI4+JAA+6I0yNOcV3tP28Kxgz1k55Dhpc3Ttn76GqAeWk5k
gvuZ+TKzHswQWYa/v7AofYiB2o71dGoh7YlwaI+t5fQxAHrU53NrsodbeQg2nJBI
8rzMaDmZg+pj0KplqCGUq7FPOJplmMxiz4O8LSdpMZn0ltPf3IxbVxuX/ofXEnbU
6TCSqjESy4hXmO6iY0Sbx3lVVouIT+9RCmVIYa81CG9snhV8N5NUJDYweImBdZLF
YvN467zkxU+qD+/eov4VSE7/OGi0FEEfV9Chhh6oA4LGYwU2/pdDXueN/2p52M3p
IIVlrbWSrb434xLI3G1pgdaRdTqn+nfYNekvv1AUhQnTD2XQz+xxHIM1XAthRJA2
skobxbJm/1jduYOCT5xmXFlOpCn0SWX4PKRQkgjvJUIcCzCTrkCHRSOuBrPcxe0o
EF1m4xMNkPWqS65sxSUepCMrY/jGlfxFaEYKXCccwi/D9mRnSh5hlZ9KlhHQdZF4
qiR/FbyiCG0j3frVnS51nRZK05Ous60+UR3EKlnqXgLh2kodC+lH9Xi7MxMVeK4T
YTlNEE224fhntfnjUwBOZ/qPXQ/Ck9Dpvtr3caxgp/mgEjsRjHQY+NT080WxfSsB
8q1VhQAJn43gO3iNwIUQ6851/gnQehnUJRdPt6OAhKzSqPFDEhkkqdUmIb9azD7F
JSUdmL2heKZ4zeo2r922L3VkXX/25X3pwBRRSL+ui54w89S/cpSgHi54RKr7Li9X
n17rg+aLmnrr0teDAx+oRnlW4ZeAwcrx3i4M6XKiiffqTQ6h/MoPpEMvv7s9K8Mb
33oSSQdt10mn3xYot2kEnNyjW8EYi4KPA/5QG+V/t/XgablQ92Bv/SFGcm+zHkKP
Q3/tve06BriMSeza4W7WPn5TbxUxZacKLD8klY+DSfRBbYHKVE+fjtYnuiuK2Rkh
S7jV+kniPyQ0AhDBkvugKk+3HwQdyXyKdaCmLa0vX/8GOtnHRffY6Bp/z8gGfnf/
snEiTsHqx9js/9iQbHQDOmCbTkmAr6Je8Yd7No99n1t8zFTxPfjYQ+5IGt3Hl/jl
Dife4rkmh4pvi2yn1B9Qm2SEmg/3BiJ4thz/Jw7jpwSUobiw7s51j+LnOrZa5Yd/
TMl9ojqjj7WFnJQqdbM8oyTQWsXX2dP5dbACwV2ygpJ4WUOy/vyamF4wdIkGgcIr
3OoXIkEtAVzt7KTqM8zw44vQmc8ZZWC9UtCkN7O56g7t4xTZyiGrN9epL6UzBtOI
Dl/XhZnJEKjwcGyAGAEb7cSceNEpOffpC+xnD87m7ohEJ9/FLmdZEezfRLiUEhpv
ozpt3lNsNFI2CTeKszB5m4TDfqyWcSEbCAMefmL2iYqnBWf4fp84rpwU4JmyM1hZ
7Mb16NysLX/npOGApHkcIN2Hc2Rv6ESPNvRErsGlBdvquA5kfaPHYTlyjLiTK//Y
PQ0T+svSJX8k4SyvUqJKWgsb9nAMlFsJGg4zX9jsxDJw682yccFyG6lvcaQZ0E3e
ma4Jfuz2GJqdEtDv5YY0sSt4MlY4vc9JPn54pBqVdzx/nUKY3Euqo6M1xu1YNM/Q
ws0+f1lDlX7eWs4Du3lpN5dxegexGt44DEDZ7cbxyVopthqC0sdSAIMXzWGzSzYJ
gE1r/FSBfaVy3dUwabJ5vwe2u2yYgOLirwCUnTZOkg9yKdKiqjq9mQCuCXQD2zjm
mW14mi+ypBifGClCp7VZuqhID2dXUdeEFur1pTLinCH3JZEjpHvAJnAheL8vk4mE
VRp/V7+Z2Uem4rAIrXZ4SoFwBM6g/vtgqZKBmNoAa1jFvTxMsXAOlXTALGad0/2z
7Jwp2C9P9NUYbnCxCZ55GwbZjgG27JsAjePovKw6/grd9A9oIYCwrCYjcu7yBZE1
95XwXU2P8QQhdHJLfUK/lghT2A5nsnCc95HQqpk5sNpxzc8z4F/jFqkSBLGr/sCl
Cj7OahLnZ99SkL1EcP2XdqyAYhFMCadoXjxOiI35MqtznYPLEPLefITqwm+VRUvW
7hje2BY088e5wj4lR+FFrCtaNz/6nCCwRr+zISN0NYIN2NnL1meZKzswrj0viaxC
djz1Un4pY2MevNvIB+FfB66rop8Hg7OAO7NfeQkZB662Alh29WPOogLnB+kv/Om+
xWFp9gPbDtQSgPafLTgFcRJJNQe3g1+ZJHWUKz1Hp7Ddxw2wSawREs9BSzoRgoTT
YDNffDMGQfv0BkQgK+2+j8Bv60CUiFshKSP142XSROb0STBVvVL8C7MTKTx6GfLK
+2az+v5GBl9S9LRJdyzm7dWeeEeV/nz+MydmoFldX/TDIp5ctzT5f7hCr1y/sWoh
WnFFCTzhhO06GMwtxi+zmQCzXOI02ap3LhXXFOD+6VnhqQEzlGCJOm6XTxkN6YAg
SoN9f1qwqrhyHQVBR0nYMAIFHPXuy9TuTlIuKg4pDmgY6HhdQpG3ALNDEKtrSP8c
0gX9VeJyTStzXKSigbmXMdejHNdy0N3U2vrcv19SpZw/PZhnlDVDgOtcccFHPlyk
Tu7I+UNbT3o14wKOuqXCXArA20b89ht/K1cGNbNgermSgu6HDSbfy+KxaYVO7774
ycWvHLRBKRp17qwP2bEDRsqQFs9XVV88G02IBbl5c42NR3BFJ46FSIzNziJHVlCr
hESp2GGsnv0R9cPIj5j1d1nKYh9alHFKVjpzLk8ntCRSb9eoHLtuzdJ0H4ThXlf9
3H+gUY6F+8qOt10OEe/dQYmuGKg5GaxJ9d6xTpUzC15yGRsyK2K6K+ol+e1Bc4RW
FAhBNGSwY5zIwDLaBr9bXUGnjNxPfLrh+dBJnCctJuZB4DqwwLqkUawAFBpu1vdG
QMB7+oxPDJJXjvblXiZdJmEWFqD6Y+Wl6rPAcYcPiKaEv/CGB287SZr4qUL6Uiai
WrxzGjGvabh4RcpJ6phFaJBAQ8bDi79jjhPKPRgfBBh38o3bzrI+OXEu2oB2KP1t
t8Q2P25u4B6XwQoLeM/CLwSR5/8Fj5HmFovvnbpChKnJ6Gz8iiqMKE6z8F37u+5V
2t+Z1Cp2dCbxR+k5muU2l+aI9onktsXLkYI4SrS401G2XyOIAD2a9jdA/7WyhU6A
YL6QTHqzy80H7WIS5j/jreZoJpp5GbxIqDQCr5WKI4igBdaeRoh3BxoMIuJVc6K+
oKjrnAW5vpCT/WZS4x0c6wcHPuE4cyQH26VUM8svU4K3w87ZeluYezB9ZHC6yB+K
fLEKx3ICbbDIo43JZzNLS9hnJcOq/jvxxp7KGCAsQ4vqJ3VPRqVUL0SUt0R6tSXi
4cRGd2Lx+eVx2/Cmd0G5ylVXtDZbSVfbrNnYy6FAIxkDZvhddDc4QhGb/j5i7I4w
o+wuGJhsAfZ9C612p5oKXvpIHfg214FfraXwuSzyrN+LcMh47Dsvhs7oS+LHxUGF
xantWFRSzlhdXCnrGagJCllsF1e9KCrxsFMx8rWValMlVxYkYU20qpC27DN9+nGS
iOh0xilN41M8nhLRTKaZ4uq7vRrJh6eZT83P8y77242S0gqgVWF+IheRdFCaPo8N
RUGw9nKuaahwaELOQ7EOtcGX2qD9JbQPWbdsK2IAqcPMijsESMSF6g37iXnjS3vN
HU0qQUaQi+s4Osx9zsg9KPGDCkuWtATXTAiCmu3nBXfd3GM0YoFfSxfvhhnUemk1
2KqSGZEXTwpLFj9LCsoaKotpdXse2SItzIC566uuSQwteOQfRwTwqaWq09Wihqk5
S84QQY3li/IGrew1275aQhATJ23v4RZ3s74qnbr6F9ysJBSWuS8FviDldJpM8JbZ
2UF5Hai6Z/xa3/IofdWfydmQk7AwkDY/O02kCp5t6aVzuf/iJMfVmNBrV6hQ0f7u
gutknzp16CW+V2cuUKGzwDrpBtQ6xab+gCw4nrI9jIxj3Kt4+XN1GlJSCFapTzR6
guWBgIWBGkZsBOhaqCxqdUEFOZhI6VdnsdzU1f/duiz3zyTt/ynyqJufy4nejSVN
u+uNlZ1dvUZ+aAXdB/K4nPtVZpJ4D9M2nyoAtLhuE6/pHhRgj/xJl0l9MgJcEat0
7ua0nnpZG+Q9U/a7byRmo2ZXFCrt2NktMp89k/HIOWPaYnM7akeh+kDJG0RbDCUy
Px0+FOTEpIOKI9ZKNqfkImIEQ4UFVFBRaiJB8oY+ZKSm+lJGvreIdA6D7fLB+gIt
2orFoDQ8r5yOXGjf7U0OY+7opuT0JfHuaWOW2pDVEQ7uBpBnKYWc8jNuEJ9cfDZg
7CZQI2sG4KhJdElGEffJ25BSMhg5rf8/rHyyb/XDcQTKsEJEuI+9ODI9xjBFezVy
RI5AMhfpVMHuu6lxx0nCeC3CdDgVzS7TSvvI4aGwcj0fJb+WKHPPCX5RYUFDKWnO
x3Jh7yDKVxB9HW+RNj/lSef6bVJWMW1lFDNUjdgNxtr056PHCC2H1uv3HeIzMVAD
3C2LNmwocS2lkkZOeXYeLxO05bgOAFeyjB3EUA4PhIhzFMDLSu9D2wCpKrKBVBL2
QyUTQr2NDjzsba24wEh8E8EOgNCR6PlzGf5opZeNzRgDJWGh2VQfstX7+u68Brzz
SF9Xf7oGJtMVl1B5YCwNuO6LwMX+WCqoXZhfVguSFVjBUCG5YgjBcRpbQM0olhB/
PMlOJyNmyy5HARXIpyWbxS9WSRsy8PdBY/4EU3inI7esqxBcMCBCwX+hTbbNad9M
Bp1KcxOUINNeqGQ2I6PvEtEiyO5p8X6ZJ7mnpoMkJJk1g7MVtPAdxr2egLmaMHwU
Z7RVTSzzpPIoxI9tbs45D/ZhLsdFtAT+t9JN6R29+t70rgMz7kr3UUCcAOFkAJgK
PaVgs8WBVy03Sh2d0K6mXAk5/cxcPyvNqOjhpNARqXgGSyjQcivw12yV4JV5nkJ6
PmCwYLkcEtDFJGYsCQ2qgXwzD1YRdhbqnwDDHWfiGhOd3VfoEF/Puy0KWu/+fUck
H2WDmroUqjmnm0yVgnBl5GJYcKbwAxH4FLe3z7I7TGYxiBuYQJH3KO3sJhe+41xw
NEcR51NIyZvRctzebn5R7BpQz1VtZ9fAGNsZ0m0BmRsddaajvV6EwSDTwRPzGtlX
BD0ilYglvxzoxAPJLIAvMgMOZuN7NuqjByymYmHN8N6mHlk2pQGFsNp2+XvLvmhT
sMeSpzMWktTnWQaAvxCdZkoe0SMIX2an0vf+TxmFyQc3t4ZkLxEPvwm2sK4+KIi0
zGect1wXu4GeWAFxZsec3yb/oWqtCLdOgHKNLTdMUWFTSBYnVgMtgSrdWjLXqY4i
WP0tcvcnPxlWLh4eE5iIQ2RRFweWykLhs2s6HIyDwkZqUY3kqbH/UkhBsHP/bJOc
T0gVQChSPopYkqGeSsZ5qZcygP5CrLqKVjYRbqHjQqKvqPSD09eYxYMDSHqY8P4A
226s7XaiibgeI3WrM8t92sUFFcvLcTJ2Wrlu+IO6sRic6HVNM0WflKZsyeCb8uDX
iSsg7SxiS5vxzZlY4NbWPt+n/pt7xzeuzM+YhO52s7hNsIIz23coNu3L4fKEbZkk
STB0u002G1O6ykaftIX2F7x8HqUc6Wc5eWxg2fZCLGAa7fb/olQiH6be0Mvv0/Hx
29bBVeCob9nby+10W0XTBfOklB+uuDkwfUDpjvFDeI33xauSMtTOdYNRZy+E0cug
2AT48aID1VkOR1w8WQYmf8gvm3nhJRp9psrJStwDgOyzEzheVPdGRRQOmuCxDu0n
SZWiRHop0RQ3LHpbJvT4EX7njAbGEj44vi19pWXdV5iBz6HR7ThWJMlfZtaPVObc
nqNKb7G4i/qGIdFWG7Z+ofDBPMdXCdBYJHbcKL9Vn6JsrYdJd7fN2FVbK+nJE7eL
kU7X6CP5HSQJAr4JZhC1eJUcPjuxHK2HTw5iIJBNyQGibHrCuopshYWJ2Wh3CSDG
wOC7qFCpQdk9agKWLgfUB24EdvGF25jzpE/8pnQucM2ds0nyuhP71QZHq4upwUwT
Vm3RYAUuY7viRSAbGfW3TOZn/6nFHE0JhjxZlhqMY1W/nQdH9RrutiMjyigIKj7m
xZ+m8d8vSQMbfbAKWHDQKA6dHgO2nXgDtivDmAONyQPCfdIgtt1hOCRmQBP0JFkW
UBygCSGyCnemeGJ6/LVZ5+jDYmjG4rS1C5jRG4oKIufzi+XGk8RXRmecG8dcRJLQ
TujNqLEaBQl/k7ip8AqpDOFaqzVxAUxXuF9u7TeXYTIKfW/NtrgMQE95klNIo8LZ
+9wJpF9OpiQsetsIWjjbEEMAGp2ZaaN5N2teP+uRTRgNR3829f+NVTauDbXYnjuf
LYg2VKS3edeQM9CH5fdndt2fnSM/W8OicfrpdDN2IkqYS8VjxkpnNzHXxLTyjZq3
/7U2TvF02sJjLSCwmrt2A+7ocJfeGGMXLXGLRQf3POXycsttksn5rWr7pQFp5MM7
LhuWvpu2bLrq1BhAXlL5/jD2410r1CDq/ULO0eG9atJqudDrY3HFgmnYWP2isJlZ
1ccOAT1zh7iuSXoPXniI7hHO03NTE5qMxJzEcocNJlP6qFK+v7Ygl8C7H4bNXtZ1
ibhL98domQnixnr60rG8S2HcVVvaSH6hoJiepCQ5m/hlpyYJnlZNFvE7SPXhKT9g
idknz4iTEmCWEU2ACT8MFTJ6jhZgKeREfmUCvFluvwLrvTlPjDEc0R5XN408yx+F
VCHaxKYrZlkzEVwXV0/JnPpJlA6MDwzl++8lmVuQ60+qct6/Cgaau9E5c+zyEr1u
Un8gE8090d0b8YEGWPfTDqzfQO1UkwaE4V8x1atXC6Zoufa1hxuKZxY93TCLi7B3
opNF0m4EP4M46uoSeaoAmuX02xc7f7KG2/zPNzdTQcsJQb8MwT+OEfqq1lGxjW61
X+TfWPPXT0A0cb9vd1F6IbY+JiBm07PNbTVrjucOCuCJAaPm908ntswOkOtHZ4Eh
LX6eqqMH8eWDCil+e3/+cpzyP7r7EiayQfJT3fOGqznKFVbzGLhzwVbpYxtt7qaz
jLh6yFd+g9oHnwXk4h+wMkBHpsV9AtTgF7h+LibiSXBRpHGTFbpmgDWnPz2MOaak
t10E2Y6NWwYEfvecHFH9uXbCZxIZ2IdDbOk0xROQK/KoyQ7/izbdDa1EFLDS6hEn
v2nL4wcdDaZW7iaLO2B012xTRsmwi62iAG8JvL7zY7y/dnoSAXpYHy0VCeYgCZcp
rUJgMcx4XjdqPDQcMTxkMvTD25glhk8ltLQwYrNPNj5SmDzC+8nHcTppKP6Y4Kh8
XsI4thkxjx06RknVU8r0pMHwSCWbYlub5jqbkQReoVBaeZFqYW1SiTIOmibaWE/y
3q63Ha1tuBic5PROwGI/3eKPx7CheNouOepFEJMxbS6OU/+6+gMdfmkFdOJ/o3nA
pJlBV46EPVZgwL0SSS8VKHtVKdjLOtI9TJn7ZcQMm5ZOlxruos6gmBfzqI2OWAu/
xZ6ty0lnSKOm2kd0xvqs8xBE9ex63oMmqt9tsZLplixUycTxBpMFV1Ejxx6lM5e0
cP2OJOaGEFo5Rdb8TxgOo9N4JreEaUqIr40ZM//PiRVn3bLuJy/KkYvWHg48OgSB
ZPt33+h2X3RF4Z8Hzct8pAgF3Ds7VctB3ktXSJ1/tfa4qCrm70J3PAlYmLkcMU1g
iYhX7D/NFkPBm9ppDXGApmGEve6p1Pqh/v68Cs7x3DZDfUTa8MEMV9OzZOnihHTj
Gr39A/FtmsYxr7MO9GGul7IgvF8scT8nfG2jEARCg3ywMvnKHBhfZkltwt7hKniC
OMRrSixSOJjYBssWFXUkvs6jXXbd17nau3jM5nZIDjNkzjCBwG5Ld+SF2+UFBrfT
ETKhvLSm0boSEkHiXaIxIdwP34mRtwXTN9NJyRB0ixfiHKc5KVg2mApIQUfhAMqf
X928qi/LI8JMc03BTFf52aXwzngScASQ2St568QfSCYSSAt8G0ZaIX68lD8o2NHq
NV6ZKY+JieV1Qo2UR5B2o+LrY5Eqbff5nkQnSFjgKunEJ6dxvho9rCaEMogJzsG7
ara7xLGCyS2L+y8GsXmVI9jSQVbhjUPRLQ9rSpzlkl2EVyI3sW6UrgVsggJ8EUCI
bCI2srtZ6f8Szw2lmzbL6ejZh+xsTDAW6JQ+ruAPN3F97N1zAGLLGrRvRExFSWOQ
KL2OE2IpVrmRv+RQBAHw8CBeTeGHdubPv6Qv+WOgVncBx5smx0wsxZN6CHEkNWMC
bq/tHIlidQX/Dp594o4o6fLoV20PoVshnJPeP8ZUs4s5veBaayxtpXLT4JSeYSg4
wacNZ6rtUrmTqw17gNWJmXITkidwUq+Dn6SHWC0LswQkOiOzMxCUvkQ/OGMYiN7b
VDmgJrDGw0VelKvmsNM81ZWu7eG9oCvf5EH5Wx+61NAm3GpzPbzdM3l5aCAGgc5e
P5bo68HotkzmDUAg/yq51zIoRDW8IqQ2f1sTzebLJJ5vw3ncyeWoih4lXgmHjei9
8PJHGtDyyrpmELDYNNtK/ybhEBFU8vnSRnK3pmZHdT2eb5F/vPRcsRp/KrxJlY9x
abPXO03jMs+gB4EUZF/pu+VYBWz4iYfx5CU2KueUNAJknwdUZCsIGmVPt2CE19jI
PHWdAMQ1RYgbZcYSWgJTKFkw3jfMwy4hGlV+JCOlrmeYaZCj2p0G3+U40Rb6nqft
SLZLtyyqzS/zntNu7KXAi4Jw4X78Agv1Ctgv/XS1yD/AS+joldc5hwxWBTLEKNuH
A5v1Ti81DpM6Ye/pZdpYZb8Blr/POMmXqHD4F7KEGOw7dmQzadknVBU9z3iPVJfn
3WgwDl9MIaJJCIBr7B7xVm2Z7jPI6hJ3Dqzw/Lu97PyGt/unKSgr///uEZQjgeiw
Px9kdkLBaTsnW/WpszcyAHKHOBsVPMuN4/poh7LseOPkRcwGsN4Skjci3u5GRcqY
YYJ/LUkIwx8+bMADytfCdxWEM0vBKrDWi8tvNG+05WakOmODSSPvog3g7z6F8+WX
fQDj0tdMgNGK6OyqzloaiZfq2aOk1jFOW/h6DSy9bubRfZEQd85tbJ0JWoY+zhJ3
+1uj9ph9ZiUujZxhqz1inoeBA3mvYP/bA9KrGTQqYio76yrw6TT1d6bZsYLzLxGl
Kd4W+VI5MXNzXzJ/vZi8fJOPFZJVnGjsWbT/LCbiiZ+6mGVn657RT24LSPf2S6rf
ly+o9La/kJ3rxD1xNrfFECvuGvlx3Xi6iY7kYOnGtKuyQKCwDR7KEHSycoSWa/Oa
b3T/ZVhnjmWtDldy2FWspqyu07gKyIKdmelYapMTwpq5Zh5JRbf2reRo97eH5/bh
uL+IIeQ9yRyUa/2ozQxPlinNgBVhMAZsIPTp6E4ZatzwDqTajU5cvwtzCEDiGUtZ
t1WfCAYpmiej5PYuDChciIYnVRZO8V9ruTm8J6zbzebos+slubzdI8SocbYdYnBn
tAhMkwoaXPfnKcJgUGYYE9NLLDYR1jW4cPD2sX/lCQm9OhoHN88hNkyAbTjIpnDB
7uhYTnrPgCLUEM5SSJreirdqMfLNb05Br5F9qi+/uZwVSkG01eOozjw95sXAr8tX
Z8dH63lkwAX+OUgMg29rEDc0P5wQ+fIfeTiwoX/n2GTgztZ30HI9EzAQaiCcH+lw
dxrhL5kdJT8FBLK3NqJjILA9CJwMqM3vPD5+q4TCoUiKpgTgeATMRwhGy44lyJBm
MnAjd6wfijoaG+WdqDmQHHvDuknp82TwE9iFqhd2x8eV4CSOh1BXE5hr0hUVvYld
WYcSg2dM/LO1+o17pmsGODZQiiYmvYEQFHOM+nQdiiXkpBYPCTmol19vS77rLcjj
Eb467tGOrPgm0up8Z0stnfeu0dGQbEi8ydUBHy+SnQiT/5Vp9qKAYiX7poDHUUO6
V8CH6EoLtU47eBmSixz2zNNSAVe+LXppiaqepI0mgtuJVHO+28c6st5A9vO24+c5
+YmqM8tEfLpi3EGpcxU5aDaSj6ZN5c0xQwhkPWAw7eUbm+5z1i65gBy7YyFnrd9b
edFzmXjflS/gv5wSqMPfVy/085ZrAAR1hntG1iud3hz9IDh+NSO7qvA640fNo+3Z
smjLWM+5igK1P/HZyI9DsrmIf48taL6EgQ+SC7YdaAE0e56u7qFZVB4nLTZk/mQX
2Zx/x8rAVpa8TQuW5xFs8m8t/6BngxGcYEWB2QzlRLivyC1+QNTSp5pP5PM2zE9d
yYaf2rk0CMgwLKqkJIwblAwzwu/heYHY7DFmynSFxXoDhZj+eDFOqQXArQlkGZoB
cpEcwG+/Hi28IY5Zn0wzn20ntyGn/TgiVpEAj7jIvPgucqzY+xwAkQoqJcPjnd1M
FyC3qhf/aL5fhhbbG1FLczQM0g6KEnkbFRhLgl+wmHDHqhG09001UrlDJVwFTLoG
uddS9x45bPNjbL7RN6nXpIRQx7DOmK8FY23ytfGr/C1FMmBzsTLlTPkRTzhPpjAo
B32niLNgd7VVnzBLNzAjE2Xt0Qsl/LWXVUVukP/Vee9ThHWHm+htZ/o98IrMVZeg
kD3e7h8Y8UX5V2WrXq/lrPmtb01Gb0Gq4gtvSuevtdM5xnGF6VNohtQFPudjeZJG
5y8BfjYXS0RxpQ443i8Oyo6MFguiAwowBzqlXoXJJxsYbloWc/g7MCha2SOcZuEc
Ss7SJNrB3aD9ETNod3I4tibhXZx1p5JDC+M4B6OAykbsbaCS9dAr/us2aiOMvsRj
WKLN8KBy6iRc6VgjwGchOgUpunWbmM6rsE0+t9S32lsHIJNEkXrQDthmxR2wGkck
v0YHRnsPth8tjEC+gLk4EkaogV7vEqbq3Z45kWtPGZhpHxd17EAuDSUOhNO8aJLt
Zv5DolsuS3OZLaynn3qKw20wfPxNnaP3tmIkgZuJ5KDrs6z3sOKKGTKYsVmx+5RA
Ekwktcwa6C6Tg29sH4dLDCVLKY06i2wlrzglKZNRQ9vjMD4YNckRXksFV9I4xOKE
86FMa1Sf2H3Rw5Krk9Kvy66OiAqahyb3YcDIfBW+4o0Qp4jB9gWnl8aqb6IZ2JPY
OsYdiEsFrbS2nKmxWQixDqOBVoUltLnUZEaBR6y+4k0nsRUEvbm0/oTX5MpKSN4+
JCS04lSzhpM1rW6uf/dPTUZObb1HbTPUfV0JvGuFz9+tjeK/8VC3Ngg8K4n2jMTK
X9JGabnEeNohce8B0Pfxe1XjyjLQAOzTfXqOgQy/qwrjZJ9OAR8MYCfeWQrGOYMi
rhN/U5sO+IerjsT0JAUe/chtPC3rlUQV1vvrRMQLzcfuUAsnSICktxwsYaMMrN7r
BtKzk794EIUSyGuX8hlKvTv7uXrBXG4fb90s5WlcmEKyRLJqek8wSRGK6AlVZQmw
aP07qyPdCNzDVUJGQkZDfYoq9EZXJ8+DnktClFJZyszwwZDzQXT0tngH2c4y2NxB
4koGCQ5xparXqpt60XdCpwNB3ncplTtkB23mv9u29XojKSVccVXaWX42BrBiBBB0
vCOYCvFhCt+JJ2my6K6wLgc42SwXF3DGJdraPe0RgCSN+TKtM40DkKQ7r4t5SQbW
xLXourJSMCyhgkFc2PO01/WK1OB+adAtgi0sfmYcrXUjbrWrBt6pQUPPNZxZDojl
jlM8grCyOxfyL3SmMwmTN3kzCBLnLqena4Zu9gZipsZ7yNRA7BcO3/pSAqUoqqXo
nbL8COyrkshqhCwkZkiJzHVFLLLsT3tdEu1aGS9oYSRjStPnDkFcVOF56XyKu6GS
bsf1BVgSQuL0HhBMKY0yjaDuM5d7RiyXvOOrgMQK1as/jPUy2Os9LUmKOAzAplrg
ExIVBUw66AP63ajBFaBMYwy12HGlrfA6tPncRwQTpkvmptn6FONCyN2OT2OuaSYL
Or6lHLx70SrL7Unj9vcNMeV70pa96ARYm+cncrAGGdlQ0eEWXGXIB0iEaeWyxbEv
2uetScAP/f6ijsqv7WkgmrrGFqUP0Gnl3p5ouKJtmebWCHFwiXFnsvGD/2X9cQ7b
iuOm3mL8B+NeNtWcF7w9E63yW9Rx4Tb1bVYiEMvXOQmZSdA4mU3fdIjD/Fwiw/+q
tvqPAOzz3udYbVrsi01lQ0F1qB9Zi302GMrnQAWR8Aon7vnxopTIg6cr0ZNbdJyA
vJUVHCzV5YHBIrxpGe1vB2t5mHgN5pZDAXhNh/F7by8GgBXbrTIT4t1se/3x/0O5
367DxSrIsQQsVguhX65t4pFfPjXRkaK7QhNNgGXQ+cGdgrufJAlVKag+mnfd81Eo
/rU8tCH94KyQQtILEOBcvg93caFOBBPdgqjwU/LBenjiQn8O3upMpow8YamXwrLc
gmm+uNMqjkLIilnvBlyYrWwbPsZsXimq5sycjYGj3VmNSSSe74te4hUqJ4ti4iUi
Z3iVEbsjiiUjp7fBm2UU2B3E9yGhhSu1mr+dLM/+0bonBxBEGXVEy1l+Acknh377
//v8ypg6TFvsr2s7EtYxnErlHd/2JfrZCPFPUhCmwCPyoLlGaykNwnEDkTamDNfj
v6+RSF+m7lPtQFLrzHM1+VlEOXfCkjAE1d1de/pIEcJICLNukPbCcexH4CCS280L
fq9QIYw8BErS0akxF9CdKPytzPFoN1FaC8rcPswyf2e4XGmtdVlCD8k/S05LWWym
FZx3qG4bb7J+3OfVLpsPx/e1X5e118oKyKRQXaI283b6gY0zoZYuRMEPt/4RJk9D
CtTS/1PIwkcrRWIksBVunXkwVkDljYqBY/CQik2aP0w054ioL79jkxH9o8qa3Rp9
Hno4Kcp2oVZE8D+oqYTNMyp1J/3+xOa0WRHxLp4c/MxbRpeo6jHT1a5M5/FVpg93
r1R3TlPgcz05/giQoGLpyfOO7LH+NNC41EX736cZeILXsWnek4jCwbzRNTKkUdox
t3nm7Vh8r+leU3ie9FachfymaOldv2x4i+st1d/rkN+oTMQGtND8a0gWN0vRJQyy
BIj8+nU1moDDMxDSdT43XeXngW9RfltfU/5Taus+/eWd7NHnkfu1TLe345KuY5dR
E8YTXqM1FR0nEuk6LKdfkrTqbK4cuRpDATpgreHj4hlWXAxWmtL24CdG6GfZUITH
KTs0f2aFuD5oAd4oH9N+N05QhNcYh0hAqKDPk/P+xjjb+2TlS8XvTFsmEBt6ESG0
rAcqLlq6rLbWxQf6wxuKHavmq4y2w1ycNz1NvpUdaSeerYg8O7SrNnEazkb8ZbLR
JXcNDV6VTmmdhJGALN8afBnm7jro6WA6Vmx37yYpAfORdwGaPCwjFaav4bCzp+PS
xxgbLec8r3TT3eXVuNJblSL6d/2k1aE8BQ3bJmsO/wD6C/7A97zyXyKzY95FOkdq
HLgkI8UilyC+Z9b6M2JECaZeWke5LhT0pGc9qCUZRCv9JwWnv6K8L0CZnKOJEoDd
jWfM6mywmTE1R0nL8LxHFAwP3xnLBq2Vxop2XEYKYZezaO+mIHWOgjgI2GFYytxg
2FSAWwIhidE7/hvwmbPdl/XGvPEtq/ej7In7F03n2IDlFCY789jpd3eDn5e8ib34
kPODx1HiK0G8qSXhdPOTy6OM3TDpt4aRel16lAo2yI/CaQlX36Qwx5pdq64JLOHw
m4hxnehe1jaeyvxkwj7+0zb0yuLjaVXJ2ploHNfdGgcbnTdzgRwtBPa9J0rFDkU+
M/h//TdnjwN46edSWMAubwPGbBWq6KhNdEtwrMQAcgX4SATYiy9Ibm3L8D//ce23
nUbv6Uc1npqQ/k+v/crSaTSVaqjLXZKBUVQwCc1kJXQ2sD61pR3t8Pog59XOfBuy
s2XTCiAxwEEBymQ8RDvnaMRn6u0eZe4afbMWGYquXzLC91feD042ojMbgKh1AGxj
CvMW2Xirt1+5ABpwuetein2mut19uGGPz34X20WlziPTJcN3T+TkFAMFv0xRWI4J
8OvBzJGGhly8dDxZL/v+QH5hDJcQvVHm6mHfyBq6BXxcaxgOQO/XrRWv2ppOfBfu
lygCYBz8XvGv2uI9SWomKYwxg8+L+HO6ZJbNXDXC3U8ybT7IuQh5fAJ12j1AFN4j
IimtV6x73GPITVYzc0Eo8CdOgcfbVq6643H3DwYfc+1EDB1w+NmG0LsyLcu8hYCZ
JgYj9h7t5YQgTl9oixpyRAbUFUpJioePMWpXJMoPRs1NRy63n3JmKXm4UfBcD9Pp
Bx/BIRV5RQAg7qxMPGn9jOCRuPiEHNeH5NKkNscf0q9tx9/VP7MFXY6RbiIEtS+F
ZvqWRPi9F6X3LNVppGCsI2Pd1gIt/psHmgxQJ7x7BmXuaowc+w3aPY7St9bCvt4s
KId4d8uJuUVnATaE77UZTpgm4sdAePqSDSArCk300bEABJq3lfEMmYE20ifAAZ2u
0KRXxAOvt2Ts1ROjrtXTf0u3wDOlD9bTyUia2mi638mt/Sct3CNILFEqYzFfY4O+
QgUriO4Z5phK48f+lJYDEOJcv6bBoFr1AzdirVCl+Zb1Q7jI95rNmz5Kvkv9OjEb
cDTTgO7qUFOYn/MMjvmHtO6Yhg7xAZfG2AfmMQYcKSehHzgzpNmzqNzYC0jsBTxq
bHbW4Bf19D5yEtD9alnnhO8Yn6h9BT33MrDAjY0468J9MG7K+23nAVG69UXTjs9V
BQ/dOffI7bkyTo88pX3Pmvi9KC9REXy+6ksjW6vlSaRFqUjb1ZoMrEAagu/q63GL
lUebCzh1rz51SJekmalkWW6fe6ZmaXMmeLLrM3nfHJq0CtoxoqW8Irh18+/jh4Y7
N0mVk0CMzKMAMOi4/Ew9iHcMUGc5UQNUrLkCMcfCfEg8XcNCpxbC/A32WZJJK3Jt
nRaOzblXZk2gCHXmOGfr+/unGP32zve3s3kDM7aCpSzPmiVLqs/NVT1cRMjz2v20
vftQcsW4NpsNnn0IcqlGT7zGbnM84uEuqlxRvokZVfyFYT+HmCsmdlIaXix6kEst
8/gKT5NYnAwHgaT+fD2GScRIvgd/klmQ3246Pihmh8F9Mg1gQOFxSuiU3soSmNPE
HyKPls2wogBs8KoM3+8z8dnfWd2eKiOful0HiBYccsp7GnFi1FJpv+uKLSlZQNye
tB/FnR/i/MKh5bhl7HJwQ2UjJ+3h7O+prtMv2cN6Rgt0ySqkaAvXs2LD4n1oW1to
qkHt0J9Yvs4lvZ9XuoroJMSpUWmB6jpgPNaPQcskm78q70M5CHfj9bbrgUz8wxvM
QYWNttS5DvQvrXQ0Tcoloe987i8/LTAQEtV5FxBN9C7VvOtlzjTKTgRAEigcbnYY
eU4EZfnq8MZc6V3Zl2xmCk7epV6m+pZ3cUkLjOXppLyQi8ML9iPYOZG4sKowEbvB
CrYWslr8XrYKCN3Q5LTDrgQbXVT4bAcGIcGKxv+vvOis4vinhO0n/bQ1IZcun7FI
81qt2Dl8qJydAsQ528YJGryHyaLmd/JWxNiFaZcYwAdlkfwt7TT6QgZB+ZyHeajE
uhKpa7WPUw8Y+NKbSQZWGZEf1xNS5Aqlkz2N5drfTAYr7y9uwMxx86DC9/7WIx6e
RIK55Dk02yLGELxw/Pf9nBaRBlNtDKX2BZFEFdqcYreupnzornrhTQUGRcZEs7eC
QV5x+z24n5UP3qK5Gbqj0uVSf2AFVkPSPQvyPAYznsn6uBwJIkmOjGsp0OJH1428
5gALwkO/iiKhNNgCX15J/xwV6HtMJ9Vos7Z/yiBPcriUIe0d5eMh5CI0Zest9OA6
glgiRGe37ZPmzevS1gH9oJ+eUe4O5Qa2S9QbSZ0QJXyXkAl8ZFy/gtxyOWuMSCnN
sAAuOnN81KcCY4riBQoEYutXGjr2LxZaSR7Y/a6V51g8gbT3tQni71YdGah9WY5Y
0A+gDErQUuEust1pOkxsSpQDc3cZe1Q40GDw/LA17G7lwkQc0hg4W8bmR+z8uK7W
zn85oeUMrYJE7/plTKBV3NkG0o6a6hhubVdpzoaXoEZiShXTnWjKoBAKXQRBKdP3
JtZH66/K4eNbVdeH1FseLWx31f1funKXTKhJ0uWpaeG3CcwTGfQydfBvsOjn5RuM
MkxhsTrPcuAo2gDdigjBl6k+Lcm9rEc4Gc/+hPgxNibDE6NtEX7XBAbwVj3StFfw
O9F7w9eMyzrd53OejXNOWtdMJ9tnrK1Fe/nmMlZUoELqISt2SU/h24Wkk0b/M4dR
u+BzKMKSgimgHV/xSSqt/535wA7AiFkglEeff9XILNMJaTJMwGQ2gnOray5PrTQB
Vcxj2lRSOzu76LpOWg+sVKX0qQJ34TnJ96YmzHj/15k1F9/u7yiW8pQcjInDMJot
1fEqutcJkeUmrggK/Jay/8NBMY64D1QF4GwbdvDO7vS7uLxc8UeCiij7ZQIaJxf8
bH+OrI1bU6n+Zh8M1bdSTS+F9SxP3M7js5AQd67J5ssyx2jrqa8fekab0R4w3u4L
3+DHtobUe2mCdVq4JC85oJtioyhdAYO3fFDE285UU7yBXGi4C4Gvye/v6dbulHkg
1MNUdRw2/5LDpV1s7TxPxmktce01afateaC8vl8immXN5CTxa2s325A1TEOCYBeA
h9xmup3vs+KRcSwsBY+Z0L2FGWSmrEqgSYkrCXXTvLFOnPyL6KTtBu2gI3hrVdcw
CmPwssWoA8UHqLq6AIJpe4FTa078BgKMKdq7lpthFGbGjccxtsjYuqQ8XzraYIDG
nsJ+GUIW9+D5ekDu6Dw4hJaGrPhlCGyFX4t06lgj5qHFlXFqOhc9gNVzeZcYCqZI
0Dmja0u/hnUURq+c90apPUyB68v+QjQ/Gyvf7kf/B1bwQvl5x6Pi95GutFiw8ARh
F7vkSO/wJ85i/bayZ1hKAXVBDUmYT/BH1Ezi42Ndg0hihXbZSp25qhRjaWK7XMy+
mar5aCwpkgUSpxy814wpUJGD9aIWhsoVAom/r0LdGM3YPl4yrEuWmSpY8cYM/XKr
OiMN/dpzzVdTgN0a3i3bo+G36++P2VMlXRwLsm+FbC1+fKyUexRMUs7y21vNm+bu
TfE3GhEOAP8N0VMcddMgvIHRmbhpw1wnURbMtUF9Wi/1o+nkGTtC3awmDkdTmwNn
Ux92S1e5AjplNQDaYcC2YrPCmiGMGzLXjp6CiudTq9eti40DgsL5J6CaIRiUWfu1
qTKkHJkNIVopLp9BpABJNqYeGPpm6Ds8f4lfUmsQSogxOvE7z+DrrpHXLTDsrJ+Z
3NEN7HZWQqj7n2BDobpZu89A8nQ0/I5005DJOL1XHESJibmgDLh9QRey9/SXkb7A
DOnlUJi3pRESr8MTQNKaDlsxhRKN03zehoKwWw+i8zhaJdnLODXfAY8hqOBMm4vO
ZDy7cXh6Qhzubq4CQ/O0KtxmBiYdWLwgbERM+Y2Z1c7dMdpbcfYjyGv1iaDunGGt
RjYX79lVyLMsFq9sW/JHg+AzEbjYn0Hbel4sOP11HrZMGWrW34SNL05RziQKXv/J
VKKjq2nYAe+fEtbyuD7O050vP/lXb6EY+Cd/NOHs6kUN2cL7xa4KVrb+4Vs/ZAgG
cUNcG43djkicuNEsHzAg6TVSVpgVF7An3EtyNbwno706CYEFCS6ta/M9STuV2k5D
nNRo2XvjrAKpmMuGosK7K46xrACP+QkteXsfx5UzrpnbgsiMxf3HVxFUWJMz9Cvm
bNiz3YcUDsRLGddGd2yE5TkXHZh2AGtGhI55KF0gyOoD2odJIEnBtpqsZ6GQxu5y
h1iscKlWZFagUh6rdeKv8YIB+WHtJMmVtCstm+ibhJCA2pHD2CpImqeW3u8T9Dje
VO7HpSh8oCEGGIDxhhtRZGzBhQmI1VrbCkpaBiuL1gm9GDAUmhZ3TN7NUy1uQU7M
iUjUHzTbeJF0V/89G/QrO0X44lbvWRVcS/Sz0+/9W8OtYYduMrMMCANf8uw6ZaCU
qPlb55VBrHc1DnMURk6gb4t4VrzQt8fwn5XtpthCFUdyJ27OoagcNdjckIqsbtEw
mg1ZcATj3EXoHyyZk4Bv5s2Va0S2azvbqKw6wWshLpJnmfxtVxJcc9ryQ1EJq6BC
GG0wzkFNrh+6oPrSaJ7WQpswYQQbBRD+KyZ6HA6ISmkzOg51PsfTHYn3M8RW7JuM
Uwt6frIquJDi+VnwlXfgeuPT7k+QVYzFwQ7FkT2NWDZHe0NqCdZy8wudDtTzTP/Q
3oJB5fC6cMJd9vazjdQ+VzeiiUJ1JaLbde/iNogEh9XmLPxHt5+7kjWecjmKn7iB
qAkZuUQoxomo1xmcAO6gFebcSeb3JdvKUd9TtX4RHlHI6MialSwelc7j0Xh8OdtY
HLUeRRNelFS727p1b7i8A6s6rA8kTQG16MRdiXB5g1ZSaG2cIE90cUNy/whQ8iOi
JwlXmksLr1uMwDKI7XHD4d30tUzqcVtSOmWmVuFT4Jr1eb4kuV+WlPM9PIt6CGKy
ju7QZTbDl+mXA5xcKKeVRwNrbSEcBDvQRdPrqSe9tPRfQCTCoHlrOm+oclO36bTD
KqGdfhTgLvFCjyz9gg2n9UBc4XbhSWTKVuFdifPl237NuFchiEYrp77AqLHZDxL7
VOOFW5oKLKGhGEW7i5GVq1AFIoBat2/iALEZi/v0OPzDyFZWbP3KFUjC9AxThhVa
VqmozhhwJfBnBQqJnQVN8B0q9Az0snbh1P177NhZ0V87DEPRNgauXKsqD6g2CbtR
vwMPJ2cS8XvKs1/jHThVvpob+Gf5hepg8FnNoogNfFPpn8Ve5pYdde9vDK8zzG7H
gxMWI98zqWENsQbaoL0DwtqoUPYfbjM0WALjEHEWw3ywH1CVuNqhCGlC005NODvB
iG/fGxtOYu23E8BGgnvNo66m97Fu2CCKur99iYeA+aQ74EHwqlIc/P/weyUDysDB
6Bz3rJf+FotQS9IoQoCgNPT+bV5KCs5jlMMwwtHlzFwj7FRs/SFLScpgW9/mlZhD
8dMqKRcZVRFGUHORc1SkL/DY9dCWsEHlYfFlMxOSF7Rc09mg46EAw/4LW2Tz5ZEO
wyOyITXxX6i40zHquRXXTqdsg4zkVFAvZ/hOZ767nb2Xlt+lOuwVe5b6NWXOS6fe
tWOJDUoDYBTROEJKVwcsgLpHobPr+2u5ceYSoxUYRPUpa7IfrI7d+mUZPDjyP5e9
d0I1+sEY/sxwSlBYddqISy07SHYAFpzhATRCLqc/R2+N0QxOes8mzuQGGUpFgaGt
kpSu/px6FOS/sBIxE8/9d25O7BHgOYnK2UwmtjgIdb+7Od3aNYS7LZRXO36HnqLX
gX0uHE3Pu3ioj2nfgP0aqn/etvXZmnTiNiSNlBrnRnt6loOvDnnKPCWSem5RosPh
+ZsGum7tjvWEgZQCU2RcodmS7EaGeTne4QAfYc+NlM8ojkKsJwmS3gV39aWNgbaL
c9OCMh9i5FLX9Fsf7K6MgWufiMCWHYpgDBvi7AnPAxHzryZxFDAee1z4wX4kiZQP
pNw5CnyhprfCfO8SKOGkJpc7mBXvSU8cbyBA73GpitWigr96ci9zUtTPJ9igRTvh
N/B3rEnzuIjHvgUgkq4zsTr4oHipVoUmiYyhJZmg9tH8NRRkWNVkacC6d6Ajn9Ro
L1ekVP4RNvAfssqTMjby7xgfwQnbEJcNOgqlRJwhjB4TrtOTzkMIUbnRht0MHENG
evOz3jfw4gXdD799AQF/qLe+SfK2DrdhXyb2btrQH4b1w/CrqpKMklFDHWsr0SJZ
4mRDMoQWU39b9lqtvfW4EfuH0Jwn4UdvEtcSvWY26J5V2qHYIp5q3kPS26MkJwDr
98z2JRjqKeFp4dApI5RNNnEn7vuOzUxL6qfv9MLptB8e6DPzEeV9Ie/zixIXcD5h
dv8VaxSWwVmW/eBe29n8wU57gNGfXFHyHNToSFucBWkYq+9Sf3ocdyUg0vZPV6vM
Q4qUfySIZhl/UoxxvdZuzC78Iis4g/tYmCLqg40sfpJP6+zlHrZEzpkQzcnZOI1/
rCvjSQSDnspIgDUeFQaYn0x5OUl2IrQZ9PSvn98rppl+PbhkXiQmQHB56qtwPI0w
WRxZuGWihVl3t/7Sv4nmhxu//AGOylbvqrXfJrBmHNjrgRGql/tDZisbzlTEBhmv
Vy3Coh9ICq4QklhUOcyIsgWFk10UIwKuK/pM325BfwLOnuYptBfWgaEr4nWNZybQ
kNoPgXpVpf1A9s7UYG65NMAXeEl1/NBLOk+cctpqYzkPDdyEPrdQr5zYfts7dGxc
MZ/R3/eviN3WPpNhU9/R0yAPPayseVBThGWe/CLwi8thnypoznxkEjEWMOiLRVQt
XiCQeyftvBMlWYhf4ViDbOQrdqXc9mUsepDzKX+l1YE3k7Fl3AtoDK+h/dCGeVU7
jcfjlqJQnwpJrxwzT8NXKMJEAjdAe9IqAR6NHfq8DsSnml/BHM00gDM7jRmFlR1V
UYgL4SOSD/PnBtXso7UNcZMe3Q2d9x3EuTrtT0kqW16hU3fXafOeYxsct0AN2u+V
qt4VBGkY2TWEgyq+7odjoJoHZrlBwdFKczDEdp6RJCQdp2mmr/gTfK1Mwj18eXW0
BcuxOYn+hMneWDGKVZf5t2lWIz0CRqXv0AYnfdOF55IYcPqMD3jqh8t7NKSgy6MB
o3hlDX+uH7uCD8KxgBMMnnjT9tWApVabGw/cqOub9rapkEmHAS4JGjGrCynEQp0s
cwNaaoA7TozpQQ+2ebDPqJyB+J7B7NskhKhwndBkoNYDk6/bKYTOxS36rBKTITkj
3KhvZqpODo6shPsGCh7xWGJejZ7Q1lcTYsMte9D38FGOG2G34PQXGC8h/X1xavO3
TqLiihw8FHDXqu0HXX5eII69x7gJs4SQ9L+xSWPQiX7svpZuCeXs9OzZRX5Pcus9
5qorwULjznQAiIkFpZR/LnndoKprskZA5tc5iLTm2dxTrqgqjzRgpuGN5qtrhgvW
GhzIGSr7FSP98DkQas1buJ+So5QQHwLZpgeIgp5abfVTcszD2jxd+PrJ+cAu/xt3
FV56YLwTjgXUA8Amd67x/UIFKmu/lz9A/e+Gno5hS9/k76oYy3kc3c6L18xCWtf7
I6eisMS+eKe1aZQFOgcYzCreNaYOz4borgwujqjRbSDYMrlplnCJ558ijRuB+J8b
CoMgEN6RD8n/7EoDJRQQOngEQE3us5atWzEtARPIQh5StTy0GhRE729AyH9yRo7z
Sk+QIu9c3sPuw1JDuV3fU+E1kpThKlyOwR645n+sB1CUpofzuILxNq9nGy9Mgh7v
QNoi6RTZrLhdl0w5gJXcq8nh1dMRJZZskXydRyShdN5rXecyGfZxS/lQI7+QBt1H
G3W7L2lE7w06GaUlXFqmDrrz9gKDCuN0TMz1/jP+iYZCjDS//JdrlHlO+Wa/SisN
OlKCglKGvWLhz0rUk74TEVNKsNa/OpE7dOEW7g8v1tuFpRs42vFdIepLPVwcuiCN
wsU8l1pua0x3LOUz7tlNFWx0HujBSSgHr4YOy4vlNJoRXVXr4Y9L3tYacFbuHoaS
gWz9E9Mz4FtJNppqfC6JzHUOtWTuQde4i8bNx1HScnK6HF+ejvjWFLnWieBKrS6h
cx9jXfg+WiP6ZE1B5cOQ7ol/c8JPygBaE07I3UMSSqfLc6dOobrluwqpRf1z1cnp
yDQSU9RqDh+ds+3CAekNb+br8wYX1LC5vmJn1jBljrOPeu2hZxPupxxTg643CnVG
2v1tu4UMv8nrR08BRQqprG09gT1QHfhFL8+w4O9xnNXC/gC9/aU2nh/yoIRPpqZw
E2blSsnlpk/bwS3nUx5zyTiwkfSBIKVUTifc2lRZvhrwakgp6vaBffYUycjxKq6N
UGbUzyDqX11JM6/XIrym41kq/klVUAsqPa+qGHBGZiamI24Edz4LOz1N0iNWjMLx
OND9NK2LNliCqXqQmWpAlbO8Uvkojk+QUGWgik2YmzrFEAvbpFPOPk5GwfSdftkK
ELK4VxEXGhF6rDTULZvb2EQ6bORc6Bbc2Aded1dNuBuS9qS8NBt0a5vnYSotx08A
bwxj1USglZbRLviN4HG/BrLlpfMbjUrIFtx0kVMmztwOBnOyNg5EPnkoSsKgMxhe
aAbkrhkUZJUeYvq6zqmGEzxusTNE6oj4fzvRy1BQWZ0j7cVXnXhWWdPox9KFVpES
Qov9PfNJCiCYIWFGFIQ5Y0JZi9WF4AY2Nqmqyv6W8CFVj9A1MGXIecBS8sidCAtJ
sJaZaDHI0xJaRPQB86iQbG+4/aXWaX+zFETML36JRKiphxu/fMAW6gXT7/tg2NuI
3xYMxmfuzd+CpJKszXYMynu+2m58B7zzv0yXrqmzT6xJvZ2awp32Csui3ccIEaMs
+2OxQznsIaaNe0Kby1NzBQvttMLIR+BSdBtHSqwQNUaSIvki8KwZBHlvzmL/lxJj
CHkb4ftwr6q3DnM6IoaXyd5JhBMtCfAQpYApM8a7nzr8ScrdUsXHfKoBOaIDFOhI
8PDftYAlDyvsLch/URH/X+FuLMZYGJODuJfsui/UfrcMGvu6MNPJnTO/UahVct47
303taYIp+4lwgZXyhlas8aRxTwZlbvVc36v7RyXsFezxtQyE7DINSXWYvrEQYsO4
fB52721Fm1bOuZZrmcow7XJfL5vzHvp7zhFA/pNqkSTIfLQtyX1ktS9Tnq8BwAXB
Ll2SfZJCNq6TNTRI8EI8FE8biBqdvw4+cGmLjZ2Zhzg0c5fTnb4e5b2Kru5j+3o9
n+cZmj3EmvfB+6d2KRokhDIRP89BWVFtiV20VvTZHBeiH+CDiQdFTvdB5LeD23Tl
SkQe7knaOJxh7UPG7qUxUh7XKuIlTDipO+hK4HBI5Gk6gyryTB4mgnfzu3zbXaRk
1jBB8zOdm9kCvToO6XDyajFEAzURfptozjmOnlZ6DzJchkwOlXJHIB0DP96pTNfF
u+lhLJoQG4PXh4gHSFB2GwXGNOrMbdA9EQl3clGjT3YkteiGZ9m3GMtsGkisLfBU
owPba70JhbkyD0hpFP/LfA7qUWh/BhCMlSpNPJ9BsS8/wOSK4hdC8uX/+hCL1JMQ
QCMfxYA+cRprLFCeMtyUN41rzcwsZwRJ+9uCUdDvMOnt7/9l8Eavw9+BcIc9Raf5
nvzDth5zQPpIPA+zp4WjS1GBfXzjeTYLCjGulMZleIOBLqgmdSUpi9Fy4DV0Ts+Q
n6oeP/q1AaivFOLURiYgwsF+qsGqMD7oJJnsScjxN4kgnKyb89psgBxuT7J/vXd+
yo7fJW7aRolCDYJfqgt7IuLZyA7kWI94Rtu9WI3hYUXM/yiG4njGqSwKKIi2wA3w
dubYHuZUEGXQeGza9G6O85RNAZe3zFDUhGaMA55+7l/0VaZoqqlzUJOnpydWA+i1
ot6jjI0hwBPrMfrUJD0oEfCtzIdrP+QJiu+dmZNfAL9bycNBl47YYJipPMnZ+YWh
OloeJwhiL3Vyr1QJYhlO2urZki0dkWYbV3pZWG4Ac9xotHj2kSt693iOfMQYSrxK
7LhGrUuC7/gQ57I+9T1etzuDbXlt2vxrY1FeEDTUz6otMBMCWvFtTtvShrynyuDg
HEEXQPfS8A/Uj+vcEOid1cAk/Ek+3OBdxiibEVWWXWs1X36C8dYl8n6+5OfP6l1X
KttnhoEYb32+I/AHAsexqXLvuLNBZBn4XkRWV31npd1T2gjtgsU3F6vuNxCw0Dou
2I3ao3eMyhzlA78WFhu2C2lmMyEWGekJrZ1MB/xVbE1kQNl1DOk5BYHkq927LJ1g
/J/3ufodJJZvzGpCTGZyWKUWpNrIH6lyy7Rfvdt+r7cTIdcYbWzjP8UhTiq72KVU
OCZNpeT9InyPQS+e28os9iEecKL4LXUikoQF1mF8+XPa3xA9O8JXRZCTyERpIFAk
qyLTdec7YhBG+3qCOwFNWWEvI/9FrLTBN+x51QjUdEj5in7Q/H/sdijPF5mP18Jv
RcH4ecPxeBtdCGMucdWW/2iVR5Qe10VCqsrB+iPMnM4mdQwRStkkPU4c8gcL2c/D
d2dk6CFNEE4AFxaRRoD7CarYf3x5SX3sKtzbQdH5yR+kWr0LYBToz+Sb3WjApzfe
m9JgsRbfeGigtx3vDVcPmrcmCKdE6uTro2MkADi5Fuq1aVIMhDrxYkdN1pTG8FaX
33ed6PG38twLAKH4RKiWMU71KmKYtmxDpFnnc0VZ6E5xazcj2M0OrBcy9ccYKhz/
c7CtbfCAsETtQReet+N5SLeX9++PmX2oto24LN/RXX+oXmlxVzxrhnsI/dck6p/Y
lX+mp3EKIgrmM/VqWRBix792hao6Uyi2pYIUJMFMqOOMeekYcl7qqSsjcJpWSK2B
+gHhuEJPBJT08OUwf9b3RtumkXpyYLPEEocZigv0PIf9kYPHWdB/aAmNbget5a1g
t+QW2R10sGNucVzc/zCe3SM/+m2aWeW7F+TQ+pM3sKJw0JJK15mJtA3FzHZufXR6
i8jrmf79Sp5SbIXAXfAYJlM1q/Dg9pHYLmLmUJ8dXLSWuWZNk549SFkp0Ep7+wqc
blFw8sO+LdPXK+EBJiah2DKr6ba1DwXdodZAhF5chUjpAAA4fV2FcO2H3nhPrJ0c
hojzeJkmiuymOBhEDkV7mM7/ThgR+K7LSq1Nvt4iCNDDQJxVUYfwUjEIGPoji59B
8XLItkATLSieZY75Y4AKJ91jgNYStHRtqKky4F6PCympwexfq5a6OwcZmiNHIvWX
qN3hCfM4tKHVkvQrrYXTaNUm0OSdoVgObABKdKqZkSXNHIwA64Zj3tQuD0EuzbHr
2lCq2KfwOrpCHkYJnnfO7oihr1Tr0QL8M38WqaTcouWBBENsxFpgQvDilBbn3CCC
lvD+Gq/WS/PDIn3suJzUmR7lP/mW8GoBoLUyErQ0qzkz9P3VeCjtOy1sbChvfppY
kCLfrHR1QB4oIYfRU0X87AM0j3MFRCiqx4uDC1gDXZ9dRjc5JRzqO6WuwYk6iOsk
eF9feKQRL1igpZiymv/uCzp4vobtvFgsC57Z7P25nZnhGJR5lasQGINKAPyj+m+9
8syZ3E2G/x6QKg3ahhAEtEtJzCwPOwop8JmKv0nOkPkbtFma4+sa4+CH0HQcYXlR
RkSoC7cgsrpLiyb9+U06FHh05Ggwi+TJYYq3MrVnZQwi1M2nNN3tglo2xj5IixuP
oy5VtzahV+r4N6ZQVYCJKV4YwCQzLZ8EO/jzhFxUpKvgaDvqxNfDnJRrNTgwPYyo
yy+kk5vhh/yQIDGBFfE3Ghsoqsk23HVLeeVfv1pdouhV/hQu5hznd8q/eYLXiBWW
Q4sc+CX1+oD6FG6O+Ed7krLMYoM1hBfW/MOxr+CLD87h4IDuMb4NaPBXk+erET0E
vD3IBmBqMBMzlXaZwCtp+PSNPQRCcPdGsuKcHg+b4YqPf3y1UoywVXr6Xgml5kwh
VdrF7uAIfPg4iEEVQHm1lxLtsatP1Y2naKdhBMOrVzAwKlzX0GcQvhMhAO/wsbfJ
i8YFKiiwkOth2816NcsGurUH+YUom6A5MqPQbydd98KLjYViVNfwKSlzRwCS29IU
h9Bv2jgX8lPe/8e/qgXYZUw3db+zbDP5jGrFptZPzKgbFB2VRf5YgbvGui5ztv5w
aniwEdYT8VIVkFzVO0VpHnnw/QH2RwABQjYCSrax8dks4J98QtAkH/6LDZHQgpGg
pYwr3HXch5rb69ilN0OdLh8V7voNqUCmLcXqLam85l5ogl6FCdDWUYxXj/Mmb4+L
safgD7GGl5Pl0xNcCFUu2klS8SGpwpGrXRQ5yUCTmqR0DYrKeuh4MlpG+XeIu7YI
PNxslEuuebqCQUpVs20w3FIrMRzjxZrsYSxgDr8uYJYqtvoDLX7ue9krobvEmK8E
DJ2i5X5IP2p/0toAQuSaLB/iCAT3kZFeu9qAmfsG4AbVXlHHWLtZZqNvtFU9Ex6t
NVeZT5e6gDbA6F5tI+cgP5UQcrc5BelWVYOogwii8QJLDjubvZcEewVnHCFRGDIq
zzAYW0mKRL3hHiXEsBN/2ZYE0jBq4OypqCNsb94J5i2boJ2IomIglj+6DZHV7YTZ
H/6RdOZhgd+PULzBRLTTO6VXRlGWt7TUQJzPjmg5UpyObdmehM7qTe1+E+E/OG+h
XK3JtUBgLVhSXPXzDou5V6oQLufIaRdLKDmPZjxIZke7GOCngvYCtznhIy8P/KAG
Fea8U7IOQXymF01xdF3KccmPfwH1TWpUMiUYJvysHn7NKiOapns1iJzCcR22tD2+
bjEJg9RpD3QYTfTocj75qMOTXDdxQd7WQ7L82xEtd/nH/PcnnN9whZeEJ6dXnCnQ
zK1ucYrSUBPR/HxRzhM9RwfiXxeYjAy57v+WGLUkkngbwIMcWf/38PMEG3cTUjoM
pF/RxpZiDoN51ZvGnzAem96roVIFYyoaajZnZh8oXTcb7GsONB17ZCUDdZLcfP6K
4Zu4WpYBNDBI3JUe15w5Oy4rdUA6errtPxz7inL9TOQKM7CVSrhVuv9L8X843EZ2
7h4mjwEs5wzwAEX8G8onf1SOBLXcNpTYnAT7Jj22mSb2uPjUraZMqORDC3E0q6kd
Hp63M0rbpH6dFXIcm8+obXmHZ3+8VOSzfY7SEj/ThoqvlTY2rP+tGwB+a6ZBEVyL
qEJRTNKf6WUjodqjycQILsuJ8xYWDg6887ya0JoYJ716RlPedTBrHlJ9dC4WEScQ
s4hO7EyX+scYwR25tSD2qECzdk8PtA793kEPR6sFflyAoUd2+WpCK2a8u3/3HyW3
/wAwHXyq2td7j54M5ieCJ5eqsk/e6P9eD37446MFmERHk5J49UGE22nYJDqJM/Z1
RC637KeVfuJ/HKeExpIJpPJUqSWb74q38eg3bbk0dRwyH5GOVYkWjtE5uyZSL/1Y
OYmAGZY+t0Vj7tOGigwXkp3UqEC4ZXgIPCJZdhs7he7H3HV6tHnMXGfON4uBhzXA
uzDkW2pe49MQd3SrJyS7+yuEb15s71Q971/zo/JKJhtniAdi13VXwvFBU/ExlhKi
6HrUGXAVxLJMgQ7ig6/hunqJVuG2SuPjCcAwU0BPX7K0DCgokFJfc8aYdGEw/Rx1
PfrNMv9dQvUzNOq1w9j+Q/TX5+LjpX/nBQyPhwWYgv/4cj47h0yRZcCP6WACLIP6
kiX5AFgkcjgprCyuYEIHNd2HTYPEyFEDO4LyyvCtsoYtee10px9HeLtuYHFlg82g
3mWDBl8Bb9QW3gFO/MddiUOsTryZWDWI8JOrwkIQeobEBEyNAiCHyVod2x7YvF67
EueOihOdgONu6cwmDM+PEhjVsK/2kCrCE+NUiESUFNo4YaYPicOpUZc/6tqvW+Qk
fC6mSLxbMWnDteif4L3Y/jiD+lFHtNrfD83Xy4TYPS3rRcxyVK3jMmtEyvKyoFSe
Y0ipsEX1EypIQg/LB0B1e0sTYP8B4zAM+3D/8bw80Dg9QexY0hfqACEJe0JaAxeg
Io73lRI6/TpL8rOcmGdr0+zfQofSTP22l+/FZr+Ga0BOlXs5znQ+hr0M1aXBuZVT
V4tnFFyEvQExz2v6IQRVyywCP6erVKUlv5rhLkHUorwnNldzFZSubNtTif+5TdUS
CCKy42SKE4W2XmlmqxDFE6xa7rRDaYm1MKsK1BLaev8ReCfvjTjRZ/h0q8ogC6/a
xBroT53zsQUy9eX8zxwgKf+9Lx8GcQTZJdw013GzHSHyhWQUoOm5wsE8UYx/xjQt
QHQQBGrImpXtXnZbADrAL8vRgxxCVuDSDXqqjUZLJWQHhrdHHs4bVG5vM+6Bys4W
fkSWFkTb6YinkeUCTrmPbLfkIIR5ivXJnDpNSppawDqpMbagNwrmtcQpmDmk2UdE
OOxb6I0dYWFnrSKGvSpl1SetLBuCmggKPM7CJM2NLB3GyPqfjk64xU2G1kb39qLK
iud0yqBzudhyWxbgFpVCVUK3cKa2ri8NFnk/3lwgiONop39NFfEPGF+QqVeHIKGg
jM2m0xPGkB+iwoKPKsR5G8pGQZC6hSV/S6pbJ79zKLN36BQxUPP8738si3L6nbfF
9xbcxYm72IB58PeqlL/vq8PXhRtfoNH5VFEUogEEu5gTpThYZkSSnpLO3d+GlX4r
Tk15jZxntDB0T20wjKd1OxAXbY8FmpGCd9+Q91Z8RpKn/4ydVmnueBCWkF3ZRK9+
0VVjRYnOqpEjbTk6RvUZ3Y+id1we7B7p2bYlJYPuDbVw5aExtKXg8ZVbJqQ6Ubly
i2vQDijU/alaK4wM3MKqMIwSruyp+Ee8su76t7I7ZUY+iSqEMXHR2GU9ktEe0ZzI
HKnrjr7Q6OI/5GEZty5Pl4lI+nj8otVBPIbaeUAPvDDscMDWeQ1Qz+3VhjYjlc5e
4oBM22mWv+YZAhQUg1S9MZCsOeEC9oExnPWPnohs0j+eLAhXKR82qQslCwx2CG10
M2uYV+wpWqvg9nisb1/LD11SdZftHl6VFZlDXIxyyIxJrrNejSkPB4AbTIY1ZHzt
ohMMzBcIkrLscuoOgKQgLlmIBqEgPJRNphulDYGA7NAg1XcNtmI7ruRse+T/p0Cv
0GE+mW8f51+zDIHK4Ogbt8vYc58CYyidXoGb2SBpf6H9knaWltjnUApsw6Gptt7v
f+KVUfigFviGnZpLE/EK0JW69vovHKzrQXw/hY68OXNBZuj2uD9g0F6D9gSeKc/d
HamD5GFfrZyUiGaKjB43vidUbVm8guFT4K6/8AyVriJso/d16AujyxUjNqJRGoRc
eBFkZap2yN3ykqD0D6nccrPhjbmW48oDTCXtBgRS3dHXJaNsn2Zb9KRtqr+hhhGJ
YEkcu/jfmO6l+aQ8r57dWaIZa6fHMwzvjleZJKNWEEkz2o67lXhmCVe+P6vrGW0+
Q0NkVYSMn4syJ8Q1giJKEWzQhkzr/uz285RRrg/iFQUgyEoJxQbuotpWgNPl84+l
BjQrjObQjEW0A0ci+N5IoV4Q26YfsjULODkKtqeG9/pIchHRKLTw3HmJYjKP/z8A
N/W9WSO/cgRYqsWsorM5g00EhfkbOWnkYn1b7qDJhLHHauvrjLE+UnZ3zHAulqhc
L7ApybENb3jpSfQqUuaChvbBdUGz+uHilh5Rz0RjrMrPJnM1G5/Tm1+YNuxG5zl9
qqeOz4/jX+5piUlCYW3JD03v6K4lLmvIT2nwra2W9fY+91tiMMim2QCyB2tE1LSM
owb6pGppAHYLoaKuGKh3o8D5edso9thUYHU+dSjEQT9pY7aH9ij5QSBE9gU+gXwB
EY19vJa74WbzCzltKR9gsQOmRDmJl8W9CBfm/DQz7SR5u0wbWgwwcqSxv59ve/DL
UZ/bQqwFuFmTcuOFTLxnCEgQ9tA7qWm+uYfTApoISI3HjF/Loa8euTxz93PpQf9S
l8mLEtx6rOC/GUMmyvfcbut6WndG+toER+HHUndJqRG3+UNPghfaX+vDD2e5kHQw
psgUpKZExsaKjJ5Ep6MIuWBLLcqEbuhBQzixdFcH3hMuOwz3CN29h4orq9siW35G
MNXyt8thOSmO+BaH8ydLITiIuHX8IE29hE87TcQJbyzD+ulpRch9g1/p/IS565IO
U1J0Bde8rgmNXQaiW0BWSUdKyZoUv/zi1JXmtJJfdfttEwJHb2suyV5+a6nmKKXK
H3TZiX6mtzj1RD2NozARIo0wC5L/s5LwJII+LaXUDlTv3N4dJUTIIUfTMJjj/Bh9
RV0Rij5yDKnTQtY5JMA3HMEJJdO7nigqS/GOafy4d8iwrHY8DWq3WFvx7Ku+Qg9Y
HLSQZQMc7BX0qR+zO9ohBxPRZg4m0TO9I9IJ+zMNN8FYYAM333q0Q4distnuBABD
AXqfgRUbY6chQ/b/9VbLAXlMawjUxkP/aeJhw+h1aOXOlcDZ/bPyDErDTQQutjh5
C5gLNcpoN4QeebCr33CemE7tW4tbd9XsHUUejNJGynRc5LVVlpYR8WBTi3fXHJzA
dUzTGth9bD1XXY8BWB9Ih4PeuRs3BRzUfo0/WjIaR0LoVMokCeJmxZLnw5VzG3J2
cio47KkPw6CgHYBo/XadmRHL4HgwEdke7LaiHVjC+PKRjmgWWZFeek9qVrUjoR7A
w2+Yn/30uwtNvDOqQR08Qbckv1cLLg8C1PWL89Qz1m6vwuYaIEpB89+zsBzxY/P/
y+clwy+tLzHnmeXAq/HRUnqWaNgnC84gXUZ8GcnCRgQAhITIBL2VHaEP4UzLtFR/
ceISnfc6FWFmVcEZ17XpN+mrJidhVkZxXXDTR1bQl6zRJO//l63KvdW7JpLxERaC
2viSXbTj2212vGOHjMXnwfgVRVvv3Hl4vo0S57AGRYx0K42TKMmtWpqpxNDclKrm
qRl9XuDLkPkqHQHwk6wbiMyFEUE14dyHkqbTPnkB/hBHIHrWlgZFY1BNOMlujcf2
QF8TwzxoN0XY4kWezj10PRxfqanbGxzLRPXKNFARtBM/nRaSNZtqXskyfWOa7hok
ZrPQYPXW01vH0hFj7tu+lVsrM8ycv1UGy2n8xTDy6G1tgpgBWZ2PmgnkrI5dfNKq
cEM42jaRjZhB1pKIE7YbzMmT5DZn/60ue1ifJPPvapQt/oil9Yo4dB5Z17akRplh
VBWH6g6U9wkHQguqkrDkC7qkZDz+WrHotrqw0tcydmQlhn2S4YxXCgJXyXzh14Gj
zOu1G6hhcbGMyUAKE0X7V1lBheYlPYHtmE/DXB0B3pbIunlQsVMIzQc35czeYbrw
1QSJl2UKUik9jd8EoRJvZC9hb08k5Fd+SfAu8kFKQWrQtbXjBVVwmH7C+DqXA7ra
JaFR0bIqL+xvsofcZH+P+UV1xrzhdVAeQRqZZ1g3lolom3kuiiZPVQ9jGU9nV+XC
sQn4o+aDZcoF7ZBN7kDWVVBVU8Eo98Z7TIYw3cH2SWKj6hM0PRpTgWkJxkJGe0y6
VZRd4XowsFpd1T93jQLQzDe8nEBTX0d92PlJ6dO/HblGdkmcO/i+N18iZcOtLPib
CptD4RtDXVL4Mi2w5rr6shebtU0psiuHhOuKbp6V3rHdET1jYyOt8kMsGhVBzbDT
L9Sr7nbdG+MBESeGE6mN2l6vRz0EAbOxM2fxE1nD0kqQmHjkh2PwGwMXGXsCPJb8
sZz+4uew/ErPk0SzvjfsK6aaFbxGJdn6C72poRpAgkelUfol7xbqVxSwqetdjTwR
j9O1b2nouj80zrjsakpNgaJz3m3PvNz29k3kM4iM95PJ0+kKVA4QRv7Xo3prDPWq
nS8+qrRx3YktW2rkXxnXVcSqm+zfgFWDWTP7HYYffo6HoLxvccvSqzpCw0ubIcn3
d9FZnRaSpQrSHoxmgQ+TMIXD7wCpov+sHT4DFt3mhZ9mlq3gpp9gWSN4MVthbBBC
yBO8Buoo0ntwHxprmbpqTZVsob6JBfj7xOS6qfODN3qL7TzVFQRCtRH2F2JfX0QM
lGQeLtod26wFdY+wUTGqSFNrc2YWBoxgugAId1YLB/0BlfOUUoM1OytaaVKp58WB
JC8nZanKUVQzQOpgXM8PsSjgALNm+20Pk3keowk+3UXSpe1Vma1lUHZ6ZcywGz+O
8EfVlkHaydiggdcUjPZxfAVUJ7yrgqRDtbFHnT6cfNOCRzq67MtayvrQN4ZYZLYI
Yj/I2WIdXg1W7EfC6ctBeXExVT57I0T+kw829x9uZ3RYGdwfvRdtGDk9+qYhqqkL
PzfeKipas4pCHXMMmwnA1odU0SYL+p7zHKfPX2AO02C4dVMg0TU3OrvLpmgawUP6
PEZ33F2yVgtc6CavphGwnKo7FrzkUQN+bAettP6a9qrzdtyVnYJOEHD0w8rt/y1p
MDn4MpVz6WmXzClYnJjWQRzZb1aALlyg2R6cs0C6xSBrM0GVdSwg3RlInlEUKVjr
864/NsQSlVZJxO0+l37GLKVNkOVTtF3go8ZLUB09Y+r2zw33D0+hm8cAO2H65MsV
saowJsCJzTMQqDKxIIgv59hdbhqqYZEwfsXG9q0IrY8INARV4+JkBbfrrfLLEXL7
kzvuy86R/FSVRqPd//kUdFbKRP2Vdsg9IV2Grtl+CniODprElYTLEKdhy9P08ULF
/R1g8NQK3Nd30yXVi+lhbwJCNs2bDhONknov5dreljZUCs3VNf5B2mmiYvWQLWN/
yT9e4Qm1XafdHryjWYdOrxZg5uob41gX2V6r5prq05pApJP40MyITqYUqsop/G0M
gB3g9PvCOwWfSRs7nZHExlrFaeaBWdZXp+omlP/h1HMHEJs0X2xIuFE3zNLKiZQr
k4xQZjyosjgFzha99V5iA+rk2XBe5plhM9D8Sv/qT2FSlLvHDvHd6RG6yF724WqB
1c1BhEltUmlCO/ON5bdoSfSddl5JDrBjU0x7sgTimwg8pXL0YqT/0ESHMlBT6DP9
/NpmeTAdW0yvt7aT4WXZe+8JtSkvzXUcIH3Zca25iO2QS9cE4Q2zbT2a8MpmdPmq
7hgT8+F71AoSHwpBs5qvg4o7rD8ZcCg80ZXdtnxhY/4EAsPp9F6FSp+b6NY1+D5K
jFCU/YDR+wdwGmnNQyZ7+UE6ymlXkIZ2S6nc+4pzhHbgOUNlx7gCypc+/PWpFrAC
4adt4sMX6C38FX/n/tMAE4VGiyc12npFU+jHpsVXjoOyykY86/E6z8WSlfKmzUpN
DkDiEvfi9+zWxgjA1gzjxCceHiXQKEMLFalm1AapPbOoF5NhvfIcYmUAzSlzuwSA
LLFxNTx679rpGO6Mf93UcjeegK3M03NFhNbnCdoU67GtDqGCfCu4Unp9qHUbcVKG
PPtY1zrgFlsJKYbL9oH4WIiK5b4JFVbF/WvsguZBhLkKU0f7S5nzbPAibvOa6+OD
X0mBt4nMW5jj0CPxmth9eQbpqB53FVZf9UGuZx4j9nPFvpGQaasm56LyLXRoaNz/
rEErNVMOMn2VvIBR9zMjhlK/HC29j6Jh/uOBARF440y41aEUhKGr3BpB2ebUk/o8
2DkMUugBBdGSwB1tPpfkFObAWOMHN+CciSl5EBDdbMdwjZ8BjIo8rHrVTeuZc1Oq
ofuxhnN2goInShBg6lqqseK6L9FxoTLvHmNjUqIXv5J+4D4HJM5iL38IJZdpPc+C
+5v4XoiJ2LP3m8PkSDKWQ0AAGTH4CMlbRdLf0HE/7SZTKWOde4yHTcCsKKjwjPxr
i7hTycUC2zQp3FgwCSYjpFCvdlvmMaeGjw45PvwhPpW5QrXEaZoB01cdmitbHOql
EmXyEJ6KpyuDQH3/CACGvItbK7yVh68VzEkd+XVFRBUwXdPzT+ChPwaxMjPhlWOS
McMOvV9khVnrJ3TFO+/2i9/qgsuaQdmX/lisiI2yFODUzq0wRysRd9GbpvXcxC+m
rJHMItZGWvRBx8a1C5pkXsJeupS/jT/dZ4NBiMavv+clX8EH72YqXm2ovopHfe/0
lVfE0wYT/QIYNXVtR0SLVWOECfFP0yEPsd1GrLPHbPY0x5KfKJdsqq5K2LsFhV5f
FGO9AFm/vpRhop9jyjdsXDm66iw7zyhba9/jPWGLoxaMvdUDDDwYXmYzBhzluxvm
yHPQ49MKT0tzIMaf/XvqrXiQPt627PmUQuiYuHnwX/xR8LToQ9ClLJPLaxRYFLm9
DLdqKmgJYCTW2lmMnYc2lGs7SzBirmCw3qmWkJBqsrMN27pF/5GpO/7gtOLOYahZ
SzrUs0GVsYPRorvIS7wpGfkassk5L8nE5+mH0JtgO9t5QOwi3bhmIspOuTtVyCjv
bc5Jv7C2PkCr1gU95aO9Z3AmKpUkMvxlIr6R1JWTFyXlRBcQPl3l9LLBIWK00RLb
0U+dEAOBYq7H5xuMil6Nr8HwlxdLi2/4GnZqZMgaItwWMkAFqhKFWV5QfF3cyOvK
CALNwaWD1MB517kR/s7K2P4SnoSf5LlFdEfnMhjY+yPpFUUje8KnWrrSuEI2BfrN
0Le2C+elgdHNC6yZlVPSOEoomXXdf1Mvrkvy6TRJweZPAnxRa332tKHhHP3JSVwB
9tU+ewrElwa5ilu9OiMRIN4osWj9UjwYbNpkRSZ967nNz4/xMFFA68KlNeYRl0M0
EbWZ8RrMSHCW3L8z3CWiqKpZ8qTtSnM3yLdw4EQnmMX/RkJBHFlJX7Wt/X09fIYr
/N+7ilZkpxtlnnlu+xVAEZY3E4vss8FkBS9sm/7cSPzumHh18aBsE14bsoytwcLh
zEuz1k+RdbUW94Uu1RlgdXCrkYBe4lk+kKsWAU8aVv5/Gy2xrmuTy6NBcXyhXdVA
y3SUU9Jgo8EbOp3jIJ039dyfjrsr9oX5HpNrfnPGlPxOtRT36sK4S0Z+/m/dXSJa
E9UWkGF4xdZe/bjgOsTQ97qG+SkzbH3+7owBdB5FmL48stf1GWn0oAj34h0Hoo/I
djdbji+lKjuW9XwDjWQA12gp/VCD5kNRGTawG3l6v5eJlPKdL2mXljKT6sDB0YJf
2a0Ru9CGTQnPFJfMN2sIhRuHUbT2gk8icdRVQxG3cZejKrekOlCCK1wUQK8JKhL2
BKtkoc9awgURgGhJBnaen+VC/k+rOW3RAlwE59eiB9uB1gbjpJDU0wI6dofLfpfL
7v6TXE13t6moF0VdRHYD1OKmRmm5fKR4ktjCkbhND9PIyChCdgdQqeKP61KR8TWg
qdqjh9v8Zh1mn43Soli9yRiG8wZGpL7bHmgOY47/FUCUAnHg6/P+08eQN7L/DOrQ
a9wjgYU9NYFkfORAwZBENwENHZCmuoq2EXO1XwdohXQTvSlVsI4baYr/EwZ5gYOr
SfDE6tMPhMTZWKOuXXG2VRCbaT3uMtXTjHS9YzE9H8WstPKLxy3Ec0znZ2DhN5hz
gvgOyilhEoQNJHxP0bUZ2amj9BzQS26qPOklkgRK9kqitnYgmPCjM+0SHuQFQBhE
//kUn5tqyjse3mncUNm1NKmuVEoNNLmKpSiZZHd86Fk/qcnWUYFM9z2sIJVx5pFe
JGuOu3Ke+bIfl4G1rsyArcRmmLiosJYLcVR1gWaAr3hw8jp1crjjBVoY4zE4UhWf
7q/DE8zhHoZw0m3Q/ZDSM9Fi+bc/S1i++EVKm47xDww85gPEKXDgu16s6xpak8sd
oozDdOyRXhptbYaYZyR7sBnaUOAuVwd9t7PiLd40fzUuaKRklZlBgrMFKmI4xVKV
ZsLxznPFsWJjPlA9zlOwzTvztU1VJmKam259eDcy3Uj8maItD7cqk5/AwSKtC6Gc
hbYZsjXToquN4U9FDEY1UHswps7b7bqksmK7VK5lxVVQB3wLnYboCQBBxqtrSoOh
Kv8rzU/BvUNiEBFAxbCrul9XQqsABdev7vYLhZBfr1ydP/LgldU+7EzrDQ6glRpg
3E1jFWUtpyzM59ZVl3uP4Ej+mzzVXJod0F/9q2pj+EYttnS6SDHamUdi78ISjJO1
XSaemg+jHx8jKu4llT4BlWY+G7c/uZ/0OLNvDRGXus+hzX2TvmIDT1DBIiNIUj9F
Jax67E3P1Da7rE8V+Hjzm2CzgOYsOKxYsUm6Mw0JYA+m9cPddEw20C2txMwjf2/R
CkX2j6NGeECk4NkuOLFGAc1Irm0eG9aO4CM0FXbevZKcOV30q9QSfsXxNJWD0sv7
Vz2+QrVokhmwr2mvOEr89L/DL/lVrMOd9p+4SUSknmtl3hMC43jLlB5NDjhNTd8R
Qi2S5EDXCyD0mHvRGqIDbILQDXWU+W8FH9meHMLDh7swAd/1MHJ/meaP3RZIq2h0
zNIPFKQuKzeUbHtfiXM4z05IcRx6RjU4V3B+9sTEJXXmAsXWjk8r+TNR4sFgEtFc
cW4ImKpHyyP1m9gdlEvF1R2xJVvwFsD8+G2UbGTmZBbCo5lq897ZB9sTiiFtQ2yn
c93R7r7PRoiJS7fEwWaLhmjtvUJFyJ4LfGyLOjQ+a0C6Fnn1U+R8djW+dfETYCIw
VKU/SMajtyvHk/wUIq3CZg/87wiXeermEocD/W1fOhu4nYXwU76LUbeOkEY1CVz8
xTxHW76jfeVajsoOL6shD/B4HhAhW59i6ViYmdKdUQ8dmyIdHzEIIWbFYPPSG6p6
R9dBlypN1zRxEPvHec3SUSSOjxqUUaGBcpmAA5EuzrkHDG6+fKpHslyo+/WFFuc7
eo0VY2n3yePucf6AFLsnGVq1IMI33ZOoxwm+yTRl8y/+tTwNqcDpieJOO0hjJEv6
Mi0nxcEgpS2oad943A50Y2hWYot/P/QJdsY2oG04OAX1Bq5GX3OHVLJlCUbOi51u
9W7E05t8hzB/TJxRubHlqxKTy09S2Czgpb0vVwDUghW54LmpD1mXzo3V8wBMbFqT
fkaJ9AMuOk8T7WbH9ufcitrPHMyZoT0/GYRtI4C7WOs+z1gAr/2wQkz03OELxk1V
+rMsPxeU4CjbfwDiNkQJ9ms8kX0ePGjeHpKtnpZkCZYaZQDIIzb4ZNCJ7z5N/hQR
yjE9tAE7i7G2UhiHWSTPYWXXtvoKyIcDnqnblB9v8k+RVJYOEsrQhKna8i67HGZL
32z2CxhcN0BWhpcbcGGhtvR2HMFdqc4T9eCZhH8bwagBLrnqjTzDqN4gY2Ca7ok5
AnbeS34tfeZ9sU4f0CNC9arQ04NbfXVnllDAQXtGPmvnvrWGY8dBP2937A207K9y
ALIDBc6d6mTc11HStsHsp0B1iWIjU20OewYk0l+6Fq9fFqV+3jgvVv2hCJJ5fAQd
H0aSVlLagcj6+jhxlMaODCTg9fweqaW+z2URyz4UF5McOJGVJGtqBP6V3CrGaTAc
TRXAN0F2djz/tPjglAysumFHBmGREnBi1muOfpZhw4BnerurcL0E+YvNNX1zOagU
j28+v5Be9bwtDf6nqFdudDazI3YbjzyaJiqOxTGV1CkbBkhdVKUCwuCJaLHLP2jy
5HuKKX/ln++QDCzAUWm2iUnebepJb6+CAOv1zufwZFfalKftegRndCj642gc8rwc
BAuLf8+ciCIKb9w+Cmk6bNj0k1TyQfeADHjY82k6mF3WFbCZfMSml7lp2uqWB25C
hDUUBQb1dn43aoRnby/Qe4JgogEcwwDINzwg6KDxdW9ebj+PnFAa8q917P/TzntB
tKV//cTJ00dbUTNQeJk7LrGK4kQ9qYYctuUEnfyp7eYv0LNtPYoZGtMgUZloawpt
c4DxzJWa/u+1xKXYoqWF5za9Pft4lGAWSv/gAiF2xaSidE+avszYZfII/q4tLPi9
g8WYZJRGJFaK5kdJU0MSerWRbkeBq9YYp0iq8L7hobZdlItx/hNtD5tZzbYsj1eY
IA7V0rHg5zWt5qpsM7tYHiEjvAMqtgHW8l8qvu0NmJ9+ktMtVCCwVWvu5ooYQKmr
c7Ie0zNGADiYaEVKpEzhXw2PhEtTMkqbHmm78S+N1yYnwCc0iqBncEz+EsAfgFAW
/nVgFeL7mkkqZMyny9wMNz65NTQsZ823k3AsauGPYrlGkxV3oEFBe46DP+NLQC3h
HcNMRMUIh3T1ugSFA/gKhnTY33j0oPG15GwPDBBZ44dbK5ZGyCgz4wzbHXKEOL+x
UdC24FK/iD1YKJHniHBIiyQoQpNiVAMvVs+WG6acBt7iLlDJnnhMt6f/yzlCJaYG
wbIO9XDYmuH4DmRxCkDs20092PrYNytOpETSJuRVKExFQ27W5tWkSIUgKqqZtDhQ
IKluk4PIgSqjv5ypFyrko+eIZ5Nsv0/dgVOo3PoM87S3zUDQrFTHl+fpf0kngttI
LwQ4yMxZabnFSHpsSXKAmDKRP9NaHJdA8C2LR2G88CjgOnl/386qRzjl8qy3LLkB
ziieqFkKmVt0ufA1PeDNFX3pnOpxJw9DKtxmX0L77jhgKzkZbX+2pfF/RnWey20R
BVVQPoPppK6VXQmS+sBN2QmqolaXy8DfCyoVZOEtDm6xXkIArFS4Qj4yJF/nI7ro
ywOcDt+p0tUVr3OLQCfGbqRS9Yj/JYc/HSq/IMkiQamKPs5JjwmszW7Y94L/FxFc
x2nHnorwJr9FYFJKIo3aoHH/ZQ+r4aMzPTqo2UvEPeOeUYxhoVhHzpXT+pBcJoIa
uzBJB2YVwB+hBfq8kDgqoWzmtoGKLyT/Bb59rC6qsj1nLS3J9rMR/fdyAXCPHtf4
UlIaWj7BjcATnntycX0xKH2zddwzCPD81GUlgF4xdPGvnaT9aFlv4D7yy5b63YvI
TsgxmhkFgZzVImmC6zGTnZ8VcDBLn2D9c9ICp75iJuwbo0e3VvKpfJl/1a/fsKuS
Vlho1fnQXrVoLAJvGklh/1VLTVBRRlXW+TzFUkEhJhMhyySeJcib8iHRiplfTLuE
JdCzMuTOqN155zaW2TTLYwzNOXU7PHvxnUhsjm64Fd+UAXHBFZs/KP/DO9zV8DHV
5zJqOOYmiFYeQNhWikbR0yOW4AlCWxL8SoGnUuM3p+Az9AtO6ivVbv4xFJdUPTMU
akQ6p/geLOrk8QCVv4DluRpSiT0x/WsFJJr2EtsR7Ntm4vMjMT6IrjH59hyq5U9e
9tlDfvwv7E41W/+MPvjEGFxHIaKVM08cz/zzMd9N319ok0M0vSQ5R7+3fV+dV2cT
uw4Trwxvlhh8StWPcuaKgMKEGopCVRdBcqywyx49xFXqPt6AWKD5gelNO5TmL0Hp
VjUoVPW0olzxdvvHoR/+RkjjWqyZYtFrpffHnNwO3k7vEm31Fo4rjnrtHdgMlm2z
tauiMMUFhn189+p4SV64MxdY0dM5scLkAClXnLlZHSFQqCtGIOtmeu8ZELx92O+l
+aAUHGkSmWUXYpPnaUEysyocEPo++tcOu9kJVDnz7iyyCbFOKsEvw7vUCZuy0htB
btjDohjTNbe2Lir7pHJBJiSTm0Js/YZpAqVATwC15L0+Kn73iYc7BJUsXzEHBMiU
LTdp1KAR9lc7UOmTfPS1KDLd0EQnaBylCWnx5v40b2J4cJHW8ZJNdMdAHAhOxAdV
5iZoEl5YRA96GJvluXWP7GqICvR506tHjlRM+xH0cp8toJbQ5AKfiejXsp5Wr8E+
N9rKZ9LcMfGZ/7utjbfPH6ihW9o4H2EYeao/t1ASTDokotwMTfVrS2YKXT3f1EFK
ZkS+zIN931qTIhHfNTn4asAS6VhjWzJJkPy2eFqCM/fsFPqjwm7EV5tCckltNAR8
LyJ8rPdyjNpIFsmQ8aj9RPjL8Hd3yWttgDQ0WdPlU69CcOrwe9fR6A2wl+QP7Xk5
Pl5469kqbloLTQUyEVW43z6a8BxbYGZMIh5o1F4K8avECPXSsmaKYVMUqEDYAhKU
M4hwgMWQvjSrajSLZ+xsyMFfuiW1cRRpRg7umS1CkACA/PXOUeuW3IsbchsimagP
66RPcWrhHI8tzvQla+8abXMB/yVIBYfXJ277GUcY4mN56KxnvQSMXt3dt7JNKPvU
1pbgYPsHH4yhL+3D1MI6WA7+Yr+8dyNv/nj2yiD5Xml2kjJPw+7BzuQQ8MZTkSv1
HNG8Ka2xR58LFipZkXyW4D1v42dHVGfheHz9JzTTEXSEqnWC9QT09+rezw2Qq1/+
c3CL1QAz6CPjnfCwFCPsyCeF8wy0vALToOyOWgJaJ78GM7cq3noMBTHB3y5nQxSp
u4oBCvJGryjn8fGnLgdEy3KEowkCh224+gzySCyEUJY+jJF+H2AgDtrAUk8DWybh
oIH5I0fG2eWRCfILJ1eCOZSfGEbYyABgR9CFJVzWdKyzmGbj4gAfHfmA0hC/ia1p
UBJ7e1iF/a3sYEwYOIiC79nK/znvthOze4HAds1TBQYADe+rFzo76gEqMw9/u1n7
kqvvnOoauMsXt7jPhDM9ABxTTmv1f5lpfgI8gYayS3du3qeWcHZtTfg0rjylcbzA
Ar0G5oOzipfL4E19tZnZlwt/vJJsl+yv/GYspg9Xcq26G2XMF/dlWiEyiNBozWel
lGbwDCDw8t3OeSL9dMj6mWjdsAn3qL++DXi2I/8CEdk7k6lbdpkU4aS8aA1RFutU
uzIOkfK7EFtlmpESKmPRHGHVNxx+B+LVxVk4+q0o1MJJWUs32KV2UInqWLTJn35v
ZkoBLDxpwTcj5JH1rA944pE4I422jRFwRAWnTidAIpwTB18e3VmECHOtbrgT51QV
eJpiRl8AJFPRxT5IuhcvX5ZWQRFrJu3gWEeylPJFH4zWRODlVf/uVd5WVDc6NIPA
olbjiSvYZhI6PbQce1GeqoupNbyyaa2gnRYwFVDiq1tMajSDygX4ZsaQWnv7c8u0
bI4WV79kGh6Kbg641z7J7/T5+bu7H7xt/al69QR1pFR/SEpYPTg4GaMWKDZq9DAa
RgZFud/NhwZvAm8pWx08oiyTJX96n98CDH+is7TUaU09mgJZTZodoPWcIzuKm4bC
Hj1MF1sZGTHkjFBuBtM5XI71rDKOOqbWkudjNfKsODveJpNzPBBORNnbE+zWmYh0
ViomxwmbJaptmQU2/23TG1qpYQe7xAuXTvDnv7km6o0YtMOVxX5cLrHKNJX2h26X
V4zVejW9jS2/d7nM9keyebH/BhWLkZPju2aDJfU60Dq/V6W4hirzZ+CRINgyRbtG
XMmL2qY8vnsH9wWkc+hlS1R6bm6C67LiNbdtsPDFiRrhLtJNWScXMEjENl9/9l8s
u3Kh+fuEHowzuEgJ8EzWOR4goiMI/RWPpjvXixHAhF/zGx79LfOpbaP3ktCtaNmK
LyUzuLJpmPsth0YJGxRQjO5nCzlnzx4HjT0QvUdCTyG6LQCDAEnv+KDPN/SOxyjJ
Xib8f60/EN/vtB37ItcecWGT54H74WjB+7Dv2ZcE9AJuoCxWuBROZ4p4+sARmlCb
Mdjp24n/DhCj7jp/VX46btIu0kYyzQ49T0AO17sJgkdLq2Vgz+7VCN7u5Ydalebd
LTs60tWj0ZQ9/psdIY9vC3WzacbqhaV+GdrN261mrOj7oNkQTSngqPUT8S9NKtx8
H2jOIuLAuD1tR6FHHPHmaRrNlEpligMw+T0FtOhSrooJFF5Gh7auUpL8bp+MWr++
H0LC+vVbpRUe1iWLMbSFciYfN/rPTc85HcoKDSRLMnN1dP3yEme2c5xZSEoydkfr
Cp2+h69tzVN4S1xrODEdtod6vlrxaCpYOpWGp/PiR9jZN5ng9nl9DRX7x9OhhWMm
5Co0V43+jP4ACrtmen3ZYmZDjHbkBRlMB0fvDm8Fi6gr7Tg0CCFoatCJaAATcWCt
31puz93bxakphbISt+d/lq/WLdlh67+oQRhjt5jE47hMwSx3Tjg+TlgiOpmy+SPo
37OKg6U2fi2oqgLNkLLbV2zgR0L/zQJlplpnsked8pUC5CEGltCymWh2rWOaONJL
CHZs+hg/4zM2zbASOzGGkrFzoQY3pOCi4J8nIXicOtTS4l5V/kh6E/S4Duc9EWqP
JjvceBNkAwwro6qW2VZFOlqIE4n1SiEPjXqM3RdovWexWwk0AcHchRlJ8nBRui2b
ETyV+clPZR5keaM0WuJ4hDru95Xq87Nq6AocMLkDxLmf0MJbX/p33Z9JHeu3bvPP
oNaojxm3j5rJSQ6FPLFWM6fv7H5cy1SyyhZa1mjATXCPzxf54InPqmwkVREBL7xJ
9KDGiZf7NsArsm0EdSIBFYKbVpHY1sPJuvptocUpXxMDfCh7sFxKWJADqNahd5qk
CIZcTAOQrr/9qI5mH9KfxvW6dL1fhywwLOgWdLZlHCzqG3l6CFyXiVBm6vsBpc2B
U2dr2qXBlx+zMbHYtBD3cG6gwHxgVbDldhZwxs1Zx5jsIOnP4I8ui0x9crH7S7ah
U4VoB+LByj+g+YnkjPyFMfdAeXLJ2Sy2s1ABtyktBUq3FbK4tHlKquuxDLDp48AZ
sKcXBeMzhmyt1dvAxsp3zNm8EI1pvuxtd4IcuOdkZJP2q6quAFQvavgZIS3zPJKc
zlVRpTq7FcNNZg/1e9Y+HtI1vdqjpE97G3An8vvL/Xw4WZ/SK6561lIa46a2eMN9
CzN7R6YQ4fNp424Xoy2M2iq9yc1l5hKahEm4ZOOgCqWKF2gg2QvjlLWaocLCr2mQ
PsPF+/84fvdAcVwjhM0jMi1+ycjnb+5HsoCjJhwGVviFp5Dfi68FxYt87f/UD0Ce
KF2NMiGNaLTHSV7TNZA8DgzA/PJp39Cu2qB9Kz2RMincfRB0OxNcqPwcrhuQkdn/
HLMwWjfPkBogtJvSbDeWKApIWU0TL79qWKXbAcDARmLSVTmypTLR/Vgyg3PFI9lq
27WTBi8Kxj0QYkRvc/KkPrtXj+2jZGrkdHMODo05mpdLtKbqg682fnD/mYVIc9gU
AC6M76MnjVH0+56c1aMXhOStWX5noNDA5/n5MyqkwFrpQUYfB2jkMAhC2mz6ioDY
KC1J8WCTkf2LWmgdNvn7rWAJyi1XbE9j8NVVWbjdgTtWhQD0USCGaVn17v+llvoG
4a5lgnQc0Zh6w9k7bJbF9eSkFssBt3w4ft2rOViYWTcBxe2xnz1W26qv4glw6HSV
j66yKmnMc3lvCCrBzEM7nFhqHLmZ41TW7rSP4+tJnR2l7JFejdsKSUOxoJysU/fg
8y/jMJGVk0JrmqUgA+b/5ArRHLbo1AMFBbEWzKm65DPyLgOrxW6h22T1nRiaj1oO
ItzkRmrIufoiFOawnOilTMhp0DpXciBNKcaBUM5q3cnNasAftav90MJgfWlUDKuv
FoKOKpYOb478sWzGymGEXOu75xKtjehAjtSYaMd+nY1A4gZmgDKnSiSyiF5+MWzr
kzXYWoVdfTUYA/3ecr5w8beNF1bj0gGgEuBBtSSL7KZTpGJM07p+AUm5CFk+vfUl
gC7DjYNZ3SJ4e3s1IAecH0l04zcFafhi+xR22oD629mGSn2ls2EucKJawm+YFo0l
7G1MKM3/SWT0fG2rk/XbpZUMd8i20Nv4K/yDGuYgijfnLffgGPNr5GYpIkdvM2PQ
PEjGhlMYmi7TL2c0+cexZBqEw3xCm4L7SLzH5KA4ywoifG5DTMKyuxoRN28pn3wJ
2X/oW3HyecQyucvhGaKJugqnK3+pkwKpLmGlVXvA6HWPfq4kZcuX2ozGp4fM1EbI
2I0kQSw7BFJgVJJKN+3a1MZExa7T+3fuNTnqNQ4afrXhOgXZ41jYTr9gmJ61/bOn
omPeA0qfZlDSwtNYpBL3e7MPVUYNsABvKn6+k4xTzlNt+7V3PFLLbngHl1hjbzJF
E39wqXEOeKRq2x5rlOowCH0z59By7v1gcbpFKahFKUrdsf4GgpA7QUj+xcGTSlRg
XWRzml3oq7j8GotN8aRFzCFKq3CP9EbcSXq1wGsEx3v44qz4uqqXEJuqk8oErGGs
eVfOVxoOcrsJGRxkQ7nAgFL8zTPI7+ngDKpKrgGWfA7voDs27LcIUCLSZS4nsSxU
ccsrASRQ6mDRljAjVhrWohtSwRd6JstnzhnZ0n/XS1N3QOyPG021LudroY9iRgqU
4Dz10kk118LSCi/xGvNTxc+FLrSO9CLFWxR0E9IFnHbQuIOKCnSeCc4CwbZ8kFw5
giwYiwESNZY/WzJ5o/Z92mmE+xWxQSkyHp1O+Tm2CCRMVXuoOKwkRutdqR8d9gQt
PJuLXAhlOqRruYzUSMB1T7AcjfVfFra/ve0sMCdUoqbSbhu4DQ7Q1BYn6i2ps+nJ
WfEjmI7MNIMru7327Ff8nAJdRkZPo9pjdUlxfEOOgAFLpnJzKZppAcKvzGz3FXJU
aXbyGo+plBZ0yllkjva2KUDVtnN36JXkjYl1KPgCT8DZn+l2S8S2ldkhjS9FGakp
ker0jCSVD5pFBQDweX6OjcZxxEEzKa6e+P8qEvDKMoL7iR7tGWfHEwAo3IG9hCFl
TXzUb2ItsdMw4bXMsGmqzAsopuEiaSmLqzqvSp1TMLl/9iAj+gEhCX/OqQeqQUii
jyIRuVZfqkH1aRRMv58MYsQJGORFRKePiFwrFwHBSu5Ek/CwyYxYsSgDCqUE0ALN
55gxjisNwhxopKOu6dNj/9xKyyu6Ybk05kOeYEzCoeZF+jNxxCHwwE7gvynGJRyG
SJ1Xd6Ob47RApE+sy9Iing+b3l5LKWFE/FJkQQjTc7gq5e3PjleP1YQAM1Ondq/D
C7NCoIiR+2tNm1OB+7DJhgdAwpu8QBnrYKgsUf9ppv+6Cdy5xJ7fBf/P4yvj0Uuv
O55ZMI7X155/+1veAh037C3W5HATetYgc7YvCvOiUXVdheQm1c+NZMDnyebKz3pW
78wVfzPPKxhcKTF2HC/Y2y7gnXjCYr7kuHnO64IzGiePwB+XoZO4q6lFLkBqLomR
lQV7EePmSiFd4/CVw3LMc3qZznHKwoaSfR0VadlBtZv6Wt5fLvYL6KpkU1SNGg3S
asRtLHWxloo1i/Y/zGzF2n+em3fb9UMKKrex0x6Q/mXbNViiaiI/Y6F2QuZ6lEHm
deDWJ3kAJa31jadBQMu3+fDvDMzAWQ6K761YkmJ89V2MZTlJGIp4jGQbSCS52BLa
QD73RQvTpDvYIz7yzpD5UZtaFqffLR6ixm00qbw4Rwm63iOlrrC5mY1D6JmKivTy
YSg8ANY6yMwlhJePcSE21e0QJKlJFMc9gPF/k5fIZJIR4y3URmeFX7E0JFi04SLF
PJhIwKdDerWd3mZGrnSOjEWf7G7NKKLvqaL8ABuo2lQeERC6yv0MQsYSN+vAiCgH
Q4gup8YsH0ojCFdT0lgrWPCGD2X5CGwgOr0BjLdBRBLmXmmdBavahy8fsyWi2xsE
huWH1iYzTsTkkNV1Sk4UMcAitY9qITdtVSwo2a8bKEkp7/+Qd+6tolICXxoocLaS
5INRnoXElYU6q8OGBGUs30LQs/WDLwmQrx7JtxJYZy+JhSgVGb+m2CURJHeKTllm
r07WmKh6nRxEPkMNdcoEpOz8WHhQawyGQvgmB/9H15pE07IW2gYGWLc98gWsSekP
xOMThGS+i9BC3Oeex/Z9niAIeqPx4y6iTStGgUI8Zu0KXze1BBPFQZBSP3N5k2Fn
tfufhxf5FBbtmsKkNcb8mmMlfxg+qmy5hkag2gGG1jS08zHVLadP6cYu2wUghdSr
HmyS9vqIj0/bwBz1ilGMRWPW+Hr+WmS5D/xiTSzMsmvdKwLFoHbGTkZHWFquvJZe
w2UitaIPON4FbdNr0D1PAt3b4wIvzk3ms3W4i+Bn9rPytNSQhNXf+zDS8QPmLvL0
S6LBSmVE7FGx5nRrA+sI/vULs4dH+c7gfN2M0d9Dn+oA/DkZxJ+XI2ZoWOgZq+OS
bIq2Hbpfod1PC4ygcMBAZL5R1DAAZpQeBfcmEhoCaaihX4EM9D+1pmcszF5LwbUU
QbJzDNjTLDlhMgP+4fkU6crP6eoT+OOUb2g/p8YGqR548I1XWG+/QhWHE1oY4oHr
FGThDyNu7AxcSsx626fP5E5sKOGaLj12hPJvX0QpOTvhyQeLHmyTYm4QkWxkTLay
96Ls1qXN8qv0xnGsNJubeY/Ko63QUDmQ8aZqXVTao5IWgR0Kjl/oKsrI5XPK65zb
Ntv2/S2fvzsWVcPOeDlV2AtvmiahtinnDO2fxMVxr0sT4z+2aUn8xg8fG5gKBlqj
khntqLWizt148PAVkCvfOr9A+x/N83VZ21LVeGaRyuIb3UtXyCEsjcFeXOKDrQUK
I4HKbQkuLfPvEY2n/lI4f5USshcv8vt7pb8bUGmB8EesQvZ+0q7MKkqLCIVD8m5t
0uPyYCgR9HmynCi8i0pap4/LTZnRg/veV9ZZ9hCuiDhWzUcR8eU53HAtZuyS857+
Dgj0n/06im2+Z1cycp/UsguOWpXBRnBYvZuXKJ+QeprQ0rHW3hyJoc1beaTvpmDv
qlkbdiBUg0HL6vNeU1VH2xzdwbxr9cVNmebC5Cm6RIyQDT6cRXek6DSjyRMmOIzE
ITq8kh/UYaYU20q3TV/JX+U2ZmhoUhwAR9szvon+2kTneCyoHL/4jYUo4tFcZpoz
wEnWwg4qXZT0VF8sofSAgWAKSdVWl5603k60FSFE49r3DWXYslajW/X05MOEAeft
YSZSx8Jh9j2lCfw/0WODCRBgi7OUDtH6HN6Liojy1pan/s0/1RzPij/u37ZC2P1D
LuhQ7/0q2m3LWINgtx3P4hsUQrqzMauTcGs7Ghh04YSeC/2hXinwqDQNYZxZ7Wom
FklyoagRUG9LyWcPcEZ/vZnavDlkYPi+V7bBMj9Hl3vQQT4gk1WKJe6Y434Knsod
phVC2sz/Io2+Lt+KjSZvxqi1TRPaVesoJjjXiJMe71REGa1JqFSbtugLEMmGF3nt
xXuiDxOlYbkTE8UUjimzmD75TubrmdYtSxiSgjINVbSW9G4KlA2rycUDVD4WiYAH
YomoMVIjFqg9GvFpKMhbaRITMsnghRwf+nOYUB5KukH3EWUlr+XEgzzslbWvBtSh
yAoIuTaMDwvPs6ACglXuM/3cfvuSwQPzImvbmA17mN3TEmlUVBpYP1pHctwZUnKQ
G9QFKlg6h4MKAzreTQy5AR73UXc36Gt9CA3VRF/C0WHmW64iVqreZhjmDp/z3sji
Rk4xDR+Ho3kftO4wZ86ctekYB2HcCwtdk64X3zpEWXbCQOzFw1n/wHkkTMVIg/Da
dbyhnez0Xblt//t9i8u8tITRYme/U6ZAiDc1yyHmdwwKpO7xyz3rwEa4wF0O6EsU
if1kDxiNbwNqmkJbI+s6WoqDN131YFER7Gannyg8up9pHzvOKca7uwPjGtBTT9Fl
2/TGQlD//txXe+mU9LQlJzhO6uL+oeLZhthZNfZun9ZTVD4tcSKDGcY8DExZlekc
cfIx2frbV/FsER0nIxTqPNu93v5J/6aRU8iqu26VOL/Uj3JVKGyVJbNk6wYPIZmr
xr7+jOGdmrKoqYvwNGc5jkcUDDfQdl7jcyAK8/9R9oIn1qmD3mSNPEVZDqSRQKbV
r+dOrdXS91CRmU57J25kyoEQnOyqWtUM0NAraLJbzjR0z8TtpBD6rQnPDY584dx9
Guy/SdrBOgiCJJOtORwzgfGrxHmb16zRmv2f4hbO3K0g5ES4MquYJFjSWPOQeYx6
G5vsfUZAs3Zc4fxBcYr5tLSi1c1y9TYow2X4cXftrz81hlnKwPlJJHu/ITrF5r7K
rJBWyDFsMbv8A3UU5QRfY620KPD5LnMYSNsHDOXtRxu7lPuTX87bLYjWGdOxjre6
Sf+2JLpwKdMyPHw1nGSBCt3bqkxlx4eawkzvnLAZ8SmOHFTmN48U+hCQ1WXLBQpC
jpALRziPrl4nckwrkYBEA3qNdw+38eoqI7alxevT0Af5N3duZS8kbG3zodHi3SXA
mcMkIrAXcMhwFxyfXImOS13lXpymq2iIdqv1LvteECSXD78xFyNvfuE7N8T7IlbF
ioRpHXDVQBClSNdEjmrSZrANUnIjlKMTV7/h5usWlYjrIEzJtb9j4wRkCqDNRew8
VZOHZ27XTE4WsmT8Ru3VluxBwxI9QT6htEuh2iv6E9iFSSsJeyZuWdB+ZcFraa5c
nB4NTI9I7hWLhx4DrDAAanzBZgKhV92JKaCmvqEZJMt1bu8uzxBc801hxfAyakhO
D7bkCzMLLz4k4MxcPvNQz5VAUnGcLIPxlHKpAyD+fSknXA2YExk/himCO/G5ULdH
+M0aCLET42QGXQO1Trl7OSY0fa0kzz0wCvpAKqFW/PSww21j7S5succOH63+k5xS
kPu77bfJ9vUBfylznnkTbw/hZ8b54nqZWPYR4K+Ja0P1CJVItBlgP0+jo9z+euYx
x+fB96oS1gumXwNu9Qris7OaIIb7fhNYfY/MZHrD3snGsSr8rukIUcCXO12mt5ZB
8uMolNRsRx+klJ1XZWCB9cp9WThuHx1ATnE6+fjnyKWFx+rAH4N0YC4uqCq9JNNW
9QF7x7qTF2c2p8yEpy8u+6ID/7MroOtSrvslylKWpHNVzw3vSL7iaIVkyYsIm42I
DeRKs/7CDhCuSlOAxqwoZAsyoa4unG+XG8TU47/+hXyiXhfzZlP52IsUCl7L0Jto
vLs7dpIT+Bn1FtOX7h6s2SUjSMbg+bj4al4wYu34Py5Ewild7/LCb0yXqyZnUMqM
rPPkQqQS5XJqSZN5qOJDciImqhR5pqFszwipjsFp5/bQd7CmfogUFBwugkaXFEHJ
qA9iesZo/P9beVvEbpVx2XsAF9GjDIgtx+S3coQq6Vc2FwS2JosIfx0U0szrkmCE
iahuUvkvMn9PscQqkGsvHDpNd40k+rr2cWhEU4mcfsziiJV7sRJ/3AtA+tIcNCG5
3tVFJeHSOc5YLmv9Zr1HmrE6rb4eYbeVSKna1RhEdsVyfdvlGd1KXSvbyKuGKX6H
0vbN2dMnebtGGxBPtm9pB6ycF14kOL1Ren8BE9KugzDhRbqLIMeXPIICV25OHQyH
Gh8QwCmGoTMf+1vW9LhSl1e9vgIvFRkasZXWgeM0b1UW40kpqavNmIfl7PNjlPSs
QGl8Pm0obJ5VwVzUp9HZYZyQiyfyza5hCn14VLk0VAxzxkvWku1A33WsDqSzLMAK
4BxsyqMLfJ7bzfA7m98t3ofUMenSA6H2U4S8++DBvn0ImTXz1gNcIodXXp+S8Wc4
HpjEkx6SXSjxjCOEjEKyGFdtYLcHknbQRAirodNbO3cYIfaGmnD+NyMT0YCPJXn1
3t1MS033cjbpJBCUJbhC0X37FWGH4W1K+kQAUfEOinvB80WBGThxDhkf2FAk3lbt
WDPePjusEbAH8nP1gO3yJuFMFTxXrqZKEFH3b5PIBGPChwBKPGR8syi/6x2VLhG3
xmz1oKMbxbmCbFCsYBBeoXwatltfO9iOPEPSS36zCNyNW+G0pLtNogilcwbMEV4N
ziZ0wT0awIxVHtSaeXsNuAooauOCGtQ/dQfzsjdfKC1rBpzyLbtELx2tTmJs/wtG
TA/sbCbFmZKmUGakIf0j9JBYtfsWR9Mqd/C+kYmbI6rpjMy0jZbymag7bXSwAXlt
wcLaaYX0GClqiyUgZpVvtvpfOju84kNDDgFl6BJ12VqMKVbNTjzYVPoHgRQEULYh
n1Tqw3buEMEua3VJZ+pX5X7eE/WAl3nrlxSbsHRzb+NYu5Q3Q5nxkFWpDbPDYz6u
bpgLIgzwXR4gStTkJab6qkHBnH1eAzhO/hJp9ORCOhF6Jm89Pzg20th5Ava4RkFC
2Nmog8KBG0fp+e4IPuIh8EG3Dn1QkLaQqMO/Wu5+pLnVX6DKs2ICWV6urdm0mjL+
xaXv82QADPkw+7bPrfgGxNAY2D95wDE0hulHtME+I9mUf9rH2hZyFbFuznuDJYZP
QR9x9nFx5NKTwJUTury7wxOA8awE7f1oDGFAWrBxlmGHC1SLpRcUhb/2Qg2fq5Ba
cHUgkLq2xY4Wcl7pUowblvr6ye4I0RbR/xs2hzglc2+L/8VIYrPMGQBa1ffa9J88
gyNCbaFiBeoAoVFuZc2308kcmr3bL+S11dAnq/WJGbQBMSQsIKwxQ8O88bv1IkW8
8KE39CfovTm9jWu5/sF/LEqMmdd9d5W2sgBRy2cMB5J2J+Al2X4k/j+8BSoK+Z8k
O+4wEgK78Ff+mscWrjSWOeh4W1lIIDh6r1uBsLfuS1oPxWhnCkrkj5jdzXIlmIvc
VlEwhhWgZYy+zsSz4N4tVO2hQkdZASk1qlRm6kHpmmA1ItyxRxrwGY56vJr8sevx
FRKLe+yKz33Q6YBn8sfzTTuWi+xNG6ZpUDG4uJzaG/Xb4CQxKhG+HO3e0hDUFW2+
TYo3uPj2Tn9vYDkoyfclpx0nOpQ7nXrjdGxdZwACCUzdD+5LdMx5xv8N4Eyy1RVc
DcKic+27lpvt1hijATRXznn9eRy0dy1hmTGKr8Wxy4OuhhWg2QKKxF45Y1BFK69Q
6K6yphW/mVSgKrCyZS4Two2sZbUy7VyZX8TFTQAaL624NdKcnq+QPMhIsbimtllB
77JmLREn7h7EKwSmB+Bimcfcoo2RD18T4Rux0tauqfxaT0IIDCnT8vnj+Z1G5Zsr
o0NBBBaVUWmEH8tEans3khFh5danSCFwB5kuSM1tMJYDYgzAINzTexCKbQtA+QlM
dmD8h0bfgu6JcVT9EZYwfscnREDCvs16ZVy7t63WAhXUU+AHQI2YhnlSxTrPb2xq
VucjLEngtYqg2eRia5FogXEKL2KrOplhLQoYHy/48k+idGVtxt3WgUFpi5hcy0tH
Cv6O8Y6PVPuOSKtaZ241R14iLkcnFZ8rfZBRDMfLkh2Jcxm6RyYdd1zoEhSx9L4g
YWecWqooyU6DyJGfuYzRcCUxEG6PXjOGmeFUqc+qV032U33siRDl+CNGzvCdIJLo
ebtdrkrOPICPxdNicQYAYv043ZODJUWgU0MSAh0fBAdtG0pdEOMxbOckxZKg47LH
p1xqd0vTz7qvEtarZBpg0b8NN2KsyzvSbmXN4G/p7ybcjUjg7PDbGc+aJ/iASdIM
a69q0zP8SJZJ0MLWz/WTKRdnNTIk7pKcu+2TrQ7I51zO3fdnpfqZ+uUcOpIQFB/J
koGOK6qys3nh63dhsjYJP3dfM3QjiRM7zTiVFQHaCmOZn++vkTXhC4FMbpzQ2DH7
dkoDcKbg9oSLoU3BHltWjAmT1hfoCdzhye3skZu+TrF9RBG0duAsGMqAVQeUP2gj
hcMx4W8qlo+68fdKegsMURKZxECv8zy16K37eBXqn0GjIEQzNecScvxpT1vMFzS1
sVcGI/KJMUiRmOaOnfpkuZVcGRwBWwoaskJt/yazvhuKsGZ1DxTiW7bxjwInU+F4
2JN3gpkKqXE/RMKcDMUDb7v5qGBTed/QEWUf0dW817uYdm/w2unfnWjdWUdRaDlE
v86YoH3ncqq+NCEPPoNFSydfob+vdlSYQfAfnJoKCJ+CmdFn81kxKj/uxPFZLVS1
00OsoY2rMK/PA85Rxf2tp39z6DggxPyW60d9Ygn/+bA/mnZr3X9bAf0Ufkec2CM9
NvYa9Da4uozNVfRhd/17ZUc7Z/XQoK7br63uQimYYQc49QJdPIPqLVANwe7gko8H
7uXmCxheAA9RmQKL1OrjRkS2NDNr94zaujsNRczd26YO6xD9Z6JeUq6Q5OLgIVwZ
RkFdjW1Scxicq55uDuC7jNENQRGIdWuFywwNHphNYceQiwPYu6mWGSHqBbhAS43a
PojNK1r3pfznD9Q8Ko7NOceh0QvJwBjXfLT9pRHr1kYQTmZsl07l5h34ehoBBD0X
9btTmrlDCdJnjWUaynqmhL4q231ibDV5FoXYSyrJAjGg1pBimZmDLPzvZfGsHd3w
dBnJhGbqP/ekGcHkJ80Kn9AgPO8oIoGXu2MwDQgi0jvH1lYoqeJz7q5xVDRF0Vqp
CJtp0AG1EgO/Mc5fDt1Z63W/M4A2vt04ejZ/KvxxCtTZZT/yFTJVy1OW0bO7exf8
MbnlDIChjxh7v8sMaX8KHKPQEWE2zBQ4WT1KsKt0L5u3OotNe+T2Y72QPeXlW11r
dChrCu5h0inYEuxeyBH/VYZn16QW+OFHR1VWz6E+wTYvhORMwstYsD2nnLnxDxDK
oBWOabj0lF4o5cK9dXRHdUgcX/9lvtCKfKi/3MLhdo2T4qi/PhZqlQwVO0AZ+bIk
7rrwfk6vZieHyjqCkLnIF1pHQL/m3T6MhNzFnPxdbmGnR/GPdoiI3vDBRu7R0sOv
kvr2rXH5PvsBLAZecoCsEpPn5Y3IPNitqdaMrwFgIngSgd+X1TSHNyCwYTus84tn
EHtlE0tI6uIM1ygFGH+wEehb8qDXXQcj+O9PaXVpFG4MoruPdlgtU8QVQm+S/U5f
pY2bnWhYa0hyVvmW6MpEbxvJPLHkveQM8UKXejYvg23wHxJ06Okz2fQZTBTDk95k
qwgcyoBBCyQ0PwnRLbfRDCzU6q/ib1Xfnj46rgFvTbWgvTBlO9ZRhOr3FwlP6y+7
psVZKiqLTwifEoFBEvj/3I5NgpszhfcO6/zWIdcbrFyYVf/cr/nXWjJE+oevdM6H
bMDy1uszLVS+sgJsyOKnCkIddu9NiyztWo73kNXYsoPypKZV3ieuvbXVZcnEN1aV
TkpGTOQFrNi5pnJoU0SmQLULzY3inkUgCbnpcLM2R2D0fqIkyBil6d1w5vgPY2Oz
EcPQSVqWmY2X7+PPig03xO164bYCMtmAsCBsTD/XPprqnjB2cFo7H8gUfIF3KCPx
ICMWw4NZLIMWPmq0iKGJTXanRjGQk3jCDT+RuL/hCAmy85GT/GXIyXG1VRgC3HHj
bkU7WYzvkTvNVcOSLHOW9m+bYrXMGv87TBj0W8Fd60GFjogKwbkGgBRE3ZDZD5rR
03y1iuU6Fuzpvrp/e21kc9SlSxN1C+tC9DdKzzJYYukFSj+7NnPVJ6f5e+DNH0DH
qZMc4pgwkFaH8KqEhkMMW0eVO85hHtLRZv30xGuA31Ze3SOqMWQzfZJ8XaBqI//t
9anVi/uH4rjkljdZymIMc4QIMq8JmlB1VN2ntlaDXsExjFGErhxSXtNqVvSfrB0b
T1DQLfBg9bg0MRbipxDQ6vsnq45Ls/RGhA0oMNyUU6HC3+B8LCjnt95A9XlS7VKs
p50Ztc8Pit5Jj7TpOcOm6V02xmAcqZcVGr0mcDP+ICS26xFPFvwFTmH2v5X1pbIH
EE0Dfg6FKSeLd1thmX3FeXLN/L6svR0mBziBr1PTHBrSnPKSLTedpzTp7ZiYyvWp
uZHGB3OIXE04HU91du0zuZelxdVyE5f1OQoKg7qRBe88T90P0IzQ5kTlNSEU9aRh
r+oc01minDjTVPu/XNbv3srtOt9UE+giLRlCXLEjkkAytIj6EtlmodxA60GhxupO
Sslc0GDokb7bMl+U2THGFmzYt6ZksDRzbtgHsaQ6wB5Am0XpGexYlvpOxJyIWw7c
LGpti0OwmZxA7m7G8CCU1ZZKwesjuiNmx73GIPOdEd4jLRfBV+/3d8BU2dR+S0pv
5SfmYwwz4Q+K4tpEoLb/4LLN5ur+Kiaq3kXb/B3DudXN+rVRv10xBg62zy5U1udr
dnDDYSrwJEigUK1d3j4uOLt5YXRk1o8b2zj7VZcjbqdyBRyID/z9ep8dWKthz0Qz
1dmBPSE49w+iceIFVjf8ZuCTtEApcoU5+SYcVUKlU60HsyGJFwCVMhuefvih0U0n
fkL3XIz9kKh+8RWKhN4CwkCekX3myg4+E9FDZWLxBW5EatBQNWs8WJO0Ur5WiqPa
QGBgo7YohrUbvKk64ir+fqvAGZZoVdVyjQkgdYIl6DMnLRu2cB2U+exczuCY3CP7
H3UjBHFoiajqGt1gMkSjVZGAhyNrfT7VkT8jp5E7r7z3rhr26gzJC+8DyHxgvJeb
AT9Pw7jSjzsSIr6vk5HNU5yLEqTc9AzLSMUzQqlGfLM1w8hAa2dz2f04wRm6n7Yz
QdNLugn7J/Difom8wRoWkHYqxEnMklaCxgSUZv/8dUVW/H1F3yKQkduNwp9r+4HZ
HUfbivY6sBqi10t+fX57oABRxP3mS70bG/4NDbmoyo39kVc1E3/1cQK1Efd9HFFp
S8BePtmniA1ng8I61MfCnr3FaV4fOAPwGzR1b4av8aCo3BYlhrxiCkbLqUpahIJ3
KznPdyi4xBQr2Pmk5GQaWhavvBihCMqiEwKR7aLqgreS+N0iXHktzkV2JSESG7Gy
qwvy6O3vLfk33JmTSQTWr3EEibjv6ri6uS706lb5u4i0vFQBgrpUx4n29+gFlcrk
H9lbGM0Q8fBKrqSy0yFm548N3myFfjP5u7IfmfW+rj4RlrCa7+Q290vd3fdsrIGP
Ok9Fu3HQ8TVuMySDg0p3xPGPI4uzfXTmVKXSzG1kPB3FVIEejqtR0oF3fuW6tYKx
+G68nXv26t09JTK3f9GSc/IFZb9uTXAOZ/123HPaA01qJ1npP8J8CksWtsPfLRxg
Yls44bEFlvkhJR4LLC2FI7/jAntSo7IYsQ5NMGqwhnGbCRWnuN+8RBWFX77hGxBy
IZf9+9FHnBoSIZCRBqrPl8UowD7XOOahJdHxCAuSS42R/OpsbI23OQDO80a3oNMr
Sv3POB4wMn3L2QnN5X0ezNwPW2VZzRWcGhn+DUZhLGs4hn/meV/UfP8aW7UGV9q6
EgfUvj8OfqxdHoRXtBHOuH/c9FHK0BUzfztU1QNL0ZuWSM4PTOqHSaCbB+uMa89A
nZUWjuTCjniDpO2E090Dz/7DrqzXLK19uSMGgbYZSUvIoJag5rH47txPwfFe6S6t
eaWh4vomyqDcJbiGtph0VA5y27k9yWzNDCZPscnZADBMPUug0aTP+DHDUn6/pN7E
CUVgxnaLWY0Z+lh3ak+jZdMfabd8/PXkXENVQGVVeGuhrT+8gEzVurIIjkr7mHg3
vtI3471r13N4O8KgQeFKCxZ7G2B7Vldpv0gDoQsOkXBjX5m95+Mi+ad++LTPHFO0
sQtT/KWzXyYZ2o7IS3HfUB72srefaJF6qatpFADK4427hh4kMhYT0tpH+zgaJF37
EjzT+UY6W6P0dEtwK32kcJ3mOxMzZPMGMm1T8YxbcY6OUQIwy3cMU5iKfal9S3aC
+X8xK+/6KHG4C/4j1WbuScOCCM+rYyuuC/xrfSbAAQmi5prYA+W0fqWHss2nOeSs
t1uI2SUCKmX7fjULPbQzRmeCeQnibBouBd6jI1sJaJx+e0aldk0nUqwxrMlsBEiJ
1BJ44grU9A6F9jSUiORJ7J/ONqPM2qpjNobzJPqTv/44ZvSvQkjznLc9odcXpBT8
q8A3vNDGWBuX54SQsvehSU+kOZnlfbAlRnzIpwxTPIL1s5S7AY0AIsJTu3OIQiIS
mdhnaNFYlelXB31wVg7XgGSJUrxtCLL9r5X0F8h4i0rmKarCZ+VgB+h3nYf0KK9D
FJe68k5LA9GhFV7hPco/DsrkH/UsxtvC7jYXlLdI2tf7Pnd04TLuBCyaIpa3tO/0
0caUfKfnpDGa4s32IRpfn85mmjroYUEfOibHBUTsl70PO0T9yxWspWtoDYtxzS2Q
PNIM32jLAekqd1y3MWcGdI2kYnMdxiErU2KBwvbUSeFtBg/IfKVU8urQzPepDW9o
N9AGUdfb57Oxcj4iHpdWIazQ6xxO5prdPcFELe/+TMEDKLVlRHFDGuOjPk+bASRT
qmjzZ2HggB1+HKneYsqUCaBZMA2J4QXvlt5qjsajKqrw5Ds5TUaLLRlUCPSsgiYI
q1jgqsfW6KSzYvmrgEB+S4A3CRFA2QR9neRTcPBpFjBPdndSWL0lFDSzw/h+WjDK
u9/W520uJn2XG43apB3KONeSI5D8wV0TNEEDgwMIz9ooXXcowIn9YewnWpwGURnA
VX28NuGsVXDsMDG0w9Oz+tZBFGtSCX+dkWbvzDPxyRFND6ho/lL2XDyhCNXLoqpY
kKdClBfHprlugVbfiISBx1JFpv3xruZ1ocp2Yigaow67nD8C3roRoM3FaT1/vcdR
zVeIULMsS3X8THI6IbeWXPrBiedeh24TH9om1sk2LXdBJUGvInCqTAAcUtKkjksi
JIa0ufPNb+y9CaYqVrAEz4r4+OvEUfrUnb85iQLhaOlJMJisqUwRHxp5RJZR7C9o
/1N+PQGRMBapMNVpncjpqzr64kxKV/VzxvAR6zno0kCb7IJw2AfZ27v0asxaEsBy
teHDA4qFWLzTUBwcCzQTORoHNoafGLJMoYecnt9CwNqm4G1/uJh95VI2i7YO/y/y
f5JuNDln5dNW/+z3p8VFmMMJIastFp6lyavL7lQY9wntxDZ0Sf8Nuz6rOL8NqQZa
BHXqxW2Tkj8nSwftcuBLF6kQD19QWdIvczXxpvb4AND5eiUHRdgnOsYFbtk6G84Z
HJZ974U4/dpBHHg2ZvT7+DyQgcDId0E/wy3j/pEgl0TtrrUQ0p95/U2vxjC6HaIX
z5aGXm/q7oqwus4LJvviPMqCHdSyVKowh/qjNeojYy1HezBIcoCH0E28VkvNcRU0
0dn9x5poUXF3PuhBnlQWMjhi8TrBr/ha3SZdc+0/DZl831+beqU8bWZE6hINGRKf
FPy3h6guZ2ffeCHhxG9NXsS4RCUtTTo/tKvN9/zoE48sGEik23vEuNgnGadK09xy
UnJWk9ir7aYJHA+FSlLyk4EvuwAyexx1AljiGCeQ1NNt3to/reKD5b2ltRwXyyft
9QGNdVSV7kgnFtt1kjlYC7eh+qg9YJ8JRmmkbPPmRX1mqSPyj1621cKA8AZohjsU
ggOZn6mZuxk1bDUuZ/xn88k0+HOM2dXs8+1RfdGdayjkXg8PBuIIvlC5MgmXRREr
SjaKXWec4AHlrrF93P5PQV9NsNMbD0Bfol4PPDgJNRrcnTsUx959dyrrK8DBVILZ
06/tbQAmfdh7ArmTKKG/cQjfuzPvGqjDvQG+fa0h9MxDkJVJiwxGZSuecz4idFKF
z30Ha4raLFITuZ/Mb8hS1kCO/ak+ywxiL5Mygj+lSiIzKK1EJJySVb9KlzLgwYUt
sNaJcOmMQ0xXfE9s8Shjf0MwFRP7ZWJ+hUrhZPzGmleabh4E23Bf3YgQslp0RAq3
+OSndZB8daKmqrB0RgSMGrRS3p1lKpoLbhjubfVgBdT9xYnNUfj1lB2PP0zf++Nh
gYKtxB9UTCe6pFMnO6Ulg5OYKTcYn4xio8OFDTJJRRSis5wzdsZ5Q+MDgq4P/i1t
9Q4w7CCz3dKCiAAPSv7d+Er3vNtJhvxqVxgSye2Zy125zEIZaPybAwGrzG3ZmQag
XH71C/5EluvPYLlAtYlJKn6Lo/w2+3RsXY7sm3toXm8B6uEM7v78S4qCZMHjQs8A
+9pBICYppJDsbPgWFqAbqBom9c1Osu3A+83GEWKhQk0b9VXod8jClR0Ip5N1qCnx
p4AEF0ums2VUh8NaD5VZ+dOuUVf2FuouWHoiZf0Jri0Hwqtgjep64w1MXeO15keh
RTLYWH2C5N/xInp9iSwBvcTKUEEJASZI+KA67OwACB60VsYNGdDe+3b//BmscMCJ
OCgeyA971IWDgawCCdDjMvcYqoGnR43PmYAzanKBIoFnZU4YXht7S/b9MwflwrwB
uO0H2z9lHlJ7k02ow/419Iks2p15U4x2t9C81S06V/zWXtM97PxxXk5W43IUkJIK
G4iZd97oKGwLMP9B4M/U20jpaJkJY44i12OutimHCEXhYvHTA/dJ8Py0wes09Kz1
GCUD98pnyA7AoRbcxASo6e4Pj1QvS3gC3N93TmxHaGi+juQtyz1LxoI5w/SibZC8
ijJWP9l/YXT/BXaY0gAvFn5tiJ9DFsH8gRfGiSl0vvl/YZB22byrSEejR81HdjUB
LsXo6FRyiz5n1uFE7t0UHPksZ3+edpcg39eM1HfPWLfdfVHObFOxappa6eOmuTSv
Kxty1Mgg7l3nvAAo0E+TvpV5eFZCMXUpfCRozn6oINz7Xlyq62ZDAlf2OnSrXe7+
TQ+Sz3jVXooWDw2oVDHwGKgBuP7P58IbSI5g3i3ul5AOW+DqKXW2Km8rNFgrMSSv
+i1O+5L5PKal0dDzE2GAqtPHR20/DPkLT1koFrYQBI3rSCGhwfGzBmGUBiKnRwZP
n4+K2OBDPc9/S6yo9hCHDrEJvqv/OwHKlALvM1WLopHPmAYW7OGFw2q4l8to56pa
PRR8QMZcHx9vp0+u7RJAp2mFM9UrvOGFb8uGaLqr74KvRpVgRwWXH6earbxI/QMd
bFx0C+YkPMylcyIVmDHuaiQgcq7Be0BBKJmAgQqHRanr/6//Fte6WuD+0IVILIJQ
EMZRAhoIQk2GDcxuX/msGUDD1DQVETpjTubfN0CsZ2CtgI7y4yucp7GAMx2cEZpv
Yy9y/LhNdWna76r3zrl3BAwqZQ6L+kkdAnqo79KQWxLNs0p4LhTd6lIei8HoL93i
l+v/d8HWJxMfgtMzbVX84Zj0opcreea32z6xKZKgQLYd44crH4YN914RrTmMrfr+
WROMWZfpAhomimGUbi9J+268LtJoDzPSaTaWGLlsoZNrVXJ8QQQLuQwy83Klg0xk
nwjeeW2tUoYFkyRt4RMsBdQPzbLnIQ2UROMDUl8iUSWI98Et95QVWk2yDK/Gndki
hSdYNBHMlviTITols9hP9Vfe/dV2K/UOonx4io04J7T164Allq1KwwILP6lXVH4a
FYTLeQX+aVsA7nalyCV2W63Z/fwLpu1EkN0RP7ZknjwAeRPk9l0F+AYfdCcCIbwV
d3CcSMXcGinc3vK/rWXSkoaYweDFAs+4J0eh2KFcmJl2ySup6s2Vbg2AFEGJUNdN
N4FY4Um36zc2Lgu+nA9CddtByDek4IiCcPcHv6NxjQET8bhKDR7KDKfx0sol2UvI
lVGxNMFOnq0O1gRXwHdS788HW2CSyh8DgeQq518nQi6RkBvWUmxp7F+MOochpiFK
TB5xr4rck9xg6mbGdjcyykN55DwYAU3Nxih+jsld2D9elURJawxi3Sl2ivpz4950
c8AJ7mOoSmXABX0RscpuqrulCmYJm0SQvxlIcyyJnfxFwmUgdiAwuGk48Xl3etwD
9+/WZd7aXFDbHyCg3eu2X2nb3s4OurDXINP6Xvn9HcuvIwGoHue7ZUFuVhvvBooy
SNHSJVy3HIEg6rvyl00ezZd/XGHQj5p7ait9Cryrr2cqpGgCNBj7BCiFbe+V1UWm
8QCwS/jDL9ODkIO9QVrFpcKtGywEABBx9dVVdtwMEBykAHJfmxnPguH3h7joee6C
2yFQuy1QNe12R4Px9T9RVPkgvicnIl7sgie4aX3K2NOiQhiotv/zVZstlFPvPQ3R
rO7aj2Db3BNMJR2TR8JPOXfV6XdjleV5TbRIslRZPFLVKkOwp5/rNo4mFyuuLT8L
INzEuBtC0e4P6w7ouHuz8Zj2Ygc+GThaAfJ5uGE6FHzdyG5WMOsWx/WA7Y4ZpmOO
ypatz7TOLqGIeAYxb8V0LDYbpLpF00YMUO0TBb7YYx1KJR7uum24xmsy/u9iLNSn
RdHVOXMqNL7SyivBekN2vSVHe9KCfQA2U4DzE31uKXctoQWS2UsHDqWErs9LTcXN
sdgAzwJZwzCXW8wwFr6hSTi0hFMxTe1bp6MhTZpgEfNs9ir9lyGObc8ReMYLTqlF
kdpNEguHTP6riy/pI4TZ6w4L22LkgVHZQUoiK4kLsm+zJnIb20Xx5f67nabyneMM
HrQIYyuVZ9L5GegAFcvMjTRq4cjfwLEYAOMFW0KG634m7ZVESz4TcBkWJ7emInSN
qf6lqbr6JxqRhigHI0lZvaoYtOv7QRcE6AqIhRkOdfSh7PoFA+s1OPpUNtSjQwG4
uNZXj2UNryoo9Z74J18xcOVMuLejtBYtcPMuQ9qYpR2ApNaa8oE51Vza+8cb0kDe
Dy621zq9tiPGSpQItBY7iWKGUPBYxiMP6UlatmPpaTSIpHYxUB8URKUEdb1ZrIUl
awbiirHKm04znFX0HJhM9JB1NFkN7m7qY0SZ20iUhGQ0Aw101pbkm3KKXXuHiSBZ
ttAUVUcfqlM5cBB1bQswb7lkfZqxyvPeroPQPcqHSkCedAxUpN7cFqzc7g9W/vmp
h4CJcOxheMmdl/IY25FqA3Bl7A+fXHKxjAUBJMEFIxR8ZRfgFhcBnlb3outnq3r+
VBWcF+B7yc6QPSYp0MvfhkEhxib8NH8DEjQMkoxlfSXZ/aJaTDoJt9P+iuA9alJa
MCwkEj0lyH3syPFl2MAPIXgSXpR42OZSWbfvM2Rzj65D1EOxE7qgZ7/Ke4Kz13qN
NHgk9wrjINbysqsVmZWHxgeD+5wOtisk0H3GVWhldCJcvvxVaI0nWQr06aj1bvuk
gc3Xdfr5yJ4LEabCUugMGtAkl9NK1/7DUL1100gBUBA7XwgYOdSmLhTHQBNzOC0X
hzvSMvNUuSlolu9zB46gg9yisnNAqa9kRVf4x7fNxRkWg91YBLltG3t1rYk8+UFd
dPeszUS/dC6WbRULi6WENxyZn9XG+w8gFPsfqlhl9TMjzZZhJLQAuhR+/5n1TM9b
oN5Mn36TDuxgsrW8iCEriLBwbrU7cp/55+ojoDF6zGY+eHDE9ro6ib98qM9f0xkZ
fYCdImI8HDGcQy+YFlKdrGLXeVQy/6ZOm24yN8P18pBz88BKpj99mPIEbuzfNmPJ
JGPhaQYXGY7JldhdVXmvaQH6T03S4jBV7bHly18jiRKI/fahs19CVK9yD9RWvZop
yOfgbnrEbvyK3JXrNUfxcYjBqDaUiRcswwhfLG50cnyY3+/BCj025RaphUkQElMy
l22ziD3edzZnJ4GV5imYtp4uJJJ4CDE35ycD5PaVkkO4VOHXIRLebVjK00KSBv4J
4sCHTHPZfe1sELWXTA9IofqOZfz5ohGQXdG3/SzzsEyQe4bdf8hO2xs4DfHm9yFx
onPa6Mw2FU65N5URvajMn2FzVSmYI79GtVGpwEK1WVefpN4IRgeEfpi9NcQQkedG
2z8/JGzUpOCzyEyx5eApgxtqqOhSbJCPgYNW9J50A+tVACZUIvHG3uqT6z1yxh35
RTBqf7UcmZ62Q+QHWJ3sVD0/BxnXZsCxgq8CHs1Seib/dIkNh8j6ms8iQHAKLXAI
YN1vtiwjxw8xqMu9wpnwBvCtZlhlkvnOq0p/UNfRwz0b3tisu9rh+AU7oOs+hsJx
FkZk9f0y9CmoRsTAvsgY+/FOl7GVyBt1ahKTwObyhHFAIQkqGCFoEcXQGu1yN8ew
ZGYUH0vcHwusiEhuvG4ZajuxZJ/1LDX9mL89hYTmTguphDrdmxQkqE8Smhe69v5w
HAcr3/5bvQPO4eqk3ob58HUeJdJRmy1mpJ7LU8hpy5Mz3bGEpqJkG192tk6WDUQo
Y2mpScfQSCnROLkK+RZwT784ca44jKcNR5U2FTq16O3Y5Yd5eW3P4HOVdxMmYD0S
+LqD+1n/8SZ0Eii/T6nIpye/2b9L0X9K7CB9dGT44C9PQCDtoGitcm0xB4vhSZxo
ZzT+fVpUDvGUzy4C6pDcdRAWDdYbz/tAWqVfUpliTvUSzQVvdWY6V6Stu0GhG7s+
cqcBxccyCZaXzgFcQGMlsqr3iLUFiiyPj/e4BU04oGD2mYzSiINmE1e31+YBJUsm
hS50O0cfZE8BSDXDqYdFpMXh4kp8vRHfBjuRmNjlQOsA9D8TshXF5qTRZun0flOj
vb8zbzCSz7RRfGqUL7YAY6vLQcoqoSqCfx848txi2wgNfi9MKXPDMVINUBU2aAyd
hTaokB/5NUuvrYoFZpQ1QZfEOquRlc1SlKvXHWMLu715lXa+JdBNjfCfj+n9+Vpn
Ba1baZrmgkgNqJQI3B/Mamtel6fcA0I2prX41lq0rYr1/YMpK2tL6Ww28zHfmRFV
v9FK2y7zXFIwFVNOlfil4srUDln6cvhqNzMsmmGu6V9yo2lRQ5YSA3LcThrfHkdN
MfvILDjWmGBxmh+ozLtMSnr3qjqhk+3M4/K1XYqcNAvn182dxokL7p7TDEM8njK3
ljEbR7AO8l5jhfd/8uA+qWHncKNU/9PpBMucpv88rJ+d3rbR/VqyAi2vpxN5AZHa
6MoLRENN7L6ezKPLOkbfNWpBCmuPJ8aDn07O1UUzrN2TEbSwoT4j6Ey+7y4MuHuM
AiWVjgvx2IhB/ZqETGupJyQ1ud9gpNahEKYUpytM/ozRxrE0wxco7X8Ny2gFsd3r
kobaxyuVmUkNgpFOkrztvry01fJ0IlPUEFIeTHMQYGPinYbomc+dY9T/88UHczUN
vV1KQ0vNp3zzzwOMRXclHhFx94lY9cgDIS7sQs3n0qiV11/zK+KX4fJutbmnHuEM
3SY/94PhlL+ig38Jd8IciKA1sNegSGj4/IDnno0cXpOW/1gCi4IA1B3iJzdr0uJq
5VaR9g9vsZGpVfPoeK2sBFxfyha1QV9SjtEisV2200FnvhktcrdoNSK86JdczTtW
CQQwSBtwwIdtk50cZz8/xRQ2iMNlnb9ugZHyN9965PfhRS1ajuPp7jN4axmMvZzH
wdC7527uYAsv3D++X+rRnEyK62vc7Bdj9KaDEzq8x3/7/1X+6ck67TPburBLKJSc
p4APVa5Q8iTT6xBPcxtXSskJUgM81BtYxzrF9hIrKg0Gd6tsoKdxV7AVL+N9H5/n
sdclZI6CJaZP1/4Z5jgoovs1eZ3yuvMadawHNuQ9qQJ0zl206+eWZoDUSHVFKkPc
W9tYnOAaUnI9sylYS/FKjm6sQJI8TRio6kKrbmlnpZL74O9mpVN+ZcxHgz3fwROf
NWZB3tSymj0V/i2AlPca/YaAvStnxIXwrSijrbxqFzZLwpqm9cMaJ6Gf8cJwAVNW
sUzsHnibXBIxMzX0HhrVMtFL5/FFqK9tSnFkM4xCMXgNTXWfQ9iVq0Bz/PtRaAq3
GQSQsAskB1Zdj9V4Lc1pPOwyqkTn9nwUglcFmJF4AZLMJfmlG04KtJyUvU8nuWOe
vMxsViu54SoZRu2R2G7xc/dsTKZUgBDSgEPb8oAedE95vyESp4x7uMpcSe5Pz8Ff
EjUQ5UsqcFFYCsutuUMkQdSdsNP249SoO9GEQzfiIq+XwdOZzglZf20HJmYtjfRy
JjMo6ruBA4ba9If8OiJBf1x0z6pFi4LyhRdW6E+V+MKEa8r4/m0r1CiIsN5943EV
wUbXPTMwgF5HpNv4WOTFW4Eaeur7Xq3LML+y6SLuECNxiH/Hj6xn2ygiru/khh0X
YQPmNHLb3dcEjq4cevBwyvzLCqbZmOmIkBzeDenmT6TuOARfUQWFXdiBfzyk3Rkn
UBjKIPrrGH86NdDDs6hARmnSW7kT52/gvsUE5DSBwykoakuUvYMrtwhFsoF/yMQB
y/XXPCDCSWn3YaHKuvLUgNdIP1bvb3xk699WGFnXaCA+68u5BnpbcVRIikhYC5DJ
dvvgkiIUXnOSRaua1ZgFUXnIyz8nAnw4KhKLlP8bWebBytxnpF8O0il65A/U8eHX
F3aSqPS6OdLQbnjGTsOxBpraU+utsEGjQY4v/nZr+OCs94/KS+1X46m+xUizDXBs
on7pVY/771kXbhsxNgHgi6EUbyw9aqdh0yQpepSP/tL3oYIdG8C4SinsYcUYExfW
ky8aR4kRKJMNa0bz6QyLSzA9KDC14WlElyNXJz8EpX3jx74h6v2v6YHxKuftdR7Z
XbBgCGDxt8Dawk64+chqmi8xB9uUQzxEg/GNY47Oi1vcoccl88gj5TZ3eWcUnuBx
3hHCAXB/0cRxTYUgVtwQZ8VIeSrpDSeH+XabqeAmcxsMF6YQ1ab7B9DgfxOcPSVI
Ima/fGpG4B845oBRPquh/lfkoLZSioT+mFgdjN8/UkRcYj3i91kTwFRyJdSVFR6c
orr5bPiOwxFUVpAVeg/MK+SiyIcV0/loBo8Cn/jvDIPK6Y+hv4eDZC0j/yJxjdTR
sKS/oErP9wbpENEDRQhLYO+I5J7ikg9SA71UDk8Lqm6Swzc2tAR9GJAowz3oAFy6
3xdOFZDIlk9ChjnAbEmkc5lC2O9OLr4R/oinnsyJodq6p5pFuZcQrkjfcBiSFc9E
h2w5TptHDsU7h+j7KPrt6F94SSh2yKe2wVDsOadFHlXGenGW7sLEqlPdOWqJR20H
OyFBR+HYL45zUYhIiqWpIBDDjHC5XH+rO7EVeyfag2aoiWs7j0NxX0dhPIHC4jQm
KH5wfcVGpfkGSn2JfbQbyzV5+RoxrL1UogyrlNatNscP3X0WvJQVySi17lT0dNVq
20GxC826f7tYz2cvNb9orVXPIm0q+kYWBJU7Ep5fW8MZ6px8uHxfpFKroMFHCK7I
ouCbddgpV61bHhJvJkTKoekjHFvoVu13SjuqCr/KQsjGp/XDfH8tJgvRZQY9ixft
Bsh1U3xFjBDhI46Tf0KvLKG9+y2SHCqUgfOYVbrp6Dw6yvPNYVBcfuOxth6bOJGF
s9KpGN4lc4lYas8ymptYo3fLYsj/DA23wdQKRzke/akNJssCv9vz690QSXsDR/Vd
eq0Idv9FTSBkp2BqqYlVuKbFRH7nANg2QJMosWv5fHoNaU0TNkZCHRK99u746m6S
5ITtpngsFxqs3NzQG81wMoaWgR2JjBViwu5n7VmjbNDMXpFFTmNPdk+6VGD/Petj
S9B6qgQ4/FBb9OkcMX2cDBjOmAZjbiLgBtlcRLxDe0WY/2Udhg5lTwCHWB+pr2Vq
z+GEE6KFT04fszSgt5JCnu2jJEOeVfERpAjXnEf8gUgDP/m0f8IqXkHspjOEAM48
CIWNfCNdF1ZFaIBtpkiIo8yPzmnK0e/+DEQZLaW7H8fN3LQV47gVzGoEy+BG7sSi
qD91OvfVJYwsEWevS9ef1dkXQb9XPAAFUF+ZK5tV982TUoXMN5E9p3ywJSTkh1/f
7oBtkEsvMs5smA43IxpZqOvxYTDlbKfMfPspkl3dWzoU7Ate4qZDUa8tmSoFUaYE
oRlLf7liMZktm+zwAsqwUyOyfuPdTL+NG5JAx8FHOZbCRZnDsvQfL93gDv8g3X5o
k31SFVV6lzgPkhocebMK3xriiraTc2/8EQgB6YT6jWYSz2udu2/NqnRFTC81sxWp
3cq4pRhe/gEZI7AzmraGQytfD5HREvuhqYwN7pjljHamSKAMSCclZPhjWMKMvGAe
fkJbVAtG8pR++UYI2MAW0AKYqDi2THtl2gI9n6pz5YEZ1sUvrsT82WMRaW3BW7oU
r/ZrW2Ef/2ofkh7ilTtsm1sNO+lkAY19cMA6z/UtB9WLHx3S21hxEXYXhqfe/0AL
YbzazQpAKrqna2Z6bwrniH94Q0IQ0FOF6jrj6a6ic2T/sBA13TgfQk/23pe28DNI
1uIkR3N9dDZAg51bYieLK5cs9SR1V3qshyqW2tPATKIie4vDuzRkoXdab2vAdPQE
wpBDi1k1K5bl1L17hh47Xp2eka8UT7V8ClY4wtGUWzZD7k112X67ni8rT/DfZBPT
dfA5Iv83H0kYmSAF9XqEi204ySiTbBazwWfQJPlqBIeYeHFQqEIdzZHl5tCkq2n3
j6KzVxiH5JJPGwxhjvxqG865MsZ84apw8yP5fhA/PyQ6oKt3kYGXP+3EchcVJHvs
hCGupd5kkDDuYZGkB7e5m37AtzeWfzUIXzsOu4sdboP64hJiH2xweY8K6wo3Ug86
IXrZFlFD9HD2ZDXLM2zYhp1m+YgalTEs96Qv44ha/AAubG11PrNY/93ecjbteCbQ
7GGNsIwnrSqizAfxkrX+7vBmm1zqFLXLkehiOUbh2FmnaM5fpEag6CMFvvy34cgv
KGCGQW4CrgrWfCunVC5RWoiGfh0eUbrQlYTIZYBvJaOr5rZOhe1iYlUEHgibLedm
vORyGaJx8KnLPiqBc1n+qBzrjGFxnc1+Wkkma4ioWbVeUSs1Os4BYeNnMppSXVlh
ON9mXEkIyctpNfXpVBNQmfSOwvuGYb3hVH26mbZODlc2MZmo9J3Odvfb66O9doID
qm071kh/cgplNckyU7N5fqxQ3kMxn342tASKRW7HqLoclyyzqd4LJP12iH2izdCt
oLuDdIUEP1MDskNyQRnXaEbF+XEHWfBnsTwFQGFhbqF/ra1+mmuSKb5cqdaqRYlR
mJehRSMvbGTaB4dVKUeRQxRRoLu3YSexZ915dXkQenXcivCpNW7z2LX6DbNufAPa
qr2FcdcfQOJ9NxdS2PhUd/eMXHSVhcd9xrvs8kuyWnV8H//5pX3GutUWmkdQwjxi
18BCQpzchbH+9eVxcwCjlXc1JdO3wx2CqCOl2R1FO9w50xHXsc1E2cdJ/iOfC5bX
g29MkJ1w3eHeKI+ymlmIYYha8JvfddUBZj7RP8iJ2hxx1HXbx/fS1Zt2KVjnEnh0
UQh6MSQYoxaeP0VlyTLvqfXdNn3KBO5pqXU/wXLMh53X+zsVWDCdcfIn89XWcihi
zavqPzAySxwt+Ks6qJUKkOpeADI7vOnpF9r/5prm/GlHYjQHKFdrhRWiFEUTiFNv
lNA+nnFmtWGX8MTCa3b3sl47j+mC8pucFRE76FZjTRNJSWZm8sgZuJydrHxupxpO
xB9hflVYcrBZtyI5eHABgUWE5ZRyaQvCM+sgB4xLEI6IrUs3kXb8/lOyVdVZQdzH
sLfeHyvFLzbF6pJFZBhGjw78mI5QHLhaYRE6Mw3J6lJDx8UaxjwjYwkiRzB9sMeD
/BNp5tNXJud0NCiu0OeH7Nb7YKSCvsBlt7ww8jjzPSkBs+VC2U9L9Ap8RLGfdMcr
SD6lpPmECNM7wVUsGEhzR6MM/j9WhlvVOTTDJHSWYHW7G1eRTX5XklOczX8IIaLX
d3s5bs/71AQx4e4psYn+OLuYPgexT8jURoy/Ak0tCMs5z0DINRUAPz4ovlUFWsYn
HcxXgKxp8x89DkgceP3V2Q4oXByfJbOwJ3eIqkhneIXsR/0gRX6ugb90rxm2aGzV
1eRsyL7ZZRrVXMJsOWa2NJX8PkRY8G0OWh/opmctq6LTjnT+XT4JbJLu+n/y+nI3
3PHX5c6JVL1RqhpJWTKKhxltbOdqppSyizjMQzZ+TYnmWoKmKpfb8iYsqHAd2Pol
rm3J9Y6OnnkjGtmpUjPr5LE0dRONPIo8UM9ze4p1epiXKRb4bqpf9bD5VPYm53qJ
tRrRJrH0l0CqDR5Ifoq3D3AtBFNPzJXDJSyXcaBwYUHkYZUsbTao0XbqF1lNeIpX
uuyaASspVfsQdUMPGjd8G01ab2lS0vV09/+is+BIYYIj/R9S7uPNeiK2rSbTIPxl
s7BWi5m3AbL9btAgPad9h5MQI9lbv1xtPP84Lskuy4H6dDD/PS7ynhyzsJi6FQM3
qoJq+RhkAs0QatMYForYVxmbQ4pJzAOLrNP704yjTKWiZKCHebWJfolzzfj4V0La
b7XbwDTYGQ7dgYq/YBdic5/c8oRHJWxLbRuqoDh00Hw3z1spWyVmVYb7Xnx+L85A
xK37DObfA4nRlPSW7SWr7QRDoBFyx2YbNWAHhKjfu7v0qkksHWvjV01VXUOV8/a+
C4cIAu2DhtURYjUHp6KgxkAe1KV1S8Oqdi7WfT29Zi/4B9W8PqRB/QodDXVeTHDi
tT1f5bHrA5nm9qckpcK0sOmRHJI4EdSgD0iBofPMhikzADnQOictSdpKVSDb4FGF
w4YUe/DkNJnMFdoDWV76Hix/9fiq7uihIbAz/sHKySJc9noF2cMfMC+S5Jlp9s9i
CxESzT2nlUFmdSDvCSAnclqsz9ZmVCh91Jyrx7q70pLb1JNowraanO+dddyECMem
bafA1ht9MDA96YnRjrSH8uQAd4HMdIHDXDpV+J1I6CDwXnc/WHtu/Mwsdc1ULf5r
NgGJLcBVhG0vVYAX2Q2wlYNX5X3fSlZbwVOu4r71VxTpWHuMh0+bLNunyiu8RA/m
i292RhFMISjd2Ues0t2/TYPmYWxow1AU7ejepY+eo69f/v1k8JysHIKnMTxpwxA6
faw9qn1eTKXfeYl1530dgoAaUl7s4yX2cOrQaqNMV3xMQOLItsWUAi3kCJYqGmMO
zeZ59KJpxNA4sGgshIHk4s6VI70rPcCtRBwhp2XvHoZ7+kKiwk6ngt5sRDKVuT3n
dgppJg7EVMvPbdVQi0+OyZXYqQd80JqNqj5gkVTCHztH55y4O0da4IazutGawqhe
eY3bAF3/qEjNbnrYmWFoVKW2CmBzolFypXuJ3fVL/eiCFo+n8u4ez8sUIXmgOUH3
h/O/aiS0TznZmI4N+TWtxBAgQtJRgJR0okZsdWIKaRzdeFpVPOx8/gwkQYqqEMu5
GUEpAPZbjvmzx2YD6h2LKyLrBLd/UCo0w5r/86nKAA4kpqiph49XpKENoWRcolKl
sv3XX5mDn0yZoOxY8AtcMN7ciyyTJBiaAyuMId7qqjUdpbT2yXQv/JXBYFyuR1IP
zbM4UfaVxm28yfd7aNYpEQJ6g0+m1qgfIvalb6FNqGw3FmkTVtyYRZ27kyBE0km7
Qv6+j40gKO+MNxd5ZBQ7hMZ4VfOorQDcSr6rOE5mVt+QAmRWAeWp79xu5Z6RE6JI
/wMbCCo+dA5Oo4Dr7r3MZibAQOlobf+bL8CjgyQbyBBO91ON+93zmwug3VV9Ag6g
rvN4M8Vq/8tlO9Y3p3UV33uvZy12yGbdCSJLeJFacbDGq3AgOiRlFg5Cvweb3z3K
ljzogJHtmZq62GT5Q2nA0Jt5P+QvZ2HWdlop6iYYZp1Ti1nnIifdOLucv4D15VPq
87urMRROdPqvDuk3uO9BkgjcrxlUiiVMII/AFbuHop2ysR1DlvXOFvbvs8pxd4gD
8Nyenx7m5pkuMnpY/d1La04xqb//CkMTI8oUNnzTQVaSVdxE2zfapQJQJkPi64Kq
lOjgwmvvgVj9ROVyuBY07MB7UM4qdT7npySy2psl8lLdjXC8yOEyPA+Gs/3TaGDE
h3eOEgbVc4jsWQU9Yxb2wafar7+C+vrpTwmnzo//D84bux+MVeVNt8uWG51FHyND
wfm66I0+Z/ub/oJrDXL1b5nKuWhVvBuy1khmpAIqraBLcCtVtmxEhGy6SzTswGlr
MYJRH+kJBu8qTtJHc8Q0D9VAPrRAQ/M4gx5Z3InYlwPpQ1fvlEytuYaXfhcz+xq5
6Py0Zpr/+a1avTcSx5cM5IDr8G3BiYCbR3GgYsCJWmgyX6IpeNd+0eMC4mwiDb+R
WVubDApZbw914/LhEj/5oBDwmil3CGCkbTlEgX7yhEcoO58FODoAyGHViDYYK0fq
V/E22R0Ja7CvzLXWrIlRxqlfQ32i6d2B3c7ns8RlvgrodP6zSxrcBEMyBF4If4wa
fcSUaQnzmQzSyNli+H6P3+PZ1d1b2g+3imE9rp0gUFKNIy4Cimut2COndNbClQ5Z
Y5tChQW+iHDHDN6pGNf3E4UuyTslLtGbCPoelMrSlD/Vdj6wi7gZWbye0EfT0vSj
63BsETefnrRcQh5O+W7HuIudYsI/xTB5p8iKweAjh+W6tWpcs2qJchjkdYHIdaPb
zqZNQApzzww3AKOAgk29ukfzI6ZJAa2x86bkwZoGu8b/tmpazBFxkirzmilefJRe
8nVIU6cc4Ku3ifriu5gDzbkpCFekG9Wpi7XQnLiqXUuPqkpkmXxbleIBkHH3Hf27
Iyg8inEHjykFXnCI/9RcNLGskXzTOeecyiomysOC/Kj+6/hKcQKenLw+LDXiXfSw
jzYCFDDnKdr9Pj5op83nEsYROGbP9HzHYo0HaRx6TbxwIXeGq+2goZ0MqOBKjvnV
IMcS4NPvqGw9oVweil3HnkYmseAjBBcEpoOljJJSimLI8SJlHp74kIafG/RjXE7o
/iDJVL1j62rFWstQjppM7DMoUAQ9XWCsE5b6Wcjb6Fv9QKEyP2Kd68ig1cLaQO2c
yU2MaZROTmGGkkP1vzT0N9p2vXFpXd+cIa3xAvSLMdnmNtdMdkgeoIMrTp59PClP
NUGrAiS6nxgvfS+abjnFH/5YDq5wuyizAQ2CCJJuVWbuWMc5im22aseL1CPAvDFl
PA1zYKdWBtCnewKr1467hwShlS7iASFt84YCKnAiZr6kyuMKvtRK1N4HAQS51dCO
2flP4Xekbm5QbTwAcqrmfPCQDE3szCoZXQ6ceaZ2O2LYzZ/t7bf5cZN9gbFbQBTt
bTDvNFCVdjbbfFAc9H+oa5gtA9R4djoMTUO4Td1WqQxYPUHvBY6mJ+md2FvFtDuT
2Ciexo9d08Xdd+K+B9SLYVkURMyiOq2sXrDW9/mWGygtpO4N2C7/g0vBpEJ7FGjf
USGjX02ees4HHT3GzWE28huSxcTyahu3fLELiUH06zvBcgQ51DuF2//2ZGjikhQV
2+9stjW745pSAhp6djUSMrNwiYq06T6rn8T0pQ0yxD0qxkjMEZ/CqZanMMDRy/f4
N3c3Qpw+S2YlCqJACARnOKzuzZmegAUWfdVi6TCVVJiiFYgv7tZT08Wz5ZKSJdJD
23c089RGmAeH1h4o2pT7ByFoZ19EQjBfzxLzXLpDA0S2nzBoQ8s0LJR7GmkFtwda
Je5Kvvo5HJbTumvcVlsd3LnIleNaK5qFVyC0rGP3xnX6CEBfMcO23J2C2l9Z4MVv
LVCsgQ+Y6BAY1fYampBzdEVt4PMrmbx5+SOMpMFLMZdlyqjywWeDHCR8d3jpbeyB
a2YQ7NGnEJGpeUek7GMblj9FkgagOIdmkSq0ErGGszLkJWOq6/2+2zzbO0EjXjCM
gWQkb5Km1MYluOn91dFlAxWmBrXIiaQ8qj7Pgaa20i39xSIwZ9aTHxlgtYx/2qgx
hRXUOoEkLMiYqyJmcpU9d0WuYcTNyzS6uRcj/rBPJzRLFrR03NMZOaUMSinQzV+a
gZbtl/y3deP8v/ZVg9fiYAwHqsA/mOSgCXXbxH9Hoq1YgfhkMUFlTVw/+t0UwrP4
JgYDHvgFd63t06h9ZgoWDt50qtsoFMVy6OELCuwH0sZQ9JwUw4qTQvD+U/0gM59h
RPslUPpgygIUKL/ZYc/uhhAuIUuRKknlTTmmMW0NTXOfwnHCmmI9LPORx2wObtDD
rNYW/mTle7TaIF6+IY96LviRn4ImJ8101P04Cu0zTI9Gv6H68P22CnNxieNenQ7O
hJ3dwmLjGAMym43fpv8yaEs5+nOt3x4La8NiEH16iLiQbpsHgQZqgOg1GFEvf9JO
T4+jeRhM2p8soAmSWHtPSXIG8zhIKyDTVbKDljx6L3LEZjc7ngiZIUtfg3ZHw2fg
soyixmxDkiZaPPlIhaHgwfIteVU7i1aWWIMXE3ihEj+b/hjdKKTw849crBh/x8PS
et5MsmEmPLR6QqP0v48XEONOXV+qDaTVHJrD5Wr+SXaics0end6LoITwlk5uKslI
4fyMLhhN6ThUbSRB4idxWISfutoOhDz7AEaWhm7x/XsqRj0kwtfmzdM+wKTEhRUA
a5kS5KeCziptpJEmyuBwKoI/eH7XztbnW7pIiVcGGnKih8v3xWreXZeRbhHuuFoz
/aRFjWgYsXFYZasZQRLWeIa8YWw73PyzePnbFvvP7m7fTAyTbzLNuOtrWfzyM5Nr
TcFbtFMXEPyFriN/85WH3GSytwgOmg7w2MXPSPAzrDm/cpYqCXk4Utelu6EBOxQc
Bi3xkB5UleinAZO9mGOgC1L4X+RCQ5M+j9HdL3Pc5M57lOAbGipdS/S9RSGStYLK
AAegTsRNjhdYWOr3BKBQOkoXEf0f1IBwEt56NvQdliZlYHJZCEkHFs5IsRRkzdcE
JSSMkjlhPifWTSoBMuVcghCFljeWzxLQrJ3pBitbw22Itb1CfDdN2lSqZliO/gd9
t1h59gk67p6JZ3vLj5yJ5eFRu3iDxm/9Avq4GZQRta5uaFEIwla31eLu/ZVsw2g4
e0NLHa4Ccvls/9VnraDouhjiZWUGanAvgSOB5VGxaxVmhhx5hF9gCAlLQrvctJmL
tNhJ/aNAnROudkWoCpQS0kHhbTHBe9Et6ayRTrVXzjLKI9ieLxzrPYmdX2yLbVxP
XtOV4P2PkPwL/t1tLRHDmCmWCp5Oq3YjTvWANyUaAcnixyggAvGnf7sRAf5f8yEb
LkGIzvLkYLmRjHxd8ObP/glWad4ExSe2WgzlvEbSAZ62+W9TaNPGRG6l8LBCdGzp
1zFlNigvvzS0qpy1xuB7KVGFOpXvTyNK5fY1WkBlHYnpf4G8ti6wGRjsffrQbwV4
nQA99p8Edw40xxVEpgIWarl1ugWA2LLi8Ad7/kQfYjW+ZyubqXUMfHCjGcm2biJJ
hlJQ8JoKU4fIIof3mtfdVS81a0CDgJNqDAwbJNTUythWJqkzX0k/qKcWDnchNoO1
AGoxw0T3UhQ6ojKt0GNkikgfld4MgFUbu7OEzh0P17WrZ0tZDIgn9595IZrUTCj1
Xt4+4iu4iDt9aCHNhwAdXyEV4zSkiSDPpNzXavT2xuqSZWmLIZhv1xTew3L4yuAr
a8vLWHknv6mPlNdlVUiXh88QgpTyVFQ9SV6ce0hTppbFF6T1kDELWN5MfFiK+LKj
kLFU8FNhs1BcrCYZUGW5qvj6eaX6mRaDm3aVyk0uYRXvungsctgUyWwKpMSNajWW
u2W1sL6te9x7G4cJ/OT1oYnoAFsAMsylGfsQ0i4Era2UNRq9erYyocAGUcRVbIUr
latr8Dv1Gnrp/lMidM/RuhpcWrieGs1x4e0zXxHLtpZwC5iEH7/RRIs8ZZA+4RxR
/ftNUSI+VF2bITvmVzwZ/q8lM8HXpX98kaCU/P+zbd5tbnPhaagUh+MlsbYVvvoq
CUfpVhaxo0UtOdaLcUJkA4PUytuYg0ANaU1YOebVsyRAxD+9SmpmjWYIwCd0Si2z
8i44fNxAc3I8s6DwHffkCIZosZ0MCLn5LCqpo2InD9GBh0i7r5VRA24ulUVZd57i
n66FOSqTBNKo1XxvxUzX2tY4vqJ1xZ8TE+0k9JW2WAYF5JM0HG7F372Naw6wSdM5
2BLH8oVDRxxdlhi+2oHgI60pkUHwP+YHeMhx+RWybwu86KSB3Dv8My0MNOMn8S6S
3j8Xv82/iPffSC6+RnBZRvZwaykJFxqmnNJ7j07FWo9lLp+33tRFRD3x4w3nE98E
wKGThgYjAowYtl9kBu+mH6p9QVQt/7KLuwUdzvqBOXsjVrxdnXBphkWP7uPtaKLS
RSt6BxeXY2rcMozI4n8F1qD5pfwj3ICswvJADyNrkO4Z/2WcCbojXHpyr9CkVe3Q
vnIdW5NUWiF7ZLZl7CXMhPxCsM5tdiuCSN2JdKuNKleEIcm7QhpV8K4J1m2XXqLI
2E5v0wILJXK8zSchSFCxs3iY724rGCm126PRpUHPtsenutrn6HiOrppN9bMFgJJz
LZtQVimJtuAupNi9JKrOqzSVMHxcNQ9rHyTkf0wBf/dzwauMfeiXZ3DIBDEu7Tpp
udPDKAeQ62/NkJCPX99noLi429DFIF+r1dtIa8BGIe9SaxsyCVPAg2qcjtnl5hvu
enOczb5WIn01yx8c+Lj/+zkYqYOOFXR2HMaqKxw3/7GPh8Xc7wc2KGttlXPprdFn
NES9F+rR+HQR+8wGDipIpsl+7dhi67y5ZIb++XqZBZv5819JiMehjUezTVhtRALS
FoOVjSo0hwhs3D3JIrT8e8UxUBpWA7LGtCe9sMB/J06zp8OVuW8YAfAT9QKvZxwn
XS1zxqXD7m/wbU7ZqRTDAb2tqXtOn9UhBcJ3eDWR1LlQC77sTrYwSGXGwtSPIDEK
nmTtbxTYBiuwecPT2xd8QdKBUoz69UdRdxKw1PgithkwG/mubNOg4ymBceQlzia6
+JFFAzr1tFataTfQxmP7UjtonnC7zEwz5tBkEgSSnbxm01MexYs0uvkeCvMjhltl
kEpWw5yP1TZbjqvIpdm0rhn3P8Q4lkbR0vwhgCZlvS5hRwZUFOhMyo7wWp/zoetp
lwh0EMykthKIMZY5NzeEiCBN3KzU9PFHDc+z00BbWwnpff+bm1r6NVK5/FqNqOaZ
F2fIfKR74yTAaOuA9EujIyM6IEw/Vvl5bKU8Ex3eEmCAHh79dcQa18uaqFCghzvi
ulLqvACPJZBwsATzhplnD1h43ZkdFHdOrRFH86HELxeuimzVMruS/fpuIcY2IS/d
mFjh2D4UF8EGLqDv11/jc1tkQXysiK2hEeE/iA/xHEoUcK0ynfLSP69xaK7XAGnY
RHb9H/TJHKinV9YUKg65X+2fBUqWWHw4EnswHpg8y8cO18+s5h6meHUmHb/btHXg
gpHQWDfEWHWgfJFXrgBFIpPurDOE4h5/ri0CqtLhGjKXFzns40H9FQNTIzJPhw6l
ogbTsRtpkqua84LvmIaBU4Tf812p02fyQzFggh0ujPc/E/XjMOJrjlFWMY3ZBRJW
zcP3jPSNAi+265eA2auoEJRE2Y/RUVbeDDWwT/hZrR9qF6K/eHCvVYSPzm8Zw/pq
npmq9K//buus2+snZJn1IeR2ggQfv/O+nanKxUVs2vZLMfWFfyGgk1cUpdzW2IAW
aKYdHGTyvaU09jQYFwXbFcRdHEDZnks+Ht7cCZ7XEWctVb7ncrqP72CDGapA8NkN
NXURZ0l3bbz8b+yodinO6yGJXiZsDxafdOhWQTKMLeyYc8ykuVxz6UDrtNf9HRai
XzdsaVhhAXuP/P9230ZuKthWtO06mPrwAk9n7XQ25z6qypIywkeaAkgdJK9uP68Q
ZHo01WcH+Ny12D55iwpobf3klcQmlMAIqY7OZTmG6bY/kmZOXseDxcVSKTJb45EP
L3Aop1pFHwmvR+Olp4iVLKv1HmBErojrZS/xyE5bKkrt57wMS2rXRan8xPV/ZVm8
vQhRjxqEnIqlBka6Tjw7uaOGpC/TYvMg+Q43RJeo5wd3kZnKRMbpWDfqm3Jho5fy
DuSx1DmVEQWHwV0eoc/F/0REtplvknFDVsQekYD26oUJsqgZ1fhvZBdV51ebVRBl
5DXVcdrOJpBUZ+paBknPm8x2qIzBIKORIhxWnhZ43A/vSuGwJJDhu2S6/xer2Ddb
RHWw6AojXJADttjJjVA5mzUof7z7pwiZFDe+0tmNjHqInicN1P+Ghtxtn++jVASx
8KP3kgJwQwufWUmJ7T5JIN0jhKiXVcTWGbeINYZ/+2JuRcRo/TIrLYJmpwXQHci9
JxLJH0lB5tQncRFH1DjpLg0YkXvDl02RLAVVWu0alI94OIvK5MBU/CVdpsmIk0La
d+vfXOZw/QYwfKi4kAwvemjIEw79pgQjmAg1RAjmg7p0R7I33Cd8ijyjiOFYsDLQ
5bns4sky0pFv45jDSKsdtDLgZioUmCv1E+x7UhLWfQGt59asIganIoMp8S8AfPMK
kBcMlS6BqvDgWdcB9eYOGAZKe9SRFUhCgzDQljUYMW2H/8+CIEXdTmV4FGAJmJ7P
gGnad2BiljixssTWVGw7rjgtPSillZNpZYyH8X4Z4E8yHpPQh9oOygZOfM7IV9qd
fiNFWkQgO9RGdzdryFcvvumYPhE2B80vPF+wWgID1s3qkm8wasVDS1zgmfdmhRQD
MKPKKWujewZ4wNZBwz5D+JUdn4XVkuw/bm5uiHhDQ2hf1q1tYaqb1TCqSAFmsDf8
7pUcLo6iuyIEGv7IjbpE66yFaF3ABD0V+5X3J6xWVrE2aHlJIsu7xBm/ecUKJxYp
bTeFBY9iW/SKv91oNkJiaw44o747kk6cLEdegGa8AMGW2MPJ5knZXN7+fLB7S3K6
iH3mIgz0zX2EdN8q4yo5Yy+6m1WIkVtEETjojzg0360jZOt9nSihC4rN6l+appk6
ONKPPrfMoi/p8+VXyaYct0scIW087ba3u49VANU5GIEqUWrhdSDUhBdrKypukC4f
ad/JECvgWenftn8hNunQMe/Gj3OCTdMIeemm6i6PRGmGkF2vWTS2acXPSS2PoDuG
Bxg05cy5RC5YxpUZUwhy+fq4wD6JqkPcZym0WyGBxfNzD2nr3gVZw17rxBTcrgju
eC4PhVLO1os0t2ORq4qoQTkJQbrO+DX2oKWS8Q2XFSX+V+xsywHbVBABYElq1tWV
8BoqnMrBLV3PMWw8fvKaVPZLT9A0915myVHhHjoUyyZTNfwn2kZzu3MubCcrHivO
okrQJaKHgp1nr69sPB4nzSC0mgsP4aG3FAma58P9/8F/FF3y+SqPkNJXAbDUaojw
GR5IsmemV4qBV/TrWvp1LSK9AcSnB7LI6gkYZtTne1x43+jPiM/j1Bm/HrjjM5r5
egzLCoyBlkccEbP/I3XWlOB7YKo4YgkjG+KQJ2BuK745NW0zVDX3M1bVAnDwSrEA
oNEVlqVZUULP7sijvL4L4DwPtQxesQgJk6bh4lj/IFFlYczSBYStFfdbn56DTz+/
OJSGcxFK5SiBuWTaeK0KZw3tFTtTtNCoO0O5w7gfJYAXnaV6oqyWaeH21/AxhA8f
yq2wxK8aHeaVH114+7o7aF4/GPUUneeBAQUfK652k5kRHl/XCdJwM9SsxTGc85kK
vm2GKUusrAL9i0wjX3+H5tq+B5E1W+TX1rYWcaqxdpWtC5FTKcRjKGI3rRPgEgIy
P3LJ1csVz0TLTCqQ9V1J7TYlvv/34zTrYLq3G/dPlDP0zNOvWevLL6QrTHX7ni+g
QquJkbBh7TBTojs1taD4qjBTYoqfBGSK0EvGKoYu0ErxMvggyCUT5uujpAbCleKU
xc1Xu+wJHZpT1qvkkt8hv/m75HV1s36G/QQDf8R0ovjVYsy4w91AuhAhPZWc/AKt
9FcKTn32ynI3Cmvu2nFZmySrJX78JYuz8fVXGuq4skTPvp9M4Kb07J8LL7tXXLQJ
sV6kkxB7L4ip4hbEJZxZG54m3d+YOSJ7zvhs3ai+pHyDl/xb8pHYeHd2rj/AP7NX
fzuuiDIru3gND3g59R7QhhOVWpXW8I6UeCk0ABvJzq+ArQasKf1c8CjIxzq4tw6m
pAntcnYFqpyEluFCqZHwtcG19SyhvIAkngMD+X+DeiAmqrYh3AxL+GvdpvTu3exE
2WftvB/sie/CuwePBHpuYQe8ugI58NKu0ZD94m+HNxngB2z8eCKGiXDiXKV9kF/I
5Me9b05jYKjwMF77mecNqxNk83tdD5UJKoOuiNcsAFaccd6Iz5Yz6Z7iUnyUD8S/
aVzG7Xz9FGmkshFddj3oGauUy73TmMZfIykt15w3XDZIUJzutanTQxHachr/G4sw
8irhvcVnZSPBXkLXPA1I71aiue7r6ZJVDV/rK65/uudLEVNbhNGkUxYhszVwx33I
ygEZ4rkGEGbWM8eOQFlh714Tk599o86mmigHOFfLB1+QN9NmC85t/knrXaNdHBnr
wWAsUqPixvUrQL/HclbrsnH6G5EvF0hEoAZy2fF/EEknYKuwpl28ok6KGLHrYWwu
6rktfjsOfvFRoLD9+xr7b63vYTsSAftVQL1w0fiQ1rJaLSBO+1lOdfweTHRW1AgS
NWCpfOjM12V6oKMkYhJQBTzlRZPyqodDTN8b+IWQzNnEI6PQ7nCtIbQ1JhEwCcOH
/gunwTCpvB9ZdxxPRd5SPdGxMtLqYVjWTSlya4/hULwgUMLrfgQdQnU59tgXA0LV
BlZVGUepneJT9zyqGNW7ugtVtSfN7kNtCW9E7ogs0k+6SMFXu8JBXKlZcz+1P4IF
8fW8K4KZjBe2+GVg6CUg4PqpFBv3YANaPariqRSBFwokqXkjlPD6+z9/7XgUadLS
sh3HAen53LbCOz11iQstQJ3F/XBMrpV3krZnm7oikNYRu9gRJ5H/itQ2cm96pVLf
WvL0gp6OdLqiJ9BeXjg2PUrxJ1mZLez5Wblm0J6l8oPye1VFAyL7mPfqxSlFBi0A
nRxSjI/yTGlWnoi8OgYkJrmzcZHUMO/bqJG+gg4wPDRZ4zKYEn5SYf18Th16USyK
E8QB8jgYPx9kd0wvttSjMPzX+zgvNcuh/7JLPOqEYsx8fASJYXAVGQ2JaAbA9rGv
E8xbTFcJ1gFkgS5rGVdlM2itlY+0HB2fLEqnx2Kf1Cfdp14Se/dt5E8bPhhbvD3n
4Sum7zpvvlLbNb7oCgzHNLkXOi2qCwj+fgE8hXKHHSG55ehj7WvjrnFJ0UA1ZMGX
V8eNEz/jDFKiTQYoGDkBa6OhQI0na1HwRUb8+fv9tTkWV+t+C8NvF1czqi0HMEL9
gbQ1g64+dPhcBiQOpokdgmjUNyluikyWekHXIX06B+nAQ5ScQ0NetQxLvMdVLRo5
d4dfcX2+Ja9bgldrA3JEh2Q3fmoZoUCM+6DBnE9XCSpoqrcZ2AYB1+C0+dUfcLC1
MCgU2slxECs9w/h99SDy1HUtOuFuktSS/3Tp2qlrnybe9xz3c/GuRDTTgYzeEwhy
4sYq+FfCIQCjhD1tbdzLfTwYvm9XZssap6iET8cTDMS0yS2hT3ib0LST2rI8R8Vj
3ntHvnYSXJUE4nDWLZc41nZsPyD43kOm1Skk+BiMj6MlYGWMoeAgZCT7cVLe9+zk
ZUEHYhgpXEZ65Viv8BApa9EjdQOu2bfOsZbWE+XWcwXqTH9iWvtTUXTMQRsT6xM3
pfi/6GkLer9TlavgJWdVMyurdNnIXZjs5at2M812d53Rr/iQ8GWRT+9GAZqmoLAu
RjgP9O8Ti0CXgt76RsCRKMFHxBHC9no2jisAqitsGVCVM3DEb3omYjYZIlHAFWyM
+ECqVXcfhW/CJBQ4EVTFXcKOes6biD3RAfz2RXV5sMRr4zG7wxvcLOURcoX+7mvq
AgUkPRBCPMfUmE4jvs94lt8tHj2TWZGICxA0b5wo28Ka/WOZrqHRUFVQC53XaauQ
m6bsVJRdCyVgvRPRNYZZBo1nO2F045cco0bt6P6TwYBIyWnsoU5dKEnkH/bmpZIg
/OG0KtJw/69Jq7ZKBK55k9IHy/eDja7++hvsqlBOIycVX5ie/KMzEYDAOApjOAkm
x3r0K3O1BvfaOt1G/MDXsija8astd0IApJDv5nB0797f2fGQZVQxWLTxCfWj2BtO
2L4lN7xfCUeBlCi8ARVev4dknQiJB2en9jP20wtnr4Wi7cV8+/ROuSPUArq+Lj+/
MZ6z3OMiucvWFUBfaUHzBH9p4LaIO6d4DDFMatOW/SMr9X36HD0efWuD9+vUqHp1
zo4+xFLFhczJxwSYYuI4hSUdt/IFsqe0Q/2s56EMbd8/Y7IkbDH6lfYzWk7TGM2d
3h6XKK8bQw39wL8D4WRnefVmvhfnQCbNZdyu96bKqDp+D8++STnvFVbs8yfaKjzG
fuUedpT91gsYre3rAF/tMExHRGJWIxwNavZaiudMWb0knREjWScocWA7fKnNSDSd
3st8M1nsn6CWnUs+SMDC4KZ7eUl5HP1NxhPQyYr9c1bluyuTySCoSLzqAvZCwZZi
sJo/HfOuZQQmr33AY77K3Qc9Hi2ECFTSrLwcXIKfPl7DqM1ZPrWMtZgFs6fDhFRQ
izpie1sFqdGKO67oz8Jb7rBOxxJgjT1bwrv1U4kNkZiXUvnj2NdtOFoTp0tt25WL
imanx06oCJH1u4qL4+k6805SaD0qT5eknD8GspLRyCMyA8S4hmsyc4uS8XSywZFc
FZCgpMECp6bBfcGp7SZkXj7vvvnCU8vk32Ti8NFW4M8JJv1xfkm75w1bETa+H1Q2
oDkTwRobtP0T9SvnT0auTN0e8cNNq1e6SHjWKqAjfs4GXaoVKjEgydnRmvDAos/U
1JlR6JOho81QmHI3qUUGjTRKphr1O4RjTFiPO9WiZwHUoyvu81mnpFqN4tbM2UE9
NR0VI889JGJXqqwOoxe4gjiRI317stC80FhKEYilGeaPQyEQXFLgfCsFh6CDjp/4
qA+LcOdVnDVeOkwGe+CXgdOAplxgZd50lwpJTw91lMcmUoDA2sG2vFG2s9baEQbj
YRyRoGFBIIep8RhJojL0bPqR4Ih5DsvN3iwF3XA/Yn02ooeCh0XalLrE3dtZfrP5
fB6HhzyI5OP6I/630nqEr9KuEa7wm/d+0V4RcmU69soLPmc54Ro3MSevQGlHS2NP
jG/p25HirqEdlkpOTfOZC22BeXj+wvsFaF/0nEsqnBZw2sijjBLbWy4QFvpnDReY
e5I62hm3b6pfpBpp/AgId7kAzqgghBp2jDnOl0ZTmNrlaCJJ9kVLmMoEcoyFAJ0u
u96EhfhuOpblzQLYCSXlXJjK47VPbaODHT4/paDei83iWGl8Avf+RwP2E/nGaL+u
UkdfuVfWcatp7qiZhBdmFxOsDBZ9ozqZBw7oETIz4gTKB0mkGbGczJy4KJmglZjE
31NcIJaBw6F0oB4kBE/D4M3UVPMeVG9LwyKQmz3Omoc44cThahO7igzK2GINc962
NqFXh7n4e87drn2aTPQ0kP6hAj+84PIdAMby5BP5JkpvcpZbmzfV7JqxX3S5/34j
Z4m57JrLxlKimBGXPlEkGkGrDm5fiMbhjHNO9V0ckoIu0OoImu3faYfx0Ay1dTQy
+8Dz2fZfVH69nEU1NcX7tCx2IdlMP/q5Soo0zSH0kQ3gPZ/FKuqRdDHfPqrlQEIX
03UU5XYGuxDXv4JeHmNhVSs4X9smRsnxvs5rDdK6ipIRKsrhAcIzl5aUtY8O4pOH
kRVKPrcmGdoWLcLDzhniA4uz0R5VK05HHrUJq4FYVPjFF6jYh+uF/wW2NkCNaeI6
E0Cu9taBUPJ16Ju+zad7V9kvFTuxhu6yXh9FLqDeb+u+JKSbzC9/it34oVSleuF4
LnupVwG3HNogQMVSjIQQRQiwrcPAxLLDw6OeGxHHM+eJtix0F6jkEK9JDxW78lj1
ySJJpVJVzGC6emcdmOsn8svG+qhAX20AmQD6nW+1gPHBFoAT+IfxagtULb6iJu4G
SMgKJyN0IWQVe0yGLwU/5gEFUOcwmy/2zC19qav7gr7gEO7bABjHYdVP+ToY896t
cgLpJldBkjK/gs5r1t+i3+t/EDDRTmsw+rXET7uLgirljJ0o2cTtrg1w5ynsOvA+
5mX66DsZ65/9Qh2Us+YweJubg4nb7CxEWYSP68m9ro/Qm4GDmnIPT5CCubrnS/ds
ZDrZnfuySs1iE5ObdQ298fCo5m2ciWgocWCO1LorGwLKZnwwvlr+b2bKg1Is1gWW
At8IT53j0bVAfHYTJb4YU/ox6pNcEHMrTPqC7iDxigB3MvNGofNs7QaBrbjQves1
UjJT6ZAaXGuF+kd1GdTFpHzmeDYqTUB7qouU3gzxZrcAccuIU2p672pLOC/eTveL
SOXzm0hw44Do497KY7VRMQ5QvOvBpioWrn7I8JzEGJjTfsfGDnvZa6jH2LrI55GS
em+LIoP1L/xR9sA3m8AE99dlNjIn34AXwCSp7OOwqu9wijvZJZz7UfqV4gqnCD+z
hU01Iur1ep84I0t13zB2gSXW/2A+TQltWnmmcxYJPSMvSYRT0KRdmFgNUd/Yornx
pCdlF56TD0KaXaWJ0ksVBOO4uUDc+Ed4QXoxcs/CFXmAOwsOp3PVrIz/g5L4Loik
ZKEGbqu8uTTXB3RbVbYUwilk6kmuVKfrPuJVTBPLi2fi5bfmkSQNuC8O9+igRBgg
qBU7QfMJuEcMRhqg8LWFsyskirNnQ1JND7vBUSqZdMmySEI4jfRA89ZXd4aBMiwl
IicDmqBQ7sI1BXDtdDEumYVjA0qlOM7whyZOEhUowt9fuV00IXDo7qm2StTFWdeg
pLpV4OM6KQ5JWZm0lbl9h2ELm9SnX+epQ+6N0JkG2JcA5HjPkg7vUkGZK2EHUqXk
CNRaIoTrnMB0CvD4BWnaGteV4obiDoJrZ6fDhuN8IcIST9XQw5vkcA43s1aKdPFl
HeToK0RJZcOhKMs7mBRC3s5SnPRocXeK/mxeMkYpbPq24+3PflJqOeZBqUEMBNbT
XJak5OSRRMpjB8mwaDF1QyEiwrPOAd9Se2sbO+EbMGBFHpGHZR1zsaDIwvl4/XW4
JooH5P3z/Avh3Mk2VyxuFdC1+la0xYkhGGpcGi9HvH3Mn8hQ5JaUdTIxqXOHlhbe
tZrKPTsHee+jNplia5ZYHnomtvu1xv2CfWp0BM/bCibL3+mWmeCgFQ5aeyd9aqNw
ABt+hUSPgNYI9IXrs7piGIopCuYKoThNjITESWMbUhiYIcc6zFtjpJLKJgltiz8S
XaQAoxFm/Ws0ua8r3b5aBWIR+O2zhasmH+zPUq+ww+oNjXkuSp6sGl6Uk8N196ls
nRUCy/PaTNc52EHHby1tQhpw3b3RYSPrutYhOVRAlL30163rWYW4vWOkwro/6QUB
ksO0p9B8vMQ9AiIoHl8jXbCTEm4y3E+yvy4KcBFbObUd9OoyAFEXOpRZ1onT3G/S
CH6B43FZPsei4Qfb1heG+Voymio8qvAy3yUmCmblezLWBpJRLCv8aQhkVJHdnnbQ
gGkR9Cbr0VNeECSOJrMLKuWgW6KF2M1BEKuQZCFT1qMu/n0FscGxOXpkEx7NCOp/
36OGFjFRuWJ+XV2ZsVRNv/jZ7JYoQrB5Z074FhFTbZfQI9nZPtl+22/++XUn99So
iZ5yHSKoLrAV+vGbUbz6cetm+XczwCHb6PxSI80JZYHE7nUH4wtoFVeBf8/7YLvy
VVPtHh3Ln+paj5Jzvp2G/ac/e0w3d6AxbAEYliQw0lutVWvEW1MPniTQWO6JZs9b
YKxRW0F+49GB+jOr71QkVFsNfNKzp6WRPU3nPrYXUQGmQIk2CKXFtdPhOXzR7sS5
Zcy4oX1EgzWA4qDokS8cWQ0m6mvLBjeufvWQoA3X+4qkFQr8jjWwkRRkRI5UDBYt
7iTp8Y96u0a4muDasBSseO/res5Z9ZSSv2IMMUZG9NMtmQVTKYbvE7bnnmNLhnu2
gLSltskUWpYQYhbEcoqgpuMcOoQ+9D8rv8xYZh2gRy7s6lKY1rBdwHLUWCPyD8Tj
2ypd8IMMS4EyvpUJt9MsOxKo/4ZA7cS0THPSbFNIm2iFlIK9exsqjtvtX3qmCTtH
CdeWa9y9vShMsIba3ChIazdjCHlF//i80rjuMBOJUumEWxBxhI0lrHe+mP9PrKMz
oiOGISiyuY57yFtaMM3l/6ER9+9lKyxUlIOvkc3mY5t6BdWrMsMm3M9D628ktpda
yibijJ031x6q5xk1rlb5DK1Dd4JE4ehDVGKMgAAjnfX+lzxlTp4j0yciiBa2D+CC
G6igDhcC+psRsAFAsKoVCnU2OXaSOG/2x7hmQpZRHR/QcejAQLOVGmVd1nh5W1Iw
WN1Un8HunEyExOk129/kRA+UY2QlqfWyL8VpSM5j+W776f3HeYjeUUNScpBiIacJ
pupgAQc7ubBe+jTCorXDJgWYgd2Zu8rs+LOl/qkwpHkJkdfMO1LSp7OuLphYR4bl
psEChltHhw2lOFQS4Uy7EFCedeM6Fr8CEUWBGHB6DgJt3iOW/Owi1LFdTmn+Pg4k
RoJiq58w0y9eaUHAlKERyk8juqp9DyHoZGYHhi/7qXgqb+4iUirVT9zaW0nvr6ZY
SSgdWWuSdgyKRhuwN/iWrwBNxiJRyNxo31nVh1h7Y/Oit/iypze71wHmt0zPMrCK
pYDiDtEyB4rgfLywXZxhinL+OAlYT2BMT3OIxdWxfcJYvBQh2zNXhKzZyT4U+K3W
KEki5VngcxLczrBqVGgDd1RYFHgDLdLS+QmpxLuVH/QkerFLtg4MDj0dtCXpyXA3
vQ2ytoSrlYQSM/lS5wvgToIngCA96BodD1zr/uBTgW/dANVZqfKVIKcvMwdxu89x
hHPK0f9FqXRflZToGU44gLRYepQgQ77j4bU1BZp/rQfRV0KB6PFG1OELsKwJzQcN
tQDdJPPPEoQILoIkP5HCNnn1OP/FDE1JCDRKnsbR5lZzeN33FXBoAg2tQAiVsoH9
TNLFoZgGdNsjQlY7UgnZ/iDXWQpf+X0VvyxJ3vhBdrSWG/rQQMNp5dPRB+hBvtrh
+W4WS2mrD6zAIxNsJ3cTjwYxDagmC1tsDft5ztmGbo7HwOVh8Q5llROYWDR2T4mz
SlyqwYEYJu3TU5ru/EIhy6Sldr3OyzuvLsiEr/W3XzZtsrPQxflQiv1xBXdLFoUm
ULI62iFZMx8ttp+/84NVMCTOAyeiBekBKIJbpZHhNc6emOtCavLh5iZ/iHUL/EKI
TiMXS9vJrd0Ong12gDRbUW4F1eoR81dkowGWu/zn2nvTekmgF7YtSs2aKrPIQ3Zd
XbbF+7odPfUOiLi/+WUDwDDj6exeXoJGQQ1/EtTjaK7TlP8aOBpmnzDp1e+k43E5
U97FWUf60iw7z0Az2IqMmo6GLrMutqOmcZzi/HFM6Roi7lXdvywZJfZozmzCI3EI
2m+rZS7BO21HC3UNT/hLnTZKX9HwCPOE6ld+yCe0tVhQee/vjCTpyRWywQ86vXeh
qiyVq+nccOwdlvBD+FObt/HzlGeW3bKWrWLFVnSPIALGYVqqiSxfIwKtFSFWieEg
OEDXqTB7Sxie3W6AKcdUmOQGXiwIBNqzlI6wlikys6L9Pu7krgBbkkfVCw15k30e
RvsSaO6Hy52dzWHUCAuttw0cuCujKcaNi959fjniH2xlIEOFuHYLCYP8bKbkyqid
vRj+uMpLFgX+0sHsIFpqKZC4ndOJ6D/HmMjPJGepqLDn5NO7R1KFNuSxh7dua9Ro
PjOfsOFlavSUSA+t5PA+k/JEe8zWG5SEIpZI/h51afa2Po1thuSfDUK23Ha4brTS
7YnJFdhDm5urOdXbUs00hmaiDNweZDNk0Sss6hbvXhzE08OjduUl8Gl8274PyZ/N
tmQvpn4aRKatmcMAV9ks9FFqulxFoemqoOJkuPEggMUeKeXPT0VBqVPQCL20QXqI
Knplzg88IDS4UIal5pZFRUkeb2Gsbd/wBg/wQM50q8pG45G7Q7O1+GUsvRaaB6e8
K4C5rvdmvO4iUEKV5hVX7FTHNTwngnb/2qRegGhpbwjY0K8mXCqj1tLl+TaSqgvT
7PanLWWWdXdFZBl81dSzdzDfhG2EGpe09wffXv7d4OcqoGqD+Vg8qdKmGHORlDt/
92HiJZ3zWf/2TNjPl1g2yF0ELGyVPePsyyXhiIU8SG8bwoEPL0j1ITnMBFr7hNcj
rhj1OcW71NuuBJyaf1kM3B4EDZ+VWMFDEOxTxeJaf5hkpZcnbEE20puygOcNO7N/
t+0H6Mgj8Y9Ekl0yGlle07EB1mt+QqzD63UA2mlx+AkRbvEWx9ARm7n5YonSq5HG
btq9Xdylke/OjQ6shdIX6le0z0PG20v6eLq26I7uQ99e6SU2wkMk1Dd0zmiZSwtz
ZXLOPQ4Go38jeWvFPC0ljAgavUpMtQhMSea3PjKVMhxnIfrGLdFBHJlSU2Fqm9Vg
pMUXwa3b2uxjGehkGbrFiZKaEqIZZ/hodRRgndS5rJnqqm19dUWJdtBp5ctHiBMW
vmaSjKEH0uUaoBpz0emabq8eMMm84l4+/59yrUmNqjkU1z32E9X/RUMww1uyng8g
VbnmslkyWM1DJ74tVMxdJClnZweFf3d17B36ZZJr6tnEGl9X6COyoR2lnN/5A5/x
KpGfs9U9KcnyjE+d5I9melIktWTTWilRvEUlQY3xmc9Z/NEevw69lR5GMn8vLBJP
FRNZF93cUUHhS1JXcgtglLoauROBKVKZZ5cdYvzfoHmpkiujY/8fcVetEvWxrplU
2g9kkxRxojoyU2Id1w97fnhgoKk7NImy0bPwI+rbC0VRmoZ2SNDBMRBQ3k6aLRsO
0BTM44WFbLofaFfHQzTGbV2xs/URrV1vBj1HKMI5BLCnHWx0m3rQ0POF3WWZVanP
+zDEL23pGOC9zZ4Ov8KVzJGOEwUhrhmj8jCu3NDX0ebuXvWmMAkn+Aizv0o0DF0P
zS1NpPx/riMMKUxjwloPtumoesR8iKi/DSy2+QtdSX57Z5MYLoVYnQHRnaYWE6Pg
klnCnQFPGvgMcoc/NiIFZh2LI37bAd/+muNKMtnNmNG1rRzNj8Io+iT28mLNLsMg
xiC6T2iReq5otii4raU7tTCfqXivX9Nw1QhEQqmnqW80XrQfd/mYN7o3dDqNu64A
bUkIGfM2Uzv+N5d6yjUUU6ZL4cCauQafkYZ+BQs/BSt6EjGX3YgLS7oYLSninrT/
ifk/xN+bqCp8M46jtG8rWLXtp7eDTNL5LZVCgLzotz3F3uT788YIHLDxPE7pYSXE
OYp9KVovzod0iqEYOvRZvUJAkGGShPgto4sIDE9Xi8rZG+zpeu6VLXrUElVTf2za
LpfQZ9cF5gkIZyGlPWjOe6LRNQ1vd4GGNVy+TzkVi7L/DO5ApU9Q2uVmBQHkVjQz
DEdJe1TnDAl95JL3HssHSc+U1saY7xi+8Dhs5LkktbjTFL4uQG5tJcGN9oJVv9Ym
sDicHEA8B4WU7wUeDeTwg4odAAz2ivfUhXphAUirHzFrUQKgZx7Y6hzwGJeH1L/a
z7zMUR4zcbk8h0O0ZX/Uh+u1Qe3MtbcC1RisVBj74ujiNvB9Q1mxbOLlmdCzwTZ1
KiVYEU28nw08h4oD8LPFNmdRhnrFfwV3L14bTdaKVTDjbYvSzupjAPPIORqiTs2R
vdYoJE3VPDjQOwBd/gGdFhMoKoicBw2hbtPcgYTUtW6Cw6u+l8NzNF6bXsXJVANq
OID3A/vWQxfqYB9YNvy9LlO3n6WXpFgjDvq4bUqog4vhth3G3tVF8m8c9vbFCwAM
marW5GTkcwernxHStddZW/EwMwwo1Qfl91mqGdlB5mWFBTJivow9hHUTB5PwxMVO
LKyp9TCjCfHcsCNUkDNPxWNNi5dNCclkug4NwfVV71o+RKU7Sb1oxHywnYjs1KIR
qr1ffZU8i3W+b/Wlt4ErgNtxd/V9wqtD72xcciAMX3EjgQzLjL1H4zBfmc+vmTmC
be0OaQqJ3WiSOcfum3dtfcRSb1UDzGK1Hkj1kaUEZRmeOtDhHqwY/tIxuqRhgTgT
RqdT0n0Elu+fjRsstbhVA/2lmCOO2gEDfytoWx0fgEZZO2bI2nE+jEU3DKAuakIS
/8tFtP1QpZBh2xXd1gUGdA/zdBOatANJL6mlM15cQXVVnr6ltEJqek64JcWc8hpO
pa3eYqPJG4dCb/aCAxZdgd3cuezSN8/pouIm3VYUBpO6tUioNXR5k56tU+DHnmor
oJFTnWjRn8D+RyNnMB4pD3nBErvjunwAygrjfyfZ044Qy1J1Tt0g07A/69Vl5zU8
KX6HNEJbur1TxNoW4pskQ46th1PmsMGJAtHjxBdKcxtJx2qnBVFx9wLY4zupX2FL
PmFLvECJrvPJHDYFoOPL8We2dZ9sXzbBZixAZ1d76qcFumuNtjLBOg8z/fYovbcX
RO4znWtrF4Ac/ex/y3RNm3crZ5cjmQlGt9qWkeEnN7su5mmNmKI+P54vC72uKMHP
XUklfXh7pTVXivnFRZFHOfCNSGz+dPBoHgZ9OcsYkr/gz5gaHP4JBwRSKGWu970a
ERkO6rW1PRMSVqe5slIzT5lOwmMUiJUd3u2jf7mrn9TH6Urr8tTdpp1nq7zM+8OE
dNEFQ2/hkHmspUoFOD6E/kjWCrShJS/JpVQfHEzRraFfBXjh/yvj4GSqSEjBiGnZ
O+e/ESNRcLG2JPtFbGhaM9iO16ONRjgjkPcIYNpI2XMPFQNVV1t7qZb/Xgd5Z+PR
k9V2XB5oQCHsJzLjEc48kuvaNCgLkYVEy01csJrQ7Fx/yx3+21bG7Pe0bAzaRhHF
vMIM3fRMkwAmD7+73F+0wOb229JOBMa1NTjHHUq5GhyjZ7+13C8cKaRQwIR+C2Xx
jKqUi6sdTxn6RWeD80ma4tAJDp0mBbFrKTbBeHDvCfpuJcVUE5QyVipYmqhPdbZz
46Bbgr9dP33LPskTh2lpYsu3gC85zeSTW+mKi/49PDkLAYsxeURBtQYdyCmwomcy
9/g7EIQvZkK9lN98eEszNZChPQDLV16f9XACrxqK597TRnRhdVjabZoT1hNCLwi2
slHDPcX4Fvqkq3v6hbPYSFaIwGmcoj+GGP7A7NDZV3H+Bjw20BjEE0ENyHtqA4hH
gta2/uEUJTeQWUMwwTmgU+gjBZDovqMxBuBMsCWllbhY9SNxaauiMnmf0/NrpCsH
uFrkzi555xbVR54bR8o+OY3/EGY00oCHQdmEb+eiMA9g9rQ4cSm+NFYMH1KQy6d7
Nje2PJ8fWpQIG6P6BWlIXGHaD6p5vLRSj+czE8bURBZm3OEFtgBJk/hvKUIfbH9f
SQupeYDy21SVTTtthnZNk3XTytVxQfe3K/lPH0qZpQwDBWS0ICE2l5sj6Np5pbcZ
rTLRSM8mOL1PzOFbLi4JrOoRnOJHLYCOHex1k0C9Xq2B1sxtVIhskv9M2tnSBC+n
7H3arvG6GM9EaqgUq8cMMcXzAuW+zAag7idrSPewS0bpZIGl3sJDQRVLIETCwLfW
TuFHhPGxjtz/efFEtuCj3zGcJl8saf8rc2uvg4a4lUs46qE2YFOJ9ooUyD9Zp9vY
G+ZX5+Y7KaqQD8XTFw4T250rRfXEH3Ap8y4Pgj35/EJKg3CinzeG7snTLoTcAF8d
v84cCKpqPgplZl+fDXRMHLaK+NxODyVIDCyzhBrzFEZb7bxSbyxiKgSoelcA0fdm
o6aSBNaP7VlQIu7NJjKA4bxF/weag+O/JRdxrB2tz2CEYguPdAf2dGiLNJKzYCA8
LQHWgPzHlC/xsk/iA77AUFNdEk0N4YOeybTzdHcB7RPxS26crbHyv779DLdjcG+M
79se9f2dA5xNDpG29wktnBtjcG3Svq/KzKXnFgw248JqIy7LfK7wobge5osdin19
gc3MkeVHUGlbmUGjwKsicYb4PqGQx87ncMP16CYhvfEFLUfDCr0duZLzlIMb9+MM
q9UW6qAZuyn4jxGQVPhXwVH5ZEgR+gQPOpEBEPgTZcSqxBEFtM+7H7tiToi8cxbL
H8pJL7m50H4iN1OIiSWkcnpL7g47p3XSh/GBBr+km6Q8dSV8s/uBaFUXuaLbTR2F
hZ/ST/b8F3WJ2mGhTAytZjIQ9s4GNw1Jc9ErIYraMfT9U/6LGMXy3UmqWhWmjbye
WYG7GV+o63/Id4uk9Dz7Y6imRHKoGdCDDhPnGYEbnzBtwIkwuWgolcr2z1gJCe0/
uDvDgVtoyCeDRDezt9xQiUkpn8wq9YViO9nNKmV0ov6tCyZfhzFGBHxLyXRL9wtD
5XfzQQIX6WFunoYKe8O/tfW1XWSNhFhz7w8s8CiFQ3Cfzj/5tWuBAuPD4snr3vbJ
agqdIZ1XLiyT0VvcYayOZurK71SyiiiPmJBixRzOrXSpEst6BqELi8D6pbPRgdvz
iU7lffH35AP4tIwnMLfkZaD+UqZpEURVJ1osPfotjK6pNJf7zk7z2onUHMUC/xaS
lga+kQKsAFVRZYyzJIx43nIdptMv85lCIYx9OLX62XgPMimOdpwGMJYL3HHqad6I
lpTDAOR48f0DILpCWHnzlhhXH9c5uIyEoybsQiAqAo9AzVqgV/1gjnO01uOzsB56
8AroNOyXu0t9GckGduE2kb/6P28J4dqGS00zKYVKc4vwZ2JOP8xDl22/qdsFOEnr
IgAI2VXZKNL7eCh37G1U2iee5Xsm4uP7XDVz1QivemK5hmEekV6HOmglYJFIEUE0
ihZO8oExF6e0gI14g6f61btExTimq3z4lHQ5mgGV5FyyJ+VLZSU2TNd/uEunIq8a
Mt9qYlvUtL2MRx7Lmil6Kh9AWjDAXJGmb9PXJ8cjP3ZKt+l4+4Na/LeUU1oodJNG
e6XMB5xCTAzMLueaYRdDAa5I91iVZmTlxF3GkwTh6JPSoKs4Z/Xikq2U/oa7xvzA
DB/ESow6gb1l2P6o4KnoMddn+zaiVgcZXPHsm7UeN4roU+gxbnjBbE5hWn1J/wX1
0roEouMkRbLwqRxZyoMK4lUMbCJLIEr+KaZM9EYY1+Mzsc2rgS2PpuFfNOwpFfC3
yC1nxccs+N8mLjYjMzCFqOCcOb0ufkQZnR8uQAceeDE9BOKpcBzPr4sOinaXyFXf
XlZRABRvozUNbBrZN1IMo/mwmwK16zb3QREx/EBLdd0f2ghQEsIuZZWoV9T+Kq0w
7lEwb3fjonK6db4JmtfAwoho3U+Ksm7HEv+OlG68E89hVsqwzk72sy/CEEOq+aZd
tRMp11O9ZbOmu26UbqZxDerNN46oAFhwIlJHy6GfkZDX6Vojq64VFffTTIgcoEfn
E1wn245AKTMRL6jV9Orz7nHVdx8NDKmNtEZ/oMb/87aAKhT+2I0Z9cok1pt7G8oJ
fKvhR+ElIn1Mxkqh/myJwxEGYjx44+qNEY8KSZzkaZ4fxhHi4E0/pk2FEz6v0r9+
pAVfn+2RexjDBz0BrzcXgTrqwIXvL1qjMuFPOQBMK8Fjg/ltSZd0gyPO1AKFXRMW
GMHIm8V29uDIDi7b+lYmncdwO7bfFjy7Pz0AzQztNUAj5UNqLCPIupZtLHRpeQgY
0UMU1hFIWIBtu+nTdo+QfabyBf/YXd2eghkkrsyJ//tnJVNANCB1lDpKddpDKuyn
DHHEnYrGAPjFdwZLFxyidJWCAyAXZ/In5l46K1223QdkNxiyh+O+oJTkj1SFrzHG
HlxQbG5pjBehukJiR187ZtbgSppS68RY9hFyksSOqmxI+in0mRxBfPOJqmeKKgNN
jbvZ8j1eyt0a5j9FAxlp9SmAX2MZ6+crrcaGXOZCj+917uwstO3uiA9ovqRP2uIG
CZXOmMElrrkrtVFP6EhNIiPx+9Z/+5xroKyQsjyaJtVpTbNOolLO5tZRrp9QZSKp
zLu2lCyDKgP5O+6mf97FqaK5JoXjC8EvIaruQYsdFJfHT/PTkrhhnX2eh5FBZmdw
u+USDr7RI+KnmLuO9LQbfK4shiarpVFjBO9WIKBn298Ya4EIWlN5NIYswra3mbtM
yC1OvYg0jrFqWm6p1ERUaD92m6rUEa1jEjUYQI437QwXVafB5Ue3IIHdUFABM8Sd
V+eBRCjDv6p/19/LbJBI7X9afeSlQCxBLI4vsaFNORSkBfwKN/dbPRTBMuSJaZxs
IkIkVsajd/jS24/s5PLjx1NWw8sZwMcDxJHt/Sggaz0HhU2JwayQH3NPKs/o8zPJ
46WpB2bFPAhg26AA52L56zNM70vfnqYnBFs+pzMYih/K+5sWsnJmH66IhK2vmAar
vecAvnPHUJIBab6c89jwYT8/HgpeWTQB7Uh7QnROk5Xz6luNddaDmlxUkeg2F4O2
R3Wm8sTX+NuK2T7b40R8h129Hl63ACRVS9RsbmrRZqZkck7TE5wDghaqr5TaMCod
AVaSPkCYLIX1VHX32f2r7CGKiqCjyUpAWzFZJgMCe2gJvAONsH3yoPAuON0q+2Yr
fyjexv0GSxl+QT63kqbr6kBln+DLn5f8NC8PIg78xRGBRIY4vd2xpK2Yi+Gx4dow
DNt1hcRCa1TKm0fyk0cGCGc/3tObfPC4n6411yuYLLJmaP/HNKBNbB8WczFp5PlV
ikNPnQDwrXSNMM1QS1aYBHLZsW2WqPPDz873p63rmoamn8xQ06YNhGYfvZFDa6RT
SyxT1347yq94beyUEbPXX0d49nWL2ilXTNfprOlZTeM+PwdaUSYh45hkbBU//jnU
21Z92XnbTg1uJNwj2RIshCGTNPVuk6/GtdShfWKC7ibJZrsxk1iyV5i9pJ+cK/Ue
nLbcTJDNm29S9lDhwCYpDKYpi/6FEAizhRoIc7D7eMEy8MlLRCfISyvh/c8h3YQ8
fvf3C+T5BPGSMWgWJyH2JRpr+/IyUdwbh9t9knOhlbFJ1i0Zh2iFkLhRUEZXs00F
lgKh7g/YcJNcimnduNsO0RePb8mu1Iyp6qUK5XjjTKycfNR+73tSMSmA8Vqz996h
9lHFy1d30c+GxLzr/L+fNtIt7bQvB9L/OI36/9aO2k802qdXICybmM/8n7tkrPHa
K74UC2wva3gpiQPXimHsFvWkXmImPKuA9MARP1L6N/KDwJAwwZ2gk32vXbvszjEk
RsKcD3+iZbfNjp9BIjQg4l/gVf56ifWn8TqoFcNRzMbS24faR3rZ2WZm6POOtxjp
GtYbGAZT1ejDbgaXCN5VMYkQk/aReZnWQwy5kZiEGqVhCVMLW/1Ho8cspR/mzW/5
Maz08FoQY8GXSUdMyli1VC+EPCRv3wxZp5U46SPzLA3hAvYi8Lq4bJ2adn77WAYt
fojNUvBOlBGuuGkb/ZsrupFjbB4z/zggU6+mBaM17Se9M0iT5GTts9jPyQ5nSRRI
1H287AgcJfYpfraZrEhgven2ImfFeD7mb0n7NxVS6W3pkfvEXQwMMy4o+kX9IQ1F
EcTsVNJAQ0PYP9YWaSSXygqfusjeFmX8r6OYvVFa14avV57Ish1x/8t8wzAjrsBz
im7NHm1mHHlZTNA9DlTkAbB/CmVimo2Bh5bcdR/XkOFKE9YTmGuSlCU1aYcYZq4v
ja/AA9XXgTsGlxqC0ju11932aXNcMFaXazdhsSTyP75by0pA9rIyd59CQQ++jq/9
yu+9xG2t8xAs+hAHynjG2vWXhgUtkG5KM05VAIrGhhOjkPhvWqJgpu+Tg/gKYSsL
zn/OzP89y5/srOn4ie16SfMiCaMly1nUTEbe7IpXIyzQYDe8nC084gwffy+Bhtzm
WhawlEk+b0kCeWn9sTXbvliYSIVJycDGpcAUfHou1K2gWEl/W+efX5wAZUoaeOHi
N9pmvQgar0GoskFEmjE9DJSewoffpmNlK9Vji7Y++78wSYcE1pSLFbbgrSyEfgrK
C8wCElvNoVaW5sfpVk43hA4yh7E22LbratYVYR2UToXNMiBeEzplW24lLpfOvqxj
QsktAYRbll9epIjcBYpEtMSjH52unFRmPlLBFw6ymEFNyx2ULVp54VDAiuUAC8ok
K1FpryEOq+sEniml/ece9isPdlOOGI+v9Zd7xFp+RC0Q76ELWzLGeLS949PKd3Im
b/AKfET+MHqxF+Xg7mhsY5BoNc8zwpuxzbXMS2crelcBIIzkHzhIEnKmCd78Cr3K
KNZ8sVkXYdRQryTb2PMcm6CuuejOPFAbb/PbBjNbHukRkG7i2cnMcD+jvxrJUcED
qUC2ZZ/GQZW1jA7uKyP9MET+IJod1yZADyidG3ySVmmiKze5ZnJBrIc4SAoREa5F
KLEW/KfznvsM4NL8qfB1HN8nYlrlEzhgEAP90ir12NjFYd1Vrb0nMft4LxASdF5Y
vykpKQQFs1Zc+yRFLX8F8f7IyhZCGLwu8G3N4W7UvK92Ptd3GEDc+9reyHGHfVua
P+7r9QCtMOfTOS4yMyKD1vkzCM+bqc+bPRjOSkkHZsBCoDNLeW5fjhVDuhLNSxpa
vthxanK6HmlDc1g1YymiIODDlXNYGH43RUlxf4y8h+02nNOKo/CqzypkiaUtk0b1
hQxrl3DCkyquUTqUl1T4ojO65Gabyydznv4Mv1ePBLKDoM5s2SpzvH7N/istTfCK
I+K+rYCg/LgbzeHucO4y5/QVE1ug6Vay39EJNwW3ckyNSDpwCUvcQyWkxLz/j6D+
JeY3i2HtqSNsxxaugk2HnV6cINbJ7HL3IYgGicFVBMROvggycMGWobJDPCX7MRDw
nB0XTQRVHiAq6xB3thPtu0RCAnjmT54V8C2570kqAvIh7+RBeqZ532YEs2Nc/ipN
eoeGirmtl6QdJnB6FhMxQr7i6d0tzvl5T0bt5AmkLP0/nTwEKRt2Thpa/uHaez9M
K4zq+A/ocj8qycYb16tM4obbRA8W/6Fkow/3e3PKKe05sFfHgfKdkiAGC3YN7WQm
GKlmWfdNrPXhWfpfTodQy4ENZbSWhG1GZ1QfP23Elh6T1MifQyWdK9AWgdMmDb8y
nCMSMy/ofcXnL3/4JuLmGP3RhGy823dGYirVYQ4CqZvVN7SLrA2vEkxEgqDumgVV
mSqBlUt6aMWm+jij+5ldDp6nnsTD82p36WL3YUV/2boy3BCh9DgOwXSEVucGk/F8
A2BAC2oCGa+jjZbY/iAfsuMtTfGCgPbKcv7oWKhmEoAAF4M0mi/NGwm4n49FVaRv
qMShLI0wtKtQXAUyFtaL/wcAHmRKO4MwoTeYhRy3M7aUZ1x9PzeQxcckM8wkCYVi
EKkvcA5xjUXdsaeTwXasHzFsC54Y+oNUX8NPpIr6e6dlLTMyq29tXHhVlLuxqBQ8
fIxoERKLM22agsJt6fw0V+zXJOUj1+R2fNdXLUvDC5FOxNW/PPNeuIC07NMGxsMF
P3ggHIVGnpJRbJ9/Q7Sbze2DrgdW3PoZitftX0oC3MDd8wmR3aQO6H3jlUDonN0V
VRPM1YwrgyAqf+1M7aBtm+0tnhpyWZXzuVDLQyo2ufaaiPInwnKThCcBG4FHPbap
HXmYsRBhwHEMm/AvbLOIjnPhCgJVRGMUnJShzi/A8NLNytdp4izGQOs/XjoV/ORg
TZFTBbP+0+UcCniI+Psy/s4Xq4JdNTs6TLbky0X9sSP7M3/m1JBqFWnHAo3GLXNN
fuj253pdb3h3yVzHtCKl6mVdfk5911MyljNGnd3YUzYFxsRMhlimiiPuuSvMWb/M
7pZ4LRfcKj2anT5nYvJOib1msEYF+4F9OhK7D8fU0WvTzDg0CgkZPkg6U+LywBZC
SqzhmTORbrn7cYqzgXru55tr0zHUA7IVJAzaUOyw4uBWxVGdLtOdwzGEN6oX5oMv
itRrzQQQb9lAggmjPoEPOF87lxMTfy+w8b0nVI+1aMl91VMihU61ZMe4tIFr1BcI
EPitfTAv8Bb+xh89U+ObS/LU+jS3vecr5+GUbpkPqz+UAdVpjxdreBNXayQ2mccl
jibd7GuXl4DrZNbaCiGVJY89J1BPlRXswTecwumpvmjQedSmoUPO71LSMdoa0ih4
ohFgTJatJ8X4Zs8O+Yoalf+RpgBr+r6evXBtPrWvm3GuaVcqp5P7IdLt8wraBE8r
JLVLsWjuXwsE+aQmU1HIJRe8JiVGiUGKpk1tsxWDKMCPI2DXzfvx/6P/041sqHCv
93bSZELmkpRstDUbJ33p5XZoXJes97b/QINnKrmMVgeVT75qZkkOsoCW4d5aVc3V
lLPI8ihWdRRrl39hKdw2HFvZSiyIeqPJdjCSL2J6o8ngEw3yz2vk+W0EfzNYCQ3w
83FpIUG6lw1oyPGy1F6MHHUG9MUJzu+5OokS2NDi93KglEcXZOj5vRwgvgBUak41
DwJj/JK/H2X23D2IuGq6oZFrNfpKON2ICApat/A+8V/gbHK3Ej/Jkoiq/SE8icje
uz8rpBJJXxdpbsfKwEK2Hcy9zcv2l+0j2ME/7GFNBfhKf6PPjTf90P5juDNsy/Ww
qbI5LhCtm5Vp+OSDocbfIoo1bZXdK5FkMEayTD2wtyAboQfdYhjAQMrE5r0NgT64
s06itSV3ABZtoeu+Fg5IqhWTjRRRVTnPy7o47eYdfof0/MtLGXJPpnzsKZ4ehMVo
xwxjxMKNOxq2OxdH2wd4siNL6StQ0S6MGwCu/po/447H5p7iqMrCIaRk42OrjhlR
GiB/TBNk/94Naots5szcxx3+NM/YNxb0BdExCR0XZ9BFpX/wMy4vl5prHUqfFVb+
o7dOO6Vo02jod98fJqTgfBplMwJCG0blTdQDoADWMWOt1FgqNG1VGmejylAvTwmi
guR6keIZnPlZGNcUDexndXG3AaQASN6OwVOIdXkyHm03IFLD6fH3oshb7dzz/bd/
lUSTSEh1QrAo1eBrHbv8hsmlk8geLt7xMIBxzeOIiUYKO6g1GkNM8TFFL7nxnR8r
w8LMMO3VDwBvwOMkmm7B5/P8txIuYtJTHY8gq20VOMJIp1ILk+3FFBlzCCmSRgbP
VHpf1qhC2gw6OSWCRsHZAcOU6mJ3Nro/Pt2T6EfOC4T3k8wlnwI++6mlXUTgbNoh
8ckpVLifIx4NAJE7R7WqXXzXi3Jhaaxwuqf33llQxjhudpYO0nluFyyTRtFjJRLj
NH6o4VLREmuMGf/dZCiff87xPAXRgKEFD3iTeUQ9OKr9Oo/3T+S3A5h9wKy34ehK
iJUFJUmNZxUdsHmDxdQWL/x92mJSmEAh/uR0/3jKDZX/Esea22XAzsY+nBO7fFDU
72rkVGQJOdBsIc5dg4DdG6lxlH6bcA8PeH4NhkcStz2Y7rookhwChtIaVS5frKTE
s6RXQw8+dlY+/uKRRuhBzl2LdKc7x6/LhaZRfcWg+4nKXmWfq6fUOi7UGebYDwI0
Yy+FGFAZZEHDl/3CkZU7CkJVYTsCiBeDDAzrmZLgyfv3i5RNvQwpYYpA7Ku31tbv
2w+25cWtOw3aqzdXh2liIkkt/nIxspiLfrFO2wsS/Z4h7mjsOQqaQeB2Kl0B2bGL
FemO1MfGPjzToBN/m+iW/GuVutkODUyX3YKrP1BPbcZG49sNHpt/XrgkZRL4JxWw
w6nadEWanoZEi8O9BVVr64GxZK9l28i1hgGg3TPWY3xERf554qOwXgosGSmoGf2r
RChX7VyVVvBOnV1XNZi2aBs9pxc5+9/7rfsRFrqphTEIrjrdBSiEt2Ik0cz9u3O5
SBMyWdBObIuP2rgI/+iQsj8K0GH89mtjBKUMTOG7tREOXkI9B0U3c2Zuo4RgjaAJ
6QXTa56KiOwJNu3pIK60wIQ7lynMtKV0juXKMpwaeADkRTU/MtL5qKaPUdW42ZdN
ejNrlYrGngorBrNqUOJqVhZT/pzS4tbeJyHr5YZvxKNiHt9yJWvTMbWq1xHdBHS7
GB3izKPjivoL6eYZi4JSeQh/1ba5mrUETunvCJTYhsp1X6ghDZM2McC5l4Wyomrj
qxvJZmGp3lm3qdPsLFuLtG5W84N7VXiXbWo3QZvO6CugpLoiNanmLqWyyWYRFgj6
2fjuVqwAN6yZ8vJ2z1nc+OPyQV9NgCTMk8jmnh8SCrGj84/WbFdxtZq2gvP3nRzo
axQcGR/+BM+7U9tUYhF/TN2QgIJAK9/icpMq2jpt0WyKHc3QrNagtx5QEy5DauQ3
0Emfo9uqJBRJ0ecHL/zatNWVSmt6+QrO1yJhgoMr0nGB5T/R0OWayUKLoBLSMFuA
8eQ5uIUkbegqfylS5XLTqKhcxU6IyMemWzTJsaLZIfiAfSvoeTqLxov99U63fem8
vRvNA9cDyXoR/GSPWD6lIcBJ7dXWJec/AerWIjhIwiJQ+FDjcN+Y4UMCgnbD84df
nRK2jK/6ZxR6jw5gClBJ1/bIeejXsb9G1Cgguy66H8/ATMhkNGPmHujjuTQBCHHm
NZz+Zr5Kru+Fv5Gb3oqGhPeuqK5IR5EYp1nfUqochednJeQiXw0ijpY2v5QVt+cB
lNZZbfMFoUNMGtzWUwplA0hIqhWKdBnrzuN6OM2m2482fQjIWMQ74QJIAJ902cW5
4aZ7f58lQEhvX2/OwBE4bAwJXnCK7XZ6D7BLc8IslzQdj54WUxl19e9yAdUqMEHd
+VcmSXwl9SvwM4RwBDYIxHIkodW9xzIEiESDfqyTElSJOU6nJ9iTNKC+NsInlZiP
LktKF2KumSjQuy6ZLMEaHE5NWk6d3g0RBLV9gWMiNox/HPmqtEDeUJmscjHoas8n
m5pQWxCfqMziM4wGRmzOSHcmaPdFlOLuvKUuMDXI3GBSSJu4isrUZf2ZoVsmI3x8
MfzHm8eu5N/n2sQfTcrkeGoOgSiBh/GvIW85vGLJeCn6ACw1MQFeSSiYwgceXjWl
aUZ3NGZCFMZnBouOJED6JchDnZJC0qrAx1lyIEZ6iCwR2RQlHib+zJskf98iSB5D
akpoXvNJprmeFxPtrc7JU8EQsfj92doTQJwjshtFfvsImRSZDqLv7wNZVkTK1y4Y
WyjBOI9WfLpcaarajr1Oz6JKDHcULOc9hrCN3MNR17/uk5h6XIeIsQahe4oeWGfk
DGP18PSjrBh2/fPXUnUqwQ4QBT7H56l6gcmIEYr12bP5vY6xQ5yVknFRLgxEah/E
/2y1obTTdf6k0GhgI6br4Kpq1ldBLQqQhFnFjGxIS/+eKcxye0HEDHGeA0qEUYSC
6UoxGDVsvOj2WdwkxjWj8G+9h69cLUTqIzFFwU1eFRcT6Fdfm9cJHKVlhocRjiCC
Uh4HL8uyFdvlknLrHaUfnN6up4d9BxO/SNm6sHcaTEeJzCcH3Du4Z/wEQq8qMJ9Y
jF9H8dASGqKIV2Z7cC5hOG/ATwaJ1s5hf+gAoPKXl0wZmxcMlWMJxk+BGnIMf8B0
ulI1Q4cuZqSUXlm8iAql0eWCkcijvvaxRTukPqiHPfEevmlbEXP7qOWooT7vkQto
7TfphP++/T7qwSMsFGN9e/LjqNz4I5bI6ZoK/2DKKbGH4MtPHe2xYrU2IeggbRLN
zcVDHTQvhZolmMfgxAD46hc5ZKHFjyg4hPeLRe6pW3wN4lZw/Q6LUAK/KCH2jnRr
C5Wqt/tfaA+3676WZVIe4q0Aj4UulSqK1NWR+Ouw+D+vj71Ejluxhmr9QNhaJmML
a6+50+L4MqY4RmlIDKdiexFLjviRb7MDazedxiOjanuruUM49KlXnD5W4P7zgG7M
+2+T3hukXh0abhh21MSkRW6W492IojcyJxJtrFa9hCTb7otAmWpi9XlfzGArof+u
I2Vi2rC+w555ZVOI7TVTqF8SgWvYDkMPRZM+ZdGB5odMKB8xVmorxrgWwsyvEsDi
LPRTYJwzslZ5YLSkBz9Mks3kq1A+pUi209/zb6MPHFcvOTXVsyetz5qryf0KrSa0
FiYSD1gAmRGbN0pDELOLJ62S4e4Y+WkPBECrouad218H87vFWDqSHx8swIBJm4ud
plYf2Bk6rtLy9cAYfzFmkWBgvdNbL1+FfwAuYKOgSIxczvC3awrU2baDPlkk8ffY
5Mp71JB/tIBPlWhvW503Ueec1UyM4R6shCuNK0OjjqwlqzvpAcGzzC1NSgiLEczK
lR+abz5GrWU4is23s5UURTcBUj3bX5BA17FKQRkNyXiA5qhY8n6kKH94ytQws8/7
/uYAsqnkLXACwYJapk5ZssKxEF4np/U3oBYBGBcJV+ih+ChZUy0QTEkEVyLnU2X6
kEI0mUpz7BSipqV+gIzl8tyV/jET2LF+475grn6dgbLs6LmYYNaywnBT13jFuY6m
CYZmAbU1F0ap2dV1dFUPvR7/NXLSzTCBOqbC0+gy7mrW2RNfCLdF7r8rk6w2bATg
xgYEwMomMUQDeNceWOQ0gyv0zllwMZO+PCkgQwtGTA16RSuLwRi169oWIlJeidj3
J/pB5Xx/B+E0RNJinCCUcs5HzZk8Uq5Q8j3Lt6j9CQfL9HWn2QKBeznSTL1tzy8+
PP9QM8THNfTxnkTTSTNZf+01xgDGa+0tXX7fv7l72z6cxVeX92d3uKdkxDLWVm74
nC/FM/nD/adfnw0tZ45F/722/mVcPBZdkZQUmSJEx+gBcQF/NHk1WitAZtT1BqpJ
JIf/whZecH87x/H9MXuhaf0lNO4Eogtj4jRRs81aZRiPkG3NjF7nWEsy+6M8Gp8b
GGH8PFoxz6DnTOP7dO3irMCEZq17jVocP8j/l3/t2NxujoW2FwulD07pAQk2uCOY
2w8jD/fUtAETecy6vzM6kkCcgLNS9VsEGGJZ/G8kBq72gBtLGYz4+Qy1GA0YQQzl
pLHhK1eOdEBHhfq5+lpcopcnoWEUdmCcwONxIYVQZGJmH3W6oSQFZI0/U3B032oE
/aIp4dVkIQCmyvyrsfU7c9HcC/BkcDLAVu5TpIJdsPrABf/CWB5G45XOqjPJyQkJ
yRmOYFSvrBmElGADm4x3qGnknyWFsYWMmZBXPLvKm2h1SjTuDsmrcgqUKbzBiQix
MVoKjszWYSp5ddKdbNFqW6qeAiQIrMBU7jwXt0Kg9xN1xcYVxQkV+x5zaDvPoOkp
DQzirmx88B1Aa1Ri8ANQtRYReVjrOFeRa+/HZJiAKSoiXUge8auDxPek9+19eCwS
SeLWwParGXO/Nf8GkpLyP32zw3w90qZihalv2DE5a6PHLUBT/H6ehR979HtQkVSr
tKFgjCKP5cwarCcWSL3+x7jDRa1cLaJBa4WfFgdQcTSuA3V/Kevjb7yn/SHnoljd
A8ulD7K1KCwTLBoHVIedIOgaZw13DyjYpb9ucEwXyLw9NIe3mQQ9Lb/rXuymX5hM
Ta9/AQ2O1hn3/r6qy6+W6Qm5+A8xDJExqdmTc63/luc2avSDRMx9JTg6uP1IVuiU
odcy/nL4bGWwiQXvC3w/YGbTus15wSXbtJgyGn0AuEG7j52BNsDFEyLcJxRkIK27
eHGsJSmIPxeqXnpJn2B6LFcuzl+Fnn7ZmwEv7DhvNks1eJICsD+xDbQNAFgiq7Te
lZs0Spt6AB9QvprUg1PnxTjD2oqPL03PN8mMpl96/jT40oIvdyaKL6YYbwe4M3HO
VlNLwa4B2UfnzVoObs4sY+GDSdtZ6ChpMq74EFRegUuF1oTwvPHPoKqhNb0D7Ca7
H6MNPsbxtG58icVR5ZGaA5/QidXQQOzTua6JKvNOFuP6/waut5V/GJM/QPmPr1r6
40Dg1Oj4h6a82voG3Xr45LMxY599yeTkv6ja9KvU44kf/Tii3oabegeiT+3Jsnu6
pKTHEiMKuaWq6uLcC9gYycla8DgsD52h9PF2/0owp5zrnK/JMma73HQB/pZrA2+2
8eOBpwfLaVOLyRvW/gj1NnjqbTaxBt9Ka9jQxYcm5Qoid/k1AZoW9kQg4H1GAK/1
hcFuLzSRchE4Z2HowB2KbKG7MwK/0zkpFa+hCaZYAX6qFD22JQ90t0uCUf0Bu89j
itlsexMHQDDMNtvSFGhih6HRNfC33be/z8qstGp0Ko5DY3898xftRdl/+ZFGwEZI
9tx+mUOxlOUJ8MnFrxBiFkXBKGHeh0UYtGs3O2VVjPIODzgxWJYWK31ZReBQ1Nb8
QGuwEciktk6bgAPFDEFOlWLjG8mDs0HlqGZXAPnGMm0dwa3XBPGCv4opcEh8ez0i
61lZbwvZ80bdsNjhJkLTpN9jGfBz0cQ3ofnYKtDnJs9Yk2LyczjtIff12tI6moTO
LcaAv68vEALCiEjcXA5ToK4/2DDFTjabCFfSqM8BlY23FTSs3zi5LxEmncVNtxN5
5htSlnZ1MZD3RUocUJ73taF9c8W45/+zHp6u8gy2iIcffxQ1FgRJ/2omsR6URze+
TDEAetUiIubaptB26nCWluKr02+sQJRHtrdwny34kHQ5aS3DKPfJqtTWHK1EXGeb
GRKZUq3tDP7oYd/zuQP+o17EOZ3l5SutCHEN4N8ZuasdBLpwNoh+FhGFYQRSgwHo
2vug0FgKvjxeC1Qd1QGkQ+Bka1l0TCveOV7OUTFQUWYIO4UgC2T0pIJ+qoeSVndC
y8yg1e32PJF1DA5BXIxW3Q8QKWofK+QovP9VsQ0koJSWqjee9LOmYn1DUY4poJJH
LR31SGl15BlorsjsZgkfAk2+6oG/vrqRr4kNpLDPr+jwm3B6PbqzUuUYdRJAQy5X
z0YnzwE9KiP8hzWEZRbQ/izt+MGK2v1ggkQ+erSHuVqw2VprtZhiEkMB2JpXk9T3
WQ5WEojoe5h7kJoVKW233D05J0MhIkUUbCyTl9spyJmxZM5/n2Sm9Ckc8mpstQHP
BCk2PHXWmLQQ5Q+jUrNVO+HKHV9ljtnmPj8nbuOQGcjSEAJjeI83tOGZZzYJtXes
12HZMtJS9eWKUTN06mYVIWMFlpy+mYr1OSz1pMoxi3jBqQaWQWEhDJBwJ7mF9Iep
aTYSmmk4wHr/2mfxvn4TZLXYv5IaSO1ofUOqZf3I3A3/Y4aukf6E4/2OA+FWGeCf
lYvnPF6WaHMqm1jiNtaXa8ErqiI26VL+N4qxShrxJDOngM+9FiTlFRDeLS6BM4cd
+8O8Y21HWCiO6LNIuYt14a6LrXqeSB7mokUakqCJ25VI/r5B4PnTGaYSgMsQJ3Bu
8JAao1Mf5CXudQOSE/uwdMD/N9jFgxLifxLd7pXB+BXOQHvkfMSjLPAMzZj7ra1O
akDLAIoTiz8eMFgP1AJfdbkCiSHpcTLlPiIwGRdVyi2aadFjQgPlbI80RoIbPXTs
B32jSOCXHhblLrTmFhgYoBX5mZTGFGR34XLuCVQkS1DC18PmaEcL3IwHs72F6qF/
2YKumDgdCKsFuWYlLM/Fx/DNxC7vLkdGzRtyT9K/mMIaKEE4g74K90l92cpup1Z3
P4WNhz5EK3LeqZefK32deTWNtCXzQ2vzFBbB5h8gzkmWItBnQpCONOeDq7tufnlO
qPWJ4PL0mbzgKSBGzUKunWjMVF/9+tp8oGd23emRE127TuzxYUHN0nrJL11LHu1p
wo3xhpX+MGF/nKxj57u5moxPqAxZ7chEAo66wTlcKO5cIze+phqTK7EXyPHFkdlo
feIpfQhNs1oZ70fsxVkFZzlxR6RBxDaDnVqIGRRDKkvoK6F6tsDWIk7wQzz+27mj
9RrGAl9YxDAOJ5IW4wwDBYMNQboazdcXftW4gpVe4S7FjnhaEhB9ZR0n5cWUCdaB
cGB5B7rarDRL4M+NjZEZVAygWGciCCVlIQIoCVR19DkG40S4svm/nMq6DYMl5i6n
4UqzNyp7kBkZxiALtuEir2DpE6Lw/20ngt6Aes488X9RZeCEBVuTinbXFk05DLpF
MeqkjdP6ILA/GHYJI3fwH6a5sHHbqdmBX/3O/XFX7T2Zg/zL+RroBlxNXiqpb2Tc
KKpcPxAOrQkWRTkEtaOP9kULr8XQPkvYmy6yUgQr097/PXs2ygbW2AJ9xlxtYx4T
Rxd5b425Ev9GUQ6IrPZsBQU0tJ1aGQAhRUpDNjPNFi1lGcDLqnzCSzXsSlnW8XI0
RIP0mWaummKVC2Fg8pU31G/PM5SDL/9Dt0QXRxuBKqSteNN7b2QYPgWqDPbYW8ox
yzjB3ld8FV99dwwXkz1seeGd6rAtqOsuUAHUS2G9T7HokTPkIFNVS4QmOvJAcQWX
VvogSPejY0qjjQ7mF49oTtfiUCpODuIBP8EopOeL8LZ3ZdyFzySlJC9GCgd86ht5
gvCHZXAZbhy0xQDfSmvwt+O4MlrXjyy9tLrpwI95kvYmPlAQS0bKgo+v5B2RPUUl
OaJCeHlLQK8mIpB7KFXyW88z0ugmUfjJ/P4y6jZNwo1l1AX8nt3/EDDXn2D+Vkvz
sn0x5Asl2BWgulzoRh5qW5sQ+gUKNRZAKl9eHEnFny1TNGlrPl/wuKX6o8AUIS2o
i0aYdHoNQLydBDYX/04cBhk+yVU8m5PIDvYuqp/1dScdrVncyQ4iS0gw0V62AQvB
s6cXCaDXUwjeJUSF9akUUFzmU1z+Uq7LcDR8qApA0Oa3Lotb0T43NNrHArG4v5LT
zlONUIgE4Os8H0j9imze2b48mqWpHZKUNsFQkHbI/hEFc1eiFiZWVckqvgRoOmcH
n/AHZNUYCL3DRFFsgRXs64TlDhXqpy3f3cZUFIzbF89gOOKH9XauzI9ZqfSpIRit
yBTLOfBdrd6U6AYMgx5eI1EwtcFW1EM9+y4HkFPgzy3kzjn4VaYGFuMzwGsDExz6
wkJgPhKfZmkyk6CTRz4WIbOFh100HQjOy7G6srqpmCkNrQzs9vGSKhIye7nhT8Jh
FJj68lJ+J64p3huKi2rY9AcTv53Nk5HpN85OqJWVtKqNkio4Sk2jUAYubsFAyLqG
9b1nJeInhB+SaWlK0Fq0k0i+iN1ZWDQzq25SNQ6oasiqd3qIBLf2UKN7xiNfDrbV
7DO8zbjrDscZKoZ4ah0OFiImgFwRBRqV9a96pnXFI9rwWh8u2akXYTtg/FuW/U5g
SHN5DJNyFgxVLesrkU4ofqpAf7CPGqlAhM9Uygpv5Z53RVltlzr9EV2QoJEu+jSN
ZPphvLlU7rnv2Qrqaz7j5YRcT+JdReoIoOkKmErMnUxKwxQYjjQXcz5iqz2UEDQx
rBrF91nPTKVpIGbSvDf3kOSWnvweCSMotJSkbqhy5I/DFOYLC9FBmcVe4wJ/AyU4
svyyvsn9Vg2tTgdY/glGYeA+p0FiRVRyPi3MqdtMc99eds0kC92RMED4lgHLZHxl
WFz1iVTQK9Bamh1X3vqIFCBphrXtgxnq/G1xgk617pX1K2ZCKVoDk48cUqX+Ba7f
WCi25ROCYJ3WdrbzUD6j3g+zSU9j3Gl6bIjnAt+g8zjSh1u2j9tXVV/+bxZSteN0
ZsgN9jksMll4SWWxObS77OeY/0GQAyzzCTSAYG22h1vVY7Ny/XS1LQLT0TCPvqcF
I/cO4QLJGZDlLDNxVakiNiWfxpU7r2k9KPlW2cyc+Gqe001uPOC992T0FKAkFqNW
hcKs72B8lAf46Sule3rUAKif9fmORisJyaroPp7W3Q9uL0fLM6RroSrkthAWAkrZ
i+kOZQ66nGRYJIqsTfQBjYjCxgv2p/60l38QQAhXw+Nv99OqoEdYioL6rpW8nOHX
o2ioukOh0KJcd7O1KjvRLSPqe9RViw5UMseZ/9tt57eWfmG978U/I9hWD6j3PF9p
Z1Ynm8NXu5yAWH+/Nzh7WSag2wNci/lqJdAprusSkyKxAftDwFe26qnAG2v55W/B
dolM7o6eu0l2qFjv1YDnnhwDV64gePonLW9l8gTGBGUg4ZojYrRVWJT5E2Wv2A47
RhByAqHM5AQ9j4W5jBf2p4fCK6MN8cBiTdRW4uE3l1nCk1jg2UdelzUKeefR8Z2E
q7IaLfF/TrsFxjcwv5UBDSeiZEuYaXTTj8rkwYecy3DHJDdFyKZCCz/Jysz2oKQy
3QPcvtKQY7yxYA4qH3LTaNG8/ejFPeMed/cjDaoEk09AjIOPpqgAWxyC3eWLbUBt
pYjVcY7L9Jo6U0CeMwPeTVD/t6/X1FoZgiEO0sb0U804mcMbYY3ulIROWhoiek/L
HYx26zE1ldwsbvJ2UtwNfKugcLKnFg/w0Ya1TO+EvJA4/sc8r0QLOSC3nSeE1EFD
+1dyg2wtxHfB1g0bphXLNP+UWpP8B8qGGYjF/UgM5jZR/1vpbNaLQhxqV6MJ2who
qE/E5iZtzeP1EZ/IgjCkOn1JDc4G1sOFbS5IXy0pz1oh9aYjNDNrgoQSX7/PQfjL
2bdV7tEZ6WMZeo+XiI/KsmiqoPLnSd4qwlOSRadoOz/G8u5snwMLOooWF5iGtTx0
ST419hB0Iib3RT/tbcBLz8MboPMpDoFi0Bnni+gq2OuE2mJ/vcn0PRSNMODGWImP
tJuBXoTEZw8AvfmtI7ADVlGyf8uNaV5R5sr2uQ557WPoROuzRtuHA5oJbiRwYf+E
Dtpa1H+E6VQ95/4ID2JIAQDeBrH1UQqfRX7jcacduMh4Uaie9Tyb4PLKJkvcOWO9
Co96ERHhskIVLpm6KNbgVb1pb5zHYIZ4r+r4VvSB/xpMhMx4kFVEay+Y3h3PHmeU
t8iPbNdOP3ye1Ij7QRLj7LLHjwTzB2J03lJbE0r4ZmTMYOi7nT9ZRDHV0iGk9x3w
D1hBR1BmCiKB1eC40SD0hBWEbozGLu6B+4OuZNJQKix1szCiVKJjurX3IXE7GjKe
WZa0AerbAImbRUWSY4dQ3gQGYqKH80A8pQlPGlyW7q9bFHZim4epT3DS06oY54rw
kGlbCXamCki6Qc80H7d62KxqtfYDiKnl4pCr2mslDpseJryjoPbz2gC8kP4wdsoh
kjHLAKirC/NFCRUapHFyOcP3GK+QJaJrL8uJUfCm3YqOvLs78liZZawlUl04JjiE
u9WOLMfvrCZduPEJMyFhg7FkBbBhFkShosDlPE3303yeAB+8GIjHWDP43EknmFVB
aKyJGC+nPIPz4qrgzqZit5W7IN5lmCTPX61lKsBaYs/HfdTe7UsEcyu0UqyE37hK
p+YL0CUj7DstXjGYzZzHHEOinhb3E1OXKvVEduBHj/SZqucWBQXPTk1Oskx741o8
GuvL9CNOgKjnSa0XTvTvgVHG4/MEDeGkRDmq/BRG/PBPwW3SFGJkulZwY2uLnlPf
/VVOKsQl5by/K8F+Z28JcDG42da8hqp/Fw1X/tcqgfCd63sbD9BYP//BuNLl3jrx
3W3EzZ65bP0WfptRJMnDYbRV0viRlIvgsmoQ/clVEzUBi7vWwE6r31OLb+f4Qs6q
Pbs9PbXTv7A0TmvNVQ6G7HhrXmS+sXCPTAuHKlzWfRCBWHSXuctTdhWOu3f+mgfC
DQn0NY4ryGhSxTkq4aBVd1BLw4IhTGDZbd223zcWhbuuvmTL4CRGXq6QY3Yxd19r
4OQ7uo86Z4sx2QoI9X+uoEEc06MDP7XWsw5ZyG9Pvjzti1L+ZlRx+JUyIyt9GCGo
oqTDPxn6kqbtb9B1I/gZ3OyvSaL78AiFpLruTE83JZn8hHi/Y6+K7OXoxi5erfnT
b1J0K+QHTQ9W1cTTnensRbTkD07/tH69eluMNATyRSdgJ+0bmLzdjavBFWJLn0uo
64cNbJrzHjY6iXtf+lVNvIKklwmxzFEh1GCY8Ct8te0B64zepX+DqWoeZczS99Na
Sx1g2WkXWo3Xlf5tkYgWG+ZO0/wzPzLjCAmxaUx9B08FercWnw0eLWixc9ABSdDG
/c2TMWyg4ctSluwsjAwTRrRMTMqxx5NA6fcrBpL8THuwq/+QKNwr7PhiRQyEI7w4
VufQ0xW1ML9eSR/haTl0DIuIWv23cKhw3N4KJQ/twvV6LHahtg+Wsw+ZecM2L6uv
ikt9BhkoD3eLsDVjwGIwr/2s2gcdw2jLz6Al8l/rdZEZOnp49P7ZcQ+nY/tvTBzy
ilTvt8W8Sncj6X1JWeRnRDCvb6u90vfLSOwCXXlFUjAcXRWs9H01OcZ1ov3TJaSi
e16vPNtW30iDUIV/nYc2H0pFX5TGUk5OPHgK0Fo/4jKmjmJSn+pLe/Pozy5sqg8u
QcJDJiw9Lx+7X82JbWUoTHtLbRA0RSrPVuZnt/z9+YJzOuc+Z7zMcpmtGxf06HJa
oOSmTSmOOBfNzgmUj84Ko8R/ll8xC8McKiAMHmjaVviKm64vIpGDLnkgLA710LVf
WKfzuLuIILB5vZ5AdmGOlbqS7fbCHgee3FL21UptTp/QyIMdhhfnYKor7jBwveMV
Z7+w9ifs1wJ35ESrcvZCiuErkG+fI1ER+OdK+vxMFfAoL9j8ZQphebDeVVDsPAEH
wWk8NHCqXZZWDJG02uZIZUCEBl6hxCdNQ3xZ12yVkjMAQKobcHf1EAAxgSD/mXXs
1r3fiFLuNLkeMqDmdkuzpAQ7uZKLD6RiACyI4VHhoa7rZjll2NEDl39El2ftUBsP
+1HXe4S8+PcWgGVzvcXUXZTeUUVDriFQ5TknSrHK0YcBauMpRqW/HaOHYWpzl89K
XuXhh6IXfsGsN6LAGt/pdOjiVekyzqjbPkOQqH5bANhUtgXI4bDKVbz9Z7kEUqHT
3U2IMxICF6p5dAH9aHctRCEojuNqivZ8IX3FYrGOEJp+eNoQzKiA9eLqXlFWSVrO
6xT4aMiBlb0O9mwIkmdRliNso2AmsCn50T5nciFn66lxTmPXINBb1ymPFp1Eu8KL
Uu6SmVMKGcE7O954qefHG1Rlpqp1zq7kS5LarkHa23bDesYReQIPm+8nKVKjpvvw
vePSZgxtBP76OsHyUQa65UtXk3ON1zX+L7R7u5aTkrW9z/afrDXUi9M91v2LfHIc
QDmkdtW8F0lnggeXPDli74tznAshFw5X4XP9OaRPCTNhSPRDwzS4Ng9WjRkhrj7w
F0SYudgtrCgGwYQjtf5ieHTHKCawYnMVi3Wc6xUosmKbnv7iTxeT4anUJKrarg08
Pz8PbTH9EuvM9p1NYS38LfvaTxN4lqcvz8pTDlOCQaK0DXaqj23U4F4BZwaueVEC
rxsrrU+VFgffZlwA4Z5r3Mp7gZdrdyghf19QfpHkmLv220w4BNej5By/tyYZIaHx
lQWG21F7PPrM0r7gz15QrRKDuSoJ/1Grg33xr3cy+V/r6a/sNfzeLjYMmyzRKUgW
aqUjd0VqI4kZ/V6NNlLesvJEhm9duBu9ABGMEGBbMHXB5SPp45D3L4e3wmDnbxbP
nVbRJ6k+Oaf3sKNc8rVlQeygEek6Rp8Jx4WqnkJ4TNPCZ/OaJGH2RiPjRI5bif0Q
PV+W/rW67gD7UxZakgT/TVkizgppBNmYm6u382cdKdCuKUs2GEVn0pHrzJhEVGCz
IGibfF0Vg23is7qf9tkDukx4mzdnUPRsYlHBJK8ra0aM//OXPEcRLGOB1oRAg922
NCfIe20rRc1c1XHwx73mPUvXaoaZk/TOx4HL7b3xGdYGTpEcTtb1+z36P88iIKVC
N1yzVmGrKrShuERz3oClIYIpDq0a+GUsBWmqYqBBIS5NIz8NfJDbkXfjkOL7gQoN
m3IJPUK3tp3Jji8ufc9w8+mffw5KjHUrtyMk/A6AAYSlXtXQmNmzqdxk2pZk8eGd
rAXQ6SECRgs23PydoqyXIEzRc1U/GSDTb/nBufO78pEWiAJPW2pjQjp52vy7UDV7
UaSaCRdcrPEtlcj5R6e6STw6bhRw361o8ibMzt+3VpHTGk0gpClF4HybqovBWBBJ
jKsUQUajnEH7OpFYXKBWnoueaCDAybwlSTOtizSulihwE0cG9Mc71b5e/WYKHuUl
cFH46G98cjL2NN9L1pCFvjYgsiPX42o44qj93v/mGxeYMSDAECrOIk6WyvyBgiF/
Pzzso5/8Jkde9wfc+VHq9UnzA3/5GNinf2jgtq+OLtaQZrRLabfUn8VPJzRTTHbR
H9X7gG1EKDZZXsrY7ofiq8ecOTtJICDDyc3M7PO6QV6LiLUFQyyAZ4UYBW3liQJ9
1NY3fBbduGNiQ7BtPdmaGt/koSq1O0W44wKceSWntTwFHjh6KuhG+ilysyEEP6vc
uFjKPSJlyxjJeWPbD57UIJY4cjzKuxtQZH3fNVkQjaHcA77nSU8l7EE1dxxAIb36
B16MOK+cJOiOfcAmskjGb/6uE0aCxMxcPjPvzD9MQL5ySRpmxS1/h5UMpmxCpMz2
uCs49Aw3tDd4FWQUNAeyEAZPR71MlRB7Q9CvCZiqBN8PMTZc8kS2uHZZ9leZr0c4
IbRgczymbrLIZi3fiL8Sv7Qg0RE5SvFodh3QHNWo92pjqamrekDC9BHICREtj+KI
9qWnlW9Vzl+mGiACUOlFrs1FwXLXZg8KlIPcPQbRMZ8MMmWzndRIWsU8/t+Ifdts
3hcPv5eJGWB8mtwsy2ytUdqAcSARxYIIu10+9wl2YM2GYQGkFXvbcBQVNNFzVvFl
CCBd35NuSb5gHiJNokHzpbxPh9GS2hyBHC6jP1SWefTpsgh1yhA+RBGriN2/9kEl
DplSjbEf3gHpiWEbZEDLU16PhMQ0edYZJPOTbCcycCkXNK2mhAUJnnhdUpEbDguj
AGDBkrGDO6V6rLbfcOdDjubSE+ZytfBEJUeIUNj9XXpp/+Lsi5Uc4oY90kiXOCDf
dLghGE2cVcWpGF0Mkr7Wd1sPBvIn1X43KEQDV1zpVKjSb01DAatyAELBBAUe3jNQ
Au64rtrCdYkor9Vq/5l/Afm6Mv60JAsBg48uH02JpGd+o9j9JQ2A88QFLU4jB3O0
FJDZtO4hx2hLIFSskRNBz9TNyCWEuX/cUJGNOSjbelYz2fDlKj3BgOkyGEd7w/Qi
aiJn2AiQd+G0h5wuKEUajSKH9z/hJn0oBNqHaaBFWKHBWmoQb1lDV5lzdLRu9l5p
9gGtEkL+L8H++WfAPIxg7AhRkbaLFHJTLRUJsNILurH8VZX6ba93i4sq2rcvpaWt
/q/oaJtTDHLfiDbVv+APft2tX6r7/Dpl4ezQsBBpKAAbxkVBN1Ldp2mCcWUIQICh
AZXcuY0MI7gb6UDFpyUYlXegnC/GLm5tmX1K5buoGt2Ge6jLd/ghdblCx3td3dR7
nDarhN53cH7jOvqpQSWPxmjK9fmcj1Mg0rgdyd6HvQ5gwRChPo2vr1u0SubzOQiE
SPt0V8SyjIJc4gFpMh5tPaT5KjY3jQOv5wAUOLVLlYVF84DzCpP8Es/Y9VXPhJ5M
9ZPFXz2w4PQlWsK+0uEd2aCURNkNYqWhZYIyqAEEip2f8tAyEcA682e9xYylM8I6
Yf9xhk9IU3LMg4K07mb0yOGl64HVsTAv+5wL++E8ZDwd/pwDJZGkY4r/tZYFtXAP
6FcRBInaDph36djuCYiTYuYD9cThcZgB8cORlUTXAKyZPqKAoZOyf0Wlygwb4hoO
7064xjXNvecWPkcYhucjIlQvyRWbda6ePL+/3xllv0jr8RreKPxxRXTXZuXWqaN3
y9x733qko/tiSJDGzuF4NeKL9TrA4suiuJJYFIFHRPMmFyhPRYOlXO5pKJSYsiw1
V6u8OetTuP5oXDzw6rPwCSK4TxNhd7JIxGU992Zc1D17Lmja1tPDBu0gD22P5bGG
5sbBpEaEB4owf68Nt85f/49IXM179zsJ6hXR1DNi3DvRkJKCg/7xXDnY/PGn2P0L
4iT7lFprbGHJvhabDyvSqsmlXvPQKmefjbRMCU21xgAErdpH6F2nV9vqvvvATod/
9EGbS3fe+2oRI6PMHHaBDhv59SeSBS3E6DTXZn/AHNXFEUbJLeS7NOqBX78zi+47
lRhiVZyxu3yeNdRm0Bj5aBVvKc1Jy6/aVcNGm1xsKEzl66DTO+MyZT3ykEr8rcqC
SgbRrOo3USs/YrB3+9UvfoElGCd4U2AnbtRBIEZuYK+8RzhutAvWPut8I63UtHeM
oc4ZU4j5oN9LtJDghr7Le2yCZNBuc/ItsTs6kLmWL8IwSp2NWRNsP05VO/iPdsA2
FgytX+Vma1IG2ekBbo/FF6y/UAh9AEK3FH5y0fgoyIUKiKXXFQe3U/uZQFiBe0Qs
fzemiSPf+svYA7m3qZyKMuAnFbEHuDJaYp1v8PUqrJdqz+Mih6v1m19RWzsmBY1m
ODSMqTJ5XhJvnDIQmpxWg0upVMIUmGkL/q7pTdeX265VD3VbS6c3eteSvo/9nOVX
uSstvkOTTFoyBQ0QPZvjTQL18k1wk03rgnSe80amMhYLbh/4fCZQCsdNvxY378Wg
B6/C9ryDNzirN6dvL85GvIJXkBLHWut4b9K7sT9rrcX1pYQMFox1llIhGM5WGju4
7VWPSqZbdYbcT4fRFmUt9N93dk4tKxzFlmewwvwknsHNklOOGVt997eqAMpzZW0h
J+tvjMM3Qcoit/yP2iV4ZEAg7zV7nm2g4WGiZ35UjSode/5bfpbeaSFt29BdK++i
gZExJF5+DG6f+vf+7XIHjJJDiRAy8nIpnVyDABaCfTuI1aGXPqeZV5hwzYl2AREZ
VH/pKtAeCDGSH37C5ZLRnaYoL86tV/ewI3yfGgln+l4qtHCa4d1g6Kikb1crf45b
4xtCukOK6LvdjnNKFJ1wKbfhU8sSAtuoPG7csnqoTPOOnfkA7mkmnOfhJl5fh/hK
vf7k1OXeF1ImFr1FYIEBdKrFy8gc4KSLiA+l3phS9WT2Nm19RyQpjK0bhVraE3Nw
hO945fg+It+y2EZwIvVhojaJbCXaeN5H23G/lAHQdvcCEgLdBVyTLM6qEVmG/m0I
X2Jrxk2oW2F853SwF8sVlNaTK43A1h/RDGdS4TCoGAqEKq4fknV9Db0LfQTESUR0
4KjLziMSp5XMJgXuiY//G1DTs5gCXS3EYEZQT45JFjfUjzr7KSWb/A0AGJPIFRtV
4wTNXz9TWaxAPAIvU1fztSv4GuxJ7g773oIFjM+LGpZFtKL6+53PUo2YJjK0NB9Q
DplgU0BEdW6zTcDyOdPFNmCoKLrnkt96+Gnv6z7UFwJScaJBEe0P1R2l1PBPWVOL
X/RJrKABYEQfm7vGnHDklb4ePqPQ1ZWhzk+aAHsv3Ocw0V5szJRXgROt/QJuaw7H
RQ6R03NN3gciKxGnxfZo01CYXJyI2wvcFtOR6/SrFcYFp1Txwo/ZZ3Xlm5vJeb3I
4kj+FqYsp1YcvJDi9Xu5/yd8Y5vWbAr2dDd+aq60vFEzWEpWUJa/F/0tWqtUEdOC
bJPdh64dhmf35cI58tUTBnQwZ9/VcNl/MPgYVACEuAyAdYzMDnmmoZhOTZ4RT+Cg
etawJ5gLbweptsJeOnDXnGFocmxLRRGCzc4LtOd1sYy2bemQVMDfbMYzR6GILhXE
8CNgy1i3FL8VFf5qouqGWNRNAhckYL0ohf4id/X2NIriLq8wpkoxZOMmoWg5O9N5
PRG+QvmugMlcB/IyY1ZRI4g09YM4l2clXcNxwGaqaLTeWFKlPGwLcVlF1edFuk+6
//YR8cuCSV/6o63h1wAhNb6/i5+3/Hd7y72suba/yoRfHMzLT7LjLlugybXpd14H
hjM01bA9b0s7penWGK1IVm6zt07USF1tOvc9T803L4z905YKN11kRF3b6Cb5Z8ki
nNcVUmOXq/0537fOZcr1I/7mC6R5qC3Y0tpNYoV+TQvTsrli+OqD4sLeYyqYHJTe
Qs3mqqbCw5r77DBdz4nFt//tac9kVXDhsp/mrKe9e25FDDkjAN/xBmI9F5QbjQtt
wDfxZuFHN8D/8jp1mwS9yFZ2Mwq1MyqcexkiHLHHF9JyKcrjHUQ/+wxIYSoLPvgj
bNQ/phvqc/XGZ7jJguuDFV76vpsRSOgDhgmNmjlM6bJNMBMqOFobeDzcrZL586r/
E3IR4RFguTQ5eBk/K4eKv9BdtqjtnSX78O1PD0BAIM7P31tMsIyUPsOKqTyWWh+x
+h1kE+o7O1LRhAHHVzg8EDzM6d96tbjc7MQF3sY+dSEsMNj6Ev1HHOyStjJUPUQV
XWydKm/JpAnh9iGTOfCRYyMWZPIatbZ+hLEd6IKeIsP3MvjdnPgxQXaKDnsc5lQC
w4t+8+en8e9U80W7pvTPyh5iXqe+A+EGjk/JL9W+42l5TJsvag3HIBfF/FjD2Zts
i69MgbN00BaNaUnjaco0XHIMjGWbWCE6CNmtollu4GuAR1olaTVMB9EkNXOxPKR4
AhohBuRVv/WGMCDZgz3sS7jfxKU83ugB5b9bN4j4bR1Fwce+ZR1iilW6/ZpsoehY
pEp00grJfN8v7nshEEynYNwjt3wvhnmxxWojyj9cgVCBxlTLRzADoJNk8R8ixJgx
nKjrjYK/PlAWauI6jCtrhzUlyMzGq9jxb5vJ5Zjs1c4QL9keZNcI+BhxyaE7UwYy
T8Blo70pT6skj7QvK/vrr2cggw4b9KE0AZePuRkygSiWtou8mTMs5o63qQH9VxZO
SJXi/jS14SmVOlMaOVH5PqyaPld0vqnAx59UW+MPNHkT5BDGJem7gp7fLxTDT2ct
V+HHWZH+fkQTQX4gsJ1CfYBLuZUJrBG/YhtlXfxOIrqP569pMAjoNmY5hg11BSpf
AsisVXrc4YHJjqt3k2FyKxu/BxNlLoi/jvWihiII7z1luAc0zwTW7RE035tgUmoW
g4ih0PqH14IMQfGrVa6qFm8/YlekT1Ro0pxdtJewq2hczYvu0QJvVuKH2M3FQiVu
uDSLktRicZFlj0lGLLFB4TpLfeLTdzezc56bx/0N7+9KvrZxt63uPAk8umYAT+iH
LEJga1fohDGdAaLXYU+T6iO5VYVY9PHlqmOxf8n1MoYhJ14gMlL27BZFKxoJu9xh
uoUWmK2HTayOGrarnmE8WOlmOiqQNe54QOjlFIEO2BrJ5dxVfENM2Dzh2xMjccxR
dQHKUnc+DecvLuv+aZevxf/fRRPCWZVgEDlx+aN/+Si4OXzrBWED1l3cTBtUq+Nz
PxpfUFiAPvJjpo8pKyacGlAkNIC45ZGjsduaWUFp1JvAbXW1y35dDqWhafx5PgTm
r94XJ1STD7jpYVmFvJFSZPmdSVY2fv1lqVaBPD3/LPEr59huWI4dKNdTx8utcmpM
RdZyL0CYBiko5CyEDxqATwGxBBaNOsmS6livtgVaREIEO/wxgR5I/PVmRQ8zXRtz
plprU89W8i93EmzmLwNVsQAd0Z3TJ3D0nYzoW+8aJ0F27Yimpxewd0IoiKsYItPg
Aft1CG/fNdeVR6hGG0wK6PY/8O9qo90FFgQZMxDoZcomUv4A6BOWhkdM9FsDcjOg
eKkdeHACBfNbE/tcbUG102DMhAp2AjL17Y2i3WSJane0vJjl/+VkAcYE4JdxTUxE
VFVNo6i4QY+opnHkZdjriohh0BnlTXlcbSZY5aihGSJQiLddE7PZAanLsYtma64f
0kbT2/QXrogOqiYgdIr+R9JDYjpbDAIm3+rWX0pEdbLOytAojDRdFKvQp0+WxvBp
iE/zEq+GnhMCveyZC345N8J+cdCc8ls3CQj7z00T8buN5H6p7AJ105Jyb3uzgw58
VwwntnXRPhM9lUaKMy/XKNfkHl9W5tCqBH4WriVp1zIbaJt7F4jilm96DJnFBaIc
WanqMwO49zmsokRwBr5Xi6/6FAdtryQIHgjdWn8kxl5tPplpOyHjNdexjM5RLP1k
RzlAXlPD1Do80vNZWDBcf1JlGVI2OXtkStdP9eijBldh6o8gIqhL9Y3oqQtbHue6
IpzXtb3tUIdRMjJaqnj4gqjyiUm0KwmpE/3IjvAY5iOOlzdZsace78AxFznv7CAd
2hEYrOCQwC4xGqtM0/X/0etOYmvE75nP3gfoAxLKRU7j+NUEUS5zwBGvwngVwJcT
kBvfcJBr3rX7MlvEO1LYH4ZXwboxKGrdKvXnlyNFunOsnvXX9zPpwGO+D5amX8LV
+9bNdDpg5jj2IdvpwXRNrt88l/uL7Mi14ilY6on4WsHKVnkiOOR+TRvB1gi+dtBt
MB7gJLhEsvJgAno9JtC/rESCsMILKbUDBDNrtu/zfGph0YA+UjK254Nd+6uYOuGH
411uDt2wEzsFM6zXqPsnSvMNhBxiZqJHTm8V55SIraexjhr0IE7rLeB22DIDe0HN
vTa6aaqTB2MFog5Xwz/WxuhydVIUd7Ifhp5A1yJFtXi0hJdFyfVVMhUbeIvyCm6s
ypM9JkaCCXU+LwXDFdoYib13JhDlbh/bXi6BlQ+i/gaF0cTkBg/0huaCpA56gTTl
iRhR6dMZ6IIue9VOizI3SyvmW/y8q6H7PWcUK+OzJlY3bNAJ2XB08PSFQM9PFfWP
w8Xi/nzYufa4MaB+KH12kI0XW/+0psAXUokXEho4q/SLxosMlEzWK+twxGgE+fRA
TFYNZ+OSlt5s3v3G0Mi0G88lFDG+xGaSXkVirOWv+uid2mk8ZlqGpxqlBCeJFSf9
aC+5WmECBU3a+GPgxYB1rQKTqX+sdIDMDQyB26N5661BzbT7bW1JTdnJONPdfFXX
mhDRHpBlnPzaBSixUU6ZRZyqvr9MFM640R1cPNh6yPDgbzMApSHY0X7SKNiIK4Ay
RIP3iKDlMzKTBnnXUmHVOUB9HIWcODFNIL4tdtTNuV6qr76sl6Dcf9W6r4/f6ZPp
rU/8yVfubHXZNpCp/2EEWCka8/eiTd+5+pL+NqBD+Sl5q04XfNqqEM/Ew/KB9nbC
NHPWFLgwr5lEp1dM7NF+o5GHD38+FKwIvdncGWAvbMHVot5dvZft9lvnWqpRYH8I
4nnJSMKUCCN1EPMww43TaJcROuUPW8WH0h0xuZVlQF08IuTcv/VQ95qMUrkzfWeg
hug24oYvdb3W8laghYN7VCzkxHlI+YCY+T959KO6cAeZcOjvd6rt2OcHhaQRcgak
yHdHPfjweuNVFL+3LXvv3yNSiTDhU2zqmUi44aPXIEvJ0gHrtrh56bBIGMsUYAlc
AjRc7e3LCZPClC73ik4HrhbqvXVojWV6rbn3WX+66uPVM4CXX2/47YcHkq73LVIf
0pRPnPjP5hK/PU6A/QfxWhjljNl8ThwHNxOuDJ19N3+xN1gM1rU4sAIXofZ6jw2J
+8YtAoilRzdR9Qddmf3Q+/rU+1dTYk0yj+3Pufah8HOGxV3ipqDAFxD20ajiAALj
iWqYL/Z/DkWYG6DqeE/+fwV1uhXU0O5MS/LQNZ/zThShi444/6C5aZIvDA+trYHR
niAkNwXHT+EC0ct8iy5zV3UDdZl5cHPYNQZMaJ8TTeKAn5PaZhyDhBtkN4UpERu9
HWvYrOY8xWFAI0jiRhLQQpW0U+1Zsp7bOrEoZd+e75GtXU10qQLYa5iPIHMRDWH+
o1Y/CiNK8SUHunTmDqImuCkWfqyPUgPty3t3rvsRODzooxg8DubDBcfJHztS+PE2
BrQ27xAm/8cG5OLxqBX7RADkvkvc6wBMTRUR50nc+RPX6nftmNuLXroZOiEQeLis
/2ARj53Q8LGKLX1nohLFBMPlkYNm/gfccK0+AR6osBLkta7ZivDpNtkiIuEZW8z2
jHALGv/73OzagAB/wUxyx7aZ3Gz13aIsCMD5n0mLNbMJWXrT2V9WVdLDvMKIBtj8
V4V4zJkYxhFZN/WJCt7iHeG1c253ltu4Lki80IGPP2g3otbZrIxqu7EVBvAL0ESr
q0kvi3mNKKyFt3LN5e93ZUR+4w9pCWYrerha4hnyZFJwfqLzztv5WQtHegXxVg9h
sfAdloAet0NZElX3MsGobnp7HGEKxvPnplBrGj8XKaShvRwW+j/Z1oObFXDe6GiD
A7alKZurDASq2WHqNP3HNevK8Um6s8Z/uT0f8mP2GLzEEENkVw+3THWpojGh7OZ7
8ISSZGefdeCSYeG2LaL5sgQWtZOb4RP3OcDQXz9dFlRnU9qRkz2MJOovAqwRpdS0
SPlflU7EC8lI2/yKoITlkjNoY/uXrKh3n+9nbTEOgs6E0ycrRV5DEQiyiwVDYP06
VLkQx1jJpNNa0LAcpgHsoJmGxPi0UgGuIM6rPe7ktvZIireN2Meaya9CUlTgSXjk
MC/ndbTxFN07YqhnQrQlIozfjtsxTZkfxGxhOw+DkwCUNgEGFzw1aRhhRunWx50a
beH1jhFl8z4ZHCRtW3X3iZY9G7Ghrwna4iDJ4VWCt9fD3JVO5rAJnsB8Lh5iWbHV
wg3339djSC+l/KMRIZ0agbD4yqbmJiYlcoc2sgUrMnVd6oKt8KGPvQBLc3d3THMJ
T9mlCWUNTDomA+cpKluGFk1HVwNITqgbD5RoUkkDRoPyAZl4UQBSe5FamrahGccA
ZHGjms6hOzLs8+op88TFD+l0zt54oWFYRgcjwrpV7HUlmeg6hRT3XlabZS2Ob2rK
o/dTbun5LDLsvReaFiU2QDmPMlntDlyzRBSdnAnU5ZyV2LKuIAlkww1r1rUoeVbL
KCpASvCTuIOLx/AAyoT2JHPXX6F/h1ULccjZhyJlz4yKLYuMCqT0SErKjSTd1e89
Hq1ssQkV2wFZKwTuB0oH+8hdHzOeOczMio67GDijTscyrAB/yCo6YzBVLYEg0pxx
W8S+nyvnFs9zzeBjBBvE383b3hNUBS9mPfVy3+8ZgO9XLmtT/U6USk78Nf6k7Ikw
mFuNNn9h3uTteezvI8DgrLKCzQvjrHSFn+30TCVT1QNvzny6/rTkuwbnl/mY7fPt
r2731YQnZQAU3r2emp0HhQy3nPD5gmN4R0TZKhN4/Eta9rfNhCwam1oUaB1cboWL
p4i5Peuk5b2zAg333F0JuwEWKmMK+Zc5EVgoNBh27w+GD48Hx6AtTRI46oe5KCoT
S2JUU7Stg/yZqxCrhlHN2zagUb567CkvW7knCoI7GFV54Gl2T8FoJZkETRcWaeAS
X8RH83+qSMNaZqVOiUSrlJNRt7RSGTr3MYc3xsqmiSKIhOmOREsawcLOlefksqHq
j7u+YAFmczygG44kgPx0aA3cmZ2j3/J1SQEEkDsOOv7tzMxSc0pCfqENi4WGVz/+
XHM+au0RjaLCpTK/CeFw5XAAMFzaLLt8uxKQUzlxjLdViXAPAnn+uoPn3bFFwi4W
+yhimZFUlbVu3I1H1GnqCMrfx/8JxQ6JviyEDnjArw+m/VbU5UQjAUNZNWZX695g
2jQ+Xz38GW6J1S0IMchjgpEmSVt6Axn8qlP79CQB0XmOFP6J8VN58R/KRZGSuXKo
ZRVnko7BdLRLEpVylvnWKgYPG2rpvJzbf9iCy82DzKKTnRvYCR+qZfSa5vko0uj6
SeQTwZJKNQk2vzw2w+LMvY2zq8snq0wgPCShT+9CKOwgIapRkGkT0Sqx8oF0lqsF
4DBAR1L6/J57kbe9uQcm6/jFvl2Bpy5f6ayeiCULRPFJc/d+XTZCYU9xZeCeUs9s
6jQlbuYxbhD7i+LERivrO8+vvsSU6lgGltzRWXs4XnweDyzgiHGNxJUbKQkHGpoo
az0rGQFoCo1bT9GwGbzZOiQIBU7Dnb2hrCCNSmBHGoAEYTUnY5Z+4ksnd7frevWB
RXzUYn2GKIx0UWaHlPSCFAZe8I4Mu219sfpCKk1VdjOy3Rc5bcFDAgR5dEbTvt4T
28dU7eQ4ZQY+39e1zpS8sdcMP8I7YG6QD/0BvycaGCZkzwlTTM23YespXxwk6r9U
kNWVmKEHbjLYJyGrPP8j6smoAZJGd7l5vL/rjQq+bh0zAjfq/31ABwcq9HvoJgMo
HCuJa0JVHtHz2uQNdLffN3W+xKRNk0w26jhLYG3R2jHLYUrpmKpLAAzXEDCzM6yT
T5gVymj8szW/Uma1vIOmyRW1JjEdK6+vHYSI4azfC/Kq4gzkxdN5lOKQEuGCAXO9
/EF9Q5qFz3E4FNt6D7Z7fw6yLaWfeP7vR/efP17LoMsAQOOsw5ieyGAf7Tk2On4R
9UBrCCTb8opy3lPbDRrPJLWt3tt3cQ/xpyFqGd86Spit1G8op+AbDtJdev8L9StL
/nS1xfKlBVtNnDHml3FqJfGCoEVlYx3dSzXS4V9thH4VpiHkxNIgXbrKxH/+CeyG
deIj0XPXlLSGCT8JdsIq7qAjt3AhvS1EahXuGSA5GgHwoj4Kerb96i9rGwGUdg9n
4wYnrZOyfLMAvxKcevgWfpwgyMntWcKxl+qfIqxOAc33Fp97YURviyEoOQD0Q6GP
Mi+4uoT0Qp3XqVA0n9gG75Oxt960M7PbAiZjefllBWQQFElFrTzdMGxbQPTKK1hA
FDl5cRlx/XCMTUS6zIUiHQw0p8csfjuXTfmQJ/n6xgY8dNrl5X6qU1mDIQcZrzLq
0o+zdJhKftlcJs07PLcI+Tv5kvo5k5hnqK1bc8m7itav3DEgmltXhcHZJJm7QKBd
kETlt0vrDhO6XTRib25X3sjFumJePJxwcvFThN8/A7mF57Fv1xee8VDv3hXAy0Z0
iD57deOrjaAu00AYs74YuHUYiE+uqZ8uiPgdutuJ2Stzt/jkW+sUUYnJxparNnsF
HAiT4r/ltXpAb6GdLuGv7J4+ybgxjoP7ldNrjBW7t2/Nd8XXit68K7t4BRumebQU
Glu+vdZ/8UcMYAYUFBckD7ErYfq8Ad2gYm7IMQVJUvjZ98hQOwD3zGnMTrkYTlxD
okdS2BST+ArnfyjGK+loA70I/42PmX36/SF8RRjH2sI6irdEEYanqT8bcCy349k1
kXqsGaconiDYbblLZInKKwExVIs2toXuyZMi2efanH8hWaFKH7UGpMi2Uam8YWQ1
wUVaXCJ6CU5U3RJYdaWDab3V3t0ZouljpXXV5Y1IIkV1Io24gyPqXHGBhtfuMqyb
BOGakIoP+Mgol8XLoApDUODUAJfQ0GTr0GC/YgUz6AkTQ+o5A2SrJzA9iTHQtmvv
tJCHNeL82oEMMX1qtwL6Kc5c6x7qXkM3ALQFqXfteDHEfYik/Z+C9N7WU5BCwtj8
UeNeBn8xP0GQ/T4FWvvQTrLNGUQhblhO0UPvB5twfZQgKMHhupG1+vBuBjUsnDVl
tPSkBrckDhPBti5ZrxKOn+FpetVUuQmS/iRfIG+ojogfQd568353PvgdCHQNQQfR
sn8MeqYdqGctIDawIWkzxVSntAD60ksoMg+fV4Yib7syehzknYzAP7YloPjrfW/w
FQaYNnjT1mHrAiHVH/Gv625YLajyznWrAqtRZaAoBIppJtQJqyaljENFVP1X8BLH
FxyE0tzeRWtQPFoTjMqu5k/v9EmjWRjFu3V4pM4sgEBC8D+taIpwFfz+vLBXeMIH
srrH9dVjF4bgw32mjNWbBwRssNPhV7YohuG4MqdjFanP7JiiIBc7EUMljU8Pf1IE
jKpTUPv68G+ZBCzqAW5IwG520Pr3bBd+Vt48+ynmsTI9mVLMr7/ZMr3pMPkyYD6G
SUM2FPmh/d9y6jvM9rZEUHWqDK/NaBuLGcLC9opSYgkCTp2EjJ24HB/V6H5GowyK
UwECTHCgA+FB+u6g0NANg/45N2G47o4PlnO+uJofgEBLEtRsjQ8O4OmAxQ67GoL3
+mx4Ed/3zYIGH4cen11sVyFXYXW9bsPDwpZuaZKXBXJL774TdzB34Oz7eM2xuDjA
Z8hs6AYTZB+TTJwMgAZc0l+CinG6/V4l2/mGCNe8vNvSxfJ/RNRN2l9Um/DfAwmB
FGdfuw2iIlVErz3Hqhf5nNhiHkFPQKRMH5aw3VTXihBVV5c4ExlfrAJ1IheGH4jl
gvw9ngcNms3j3F9XtJZP6kFlPBIAX2XgVFPTrRsCOsFLWaRuwcFpzz8lhZ8DGG5l
D3MBx9ji+nEkgQOnrnkyW6JZqU4fjgJxSYAjGlMRkx5Ln/LnS/ldAOfPxyluUaNM
Mw6WkasOaBKgwuh0DRpTix9I4hdcuF1F8+w2uH82gL62/4Hq61+laB7b7CXmq7TA
Xeddhu3ZybUrH56JpCvBaM8kHy30RX/zImkKIeg21VmszoAgm4dOaY4TEZGb0lgO
c/zMUhoBdY4Z9B7tyZzZzSGMa517GgEn2IXwvg4ACWZlGMSK+VbFmU2hSOiKv5Qj
pToETBs84XdLIjLoD3RHPIXMqdixP70A0DtB1I1+mqVw4qso1Bp4tH8th+LJGo8v
0y9uY9d/UrrCpYWvYUrGdb16Ft0aE+pRs292GfdEDZvf5IQjveTvGBoFaWaacSlf
8BemyART5ABcjyW2sYYhnHg/InQGzfTZ07O5VdWBqzVkw7h1x/V+VqJOF47tR75x
w9wUN/2kMe62T7UfmBW37T5sdiDpT8FN53AzPMd133TDKfU5If0uiDsQWxrNIu1o
1CMZbHicpDh7CivGE/jzfmdSEYZUO16DP4HOnuj5OlwXUOR4rLOacktPCnQR0ngp
AJwHmA11JNi/8vF16p3lD4wPKthVb7sYJjP1lTndmQoQGzBJHhJwvZKo1yd2uV6v
QC9LCr7yvQlPeHtk/6CkR7cYoV/GNhEw3l9NipdXcxQ74hfyqAquUl4ssL1HH0d+
lWA36po2EQOi2ubj2SG4cNjFcuPLcjLfObXf57EyLycLAtZHeYwmdLw88aOXPXTj
eDkyB8KoOvcpzAFU6ZyrMFOihfjd9yg1qPFDKJQ6zZA/smESBrHWta5o5eIAvSpD
qMRP2C5QKvU7Eg7yDBgu/zhXjz+WxcTWHIcppJ1Rm3Mhp8eL+vkKbXDUt/ptL97s
3wZ0abHwrrvttkQRGjWmH7VgmodOCegXPDwuTFcMUpLmLlFyiILzpm0bV7QcL8XS
CyrQr6uQoKHo+qevq3sg27sYYEzhq7akQv6mN1XV/0lyoVGsmo01qm5VU7kFGiqT
RlMt5Yx94k2jiRbfWlIK07RQFj0d7rDhP+OVr1sNVczXBvxWXs0CGkbcWlACsAtG
Q6Jg3Hp5vtx1l0LKDGd3Ttpc2nVs4A6rJIK5slqGWfbOMLKcdS02X6h6KaSV2ntN
8TFhPqT8laVkHsdF4BWi/FAvamwu98qoCaWWxfov89lKkv/7oBcgHX0KtkJq7Y/L
xA0+yzsrgSlzcRywzZQarOox0J1CgZHxBCZKt9nKMgPQRNHmyy1k1if7NvJJIaVY
NysWf+nZCEqCQa/9OOwZEkrSk6+zIqNPloP0i6zFwy7MGxZB4Mrk9G+PRYiy4T2q
sBPviExx6580hxR7BFuPIb4ccoI767z/8e6MkYpvAqUmorPmZQxMfPam1+Xfp+Gt
KFSpnRKTY7mr2tL31+a2shz/8gJpUyP2Ax5k3V+YDhu/ngmgjYV7c4jWYfB6xlQK
/ugpj3D8tz4FJOQJjB/z7oOb9IKBtt/9Cj5Hr9Een+wgn2w1MZeXDAuqpW5S2ibh
0GBOcIHw7RGOL3gxCa3zYY0yXtIXhkehtkXZk3CHnRMsSkNph1HrlNvdfsoUn5NI
oZspXWKsNtqagrNs1fwNwD0XarqU9Au3gtTNuGKDcgIvcWdJOFkiEKHB+m6qXtyV
1HT7+7UkTBdcR9u4hZukFjnIB4Cvdjq4vJxCiKEOgQjYSObWBy5MQxktFIqVQEC7
EY9o79ON0HpZmbxw58EbfPGcGURc3hCIz4KToGdqMM1gE/MEn+1PPi0vi12XzuWk
e63d/o/afIGdwbc2ECJOozFVAcepUmAnpopELwmOeBS7907rWjUQjase3ASc59jE
DK/n++2qnL5UTRiOjbpZsZSEx619axN5kxk/XoUMHtSNW+2vo6+ll7aQd8zWPYWB
lt9sat8UhfWGH4OlXTsAFqRqG2xf4LhPh5OO6pWZH+d/M+lzZaoeeZHZDQ4w+be4
zyA9Q5SnGDvOlAvOcY6J29lyMeQ0ENiytjDZ9JQEHbCeCtsGbyGs/LpdIy+qXDV0
6rGYUHumd8WApdutoT+2vxMGcLN2jmxVYnnK0fqpRjzPJKB5IU16QAwelZf+jNE5
Iw/IXVCh6pYqeqGpg9h13RPaOMErZWmWeh86JglgXCr+AGmZ90dNDW1VsOcauDaW
R/pItcuK7G5UZE6JTELYGbdPRpm25Lg7TrnpYj9uhjKABVq1lh4hf5+AcLbcHlM/
oU7D2qteTgR6CgIMQ5qiJ7TgnKGhIjyDfhu1UR6R9qEWXVL6frtGaw3X8hDwZJlh
gpiiw+BYfiqfPSfloASwdCEWXhn9ARx/L/HJ0e5FGfMuKz3kHUNjFuq2T5t8MR8y
WLxTZ8eEtdXjBbmsTU/R1jaicuNSfsa8w2+PsnNSlzp8w8/vYScmRCZ+yAlo4EfY
+siyEvpMAj0c58F0J59UGIq2T1503/A9aO1dki1A9KlqirzvbSTCkPbmgn88V9ox
vu7sUt8ZaWC7XfnH0N8XzGhvUuKaoGlhyXXR3x+8zCiVVYJyWVfRkUpMEUJkhvwc
R0leRXBa/MwGZmWag9YHKo8QL8+wCcV3jdsHGSG1z5WsGI1t1l8mHZDWPyuMfQCx
Iy5lxcOAUYXfrWqSMh3BD8VNBtTQlUMZymYGLdGPS7RGdOq/ygdjevyvaiFEXXH/
N/AaI96s0I69Ek3qL9MlqSyBEAn2B/RRu0HZVRHKQXEjGid8wwPOs7DlLM86n8Cp
+Q0ES8soupCRgE7OoaQM1DEZcWhdbRDnjiHT8DuE8JeMGalp6BN1DxuXqlTee/dd
Ec1xbjWMpvG9n6ItQ2/4UsJhwlpVpi3H36Mmb41j73SeqIGb/QQ1LkhS0el9QXyF
X6yjxghCO9SRYoy6SFpFA2Bo6IianOpGSzVLRIiQS2GIXv4842xaXlsXGkTQ/dFF
zd2lLanK3ORh5Kj5KpKaSQ8YEcl8wElvGN7NQi6cBcZZwg/zg+dfUJyleSiL/rHL
5cbCa1F3MtA+MbSArtbJBo6v7rbpkW/Uxqlf4XVDw0geZw/i4A/VCPjrXX/Gyhx2
jwW8zALcTtDOOn4xFK1eGXoqiccqeHe6dUK0hIzneUZ6gru/WU7eCSQRhr9oPxtg
bb87Pyts1Zzy6ED1iAZxokcGH4kdDZHQJgKJi9YmBCyb1tJBRtZYS2DL2GECMx8a
+d9ZX4uqyaW/XD4Qx5HB5RNuu3cB5B7JgzFQzvFQogAA2XqfChSAkdDGjAZvWfK5
1reeOnYvvu9adHaIxn2EV8lX35V/FwqJKXHX7fSajo4O+2ExUFo08YlfnOsaz/CY
CM6k5olIvibTR83M1mZ14ivYT+sIIqBHqe1EZ0hGVdxRqzj/3F3q2j38DBrM2aVs
pHKKS/v+qoBdfXXTx4fFqAvAUGJ5d6pyRY9c4KA/LoA5bt7cCfHX3sOYH39qGMWu
yKo9b0nXmterJ/1gtCVOS61QLUZ6hpVnG8cJPKOZSYd4U9qPYWafF8nQiMdhDHPq
Ai5L8NEjyPGB6r7gwhuBUNJoItLZ0D0oYA9U9lMMv3hZdSy2TPFNf6eoG4c2Srd4
7cqKWVXgvSOr15TOYi9bgrURr8PW6Bba6ZNH9L+9mQtS1riV1t/t5fYuLMQGXbuU
d5l6F5Me4W4oS+lTk0yl1WeEhFziiQudWVsCEDHM98CuO+rnM3BChQKwK+Nispa5
V7sRejcu+Ky2TvaFfT95iw+VRh6duWfzsY63FaXa4V8BzGtF0efEEbsQcnsRk5+k
FDH4XL+qF/K8Ps92sTJ/TWz33lLIL/v4vo5CxJRUnlb7wGfsZLri+8w5GN6Z9p7/
LBSa05ykwDlTpO+vFgHirt/6zYFHArGkRwLuf2MlI7IauqoplDnxHyeTECM8BS/p
fjtlVCTLtw6774MXQxKXVCNDEQUucH/3e5O8BkDVRnvVg6LieaXIdIbsZcYXyRun
uneHJifXwgx4Z2QXqrwaLV6JLrxVBC2GKU0QTrhkX7TQgRt9z/aNMWy6+qnpoyTD
y9u0ihY+gWMJMUZqu2x7ovazvXC2FCEAHG3HJI7PKK4famOFk+EwagNu7Ti0/YWH
9c7Soac/I34Ozj3rz6fCANsHC1MVaeUZQcbG0SgSNKURjXSmuFonwNB7dFRwudPV
LTVSkcimfUj7bLLVe/Cdgjang43H9IoOTnX76irqqwBZ/Lo3mZkYypYNtQwJiqtv
yBVHE0rjA93y+R8vYV13CwFbT9HnIQ9pu6y1uvsxoy2u+iRKt/fdfgZzOEAxeTtp
YU0EucsToCp+fuN1C+JXk/wzfIY6EkFCj8+TYy5l6bPnOtYK8XXJXi4w7MwnjGKv
sqaUFl61wdVqurYWOsegcOKA2VW47CvcaE9Y3hKuw2t8ZrqHeJ+LWsYrD/4lwQBv
Vu2WYUYvaRxIq3d9H5t/s4Ud43WQuzZ4ZcZdcEXw6SxOUyw2Pc2L0ZHdQ/cO3p66
JPSlguxEqJ3ISEn0NrCSocBKYWYVRXv1VRl+5E9BcPeS2ufT+rpVcNwEU/mNPAhq
foryoKwcT5EkSDFhomALRSaa/gV0kE6LDRqlzgubugYT0rJgdsFkjolyVfUR21if
FU6K6EIN7gHn/Nh6IT3YCgo9Me7qcphL+hrYh9mMjcXhg+oAn9o1nmbUfRi4BxAE
yoAtGTmSg9HzSl1kgI5luG49oz7+nzMcMNOJbn8hN1/7jpc5LgsA87FpcQc5zHL2
xgpnJfCkiW67iOBY/LVe2tiVHiMyRACu6Q5R8GInA9O+8abFRUmkNWKCbbUnBMLF
sMxkq7sFYPMpcGT2jOgklOuqBPzPTpj4Z1AlMtK0nXAUc5rmkmMlSnOowD+Bqxdi
opDBhL5+PBqShcAwNTerXa3/1IE7FPjUTxjkUgvuyfrI1anyy/e7AbPbHUoZZc9y
KHM+OObcLdOueaPx4kZwKTQegNU4f7CliMjDRvt7lnJk2FGWofjbQS43Q+w5GSKk
dIMO54WcHZuvgposWFXsswk+0q/RIrxfE0OvpGSwYKvyJdVLchVv+zx3/YBh1fmV
SRFm/3Ib5ntT8W9GEyu0PrpMAUN5/ZCvuzVF82PYY37zfSq3lrrGDA/i0mJuERrn
HTRaHwwphouV1RnSzYP+b5C0D8QeDNnxNu8NZaNIDMznP3ThXGu9iG2hfWFSL/SP
Fc9zbTm6nkERjOY+vZUUBZC3WjrauDMb+GeOuASp/2uPqYlgVrA6bPsHf7otn2as
keI4NdpGB3pqVF70Xo72F/D/e1i3dBjnNQq3hSnIpcM7O2LznZLp9U+Pp/3cb5kf
wvfHFPiqi14BeDdupYkIvJlDAAGvlN9DJotGZqqyv9fpBY6FkDuNi4oIFZQ62mL3
NmQmHT2Fki/e+RHcfBwtW6ep8VARwOQfEmmjmIdlT+N5Xsc9YK+EpgtQge/7UAgS
VvnQ29FgCy82kHE6gXKWNx9QkjO/hsdOzNK/pAQhCwnKAasq3q2wWZt0aAffJ10l
M4UR5DO3bIhi1qRZBMwusP8FZ2AH9hvMEi0JIqGv8TjUP5F1fJP+ME2AWMKUdMP5
dSYGos1LQpxge9qd4F1ZvqpSbxudxJR8Kc8sDmMHl4OSO8ohhF+guemmqjQTYmr9
zDT5vVDI1VNFdq2ugUQNqjOJvhWd+IAJvrj6ycC1sIsRQl+hU/fGOJPCJL7388vS
/PchzVUZeV7YpDNa36GIGMPQ1sM8Wz5ns0fSc2mSHcYV8TcaqkcnSsVJCxJz+29f
UI+TJv1dcssdil1k3p7tHFYmxmrDlTtIrCbPc1D41K/omBcYOBoG9UJKpeUsK3/r
GniUCj5XiJs//iUNZKs8jSRyi95yVHp4GUDpXiLoilELMV5P3ujy9FjTfhOjlCky
k0HEJT62cRGrNum9GJSIOFIefcTa1/FwWgYvri4D2ZATtD8MOmjVDAJRbunpt6st
aN7CKAp85JtXaC6nFIVm6mToPL0pOs/fU63COrJEb4Ew2aFuay9kFJz7Z3N1+p49
E3DtswSgHiJpj1+KHWjoDRAtO9I5QqdqlWVPhbumrp9kRua6KsucYqIj/XKLyqgs
+WOCTIF/rHyqXYtyCzV5CgVsBxDODZTuSMk75IL5z9WYHGJFt3db+m7jVb+ECTy+
eCMYB/CDfkOFdYzQ4JLCWLQfJi+Lb9eAACco8DEOfrAW/F5kDzEAd4vXWfwuzXGU
Y2hp558PH0E8/vfG8UETQ8e8wdScp2tdhrBmZAZnuYCMwp2coZAXxGzblVh9Ws+2
X5EyYiOAMqg+AhQoUrc7g97/G93nhGFGwPkr+uXD31GyyCVFKwjkP6qqPFQrgtmr
VNgHh9UDgtl/FzW1SFoyF20jcsIXu7u/BqMvBGlQkwcGz3zN69MyGf20pMVVqZC7
+eZc2m4XmQ5byqmF9KI4m+zUYPM2sZ0y6u3mTF69N7MBioi1JkoT+QpRYBvi8gcx
o7I2SxN+769AyftCgRLdPDfVnWmpok8RFgeCPXynAHRUveqoGGlwcc9z6BNHQ8Yx
WAW/iRpnc4YQr+63Z8qBGub/jensi82/cWEBGZZNDNE1a+aMWMepjranGahTDg4/
2UYZYUeJrKreyhSbeRfe9cFCrhZPnZD9BiEi09uOOoW0qL1A1Ed4FYRTEdM7XVEU
U5MSHesk/SMw/TcjeoEq7hBwqKx+Bi4vjjE4WiHc+uJEttBXTs+t+3po0F68vnnR
+20YOamEmTX2fR4MRbSbMZoVQtlOLAeL6bVIoQ+/5bvbLIxFTVrlNSVn+6mbezK6
poP/Oen4emJQlQ+zgh5pmqY+dXh0FLOOuPyV1uXJs4bWD3I4X0sthzqjQng7UR0G
A84Gx5rvtb0vEc9etJ4pT2d/E0dlIxYZdsvO/8+pYQjOa+V9iY4X2dUqPSqc52D0
clsAww0DOSH8OSw5kqJ0a7nnFdKx4j4hRpwzS5RMVCXkGJ3VtQ5aHnF3eM1WVDDT
h/9iyCBSvUiC09liDIHOFSPk0BnLK11gxPVgAzJfhT+CeiO6MsNPMxPUIQdAfZku
AeiwCRGP+c1xPdxZ7IUQ6niSjj70mRnJBKCWZ/o9ZFYl+kpwv4W7rfixy/kRxc2o
fTQ/6Fxv5mgwgiC7pMhAV0kWsKevGzFON7FRFHfvhPFE3dB6ojB7+rYkCIi/mKnF
+fIVJg9LOEy1IlVwMnrzNiChrxRViwSxEq3Sr1E31Q8yveVULhPsm4XNb7S8xf6f
ZGyPlmdvCubcf8JXMk1911r06zVKE4/JxWkFAcDTo6y+jI5NKwtw9MWK39L84xXK
Xa9Wq1ocW2Oo9jVT5YXDd8Q2VUN9nNY6pboeRw+vlHkme0z369kAYftf0ZFoWRhW
ixKwACn4KJ/Q7vKjXIY808sGsL6gVZIjO4qZdK2fOdJ3C+zZ3K/EJ+pccF2wrjE+
aq9QDwaGt+EdtLheR4TzE/CW2IIjIrqpXodysnYOxQTZUejv5f/6MlDrP5KuZi5D
iDYxrKloqjt9ZS5Z/Sh3+woqJ+ZXev9Vlslp5aBPJBFZONkWR8Z/+J1K/2m4mv1/
auFQ7HxBnWuOL40u29EExKyZ5Ejv/Vj1hnzcYC/Lcu9XJ0DTwAr+emDprbuGWKgP
iIgmO/l7i8QqBVPxr1+JQNTKQd9WwUU6ixq1y9V8el3tLKo/DyU/f+hxSpBIHymJ
vflZACdqsc1mEFpqCn39+8OE+5UlDGX3OPAHg+KXMkhyP2j6IUDeX4hT6KwuNg7P
T8q402tBoYLqVnAboFbjs2SL7cBma7sC579P3lax5XuTc4Cuo+8lvPwLTH8R1+ON
GtlSNFKhFzb6M58uSMKAt+lhFTerT2z+af6AFdJmE+46Td4j/Q3hWG3fo8E+kjYY
78CIApovTzroLykIjfMPsoWXd5SP0VZbly+SAR0OrHtGZnPTKmVUB8Ab6JdLeM2y
dUWvSZr1m5cu9l3mVDV8w+jojrq5wG0IlNezjvVszl9qR9xMNNxURTZGQ2tcBYXF
+/Q4Wv7nezqjykDbMzScL+ICIkztup6nbYfp5/dURVhIKnY2OBprMHswfLLgLvDR
4pGdd2kCqG47unWgLk/XAznTSXKcBazII4unrk4GnK1eg7oKoD4ekSdML4+0w+xG
39aFSyAlD2/5UhGjtbvHhR2Uumyq9kIbIABnW2FZgYBzy7K52bY1r8EH/RO/Jqx6
n0R1NeGYbP3BcTEU13oAdVc88KyD7dZbTgiAUKoI79PjgeeO73HUVqZRRXLD1/03
71qsDYUuybaPuj/joGonxt3eDyyLXoFYZ4Uj9GxfDpz0ANMmujEa1EpyAI5IkkL8
DfhuCw299WEFYUBjgdFnlyCQwF0KD3glTMIk1pIGJM5dAUrZZW5g9+9+PFbgXcNH
YHR8ogKvCC27AJtGMa7nIsFIwqwSGvjb7uC+Z2THPmhru5+PX1Y9Vt4pMzW7d8lF
G1kk+uQVtnDMJR5lfRGUHEEz51GnIi+QXoA2jKFIHR+xyp73IYxJ2D+ALhpOFc9O
U4fDNJHXmEzRSrIBRX0TjvtAe0myApXm7cBgBSNWDwhiTXkarv0rTfso9SNnR4fv
XuRtmRXmN1zxElkIYpimwVPSEVsugwZjrCCiaZX0b6JP0R7QiBCbn8sz9u4BVJZy
qocJvoJj8TMgwWA0/GNjQNLN8Agv1DgcPGoNlTJrt99eANDroyhM2m+cZJwvaJhf
pbhiO7px92KAHuODJoLuvdBc7NQmhWFmY67x3MnldAvzD/6IH1z2A7pcl+S1UpMl
v4/P0KwFr/sDNqausj0A7ae3PKpRxfBxhwdrbba0jXaao/l6n+XrsYSEaNv94i91
Qs4VrucbE0tQHQZ036YZZV7fzc//ETaj0phOtcgGEoIjEWMxBnISEQbu5y3SWG0F
e+rkfmaoMYGtmjdMKi6Cn1MHzd/vvdsIelZnIOKDCS548TG1QMEOtZFDTodrWMJk
wsEU+r/qcsHjDfA5f5uUkbrz5iynjB1txxDWdlr9U4x2EbMfuHBKgcYpcmbIHzD6
C0uZXxrXQH5aT7vN4Oe0272CAqNXPzFQfte5kYHGW4kbVPxkhzkBn6tuc2guKEHu
aKu4OLguoSPQJQasJnivwvdqpGIQsuG0A3yXNybL6C4kBYeMVOwCHzVyrKWYuNz7
/L7ataDEW/R4CqS/e3nCcz4ds3AZaeODJDaKtASvWr8vaXB1v+B6erDX62RgwEUS
/h1Nu5jLP8FLwEQ1WZYfWITAvmuGHcnmoRaWYV+cNH5NkckIUgIRSg52J4mOMyDQ
q/F1Qn3eATgriQYsqoaVUoOPVWCX1DvMjLqOrpadGw7Wy5uZcYC8ZSNPKnMRsEDd
xcA7gHfIIQBhqLpZDjqkHb86rs8R4Q/dMQ1C+GY6QJL2AwDQ+5kPfj0rvg3xgFKq
RHjaTwgm43LAKjnC8okr7K+dJghb8hh5WyJt01s8IgwKAAAc+wCVMsvn6GHot/SJ
89vN1aFp+6KFG4G128e24MTHoYd5TTLUzddpBisdmuFkqZYRBCq2pkDo+icF3O3d
GVa24bpaf0UxbWTmKJDpanhm9eR+6rfVFzQ7tW4X/uwvQc/qclEG+WyDB2OBHpH2
ml1ZvVxEphOpkmCpzl6w4ZxC1IXXFBXWOK2ddo1zHkirbsaBW/b4pn5F7KQL/f6r
AHNEbgBjvQdk9sA640RjCvagcmhz1uZHBruJ5S5y6MP+4glSZIXl2ooFIXR1VLfN
nv3ajJVhqtXjbTSC49mOtbuuzwuRVyWfqrtDC9cgrNdtBev359ZhrzBu31Skzzk7
+0w9W3qwexUN3303ZwjGgwKb4hwA3bx6DBceIUb7Eaek7LIoHwoOF9IdgdETLXaY
ZZw9P5mdVAIs9ZehYk5xNluBochN39bNcCfkp7+6nTNoRX+OPaA+ML4mZTbsZ+ZJ
EJb21DNrpMosEvBzszSQuU+y7BceZSqng3bUgit9mpsCBO0no5asOhOqsxnMp+bR
vPGCO4wFffjnP1B43b1g/OnqzNV+U0Y+oVOu7gDFmnXdYv4Qmz9MI8hOeUN/8du8
zeOdgfA5uh9eH23gL+zxYU+/zlPsNEbdyFFlq/ozGJd3BUw1PhTktKG93gFEt/4C
tQP2jFQY/hkmd4x0k6J8C6yWz9/n6JpQxmtqWHdxpj6KiLeiroz/92nZDmBOZC1X
AQ2bHiiQbpyItS3i/CK2/7w12DmgIdx1ew66PfJhOvyVGKJhrYUvKH8zja8uvpV0
Qe1dmyt2PNPNwIyA5LF7C05l1NRZBMYj7uwG5HA1dX2fPvG4ZhNNdfKZK5ac9rbC
lCvfd8rRDZ1BnSU29/Ne8ESSwNZeO8jn0sbLytOiIwkl8FViaiONcbX0vmcZqOCI
eX8tHNiQVCiPHw2PjrIeaa7Y6DxGJnJP+YgCG8G7VokSyIuc476KOsHv3CG1UGLa
MI+/VQ9ZA7EPSTW+atpczEQQlvrq443ATF+v2OsBks2K8FZrcXu4KrARkqtlC+VV
yz3UUgjgEnz+zJ3+4wmWnexFv5upkGN5yjU9Wc1tZSDudsd7PDMM0+VSVGem70fG
iTwlwYqtHFz9+ALGXb1sEGcbqy4YaAzgwTUJ/RIUjeWyDwcQNoeyeYxYnwSbhEGY
TDyA3iNkScvHMWXR2rZw62SvM/vkK/IvDHKgQk6GECcJ/oqlXnZyqFAq8fM+Ycl7
vUdaozd5LMQMlQQ5q4NkifIqE7NL4tg4UqpxDwkeMcPHlwyDppK5LjfQdVTVNLMj
RYDifLqT/kfcj1dXM1JbNmXwwEZlJxesOdxa3mjmO/HZzVrZYsvDHSOCatqFC2Ys
/3djgiVxdhMNjt75dH5T5VVqsEBhZgUt5A/kaXp/38273+3KjdzpbkWra3sKf22M
UeSqfdaL22wlxczT/BeorMRqCoVDLRMM2MlxrQjfMCzhitLH0ukyoisU5aeop/KF
pAYzGIXaUs/WwfX/ozm/oTbc3ASELLjqLYj5n7gs0bOBewHhfYThDsIa8ZM4UfL5
R6XJjmKo6ee5vaLUNgxC8PiEWvpnRYoHulM+SGOItEicVR6dyYg3ac6mrFeY55v+
v2TwtF05jTG1Yan5cftSjGPztgawUaeSAXAswwrzNzizUv7b3sLWXKMbTLzRD8R9
cnZ7zvFuguKrf16a5jjk3BWMLN2nshNjOdv0MOcnEVd7qk9kAaYY02lc1TvW0VEk
/4zngEWCxZp5S47TFPDISKby19Zoeyn8RrrriK/f3lAsZGBczU/OymWyC3K+SMM+
QS2ZiFm/GeXSdzl3/wIZJn46AgVCJUkXMku5jDnHsjh5QlYnUByk4ttANmIheu0L
YmMQhTulAVQnNZ8OtmSceeOOubpBchDsETGhILhLumPPt7MKZOppkoVMQXnxwN0u
9oIMt5pXncWuJjxggPlwOobdRxdw37M5cCvhtkrbAplxGbmfYyAlRrofRl2We4Hg
OiADGuhJsy2D/uJZlEQmN1ZKDM74ILY3+u6Il79ytMNi+HYJlG+mVlB2v1M9BrHA
nee4tVrFOoZpRFzWN7Q+KOQgehvdVzf/C++lrPBqajDdBGcWlpt72l7obCoEjM0g
RdEDzrEF0xl82vHWsoyDYmMS0f1z/lTTwj2GsScwj3t2uV99guTyTer1aJW1gjRx
Qz2F5i4Bgbz+1wshwlsF+XEpCy3AzYfTXHqRo6TG06SqfpxSrI19mZbcHdjClgGN
BuGDAFQrVy8hLVoUI/pIOO+M8YQNAEjrMduF6s1N6+jQHc2MNIoshl8X1x4QCqdR
VjVUKEVLD3uzcLS/Z6+td9kiPmdjlPI+RwCKEL1+ePZybUf5ZpAOVERznUDxe22D
wEae4fWhW+B8Va9D+dWuhxqg5CefgELHLRrEpP3/QKQcZKn9tOMJX9SXpFdRvr/6
5VWHhXCSKF2dkovTUch6Ejf7Seg+JCJ3Vaxct2hLGDn8xLdmReyuQLhjdlo2xs9Q
JQ2pbIv9gHxfY2cVK+MMn3AVSoY8PCaFPb0IdzLyp8s7m27MAoo0rNUa0XOE7MWd
aOZvwSrISl5XFPBf6rcUcsEysPYcz5aAmOEk7BBMrjZgyHCSzCq61zgqBwmjfc0K
SkTpMTgfss19ObZ7rvykpHXvwiW0cpRcjwxaNrxJJ/a5TJ+sg0dR5fiEMRX+HjGb
KJBlSubYClDMN4gWOFxKkmofwng5HgRFTDDv3CRAU8fjpJxBToVJqTVAUxGsGxr5
wXgK819atibmnuFVw4VJyuzZF9FWPZMAixwA4/wP73xQcFCJGcPrVPk+4/9osCzd
jlbd2coRp8SZLmPqoWNe8AK2wVM+pxU0uqLa2UdlO+C/lenX/JqgtceblNdtOtzU
8olT6IMJR7DLaeekBReodNqia/pcoWwjJZYzUg7R0I/3SBxs4+xEVtrW95POZJ1X
wNt/DrmtXZEzO71y82Mx88LAPid5fkmywNqfVjv9LcpdS3xk3albLy2NIusDdAH3
s1zIZrGzuqrEQRoVgzhXbHwp0mHeqb4ME5isMvQr7LnnX+dMr0T27EkJpWX1ItAf
ltfJoWBd6EqwcjcSjUZ9OWzdOgFVLMElhEkyygUXrTTIBakoXMd5pLGoluQs3IUd
GY2TG1KxKK3wzQJkqkvq54Gla/23JRlIiuyvHzIn9geT+2rJ/ChvlaYKKEhxZWLX
Z+88cHPYHJvis7Je094P5bpxsinF1FO5gpG4CIgtNjhivWEkqo9M89PX9E9+C166
FgCRLhHfRRTaQohgVHTwQNu0JlpH2VSbPedrX8quSnoA3kuoYCDxJGSKHtVCWHFc
9SO1MItgsfQ+0PeB9ftfzemXROjrRoouQxU/a6WrRYvylzK8jthWI+PlERD7mo4K
/Fn9lWbGlrSJTH3Pu120XLS6paddxTUIKzpbg9T/+8JWDdC20nBNsiUOezIsUt7m
swyXFkWtei1Y79TuNTo5JpXmhcfwkXxl+I5Ek2srPBPmLo830vcywv9O7BorKpdv
V9x3pYh/sWvBX3amqnQxTQ1orfzD1mxafjv/dHZ3wK6Jdk3T31PlI97EyXhVpV9X
CrH9+E6Ia7PPuRl0QpJMMzkeOwdaDUepB0LTQHIgKr715kof9UqiwSztY0vIbhbO
1pcuhhAvrwYUroFvp6Lowfeugx6sO2LZ/mFKv49ZcqFfjNjxaTzd9ofGGD0Vxagb
/TbTHXdxWCM9iV+vQP9PAM6s3xG+TDh+/vjEW1hLEBwHFIwWQHqsMz7EWp/V3wqu
ZGM+RSfwv50rUuAtT/mE2cYSrcynW8A0oGG2bL5jGLtJl1hTs+6jyEV0XI9Ad9Mu
UFp8KCkOB7iWg9CFOlFUM63yI8T2o4VmsDP83DT3AqgAQ6TC3kNwrc6wsTh76M9d
wjBX+cLawyyXbZ6phRKBagv5qN2BJX5MhRj+V+YJKlQS6l8ZN3zKzaSeg36bHhmL
00RjzM8VSx6q7Glir9z4hfzhoaoStIl5rFiG2tMFQLn1vD/tKzovMQrS7MDEOmd3
o46SCnns5u6TtjhRysQz+V4v9cQFo8p3MPh+qA2oyjz5SjokpunA5TGYgCi7R18o
y9pES+6FzhREewhRBdn90WixtpAq+ynrXQbykE7AQa9xlheoDgrMR9F7HPNQsX7q
T2zsMsn2mUQs2CngQ1azY59joztPQnizz/bqtZNoJYZF4tNxJGriks86LgH7T9Hj
ZKeMW1Cbd4xNYuTvv2ko9x5a82n/yfBpzQeAl798A8QwTj/INQW/Yi/NHRKvkdLK
RXm9/6bnIrNw5ZriuXpg0pnT30bsPzuBltGqGe2mQ4MCwT1AqrKjw8wJUXOVLfTR
DHFx8nWe5efcAYJ6r2Ey8wLWI1170ST1aWh0HDyJBMbkTt1GrpPXTLI5nzoLrlOM
2R+04qNY6E4rb8SGgeJCksdzTn3zVcbQ1V3Q7mBQaKLvtCB/QtqwrxJqKUApUeKI
Ak659s91MBx3M8MaF8qKGWPNSDsD4Eo1F2n+BqWhOQzRmo9LyJ75yeHrARzEC2Oe
ZHhX1F89Q7hMkMvq9CoDuMkBd7KHiR43zIO+IrOmaWEPp11I7TH6jbBgQSyTc/UO
AkGT0GowYeiuupE0jWlg2AxAlLOTCXWnU2H7QrN7j+UUJopTS6vnY79KvdTiGjCa
fe5SokkIUq4/RtRSAQnZcYnxoYInZp5uF4QnXoRIHP1XkM+DCCimURzxeuXdC4ZD
m+cwO+c7jrEhXw1Xt3bRJ8flpVexgzt4CDwYiEgKV56jVTWHocD00T9gvbMzCKMv
g/8ii+N/DiNX3DVgwnWERfGiuFalD83ldA3XvAxK5AlF/LKU46pGz4ERuQF6cjqD
bcu7Jx592zo/aSlBrEH8h53OE8H9UTG39vnrzm18iU1ECfO1H7ooS0LIbjyRpBCW
gru0D73FJD1HgN+DOBoYsO36NpfnKADd6I1s5J2aJ7gg/m+z0PtXaUtZwztgFGQ8
xmwfkeH1oUx+IKyy7Q9S6jTEKzCYLExBUu/UP8KUWNCu8J+W1QIq5WqGqiN+VfsM
EjLER8/L8SsVf9O+Ty9xT0MiF0ro//YKSxaKeXGhCcCTXL5N/5D4G98C0AW+ldsO
jIdB1YnKNCP23o4VUZw38x9/ImjO8/6GQLU8v5lP2nUqRBLVwQWhDvaLntifsAdN
WWfmYZt3A+dbIoFPnpKu3yV7kuaVqsmgy054RSGtBfvAvWHyjlZzi9q/Vqh1sE4Z
zmWlPu99llhkUu7I+sVBI/9zhoFPL9CXDdePSm3nKTlztNohJ0CDjaE38Q3umPIJ
bheP89JxpplvPCR0ECYjiBOrzqyeGF7ZQLJR75HCtKYcufW96YhFL0T2fM4/pYQx
vvoPM9o3Xl/mX++Z0wEXWZsfqVvvVMr8lpeTTAq8R7TyULF90XC1NyV0fqrDoPuA
xNdgPqlq2dXJslKaxQq7MNc7dTZuCjU/IjF6J9UhzwqkaCZFCFJnvshkwIuacp25
CHSHRBWCiFxSeIsAcOeJenX/Xj6aVb4jSVuIJamac0DThE3Hs2SaWjGpXNZaXLy2
J5koJnV8GZ8p/IyyrZOx236pQQFMyTqAbTqznUTfyLYY7W8cUWtLSQkOqYxlhFWk
YkCxQQBgsJXotmoOh/zLfU/BEcZEtvZBfnJ459MVM7phV48MHrxTJ3aUx27XYqSb
KQLckOoAclFw8M/3EDHc3w0tgbUa8j7pMmsCDbpYv2jtN4EDtAAnhpgzgfUC+6s4
J76+1BJCyGaygw4q0j+rlJy5BS0OPj62Jo8MlOKUBp0wYP4Afms8JIi8V6/b1W3Z
PApORIiBTnK2SgIT5Cekwacr/pSEZY7ygsT4omHgA8nZYDva6lyl+LJNEwSYw2Sz
9VbTJ9T853jZVJbvX+PkQ66E8+POYehQv3BXyJqBLtEQh9W6HFuwY2C9usxqH7Cv
FzuEGjHfBbV5Zwnl/eX53zuQe20A1gjeSqvLpCMKEUtshk5HDMETD82E5GDm2e//
YRU5/nXmgusCXJswO976Ik4YR0+Z6Z1twjBQBCR5kfrOaeuAPoQiulc1MsWBq9Vi
rGJ1CVDq3oK+DolSm1RcGt9hwVqUJHwuS/gIgWNyXIDNHgIOl1dP2LzdNSldPC5B
664EuCEiwROnEHgfpMW3YvbggKdeFq8/Tsd7j6mIRLXJoposoXgR08ZNVJluxDxF
gk4vZdQ+1koIrSFbuQRcLK53WpT6WTvxCrx3PO6JWvcd8s0Dh5wBLuY02mf+dBXK
DiMuQrut9MSnVe0AbtCVpT5LTt3BeT2GOMTZW01MEC8W5Y2sFMQ2V213fJYPkXWd
ikFUKcUJJ/B5OyMPwyCC1x43OhABSw5ina9x/rvfybyZ5mmgoLRUskefYjfJ+5og
OyMfHuIUHIj7Qkqx59csAptb6BFrnIuvTCXeBCzvdDE2PcVRaF9Jk9vhtKkRRQN+
sxL+ZEBYlHDa9OHeVbPaCMQtapPY3p8Z32F6sHZ4SJMQx7JM/2QqLGhfaE+rgYyH
U8gg8S98WQ+tpOSJ25zP3qifs/X+huFoZYQi+edzfze/heNPCO3lO7MamtXmqPI0
6qj2Y2RpL8sdc+1diCKi1ZwKGG/5k4s6vM6o65tcgstc0rzIL2xkDMKQqHqAJMYE
s56I4ua8ij+sjvn7IRIvqa7bUe/FgHmdNy1ff/bvFGnnQf2LQ2afEO0eLlQ2Tps0
BZSrjsmIADNw7nItIFhbQQWzi2vJH0WICzzQIwL6/f0XHlOg7VdG3Owwwe9fC4r+
XbxbJD2ciYacWxQb3xk84QSQ1TKCt3qpo42dKwZUzQguo+rDnHP5T0evzH4WfECw
LRv8P2Edc0Re4WKIZlbrPyq1JNObJp7e3mCCI/IjZyyrPg+401lnqK29mu10qnZo
AyQN40HkVb/FINEVcpZwXLGPVmESCdewPbJsE2PiIIiP5ZpYh9z+DkaQVJlrceMr
jIzHy9fAcZzu4GMZCBsIOt8UcJql+ODl3hXAVWllOAQAaY9WimrVm2bNgKIlV0Bb
de7wXra2K9L+GyMSbquUmYW6ACbrwR4I23RCY7jp22HwMClqy4A9k8xl7Swhtgai
AzkzEFrxRkzy6WHqpCWjeFgOEhcuuF1qxqDSpHVGIad+z/tbgtdVQyYIuISlX3h5
wGmaJld1lwQ45AZLmBQuxTa+oXWPtLf/f0tqwJ4vJcQrviBg+2LPyoVjSRq7crjE
kuoNcty6xDvyov9r2b9DUlOSqVvjkQceNvF97OjaKONe/ZCMpAFAU8YhTtLdQrD7
TUazJEx7MhbX8i9sP/Lz/A8QVfo+78UzQzQQbVxk8KqBNcSrEN6X4BiiAx1TdzfR
VJqWQVjaxXOw1hyRAoe63lGuO+mDLS1cw/3kiKGynZt+6LaPYAE3OacyIfaMTjEq
hpF7IpUO7+nOuTeQbC8clWk9gaHjm7PtCAqAkRqBmCMM/FqNYcF3kXp/6JcXoiNu
s0j+yQsGfwC2LyYy3yJmYARhXysxp3Wx0HiLYLE1VjhrnN1vv03sBDGzmYr+IiUz
Z3E8C6E6RezM35BmbVC3HNO2PTbeIIlMRrEjIbJoE+1BfAlF4DAQ1QMAUOBMiJH6
nxJwan+4HAv3SLIMOfyHXPFWjS8ljpGOz+xV5H0pmd4NMQ1l04dXON6tFT1NBiH6
7Pi4pnk5Yp3BdJJOI6+XgIsnIgmai5k4hY4xfJ0ptTvnja1RteUjtfAQi+axoTXy
TIg1AA0nNcmo2h4LCcAPxKMzCE5WC7mucox7GGNV8K/X/jl6gHp7ZZQw6W/Baadi
Vp9CrDyLc61eZZjtDeOtq2yGCEnhsHN7H/+WnRJQaLH/dILf8wXXTPXKdZW102mv
jgKs4OMvFmdXUoRrEwKx2rKJdBSCNFtmYTvTzxcwZgcarBO2Yp/tPdrKYm3A5/JD
OGAyT0eSf9Fwq89+T37sg88SQtswB3titlaF9wAt+S4GwrEUuLVXuoTeKLHw/62y
fYSOQrQdctanV7uFo4ZxWQIvSUmTUuEm7rcIbIbFp4c6ejYGlIKbVqnHPqCyGr8p
iVHHNdX+j+ntNODViApGX2Plq+fqvDCQuw5nPgMXtvcBDprV9bJKzQZYQS/1zq/x
f2vyVhHiDFivry6z017VgoKGzXru6lJ/xOUIR4pxSFOh5xG/Y5+c8FWkVnX1Iyz5
UkVNxeM6f9Pyaws7Dbodao0jVfezhep+CNgAqVJoLydqQCmMV5FVJg8LmUipEeMK
9C502aDHhhHSL/SYxqD8Aq83qmvxp8Itmky5jbcK5GhlLX/3rUpiEeaAYRJjl60C
XNnk+03uKfGe3Cbmfo7UEjoDHwM+2fgyVlUJ1T4aGIwGSL28i0lP+5Yf1FOXxTBq
UJ8i1xoL2Q6ooma45i49MeLNHzO4kdu3i9yqtG9gqV2BIII3eEodNXVi+uohKDjU
ub4fAeoerZP/qcS7bDzMaCvCvkz1Er9RnUSP1Z8o3Wm7cs+sppGb1rHTXTEgMhIy
PSknUBRS3Z0IKlTkmV57X+ZgvfoPpi/0lnFrHkCRmrPO7HCEl4PDebrhbZATV9MV
b7WEK4lwuOBj1cWZiNrWlD1BVDq1kHADBD7wxWBMbT4kCNRL474VR78GDe6EY0Ks
75IN8PG1Z34J3zRUEZItrqnt6aE7L9n8UnTUYVMRxJoh3cRDDI+qHuTM2eIzAotY
I7XLstJflDJFFndaMYy0P8qRfoAs4XecfuEJZKYZfoOP7SOMPH/r46O1X7k773C8
uNYXwN+Mz8CGj9K/sR2LwO/8G7kQQIDItWvvs5/5zc4sEcBt2jCciG0V0+NNnY2a
LVtKcOvzSrquo5tO8uGEQG9QaW38dXV4uK8A+f8j1FLFvCf9lt+RdjaqBDlCwOII
gFsHBDN0xTt2dbcdf5idBNgprYhxSaIajKL62yDPDmjA1VLw22iuYQP7IX39b7Ii
IU1y4twQ2mGp+CYsJI1SlKdln2OmthaMVmCwRXup/hFEBiiBXb+O4etVp4T4vAg1
lx3J+g0s0mUqoctDVUThOTJYoNcpoqdSTP1KyBsnC1MWidNOqfMjJIQSQQ8B0Vvf
+129PPLQn9dIK/KCjlOE8yTyd2bKLIWeiNrb8y975/BrCY52HwAx8Wb7r7IP0uzE
HJaUkiB75fSz2kaQzkyxBdJrRq0sT4HWrp+Sxg2F37YqfNjNURiV2TgaHketZLti
wjHCOC/UxQmIjLgm4PexhOpH3Hg2/Rz+Bx9BW7VqzqI3Wr09mu9H7ClCSykYqOKl
UJNzhacpOEyxUujhhm0zz+uF/eleGf5uXB7H+xXhHINFAK6ABiXWIYPBRooBCwZi
pYQt/rAn5hcD1CZ47LIe/9IJlkpopW5++pPs0NXSAndQx5BOpHkf+nwud/tiNDBV
eQTxbMrNYvevARCdkX0yUZeBQwHS3k/tssE2XdrNKNMFaY/giUgUfTPptnxrsyIC
D3x6fRkJSza0VoQlZhtOfXPuVMeCfMItDu9dOY8LYG+wnzzB+V1D6iaTgEmV3MZR
FcKt1G169L20eTII9th4jrDOYTXUN2SMfMGUwz0W0eNV/IydV0QskTtgzWCED/Lm
fWq0SKMtJesLW+NDGctk5PGzXYJdRHPkXUhy00MU9aqz3PIyHYuIzEjfxV6j3wL2
Otag44kOPV0p8JeiUp3cosq5prXNeTNirjbJyK00r/UIEEIefrc3evinsRwLfQeO
I4DYjkHvbx7sHjFfpmyrNN/zZLW4/p97N7RPomBrlwPqB3NSXyVe5tmVk4jsDMPE
xu5wWJcHB909p5Ci3mKUqRGXz6tUQpLrVzI4RZ2C3/YPza17LIWj/BLP4PLZ8ID9
O8mAxwOP0XtZ6dFj5QoMtMlybIwbm5qAR37x0OQgSb1z8VXslrIsZUYf+xqisr9k
AqpG5dRxMGlczcmsFaZgmNQCPahzxgCqVtj5qI4A4XKeaBN+bEknAOQxfz4kD5E9
G2b+NNHLU9iLyIkj43cmhOhGay1j4pQOtLjGo3BnMrVH5ZpDfDZkAb3hgY/LDopv
MRTutIZwFaIhMjG4rV3Zpl4p7Ix8zLZn0oOTvCGnsLH5Vs4FW+BiTQ825kLkal0a
HkFBvwGf4aDUi/hKT6lC+s4wexPoSPDggOpqm8xBG3HahVT+V6v0Bd/Od29N1Bxl
+aEdYomFLJceiyR+XIxXpatvAsHK/UQWeRhCBgdghNqWpkSmH2M6vcz1wrbltzfh
0ky3gt8SIYB77nD6YPMJ6lOATOqskYXwBF9FFGiPafkULp9gajEejpphB9VayHRE
oP3GyMoe7+OBg6HG4bB4DB4twe2NV+mypYOnihXrK/fcoNNlpfU6Asi7X99M0tQc
8qcO1ruDcFG3XdEvlYJG6MVKpekZN607mVxWQns7dcj3f1pPI0ZDh3dx71X5Tc6W
wKe2MYJ/Eog1/AJlvJ23MPB4IX6UC2H228kf72EnpbVsA2Eg6uJQTZbNm63vsKLg
lmA+XraQ0V6suOjVIJh1tzNu/E2vQsJSxaz8K6JVIuP8ag09QZGwuprSVH2v9+4R
KWgD7qg13zXh+fmyNtbw3qxNi0HKQ/MmF0D4huQR2L6zKeXFmxaefUzyFKMxejNe
vPDLLs0YobROmUWppZas00gvZqpu8odOJt8QLI4QzWpGJxL7tvh5gcRQhbwn24RH
Iv129rdl7gT2kMlkXDrUGQgEV42TMmELL/op6Ej7n8tDFDE90TG0k9OpxWHAax5U
VPyJEDGh0c3xvqALmZW3mB1mvtDqHc0cC5b8KbQh6XPS3oxPqEVZBl8FEAJaoOrk
Aw84PsbiRyVlZxSJFZI7seWYofAMYV7as4l9qTwEO9OUFt1ZlHsxk0PrSCfS+C50
8OqrWYn8/LqgqDljj1crIK9PmIO2qIvMNnys5fW6QqPUC2QCl63EhtJTuKjhBrfU
228SEy0TEDw4vYgbLpDARA/q/K+qS8Q3RySgILabDkhzz15RlxR+AOx7c4x9s4y8
vsMlA65HMF8765N12y17oPr7FMc7cSHcQRCKhAPA2xNV5P1zQjNM5i1p06Gtj1f/
jOmF9HWnKCG3MxNpCO4j+Ns2GsPTh3DvyrUpkefe5WiXLMVxL1au6EywRYVyVG5S
rsTUXtHQ2mpM+5BessQuPAEohpctRlfW2M6VtmBn6P/UWeWGlo143CtcPkCS3+Vm
NMyeYrFTEH8DRSpciy4k0JbNczYpqZR2yhhN8c0LsrpG0Dpl+XFf8OBo5P1Hr7in
qizTtMYCVXma+pyQzHkADaj1ewNi3DQrgBWY/OI2lwCBIDz32e0s1MPZxqqmeKsm
MP1PFS2tkrO36uP/NbMWoZsO/uoC+4/rrDk6s89q8dP1fIwsF71nbqsoAKdh1oMw
RXyFlP+hT2Q2CV1PtVpD24bmvKIymvcmI9vjibE4cv29gy45ud+mjse1OpNOpu/x
81s/9sXOvJkf+AzEBvIO2ZXMbCuddM6LkkQHhblBSeTaTXrww4MisD0PgpKH4jUb
Nozh+nSlxruenps4dncZ/lvgPpmiBvTTxrNbh++wnRBPyBHww59kIssVAE/nLq1v
ZpsKO93F5uybAfsJEhi9y5Tpw+W14xBS8iA0W4kChlC/ziKNPuClFWd09omCDo2m
w5Rxx4WHcU3V8BQYBq6MPya1PXKNLHJIZkWRxLvko1UMV/O4DmgPxZnIU/T4taoV
5b3N5gV/PNUsYqjDzyy2YAyKlf2v3bPHPLNSzsrj3jZRNaqkIOU+/oOPeUqzv0e/
TRV5+ZDk5Dlupvco9acpNH0IO5DADQ9N5wIaWatPEKLahnwslkjgVp2F58PRa6Bc
dh42QiNea0f1N8OpSOjMcnt0Os/UgOgJj6cNXB/e5qnXs/R3XlWz1MTUsp9CZRzq
N8s4qvWHJjKPmuXvZ+Jf9x5BJSfvTUtXeucRI8qysPdIVyjfLPi6nyr+hnkknC40
etPTKL5wabskwNghuOcVYvbVS+AZPkUcu/ggOP1tW9I8t7Nh586Iw3qfJ6zu564o
GRTbhlQPJmKt26/HZE7ZH5e73SUBuo/sEzrJqwWxanBRixT+sQt328WqvCnIWzok
xmdQjPjZ5OAwNg12PUDydB/GEyBEMW8VdoF+ACQC3eNpN/h++RyVwmLoFPaEWLH6
um3vnWs/XYFqg0FiTDwWxNlv0HoUGOnVg/7k2d2/t+4qmkea8vUpvr2wcGSmZ9Rw
LAHRjhVsITIVnP+rmM9XraCKyfBcY1KVSt1TYpe1ZTLnjyuUbuu8f2VXSKyWgx+l
8ci1JHotQ2h3QDn3si4QeSfXZ5lvsqK6gOLeBt21JA0DdJcgWF0DE57MpuOrFhEb
Ak3X4WVeROHiMV9v4SnSOH6O2YwEKHXXBa9kaSf9I8hud0Dp+MywDlgcxiMs4c/S
2BmFfichJVIeOvqrm6g+8TMUX8zAQnaTOWgVy3MGc1XG6zAIwWQPJXQbhGD+Pm+X
0JRUklDVbL20BY27C68hn7XX3cK00V75Cmcq5C1VUR8mfktp5ZaWla/4MZcA8AsG
ix8QTAw0vAFjskUIHwbYwWub/gu6gSCJRYDiirPGYHaJ7gtFtw37qhTXfHwevRZg
8jhZfy/srcf7qJxo53sHthPDxWUbJwq4nJqcLpVG1/XV0alD7AChXlYOUUgLkJ91
kplGEx2j/eZlgDk4LNT081I1PbWxUXc1KwtL7UvIUbC+uifU08RHuINC8ZSrw3sy
YQQtkX7RBXOI869x/DmN+SKaL0TaRPjCKqXKlcbVKhhaUWKp8SBS679Pwc5mv0eX
9GRbQSse9ena04zYqJRvtiT6EW4Vgv46pUdhcCE+p/UtDLUwn/a6c+DEW36xBbSt
qTKadZGL48y4G/kzk7zOAo/aoOOdQoT0lBQ5uTCf5zhcTAyDFZ2HkZjQvRCFEIYS
JVpW4Tw0gE3FDYQD70C/m/xS2weSD6RTZWb4SIoAoCvwIiMtom+A0fNTKB/CeDYs
92hJHRkmbQqQoJHUa+/AYXa4BYgRncqxduqrKfOPVF0ecfbzFKoY3lOJEB9ELtsn
xjzh3JI64oZns5kSd127CB7X/0+6Xt2LqX5V1LnxWH2hrx2lomOFw589AI0zGSdq
Inp/MIzzk+JOqCl+aokY5ySXqCnRAJ5L7Qmq/QZI6OuB1ZAQ3wsIMyqlE+Xdg6SF
FEoTEqVgLe4Cjwiq0RRpA/f+R3jbzeycdW1CIVjRL1LnaCVyDFpf0oEqMF5yMi5d
xhiAwGuYpmz3QipEavfUeMnanyjvoR2wtI21BkMwD+T7LQNb+M3E3tMhB5gsofjs
KwUvjgPWhkVw5tqLlNMbVDOVQslcjjZskJYFmF5+DXk7Q7mYDV1E4A+My2bcS8wy
p1X0Tkxe9uDXxIUCUp60Jub6BfQ2laeC457lBo9Hoq1a77RrbOpG3fR1m1IwgDDZ
tCeBNkNX7HyI6mzQHtzsnDhNQ9iREDEG4vlZttLy2F55kJh8YefCu69rZvMLMwvo
vqBtpVFQ8oasc5tUjMvDZ2EMK+disHSIcxnSKyKmt/P7DdXOKXgQvCMlyCkHEsqP
KGg3vrLwU0Ee/7YDiG9FuQfbmCp8E6aT6DRj9MAyDPPjaqRg151p73XzXiYcmChD
Ua4O1ol8hKUAcCjw6mnc4fDSaH/VqtNDWhFMWoZ2x2QPUiCnjtQoK81R4hnOjevc
8RJMVp0GG2Yp9zO41uZD8TmKOvem9tduXI+x03d1IKZXh0aJWK9UEQEZsMUcWUiE
iWUtSK8hmfUbndrnWQX9S0aboC6p00d5d1z4cTm6vbFwKMD/wiCVDgVTm+ffgbUM
q73dzaprLOeCedKC5/Kzi6B2YoOKqBEt6akAi8QA/A+EzlVQpDx1pjDCunzLhJeM
uHI6jdpUAlOJcIU/iosCw33mqHYL96TkRs/+O+vdw17vFbgKtyEO8I9AdwCRnRXi
t8JI4C20hAlWsmg6gwRsTaJ9TvAECtKRiyTMoS1psgVnB15xgjKiqVr3U38qhM3c
NmaMdThCKljqNG5tUW862cYoKNoi8YjXh/TZQMBE8HuUGDra56moH6qc6g2C1bCh
zlWkuGD2crINQDo0WHZyJ7yv86LcIPtAdMEmPW7zFSJe5h7U0mPAfucFfC02I9DO
jyHWG9Iyc9sVAMaxtlosoNk7A2nvoPr3NN1Mh9+Crm1RhfFHIMG7oUI7zU+QGss7
RHBYSkBKQiApdVOOTPpY29ayQJmbSRinhCG1ymUftJKi6C8DSm5GtXZIVTvIhPxt
jVCpWmUgPISE+SUx0XoteaVnxj1iTK5gjUXUn/a8hdY1o+aNS3Z9LFMXooz9Uh/c
ReqT5f/hprCnc5zsu/Rosv+02v1b0gQ6hNJNH7+SEGqyMMBkigWlBnuoKCMBa0Ox
XLZatkUw6+T3UJ0gxBCekDDU6TA3raLzid//mpeO15KKDCONE7paQTqvUQReAeqY
N2eBxkwR1ZCD24rxsmbZl82CHSR9h2l+BCCdiX6HgYZOQzo0KsfAt3EPEMEK3Csa
QzxeVHB82qbRPTJAHE5ybgpCWlqfX+XZouOeipzdFLC5h1tgZF17Q0CHwtiEnHX8
O/TBUv9Iz07YoT7pbRU9jOjpAT5S0OJm9U5+lnbl7bC/hJtOL4Q73f227daHVupj
qVBAHrQhVCgSXC/xEK/fGOBoNoQ0wMN8PCRBCiV8AS5EA6Sw+DgtK0aEUGm1qABg
+hGCi+OLk4aHVZCo53c7EMAzGZ5JXfxAYvkiVGo3kuw4j8c6P1NpeOL2j6PPqQuF
JaHi32+HpVjVMTRWMjFxWn0bwfPsvBixJ05hk0Jk35tRyGIUPwc5GLqpInbPr9xI
RoRcdkX+3aeNaSbL7su0W35Pqdcqyazdap5PNUfKQEjNXs2+7T/59SQbgld+ATjz
0lrdHdStDiwxuBUz0E4Yi7l50ZcHsAZCUpVnjrV+6EHBGtn2MZFEcMZ2xlZaSokm
oltpD2DxXyVMAhdWEyblayBrIVnUDSISy9kp7nWZY7fuezfX3vuWIDuqA6UuoSEg
ywPJzJf/g/ijjLkhtoEo5HIhJgX3fKaEtLsR2uzvnb70CVz90XnLx+D17JQjWyVp
HPjLkydD5jm9P/zRsPAmT5PxL938Pmd78VQcxP6SLqEi6JzNRlEuesE11B5O1BiL
Z9TUEwXhxbYL9j2z4tU/Dqu0QnEklC6KRx0MpvRVfTOaHx5bClCGw9RWjS4lanPs
LF34ZkFsAzRG5Y3wTN7TrdAKvWJ6odPyeURBzxAxVa2aTu+PHwJxs51JxGUWDdxe
9AczPLRyqQytaMoqr+vH5uGAnDgNq0/MNAoLuHVLsODW2YKn/13TM7SuwTWU66cm
Mgl3nrNwDpyjq6AYP0p+a/prGHGaDMqfK4h339T/qmnLWyITy/KNOcyv+U/a60SS
/lXGMRjS81v/OC3WGCb6WjBDpt0nNbYi/BMso19G8Nds4sBeZ1X9uinZlL5PE/Rt
rLsFrdWVmX9qoDkqMhVlmLpFVQkiNeuVlCx4ZNbb2PdzzAb0RaivORuabJOqH97j
iPwWwk+Zg5/WOVXK8JKJXDrfkPfDhVbSZTkhRyMPX4oarp/LAleUq5VykEuMfJ1j
gmSkIljAjkCsWJmfxUzkSuhmhsSUoyC3is9/WvGT72w8kvsrdUd5NWayPgvUxwhK
f4eebZJP/ltVJFEYmB25uN/Q39e9bnT4jY3AzYvSArRQzaQUTTPZIndZQznAG3b8
5b4MasV5U6I1jg9EiX/Qkbw7McdMUnvo21+RoVawpDK08Hp+eSIOhLvhnDj7su6l
KcdNOZLYacFKVWF/VZvHfXxpcMitIle4muArhHgEjYmrhYE/bXsN35+9wtnBdBur
fMtPDyQYxHLqXEpix/Eu8tVlI7HwcpNhLqba+tGz5McZJeHFTb+MmbcxJYlErTuf
ZdjBj2RRE7c9eFx5aX7lRI7znyXG8Aphl9kTWJ5TyMSvfoEN4duDwznbd2OAB4NC
z5xGoPpB45oymdnc1pnjokLodOdWexiVaQyWBmSMwviUrHdY8uzmv+cTPRxi1tAb
Vm8hbFlZx+V6LyoX1F4cEeTps+Ih2JyCObBFbOt0tBrgdG0gIaKYNxchokRh3cBx
YVmhDhZOdWtXjtKCjpfWOEltmjj7pptXNboBU12jNMtwasZ3Pq31X2IQGzJFUvmQ
st6MkfG5R8ffhvyThycE1Qx6aRbOb2UKfBlY6Vg/h0AgTD0cCkGjsc7+I9a/rhN/
h0D7OHkdaWzqHkbESsVEXW0bPMgvMRM5FckY4gqXoPHOMflmUYiPfZdBrQqdwc7m
/kbka/5H00/nDm47NDBX6fGvAf59MaYV0fhvQKg+LmzDlkwjGT+QMF4xzbz/VINi
ApWE7KZVTvy1I1rCdrZMz3PtLDhwMfoW/SpbgVKeC8h8znyCRNQK984A7FoO76EO
D4CYlINxhN2l3HVy4D3v50LBvdD7lLDNJC5/poci5wy0C3vs8aRGn7ETtU94zp1w
w9n/VtPqwsvBWr8LRVmjWbSFUgBj4IQtVrggUP8FFZMF3E43W5PwagF8MUduufBl
oB7F2rbSic/UDbWejFZnmtINkOstDvEV0P85moTDGF4nhRO8+TFFCKcBkpB34VvD
C64iS7TqNNJ4EX0HE7ZotWuqEZZMq0IOm6FvP28iwluDfCX5DLCnbS5mZN9rALn9
i+SqpcLopzS+AilcZRW2tHzveFKf1QZqP4BkvtY8oWsFjeb749auTcJC17XIfdKc
mZOPcGXaOXxcz98aHAB/SByVcwja3yAE6SBN/hlcwdEszUgeY4Wdq5ySG8vQvzuf
cdqIrww8fsTzW4Wn65Xm2xOEKn0+/gszLD2RHZ4FO8aoFIQEu9o1A2OnHvBzsMhk
RVEg9bXJiEQ7h3+f1P1UEd2V4GB3/zk+Kf/aQZlrfLhQcFaxY5Lm0wTtGzFCqroX
Hswc+PY3axBVGbh39X55AdXY3MvDC/lV4CWdCfDoqSZjPcvSua1JSdQELZjqHOQh
Qz0sJr0XvHjAxQwRHx12wkIIL9D44eDMoqE+RL5G3c3Z7iHNGA25OKInzLxdQBpe
/r1eR9VM5RIdWKsJDRyg/P8Bj6QVTsGx1oA8FECxn4zsyQNkOZUlq1dKjO80n+ql
LMY4PDX62H1IFfxLcMBTDjUVrrTNIutV/cFEiTfubyXeCBoy9/mQlQlOp5QCQQkt
KN8Wdz34RQDmbP3B8uRA09sNsrMAc5PKZ7DktTLnlLU6tu40a79k1bFba1ShWSeA
lNrCKD+HPULieDyttJbayaftuTq7hGNnVzDFRcIR4p66oONSJcHtmjAOcRSxYUjz
eJ+bBzCSrITymKIKKgw1MxU+skBsQD+wmI4wmZC3/CSqJJ/eyeVIMDveGEKlyrwJ
mcX5lRsSjWKpxmTYNGc/dZnYyvpDacsnXwGna4RtmGuY75WoVhf2AKO2+kl74Beg
POABmWb2RJvKYZGEUjA6WlWJ60qv6T1DQQQLg7BS3r3UsGyfh5k+SVxlIY1yZ0gU
GMfD6IRkYCpfGj5ljp6++zkxniEKzq0WWD0F/BpruUe7klZqPYER/gq4BVGIrEBt
3UyXLq5LSDoNntYP0BgPZj032MGAxo4LwkY4lhWmlFumZWEjnyNd3+WUsBKaPc8Z
EsGFzZZ8WGaS+bhC6K/w7Je7hFNXqi6Wm94/DSXa7J1LWihebb3MwLsHm9AGsHC6
MNwMX3bS//oyZAe5Z03ZQSt8uWHhBgNd/JrfirkY6zWjfmV38UchLV/9ThiaEGqV
g5P/4cgt4PKkyvkWDqfawqiPOhUyo2NJ2bG5iRYUxjINb/sCNCrKsqb9bah3TTM4
ik0WWZhfyXGi8ah1miCStEtlQvdaxWmbhBGi5ON+wGENmjSe4+A4QYvmyUtyqCTG
ciU3W9oJ9m/j57cq5tr6ARBLLvXNT06e1VX7i9px99O1iXd1c4qGHBiakjnJLDsc
5FTz5+rSM3UkDc4bQm6w237SuQWVQ+F1klel0nDVttsV0ZYBrYfdMaBPiiPCmwvp
F2H24NFFABNajO7k0tSbNiAQLVD6t3MgnSeUMZAL0fh0wo+Lfpu1Kcg+RzlIgEfp
rxcGi1KBAZjKf7/FDsl5ZOnUV+il1U+BZYtXps7a72+M9YAUeJVw/7ypSGOBnW4W
N23jqGZsy9LX7YLgElHLCXhO+i9O7N6vLmTanXjuqKYVjitgVu+vZwpkTPUVOWjM
aCf3Q3srgQL68nhYypDl8py87IqywX6hcKMMLmviZ2DMa/rMkbpeq+hWsAraft/I
Ccp6dr3Wr4kRXG2+gcVtkk8fLb7ND2X8HWFa9zwBHLIxyAj7JxZyoofwkk4Fqwo2
LdSiJPLnUm6747GPItX1Z1/F6rvsG+CVsUopFcxYF2FJIJEpINgSvMNd2YmnUfZV
8wqip/ayszvvTzifTh06Ys0MTw5zLu9kW7pp3A/VbKllywcgVJx42XkaAN3XKFXy
35UijPZGFJQhpUd1oFhF3JLmGU4sxkeXNwzYt4/e3cbJ7ngWVQocUJicQfC6epyw
YDa/4JFYjom1pM3tyIyO3yeAJQp1gPEoLLFX3CJ1xOUFaR38VZF1v8XYEWX4JAew
zal/s551qBdV7MoLH9Eme8wAFEwMoxBtcbRgYwbJXfj5DibxF/Kqys+EKV9dD1oN
yyCV6ZqhgaEJzi/0M+ocrV9j0sC0EIorw4IADDM+Qp1y7rHe2acSDNFIXYu19ZB0
Xki80kgYUlAglfGi/yYDIIJlLEkbrODeT9GryTiXhpp1cVOKcTV3ZvmL8sNbpv2/
PA1dxAEJ2QsvGjfj2S4cVvPyiNiuHCovSANelo6+OUN9r0B2Q7U9FJaRMYo0YHRf
DQrCvtP6FbO8LHPiIcpbVD+VmusN9jeSER2rEUnR1+qyCzdRr2+4hxygaW8GRpvS
jwhNPfFoIuFCByR5CGeLiMaZIk915EuhXaRUDnsXuF61lgPTTml3/haxT70KYtj+
o+JNwR45gsHCd1UwMvFywA9NxjNQ9EzgZz4V9v2Q5YVQ0e3maEmEb1HX4UzHfXpm
vaVjda+KHlbomxliyq59bNsb/8h95ZH396TFiwpmXOqwot9kOVZVFMpa0YoP3XB0
y5MtlM7IX5mzle7Z+6BJNbTszcTJRvU8E1tJwASss1j5bwf5OMesS/Zq9hkG2mlE
tqM1TjJVM1g1OcmI1xGL0doB5qaS3PxAR+jBFqTH6WNayci3r16H8X9ARoEitYuX
pN33J8KaIVEIrXZWyl96Kq694sPqIFc1UN3MsyvCOvciwhaX4YuKvIBuD0KxaNPV
E6KQNcE7EJ+04K3Ox+JcRhebLEFA8O/BFMU9x3NdcBspirwxFNrpuIZPKKgevJH8
i2SeXtro9up6pqaXhh8f9mr0xMcozb9J6GP3SbE41qn4p/Nb8vTCYEGgixWkkE99
WPZDr+SFNDwy1TXjUXrysyiCDW8ZXnglUxuLXOcWISFQ9WTjexcRJrb5nk6R1ZUJ
/7UN3tH6auYVJPAveO0DVxyaL0EMcP3Oj1fDF6P+uRqPsEsU9loaQ5bKSX2Ek1cT
51evDUwwcIXmgumOZD+Sa0TERo8OPFMImdEhv62xgpt1OIaCXCuDhI59ZjcFGCkK
55mHQIWNzFOjY1wAJAr1MQL1P1HU0euYYgNfOEQQmNxOcBOmB46prL9UargY5TI9
PT3MhZN4+4Xc7HbGKTd9/aePo6WYRjCRNUr9QdtOAMM6ppZXSYkxC/5sUQZpkIax
xWK3wfCGAYkFV0jj7Ra0Ole4Kcp9z1z/V0f4WapLJ8WjF9P8TqNGIQ0/0swe6rK9
LFHvNVAk2KbfCaf96qS2RAb+xO7q1dIrO9rUAOqzyG07EdScf9s0+rtW+F2iQQ/k
c2QTxDWErKXLGgVaKWYzYmYSMhe6LqXr8aeFs/x2WJ/9sfCL66nx8azynm23y193
IPg4m5F2IMiiFHEg+g4qafN0NKAe0lBrfhmWVI4FCg82x4FohtcAHvZr9RzbKDPs
rui08FgsGT+QgDucw7eANsPEJZ+LGBqHh/dKLsdNWjHNnsSu8x0j3Iqeet51bVVb
ZWdbBfd5vOqdK8ANX1h/TclEmsR4faCbCEzPOXNzrK2vs7Ndkxek5MyBtNzp9p0o
U/Su2OKpwrGsR4MTZhl77Xr0NHtb8VPbbKVATJ6mAIyBkl/g2XfDaqVP52X7SJ+a
bpG9z/lcwYmU1rfiyxM55yx2SbRYVtK7kQr+E+ASDOCRdpqHnISzJEzSMuymf8JW
J9Cssyg281dQh+a7KQQd2Z2KsQXmhn5eFUHnd3j0tm3A85FDhOkUQXFdqS3/8Nra
FZt71TH65np9Epl1JgLdm8YWZtf7xaleUmylp95OHFdMmW6ehijId1A8xw4biqzi
nBCFTaW9xIvGqjOGJ0axN8hyOrwjKwxNWpLvKCV54s0uj5OCoGCpEirGyWDEwWjr
nD4O/9cnQ3UNS+eY+wane1ISCCVt9aI6CXjKw70onEQ0/8FpXv6Z0Mtmyx4edGIW
YLRCO3fBmsdmSryfcWWBFE/jsiwbw3PyQDOyqAvb/jWvFk/7n5hQC/e0CP+haoGP
djAx3zoc6/yDh7Aj0h0O/075hDcHp63OYYFnAcLA2V6wBBby1IFfFDHm/8tVyXdj
LYpxxAVB00Yqp+eoBI0Bwn1zDqe+yIuNT89zXohgzJSag3gcVW1p630e68+0cQgD
MAX6EHxT2KccSn2bxE62c3t0RXlHmAHIDdkSQPA8D5oRDwL+VfMxY0uahEa59J2h
8R7Ozy3dH+/q+UwFyeieyN0cvcSoh2revbG29Oc5NL4+V73o8dY+NMZqeO4UDhOR
3oe2qUv42oFHnF7TyXfQ00QSirU3U20oQnvVKxAloXtKpN3tlK1HigLZ9aCA/Ns5
Ix02WoagZO7gy0MWxvGnpN6IdZ2W/1n8LQNuHZ4gAljc60gvfwYtbGj9UiQUGA1I
ipkSXwh+Nv4VfFCAb121Iz9gW/zWLkHYOm45mDoB1hRnapE8+kDfstEYHXt0zf8q
E8vZmdlHD898BMV7tbqQ1WD8DJaY68We0OjCojh1sUM2FPJjvq7OfJR3jiak1UMh
3UY4EwsgvLrisrxJKna81oc0q45kKQA5s1k9rnU5g8OaZy8uZ+njyJOmBAbmw8Vl
OTheT7XhZWzH0uaTNWe4IX+uA/6c3W++2S2VWG5lZ+stzs9FbMppQJQDvnFrRj2X
BQbHQlIPb/i1ueWh8/0wUewiEqEZCq9z5fhEV21a9Jo5P9ab+i3EefhPEAbTSoSu
inEL5McHQenl/QuQo7nZCwuYpDGQobSwS92f/KwSzGJU3XUmsmRhQ4QPIi10SchK
s2Jpu8TU/9PYz5JaiQNPqVf9clSqSiC1d5iFABwUU2o8FLWw5bui3+bzMpNfAOqq
sL2IyyuB0S2ZXFssVGQW9kOTIGrzfs8KyOyPrqekhkdrl5eS1GL51EAtZJHTHDH2
9DD9zMa0HmFy86eSv7bL78AbfJ4ETJZAIxfp/LAbQpZte4iUEFZ2geQ8k1TNKvLc
uMUDlWMPxH9d9SaHHDuAHFddIHAmkULV3/wlhIQwhFNnd+UzvtcJQvLCmuHDh7Nm
HGh68Kjvp+no22ZNQGEkwLab099ZWSAk/vRnYXAbdM0hvhpF4F/WaRnoB4nq6Aks
AK447F5GzJZfeCQ2V1tPrm/j8O1vsE5g7fEMXf9NxJIPq6dQxfKM3kZy83gTD2q/
fEGyK8abIU4pfGOG7/jtmPrMTUekHcpN/GVCYbt+0Joz0DgmaYEMBBt6/6ejMG77
BWKdEvTt8vO4uboAj4efrzXAXXa09FKMqyDeOtpGf+T1i9CLkluVbMdVCabT6LwJ
2fOzrbxolVpoEDbd9bg3MekbqIETYSa8aeQk3ik9H0MbRdR960Iv3j27S2rkDy1K
RAPP+W4bg4qAgPFPNdcEkPptXRns0IoJeWVWtYwpyjcv78X7+6K2fBOLaPicK9NJ
R9qMTSlsGOZhx6rDb14Ve4dZRVaFJfL8d7lJizr3LusU4E/NZytsLjQLBySIHu/t
Wdg6bVN4bfazlqaCoMlNgUTHhMimc3zrZYcreIPURE58NN4NkrzkfXx1XB/T53Le
KOSxTg9ZQp52bAvn/AfBwu6NrvHp8dWcrD3huf7Qo90fBF4k55ysvXlDNx3Bttav
FuNGDIqxfIJqbN03q48dUoccnA87k0yEf5qLja5OoWHDbbOQSDhJtEFUDINkPz5k
LnPWWv4xv4zvgvXGqMgeNcdTM97XHx6MXdnfZOVl8HHPMD6fh3w+CxyhUFo3OQqQ
hxu9LhluJOfT+pNKY7F0WanYSbr3G3lzvjHOlkVaah1dE5kOe8/U+BEAoNc7mLbK
B8hKFsYnmasjan3j8B6UGCjUI+sT/Yq+4aMwy6sOHo8phOT5KsikWlI5clCBztKG
mIgjsEJnJGbLDdZHe5MFF7UTOXIiWDdnXccfkTEhsxDpGYab35HdNMOkbTymb1oB
W3rVio188ThtiW5u4zDNAi9U/NLl+fq7MoN/DN4zKcMMzCfwRf6jzfT0l+UENB29
K74oh/G2Zh0AzsMv3l9AEs585jW5thxJgmfTLoL935pAImnKN2TIaV6224g/aaHo
IXbehzdr1QeZDkQTr/Mn/F5q7+0poL+56Y9n8YZWgq2YfjR3kWq+FgaE9ZU6iVli
36Ojli1K9lITnoU7FX8Pr7fU6NSxVZmv7MvRFEctWLAFjUpZoMouESFxsSuY26NO
P9jY5spoyNuesuiqYXwyxdtkRNTkGw1WHf0oT5FE7evCDuULpaNdN7f8pXv5MpTX
onkAywhnEua+RlCXAx0+mL4XURtnB2uQy14p2mdriLkq2eXWjZ9kPufoLXJt56jU
y+zwNuR2B/RY23puNWZP/ypU5UjXUjIyszS7FcDd/ggk7gRZO9iA+Ewc0UUXU7wx
Xdlp9ZfSmx3vYKp9Zc82rH3ITELCjQRxsKMk0jPDgvK2NEKUsPJcQ2oDCYvuIz0S
NJNcNEE/oEIW6zWWvN8RW+mMLCfeoZTGDYH+CQqN5VJkuRRcrjEDUMsZh2OBnTuX
zDHDsHUVl7V0I09hWjg9lG8IeMHiSAiullSFzAJpuc7ln89kbC+TAFy4fkWswE+Z
/EZiGWZ09dK4qYxzswyhZWLSSM6BDK/THulJU/rvIgZ+46Lr2TQRsesk7lFtKfPl
ge3KpLbYnyRQVyZE4PxIqDrH5GMMZBcWkZPcILduz7OtMY5sHyywOrLYwayegOtG
H8cNQDrJp/eWu3+j7WpY7kFQZrZ+ZJM+PLmkB5ek5xSTBcUmWJ6W2NphIN1YegyQ
YasIPo4gM8alxAYBhqLpAfpuDBgfRvaYH0nKFdLNBjEgc9l8nRBB2r8E9j2kcqwb
zXS5YdApP6uk0PAswtuAcVDyntFHDgxYBX6kf5PF4vSVDQStSy0KMW9homqqDlhC
3n/u7ObJp8TJDcTwTwh40p1UwEOgeNf8LptZKOKDDu6vXvBG5psJtYKFfZdmZc3n
CL5T3HLtZz03LwikA1w4/elM/IRjF0Mer4J6m0XLJjFlr6e2X7ZoJyrBuFWl5dY4
VuLrN/GZUmMjlUMWeagYWSADYwzR5Of7Wm83AN0lcrWt4JLH3NBDC+5p9TDBMjKd
RA7SY4Zvzgfo8jMgnY7rNYmGMwEJ4YqESAQ+m5bxcecZlAL8xGidS+ly3SB3qUzB
NwBlY7/ZTZsUbST7yX3U6TbuKvdbzYkhX7IjVPZJ2A+ROlSqqjqXFkGVRiltVOMo
smIQDJHo9lV0raCGSaWk4qjg3NyY2Jzq7h3CinbEToEuLaZvcUOS5KYKWpfERxed
O2TEfQJYo2hciJy1TlO7/6U5jVFobYIqHQS/a0rmTYTFN3oPeLcJSVmMnqEj3dX6
40kRTaOcul5ISl7y0JgLZx+kD+4JII3ICGM5KOPZyFP0bx8C3Ggn9bvhNRdRP6u0
/3k1gxbqQTsoy47sN8tMtVOW7FGxmfW1SfSN7hctVdt42opRGq1yg8gnl4bURJVr
uCN1DBB/BiRflF81e+2IfRGqacLTjiC/bZsUTzovluY45p6TXzwhBAmywzj/kvk0
ZcWzTICAByERiZZ19Us7omZbIg7sxj6AP9eLgAH0D2zgQCwlFqcgeEj1ru1z6qoQ
8Is3u31A+ZYwMERqq8S4CQeMrBjohFFlv8kWybXuG9HpqlARS0aJWds0VOxUdfnE
z9oKumglQx7lzfspTAPb56dUBft5X6/u2/upbp9U2XrMbrbIdUnEPBgUSHLATrpK
Y6GnlFEh37pvqUl/FbzbjuapZuq8mXgoLswgCiWkdv079VXa3rsU+6yn7tHtS2ZY
q9hHLIcTUOauti7NXgHaA5Z844CXEug0FyUnbY135gvMXgWCquiXSb6l4cpzUxWn
ZKmMbW2zsDRZsOQ8r/lQn8s6O6cTrvLTva/szq2ZEFNGR7JeXSUQjVYv+S8bD5S1
iBK5I1YQ2ysePSdH+6KS3jCOE9tA0yStU5DK4ULuxSqEmw0ZVxNBNsLz9MvZbTgq
blC8pnxlZXZkyKUVSWVWniqZzE6uxxQIDrXVhMHSt2MOoLaFdGycaWvNTmMtP6+v
OEjjfk7GBpqKDXzmdtIu7ZsHZDDM90z9tgF+TcGfb+CJLTfkKSVV1sW6PPhxWO+3
NaQo3itorycnaqw9peZRnv4HufM7YOyKWld6VtE+LtLYH06YLOftVUrdDruUWQzw
ljN2YmKXVpzuUx+sDKtW54+Ndu3Qx/L8F5YUaoTDPCb/o+50SKN5D8QIvVaOhZfe
qdcKvxhWZy/Lb17ydyGlHtUM9U4IOWFdJxRRMszQd6F9A7risebx5VHUc4oF2zv9
r5/mjA00ClWO9KIeLZ96MMO+bkOu/ZDcTAQp+soRkhBt8Pfdefye0qiinS9d7uQv
i9xB21pnU33e4K/10nJ6LvX6WbpnlDZEB/5lC0IjVSRapYYRqKOyV+QrDVBlMI0x
fCD2REQuxyQbtxiq/a8Wr3gTAKpAd2F7ZtAkrkJFqCRFpgzGzoccUDKwhGvCqxK9
Bpctvub5X2iK/qulh+miqLLpRrh+n57ENaZl9RxuHVpXB3ZJ7fNYOSjzspz6i2eP
7M9aCYx5+jKMvyxUsACRIFn9twpOhwJ8AWjn2L0nj+fBzqn+K2UExny5o6phQTlL
PjjKunPCe5tyHluWCJlyc6ul09vLoZzhHXr8GPt9jOn/8PFhE+lw2qWdy/V36PFc
otqgtasosRtNdMCxo4tZQIik5cemjeRAg2WLY0HVvrh5w06EMZu/BQ0VmL99LLKz
kKX5LNyNSY2bi6ctnTOa9mKrJQ64ABRWLZpqfm9bl2D03te3S4e4R7lfeICNZzEd
6JhRd0hDiupQoFbCtB+RBIFCPM0MOhEt0gxvD+Tc9gNoeu4PZ3ETRb7cLp+zPiHi
6a8LTHggj//NsJ6nQua1EZ0e4WxKe8+WamOxPEkVX102gK2kUHICobOLtHsO78HU
jVEQUbvhfwerE32mOrYVtEaiBaP+KwaWoiLuikxdV7anrlQAcaAyQ6sJzmhYS1RQ
ojzmQTcaGnZSK4q6/6lWrWw4a4j8/DjzcP4frEmO4O2pR5SFiISOYEzOe4b+xcM7
YzQ+FNpN2xJfTHgg+oHLpuuS18s8e+oYjJCn5bHx/AEwXIVZSzOZoBTczDVPoDGA
DMt+t0erWxHuolcZ52wOqOBHGYL3DCcv2NLSvwfBLRZA1KuF4iSfSN7imWgaHXMJ
RcEBtR9Dl/TnK2Vg2nTs+B5O/k2Btfbhvbt5MNV/98FbhFmcfqt34KL5vpbVghn9
hDg+rS6kO89H8RrzvDdlnLOSIBVzUmB6gY27jQSKdBG70NlSm6xIFQcz2wxKPpj3
Wus1hjM9no3Ao0JG4Wyz+/YrN35ONqmCGkvHwvTyk8wlZAy3GCw0Vra/YqyFXF/5
+TSfZy7K05T7BGLIQvoto/GnjDqZrTXLw8e/CoBIH1CzCpz9R9vTYjnlt82+21NV
IxvCEwGDdGhAgkfMCBknvtftv+uSun/CPEJ5dqlYVzR7ZnJhzt+eiYEOv+eTBwnZ
7mQrYG1TjyqnvjXxg/cEhgV8WoQ7qVnRovLpbwZyBglieC/GrT2ru+X2b47Jn2S+
4MePj98mOM0Y1oZfjY4qkHy9YCJjgh1haY5B3+uHDVsOTHWu6EIGza7joONY1QWm
YhxKoNAwijab/tjD/Sgzmq3c/BLKxl3Eb+gYi2k2tukFiSSglNLxMjPhruouyszZ
VzqNqZvBm44JGpCL4+du7+FE/LY5UrqEBaTaMwKeCaWK4p5V3Df0Lsub70xQlD4/
ji4UvfVD5QHqd9qy9xKEWMAyqIqTArkzyOw1qUjSwC5asnEWWdjDfPnPlw710OPd
wwV8phDlezEd211lWGeaabgxXRTChzf6iUg63m7dlOpPBQPLAd6zcLzvSnyOyIrm
9UhgUyJ5KyERNdK5vVWq0cyLQ7nAR7lif1ctvEwAJgkU3CeOplZhRTN3j/v2Ivto
9BVt2mSZl0yVHJKqlhRsMTXDXYcq2lKhhcVMwwQwD9B1334t76TJ7pIxcweNEF5Z
FxhZIlfX3T+RQ1d0dBO1M77bJ/UcbMU6tW08BFWF8o01+IFvGE46EjkHjpir8R9B
BvsxjZo7fKrZ53izdj8hZFYTod0giz+cMHRAJel7fpdthds6uNL7GluFF7TFT/0N
cA5HPAkUwl3QkDsg+gWUo24Mrl48EhMn3dGlvAEie3vrgW2eAlL0rmMl+by//P40
2zIgDegOoex8Y5NEG0bYM7osuSAPkduz2NEc3PVPxo54KUFLGdHpv4LuLzIa9hDZ
m8i6cRbY8xpsvbVENkoXffr7IKfo65DD+UTmm/kOkJiseZ+1+8WPnp7ZrYIobIar
jxRbD5g7zO3IU0CEN7OsKgJXu2rPj5nHu3Zwynf0AuDN4k7zPX7r98PMoGkaDw1x
sMJa3vEasYlnK1YSXeg3xpfcYni+Xm1sSz/H9cQwCXnyW/gg02Pj6esHFN+vgH3S
acfLn4TVoKJRMoCpJHx2t7iNKp9ViueuZTeBiNaQ0/KcpYunFOwefwK45mDuXv+/
ROR3+stnG6dsTEZsioHwMmlM/NhDTQtquJv2u2J54Pj4mqFHp4cEF7I9D4DwCEpX
WCdQPf4Z6W4tmQx2cyxzkfa2alnI/bRuwL4vObt4FE1JsOgGM/9ppiTCp3z6NZ0G
nEvmzZrpeLMJhR3AIL61Mks1XOIjBpAB4jW2Wbn5IaAEtqmKkskQL7acTHUn9+tj
IcPlVM7/PX98Od3Z1vMpRS7R+hO4fOUSawNcRcxTTikQE6sxmUQnmPrchrnQiULt
4u7y/0mU+HBT2AxOKlkU67054rYsrHfizJPRIowTbXhGmR+zw7bn0azolOHzCxHU
TBBvwGxUty/3wDhSbznDYiEudFK14GyJbHP94MZZL3dkl8YOWmYuH59rQBAX4WmN
wZidmeqtFWx1iW/dhW0bSG8QdEhDvhv7X1zLlF1luTS0p9lOSRwHdKZj1fevPDaz
sMOgLQiChi/G8hywSF3ZgWOM7yFGbmKJruwcQKW9OEiFCWZQrUlTXk0kw8DAU78y
yv4lpWzK4e6rx+/SouS+p5S99467awiidkth4oa5V52esRtQo+kmcPhUF6MEM/SK
zJ5IJ95vIsppo3Q/F2ppG2YHDWuMjsGrXXW5sjSKDdCMGDvgMbB4cUCrB2ff+NP3
rZ6d0ruE82nCzGyTYU78FHqoL2Rt7QmFLrVArK8bvGeFEKRpPyyT/N3OLMMEKWQl
ntPf7xH7sMNt72aufesNfBJ5Al6UVLHVaOyKQHenB4jB2bS1BZD+831bpz1lQPDF
RuIX+c9KPs7CCJ11PGHxCNIxMm3UT0KbqhugJenZBLIqLltzIMtGhoH93gWMoDA7
vVskwSa88PxnGrraRpIrwjmLxX/k/47gSOUfPuZYnv6wZyTU2YW1YOhaX/JT0QVb
Ynw+QR+cwknbUeH5R4x21Z/qCj5kx3G1G6sANi5tcB18OT/vGf9bbWPIHCfytRbi
/uNDC0R7QAtMiWNS3h9ccsW+HXJf8ZwXTZWjwEr1JYJo536jQJCVh2CI1zttsziX
N52NSmFu9iUa2SCx4F4+JmlMb8A3PI4CZsE2aZM0ZAjxec5amJYfsFyEoIRo+SZI
5Gaz0GQOd5wks4NEAbEyuFQAwj+Pt69tV3y3BtIdk9JkTw/brk1QEtazPAEYJPQQ
tf+8o2Z3Tu5Y8UhZo1L8yjBO5r7P2bFS3bJpK17Kl7X7B+dDQb+nqly3E+MX6n8C
Vfr5Prxn4WxLr3kadfLcgn3b3zFrWAXCtQ76zn3TtQ2EOHBNETbSd0WalKs/iU4X
XXi3cvpds6eyJqsg7X1xVZF3urbnwk4UpCa94i0Ymt9ufCwkBE2YujIvSSy+C1gQ
EnvHf09EUJ3UtCv6j+/wmeLn2oNLgXnZnGxdIjTm0WKjrZ7d0haMx//K6A4WI1Kc
kvfrIiBd/iNC1GD1f0kHS/dLxhuKqyRcda0y2EuNIF5vRQBeZrsFkpQm12gqbHjG
jn5BXBXLXh9IvSmD4ydRosyDk9nVwFLVoWO5CsWO85JVquCtym0rv5JMGOEqmZN1
c6sjt6PBcOoRoGV1iLOXx/OsPCt5CmvLiLSScC48DCHx2qxevxyeToM/bkz4XVEq
5JJ+OX+h16/OlhF2fe7VOP3kJ6IU84wvnXLUn4ndZYukdT9Rm6L6C0M8jLEAz7nQ
y6JInQ0PzZCH9H8ClM7d9VqEfVzzkMiT3i4q+x+7KkAQ+yklq+h2B5hw22jsxD+/
lJx1ISqpAjgD6muu/jj54GfxVKNUqH8SvlV4h0zyx0zuGDfr/ONWdayHwD2/ShUB
8/gNn08uyRPvfjclScyKCFm2AtQzSObHXZ9ivO73sQA1hnvPAJR/UUQy7WatfXqw
2e6rvvXZG5cz36qCKKUoEjiOPQzm8fx1szwF7ZDOtQPbcJNi+j4ATIQSjQrd9fB8
S6YdwfNDBQwo2Rt5fI7K+6Pd3neOjJcGDDEgUpS4tPyurzAB192BAZ19q3Ovr/sW
hFsDvRo5zzS4tllqnPqNnOHuWJePrxmXjKCEzL82FWAE2jFOd9cQ0DePlZUjnm5G
jvHn78nkVMiVNFhlmpgd4PkSQtN6uqF1kqiyd2x83P4cUT76G+rRpS+vyn6GVTrb
fDh2I7zBiwHOx82iU04+/wUN3jDqND3Qb2Faf+9E+gFNeu6f0gwqKSt2xKTj0FaK
GKeE/JwCunZJ9PiVLBt7SArmOrL/P+IUlghDQxGBT+0T0OZNTgIo4TvPlrut1u84
Gpze0S4ME2rSEdJdqCjv7ZLBOueih4jORSAjV+V+OZLu/1TjItP/+fvX0Z6+4Mz/
YyTrBjEBHcsOfbv7KKrpcavf1cncNx4OP5wf9KJJ6POTACFu8CnID5CWysGQNt6R
y0L/sWxfGToaftcRWS+YeImguFEan7+d0HjV0bcqaqmFtQuXoFtJfmz0XHXqt/vC
HSF1taGddh6xkNHHvcA/U9E4z2gIQRx/u2ZquaqGrPSpJ/DbBhjO0VEEKjLot0pl
y75HhT3gUCScm7/gytT2n5k3itTVt/iJThloc0NdQTiECLB79QNkNoJwJ39rIa+K
VTsRw4HseBMW9n+8pSN5A2L8r1E4wxP9/wufRGpwa3qLoKTf9BCu1TXk4SMw/m7n
8W1Qr6YRy3ctDNkGLnGV06EaSH96AcoC0hZv9yeRlfBc6Da2ZlTE2T2mOxwYnRYY
kBjVDAmWdm0NqUiFGbNAsWQQFCIKNFb3lNcaVpGmQnBWNj+8eXtZo/Ihv7mNhK5Q
Jf3gN3IjYoKzbdvOUJn0vf2zsKfpdu4IUNQrHuOSqXQX/zhLkRdbRxrT+FWakq0S
Jn3YwmF3ZVO6/gOprResuk4frDSPBbQZEu//z7zndKh/vR5OKLvpMszKFaDmqf+i
5HiV+Y5wFXgJLTs6fIJWYpjCSpVEBzP8jzgEGxw/boCo4S0ozp+SFP7rJs8NoqYq
+uupzp2yXu1LmLPy8wJ0JVMqiU4uufoWxj4xcRo4nVeoQnLYXlBTmyMZEqsRBprX
jOY6kE5RbmGd+x2ruDqgJy1urO5WReINAVvNa8rr04oV3cbXjYjVv/oeFTQsvVAE
cZb6+TJpbptEEiHM5bMt++lx5KkK9VpNPwuJ69cvikc9y+wlxXNp50e5pOATy1vn
HvCvi3tJOQFIuJkNtNDQJRbOD509ToI/+vd5pYzHjRqRGp/blSKmlRkPBsm3oy7I
ZuSXUgHpXYlIt2lZF5HFdiy9taq1cnZqAE/Xvgr2CR65xAVWGOI2mS5u7RMHwwiL
ZwStvfArjJkCwTgES2lcwGiF0dM4J7o9HokSFEHIg2Cy71YT6n/xU/hJgsKb95F7
I6kI4fdHuN/uGzDN+0RR/n10KKb4kYEFIhOAJWlht2N5W2qzr/YztqxpNZ0WXO7N
JmyRC30lK6dTgkkY4Imv+dTSRYfAUHUK4W9T+MzSC/TbRXpm7qJ/5Zi6cKHRtLo1
U2j4XHwP2cUJmC+AQH6ctphmHccb5CTlcmj4kjHBO1kj3Coj5y5EdoTPVmR6bqlq
SGvU3SUy76nbzYYml4I20d+Cs/RN/rnQGzFahHDOgtPeqLJl7cuWXyVwKrHQKPmZ
FyPB47KBxyDTrW3ltE98xg8IT4l4iXtGgwKzKgIkVu8zjDvUv5aerEJkGCnoHd3u
Xaosu0HyCAD2RsGL9OmEPEYZsDj9BDdQkPFyIMkx6uvAjdbwi5x7Pzg2RR0Y/9C1
vRWuxj7oXQHZzM5x/Ntx3tSvcyBYhAUd8GAkgPFwB8mEmHyhT5mfwwYnngz6ac3I
IQZFKPe+/HCyA2qARPIqhBOccuJWMmiagGFIkZmjCJ55FLY0uYmJIGXycBugVG64
KEl2mbn6R8VrTxgzj/g0JedvWrsF6oOkPsL9iFig4xPRcqqZHzrzfOrT7KpZrTfl
Zbc2HahDKSoGJkvGa/xQG7Mec61jHTCjPaXrHZS+jSVT4snNyyk2Vwc/AT1G77J/
wxwHq7Jxy6FuVj1TPb3U6/P24OmxgWJWiwvJcMR+UQq31i5zjj/mJHnYICFwdKU/
bHY5V7Z2yTW6sAe+/9qupswi+F7hPZP9NDLje6jCTe5bPJsKnThEjPsi7Qp4bLhF
NOSV/x+TqWDHbcQpTm6uHiPwOdN5Wha5B0LlzoBI9bgIfWjaUaCB82YHYC86LRoO
WsUnD3wVAXIkOWk2lNW8fIIDpXUvOFj/gZzqNVck350ZhZ/OobA57Kt1R401tpyk
Sf+IVcr0gEf9zXp3Q9nPVvP5Y/4suuGkTpeJjT80DQEzycwMFxQXwASEsfCWyulD
y71l2BXe644t1PiCrFrCR8ZmdMyJCePdtSNStrL6rCuNfdgQFk0WXZ2UtVlzFIoP
TzEbBI12ST8fYELvbi7E7YtumuYyonXFq7Qot7QCVjeGsX+SwBnuWmaJp2lCtNmS
QOTMNZMXrzfsPDuji56dsdvYueuB4kI9qAKMCFio3JnhjlOOiDA3v2sJggASC4rw
066mIDjIrc9/SYeIfRKg0dY1Dvj/waL7qvyp8hwYPxI0+lH4POzPWe/Ixda/31YB
/khXlbLbH0tT+ORBkAEYyUFq9eKZJWBblobg8h0rlJVXt4+ilS4xpYwhk3OcnoTm
T7mGTnSTKgLdWVfBXlpGbfZLjvCiI83RsSEWuHZ6tOX83E+q/D0ROEMM7G/LUXBj
Ms5rT9zvdYZVdhJBem0S1svCdiScbHXvHq23yVdP6XzytT0n3W2JscwG/mK2365b
eMm9eaYbXpaW4f9sZg5VJKwQJC6pmfb73TJmsBCL5eubCPSFUnRXfEQ1URix0+AR
OnhcXBW+8XfHZdOtMK2rchjh79WJC/xt/afOAPs4EXozB0bjqtVKMcybYuH9DQ1t
dAqwsJu1qIox8ocw4x4CcX9h6FXUpnmgLrnPcC8U6tXZZWDIzVUN/OZ+RT5eapTQ
SfqDPFKA+0VtswWg0aJvArWCz0qduP2KXSL6p1oKn1s5xlPHhLo4qCo/JwwmkZCA
Jy/30yKGNTJHk/1mNFSQ1rZrzWuWmAniXrldV/I4VbzuPc0YIMccRYslAN27EpF3
ZdBQQ9kZthEdD2sCVFSyD8Xv/3oaeud1ki4CI1TVrmTm6zNF0ER3MX76H2hIIP4x
OaGpjpY92P5H/+ynzr6J4io9CNOg5gA+4bPsJ3Mr2ihQ9FSnU66wFCJg74e+JUW4
ovMLxV6quJoFMLNAY3s1maYQ1zLqQbgVhN11OkE7VwBPf2vtEFzak9chaQxzUV9C
H5DCw+IkqfhcnYVJ8HfmE55+eU5Vh1sXQZbHjqRfW02T1btEZkyquBbhL6byA0GG
OEfydqyLOOtA7J4bi2bygRMUAr44EhEDUM1UYu7BzogbiSGAmTYGfwTH6SMkL0bg
sorK9355Oz+ThN1obVKninuzaI4HnAQGJg0A0LeZKTkSl9fOL40jIstcywX+0ixw
HGXFyFO2GgnuPPb7LhnNLrpH3ZwaoxP/dQY4BcHL09+8z6f9SxXTIrPoVSSGFvUP
dOWZHVbND8H9EboYFdIYn3uEou+Rlg5wb9rDNTuWj7FixfQudET0G1wG0FTE2lnY
z98jOeVDh0tGZyYlmklJmFvXgjCS/B8vhpSZ9aUFLUlMQOMH2WTpRzjgrI0lzKYq
wHa8BxDu29ra3TPEsnAhm+hGjo3WPI2uNmAYmObA9/p6m1pkwHvewl9CHoxBNhhD
WHo1dfQtlJCvoQuw0qfNWvftGq3seWMZGqAb5hM1UqfUe5FVuFE2NdU8qXILC4t+
xlgjQnBJy2T6WuCnqftrL5/LntvH+IgeVISy2CZhoH8N7dmUpyKM+mVoiys0dPxs
5VNmrICKoUwWuZvyqOnNx+Kq0KOtIj0yKEuqaeLAhLkJ7bTfUWD112Qu1yn8jTX0
71utlLouaQ+lK8vW3bNv3+QbXXKUimWDub+M+SfXCFfQAWR+88qUJWUv+sZCQAaH
v8fAv2ps98IvnMpifHQgfABUJFUfjRySHunQqxqJPN2ShOfjfouszb2/LQ5Ljox0
FiOUY+JZghbkh+eFGzuRzpPYE8n61orCfpmpYzAWyEFigEp3GVboQLtJpew2oHwU
3Qw/e7MzC2mpbOnpQUoWeLhNJL4FNY3BY9VJ8DOtiDEbZ2cG+EcJa/ZD5wdPIqb+
AJk8rxdb0AJM+XdPIx+9OxcXjUaPnaOkseHseUWqFnt/PToRbhPKg+jZ3upMdXnW
kAL8t2K4ZIHxexKdi8w44FVYrnoZnrQIjKpCr4yGWSR4x3u0G7D05PSuimu2Kpqn
62HWBg+vSDXHvVWbRUTygXWQKNONZ1ME/8nLsg/pubbSUcYurTh8WjHPO5R0RwvN
fIkowUrjsVxwBkezieXXfGPnNIh/FoSxuVvg9xdmZcZarudAf80MnLH+JHoK6fqH
0Hlv5XeNm7wK2/QqF+JicOkLAX3rRxrUe6UGsRvC/FCB+CvU9nR3yqmTSg8UDsro
GKu4ONIBGrx0yTwBeJJARoZC4AN+K7XT2vod0nSiiiS9FHfU/yz63rlNLlTIhxsx
EkakaLLmCCwmZ7ebXWbYTnPt9FmFX6bGg7ejTX/OTlVvmdW23Tomn9uY6Ai6phE9
9+uAAeaMltkr2WEZZL1B+wmV+U+ATRfXYLPNhs1IIwYynvKavLfMO/6fVPIC7Ifx
RHTE4i+oJOPwERxiyXURQxv6aWjS/w+szj/kMYAPyy8JY656LDiDmBApsto1wRId
+zkWxU/HKshMXDqgQTYFbOOKcgdbnRoPpw8s5Qo69UZ3yTi8X4SUgu6tSp51NRs6
rGZ3eVvESrpEY6J+wkqm0jzbO7RHR6q9OjywmJ/1w7t2spyKo4d4ShkrHIgkxKvA
Fd+L/rUzo0Iisy4q95mJdXMjpaqdRMcYyK6ot+F2Zj24zvfjZqHqOr2TcscbtWSZ
rgyRsOfrYgq+spSsacqynox3BQmq0W7YD9ie1PfoZ42lQndbiWte6L9HI4ODEyOM
zHcxEgQaks79hs8Kh+UYFsZuMh7nnP74CH65P11mX38bVR3PgVCcN6jBxUnmuMuC
BKiyXRpo0G/BmfzFlGhPLarWZkpknL8T9hkZxZ7xAyVBU5hvR9icOppUzUWi255u
xB/02svCITMM+zIUGkWF4GFx3c+1WHvFWMaxEeZaxDc89NaUYT7HCyn2tROadUjZ
UDo8h/eOO+2o4psDLCcplrAgD8qFxNgUCql+NlMEs2OnAIalniwAPzL7GInwE39C
BDMExUJPj04FfiE4ysrYvhHLWUhTINAS2Kd8f9f8S5oIxaUbI6cKxbkCoqnStAyc
C1xV0e9liDhKzm8nZ6Al+w7Eh4EsC8i5TwdChx1vg509IbJYROdhakCFrTDly9mH
xuQy9tJuw6E3utFcpvvnJgDe7VOxT3yyTnHoHwfT1z2oZNaRjX9DNAmMXyXB+rI/
EyHYhzaim2hvxkdyGfRJlu+PqO1bMcH95aUxbVBx641JW3d9EwMF2ZqRORu2tWBO
OLtas+DHJxbuPP9kezU/FnKtwQ664oF+uAE3HQ5Of189LkIH6iNUsMakjM0d0v/G
5bNSy/RI+g1T8QjgYc8A2Wk81KiCrA+PM43Ls9PMPMqc+la2HqmNAcmYtneWx8o+
ZfXvzjzCV52gL7eqhIJBHt/ASafZz9xG/9nKxaOD0iOyCBj9FnNDM+80dEJBg7yd
rjppJrv5nlUV6mtvEAZA87qD+ktIhrWcsVpcaUitmIGRjxGTN9rGecEGx+bVZQkl
lhs9fI1Tybe3LJqsBgqH/MuOSrmHjHrWD/EN++IrZFrY/ZFKs8AIsIls0/znFoBu
TU2xeP/456aald8fSdT9qh5hsD78C0pJ6ukinSGWcbSukpJv3Sq41GfIryyoDuaR
3RiUT2MRgAgKCIJsdGF/KMXeXF2b7h6ko/MT+nZJ9TRu0AED1oIqfdGZlReXC9AE
Os3KWDJ3dg9buyeCfBEeywMMH8sczgf4TRVo4JsXUtAe9Fy71kW4YXqUteFq+Y/H
/llZXbX+JEVPWw9Nf01X/ImxUIVntmiOvwn3MrC1J+0y2ITnrmpKEJy708e03d1O
ZQle7nY4Y7tS0wAf4xHQsvasRcNA7efM+n/q6Re4bsqlzRzwn8fN2Yn5cx7V2BrY
CRF9Y2DKHgQ4NR3lWqamAvCUidhg2E7oNH6NzwkCcqiyvP/JbbbdMgO/FiSW9DUx
u5bgedTXuyu9mWMauxfgPUIeDyLTQzHq8/lPV6otaw6v6UztFOql84qGS+7lqdfI
NR1xqr2O6jNDGR94JlDD6bFf4NgD+8P4ogC2fV9DAARzrXlxAbwGMtP9FsL4UZpz
glm6X30rwzLr4k/JA9IXteGetOtPUnlUNo0vN9ZIofEANSgi1h3/n52VGiwo0FOX
ua8DFiaECrdxRC+nRgsF9bSawFmHcoUT2nklGTOIm9ivfzfE7FaDDUjudDFE24lB
EhZriBE94DBqmgdXkaO6Zh57U0xXEIXxQkkOcWHNzYrrhjNWqDOhjr4cLvVVIozH
l+1oapzOQuK9lopMq2Rat8hvVCuOeRr5cG+uAacTpgRb91m1zXvp4u28V/+M7cVn
7i6UPMfL1txHXyxh5PzrelGgmnaw4c7dvfj1VW3eBKqQtY4kE2KKN71qZtLZX8Am
C+BzrSLKbHUQHS6H4bc7KAbiSXLIBz0yLJrF13KSW7M7smrgrNUdAH2LcZDzAUE1
8aTLKaiL9xzj2AbC3z0HWZ2AZKph3xwsCtVqE3iD/f4W7oBJ+SeSUGdeMxni+2hQ
1azcAkV2GuRyMmaNQ+KIDh0Bak6ubowc1G0MBTOi63/csT9r8MpjURe6tID/Ielm
WtoGbcE3ITnNNeHXmp5ps5RYIazxxbna/0AsDmdwvfbVv3KtaECFKxTwtmLi20qn
4EXmDhKg19o5n16hd6BfAU6uF30aPZeE5/UJziW9uq4AFqrBlOzSImTdXD3UtNJW
sIRSlbzQ4+fAeF0mr/9n98+BJG/8l6uG16UItpyo4KeXLLDvbwtZFafiNBoSrrHS
bHWHbR+6rn2kD8zZlITP3JvnVNbvOaVfVw/voqF9lL7DEFMu05JXvF0iuT3uvb13
36Kzqbu5nE/W9/BsaURuINLQmnJJhcykaXT/5e8SLw95C5Ouxj8u/xaizL4NYg7N
vMvyxb1jmXlcR00WT3YfuvFRaTEDPxamSBUwd13nXtusQqHkFuq5v6aSfTN0ihXy
HzxSrTjwhJxiEocf/Tkl+yqCB+goGnBpTGeero73w2ywgOUflSffE2FTHQC1wfqB
1i+xp3g8jplzV4m7UjB0n5yG0Kf1JF0D8XfnYINFmL6y4HeUGcuWl+JsbABIkJJT
rss3Vda0D5c4hk7M0hkbBSV4594HoKSCygJ9Ey+HaIvK70cSbgDlzZCDq6xE7qCd
lYRruUXka/piiRQKr6JOGRg/d8HE3Nrq1zVOVnQO0YWrfdosARllhLL2n7JeAVnf
s6Z1cMvPzAZ47RUeskxk4W/t9SXxCnWYAnVf3hOJk3XD74i+s2XM5hF8tBH/DvA2
Pnwa2ki/Efby3SI48eUbZLgZ2rNQavYeoJ9D9IMnVQCAixjRWLQCSWjSI02H1YFE
xIIreHhhfkf+uK5r7ni9wAqH6qaHtZTJMK0qeKgwXsPRsA+4E7NR0bdNxE05fq3B
qDFH+ZG5v+0zkBm7nOFVJ05Oc4jkGImHuTk0DA/52IaHeY7oipTAO2s9g80TCNWv
DubxN+bYJ++3SxlGmbLFX4Ih4cK7iYPp+8pUfvFABm+tO4T6XeUEkSPvTt9nJqcJ
pHLS9+hZlFBNEF7KvZseq9mHSpmQwXJ4vKAU5s/iV5tq2Bpybm1qxnlUva/5L/WO
PObLEvc6h6MW/7hE4uPkN4klbUEMtbNPh3Ix18boy3mA2yyZndd4zYVaqgrCHcIP
Mc80qK/mGQVNx+U/p+k9xHF3jbzpQW6F/XIT6Ro4UDP3tf+hl6iB+JPXCGWUKkjV
2l90AeXQdnLB43iFyqnlmEqVLkNQk9hXLcw4YZ/JtbDFD7QPBHQZ7rzlN6wYlar5
jhOc+pMAhei7dpqIORj6svRPgDP9pSHwJCTsuM5Mpmh3UYBaG2Ob0PKrQlrT2Cf+
5T5fH5Q6ucZBXsvBHMvZwuMKRYcb66VgSpu396Evq034jYF1LJSO1aheOfSdYSaW
d6M1WqM3tMeGC9lYwJ8zEn2XdEcDYTwqFE7djn8ilhKSw+N0XeCv7czoFRZHZGZT
1Nrm+PdcTfRgrhSSQxI5nxfuTRJuUlcmkj4a5PhJhr/FGPEss3EpPFfhB4OhaMzb
/fDP13wr4Ot2q+yBS5qFKQGQJsBRuC4Y3kOh9dmnc2OpL6ZSYqIE6miykpLbuXsK
HE3LTu6n1bMiuypYvYzBV2Hx/4X6ES5xt8feOnZr5Vbp1AqPubBiomHqV96SBLdw
JalJfuS+MJEuYD2ZNr3/oOQkDUISr8mDWTT6J4StrcRI6HiY5LJ7C5gu4M6lHh3X
BVjh1YmGZV6OfYwOkAGIHov3EhkdEe4ANvRJJxc+lEHuJ/qxyeh1eUOMO5PLmkJi
z0sNomKwy6qNepVResZOuETSIIY1zsC3QAVyjU74FEB8Yls+xLQUGU82SwcUXRiS
wxF0AQBiAuEsK0vMRk90J8xxqQSMeJTTgVkl33vYd3DIlIvZLp7q02k/dZHXyf0b
HFLd6CuTLCbORKfKoHGyPVuzqTjMdjJpy8B0RO/EmDXPOX2Jgvy7kz8gAdtgTBsW
t0MDEuGI2/1XYmvVuQ8a4iWO4O7JgaW8KxGZGmA9rB+cWlAH8hVkpD2xt9Kkt6MM
i8/AtcuI6ony/9CStteuhsdFykw0iiCcR04BXunA/cvd+Fj137aZYJR9XOOnHIAj
2I4kH1dqsyVsSztg16NsGLRsy/n3STn2VN441dhca52k/fgx6McbZ0URieTc9gTR
JNBFgBlFaW4Wi/DcH+x1ZbOsrDl1S+f3A7gUknL2s9spE9WJ3j2MPyT2W5sWs+B4
kkPPvBCQ8TfCJOTcL+9fJePRxTipCbAI6TLPiWBU5VPlXlt7JUByEZ+Lh4P2BvjM
XCQpICojkVUGeUgc09NLmkMR6HaDJzW+q81nzKby6qK2WCTjoMlTY7YSmaCUuPWj
990v/V2n+D5PplMhZYpaq5Lz1AEyYZeBRtIBldzLhWNUzacEOYvgVP/4i3ewCByG
klDouqF5wY1vkL02x/75tjPGD4TRfVTX64PGoUWvYBg8mA5X6LHG6QkCwG0sOpvJ
lvLDvi6kRbKpDcCken+m9cIFmOm9/xsmlFLIIxTUhj6kN6bFmUqVBycACd2YvmTx
+hM6h1SQ+n+PN0vv9oUgIQx/iFdbN55Wu6gyPZDo6n8M0nrpKf3uVFPjubNxAlD5
DGmiBTTP8z1EWm8p3gIwnqqEN/fbYkSxuJ8sglAl768D1lfgclKOhl7KCrkDnfJH
CRS24Pn4N0le83iy+WRs7GUWqme7FjHTRn0fdGVxFBzspOYiSorH1s7BYBLTlzLs
CsRnnNPTL61i9dkZ93pTXyQEONSddLUn6rSy6FT8KiOfN172wbe8e637XGJxTp7B
U0atXUpC9V48lEn4Tmmj7MaxvPoaOv7gNstsx1RNYZcQlEJtwiKxHoi1eeWBVCdX
yMI/ssOp5YFE7RjIfGHTaaJu9h8O0QD/+WpMPctWr4BQ2BE/FU8gHoJfdOi0QxUe
mcyTXcbMN72YcEznHdJqh9eaqgAZ3ML2p71y5HWonFCZ20H4QE7+aKblvoLxVDM8
rG03BwBn3Gma2eSIYf324X756lOYINpVBYS7gto9ZyphTo2QXdW9u6wctEiDf54E
txO0g0bfQInLCTSHeTfKAHYRfhHKDGt1+kQyD1YMx4HqO44QUEpxNyj8nEX9ERLP
ORq7b4EUcBYuBaXaua9VZ88kdT5AEkRJfrMGzhJvrTygmpCreO45Z512d8yzvUsy
CVj5u0sR7nvm9+BNYuhjzT5ABRxAFGUH+qoSSgx40qy/xyUIgZImJGxJGA7mVh3A
nA0N7tfPrqbO/PcVIa2JyAMFCwovzZsVygqwnrdrpQpIsRaVdDb/yz8jaZiUkK3F
Y8aOZetCKoSNmP0Qow5VKzsaF5uQhRjvGVT87f4wHSeBD0x9nNLABh9bTD2RHrcx
jORmlvh1DzOl5yNTcyDo7CFy3XHKkeSsQ4CgalQ2y/5lFKi95J1QJinzrT5c1xUL
M6N9mwP3jAdfuko/3BNouKtiXO/CCfEsmQQ61uMLrtQgiFi91d4ebw5L0jvMNh1X
Hd7Frwz/Ztd2gtRnq2dFVnhBoSJ5z7Av9aPaOPOd4PBvFzQeCuRMaUJh9hnvZrg4
rS8fpUPGMzfs+SbOhGsVFzZCYJ76x2ehi6rIb9xtcYgytXAwqEYDGE/aXU/uXpiG
J5k+w36pCgg5JZt8LsBCPzu6dGWHd3xduPBStw18V3AKtUx2y5PQW5VjdVXd/Dvi
rTTK49OMPWg6oqOfzHl3rX7qG8eZlO/698xzlfGH1C13F/bIrdqYe4XREHCIuzBM
uxkZ4AolNjnOyg23XIdYmovfSIpH23dwn98oYztl9uyDcIvbE/WQCd+S8NJR49uF
KfkTkM+7m5/572G0r2Vn4jgr/vWSMY6u69sazQ+pbMpG8tFBXI0bk/Cvbgm8xHVR
DSwQsnM/pRaCFRaKO2HlOXsMqL3d48rFoGY9SOWvc8LV6IaRnKis08sNPkPt/da5
nfGj5b5R/JSJTY7KmMMOWTHY17bV1YkibftETASXXJLIaCM8ZhunEdGXDcA5MEF6
9l7EtMnaRr1PFQuPUFzWkE9nc2w8S1NEVlmRv79QzaJrZBbFY54RmaMtppyCbxZ/
xQPNcCU6dfCp16ZW3CElK5Hd+4hMKo4Pwpjx2HLEZk41mzMepgk+BH8rtnkD26er
dH5NKjbpTj9JgKq8Aj1pSMTaM+pGCvPdGdgRjzkA5llkZTA2mEii+WdkRbqQ+tvr
AaQEz/nagoG8RkTv0hGU1DVQ01jupr080qB55XnF9zCB+9fcy5OnmVopNwvgg9XX
DWSovojDchHsOLxsAB8M2ZuBWmq/a/gSaXZ9SkvuhLASXjwOcRRjkWoI7GMIO1sI
rU68qbZX+x7TUFpgO8t2tdWiIVFfB8oPoea8DvK6RXRh/kP88Q3x2z2BePOv8CTm
0+dx8+OUyY8n4AVGIsqrD3unr40x3a08MztgkI0i5UrLxuKG+FTVAU+1aknDyCDd
SuO9F3IOectfn8UX+MjlsUukH5ifKuXZgLzxoRRxTpVniZ5cFzNUC+B28f1n8rKO
xvRb1MvJRyRF/S7w29e8buM1EcLeHzcOn8DgQsQqNAxzmJAtjanqY8UGS2ft82eq
X45y9JKc9/30xcM1tW0jfObouiPsCujc6owkYLuObq5WrvzySCW8B6+dLnzDfogk
hgzI8Z7Y6Uj4GC+gmenOO82+tn7NO7+ewcMVF4i2oPGpsQidWEFxcWP937rMc4cT
7dqyDy14GU/0MF328s8+eWtOzAXtr/wWU5LfRdcRSsFix2jOiwElWh31UNzXM++S
ZpiU0yW6tE58fkhYMAoBDwQxMF+ApDMW4TcahHlKJBDsdNS0IEp+e+bXjs84Gvq2
1JJPfJXZQnf5lLC+pghdOhs88j73ZXm+ig8SK/KYa+viQ1NAPuevyBP2EW5+B6aX
9LLZoc4wkXVXAHEI/2ccybYwrYKccvBR8NtQkuwfFbA2Pt3FlWHidT2jl0QcCJRS
8jrpHPaSRSx1Y6YjS/Gnxo/HT0oXXak2Q8Z4dR0C+c/FpajlWdUyJiqwJrkozwqi
HkeuItYGPflGnKJ6kIUttwie+uxDCLarBNT1peLk1KmI9u4Y3qlC/f2t6kY6gmxf
/BrY2QZ70A3SQHa2hDjuuDK/0jJNTlOJG/6Q7wUyrQxdRPyuz6dkRneyWxS6Ymce
O+sWvx4icG0WVuAPorExSsiEQVi6dgods0fHwLv26Jj/5prCafN7oDB9RO3mO3gh
7SDNDjPKL+yLE8MXoEGKg2ZuLZmla9+0kEQ9lS+52tvJKe8Ax+ASjGt8Ot3uMBEZ
dLDtTDgJYqmVnP9mJ7LeQw2HCySYjtgqly5JkXERutXGFmPiXQPU0Kcd6BaTLMo8
l6j3D+m/Dl1NHXs3XeSjvB9KQITMPiKpciOkFllJ2iNrRFEIaGJtLj8JpL1UtFMF
lmvnM0Hb60vVClJhC5T/2DVSpYE1AeuTMY77NAP4HKrvzplhFOigM2FsnbTGRhmR
VN5Bi40OOWUkeZZTrxT2wDt3+k60phU4bESefVgWdoNDzVtOD09RdcjcaLcPrdPR
QbshAmh0+Yg7wrAC+DQh6Bsn/lAd5FbTF+uffNJVtJTpzS4qCbLE5pgj1TKo9YwV
9xXSmY9FblNV39rQpsIO1YhqSqaHcbufxNsWV2kJYpOhoSmaNMFDklC4R4TYPx8E
ABWFCSAuElGOJUnGlTKC8Q2Efd7Oh0wGTp87yb/PrrSrloCpD0IicS38V2e70+Vi
lTlFIByCEn2AivG14VDMqV4+dVb1MHLsfrymYGT+n9GvbU3CAPkd3IaJAp6+RTVi
biMg5ijQlr+JBvuQ+0/2L8bhDHtXCGLkpYQ7PMFDC3E0Up2Ygpoze4X6BvEXh5+d
e9URMYsPxjwGi8LWIUPFdMrCNzIMkA99sSXqR1XQBm/FVsiivmcPXAkdydd1qFYU
Kho5yqg8wbLJE64pXTBESTaEMuLm3LO/OtqPnrhH2A7RkAiymlDgph2o0Km2kqUj
rhi+zlT2ltkgSsH65Y7XhYVfTBg7oT3Gqf1WjsPAQggE2xogBvaDBFmm2nnolJ5O
b/p6NTFKTi67cNYiFvV7ix/YnGutgHL+fSRgLanH0mRPaz+7FHhkQMf7zIKUPwAM
6LsB/X4FfceFq9MhtcR40j//hz+NU+Ltaj4+jT2JC86nPYDUDsgfL9Z+efMhk3WX
kHm+Ak14Wc38q73r+mgqyHCyl2I6EdbqNiWpLVewHzUByuxGyrNLPw6ASlOb5lah
ST0fwFbUP9yNmVRreOy4ar8+iQmCFO1tIlT1yj4alBQ7Ofoao4l4UdfwO7TFrjk/
YN1po8YbvY1GGqErsgbwPfac7fVsoVCunbY9PgywFr4I/HOSIjDImx09IyzIrO6W
zOsY6xxQjGZq1gwaMebWnLx5BuSVtpvNe6/fXAfHNDtP9EKWlYzQfx44C1cOGpB2
kHTUxQmziRgUl+aSn6BKBAmEkP5yvDc4FWcwflb3ZCYxO5IJJZ3PMzZmEsGwdgNF
i1122pjFoazldRWSmU6oRUqI3CMkRCMFApjYkooDUESoGTryrghcqpRCsISUSoBU
eoDW6ArfB+RVTfRuEirhxs0oFsZgGai9ugdKikEbFSHy+SXDVtrdM0E/vFS3yUUv
BQEKmRFpB4HiyLnwPFZw2lLTXFoGoQj6ND+rAKycLp1kMxroXMOPKmaAL9O05djn
i9dFx/Nsz/jjVIRQoRD5W/XRvZtUJGteb52qKBHBQ9qI7ieIpJA7Bb2TINIGEx6L
18dD32k3pa46IP6as1+YFqvBcdyJzPWoilQVqnSYph3zg/wT0Ho0TnlQPh9r0czE
T9BrRU41y9na4M2SmM+w/43ibh7OwpAD2BttC1m9dFcr7xy/ZZMiJzmb/N29RlQi
Z2jbnXUlg9JqGaKrk3wyH6ViUpAncbgLQsD2LYQoxZlfn/8/yMKO6BI7edB+ifNm
t8MSLGC+ZiN1vPevC1GwQK2Nc8Xis1c9RJegZgivvGKK9BkJk5Bf6vcE4n8Xb/Xb
ebxa+9rX4kIREqAibQxe4mrs7an6EyMauOgR9hHQAqU1qS5+3CAtEcvfcQIIWNa3
UfgsRVDzMqC04vWIq28GvZ/YKfv12aZHQhsUQvM+Kh1NXoZrS+P2EzneyYzffuyU
+tGQj7j45XaooPtn8EwDUNg1yckNYgb4LlCzFKE2yDRK8dbKDm0PUpI2iKRQyF5T
FPKbn64HrZpdGl6DhZtxqXPbEMzKK0i7x+yKoX1Zw4wDJBbbwGsUaGF6v7AEaZ/A
ui4glNd7iOgAy408RmZuVcsFxX6djyksp2G3puLKdId+zUxKMe5Ixl9o7vb56ajH
K0TqIcRcADwnUrdo5gxbOPo9HBbl8MtmiQWKJlz6ZCBR0ml8epjrmJmfBcpBoj7A
Nfpj29LF5p72oPYNDMEhy8PrAbjl2Z9VWQFCjnKzeNgDTJb02+eE835FIMu+7R0Y
IxI76rraxqmlA+kfmlopdaNCqh7sNUuKHhxkpOvewe8fGJS6nkXCrML4S8ztnA+7
QHmj62xvHzeLfGLTIlhMCIOSNSYT/WYk9eMoGw5SGgXLGZGwNzXIwVzv9mEH4zth
pqX5wuXf10IUKg9xg9RS/HiPkvWkLPWie64yVLPPF8eyJttLAm0q0LEeL4NyLKzG
t9wi3poGBFsLEkBBjOKBwqHTW8dJ44/X8PMABeTq1ORyia51Yxbvs2G8yRDVcsy9
OPTi3f5Ondx+183i9d4II05A+GH2rXFhLfPP6uOw6eauYfZd0XmkEhEh1h62JTSa
6k62bTJ/eCO1ANHRlA8ZgpVWR8U2G3ROUBv7LRN7cAZpOrnBOey2KJT41LxycKn5
LbZVn1aJzv8P96YP02IFpL9DBOoTFgeYLh5GkNtDp8G/eUeovfJ/3YWnvg7lc2ia
ZmNeAhOq5jd4U+hKa/VhiZ7Fn0nv06gUCY0p9U64xeyxHnEqEhuE42lJ3dKELlED
GvNJ0d+lWfQN7fKJrbiGlz8OTF0VeCLUU3niPj4nXgYQLdgD1VHpFX8vJLKddnfM
p3gg7V9FAX/SydaOE/CsiIl1KrMt61CY1QRAzpketwtl4G0ix7LBUZykhyul2nOV
c6rsUw+cyLYGRsY9R+5rFnZhXV+czkF+O/up59zA9/xwHl3KhfKkKe+9c8bt9ct2
chQT7C/3pO+r5sdp9NDZtFkNbJv71MK60gHdIobQ/X+wD7XPadANTmbLA32kux56
CbQg6nWd99SXu9mzeW7kfUrqJ5TAfSCu+iebJmbemcgyFpzWjrAuBccNgSofpNCj
15RS01BijzvYBUbJOU3c51H9aKiA1M0Oa1a7TSgy9njKOmsLfHq/JNL1jrf97mE1
A3x5eNHRdVkrP8nAbrSjaxz+iMehqX+kevZ2TUoOueWoKC9WFeywBEbLrNWSFY1K
AYpu7Y6dw6t2iwlOEyEoAKUTzx7pKGCkxAvnhW/KnVI2VuclagesXI4ek/P/aoK6
miOgCXVXu4t7pGG7F0im6931EXR43tcgN9HT8lTB8Yywc5lxgowU0w3lDfIKJBac
towIenbl2t7Lc8LtqL7HLeOGef9neDz35U07cEXTZdwMaIYjmGzitMBUyAmGsaZB
A08qpLVTYIeugs/kGjw09BuS/xtxh0BUThDrjpBKDiLJORqHgKnnxR5UxbhaPaLJ
l/ZLFFjDTxJkSm5Vcll6zsPvV0wmep27aTw2WoRcTj73jZ1+LDwqP/NpAyVOI6wE
ClyUNmHNvPT+FLQM482J7DprQBeu7jfjb1rFMjRcp0nn41Hfg6yCo8VA66mvrPML
GQnaEAwqL9pt620c/2Qa7GlV+sABfk7aqFIEKh/9K8wyYDs2lCy9pQ9Pik6UYgtC
xQqCUplEw9vYpYZ6Wuh764tcn42A5kzceIPU2e95nrUrJFrkG+gsX2HUzq4OCNZX
AdfMNZeNZNrb2diJCGgg2+KjMu5l+MnY3A5qBkjAzQLm7/F3pVtheEGdiEPIxJrT
hAAyWKmX272bQLbm1RPftJJEaHKa4h2pKisZSV4m3PeyqY4SOlNC6dYZJ51qUxhu
61AFBVk0PKBlzcnwI/y0WIg1jfhVpUnIZ4U7uxrDv8w0eIirh883gHXgTpTApvUt
Vn6mAJIREy7VasFutN0g1SE5vQh4ZPpm6kDhz86bWcTb1PobHdfgkSF+LKEdHGKx
lZcIYv4buDTsZ1MvErUAjMx/qK0PJBjQ6czVcMGgAlUkML/Nz3X7q1TmWw80O4Sd
8C9fumWL6XMjk6RYXKEqMWOk4bojcKBKsBkY/1JYOcxsAYUScxb70jFmY7OCREtR
MuKwozWz0jlTE2OxESPbO2vOgox/Zhnugn0rqNkRNl4QaMg4UQzDwFpCzEQPjjau
EiTt2AE3MtcZTnM8e7hA9l1/9BIJO13bHx45M1NY9+4N+yt4D0E9pll2EwS+M3MR
tUqAoX3Wd7tmOq/H06DENHbQ7kTJSh1WeQ/ZVTk7Vv+u9SAuRe4AiPVazS5EhCgL
orTSw2VHTbWMdnCUmchlmZrXARy6IlgNFW9uu4osMosFnEAVZCZo/XDWTHPkMAtk
5lViKe311UOFNUbwoO/GjEnKtZy/YCsW9QoTfxDe9pTk5o2GZ3pkkDYi2a2X4X14
VaIBG6lRm8V2EOvmnLz6pClC2RIog/pEUvm1rP8BYSJ0XUlVtzInQ4t2tmWGelk/
zTbppS0J4y3sbm0EecyOyQW4IJAeq6MrPwEvI5D+WGWr1ACS6j47sLykywuLOkZc
yvZikABFK+h+h5VOPrdY5akSu5nxyoQM9k/mWBh3pR52D1LWrz40e+t9X0ATVLTw
K8f25ZQVWFdhzbo81FKJNGyfxSgo4eNxKZy2Vxbu5dnqO0noYddmA8T9s0orsoaZ
v0N+gG1yrz+1gFOj2GzRnG1p9+DrOHOGlfXVTiUVc5ZsyjXul8HBzxdP+fUhhNNv
fbIKzwNgOXVt2NySxI7AtUl9YpsUAN/nE//DmaYKhby2odsxSea5GjK9b/hvi6pB
Qr6f9IOoM+We7GW+OV7JoQUqh9+pOCjfXWwp2BzKAmROsWw8eCLZ1AJ1rk4YCzdI
d2njAHibHXWg4YACb6c6ii1Jtf8OM5n8heHJ9zkrtU0TkTUU4/VJBCKvOxnNjR7P
ayti1z6oL9L0IPHCq3IvcA1YQKAlWSca8J6hi7ITBoHCXCcy8Sj1BfUOm2PZ52Qy
NLvT13LDACVgOLqg3CtJ4WFHm33Wb0h8acEcUISF1HWLcJxXmEus5myuEbVKqK7j
93g+lbS6DC+U0O+ak6RjOCQcPvfwjjt6YjwPxWNN0JFe5DAyS5QK0I8NbQkTH1X5
SRflo4tmJnHmBCeF3N3MorjbD3W4Xl+Xi87eLCn/EayLHI/4nVG8qM6SVRUfGC6N
JqCtYPot5QSqmTeDztjKF/3fGSW3FwskXd/uT7T1xrNbte0A3FnZ7ehYBTkkh3Ba
NNktH3z36SXEuIHb7BfJ6KE4ZvGyY9KJrR/ZhSCCZJWajpMKKU3A9a4Ag97GpxMu
AEIBq0xxVOwIy60Oz/PeJwqft827Lv1+mKhvy3qL3KMOh6uDmW47MlI4ZY+xtzXL
O5CdMabNXNfIRPL0gOuK/92EGfG+el7hWgCpIMlwmwjJFZeMQum0CZgR96uIeO9a
iZOlT3oTAN3bb3Z7VSxzOypbXWPsCA2vWGAJPp8061Cg1Qj297hwGGhOKtHJenAt
dW3pCu61vfCqY04SbEjJ2uWrtU9hhqTajJbVJAt7aDVlGftJ85bdBBlgWJdv0NUO
TwNGSawCEXA3Fv3dInbpfDKFTHoy3EUG+kyCRcTnoei3/EFPkv37J4a+YIdnsi4q
qNmaAP1Xxu3A16+VXEtZqRmzgmde1blNc5u8byqfQZeU6sJUx9POCRIA+DBBMqTt
h+ObQ0Edoxkg2+eRgeVq2X4b0djKVQJ5+uci+6+BrYpUgUV4/oARAr8sq82EVII3
CC2Yf+n7sfUYmhP3/kERM1BmLPXhombXPRYQgWo2VVt3SnHLuWpyvHDr59Ps2Csg
F+HZIeRBABwFoc3vBfgj+JDK83EJAQ2OyNyDBzsBy/iSShRjhENEkWzWxpK+9/El
B1zGGJmuVttw1KZd7WLBl0KLpCcaV6adgS6IiwEMG+EGOrs5AH3UpUiCRGuNLzdI
IVT8hT9h9Cp2Lrn1frKRJS0r+wGeU9ex3BiXkhzkLFe3ovocY6Lr0cmeCbmmiC8m
O2O0nH8jkrL6WPY8BEGDeXq2to1jBJlHgg0talf/EzYgN5ijjh9sPqTorsnp7OV1
elKNb6+8RQeL+w8dB+nnAUT8KmyweudRfTzdRo0yCSko3cfiGxtYq50/wLOmgEL2
+iHFXPQrZxTCJafRql6ZvEXtF4icW2MfEkhHYhQ8dpPBt/FggPe6PNayNEIDcSI6
/Bn5wMopCUR4HLb9FBnSI+4gaX3EMPJN3OjJ/ciX62X5dhb8z1Y3f5FRV4/n6uJJ
70sRBU+Cxl4gxfJMMEUU+PHausbCBsA/H6yRDLyMwbZGtm40KhUlF8bt5feu5S3K
jOKez4UIqeGiTj4vEpCP3ndGZ0d03fKiw7Krl86sSNWhwOi6HZdKODa8CBFms27q
dMhJWzYwzGIgw2/Z7gZVMVNKXCKLf+5SjFiXGllFzQyjCDVK0cQfhekucySKtxHr
Tpy1tiG+rFb2AsWpB09Y2rMrEv83fLwG3wEFo4kMTGKYRnNqSHuccq9ozSNtHDQ2
4rd1Rb2g1Tp+XpZd4dtkFWsmgZCsIaUdqkAK1TU21dFTUx5gEdRE8paAfSH6bC6t
G3fRa62NaalXPxGSn2tqP2c6SuNM6SUl+Qr4wJYkE+7wM4eIJ5wCQoN0qEX1gO8c
5G+agjKfVnyNYw3wqvYlvYGa4jKaHRQTXO3s7P2VQhpbq5GwsBQsc/qGLt+ULpSt
SEsMuIKcl0QrVWZBZpE1PYFdwWj/PLW5yml7+bULjgU99PBD8clAmUF6zDkFzRVT
Qgo8ukeF39CjjOFg5I/ueXozu5i3aAxPUD1doHPBJdF4ncI2eP+XHdXw3Y2B0tQJ
rl0Fgfzn89Y9jRfae3iN6hLFlF2fUc/SekUU9R3v/fiWwYQziO2wdqAqNNi+LSTe
9vl1oPE6eeR8/2r1F401tMSPF6U3zT4k8UVOAeuvQaqfHNZB1eOCuirUXXmtKP1t
tC/191fxEBC6OLgDzq5uePeEk6b0YElMUmGDNmIvNRzCX7jG1aowoFBSGTIKXJ8B
+51zFPWqEu4QKSces60OLZcKQm6q35HRu61YP8eefn8vk17rg/NAEydaXVNivvgc
i7Bdk4/rXh5AOvqryMxqf0nQuk8fd7vuNYgnxNsi0oSNqdU0EeG0s/pbfPaEWMom
H5R3COFlnfvdQhrFeTnS4jfAn8LVBWfU2UJfC8LEFO+9clKYd4GE7tBw1CPHj97/
2EwkN7KaeY0Ycxvck27yqci9U4OBKJzIkck5oYGD80oM2CIqL8QsCnTqCRgaJxzq
uuv0vNikgsM/qqfsdMBaOkfrzMTzHnYIqwGvxxPM9Q+vOf9fl+kLc1DMCquWNRD6
0vnkLf2EpDuTHNNhBbDhA1TLWrB+Naj9Fq5ljkAyyfFetdNMXJRN3wlPFXpdpbSk
vW8INFEf7i8bED6wh2qI4tjXPNkYKKTsVxLKmgzUEZriWdx15UKFxcJVe/oeQoI+
to1ppQ26GKf6UzL6FRifzz1WQXSi3saUgJdRRRZpWTQui8AbdJM1YRaKMWZ2ZboS
bm2Yxy4PDwIW9ED3RWO6HWVKhPXn44ygCIAYR/kqvJXdb0OgBb0lxLzB4FFQzlZQ
epvFc/ovZzcMfZ2uJuNOyqNBAPTCpeKjppdYi3MM4X9Mtim2+4dj7F0+jZhEoQau
utTGj1YHIHXT04NrHCTZmjipEJ5WDwCfKvTfYVk0IUhPhqDa13K558hVuCO5/XeP
zLs4OkPwerLrqtPHg0RXYeyjpCLdr6t5SbExa85/IDBPW75g/1gu28C2V/gZizIX
AELoxEzLU3AnER/bihbco1JyTsbLWBIKwtrLIGJ7j2oUP+5ZjyhAtDmekdKF5gOT
QAdbLXpRi3sIFjOeY2FNvcOHghvW8Y7LyBOxTg3v10iZYTZVunP9FOQzM0/z5pUL
XnInhmMFDlTsk2y5vMnainpfKMXokRz7wFeUWwHDLmrr8sMTwynf9hbf9G8CkZ6J
I+g2+7wkOdDTWFovWI5/NPMznvWax6FwolLeY0i9ezPTQvE6Mpj/clVLbPZMhyPn
KFY5KgtxrO4M7TOj8Hiq+Df4Kskl12NNQC+3tSF5lGW71Wz0SmdLDEmHpAkfzMlh
toOwucyIj6pPCc8acPXxYsEDAh2SV4GYXFJFBEV/RqScWPhx/rIdJreCesUGhw4+
tBj+JA3DHrsSAcwIuilBfirW8HfBRgXbMxJbop9tW2kqPgZ+l/5SWOrACJcoXtra
l5jzvmoYC6A65Cvisid1ko3Vd941saEJ2nZtCQrmjlbRqV+Z0F7QL31iaKFqX48p
KPaCzBDMEY6uqA/6QZgzI69SWoObJuprAqz3CJtPSnXiXh1QT0Tzk1pCkCSm1dNW
4o40/hLtfJ+ijqEhgqiq2Aool5dKDgAysC91fJaazYBt2sRhqgD3Fw4JNzlOfsXb
qXzqlYtE3u4Ac0hKrL3pMPetWwO2L4u+LpsDghl79iTFrh96HOfcepDuQnBShrAt
/XS7m88jZoRVT19aUdlL2l9hyEjFjhWNLlkRgqsS+/6BV75qBjqvcJP1ioNUZljV
mWxgafFt12Vc8dwNbkNXP8HGn6S4wXXs0UKLN5VqPTK/cLX2/VVH4Z0BkBYKOBNu
PMqug1NgyNZtxqxEGYad8xHkka/TKQC7QVvEEkQ/4/aIcSqzDkUpV0pbN5F3D4Ap
qohfYfzXRJ9wJgsjR3xunB67U9hDrL13pDLz/WtskXIvEDyB1uNBOxYrWD2FpsRA
RkSRTQti5zAtUV0dI6KXyD0ZYQ8WItinOJN1V+ZTuaYT0TVpr3maHu4isRYtHfGh
wH9rS2p/BZaGgrsZt5mAsi6RoGk5Grltf1OHwya8w0PQLeTDR9m2DYYWl+B2bI2n
AVGHRxnRdpnFrKM2ekv4k+8B85AZfEfMvmYOqeHJO2c/EKeH+l+nAAlLSMz4pHmZ
EPzfxGODXtux1MzDN1+aaY+JtcpnKsqcWOmIQ6znPzZ4Okn2FgdI+jg9oCMsDWCO
n0qKNVy/hXGUEajSp2Cwap0H2gWqXwmxF8VhqBSWyxJ6CaMP1W28rOqJncWsJbp6
8Fztrr41Th8JwW0YggNslNfckZReX+KKG1rQD7dMB7LgVI7CH+p8RYMrcVU7zTwb
T/IP2lZ8IFSLp4AEknf9sReVIcv9IUagPM+X8wG9y0HGRK/+glqT3chhM67MvENK
NOsW+OHHMpPknfGKH5JDRdYQhWCC4waX9RXeENIxR2CGhejWICem/nE/g+rQM0oO
GFIMDtuLsx9af01lB+H6g5bUok/cpiquZYcb1FFYpeyDhZwlopOQmTD+H3kw0pNP
Y2CXblRJpqg+m73z7+OEqFBzu5mZ6vE94eq936Ag7WGfoWJfPDzRVtkLP/fN0Qgk
5z7kTlG0NlOvjs3dwq8/uqaI93c2UtvptVYNG0tJaDyj8a6ef0ynj8eAgrHMPrrF
sicBpneWblzk99Lkbl+fNVux8InHWEcWGlG9z5xankMGqSAkQCQVbeRlw+rxtgvd
THuZxsxKTscFJPv5e7t8Dj6Snhu4eGPx+CkS4nXRG091BS0XwDur0ZaoI9Dzgi3w
b2HiyUZX3szRYTsNieFDnbNoZNMpVJHGATEn/6iby/ZOm0QL/Pr18nC+ONygzl4i
fxIQ0FEEpre4IT+FtGz6zFjQ41NLYOw5RPLCDMhyaVwzltkVPOLftFreP3mudXg5
xkoefQl5fe7yHUV7wHBZgRa9V5Ylh+3ja6xiMJLUscKGxkLqevlIWfwm+yE+xDpq
PkZgzcbNWOURG8liXxcL/s39qhm3tXyymvQ6wXr+2PM+rSPE8+yyPYJhw47HPBgZ
rPdoJLZNXWPWBolybkRv0u2rjjSWTutFou5nR5PpN5cXhnf/p1RXexuVZIQ47Ynk
P1La26heumoWUGIDuwRdMvYcbTxRSVfpXaaKJXAk0503M0E95kCfiKaM9/IbARP3
QfOfMzmDygw8aYzfqCSXg2Y+/Ni23Oj12JRWxtcEn6BsX1eZkJw2ELOp/IePP7nh
j/ePKK332zZcj1rAj1EjmAZ0MQ1m+JTjb55LqwtOpB0/sTnPEEPa6+iZuCQ/IJ1G
D6Z0PkXelgm0NfAp0DWmzJckqyXUD72+5HdzUCjIA3cULcHi7p80VxSYw9jBPAUa
sFDO+c/uYbWv0H81Vtyd1M5it7tUA3usNd9fRPkkRAoFZcRd9tb9JHxqqfBbEzuF
z7MyNHlVFjRtvdtyk0mvLPyrfU6A/KBX7wmF+7yCIsMJnw2BzL3/1n12wLbrB2Fc
2J3nMof3PjCJN7WRS7WYgfEhr09ES6gpnA8/Mnclv5YJkvaSsSKY7qFXobCaG9TH
hRXKcj/WT27Vaha7JBgybOD+fUu8PCcWQ0EGkvyjxzxobhlF9FaNpPKr/FHU3sRz
IC5A719tt4fzZFK5PlaEAgVRxsRNqqAPFbA/qfNkP/fDjUF4/8HaBvKwSnsxdAxl
Oo30TSQQNZK/EGLX1Eg3pHc90EBUf+8JB+M8l7ISWOl0T6kryOqfQo6wk9k6YQ7q
OS3X/7s3NoTfPG6LBeEDt6Mc/hb5RKv/hAKh174VDxCkPnt2ehcn9yyPznzLuqYU
R1yPTD0gF+fGrmczWDJFf85/xtAZwyLsE73HLu7CfJ9kAXdR7qhxH2+VVh2rFXDt
miMRHOg34FGV4H621ttnQRCJg00GPbVTl+rMvno6RSKoZuMHgmAD3EOZYD7PA76B
XSvgvCe7MC+jVyJPxmAhlaTPi5DmKLQ1XIonNs2kcd5ciTvcQWktmSiPH5+SN6Bf
kK+TBYjpQ5bwZbBag8K8Kl+S/qgU1MfCtzUrr6IY/hZlTNs6MSq3hu51CYLFWuRw
SwsVBl9F8ZW5jnPPTIESecMxZG3umgft9sHlr26pWIrPva6mK4Q1f0pKhocBPFn+
kwaJ9F3RKqUzZxA9GE4/LmJTR4Hk+TBwkgbn/rKaKSa83mVnIwXIieMoXXFGK8jy
mAN3RtedjYbeIch2XeJ2tML2CzdoFHntteB4IStIn7h3RIf3LpYy6/hyBp9TOOee
SKGf65t1Oz4eewomLnQ4vswg6ESfhKm0rccUm6VIubbfgB1GEG7iwhMx90r/hEgP
BG0QQYd0sTJ0kMo/z4cjbu8wXULu5Xh6u6hrs+FexoIgUxDlXK8YlZdy9voYORcl
MpNIFT+ro6f4N7a04wDjH6f87Ut3yo1333vL9davAMhMG7Vp3V+cS42peffgUWVn
cLKUVoTqFMjF6Uy4+TQaV+Lmb/NhUY9PgivTInasSiDdw70YeEHGQ1kSZGUzvp6o
0ni9HZkJrNyKkQQGhUcKPazkLpmt2S6574FTSE/yfwynH7B3FySjEDJ2Y0Yi/0zv
a08+bhGQNDBfkmgZrmyEApyvM5JM/GChDFP/rk2piwWPhwW7ad6C00MxjBqn9Sdf
V4dP0oaY+apklOCunkGvDInMG8OkLVFKLkyskLE75mOrwUze55TXQr/MtNtcQuDK
xbS0ib7vZ1sIopZYUWHO+NFA5gSuLNfZ22CTFyrfneePfTial7hnfjXMGEU3nm/V
XueczaemEUZueq7Vvdrt9XHK14mt8qIDeW8WAneG296QYq/fN2/ZEnwnzZNiVcfd
mSJVoXuvfHL+W2L9AVqhtFODdyAOL0Yi/huppCREjjj1RGr3fRPHL6VzmVBCmUMO
oAUzJ5T3u2Uno/LyDbICnaZ7xd5rtssV2qr7fXptfpNJdj0EpPywcpP9cIrgViqo
aqAAsWm922hoKrdCAdeJJREuboveCcuOnNZxwy8zmxTTxznFu0IBk2+biOzK1Y9s
AOedqBX49IJXZC2wCmyAfYfbhXHlb/0bWPGE8nfhhdFRaxaasLUeFNblVr0ZwtNZ
ANZcVeQyQqGStyzhVz0iTk4P+dygsdjKAF8UYYt1h+Tcdqqa9A2i+J/wVtV2oiQP
am4vHfwpEyhojhx8s89YCosQVGxt2sTk/059bk35+KVqb52EH/modu7lHz83IRFF
2fBMhIYRtSwpy2IRplASynONiVLJiRbbg4Uvk1ksfK+G2u/hUvRwdSkbKf18xhU2
Aib4/ZMqcp8HRjkDMxO9BjD4eSL+1Lam/Y7yWoCWi9QqOw7MEr2vGPZJTTuYB5DG
R90hfbi4mOatXZNuchnmX9Npvqk08zXEWYoZFFzWnIWb2rLfiJx0SgbVbCgf1wDi
BsWIuO5W4i+sKjV5CuKCKLfw5xNqpqtEDpnY8jHf6LH2lrZE3zo37H+0UTYSqZbi
4O22/fQH/fHS9vTLOrRycjsW7+zsdtClt4jK7r2/q3rzG0lTcmMjK8zVDroyqvzk
UDXDC7oTryHL9Px6X1lgGnEPFIM7mi+Saqdpf8rBtRfXPG898yqvtJAHOWOPqesp
3svt/yM2GkqnSepQ0ogqGnu7sKe0Y9jdIxGtWIV7O+AZdXNnjdcM2R5og1WYnIs9
UXeejqxaTTl+Vt6gPyVQOUdsgRUQAT73BQO2/HkAbSJcb+knPAwa/5UseKagaqan
7F7KxEYolsR0CMTngaj5qHApwFEjhMnQzNGs2iKc3naoKyRYtpEOSHN74lcc7ROi
0cc011rGMYgbmgqm2JUDXcmZNcrcFJUIRwKpZZQoC29bq69VJkYfN9435HG/W20h
qurEHm79DDyUWoD1ksqUDnMWtTDtHJQVV8pK/m0eyDiEik433HwdVPp27Hjv7vKo
gVLs/gTg1TLM1vnFIfKZP+EexOM5TXcTRFbwhG14NE3tdfja0qLIImCmpbNusHko
3C8sTQoRQcvGWThTvhzcfzwHAOYPoyCLTSFYxYuTltghBWrOIK6CQT1FCY2KfL6E
UKTdsh+s3r8OKSYvQHuMhBKPepoyPQMyoXr1kJKAzYo9RyLG03bqLkW+PVR9sXq3
oOGWV64SadIdTga6e0+xV+f6aJQX4rhmd7nklsu/6fl5rN4tJm0UF4AtuDdWe95K
/FkdU1IjruLZqLhV4ZYuyfOaxqHjG+HA8rOE0JTpMj7Sb1z1esf1qUSJPXrHot7R
j2upUbmPkjLpN0R+WdHPcU7vt8eRV7vyqQL0qHxQqdRRYE6biGTiuMws/N4O8W6o
sjaf310R0nIWpWnhMPPQjodEmF5BfI6y56B42roEW9Efo/TdXuhMFwjOdXENWcI/
/kiaqwZtmyfcSa6IQz646jy8coN6IJyB0mm2pT7NMNMZHZOlGKII+uzBr6Deo1s7
W3lOXophFBCWPrMig367ojwulDbg4xWVWGVNXNj1WTfvwovrk11l7fiTY5KyITNt
3qb1HDQ5IM0LTxBC9pj6HkxgWgxQyiZewFa6E5sYRRSTp+xILw5kULW6efJGNt3X
RgO8CAvtMlpt3uBbW6PkRlgzxvnuUB7HGSzrONP2Q6Z/RwypeLm9eUk4PWowctLT
3QJ+SEH8ikFeAT/gzy9u1Kd1268GGBv2YyxihFztWuEvGKRYxFKNpNkHB5tpWMfk
rXi0xOPJ+9Ly47d0NvhwkCp9jRX9FG9SaS7yqAjknPeT3pPCIl29zvAH7PYnV1Mw
dBUQaOrx/2Pbsdjfn3S0+CeC9hRKgE0qKWV0WtsZZFiCOvuGSNK6jfBqdvaO55Gs
8tP4TGTDGOc6fN1mZHMhb9+oOINoonSAD78LvOtK9lpba+TdH3x1Tzk/CLNI0x8/
Hhgx57NqXoms3NZc+5AR5lo5Dai3KVJ3TuoEXN+pFIIkyfBhG5S0pCHce2RfWkJu
I2Zj4mzSG6zkxtQ1hQK92+T+FZjslXFaTTbTh97+iEnKIcqlwKrwIdQEuMIY0AcH
nWi77Y1/Fmiq9KQq9yVg5BzI9ZBcEKFirrSnCX+7vW+8Baw2ifsCK5cfqxVXtdz3
CIb/QWjhJJqm8oOUp6xvBgjfvKskw2I64BjqWfKLQUlvIAzK+blYG/MTtnbW/Esz
FRLWXI+JB+Ce+usKvCkxIa0sa0uhdjZ0Qg1Jlj4nN2Xgz/l/r7zazIfsgOikYvbt
R7exJzQloWNEkyjxX7PDPIEc1D4VVxbbpk+VVpaj8z9YjhbvRxJgjq9bK8jJyrwW
hHAxkzXPjK9S9teLQF4bnFJ3yeLSdMtK4vhOO2BKN+qQfThv6j5XS5hk2up+oNW8
OMzwS0GSg55PmkT3JoGNFS8XmN74ZQmIYgSDeG/vSTGQhJEqnO1rVzxa4kcvzDYX
IoKE56CZoLj7BOw1DtI3BAlmK4xZbTApWRg0JbPhbfxQSZtg9zO4EwgK6jiv1EFe
fSuTW1Alwait/fdAx5oqAMJyuPZT6IL7yr68flhpNax3SG8EFYImInDvNFnOZSax
rZgExxRgy/TnOER0+PbMaMVuuKLtiYdoEaAKjxK99TFgQc/CFRZLBFCvbjV2yRDz
AVVTRABJzNmaRbfmJwQe8hSwGLFol1b0tPtTaWgyREzj7n3ysUH85hURFmn8ul6S
5b74BfQ7pgyOAx7an0h9WF32KdoJkV6rCIhc2dBA45b61GPU9VEDboNp3EG0LuaT
//szckgnzvyV44NKZPqkjXquYvJ04hZmeJJkXQI6qj+p/fU1QhogXMc1etLRU+Ud
vWVetJN4eYHPezGrr/RWVGpHE+riwLLCJo0W0gL0+8HZvTko8JCoes17rzSUu978
0dkxDajjsPtYXmbGcpshLHUXC2uxa/qvuzXtayt0K1OQsMjp9rs99kNOobs5ndWY
zfqQRuhtNDrTZyePPKWprN8hT+tscSIcLenp/z3GP4y3BWimaAWvRaM5IRjh9KiQ
O8shG4cfXM7g8jKediRK3p2FsXPa0TtG1sV4RuhvK/gTW4Glb5a3+bp44QVe/Nmd
xwZFXTqdcRl59k3l/IDZp6FPaSOwE0XPevsbiMo1UF2aVCmKWAOfnpd/HviEWFG/
a5VDV2NxFPt/OISOMaV7jma81wuE0nSupr7gkXCePQ7/pf/yvAerBJ4XfJjy2Jt/
Az8ZPut3tX6Sjh7v1WLrOU/7CRCZuv7dD70qBnqE84UEGI9YhMjbFvMBOBitYXGp
RzzvP3XBzaRWJ3MU9CzT2pg0OOmfi3kS3oMiwjpNHccF8qHb60sj8oluKCZCeA6T
BZLdmPEnnzC4Jm0dJNGEnwi9X3eJ3HYvhO6MzooaK3NzJ7OFs3uHQziUAVgAbeOU
t3bBeFT4v4TB9DOjrsjPEK3nJqTbi/vZGtSBB9zNXl4nDYxunPiry/jzh/72DDD7
QklBM4LlRlsyTkfnulzpz3CJ8faccAMFbTANZThXc0ploOvzshje8l6zFFXP+Ak6
sMe/txroZCA7hC1rVqeU1SF8AaAbV4eFMIq1eOxUO/JXC1/hCe/eLKePvLH4bZH1
1JC/+ZLhp3fgOmb3JEOm2nVtc1jJuiX8qenvKReO8ArLfr6gunHxcRjDONVJw7Bj
aI3lYx1IY9CaeLiMLcosztw6pdpFiGJH+fOWJACpQLg6PPHpeImqFAX127k1N0MA
tdzPf8IEsIwWKX0kSwG/QIDPKRupr6iUHsAA81/Unz/ixk9V+Nn7CiDmNKp2ON6E
C/ZJWCpyn6gVeO8RO0KkxwR4v3oU/d3DQxdmD1/pRybn4KQ5EiYJ57sWF82k1pzU
FyVwdquXtLZ3zFJc3vBpmPem9mByXpCee9pUgHlaXrFgI1KiTXc+0OW4s1AWq7XR
dVb71uW3seKcRymIdT+ff268A9p8SYZSjr6VbF1XnHjlE5idny2i/CdLHzWuJdM/
iwFevhvTw1ckcrHpVw5Vq65HMumbRvGtTSdDL8ZUAJH3l83RdtsK3rx1jnoOO7Kx
UXXOCF3npzf+MeoJA4PeArhjPPtQTaJVj5Eo1Q8Qzeu58xkBWM9nD2s68+eWwq85
5bYr+hdFqPpSZyK1L496T0SlL2aEAbSMxWFRVfCA3MlA6KYLaWHe1/Vbbb3bsYrJ
yu3WPo5+eBcIIFmJmN4TI7HdJtlkUS0D+PdUvCpOC3NaGKtVWw3CSWQxYd1cqng2
Jjysp5lmtZS2Q26HJ1lK4wA7Mc1BS8/1NeWv9wtPdJ5uMBawiWoyZ1DBbqr060TD
E0cwTxCA4sr+DvEml0fSdCQpNpvbiHhmPu7XQoWWSjD7/PW7qpgLTLMh8K5aCDHW
ssmMHIc7B+EdZ4GVGewWvmJ7Anmwwf6zyzr/EiV62WwaY5UFJMX7UfEA4647uV0Y
XeuOghxNFG5QSmWpYGLev+mzv0fkWVPjLzs7uNUh9TcnHS8vHwKMoU2UWOUow5qo
pSNduSFVORdM4E7ljM+x+Gkg9+jM1SMfJQxziAO9E7sRPLLea3dB83YiGIMZI8L7
ApPseHNB9CRFXi9ym9UVJ4fRxof5DXZdtwcaRCy44PLrLvJI8mS9m8WpWbyF4ulZ
7AUt6Or1c3JbOU8ca+8FOUty3gdvHDxnFWapjZKWroBIvWiR38kRhIAIf60G8aay
GZQ0L3Y4/Us3chgxjLaZDPCQk6+GEHdC7K3RW/zckhg+2+cffa1gvBjMBaayyS3M
tXR/DAFeKorULYdGgiv35Kw+sUCTZUclBPfjzN1wFhw5CB9m5IRcekMTknH1Bdx4
nHeorGnIxHwAZbxHXDaiTOyrA4jCmFbC/oGpkQuzEfG/ch6gWiikHQw4LLWFOP+U
86ZPIF4/dGV2I/R2qgHz62DQgTqrYggWIU7jWbYmXiDEU44yirmdCQQbzBiTP0tX
8k03Z7xU3cFxedkGBmUAwZDDFBbM3aG4ucrv+9MCCqxxcuEknAAPRq8XZF1/5zCe
i8wWZmUeBXO8PsL7fm7XphZngRQSZbeV2/TIcNskGW4L6Zq4xE/zNS71DoL9eURB
ffO+NmX+8HrfPFSaGL/V3tGclCBsJGFRu/A6IKN5fQ1RlfTOl2GSFB33XojDMYL7
L1d3nm4qTbWlOaDFRtafmRnz15YzQDcvMVVkjfL6NqCk0X6i4XwPfkKtZhB8cnFg
Pd0HPRW17bMzzJM8o3Pez3NEBC+9y3WD4CwdwareutKHkQ1o4d9poC8y52Xqu+be
GQvzIqHJG0rdHVKJqf0O84O8xSHXKWO5orztXToDVbSZDlfCUGDht3arRdSjwXvG
rn9lg2gr/Q9eJVYNboDI3URDHaJbICk2JYBD9cz1xWuyx8kSPk0xJSIiIkzcewJy
GRThO2qeYrmQtECfsA+l3Nxo2axNNVzbJjIn8QCGCOZGb4+gIidsb8zhyBr6xIPY
rEttMOYnrVfvkLH8JyCKuo8uNALfimK9rO1li5MjX52OYT07BbFXPngjiTbOSNSS
eX7kX4OBUY4MzqU5vNw/RSEL1V12tcAfhu8//HYy4SMIMOd2eFvGsZ/EP6e0sSr6
B+iD7v9By+9KkFhWPfctXPzlYKtuyoL0s+XbymnkBSmG6H+DyOPBoXziRh23deAw
REROlhhe/YPmK00CX+daIoFwMj1VO7ywuVPRUsnXqR1W+U1ptWjnx6RpYEDCu5tO
CtRIhdRSWmRX3dCIBUhHF+vyoj7uINuWBXv9m6pedGv4jKj/4GTgbzNezNTxyc8A
WLvajHx2Pn7KrNSDv/REekNS2UXTa1/VArJFAXHB88zJZu7HZeywGP06XF2dhzXO
+uXQwA+eXor4W4AbqNXXHTjz2tRzmBo5twHUsQyut24PzcXi0Oi8WIVN6tSvQYxE
ErHlza0UYnTLJED9eQpbt8/9EC9AxCNnA7deA0a8DJqzjYc2fKVnDgWVux5Ntw3e
Z9AFTu9QYbhh+2frmqzVRGgLmR70WFmp7Z/4xJ4P4n/WxMErqdGrpVUqBcP5zjXA
i9s/rFztyYoTGdWYGXxusaKfLVk9pCTS7Hiz/wDWY65HaTOMDg7CtpW95pt7Nxzq
YsZ7cpH1+0ErKZ67y5Rndvk4NxldCLFZMKBXArgJd96ih/R+0UUM6Yc5evMONkCk
GngqrACLT/rvTpZ0KjIv9njE3U0GGNBGgKhgf6U+G7Y/7qzyTyFFFM+4FafZxUOV
9ax1CrfVQSh1XBeq/NNiejjDBnmd3COCMKV+Yjp1qEIgH/YxJsT9WWtLE11q5wNM
7MITzKcyhqBS7B3ZHzhFGmFrLaLQe9sVJGQjUis7stVTClbIqu0NlcCdtBU8k927
8YUanxHrZq8qCsYZFPBaiQw5K4++T4+Ck/F+XNrGb6z1pVGh55emhaHnIGJ4Yk9B
8oYoEFgKtLEbUFAg6pMwpm5BarVuWaXb6BZFQ4XxUZBvM8H1fCJwmbCp35vDkk53
A97cIgtKMeUXeeRQ2y7tFoj7kx9EdSbUbwG+dU/BYuTJKyv4LphsBYnGpJIbC8ii
QOAIikmSsMyybkLJa7fHAw36QLddKgN7eEf2EgrKwLwDWGZxoun4W/npCWhShh/s
25q9mM37fowGVUZgUcOuGyxGlPKnHDB7qTGC/UFYYAZ8qK/ZI82WVApNVo0kYs3+
k8tY8XaQGu+VMnWjtjmQZwBIoHAtQ0N6puu8jNQyqOXE4EOQcjJd0P21XwlJk1Qy
xUdVEGwxI/L7fZTmnGQeFMcPph0L27R3Ug8hHf0JjRCaxYBvNODSNLNVJQsy6Ebq
tmvqPzAFS4XaMNF/ZB2sQVmQdtUOyGuZBXalXMytDJ87xMvTSnIZ+i+j6q7Nh0sK
tjU01rZZM2ntu5Vgn0qAqGPlLAcMVgT1jt1K2PEsa7pz2qztS6cCF4QzsfB4D4pH
S/MfcbxxKkT0lYVxyqf6e3iqanxBjvnDtGNqJRbbAr03Hn9QyhhVAyAnxY+XhyoF
zZQDNuWxAssD39QiPKVD8Z6WzSuaLRE23xt86E0q/qLkaCJGNOOtqR0heUPr3WJ2
DhCzBBREOA5ntkaG7nN+FNh69UWqQ5/8pc+VQEvVK1eFLk1EXghekomWT04N3ZEK
tIOieLJmdvngXIvXhBMYP8b2L8LbMjCvzZXVPH+8qBusC0R1n3SdJrzaNdE+tGW3
vLdQ52eL8oEzOVcSKTHkFEfijZtf2j7tSl5pKf+t6xn06mvsjVUz1emDvL2mRrZW
M90D/Pa74juPZDmZrHfpGr88hTDGQguRNpNfodahFTND2gaxp+cEpJutnsnGKV1e
isv83v5VlFGO9kIKqJgqTcI0+1eBMb+f3B4jDZoqm48OLNAEjrUDeaL7qH8qQWEn
QFk9LOeRwfTAqEyLCf8ln1WPLB8KxlzBapezQLwJ6kDmjGFSdhiAl1OEaRTiT40p
vJ/fSDu8tpdnQFO4e3AEBRDDsfdFdaXJ6UC4WAgi5976LOTAo4komyJXgTJZ4hyP
iYAGd6vmsFieF0s4j6y0FVPgClTEUP6ccmzB/krhKjx8d+9XnHpWO0odM85mI92p
iYLrvImtikidzFEOMSSKknSpbFatuZPJJPKK5gFr9PfXAKJ/dLXnjtlv/4lEcNdD
vLUevssSIkbOlvYdkIeeJQNU1ODW2WW+ykKW7r6yomp5iPVhxQMnLCTnINaBP+9o
GKJ1rAjcqIwbnIROqRjFik0qM3N+ScLQse+HM7QfPKNwCyernW5uNdfcnVntoPkB
WWhWgcG9EOYnKHCQXSZyuHpQyWGTR8+yuMHMl1WGhXQRLxJrY4f3dm/ztlywFynt
6XeizjNEer9IB/DPgYHvzoDe7dthVs0GlaiRPrBIlY5rTQUPDBfZYCvmt/S1IZar
Igx1nCBdWDOeTWciNym5UPsbeCt4baAPpjzqnZx2XmdzVJL3EDrMWYQJSQM2M0r3
6J8Sts3L7KCFz3YuZE61WTKDspAkxHG0Blnsr2O5UxxD5OzqbRN8WC97stJNF24R
OPdqZufZ5ppxIeWJRfKIm9XlMbk0Km/xev79NEKEWFdV+fy3v2xJn9pZE1HwfplL
ENpwQGtUSFzaEIoxRSQ5fQwhwl00+4XuG32LELU667REK3n2MJCF6Dqpksk9QImo
t+6I14gQhVZJXbX08sOQp/Mwt872HATZf7fmF/3Z435rfair0D9eU/cWAF1sUyKP
t88R+X1hBrzogA5sScm6VLRp7/c7nnE0D6Fu1qy7U91RP21C87ctkygJ1LXfOcyr
zTyuZ8y9n4Vg9zH+tVxfSAYhAMyXUnu/lEw8OmMDjjX+hcI0+5islZTC6OCdwtD4
qMLYAgkUl2VszMX2Uuf7ggLzm/rYhxljADpabSPXBQIRrLEnba6RatVOiQN/pNn4
ZVGR8NjZGDO3TBxt+DCYtv3sYJ5lja9XAOb5QKiw1HfqpBOCp/GSUo/AmCKKZc/U
S+wfpdqw30jnT5WsytFEdN42Ay/v12MF2/PhN0Nh+hZd8po/RaUCmUB4g4rGowPy
BfEDEJOBC1cLpynKVtUiOlAKLgL1QlSl7asmSg3Oi6+7fgtW1k8q7gcBQScoCcdY
sI55QeV6a6+/5Z9zAXsnN7pKZDUnSl8nfOQolw8dKoPGL1t2o/VaqoxWeJBXJOkk
wreWSioT9Q8WPXTJpkEsq21NqwXbFCxHXtev1iTJpLasRf6hF/2ap62Rdq2+0iit
YtjhxZRsiT4p4S3D/UZtZ8HrqmDObsrQXOW7b+2Yx8p48FrGAGe84PCrpx+7/yoZ
RV6JJxglZ6psAQmFE+awDZDIT3020FNzXIfLtV2+8kkFEqqcTPwstskccL6Jcih4
cM8+faObLBX5K+vwlxAgPs/4wYIJes9u5dQ8poEXULImyOTGA+TcC7OVNb/w5uvh
KI++e7LXFYjbGpVrB+NMyv4o9SjABDENMRTC1zWaZZXfhdNq7emML1keYGUJhWxL
XQb9ysMhTF0dJvwM8Ix5Dyra4jaOF9zpB1HfiII9mgg8efL9fnkryxd05RPH8x2j
qzXZ9aPofzcOciQJqvzO6CPharaQosY3bloT/XuwCjMaFqvmFeVr5mO1Yn+75WXP
e9mkTuGRZXeAptMXqRWxq6cRGH7zM+BNZuyMk//Hi2RpfxHdfRHoLS/mY8wuuzdc
2ooKeeXoK1W1g6kfBXHOLo93k9CFk+PZ/N+Ap2YygyfT6TjEePw4t/6jUKSkzvUJ
grKxUfwnMPLHE1Ex6FiaWHOX1jv0W/q8hLU9A46PU1N/TaDK9O98vhFoVtgIDil/
887n0xQ2IP/5vNX8cVNF2jdF+lVZiCoT46RnlOXaY1eYppcQmLRORb1aAfkiMTj7
95TRpB5lUfGGS6RraIYAVsuT3EoJdO1qUSRJq+Wz3TpOKxeL3UcbrO9qHh2nkL1t
GU13jDcF33cXGPTACBV2/fEAGwDpyLI+6RWSM/4I8kAZRbMneTiMhZz70bds78eR
lu6mVydCGM8obOb04HsWPVzZjwu61W/lmk1eSXsk/pztBCKHfvcbPQds7dq0jemx
qre0AJ0VugrfEk9wzWGF1DjcGgi4RX+4IOH55PG9ZA2WTgNKWzOaFUMkkaD0HKmE
6i9dgpRCuw/pCnQoaEynKj0NIVeaDE9gFC9/8i5dj3ijY0Aeu48Mi/H/pivIw7BP
EoRZQZg8nORRI44D5Jso/8kqfe/ep4RAnk+Odw/8A+0A81X5151asBi8WhRuenlc
remDsI335JtCgf3J31ppWn7NCctFzFr/pXmqDx0SAUTE1O7cWhFhH/kIlHUlofo0
L/CZ1gkNK4BLqkdfY0qNGwl8MS1JmWM/ZRddQtBJKWxJ5tzdkOQ+hf0Z62NbhmH7
iDmUxeGiaCvN/9A+pMi59FTskBTT6Xt2yQAl3hXCsoWIn43bpzclzY4HckPH42To
ibsq+SvA4MCmEP7Jr9Yd5INeFj9KoytmpvthrHGA096wWxMAmxFLownzuqSMTtAG
Oj/A5p0+EJ8jS8lCY46CHqb+gBozElFCh4OldVWrS6L0LD3Zk51E8SQ4A9HsP1//
BwcxDsDWx/KBVpUWxX3oLzhQ3lKatQ2A8R79Pp5rsxuplugC7gIPpanzDBfRLq83
jgIOVGhaLLhuIgHOLvU781/H3AI3wkxb/U9S0QLIsghl48u410JiafQ3iBCDKjK6
eOc/gzzW//pmcoFaDrAi6/rg6ntOSuSpx7SCoDFz+GYaxKeo/8gQdOP9HcetadH2
ofYqPXI5cVUHQjIvkKq2GX8BislnBAUDbWXe81N7AOSofbZKVl2hqHkgV5tL/Pjt
TKdDH6RJwikXc4lBjwtXbqUSPros7ydxIdyFDhkCGJZssgT7Z8+t2Nzl7+WQzrxb
AHzrBkmfwbh0alGwy67fr4BWHqfyyWNkRtPfdPawswk/dYEztNHnqDO32G5B4awF
sKP6Sn99fqGy2vQIzSrQP69/gkynTMnUyl328fUCbNXPA/kQ26ctLf4qfgRkbaRn
3IBKiQPkcOz7WnT9Woz59rXdAnPjuyAoVWk0qA1/hUkINHF8pQelOVaQVF8C64dm
aks0KqEZjpq66DEkzY80RMy58H9KoupaM7EoX7X2F9dvl4VtgntEwUG1R2RSlN5N
B30VhFDfA0wQkrU/N77sJkx+bU/5l5y7kvolfualFxuFEnRYIHYVpBl3eME9NGHU
RaGZU+nxvxfW4Xbvw9atLFGGre2oXPJjaW06EbFwlePK6V3Hzzk4VId2K+/vAHCh
Sb0IMRfvzUd5DDzzkJpTMHo5NAZzPLyeliAOe96nonxq6rhgeAmLe4Vtl/H7pEM3
lrGBK56PIyoBYTy+bB0Cy/2j/GeWlnnhvraUtahq/yKot6XRcORMeWqr2SkNh6sB
tDxid5g/G4qB3kOMApV+2AmBvy73t+pWw8c6DwUYEcnlx9CY+rsKe0DFY80Fhm23
OaqAGDMbb+tm5vL3O/SsOTTMnIJBdRXXQUFk41IantMJUuwzSjarJpE6NnfuBO6o
0//IymEy2DskAypvmQkb+ilkdrGYdkyCZHhwAb/eGMZ3Yr17ErCIm+b80qEvE+Up
lzBlZCtTQZmL6ojWO3tfHTvVhcNS/zZdAq4Nx/NHLWBnGkSreHP2m3LkW9YAozMV
VbObOWYjl2T2Eu0DTUKnDPzyJ3KlqHzIcJjIY/NlAcyQqVnbJxLcDsT71rBdNgPN
sGAxBD7GdL0mgkEjABnCl7e1B2H4ahqvWBqBsuY8nWRRp/RbiLch+y3vxMVFK1jM
P5MmppErt0KMxNditATWQJq05B0DKBCCO+6ZaneIkQZmFo/CpiXblzISNvdFh26Q
x2QJaIfvqlyfi+eJ9lC8XM2AuO9eSPl5m4YxIPuFo8WXvh43PMiuEYo7lMbsRmF9
WewR7aI9XwEABYL2R2gJ2NK1+DnZ3vMpuwhh4dV/c8p705aQdsZonqN5LBuY690u
RXRfucl30P1xyQn0SotzBRV6ZGQfINKkQPL1vVJSajqRP1lRe1aV1Hz53bBghm42
DTMy3oLYRKpopiki1yySCD6kIDysTixliPZ6pde0ye5IFKfTxmUejUhcFWs20pj8
fzwixVs9dfKVlRHH7MOFdoyucT+mMH6OJWHXzcOJIvh2kp6qj2lyX8Fgmz1+GhGF
e4/3BJEm87YaUf9Gdlgw3ODuwzs868b3BwGjPgAlPSPVNbznxh36pt3hOGFLQhA4
lmqp7QfTzWyiCLV6UxgQtBxUfm65vb4lSmPumsQZBNcOzzj3dErs1jHFJP0eACIJ
U2KnSIWOF33S+Yo+t/JLSucMFPhc+rxR6eh6qeox8MdFn7E4x9EIBEez5etCeBMU
Gkif8RPvN6p90D1c8iFPGHWO/IOIzVIvaFtrw9qbIrlmaC5ZnKWQAlBXUyBqPnnT
95d42lQHasdRC40Me6TZxdqGIzwDB2d9dxgnKQVb/o5wajOUJlOk5NLM14mVzWcG
t7tOFQhHYjH2xE80hOBG+9Qfbf3cXh/T+m6PN/kWb4Vnl2FlmqBVrqWNovnV1LG/
tWVVdTtVKrbklfl05QMSqsTFmmPkkvG+pF42Jk/j32jWheN4wgtvSTjW82pHqfBp
FdAbg0sNLD63TAF9tDv3zB3QIlvzciuEEMGyUEE/BqCgVp1R2+YgRfrJy06/TClD
nNjZrNoP0M6XdpzeppWzwk+KDqcB9dT2wiFa/jwcjiS2EuLFYUSwmqgVMG4QjZ/y
OEI1bIS4m3JJbgkGz6Y7cL9T470ZflRE77i5qiw9WokhldAXhvmtrDP6LfWwE+3T
LVLUHRibTaQ9adyH9Vr+tAqpvN2qnDNZmdsC+cQtMe+xp/YYVeGrOzyksXRjVDDq
YPVYaav0qx+xVlawdvd3zHLKpBk+95o47OV1KkE40xqj683sfVjk7dH34KBsSzfT
tW3XCK01WD2oa9sW7iQTtAotHMHoJ85pUom8SwVRARQl5KlIbbiusQgfnoeGoKQi
3s6Wzua6QmFAsWKSIEB75EvzA+PNDLdT1riAmG2xYGOITwti5th36rRdHETD3LjJ
MuS4zrrllm9LjcGPgeJH8UHvv3OjbLgz5zH6mJWBR/MFDq9rSd2Uq2RTlON9n/cs
rlvYYka/+npLxokG7bYg6mw9emguFfFKxxSpcCBGs5YPG3xRsKl27ahWXc3A5nBL
ZidFU4iVB7Zwe4iE8UwZ3AF6k9dur7lY2ARgYJ1KOOzy3aOIt3TXxgaVnGOntvoT
yttAcoJthjrLD7y9wf1YU6DVW5uOdmmErRc2c09OHu1+58HG9F7uZjreBv90ZDLp
jx4VLcLQF15Lnr+yjD5p87jCrfv6MMthuoBEyxZ05K5TRx8jTDr9mSbbpc6Nt3dg
+paqPn1ve3YPSOe9fMo/5ypgnSlC+Z+RabVQwI+I/sKP/3sn56U19rUyKcEyrNp4
WOU0W4QvqCvhMDayuLCuteCWjo4UspXi5ei7cHqCKcB8p0N8WfTGZGNq+RXmzSRL
mb2EAULWYHUWRInppGyvSYU/Nf8E4qgWi5H8k3TE6ja+dC2mYXCleVE/ZX28j7fa
ysp/5a0ERIjiye9WxTf3Z7XKetSIZTOFOaWBmVwxYlXuOTb5OznnNUHq6mteC8WK
dUvSZhWYZWfbIHqIn8O99EI7NnRHUIuj1nLbcEHChbXhRORCoc4p2p6AzRHXJiLS
s8UIFhTM9q2L3ZDU3R/znMM5Ewp70dEcDFt8NvWmbwW+m9b8JMYAQiC+2OJceDvD
T4achq3IJqglL7xfL5VS1kMvBhp+D20+8jzw+lgBusYcGUyOuUuOk891KhFQsuss
sSK8N+lnXZgfZ7/ETMFhug6XE1Cn3Dd+VHFSWI6nHZZNeZvCaWSO75H1gNjIBuEy
ig4VIcZFQjJTgCVX5kieGLXLQi4ZE7/V66A9LiLJgMNTbvTykJORHwxQqlsehhGE
z/caY4qQAvrAmY7E+aITc+jYHxEfgx5VkifRXXUbQ9AjsspsCRVAzN86KT96pN7Z
HiCSHluh8JWFbhr/G8fmmMIpo8XHwYdMNLG31zEBhvmrizF6pXBbrE+O8R4jfCFB
DawcTcsR18K452JnYKBMovWZ+DR6lXYP64keudaZvprcYoCE8zOMtgFmAv7kpGAO
0BSmoZrkT7RlUtm54l4er5bICdY54jNHawTvEB1HrSZpXKWlqSjRM/XMVv/H4tU7
7QwjKJldDcWYvR0inJ9GEnwYcTZUlPH3r0V6wI/eAdjUPkUrJQ295UMVSISmCB2M
mpLb9xcYTh8FfPUE+jNVJY+W0ZQuQtDvjh+gDNjEhy/oNp3yn2vP1XhKinJQxkpn
a16bOPkPBKpA/9+6nZXTSoNzDo5CHDkUOhJ3sva8s5P8DE0PEsTMwXya1Ria6e7N
Q3C+7lXbc6UNQcsiaTW98mqP2vvNajhGfdKmYTKZl6KLUDjG3vmW073KbCZyXPcr
yQ/7bdBVTN0szDdklBedlapMJhfyfWuM+bjaOSoUys/0HH+XxKK0WLKdxaNnSgmC
8hO4eIAd3qjoi2WqNBwQgHcNPDu2fw1sQNMqctqrpRMpjedzkVgz5E52gZIXh8Bw
BwNNFKWK35dRLRKkN+m/S0Lto1DY6VOlP+sxu+79iWSaJxOUDHc3k67MdRexG7r9
CH8weobmr+NaMuLSvffaELKOBlmv8bsJW7MFUGuI/1DGrRpMjXj5q/Qy/PLzzFJS
dAzRGtZ01aBoAhY9v9PRzSBGXhJuUFGAif5ORVpS3ajCxeUJinAbihgDFLtL4fmR
3gZu7UlsvyssSHa+NZC+435jvJMzGjH3cQ/hQZjfKbjZyiO5TiqEPKKsMyAzD66o
xP+H3hTGHAS73Rg3UDLRsDz3DAVnnyyAbkUFDhYaxIcaubakxW+n3yC8hhlmBGxs
3Fh2qN0CNrQDGrQAVxaibQyTXLi1WZrTTBggJWqJw4dS6YmWJ4VCw+SMLcNNWGeJ
b6hONfhXoKD5HZ/EBx99MN6RZSN6pNcsFZQUSXsOLhQIrbR7LmQo65G914Yc3Who
EeJy9Ckocwj4PfRnsMAq26DPYRxs1s0EvaMhXZ1uMmwAibCprMl55L1DtGGUOos/
SSy3pEOe9y6OioUV75xcBABoDH4ghDueCf5mdU9PQdoqS/uDaM4/Ppeo9GB6/wyw
IeE2Xjwh9Sg3XKJfCyfIshwN0h+6uVmdP1Zq8cITscEm1M6xFXmDO2O3MW6G0XAt
oRJtCrXehulIyhF3trzcOEBzWNBzrGM+oMWOkL8dNlDS7NXxQS9vC3jQcYRsh4wY
xaXIqyZu8uUI+q8fmaIQ2D13M3U+hGP3ewK1QjkZGKoAKJQYniBxMLPMKmwDyLRu
9ipcOzWyy+d9JwV3uoX69iVZRPG8QzHrAqszv2oyVFbkeOLX8WP7rA8KBSpLbkvb
wTSUmV/GOphd8GCbwdzZSkrEjm6Rru09mlbuKWIvuIXigoIc/wKAXZMTjBJ0dT7I
MQUl+imSIFv4H9mcmti3jlZuQPbCvCapPFbz5u6dbmEkShR6pOTWDYagKt1F2Pj4
eJBtc+ILemkT6migm2FZZd1s7maX+rnO356zzJI9vUoV27OxDZ5RGqKBd6TCKMw7
PNrR1cVQaooj7g6+EIzciVNFBL+mjCLmdABM7VsesetLtwJS5RdoQPl0AhhPNr93
EgIuE1Hpy7tJOegPi8AdQ3njmbff61eYXofC4cT4XKUMeI4oRyC7CQDQmbNZPPBG
cYNbrIxkTO4YyqwCIsxaW88Zq0mlAcWFeqwvoSPu/nc2SwEidEQOnmqOyugjomWk
AfVpyYHHUaP5WHxj3Rg6PTSi11XyS6AfqxKix4Yl5m11cf3tQDEzW+XUdnjWC4SO
cPFycgjK0B+2YqlYh58vvlis7WMaVKlpfp+PbHV/KNE0WqCLc/Cv+TWM1QmY8UZI
iiteMDgFh3cikrNta3i7eaH+GCZgEbjto3gaXXDlGy4Eeo/mnCLdSGfCU5j8iyf0
u74xE+k06lVuKOcEESkOOGmMiW6XMsN+EMWgu096ztzxOOAc2thvBLKGHCgINQc/
+r2Ib9NuiCJ9/ycV/kKja/GvkOqQJ0u2lR8Y+xV3iSIbKv6+dnay8xqMv+9JEHp5
Aquc1oX2NGCR70qyOPIkzaLRSfFgsfvX4t0EUVsHWBbm8w7gLs3ZJTErNpoqUmj3
4/aCLbQkripiR1lejQwuSbq3WIsu8FKiqcPKNvy+YTGFKz0uf9T91GxOegqyocfV
uBwz6ulcKcQaqcd7MMu4YmLOnnSnkrzE94F3qtZBEOlFQhznDWi4/rlTMDF+RZ8t
dCJFqn6sbrLlz+SZLQ66y0n4zUisPVoN0AgELuaoYsfmBPBrAlihNY0fD/7HAErR
p1RXPlORUfM82scbFrBLwu4o9N61nUiTTRU98m/LZLEpf9vp3lARkMnh/bVGJfMy
s/H6PlhsgGgvrLKhMB/eGVMMEq8MuNIEt2ZtWVyUAZb8CgfVejBQqM0DAJdXef1s
oQ4qfvZsSYBRGj4CL6fsbK7eMxiq9I6QFvLnIERjj/JDgSvoarUWgH/j450j2ex+
+YqmlwqsZ/cKrbKdKirwqJ90KURitPioYPDdBbOvQSEL9DzsmNMr+cwoS8ZYaUKr
PjTAWKAfxmG6PASfP36O+KSOA1P1eh6xOFpB2Un5XqYYRz1hafjtQ8/P7Ca1mU6f
BdWEEycdpbZgmep4FOl/k08zQpZaZigkj5phUYn1297AhwFKBvS5N2TqppS7rlaN
IkjYWAhULUPOq0w2+QvM/av9o545G+djrxjTXgUY9Wx++fWv05avTf+H04qKUM96
8gOcWMVY6r0DExMZyIpVSXgUzzdHmFjxmB4UIFebJEqPphTteVbYv7M4gWHkZx2n
J4HIdgdO/mMs+H6ByOPwcQtzvLmprvN61/udQHPB+xK6BUEvRZkUGSUcX0dw9XVY
L/PeLZrEl0pygJa7GTigQWNMnJLoojakzJibuExtUjohozdA9ix26dmCmYXeOdQz
QwrAZC3UK8gwoau1J1b0OYpQXQppoIuE1ZyJspg8fP+i3k+xjuaLq/kuh828F3yo
wVGbMVz3LGKCpXO2/ZLkErGaS8MWG5YCvcRP6yuqo5UPEGiaXwDOXj1njpqh5Dbl
8VowGohBc/1Ej9xSGYgEgZB6+aqoyIOnMNSXoPiCWarZwF7HYgi7iTVHSJE4ev5Z
KPvh4yyyCnwE8S6TyrjVjS31YrlosIWzSvUE/5jKDqEy3Dguw7/DCBh3PQxF3NFi
feadnX5JW3F1yyDkRJRQtRPCAq0R+ymjXLEdQDPimqYT70GEnAbHOGxI9yukPrpB
I+Z6pKiegV5xH2KYKKqu9W651ZOnviHCsRi1rRWYpDtbStUVBZmTk9uK9cYwvWXz
UqT8cZkCgUEpcDEEqdVhftMHAYmD4mhNm97aHBus6XoBe8HNezwNTGSozL5co0pG
10lfVqIW22KqSe97CkayVFjpz0u0cGNsLVNJqwTZvhSC81xTczV0lSi0RJLuOJ+w
SIo89lYGC2mgUTbmg1wGYtsukONJYy0X+Awf6ws5kJ+1iTKgRk3NMHgGKas51QHa
gbYkZGuOk8HJW2PbWWr03NYC0ju6c0x0hpj8idpIQgjeZBXsI4lADucNbB7Y226c
QkIFMMfqVf77kmNS5LQbVxk82jx8TGVc1/mKiW8b9/iiw3SJjnYXpFfxN6Zy5nxm
ViOvZfDgM4HTOYZWARnZpheobKAeHnQJF2yXNEvQPekU+fLXoNsaXLXH17LJ95DO
2xUpIMSKFekqEi43GJTiX/mhvHBsb88NgDZSEgV7tqyybDn/R6e3NOep3JcLg32v
v84jeDdVA8dQWW4QbKeJXFa3bMqDF9LMFJnD0w5SbjsdJWXmT/eYmqlJ5nxcl/im
ooA80ZdM8e5j7kTafuEQWitdCT77Cj6XWQ5M/PuISl5Ayo6nt20QvCZu5ueHg5aE
qjBa1ug36eQoRfvLAGvCYnSK1bqqQiPic6Ma1SfwRKnpr37G4J+sqR7HXG4VEPns
EOo1zR/vchqe+43X6/IwCczrCP77ZZVvV8PQzew3eifXhN0DkfylR8iwpTg6Ge6P
uVC7yxa9lElsTlqnv1Lem8JveF+cWZtz+xdceKocemqJX2Vug0ueWhl1RmcBz4C4
XmcHMuXFamtLwhfnUcofm1Sp8QqwnD1ic9n5vQ94UegnIDqP00Zal2OkKIpMRGOj
ej+fllhggcLpDODcIrV69hHH/st5mPflqzb2kry5WdmJUqq4akYtgggK5fUAgFfH
tjoVqtx30SK2LXoPnkejdcgHCVpJyA9jO/jahIt3iuM6KrKzHxjPbKJhBPiN2o74
YIijbmmF68ritJh+wqrXMz2lNeOXZ0CQiFkOqaprD6xUFut58w/UtDMaq5mcLXo+
G+E8Q5lqwoUt2ZRRurWuWM4V5ItNJ1V8PV+m3i9T3E55ll5VD8hGS2yNqOa+cIB/
LCUrMlx2r2l2ULeR6HaDaDen63SZX9YRsqKsI/eGF2txY0/QYWTjSnUYdrnlsCfg
M0ezxfFTzhYyhsjUyOyxVSUVF6WBgxBzQFHIgyj7x3QyDfm+hdmIgUnUbkYF4NiX
g21u1kPMwBc16BqUhA7Ir4fth8oMGEUCeTm4ZUfF3Ui8OPDORQnAGyDLNhcESs+w
1IGkV+opDrVdZ1Qlyde8Ox6i2dU4B360JjbQve6iMU6qXznm7Bvzrf6FxEa6mlO8
8g9r+/fYvgl6c1Gu8XFOYnBIUGMO0tuOwrKOoGHEjvYx64oXzjeJhQOigbEyQmX1
FpRxX8e14s+/Q5tRGzwnEXEyKzzJ9axJ5goslj6i9KRfBvVoXS0uiDdx2Kvk4pD+
9Ji0jLcT2gV/fS1BUgyAKwRFKs6nOSVeAWOCkVecpGiv/oQcoCeNm+sJ1HiPwlC1
ZqYPo/BgewhayeLdArUc6PPLrrpf+cPzv8QULjo3X26bMdS3wVHUfdtmNnkbgWy3
LvLxZKkXV6+nvXe/ZB1HS6781/P0j/HEpBQHToqPKeYQINwftKi8B0UEKWczVc8L
vMmVPmwc3EaimihKEJroGkcYowpfFhYLVpUQ8EycYLow7Sh/nshPSD/XnO6SLppS
kd1RBYWd5/rQazHikyu87XSrpmOoLW1+Qjo2l0ik2T3UPZljEFMAZelqIoCcMxwF
cOQn9UDeOLEwIpfdR6d2xrkGrK9/3zG8zvoJFXCxifvEweJVFYD5qZMKGmRxpzDV
cman9OunoThLGHFgyv3e4eHtifozxdK4154Lg00XY1mbsTmogwqUmId8NNCWlzLn
rDaZen8UtkTEDJLBrzflsiNGWP11sqYjh6T/PpGuIIALnmI/br6EgjKbQDNQQ2uf
RrxS1PvfWcrz/FWndKTPKCd4svm+dSTNYVJ1gLq4vtsgwF83X+Z8mdfzpo20oJ7D
vbh+0V6Tbxls9VAXh2WIo1gs8iDFx8DVAp5a4v+QpTdx4E+frSkVuVkyEu/Hlqge
khdC90XLbLPBCPkiYCAG83/bHHcUb4H3rP8GdPe/RKSnZucoLN3fyNmZoaH9/XR6
TOiMwZ1FJZRV3YHcYL2nKAHJayvwWDdloglRutuA2yGWAbzRl+5V/m1/s9/iTxhg
JhBagGPtM7yQEapljQfLBuuHXX+AR1JzER8KqBQQCEyMf59yZwLUnyccH+dk5CS1
ZyONohymAvb5j9EGDM1/XPmAKxelgoFVB431ojT+0hwGTZkBunOJtvRhKKtyWXCY
huHfvcLq5o7pmoL91gF9RwuAASA9dX1/gg2txkNu+Dhxhq4/vrfXG5YLmAq7E6q1
qDRIH1h2wFaA6HoWgkVbb/T0XBLVr1/6eq25d01A6eSaCnPKj6GeVi5DuUQGxbur
fUbvjtVPpadrX0v/ATo8pSXuzHly03gkRiZI/6dcsa7IB3PAlA+Dy0xt2kcOmmyb
O3VnCmc/0qwShaDX1XFQNIYIxDlFmultKlb5zx4E/L/Lm82M/z9W8DoBPsVk+4oZ
owYA7hukS8iJlpxhxxWTJgrDUMT3KiJrPvMWFHQ2t3XhnHJS+d3ulUmnGKiw9R+5
dRk8H1DvWa3CO3BRWun8dpBa8sfR01UPsprc9KfhxwUes2t9PCRcBpuv/7n+Cj2r
QgKEGpKF0qagaIm4Icav17I2zjm/fOU9BpTd7nam2nMNNUXKvuzg9tWhhhJcxjsO
PotAZr3YeWlDKHeQg90pwfItfeyChwuCQ/2GG2ZtQk3vhrvrDmUDn8Q44BZDy1cG
j4d+71cS3JgYvIidkGdAtGZAbz0Hl0A9AWK6sAZukhwKZf3wYDIqj2lejTVXQP5d
0dqDSNPSRbGyt1LLxYsKBpG+PMGxGdwC8nGGvCRTVVWTIpnMjBKh/F+QIA1WrT5T
s7/2eLxhwkqtQzZimf+n79FkNnWd2U2tUHBKyr3BTbVsP0h+4kQQgWgMtH2OxsDS
9W0xJcq3kwa+n2Vub3GsKxMAeR/mMPhe2JiaDhsoyYJCrq4bIAwDDfV/6Kh7cuMg
/sKncJoI451GRTJoTJ2EhVieyPAPvYDmta8DccydP1iwGgX503beOlfQoqJ+qjcG
OrZBxJrRihELxwse/+NrvDINe9iIzvUm4+AEcnzZy6/Jvn7QURVlcFoJz5hsyCUj
MwjExW1KtxH+IYCX1L1yUdDsFg9Ldy65EDpi7hgtPtWgbpCXJUZar8s8cttn9y8R
Fc7RJ4AgCAdNIiNTgxxKwJNq7YFmRfNE9xlelEQmShIaSMUWbzyVcdAfph/gOn1P
teXQdZ/kbUdcFoB0CyHInAOSxznr8ewvv3rQHwFZa08f+tkpGWgBXrGoJGAPuQjn
+ZxBfhPQhqqJaRVG+noqxmtT0R5H/pmqBcUUOTL4HKUgBnqNKKmm7YFWM+8BKKgZ
Ii5C+E2yZI5U2ddEEVo6XimyuKfZch4DHtoLGVgtfhkGfp+XnhqFVrr4ANxNvtEn
WnLZdWfAF1csm3GmmowkSO4fHM/WAtPAJzbDrYh7gU9H8IWH+LqGwgA2pzZWvFDf
EzWqicRuheskWZZQ70VnnVTR6LjL+zm7jF6tR5fsycdlQYWnQs6j8siXFZUunuKQ
tGIS0gAdJE1YfdyuLfkeYqf37i8jHchEa15RjtfabCS4drvZSDSbtwN9IESxoaAL
dPBOoDv8dvsmQ2YNeveR0pjSGbzjTHZHvm6CXsIEjKIe2yjjkShSm6glLaDsDgDn
rhc11AycbPJxiCoNKhS3HXm8WBAvrTyTCVMQTGq4iL6BMVjoKL1W/g5rS3VM1X+T
hDjTOXGarOBzMPTnNz7sSlyMWj/VjS0eTVUAIuCEK7UJ8QBYOmHup3hDoV1dLYZ9
tDK9urm7qLHmXP0nCOBWECrYzjergmNE06yqMMnXbdul0b7LTVBcK6ntuZnAfnew
ACut2mU18EDNRUCotpdBdWs32o2fdCt9rcvaR+tgu40FoTAM86CgBIJc+9ouMBLu
VIvsHyHB1vW5c2P4HhpW5bx4wjGZQrubVAcCUBZtgdbBwwM02HalfXFeXM2SkmE+
ArRIp180nY4EAtnthxJNGNbofOJCrWr82Vo1z/z+n/59e9wTR+ANPmIhFY2idsXt
HbiKKfa9ZuvmhYkoGzLJDaEZOrMjRoS2uYjweiZ/7qDAjNwSi/LcDpJknwT1jdFn
i5kAjb60GsDIIcjh2H/kXCO1nMR9u1Dtt/4n3RcmmlfS2ZIr9JAwiwJq9R9nCTL1
DWNpAXcfZom7L1QWWe/f+a6kIBOvYJppVsIEI3CuNZE+J0ua1VR5eN6KzqNvEpLN
1IWxZJF8Zt3MsRC9WSLrNVAmwdSna/O7eJ6ABwI8QnLwoOVp8DwT9pPAAJJd8lbi
Ny59+Mpci9e4e3rMOG+5hsb4T/EWyNkSI6hyRabS9NRwVqwKVGjS3Etie+oJOsiv
TV0/XZJDoNhHzDc9oGw8MvJEV3VuS67q6ayAQLZKTEd1KTdxFxJ0dcChKEZ3DGx9
UlsKXSWTSrqQveRpArxrofm8AwPZDuZyNEOl7/mCixlL4+QUrm23TyPB9npjc5lt
eOfUQe4nqEmjmnFZWzMI9Jim7JrOZXvRqircyVYz8NxfAu8NaCWLy+J3K6sM/j85
cKl+44tKF3tkLKjy4fyzDzYD1TY2k+bHp2EpfnQ17O99txMJ5TeDuY8e4GKuUoTG
CDEYW5fEJyvKTyWUT3A46xZkvrk+IfuaTRHcIpxg2Ctho67my0OKXp8B5EtSKwU2
PCGePyKi5ZhaYF9312ioLQE3LwGn51mLQ6Xq2wM28gE0mtufVSH+vS7ItFHhLo0n
5QYwkwhCWTrRGCUUwmDnAKjbPO7oCqMiELnZTMVwEonNKzLEwnNC8b9rZogOTSrJ
dwJT8SxpRCpkEW80eoTjnPbpFYoG4NfpSSgDO86JehbEa02+LfRn3kVkdMRzo0KV
qVlcXEJEzsMeR1A3khJqUL8nw/h18Alz5XtvVp9EbZJu+PmaVdOj6AoeDV8dHnPY
0Rlltd+kDzuFOBJDQpeobD2H2IdE4E83p3dp5vhOFW1fkMWNn1C17nytq0CID0um
E9Q0BHiVJFw1LXJ7KwZ6LAgv814xdnsV20LDveTRozYLfXhf5yV/yPVdkeC9YJpU
5bmO7z/0rokRh6SHQMH0VMTh4/ZE5xz/NgDpn0V6zxbF+Ox/9zDjMvwL3stlHF31
XiqkP3bSd543M/J4igCUTYGme96zuJc++2f5f8KUH32fnas2FKkeeOf68iWgvbqk
0DBpgPWaarNx1gN4L9hKrCSbvHakkwkAsDA7eHrXoXRxntCP72gplFxnbEpTkV/s
DMHXfJhk95Ofs6aWaViyXAc9+9IuCsIZBXfd5CveUkQRgUa4tmp/xdpuQiUHD+6w
ozUu1EXmwHQpcJW6JiImPKem/n3lT/u+DSnHhUs8UALwOKgtYyrKns03i38PJPg1
4DKM+cOuX7hdVeQbYkyg2TRg0EOb1gX5zY2BVC2EZ+0xXeZ8sUiuqWkQmqJuRlwq
2OllaoRglg9btX8lkL6W2nkp2WfgHTlncbMKm0i88/bHRCToU0C2q3cEzEr8PtJu
0OJgZ1Jucm1ofthxkkZaxoRogBlwEV8LstKm3dVOvcdm3E1sGW/NRfYBuqWthD/X
0glQmkD/cEshBGTa/9TLV22F4i/Ms3inCGtZPHLI3GZzMAooFYqhL4ucFwARjWDX
g/NhXZWs4eWylGdBCNTECHi7OcO8XfNS9kqhgwgc4pUCQJlTzVUZIxUJ0aOPPGHq
dyfsJC32WxmjVl8coa0NW+kVCmH1ojekZnic/cSbEmfYE9pe0yOJcxmEEacp1q22
i5Gu6agsmU17MEdA/ob2twiMnjYFomoB7c8aFmNg1RogVHZO5oOXlkSyhjyB3tix
vuswA9xXYfuCBVWxiXu9/3FBO4HV2LvNRYmNo+7AskNSDXhazkZzWr3dGWu9rAJw
GjAo/CONWcWqU/EJsUxx2rBV8MLDVdpWKPrkScVSdfFPYnDy1bt8j5z+lscUrRie
/OP8wZ2RNtKhgeSN3n/dgRdhMiWcBXEMqyuo8soreAKR0Tr/ZCpZ183D62+/ILsQ
2o55z2EJZjttEVG3IYkLtJC+uyGSKHymQ14vgSgB+emBJkzEo3mawCrFJcAFnY4a
bheLubMlB+tI/+QgkIv8rt57c3gCqu3GmBmGsSy7EBRVPsr9QRZMWC9x0xArTm8d
VK7t/bFcRqOKettOzykLlr3ndSMqCXUuytCw6egPLrZPszIlGzdZCt08e7fTgfSS
roAQXVYstS7BZnxVv5nkvtsJ2XvanUOiWsZ1ECtSb/+11Q3hBmP0Hz0OFZfmdEHF
Flkm3S9B9FlruhDNu+g8OeXoDRdqRx9uk1gUYV39QS1qT4gzCR1ykIac1e+dvxf1
FNnqIgc63FwRmtYnwmCVtLw8nvwj5Dk7azR1AQpX7GWeAd7cqV9PWu8feSfpp4nq
hlo6IKstX45k7Reb8cQG8UazHqgjSPjxYgvF1hteRMD2TdIXAWcY2Q9f03/+YYtd
b7T51nfm021z20TY2Y2CNx49Yb/21gdCnQ7yiESPBTgOAaDU5bOoXbzyNK0l+262
ZEKVi8XYMeB7QV6dxmul6ti+799SKUItJCpCumQKTYpTUGZxGBXvLPcKwNj7Zb58
8MEr16S40vX6pFe/Ia2yPGBoX4+fRMwB9vFAOl5F4wL5e1Ja3UaSZzXPyaLOOvop
v3tMxlvFdHDLAWGCsubQj/r5BBz594bCSf6bPCoL9YasFpvwsjfYwe2H75dH5BdI
vZRktRYauXgwe4FE3wALVtHNHk21Cj0g1fZbKMxuhj/R5uRK3W6wpzLQKFcNZ+A5
b+2EnYkYA7Hua6z3A1mgsUKY/MMCFq0/SCpeH4KnIESvOpqzb1wsC9hHOeVXsoB0
3isvb/hvfqs/1nbYYq2xW6AW+HOLJUMKRuPpfMV1nkZP8oHUgWMgWGhNpvbprszV
gaOOqV6lM4vpPVtbJ6p9+lHdkPIPzHsNxklZ8xmuLUMjgVMrvIsb39vxMRNYMLFA
MgpEgzCJrnFwzXapiMa6CHS/NE4iIJoSQmZlOlm0P3iuED7Xd+UJrCCk3ROK7rFB
BMhOrUsFvi62IrqZWr1tO7quhD79VnRz+/PcyD0i3SGusips8t3MKAxY0B/8dl3b
UELkOmaFCgMSq0gcdC/8p7eQEXlMgHs/HdWui1Dw9eHmGY+6G3oRTaY//6BPv3gr
z3HGhktBnUkg9pPEqNzEWf46sL4d6RzxCKvR1SKcBbsFKxfxrcZ71AEXdF8PuiiA
2s4+5bBcOYyQu0nYUJCg6Uy4Y0NoXG87VV26DcpWsH4IEpNGRgkcPUV08cp0xGoM
xHbZeYWhPwHFTmK7LcKTAUS8BiMAchn7K79wrtgoYWgv7HppZ0fbmq/gRMRgeGyL
l1jTS9WLsgAnWhCHiSL5wDaf/6x2zRoYKkCCnl80Q8Wi0rAayYU4LgXR6sayR40X
7p+DYYYBuD0Lri1wCPMqtmTtp7XPGqdnDhATkBhZHr8ORHXhVZNORiT5Jo8dE6o/
7Q4BYxWyl8TmYPgpczgIDi1qSn2MzdDIE6x3U/U30+ND77AYQjgl39PgkVyJdfHl
uMirsBBaQ5z8KS9IyezdEGiXnqZywwajWOfcYx/gRHE8aRA7x+otsvu+KgUKBUj1
Cdb2cvM3vIc9qJnJ+SHX78AoGWcD72HBD1YPLHZLXwfn67nn4kFMORtgmYvDClYa
eFte4aZZ26Si1W8AXlCayd95tzLIoGgA3nEVLqF7v2UaIEELsODgb4uBgT8Rea4M
WWog89sO+mW2yrV4fkMzLiEUFMvsFNIbTGsSflayJ94/GjK0eOQQhYQztW+tuHgR
Xh3oX4AgAAvcFFPAj83+/zLmvtTrkcwxKFdxOqqKPqWL88ouPb13VfFs1SRLYitt
5vULdqTean9PdNQ3w6RpQ9FIfRk295MFgSl51ddLMr7GnAGjfXmcWNgRgz3MY5mV
S0/kIKMR1R2QW8xidIn1yAWw1ORfvg1X1dUEfHvKHirxOsCSUm49PaOIojBjk00q
qbsYbXUZPAMH3x+WTEFg3wrz7q4qmR0vGEnFuX1L8EpXZ4EB44SdRikANkLJAuzw
CGbtvszPts/H/V7ArJyeDtAcCIBL1ISlLMiAYBezvC7kiB4mSk/MPPeAVEca/KAo
NHRP2EWXSCl+h2HQBmB5mCU2RHJok9EK8y9yD5LzPe8dQQuOMZ2NaNArU4L2s7Zg
cB8xl01c3IPQ4GEwlews92oLSW8ShUWSUQ5tKoPBHmp+9Zeb6KFP/RpgB/JjOxJQ
jf/3TKZ8Oa3QwW9krSJHAJvh0DqCjeCGdtepn2+wwFA+ZS+Zv/WL339karTqk9U6
OyxuPlzvCAO6vLoj1pR94FoZu3Ua4BoHqiIm7GO8iYj4jmHhm+SW0SDY+2u9EofD
KWQv9+uHbRyPEFiQ/2rpbBKLpEG92P4txQB08W5XrhugmUjUKcN2/NpVIGJGyNHQ
J1h/svWbJ/bmQ6XMP39XWXJ7n2nJf064r18KI2DXqJV2E17RiSzYSmkUO5zU3Vv0
fsPj7IWOQWjTjC9xeLK3nWtNfIkHYhMsT6/lJeVzxACrUJ9kx1Msso7f+XFcqCCY
mp2q8Y1yACoC4wmc+dRiM0MIWtq9D8G28s2pmrVeE0rV0aXuXw5dpRmVHzjgErEc
a1jDQytsToH1IOdY94O9abVt9NfszETsbyAAcEs7XwZLUezdphH3i0waGkB2cyLO
9iALNOzfElJigoZNr2iAqqjU3tSi+Tdh5Y4wqMpMiwGz9EduhJuCsY9egqkVthGx
jX3Vq040bBWAaBlE3IgtAbzp8pZZygvelm+LSkTqlxLB+oJU8tcKu9Vbe7qy0o4y
/SMXsSKbqkIzncJfD0wx8cvH4a/1D5KUjMqwlOEywdqS7Jj226bdJ7YuEjpLRHcA
mH7Dy4PFFeKb8mNXQkE4d9abNLXu2NRFHLxgUxFJ4XvKARNa7ddbjBiDDgqrpht1
foX7m4VLnxTIkOaLEqZU6zY2Hos6OXf7C2zXphUWGh4N1zb5B7jKAqBnwpiq1Dbt
/U+DJnJ+MbYQNbgOY/rtEjZPwqXabp4RDdVI9yfMFWgMO/IOMYiZ6acDt4YnFy3P
nHGwurBvCvJoRPCZBUyD0AK6maKceh62SfH7z+1tD1w6NgGsT08kF8Cxv9Iq15cs
erA4s0b6d7gUoTx8V7eVCnFPfPBg/RXHG04CAjRD6cQmiA5hOiYUOwBDN8+MItqG
kks/vSNNRg8vPI3KjNGtUhwGNktB4adzU4UkvJQad18dsl4yF97fxC6USiZTlniP
l6bt4o50G7dSh8y/21nsYgtHR3p6zd3rdQ0T7PXCGISAO+bv7EwqrVsl5PBPldcP
XsSYhwjq30tY7id02bUhdlzgLKecuSNIxrSUiP2S6QXC4uUqNpyLu/KTzCQnPfZs
vchm5Wp0p4Pdo3OZKtmSZYKDIjecOyMDTgkHD4xUr25wC+Nu0Ki07RzPk85dQ2ti
ETUbqdqz3OpY/wL9vdpOl+SIU2zdjtO2kbGhNM16PGtr33LAa1h5jL8LcSZqTo9a
jvWGghTSvap/WizoV3bl0qCzSC5sDnl8ee9tgwjBZWNyZtO4Vj0YzjR7JBbIhPbJ
nQsOLu7AAHwIZwoaIvqhiN5gFLIAVtwxdKLgKlst2vfbF0N5iqiBz1bSEPfVWPxi
j13HuFyXLUkY3Lk3NVTfZ7sfWiW+OwzdWntPY/6JOOhuoiDxZoheDScWdNmYmi4+
Q6PTqmNRNQ96P2s6JbxFwWh+ReGkKGZr+qiZ+Tm3d1Uo0P11Ru2u1AXC/xFnJx0r
ROUGq1c9pGXY7fZsJEL/G7AriBjdLxynMFYW1oYF/BWPcnm8b4RXkDm8jsBoAeb6
Am0J/nqgLUIiWqwB3anT2Ndu8JxscGhl2v6p9S4fX4QKG3hfi+tlvEdQ1tMhfpRH
AH7S+1nghQLAT5cEaWOhmZ8gKQOWCl/b2dCnWWtuInkthL6DAagPTAPee/ji4F9U
Jm6UjbTEC/i5lA9TcN3hz6YEwIOFNM1ZO5K4Zcmcetg1j9qCleBfX9h9IW4Ktf/J
TANmwNNgXnTcRqNesrKd+zMx7K0bvQZQL6E0RHkdA1/15xt1nwxDuvuQM+6wRifP
aI7F/JCUoXwK0mNpN8UjQtRoZdeFJwtNs+s0ncAYyFliKGqr320nM5kMYLDZaGRi
kOdkj0bub8cBPuXsRAZyKTLEn3uQjmQrvUqczhoPyCFWwGP8v8FuKn+e+D0nDzUB
oX75UJSRq7v1Ur37XBQm5+V+0/7yC30qZuQBYoBO5fjCJ631h84sA4q6f4GwBJDu
1keOR4GKC+Jvd1Q0gNBvkl/axxu23Owee6VH1wEu9eTZathOjWXDw79COEFekBaT
0MJnHoTpHXfJpVxDlI7u/ho7L7qF4fPugh7wggWy/h8gSZcVdkMf4qBoJkBJ5JK/
hvuTNZhLhPSSP7t+WVAgLAh7BLsmiIS68BgZHOl37cILoxr3yuMN6Gro+IHRjWWD
fInD+CxSXQsR3NRPq6Tg2VoHwLPHEibzW9HSMsXGFephEHNzDppHMEcUfwGOs9h0
HIntAscq2oZIx/77m2OhHkVxL/MKNxkyIjogenoVXG9gFxIdqAzCaYK7oOlv/17Q
dFitK0LxKPbGeVUEDlZWZe3+Yj/LbmfeEjpMUXRSX8LqwHQG7Ztwvcxrj0MRhJSa
X8oxfIIhznjN3sCOj+9Fm+UVi054YzJ+64ccI7hlwePhGfvOs4Jm1jspSZUOwLpW
TsYiNJIPpPbd1joYDTgZYl0RfnkFsK9Le6/ZU4fxqNPzdcu7CZjTFoDLex0UVCzn
Y2Sn/qFTrraOyrJJ/sCkAVFlz/lyYEPBV/zS0pKWofT6z+Nc9YmmZmYVgzXpz3Em
EaLc3jn/Zk1Ol5veURSyeVgkBVBwrcDUtjxDAXPhfzsg4CSiyn2Qrqw+4jUwtF2b
5MDYBHlhmdvbbjoI9Fz3vjVOI/Qd49upFFarLfiEY/AAn+/p04s8gHwWwY89Kdj/
X9wZQEumBwYLzWztVjoycr8BYapvhosar0GP0ctLqh8ojR20Aj82QmULMum/8Z/n
xXDXBnsK3crTQudbQFG+f9EE60o7xv3zQjhDzurOTB7D6pCbIEZr9WoUlq0SVuj+
cTN55uh66NAcuM8PzUcuUJfX663SxzT8kf+eyKnqjb/aWh40y3gEBXuIcf2/FvKs
5cv9aw4GKysfO7XSJts5GFxAUfvt+uZ8X4bkuX/QamnE5L881cAtPz7d7i6CoIx9
BbLhrRHip+opFGeAhRwxFXXvJNvIUql4J49hQXFLmrQnTEzH1cDcegZq8RXa+ZE4
fUCzBoNfdg1F2pWLIr4dJ5ogXPoFu7rywpP5ysahs6hPsemq77boGASiRFfHD2Vx
+31wucvbASVKwftpUJYo3DURDTgeBLgsqX+pnZ8rXg1u1BbLSMA/P0qHo+VpILZR
aeJjzIh8yE/LQXrOYW9ucKoVqlIlYAHEnFH1HrsVdn1DiPh8SPulBfQMJEp9dyzH
OBrNgO6mP1ISyuUQNwohBz1EHDDhWnoo3SA+AsQU0ulNgfHsWaBFp5k2BZ0XEvV4
fXX4psPGQ/6y3SShvln4/IqGFnTm7eq79SbPxurpJlu++V0sNSE3mtCvinHlRMNk
3uHBdaDpQrin9/J6M+w2TV9o2eZfR52/xXHH7L+iJT9r6eRwPHFpjokw0JNoFkFD
/ZXCxm6QIfl2fN5SjIl1lsRi1S8+csCXNRwN6sptMpd62ixGpjNPzVfYqqXvIkD1
sVL6FNfpVh2ZBhlfK3U91BJ4LLFa6cgwed3SX2A3CaUQJcOpEJWly2P3242NtgxY
3JKgAFf1RSR8HO0ATPplzxNcf9zsjAGc+z04nmIVDJqMHI1rBFAMEyTtyMfFYpyL
kPgATI5ZG9VFEYZeiyGa4i1sl2Wuvk4N3m6u4WCeVlLpiGtPrgztxsqDsRGnIGNF
+FYiyYAYL5ARMHS5YuwQBvm5MHsX2UETeVd1JtPfocs96liHAPxzG8zGIVL+fUG/
lw4sBtV5+YBRRNSsqBcna8zEUJYt4NMV3WB7gOqJXcJPQBLPPIhct7C7FI4nO8m6
oMKfim0pdBvBSuwZrDMzyUM8j7bUgOksrD8httBbGiacGZXwCAwS3+i4zMeOQcd+
jgG6Qi/HeS8/7boxrNogaKu5cpq+zPvtHLvHy+WzkieQoc2Iith9iUtnd+RtjSoV
7kayAWQZDOlCPs67deopiZuTQnUbZTqQqeRFDYk9A1nW/ziL/RHdPlmNvLlUcaYY
KQTUgJzn4xFCZH2PkZKWYoAo3dvV9CjZhJO03z1YVcBAuCqpMH62V0/E7SNsnLvR
eE/8s8A1LqMtyuucShBE7GQDUeai4gMWKSZ9+4UhVvyYhUFirSEp40uE/cLwf9Y1
SmDIeJ6R/kyrMAwxR8HtOwk/MDGRongwBEovAB4mJgduQcuHfEER/RxvH4bVpiEj
abLYKsk4V/RMz8NMa058UifyaLuK9BaoSSYHiO88c7ZyWTjXl2kjDp57D71JnZDg
gLYlP0skwr8JER3SZ+24rW5qJ6UgSIZ9SSDI45c+AqnZwbsqnOVfrfayG0LdMVyo
OywDyMMZoe/UZBxFa4FSWExRdLvWxH16bVynjngeeog6es9xGjjcWOxArdmc8Wx0
EGcsf2eRhMt9Ah5F+suB8oc7Vry8cNNkTil2sdzZovC+RGXiFoFVtMOYB0zltAdm
tyz1h+l6ztko2kD3Yg8CZHVKiL65miByV2h8XLDknLFjy2ESdq3OffES+12ZGj3Z
dvEhjvdkRJ3rVXy1UiLsdrFzMBYT3FTWtOIeRHN0SY0plYEbetEBihQWfHaLUhrF
DrH/JglPMu4vje3wqDhPOM85FCzjck/x0dbmWl7cbma7rHW/BC3HKQPZvBQcnt6D
yryHKc5pUc2/2jxBQqRzQbu6t6uy0Rey+/GLGw0m6bXvkyf1i5zf3AQ9Si7YyQAz
6Rr8YF+hl2SMYF++3w+A7qewY+glr/kZZ1UmOTHKJnqqW7u370wW2zGENREDbotQ
KJMzE16w1GV56j+X99FFQIogs/OAwgiMCvtf/123tUOVbmLJOYO3k7ZuFyS2Sjru
cFl8KAKxzA3sUvLXURVDx4W59df8Ft7Qqhw8V6fP9lJieIlHjoxhdw08P35hGpGI
174WmiievF7O0o5oZyPYBXH8Jl2jlGF3owzPzawBMBmwyjAVmUC97fztP32WBt6W
xT5gk/MCEHB5n+RXY57Yl55RC+ri1kqHBQD5jeI03B+hGH6MJP9JN+cw7b/nx3hh
6qbw813swLIe5NIZt2gdW0khgdG31HUBpREu/NZTugpZKY2W2zLGirViM3pG/UFr
34aF2t3tTZ/89ed4EB0NTSGUDS9mUmw5QuuRPinlskFnjdSqJs+wnedIxQhFIt0m
2z2TjzPcTCcUyGKuWoGrhaJfRuxz4o8DFK+oWgM4pg07WSRvgPtmJbp78poM/uL5
EkSNXOJjrYzHKBM4nENhYsKuly3LYUNaSNRnJ9CNylIPtHLDvydH8N8cDzWi6J+r
tXfJ4VYiaOVZ0Yc05ol/IzxkJWSkg7J4rYWP2TOU76QFN0wZWpzGBsc7ROqjBtBr
a36QRQdukhPIk4pUZ6YdhAgadZ+zO6efZFI151U9O1ZLoavVT1sdc13q84VcIar1
0bPReQS9kcZFe5Ot8FgdsLtb0hyHiJ4Ok7P8jVX1XrmgcY+06wOVsNTRHOrU1y2A
J12AuwxwFPIzF9OcuQBgtnSG8qf7I5W7UhAZYigzjr0nhNXe9As6GjNmjLKRENvz
C5wJazIokpKQ8idOpdMAQevoelnpU+vD483p/T+4je+ArjV55Y+Z+ujG0Cs9H1mb
CYpKo5H0dGS3Stbcm8M7Drrb0AgDLzGIHuJ3sClnZ9qAJ6gKOzonS0XOEfyV7OUc
ovJErVTeCv9En9+epINAlDYk4Hso2PsiyHrt5vn5Ld/mLAYUD+VxixeIKR52WmUB
m3iEgt+ym3C5y8aB+UiaXe+73gsP8DcbxrIDAuMeKNgyKKYDm3eu+LqUjmdQXrlQ
cRt54rgU/AvEfYUj6iAj/NRNv8PJqSARpH9rcGuljDKILmhIAfYeKtsxbEciigkj
BNOKfnCta51XlaxwlKI43oX2kaV4y6S0BeHEAkn0T6SBYOQra9RaBQQ7Q6WyY192
r1ZlMrzJQ2g2oFcDJ61jWEV1FKmZzjy9unjIljDxHrcpGqGTgptAxYfAi+fBk5yN
bw/QpFHcmqHj6VT3cf8VBLaOaJ80wtnZC/xR62oQNgZuZcqtrvlFMY9VwN7j+ZrP
c6YVwcLKg99pYIhYd4fqXohdsftmh4zfCrOTiVtsZN7y6ZsRalvD1a0K6fWUSdX9
YMVU43XO5/pkFsInH+/B+vlHsoO08kubiJw4t48L8KXtCARUgYpEkHpGgv/o1rqy
UpkhoRW2Jkus9DJxAh9jcwgtaWXhCMctNTc6dOtLUGHrNz4Jba5VvBCUyFSm/6iz
KdiItEYwYMSaF0vQ7dhkP/+NFT45I2exzGfmq3uKAr0DQ2cnJnEa6/em7pJbNmVJ
RNOjXSANuByqNmBEBgpTbt4vdv6ttmR9AphxwVlS6rBu02qC3LQCQJPq9Ow+OPUi
tylc5gQsqDYmav9XXIgMBauzEAQJYBKDPUs2gKSJxysapWICUVmdn17GOnge7HVw
VI7XvFipJfJdFVWEmzllNNWAjhm7typsk4uwuo9StApa+9HgNc303HNEBPTZSOK6
woZRMfOqYaApHCjapMj7VqmQGrdgbbCDtVvzpK6yyhlleYWcQnCCCDTdhOOrkgUl
7HGJrtWE1MgxFHqY2kLtJAkW+zmtPdsAMei1rocmOosNVK1jkevC0oSt8TfAbsRi
bmFWxjRj+UkajSE4Zob8HgbCdmd/nD732/3DuKbmT0VwsJ4ziUJzVaDzx3bP7DZT
QbRrhRUfQm9VeTg1FgVcybmXea66b0jKsAFP5ii3mHnQmunnT+6bQrPYoFPKWwUX
hIb7kE4vKcaRYhTTXCsc7Gnpz88SaGAU1GDQVgxc8aVH0ZuMDTYRygoWBWnWXHjw
NXTIPbl8cIBN8PVDqcddFrxYwNc4wdAFJKSKTchMaH6WVn0RLBbhWIjsYmT1K38G
tWRDkPSowBI8qTs1A9HVRT+jWl8KQnZAZ9hyY5hLX8nkfSGhgQ8J7yYZ5mfTJMRz
LFFlSB5q7d7MRF2i8f14ayIT74lGB0wCMU5hoVPx0B7cAlDGCtEzCNnE6PTZUYSv
CNNU9hEl9E7pIik0xWMWUSRjwJ1/Tyt+j6d9ZUOOFceMAsqyCrah17QDPBznexcP
KSmSOW3Z0zzFoVkdJHArVfbR8yNgFbqtkjpOkBfg62M7XLWYmUbeeBAbzgSKHNea
DDEeZrA9vbp8bxcTDvRqkljKAhCoSh/3VFLSCZSc5J3LyZxfdmRF+fJnYpnbULEh
GcW89LpzK/tyTw6UhFaj7BeSqXMGS7e1N/9aVdGCpucq8ashaCmeroTSVekh63Wl
Ya4o7ZFVAk33hCkcWKYPLEeA2Qag2zq11vXtYnCN+qgTCf7lcoNYVsI8cf4rKN8x
m071io7Xhy44oC4kAz/riGuE4pEX+imsnt4xEPTlA/EzrQsR1xVZx48WKGd0LZim
N0+KTeD9u3wr44GfUqOC6Mh6qMUZb6pQbS62wwD7eC3i5CHxxqtVbDKX88/a+xBN
KtZ0Ozpki6EvFDzLyyKxg2P81sC7+z2bepwJXs0po4OI+wZ66mN4J1QLkyCb8w77
MreQ/4AYvjGWq87clsV/lDF6ik5o9/NVp2eImMHjfmL+zPgdUK4luVxsN5E4/hFo
8OS3m4cPf8Xkt+dVwJAgtwANX/7u23z+LnpSpkj6H7jSwn28lCia0A3WT0lJCnjm
BLAQvqp/xwbp8aTjB3xlBgf/SIwUepd1Z/F7m+IuXMTj19VC84VOaG9o/vOp2upK
ATvC6s/1JDLLriPP9lzErEJKPCdM1d056E7KtxDO32cZL5GZS0G/FbQKzwWua14d
X7lD6N8yYUWVOE9lPXfu6F+i90mPUSmW9bm1C3W4LvbdQ5LnuAAFZNl+V8F53uFc
7WGdAVMYjcxunmBS75OXH6pTnT1EdRoJm34gV0RPvm2g6nZcqnUW6491kHlDOiT6
B2mwgO4nrJG/bhMY6yNP3rUZEn6VzkfNED/QH8FZq7zyKs7C5k4eqEeu4bj2GwkO
S6ondMJgWXZBZ2iX6M8iXeH5A8ucVGgrm/GrgaJrLVedRZH34uBZS7+7rVlnosKB
gbSQON4cDT+Fb2HaL7vgsXxzCcRnginbSz8MEnxW1PO6p+MlJbECVtewU6yLcz4q
fdD/NTzDW27yo1Y2P8RmDhjS2LPChvx0PsUNdIxaupLLC67UQCMa4LdeB+S2f2T9
IQJt0TYB1rj3qQNRUgA2/XJ5QNQPqxjYo3YiLIcW8SmOEYquGoHWnF5dP4GwKuhm
gA9wxXS7/AP7WZfBW/R1RYJ1AE1J7K2f23LedZfS4e8BSz+/YVX9fGzIYJGKX1hO
zi1/PqzCrzomoZyxWXOHh0oK0kALP0Lk697yZTY02Lybd7ocwQ0CKp2j4yQwT72W
V+EpWC3khEhJXxqMw3K1b6KiuCDfF6Bc4w8LBw9NQsqdp1mNF/wybdSYO9KVgaLH
L9h4wpH0SzfJXW4HRGcysMfmorJ7tGIwKx8gTktoJxwj6PCmRKfCqQweOXyDbero
PAziB9W4Ssb04N8JE7x3lcVqIkXlmgBUdzbzUP+CA+9DO9jbrrIQtc/Oz4tanxjk
8I0Beo3xwjPVHKLvZlpdtb2VH6QCxyN42FdhzdsdRkR+9YOllsZasbMpTeHXQKyH
1FRmoSbVF/H2bVj3qkHPKAxmSCymEUXnQGD0FKq10I2wkN8QeE3l0Wc7SyhzUZvG
93xn9OYdmfgSkYnGijdxAOgMrA0zt8Sk9ufN98hiKbRY+o6ZR1osbOGFctjjpqU1
zVG7C/e+6zfv7fYGDGG2RseCo9bTjzCItQSbf7T0ZY21+cpxgkEzfrBq5fz6M75N
GjLCxKzeqiOPTwFdC+8T1X/Gzns7YOtUkK3gUANAbshpc2JlMX13eq+j/r0FU1lM
qyOoXJD3VNKtAwBDToICEVg9jOwV709kkp8p6AWHVdYEjw5M8omWSH83kmqbiRc4
m4WwZ5Az5Dd4LQxsJxndh/LHdBX777RjjhOQwJQfUQBV957qYA50hBxr3v9XFp/Z
lMtEHLTv/1Ys/c2PS6KJHPgmnpkmjrz29UqvWP9yyIvte72eNlTzIc2fa32+HA63
UDRxDgwT8pjCKKCtmS9elIvaNo3nI0WbrkWrbqauWf2mat+gw6WkRHnG2QJm4OiT
E+yWDvn08iG552oDGNxgJMUrviGMvVouuARt1fEPI7+Pmp3QHzmDjxNPZbhpJHDX
gCAvrxUTG0wZuBWg8w1ckkGuAr5U7ptQ6zWZjC3g96h7vsvgPhSwzqmp7qCVEFrD
Yez0+Cb6Yu+1G9/9pMqIdfkjD6ilG8G4Y8lJ9nW6iJ5O7CdaZTPrkp+ge9Owsdfv
DggMPXaLgR7oH8X/Wsxe/evxuVMUrACM2FAPyo5G0fZMwae6ZjmGtGn7qhVExITY
NYrmSTwJpUVKDdxC/l5F8Vhatd4fplWPJAkeX6CloLK7ux7SV1ah+JLT8pC5XeC+
O+ZPgZ6jPZpVC/DfCTpyyNn3+OcLhUnhYm1qhryZQeOq4n5LqNSBPVy6gBvjW7MS
2zGqQoqrDKRZ6bRvKz1sozod22l+QeNItUSFa4gf95qrdTvcJ+AcHreIt+y2vWCu
xQjSlLr3gcdH0QvqOH9fGd64Ky/7zGEBfuC6nICvzX4T4d00aQqu3rr2Ooa0f5+k
brpodisfPoRoFxag+8lVSow1ZVhN6wNuSbskrt1Sxo09EAVDBrKLwGn2Qg6oRBje
GYiILH3sE4gzwhVg2kE+7MxiCgKX06YDr+CfTbJfLv+ch2Ao/xd0Sa/bnwlCzY5f
3O61W1cbfSRj+IP/mlz0lZHuIJAdJXkhgT3rel1KJLHc8gl+9X9MRDlXX81fX8qs
BkoKVuG1CEDetfJIsStueBSPagIde/p1ztq9cKqs033QbdgJjRa1jaAxUXxoNvyY
D3yyicPhLADCp6Uh0as4dhZl9nBBW87TpfMy4U6+A2wKW0z392qLDnpGUiYEyACX
2hu1dOMBURE7eo20c9+Pjd9qWr+4r70IVa0F+PxJYJM2GUwQYULCYBAzWTZo/Neh
TSVfOMfN+Vo30uj82y8tuJ2faYxn3Oz9FDh39TA5gEqUKaFtG0moeUPl00Zgrh7y
TwIMab8gjbCffJxvF9or6HVnTsnIcHVpzoR7tA0GtDgrh5hDNhU0IKfERkpf3fQJ
49d1EBsGHmoFT6tz9SY1pUP+fjnQb58Vo6lEClBcVUaYkfpJ2d6Nxit0wfH/+nkI
WdiENo2sfUZN+UvqILbdb1WtgIYU02/0DOdxlY6FDQn+ECqAIm/RnsKJCzIrIBpp
UO1N1smR4PTgmVl5EHdAV93J9ana09v/IoDQK2V1qlZqisgjmSIqSlPzdjxEDZ46
RhLIPvjh1AVpskVc5oM2GPsDSJMvEvfsisX3dBQTXXE6Mab6TBMQTqR8T14t4YC5
Lb6stq/WI6SaWlH861vdHcIYKkMMjISfc0nhks+sinjnLUFemJW/jsxpf8QiXGnE
doW5tQrRD19EFcEmYHsr27e3Q3UGzFLs4OXD/8xSCzR7DltyxvCw+Garyc1W4+HJ
ZtwDuU4Uf8J3Gi1cFIDh6xkB8W5AdRJshQ6qDispRhGsBmDRUhfucWhXgD/kAsoF
+WDUedfQYnI3DVlx5j869e8VlVcxvBpmD2DjphWifE+mPNyI5uYeuUAkxxnYK4qY
Ujkq8jfiORklr6kszh/+rRi0FcHPGWraCzk9e6h+fuVK+4XC2am6dIzAaV+wdsuG
S2uPpVUaGHkmKtLI0lyEI0ekDVDqFUNw0gHl6Y8j36HP/f3e5+jGKIcy4fev1rol
heqnJG2zgc2ho0GRqWA17ilXGr79DsKRN/8UaUWeu0hQzBRvZxnzANJDWhiHutnV
93ehFHkYIVcTVps0Wz3ghckrOAh976IPXS3iHMY8ruIGFujn8SOa25dh3rJ+kmb+
SKL8KvIo+2EaVhKDCErOUBWFn0jTTA4B57erAkY6kDSBFGqxhybHa/vP5CWZhSbH
t6TZy4vnz3eWI/ShVmuVSlFr96MXaAiXwVAXIIW0XfHrEEiAl8vR0KUFpY2SqiDA
/05KjOsi635q9tKmFL/944utGUZ4iaDWqlzbg/6F9FV4FCQX4If37eZaZcEA8hxF
sabBWZDUFkXPlLHqgsVCTuCteG5FjyDypXXca78EFruuUEjxTNfzfmfCGRX0ELpx
q/JpCvKOGnQnT5lvDXKIu6QbFINSzwS1hqBWrlqODlVx6TfWA0mO+nZlwZOrcwlc
VJdg4rbR+XIn/Dpk6NLYjqweKhu+/K6EmHmAzgADTs4LBI9HC2cnguqiZ+gkwMUd
JbFu6irYBptdvoaZtb+xaVZ8qz9ofjjW/s+rsafOEZmojv73EgiUe+ckKpbk4SYC
QNyW3V+SfrszFMyvXA9SMAbrc1MYVsIhJZgO4GjX7um7x9x48PZD+zR94D0Ny/1/
aL4JQt/JKSEz/pFt9ZiNsYWz+9Tbbg1JIW5/vRYVrjwlFDwQKEIMOwnJlAs4YzaR
utTCsuJkIK71KJ3dql2eg/Zd4dpM++1nu4RRapUAiio20n2jTXEkeTLAxSAgVQlc
h256Sl9bSkZAIDjkfhRoIVs5x9rcQ/gYRWhZhfYXBV8ZdaXtSxzR1sh1WeX/3hFL
zJ8hW4DReIiWlLHZgqvwiNF+w/yeOg3zQDJkKvFQ/uDWXCOm74u/UdVHO/puqFLV
CPF6ZfWEJ31RzpkA6YYJ3fczp2mkgORUpQQoKZ093XQNaPZ3jRjkj7sP4qzcKErs
4G9IREvbtKjhLGbq8TxVnPGBJ0aVwLY3ifZzRBwtISEBZarxhZq2p3FfJvAq8b4q
ZGJUfuJJ+2gBubq8QmdXwJYgL8EuAWSaJcWoHbzJRNYoxN2EMDRMkS2Rq6YY6aEE
lykHw+YqVSN4jbZyHre2610LcujVFG6/T16g+Nt4SJI73HwGLpDlhmBGjsXQ7HiY
L4GxhyABYrLJDYF7Qy4BArgLF5+5aQbCKGKqKLZObYjtuMUq2xEz4WYEiey/6+gk
E2+aiQIipbFWAedQfLXrPWvKuxgTbNMXzvnMHjcyAH7PtiER8U6B7zUIAaZYhgsT
MSbGe0pQ0n4LEGev/2exAEbQPsOKEVhZJn3YA+zzWsfXriz7RzeYba6d2NLdn9XI
xBXqxAGG7KW6KwLT6NCCBt/zQzAzYkAgGeDRxd7PQF3USL8+/k9qAdy/AA+7eZ1l
RvljYHwpcQb2GjWilFZV/JZGJAUwivAoPHKlaOOvatg41Ry0ObIWASBmDmwQXKhn
SM8+VnM3CZ/PSnQddPPTft/+kpm0ZFOburw8O16zF89lxD9b5leIHW7bTEfcOrK6
t4eTiFe2kjI/SF6pWoG0izdLd92Bx399ozp4990mt0lkMOVtWrUwt86MOdpHnJdY
14SGv2KmLTH+qscpv7nJwzyXyf4i0IyDarHxHgQPZAyAzZQw0iMEORFLuwOyDdbj
UHb+1FohBJZMYaOJTa2Gs8qyC2m7pffzl0sjiWzp3ISUfpWaH8hy9b6+InBSmOS7
q+IWY2IUCU7imH4ngkeqOf2/nZ9GDepXCID81YKISABkX0dnsxcmM0UuL/sRFOXZ
YmX2txTioXzS2CtNVJyqnuOXKa6UeKPD7MthoY4zPHJh7bK7a2nsqSiPReCIy6Dq
a9xYaO1zFh+6Cplq0xoafh763wOy2vSnBcF65h5F7szIwirk1/E4hhpdUvrgc5T2
eAd8NIiVtFQKTX1UxWeRSpPHQ6zRZqnniu1uMInf7r7uDXIzO22dgG4OB/+YrT2N
F76QNMVEN1zxyyex36q2ElcrfQcXqHsZGbS/eknx78nop4tvkUVolpgEOZ/h/25r
SDwjQ2s8jMo2FkP3yhV+DAbOBd2Mw4K+cb33sCSOq/BUgzfxJBM3mZJWhEDRtBiV
U4FXUmqdmhA0rapFAe6Z9IFwVaYis4SsOhK6varyBHysP9yZDr1XEb1cXZKlqMfB
JWKYWVx7dEAHd39UfbyESh+k+ULzMoDV1nloh4qQqM28pPJiyPSykA91Kf0ITHK2
GrPD6W+4TGer0tDvskDG+dYvb83HdMJEhD+ZbiyVCcEAwJyB7IfrGQWTftBYXK+A
0OdPL60XSDRcGs6Rgd8r9NTlzgqxpgbDjrVfoiH9HjMYS0MU0O+A3VpgAfO83bL2
e2qQN1r1g23Bw0Ei79y2yJnNQ3RyIkn9Ixpq83e8Hc4NEStUjOIkygSOR67jfXFy
u2CujfCZgTxwpCz7WlnMIXKZOVaSZaW2mutoYftIZu6nx6TyiYa571yvTCHH+nqW
aBKoEotE34iM6auso7TiwrFUeBV6hWnJbaAL+Pn+FJgF3iNq4iPytH4pWCySzZSO
rTNfrZ9RTcY/rApUYri4LeVN6j4lXTqyIWcvtMa/r+lQnnetodzKbHBpUWsg08X7
TBH5Hrvw+NiNdODkC/IT5bFDk5bvieihNY5yWHskqkEyAwTJXD+WL5NrgSlqnQ81
8pi5yYC0zQkXVFXdeu30X7cwHiGQElsyO694mAkA2PeHcDNDq88kAXIdBhDiKGY9
mJsHJiNdEU1n/+uecUMn+gkXcsDaUO6D6CVD9EnYrCxg8SN01cWRuRaOrMtcy7Qg
RisQl4iiSsonsIE6SN6qUq4NdtYDawtMK1R2hE/UKfbA3OlEdZwrHDPxRY5Vncuo
yvPTXta4W0mM7JmvXxZ2YmqDwtxkYQkMQvdvz0lA7bBvq7ZU6xnFd6HR5xJ5YIqW
EBEGxatC//SIeTVHfhsPF4Q9ChHjQB5aF7x6Hj+lSnfrUms9d1GJjCR61kKwc7NZ
Cr27kXHjxJJCxG1EytKxDlA7HBrhwaK8TUAjqApyKYgyALgEO5WU0hsowHeil2Ry
zOz++oLCpea471lcTzxUq11Y4nIqi/45wK96eoVk7jwGug3647CsXzrEcTjvg5cH
9dTloJuwzO4IqU1WNsSyI0JBTlMSuUj04dogkO73fQzKH/V78RIzH49bWIu/QUUX
G32QpqbaDHEfapYJag3uD8VRr8WmUiiMg13tB3vgfP6J6OXorJ4rKAgkCi6JNVOW
uXt6mT42GwN1IjMlZL6rR932nXB5kX1WEH+QUezQAi+uQgZ32GyG+5L3TSKT5ZdW
cOL5Bcc2ttZv1Vuge0/IvxCqWNi7qpQpGnyIQOgxnhf3EccN+Cf2rQeDDz0mKhfY
zpdvaAGttMViaBgKu0sVC0rzlbu7i/pzsNlj/Xl4sT44CKTK9cLG8yJiATPgSTmJ
4kHU/KP2vr4U2Oy2KJoMTrtvcrozvub0YdtUsPD/wF3WWZ4QK+t/8j5rVa8uw/AF
98of7zJ+oefqGuNCrsnprH7GiSThBzJh2W0HeYjV+7rZLOtJC/NDfgJTQMP2XuRj
Xbs6fZlWLkWKzqPnZQVRZ3rZNnaNgd1qnd4Z0WOrXfNQhg7o2HDyOd40EOhTUyys
YiY1SjIfxVvMKn67tLWHEw3xS/4EtGZA51n/eUbUxOUOasZoVNNj7MD7zu2WiJ8z
IDxU+SbtIRiRD2EffovCtkjjuAvCI2TjLQrenTZ/tU0vkQJ9ihB6STgxFcJRqIZA
2UgHA545YEzt+zzMWxzSo3oKWqwN5AHJLNTUWgrDWpaEHJmtn9vWC+8i1qscI4rR
8TTKQW0Q/B+7TQIjGRvJCTSQ79e0Os50nSUhgwrNEwe46UlRqH2dALzvnfoKnXnx
/xB+J1RB/8aoqWENs7IuMeU9jM/wcuIcXHh2Gx41awXJxJ6v7iMeIxGkmdqEHgM1
8Y/ZtMF/+uZ/W3EbYCv/CcWI/9Xp3sByzNeojmV1Ll6CZAe3XZoP5fK06mmWR+C/
xMRnZjqln9OclMYTcKOvhTIIGQLGXYa4R57JjvInXPhIW5t8EsYHFKlXSoFWdsNN
G1yP+WR97hgRqxrvpi2/Waffp/J/X/K+TNH6hEmK4uEbdTYlkIYS+l6i7gnwsOPm
rnnkYD48Qocpsj0ZF93AVkmlYWwHM6GG5XZJI+E/DrQR19a6KNnI2/nIpGX/0GoZ
txAeEl8McynlkmUuu67vSO6I8qmH//eruAhvEoGEu+gCuU5mF9xAGIdwsfCalNyL
S/Q2mCDnRE73nwz4HMw9hTRkRkfIdLafEcdLqxR+kXJowVbxvKlEgeYNEl6+zOtp
lDZGZsU4sHeO6WhCyOGXXVRYKDK4R7QoNJ943xzaFm0/GxC+SMLtEkMs3drFN6oF
v+4uJIHUBwo41QxhMUyBrbOg5i2f6fX2nwAD5lfVisW28mx44rwjQFsu8JNQSI81
0xnJH5WXnkK26AIdANTm1/1mWv0uqNbxxTwsTI4znzMJ2DwQVRNLGtzAkIXR0n7+
P2cpaD4azen+Ha+aXyq4SmCbJTN2QB9dKOdDZWG6gQnGI7Gprc7lWwm4YAt6XXaY
JGeiNbFZys8VeWcZmFeNTg8vsVsNIUa8+1VORog/zcDHaQpJQ5pSZmq7WrR8rvPP
B98fi1LkcjVR0q/jccf7wQRTFKiyOqnBblx8t6bOPiYTLn2bAZtK8FAhN7Cw4nBq
Qs7fjBeF4a2H15aTwNeUzN40H8T88677hPclyhUbkucjglj05k6XNWTACRBaOe0g
DhKyfBmbr+wxnjS94k0ZP0L715uugTqjyOich25I5+NB1gYpzJfeVTT6jeEJxFJU
tJegTMt0upNiwkajlHzigAHihoDl0AMq7BEpjndVDrmFIBOEA5FAFSBCEmYETkfb
f0fwbYKOU7WWpiYoeiFxkR7yTRSj5NFQFtNJlmVLCC8eQxC1UuuMk3Nz21ylC9eT
2h9Z0kaxzJ0feFui3doBGUOS5fGE//V1K+8Ir2ax5zchLw7TUYVU42rzLkAX46Vd
l9O/4YpaHUgNRbzVzqi6NYRIwXtmh4nUxBN5pcvJ10Dt3BY1obnjcPlVv4tg/rP5
DOLBLmaN7WcVqfve5MMst7lJRJWr19bJ3OVtaOeAo3UoY1LLyzQsmFiL8U2RtWRN
pK1f0pTr6EVx8XBP7f+jvZWtKgCFuIwC1zU8pPn5g4OGqePvjmAyIuHK9BOGy67O
tp1B+mjnDJq3LMbAGTEpHlbk9DdHQDtuuI6Pk3/oIOUvN0noH2AQgy/oCiN+ydcB
aZr9rhJMSdmV2Xl+AGEq7HbhKP78PcZBIyPCsBOFUHV+TSEu76E9PFz7W8E3By2W
AQ/tPPxbYssvi3jPuz9iPrjZCfcauXoSdHj31QGNGdQjcxgnTsRHtJkiuosURYNp
TngPRh6Iwxeka11/Uwukf5mYCbA92n+KiKJkXiE6Lw/Mqsv0Lf0q+O+IIMlcYvXC
uaun7hwmwQlDT61V+UxbBqNGhr63arEgZcVTJaEk5tKhmaszWqgRkk7KFlAIoqzM
SsNrodhiAxritphpSGlsKTr/qieegsh5jSstjD4U/abZExloPPgOLIvj/8GjR/Fs
hc3Vh0ONqVzjyk0cmYJ6WbY5YmAUg1dySMTVsGEiYykOKYhPBoK3csjtVCcDFqCG
sKvsm02Kn5SZ0s97M+qZnm5c8QJ7oaZy4YCu4SBQ86dBPaLbVUmo3Og8JmBujEWs
Y4XwgR47pH7EquCgnwRS3rvFMMBl/BF6JMS5x9fxjqGsBS260PROvLxJ6KCpdT35
Jgnngv+0Rxr2VO8kdpIuDEgXylmoG9fmEt4kyWb3v6Sk3ohdnrlO1VSfYKJH1wvn
Vp+D8xynQzygkO+uK0Nj5wG/Sj+Ttco7u7S/oyzGTf1jF2yEP/ZiBdjhNqhjYxwk
DuE8fCJ63TTRn2jHH3H25Qvfq3D13zfQ0JinsI7qpj1N61tByLh5ZgNjEbE82onQ
5o4J604BHGDXsl28bdYlGHXBuFW9GN76rMdoqfMYswZ7VUT6dpX5+xvhyK7eRfZU
4ECTZhfLQGpUqs0SyIN4XmKtYgY7I5R72ihDGtrjng1/S8Te7AyI0yZ7xgJakOCE
AQAerVVG9f2WXhU9pAENAf6mL9X7a6ZznX3BwVao8tf3pnBNMtf5b7UlwuBNBs2D
1YW3JLMb2IfXHXHFjk2/qC15eqnZ/z+0G4pyS5/eq7VKgbVwoP5AmyXOrv3rv2VS
ZqVMxefymSCJVvpJH2nmnqt3jybD/IfCAXhSi2GanaxwdwrONzj3JKG3eT7o02/k
REfl280D/IjUngDsIBQYbGE6Sg0n9xwbQI3ZksqYNeiODoOK3rkAau9iYQ6GbPub
f1SRraZoGVJDadBXOf1BAQxtCZvvJz/ASimICsBvg0+3Qe7jlOAI1HdDFkWOvAmL
xKDkketU23O/uPXdjpMpp9juOQrdg6nfV9x+5HUONMXA7/hMwDQX7sh1V+YAiXO1
dHKBu1ZMrkaa4UtJECPD1C7cHzxIiZnSgBjqqbWZ15r6y6TjkSW39soj4ccd7F5V
IS/QiNq1GvqJ0oY3CwM4GEtT6utRcvIWXDSw7dy5WrVpc7iM/2nugtPVr5EiufhB
+QMEcro0KOSH4gxVmF/pmoZBBWc7NRw2Bu+zWufQVbzmFRK3adKOMWj6vco2i5Zt
eGP7pKhEitkjgoTrluRd4QjW8j+10T3JZRj8d37PuBQKTy0S3uk+FlpbqcjA13YY
m8gX/xeMCt36KTQprzTrUVhdPut4WbEBzzdvQ3L7Qiv0tb6Dl1asGPGOiyaG+6zj
80VOLL1iFfDRkyJNTq6mmiuxDE4liEZx1rQKb2K3OhJaFGXz7JfoHTCa2LrofWch
bCpZAt64vLNNXBxK0f+tqttgtnhBCdx0sG18HiVFPKTbJJFgJ3luOh04UanW/jzP
B2v0Ls+HbWLqQ3MM8ZTGzcrbSu0+q0JrQcUopiTdXr+K9WMXPJtzYwiqs4ZCGRPk
v3uKbCaij4pSD/IEPmxNr8BqInPXtydYx2l6cJpTRfBsv8+oANQhMTepl943meUO
n0IE+HiRA9kIAnOKWlnDSUF+dxNbJBVb6Yb3/xVqKlWVQHI0TLN05LKy++/MRPO/
1OmXzxwUboyJPY7Qgm66Wbsm1GRgKqrn6+KlYsO/0FSR5b3L1qb7AuNAUOKLZf0y
Am6k96ewL3sCOvLCx9L3JkoMqY1ZEN8t09JVBLOUQVSm9qxcp3Si9vVYyqoCZ6Xi
HaMO1NbLGL9DGnT3vW8wQpuB70ZwFWJpf5X2lh4CCX1ZcJ1zaAwcHZa4mciq8PK/
4E+/kH+/wizGhAqpOvgvobPbIoNUUh/tTlipS9qQFzH4LQ0HI6hUYZE+L2/bRj6r
Q8maQibgnmcbWxGxPw6bmIZchCHhAE50r5/p220DC+XhmP4zRU1c7vk3rSwWUrTg
tBkmchxurTdCAgw/JqwoBHeZVZVmDiX0SElCmGE9Nh6miSDtO2PTVSgJaPBM10RA
WSnO5bv/rPTLFLGH3choJP3jnijZUO2kO6lL2OANB5gAuXAnHSVIMjqxZM8WpabM
2DDoKG7YNKactsnnElOICTVt79caXAZgnZQMtSKd8+xSD3ZwBhx5+RfXGoQKXjvS
lIM629uKBUZw/aAWzJwAqXCGTQONy1hrzqGDrgFFISLj29vt55wYgHY28zBo8+QR
PEBij42S39XMcGQ2WzJhndrou7xMNsYUuYfRsU6s0p1saeB2Z7sa1i0oyUr/lnvO
P3xxry7RQLJ3XiKArwE99MjQJFYd02eb546dB47JzcDLMCdW9YliqWpOz8K1X4Ab
4Bpm3kK8f77X10WEEEiivi0Gfp2VPPhCWCR8lXQXFhu5FAlBZEG6xpQLvyWr2+gv
RP9FKTq8FSMeNcme8b62HlGZSSHgPLmLoDHCShO7aVwltvO6o8K4BQMde5H4kFQE
+pK+sgyAverVegoVzfiBS+s7syviJ50pzRcQ7vCu//w3bL5h2iY2cvyEdm/wlfDK
QaFWG3zNpkW5DQH5f/tOLWbbdeGpr/2uLoKH8UixMQinmMTIWVvjXov+fn6KgczB
dF94zjUvy7Z/S/23pgJ9HpJZlhTJz+XRE+df9dSwJi65kRE5CQmTh/A5wcI2QgbM
YIACebSskooPpJhQZyz3CYDm2+Lu5YzTDsry8CP61Z8cZ7NU7w0Irte/nk6kqvUY
Y/BS707+9QSnIsfmMkxl887DQcK+d+eIXXfEkKut/9qEKpBql1I6p03dheCxV6hl
RsvYSdsG0p7Tg62pcp/B8s+cPbq2DzLBjSblcUDsadfeQHap9W43LWC9El7Odt6z
o9zKj/x2O79GQArWoeiWBC2W7fofp4LsiSEOngQiCxITFgmcgOv8vg30kjOermGu
v1EUn6GGzJ5Z75thhS/N4qpIKhfEDYVmTExuM+NS+Rh0jHzaSRuqkFA6/Y0XMiHD
EyGjVHsnxl4MP1hyHWrvW1zFwKrkn42mvoDucv59oEgH31/dui22YV4TmueHoCOj
2qiPTYV9fXP3hh9h8MzqCdH2X6+Sx+n3mv4JbS1gF1aSgKPNExHgl4Yf5h+fi7Qq
iSuafA3NfVaZffEp3dBlCHRYPbZ+IvnE0iDAT8X3jMaUkc7Parv4PK+URDAhTE9A
clFpae6NYHJRfHdJeYR3P9Sw94/aQ5WGgiSaUPO2quVpdDcaYZEPiHeCnWus4mBJ
9viuBSuP36j+BDuYK3eEF8LsmpHxtOI2BvFiAG0QXFCkgVKApAvHrtd71+LvKDLX
C1R2rCxgbvyAQnDQECoM/VsdozU3E7Jd2QRLgeIafDKO37pAHJYlhhVH9P5kRQ6P
fC89swH0x/bqyB0dToY/F6AK7427WDeSe7aMJsV4mfhp8eGGkloDHi5jogZAlIt5
xpV5O0IZrBbsfB1Oe+7/I9ZM9KzGeSowbPT7y+uNmYW77oaVuiZ4RACRAm+HPk9g
xrZ7msqYjLsuqemt3I1U03pFVs1mXZhxXtLQOBf4iuYjyx5vqtKEkCOygPDGvYRI
S6LgTy9VwnAy1wPSmWurfMT6gEzG1rAJLFq5JM2I2zr9SQEmcwD6J+ZqdAsDWgo4
8UdRHgckOrU+a+C9sFGJV0Y7jnUAIwfRZsmctNxtjNwFuHqJVFEtK1SMUBxcI1/M
Q9SE/Woj40pP3SaLgUhHaGhdRnQpiIUNsF7cvqRnZN0T2jG902sgH8TAtzxMqJw0
XFZfBY29Pu/oh+P5UCV6Ey4nN3iMWSRqDoWf4xC/5Sef1NLws8S/ObtPsWzzalgB
QTo2QXfSIRI4SPLTUfyM7JNhTH2mJw/DPiYvva+pbvGzvy0yHP0e2AA1mdZqJM44
75inoTEc88x6rKAMp+wsdZscoWVxahMTNesum92PAVWP7RiEpzJ/7MjbZCK1wYUk
OXieLG7pg9NrGAkx+YSDkIPm+vtStlBaN3FusdZRQc79zVCHrH3rQQr9D+xL+Agj
JT+R6/zE0hb+mTfxFj9dLB0uUGaSYipdvyvHZ+n631qWUbH3B9nrkAMxO9blLlsu
uInGe1lFwlqjEWW85sfZXVKooRATYMZMkYSya9Op9WkH3WL/45cOUaYuejgsnSHP
zNVZWqyzqfedHN8Qnhkfy+kQgqMLRrFycEH7WJysXZkz38MfyX+5VaXszQoc1sES
JLaBzWHzUxDR9JvmA2sDqNmyoCVnGVblZI3cNZfxN7Am3RGksq122IYsmjMupqRM
Bbtl9IbfEPDzvW6+VCzlO/U40NqrGJqOQGdrxMAANh3c71Gw/mkhwxaOq0LzutzZ
mwL/E5mweREXrj10weatpcPCTajbkA3NG3VEBdtQiq0oENZTR7zpZGQAcMZQSZpi
SiMI3oYj3YPiG4bSb7VeYBF6PBdmnKbggwNfcyqyhJZ0lrJ+Zj0VmSBZ5MBmaXdL
ZN2hdnu/DAVbg1j4bWjhxs/EpucwEe0hiROvqjiBcFAanqUobQrsQAsNvCktXNUJ
3KCuU49AdAO9I5SJQG6e0KqUqW+yMIbuUmVtsEfJnotud4vTI5WuVRBCkai405vz
2qMFs6Nk2X8I4MI6PDHV0Ux8u9HZTW6yL3tfpBCUpdW+jKQ2tz6TvLRbcVoO5OMr
++QZE+stIx+pm7PqXrYPDbmB1VmvpUbwffkla/JBLchDvZ0C4s4X0rD+fYOABGeD
Bu1raUnVgfW4Pl6BZrC8JyByt8+Vd5wvt+NqJk9ewfQJziZsGv+fnXXl98t3lZA9
a8XsLgGGHbpCf2kKf7hiRAUnir0odW8TNxVrFI+macVxSLF/5GPPw1uJxsAZIohb
rJoDrB04dTtbQ0GIZrHw3CLqC56f7l90ZOY2GoFMx64mxYmohYhm8nOmoWFPjACK
6soFt72V2fbcryBGGKJwuWAkCMINPzgy0V05QnmSqjb21+BlsLExyLxuvC6rK7AP
ApHr5r/xJDTGCAhltPqWCJ2RWaZk1rIltvkm3L/leHRxFU57p/mHpYjkGLuinCJm
Dgp9ZIxLenMDnHYvpOeFmrjd0telT6RJ283wvjtuGzru2kPBa4ifUPmZFDWzxc0E
ubBqrOuHXJkGm8dBx+VgL+R1Q6xrJX80GDN5Ac6QhloqunFBHGbTKyl2BqlQnKz/
EJ4bzFSjm0m0s6Ri8ksPb3L6sD7GG3KThlDDTAJRwv+PpoZLkooDC5XBmQ7mIS8Y
Rv6O/Sa8yzzvXbCAEdR9SlrsNI89Em5YHbO4i2e0kJ9s5tniCIBwA6Msdlgy5Pa8
h/15DOhRfJOj+O/J/yyO/6eSQWf7hQOAm/N9xlH9wvBupx12DsYq09jD4Tqslibz
24EguruHEoWr0IKQE3Q+Xxxq8K4JHN5hnYpOmYTh+FCvfrLxEGuHeDe0iW7zIP+s
qBzN7Dw4metw4Qbuvfs7PrsN30eoJD2m4yNGXsxcHPUKRygo6I6aQunBYzuCdwes
LnH4C10VQqhShLtXHXNBusXVSkfrjPMkM0xcLvHmspk1oa8QdA9MyMnAdAJR5wgw
g4TBwgGF/lrP3txE/3X7BjZ4GyjFC2jAqsWjcl2anAOULDnxN/It9bXC9GS31jUL
6TeIrSE2abtIOnyitRCsRhJI5vjjdvTwGTszEY1TRgYjB+z/uUt13WbIMH6zs+4+
JzaT7VoUG0vzOD90QCJCPuMoKNdwspxZvV3lKxNoVhZeLrlxjzDxj+EoVAXdeJOG
2FkmED9IW6yUyFUq6TQ+UaRjBYgtDKmeYa2dnsCTmgvuuO68DJoTOeCu98D/BDIT
7oTnJ23UItDhdu1lK2PIzAnoMsYsJPChOhWe4c5aKLXV5kZ+lH1TzSl+p1BLMK92
0w5s/DomADddORZ6VXK3KZNET36/zbca6LuznmB8CIFwa/eZZEiqH9zybFgCj08u
tTXrDPM2HN4+AbySu0EsOiJPANv/AuREbirhndJm9HZObGxskhHsQ4uN0TfC/LUB
xXtrbBG18E/iSzHhKd2dtDrHBvFHgEOSF9x2EfrLUPFRp7ApxnaiPA30tTMvfCsh
ayvFAO/d0wIiPxR1XIxB3RaxDuDSXsS4ox85dLnOM3JsalrPgoQaO1mby0ZGWdvb
pLG780fGyrxC1uX6KaHlXNefoHe206zyV5aWzyA5/ZHRC2y87UTcEhe5ga3ZJWjo
WgEmK+9sV5PLMNj9x4oSsYDCrBADnWNPnkntlors3qRvtVuE9mDDtRNDEkZF/tat
tWz9zy3GWRl+DKlSbMbnYljKySO/9ss6bdVavhu8g/rEUTOE7CNnWWK9Q4IV1LXV
9wxBdirjCZKe0gt7DQCsYN8dceo+Tp6lP8LdY6AW5s6CCfzEtaLetc7INA/LBaKL
Z/6TFARtLTEW62zg4i/x60l0ZGNDE06UDNWV22fKb/H9IOk0mbUBs6rozZWvOaIX
3l7hF4VxrBh5ECv3ARV0xBmPu/Am8rhNQQcoFIdeP2Q8vRjUajW+geVtLSKUcylw
NUgrxE180GNgylObq4R3cg3jlGaWZaPJCneqI4+OODe1GtnfrO+VS7qy4Wn3Y9os
0A3GhSPby5pLjQQWCqVXGDZmuqXQBcXiyUkeez3yyMdLEYq2DuAmRHlihznXgW+l
GZuN5Q73lvKP0Imr2xmJMrOzus3KpLPhESALBrfIPVUsrcXI0OiKIBRpe3bempiC
/yTtIfBvj9XKl/7sOUmi4Ne9cwWnFjI7S7punzYo+Q2haAihS/4lsfQX3NXxUUSG
D+bpGCHJZvcC/QHU28wBOGbt7uuX6B0TR5dwHse+9LHfZBaIzUmpwrucHrid6BlW
gYw5uBKpfCo2WrDz5X51fq09dtA79AG/1ua4q97B4Bw0+EopeMsysvFP2tcfF9Ol
UNHtjVu2AAiMkhbu9bKI7Ki28IXrGUAS7udDroa0XAhS3Nhk0FQf78DcwBo6kjat
Eg48rY/YykQQMMtAs/W9sT3sylhkrTZIq0CmGB1y4O1qDk66Lpg6yjC/iZ/N4JCh
CCnLWrYUCNxiBWdN8IIfgZDRITvzySXQYoyAYZj39kYKnjHiTkVM/UbXhXl9Pw4Y
GkEFs0zAYE9tkl3KzPDpAZD+tUNkn3ijXOQggBim+JajFMZPmVlUTC8ggOMRAGL8
8JwfXMRCS+6a0/S73oQAkBwvWZqJvESa5xDnrFRFZgTGRvpwC7XmHJAItkdnYzUU
/bFc/BC6jejxDh59omGokwxhqe1qvC8OUnvhQp8VmMP9CdOV9QUHA+7nKB5agSyd
2LExbWu9ua7JA02zCtx9TTyTZ9zJmMmYORuUoR3SpNk9aAzbgdoIHcQmBQTGmFRa
a/pDpLc6WkNbDPSjKClA80ULlkDZvs21OZu7V635kHBplkyM1a9Cwq64SQqm08wh
kVbti/HQGjaCtvvLeCdaDxY5WMP4Ye2ExEjVJgE6I8Le0W8n9Yrhtrb3M4Bqfc4I
bcgPlA2qc1k9AdSn9ik3LImViuM0xosnezJVqmjPSS/it21Oa5q9AW1kngs8sAsA
V9xrhcBHKo/yDr3gGpWgRR2Y5qNT3fOjjwka0zsMwaf6et4PmKX+n587Y3dfDV4u
IDWzax/9pFuq4VKfHnfHExFirK15yjNUlZD8/3yp5ra/cRCtXNPFaNwwuBSJLVbL
+kaK/A3lxagENW6LFHnsTHN88c01IaS78C76uZvSFdCKT1ZA4F04EzW2P5i3QeKk
FjAucszlY/eCjPDMZy1DMHcUP5yQGc/RaaKkHPdqKM/lF/gYUeSv3qHEl370r0du
SaLk1+s66NGXKPxVPHM5+COGiXFYz88A00IDDahw4Dlcq95h942DMltvma0jwS2D
aN0P6xa/AWrmH5mXaDlWQvwXM2LM4mgWUhECwF7UCYzqpgLFXN9eZBAIJeZVst7H
gLau+VkTtqinBQXqw/qsBB3QnGV1Xx9A7kRWp/YiE3L+GDlMTX7tvIdlt2VE73Bx
zZE23MbFJm012IqfUs6bNZHZ08eoe7x3JzDb+UgAAaKpsm2Cv/XHxhMs++cTqqDC
xHqKWs2RigPl90bdfw/KJhpDhzqL4eo1LJ4V1VjInhTCCQ/ElkH3K8ghPzLTwZLC
s2AGVzXTTMI21SDbO/mj9R3vDUIdL93wl++ZmszVKEiUusvwuOxjxHVH+EPCjPLm
bpt5ROWuxf313VQRL6yQ4Po7Ce+DcU9F+CNLeiKnIM898oqgYhfheqHD0HF7x5Jw
kCNxATIDX6nj52NKUxVJGLYPu9AMeZ/V2cK99YRUuqCyajl4cBNT0G24E8UkqlGd
TSGeoHXLwFMVXsk/143wABmiXrTXpsZqmbq/1HkdKdva+bYATWA0grNJ2VaUlppX
xB2oWvKhkr1nKBmcVf1Rcg9vBY5FO9mJJQk3R/Ws6qfmEOOcG8XbrSOiAQz+tBsn
OFffWIT5/54ZasfqPgRr0c/N05+rteivJc2RUAmd2gyJVVNQF9W7NwP2LJ69jZCh
eDOKAFFXp0xW0T15TnIbXjGGwNJ6+hmbokQkSOzr4fZCyT7dnuDGo8KcLBXiSZ4a
q5PyPLc/ZovDqNH1YSw8kIwy3qQpJq/Lwp3h0Qz0bIm1bcPFBO18OLK3UeGjapML
3ekYOOomLYHw8kVhejh0aw1QyN5YhmMod6hQdBbUJJBzynJxW+S2O4rEtuGkkM5w
qBmiy35kOzuCn7+xIXv3ZEIkfokQOJj7OyMnh950aDBAkuenPuYWxCd/crJI7tWF
3P4XsNXjbS8GwgfRKnmi2e5e8vjlWgRDRyNfiUqDAt4OezQxcbczh85dvUG4pBqm
hEjYqq1oTcq4nJEX2jWmPVU5irBaQPudV3oZziCdl5IXajk2hlqoOycxOsFrgBpC
xwi4688cURk48E81N4FTgkR0k3hddBDJO2oKqpJlm65kO0A+F0n86jVMXEZuZ0tz
AnVbEEIE7bGW0hXo9uueDBEFT+7Fwn5xfBkAmOlwnCEQYHru1UXF5ZENiTXXYx7N
Z9tN0kBTKhLgoqYy4/dT9XZDLjzI8Zhq5vxGyhPSejfX0iXG6/GAcZxvhD/VRD6b
ib5oRnJEMxE6YEsYBokrOcyy3RGtyuWBPm0JGNYJjdtpxBmo3xcliyduOW+IFZvc
h8+Vxfce4iiEGfcgpf4B8BqRApvikTnl9Rg0fE7IcllLR0dYT+xxInx2ODDHnr3n
vgiY+tInu9FlP8gCSu0Y1i8xx3tWMebUQqi6GX5K+EbZfBQ0LaJ8jVriYglIzYXm
38jZhI79q6F4M1FjAodRdEW0HLUt9gO4pbwWRiVxTEIp5+PJag/m9DhGlNJ+NKOM
EzpN0r3hl9RVbyw3Ulb+RQkeGkv3HdCW1oPmy7mey1b6pemd/8seYYIAWxpD47m3
a3rqr2LtJid1HNP7lIBi+Vgyyy7ZhsZkRsNX2oxYj1yvx1x2UY+VuZohrlfLkRrJ
uhF1YTUDIdT0DUKL+B8o313KS9BpgrAqP22d8aE3IJROvj1UNbUSQvr0eq5GbSZh
MkwzB1suBllDMwLqFiIbof64pP+dQeivCDwa66bLhdju9jcG9tecMGNyt4pal4tV
dJNUp+wSyvE0HPnNgT1xXRM8sQhf5Lde8rchn84hOYT8pP9ZJSzfgIgZIs5ULBQH
rM8HcY9cGmDDvbrcqHot1Y4DSDCHKP1C8lxUTYP9cLzovjzxpKzo7WceB73yRoDO
c+mSV9jA1uoYmtM6KbDHaZQhr5RmpCvGuYFo5sqPdUncQsT1xt3uFFPpEAVIwV9B
pdD3+839MbiLdOo9TthwlG/cTGS0+hYRh8mTF/YlGxe0+X/T40OI/yjDRXM6Nuk9
j26xBbLS9LtXtWjFalyjQYO6ecarZ7BrPnATfui1876zDfn3buOfXbVWu/B5tECx
78wBqbFdY0975z2KcQO7dAGXxquyBvZBtCfrFrauKkji8/7EOsaVJuQYCct5aQgG
y6YDfi1Vf6oWQR1AISjWiCujmTl0kdikq1Kqn8P1eNno3icyzAXJcM8Z6FI5EVmU
De7fiJu+JBei+dB2jDu7MEGH92gBDs1xKJwNF0z263/MXT6jeM4P9eZSQgMEGj6x
6FyZ5zph61LsKssaPCcjZqufk3JvVaHFA4PpFEhB+481BSOy4sVahU6TH6tvoBGZ
R5q8QyJ6376aXbAzZnoKke373yuFmzhRdNTu/vuzUBi8ZhB/IjS6iY0KGwqHJFIM
ccRHSaCOAqw25fizSHxYjm3Bb+P+EHfqC3WiTz9QD7HLoq5QeMW3+GzSTVbISg/s
fWTwPpJupAapiMRRyPFwio855hiBjB7d1ALtk+6t1jqgW408HgE1k5jFaMJDnWX7
Fq3zVQiq7k4U/bqcZULUiATAUb4gs1ZQNfpwACRVwM60meoWnkpH9Ld6dN2cXCgg
JoS9HNdUPz2myMLJojkCPRXR+tnLVvMo875xl4eCRnVIubyHnAFtBEsMj+hZi7UK
lB1Tj8FlwP8YRq1cFLtOs0eYn/F6/ne1vzWsZKlfL0Prx8V+tnif9abXsMY7OYzF
YyQhi2Vum0pKvLogDds1v0QeNagKYasI34Cv05N932WHBEhvqNXKb3FJLVBc9Jer
xWeTj9exEQgDRbVkKthHSOkMryfLuRuUq4KPK3N3ViOpL+fpgSedkZyDNINbh1JF
DZYKfTU/EA8xyAiMMUF/pj5zEOVqGFnodS1C/NiHEhuWqW2DKUlACXiISq7/hOa9
casNYvt8pgeKhWMGysXHKTfjHC61EGDTBb3R46yE7Bea7+sNX0al09kfmjAu3RrK
w0E/V1kGkcv3C8kbht2EV6IatuybEq4BiSGkzfKrkw0m4fpWtNZgdHkH05F2Mf0Y
nRbz29Lraz9TpV/kS1LBon+XeRQDtC/CP94ElIcJbepEM8oISxKXlmvb2pJGWdmQ
4LQaXiB+4zotNxF5FbxxgpBHBYeodHE9xquHo3/7P2/egZpqcLWJyfnapqhm6ttX
6K+BUCA5LHR5I6qj1WF4f34+xfDQNIGHQtpFUHi4XNubvsYx3uDzVgRECdZxOvLF
9QEvJXwop/G4yfiWsyAzzJencWfQTnbmPVCInZgGXR1A0p7GR3Di/+0VAW0AJOzh
VSSRjQEPBrHDOt4y1lZCGa1E54+Kh5bYDvx7P4t+IcNKx035moXkYCUIPIhrsqjf
U8T0bz8FCTphVS0zfIq00c8avtSuMH9kr3XJ6cWnwMc1Mdb4KJ9KuqshlIMiza/q
J2GCa2NiRf30m91MFBE9jCTeUxTYlAT4CgfGUI6C7e8L06lxhr2+LbSR/RQJHGJx
dGBAcY5XImoN8DpVfZ1pcJrt9X78+JczHZ03NbhhopuaoQUd8TTsw8J2LJypSN1o
0SiVOYU8sJnP+nRcZfZoHNM3OTFcZnH/ZOLlo+jpLcpblvD05fufUHd3zDFI7vs0
xPuMO7QtYxmXMGdfEIzZE6Okks1zzUYB0Myw2stRtXCodzJVpHvws+Ygl4siBhd1
oBOOSL7LZ7hO+ZwE/YA6TCUFOy5RXDEy7KvlGJGjKHqMbknGVRAh82FMeaA/+MWt
ZuYHN5rsG4Sqnw/FChLnhBLlJRuATKdElSUsRL9X8h8s9XaAYkEaPnGPlHBqNgiH
dT7e9z1h0nc7Qs+PAsDcm+y6oZqpJdP+iOvmoWn14aPlE2kLq/kVZsTuGDLCDYHJ
CgqTF9fYJ91rjClgNPAbV7lcBSBb+7FBB6ZERUxFKutz7hMtHYTGLGbPCSFRY0Qb
qGqDwUPc744l0pyu8LgHK06emZgKB9HefwMftCZ/dyeb9R1IbZFhHfHagHfS+au2
zxUXFkJz63kwbmO7mnQ/SSmo6ddrFnDmHphdUOtGbmFR+EiNzKL3nt5TvaNxGnLG
NDGZ+BvBMu7fbbXjhjPjYelmpxFcM4yQmknyN8V57IBG01U4RWGAfiJc0ktmIgzA
i+njdkgAJd7veoVgEgdH0NZdg7OGzLTLr2Nob/ZbfrFTo7QZ9GHKKe5i2srtKl5t
RFzdzzhVJu4qQAykGeAYTdpEu91kj6Z666BEev72DDZf+5kji8k3axFJAKVekdL/
bzx3TN+R3fMHMjRz1r+pi/51y9jF7Nt2Hn4ToYBWLjC+jWyOsMq4CRLZR+Ld/gwY
26whnnEDmjv83MNMBKuDrkD3sCr0oh6rOZidO75cNrNC/OVQiQw+Hs9DCjxutHNu
XnPqDrSy6Pqob3KXthq2A0TIZgYfAPVnN9IVlnQASo9IGBhusbyXHW9HYmjkYlGg
lJS/7JmMcEaZOJRO/nJnbZEIjQATGpTkJTrWU7egLQ+SBHafoz4LHXcWMMwiSsI0
O8Zz+A+grVZzvz9ZrMNBiQijTe14VC8yP02UWg+GMonyGM2t18JbGg17V1ZQjlPk
UnRI88nHjFHr3146FiB9UvfZf87uOXoSlJiMSR8s51h0AWz9oYgvP0N26VzI7G6a
kREBrHrf0xMoE8WmcM6qIVgI6cCmY5PHIkUID7L9rT+h4PI1SlhypxFHY4YvP7P/
N5JmzOPyvqsCiVOMKsBUm1JNZ3nX5EP0MddjwWvzKYd1WR0wL92Aspyv6SlZVo9o
3CQmI81Ka8hR0bOZXNXBdErZIfB8JE7jMpdEdZ/WtQd60E+diaBN3RY6hNuYevJW
5pnc8UxPLYnOQ1eubUXhwNTEcNSBraHKDS7ynViKm8deYPK2Oy3B+JFAhNOrHe/R
L0WitM1AuGRMy+zzCHWlCnx4MYSBnWGCGTCJ0mL3poyCM2MTALSbChxgpKIELsad
5YBY3iZq1HTETWuilZNs7K6g5to8/Qt3tezKUAXPbIBNNvMP5tn3MJWFVc/XRK6f
ju0i/TXJaEvUTmw8j1xbF6+aYeKBNkNUiY6tneQPfi3QQSl7XwJYXBdr9X5jxrvj
ahQSFjjUEfh8uWTyB6AupO+7lwAPpjDtn3woZ4qI7qH57WSoRASQbpOBZo6lbLZT
JowKuiUnfrw47kljrEWsEE2/EEwlfuyxE8i4LBaBgwn7qpF6qj8F0IcRDP0HnDiz
dwrLbUeuxjivzQnNPNrYbi4CjemhqHUH26TpqUhOhd9QLKjNEfvBaYnUSh25tBQg
xNpWtuFYaj+wCxQZQgX5wqccn+lvnCHzU+UcAhA1IZplbUiIZQ6QXFspkzsHFBZN
iCLN9mJ9mK6emVNexAXdogyfqWCIzXLe5JDfDqD6YlvzWp+gTxSeB5Sk/J+40Bf7
HCSMjra073eSlepkIQaKcc2wHc6LTRSN46AZFwIt3/s051x+iy8ue/HaA4NN45fw
j80VqKcedU9lOcwKRraG/YdIn/UAOjDFMu/cpVxkkoA5a/lTk7Z1ZIm/TCHHtIrD
ax85XOGKwJEZAqYVPHmMydmNxP+igqNOdf8+KY9j4qyChnoYb77wWROLl5Z7EbYw
TlH06YR7SjiM7SRQcWjO8GACvSqmZoq+ztxZ7/nBEkinJlzgxJL8VXbCdciSh23V
ekp9xdhvE3vB4OEI66yxx/PLNTrpG70/5tLDp6jvVs6obweQjO+StQjRw17CvYGu
sggN/Ioijrjr96drPEdFSD4B9IxL+I/5IksiBJR2LKHdCMkasG8XTgluWkl4AeHR
Nw6sQVjSAojQwS48Yle/QwgzoADWpt8+Jo1MGmVyO7erjUXMTqghm+sqS+NqzpRr
XN9PD3teuq8SjsFsmDMNV0TelHzAis5vYvBPTwKKfza3p6eytaSfydmC+ece094X
PANdkNp/YNl2aDTD5JmWH43wnVrAcqdhWsJzDka/qKFKQTVY2GAaKikpqEq3U4z0
O2UuO4apoC61FBE9++yk+cqg+KHwCgD0he5Td2XhucERKeIx2NFFCZ1ygd0Lfz9w
Zr5QLJ99K7pFwOX3PLQ/TSykAUJwkYHFqzYFcOBVNA/9ES7qzUQhCOcEvGbeHpZr
PXtfKdXK3SI9wR2EpFfPABL15M+DDUG3ZYU/Ldf04rIFjHyF9bh5xOv4Ds+XAxtc
I5XVAwN8lKyR5v4lTB8Ar88F/T3P65I6fDTZ/a0MuRmJ1xwvA1IdGO+hqJydcWil
TRVCIybwIem6cCRSx5veA6iq3pC1jTNf+N60PIY2zesbX84J/HqCAvle3tIuvybZ
NS/faeqnWqB2yEitDaqV4AwRRkExi6qEdMQtlo4cIY5yp7b5dkm4If83mdhPk14J
pG1QUm8QPUad0prpoMSc1o+AJAlxlr1+DJtEUoeC0eontlLuQOrqi5VMaIcj4MLX
MoKEQGpv8AZI0g457l05SQf8r08QMGEqSqcOOCV7gE+aHJnNsO5ims8/U6umT1pZ
Ypqf2r120l2Hei0YGNJpuT3mhhkUtBkIBQ9KPze1sm+7Zi3DqeX3npTOI6Fwq7PG
31RctB7Kw1u+cvImq330s0o7ph/exML8dhG0vhCR/kjQT9qV4oGvKC5oaYM1qZOt
KI1FTmj1E3SwEymKlaGlBUB5msXTjRekTnU0KLYQs96BcF32AQQVws16zFTDRZ7F
XnA0Rjepv3BOGdpe/JbAIZTAMxjgTiGNRJ3+BQDrjHK9d3zZmFH0Bz/Uv8v3VBlh
ELMvOnPUA6Ei3lbwJcJsNmD5CkEslU0c6k/LEdGhWg93aUzlBZ1oeoBAUQYWIz7F
5Ce8wYNxDhz6RHdHOiBNB3vqsSRufoLXbM7X7FD5rT99LV2Kciov80mrq9A4U6Cu
NpaTPdOBFEonYlOi7aZMVd+erdHuylf1LWNtmsbRjvTnPSFcyv+loZENkVdfVi84
pkIzxc9ULdDVihjmrybWVlZX1UsGScjO4qCd+u7rOFs/Xvrwd8BkzuJ4plZcUH4j
lpJX/MmcOOWtLC68uggE0Gx7gmXFwv3m6hszs+uUBjDRZqKLtBnXlctCem8GSGYW
JZQ7VPf7N4rEUT/aGKpzgLt6Kt282rXSQzEY+es6659FdQeg8hkcR4IfmSJ0ClVv
ycAy7ftiBdgpeeqrlZd/ZYtC+MufsvUFsfeyBAFmPu3ogDFUfLKwj3O4sSrlaWN/
qW6ahCf1w3yhNgRmzE/RY2/dtargiDSfb10s4CEZKisWtPyPXbK9zhEGHsHSVR8F
28uDiYyzJRqqy1pxVD3W2gNxZlbfNzrTWPFv5PN94G63/C82a7ULTnbwffwwkdpg
ASRUUt4vV9F3He0gH8TuGV1JKfZRI0IKyGoG9g1yHTU9CNk73W809zx/JKVrWYhf
D6fHS+EqsriEk63H2IIlxIrCFfOnCoJU7d+Craa/TcIGuD8XHDYjAWDF8l1P0gpG
7kW9Lu2YqY/EZ8PonNDQw9/zbghclmXCZJcF91BmjjKNvQDX4PEtRRqU44FwxUG0
RYkCkfVYh1MtSXQH9+aTYiihEzi5dVGxcxhZIiPkWIRGNeKp3pfuLQIii4BCpCc3
b81BMlu0wWQToxzfvrEsrDzavzKa07vZlW5PP2da330kaJihBi4CbezMvIROd9C/
+ze2e/PHiE1Mi7St4cnw4AW6HN59gBP9eVe+nqqmYuFqimKsTXWjwCa6sCmqACLM
OEqmMmdZGKkaEiNCWPFVDLYwvLSzmv9vP/Lm8mA0iCMkquKmYeUCFHVsEE6vj8h/
TjyXYu2q+TZoMqzu4dlWDojhH2enLOnBEVRV7P8YJ+KuNEzkm/JBGcwdXl73Zq5f
Im1ptfYlJc0g5muYBp4HkhcczFW42gexG07GZO6ssgzolDJq1H5w1LgZxd2qC8xO
KVvzH4FcC1cF1o+NiLLRANPJoVhzdiKYnNr/O6E7sM6iuLLP1HvBBHats0WJRGs7
yrm0g2NzsKmlbK9xPDxnNGUv1yZfErcU3XMh3lAZA/GzrWiBDr6/dbQa/xYEcgQj
ry2EGGAf/uFIHrLLyVspYoM3iUlyIr3XO5TpHPmZ8wHjQyPmtIy5wqma60FX45CZ
a7RJ//I3nfM22hG9OW4DD1Fyw33cK4R1NiuQylC6IbC8ErLN94SDCZH4w77//TfZ
s6DHq0fjljs0JYd7mvkSR4zdXY2JXsW0XtpKvdaHpRvtERNBg3l44ImaEq3iSTA1
wTlmaUJryCG7FfeMm1hf1TikeE0UHS2ynY1Dq+2ITqCmvP0hxXzljNkRXIsY30r4
2rMCqN21quHQEK96o0lQq0QdiavQLO2vh/mcztCW2dZe3QUk6c8uVPCuTo4dfOzU
6CFwdDVS9Ao1j3W//Ba5bT3nnbYx1XDxOI7VRX6v/rFGhpwbqg2F+OnUQIePb6nr
ZoKOVEBeCcRmlPLT1LrEqBYTNnYPC0WokjcTz/muGC1GbYEnsrrM8IeIgwKGQ/5j
6GEgsCvM1xtA0XJYQi48es6P0Iun+CqCCIoOKGyC56q925epfsfzeag/RgQ12/Y8
aFf5PFfhG1YA2/EqUrV/A3o6YtpsaYR43GunXI73dJ8+3v0eLVEeKLyWe7u5yERs
8Azi+nKWrwfhJG/u9wi2Ioz53Et02VBOkhJ2bopSS34zn5Y9pljJvOns+9g3AwrW
ejh8rl1DmcqvUhxqWVk1J/RU4OKliTqw2NHR+2ssvr3Qo0yMwQYHeXH1voJGbCUi
ycozp0FNnjAhno3Rg8deXl4zNsWWw1t32GCkbrvPJOzEbnYiKZv/04OholpHv6R4
cK8QmdaRxDNbZwfY38K1fXMMwmZd3eKzfCRniqIhSguq/1uHAwbrHH+WdrOvYu/S
RI8DbLcDc3Eu9jYj+F8avxQph3VLkGFSLuuyInDqjiXE3DU+GI5auVRUQd9Lzhng
m9B88FzsIGQtvkc6suNSJYxbzq2/FQr++S/euppGscdVw7U0JdCQBkCnAe64OasH
CGDXh9rdH8T0CGVIF5W8xtQbzT2kRBajn2BbKzWbMLIs4Y9/weHBc8TXegN6dy9M
3lZJ/KovEsZsvTl7CSOdsHA766bFRhxgItLEBTaSbwOgE8UxoP0QleP0TR72+1ss
SiRUvobvcdxwCmjfqhvgHLY93lfGe9BHwOfJ45wY+QX+DcLpFCA2RcYnm/gEO4c7
aElmFp1BvCqAKEYoo/++msTMMfDxpp7LtQ8ta7/33iUWPAVtY1cElIm9mijvrRki
dEth69nYnyw+XjAFyIpoIel0GqH7h+ldJI2h1OGyJ48NzGNySDNuED7qb2fdc5OA
DGvA3TyNt2eAhYvDAykMhv+NBBbvERQ/QUhgKf5RE7vp3wsSOLHbKO6ueHRHv9I+
Gw6xLf6r9i0PQDC33uEMuB8956qcmYR/UIqoSqFOGNBfO4jlGnz7wHlH7yXhiayR
Yl6X4KVpDZgvkmEQ9UwveozMG0sZ4ZLlEUgv4VTmYqHZh+DInMieInhRlRoFmkuZ
ZxlZR2c6012b8MvvyM1uXB6KeF649RZK0wAFoIsKmjy2p2wbPjznQU2mvkSn7YVg
ivsURM09CMMPk+t44ud64GPzsUDCpnhpVA1VSGnyAJx/g8BM+uv2NrgLCavYOaPq
x7NiOibTiqlOPfQsCe7f89CiHGxhnvoGETl1+0zAig4T7Y2W5PsdsRG5xnMK3f6U
nteCpJ7d8CWSPQuiMjXSFsnpN05owTs7U+iB355JPvaiJpB9gNWn9Aeh1nMulaQu
J5zQn1HjpP5OkdnkmuYWPLl51McpGLOp4+QkRPubIMMdqNwaezzuRptHiRUrIoC0
u/B9p9yH/TbrbBBfPZQojSogIPFkpsB1m7koI9pBCRRIIXbAeyiw/cg5mOA/3P3z
0KpFbNq6QKcDsUIaO24VInNJTHue1g4MxgrHa6SWSx7xKmdkW1wGKKGgKsEcHqKp
VH+6DArKyXyNtMoVP8saltqzhE1vbSgBtlN9m8tx0biTKYQ9ERlPmhpubyOmcnic
dRKAXG1R6SJLo6uzQj0+7aES6GvkcbAXX9wGgBB+Rbx/NL+L/KU8qKcRxwd4b0sC
01ieBe0ItWneNbcLLI/eD2pUWk3mjjYCFuClNyGUlB07p0NyH1NXNHiQhsnc/Ux7
Ynm6Djd6QuP5SWRb0wB/SHncA0Yelp86+Da+yD39GT3j56dRHk3f6IE6teTFdr5D
D5Zb1daUrja+ZdlzGtLXyfgjp18QFumL930PeBrER/KCMJtzRLBz4kPWs9x1lAYs
K6gYfmqh4smWqiOdqpO8A6tA1LXLrAaCYQCI4BV4EZtJkeiaY4aRvAtfantvgGvp
Tmf/e5yIiJacckk7/pEGZ4hCnSjQCpVK7IdjtBNsnwP5slsjEMBiYBJrxFWfxd8/
aJibkj3r5uF6XvlFTm39TjuE6BVs7R8j/eW30dq8iQqAKlYNp8KLuK6nEwZDGMz8
Ut9TdlEMdNIBkS5/z72qf62BAho6NichyCgLp8pgPoywVOAAe1jDCgy2N21PMa0V
UxzgZiH8cW98A5TGqcopocxXDv3xeY8KlAvIX4omugcYLRmFwP7svTiOOamxs7uX
20uC48moPONfBwp7JkKniIYsaktIE1HDyfVvQajlS/6MPKiRdGObGmV+Z3fq2Lyb
jq3n4IW2rZCNJ8a/gaoX9aNAA3f/tN0jxuiml0kFlQKNAs6t9p4oLDoH0WVyDdJ9
uczryBfvzkWGw0yY7S2IA2mvtqY+bY3gvn9fGKtheswH4UBjfUoTyenNDPK1Lfub
tU+ItWf4Iev3VLpEkKqkmEGveMgPg3UDedim0N2s+O5kxJNsTv6ADDS7j/xibK8u
KSiu6OxV4yDSMEHW7B/63CDff+iSwauqYKcAy4a9sjx9AgfD1Typt+DvSvqsuOlS
Q+CxMOSHBVGuBwrxYxwr6H/o3SKkv/SPabpLqL1SxsWC60+IDnRSWcBGogceYQ/3
90YzLwAFSUo9ngRHbt3kcE2BVhn1/ZEl7D13gLsfc/F0p3+IQD4D/o3eE23Z/Fc0
U3tf79hPyvE1esi0ryJLhXobAZwhCszVUyRA9jTjJNs3H91Xg/w+NtJmRDwa/tK+
zCjs3+hTQKyWAyfIi4BMROyu96hqHY/Wncw0ElQ/8I4nawKZdHFXKEGHDz4PJL9L
/dwQh9GkeKWm3p0UXebJ0v48bCzIqIFhuTC5fDbVZXMpYxT0HhnBE9He+5kF7EAg
V9+gavJn6fadUSktJQHZZhWyWKd0upz/n+x+rl1bUm2DN5ATkv2k8B+4qiA1OxNC
0DYnh3vaXjEeyYwmvpIipywBOWf7XJZVVmWRa91ycUi3ditHLbQDgG4PrOKD7W3l
fH+rLYjI048r5gXS5Yvls3IGgOLtrUEjIZ+mYUwFRq1oXtBYiKcKEGrskR6UsS4J
GOTWlcx6IVBn6IGLeoDzuVtCPg5jt+L1x78w7gZce3RcQ8H5rUEyQ4oRcbiJZ2Lz
/pQdMdytwzZscgme6GWOxGWxe06U/AGxYC41Qlks7dtFP9DnChj5S1tLbTTyYfUh
km7yVYRwq0eqwwk90bRbPH4v8hz/m6MgxC22VcJj6VOvYQqYzF0HIQx6jviT8TYT
jZdOFm7p7PJueSdjD2lf6fYpx40sApy/bd168f6GMMydrYYmcIZFAGvaQn2f+SpL
9Wulv+Oc9MCHHHdDZCRNcAnv2ohnOIksXAQHHDmbAPtKSdbvVrMdxA3JvztkfggZ
xLTMiTkzsChPeQ1F/4JTGIm3HWSrW1B+dU9ssumDF6Tc2B9e1n77+sPRSt6lck9H
K4lotYcAXMRdbJKe8Fx1hTNz2i1B/SWzQ4muJKwdzOEdxa6SqZqB/JsCN+d8F5Ej
lPPeX2QaVqSv8sWGXMV5RPVSK8dCbFTF5YELh3fRxT4MAUDt+Kdp3s5FdrUI9p7X
qGyhlPS3gt5bNphiML5bnBe8BhlIqhe5EDr7zmynEQbx28XPvi6KhO7zW8pswwKT
anE8oArDwQNcAhlCVrTnwZJzA88UQGBeJ6D1lr/QwoJSlUntaGLa3paADn/2bAtv
bHoq9IAy1282AicdnThTJ0gO2yHFb+pKaf36owyBEYMlLY5iEYQ6D5jThZnQd4Sd
ltfoX5xZQO3hXbWIyYe24Aq4o2WY7J92oBR/eNOsAOx0ZHzspMyB2U5NeJQwCHyQ
zXgvN8EekTilzm9s0uhNC9HTk1PZoCgg+BuG9DWlqFaovlvlRx/cbD2XevodYbxt
RhdHEgFP4cgQSjv/GDOPbp/yyvMtGzSe/eoYZT42GbQktPicxxrCgK/wcf6p5T/Q
p9wejOha4oldiK50kngYvIrDTEwJlBIl518SyP88yWqwnsfSRUTZKDV7gy+MDpmj
Gn5mhdDopkrUeIAV1rCshNaceI/OM8nqGdlNt6vcSww3HGLj77yl7n/2ij5G0O0q
rkliyMCGSdPHIF2iKSHWTCP/Q52DoPEJCJTWIqRDNR1wWqgHRbYG1Y4edJdvoaIi
QhQCv6ayAazlJW0oLufoTHN1FQnuHvGPLtqXRWqbpCH6a4AlZymg9mAuYZcnepzA
pu0KBE1r3tO2Gof5COId0USV7JfwJDyWSekmT6YNqCHd9tJyz0z38l4O3mjqC9q6
V681okObK7mGhVnTIhzIxd5iNI9hn6dt8b0YTsvFeuhg+3n/7PngUm8u77vuxt5/
RpFApbGy0mfDRXw8eXmeRjMxsDdpfm918ZcWfQw8gAhg7uAw+bwYN+ceBoGyF+Nl
eS8y/aoezm1BU2Sv27QHJXnOE74A+qvy1n6vyq9o/5ooWj5DRDY4Y4MnxcGhhlLn
Mmfb9tqFyPR4BCyFqHemUwdSNMoI+/kQ46zLc6azNDY9fCjoaw6butNGFqm/sLM0
lsEpNFvqjtAQBlcTso6YBZZtilrqkt5gmO05cfleHUf6rUAmBAiuRDr+8LAqIxFS
wPgPNMlMQcYAPhcvpZmFR3u0YJEuW/11ym8Yg2dl3sHUSU+7LQSWb2qZahDSbOk8
WOGGY9y5VFOYhvv/iRAk3SE26isdA/N1WW2cM+/VDPWOT47qVQoIbUT4y0VvmT94
pkzxxkGgR+CdUNIpgHkRUFqW0USR+zji3NIcmOCBUG+3w2aKu6hTUuN+T+qt+3aR
9JzsYHmSEysurrHPhBKAgi0XkP6TC7yQfwqosSlG4u/iH0OBrLKBU+AddTt41QEw
gK3daJ3ns5vOp1uPXiZhvj1HyMEIl45j8+uwAq/ApL3nou0F3NXhAbEBI//uxGR2
oudiByns2id8bht1dX8WDbMCVcEQjheSUjaqEeR9vfRQyB2SZbAonnXiI5JUARc/
ptQNP37uU62DeSKpIrCXYiXzr06QNxRvhxaNp7z0I5R1kiXSqHfa2/do6Z91AJRe
X0LTHbujQ3QTsT0h9OZ2m2nsJgW6YW6fYJd4p3pxLcqOsw7Jzm1mn/mHOHZZPLW/
G8q8k4HjQzXYnZmOEXgk3r7fHyTXq/tCUDn+aJWDx6PjUqXM+9IshmK/wQOj1tAG
cS1D33OJfq5sb/FMtcagZOHCFrRTWvqXIbVHIfx9KvF3WqyBKg/gF7pPTCN5CZty
iGv49i4vup8qa02LNhMrcgXNhBddTBWveMcCeZ1Nw6oZx5cneir8AXeZqLwG9KH3
AqP+4QvJGh3d7EsZ5nkrR/3JxgMvjp4TwiWD8Bt+nwpW9gPMPqxXZTSnh+8++c6b
n13z5g/zlDAOvervfJYRKGhY0XQ4B2ZPXDstqv+qUF4hAaraPSGXN0pYTBSx60hm
xw29NKp/fc/7OwCgy6tyzysGU9kXOW1flWoNbgNQjiRHCto9E5msBwGZE/iYSwJJ
rZJw4ed9EpCV/ZXXCpFV6TpvjkzoarDVQ6hhuCl0zTUeLNNxi1WAzObIZWr1qtwu
7yqIkiEusrDKntlo/kvJytGR9kCF1saBpEYnC/VJIsq+wifP7C7sT9ci1mSkFEAU
NRohkbINJnie3Idb7mL6YiwLViWt3qvmPrhFZnoFuehNewtxuNCbgXnPJjCg6kUw
1cBwU6z/WTdqDonrCspkYn/MON0Iai1ZmHsAeCDmih/L7VlUFyL9o7GVMPUZChnq
rkVh4LU1RyXim+ECgR7YqBFfaua4sKzYAjZD9XKKZXBvIJOgiqOs6zrqC6gbDSWD
DDSn2wPV5Ek4ZSgXeMhL+v39FzEMG9yEfRh3yoD1yuiInooGHf9SMsOU+XgswE6i
vwKY5kKLvQXJ5KU1JwBfXQhCrduA1quzLrWTMaCit7qT/vfXBnd20XE2+ebbMlDe
dW9meRj2UahbxrYPqtL4cLdu9WCysyvy4ks9reKRX62ewlavK1SnZblqfubfp7wB
Gih1SzViGLW78RCydo6O9IsKjudtNPxnAeIyiCUmejU9f7BPAkUUUOtTA3FOfzoi
iGk/n7tGPR15W3HZfBfXeYuDxxW5gAGkwklQK+suA+8QIY8wMu+6fDEfZPP7IUiV
Uv4HEX9wr/o2/DTp0z+6VMXZUsL/cWwvQnuf30OLRusZ0CMHsKDae5u3j2qdKVSV
+C4CqMEHCWhuvKaCIZPn/B91uhX+rAg0IXszb7ZtFIxRYgHhDyKExOcAOPBfX5EP
GTn+w3H8chKeYYbLJOFCZvAb5LGiYoabQZ39GLxNLaG1BQfhtd/fj3InCJA2P8F0
hCmNmbPhoi1zPHnaMXtTXaG4aPwXRdpjPJAfEKT8U4T5HdGMNWgsv6WQi9B311wc
F/YBiDfEoAlDylH8gScritEy6GGu6ew6r7KrEIse78d+WxtwRQZAEzlILNNgjGkg
daLmjcNuWvIR6zkp3bajIEFf7p/gOc/nfkhx8KuQPzuqlQbyJ+6izvdhJSwMqsgW
L+wnRDSGfwzCyO0mvBQLko8JSkOAtNiDsb3Rlxbe2S/gAtZ1vY07db87buN65deB
LS4LA+KyalUwMmupLlk9PW0L7NZRmzT/1ggguFMSWgmruZWnTSRjPKWhnUHp/cx9
JnB+fltG++svsjq2Aied05wd57uEHgTS739gIwIqkJ0ssNNioxait+07ekSgfFDY
2k8muJWCeWQYj/MyJAY3JS1MnStWRXFr6obcCYJNoE5whhOXfpWC1sFbIfGy1ov0
unLvdJ/IC/BlsadfC3u3CyusdLdwyCgeBrvt1aRiz46xu8suv5JNQvZOHcWkyoNK
1opTOzrfEX2aj9g9OS9R9n0inGPURAXJdWRH1ebrnXcel5lU4dE5YTsqWz/TmLI0
iYW8wE0WNKQt1reAQ+z8umnMqV4BogBXMsh+yTBj3WxPGG1bnCjB7v/eWIXqMcNy
wylAuVrLGAe7GV+5d7qdwSVM0gBrcduYsfvg7shOeUmZ7e89Mnb8n+5dXtMegIu8
C0kSc2J9uurvW7aJxL+YtqREw+kqNmf3QBqafkCUkJKcRl4Kd5905uA3RaQ2/Mfz
aSbHgGKK8padIgRMhDhsq95QgCeHlMEJ1F0M0Pk3ExNi//6eJnAKL2SN+FwS93EX
0A92M1pr84IRbWufxJWOyrFxUYv0BKxy0T+2jL7f38jU+0N8Al/sQuo7CD58REVO
qar+OKLMYI9eaxsix57XVQrz5Kw5/XaakT3Hmts9m7sPUa7iSO27Xot7+W9EPwy4
icBHWMIZ7jwjBkobPOXyzoClfiT8YXpSSk33VtzUO81wfBaUOEMU259/Jj52xzns
Bp4OYk7XMRizqLOdT2PEn9LLOYNDxvu8YWLhrZJQsLTFTnUBbwUot3dpQIZMHWzD
199LI4ir/s2zHln4Ibr/Jb7cYQ8mSy83Fajd2jeMahB96GqooZ7nD/gSgnF37gqV
zK8AOp7UbNDwcuDnUzZv8fe6Pfq6lF/tYT2EH4BUr/3uWTUn5IU+l+IDNX6RV3iw
kEgpMbwDg65QMHFGouj4mQ4zMWGnLSq0VsHL8/RKbI9kskpf44pFa77RVuaHBbNY
GOeUQjWRwu7lVL8SfzPF+r1yfwZb45s7ET7Q0u6p5GTRdSwjhy0dSEMGN3TFGbcl
QMebLXJO9ku3biw/MhFLtntZ8h/EMt4i46Fi/Gd03bKSBLidRTTYc/D9kDTKscIP
6sjPUQRo3pmgcUjTEnbIxZVLrY4NxSOBphY6Ivdej3+LK6jVEsMeYbpJ3EKBDKWi
wo1D0HiJ4F/BcFT/FgDs0ddWmyoxKiozrL+BJzOq6EpSQQwhgt8jpIQzi40zKtcC
a7hSj7TnCixJ4Sr4ELSPP8LWucyuiy+eKdg87FtDQ6ldw6EyjeYdUcnzE7hfrnNm
E8OH0aOq8/X+vZ59UtsYBKjAE9Dgsfd+yqlhLBmGGB/y1FrFKT70au/T0qjWwaBc
nK+0Cem9nBi0csUm3jB6GAE2fp3MaUaOrPcJ/SAe0CP3iA1Cdctw310yxYxqnsZa
fXwFk/Aomqz0IDHGnVv1gP2CQm2Iw0qxHkg5qYztgWyMeIEpJ683h+SruDtH6f2F
mb30EnFf3Bdpccuosundg/jQrjUOcM6KbjVFUCVjdJMiYjCwzX9N2RY4eUuojO5i
OERGaRdyO+AIYoWxIQubidzUuDjFlpzBKRsplkAK7LiQzEFmFOgvFrr6ihj2aYsq
Ow1KA/+iw2v6v5dD2G97ugh9vQ88EkxwJuk7xcUuqkcw7zBnbrk/aUIG0lchslxH
QBtrm/Lq59/7A9cSDo9yrBGv32A8gTox5ROfVYGIoMe0LEVsc9hzf0LuJqGRZ1gN
4O1DbSctetKJi25/P+2ZIrirvPMoZlqdaPosp5f1kNODmA2mM9uAmpC2i+bOBO67
VKKe1s5HhqzIrQM8reVeuHct2By1GjQH+8PFTwuY6sn4gfBLYKiF6F47aNkdlXvJ
7dzapcU19nIpMiBcKsaIkEyw8N7+KiuS7VvNus6Th+D5RAtL/SZYGY/7zcuo2kXu
VIY+wNCeGc5GB8QUHwyFvM9kYOZyZDUDedov5sFlQc38Dk8ODFC6uqwx2bTt++Fc
5S6Amua+d5bkcM5Ih+1ZiGYhfV93TgzRUGUDfowHai40oGwYH66gXCTGwlYsIbN2
BH9F7uAbnMt784S9w1RkbK2D0M9T0pdpgS6s3aSFb8d8FoWM1Ter6rGvI7EZpRAv
uYMYqis+PV9/dqRnjXoW7FmGQRCxFql+AkLIoAlfEG2uQ9fNsjJMr3JtMsHie+uw
9Q6ETabvfqbDDPkcrcqMooQjcNO4wxD3nXDbCv1Dc45URVwTvr9mITg6vlDfCBGR
5Gg5e5G+7CFVzXiuMS2+49Q7RxjgdDcsY2Jpw3FLObjlBQ1eLUz3QlrCX/elv52D
AAoOvJFNQ01qA6XMz/SVC2drDGbjfMoLjno28QfKHIzs0yjxkxVlI7GZlwC3Yu7q
aPUFb7Hsi7Wo1D1q7i2USO00YZ0B5Mq2iZ5qWhcuLXa3p0I1KWA4KtlAgiMdjES9
t4HJyUjAqFywBYMu4DRPN7SOAcDx0fQcLYlC8PNPAjPzSU+GKL6fCoOifxvupy+8
sEVYtepozsvAW61uw0fKAEUycgD70JGG5CdyV+Wt1bzfDiVYnL0pYKaKIaAtVtRX
kljgKGGDWve/58tLSXJmyHlkPjS3bn8Za8ueZS7N9gzSgcTqcZ4bII1nz5t8Wfu3
JyO55FF52llAMkGllc+PYqBxRL+jqknaGkNdHqLmHebeyEufadzJubdbotSxBcuz
TR+snY/yG+NgUk14g1OHILokwgsAJkVeZ/1na6Z+A14hiTljmMKIglYBC3hdP/iO
ArVF5jxQiCmmVntSJBdyV731pIYDy53MwpO/Xz0vumv7wk1bWIJ4EU0SLrHMuPO9
gyscYFBgNtXn0Pk1QRRa2ySPXYT3P4VzdxnCStH5qbc02mQn/lJqIskhtbqQx5iV
cJ5xeVwKNuLKafo0cqjPnf4kxao48p+pw1tKfAXGrGjgMTqofEsXv4aDAnJ/ntim
85QjV0raCx0zyZyVByC91hYs/oBckel940PH4APSpMnFsn1WOuTmhqbv9J4cjTf9
PFww30x6Tgq5fQqTssU/6rPJ+u0qhClT787QwEAUTyWDNfo89fnZ59U0Se5Ce/bf
NQ+2paKzbbOXTgpdjUeOhAQX4wVlDsPPxm8UOANvC1k1ExWANDQvK96BZs8w4pwk
e+SZEg7LuyZnsK2ulBOVNBIwBrSoahDzGo8OL2nJ0/KcY+qkr2S1u+LrBBDxocjE
8k0+BwAaU0kydA+mJWnzMyJaNhwNMr1uIEwrGdnf7O7h8zRi/qGEb3YkS1QJ/U1+
q8NcAo3MCU5N3oKq/E8Gz5ScQpS4t8CR8DaMX8Vpl83LeHBGMOUNPeP/ZJbNmsDY
cJhRVYIG588GtGvoTTTXFkoBFTfn4FXjZGLAERyB2xByY9pk8TAkeoeEU/HR36uO
4s52BKigHKTztJz3H29g/rHvutHGiJOn/S5Wow8tullngn/dBlbcvT1grc0iFPyZ
oFSpH97c9O+9giK7KXs76X72L1ySh5HFsRZ1A6gwl1hhyQrzwjdYg4f5fxSXcZ2I
aEdWmdro7DTTxmdYDLClGOzIcIGJ9ZnhzlGVmWVqTuFTybSIPLlWx2N2Inue9PnB
f3/GYg8mrscxxudpqnYnTHjEFiCIgLE1XrUsGwdKKLB5+Mihjb9fb2USaDF2sjvA
lDXqITp0IKerO283I5SX24ORk4FPq8/SNlwg1yXEG13QUP+uRDnDCt6yopZoNflD
4mVIKOGvkcMl1MkIhj/Jc0HrLK+RvwFt4JXl+4M6aTc2fXFM7zwkuskzYc75jxlz
KCoDk9Z2b0/YJkg6/ujKj+EOY2os8CqBRF9rZLDKnGg8PpZ5Ml0t2cTJxxyyvtoz
bjHiD4FGOtyCM0QUtyjRM2quyPn8l/Lx9s4pmW+J1EZLKMPRPWiiCc8PtX1QdLDc
BYBpE/oxHV2PNHtjjiIn0F0ZYRhx58153HUDW41m1D+5TJyCrcfO6T3dd3BOTwN5
pmFiQdtyLwZxPXH6CXa1u08K2WcTVrmfM7M7OYSPS41GglOkeQuRs0duk2WcN00R
y0yjKf4W5oACF/4O9GCwJg5GUdaMurMjkbkmZx7q/0z3Bldsw2IkwaMR+sXEDb1x
CacKGW3OPv7j2jjDMJ7oNFbBmz1zCLXVtzv0XKbJiLYLxNmR029nCypf+/mqRQA0
Evn1f6ECJUKF4EzsvmCy4SoiBk/Z5MIqGB7V9UqAV+M3jQSXFx72SG7bCKelSCwo
LNTWL1AI9AXlMPePxEgaa+kUUa2y5zSTuC2VZZ87+allD/Jj7gRmTQ72YWRwIK34
ZYIb6xuH5h63CbZuPKt+mcBV4UYSb3DMscEYKLj3v7M4PBia8PU0+CHuLaLjcdM4
wuySP6WUTBo46bm72Dz25ORzUwiUiFoNa4WXc2lXrh/7mzDtk9vVoWsWc4lmff27
UxIUImf8aqa3Uz3kkcGGiQFqUl0z67iBMnjP6iIwj3xpQO0pXNACVmVXEc0PkK67
DmlRI3aP9bF7KUTQypPGBMo0Xz0TLSEzChzQwSm+5xz8Gc0kiJCLJoYw4mG7/tQ1
yjbx9RZDl7AtcAqZNm7AhgzorQBQZ6gGca8+lwYbdbiRAkM7sjHvZHOwBjUXi+2A
MqIIsJ6/Yoa5sPKwu/wcs4qYlIp4iNWwu7jRlQdisOynh+YeyIzOBJb7c8WgD1+J
+TEUeTABIoVHh12ztIDu94wmms3i2HOxz0pjUsu0dg9HmXJEB/7nBLOMOOOxRPBd
cDaMM/97u8RxTFPJLhs3CGcYD4ozt7Lzq/hhIzHqhvNUiTSvcRdUvO5xTtPdgDie
wtnmTjq/xYkgKS636klKIih8Gk2CyARUPL2INgDFu1oIaFRMNPh+Ldz5IwH9W0m7
d1XzRwhOZvjRzAkAdYaamYwdCcYi6UluHDRCmWJeDKLjdzOLmcxq8b7VNJrbamxs
9ikA7bEKJaxutrC+ZWTEieqFiaPXjcYwh7aLOoaJJk/ZAWB3tDDn53AD6hP5DnTa
PniBYP/l6x80KkW3Wmh7pj3HWRKKEi+lgMn6w/+3GZHaNO3X1CKiy8SurgcnvcEm
7PAZV79fXZKyn9whFXeb5n6WS6kViZiKMf6Yxl65ewysvdI2k4U1YUN2xCtT/R03
TGCJ/k6QuYzbgBe73dn1BYJAO/nimKj6KQqOOc5oVpRjMuDULoHBogj016s+YfC4
jiOxn30sbRhIuI2YSbUykEevnNx3IUPnly7i7XapGD31Igj0JvRMisIVCiJSmSVL
g1RVBAe3l1P/UmK4FwwD/ll9u1Y0o+r+qo2fM+tB7vVW0TRmNvCRwyH+gAhzsKKV
QZ3qKz5gYNi4Ct4xdDsFT2UVU/g3wm4WFg/rVlcVrLNPiV1VmXmDGk2ihwxWNXUm
sBjFcO7fWZA0+6YKCOfTe3ObV2978Pr6CCbodMm+66FJctzBd6QAnJ9Ypx2wVzOt
eRA7nL+b0+Mhbe8eAZiUL+7Dl3V2lO0MkDCFUuTOWVFwm5AQ1DWM7J+WEfXtP+sn
VZAv8mo2X/v3TVnXCRtWQkZtNmjBAKExaLZYi9nkTapgo1Ah3lpj4YjVjmAbDvOa
iH3J1uIbDh4Ln5AXarstc/6qcIdQbtXHcyIkPP5Bi/bPnPqJmsAnySnVvvCEpee1
j/3XXN4TvKTh/6Xx9n/85lraM8S42uOLZ1yDvgN10/DLylZcUBPmREU6vBKpWG2c
gLpY9hDK9pP3yiZ225OP+mCdJGLdiEmoJPfxISWF8smNOR1u+/VAXdeHssBqPGIC
2byoVT/+hGgQ8LHNuoTG9PKrNo9A2DHuVFu9qdXNKvqR1sW8AqjV0dt+sHtyy6lu
jbPkSrhjzUupqZRtFDu6wuWSuY4EPGkcCskLJ7/1419mbqw9UbcvtFTfRuku8cQx
9Nx/hBBGzjA+ahXD2M2g45zn6gvaK2sSGON9iEIR280Elzi2cUp86hw1UAPZaFOq
mbWHnRo3aIIXzq+InfPJs+0vyfJbw1yPtgykjAhHdTdWC89lmrPwc8XdjJEkJ0q/
Xyz+fEbZC/c4EnSibt/JzMpWOCS0Ru+2+tNudavTP4NIm2vQ9Se5Cg1zEG6guds1
kAN78SP5h9E7UzIpYp3gMqdGUAsvOGUdZn5LU+A7Gdhxn98QDwWvst3eNVerQSHC
TKlFhSxtUu+2QfM9R0qJqOgL7/a21d2T/C22mOuy5Q7U94OplS2vLw1WlUUkNQJz
tkefTmWVHsiuR/PEBg9aCrgOxlNzTVoZDFIIh5kmbL4es0nNACBS08Ppfr6BPwaq
OhsUvaJuz4OVvUbhFDjeI8S5Q7rfFc7XBs/vs3AF713uNSMBgbKsMnVGvjdLFiZ9
e6eJdnnpTp0eupquZBQ4fNIBZYy7elC/8lYN6u7/jhsvMbGenydpULIHZ+AV9EG1
rSb4EPtDebUdI14mVjRRSa3JCWUvg1DQXwPA291gvNfOr5b0ZnYP8Tlqy3qcxsa0
3Rjq/k3PkNMPXRjSQKOtPzpPLO9AMi0OIQU/ZG65dmk6n2LNyXhf0CU8EX3YgoR9
3r0Dh2CaH32ERIAr+3gWlXBd+mQAac43vERb4c/kpQeUwxhpsovVlg9DP85KO28p
Emyvtnb63ejZ3JjdvlQHKrl545dTufwS14zYEpfGtmmoBKQrcExtI9zq1H4X5BRs
Qr6+R2PYok6ssU9jqlIFalFv9l9QppMcxfewnANeA/2r5j9vc9jAzpf4Vh68zKSg
XyxVnFkl/Sa6ZF3yv9XES05oCQ/1GfoRUxZiL+1YuE7c1vheLueTR01/jbeyilQs
ywZqaJGuVgUg99YrOsONvzCBguFOdTGe7ATahRIkJUuuCBMESlYuVsdvh3Oh/GuQ
3tNpgodwDmrewOXaHHlXJRj+Xg+EP27j3UTinNUGvB240zSjj9DSrePMAWIhCJ4x
Kyd8i+2i8rsNolrOZXuFGb9wfl8cxB/0qpDas796nHVggArzHp+YHCXXUTpLLl55
8oCy946iNihiFD4XPC2rknTkpJ1W8lQRFA+BS/7RmTmCZvnnhczaBoOKM4WiQDMC
PrTD1flsQdOxrDv5Vw4hoQzq0K3KQBth784iOBPkwSHMbAGmesgXfo6o6922fmAI
ngnkgi44S5c1VvqBQkHUHdxcg/M7ssDqt2ZwbvFtChhixJnLb3+g0TopqxXfPNum
B9OGKbIQgn8SNMBqT+RjtKO3Dpw7V8gHbYPEO5lJV+9Dq7EG7GlTRO8JKAl41iXJ
QM+FcAqdIgGeXmOVwbyZFgBEXxKriAK9fpLGt4qwIOuNKwXyz7Mzi7WGgHtI4Khm
v6KI+5uM7FpDw6223nXu/NZokckBkf3pkZn0wPfVbFbtwgMOp6TsRMVknSzkaaKJ
vBrF1bh2sifULg4XcUlJwnV9ws2CVcO+0jNuOyz21UpEmj61R0PN7Y9aUSVLGCVc
v0MsUfMa6RaoalfLqLvZ/0YC3PvqTL8uhy6468TeJqresghHXaRp34X6+k11osZ2
WDvr6J2pYxog4H7ANpYXnnIfB+h0Exp7rblRvP1yZXlyjFD4WDJfUaQg+Z8X5yi7
kOnuZgBQfqvTeO6LMsKednZnRvyG3y8ObHAGU8FPTOxXPzMTeWPr7AcAX6LP2OLp
4XnCi4xUiBfKGkB4yZJjlQxGXIByTkZJMQsLQF7Mpy6s0yXB+pdgTTF1845vqPM0
GhBGvaLa13L7/kK3KzuyAj6ycax5hax2IfqN1djaflOV2TAG9s5Ko97YDxFaNX5K
JxH/NUsb9ZoQHxQ+nv1FBqumvG0LWPXihzSNgxfyVM+2YvbDUZ5c0JHFRbL2kbmM
MNFDI2qFTdELWGgfrnsenQwZTGcsjEMbdoe9Kz9VD5HvlgCybcHysyUWqGcv/D7q
u0CSFbfZGLy7h7IVeWB95PnT95fOHciKLzBaQVXk9r48XeQcSTTc5jG1A9+XuH3A
ghYv/Z9sJKwKI+8/RDa45Dos9PGd2e6XntM2vk7mgf1ws4emvc9DiPR4ZgoiT6lY
BqcETlmz9n9ApdqLAhI7EwygqJp4G560q5J/Boi8Y4VfpMoIBLgk2JhduuWuQWkj
1OAeC9H2IWTcTEguRpNH+9g0Zg9xFGfIYHUSG9zCRd18gHrT/FgNySkSxkeOeqdO
zG+1Xf70XhrWMm2SLuY16EWjbhJL23fLX76uVxB1cS61P+Pgw3M27RmvQT/uDtEw
KNtovC/Z4+i3XeSEBWgrBt1hvo1IASnlc2O4XS3ixMJC/efD6fMeXNb6voSz1Nkr
kfdFS2d1AjS7MTLAEvLGp5OkSR0VYoaWvs//fHJTkMUqgdR9GrjvvQ23jAzld8H9
OJQD1M/CcIeQuhZQnjNZ2NsqTwv34u/YCnWFRFHq8tgHvJTuNnzbfp3f4A7KkZg3
7ABmYge5eVAcPXpsWILYgGnXxFp6k8F3Z/cyv83hU3bwYaetqJH8itFmR3cYksyJ
tn1McOckSnZYqU8WbcCChhNHIesNsMz7mmYMlkdglNg00LLL9MM6qMY38Q7azCwh
JPH0UldNAIW25xMyjxX2Jklen9JKsWsMCWFMe8Y1V5KizmHb8wobgyYGl1ZDKNIl
jia3s0f6o0rexRGvorNNfsfM1NSNhX1496qj4YqAPRyH66V4mdEfMAi0BslN0ChO
Ok4pSyHWm1gImdHTIXxfKknaUmzwb5ykkjLmvQaM8nW8X53um7warL9vm713aPPw
PGCyvkgr51m6d67r9aSS8AQFeIPuORbl3NVmVneTRrp5ooUa4It/hGuyJjOYDkDT
aM41ksF1tWojpaOOacTz65Ce2sVVeCc4tcle03+zcF22NyyL7qgmFQ0uc7iR8ikf
A6MX/B4+r8u55TyckKX0KXCteN6VwIXX/18sRv6NA02VKGEfr3pLwJJFbxzbuCGJ
VVKOk/gsT2BdFw/mvLg9OrfjzFzkF0PwhOQvXDim7A01ArU1QFsmvTqiJh1ukQw8
FD6S0iIbOCNw1aTF5jVz6HpRxE1Xwy1t52TLXSgcZqJxNn/m4h6gwrfw76+iB5EG
wPRL5z4SYSJaRnliYhNmsAr0l43zlkehS5ZDu1KPT9L1sWKI1uMw/+/tCgqegpzS
dKPoMFppp1fycd66gFZR3RXFBgtq2qR6L4GLUjLQdCUdnBsmRO+Ed9FlaZTSv2wv
2NdipKwy+iTOO1PvztHSQB6DmEMmZ7Wiv58xuEoUNpYcWwM1C3Npu1w86bMXFsxZ
rhKuL6nnU0QlsdRoTUgBg1AzAYYpu2cSXmfcVBl2by9I+v4HFUN+4Ysgq73HckKq
bPLW0pOlFSeuxnV+gtbRUDkqc6cEmUCs6mi3wZw4PlTAVio/pLoQVAUDhAyWGbhV
NKzf2Y0DiWPgieqm2dbxEqrE4V0bLbr1fzWZlioZXQElpbkA1XdKj+Bzm4ioXhMP
uxLpBJ8Y8h5YY8vDCIDCP7LKI0soAuunQjYyd4kmk5Uj9pLq38Uc0tS0xHZLjDJJ
Iluaj2LP/gFSdqjchxIxelOPcZoandwNDexvUY5tVYWYRVP3je96qkSt2CrzsnRL
no3aX5GDCiTsN8wKUfRJXmLaGe4rY6Rr+dIgD+R8+RZb29RhFatyuHB1h1oZbt6p
STXAv2SvZhPbfo9pmS3uG6XG4mUzitycFX1RudWtUVpOsZLaEcF6K9rmRyxxLM32
lhrBrQ+asziZFCHM+Uy1qqpIlCjbQu6A0NeR3lAbhS5k4PIXJe3wRd5dDCQ1fG9Z
P51tqLfqk6Fz0AXXFKoljp93q2pErkfpKll4mDCzES0NwCXNENtsEM0182gtb8wN
ZYTpfZfTldj3M3KUJrdub9tdiZLVSHT28nVrqJMrn29fhSNmMtdh2ghydeC8X2Ev
59uS3H2q2NbvIrx5DeqljnH9Fj1/mxSbQRFwtLQLcrTCb3sIHISCVPQRloUnVbyf
FmljZcCaFrpoagxblYJAYzoxnzGjsp83oeVaQZdyfDl61aXPOZOmQbDbJASo4TPZ
LQUUe4VoE2bCCiheV+Z/gl7M4D+WEkRMsXG3H5cG8jULGwxbcnuUb4UJCd4XZNfm
6meDRp4B+YwFVHC3qZwcCMJ26VT/kAjCGlNPNIktDovJ6T6PM4Q9TCwjdoKvJHXa
65cW9LqOX7ZfuATab61qjbFlNEE/1YnWoT6yEfi14YN+P29nKgH47UWpC+A63uWe
pPav/6abngcjRsMAufgCrWozH9g1aX2WHI7oi0LvYJAQ2KiHT447xG+M/4im5AHx
1GmVcv/py5S+1iejmZ/hu8f6FGrHojb161+xI1zslvVekOodbaBwwJ4sSenXHgIR
f//L5YQ2110+ajJaHWQSraUcWxqXWFcBHcPAEQa7a2gooaGRQsm0Zk3WabLPnk5N
z8sISUXklmWsItxWz/EYqbWyLjaBGF72HrD03RMLCXbIk9cAcVtD5ocnCPyhxlFN
vSxksSwk53YpA0wPK46CkxvOQB5ljbPpMonOwutIqakXBLE4ca9S4Ised34nScwL
9mRshD72T4vLCwNEfKaQ5HpA+vO7X8TDeKhxhVUCoviJZDFku26LAsdihPrkxbYB
Gfo8LwteH1Xe2ou9sp39q2ieR3q4Y5+EO0TC4ysEq/yyvMjZSOenAyehcfSk4n6y
akzMQuzUgHYkjDvqmSLjYIDSk3kMEnXffC+Z/MhS7OlOSEoEsDIh4LMacBJYeigp
WfrNpsfkH0sN9I2eBPmZ09gAJLn6U6Hlnav7gKJQvE0ISokNVYo+9KOcxlBYIBCv
GAildbTihCrP3Jane6rK77QNnytTMBJL4ohrg17xKrRvwEesiLtrfixPzBvPSINg
Nww8Xrvk5HbId64BOx9aGVsHhJuPBMA08oIQz7tqI0ZAGYwcv1riLzPd/r1t4YqS
SSJUL4FLTOKw1DKASm31D3n+Z9i2S7vRKR5Ikx1jnh5ZfU+jC+2H2IcwYSfJ8b8b
WM0MC1c9FenPNDHcYgBwNUgSAlUWNCB290LKFy/0BcvdnUNfvPW15WIDHZr5rumR
Gb/LF5EV590N1LpHT7mzX+DVgFGhGIXn64HCXSfB6lNbcZKCZweWkDXawVQvoR+Y
BWPq7TrfywCh5WWak30zKSC7EwDLfP5eKQ5Squp6HAlb6m3zzwyxy5HR8VYT0zDB
UTcT9EjRyD+40Rc9HRVmC/WE5yTK9zGUdX3T9tzqAggCFSdSvg6Y9x7YAZjrvH+w
L20+wtq+nqB2v9OU4U4sIJAPRL+KOPqu2uJ2ijtoIR2d/nOeUIjbOLUy+Hk54Z15
52rzY+P9EJsPn8UFullA2dDLjckDnFFkstejPCP73PdyS2gbuZRnXTIm9ECTF6xY
kNR4FnLfCmoiLAOFknDtu0OoStbLHA9ytuMhdAdMkxP7JUuVzpPO85aAmp7XeLs1
f5lJW+JdqA/hw7OMpI7Shu0ABv5znaoUoxz1w0YHUaKTwNdzPqH6LI36Wz5ayQp+
gy2K0fIXOFMppRqx5JtU/d4oHT/N0p51dEI6UrC0S2MWzf8qEPGlOstYgu0MzzDc
NNxeDHQk6jmi4fl101tDH7T++aM2DUbhx8cF1dz54VYAnuAXLm1120/95aI5Dh+o
aRPzIQtkOVH93ExX5ad3m4ZOEYRO/110HsGXRynVWea5DXfOdbe6dPuCCzRkdwYq
2kcI0qlL8gh7OHW46UXMMrzJL2UfcBp4UfbtX4hCCYVcZi/TrZUn9Nqg1vgh/lyB
nOQpOZ8oLA/DVsoPCl9VXqV6toDtfulPdgnp4pokhhKlDxPwVcqMhBMXmS6VtUZk
kZoAiV74E0l6e+9cWE3jITcZ273ovqdOIyKC4/WDq52fDg6UOHc5CijFBzqSZRlE
5FelicBIB4+Qc2aBqxqXpc/TFH11HqGd7c8fczOTPhkA7M1JncUlZSWATZEHSl50
yYaNtSUw7HoV68M/C8F1ENTPuYGtVWWtw/h/2kvrKkcy4hFwrxM8tk3P4yDyVswN
3ncZdJFGxcgY716QkreRUOsGVIxZp3UUEXNWwoDIMVIPwjqnWaU+xRkfIS8Z9F04
EaNKdsploBoy6vQtqnYqHO0FcUJ6AfudaM0JeuO7UvZaoIWvoMmN0in7GPVGxyqE
IQAAutUWnu9H2mDoUgbJFE9ORtFfF0lvihDrO00C1YEEaID4lQ7ozVgTnTnRdWJt
ZSsbikb3GkUQErKNhuHspt2XklRRVd7bBvkve/ZUEPGwd8NV2uRJRdZE67lSQshA
bQUnoEOpsZt/23By3Jr1tlUcpFBH4Js6T/IEa4+Mkf8sjPOAYiVll5n3sJdfLbaS
YQnlnIrzhdUTMhDaOL0xTjYj6BqIBvBFVd7vYHzvQE+QKM5oOsp9o9hRKvNERJpS
8O2Ref8mx73Svpb2YM+YgUrcHAXBTaLj7+BPb+lB3XARn9VXmLeZcQ86etHDvCM3
3PQEUYPGo5OOIDFYfu2flz96Ztfuj0KXJTHWtrddunXutuTDcN1Vs8utbUfxNLOZ
QsUau07LUXI4ocMcIEwRBYsuNrKKoVzAgnKO9iksY7UfZloDwNNDvKoh/qAXw6uU
B4gfMOllPbeob2L8bWt6o06cvpJIDdH6b7nEY975SHArRRL46hvlFkG4Nd6GuWRm
W3/YihdhgV4u5oqGaRRE5jMnGSIGKe2L7zoYbVRGPQaji40vu7Qu0tFj9JnUR2Oc
mKoYwAz9rbcgVcSZd3+3uHQEyhxR3805/D5fd7qZsP2FgG36K7RPqUiJ6TgDAwhc
Ic893PVT9NKQHJDzda5DvQGS6MEwv3dbbUB7UFIz/yQpUV7C4eja5697NfWat6xy
j1ucrejpla+ZJ2RYcjzkQsRuJHplwXxVz45TGOj/nuRmX+h0SiHR3zV1hO+2ANRN
UBnyAN52JHPNIcWr0+EF+jIx2DJj5FBkmEFuqeYpy0Jbh50shBllDxRSQpB1HP1l
dznsHmBSgeTthgGiWFx4ZQH+b3EtEzJ82CpGE9zlamoMMVUer6vIpNjmHzB5g8E0
yVeedhlS9RZVglI6Gus3BWJ4zcTdkN71tow1kkB8H+6uH92XT6cCnalkADhIXuGd
52BpyZC7jtXnexlXYT2gikc0UTde246zM8ZmZfvKyx/5xpllELDAh+WQormvltxB
ghe3+Kc9unhcHV/yyZQgdgXJN3HWa3J5i/cIbm3MiEcU7YjjUOHEMw0cHwU8jvY5
CTNQpCwntDS6SNG1LzqnDrYeeSVI1isvNPtofUGGKolIanNVwNuYXS0ulta53Ie1
usf1/9xtgPPw8fDryNsFOj9hPmybgfgjTZKZEaQlhUVx3cpGoVNvCzx1ioEh0TUk
8B3K7y3YTtekv3t6aa/snX55Y4kqFPw4IRbjcOIGyu4FHRMTBonnwFzEjfnQJD0W
2i0oGFN1yZmjDaIfuytoJLE8xIvIhpkBE8aeIfUHjIui3hsF+6PbnBHtZnXOyei+
hRVZmFgnb95JBDnCiSUIj8jRqda3VK+ve6v/6Ral+TJGp4dJBLvZrHIOrIEgMFVD
cbuLUZsK5VnanE3SoYrkZ/dFVYiCHuzu2SnSHqO7dtbnLoAjHHpPAw6HEFLdQnLm
OAC3UA3TY5yiWB/D68GrEJK/8OD/jmaEREFWC7xa+6dceEEqGvEL0SO7oHb7UpUh
+iPdNiU/mdHvclFknPXAJZ/g0u4rwN9YlowObuYCOO7EikL7npVuyrxZ14CUw0Vq
dY3ybG5marZl+Ae77vAORxbNGnteXe4sqnl2tbHgGN1/V/2xUoW4DzFIXzfN2Nhs
YcF2ZZJNSWIsGYFoV2yz2oJ69ZdvZ3J+n9VFEtldYSjQc+0gteUOGaYbMaPjCwmP
HgmOHmHJ+JWX/33skr/GDsDNXxXNDk77Wz1Nj1CqK1/4hI6yhwd8lfd8WgjEbTy7
IzeZQbcUCrM//Ye1KS/ltXV8t6SV+md/ybn0G5rNH8LfqiXcsbgK6D8xJdHkD1dW
4ggAEupwDqop/kChdbif/0iCeRMrg3yENybr9IZngN7miBamb9OCEl6P7u2sBN2N
yAwOT0Iy7VdxMCBLPLMLNYpvoZqb2vlU+2wCPVoUUMrKUbofoYH78YfPpdG/cjY4
bEGPBAL/jJEYvAmccz+No2fxg6bJhNMWifII+YmAb3e60QhOESPPRXd8q9X/inmp
nJp9sELzwpfuDQ92x3BcX2c4PgH0fqkT/Lf41ueam+bfPbpnBcZQoiG9nuHhUqa0
CLYSMgZ8HtOtKsrqCLi9j5bgK+vQaNCtWDkY4zjumOcRfgHquOLF1zC8LzlwFxLc
OEYKcmJcYVwBg4Ca+KhVYrH2R3ZUzJ8D6JzsrCMEVWgvtqn3lkTsMAsBxVcmVJwb
R1Q/Cdn1tieo3eqTWNlp60dkZNl6369/IYS1qIppaV5zK8N7gbMbKRCktmc4f4Z8
X0RU099vvzJSA14cmOKO/CFJXb8XVy+ShdQ8118nxQTRZG+0/d6w5btimEhswDVZ
s1fOxa64drf1TVB5b311yej+ft+c86GxBaxh3FdED7N9YQav9y0ieQhNpkLwCMYk
HgS1PYcgYj+Aal7TY25+GY3SDVN+a2yGnOF691HmQi/gb/MrMtc0ow0s4kPI5rS1
hIJc3/0uOXxlzlQi4OO1BBhAnmqokKVbaGmXBDwxJC+mOocQEXa8A8yR1UDvupRP
+sVHsmA0CMDeAnFR3f+MqbE0crQKwOqmAR9A0dlk5g/uTZomIDJmvweQRdWkeHdF
49XSM8NW7iHoa2IMEPOvoC+CvvUuwFsYTUJIwWFdG3w3eyhgWJfRWWzvOyX8HKXf
u0kK9TDIh93Z8VO4HcwltY15nl2fLDC1b9/uBqMzTYiviJIIshiIXMCowKGYdJJ/
Jrdy6Zxv1ktz7dQBZdqkccZA2U+Ivk8m692natcDpg6ejE0wAm2oaUfYZnT/QwsM
QrL7zL5UPclRyt1rzuwy6EtBmzKv3uVi+Hg2H1hhEnwPPmuB9kbQnnDFoaa8845X
ITTihQyUaX7BJH1rkp3lV4hNjZLctEn+o/f8spn0RmufPN7MO+8sx0w3sRYmEUJQ
qnmc4K7p+WlcjITI2igsuOdIO5IOaoa+rc9EPF7Wres7NDLaJd0hyyk5Phs3HWvs
VG+3XzGQru6SWylySEetXnpg6dEO+XiMhltpf4q+SBaG+29Mm8qSRsEnht8EO6qU
aV9v3roU3Z7I34Yi1DQ4vNUEcqDDEQLPE8E8/XXNkXOa64PpfRGVS6+x6g5mYnPQ
fOxHidB2gwvOvLqIKcoO1mXtL2hH1BUBS2NK2yg+t4JtckE7sl9Cvtl5BHMqwz+B
ISrqy/1q72f8aSBSKm7uM9TjQzkFo6yxJcDdDP61pVyKTa0qLC6VoVMX2dGoVQYf
SKX4qPwvtXSkKbmlXmFWbr1qd/Drex1hc4j7NGrMW646HFMzJJ4o70UMGjg/Mo2t
dwPHcpreCBNZcyqEx6yQN3PEESYIgVQisNDL1xdlDE4nTEJBpUGixMDbssmFvg1Y
nUXWoefUVi7b6buhL3M1YkRc6GSBAWFvuGUEYhufIKqhPesxQpXAGJGMeUegSdo2
Lii3qkXrBa5acXvU/JzoNWw+yCZVcnmJ4KeZBnfJkMhZeKYI1qZSq7QpOokVe25y
rmXOSSKT0B/eduFVeoOUB3yB9W2wvrnl9Xsh1kGb3F4PUjeviJS2oCTfFK669zph
fJYkXbppUUdIJ3Syf+BFJhJtGdRz3fFH1VCiEOj984zxAIcwAzUeg4BfuB8qm30L
89o9ByieCOTuiDUMgz0NEIHuOJdb0g1pbOcnU8FlfnhYf14tUQtvMJDFqBzbiXGB
+vS+qHdnr/TD3CcFVRVupVno81JcBcuJ0J4PvasDlx4VTEYFa9IF5KAAtWOGAXc7
d9YNpaWcuuyrjR51cbIzNZiGAc2vypQgHJI6EtsFp00kgLapQL8Uyv5jIArdvEd4
Js7MvJgWMKFUfdE2v/Pg8K5Be9tBuEGQo6H/SC3NfJ+2vEMGEtPwJWn3KWZpA1Be
lnK819sCHIkyxENU5NX1LPmcgz8C/sWr/YU80QFVWM3oKOBmyxRGo5Jt46XVR2wk
DQ6tUEMZzx0JSMvhGe/1N0RJEZ1kukDw9rfczCP5Vj/u90mc6q7BOJ7PEFBbh+NL
YmHwy1dRz5NFYsXj26tLN10tLvTf3tXm1ObhAjn3n9VeepYgCLmIrQmrJOnDL5Pu
8AH7JtUu89vVxD4Krw1lhBJ0tLc4+sAMk5bIq0yPul/v64DD2YyXT6jk5rIr0mdS
B745n5tRVWFl7NJ7DMQpIuYdft0AhC6zDna71L07CqWkri7CQa1p6hzBAurJJq2A
FGPCP/eMfoA27WIGTQgiVQkfKuzFG5Xgzc2pOGLgbpYmjnCrbsYPau/eqwTkHZbr
Pt7ZBE9myOrxTnmeq1y9X0pQWIRFolXxGSr4eJB391/DGM7yUn8Y6ZsQTh0XU1zX
Vkzk4vw1JWN62hoCk3BC8apuTw9KNrTXbZhM8pY7tI/5y0zOfdXsZo2xLGPSiNsE
OhuO9Bp9SS748sepguz1PRbdHxpWG/26/feI+UvCOa2hyoMLRBMZDZAfr82xnw/f
knqH12BftE+rKL4cqXJw8LmP6qrXnLIswzIJe7BO2jJAtCvcUKZvRmagShE0ygb7
ICPbtb0XCDEebKezRENvmpoODuie8Vr/l81zg0fS5xXQIyEQ+h2IzvHiTgalYjaD
Z4vMwLdxj8EikTJAaQBgr3wDtnHNMOKQEfLornCDlN/PU+I7JD2m6uMDgo9kbrv4
dd+7nqto1q27Tcfs7txmPOEfpNXqPaZu+8gnmfPlW2r8Ynh8aHssh6ont/R/IAV8
SkVVy1q+uxMgCaBpR4Lsuww/LGxazZWMPJQHzcBVcZb3MRuxHiXnT3rf+bOJJheY
N48N8sNaQyxUMA40mE7Uyk7iUSejrwdtgmV1EgLN3sblt9VbtFxItuS5aCOCscS/
Pi9zH/7FAEdW+oNwddHoYSK0B7RXjynQkeLnJC7PKdKFOwd5raoyRsmYxi7x6+7W
dWxenno0vD1L4fBDFWjvsml3ikiqpkoJ+yGFQdpvfZc8nvMSpXgyWKAn/g7zFfrb
mJwDgf5/BzSOout66Pg2limOojtF2R095RqLTwPuzoYCDY9qlrt6DJXq5siaq/vL
uVOTXx503CdJgpbOX84ovvrEtfhT9AHPykXGbcygWJifEGdy7TKF+UGXGIZ4oLlV
L+Dekaj9SHZRMyDItOjMJ/HOImvbJTCs0IEiRkIqdbueM7RTPYvPILr5HdqvC1NB
B7r4h64gYdIUrW98vq6sax4+H61FVQSS9Gi3jTYjF/VpRx7Lvv5A9HwY8+dUVZ1O
fdyR4T8xbU7WxUdSrZifT7p8saR23kb3WXhIM7Qo68mAMOTMq7RkQD8qyyC7P07r
Vu7ChIRGBJnkes68INO0lfyUBZ3nGiUfQ2ejtAAArAVpNTlOc7hxuHrxBltgtGj3
5TsfTPhmV2Uj52SRLvPwKzr/b29RHTen6QU7dNwH1xbsdA4u/KLzpHEIBjTtjOx0
IhIr0+KwJvcXwUJhmMUhW4PIKNMaaKBPTA5rDy3wkgllYn0TjcpVPQTD+oIEc7Mj
zwsmebBmgjiot15L3sV9XOrU1HtPcdl7275MstMemmSLIIQey/VddV6DhoxUD0Jd
FRP1yl0EPlBKS6fpk2nnJ2AuCAYeb14tk3IiXsTfmEnaK4urhLDRV5m8O7i38L4W
T/5FASS0wOccFmHGYAe3enEvSWApnbbmFgsSi8rqyiYW8YFwqgUYg9J1n5oXIbW8
rzAAEiBqA4HK72+kcbhOKeQXITnrI7bEH+PwZ8msnMuIolJMHq+ye0yJaJVqytqW
ZbGZNvYxNEiHiAeP077qMbJVyDmSogBd0/jUgPDrp8gcrtJxL/n793QoENoOdkyT
QgUml4d1G90nYwQjbydMom4anoRKz3LV8rGiTqCUcHA5UunpgiFqsG//5FVArbHq
GbYn0vo9Cdhs6c2d3xw+SdzPaT6mkcIme7fhA2bxl9cRhbfCgeBHarzMXd4bQ83e
NpyCypRiicexkmso5PI9T6LU6kkVSDiCXG8g124uV030AO1Dekgb8S9zyBQrEr6X
hU5+/GTq70+O6HB9NSzZnG2u+9cGd/PGwUhimhE0U6nnNfZdDmHnZht51T9TACGq
A2CsYG4J7It8mgLzlTIbwdaE2Pg0rmEG6XFbLq4M99z82zKsPXC/yzutN92BM01R
QyDxmjLjxCpsLyQ+J/fD6QZRj0QvTNmb4MElHhM8PY1/mz56fBQcsw2l+f6Wvmbq
NHjomplEihspCHeA49OtKM7kxsm5XnQQc2XzD4TozKoYmLb0p+zpwKHo5hWdP3km
AUUVWHp+sJNYaR6V3gQxsC85WgkEVgKNVeiXCx4q0kVIN3NyUKg3rxm1dWwvjzMB
AfU7CczdcxIGqH1SM9+DaUmRgRSHDC6+3tFsDlqhAfN5AM7C4sYSj0lsMFKbLkzF
WmFnAm4A9rXWfDOd4u3YxTWtKkrUvfXe5e/njf1WhyRf5rn4r1wvxman+Te2aTri
ykC0XK9/seRF4Ouu2fY5uveN2Sdv6IPcrtof1XimOPLr51GpDx34lczrEoMYc3WY
Ur+SgSRg31MfR/Se1LzCC3vOvv+kfhenOx2EwxCkmSY9Qx3r6mQcCW8pHIgUKboT
uszZ6NbZrF6n9jQ+j+YGWpSUnCo/OGWF/kspj/USWQVqqb2OJ2OK0KBA4/aETkdo
D3WBw6k26rLoa/t474XskXNt5WC/aDvDiXfTcljkFS+kjS5nmkYfH5mEG03MY+Hr
d3Fl6ZbXeWgQ6JlriGD3TKryS6cbb7KxGBshOJ+/TW/hUYinkU7OTwDsXWf4mKOI
RjyDwDfrFS7YsEax87Gb5NeFHfz7/WoxMD8qezOXcBQcg91d4FsemXQMKgL316R4
GtqP9/kwMFIq2jSxhAd/rQjpJjjDr00miof7WX7pZ4icpt1AiYFioiLGVY3RoJY1
j7cd+HK4w4lBSzU0J7SlZjCI+FCXdupXV0QwGhQI0gZNkPnz4xwOf+IFPrpSPzv8
Dz8S/EFWqVJUCVrL/ikWsQnYz6skrMP6gwmUQ/eU/wyni1VYpZzZBQ8D5daB9NbD
l2+i2BUUK7bydomT09X8FbUvQSkiyDk7gJeI/uhMeOghLD0JlV1gO14qwMsp7NZl
UbdKDQtzsvOi2MGpE24+BypBhvjohP9dZyWVoZPsUf8p24nq4pGptiY+kAZ0i4+Y
vsnEM5T84go8DRpXDJfzg1/ZFTNqztkdsqDHo7AyRsUUN1B8QR4BO5NKTiCmrkBR
5lXGqKfPe9Mv90ebDaLxtJ7u3q8G2L+GjdHX/WHXLvhPGZFb6MEHYvdsuPNkOaxi
qd0wEZUd5EXsRch6eanJZxDKu6+o/16szl2Q4JemJcGBfG584HSJl0Mc31K5Oli9
sq5z4EKqKHLG+l3q9wfuS07hzuI79MxYjm+kMIhM5EDKzM5zSpAo+At3zyEWXfsI
kuM2HRI52RC3vmMozmjNAfFuv7q3zwcSUOtq+/nyYw25FKWgYq9SRKxEt9GQRucQ
PRFi88VlTTbjlx3WJhx4+lO8/cldaSUsNCzsOF5pOS5ukIycq5nwLMwAJ8QBYRCC
A2Rls7BJlxDZN/aO+oGs5amCkO2asOTHm312K6Sx5ZD5hJyKoZ+NxFj8IsI0EVti
0Czo6vHjhMBjo7NSgTzErM8dWwle32bgj0eN2N7OZ6DQghPloFQCbTdJ267l9a5c
B3u6vMpItPysbEqMDxKpS24IEBGg7firqWwArURB81P85gPACgkLZYIRg/M8JLHQ
Qyl1AIZOeWKY5r/0R6Ph32aVBZoivEu3xwv2xi0NtbXV1qANF9bKWR4Dc4PieIno
DfERw2fuEp6T6tlUT9CvwkmrRZHL5+goyrUYXrPmVTcO2F6j7ZCIsiAk+HpJ4Xjc
QbBPM0bK8+KNR2A7x1j4ckkgIYf+tarvMOgkw7CXmiPtTrG1nxoEhie24HGtoKaq
q+KDt0RBjgvkBa9J5TFgN9budXaccLxBeLerBFRCmovNaB/SRw3J9J0UAFPfZNBD
7mFWtAWftlUmjlJRX+b6lNAjjRNt8s2tXT9UVJOkOtGKtT1WQUzgqkNuVulow7Yy
19npNz9G9WruDC2/RZb0LD75XGw00zdmiiWvSXpObTuLR8P34SC18lz8jIMfLXkR
T4ccWpX3beZ+HOd2Y1P4POnwXJpsiqink19+qyceoU/qNZxOLu27V7xpzHHEyMVy
FE9Lqmb5htZNP9ssB05ts62Mc6N3aGBaaEsu9TKKSHf6jC7L4IIyjh0kuPlEIzFc
0kl+NnV/ZpgUxcRt59320TCeaNMKODIpt1Vc3+zu57r4K92kaiiq8v8U14QLGbEq
koSW7N6i/XU6qT+Kr7Y9fbX/7SGqYy8zBl/T50EI1AkGVt1s/r7YdTex5IEny+MA
SlB0xhfrC8ivCNAOn/J0uHtbk+gD9LOcgMtYTV6gBrtN38G0HAtVACQr5m32CXiW
cJATEn33c+DI+Ly/3K9jQOh9AyI2kVGkiEjEMcB0VshGs5X880Eh/BSlU3VMTsyB
bDHpLGrfF9wCq9BBeU1pBDh9syKdDK5HlVTXfgFYB456c2eVkEKInXC0xu9HHQs/
punSGjauQM+P6N3qp8GTC+ccvRh//vFtN3q6GBEfPFMlkQihgxsQDTe7FnuxWaMW
AYo8qn/uhFuO3beUU+9eNumm7zrWB0w4MB63BuMthLAqinwMQN7HSBfqFavN/f98
5pFTzn8UxiK4lzQjI6WQB+9zoxn8j0e3NnH7acLWKm3ufdZCYiWTaZGKu4OLFTsq
dT6etMauVT+U3O+6sAybqAPllhHaltBTA3PKRHx6IWbHul42bCkn1Uq2p/ASRQWB
OOvww26Vrgp1DABTxngeW2uMXrZ/fLsgzh663Yd8E7JFSwyg0JlufaMOaI1SGuHQ
oTsyX60or9xC1NosrDKnB1lt3JG6xRssP7CMpJimwa7dGaZMQOdwA22aVOBpL6N9
SNqK5GrllOUJkRrQeQZcdDA2HQcHJxuNr59W4F2AdMO1Of8w5sKYaXWM+I8V1bIM
3ADn6DP/K6LrBfMO6FZxxxSW3aBstV+VEMtgWvj983LeCQQhJkXFYqEUjeDFj2ku
P4Uwviwq6251r40AkHrrQ5DtWOiYff87FUZagSvYqkP1H2DpaIJVzKaJTSCVGnla
IU29BZXpIaDihiOEUX6ViabVn6BJUkJl3KRyNR2TaxDW7CBglZVxBmAaL13y1FTS
Q5YfEa8mpyiHBP196tt9dTKpclDC0gCptrcNHRbYUJaIa8odmuRnRJCe9M9sn2hR
OUu22DaWDGlE+oWLeHyxPAmJ8Am4Re6NBG+171BnL4daSqC8zr2GKbGb42l6hLh0
N2KQKkLunJkKRk0OxFgQ0ZHCJwtauxkDbtCdSZSszKiCSXDpZFQlgFLBGiR1YPhy
nyYnOHitcMJrhmjkprFx9BU1a7+djXQLl2fNpc9iFDBJ+f3Sd/ITLyTHGbkVKSDy
Ds5TxTXfUL3rebyqDVBe3nPJmdcQGTZ5nPG2OJE8m2+552VCI8JjGpiuUh4xqKS3
Zp5Fm2DgvI+Y1vwGvQe7dY15A32hoWPQcd7S+NrOLecGPr7YpTo1KmqNx7aI+hSx
e5EbNPdCTeabPY8i8lkcvHhLgZzpDCQpX8sKsNo52GsX7lKC0N1RHI/51hc/op6J
jdpBdQw6WyqBiCHbVuRkwnxWVtDFAOr8yTFD4ap2in/eTGrOjYTI6e4K2ReM7XcR
SDwF+M55pJsvzhj0wVG3jQIFL8pwO8zxAgd0hCPV68DH2qmnQyeT0yAhJZFzJklU
JvUYa2vd9SLYNGMgCBmfQFIHhKeaFoMxda0mhJZXRj21vsHlOU0RjqWb58ZJ2uxS
VYLuAlZ9C1+G1hKEu8cZ9oIjCS4euepWlJxk1OPpyeGRixTtB9iRMVQKmcNS88Qz
g8NhX4Ibj0xjPcD50AYBoOLio9xVFGVS/fmpsd7ucNc99NsHRcGYGArkhztTy7Y8
wzh59HVlYKir62tM69GwKc5edM6fqtwWeep0L7dbgP4Z2HY0FxDvfKNbWzMC4wIS
FZU9S0kmNnAkim8y15+lJF1+RDZ/d884X0HJgdRzlppji+GUMzbdKwo3vlhRUaUG
gzo6S2WptvGQu7GDrUgTB0735Dg/+X+AAoPRf/xyKfDAmAm4iVQh0YvWtNHmz6r+
egCNcFtrVT2kUL4rnNknqfFYjrOeWBtaIJeY2u8N+SuQPzMbGgcPRjk5Rfclig8V
S9Hw4oieM6ZwbSJ0EdyzuXzGa+bbvO007C5NtksK0nFfJBumdZBME1nI5emG5NTK
YI1lHgdLN4RT5cdtZBbzo1X44H7Llh9Gjgsn7mJwAKg5U3tmKdjkOzBwqUWu4/qB
gLidKTwFBUFKcQD9jz1k/6oYy/YOOluIgdIAcF5QLBuEzyZTzeptpilqSW9NsMHt
a6fwexyDSBhOcr1ZU+MvfIzQAtPluTUq3RQFy/Bi1uMpeGaQplmy+O6Nm+ILy5Om
WAgQvMfxPEJzZra+4QE1cPFeldb+GdjFI7t9GcnKQZLTTAa4W8dyEU8Ya1vsykF9
k117CnujKusOImlhnNWrTnpTED26DJM2Uf0B7rNVFnmM0Q3BYS8r2cnSi2u9+o2m
VtCPSkI1zrCo9xx0yb4N0neH4AcoM0KqwfwHkHBO6Jy5nRMqYSh5b7mTf4PS/cTj
/1aD0HU/oX1yGzlAt/HoLNf8lhJE8y7QsSMnApvDqk/KXh1g0OBeA4rIh7vBCEfm
aKqJ+ZM1njx10jvuIz32YN2J2bF4nsAzWYgUWqhFSHnCMjhG3y/CwXK11LmaNsbz
o+vvIvt7OyIrfPgqsM3RYRPF2dPyyJj0MpGvJezOVYhzsFLcUHZJ4MySxkxHa2bj
zKI3encQOY/hGDbb3CUUDqhfoM1DHTJsmc+17Fm3TqgRXbxa3DPpXRticiHybivc
MIEQi8C0SDNS4Q8VvOr4RKLYm/iU/5QfiHXZPfwQTDMCh1fFPWEXF3OkmKfuF41b
N0e19Sl5HMez2CEq+ptMkzO29liuEn3tXu8zouws5P3vhIzpo6eVpGITqtfwG2yX
shHppXVqaFruCFuAqcxHIJaJhtOgcl4VARKF6/v6425T9/oKNEVwaEPDvV+lpqBz
DzsCtrXnQooVBzN74BycfWQfQioJV1fNFc9JvHbNrQ9TobqC8Lw8v7yYfeR/hSBs
w71gqTDkVtY7SP635ApupjCLjdN9mWJPhQ8owOOCuhsIkso5WWv0wBUYkNIoieFB
HviZVNtDZcpzG9UyYS+vz+0+ihf9PGdHxG8d4w3QAC7DOhPcineRl9giM+VQlz6B
DjksBqJ/gPOCpK2tfNZswOtwPW6q8Q/LcHwUjFUnD3IN8VxeHKJv9w9svhVXPKmX
yEa4xHFiODZxvlzE7BkwYPVomRV5bHHjjuhOHWJPzlsg236a+mYADn1toCWy1iDa
FOLSHOW/JDAAu5E3tiwmN+yACpO7T1ucIA0shJjog+gmgB5cLI8jwl86J0njaRjG
YR6a57jQ7Cn+QQJ16jWCmzDygHCrRZbGI5uiSBZvkYGeCP5Ihnww1RGd57O0E2aL
YZ72VBPUsC93Azi1iCOhggNIrcCYKtmhqgEm+auku2fJpdBsYXqIZo9OqPL346PG
jsM9HvedtDvnnmdiDn3ZyR4lXxxEhY4Mt30L5AkpUMVWIrSJWhgDg96/y3uPxe3K
+K9f69tEc/r/I6dELVSsQganrQIk4tetEsVw0ryEyg6tPW/KDG5jmlkmCMh7qu6/
yoHT8fuyLUv+sLTgGRxFlfEb1oDBl8krycm4eNrhWPknLhlNkPHKW166nBjQyqRr
i7JhKUdhNmXXWGwyDxAWUplQrp9ViVkyAsgEzkOmR7mO3iU/rjciepOi9rypRzRo
1k3/+DarzrfxcD1FVFLSBMT+Ra97PeDAWpS6WjvAAMtMirBN92VUA4Rfle0/D7Y3
cjDk8FCFDXLvNO/hb3au3TsYSJe325lUa8IUyCd0tORYC96zdUE/7umzzAjW9c/c
9Ucb+0w1jCxFRnjDa2YTBGsSoMCui2Uu8vFfXhWXRykGbLJpqA4poI5+zMxhR8wA
DKW0ArSzRHuG+RBhPDtiomMqQdM5NckdmjfsNjNmiemAld348hymmohWewXZVwwO
fnFzC1X6aqbzMV7X9AhSUniDTr+bgOgo6s7MibRTb7QIyv1DW7BvgGD6SQtu1Trj
Lp3izP/5TsgfLoDhmYO4dGy4Sj134wnFYU4YdnLHVe8yaLPFExyjWah4/XJfRHn3
nO3ljJkU48jbK3ZvTu8ZsWXJ1cgqBxDGs0B2OeI/OBCvzjyyu2WUku5RWiCYUy3x
jyom14DBYaamHA7gXA9ZcDw8kTb9p7cfd45Te8V+8QyqIJdLvvwwgo+5r5ltWK8Z
u1MYVNggeE+3TglhsBef13BkUjpEiAJzHPaYBEpThqTE0GTnWrbnNbEVink1xfgX
jvJEuhn5W5w5lUI7fTyMAUPYkwf/64fcA9ZF57g7f7jszKcpHgVHxH23yQhTsn1D
EdjsaKf0o82pasOTzrNYx2z3X6Mru6myTNFIGEmrQAoBzE7kH14BVFP0S7wKYVxC
bvOESEUVEllSpyZMuV86LG3eKBy8QqSsn4IvopFX1usZM13rJVltkShoRKNlPmak
932PFn4fLcoOzAue7BOyCranvZ1MtQV6veuDL8mJ2aLdeoL1t+mwBFNIRFIVWW/j
TANFt/5OWBJ5vW4tmSuJ2e87vlsJUOJ6l8BLukoj259f9DXNzKdIA9lVTIRk9rkL
pbg70IOfRxq/pqH7VNd3u5aBPlwVjT+GywbPPmFVKFs1L0lyO+IUp+x1NLiIfeA9
p4MkpTEyA+G1VeWhKQI2D2Za7yD9RFEivV+pA4KDIcUvbr6xxVCumzYKa0W77QqJ
sHoa4fOLRene3oSwLxp8/Bw3QQiW3PIWrh9ZzBmY+RPGq0dyj8xUi0MVEzLLSrk2
RATDpMc58Zi6W2UzhesmzxaprRX0zh7ugHun3MfO2C0HboZXlUPWIdOPfUVmNevQ
4KyfUVdC9LxDQ9NWt+v561Jiy3UPo4+xq9k4mtd+AHUAD0/x7PTgaVBFVqqZNDF9
MdQt7WTRjPf/fkywHd1VK6utKNQO6d8xvmuzPgKqSaqVcejJC4YqT0JpxewL1NA2
2ebfhYmsmfBH7G+5ABgyYN1DG+x1yR9NeOJexkeP5HlnStCh9ffWANwyfH2FFfTU
c3qwBgPqBEiy4hjcgaZXte5jRwK/V4Qm5QMmUNHm4PokgBCY12rGn3y/RB17uuBP
znicbLS+ty4fgqGf2pYxE6Nt2N+WxZJ/bYvInjoc1MOfRJBp2NDRTxo/cdQkV1ZF
qydQBUMNiAnSBycCU3fn9IVWUC+ZkJ0WT4BLpXVF/5D0yDaIYzEDfWdvpr/zkX5i
bkLnazUCgEjb0UUO7YwhqnESMkEzYG78AKcmCxIn9UGD4cAF5WnYDH7B8LYr3IsR
oOnKKDxYLWdo7a1z2flYCb0Jo0qOZryoVcqkB4fP3WgDj5BC0ajQ8RgrgSTGNi05
xaZa3HJN5/aWB102qB4O2ryQbARB8vw177Mew6ijAu9MCw+3bZW751CScDGhRmZS
+FWFizwHeaq0OQqX80s5bENRBWH0KROqh2vkT0xnQ4xmhwcGGemqUDlEsx8e3wOn
20u3Tak/uaob9tTz/PdMvAyt7SRdusCuZMYT1YUmYktyaEQzLjQad3h/pRGGcZv3
1YlJ3bhCLCWGnMPlkYOwpypRrkpfNp7jc7oyCOcf7RcI0WpJq4LM/N9GEJDIsTjP
thTm0JBhHIZRd8Oo6smfsAgVwYp2fNiIyo+Xe1BRpUG3klzId4HBzpMixvwYhGPr
/1IsMHuoRusmIfUe4Lxdpq6jZ6b5OniVm5Jl8T7Libb6U8MbE9Jruclml+7oTQdk
EKyKm6suKx0sTz60QZYZ6OavyKiUO2ttlegvUxOxnCin7KmnvjCnMleNIj0vp37g
hmEU1KG0EV//nV0PC4i/J2Rd3aPIYtRt6GQY3hkqIQ8nQ+BOYnuj1lbOv/Ht+YiW
5qYQFLmLYPmmN0avbvcQefmWdS2ozx3Uyy3lNWGWaQvn/cn+du6TYKmcFHSyHHsh
pDvBlnsd0L00e+BV9kDxm9XSK93qlrz4/ee6hi3OoObkDx1qyLn1NihU/zlNoBSs
DSTVGburfgYLnBmT/gjPL0Cdf1b/+JzaAF5aQakde94p+zRkdRFW4Bo1UY0Y6p45
0XNgrDI59ZND7PVJpe0Zf3ZiDiDkVkC12ScrQHoybrDGwGC622pGhW3+GO/7YT4V
96urDgQTCDgocnMwFLkLnI72gKzDsQggfxdfvtvxs+/nrShysp9ENahf7uXZGw0W
8KBfbagmVM0B+aeqqxmnzpDrq3gZp4PsNF0zpHYuho1RI86UP77seZUAganj3Woc
fnNNRir48oTbtA/j8jz1kg4MNxW1Z9tNSzuAK0o9IgUUf+XvpA8dBKIKVUFKAzk3
bUdP5hsZs0NsieQz/UZa9l0iFYtdqz405KOumT+m/jb/PCeV8Ki6HWIK5K7pFZte
uBu0IBujRSaarw1JT6abTDVI6CW4bIC8QJbgzmfaueVG6Su3QOoIDNIqXJRKnwK1
rmpAj4ZO/pEfCWWbXsI1XQA4/PKgZNW7JQD/k2mEXhaeVqVv85kb/JFtyK/HEtt8
u/XPjbnosrmQCe8CMn5Y5nU+ajyioytXBAip+R7XCKdo1VtHScOmcK8jTeV0Tp4h
62HAktB7M7EXIl3QAh0aqUvG7ntYf7FJbJ7qE8rdS17TuRYcPP/9mlBzXTFBw0sG
oUCW1xUzjvLhZhuDF8EJbVTyuVWxR2C1Pp3ddBBPtuKpKxD7bMC4ziIxs0Y9baew
dfBJe9FGc9p9fsmn90gR13SimwWwJ9az4p5uz9EPMCzD142YyrQEgmIGVKfbggTi
csbUfBY+a/p0fomItfDiiEe1E+jfKeqv7jEnn0aNWFEnrY5Bqq1GNCoBieDoEFVZ
e/PB2v5HWX6+4eRZOk2PAUVYTeAJoTF5kl6I67ZjmTx3MIwkoWZDxDTcAbJCDNSI
kmceCiEpiBBblgERbFgcWNZTNvsndeI1KW7gSIjqdaRTfs92C8uG7nmgO+vtJ3tQ
feIQhFblabMO34rcXBHlZMvw1Prm4vNcr6avqXspBC7DSdvlmJapd1AwhRv6L4UU
3pziVMkR+LHGPzJEbJmJJZESSQ41HGLcR9Fgu2p8MyYHnXyN/OXgF+5l6FS5lZZT
CTZUnF37fgSkyrZzAgEuMrXmJ0Vw7O3redKiLfgZm+/OgD3eEea7rN/ZdRD3I7NA
OSikDEemTfd2EZzaBcG/1/KJ5pMtBYoXD379qZ/OKu3T7Kd2ji1/BCjMERofYFwa
TdRrtMbXLODWnesTjugNhqF9yRWmVdie3AS6u7boa5PWeS1Gu7V+fk06RBNa2gOp
tpojDv71fipTIO7LIk5ybf+i6ItkD3uLxPo06/wfTGrvi6TsHLlDVHATxYCdABGI
gFdjpkS9EJ5br8Mi63+pOiiAxySd9WW9pg1n1ZFkrHoiZXLdFfmzoFQuwEY5BGbH
6dQDonExKDhfvaOxMkvcG4ygeQg458yp3MnaKxr7y5nSvtv+9h/qNEiUQ2Z2PvUK
1XMuIm+ShkhNPKAv4sqlZoUz+4AqpWmaLr0s+HGa2UUsqcM2fR68vYtlF4SakubZ
vmYpqw0mFPzejuNXxNIkH4lpnCid5IcV6XJ4vQtv2dDF7h6iax9keDHBCs7IvqDO
2UGthU1TJJimBWR1YE9ZEvZlqpXr2kBPa+b9hQrT09kB0vahH4n8PGbztQ/lzZ/C
uCwWRD7i5scfOsDWoRekDcNQ881XjufNTkQ5xQWAz1TqUDjOW2qB+GgdGLJ9XBWD
WPBeR19+ioPHwc90LPyVZeXkSOOEA8uEOCaKMKQkhzdV8o5+ioIv4SZ/g3nB0Cse
r/yzZyP55JWQEvJU3Gat0heAucNH0PgU/o+BP0qSDkJzNVFQunlmn3y6DfyXYj+J
jmiRl/JQewOD3AObt6X856PjbtKB/+mUrV5NY56wuVzCJ/22pED9DkX6LCvzXn9R
itMjbTHxaOs2QH3jm6iFo6pAeopGhsPeRhSRso6T2XJ9duoj6sUNdvqHcTomd7eW
EnfLzZUzO2E5lLi8XBc4sI5N2mCLmAnIyvow/uZrzuPfEIdj2yEvHi11ECfiir+j
ZXD8pgV4XL8XZuFxF3ZoVexdcZvjowEXXpaexGeyqIrPgJEZFyupg8wJQ17YFepQ
C3LrFAp0WxmErTqeo5JSi6VH1mKo89Jq+uwQuIIlSDcmYTDta4rhkFcEKfKbHU6W
ZzTFXQ+4VRLwgGARKvy9y/Vn0IUzohrePGaeyBelBj1SV1d1ovv21HgjLrpPotlQ
bYYS1/tlt77GBVOVbWhMK3K6FsPTdk1Ocl3YmzET4UuyoDiLstZEYEazU/1EQeen
tCbTUhrqI4g+MadTWplXHOrlYTGsO6HdMvujGdqPs5m22sjMgHB4f89mbmR+VMHX
5xlCFsfkvM4y28aoCoBBWc/P97neVwZKRNDwuDVpeX1gJep35WGKvRZduy3fcEBr
wVzcXOzBPVK18vU+jeOBYzf4x2nKsWNoBKWTGIa/zumgzz23y2Ijat3w8alODI2Z
PgWuOvY5tMKJOMKAuZcpDha8NcpKa0GHNNh2SGgrURlgY6FGaEJ2uOtcfbIggzLA
mX9ZZLsMItpE+WqISSuSJAzYwtHEilMNMFho9pT4IEbxPxi/uuJFVA8C+vLAPsng
hTlXN8GWbzRDscIl3mo/epneoWo7vSMW+nVCUUIdKzzdE9CHvqKtLo8tnEJzipr3
uV/fAbsEXt4AureWrO5GyT4pgLHYOCMjnwALcP23lIwW12r54jPewh3/Gkclj8Gd
CQKFAbByCwsnl9c/2DIsSbKclxmaOCS1olawT9eAjujm9GDoom7o8kgH0flqeO32
b2wT6QFvQbnMlYOfcy2Jq3pIug7v1z4tG/6t5wa6wC/9Tfx9dHjMIodwIhuNCY1w
NsdMsnWY/7kUThb6sY8wpIBf4WJqj+cehLwos//woRYIXN403GZ6JPZTs9u2voPr
c2iVaVumjaSwrmOMMxdVy7V/eJ1HbAJ2TTtZCgSVNYHlLjVIwqUSAZpV+ulU7w18
3J9B3aZDsltYDUCVFMbdhcnu90vQ2J8jXq7bqzn3eFUM5so49lMZLp99Jb9gevjX
9Sf1tMWQpzS0b/X85vfBkieCWpw6E6Li3RsKxu9JaW01jwQbIYjVB9/CUf0fWoP3
nMEYLuI4r7z/tg3gpFTDfYDNVyFsARQfySGgIFhpaEpm0JpYw2N7D683l1xg1C3T
LOUxM5wu7vKj0wGw9IuHB7dnvFtA03uFQ2zDjtgyoPXAIS0m+oZwvNoODio7+LA4
vqch3CsUn8x5qgCx2W95S0PutScL7AB3Zgydjd1aZEaNFi+mHYfY0cPvuuNd8Kxb
H9U+8e+TbfFgfcvkjkIqoJCxfCkBKzENyl0suK8uHxmah2ERs2icWVXiOG0Mgn8V
zH5UsAIAV5TB0rBMyG8Upyr1wE+puyHh5EmZ3XK/vD4fON5Sbk0Sa0fhCBMm3smZ
rCgpCR3sFFiBu3ywRH6MRy1bOuAnzJzVWQhQIYmdNqGBmKA9GHkHiqCbnr0+6dfU
4Eaw3gHfY2VklfgxEobrmiRn/orPH02Fh6oOy4B5IwVfWOFlygFSiSsuJ1ckefoj
HP0u7/JBUlGZ5azOTDB3CxH5qv8/zidkbwuFpi+PnhhtiSpGwn+CruwnfzZWNB3l
f+cR1r6e56Ud79U+/YYNoFiXdVwWl84UQMEVe/HCNP3iDtb/tBqG7oJxq1iXpWew
TL0fIHTyap4xQrtfTYVVDGvNIrDM0W3PMSW5Ibq0Zydh21mlmIbd9CAYNSt/rJ2O
KAkE03qT8Kt+Q+yjzflCJHg+DAwe8w++kunvZ1s5C2dQI/8hmY24OixqLr/T7VvW
+wwGtIkk+ml2IfDqUCTb/IvxqiU5eVHBiK/zVuTE6Cz76K4nCuGP61bxn4WS37mI
WoWXqQ/suQATQqIH+qzzQaYmGAFBSZ0911CFJdgjSMN1EweFLB2jxOzAGgmxW38B
LxB0Tg0x2RjLW2Tazb78FMKZ56LQCZSBzIT27CLvu3pRmNMud+6axKUZnRoaghAf
5LcsQUoXU0DXl6PfAc/CVrQUWrlxm5ZPZoGgml5etqHJDzw0priVoA6dTek5gkNV
3k9auHQ5Dv0FtOWXICOW7n2+DfSHAV+hFvicEFJN16P7/2L9pwjkm8r+GUfmFw27
4m9GMM1V1TIcOp/eS0Bkh15zwmYbMeiZG3TQMujGxIV9bTwba+MK7bqIpYG+L9Ov
5FYttaGmneOfmnTd5prYTdGKgo+k4KL4po3U6bwQHkjYoa1YWfJVaefamzgZfTs4
5s6Zc6xc4am5gITCN7rxmrqcOmoWZ4JzWSSsyuaiVTtoVEs/nKHr/EFQpwBsESOJ
oVsv2tW1mcrRcKzNGD7GpZVH3MWyUCEWm9cXa8ulQ7GfQiZqY9uQ2L0V0Ml0I6te
IUbV0UUQzliW+FreQr6N5ympVCAlvjCUXUPssU2xVG8x28RF9XeFHNVj7aTDvWCL
LI6zPJjJwflL5qDUqoyNoootS+y1tP4Sp+pI5r0ayB/wz3bbLpw0KagmeIA1I0p6
3siGXRKY7MQ7IUswwg/ZLnHcPuX7c69uThnxuDm6cBFXvDgPo6RIjN+xRPy6YCqN
YmVM34mBWnRe3l9MA55bzMal4fVvedLd1+AdmXSzU417+PWJfBJzsRACiEMOKsX0
CPg4r1d+WDtLQmdK7o9JQzA0UYMHV58gsrsJoHeetS+XRQMkbOvpozRtCA5XwSqL
1JIEpkAAa9cvWqgTQswcyVIHbTaiN8HSFkBCxLNIarA9X8KVsKsqSBZyhDqfD0JP
/Nv4aK57aEi4QvwnCGZvJw5dRCqU0d+oH0dYpecYCYgdvTFtZpWYifIyg8ygGBkl
+NY+mHTAxgDvmnP7kYJ4CoSbuT+H6HG0jMOctHCQq67IHy6ETjVXbfD7TdMn3yRj
PFm9FXJmJ9iNy2AT6wM485DLlX+y4FSf+72iLyLgtLHzuRTv1aTuWtqLUb2aj8Po
iMYL2DZCXPxizdXxyiBrp8nBS/JQqUg29M3HSZkRJDde3312d5sTtqux12BjPXHd
itzCPuJtBH2jszQ15XS2FWRHabDE21C6m3IHpPPLau57i8MrDabz+Lb6iwd2NxAN
fzT+ui2GfrySBuUBUPjSSd+FVJX+fm8uqbC1KrfJHCQHdCTwRutLQHNElHBHUeiX
QbxKR9AtQfNvUaoGuo4WMgojFo/fBjvZGthBqURxqH3Bj6Mex9YBwYqyuEnUEjyv
XijcnpSFavh8qrTp45BATATMSRWBsaq/mcWm23XX1IekCMJWiwaXuY0ZEXGrQAe9
e+azIbbuRUEHEisBL5PKtzHpegW7m8D8RHNR1hC1HNFI5ksV2JLCQOLb6uLxlwoo
8/5ju63YOO33tzu5lPWdqlptFVrHG8khl4O8Rz0bztsfPy7dmkpM73KQDFTjnM4Q
+Me/QtdlVrwAqD3U3rwVodbouh59u4fX0g/9saSWVSgh2I+ZN4eunZJoiVZauZHo
oqVyRSoTY7ElFiQJe+SjYRkFcE6tDZrOBb1UeK6J2bOV+XkPDYaAr4LRM8VF9fhT
5sUUp20sw+Pfs6HYAg5GzsEIQ9Qvg7xW83oKmiKfcdHqcPS3+nvy5J57D/76bRaN
eqrIwouxqmX1MGfOLEwDtH5MJIkYsM6WBUbMDTtZPcpEvvzAaeq9iB1GnSWED7/x
UY7St+Lzv/S1MTbozodEp/VbCnxjbiRkQ+TiIoBis/qCta9FCPiT75PdxZ0gQkuM
X3DsPyr/yVARFBaxHYf03XzTAIzuxuvLevX6dwfrIPvrDvzUx1ARU2JZnrusUp4w
5vm6QKe1OcOXE/xzw6mKuSpRptXh02sLpWDtn0RTQauc5iMbPfCPhY7As/bMkF4M
mTirsFAij9gDrCLj5zmatBPZfYZbNLVndMADugF/Jz8a6M3YVXPdmAeRl6Yf1bxf
Ofv0zUpFHgSNCObQSGr8eBEasa8VA9GcO0a6RZFC1q2M+gEbwuSJKMi6H/rUZS9z
HV6pJgKR4GCWq+aoEd+9G8yCFiA+Gf80JDnCl+CKNlTKUlnwDYdLqcG37gxmfxyD
E0lDTpcgWaJOuClLYcsjOxRvcHyxaMtT3wUr4aVUbDfXqDETK+lvsgzFTVO4OM8F
zymQP27f7JvBEtjkLXmH/+RsB3CLRdFJfjGutU8sNFz52Zp/KRcHrs/42XwIMwyj
y54za2potq+F2WUbwaeAoarXLGvbBgL1G+YHQkZZQIzd07fsBke/Qr74nAvCMgN8
h5btRjk+54Id/jBap3cStOKx3Q0lyoFVSMgvwtuNRPgnYUYoUzVigbSWjkI06w1G
I6po6YjYSNU+xFjZfckIzPp3yqYVUf4XZCovPBMCeH2Kl0qR1Jhlnuwr9WUsltZi
EzuoYtdAwRmkGjEcKIWpZdaxq+XdBralHrBZgTqgfQYi2A6Eh/TYV/GLzhNq7HJX
PvfWAvD7bOiV4yLd1eiTvWjc98H77lR4Rf9fCV6dJ8Ir3quYXx47dHrD3e7/+eRp
Ejp+/nsNsXwOvLQovXui+KMPnW6ggDxIfiqABoMzllNScx1P11eZlmbIv6L4+UeA
MVI2H1qeAlcdaeGNmpiwUXRNbdZkcWEhL4leC9+zLmFEN+YncxNVLddrh0b/A8/y
siFzFItzcWh4GWUHZsV98Sdm/5JIkaDKHPOizx8GOWURFAss9dAQQyrz2Hw3eOYn
jx8fheGafBwwUsVgNQiPut+ItW1x9KoS692216UOuzQ7Dl6QOJkhw5VdLTSwAjQk
+7KR9R74dKr8twUabt/MP6jovtxEqndCA+7DbCnIo8YtH6g5EfP4wsFPCS2hUowD
uwRzqxnfG/0u7UZmWJl0/MChpcqgLY89mUgBu9CdAkiC1MIadDbVvXKkq7ntre7r
Bwz5zvgpvs9xP9taHotUsZK08XoUQ/V8HpwdRgghKwQ0Vx7PdWhqwR2aLflAU6Lq
s2aC06dDqMYo/IfsSnmPSt1aaeBUtSvBe50vbA+ab9wpOFLd9YTJlTzY8k+EPFZY
sydtoqoSnKA8Nvev/qHSti14n4HF2/fgiZikXW2u3m6IHfUESlVd0uyaJHtLbliZ
sV1KzcnfMk6cabFvi60vVmhRnwizZH65cdZ4S0iqktF4OiEYuQ7dn4ewsMeOsi7L
xEpOPFpT0YsnHeJdQA9JgzESfXd8WRvyU+3joXGG9sdl65leEoGd5O+4LU6bSmtU
06YidsyDbZUelc3quOWB8zX3xZeK2e4+z9x1HssQy9mwppAmDJUmLauhKti9Igi3
z/hGgatYhII7pweKL+Qs/IIPrymF7+7zZQ0NObCDdkQgkPT3cGDdA6K2PlZuoKaY
r1MW2wW92fM71FgaQVuXtvV1qqrxqrli0Tp22CT/yJX1QHcR9/QBVrDClZ7EqecT
qYq0bpjxdWNf2JEs214ZWRLj46xum9N+1VxsEK0CaPVkf0HwlMw4n9bY1G0niuD4
0jZ2jtEHr+Ce9B456v/0i4qskImPoBx1ycEYQWd0BgvkrncnXeIwiNGqeHvse+bq
t9+buC3NRGNu9TCYUmGwJv4jm1+hYTWMgbMgB7Jakn29vcUXaEHu8OLLw5uCjUEN
MQrkL+fwtfnjwTpf3Sk9Pu9SE4Q+tNYyvfS/CuONkJExmfQv4/5+gPDiPNQIpEzy
FrmlI7Qbm6qvSho6z8NZEk/TytAPTlPP/lHBnh+BOgssu7y3Kbf5UKY/kMQBNEOr
P9DVt5EULiw+wisxL4Qin88CXdL43dki1bSr4QGQLZAaNZBS/vtykrdpyO+f6hik
6ZR5L8pJoJjbAF8sDY4ipA7VEIk+PPpl++bQWShgSkf5YbVOZoaOOT957pncaZzk
98Yd8gk15DBmUvAEyBBAED8LAKg90tS6a+kJUZa2YLCDc4mRKthnwkCQOSxIh6F6
hABLpDzAd4EpXmpPrLbdkNMHjv7JhU8yz5LJCJh4RD6/Dn+7ylOf9YdeMzCC6yQ4
32/JnQQwLLh864W5yBKFo++HfA1ZK5ItyMR/Ih6+94mmjKh1F2vWJv98L++efc11
2m6sgaMZ43Z7EwsI019CMRu8zRcr3rn2gqLYIDAD1io1ynRWc9/eQFIwwv/mLiHk
N1ry4xIgU2ek/fO+YqhENs+3hbGr2BEn0KLLotS4t1f9df9RRvS90QugtoYz9Qju
1+4nQ9TlN1UBsBKi/TUjialWaKqVYF1eXa9m3jgllJ7b393xeUfYp7K2CgKt5NLr
6Y1456Lyd6TX+r4pbIfCxHswl8hCjIdTjWU/O5W4u863BEuYDcCQnxlFKH/FN77A
XfJoYtPkzB9UPbfce0r7l7Pp1Hdz4kudmzDla/EW1EKbvFG2fgBKlrIrcQI6wIWS
Xm4rZKwFp5fZKZEaFlPp2LybmUJBCe+wP/pY+WnweTsVroabk6sOaAc9aV0HKG62
KIOuS4kzS3o97WQ2V71oG81X53glA8ZFwlUMd/9LbOKQS1ZrldDZ3QppSTSlYkWx
+CvnD5ce+gMlZU58wafnKSN63xEpuzf5r9pkwj7JO4/e96bOtd/7UAsLsJiya1hp
I09aV400gMD6Oe8nqm+4Bzi76s8l9lSS68PzYSKCPlb9oRz2ex4A6GtOiGrzET9/
NegbDY3NpugNX64+eK4zAYrscmrRcyS7dvCx3mb/aASSYNqlg/NuJUk9phzhonT5
7rlNZR30hZfl3Bgm32vlJOSU9zGpDIkbKX0IAnZEdk+ZIIiK97iaxUkkxbeUALeo
qNxU00xeWTDEUQnjp7M955xv7chIY8+BSuRbgY7QFvvQXG2MoQqL9hb5FIP809gk
tE5nAw8w2fd82j8oxZEJG5nTFmNd03GtcWOCLQQIaE7QfnAv9gvpG/WxjrDh9IbF
oiAA7ZZPnHH99aIvO7sxKYlaLogSuiCMxUcpKS9cvApi8PR7cL9u7Szlvdqk+O2v
CD4j0sdHOikP0Fbqn4a3MMGofHkPTKP/0qAIpRkSSWHbVlnwSGq/8Y+6WS8FnnZs
Lh+CalN45uyqsHH0p0XfhR2Q+8OyxFlORRqJCF7FTZnlL5GSLpv6jld7IjNgGwNM
CZVwDymEmRX7tD3XH7c0jqf5/h6Fg8XzG//Oh6dSIszd3hT3mIDM1Sr9dTjOSOzR
FLEa+c2fGwzuZS/roFm3KjCDKUvYJWy1P7VPhctH6F7MXMX8mYCD9Zk5rdMNb7eB
CHvtxGDvZgpiLikQLhYYS0tg8MGO99jXmxz5XN3is9+siVD5OSoxqhOGsAi4kZqW
ckvhVHR7SM0DoT78Y4khgPX4saXrtXRkU7E2DviRmNZrBfGdWdZIA0Q/wrRsFgJb
Wq3k9AfEHL/47x+8OGMLDrTF6mgtoGPjty6OcJw8ohLy06p8Cmz1a2WKIhJkDVA0
+JBdFrZwZwiYpKQC3LgiJhgsSWFMp4bH+PMsNZC8kEiz1+SFnlbW8zwVSd32aj+i
V149/7rSFwp5otHPbcDx+/COb2rgn9nPfDaBkofn9cpCqH25hik0t10lFbIkJHmx
YZ7CBKXXeZmiNERWcvjB3DM+HfxG4L45XeRdNQ5FHGzd0apthVzawaF20XE3LdCY
y3aIoEFisyqcvujass8qPvUycHXYAefz9emvd+K/8Capzz+LqVvZP/zLryjiNNy5
VrGaeIXbUFS05oHPoo53YdJsgxaF4r++dV6BlIM3RdEjgVvEtAmFCbdEsIw2dvjT
rmba295whRZTYzZj8eVRi1pif7Dm7xNUvJ/SaCf5lV3oiyH+j1lpyJSuK3TGjkds
6FD0ZmtjG2O9Uy5WbbRH8zU8SZ4Y1umOHc8ZJxpNNGGvw0vDBnvv50+5VrOpgJxD
S2svYIuhyatXeWFYBgrb7QhjUENoXtaBcOgb9sVPG6iwJ39YkN5kuTwtVx69jsWm
VLFJ/Nq8iZpc3yDE6hVYhN3AOuwFAQqs5Ct1b/d5t+MtHtYbCbsHXBwWpk1pBdMR
3s4YM2tq3kaGOSnL9LLK90dN/FVVMUKBImtm1/BF9AmdAzogZ076jyDEgHzxHYI7
uLo4w1D2r+KDbyd4sHSkP/63p79fT2oxE/8g3gjP6yq2WXgIvWYVZLcjNpMTbKLW
sjCquJuCTNsJ++YkxEv0lvqEYjVOOy3sZIwU4o4piCgcX9x1hehCm3Jnd4esWsAF
TKoJVfk7XPQmFvkISJGgiAdNmlqIyTXDReuS8ggWznHT5qOvhy8bSxKMtdJhlqx+
3TejQUojVcdVZC2l/Y4zxam6w1iaWOuw6+16TyF5OPM9ILoIdTUAbjabovAixpTs
5SQ62/P1hBTiZInrhK/w5TgbPpqfULC2BR1xS/9Xp3OUgScJ0gv7YpRTHEVwEMSp
+KCKjwkb++79IOGez/JyFUnvZvxV6iot3SYweLRUkimRqTJQnM0b4WK5OtFuCa4B
YcMJhJoIufu17k+3HmmGYDyyWaUEvSnMJ4MZTWVEB43KCAE/vd93sGyu8edx0IIl
7f3RFcf0Q+DS7GtFbKOkJ05/iHkl6XlDvDvhRaUH0RlC6yj5Lg2+0E+rbCPJqCLU
nSLz5hrap3O1PKl/UKDQwlGKsYZfe2XueSrGqFYkb9/tjnBfkjPw8kpA/xuOB2sd
VoN5QOaMYjwqHgheLiVfdBhEymZGQSx8YzznhMOM9qcwH1c+IytbD//zmjtlRn3C
zuSPt1nu6UdEPS4i6dA0fEzwAc9CW+WEygnYtXF7TFJAj1l3vGKCkoxyDVZjuE2m
G7mAZU7gGCSeLT6iUjXUBErgylqoRokD8ZLuLGoqkCzcfUMpnm5b/zJ9MGDy/xws
PCCJO6QtUT9UdY3UFv+sM2CmWt6p/bu2Z5/oOxcDw4hgt+wn4BrhbZnLsrRxPNgV
Kf9b050hHrz2CXMc81vHMRxnLnrF6aPJyg1sRpkjuDqoCnGbTdzMfjpfvu5hMwuO
1TJgaaxvUhrHzLwgebVvj5IaK6pqVwFmMm5+obUGLQr+p+wZorOnAFgR1R9iuTCH
IvGIGB5+Acsrd3ypbjdNbEYUhYbBCY7mAjlJlj+5STnwxaq6dYMWT2tga9nrrNjo
/UMDKhpMzkhXbom/E3+YKBMlyX8bKqKy5oeHa6TrBtrYf7OIJfirbbArcJT3rPai
IHVtiKGIwzazRtlUmN12XLvh7aioW3mKnHFm7sU9CeBzByuP1vkeb7M/uyM8iclz
zreRTU5VepWCzGFLzLZ9cgF46CtIZFvvEot/L+crD1/xq59H3DRjxfE9aCawdoCb
kI49VWou7cMVLXLhxLhZ8BPdYFsCkYFsQ8070dylNvzhxgHdiEg8EwGdEnt+mV52
5nhixS1dPUA4Yln0vR2Up56X6nMkPWAc3vBjye1xaMewBiRgCCCxhr5xoq6gHlFG
3Sb+VZKHQQfyblOMDt0TeBxeLlbflZ1qZ8KCQGA86+tAQZopToSQJyZ7iJ3TC9q9
CCYDhdXDiwf8v06OtKkeQH4bK4PZi6i2j0ZyAemp1U162lwj/1jb/BckJR1etthX
HWLis/g+IFkBJ41UREKYM+5pqtCFipNbbPrdPruND5TXJWkBdH0P4ET61MvTK2dI
KjTTQ4XK1o81W+/XlRr0uPHbJuaDhd7ldAzakkV3FKx0XlzZeN4HklHhAFK0nyLR
rg4hbEOSd8O6GOMSXUsKTFR7Q2D0TgNtzIzB0v6vjw2sy5qwkHy+gObW7Kx8Wbj6
cPra+vwp8jkx5eyuItv1XZ5vOXFJDGIE6pWib2aN0XHAv08wG7zvy1X+0BAT2HBh
yFi6pG3hXUIIMHGLfczI4Bh7lMz6AYyPDmIHsut2nl2oB1UyTBGslgGS2jeorXKr
y2f+xjiE8lPQWjqECT+BndDnJ3ifOIiEB/FRXVQKRA7dC9zvn79KZ6pv+dbyefs/
d4HSx5m3H+eBPyrgUvdqlX9NZ7TUn44kOeiNewY0aTEiYRSSHW3Ogoy6X2EMflXh
Dhnp6U2f/tvjPRnVI9XrGaMyBY5bSWSYb0x1Oe+tuZO8iL01zwsAyKjb+hKUL6yj
segVOwCpasr2Z6qitPZjHSMXYpk9JpI6GyG41R5/4kwj+4y/NuHapHhz5zThZWSz
3ct5gKLZ3SovdLm0qT71ZxZalmThxSO7I5Ik48riMHldBuoUL6ATJhQIUXg5ZFhF
ClNCFz1BpXcyYpwAPlYssm0flaHq+nwP+m2+F/QIJXdyrgnMrY+uQB9y3VZPAStq
OPnT6pX+zBVrCZpyaL0Gbv+8nsbt6N9RTOBh1BPPNKf9ubAlup1F5wJ/uh9AmwLY
yZ3PRIwCkc19wM1PCLUqsMM8jXYNWY2baKWQNNGGQ5SJpJCKFRSS4qYEAmNYqx1I
H+aN/P8ZrLANqkQRbai/zOq4ohgBMAlyhjFK6AYSLD3nyFsZum4XSi9biEd6ANap
g2RpkW8tpmTG9LehteZjf4+/v3dXYYv/j5KN/J+Of0btf0qpgcZtO/5ucieM4Wtl
5iPJPyWkT/J6QGZfWlGxuH+o6aJbvwPjSYajx9DeCPpcYffQtBo+JUpMqJBsqHZK
59UwtrjzV3NqbXjs5sMWFyaEeOVKVwicJhVd2WtlWruGeEzcZ6DADQmul5RrJ2qL
CPVqhXVy1Fth7/D3gN0+T0V2JXXymNAV2eU+I6MmI568hFKcOCAO91Vijneqwon+
Ix0A54yGO6sKBzQHkNzOw/9d5PZP4jq8cxqgGUMY/RP6k6BL/tt7fTFAGNHKQxm9
REVkmmNmyVaPrKnKJNBWkISNXPBlqcysFkvCdYsZBZZkMl/5wNvfPmt+Oxg2DPlS
KF20pt6XGru8SZZJMWQOYAxza8CA/5zJ7RNBpO321Op8/tGsmXH4K9iAMG339HMT
eUhzlKzypmq7Ka5BzNUchheZe8GA3Q133X/qA3BMyz9Vy8u4gzuNjB9sks+Ae7Km
0yAR/Keq2vI/imFWYPW+dwMd8piCOVKLOsdJRUWSwdSzPBpCjBtrhPd9NWP6qykm
W60Y9wmN31HSS4SzNLCP5vXOKJ6CuUAIsOSWYBiqu8/qFQ7tYRbytysd3acPnKBF
W7zxG2E3C0xswJZ6g6MuINvE2T3pXMcrekbpe+GEEtcOSzryJazifNYzq3UR/CmL
rEkjOAF8ivf1RKNRArTsgfZJ0Momw13XdJpejflNXI3JmTXy+Y61aGCgzKjBR1og
tVZt+EepG7XQnVL1RpxTQKIm3xAEVzi3k1fCiG0L/q6294JqFJ8vzpAb0/daBzvH
207Pc0DyFh7gnviSREK4rfN5f+aP0tAAqTxOG4h8yl6iGB8OzX2MshGtZUd2fGVv
JBdm9leKNmHbpSLkjRdZvFuvFLzrBBH0VONjwauBq8iQ3arjDPpnAPcZFU4lIvY3
NM1M8nRITCDq2o5Zr5gtrdht2+B7xY/9C318Z3FpvKdlhqOuSvBAKAdY2FaYYLGQ
ClvixNq44PMIuXiXreIWPq2IFM1SovbiWbDgB+WZ6LmPl0fhDmQ5yPqFm2syU0pI
nETd8MPdQStIZkF/IDFJlf6Semg2V6lMY2MTUIoLgu7D+ZZCCgDf86RCEo//WSqh
DA6PmYaU3t9CBDZa8DTyyo/G5Yt/7YgXV/uOHAgkN4S4vwH+mtS20oWcbzujShR5
Dk5TCL2O//JPEFIzNaJezel3gYquE0pl2eMrLyAp/JW5orrklJVtb/FpNreqTlBa
QJCWu0diuExk2V0p+yCf5wgNxFsyI3ffbU2yWSj5tBZp04qP/eSUpkmSNmD7EWto
SEWfWZCGJHdX9iUQrNn7fw9zog6jEis4zsAsiz/rLNzuI0ayVCANm3Zg4qvFvDP4
IEOyW0cWS6IbiNfdO4te2NTLTjySEqjW0b7V2HP/v9fKmzKLrkf20RjtLj1AS8CD
M8Hxs1ZOUSmzyXYV+vxQYIA4eAs/UZMxApA3r8771mq8v/4J6kR/60f3wXQti6Fc
amRgmAHP9f8q8Y+HqbRacupbuFWjMlcRl1E3WqLn1wnsZjaBB1kIE16JqTGubOHT
22iL1TDviocPFrUrUzjE/9u9SxyjCYCD2+UDuQOYsrkWpIRrUk/pf9ZbGkzY+Phi
ZNqa/BYlJDODlrfk/gQsHzrZjH2wuDs8LNJEFD1Papc2YtGUV8EjjWQkOzxn1LLS
6EMNX7G+1HHwNTb+nxZr4b8EEQWoFDrxXDYJvsYZ1MtFh6ujvY8e/8zsUkpxGVWm
yjsHMruecv+0Gz3jn7en8RC0N5MEBnSIE7nxeBc/9xG8ZYRz9w7VKfbqGPFA5Eqa
HS7I2DYjHnK90WflLkZK/dIp6h7DkavWp5KjkM2lHwtqnAao2BvevaPzQ9ahywSI
3eX5uwvdj4PJ0Ez7V7VGWZBVK+baS8wgKB4jxiZULwE8/O1phGhQAa3BDFD0iNAr
080zVXdAtK1JcPnoA6nwthJWrCmonC0SU1hhowlaNcZoKaucko1Qq0qZxQR0QvAA
1/tcRGadkufoqnGT1U5HisH8wYlCE2rz0zBjNiXG5HRXDQQ8tZGkDY3IuGsJFWuA
yeoR1Y7ajO8XhnmZ2lPqRGXcWJx4FGXyViUxM1UTLM3E/A7Q0pgnXLA9QGdG1kXS
5hbwz6HZ/2t5DBFszMzaqEo6LBvx8F3m6uGNFR3rXv+KQ01o2/Rxt6qDm8IZ1lJz
Ni30Q1Qtg1Jp27Al8LuFJmg8+vIogtwLlGy0mPmY7tbe6uzpKFZqILmWjspqAy9w
ILlgMdkG/YmHvSukaLXnqTAkTZRF7UC9gKBcU/Ay0BznUjr1DfO07wlqOvSFbl4+
5dyiifCGBqcfrPM+MxhbRUiTjxvtAT9IRDSgubAeQyBavbEaBHO3h9qCnAnhgmmc
8g+rQf8axHUuquT86HKiU91KZgr+OQcSR4oanmm9FVZcmo+Aa+Y4xXtMHoHRTzSA
UlbA094Eve/Lr7IFY5Ngh1IWNPWLn/LdaaYNnm7DQ10DDCYB9lsMO/2L4zzNLbiO
jtcamjVPurhzVO2/xtey2/66d5SEX0n0xiWtY0onb3FZ+s0W2LZda+z8bAmETveG
l1EGMjAbmr/ITIVCj44SA2e2KvnspY4CNIU1g9mV8BDDVV0awOHV9x7JD2MleqBP
Cd3XG7Xakb41neivdYt53M60KC9VmHIaQ6Zp1gIkusvyGgNFX7DzwbDBrPn+lSTv
JK9JikSR0psFfWho1XN0eQoQu8ERpmCmE5Xe/ipxFX7c4qLC+hlDedHj6q8dOBVY
aVGrxY9gXLWY12tycdPOpNcvgAiCbtIwyG8yCHt7PV2nFK6YPGsyqWVM4XGzQIwt
HVvp8dj4JXWOyf90JRj51eO8Dc8PDWDUqf5MRmSX49H+1HGIaF+TvCzaRXyl+sBk
2605twYYlfQNtTKqQOLg9c2Mq0Vtr9gFnsN1YrLGPuhNiLpP2CtM+PwIa96aoGyk
mpEI+oLPVa79XIxaTpsoG5ZGkR8PSUnzrYbGt8ssWsfmWrYvr5RcNKKJF+h72mEL
7/9qyB/mPtr8wTPwpWxIPeOW1u8OBh9wZNAe2TcBkvRKUfY/9NFDmZtrk0BMmf9h
JwQ6rvSs8F+TX/eusXftaWkRt5RGCe3eM4xnOUB3wcjQ6TgTv16eA7Sl9693RepA
maBUqCqLQE8TlenbpBk7ZqnW3FvTKCm9dZ7dn9z8oiobzatXqDya5E+ly/uas5D8
QdpRgyXgz2P530uT0u+SAjqAv87c+0K/F3o4D930C0TwaEvBv3b3fQBfb3+TkcKJ
OND62olj5hYycVXlqghvVsK77PiyA4iovscV6vJsjPbd7H7EmLr1K4atHofwYXYN
AgAvM9lndaIJoNOq3BZmIbani1reKgYa3GFFqFPQjj/gfQhTt7OOrA6p1lQxkqhI
2OqPrW9ZAb6T7MRUgQb2tM5Z1WykuAbDctCwVdgT4L+5+OxZnnopB4Qznftc4Myr
Rfb56kaGLP4r78oKOvjakNduTmEhU8MPtGB2Qev5PRkVz17ujVfSmlSxa8C5mxdw
O7jvswkvoDhAvveThW5J4t7y9kwPL7eNK/QiGsFX4DvEqn3TfgQLsb0POk1mxCxo
XXHsu3WtNJNvUxFrGsElLFr0o0+RzjBbkVGpKanDxhnUxgwDxTILx/uv6D+b5EWc
F6eMONjyl/61UIvzarY+jq1QXawcaBSyWniIUmycA/osXRow3Uux9s7XUP9uytR/
L/t1Arc9TsiTySaqlPG8Ms54vH69hSM304ZYCDZ1P4Meqdx/gTJuWKiFhbnTeymM
R9XEtFADlG5ZiFKU40CgJQ3XalEZML6XwfF25N5G800W6zAuWmZrLqu6yIgkdIJS
OnxievJwK9V/iQpLGiTB+B7KOBCR1ROr6ZolvilB7V5nk22mNYGL+i3As2AFJ1ZK
Gg+PwZ5p3ZKQKzAlAOhjV/JkhFm4TyDuK+5xdqHm5JJEammVpBvzUiQaUsE5mInr
dmQq0EXju0axkKZWNK8a33PoHDjL4Vk+y1amjdEnmDJ2vhiaEBSh4W8c0r4yEhIL
pil9svY2B/gei1gHJHveNRuvmJighK0B5IwrWj5zU91ZxBdaonHn13FShigcgtFt
qviW6n44wA2qCU1Bl2J56rDU/KnJhbEZc07txk3VvU2R9K8S2yjOSW8ag19eCqqX
bJ8jtXA/GuUunDviPHNL/sRKMS2mcW3aPefevEpC5AEfrJpxVo+wHpMjrxzxC3Uf
c0Jwc/ZPQdemv0/9vz7Imroy5PTHG7+AYP9IGEsnV5GVAbuecLq7b4BEIHfHvAtt
BCh/V/sDXBqKxRzYv1+0Q60gs3DlwPjuoV7zbXqgm480M71z4nuxV1x29zlLpPSW
TnsxTSEByqLbS10dTB5H5mYKTX+euz0FUpiCNzYTFBrAIsFJIYe2zHQ1/9rkT0o/
hvEnuebBc5UU9h472NdYJHf/NnpTWk72zzjYdgfnHU1O5qFoSIiDwTShibD6ogni
jTT4CNRyr+/Vb18iOG5vbjTvYeSxIKVUEjLnLAjF9WfWlXp+Mc0Ox89eiJXtlaZk
UAafTIJst2UR+XM13DJ457e3+sDJngjj4LOK+4Ukv7vScko2KaUtyn1g6QqivVXJ
I/Rk1//T6YGSxUiQA/AuivdDR8Z5R3oNywMryQBAs8xUrAgKvFDpeq9bAUZS7HwE
v76n+aCDxCdE6Eh2s239ZaB/T/IeNN2vvzjAcJpPZeagwKhs6NzKqRlhIvJCiSRn
2khOVMfF/i2kIqlfRTdcwZqBnLG3CJR3EUGMFSuuU3OA5O28isPBphTwpH9aaoPE
GlmF0+z+OzWpQhW3ruViG8wEZj22dHmUYCWeOuA1Qh1XK1XH8PZsiSA6aX9EL94T
phPNwLUmzZ9Ge3Yw9STzqREXrbliaHThAZyVriv5DaS64BNZLhsZZJLlMEuKOSzk
Xj7na2Ns/uv1w6xJvS0AEpNPfXP0x+KjpNL2QxvCIk9RCcOiZPJM9llAqFxnnpnO
F8SLvGj9DNoOdhFBPwcHz0cV3DD143fYluJDDKANXG4eCwl5XcVRA6M4LNGRacsr
X8vZJN7yX2yzmr+w4e3iHUgjHH9GV3Ij5lkvZZouLEdg+9fz00XMumYFy7yEzn3J
iPdbpP8V+vSSX6Dp+Sukxg9wduM3/tW7RUEyTCeTb3hOIIVs8JJAXR+vKNgzDBbm
RZGeLas2B3nv7LTGsIjriHQ32GS/H8ZGMHVvU/Dk2hGxZtwBaP2lg3zLdEx3ZNqp
h7yU14DitUmV4vqHxjaDFGZz3tgUWFUvCd4jMMVWrvytdf/2qUCdVnNQEOlhIcwf
sW3vqbh5HF4J2cLgsqXXRoDrMOVV+GxObFEDuOV0imZLpLh9d1sMdQ2yNM8ZFpGh
EWp+dQ4pjBpAHnsCKgjWL19gVMZ/QV6EVenzQl04gMeyBC/j5sIYkAVaFtC3qG7g
Hw+cbAM8OqIQhhOPpTrOa5L0vNdYWOfYdatVAH71KvOLuSfECNmovYVqWiP51Rdu
rwkWVIKITquSB6wOOgCdJa+D4K5zImYZ1ECqrQWLPFhKpey0z6cSsX6gvPvt5YS+
7ALwomfODkiHpUleQ0hMWGCARJx/PcEObqRAWH56rHr5ZQQjXqCr0sHrXyE2yy2Z
yA+h4mr0f89IBx/YggiqQg58hdis2H2D3PS8L8v664EyQLOjwTYOmwLoVmhiBQVk
mTpla4mUzchbAxmFLcs5cdS4ggx7ICbcEOu0LowrLvsiE8E1HlRGG2SA81rv6XU4
rV4tTuolG0O7nJOeKQCO8sBanndViJzCrfV3XDmNGE3YSxYmgetKH0DWw+Swc3kz
Rpq4V/y/M7XdW3ymh+ksGXrpbKzgvOzfj2kKKacTRM9uWdRMOHTrMGkd32AGaXHP
iOiCWZOT8hc0BfeuaCdei8jYgxG6fHxtByGC8Q/NSoux+cqblJhichKq7xXOjf6b
P1gTKvrTtsWl3AoFznmRkue8CPCyNhZesD/ke7V0PlGupWVJqj1Na8CCvQDaAq1+
LAyhoYMfNc7pKGCxTamLdf9sJnBRWtsh2Sy5+OdEioB9Joj5E3LyuI8Pxooa6VQw
oLz9FqBNfButKMO+IVh0EjHwsZvfW9aZCO2W7Ld4GeUh8F23XKc+tguPwbh94cwk
2CDmsgB/Y1550iORShTINree1GgIHu3kqEtQiH3Z0w12EmJyuVW/75bUZ/xw0bB+
msy51+ffOpwezGOhG4hmwwMWmETDyylO137iC5c85dg74y1vaCc1iG6N05KDaM4n
/hvV5skynXCDG3XELzx78CAjo+ZW8Btz0NYeY/Z60N/dXpQPlQ1oZ2cKGj8iLRyU
x9gWKwr+SyTMfVJSmX0/U+B9TCTDfEFDbtkzAt+yHy4/f50eolOOSBKiylT+ituc
i6HL7a+3lKKRVvqgjD2C7NjpNETw/e6ucRDpqZh1jZfIDNl/VYo3Es/0KNS3x2l6
epPMuRu/unPAG5iSARPOLxb0hVvy3WrFnSbsE+6NWA1vrpt2IBj/jEaJwXhd8f0S
BVkkYkHnmtybFQJX5FfHd4rgYfuTVl/BoEQIKLstIBoODexfzeqyv+pEXOD7Et9g
q3dAwLUblq04LoagokrCs+l/1At7VLCfAgsAgURR9MUqpmYvHwt3EbToYeqmPMNj
8vkbtZUtc3FIXK9vsBAzs80eFRanYbRwtFN30KW5mJdPPVMH5vtYFiv8gRTMjaCu
DKaNYrL652LfN7WQaJ5EgYYdmMpZKsp9kiILRhkIhsQShFBRoVuRqmIGeMP+Z0kO
+wbzQ+xCUCULj4Z0xjvG0SVd/to2dUI0EGlS3Mk6YqkhxZom0cQfy2mTUpI8nklk
LplyXRpe/KgD4sxZB3+uy2BPdBEdi8SixFmSIcO6uLUcBcdZoyWB2n1dXLSkc2rc
bcJOHJAFiGoHQJFYJ0sLml8hRmJfw0fUCUOqKnNTo2yRsumPeqf7FXSaQlXLqfYO
0Gv0fVAKSSkQkKlLzjmNEd4WjQiROgrB92oMBLqadfgGmXFl4Xrzln9v7/h6qlMy
pmZMl342r9XbAsa+HT0OChmIaLdlGbFQO25Nr2g++uZ8egBo95VhCAIqjClgHGgm
xlZytxwWQc1LpkYRHJAiNZ28fTOqKbR981+K2FMqzmwKzGIfp4KvK4QPqqL/Hnra
xaW5fxVzlrsYxDUGJRo/qi1faPq5s+rR0T+g9AVd/CUnnvg0pxd52JgRj3Udws6X
IjI2+7oFTWIvkPPMB8otYFcNSudwjShVFaMBYYdUwuIdEgHNOdysfhqNDrmkuID/
9ddY/sxo8tNPAaiJDL5QuAnoYHAY109RA78014is7H4PUzqu9cJyGjvKgEi3fZye
tqlobychrKETsvTTUr/13aSnZbM4HnQ+5fKCUX3so0swglX/8tN/B3ohCqQ4+5gs
Hlqtl3qQOQRK6jmSUgxWFei6cQfXHp9VjRtkwycFe8Jw2KnBFo5Pcllx9wclhc+b
OQxqIOpswroGaMCOFtBPi4ciDusPGQ29oDl3G3bLjL2Mzo1x+dbKVsbFP1LLFsjF
9usm3UZ3lteKemKq3y6jKqRYH6ZQUj9WSkQcHzJaF/KMapJNexPmNH2CaJH+tj7l
ABsF+WxVSZvT0jRJgCRDTtrzJFl2HoBJg4G17k1qafcXzJBDpZkw9dLXYJW5iT2u
2PZCBLa2cBqjCPGAM3Up4U/vqBnVp6tlYnmIkgN7hVAQI9SZjnLKGgWk5EhTzUjv
eaSU3sOHHFUpHm828TjbvNBWguq0JMXYWp0j/VEN/MZRbMkodJfemmPpzAQffJq+
ggTFUGxJNz8cOWX3y4WS5+0XVn0mnUqlvUKkHu8yp/8nQaDsWWzvtXQSnYFMKZSa
gQamN5cpcMmDNKTZjKp88923sjXDhyNYBUuE8s8uc8aHeuOhXLksvDXokGz3lpgw
DjmDCdYz745LUrVS6CPJhCHrtYZGRHzCqf3Uldbsxym/aVTIi8Q++DozfLfRTnn8
0mBDQwkRZOuj8rjDPWT0AVobZ15mh8vCtQx4L5WisyU+tUHabNXa7pOroovnGEAW
WLXbKH+H4Y6P5mej1VMGzz9tGHtEozNwy9xFWCWxZ2IMNio2VK2MDNBeayaSIN5y
DdHauRjGHd8KRl2WxFRW4kij8F8rx/nY4hzSM1pVqqn0Vgkdaaorp2byoEQdqplh
zLGASE4Yw+RyWazyyNDq+/zsK2UHOCnqBn+n9YIcBE6hyFgGk5iehknUFC33Hz7x
doforFLaR9w1cEMfUrkhXnc3vq24A4IlvjOwHJAqf3UDuTlD+zq9JmnSUR6LtqUY
rXV4mwPkjHh9MXTswiMPNBfNvgHZZtHkeZqu6No8e2nxeqmhJMY2J094LOc5Z0ts
w1LYG5M0cBBOWRakmS6XrAJbSSgoeNxbzZbXgHygYQyO/TWoV9isfZB744emDVLF
tKj49EyKMdxi55Oq6TwYENVCPPLqkv4h/ugoFoEoVr20lBHhyfq/FRwLMfiFbwQc
VkpyRpeXDKmIFSqNq0rBw2irvP5DW2AAONM2t2uhkpqaaq3/9HNrDE72ijyZ2LPs
q3wHSpTN1YC+dim8PREoDThXSUrhrs+EgSMKENObc/GRBZT3KYJIplix8ICnFJGg
o37DPIea5Pc1wmEyHg4trJpwMKB0OzIC1T+y2t/uOyesDTvpUrV+4Yfkx2aL8P5M
DygVAvF9SwpuoiYLuXfZsN5Hln3CAOZyEsMbqi6PS78jrsQS9cQrrRouduMqUX0B
STJP47vnGTw7azQQduQmjpbUgGgCVBnPufKtUm/HtgbnfTzWr2ZbvQz4vtGLQy3n
tRhpVIIiNlVit3CEJ2LufjIo/ND9M7sMEOcpGNZw3md3IkbdaTWnCLRBtl1QIIA7
XI+5j4L+F2RMlMOyKzuM00kFLMt5i7c722VKI6GctvR12n4MgkPnOjZZCEmyw8Ah
aa9NbnNGo2yJY/t7URDJKRbvxqWZhPT3sFoUcn0zRytXD1cN4aeQJjLX2O1lGfn9
wbfgEFrPg+vXCvoury0xdxxyhmDB2zdmDoosCm7RxDrTSHf0Lybgc84duQ54euDe
aCRh0HJ9YwKNuq2v7Ziae/+9WvWTMot/pvenhVVjPxylJj/87m4lxhCp0+b5T0fI
e1zyahts1bMK7VKAQvAy64qq7pc5Z562LLjN/mvN2RqZDeyfI+33xNjI14mSmvwq
XQOk7CkIyNbIal4InuPD30aDMJWuBJxKhGskHO84aG2yWP422s8w3fPPEQTMBmQZ
tHFvNHA6xYrrferPRVTscBpz5mb/DFIfRL1uzHiNmYACiRCzgmg1HXV0H9T099S+
NGTy43L9Q+EtkJVEOeecAXG7pTmUIqUqwpnZU6AfbO2iQriJnUy24oOewKhNv1pz
34opALFBNtIINqSL+MbOSPIUpuMuwIbYmKitcbGnzalg+h9Vr0OzSfrhZa0cfY8h
HhwDh3zapDZB3vPR14YibxIoKTotrlpdsMOkV5csiaZGIvtOAi3bPHMmRw0rYnJT
jIcOJwd2YEbwMbowugFIQ6kRsRJQ+Xy8SCl8cU3i3MQ0BbweqAcZiCVrcYqlrN+L
iLggsfPmkbKvwJE0pfViU+LvlznFdB7SofJbBGVoLMRRuOYbl5hIOLEcEKm3wz1g
kWbQ2Elpm4b52O/VMmm89+0AMqVyd3Xf5V9JrMHm9NPf2NDTEaIlNOBDq9n5RNg/
7tTPmVFs+TOeoKjAwefStQL5l7q9ZjksHMPuv38fdyeyuVhG1WGfBbT9fMMoSpMt
umLbQr6E61e1sQUTVM4AyWO/vbB9sFCkaNmXydG9LLxnucow5TSIeO72Q2puHRdy
kopqhpKEltZFLcUcZZ8R/Z1ta/tfbeyOyJ9/M+BpnMwFaFyOtNFuJgKB5dugV2Kl
+aQdfmkvF6QsOoHz1CvIwr4hTDGq3ZSJHoNWRLBUxTb0ZAp3MsNPMZ3u4inq5Vfi
bcbI2JTvXB4Zd+YbeXHXpfQjltnlruYfC8LBZ3gQ0XK6g1WY4iady7GdmhWqrRPl
u6fldPgsPkAzSQVq/n8lSaOF/oe4E7ODTFQQJyESKyPC4inPJmH5x/D5ySEEmlQJ
tgNSkrCi0GcWrD27NudSQ59VvvcUNw6cmBJ5YLwJp7vOqoVk6RXw0ceAvGUNQG4V
nnVlGzg91mmqJDlXnLEdqDaN5rv8B+5bMr4yFe3POxCymlcc4xj+NWUBr3USj/cy
P6dN4lr3Spp7HV7nifQx+pmy99HkuOtc3RPwwGO/dpmOYRTZCeTSM19dh5orZGug
y4xqRAbQvHF2/Lki563/Qxa+8/XhqEixVrqUYWgVrnZ9DW6utec7olUQWv0Q3kwq
CsL5NX5he5rhZYN0B+B/xg3lk3GCPO4ZLdPUk/jy/93w4bGBahhbceN3jI94Y7wC
Db0xyVnZEHtPhtP5z9EEtucbo230dlpyQQv/e7c+rTzYql3C58jReRDbnaIhjorh
y2ok9zLgo20OESd5jGDvYzs+R/Aa2LxiMWj/tSPAsMJn+bX3F8NT49XG+8xZCTtV
MGhvmrZ9Z60CkrxQCXCpP1/Lwef3ZbzETJuieFepvS2TrI2nd8zo0ttuS6kDcZDA
jPrx328jlY2a1eWAyITzhRfdxQzP2hgtiXrG1kPOAyxFFAwGtAU52dMySjs6C6Vn
buVHh69qW40nmFd7wAXi+61XB/id3HuXfU5Z5YBonBoTfiA1gen9hCUt6TPArk0v
oJwmo2ELHMX9FnKYtiFtNTpUfW7OgK9bxRqua8cu8AwQI0lZj6kiUROk3ooNDaMP
b8ZrovXPbhpr48wCO8FR6f9hbH/dK0jrRocMFgIr6J0N6NIwqGr+dmxqqknboplr
h032by4OJ1Z96vXXPB0VOQdi/QHWXqFgKJb47/SFPJLf2ApbbSkJ3A5Mnba1/Uu6
9pP/OpEu/7glQkq2d8X0G15L1YuyLtZ3kxfE2rVaNlbZ9YtG3yuWks3vg/8pcU8Q
nN1caEk6TYHiZqn8k/IEmzaOqiY5F4+3yvJscmfAMGZNafXxZu82ZOY+GSC6KAli
AK0PYUUdrZTu4TUkLyBFpT1aEODgTa1unPrqKZfBx8zZU6njFRJi+y3fM0SXZ0/T
LG/+O5znIoEBdkYhSThXKNG4WPL5pKYMTc2vt6lApNyBQYgNuLpH3kGgtqaSdUMU
sdUuUFJJ0Tn+IeqD03cVjph2jFijZ8pOdk6i2UcJq762mjcnwPaSIaIchF8btoI1
Aa8gHuzIf8xF64agd30Y/DVgfpl6auYvEw1jaTARUOmcYQRUcciV2d9xrEmLSvjb
uWxGpG0UYE+J4uTLsRNZyK7QbTIljyj/wiw032as4WM8bWWjZ+B4tjPZKziA4/cJ
ZjXrzQxzusm/uzWKSCLyZax/f7fJBwpXOtvZZrSfpWN7T57jfvy1yjtB6c7j+86n
q9glInmA+2CMG/C8jGuCdBXFU5cHZvQo/KpDTKLQOhPzEn4jt+QFJ+jFwc3IVk+I
WJgTEbtmNW2CwpgMuXDA0C+H2MYWudPGJfDSiK90QuJ0LRjU++IxsItCZ7kpZDu7
LyiT7IEV8bPVoxynraxWm81WFepiFDBadcEZ3Eeo4gwhOfyrHTnvb4GzJZBWgKZl
HSC+KIeWHiAqCiP4u3p+zMX+N1RFWJO6KwoKUh2N4WkqjoPjpUhaA5RmyVOmJdPh
UohPeS4iXNUorqF7ikM3GiGbYzhzRNXJ0we8NGJVMwoaF+53Txsmh2n9jLUFPIR/
RtRJrM1YbKDwry56OPMQKtRXXWnwwQIMSBt3TH1YIk/qJl1GOlh1zjA6Gbb4uE4M
RvHBjxXvlcfsnMY/eiuYFiqnQEZxrsZEVRRkAEXd1H0YsTFgM8f5b6jEB+PeiUKb
b2tmYYGpVkgbm5/+CICrbV1sDHcZ3cHNbfRyqMrhyr7IxWVoNL51UcarQqZhW19g
/Ja9Q07yHOgP1hQgCr8Ar//W6UzoVHIlnHuSASmzvwY2rYOPbeBfVNKXlnOtZQB9
mQDV0BsUgnU/JwvvP8GbDA/HFKYmtONoUMgUUwXqhpT1Y23onrtxukkAjvgcr+XZ
DMXru+xgt64Pi/d5ZVo+s7roRAYY87HctvIjBa05HXYb2aZoUy2NnBcWDnTDgtHD
caAq4Rzds2L5odqEaw9sHcY9cSmZpAiI9o7o9g/OLNnDn8e91Ko2o9iEtUS0aIhJ
yJVt2sHKkEopefY4Y8WTgR95w3SUdoQUMvOpFHt8vncQtsLRuDH1nTI9vhhqS9us
7GdkqttHYQmv5o7gYQh5ycuUoyv3AjzuV4BuywSQtxZVTb2lBUYuyA1vtVUZwVmD
ArwPdX5B8lwGvLMIM98geriPsIYkw9Q9oXbkcw+1jLcaXg9dm3USlYwK/NTkzPob
qmsEM2MXsxprBqN1915N7P613SNBBe3+6ID8Q5VR5gbsYtTMgOTFtox0lhXM1mMT
ucYxOKtca2bfsSFIyBCoMJLMb7guIZSAwouwn6oOymgSfDrNA+Edy9wY1cn7gRPu
HAGJu9mcLNXH4DaRwnpTAohkQjjFVC//0L9BeIQVTztOtdPhyvppRxdrGlqercZQ
cwyecvWYonjQoT2I9iDi2NagATpMiYyfRsEdoOmrlWvR9+JWfmZwx/18wn5VNwVT
0UVF01tkzfT/Ow9ltjIYoz7J/sG1Jv/00vD8rvqqOtiP7wiDEYefL7cmC3WvFvqG
lUYXcbru294kvy4T1HJGyiD83Z8LjkZulxvgkai/f1ZwYZQu/gGZmL3HixCMQojk
E3xE+s5shlEXworeMx/fKUuwnquVEOz4YnLfJ8hPGH3bfe69SzKap4jfYmd53JEB
QRQ42iLAoOOkMeWuU/uVjDEQzvSKkzKqvuOLpFWEu3cxidp7mIpontAt5SM4T0pS
PjTLvxya190Vg24FAewaNbZyHfbFNRYZUM0t0PKtt4zSCKg/v9Z6QKOa73/AnDli
vXp+BzWs9yVYhl5La76eLhmv5kSMm4hnGkwnHpP5xCQqaZq2MljcUPjWOyNvQzjh
yHVi+UEgx2fw3T/+1qOKpxwDbRAYviOM4P/ZaZVibWLjbsbJCVo6Z/ObcfUIPSj1
vMDMCsWSox8aJEx6PZqquhqpjDFyVfqTu+rAMfxnKHVipq8fgznU/wEDpDkU2vo5
1TmaqhQSbghhRxrKv09n0/kK5JhC6+cmOYGZ0vOcxySXdXoQsD261wSP3FQfPi8F
iSvcUm98VHyJ+5wKrjLdBuevfMfaUdjj2PobeISpwgXRG91wOAq0ki3k3PFR6pDR
9LghB9ZI2jQteeuYGfjmHttQhp3fnUQh6aso6Ou5W8eBOOPpmyLj4Mt9HWWEeTWb
O4/h1vLTL2wNGOjAq+BV3X+TrfaWPgmclOeFXVLXmePKN2japPxr0HZn40ls0tcD
7znKFXzb+caLhlgr4HdA7gw4uMNeycd64G5Us7rjNigz9KeeDiv0nuvjYbhPm3Fb
MFcoErThpke1XVnOuO4a/3q4kC9l0yffpVX+1UKowGdQDNZ9fqwHMcG+Q9JW8f8d
7UnY9iE2//R2hUd9pZLoLnrqf67BVeMQAsAe3VzIqndoR/J/aAEe8quE1ipaZ42z
3w6D6bDGBoF4iSA7CWvLnVDn8SMk/teeTFhut2nwZTFB2mcBnMOgRmTtPLG6IopR
0PdVc7Dy4Dqp/D/of5C5412S907iJ1zgpdZGfrRWyVOubaQ1757hBuhPvijUUqb4
vzv4Gr7VvkSV+EfGCq6rddeiWzBJeNjn0yK8p5QauhCHxzXqMzsYFQed7mi9MJaE
Nc70Bgdznx5BB8IQ8hMz7dDjjaChyTGFvxhahZxl8v93YqFw+0KmMhsRLRYb2jGK
jEogwp1UFertF+/KRHjRIfvsI9EGZWYL9pIlE00uwlviA9yzFHL3Xk0lde/W3vJM
bNrPcaQL4jn32YthBhvGAkffSNLcsgQjzpJ/LJ7PHTQErhF9QDAOhIT7qOWodxY6
R2Lw3SqhvYE6sCdpaFemV755tksDjo4wSvgWguebhjIdzOZcZTbqPxfr+rKHM9mF
MPNQ5VCjCH0OawdPKrMOkZ0YcXuP874XP8JwKdEl8bUvYTEiEXGgML1PiuOGJ2uN
1xLuDl+i1oltuBUojZ94LagW0CrC2ADA0VEz9ANbgoanwYlmkj2MPiMzLxEyU026
2u8Ah1GZB3RCP422bGSGNPzWoNW3t5R2XvuwyzjHzwoM1qmsMBY0JmWy0y9KAzOj
bNHrmEv+p1MefnvGTXlssX4XzrIzuGmyIT6Rr8AtpZO5GuYPM49lUBLatOs4Fi0S
jUSjMPADlvGLnpgB1sRsQhhzf2EaJBQ5x3KOFFg0C5xMTLu0WHMf2PDSLQxA+zJl
THGpabYjfnauyTS1LIYDuLORlsZjwRFdMxtyZeSGDkbB8sRiHo5C/5mLUUWtFrw9
Y8j/HhqM3r9cvcVZdr+t35+CBvzw1Ef9s4scGYi6RP6J7DA79XqbgqcAjS4UpEng
Z1FCXOBEGLIzOzlat0m852L0vmy0yoUem5czgs0tGAjeYbLumCirLCjKl3aCfy74
auCPsgHB3Vy9o6Y54k7S+MzNp5CJJXjnpDgt2k9BO8ugaNyu6MJBmHjEOo+5aU0v
yJr6qgLMN/qDILguM50VG2boml8JIZ7CW6N0mG+JxJrVZWHlrqAPBy7Nuq4wb8pF
iAtPynVkwJeQuzsjzauQ2jBIbBVcyANjAQVO6Fo4wiPMp/ZP2pnh9qgqhoAiKXoQ
MxxY3xjtEz/3yfiXgHLc9wa/noEhO+Ke4QEA8t4iedltERR90ER9hP0bTq65i/bE
2w9zr04MuKSj5MaZVaj5tVrbD+RGtxJVeu5eatPkrAIVl5fD2QST5LPbvO+CS/9c
y8yxA/87nahL1EBhbzycFrAup9a4171SmZzKHOVs8pbw+jpOksLX/INQ1KxbOnfv
w6hA5AnMwD4S+mDRhckXYvjDDGqQzVk4IO9LuruSQy5FNiOknZ2PueC3E+9hXbBl
fRO1MSsA2uX1fRawIDC6NYjnTxua4aNBZi7358S+0nnuncQb+QETqFx/otSoRcm2
PVWwBq6SQ1ujOgAcSUpjVllHxbZDzP0BBKju7JYGF0C/pvH3rQkGy/neNIBDNtkV
dWpc7kYNmTn6jV8vvVqK5oaX73blcVeWWlf9L2rMaMQc96Hp7NZskOeeWShdFvhL
gJGP8VF5NUfDOTninAtExB9DtIUFRIalcblK3A6S4JzwtJfBHYJ2UTAfGXTIFRvY
xL1CDy0biY5jlhxvkL/LGB/eSUrTBpkVL9spXxf+FDU0WCFKgHSD4zGSzA7JNM+A
qisTzQXycvfKqPWl2KrKSe9v/IRGUGFw91CZyk3mCRvOJg1nCq+KVSJaWSLTkCBV
EyyTAl5hmnaXPKDb3/Bjo8rf4oP3h5JxMxylfjjlZS1glMn8D5NQr8KdzQSo4o19
WJsGJBQ4Bto4R8nxOMWDJh2oQv+5Qna3JRFXt3kd9bMB/EdZ3GaHAMjyicRss1Vj
3lz/NuY/1ckw+I4oFCT+PQUXevwoc/ANIOOKz0k/HaIO7H9S7C9y9rVeQVuTjVyk
dYgmayRx+I8H3DjHFr22JiuKpk4AFfr8oFVaZaYr9edMPlcGB/1ds9EAt3/+/A5l
hRQu34Kn80QILCf6RNR/btnDLxrn7JFWGJESlGtO7qZ+DnOJ/sxSjG/EHpgemj76
aPbxE9Xrv4QjWaWs+pFXmUrZEWY5Vv4F3cNpPCkdnGHBF9vHtCUOgjb76wc3WH7c
ZcHMgaElBYkf+STh4BCa9B5d6W2ssP/JIXtPNBjoJlOyUcclxZ6zTI4kQQwQjqaZ
EwI9S8U1+PIKLIhltpY4oIqdKQ363D/ii2qM6Y+j8Zf3oS6HvrvDQn+vSHlbt4nv
UlUryf1Dj/yRjyRHl3v/TpvRAEGDNT6SOfx5mFRxZh6tIrzRI9qU6lLUy9C4KzUb
ddn628/5g9omltlPf7kbEQxUMiKjIpxX4i4wtzNPFxfJbny50bu03l4FI28DAvZT
4AtGpP0JHfyB4+d8fFVzHBU/2lfhtwic8Q5H09xZrtIRfs+b0FaTMfT41oQclMbJ
Xlbn15a4aPqW7XmKeefsQz88sO9xEe9P1pLFqZEo7HveIyeu1PTF3huIiNz4vpKi
St3tVA6a5iMnLoSCfMToFqS0+SmIhjjorx4KxTYZ62B+6BnuTpl3zDcReJqfyhaH
qZUQszbdPq7pKZhsgOP9UYFXc2tvfrDC+mMDtKfh6Vp/wj5pf4jVqQIKnjrcMpJU
djKD+6vUfUmqQNv/kjMOtmS3f7tLH30gTh1YH+P9P5Y3fcxDx6CR3EofowK1dqyB
/G2sXgyGW2C0PPmZmJruo3xWnFG3rO5g0abTnDxol96acSifQsXXasoHF6cB5jUk
95x0lyigeSS/iqZbCSGC9IibQA6b+fIyEvtybpocFTlATlHM8eenAv6ruFPuBic/
NdiE9UQo78tnJbmM4d59YNBxJ7vmVvcEOk5/sRqaoa6AHZli4nIQjX7fQ4yEwql0
TUu2rzURTzTlnsrYRzgw61kXOJzQIzWOL81pJN4bk1A0w9W6fUAUATlLXv+bSM23
IXtKhl3S2KewYKNXTGH17LajmBxpuDH/VOl8inqBS355NZi6XV1D5fQ+D5O47uPc
lpjMlN2ZE+D8GOrmj/4gM4AqosLxMjTO0Ve5yM9nHGyxiab71Ct361/kQ+GIlq6Z
uEmrK1K3bgSIRikRGzNM0hGENi0PRCDrJb5qLoysq06+txvMd3ygDjgrESvAnBS5
hZKBR8tSkvlwDCK7BXE6yKwjVPZfMH+HLzBii3GJjXq5Tbj+Nhpti5oa2mb/Kp7M
4+XTlZEtdRyI5zBcxAOkLVE5sim/PCDv+EsUJpfeUxVNp2C7W/O8IgTCcDc4fg5J
vXkczEaPV3L8hk2nWCyzOpN+9A+62WOQALMcR68DuxLVqBYxv57abbe0z1IeXxAE
n2KYsQ/hlblB7ZV38TtJGznxtRgMi6IZVkHiNAz6riM38XEDNulanS7qOQB58uV4
kLA5I06ufbWrlrCBRgZvNCrtV0c0NhG6af9XIMCTGcSCHu5BnJjhL+eQT5D4RX1v
2h431GuGRMr9V/BnwyFs2v8M5abxBKkjRelLdNTtpYCEtt8LGwj6Gd0AAQhJwOe/
mOwasHghqUyFkrHHr4bdxI/6/SVpHKl7rJBRm4KZChtMiBFoSQqx2kKGVE2cP3hB
Hxc+R02g4tbiQaAcJEQ5nNicPUTiqJu1+4gExSAQBF1bVBIwOuXhZOB32xDubPtD
rRVT7m+NtxJ+C90ucmg0XrSAq+rlAT1izqCJ88mWk2F+5eBRPIVu1YYQ8pQ+MXj3
og44OtXxyrusd6AcRFfjHqBUmcDMAA9pB+dHkwtkN2k4HzsOqdkmT5pvJ5qPCN1z
gwsX76ruBQrLhG0nv6HwDedJRkOSNpWew/AB/MgM+pPZUQYON6j7c7m/0/2K0lzo
3WiuCRpjMwK9PrNbLuIxG1dCQrPIXmG4Yi+p8GtcyxEuWNEp8aioT3+ut8+AME0g
vZX5JK4FAWBvHf7MsADyrpF0/EPV6uGtyyv5JAFvEetkr2zGenGskXGot87197MB
TrFhEzX+uv7L42JBeF8wwvu1S/gEj/N9ba16Y/iYXBav6VkbQg3uxttScTocIOyh
BIKtRAqrEg/r7vleJXR600tz1RyBQuKrsSFNAZZMeOhed4Sck9TtSLZ8KCth+7kc
R9HNAACMP2BFpZaClGfGRCGejGlSMPqjSPZ7hKeji+gVaYWtPCpM4S5Nfv4Y8FOj
OU5DhfSHA9NjyEg3ch+U/NsB7D+z9GqcBY46iAg+f6FPHW/jhRsZUOVp/o6VLTUx
m7ljuxMiY8xczdvcNGGSR4jfSHcy/7rp2KZVgXTpTpvy6CV9GXdSvWCWd3F2gVMO
/d0AmD98RZraXQA3brHaw1vhl5oOp/UpY7N1vZAzxm6eGVZxI3d9OauCJO02o95p
ibBTEfHq3x5eBwARYikFbeElPDW8ua+jDVrQHUTNxaP7I3hsOfA2LOIAMB0pmFcj
Zcox+FvkW7zuI7oUyKnXo6DcS7pvGBvg6gnb+1lFU0ocQ+zgTHIkan//Xf+TsqvP
YWKnPChIl+lCANo6lLE1ZRunfGh2370ACvgMzOELaSntwK+A+FwG+JAI0yLiPgc3
Vf6IhNaVrHpfrroxj7Ntpnkacw5gGZQyFeyol/sZK7T77gg/1l1WZD2CepTpOz2p
M3idhjo1w7ouTZLgr3UeeV44jRdLXnw2kADzCdpIDPWOAxxp1N5hDwfm6l8VIg9h
Cl810eUXHGrXUy1hX5X5od80T0iOo1JMYPZi557W8yRIi/viUl0nqkGvLc/Mlcgo
Hdr4jtcR1Tyq41kgk9FE6/R8jLs0phQrk7V6BFl2xyGIhPRzXStHgtGgkz8ptlzM
ThRMebzrpwPZBmqkaAnzKYNbm0cd4V6y5Lys8gZmTwaprJA6gxAnJNc6t8VRSsGy
tx9L3hPPdBO0EZEfiSUdEAWJjB/yLq0B3F61PBPT59O72VS5QldvhwACY1aSpLAO
7DLtaUCDI5RUazFG/MW01fgm26uEPbd8T3R/7gTBTcO08murkCbuqIPeELkB7c5J
uCcfsVea6JF54zUXfNnvye+PrfRxEHOeUXiq2CvfYekj6fFogyBzfJ1rtcVsFIzE
jin/gVKPUOPEbPMSWe7aaRJ/V7EZycycQef11NHD8HbATmWZlar36n7ejCwS/wIE
r4bepY9riKfIfX/0jkEH+2VHdHgfYolwbZuTxprlXkWpD6lXEbz1QaLYOUgA2CbJ
oo6ORiQiDXVu6141pqaPIMZGI1eKzMgUbFGlEbvClKvhfIEsIcNlh8x9hs7QFJ1R
/BcX5iKULYYcduDCa1TVmfoXe5AP8K5Ptb2p5rXqJVZ2VDRzJgCO0H29ow1q+Zal
QeSIY7sh61+M4dOeGWEkisUsTRmrrFAmBrqPnKSQDVXZv30hgbGMdefQE3rUwJqc
HVPZFeSF7JZRigXTXjPW6NV5VujmVxjomfrp3lEcPBo8vrOWTibqnc7OsvosXaQd
KsFIuOz1RCWlQKhr5W47qMTJT8dvoK6s3JBHyGE5qcwd3NztpjWUPvOD+ik1+cXt
mnA5WA0Syj1SrH6vaRSidmqyj7MBWPR+6Ws6J9nunQXQJ+VIIGVNToZHyxG9hT1R
qHGQilTXex3Sy3pNVxFkwBMIQmU/uYK24gx8XUn/uCpsxKGhPSXDCiHDWIYygGAz
N/yOJiXYyBdMfr9PJjcRDoWMUzsz6xt+Z76oW//n1Nu5UZmEfBnBEFf7uN8C/qEW
YVUGIH72xBEJ18LkbW0Ri4SBK8YTjj1C79lxHIn0816LmLjdNylPtwmrwuQkv3Dn
ZPde0rcv1tE+U2HPluTDG4XwqH6cBMUeURN+F7csY7lNigE/Hee5CY4SDxBSHF+J
l3qYN/TXbdflD15NslThzY70FqKJxN0hakstHUaS4PWUDBWk+6eLs6T9sS6vXn6M
TZdZC6Ebf+Yf0RK2h0nNHr7UwYxXr2ZprIw1g4N7uxO5FysAuJzk52SftAn27KUf
yotWHNyMGKx7eygSjwIh+/CnhPjl8C3PMqi06IDSXl88TW6z79gdDlBeOMRy49oU
HJrrXugXhM2RQob3A1y4zHZKf6DRpGR0Fz97OH6KQ1i2fN0nW89K9+OkSqbVONDP
3sxQPY5BriAL9NYHUPaqc3sB6OLVILjAAMUvV8++fuXOJdQ9u0RvgDgtsnJkzeNy
pyCgjNsKci+Bd6PYAgRuI7yxruPb8OCjLz6noSW6Je16pplpzsH/BLtaiMjs0vmb
nYK991xfnYH4TE2VG5r+w2Gd2sNyc86K7zyfcoj/iv+swMQJM+KarGHOFwyy1/xB
lou4xDcHqiFiywj6eBbGC/UWtkTlwLTX0EREHBF0KDvUZsluBmrV7c81CQYK/OWv
2R/CwaJnkq4p+/zDjF/XqSko6GMpoY6OPwuEs5JuOgFeIWuZvGMO5k5x/WjzhgbK
p8DOu/V52TyM3oIuthynKOt7YkhN9ssR1DPmjgD/Ma3O92WAb1opX8M3GMsdxIpy
jbczNsjCz0rfbxEPjcoZ4WFrWFb2WhybhftO/rRk2dGf/21YVsIm8hje2vN4Gnza
rtHnU0XnwOfOJDxlU23FGyieXrybXcN1jUW3KER6+zB6zYqI8WZKMcqcBXmxAkHx
cfsUhdKGNhra1sCH/8RSqZaM8dqkn/XNFW9Dh1AewOQUb+o5TG02bScpru2SXxHp
uFu6jbWDAXJTHg0Zx8N7AyZRtOO0FCoYAuog8WhkDByIdP5Chv8iVQ6cqA9O2gVb
YJxwU/CZWxDGrHauUaDlSDiSzHbaCnnUNvk8NVBMFICt9ZQ1TGjGeY1eEYuqAiEQ
2Sm3ZLfcNiKjkQEo3wPB6XL/Li2WKhp7bUVHBr4gAt6LqS0UI+JTDiKJ0Wkmysut
DxoRK/slMjDzNRTPc6Zsl0K/QYb4iUpeJKG1MYsW+0SUuT28GpFTYjHVLrb8H2DT
DTEw48A9Vl5cGOJQn6a2IRKcW6SH4ivq+i44DS7n2nDuoS6pyz8cmUalKuGuaUpZ
6LLcUS/ISeLHHJUlBkA+2S4lxDvVILk4odF8kUeCs+BNiBHHeSXavLwu1UB3beAk
qekBPgJzLqOd+Bd07skMC1HuF7LhM0EsdX0OpBUqW2/+eYvVjL5mlL/RQzOetjA5
adNgpMQoMNfzGcEqC8M0F9UQp2L05ese2RWxHB7OpmMolVvR3V/IQjN/+UEcsI9u
nI6R+NYe/Uy6G61HOIrsTiVPnaiigoXzAgLZUqmYBp5p9PL++qkjGL7X3SZ0afJ9
fiv+Y7GnUpgwDKIV45GAIX6UXoV0JpcW6QJA/nf8LjOZ9TeQTVGO6LNwHPlW8XZQ
p3tmejt1OauoCZZnVV4OBYndzxAz38IjTynrEgI3Lvd/d2Eqga5GDodLKputLTy4
7zM3xBl1lJK0jmJzH3KPRG0TVaJoxzt6Os2+3aCBkUQ+s9SaQwRoB2+Iw3PC06xV
4Iuf3vOq4vGzXHwhEBsCLRFLnOwbv6CiyC4JeddPzl++sHPH1vhws+Ls4X1AmEHI
KMIi5gLuKntQ2zsaPWa4Ka57GoI6dsNaUkKLKJlsRTtdHBqIAdX6QrnprAa7rcSL
ZPMOz+/7PSV+0jT1+BV1AR6s0AbIevWQZsLKKGIqrrsiAS13y6xquk0DirHgvZWl
djmZYCKnk0UAmPSCBoNmXyNwh4TVGSkKUvg4PTB9CyHZxAbXUDAixxX+iDA/I+WU
Vs33pvR7PjrjFk+7Hs8U+QQ8X/cQHCi/EoFgndzGhI2l2ftoqKTZz8KUg0XtkG+C
YAdAX2x8/cYnRz/HCxzOzdaeTXB1Eb3Df9WZnre0Q9ToAX0DEZtw+c51z5oFqLhB
Jgt5tUeZONNKk6ClU/CFh4jSIPQwXSgvc7WiKkynOmKNarscbzveNvJoV9cQ7cfF
N6QSadh1EiV32IMddIBdr+qasyVcycoQwCKTpIChjViEvJGIHacIqmhE5Cg8TqGd
3GMwBgdJP3UM+MbUFOk0jS+iQQrK5akEraJ9xj75WvhJQP6uSXYRBZbuGyvx/uUc
X1ikHkKmTJWkrA/Y8OCbvdIg8RF31JLO54RRiyhxjNOtCrsk1Ze1bPFJSP7sO/76
gSb776jjXFXekCfUiG/wimsCo1Rh18MN96kl39YHyJewm9UsKumuA75VUYBYpx7O
IyLJgTAXdjTVG848nIhzDhlYP6yHQdgRYMPE3Eg6ETNxBjRgcdpzn3eDUOLgB3sL
yQtmvqOc5wdH1l7+w3lfJRRnjh9IEPfAE72X6Ufsx0lMYkWjnZaO6rSo+wlx4pct
WsQWEy0h0au9sxcGEsfEVlGQdULRViuRze/Q9IfmErdHLRl8Sw7KTKSExQPEXugn
6a+THx0nifJJ1hS6HgGf2v6VZ6U2+4fRViKmxTXelPEyTgOfIse/G7uBD6Zu7zaS
ub86W7YRxixlFdtrbrUiIMzkoPIITnzgY4gMuuykhXsa1ahhTgBP68TezVeu6bjt
6KF/sWObpWYTFstqxBhH8rCmj1CqQkfgg89QlNI6oUVImDcFuN5EubiKE0YvjgJH
9/HsI51m8ut3MwEwCvtLtPvTPle5MaiaWd0yBBn8/4VwewZ4SvacYDj8loo5iISo
yluzzmv6uG+/o1nTO6Fwpkj5zsu4yER20TZ132tjpBeejgtyhHmTvrbO85M6Ip2A
MC8pJHxbOw7ByPSRQewnqWvi8rRifEmsK8l+Ft5IjxWlcNnWR1fYGtdZH+qS3y+E
n7d8eUV56RuTIygsyLE3S43u2D5ve9iTRGq8v47QH5aErRaUBY8nfO6ZQhOI3xhH
6pXamqbkTh+xBaXKWuqKx/lC4FbEWV9mZwpNb0eovotSWoyu78I5/Vsd/hXybiTY
rAvkc0ukh/bmeikBxUD3T+r5mLvflubdz11pLOyPbZJUxOhkhHwlP9FzV50qvr18
9HdIS3GNWQ6nlEZfwyzXjONV415S3aHr8jyhercPX1lLsHz0ADvwQ5OEtSyQworf
oelRooxFK82bi2OeqY3Lk+YU2celeOWGTRFIbsyAIBHn2Rt0gitB9yBivPAS8XA5
PEAFVOnO8jQZXCogyDVRecXKLy7wjRx64/igL+/9L+zqPsFyvxdLaqs+xq/RvF+S
qvJswVgRyeAgeSEQDWMXx0+LTzCC+kilGn0Mneh5gJ3+bpnnzhG3v3vUGYkJExWS
mmHhVaYGznssIsfrgl3I3dlv8/RghltSpkU4tBry7Mh6Tsd4YJM1HNuGPDrGU0rI
ZLrkXpx4NaZWm9PRsYzbLaFqvdW9ZCswcPUy0jpcBltNTFQeUZzfAIUOkWKJkfT7
aJtv3j8adUDD8wDi7qwIEhZoC+Wri7/Up1Ta8NMZhbnOSL2RrqkRX0zssfLHw+Po
FWsQH2oQbxJQhkN2QATWlD4hUFw+0OBqxBp0UKKhvCsLTNP386yC9x5fwZShuFpC
y6o+VACdqcSapfxYGosdnYoQur2Ra7d2iezhbZueaakSZ0HnnKKmmgilvnNT12at
ob0Zah1C7n5NOSoNJua/e4DO28Db6+EG2WmvolIc6gTvHF2QJqECqr35j+hPLeJI
Rd5L7zzD5cYVibxEHyIvTlLwNL3sSmAXGNnHicvSR4+yIp0CkRzx78Jlx83T8pVx
0bn4GUTb/fi3EbQS7fQ18EyIJY9lVxmIRNSfBXnB9o+hlwL6GpJ1+I2evMlDo6uE
Ef/ehmW92Wkl5Z2lBJTPyyUtlcwqFaKOJW3Ou4M66UisBZBfCFq0esHqB4ZUAuq+
kkXW/1x7hrGItW0wHEasSgk7L63EE8GfvWtSeO8iua8s8ULXF0Vye482gW34Wxpx
Zdsz2AiD9NafBSkX2E2lz4XiHR4oiCViAstJm5aIqmk/oUmy3l0wV/IebvVZv4Hw
9jmprgV/4zfKM0OAZCaKZ1/BTC7qc+AO76f/B6olop/zecGZhZ0Wh2VlumUm37Ak
RmWqI64EAiOjW+Tb7370CkY3zRUWDRAn5WzwOv/7c05QiEkfB+nZsI4QTE9f+Ep/
OKPm+NSKUj3sb8TQB1JQX/K2WsI14Z7OvELlN9ej4lxSxPJ6QWDVAMOVPX7Ur3H9
j4SOh1kvSN/BhtbU4sEyw43gUxmTYaUYHknwKCBa5YGVIERs8JiZ6Ur6l2T2Jh+P
PVSS8g9yps/2anzMPEublCdObt+8eZfuqrlk+b454pIkmuEMyRTnro6kLhwtUXTr
HlzfMbMnLq94n1FM2dJTnMRG8TovRt67sb06NzgouZMNgK/88UNWcZUWljQo5IIX
pwgc0RR10pORo9LERP2CnmhHrzXWmov/G7Zgej2gjvhjV1cgsV8doe3ruhjQw0zF
LY3gNqwKohYTjMx+JEkL269ONES2iju9aJY1pNb9PpFRa/hqsF1ARW/1lLr58oMV
UH2hriCxD7w78XqFAmOuw1zng5rjFTqK6XWj/+Swv0yNMlMdWfwH3up6uOrDx67V
kR/LZCKmuds7L3isyB/7n1GGqL77XWHba8jicmKQsK+w4umKKVZfpWwRa80h8g/O
1Ql5iXxivh4WxcKAlI0HeMXQqZbznuEejzPZvIUfw4z3OjRojBQhpu2DYLWVS0TH
fgGJMF4anzMciFXVT/f3NQ5Z7C8gzK4TE2hiWzsVDlAGbnC+AtsqdUARjj9NSomT
yieuJ4vxNmTKFHV/atYb0ZvWETpfkHVRpkPo1xMg733nBSCJqwOewEnGIPX4ZaiC
e7nExGv2NYQgbv1D5vnpMuncUmuxwbMvJfqD5h1dq21YrOL5sdpBjRvstyFlwgvd
/mF0WWKQadS0ro2JFny0Pb4x6zvU+uTqcvqHPFml2ebe2OWzGls1HtoB2hSe3h6/
/fZOcCpsq1Sd6Q86Mrdz1VIVNBG7OkLSYO4heOAOYcnCzMRz+tTGrxV8J8JMOvgo
+OwMLOaDtmsIuGJtsVS/jEELGPgYs2bPVVuw8U0RCB7RZjRl+6Wrlw7yiptuozLZ
1FKcxoAehX1/nLxLSiNGRKy5kFVBxuCIzroDVaRfyQWnfcAiSF/wTnwri3JAJva5
Twlj3/lPqQRJ6iWScJ8EUPOVlh0Qxu5wQ3xoj+AfdQpeZTV153Eot6pGUlQIh6q7
7a+drpsyEZxUe6ABzwm7i7ZILUPbUuVpddADn79hzkru0Znqq0qfOj2f1m//P5em
Wp3CgqIH51G3A/Tc+uq9pzzDP8SAhG+pvNTO5UMzE7Yv0uW3uW7f0i10ZiEjopip
hkZ6Mrd5XT3ZzlHcxmGEwrKp/LTkVBFZxBa3KfLP6TGgCmQ6QVIUgNQRat9O7mXn
rRcwM/+gN82h8DlTt2KNC7JRSgJKr1WS5/d02KisYyY49sZ1kWexicBt/iDde5+s
92U+is8HiEk73S+V1Df1iIuJaz0eM21kw5VPJ+0kqOog/goroMUdLI8bxpT7VrBB
/fv8JLUOTId1x3xb+2zL8XEysY9s2OS/Qgldspe6q6aMQmVjyiNW8TtDPZ0/60wD
57jKcOcGIMf4wsmlOH5JwUkdVuqYk0y5JTwJ4l6z7vu3fiZwDQxpmb+r9DhT+bHb
niWQ9MO5UnIzXvLgcKUnvipcksAvPzsWp7mi6fkhCbfkr0QrwZerNaoU589jtI09
7Ez5hna91pNmhA8vt8YcUZyYzseyhqs7OVALBhWHiT/vCaQJ1/XGAxB4VHWTfVRf
riJVaUs4heehW9OpyQAna6RAk/Gdbk3bcyJExB/++Git191nyam7hxiuW7dY8aDB
HZ3dklFX+4smB2982UJML4mLCdclTO8b7L/fh15vp1erHBgJjuyblK0WkyZecQZg
9JfE4G4WZX2m2ypDOoh59J+wMs2EytnCtxkIkQF9vqghqWDmG3OfFwLU8hA22ReQ
m3ckDfmKs9+foQYCsFOZRJVP3AuHdictp63p1WncHOMdgaJ8f8pUSWfAokrYeTIN
+m0owbLwevafSUYGbD+Wq3QshL4I1N1wAsTcO0ROzIIv846Fjk8ztFJ2XvMZH0FT
Ky6U/Lvk5ARlusdSdZW4uMjfOb3tIcSIgHO0DXZNaGliGmYrWL+LD3Xb+bKO8vjo
sxAEM9Ex2Jfq3s/GE4vg49yOqErz20aRuZDTqRyT2nB6sBEtu37cf6w3PG1oSvCh
zOFMfzVsd8t+tREFEVvs1WIX029jgex7NtYMEcRfE5dfXkkYuTvkVFkeXEPkwUk8
YxqPXdw6Kse409rlW6UbRWGU4REk/lPdGCG66MrI08nZ+MAvWa0gTvV2YPidrDLw
UwAJvBERoSXgb7vOY19RJruezFP77CZ2Sp5Gx5jkvxlpXXk+pWqQw8/DWqkKQx1y
Z+ekJFj+CwHlhISWI7e5rYB7GDcKZDJfVLoIZxHZce/g0z7F7/SufJEpJJskC0n3
giRwn/xjQXyHFEEttkQDNJRrlPfYzCDxnhTfVW+p+8H3RTWV6YoY+0vkRpv7dswm
QYyS1UX2TJiwAHpp1vFli+1Tlyw5sJAVz8Wekcjn6Lrq2j+qGXsyV9g9DWtmnJ0Y
m694KlQUyphR25OHNzxTPoMk7iU6WZEnjhcKe+taPJxSw5ejZCI5V0+TUTWvzuX8
FR79/wl6f/FcNtgUjuNpK46gXyy39IAem1Zn/GDZ7t2QpDoz8xCKqEF/EFhwJH0t
wpVHF4hYLcdLbv48DQrhcUmLtU5Tadi5oO7UdKD9FofAm8wYwQVH1gJi4VI8Pxc3
2K1zbj6xfpRIN5oJvjbW1Y1cS2kT+1/7W2MsOcO87DQ4lhdTAcBZtNYKuNx8zXoA
igHUrjPTWKbvMa3gbCa3U3574qk5nPzt0Isu6Sssq+LIgJ5j/ASBSvjVQaPZHHkO
ffdV2Dn35FPomCS3ucMgDe2XkXyBgvq7Q680Ywh/PwUIAOWJqdcjA4c+7L+cXsRl
P/0OYx3OqVCPY9t0HVoLCYXba7PXK3JiWrzPE321P8VA+FbB+Q7F0PQSTjekemL5
awMCpxBScNyJRIrvt5UWySGkacDAh9d4AjUw/PBUr+jSO2RJjZ/DcCU8iGFEoEkv
IaWB8ajAmynpArUFlUjDZgUOOScxUHtGFnvDB7RPw5fAxSx8No2ZfU7kzzkJ+5wl
fBuueeRMY0y/x9/FLet+b45EwRleqj4JYwLMN9drUyYQWpD0pMmQLI5bHbKHA7Dp
4D1/pxGolRh8pAdNjst6BgiBH1y0SR5wEM1kHskngnbpV5VH23rWy5d1d84SQLio
vDpyjUvvekoshebs266JOwxjw2J6+uw5k8Q8Jo2uHV7/PS3y0Hfb8xsCpLmTTIRT
fIGt3p3fwlsqcxQie7ylJ4SWjC0jnmFhqUTXAUwp9yER9T3sLhWGVtWwRFAlHdIu
mKVKkSYuBJjqDdx3Ba13BYrT0EQrCvMbYfvSzyGLvwp2vSbvQTn4sGz4iXnP6vRB
fBOSzy6yITX3fdrbmtqMXlYuHtFatg8Q58KYV7Y5Uq/720WArHUkBuZ6x90SVdtO
y1ztGAaHw84U0cpfVV6bKOt3aBdIuu7PSzBIXQRrCedrsgGS2iOGCq+/jZeg+nGE
1zbcGli+lfpZwqvGjy6NaZoGVSuaaWg2JP4bXC2czgcRt3QX/PAndB0dkfymNH7Y
J/nzPP1apWF4Ek1VHrSL9GboIP7bW6/vfLkdnd40lqFYtEM3pCAs7emZGozxqIGS
427R7ldK4RDKbRl7nNmwDJB5r9d5udLBAAGbjhzuNTmtx50S4FzP2HpV9zIdjWZC
8QBeJSnMly6s9ZhJy0P+MpRq7zN20Fy1BoZYekMCpruhSDy83u/+QWNqbRm6JJnO
VIHtWgVrGFQXBCApnnG5KFT2PucHXAnTTmT/kypSizoDPcvfnaWkYIT/RAzl9XYB
XIRp2AOaQotzIW1xPMR6a8o0YX1QIUTUlWo1iVTu0TuxDpGEk4AzPlSPXVCXvZux
po/Ei4EZ1lPtGAxMmd7H/EGQ/dZMo0AOsE7gHkbyCeM7/T6zOG3BKIq2HJgGhNfh
03dpeXJWEtixou1K41qkIX3u/GYb6gh3V3UhHWVz5iF3jUi3XuOFa+dEpAOhfeAm
UdTM/ws9hCIPU6WDX9Z7DGMmGiAyQNi81K6nsXUqwijkZ7L124UKw1yTuc7Lj1Vx
i/NiniN2qvyTviXLV84U/KTHmdyDcmfvh4yTB+8qDx0NQReotPOMyO4oT2fmhIzY
V4rrX0oTbEgijUu6BqKFvbk5ufooHKQcDY1DEXFydIvKj9iN27FoVUPY0XpRb1d1
X304aEDZzk6YeftCunFwo6N2qFserakvYmC4V90ENWoZw2ELW6U2tmdl7csluQXL
M7cs+em8aiLfe5p3b2uzrxCsUHEvM6QEiN9cvHee2ysG5yx6tfv0r2lazKQJK2d5
rq+UjX17CVEl2yJJI8mGjpvekFe+cetEAzGQtawdzr+yvdNcn9LMi65KD/C1oZ9q
sWTsEshuvqvrBuRW8+t9ID70XvfWNIpU+SixPUx5XLNY2B38mvfZhI7VnPmGGm0q
BD0qpIaMXErCVkT6snSO9dZw32YYrM3yHRXklJb5eeECzq5m4xq3VGzRhc0s0Ar4
8nRkF7EicKEwqm9EZMlolp+8kiyaPzjdR+Jovox0N3GuM71UT4N/7HLJ0kzH4kxp
IFpV4wDLhO7ifVgCNPpsH0eU7qGMK8OPxct3Sm+UlhrLrpeRqE0wgLYD56XHlN5i
0mtBjj2Uip9hSmXwRUs204jKwsDTPBpWbwgkP7SsguG1DhnnLw4+7uO6xHB9mdP/
qPL5JLMrYRBNhWEKVw0mBiTE8BcqlavVi3Xe/3EyUh+LnQiLSjS1mGHOQqU06k3s
O+39aWcG6kC5/Sv4roOAoTL87L3na33zY8O8Ag4+Hib8pXbh382RE8sU9tWk+hQQ
BqO+6M6PtfeSL1aoXp1kWGkKgC6JOUdcVdeocaK2Z3Z2RWKg32itnlWRfOixhSD+
X1CLAfyVkvn0Qum0wNy7h4z8+2ljuAxgsWKZMgavvoPF1o7mFH0lyGjISIm7HISS
Qy6GdIkwOGR/jA/1Eo94BQDA6wPiui+Binn0oJ7GQ/2MK2MDBdf8XLcuprICbcwC
okq7GQbkAG1JiewnmHrfdHCybRzFGU/ttDbWYXKJQPA8WRg/muMpEEJ0WUDKjt0Z
OF07/ZpWw0LcqZ5rCsJQlTo5pHhQcRKOfhD+DlSCo39FsJUeCs2lRiMO7h3C+95z
h2+dyS6iEwxfs13/0x8a/RTRM6IxsPUTx+OJ4kvYXoL7sqetyw/8gW9YlqUO0vJL
zV8DrJ5MC4sptk8IIsV21WOoJ8Lqa2n9IQwd7//obVU7X495ccxNrGzOzAj7zr/A
Lma82dMLE784FXxk6qT9kSJW4o/j9u+hlS8KaxIzcssLtxfUTLTZCrclzicXoifj
AyhcKfl3/ohg68O+QeDcePgJQlxvQoC1RplOEGfiKYStf7YxKvBHZzdvzWBVXazd
ydLDsp/34HltbX5eCa1lu6YQ7v8Kt8IOHTLkPEwrGJNiOIiQJ66/skNdqn7RF4Dc
+byGi+MKY+JrFS5rS0yyscLcRsEPjzBT2k2lgqHIlkWC04PTU+8n9DbHex0jyTRb
6R05b7PydXK8+mWl/jAT62qx7nSoXXjpAlWuTEs1GZ1vC/kEbbqYzDLGZVj9Pn2x
ddYoVNOpq20Hxo2/cmAQJmBbyQmKDVqwc3ai9EfofrQdYVtw2y4b2cEZHRq/Vmds
zSI3nOX6LLFWH0ncTHEOSUbJ+Kusew/cAciRC5u11mhlz8PXB9WxmbGcJXSFxECe
8cT9AZ9RvdQ/ecYCQ3QMVDWWhYyEg2EfPZA47YUQ145z7pajVLBnSFHMpgvgyWti
FXmnv3icxAR5ZUGJ+fqrvyW4zrodOro4nfzKwVTQeToPJSkF/c3FlsBjyauwp2Pt
bMSXHu+C2IcKhqJQ16mhGJ+jSI/KzS4sKxDkCvJuqF8oA3I1wj80nYCAMBuR/OkZ
eglXnlQMMSgH7mZj/0h5HH2jzsIMVLJIY5LKdQrXHV9Q5/2ZhF9b2TGGYPMmT+1i
vvFNjbBsGmgockdQtw0I0cOBHYQ4uJVnrPxs0liLcoojXiP9f+mMz6LWKuiqCWJn
H2hBZoPUMm6jN73Kf16ZwQCW0wqP+C6StYpfDbaumRYe41OJgi0qSOe8PaNJ8+cA
Rfemci4sqy6ns2nmfDz5Ep+a2m8/gn2x38gjJDSiwJ11ZY4KDDGT67gfclOSSsdB
lterWgPYIDsgsjiLj2rC5tS9HW1wWAskRjCHqAo3e2LMJMNXsLdiSQDifw5sOT2q
Wp4C2X1WhoAuutjh8qK2YAP+D53nzQDlOhrayh/3j+3ryTulMaXPFFO2khsVBHst
q71ijP4NreZUgM6MYixu7pALy1vKoXs2PHcLaFl4W4WBI5WLy3jx6xRdzk6zS1ws
89cPJ2xaLZabOU5MUwjLaDmNi4m9201CdKaWgtZP5bgdHKXB7GZRJTRUYPAxb2Jh
fn0b9g3bncNCULrQLcEQj9GCXNtWWxCpjYq3dA0KzIzscXpUrnVW6dkdH26IcX6/
xO5XNZrckFw22oRCIaWYNizyCul+TBuzeChN2D1WRrEkoMzgFmrrjhPN0sA+7NJk
ff35gPXUL5Zx0HxAhIEP66NiE8NvpXPSys7IcimI3olYQ41tc4WGznbNh3IqrS3p
3jY5GQiWMTJpE1LBEpfAoP7amoM1IpSu0uFi0GfdqjfOxhchQL4pYvN1fWZIFuvo
yrSzwcdElS8g0axlfwyjtdCQKBAuH0kmbY3zClODKTFOtwPIH2Az9RJVI5tAg5DE
6NV4KEI+ufo1z6q5KpvgrmXMri+CKvirzBAnAiiRSuDYqBzNcmHnDifadqRuCQs6
4UqaQkBvim2E3nBTMO1glmc/tQRywzZnnl7GVp1xMjnhNnm/RB2xBDMH03f9bftQ
7fjS2BWz3XxRJUqPOmCRJaBycOM16tEj38zF615JE40t4aJKrRmWSaHd1xgr4nMV
qXElkgYpzeTc6n9+rGF21gZwHYxL0+U2Bz2GrnIcki310A33c95xv7GFmbok/DzW
b0wtpKlVpM9Zd0xN9X+wElEvSHNHOl37B5Q70bXnj1iTt7AlRpOAqZRN5CgbtFuj
E0cvXg7gD5rYr6JuazMwcDBgy9YjyNm2bQUtBZ03o/IaludIyTH+JjgooWkKF6MA
+YmARPprRMBjzve7TPdwX9dcVzPZvR4zDFi0BQQo102d618QWEtG9I1gLHsngmFR
wluNUHrQMJOxZLBh9AWf5BjjQ/qy0VbtS8R1DdAr3Td5eVKjv+YCWMGUKbrCGSK0
HiNqAROCi0gwfzZ7dToJKhVPAClX0RuKP4odSVw+FJnW8MmVOC00STV6IjFg6RBz
UdNZWKXhIq+Cc0ADBykwA2gYJD8HKJZuwTie2z/pEfJJmN29FEcITkxhk+fKL3HP
9+7UkbMVRHGsT7dUnyXClzhIhLaAMWwxHpMZskP7nCrWBA+POSbsiAoJvuLvbwv0
VH/7HOC2AgqF048EHpMy3pvZKvVhAuwvTLR5jrYtLJWjEi4cznDXaA/VS3bChquM
+FJy5igTJWva0/rtCVqk/yy8yonpEHUL94lgdKtJXDbBG6up2S9cFxvSV0vWne0v
EKmR40FBqge5r3NZttcGEE7/6nVoyxvPOkozcGRTF+fGHanBUa8th7y+PWU5l/r/
pUa6yT9VDrYuYLAOi4vZ6H4C/JeSOYz8F2k1ROpVhyFjluRPA0QhT1FY02a107Yr
xhW9suqDH5T+y5GCEwKi1/++3ED3S7Dh5gDupqhhuJ4dpTiaIyKI+AUa+3ykC2uc
E4EM7pUDJPWRsNcbxpQO1Yug6ZXfxqCshzdgBWbKqD3VVZ/pQw6h9RGIZta4+TCX
r3ZpCAjJmiJQoWmRY3SQL4Ice44dufb46bzQKYpfL274OxpANhGmssq9GX3qXoju
dngKaVndTEjxCvLTIy+RSyERbClVdiybsPs2BtLUsEFixoVDvRb4kjg+ZVX0pGYu
SMtGJ0HDnihmAmFdbxtjkv3aRvJYtuNvkvK5vb8M5WM9Pl3UB9aysi8WWzApwrJP
rmZnvXFFdlsxKoT9RB2yH+N0pimVUiPElIWY14iDHUpOIc/4F2+eEigAIs2GDKvJ
7NVqb39rmNh4+kBDsXL7kQMN5QCflEVVIc2UM90h1tTvfK9OXgHc+4eCpMnA0ldw
jeU5YqNDs5VgUAeGfWJAn8b6i4KKFkSkm81lPKJNfwQV8gUk3NOwuqrRh7+N/a7e
/Qbxk1kkw0KvkatUJxn4l++BG8vJZNVtW7zgybX6mOn0Ps6AWwwCzrnix1tMnU6S
Q3StzLCShF2UL62n9AKgHRf7gUptQIj5fC+CFZKaN2vRRPvplXu+bHVPVknc9vNP
F/PufCPVKI5SJveBBom4NroHIyGRcobQoxBRlnwnMDPMP9RlAdDyCIxakDCo6gtP
5rg8bOHI0J9g7TKd2LFhT7m9TlXG/gORGaobnCrp2ltqCjfiX+CU07Bxbd7zUSfR
a3RrUqaR0w+htd7YaBeGMb1o4pz3o4ugV/EKMym0PyIdLj2SGoI6/q9MUHUcjOg0
6JBb17eJB3ajsGKXFVb9nF5Ufm4Tfux9Byx4EQxFTtiCHKEkf19sKGM6yxR2uwad
3ZP1N2VCkUMi4evfsjrQ3z0WpJkuuJTnPO+OuE67EQeHsgunWJlh9XwvEF2dfFbt
yRxW+F/kYyaxM17qAb+qTsbe7jtVgTdf3J+VovzZIFtMwijKFJdMejHr4/XWpDNC
JxLFiJJt71KHmanRs4RgSe1tfLYQ5K+TQPzKQy3LUVJSpLFW45reCHimYV0WH+2T
bnCWOlnZ6xTVEVAUeC17N739YK/oSh7f+bUzdQ/SQYP+SiGL3IoJ9rJSE8le8ufP
LuI6LFax9pMPPMBjXiQ1B8tSL4g6tu1RYxYIORUAAN1CFOhfaiP6ov+65Zc+S67u
DjPA1IX1s4GOpKnBwHZORo99t/4QHb+RQD6dPcMWxI18JAz8VIBiF2XYqQpEu1Zo
3bQAFS3y0fuyMlMHk5lC+Cma6w8XPfLHeU0Fockc1EEGfAhXGO+L+z/9TuOGOwez
yuiLGckoxJvuuADnFBoSLK78JRrFpHJnSXfiC1q8ulOFNn75kK8HpCIB6LlS/Fcp
w2uCa8gYXmqX2AOQVF5zkQYGebsFEvWjtTY6KRVaKws44iF2rNYtixEGF3sY2Q3T
eWbQS9KiWxzdJqutemuJ/L34oXtA2poUtyq8m6zATakJq06jtzUKqgibKGc4qaGV
3TVa9ZTD6340JCKSTZtQTONrLsVE3/jPAHZ9/TcXwZEsVbnn96hEao5insITW5O2
IimB2HQK9EzaWd6l2aTwsUbpUbn6lsucgnXz6TZT7Yi2wYD4OY6xeGja11OMGqpn
opQd9hHh3grt3SqZ5DCOddgcDRt82RZXL5qTj5Fd/PGJTroIZh44v2dnRy8OcZyb
BcMkJgh822gnVfzZgXjcPpqifJyvI5J+kazcGXscqBuAVAOwOs9hqr//EoxzTUc8
SPFexeq+eRlCCHpPwegYd5VQ/kaoBivbFk1nG8D39sBh8ne5drooucdo/MNc66kh
1u/BRt+TnHx0Av5yb15XA/wUhbn0OXFoZdB3BDzzg0TVPqqZ6AU1odAttFEgQmXi
9p2lLF/9v1S1ymnM7IQdz1XGox0qsizPPaz9EBgmdIQd6iGdVXnjjqkCpXAFV4vM
Ubbx+ZPmwZx7nXO6P+im5GYyKa/632e/+vhdHRyTHv+AcUH/CH1Y7utdDi0J2ei6
609wvx5cxtLo9JbQqtx8tASEZ7ydg23hIa/5eDI0MRV7yShd4fxM+y3FBVYeiVvt
Zb2tGJgqjdo4Qr46YsBjvQCJyUnmMtoAlDbSMfo2pMmLuvFDHYI+iucd50IL2Rli
iw13lf19ZtEbnQNVE18zjwK5UHzpTgL8ycv1sswG6gAiJKx5YR6nl2uPhvg20NDm
RVBZC2wr+o18XpxFHmuKx2JgBlbJdXCp+UDwNaUtqrADc+sp0cpf+nwaOA5TPn+O
LcIX3QOMo46x73C7oqB+EWgpiPv2TJF5pvkRo/KfzDuzycs1y1ddCq4q/sMZyLL5
bbphUg3rZfCPYD+adR1XXnc5HsYz+d3S8ftAN4yS2aR4VkwKQ1zuR4EkTWZGkwtz
GeRmHIpMiAF2nQorG5qjEtwMLu1sj6JmkLPA7VVwq4NxCtLOtZnU458IC3kQwUir
rqEPTEkbfPrBuxVJPg0Z985xOP4vtCghTyG/WAb4H3cfrayD5zVvnktgYWIZb6tP
fpfN9q5wTge07gwiw777Mj7RgWWBEwBLDOnTgBsQhdeFgfFAy/EZYjxDMARqBFTG
Q+Yam9d48r9+FWqTcj8YTOpGCbR/wgtuzpJimf75F3eTSEjeHIXUUGLS6FQbL/li
uEYzerLSBfrUB3j8R+nCrGVjmiF5pRw1fhW/p77Zpyi4SoyaU0cD0NLG+/t0JMLy
4kqi3fS/HacDwcY2uWZhpyyJT5gXDGDAVhF8m5gENsC7h+rVlWLZOpoc70T8BnVg
1u0OJVPHMal+OAUpcxGQsCOUhx3PIDQ/c2ufwBlJJtMqUnf5JolIkswUwLldumOU
OF7tL0QB5jYSlIDIAylGgvAUBRMvIRhGj4P/QIq1jXhTiP9Fsa6I2siUVpGv0wVY
8tImHwzHTolj3WIlDKOVUS9xMkI0N0A66pJtkJ/lKRwmBj4tDck0bNWdZxUttxB+
6+IKlDBy7g7P1nA4C7LjtAjIroWkaUSb6BI4bh4Kdj4we1dyZuboAA7HibESnhQL
wcpy2mwMcajte0mU+ly5kWpRxKLy/K39ANjIGP7NQsMnbIM2pgrF2Fq6B5jWGXIG
EGNPxda/d9eOqzhD7OClIvyqAxT6nX1b/+ySb2h8Hr6GS2XHof3uzGu8/1k/9DHd
f2NkbDAXjThDmZvjlRn/MCY36ybLCjomKWtaiei+oVB32nQjQXZA4CBdiC764x3i
m+iO7sYmakibo8vQqTHP4QVDMS/HYTQGY+Kaed3Hgl1xzYja3udBHddnszwUMNrP
LKCV0B5lUOC2Aomu1zMx1xJohRzDNw/tS9kIp9OtdnRjO46vDUOfHtMkiVB29ws+
io25aNTi9V0DKi8skGfLgMT0at/Yfbyr2GYoE1Jwe6hkULTwnuZO3d7IIIOx/4fG
PMJSIN+USffafjBZsKioz0S3A+9lK2cMln4Kbvi1TotDsV11Th89scwSR6rgT8I9
KNJc4eTHf+x6w1l5unVG2qetEOjNSU4AS2mb+kX2qcYLbFUWduWV70oah5ui+TRn
0elf1d2/T+FgauzBC1A1Aqe9geWbfLe3GPMAj3VLZBfwu8Qhk7BxSwQciZVWg651
dj69toBQK72tlUzoYIB4bSBPLrlP1k4LuVPyCMCVYrDFEm3N/9uFryzA29Rf07z6
M7vibHQE49UghNJN6LkHncNEqvyHwEejFBFOaLK3d6O6YFGaHquz0mmM+UeSgMwA
G3at09HCEqg4HpVIS6K91XZAJwRtC+AptdXl4aAy6CODog3Q4vQInXyKsnatU7iM
Pj2z3ibV0g8hMDLPxtZfGEFqKPlJjk25SJW87Pa74MjJw9GNIq59ioqkt/ygoOwz
VOg7N3hfUZ+g/u5skFU2wP+KPx+cMGf17tUtTGUhP+W1ResygGprI+ugnievlUHg
WjEcLGB/5tXMeX/K409f2Km+IU/ODgS3xaRbZG8nLGG4q+l3N27/Qq3qJQE+26jl
tX4mKZ6rMaYjcuDR6ieP+0bLjjvj9yK7CdF57MBSOQI5z+Cd9uITlLXnZT5yPi1n
gGOK3RwbrOorPTGCR1YMegl3okLyju0/3H8r4l+NbtIAOOPbjF6yTKLY2F+CAqbI
HxHaEeOob9mUDkvE0xvROLjQzeYLF/d3C9dwyXIZ3tOl8VEr7JGC9XI3ZSf3KkOx
levHrnbDgWVPFGcXXEm1MNcSV7fwCTWMWkL5THdJ95Tz/oYekZtTG3YjqqeETjuG
Ayhhn9VEMyj7JeI/aELBF3/4P1WpR5cVnRFgewF5UlFfzZ0O1lKv/wM6e1bKorUf
ZXpw4ylw/bSyV+nK4DSsuxc8eNd5Mwjp0fp7+K+8vmYpwkylkSZ8HTDtt9EYoc4X
HIwWg973j8/uFvSyDkXPn1q7HrtoiM0/58Id/UnFdI2JQ/8fcp/AZ9OJg22fMJhD
krBSL6T+XQdFe7CDEL3DIoTkNzgvH0oSFYiPeNU0drYDanZap9upABv1gb0n8gN7
VxAZ5O/8NS287Ptf1QZ297StArqVswrxoGcPt8n87Y2OexPbABNi6vBwAySIKVc4
+HgSRIDMyOnZN3TARy8MsxxpQdpb7Y9nJvkS82TyRdDoxSSu9FyfAsP54TTtuLyM
/MXgZlu1k91giMSfP3/iPoT9PRs7r+F0iDtWyqPFVs/4qLNrV5oICVFV3RT6BxRD
fgNDz6//s2reJshZTopgyWjp4ihGjtNidZHDeB/MZFBJSq09WoPXzqGaczKjaGhH
rkezunHD2y5Wrc4QAf3dHqBshoM8OkYnO5TJWKlZXIKchTM4rjEs45nAQK4U+5Qi
vMACz9xXX1MiYV5A1qLSQ8oD31O66fuNUVmPRbgPsiNjQuJn7V0mtS6RX+mAaabX
oOl+9oEQuzESDdoSdDcyKaRMaQWaejVXMBEneMKl5xBvfs8NwWNyVOO8Zv/ddWb1
r7aORn4V8vQ2Hqv+I1i1hdUsP2D5T5uuZEqG2b1ZlRJHZV+3IPmGmDVz1Hiyea6k
YeDf316FoymYlEB0T1QDtcul+FepL0Iv/0sev3QBO8fcZxraPGwmDrJH6dpLoGJO
LyCaI1rZx5A4X6G4dCDpFGufgtwfnwJcTNNxu9l7TKy9HUC20IqqD4Uk0llgP7pa
aaYqGLKmqLojxU1d4TEs7iWlU37wm2tLlQZIYnJ+l0h+Vir9ntZd8TvpRhNJ+2WJ
ULZ/LSxj1+dpJbflgmAFlRPn+6cMqjhRRd/6fLpNmyBN72xx1Fa7N5LwjiSCASWs
Zs5OKVDvpO3sHB5ssdHP8SwBxksCBGKBXzcmgfgMP0n8QOsUgY7OJOfayC4AlU/Z
/4+J0YNsDz5q9lYwfqoD/fHjumPuj6AMmWkKhwnLgmN7rtLb2oUqOLd+3qIDPKjo
rhM2HRs17FhyxfyPWkuzgbc7u3mmYGpT8tL5xALm9NYX74ns7saSkH+UpmNgN7o/
xyu7uU8qaiMnhq5MpFwAXNOdjIjP60Ov2RFECpcNcOvXY4QTqRV4GzBszAqMCmj7
R9vTJ6O0ccIP5ldFOd2Huaqpzmzv5gaxXqgxJkvRb8QVJ0kn4CcTM7Pf25RKUYYK
bRHuj96oSjmM4nEsXKRzMwnTS+MPId8neE6O56OBtoW+vOs9t3F9QLFGswVTQBcq
9eAIDFGNw/qDoVw0kfpUZ5XJjrym2MxHDe4EdyVaSSxY7ZgmDeryXWL+Y/pn7wIY
SOF1zel1QWP+fYPf8CbFLmcko0m4pQwicne0sxb+x2tv8FdWpC68DspCOdvFI/tm
f/eTFgw7bGVj8+zaswnwg8nswBfo0narNTakRNFnkOnwG1tQfRQN8/vQjQwDNV4z
jd2EP7a+gILGRLWBT/7op9zIWsxL/tvsdB3rZ+4MD7nVxnObQiw5bTzy/wcW42Or
Rs26ayXB/MdMhgKB3xQVHtwA4eVyjBQfrUxqtXykHnGaw/LY/xxH2yOfxZzolsff
PPuPehx6WDtb7k8HlLbqDLn/W/KMw6Wqjjx3XuBgLW5iBEdrpZa+SyRXzhXeobAy
Oi2ZuVVMFphkQKWqPluHuz9qedUyT8sYsDC7HnA1vEDXskhs4ZzLJmO5Ep2bYicB
nqHEawAuFWO8ozhxYaTUyA3npCUQhxDHnSnYXoNsSa/1K05pA3gkuZMpTKYsk2tO
opSBMI7TQJNbMFNaiz1qmqqBMRX06UI3aEgWBufBLuH3ZORQuqez6tZmYbHdoI/e
n/rIF9mFtxqZzCQ62+infAlcVGlFS3WhLAXhVZYqQh66rJJQccZk0xZQy9rJivc1
xKx4+KH9Kf58lz1ULRSH7oTQNwi8+VHxTPmZ/aGd1PuJJvJgufF2EDjoxxMtd4+b
hFgbB75Lclug7txgfBR4OQjlOHap6lpyBWk9MKKQ6PiNsOYjlRTBYlFWbfpjYfwL
OXbR3lZ070DgpRiQ51rA5flU5WUsRXIu0+hdXZTvaMVxyBcMWvRIYbzFxxSHKP0X
oWeoQ2OgS00Ywr0iv4RoLDpKO4yfMKQo8l5TcqRwvthsKFOh4Sj6E1m4rk4Xv74e
mrcTdiH6WLmVXRXM0KKI3NPaHHZ+xrcjesXu9KDGeDGjwLqDZEfqcfslKbH5nguy
lCA6DmNIxv7XlKcvQBXT2ASimexpD4nWlJujHoehmloK4tr7dcWO5ElVm+MAs6M9
0nUoXGavc+XoP2iP34+zE8GXQcavMtd5081DVuKAV/NwYbNk9F6X2Q+I43KUZGBZ
bLaAR2Imqo7TTc5GAyv8vpM6rtWkVmBGdpYOQyt+PC8w1jrFdGOvI8QMJWM34507
A6EIc60DqL9rJsvQ0ug5Dlb6ve2Xh1xgF+7pxXIJ6lNkd0jwpYcWLL95t5pmUcKk
LOPhY3YZstzXilkpg/EMppl3gG6+W+/PLgEDqr5ejO4l2ltly0W4WPZLLlCXvfvi
j3SJ7sePzvFVKGw35cBnFyy6Wl6jZeU65o2as9BYGlv7wsFev+Dcm6aL2ZgAbafV
bnF/q3FiIrfNR0Z1xm9B30vIpCXP4BmR3ZywFnaigBtKOOHvKE5O7OYSXaqEG9k5
bWSgCkkqxJSQpkrFMJIPsaaBf0Cw/3jMp12Tnw20XmMLGUy8tbTgw57gnqOHrrUe
cIGc09nsvS6JgqYVsFfGn0l+j8Sa8Ca6f5Pft34U6KaGLnQrNFVO/Tv7rEBc4u5j
jjQ5CPHmFtA6A3WJ2q+fWmqAzXpulLeStOsMUmF8RZXZ9S0GZ4QlvNzXpmqOkXx0
h37c34wAF8Eh7jiTaygxChBl6eUUKIVpMirqAeUOw8BtIYklDxg9bbpd+Tyzz7EE
H+aDIDUjGur1IGyPtLhaLINO4nHToP+RcjHDWJCFHdNJd77FSRP5wN+PKvbMo6l2
6UD0dC8pmoqOvtiqFQ52UmtYB2poKQcwYLnBD+Fn0x0oYKvVxrJC86JQfTTfnogl
vZu5g3qETY7q42PZv7lhLjE+fCwg7zd0+H1nezF9UBRjZTqZj3pCuEG/myrCHJhp
cLjHgIiPEcUXe8sbvC0zSedteANhj/Mei5m87Fh/Hc2AjwjEcq9Z2TbJAx0Vt8g5
ZsWq+rDcyhe9o1jJpDj7+1uDjL1/ds/UWxeBbPTcUlWd6RXLb0hg286Yfs1esFKb
l+izRHHlAK5y9jWi/Ri1aEZBJodbcM689EgzmYowwbMc3wwqDZIqqcHRAESUbhXi
GV3Ef/qEtNMAgA3JEa4IFum9zyDsQrDwECnIXEtI/IBCfJ4MMrBAc3CO/YEu+TgQ
sSPIKyxo5vVhqKwhyoCtaj4a0I0ZTF8B0McVVwLrMH1RJnKMH0dFLvoW4WfluPLr
xTCZS69Ln/nJIeax62fg+D5N/sx6a5PjtMHA2JgYnHuPPiQDby0Qi2NyN+YQO3z6
jjp8X9O+lxx5DKMMC/MgauxxixpPc0WCw4RguDM9H+ymVHI6tvhhLys0xQ7mkOHN
XBoTZLGAxwc4PhahOOg+YGnJCpVDJJ4KZ+LKKPD6u2kLlJl1xJgswSG5bfIvUaUQ
nx2nExIdmlC19I3uzO9fHatLwK0i0BaKykqAaQeGAeM/QHYho8h2DF80S4/l7/uU
sR+olspd9zPyWTW04n4KWEqV4mr6igEXKX3xUyHf9hT2nz8YYhrc3/NYbCrUnHFs
bHeDDieMYlyeYZqPaWCFUsoG8X8LhvYt2iAdhiaD0xAf4FEf7+l9Qm96alEM0G7U
H8m9+lHywvax6zwLVJJxq0Gy9wWc2b+tMKgLKUo+iLUPxm/ACF3GRGwvS9axoCy9
IK45Y4I91urXuJ/b1XRFoxst1Lc9NS8PO1UUBgt/Difg3DHJujaByLR+rSHAb/LC
qLX2oIj5eFW6rYAyDMxGhaiJxnnHY/d52WLjyt4eaSwL2qpQfOqgKkS1YuPX5bkX
gzYzcaPTkvaMi8p+DkErIk5eKciu3lAhOAiEyJY9aCtEV5MvBhuKnizTHqk2K0fs
Jh2E1eOv8KBhd2m125wqXvt20RlNah1xXnI+kVUUPWfPXpRVVQb8Sok4VMqAfIIW
dnLh0YLf86ILeMViS6C5KKEqcC169hxdZ2wjKjLQz1CWXOY6wALCLO/wg0AkpRDc
vdx//OFYFDPJeAnQdpTtQp0eWfawk05opoZivCpOglM1x3/XZE9L9uAiLekIR/1O
6JxBkwY2w4tJ9aro2035DJaZZeys8DY4afGELB7o5CrP1XbG36Zh2PFkvyzpk2Rn
pZBfIm7MVeCtxmdTEzp9Lz9dUrD1e2z3zH1ETlZjt32uK0l/dHxaXUA2Fv2prWqC
XJlIIDh5w6OeizmQkyQF/V7K84cdkYwYJEXfMWuZ7ICq0fdqSHFQ1TU4hUazeBHI
nTafwmlhpEh2pQkTzn7qr4JzUk07C39T3vaSvfJNpeA/P//9dksu7Om7eSmvH6rI
8iQ3YXLgwNuTKJhVKIL21AGiSmgO0o1SLKbqtGoASH2De+fGpI9eDC09h1AWASiK
/E+EvOi0jPsrDOrInQ2dKObhueGyjJExemqtsX+wWe5K2S5+0ptV59Hmw4prEMGk
ePm4Ovb+HvWiygS9uKaVzLAQscLCjEe6BVGz5Mtjh9fyKSap/eyDgCO7i8VPyag6
+hPY3wtQTOz6ovueI13nk8UjaekqwEobSxHORSyovaXyZCIOyU/3PdBOts1exKkj
iPPupSC8nvp8dGUfAgGsHRRAIaF67r1SPMnbpag+E50bSxO/FrcdfcUWMMUQWWqP
miV86uFwzhMBEn48nnwgJYfZjBdSkymxTUx6saZzCXlgcWE03crp7b+LLsxHpHFf
7YDW1bTxTvxdqcSCuvipf4ShW47BVUQQ5tm7zcjgojymU0cGSb5OBU2wGQcMqgOz
5f+jk9T3fHbK4dRBzVmumnyfyOKfpsl8Qfp2oeBU4Oi0/YpqXPxQDgrvcc1+pviG
93fvrc5g2bK2AMUJ2fLWbq4tiV6wltBFf1h99c65x/IRL5cqaA0jJOu4BpINBd0h
E/OEWzzKZdtPHLgn8x8rGLfYOZdV36u3be8kFAnyZBUNPbnET5fgX33vyQsMH8Pf
hNIr08J8kOPJPcrCHMgC6joB25yL35RmFeEdUeSbZopfxw+qdoQmfsnJ0un3o/7t
7+dByHb+5/2k5mp0pSCmbKG6IC+ATZxRx6prFzKe1iqE5BrUXbDqbiWwHTW2GhCt
M3jo1j+d5fSSm5TD1z3fu9GgX3uajX24QTgPJDiZRryU5lup05ki0D74rm8wNtHj
pA6R6iamcYftEDJgKbnkAlszyc7qV75uA1Kca+Run1rCpIvm9FQad+TUn0545bsB
7EWWlScKzCzOPGzOvd90cq+g3EPhNmOU6K2e2pvz2iF247eLUCc5vG6mh9PglGEY
sF9ugyHKPniIWGV7eLkjYkz6O9tZxfYRR8yspjUei2uHhiqemtgaj8mhtRwfEhQ4
09tLgvbRNl2jKKhrwomAH1JqgtbGm7u/wpmNlOJNVSQ4M0o0TPZ9WXL5hdlsUZNV
W8yNRBU9K2hTnpKhNlRmm77clWdsRBeN2g7PzEkZXqTX/l2yDhlhZqwkkGSe3eXV
KGka5cQufZqtQ1ZEGo4m0gYToVsrVDwvpuVNYnI35FoKwukN/yOAOt5YEDL1Buv1
49ABi8cRv/YFTnc5Exfs95KNuUQOL4DxyaP8w7cblJr0DxIwkgZ7oq+PQ5G1J8aX
0rTJksbtdnm6OND6MAeJ2Mz9xYQNVuSow7jbrC/x94QlhGg0EwbmmtGuB/nfzv0G
FYc2SkDFY4DYm72KwCdlDyR/kxalzFfwZKRhrHNfld7CToRHVmV3j0d+y0WJD5AJ
oqZFTUm82S0/uhEYrz7c8p6rafVG1h4n9El7MNm3dNnuzzK/fZ+MKEQFJWtSb1BI
rRw+cfTerhxZkA4ozlmdgaQkwdw4DgTOCuGgsC/YYPQvB/4YLHU6ot+ww7wZdLBq
v99Fd0nEZb+rcSm7P7WJLvDmSUMNsw4CnPm/S6xeFfXaKao0sEfC3XQbuZZ4zGz2
UlsT55Dd/9gOol6+bfJNLam501esVGwv37tX/W5Ww4tu4YLGzYqmbJvKg3FNLJoU
NEtrVx2X3q2dgEAOngXlc1ES1l7FqQt8HL8QybAzqhpWzUe1jpw4bW/yDkD20hgg
j8wVQUoFq9mGp7pNuYKJFUvTF6FycUqzi9HhxYNBQYY/J/jiLEDC/GQ8XFp4VAwp
2Z0CY/xA7uNbO1xMBPaY/fSNQDHLrHic+RyVp/ZyxRGp+hZn6VJ3DP/DmLolAd9c
7nsZkiHbWzu7oDnQBx2ZKfAwSIXAV7xn5aoj2RQp9gzRduokhCHPoCq2acfjYsqq
yhm+MB7H3rlG3vE8+M3pJqRJY5eGS20yWMNGVPuZzVwyqqVUUNJOrp+kBvicveH+
0SfXMAscDJp36nbjgXCSBSaK0GtgfkNVOim6wAFNlZk75ala1Tvz/6jbWFk34gtj
DdkxKbBiCWJ/0eW2/YZItLuosLpzLtJO3V/jTzL4lZeprQSNBpIzOr9C9bz/GAR7
0fqNv9eQmW2iEHonF7elbtmCY7uNPBal0Myx1IKc4Q3YOYdbhw+HTo0uyp/f4F1/
Sru2awOiWbRbGFiU1cTuAzeIfS1tLACRDKWK9iCw+L9WPKsUDS6qBqKC2HTyyIhk
fZe5dlj/xPF3Yf7wtZ/7WjH+nK3g9f9N0JzXZwNLqEhlVn5tMdZ7IgvW2KamimHZ
KtZ/GwM0JfhpyOzKYUAh0nGYJ6be6TrTYsyJSbKBvSqxyYytOTZS87i5Bn6FymJG
vS9RTMZU6uZL4NjgY9i1wKbwD5GCWHmrqYVFeSMBu/1CrXb8QiPf7Z06wenpaGLU
OI0SwMPjIiJI1W++6DmkaXGFd+QRsYmzCeA3b5i866Bj0smtdna37UowST3zqhox
fngQzoaMM8E6wnejjGwNv82ymVFpPCAl3/m32DYeGke88jRmH84bSyL/1/urehto
8BbEEIYjeooVLubl1odNxjKte4TrViGTu2189ff+Gj3iXgf5cqd2+/zhzaSh7NU4
DazAV8OWeJkvnfOASCoo0ST2vi8UA/wJReJ8VmdLrpmKvHDXN0y4L8x6ce3ULN3P
k5DgKQcdaLJk9ypyDP2f+8U/Q8OEIdn58OogHWyBoK3VmBx/kiczqxvgD7pktUkw
W1FCK5pr3B+m/EmHEfxLYbwRklyDwbTvnw/7F1ARX143fStK5DReqMOQ/E6392mN
pnjaAZUscdX69riLgpL6QcF1ZlC9Rbv3gq/qplW7k/LJQUHvFKrkUvBsPFFFP/PS
Ji7NJBMVQIrDEeuYFz3tMG5MxNUIM6e2pOJo9n128hfBetPuQm2YFTiTxg+5DcKc
wnck0zNxzcC7BITIfCHKWS0CmQiP4ZY8fA83M8QFDFFNNW/Ec18a6nA1BfF2HAIi
QNJ6kAKV1Gj0hE3fEfUJ2Oa26HajSSwkbLr3+WQ6JHdliFiXrZokcFY65QdSRrH3
b35xonMZ9TJnIkWNOhRPq85z+OHYgx3qE/+PVXMlnadkKNu4+qFQ5IWwRBHmhlJa
qIIkuGXiuRdjcbw65gTBVmSqnshyQybwyeLRSQ97yC3ZxjIfy7Rtuw6Ovc1N/HJa
FgF1G5TlI3SlVzGGz8OXepHfc8Ei0gZqaILeufOQhB4ZMe+/xCZn2n8saV0bjjIM
pnqaWVf87Tvmqsxu1/n2jqd389cBPwyIcFixYWrxoi8W92DGaKVE7qbC8lTslfz8
8ReNop4YTEp4PmK4NK20S8SEKS31XlIhX9d8Qm881xQmY197yln/TOgoz5Qtchm6
lyYRH2A3EO8je96zy91EZPhZ0s4yWFa5EYoExMgMTCC4HXFtGqi/pH3ng+kswnrc
4WKrzhr0qjgx/yS8udE7T51SJ/eaDcE9b+3WCtEUuGezwbhoPzXGlD9IFAyo/srx
2O1atxgzcO9Sk6rypYQ1qdTGD8lpxdhkT/ySmksQagtYUjbfqwqActnRCpAQtTCZ
96JEgS3ltnSQ1EoLP2grprE5JrXXjDoE8GLS5/hJVphtUr04VeBR780mrDfh1Mmn
6fvbzxTClLZcOSZKNkj+HYl4rg4vdc4mfw4LIKld5Cyc/egcUeHOSXBd3sDoBYR3
6RqXl7ObkjSkhLTOk5OzUcaLyw62Ak9dB3sraN/2R+25iIbsleLn+me6e4e7B5Yf
oM3KSO+KG8IESr0sbfhyUZImxRN1Asb66PRa7BJ5b5GVqZB0sQSq7iNcrSuchrFq
/gtLgA21+F7Jy84Sk0Rcujod/19PmuVz+fT/zp9lzu9It+Y689HwDSNc5LIc3K8P
rAYBmoFHm2kn8tTXWLegx8wT/WQ95+GFZmKV1LImmCz/QAQLtlKI3sf4ttkxYexC
kfsETqELQnoiiDGR6+uTYKPqFmHEilXWjOreLbz8f4Zk5O44guM5yGGB2TTWkonp
NavjoQxS7fv8H1EfA+o59My91EzlJu60wTkDCKY/TTdaPrj++0zSvBuL2vsFpkr+
7LAiw90oF7NyXP/ETIDP/jgDipobEuLua7WNoB9jqIG/pFtoXy8ctcMlkXr+bqEA
3pmpLRcz/5wym4zmB9SckzmPqMkkriz1+L4ob6dMjFJnlrjJoYmZwIRNEOUEAsu2
+pXOymyfS7O+tixw829vUTtccj+/4R/RSGI/wZ51pFmX1FXmI2kVJOt6p1dAqq6M
xV6lm8eBKCkORHAwhY1NEvtmdtmjDK7KF/kQhLzR5eqGjSEv1YYEkp8+oOdex+SY
PVgfZM5iDnMqOO06DWQdJa8aREOsowixfNgXisU2oRVcEupcOaXXF8FCONbxhwI2
wzKqrj8hYe9A+r6cxcTXrNJhtlPVuzfBFoxryp5Sdf7NyoTqxAJFbcxCXXETxv+9
cEkymM2K80lNEMoN7jdrfC/egmL/JV6yiQXpjyEgx7xOpOK75gKRW/tnSzN/JxI5
Qtu7wEkpKlDeG+HiGP6ouTFztiPi9DTOlwocLKUYMaWrLwYLXJC+YyI+peYpY/Vb
mHDsTq2564X1GblxLwvAer/l3Tvbu97L5OiHwuRGEeZTMJM59orbtjbYhEP6W0Wn
Egac22M8LwljzLSfnslGX8d8ekBx7kqAz/y2w0/El4dl6chd7E6S2PGFvl1G/dsU
PkT3JOI5ScJbMEHFkRUAHeBevUxy17RUAnDc0FXvnTeNtLzBU9NWsTxAg561VgoZ
A4OTDIbclYHY0xPut5Nvk7eebJVCKlmMARKLNC0EetFWHInY9oQfaWTxcBHlrDd/
q1KfWraqAlYmKcY80X3L0bVR/QdPM1IHgdGom3JIox7rPYyY38NQMSIaJZ6M0G+C
NfrL1GixsHEZk7epPEX2+MBPeWKnnx5fUB5qeh6wawN8zF3o2KpQz5XSGCVpfjpB
PIFjyfcXd4In0niwBTtLinPeUydmMZcg6TG+6FYlR7v1K+pcmzZef1AAOnzWwGO/
aYsY/CZN8xZfFwswNhn7BSgCX29Q/s3NsSptACUSc/SKyfepjedWxQE8wcNiujIl
y+X93A/gRVhO4OjXsYLYtcTU+EuxI3XESbo2IzkqzASyG4GrXJ6ZySBRn//6SU7j
FVswqw8NVcwLbngq/VGUFa66eDCtPZYHKJbpLxKe1XahMph19eNjGIWaorYc9Tb5
IMs+ogwMF42qv5g8ouAdgSgfWFARvx4e4tteBoO5BbN3Vpw85mhKlzh9x0ayPPVu
tMpsf6Z52JdokGM29+azF7m2C/E1JvoioKhrg3IeWJbWETig7pXfDWOVLeXKERHk
0k2T1YPPs7xwcIX0F+83XeegGSKxz/x0lcKdg0SE2UJiMIfAu8tlagyXoDM89nPP
A72ejNkQo2k3jH+f4M1p0FFtxq8ecKZOLIjh+Wv8mBaG0F1AvYgYmSrDemfzW9CG
YtjkCZ+AggxeDHELhg9HPRf0QPAtMWLrx2ZUTWB1n09aq6HH1iy/JAxEfXQdbezb
3WUy1tQlmduiMcoFQo6yADSQ0h7CN15ynvQCtNeksPkmP5EfzIsyscK3OXXoqB9F
38uAfju8mJxDWQho6Vf/Kk2t/4VC8QCaSURpSKhXOl2BbBLRsw09PHoiatJCPDyN
MKcTSXY9qvQhjVumRmr7f23ccyhUX6mejwdTTwWd8JuJ6QcL2Sw1fFcKVjxa8U/y
/in/FwJb6ow0O2206yez1BCvhpgplZDa4n/J0KhOH1W4Y13gxVUJPw6fpcLFMJjV
Utqw9IL2Sl1OndBENYEXY3QPIPiNZMkFJNapar4V7ptsASpJof4+fnMoRLiQM7M9
6OIVA7eqkLMfy3b3rk6t4SemmJd6vLKL6YuuVvxO5bPTgHHolYsINEsaiGxofMwR
+8Zgy+SzPwrkFqZQUswqfNzWD3AMf6T9LlIYWE5/s/dzbFnqWEHdoWHL+YDshgKi
M79eifcpZT9Td+B9r6Lqj3jP/RaLdX3hIEH+hHegKv5Fly85uP8oi3br0keZp0p+
yn6tv7HIiJjYuk3mlmlNOlmsAqFgNXh8NsirtJU4FXSY+oRcSToyr7Bh5s4mCdAX
3ulYKFEVwfyL6GiNfhrfB2BGPqQmrCamkKOQpxpjZOyoX5x2/dsGGOq43fR+BPmj
PQLMa0P1q2MaA+pA6bHyej6VsGaKEFeZkVUm1D4+PtwGhgCwfsvKm6oRUo74zzPN
V3Yh1F4GZGAyvDerIoLlWvqqcGzBivASQxdMvGqdrWegHIXxFCb5y4Xw470EUGYf
Z0xgOt8kBRu4zGFSloKS7hBLDAyCzzy69lR1OE/YNneCgyDSwk5qKmp6InJQH/86
K08NdSqME6iQoCKC9Pw/oM2CrirIXRQc/VcVOYUjbf5Z3tSr6n8JIf/MbRQwiXqS
8xDwORoNHQSLVrOPJ05EBSdoUvT/LnGF67cbpC33KIgkwpzWM8F9ek+s7h1USLg8
fmKw/tQDd6fDvrssH8Bfq3mTwVNQe2fTxHRTQJExwaz1SaaK3wEAMCWq9NNgYUv1
TOsPGkmjAjbRlGHOjRkljwidL1hR6WJkt4Sa2gPHYunGQ+RE/FimOwVF84GBVUaZ
5DsgRiy7S8zKxTpscAk6gCU6+6aEvDuEP0dmvaCjtu+3rzSKQ6z7b3pGRFDwWjBq
zx452DotkXJhOFdQx4Xlq8r0kClG6fCtZqh6iBaLUtJO0VQ+lb38b5Ukx0InoSVT
EqtmKBRLse4oYahzvxbhTB/blMQH3/BOL6EbTtwf6B8yDYL4sH3MT5IpVFbwzSJY
f0GjuHmbdOBZvyHvxB/8Quy+R0uw1QOxwIoFJEytg2k9NjGRHNB+J4iGIHRJVSyV
pbX0mzk3KLeazl0rh5JLGkuBdhJXHc484fduxgCLzUHVLqYpTHvhSfvQe0ciA9Vu
H3mBTPpZLI83uXOVKHoEMGAoERKZLiRjoGreYTvl1YzOa3U9lj0gK5kOtBdS/R4r
iljQ36MeewE9uInpm26I0AujmTvwS0yt2glSNy4nZkx38F2jpYY2xE+IF3kX6vQz
0EgvAyL7mzpL1CGRGxLo86Hj/V/jNmbUqyCjYvUo/x3Ngr+8rFr+Owu3FPPF3/mu
JRFA7zPwx6glxqwcTby3hlVuBcHOvVJZHUasUkrYBtL+7NCMQvqC00NCZxEfj1RV
xFjqja0S7uGKgPuCwOJGnTcqD3dItLsPtdHGj9V5MmKPo5UFRvWdRxPqNIFJ9Fh9
XFncuGmEULBC/LMoOsh2v3XFFlF12fyZp6sQXXA5LyqI3h2vEnGxrefany5kdF/2
4BwwGLNekuEnlRI7cjAjgEsDXKpH5SpWQm+rdlmx+XnnyHEN+gpyi4xJdf+/ry+R
82+UN/9K6K2wttIkJE+DSHLzzr+RSXj4tiZBjAl5PwP1IGRIfBzuEAkNGUhpFOOe
74nwQGQ0I4K2nPxkCms5ax7TB0KGkFexMF0DSxyKzacjZuerw7833JaLW1wRTIRk
SPiKppqvPXIxJqBHzZiIOvWp8kZy2tpki9p0uMhoLeZRDHqZfkdefapt/ln/iHrn
H+V6DhQyFHAH4XPcCjkGgRwhVA90m2vAupqJZMFDQgWxJYgXK7fCuDsovwBk+mWG
zE5B0reLanUSnlQrflKjhJM91aVWHwK0jTDFDD5cEBC2T9IOdu0pErFV3r8kVuPt
LgZsACabc7PwF4Q1aNAY+d8zQi2saWgy3ACxHWF0auGGWb6z2Jo+ecUfg8fCB8jJ
mmzjgxEjH22nbSHUeUllQgXGwcp49vaxSYpH9EsWCtFrL7FZ/hpTIWVdIKUaA1cQ
0DVM6kFwc0FHJ2+6WWEtRVH4Ij/+0pj5MRLrUHGuofIxX+dZf5GE5rRHsaksUV5e
kIx7Ws98miATGZXXAUKvuNHX7f0fa0GH0Go0gLmemNKz4fra3zHkvPlahIFiThZx
8asClMqNNkxyiAyRDXbyZ1+dcmc6eoEjpAjV4kNyQ7H1YSmEp8xXyH75x14XQZAT
ho5xFHeaJ1jHa+bTb0njXUEBffUFqPthWL9xs1dWzdoZIUjWuVRjW3ahm59M/ZFX
2F+zv/fhdWwUTtZMM6m7ZRR850htKCNq1rZkBwLwFloQEWXF6PbJK+uM9fZyfNM9
ghcKMiLn6uX47B9sjqDpCgoAWJUQn6FlcvVr9D+7GA6uy9OXPP4Mr4Nm6EOQ2KOW
DtAUBmvvHx7W9lN4Xb6d2VuzIKnZK9U91+0HVqL7rg3kz03fQ5HL86FemXEKXJQ8
YrJ4Y4wUAEeM2mfPNOyve7oD0kuE9XpXeK0NQJD/K8iBK1R/nB3WZLzvdSj6fvDH
YBzgMqNcD4GCmobdIeZf0veiyJNpvlwb93oZQ/CYVr+Y+uAoY9/hM+MhW7gPsXFU
2matrHsqfhgiKq70Uvq/4RqY8QwB8VyDJfhyv7hHlw6CWPBFiWCA2jQPEKChrq81
nIaDTcqX2LzqIF4Fxq60jSZwEd3hG9XHp8HXI1PZQZB4q4JW/GMq8edDGTfQSiu5
zKMSZs06BcNs/v+77B2Bghu+VJDonswy/0uEj31h/qPYDFFW7i56IGp29SHelQjM
c14G+tBk/oPcDoODbGHIrpKEsxjipNGChffzUbjYJz30fZ2fW8XEC+Ht1L8zd5y/
dP42LhL2fVZ9sNomKlyqAIBCefOLCi8SdIltin64OmLP4coxehbJQCg562b8CnV7
j2WEecblK66I5KsI/TcABmWGatgH5WwQGfXRYzsutX8VK7q1Ns4S0zxaLcd9NDqp
nm4SUvMRX3vnpxZGeJmb8J201ZKsKiRohnEUb236avWjmjadrktDc8I72EuXNNFH
iJuTgAg3Clg9LbCO2wRj/nPvkhf6J3xWMvqL4yzpZd370oSpySOSwwZb6Rrw6XNn
hLL6O1yxfcNlec9EQy+6xQKqo5Gbg8MacS+qzFEL2TVPNenUpb2I74VhTIBM27Co
iqSlFH7W6GjLX3zYFMzaGbLvBzgc8KYJplVk3AlNJTvl6MsOAy35Oum16vrspBEW
s5NFHIXUqR1Nnb+t9ZncxMtehOnPVdiTGCJYGsZvq5PvJnD0baoIPyiKsdafF0O5
2nM9DTJGRrBpaWcjg/vUgExY4mGRpaVHx6HqBO67cFf09seZmuF4IOAccDYClRPR
o4YPzh2dXVaZyA+JMjso6m/xWn67zZv+L0RZofa/LG4JGmcq0297tH9W8vN2DUpn
MCkazpU8G3ebg1Q9Qh2IuXPxX8U7DWwcax8VE0DELc0aI+5ek+1GXISdiiUwULWF
JOYVvOL0Bok4czzYW8pgJe6oQB/TIc0Vk6Ra6sXGdzRAUf4yMEOBFOhg+Uj4e2/t
0juYajBnM8egpPWlPjPcfKbKxb053ueMHIV0SKBxf9UyCjs30S3OVqe1xRmcdyER
RdIaOp2g6BSPxojmYJxRimnGAvGY0yXiaecgq5QgyhY+YfO5Z5MgGjlWZk2jZVUB
ViDImhnHS3c5BcZrfhEjF7fJRKvSsL4fh8B1t63ajRVX92YIC2/ILbC5sZ7BCelL
guf3PJKIuLq12+SyoqT8cgHbFnYwzrpFBUh9TZrKADBhEjHuQEUouTQ+nODW1r5U
N8qoAVqWr3hPUYhAzbHwhEPkM4lltKjaCRp7Q4IdPJ3QqZa1CzH6EsuEVsLP9be+
Z0ItmJHXLPJNlmKavOhP/joPcN4QCDA/HcBWriG6Rhz6XjKWfh4B82f94/wjm7UQ
IeJZ3JGKizI8+cXtf8N3J9VDkPHSVGKRhqJMklahvAnRuP0xv6PUp/qr4fl0gqDY
Cw4gaQ5nhRWgPSGTXCX1bfUGPJX+I2MkqzFwJ1aaKjGCUD6OZ4Sjm8iqzMJ9+f8q
6MHXijN4gHu5nvftjdZiI5Jq0n6J6s67Z63Ib4L+TzY+/c4EOhbA0k8uDcZZtSnC
Q/NF/UiNRs3TbZPpiqazSSJ3z1V8QdFt0XnzkLIRKJSRnIAXFz+k5tsQo002oIAi
XKSibnOKwLoo2k3Wt7AbyNzfQVaWUuae+BdfcVsWQqlCJ1ZH2LddRWVG+LY0rDsj
D08oIMAiznJWPd6CNqpOfgfxQnf73+l+qVwtfvlN6RogQZDyJYVsQN6ZTwvnNWJN
lym027mf/AmpcrWuvfFyNOqyaICUIiZJgtycbhw+SzV10Mpht/4RFBZgT4EW4owa
QRtEAWhwGfzhmifwIndWFNMf6S2wcSySmHxDbKSGqUAVXVMcB7YUsLq1eRZFhyk9
FCW70EsxrSHfgYr4wJoIR/sW4R5t2x3rMwTcISfRrTiaVIyN9jGIrRj/Ak1bohHQ
2qwTPwOb3ZDudt4XpKNkdr/qNDtoTR27S0Izkxk2obSR5VGoXaABO559iCKVCfCg
xSNXXBcdt4aqydE5610l32hE6PxPXIqL+3XCAVE0tKKVfCYYmahgRgpx10MXdoF2
+LB0XcSn5oFzJLuXhG9MNpyz4ZV6FaXRLyf24SvNusnayqtGSAm1bYkRWbNRSjfq
5YkoED4EHZhM5Ki0uiBUp8ZTnjoqXV+6Dp/EOViJ6d7dP6X/oihscQD13XzJiLBT
H9fhc7/5U4nkeMSsySIGvPUBl4EUjyhlHO+VG3183W9VcA7xc5wDC3XoflUAR3P2
rzvXF0SixyB/xS92ji7/IWDWBTE67nB0UxOGXYwiAHvcGzV0RppVShxfnmUz3qnS
jrJPmV/UyQfV/qS+eovJuFyXpHt9AH2HladN8MzTw1FRAu27DLAHUkn42+e8YdjX
TJoevbuIwKP8eGvTLOqpaU1zbJqm6vfDeBmJ6zgTBWJ6QhQu1MWm+Qm82EA5rDqU
ExEi+E0aCYq3jHJUHYLD7JDroMCV8foO6lDL77plKKPYIItKQ+OanMPwAo3nwf2l
YeBMax9Or0R+62zwYE9v42G8l970d4IB6jGVsMVoGIYWr9NHByNQF8iCRIhS8HNr
BYFv4JfyhyoSp2yX7qwVXq5XJuNHWftBLFGcISv/wMZrQwF101fi33d1D9ZeVJMA
MwTeM74oVc/Kh8Wbu3hb7iI36y7GhpKdsisLP2ALPU6jaZIAgA/JSdnALmdV8VbI
z8bOT3YHihSNR9Pg2h/EXQks+3FMvAANmqoy8lfypmKf3MDzHPf6O1Y6fWxonJo+
v+k8EYk5IMySZQONLKW8lehZKAbxNxWuWiCDVvclfSgikrPAQyZ3sh1Pb13DkQaq
IU5kBrq/7ZrjquztDf0IVyp4RXQMlcWFlf8XasDmK1SkFcW9SIJsEnCybWa2zXLl
uClxgxtauqx3d1MnRv4IW3nqDuuOC3+KhaHCVKZUy3kTFa7CyQgjgAgSipRt9n0/
ipg0uqkgGsLJXr2LOiilfRXncsUntk6J/DxdcKtbMGVJG6jwCUSJDupqZ7H7LKbk
Kvdyf1ieQUvWFRWHXBFiWvdJQMASzEWXG4+QOymNeeJR2hsFYLLUDvkKeoYGhc+c
Irx2wStrqOZWj3bhpV23c7gh6YwTX4Kz6wTZ9XzjY+x9NEaN+D/jfgZTZrOmQSnE
fg1rf24nJIC8NlghPsNjUmG8dT70IvG929QyU1DlP4Rw/hZMtXkUh/wmYFeVyWdY
qajiz2+MxSrl8FLU5GL+lanmbT8yCLW0BYFjw3fL98V9R6QO1RVVdyLrczQ8/JUr
x8eAzK+zPkwdvZ1MknJFyWS7IXiEUOHsedJtSTpPCt7YHd23NS9xub2O+SFDii68
SU/rm41tFVaQ6ASLiw58acgqMk/AyVRoGHzWWWzsQb6fh7UpU6GlwZkUyLtrjURy
4HZlVlbN0FQ9bWeeL5+n+edd3/25C6QXLZX+dO1b6EChBKIZEhZZYOMjbSZIs97K
scdbC91W4D13owUrtVmgcd4Q706qDuDfSQt1vYkbxNxMx9c26UazFItUBcXsJ6Ys
pnhTW+ENICBaldzrCxcEQ9KTzpsz9S5uvgyoIqgkTuN0KBo5nb6jkAtd5nL4cP83
WgNJXXz5wLSSIduORyGNi5sXvCEXr8RuWamjY+Hw3DQ2C61CHDpKVm9/rIogJVLW
fD6ASqpIkXbAGGDbicdXpIV23GAnzABGAjVpUGA2ZmgReHoZscZO++NozXuAwGra
pQj/KZ7A6toNxjcz5u9MSS2KHJ7OzicevfrtTeAdf7ZDjMl7akYujHX2jepQVDmf
jzD6/3u+IJ9jozyWfZORUGXRCKXQVeobnVjS29IspPvckUvwme09xF/M+n0e7f1J
w0eotjOsae4rh5tRmf6wOa3kyVeX57gchoA3/oxsYrqZtTBGUuqSlkr5BjxWYEYz
T6uyVPNwY8nFuSLyLfq4ZqtbsTLCNb3UaI9uPqcmsITDXHnSSWqbn4X7rHnxKsrp
nCQuNbPJ4ns8Q7tdBjCPK6DLaeKl6A68OVukfzn2ndiZdkEUSCev5BhM2HtQIpnT
u/QMk8f9QDqUNcRp2yKcgnFkGesVL6qhTrlUJYwU7JseMY/SJkm62yYRoXH2PGRo
V3T3DLURx2RfFfd4gOBLRdyH0sIzgxvrMykF+WKEoVbj8ZrZn+ibBa9hkoDc12cB
H2lA7u3JgGpv8wcd4VB95TIeQ408N6Fc27wPDfMsdy0TORdNuQERVKXDVpifUNk/
2isjvL4jtsZRk1aAzvbnhHIzbuclBiFJ4UihGTkG2Tp0klesaw7qNQmS3Vg8qWQR
s5GLojHaOA31+WqfgjbJpYHCfBiwWyXH6jial+R0vgaWi7OzNPjSVwid/5Tl2deB
T0N+MDmxP2hXpytDo5SzhX+4DQ/sreTcgY001IGgtv32ne4W1FMMG14mfDlv4Khm
qZ4XUpkshCkj3nZsplK9ij79r1Atfg//K9hh8CXOAHKlKAyT1Tj6+T10qKiskz3y
fkhDCWeRbzxdOAlYoMFXM//dTmhLE+15rLfR3sbmGHwD6IO5etnMoAyj7UjHCxlQ
ahk17apvViRCLTtxlD8Po3+VEFEIc8QYeT7ekVGqsfmdG9BYrjH0TIVpb+74nKbj
OuTEJ0tr6OhQgE0bq1H57GkJxvDX2ro2snG7CfVBsf37mpcS15shfxUTgXiKB6NO
eRD4+ArwD2E2cvG2sQ7X+0db+gsem46M+NfMswcWJSDtj2clVmpNo3I1WIIcX32J
QdeoMPS7+NRUtm+p15Q3NhW2QR/tlDt83rVr3wt5adZGvfZXB8gt1s98vQB1bT85
k6rq5WViV7zazgMWmWDWY5dc2KTEV2jePnYamz/GFvBxucHMCMJC8fJ4EXx7qL33
JYg+XftSJrBZchBPCEgU6Z9a7iPWHym74+KV+ooybgigCerJOKF3t876ijcDKgAJ
gfC1WcwXiIy7XGLF2zqQiCJiin/AR67/FvU2c7hb2xhVKkcrd/8woWc02PI9Jvt3
GbCXObjftC954nKGCOy1Q/lcakO7a4FkkCfIV6P5f1oyLlVNlfkJFzImp1953v7r
vIapdv1U9XnT+VngFmkjtvI4PDnYRNrmwNzyhL0+Hr+hAJsTB6MTbExd8CoIQAp/
0J8FnpcHhUDCBiyAYRA5bSk0i9h3IEQZQOlKGBQibKerPK76hqfV8LPPJMduKbZt
utI7kU4vpW5+q+zosji0JME3XdpkFs37fpMEgDhWiXjI3HOgvcxOGN6DJxCn2Ez3
0IFZ4Ydwd7snu7ouzup231dFwACWaEo+Ynkcv0/UppV1qmrNPe0oj5ZlgJhJpkPr
v7pB2OYAPCcnx43A1fad7LyALmypxBKp7Nyk0ITLuZnpm+C/mAKC/1KJOsZToqct
/CYc0z+otw6jdMIP8ESFYF0ZZcBWamWPj7XIR8XQPjVdDnboztO4IDxIZL4H8BCx
7ARn4EFmbkec37pGxV2XMtPLIhS7cgMnncn9NngcBEW5TCfYGCyavqB/IFFDWiaq
CXMM47bhKmQNWMhT/W0tCLklh1M93RRHpRJ7OYDgygg+DoYzjJp4pKaodszlS49R
Vy2qpvo9onQKT+pv0x95UmxoIylHJJt9FwYP0oad9x9Hvtq5G30Lxyp5f+V5l1ED
qOAx5pZHPe6i5cWaK5saJTeK82E4hAeS2iXGhRlUqaW170aRWOjGjTTAhyEPFTtV
yFSq7Wsubn0WiFfPIOPFTsXC7P7BwQZBJOQb72Tu+WddUSKX0lbrSgNLf2TaYkiP
07W6TWKO5xpPv75gHkrF+LT+Ljm6U5pU7HNHEzkN+AD49/Z/HkcEEb+PO46SeonU
qTcjVCKMxKjUdeJEcghUohVowp6a5MU4WGRK7keDiajT5e3RWd1DAcf2yQNjLZzC
eaogGOr10eTyP07r2HWkJjffnnpKwWGZ1oLWQb8DlPPl7PRXj5dReax+DYfKv8c4
lz8ChMvy5je+Z5x9O6N3hsvblSl/kgFqQG2luUuujXiRbYBsJ9vio8/LIgM9umst
FbgRIukqLN7c3UNOpnhvNS51tDOIXhA9S9PWgf91G7WzicFJDgD1ULmEYfQGQfxo
nNYII1K671MesiHh0vIUXEk1llGvTiz1oNLwnvQ7XmTrrUtX+2SlEmDASlPZPm9Z
erOwPTyDBmP2iE/rqCGxYlGBH1Wvbj7ZfwRO7/m3eIuHUuWMgggkVqYoVC0nBUFz
NPQBDHrP9jeMTG8ZJnxRlVPVB5QlktidR1lUoWs6P0jwFpnZMN+QpZbXf21WHore
ji60CkphpkNMBx7LY18PdWypu5sWPu/Xz+6C/KwI6qOEH909sLNkgy8YlG33DfR7
OaTZqZ+FV/jQQlxTYEmkfs4nwVRfAlP1OO0m4FHsNbHM6XXSAQqQTuCCzTCTroHF
L0v0E4u7MnAhL8K64T7mFTMZlYYhYnWG4wU+kRxLF9H0DbGX0MUgtY0s7aKuqJkb
Ym6KpPOtjVauNvyndIUtWx8kXtp2hGcYq/x8wGiy1s5A9NO7HzA22mBveRyJyyhm
p61zQ6LrV3ajrwzOIO6YFUDB2H5YMylOuFt/ul5zYhLRQaJIesUWa+SHFiMz8R9y
7kGAdvtNbaA6QSh23rh39cbeqPmWrMhC01dnK30ojxAEKlpLjgX8Pej0lnNGqFbT
j3kLGb3ztQiGp2N+dh9ANM4EqHVA2vkTU9ViqJs7n0ypfCtzCrYcDnN9GX/XDV76
2PunxJxDCA0YeANIsZsUm8PKIoty6TKOfHuFQCJwX5EEHncRVmrQ4biKiv+koklc
18Tu6xLRsHCKTdfWeSmZR1eXs3wiXA/IZ/PX1gQyufRgwCJ9vd14ry456MA3sgV2
6JrLDE6thFuxqpLdHK/QSmbr++hTKWDwtLqMXi0O5p/NdzYW9cFfdQiFtj7KZEaG
pNRUSFKBNh62YqgfkFxIHggg/JA4dVkAJydA5szRmhzJ81WqH9bdePZPfAuKHOuT
WhfPrd6v0XjGxmu1IJIgYwlwV506F9UTMUSM/zRMImWAot8VqiKeb4p3L5A8qXfX
oZQ/Az3Cn1NCJKLWmKPLwxdhiueZgR6RLi1GCwffIvaXAmaY2PAkuZHw2RpP5RyQ
SCGR487vx/TWD9nca1+KHtUC2E8CjddPA6fS45nlzX3aJsJ/WMAProqMgq1OByiu
FDCmxAjTKZefbivFet1+WkKV/0T/fLlE1nupoB79TqFZZZw1NRnxHShqIT6oqODG
zxYW63A7n6ZOHgV0/hl+E465UN7OEt92rrBbiBui+XoWq7CdsJMe9nKHrBHBmDe2
5RiRjYEodSEblKcqLRaKU7wVEUYDbVAwxDqV3oFlEPURsdFG4mPp9iIX4NYMi2Sk
GMXL+9VyltmBB6UKR5vvMjJ7rQ0nfYS75NsMfEzF0ZkbcfumIHzjvT+87f4AJuF1
yX1rg6rl24ehCrLo3Bd59NQrdPEinH1Bwutatrl/3CQA1S4dciWFOH8Og4PDUpdy
Jiel8VrQKSjc6Cc7Z3Qku4IcaOEQnK2yd7Ge+fqDS9oE4rvKKVDbCwzdQ1MyD3s0
b4vptQxLM9uJZyMl9vgtIBbItvsrrpu6m+cpNf4JEYxe86KXRbuSb08/q5tRv9sF
8LZO4Ll9E1/P+wX2IIMlyYwlwBlit+GldvfqZmMBUBDc7eq3xrxSvbDABLtgFIiv
qXsOZgTYcvqCY062/NrmQxH8MIFxnkxDy80hYQ58ogBE2LWXMFrBxUpB529EmShq
3xy1HW72j2HCyGIDdBgeAxbIIJ4iVwocBRm32AjGnanzw6dCNm840SOWpCdjl3pk
sYBMRgujGS11nB/EYNaR+BLHptqFC4OaNYRkFf/kY81asB1WJmzFQeJrmllMKyuM
xVhOKIkR8NU57lfS2UWY+mr5/fGscOibKRCFeTZxat/ujiJmjKAapMQhqCVXLL8D
1uG651qesmHLAtAy6V7CJ6kIM40prUANUU82dJiga57JIwKiEQVtO/hQryv0wpuX
vl3Y25BWhBYp5TGgZ6clNOthKbmMv88Ew8WPh0Bxgs2yJie8WDIXT0AClEfUmlw4
V1syMucKmduyq22hsmT3jaBwW0FrOMuDoSdJF3TtTY8HmMK8tBy/e5r4VPTuMf2c
4LC1FeAE/rumCxYZuYWVwmdxLPnGBEfteVfYBePRn0CTLB4v8kj+al/C9l0MBKBl
ZpGeDAM4vIwPQgSNB4oMn3HqFS4Tmqo+kWxmhAZCP53/LLOnSESoOiPIcWupiXop
WmJq1lZans/PxwVGYxvjYDuLsvIifhRUZCYYE7FlTjzpF8RpxTPWEGDmtyGohCo7
hpwvMkJB3x8dZFyRxKfku1lsXfhdR3g/WjXLmqAj2YuZGoWrU75ssny/YlZsmM/C
m2sM4cfRI/SK1ygNsUZc3Cez7DJES7eM0BhrPFVAdNqq7ZYPB7yTPW7IKMPKdry7
L/fV7Qs2Gm+Yp6KvKgIWGmGANtAUdfGVJQGpokL0gnh327FXUKqTHNHbIsKkPImk
P7Av6k7ByULO92vFjiBJBohlDfCkMs4du/1NQ5dsNxHHQwZOYsL4fmjTeAjz9UnY
Z8+xjf5JSFPcvvckubaMQqumFT70YP5en6Wa7j3egmIBKDjr1m1Zv1aT6Nazkyu9
9DQASFLCJNgDOukr15Fd8StK7K1P7nfBgmKDlBLw+KaVQcw3gHzkfzrwxWRVlN2e
pb1E7jf3XHkV3E8b6G0QdQ45yvdX16/NToUg1meIp5l6gNAbuquih27PVEvyKcH2
PjAiJMm2QKo6ttGFQ2ScNP2TCe/R+AYU4V9+i7EP8VVsRQ8ocg179GJVnlhLY6/G
g1kq78XJ0FI1sJsKfdTCPVLVP5el25CJmYMfIErKqU7nnok5G5iD//PxF+hRjPxk
utteHsSuZOkFIigj4AE/FaWtniNM2nnOtqAJQkjgbFp5BpkRy/QC1RHDlleM++uw
owpbk/rMwch/fTQ+WIomhyR3XeQnEDtECtf+YE8usgU6qDNAX+Nr2du+nW+DbMVV
jdddTWr/QtetdAYWAdCd8rYZ2GiPJBfO8niNWSoT0WlP5nGeoQLQLqM9bfQGPKPQ
WINsvcE5mNN2E67h1NBwgtOgLMaGlwWHom88Bo5mrBol5dSf+KjupJcuhIHHwqln
xjk2tuWtn4Uk9cHqPJ+M5+KAXhRy1/jJlLrKXY37YyGpOZUO09AHDvKuDQq7UIjK
UOhbBcSZQXgpQEBrr7OS80zy/oIlPpeXxuAgTD3CRPdPvx2K7z9lxVHHpl8KOgku
vvCmcbzzRQk9PxyCUM1WLBUB9Kd9UotOyhPwI+RoYIkabrjrnynoGBjYowKsjE8q
sRjUcR0s9bFfVZr4qb9keNxP05erNwDL5LIltepnCfdjVWzLU234jFb3UBgRiezY
dq6gkp/6dV4ffXwyAOA2XH9FPePxPM3/Z7oYsUp5onKcMtjopbyiCkH3e6kgW7YB
2Qh0gB06QxmuF5xf0NtMc+1yxBTMAlXSTpmOjYs8mHaZfScJtB0P9dVLh2l1rF6J
rLDRTOf/81FBX44P8oZJo/I5h8hVvilMjoF7V20MRaQqJA98/ia0G05vdIjiQoxz
PEHjZAeoKbA+rZS+hsTHWdWdouFpiqFUpxxvi5r0laz8zQ3pRD72DeDKDPVuNjNa
J4TW49xk1EZof0q9GwkASzE6KE62VcFoZZn/HhIDPgeyoEU3j8iD10x1lKJT/Edp
bYsXWVidb8dXHYoQ7siS8Q7tMXmp8QWHRtxTP/emBANVyZ9Rjkt3mPn7omOn8UYh
iYLbc7TLrdgouEeB4HtAHnCHeuHb8Sb2FTWfkBEj6zdAZ7kuv4/3kcpOAL00X9cl
haTnxFKgbk7LQEQFnxjON8krnRw8pVjUHWQj8PTssHsQEHvygS5/n+1zVF+5E8NP
6jNH2ZydVzYjHVlFKQTyaTQDFJr7YNctxWQpt2Y8SrKhgnoOrts/UY8PFEqRATL5
Y2gc2DRPknj5BFCTnGHjWtgevaY9HKgoDfxrdt0AriUM0mjj0lLeRXtH2z22f9OT
KR2VXsz8fGoUYyYCzJohZHhYjYkbE6jHJRbmHtxiDvsTmALYjpugN9nn7pQqDnO6
ygtozoxBgPmMhpCUUx+bfoWUigbiB8ZrH4Dijoj6umU8EZ32gyIBT0LAisdXoSbg
ho7pRjtYZ1eTsLg2cDaHWcSvmSynTlmhT0VKmqQvHkkt651CoRJcnS9j66CW69tw
2b39YZphOCEwnFNwuhME9Z5GXT4/yFhyJXzar7rwN44EzztcCVZd9ZTg4jPqb84z
IgV0H6Pd6R4F3suj2EBOemY2yCj9OiiAZU35ZNDKmGus5vsrFzGWapYTFKTSWjRM
MIA6fX+Bo9hRM1ARKMYFXxHrjH3zoqg4f4U/9y0hvUM8ZWJHtaW+cy9UWELeVJjM
YDCQB8r4LXY09nGTirMm/Y2Z+Lv6MCe82rnspWdX651H+zQdmOd92sYffecssplU
sgaPMIbm+0DcXhTcM+EDOOvxwjAB6lmivLIZ5DXE5eCd0zmrxsniLmXGD7B8SHZm
uyb7ity2YkUd0Ot/MfEbAzuuGPqHa2UvgbWGfCR5Ac3+5iX7vOl2KkmHfzD3qbxj
AAYyeqvQVoL5KLpuGD0FmksCKjIhu7wRHM9+gTkYQhXSDToR5ofrMhGu7/Mj+/AY
QhH5G/1Mbm8GaMLOH5kxEusyAnZe3ODUsGf1gq7Dnb7gwN2Vy36zrncv3rWqaWYf
H0uvsY9XPYGkkHBCB6/iBSIFa3c8NLRoHUi3S/j2xnIYAzbuDEqfEWaMpuXrVTlG
V0rlWjy8xaqk0tRKx0tT1fpLCNJwYiIdShdfi27dznCNH8A88mjt+kXRZ0FsYB4o
pB8DhA2uZPtc80cefbf1u1xztzzrz9ZmP8UQTEauN0S78A/TqXvypF40yWvpT4el
+DDhBBo8O5yI/McbybjTWoDbQGoz6VEI7ma+PC75bKKg5EQc9JfnUVp0Iw4EfkTb
zjHD7g4i3lmImzSekQD3jBaILf9UvKwo2oD2zYmiwirqNPx0JOIa8BTbIYFwDOFc
dLJy6f693g/jH2vLIy0/bL6hj2YlXLKrqirQobTV2fKuVz1bI9ZIOmrvL53+FFNF
yoWZ40l+Iu1TyvIGVUDgNv7UCN3ZNrDV89tHN8U29UmqGbO3egfJWxfy/EiKT1hX
ZiC0si5dajPz+POSs0b3Zc4TxCb8Yj0qK1vG3AjEw/fvSmTkv6TQKMVwzEIQGpRP
G4a8Nnks9s4UwYuooyn1BN0cd3cyO/hZnhUV0eZUV310LndE+1QHkEAz66XfD5R7
uBzjYgu9bG5rlh1XUbu06Bhbfjv/yUjqwv4aCFcAn0CPQQfwv/OyqtugBJjx01DO
efTovhoxGNXEkTAXr93h1jLc6H1ls79+PT7jdTnujuXs8qP7XSdQcEAjLflK+M8n
A9t4QGHrhHnvLBbuZHEy7gBqewQGeqGZPAHIIQF2P9OJFct/RG4UXFZhx0Gc5izK
9qUIYpeI9PfVc7g1JuHjNWE3AIcbNPKGqzrB6/vkWY7HG7ld/kOJKbxX9AJ15PSd
GEXcxS+3D1tJwrqcqYSu5MfLKFMnJhuY1+e+dLxomk46FNPqiP7ZgeE5iwIiwECN
FAL+U3TNrVHTxlOA3lz2ox9+mUKu2r4KKkEqdpFN9FSggI2Hf3vJt8JUf3Axsbm3
4HG+Q5F4Rp/Oa2iQ3zf2848nUEF3Phk6XBxZcfco+t1G+WfudgFm551VDnDhaBTQ
kqCK+d79zf2JXRNhk4FEv6IpWPM9eCh3oGxlwp+INDTQS7jYYLp+6yX+KCgGqslb
DQT2HyywT2XiRh75M9VxCS5QN3Rq1+SGDcDdjkrigljv4thxwdUgFT6a9FbCgTdC
rOvsDuyspVjYbEF23GUH2C1nKhD3FYw1JqwHQdCJIBNxZDxK1pk1uHGiE5jhJ+e2
mhOz7jKzZS1cOG5SygsN7mGi3u4M3LdPghhP7sxN0EkUf0FrRSjdc90O6yw6WiaY
jOcoZ5VhHSEEqV52A/AvzpGbhF2K6FDaFOyfE+YjfB7VDpZAyoXXLjGSMtSoFDMe
eH8KvcW8yo4Z3RFQrUgJ6M+yJRtwPdyW/vl7GU7OmJt0VTmC/VO+dNQl9PiQoVyr
30JEhOIrtnlE2t9hAm6NbaHs4ZRi4lvRf9Pk33Jmj4Pr7wU6vtFckxE04mWKGMKb
ASzOkmypXsEPapTAxFkteVWrpUge/Uolk7mi3jIAlzShXolRCX3b4AkA6exTXOiF
Hd9aT20MXgxm4JE4E5mMtE5V3GXfanzx0k/M/4CGzlXAYLy+mlrkh4t1ZwRQTPXm
XuhZVnEE02QKteXuljd5RJBGLuYvEvxJ+g+KUJBwsboHwHCPAH9HJnrumcmPgA6b
R58q3kn4YNI2ctNsWUBW+iWnwbzkK9ciH96m00aIjD17wUkvaujfgv4lUN5Cqo+C
qqp/PKJx4rr42+RyORS6d4QOlce4maOZVGaFjeUS6a6bYLToi6xbkWinX2Tg0qEu
KONfqvQBm9UoIEo+waIl/GHK5FXHJ1JvTog26zkYkWIU/KjrL2O29nCT2nRn4P5N
0Y30aDvhC2j8ukFNm/VOTM7kLcuh0AoojWFK2Q1+O1vGkSHi33uniiZjeJC9B5me
HAsN0MX++TBoy30kGdQcKxTR1g7v+/CxXqqH6M4NNc6BGVnUA/OSCvk19Sec7CwC
ggCl6IQXiyCnRNpP0QLXZWVCAMGwNNd8UXNtYelW5H1U4bvf12fBHfyNjUfVyg5u
yK5LuK69nffIBkeF8iPjWn5sWWQiB4SkJokau5BrgQADvLOrgJVFID5S59MFwKTa
6BXm165aQydpk0z2hxayF1YoxK/lywsdbclhdVdH8DrSJNkGB2xPB4LvnjkaEUnK
pY89FzPH3/UooiE8gDmEhzlJ8K/4dYBZRIi7raGapuNIgYqEW2aFrheFGKvB8gXm
l7TXz37xFmaKStkDPg3RpdYAG7mbjYO3tF+Rhl9DgOem+nUW1e2JEaH9stiSB7X4
GlDFBrcrfK9IT9zZwvigWVb616+75qHUFt7AYtbwiDRG6OsTRdOFDIsD5yQyi/5z
+TGdWhspr3ByFnUV2ldXyjXz8wpgNzuP5P1pDth3jUO+6u4rBRXAjHeZjBH1vFvU
wRQrXj2HJKKLubCu3zm4DF4jyXN1OC1M5B5wdDAfSvJhi09TbeNF6GX2Xs/AT8Fz
PCjwFsk9SN7B3u3w8qNhbnQKCUx9/k/TbbQUI7V/Jpuqcs/qbgvawpWPuNcm44Bg
5mIw67EWOYLhA2V201AFeFe+vAz9gVgwXQgbZ1LUe8bKG2EOx4YaIHvBq3cpB85E
NOCEiUrdIIqpFxhSCY0mAUL+zXq8q1O7zaVQIj3F7gg4qildUreSsHxCX9xDBcs5
4QxK2OAXObnjtm9IQgVCMAVtIsxj1iMMyjRohB9YOj64wXa2arMKwB03sQ3r85sI
pr+Ai+OVKA+H1iqFYkZCQ4L6CNJg3ZyXOZLEXuGTADl+TuTqfLM0bQ0u8oMwpGxI
OB/9sGksz7D07ncOzjdNpKJZAsbZKxbTnjrPP0Qpm0iRyy+0Ua5Mbz54ZpCjudQR
yMCiTrk3Aiq15f7kRUYoKuqaYcuRuvF1HoUd6PPcnuZDyDRpiCgr7/8lMSC5qUMw
2+Bk9wypWusJplfSdOQaYKq06teF8z5FLGW361MKGPa7OValY4YOaP88XcoOsagd
wV/7KCjDEP71pME9XTp1KXZfLWfBZSizpu8KWGwUxkVjVPd47y1znHJy4OENDr+y
fs5soPaj2+27gFCpeOEbgG/cJs0cSz91AEaYemwY+qcZ5ETiIp+xUO0teMqPGq/M
Ph8/vGHWJKUICK5JytXM9iEE66pRmts4hRZKJ6oJPRs1C/iEQ+0nrYTZvBb1IzXX
Fb531wN+uYXteH89xLrDnZ4a3q0x7hHpfhNiigPRmt2elaC6j2r0PMHsife0Jijg
QhX56MX6tiITq8u8s3Qi7WJOSrayb+n4HsKZMpXNfzU8WwIYZOBxtlV9ahq9ctnh
5LWyvpMIfArfy4WzgoThgd5g3jnjZhda9At7q6ksZgnJX/h8FJRr2crxRvRxYdO6
kC7vNiSmTP6ye+jObE15PwHqciLYrcIUl+I8Ilf+Gu934DFl5NWkhT6L7cFOmXH0
nok2x8kOv7/I7lE5FkI6Rb15ht7wYbkrs/JW59fL0SluRGV7mls9iLzeZNjRtCs1
NRJqYKWuZAhkAenLIC11vxnkzmXRlH6lGnuUJomUye8hMgLwXZQb1rnRBhX9T5bU
Hwpv/3T6VdGWVyz/zBYTgkNv6fv8btb4aox7w3HmVZWlEePAl5RFhs6H59x36oNL
GgmYOkYM9yvdBk92jq2rf84BLPG8iUodlR1behjld+1E0CvOZXff+UMcncQNWQGT
YBF4VXdXXxWR2mB8RLOE2mYegsEwjheYLH9PBgfdH8EjwCbLYHQIJEW1aDLlXHpS
3ZGsyacZBgHmdZg/nbMcjZVePzS3XTUiZiT+EkefrLeDumAOrY2eKJ/UKeQwi6v/
FDxbG0KstYwRXUdl/IU5ONS7rNrNJzkR47fVhsoU4gykNQO8s3flEeBaoSeaBvU2
22DkB+QLXedWzQA5rccaYwtyDQh6OmXldgXypYJOF5ixikECvrnwAk2RtcTEM9v1
f/hUYG8r58bWaJnH5kByY6643kdKQMp0KO3BwYZTfWbFz4en4hrg0GfvuDVfz73G
A5SRowOddoL5d4OloKJ+ltEL0Az8y7Z1SbolRwnPaKghIH0qZd+5IEnX8oZ0MU2O
YC8R/SgQPTRdlCulTmolhNAfu8UJJ908iAwdpAwj5U0KHG06/Fcj0iOLD3Ha+CKG
2rJlIBTKRhIim/q0ec+SFDj9kaPauUPZhedK+EWjnAv6qq4mHxjpdrGaqzV69dRB
n37O8dHDLDAgALldakMmy7HJxC3/o1fHNxSRSvKZV8AFuPQec6MqVbF+mzs17LNr
A+OnY5HzEpujKLPB05OnWkIVRmEFA3OniYYUlEkRnCIesqEcu9+2Yk6Oq6qSOjFd
X9CxsXQJWmaWM8RrdU3cdiHd7zm9GDD3d5PnRebvRT/qukmAZNO8HuBzOU+nvF4z
lFY2ycLB2P47uTUsSXPS1iYhcSV8tUKh5cYOv+462E+R61BUpXlltbdBrPUbeao3
1aGHY+ngq1K4kOlgX5K1FcKkpX398N98CkAAu5H9Db3CIdPMC8A76pME4w4Z7/xv
u1tGHcpFsoHzpHhJwn6FeCMCms/CcJa6juTlHzCjIoDxB/fZMfObq2OHsL4Hj9BD
TsH2WOplwZ7KBPgrj0PffHfczihhRBoopKLZMqxYoy+kEbBXmdUXavyhxTsfbjNG
F9PgxprONAwcscHL9zPeFtLRsJPq0zAjiJMQ9J13jroIsQsFfJYbVCQwr9Clrzv8
NI4d2anRgce/tR22hIm6zIk6ad8XeOlFe2qpU4Gp2CFCyBxQtlrxRB13WmYcCmEi
IvrO2pU3WKN++s+G4U3fEwzyRj2N5eGcMxZ22UQzOovhI8Sp9zRlhBs0K+OSxlFH
uXBssgaHE33hU0irvwtnYntG37DGCB5YTG8LLQg5niqzQngTPFs6L1030eI4NDGy
+iosatpEF2rmkQKLkTEfGJQx/1u29OcDygJM6OjYMhhXhDeSatKjxvp8iLHoeldn
Mut3+qXHhgc7ihJFxbpZAxjDfimGtgCNe8li5urN5Dbp341LwEur+fI94HQbJ6Z1
tAOgyjjj2rR/3LpPMRfb/+Y+CVVo9itokUDhNd33ntjsIkcjpdANZoidgGWLxJkK
l3h27c/Q3nXtBrR3nF9mCimV0nrLNWmWpFcu5OJtX8Oim8cQv4s2gSIdTWxwKYJX
QtVXKEVnvWZQbcMkOUSQE2L4zTy9x41JndzDyjpRlijXG6d7NrcycHcZRl17f3mE
3+SuurBQWB5fAY17fvT0AQS5hcMAhiHSqDxzuu3ptwGKIyamxlYV/xzSmrzaL2Ml
zmXRfhdtgvaZCfffEPLVdK9ILLSQYycMHj5P6lDBsKAQFR2fKijoqM5RtEKMcNeg
3FHIwx3DHZkoekMHKCcMkTIwNGPt0RilMnkHAeJTh4R2Ia6sAN235ziA76dUtaie
5htt2YwxyVcFi5mOZgIZwG2FAC6t+thEhdrVQ04EhVd7SKekMzAxlhTIkmPZd8Lu
WWD538QpndBmN65nT0xLbM/HimueAEkuEvGF8ucrVk5zTea2Xfcxb1v14iQZ4hCp
Vu9Vy7UhpTUWN9Bb7+/tWOHSztmB1vDzm337sRkTQ5Dg6y61HW19wxmnz31ajmjj
Z0LVt3uiOlMnFpU6Syj/PJ1jXAYm45cE5ZAOCRS5yyz+WUMZzKRaxjDBWafYrT4h
z+huFKZJ5s2rtnl/A8xcfLoFBgERW5bdB32WO8+lWy0pPdZA4QRW3PgJ8DFni2dL
jPTzONIrdlDdSzBXfMw8v1xXXnMe63Cmk6nYZVgEjrDlrIjNgIXWkJUz8UHGsrvy
/uJ3n4ecjfK69j0KE6wvOaEmb2Esy/i92tI7hrAWL+BF625gLE8bgyu1b1f9ToCw
RWOMeDRVhp6obX9N0/L/TpyDGPtPF11nDdkHzZUdZJO1y569rghySNL6F4z7Qhd0
g9D+mCShPaad7XnEJVgj9QWsDNwpDy6P1/5dhJ+HPpvaR5vC+nxHrc7P4oJB3HHg
ob9VJ+gNeK5IMnIEREAlUW9iUchSeZPT/yU32AOxVncA+c6zP8ExaitOmZFfIrJr
s+OiApB7FHcaaAMv4uuZcA5KfRD3GJi9w3Oump55CO1iMeQt7wdHIxvKrtrQeRfc
A2V8d4h7AtIQD5IVE2Q9HMW7eOQ6U/RXzyQtI+F4rSYSz0Mz5iTYdclD61QbYVc9
XR5TobmJHYq6dDmtiOkfZzdNEcbQPr+cdNe4nhdXcFQQcN+z/TkrE3lvjFoyP1Yo
q7Ex7vU8hPzkMeWQGpXgyDk0FogzdpgPdPCCwPHx3LMky/WFL1TjmiBPQT8v6qi+
jPDjXRdEV6EAQe03Q7Zb8aUawGXLxHJ6dgxXLRZfXsbBEK6H/jlLx7zvY+uuI10r
1SlvSEuj5zdtdy7/gBh034t/rE6CD8iYR4K3xwcN2NRoyNS7B0LWpKwDHQPIrqQh
A8RogaMMuQ47NdAsAAxpcEk7D+iEt1xyFYdVoLds6MMXnTgsp6WUp7Xb0KYoyHOJ
xvoglee14kXk059iRZzSozdLyc4mquWI9CKqzSzYDomfCFtpURHbEt5Np442rJuR
3KSXEglDFVknftLv/ZOrOCdxYqHodVZTqr/y/HtEELGnF95l+6ypLMwipDn54UkP
7IdiMpSYY+98c0zE+3jt5pGCh8bElyM+bsLlnwTM3cUjqxtPUc4whoveG5fQT1u8
W+R2kWtDkF/nO04v8OEWQa+kKAR0Msi9f7qpcCYF9QAJC76OCysAWxhpAojB1tpB
ByffOfQOt0tUkq2oQDnqm2arHT0IC4lLCC+u1SZmHPqlisz09BIYsvlh1wLgbgYC
bPyV0MkLwlJZ/DP0Ukbk04pymHqyf2QzTpk3HN2oE/VOJmpmiWyhArnUx6nS5Con
CjcVTRYmI3luFW2NOistGH7H/Qqotp385jTRluRhPqeO59r6c7LTDghlrdIG5oQL
z0zf2AEFA5PgaUZINUBAqZOh2/GXqYkBxl6CgSK76rSiqY0YOLOwPETborpQCLL6
qHtKvP50D4VM4PMcCjMY8aK65I0N9hK3ukb/UhMkCgO6MHy8/ZNkLGTq/Z3R6XEQ
ZmJZiQmt4072x0fGRMxwCg2rVu0PAhUuSft9kjOkRATe1TQ68+lND8ziBOfbHnlS
ORvzKuMPVIH1GMJbBiSf9NcGqd4zhD7vu/08KCngZPADGQfT3CZ85fPIYibEVs0t
TfqiQHsa5JJyNsS7uTw+lskzQaZjhlcGdgce0YxJNPPrIkFsSl1442m1C0bijHog
VgfNrzCjPtnehIkjI8nbe1AWdpX89y3b6uVeXgedpbKkDYiq2ylQfivMAkuwinzu
oO/7sijnedbM+bS1S3m8iS2VqarWJeZBlF7pwyklSr/JWl8IdqPK1RV4RPQ7cz5a
1UGwsp6iSbABkzBrTOKonP1lXiGy/ojfZ3XP1r1M5LvCmjw5Gsoke63kB2whZ1U3
kxmwKcFReWGXUKHCjAM+fmfxFbmo0pSPtz2sdt9grqq0SKHvUcq2y72s8Up3kXOI
iUixlxZHFBibN88p8kt69swFSwrgmES4vAdZQPURTEw9DXPODrzKM7BrtRilWyb4
k3g4Q4leb3CYLMW7cn2sBugV72iyt12pazK8Lc3mD6bDFbCW4z4TEY4FgqNkf1nZ
zRi6Yc8BuyZ2Js8wA3VXgHSmGWcxNBUL7JCXnWvcKgPnkc3gyLeSlS+Bju+mm9Bx
Kg7I6pRiEVcLjMrUWGQwNK+GY5ytDB8kqQlR4GkWviuAX5nBMV+2Gk13Mhm+sasz
Q+Ro3nPC8sl7L4G+QvyNs/SOwFtxsZn6K70I3ebqSggi0R9uevyF1IwFLotA8GMx
0zDYv8ENF6S3U32jSteRBTwcJD8EcbAbPc4vTwaHfaXdMGSmXDEHiGwN4YCaTbgb
BfeDISXFOJNwSVrRBkHPMwZ5sXMk/3WYAp2ZtELMKYDVbL9BWizxK13el691FHO0
PZ3W6UuvQQyPPIFn2NcskS/l33ssIL6GIT8E0X+WZ0zW522b8/mSg+JzntsUhVDg
tLdg/aJIzLC9HlEqC9ZSuoSOnPwJRClmjQ6FJzSIUCB1HX/wpy3li2R62PuYvhDa
Q4qrwU3bBRwx7F92FjgAcNdO89FUWr2zM8LE9R9piMETpPCtZWzyNd4MdNICyJxD
D7g5yUAcSfXJR8Ce2MvfnCTrX6AKEyjRzmnYra8061/Tku83+kBwD1roIXeFYVuG
df0rTSOQZkTp9QYyTHrJ9zgm0WRqVX787JqZnGKEPpxqbiT1Wr4G4geDDiIXoZTx
MoevdM53A1JQlSGyjpANeB4w48mIMlQ5EoGHgbVmzf/lGeGCtWaCRMPzUh+Ngrkp
yhwU+YW9GafqSZY0eLMp8lms8/BGaMt4gzpUAgrQpJpIYWKmbqhdWRMv7eaiN0q8
e234FJHupXbmamVLbiYyE5Is1pp6pAR6/rplBLfX9d9se803E3CLBht6MxZ7mrBb
DvoZvrmqxmeteF9znjS5BBxTClUVdy5juN6rVTgjHTAKSaJQvaiMASe2WbluhIfw
zZWVaXXfqAtc1kdSEUqN/R4oQ0tEjxHX4kTLB3lT82jnZPDdKikxgqX6HW2O8Cfz
iOYMEz2pIquf6Q5jPIw0+rHIAeAOF4ZJov/+un5QlMgEYJMqD0fFPlLoHSx9hxUP
ft/OCbv7JJZuB8vJftguNkIGtxiot1PAgR52JEjfWJKsU2YCikVsPZXlpwmXKYcj
cOlkqyVkAPbs6g0NnPjaFHcgSe3lWrZzsJVXcfteKeD2UOb3cCfIUuvRYW+LpDSW
0sWPd3tpTG+km5+2ilZRvmsmB6166fjU9mvgHsYH8MebZSH4KJG+M6KAnl3Q/I0x
1xn241tDq94VTLJQ07DNA1tkARX1bo3q92fL5pqZAD1ZdiWA38SAezmwVQbg3y5Q
DZGWP7Lt+0xVdSI31CbxIo1Lr128/mfzLU3KSENv9tWZb+f0pEZbu28TSDDkjN5h
sKdYF+0wbcBE3yUOU8qN5uIHuS6KHu4j9JrJBZXZ2r9UvFa3kAErKKLZAJElcwnw
ELOc3BtmROVRLLHnSb95DnhVu1cHFWJZzzJ32b4QezlDenJEatMCyf3KWoiYE5Ag
BQ9Pcw2ONsyOhWzZyKbXKPjBajgiRp+rS/GnaGeVZFdAf/Rj0E5qstBz4aOhkvNl
ldcIq2C5L+RXGflbAe7XDUBbUIyibVo3h13e7pQq1QrRme4EsA7U4hnb0r5RwqzE
jptPqTRlnjnwK35PFN75xE4oJ5xjr9Qz4wtJMwMHJC072fxY7VYDA62oxhlNukvR
Fz9yv9TwPE8e8dhF89IWvPj+HIFZJi2FOPFSS8wevNrsLzq9r1cvfabOniju05O3
QAsDK8ulwNSFMIs9JUwuFUwAhg6YaMJx+yFWAtuEpvLLtP6EY51h9AQB+e3H9HAJ
THMZUdHYK2h1fcEVWgOzlIu+r+IlpRovS/ZN1KRQB9SmHPbHm6263bPC4/qsec8P
k0T43mSX1VrYL0iPtEJtWqHqnVEJOu1bvr2abn0xukgRdRcM8poPY7ma0zZ+8ZxT
/XLmg0qgpc8WNdxse9XHK8mMVkQ2Nna6BjKwc0gpjz69U+Oo/m0VyOsrEo9aueaX
xhX2addBvh4PT9Bo+pjRR7WgdwkggImk2jhnYi5sB1UfNCdT99YDYIwUECHpvJ5H
8hyvSFr/naoJWdGg0IPYSgpyC1OuqTy4OVhGKAQhlfsz8gWu9qLza6LVyzpqzmxR
5oJvMccwCaO+FJwEgcdidtMnc8Bzt1igq37hx3Der+mv5vBxomkDpXmpX4phVtdz
NhLfKfYaHSp6H7qtFBVHGAniYhWMOtEDFf++KVg2GlSTyglfYfDT0M4CHfiel+6W
SlMpnQjiYaWWvLevxAkcNTqFYKhVKve+cBaVEs0AxAZblslUbxdvrNA+ngVVKjwk
YQfPDWdmJMmQyfGo45PRxoPvnDI3CCqdBIB3gAbz5vZ+1M+6nB10jLlZJXddof4t
A1zfV/t3Bwb/3M4MGGU8ZiLKVGWFmS9WMqHUNQDjUSRizp5YvCJRcvliCvC2nWOG
JTH3kCi7ABQbBE9XuMlSPAzZ5E7ym73XKpoEpqOoyJgqq3OORiRAvKJqc8AMRGTR
RKGbFYKUHSwXEwLA4AKohwuS3GYrxVMeEGDmAgRL/lB5XMnw5JZJCtroltO7dHOV
MaDyK80DMKW4j0L1ZrO5tmNcOFeB/R+f/+6xL+Y5XKTWz2Bc59RKXf0cOSpr2Qbf
VpRafwrUo92x/0sPT+nYL6GJAHfEO2rhlhCRoVoJ97joOELL0u3wdW3b+dVOZk4l
HesR//km6b2w8WfeijAqgxY5hGioT26YHQUie3/kPuZO53aLUcwV/iY4kJ9NWWQy
4VYine8hx6TZEa8XAdc07FucVl21Y8FuwnWi5/WJPh/NlPd8W6KJ1zhGT24ILSew
aBpBuWL0MiEmqVIwn84+0oBKkgcuFWMXkznRopES5EtepxM+yrDNSvDJ+zSvW6xe
B9SAa3ZCPaUTb0K9QGyd3Fw58slZ8I4nDTYhHB00bAVWCjzVRizz0WFBp9vhjvST
YBC68+t1UE/YcPIU9iWS2n0nXDNFlSGP00OaP2uAgVnBeE0Hwy0d3gTOzL3zXNao
n+T8BDCo8WWsR8kjoeqyW+cvevyckdWSRhCSkCK5TlL8zvWUR+LQVHPiryQn13Mf
coFG8VHQ/D/ID9afpliAyu4uJRFIDmg9GUU8lq36EohyNGopaOQOIviccjJg5aDT
yfjW3UUMtNj5t6aZSJbMVSUD+elovJbClV/h1f/M+6prYm3D8zB/QbNy3clsTPgL
sX9vzUbjPwIgaqfeFlodBB4y9BiG5k6477ON0CGV/Nj82RoDC0RYk43sxZ+QmiWN
QGye/vPZ8ApiTvGCnEEdlRmPuqDC6oQQ1PruxzMHJUytB669roKutpICRpWmgJ4O
4jLttVK+4U97yJEVvqEN5Ow3gAmvy8sZcGXVpfwOtiaLuWLyp9XBkpNafIm8ESkr
hmozzlCSq4ZBK8j+Y7KIXH8WR/8VeABSAP4ykF/2vktpbjdAi/AH+wg680TDuVIV
9H4edGA2pSjrvbAAM33CdkjvNZeb86+tIxIROGGRqLo6xHjb9+6fkTYUBp+QUQhB
08gEbRi8+86haD+kNlYsV8kxrHlOIgecxyrLkCHJY3BL/d/CdINrywp9gxkrxXAV
mACkjZ0dmaSFSIlWP3ystkXi6O5mOIRFmwNGgPTYkTeNnYCfo1VLgYRUMxD92Jr9
iMPuoSyl9ZT1PrBZPHgJ7BJuNCfKuFqWmrpsOToYVI63VB7KDEpxLOOc9Y06VoKm
pNz8lBXOLSxUC5O/2Y2H9UuvNsHXpTr8hCt8bijz4Piph8dYo9n6g3rujHohh3To
uo4g5AKH6n4rtdBtuRM5ke0h+CAoWWwJjwepV9zKxxZ8/Bxfa/zBWmyeX/IqxVZd
UDIlSBsaiBhW07ctJ9G2a2v6du4VCvIkjbVJZ65ct2nufDYdXRIfmCoAa/eZ2xDk
AfKSAHtrzl8uzPXeqSP6Sf4n3T5oJfE2RFgyZJYz+81UzQAheOEqruT/5LzYiuQ3
eqLte9ME80GZ5ORE4mlJ2Y9S/EfBg+qD5a8wRTqWi94/qsWi5qBmWNSIB+eaZkfj
JZN8QX8KPs+VaA7LpP5Ge4HfDWlqfMxGuhlvHuqywxtM0BYBHXt/v0Wi9Ed4hB4r
TZCAj+BIJ5QMGfO3VeVWF0a3N1749Mb1sD2IWz95otAPdqsg+tD5zU27Ajy9s7IP
WdJ8ny/zrD1nIsWGgYb9ngD04IM4P8c0aLe/aPI+2AgHHGisCDolW8Z72T8tVBFG
laUPUbrxi4J4xMx1G0A1QoL8mmXPmSNokca19YuhAgHoibDzmnqii/85gOxpZNcV
2HymhbCdVpAW49wqUo8gdxm6YyDKMAWmNYWRAc97TGJUDWy5URYsDEYKAVyrCDQC
5N8NMwA53HoEPxwbOZRm7d6SXbp6MtWSb7zxm6V0lWzzWHkBWd6RdVwrVd1vs25V
S8eJto+pO6532rYnLKhxUYq6V+YId42FhEgI/OeI2hGIH4MkunC1oVsWqVyBrx48
5GxjevyN7/bNlZHH3omJj3nmaoiJDGMacp1g7O5dVJTOf50k2gWeLC3i24jD3dFP
j+F2eRqtvu/6OSMIo6GYE5q1OnWLuZ24PqDWtQFVUlAJOV2/DeUdZu85PGsL5cNl
m2i3Zytg6Nx54EDOru6ESeatADpbmVvqCtTtdEU9WYWqDYwylpDwu0LqHNxaDny0
cna2+9P/i66nJ3IAquazGW0aCCe7l94ozq1FFCtLOjzeBMxrOA8IIwChqxKrxeDf
UwdaLyrm5XXWV29FJ+MKR/PK+6k0HNXK/LzM5lhHUVwnaVsYw14QIn0XEyl4ILGw
cQL+kDccCzrz565CKiaE0vB6vpiCWfITR7A9e7fivyDmorTwCJBF+WC7Tf4wUCoM
WwPaAyh6o113BPiQCqf5Jkyuwwcp6P5WoRuB236+uG7HQDfi8G08soLtg2YIRjBX
C5IMjMjZrc3ciPDEwNwhmxJIrrkcEFKnfIvvsAarm7IEDbeH6yVsrjjL0QE8b1jK
AQZ7BVAWpwnRN2JUCFmbvNTaPmUOa14yLzxHpTFXom5ELkVbUQo0gv3PwZxQ0yiJ
z4HNIPGRoLEUUBe5t8Da9HSDZcFuGZJEpbngZzsVoVEDIbt2c8R732PEeF5OTD3A
0FChJvMmhwMvL+E5E1ovCAgjFh2ih2EYIL/WWvBDiXFt6Y0AejMH6P1360jfxAcB
J725e6S7ivO18IQSvoeWCmPmSZPO66AdRdpJRXr9/ho8Hku+r7I9O4go1fgh43Xe
M6CY8pshYo2P2LNipxKO+evCS4pcAiJeh1DpM+hLd1RnFOZgpZlDhieHNDkXKqK4
jSccBb7b70gcHaZzTnSSuPIyyPVLEOOzXa4sBkUYyd1IhB29vLeBzYwjgjTgPex4
N+8OAciWx05bNe1tnR3HW5YRog76tcMa3PujhV8fjoBDMxtwb/5E3nkyWwR67HVr
6txt7WKrDmoG+r/Z+QnqkozZ1ZikZACpp6kjPIa1ma0cr4FDmErf/2iNTI+/zm14
LU1D5YjPrxhHBfRoPupZDIpR5z1ujGtsJeZFAmIH65REAlojD08WmiL/PSZdlTH5
qIjppvsVwu8HXlfy6VMRq7ecxEpDmwgqT9A+NNDCMXliPzUjKQzGxHaymf28Qfwg
D1Z1r5xO1xhtLXze4Cdy0bBsbhOnf8v5pZW2z28oYzB1mMB0eQMPo9rXshowQbaT
TmofXdzn1mIdXucCxIig0yjvz2FR53UBh9Tss8q5jOseFUYTYSHo2pbD4z4QgdBU
MlVo7RDZ9fRAFXpYGZmLi0MU+Z0P3IRKId/4f/+IJGZk0X9l+1y7Ui3BZT9eVYSP
gfuQ8ajoDBiYcgzU0QVIr4YdMoEvMSRhCmnnNmQnKFcibPTkIr7ZAKajrh/9hNNE
ZAi79YbURcJwOY7tlLrWPtqxxzSvTGKpABDaOOeuz8f+kGFbWOt04XHPzNwwokGe
CGZd31pILalfG24EFKR80o2MvWBByBSOtLvE0QQSCy41SU2Ilf8xML1L/FVcKmMZ
p41qN56sj6CpSJkoPL6QFkcfWhPC+VQfEDzwLgljhZnZv6A33/XwiZUuCeILqjSL
QafENIwuvr8U0BMb5HPELpLe33DLYg1OO/QoaxCGFu4Ong5lVbAUVoUTIApce5Df
MdBctVsbPjLKLZlVTa86QlXpNVabMhnzkIP97aVcGrTXc2mYzkMHiLEgcxTmxJ6W
+wu8SQqacBEGyXmbucIDUk5ns5JJkERfHI61/rbEzjlFdpjnCjZv4yvYCT7OUwVt
ivSlQc8byU1YKYU9FYiKlv+aML1e4+dDln5zXlAVSOfSewXA5NmR1s8EtUC7//Fm
COuxkqDtAs7OTIPmzN+p+S1qJ1G5WPAY6KLeCIHnVRfZEChZeQuZLPqjN5R2/SYQ
nf8iFoVIVCxDaA4BDfNeUCPtridJrZK0SYiyO+dghGCGRaQj7rIqFbxPL2bxefoP
D9PMl3ybRKD3l+aBWOHZPoV8bmWvyw2TjzBXrbFHbkpa3US7RuQiEl31odTKsEo6
+jL7UnSEiGWu6/tQ/qgSdqNJb+ff/aR/3h6DwGek4ajVzqAizgwp7Lu8zhTL37Ph
P/KMwHKdv7AdkHKY5Cp07kz5c9z1OXjfjsm3uR/FOB5+Y9MDMuxNM56LehQcztzQ
foriFhuyuzrrA/WS40eK5ieqSOTtoprcSS55thAtBoJWbu7PzfhTulYvtXfKPDCz
sqW2phHLpruDJKneXlK+s1RZr3KMct4BPbjaMQSn6RwzIapS0mMvIpZPBKXuQjuo
2VantPIYVDsvrdlQgCyrZyRB2+9TjHSnfPv58+cUYSg34xDruailg+XofzGRCwWZ
hYwNm6f7M/lF3pFqrnjfTYAhWLP0JSx+YTCSj6D18MiSA+qmD9qW8vR/yhAurWhF
/kp4D0Rv0NfOR+Y8SB1sPNLs5N7Vo2dKSxb1Mbb0VLoE5UkvEn81oAfIdHXjx0xk
KVrsiFfmw/uwrvkgZMS0pUJkFECcW7+lTXJy6XiE0MvN4Y9hqdVdCYxS51fuMKiD
osqA6b1/1pAZh3yvnKZ8CbAY7ccXnSZRd5pzPToaAHXUho94MQsLMzE90JYmuUN4
RbDjZE4fvVo/A7znTADZtOOuVfrh47k82IMN74S2GrJyd2N+jJTJ/gRtA9/CR/+9
2y3CFvwcKAwZdHXwgFR8rl+cXaV6UGUGEU8Jpr1ZjFRQArbeufrVYnXWeX0CcQTh
iHfmP2S49nySX9eCeA0X6J4OZGdeBwHAQEkx6aymyQGakDWoaLpfPoWhT+ySxc/+
WwO4hRXwrelBo+1mjWq2ZoG0SpCNE1HIQ9C9vejP2VabS6NySEFYzlXKVsnsrT4+
f2JZIACwqbXHLbbavvjbQhb4nNo1HsjcYzcov/5gL/Wyk+KZRe7RWMUziRWuNGAN
okSHMVhCvsHPDmHTtFm9ivDaXewAKdCVfZg0IenBE5z4ARtL2aNn5PeNRwYJcxse
UnuATckrHDMFhCqt6muyf58yXUPG3518QlF390X+crg+SHuo1lIZe5qhnsrFBw+/
o+Ysi8d1juHyE3rs0GO+tEyFGfIqv/+qVeNDCoxHvJ4B2mIcrwe6eYzsZ6bx6UsU
GnnRScwoUKcNvSFw1i9lR1jnXsBNXkBax+pp92PS+dse94Y/pvCYXJUEKQ115ixY
Te+fZazSb/kEnweV5J6nIxTZJ2E4UQbeLInxfGXrieQV/OtenKIvTyyD/716aLDF
UC1zDsZi0sVxeBKl36SwIaKryFYKLNxQiPhGivnUsMetbBMsjwt9RDarIDCfzVoG
QvKy0nO95S+UvDaBstHA9/ZKuv+rFoozKVYXe6gEWGEoZXiJs8Vi5HoL4Q46jfRA
mr1X6WhFO4xUYeEb2U8F0XeYha5QOiTay78aXq9Jy4+6wN0GuVV2BC2NqoKXS8aX
9sv0jCztOwxWtw2hmiTVhypyesG/1AC4bdZZ2/M13ph7Myhm2yxPWeoeZ2Qg2Xyh
eLTBMBmnQzgrs1sX/Bt0HNEc7CjjceI6Mr0IqLjvZATThaLCdobPWPSsk3JoWRqv
t2+wL1gSj4fCKe4EbguJjUnsUuV5kwZfBN0RdAb7iS9mwyTM8jPDwq/iQrP/B9ei
xZjspqXnLQkoep6cNcd5WUPGE8mYs7S9rB27gWdMGSVJxdVN0LGrjro9dSDXNyUe
r9+uYejeRRNrSB4WbJ2O6Z3Hq0qf6MvdyG9Np510MHCgbcCCWUISZWsP3znD5L+k
lFdNWahyAB+vEdhpjng3EKC5L3K4yjtGqrCZSjD8OdN7EV35iZrw+zoQW2w6+Fqy
a3dzttgDSmjzQo5HGttPchFsv9tXXNDscSf0kOU0nkFNXJ4jKl9oMLcUWqyd11c9
gbU/SHfkLmSSpm73HXRXayCjUIruA1grgF2TUEJggFSFMsNNWdU9Ur1IoofVkLCE
LJVd3OVqwPdyPmUEYI2MKaDtVVmhH8fCv+7HLdVkAwjg7sVeGcXJ3tZiyLDMSHqA
ecSrGvcNSvTAWrCvrtYQIMdqLY+iPXTLE+FMqbPmLKJw2pm/pTMt2YAMYwa8eBnj
8RLgP8PSLsjDxpTKFZiaw7uIokijsreT+NXCyl7+ETOyZuaQaBjI9ahp+bfCvmt3
zPSkJxJjpFOHpjyHGYnmBb8pb54YepOVtgZ7XFHV6WE4ZI0DlE77BRwcWbd8ptlP
2T1xJOCopT2ZzFXsmYH4OZn5sAHF1PjYCq+6DfX25VSd6DjzPqpb7xIpg5/LzJOB
hJC75BNFXhEGUYYLa7PHb0mI5ODfUCX8GLYEf3EMx32ohfd6PGfQ+YI1lvk2s0Tg
sfEc2FOqHwOAA7XNzhGtp7C3nNcNKz9zIn0pV5XBhnjLe2WkeN4IJ1TSxNT8QFsF
10CM6UtdzsaWLiQmrc/EIVw6gHE8BQyvlff3tMkC6jqIM3DpztnAlsyuS6jvtunX
l2iC3RADXTQLE+ZeGXZRZLV9aULOcgV8vTWAlQ2qvPaBVzXsnqyq5uR5G/nE/kdW
vVnuXXBQJyfrxaGi/b4PzCkXCJ+9lIO/oK16+cKsiW9P2XNOuG7oULIL0cDxbjy4
XoyFVl8VYckV8dmgCysZ9q4RuDqm2TvWcU4ygTrqHjKqjl97sb90g2ED5YhU3t4f
LJwP4uQPrvAgDbc+RszBA42Uz5u0kewOqZ3LHnV7vuTW79JBWYSaowIhIr7w2VHm
dcwyFwQEVRejxxHWkDiyOJkd+HpuOWs+bXqSUkwK35roSDMHHUWLwLKB3arK285p
11pjLk9TGKn7Zp28KfGqrXnozVLfCNrIR1nNkr2bTkKFVTbf4q72O9GuQdrxhLSg
bOBMR74XG6FGMQAqAfPOPutY5tF2xpy/cjQAmTw85hYMQ1JYDchNpAcxW+o7sn5n
6l8CTqjX+hLIn5LQDxSFUpE/6oBQXHAYh5JXW7pPTjnDgDDiSLJuY1luzGsCXspP
WhFJ/IQyLa42YvsJtnhcTLYov3+ZaZXdMmFGG5Zo2Ke6zdHY9OlHoUAcQv+C5LQn
22rcfTbSc1pZCTtulb1KHRCVP2Lw1DRUrShYsEs5nuAqdamtuOyPuRBXTYAcPksD
HQJ8LpUmkfdASpy1AIFCv0tVKGRqjStHmrrDAw75zmzGNYJzrXKjcvdHlIWO+Dy5
yl3AvZL0OdwaOqpXSz3827IYrocYQnOiNDbIRv90IzA32zie+7/ICAW1INpOqdHI
A27Jw5fcfNam4sGffX46p+JoyJO1AA2PbAMCzMKScYPoxg2bMFCQrw7l+UtJdlA4
R6gghncKYCgYdZMIuD32+FKoSAwxpDPQrSS5WYIQu3S2NNcdCOueHWvJ3+cNVcNK
QXdsr0QtJAiWZljGpiyHvauE3d+j/g7BWOWDKUMXfRBzu0iOOfcn+dtC0aR9fjXn
GJY2oSpzJcaCq71xK3jX6GPRJlvu/Hv3aIXBrMbnC+pvkh9SMjPmiBRXk2mnApJu
4KfnfQkhhy0HuolmQiOCy1S1OFUI+4ln2QOGz8ZDNQwCQewA0Ah+ybcwDTfsYxq0
dBvoPudFatfqWTElXKXf3FJhRCgt+O2zJS6jxhArJ+n2eKeQKhnShBe/lSo7Re0H
tMkNO5AT5y0Y+WpnNJz7aN72uSx8JnACvXoGuJePmddUB/gEh/aqSI/+gsvw+dRG
YcbXErBu+ChWwbFxjRmHQo5HjRlc/ehDjYSvFBhufFYFq4CfNxupCrx30Czn9wHT
/GUGn9x1QuxL1mp6h0WyzH72/3VS7Fg3MtD6E2/B/zoDbgf5pgWwjVeqgih02Nm4
U3OXSJqfkdZ82DxHxmH+yHuE/P4YG5t7uzYd9i3XKyYcj88ejNL4y0O/B62IFZlf
h0PYra1Rnr+BCMyWkoWuWu7qyFcptLdUGuznDQCD8PVNXsnP1mz98t111MA8HVAT
zeqcekVz12fZQah0/dMvCCX3ehKU07Io9Cf4cI+42gIzntwCTpiDZ//XwhCq0Z8g
v2l/1YYXhSTx0gvnKr3Qc2r3l7I0VWw+1mB+5vqtn1YgoXnIHnSiEwatKWy2LXty
wopMSQcmAcBjp3hA0ZISdU3djGox2HuZ5HXa4+3t+53DCPyg3bLYgoRdnQe3nIoG
fDa0tFSsmc3CcPAaXm9xA5BYUA+Qf+e5+MpVgra4CRIFoaTCnhKMUt7dXQ5mha6c
9MV+LTD/OmLp7gsib2j1rZjeC3T6T6c/pSXIaMEZKxBfs/H0gb10YC1HNgQtou6V
QQNu4uaLhy2EvYwGOaNomkjsPsfMbToXpC/Ba2vlsxulIDO2ikuljg6b4KFka4Jo
SJBqi4mVBsFWRS9f4Z3gHn15eM5S0AjjFQGLIg0iu3Wa500nvIAyYyDykS5+ARuE
/f9BNylBJsnFR4qbWFRYIZ6FffnLdN4LKkgNPTSW8A4t1KAim2hk67BcKZiVP5uv
ExV4SVyis/vm3KI6nz93zTqoZBEXqT7M2cee/0+8mAqmjpB5P0fgPnsCLTOWoXgr
/xTYjL9+GQkCPUBshDCnxmvB4u3SNr8XnSscjWNH2DQwTVsabW6/IbLi9VdaQclX
SGn6h6voJWEgK7pHNKv3fZPjThXdfVhzZJ9ODqu+YAKmOovVBfQ5npCbYqTMfzBu
d+SypBRPNPzJXhqlozUuZ82rAmaLLwT961PZZ/0F+mLdyCL8Phy+iIAqxiTkO2hJ
qTFXP0lC+K56Tz4yS0THZcIjT80Diwu/G7j7+WYL5u+azvY+9IBXzl1gwlriLK6k
myPvvsWH0KDIpdTJci0jhcvzP0blqRnikZ5owYvC8E4X2nOVR4qnkuSLjscbFW57
OZKElbUWTxhCSBeJtPyu7HKBTjZ/Cjaq90AKHuctPfTgtFrfBqbwmF660b/9mEJz
/Mr1daHXEbV8nI331nqfHIr55h9pXtkOIzJOWpDScyPlWaVO+Gog7cveeNaAs0yA
0h47RUMT7KhVgQi4wxSs4DR2AFfi+MvG27QtoGraz/UgbBZLllO2OcLMy+bnNTne
QEYdJKza4aKy0YXAUaLzGeztwy2CtEaLxCs/J+l3Ewjr45f3k1kIEbaFsMH/ju+F
6uTc7QyOFE5ioBNnW1w3vv2hfr+cfTNVVEL2CT7Jqe/rHXYiwkYeApsV+moC8yxm
anLmfW6d1Ee8LSJMzjGYinJh8FiMIhtZOh/Jhp3Kdeydu1nQzFgiaq9733DkDMJJ
TBHJ/yECHDFi4G8xezJ6f9MC3ptO8Kg++zRhX6xfR70jpp0ZWk+RUcvZPmohiU9X
N1mWFpmO83275UDsrjQycRAVU9Ge6WGpYj5KvSW/zvM8wWRC7MBLAjPx/KtBQPvH
JlcSVU6B6dw0SDTjRzSTi7zV/NvxtEMzqL2QVOkcleETeJpF0p9LYFn4nkbszLin
walyeen4Y8h7SmU+ETNEnNVSRCUOdez1GPbGKwa3EBw81xBsXj/sCM+xN4aOrWBk
g2rnmAc+FBSZK/nfGJwduF/7Y7fnX/IcsCFd76oPq9kTE12ZxhpdtsjZNCtqjAMi
OaWzOwnnw3EZ5zKsrxS/uh8XPbmlQ2FLfcwMJE8vR22IYuxQ5E6h6BoJ/o5L+Osi
FDjIXJJ/oQzvQ5TDzPvoEtqYu6/fPRvuvqVWy0MB4nR2d8VraqqLqK5rN2tY+pEK
C2Rm4x4fjnF5dz48BwuiTVXqkcIej80GFiyS/uLmykOH7rMFjregOyjjB3ObzH1z
7Q1GEMzJO3kVxsL8qw8doYRU8JGLaNr9l2mYPM+Y+fXTzzIvqw21XU8cQMWHbasD
TjeMir6F9o1ENK8vjPaVvPjlJtenWcmb5WvuBi9uTCGU+H7s6sh1bXOHqX5dY9iB
gz7vqXRySGp+ZmuQZojSghS6MTE6g/5ekdKoVczDK3WpSh6Af8rGZlUqFxpr3U81
SWoU9nu9w7z1ZurgHd4hkVnm63Uxvm0bgufvJN3pBhWKlNMB5bi4eaVDp6g2SFwL
PGn9/gzclqBmyBg5ckPHSC5k8sO+kaJqTidXwUuqhxz2plyH5FWoe+HajMHAj/8n
/xkuwrByvbMwFqcQ3DWr3R3wPBHYOu0/bCyJ60pqI1MqFqZU0mXLdarUI/PvVGVD
fX9JubpddRoA0VuT1hmOAeRJwsPxRzy5Itu/bHOqJPc4QH81BSTc7gJphHijzRWP
02MtMrSYixAY5xWlhVh2dVZwcEptI+sM81+O2Tc9UoRWiSO+5sKLYHbGeFFhatf3
xH+SlNW+u329JM8DXhKsjxQuWA+kzHnbGaFu92Hj302zRAYVfv1Spm6/ant+ZLry
830H/CoU3k6TggXD3Y6T4RiFe578cxPwP6QRhO9m3rjTHcBlK40OEDmuYWxnTxbO
G9PkiJyei+DqkU/kNXCYeH0F1HHfcBbTJQPtcF1h8TKDeW/uvTzcq/zv2wakdwTG
PDwCtqTzL8B2itNwqH5v7Fo3UkYK3EZtB8XKHFpWTkJtbdhxyDhn6MGk+6Ln066q
0YEedcssqeIs1WosXTF5ztxu17/7/LmShIteBw3HsjJOGqPFwX2ctRIMYW22/re+
gJdTrMImschg3V3tl6bjpOeFVMr0af6kMUe0wU3I8cZTOsV2BQrMwVSjfYuQT30y
1xpEHaTjpClBQEwEonuUTCGjORKMds/WMg+9yZHqWlVlgRqgfzx/hE/T4nbfib/P
XVYplL3S0EmqKKgHmNX28yAZHPBgBvTroM3eDh/W8UIUebYs0UYfx/pB7KlQJ/Iz
t+DI7PmOoSmsFrxDDL3DJ6dFQqenRwj7tftfKsvbab5oWezsD4fts+snDLV6cou3
2+bruQbKYdnvSwOo5/hfcYyaGlGMKIC+wX+2uV6rMP+hUGi9SmYWmQufvHTmHQqf
XOmzD5BhNgzj965YpmFUR/nKPvbQvdfKE6WRNac1ubn+06WoA6bt576IpaBlJo/Z
jRCjrlcxpvzYnVTgrMIpgpwUZXrDcibMNAddv/XFDsqnKaJHtEAIAafbz+IxpBZz
We0kneKc53lSBXOMusFAmzqsQS4EeEAjcgPrFhEqxVQ03LpRX7yNR37xPrZUJx0g
NADECULZacOTzhSeeC7tBCgsIKAmJeHPAzC1962X9WFZlLo3TxkyVF2zfOMLPqyo
J/PA1IUosJkAuVnV0USYhbeNWXbSBnzABABtcqYq9P9RdYLcCdAEF1aLgUpX3LKk
EwDfiFvb5pnYPW5WE6guSTD7B/5KWKBMu9lHQMD626QWPhAyv2xg0wHI7OAZptlG
UcFQ/iSMMeBDgstkKcc4H63TB9D3yGHnB4F/yIaXWzaC/1Gzj4AlrWpMiS2zj70J
JYYoRw5Bchht/QNoo0hZDPb+Y5bUYQH3y7k1CJZ1m/fczVTEcEZCkJvlHJr091MG
qI7Bkn0Eniov5jseOC5EQkliphkRgUadFoYxTKTfs5SC1RyzT8eBpoD0YdSeCUUV
R8NbrVCpaaZV77sdUPDgeZTV5qoqLImyBANFWU7/WLCxi4kHHVx9BoHBAxsD5lR2
dX4HSxWCcGBWf24Rg/Y6QZ4HGVwtJPKgOAVzvC1hYRQmxBNDyyfgy84XxEZw0c7j
tqu1ra9egCWT9Ubq6XzSrNy7dndnp8191DORdDw6hBMnUtint4MajLnNLLnbfDKl
Y8g5XpjFW6yIYdZB/joXnW0nMkFkWIJzVUGPaNEbxexPjRwtqkkfxHNWqokdb8K3
qPMXMMXShnOMeQIzDM4XbhrILFyoA3hhww1pZVdC6esyzTYI3nserwLyrkjq0yHv
LUXqkdG80HKF0/2O7xt5aut6Ovek3gERalOPAUo+XcBPSZYGgYwR3hJKb94Sc2VL
VPjNB47hJJ97sRVnoMEZqqfhTHhMfsWZiwezA4K+TaWbBJNdg9R5kpT8NqnwwuIU
obWBfAwlrOE2C5XN+QR7Xng0u4vjjuUNFnQyIH9Dwj0t0Fr98RP1qoQffGmbn/hH
8E/XGoJXE7OqK5eXLoJ2Iq80o1XUcUeVPoHK0O4ddWjjTYRdcyNb0YJki1kA23zo
2yw3TwualUGxuH8REWpONQyNVGgXNIES6j8ziCkgmLdcRFVz/rISoBGF+SB5ZP+6
tyVmRBLqzpEUZ+JTgJZEGCQzQQR2a9p2PH4fgmxQ5zFNPhjSWjpBYESoUNYlJ7QY
tLYWP937uBJ3qg7UAr8fBOQEMWXBBd4yc60WRa7TYnFZ0CetJUL2u5jEIDiPRD7D
gJ1eA9njODcTBUF4JiV9oI50Trb0DVHkoLPpNrt6/xcIhoWqEaaYSOe7EFWFRxF4
iCph/GspaGUkOPPItnb/7cTSudi96Fsd2GfJzJwLuy0Ehd3+uX7SFCD26uRWsSjn
TI4vM1EH197huq2kvYO02Yx3iF54l4VNwlqAzepmRFN4lh7lgcNQg6FT0zEiCOcM
4buA6SP4dGcdG1r7B3S7DOga+dVZQW3o4GKOiOIFpKdJtDMfMwdMochr8xy0YeaQ
9T1n3oXB9eKJOBWp+LSZWKaLP+J6QgX9iXEQv4ACRPimRunavDvlZtKiG7QngTy9
UBmEIwVEGfqfB3zcrwRA1n3Eut2m3fBXleKiEmiEaWTpFbGNUQMCy4CecXYlQRfl
0TYt6ojxbZL0tVyTxF/gfiQeuiCLvIJV80oL1g7h+T8edzldLWqd04o5oYjb7k9q
iK47sOt5xzB8nca7gTfxaJ0DL53I1zemdrte7u0ASqvVeufn2OkoeyVzi7kg9gL8
lLOf1Q9Nqz0K7I9RFrFkXPpP0h7chALaW3nlxXmlLKFaGErFMzZ35aZGUCXMc32r
7BWdqcCV9HDOxpnx32wMo2slMv8EWdP+ENDUOnlw7ipMuu0JWxNrhEGhcSoWWZB9
lUX71islvroTHihLnkAI2h/xgzzhu/VM/GOkKx5pr+uO6OU/Ta2ehykD1+FAGHjj
uobzfqzu3NOrhvV6tOWJzrWtHyColR3Yjjg7r0VMrpqBfUYnPBiePKhLWXM3XOwC
MsHRNsbiB6VyDWaR/ypxqp9pl5fHvK1XB/j38gD2fMXL46YY2vXdu7kDBP+DAder
rKQRZm1BsfHBpWPZU5f8wSVT10xZBvHbN+IMuq0Y6BECUjHlFP1PDhlIALvuxKoL
sAsp7nSKCbLh+ztugYVCE1sCrZJeftMlcCC6pTpuvhBBVJbk63zKx9ojh0yvwo5y
dZ94rvn4B/OzonD3WD9DbQQbkLl4FtR8kVk1kX2i75JCgLS1AuY2LZDuLSA+j0eL
k2+cJOWYEosd098XULVnpMpT3HebhoD55qHz0wi+8+8UHnvvzG+I0WGzYW1CLv+/
sW4XyePC4KVHHwRqQjb/YM/tmSQrkx1B+7Kyu7YQRATUy3zs8vUY4J0ERKRGrBjb
tD0XOWeQSfuZuWtwm0TO/fDKp76FVzQZzeoiK0avWu0YQnYWGGGYwlu0lKrIQ6Hf
ktNvWdpWaU+vQfZ4LxytZmqKofBiHFIVfSvflXrHfjo86H+YOdwZS5L0bYYJBoE7
cjml+ckO6SzOUwp2REr5nB9NdxYTQvtcQjFUu3aZkXLaxDXekbeAF7AXppGHumF2
6VH59Uqi2dpIEQVq46sYQR1xVPst25ExTNf8yDFpPzE9PzDTlBFJ5kA+OzkdP9AV
ENoJVWTSUBlkH/p+HxbwOF33vXj5ARFLz/11dOWrAc2P8gGBAHCH5hPSU4kWxF+v
DxJBTt3AHo8TCXdJC8V9kbH2Xz749sDOaSoDT5u760RKsyVqCNgtRPPEMy1LS7EA
oVu76qxQpiS4WEiG2DbZ7KqnBz+R/9zIS6/CtWDog3y4gWhZlkeA4sVON9f+GdSd
pKjksD3rZ5XDwG1BH3eUwPi7/x0F5P2X6RDrgxUWkjk63HvVrogXWrf6UssVKVPQ
NA6MUgF7QRQJK21CmBLd3+oWkLXlg/M1pvI6yaRs2dGtumeZ/TRZTQIR0GhMgFFQ
U9KLpzchFX3xqwOKv2NjOJgfWD5Kr6yxmt4dRc0EWkQh3bH2MthBNlx2m3XmlqsD
ZsHzRuf+z3okehKH/0SOZtXYYWS7Fb2e392OWhVcGag3VdMtm1EVcol5jBDpwfGF
1tmHt+kT+GGPTVLpybNYIQCH+tXdwDyppjjnsZ2lf862r9j7uLoGagqKMPRYl5Y8
kGs3Dn3zKUh6s9pApDezNMxYtjwjuuVs2QaKK1bZ6bB2UEsIj8C32dFggfevNgre
Rwgenl+7pApwM7OsaJAWYUTLw6tCKD8cEi4XZC4n/rHikU2ZRbqSPFdu8hU7zMVx
K3n8sycX5Q+62hpfh7kH1xWRDBdpeVFKOvElmrrAajottS5i0Mfn3QlTGx8rb6ki
cw4qBe+THGEFInNw8rI+NZXLuLEGaT9a6u8LsfChR7NjVTywPcmP98M/ZcjL8ywm
zR1nd70/luQbktLL3Kf9ypS0r3lEegj7c2TjgPY38unFYIcbHEdWNRAR10sI8caF
JBDK4F/QMdgsEDokrJAlPF7UtyWVDRsTYyT9qAdYFa4Zba0aeCcVlNq2l+mgoivS
3vYrIQ7e6gpf1YE7CCjqNmfpdjs3UxfKEo7N83adaXLVTqDdZ+TBkYex+KXiGh46
nM094HtfNCQr9qLkG2Z25hte7Aj3kU8q6StDwfEr9sO+xynZF2NSpMykaTHU1MbS
3vgP42U6jZ/IwCdLXnc37ItR0sVnVd5WpF9Tij0Eamb0P1Uc/9S6woX3n6UlN6hI
5NTTygAvS6KZZaadYy9cc1HXv+TiJb1rMUyXdZ5/1NsfTtc3UMDi15DNSV109N0Z
WqYtN4XneUYvTMPsvbGd6s36+aM/mPWihfmMz8dAJHywi5Mh1Rpt9xT3ex1eVZ5K
GqyS6ENAYW3G8zNCrxjHHJOxv0jYaoG2AiN9loZr6N9b9+1CoeWOdS1+P+xR/0Cd
oGYHwPnTHbxHln3TV7EsYGMxMeuUpbzCQQVcUdlijqndw4zcbdqIc2jmw0nVPAXJ
8pAaitkRgH5SUtf+Zr47IfipalHY+k5IFCxMONRAL6TsUsmU1jckuliDPkUvjDnU
lyyfWRlvtbLCTxKo5hIwXOIXyOrSzEb5/eWKHtVvqfivAdXE3sXnsb1HQa4GEAQs
aSDMN8OsVRX0jcWYuQWA4W8LIn8skMI/IQJqqkdR64EfIpIViwK25dPzWn3o81gp
GoYIqcy8ZDBPXzU7jN4SaxnE2s5OaLu6OPTwGTcWqE6D37FxrzMaPQqdJUVkVyga
4H26UxDWpLbbSPf0cL32/vUSO0LlLGLQQ3iDOWnUaCpikClp5XDijWOvBSO2Ohlz
Fng+5wP3rVQMABWnATPleEY/1SsPj0n2odJ3MHyuFJUFcFyuL6os6IkOxjl5yXdG
NfIWxkJZ7PsyIfmLr+pSVEttxKrjM281yAjKgXXJ9epQTvHJmK6h/FTEmq6vEJ3N
6/DSioM4QzPZuWmZGUW3D3CDvLx9Z8nWw9pJvfP0CL0bWRJmhYcGGJ9AA4K7NOe1
44M86564XwAHu14wclERKckGJXd3NU2FeTgR4/8BJR9HvRP5uDrOdW/58LW9z+Ov
AVUah57EySBjTLKjCWhodpUz0KwL57417INMK8Th5y5f7X1pQjlq+MUzUhTOBR1h
xxVNLYTEQ/jp2dO3mk2vXjD6HdJ3siV4AYwF93ISkHrmcJMVfhsbLqJyjulpNMUs
i+QujDcYXsSygYn57kBQYau+7HDwcM27OEk0qI20WSL5nc1DR4w8UDHt/JygrJWE
91AT+py1ZbGDkruK1HikqyEqWbwJnApSf43TRCwziIvOCLPT+CtCRJtpaaoWYKz8
/MOJvV8OIBaC12qNPfdgNZEAmHdHF+14KzmScxlML2I73mWroW5uGF9JiUtuwmEA
JOs88B7ezx3hSKd0bMJKHhQoTpK+GNAB13kFZJvZD0ZZ8XJxHmjX6PoAKCiFJCDz
F07MN24UUy44rlJzJZilNkdPVqp80Wi4BDe2KMHYUiaq9M3HSiOVeR4QkAPn+2W2
P22w7zO99N1B47Bn0aPOY8kfI3e09PzZVXuF6Zmo/5i+hHTqj0SpIOcMFGNJVg/w
yaoFZQ5qb+DSlAfpltXsk77NiCyeZE8nUY4YTOoLbNk4KIYFg9JLmq0+hYDh8RD4
et7FRsuy+EHtXKbbqj6ETOpQ0k9owdcNCFx9vr05toIup1IqAe29J73orVI3jy3O
WDNmkbybH1mmbaFW3pO84i1HFj7PpjXMbjeTmpMEgb9zHc2fp9cnybi3u8vlh+d2
wrq+bO/dRpR7FGqPblbordPB1GO6Rszj7L5Z7AhS5PU9LubqaWTuoPYFNJCybbdO
nrf6Qm4lGGRkjUxHPaADDepcNotAbjh32gR5tw070gOZmvaJdgrQNqSPIJ7QXUU3
lDgK9BdsCKqhvOYZaQmKmuzeKjhEGW330gYr88qsqC2TjLxjJYGG2E70LQhHRYaL
TDrPZU5p2Nc7zU2WLcgDm+oHjwO8oQf/a5fh5phIvHN9KzGieL8wbHnGL5f3cJGq
RKH70s85O8RzTCJnnlgcWDm/joLfZP0ejC7EDF6h3PC+XxGRyldfeX1AlzTmJ7lG
6f13H2ri3Cd2g2g1qj7I2zTet60qWjjR5jiqXG5SPd49IX+Bm8Ealh66AdVCzHiI
pDgiPJNT+ojgK99IKw2ZxahZ1C1je7yxvBQYD/pmHWsvP7tz9HvwFpo5ye79xmfJ
ot1tcVkh2FO0mFwvKccxFayCdJhJntKLK5oljcqV8fm2J8aomgKTac7VZcz1wQDe
jlqYf1z/wRB+eN3yvb6MWCB5xvSwZ6ilKX3WJABKWHCpaSNcjHj/lZRUIY3bnPSa
hXcmz/iMCqYKqpv9cGzT/OkZ6LfS+dsFf+fgxba7xJOPin93BQ4Rab+NLfgf1K0J
iNk0e4mD09eUbmQlAO/n/hhAYLBUMNhkvrWaakxIACvsliqtooIHE6PRqpG7ZFcj
JgQM+Z/5FIfWa55W9z20krxPYyf4olt3vfdDEZAaoTSqpjG9mCiepVBLIqWZ0+HC
TEMSyz8dPedOwuiVJN9z7hIqZtMBa00SVqUxm4jl2/k1xcAaItgYrNc+OGuLJdzL
sUCMOnUY0lqhp2cN2qLS+MBPCP4o+C6KET6A8x8LOvrSPsd5LBoVW0sBSQvzPwng
BVdQjLR8ySVGaLZAPndz9ANC5aF9MT3ld7vlr4UHOpGoc4lTdxSzarZXZhae9HIg
fxJQuUcdx7e3A4h0OVdmGgLdn92HYYTvr8ctcw5ma8PDjaouXq4TklWrG6KkpDLo
XrI2ameaRp1mwrZC9VRA0g+yw/M192xey0dvZ5YNdikNOZ2Qp9xsu3pcYplRFC44
wsZk1RCa29vl8hisWQNaCME6XUC8m9oXpYa5xnF/g+pNr9Hozgdyo7kjDoApV+vC
2OptcyG/obxZ+sDkKHC1/WTY4lLEoYDVWVnMV8IyI2DdS247n1jtxRkE7sDrxwv2
LrrXvAscaV4glCRfn50eNCLv4CFByzcIATvWbvBgoWrNP0pdz2aGzcqpOl0Qwva4
wV/v0YaYxf+qGKOxUnUpYjBVHQIBPBoogrqOJ2Qs1BGcRoHkNDlZty0MpswcVkAu
K8/2NMiT7TNd+5lbyMicmaY44v12eb6OWktIKlV9b25MVpUozzKOqDtCIwyyvGWH
gytM/az2/rgLk5Sv+GMFhNOC76N8SS58n6EsiEU0uwcoB43nzXnv9T/WhHypOfvm
5c4kjwng1H2VcvKYHgn4GyD1/KCDKMnTCJtq7dF3W2XKVQ82HY+eDalS9KMRnFG7
wvrL/QyXjZl79d1zBhOiDBr0XbxdMxa7RPotlxyp1Q3DuLPj30CCKiNc6CV9K44J
0TPXKjMtcT+W8sglbQl5JB/3dMLt6v31Yx/jon/0D4jp6xDS2xUWfCsfELKw7vum
XpyUu+MFQFQ41iZZSUy+l2J4ORtsgV/VxtPQaGIIUYRjiLrj0yS1URm6JDFVmMiW
UOOwcoxKAkbehYyo25/BoLX87hXyHwGAxnVAfHjeVUKj4Zt1knYlsO4Yq3OnRing
GdjWn6mYZRGykO5X6fbXBToDgbR7iI8/cJGJRBcZkzCGUeJYSQDe9MtQOx3d8bak
KdLXc8SSxgbPGvkzVCeFtTxOG5RNeleHyAvSKlR7rwMMymEp8wCQLRix2+SDnoMS
GIfmAtYBrP1KJdXPykoUjrrP5izPRdgAAdrDLf/2b+WuJltHS0Kb0SZ6lY2mdIHi
IT+8u6hhPkEIxAjoHENqjiujj6XUQQxRVgBU/6zTuwzPCfUsJmJOnaHIweR9lg3K
aJCDX7lIsf3pRuTxTkl/BK4v4DBlx8CiIacxZsutd7klDlfabLBn0FmMYvWLO3hD
+Kd9dIzJ01fZF/vvJi82FrkUDmuQ8L/4IpAm2GPcFEZDVNxlemwWzEpmqaWKM4xl
3Z6Vv8zFhZ4agFdTS5CW5frfhCGSuG/F8sHNRPIM/01azHdzsk0UHpyoa8pd50C/
WDLqpNc6wQ6uBVZUFstOJkA7CQ8mho/mJMNXhNmXjPAVTrfFgQR41NDIlPQShGlM
IhPgdXfXVfvOTOxJH1DJONOaxNpbCHoz8NjmuNWIWRWu843+aTQx5mQo7JhNqqMu
VkWm8x82Fb7MOIxr8BfOLxuXPdTZVDE+RrDkqCNhldiUNzIThI75SpXQFxL0fV9g
b+2LJblFizbpWpVAaqvJHtdGYsEuvhX8Z7QEINFJDGJVcxT1wMN9ipemxqaquMYg
m6vgTwH6bS7mjalxjLQvkVXQgaAh81J9dB+lHckrhRVTtfQmUoeAyCdnkIZnCssX
zgT7Bz43ajAvtH7CwYf/qL0JRoTEuionNtoPX6J3TYyIYuYyHmwhSIiuILcfwgPv
7Xn+M5WAyqKq61V9951TJgiNta2T1FdvXjMWEdkgVnS7m2a2nF1eaJlcQcyL81RK
9204x/vOoyEfB7HGt067qiAcgswemCBKWgPhOjklf4cM8MRwjcdO4PPTUctMhVnw
I21COMDeKJl8SVTU8pG1MFui2S3tcoO3o1Rr47e0Bffr8ORZNxB24Io6jbzz54HN
PCbjX4qDfCMvW/5pr29M8+cGH15k1h9Cv/QUmFL/TJYweqXTgX4NUaSJqs9WF1ys
MlC7ngkwP2pxW7Wb6ISHC9p7cvP7eT23+stCachOLDbmv6RpFZE5//RQGRSC7w2o
NXkCrwg9jvzpKLZ52m5JnBIeKO/2WQuoVThgLUUX6Dbditb+tnDeC4LgAwV3sQU3
sQvGfzqOsS/j1D+eOgzUj+bGQBYrHOhARxW+WZiCZoyflM18VN3qSZbNpBmVbgXR
OP0+4s0aIkJ4SBKLqQs/LEBwBOdvSmD9hqJYPjLnIU4HywQeodar5XN8dDNLfARO
OTjtnqK48M5ikaDOPAHqj7X9Aka61fHHvDFeYKAx0MSr+8POm/fYi2cvMbi9nkhF
nYDXSeMSCqlNVrXkd2a25ro/kEUJ+xWrfLp5hXmoSQTq2ZtaZEbC3aifDl6Grih7
0OZm0BDnFcOth7TsUWopjBNP9HfC65WdrB4koZ+2Sw+0QljuHOCN+WiGcxkUT3gh
5kGfm4yR4ZVFgF6LnGTGi51hzDBewGY654nPySI3iLGvdaadTVcj1DFVavHAI8kw
QCGWWIOXPi+DHKcOd0kBWuFi2Cmd5jikf3wAYjBJmBkmec95cKbcM3H+IL6RZw6G
Jhz/jNTZtw5K4Tn9BNiwwvldzz3YtBx3wISOitW+0L6K+fX9MYvHttTE462Phpvb
Ol4RRAKiGDxo29vsLxZVtlPBK5TViWy31uA1nEu3IkKj5FJm9k60uyc4qt01bLB2
wmyWCdAdB0ROjk0pSTaR0dyP5gWqRoCURGraIPUQiDxxlIDp/Edde2qxe6AeoJKP
w1/Eceb28Yivw/Yx2XTLNqcn7g361cEZRG3xK30wok7ow/NCCbkWmxJ9WCgsG9xp
XrFrPr4HJ35Jg0QUx9o6aW9nR8HXiUpbMhact3bg7cmJkrK328ccjJM92kZyQ7jV
2+IaipqIudNrp7Qj3kZpP+A/HEIig0EuZlteeeFBlVjStY24VVT4qyHT+3X7SkhD
HM4gkt9YIXpDGatBA8MDqS4SimfyQgZT60kGPWAJDlxtTEU6xKBhvJrcE4AOTb3a
5Ht+YWaeZ2HiQXdynwNQTwf1GSf2+3P4tW2xX23KeGxyNb836G0OVIxs6UNoowYb
2xY9QeLxeom0NZYHHpsjj8SNx3BGulzVFVJxgIgHGHoSALDjuTjLeAje23GXWT35
WhABTVx2J/y7fT6TXN8VGeaBwnJBs0SSciVccf0SryNvEVOQ/BLynPZoJjEg5Ga5
N9NC4iWa7BwcBv83UUCi1uQHHYZYDOTgtdcjPykx4LcSRMnx3aT8zn8I7eBgWkS0
XeMVqGu5fdPPRBD2Fj4vijVvzAf8zcbN83GV6Tft8AcQ1qrkodLYOpQ9bhVEeSc9
8nRNxFcADB9Zr1kf74yLObjnHnlIs9iQbF3KgUGlCNfy9FWm5Bl5i12mmk4ua905
RFZOveCuOL0D1oWOUTRCDzOvj/QRyc3+aCewjd0FEATacrqPyI7CsL4bqXp/gDob
S7bqKzTYg/NcTVyNUxSnwUnOS3lruwNz65F/jeiLbJ3mdr86Yt/BatYj522ab2IQ
4T3QkSuvvR3ksFzcCXxrVZgzDcYebOIx2BbnDTiTtga8hpiXhb3XkowOfNkNSWLh
3k35mQyfUmwt3Xdqo6OF3mu+1z+r68vsnh74gbI9ohl/FoDw9bDFobBehuOGPto7
YipP3oJP4FJfLBea+nRWvAhyUvhwcE2EdkIsxy2ZaD3LvgIShXWwJqeaEEsFTHCJ
WuK6G8E3a07NblheDnZbvYLHO+tYKZqtMQmtEw1wQ4+AAUZPQjzaYgO/nENLBpD3
e0V/YSoqPN5LA2rmD79Qdq8QWMdoxvWoF15t9id9FvkmrrO9xEhiTsHusl+7H5JQ
P0clXnd71OUIac+CNhBDza1qq+2JXxK8iN+8jfWTwb3Q+IpxEXeh1wtDGBqhQ1S3
628Re9P3/mPamp+IT8BH/mlFh9UpfeRPJbyyYMIqJPRbAG3uxpvf13khhZCcJTgs
qr43NWsBRAwv2a0YvYv08zLHUIvpPMrer6aU9f6fm2tN9rPHtGcPahdSU7yX4L4s
MM+7QSXiaoyiGqzFOnECvkPOM6TTvmi894ctZwPeA5+ktPSdDzmOtMWlqhVUv3lv
oKuh+GcVFFMVOA1iD3+R4Dqq6FMMtr2dZY00dNEcKCw/WHIKPOIJoxugsm9QQexr
lbfqw+JQc/FB7oROQc6ErmtRe28NhoL+xrDwYBb0YkcAbUr04AKZltzOLtybtJsH
1NHAGs3GJ8HOvE4yxntJHyC3Qe2q/HQuL+FRfmrWvHQfaQdCeuMGmpFBC8R/qtO+
78xVbdl9L86zky911KOAD1n2AgDj6A1zl6AqZV03S8WlZx+n7x26mywnfjqkehhO
y/3MrZG7ALVfknsNAn11iBO1H9zALtJh8d3vI9moaHj87AZIXeUIAt1xIr0aHrMk
GTt0TtgX6Okx9ryImeWa08o2dM/Jkl7uxBZ1BCgnJ4uRe+fOG0jBu6aysybISoB0
vjwvMmFMRxZJHeFAituQB1eE8xbAvLKzvL0BPMyZ3TLsctnGkr3pxBweijZOa5SR
CWPgzcbG2S0INt4ZrC6imhUHdQETz4C7gKBiQoZnd4DtQUxr1UmD8DQKJrql4BNE
A4DAGQp6gS0c7jI4KWTaL0AkIYAQAPtURMrOVmuJDUyrjgSBSOSVdA1Tx/GWoqqZ
K1lIjGqYYEc6enx/JR4a8kJsfVumyzGdQnxqbYqGy4aODG7R2SyIh/GEvntsyIsP
LdtIkFuTasJgQNlUFZNaFE/wZx0HaPJAMOTid9HbNJk/s6JQxqdDCSwXXmDJCRUQ
hVxXmEXvjqWjhcKzXs09IZ3CMgF6BGM8wIsx8PfmKI15N7emu8pwzG9akEqLDGqu
hmGQf9nUxmZ4RGF17CdQZvNq4d7ktHEzsMLdzOyMnoOTce43uZ0Y+vRPht4y8Q1c
tTbsPQp1T/Q9lHxVEvwl/H8LJdtnd/HTcMxHY+JNM+R9yVAfXeywwMIVQi8WMsBY
3OsArrsBb2jHIoR7XOAN6BHHPQ9ngvldJrfEjqMSSDhjldJKl3yBY9YGMg/Nqant
aekF2nDnL8eZWNO+q5t6cTS4g/bFTqBJAvjELQgozMo3GBQ7Z38NG+oj1WIbGGQc
CwmQcNVNlnUKcnxwDkmcuE6cHV+qlruFI+10SqI/dJ61tOO0HC+wgsh5zYxVL4Yr
A+ZJE7ao2cDubuYV2kCmmaLbRBs5cN5nRMxwYBikazI/OGKERpP15NKuVOq2F6QP
WgmdT1oH93Qazsu9nwDMkrn84rIj3ZBv7PJV53mDl+oA4JqthIPNsLlwRHkTK/Er
tUmfHw+mpKgSWbxwlowYR5OeIUjJtnweVcazE6knCfchDWMyyu//vzADgd5sl+RC
42eWy1PLPLUFfsAu4+h6wciBQaKIHcPRx9IB3jhzYyqovbhLTOlF9hA70tvrhPUg
iqZMc9rCOmBbEIl0gsjdLKYCvrogFLM+LzxCBd4dGlT1wdXB8p1uHNEZUS1TuRv4
nbyxSpOLd7o5QSTvGihKDnp+TQCAh1MUCBHMlgwRbhCoqrAkpaxggY5GO2iTKFec
tafL9S5RxrX2EuK7FljZ8eJvc0NE5xlM9+BYd5xWeslolCgrTVwUT/jJt1RLmdLU
EXDGn1/mQHCEocFhD1XPPC6f8+GtrBTKCOtleOev0565HZD+4/QR8Ksuo6PZb0is
awcCNiVK4rOWlKIvJJ4Hi1t58HyLClfO59qQQS7TPc9TRobgBdVfAZE8Oe9qphGn
9ccCFomhaC6+plUDJ4wulM1nYoBryv4h+WkWSyEZI3AN2dIPeAMPfpw56cacPaEr
e6trA+75WD/GO3ZWv7aseeVfpyaVHcY/656GnmKWDF7RLBIOcsfxM+YpVYL+m4Tp
Dg5tmTV6i+GF8kAVBdmozgEe2lc8ak7wOvPbeShuegLLZj2mdgdop+pEqjmXkHDQ
bJ4wJLdKNkS2BMlegfLN0qCjU3Yvl0GCdl1x5fnIA+ZYTl5yhIg4vO9DPoX05cje
m5mzDNdjjUdji8/l0di0DYrwD59HKIO8nBI/UDO80JWmyadh2lkv46z3T3XWh5RE
nsXu/0g54tlnCKjiQ4UT+gK1fb9lmmF4BLecLYy9eusJLSJVX1WnxCi8lBWpobDC
7bPpkU78X5N/cS0b9M1n2ubrTEih3/Y+gZWhMe9MZqGohV1nKH8iCpjgpv3E1+uT
5ZA8TEsA0jkP7/tLE+78WPAhKXVoiM2lOu0+h2DHVY4Oh9EwJ2/tRATYtMyIK2Ts
d45874sYFDnzZaaIbY/PbF1lFa4UpZSvARx+vVKwS7ad6H9PNdIYoXaw3XThRnjv
XjtSxev14cALRYb+0bVwLBOOlhSxvNxwIq3GVNy7ZILQ3ROTYPqmCLzIHt1Sn39/
GADsJHDAmhS4eXiuXKvqKYW56e9adOC8W7AU4Ah3pzYYGBtaDOQv7iQIXWJeeAey
OtkMxIfvgaJmjWEwqAWjj1IdvvYPjDh7aWHhBOO1j2VXMQmEN8RjfuTdTQG+WYQV
gYaN4UQ6ocEcSEdTv3FQ2FYy2B6lVzPDW5iySkBLXRqrZDeZ3pb9PJywAEcCUEl/
tV+i1+BoLBafF9QHY2vJ0TOyRJXR1bbCQzJcTcRCC7C9uYdqTV+omS3/6TcI9kCz
HaBhwkArztSrBjCXnmvaD36nWF/s+ElJrb9eZG2SmHyEL1+ABIi2hWdKJftoSRep
kuFf9ytBjIfbg+sWcYeA3iACnlbdch14XGKr6TlJMUbWXT8wWY0+EAltWiIdkNkR
C5YKNQv2EF6tUm8lkmqXk8NMeyEasX+PILr3b3pd2xrYsKU07AOVT2k7jta7h7CV
e+prexln9UeKFHHRg3/KYz6tiZAHMQ28uPuV2sN4niEKcc1w9qBFCuCgB3AAme3e
AlGYtvHigLUYJpsQS7PbSOFSYe4o/QbtQi+ae55vTzQzLr5MtMa4doLm4MwGpQM4
kWrWxQAYAEwi7s7aLkPgsT9hPUSLKMIUzYyH2xPPyx0JSTW8reWl0vI3BOBQmyV4
0LtFNIIChU9uTifJK4XGHaDDWIgYiZIQtDniOBkA2wc6AwvllXaOAXsYOUemGZTx
4Akxnh7AT/Pzdso040/pWQmwe0RzoDrmKCL42wC0cpyZTAg+mD1O3vi2Z0I9BYS/
ZverNxbyBMy1ovQeUNSP/bgLHWv2UIaQZzxpAsGI/iqENbRmcURPP9t/r+Lhx7Mi
BH4YIH07Xb3IndjstMTFAYl5bR66ajCsGDGkfF37KQPGmc8k2w1hI6Iz2KPuNP92
0dWy/iSgV+Jmx+UJ35zHlPng9OGkgSAh9tpRQksG+JvZRsXa9454mA/F9/aOWaVG
AeQhAYbpw23bb9iD0qeJCdueH7OUQc+e6XpaYNlEDpUwbavnmuehkxn3b+oN/BRM
hGFkdZs7fh2+SJGsjVH/BFnX59pE61QMtKilBi4hDV7gcHl6ZSS7Hvx0jp8vcU9z
ON8iWZnvIlbsV6xqqbp42oQjDmDrLw1pMgeOMg5yo5BWtt/+nR1lJTyAkYM6fjRP
f4v2AlLJ1FKq2FWzUAfeLxlIAelqsMfolEb+BjUw4W6RilgTyxPCQhQQ3BvOmUus
pBtk1pJtsYP3MMYU2oJM03zeMZed1ZeMmYwXE2OTT9GvanW11VZ0g9fdvsqDGw/F
SRHVOwJ5O1kRyNpay3b5m33QBuNnbnF/fG2t4YkDNMvtKGow81mafm8y3LHeaDt0
1f0hxh0EwGLlRKIuNIOMLTKpc2ma7knj2zFdi7I2wJ9GRG1xDgCTqjRqsMyTRBpZ
T+H7PdTwbM5T4bgfr36GPRkpfWh1LzOxAoLe8mhwOfdTWISRio45cgHujxcDlwU6
1UmmRwAO8zVPsyLZN3xw5/HHiLqxaFeyTuGKSmBG+bsOqm3JfzRBCmw/nqDhMNH6
a0d5zLpifiEmgM85DDVI82rxdwrFCkpm5yctOwwxX9IqS7jRLMclWWqyELerwQ6Z
MflWrwZLNynEKD8QHJLS0cQqijnO5ZIGxGIDPVP4GZLRqftY6ZjzzlXiAaweQH03
Ga5uvLYepQzpwrP4zsvP6lHq9KEdsozOTrIcYKPi/eQTDpBBHbyxz/QUwEQkTCru
nV/SvD66JhzNmMaP9GsjsfCU1/+KhfUJ0tLm8w2ov4VSHi/FS/+SbYg338TsC6LL
Gm9GQDmjG+9F/IyqsX/4fRSqxmN40NAFOJtnr+5G2ExwgsQqJdRiSEcX5UPQ6EMy
nkmdi2JemcYlpwWlXDQGFhPYVGsTMwPFKFOTknYJQRWqh0/eLZdqNWkybQXbKSKV
rGWc4uUIz9ftvvI+vPg5IRhgr0Wpo4ZZ3U9XCZj1ORuqIXz1rH5x4tclu2rDKf4P
+pthRQTa4JshArYJMYj8Fwi9LjXXX/VDT94EDZchOSivAskqbSOFYbcwQdJgpfvz
ghn2CPOBbiYIQwmD89HfkSpugH/+B2+AcOcgbWgNC7TlhmWiBGZRtE+rImVt1t8a
k+XutjC1/LNI27VU6k2EdHRVjS5dSto+X9g74gwdXtKCb6GSZFJ9idnk4C6hDg8h
+72mUbdYSRr2nSSUjPhbJCjt9AsUSoARxXnKkYvb0PfwdHk/kjH34JNm+oWkIbmp
qUaEGGrjyAXfNAu5JmiU24trMSfc+3nzyEmkS/rFHcEexwAkq/6VuVyfr+DGbnJP
J0OmG2mlIMs+cEdmUYs2zMtp3JgWCEfL1C3hJLx8HQombwORSLHO9BA3oMnsUX2Q
WQ0vXC91DZoVyJ4Ja1zgGisj8Me3v9vvEnvmrNeiayl24Rp5nAe17fqhLdFXKNjB
8uKEV/i9eWqcijQHcu4gA+3IuigeLLs6c6FMR2wYqTRIe6X8auZR4PNdaub1WjRG
6gQnnuJwVOc+olKFe4+S1ySczZwTthboRuu777awG9sZbBZfSp9s3H+qpkauSFPX
dyAYJ3jcMhZFk4OClIwwzcr/Ef96QXbGDWdvULAMpACRznMtz7aAOVwUELOweteV
Vo5WsGIMeNfE70zaMeQD9ZpFWSNtGi2MB9AqM1sL2WZvWfAoBE3/hoMVLmWY6wKv
KQQowrA5OI9LfcOAsxUW2V+D3QKHB36cEyfmxCG/9aZ/2Ad9sBHRiMRqct6I62UP
NHbbv14jN3G+7rCHQxPjHRKKGuboq+vX0FazS/KKy9hOFZYvtGwkS/cp5XvHrMiO
OEdVYfUCEk9aXL4UWqTb9sHklnO0X9dLeOGl8qYeQBf2EfBO2nvITMTj0iPWHyHN
C/4zawksqYtLjmXNhudn65X5xDQURD14iQqj5IOumiadjrfM7EUGWbGAU8Z+l357
LRq/EbxJeHNShJCpaDecdLfyvGX34KUsRBGZX3dWKOoERS5H0Biw8i3JFj5Qnmv2
gpTvT4LH3b47iNN6RmqAYGeiosErSDsqEClyMWhokiT8FdQW5+3yV/ppNvI85h4x
wY2qrGGRzNqmvh415f6r21zyzohNH+eJQYs/xvELLuJ9klN14hIvgs7Nidyh25YT
FbqI3cFPepafGoXQBaXVTXpsk8XHw6dx/kGb4tH2Q5cZzNT84VkGSzg44Yvz7EhB
XfW0y+o9SCC1tv5gQh9nxrDNBOkAWzgjtix0SA/nGYmI6ZgI9jNSPx3upsEAj371
7MsccjIs5ChX7TP0GwRxGEdzH8bFcEDoEShDfPTa5l7SGy1n5XzqZkkTKhYq7Tya
2yvDOwqV8hPk5HplD1w91fme4+51qmY69ooJhFSsN1ZWLE3gfHTHhKe7xpNqjrFg
kh/env5EiUiZwFd85HFEqO+Z/+LFNper9pmy0s/JsofNWQN24vt6/uRn2nMP/W8E
a1hNNusxRmhuCxa7nw74sKx9wzpal5zgRqwGIhS3L1+Gf4qwEwwsOSTWeC81yh/E
/HkCwaBleGDvNY7W/vYJ5hd5/VSDUSAb+Y9MvDUp9kaoTEkQKUDmR/W3IVPqTdsk
GT8ep3Y9410JRx+NO873cuz4e7NC+svRCUad/xMPrlz6DSxrkjHiOR4K5OoAlo3O
8l3sjptcIq9/IZTHB8SZMfO6vL0MCVgUx5Q9NInOlgHSrEg8FVbkjuVjh91l5sHC
TSZeoy72HBRY9ZxTwUEH1njoOPnz2hg49BcqgrkLh4U7UGtvwmWkMC9kckxyRBe+
4XNbZJkSGAmdcr8shn5MmfupmCG071T0skl+WsWohqg2CCiEkWIsZL8vgmHvPN8M
dwitkgWfW8UjdAnbnTyeIaFa8Bat914trsjBbk/hr8Vi1fxBsQW6cr5o16VDZsfT
GclcUSD8jwHhfj0iudIPx8biUtwL+Wz9bYthVigJc8JfQdoRgUaZCnPt8wXIVnKA
NnvjbjH3FU06LTjNcXFhqcS5gzldPl4lFCDUu/dPIfsf9eS21l7lbNpqeueGF/ur
WzSQ9uHS5LwcuEyFbuxOwGK20XeaErI1qslHZM5qaANbd6F41odojud0YXAUgs8z
hnJTCKgO1wLkBst9ngo5IKDfAAmweNGMBE6MGzW7My7WKugzacs4NnMulqByx+hC
UcbySB3c9IpnoreK5SNnpKX35DsWpSk+SFqsnURSWxYkCbRAJWQUcIzBg891u5Wo
MUjDYDwa2iR6HBO/EUSEEtMLAj54anF4e6BH/xa9zatgZqMPzsmpi4nA4tXF4uX4
YgVq2yduqwA/JUiD94m31k5FLgTNKGQh1cyrcqUpYxhqzDx0oNsZpqt6GDsYr+zf
NOdnCLPlcVhasuecpKbFtp3kNBOGS6D7SA5gvIjlJowuGVyOqW2T7YOe5rmyusC8
0tXQU5xZv+4iVmCHhJSzfj2RPXm+w5x8cSXDf4d2cMpb5r92ezdHo7nXaC5f8fTI
tMAo4e+M0eForKxjMz5Zh7rUXPWw5x052syiz01jKycKhrytCO97KL+J/1twjstA
9N8Y1osWMgDdBpBrlQEfPnpufnZmv7LELZMXRpUOVdAbQ/ImRafzyCQj5xkfmzzW
auExHnmv0H7jkWlmTxJuuBmo52g7xg37MZgtFDKeQPiGcvgS3oJExj8Ii6vsDy/o
HznAJG5VwslcPVZ0GuJYyLf1rG4YMQ3zmN7CLXcxIv6dLKvlGgKh2+5NLHbK4vrf
J2NrXzKgNtMAXYeNHl65pl1VHnIQSiuBVboLNULmzSfUbzchyf+FEYJDs+30/ul+
b0AHikK7IP7iyhHZWRDFXrkmLMd8b4gv76NWqHcLuLCH9joP2b9nhgbDN3vATi6t
nTIG2FV6YmeQcDTEm7tNmMJj0p9wppNy2KcCzH1xStG0O/4Y9MfiyVhVuIy4SAJC
+a3UBmRU+3/DbpVuqpwySnsHBAsNbidN6yTrD1fQyV4j9nPnGe+7Op/yoXmzaMuR
bCPYjntOoP0cw3aPfHYSX1zp8kCiZizdTCGpem9YTd2s2vELssKHiSfsnzy2hVWT
3eteWw6AwcxbP/SZDQlQ+ILZXY/5ydMlIHIATO8qUnZVWzT5iH98z6jsZJ6mPUuP
uiO6ckQcQaNtFb4576ZAU2/cILIOJjeUpsskBekwdZ++uI0gR13U0dHTc7kjAHZY
lY6D4+VPqsFp60jSmzz9g8BcohpH7KE26U5j1EUq2bg1a4WG/pp9OgKq3pBjhpKp
ojFk0fF3jpHW/AcnzvkzdD4AEhsc08IutEEFNA0lkKlDcCcY9hlqX8vdfd4Au7s1
kG0zEBoQ2FDJCHZHgINWWnJJKKs3vNnNXw17+uVO1GtFliW3JCogoWLhy1RI880Q
s7XpuTk4Jc/foTzV8MZClrdKygQNj1V5aD8N1MSeAsr7ekMLhwL1IE37jfdGXeD0
LQ/PIx5/DAAfD0eLk5IiHbILNt0PnHcGrp+EYI07eEQmaKpQLGcjsEpUNuEbRFUQ
0DZzDryUob57MN3Yg4j+G0Fri6aaScwcHTQ7ESlyHdVArEgaGLT+R64O5n6h0kig
IvO9LizsCGj98bVEbqjuZ4No+v095D8ca8N22bVC10QsdxRiNiIV+qPRAPHY+EWK
2vTIqL+2mB7yGQvbh5WD4kggH3fqz4akOlRW4+WJBmqVAJo/AtAKQa+hxADNeOHh
ZRrLfxOxnFfzvNbDhbljptZhU4L8UWdvTwN92KOlbq23y2ZgH6g+y9qxSGmSfhAz
fAd6YsG2J6AVoqRNtVy/mn0mt+5/T4250tHOq9ZjJZCvwFs/3H3AXvcYgULcZd79
Ug44DLdDkejetV6PV/EEunyRVL2+gUDFdg2XBLy4qETRn/CJKFinY142XI0Bulzz
WrctJlmQ7Lqj4cyruKcmU7mh6vkggZdJ+J/24s3yfR6YQIHG9WkmCLXpGW94cxML
pIPDi6soQnUipWKlGQKQCgk/b9gwUx3Xw7FnwLk0qi44dCfO5BssTVJS0ooyAGvi
RlPGiogy716SjPpC5DBXY7O1fi5HoK72QLOjRmjfAVV2wG4dpSQQNQVxegObPRSi
nkT7ZUVbOz+NcwFq3TuiVDIRa6q2z1JpUfN6MoYsrmAA7VqdEZrLej1QuuERlaW8
oD7lBPB6A7aNYhWgx/vfofxFLyL8uWPs7zl9MD6zAqONreXgq76CUNZcHKGeaViJ
YcQU/qdSxD9QMWtBgBCnestRqs9azPSWki0Z9hcL8oYNoxi1gYdahyadPZ7t/Tev
fg5L0caqkvSUSFByqrp3MERi9/9+VKpVSe6XtdUvrpYCLdhOKSA4KyToWH9lxLm5
KmBX1a4jovQpYcFh71hjedB5YjY+6CpLZnYHhcmaX2Ijs119GQLdvHjUCa0L+0hd
nsc7RgNV8dtSHzPNTPY2ea3apPIkOahT3xK37xA2wBvQf0uzc1jABNRUkJsRle9i
ZKh40KxMU+aV3e9DpSaifW4jdKUOmMREIgM6vLRO/6BFzQXLNnlHxc0EM5uZEhzT
rkSi/DhTPH99N72qOrUjrNUwX5s3qZQ1gDGW1s4b9xs+v7qYMVQVQp33EHLrOw9f
BDU2baQ+Dl5ctVoThsw7v8eRNl+gUR6qBY/peIJNdqRzYmEOnRQBHuyqd4kpwVKv
7Z/5vOMcegJRFZJ/wk9F0iPpchYjlVWZMHzdiZ+oEaunSLjMm3/75+ij7RpKF2Wi
iBpwMmtY0Inh75hsCYQsBBXUk+Sd6MJSaF64FdvbMTl98CZuCpRaVgnVUUc9IIgC
KD5SjJZ+5PDVDp6Nk0AGxM3xtFRIk5B4BcnIxfqLPzeOz1B3hK3XGwCjJp1nI4Rh
2TtpGUhYXWL5XLyNPKx1B8BhM9cnfDKfaK62Sr0n8KS07Ei2T4vBVxmbryMvEgoB
CrDxUgeMDNsPf8QPNW6WXaCftMBGNspstTnh62s0DeSnjJpVWSqHBcyjHB0Mg9Ry
qivX6pJNbFq1neAEe4/a+7cPtetKvb3hAok1PRLgiiNQIGx5lFVwLxqjUYeimgeC
ynON5yCAyzmtACIc0iIHP93JXUTm7GHehx9A9mLDyZn2aLSxZ/bSJT+DvZx/bm+j
uoNhcW5c8cuI3iVik2bt0ZiBvBU8V070L6Loyt2pbKCoO4FFaaVPyNKQEhugE782
7qv6JZHMBsQiX989FjLU0I9G2OP9FF6tUx9CeN+n/IBSQ6mhSSNTuHJ4PZpIlsKT
PF1qZhGyaOGH+ha/BV5el9DE3qi7NoWjEcMhKJ/aFaY5PqkICUPDSVK/Xx+btJPp
5kGqnXWyeFYUj11HZaKx3dzoh6oWN9EaUDaNmGOcO2DpPeE9pSa2r+ZIYaSfoWhX
Svt1F1vTzSSho12bnamLjFTDhk+nIl8QX5e4RHMQAAYrykOzGMTQJO09Q6fj0guQ
s+3aXHlCt84i/GiOLk+Li57J8zzThMs54zwG/ui0E8urkr8tZSTkEAYYmLFFxQ0S
yMPwuvAjwX0NTZCir3sBCRciy1hIoAN6Ip2F6upuGPbr4tgCoQ+CfPM1u43V5QmW
C/EeamQHRL88tYxkxMfVO0L37YnoEZ5SctuYlfPGWaGt15pcHRqXbetuuLWnhOVX
3lQQW1m67AlrngMyK4liuQ9+vk64Ac0MBhTxRkN0lWTtsjcW+Q7zitUBFT983BI/
cJEycPfny/vl0jWf2YprpH8GSNNzJZVr+eOmJMUKoAv0ijjMH8Z8Y1eCa7jPBc/r
wJly/tca+AUAQwZUmqxHHZ6sGpX9Cgaf8gZTRtZckQZS6GJuimsibbFYs7FVtrpN
JfKkFifNFD/oj0wZgWtiqFIidfoKo/UFyF8Ms9PVRg7n/aoPmrHoCJNx7Ju6YQGG
PTbK9On5M5sjT4CSJJQrizDtozb7ZWZyuOihsNEMWb/Y97+eMRd4RSnX6AqKiuzQ
HGP5KdA/+/myDGIv2Pcn7GLopMEWX+nrY9OiUm5nVKqNdNrkAjAmUpcDy0VK5N20
YVuh+LY1Nan4+peCV2eYoWG87JL58evzMTzEwDeQmZiFqKEAmzymT8Hg9Hmt0lyY
udPl6J08HT0eg3dT7CILoE8VH9/z7d0C4+3aYut1hCarN9Dt35tlE41ID1FPl/ta
6TvA7PxKsjeK23fvTxiIIhK4UAsKIo68yNtALVkw4M7rUPMBQtft+ZXAXjKjrPXK
IFyV6eoUXqBxhsMIHaaxKHMlOgvzCJtpGlOmdlCC7qc1I8rukUrxGLlkDI9TR5Df
S69dN21uw+pa55a1YZ+bHf8ftWu18sCCB7SOQRqQA7BnC0VP0PcNjRyUepLkC4s/
Cg8TOZ67IRofNIhWUH9+ygnUDX90oDO3HVo7h7hAiiiiAEYtd4tyehBMAd/aV2Bj
6Ba9RxNIQ7pCn3ckJBvqnW9B/9cXCUwRhrrPZi7ZRxgOnZt+qRjgHxofa4kiWkly
c/Rko4/RxZ26EKKWZXdmJTA251cRapr8FiVd5tqG9nrtrNisGlin+pjvLBCBPPJm
aognhVB1L+UlQCr6+NULPT85Kn+YFw5bNq77fREz7jg16bQNWXlqW44IMdLX1lXO
605h3jQfYwsp6YWLMBBjMUzcF6plyduHL/km05EDZYz8xRg9JurwxTxVjjQseKDS
bI7G1N6M+id3ILqQsdpdDr8dGdw7Bo5dV9ozr4VNh5ainic05p0BwkjQLi+3Xkjc
9EO2vshqc1bTQwiLGjJoPv1d5a3Q5jygi6PG5FiuRuqiSHPJUDYfD3rFnHzs1KS6
tCbBp9j9s95kteCtAsv8qc6E0xXouiBWHri0fXzTXlgQbysTl1njViSug6FKjA1L
68i9zy0HMBxT198pRjjvixxg6GCX78WYjwKigSSBRx8Cju1jQNJ0zwpSGszHMs6U
mWGFFFbu3/KLh8Q1ETIpGTWMA3++TcLnsz+Q+duHrViZSZoYZCeaY56sU0fSXYE7
cH4lnB3zhsi6nHRbfZXqINYrJwJ0Qx3/PmlQMorL0gNRXYcL8ZTTB4gmb1+7d4qb
PVJmtUuwoMj/dF5HDat0zG7DGesox/PyTPMlCObgi01V7B+sjaQPeG30AOeHRLNv
lzufWxC3mOb9UQWSF7yC1Z55M4+fia8bWbnNuru/iMtgt/ewjpJU++RYUQLKw6RZ
TJxoeKqdpQDcVNStuOV/iyj1Lb/8FQP3/AZ5WfxP6Z0mT1M2DYbX2BceFxARruOr
X+2rdl3II6ELqV1STUniFeG8GRouBVm2P25E0GkjHLDp5UHzxK30v3KiZb+LbpmU
I9Bw6ewZX8mmocKRI+8jzGjgmBhoSW8k7WxVXeN8G3H8ox2XRcI81mXKkmhJCb+k
J2MAPppnh/+BJ6twtCyPBdnlXoXMDq0AhLkTlCD0F7NJcgYT1PPUXjTEPlkWnVg9
YKMFO4YIiUremlzR766G3nKIAYaeT2d1SZatJ8nClPkatp6SZaJ1eUcljO0sMoR0
nbFN76oLhdwJtklzOJ8kW43MEmw3trP5riyfTKeJFHcCex1kqYHop9id0DFFAG9t
yaRoRq/X3gUNSkpU57x3oq5/nbsF4wi3U1/XjKKxNtvr1/ucnYqI1AfCs3J44cgq
eWSIf8frk8AI2QEXHKuQYFPEikLBNX+GrQvjb/Q6Z/bpB5JFdm0hienzn9UT1uAA
aXKjxzuopabLVehqYesF79FhCtHssLsG7yK43dKYq8GpsK/L6l5K1Y+CLkp3cPB9
QvIwWliHwkZT7kNT+vv3CvW6wO2cxo3eEngLVAxvH+4Z49d/oy4dexCguNcS4Xsf
iwsv8bHnXK+tUSow6K3s2eBtmOHCxwyyPRAGV3zyoogV+y8Fy45WzzO25Tg5TxNY
4+mNZn7ImbvUOcqurRdZo7KhxhB5uuI7/YZdeN+f2Bv1HQ/2Rm5YCM1Hf9+qqk8f
Fo//0E06pZPY6PiohXngy6PJEzK3+yKUyMT4MAVPNVP7NUqjYNODOZzoOZjH0SwI
4QTtA53g20RLxgA4piG0Pe0RrYz4ds856fafVKuXEhtxFRNcCiX8r2oJOHQxJWAY
x/Of/xOaGdb1k/l2GMVCQy9sVQxRVztmEyUPyhUsinlxjMqT0PHunqeiy6vgt9dj
FOXagv+EBWQIp4xVxDOSUEoctPs4kMOY81HOSXBazEmWLOqpwteIdX8n9/NlEmun
+mdGB1yHsQl1J2nlnh+vqgq1efJTTQgGMkYVtqhzRYRa+Rg5YrWz+TpqrVhDjCxB
edcs0zRdRxn7FvZQWbK8EBK+iZ2TR8DMWFTeTlV64GhNXJnC/kHJRxZrPqPSY255
YvCIXNmmD2h/vFjzLaSm6UXDgZncvaI0uFU3ZTspSw65E9KXYISVkCSKgWr6dpA7
04xtFEga903r34l2Yu2IrRpVaHgMbPpNPfzxeyI2b+Z9qnFZ/HTqca44qWNPnHPe
hy1ahcKsP2E3AsdHr+gQwi1kq8KiCFJftK5vaowY0KjjWB3+pAjRgnvPKlRWvdVs
IfYZVC4kSBHIQ8iQXDIuqmGfFVilTyN0tI07d1frYsF5fpf/XI9z+t9JsCzKl4fV
TVE1QJBFa0N8AqaRSkWfn6u3nr4VztNi2kpx7D7SL6PmQn9QHpZyGQzbs78RuImG
hiCnBVnzcnhELHj4DkxAUys3eaRpHJhKrC3fLS6UQaaAZIoIbl/xwRbMMShyyyqk
zLAZ2VB7LaHiPsp3dkA/ioNV2r7+Kq6VIpEwIIz9Qd97YVsTkpWONYuXVIDcWTg6
Vz4byUG7NuQccxJw8qbQ0FkJszg6CR+5G75Eg0YNkDRua3SbuK+FqdIJWeuW87PB
OEEMeIoHW0u9lmvNOzF+O/ooEd67455EXEi0gAkyO2iecSA4P9pV9Bt1k5pmyNNI
0OODTywmDdJLxj9QkFCYYiteSmKO4Pj5lEqwTaIb6m+zOQxDXn8v01J82eTnI8Pg
FUpjmCVw3mua69uT703HJnVGmX8bCxby22lhYShPY8+y985GlpcTUf8iA/+btCSb
bUwcRdn13MW0fI4N/81AxSDfTe2w+GYRmIlk5kEGudoZT9qPukH6ECmOtbKNlNAg
dnG9n0PneTDDcCWYkKoJ4os8b1BauX5oiUTJc+VQsjs70ZyjW5XmlCk8bmGZoW3J
IbAOe75mss1hU3+AZahRIfMqAR7cl8SlSP9GUBdly/P8y55urRBk9v0eaFp24IJL
38AVKR5y27V2ys42i0BEiZ8KyFKJQ5zdo1tgaboR9vYWAZoFph6HdHK29FyPJqSY
cSxaVh9NViSojIQYU/JJ//toStxt7yB2g8lYx1nTatk55YCi6jESFcjLL2z0RM+t
6r6jSf3/IBzgJi2Ze3kzJA4qTkeuifC8cQnflTlg3Sw4hsauk8M6dxVfq62RTJi0
9VdL+zm/EaoduKMyniRjgW9B1W01FhS20IUwfzUwL+Z1gOSaDG8iULtBg+LT5LGb
fVK2nigsapCNYTa7isDuCVC9s9L+XHoA3AfiwEvd8HVVMgpniJhT8ZgWryoJSUUZ
lS8+6+gYOl0PUfaS+Xz6PDIFngHNF7xp2oV1/cdF2cK0geIJyW+vAap9VClh4BQC
vYh5IdsxwlhCGZ+Tq8odNjMXyYpWSeNFLoYtOpXW1Ugmlq47ITlm9ioBon2+gkLA
dsGMB4vN8FXppfrzrm4bq722mGJVRwFAJhvh+bEG2jdqmI+v6qpH3HjXzc/QWlpT
7JBvDgqrXS+oHgNcN59FdbjCBU/xpMCrWhI0iJBQFXXXZU2hP4ACqPfrv4m6qlVi
b5yuhxFLJP7T+9FrtfjHD0MlMCgOcrQe592TJFcTrrEXPkQulP9AC9icluhu9d3R
gHpfQX7tI41LK1WKNPReYdzPJIyWUDLMy/par1OuZJ4Y735sBDWHK/84APFFkdII
7SzOB0bK76BRTKjTLUsK23OHqOH/bdb7xa418JlKYVCy9uR8LOxhtsow+3vmWgo4
JhxOYZcd3g6dfVBzZBEl4IdcBvBgW9XkJ0zX8nMf6+X1RCdO4eCwDhECdHj5QmYU
90AO9FqGOTcXxi/Em+kC9HNmGYy2LwexECRn555XwDA3vrQEICEIPmfz67dsTwJB
INU3bQX31pat7w40LUwuCSUIMMNwUZ/uox0rhcKgDQH6oMUSramSQLApaOxJjbUW
cqKfQiZ/glI40h8A+HJ+bSyGYD10/ztHGna3XL9N82I+JP5y4wIKrki1GtxXjULG
JP6wtj4yh7NhOi4Wt0SMYc0rkrpDuWv8AtAfe60tDuWGIaVXE2cKLuVU6kk2tfjr
gdE2Q/B/SnicqCi4nTq4ZMQoTMmhdLOKE5Cf9bhds8rX+jITQOTLn8UC5wYUano8
3CnhF2wubk8S2bWZbvyJnylyytLjyrenz4Sq4HXR01aH1ppyQis+W0h52uI2HyzV
2nXLNjrg93a6R2CDCAV7zNFjfeJmpOUky1CK2le8HZ6GUrlohACC0Mho/gEUW4iJ
8n8XClHSY9v6YQbQ7juSANwg6l98IlITfcx156c+yBdXBLS+VSdYZreUEpv+s4SY
wqLNMoQBxJHt/NCTUYvjytDOQ0muRIksqMn/21kj+Ha9cEBNXiiBgVwenSoZUbm8
szqWD4HamRoTcW1TJ+kuDBkM3cmgUZ8r7JZP8Oep0T9C3MLE0FepjDcrO77KUc8S
9rkodXSTKyTXaHeoO/MY0UQyD+mOTrZteodp+2nTYDooN4NuotiBxGvI0ke2YO9G
NVBiyXzOb8KmyCjgw/682Kz8SmyaFmDyzIsM5ZwLYn1ly2eLWuCT3U/1KieJnzAp
2KUyKvRqrOjSLHKrlJm4ztAV6iQ14AUdeWXXidcA5XPhdE+nYNxYqANcYWCazsPu
nnrgJAkhvgNgt+XZRvmXKSdBLdLElHw6TJ+vI50qf3RxP7ZGg0qfzgQMNxUTTxrN
JjVwUX0S4n6erP5A/zgAhtvfbITN/gLEIEYaRbVYuefjo33OkXhYhgpXALIJT/QT
zADhaJtwFsQIJWt+5qPQA8JrJnyg322mLtuEhzCZ+X32QZkPT3rQ/axLJz+PbNBH
yEEcHLhEtSVralZbtdSMRHuuvDmYrr6FJiyPWhjsakByUKmFSyMn0vOFqvPOvbOL
pk1VWQW5utylWWHOMaa9ELrrU8blFArgj7Tr9MAYRP2X6IFyeN+R+OqhOYRG/5Ns
WQFqlpZ1QXnQtCCbUPYhvpw2Dm4J1KqO2z0/LXixXXE1HRe+olQoeoPYOZQMmVEa
90M5Mx8aWvQDMUtumpjA+6sWJ1RqiP9ovGtXQME5fqsD/jlMbx6pfLA14+XImqIC
UfEG73y0xuho2dZTBoKdgQLoct1MNmOLAIcDk98dxZ4jI0tCfoMqLhsm9MvcM+lk
kCh/6+xb79n4YhfZj5uXXzS7jHDqZFlxIma8zlqnKdo5DHulPgW7Z0455SAPo3q3
qdWgxPyxB+l/Zro1lAy+djalc2dYTNwQgA0aKFbzPxeF9ihnvprWZQkenfZ/GO4I
eRTnyedXiNLK+5YebdeQi+DWaJ4eva4KdKLdsfqrQXMXmFkPBHnDTmzX/9aw+yH+
WWIVNGs2txRYwyfI8voLwJCNKKUPrC9BpUWIe2CiRIOB6sgZ8yLveZX4RX7qreED
Sf3FhMYwLsh31a9xblNdOcuXGBkFFFEFGQqmXMyBe5fzUcqUHO9rnKwxPFNFiJoo
jZs72W/BIeHW1Ju66K3U0UfpeQpmwBYQxDhcghX/kDdj+/qTBDIzrSDhC32KPkKj
ZaV1vq4WlgxlTA0HFHwXGtAtC/bwnTtUE3TiWqw0Gn9I/9WlAFhUVY2/yua7Mod5
upl2lf0+trn6vPhN8JjHSmFOEZmoaJHJDzNXy7yjCIs04Kb4kg2SmsogzNjDx6vA
tdaK6NlTAwyJYi03fzxn9Gdf5WzmbnLDqDKtqHcG8JQwJBbT8gobpea9RwHrpYgP
A1PlP0n3is8YgPVVYtU6voZbFY4++lD6QiMhOAayal3fG6Ro8N36+m7LRgbbjyzd
hL5LVxqhUneeGahTEszjF7PWi+Z2QMKOuGq3OhAku2Rndq/J5Ve8uB0HZSGyayfZ
yWqfoWcHvY0dX+H65VwjKM847Cnh3kBiVyAuk97Ev+VJvqS4qNIMiiAvjV2TIQPC
vkEr+9a376ROcZLwvoHO44nXUTfh1phX8WO3g+s92KvijPX4Y3t14gFfhTVbL/Ix
ZEkK/zBllNf4w4gOAQiWpD8E0MQNNCsbyUxiNISlhfRCO80R2xXA9+kMKS8jle9s
5W/z6zIN1aij7H6aWuK3ZSlRoOrk7Fhyvbj31BDtU2zqXkGoyJOxN3fBjd/djRZg
WFep0hH2bM60gKL42z+pVbjG8iatdkp6YrrhwlsHbghnn18QnxrCGfaNwzfqsX1i
+Fe0Ke91Vn46awfOGr1A5UzyScX/pK78xBzr3ShDUihFKJtTggvXvXiB/Kew1lLz
KlXUXejLC2Dvz9CoXnYyj0pew5ajDgYR9BWonO25o30YFHrMPpQ4CNDze9DkMIco
wuiJm+VjeWMaudLLKUoJpZaYKiRExCWDkRVLFnh2wBJXimYxSAsc0YuLnwK0gE4i
JIXZub4pzkV6b9pOsq6vQ34HNQxf6KycqdUZzZRul9qZUMo/dOHyN+Fyct3qC+9W
cJP+RfOuhSvdVSUBNhKCqRE7XxhspbL57q4DUd+oM6m5icHQpFnAlksxGPLiOsUu
itykq5Vf2k8u3I5uZX9m1cqm7yAl1nyC7kybmHJ5gnPgGDf6Hn9ZhZFY20PeBOcj
h5xFqexHdMnDYOSRPwDfnQVSh/+jW+UuDSXrq1WScxjdIZugIAisUXE0D1X/S5EO
tpT8sfrvlfSnHEm5R4008+5TrkUGGO/Bccyt6ywsO5UcixWcjSjfI9hWmRo1ypOR
eOP6wvvWEkPu6osOE0nCtNv2r+OPygRd37C4PKPLDQ6xsL2CeOsE3M58VoyyNZJi
eOyTNehjLRt/DYqc9TKpncwZFPxCqYlU3iVCK/ufJjX6NJSuFls7GJX5yisVHVNd
G+Mz9gjtw/fmGercIT89+VL+r9twhoEYXitUW9ROe+0VKfsVnhFC+1ezWrgBxQMO
gFKb6uEEfuqHOomlRryvBc2rAwZcOV2RkBzX48xwnG987VcEvq7h88juh3PG/siM
/qCneBGpkZi4bC3OF5mpwXdpUFnZyEsDqsCus3Cx3PI1mFx2OW7+OCBFyzyWPVmm
YTvGZE7EHjxCarjtVJTxxmosp6GlIFG7yKT8hh6j39x1t3/7CxuuPF0mrGyBHldC
mT3deXR7U9V8wL9xFy5xVClh6y+o54pAxbd+0eucG5wZ/9CYa6exBySks2xYel30
2wHxG32W3mw9pdTmxMD5jeMfklmD62vLtcbwzhsQBFZXCrmPotQRMyGMrGdCuuQ2
A3wvtvnN1LhOv9nakFFLXaRKXFjAZ82j3yfG3Ndb8ofGm0l3l8VSJc3QhUsUzB5t
rf7AAZq3R0rmZOXQuD+JxWCjxNVTCTHKfh7OmDGQ5F4ACl25UzhuBJeWtBoHwYe3
VzCeo3+hcWKDrUYJuK2NNJ8z+QeHmrjItke7XJcL1OzaDy1CNqVhzKCPKn1MxYT4
CgqO+e0LFu+b2URqOE6uUJkdwX7FwvKEOCsq6q0GAYfD/d3AgOPsKAhx3J9yVAUw
a3KW8NoVnB4zaLlPKKcqX0nSZNtlu0BvGQG01L6zBJPd23zit2tokJJafALGOHgq
GkihN+zrC6VYtL0fJV/F5nkVIwmnMB3PUQFeYx8H9G4eL0NDEsM9AF46XsQ13czd
yWnEdCPTEB83vCFVKq1XJ25ymCywV2N1GYuYh6S24Umrsw5G/HRL05atCA0qP3Dn
/CJAGP/zBAGeK53xcFVwgpHjE0IkfSx8zt+1llxtGm94cFP3EqRiFsvjcAXudiDa
5Icbof2KgfvbQEAiMjPMAndxMsNhAka5mHCe3Gw7+bBQox2SDJM8iJB5vCjRTNuN
peFRDcuFFEGSWjWMG0PQz43IgMFe66cITnVaY6S1PNpDjPrzT5TUdVXoLGf7LCTa
ykJAEk2R8ekIrgCqluxRFul/pGlgng1wfe7Wi4K+kjaZnCoLvlaoDMtbSMBhfT/h
JtRkLX4Tlj7AQUitrLtSqbsb0Q8wrW+Mh87HSO3bNCdgTJoPdlHse4Y1Ojw8tp5v
IO62y7C0ZkZlLHPYo3m/BycigXucBiBWk8dVgvn7j86uxN+2NC55cj2u821sRpmM
Jfnref//3ET1O6t4N1wIH2lBxNk8J8AWoGn+FPNm4mfyp8RYJTW4TXG0xs9WSAaI
53ryqbRKN5QBt06dwr1mDjhQs4EYDOqTclpfxQPsOnbnNz3eA7g7rzTGJCoy6pHp
iqozwVAXU0R7W83K9pkVDHyjmIz9XEhmA6RRWmSMg+INX4CRMYWMA9cdpBv+FHTW
iLhUGXzXKqf6cCqFWTfN73unh1Y1X3gCGAyMIFfuHTtitBpc+p6oi6D69aVjo8l6
k5Jlv5lAswDBPR9Q5t5fUCC669GMqIluoiU4DOl2RoR2T8jFdJk6UkxM6Tn+nnD/
unIJzaql5ITxe1WibCFv39R9he/U+KANeuhADrwz88vwDB+lSAliG/FwaYB2307g
D/gT9vHSqquh6Crgltnv9gv0f7lrkwe7pphhYGmDGJ18zDBnu3FtulnNO1n5ErMI
FBqnOBUuFnZSZxEXmnK9Y3o06AaCilOXZPXDDcAeaod5qgSM3MdBrzB7h4C9qpH5
rS91J7nEC+4uOhfaIBjwCylOBAodYgyfL4305LLjvguarmR/eo9w5et34OtoCL8P
VkRhiWjOpI4czeYmtvgwvk/dxaV/LvvOQu2npV1igx7wkElKHx1ChLH831mn5Akp
V02d3mhAoegPHXdUNLydALwGDxLJ3kYOYeL8UOFx4ioq13ToGjpV4mZrAULI2OeO
Rn/Nq+kA5cmUpEsNRkkd6Y6ttocHygP4GWMOszu3RM/vflSFIktjDWWmZttm1Uq/
rkOm+N0pbf2SupoE+0OTyeMrECt2dGsGy1Jf+TZonkBKD7IgR9EJo//mqjCqoqCO
qcF2bE0wn3dCRxPiXRCIsrm0NTPQmaGCiad8g+dHYxCDw/O5gnvAG5gliXHc2AIG
iiqWcrjplhQFj4l2Au64d9bUN//1HTx6lStXsXcy7QBMKKGWoITa8ypw+Y78JWNi
2U+bwjUqYtXajN1DBr6rxUpFYGF5FCqUuT1vKJV/ys/Ysk9xzfB30TWqRSHrTeXa
rTkvnXOV5AnJBVHhTlW9ZQtksc/3+Ft746hjTgkmqudAMygSbfg25RQnU/xwoj0x
+yc6BsLgs8g8iDY/HdwHY0AHgDsZdW7COV4c3BoN3AEYgQ4KMLMO0YwH6sK8fg/q
axHdOtmZQqyOCZ9H+pthtzmWc9KEJQDdMhjgcDo7q2TPz3Vx/yF5aeZPPZ1o5pqZ
Xelb3KSH57zagXpqDWv81Pe6RPJ8HHXtcAFxfiV/pp1cMZn5swx3waFGfCfnhM78
XmBsUiN1mS4jLLB/75WiKCQipwvEfUEJqP4LTuvVvJiw97SE64idH9P48I9fJ+8F
Qk/krCEyPeN+ZB1E9EJZBX1muGMOqxpWpPTgNKzoahSOIH4bUCHFKtgiUAArcksc
ZCN8K/qVxLNkQV0MOB/hf4PjS2mr3wM5jO5sTW1/3YAvrGshxyMjU+3vAq2GopnS
Jn+0cGgtJmv08KhSEfjasLBEUjey+LIowVORU9pzbgxepnFF6/KMcBQ2ukvubD/s
VyBx0gbNohM7cGHYmgNHDSJWrb2Hp7lDV7Xy19sgaIyT3hfMe4NKmiIj9qHZsBm3
vdeYqDIMmrVffHzUkXNI6FCEwLSseAY7y+vecIwXuAkO7qYvxgZt0X27ENohZ5Yp
SzZ4V9YKwbPLuYqLRC2yYt2b0JXeGEXL3Xw46UP0rRqIMQ8vH9ODb/ltIIj04Hco
LxFEPuVJgupLCkjv88DYmM4S9R6b3BJ6mRO0HDWP6hYVPOraX4mVIYcH6noU3QOo
Itlkq4dbJgRV9QCRP/A1VSbYzZqr0/1Im/EwB+GasMG2hYeeBDPm9R3/stMbD0gx
mpN7Pe5cZL0CEs9BhyetqdYewzeQQ2OU0MfeC2nmKfc6vrn380lCHVfj0f3K0fVv
PhrjlGoKB+xYezj3bX0e+S5OIpFfvyeEog7x3FiSkaju5pGlk6Bj/pLo1ARkKzxM
pP/Bxobk7+UX1V6O+VazIodo8h2hu1XiSe8/2jc/Nkxa8Jjc3LlEDoIywhPnL5Ta
o+b4NC4cZf1f2OaZw7VoUDUmzokmWmsFH1MNqOJfBPel/25uQEG1n+CP3301GGWY
oK9XdBz4DkhL1T9RMT/ToLeY8ALK6cKR511LDG91+4vDe2VaOYPUzwXAr4JldlZk
D8bQMIwg5okP8EdoLAiWrdTbt2XOdo9IKy8DHYDruAVSKymZD6wgF5jvX7fQ+dT+
wvOoBQoow6JFI1HMhcXChtoSO+rZnmECbcdNRNG8EivlOjjRMTVMyGNVP4kKn1CO
mADD6bhksKHiDZlMjmlIGWH18EKmIyikj+wtcJIfSENJ5xiRRfTJhFmbcAZiTF2u
JJddExbGmvTachM+XGqr0tY7NQLu3/6/RDOoAKpDD3P3l5LVPpT27wVTwfebGXv3
mfxmjVsGqy+mc2Vm0nNXLfo1STzNqw3KVSzkIqaJlmyKZ0yDJfCvcF/rk3LbuMIE
u2b3168q8oei4coSXqYUXHbugOa01iyvOar5tFNabaHvX7BBSyLS2RpwaLarneDf
mVmkrZVVYP4T6+0UW6pv78WHoC10CCXoLH3M0vkW83qO63qDTH/ng38icit2gxFD
xZiGLDBo4EzTVB7i8vQj4Ba0+XhwBoEZwmh8z+72MVXG9jU1z6sX5msgEr2ZzuKw
6lBzQscxuUYvCZ5qvjfxKpxWoGVw61yX2puANUleKvkdqKkSaGpkwLoiiYzp8P1r
qyp3e/uu7eKYOvVzaI6UVBki46W1pjaEji6PDRJ+gXpCOC93J82qO62u3vGyocsy
m42VHxZuvFD9vdZBtUU51C3p+3AepvevCzo4sPRfdNJxG8X5SdYFJf2gFyZ3sgY2
A5N0d4ya+0EElh2vctW+aALYbxGoXUrQPe16pCeH1PoVoI6eSNSqFh+RR0WXu2KA
cQIb/FqHnf5qw5P8S3WOnAff16mFVF3++ROYvBsPh/rMjYNleQ2xQPNbGwZ67eIf
R7qfCtmBtPDYxI6toK1StQkdAOZP6VyuyqiafuWPTCy7aOnrAeyzWhXzS21eJ7we
XLVW8KYPNn4dKRZ3VtmVKgBZbrW3zS8L1kRbYwR6speYXSe1cLT5Hn8E8/kvRXFL
OirJEanz/aNTutd7kk04g7lmcN0VzMj16a7sZb2I+/4RyT8Pyq1kwkyd8CX0XZud
81G076mzkHsa9PXJhe60VloPDVLXetUVUvAM555yd6foNfMjd7ZnIDQxdExZJcZk
vz0ruMBLmW6YNTDbxhhtF3QHCvN7x09chGKRiyi+S0QbRP/GAA613Du7ywJRAtWk
UGK28jPoghFQkDS1x08wLXjAzXDkTYGwgeueRjdI7+xcK8iCoyou+FV07L/e+iV5
eHiD+VLGMTebTHr1zrJIS3nOTIFYujo1Dvlp9299Crr+jnDVRehQvqkWhsAqtlTN
wPEfPzqfjc6Nyyaksix5NjLZU6Y+1LA++9WzEZeZIsqBYMY7/H/uyKXxHK5b3Ehw
ufC4vnbzqrkylsQH8XuIQ8MUEUhBlp6T0/zUPfmxF3k2IaTrtt5BXs0deeVPIOqJ
FGHF56UAG8YGPbuW6qeg1wfc9KKkLuqmBwLKEUdvS27h8c9KuAij+bWVhf+RopZZ
5Mg7eF5tU2EO9YW8oLZSM5hnT1cKpndNYvZEptbTicLH2xe0GeQEBW+DDPJcYQhJ
FQbyZf+fDSHfT9o/EGHfQqx5bLA5EN92t3kTHkwLekf2/nqaHwqBawpXB4HSNCMJ
ONjZObzVEfvilz4DrEjyc8KqPuo5nzd+XfW6WFdStxaEps6wkh8YPk0O3o2RZ0lq
2iQqrkOwPvfQc5OIE1z3YebKO3+dr5J9Sj/mGEWPPvwI5Sdj04rggKDISG0KAt7H
XfeGf46TX5Xr/STCrPRTGHD0ezlbMUY6MYNOgB1t0J/EUHoAliW6KDrubuUE95j1
336/ncp3er/SxHZImc65hJYqY1vbdQiDXLQPoZvId5TPrSHWiuP7RBI+SXVHYpWE
GgxTCJI6xQC+il9Tn/jaND1iCKRq4DEOgMA2pAnZ8h7s+dey94vWsggDN716tupL
1Xnl9PTGwvp9tixCqkhExZjwGT1snymdWA5MbwlgQH8NP3IuPmy8VzizXhXNppXd
A9TYt+cyc6TFAfer75Hc5BfWhI4fD1PIA2V4ZtUI6Etp4wu2ffIOcG96A5vGtpOt
3HaIM67Zj/BpqTvafSJDKoEsx4N4pqGCJBIW5s8sd3c5q7AVukHHwlYX+fKtChge
uyZLi/lVVDcaLfU/UvOecMcI6kz5lx+3XaNw0h4FSrfpZl+NM8YXUBvJIHLceRrD
8Ib9bEUGLrPgX6LPRYMvdLtYVrxYhnyfPjEd+dqnrOjPtQPyQmsuY9k3MGdYHgBg
5JyHjL+xnN048P4e6jZEGTg8DaliPQuWVFxTF2GxxA09AMMTP+VQr0uFuCiEu0pd
uAvVPzfOtvqXnn3Cb73JqVvR5cFMVR03XVhRMe5RlBDsEAQtvEdjem8cvw0zyIoh
7mWBesNcewarYEfQMDnbdQrngW6w7n3ikVRDxAFmJ/VlOw5UUVqicXiUN8AtCxyE
cyOeIGSGXlRlMWXZx4f/PEJlRShbSZ7V5tz5iN6LUyze1pVCLDrfou8y1BMcqn1y
+84ltBlzvIlIU70sWsvzk4hgndQ0aTRnP8WlPjYRW6UI2JF7xHDrELny16qVV+Zn
sb9Bl8WGSXjy3uT8zSvblQLG+gnBqUj8X9YUHkR3o4GgYOdjz1fOyynMfTHKMXb6
yivT9xzMC1dxZrgkRi7W6ocot2EHVDL4fKREFKFBjqG0biZzCEEgaPViISwZ4E0B
AbDlNmSr0auRjfOTg/qskd4KNF3buW41WWWaXXTJsk5uR5Ze4DE1y/USeDALdAMF
WOa0CiB6P8D6yP2xh6BFeDRPxY/pQjQIP53Lola6hzAXnadZfQptHtqyMOLkqvWf
5+vrjHfIY7vY3QGLQULTt09ChlZrgNgp4QNaAwhh30GpYuMHiFxmCcXqgd5WqGy3
oyQMsQYzBpNlfeeHdQIcUDt+m6g5HgV9Tkzs3xEELwqQ30PzcUEjD+b55TmaQzlE
1q36XCN6hjzOb+zalBQKgZLCUG7igZSI/u5xJzXL77L0slGRpNnJELe2F0fbc6cU
Ll7V7cbXMDuzg4gtZI/7KnfdmDD+ogR2PVIi9OXmbjnIJNN6X9g7jpkz3dvE9z/k
rEjkDTz/qv9VVkfA5+DZpMD/MSt95iWnBR7xg23tAOatGTL+GaQd2Yyc7ETKa1em
A87k39VMMrrq41fDQ8Fvr5W8vCy58cwB+Meuva3zsScWSSBVoTcIOcBhvm/WnS+U
pWfaQjEiPzhoq1fTBQsqoJybAFdrh3/Hzg2vmFNB18xrTeRYiS8iEOtSOXHiHA64
mRmnOuIMvGQ6cEp3xbwtlipOECTUpJuWUxRtKK7D0M0uS3dQXKChhA/R2GPRRmoP
wOLjzfeV5c66KvgRGMQzx8GieSv3IuB5U/qRZ8NNlAfnnGo2frph2onCXj7F1wsJ
+RWuCLbcCtLly/tbdzLWp6j84bBwE2FrwiA3rRJxaT5ajTFB0bPzqtxN4DyscDpa
+WXBTgzp1r1s0+ux5lqq13GTczpQso0mqrKEUfSGYyYnZrjaIrz+MixAUBPMjT9B
95mQ+2xSU2eUVvtKIbTnLDxJ7sBrJYNQj+aJEhQz0jCbwiRVZLVgAXA/QaJc1t24
DtJGQSm16pduAnHn92LcOleVQe4E2rIV8SS8tulz+a4p0oH7KIlAiYjkss+ZXVki
+G+rgr5Wf91Riq5ztuDJCl+KNEoZXqVldV3UlyGDYPZZbrmOOwpc2x86D/ujoahJ
7WmIR3TybxAMOe94fhlQDlgJ8CTJ61UumgPXCbZ8GSwc7l2UohkIr53+wiSNBlVV
wlGqA5Uchd9r5zYXpTP98KoTaUQ8TrwMwUQRXryCo5nqty7X4ryh7BF/ImOwH+13
uGeXb3ns1jOMnR8Jj8pEZpUThXA0wOcwJTk5HnrBVgten7ym/RvvP1eHA6CgvnXF
cTTDfZF4QTRKjJOtlRsYFY+EO8FwNUZHRZco4bQVBZBKl5tZ/DsyL+j8d823T+Ue
zME2a/cN5L1G2scZOe/mmaugpWNJjgXiC9uawWn0ZgmC3jvXUurhDrD2GnkzbAMM
YttoSFsjPKx6/zG/y5l4ZqR64DsR771oa1AJALRwgfoaAuDmoGfZ0f7LICw5EqqP
nAX2kZVPALE1CdoX8klpTMW9Mp0KN2BjSm4brmtLxMPftDs3NPbrP1cxV7JjJDCf
xRd1tyK5gFucAuEHhHl4/ZU9BnVtumoWCbLDg14SwTpoSLO9xw1YBd/aO6MtDbA/
gMGxDyd+swjYp0wc90Ew7x5hGdc7S6ZilevT6iBZ9MbzhD9HdhLtfW3EDIQSSTrR
tU0x8XHvCETqWYk5DyObT3UAgD6unwCCRVX/KRC1450xftMrEDHgTEqobNyyTl7c
ApGMJeX1sjcYBIasn4XxG8ozbQ8VecLSV8cjxXpL+ih4pJpefU2t4DNMeDVVFoEK
sDU0O4q945nmKSeLX28tSUQvyzjQHFw2lq536nbXSv7l7TxjjYTIG4LpRA+h2QFR
mfX4U2SgM0DF38cxGDvAVgT5eM4pirFjlofSUzs+5NXbw0iTGAhUpQi4CL/daeWI
0TppX6RaqxRbxT9QjQgm1sEIM4LTqAtvlvYM5YR8Jwgdcad+44AnTHHyJuGx4VpA
bcfvR9ig1xsTGFGkErcPUYpLgDu8gFe3cG4GhnGkBweUTLoYZ1b/Yu/FT7AWs5Mn
s+tkW1sH4QGkW/V54zcJdrrMTaDyIdJg0GkQiiVdRHH3ESO6dEDE8J9OEvgDrz7J
urewzZwpg+KWAbp7x9/zTnr/0VHSjjbAT2mLSuMYdKU49cmFFrXasbNmy1gzlo+1
CcHlCm76Gseg67lSYU0xE4xyy56l+kCId7fKtgd3YpAlJ2InzqHswHy99izBYN99
kQPDLFvciPIjjqM8r3UIZU+LJCAWJgF9wkPAIyZmmSnfR3VNLZtMkH/BcHMli42+
5b3rOjkpRMLRmtehjYpCgNldz0s0lAxSqqfNqoS0GucpXLNXMAjY09nlBLgIGm8z
r/eINZtRlkbD8QNOWDyBiMiWG6bWltdrfFmEmvaZGpZ8wS6paCT5UVvqE4MfvAhu
1MABJai5AEsMif/yGaDaMdmiWaxOffJPZIti0okQ4upLIrh1j7OIZ6Q+H20l+JlL
nkUVMkz5ZEslQbjdqkbKkHTtyB3Uc/l462H7sVlRLFuG0ecBIGQE1SJppcA4U8z2
tyo2RIvH4wpbmfnvN+cxZBdV0zURJkc/u0OszTEozhou1zAC8HZeGPKMKs4iaBYx
TYHwrFr34eVDZQWcbCPwCZwuSiwnIrL2xxDd3d2rjbTfrYWU03td4AQHoZ6RErIn
aDYx0ND114eShdwzFEjGYzgQwKLAWZ7P267AwZ0BfdACiGfjP89Ywng7THeNsiNg
8aZjzUtJSLLbGovGyKgap+epI0mKE+xfYWvfzaP3ufjAChgfXUD0IL6XqpApG7RD
R/e61qRGCOUjuZ3PgOi0pbfEoqj/XSK63vj6Wgl61lIYgus1Y1JRwB24np0NhfXi
Kv5K7Q7Bk8XVbqIfLuD9tn8dZmo8c/at1xSNmEBx9bfW2o/+E+8jF3H53/7YijPI
no0po12We+rmf1sUXonwrOAkrIuIkugsbpFNdV+qim7aoX/je3kuffV3sYjPaL76
vKCSpAREYRPH5oTd2ulWD/Gs7b2fK7h+UnSwEEG8YRUfto8k69NYk3uBFsFyg0nA
kkS0kmJDGi9mIzJ2BfYYcg5hxhwiQaxLaXza78lDAjYtqoowHJwRKbEbjopGbdeh
Ed3erSEDLunUvia68cP49Y5HZo/lP//VWL9Ebiz/KW/tOr6sL0v2VMT9XTl9VDg+
dORqgZIQvtq3iaY4GTui9ntrSuFKW8aOjZshTycFbPhrGIlm1E5S1ktu7JqUe+FC
bkGHj2DSaXXgMYtym/MU7flZKu4THC9BsSmgYzYfo4wzjgk0rfDVlxehJCH/B9pr
OiS9pUARWu6ZUjN0fB8SgE6iZtflOSAZDWFMZS2hfFMedXZx2qq6RAdhLUl1Y9NE
vS+zKKVz+YsnRbz1CWdhghtJbil0EZ4mS/ori+nJBbn25IOieBMBN+9vKSc9dlSH
jJuni5VQYdeTgBrsOr0KW8rkzu+JJz41SpEmU8cOeStVrWN+no8QlisBQcIZIyz/
8Etkl5r1ofdAPDgPrxMpuRchmesoKSnod0foT5GM3L8tO9ev5Kg136FPsypRyQ5T
waTFZxmkWnKR3KLez6MOT2gF3bdFYL+q9Uxbc0pOK4pJbTt5pf3Z6OklFYqYG5nw
awlJpOTP25zSTSH8OYdMQ9J6gfF6fDIdhl/7VdMWmuPD5DhlVOCz/6IP7+QkaXHB
nQROeN4nF3qZ4dMFsjSZy58qnQsC+Wt7ldMojVZ9GyGZ8XtZbdeiM1WQAgBm4fVK
CYWb3wRt8itFdMnncSCU3yzr5P61cASkq9BEUBSy5DDULzZ4/kpggP9xOBYX3O2R
yhdRq5jX+FPt5kd+18SCsCyovs9yITwR55Ar8EchYFLLk9DU/sG5VnuPJ5zq5JWv
ybjqtrg9QNTbcHSEmYJH5FMa0shKwWKmNEB+yD0eFTLQCdEUMdd6nY65M47iztHR
CScWsB01uUnT5TYnySQpbwGzYvhwoXcgSZaM5GUCU/p6TncOSYwTKFa7lBjIt+aD
9F+ntZOOiTW2jF68JHpvK9qeowOXkLZMRH15bdQOqjRQkJW2e9Mts+WVp9vtha1G
FAUBUzMhJZl7X0+n+3M3vOPFOjvdFfZPDckcWHN0702uDwBffRTxIrIBtI1xIk9t
5/1+3eAYuy3x303FFmowm591h9wkG0ZgMDP6EA15JzAspXieTaq+MbQAsLXaN/3o
yTpQHrPTpT+GZN7N9Ot/CT5+/e1qR8yFX/nLs6gpJj1TmXeMzPreX5yexpHiAShD
tC3Ms9M2JRq8Tj3fkenYclq22fhl66hm449QvSANYWFCT+JrcE926xDEk+AMgE3y
8BjG61CjIcrA+tIHl5N2wvlnjzQSzIAeyiRX2zGH+VLO1ku2+7ONgA0fgSWbnVzr
1WsYB30kI/tlrNnrDVFXYLucMRlcybUmMwlBIrbNVrKeHzfxuC8on6kVycVvNfRM
03wbTqJFrDMip+ZnQoqdgpKbjQsUSmqAj90Vvum7WxiGlqQwGR6mH9BlcZuhTvv1
pAAjIwT/RN3D2rGB5l1qbGmZN/fPRkOUi7BzcL72hyGUXt5YlXF52WszG8ZTP7yJ
/4JhfNzakGl2eOQdC5/SkEX44Z+CYihY+CqAmG14mAmdU7xIRto2gaXzbqd2ovOm
uR8S21moWZQrHLm7igrb+ZuOtRJyNKWVdVBpXQ/b6LspaqYRM289lYKTC+1/ua0N
2MJje3tHdHa2F+2iFEAQacMwuP6E8uW5WIV35N0WNDejevKnazyAMQ7JRNsUJdkU
GEErkt+myuKxZ/r4tYXwRPK+Avhw4ZVAVwtONUw0Dpkqy6BlkTOUAmyKXLdc/gZE
OXfSorTvhOOamLUBELE6W7yyTWX/k7Eu5XO7cg3Vo/MzZ+epvSUiyHeC3s5iaHj7
iZE6ohccphImgu7N7NPsv2ObGpFeIa/ePLs6a6ZPYc0WIonT4J7AK++gIiU0W5pZ
EYxyzWfGhkJTe97qq/e5ss4IWaGh4BfFNPonwGyYfYLk3uhaf4N6ewwmC9UL1iG8
O/G3zWwX5jjlzuzM7ZiJhnENFIuFL7S4ByZ77xrMLtXXs1/g2DKfirdOwHksx10k
cgo9Qlz6WonvVG1Ds1VY4JeZLYi9t+JHXrl+b8C6/ds54hQphLI4hx6dYdz6d7n5
/Oy89dV2oBZDofcGhd8IqFKyPP7A7tsN1qxZaaw7eFAnL4gP9puK5mfR3gRPBp9r
85Y6PgjJVFR++kpILzVdd//nJWUbSjG5nDWsJ8qIHZ9zrvc2lOyp6jVC4FVvJCGS
1wMHMPBFIYfRkRdtjKAXBFbIiy3DpA8hiFOuYrSQqOqpRz5Vcq/pavsGmCKHrOoS
Jb9Xor4FeMc81Z17ere8UCwFffGBzFTvVa1flAUIzDgQ5Tb4+INnKNLEYLnfrbZ3
IQ2u2nHOmIrvQJLcv4/QxbCY4DNUNqTAUX7csnjfPvH2Ov1OAl7gamLz0nqq4aq+
gp47JDb615y3ZQcR4ciLle0J+F0USTv8+LJjzVOym9RnuJam0PZbgMD2juXq+Nla
fRtEhyWYXO5fm/fhOHVd1GK4YutOCwbwbM1ZTs9xQ7Dgjq+Kuax2Iv6K0dxEsFRV
gLFKMSPb/riY904ZYxuW7DMdDiD//AFFxboaXs6KsNac99T2ZIFo780K9kt4ZVEh
7LG7K5b+/FHJst/1d6Up2cv+1vlqvUTx6wMHgJ0tX7c/2yzP/OgFHkOe5MesZ74s
fCkyMHTH0liTRfXCV11NKfiJbuZyFpNhAM/On+F6wsn5+z4813f6KstTu9YJTgRa
nHdluEEqqWbXer0UPgLx8lu34KgegXtvS2jelD3UXbzzA1HZV4/Si3M05sLm6tb6
9ZSOUuJHk84/QvYIhy0ANoU0gzKisWtJ5XX0Of7la5X62zsCdQ+4KBR+6jWcN40W
LL4WEZH97D+4S8JpPKRYuzXPEm6gI+oNeY0gS40PYVFVdbdtCg4Rbdv0Cn5hK0aZ
/MBRGdGs4uL/oF4MFe9OEojpaBhea4MQlWgL3iTz6v6UPKValcYKWPoCspHSYLun
qmAsxp4vuTRONoK5lPlcQ3J0cGlMv2a/zhVc7GxXO7DWiN7USQjUT4PQx10LYzqq
IACzJxD7FJF769IqqQNx2zqCGx8WXuRtyezC3ODVklxWL3sUaXQgkuSyD0+ZxSz2
zlEGwp+EIxATZtDc7k86rkjYF7UwaPw8+Ba9meDvnGuAu6+79OfKhecwzCHF2Hds
fx6dzJbMeOBy3txNMw8qyLk7RGnvYpZqhejrKkZy+7I+zK2dDJibtYcs2cbkDGmr
bBaEE9964gKi1GUAhroAuy9wFHl5M6L4GigDRy1TGygJ4cdLnfTqik3igEreZTNq
8gFiio8et2IKLon4IYwtexH+8ZV4WkVIJdGxmXpZZyQzmSMZuT3AQeGQxNN48Nft
j622dXcBF7bGqv/VFxatEDJuVZuGHBRxrKEtn7lDOpYko+Al1Ggp3JWwINo9WkgP
sxYW5IJQZgaExvanWe9nwoLZH4vZSUQFcOb6dfdQggq3MrUjwFqvxsa6JrhgcVVm
2eC3BgGm5k6wZVpScgw+iFNc0Es4UsvajVfANzY54QmzasDA9clxBXNoiwQTgQpI
sCBacRq9v74VBzK5EENNzcJLl5RrIMYlKEfvw56eURx0l+cby5EHLyCI3SK0zR5Z
4M4A01nJMxo3CXDlG6uk64EKRVq7nkaQZLSflIB8l8ehjxzmCU8e4KN16i0aBWqF
1sjhnzCv9hWz9lhO0ZoLLjYwiwf2i1+oGzJ0yX4icB0YFQJy6jwwg0U94QiiJRKP
gehLX/p+Hw3MR1cuRVCgcynMIrS18UMSacqaGnQlepMNEksY2gnxJBin9lDP47pQ
OyZhoifrshxjb4dM+2tA0YTJqvIoGmZvSY5Ars43re3APahiUDzdEKjMO2K5vBd+
SlvfIsvbbXaEHFPYj5JHSTOidnjvUaq3ZUW4rkJ0hKgjSBr8uZ0WmYW8YG3rKySH
oMn7rSE8SfH7KHGVSW/I/V27p9wW6n9EWQOh9O0cE+PXz8MCnrRBo5TibP08cl+/
tBQKDb1uZcyfZPxuXFwZK3Hn1D77tk6rL1fSMOd0rRd3iNOqS3WMqhDXzT6inWvQ
WefW7JVK6uRXkOksUTVRZ/qSmC3bEeLcCPmSZomF7meig6g58VuJsrNbouVs/vJ4
Rai8IuvmrNw3Z2D3349IEFzTnBqUKTGb+jg7c6YUYTWdYYlCKoROU+k7qH3et2hs
gmBL0XPKdsZk7Gz5mrwNwVsi1z16+sXWHnhnWrffn0u+lxG03z4aYX4JbVh+WmdK
68FmMvrEQudoPC58KhxyEyYabj1dIfNfSpLwDgi65U5kT709GQNa0LP7baIcHXzt
zocjrlAiFVq4nwflvs4OMxVcJg7gsTBf8Q/VJ9afGg9U7CoyOmKYlnw54yeQelbl
xqfVJzEe0d4PI8X1bwmZKF3iM0bSUOeuzv3lGTJEsVCFQYhIgebJ/BHlOH09fsu3
zoPSAJ4+dZxJVGuTqPqh75yqnsI2YDGWBALMObUrrO8BPi1ZnS7mBZTLo84npllL
Tp9C+/BUUK6OjkHIQLtaxL3gZjW778qYXRP1cMJeBtTGy+75nMBXbwzokfyE6Z0o
Q2O+DGM5ZeJYq5gwNX0/tcle90GkGgwBq5x/6x/joUzUW5d+3MFMLMhJozhL6v6O
DfxFoyN1nMVBjKkFVBuOKjkF/7A2aauZ6pfeSMZ1m9m0zPtQXduE4J1ck6+YWDqr
sAaZm0ymGMHaRA05m8i6aVkI5Qqw8MMtYVDH+HdGW6e/fcPGTx56CFhc1rVkwPck
mm+/zrqyyLwckCDOygr/GyNNwCAjRCulXIX0kbSDOsrLSHrIEAHMuPMKpb3uVN0r
HjUCSATVisbiE0R+aG+zKxvjoArLB65gNj1cIjslXpozDTHD0p8xnfUoLxea6Dck
N9B35oBYFt6c3QCageG9K4T60b6tm6n6k65BDXL6dO4fwO8UjF3Au9pvD5TlWR+Z
7msmgwgOy/ACjlb/TLyP6Kctpl1NyRDmiO2GlTId4ghylLtYtWAdvXCSeq4CkEhM
BCp6tHxz4r0Ue3fzNS2LVQJfVuF/9nKqdhh17f/Uhde/3TICPkw0P9Cz4R3HcphA
l+XBW90qlK6FFfu2VcCmsdnKFBedUTsOmgesVNYCZzR2BVD0TQRdaiK5qVyDV7mw
dQ+e/m8eweQHH3dG/SDmPtTGhvBw4TR6Q89eImVEa5XIF7Hsy9l62Hez7Fp5Qynh
wV2LmMMmSoVnTBl/vu4T+bvSpzvMdMuUhv+5yROWgpSKixwA7BXxNpOJCRGVk6jk
WC33p6+LxSKexb5lP16XgmTsg/fW+Ovc5Qo781U72P5FCLgKoB+DfDXgCJWH11DL
Nhq4a3IsomGJ0YQ4WMb8gX9m+8JxWgurV3BBm+PZYmm7HBsw1PicrWaZ0eS0WQTB
mOMQ9YfrXF0/aMC0ERdOyVyt/b6XFbALKWduwW+eCO89j3EpDem8sz251hwq7XFR
t8Pe5mz+1a0rX6j3JA+Chvn0MLO4+uqi9FIeASKParWUJ0GtDwKsnM5+6sqjAF07
srEH7nMg3qq/1WL6bbIUhY1Zu5y31KJooO3Hjmh8/wWCq/pfxqkFTi7FYJLwarLS
rWgohVwcyi+tgZsefqKxOkP+dEvqitDEu5yyDC6mpde9C7PeD0Per+lr5CH1xyWJ
UmDezhlQciuyi7oyQfnriO9VOBLtKm6lPJnr2/VMkmVIVLNuY06ffvGIuD3H0e5A
fMwGCKY7a+v2AUqXEMro7oBL29X9G9dAvVuTG5thmuSQkV80q5ITbE5rPrD4gv2v
mo5p9uQ+5EqdZWH+RUVBWIoLqkwX/jJ+JJ4dh7BHg01kE5kzNrMUo8kHu0Y93Wer
SxDbZx3nedxj3Pavorg8eQ6Sl5I0jPTNnwVaOUYEcYayNxZG3J6ytEEo+ji6Pvy5
39E+mvfWRjA0/VRuVDXTjrPkYBxKrmYE0iPzX2icBPB9smcWl2rd98+LXCfnlLsn
VzIZtNBpOT2Tkggzvda1nusl4TU+5HovBWCT08LCjlHzUhUen/8fJw35GY8Mk3tB
NWy58iktlSTljS8gQ76V3OsHnWtj/OVLgtAGN6pt6RgOIERo06z/Ey2bQKU7IKNU
pu46aRxOdZdlsu2M1I82+0mRdRTAyJvL32aAaqdnzf7qPPt6TKQrrLgQsw1bWORV
coy3CkI+NzNj4FvV5g8R1NOqezQ+a+aI1gXeSUE/kw28J8bdwvfgd4WzKprcRbZE
iCLwlc/EMo/ZaA7svO9fX1rUiqqd9GmWfUuZQXcVi2IOLMBzDqGaw19rIGmFg+IG
vyonCh0yuo25KqJ53buU7P/DUHuPXp/NqE3YsYk631hIVzFXOqgVIBgrM6Y++xqo
nDtfQCkOEhACnWGQKAbl3H34NqNai1pjN9Xz04if46725CmkVgMs/iOKrQPfJUow
jAU746i8ltPOl7Zz5CxJQVQuI+zQVnMGnIqRZO0h3vz2RtfdABZzus0qTxocpRRq
0DLyYA5D3JdJTtKC3kyK11VFqQJvkyMXxoN/Yn48NkdA58g7M797L3eOYrI0KUG0
pZchI5UKIRsbu/QndhSf1kCAs6ugjO7/TPJM0MTDcHaRLWWZb6sJD+0wlDjxOP5C
pZ9eS58esxNUj/k1lEiekVbYfTdsSmtAxg4KQDI/soBms+uernLB71NT+qUC+0Ie
WYZ8raRvW2DEeS2rWt5n/WAY91t2zksNEZ8gWRa6SGBtrRQQQv2kJTWyVvoUZGjP
/4wikKnXpnsCNvgeCRXezvmBgOek/dsuAYSWBTecCm7gbEZgxzpSfdA3WW65Lo1v
qX1Dj8JzbPiUF5IncR0COMFlrcosNPzJLa2Nn0C1XAUS2Iw8dKk2GP9zSRgoGq88
EgiOB2F9TmJuEvnx1GDYhAxl8T7zBauRLq4bHJlILzyXfuTN1vDWR4tGXYZtY2sB
IG9tXSF/pULgPgYxYgYxey3cU4n2PrKwD4LhAnvS8LmS+7VgLZ+udTKfh8Ku+de3
mAX7qJNOTqyfK/yEhDDnbbMIcvChlrlzQLW2IMDagU9BsPCrbTeY7rBxnDx1ybig
p8aKsD5csFpis1Cu/pXHt80v4iFBmWT1k88hQ+DzY4F41KPOhSdqpMHpLxQ2D431
oWEdG4/bEbQLBB2amuiR33Dn+Az3XhZfudlrQDUW4ZKMGSrEIsdoGtezX8g6aqXL
PWq3Q5lx6y/C4r9e6b9Ji1KQBcRX7HFNcvz27miwFu61AVhe2zM15srr6Senx/nb
91r3pcEzBZVfEbnYpmg9Eto/dDaCFtbobCh6tZ1QFBeEghj83pi4heAEdm5qi21j
YIM0AZl7G2evl28SV2JWON4auDSYeZKplx7SPsk7AtIr0usDq3CrOLz0/0ndtVpj
n6OOeSEQzPMj4qJi9V2SGxWUTT5tu6/zj1cTfHpqFprxQIir220TgXM/yEzzL4SI
DC25N4wgvfVlL0Cppi8Yco/1gvQVNerEUU4Eu5+YyjHiagpsOPChTp3Bu4FdRinH
7ty3cCtJgA0AHAkoP7rCbj6yqUpHn4TZ67w4TGKiw8zivyEuqqiGP0YDi1g4ul7f
RfBhibYf333j/agD90IbU+mBasdmOwldlGUc50YOSA3TE7or627wdDxfRq+cVNMb
nBLrxuslPEYYi2u2A31od77HTLyqXYk0x1qVItNvs+kQthrYzh29bmIC0ma/SEuh
ixBS/8tGJ4ysV6OtqrokYhI76ujFgP2rr0Mb38tNttq77couRk5wSf2uVgM/iJAy
ANaar++HOW0kpBqshF5YhYD+GIeVBKGo3XYfnOisVJfLdBR0s/xvnN5OZUSmHfxq
Rho9vKtfN53vPLghfpV7popLgOGvDjJy8YDrmx/h2mo/XW31XKEOswnXpR0OxsoX
Vi9jI0uLm6ZuiVlNkeuh+LeTQwBcO4bz3dOV7/yB3bfgNamfBrLdJoi5tA+EVII1
VqUUkKTWa4QSLwjDrhdEitJIlDTq/I4EwcGSPlLYE7zIsjE0m1HBR1wPNSxS3MV1
NK4G01cfzNm/7DC58FvFZ09SBYCwUHUn0MRRRlHoYMR4HJLAWz5OQ+962WCy1shx
LH5HO5ZpOASfEGhsfxIz8P+oW/lz5mnTI63SqZJh5fveXkVPe3CiBbK/Qx/ItuT1
gj/jdLnCU7tuym7+fcHBOjzL/WuK5tkq9zcSuk+tNdNPmmqCuJ2h/C+9x05t6/aC
TdBrgaaTozvKALonOGi8pOZwSSIXm5c+hTY/lerJsPaQ7wxSC2tb95yJRaj5Y2YI
owyWHVS0dDhP8WXOC95wmafxdVa4LnjY2D9CmKEb4e5cm8JC5O6Dl9K3+1a7fbfx
Yn8VDehHYCdkQyj2vAoqeSJ7jMObKrkF/wiOikV008FzrQc+Cd/ZKHQAUib66pdB
WPdOHahrXC9P+78eec/sGXcB3PQaTQ9SgtOXL2D1j41AuyDcyRZUvfYJCJjTLQc2
JAyr0+n8GooKyUg92frwV/jccQxIdO9NzmkAIGUG0RVsK2H8FeXzcItIM3E6wycW
NXdsAHDTa2wIJYiECc1mk1vjk+VxsMJUqqbs5tzH3RT2grXi0KeV/SpSJEYKSuV5
wkgjXuPNCoo811wwCUe0y/EdIDCjzTPljpO73Xk/7eFJTyMlOKz/5oze1ePJZsqO
VH315HOlQqO15etn3xiPb6SWc5QhH5XSN+lRIH5VyAtIcCpbc2ZxseoNIUosawYW
W21n970cTkhNX6lY+8HKiytQYPnWfg1tQzwTRRjdtqYqNX1thNkVFGwD75Ivw386
0MbO+PlTnJ0fONcKerdKdUg6xsPQw+HnsRA2cAVk22sjK7gkhnC6V4bF6aVHR9zJ
DHAbhT+Bhli73vfTGnk+nyVAKNzaFvYBDFgrs0Etg0wQAbMCTa8rvFWX+bIFch4m
U10L7+FLHcfcFwzKANGxQX/YsPjfst2srIz2AARTsJ4AiF6WWOygxl8DNYhYlQ6Q
pdN4mrj2R1TgS7hbnm4oDPWKhac+33SYyEu0Ru9c4FzVDyia8V525FzOG+rhxecF
Bv82CJIiJsp18yqtdrXMyCMFSnqu3lK6yLfHyAX8w6fgOz1HeMi4t5ZtwcjlSAUi
MCQ2EXY/bs9LLTLfWenhMCsoPDCQ1ayatZSkWEUeBbtLbj8rEZYzGMOEehYwH1Cq
EG8SxClBYnoO2y90C98WjWqlViXmMGIm1Uu/cmMM2rMHxhEJEuzk1ajA7uaRmvhB
cmXL1n8ngXcV35yr2yWA7zI/H7f90OIzSThDzPD8h1JXA4HMj2OJiKdci4N+4QYr
lPBYlhvkGxuGXBRcCN6JqeTEElhVxjY1InN3CXpmNbHwY7HHfcKoI6ynj6KWFj3Q
hNagpvkAaUTJKv96J+NZOb/Jum5mrx8IRzHupGUc35DCxz7Jt1LPT1Mu2p87SRkK
pbBBfdmFKyZcZOBH5aVNdEcBfjov1oBQ/RddPlPNBNsSCpBCPnHVJQlI/mGPCwEV
yGb7jDqjdMCwcJOoPvqQm7Jk2sQBQ7OHMYMd6rb1XR2/ymzP0anPilYACX8O0vUh
1NvjwTxpuejxiKsXBgTB4goD3cIDnsF5vR2JW6yK0cufPIc6vXPCNhqvoSOd3mtV
Bo3YrymBTvOOxFQiUle2h2htIj7i9bCJroSCDYxJ/vID+ZQPKuXNMqvQXC3hORfp
89jIh3CUQybnAH+QuSX5pcZmc3A+dOB0mL5m6EEeaT3deY2U4w24WNl+UexgMYC7
51DXJ3O5/vV/ltnRt0/Wzwza9x8yeWVQyBZ3Whjyv5M3ysBclwZ+ztN7j4iSWyEZ
iuSgzOkhtsl6bSrasbVxJEWnjMaYXSOYMVCs5FV9gOcXqEyaunhXfP+9p8ov0JS+
w6AYaeyghCG+ggyflRhi9QdyXBLPcOSsmvwYrO4z6V8MDToKb3/euGV4FjkR8nLG
MkebsLz1do4fR+XFX+WZrrjvqBI6VarEc1racaWxyGlx5g3/8wya45ZIBecQ7kym
wFNLcg5b82j5TPCWhRnUC19DXjrsxQRp1BiWXChtukJ3vsnHn7dSu0a/+uI48tgL
DpGvf2DSUlWthUVLxYFpWvfLqw+NSpJp4LQiFgiHHTorA1QkizAxnC0Tgkt2GG1K
S0Pkyfe74ESR3FxssReU81G7EdVNNT6WQjZbzkTsnNCTzDLmcS0xRQFBROZZyPBC
Q6kFNSqAVzSoXnqV1mFeoC+rx34xoQJ9zANCUFOgOpnJ1TcN4p+z199kv/G19ZUS
BHkTxG9Ohg0ymTOnoL7cMIkzmWja6BFvlZvc1kMTq3h5qIFRMzVA1L0wT+Pgas3k
5nfP+LDyUMW2pF7yKK4hp7/CN9pUt4H3HaJwEvvFSb49fdP8d/44UM9oDUN3BFbR
GjmadmwXRCkYwVL3Mz5DrMIBtw2u0H6MJ/viaZj1MD8+Lt/h6lORsbzP8KlUNi0e
C4OIvHeZYg/XLC+06BpdVJ37W+xPHo5KtJxQEVpLHU8FU2bHQkz0XYXO3v5OIZZq
y2X7lXbWYrNlm0fj6wjfsYld+w+ycKitn2RlHihJBGOVGhPasZpSjzM6ZjiOwXpS
IRS++NEmQHPj1tW6mGBiP6k81T0JJRvL+eFr/wHekIFVdTuvBU3RIHnjH9LyZ7OL
RRCn6wmMSL0IKnf72fC+ZYhLXTHeCPPlBbQ8WGNndV9QWyGdy999aLhDcTlZ9J4a
qYvrsCiHDhCwiKluRyzKFn+gZ+qgXEjqUxC64lI56JrT/N6Xo8HorJg1fzlupHnW
TKjUIBNArE0DiM/+BBtvT9wP8HHfr7fR9uIA6ICCSg4K7lqKCEBf/KFjX8Hud8oz
hlXqicSCi4juyqg4TTsrT/eH68n8MpkuiKuUSAAVQs+syttb06ayOE3Bk1Yoy2I1
PD5/L58kknPQhFYz5rgk41QkdXtWu0R/IjUi4bMXfXNZR1wkUwZ/TFMFBifnZxLG
qTSnkyVH9wFCM4rfdPpwbMHCz6xyMTIcqAR5ok6uuFpDT8TEP8SFZ4/g4Wyov4Dm
gIoPpCBhLe2Sjhp9x6yUdYc+EzWCy7S/f3Zl0eIyaYhA3kVITmC8flBJltcT6p9a
ZEthjHTxGyqH4keE57OLd1o//2vzvDwyEFJzsBCgGGVDLPGIWs7puwHBat/WeTkB
7dXurzcPwq5WZTFEdRkZY3RmI5qzVGHbGIVY6gFf8lHUsUxYUaddKVuBJaFHVNPr
wpuMfS4aRXc6LfZlumQknnezyukAoe9ttL2Fz1oLm9+8/++kMkq6Iilbq6NwVLhS
QyCfJSlS8CfxAllg0LAxZ7SUWPwxSxZDHMzZAdw1z4RVjlb2wfeZlvtr5Pcm7E87
5BoJbjReGHYmYdIt7BpGOqi3NAa7Av72zfrK1Kwrga9Xrbo4aH5f1HplHl+lKx7Y
HYQQYgu6vRrYnW6ItVcsEWV7izHDPE8yTzSGPy9wXpAMYRQ0TByb9RJdWLSOkCEM
lnW50FoZRLr6shs1GELb6upfVX+WMagZ3srjuKZAmD+J38gceNb/32WJgoU8p68r
kYaRRmJgi3IulXVIZWpPkmr52nUwhwKHl307coj6pe0rFF3+KSqv4FLi90sVGhQ1
vatqtWKPGbljTnpxSsb5N6fawdWqpKlu7myysmRQ6gU9jpry3Utk/cZgig/UEWHY
tS3rQjfri1GRcpGaXH4LJCYhibKc2q0GS6EYEsrcpyohQUe+tTckKsrcuSwYI/bJ
DH6aqWeEjrxhFCCQ2N4VlR6S9lPC+0YlqZGUZR20i9EL6n5apzKV/u93p4RRP+We
ClYYR9Da+6IqUAOeAuxSL5kCfpAs5j7ZnjaJ3T343prHG41CVIIgjO4cE3tiEyCy
kfacESEPl0yIXr6KvoSYY0ML6Mc35cGVIrv+vnUG7HETlIxU5TCEy5vwvn8VZ6El
/O5VXxk9uKGl2Iq2I7aMl5F7xVhIHE2+R5ExfL4xisBUFtlVKkVjWfiYFpwoBEAR
pbxwMoD1EzZehmdj/AJHfjwGvI1KjAHf+N4t2IdjPLUgMvs7MCLE7qS2xweTKHa6
2udiNIj/sKrW2MBTjb8BECBlRvhsNC9cpJMnRiZ7GCAhdLNP8VgvoOV6TG12S5qo
yz/jKpgL85am5K+04mdrAuPKYQ+4MKFVWG7CFeFsa2n6/M5xcXZuhoul+p2ruwFo
EpP0UXJrKUPbwE8TZAruFYw8CFqac9m2Zbrcm3LS78s+JWh7r1I+prgAJdKReHAV
ycBbiCW4s7+u9lT46TLGOL5o1rZLsUD79BYR3aJFzAVkt5SdSVZBtP7MZjnW6vG8
jcUcxeCEcnqH3w4V+Y1tc2IqnAhFuTTmUWAf9iu8qwxgvgAxkTE7itRctMNSCp5t
PuwJjKgU6MN6LGAsel65qyg/9HRv5mhtSCAdsvt7DzVbson+UvS9CHSaqY//iGyl
V7/jmTn2KOh5QHgxM3wYdQmKHBBk0QrXm0WR7cbi9qY3ayXB0/hM7PiPBnz0MppV
feHAmHOhU6nzUj7Ri8r+/S7YDBUk/tTUP2wkmNiEtmqfL2LRhPftdsw0eHihbdN1
esd5V5FyROhz8GMBx3ivVOiLSuE0fjAUyzloD7UILnW1Ak3AhVvIcTOvnUNXEgyb
frEIFiDhhiGh9QS73fZTcN0ysX1PGIRjIdXWUXiTx/wkzCVatWAKLclWZ0cbIXIc
Tb4F5O3yZJhovrL42vFow3S2wbhM03pOWRNHBXvMK0dX+MM8C1OZw82UeH6fJyoz
x5dAwHSXXhg7RJOllt2b+YuJx2aFV+cTQdxdbnfkF3g5QIM/aPOyD4UiDyCNNl9x
tpRJj948jrYRtiNt0LZ82p8EBBiVO0kTaX8/4W3cafr429rbCBpJSsd4vhU4jpFB
+NsI8kqVOrbdq9iwQ7CbcVZly8aEUQHGogg+h3V0N0g6fiUrWDlw9pvd4XF1gDt5
zGE8V4ubV7UR7ZStBC/NWEVoroEkQa7l70RqivDySb9ZplZD/qQxWitZ89YYfPq+
9UsL9f8c4CssgG+fQ3YuauGi8s28HOTn0vfcaCNaklkIciR5jsISw8oAai0o/xUl
jWXTxOr1IS9p0gfHZ/Kk+8lp5SkYE8faVHNGFxsIxrLx6psYEJ/LtwwIU2YzRXMM
uII+bM1fwSN8rxV9+4xVvzkQKM58Saxmpjs7+cuBKi+KUjQQrPtMLaaleILI1nqX
xy+F748mWfSHsbHbEc6xbp+Ffo2B5JP06YnBMMNe3lCkvn7d0yy2PerXDZp7Znlh
K+pmvz9k08O3GyDxfeESt+rJ0ydF8nnJa4y4r61s3gRygwrK3aLwpebP9IE/XXWV
H5DC/4tPqjjKzzB1fURcmg6JFDohSe1QHgecw1WjDZOrCaRUJBTyUMSN5+fXwP/V
lRa8RiQB1Fd1dJIiM44OdEowskCn3o4WdoxabiJ7SNevIXh2Lmv0JPsBQ+6EL5J5
3b7Lvn0i6/bBEb1OlNFA67onVMqQZOipT2A1xuGWsz7UmdRb8ME04KDKenu64Mix
JVgaExa/YS+o5MScVu0yb1qHQdvRGvlg23JhmF2zFyNu7r47IxUCIhNxHZjWGr48
ogggb0WoNhDeP3pAvdnntKAUWJfUJWuBnh7O+yMTMcdSN4Sr2qHLjFhjv188Cc+A
E81/sIQweLE+ZTmEeOBJS2fj23uwqScvUGU3tCbzWiDaGRcGvQzcXmR2kIp+YNuM
0lkUJ7q4EM5StArVXcaIHS5RKvdcJvf66l7N5ptsZZcaViDEspqVUQVzQFJ1/+5w
BeWUHXBl/eQ/TOnh++TlQUZayOGMW3L4akd4EB6kjL+/56OSgnkq2J25MZ6ZoOkn
fvFTt/utG4J1rzS5zCzpAcKR4zLqMvOG+Nlu92yfZ9vanCQqEOXG25y8detnURsg
x5HEZ4qYOMYNcFeAw/rqkTOXPgN9PPPonCB1SibcA9zuU3PyYuX+uveR/zejIOnC
ig5/7StZZpzxTnlkUaWAftPdu8olH2thuLVkurms4XvD0FQ0trNk9RGgXO0tY5ZK
NkbFwbrdmkRcyAgCvsF5Dh7UawMsOfC7Ed9+lw7FeoNfRDvIWjBnH97Qyt3EwVgm
gtrZZ9xOOFeMitx+9Zm3Xi+1gBKBS2BS0VapEZX9GAkv83kjG+hKWmgXWgYLzywQ
qxYIeH4IpDjTqSKkzUDdB01MlWzINg5qLP8ab2MTSsjByPaK3TtSwp7xWPkxDYe9
niFSnTmpe33157iWVOgYkjgfOqqMKWT6vSUQ3VDcP6Hu/t5Uead1fX0Q5Sn7cOJU
e75LcQqiiQ/UOrzs1zKy5wLtLgw5oSzop8XbJp7wIZ04B0IwYF/z3osa+LfAPLJt
Mh9UQAHT/cd8H6IqO7dxGKiVNO9IU4aE2j7fDUvXOHco0gPhSYRa8DV5a2FzSLET
6tpAjbjKHfL25NidbaJPS7bznNMl/gWKfkKfV5gfAU2ZRe9FrMCyTyvkBKadA80Z
g5TagzY3Vpu1tm7TNFnhvjG07Lt9nuI6twO5+5EbTOdZ34hh30P8ZDYdJEhrWety
+yRUL1e3qdjP0TJi7HwAxn2RA/x+/XFBSJAKbFba8xu8UwWevIhzjjfeL6sZVb61
A1Z2m5ZEFqcHIapFVNJ9K0mEnRMz//36zbXquf6sgJ8VXN70noNjaakE31MfxZRU
2LeQQTglFpq4xz4GL0oawOou1r3vP/Dyy8XjVTDr+P5enDCSbhlcpzWYpOxBQol6
RTPFg0A1uqYBxTrQ6O4CPXVQAhNpa5KOE/AuwdU2gb91j0mxnspZDKKTQv+rgVjE
r6p0NCFaeUTmeWRmkaQ2SYOw/4BJKlAUl4UplmbantUnNwThFmDbN9sjy/Jo2yZD
AUoiRihpMNKoGqRnl7luYGKcjgtS6/poyFfIwpzQ/ra42saiUStWMHh2KUHfeuwP
B29zyA2PcD0E0YTY8YtsiFat6VDQ3/0F5JvJRLZe4HIsz744A1jCn7hf71iBYGjS
IT6VBDSJQFYJ5kCgwgqyZOK22Ky7e8zQyWRTw91TQb07GMpFPlyiV6WJYPEugRob
kl+Moi0wnGglEM/eddMa5GX/loy2/NPSR4hNkovFvuxMD4/W7G+wO8/WCzn0WLCP
PHSwY17eo/umczMXJ3VdkgrWKoT9V1vw+MPPJvvNNyb6BaH4wkW+ByRxmGnj1iZM
+Xzcic0qYinEtfXyhKdeVzozemPo++QVZs7ziPmcNnIbyvsM88Fu9urC9grObL8Z
vMsQIteWuEU5hhtTait3IR5RIZfIaqA3lHXVbzJLXqbIbwtEYFFg6IGKMe5ECkjA
j5s7HC8apCl55UiE3t/2comEgoFMkzaA45v8BaXyyXe/U3egxyz0HIzud30HMmAJ
pJtSs8wJj4NNZfH1P1z3kVBFj1KOruzilkkzYQ+VxCWcFwsGemk5cYEjHZQonbly
6uxSPHN6KFXPOZkkko7P1uIuosViQu2+q6QoR80H5+qTXomJQqPR2kvYn+l0Zx16
TBV81Ad7dWvlqeywmc5osYdclD6qIGUMYrAhahBOEVGztaTL5IDRFMBvjmVoaKzL
lSX1PlM2bofwz1QtUjggf3t9NYum9h0HpZGJWcBJBWD1sVZjTqBZWMXZ+5yx1wY0
+OimjL4xSAO0vA5mhGidevW0ezHu0qecR5/BQr867UjD0IUH4a17EhGuhUBAlIZS
X36QvbSzOKx6ola4UbTLbYYUSbMXK5g1W4lt8C2DGmFxSjAYptQuBBhLdbzckUKu
HW3zI2n8RueERpGRW4EpiYePUzWmMVD/rWJ5xGyUZPQe0vvov0kYVbQHU+jWF9ex
+qmxVLguJWWCW+MkKTzNSukJzGqf3dRa+jkbyXkJYtPwo1MRiSI3mOiVhiTgKSjr
DZoy+190eX6ue64wtEv2Z1EI8rCqmvBfNElEI3EYNMmNr22nUOARQh6yC0mrpYC5
3KVMlVaTTboYMwBmJa61nzUtYlLYcAseTjWw3DczjAejQvNwSQCM2eLXLxszaWiG
cd26t9thbyTDa9DsPLdv0NyUHzPwrNc+zbZc1Z7BdUYzh+SQ00sKmx5kg9XbwoJJ
KfLO+A4DJHY0U1J+yI3GbXr0t9OXg2r6SRxLjuBG+edD7wse6gxusCZtbjaN5ENw
kzogawBvnOeW+vusIlwVvevfS31J2mLsD9L4Jr14lnFCbGpxjF42zPveiobU1eHw
6Vhu9PoRwU6MGmJPdP85r+yd8XZPF7XcssRmo+NZyfbSeDByM7RzF09/cDijHT4B
Q9Y2ksh2d+Jhd/Fn+z1KSn4Oi8w5PiyIqfrSVUSd9PnLs6gZ8o+nriYjxd2/Y/Wy
lftnbanjq7Y2+mqxKI2KHkQOHP/+dGm0wu+mabqeZD6mm2GOVEWqed9ucOQW1v1w
6Ig1DB6vI15fGE3H0nmbbIHAbqVXWw3+4RZ0ac9H2IQriTm4/DFZV9EX26+xzJ8K
KXFkoTViALVDtL0JSlfNJJ1eNdz59QQUmX7nfclB09ATP/w9IHErkb5F+6LnNFGM
mPNzQj+tXSyjJLyVNV1ZQ1NwPT/Ze3DYKYdRlmCqXQtJ2rgUC0HkI1OPTr4JHIvu
QXCNtmynm0X7w5OQ2t3jr59wKCMAH5LMMMU7HSTvx6ZzXn0icQ+ZSkQYMudMgIKY
wz0Dx6dDDw+TRymOPRREYTKLNslCJGtDsdaMnQiZePW4Z6h/XnyEzxbejFOk3qeg
bg9sGLEsJVqoBiQVBH0yaHM+5zEsvGKp14T2wAUVazkMVodNKxolLwf4wUbfxcvh
reweIVEGS59rvYwHVG9JR3zgA8EebFaKa6vAAKt3dHb/Zfjkjrmb4lsC5mPOW4N/
uvt6x3Xv1EyHklZxhxE/qGS0D+7/Mdy6eTIeflKeIXGR99CG5aXF40WCUKkIwziD
uf/vcL6vOprcCAUyXdwOnw6mS0Hzk3hnoa5SWCTGOlqxeSNlLJJ9Y4uQ7zrHBgAk
Q24NAiaDEydw2/4c1eED93RSfxNgSEtQWUiqVzGWSsy6nCCaNJ48Qs6Xfa6S1Wgm
Nd33BGbkwRW7PhGUbKNfYaXaBaIXSRrKUYqmBTXhd6nR98+yXS0+24Tn/zApAQ6e
gbZUdFEi9FswwTDHFdcyDhYrj+AevlY1rb9eZwTyfRdzQcsUgKTnLG0vj+ecF7kV
frKsPfBla8b1gfW5ZBHDqRN6vlZuQovkJtxHp2q573+wJIMb3p7B0cyeWeKuev6P
aeTRRL2LHAN5dA9zNnwRPWdv4By2fjzsgavHfz5O3do9zZaTP3ZF8DTSDRwxXmWW
6fGRqLstclD4y+ZRA1gcV+380gfAPFzc+bjKbQ+m9VgMyQEo71VD5STNInV9dcrz
cvU7mUMFDfcR8vIwAMCCfHsFMTFALG1bTw1eVCYXhlAUnfUCtLOzYo59zi/93kOy
VyATzSE9VnGGPTq6kfrxmvRaC3LCiyOUn7YjxE2URjbZ5LOJiQGpFsCsax4Pp5x0
WokZDvF8Sky8ZRblmVoZ7yili312/5ZYGnqzEhsC4bkganrnMyOs0j9MFQZyFgcS
cWQvGOCZYZppbET6hlg6JCxDQwN3Nhld8mtwka6utFMYovM+HKDpFsE/ykmu26eW
hox6Rgmc6wzvWutjoyCrwYz+R9XRwm/X61G6qA+FkHO2I+xRMqL4Ehn6p12fv2Yu
9+g91FTXj95x+dT6e0sg3M0SfLiIx3IwMWmWlGHphbmstzzO2okRJH/NL0nqhDQT
WlGsrXt/osY911ciRLVuOsNvD+RDWG04E6wLSV6zueBczyowGrQ5jphv/TNdTHwu
IJkek4oKyFUMeo3ECe9Y3iz4X7rResqNV7/Sj5jbPEE07Iqs5cRv8bLyR7TGUQoX
KfAlSv3hqeMISP8aYsbZTcqYqFeDzyXIDEh+BXRjWcEcoiaLeBcBXlBFIeQs/Co3
SAzrbeoYn4/aegwGVaJ6YySOyO/nyzCU3hbbs+z7VPL3D763F5qcSbga+9H8e/8B
j6LMFCq+nJv4rvmBb++2pwchi/U2/8QGyb/qgJ3PagKqXn6JUdUhqjmufFH+MSXd
QaFfE5YoZ5vjkuN+liUlKbouQo8o4rl2YMXdRDUv9OQGT5GKFfzOHCciSQzgzMwR
0gvPgFDTtkdE/SMohABWJhIWbfVbMPEMWqRehYNFzJqlhCGJ9Lph29jecTdmuTPy
1eddJ0VnyXmk//4LO2GXQvv2Bha/DIHbiu8zBlMRAk4Clysu+ir76gWRq1jaSQyi
hYbD5gP1+ioQWOuL7zetqcwAcFaV/6W7mPN0NX82wwp6TyOz8v6oPHZYsHJc/AMq
ktW6MzOvPSwWDe0Ju+lBYK7Wui7PCmqNIdBaVGg5CHvo3N7IHFn83eZiHl2uufNK
Tw10AN1U9tMghaChNcdW6UU5YfXagbbgpKIpLIQP+fyCk7HnMgPPxddfq9SC828c
UHU3hv3fVEKQRt3Txgo6bSFaCrShB1AsjD8dXG4XEKT88YbBO4aIsLOOgoeiK2G0
6Pvrdo+wzZqVZRZ3MUa6rVT07otumZpRk+7GBp6iJofWy5W+sYWw9xFcfCzEoR0j
5XRIeqXdVOWm6Ebw+lqKYjC3KQDKA5tqMRCEseYTYLfo8zBCT7le0NZ1g/V9w8FF
hQvPSRYWOg2EdF67Wz5kfMnr6PaaAX5hyat+hfplMlY/BmioFXLPAB4VQQfhRF7/
+sHZwkT6XDYaUlECU8HCV4ir1dyVrzLdO5WfMbMrPihX3WtJ4K9NMecygIgdxysl
K3MBwHe5caBxwaujw4lrXP36D7BZd3JhJwsY8m4NB0iIa1G0mlIAtbMrrrVCXPzn
omfFmqbdL0ylM9XoXscjsqT7dTwH3ilBQx1kLrzYNJyUFuFIqqZGAdYwLca5883H
knGsXwF89rs2Ph4YnaeA75iKw1Nh2vzX6/4qAPuqzHESxgQvpqmZwEMusW8u6hwW
p/5JFjS+PHbiq+UVKoX1E/JeY8IdY7DbOKbgcOGsA+joYV5JgU3yVnMalypgGqnR
YxCipmz0hcGmwldIef4Bs1PjOWNytgG/Ol49TU9QeVm/hxtWMxvCvAeSZPhI31ax
kLBLohCH7ULuB0xliGPGAgqWs+QTTl8Z1Bb0lM7U1B8s6U43LYP19SifXsAdNlJx
2QWd5Z67/E5lQXr9Q3jCPGPxUbO4eVhvt5+C3UIpj31d4rHuehz4g8npNVPgD1jG
KzBHiCYlxuUJ7Hd667AQVk+e2/575NaawtNJzgqmzoJ0SFqcGKnI20wE0zxoB7rh
ucvym6JlwtQL4OmCZF0qvHBhwXlYLqnUvaYhaObv08K2XNNYjPsPTsedCgWQIjf2
905P7fRdgohVOybEySQ7L3Y9a90eR0wDSXT2gZaz+nPUrwnupqpt8FDF4rkf/X+m
iurGX3AiRijoYkYx3aAkBC1riIZcdYintVkFmOPBKHX7wlyfx8eV+J+EnNYpkRl2
pJPR3pktCzFizA7BzBTt5JNCcJW1roatPsLvkqtmM1rraT3t4kc/OI8rf8bUv4Hn
BZ4R9lgjCVk08yROrQ6M8I+lHC04Gcka4d/Mfk5dubSVCK+8gI8dPEwJ+pciHGeP
odI9x8xdoc7UOZyufEihtwbOp4cKNxsjtlhXy2GtcrPA/a/Eeqb9nqutYOXIuBsg
j9Jq6aAep7ZIYg3pBdjBjeNVDlYKuL66KsXARlnGmGrQi3UFOg2VDzheQqfCcBAv
+qfes3MGKFulnCPmjswiw12BGe3vcaYrejPms49bSV42ZlB9a/YnlHGHb88Qjb08
pzzxe4jAo4xrHAa1dE46HRFluehHY0YfxLPKJy5G+vWWfI1S9lnMbTwPW9G00waE
lje30zYs5cq6XBEFEkWhFQ/hGL89s1cGmwFGE4ojRDLAUvJSHtK8TWsiOZgStjsz
DB9GZ3aOl6JFVS2aHD9ERyVKPeUInjkHEeGTNHTJ20iJOF4yBjt1175rm5Xpb6+U
RTfMOa8hsQI/hR3X5iRJ6LLPB2ftjopB/9kgws/ScimNxocVHkCcYX5mXatvQADC
QWuYgftDg6J07qGK5aLXB4xUu1srJ78DEZWw/dX5PPCpxSEpGzny7T78Msf31oF/
snjWpCNYJtj/Q/2CxZtSTPtXyBNkHb2vjWJeQmmuNC1V/Kh4WQcDO9toGhKpolPo
FAZ7NQUH4NzUitxIJzpmLg2Lsdf6tA3SdyFQqhnNDLy70V4PlBQ3RmXDqW6WzIbz
LOw5DAVMD5jeWGIsqNMxdFp3rg3bqqz9BCUDbnSZDEmjofYOyev6W/wazQc7D9DG
7QZ2KuiUqZqqOuq1CJbDYZxIcWkK/elyFRTi+R+z20Nu9IRp3jb028ocelmhPHyH
pu2HVnS5g3WBEPLmZSx0uplmyMee8gbnEOLq7XWhSi8DjLzNZL5ht2oHCnIEGlmc
Um5FSfMDWHJvx2L04JZE4h44vfb/jTEEqewpr0uo+rrCJh78mb+RcZD1ViCDggoI
PJl7KEnoHh3EyDWyN5J4adVFMx68T8fc/A0QUJr22+Mtcu+2XxJjgEzYTeypgukW
EiWhJPIc0dXyJM2hJGwVdsoxYf+DQ0r6NT+diqc8O1lzSQKEBE/91fvNWbCqwNh3
Hvy7+0NfpE9w6ASuaSvSbbU+aH7eD9TY+eSfxcrsoc/lTsf5gmXVg4bp2AZxco7X
m4NUpPuOleEQBL3XRt7TH5N6rRhw8lyLAWOSaVxp6WyC00OmjtXSLwsV5fa9MoaW
sOj2rii/A6G0bns4UVFP0e4nJer1kPjf2tc/HU/e0oP51m3DBQrKPOF2XHGuGwLO
yNGTJpQSdS+BlbD6464qVZEMSg+acaVDjdIpCzGu0Jdvdp2/x41pu0guiwjjtMMZ
66qrgpFXHfgXutoUggY2jm3bcLmw8FlstNmRRDUqueaiG/80uNRTqlSbNmqwGWyB
abhHsaiaH78knzO8ZJKCbCsb0jbhc3kV0zoouLOYGcpRowkDKizPNfuB+oFA1l2I
UcAZ3QOtLVJaQ8XIycL0TjM9fjb3Z5rvuOoA79GPQDbzM933H0yfuNEjAvRfA04z
hbFRYB8YH7LsoYNlnu/gtyQnUtbR0I4Msdpn0O8QAo1LGIOxX+Cvgzrq0YZLa5yt
O0SlWxaXb036sYoL/G69KA8atDxwdkBbABfuMp9fve92dajrJamHCMrajIxXUPgj
et1aHGqMsGY5ecFndexAk/jr327hNJJniWT5dN85wTf2w+V0w2TIOdQcXc//pP30
1DojjVBl9Da1Pj4FrJVb6aSo3WEGC2ktYQ0PhniKXH3p80cdF9/2lSBF17Vrf5xq
Fxm2viK8F4FAI4dFzf2ai8k5A8eQU8m2Hejx6dbs0/yHZflzo82AFNw5PztKqTr0
NTMbGZMLr6/6+n12cj0t68kSk1+FQHDfvgS8cb0S39YuCpgy2FQBgUhfzxUPaxba
8eu1nIJaBnbWm55zNuS29DwFLyKoi+RecQ4rYEVpzoab0WNXLxOVQ4ti5syfc81r
MZ/+R0dt0LxJyssw2f46wwMjJvQ2H6oAf25zmSVZT+S6zRswPug6nfdmVjooX+U2
eIfKjkcUrS8xf+RosLsR+ynpjiD0Pt1c0CJQMV3XqNQPiwXI3YvXwwI7j6mInLi4
tGRNpe9xixZ9qPUUWScPNQIOGwIuk+oNoghbaDPjWeZeYJaugMAtpB4xG0A/sPe4
1AjLEydvteJUmt5TFRAXcIgLawd5fU8nwssQ9ULtJQ5XO1cXmZPKiiBUEqqTKVxj
zE1kF0nLMOfcOSdOSseVqxN1wWDuHpHU1ScF4v18gkO7EtHgIF1EnSbFokiawz4e
1YpPw6wUvaZ8E9uOM1QG5LBigtW4EEkdj1CK5cH8c5we/kxLT4Dkoeny1GqVTpNE
o4zfoVI9mGPXrwY33G1xkwEh96LFRACWTG6v6MCMoA8lfwWMBkKDC9FE7ehJoYVB
bFmNkLvYOpq+sRY+RDHb9yZ9oE8vcvuUr1p3cNLerDVpRaL4aPd66av440aOe2RK
jx5v8eI9cu5A7IIiKgJavqbT5T0+pl4oy65JpTvEKyeGSx8z6tgJQFKiJEd+h+RI
8vpvJscdW2HD+jXSXFuYn5K+GLZD3JG8+JbmtFdvAh5l3H87tw2JroNHgC8eNOwB
k5UdXFfZVpmnnDul3kR5f2VrX13KHiiL65r61fWrXovy71yd4UcDmMFdRbUvC6ed
0Pck6VdJpp5NzsUq3ig1FrXDo+/Ol0VojeD9FFdpb1ArMzHMZmujK4O0J8d4m/dX
b6zmXp8vGMbNlbJcwkwROcItqHrfsIxiv0KLERfqNRVlq1d3XVTLETstmSlDwx2V
Zt/oCyFfxA6ywv/9U/jBTIQ0F1BwWacsp3m04g4VaHgWpr/q19Tr1LcBHBb0TbHf
IjrFBakbepdD9ttjGaherWMTuyEYllI4Mx9ZgIhmgA8SwG9H2mimQrnvKNn1s83R
lKYmsNa2ou+tsEk8rprN3IAgR6tUicmS84VT1saIlYJN6QYWQrLY9EzN9WqBFcCL
kziFUIZnf1ptxGrOCQs7n4WTqih9AEnVjiCSiiXsbztAHO4zWn3j7VImpYMhwLqT
ZEheBoIadcajKYwGXyxMzL6COd1a086vaV1lDmQGAVfZ9CVrvskqNtZ22sazsugn
4j4vRotmoQjDxOYhH6qrzkNIyQl+Al9jIVNYa7cujNhSqgjEB+Ipj9eLGGLunQpy
sJ+0dhqtmD1hss77q7fOC164ptAF9vKew998OzHFYHm+DOzNmw+9Tea+DW8xAEY2
Jr88gIbrbBCDnbaLgi1vhiYPJGU80RA6UJ3PdUgr8Lch3b3NgAKJ6FPH9QnLy3l+
dgg88SwBeAP0cdonsEGrfrcl1QGF3CJx/cJMWc6uA5hbcIvcBMiX+Fe3rK5LIPg3
xEifXJgPlhZREPqAs/9Y8SQenQ/eFHBI17yOEdma588OblGBMGxq0GyuEFvRiVcl
Ej8ptCBWOXdC0akTNESc2K7CebktzviymhQkKdJaxmfpWIn8HPl0sFykujTWQ87R
o74ySrFDqfwR47PRp3ju7YAHhQ7hcp5AoixEnCHRJPupgocYGFTsuOfO5SZvUCOj
iV1QbdNj7ZBlN6SGoHZ79bwAHWmm+rGDsFdZI8Oegj6jBZemkfWXdecDEfanvbaz
DkWLosApgeKlxdIC9g5AKQCVzYC/hkc8OFVxeK1sOXGdAafux13noCMRiEvjyn4c
BSKEyoisXGLVpwASpQKM/fXFSc3T10tae3UD0Gtszx3vpcyE7v0+Qn19VoyrtdlV
5IqsKz1oToZXkQbJobGfUwLi7gF7UsOKgD8aA31Li9p00gdbJibeTrkPAkVyWv0J
oEXybcHw7oUTwGgFH8+R6pTC1f9bTm1GMxYrMAlJVNCJcVGcU+OjyuVpiilkomOR
wAQNCLEMlfr2Xc7HDflG2M80WmgW32bdE3Dn1loP7tuK2PSyljCA+wBvbiocBRVD
Mpwkg4kX0s7nbRfRuSckjh6fMr3No9H81jegWbaHSYvLumUJWwgzmOJ7Vut9Xdk8
Q+A/X3idgf1g0yuHtI9C7h1iamogmWWhlMeVk7yiXWJroOUP7FWdhzSIuMTZ1you
0aiyIxwkZDueXohmOhMjy+AuQvymjoIJVHJSXYHMHiqPQVIM7mRzkKgADl0XXO58
NgBUm2hpq1rcTAQTLOx4XWc9R5mDXsweyaUXGxyj8AJMP0e/DTptkXVPzjWQnSD4
mC3HcqJV7GalEnPmcgLhJSbZXZ+CAir4AZgUW/wVXW5enNgqczaZn9vdxwwVwXEC
ApuSvKER1b9fTR/Oa96zS5mdIyfoEGsQE+/Atb7TTc8KBI4jLkK9BDmrUSwXNf2M
jVG3Zk6NdkOywrGyCxe9TBIGeW8nPiDERchKWb1vUpAZjfbzGxMgjmR43g04wXY2
PsapCAuL6UilYNQC1tt+QI+IoCtNGT2WVBiwrbIFVZMKW1OlHzp+58gVY0n8WrN7
a8sDXyxUT9xelGF0niMz4/7Uk6JnDnQ01mlvOMiWkrBbEAfjnb9MFpy+b8IepJku
pK3zQbNzdEOt57a30RSxucMyXHVK1lQKG91YCMLoNwBPWRdELmS6xl5C1wx8CMsR
ZgGtqkTMbpaAN87e/OoAftb0gynPgtdMwZgYaEEyMgX1pMoN+Kz6L9ApBkc9bDYB
Av0heoZXeA3RWg9I37aqPLZ7ejsYknJgHNydq8wTfhMkTpUtCKeevpUWEMv0DtLv
RFc7ahZpA0FS5nYHtAHd26CN4OUiOLikz74SK/XIfISheAg7TxgsgjEa9qjw2/zt
gNUpLATBOpm1PY6wBIMp5jp5/E07JvdYo18LEpIrjlkloIbGMSh1M+eg4vjY7fzv
1z0dLuEQLQGg6kUppe6cR1GV5FmeXkYtXut+iVlhBRIJ0lm98c4nBudCMrN11hQw
ttWhGaYds8cCkvuWWcNi+dS54n7vWEI89gRBHgT/WW8kUNj/KZAhCvuyS8pEUGMR
YbtUrBfGRDOZOZ1PLXSrIYGddCFbf6ojJDkQNVUkmMeS+suShH3H5uhaEvsZcp8Q
Ffx9kY9DDfRy80ObD0MTmDHQLwT0aqKUBExHhWc+xHK9C0oUM5v2Acah1s34MslV
+EZ3a63lZARaUHsXY0hZ6SCBC2zhEAd7+XjgfQPhIwkfjdZZKC+E0mcOQsnFSE4H
roQ/SbpORRzaep/V0OkSEU5es5qCPcUvT9mQe6T9UFjrlxCUbJdq0oB1Gt49y/K+
OSn2jnqyRFFCxhSAmiebFnwf1mOklPbRTJsAl8uoEAM6IthG2HdMxRWrIvFp6Wdm
0kYV4Eq+QQvu7dMj1eUUw/G/9uyIMuNupP0nDAoTEOwSgF7O+toN9jyi0WFQsZOl
VEAUfDwyt6fpaBil/SNqAWESd6jyZ/n7CbrYeZLmNaapxwoYDKHfjBJRXEmF8Kjj
f+duSZ1ZxL4s4wd/LnRRG9LqHNrl+tehda4s3q4Dc/kfiex9stS/X5wB7mmoWEmm
3ekTiITdhg0Ysf1ADbldeNsxp52B1YFncYuruqX/jdrSta9Z35TBTzLJ4S34nc7w
W87qtQTGWoqOTYXGfJhSMMzymr6i46gVfSNBk/Dg6TX5NhFRhfm9UEhsW6B6z04o
Ojcv+7HOnMPNgiLPtP9c1NoxQIlbSDQnaAiREY0yogRsuIHBLqS1dH1cv7+ft1oS
6r24OLjHW/mRq1kLwDNsG5ZbeOq5dB85lcAE6ugGWYz65yWoCub5e2fR2YO8rcK3
u25BSFxdaexy9bbEoAbls7f3Q0PhD6/QXdvHjJUVJHQkx3CTIoDhYR5+brhvA+0I
HHTMCahwb+Rdg2KvR0pv6KpEHeUrasbRUSYUbj4Yn8XPN69lWL3GaRfn9JjgnyFc
mbdhldIK27IPbV+e3iJmekbRC8zwgLOU5wKgxH/ALO0DgDH6YXTNFw6gCdMRYchP
ffQTy0TjTWsJR7o6KLMPk2EWNU6tLpGdlysgTvXJ7OEve1kgdOvzWNwoK9vagfmv
aeiS2V7VmyBigREZrCH0qguE+lTnzdgi0LIKWDXwGICyLhBK2OHTTivskMdtEEXa
leDt5BtOr8tDFBQry0jmGiJ6tQ6B+MFVWkEzLMtxTTvD2G/RAusINOOd+kdlzOFz
yBTXoLbx33uUVhJJZbWvw/lO57Ny79Y6lSXjHy/wrzP8yJcAvWOUC3lPjGWfy88S
OoOVP28bwqxNajYilrirqBhkMyfSQh9idWyYZwx7jtba6vaBbOHJFL4Y4LXnZHTQ
lEP+BEaoofx8JuVuGDyh2++b5/CiOxcKKMAR+Gn3QfIqeIDlLl5Crb5ripkKTYGx
S/fNPaEsF6L/fhwcMSk/CwXobBpU37pWVuWd1ByYhA21Lca+k8fiPEdc6VEzpdpb
OioLy2Mn9xUGBiG1azsS0nY6VfEKvnAvt2AQLzSkGZvEQ8LFDZgq98mO8d4yS5/6
s8Os6cJXh27TkPDJojcoDakwoYgbQ17qe2osJ7Kcwl0925KdllxqutOC64cSwcvT
qwIFG/Sv+R7tNVXNhajCp1ATSkiSR9+o1ouC2Q9iuRZtqUC7F3Z9XGHqUoi9Fu22
IkbNfyfzKdrfG/kzuTgBUUnlEqPww9FjHGgGrMNUuwa4BdtcL5zgrM34gmFp053J
kPvg7VoTE2rpbXjIA4mbkA60oRpLKq8VIQpVZoYnBvN8zz0jieBd4osi6o1RE6yq
WHiP5h9fmlWFyhMXEgz2gATiIxH7LChcGNyNSYL0AtVmwhfSuZA4bJNIo5BmKnM6
0ERigXbbf+dqTzA4HOArZjdbCkKjOsG3KWbLkobXl3+xI0DnzINQu9J5/ioupRdR
Ex8LEBvx4+DJjpsuGQEwQ4wkZ6Bzt/LzGEgxi8rb47R2mQrjpbuPbwmtihASfYOd
n0pevByjXOLWRE30k8dzyE+1CR/6J1ThhnG1GVsy5HH5khtU0va4OQMwGE1kZwCt
RBLaak7KwI+8yhY/ORa0AEOZahRtqEg4rAmQscWF4w7FGg6V/SO73eWCxx7sF25s
q8UnrrORObgZziHMSFI27CshRioyWtzvt7qcS0znDUbM8gzREX+XlFK2psKRsBRj
I7ebrfHJoX5UprxKfbPumG2s2eoumePSHuSrEjOLNE+qIg7u4Bf+WZCBJlNSXA71
29BRRHB4Bu40fJT2C5J4WO3O3b8vgCqy6T4m7Vkt5FE8sK68NHzRuATZXCcA5L8E
R3ZPfXepgwckUHhxWzq7wZu221eXAK+IlsFB/wQdTT2tf+w9I+J3Px9ijr9NUsFk
6J4k40wrLUnjj3xm0CvfVP97NlIyNm/nHKw8VmzGlrCtnkOxEMLbfC8hqwOwjFi8
p29K/xdgmw0oo7yUql42/gmgSStoBihFdRULI/KZH6qKjkmcb2tqlyUnDRLwDZX5
HckJGAsNfVG0u9GqFfo81t0/fmqD43pwsDn8vWCAiSpnhwt2V1Ms6B1uzWfgSDK4
lsvEoUDScyrNEwTGHeIqhBO17Swwlx7/gEVixrRD7MegIRcbguItl/A/binZrnSd
Lf1TSe2YGpjNOjCOnSj7Fun9ZS3vQyk5TSZdzd2GtJFiXAe09ypus7gl3seNqTT0
5gQj055ckc3dxEzjlGABPVOOxQSzJWmXrXCAOKAVBXIMX5IPtzIpcdKqCCK+2bSC
+glYwDFf6Yp7f3G21rnxtOWpmIeYBZiNz4OTMAQqrpsI9NFgojpAEocVKP0e8UYZ
bEfdWwP0+icqJ9lrtDmitaSLUawcvDKNHCJH05wqmb8JdTLgvwr9SfZXb0gnt3A2
DuusnEVek3kBxk2AUxIERJ+Wbv0cwBHJLEc6KTdcctpU102gyl0VrDGXZMb5P22d
vjE36WJPMnBEItRfCtScfSOE/BKRTX256F2jnd/4VmcoSp3FwyhyPqfeZKL+QsyN
YKEee4601HoEDE/vKr5p8qW142/t7ACUaqEj1DZHxKxQzTxMtQ8hucu4MEdL2B1E
t7BPRSJyu/Xoy0lUe6oPsFJFXEOcKaSkVZi3ivh8C064SZpzKNUm07B+DuqSP2U9
paU9gbmwvyxIIyt8BK6BVyUjeDmy0HFfJCOJwc16MuO7Bq5S2cl9mSJy5LkITgyL
95MHyvqhoyI+kASwkv19FyG5AbTBlTHBBhp+1UpZD7vdrn1EFqnK46ht+GWuK96O
bHVr9nDZT9W7NFnMtTCgX8VGhP9deM0l+7OmfUxrPBSy605qtDDgDN6wi8MUYTBq
GMDc2VVXqMK2bUYmMCPxkdEXsHZTboXA3jhzf3XACeC4fkFKN7OnUir98nDijH4N
Hn/SlDrhpqcg0EeuISB4+YG4I9myXDsD7lid+x7aKvepQnpd0mODmHa9YsJUa1gR
Cmah2Lav5xJkM/h680BFRtEre7C0uRdeQTE6kJoS7dSMs9oqPN5un45q5fJf6PAc
POfCovdiiQ4s9UZDChgvFCjDiR9mpL0hQyh18TINqPfecy+V3eibpkdZjJmyrqbd
9PSkVzmt0avrobz/J/U5Yya6o9Ee0VQlfi8N95TMDZSOqdELp8YIqI1F1t9beAal
cHeeAoT7YOxfrIFsMUhLk8ibTQigD4e3tA0mbI1mUwhI6F1X2gCwRRGbZ61j3+gA
XQRUqJS6wBgC3UkYeRP6cGRvrvOBB1pfsyWwqUVPuj29UYlJ0yK3PHbpTEdP3Uuq
VLUTaeMcyWb1ituNccik1wfSGtJXzxfUWdBAAsDgzTBdYnrmybH3qk3+0VsgPUyr
uZwB8FmuBUY3iyjO5u1Q9XGftbB+xQA9+pqRhsSjumjdsd8LDTg166MZ9gvredhz
21fE/NxoRzlbXx0/6YTu64NgoRd2M4BQPJ3ThYlapn11/SIA6/hZOowwV2qhBwWz
Y44puFj5VYgwqSo9nraYBjAiP06hC9owk0Hycrpn6y5XtssmJd8eMYlJCA18LO69
bCzQZ6Ng73o13LpHPstn5O9O6NFs060YCEM/mYW36CLFYsMb+XikM6v4YDFhruqY
FzuT2OdGGtSaLv89/Ra/53C7n80gyjwokqAWFf0lUefZRBwSa3VktXQQAKUBIZab
uzTJJq6PcCLIAhDsjrBfKX4e9i4q97SuOvvCnw1KkKMUxQcevRX3FWX4YCrjqfZu
rGXB77FcyJuo+/A7IeCow1z2CEQn+GCAF2cJE+s3EzuicyMhtyG9ZxxZh/LEvGCz
leeVS4NtJtPHED8J/0Cpv7HDGmhD5OLTJe68F9105h5VymMae0bA2JMZYWvBGVEB
aP36cKNe+i80XVQQByDr6+GVNIk/KSejgr+HbibE2pISXGHYMAKSLxvYSMdcK2jE
WjrPpYaIdNpIYMUEGO+GwUDcLqdPWyOANsvaRLcdwC40vWLYAnUfqoIIBJ5bA5QR
lpEy7rK+Excz5DqrYmgH3yGtEPhpWacKAhgYGP9uj/DsneBvIVYzPB6A3XRg7MPv
C6Tc1aGL+uL6GBf7NZ6GdsyC1FDfsLsEF8irizYcrrERfsZw4nX3FEXf5wIMQPRE
lRXSQZuH9Y2opj28JJudTY85jWkEJaCUk0ybTswj4soGsodGba7s3b5zTnkwsZ9i
fqbVDKjc7X7h8grh3mufxaOX/xqcI6QiSvIjacmagMwhmVMqL6YLN8u/xMV6/qVm
qKwe2tewA8LyM8M00s8XYR+Ygh5Sy7W6IEBnuF1E2eMgpaqfKzOeq18LXc4eiZYk
8+/ONa164AfggQcwmIM+oQ3tC/qn613pZvrevf2lqCmVgRU3AS1ZKSiRdRdhA1F/
PsUEG4o5PgUkYhLnzt6a8kdGb6+V4DJq7Fi4LNxwWz0vSA9S7LnEPfHm0HenQjXX
QXvWaqApfv1TGzutz7knJzakBgLqzYA4p9RUU0QzYt3Rz1BwtPTVMJ89+6olDQX3
bwkd0NFYkdJEVUSKcG38hUheELerfqO7u/lA93w9yxmvlGrDvJieRrG6HjcQIcv5
Lw4iHqy6+y1nK/b8dJW879k6UJx+nXAU8raWtf8PxvjFxQE6EU349SYBE+RSH3Y1
v9jhUGuUciW9g/d1ENcDGUxP8wArvwW2agt51mk6k/F2Sm3P1WEqkFE82+Po+Cnp
4LZnA4RFcK2ZnUsmggz5+f9Utdfdv12Sg33sV5GMbgNCBomYY2dUuL1s1GXgX9AH
iekELpSlrCQV2y2L54B5P2CKScQOTUfNoPk2waVm0vhb+bs2tf8Ad00OIZMSF6oQ
eYSOk43ew9fR2uB2o3iQJxZUV6PyiYM7W/8TeMXyqlw4PyxQplooisTyTdieh9MB
Mup6xze/vJRuuKf6OBiTJxTZoDIJlsKGiFgJzfWvSWNOqHMdEaYtGz2O7QF19KXw
CpgOQuBJoKfI3G7iHpBLBayX4byXjP2i0tGu6rIE4cXKhsfNN9n10fakSOARkoaX
o3vvcqeQipKwnIGM1UfFOaZdqPY+24CWlDggKl+R7J5M3HGYoeFzxwbuHjCZpbho
jfnKlINqWmzmvR7GBr0i/JpXEMJN6b7JReQZrvMNoF/j1I6CigABL9P+7owSv0+y
ASOeX6YXHDgcmqvIDOXCtWqr921vQV8YmhU+MyhwMYjPT8gLmzPHLQUzL0zLwyr/
Gh8llKkTkDfXtoZTcJGTpkr2VfR9fqX5EntRjzvdUUbAELMQLUT7m0a4xkWF4+6K
W8POeNJ4M6KyrMYxP1VNlq5YDuQXd/sjgRoVb+YrvfTnCiG084njtZ6At/LLkpAK
TdkpWrnvNXswhIYQavGaxKEehptVnhH3/ICTygLNazYv7jDc5lJQcZesc9NQh6Ix
d6rUrupzwGybjD7t82gUeQBXfIMNj5GUiiuUF6rftlfHmi4VQ9AxjBmQT0r++bMi
2Wh7QEskqE2LcNTm4ZDCREN7b6xVH7zjkPEOQu+qQsKACWh3XxtvYzbNnLT2i/1d
afECild9AsLz/caeudT0SDbVhNF/AtsHWghzF2FcifhPRvEuT+QbuFvJDfXjYBzm
1x8hQoI5ksI8OMMVVH7cLCLj+w7RSdTqHVwpP0RoMIc6HTEY5/1MZk8y78ENpSUA
Ne+g01o27YZWNyLK35HiMoHNMlQ8peKkEGP7BZUrakX/Cczk/GevEq/nyAkfBkbU
yRGrwoQHnEA9MDhGwh0uHyDa63SLT6sU+9kFCtQRFck8aeHgrvhZ/LBDsrYg+R8L
N4aKYIJEd5fbuG3oDINJH3EdWeSMIkQlN6lMNxI71XGM2KFDc6xLMFJcHYhEukp6
hiTxzudwszuudkcTM0QzItLfjiZLxqq5m/jiGfTSiaxFUNxBGfBfWRTxDYRTTGf0
NafQNYaA9oATINdNDUZFDsjgLIb8QxJXxxHPZQ4JHOI8/tFIvF5ZYg/joOXwMSHd
3cJzUgYJSNppDNWeapcDnrBpW9OrAXPjtYI714aSgaWPbIXLnZBYBsvBEt6utACY
AiZmADiIbxDDnI/DMuLazNqb2HxheTrp3c0bWsuuI6+R7IeWLCvJHO43cz/VZeeU
Z3uS/GYwXcQqaTab/tD4VjcpYKxMOUH2CGXph6RLMzK9fPqF847Lr+F9WKyhFQcW
IiV+ljy1R9ReR6Twf0/NTDUiFejVuVZpRs/BEGxdQ3yIpwNA+hsjLQpnQMZEh1Vi
uIB8xqYwm09EO65SveBtmR1NlhdrDizMPhMXbu0U+NEDwxmuSiZVHD1QVai3S9rF
ffcWEi7ghzrvPwGOeSnxC3hTzgcd6YKHvVYAZuTvUKV0OmMjWZbAXIwJBX7nhLwI
8qpv6X1KtTs3CToruWBJDkwlolcfmyLM+AdgwSNk4nGgBF/E/xsraOT+cp+R04Bh
vdCIKDUJIw1fwAvOI8tlFXL1eYEOgsNfMV6Xo6R9tTfq6kfZdRI6R1v02PF/x4e5
ACe0ZIyYZJe4fNG+cA1k1c9Nxxx57AbZes1mD0PsOtbllibdlZ89KrPoKqtXLcDn
HU5D8kg/w5ZlEbjJ2FgQJpbczwqCu9zjKkYUWDUJsYU+RmXv0qeMIiUh0Q/TP3PZ
ZNlxsG+IH5hwAvBZ35sSJyrwxjhCpKLF83EIC0UWCQeJx84mM4yMu13PNw9usHJB
0vdyLxFuCwBawIv0tPxOpa8D3YsuA0PEWfW3GtHTjX2q4y17lDg+RsxK8qvvEvlo
IF8MDspLQG5ircJ//bj9xECNa6hHw+0kiPgx4pYMYusyB19jJzJXIz3r1USZQ0wg
xlwZOE+ZzNCqs29RGw9jeqLaHJmXYNA7nMNFkbBsYwe26SMDHkVMTc5nqsr3Q/Xv
hJnAZSBEOHmqHs7fycyz+Aw0/R8N+yPbTBiwkGfqYnYIlQKc1atnCMoDuji0tHae
ln+zJo6sHaJbpqog2012XP+aBNE1WSqh51LiTyjiCOicecIJMr2dil7eMs45iFn3
Q8hDzLW/9aTu1wttbZfywYGfV8C0hCXO1g0X8YFDtJC3PcBBFT4ciO1j914YnGYV
TT1hDgRqSwYRxO/Q/A7D78yfSRYDwrxDF9rPYoGk7Fw8cUkDahYxXq+TZt+KyRhd
57HeG8fhPVBg5tqTHQzslYzoXyKXt4iELco5xUUbSb5RXnBbNWkrQl38XLoSrT7Y
lmQD3mpNrMIwQsUqLtD08W+CxYFFfdg88cnO6BB9DN0O23xom3QbIyUey4yJLE4Z
lShh94ovbmOW+N+V28DlGr+OhofaStEZjyjb9GYcElC7V+1rzZl1dTkM/owwUYe5
aB0i8RX6za8NmCJ6NvrcJhgRj4u0D6G0gPXDvkaMw+3y1mFLii0oj4XWlQlPle1R
Ofe3rbnwiKSEKO6NH400fzNb2n514qPodgOqEYddEHuNYO38LczFME6zFDouqExr
neCK5/JaQuIJp3xTaZviQEuVf+EJ+Mr+MihOox6O7TbY303FKohISR3nDqbMwViQ
NyLCtymRn6R3cDP9HD/8ctXPTlsF9gIOGxt1pRU+3Pg97BepWOu+X0HEy3VPagzf
ghOSGpNRNhRDfkUhs6MiGWgPBXFrieox2xddCJIRfCAG9R+8nBUB3qd2YW6avKvm
Pnm0GTGm/hT077aR8riUCAOydDE/r8KWAHixruBOTjcL+8mhYPU1Xooqg6nQiM/j
+xOtfiW6oYU/cesKO3ltG3B3TBZuBboTgea7CwRHy5CuAEtEC86QdBeYBUhpqFUa
mD5tcdWAZjCXlKJTa/+NNG1UXvciRsLvAWJJIAuR/zM7lgJ+W+YXDWjuPSsExwV0
JhgwqkWRuADhWxuNDFIccYsAqCZj+GnWLrlvodukwkq0+hAi2sgobEIwAzPiqUrq
KluwxHX6vRJKFAN9AUkFINwCaVj4Vf5z2NrqZFCQ0g3F1ID2M8NcwPScJkOjCA/V
o31UA6+sr4y5LaVNfs+5sHeta0gfIiQov8J6E4rZqg0lrK5s4MFwVfa7G2LxL7tT
Br9Tp9B0Toy7DJSejbvOuv5xum5Habck4wfAISeHe1cTQEMsUK8uyT6CjKoOWvm5
Bw18Jjs5/NlYx9k+B7kUbUWoPzQeW8IFrQhU31q8ZlATPv+VCkh6Hb6rSjj3vwdV
YLUVU1APMqayvDVgBLqULxbSh1g9e0B7HZw2UOwEP/gSwaBrP4cvTYibYlN+NauW
cOcMjioqSoyeHLehTOGbRIzWCXZKxFi+R/mG13MpskqVe4k2ux022hplaD+GI+m3
m8x52BmOgC/VcLTpb9bxhFXsqZW2w/61QIBHzvX33BqBxm/ynXHYArmfH5B8LhO2
8nheeMFIVKWyYPnclaE+lG99mvXgQ8Mzlf5KQTgO5OguES9Ja5/gzdoZ89zdBH/H
9gnvRSIiOtH3ocaAkV3PebR6q+PwaBb1VDiL4EAP8h8/vSJnJuipUD1ZeYWcQWBl
K02rTQlgmKg+mt2fYXGYCN6Er77HMv47gppaBWTplazjlyd1DyMlnDqrxRDXB5a8
rlg87i3LoMczl0FEJrBgQ6vbeLKkI30lFS+nH4vlvGHzOKQqIkeAwS/BXBn31axi
pK3AaBSuVaAbwzNsSVlcwNEFlH99ymdLG5eYbsJzM8Cs369uAFNMAPwPkZQ7SoRC
ccZzlDx+HvdHnmscT+8fT8Mf+vCtH+08GIqM+317pCYZj3KzM7+fWykzCC1UHVO+
rFWWS7Ifb5mXS9Bu28VwaU88P65a4HxmuQZstMsugDlJ5KKQZdyZKECxQY6tApQZ
bGmVyXzN+JVMWA6FoVa2yzvjYUwGSZ6z3EjbXUVRW6l0Ti/hn9AH/crGm5w4tDbj
Zya1rww3Eza8yfigQK/AxMjD23qqnqiKqrQVUoZkVmBvAu5rkPt0gATgmofOP+kN
/QcSR+aIP5r8TUmyo0DQuNzEMRTLbnACUyO15EkyS83zxq3aVyaN+7EzX6j8rZMN
NM+ZO63FuvEeWRn5iY5h4c/1gxP2rviQzHSpj3nBYxxZcC2oio27f3K3NBRlnuLe
Xgv4PjVGhRIJ6YNuun5XDNgn9jJiwZrOAPEhOH5EDIkSC804ByjH1r+I0jnI/i0z
dlTuua7NbZ8Hykp23vV7HYZJV8VlyvMjakjBHMo/yNPx+B1GBkQRX+JfbmSB5d1F
gqnoY805t/CRaU1mv7/5RJQ9sCc6gzD7NVR8oj/TfnRAVX/50u387hCwkYYjznJr
UdsglJlVm7G2Jh9D54OL6UV1og99mAXuaoFU/W2IXdVMJyKrogKJvBAB0gt/miSz
VYFDXKAQIQTx0F+WjsSkGACgaFm8jn6eNgqiEtbK0cslhJrkT4SmsH5qZELBGHln
1Rm/n74nKZP28QRXxLUF8WLw5vt9x7gIbBMgsjLiQkeeZqu8AB4fkHsRIL6awzYu
iZ6Ymh774AErvIm8QBiu3XbYQPzixZOOxNwD/CQxQmYF1np9PbTbEtciZJ7npymf
bh5NyjM2VzEtD47Un96DN8uDHKSIBa4bM0oeENGvTeGEObBPamKbKyD5u5MgTXjJ
JauM2tB2zCU0iFbIOBcFEfTAXuSqwQdwMW2gcjgI5OXNpaOlM2zbAv3p5sjPPlMK
alB7Q5f+l489ZpePdEiyjG8/Y6L0h109FWW+tSv0COxrCx4yHJMbXy9DmHeqyc0g
rrdR2puNrerdQ66A84UpjaucPPyeZJccD4YOeuRHZB64hKQ9/YCZfMQndw3Dk0NL
Lofc+MRI+ZYlhYL5YsBuCAyF3Xria4XCsXoqHVI5VqDSqxqt1yE0/4sxZ+XLFdLF
EqOCQHlzrkKoJvd32AEfsWQhyQj6gdojERDYXDHLqcmiOBVj70evbFVacj76rwDX
kB3ZAVtGFBDml1X8c1eN29cjfDznrBaJ5L9ong/qRn0jtrsQqEkS4hOZLD5Y1vj6
WK0ENzYTK9GF5iY3cKIS2mhXE3JED4PBFG+6G2Eq7EjEKxliTngopVxGAfLNl55J
vbgyhpPQmX0jRA9a4wNwL1+n899KDowEFJcg1gkT/B8xAX1siA9GebDmxw2Vx/71
WLnh1UN3HveVV9S5crHWdqJ74tHoAS0W9ZRN5Hj56KqQpcCsU75qBSsVKnTibmDK
IZRojxAHN6ZFXCo+aUI2uGzjB6Id8A+Kdpq4UGpvnGGutz+/oT9AcqQO9w1GAIeb
RJMMrgjfI3X4Xcs1amPcZ1Y/NKSipnu6y8OgopvPo4BlJPU/nGe9La9jIed7X2Rk
aq8opwnu454pk7rMYS8wDuVOQoYMXwo01n+YaV5AwFxdNRqOG54ocX0FlFskV6E+
J3z87Q85PZhU2bIaMXMJk+G/FPdSSPRyjDrrQQK/wfT+E5wVcV2lS8gq5y+tm+jH
3mn5L7oe3ZLmR7Ghf4LT79VUY8gfvmHQb/p91/KXcOHRhAKmhoUwzBupazeyZr32
cR0qilpe2wujMak8pYxobp3KXBH8nHIsOpr5J/O3zp8uiEplo7aw27plKKQq1FE/
9fbizuGDeKdne7l8mjQl2T+0Emw61Mv9BZXWclYCnFCAchkVAtwC+SEmgNRVjTTW
/Dzqi7PWB01xmXdGgM3moogaJ2sNkCgGm67ur98Q6nBiTayztNrph2x9TC20n0BK
Vd/oKmdUkfiRSjbU4U/CHwg7EIeI6Vg0Jp8mpFJCZiooPfEqy46whBd26eChx53z
5xxbP2az+fSiswYhJpi0SwWppsDkFs4A13GZ/V54btSmk8xgjbpxxm4iDL+NxvKT
+IBIILTQHcO6QsAmrUOaR4BaevPSQ8aYJFyTHK9kxv4vgwFwo1lF9Mnd4cfP0zpP
dT0g4wZ2dBYr5bxPVQ4TUCBR4lP+dsKYO/gKcsafHW0VR69cZHkIwMeO32wZ9j5t
+18jhKDpniRXMgQSBx9s4PFPmGcIBeIczluySAwWRV0NppOCezSAbJxmm35gmwXg
WeQcuGglwboKeP4OFbEDn45tICV1I1nfR+vGmAKvfQ5Vtc9OevdpE+AWKDeRlTGZ
OTHqRDyaW2wF2HE9IRSsumOkEd2X26Ab6PDUbkRfUOeSQnkIXOBUvjdT85YBFa8Y
XWG2ZSZa9/mbzAnLGyG+rm713iQHe+VyqiStj6ecm8UC5NCveB4gCdSTkm4pjSf4
2tlv7eOZzCOfVKslR/rCRmi3rVccda+A8pU3ZF6Phn3sn4C+lH7eF6Lbg5Jk0vH5
wZ6x7DmJPq4d6hQnZ2SJNwNTHlXzyTVWBzxXL1yKpfdRYLHleDy+vB/1hT8ejd6n
D4CIPEJnLVZYC0HH5WR3kMpH6eshRNk3z+p+z8mRHi6SkPrl6ZIO/m9Nr0AmNj1G
ZEJYv8Q8gSlDLM4inFEwTe3fueRSb4GRzkMsFLkUvULq0S8C5T/8LpnW4I1fIsm/
PFwnYFwGFbMR2LcP2zWgWgMQ5+m4pH9tp3mPVUzgPuj9g+aXoizr44M05eKX1XKP
G2OYDPU8zC9vCOmzv3G/1iCaqkkZtmoNL/3LjNm1xyo4Zj+34nqZmtlPe+Fym4Cx
yk/nhrKPFyiGSUZiPdUociMfClfS1c2bXeSj237DLUXrwYXV0g+lgILvLxspaIBO
2+EEIK9DZK0tDGTQfBF8zEKbjb3samwLNNnYFRWPWxSpixszOd/E8AsibVgiQSln
Pa+w+zf8m6Bl9VJhiCUMOmCwH30+AOFvaJx+mRyDSFaFsh7uwY66B8jP77D4lYcP
YCnwrNGzYTOgjo/2wfid+By+H32N5/+gNlB84IkUk9x2M3+Dx2EwHZgeYrDpv2W+
a+GtseEy2UrCRHBpvpWb2SsCxTVMNIO/bQmApWdu7JeMUcd0c5+dAx/B0ZbgBRiz
DqnePqP1GOf5HYY9UBIIIg4gOTIW4KBbMFZQWop2WVv63Z1hmP8rmN2+xidRCt1h
gNNsJsCC+C4VjhIqxA0qjqn4DG2p10ji+4gOr3QDy9HBq+90Koq6z9bCjy28s/xY
2cEHCsdyIzkC8CmZJQMgMc0Ql9Gy8YzIgcrKG8kz0JxeTCi6yj40td2MxWh4sw71
EzNV02ih6r4Rz9E/o5GPrBTJFlVFK+djkard+iK7PvsqosL0BhPWZGhgNTXKV1xs
+fufoyP77or/jmm6Q9uEtZz3WxDzSyvFg0Yw5XnTqI93AoZNA9WVVY75+8mDf8pZ
nfrlUjaoKDwU/Dy4VVeEuC8cg3QFue3qH5BKcMlttahHReG9jLwAE4btcpOV8yr2
EXZc35CxyGkzFrPlDYxMgYL/IqLltFiKbV0A7bPViTKeZ1jWqrrzvdQERxV3z/Yf
ijKL+uvUPreJ3vHNy0BYta6LDwQGvNeXzxyRstF17fqoW0JfBS/CN8zdjwdurrg9
22e0LuX+ZrZ2ClHCNeoEl9Nj7BRJFyf5tUMcCxDwn8LU0SzIjCr2Z1ylyZEqupUS
Yc9hCym+Y46rYpTTYsCYeiQ3keaE/dR+e9R71uKtqbgwYkAP8GN+IksN1y4sYjlC
RBoKpVpiBtXfGoj3SYuOLcjyaAe7nOZCdzfGEL8rM9EVP/z97FXk8DOP7PaQEKdN
NYPVDIlMgvpZGPZ1Zeg3H7qTvz6fXIJyZEtWUw4vaJi/u0YcFCuK+rOQXriy5MNT
9QHi+cGw28CKMxYTtn4DRTioX9EIvqrRSWrzAsPJAJ7y48bE7TcFUf1ntLqFMSfP
F/vQDpPFZHHzwOS5hdasx0mDHFLvu97CWNsHjB+GBxTm+yMGvLF1sco+3vV9pz9F
3WJJ21ygz/MjqSo95l8bS2G22rKQiuBEH6v3jwk4kEmhvAsqt/DvIND+EkOuR/0g
wP055X/kuNxV81NoPuTRTnWvsDa/Msn3fHvZpvq5L5mo+jjHTSUrUcmWUW1lEj+k
TsImucWlKb4QNv/Y24czsPiI9YShk+7dgbqewnum+8aGLRph+We0KZpxpG7tjvIY
aVOiQLko+a7O/j9qSuR9h6zSLVqEZzBfpi1d+6hNnVldT1iOfA2qU/zTfMr+715e
eqKfE+UnaTS+Ag9alKUsKD7v+VIOXBh5e/JrgO/+YFX4v792MdqNdDVsmThX4mRY
Jgl7yP9yhtFPjdcNoDrCvk/Cl6zk+2ek8ZvUlfuLNPY/d4HqbmaIH6185rgNzVb0
R5DkZu/6bzrGe9R+Bem21WcHaAfl5vbugJcOx1vGaCrJEzqo9VEzRMBil0EMjpho
L4y5vqo9bMrtIemv5b2XHO3OZW9tC7Twjh9bRvs6+n0uAgz3JZGqFOC+a3n5rA1v
48IUYmaPzfxJPiyyuBlo2sl0SWEVbBbaTX4SgAStHam4+qS5hHvN+HEA87sGsghS
kkP9r5gOrcynZtBSt9yp4yggWr+hpYS+kQ+xt077/vGiTTv719qKhMUeqDiKNE2H
a4EGa2sVAJSWRvxN7YFgq5vVeLXLiR1MDAOUTITbCeNmYncFEKcusfzl0AZN2UJD
9V38hQpohmO03nnoj27JGevm1q2k1Rq8fnbfRNIuQ2I2fZ4jx6pKqFxZDEToLk+G
bt2PD2cToifNiI1+XYiZx4pAHuUx7wVNxVDzz7m6mfeE2Mj2Gb0h46o9cuZIbTv6
EBWCEQUeuWYt67Ap062KJB/lWY6jKBm15AejfhUfN9SRMIe7UocNAz/aZaUu2WRf
I8Gk/cRJuFHMJnHydla46w+pZeDT0Rk3lFijORBWG4qDuF47EBpGAMm1wKadbsLk
Zz2bMnR/vspUc2wQR5fvLZazDkuUkJcQYBpijiqZXWSwZj2QZq8GxyZpoZbBQX7p
ncal005Xo97dJQ+fuBVLgR49YXqvjVUO5B/G4loYcGLYrZ/V8l8uCsAP8oFdgLpx
72SQj64SXn/qijGF5wTxKSxMvJW1gpT/cvqGtqLHO95ZiOVgcwPJGbYGdv8gB4Q+
a0TqRTVL7nNiz6aoe/f0Zfm161LATakwynxf1pDDQHt57HxMG/kguWjC6oumbiNd
gYDNuzyJ9e1scma67tFIAv32fI91CyFUhAj6RoHC1xZ7vcWlUFHm3tzbA9dW8bRd
sY3IB9Bk5nTTaCDh8mLyOuqxvVRAkmXqjIbB9SDAbttK68tFVVPfb2gomzsp5mSU
GUMnU4yPPaeSVLCUd8E8GQTyWnXZrglWIVBV0soyjMgNk8GkHYkzKErMae2XAcAm
8qvBn/18KJNCpJ/Ibja6tNUDqY5ZNcvROict5TQ2KroidsGGr66dm8ghB2halLz6
83587KLrYd8B49MMgtpUS1/AN3KssXxMA3g81rH9XAZ9nSByl57ijJwTXikgyVTI
gb4JhFt/U0ZmfMqG622l/otwF4TROS7XSsogGxtMbxir8GcAxnRAeuuj6MfO8+kY
d+PMxpvVmSlaCz1r1CtD+aZu8SsRJaEfHef8mOo5kbYNFWMgxo06BaNS8xd3FKtH
ajir/GOs9eTm1uemZD+rcvzKAZn7IFQGc5VoZ5i2QiSVJsiCcPDO/5VZnGSsfVq3
DnWtExZVNSkvNKkt0yDv3WbRMIfN3ncLoZTazpf8q2okbY39BUosvDPAW8DZSER9
Zmuqntgpi/BxGUj0CeIBpY7ycXy9tlAuTdOr2gtSFuUV3W49eF8D0TjfuHemCpi1
Uq+NbyaYLCedTcp66BQU5dvEthqETIIGULyZz8stBU8HSi8cNnYsI22VU6Xyd1L6
tgpk+yoWO9Jq8curNlq3LZd4UbdjYdGWpYG9Ng8c0FDWP6xaHNhRrypqfab1QcG1
tkZqQj21zz/zt50SqxNRB/0fNgJTNjqObC/Ughgw86zvELmHUhnCQdjzDInp26gc
lgt1SDOR4jzuMhdTvvRK6dbfWbBPINZKEkbpMY4u5dIYbyByU+yx5KDCnBisFeUu
lCLMiwf3no/Q6Gm8n7XLdUsgGXMw3iLqsA/J40yFUeaYoVWgnp0IETHNoVb0vHjF
EYMQBrEhWU/whx6UQvtR383HwAO3TfnmGOLqDItoVCSi7xbqdEALXrytmxRRYYcz
+pldQxEbimul55yPHpmCQJCND2EvjNvQ2B5LAOLTb8u/zGps5br+FKRRrzeIufPq
6JJeXoTJdeH/+uffAhKKS87NSczCN2fGY58sdS09ARklfiBmfrOwSMWmhBWnYFay
vYLWI82QPhuCKVJ13fONwO+p5rVB9ugltfnPopJ1HA7JI1UWB3+siO7zudowvLNu
lD0WVVUCvLAp+acr9A9105/UaOSqVg6vbr64gUn6IY++GxyePIA68GgWnfcF1Ddt
XTNQbZCapCKrxTf6rgvpghcoiNCnKP/NyvCjj9Bd8535inQJ3571aRCzpUsNBDo2
U6iQCjPKTP3i5xLc1mRR4ar1MjeZaGMIlFJxQy9x1RFzapoySxKW1vFxwdyOLEKm
cLCKjLoc0Le31RQUkEyIrwPNe4goO3/lyCwtPF1ny4vWu86oQmf4/9jGl97FGwfS
61hI2gZ7itzjJmMBjp6rKFBs/6cqTRCZdgmAPNbALW8QE46ywV/dqQyWBXimXhra
us8dpIHNqAIaihot4RCSZcT8AllAtwIwwpuuFyHGg3q1CyHbYLdeUKZ/8+7D8kol
03w1hZ3C9hQ4AKTGlBN4pfkONabJnUxgbKfcyn5jaXCDZI8BOi7wWJElVy79Eg4Q
EdjzUzSyveO+SuWz9cHHLYkT3RM9kF27KkOv8aAcOBBmH3pTZkkhLgxySD6lX9St
Ys1+KA+SiZTxuqvRYpPkMFEXyO/Fe14omOe/99lXr9gUNG0QM6uBTIgIuDDnlQDu
Phf0KgacEgKFkIRazpfLl7plFNoB5lRU6OfgonOYZnj5Rda7vFPGZYwuBLBTylzz
zxKwCfLytwl1ZDB5MLq4R2CqYY7IRHK+IU5+nVyzqMgShpf3wrCuYlG2lCxDH0CD
jNCfKEffFdp4VfBy/brkxGFti5cGloEsQWsx3a3jKth8cTLZcCgPuNuZkcwsO0UJ
p7QVEn8Dzg4b9QmdAYCgWEcoX7eZZYFYmNKkJzNKRj/BXEEQBhBbAPuq/4ztV8Lv
rBEBmEYTGvTbtFO48RYW6KneXmqMONieQjzwFIAsJ/Lw/Bgj8uK8qk4ep72ROUke
V8BZlOk7pMdUZ1It3Sii748HvAQ3H9qVDf8WX3ncNe2D0m7RBD1lDt7xMQ/VrnN9
csRsCHNXCc0iBc84b8cafM279U4o6Mfso2vvtwqZY1FSkigbMMQCu59GupN4PRuu
zlvldEEnzhFMw4Qw20k2CwVKU9dwQLnPnDPcnGswncVoy8+Ktr9ncQDqG+gnIJbw
AZCM2I+dyi3DK9tQMdD6W6IdM8CbFfgbIJYixQz9O/JoZBA7/GnKjz+luHIrO/8y
r1CR3xbbyXX7vTKLwzIur7N0zJate0d6rO2KOacRq4z2KkoLbpYA1ElDdlJayJ9z
thUDi1fI5sMsLybE8NZBuPaB6ew5JH4KgOpFwVeVverwLswf/JR3636LKMGAjmt1
8vMvQ08eOo36xgQ3ZjqzpQPp39e9G0alFLIG2C0tzxP+7wCFVovFb1Cx35CQKtep
cx/gxmppe7yDmvXqSc6oVyg7Gjp9bKxkwZIXgZ0z7soJ1tUH3VWIOCArnNQsZj9o
0oDFkm8A5P+lBSThtaYnkdUey2x1nCbQY65ljjtwHr8cBckPALVNGk+VfPR1Hnmd
BrAa0b903VGMG7Q2CYIuTZgRVts2tkwmLVHdL4Y2yikIzgZlRwTxBiKy7kQk2oRP
o8mJ4RT/41X1wObjDUsSOL++ciMISWSSLEerNPfe2hnkqammJ5BxqTwJIDVOpa3W
xFa8TwI5ovWN9vdJmBdD+FLVj+IxXROVxg23YISNwaLva8OEaRv4YpxXhZYaqTQJ
vhgFhktAfnqqSl508XFomX9Y9TEBSBTJltGcMeQQW7vGe5CgukUmImvtxXiKiMN4
NmXhEYQlIP7lOD9+wPXojIxbjz+g0TVIi0rD6r+VkSrWmVsJRmbO4ZODF4jYU5au
F7s9Ot4MzJTYqIv/IG6HF7nVNEEB1oFjv7V/umYd4Usne6xlnGCsB/2TnWs8NxP7
q4DGTM+ptQBBj1MYb0RUVcubqD0hSYjwUBOpu0ERl2EHOqXMdwcmb9dAjY3EXofE
Wc6aHPB7ONoxSEzc4DFDEScYbid/BxpxrQNnCvCyrdipxyQMpIhAgyW2Y6vN5E1G
yauH7R+Dt4zCu8iZnp+LO3YaF6zAW64LSLBuha6UtV9IxVJ81CelISg3M73tz7jr
5XUMqTz+Dc86GdrzPuxMgXLtOrH51JFyhaG4A69FrTBErJ589iLee2ZljMq0/lGw
ln4aiqp/wI81p/efFvOTN8uSf62ZwKsTpfmoUQWor6Ru5w8+WgCMHVFxLGskPRTa
P9YfmvdKTcwNdJwhyk38Q/e79h+qcTEr94M9sX6wrPQOoQiFwvDkoaLwfBMaSUm+
0IWoQJ+RCF2BxuchXq9buFrd/1aijCIeXm8NewqHlvG0p36gRYkIPLahVBGUcqLo
0YAd6UZpavWH/hm1tVxNexP3/az+isHl5GJ+8VfG8EzGSS7ypgaWBpPeemTNsIGc
ALBzGHcCdrUWOqTI+oj5wWC0bWgH9RrnWlLM2clohQDFosh/riHoLm/YRpyzxjno
KzLKkmMf+N3NsfgvDKRs7oLP7en+X85l1/niM2FQWyFSaL8VDw3Kk2u1FPvKeFti
F9xZn3UYuIRBhmnhfOhUJIUkFm9mT/XyeAvw4O1lQMmlUs5gmKlO+oDSImUpkdOS
anBRSDZq2+7ZWYuDD0RbyiNxbop59PA3E+/qzSdEFIzaJQQrw4ms3e9X9EYm86HS
hQOYCFwpFnalFTDuPOhlxWJBsWx2PDFYa5eKwCsibpN/wtp89GXpU5nfHPHr16gA
aSawkWcKb7v99glAEcgunh70zWag63i60dfjFBMFCfBnYOaLPpmtAvX1MEjWsm04
H08Fr+j0qKvRmv02JIL7sxDCv9mIsDL8pD2m90+djr5ldOb7GjSOaKP1wDOqL6HP
ZjcUVUCm1bgHQ6y3LOR/1UdFDYgUtIzrtAyzmsX4tQkgFuNWdIau1krf7cGPhjBT
aGGIO5iFpfNGWgYWENjZAvojEtt4xolDWyqbpVh1zUh6VJJXdWr4xGWf+SBAVKgD
sI2dWtIf78xuNgFtrvpUXhSoCgubNeIlo1tEui+l5XAKT+l4IZmVbp7CRxdoyAN8
FAiUM9PfoIvoDW8KUNxiKDVxmlOQNFcwbKtZKQL+JF0Em8Mlq4CDp3M9pLQVdTjv
8nD2/NnAwFqV3az6asJP8Iv79ykfM5HvjyrhY2G6rGP0UVplyQfThojrvDJahLed
7mfVY6XTfu6/PfurpmG4jYpK0t6at0dYysG38iUz7VaK2AD/pWPWbqq7LRt3RxO0
wFhPKvM8YYNEuf/upD49izq317IrZPskbimRM07TzqTPIDvfop4+CIBKw/D1IV3q
/Tg2U+vh1+8wRxQGdbA+WVsnyH3bQfnm01fLMOgdbIrGam1arsi2/XvMJlZMZGTQ
g5XAp6dVv8Pet/g9+QaIU2EVQoq67Whd36x2zMH0ogObkBIbOl63vMqCbCxNtdBh
wtFqg2pJUllKJD2UVHVUmaLjLwgVxL8nnwzpdMQb+D4aCORspdBC7BPI/cy4zGcf
pcG+vx5ciV2tHLTjAgD7Y3JtOzwnEo/InUML/MXLP5zBUwkXqo0qC/qN/PhlKymb
NzJwQO3QQvBA8YKpw0FF6/Lw43WEFv13trUz+O2auYtnh5Joyra9xl9eAznluDrb
vhwq5SIwA60wC3CvVQpLZg4zx39oy+xsfi1Ngj3Ghun515IawL5wqQyjyVEn9wH/
0Gbwfzbz9/P6cFZl5Qdh/6H9+iHsqRRCdZ/m4nT9y0Msrj6u9m/f/r0p+pAtGet3
AYT4rbrFbErafkFxKr2rSNA+TyTAhsufpJ6tN8KBJBOwIEQECRJCNSFIvd+nHP60
1Rahlhbdak5EKNg5Medfyj3i48ndX2AL18smKT8sbV5uY8e/1N6LcakZAL5NHYGW
CeO9Wv+wxQ/IBwdBdnuxBwJbQXoStb3nBujQkkfJ2m6esATu3r6rJC+kNCGOQcAD
eY6zs38gVfM0GqCYIGJSfb5mrMqj8pAr7Gggm58FEgv8Fq9w2UYdFNSAGHug2rE1
8Q4eUljfFfMo13p8wmzlma43FpzNWkfrWrHznZx2qVo3g68YzKrGIpE7IY7SFFJX
SrtZKebl9e9kHdNyUJ18iE+zEX3oy5Qw/cvtNm9sCVJ55nQ9LN5rk+Nn0/NmFOZi
ehFyhsn0vZpzYydABFDOdtfOBiCyNwhoyWscZi5lioFJkASkr8dn6L0DU/wndA7+
l5HRhOu2iJJifH1Dpa5xHaeZAtejl+xLDndDgPubJvqxFtEug25OXTQdHZra7Xje
mBxbeREkjEg2bqf6RZwTzOCZ1QjX/O1LIq9N3yJ+37l43Y8CnbU9FXZy1ESGfXyi
1DhUQlhLLQuJLucq74wSbNmg40iJwI6fug+hvplKn3VXKUtT/f/hFRXfIp7TndQN
2UwW5JQAvUFZ0cVOdo1k5o931/0Z4odmmu9r5Sd/JSETrHzjQpbHGHW188BA8IZe
+UmIx4+tOxBJ76uyDmnI5YWN15DyKv4KtNepb7eXCZifWzLBa9LuxzUD4r8izaIJ
w81T8mDI9EOPRWrDHM6rrirgG0puQx5KsXwOSPMKsE+kJn66Clipw4j/jPVVJnXE
m97hijZIS2LFblRd8kYDjPuDBYa9eXUzup6x25QjA2e7Wc5+WU3MSjxHZPDHQ99H
P+olClOOoOmRAwhbhFE0BLGWbGrxzXScguZTige9367lFJoSg4eFp4qEpTFbbgkX
2aF3FbFVCjPTsBDA5RTpnp7WdBacS/xALPw2YNJ2ZO3jus+l9e73c05rSLLXq6J7
KBENMiT2B+RD5RDuowOiv7BMB0jNUAXvPeQApYO0DL5vhbsjKLAJ5W+JTiBWk74g
lc7vgLxl81fgs2x8JGUSe0a8R0bGDghw1g+2by55v5armorF1koLeiFFAu+qDrex
vBZy9S2QqE95wwp89LzU8PQLbKERkd7VuOOK+KvVfGVbQ4gzlH6a/yZE6D9Z9xkv
Sao9MuP6Jxfhtw9BV8aL6NUn0M4Lv4g6+HPJMVnNVF9hS7wecrHhH8adekjisYg6
fEoPDpjvzyL+epinPBhPyYsG9O7UWcAILJnUoYUdFjxwGuIm4p+2qJTTBb8rD5oN
jTuoiVIVNBcasQBV/glcf0pF7IBSRj+y/xDiNKw0XDPTIcP1cV0UlMMZOIqzoTTq
cnQevSHs8nrkcMS2Cm94mBT/ikBTxYes9mtH43EL4Jx4YAJRUdSYLA05JRyGd+hP
cOpxUwkPu5+yjvU4UbrNTq94ElhsuJmIqLaS9jT2xcNiznFmUiTWG1FvfT9wVukX
ya/h0t5XM+wEp3UKYNRYxhTU9GirYOJAntl4teYaTXWz81KA8kPQkHTqwiFIYfY/
ZxltwT/gnPoih2gjAAWdQWa7Ji94n8QU3jFlYqyXLhVRL249lskjAVXiaray5ApF
ZFzWR3ZOmVti9ZS/wrGhy/9nYTGWdmTEhVe1c+A7gG9lGQydcTJfHvGiGBBAw4/A
5bQy2ZZq2mpdQduLOpsv20Sa+0UX2abiSLZ8HOp3BnAFNsZLt0SYebBTYp6dFXZE
Sp7uoJ0G1l9eKLo12ioRJ/fhUKzSLrZYUdZPTQ3iiESkeWKJjPzWBGxhOABFvkIH
w0BwYe4fXjV9nxDEEJuHH9PxgUEX6rLrI3MbyTOIt4v+rE8KyyuWvFgfXOSHwAYp
ZQFYIr10BLnw171LTxIrCxzfPP3Q3bisasTlwdSqUXCSe7Ah9RgT/r7g7PMWubJy
h7uDUDhk6e3QkYpgy2JP0wKoHK3haInpD0UDdFSht//zTL2nZlLD5zlwO4cj2Mv5
bI72QV0qeX0ZX0f1UOCCj/kozldAeOaQOHB0f7K7OMLcf1aFujghSrbodVOqaVUG
s4dKe6MjAhzERs0TbbvjUXIw5A1ioZSBpU15/dOsdIzZnlCBxorJHG0UADEg00/v
2as9xHJwXw9WUpg0Wv0JwQZF6yU2qpbXLeWIPCbDAVoFnki+TfanAdIF9obIZJWy
9seFrqSIX9UHMPljmB5urnrxzWeNonxznOTqd3UoQmXu3F+646RDWRHAf4Z5yw3H
vKzLHnrIUW0wfgFIgIbU/TFTb7YoOUbUmjK9lgZLCA4qzyjGOr2m2Fe/THKW6L6R
uajPaU9OXtNejGSy4eq79xnHv3UmoqgjSddEhVb+oUF2DZgcvE2xXDsM9Sdbpbpw
vUXZBuKZ4FwwbzxdosLvceedabaBE4CYbtZU7Ac2pBKaNSh4RzY/yAED/3grlgAb
NqgkN6kXpu/Qmon6AFU9RNJco2sh/En0O/tVG4pos/y32WOudgIMvcI1JiKjdJ9g
NZ7qkkuAf/IiOHh4W6/VoeEkPnmXzXdboXoQ4OuSD8/RBwx7qhCfCzkBfgo1I6Ck
48UPijgawbRdaA07j2ALr3iihF2SUZU1SuZsnnFojREKNTmxUrGJJLbxJUhO2ipW
JU5iPHdue2wMSGXgdAAhJdCr4GJjR15VpgHgZ5lHZgd+LpAD160V9MBCgiIRyJJk
AlLZtmSjnWzSsBTcqRkpxyKvShiwz6MoQ2wVx3uETkQDGJMYglk4KmTEQ5Y0CYtZ
6kmqZmDKeEPL027QGOzl2vz0gHC5ILblecrw8CHBVZbz9lBuAzo/iCw1U9vn8g3B
MDr3zNtsbhz/X0bSzZiUyf/h8Xfc9l5d9bu4tS7ak/NbmyLnLfONG4lewkHrE8cT
H/tI3cZ43jOjFtwEImwd4EjidQ7sy3n74F3XAk7jv/UflvEnpmGRhuagv45Zfig8
l2kyr4L3nIqmSoja2UOPTQ5MQQgZg9Gz2ImZIq8/I3pIbxj4Z/T+yYtnzFEuS/Mv
HInBcE2ZF3Qh2ftw2ax+3DWr4RVb5jZeZxoef2h657CRURipPkiy9QfBLTTUus2P
aK87KPUn2oU+XoQ1ShzmPaSzRhaiVSFy5ZqVov43hsdumnX+VXV6q4RzLKqVs7M0
9ozcJ+wDQfQsbLR6f0lTRC2bvBGFAR2xw0g09QUy4OwOpINgUA8e8PPAuJp5a5m0
oJIyp5SqeiwxRcRjwai2rhU+5/UVUdVwWAfxZNcFvbghqomt1r7nPx5VhzVUvUZY
jSYnnSdpKMXe6GA+UgD4fuhanDQdo3TdNWlqdw7ny8tNzy/aSk27GRfIhKzY+E6T
9Cfz/GqLUZGL81WjrFksSHqhqcraHJ5leV4C8nBMlgtGPXdQJR93YzEcoPxUJCC9
zvbeoMhHO2LAsQs8GsVWumLkc2PdGNgBvwn3nhAUI+LnjoSXLEHLvxbdvlLSv1cD
80UIgBhS99RloPllnSmONr0hI1bQpxE3kwAkKu40zZhmxmULnIRxYxSxmdaSiuur
ve8RA29YFjG5vc4SX8fzQHCwqbSG3AGUDxL3wzR45VClZMJrPzlceLJKQlAfJb7a
YjgXVMk+WwkeNIF06Be/lKEyKc1vC3hXKAwBFUvlwA9UQ4rwZzKjf5MfJTE2KrUR
It0uysRIG3NWaPRAVoXCavU811reQJDpPMLYFgrxVkHJr804ek690KuQqBi4h+N6
ayjXkspIuxtCfTLeqRxVhGupCMUUHj33nQXApuPgAiyCorCgbvZ55pImrXxqShiV
4jP1+wbCQZr9yqH7kGyom5uFfK3YRp1cuExZnRuqP2y+wOf/bsne1irLdTTZbpQL
tzbhCMN9QVNEZ+8DcZORjGgNbKEmkMf/MKwif3itmLaDEg/yncQx1b54nJzQ4pTJ
BncuBAwCX4bHOqBEH3yH2aBV1R83MRwZQINUqalCGXABfcWxcZ1BsuZ63qgO/1Xj
8h0VJiJsTFWtIFNznmNGSFyE95G6wdXerkcDxtOkicSwFFhL1y55zLzFzzhZKWl5
KQDItulvjx2YYMSViEHULp97HOw0fHNFoWBeqJwYwifVoO/9qEO3SrZRudEvqpof
PDY9yGAlT79zVpMUQctaYlBLh2txLVz2s+1XdP0zJvGreoUDDp2TQAxwbKnx3Bz3
0+bmTwzQ8YqCe1osnvZl5cUHpMIrkdPbQVGFq3Agi5R5bE7AzmqoiV7YaXxBZ5PF
sXIdrVzaLndHXiKzkSqcQD1y5r1fr1VGsh4nokGAwSAC3cKt2QnyCd05sUEbahU/
Yz1208HBXeLUWNRCjOktr6cC4ewCIxuOUeH8DavKMm0ZQT3CMFhFi6al6GPW/Xrg
oLq4v0TsGdxBt+j7svGBlaG3fM8teHOfU8E45XDu144D0gK76OoxwEycAqEDbvWV
plLAPq+kUPpNFClJncv/w+MkvP3y0RtMyspKBk52tSpYkhhVux92MQP29zQ/wqmz
N4wMdhwNtKeAuQWk3yWVGF7J1wtM7z92KuydKZDMWPetfHsmvpm/Tn7guHLmdyYj
GoOWsdy0r0nLv7CVzriE0fVKfQMMqiHcVG2g/ZJzpU5ZomlX4i5N/XBknFR6ryLg
8IgcX14wZ0B+IFrnqTU0olkAKOlUSOJU83L8mJSdAdeqC0BO3vnE7h1rktnz44bk
CQbmo4lBaxLLv+7GaRcUY6mECVtXPZMzW31mjumF9RwUOhyM66yjWeQysF76EBdm
F5vVLDIg11+NZEzk4QqtWuOyotmL5tTROptH1O0VeP38NIWujpZ13BQHlj1378yY
ctgxtYTwOhfV6ZIdL8Z+4xOz3Pf2eaxa4dFlS/5KwqjlQs/3Eb1S6f5FR8KNkV5I
Y3UVOvickVmkFW6QmO4iBUJf+Lz4fG5c6h5Kkj/NzFiBcuEW4fFV7qNAD4KMX+LV
+lSHWv7LmXKcb57Jb9rDuO210sTtYBcn1GTcr5lYHC8sfzYTNftcVDWE9cyJ7/C1
iIkw+0qIVfMj646LNwVJraeiaNGDddWl2sr10ehiKVjwpy/yQzdI3c3+YNK2aA24
7KYPefxdehDbzkPhdwr5PW3BIl/q4gPb5raqtuye9PbdpR+GUn4QvmhCzdHA4EYu
LMtDkwyJyjlbqiEDjuDYAZHa5akLxr7n0+wmvEu5tn47ZmRDqTQS18dNwTFgOv7e
dV9kkJDOhxx5qYOIz6tc8R9q6mfx8g990/xyTmAWXWtF1m9ijmPjkfxrG9T7m5Gj
NWENe9mWpjhqBeo2j6K7cIvDQy8XiqtVS+1aE4/TYfjVrbnCFQI5eM8PxuE8QJnW
t3XfVQzwJYvJpBkXePmNp2niFs3DlyAW1jCU5X2I2UvjyuzWQVAtO+VJ/v2Oj9i5
v8xrCmfKXv2+9jcU7P77PMJVyIrtVitzA03ZXwMlNukk2KZ1u3pSEqXbO+F5xi9U
I2+dOmDrKBVN0Ps8hyG+GmoAN2i9MIj/7c8JRzMTEXMmeZ9dN55kxSM6lk+JfRrp
Bz5IlSPmPxHkcFf1VnlkAlrPZfS/lIWiW3hLthTpdl7FIz/XLwOb30eRpoEnAi69
eP9wdDJUWDn18s2hfPQiMNbzAIhOxnlwuh6EwXsMpYr1VNVAsj2MWiU4BkZoPhcH
07oVZx9T/1aUvwz5PiWaj+dvmu6GIhIgiAT3I+62qNlUbu5v9wHBdxlmSdfu6Owb
yavYC/S4X5h+pVpdQwUhXgGkREKWWwXr1s5N+Z7nkkkGlH+fwE/0JSOLHg2dqXfQ
WudvPwMTPY2BdDdbASQs6L1LWGxcxWeCgeDNAH0Xm/cucd4Ue7VIGP2y45G91Fsc
M2vVNaIRsMpfJ4rrBBRb7AIx1nXbjWZOEl+SYnlhcL3njrdESBNEXT/lsKxzqfGr
16AKGv1H1UdCqBZWuejJKp/AUpBtZGnCPwpzeWbm7t1Gatkpu9VR7WEl2njNnmok
EUfF4mDTBsdSblBz+2zNx9O+zy4/GNGCvk7dxkaPGysvmqKfXSYFHr/mkxCbPQZ0
vjAkUepqgjGdc9Ttdvbs0De79DXHrrp7cXFXT19YSU2fkUYpXc1apGFvefzRVO2q
gBzkrWOpYQAFG3o5yPM6Tbo8fNmv15EfSVgPYum2BaV8xl2/tVBraFrBX4dHgvnt
KXssl5xj/OYkq9IrxmHK1wITWQpG7c71LEbIlw1pigD/Q/daKLjFr9pfw7TrzsMz
p7NsrfauMlZ0HvxjsdxBn1XzztewQa5qxp89Y7Z8+gT3ad6y+FPc3JPme6BAXc9g
nxEK5r6pe9UotFXKXx9eCIw1IbEc40j5oK9icRAxN1aYXFPpkyI4JTOz8zYYlpST
yll7MBUKYkwHH+j0rdERSnuLXjwPlZgaqFwYN/LwAk8wDMkQX9Z2vLoUW1Q7wm/R
D0AR8j/vIt95JTLxBkDiBbanWnHaXqNsXhUBBUqdeP3VKZlharv47H+yNfWEFzkz
RYB4kqFkStXfMm3IBvv+7WCKflHmMTO7jFA9Z6CcJt3DEIBDuf/Njt26gft5qC0m
75d2g2buNAWuu8VBbaMZyHE30IYVQJt9xhtP5G0G2tjyoLzDh5cZu738nxdfRCg0
UPuF+JrIw2PWXNXkbt+LRVLS4Ll7B3koVStnYUtB78aj3vyhD76s6dhMq+UfHkwM
JNzaPBOzpdCoawFvjxDbBNov73+ABJBGRE2W9DVmk36KaTscqU9diCunj+t1uq32
wsShzcMoOWuDs9HEL3LWjmRY/tsbBhmFuHwML3ajgkc7Gj/yBFiVpGu0SLKwvXPf
OTWl0qNfGOG3FU1QvlkL/K0kf1XQWDXBbcUIOLorUH8HBJmMRt5bT5Diz5olNCNe
Dh/PhMUBQfH1CboT7z3IJ2QMM8U0s29atvzPDfLExlsL2BL4UjKy8A4ennKwOgWa
asmPXt+Tn4Su/Z7V3oJdZtDw1nrFpQ1dPRUb9Ri6bp4d/ig/CGFd6XCk1nEM/ipN
9zuBVAJ5VQB297BwTv/OPih10/y+pCZAEYsAOJyfgoB5ck7fcP2t6Q84wzVDiXA3
N7ArEh3gQSbPYw0bYxHp8SEfhqPe+3zY+p+aT4/Mhvi3HabvWeGJeaCB9VeKb8Y/
3ILMbahVd9/gVk3JMb3xfsHTmfrbaF55rp4ArkFx4WaNWrAhgbKuSQYN0IR/Ps7b
301WzNmtmK7uywzJz4IotV0N1ifU/mAJ8ORffG3E0/DCEczBDlwXI1M1kIAn3CWj
oS8Xl/mMP8DDJ7a8kh5cdht6kqi+Vykr4qCOWPzIybTIrDuIn6ycIE/rsLu5/zF+
6t38RI17vk1RtCcVeeC9HqpllNanvao3NfltvbPV2peTf2XoZGYbzkOjySnuItud
VeaWYFbI33/tcduucCLfKtoEnfbsgNnWHPji/w2ehEFhZw3wl5/I56dgO1vwuX+R
tLG4pL6I8O0KHmL46UyHtZZkdCF/zs0m6UayYGJ2v+O4RQ4IViuzN95vKLRYaM1n
jwv0+7hF2OilUW3iXEoczhsQay7hF2kDfD8QG2DtOOlWBQgt0BSzF3fcDQ/DvEox
oCl+KTQ1yQGUX3g7AcQlR2a1Snim9fmU36J7W+lZWdjTDNZHr0Mb2YAcryAPjGaQ
B/IeV8jekZddEXjKwrGrwkM2E6WeSdypdd0j1VQc3ofOoshQM+Y3RIKWl/vb6DCB
VkerIwdeAvzhj4tHXZN0qAgoI+uMDrD+qyXWuYe5PUNqI5GVhM20cfkl6uvMf9vH
3NxfMNUTLgrXwJuXAQBh6sW4TypS721oRCbIW/Ij7xHhAIVG9usvwfG9gC8hGiZZ
Th+r2Z9SjRLlWwW5RKi6yl3/peFtKQs+krYrXvIlDJhwA9RTMQI6JfxpuumoK4S6
e0erXzfSvGnowQCCDOSzrpMnOnBh0NgVteU6yzRV0XvWxFROXbw00heuiFXmerDs
f2ZmlKA7i/mKDG1+KZan9bDm6YkmZCTZxpIbNGTbxpZQKI+ZhmbFvWx1X86S6FnV
q08KwspYsFPtQlX9eTdHHYnH24VlbOqi0DrnB+hhndTHerZbxsRPA1AheYTuFHQ8
Rzkm64X3AhDjtmZK/tk2JyywNJQBVSWCjcDT5fpW+0eFtrpvWX7Au2qE2kh4L+8i
B07Co3H+PpBGyG2eBSa27i7uV/Z7Q8gx8XOldA6TCcYBStkLfvuFjCcZHW5oIeD8
GCiqzn7yHjN3siiWskD9gZlHBUhc1ao/FVY/ezSUtqry8R3J+VsO8H94WGBPnzy5
AcCczyCbG0kvmzcPWxj6hIc0mnVWwGJ9qLSvwZ/cYdy+XV/uLbu6Y+X7OgSdUnpJ
xcKKe0J7/huh8OsyYMEpBl7F4IPwtmFpd8WS7HIUNfjqtIMVGfkdOBQ0M/3EW/eB
pNrcqobABuRV+k48AVoscDia3L67R+puymbtW3oEx9mYWk2qJDftmlM4YeIcgYTn
ZStGLaD9fIgO9tYrF1nS6VwRh+qAe80Z+o8ek5Kh6MJugewB+glGWaognrmvQG74
6b0Xdxm6B8VLP0/FMVTiT0VBDzo9lP2oAsHZWBYCpPPsJIJKzqJy07cch0B0UjVZ
rQHLdVdHsuHplT95lnG6sZG4JzTCGu6Mt9yjESzo0n7fsjik5ABSDNWWU4AkNS6V
cYFHZ8642AZbbnPRNHoH9RTwTSirn9iAwoL6M+v+N04n7Q+YlYiFXGk2uCZXOTaf
nj5m1z+bQ/jWVOFA3XZCv6j+ed035a5pGZ4en0aVvycEMzIqZC9V85TIxvKZKLCd
UQSI1FEU9Gn0ENes5yQdk49JmIXF4yMibgASJPST4+JHWayANWVU5kjCnlfh/DES
jWjJKXYs8h8AfTgBZADOEbnryyzGuEoEiiY4m6jopN3Y7rXUcCv0msyMdnRDGqq0
m0nvXEYM098GYLKj+io2QbLeQ85ul8oMSfN6iaFV/M1z3qz2OjstGtAF/N7s22TB
WGgpKUqgF0o7N7J6EYvLxyFC0rz1DdvG+ksLJMtPVynoERfpBEIGKuaocfIHrl8x
YHOZGb76ahW4RNiV2nGP9LwErVEDTdS8KmIf5H+VMSkkZ4/OJjo29S/PXAgcubFs
Cc3nNSBYNL+4CMyMBb6xKPMDsmr7DxboGvIgswqwMQUMpk3uG7pXp5caydAvzuUH
K7P/EzNNgMQOqeweQf3ggHRE/naBuSZWzcj5WIXmmoywvrfvUR5zktGx9NiD3KfM
UmQX6T8H57pXGLj/CF6O3RureHKAU6rtpuHRIo9XPt41rPZ9ZSOEjFI+18MwZADq
VdQwOJN2mqfJUBHRiFSnLhZd0rtKUGhxSSK4JqHP5iTgFNpUDHkaOmWq+WJ1/5P3
7k9mmuHjfZW3ake8smN1JWXPfx4p6gqj9SFHNKpomntB0D+cufgamlUUo2rDtphW
gMuEGot/LnR9wVM8hvJNeeqtIHPYyyaTi84/8FY6fLZCiGcgWuKvwtqHLcUR6jl4
DlEBC48TPiVp0+68pZXj7mNvmlKzsqKH633wNIN8GmPkPnmGw44gA9O6KDHiTKrk
sPCsYH+ZIv41GZ7eYMk23OcVptsBOkHKGJ3akuEN1MRDowbcBZRQTc3ZXsF/c+mN
aRPuu5gBi0aKjhh6bUWh8+Hr5VWtp33L3YCgJRB+GvtaWpKvMONHMhD7UG5H1QkD
15b/kDjlMwsjy7R/z3OAJOWcJrkHEg5Oip+nni1KikLfgr7XaOJ/qn60+wYx2bl8
GDetpz7/026BeIRDzCLwl633Z27ObcgsGGSZbA8h3BZ1RVIFMzYoiyt1s6UO9SQL
KAM/bDmLmrtAA43bP8t9lGENCFTXmYXxjGcRkrwTC4aRCkcrCDBEFpccQecOcI2l
3Yi0E6T54Tjw/ApnTgBaRf2GX+19OD7j+oPIi9vyaeN7GKc0Dy/xw9wpKLL/lFf7
F1oAV8M7rv5BbFk0OEfSVwX1Ufed/kJdUDVkwm/eXKekPtLp40CPY2IF6EeMg19+
Cfuc0ZfWOarhMOUwKE6avRSJcJ1Vcniv7buNYwwtETut2D34invULyl/c0Kwvjjg
0sHdkVzv/fQuOtlu+KkuUitl04oYn1AZ4IFWo30T6esIppOuXKLQA0BAU0DYd/ZV
asR1EwHgcvAAM8G/XU+Mu6SHVVT/KJ5X8DUzrrFn0xuoxL86phae7zugwy73o1kr
9UfbJqBU/agfvPLCMPG7PA0WpI3q0U+G4TykxWBLb5VJoDFlP7XiBWISVD9fa2sM
NKdg0WPeIzfrTN29jpOdB9P/RNZ/gkNUDjh6VBv7wvktFwrge59OCcZBhkqGQdWg
VT0Roi6VHmJ7NKftmFGN9DFgYMBipqltnP/YJ0b4Y3sM9RZ0vjFScLenvH8//3bJ
3R990M9f7NV508emDd52m0uQxHqW6YjzJFA2HDWL6XI5XHGh+22iqc5gZDvX48DH
mhClQllqbibIkwAy7pZiDiLoTPXAqda0C+syT+kS9+TxnmoqVpRIfx+fL2+VEijM
deXl428C1BFf8ppKwlvdAF4fYV34pXqJVcjdLwN1B7wcoNbv1z7ragjc53qgEPDq
qza7j4VIJZYTq3/fmZ6IA5ElkzrZvhDm3IgsabuLDG8Vb8tbp+MhuaSyAj5P/IVa
1VlaSesJhPPUwFjz6AnMkQsbTABOxmzjaD9Y/zZox8YTdN5YRvTqZt7CZgOaHTC3
dUb2Nq9KDMkySrnQNUQ4qzJIUpM0uJLOinyFB9q7RakiCgea/EwiEYvGWCwIaxCm
N8IQXtpBZUOw6axs/E3a5+oUANa81J9PXM91ggFO4clHxXXoMliw/uRsIZDPGoKy
QKkpV501pg8gD3rzp+R3AsfImLNVyCNg5oJkGL//yL2RqvnDFcZyZwDOhQZ8Xqzx
df3qo/tFLXfXvwXO6ceQGa2u8ZmUD7w0LazNKPl+PoeTIg8Jynp3ZuhUm+VBp6nD
xXO/85wuMWXPckn3SQcqnVhSjwY9x7Ll1GG7VNzJvOuKQjQbC19HYBnKXqDg8oIC
EhA3gvw1JvTrccde5oegevPjzWPdMTnyw6wO2AdiVdezbkdNy+Zj2LDoUtP0oIDf
0HkGrggO5Udr5tzShqvNKmQNCr0SnY7Hs4d6U+BnS/8PjwM1fG0stYf/UYnllutF
BtqtD0P3ny4+Jiyd787Jnci3+L50ehrRKZdaJlu51pGeT+OE62NcXSzAs0LSdI/C
JyKdYd8LOqmEFwV5MX7PkGhgdl20rXnmrVRFBEEuTrOdFydOGSI9HuLyGWyWM1Pu
bIGh29I8lAz4/sR1HHgFuYvHi1kUyK2fyv4eSnnNjIEQLNq51yuvmFUG+ge2nCqr
Ew+6hxDFGV3mBGsFfP27pYB0Q4GJqW41AKcdq5CaLpDaGhVezPltLygBCN7JEGpE
+6BSK7PJxdiDdElLOH9+fnGXXYFCrUC+6PQw/EoUZqH3SdEltRhP3y1gCb7jKpzS
+yc8NvK3VpX+eZjAwddhO4/BipO3/S4dBR5v95J/XlZz2mvwDHDT4sx3W7+UvEed
sNwTBhEZHTN4vltrmUPpJGA+smhAVSF5rvnISSLNI1p8hErGWcRHFwpPVQv0JFBs
/qKGadIxSsPMw73+UFIgWxoEtA3gz58wVTsNuY7bX96+gWK2eylnI+oc4mZJohU5
eLZG3Oo61PJ00PlsHNRl4e/q9mxDxJoG5h6Ag4Bv1C1U1U8yiUNNr7bBAP7189oO
aveVYjO4onr/g395wUofRmjwCs8NUeYhj7jnoWW89aaX0Qt+rMLrlQwKyhZeyJSW
nL6y7B1NrQjjib/3B59Q76FyZWRkW7IQ3TejNR7zaObBtiU99e8yNcwOShvfFfUu
RdGx+39lQfRrHZFa8sJa5GDjcVVJFL2S+VIRSs8s02fjoQQrzbTBxR6DxKQ4H2t8
RsU7BKpGiIB/xObYQ5cbNa7Cowbt/2qHtP7ZB64ceFRz3Gypd9jcB6+/A7OlQx86
rfqEhSKq1DVslsjG+NXhNLGKVbjTuYHIjncqgpcHJ8Ze6wqJnEDboiafbgSHNYgO
EnGgVwmASqhaiB8DFOst5JsZQQpFQX+MfvYuax6jXdkA8lhgADdoS7XEhYDdduu7
v4BB61I6244MuXkbhBwBZNCRq08BQCWbCIAoCYrsHkxsoZihnb8Qz8wFduELhOtp
7zvQj5rSn8wIZ5RAjjHTBwCYL+NQ2MdlSsA/tA1F9YhoZ9kNIS3oWGFLcvIXGEZb
i13VKLWdUO8CJiKWXqyb0gckm5PhOJ7Mg7eg7ltUsmDBB/ogfuZVXfM2PqGYd5lZ
T1QEtpuuNoQaWCuPMKwi2W2yE0nkET/7DDexUrMz8pNPqPV8YYvWDFr1SA0skutz
lC8rYI7ROyHGsChXEQycDZLci51V9fzcpz8A9juAEPH9MiQW6Mrw0OnbPZ5UEc7N
WQelVgwggYuZXvZ2xSf8f1sox7UTQniaz37meXEvPKwp42E5oGukFWSMgXXA3h6x
4JJ2sLIn3CecPBRfXDiUDcv/iIDXhh9RYs4tTGqxVVgqFG4f7PsBex/f91ZpYFUF
IvGV/HG32klifA4jvic456bTCEvteepgeaAP/dL8uBaSLRGz1ZGYHE9bcRr3giiJ
QlZOkGPL9UQfCnEmZICqZdU9uwKs2I3WD0nBjhhBSIGNi98cfQLh8sw+Dtx/BbnM
uZ6Dk8e31mYQHiKWEkOjj4j7Rv+wHmKWKjwAX3U+6bPRkCvBDXIwG74VBaUkh612
AF8UISY0V+MCBZlBx7kmLy/lk8kv/Pc3oUT0KTDzgVI1d3xjvT3qfzR7JY2iYDwB
4XELUBxoOiMYL/m29SI+nRB+WZpbrz8J5/PQJTddRWDrzcfM14bF/eeO6LoC5uu0
0GdT0QILLubd8YmFKT4oLMWjlapnD0+WvT0V8nCiH5zuK6N3W8SNnD+EfADZCxOc
eY+RTF/HMrpo7+8blmK4lzjENY3QbX3WA0UPoaNloYgBI6V6vVzhHLSlZQODdYnu
91dux9FPFFOjslWa8RVHNe2gqsLCz2mAeJtBbCytXyZT9s528ucg+sFH2BGIj58W
ZpuwF6b6C+trvBBeXcWMayGg2boMUQ1OhY4QIzAtyFY4aawWwaXUInxNq3byu4T6
3F/d8cUEI5MRi9Z8fG8Q0volt7cz6ZCrF9SPpYHhrEM8QM64QH7l0eOxc/6dhYeB
5WnHxlcdwOWvx0Hs5FzfBeVGvXWlchDfLqlYw1/keMMfnaftHsD1xLxCorUV9mGP
FO9W9oJQUxU0pheR27D4yVv1eLLBuPHF3jnlrxRvyXpUG95/+ijaPPvXFBrpzOEm
wRbFJx3GG1NNNepTr876eRPcJGQQktgZ6up7x260jN2XBA31yXIR/8o2qilIpcsu
kprMeLVoCfWDF3K1BmobZb/WL7vIHKRSyW87MZ0sBWy8R07apPW0dLUkayJiT3MN
YsMBGUJUytGECPFNSdQuH1kYK5PQITfn28FIsyq6/2QPWO0PZY1gBZlYXIqkuuEG
NQeUgFuo4SwSUW/eFmz9/t6npqRyEkqapB1j7iLV/iWjfNRWGwTVCM4jN6+hSRUx
l+V1YYOCpHb/d/r3QMk/QiDINtYnT460qoFhYmCHpwgct592s2yh2j0R0sATBDrN
QyqyaaOF7riH2yCLrXZgl04blCyJ953QSYHVnyWRStFhCZlrI0maRd4UPF390TYZ
9guonfkiqculzJSTvIVyRyD/69yLDCcKfsHG4wnVbn2QXwKvyO4jE1UIpk/remch
Y1DdLq6r93Qm4Ll25dAuqLCIa/89Twr8PVDw43F1Z8y+rZqwdOkv8P7YnJQAVAUi
nEEqU4RISkTuwRUYeIPqE1W6L9PTNuRliwWE79gNwcQmocZO4uxmL8pNibuBnEpS
0sQ30wNX1n2XQ7Xagxobar33YvqkcKOqNLnC4UXzbNdo8WIKguRIzX0y5x1hI5sX
jOEJZIggmXJRhtrjgaqT1pU2BvxA3JHoOl5NUfC1SqwE6py3lUhKWqCwvRbaLQts
Udb4KjwMwgqf9m9571b5DffVW7t0z0W/Lw1+x46fa2aIgwNsbprSarPJHRfbCHkt
vyCIDCbK745jW/vvNAYLm9wuV5st33RL/ro3nijx8ORZPJ/yPTwB3LmNkJJwexdd
ryvRKaBLF1J0ve/mt1Lk/H5Nnvu7wi9+S3EQ4YEtlUqc8F62ZNPuCYi6dabB1iok
AQcLMz8d2fnygjXTbWdA2J/eGcPNwSErZ237r1Iw8IIZn2M55NruELxBwKQQ3u/o
9KqmsFN2wzL9xR1tQbFrvQlwtwl0XekJfcm8gGn65I6IdYfRtxPzVB10CMJ4mSHO
Jc3wviWZUUtvJugkaiuVvZAxaVgnuh/QEIj3TGqaVee8lcYldPlrKpEfZ+rjp+b2
z9VW1zHAcgkhYTGoL01d42h7epsbbb2Njbkh0Z171wbTqyemn6cSI1CpXGOS+/4F
kE34w0/oSZn4IaPFUOI0iubF9GqEMxvyyq2dKiVLcalHfeC9qlY8WKv2eZJOm8Mu
56ohEYeG/SzY0pu2TTqXM229O/hbrWxh3cs2HKHf+ZvATFRy0mrlZcb1rguKYIk1
bbR6skmwbrsZ/0u1p5lsjlYzkIv+KFHGNNTqt1/6dt+ioajghboEtuKTzzNfvyY3
AsgNg0MLmluszOJDSjdukzWEIrpPnwUTZlvI4IwQMRrhvrMU6IqI207lBzr66wKB
7yF+YB4F4wmVraTYQWkP9qiF8FxzOYq1dELGZSIx8sAtOVNHFyR42jxyBrwxe41D
yZU/UroyDg1ZmouIqD31W+MrZeLBMjnsUH9e0g7oWN5CZl3+p9vJUtNN+Sve8UpE
hUhKheM7DSLa7BbP+eR/UTYMLMvZv6Htfs3MPCEnKblgqDnsCgD3Xb/C+HYfIYjN
L3WrFZpW4NZAUD20CZZZHrFdPH/piIT8oB2Qjx0KJiqXTBveieJ+a6b8heqBpje3
KRReYAvfvprT+zlL+ZFnq+LPVFBWSJ6N1QKpuymCjHpnS7tYmZm2x1dK+fSA1KHS
CWfyUFOT7qtycc5N4SPxAJhHQW7R4eiPNipR16IBrrXJxNFP0T0WHNqa2uAMAsm5
SqchAW+d5KRV++H6EcPPPmrD0PqitBCn+VHKAqb6jeRBbWYRebRvhZtkZPPpD8ec
H8lVFaEDVTqESS6xujOIwVjLn8vOqMMRQrhzWQeLr9k/h8AKEZqNaD11AORC/Awu
PHpSnWjbrYErqP3Ahp5irbh8ZHW1cb451rLRzZf5Cd13uKQk4T/pW7pTiDwkDyKC
UwvJOpVa7LwlTgE5d9I59PjxtNAFZEf5Qh8i/BZI0FOOc3ak2NPpWtMeDUWLWO7B
E71yRXA1pKzW+Y0zG+i3nWris+5i4ze+p/2dPHPN029KlJUWM2HScS9AdJ2MxZsi
w4fUtwarNYon0508V+DgPu/apSF8+WCka9cxKyN6LPpJsF+ecWNHaqSec/3PFjyp
MaDpLFW11p6zcNdLXQ5YDLDWWgR/AuwO/+H5taUHVZOYFuXP3vkKaoCxDBcMu0FS
E0vEFP5++F/Lii/Ek/nq5RtKeXhR9D27s3+DRGmCY4bhBqZq209XUn2Kz7e11qsm
ZtDVHMxaoCwwSBwqRhjvwc2a+v01AXDB26mZcRj6k/Y4RPWWbSyBk/PwSTWTgzyi
YbFqEC2kSS6sMOTfUvJ85QeivWPv8ZJ9nr3nxEAekPRhvMwYHysae0ySt/KARwsz
Y9HX7gjebwwYf/1uCv7qLjOv7FOX9i7D54+rwQ9m5QGKY+/Nvxal0ATjgvuv0Sma
6WDnM55uS36L6fnMnJZJI1vLYUFGoFXV8Ab325zr5O7uW2Ir9MmOOZYpZOhQLE+x
iZ95eEacUyFlQhR8cJtHJdbhYAWmk17+7YZLkAKSMcuSchObqtIF+NeCo6LQ/cxc
n403KYdPVnmb4XvvsVLHpd9Km1u/4kvW/+Ym31TE6dOSoe+sDsK0mfPKXJEwR7Hp
8L6wA7tVSdyZWAQqFKcHf+lg/S2FTv5O8xnvoxElG6rJbI9tIRJ9jHuWISSM7eAw
0AjgK50xNI+kU8q2ZNGw9VCuZTfUMX7DFxEkDEAf2ptXoeGz603I9HOUSPA4tAi+
n53pjMN1ggCq0KFALyPQQRXS/8T80O4bg9vYTmtptduZJ2gdHBXjFFSpbHa5u4zw
J8clvTBZB7tuMP6FLp6eg8tIbGM9yTPOC9eAT0t+69KxGNQLGfvwUYt5jtP8yvFg
Jc2Ox7/xH520tONe7wKSp3zrCK7B7hTha7TKpBSzFpIMCgIc26wHXAyaiIbrZOfi
QL8cmUpk+7l0jQRa1ZA0Gpgw62BhQ5zC/KFHu2OV2L4YfYcQIA6SVmNlNjYVogu4
jKcM1a28GRwiU4cYbBYiI4IcfjVpV1aNUY6dDAuQRwVS00LicyOjtpfqOeORn0SU
fXB17FFRZhAXJQ8SJl0kyszuAYbOGaT1tsXigSY+cu8BO8lofVR6Tw7dfKnbzZAA
dV8kYvD+3wP8dc2fH1FIIr4uRgeUQGunoF4lkKGr0G3RGL4BbryhO3p/DPlhtQ35
Wz2QKvxGEFzpFw71pVYSqASNkSO8Gbdp6YJ9buwwykKBmH5aVbv5dGV2Dx1+6+Hd
CJS76ZR+/5UvcmEN/vyFTaSNN/OM6ULbShGhhFOQ7LGfexle3T0FW1cfRmaIpgEM
kD1BOiMqkXD4yrcVvnLRvUhsV8Jin4jF13rDdw3e1Ft665l48O2x4kgomP22EUxD
cJ5ZfYYCVWXav9MjjPfyprLLhm0OD4X6H7PwLHwdVhyhqWZ9+mLgIX6ZG/l0rTc5
cPB2nJlvPy52mg4lKj+nKfMyR+eKbr8pPtJtD4VxHU6cgGYrg9BDY8zS44cWvyCn
PcyKwShX65HpSImzhwS1XjkLMFN6fEhCMom6M2mdjVxllUK/3f2HyJPqc5jCpm2/
xTwfo5DfINlB3h+jrocdteazsJEO7W6CpZvD38f9r0Vp/CtU5KntMLZFNyHPr+Sa
sNocViOeAsXOhWvBhQuXeQ9CRUJH33L/lq5pkeo+ldw0XDuaKxXZVyXCOTzpp5+S
bXGKhmhoNWvLqkHWMhTC8AqEIYp2Wx7chdaPING7DoAwbVz49UbL5BPDBPX+Lgff
7dtS+ZDzHNixSeY1qJinhKpPNa6WZidXvtIvx2cE6WKYCMByoOFQqiDRtPQukhsg
BGKYZXiviVNJMX9J/CBQMBrQxnXkasOPksz6gs4Kx5gzlayS4PFTGHVpqd3ZCAU+
TfrkvAFHcAkL+aggAnB/ltUeOVnwzxVqeC0MtW7+GG9glOr7GDabhvr8rjYapIpN
+/PL0dJL3Moc3o6mJY2wmIXwxircd72Dd3E8duBcwyYtx2VoybJGaz9M68kIsCbt
CU9XhsCfP67Yy8UPtn9hkdMrXoM57gx+uqh2+OZBTaI1UoM+3g27/I+J+77lLUnp
YSdvMN4+5CU2/72PK2JntEfw26iqEIHxwPcZEHndTKt6GZpnhoO4MMHJqa9jgmlU
8cgASMwwM6Xa9HAhDD+crrxr9juaD4PBiOq3lWCbLgA4feHokMqa5IRf3dwj2zsC
kM2wZwo/BpQlfmVReUsyu0rUqWDagvwociv8UqKRXJqCb8X1k7HICcGuSK/dj4VR
N47mguE6QCuq5gLweVPmeYNgM/0WVBGctpQcXni7NZydG5LfixRbDLpInzyxbtbV
zE5XkqFBvZfDfqqpeaZHnAVMmDMYkvvSy3y+9kLEC2DT/h5cl5p5YadTL3bBF24O
sDsg3lo3QYkvXke4DjxRDmZUulcAh+wxRdRGEP0D8B4xI094kssL9rarG5deW9C6
maDBbzpKbXHEx5vXocSHua43kE1FGzr7GukP16nkL/Rf8Z5hb01j3396nx6+Q1wj
k/UJ6/SAXSqoKeMPX5wykDfPafgk6QQmF1FVWGeM2SrTfSEEDDSElO1wzcT9U+os
7plAqr75T6x/OlMVmoHCJanZ8XjXQVkv5iUKp/iqAKdL0K1Ir35FSfLPHKq41F8D
x/tM9EGxC30o6Wgtd3WysjeEqpu2hDJgYy/pstITjga8cvJCdiKQ3dDBhRLFiqMP
iq1y0NTVFSGhc3y5lhZKLIz0wZ1KPOD4ziwNgHbaeq479ClpstP5WrH1MZ+zj5No
1ChMSipNFQN9czUHDZ+N6+L+BDmA1ji9UkrqPxBW6APXnFRRjiXzhox/WqQgf+S2
9yR3oDEWFqbJP3HauUZd8RYahrqf0pfYc+hZTI4xEVLYuav1j29qU5qodiq+2O7c
e9XyhjbR87uKhLAkDZqk/ogUezJLEo9cKQf2b7c45NzotMjttvnayaRtgCeMbyoK
E4RrndhoVsBuCtsiCEmFvMY/a7z2Pq2J+Jam6h/u23WcJ4e304481yFb4NSOxxhJ
Hd4Ottbt00B5Wp9Ubto+ecB7RpMdNldExFCWfk5kbYb6aWyH8YJaN1G48beFnVUh
TTMf1Y6SmvNBxitjseNjTWbzqijcTSLjmYr/VXfCGEmw9SxNtpqlab+c1mQFAOG2
fuLf6clX14lreYjFzWbMC6kHs3nNVtR0HdnyeIThIoiPr1gZmjdyDbrowzQ9fI6F
VzQSsWZxuBYdK8TmfqpGPN+aw7IflkosKvCRLbhQ5knqyRW13YVimY40IIRPimFq
pI6uHlEEvLbE93mG2ojwOFNwTR3ctLQKkNquZ2WmDoCzw6W8WJsQ8uLGlcHGaVbj
VohMrPnRfsnReG1jIRwxOz8RFxxy1i+5bVP1dPwhiv38Hl2v62uN/8+xHuxxXFgZ
KGCXTXJayaE/n0nP/fwnlUGWlTFC3sct7VjNqVjMRbQ2iSyaK3B2A5fYTg0OEyJ6
Tw3/c8+Zg38iUOX6gCw6Oh8PIYKA4n5RY1xx/bvHTkK0Gm2oVrvMATlPLLIef+SX
FDlvSE8mtSlHuTX1IeksGis4kfOrd0B1iocEAjm622wdz80D5OzM+uXO4rld2QG4
xN48f4NoqjmgUO7Zp1W+VbE2wGZksFhfWtifT7ubHyEX/ELYM+2MFH0zU8gC5/2A
zA6PnmBg4RiImFyMQ9Arv21tPIcZFqYjX1w9o5O34qOg2BGxrnbPsXiR5Hv6kSlr
Svp46CI9t2bWhix8QNuTj9tAl6gu3NZ6vGI7+j4CEvr+RKolFrKKyFxRi4KnmUlW
f469YpZ29exkTSfWmsG6OgcBB/sosgDcpzclGh+WLyb3yjzEOfP72Ga4UEPfoHRB
+AwVdiUZQByqKpyu6kJrzBoHE9gaBEW7a1yQE0pzhN2hKPmklzP0VQEZbfdq44gi
AoU9xxjH3++byMc2FT2e/Ai1qovwYFhze7oEzi2kYiXROhVse2b3zDkZtq2+WCLx
1oc+cKapvEcsFqXluDtBjxr0aULiqS5g0o8YjTG3jzjW/QgM+8+0JvBbpO8aLKna
9Ph97i3v9pVuuHKsPbfl0BJjAuzvN16lmMWAJVJZ4SzPg4UeO8acQzdyMxegIAh7
oeIKlVs01WYv7T78/1zxutWhFv34H1m4OLUKYFDKJE8MBKVvQrfgOtprULsTl2ig
mOIKhHnL0i/mlDppXbNP4DQgJ1Us6uwSZhbzsFXzRQ7U4/xvbR372y2Ei1gP3T4y
ZYvTzxf4JLIA3IllK8Jx8EFZgkttYO41cjh0hUeMW9pLa4Qs0BLub+q+mKb+uxcQ
QetvDrJdoBPInyTlV0i6J+QIMfF02Cu14P/ec5AIjVgFPyYNFJUYtFetha9YXP7r
2v70T1eRw0apZmZ74TIO0Sp4Rc6VTpW7LuudD1YxB6JQMZpJT49CAKqkrspV8ik5
rL9XFPLYUuORW2PYDC3mt1jHJAjlL+08rjihnfgpQuuw/jDN4HHaDBKTm2cWIs5p
OYDfxTXS3HeVjilaGCX4FQK3fFd1KPaezDiXiy8WjSReyl2KHOEqzhjc3Z1TxLLO
85qHdWW+Cil3auOd8cGoO8fw+Q2C8TlJknQqZLvw/g2IGtH64x3G+Kb5rtZOSgcN
b298cXhBNQoWNkqBrfo0u6TyAbVNAQ4hkYvXGo9DR2W+NzRsypX/F+dDTVkHSOSP
ZKBcNSyvx57S/1Bpl/WMsN+wcoMfkIXeAdcS0CS4JwU+TJV76QJshkApaudNJK0u
Kqts+D/jJL5ztSbg+Tn5ZW5lIvd/YlrRkoIEbxBP/S9UwltK8uNv57dN18D4jEKi
7ns6vA95gk5May/lcGiNMxx4PHYn2QEenPCZ8SPjuQwXvuiW69RAsI4h/efzCqxp
mGSYq5p4mWyk3eRVaJ40TlAaWMwh0/XektT1h7kyMvM8sbh33vI8SQGAw7A4agjx
Lf3K3gxuepDI7K7G7JKgZhn58f/xiczq9WCusVWoRxi8rXc7xxtKeCC07lfqCLKV
138kG6j0wyDXrJQOyIEbmNTIGsKXVDJDF/UNVIDj/JHW4ADFYB+vU7Gb0Cy0UuPJ
V2FJHMHwfhrWW9ji3miX155eQ5DMJ2R3If9PevLnI4JdjoGTS9WkY+Wy/BiekcHo
qSCIOM25akjhgIjOZa5tsDzXahfX0zSs9Ck88hi88eUjZKlzeZ9TMWfwsT5BOWf+
QvSORmzKnkrnqwgS3I6E2Iqtw6uXjKw9/xFm7+ywRtxq5BaSy/2oqNH/+L++PQTJ
xxuM9/T01Kb2c2ZJUtRVVD/sorbZVRPWQQA3Ngm64guoulyLBO3EkskCqxK2uFOP
aJy0LeWt8zKznMuvdN3l3z8JlcFm/EFtyH0APLLEQSJQ61DbyBTvY6KWJjIHEVsZ
A+4nQs+bkDStCdQbLJC7BKpJ1gJPwR+mlS72/tTPLSRRvJW/1nfGt2U+FhuAYdxD
VbTMDkTYT+5b1ZpiJY5/e0k/QFrn9djTYCsYBCtXCtBsz3i6aoUmryP9u90GKJaV
eKZPsjgxdPlpVxTqQ5pBQtmdYI+SOpnCCpm7AX85O6fqtx6I1emzsSz2rwJsLB/r
dCyfRYs4yFfUuAe/MDhIK2JaE6K0k2/38zNv4lpAUTvrmyZlFNr5wke19JQBNjVV
LZt0vmUMMq0jqdcHfcCR8fQeR1/7EyBEfWkG1rtc75k/3bAaiE2mspLezcEW1Ci5
nM7TXMz0q17kMhHCoJUloe7eXdyI5/ZLVWD3Zr8ZO3SJvsr1wX2Cir3pXVM1LuRv
VnNhyTR5UAMRR5wYGMQ0KJ3tSyxjG9FzPS02cCm1Fngs8Ck4UbTczc0pNcy/rDrh
Ie1dqHi6MogYJbuP8EA6iY2aDjCKtfM4pSPmGRtTh/2FO6X41EU8zZFMUm4G95TH
RfuTh/Bdoppidk3bF+2fcvNSv6ZYqaj1qRK0I68/zZczOPZqG4f6l0PdxatRT/g8
EL48E9Wam30ZGeU2iBPnWZvPrJEs6xbjqWHvkDIffyE6WIkOB4IORaxVdtHGuEH5
SlG3PBeq7kde1vn2tFnx4Ir+YLf9w2b4OSNMMot5L/N2wB1WsAk7oT0M+2krPxkH
tnT/xykoRip/tjys2EIxDmSBo8OxCc2+Mt0bwfcEDV7/Kuq0Yd25bMrMrdDVohT0
QHrQbTB7nf9G/V5zc6WBFn9zK8As5VlWPp8vErWeuXRSZd5awVhoQYSSlvjVuo0T
5h8eqQOrx+QRObEHthOuDX0t8M+Z+oowmuo9x0XvCBF5Shs4e77NEjGXhVGjUex9
oFmMDyaL76PT1Y+Cp9bIgsEgSjtnM0rOsCTTrNbgxdCNcQMRWtQsMoCDT/Cbzohk
M1xtKxvbSdZIGt4rxHBE0Z0VWh+I2btsNugEVOFDoqxekamrBcjqdMHB4KmjH/1C
bvvEWK2QlevTiD7/ZWnHjrdGFls1sHza0K1jCP9bVfeZX35DGi4doVbTJwG4+Rb1
zDZtokmUg9b4cADMRlzOYXQ9MvEF3XTolR54BPovOtZeM6YegmuiKwlIM/v8SRg4
n5WgzfbPckTBa42hexOdvKn3O+BNFCfbwAOGGkaKiyszuffACrFNGzIEygWQw2O0
G2+xsSkRe05Czhtws051U2+WdpU/7kxD1YCzB4UoLVE6BQpFo6mQKa0s/VIhaXee
WBApC18soxDqafGGRJkcGQbQdnheP6NAH+T09Kdx/06JJxzG3VO5GBpwKelef4yG
Fa/hhg1ll2/eq4ekTiH7KjQ9LLig7IXrZ70MrDRWw1ymMpZzhRx6Trg5QdbpQuWV
mPqdJhjCbrVTtI/8cpsY9K31EcSBbjP3v4HXctAHhk+rRUWqcKMFqpErdASPssFy
iOjtALmF23VP0SX+PlNyCtSY6cecZUHoVIy6uFF9WZvJgd9LP2qUfmjvOBF6Lfyg
lVFegFabvKUlLw6AsJAIl6qqRSddOcOOngivsuZBABICoTlB7myoh3WjBCDaIhPA
F6ByPaLMrobccDQc+zyQ8J6cVPaYdyZrYJY63fUcWK5zqYKQOBKqJZ67n0YEfNxh
4w8gEif3R+Skc3j+aeN9YNdODaCHBImW3ie5aQ8cD3Pka07IAkRmqeB8wcLXGrE7
dS9Qh4W6JB1Y3K3VxLHDUcv0rgT65j7KoiBzlFx6W7GScg6uIPmPrO/cG2sGqQJE
8rb68DoadUl6WBOdNsQpGPLht7WU9fRalu588Y5oF4RkxY3m/w8lYgXoU1u9GW5b
kpcNTHAtg1mnmJEhifGDbdQwK7zd8nELy3U+5IOdOzwKvy8LEPDhly+FQRVvatk/
xy6sMID0A/rBRTZqRjFQIUbUIr2RVeqv27jdp3P5jul+kAWPiEUhTV4LMbqsvrT4
A0Viql9tjMe2xgSF8PWvip55WUY4UyIrdLva9NcRehk75Q4ILXGI2SNNjyjuY+xO
V/IHvaq1+4cT4/BQWyvIs0eVN39UskEg4ufFbvip/uQN8iaxsRodofOErPRPDXVJ
y3S8RYsDcc7Jok4B5uC1pGBcvPiP2I9emdV6ko/h/Gf7+su45nHmK7wqLu7G7hUq
lIft7ZkTgNYxHx9sxuPlwrDnaqg3lI66WLSKCFJErSjNgrjouVnahDiOfHWGDz+r
lMGQgTl5HYdpnulsrHGWTw06aGZoBWUiU4emwHn8J7Qtn4iBs6p+QHwEmejfjgJk
jkjC0gQHnBZxCfNTeY8HK2uL/6yqKyuuOw2UQ2f13smk3MV3me1VZYNmFZkjGxqj
UkOstktGETyoZWpRIyx3As5oEA9rExnE7zwlGPqRL9Tky0gB/lR5LTYAZgSvIoV5
jnxsVgOUL2XB0H5iF1tBR8K49sX5kskPe0YOBwZQ94qcVm+2FUIjZhD8/DG044G2
gXFMtdBICknw3qTUd5+h8aOKCAEsxAbeDJOT7226NgR8DQedZ7fLhUZWF7+dkpXP
omo1fZT2bswi0mHj6jc+gROSQ07LTHjv6LMDcF8zVsPYxbfZrkrwn08qnokG0REx
1IEyP2h6k/YociJRaHiuHwFd9eYThxiEYSVPtAemfpnvg+KbxYdnB6irV9j5DYkl
H3EAGwaoHmHBeFjeafMqPurxkglB78FgZf2B16/G5UBGIwyuz4up5bHcI2VUzp4H
dLGrH1YHukMxcQ/QMtbqWHzf6Y/TXdth2z3FkEMnX+zM0gTy3bB2ir+a5v+czzaA
pzoSn7WQgaienv/N1Wxl+1GkQPe5OLa9xOJilaG7o/zCpDJkJjyHUMRTiqg66H9L
aLu40vQN3uAgv+wbZBttJg+EGEGxUKR5dW1T+kYSlg47+FzklUHsjxgPL+CQrCAo
jYR1rsYzVovZz1w3W/h80GHqXTyWkSyqIELtgnrOl+6AcZt3qhDyfpYzSq1QWwSr
wD+RQJFxCIKlQKQhiGE7DMVuhiPMlZwur5ppbtojC0bl5yYu/xCnNfH16QdqCGyi
EkYmAvd8b2d2b6W0VyFu2IQQ0N3tV9WMFHRR1mYghMWlVmvyKtxm8I7b5lgvqqU+
fUcfbtg4yqhTYxNHS3zMcMjxOl4LffNgdYDBdrWYSJc6ecOTtD1xjuhhF1Q3eLkk
9PyTMYsTaX9cT+KhJzA8ThvN2lvlLp/wKKBBSiogRlycXvqiYIBQffNuSAWIz2vb
PxnycAkVBp6rcR9LSf8RxzhohWb+O0M7w1nQghdS1eN1ueuQgxS59+pIhmOXKqD6
+zHDDaQ8LRnCmJUY5tIxt3yOQWD+YCCZiBiAaeCPiwOlTH3HEEgzdv4RN5yk/62N
HwjDwOz36Gv5t0JKhxYnZNHrXgnv5NLUL8/OkJ0uxIFZBb4CwzEq+XWLjVQPC59b
3NorVwjU7jmwLhJfJPpPJIUSlqi+h68JXQQ8QiQMiqC1ud/nRT7cPYv3uXxUcvHL
mliYe3oR1Sa5m0w/TdFM+YSYweSwT/SyepaIr9YqhkMomX8+HZwUKVAA9jUAWbBW
33k/eV3/EUNZCQhxztNGFbXVZOkEOXhDx85z9ycrEs+vkvl3FwQTuFCGs3521vWy
zoaonKVu/l4D3TRP0I32tSWzJb80dpwOyC0vKc+zNfnKYN1vKhL3JLMXaOFKM4rn
lLi7iUgBi+XcwEaXq8JqpmxGw8Lm2OEy2+Irm1SVKoGUukIHqMly2Jjra6LrfJIB
BjsdvDdFgsxtd9eYrCAs6dJWVDptLMTkF8VGP5qozhzaPJ4qfEfJhl0W65a8dvDX
7l3i2eUAm37D2tYrAr4atzB6HazJKu8Afy0paQCxnJDKgKVoH1CJo22q7FiwyjaC
wroNR6gywwVV9ThmjkFnJV+M7F4P/tQnuSw6G4OMeewr/NT3qVtZVZPv8KfjywR/
27YgMpoFCZzf5FwuNgy0wamk49Ybmvr7UkggnBPWBvoFJKjfleL0bYpyTrKnfjb3
YYEP11amB32xtB760mVkO60sZarD1fXdlS8wm5xK5F/KTs+bQLqdEjd6043RZlsV
f0ZENp07tNJgdTysxbE6n3wgYoEyxJD+rWhzHCbyE75Dn1p5ASwFoEdmWhzgLNsN
9i/uEuogdFrWpcVqprazznzPvAtEgJYRVLBHtzEXrlTHy7iIVQFD2kyfpLojpm8w
Agx1b2JuhwwTNxoN7hmZys1Liga2vwQFMUc25e5Mh5PoFcIwtla5R8Vxd/KMWMNE
62duU0moHHO0K25l1MlBcu+WmfH7c6xp2rEPmUEavDLurThB0W+bfUeMN4of48dv
UqPiaihJaG11mqOTrTGPyoPu6RQc6iqBIDPpZyJIfLDfOAe55n4QtiQ1pg7BgELP
nJ+dz2lByzPhb+E+xqwdi9hYyAK/uCwEgNkc2UKEMrHA7S16ESB0zDLrXDFrRuaa
cv52DuyRqaum0nL5U5BXvFK+WBFxJu/6DNrUXRtwOPu/k3OWuoz8jpuuOMzXMGZX
WPFwkJXgjli7dYg/lZdZl9U59rGaXBzqINJUuwjFOBZnQwo+APP/m2DxGKiRofhz
bRFSIWjx8TcE+X+AzhGypM1DJZ18SBeJ76gCvd0xwUuhiy+kXC3/L/6QrYr9tjln
DL0iknPzz2u3EaL/YR/0z9E+I9JUvDTNdINXBGavKR4DuKU7YMwiXsSuGEVZX52D
s7JeD5DxlCmvfSBYC0C5T/kxVI5Y3QTJX8QafJl/FSjvZb/F+dKu70ol44UxExK9
GKujKTJw06xYHOIOTp8g6VFMlEmUfOj+ZjFj9gZBIQeW15IpXGoldcHeLGMa2j8y
5mE1OUifdSvlJMj9vnYF09YdxADpeUK55EdXrm6yuOM0nKh6OTReN4+C0kDyTc02
XAZ7S9yO/EOANPUDQ4qq+aV0sYAPqCDfjrOC4lyn9bpbyq0mTUUU4tHaKl+Hjakq
ru1r4fljfkDrqkO5LS9OQ2Z4j3cXuUPF0fX4CbuUJQligP5UNPueim5COeOEe1xy
OeAKJaT4WZu1HO2LOkX+yuZfnvWHryhOFNNvkAkyg1OU1pruvZb/WDmEgdSbP4RV
K9YIPz43z5FAcagQCU4LccI4ZvDQUe6H7aUxrR9ipCYwSX+qtgrS3mMpgP6NYakv
nghCdZx9jOAy4MZtTaZJkPzCUdJNHfdtjTbfMuNWM9tPLrqHKk12BlxZnkvMMFG7
x0NrR/6EgjBMeY0KyrFwmNVNlOR4fPsh+L4yr900/dqhjtjgUmRhLffg9PUpTglx
FPSDGZLCL3VAdx7VH9Ie9XjOUAqnlW3+CalRkIlcTjk5WGYplUmV1KoDjnhARnWY
sQVaUdcqKFH14MmTAaoPTKG43DraVfEKMip0f+pbGsD/OzAI1CCm8BMfNLb1R/+I
gYAsObFON94OF1mD24mhf/jGGXSFyWfY6UDieJk/EyZ+zmgggdoiP851Fk3FTrbs
bLHQ4ly1AJVrVE0oUYalRfvF/t+iQ/+uNiLaW1mgu1mTrCXIJ/gSycJ20+o8X7N5
mUKg5qyDtg7b91esbD9noxgpNtXNAmyfVjMLNH0DcYDpDgDDWs+9MKNTH4iRsQdx
oCm0bo0UTjIPTLQt4wOVD+rF1Cbw/ONefu6oqI6jSDgz4LeweKbU+lnSgQXbzO69
r/LPDB/uqetKgSJTAfnmF9sueG9AMnr7WNB01cig6/I4YdAB8YFm+G29qExTiiHD
AbjtQDn3lxy3uJE7rxGxZ/44xf2HhDUaoA03ZU7rKlsxuTBppfsJ+ZpU88S8uMmk
KTV50moT2qelcRlnoLuAOZMk0D1MAa+qfPXYWHbD87mVSWuwaN/zZ2AI119oyLIt
DPTzPJwE7UkGet2P4pD3g7Hig64c7GmaQlTl7Re5c41WSFuY8xm+XCCFROxzGksE
o9xRO0IXFd6ZxeQu6haDlyYB0J0vIRVRebB7iyqEom9UAY0yIObvKH/RwWneFOmX
vv9d8wstHTpsmCGSjpvpVIPI/JoiQop1xVmAETg3TnNBBlyRl/Nfzj8rBTg2Nf7y
PIeTwiRO3oxDa4Y92zcF4fN4PZhF0FRgBdN7arg0d9FPe62LjLOufmTomDUDS7/e
Vp9whLP88eFMtqTlQjPLVE4v85I10VG/3bSByiDfIcoVF0rZlJJM/j/AZpQ/rfL+
qmq6Ved9qMy29BpBPFI/fiIIuQXt09y57DoyxtP/0YVWIZw/7HEWbFGmTnLTzqS4
UwXM508d7eIldQ2RuuoMGMVlvX3P+0JjDCjWs6mFakM6TIirnQInAunNoLpwNcPx
q1ATI8Jgj8SMsx9K1tYymWwZ/55Hk6LtaFi4NJj6gGTaD4yW02FXF4KAB5sCAoq9
5fXo8WOe6i9AEw/B9pNZR4s9MxFxQMmAtP22Jpud4Ypl2Xr2Yn2hdtx32cpmtI8W
3SGjpwXs6i0TK+iq17XC+rovqNC/iMn0QUG8ZI6yNso4tlbOq+/oHCAeSTXDrEHc
MsVvz3IqrQ+mMNjDZ13BgJRme/kpwIsH+EMLvgj/3NzaWIlmbA1zG+q9Kk4ie67S
AGS5zW94QMg8hzAaSKSeubOwpBSdGEL3SWmqD+e/p7+HWQxI+SPVcOo74gnraUKa
PLP5P6DJfmh51YCpdKbYdhPtAAJsGBmRGB7GgvM0RXaFbyhRkJllgg0RW8PRDNUu
BIUhU9Kjq/hqzZpc5Eh7D8KSncYSCy1C/rY+LTtQh3+24TQpGAn27XOUL11ZDVU2
01j18K+1s6qnW6JNoGA9J3aplomF5ofbXsmwyp+lkBCzJkIhY0hD5xRD+T6STIqf
ING/ORWKTG5bLK4i2jG8285F5eCGiOnQfflUPiGuMyV+NACbA86yetlJdGcK30vV
kpbsiALcY9oMWuYhjeyA+Uuw9s46v517SJ77EI9RzLgxI38+kZ8Bq3yM8EnUO0xg
RWTYPZVs/AdqwYWFrBFN/Alglkjd5/UC6dODD576Ll0kPQapnzEdhTjXLyinojTz
lHAVYHcFqeVFVexGkb71M057o0Q1zwJ/0mYjRiSJzXBqYL9rTFfuu/1DzdF5ALQk
P2QScdQHFZBNzO46gAutw/MKSNYFya+cmS1BnC+YpdsN8lS0UOeC/X34kD4eARML
tCkTIpfrpCK9leVxO0ush9o51xCMm4MdUbXzlEb9grq1Uz/YztZfIGhkeqJo0HTZ
Ko+QBSoNZptVptWeS3HaSpBN1D8tA6VfJP7NxXCkzvC9C1EzGYwIoHfKNLzfeL6J
lcESckNYFfkV52yIciWdAzOexBu008ppdlyjRzl99TbrTbQPMZLENyVwX6al3GqT
cB58d4CQMczKQPZlBfq9WclX41NPsFDZrhinc+0iscYagtQZI7sn1jQApK72tSj+
dyQZNa3L59gsm46a3ZDKH7wcqwGMD7RbKGzoqWfSxbKZrXCL0UumYq6GJo9i5Ocg
/o4ti1u7QaAuDrObE+oGntzc0tBoI3vMEdz4/nTH9ywfjr0gzInlBHsUamKFa8bt
/2ymlmkUNIOMt8XVlKcnZWMF5uObgnEs5UZIb6CkR9ynxMRNxK/u42EG7rCBwDZR
7SE3ig4vet739MZGJ9XoMsiFh3OtCN0y4gyB4YySg2W7l1w9R98hWXrkGLB0cFZl
WoKnIL/U5cn0iYky+YMm7sy77AlR0PALGTQ8L1TrkgQStTyu7Vqu/+SoR25KSiPg
roKKNCRXt1/AzD5s52OX0DOn8BgMDmQ0l5r40siACul4Ih9n+oINgk/joJVBwlJ4
WeFGn26J7pbUWDzzubMXeTdxhQDty2/3C6lcseC9sTkadD249LwlPDCvYj8afntS
vnwFFa5xXh2oCiXQ99RF0CZtL3PbvwUqtgLgba9n86FSs8Qxexf0n4NjLVV41HgJ
SxWlvVvt13hrQgqthPSbbsdeORsUgwMm31r1DM7rVhCTsyVCIo8pF+LDQqiJSnCj
pNEM64Musyh3nAJVMoKF/nlTh9qwYjW3i4pJW9Y26gnfEa3Qe9BjN2JWlQwZ1uu9
lnjSDKf56TRRVuTNbqcvV9h5ZQDzvMkMaC/FsMM66IapR7brjRtcpLuPxguAQnqA
xlDILzz3C+wiRbMAQNxYnLt25UrmxDw3eB9X1cH9TM2KmM2cUMbAsyXBRceNElt1
wMDg1yxfVNnaPgmkzxxb0fbyrfGjPMhiDLVcTSqHr0W/ycNsO/7e2FQv91MHnWmu
qsiUq/GAmwjnBYkZaC2/VwbSX3+e1LX7sO+px1BXrLZ+54vI7YTQIaQvH9bpQjQa
DUp0xeqO1qj9NsLIp8rmDTx78inVfKR4Crvz27CjNzdzJ5vIQf2SnkMSnBAgZOnV
BfhLE5Pz4/NnaStKavlnlBPAODrkapGgGcZSjYYcdN4ylBdDRJcZ6lGan546hGA2
8zGIa5wGhAV3jXi6r15UQRpGlLlopW4rnHT56HmaK6rSPlKqzqq+I4wxF1NM8QCP
SH2teKhmIIRUS1mGLGpIsexloyy7ZKhhis6TiVDT+H/vL+eaGRK+kLFFrR4AQoB/
QejBhAlPuqMbfsKn+JMn6BBIfHvcMiBeG8rTbTeV3KoL3y9IJRY9oi5/LX1ei2SG
RbKq/TWFAr5VcMeYDH8MJI834C8fOx5FErtBAvvG1rRH0FQOQzV2oPYg1ZA7cNm7
wB1dq2Bcaw18KayMOdCsjmTlSLmgagCshU/8e/linXPZBRB3k2UWLhESdz4O/mXx
4qQL65aiLh4Bv+NSmYwigHGpIxSofpml1tjICpad2/h1yzmrtZGEtFGFNxgdmjpT
Ljc2XBMkXBNRT4F19Sv7kTnCRbUMCl/kTPjbjtnXCDT0YGm9PMndEmTRNEEYC2Zs
dlwCuumG51RXKEU69gd8gk808/8gn6dhaWtuaMss7Ea1pzA1Sa3qcF5aEV32H692
lm2NwEreSFy625fhJBAMvjf4eAUZWjDSQWW/dyaQzDzUWpSaGtXrWLw3lXdDARsO
Yr928dx9Gmdw4FMDhML6bOU9UKYodnoCG6CJ0/Uk8x89EIzKmRUX9xJ67pXvc8w3
NCoO+qfiYBDRcwYDVmSHcZ0vCGL4DUMlTYP6D0wK/Q/hCp7VLszl707Dtc8PCg96
c9PGKVdgAXNMIl6Urc4EEvVAHohZ25vv/Cii6+P3n5jljUh2CmooCR3iLgXi0iJv
TbAmgcWHr2FiTOXztK2cdblr/XZlfaQqMj7aMzf8HgDUcvbaszSY/VYgO6XseJlt
SPSfPY6SeX3fBDDRaNjDlOeRYIFyaLiuzWE9sb/T+tbcGPB8eiO9xGitdF2rnvyA
i5KhJCROzglEnqmWQybm1AsR6hf3l7KG2vsiC4Rr8mRsc3BIHfhRH0cOgtr7B/GJ
pBweGWzs3Xp2qkM7cbC2UIqcWxZe0wqu6J/HIVxDsloZLAfGyUQVv2n5nhc+ufw/
dPbxM4Y4ell171Wu9HSdCTCaASVyCC56CHi+xu3rf+xYzFbrmgcEg0Eo6jhhaXeA
rJ6VqRlDMW9aqipaFUJjiBFhudgI1ykcOVt/z/KXomCLSY2HO0wQK/KNiMUFDmwY
3jaOMO/tqcAnWm4tvVwqYhlb0KvEgmdCwVxUPyU02srkXuqZzQ7cQgrsIXyt47av
Mo+h5ra+6gpVbGwiK4PwttYJNHkSzNGJia5fSXo+LaZCKJLzsmNm+5FF80HH8JOr
V8FoHledvm0YqwwoUQr5vGkkR8vdQhiAPQoKR0IdKcy+rvIeXy3C41QUEaxn6F94
LlAVuqmOOnsun9UfMjbdypQ+6+D1CDYbjJXjbdx4jzQ1NXB258NJ78NBT/fZC6dZ
I7SWt6uYwQIWcV9oyG7P5VLK//DoC4fpKQCPLYH6AMH2ykH547PYn+T/JG6O2cze
xuOnOMhhVw0F7VKB4CUegsPyB5v71NGlkhopyIrVpvOX+OahkIIx152+Q1r/B0tI
nfGMJe9HXjZLl8eebcvGs7Fjz9yDi9FINXq3RQHON0jhAaYLeUzPez4Q5e3NB/3s
6JAHsqlVhBxMuFswT6OKfE3N5ii4Ui7rRAjP9Ente15t8rz7ZhVtLoBULjVrrDe0
80Pq1ZXfMQ/7nSdfPEPLWSVbrd12LiYTatQPCiAYxiN65sqktaZnUSYpTON9OSwm
zNOoys9k1e5GT7E8lvIeamBTxKJKJZCgpLZhoOehzedxxF4/MRZ0FKHcLCdm3AFy
JWlOiCvGnP21mwFBfda9uSlswujhsyH9mUq+BJ10yuE7Zz3UlEIeppkKTuOBEOoC
jzXYJqqIX+9jrEd2xeoP0YHGTOueAN44+6EPPwDZHkGqIKJYC9UbP7zfZxaXXKD8
+9aie0zk4DjkMzb6psdPCh82bRCao3Bgf464n6xlCJ9lesyoCrlj3XY1aJ4ezlvX
t/tZdLCbO6eM08GvRNJ29Sl4/QsWsOI3twdG8NqWHNE78844qyXQYI8ytTCu36mj
RXvfOWaMiahgcbdsYE2GIccwwOdm89Rh188DDO7KGMaOK0ufUW27gshlcn9cV6W4
iN3KxdZkdvLq0jZjRybReJP9JveHGEMv0r4t6X3eGdsfpnj4FxK2LTW7XJf+RSNd
SjN2FGBxYWm/q9JsxsBT9A9JCtSxFTY/uDi3c7n/CAf3v2TYB2RyEvVWRH/MDwtV
NIBM1ve501c2GAt74ie5g/ggZsHNTW15++AEL5LUXPJ95Khj1xyHkEKNNdTBOQIt
9ezRZqumGivmyYH5yBpm/C2ftiFj7ClMcmMxiMAg8KYoZScPCcyKRLLGSlDQrPID
jcEE8ge3haEzo027nNwqOcDl71gV19LdRXCXNnJLm8ZuxmfyHwNPvkEhFX5ShRh6
snov2wKHoIYfYmfK9V1q2JfOHhxQm+lIAFBLRUcAg/P9R36F9SBWlAopSc6/CMym
LuHZQ4ffKmboa9TAe0CUJ9V0sm3dLz4Yntjly1KWtVzscvppzocwVwigzBFyALFQ
XW12xIMsj3nfvH/vq5yFSoJ1ng9D2jJQh38aGj2vqZAacM4/npaHoEqBOaG4JFcM
NkTGS5fWeLiZYQWkCTMpSv06QqOMFVrcFss1G6BzPycbnDmxWnTm7vD3/mY0dHdc
huewqjZynMvq10oKUgJmbRsRE5QG+15X1Bbs0FO4nPByO5ypFd1Z4190XzA0s4Oz
SkOPjUb3EcqcMDhdhP+6EHwSrTOSKaa8A9rQ2QeOznFpjoiyZLnkAU1g4AhR3v5T
c7sZz339sYOHfnGc+vRmG3wVwYQ/l2rjGEk1oqp9Sq8ydMbGaT+yrJVQ/Pmcvo03
Q+CXDsuV0FwbJD/KAslmCk+YsJVmdZmlX1DEBoA81XAV3mLUnTz0SMGX0Es7K2jZ
EWG+oqMl74l3veBq9mJdV5GYGAVBnfmXsHE2MtMekF+2j3AFilGs04NCfJ8WWGB0
xzRmCeQ3aKF/Qk7L6MiTbfVuh+t+3pATw7rUjmJe0U/DN+wBMQ2v6lEfEBCICpVb
QGHQ218Dcvt0eg6ydk2Jg2D+v7rH7OvsPmcry27TXeKlhjv7Okzvg3fc99tujdGl
tot2ys7spSeWXA0UiCnp7fq+Vu1JwLtEAaJ1Jp66325G/kZ/0feFHQd2DxouAZiU
QxDcCmDA88/5WiPhqZ29wiGXc7q/YXNmgqj8ScLbmepic5PQxacxGKJDobElfaCg
9Ta4Srl3cHWab+AnJlUNJwhwwNQHg8H5L/eP4yL6n3NLawUa82+og1oDQWcWI1/2
Qu4P5a4Cpl4GgZyZBY5ujxg4+Udyi/YWjFMvXlG0+D3R717Xk9Lk+x+UU9zDSUDn
zt7VZTrZbza8oKPb9AikSajQzKCpcmfhKf0Sq3hPlGMWEe7qh7lnJArDlQ+UgCDw
3WATDW4Lbrw9Qha5jLXu2GClXRBqsOyqKvlrMDponCWAU7tvt9kClnUREn6G2neK
aHmjQ3pi2LUn9ADf3CgewIrEU0jn1IEQy263rWUgAlDZzhDvzRXmCYgN59GP1jXY
zNi8Udc02m74B0FrwOHRUdXgSw0umPreYtYQXgx98nIXgpmxjGC+yPI9NHL3iHRk
g12yzKGn+uqghHYZjjLkNmc1wGWVQLENK2ybrNDPvIPtTYO5wq3o9UF5fQH2Vt1+
w0tAcE+8GV2GToT20g2rPtOJzVYLou+cRjzMynOkqs7pXKrnI9rLJplrPOS4vmPC
KheWp4uzRPuWvnQMUw6FsLJxFCQQMdWSSAFM+uo1KuKjOWlpppGPYHPFH7xxZFsI
LSAnb5ve/mOGIwFdHoOe3pcvb6dZXzSYQWE6YFoovQWOte0bnGyGYl9kcweRP1vR
S1Jky2Z4hKB5R62O6xJTXy+DXfbP1vZgwnUkFbNimn5kb3VaDrK0o/b35nlFlkvC
WZPUv72C87OAQ7TKxEWpjz9jCpIFJIy2qc0p5krL/9qXdEHV0yKGGl6hFgEb+6J9
XLfit57jciGST0nyNdmWfd6idAVwLzErPsvn7BSQ8Phu6oMn+KyXyfGch6fcA2As
WiKXG+tJ6oWRVrShqMGtRpMxZ4MnpQQTQFyzx5zYvQng0+Yv78cdRMPrcughGZoI
DGdrVPTQ1Ot5B/UT5felf+bcu4kslgJVXjERtDoVSml4xzpIlV1D4uf7wpB05GW1
5Qd6Qsx5Q+4I8j2qSAaYc0t8clY1d3/HXd8hxiqifyfLND5CITHyCZLdFnt+oGgC
7c/J2pLV8AXplgFpKNbh2kzJxu7o2fPIEm6hwbVbBwytXlZVSs4Fi47ioWc1Uz85
xmc/UtwxndhN0BggQB75bN1ZEIRX7XRXnzjmIaXGGakHGaNn53SKwhrX3xh07CYR
4hFEgkVqAv1akfsnUapczivS1wNrGh6oBRo1VnrklrqvN3/5izuDLbExgNhUp636
7xYcTUQPVHV2uM1EJjfPrZ8yUDTA26XdVj8JPGO0tBaS8A+rr5bwPlip0jl4RRt2
ZOC21cZ6EJmh3tIJWjrtoY/c+fzl2otR43tJrKpbzz7KZfuIsRayFrafuU5MDnQt
WSevljwtvhwIqb1o9qwHR6wu1D7uyQdtInhJRrm3VuR4euCcj+7aeTrnqTlkpgWx
rA4MZn7upcwJJ0KuoE7/OSDI0IJpal91a3Z1vx+xSEv5XgFOrSH0pM1HafFzrL1r
c3LA6ojav1k/bs1zSxMGRNXazwqOrJRjiBL2qCDB2JE8y0aCy8gkGdPbpPYf/Pl3
Hd/tfimBCgDpUFBRqrg56cAe6Bid8qmTY9HpHYk2F2cUPiBKphVE0PXTeVStYPh9
LXkVKaGJsFd1Lhs27hBYevNhW4lVAmotTfD2jMPne+QFhz53KZmrQQnSf0SxhfDa
nReKe0ZrX2dsXOWwDJm/WItfqUY7zhRCqqiZGV50MDoEfpsCOJNb75qFyd2VvQqI
zY+hgupouerx5OdJ8Dvt6JpdFxlxrrLpmfr/BiteRpSxl8z1iaiNMl8r5CuiIUfe
6Mbh8o365g7sYiuXv6U95PaG1HW7mF5bz2f1WQ3chcP6rQ87BKppsGZy0XF+i5TI
m3axP8ErWV/4F72r9TtUPk+3Ki8xF3M2do4Ze3Fraosf8wV88fUXBtYxcoPLOe6H
7P0rVNyTFH35RKqXatTnrheEEZD8g8+mfqLzUDoH/KGMCe5oRWVYSdAS6z9NZnTx
ma/R28HkmVzsG6SXFGNt7CGrP7nuLD1CAC6+HhYaZdl8wOx2FrGDLJlUpnduYrnH
yea7CWWHTt3+ix1AXV0bZR+DCZvjdicO0KAMH16dvYuvUP+X0rybGvJ/MFIFDWFQ
aqozhnw3MzSWyNQ3156kdZ1cyosXPXJxsl02mj3QtfIi6jAAhF8EgtsXVUuUnknp
InmoKxANUlRCyOBRkqyzuD3a2v8HP0Nz2B2xegBMFHKKWg2vupcWU4KEek5KX9Sk
mxjoklc4mLh83mIXkG0OZDRZNqxJI+3nPw6bsBvKN9AibsO4Lls9rDwSaRyossnK
qFXvyV6qdBBi/8eiTALhV5/7ml/nuy/nvjGcxIzU9pI7rV6ybKanpMbsiILea7Td
ig03/pgJoYEKdorQjIbAiUt2CRRBEY9HLqj/BemMNV59ziTfHYXgvMYfCyPO7RvO
2j+NyDo2ZFEdfe95PsJ7CVwhZ/SteKA7QaU1HDur25v/pdPZWH/mH+w/OaXGvbEG
/5Hbk1Vx9nQihkPo0Ovs4ejneEG7RuMwyFNNvG1LdMIiz2fVCPnTvHaaTV84UkA3
z2FpjYh2MZLi5sXHUzbOUcpK7nFM733A/jSpV2XiuF7tzVETeQI912fiklhrHkjs
+S6SmoxiGkYyGYqyLXkLZrfli0ZL1P+uY+FFqJuerg6SDrve48p+ZWMms2VbSC12
je5S18ZQQVSXXuzsDBx/VIe/z/1MNqKJJ0FbYQCZtVHJ/YgVC7zwcLOeaPyFZm4H
cb5ZzbkbiZr9JAwXlA8rTQ1JlxYs85GINRLmi7JsRiSo7TW3G3kBzQJCtA2M94ym
xT4x9Re2SIetg/I+k3KofAfSUWXUjUEYpUb/x/bhRndY6OtdxVSlLCPU1gODVerh
JjTO9AmNM+Aehu8FXnDLfHUBS3XwjeM4UzGB3FFqSaJ1DgkzXq1QTzxmkG5AhnQs
769hjcsqxNoummdIGPAM1Juamstpxsze/zorzU81VPpzaLuiaECGjFl7N9Akep51
Y4dJGpTqFzTCMtDOipqLhDKXQj8FStDC2Oc4//Dx7Zhj5oRogpW3aX8PdXzstCDs
LKdGomk3BhkuxkFIJrRvEl8+cC2Ep2ULkvX7pNwequWegjEVyRpiPLFXEKRxVVur
/a0Ne/td/jfL/nGKg8BZyYaC7tr+tYKmG4bJs3YDmAq4v8G4q5P5roE/dGACzT9y
kcuogpfPg9v2rsu68b6rvkbFYcicpJawtVWNhTBF7Sms2Ux6m7bjniDxp5cIqLo6
LOgWXWWL8c+qdhRnDhWvkscb+e28deJqLGgUJhXNEOGNdZ533zkGbieaLhXQWwEX
5a7sc8HfGKZ+VwGTqEEkympUCRmB3Dp7bz3plzSiagMKZGqL/gdIUr0A6+ajdfHj
lUbKZU1IGPjpCiYeL6N17fTAdMeH0PrCkubaZSvHZF6LGHigL4Yoq9icx1fFrLtf
VOa9wb9szhVoSkbESQ1kFT6IQtFsfSUsTBvIYAVdG6qrdV9Z7suOUEXcnd9nEcmr
hzAQcRcgA/7tlAeYL4MSGgz4TnSpCvaPL9HiWO22KU9N0jxP3zULvKpqsfTpwKJC
kIfNxwcnARJne+RI9ib2u0iulLTlCJHgZTp87sXvu1aQfi5dFrrDguwv9fde8f+n
HXJ/+HoGEg+aZhJjvPeK6zv3q1rS6LyMydSmnGgqs8no7D6qJPCKfHnGQh1DK1FZ
OAQ565KOAPXr3AKS1IIJVGBODD3drpiMpfPhmi1XfxtPujRjPlap6RYP8agLd6K6
ApAo+dYNAFYEsKfHJlcVRmqVqi3ci7BQOGVcprvTxQTXOvyqArtFdSw/mOoWYkjh
mpQ3vLC7U/Y+z5jPC6/uXEQ5PptlfbTrI6XiLT+Nyla0Eo6HNjT6V2fcAA7U5jkC
+NnCGWrArkkT/tnRnk9/3ujnuJT+5IcSP0dVqWUsRxfxeLBIhFRpVs5agEMalbRs
vVaMbYVHn81k47AXNR+lJfPBl6DUzizlmFH4UI1YT8zlIp9gt3bRdqxQbMJDH0RJ
volrxzxYx0PXOI3R/KhEGPDWiGX/ajSm8tm5s80VFj/lOZpXXUHpHyA8YD0lmV6h
SWHHeiNcyMNc+cJT2xmy0YLb5Y4cJ5MB6Qfdyt8Gst4wMQwRpKSkzINqmJIwfU6/
pIffq0/ElJf4EhtYvLClqFpqkrIZ6sWnXmh+AFmNHX6sd0Q+nXxbYs8/rGrt/K4g
NecP4m8xuLbRpBPDhh5VY4keYeQ5z/tA4wP2lZ5H4lndnJkIpO9UxXWjrxPv5+p7
fDnc1hOJDhsJh7l/zNsTq5/mI9m4V0e42XxJczZlDflnO6CVg386zHH81+HnalmD
vTNVFMa1LFoAcTicG7VVBWSsJfOJ2v5tV7BTntcQ0VjqA96myKv3dlb8++fcFsYp
TxT+iL6PYOpusIIL5CuElNCjogi/plNhVRPfm4IJHrq2abxtdZF+u//q6jtGq2yG
fnjnxoRWJYzvOQc6KLKvlkvMlnn+YzyepAyQgGKMBQbiQAgwAQ9EzYQvrLjWLL5T
ChQrt+pg5LSHA2GsS+nlk/SWdTl/DrPXvPsMzZFP/0pZGHroKml8y2q2LkxlmYnJ
PeZFoloj9JlCZKa2nkpDOPoQ1sZ7Sey12/Vom0ugV67fJJpaGiUfY8gdVs32vquv
W3/Mcz28wZXFxeepu48X9PI0pNVnrYc58v0HLq/hebl+KDz1aSZ2yk+ew9IaNjXG
HC0FfYs3jovjZwZ8cr93L56LbktZatT4RQkE0tD4LROZWA2A5Hifb3u5yWDi8Vva
WmezLwncJcUZKaLyggSUOG9hd1gc07bKpzhC7Isfn95wapBfBtWGKPFu0AECpawi
85+jqFynr3neqMQic6WdoDX884hW7ZmYnHKnvhAwHBj2JQD0eMKasu4tPMo2jySm
KgSLOTZaIhupBTIn1Rd8El3FNFKaBufvOWbcyCCHkOfGXYbYdTK9Z2RTH9zflBj4
WO98WEhue43qxigYzXPwT1SkkYbX+L4k7z+yWUj5P6+TQ6zzQkNb4OBRkuD+ESYb
/xOVYk0UFL+QuCrYYrZKXezML6BY3xWze+psBxsVEdeF0kltsP26GmBTmJYx29Ji
Rdy4MbWhyT+eaz0hcacUQzZ6tupaKZfqHQEh5YQb8xfFT3O+ApUzX2346a31robm
d3TncbPaFxw7EF9kHPdezPxJasMkmJZsx0nPqPtzBuf07WlvNda/VSaLXN+vtERy
I3JxHJ+Kvvs7cS86o3/fFWy46eX2oFkPIpJkepUh8CqAHJTYwq546d5pIcBsgnI/
jWSECALSa6T1prjeES3Y3w//QyUHwj/JvhCF/zjSED7jEr61kYKN/WAV6iTgz0j4
aKuIn1tsm88Bgf8N1s7Piz00bTUQXwrYSFfctJ7sYbMvpMvJ31aGjI6B/bA4FwYt
v9yQMSkWYGtNzfNkVV/NxDMD4vQ6QxCsTFT3QeSY2Dl0Oy5SXSij5bMo0apHVYXy
zAYLAZIMe6SwyCN+eL3rNFo4szgdmctPjlsAozmMaYSOnAsb6k8Hgd6PJoa15FnA
zrhOaZUxbNCMVGKqzaiTJzPruIL3bwvGzlphOeyzXO9Ktm0ldxhPYZBo5tO7HEE9
bLjN/WU8VCUk/So6GMWizFmv71ORyChcK8a2AjKunXNvnDsLwRmh0L6QYd59BegB
0nWfI3k9vqg2gWbSIr2YMs1+wD3zAYFD2LfoRopGi2Zxatz8X5aF0fXusnc43mPE
eS74VnpokFFf1T/i4IVks/zH+A9mIPmeoEOUVOR2fyQ0qzfr562qeR288NB1H+ub
7AK7P9GE3al6ewzNHEsDYarUEMpp1D3IXZAjbCA5ewanNlh43TDvkgFAQK7wGoBZ
gie5YQRUKS6ycRAg00lNks+RokNR+ewTMVTBWogWLmX8Sm68ml6W+BTMC1WTWHO0
BxAg230Oqigh/0Yc+3gxd2uRrNqL/ZUil74khJ5jyruxzPqnFsYMSujp6aq1n4Zs
voUih30v5ojFKt5Fy6L0uM/RrKd75+NDi2U8y+krYN3iAgDtA1XDyyAOhvwm5ng9
NIurtiwbZYFgDjQswIKz80tKElwyXy6waFZ99xbKBbopuxpPAsZb24lqRNRxBc7f
xEJs1XqmHaKS/g2rYgn4P2glReXnJuak/95RrbYEZYbusx019IiskAGvPGcnl6gF
iyIRhCZi+GLY1TK5pdbBX6dc38xhs9HNxCqGEkyInJsSFW/AuHlt9r+Ul90sBBx6
YVH8ebX14REa42vBNbLFQzSlCts4TUkgKp/8hIT3lgkHxit8OWYoxrZZBswoadsj
fexEfFbVEjCcJDfdnSnTns+PqKFwKO7RvXAVZxOQ8P6PlQE0ikqwBx3Hz/c5/Wgx
L8xvabeZvvF1YEHfsQaKLYWjS+Ks4PokEMA+cXh5pToB56Eem5JTlZBuhp78/weP
bRs/8Nq333JPJx2trkGlw4wpVPrrAySzEUpru4XL4gsb/BUybGaRfffoUNU4Y69W
mbuFcuytHMEWk4FGwuH6sPRwiZ6AEKrAdcDW8sJp6h03nHqp9+74+KlxzvUBoWOO
tbyGYf0EYXpT0M/NZQzkOp4VpnIk7ziZ2d6uAyOYhOZDo4EO6gVhzhqVOPTaPIE+
4nBEA2/PHcTfDrCLp5sFbn2GelhlnDPTsXRxjhTfd2nqHlp7SACw8xGLOE/rbMul
BcpBW0zHYwYkVEDo/6WalqrN0qi+POKbncFN4WHBJEV8IQndh/2T2iGIF3LE+Yld
i76sP0OgvJENce9TXiVj6fl5DKr+W1Un05MTYt8KPdcA1Fu1w/+hL4WBwtKCiab0
6m7dYxZ7eQeO2onNOGRwsykOIXIASVDBSzlU8sK9KVEDnHuC8Bo/CGmBdJ4GGNBI
aMQrdeI1sdr7xuLbsU/PuaFg+z6UHtwrGbgDWZXZ/NECiLto3pnLeaIxaTAXtRWy
6waPVUm2lN+E0YJ+oggYD3fTCQWn9h7xCzg1Yph52M2XwqTGVHk1wY/ffFKqQ4f4
ybTsc/JB2i4eHrPpFb5AFgt6I9r713/kGyXFS8TfV0eMMWOKIA7Kpfc6Mmp/b2eR
8ifxgSF//uR1+Xzg6UHNUVmiYOD/9PgIp76dV1Q18jJ63jqer+giBKHp08uTJ+hl
woKS+0a5BXcKwv4LnOd6fGbyZCh1aZ4MquzAbyPuAeb0PK1IuoOvyoLl81AHZHBo
xlwEkfg+23zfMptUI3kPK5CirAyvOVXPtMRXbIaJYUjhHUnWUUYmyEDjtTTF1uFN
HQw9OoFJX66O/rLAVfwyh3Nmyw/LaZE3hFAryfrgx4cvudzpIyh/EGqM1ym/wusr
7T8e7+PwIcKNVZLhDIFXd5mhws6v5gd5KYFaDuvUSa+DQvf7GWTGk7LVPf2TJUm5
0/VlvXHBMmAtBgZjy20g45eGXkazquloQoV4u1ajF5c4ex7MUYHU9rkvt52RM7Az
9gDDsVt0UaXpaLoXsawMBtLTZoxZ1PUap1vrntdBykBPoXyBBwKccHdU6ZmoXNH8
3YXa5TYmyR+TuFBQxJa1m3p8Yp6VzQYaH7rsD6PnD9JDoBFANiDcRjKVGCloULN3
C7DwJYYMUYCchdnhcPO0Y27NPH+BUayj03IUyyTsV6e6P5bjQZS/JxendUKDrHO+
YfKWG7RGy9JRkVr61BCpB1y9Hj+eZhx5197W4+Z4Je4J2FPpgoF6IhFxXpmL6jNn
xaqY/ul9F2DzS5QOQak8fCSTJlkulrnJaYL1KwWVUAOvmoEwVACSt/sQt/afM5Vq
HmQAMpCXprESACtuU1RCcydz6K+YYJReLMdGvRW1DYNu/vm6sM7TA0eVk+o3RThI
eCeHqLN+QVezO6OwISrQUdkUAb1f6vfgGh3EQRQcESwNJi9KGogMnS13ZCQa5gJT
4LTVmjiWwMBwoaZ1ggqgYrJdWQNt02UarXk2dqP+u8E7I66QW8JzeNYuKiiSDwL+
bOL9sQ5qruPmDpInNqPliF29BDHfWQyxDVTZnD8Ip3kU3SSfu6pWFuThDuPnfXou
oSMeaG29+MQw+43Apbim2naGjCnrxbj0+yLvr2a+/gusA7giKC0X7U9JzU3LTf9p
xDq6+Q7gN45aAbcvOFsETziIdwExb8fEfHmvKMCaNX5yPcEbXy6+vERopbISgZ/6
uCpWPadxe7JUslViAza9D6EAJ/D277ftgQn5XtKI04TfqI9Z9bpMAZTjZGD8xHxH
SAROm7QrK4wDGVMh3CxCxXCZx/RDIhMvncXxI2549HBxd/pzTS2aZiXavm7bGUN4
nVKgx/o/SQGHJ5FmwQTwsCutIAtt9Ht1In6Ue6guTXFcPUT5eycVnQFl5zwxrg+o
e6mJSFowpB8q0o/PHiVkQye3//chzIiDq+uTDPHtmFZRK2zfUW8rLkbLrMGPkIOi
p5D0Gk4lKM1I/rP01gH5/JcozdVhZdmZYKU1yRYXtRSuByriWipx1MZ5a8TXsf7x
1Apr+1YswdTprGoamGx5SgB4uvDmSbg5QPGq5kjv1b1cRBU+i4Qy0Yh+jBzmRfz8
a44iL4WTlQ+9TnkLXN9j7F1DbGBsOhwmYstc2GARU1OHIFbCIdo7qlYWyDipVlqd
3JaOhmM9VJjZsLV8ogVgU2iV0mFwWLOgXZ/z7UdTvp+AXUkhv8ag17ESdazq2SIO
J7qM4wt1m6YtPff1nzuNuiwfUUBajji4IqPfGzTpuAgSoULRB7votVHCHDxIsR5H
tdbdJq9ziRU0sbry7SENGif55vUbKbrPNYR0VuxLnv+rAma9l8HamAfiOBz8mQLu
EzPV/Tk9IJWaLxx5MlTxGd77Bz02qn1vvykoXrixEG6E0OyXshKCHR5hYPn+qLeA
kYFGGaIFPM8n1uGGr+onboVH1zIVfCXvqnLzaHEGZkQoHVrK7FLZIo1+/IcTa7VR
hjwCzyFeM2vwJUv+baSJtru492c4LQ5Vl7VTo3mUk2RoABaWuGCdgCfX/MsT76jq
4ocyh2/j/dLNHLOISC6Yi+BMUSLzO19nLVOf1zKoFMPpodkNRdcv4JAA/fPyjFSo
2hBi1sRj44HbXfPlpl1OyTAbFntKEFRA6V/WMFhJxJ+OMU6LEZ1kI/O9OLtcotYJ
NF6qeDQi993c9FlU76INURh/OutS7BNK6bD9TaIYGD53fTaahCIAT2aazNgDaiSV
X5iHvJPOPkCgDr+4ltQ8+jCiz5DniyvA3hSw7/Ia+0P+WMdWyVgXvU0aoYKBYt0h
b3QVyekXinuNuTNEjXa/8NE5OO101PosbiQNCTtaa/8Odvj3z3bi3jcIvErHmXhG
MPNtbGN6R0oW2WohgS7zez2McGsKJK+xgMmkJcTr+5VvDwUbScU5Rnbf3Pd19Qxq
IXL1T8UzvRr82J5iyQHiI40G87wiXYDOxnrzTW+aGH6OIB7lBHjBjGjRTsYn/XGB
QTvux0Tr5aFbfNzAFZiizNGwZgaWKLcS+GToKeuneuMfhLAEqyrDIhpbc1acGleA
IG16qpeFIimdzK3zhrBBaVGcVdaHrZszKw8DUs4Si2YWTGFk6Z5Hpc8XiXSaqx2E
2op9U/4oFD4QG5/jO2B6j1t0xk6WM48UmgEB7Rtv2T6tNKHM0BpZeh0sFaGkRSM9
yneF0b5lC31qPuc4QfZqLXw4B8f8VdM3ZtGvI2JD3ENOLc1GfhRZ6SF9zHrxBxLI
dWFZyw6+ODtmaCnYtKbKbGx5Cix4eD6ZoFYT5T7nH2sQZXPphiro2qp/UkDOOkga
6F8oiq8UBUSaM1TIWxZg1Ny+3QWxAX32C9snQ++6Dbr/mU+RHTqjigCnH8pICTad
+AeLNcqdePMwbWMeifInZ97YgRiYbf987H0b9ynBSzRrvpT6s6DidYKrO6IgaNR5
oAvIDhcorAHPOYRv1FHD7JsNC9LlVVLY/6k/VRm1X3DCYM8eW0oy1UTiFJMmZQUP
e8xtbW2jyOSyNENSOJDiDk0UuQZWWY8RgxjlgXU1l9Bbaekpl/l5nUcg1uvM8sDA
X1nHImjnuNaARoQRtU77JbAQZz+BzLQzpGTZ6Y9WZsERCIUbJd2e8m+mJY1/irDN
xaa/jXQiptDxfy2H8Ewmr0CJwRvz6Bz0Tf8vR9ppfiCtizPFZrjQvAXLrKcKB0nQ
FvnqsEAhFlB3ILyb+KLDNRLRAP9TJUZ+7ZuVtBxyxNeR7dyQCeYilO4oTknUee/d
oQO2Aj2GVEaqlWbCxVcgCpx0N4uBV4rkc+SfE4BtgHvhCWFPvtgRkOd2ULKtJzr5
ZVUdLdvRWXBeoPSmYZS3ttRMVfgfXAZ2t7OHYqgRO5o8Ia4Ss+7edoGsNW7RAn+9
+PZUpolwFD1Huf5bjOLb/HqmqcMJ6GpXKVhE7W5TYlYMV+5A6Zt6/xHURzJNTKVC
lvSIE7RP057ih9GeoxxRho4zk1bD6MMum+8G/hdecbhTlDHy4lsIRraE2eF6ASuv
kpl6ezNMZgQ6DFQ2m+fkFohGj5/S7hspEGP8r4Qehz6h6xsX89xz8jEBHGAa3xmt
xtH0CL5dO0JDs/R7NIPCR8N9LLRcwCkgNq4HFdFpgu4rLr0qxYPmY9RvkZ1huHWg
2xNR497ZCfq+bd7730RlZsTfbk08NbuCO+qwwepWsHDGODKqkLFPt39LNR14GH+t
ZfzJonUIP2SNiFAa5qbGwZQ+ARiAGwnIiyCQDD8/Ad/uB9svLkrPzJ4Bxw8QAyHx
l+VQPO3b/GUWFc942EQwgDnjIWYWOOFZGeHxW8Qad5+DdfsbYGkBZ7liwXcYQwEU
LBYQosDy1MOpyQifU/+nymL8qoqbmpXYtQ7eT4RzQH9MqvI5HelEpDgIgMYXwjdu
+7EsjfNe72YkI9jxl2PLOBiX/WPnuPv947f/mEV1BOENdU3fD8ymZ1dLFMJCtHNU
PzJ1hmbtqaKkhw+LmWdMCM4yK4wevo8PpUSmECVszoOvrnYFNiTRevPXQKyjgzkC
afWxriFLRxH5hEOt6eclHi3UIQwl+hsmkGKgp2yJwlH4euHGEXKtF1IsUb9E5dhf
THJQh5s9Uq1xQIh7eDSyWD+CRLWMd6/r9hyhUBqq4t0oxtarRvI0In36Xujej9kT
0PfNNljDmnw6onQjoRdoq7DIpIB7vl06pNuibuLDaDCTSrz807k0yCFcJ89WwuKb
7IvuTR780NYo7UaplKqQTLxqmcBFgI0M/ulQvZzCmMiKCx9xvN0WuJhSghJYLGo8
YCZ/LLsQ0Wto6UTJk+U1xzdgQPxlM6eJWGU4ApGCVWtUY8i41VmnNGYaWjDLGH0j
3qK3fCdwsmUKvz3Ibq4Re/BLv3YA2+4dLyL1UrvlNa2TpsI5YTCdiEyPWHKMG8r2
Enleya0waX/Qn2w7W4payCXDrVqgwF4FAK9o5bJv0Jsgq6Kio9Rip5/T16Fu8LKH
7vOAcb4NjSxtXxpElCNkTh8L81WiiD02/qTxGxTnd2wfewGL2/9a1Qxdu+JkxwZp
oo8PaEM8vhSHS/d5wdEDLuFHh2eOFtvXhIrMPBGphFiVQoZZuw7sdJaRgP0qp9OP
iU5v2w4LiRBKbwXkLeIoHF0hYcdyjULTItMLeiUEyZR1uevpdWEYsXpGtSpwcySL
kyMYJocvfmiTRpLN0Neew0c0S2jnfqDX6uDz9VCl8evuFpL7SV51h3824HsZPoZN
VPbU8xuOuAUGLlTlnsAvmE5rDZAAPm/t9IX1eNDlqzTl0ib0jAaJmU3C8oGaxP5c
O7e5TpzEqGtbdrj/wA1CA8eZdqTLbsmH6wWv4Ny5/apPcJkpuBDNzr6BMdV49AEM
KVVel++nIxCZx8bSrI+oayyCP/jABxre7hunIbf2wKr0sme7dDjJKuHXEqnwxKBk
8DIyWkK42jyDm0zkGEs4tY/F56ejo+kDc0nOK/4a12fBo8DYMiVubIULOBusuGbR
qeoEznBhzbXI2ybzcRnjlj+zsXisDEAeJz6fpQYnQ/HxxBc5oC4Ct/fNIhoeOKVD
/esoBpSZW3FMgR1iH3j9EE4O0q5lzdb7/G4Vg8Gok7S1gr5yqM+0QL2uzk80jJSs
P22R7zFClvDfqtqvSCwzSru30/Q4JoHg+nMIHVluPCrKlD0cIoE/7/ibPUgFyU8u
vnTKOiYSOx7bnrly2R0sMltM8TTTJES8p6POfDy+TpcxiEUlWrfZ+MnkrfyjDYN2
35sUiBeQJk9dOTzAU8NnvwXsrySXBonIcu7T5Y7hcfDAAmV1Um9kJ+jCUA6q1o3V
MbPwSmoWnX8XfelhKkyugwNDML4VFXtwTvbbqAzHbcbULmCPFMjIykphg9VlomTV
eID8+ByNvgrwAZlJ9R5GjntfOv1OEFbnIEKCy8u2oCq8UQCpWTIVc4KvBfH/V83N
73Qt5WpqDcmpGGcgaIZ6Ww0rvh8MuwcWHnPeWHmUhUZ1itUKgpHCmtpq7dH5p+E4
fP9KntI28qiF5cR2CR3W3zJjeCDAN58aiGpsTxoN1tuY2h7+GF1Ueeque8HauUOU
+HbnPLlIkc0Cm9XyMHq9Z2dbXXBbmACJTtZkuA1sOcDCxAq6p/zOLkwPBNi2+8KO
azCBhdKlzTtqE2xtCpgFqYFL3fzQGPcrzx0YY8qSGFKrs2uFzUyMzN4GcjuDpsSN
r3hYMceLq0JtuZOd3sMC1QFDMe1ZK5MUEbFsObgK2i3hS5A8LOqyYbueFj6T0jo0
mHtMJAOlD5TbcD6FdwJpGtJxRZOGPuPcIAYAmb4ehjkKKeZndACZRjEKkcIVmQzu
uttfMbwNeWbR+20zFAfHhRotNao6JeQaEVTRl7s7i3GtxBy2uWr8FrNKry1WpINS
6ivXQ3yj+7Vm+kkpuXfK52pmVevC3xXrWeIV9pnbs3rg8c7lOG0nfSn1gEtaiWss
Hx/Y0y2PxVdka16Q+FwjEcX9TyNEl20beYdUaP4IxikYSFm1WjdLqT4cBJ6Ks7HZ
C91qyBZHKaO4FtnoLUpV94RZo6pq/5WZYBmzDerzYXckmFfhJYTnbYrCnNtJIrUR
IeTCvcpWfUNpBl0jbGk2D7SLJwWA1NwLLhSRHGBbbNf8mRNLzQwYRUV29801gz0H
oewo+gUGo28oSOJwbSecuMLSz5DsGYzVwdQkFONDV1ay7P+g4ln2+IWydA+jiGhl
so/ADLTDVuIA3kPLm0xFdpv//CK5sDI3AceKVA82h/Q/of3Fxufgxbg1yXNE6i7Y
ftK8ALSMt6qieW8GNC1lz70dpdr0Rw901DusFfh55uo4H3cYWTOnv8I6zPG3BB5i
KDpfG3BtSkAjyGn+D3xDn67LuEOXNPGeKExUW1DxcXXbSd5jdcIeDT3fNdn6pO55
mQtnu/Cuzj0ZwSD7k8E/9U5DLBbwrh9bCFzGK19R4crAuQRKpSzNThoHvQcbJydB
AiV+zJaV11bTjrUil1fFA4dDCpP2o4woygsU0dGzgjC+VKlNIKgyfqkdBedWNMBf
VISfBOrmz/2PjBVrrFs0GnlWe1+/X++Rz8+zJIC/G9lMMaWT3UwrdWJrrgZTF90U
dnXcKzkWkDYDWbBMApcF45TTc6RBOq7i5384JDfFaZelnH44tNi8Wgmmip8kr1OI
6nVdmU0VtnfIE5dX49LvSaxTOwMIhwTpoluLSQOegDgEQvZuT93NhyDEJfBYwgZP
hb/FbQ/8mrNcYwf/JzINmCy/OPSt50avnC37C5AIFT9TUjCNvBTBLVrbthhqT14+
0k2mwpuVEWhG9prLcmFjRGfTjiXA7o1RNH0SzNs+lVzRA7s2QnzszDgcz7giJuME
BnW+jth8jqrfnU7ghGZV3wKB+3HMRnkEOkZo3qU9f3wq3lcStWxwylBf0ttnbCv2
W4SdeKBsodVo6JC1V8m6g0LiMbTyyEZ3XvZrmu6iu3IbBKTrOiavAaIiZYPZIwMv
EwA0RBx4xWPcUF0ux4RD4hmK1ASKVAzqFA2ee8Xmg2ELZ3vJ63ZO9BQy0btwZ8tH
3Lh14GHo22KxscSmL9BdGRK3EnRvxtJIiGbAx7Z6lU0x7ZDpOH0b0yb6uUQLzvde
vSJE1CWizrfSpIqxmmfwFFYdxgn/zIiJWN4oWalKDsVKf3U3biZaAVk46ot+iu/i
cCrXNND2SPjdtrjFcsQ3toOqmcqw7NlafCZGufdzwP9YFHxV4gx4p3tz6mwdWf9g
c0xoaN/pGyBLoYmYnqxwqGP5xizfu3nl+J0O7GYAcPiyrjWANOm0fo5cJV9J8Sol
aoE12T4M00GghxHRpLGQuZZNKWYW3bV+ujczG+BhCAS2lZ8cvSyBoUNcBNJUgq2Q
25ZybymlzLzJDMmiZ6sr2h5s0hYTUNCs2W6BWqZsH364fsUMx3NyhmMJHR0v7mfa
/bstLlJ7hoh3YUARvcj23Kp237bfrz+fc2DgNz7ZGcCUgyZ590mn1ELyPD/aPRhY
GbFIuWVGuH8bd7A1Xk3LLdIGIUd+2i1usDtWfj0uax1sBfv0W/+hbPECesCJhIDe
gRAN8Kik8CggjmtAQMEM4Ea28RWbPsFEWFLnFqHWu0yPhpY2f4wbHqDRWlb3VfyQ
c1YdlMmNO4jhwRmzwd4xamBnQkDRPq3SfVJk5dhPH7gu+FfE9sIliv95NSEIq/Ut
qbpxzkHR+o31vax90ZK/NBo923ewzh/9aBCnt4HZJsTj7vXKpfwJAgwvkSdPQroR
PkrvqbRQ0GCX7vWubF6F2+3gF++jiju67AuA4JLyIOVJX3rjaNY3pQSzX1OobA/B
QmZT1rr+N7uqNDUXL+DlLswSuhwmmv5GseGO/8430EBgDKhUsGBJufiEEYH7KLzN
zYLC22lgT3LeMZi8sbHfQI8Oyx/10qOrIcSAIBSJ7BQJzNweFAct+Cwc1cCp2bA7
gRcahVP9mHUwMs/xocYhfmiyzmvzA4mb/uSV4u8zL3F+hmeGQrQZQd7Dx9P8Nwg/
uRl4BcbqLkqg+vHyYQeTEovy0pX8bzLjVd37WNkN3vSYpCiCbOYaITRjKa1Tj8/6
kElTY8J/mEJ2jSQA/a1y0+qBzaqalOMzm/U6UYLuRiUsymT6tUW2MXrYKDrJodfE
AuiBXy1ayxlr4W1ahgiheUED8zEam436v9xDY8wGVhbitmAm5F0LVBQfypO9nLJ0
nUk7NUIU3EXgteLpUP6WVCQYYofg5XE6IRAzNrPSRDJ98U+B8TvTWSF/4jhbmxrK
gGylHywj4xfDntJk4hdjyF3LSAhJCcd82AUkduJUXpxLOfJI/W3De/kTJjG7PbYs
0o9J19Jxv3WoKQ9/aMt4op5JFDasGKi8/IhymEV9ET4fdJ6YyoMGk/OWR5CevG4U
ZCluOVXI8e0SlmuUpglr0bTW93u7KyEeLdNUc8xrQIYCvrwEBLXwe2igPLdruL8P
DWIf6Uu9HLLxTKYidrb1UZiyh/xJUW03wDwpfbnYTL/o9/pVMn3mfItNorIGcrHC
m/02PoRlEy6aBQpDjKeNM3U3HAFic6vSraDJt44/JofBgMGKNF6b8z69jNPssRK3
06DUhUzKHMMLh8G+Q8kJCLV/8Dm7Th9QrdoFOXruTWvEwYZYy6TKgp2JFG2z7UPN
Oi4Lim1mGiZFPpQIVpzIE8i6oKsacXrWRl99dxKkmj8fPGdxwKGdsTFAuE/8ffuh
YBnbvsDbBBJIJIZ/6ouvcLpRMo8sTMloKRmo5bYhyNK5G90zQa/eCkoOaRftjXEF
72nidQZnq0PyRq7fQHpgI0Nbze2Wj0W7ycGjt0ZoWAOasKMzFIYEfiO9WeqUMF8x
n5xUsiwiKFqYrD/PjNOjEylHtN2SDN5SDMQS0y7j8NoM1utGMUGASjy6HMOwA672
WY1cvdKem6zrIGXhcjjv6rfMG39uuGAkVRydv9CvzBJh/hBCZ7mm4JDJ07BEaOgv
Y/n8abucw1JW2gSGU5kVUhZ+G4EczuzvpPlX7zIngqeWeMybT/a81rFsiZXb1Ws9
y6CkQwOi8EioCmlNoPvCg9Nuz4lbM09TIeqZeQVWB6wg15Gd/3YYcSYfsRCZPAA9
mPskcjdsp1XQIJ0ZfvjxAlRiQkR43PrrLPTK1+fuTlP/Aos0ZgvPvzoc04E+0Unl
NsXq9N6Iy2UMJAG9TZ3x4eicDjy4e+kUVMDKghaekkHkf5i9pTx8MTV6gV7kbhsc
yYhPftK7Ko9U6HKcwE4LsNkwH401xzq09HkS+tFUHTFh0ZqbZnzpPV0Mm52HHe5k
WgC24NXvkX1uFZxryNKtnePb3ZICE3xxqdd55Z6Mj5E1dcIrODGhoNXeJvRizw6D
IyUZG+uSdetcvFVC5xrCaxqUe5HwLq3DPZGp00bX+gCh62g+wlAZnE4CO4xd3wnv
drl44nfo2tYzZ9JSDS6O34bhCeGgBiw8qCk+AUc9eLjuNIMWEewYzgd51BEM05wF
zvBHRsvG33MTOv3XnHoKcaFAwAK5HeQzet36njekDQvDua6TityJ7R4uTdOohbX1
rCCvX56wXzVmqCBrCGtvPDtclgpMYYdVX8Ufot3lqfDU9nGupASt7Uhvd1F25pX/
ObEVQ29aiVRYIREPVggpH1nMo4sP8rJUXCUFw6SLEtuLn8KD1P5lFO7CZ4+qbOmM
LG+Wp3GBLkFJKq2r9WsrlRWthArrUL4C5ulqPgfv9jMJjsMwT5mUJJBGwMNqRKrV
edvnfmr+TexI71+TVbhd7YuCP7jXDvogghKkdyv3U4yLO1r/9HFjclN92LPhtNgi
aWnTgtzAjD2J3Ef280tpBty6aNRoBx5N/WHKdotrBJX42hzPzLwtN32+vmvVlAtU
0LQBtDtw5r0Os7v+XYHmvBookLJ7KArQzK3NZuG+fVEZI7nzQHaHRjlw+UzUF9A1
HhOqDEUEOVnFIgbpFYeLqCuzv1Kzd2zzpV20+kWxv35JCA1HkQky8XXHMO/c6dBa
rhwyDtGRp/dTxTcPBy9/JZOQdqz89JjM0ocK1rO37sA9uXl+uRhbqYWMa5rETONN
tkPFCD+eqeDBgWcoTLclxWZiphfjA4jnewJbcWY7bPy0ZWoqowfNJ8tmdgbo31dj
ECJ7hhD4aEI7fGmfwMqAgFbUYjj2LpTQeoTC34Ha7FBBj7aWd8YR2kQH7uwRiHeF
xUS1syKRwdpWAIn6fGBCOje85vnO7iDa9VzolF1W7Clf0re7aGVw7YKRQZlYB+6M
RiIa9fxq2Va0xQ8c3N1/YdVtGKpooaKyWU+qNcIp4Qc6lKXDHnUAzojfPRWhdtxj
/tNcp3KnQSipWsXKrkhDb/aKFh6LQtyzFULyJxYjTwKPWLc5VqSg4EFbo//D+6y7
G/HBI/P3+VDbbbFXKI9Y7BE81Hh/xv7TD+ESX+wHAawAYgPQTSWRTWh9wy9BF+Hm
pvHfqFtti9regGI9R3oDd8IlnfguESatTEsZfbb1riuLSDGaCPuSFrr7P5u89f10
4cIqDB3vEkTFF5kcvLoZyGs/EMIatHwZP4QDDGWzG1b6b4mQ7ZdYTeVANdzuvG5w
chS+244T6RhxxyJyzv3cs68HXN49XSUw/O0lhR9tsW0G/pH8k8gnHr+D564HGnJR
N5OoofQCFGzTNf+0cgHIKyt8DSAjL4KipiKluzsWgmVrwCHRe5e8CfjF0u2UBn8F
aLDpArLE7P/sBY+lwbfsVGX2SmTzRzVAHKbCWjnEFwIYDUAsiuMbOYhcfd31D99Z
o5U+wGpZjyUJJiGzYZTCW3xzgXVznnAyeGWLI589z5fshyf92yK/aMqZSlBLu3Vd
s2R3YhRdpOLd8yB7hRpVCm+4anXddcmyMURYTVjDEzV9SSX1Nv0fc3KTOop0FwMO
v+oigfHhtf0S1KarHK7WX4emr++592algyE5/qRvN0so0yVBF4F5oAAys0NT0qzU
pLnsczQZHtCDWlW/gng+nrqbf83WJtf+5jP7dnOoM7snhu6qGL0/8yOz5kwFsPM8
7SMWufNNCm9VpDhMpo4GsQFZ47lE17vJLM5RSOrMReuNpc0nWGtDMPV5IXIKED6a
Z7OmVaFhbmNERdcQM1icRGagxFQ+eADlbLYFxCtaKhTEJk4Dn+cHQYG1QHxhvwBL
aaCekdEQjW3vchp4C/UNGFAcxsjEK8MXPs0dxX0bTH7CjcFBe2rU3gRN36hvt97I
upzvBol/3+ZxMnRP0C/ZYOhfP4cryatrZGJSQOlkxJ35Y/jhfzJSc1+I4MVFcX22
ydtPGbuVb81rJxRwbCUYbWAFjQQHdoZIPLYDp7VzstJs47RZvWS3ii6SReDHEDIP
WwF4VC3Tz/A8/TEj30e6ZcMMUrg6WfNazkPov2wTPt3qQOBvVnSYI0YZQI4nzezc
YTVQeiKgzbQetLnf6unItiig0THMUT0Tn2KjAMGsmJOG4OaGx66Ld2udBfJ9cfWN
I8ivAMNbrDquv95NWDSJofsVUMbyjh+l00IkE6vCo1ZdJMq9FxSBiSKd5905B4mD
glStaWBYjBhqMO0A+KdlyBnHTfEF7N3QPH5nPz6t8IA8sRotuQV1Jj/8sKf+8u9N
cgbhomn6J2sPuRliTv2r/q4HWW293hFIu24VXe7La5rlT61sxgeqbf4S0kXwE89n
vlrns9KOUulnHCxVhEKMD2vVtgHJpt0E0IN/2VJ7qQWo9Y7gNxzIkauu29ZYHi3x
/HJOCC6iC6gh4/pThsalltT0riaXUjzArK5nwDBLcl9d02f+40AqdPn3Maw+3RhD
ow0ckJwcNif0Wy/WpAGCcQiE6ryu0Y++AF1ByGO5bxUMlw2wstl4CFNzX5zI0SHz
kd96zceW9CEsp0cdnCfPconAEXgsVE8Ae/V18oWobPxJNM/vK81muDQUlLnuYo9g
IR0ty6wztCMdPzFWtf2ZUmOhWlX8UCvk+bm29GAvtGqDLbJJHp3oQ44PhxEWAkCK
QfBJ2+OLK3TvDsO63yl+JTm5cEze7tHtzD07l3hoX9c51mNnGgojS6HHo/ZyQC9/
grf9qbNMYo597x1H/wen6NPCtBYKG7T7n7QMqU3nq2TSWY3Fhg4dY90g+ZGOqPy9
/hpbsFt+45yfOcuxK2nSGqJ63IYp7J4fDIIHsVtpUMEOsXi/vOmgZjmu2AU6Ic29
oOxKVQOE0jQBLOJomU4sUoJN3j7Ww/WmHqMDSvsSRYLA81YoluOYCrVa2QgKVenr
KxTtBZYFFhKENDI9q9aKI45+2pE1c8SWZBtB4RnRMfU45YSokUKLWPq4v7THnX3t
ua2Y/vqmn8R0RA/+sB9Dg7GazfULSGpTKSuBeHM4fp2OFPw5UE3fM3EmRNNsoXo6
iP7Or12vQyCDbvhD+QmNNnn673Ce9faKPvhaY+gNKXtipW3tur7cAFBKHTPZ7JlZ
/r/1osNF/sC4RccF4WOzl1GrfLL4S25EDlwbUQlFp5NpKnSIiA7z09VfxQO9F/Bs
ftraR/CICoIdM4gfdulCsxmxTXara+4jZV9cS6m1tmcpABGIf2BzRKEUESf8NAvJ
MBXx1RCLe/4dn+sKRZ+AAEj/Q4jXb+UtL5nn0QCkw2vN8l3ycyZmmpWx64SOPigz
JdHSgSIH7kd5zTw+MdtCYjy/Bh2ivIXB6ZQVeLvGzC7/cRyhr1emg3EjcF+9FxFY
sDRveTyRyCCz7kYaoUfXng+4Mc2MmuhhpffkFJFoGLK9Xc7cgCF5tAoo5RsN16j+
R2Pulq+QTRTX72PpzEUUxtDiBdpVAcAq1LCXDBE4xC1Jv5dWB/4iUlry8+doHL/D
ZZpB22oxC1Xr0kKJOSwoGsXrXnHP5F5B4cEf2BDwT80hnxe6VnKeHd+iAl2V4eq8
pRPxN3wCrmqO1LEpqLMy7UNrPyyJB3uiCSwgCvUy1w6hLqYuERuAfP2gO3w9Czf2
ZsMISaolLknWsp0iGeh5SgMfQ7hKXOGWyz4DaF7Q+3N31qyy5wvvnVHvNyzUO+an
+k5jyPtTHB4nMT0HMCN0ZY9ZamIVCNd+uMXxoGQXCDJLQANVZ+s5besklZ8YTGsU
wm+fzrszIsgDlAhX/78EFclErSI50/R0gak/C/I+IW0QRvTIPmz6rJk4NX813fK9
8LX7ZxfOP9WWLJc26T8KCNqvQW5pKZ4VyDxoEPAipnjF+Xm4h2PK12vKVIq8Ze0V
i78EIh5f97YT091nxbCrxDp4+NfOvLEYyycY55XKhxo/T8LvoL5JkI3gRuk520Be
F5+cTqzTU1sRBBwHj6+W0FI5Y9V73tBm2tOeeYZJ4ssvu7fu4qbJO2ga5PhFlhwm
Kk42mxkaT8sFlxXVE8x0a+xWTy9D5eKQjHDi+/YVxoZ/SkUKeMoYB6NTTCcYOwx1
zKPdEJclh10WlBpil7CDA8Ggxv5gvRWFvdt3Xccrcs8UmUtj6ni/sREEWgz1cCzZ
9ACNXqaz+/xGvJ9u/oIBQsOICF2wuh0xEugisTGWIm3Bcsbyto29Pq7Y6OrIEoBp
JG8ykRfyVlYhyKRRexc31h46LaBpMo1FBXWsYn0C5LNqV/ZIAdc8J/DrnGwGlh2E
1QBdbCaH2Ia1IiuxGn5vcaurA4sHkROVs4GswyWs8QcHiQgiWWnzMq+PFM43S78o
2+IMK9W9ltZZ/rUNoKWsr0ZxDFmGucEkydeVkWnRr+x3QKR/o4tjy1+DEI8oLMUz
Oe5NGaeqsmHvLL8txJ7ypk51I0Cpu1RnObsYl9cd8OtgQhx986ukv0sG6O3qf+Rq
f/+XvqN417HYCLWmDI63WBUC+Htyh/rAEZ4eYLl19myZGgtpx1VqzbB/H1qdUvvu
rfhSqwbprvBwdIurXok0P2te25ppHhwy/zOKpciZeR05wMBDlFmuw++jtoajgrbD
oYH5ymhu49pzcBlY3mKdIpv7/xyNWilSOxaTIfVAGtyD1hC1D1in5HPH7SF3KiH1
StYdo6DeSCz7RPp0M+WG18tJ/+IUA07ktUqLugs31vZkVr/TnxfFRjA4XvCMN+Gx
Qc9M4IT8+U7ecYYSCW+EWdrNYeiwrrwj1/nMYhPpVrwnlNF9t1aa7z6sJQfzMS7C
DiRvtqsLbceY9uhnEst8UmVK3wNeW/R9SGOOobt4E2vfUDHFE2dypKgxcvph/JHa
XnfjOc08hCMUebIZ9zcnM+vCx8pvPjuLPuMcxhCPdeDfmtoVvur7F+27mPfFNzdf
SCiEq/K3BK3DIzpQWZij5H+nCQxfyHyR9kMAxVO6k/v9rV0SHSOXhr9aifMwqzZ0
QSCjQbWv0e0ePbteesXuIKz3LFhk0Z08ceetIC9iEMfbPW5CHAGnxwpZeK3u3R7e
l7M3zTJbI9zaJYbx0p0HgUJhlD8eZl4FEn704H/Guu5nmMD+QmHeCrFGvmOSUQYk
XdgtaleW4Tqph3ZV+unSw7RRcxqAFmlyBw53KkAKMEwY6WFeysuenV9AcP75kK0B
XAznUZiHyJIaN+9DVeRgVx+E0dfyt/1vttvkFukp8CxTSBxjAvmkYMUeYec9x1SO
Z0Msikza8iL/WOGNF5KfGTmyDek28ueHQMnQHMTTGFWskWO18ap27+9bXkcwIGLv
F0Ah0Wznmb/QuAD9kJW+guvOnhwKSSC9BBz8BGa1/HWCC/U9aw9VM9ajabe4Up5G
hXCWETmOzwvrZMoWiTnQlUJ3G2WctixKsnOsUym0ktEjXS9xReYwXhG2DPgmwe6R
QQr7FfN4YZM4ueqKtEAkYamkL1seYb1GplxwJl3miqzMKyyQPoxqGRveQ4DkeVgP
NPOX8DuphOkUS4+1FY7fs0kIf1DTMPo25/sEuL6h/rh2xqeInFNN66F1UzkBBHwn
Ub+vc3G/s6yzZWyfG4ar9aSRXrTrNG/b3vVrlg9LjyrZXbMWf5jFArM8uqYzexh1
m6FPeNwY5ft3FK7LHkAtsdBME5P71T0eUbaru3qKo3uFg5phGtc7KM+83lhIqz0W
6zq+wXiLDp4Yx+XFZBKffW6CNQyj7NDgn91uHAv6S7aUl4DkbBxijnOXXh8JUEk6
c/jf1zA4YC9DDyYlkk5B4J/TW0ZdOZmWcTLZHk9KPePFturi6d86mgZnwT7I2Uml
T4a0KpLxuBnzj6erL85cqDGTuRSAuaB2PEYe2S19l9ZZ8VU12rOEI0/4dIVgqQ3a
+p1k8v2PhCAsaAhlf2MqCHRByz/l3Uwpghdry/m9Yr1tdat+L/ofUL2H3SvQpvDt
qN94Lq8vDafrnr93aXtnJB/rlKZEOj+Ol36GiAPM/H3FoxUDiFKpJT/LSyj2rXC/
58ur+uDETmbZCDtG5wRpVapbpfWzYS0h+vtQXcdrJBZQazux9+OOv0mn6lu4zUnC
eoMh0NJyLKDqFRKgrNUW9fHuHop7cf4G4YOxLyoXUZyfOeoI2aFgnJSgks4DlJXU
Fr7nX1Coy1xOx1n2x9VjApwfwiQSJuTO/j71CeZ8S55V1PM4wFeHjqZHxCuQFpWg
zORMiSdjcN3s80/qDFln2KqombqIJfAaWjX3Rz3yrJ1QY2VOZSFr1HHcqSeVr6BL
5ltGJYsbfjqaFYQFWXrGEZEvm34hD2kUc7JfJbaX9qb3L4s73tyiIXKZ4CAecEFw
wIV1YKYcEbvzuDsCNwCm22ABbSYb2uScDdWNTuJBHlO3GHmn1BfgKVqOxYCjb7i8
QcJnA1QQl4soU9o6/mi24nNyuWo0wMpfAAs4fko5dTVw9IAFSpB1fJ/Gb8IZGXrT
u1OEpn7VzinUU69iqIqChEedLDURpk1EtWCoKucxi8zQCoPggXrCCpHAz/SEuUr5
LsBweXqXF6ltgiTJly7q0qSKZP7kcLmwqkZETvagXVSiHU80wCy31E3VdvltphdQ
l5ChWu47ziEceEiYhcTpIjuHtwyCp29pZAqnkpIPEeD5epNWGSxOIu4MWGQD3VIw
sKNp71qV74yeIFZ8b/f8Bgh3gbn4C9n7tWlDPWNuiXFU6GtO62srOpxg7GOAPXCH
hDRReMJAiFblDlXxFBdnce1MBUp7D51VEF3VzCFgZA5YhtOpie4VA0uUG3xTWDME
7JTxMxheM2mW4hOejJfLQem1sdQbmlwQovAeEV1k0/w89w08EuHkIzH9kUMaAZGs
BZ2G6N/WvKJoxnYIhJuuOpwbecsnn+WCIYADP9hEH+kSg/ZmkQ7ILfiv0CO7wBpS
WvlSuBiMovG2gu3uIaYBSnjudoXKkBXY/KNC7xzE6vAPzPgE5QnlBX+YVjpOBkaj
EpbhPSfGvsvYFQihEzwyV34rBNixhLgnPQz3E+Y3qeGnZid8dgwLvbLggHzj33nZ
RwoWUZFcqXfdYwjCRxlRWiVOiU3ngFztMg0xNjdBf7knIT5Ma3dQ5Oyx1AdbfuYV
bZrM3YXGnpKpBZjZtAhiymTENums+R7YwVX18g+O1Z47kTz5nk7dyoDyEuGunHOE
8flScCrbL6h3dRrwrY/KsBLEQHICzxgJg0kyXLIUPYzmIj9Aneg0FDx4UWyxgqMA
H4wmHQUjEStBo7SEezW2LCNU6YfyWjTwFK+B4I/D/76btoU71AkWhZFx4f7/u28E
axac7jqbvqf6BXgq3jth/wOKYzFJVHPfjpo/kILA1bMH9VP1BdquZhHJ0JYBD6r3
6+YLsdes/57W0MCj4XFl7P9czweoR5y/isB+Ip6ZrDL2pdDXLKE1UK53/1oLJcEC
1LMi5iskG6nBbQoikR1bQ6BIZanQnuCK75nZN0gUA1knAnJckvt6DWebrTqmUkCV
GkvqVYRxpu/1EgTwoBIjaQGWfaLcmuDo9oBG/jsRT7vuHvYv+IUB2TeJ2RWHIaZC
ceBG8DsA9pRHSsT45PRBUHFa9pUURV0PxWenz3NtjA2fc2WP3YC8rvCUrShNMhV3
lArS8oIH5U54OqyBU0/OiC09sh0hhvddngvyIWrpigfeTWXGVfJPXIn4mbGZ37uf
TWoGEbb7j7A9AOCZNO8j+aJtzXtubfFT26Qq1vQc+EGMv9cjxUYk82PBXq8OoBLn
6oCu/lzIhHZ4pjlbqE6v/+LeX7XguNFydiFolBayUY5dQ1N4J+LnebDjIVKun6Z4
XYbbPUZQMfAnosCBlsOHo2gR9IiTbOCEzo453JtjnLp4sPnO0SksUZGT+N//tXip
filpCTINAhPI07I+lNnlZcjr1MMF75Xpu0j3l6GqShJoMo97GrW9BNkNClXQngip
jng/mvKQP6FRC4y5X/xMF1BJgsX8VZPCC/RODhxd8r/UFuXzB+Nj7Cf2wRSQ138A
rhNRRofqr1SBTUWeysvtLEp6efYiJA/9kGGjTGwx7qaK22JaDpCTjh1a20zuAsbw
vKYPY/epgDoNacqqgWKC7X7aGAQOekymWcyUzF+MW0xQPlIqkXaWs5S8S3JRbyat
vtA7KJBZXxM6wVtNGZEQqcfbAjx+QFpV51Xjj3NtRyV+hRcFTpTJ9Mon08vJfiCJ
Sxh2LrH2kMxSHVnCrsSLHcQtuPTyf/hgb2pMUJm247eWvpC9gDw6QXTT54xq4673
i7Tav8JtBtW+mBSlqyQC6+BCMEsH0t22fYD1nEmO601ZXMCw4/wgoP+Ae/t9Q9NM
EKtGoj+jRi+aGGZ85d5YinXbWkM+s3vF57Y8gUrUgTytJRWI1gv40ud2RqlUsMoE
vPhIJ37xIu++eFAR5b6XHJn4A6nS/dd1uwE5lCHJqGGG2r3ajLkwZDVpV72ymDoJ
LGLQXs3uYFGWU/8uaA2v+xliVza+JxnLB/nDEToqa2ktjqjPcduU7iWesLdg9Cp+
9IGJD1MCXbuOd4eTYPdxjDMGkf0VZz83T+rt4RJVZPXa13DI3isImskZXEHZU+ze
0NIktQdZvBQjwurstwxBzMxVcCkq0zHy1svukzWfa9iFRN8aT+yxj1v8IgkdWvR9
FScnOReGAKv95Z4Nag5PAtmMkK7FaL6KTzNLnozYPS4/IU312+RSc2M5aR8F4Egs
f0Wmlwu5rSxvR6ZXC8ygqQZRPTPOmbzvfP6qHIXkVbXkihivBhX+ZuYskzqwdEfa
xT2jDLmpxiNGKFKleosrR5qyJnN3j2eO9AduO0YSONVWdKRkBhPfUgl4tACLIA/P
0JR/DPOZIpkUfij0ybcEQ5FE4D546pfaRnoTYGSVh28Q2ECKMFoYHEfWQVE9uay6
x8SwRmgj9C20iKszKPEQ+OlwanXgOqzaPkb39gVrK/3ySuETG994/aKfqkcdzeNC
rrbVEusYyQm8Ws2ft2D2fKCrvji6CbQvMYCbdMP54mpn6C/NfHVzjoOqvDlu0243
Wwr3uNTzuFBpl0jjWcp79ZdvNxROAV0Za+MkSJ3ObLEz12VtuZmngNW9iuxSXdnh
TYDYwSy87OE1u563mt9axdqgHNefMgkKbq/bTVtCzWVHojHNoGr5j2SmVpPQOG5M
NFkedY065VlhG3ja1b0b+NoLeBC1a2Dt0uO+DvyecET0BkYr5iCVz1KlC4/MBghc
CrzKpOGudhbsjzTt7rDKwWmwtZTlzbJzuilJTd+az5Ro9bVecpzGXsrljMBIo9Qu
FQFtPxcUWXxkQNyRL3MwrosZhXvkNmUJ/7KcXSebnQV6BOolW5k7N/HyGtaQNqrG
GHNQN7NeAhfqX4Bi6W+OkkDIikHyIMabAyas56D7nz7Ri42jM2YAZYDTqqNt075V
SMl/WiTcXB/70w+m9zSyS9ALM1cixQsxeUjvuuhQtWNlcsnd/1RCQ0i3VzFByw+3
XvjKF2aM6/vcxZmWIXgrqI+Pkkn/lYw4iFAyjiOQzexZsvFUAzbT9pUDFdlJ/pAD
28Db+vxlsfUWh6EedAKJJy4RENoHmJlTQSzd4vfVhUVKo9X7QfKLhllJLA06wJbB
J4qsk/shUeAA28uJ9Spy/vt2X33g4RaP98GSRD/+EJbS17axQ6bv5iMyOinm0Sp2
4p2UCy/lwSlmoxXUqGg3TrGveFzl7I44iq+g8JWZWP9utizouYYNQRYQpumI5TfA
YQEtUYHzLQUQFF39v7qdixRHwisrbfulO2Y7xyco3mgYFGzVNVTXxRWlZOZyuXmU
l7MprIO3GJ3e6nbHe9ZDyfUV19x90l/G2VhSS2Q8jmS8Ig5qsXQT+M4HL2m4b3pI
lY7H7SbYFHM4m22UBLZrOKsqnZeMqelCjLy2kS0dFWqMK300k4HFDaSAVN9tPvMr
eD2pv4+DflH80TOKqn8mezQr1DkV4u6e3vdTA9vzAdF5yZleS7L0G/yWHfO1i0ng
M0kcOBUKIEZybYg/nDjJQZlOs+8b60pKQjOYAlrL/50nsTcHnMEgsiGs5hFasnob
aTeoehwr3/oMm7foKdusc4Ydq/+c0tbBWtoaZRgMg8hw1zLR2MwYxDnXlEJSO0cq
g532Cg23feFmbMu2xIIV4zUq5lKqdxG/9P4KVOK1PogBOk4iuWN1KwhNpctYZGet
bbs3XcQMZyuMSm+n4jUciUsoTwS996q9rqcBW+Y9N3ndUxSLULUseXot9JpuWtiC
2+akx4iA1z4RwrPnd52jrliPEn7MVFP9qwupCgin29DS963tCrAM8BKm1nTI6Ezp
tPNefCJJdwRaYd0zjBMJR0GTvZciV6FW2dsScwIR3vwrozGCissjl4oMIizlm+LI
Edj+hhEvygKgSo0rpqof6BvXfwUYsRy8iJji+Iy6iC6z4e8Pn0dBXSgRzh2KLx6N
GMGSDzNLYTio6mfsSwX4TonEdO8FTclczYc6wTpGC1X43pPzhff7WMDXFtzXTDGT
xybn0EvReaJNDBTMVcQIDNpstHCLpQWJQM2PjrTHV5dSflv3+c5DqrQLbUFmXPAd
YqZJSJNhRtTvcolBAPZE2kU60FBK2a3HRdfK9C/4F/2XyNS5MhFdZPr2E9+iv8um
bn/QEBKnm0yfxO3pG8T5KIBLO4sVW3pQhX6kKnjL97DSLQeUprHf8NUUe7DB+jIr
LWHhFZrlRliKjl5SGTXIUL5uyOUW9dK7pTHb5RSq/+vKeAc7RK5E16m+uqfZ+6+o
bztzquw+9qk2h4gsnwPjBk6E7CMW8vfhw6L7zeVHXNT5F1viPBDMf5Y2I5F7Ic88
19oOSxWM0vUgjFkoPycjvMMqR9nJQJukzMMiPO6ZkfeY80BY+Fv7/popKwnyw5k5
BNnt2F6TVF2nRPFHkMjXu7yKW4aCCv+1vMdaOnknFfUmU99SNmwkJopRozaSH25s
LXPHFPAUtII4YT0LE9yLMSrnqI7Ho6cmdo2nCpqfU6YgdOpoTSJlmcvGs8Qi53YF
hmiADEZhZjuEIqdY/nl3c7Ax5mfr4EBWxIsdKzGGKDkIc9phjhp8uYcpFrxpieGe
3YTNt360Tp45Tf0g8eHfiAwJ1CS/LbpzJb7BkkQXLj+QjaYOoteB3Jw+ssK2cq60
orsEZA1iYoiX6efg4xiFtA5mKzeoV2XG+t0INF2l75l+SJJt/RG2o1Mnx1otdDoh
q94wwolSt682TQn2XXwNZ9uEpixIsKUocqWpDuwRP88iX9Npz1syFz90ZufSeMV9
bSWsxhhLQRj6riSed5R7NN/ap1WtYg1jA4mPcsAh+cAX/jqp4jDTMJ6gVHAiIg3O
NBMWKjM9owZOyQ2X0HZE+X8OPXLT3yUXwypjKr7KmgO+o5QiZOELyDAk20PNgxOS
V0iMzrZNbBlPunnLbKWIOZaHWTIozHxnQIiR8Pux5c/+1qur2fwurKpXId1OWlSK
AD1GdBUmmT7P+XEhMN8i+q1GnYPKuFrwtZaJNfa9q/HhdOzFjpXSta13B+KYm3NA
dgLJCcn87jHCltFP63Om7Byclma2byR5uaBifjRU8AVKDG5pEqk7v9bBbS32mAOW
/UcIavfSGvJZMXxCYN/6JQcLqLnZojz5N1IjPTjj9cJdrPaS9xXSk9vkVAoQw+P1
IygCa3q2xT53hXirlPg+pasbE0X4XHHjOB27qAEpcub7dyjxXmF5BGZAm2buzaPI
JzpOnLn8T7XxblSgb1zXf/2fep5NN+mVOus4vqSd6OjUf9qccA3/ijtBRQ8at6cZ
hUahfugZGsDaEcVFFJpoZsdfKklR4M/h1h2RiPq5Kyo3yvqcV/PAXno1mulFdkrY
KcSzDMdHI71hDqZqaEhQx2LkpMtD/QpmClCOFJm1W4MZZamcpAlYPpuU5YBmCJwj
DVE+UaiIJwiqR0CFecfqktEPu7hLNWhOS8O388hOcwgFJgvn3EfJwVEGDXBAqL+3
Z/0mLzKGTV42FEp20epAkdiTVEt+pdctU2UNyjfYAf0o9duXovCTZ3HxgiKc+YDQ
Rm6D2LznTQCetwWGUn7ZySru4XTOd++u3sHXAEqhnNZb9x6tEyGo6faopuV9FVxP
jiPwF3Ecd0BKPfqMUXHp0zP+zev381Gag1d3XCN2TmBXgEjFWd/8F3vm7hDnZVxZ
RuV1CWpCX0gcTypZFtUSC8i3eFXLHk7TQ6dX4YBmKgu24JPi6R5gdtuawEaB+jqs
oxWj0CaFJEETJLEadcS8s90xQ5P8fSXuJuCGCI5n5s0l9dzoTxPmlUmrGgRlWjIt
EpYUGk/Ta/MdjBxUu2OLWAWLMFcCw0+4FR4BbQWe9S7jAnVA2/RQRZOdPxb4Mmyy
GE9rIkoSVXnFfixqUyQCx41fenNI8xudkCRrQZa4QRy/4jkGFsg8Gho/Fqh810Me
mJnYyMifg5gbPTExHSrfjotqKtpPJnfvutfu+TbmdHRyMj2QZYexFJAcEE11dO43
j601hhLKWfbTyOQGQHbbiiDmg27bAOxqa3egYa+o+w+THUHnIwU0bjzDY74tEnB3
ukxun79KPK0qu7kvnSUZAIivGH79/RODO8KdcyAYM8fHs9Y6mp+MEOQI1270vXL3
RgP6244ifkA1fSytQb1i9DacJpCVAOyF9yUpbEc4bwK/9RHUCqfqbT/+yWuQiqwT
n1qefIJCvhb2QcgKU8BWyMJqkgYi2CHLYALbqRMJWttbNsOt1sqGdPTb1AC2feXP
peCqBNcTwoQ6Y0pptugw2az4rHYCtNGNWfM1x440ryWVfGUxpxhM0qa7gjyI2E2S
zfOO08Ir+NsFQiwoeujSlDnZKN8sOTzf55QMYEkBOnjcaJmWCyOiYvun/AzMeTD0
YLs2Ka7O0LkfCCpFuMWBLwj/vxJ2zJ1HqPMBAPetgjtFI8+lHC93lMXYrJyHvIbc
L4AQknw09rsEd0Dg0TWkpmFKbv2b2TtLJA3NVwXf3yFQ/B10NLGLGr4c6QKWieYB
jfN2E6OaccC8KnJMe/QdUdoTivliaVXbVz1Rn8SRiw6A2/BePPTYgcz3OS0L6GNe
S1J2kt0YfrLAOja4ExAQdzkYoVvnZ3+txGJmV8vEdDHGmm2UvD1Ndfejk9vAArPl
ajEMebqe+hR9b4OJ3/eZSp9JMmHT9y9U2ovP00AjeLtjC/cKcgFzAiagkIJLI8Qq
xTzXy3L/iUwPu1LAni08BSpa9TMHrdY7UzpM621xMXoafVePaSiz3YSvTsIOuAPk
M+RwIrdFYaP6C3uq2J1N9CgxQRuD3Q9pObmJqY0bh7ddJxLVAZlY7t4kgh6ZP2yt
OW8BABquuKTmYuNqzO5qKl/5biAc9so2nl/z/sRTX+0Bb7QFqrK3r1h5DYUSnviI
TWSaQE9T663ApiGHVbQ4XmelAyEbMsk1lsTK7QyqagvUZinmVhYGghMMOaTexPbT
PZECy/r1RRYBCkjitlJRPBAXvMRd5B/ENm6TF0F3ooE3ijRKFM9aeaSz4icAZH/6
yAHZAIWN1NP8kLKdM2cpf1gmbmCOsGvBo/J5DALBaFySoYFuMCJPnoxsLAfjs9RW
+XeK4Rtm+cN7sI8VS2dIO0OmvgzGsuoYvj7tzZyFEmmjuw+dhNiMmGidbvoiLsV7
fA6R1D9l1Ie3DYqj9AYbgRWgBRD/GthFa/qJ1owjXEZcLcNRdhaTdqSTvc40BwxR
Ors7qyXxCSPxekSGuKhObccFNwWdNpF4wUq9Qa8IEwx6KrDc3LBxdollTBD6qwH5
X0LF+/C0nHsRbZzaDb4aMjcqg+InYAngnRstb/0NFA6aKo64c+f1j6Oek+WmZy48
5iBy/ijfqEOe3UEnH2LRyGnRQkWNBZEvHe7AlgzVjuNhScv2oZMfvHUQRbDLRnds
YNd4owEvFoYhGBJuMe/e+zhLKwdvtV9+kvaFGxqJ5Vhpf3l8OM9z3o0LSdLlWTNo
Kte570NrVsuKYurbzZ7l5e0qfRepWndG86geOOXBh2esi3gwCaa6s70Kf+R/ey6T
febNqQg+9hl86e/Sl5OnQFYFDtIBzGDv4KAYblGXuORrjZcXPlG9qPDiTW8u+Ri+
Y61tUP863uxDY8Keh0qqpWq1GwyIueMcihb/yVa+1wkB9mzwZ8EGP/X4LCRMDd3z
ZIaqsmWqB8VjK7Vo55nf4U1SR1ZrA1vF86lyDcMV5FniRHynYisYLouK1+49V3ii
hSJaaY2G+OAc9vQhxaAPH5b/Npemhcfu9Ls2prUWOET91ZsnnIYvZd7ICA4Nk/pE
keX0zURssrh8PKGOjwGzKz3+KzGSDm/iEzLsZpD6nVHVO6IhbirtjXFFXJhKGR9Z
5wHpmMp0c9drusx/Udim//rPOcxA/kkDpFlrnaXhr3MSp3ARwBEKFs+gjt1FMxCX
1rHfEOUBkHe/ADhHXnwiUTD26Yz5MC5iU45hmKtAhC/zTZNilmQhoy09vtB4lIAZ
jTj2vO86P89eY02Kb3T99bHItAurh0PCrIlU4inmPaVLH3zsXrdYmBlzxcL2xg7H
i6f9+cVG+KXpBmGh1+1Yo/nIPtm9Azmxuxz9Z3MhWIfISUQ1G0N0SPOa2dyVCEgw
OlBtVIJg6vLPWpDP3xFvtRio/GrVViUkUr1FyWCTMqCChVjqU4W9Tg1jvbWcL2ON
aDxtogtgCgW0wbt2RD6nG4odsk5f/MF3GqU7h2QpICqffxPW4wy3pIpkQtD+W+XT
fosk8HIiQhW9crXLd3+SkufzE5qUeiTh7RX/DAehG4uly418sJvtdSMhee7Jvp9k
0kY7GUJlcbUemBabyzNpxyxQK0pft40bCdMPJZhrDX702YDT8bajU5Wa6g+EK6Oc
B2Pf65HNFlT/8ckQRhZL+1AovASIFhV3J5W05vPF3eJ+d8WBnMy/6mMy6iR2gPRc
4gzSpbARzhUFzHrth+qJ7+rXyCN09z+klpN9P0NlcX6UCfrjYJpY1kmzYE5n9Nr3
4XMTN0m8UPMJRWG7HNrmfZ80Vom5QnzIo6nl9CpLuaE0lN6UjMvvpMEcGH3kaBPe
/BgAZ8LtzM/Hgn6A8GGPJn/fFT8pyUkA9n0pRRYDbgxqzBYxWKPr6yzpT+ScY7Iv
Csou7xJDNh6DAkBYmkR2I8uVEnq+vGfNyqVfbNfp545RKnA6aHhS7d9x8uewfNVu
u6QBqrj+wx7h0tnZ6VR1k9v3DK9v/Jm2gnBD2R1r1Hkzhl8GfyY3lQSwkoE/Hbxq
EHtU4CIuSyMwcrAYlA4ZWZRRRfy1x7nYSOVNMTOjK/CtqFJ8KHGAtSQJMpVCEgvK
5lywYCvk3zfjoL6L1+oxiIAaJfVJoLX/N2rvluYD3UbET21XPf9m20Ma5vVFEJd5
+JcUAXRIUyCcUJyTlBdBAP64YaxoeHDSAlxCGvNhxaguB8SZmNT4rlwU/JH4seCb
ywB4vyFyp/p7oPwi3i6kZHChfGf+y+v3II1ZX0enirMWxWScOD8S7eeJkpMB+5D+
4MEALrnorcMG2GdFvjpQ6+XJ/6xJhrm5mEknREmCVlBHvgFeZY5agXcMxMwwQx+D
heDpKTbN/nfxsT03gbkZPLVz/BQ7Ee9drolqD+j683ek4N/h0f/DFEHvu7Ldt49G
88sg92SM3LP7NhREU95h2DSXRxRGrxgDhvq/6VpT4ualoDocbvJpa+2F69g7ZFS4
xDEaYGlF9UKPoCv5fUOxDgTMqGT0YC9cK/BBv/4Wz0UVAfd7VqLcgBaJOWchuH6o
gqDiWH2wt6mc+Dh0fYRUtPByIoRBIGvmmp9PgEyjkqluw3DbQhyogrYCgOR6L+DC
2FTX7zc1Yd83/qcW6inxl9+ZLtWfXhnk4j+jOIF8SyElO44tvllFg3J+LG/+iihN
6SWnaZCz4VAmQn8zE3XcFccvEoJ1sc6GFF45ofZYne7y//zosHBa3E8+ZE3yzw63
c5eWls1uNDqe4OIFxyfcsxY2FoCXEDQ7Y8nr4krToXZS5iVgWkokwTOqJ9wnfXbP
YEG4jtEMkbOh3q9Fv8m6pF1zJVdKpJOnuWdkn/KyTrLF0UVGQO/ywht10+llRTzd
elBrgrDiKVQwmcniQbnrOiHHilWbTAhzZdKIv5VPlengADUrfhVkhNpL3jb0XTj0
u1NhmVETBQsEbZlyRJLXgrJzRbvd5c522YAUmx5z7n1jjLNPN1fh2idaBZTF+3yP
4ZdOHdLF6gWRrcG0YATlJJQcdRVfaydB1SYHTZ7RkDHqUoezXyO2TdihL4FRf6VF
l1O7xtSWnKJ7b8UcmRNLlnG8T6GRIJ4kwfPbApP8cA9j+E3ZrYw5nmvxubzFEQwY
z7Y8samMNgiOARuYZO8j6AiByPNuI5Q5onBaIzHjesw4kqqWKB0BdCfpilgkYe0q
R9AEQeXRlVRTBQbrMOOwgy6Lwxud0OK0AVgeGOyUfFlxMbCFnD3fpvsskTtAnwrk
W1FpIBexMwMsBEZQfNrgE57M/9mRugGETlo6696PXZoACtzGm/WwHZnl7immjtrU
7E72zFQ1d17S5hI4acnD0TQ9OuP4R+K6MvQf7Go3pLh/LCQFu/sePwQ9/Ezelr23
kigbICs67WminkIqfjMW3+1dHeNgPvmuSmJKg5xoNqWNZ/fP7uooCDgnT5XKBC5v
lVM31Wdf2DKRcxyzIEyi1klcgkzpMe4opFHGDyP3oq55FtFVEtHDl5dS1bcLUuRj
JZKEMumMF+J5/CGEqch/RUgxGfzKd30/M3maoqA+Kb3WowwjNrLeHtQp4l8gsAUs
igPrhEyC2J+IEoKZ2VXyDwojQ+RRmSi7HY/jmmHKihWJdKglyHfGxoVY1rA1K8gF
zT0HuJKel9QIMgS0LyS63hJu9ckTvZnG4no2Xze/z1fj1D41lapX1wteRLONM7ZH
1b/CQQHFTU6AdqU+23BL/8IaRkwx1Exf0WmQig1L5YkbhxxDaTbqtz5fnQxyPPrv
QKXZ/V+90Ct5/RftPgoSe1+HHyV2bHYmx6XBxD2peSbVzb2xea7Wi4lYfAaEf+Ry
06lQ3oiaPLVkP6DruDm68lW7nnB9WaxFEpSem6ZAkCPZrMzE0OY0W3TGgonfCcOj
qI77xRqDkB4WiVp79Lz5bYV8/ri9KnfoXtAis7cqrWVbvKVeac7ozFKgAOQLleKH
f7cStvQZW2l4PUAL4fzWesDw89keEVciUqOGLAJu4D8V0y3Is6qutCLRU8c9Gh80
NRQWZcoR5Hbv1yg3/9Ep+x7wVGjZsDEr4rs5Of7AbJutdUH6ed1ISYHwRocnAP2V
1xH3Kz9MzGmkztIx5uOOV7W+P+d0u1JFnpgLtl3T0iyF8eLn3ObY3CWJKEs1LHLf
OPzbjZ+JxwJTgnFJPkazvRdah4c2uI+0r6KYyqTOtNAYZIu8Ir0fGhi9y+A7ZaM0
Dn9CjJTidGiPDJufEqOywnS5PSX1fEUMPwWe9+C3BQm+IKk4VZUDX+ZySNeu5MY+
HwfKVzIrmjJBrVUJYuNhj2xNL+33gBS0WiVKBHmLr0tK7UuMoYask1r3R27oNuZA
Oq7IJYQGiHohbitqsaIbzYHiWjV6Orf5SaB80nNBegNg41XOMcJw3XIF8VVf7hTq
vPIyHEpgGLCuvZMu0n2fJno+Z9Buqy13iPVr+fVpx9wcLhU6pcTXEwB9NjGRueB6
rarMnypLULH51KnGjw8L4cAKZFI1llx5oxjkWgUHJIUnlf6y/BGfZkN6bxx6wGMP
EyTU0xJgiyO+qxaAvzo2gl0WGZxWADX8S+EfIrdsIzYfwloFOC9+NxenAFbMNr0X
Hh8XC6r2EldyPvYxOgrGy9YOI5yyNyupK6pqQpzI1c5ZZg9JnHDb5kgBe6/6Ug8K
ddPnfuX67wazgUi6i3DNyMR9Q6tk7g642c63T97HxwHFsipCGuuLsXVOMNoxKvq4
+51wEaQUtjIqBtCwqiBtPJFY2G8lDXrcAmfKJlKlsre9BlBQTvA2DtnFSgKaCOeS
45UUm3jAcme043APhK3NY7o4ASeayat/3fj/H2CHD4EIpTDoGoIhop0wM8ycnbRL
4/l2cQQIyHIecurD/mZMVgvEB50uVf+JLa/bUwp2pQ4g1wti14cW+2v2mdUK0ujK
a4cCS6Cs/ggECOEwnrlz0SRsrZdXBTWt1zoibMKt0IVuQdJEmRcLCZK5r++xGPOV
lIj46zgOoT03qkUUXjPyQTGH804thRqKdSyKMcDNVVTgYdkuU/vcj78NRKFIxbE2
Kg04e0zwz8wvTteu6WUR1YFzqMnNo1M6m7Hs+2wv9Yt235KcW6Zs5Yw358e6BAx+
O0ai4RPXZpZ6xtmofH2SMZWsHZ4bQmZeq514TtqD5Ou8JCf5vYYdZp0txfBM1IYK
4CepwODW38UxMztI0Bke0SNkRWmKK8To8VknJ6hpHjiDyPowHDKuPPcO4gm7hV9O
evfOsn62Blfaqdyia7B9tH/kkrorJjRm0NPP76Mjnq+WmOvpVQxGniY6NJCmpvW6
EdNVBvGf3D/QKuTGcu0+wX2CCHrUQjn0MxeI1rTcZE+5OsNq0vEAXxNW5itLMGbF
rTS9VVr7SKtHQETekxX8OoOIZ3Tvz9yMbFT9CoVXhH7I4/bE0CGUJ4X4ouuN2dza
R2xam6YmRlkp6AQSAdxz2gtPt6Ld+vHwusENNm54nzI6m2AWTa9ThKORzy1MQQWj
6oFabZCRT1MOr7UD+nEa0KMrgrA2PIwWmMBN6NPmASAfnbNzCuajEqSQwvBTUvxt
f8OQY5HjGiYXcg9rcPLMdBvYi8fBYfE/IFQr10AtHzLGSj8liHgn3k3ffSHU91f6
KF2bt4AlHxO5GUNGW0hoC7LYNotSTouBx/JPz+w1y4c/tRW2UpvfH5oANbPTm/nZ
7dVG2T77ClkbjfSGAmkozSmXe4rrSTRX5hZMFHWKE9ROKdftDjMTycS1uAmvN25V
3EQjoOazfk7YCk40H5C8hWyGlo/G/gNpKbszqbNS2skLsFancLy0L6tQX0J+3bRA
k/OjOCEviIIrBW8YClMO1r6unStdSobLIJDvXK92nGNQZR5+rO/7x5JbcDJb+OKB
JoyrgciNBC5LTl6Y3oLFiCpwoHXcG7Zi+pO5Bbvd975fz7wMYQex9ekHwCogvwH+
pOx5ju8pCPBajavUqElSm0k60kB7qojtjzwRzGabRJGiNoNAoSulzQKIsl9+CQu1
X1v2r2TXCHQgG80qz6rX1kwd2CJcziL1KOpcLQsLnR9c50kTIN4P64aKH2Cggg8N
/5G3YEUcO/XRuv9IJOu/KP7QfJEUuMmw0rfTek8VjvkLmsSow20soKo+cbMbxRC0
Y8lJBYw4To+LJ2fUnbb34bzEqSurZLuq+rNXX+oCy0fXj1salWl7CKGRz9y7EcWq
Qc+D/ULzhRUmJbKxU2Ja890DNPBFik95z8ZOeJ25ystRB7obWbIg1hkdGrof82JJ
2JG4g3zfk2pk2NpdQw5Pm/m/np65rkeahBqa9Z5mS89DpswVm4xMCI8GKZxZy/dw
DFWTdUyHptA3/FXGBjfEbenLtdSoBONVIiLbMqlMXGdzcz94c1wcuTNVMa8ba2nt
908qWsVj4pAh2+sYWPzTJ+Zeaa6yALrDE7hOEYqRN7Q4fhRxz7J6WrJltMeFa4oG
7/HfsMc52jdrWjtBMfDLLo6HTbk1s76guoJGmvaeZj8fagugVsGtJg3sexgWMjB+
Utej7SyKg0m5G70Wl/+hk5qy0wOKhEo8JAsiExA28otJUIa8FlSqO9zHHjSoepgm
zYL50ab1P+v34HqXIopKdGZA/RdS5fTTOGZd3K1FiInVaVOz+0QXU3Xg6Tt//p7a
N+XbkipWCY1l6TghjMwXSP0Py4GrQG1Rtmb9R5ZTmF587TQKm0iDlhNbfNVf9xKH
rU/Kosx8q0S86VLQoUKreq7zqGmeX3akowe4kXQ3K5AAHtB3EORiy/DNc9FhOFuz
UU9fge+SBRgBetiVxiRm//pFh6Brk+mrtdxcexySazPRSvJ26Tzc+ucxpg1WcFT3
SNPgyHH2/QVIWvbYS68JAV2GfATvpTYiokQZIQvMh6FgEYbWiRdh4006Psn0zt5I
PqCPAogPlKXR37tigeLhYNpHBIgK8dARm5xS5wYGohPZRObqSOmK8crU57BWs63Z
mDYGXdiooZZNwkqtSWETYTxw2GxA4Zp53aqzoNaYnwhap5ok3Lh/JB86mX7b/cCJ
adv5cvotuT1YZWCnTLzxvxBmUmCWv9HLkGwiEEcsCiAWH9QdvdtwPrdZ817qS+6o
ViCGCc2WDwEDyv63V4CmdPXpYy2okG4+BTfrTL2I7nI5HBayR/grLKLQuJpqQYMR
5SCwH+4yKTDzhvGbAWzXcPohY0SHSdxLOi6ArxxHvTYcD9vhwo7ZjjjxyDYhwXL4
akf8sdOMXoI5id9ocdwbgW/uWV4IMtUhb7ISdilc9qmA5DaEOMJS2kteZ9mB2Odb
H0PeYDvBIGdzu9kwGB1yaMRO9IWo4m+Fh3acIs1VdGDYzm3VtKbHd3Cb+pWnlfgW
K8OqAIu84jc3xxQtA8K0lkCOBgq0jk2YESf+Fvf5Fcr9RJ7UxAPXtmbAJ7iezSXz
XbtRQTTxV4Th6YDVU2aQpt7bcAey8ESFC62DTU1LPtGLsvwzLs+QdzwE2fRGzHaW
sr1hPNoWSbthQQ7EESEDAFgCh7c4YzebnuagXh/qwyweJmWOzWOsDuGsnir6lr+l
eq1UuEDNTRCGzsre30EyGd1uv/psEQL2dxHJNnB3L5C4JiFdzcAgWnur53yI1R09
fMyepjCyLhrtJTYGd9O0a0R6AJV+6oLwyH+OfIUUtEJ+eC6EVxNdHsvnOdSXdI09
m6FhEMGuJQcf9Vo2pftLvQ1le98uA+YYFnvp+BrXsgjcUjcLT3OpseHb4LB3rtia
DLQnaCstpWiupI4vf8JhroBkk181au85phts7k4XouyfzP1Cq45iQXlZhm2dCE1x
4dRK+jkC4UMCHLf7VetC2SfCXQCWQSPQaYPLTkwz7v27FVly1qm6cTM9W3mc+MkP
ZD/UR4tw1wfnHbR2lGZzIk25W/1D/D+OcEoVdsqlvLxFKiibejVltd/5dxEa7wP4
gZAfnfzlgUYtDHaoAbgT/mVAbjD1y0B8FkIFeBDTArHRVS7R3RMdZp2pFySI2V6f
gMfflUM8nU/3g+YwzY1vSMb8qi9ojazlIeyG+pW0DxBMeoelr5POHDuUUbg07a2L
OSIwB2s0LIog2Inm/UbdN5ymHSUTwG+alDaGs2wExolQxMJrcsfbKRVXZU9qNNgw
Fy9SRpyBJH66gvaDICxi+RvFoNwBZE/P2PZLh72xhP31bOcQuU8HyM3z+d4lmPtO
Qm8qt6EVv/zH9OX6r/wVBNJo+dwT/ov6Wsm9carUdY5IsFxmNwRnjeajun5WEMmz
eIjfOFcoLqpVA/cZLWuLK1KsZJEzd/eT76B2QAyDZ17prXCUs8IRJjENJYn4PIvi
yyO0r0tCpJ6vl1fMflMf/dK+7y2a8pA6Q2hsGq6jI6x/DNN8LZeRPrF8JmdG6jEE
mJb3FSNZeLv4g6yQKbSMrcZkIqHjQh1jDgBXLApptzMMWVtzWr6RoBzJoOWKAxSa
w8ZiJIMVBPeYkUnS1hLwvLEjGSzXVpSs9ILB2N48w59bsvJ7LqyDw3hqwDt8src+
9hsSoEu7nqRgpg52If49SAp4I62SnUsgteOL4VbzlCfBCKK/YZ+IMSmwCJoUa9k1
oNiK0kE+iAon0Jdh1k5TsvwO1C2O8qr3AlF5p6GLCLRNDubbiYOx3rnJL2QQQ6oc
wAFssuKSx9JjqniQmDuVMgy3HRuq0Xb11cI1WxHqqaTCYxl1fhR/divDkP9YGRJ4
xVWjTiIcRdiezwLohiWL7fjT8BjVyTDoAi2P3lFvGR+mB0wkoBq9q8tEUacvRDWR
ni81XJMOku0alYs76CrehRvij17CgXRCmjZG9iocC06qWlD7JIWo+RJUqAVw/IVA
RNfJp2S1cECh8QIYK8WcBkMjUBgNy+rIHuG4zGE1syzJ4rHDM5NwyuzLflDOTcFJ
nY/BwEuS130hWFD3RXzhHlNBqi5J87o6SVlfoTyUMX161DKW+I5+No14q0cbF79S
NQfxfoLt2plEJvk7D7Dwfg1S6BsWlTXUTiEO+UzLW6Fkp8YykMmJNmYgZO5Ew6SX
DHFoGh0PbGdzAPwnGiqQRbgP6FnWkS8UFHDn5gsxi3EieC62R6Fmm+KSFWTo4xnQ
GtLkmzoxgAC246E0ZTyf8nLEK1D1LTcC221Uh4Wd3Auo3xYhKxqxKl4CcOft077K
z64UeVpET2gTXTWuiuDSx6tX3USfA9r5dkPYDJPXrYGa305OueyYQFeA7K9dCBLx
QMyUWwC+Dr075Re4EAOV0Cc6L57+BgvXXseb6GBCR+H+i+m/2S3gTcpj0ofJJbsc
Cp0efstEegXwjyZnGc4AIM1NdzPFEhahdWB2jTBgEAyJAdIso2Ldt9xdYBijUdns
zCS4YPDP7Ry9Pi2RF4sY16QDbY+2IQ/liyyyi+p4XJOW3BZzmE0u4+KFVytZtryQ
jhUmR4Y8cWYpDgrSGlPOiu2a+9nUtGM8LDr8OUCuPFvReKTYNuj+7VXvbgFmPiTO
4zVw6WMMswa7vdAYyR6hVmXfWMhHU0jxBwGzFHiuZXBWSYa8CXkQGXW6DcO/8vPZ
maknldQ0JAPDPNdeDO5RdRPt77D7gEAOr+srXTExXyuDCapKz/Xj/ASI7qO+2d9N
qiojUJr1B1LhgE+FQ5dzI+GuLcZ2E0+ck1CxQLNCvbzYBu8zFgknXUw43ehOXO/N
9tl7FurNULMLN6KngWr7awfOenasRWVMKVnj/9ppV1/f6qgfv68KnBw69k57f30D
mzU4ITWzWEnoS4muMcPR86zVpF4pwfDW7M3JB6MraLMolmOfTKa8k+/ADtIdnyHj
0OUivGE2Lb6BFnYq1UfjRCODNp+o3IhbzRpVQpisRvR3OoOmgmPy2gpFfxqArJiG
wD7oD5ylc0RFsDQUVNCPXsTdv1j3H41EsLcSDgpmdDyBAB5aOyFW68Fz+qln/6Rk
7cledwk5doGVa0ylAd8+NNEX9uX+arkDfNITUWNy/pYJO0UQiUTp7xyVixCaN7xd
4JbEh8bznIDNLTCKI+PT+lEGmQzFzuWXtAZqo8gT+6eKNirIbBUQttQzDIjpYLRx
z5rTc9UrRcadTyBmbr3k4xyLv15mSjrIrFg1/o5EXLf6q0m1KxQzvJXvElHSLHJ/
bIO7WPNOpc6I6JAMVzzcJ5UCQJAtmU8fmiDM7vQmpcKh241Dyf+272llg07Fgw+N
y+VFEEoYMqAi2l21DsNgspQ55oop9X6cBhq5k8ojemMaNy6ztNbIbGE7gGA5xCza
Ei5GdJhijbp8dTjP2pZgiUpEW4rTYShJofOp8kMxh5k4P4/cmD9BPRkxPYfoSu57
qf6I6dlRZPVcv7ZzzCF7jEhPghiT/PpHNUDFww1nhf17YCG2KtL/ahEswC14PpIA
C7r4mk5Jhy3zZYnh8K08uy7+LxAsiTXNaEhBQjDCE4DCsaW3areS2lc4pLCSwkDN
+WiMe4+rgBtNPZV8c7Ucv/NDVM5/K03HGFEuHawp2vaJj2RHjZm7HkABGGrJBmkd
Hem/pEIXlvmaLVJNnDnpmM3vlcuWhjwVrWSdlgoFTKB2l8YLCHhcVYZ6VmDH30kO
vHQVE+s3zZoHoAngE//ScF7xri4Fi8LHAuotX/d5dIps6M376iHZ4A+w2AN3IXqQ
QJJSmz9qeZYy49Mkzi3wOTkXtUY2VnxK8XuHJreUWddmTdUYU7tLdqMUIRdxQqSz
GCO+DdXhz/NwgwBDGH5t2YzxSm4fryBKezf9bcM/tnziHONS+zISyMPOgVok6ter
wJCGe+kBzLlbXfKzObuuUNbo2itmdBmD8V1VsrzSRR4IQk7gxEXXIXcxlC2G2fdF
JWaVR48PpomHYtZsKoMJrZltakc33YktQ+4H/FXCS3yY4t8OjF/UX8+3GPSCYv/E
ow8VWwJVM/g/28NTX+g0s4PbcDtOrKT7Wzesjz5JmJEhdPsPSnqOmubH24tDiBLV
bplTXUwuFTWfUMJD1pvKWNsTdnpcHiUr8QW9r1ufpf92UX0YNhHC25kcjhY0+eSD
VtIn/7dCIvKFXiyw3DqqBSMdrTae8ICJrn8ysEjQa4eOqM/UVTxBSo9OHoTC7OXj
L4IXjb+HpcjVf4EtyU8hmB/cowOp08ymkGGJ6WqRbQDVU4iplyzGgUZsjwvoQuX2
KjnEhPmc9Rf5H+rH0p0+l4fRlw/bMG4ObauQj+xF1/n5eYvFd1s5l6X5957kmCyq
mLo65LehoYHTXzXBYFMevnG1yPmzNaQcfGPTENk7GIAmuc9xCCkgNud3Gi5giU82
kB46fV8Lcy0GmLQM6rwfo6PH1vprliyf3x+tZIx5ze1/SqylL++PUzUc/HwLNzrU
bgeHaCp/5vgLifmPfdTrzJrXuLgZiJb3YBgq9sduvE9GGu7SLJPgB6+Bp3pxDsQP
hNiN+OrFYIiYTnd/DAIi0XWGiJRCIh14vVe3AIkEx3vhGvYVCXDKGTwg/I7N+ccy
2YwWdObAi/RZBisJETtqABCVB3HpQ5qTgHvXhB8UtSHKui7E/gvGXIQ/wJlfv5Bu
Y8MRERzDO6TCO2vxGs+Ga8kYWBd3/yNMJQz2vjShf+UOSjUvE6WwsU1N5NXe2ecM
j6GjdYrcFzThX1e1bXOpPkG3IxsTrg8uYgZZ0BaXYHqP5y4IuEj2UtE5EHLhzPyI
y51ze6BjfEPvW/AdLmWzsm4XQNTuuF1XbNkp3uMyqrGHchbp8AQsH/M+4FIS7vKb
9fNfDunlXjtnzp0uBSUL5le8z8HKCF2IlZZ5Jeh9EnN6sU/EkpnZphBU+4SB/uQO
NJYYAkE44/RYwe5P1KQTUJ4wzlFzbabu2jG3oCAHa+4vUXCmz5mf2PIhB5vY2MX8
5F9ckfuO9DRpjS0WO/VdCwldQas//6dsX9L0L8logkZP1+AnApk1U/7IjytU3hPv
qsasfjxtAaf+5sTCR5OLISzq9wv/0+fxHxjCSybWONpjk/PBIpMfyUtntpugAM0r
qP76K//rS7MTeOcW6gjIP0NyxZR4geZvQTf3nLmCtF3dzoAwbH1J/QGFwuuvl/Bg
FIRnITfn9QlM2br9z0R4aaPu3orHxfYMPm7sA5ZUCw92UKa91qS1o5wKRN3Yhovn
WF9OfE3FatCQoHABRkU2bpLCqTd8LqEXUupLKft0KaQft/lELcJV5Zl14DxPklo0
GE80AUOw1KOHGIjtj6VrjXrDHNGoluHCt1azaO8IIsX5mFjUpI5bcPyzpB2Ga3E7
qRjqA8GzAIA8M4mE79PDJw8vx2qn6/OejjLMUKKLOEYjef/UPXhav1KKzqMDSgI6
24rKx1iD1mc7dCTNwYlgwFvfPUdBwRduqeVJeTvWXEZv8P2Kzdl33vKxWqfsOd4c
aRNluONoUHuGqJOAC7at+OYglgKyrBDdqSELwLTts345tUH1szMli85c+TP/PBON
FZvzH84RVNCcOb+tydjdUljcQEZnVO6rTijNxodIc6fOQv0FTSPojJLmw25ueIUm
epP6UkKkJWbTlSAQJ0DiwiftlEDgbFOS8fdTgbuk3iYlZYDe2CJu9gcCFvvAmmfz
x1o+cJeCWcNbBrV6sPSuXn9IfL203sCb7eououWKZTHowp+zuVxg90OkSqCjdiE9
oVcQZti+do3yg1hARAo5YwAMO6BQL6GOxeCtKFGf4oCWuqGmroM8dOaaQrdpVsKF
xeXuB496TZTveIlydwOF/dSnNULWHBzX1+trJHZamA0VMQtmC7Db2kTDvB7DXW5R
M7FGisd7i9ADeJ4XfWM1g6CbOqJhJWHSnohMm8Rx7bJ3fPnZro6+UYkcgo78mPKg
W9RLGJJKIDMkmUX5BGr/ljH0Hl4+Cd5tuAwuzj3taIcxE2Nwd+lM/cVJmSguG9+n
rSlZJKL6J6o+uPekPEFNURaNTF4uElHBBsdHkDY2uJwOl/nsAENXMNKB2YLmzr0W
rnjLFjMEnb7EwK8K7i8sWbJFApw3t6sKS0Y/s1SdQxwhPet268SSxjeNywTyVrfD
cpqX7fgRIEiHKIrxIxcMLflyhuJhK9N/wMrDHJnVPbdUf0FA8h1+Oai5xCtg3Q9M
+/I9mDJEm7+XsMt7GLRGMffEiFfzlhUZvKVyUCiCBaMCcEuDWCOhVNomxOjhHWZH
cvyrl84F3E8IeEboVTtzny3b4RZVifDm4ceYgHCwoZ7qrsnvHz8MDnP//9OkWlNl
pEbEypXIKN1GVHBqslNQIx+3sAKtWuYLdxQ9ipsIvruSYhgT4zzVlqOHhCrt1P6m
G7T/uXKYUpxpR34hqp1lNze8mkdMDkeVQOoKjk+BFgtJeYhL8xhuUbmgpayBFdRc
cEBsAg+Qb5gSc8jmiRHFDTZ+OYXaVXu/HVBxQ4RUzQSkHu6jjMXqlkA8scnZ8cLr
f4Sm1/Gtb7iHVj7W7ddvBMViuCBOKfH5YZq9NAop2me5j8w4m3HHyBqqaEidv+f3
i95SfDCTVDP436Yc7cLnitpHmkMv0eb7hYFzmn5YINyviFLENXaEXsLOwd9r6C/Z
Gsmp0hFajd1If6er2SRxHeKQlWLlx21a+alORVxZZGNaQMQVneOocpX/fNMRnfz3
8x7Gyoq0EgiAc0KlFf0z170ALofBgGW5Ba9c2EvKqjrBKEsiKzdaqLo5LAgr/NSe
SkNsp8KvfYuQR2ngDNli/bhg1ERfJL8FA0n6YDFyX1SMPV/9QHpxta3RDI9ZkWV8
3Ix3Q5RE2FwYKZBv2a2IrEzIPbGjZpXBP7kSZyDKccZDOPvqui2pHUbqODCC29pp
Az3jAKgwMmuBFTkhgb6e76ejLIvcEftzaAUTj7vybp3Ou1ykUSmhfUZyx2ErtXSp
cvN5bCdFYe7jDUDiclnmSro+e+ctPzq6GbxhgltIhFzMbbGGsrkGOK5O0SVj7da+
Ipcim8Vaqxy5X6Y8wu9iqycmgpRk4fpLlxf/I5IzRskRjfPinYybXgKPr/uov/8w
DvOUMG3I4zdFMhLf/9Ar/sCg7wX9QQgMhhf7VfEu9R7NyJY8cJk67lWPVDU0iyie
xOVDZVSH3F/w6cDVaXa2eb2rXL1ijzpf7wbkLMDkZabW/G+HzWfcudeyFsoFtWJW
+AO84oHeFmWkAxEzG7v28afWK4uMKjeUOPBDAkShR5zjZfgoQk2vm/erNlfblDk0
Jlv1GPVnXEGVFYlML1TgmI/w5VVsBqIDrBeKvyABP1nBuVKD+GFWtcnSyw/rUrU0
F9DT7KDG0hM0gkTFGwwH4O8/4CQY+JT3vjiWBl4oWgrXmkMpmItb6qXA76J9jziC
d7T5kO6Tx9jimZ+pir00jRSAEccd2fvTad1jjjBWBsB6Xu0EumUYOdJpTCwuyQde
K0FCkzJqot1hn51OTbJNsob9YRZbtBiokVvmYAOGbOWGa+/ckV5ljg9H3bo+eI40
dAoBV/FrIhZ3SU0qoj5iO7K+wG0ra4NYMeakkng0LtTYwV6ZutM9+Q3cLiJrrfP3
s7XCW4PBn966y0iYhh3KTaE3JX64oXEzLsoQPWyHek5iDwx4f+a4zoDS8KLO/GGE
Yc5fdOf+GD/ali1wAbUUWR2CAGzAbaG4FBik6XBjagTdiZfUO5klgtVC4BgW1C0r
SRPku566ip6TvY1fE4KN0NOfbbHEAMwaojtDmjAiw0I7dRSJTyEwMFQvRGcfglA5
VJDruGWS5QjIMQuQv6iTh6JE9V773SBaNSsz1pKNbua7c2id1fQPg60tYONGwl+c
apqDVQz4gZFvSeqtRKPdrXCphqo9jzwjvpfVZnNC/EKrJmXAGzHx3T8gtfYsCt8r
bA1LDjQw2sw3H3vEqLdN+JoXrNteHeotgkAS6+g4MHqQsQuSKqaidpBOWwRENmAD
FcgD3UCup34OW/JFHCAZ65Fpx2OH7jMGeLtgPo2voGFSViVtEyGV5B4nKyeesHBb
FxsVEUTTmj6aa2anlsJbfKHwINg5foaR2RJuw1s6qdurEGfQdTg5rZNImhTBkV4g
2osLLC5fU/KWW/qSM3EKvMmjfz42OFpz8hU5MPWnrVrpY3M3eZh6gY8xs3BREE3Q
FuAE55lAX/RpqYo2QitX6TcDlpVeRaGGPy9Hu7yP9wsgPTyYcdktQ8ND2QLXtPWz
sAVWuUJ0Of0q8dGF8iSq64eWIFMT4vuraKl/h+QFjZs2YfVr4YjGx/FzcSrMBpsC
ecvZUVv7+H+ZK76OgkA51gLmkQKQp4mt48XOEkaFFcN2Vbo0cNQ4DMeR8GLM/KFR
3ztmbXGPOu13hYa4w7otQkyBmn/AhedvB4y04CUsdacnxH2Ut442aZaC3z94OGuN
CHRip4AMZFPlYtfPYbiV/44q2NGux95mzZPsnq0fciB4KnVS8AbFa4MsBwZsW50y
xBfObgLIuUHi7IAHal2f0nFzl7CsWgOCMSXVOXVI9b1pdJyY3JpTYEGcB+vz6ZRp
I396x+xwBuzgLNremfEOGeZDB1Xwq4eksfzhDzgK90H6YZQUoCpHGmL/8IZfqDCp
XH4lUKjOJ4l9g06SSQx/QxazpmySCsE0dhOcMYZmgQJj4h71ZVQTcbMa4XM4Mxpd
cAliaCaRPE0hzCmYiMzgoVDl/rHhxwdqUBgteijIhgRUJ+8bbRtewVUlnf9SeihP
l+3xpXmcPnzYemFdNhFDkCZSve11RiAeCHA6Ebf2lwI8unZ5ZCJUo0H+xtJB7lcl
XB5Osk7y4x18PCVU56H17NnGfR5BiIHj/tu4pD12jZrc+q5hZgGOqRlAsa7jqYls
/WX0QAAHUUUTghdye6Uyl8pQ5aohDPBhCWeWwVxlfpHWBAwd4ivyWLZ7XBaHBx2Q
6ggN4Xlvrmz49LMQG+SCeX91Fkx5FYbiUYZwVz6fvdvw940Q5Dh5YnBXpVAWfUht
Fq2qSRnklRurxHPwgMzMhUSHoRo8k0ThhaFgQNCmDUpjc0L5qyBdSnv6C4gocMWU
y/u7GErU+41Yx060GOZhUj5mhRYG5hc20CAWePRZ2OHtR2nbmRKAURzOkoXYDMGC
1d3DyeIrNeZBnePafHaFLqw85rD3mcWfBko/MKvYDYwzoBgo4SPmkRcWqa4r1xGj
uIQoQUYrL2f9mop6dt/+Rhc+Bzrtju5469L4XErEOhEiiQwL3bv5EMKqLUNx2lXG
qtsjH9tOH22Tos9jYF0sMsQlbHi3AReMyP8ke7rciD5v/UO4/fxK4Y3Sb+er7uv0
Tn/8ZK7CGuObtDCG5n5/QXomumdvXcKO/bL0E2FXtVndXONQyIxmtApeYU4de8H9
Mq8RIyJzITST84Fc6VjOqBHcMQt4iDqtWtW63h+Ty+imYVMvVTTuC/Ubznm8oMPJ
kBuwUd5nqlC/laH8X5aGQ3+xPgkhVP8DUMs62t1aDEQRem14S3wDMAUHpJGzBrTN
Ocy1gDTxcSKmOOIrBC3+vUt2brdnfdNir7fZ/S/h/gtcGZCnkpLR91xaiULjMmz2
doqSs1cw+2ZLT/+dYfLMvjk/EwNzLQrLqfCN/eHhCyEFP30b0hysApyYjE26JSMj
KbVgt2/5XDsyhb8VrySj42dFLgD265Woj9v+r5x5HMJBg9OHk6kkZuvrWAGe/3Sz
7Xs7wVBRKQJCepCfi51stn/WDVzaOpuqg531iO6PH2wktu3wI/MVqYPhcmnmyfa5
NR299aETdKkZj9jG2qWM++Fq/somEHCwUoUYMeLdJhxu8NsgrwVsZaBMcyPm5a2E
icDer66zgUcY8olZekb9UUsDaKPnlGNg1hkz+Q6vo2ai94QzDhLUL2bsO1IxFm2d
f0PM8lhvKRHarlP+jSWy+B42MUCQeKY1Y99IGP7Wn2K8kkA/qJf85Sdkk9cQN0De
/L2ZeULZjYduKtZj6pXUtnL6zv1ZCDC3LWtQ3vc5OFcyCWNGpRIsXJbToJDdeh8a
1WOSFyixx1BM5gz/AAZ7gDFqmcTvXNRIZf/CXf7sqDYbmT8/wgLdKRAr8nAGQsRK
1xlJVyB2vDarDT/H153231N//7p6sMjKtj5FnFLy0CXA8UDyFZOFBEWN5Y9gxlyR
nENE2UdBHpPPqOKwvzEU3xiKUgIQPwmTqEX1Dq0EcSb9GlEuO8rHn6qXR9H4C8jR
lyHGLfzfBO4RThNZ8mzVFmO8Bp3ybrVAEmJEctKDvzkaRPHa50eWarYRZxGl7O55
TZXlkSi+rXcmxLR99bDtTH+VHL5tin2wKcNsvU0JFGHz/j5wi41VAJeuNqnVWqMz
Zd61lhB3Xa+ZreOOEixm/nk2kgjj3OS7C0afSYu+4XzSJGITLQgbIEZkTbul5Ban
AUZKmjha+61rZ124fD3Tng5hFdsLouTFCZsXlpMlOFw5MQEIgyBZiXWT6zMPzyRP
B7GG45QO700Q8P1kjs9vKeZlI/8XlMlI60z3sbjSlc83zWmeYFwWUz81OTCuPWDV
z2u5XDBE88wzn6I3b4gzd3121ePED+We4NU/zifPANgaK3IjOkOA018wfUdVvAQg
CFh3deAm2GYpEExliIlbX1k6lMHDaKKmvESQJmObEH4Iaux8rqlbzGQdRKQXm0md
xI8d0ymNfJQLxA6lCRZh8d3v9W+KouIzyxsCGY7MPgo2HrTVw82ViWn39l6ssfD5
qU+Uiu+Zlp8PxZOEJBYouoBsqVnJTmi2i9YxZYu/rhoFHay7sr3ij8YMghT6NHMv
cPeHtJTFAR8+N9ee9hBTKw4V62O0TQxEZDlVfgkcxl9DYyBah1j3z2P2ylE2eODo
qpZdDmodLrxOFmo0xorY/m9S3Aj5wb+5guRp/521lzFfkcAx+Ut1zDVOkdp+efTp
vpASWvHMHiCGe7WQLidg3920MogFiRxGGOy+zjBEDx/exWVBTkpnOw/8BP925Ok3
5ii78tMrrdoagrHXKfmYWW2RH5NykQPsGJkTgMvrM5+nJGo4kMdKM16nFx0GW0WD
zVtKdnymFWqb2/TKy7jH+rmyLC1j6ZV0bLwVTZnD+BqUfERQAZ7S59HaIR5+mC58
A0gDPts6zXO0JDksuBgyBiDYweh0tNmnQ+Iv9P6DiAGp/M8LxQ66xNnLf9JZ5Otp
yQAU0OriCWnfGOC2xXVTOBrfh/EMCneaaayxxrs3IO2UC3QaKLjGkcHY2vAp+gqU
A3S6XisvfGsssuMz8VTOJAw9049B6IrXTL9RQFnydhfJ6bLyc7V7OaJqoNagHTpL
0eHs1Z2+czvz483gQ1ouMkdGzGEgq4Tgu+Jga9Ckocqx5mETWmQpaoQompGAJk8Y
cdDGkenG05UMv3Ry+20fnvxe4679EYqXNyij2fz0JQvrVRN7/zmP9OGlD2Z/dEYV
UdEaN25Hs6tdQ1hMGOV37TT4VpYbv5YY7Q++vAinvqXO52TGZv2saB4l67iwC1jr
PVjSEt9t9ql4jvY28YMuYbBqxby+KkZIZvuECVsUrantOfsNGOpaf1UuEj+HE0EQ
MylhIZss3rIEKrNX/9lrm/9TqQZZo6KFdlzezuyN7huEfb6e3oVUH/T2XA1Ptnb2
yPLah23QNKxlEByyWwA4Lx5BJr3SVcl2A0Zq2V9HHb8ryu4a4bUZQHnDaZLsh0oY
03n2ZYtEe74veuEpV8PaKYNyclCAsPTeW/1A6mLuyH3LCwqCWppLHrApjFTyQT7R
sUcvGMaiWJ/yFJ6DFVUO1CUEBK42wWUUOzwDgiJE1aNvhNcNWFWIHiwDHSpz4HqT
+aK+tSyIBb8s4RWrx/1b02oJ7Y7thlIV/blkVCy4tQakGcLIDpR+yyVyy4hkFRxI
hJdTUoaevvSygm41+GGENlKLXBrv3O0dDo7OuTGOuqAx36HDVXaKnC8MtWVRhCBa
6ccuAb0Wrc6tk/3xC4miLZVxTe9tubh/SMQscOMcJ8f+JH6dKZoAxfAVwtQYu0VJ
XNtjYbtWlh3riOcVorBtYPW8FAvyVCc3sJaN4IFy1GkV7hXlSyIunUn4u1xGXARw
twYhnD5C7h1vYNGLOsJY0tiaC3qTvsrbmSSpIvAvEnKd4KlRu82P71Nt7cDMBC8U
ftSelgXUBlOlaEejNj4l9GqDimy4BH3cU1jC5DjkSTOL4TVBVvPu8hvGcGwzga0K
YDf0pxb1bbIvS9OWAZJgnPSYBcgyqn9pwx+OdYrDUpxZzLDcv7dfXyVPott+MlZ4
8HjTAOVmg5Vo9Ii10vdNQSjeNux44rKnOnYaJOf7rQBrgbwrn9MtaddDa/acYOaZ
hWx3/d0IKwKOzsv7hxguZ8qh6DUYs33jSGHwZdY/QpRFwGICp1HaQPB2wxtU3wk/
BhTGmQ05dr0neFvemPnAdtj/w7CmEku7TbkGYM2JAFrLItzUeudAjGmMQ5RMF0Ps
2+nEwxfHw6bAH5QyB3Tyk0X/tY/RJAnhxc1CTKOZ3V8ckqjgiqYEX42tGBJ5ib2V
Pnghom9QvGVnf8XrKVoTeYkAUTY/BEScgD1VNpCRzGmIwXUocWNGBId9Efr9XlSA
brgusLsDz1r1gLHG0zq4FPppVY5BKzKOVTN4CenPui9o7i/pr5IlhKXUJZNzv2V3
WrOEO0HQ69ALOPpoYmdiFeTyk6CjVfqzGxeGYtkUBIESy/lmYocABoyJ5y3sn6vl
cyQTe85iB2fNU9bU/Gb+MdGbMByxiU+7NAnMYLijMso3m33OT/X31yF8L7ywkc6W
6iH0mSV+ms4Ne9tXTrFvHz6dFdgoVCCKXJwFF3PiLZ9ipiWEqsfD9fwrRuFOVgMO
tnI6zle5FOjy7SnXFpF0JpBGSZ7ijoQqhHEXh3BbObpo59DJrEVHu0dEevf5feCI
HTUcAhKAJbkPSQPmgVqeyztWF7G2KD1D1J8wYbLAiFXzFLPP6KbJAGWlt11HUpU3
hxPzglEHUxT8gR/RE2YTS1wo4qEmZ17VR3z0kLhK414uNecAD92zUQ7isZd1nt/j
EY6zz/iy03GNAmHIzlA1NXzCA4JqmpCdmiokStQQaL3jnpmtmNtSyprsEYCYlb+R
ZI3mqYHggTeuijjo38rxTZoLB0hVQxRZSXGotiQf+dS01Rz+uj4zGGYvvjjzW2Dc
qOYExJgPRXQYer88WCMNOX7hYVN4xo5Vh0xsNJ6C/fKJA4P470KNkUUB3jeTvZgM
C3/KOer0Rf8eDm02RcQRQICBCHRCLiD7ObdmSj4QG6hNFxcyfSpfJHMDAbZaj08L
gSJeTO/Ca7h4MqvHubqSopSjp6LNdHgFpGzNIm88sIOXzq+aijNvXd7iyb3cVKkH
FC+r2LEAJp1nwMTHr8nHfAHY6V0sMekiJc/QGH9uiKKSURLPXKM7kOtAsUAoZ7uO
YQgbtPhEa+7YcYDcuuU2+LdkQWdYSIrBdQK6Kw3jui42UpzNcA4L4ll9TFDSFHAR
Vd34yZIHljfHQciGSQ5WTfJQKCx7c0vY9HqgptgvSW51kP44piOJLRk/Hh43tzlv
wSAPbfXPm5IvsC9eKKSFeDcKEcyHe+6XWWqLmBsC4VaqEjpA18lOaXWsr4c2g5KM
FwZSzCF75v7THmfs3jSrtvzOopJuEdJUFhdnRFVP1Ut+IF6K4VHGIam4Dgwpaczz
ltgGzjVF+oI6SOas8WPdZG2eamnBAuLYH6CrwhM9ZcUGO5dms+ahAn/dD9Um9TCJ
GB93nnJnBcAZRd5gDN/0tiSRz+NRQ6QQ1doUtVxAe1Vmi/zYD8bfYLZOyA9qofAQ
FK4XerT9FE6FrOKo9C04M0Oh4e8ner5NxbcIHLm/LZ3uUStdq9ZLC/OmBHhMNY9k
TanzGXiarIaWRZlicKoDevAGuI88lLACexQPwlEuW4uqcPLohV62GB5mc9XBFtaN
V7hdL6OYTWBl/1k4QCq8Vsr3V1jLRowHRMgEYCBdsY1xnytsVMwFsH7lDmNYFBOr
p5pGcbnPApN99lUgQvAEitkc/vxJV3pvX3lZ3q2TgsKXgTFDmDXggMIhFpNW/+P1
Un4g3B7RZg1G0xL2hnt6OW2IEU0DG+BAn5r3ruOlZpCLLG+m4w2E61viCw1uDTBF
Ol3jURStBP2rahKuHusjiFZTme1hNkFSB5Cas7+S9DR0Yt37wvV09DYTPMrMsJjk
j1iUsXppGPzC5R5+BCq5zWeXID5SbEgDyfNBgex4YTEhSvEPltiZbF4470igIBSG
KwKlTzCD/4oRlyeVjdpMFhYHJwnzkNl+OQ1OhVvGnWgSmX3C8aXe6zyDi8ntyJOk
bt3AKf3duDCi7DxtdoOCFFqffa7zJBlZNi1Zgd2GP265o6sKM8UAB3SP6Q6ew6Yk
92qPsK4vLVacElAJ7an+Awl8LJ3fHF6gAjY3A2vfkcTNXMoPsk66Os8FBrjq6Sug
9IOJQz3vzXjOwn5iK1IvWZkB3I656k+pyE7mSgaFpcZT1QzMGz9J/eRpdwxO/I/0
xg76rbI5mC3kj8d+42EPE0d+nOHbx0pGUyvcQIhIUwhfKaFhXY8kecJxCxuU2EWl
8pdBUIYXyxEmW6VVO7Q12WNKVn1vESJia2CFBT0UGNO42SfCWWvHgcSpF2Jnczqj
jQiDUVRgbBBodekYcsZKTS//YAFiLtKkVtOP6HKLSHido2M2Yvu7x1MCeGKXi8Id
plFuQgBMMWrbK5mAjX8a+g9OdG+mJ1yyYHe1QmoXZ/j380onJZP5Y23WcKIkXu38
mkTjcZEwWSrvt58CbfyGFhBVpih7O9QmadEdl6LVhOubQHBQb3jRL8AG1tnAIX4D
KEME5Rsy5EC/5n3eaIFZJWEZLgvkYuQ9Dsz8etbYwNmPd9/hRcPpwQ/bFLX1uuAb
u8XnkDNCw4nzuBEBsqG3Alcn6KlAAzChCPZDp8cEfC0Ad5unTYchnC3LTJ9ULqVC
sMfkmwd5n/bOr9OI1rZPoByief7p6+yDcsFsGn37AjWFoV5xvO6HouImB2WHphKU
NDFJhbzhy95ubfS+0vAvv499yUAFkxV1GMWL+JV4UDIxrBcOa4MDHzcCm6sp9Ihh
EyJxMAGJM0ShVjCkBFCvVnwX1a20Wd3lssmSxpVEpnUXBddbXwV8G0GSD1m2T/86
PeBiPpLFFdz3hBilpyI96gxQh8W/F6DCunUjVAwECAk4mqzYFbKfBdMbF5juiqCu
vxkmoZ2A2833kIn6zz+JDJFMcekfrhNl6ZxwmrT2xmlG0+C1V2ZM70lXhKirk6W2
ZIyXxz0UKDCb2THFIoslloR5OAPHi84irph7Y3BgwWq+vc1kdfxgNzLTdmHk8DcK
ThGQKPJxUhRSQkdLRVE10LfqqVmaWq6dBbeJLJH+pxuERYjFY/7pegBW5X4qVf+V
c1SD/HPFGnbaUHTzYmTOdYy2PEmVR5NIq4ADNo+SVaQlD28HY3wBPEGcrQNzjhiO
D5QFm9H5cu3yK/MRNA9c+3QkExgYZ7AXu9/4337oCCuBj6+3QC6/XZH3AKmJe6ee
2az4gJTA702plvmQkuiD5juJPD0FHBPSv4yTc0Za0OXiiyVWuAxkKW6n1aCR9dbe
Qr7uzNVveETswutbR60+r0MJaz17u9AqkHnG0YwnfgVZ9S2OvZJXFcBBN/r6zaIn
dClg67fQvgs6GY0ZVQnQOwVu/yTp5wzQMfHUuUG+H5MSM/bL6+QjvCasmv8hPjL8
29zkxQluGdHJB39q75FvlrMAxW2sQEcipaM6ryOOgXkN5aszIHNGWnR+vH7Kjhbf
cUL/7FDp+tFE83MMauzZ1JPTygOi2MJdjy9aazWMCNFAWsbhl6Tr3mRsisK7SF9p
6n2NMhzWzGopaVOLYs9B2mjCvBefyZ9ZwkY4WttIzCH/PXuAeIwAIdLgSO3WQksI
aPr7k5/eHlokCpPYHfqFUQHDBn8khQ5yYuiUVrQF/gXpWFxJpI1fftSfKTyhPfVK
VAptb4/4o4nDXEL2NZ3UDGTyIbJSmHFhkModj4ezBrGRFEDYSrUOPgk/3l58YjZX
TEpiYYRGwweR6EBXj/sDlpgWDFY9OnoCVO8Wzxt853okO3XGGj5mgtXFX9uRSbuv
9AJFwMdmlKDq+cTOYSd/8J4u2XYXmkAOIYLENMn8fHgxZP8eS6Yjf+1GmggGS9Nj
0DUCNcO+otl9rpMGbDzBqlwRwWlXP1eaZfcEZ4w/mEWDAW8lo6kllyvJ9YrmqYsk
ZrNCfWZIRXholvGso9OxYjhm93Po+/D3ADUaD+R8g827E8JD+WJhXQwSehLCf46C
0k/Dj5RnjWkx1RBsTE2v0a64WrkXqf3tD/i07I+MWKH/Czh0yuBBogdAM+QEsqev
IV+UJ9qoflAxKqSc1GquBb2cc18SLbXsxpxvzx8iEkc+iIgioo4tanK/aeflXUSh
f9Hj1ikPg2CwfQrf6vOv6feeHhjcJqrT4qHEO97vLDbxy5oT7TFmTHhbhcTnjml9
6fzCVbnU5BnrZnrr4LrWE+pyakwULK9aWpof7QfFrApijh+yl9iWfplmp7boj6Ww
hek++MTej6v3+gWqlpMkOj5V7wPFIb/+mQHVsqdRoL/GedI3Q5Q716J0yzvfg3Ie
LnuGjZ7ajE7ZRINTan8j1AcO852ZBDc34I8gD4+UNCLAZr+XXKQI0vrrKf95rYbC
E/oFCjpc1aDUxQEObRGvGbDtLCpRYO02B/tyHUB1WEf7Clg0m9kPdGU1LZlqTqag
gdbNm9vD+3rk/jovzbEN6YkvBxCwz99OyLDKKt2N6hv5zl6aJ/4hsPUhYa53Sgs8
zitOWJU0n3586oqgVx1XjT33UUjkrJe9YcBzOlN7DSovCUPl0hZRrsk3vHFfJf/d
zXeh0urOhmbWRAol88wQ0CJFDCTltJ2VPryzZLIWwycUFzLcIUj93S1v07amXNET
Uh3OfPQTYx11lCrNIvWqBNnZOYoi55LOXpPVl0rDpKS7cHnsgmEiIKbjfLmmlyP7
iAFYLON9AZBQ4qiMz/OxUuyoEiXLuZXOQKFFUcd1+4V8hdlgN4Pb6CHsYjS+KH6i
jEsxuDhPa61aFoAa67c2rBVJO6y3q2eNe2jEmJuAq6mLRLgxCIaXKerd1TZCYKbj
MvMxSytxdGD9ZDAjvj+l74Z7pmbQi1+HTTSA3JYCNa6NRYH64z7XSZ/fI+9x/OXW
LHp66xpjsVt+8A53XG/c1UB3Et2DwvwzlIACpHebcXPoNux5kz+O0mNqHHWlFS0f
L8nsXdWooTI+OJfsFOSwsH4/0f1OfB/82TQ4jRoT15r1Uw5aRuso4M/GBfsz+IWB
B9qhFswyRF+hgvPUP8S1cW2fpZDt1CAzJpIKz8kos/I7GF0f7pwIvHqal+JLWs6M
81EMZb3DBDkGPVrVTVdfGNlviL/6GiptL/a2YzjQ6yaz54DXi6MzEUNs9tMPKUT2
tJDRhuO8q/pDO6exPFxOjutAyxHDp2MtLSMGsfOgLJE5Sr6ww+52R7QfgUOlYKnu
wKdu4Seyk1cifbCaMmf9yew++t1JvIIstj+qYMi74QsxDhQzGF79mlTAfoLXXXgd
mnh0uGkUZyvDFqH8FxVbhKg6OlKC0ftGaxQ+aWcYAJIll/vCOSiwmAhNXrbJF3fS
YD+NO7QApbx4/xPG1G802HkSyeyjLQt0oH0vUhOCTM3I4Y5EL6rEmV21RVh7vWIX
qPBpK59x7WEiedQUuuwEZJjAfqolBSejRpkOGZsX52LB0j1vSanE+RvNrltmK+HA
WI/jY6s/uvu5lHamgrYuSuefqwmze4vKUiIONXtd1L8tugyXrIarjrJ6/17cg3oZ
pJ4NhQj9wigDl0U8MuVJ3lReotWRoW1mQYrceVguXrbjSzCntDLqBU3gVoEOmsHz
K0gsdsn2QJWh0VY1ZMwqd6S6PhvQ837788+TtatlnaFhzJybABKwPslXOEv91w8t
M2z4Mu3/70A3M+BVhffv3fMOun4k1t0G+NPx8aiQWvXpZw+Zj+06jvIRIot4IeiI
yXRU2klOkJW3dH2TyDdPEeV1QQvDc6eSoY8RiE1APixOvIXYBT+ugTCdLUY23Sqj
qzp2hKDlmbgEawF/fRf+SckqAlvjivPFszIGOf3FXrBTiupQn7xou1j+380ialOP
av/ozfQT2Rjen6QqxeTfEx4SHGc877u1Lh891L/rSgYvHzcaOtTpHBqtSOCyPPzO
opzYLTRpAcx5CzPSAzZC80C/mxUJQC/qmIyx7MlNojyVEnK89lFJImcRqR5/yydZ
R7WcMoI6QhNO+GJDjXF+PcZ2EvxLTTLJBJGycKhkYW40OGbH7SEQ5LCpOWQEG17i
99I533wkMVzFWzTY7WFXnQWHLKZbziMJW0XpKOhbTBXJBUd6cFor++2+YpwZlvFb
Cjj1C4hdVhk882QCNotO1k4B43pyEJOgYsxZhuu5GDXxl6yMOB7RD42LKzKxSbg6
PaBQt3nAm1QdMaK6NoSqt6X9rNzjnXCVZke0fF6rFrm/MrHoSFicFnsDNYDJoYkW
2giAaq9gcxJc36f9gMTeUTTIq4LfBANTmAkKsBnGbsMmuXAQt0fcr8G34oT9YQPL
q8gop4FkcCbGi/aCvju51zJF8AwzCuJ7It6xaOw/N5lfjmLH3CJBKOF8afqsd43D
8Tjmr0WVfsupMhd78ilGCpglx2W5heFea+7CLbmiEBsgZSBr/DiNLCI+8PpMhw6B
kGFQApI8HJhfr2Qe6h8YDozjCLmO9SBdPIGM3g+9aqWio5FQBDyOuKGH4AHBML8M
a9jgUflVtJY52X6u31n9yoa0K5M2n+SUGGNg7BCa2jWlWpP4jkAiNEAecZwJJpXO
lEicdxy4z56hJOGMjgZW0LWRWE5DIMLtc6YDFIm1ACsxHqYkOkapBU1tIasAw/Zk
4CjqfdNVuwVkN4A04PmI7IdSNGssG8U884AyXGMMxoV8unVhmt+lghXHbQb4VXfN
3XxO3Si3pwEy04Mw0U0NENkrYNM9hEwQll45VZtkyM/tXqI35p4gqOqtEyHc3UFx
x4XJRcKfPMUfIQp83l7RhNLpS821mM7MZnv3gZ4PCxVUbEjlmhKeBkXJXfAbCfwJ
p3hfCVKJtZj5HMHB1Ex/6PrGeKhXDF/460HNAbGeFdPL0j3/9hfD6BY22TMYsfiw
DP4mi4oAvuZRHyIB2k4VM8fjwLBQtfsrC2PQq5OnEaxnkeK+hv70jWhfcpYdkBgP
b6F2SWHNNPLdD3zqkeQxTVD2ZNWqxOyN2x4MHjCRu8CxurEcXdqogCLAgOWbt9Vw
4wOwB1PnhuuhH7SO9R4KFFhPLx7EKDG/XLoq79WvIDItCNSJYBD3/A9UQ+9ZBRtc
ncJydZD0JmkLDTZytEsmSZp3Djwkha4/GZyq/P/S6Umj6/ErwJV3IvD35U4fFQue
hZ5RKx3IXW+YG7lgs/+8/ext8dJiy2R9Fj4/8T5oYOqkVf3tkvc46Z3NOCG47EAe
8KIDWMoudppt166oehR7y1NRcfXpMYGfnC2s/siziDD/8/IGtQehnYgwKlt9ghIs
uL8/JbTfv6oFfCP2wdJ1/8cnUOjpplrXynY2vAkcWilWTmJ0mjIS7OJaiFHPM8lp
j58ld11CkSvGAo6ANUKPX8X4GtNkEFvFpMLrfUGtCjJn3UKOb3DhbwejD3rYifHR
63jlb17BShC03KCigUvyHwZUc/JXYcRYNO3wzlufgMOUZOCmnb/ky0aca21Oqv0c
8NVKAA0/3IXc3LDR3jpip+t1nGH1EWP2IImRJPf4BWWYVIE3A7Oqqv3/TGkY32OB
kXQ8QuQFSMNnXSo+CdaysHyejsniuTaHl0Jf9Fi7YGLhxVhKIGzV+kf9RF2YCC5a
aj4bBta6hT5toaKYAjYL8l7YJcj5Edb5d4wTPntoMxSYRj64eL6NcXExTrbbEzIQ
BRufRbXOS8uPVlLrh43twY8UaluJ/yLgrqKpwcX8rb4ity/cAT0Apa6WlN3P+ToI
588K7SxUaVX9kGyH4K+zOmj2OA+b2/0n0Slnjoq5hiximqVeD3cChTn9Sp5QGIuQ
EgP915TKVWRPcQfBxW5gcS3PWRH9bRs6ccZpbgL47/IGbyaMD2uVnQqT5Qo/DM+Q
O2lnH67aIQpaSVVHfXAtoO+/mlOgMEbPRg0p7sqARvkE+zChoTUMF7RWTsCV3xob
q9CHths3K5j6sUOL424d1nw6D880T84LKbn0VF9lBr5YqJthX5xctJgcyj9AC4rI
nO67EXlM9ggLcyax0gSfzw4rNbyPPHhBOetPd+JZMd7BEpaLOnkDctWoTSYT+Rlr
c9X0W6WpbdWLysN29q1JL954kmwL7sLmh0QTdtMikJFuULvCBdt/APKx5SXtfDDO
NrrifMCEM8aFIR/FcsfVs4V303Nw2WgQkCyB8JtvRNSlkVp6luumkVoutzD0XNF1
YSUskc3INptPGxRfAHOgvPTJ1O/g7y7wOePUJncHQuTnnUQtSWMYzr79lHMMTX/+
8LZEahTTe1qVoLZ1Bm/xssDjQDMIg9IBUMQGyGvXYriITEvwrTIBOdELWrz67Ryo
HPdrINssvfdLUfhvzMCv6dz5UT03oGfgAH328+1TBwiL7p+NMQrHo0hDGNEU9NH5
uh1yaMjFf9df1lEORlnRlSfHNhq4Xd24ybzAcHEywmhCA/FaTwsGRsLOsKnKl30x
NpBhe4NGplbUbLf26Hv34foYxr2aFjmDOo7hmg5rjSfeHs1qA1m+brlW8hqhlUBI
ldZORFHzWNHmcYHYGevtzZZD3o142bslzpAb5XPySeomkQ2rId/eZuDhHUQIjDYS
cjtWZrwEeljmXRzr/Im5uJbTtVEpNwVsuNKMFdZygQ2YX0Ua7D8vVpUli0WcgjJS
ym6TC5wDx2hXmotwuYDgur0GWZSCNYdoYD9RFcuoSIXcweVED3iNhnzWql09IABd
pGgylhFhbdpd1RCJCefI8AfBOi/8JRWA95xns4QFxIbwAaAf2EjHjB2zgHD1yHxd
+EYb6ypEkURQ/Vt17p3OaGuXrhaPtkZOCUBT+1MwD1quOdGX8VKOmTVyx2KSa3JC
yyTs0N/Jca6bJIMqeJuGOBN7ie+Dj6/QoamIjYfPQcAsAR0UW5c8+tPQ6OXKFXc8
7f5wGFYhFmTd45lStmp0VDRxGh4isg4nYd2SuaaEOt/dVJF5xQWlKFhV/O55PpMZ
07QjYcWe00FQSIx70uIDnZzO1SJu3tc4+JtyziC3QDBWgAXIjfpcRXJKKE/JoGzW
35q1sC5Dp8rZgBC4wMgcTX8mfpvf1E8uvG7OmQoIspeKT1l8dCHzbMopJYZUzAEH
dfPCfKq6/9KEF+QgLsVKNoQuskf6Cdh1nO430XF5dtrX8rbdNsGOi1elnaIBgpvN
b1SiS5Ot7AIeNDONcyw6s6/DTr8AIKnXnoC0ER4nSagU9/KLR7Jup/ojkbJn/zAA
nyTz7Ymw6w856sr9C7ymSVHkWKIqVtVT5/nnTk0HUQwP565YIgf8Q0fnXjeNj3Nv
ntvSvhbQsYLXN5sO9E2xvdQxULDmnuYiEPQwVRvSoOFJq9AZtzqQ9+dJBnFMYFNU
v5za+hoSPSobZx6BZo30PFiDTkl+qzpf5rQDT6wEvBJHYg+AB6ohOAK1ntAAXIzu
iqEmyTppMBc1a3N12knIzUT2v/81SqAM3rb2VBC3opwQEmlGLHVGMDNm7fw9ZEoT
u2x+oVidlid3CI8jHu/zdYzQVq4KouamnUHmVRhBaKCX9LBLQHV8on8DZPmZjE+x
wJ/LEDM/FAtK5Y2me9e/BG/Xj8HkPmCsMDN8uVg3b7QLQVnkCJ1n1cwqi7YEk1Sp
7avMcpOAkBcd//W039mDsZaIQjJ8zlcjZCmt45xXYQEu4Vyoz64zk/ooBY2dMqo9
Qi+3KG0tD++8SzzvAFAZJiJ77iFceZbEVgWsPsztD2KnE8P3bxI5pdnO3A7qaVN8
+8VTfmB+bVgSAYIcxCXKxg/9gDc/g6QHt+7h/8V80f12JV74l4I4z4WlDxxY1lL/
oFvDIWwAb3ibBGvRSJTrbpGDD3CtGIxXmEMYA6dh57kM9mjqUoZm301c3NfxzAFl
FcDOjxG+DyuA/1OOGRNVdKEfFkQAJ9G8ALki4H2WioZV4ePlebXXEShkzesjsCRi
YEGxk+JHabM9ZL1Q1jh7PkAQOiLuQQ9EsOCgcn0YjX5dO52295WYBDY0dtVZml4k
bGJfHhar8Z16McT98SN+Fikeb1UE/Znw5i5+s0jJU9RPmfVm3ITdVqcsKyEcP+oA
KSR1lhzccb3f53WF4oQOq6FtP9S+IHbx5DiapY1nZPINCsnP1U8MKgLQ/II/t///
OZPiKqZ9smrqeBMtyNtk1oz8+AZuboJ0PdMkqZF/hcJS5I/psXkHN0zIeGHusbUy
5Ed73BZuWC0WCC8hrKP2ikVqNjTSe8F3rC8yWJgxtbT7JYzt548UnGpuwgaaoTVN
q44SevCGQdZEhXM5FjcEoYGM4bDSfgiLaIMQCk6RnKJFyQS4KxW+FpI9c/2r7HKC
igEH41XiQOzk8Nnzr1LwpJv7f8Q2ug2wrYLtdl0I3lmfpPTewRhvUU1bct3g4yXv
4AeDuFO4rJsy+/DonbIVNkHwYiDTGkRAaxlIqoRGCnJxGj+hvcP9ePSrk8OFWR+n
jQj2YMJxZoaC9W74E67pErOmKROrg8UykOjqqa0j2gd2ZRIG0yGBdZpOVa/eix62
zpOOQBJZ5i/GqT/bRIYXW5TE9A8heRi6+0LlUBtNL2vKPULDj/tq8I3qtTLX+Rwm
9uVOGbzToX4D0N1PAklxY7JO0qHbKTvT7YJFKh29+/dW3Bw+2LcNnMEaUceVlRp5
momDYwoelHmuGvzKwK8zSltGLKunJFSYWT2hOHW9l428oNeJidRaG79FZs3YCNPm
QPqeiMQFLvMJL5jD9RdhwQkUlMd5od1JLb7LiH+HO5GpESpYWho6RDsWHBX34jA2
q57lPQoN+zTSy7SDbRO9K5WM0F4TV145eH2Edlfd28eO00UNfosKsHdKflAKfAg4
MFLRmCcTq04GhYolK5MdFNfhmJAuK/n5Tp26dhQ3HrBb3WpyyYYL26eCUOkFQuUd
f+cKBpwozn9y2UeaIbKLrqFGrE1k7bQrPEMeg28Du/hXbrLi15Malhi+Atm1MFW8
Q/AlNz6dw1iYOzmpcqc4aK7Zg6Jqso2eMOsClq8MItJ2ne6D+4hkTBXbNdXJJDVx
Hmp748mjoxeXXwsDY8+T3LQUTzqFdPmrvw2EvhZGO9YfZf7FOsaSCzBgGT7LQMJt
avkURTHKiMHuzxg4f+mOh8NjpyAhbrrvMg0Oge88Lp9vSA3I8g9Edpl0yn8DSRs4
zLy0RgWUDezdfOj7PNga2VYOhrbORqXYlXB2HnOOzPSv11lMAH45hym05qev1UPu
uAsM6RNs7QB57c57MY/dmAhdRv59YZH5LWzPk5pxDXHIQvKKFbwwkh0cLUzia/Ta
G2MIWh8anj2ihCwWnc7Sjozl44FBx506cHEi2tVM6A6x6JhuoCa73ggxEpAeZOVN
zWMt9alc6wHo5whnOhGRb0TqFBQ0GAHpRc7uY1gtbj1ZY1QlMEmBla6CAWnJo9P+
//+dIvRSg4pvU1STLsveFPX+2VA2lHrzhmZWONamr7Q6BNQCT5FY17OALqw82c7R
xdmCfyms7/QC6Q7/Xu3hHe/Q91Ji69Hn87z8Baz13lXpJNu9QGLtNa+1/q1l51Ab
4MLBRVGkAzI29VPTDKkogqJbCTqKkxnB/FSGLbI0OnMfe1oU603ydPCTmYw53zbB
Wr89f5iYF8+ANDHxAXJQEKZinzfVyx0YeeFn76+zkLWOXnP/8nTQs3R90YQr1xbm
9DA7j0nnsq2jVSJRNZ5E6/4CkRh/J+EOb0uOMjSHnVA1vQK2ekP+aKL/pdOmREGL
yKK1KQ1NbBdlTNgzYT9eeHHL/v0WaPw5nhvb79KuNVGpTvqDEHnDy+o/eEX5CS+G
3E2ltmqBH9dXyXAje89NzyfbZf/63ylFCBnMLDfpEl9qah8ye31lxxGnQfoHRGpH
JwBeU+HYl2dletYqx2nvmfW7viumYQ/QG9vsjxjKwx5KTjDXU34Sqfty/ugtxraV
eT3UaQ2+eje8qTrMeh8I5YSfaQTl72j/2yuxzPrZdgVd3sCIM661o6j2dGq8fSCr
k7fqPGHDbXK6rzT9E3UQ/h5+69RhUpzzJnFEDuBGV/H3ERZl13aXlNyxJ+TdKI4k
fNW5Wu2WmxeStLxEYXNVpB986OYp+BMeSa7sKrVF0Uj4UyGVRJYGYBz57l7oAlJZ
3AlCQ1BGpI6gbP8RJAp8jss91p6JaMpnqyXbqT+4MoD2SAxY7YrXH6i82pBpdcWa
XNl9ly/qeEYzcboP9IhBF4dWHtABVX+HthihIF3Otu5wBoW7e4TRpc56xwiha/6L
ijNUOY2f+c2eKwsPSI2WnUJjTTGiUyCkhgfnNgErEWFKY0jOgYKg7thCbxf2CLgE
hPneACyXNAMhLM9Fkz+SiUtRWg1ktck8Ggc3grnOnCbn+U99fPvdqD9I61ZJS4pR
De+4b0QL5B55HNmHd9E874+Q7b2bib4DNp4Q2Ic1dMM0RYYZx/P9Fvr9qe9uk2dZ
1CEX8ZuCqrPHn1FPHhbrNSMFjNZ8er2UwxHvLMIupVNTKHNRBRFDxtlC49qMuA/7
cvnKqalVpmlncCzCpc/YlFJfVAc4B8U5DlWv/lQUFHW6ys/XK9l2QQGT/lV+36Xv
v2Xz9eA+5Ql3P/K0r4xeSH8RxQtCrshKe+C15DcnrcpZfcCyKGtQ4hsOydTJLPhB
jPIUZfoYo2wmwOTDm1kTxuoCOqUuGaAjaBcR3rqMp7q7chg7/TYz/BuQFV3mNo9g
9QYkizfhUL9VCGGcqFHS4ffrfrb48Y/NoBxlrDp/rnj+I2ScjCztjWJy5HshiyiC
9ByOtEvXuQ3tt77+nuWs6eEXkmXI+1WwROzigB5jEyo1DrhP8E3MEEm6YGdM+l2O
LALwtu8ayuLDH5veVSnfDeSD7c+w50CyXApIJh94qsGSYhEB652ze6GKM+wiEv1h
awBciock+DfOvz66raR0fh0YBZ/WCp3ofv8Y2IfGgcOBWkaPsk67i+tbp9QTKgDW
6JcWEEn7GpZsY1oPnjQxSgzaBGc97v/Au8bz3H4vfKqRkyKdob+39poaWuViuJgd
5nUO/doynrKr3cUdXY077Q4uHq/xte1goQQ29r+ATzLpCJvLFFYcKkdHi1BMi+f7
GBK1eONFLe0Nvzq/3LPK+vh8Zsd5KZcz7e+0fqrBYe+CHqbUC4BkUBqA4b43VCo3
OimOUlm1Gt0bSgBWpbB3qhKYnQXa9LxXKdOfGzHX/+nx37FUmCjz7pvnUz4RA8Lj
8gLnLfT4vMS8mB71s8P5k+z2v97mj7nW+XB68U728imfGc1DmisNz4Kkqn7aG5hc
Z3zuxNwHWmbopEvN9TekRgUZ5dCSUQDkbExPJG/rqcWWX5KJf+D+ssM189ScE4Kv
wMv+t/1+9Hxy0NRgf1agaq8S1OvrhHgfRAT719HStJSiLh9Vo0VSH5kkJtK2nlL6
07GLHB0jRyuYCQ0jHLHb+eFp/99l1dkFioYmZ+FAMqfz5AfizaM4kGbHCh+slWL2
gYZzN7wn1UOfLUx3L91yuLIzPvcZGJ2d91RPYdBaocuxZ7lWSwHrnz46MmC/yalx
BNi4XwOeZ+y2aH52GtVU0I1/ujMI0CKbCTfuvCMQUuNvoxdk9i4Ka2/Fek7wEtFG
khFQw3qy0tMeH76c/pDVlYDq08wWZwYMDrisKN4Ol4IF9nKgxNWCgjAaxEEnrIgh
EwN6XBLIWYNmi58ei+55itptFxEsOg1JSdjPQrmfqNxMeGoU4CwfbGIiCHeJtsmj
WFkhRVVK4x+LksQpZ3SQ+85YqA8drcIcduEm20NY5VOvZFJr3iJXm6bMiBM0GGo4
n949wtmDLUlNOiv2+A27yZB69zLW6k0lvX9qgs/yR1tpq1wE6U66QU5+q4Dh2bIf
THt5z6QGXPC4PCl4LJZcFdl3cnpk/Oi6iUZtK0ty2iYVRYyo4cJfwcaKwffeq2nD
HCTHdnMoFm7TQjDBj8cNRtlbTRcu7zAAJPW71qlT6NkK17GXRrM3WJ+0nNg2us7v
c5/uNAZhYUtcW9wMBZcTK0tI1WYZu/CZDcR9q5Jc1JycvvJ8TY5vyR+iydwV7T6w
kCrKKia47aIs4Brcad9EFXH/iEBjg6tTvfvfpiw7aIoNwel3dlh/cOYh5EjwEnTm
j2hmNGB+KkDWZuVrnBnIcMzLV6c/jyHmLje2FCobSBAIQyO7oQ3nxQNXe5jbGVqV
fuOTg/He/vPsKaZjGVsRlx9fEXljd5p/nkPDHcpOCA81LF5xhnzOuHHolWt19PAb
vELkxJsslDeHAeNuLSQddlwVo6F9Ym0b+slLzZmxcC8q+6yAp0QpYOd6o6YNVTu5
MUUouOsz6XWyp3oEcl33F5yEeRVGPiGJWJ7gRWq8SMEHc9Tvg/R2LIkbsf9aLcSi
yB+OmmIbVnphkwntFVlxwv6om+hUi2mWaals4MdpABwKP6hxjSG+WcHdT9fV0EAA
QmdziUXsdEPClKP3o8dY0YdNZ6v4V2JSXobPQ+feIMbts31B4r4Q0+KpZ2+6mf6M
8FNfpn17Mq6K4Gjm6WPN5pyGJu0r/4XSUDZBooiHTStfPdi5ZxhHDIllzX9hBxnX
/kQwZKO+wHR2uQ+iaTeHyHtGY16+JWBblgu+s37AJZYkjVHDYFYqFosJca7ruIXp
y6NBpaMdJR/AWtN7LSsTe0D1ctW8Qjz8pDRD7C3M7w0g4kYTWJ/qBjgNAhSOlcxS
KfcQUiiR8v+riEc1GiN9owAbNHI/qECpaNeleCCPQbN2RCw3Biol4nle2NxkomEM
V1+dm2kTmk2v8H9Tje2zHJN7CjnuYnsNhGX6Kp7bgTLAu9gp7v02rYVOlYpehUn8
hEAjnF+dltllohljFuRgQC/C6cUDB4Fz2JVxYRiJU6JTJS+jmvXkVEeaR009GvWK
sLdY7zHqB3WgeIY+8Z9qzVSBbI9soMFq2HBnA33B+Ic4qnf0CvqHawRIU5dZ9XEG
W8KFLUPH9izm6AZwyTwLB3Wm/W6TpNQUgh30YzIRkn2S1CYOiPhOYadL4IEXV2p1
lfN4pZnEowsXdnMVl5MDN/q8hgVOW3MXn0R6Cv5qMfPHNb0eVjnLMZHVHZVUAh0f
RWVkWyZVCSwwjOIvSBMVK6gkqba8W8zRL70AfvBRWbbaC49KL9IOFmfuyeDM2jyn
NNPrK48t0zrnqHoYhLWNf5ZXxEbjDkHhiGYM+j+5+3xqFrk/Dng2Xf5pQ6wIScA6
P+/aKTXftVbfmksCnsrwRGYhpqyzY7j6saeu1ZGzlVEziXJKWi8IiBbsdvGF+/L3
00JiRIYqhhaQJk2cQX5aHVJ4Wodpxy+O5vPvFarnDhj+FDZ86byptceaPj5gy+dv
h6kSAxOOn3v/Lc9LpP7VPNcmlvjY+3WP299Ydb4IVWOOuSX8I46izt8Kdhdmk1xs
VHM6+jYzPbcGM98ACWNUABwlPEp4+jO1Qs0Dk9+4blGVxZH+zlH++w245PFkS1lK
n6UF9DP1JENih4Q6R56Vsx0UcyPpxiWM3LLDslPBphrot07UNcjmdgxsUWR97Oak
dWIoGuKT2b+A7iVhbQMS5T7zBx48Mq8GBWJA0A36PxdZsxOO4bQ41xoFPIJtPUzC
WEAGehHDFW1W8mUBP3vUu4f7zb5QggeAgOshIHr62j+Tn81ELF6O6qIUXv8trAn2
/C9nqpPLMviot+99Vc9+5mcTCoFOSsK0VDerN1TnCph7BQ72dfNQNEhCp1+5nxCT
5ihCabXUIbocp1XuQpHoSc9CivCmGkOvMtZBBoKfv6dCkIfUl7bhUuy75DVjCF80
nQV/E/lqzON8nKOJU2ahP02EGM/QMMWhvz3DENfVdjvkrvuYcKssJk/Ui3LxpY6C
n+f4IcGo10CvP1mamXnv53uzC3tLA+oScw4vuDLZvkf9x5MXJeNLsPlCUjk1PPy2
oeTwkCrbJ5dkobxu9oS09TqD+gD9a3/7jjt3a3xWr6H17KXJ3eHbVBmfDlNcTIKh
FbW0yj2arJ79fdQBOGBbE+wj1ksJtEBvUk49xcKauQBYernEkzNe3hqGdswSWiV7
Bz8H9lV1Zj38pxzftwW2ar4vBvINvG+gXGlX/5mJXmdtQ14cUlh3oRXiJsnt2JBK
mDkVuqsRKN+fSTQNU7X7cBMuU8fzDElkfEQ+uFDV74yOofROMhoq8ql20thyh4je
MzLlSynbUbATKfe2djAyTBpxqmisJB2c/qsqbfF90JAmqaPZN4XXNOFG6U+1Aml8
d6HcfubZVvtxHwCwEsuvprMaE8XHLyCPIQkM66Nz3I9cPw4hu1T+zjokHP4GOxkt
nHkVjrSBSqDpRGBN/4ECLJpzRiAewVxskdw7e+gLeQrU8P5Rzl703eLgqHzNZxNz
/S0bBc7uyYiQz/KEfLkf2t6PpRvJp/qzEJHYhtAiMvJBKyoS2PbJD1WzWlpffz/w
QcbDdxkJug3H7219TOpHbpfQL911u78qpHacyW+Wr2si0nb0DkOsjMki3Kgj1bNe
qUwGNpu++IQiHTuHpRUNCuaHWxuLUMHmPhBhLFNjvZHTHY4WXIMJckDGz7ZRvT4i
nj7tsRqE4p2DuVUtqzUGa3uejQJ0qCYMQsz257NR+TOcsHvO+Ku3o+iumCZrhBEA
xcQQ69vFxbHPRwBiLeNorypvGLtiursYsljh5nuxL7pw4AW4lDvl3hKHKVbLofA0
t8UuEX7IlIV/cRkf5q1QxYfWqbtlwZAsF+Pm03dkGr1IxJufBXhV0RO0gBohonXc
BkJsa82ZHsUHPGTt1GPCY01JTjHlclx8Bey8t7VUTCukllnNWllOKdZBRFcp5866
Wu6oHfD4soOHryRSrcFH/moeIAwyr+ypJzmGVJNBELShlku9yRia01VCev49/xcP
meYHY2imJupnYTM4iHXxI9pZICFPxEKOVPD77oeI5klRuHEXdk3n3ctgCYvhIXwR
J7kerYsl17jyGswHbJe39u8q5SMHDm5F0c5JFQ67fBT7keo/M7EhakYcg/e2ZzWv
9KcrlCGndX6ylg3PUzhieo6MYJVqfFnvxDZ49PTcunw7Y0YrsYIjcFRJpAGRzWHI
jbdWh/nR2qnkD32oMW5bRZd6ZcnE/V6DdVDOX6Wuzn/gr+hU7x66NEgJrZBeK/NO
23wEV/Cy4tsg0w71q/tsQSC6VqPw7C9a9bO57w20lMIgzSYAqLBRKbpN9vpBShas
VrwRGstv1qilTzbnS+i2XXcfsVOEyNCZmHfapCsTPygpxH/DJCvu1JD0inY6XBd4
xSeSULsFanrwYeQ3Zx6JaT+PvzKuvzvsEWQg1nA8CeK5LKzsnAgXmcWpHjo3vZRS
DdXr+loFsc7Sw6ZBdb2LOspPuR/RvRwuxGjQvVuFNdgrpQKEUpZCoBmWAePenZM0
6R2VUI9Dr9uUnF8j9G7W+MpEeR97G3sBb0KXkn2FBgJwkQWLR6rHSkw9XkVkgFya
3iW8fwsTb22W8y2nP9fPM/BORdm7HTLI43GGb44IaEG1MnzyKY8gO24aVwPEvq+T
lWjO+r/e68YT2RfW+MnhvFuSFaXHj767tEYbDvSs6IDc71iBYnQoUMxU+C+56s42
/cgx5yq7f28ceQZaIrQFL2WD48J6Rke/s2ULHg8GXDdyr4G8b+xc8YxiB1WERmIX
PYvx2BwveJzySEf6Dw03HANqQKIdO/b+7zjZZyrubWW9ozVaQcKCzRPAP4wIvFF4
sG9Lt0SlHLLXSODAoAQUSBsn2Avp18iMhRH5eVOAk/qB2/6/hmf1dZ4Ezx13aGJe
eUA+EZyTT5R2W85cAUxpS3yaDaXpe9Umm+AvRw2uz44jGokhu9F4mhgKF8q2164L
Tb0vvMhjt6KieW6U+07MYfz1B497w2/hvOZ4u3kaEKlL3GH8s2emJZetRL3f/yCX
urFHgbgP4zjEOj1KREjSPnYc8vXiXa3PyPqHGKwqQevEzwD5uA1TVqQWiSmlM0I5
PKVv+Df/KthWpg1TJ9L6Jrh2IeXtSIMdR8jUENM4pIRzMivITYJ13iO6OwM114Id
So2Sn7FQ6HwRiSREIRDyF5xeqDhO+46Hc+VFC3N9KIN2vx/Miw6I2NPbGk8yNrRU
W2SNW77q+lWrp6l60XNwDXcUoe9z2r6U81aTFz317Tm+ZQX4RmWKFoRzBCVJD4CD
99X/9ZwV2McQX/XxvxvIeRd4dEUT3kLxUg1aK5EyKE48UJqetORdvRRsBVcYvqiW
+7eUS7Uxqsz8ju0R6NqiLfFuzD8m5t/cB6GpC1J7sB1b+Fzt3ce+65ZE2vrHkVpU
RlLeorOqy1zeb47BGQBSqUF1jeQXgEQ0rAs6pc7WRJ9JRpc8TStQsoWpEhI5n81z
QCFKgjpEWiC9dCEKl39XrBNjXUusxgFm2ACc4XWv8VYHVi8gyWrSeJG46CbvzNKE
3myo4s+dWsSrcoTsg1OR79eTv1hbA4rMft/EIo8S42B4h0Lf5el7amI+aurgQKJT
SidV2xUSjr+2WVSeOfkTifUuJL/OyZZlVDIq39gaolPYPFqytu/y4jG5SPKeas98
5+o98FmJo8QAXqaMlPpLVJGpJ1a2QkzRkleRl3g1mfA551TCWNWxRrY22Y2MWjdH
bik4Q0JW2qevtDUR1uw3CqsUvJ57x0J25ge4wepKuF0Mrq8GhUfD93xeQ55osaeR
L8w0jcjm/SLDytUJ8FiCKddZjJ1VyJ4xYWrzlckhxFBkbGjQtCVuw0sgDUHXGTsM
gonXTewxR7BJeNzhpRizj1nYHvfwrnKyV/evwDamUdAm8AuQ0dx1SdZyow5xwVRK
V0eApRTlBKVXMzLBCaFwLLno0CGNROzHLU90uNSa9jMI64bc3fwJZJ5/Z0jg6Es3
q4tifUSbz2OCo9zc1wHJQ3+MaOCEj//MMtuOYyFfLC7LFV8MHdIMSl56zmpQGQgT
W9M/3Ep00XKRAtJp4bjcehwe+AkMneDg3TEHFZb06D8b+LjgJjNzrai3tlLN5wUV
P+Vt4EUbeeefjTRvgugjHgFSG92vglV9tMdyuolrljOO7O8wqr8ZDDSqXxhaueRH
SqWRlwk2NDaw/neJ3Qbvb45/anlIFfSz66VeGIKfFjnXejb6fjscOdKzDtZgcA91
G6VYCagkcmZ6KIos6BYXy8JPGqP95J8ES0Ylj2nkLxjgtV8l5r6tgi2+WKo6mKoh
ZVWrtDMSiWTBGuU94Ef4PO7E722lHsEneSt1n3I6BXOSRYbxp1Nt9LF/A9v6Fa4r
0u5CJRUOqElkeMvCkEj8zAsK/kQJZI/gKBzgn+Wfuu84XjgQV8Chatgwr8UPE1ow
v6tiQi+zakw03cdNsKRPdPr5xvJAvV6HrH76Lv8hwnUzn9oOHneLI4P73Wq4wDpM
TJiOA/aHbTEIctUDOEhzNFQ1KQ38ky1AdH3pH4UBjVEEHgO4dZLhcblBmZQ28YaS
PpU2MLI1qcWVryw9fW/Ze6YtWtcUHEte7p2nPmexRePfusO7kMRO+BqDNbGLTrcT
2F8bUKGG7z6l5zYHwrREGO6fgIsGqBpvMrmIAcia00w5NuPxxqvCqzJqhr5UUV5f
PwZLdD/kN9G2hFv7wc2PSXFHZ7MZzCkfOW5rMwW/qleIFQ6NFEdUmU6cbG3mJS08
XlTfqmyEykAhGBuz4TFj1Usod201iWj3lr0IN59Vk6ZBiGUSN+JwC6Xx3XXiJO32
R3TRLWaBJeFnPvypm8YFw040jcqwOBBXGiHcAGbHJ+seWHG41/GgFk9ju0ZE4dsU
SkzlABFuQkCDLpWcaCfcIdfD2nyzruXEIbGYIYF8Tw753G1hnE2SbkSceyrXEnJC
YRzG9ZHQNW5y7oo9wYwYX9Rys4CMrjgBqN9H7UoFtjm6reQSTgXIEX4sE1TDSBS+
WLvmiLCKv0bjZpaNU2TLKgzWpJSZN737gFj6oos5NP2uyP9iGGFSBaH8MNwgYvmZ
w9x6ioB1wVxM71BkBMVC5Ru/pn+jkwOXkb5iGD1fVknmF5xiL1FBkh/lhoDey0Fm
ZHebOl35PxFRe2dQbvBDJw1wzSeE77CaktULYAbH1z6NK9cewH40dDdjToi60p3b
NI1jN6fyLL4pPJ0PuKAbI8gKM7u59q35moJmJnNtpzQev0xRWDFrSmDHo03O6OA8
vYyujcmqNVlZ6D/m3D4EO679o5Ik6HRTHgHH0+EAkUEkf0Y83PPR4DzRfQKN+QSb
Ei3ihBFqHeI2Cn6FnxOc13qfp8mWlGgcNAQztAc4drCxZVD5sIJZgrTiEhR/1c7R
wpioZyL23zppn7Zp12x3CB0ZnXaE5NmiiohLPiS2yvY8NuEC7mgAalQMBIFe20LD
uWgOmLss7So28QM43cXbNyJxHzkBMIE0BL/u5o58lltHLToVhyYIsqZKRnwRAA21
Ueimtc1aXVIQ3oBITmEpy7glGfBWblX+jBKUWKO1FAJ5xIAoGo/SIRdL1OLdRz6P
PwfcyIjnUzHp194ciaedu1z63wIsuu27qLjh9oujDs1nE2eaDnnl4buRVD2IK0Md
qfJYhz6Ar+kQtEzpJ2LiOu+CpKGxMaghUuCQaGvmFtdcJngHUzFHmI4tkXS1nWxU
vsKe5B37t7/pB/Ceaeln1pjOrWhkAwd8Hgkj/5VwG298J7SKiZKH+QEEBqhwhIkb
ydhqo5mBbU6rsnEWlNrYR6vmOmqiZjvMZJ6uVsfUdB72j/tmJqp+nhquHAZA4QjG
WqMryiW10XuuGSNX8CLrVGxouJTtBtWlnOFqaV66fMt5OFR9es8gU3dNpUw4tgHK
nJojGw1PhCD6k656Z72Tc6y+L6xzBgimWY7QhxdM7VuKHDAIhY2GoRe0fgjWX043
53iz7f23DTb5ADPlaJAKD8LE4q1P+Im/3oHy0JK/ZDikuYyMmCTGvclISvLgNrOe
wyKClwMfOysDM/U+pVYn5Ma9BTsA8vCL4ygA7dCnTy1tPIRYzRADRYI66vmiM6wo
t77ScBqpEZZFBbCkW48gmUOybxgN09zC7px0Tirtr3DTQcF0q8eeDCnYpSq3jVkU
K8eheF6DVWhfmcwkMuXrx/5sWBbjYrC7kdXCX+uqaMLoTPa3+v9bassF+cnWBs8a
tsdSxsJBr3s74mGlEmmsSQ23NOHbcsLvt1s+aileblhHU/eGNj33t8XAjQBo88L9
ojSxuX6JdXqpqxEwsyAWYYqnqR5OqKt81aYDM58yQNEAroFnpiiUOYdOBSfOtQM/
Hq+gDWcyaCrnahURRzrCavhEmlWHyRLXMTahQ8t/NTDxAdf0TFHvlWi6IvC5oZM5
Q3vaSKE3IjZEMvDEF0mZcVbRiqRAhBQmKvOlEOcCE/dGU3MhBWYmlt9SgnztFoaa
tO2RB+LiZZ8S2SiTJFppeKMyjvEB1qqtBObMhb0GxmzFbXzlqJ8hiyUHjVj7DITN
ZfuvJudyTc32RCMmwKbe2NseoLTtvvtnHUPBRr2MeGyajE5wvmEc0f4eh9fguFNn
EyBRSGE6DnOJezG8oUJzLG1bekQKSelJONmY14vjpcoWIfUDBw0MSXZF1rSsTYJI
mgSGDh+XPk5F650cL60ZHGoirw4lfcSpgUY6gRYVjfY1Kjhzophnb2NEWqw1V93a
eZcYLmxuDhcrbElZ+JhyxgQwwp6VmcAtUMIpMhl9i6OJryUfDjoq3BPIn0yAIask
PCLWdJju1TOd7Romlod9M1VXBzMRK2PGMH5Y+mU5B8Fzk1N+g5Iuu3zyPHXvgc/f
3IWPtCLpJzKvIPrQkek9bTFpjdDyba46ItUNN4vdKatZEWjCBpG2KXIFYFK6AGdd
3HInUcDC3ayZoBSO8gy2mbKYGkdYilac0ea0fl/4I9OtMfTjftCR6Icg45uHQ5Xm
DeDzppRod08ZJf9NmQjpx2VYtftO2kGXhaigHsu9B62DuAa3UscRDCg9FoyLZ//I
P/n5EfpyxrcGe11dh+N+ZCOQMUPofXEqrCsnfyr6Dj1cYKFjPvMZiie/ZaFOQR6w
9U+PyQtEzO1HcnPbGxRqdaVzRxBpXDdkZVfouTMVYPpsYaXYwN5v0PWEieKrAiZ1
wxexnFjY1qBjVJifyvssApXKLlzS0Pojk9/2dyIDXwm9kCVBy6KEUMThSzQN4x7z
SrG05YY46rUcCVfsnT0kdeewxpRKZCEllGOJ0li96zguiKTODdIO41A84coSG+pP
8yfCqm5RLyWVLkkqB+RBrsFnNtU8c81HNM3j3ddKkwbFyAp5TkMnla4xE1ZU+fnD
835hNQehB/uMWd0RE7OZLJX8MuKDEJOqw/y4FlPEYMne2Fvz5S4XkOcjfbDMlbUt
5vjhbGc995mxf9LTDkb1LvHqcoWv0Zn7k6zfW5MksN/QcwzZaK0YZGX8CMuZHnW9
mVoi5Nk5Jv74BdYUVVtB2DtPp/ocB8dvVHcAtRuKtT4gUQdgWD/QVsbRu9rOqM9O
ge6qZZnebZhb2YElslX5hgEb0NixFCyr1tMJjS8awEH3Zs/icSpzEZZVtALNqhm2
T3qCgtT5lRNbiqkpn2w98zFziDlC3l+T4isXe0SK8I1vS0jJrIJYwJdH/m2ZR6zO
1nPNiCSsck6j2CWDVHMKY2CeIDLj456r8OYk+T9W+Kw4zeZjI2FF+ADGVGJWQxhu
IzddbK6jcvzAR8FJCoJmrUjAYeVFBk/PSAWxXSAAZ6OYuMSW32NawwM7pkiigo3H
XhaN5rvpuKlcBGF9EZwUQh4DVn4llCjuaNQt7Il06uuAG1/daKmaFU0PUg023ZXc
EdX6/c1Oa8x3eO9jiBZPQ8dlqShZ/BlA7msNgzUgU85lxupdVIaJ8LL8cbZO/tGI
93vDGV6LCd/vpr9LhvYjPQ6ujQr0Lf5R2vuHRQcOnX3Cb2Q3QG3NyaIEHhI5kPyb
+H7cFYZJpgfMNh8gOv9vwHZNvtxvL/L2TWUZrds4ac5zXV9956I0mBhWAnn6qx9n
033wTQzkKy2ovxI6mIw0GPtgnoORVZmIwDRRYstoEeJCjNY4GEWTDFEcsqW7a+24
gQHb0ydd8tp0H784qrf2pP87/pZbHA79hQKJ9y8qmbOmBdeCBQrRMKdwGR+pINp6
WKl4HlTb5mZt/Qq6/mjCOTa+KDEp/yP+xKTPxiqjqD5t9Tq1v8OUGmTGjwFcpvIk
JezZ1SkA5gw+wTyBhlkmIfbm2mfdGZcVSa2VU1l/2ZP49VN7VgsA+ngh13xu9+1V
V3SrLdu/kd5HMjj3Ic0NGth8DueMaAPKvcE6lDQU/k9KJkotYXPR4n66Zm63VInv
VSLP8PED94CnyfVgqBb8xvbJJI9TA5ekS8khHuaNfSxgmWK348I6jSZzDyarqque
8azrMyYDKQj0AS0wNup3NQxvhb2Rajy5i7nk0ga4Pu3jQXTs6i5VQl28ATyrlMNA
+fN3b6aI7Chi9547lrnG3UlJLV09YJrQtexkJVKOQqtzUoGb47sZIQtgoXHCSmTC
E0T7i4YPqR37O9SH8OSOPPuQVVtYmSCnkuN/ih0F3MLZILOHGwkoc8ShuQkWJSl/
zExY1UlHzrUxh78sldOer1xMlbdL1w70Mjw9RReubfKkhaXqsmI02HrUM3/FBfPU
0O0XojqKMIVAz5ATzT4NO9gQPhc/Fk9CrEXgrLlCnWHfFZwVMuss4D7pGnQdcNjJ
ZNLZWgDVrj/QvAQ4SNfIfihyr+UM8vFpJajjPxJVXeBm3mupeDz7XtxJMTh2m9oE
iRHGleEzMvEAb9hYAtcxM9dQ9BvVADXWraZfBonnPmdZTql+e4OFhqPithKtkUXt
3QrXFh0eh3NMQLGHmrAXHbCppqxZh0zVsCbjnxCh5Z33Cpz37jvaBNKuAF/kpysx
38npm3RK87NgYTuZb7edE9C34Nbo5bdy6N4rh+DF/9K9icGor98KG84MVaHJRHZj
X9cp/Mk/jRLCVdg32YStsKPuHt2Cdq2L6E+CGOK1t2angCdkgJCNfGpExtTl9twg
XolacnZpXAPZrIAc0BH3Cq+vShsA+B/HjWGycHk3v4vUw3n+aWbOdIgoCYO9+9iw
iAQfzdSFsnFVx777TBa8Ek0b7TFHvFjG7ZoyAneZnvvSXwIpyBJIFBSEnlDgS6tD
uEByL8cFG3+42+SBhl/yNtMdeFNWpszOiL7msdq66TCE9R/jC0oyceHAH7u2DUxT
OnE8PUoXAeRDEDgLgTOFy1RxbI6S1bQnKhw00xzMCivKwx88gYF9nr9oa4/tgufd
ndjdYfT0f3s4DBbF9hd/hsU4Z4eMLlEbmJcVU+YLtVyzt+/gf9OLk/su9p7RwAOy
EBNB/OY6i6gJLND0ceHQK6bGCfWuH/W3U1HqOQk/HXGaLP5crzw9OqN/CGerzN4H
F6ZEIUMBKIDouQizsbA1F037EQiVmJ6oqaBtGqg+hF1qlSrW4v7TS1ZGXaNUCIUL
sl7vv4Tq28/jm8OvP0FhZz6loTr3mhPBeYRVBOsv/cUScNdg430QIP5XHylbavnI
lZGXer3CDQMDSTbOzBM2bGud6n0PcJHn+RHTdjqRty1PUGmbqh07QkRGI42Y5Iyw
w5If5T2b733JB2UxbPyIbMTdLJma6A6L0opgKyoqcX6CBffXvMYQXxDNqsvfMhcU
c4VBqz698edNNZXiRELliWoKz/wa9wQGOfBqjB/5pKC0xleQ1AryxNY0xanTeVS1
DAdlsCxLOQE9UnS8bVRCnKNhLr1rbThVnY1a2/bqe+b6FEWM92cscZgrsEjjnlMn
mU8ynXPiyhWnmBmkiSEmOp6zhZWkzLlq7TILvG0lC80jOPePogbxbI44M+tvRFt/
r15Dq7C3FBjSZa+oaDHJC/HfX24quIkiGDSNPeaGe7GXwjSjROa8D7JHwDgLbu7t
1EFNap5EOAzhOag7OkMYcwY2gPUa2zIMbQIICJAFy0mHP8Oy0KWTgq8WxdgAJJMv
AGk3hHUcJgiW251NvBbRon+iNsycYJmJwK2Vx3UuTuS6++fc5mXgVpPaydVDDIur
GBPcmGvbiQHRI2b37BQby8VNz2+EtxstIZrGOJZAkrEZblMX6Gfwfd7hwxE2BUno
4JGXCSnfgJwRrdu+mRjJHqSvzmOWsfR4hjVmFE0foZ/95dDZz/ZKzrC9RSUjlz2M
++bkp8ud3mSFwoyNqAgzS055/KQ/U9DIiiEfK/4TIgKa/BV88E/h71sqZ0aK+Rsa
DbUtbsUDY0Fle0PpY7jVax8N9RZFlG1/KByKovA9fNlWY0Hl1l+HPK+xLQoM1IuE
XoBw/oUb1JAjuqk/62Ds9pzkTJOJVKZwSOXkoC5faWSgoh2cgPh7n7MeQY+gcsQJ
1PCwm4msaY8k5Flf4QCkWxYq9BSaI9Jx7bkzkbmQU45v3GKRfOaJNBpTl4w+nX55
Q3coKkq4bMDtg7Ea1jvCqRGRUvnna1yW2TSMubh8UkbS7/vPYzJWltGg42zKCGEM
zTdljc20s4ZhP+kiuT8iaonC6DpTLvMGgq3CWwmaBm3WQl9bCL5fWxSVwHiTAqoS
djs0bDTAzgOUR6pwfIuhbb6ty2Li0O/9Ec4nD1+EM7sorTnSJUwThl7Mbvzq6wGh
gj5s7qFUnvza3jJ7SrY3vM6BlYD7hE+MG4papprBgtDX5luU9oY15Dmbc3MDeLoh
KhkYrxLHNsjneed3uZsq83+CxblWv49D4rE0aRVbecs4Fh7ciQ10HSNqZ/+PJTpG
545dyaqWR8eFt+jSppHUqpd/E051mtHkWEqW6ly//oNZjaGUB1MqkwfYhXksUylm
LtpDk6cR/1ANDUfpt/T6RIqFX3aFy0OcnSE2cN8miRVV03tXjSUKjEUTnB0Z1S3S
KUd8OIYuRdC+5m9cAxtqfWLw02d9ewuVGhZl73DTe3Ia+93/0BB8IM53sV1ZRHJZ
5wFcTecAzsGbrYn/uCDWeb5MPDGJXChqMBKFYcXKVBOu3dEmUtEHvxRtZ5wrKHRO
l9pXCZtkTH9vRcD1E0kDkwE1idu2VOziHaQtVYba9JkH2csx1EQOSNYvye8eV1B9
uwBM/JgL7ZR4ad91Ug4qzlmyxmIgN8YLprZHANzjuPCiSZmwqMzDYV20InFAhDan
OcCWcLDDBmbidB2Z20uDUg/oK686FC7FXsniDNQ/0lgXfieS1xW3dXjqCQ602/ym
hO3wxWHTXpurhjowYLsqg6EMECQsoD7n6X+LjiF1rDfjxisdVpvBGeeJ+QX1gg+6
dMlr9I9PNQjODQyopwXuEaX5taH6+ZEsdvQEcTBJb922gvUUWmjV1KcN+zWXswBr
vH9k19cqOvv1SbUdjhR/hRJI27ww5FJTj9c8q81ZTC/tFCDamjF8ksEOgDItUCEH
YiaKBqyrUwID2nX30zKE6VrUlqJQpBK8PhOrVSqTtFFp/dEgRn4NCMgIhzvvYTXO
T3Basgu2cSM0aspDCkVzefh5QcjA6owIF29OExjsF7GJJcg2B5ZE21/P6ZO3KcV8
iwlyB4hy5ZOBeiTa1TVK2KUD3y5XjnoK/80q9AMc0mhjvSKFjS4ysQG3m/SVLTwi
hZjcwfysGf+EfHp7BniK3+CbQfIJcsdnotXW8hkQvAGtd+AH+CJXlp44acdVeIGl
3w7Vb+FRsytjqO3IrXTnt5DEGQa2J4PIRE60XQWkEAO7hWdkCKz2RWDJ75Zyze8a
fO5Wbp3g2gjSY0LzBrHH05+g1J3csmK84zNh137Kdl1JBUnSRi0fF2zACHjtK5iv
ETBeoV7PN0CFore5lBoOLHGGND++kBfPAgWDlvV8OBaswT5s6iNUy9uHUZm6uMys
Vf71J4oWH4fE9LkAXKnyyZ+mg5hJZSBgkpXPnU+0o+UBIlvmLlk+u3LWqufkn/Gg
t7zG3Eewb5gA9XJBY+M+jripscbBNuRS1YheI/fnqszksaMShSDJeZUivW0INlF/
IxPgo4Sl14ViYA8Y64fMWVbQV5ffgTeXAtMEqwnrbjZe18LD4ra0mkpX12J5t/hg
QJ4fvh6ViNt9oqeBrvZUQiPDDGrrekSjQVaMMZPM91FqhJ4HF/tv7KO6lFn81hMY
2HGE9HEenTt7afOTi4m3O5OjKkHdTRaG5Xoq+j35rn8h+TSKIFLSrgitDl7YyQDI
xgvFhlaxSPxAlgCo+ynPc8Kpgf9m1WUSORsoM5RkfHawKiHbfiHwueG2nZWxFDDU
fMktx5ksR9/w22BuLtXYt2HSZHum1XqKVdn9U/ZG3Ui5AksXRMt9Yo8LYru8nDtB
+rh6YXAis5STfsfos4f1GPP5oi0FzV53sKarkdpoMqL3MFlBdg0yX6rUXGW4aLTg
hnk5flVQ7vFLV9z6pm/UFPSkAE2NI7VjqYxAWevw6BklvWutaFMdioOL7ST0fYR3
Fr/j23x0Z9qZW97kMF3HZaoSuiEWZ/MoLcn7IqzkFvibz1p3YJY2MDBsJM3RW675
3XRrukrFEZU7k55HOi91ssU9vPPsBoxenMWWihmTW0kGt88CsrXIIE+akxVy4ghq
Y+DAPtCNWdXkWGeQt7WzGuJDzfqrDSC7v77HcriTLPmjcDAiqeJTn9bD1EcGH/P7
KNZS/9GTt/diVgVVwJ5VdQEu3SVqc0qf5/VuxAvIwyUfB1+7RpNVCRDWqJtbOTSq
orXjEydD5UrMaNoBS+ogkGUMmKiDIBpel6QT2BATUQOOcQQyRUXY/6WKiIAg5tMt
esJ3i46T8OvsOYzePaFXQq+B7iTcTSFk0bYV8H/bTx0hociyOIOFlmJdvU6JfeZ+
3gld4ssKrK4IYhuHz1AuWmxSjQX5hisRGTt4jmvi8Qv/xtks8WoR52z/HeSvov8L
F8vsEg2JmfPHjcBZJCraTAgALqWR3uLZOAw75s/lLzDofLP4kK7INGFRQUrn/gyd
lPJiUyDKO+vH/NQDLpzpqVB8/ShLZiW7Zzqcjlxa8t1NXUCtiEnsYGYn1o8sH3zA
g0t0W5+fjmqSptiFanNC8U9wJuc0KTF7PqfsyKhMypHQPumtmReWu55L7BGptzc1
lStgvw0dkqMlWsp91z2eFxZvx/GKrqevKcdPO0Vzx0XU5ZGg0Q2NdMvjjBaFaXx+
gxYgMzoYIvnUEmAIuYfuq91tS2kidjmSsYUr8M27IMLMJ7eyVdYNx3PFGrih5IJ5
aZ8FN6AfpjJSZXnZFLdmE6uXzBPBWxLp3SIEuvCBmvyIKRuAGxzL7aZ/NkIHnTx1
eXdQ4l2h0jmtRFJCanVH0nHpNdmMkMjX4LbkMLAiBQs2xU+sOmt0J9iOiInWUYrw
vrKj0KEAUmSLbipEfP3KhqLMS2uGCj4JyyOTItR9dt2fQyjGAWqDcAgITi6t6PX3
RP+Jv5O+0BhQiFotX2BAme730SBqr19//2Zb/lPaFwDuP9f01D6DUAts41+ZOXlo
F4nipIn6aoubfon/NH6toHnI+mBSqExiDDxbKKn7ZodRAuhNnW8FJD9rJLuo5eIS
F+KOJvGm70Pwmjyn3iZfWMOFWMGx1JSaiJOMVY6cUNDubtnQxgqgdeO7bjPKYGZC
qdySCBgdzQZGQ0AFhqLsG9V9gx2kDJBw2PFbHe+eYhdF7VqdcSReAi0AhwGGZhKT
USkVAovdERrHJ/uvUqGocRHS2mKGoCHvJ/D/DU6zeTpxzg3Iw5kv6jopIg6x5UmL
o7OSHTLXWm4v21c6SqFIwODlb8HOyxMc3J5UVwqsA7ZnkqDVucTiVfQg37PngirH
jUvbL6qwXSnY2kM2SzeztUvsS0tqwnn3sIQXjrprgjRApxIBSeGPbSmyw3CRAXSO
Xx08s3VORQlrMLTFOC7l98Whbwxhv/9wjP1hEU2lp2b6nWOfhJX35HRL1b9u5oFZ
p0gaAljyhPEAcq+fBiG6SxeEikHL943OF457lke37gFMVpdppV6eSZVW1ZWgaBfA
VyvfLdaemBYJ8aic9YJAMxvI4h4Qb/gesDmW0ZWSl0kbQWWrlmFgCF6/XAEQu6u8
AX6xbfrkj2bPRQ8yCfP1vkN8W/vPDrdE+QDkpcXjkr3q3zCGbl5rsMl2k5Gc6x+N
Ha1TQET31AyFJCzEIxmvPlXsseMmfULd+/wN4zNkfaRYApAVxXkNpViIq6Wvs9SY
IIULglso+/dVlUYTbcGGTG5XNe2IuAY6cQV/c2nBt6Nnj0s7mbyrsKJRugfpSZL8
wOvA6Dd+6vyP4TkwQyObK0zvWGNbfbe3wiYnelG48Zp+kMBWqGtRAjgWs6XMPlAn
kXbTx3KjPN/QzTAvnn5PbH+Ye7Ar985y5Mn/28XJnBkUN09zClazaqeVdwgtOCbE
LEQGQ0OPSWZGDEedQoAJFMpV1Nt4kNDo3yJEBs/arjVORCmTgSpGISpX9YaGTew0
RqxE7FlUBXVAtzdWAiZKhbETkl83Y8QTVgeSIGEFaSf2fQNRfvqWq/ff4u5RBPeL
IJq5Cy/cEEVaGjHqwd/13IuSn/3o/LDURictWoBthIRji+9eZlg8t1FkP61Eh9JD
8o0838Yo/DM0NQglsCcK1wFBQltTgXOzYDH5yF+u+Lhp0eVFUO3YGwgY05Z+AYX8
hkg3NhgirXek+eE/IvEZXxdMWhxEC2MXS4oedtzv5s+K+TgZ7b0aMRPTJs1uPThk
CJ9kdYrxz1Vz9adinwI95TysNIhX9c0+RYJ2G6Ia4OcY1gJmjJLrA1mfnJ3phN1p
R/MABwXccsFDu2zT/onBCgLyUXtFFSgCHHc1SI4Ia00+IAW7xTFx2BuND67tFQ/n
6gh8nwX6k96CIC3r4Fh21hUjxDxoZPxAOIQTSbVVkX6VAo7yUJft/A6tlhTXnvVS
fqHHYWNLfNBo5b3XEnBKITYemnn78vQFSjNmTGouJBUHjesK5r3NX+qC1+Boebf8
p3CUrpvJPT3aa3u4I1gVkSceLnJDyu0/rMnhOQZq7TxMra0Jlc+INn0xGgAkFfdw
oBx9lL55ckWUCPfdf+w1NnMnNaTqYmYfmlTf4pa4PtOpxLN+EN5aJFlAj7UPzD1v
oUp9Gt1pB+ZE0zDqcgb0FSDlaxa+swWb5O49CDTFwgK3Fo4KIr+TdG7BhrT1SV24
VeZ4CMQLkMYi1m80EauWDgIl//2G5WpgdpAV1Bil+UymZE12m++WvTWYEesWEhEa
aHWfKGIx//JCqp2GZBC6jotBf7uqDUZDR6akHaXnwvIrTXf0/zm7h/uxVjqeCrd5
bTvXpwNz6IDLDaaLR985CJjtoIe7CDIwho+bBbP442v/I77ZFfx89LN5xytC8oL4
9ZBlrZ3zMIDXcafXmYY9XSyjcz1jOtOEgPiei2XMSn9fzRNWrgIRQl9f4uw6NNYu
PuY1R5U4I+QsXLVeODxSJOju+OxiWNhZ5JiYNZ6YFMbtmc7+NzYPjPRy7NddKvwh
Jq8u+EZKlqUrwVVG6H68c0xyFZxTRj26iCQizdAQJEmG78U3QiHVE7oBDtR87Ct8
7B+THkHBZubCwvV5PGEIIrj200+QBWis6HBBjIYavmsCunsb4ZpQtdSCOFFVDjsA
vLdePZ8vDODUfmPFIxOYZ2oAp89mKOF26Ugl7gWSQCUfFB5RMFrHE/9qauYXJX+1
8hrZjHJc5FxQGU7rbjEJYddk2UogKCzGI3q+Qzz6eBcUpytO0quqxXMtxwv7Gwv9
RmRA3n4OeTRcjPqhBGNJEz5Y3mBb5wRTM6O/359Rfe2XlohvHnjrf1giqNr/nnFH
BOfZxMdIyHtzA3AaT1hXlihpW3SewNSa2wlVhe8GJSfW3lNVKL1zON1cWXll/pcx
W/8nT/z+7YMLQOEk5eIV3daiqHFwYwYW8S9c1hGqNCXZJbULG3ntpqcJfSrCWCS3
yTMdSaclvz5HCQTy/NxJWQouXUjA6J98365DpYdxe/XIMdhX4olRGZbmp5lnKGmh
rsxpUVIZ0gUqg67mEwTQn19MqSgRMnZ6dYH04P/QBzi/4ONBqi/uJGFzTniv9iDP
7qaJK/svuFUYfIm+7jJ0Yv2AVENQs7sqmasPF9srg1yj2YPu3raJBWovFIjWTwdl
Cx0FAYIrXuX5zQoA90ZbZ0vqPYPdlm/5DdIKKSXxMYcET85ymGce5fJgjXQiVotz
Ya7AoDK5crjArulzax4WS3XPWyfoXz/aKJRb+rArGWCZW4h8WMUecu9hppiaNQp/
b2S2GOG8Mzn2mNI+I6PMWHuOtLjCGhF0On6bpsyJcwdAsvAYH5vgnipsT1cCqcFD
nQqc3KvDcs2u51/IU3dO7Ttvvi8i1yaPE0AsaP04BNW2ttkwOp0MNdpQXg0UKcz+
vPYihFaJABD4D7piy5QSdyxUkkV4YHmIVEuGvb2OtOgUONPkrUrQI2JN8PLtsvZl
fBNJKxemcgl30pj6bTw0tKUcvDhAK3YSTLfpIwnBYE+RH/MRRb7bGvlv0zZ4QnDX
GMUM6/1zjBs7GCi3qWbIE5AWvfsVf+fpqyjrncEWCckMR3M8HFUNU6f75RlwG3mK
fgN9bymg8+hkcjlSN4NBjjit7Aneb2VkBg9ZnhfdcGUwCZGQ3TbzCmX/iJjgTKkt
1NOlLaQ5FmSh8GKlxT7/rp7rWAT8WgdxHy6mvXU2atEeDxCMsvEAF3kLneY9QlCr
nBsDg8+5s70jNm079q751Jg920qyP+czEGPDM8kzbLiXlBfL01uGiRAXVgvkPM4w
fVGT0XCZmEm2n+ERv0vNj7rhflTrAMHNXjgqppd0wk0zyWngJ7TKEzIW8qmTbilo
p2rT9eK6DoV0arcPCChkJz351+NbV6gLHmgh+XHSnSsREM60S9JRz31wTh/UO5Nf
RhzIsXX2bFgg4P+CUJDoRuJkSQQ3t8LQWYdkB8Ya2gg1bYvZ7pVxkkog8fRFPzy+
v+e7P69s5QLVUXtuzQlF6YHk4bJU13FXsYbmWKFp5D7KdV4ju3GzatE6lD7jo5GG
dc+iDmCscYJlYncLfINcwPs/7dlxx+cEGZ2z4gfNUJfncvTN8ov3N+El9F3EAyoH
V6c3073+JGxBeMuJSAAp8Z4SzonpCF8Xf34lu6TP/IMkDllpSmP1g1L9xtiX1akr
14cRjL/q4doZy8gf/s1ZJCFptSmKN1w9hCcmUrMdZGGUkl1t1ZGJVX93Z2U1G1KV
C0ys3uA7/DX1/p3KZLNywNMNN3T9o2LQn5LAC8l7jNzRxr4KMLcd06KZwyB/iFqz
bV7jBuu2hdi6oS24RQJeNfbt5zTXsAusqlPrKFBZf7uXQfzF3qOs22BNcvxp/EqA
ilT47CMk6N9qyJzsCTtywYautjx/Hjigog0VqQGGM87DXyPHYNiN1+n9QDaL8OfN
AEgWM1YMUComuWeMekoiVAgmDVTPn5P9h4fgaS+IdCfa5AMXI6Z9qorkKmFk1v2/
g9t9Ulf0pCH7dEgpWR1ntCFeAhE1OY8QUCw+7JjzDmgpZV/S7FIqX+eenL4oKIIV
K8ERfcdyszZd7eI362VeJr2x5Z2pfnHRTRi4e2JrSVPHuojvE35xx4KM9rXSaLpi
9q3F1NPaDJiB+pc4pRCZoLYaHVrQw0sxDOaWdEDGBCFJE9UmhB7jhm1dKV0soSc2
i44ruQTa0KGIHZL1hAMrKFPkUGv4MxxzEsXJ086aFcNJBHLIDmsfu4/57EaIz8QX
BU5ShQmIwT4tP8krM1P+CAmy5kVTHJlPz3vQnOgycl0r/nfljBeF4o+U1r4VaR7n
rTmaSOWnHwHxjnubrjyf9TaVby2hh5Z8NkEnr2O65PS+oEhbjXdh9/rozFIC3ofh
Rc/pV9ceX/hLo9yKJB+BNxH6i2tIUkjgFrpyVxbLT9JyVqYDKzDCdYbVpyRE2dWT
t5yG4ovKbdmzuMJOVv+Ydhu+aEf21QxfEY84/zo4dPHrfw52Ftp9EUjkkOKqd/jg
0iY+iZzBIayc6b19b6Wq6tJrZ7N+htAQEXoSEodGt1u8XX9+SSW4bDRCYI6BzTBu
Xs+3yYr8jgev4c2IkuWp0G/bxOhqjHYvuDfuqS2+k2hsCCDJeSDfN4XMOVWJ0kio
VYnxJ+glgy7M8cbnbQSGBIHUcqpeEPK/XnCkL+xhKBq+wiCYjjaVAX1YmUCwDW2u
D8/iXECEiBXXI1/KFxV+01bmlq8DbjiTQk3UdDhj9HfkXnhGUC8FbMOfSw8FNBVl
MFVD4HUUlQRdYUi0PtTv3alpl4RyDq3yo1d8qdB7wevp9YDTJHIJ4hoF/vYnLSs4
XrX51iLrvXhTz/xZJg8Quvux3m4lpWdyAi99MlHzAlkRzNBeQbZR6vWzl8IN4tVM
oh7RiX5X9OInO2vVM8UdaQfhKeRmWavSVZau6ydeJblbUAGvyYW4CxGCaJNIXfEa
jcXJ9Ty/1DbdNNkUPVCfQNHMXj1qiys3o+CslgnpldBMzQSAcix1c1Wq6XDlSBf1
NiUVclGiuzpmT9DW+bPpqU3SmdHxlgIlj3jrbwebY2FkpAcMAm5q44nlqyQgY7/o
27JxGrYX9owx7Md2PC3Up1yQhSoFXgrKqYSZzOmTYvl8nyGDlO8f96HLaCMHUFoF
+go+jfqukwfdF4EJI0WIkeanT5SPhRmKkT2LcUX7AG5D60OXZ9sWUaSK3CCKwdKV
23Q/JE1cYlRwUarguwP6sc5yfp2eX3tL4JW3t788rtAj0dpCYs9OyFtkVMyzN5c3
Tll1LJVPwEvHUaWlSnoPLd0qA1V25vV0pweyn8jwlLXsRLxgYfddLRySrw9EZSU2
nB0z4TwpeJemPPmI/ffXPFb8UPU5yN7t6O3IxldR45Q/z5AlWFfjGgWTODUMmEp8
9srSFgUWQVDGwVzu/eAj8eBjVXitR/EPjST3kRL4SMdHWuKiZsPmxSYlNb9OQbe6
bQmTgb3cfudw7rKzu1NJPWoEbk2XyiJ3uXJIbYaPwC93idv49QXTJCAJBfiYMD4N
fVt7J+PRflvOb0yn3P2FRElc2f2mq9hj0e6nECzMYehgh9B6Xqy/hyyWYc2yHs6V
N7gsoDT/L7cCqtviG1zZ+PiidYZNPz5e7N1M8vhyNcj4E0IZtRJYVWX0BR7zZr8m
gXIEQU8/bmHA06tdq/Um4Meos+EExX4Gv0gmHLjvEB9aan/k4AfCRtV43mwmFMEZ
GEaHRGMVWuXtSigOm1yP/y/ouD7nIe+pMWeUob1FLu47MHkeajAfg5En7yaD6rD3
nWVVZgGuC35IKEGv+1QKTgChCzu7OwetNv/VEAef884vi+3luRc1c3L1K+nPrQjA
pz5ooW+qiEQaedQhN/xqn//1TK9lY2+5u9D7vvS7hMsKRKI3U9ilGci3Cn3jJ2iB
MBts6mQ8EL62EVxngw8fvYxXFk1xa5OfGdjbdQpHeSEXU2W9DQ3DSG7nO51GgGQd
2HAxz6f73AH6dZIdJVYlzwOCsQZuGhFWUn+kG3r/lCkc0SGIssTsWYCJuBImeCxn
xI8CHqqnvVWXgPStDyJakwatuFZM0Jgd7uHEJ+wUPJz/+OMx0a0X+Yzsuh0Is8Ss
CNEF/fbM9eYL7UMSs62SWusq59KbsUKhf40DMyFgDh6pQgGiiZpX/e9LAvX/HH6m
Ui7YnGq97iL6Bcss0RNsCWnceJQxz7AMtgoZWjb4q7vZQQZaa6tynAjuSe+UfYYn
w1+RfUo7FN8Zsd9TtEzfDDZ1LQcrTsKrP9cK8oLI26m9XVH3G1mKEGazvoIpaKLH
0xASQY84VPaOmVezVF8OQJt0IUe4YwWZW+zfOdPUQyxs12WnI9YlRk40lPADRMp4
XrYfo4WxSn7Td0yOWe3DynxTabGsZ4m6KB3pcYG7lrGf7VGXznIGfrb0eds2vWGx
J3A/2lm8vOP9Ak3fMVI75+4rVlxOKmTxrZhNRKqL5EbOYWH5r16UFHuKyvGGq4ZD
G2ZnBbcMtc/aZCT/rEKZQlZaDDPTi5SjSZK9Ohbsnu/lazcnPU84uUNFIaYLO1dJ
5zcZUvH8IqsBkZa1OyGJDKQtbuUxz140gnsqcmvfQUrYSe/FkV9oFLHDwAtgtGGK
szjanUKDt7itE4oI6az4IXKPe8cXMYNobZ6DTQRyMAZmBpMa0W3iNromVS5GQff7
Q7jODa3SVS3c4UyOarsEzLtbVJBSmX4qCF/RFMzb+y6rCfqYsF0Q8Hu3bJHOeu6R
gTB56Yj5haLf42PlkXUlKrgoeS5QIuqiQusElO7PQG9/IR079YUXXvE1wC9OaY1b
4Qk5MfWM9XhzgrGNPyt89bN6vN6aWfBTeMVfDvaCFzcneqs3tpBhbvXxaRbv5fJz
ae31TXva5Gq0AjM7gEMXODUH3RKlKZmPCWAPej9vueBDogIPhJzbx6g2NhNwfrk9
jTdCb/6iACuDkBmmnMfwTeyEnHK+Z5FXd6ayUDAW7oanV9TmR4HL1oQwF9inIqHb
91hFEta+e3fPRHV2es4ufr1DyewwrNTzqysi26DZm0Ch0ZVUgcKAVr49daAnWcuk
FXOsHML4WbU3uzdtCjOQHSpbXol9frsxEcG7lnjs39QRhxvgd7Tl//u4YI3D4n7d
/A5FlLLeHmO9VijOV1HTDHzHPsRAv76JSRUzVHF6ryX+m1tv3UrmCjZx+B5tolQJ
+parMLgj7WgLOi8sH5wWrIq4MCkjVVhzX/CdVNOXkkY+Z+M6ckK6UJ339AW6xN+a
HBjV3a9w319AcA8DRMwQ2sqwO/fn5+Ko+Cu1GY3ZszsHH7C0jpkrIrT9Z5NUwRjj
5CKjCJ1MNJfE4hKkZPJeuGFI2pMGMpUeLlZRKtDgapQi1w6DpQlTFh+cmkHeVsdP
WjzGtr+lY+sQQ8qxpONLbO1Ux86w0txWENiWGwXzjtwm2MRgH1XrYFf0lwA+2Tqa
T9zh0lM8T9DL30SlrdOeFCczqdD6HLPzKwPKU0wfkgzOV/meMAQ8rElI0yWowPtu
yOcHiGi9WZLpz9QU6zT40N8pgHk2Keiy8ywC2suT8OdJ7DihwDEz2kYUN8/sSsGk
Od+T/c7IpDbH//f86ZgyexWH5dl+/qogdCugyBRA1Jf0oZuVs4+wdBuwBJj4TtGG
bqys3biI96v9j6nru6Htcg/Gq12qh00W8wqGqpllvx3RsknC4Q0aLrY16sjibDdt
wEVSSTH/+4f1YsNfvO9Tw7b9kPiJHw+rFvL5rYCTrwokm9lHe4yrKRIEL1W1mRkL
NsGlV0PTwCoVD1coopBL3ZE56cVtudeB2HPISKlklc8IuNgJM1XkpM/UvYSBnthr
vazffcA4ErFWEkxtO+8cQbWS6iilhmrV0Y2fTetfv+fQNUrWeMkntLjVZcfuy9RR
noPaxF+go9ctUf0/BbGVjGGdZnAeMapi4XL1TXtqaKWc0iQ+CI9e6pnCKep7pmk1
IyeyHTmgWV/1uBDc9IslH88lVy68/nEtOrBjYK9k/3wDUaNKTYf97dt7sULBYG/T
Ix7PEzrCovY1GgPhSK+fLgMFQt7XKhiHGYRxExijr/mGIQ+K5edDnHe1PClKrD3A
u3LrwIMSEe2nGayzgbSqFufu9gNtkjyOSy25kMPjNbUL758PC5Yr5bfCA06BmW1u
etFVJHLLRJFx7CtSl8QSEDJgMrg72xdjyB/xKUp48vuv84yKwIcDLewjY8HqDOqz
jpEzIUULRLm7WqTsbX800Ihrk2eWgD1rX+u6YK5ZTPJ8MmAaiyRCFJM6VTTacGJf
wTMKct/2aOMEn8MrHsTC8xVBX6vbtV8Q+VjBimmsrl2FiqnKxYjn8Xm+LSag+d6Z
9Tw8NQgdiYzNamdLMndHJ8HMxkknw/Psi5s6xD6NMA+09EDxGRgVE3iZxoznq8rH
pljLLKciZVivDFQxEz717AYI0ebuGKSsceq37Jvl+q9JgIEfv8lOHs33mTiZwoei
8sOEMe3SnnYYBIHtbbbqKc3bA4Zny/l946U7SnqtteClu5aFjMbRVH0m+Ivm6zts
ziM6qb9cggBAnDkAUrx8TY4dM6UlQgXC2ARvZBcMsvSbIxmim8mzgAroggf+TNxD
IbZKvOUJyiNvi1rYRT+MF9fkbfjICAX0smOvZJ72pdtNozOiaLSVG/th0SGpUtSv
J814emJ4ZmSFCNoBTVfWxIJAr4/6RkX8L/EtJ7T6tq8UsLiv46K3nlfwCSpYlJVg
sQjZIgwn3bW1GYqykCCP7z94FV4qyYUQAAoTYDJn854AORlK9EPRrmCh7DkDT0rL
YH1psv4S4yo1U17Z5PEmA1F3SysoFXFom6GbcmOYvovQlLQjYfMfW09dW9/58R45
2OS3T7R37Ik2F+R3rkz73IorbugXGaVPHa2CteA1zxwWAlg15c/9rn1dvgmUErbV
Z5EX1V5miPU0FRRl0zroLC3+X2rHu74j+GW3Wz7z0ekftBj7VMI77YkzztkBQEOV
X8xdSGz7FhHhoXCGpui+O7waAT+vnuVZvoDTsjqUfkUKFWjGzYJbBtvaEtfTpu/A
tKBaK28uxWdn161EwCiP4ZBAh5BpSlQpHqGMmer/DESaeEticBLP+/+dRHTK5C3c
lYq7dI3FQfdeEhxQOZ6ccTsGitpCW4iqK4LGoh5WC8WoDmL0HMgJu9q+r4cwAW+t
XJdlZfry1atlJQwofkvctpWx5JI5ZMFOo6u5PJwHk95iDtXF9OZQmF4SnX2wz1Ko
E5Siw4+GOG/Yr6mBvHp7AECWF2CmJ/a2HHYgEqXjyzscCx3UukkDGO0n1aDSQODE
vfPpx4pxU4V0VbouY4Y9l7PZ3ri3vJ74YMVsFRAyLRoKYfnEZwj95tzg54pCAms7
OVSiKB0+QETzL4V5de77MSQe5mOrHimx/GLAc+KSHpsQI6ObpbDSo03/NXpYitmD
p9/1XHQKr9O2svBZjCr6cG6PjKIBKSmgHGF7ijMTgmyOWxGxgP1jP+Dyn00c2RPf
3APyXSE/M5e9nA1os9h3+L4Icd4646mZMN+60XOKThuAEnP7Bud0qh7ltNryIwyn
1wV7XYi6AhRdBjgl5AbW+X0Rra80BkgwTFIMy9PkBhcVBgreBz8fvRRMCFVcKqn3
Zbo/1xSY/ywHP8DoBjhIYfE/cPNMi+OfgGRf4tVFVOrLe1TeaekR5IeO3NaO32/W
rTyjBOZHao9LaEbH1G+TnsPM2c7MQ9w0UHoU6QzGgWQC5hEM+F+nWlTNnxA/AtFp
4itzFhJqV+RiFIe3rtVoby1yFqyR/gVne2XL1+LdSJth0Vjg4mDLat3oLpaEKZgm
zPyzAwgSy1vUlZsKpdPNSX4yOZc4oq0Fr4GYKDS9ARu62M6AvcfUcQbvfJj/jpTG
DDj/7N0TUxYa1+oKt8FLjPGrcn5ZBPKofwHk7oZe90AUMeFAMtZlZjOG+ZtZ24O+
knkM29Uq5NLL69llZfGabGdvkQdYPafN3L+2Biievsx0fayMb9YnbhObSp1jyzHM
noiqgUdzwSTN0CEWBPKQ7vqddSSlAoIJjDuR1rROgFf01rBD0CQz7K7wRzCzm+aV
ErxDmaJVJh5/ZJ8nHDh6oqcfgaRXzv1ZJ3te3gy3bG9NhBRsLaXr92gBBFUyq/dj
h2iWjDyUNP4i2PFlDU6jVy3CnKfAKpwDD3sqxAPHrvuzIqro398tOWIjhcujE3yi
6m6bLXMiy3i6oiHAvgfJG5KVQWLlxybquqwF7KMuMFNFXNwqdwKt2AuwxTy9MQ9C
JDHHjYjisOB4frWWahYZ/ZxGg12OjpkFpdwdVAHS9fGjfGlP+aZn2GBO4fhpywk4
3KJ0PZWzS154uCU0TJ+SFBcUg4HXPTWFCdelpkhy2wZXA9Aj9p2dg2gqvGyDpXKt
I10iMJOGIWNn1JILlKVCeq5CpvngTbNGygxlSa2O0Invz/uJxXCfSIU9NLYS/UO7
KRAXXeukUQT5w3I78j7dObES5HkyfRtgSKenb6RU92Zcw1KPB2DBD8mw8lUBRp4d
VLKpQRL1RSQkM71l8FWuH22gTR3Va5gFEpn8UHGAnRfN9Gujcgz78S35BI1fP+EL
dH61RHl5fvY52gNkxPdiPb1FKF03kKCZTzGr5xlDhuk8sHQZQI2CMaysmJltPkR/
sJCUgCIc5tPcOcchEugUpvWnYV4g7wNJeFHXGc1UD/FxAaWsBV0N9F9l4gQN6hD/
aKxFkvwiLaLq+hNumDoE0jh+yNVlMrCzou6npLgJKrnbOEeTl1nlTGxNYxfwm3qv
CF0kthB5m0xrWpb0Du+iVN2o8Ret0mUqivzkQoau/70uqP23pfz8ioODb6wxO066
YGnRuWc9hZYcl/RJsWe7H02bKbr3f/7mMcWeXJ64IWpH9+NsjG9J2uy0SIE4T+y+
Qrt8I5O5Ytmzr9B/y1h0FjQHh0eW3aIZG47o+JVZAzQ3uzXlgCg7rlT12g6RYKqq
HFztL17UsPJhyY6sKP+qBTrBpFSDgL9l/lkR4po43he+PvlRVANaUTL2wv4AttJb
RSW8VbVyFGuIjglIVQW0yRaCJ/anLMlEh0bFJeGFHVZTdP/wGg5stPDar//C0dK6
A45LWx8RTSxhM+L/drNEdutezdleVEKvKG01ecCp0pfF9SJ9EEIh11agZGDT4hvA
mtwDSRRxk96vVH1R1f1PwtedfBlSDfJ61+dbeDT82DYcb/hWTgtoWw0w0q2TNVrs
qGTMdETFS1+CtwJafIfrBMgHMkhUQ49GLIueZpgdBmXOmJq558Cb4lJv5DFLNnpo
i1ymixs+88mzvQKkMof6FjiBUpR+j2XLVf+j0Kf01FwY1GU66lGqt1vhg6+1GI4K
bEDix+K9tQNwcjKLr2h1UDdCbnMck2s6a1oCKvNUdzjz7n7yPIUbvjFFFWi/MSmH
Aw0NYeayaRGkxJq1hXBKjL63xARRngOFbx7E6ChC9oLkSbcPDpYy8pvQUUrXWse6
ZgjTGwZKkBaL5BcTebkCCiBpDwvhzAW4sf9VTgSdqFvpBblncImfI6MWBMuh3oky
EmWwsJgohQKeC0IgUeFImOmQFpS4dGFvfwEkZLbsszXnJ0ey6040Bpcze5hcodv6
t+5VJFVqM7gEvVpndsMX0C00jOkbdQTw6th0ibPeUdgmXa+GKV+9//F3VvBV/eTJ
UY40+/bhO5JJhvb48kHPthGoW0v/hgQeVWtoIto1oyxWX0RrVIqhGJlswJVKf2Fh
MKRgxKlmB//cttvO8wwkIgiR82xW0v79nk+6JYsbVeea+AeZHT3fuevds9mic2V2
ParvXHE5McpwH6zFL++hqaPhs8Q9vle6vxXRuMSbbmtBtYPfXZKosuJ1puF7vYmY
jodNHxzp3I4Ec2OEIJt14l0Cx9KT1EXVk+9IiDOuzeW2yxR42h6c5ajLfOipOfyV
dALow8ugmdujLVAq0TQwjDlnGN6eoZ/Eo5oQ7p2SR5lR3H4lJSK+JWN/S/BLk6zC
4C2ewnr8GCldThDbOxFUQ+GvpJG97GmkeyHZVsoBITBtEa1f9h61FGhwduLQwoKd
525j1AwGmqKD5UEcTA45jOvTCaSzfLiAFDX81iOqDN2YFQ6/5rEVz6RN1Ss3KpHp
FrWxi/j7BrBB4+ssfRqDg91GtxvZisVuUd2MpUxqSo4PGDfp3xlea2nwRlKZmNrm
ElOafDfRIwIJkaw/2pjTaUDNt4YdeLKeT01aRfYELsGktcZeAA1c4QWTn53tBW18
KYDIPHfhgFSezzn6j85smu1M8n7Dm3Ef4e5fY+s6z8QtrNoS0ddQU7jO9EEg+Ajq
D0xyk7tUFY85okIgVruIOOWv8kK4asAhEQHpMt6slLW5VAKOAl5IuQC3riIWLGZ+
o1dBoIigvAqrUpW+tRkRFCXDbHByJvRyxJAaXEXhsoZFccdvVWvJqMwz5YIzBq5Y
BQMTaA7cR2IDgWq8FQXJ68BrQXgatveZykgssDlfno5Au6aHksqVzpN3zAwsLMLX
DmOZWc541vhYG/ZvVzHgasP7b02ct3rTbaIb3annLdzNR9UirAgy4XAYPQzcWARi
A5j3jC16wkEVUQQM+Qbvw2cKcC8oE9Bc4LoKpkiR3t0bA0VXr7pofG3jjqk00osY
s5ULc2L60J3iAedhSWecqjA13ENepqBNNtQSsU6Ez0XRwTKQXDRgD0T7b4kEZXgF
ZQ3ewZfeetCZHusz+zThOcBCHt1QeJQG/F1v8EMnRhbxiq+WEPpqwSGpgbuawoiP
gyl6me1Mmv/0L0BRn8AfMVIFV/5dpKg+evYkgjPphVe7sNm7X7iqmK1OQgXc4iyi
k/tvVVMFFREWEGCVIo871Rf2Kx75bUkdIu1b5DE/8HIhQYrMfJ3eF6jmOcFRBoB7
cfDYAT+1n2dikYW5QGCjaZMgwCyZIvRCyCDDWNW2A8zx4mCfiCkKQVar+wYto2If
IFzVdTeXsm7VeLdLlrNRRdwXENnrS0UfryCfFxOSMaFsyn6k6i24EJLGrB+ZzvB9
10OB6XylCEf28aIL5Zqm2xqZI0SurU36Us02y/hi/i+JRpYm8KEOHGU8It4wTFAq
GCxC3M9TS4uVNIixc+838kLNRn/FFAwCAqTxVsvzz3hMtxhBH6m4morFgYB4d4LI
ZixrYMJYN+EQayimv8dRFTidIJ6NxAF48zM1TBsexTkCvQfuckZJdPO9nUwR7GpT
g285yUrCj9Xp040/cdi0a7Q2BpyNi6agZxqKwS+9GhEN/KEHKVSruTWe11F6nOfv
WCISNJJRZ7KiOPD7skhse21oFUUgv8oa9qcJ5oFjZIZFNbFVlnKPSwcukrgBZI+v
xepIlv/d4MYmBI4qgELqBtJb+VaxUg39tnB/W8UmQN5qlE734sr0tLgLI16rKpoW
la1CNcnmHRncJITQqeoX61lFI48GHTO2i20JennKPJ4DCThOUZ6pZNSYK1y/8aQy
qKcer75eW2SXPQfeVF5vDV/w3PvX0KgQ0DLK+oIh0L/srlEGMYxS04WEn/JKvxf1
2g6rZR9hIfkhm873nMHcbBsrHm4H3rZ09meA1Sqlvl+H3knsdKbxJl04mcFCTDjG
jS+ZJBJ7TV58yoYu64/s2mKaSQ0rbS1jhZMs1IO3cVUX9pt1ebaOT59K7/ZQ/gfa
/iW4NbQlprCovuHnjL86KFT3OcroOVvlIk/a1gr6rYdrT6CUmiRrJNB9TXyPF17K
nywLg5+RYfPW0sagpcGumP9wdWfOCgP9oBcndtSI2fG7Q5XZhQZEihhvBAsWVn24
3GcEozP93RguAK5rmB03D6L6DwgBXKv+JZyuuPOhzA0X+RhnFmIyJkyiEw59Qv/C
qCqgBzVO7Sgt3SkpIdsACu9hXM+H6WLLIICEh39uqnjWEZ3triF30cTrUKixp2/J
NJbjaxjVRvbcFhCg7IdJX1vhqkD+SXd36AVkw3SaHAjZDqwOsAi2CGzDrWzFFbtL
zrdXRU4blZ90Mx/ntLtRRI4oQHVBC86lOVcOUEreyomtobA8ioaVtvg9tWRyu9QD
juuxMKh7VuITQBxsOor8YsfMac4uYyjC4Idw8l7FBHMzJSSj71ouml6+5DPOiW4W
NZyCthXrGtXVKL6BvPOx/BM0Y8YozpYz+I15WLCBmGB5U426UA+2atE9jCYoUsEi
DhCkO4OtgLbjK5s208LjSt33j07IM4P4Brg4BSLKQR0pNlP2FMR9KVS7TxyAmf0t
E24YV90mh75kmKX8GsalTqSGpeoh5n/7hdJe8+1Ej67ruYiZm9r4jX3lFP/URrI4
x3cjlbr8dfdmqBnPs7ddlteLM7pCAXdx2kGY9stLMMc1FN6TEgqyuhnG5lVfTDGF
8TlDVXFwyvcuLM/Cz3QOrAy0wuZYBEZKe55Ym0/JgidrBE18frQh8kW3Ax6xdKF4
gEuWqX33IF/1PA8Hd38EirqWjb4iO44P/WPgz46V+mL6+kP3Vbo5MhcHuapQp2NY
jLYdgbPvs7TmoaU4RttCf8RYoTjy01h9zGZKZ1VzOt/zZn39KGlJNQhaXe/M0SJ3
7aw0Pi3lJ2aaeEkxZovKAlaLfLBYDEMqnOXaKxIoOnvXGODw2N1CBppp2qZzGQjY
b91REzI2KaBKXjqIu0g27I5IsJilHHE0iQRxoDQiV7BVTqbXAYrG0YnI52rCYtSq
Cc6sGJzl3cOiLo8PiJdxxTzwa/8fgenpRxm/JTMHP4xhdMFNrHm8F7117vhzMcwg
clfU5QYE2MuVmwzsyoR/KQpF1bb5NXkWDXrKjf0Q23PRxl+dkpM0nv5R5co98lC8
GCpXpaaQhVGHUHpbkIowFhqcUMfccGDRcQZvWzXUfg9pkvG8oaXJP6RtTS0HrHT1
xbL2Gs6bxEFugQ8SbrdQ0N8FXwpU+8DWPwXfUpvnlUwv1DLZRGWplbdXOyaCYUWN
ynTgDOaQRto7/FZpqx7vfTbEff5cHZynBES38rZKNATdJzz9NJ1O0wxpH6biDBlQ
mATMu2ZMkayRyYPm5vKC3C3rQoA4udm0OVg5//oHurVSjl4WSTApcnPkFNQ29XiR
+TDoLleH39i7YnOIEMv+7a6yoaS1sBgneDOGYiNwt7gycweGtoTLwlKwQkwp/SrS
u6gQMk0MeTx5a0XsB0JnPmO2+7RRn9ihiEAyMsPNugP/cWigaYXRKZWrKcaQVH0m
nABNKMnQVsp0luo8xLpPZyVQxDvXE2pCumTjq1RTbTTC/vgR9Sum0NpHhIVNTORs
/B9SWYkj9HSd5XYSEPYtvyQ1jK/xGupFCcrUhZiojV5h3O+BIXias4DYWRLxhFVu
zDfHv7bNoGsUmnaB6/fOJRTsCsO4jVW9yXu7CUjtI66Bjf7PTkhw9dmPUc8X/M1H
CdObfR6eoRROR9E+yfaBR1enI42DM04dyaFYV9zx9jH9o/45YWdKz9yLsKOo66F1
0T0fJCg3nPb6N7QX5qsrJIynGlANUy+lb5tYcrQC9TqL3clBBL+Gxyyr86i9Zygx
07YagJdPi7BAj6Y1+joxqGOn+5UDg5Ax4cWvI/FVU2b0Y1B+mklk/QISsMy+idXJ
7XyNBMn85+QfhMooQO6BOTOiQhcARKoOxtrG3++BO4ccSnZVYVdB4CZHJ9xLYjG3
4GLd0anBY/WOSaIAjAeVlObhgG6WmDhY4GarJnE7icZN1c2dzxt+LWWtJKiFE2/2
5lGScpp5QQZVD+bF64p69jvHg4SvuC6N7MLSIlzs+3HGyexNxTEXUgAqDBUuICxl
PePg8ugzhD/2TpyEa2edd18Uy/4WBUd5kWERUsn7vtMyKq3KkEL8xXjCVmOB8SRJ
Zs3GDo64+EQO6NMzWIVNzfmG4hOouNHXPLAZ6RtMQ43S9CDJbEn+Jb60YjfD7YHx
VIitrCvKIoQvssEuIzuyxUjvE5xBttxH0jM6tetlPVLzPZnMUOZbtjszsgL6OZ2i
B9olSyqAx+RYA2Fudz2Mm60ndPSp8oxz2LAbGWy1GkPW7/IHAOBTCvet9dxeeBX6
jXyXxlW78R5ojzpzblzgjbr31zISF7YbCq7quCRbhe1fDs2hIiYaoIA0nQNg9Tfu
rvBOcjZVqIcx5YsOGKarVkrLI03iSrtsX3WjkSLgVm9q4j6wCZoKjtvMeIrtvQY2
1CyLUOQMmuCcCSgWyousPgnXy+4TMl/X6dg9qSvQZF/U7H2ulhH7p0naNRzyxBoh
6X08hoEXtV7ZpJAU2+w0KzOTnmpGGqYN0kqnz+mW1sf37Y5FkoHldQGNkiJbNjz2
dneAinfTsD+MpU0UiTCHiOvEusuwBrgfRGNzHHJABk9aPi5XSvuc4bDfPo3uOJyV
mfl1XIwXXL0sb0S4NeJyPOMQESpFbw2RnJIhATppBSH0Vkye5/skqlXm/WtTizZe
eYGuw86ibbFK2TEX1nn49THVIVI7/PKaSs5CE+UVdzWAGD/vw3A5RU6JD/d1JygI
hM+Q1YzAhquZl2sur68DecCSaUEuNjXLcl6C3B1dU9z+a41LbujZGvFNlsw3zt+n
FAq3+iOQiYct1jvncgbGzcdnscRsTUhIbXQG6Kv4CuInVeE32XH3DXweLNxjkVcw
5ivRm2kK7kMpiHW2+U+GDrgEzmW93cxdXhkVx3PP4s8OWQHO7hWhmapJOcSVd3pY
kLlQ1obuYldoq8YD5oV4C7YpFEpa4/hVJq3mHZNLHxeOJrbMgoQEPABzh/DAvK/d
uDnPeVX+idFmNXgBUO8IFsjjiwcwVhogAKo8EDMIFfBylHkxxLYL/YN8++vqwSUn
mw1KWyBMpGL3bLrp+Dbgi7vQQPLoCjDn4RjF8N1cQuk6rD/VzRqaU9ItfNI1UZBm
iQVafjqKS94KVBdpVsHHD6cRZET+cxGu62Md00Oyx8E+iI2ouyu7xlAW5MbILlLu
jWGx13DpGI9NIq0aYytjZZMqE7cWfh/FUnhrgIScBJIxLHFi3vjGoYLmx2y7iOMS
pASSq3KyTjy7ikizNy3tnSxpB7JcHEuHjktrbbt9SndCcc+M1Bpsiv2HA6GXsdzw
svndrVDKwEixDYZOa1WibZ9f+nrNqrw2cKIilLmfvFZea9tn8VMNxsvDsnvL3+Xo
0YEFa59NCjcSWJ6DQPi+LWlv85UJtm0gr8k1RBhB9uzqT/TZ+XkzxnsDvWpMk7TE
Uyr9YESIHv8rlMT4Kb+8jE0oHHPx5N4gFGDl499v3BcKP9gIk7OBr1z+m4fecTbm
2Y6WYFZYTv2AWZG0mz9CnGO5oqA7FCrYSj4Y12MBXqmxxl8JlXrYlkP8Hnb6KoL8
E+xqlQrQv8CSkXlhfsg/BuxCgilOx7cRVmiksWRM3VEAup+XvpHI3+fwnqHT7/PS
sbOCuJgni68zGp418dL24O/g8m7bWCr9YNtmJYiHllJgBSHsv7aah5AptVKKlQ6f
XM5cCQIvvGoZ8D5IZG+6gn8UQrLQ3s2nICiCzSqdPFs+9grny0OjplD4BmkWxIkn
XlUV9WbzyXUCrwvrn3xH11resRpc0A7j7Ql3NBG90rrVkMYCxOqr/CVzb5JghEAh
WyxHFARcWzIPkp1XdmBOsnLI/87fs8qGHFooHwL+pjceO0m+7NEg/UO2CCSPLWMB
YeICnUrwpaYqGRaTjGnPjky30js3BSO9SYaHMMzO/78Gv/VUc1cY6deqsc1saOay
sUbNypUjZRoNAj/pfNYxcyCyDNxUQ5Wkq4twO8K62BG8PqR1qnQtM38nYYr91Jf1
viphnOlHTfRu6rS24R4TzAZkr5iVbExMxqSCqbzjIN8Moyz5A/zoaoOsbOwb98T8
usQ48BPKSDeYha0fmzDhAC5t1flPG7bZUpIAgJprAvSi7m6ly1RlHLfNXEDAUU5V
VCtrYmvSIboxsSf3SsqB3Ut2RrcNtgq+aHPwCtRnn/iVYHhaL98HeOjk40enF/3z
UxlEniNGCZMlTO28dvnYhkPLdkR79GDNoQFRT3FgdLR1hslS3CmdHXLm4gVY+kWz
aMxkCIW8OjJcWciBBQ4FHopZ4k5m3LQdlQre5Eo//Iq8vXgFkn09rk4Ti/6s6qgc
LYAfDmHsLs+UCa3/Uhl7T0ebxbsr1ab9dVQUAH0RdYMIXtjIQ+RIVNGTgu60ak2O
4N+DPG5VJKeel2hDePUkBf8SvE8XKQBG1w0siWfQBW3K+sY4EUKGNWM+sTln/B9D
GKeIqYm1TDWW93cW2dtBYo4rvNbfrDWRe0tn/2dxd44p8lmi0V3boAgsj5rUP3bx
s6LrrBYXr/0P1ake+ZbR3wh4PuN62PrJacYxQDBaQ4M5wKSjatS/F/NEiw1f1xGA
eLr4ahs9+UHpa526Ls9N/4iyy3xG+/g57LeaJnAeW6f5DguAY0QeJyJVrWTceG2E
8BskY5nrjGMUHk4H9neXnK1SN9sSunp23WMP+FEYKjPF/OPicLROSrLtyhyi5DgY
5bI9XRInkUTDDXde5vlPL7ixAUzyoFrJRqLcreiJ9F67pVKQGcs9Pa7s9Fo8r9Ls
jLtUQqtIcqhdqSapTUmaqDMqp0xWPUhiWWBMY8SgznLoA7bxDkUHFK4WI5FZjSVG
S7rztXn77E+3z5S4V5wS3T7/ZVW+aJqlG6IuqGeP+XkET+Xpr6spnPO1E5zm+nE9
5tg9BorWwOaMR7KZjXy00e4Wre361u/vA8ge2tQi+xU1INK7BYMHKlJ2Ml9A1QPV
H22t7Kzoxdfwiz3pdt1GmuAOT+p66K1ZCq1bBdicKBWNsGD55t32HnBK8jhhFXpt
NNPKNuMU5GKt3QB0qCmiopVEpP14oYWdyhgRkSLvg/8GY82vV+EzC/C5b8YQggj6
8P8L4HYrdUe3f536q+qa6rjbUVQV17/t7+ac+PU09I0rzZdknQBvSCfOE9IZralG
+zAgtGdmL+jl1zpdYyGdkdfWFAW7/aKDmnxeHR3mAyfBjB2F+dMYEJBPRqUh6D2/
hQ1dkskVmP8U99ExaHpqYXObkzkYgeev7HQluxbzJo6mEISmlHlE3BQAVnyzQ+Ex
8qyjiodH1UWVRoTCWVef01TGW/Kqr7f9Mezcpfv4DDEP+zCZTS1dg1IH5JlRz8Iz
VDXbX71Qpg+pjXiwVXkhUEziAeKrfQWg36osa/OX8qcbxnt4sss5CYfC07JdmN6u
vARBVeICsDtWMbMwA/hvheXIpx2KlToe130TR1vhYKmEkNuRxmRbnmR8H0IK/kTH
tNvWmGFhAwWWVwHT4X96P3AABQTDhWzamIViBbA/viE12xt4v2suy6gvq0SUKSZv
xDB3S62/Lnn7U0HjE1wJgULUAfQ6kWP3nMvJXsRV1yGA/kZ5EBBqOObmwBSIt03l
mV/gZXqfII3bF4OU70xhceXjJStrBJZYtHQksaSyut598h0AFbGPcCJ04oFQGC7A
JFkzJre70Oyz7T6/pqC8B8qYcVNwePovZncON4x+VgH8YOBo7ikZUf/RMLsIpdV0
UH/iVuV69RGgIXvYgkedhryUdtPTBk/pG2mg8b9YCWuKbS2udKAV2uaftH9QfDLp
AnZRxYj7ADCi+oxCAtortrksxWZaCUvDQPjtYuO+NVhuguC/SwKTs9+DD7zc0tKN
DPYAjrnpZG0e4AmHl5HiaI9F7++6CUNICiv/WFOBEOdXThHBMmlgKCgI+onF166u
sxrzkyr4/VrQBUNdPGV4fzzBmMPETuHWoH7iABcyMfVzx2fTBOMax2CKji+JDAt1
BE8cpdxkEUePa880/bc1WwHk7qx46B0KiMCBz1tCYRpEQoph63zR25D47JRXICii
HE8iSO24S+lC9qrer6h33dBFU1Qxlsh0mvCZbO4Re5eZFSWwihAlTHJ9UEF5rJ3F
/wGXIMGGuywAfAdYGJT4yAsKefXVWzcVXbF+3uDILvC+5nfbzGzZSh/jW5jYEU0/
CA1nQqVS3JU0XlN5hrX6rLB6cw6qFIl0+DiDT+VngrxrpT99+LzHiD73I+Shhdud
VD/B2Hby+/Hqzwj3E01GNijuoOwB7vRIZugxhORZ9lXOtSQFKVNY3bPtNlCqgMpe
F1TscXgedPo/zjRNRC4S7tAUI/wIdTtK6fl4+uDXD9lAAFMMmyFNvbBQhZGFv2xv
I/YkOvFoKKjT7elT1BpLKdZjNEIEuYZcJALmkBhAy5mD/bkPy7xvKjVbPBtxIBbe
78Jc1iJbV9WUxPFvqTeZtw9c3oCIiV7hLvdS2fqaR510u1CVWAERZp+BXDzPkQmi
vSkUDSVJOdSDgqgOhT8XLSAaujMyUrdrB1DV8bSs037jnD3LP4LusMhyBSOfL6cw
kaMjXmTdeKlV6Vi15dV3aWMXKDK1t8XiGWo6Dxaknm9RcyfADNeWLBQ+cLgZ6Eo8
2eTQlXxhE6eACjFVlKCEhQPgZ17K1CzcWJWCa5rN2BFw8dwJhGa4/HOGsH+DZSwI
KjqC+ReRTQ10OyLTBk4os+N6WEptxP+kuGQVCtXVuJ71eufIRBUPVul2u1ceu5lL
cxo9w8EWohGV4hdMxC6/TlImReenNmtqQLtf+4sFYknvR1rriVXFXl24Reap0ZKz
I99fmxKPbXg88SRNB/SbeqU5153aWghdGIpn05UMPTbJDGzu8nPsADjioQrAeqR+
hHpMWuh38bC8TbqA8ZYTkNC+zLsGHNfT8Jr+oJdv83Xrfobi5JRfswAvnIGRqaN8
BSqbitvrCjY3bxDIq4SaKTwx3FrQpgjEQQ1aIbfSdMG6HL47G3E6LWPvRL3jtUD3
4h0n6hwOi812IB4nYxBltM9TEhfPRez4rSrU5dZRDCRQHIUej+vBfAZLkisrab2q
4a+ayEHMfU73z7uAHNUFeJgS4WtTJS4orqnMYgIhlevrk5ywtlSWe3s0pgKJOmAp
dSZ2oyq0Hl+J/KJ9hR3DAmjxxgqDiz9nkMnwNNv2anAdNbaweMgc9+cd1K0ZLcYD
mNvtDGaoFjW29Dpcs+fc3N2Fc6dzY1MTcBiqmnTrcecJmh3Fom538b1M38nRpNVm
pI9R+n5OhhQCp/3jyBMzo7dNcoN7zae2cMahL3AGiRmBIC8S3aBF/KNafi6YTFnT
oSv3N0lB4LL7Ga7iBckD29cj4h0rKNGzuFqIKTLvouzo/k7GBJLJsGlKLRG2p41X
HCMez8WN5XXcjX2otDpYtfy24BbkPZ6TjPwEuk2+IUZi8nQcCuBORmIUxhbcufGd
BO5T1zm9G51YUDq0xSB080BEXhlrHYdY5spJLzrUW9BwKIpCTxgyFWHLaG9j7Yy/
hXoaltVn0ZjmkYpPtju9F89QclVhGDLrH4WQpTKjXmYC3iJQyydQwno17uW4uqBw
xhHFTatwSux8qrkj0EWVw74IK0YUOuRv9N+cQjWnPLuJ6lr+UXGIkIjGtwWvt/H+
5by8XFx/eS6vz/izz4C/3eLZAJry4nchQEW8rlDpYfdnwkfHumeXQXY0DsX0/NCj
3c10CpF1AflHO353/guY55yS/0HEaHBeJ+XYM4Vwj7QV6qrIl0JR+l5G7+h05W8y
D1wAbf4E8mw1y2XUBxnGXa7CKd7N5Zv3fTLZF6K9l+rY3MhZFrJk92b6BxuDYUp2
yBV5vMy4JOWsDy8Gckuuw+HaIFbT/oHlu519h5O2XfAFKjnkJis0XYeUHZfRf1l8
uIb4yr/gMV8gZmu2Otv+Yexvb4GGKVE59574FWmj9uaRRoGIaoJtP+ObeLQ6OSOx
6U0FtHrjmyKekaIMJu/gmRxaNvYseh445rPtJluVzgrbCZP1rF2k9oy1+7N5C4+v
Ip1huRqSsTwTSvpAwbUtfRNxYvu10+v+Xtdhi5ODBgehYnClh9Ss/zRd9itdAEmw
lAamVI4dCTha6OAMrGtifO7HrTduH6SbPDMF2kQ102A+GLxdxFd3XjEQx1Zgqp8A
xtVCVL+nqhWMQs7ZcgE0plTXXAfNpQzEoT3c8KnF2PlqTH6UX3Y0iZUnnf0MAlrK
bnhlGIfd/+HMEHX6db0Kxo6Dn8y6eiZ4dSl6/7nkVPxa/YKvSMB+C+qeisSuIcHV
sg6OHempDEw0bAs6ycUFVmMt/c58syqXPOk/arTRoukH4P1AVQkDBIvchsRZ0zVA
FAymF9Llwl0bFaIED1y0zBUL3FWkTFAdosOAOj33czx0e8V/OHhKKlAiux3o3Fw9
CEWB7TFHxM3bCEGapape0+jf0JnxJahdvnvNh5UD2AC3aSgkSwuqaDi2ENoe1slb
A8hVnowLquk3BZYbKoloZdjlLOqw4yCRsFS1gBRpNzC9BVkCqhh0BNTdnY8r9PoO
bv91lw8qnWTse/dalrVg/RuGZohgH3/S8M830qxT4RKlQFkZPad76KerPSQ4//vd
8OyldDBz5Ao4ZU51LzEsOM3yxb3SuweE4HEBM65H+sZUc2fMyREcBoxv9oRMmjLE
RsEnIMRBbAfPfEAk+r/DgAJw6eLjdnCyT4/ed9IaeYfYP5iPtguUGmnZk1I7uu0E
5Bw0nvAA2kodHHD4UoOhFGs+9d78sFuBN6RedPcp7WEOiPhgQtrcLKU5Z+s7OJ7G
T2xwiNbV/juV3r3Tvlml8+OfNWTYnCAkEHtmZn6OQ3bovwqjqEUAh0ZO2AZVtvHH
60XUXmj+WBo0byjUAobhRP9y/YGhA2CGZTzPaPCC8GT/+vNKafJut9R3aUKvYhSg
SjcZHek1PO9T7QqSGGqOa/ccASPjq4MSXdjHI1odfZYdx/4jO/p4XQ39iMxIU8IH
iSCjJi6zBqs8etFNKOpI0RfJ+QX7speZG4bhLiX+eZXnTsEpsizwvP25u+dkEQMf
mrlnO3n2LwnyvM52V7aoMnCoteJjuWX4S0RHg7CM4lC7k4qHCkFiKsaaKV25VxDC
MqmFQjDZLkWdDSr0o4DVusQqeB0MFEMUcV9uITsZ2SETzbmM/qCQu6STw4SFmBbg
rVOSMM2zVtzK1MANi8yF1LuIFjM6zmK5R8tdY/+LqdYp34kNLDcINAxvZlc9h34V
2hBRAUkABVuvMMLAoRWaPtWSuZ1jTSxCQFVIlDHm0A3Qk9OGx2fzrFbF/d4pdqBM
QMuVw8fDLweNmmpDRxkJ8oLyOgQpl+zn+1sJAKevO+npcxtsxBXPPQ3cpaA42PPu
ft1iuEtu5Mm54/9rwG94T64iqrzZLVKkj99Ljko8L4aWX8VMW7anUwbvA+Aa+ESg
kpgCIdlxWnHC0YcuPsHFKUnRM6ls1KqF7xYT4kkZE35YKsOtyY02pLF6GZV9bCJN
vusoSAM0JRD4a6FoD5PweGW5JkBSKpJx/t4UQfVCKILEorS6gVU3uIoQk3b4QlXM
j+/eZ5ZgrgY/g+tgs02iAjUBP9vKzs0aNSSDaYxDTel+cj3whKkd/U/2lxMxOvaa
cI+F0w38S3Il2xyNjmgGJglfddMWGSpV3Qv9s9iQw2L940mNlBskvGeO7mUJDj3I
QmfUHmSibyTnm8JRK20LQe/cDGX3gJhk5sMMsLQdZFaMQHXpv4fBBKw9ne78MIB8
Q4OnyTZl8lv+QNo9yepkZtyQIQblXruYXQmhOtdEvIZrJpTHzOzqgyqAp9vGD8aF
1a26NoaRjnZ1OQlHjCkK9K/5LYzPYJ4Z4TN8ydytzp/6BmbZGx0bC2EWTrYRQnUY
K4SjIZXL/0NqLTNoRBYFzOa55/j++MgobDRjETRKgjwBvK+m/gyMoOfR1P1Z2EFE
OU3I4Vj+hPbjVbUo2HYI+w7wwmilv+E5N1EoH1b805SVib9xZatcdc0HW+nPKdmx
meD0LMjl5d4PRaH2C8zlXJl3N7CsLX+D1VEO2OAvW/pxXr5zb8WAWMI0xk6vnHW0
G43uy7PSf/AwP9RecyPafwQA6fIx+EigJ5fuAj9sS5alqMUPN3z2uf7+cL3Am15h
ay12Vvs3BX2tqNPKOe17BQ3GpsscRBbF8wRrgJWubGJ2naLbaZJYR1bt8IK3ik8J
fMAXS6MP5B80CxXE6VhjmZhBpcmfBoHTVZrTeXCijmiq66SR3RccS/ZAwk34iAap
hICK+FUW0Ou/Tyl0c6wg5CF7J62bKkEu51WkwuYfBBkNbPyXvMnuuRnSChYP6Mc2
5EYZbtO3+6NpYKY5J1a5MLidhsHyqLE602AxHKZxjUAaZWfl32ifTtTk0QfUuVjU
V20m+8HGfveEAUbPWTo0ehNl+Zpd08z8c9jqna1YGkafrvo/x2uh1X3dfavgqarZ
fsRw7byWuPoGQyF3rDvpMzxVfbLqEMd+NszmpjUcCXLj9hEiL7eRMgbiFyzqkqNe
o+3paT5Ke25rE5ucxaENNVTUOHzJQDdQWx6jP5ReJxGLYIJwuQWjjg/cf7PAnqJH
dLYJ1z8RGY7ePvm2XJ8py8nyQQsd34oH3eMi8Zh0V5y+sABQurYPtnhoH9RfRe6f
GVghyTP7uUI7dKLUPK/lvVTyN1/OWfRGOY+nGmnn/fYIL41khJf6TpbgNijTsHKQ
GgoQqgt5BWFDNEmFvOEmOO0iOkWgzkgjuH4YhKqVDIFL+mmmh6yHW05efko0YoVg
ZRX/3t/3VfnGmgoPF1FAmRvJWY4zX25in06svU9tv//kXVy3T9ERWY9LSfN6Z/qD
12lscDpsph2rgWcfHuKuFGhQAQt/uZ7xC99MYYkcGqxzQbrJ1W7JQnI5y1O3TEX/
SOLF/JXxpRet1AoB8YYb/SkqcAlplmn3q5sllbKqZF3fsyrGt5AJ+HeHY/fkoU3n
kgjAjfQBb92cYx2jy+uwHBSGG5H6ZEBOZqULOZDP/UJjnqSbeh3MS+ZCWxpNnpYy
teb83BztCS0fjvNPEsrb38Kmir8NW5mhcINfVjpJmw5VHUXnyPBtNeo83os8bEeN
zF8+/VbY/DxGUl2ffr10iqnaNPFlOcXRsTrQJ5yIGTGyfA7b2hQ15I6ia6HKTvSy
4U7rIZw9AP/s+7JT6M9NDrKHmx6iKa/nNHHIUWYPB742N6uj4JjcderksypHX90D
mMdwt0rqoJ1ajmEnzMJ1C+UVJAY93KaIsO++RRMs4Ngr2nSsZRnLDn4yL/ghYgX1
P9VDfAD7AulIZe1jDWV6ERfMFbbu9ouMkSb43cmeW3pECYCAAbhZt5lG0qnPvHbI
wzXeoAptK5OAqWjvItWF6Y78rey0oiVbwontpEDX68YINylAJw368tOAEZaMyTYw
GUt6is0F243wzd1VZYMS4FqzAEs30dNAHmXdfee4eMWDWo+tjT0n750REuRy006s
aJth5kHJ9DV2fCfPBhmKW42hsm0tCstOLf+OtiXPF8LLI9Gk201K1z/xwIO8Vpwd
DHpaH4qbc0NTtWamNyaCZcUYp5Jn5QvJwAI+P0k3TuuvBVE4gVMCpsotzIBphs2x
OkgDzy9YGqXDtLW7vu+72IFFXiSCI/DaocOSCpxEgPOFW95to806UtwKCgMjAIsC
7BTiRaCSUK4RnIqjil7JDpAMaoL+xL/00hds0DL9UIOLPui3BHJwS9m2E5xheuEA
CefOPB/4nwN7XE95W0skQbrMyjhMgmKmFU48Yi2TFtsO3wfbZ3BwuJqzfNIKx9kw
1gHJkXNvBfjQC2IExivdkZOgorWivq6dZNhdJ73METZ/WVIlWkCGHDdrFYwUdG1q
Slaaa1VHEIKpWJKS5l7axmD55hBha9FtOzJDP26ibr0SgONDQQ7ikiUIgW6I5h1Q
FvDDjSvMAqfp+SuFIAE2EyYgMz6Uf11K7G4YRMfTYBzICzsksGDFPneJrSey0WiR
A41YkUI69053ebdo3tf0cYun264ldFs14rw9kj/cgwZEVZYCsyiP+pKAbfx9wbzn
jNswetLpqYLlm0YIRqpy7kqr6aX2n8OSAd2UeA/WiehfkoEGHxGzG6s5VycOIV72
/MZMOmxFk+ALqLUqnwrD68vY2uExFnrvQqcxXePPmfLH4L9NhomnzIjYJB9Ud82+
h0iK+EiTXWmRsanvoncQEJalv49k74F/9kFjw7tuQ0CFrDN+e4bsOkLHunBFKElp
Mg4nWT99NpMqKwUxfHSYQmBPhcugf9eVJfKZeyKG3fFxpfhGRXvm9oGkNmD3sXcM
N3tR1HVI+KR90z0ZS5v9C2VO1CoAAvVqWE7C/q0QYSbhXVORc4/EdD4aQicqVlQ/
KTcBkC1DVlfMzCt62ShpkTmJq9L5N86KVwT9MdRGHfPzyYvyrogwM5clAo/c7HIf
8nVxmRGagu6+3ekedRFPK2EbYBOJwZgpPq2cmln/XGzdfTIN6d11cOBIQhC1qk73
Q3wC1Ymf/C9AUj+bAHOj01LTs0PqRYJZxFFeRBLHhXWvu4K1FC6N66eJ21OUfAR2
tJTpY1GPHLpSauLMKvhDrJypROZO5AYTO9DVur5Ia7qZoF/zc6/ylnEeUEzGTCiI
1CfzEwpxkTwPUj2P6Pafvt80svQhVuJRllWfJFxYiMDdslnFlH2+iblJPHLp9kj/
0w/Idgp9EO8qN9fcaT5CK25lOJOqfXg7xKUYdm7RfNGP/Qk2eUjwVkTaIlk5kbQM
W3RpP+A9CR4HF1X6uTKDWE+d9HYav+FMxkd7frV3Fs6cCUddHUuDzgzZFLH3dLP9
9ealL3w8kDyxIaQ3FaLd968BISkUOdU4K4jEFj4q6teA/NGUL8KjrEiRyXsTxZJt
CN5ZIImV5JUvZzcYnt4gpuZQ3sHiXLm7HQX9DVu0NQeqZd6S7oeTmQtUWODXa7Ew
JDF/XJv7VRTuLPYPjDkRu8iUiGM0AmPQpnnEGsnW0Ftpu2/YPJOFQYU50I8zGi6j
XD/ko3pCDbRZG4D3EbaWED/lVTPA2E2hKSHwoWttxPTH7lRU/56qKi8JVRH5dUDA
mFuvolXZKUrqP/CRkQ5He/pelUBFvmiF3VFyKPOwP4twfB6dythyV0InOrYnjPOP
1vj/xWmH+bXQmrgrd3HQLk6aJmMNqSFm7y6BDqkdo9DM6ViKebF6bSA4L9t6kWBI
8dfF6Y6QJq0eIF09HxW6OGPlalmea1baqcv1SSaPHImH7fnnwIwyZcELsQgmlhJ6
fd01lk/RHOzADqXOfy9wYGP+zN9+NQ6rZY+tRByeAjcuXhlsK1U2c0GhIwrbCw3D
1S4Wi7xvrnu0aFWeUNgahSXIn5CC16yqydUF4ARqvFK61wNrRFJziYNa1drfJyPF
UxErs+NHhrzfp0gptwqej/fXU+xcOPByuK0T9mQ7yQUbe9MJJrxJazeWHR46nEr+
i/iQpFwU6WGfG7qv7RjH1fYHE3htF93eK9bCU2LNQ3OWuDdrt6xgDHOCzzu4YExp
MdmIQR3iMXa3M3FiI5zBZHtYL/sMju8qsFWQUCpfXjXEafBtUZtg19PRBUvyMqYt
rQRZNI6X9odBpNmhbY08cEpV2HkneCidmbW1PLOAoH4Wui5U8s2D3ixt4Gb7dMwt
ssZUucOZrLsKFe4zezTYIlez+m95XHXHRDWbbbbfmWO6XfLoNn6CIx2dcqLfWDC7
9MpambahqGS4s1gktWRvWhTEgzTol8uPuAff/Qjghc6Anpc+vp1G7cLjoBcFiO9i
Bmz91nLLlncZw8WLVNAqUsQjlQfaT7Y1uGKmZA9bhEaxTJX6eCV3CoOXVKBTqAM3
HB1mNSXayoiYWx1xeAAjgzMSKLgjum+YvFi1M7M7DZQF292lLAmV3Yhhm6RyBkVc
053+wAfDScSXSJ9+LXVlRGmD8+9rCrzKYO3qz/+22m3tu+XuCLbLVieCf3u8xqcd
JXWVmPs5c+C2Jgmmi9U1WbHJyyUna6U3gf3jAkoBZqu562e+SKrZ2woxbT3gXz1I
zPjxVZGPIt2cjzGwSQuGUQEIe9YtV9nqQTL6HDNIJ9e5G/AWfLGXH2ywYGHm7LBm
jZYGz8wu8sl8hcY6rBbHXuI8vMq+iTeofhlS1VXYvGjBQdAuAubwAlXCCDtLe7UW
KHGJ3ai6IC5o+ydWJ/KFKlRZC6XDthvQWcJnsGUBDGFlorYAFfyw1LcOxIkijxfb
c+q5T1f4uKD92voJ2/dlZX/2P1KyxmPHUwd0nk7vkA6G+E9t0EoMN/bMgW84sOXo
A0b71NnJLQo5duinE9cbpMti38nh3Q9G3sjKLETDhgg8PSJW9WK4sCKcqcS5l4K3
iln15pAVyGIouQy6Toap6WCSjY/wZD8Sjp6z+ifNkp/ZG7a4A0sLbEE6VYKCdsjz
uC+bYZBYFbj9ZebJvSHTCtXvN8RzfT4ep01RohIaLKcLSMnDXAX9WXtcGq5gux4s
g074+K19ke1DPNYwG/4TmfSBt0dNDLrWt7sCLTlsvKpurmSmsVmyYUWk+2gMdoD1
maFwrdisJZgyeNYUc7pgWogiv2PeoW3Lw/1w+QVxU8GUDkdrADSwt6jTnTT7xRap
hcmEOnWXT+PLA2euh3aWj0blRF2G1fzu9NPTaloSlLKEJUgXk8tYsu3rf7xzuInF
qFUR/bAKfEsXzu4LAAzPOh6Uli+rI3OyPkEpNDp/ztn04+oa+3+n2gAmnQeREOTQ
YmG4PyEwBTgW79eAaNG61T7CPYu65uqttDiUV2Ymcg70l1RaFqOkuN8bjd8tSNeF
wvUT3copQ/EhwjmBN7LtOe8Tw4SKQByLKx06mkD2+pMTFgAahKIk9fJuBs+SRyfd
HRZ4OcaG+1D7iLeZHgGffXwbZRNIBs9wwkaRSyE3iKiMeOWpWnJON3HG392dj8J1
c2TTxQqTV4HbM4ErUffoO1TWdNOHOv7VL1aOf/nwZ6C34RMZtN/a+ciOBIwhmvQa
9m4vmtiO6XSGnoRAc/WxolvbMRhizKZNk1GFe98M+I2pufm1fbUmzWVnHXX3yL/N
S5FjMMn1mzOm9aRSjeNgTcMAMeNOObxgSEtO0v1eIZZa+w13I0p5AAeDNylXm8DD
BB5yVo9DKYsHeAHK8wCFIfHBOZgip2QutI3N2RKFduIzAY5Q1a9uBNXB1ftOQzY+
3riWhaw/TploREC8IJZXP2MhB2ufIc3wSJX5waAUChXYKuuW0/i6t55SzUYjWOAG
/0Hakk3Ahbmw8dffPMNeM5TiTHed1Xme1zWkCqKS46ZnNestkwJrNEaBfIa5utiM
vugG+aghjqr/gkKcgWyEl4hDifD6M1uM3sZgILS+Na6Bh2ncACOnwwmtXFsjrmwz
bPXKA7DDs4htXfXDW1uWOIu7H4T9kaAIQVoGnsq6gywibJ/VLhafPQAI93dbDWBC
A9Rt6prGCDCZ3cvD4jmxzhrS+FOt/gD4qD6jLOVbExwjPZZEybolT1dRbdeV2ikY
teiOafquVvrGfHqquk5t4lf4SgT9sjrfX77SVGpG0G6XOMaasO/e3HiJ51bmU78r
moLPAGi/AznrQ7908+zVU0WebfSxJULyTT8D3Ask5uCUOEH5M07EZs0Idx3hVuiV
/WmkD6k/5ujtgMnMwLzdRfoI7E5vDpKrjcLgNkzDOfpg9LJLJgGQurh9wqtUOi+q
BmrZhJd6KfeiZ8ExUi5uJr1WWWlQBBOoz3yYrCPxQP9rfyDnQRSdbwqGTEDbGK6i
9Q3Ro2WHNKy3w3Ipxx8CJHr2ZtPuTEv63IAP6i9/X0GMUlHZ8zm5c8XF7CT+8p2O
ryoI6nb3WpFoxgcTtiW0u0rBvtIutmFKFEbhzE2I8gbe4VPCMS9bWz/1J9WVSy6a
IzFiCgmZdzxzQazvYegfcPYX67BGU5Kl7EK5o6tkBR+Qqwa70bAFP1vDQwaKzovk
u/ucdGMfPAfIy0rqWmwEH6hUYTVjLLrvWcFzukdMvL5pekyes1lLjvoyva6Zawcu
XVDntaBMm3OzWeKhIAY/4/BZWv/OJ0ycjoxvMtPuV+w0JuLYITY9SNEnMISDyJJD
k1Bz0Ea7Bxu3n+JcwSDn40dE8Olkox3Uk1z3HPeQnG8a6mUBKzVxOM2qLlUh/Vyf
1dFDIOZkpGGFgrI/XQJpfV/+TgX/mwK2qyS9YyLCUZCB+6tAtzUXLvQo9AhRwAgA
i75v7bl/HpH80fkNKQV/aKT3P6oVZiw2vs4yRuRxGQRSM/o9dFi8BZ3RxGxpG+SJ
9Jd0RcHTSEyCAvczKNpQgwtCHaFp8ss6L/qGvmKiJCYuhLGQuyTBTovCCjY1f8oY
IlG5xvrUiqmFeiXIWW+LBdnxRs9s/TQZ3AqOBLpYfmKsZ5Vcv2F4mjt1idERebg1
nFe/1Ngnbz8PtOxDjvVI08Z6ZZ++uXb84As7h8aZV/nMFXHskmiRQjEIfAOcITWQ
4bASzUugWvH60Sr5LalvjlLLxLQaiUq/eHUJcaFWJUKFeErbr5+d3U+10sON0ctq
klczIc54dmJJEu4B6ywsZnhCruo9UMrHDxCgSRhFbCL9LiHikTZWHuH2djz7WJfO
7yO3IIaKWjg3GTRLJp4vKH4FWkaQlFN68PHg2z1dgvPKyYLcFTCMLjZtLzkDvhaI
0hSNgWqLIJuXiyCMtAJ0apzVqIODH9wF+bVSo2nIGCS5sNwXFge4QhSMi+HX5D9r
5KVUabRqt2/b7VIzDjqvQsBeA+Vz1D7MpXxeEiO6IG5EJbcN9jPI6QQL8Uu1YcUj
QWdOjfsj1d54tNQGLOtHxvQMG/c5HBtEOdqSLNlaP8UE7zA6pv5gvahAukKAY91e
G9iIgC0aYYDbENCrK5AAIlifTuG34u3ZX6vewO9pnKA2SBp5te5EAGl797QMnnkg
nQQbCeXY4btD+NpT8JTHlPmi7dFXfsyuD4MiOfbIBZIpKFRpWyBxUO3iWrO7gJql
d+QzP7RnC3UJRgXC2TKBj1NRdym1utO7HfowaBr1HYLeS/LemtonEpmO+ogJyjCA
5FDanGzD19lvGpztTVc123p0nC3DqxnBuTCcv+xOoB4nbDI2EQbS9CF9MnSXJzpq
8XsptiVSof1wyniUO+mYadH6KbIkzav/OdutRcEM/Fbp4TFe+SQho74lHQghEziX
C/u3SKeXJr8Oq57RSzdhIvTsecXRzwyKlmkBNtIZ2/xInOMkKz3A2STOtZZTUzM/
7mQRioCRDkO8HUoWZWRFJoMcViiGB1+YjNXG+8ALrO/Rtv67JLZO9SeYmtyq+Kwu
nnc4jgo2hjAAbXqTDWEPz0P58wVhOW1Gw37Dhg4WYC+BY/DhLOCLaYqUEecZkYll
+W9DZhMpy6sY5moBo/GlOUwwoYTEiSHqhQZNl/b91WnRyu7qwe20IDi1o7V+xfiq
Lzm9pL8X9SoxkKqMLcj/u6r0968JNTu2fmHa22hLwVgWyyOxS5hOh/xqL9CDWhM6
45KBzg7c0b895f1sX1E+hajkpgOpvF57NEuTNikKx1h4e7AV+ZmHe6ZhnW6lbSve
QCBZ32B+DhBIvyho5hVc68sXt19sbBlqIarilLB20k17vVj7je7D5IutuIo1TJls
YCTLvvwFd7V0l/ZwTNgRxzNsrgmI9Qu8+mQFi1g4pgppVGqPQBJ43312yKlqp/0L
Ua48ZoTOcbNQQPv4bf+7WLep6ykjv4dUzIh6/alTOTpa2eIm6A8JMhIFIPdF3M9d
eb0P7JTkdkG/zMSY95/PZCbwrob6t6Djg5o1EPkhLSV92oj4dAkz6HMyc03XZxWJ
xV76CNUgiZ0rtuV1+qHJ21rXDXvDuiN64w5HfgOZNzWjdbQiRJWL1nl+bGz+BnB7
4jW2O44ecZCxH01E+GejVQWx86n6vywuf2Pk7kTON67E3FJ38jAF2UFOBqJyD0gr
qVmVj5zHD2jyPNMV8DVEZIO9JfMKhN7D+n4BkSG/QdQmEiis+O1jBHBksurhShVp
xokBr9NkEG/VgKrk/IfSJ7DYjI5HeZzVvsqNGanrgO26+cpcIPtTFh+q7p94iKn+
4cb2FHMdpzDNB8WrEfoKn8xh2WhfaURdiL68CuuunucJPBTwvuu41TX1Py9aRGKT
WbXu0XkmSUS2RpVXBvxAKsQTXDo10HK6SD40f8/QORfCi6B1lyWFugMBaiYOkRqw
aXNCxJVaHcuhJASCAIndD1BBwUSJXcwWNwfp0xYKXqoubbUpdO9J+4TeDEGMkgMH
Lhn0y/f2qv2DRDPfpfGSM4BAc8qkQTrh0oJ2VoNNLvJCn55H6oDMkAoLntVf/emF
Aa53u1xxhiWjpDBj8sthDI1r9IThHtZRDVqBijIU8k3dZoAH5uYE3NulGZVLsk7I
jD7NUrApsWQh1ddJ/4/otTHkxRCzENz8/y2aJAGZ6nwSANRnlwzz1CJCfe+aUgh/
Us/7nimjDS0s1fRysVqlkJIqKghFedKESNfzrMIaGMjjxs0yXQDIoL2eWknXuPG2
uWv8B9qFHrFKk8irlLzRZPRQGGNPXTNvOtPxr4hdd9OuTmW94oKSpVOmN/33jpT0
iDGr/IT0jntcLBIIXo3/fpHZRxdHLPP/8GmNIRTGw6Y5UsG3+JOE0CGFTJe4nwy9
OD0wt9LzjQAlTDqjjN2VgdOqr0ShfPCoPspppwpqVwlgNHcaJs0dzchHGQF0rWUz
9cp9mz3t2nF/oJSdOlxa3ki1g2qLva4gT8IkK2BWmdIBEsg3T4HFUbWXVzU9W+5L
jLVgrnRwnH+d0W7wMl+CoQi/6asftebMsZ3Zq7h+PJYkSHuR/7XOQ4KeYI2ZG3r/
9cUT1M4Vip1bjuDPw+uQhRtLWSH3LUiLk/fXGSxyOM2X2lHt/9mxqv9b4LhjyZqL
RatTGb7KzmkQOV2MGusbneboRkoxsuw+RV8OFmoLx52eKl5PjQKGsfKAv3ENVB9/
Alu7QoKmgBxP2OEkzeQY+OLfs81U10+9F6mxAeTFYSXZaUb0/N4VfCWbB5MnkFVx
tgocSHVeD7QM5SoanhEQy3d4VO7sulI86pixK3PNA4SV2dSt0/LtFrakSgXO2z0I
hBeEC71ZDR4Zu9dvRbpro+RRrsbfZfu4q01oDcwxj2/tDB/fVMWxuMipNzIXxBT+
ysA34MASoT70gJ2dxq6JZIQR54gffW+uZ/dvY6yctfqR4HETEMJGzIDsIRls71Ac
MGyevr1PK4jdKviieDcutAyk4oqIjMmJezOfT14vH13e03aHTSKSAMoQIQyzl5LL
HengLIynt2mQMzZO4DatkjpVeF/P7znM0AFW2I/aKhJMh4MRMaIQC6ZScgIqpgU3
uhfNa1CEZcARHOx4bQ6SxbiEQ0mPTdqbSR5vZN7sevV20OmqyxqGzsf3nDe9Ccvl
NO06nVewffDLBaBNgKE2voJKfr7bTK1ytRHFz5Uf6CsBpVsmxa1+FHT0P7EKPFb8
TeQwoxnTG1CC3LBC+Mu/2Ol5eVMjWFf8JEz+0GvAhJ5Jn5HNBzcLaESqgKKlRQI0
H4hTjC5/s9evoBrBxo00vkLRt5GNXeZOTi+rNdh7GYoP4dOQKlWU9p9tJu1oP+n3
jN6DGiI5jHVFb+gQ/ZQjN+NxNPlQEf6dTK9/bEkaek2qcjv0kCEvYpuXYdK71w5Q
/f37HmmvIcDLfZVWwS5Z3hS+FvUT0q/iGApl4RsHlnd73KP9Ep9nfriAC5alzMYt
Ksc0StWy5OOc6OcEOHcqz/isalZ1jNeVZ8A92XsvLs9ZuyMRUYXFfWypwRsQjAQS
dICchC9IItIOryRPHHp+QTaLH+dvScS3DZsBsZ5cBHuk6s7s1bXuoFETEDEIaqFL
F+jz5jpi94fbEa7is49Q7HtJQ6wmQ683yNUH2dldujUY10T0fnt6WajcA02txI19
IcSHEJdvPpA6AIj91XgTM0Ib7m2Q3bGkfg7BuOWTuVHIwssciG33mzU2JJqRuw7f
yk4V0QPa417GziCjbC+Xfkin9qHWpp/V5b/H1G8qVKTQMuWkaokbQRni5c1Rha6R
iwedDBTzqWzTBNI+boXw54Q1DDVMnNOUMMcQBoeKVTLFv1Po+pp3MNXYnJPMFnu5
PDRls0RCm8xdsV7ikP8Cc3cpMt9ViIeluxy0j+Jjw3s5tfAFXuKHadBFh8IzT4c/
rHwxQYGQ/nd/MycpWvwRe9IKI0TIpi7VBFd8Hn0j9BKMFAFMAhQ/xmgiMk2IlLs9
9kbbpdWUMjHa/WI23C5bwQb/iEpl+1UBiIb8UeUIE6JcUaYD05bEvGDEz2tKg5hq
3vF15zmrSe9wR4AK7ewUIAB9ev9HY4YSLKNHs/ut4KDr9oKMcIYfqcpxjuGT6G2P
n29rjrXegKlPoC17B3t2Xl2W3VQY70XEk9+ziEXqnNPrJ3MO3NjUBud4UwJJS/H7
knUaCuOXyuExodEi6roGRllDbGOJTDiRpD7NNLhPY8XwZlGB6A//Egc1si+osllE
61cAuAe8hZpJqftQwReLcYFtc+9ffejH7fQ0clW8zLPs3FdENofdBBlxmEs4CTVr
GdDTT9PgbEiHa52efhfcnX/0MQUaynYPRGiIiyrI/SVhl64mMPDKbABYuGHAYzcZ
7bT4VyeI6mPvfP7dUvSMYjWu3BxPWDP2se70RFc/siuWxBA7e7ekVQym0rNnABTj
HccuJK7MhHwy2h6iJJww3P3Mu2iaH52fH45QDmJNZQ2sGcdFLgX6NmNLbjkIgLJm
Qd3nasEZjLZIm5U6TGt1WS96nON0sdndMzKu+xXhqtspUDF/i4ohGZhkMpDEBJmS
/Crt1YXlaGCHcteKQV0LW/jfl4dP2DQ7B+eHDhoohYgJ7Pv1rFv9N+iEaFeuhX39
IBZnQNktZSznLdZK+cZ9jqZCh0L0Elzabs0j+HUNVrq3K+j/d+2hbuGTpal1PG23
Rv2QU2bBVnQ410S2ce88z5nudgrT7YdiNwEVrT+qoiSRErzdH7iVpyWHpRVdASiM
wHAgAn9OPFCIZCCojW6PdK+alPooddhPQ9qSNeZmrdISh+Y2QV0uXVSP2WRtzKt0
VrGUbrEOW2Sq2FtFmKuywqncW8I7I3JqEfwlhRC1LLlAj5bx9uD7crdfbMLV2wXi
Gg1NQ6D3gKjlK6kBKMJ8qFWZtb1sEvr/WVrHGQTaAvrzhBC6UYu1Vmomfbnbu6ur
GOIfXv+lsDgBsFVnur+LQhv9Eji7IVLY1bK7SN9w5yq9kyHoW/E8DL0UJQUfHAhy
xIkYgxTE2v+206s3pM3x4Tsn2uYRC+ygRSddEf6W8E5xuJopCqAYZyqZwWpJi5jC
8n37bP9gaxFzXe7aHxL8Zm582X0+hLkEfNwWwPtOhPtgI1ySHOmyuOcIhv1P4Oa+
wcYE5OqPf7t7mdcm2g1RAZ3IgAsGXWJbHW9pBbTFlMhd1i66qQ7lG+KH1GpE8udG
GRhpAU4MHrznqYOTcg4GC1xTEGxdlBpJMgFi+TkA1ed2cqsUkg6+KBWyNXRYU/AD
u6h60Oq8YTj3K7sPaetUmj7XtyA9QVBc/Eenjqb3mFYXIeB8EVVkRBmCtEuokJ2n
As/ofHuH2Y8dOP24MQ8VU0udRZc7pUg8gqIIK3xw7VCdqA3FFz2ygyD/oqJ1Zjxf
/kbp710l9iLl9d2cOgqa6K5Sd3AgF7MmNIxHKtt8dJXp0n5IlDRXYHvlgYPRVoc6
n9ZmjSNhFtT58wkQFZt3zzd1JQopwtejrc/40j9ZRyUPh89/EBSEIAN2ly0K6UWg
UIHcvEPGpqwusD7L0tV43qJ/rDJWTrvSUVWMmRqoO8ILrkawMbZcUE3cqMSKJweB
4VZVroZWDamMKZwhrvxqhVbTu2/HsWPxS+dYJpdpLHdSBv9MtglAMhS37cvV9rZc
mej+zfYbpA8SbSvj6f3AqUNN0P8QjrTGZ2+ClRI4VeDvgYTahS2ymsHfB5dn7xhH
hUAUblXmCM7DnWWDVLq1iwngBw3HtDUTOAI7Mn8oaD87UXap+g9Fxd1qRtrVuONC
N3/TTwmp4zZYzcoiRmfkkb8eziqIJrhvfaJheR4P3mlVaYwN3a82nFJRweFjdmCa
iLTWeanUKLCNjXhvzPVl3FCUN8UA7TQr1dpd/I4Ml04QiECORoekntsl01x9jKOL
FFL+8LMkUFZ+Ayos11VVV+AinAoLoV0tWfzctB8Qiz+XfK3gCn5bHtv36HcSWPI+
+/3ycQoIQBiPBNpIFw/hlDJYQujK0D8K3aT8e43J0C4yEtDpU9u5OiKUNZwXsm7v
iVtnjNbaNcon+V+P+ymAC+Ads+shXhrhqp6i6U84LQNiCpDi9x5TXcvrBTnGA2II
D87xD518+1IS710A30/hD3ipGS8Ks/kSMwgIYP9EEAyqvbWX8JqTesV/SAKOFATw
xn+8LpmWz4YqcUROj96lhCrwo/5/EMq8A4FUZnUQwenb5N1x070+mMQ/6WD53CdV
wIgOHYE6hI4lV2P5BSJLuKJ2Kt897GSOJjBjRl5TGg0lu/9VMrqc/vTUShfj1ITj
PJF8bQ3VZiXFIN1PmjwbHlrd0hqFrCbAe3DCYvy7+2+Rc55dEhfB08ktIaEQhNVP
ykf6wrGsFGCj63uJ/xkVHGgbc+kUfaBtcXtQ3zWZ6Ik2bp05JdwbolInQ0a/xTVe
2JdMivKtrfwE02IGiU7J0aYgd0PyfTT5fnrbukSN3dnvoyXdlYfEaEPJilbiP26t
BqZX0lR2jU8ol/+i9UaHiy7xcTwp4zO+ZC5w0PNDhGD2fnfcKe77+qJnalDMNx81
TtT2v0B9h74FV6u1JeH2xalkB3pyQdBqytuv0yzxYznWslQ9ztzcCFyCtVgvXvgr
QTssMeoSt+Q7lBqYb1PRzMAYOUQIghdnpt8j4nfiIAV06RV/+467GYTabRutpwFt
KMGuvkPCM1wjsppSbp8qpGkedDZ14zx3yQxVBokZ/1lY+m5rNXpb8q4tgyd0Rtdn
iCkQiOXPMt88Z9BObWfl5Jyq8mPGuxrXuAzA/UXS7HYxZt+CeHtupEI3XJ1dgaV/
ww0yOOedfmX/BtCH3FV/kbc+JiwFtFtoNdNdkomm43kThr5FrUUxAVhpHlliC2Qd
j5pBrLgVPWfjlZ1QqRnPyFVFbUdkK3h07SDl2cRhUDANmqtfBHPRjpXz7E1OMgHC
x6XJkFGL5v2QzdvwOAfSJMz4Tvj00grNGl4kv/92orNyR9YYUo7yZEl9n+6gp4yY
+xRqpfsR44A7F0u2QuMjU38WqHo4zQXVkMKvfFiA2lBMM/hQ6LffVkCBG+ckWJbv
A/KDDcIJQYcEsM9HPQVDRamj849QfwoJ4B4onlNguTtm380CqucFJJkb2HEQdCPk
iTP52eX+lCbz9558l96JGlZ8v30l0mECim8Jk+HYa0k64hfOxIkltfVENqS8uFuH
QHtN/6oFyApI8D07yKni3xrLqS4Ex1dahBCQ6fthg6Lv99rnnE7EHokn5a0Zc99u
aSB6595BMxvKiShQnEBDJYTcGg3t+fLGsxFEqn07p0mIziNKwE0pBeMAxmJfD0BM
674pWZnVhFVnfG4D8+Y/Fsp//yqoq7zotP2KK5g3WOUyEqB+wvqg+msRzlu7iRNT
/V4vB6DaXsFi2llOr0NOstuSfJCz+SbBZ3SmC4U1ktPvtBv0CECrxoQUIYe7GTFc
ZpoIhKN8nZ41DfudGGBZK01BEhbNqsgvc3SiKA3Zgp4+qABrE1mZv1DPpnwAxoGG
l3QpbPxCID4rRQ6sPMZr3RBcuMIGM+oHIoQ8bNKzE9JJZjqH/r59qIgabU33w4bw
Ylhm1SzWPW/g5p6WDm473V9ykURPWmm7yvipdshoncdHVO+IpyhPeMD3x+E5xRQ0
Y2KBb9+IIB/WVOUvOc7TkOU0ZW71AMicpXL9KUeEioou+xnE6LdVBV2ZxyZuWo2t
omwb4yzZRwvSDjWWWn1acwKWc009mjVrdMnL1rlpcquLvdAuRZ4qgx9hb8DPYAkt
YnrQA8yL/l45wLbpNb8OzdZwKHz5UULZwpwHf6RY6xJp8V8okcu0PFbzsR+EblT7
xcMSj0fhXVSGh74QcaInSPamSY9HpdJE7pYN7+E7WyJ1C5ugxVXu5lDZqYeqKY83
kidt4OfNKFTqiiDtpa6lFtC7ZVhlh3msgF870tHRzkzj5yN1+WzoBtjfwz+AthyI
2kgkok8W08WcugCTBiQgw0jid+zp1dwh53zhzXcss8k8JzzLUx45cLXZniyITawS
yY4r5wPwBGGT6oMsnJGU6zu18yiCBbJuSRPXtvEHqu48bCn4efk1suxMF8G9/R/A
Qu2GQG80aAiXyau8M1o6F7IgvAJ6jQ+IVBAT8rdWlQB965F4y0M7WxFXwK2UBW4T
HUvvDr6NSDh9g8eZQvoWnR/IoqSCCgXBX0hjsHO0vmgyyjQ1EZauj5HZnLwOo+ig
uNVKY4BI04GIY1cHwjJPKMij/fRpSh1iiHT0YPG14LLVtpG/GgQBvf3s18WFn2ry
dI1RZfLEczih1GsVcS9Lu7OaFxvfolb9jqATFtlZqN/mt94OYjmsOJ1xOa6nlTtw
rXaMcWwmuF8cZmhcQriVL/xoqiQfB6x2omrGKgFxFQrQa4xqYb72dqpkqGAxxoFg
7Rnue6CwjfTsoeWhg6NYLp70dTdoLTL3X7WkyT2UR7sdMFBlIOm0ANMXhTEoaBJr
Q6h3RtEmMA+ameFFH41A5Zy4GZqLq+uCajCoozJ3Nw8YMVTsUYV/DK9d6Tezxz1e
LpXtgkwGXghIKY7eWfnqsmHsTtJWAgwTk0igXluiuw2xQMQaa35WFMkBkah5NEal
Rlj+109u8JmCglGSSUw9zChuE+g+jIzyMVFpNjmB9iBksSeJQJ4gTylVcWcexg7C
TYp0g47GecsfCpfxTQg+ei5X6e1XygrUu4iX4czJ5Ctz9VozUSyQZFewepHie1sy
4H4yTzx3b1gxTpWlwdIOSQHLBc0a+QtertVa0sTi1QGoZfuTxu2TeZFHsvblK3E4
FoGO9uZPtIFbxBktbK0lCfTOxNCmIas+4GsFzWYjwMlhhde9TucE571tW30WsikL
ZPG4TgXE4RBs8uzzvjeEvmGJNBAGHwGjPDgyyZyTEtFDRfd8tTNkA7EJrp5uPnVA
Y/XVw+RKKBImp1FBhWIf3DGysxR7C6ggPvVBAGQMes+gxaehKd0WZgrUl1caDT/1
SXJrVqFDQoRs9XFxR6Lhuipx8DIhgQ/9OHG7lqRsk3m7PqUGrfWEvBOTFCxGU6VW
bpmlcE/0rLmK7kWBEBaXIMHSBEMN4kdcxliRfP1/O1soJCwWIrNxqTzZ1TqbjkPW
cLp6JujVM5/rmFHxJRYYcbg26szzzbe2pak2lLOMQHvWFselF1ka6GVmTesZGq5n
5WTq6NdlPtAz/dENw7RAOYyEByMaUVnP2+cnEaJa7RKq1fYVNjgnN+fpQHfNazvF
lXI1vrmATrG6uhLSCazVH2flFE6j2bpdi39MWi7Z72LW6gBvHuvqWvYWxTHGBjSm
LrWMCoDG9O8IoMgBSjuK9JdAhSN0ZnYIiqqkO0usQdoLtlT9IDs+2oDghfU20Kat
urn9GbhV39VRyOjljYhYs3JiTXn6tI8e6tsL9zW6CxH/BXrMYOaYKzsEWYeecQjA
nroDA3X8SL3MyNc88bg3nio4AePA/0HI7pgNRzuFdWNMP9hLHaG+DImfeWV86O/k
T+VHFFXiCBPpz2BPcwYqnVCtIYfqXpFg3UpdIbvC2Nzv8lkGVjEul1xjW9SWVeZz
9IePKx49ufD9OTK7+f8f9ssDB8WAb8t2UMHGt4MwQGZQasnjUenm2Hv7ThM0O0b+
h1/3N+gwchvpjoHT54OgWf5rem6KZI0AdyH7/UgCUnTeny7ueoW0S7Pujx9L3BtU
a5oq207bWnq2UR5eBMHJKwGIcwe1+r0G2p1JpUdiOOBWkv/9mmaAw7jMYVzJSXl5
rJP1KhNK1IPbNzobGMMXK94w6bcqH4JBnMvLQfTHx4kvUGKv/PrVMPK1IEcxg7qi
eMAGOGWEE0eGqXdpfTQJeDJGda1bhC2/GouJ5CGVscZS3foG5pW4T7d0a+IlEFKU
GEj5PpTc6sSTm/W+qDQWTQT5UqOVV9p1gvXAE46f7q8W29gGMebijOM0qzliJ376
gG9XYDFeNr0jTVTF8xtcnIipUUViHaskW+N4vYGwhucI1Mj4plWZL1zjba0RTUGD
UJcVLOAq62RO9HoH5NWjRROVBrJ0nB+bxo0e/yK1wEb5DAqHTsyv4yfHFHnB8fXi
skdkxQURYgnbuEeNo3bn8XAKiSzyz4SttcaQlsjBA0MYN+CE4mvvbdubClqYSU+T
WFJxzNlKlYCsoezmg0y7SuKN2qULGCruqcm4naKBsJIWmNoTY118sl0fNcagwdbG
DbPG26WCHqVuDG1lXygqhkZCWFWNRunp9o5m0goN6K0JXbP7/9lAA8ANYgp10XN2
+St1T1A97CugszXgtoF7m+eSxjnpM8VAT9i6IWyovL9vii801Lb5bEURsj9ngULk
56Vnax4we3ovlPCQVyHL1OloEAgqouRHJKKFD7C/UFLUuBpn2Gu0RvK9Jaix1eJ2
p2ZVEVOVraA8UKHaZ9ivkUSmttakJQdhZAx3IFVtNiMLUjaYXykcjsNehK3jkbyZ
H6pnc24A+iMv/fu5UOw2hQVGwXJQfnqng1diZGPZ7SbtOTfc4c8WC2L3lgBCbr1h
YzyuQf8ncSMjCo0qwosSC+hj4qzHyUA5W8OOL1LThiHsNALlAbL9XBe7acNwShOH
wT2KpwUb7YP/+2Da9i2+Ys2wlab9v9qDo9CEDsrQFCVLA9b3x5XEhuBbRSfGVvYO
Kw99sTDzo1h2qicBQeiwigPWR8000Tjx7VtUkJV8mBYdjzeqPMDLL2gC+a/n7a2z
AWWHzruuRj5sHTeHAb/avJmlUdJM3gXTPYRP5koPW8Z8T86I7A+S3KkPDHVP9W6/
GzWK2YpMFR30fPysAlG20BZc4vfnJ5jfcurGK7RQ5Dy5Ge/pAcIKDGVEFLFojIni
fhihQAu1FoV5SxSjl8htMm3dn5dm7ECSQxVO293Lvu+0635hXiG8Uls/r4z0qDQa
xuFNAGS92zDkNOr/d0yEJHRXXyzclio/psOuTSOwchBrPOpGZCGyrrZ4cTnTTRdx
s00kK8+598IkVQxAhIzhAMRcFVkA56DS0upfpsJ3uOptLKgoS83aGONNwV+UELNb
82DUke6FsFeKJyOFf5MvwNasv7M+r4X7lxEDVmeI4kwMBaALp7wI/RN8qNzF9MxU
FEtTmwXexQFEfZvOBqsPS//jsKh6Rs7LTryPLM22GIaW56WHG8aqRtUywN6hL9IJ
WWhGnJgzNyDml+PzLgktMy/9lfj+x61eMZdelFkT5L9DDgZFHNJ7iScKpaOGTWP1
nNK64TkRK3iwmcFNGnbxcnXnSrSfgI71qBHdHAo0yXPhE364m7aIXV6U/t/pHZUM
qniEEwZox1Ako11DJ0QmDwyd2xO60rlXZXqRJ4BCP+AbDWmcwYo6xL/MkoPTK0mG
LAar0Mnx1KAeHIJ5ihjS2Ed1oFGMEOmPFd4uFktjue1MfreTdPlztLySG2TyPJ1H
DWbhoZ6RzYm1Bnlv0IZIf3jID78+uzvZKiMKU6OKBXT2NeGrGMde2wSx4HX49Ik5
3lu8AXEwIBQNwSB7Sc0J+0CnmEl3SHYbS6I2mWVULURRLcy7fa6u+YMWe13B5U73
3iYx8jbXVNGduWXIJz+oQAy+gWgvVSHxbpBi8zf6HnPH5xRBJj7tUd6dBjDRzvfV
AEiXWx9yL8+cIXDWdCQ8kFsn6CRUWjZLYKAbWubT8FBbqO3qhV/uX3+NUSYLuy1t
K9+x7VPKOW4WIYsCGmxNeEaYDPgiftruuJjayV5ONFOEGxLuruIa9wJtRZUopW9A
+trgB4Tpv+DH04ahNWbwmbHOreBspXKAkU6+vghoAyhXn2FfEP7Tk3/ooqyyND8W
mS5HXPkptg6KXPVWepfq323D8Oj37nm9Pdg6CkvPI6G6GfSeXGFZkA6KviEEkzlU
MPlExeDRONgUSS7NpMs8xsuO98echpnpSJgjE3m55Kx2wKmJ95AP0izETuWx3ITJ
iQg78R4er3iuU7FZvB9z9ioAueaElxv5qIMMY+cqD796N1NFADSPQdRYEk8WidKK
ntKtOsxOfRl4Rho08LFUarpyYO8Ag61vMtXwrgTrbtk8T6fiDStfgb4oBIpEtzJK
OJnM4rajjUz0Fq7ZhfMAb7xF0TnN31FtsvXTZ6kgwddALonXm0X53/DRTO6lVZZy
fXE/BjVWbgnjBWxpVfst4JL+ohL4YJXhYmqdMnugnegDrDBWYG2jRQv0nUyj8PZP
Ey+r0Zj/1ndlsTYwH9ZMsenIbffl6RGgVlAOB8xKOwmPNf6HEqOzOJPkCBfIg6mG
p7AAHwSw1L3WTcBwMEm1Sprr1VGQE8qQiyklpcDImZGWYiWViUcLpS/iZsBiquOw
1ZwnUxATomNGPW6VgiKwrAhmDWOXNn2y1zQO19LH5wejR+IZygROjBocA544FsNv
bZJUDQ7YgBWe2upm8ReuvAoJV3Xi6vPogqSzdHYG6UtH/gnF2fuxAc0ys2O/LAHg
ITiKlzIAbZFbW6g5i5gxnu8hKlWhSn0vYQRrkxBJRw0N0F6W3YPGpqeqtuLcRR1z
RtBIIiFKNnf93j7TYv/e+bq/nraiQE3PRdtF6WTh+cRsQ8cpdaMMqQuG4nlBimcr
zke0f8qA2uktYkEQQOCpaQzvDkHBZxKx9f1pOU7vOBlcGghbxx5rkjcxVZhUzUaV
I7O4BN4roKBl4g+Ex3bY4tWAqJWkTl1ZEnjj0mWFXYbv1N/5bZszoSdc+uvuPqmm
8+7dQP6+V59mna6tlnQ15wS2Von7NKA0vNRtlIn/tCKhAp4AUPXFA4I67pmSqIgS
AkAz2tnlAz7cU1knOZCr8dw3foK1RqOOyVm2ZJhUymRl6mrNShiLApnKmFZUxuC+
SbJk5f9P9CIcrKoEGKWIweynbVXMwpv7zvhwEp8ke+SS4P8yVHrkAvVdVXBLLAFG
DAva347f5rXkGMoZbiTB0YxZYaOAwG0prjWqC3X/YtPklns6j6wRqrdKFuNxmFD8
Gb5NLhDL323TCEt3uea9fcPkI8A7mx+y4OP/XfV/vX6mXy+bHFUZjl0hJf++Lghc
gM7qvMVOhDbSb1j06Tn8+a3iLyTiRLNz2+05veF7DBYjQIWTtcEJCFiSwjzJ4N7W
+8I98tNgjjdIom0Dnve3vRIM7nZHh3TljfAbtCpP5oGBJA/k8+GdAWNtsrxQxK+l
/Wyk3YQWZmKPknZ3bXIBFFN+v8IsT/ZK4IbHrHkH9p/O1199JHjBE+HG0l0i0W7T
Zsn+zpEt9oZ/JWRj6L1/HXLlHYBNw3oSuhtDDJSLAXsrVNYVlcxLdICeEMuQNdAd
zVldhN+9p0DkyGFnLlocVuOapUQs8eeXJdAivZC41tlDv+q+xbFjsD4562cw8gf1
ja2ieWcrjfvV/1hvALfPgr+EaRZp0onrVe4m6UGsHCiRi2916LjF9sMK44LSdrCZ
uq+GKXHJAvFNKJeEJKSXlOC8Cr8gD6JBbdi1iAjml7LBykh0Tkm9SV3Po2MDPVAz
kXu9L8dnbfSqxhq8REnIdOP3815mfgl+DhXIn5qqa5AE9E+mp9KV8zlD+ddIUCNL
L9rZFIwMyE3htuovynu2/Pj3CBZyDb8VvR2TnBUFm/rjCJ1jgMdR1rmiwIhNP0xc
7rT/4GfvBWM5hVXPGRiRBH0+KqPjhDG+SZE02nwe/ts2XswwnxXRm2npJtWCLuzG
MZEARX1lmzjVwB5OFvFJTcSlx2VYR4t6iSyI/IG6M6eURGCsxFwZdVqn5rNAZN8J
W3nrLLnq5ghe81QxdzZN01diYx9Tpsj9yCFkMtKJuVrr1S1yiWfodpg1fG/JQScD
D8Ji4p882BD2AF3pH2lfl6+57fpNGNT9iamnE3XYPOtBFPOopvqg9rPmUmaAMAkG
Igo0/OBye4yPF/6jokOfVek3eQEYbKDVogqUvvavmOjz5v0ObKdTE94v5b2FXkNL
G0zXqltYWaoYOwG3S1eBvYW1IrolVnK1aBb2xi0k9Zq68sdnkycbqiKCL+gixT6K
TIsRk+EBYnS6nO3a1gMNRqD43OnFos/ZFIczwpyjBz53H4ehweBA7bWXEGOE6FNc
BR9MjUgqpbaeTKeCWFJWMjJI+bWF+MPZQspp3PkYsK9dO8AhhZ3P7H2q+/WjbB2k
tu3yeSaVIOdCq7ytRmlsRhRzupgDIJUe2Zlz53BTiBSbj2l9JVf4k7n3Z9n+UjXm
0HJvSCq7FHErLkfcCgG69Ues5x7eWcz2AQj7BreCrqXCxLgeCBiRJZBWKLjz4TVf
FHfYksyBZx7WZhY91r8R0gUrIS25trkcOKoSUsNykg4C+EZTpFls0WymzXsZCbFs
V47U/SAy390SF0d0Bb7zdG62S1f1hx+GgnCRVJ/A6p8MVWLJKkEScBxp0d+um49N
VT+7eLaO/x0WN38HhLdWeLDi/FdQHnsg3Q44BllThGVfW7n+L+tnKgQUh6Mcxd6+
2KuJQnhAwv6gdbqE7D0GMZrSTNkCBZhKQPSXCD9cVottvZWcmEjdHnTMmXOHCiHL
lg4YvSGseJe8tEcOYYk1WRrgJekH5febYg39EketWhkQetfoIR4GKFOcToBcJ5qs
D42yQE+8cAgJ29CH1jDt4+5UxMFFajnsnccoPLZmxxqoYYBQsINKBHRaNqdfQo3s
Rb2UOf0xA2W62YALkbe+R51gGRhfY7zoHdP/mShOg9gBUHThB9/av4oiJLsaKYbS
Hc1iwYJ+AT3R2AKETyZUssEjS/AurAlR+wADa4H7SPZz/m2JEPlGj/vXzZjOYTS0
oUR5lx0sLr8//QW8gYlz+W7of8u7vOopvnbw1UUHb7p4fTuc9tP7qi5NFO8dLOri
Qjp2R31xuCOco+GWDM1fcxgiwU+hLf0feWktUJBtBli63jYlZSDKUXA1M8pkYJPF
HEcmiZZyFfivJPenKvXAp4XiCYgd2664mBaEwHKRJSu/PUe1Y+aVpNPnksaEGNVY
UPNdRfOl9MvmMfdCrW4QsIR6w9sI6m3SrbQhjO8QrGNuSPUaM0EbpT/m2vV89XKW
0UM+WBkWmBQOiw0QV42h1+IKkQfxaL+4vqyO6hvXUz3wx2M9aBp8Wvj/cGqLqoPC
raSrS69muQCCsSZcxb739kKE++TLtqJqvfh3Rj4kjSEhIHTfzWu+iblxdZiaZnKX
TaQdegw9aHfDiJmYJxllDmB5qV4EUD/7kK7iTkqK/CCVs/qZdsu9f6tOVMCtDiHK
bG5Sf53AwDNB5cvuaiZWRcLIykmTcAj5whiVLIcTyUa4rbGG47Ea503ysD7sUFEV
O98TBtaIazZujGlMIhi9EIaOYFwLU2P/GmEdbiaXkS1BtNDXPRUx5Ci/GYnPBWIa
RxSbhb9EwnhTQCA5RFzr5uOTxGHwqNK8SabjAQ6Z0cyh3frs8snv3i1NNuEc/kY0
h8BFLopoCocjrZQMOgndp50F4yswcw78lDCwbuLOgEaK8SxRTOYYpD0d4+1wtNSH
dEdleUK5BAjvE8QEI0U3e6X/LIevhKzz3sDlUo9TFWavTIA33PNYhPy1qjPLbZn/
ysjmsCcds4GFelyLNAcyPdjHvRpeNvOB5X+TmDs728uhf/DkHur7LgFdHDXyu/VL
EqKXaQ1lcx3K6AbTfApOdv4h2+RzsgFKzoT4T2onQAbrJFHCb02DrgARG9UwaB8J
6BjBRagjN8hAT2ca5s5wTkAYx1CeuX//FfxDinfKiet4jJufBPhZZYfPN5jvIDKl
4k44BFa9AgSPEbCLzSASDos9HTd54dOD1XR7uuPY6bpiGf5rxKDJWBfjzcc0dWfj
O9x5ozPbuXY0pMQYvEzrlcaYVgAlRbhNTeGOLtQ119+D7BxgEQetlBMPVufc9RJD
h3oojpV1dcjpMjbOD/oDEXrvk1rwwnGZ1oEJRAKSAJoOGQqKr+34zyzGTMvzWqjc
FbPl3xYi2qhqnWbBoWhfIz1WmgLuG7eUubv9fvdXCbexx5GJ858aaaJSNpp5ybky
uW93XSIbzTWY67X+HpJz7JAjnWMswQ3YbpVnr9HQtuQEyGPqraS2+kMNdohhkUQy
0X6aGhfvPCbd2yg9eEKVfSz7N9UHXKQztFghtfTLiOELoUJjqT8u09OZe+xYPUJ+
zEZxpoOoOSA6zq2Vk2iWP2gqwpF8SRCfkQ0q3xr6enZCxCjcXNppFlL/a1wK9DtZ
49WXxT8RD6V8sQ7nIHjkKTaI14m0aoiRykn7nRq0en01NC8AIaJJHNcWgWP6QgmE
m5p1UJ2vYZUvmRcI0PtjW6xHu8CNDqkkQlLMhcoX/ykvCc7iwEQekIjtxeFjfSbR
lr1GYdyKV9o1Q+vRIHTOWhQS9HuyKfFtrbpMJiDsApIRnMebuVRYUjR+vhWQ7p3q
rJhwFz9kS7Hq+NvxpJ9Rx1MkaBbXiWzCSxg2mR0x+FaNRyAX/B7iccqsEek/GXeh
Om6epUXPwPKHo5utlCgrRNU5L3VkYhpgp87J6Uuk413ee+kWnSwTw6hFHz1eyGEt
O6PvfXKJ2pDry2n40E7Sah5WBtFHXPBgTR4fpqHiY93p6h1FHktJTmjDguH6SgRV
P46K4G4sEJnpEP9z8udpn9CaVq5i0g3tNlIit1lQzhLmV4K7VdqTO1NpG5Og96PW
L7tf3KJ1lMkmU1T0J8K+od0hTXPq/YA9sGuLShUsuEce3n33l4G+UAeIjSWMhOij
+NEXWzsVlaTRKez9WPi92fhmfPp6GXZtk5Srj3hrGNwu+cdCrlQjzjUN9IFs1CRa
mosu0QE409CDFbCpZbawH1Hu8VEZ3rh9e7Vnn6Ybsujfi61RLj4DygX+r9YTceUp
r3qZLDD2QQjFIs7Pu6SYbQJBVgl6D22Eaf1s5xwdYbw0VM3QOW0OMUfRR7kL6o4e
J2FmHOa27pq/JY89lxSS7s6Hm0xFOhPMIxdiTJOHta57089I+D4IBMC9u3OKVyS2
/zOgSaH1UFZLbfxnGKPgdEwEYy1FNuui4SELC1+4TwxIKeMSFOjAlA1HWt6Y41ec
QD0MIh2JxBhx2Dp9NIyuaCw0DuChh6hUKrDngywEARh09mTIRiBLA7fMYuIDUI8y
DGdZu3tTAscS2ja53iWfCYs4QMoKB47QApw0Mhy81N4exxA9r+Yhdxo1LKPVWBjr
ulxMdk6pNBYqSQ3pWVY7zaiHFGlOiT08NDnKqfHCaHk8ZUvDkkLQE+i8DqMqdJq/
OhnUclABJ4+/0lgQi+NOa8YdG5XxZwwypy1g8JXE+P8RY/0QOcbogdYuZFARddaO
YOtP8WftcW603Xi2MEuf2Y+Ek56jscKR6C0+FsBEkl2kwDGZPowE0y9jd6yEQGT6
no/Qqpddp/2T0QSpVQNVnuexTtq7nEg8IqKPZG9ErdgE2cLCmtTNOnUHe93JvJfS
kJzjTibWUH4aDlysAvUTt7r3HUNlglWvVhPBGowpnieWyjQjOkMJJVQJH7BNp70K
Snexv4Vw8jV2UsWIETLcNQiPmNeRVPWotUvP3Ju6xZaODH+Hqor+g0GBcG6DsqIr
JrPhloSFYWgaDASfVddfp0glrPQQLaeByWsCAldzcjAXHxtS7Cndwrxv9LN8Qn5t
pLNSuwIiumIcAdQsvyRNN9DavGECUATQzPQvr9960fH25B+t1vXRI76lHqAQXD+7
mWMzX+WhimZBmmpL+Hikr/qwaOKiOOkpgWf7rOx5JENoBO1HFDqc0coZS3I5DaNN
vaLcud0yd71wkQ07REO8CoHNAaa86CYPchlUQujytFT8HbyDSkFndCrCYPmWmm8b
zc569Oed4FofXAM3WPajGFZV3MmkJRak5o+P6kpz4vL2LvxWOzR7WUagOXm3C5Eg
P+NiIDq2ykxvyUX2c57b05TQZJcJsIGbLeh/VnrEDjzae2G9t6Tmm4Zfh9BG0Jzw
0p0A9UVfF8KRK7RLGZINeTLSZ2X9f/+8jtb7+04M+xvTEktBaKVKXSlEWeEeINB3
ZoignVp6pe/mb0dFqVfiI2pEof6tHdu1P2KSWOvCrAvUsqDPg312THKm1fgNcae2
UdLEO5qptV6aL/gtWk1dnSEhRizfUC2BZBlb3H3zBysP/XYlhZ901tlRtxz6dwTK
3JcibhJh6j4zU892yek+/V8MFFnF40vMaHzhT8fpyLh/PZgadn/fMXlAT+HIm4av
jrkv1ATzt3zv/BImpawbqNpKT8GbUonjd5kgrGtFjGLzo1bGJrbEjr0Z2jiQPdNC
53QI1yADcJuOCNv0XOxg0E6DvquP29VZUlvQdhYOZ4l6Q519JN7Mt7+dJ/q5z/Tm
EU6WPtCu+i9rJEPx27rltTkgiTyirV34HCv2IgQAM2zmzslm3V6zoIo1mDUHY15R
fF5ZS+rVLQdJjXogg+fA/InqeC+2vPIEVNtrckic2CdH83iT8VHqhxzVRpeC8+Vr
fajKP/tNT9os6LnMSTGPX2nuWC9WvHL7d/u5KS+PWwecyMvzzSDGSbwCsKYNWEN6
5b5bHRJkC9u1aTUWwaIYd4mhvV35ZMoP9mAT1tfHT1u2AjsED/EGzaaIZUHvw3w5
RiB+ZO3k128qP2q6LI0kHfJ29xvb1T3LvoWoZ6MjGpYe5hY4TtIVXMUFQX9Jypjv
u7dCv71xRb7o48tmLM02XOc8DcEYQtj18TOkeRjyfuECLQHodOaAe6ngUV5JH9O8
0kE0U+1qbAvSLh4CmgsYPZREi/KwTMzrguPHy0cFyDWSKMQPlOACHeRM8K15Pky9
Se5eKHce0WNBno9ScoACWYugXGgJ16Xi9CLr1pLm+sUhaaXwWFMhfV9f+JMKcX8o
1qrFeDtD/ojViZ1Gqjs4f0qAYdBsylyPOhSsjk4ZEQh1bFvtULGgI299JyDErioh
3oXmc1s5vCFx4fSuygTGq5bXBmknQS2n1GCl1r163+5FxSYI33aTblVgmMMoerZK
47+0Y1Rt5xZMcjkIF0NonvdhgDwBRND3y0QjCGYuKSUWuOKV5XPcCIHqsxCknfoq
jm72i6T4LAbS3ZkqX67s3Qb9BL7OE/SaahLUzsOAeDHlUvwKOnpa0q+7qcPPgsbI
DdakzU/OLxF6usKZa88PxZFwYh3zWUMp96nWH+EGKIhfS1gYEZdcJoVjSJ3/UTmn
2dJQtlmiAwxCR3gip+1rPAGcmnxzT+4PCBdk2VG8g1PyxbNY/vPdV7JFWkYogif9
SKomVXTp8oDi7p36uwUoslqfLpFNPKYmn9rZUGNToMU6mdPsH5WRkNrbHCw+EMSt
E3vcS1+RJC6yZVxSmxjFJrlqpofy1CpO9SB9ayRWtW9iG8wvNFNZv1b33dzu3TJB
f4LcbZ9mDZxnL0UonZ0YyIZrTpQrseoIQb1ELyjkWEDqJneHJw2nGur5rfwl2C9y
w9/SFRvrmUaof0GpJvv+0IZzdLAXTlfNdKmHsBQAgE5NprvPYm9brCGRIFh19Sf4
0tzL4VpXfmdbQSYv5EasGc30Af789Fg51hAuYCBUKwfmzQUnkL9wrnCyZ4Xxcw9Q
POR4E4ppKouxQDbozep++2FKtEG3Vi76w0xT7NakuK5OiBoK4WEgpJ5pDlGl1u8O
GH7FxlNBl2/ID2INeh9K5NwxqtRXHUuT7le3aLKeapmMd96NwiSLomSBy8eFIz6X
Ck9LVUPOzN0T6/5bXOZDPdtsNdGMlFZ+NjpLTyKb2v/Pfe7idfXbK3I/BOPmiVIU
EVkHFwgI5KNFVtmSGc4XBrqv/v36lUr7HdNmp5UD0QX0+EMIF1GXckPojnAdKwcM
MAIH9bImgOfczLvPJHfynKwySotb9XKgnWzxQgYPAZ41CQ4kZB35riJxrLlCOqhA
NV44T/3wrL9E6g8/unVqyCIvTynYpPoKZrXZQ+oJsuxWRciczEjqXe9rB+VTw6Ki
i8+oUTgF8zKMPcBL6by9GTiNe4vfhfESToJAcjFxyeTUFSSxMrrBht133lR+dLh9
AAbryX0poTVYb/ACjYQtRpsXYgYvXZZMYw5hkuS5rOonT36YF8FWV9qE6eFqtjXC
rC7+u7HyquGYX4hwWpGD2u2NvSxjPalScp04Dmi5h4wQMZlJ33C9oVHMAXr1o2MN
nj2RgtUERAlTEdawxrFnZAwg/XDg03sA1gcf2LsHD9+Ckr8NSPnTvXQQhF5O86ex
o5OrNDT8fwMWMgzhwQPOb+tk6ScXuNPiXj1yLxEVeikuoBYWI+RtENuVgg7Lwt13
gbzi6PbQ/aB+PvfVWxLrO+8RlIm20j2G0GZAtkmN6lKZ2a34TKN6catOTJOwucup
lfd9CZuVN4OWfkIYvfUV2QwJA0puChCMBaetSlqO+wRMZsP3t1oPeqc9bQDYyMGX
PrRHQnJ/oIOICB2lbAqh/UxsuLkRVczRJtUPwh9IpG3VarDXtAz+BQ3/jCYf/o3C
tvpSVoeQG1CbIVyiwXO/q987ii7F4Aj2vaxHgwZk65FPbxE6AKCjtWocObtSu9fm
Az6EpMYytws5mQDoD9+JBGqASZQRGMfKMFJKpxPsw2DkC/W83rz8dHGtPBzktLWN
VLl4IwrbQDZ2JRBd9STw1TVCIRdNlLEQHS18r+EZeWsvazI0Bu1lJ9dxOF9NUdvD
VcIOzT1XMGZegxEtx0bCWbYwP65OHCV49kgh0qBBHI+PEfwlIsSGcmu+11DxyAlX
TSb43VMntKhEyvlJlf3n+JZL9Mgvoo0AClaUOZ5aLt7F61/AoVBr4s4VVbRKNbOA
5ubJC08mv/sSnZVQsRp0Fy3MibZUth+EieId6o9bzvIjT7SLmOSsjnTFp9p5y5Jk
iiKkD9b1KEeKuRntET3wpJzS/Xv1c8kTgBQbD9YhrWW4944T3yJuy7/tBdnM81V9
Asw8JUTdyZNVXPje/JG18cFIvZcDohDi07c9xttcAbs5Q8s8fDc6+R+D9FsDFVyz
XgWd4X9DpGr+FjGo2aJquCqdnYwE5++gmZfVoF8Lx8MpyuBWmDAAIk9vhDgj0+wH
GZviSMQBRaV/c7NDKKesWD/HelLnNYG4rXVs9XoedDoIuEhLhM7kqGZ9Fh82MFAN
hdFXDyNmMinPFyvMLI0dqI3TQIBJE1hB5UWuhj3sSC+G+pOBR+1PqMiil0ELsmRo
HI09P7rvQM3otoubnA47s4FUQV0b0OwFYNN1lQQ6GzGoebV6fHQvmPZiGjM7Y9yd
r0edhi9sgsgJs1gZYb+Mbf7c/YxAoFxusH5U9/0/8QsQzZF/SLAVvgKfbIV0iCb9
xxPS4iIdePpgnKwAEmt2p4ujAfz0czKIESbsQ0wZm99yxrDskKzCkAZhCVuQWNti
q2GkPSVlN6ZuktcO0yXTMXqKIJXdktaU69v8H/UUY8eQlEX6Lc22tW2DJla8x8X2
ofSZmxybTZ+h2AsYUdpjM1Qr5hepOZIODS/qfQhQ/tfrlF8PqIuZzJDB/W7oFIoo
YVlvlOp/FKwU5Zkn3iYALi3ygzTY0Iha2p5R2ysLupdoSX96AtQieGRcUKE00QFC
n+UTgzOXGbv4nZObJcGf1lPYmPYoNJRvUnkULq/EKzTBO91w2+tuLSDv6go+s0+K
BPR1BOrxhjsaA2vjab2S1TMaSsKCu4hhN18ZV/YLZrb/Op4zyohzofHRd7CsefyJ
4Z+hq0FvLHuEiHnBZy5XhbaJZE3z9YCETeK9/+oscYB5qtYNNrKvduoQF0d3hTN+
H92nyQ/vS4vpcPsJ4Gh4zy6hHuRW3KUavMznpjGnRtutpkXeWpmd62C3EEORPyef
t8rZqXQLQyTM1tns6hAon61zdtskiZPbLwZC1zIiP9Gpzoqo3Mdu4HoOpvtUrhLW
m4AUDZYYxaayjx/CqyhrJFeM6vGihhm+83TrtTzmEuHtVFnD31ty7tGqxxZtWH37
t4bEregbauZkqkZwLoN27hH+MnNy7d3OzzNaHq8QJcJjpeMcDf2BiBbV9k3amn9g
+iieNq7K0l4GRUrh3aBdC741uU01ifh0lwD1Gmk/5D/uU/v6eEJXDLhGfNLPA7z6
O5k9EBrXbE9nMlWjLh/A53M8aItFjC07RZ8P6hoEZFCqaV6Jone8BqiK4zxCrjed
XCAO0deFQVH3ekK2imFWLyAzTNAgCekLeRKtXcOLS2Ft7js9eN4qjODGeMWEqKDu
nK1D1R4bA4DudVeFGl8U0UzC34WmPCGiv+K3nyIdS4M1qBZhybHNeRFcZJn8x7xP
YE9GTBdRxJCjbf69WXlZD6sBXVaYU7v8lAQzjguiCw4cDGUH2sP0TrloCLs1giTA
uyL9sHH3Ax3lJQuC7DaP+f+xBHqDAs0/izfGCIRCDlw1GOWUym06UrPiKkpXgh+h
Ek5TgCXhiofvyxr5zpjayVpld4Cx06h9uhBtL4PFV0DEi+DVylmai5nqVYkTK6o3
wA5qOmgPlO8JNp3tQggNZvfQ26nKxGx7NZsSUFH1pJSVS7ZjLbTQdtzUxvLYe2mC
avv25liGXdIm6DI0+13ZNWJI7OCiUc9+esjHvfyK0PQJ1GZ/y7LU5U1M+fSrt8Rc
bybArQmE/gGcK0vybW2ftQNWmqj1Wly1pS4ZNEWl654R8oMA/4DdM2Lqzjau1ECP
7Jf0JmRF/uAGugml+/KFRoWqm/zLvFub1EtlUKN6vcOiBWK26Me4MLXdrDA8E5FH
S4gkV7UvJMVMcpx3vpZGBSZJtUfFuDUeN7yBL9o0xQsRhj4Hx9+H5nT22tP/AhJ2
igm0jnzZLw2UCdBsLBREt2nM8ANCibZyMFqytJW64DJ4GQxAYozSfJmyFE4Bv+pF
nhBAiNDe6E0mz2H/cxCwoMtQR/PDspOccWTdruy/sAnaq0LenXo486namlDl5ugP
JHKD59cMpbSv92YkN+za0P2D3DOmG8q/i5cDOQISgNxbHY14ge5LnwWvKMoqnpBI
qYOfEXBVAAUT95rhl/rcXoKp6kHYtdSaeRS2zBxeVqxzZbJWhuOErSmMYFW44khW
4IdUtAc9j5KRASzj/WPhHSZoN2XgLRGKmpB5GlkNy1Z/lj6jQgNHphI5E8qYJzhd
lsjCarh0eDyXjglJsulIPMFGHu7cHm+cyTGZeMMfkrPq8tq7WogtmUQtQ5qdX7O7
WrD/qUG0lK82p0kgahyGBjXPSppFrTPoSFzV+2N92DoPGeKlh+wuNCremgrrlpOQ
QG0QnXMKtVsAo5/xzXTQdEmEJkKYJGm8RLgSjUExzBdGhyElJTcF6RWZojdcA3LY
N7b0lRmWgFnsAu2iFVckf3DLPiWt2mPrprDnGm/C4q2BNCTruVKMxFFmrW95ruFe
oLLil5Ow+VgRvwpIz1kPuBmgOsq/XLVH2fRWiiFBkb/20L41h1fpiDqAztIh4/9f
0S/6qtS9ODrA4wiXR6+K5qzDkatP/A3GldRkUVn9Rbj+NWTH5QdV4lsiLKJ5uxKJ
q4BeVcL1meka5n5bFsrDEgtcJmQsr8EwfkKzfslMh+MYsl8DzyYbzBlsClyXSlUB
3UZ53fBq3E2lrsfumB8NSweBONhTWU5cH/+u1KJk0CP3nnEDoALA85neUt6q45eS
UPGlHVo974D2lEdVX1ZUA2gczRFS1qNecl+CTAaVX8HVZVzgMUbl/H431ozMeG6u
9jq8NZMtyUPx/Ero76tfYdBzQxhKcgiISLFJTsHtSw8uT63lGIzMFdnlMCF+j7P8
8BSdlegNHampzyXR2ys9RJ33IxNPo997MBTh0kstm9BB82Zo1YgFXR+fwfqTZgwe
2jrs3YwngIWz5M48vTZmBK6WgrTRGUi5+6qvet45E4pd93/kTsw1RBntqyYcOGoY
n+iN6fJBs2CM0A7KKxHd5FhpXT5SHczA0BMz7186fLdQDvmu4IszvSlg99bvZJ+E
7zC/6+OsloEx0UJNYDmDUKSQGZWOX2+XdztsJv0jWpqiFrepBAoSYZ2bEcZ7jnVJ
Y55AX8QLkSzh75aOC6Q2oorhIjCova1pv9V+z94gj3c6DYlImWJ6KJs2sQam0l++
vub10km+oE1EyhvoOX6CzKhwK/2eb18HalPALPyq0DwmnoS8QmYcW0dM9he6FVSA
GHHtrCruH5vnfXWYVGHBfb0HxZcW2UegtCXMnGfukIk3+Pf2fj+ysGhp3hG/B+yB
hmGwLcRMH+xvLkKoN3qMLtAFNwgycehts3bcQZOfvGDlB7ge6tafAlBjVeAIUN6E
MZ/jjE48LEyGDea08GZVleUj7dr5dxgSC9gaKmooZtltiJCwG6YSobQhRJ31IFYP
pS4yj+UD1FmtL19McO9eVLNbFW/Gn8N5NPSKSPyIHqA9vgjJSFfJvQvIf5oVK1O8
IHCaFvzon+MPJb0yzVy+o+Rml3iGl0aG/gSUmNy8a9EzGn9cIS76lL4zaAk3V/3g
jEvm/ou1mfZZSobr15i9CxVfqwGtEX2r0XfxBgOrAfEGXrjDfn1b/v3A0zA79VZ/
efRYW8AIzDnVVqoDDpRGNjKTFQWfDgb0UekI72YwOvQ9Mro7se/HqmNsVsWmSZ9r
JmtQVP+ofRwSF4niDjQI9HSEus5HyWArx5B5dTBLyqFm8p9RtJxTtPbxX02+usH8
+OG/KkrIgZpxc+BdTKlq1ofYfFVkNKVE2IJ+9UIbGtEx1LgLlWP+TwEhd6PWb9Xz
su+G1LYdU3u9t2OuAvylJZsIqus2bcoAGhTyXjIzuU8Nt9P8+I5SkK6Bf7TP0J3o
xLrbjtYHP7BxV57dX311z/FE4/938SuvUICAtUNuo5IIhejNGZXvsxOU/fPllfkj
0zVtPQ/6KIqZMQhL5Q6hHml9yFJqISV/7Ud+TXYO7a0Vub6ijtW4EaWSImyE/v++
wFsk4wmT5J9x0Dh/upduI6CW+ofll3FE4N4tvrHfL2Kjn2NdInuQ6q7ty3tTGvyw
UWmHNttI+3hoR4TjOVqiAxNh1+nCOHN4UXXhwaWnnopFMOUTW+3NFY428MR2mGtL
ID6+Ecfy8KXcmXIRoEGHbbEC0MTx8VJSHi5/rjRYYa4swSOm60pW+ZePGYu0Ypwy
bHYMkdAZ1bczSPsfSOQWKYOpiYn0E5q/v17pYGo4cgUpZLXCdA76kw/gDvvFpAGt
ayVLd8lbgGIfMSG5FM5iBDkiQBP0+4kHODV+eTcUNHKBWFXoKHozjSFMyuNLGaQk
r8EXG2vIQLypuovWH91AyWOIQmvbmQa04bsCzrZ17CFU6Z+8AkM9Umbj6Dq/L8/Z
kLMuGMZs8WRkigk9viggfwR2d5jvMj/PNlmbWX2vJjzs+iKlU838gpdFhZ68AL8R
XupbP/EK5mfdN/o5lE07gCn5qPESJMSISYAxXUXcrKuT7BhJQILnBeYS5uUY7PIb
flXkbsfdqPPl/B3fxE0TRMWm7l4nkOqkO8wE/hJjwgSUMQmFvZxU9TZpKkrqxFMy
Qn+9oxeWWwP+g0hWAo2w4YsFum4X8NZanGbR/oYOWqLU0//4mJ1LLujeP1a1Ch8T
M+scb3b9oIx5b1Bk1waFpcFyl+yN2umYIHmRtYI2Pn9FkmSOG/KjN4w+9UFvjTkq
uKV5NY5MZP5jhE8QSI+pKqmKFp0dq8Zj2YHk3tcf/lR1Odivl5o9i2Nncv99Meo/
2PdoWb8H2vjCDxJtKeNXI3k9MG8b6GAPiTEnJusd5YWcbBA/Z9sFEj+xr1NGnqUs
sj5CFiLpZIulBlAnVcqlQCQhAigGWVyu3PT18I+JinRSiTttTvrGRdnq9BaLBHHZ
UAAKb9x+1vuGt3I/fKZWG6ajqfdYElECkfxW52IJgMkThAV/07z8nbUwiTItMihw
NepCLF8eLW2aRJ9kLsaC+k3zdsFgyFAGfpWDpBWKCaeMkbYFU608kRMd31EEdEfT
ZdNeLpJ6tqIwn+vRI6g7PS5ML6ox0JB0WHy2cltxhNbvfiKF4Tu+eezrJDtG61gD
6VU/lxj/csGA9IQJiLt5PwWl+j5nkMAgyg8+IsVoLqhMF8LiUOVTKyMYq99q/FHN
8paTMB1i1Vb+FSbJDURJ5Vp375A2yfmAaveuFofOgjmItwzti2b+pwwkhljeeNd9
gMpFelTVmQf1x4JMEwVnSdsvqxwGu4eEq8OOCfmalFRrJxI7gxZBGuTNIF6l2CZS
j+0p0LKZ4aPBE1hnD+LwmQAqGZ/qQDl5G3/YSzcddcmeZrMb4MJbfzmQrXyg4hhO
UxLAqkrnMPmTzQ8D2BU6Hu1hRFVe3x/lYMbpkdw5L2UnU5rrAgBfK7XflggcoVNf
RUNLbix+C152zJotR0Ri/La3DFidfizdYk9EGtfn8xT9gQI+13oBpZixWWbF3y24
A9xc8aumjpJKrA2eIjMhTssLOLTBjdl3JqLaECwDAP9StVjFmhCo9xP9ii1/hGl3
h2UxeS3d9uHOewXBw2gap6mEGfRjsjh0VMZwENhQrBhrnRuz5Vt9HlpafRH8fv8D
pFefbCSPXN4fdVnef4xGHXqd81UOpOT7CsKo59kLVjWP4PgHIV3WLGoncoVbgXj0
djNh5X3e1g3eydaQDhDnBvNiG0Mieka0Mc9KNzbObtamebOe8F5gdKzSXcmg037M
NIzgFIqa/haW+zPmwefOs8QfeaMEvusZF8LrYqRoDC5GFRgEQOC6B2dvw+eUCfrX
WAnmH8SjNAr+WL4csFUDrC6Y+EZCfGzCVlk3HwTSRN37ivirJpG8L0reSTVgyxUb
yM/eXhcnW4z5t/L31m4OjJaTN5i7NW/+0cV8ZSut9IFdkhKst5+SySQWR451zTuc
Zm1M1YTvwvtCbsARJrPvs6TKOEhGCOipvyyBk9f1bvwKdaq5SHEiXYi+jpoyhXor
wfa+PP5d6v2AseaiAPKsIQIvcaNr+lmGExkA2SXZpD4iN6d5OOhhhSXQ2L+2Gke5
4FOGHZqHsltblvyVTuMK28/o/v1/KAGvsNfS80GbUjkueFLsYGCOqFgxsBxH88cx
DzLfqm3Q++1l1vnP6+IV0qwO1E/Pe+HJgPWlufk61MSHDQlnOzu1ex/tVikaZ6h9
LmwNDyFqIEvZqIsvXPJVxCVllw/q3yfHd/BeAwxHLN2IyMlJlrHhYHEPGCuH1WdU
gNpaiw9ck+Yyf4cz+VLVmbVEiIOzAoChRZJUNrUUCpZRN5g1mGFp9+dNDsYKF/lZ
ZL9e1bBDwyKEX4gCZaGmodoTwsrjkKy2jfUD/HQrR9lY8sIV4CFqZrLDbTWB6VfW
VCHyizd+y9EHW5L5nIVtl2n7OM0HRzFbvxoBnpPK/mYOs3hmz650UanoSao2Nmf4
fH4Cf6385q9AJQPH8nXsSzmSccmTM+PgPe2Q6H7qsy2O+JS7rLOc0f22ivQKsyKn
ptUWC8BhJHqLY+TiIAtREP4yCJ4R+NXNkCSMPj+Vxt6/dAJPeRV+o1KJ685M8Tch
cU82LWzseMSPGs0ymI0EJdzBjRfVauVKD2WeFhdCOc3T281FXTQrcZX2sjf8+tqS
T16AqRB7GkYfpLmKgIr2vWESWqgDWTABqEV7CsGt9Bc0ugmigLmJABEPsUdIMNBY
VkCDR/0R1IsNXt8/OAJU1drzoLIY7HSTDfPXgTd44sud9rZLOczPNTbfh0zQFx4u
WM56BNjLI532sysLMs2LMMHWqXeh2Tt1AP7VH8Q7V4fe5tr1ZB3prPEYKQNHdd+K
Eba9q5YGmrnL1cdLc+AO1wTeJ8YQPtnaAn+lBx1Qp8emN1OIViC1PBqK69zt0dSt
WW/xOR69/5uGvHFaZwKkYkTQ2LJ4fvqtV1DhFiL9nuAwI+C7Cs/4YJ082HrnknhO
GJC8rXAk9X1wuaT5IRU5qXfc1MAMOjA9RQQw4sD104uNx+Bx76PoxijDkn7nrC+X
BAY9cIkb4W0MNBg+ksexfBTQcGeNs6/QY4Um/i/U+PSq+DfMALGnPeoHWrlU9wva
vFf/dqbacGZztYYtYNfGDceY7MG1ZybwwwniQiyGP398scT7UBesDhtoMC8B7NJf
AIBeEVLMq4Fd5KEiSxAuCEWDR33MgXHHFSIx3CiLFtD6FA6k/EA5c0DUgK0UM3WH
PLzATr/s85pxcCZoyQWjO2IMxXBtVRU4YjK+W7HmefA7ztGr7VERc+Tv90XH/r4D
agMN219Amv0TxEbTjXtp5KtqV7lhlzTRBxr9o22b6AJtrK6/EARI0Rx0yIaAx/a8
9MUwVN7Oxiw82eZ4u9wU1RyelOFWxeDjqgUaSNA38FgPcKu7gt5iAcfXs2Dsug8E
TgzWgaPoEqmYdw9MTuwZDIl3U5nx4XxydXCFm7iCpKqz+b/4179f03B7Ifx0HxzY
+LB1g7FpQHIcqpKnxsXYd7ejTLMvxY55/ygPXGK6UaoFRWe998LvAuRZuhgzYlUx
TEnmSMhCseSeNmUqPRFA0EFSmeP7POng0H2NgUi1q24s8KsRDQM8I0i99roQMxQN
y8hqp3ErdJjWuQyIo7mEwsK7Ki3QsjS514bEbOQKrolzrb00RQNTkWpKbAgJkCyN
GLwOOXU2+kwGp7KM0o2IXNIjpoulLydxJ6LRwONec72XC4DdAv7YnwXQ/rgQtKSN
CWFQdTn0mNZDPUPieW8CZgVRvvTe3n/E0ZgQStEtEDDansakjp50tftEDVDS8JWA
41sxzsiX/j/UAmN6pv9cIwtwy+HEso+oiO+6vxrSK7hdSvDyw48bIbmxlmOW4oRi
QGUS/JpPyj9RzG63I9dj+22o8mCdcdhTVSACqtrfy5LGnseqiqIZpMBFhz2kY1+d
N7PfAS5eCiyKLda+uS5aSBqmUBe3SeWpBB6ouSWO2u6FUZnWlDuAsXvqR8u4kwpC
34HMz3hSd8iltDdWmXzl9fg/pb3nqi1D4yUCoPS2QHqKEUWBK3D+7DVChO33k5kh
f6/z9XfkNcW9hxQife/lVXMfnQY6CUzid4AH75dG86vCuvNbmJYInjB+Xrf+M8+j
kAUGXyn//X3Jd68mE8wzFQgKTQh+R5FDSuWlmwQw8YD6oLxc+0o9p5OPE+nhI2JV
Wb1PdkrRQC6VmtN30+5619sW5pdHiko+Rzb3HpELwQEzNWoQGqs7gAy4hlG8NMuV
eRdl69zeSt9Og89LqLnRuv/nRk6DWGjyZZEKjeKabxq0mu6UNKwFgkgERU5mgtaJ
476W69sZ8duIzkmtnmyQOjJEnThccOnQ2uA3fuHXH1B6WNhg/zHSjLxbtO4h68b+
QWDiryMSmjTU9BckHLmgUYKiQ5LNAp1OGFtirHJrARTIq0HeulOoQQ7e4kens2lM
Rtm8fJ0Kjjb9znYgNeH+66KDSpgx2I2yNUCaX3eKzt7N+h7UNcwZ9IHZzHSlxTHq
i7VC/NwFQt5VaJOBc2Z1uQdG/w7y6Vy6ZKNzO3SqEV+AnxzrK94mZqXdIs9yPVtq
l7e8tjvmCflbIIE3mydeMnSBE29K0gkp2mcDF4cCeONcRNSuDF1IjAePVnftiRcb
Xl2oCK6c/w1MuCc2ZupSQBB7L4s+a74A1mYiHSGNogMNMhZuZzCEJMmvkSsfWGuU
EMSFl9jonYPD+t+ctRNJYdW+B6sw0nBwKUr3KksJT31atBgRzGMmN7Lh0xmHgfP8
tE5RBvnY6Pjma/aUwfz2ajL7JVng3BqvuDj4ufXCz6W8VOdp+CLzTotWpqeTNRww
Rcl/RFhKylI5J9PG3nb93l5p6trduhr1L5UQGUtkAUPV8SS3tvrLUFydDK6A/mRv
BeIn8ehGmULS7Awuxi6PnvdhajqaKdnhq4OnS99OSpKCkonwuQKgiuW7+EjVVRGB
gVoxzWWUNCGg2v9onpnJISdi1XuT9kqJZHmZwBGoVSlMNs+yIQc/eW2fMx8BBn/C
VgLR72gstGRi12ksowI2WZTg+Y5anDlGBlu7jUgxjAtBdAKKziDbjURhcBRJI5pU
a8TEKGzNH2seStB5mhYFSzzpw3qOIFi8gx+mRfV5C1eDRRksa1wblSXw3OFt6Wo2
AxoVAakc2sPdap1awbpquMEes6miZYo2vASPJYZAiC+oCB2EbVBfsJbt8yn81CQp
dvMVhnuvZaIH9FAglHxp1kxHzLTBHBBVg1bldF3pda8yCSux15yxnArRN+61eOAV
85hwaXRg2ds4SirUPcL0SczTWZPRBLx0lp86VrNJFoyzaP6O1J44hPKQDK8InZMa
fMX9HZMObWtiSJK8zlkuHHDng5mRQ5+KI0/32pN38MWzE7b8TaFSohlpNfXLi3d2
kM6ZeMO0O38hxHgKqYypIhzY4ipFBZ0WAz+YQeoDvGt2tUDYUdk7jcULQT2PYa+y
qjUJxciUaKRHDpqLE1AIjA+mwaM76ZCtqQQioLcrvQaSI248jd3H6zY22CdMSoss
rU4CfSEwI2kCYYNFN7ExtKZr2++suq6TW3uxo2FR5/OOr9tdoshNFXiqCZR0wA8p
ORnYuWHJvWGwCh2+ugeanxLbiZPDSKwIH/SAnzXjEnvQF6zU2G8ZZkkm32q/N1Nl
vb67qtjSLwdcqPLJrcYWI91U0jaDvhQ36ZRbbKDE6WW1Jr1Lwf0z82jGEeRIAxoh
O4CYiFnG6vl+lW3HZiHvqH0Hhjrb+WKFrXLyGbuSZ744YqwSEgVuOYSE55nPMWmz
z5TjcCIP+J5BgUenbq4w5UKJ+TxJ4E4dDVlwcdB1PyKvccHFQP4zu55G6aMlcWMP
HBMnjtzM6TGavJXbHyA0DYw1NhtryqGqWM7dgKhjPtlOm04P+5V0fqJDcYm8zstn
6RykuqSlyhoSqSwX9QY3D7IaTSqIo2/tRBruphteni0S49o+yxiCvTuDq5VLJVHt
jCIy/+WTgSaM1ObmShpPU0KH0mZ7YisdCif6eXpK7rXsWCXBt53IuyBiSy0U+6pz
VJ0gasZz9vp9YZHp1zyr5c9g8sASpKgyOtX1e8dSc27OFF4YALbN7TPB9U80CY4I
myWcG4XH0JjV0cl372Vhz2qhIAbq7FDN3S7CrCBz0RFR+5JlYd04aGd78id8MJ+S
/yT7UZQ3Pe3wxhJmjALQUjiXDld+wXb3mjNM583+UI/1EudS12Ja/2Vpk5QAOn9B
N7bzB5a81SnlFFgbAySnb0mV+jbTxYEGOXDJH+TEAhRnabH/6UhFIyJ0BvtgMovK
8R7N3+MLuN6E9/EOH+1aMNcCIl+hjgx/VgtJy5NvXGZyWQbzOODOVt75aikUEZgB
BTDQDXQQ6ICjhJaWXxagyYYbtcZLHsFWy9vnoEoy//HlkpNLgtvzHJTfx+mEn6Uv
ooKhX/R5SjlGRGAWZLn2fo6oGp7n+MSg0ra++4NGuR+1Xkac/0OupPN6B6AHuKFn
ZfObw2RQgcfHs5D/UNiHQwn2LXZf3ffHlHOW33sVbh5iXH/pK9orjk2w2VYyvOqO
guuPREYdxCMmoAhaJh+MAi6ojU5u0XzfYg0x80mpUnBw7MTD+TvmOjMS1E3Z2uv9
eXf4FsMQTsGESUlmF1q7zTaLGvM2W4KuOLFDHbePWIBz/or3WmxYC+Ynh3rz5s2S
jehSpi5oIEPDm7xwvKuDqL6jNTTyTg8peFIg9kRW08Un8JhhrPUrVGCTsdFDut8M
TfYdKldWUdqXQJSgBwIsEd5p7BGeYvCktY21K0yrFMDq2cb0qWd3Clhfe5mk5FTJ
Krj3m2Ub6AQ+LFrBJtAjLzbjYi4nqFEDwOgRCCRkKRnjCZEqRcfm56FQdL18hMOD
zNVvxUo0NL0dIB3a5hBrn/faU3aeydvWTpF7NQIhHMLUAMytTSHOtty8GcwfYEjC
UAPBgIywxjQSa1ymCijohxiJe4NWch8rtD3pBEK0CTfNHtd8atMWimFaCoyA8MK4
BSxaYOpBzKg9sYwpZ2uxP65CZIISFjDZkrTrK3P123oWy/VHBBuhM+dQKbaCN+yt
Z5J/Ua22+CocIFauZw4GUukpyhSBOyQE2CWXXlo5Oe2FGggTWsuknm46R2wFTsiX
+4TQqUGhTWmipV1gc88K83YAQAA7l+7lt9P4+L+Zm77gyITUvZI/pwKA+on4myv0
QOOP3bSAPWjQ3dULH2/SCSCGRQcKT07e9nP9XNhRx0oLgDa3/R02caU6ENPMYbJh
/HhGBxzBnvxgX97LuESvKJCM5AY53XHbNCG7b5ne+7qv+jw7iHTxs4d0jQsrvAY4
PhZfmapYy1HB1cJg0graL6MZJ3mjdD5aT3NrJVTFOfV54hSgHbKcfUr0yv38DgYT
8RQFpSyFiJrRKbTO2L/FumKdjgG9E8wE0SB++zhN3XB1A/xLxFeUG2I9Z3TNW6cC
kyn0F8n+qndtzpyqyIN2sDh1XWVvnTxIUiy4PqM96tlXDUfM3x0cY2F8feiRr0K5
Gdpm1i23YWnJLshLcmPdRFkBuWT0nDqybfifKpoMwhafw4EntkTooEvReQuQ4gjo
7MpyTkWhzl1/v2ogGeJ8SVQlAKnzrhdl22e8j/PuZY4H6X0lmNUk8UBodVP7c/Pl
Zc4jJL+ccyTYgJArnkijk9sV6f/dyLenG/JkB28bxkByUv8Tbpfr5GVhCU+4L15Z
9XECSFj6yirQNPqe86QPJ3xOCK8eSSlDA1jUp3uVB5xLf2A4zMfUQjkSXAgOlznk
KMvnzP3So6aJ2fLA8Xaytkv4nCPbgNZZrJYyjyTQZj8j423Ya9zmE57LxBAXMRp2
OrvzRBktTE1DwtgEXpH5EhL4gAdrbXKe0sdHEUV9cGonRBecn1FNEaUbt5MykhqJ
b/rqFmie6GWutRXe7tXK9jHf9Ma/rcgLEJpOU408fUy6awAyZdW8eWKYQjzFITe1
hSm8QEJCYKBUJAJtdXcYQh9sAmsPFEm0Mk72nRT3wmyoITIev/N1OxFWb4tyuvLA
SdfMH0RKlZ5N5PK00SLKZ/8fNV+HMD+QQKBKCbEi/J+G4DCxY5fyeTcLW+6NhSL8
vUkWCg+XMcd9RbXnGYIihMt1Z2lZbeCfHn5iC9+mNezbATecvEYnSwwZGC8EEipF
w+mL1Ft38a2YVGwT1FYAsiXjyrs1w2h4dTXm5lehOoG3yF43dnNOZNT/LzmQCLGz
leusU4cjty5kxjs4FKacgmQ3qmNGOyIoi4u4CIAXHeuhovQozSvUu3USpL4OcpwZ
z/maLcZHv1qSup1gO+9kz07nf5+YVZjnhCIemV3ysUtB9uCdLtQI2FVOfa2YhozT
TSOldqvDRBqhBPLxD4DNQ1w3F/SZVAeVs+gQ6/TrE5Guwv6qA+kufOidfTfHevom
ddbea79/Aw8n1L0qFI2QNDR2+sUALijC7vON11+Mb7N6MXnZXBMPU3CBHNPYJolD
j/9Y+NA3YBzUN22r6TyNFPk06qybckEE26hXEj5sox5knqt/m2kSeg7mJ6JBl/bI
ErwHZ/nj4bymLB7qdrKA9qR02bybotxmUysLPHtbvtHk4x36ss21cygFC9dMGfCW
a9h7ibrJAkV0nhmfEkdfiAaqoFgmIo6G2J+x8XiAjS7779nCFjfLGsGsYPcR/qSC
4h406yvL+JWhwrj+2BYBVA0bPcSI2VyMGr8dICgIhOAp25MzJ8uOXTMLNG89DNYN
yeIVrEO/v/eKTp1Nw0SRPHxutu77d8l9k5teSq8ZfKRTdrQWzwzi+Hgs5mht3iNK
TsKkpz4GdMG5uSKiNmRq4RNo1orlI588Jf79Vzske3mwNSS2LYDAC8WGAfpHN666
eM3T7sRbshImDb5h3hRyK+NitCHEcBZzIItDCHCf2vQhKiJBTQObqqUTep8ZHRu+
9IZQXK3akNaKPpN0FAQGC4H6g0kFwgRSLGeWMmD5DYNdC7rsSqJOQ3bqKq6h6Tdi
zvoh7SijQQhCiPT0WWcgYv05LUQ2VP/6Jbh2V5FeZFQwNmSJ3WBz/ydDMRFN/3Ww
nvW29W3rlgu86blciH8QKBCjaPb6FmuEoGw2j6tKgAVi13qr/ap5CQYECxThsZ3y
5cbeOGRZgXFTY4X+koQ/nXEKb65iLUvrRzFb4gIQ/PdyLHPHRL0HUZQCxp+h8egv
/j1DivVePzQNuYmwxCd5lIjWNnLgD32xB2RBA7169GlFaChSF9YqAsrAyh0SQ2db
wf7uFHzCis5ryYzySo4P7wMPBeHpMHUsC6C8t/k2lYvHtVZnVEeKZ6z69Yxs+XDd
DatxrwWLn4CNRST5m0vEEK+uSHw/UHpY+gArFIq9xwSiy62hYTI9ir5STDBY0nMA
vgL2vtD7PSj20cYgaOJG2VH1XcCLSd31XFGuIY4127ufzpBV8pH8dDQvbJCs3zUT
o8LwlU3CE2GNqDkGksJPRgYzU9st9tUxOgsrkqmlhiaVMtBsnmtYLV5AV0JVpU5C
ko6FnuyqcunHbXnK+uxLnMl2MBJyaUZ5cVMwxaQBhyfEZiTd7+XkKdW4Dvlid5jO
7qGV0n7/j2ALeCtLUGh6YtlRv6PJ/HNOu9V9/ZfZooRFAl1MDolu+2+SGvTSWkJD
ufyUyleKdlmSLVaKQk8etr1qgdKHk/O+bGbTB7ssxXJG7iuszfN/99SmGYyYe5+Y
6uU6hR5LhiSL8XlzB27wojpIEOcNexZvafyye63l2/oVTdfuTo13se876e/2LwH3
NY+FksLQ83lf5qe72t4ITXaYW2IWD0d95vK6d67eSvWnq6CpiU91K0DNblr0Lqty
eT9upTnUEAbPwTVZUl+p8DSRgj85RCQoCsLoXORqZyvYdA4i4z8ssxUzKI4EgdJb
gkFxvGWee5+A+zXH4ZAorRflzj5tf1V2r51mE2rXwgjZvTkuwB6s26p5VlE9nqeS
g6Ilsgw7wfQ4El6psMO0Sm0ko139QI6FF/mjCS20nlQF5Kn3hoWRuiaz6ShOgDu4
c4w4++l1DiYXxqdtlWOdU9cMg8rGq3B60O8bGuHTEcsTe0tcB3q8CdMpET242T6M
p1SC6hWBh0oKgnCv5+NO8XqRonZrmPMyd4w0b87YaPB+PwXj+vgUyJHWzsbmdIRi
hwoOAtZpTM2ly1/jJeRnRYeVsaJCyUuObSTcLilf1Tt13as2xGl7WD3wqhUnYLU5
XRvPfqKEB2iPzohrC8p7pQPdUBsYVtM5AnMLjeOif7iZDtro2xSDaBtjRvi21VPn
ZK1pI4wxHgHZitVtb4Jes+XZ5/wE6C03QyG8ae4a51nAs6YQdOuBUJpelsEq9m8z
cTKoQUtEM/YqYVoSg4insVe7krUYINcg8HVtR21SeQEpDMC85xO+YkCQJHi0W/RD
DEjhGmID1HijNPG1a7aFcrVLXGzkuAoZGi5hydjoUsqtvZrZE5dxfZaz4ZFqO3wa
dBwEUCU4ggCkCOCkU5mOIvcInR8MNlc2W8uvVy/P/ubT7QO/5hXd+1AMwNa5H01Y
HNEu8E+j8ozn9Npicear4M5Ci78ItX0VIkDGn4Adhfohj8Zb1a1JkdFFnuqxMfNl
AXxL9GksK8+36w5QZELoaoqXo4+ed0pk21kOPEbSvmXI2YxIlp8tHtKmHKs+Mw5f
+fIAyEH7g2k9mJ1WN1LY14fOdB80i/3daNbvJtRfg1d6xoUzt9CLEwp3UEYfxqmL
WrInAnKVXHti1bHWFztGnI4sJuL3rz+jmcKH8EA4BQ55o7sk+5iXSWsQ/7tvALQa
9l+aRNURMSOhHxqjDNscWzrfkmjvT2W6masYG8vOCM90D7DwyL3gTrvMPxdpfC21
Z3YqhxHF4F2YAolJpAd5LPyNBkGbH0XysFS8hYTnOfBUK7sb/8PSnke+RV9zBItb
GnW38k7uAWNqFMCWKHWGwNxGCQiAjvDKiPv6Ds3JR1T3g7fO07YqMMNkjlGhPFr1
p6p6RvjZPDIt6eRV+Oy/erjeu6JTRgzeurCLH9pe9ruMj82TXCVZGDxR+g1z0reP
7eWboSQ8LZ3PRtUsGBs7fMcLlLvLEUyuHcYHniFN5vqHjo3SwwHtYQveyCaC9H8t
moxwTIcGAKBs+JCH0bNirMKhC2hkSrLtyr2THcrYyoqM3rJxsNW+wf/Ua1Qgo+pi
RM/2iHhXfsMjaOTTBtwZFYbQ5MnVN+rofNtKzoGB12ZIuxqP8r4ppGuwAUECbfby
BrI0NTsSEkQ48ABsz8eyO8vuATJhADTClyHbMrRSWgau+HTeLrK7iPIMoAAWk6Oc
sKOGhUEXqDbkFaS2IPerxYCRUocPwOL/ZVg/PI7sUOq79S+kl6BHq0VzFHr0HJpt
IKWkXU9UpeW6KLMOMSxvy+7HOA4v+NyLX/6FoEVwYV9kTdZPlrLqCKbZdMD9r502
dc8iftSzF7ifpD/+D/lqf9KbCS1HJV1hUAzNr8q9JcWPryhiM+RAeq6N/sW37IdE
w9jZ1z7V/DeQlJW81u1GSYrH9E4JM3f3ND24fQAUgZJcULdGyYogJj3S5G71K2LP
gxpuqVKvfsOmMDj38BBvvNTfM2Yb6JzJBBCWLuoonyZVQuo3vzeYaRMCiiZ1pdG6
PO6bgommHzfBrCAwOYiYYcWJsaweYzuV4srDwkYQcxaw83I3S5o/qrb7DRt6GMal
Q3qz5GqX2ktzGebLZmSJfd8TrBbis3VDvpTc6tYzcpl8tsJ9WfPtyGUk0OvFwTa2
fxeAxs2pZL46vqMzP/O9blYFc8WOYznWCmmUlkD6TYk/LKulElA+M7I5C/SU2O/5
AXFkATUruAY2l9KclzXOqCFOmQlXZE5RbMpFwCuGiAxGeGHDkQ5Bt9nARXwCkZGd
0F6kRI2r5dkObnvOnlXU4BC/wHosNZDRN+p8T65n7pGy2HJgdcouhyFkWKPr1RLs
a3RHn1czd/mYx4OTls94botIN9l6ssiEer9380hitAsJia2HKcyUN4qqlN+aYey4
MY3hPSRAQmLoA29PKzHrbyO6GdJRK4VHTVzz1PmckROrchPDUgigdkFSexGxFhvK
2Tj62IrRb/4IShWXc5n3i2nsSDC83WseVxtl7FtIy0gXUliEc+zs1apC1sydSfSR
pQg1aTC58FxyQzww+//5KwWqYSlybOVDXqG7nd9OS6R4jyBd1S2S1S23OuooZoWU
LemfdexQJZG8NPAloTS6GJ0DHoQvBLJ3RwDFbKBMEtL5EvbsGDcpfkBMN8SQm0Gd
2ujP1quS+dM/kEY/ed49oLPNIsNQDK0l7ligKqwLTxczsimddacjYciH4IGX/T4/
f56b2gXcRg3KT0KI8JRatvHJpiafbQZwCWcQfaOJuO6fCjybTx8sGTV/L8WZn3Th
VIMvbNcVrKMJs0MPS6aZ/R0jjB0nuU03rAIpT/ycYp/7nwSoNPwoscSJFu33iRGh
gAJNX/y7mFrmKL472H1RIbzRbTmfiFjNcJ7VB/XCKQInaht4nphyrMxNhxVSaUbB
C8xK8hdOy42e64RQvz9Q3Lqx4WpGabNRTuJwN4OrKSyaagveHejNLSzhMS9KSXWs
h8tua6K2ibn1dXKGIRFYTiRkK5a9KyvBWH31nR5B/rrvIeFBqngdPpn+yfdxSoXD
B0qGaI3Bdh7/RTVL3YeKumWhtKnlEDaWlEcmH9ZFmNt818UmpaUUgjJ8XkBNnYOx
V2KVSk4vHWo9VNhtEQyt8GLh/7aYqLckxZr6vFLNXGFmbG+GnWxkgxxC+B/1U5b0
soIs8tmFFCuPPdLOL4IlilZJytDpBG5tCDCYYkrK8JeM2L/roWh+eyRZhPGQWcVi
7yaTurMX6lOhcpOcjEc+KEJg5rnZB59DbgzY8ea00jl0jbc7iVbKnNLwljd84lQF
6urnAfirc3abQVsasYOrd1512LIunmndHP38yYRWod3S0XiEb3dwV5MYiQQMX38g
t60UXpiq5kyqqNOpwnR8lLZ2rxhTsIfCmBesChCSewmnHjC3h0n7kBfFe8S9Fe5l
U48GXoPiS7sKHRTZxiSGkaKCe8QbJHYOmbefsA20+3m5jHugGJtkbSlmpiCwD6gd
4Tkt4xLvHaQ1mBbVMyFJgmpmWnhgteRfNRxm7wSFOdS7OrSWpkYDH57G6Khu1RUe
dUzkjn6pmlO9AurkQMdIZG0bjUIhVNZBBsidBu+tBJk5770cJwZzaXIiIrv80zPx
7TdQ/bJZZ/Z/TD05rQeOPTs1Xp5CV8FbS5C75rqKGMAmNwlgaEp5w2v/Q958+nVd
+pmM/QiuDEQQtG3WVpVw+6UIv+OTZZi3YOus6Z1iZ6OzlMhHhrWaV5wp5WPqU81v
nUfTO8uF6vvFlGnNDBO+nRU3EDbiPSk/M7cgXXxqVWbtxfN0R+MLiTUROH5IxBLn
cq+JyibS8+oqiOWkRFNuALw3Kx+ZaGobb7NrAMb+HW+c0U84FnHxxwMBm+4P+vWV
DPxEqfI3XeBGS6W9PY8K3H3b4dkCJzMbEjAOMExP8KLAKGbMAuTAbIpjwzeqmFBU
ygXVpWsqbGv/IUQ3h6foVQbJuPALBEzxnKkqxNNpH4Hc0mM40ozFn4GO6CDnUqbx
hKcEl+IeazegNygSLQrLMtmsARZHzExWdk2nN3fLqa/oQPun5uSvhJHYS27JzzIw
BeOTOJA3o6SZAQhgcv8EA7MHDinsMu56WiJq3p63mlHpbwlF4A2h0r0oTeayq3yZ
mD9gnAJjmeH8B9tSWWdY7pltS+FMLUfySHDBcZP3EcNK7MEorU63Rm/O1CyWEZED
npVn8QT8XjsKJ9ORkCBqyBFI62n9W5n0ptqzF9nrFc1eppb+xwDvoY8c/7sGuEvy
NKAHCrsxYo7FripBH9BQyst9mMDTbgDWh45+I94n8YIYnjaP6jhvuN1sa5XVcgaa
l5flQCOae443p26BrmuL0F3plmyHJi0KsEeqGn1IZ6A4qFoGWBJML0tU0d9VloTP
kj4zjMrOfEWVoRlLswG1elyahzppqhTlPx21v53MyS+AULtNucE0Cz7DjHBTpLza
QQUMP34Aekdik7J8WCckumaoBugGxTOOeFegMaJnKHsihrw5qwvaxlv6V6HiSO8e
fncc1C7tUBIQyYDAOKn24Pa8mxscF5XmdBAIKGO5Mk911KRpEfo20BydYafphjuQ
er65rkfAG7TsCtJRauItSm3TjVfGNEf2wIxzsFHd57bhwakqWnUaKXWCrJDghUsZ
G/tysfx/h+dj79IhmdwBacDj7cn6x0He5wLNZoFjuThDsbWRElVmOHbKUblOSWlX
7Q+XRltKLhMA8f36dnST937juYocyLPxmBB96nl74ypREFzJnw94I5H6rCV5p2/h
9Cc1oFNtz48tjk+BtIISWi36vm7T0xSWIyQCYf9InrXb1gM9SinGnJFqn90rgOBt
rQTOSwLWmHRRjkslp558E8inFsp/7ASl8a6O04czgc3DcU4lZVugqT73vlVt6GlA
24LHZ5X+76+lwcuQh9twGuELaR39NYTUPBPbPbo0gqM088TAT9AdrIfaKqaZYIIF
4vQTKkkUz3QX16dtJf2ES5qb62PUOKPYj/BCzYtUXFFbDv37WK8trwCG3BuAAJ0u
Oa0gBIz2SPyJz4ftha+jd73szQV51PeJwWsvG9OSa+v1Ok24awzqZ5PJS9vSasDo
RZOn3ncJC7EbOWc78IcIPu/vxsO6Ns20Otkj8vCa9shXPn0b2rK2AOyxfnoTmSio
korC53cv/JC3oj6ePHZY2LiG9N4ib6ooUSfcPu67oiaRNJgVOxVcpGK8rU/MU8uE
dnV4R94UNAAATruJa00Jf3uozA3YU0fkdGlpKiadjLboM3qEETVeVIm+H9i8tzJO
FXkuy3GzaUzIpbJyX1DWdSBUvBFrCS3pza5uypg5xKhbhF7pB5zKBc4s2VPhPKQI
sCxnD2rFkRoib/dpYmcwjSxqxqqJ6/PyfR8jeJCHEfi2xl+8uebrxP2cLPSQOdE4
kKtEYT4sXfHsye4A0FB9fg+uJdbM4k58pNt6Iv/61su1pIj28XQ1jv7KQSToS0Op
o2pO+l/OjFKHpfKSTQa+GuJUHeTkXEVgTzQO8UrXrJDYT+wMj4IpJH5Ns4Fd4MsA
Cmq49N0A9Xn2D/TnjvtY29H/iw2kFzvLGG2NaDNrfrofKWJGRhDgf1ufGvHr2pjV
VCnj3Si5+VFW7YR+FbxHCTquOROB2KSaviJNqdsBllT2r0WkMweJWRGiGK9LIH00
Gcdo5a3oD1Qp6ClZk7uq/7iyiKxsKx0wZc+lYszIIbJXu7wVsJ2+uW0tw8z6BHsg
2ZtSxMgs/svdtTNkjuspaxfZTGDDzjYvw1D3fxt0u40X1Pb127DF1NHsgt8YAmER
4PhB7ntxwhy0EEYlMKWXD2+SjLnKIbiMqubmFN/lf99NNo/WWnOBGpdEhqNyU3BT
6Wqo+xmUn+uqjywZRLu7i8oUOYGJSVa+KLRzYw7MdiT2Y2TLP0M7Aoo5dr25w6A/
+EmkK+0OUBkHi/3Eib028BpwcmYqebRKsG48eiNnEnrKSK8Q654RXJJShxgrxc3C
NEJzCbGlPIxfn1Pu+FFBsAZgBBiNVrelIMgZRZ3vxxaImQ8F0Mh8RqdNc0FMKj8G
d0cqv1md0gfuwTqCnODfcTLMV7jT0vBZrk9+o4ZeBAXxsD0wLV45FZJqzhRuWbDX
nyDxw1/A3W0fos1ViwHeGuKVmbsGJrYuaLxwMS3vxW8CtguNTJp0/0rheBQdGdji
IRUlCgp6qiWHHl7OTMGD3p3K8f2+rTY7IUz6Fz9rawZ1iQgS/onKfUDLWaTHi7Zp
9JFeRom/jILTJ74wEhkjvwnsh0a1oSP58C/LpBQ0CS0c2cgtfNqgnIIAnjAMeMmA
kvUelxULqjsEphHErowL5lCcR0pXQa3/63Va3S9AUBMA1UP1Y2OzEQA/LRmJAD3O
qScbE7oRXsIbh7TvoAi+xk2/i6SGDTWn4w2BWptC86UBm5uCRzV2gxq6Xz2H8rK6
sRf0ZWbQQ+ghp9gH/rqPpJHmMVvz0+KI3Ez9gRpNUBVGCCL6bGGygWQ0bj5J9cRg
0N3oq+lWFfzIGzAVBl3hwvqJmu8ClR2pUadGgPpUc9vlOlrMvg/+hekrGX4H/VP3
4skiPdmy+qm66ln4GDfdpUUwLIIHbQsleSz9dW9vnAscQDk5iNut92tq7+GeQM2O
MWq1JWg0QMXOHHhX/RUE34J4TZfuHfTJH0x7Ljl/VATbIuVJzl67rXjhaspjQaq2
X5ztpY4oFO54O3oBdp1bkvOWUgCTGfKJMxNksdsOauT2B0kurjLDytCUcH0Dhvn6
+hTmgSSCzf6rDykwz8zqkNah4E0z+zTjJJMNd/NLFRzQFRtgSn33iRWRSqXs9MbE
b7kOT1SePXK/qT16mrlCJBq+NhBNIVL/8jubVTZ6erpE14/MfNjrtUVz+5YiTCLk
iW7Frk+HYofOXf0gQsXafefWJo4wEJpZzVhZursVWdgLSCUi8fPehOwGP89kBkAD
2jR1zNmbDSvnLXK+Ibf0xx0VPgNvswaFQ/bwGHPltHbyNKZ4TJ1Vm1Mu6BxwdRPi
oPz1XE5H0XqWU7Lrito+LJmv1QdBrUW5/UogGriLZhJxcQDri1WlSthtvwAmD0Yi
rS2t2WbpHEwDBFOorypEf5ZBeaR5Zpg82/Q4DxZ9r4sYUqS8ZGn8aUyCq94/dWM/
Zv1thy4tWjCa2+4MNHYubqf7wokqv0dmh//8ZivOIC2jxF4iOngHVj9fw+FGMr0e
mZgwiMq415xTnOuxzdv98HWkH5HgfZnna6/BCZMb/zHn0+W3GPO9xqBP/YhbGchJ
pUVFZK0EiHs/WSXAxVBL84gEkJ2AOtjAE9K3WlQisUKLqZYhcnNapzeQZYknRgyD
be+8iIbtCqQ8YoAOIcIJdaxCuz/e5mHgj7U4Y1CXx7xVWt9hNsRz/EzYRM1v77lo
f/7ZXLRDhcorSzAcyo+qTlap1uJ+rzSwB0JVsrKj853/yn/M0PNtMPtAY0Fzyl0p
kOYnxKek5CerI6DqyTvlHs9UKWzuqgKBAX4uQKPtCkEurJlBgcoRw48WkzP7Lyj7
qwgaLQ3DmNtSzOx2fq8FGjPhcuBOUaOY8POaTgpzfH428yd15X3zYND6A79+lj1E
3DODXJhe82KVFd5dzWDqmH3nS3vBfnpf8euFNoDJDub6XeXSRtF13FkB/xTEXNFL
BMZIa1YG6rBQWbwm+1dfmUkE1oUA9WSuRH+x+AMSyXnaaoV6DT/My59GNZOog6BH
M6Gj6cVsgZ7rZUeq9GcarLbX7SmqqHk8HoKp435lTXTqFq9SG2IUvM8jLX5S2Oiu
wBge5s99bVE0+rzLDliCIr1e9e6KG1HmToOTE8PFK/XryTEXjs0RImkxb8Ogj1R9
eugKTKl/DgzO62PIArU3ws7aR9eJ7noLSA1OtSsQIA2qATKccgblJIk1IFNS9I0h
xfkKE0xrf4m/ZRmwvWm1+BgF8DHHt3G9wGQDOUo+z/IUyZ/ZsfwkuOzTZWWqUA99
7XpT0HEBNsWNCiYEUXlBYUTLBvlB4vHqDBaxzqj72h/K8Un7/xIsB47Qw7izQsdR
za3TrWQ79AhhGMwt1Kh3P/eWqnufZ3PaKmn7D3eJqRpuloh1AbnBkif66t5h7Wii
+g8rZXY1REKOCYMIku4zkSd0QgX0GPAZipzYNSQgfHJl93QVp/u/k2phky6xbGEj
64+LShdP2QBOkPdILFNXSt9Z66gQYHhaVlXVVv25UMOAQ8cjNGEAZ025wKkzC/vP
lV5QwFdp9MRI4+qDlPohNAbd1780y7crZZE83Cp8feBKJmtn4kCx3BJ3t948dAMw
266N92JDpPWYaUe0Ng5mQIvH1/B2mTm8UW0++wNAsHycB4fuusu0Qhy/TNitusKv
VKKFJqLNkSPsVolNoA6n0bEGzORJq1pNhxGe/5KR72nKnWyVOy5x0XJjPs3ZD9n8
pXfoQO6JIbtJV1lf/JOYnCKOcVGPyWO4WlHFyvbGftOImOqsorigEXwCBV4rcHol
Y9ACs/A29+LL7Qr0OPGkI7yKOwdo5zi1GxPROkTv7jS9hbqt/xFVsgMLfITY28Lm
ZvoBr26d4E+VKU4T8vnNi3IGtbFT5orZQiQxEWz/EIWjwZL1WGPPAVYRcVQ3bzG+
c/6i4HmYOBvnYqbiNo9GwlJg4F/5krWwyVQ4aIQdZyq2aC/e1IT6d296g9m8X1Oc
VQHchVEtjwvn66Qsc7TalRBHeWgoUXqPjodDJd1UR/GjU+PxbHv3jZB24nxkioE1
nG/y1xQTcQXeNxZa3VFvc6lAY70f5zSyZ7uaRnr1PcKn5XxomWghU7wXqC1KuQo4
fajjyzPoydvbXA0eChYlLzpXw47zwxQEzonDwhQ8Gj1VKNG2mwCD1MzyJtxNQCzl
PgjIDjpk6U3qt9n5U6NZ8MvEJqgyWBWXv/xxRiSk6y1rHCGmqhGeOE59pjyWo3kl
+vEALwh6hyhZZ3887nNUbtxdzvTtawmI7KH9o84vQhBnRrpGYic2n1ZPSuNDPdan
PmmVmxEF9LUSPArXB/sBPC5Y7XlI2thraZyfVYeMaSe4Xthk5W8jLJ3Fp0861wrT
Dj0poXEmKa8hInSBKWpw8ZyqDGfRDPww+7TW5UpMJ2NLI2pT/Ts+TEmMDYiw3UX/
TgQjheNnAakFrdpdI8CuykVv30FqSpdLHrDt1GHJIPowxAh0+DEOfuY7Nrf4wn++
n/iCq/xTfJGqOwcAiKqLuRXy3LCqT9M/D1V44nI6UBexdjEdmMSj/Jr8NJqme/k+
wu6DSuK7ggP2xA3/q/uVi+IUQUZxtJ9HLfMkfa7RJU48zoenHzCAweTw07/+1nUT
5QmOS88s4/xWoUP57uAtm6+dWSDouaInVyoDs8+umNcezNSycz8onv5rNJkTEPvA
UrRNZCiI9KeyphAj8CR/JlynaFTAGITJN3gb0xLLVEAqeXnjQ6M/2ITuZ6bjvzQx
P6jknw+UHD3niBckXLFmLifTFPjIzn7f5RI1hh/KBkI4RSmgzzy2clWsQ2JzE6ft
grNPcQzWMIzDnyWVZACuVyR+lB5ZStVOP7uC9peNmvTwgGYQ5Cn3YNhe/tXMbmyP
3QFi7y3AIZ2xN4O0cNaqdF9j1NFuAUYL410Q5FZal8muLkM5bYpms8ZBuK1U9XvM
ro92LhvzKWZuk5Mujfj4rcPJ0a6RaFdpVAmtC7McAwDjLbr9gvdY4UPq+wvanPVQ
kA2lTqSxOh8fPdr3i1WUhWnZH5oV4V6QVs3jiaHpS3aHNqwbqeFkx/HOraQL0M8Q
Xrh7eAb0wm+GdmRuApGx7PYYiUnPjdZLHrOCG9pXhQGl20AZiBqmt+1xfiQkVK20
bM/HQA/ZSvXwZzeXVJmj2QbrcmRmpSB+jvFAASkD3TzwrX/VX7CjxmUQS+N5ahFF
paxELw9s840Fm3Y3ndEdutewSvoRX8MwFPqB4n22/rxtr7d8ME9YPKIXgJpqOJmN
dm5oIaerH7HUcDXxJlm2yVrkVxYiooTMM0yr+/G7/1XMqh/0nFobGNNHUB3m0RbA
rr8NtPDNjPZaWGwRX7Sf2sDzBjGNyWFrU0rs+NFeLfjBklLY5tpR6eBDz+Fb+INF
Gb7ojhd+DlDTIZ/1kX/sgSGIN+ew6za+CoB0arbP+VnUioiO+XJxkJGjWxG3kzsm
QKMU+QR8FtXOR5WN0ofHOJCwZESu7fMmW4UU/AS5czHc1GYJc8QfJmAUEn8681hm
rzwoeLn0W1RfyraQEWMdvVn06xdW9el6uLb1l1CLbqhBHVzfJyFi6kXHHeFl7hwG
6gfwIIFKsWvhWKak1g+Tbkr5kjJdCLZIs9DADo1MNngbFUF0LQ1bkLHr0qRZXU6E
EWxuhwNMN5pDTpkzkARX3OkZQon2LnOTnpr5+da+9EKlmV4W5ukocgPV1+WLb+0m
OYk9u4zz6En5eZu361j0Ut7LH50ZkIvBoB1XGpE/RgB0LJU+RZEtASqfx8MF9VgU
tvGH3E9COb/7stJ1G9dmQ4NgOSyQu1gk8H5vjgGIfmKXVLQOhlSPrPg2kAmvrQeJ
72n4TMZ81V5GqwBFCOjOEC+u8mVx/dsuXBOnau3di4uTsuH3zfkxERsf6q+idi29
4W+vRGLxbCkmq1lys3BUoUfArRHFxn5gUgApt3WAh5zg95NRzkscwItIe5jw0wd5
CfB0Ra/Kpe017XP9OjUyuzJvFKloqu4B0HR4eykFZB4WwC8sQwoZaTQe1EqqGEzU
jxbnGWhFgMQtI0kxnpIXk111uRVCwf+pkqon1xKH4ZjFk/Z4KAFDg5yZQ3nKJcz6
vhsD4MT2feSx0M6tWi5eJQ8o4sD3Mxr8K9jh5ZFmOuS+dB5UtpeYOe11IPGxbVd7
+tFC30BzvnBoP1bnQygzIy/boXsd7RnMzQCzNm8OxoMmP8Arb+9MHbn8gcdI8N8t
knwhd53PxXnCwaHmwLIqEsdCFPt9HQYXX2hf9+lKoyGVd2aikUO0+NgtfapRhJch
fq9V9lzMVB8b3OCBhnWj1umk87FLF8wDvmzlkazRJLT8GS1uEIq8hStoE2m47AWo
+F5VcWRLTOwnZDcioqT6xXvLH8PHMT8Q05eiauVCGrPWutE4UkRybUWMa1Cb9XL+
K1ddj6x4naIo0xj3HiYOLUJH4+c3asPPzbfXb99fDVRwto00riffiU5JmsklJtYV
GYL4t08iiTVKWaRpZnSgHHcGyJi5LPpFbIqjSp4XzjIJYl3dHjKrbNW/lDCnwyz0
FBERvrlu/IkEQUhhrJwxhAI2Fch2YwR2NJeETabvv7Q1Pjhk2a4dpAsWUSEhjLNy
jUJR17KYTQPGPolwJEeVREUyKa8unvCMovbvO1SeOJNzV1oS8cMkp1bmlXW5c0w3
Gv+OX97sRjqA6o6fW750ZoxfVZrSw8QolvWpkULzEqiOEM6ODcZqglpsYRcjKE7b
prqy+Jt5Kp8mHF8G0NQhg3gstJUalIB7a0trh5IxTkj4qFZCG43WqxcfyMDhouz5
CQdTq4zwEO2jwN3kTZ9XKazVBKDhUvAK1qt1nThMXqwPN/S3ySxkOp43sd3n4IjY
fqqn291FrwKDXexSLGB316PKoaeXKRSE+roa1+SC71Mx9v3aU2TRXiv+Pa5Lx95i
tBYqwSSIUrfuZjhkQaRktU5U5MQSueJysoSZYF7Kk/oRi3IL/9gQYDGo4Ez3nhRK
SXBqZfEkVJMhjnWvYiDDoYkgFVBUDLMgWN/ZSvnbj/MbfWHxwHpEqW6q62yM9Gc/
EPXKy96QmjXSPmlxtuc0t605borp2+NfqxJ5S8gDZv63/Sk7tVpWVJbf9pYcOseU
BhKKZ1EWwOAAU95VmyKNGV1CngBM941yy52lS9pJBUG5oyr4lDpa0y3IlHSFfd3z
CBrnej8y9GUjZKDWXUxeZEJuXfvgKBFxWU/bDmC8EHTpJuW9l9XnL9sV57SU0Pp+
Hewx23wslfBNE80OoiG0NHxHv7LiRxgRzXq8OWa5lIUfCcR4SwWgrDeEOXwalROY
kRjKNn2MFFsfNoKADp3b0s3bh911LX5FljnA8a8WgXK11ZP6q66sUJJZAmvy+vvQ
MpWXSGmjk2QFXitDm9y2xrZETg1471Q2vOKNDCGXJvC+HMYY9ai24v09r3B8FNa0
5Q0ZqZ7FJ7dDkCe6eNhmQIdlh6zOTIT5bSv/YbTnsrdYnztKyNAajxQU4L1CpqIv
vYQ49mWW1uktiamgFltZrou9nIBPyo1iXIi5qhZasHfFkyPK/FISXIoPTL2ZBTjL
1gX78QPVV9jjkr0Z/juicBTno7CtTIYj4+JkCLsPE6fldUk4sqYKMbI+tofFCv68
e0NjOA5+g4RHJ1jjMR74CAhLjTzUwLP6VYFPVm0/ml8yHWx1FJe+1n+7I/VRxLPY
GfXVP7J4hv5vOkgFUCD0+WM+J5n0MJ7N6D3XFIpoCrftrqAMyI9Vm/aKpon1uj6O
aTXCpF1SaprUjwE0DcjfdeqEaoGZ5BA04RYFQ8Ey0k3U+XsCsROEna+oJlzXcSaS
9brl8cLD6ANqCTY2QTQXld8QjAHuvXYiooFN+ZVYTWjCzGEdD5qsejhutBvrTDFV
AURgz9+zslUIlQbg5+TAwTvjg6qQoIAnbtWSS5YMsL5zuPc+sB21Wq7xs/LiGYs6
0AdEwAhzWU+MPqfd4kNAlYU41S9Z/gM+CKl3WgcrHmP9Ij8xbrvWKp0Xhrp0OO64
EgeDBWoTmTAcr4tN45CgGUcj1z2ys5c2yeE0E4TmGjISJfG0mEf2HhcXsHBIQ0bd
euXOGYttR5kva+MVJGP0D8SK7ciAXuOCb1uW7FRVVGl0nla9Boytu8a4j/yx5XMl
uiAHC2JqWrwzCuDHtL3LlkqXKhiocOYdS25Ig4bNulMLzD717vX+0TSBk8JOvkTK
nFgL8n0VtOotIIrPhgCcqKGDt2WHuU1YUNPKH8K5BjGPmspWE0/YM12TfZzHbI5K
n+KXmxtZO8sBVoRfaExCtvT2QJQK+Gn7e4TwYjLfov+AvYy5Y3HZFn3ls383tlv5
fHoTEMkzkjxb95/qP9BRku09FuZGH9f4IENsL8mWJOQTKRwZh59iYHKVqd6tiFal
ChzC19Hmp3H322/zU5XExueUrv6lqSlPy+9Zd8mkExxnLSrnjqg2NoANIZUvRNA6
VFigGa69nNKPJ5WyVFkndW6t3BIbrVG2+oxC6rh4xgD6Mh+4qinQSljmH1nEhGjX
N++DGSi3cBhYClh+mxoJR8k67zR0IRq2XZdBe8O5MDa+BcwMlSNr0jru7FMrMiKJ
tLBgjJzak4lf2eeDmsCeF4TKELYYbhpBUNUr1NlHRivYrfEfhZWYdUi5dr5EeyuT
BS4b6t1IQFUOxB61sAQWVXrQtXWjq7O7eXzLxKCAH3ADBe//sr+ZC5BBWcK34x/6
LbQTlLxWJs/WZ5YnbQWvHYODb/mnl8pHqVrun9erO0LxTjA/ou9ceUCFamzOwCP4
pLH8sSlM/QQMKSOmLW1fJwIRPG+Ll6km14YcXXK51WsJClpUqtwvPPrzWZ+zGNqb
nkny0DaWu3u2ydRrEEbSvNcgs1+JwKU1ooSsvKTDGl2dxcTBUXYjtKDoagIn/Mum
fRGhl9xw/gYFchiSZTqSCjrj0VuGyy+fFox99bjt6Jpm87UGg8gGSvEIZW1TFhZu
0B4bekSCoUqYYIMRBEvVo3jlmUeGGtMmvXB/BYoKf0neaR0D+cDlsqlNgMvoSYcO
IDkgKyZ4wyhMKq0hcdriTqKn9fTx9W1eNo1IuwZjksKNiJcW9EQ/UKT0KQwxyIC4
beCUenHTg28vFJphNX1lZZsmkQE9gkFgsAgjEbWSX7YJsgQj4yYuBJqYnH7uh/53
YtRHwuRNfaH6dzKzhD5xm57FDZr+niroM5jfr006f604yYPVjfTRd+z7DqL49GHv
qRgV0oBy5Y6Ei9vqaM+y77U0IoFojWl+9W8+mNtB7XbnJlS7lyhWUA4hMaXgZw+a
h8W7v+ST4HmzCQfC1LYLwmSMMxFs5P8zZKDC/FUEMAmJobWaNbF0v9qEydMW4uhO
GcoNdZsnLJ//FfnkZmbIGqLwFDZmuJsbpLPr4BM9Gi5gDPiLlOD9lrKQKNTWMRcb
+PiV9CqPf4ycMkIUVmrXoF+ShXJL6OpXw9z34tyG7UzPQSEHcqlPf2yFwR2iWzlg
CgydwwhNkLWRy39AxLhihGASXlppYJLe5ItxvjiqXo5vL1URhpMumzXblJo0KUt1
hDLFb71Q8bJFJIpGobtfX4qXYzuibsBWcZ1lkTqBI1R0I3UeczR1rX2Y4ltQgHCP
nvSqYGHGZo3jiqPIbIM6MAX70y6yQGDXYibRCnleAuqFxBQgj5T9NBUNwMs+e79+
2Lw6D7X3Qgi2hbt+mqoDZtCI0/tM9WQPp8SKtoFEO5pMET8CBu1RmMFwNifa6avx
PnFNkfd3sV63UvJHCQPwSmvLuwPDzbDvnBzUkjMygj1UzejyQrji6g1sj8tKOYW0
qCFtBKym8AUgoL+5FECmjFZy6UoIsLpAgVhVQurWez994atgX1MASSqmPuikwHtv
uEUr8GLFz8QKlBr4HS8bZymdgOqPvkSzVjwICd/s7yV5BNezm0AeuksGJ5wFSvIK
2r3CnGKsUWv+RwE+UD2GS21g5tDSoNJIRQq4SClWmSA6qZDJwhtjmZe5sCdfQs53
pJ9Qh4H5KJrlO96oWwrL2lihbfJn/WkgQfpBx2/moPQrFQ2b2A5GBeWwIjrMmS3h
uKCsT3jCBVFJMYtl4R00hv1bM48j5mqOwGXzPGNrcauZxemT/hHwnAasQbtFlyn+
shugAKdV9XcLPR62pj+cU/Ra6Mnw9eVSfvRu5Hz49Mbwg+ap9+9e8Gxey+5MlhEM
pWyDoPMQMBvqDbok1swEMnFOlo1DWPwaaiTEzw6ss105PFsC+dv4hBOqgjNBjywX
X3+U8vhj7lYpdajEsfvFrviS/FQba7by2lutFeyQHTrED+0eAEti3njV+N8avZGp
XRf1CKAuZlEEMN7Ip/UewOBWDJ/Q0vR2pHxaRbp6rVpRCJ5+/AiLB+PsjgR2Mhk2
XRHNMt4aOXQcm4OS7s2tEoDIpvsXFgc6zgoQedR+nFhHdUkyBzWlchJjhg7OPKIU
31YPyY5xLFKzXPkDwvbK/jbUCaWjsmyS9UUQ2HrjYB6SNZDexw4exW1RzZHnXaK0
hErM6CI6VGdP4+beZsR/toWUKPpVlo61GyS97BJAyZt6+zInxyR59Aj3ATIDQTpT
Qfyf0bgDaZ6zstSFEJAlaeDwYwR/+/MHrG/JvO3/83SLXkIi/jSGgKSXKkZg/nbR
3skil5DL2aQj93gY0ylWQiQOq/SsqZoMIMsPQ6doJoLVbyAkTECXe50nZpZlbtCI
ea7n88kVarFgsj01BBXOl4L5nRsN2/KbVg6zGJ9vjZl+BgWQY0MWXO3Ij+1PHinO
LpBcT5mPbxM3hoG2NFFu4c+y9avZLy8D/vkYVRFp51n81ZV+u23sdKL5koOBb8au
Hm8GfIjDiUP00zkPKhv587cc6JN0gHo4218Rt5L7Xl2/hgvJHZjhLKuTBJFJHiz4
1TCLpIaho0l1KYgbLOmopBLhn72IJkWLmpHBPiKlnoz8PF2jYx1MY/LfY/7LG7NY
IJ0I/6OoDdERQhZcbYjWrUyXNIgo6vKmnHXiMGTwuM1yIwjiIJpX3frbTDC1AH1X
6T69JqpAYfBkTy+LdA8LPK4pfzLIqk0bq1qU71xSIl2XsM+ncKdsaU6P9Vl01EYQ
fl8yBgLHJqdTW0vZD8lvlEs0vFwFxLSR5G8WHmn977a+5nZwsOY2tEmpaO+ahmHQ
Ky1ZbmFqTIysMYU+LOQQciv3zmKYET4G+ENLgpcxvPiMgpuHvO1fz81vyUilYiYH
CHYRNdGx8r1+pmyDtW4X1k/3gh/I8EgrwrfqXFRQ3H5VB2b3S+buRoOJfaNVHip0
RU3T+TMhJoCwINySsuewhjz4i9o42D2UZ97pD/L5jmdYdSrMP2vz6OeKCKraPu/a
KIuHJIWbaxXfzzWKL2ya3aDkmI8l/445ZkwCfgkvxpcJJkJMFkgDBUGlapqv4G4b
a0e0krv5nrDL2kLT0Z9qgKJB07UfgMVXSZhtiwWWr9HZYlfJC0H2oDdHNmKzqtLi
WxE9hECMk4C7GHQBU7DoHejmFKdcJ92+InQ8M26ebCpBYQ3NaGHmmKDHvyIFMquF
EErW8DrACggz1Csh+utR2C1xUbLpzZFbUByD2WqM2kkBaZQW7zuYL4EtNtlpPynz
b/8aaQEdIi0fkkAKQvePa7q/h4vB1gNe4fSNwxZ/pCAbA17S9t63PaMwXi7vuSRB
mqIwqMf/bX7EBrWl7EMIXEQGX3BIaQKxuXHtvXpZFcDCKo4J8bIGwGMbNL1XDNCD
AUzocM5QgH84LVttdqE6z0MQea/wf8Dt1MuC4O/eneYOMJi7z+/kkrieoHU9otCd
dxfxVetmK4HMfxpZGIW7d7HcnG3PIMXa5nIBfDkEa3OXTLn6AzPWJyLgmka2Vusd
rzIZh+H1GSmpruZ+Yf50u0MfCu04/KlxduzytusQVEUhtQZJwkD63FUmZ5Yox56V
pVjErTSY7y/BUEEqW3knpAzSanTssVuiXz1F9XgJwKZhLaD199I1ZaPbLKDUwWve
joqJSP0jWAeP4PwXPtyr7dsAnXWp4grNA25UOLkmo++Ud6/fjqMTjpZN+AS602fN
e5fmFzBbR4BIH7GBnXH3irZhTKRZTcbHwA7H4eVDu3/bnB22Mxf5ggFSN61AYzVq
OVQo6fCPpel/X5XXaKzZr+gS70vCFRvIDdn3C4BOF5jpK3VU/Yo/QgQvATL8Zxfl
723/kQImxMb8zWHaph9bv07rQ5FpBSW/8y6LzIypfGTe9OwMO1n/SGIGlrOiir4N
rgb4XNxtaCBRao5efDI9pnKoyHV6nuCkxo5llWL3NGpITChNWsmWVXQql45U9FIV
V9tCz+6Fv07YNa+9tSYqNs0FxH8qufN0/tyh0xdAzv8EMKn9BkzWEGQ6q4cKXK92
4njbLess86i19JP9drHGH487JI8HB2M3sWITpyLlGEkcJE3eIPq8yePUwi896T6g
5QHe9Oe6Ti3Vp8RzZc6mGWjFMEBubZmHpzfnoQYTbn0UQsy4heaCAGvCHNhNVR/Y
jiRl1m3Lt8xM74dmXRjiiBtsAxjEFnAiV8Gf5IN6hgY+SwfXG/r78PSdkfKbI7eH
H0QcRLXvq1R4hQOmQmmHI8XBCcpOSRCc6ZVfAb+Pjpgjz27iWreuF+Z0PZgcvDIX
WGU7spj1kSJHNROzmyvfGiVGogdMKsjAdcY1U7r3Bb8wyMFscbZ1kfPozJhKRhDO
VH6IcQKUZykxxtBtM5ZUmElUig4bD/UTE92S+G/4gtBN+t7UJOYBtm7zHbcwKN6l
5IGGqzb4zj2ZqSwK9IDXbDD3orgm25L5//+LkRtKrSngtEOdaTdtX388zC66vijR
lNPIt7G84EPTkT+WCe8c8qWmwz1WpS+yAzAV86BIu6zSEoFnEOwowDT0nFNCJZYp
o23wca4l4IrTBblujcmuVHbVP2uclw5tJUfatNlwKqmNehsK0aUW65SbtG3t+ROP
jXAqPS99b1oFFF/6jJESfXJq0iKIyumSQ+8eEYE1OA0/uTPwSSGmCaC7EYFhPP6l
iMUk1i5d4qSxD81Ra7b3oTXNeYACdPCdNxD+kHDrJrZi5uAOLX1lsDXT77sIKj1E
mxFTzGVxbm4HeP5Jt6ysqKVgXncmb/D/FU6VvyHPT7CjX1RWezBk9r4x7YlwYdLE
uU9gxRRfl0tT9j18PM+/ZxAd5SilSVMSdwdftLK29w9ooX7Cj4m1nVa2ooLrvjrx
Vo5gMNWYOKQGVTIPSatDF8fg0jLED2DYbrbgdmSpXimRA7FZemPJzV+lTAS5K+cL
NGGx6N7FS8YavoKeqaA30Cxy+9ylLEywWI0P++RENRrYQ41JHSwBnHz8ZE4YP1vV
klpVfEvhk0i+Cay4Qb3kTvdHSqqrtBuAlI/WFs0vEGpcbXtxc4wFrdR/nCpotxMg
ClVDFo5ZtwdWlwi9K5eKFpj2gA2iusiRNDfw7EKTZGh1MQGmdq7cbmh1RxtpM2HP
nqnxIS+ZO0xh8fRUqiA5xX6FxcBkGlgqSJR+CueQEbSoIP+fuSIgxzoMzS7ylel6
Ykvw9CI/qal5jYqq0M1ge86tG73AIODVb3poSpt4Uhm/W8tzySh5zF0foAU55r2w
kR8eAfNVTc/5+QhZSRFCnKJefXDIWxAAEfohgC4tlXVNueau3fljg1HiFA9iBjPa
4gGAKltXc0CCIHbCXe5r2NsXxaWdlKBdS8xfz0XU5xbpxPrfYJwfsPKE0iENF8+p
zFKgTdyuNrGzYuOXVnDYRaYObporzneRVGpvv9Kwn8ekEgDTGnNqTtxaMeraH8oF
kR/DRZCYfZxGNh/gQ74KcRrLryain4S6cqRoEe7+wEWBciDjQM5IojbmlOlAjj+Y
24E7z5puWQ8dhSt01CJAGzYXb0eITu3ZX45QaFc6Uwx0+7mhXGE5Po8MRbZSx/pK
WVRqw7uvBxKwqAtFCVdkiPUiyCg0ABSnumfHOsZDBvx1UiOPDq8UKkhWYkoZlLUY
MXAQiiTchbhvTTiK8JzRY1d/ejswL+qSQyDwtYB4ty1eA5TAJQi2FNNNYKDHJTix
48A/rRt2fSXhqRNRpc9KHB15kNzqAdlcxvYRmS3MRpEJsWoEsXdMzmwY/Xd8HFnz
WkKXYzCIoMCbsu/+lvMotBg5loEDFrUUczRlAumbIKbeB57zGgKN63zC1zOVq+rp
bexSWFtfXMfDuhy84xkWVFGokvYLSGNhlZkn0J0Vvi79fiot8TREjHylVh1Q99G6
aWnlRYGJUTfZfBCeW278aRugFvaX1aSRdbYR8TgO0FA62eH2tTcWr6hp5HrSky1P
I8PwO9g9vY0OEQkpzq9PJ31l+kdqIveZfMS+dt0mc/JjLDgFM9kB7oUPWY7oAUwv
UtdrD/3y15WfA4UQ1K5NxM9TDTtnqYCwbhcO8KVWOPPjH6+UHjlQo5+OFofdoGDA
H/B+BSAhM7lDsCOUeijeIl11oHTYQ7mp529GnpSaVOwGmY4nwpJKfKjxh/m4jrKI
Ec+4WcEREMWazkXG/XKu5pPCqKb8FLjsbyCusMbRAN+WAphTz12HgPzky0naY4qi
X5gH20zVBaVlI9uhW6CYC32Ml94ElVkjhGZ5OhAevtbgpJrfZC1V5wfawVn/1Wgu
AlocifS+Qe+sGD8gO7tilsBT4QnTLcd9HvfjehHMeNoA43i+j1G9pC+Slbj87UXF
QGDQl5cNC5KbdZEalLcnP3nBqbb9SdgGLZsOqLfZSAyHcPVPMqAkDCTZecGfpSyH
zrfZD5IPWU8GrzWL1jmnmVFFjHvT1F9lP/55Tu56j7VIk+me15HWtu1j5YMCNVSY
6TIhcddBcYpgIFZzYQhiqugh+l6tzDGTn+qSV8fSP4otCrg0P6PXExequyABQBeF
ja7mwLfA1BOMpxbHNmrAqsUS89Q8UaxMn+iNW6XmAYLLOVXWkawYcqOwnA2BBMjf
+j8d+WcZwbRrPGFI1xfZZQVDcUqjSqodiF2Gcq/WKXhdUPD7oUA1/9esju3LWlEq
06/I0Np+fTDopfyUuIsOCzv20nURV3a+SSqDy697I1vpOMHz+pNkLK89icN2fMDl
qEnsEh7vDIXqa9F3lzwpgOEqNqdTtc+AO2Ojyr1ZcPpw1DNncHE+PR1N5vWv5NKo
qvsT8HyI0b/6VsKoW+Bfbe98A8jKD3D7qtPQpbYJrHjnHwlWcqIOE/miKCmUcWqD
KkUMGKqqIMoLkIDk8mUM7/8WKN1ZpRr+QO6XNTFP/aBhGw2YpOc5tzA0WVVz2+R/
FAVooyH+HRf1QC+o+XxjcT7RrUFC1JkO877hsFUmCdkMHPiCk5/vW71MfLnpPNuS
6yy5uYSG9bjYCZS15rPY1ohxw96QZHxZBVj0BBvH/CRs5TrU75wWjIhF+jAY8qBl
jK0x0nWwuTTI6eqADODyGc2/TS7luqmfM/6lirCDScddPz6PTrdzJEFYdpMARoBr
KYytguEpzAYBYSmL+EXb6XI9SUqRuKjfNQT1+1nCiAInABfxUnbpyzpUymrDkKTK
Et6ZVeqY3+UlSN94uRsu25Qyb2a0Bb7PkSVHv8g9mhAaVF9ajNF8br//RlWrQXJ/
a914nSgW/hCKwYPISYhJiS6tVbiwfgzK2NUIEonsMIjPiGevyrNDum7fEk0dqdI3
EWoLLvRQttiAp4GPHEhqiOE74nGt2yFEbEMPu7/K3AVJBDGNUQH0p2KoRYu9P5op
Hea/CJ3jx0jun0AU992hAsAXPO3ERr6DByu3CbtsXu2LaaDzKVR38YUqs3MT9Wes
d1QFcyZSYvDB0PYxRnLCfXhMMRiA4J1gaPVcqz6qzPBmskV0Mds1gyAxmk40pLqg
iNxJDUaXV76iy9MALczunX3Jgm7dBgQNNwrD3nc/gdkpg2Sc1FNFghFeasQOXQTp
dD1mBZ+SaHbskZiWE9Qf9N+uRrqtEJCr070y3E5V3HfYbqwfdHOiZWJmVNKG4zbS
8pVq68LlOOzyRblGMd7YsHTisie8Ban9rXNnBN1DQGu8SflSderx/oBl8Xcqowtk
hgqoSYhBy7mI3Q33qRMJkIo/yb9qP47xaU0v0MYQVkt2/nZ9XeP2jPa3eBnxAcbp
mC/d7s/TZ9a5S1XgOhYjGH4MuhQG3sbFZP+NsQqjy4thpDEaWe5QTpdi4uvk0rPh
gUzFBxV3kW4h57W/EaDO+ln6tkPHHosNg8eIDkmUqUlA8puiHqY0q02ZcHvXr8Ra
NRniLxqTjzK6GKTVxd0JyRCvIaa+h34Xqq6flRuij1tqfc1nPrMIg9E8qTHHzEVq
Vri7SlARfhEbgqUz3Mzy79kUJ3G6YzOJPv4GAFwe4eXMfitW1Cu/y2SNhXTXu7je
oHhx3NLFxzaP29X0InAJvzSK3+i0xbD++qXgpB9dbFp2rv7+wv8tllizuSXoBAfs
w/yYCTm7XeylqCGul63+N4hfEoShdI6DYWnUn2S+bmWYFV2v3OELrVfoWK3d2xI/
xCs0hSaEjMOjtdcobjmp1M06dbzMFprp9vXth+2I83ZAoqE4uNVb9xF3SFe/t+ZY
tt8MFkkttqEglSOxL/WPKWf30WX2B3RHct7Fs7AhYuJWnvc/bE3KkWfezpDGrWQb
ypreBFmHwg6+NRX3n09xRS+XV5OHKYU2oAUVzToe9Rjh8NfDjB1OnaAJDvEpOpLT
g5MvS/daebrY66i45mbmd+7Cs9UFWBI1E6YQVHeJJI3rLwdr3IPpO9GaVPL6w5KD
ts+fTT0mkT8eOKqCvXyc9ahV2HGtp3NXhasB6sU6IbwsGtY1mpTxTbPm8Tz6XYEx
QRDWDGAghzznkIvTL2PvTKTjxGsgzlwfabWFwtb2CayAaJubuTzE5YqGcAWnhERJ
HgwEOxkLBgwThFskQQIixwxdKPRE/Op8OiVFHm0+8DBV7w5BOYGZ1QX472BTiUuQ
JamssUEvn4vK+0h/W7UQEU+EJwSKQR8rKNliNpfWwgc75whQansv7Y7W3Gbnim5V
grk/AH+sMyk6jATTjtb7DssZGGnGbQCQ5XhKJ/45CLo1D1tbfqOCz5sFt79cXI5t
1O37UoF2AvkXQPG0QYe1RMnf9vASstd67Xk8p2cu9VAgXqKUkeaPiG9fwsC0Qh29
f7ssY8BnUVZcRWwfANGi/S9zFS3c80GqbWWxrt+MPTZT0qaGXOc9quqKtK4nsjsL
TMdvSiI7TfJxshozbskN9imEjuldQgHlUJTp5CQcW0wgpAcOIqw7NBnoP11VNVKA
QT3+x7uqN3BKNS958p41IoO2mW1JHB5LkTgmLX5X4pv3ddb9yQYsO2GPgOp+Hv+j
p8JNT74t9sRadFbGOgy0lhS2LFSj/HCP1ZVG7wxUlw3/XhtzobRXLn4Zcg+Ck+9+
BHNnQszSpGdI9+m1BVHIeIOYbaNYAgb5jqC4XEdaEaHDZjtSlJpkUXBryUyReD09
tM2iLLtUOYnDdQsUlXoyJo4X8bHhidMayIhTRlFEL8Do8QeeS570JrOZndeagHLe
c8vJIB+kB3KwZ3fXYdUGrKO1q7yNOWjUJvWVNwHV64KBip3ndkbCNYuIM5yV2UfC
iLcgYCysGgcl3vbg+paQxl7r90Q6bifoM8Tv0oysj+/tcLxI9vogNXh8hMERB65C
I5SW95XMwmRgfz0e6zuO89vDM/upyOtJuP6LwSt17TgQkA4iTc3zfgI6BjSC7xAB
l2oykdtr2AmfBJZJnAk4AgeaYP2H4wiQNAcFlt55xmXUaDTpOSnwo5HQI+CpkRpi
7B9wmojzy3Yf7EzHMFsHuQ/Z4r214Q2/NO0Ke+AoLM3pOb/Ey3SBio4L4bn/4UGB
0E320qKod92Dta63enK2S1qAoO7wf2q2iiVC+kmzOFoFcR9/tJBpAJElCgkEeckP
uPRA00qdnSyAjTHzyfX9G4ZOi+b1h8pHvsFOTqPm9x7Fw6hWeLBjSPUTggYdGX4i
FGIaS/2LWrQ+SFYoVvDKxow2zXK2Q0xZsQRcpRKca4GAnksMIdqlpHzf31mayQaO
dwSSWpZWRoH6Z+uqTHpRGubQtToxtn0vGi2eUAlNApZ9BunOKEBj+JiQycGajFNW
VKbzqanzpjLT/yyBMQld3NZGoGsIP6mODHiFjzvr3c+BfhaBbvo+BcVwENQRafDI
dRQLjcI0W8nnhoL48Yu4XFDgtBI4l3rL8Bdo4I7NB37dDlq9dkSvg14mkFhzKnxQ
46U/Z8rT6Jx9pUtqG+6zaUbK2o7c8tmQdgbDTgD/M7enIaWqQA6BARBtwxR019Jt
hGGq/A70ja02MaBKVQA5h/OY71HlrAQIHP8SUJvGJanLMsiglH2zscIFcnNQgHNf
eurT7+ucVMoqr38Cdxz26DbppzRvmGjcdIor9vakVFlZ/VA3gv7GX0tCL6sSnFea
Fb5Y/ylgcUO3wsyILTjac5GQZLL/BKDiYQSkoCjOpEtlajuKn24jFnVqDGG8XK2C
aRDkyBJJeE92Ny0zBA/S3ZXjU5wZcrTFKhC3baQ9J7t3Q3KFvrecwg152CpQiDpy
o3i/vAfKAt6ASsViAjHWN/u/u2AXI5tNCebTCZ54o6NboSBC5bBjEfjS4dUj6NR+
Lc+EeS9LWmrGPq7aRAogw9joCEdQWJZMMhc18EcA3Cws2UjiqRjopSphjnLVQr4S
9UpOyj7vzX5haXm5S1j0aZKDC9xHN8ZzjISzwCTx9kDhfleutpqFvaco3X10q0Wi
ALOkjWxNasys1Z/+n70KLk5LHF3CUxl7cf2L2ECe+ufkvlvBGGLUBIzxqZ2+SnRe
iBXLXTkWmEjyuUc9zSAvijyLK95r2xZwRLKMJfdFr0bOQ+x1E8uXRCw/MBmtf/aE
MfDuNro4RdYpK41UD/+KXJBeKT8H7mogwU/dmstKTFKcDEU9j3ra3AuOunwlEJm1
mXz/ZcCXC5HYgkPAHBJ0GFSNAdavo+uBfLpkXO7keWK/KeboQDdWssTUtV5y+eZU
eN+tZH4lSqguEAK/bIsDburvAsldBRajJhSLMga4Zq7ySaj3VKI4ClY1A4cLSJ+C
gDieXJPLBy8hcOqsoCmVh56J+Vr4iFIuJ2QGoUa+sM4o8g3FJtYwvoz/gah6J5LF
N+Z3YFc+kf/3hrw+kmRXBZYqmZYsEZKAuSgNZCf6nmaI6COEbdQv9MUMFtH+Ijs6
ThBZ1rFCHanTudowIycHvUz4W+9oSSSFPfYWnZ2JaSPzeHCpxqNIP+T6L8F+E/x1
LotC8BDnBk7YRSSX7NZS4NSB6kyN+aq3R/7mQnuObAtWjl3H5SeLzxXN+rWyJxl5
dWz3Zg5lIt7bpWljrUyUXlh7jEyTodG0GDU6CX/2k2xMmozePEDwZnFItgQLIZ5D
+S+3UvUfx7Rc8D+4sskc13sg0LewWUNgYSlwusH330XzfynzBBXXMR7TRaVB3cWY
HcNNoO1w4vSdpViu5UIqcO1ZLcl9keNUXmHDC4IN9v3q1BeLN293u/FZNUKDSPqe
ZN30lCQ9disiyZ92r2fic115we0ZDC2hZEQS4PiKM1wPV5lOOz4n0bQcGAvc8Fae
MAgoZgoLv3leTDzxmS9bzU8J7pCAcWmfnhReWTGIPdBB9xKz8sxbO3flSS9Zxxiv
dSthPukGo942shM/i6Z/ck94WyIOq4BMnxXXjOYk2mF05KEsF3NbxOsV6tt+RRzK
37weQcYbiQ0zR3/4OrHXRuPapKXHdHbLvx0Dfb8KU7rwRbQyHyggbpx24yPnPbYP
yDTKQZ+34Y9hJC7ZI5mLr1ZXvuyo++c2URM3oTGNXtB+l1lwNXw341/oB3hur5QQ
n+vPWViwpJk6gfL2taPQRM4NlGuQXJKYMBN+A9EaWFagYbtOi+TJ6YSYeVAmVOau
DXvq6utFLEEVYrSg3hPfBOmdcg2omB3AUOJ8uKhe5w2H5RQzqsUd2srLYV2kSfrW
QrSdR0lwSJC3Z/A9fdvQxrGP8kJSNbKMbt5YFSaNiXnMA5WKp+quUEvwK65bJduD
i84DgRrDtBcPVvE03DgG4w6lIAEYOTOvsgtsW6/Rl+LwAJfc5IWWlUMcRV8MA4VY
xUXqBwTSGDiNybDudHf3C7qVJeFSAj8L/h3h46KiDkiRrF3C/gFrvO3AHjfQhgeq
TrEC3BHZRQW0r3SnzBJ1Sxl0HHmSrgbVg/k3erZWGgPJQZEcBTJYqG2VML9ldEb+
geo5u/AvuCH0u78t/+sDzVVKeubIpaqVTtEn0w7KM6W5B+OUwat3dTtkD9q/3ds5
xGZbKzPP/61DSz7dUS7nZnOZAZg3w/aO8u8fGhV5wnVdSyDX3dev34/A/NFmJnVr
ovzxl/efJ0tub59mUMOUsA+BWYvtoNWc97CrA46qr/AKas8WI5uLuj6P4XgDJUdJ
Dwigwt8N6gD3+dxVjAVgsMKGsTd7+0JKZRdEesIIgAh8r1CgybVv3DVjuedXrD+R
Ww0NPDR6mTcWUwq2++s9XmkTgRPPW6Il47S6jGLrSqDuOiY6H48hN0vezspRzUlt
Oc49J4O6o2b3hRRiJXw4ldD6XVaGSlHYFf/KgeM1Ba/AquZPdu+HPkgbB9wS+pxH
Y3zOATuhPwOS3gKMOpaoFyKAKlztExGXnz4KVSC3ibigwfK9Kkz5sJZYJjKJXSV5
MVuJRSwlwg+eoXR0HKxkbJISlM9bfTtRU+yNPb5LhRxNCdGI0QmnaC4EVxH9bMc3
dl07dQDF2bHgx7x0GTfBNFjiQoK/Rx5OcO58BwQyXjEAEhTlfab9MkyrpPXQ4Yyr
EZi75GayTAQrBAEJoVIevS+S25dU/92lfIALSeMqBh2FhWLyykvI3hp3ONkOiTNC
HhiXszypXeF3XB25zHcCc6veFok7LQNHOrIU3udS7VlYqQH+KL3lG+WDpGzpgozA
DdcyQIik7d9OKQc4YmjSzYJj7YDzZfiY3YRY/fRaYao6TaNnRJcBNzMPa+rkDqG6
Zq50qQuTa76C4WNtou2M+0Ch6ORaayw9hLyU7lEbgsGWsz7c3S4V+e5mkNYc5nt2
EqapfQLRFkLqHghc7EI1JeLTGS2vq/io+57GwGBiZB1eerjaACnCdSD4Affx/Hjm
H4Vjpe79V1YYlaOixNuHNLZvFOdH28pPXAJ3kFQjut/BkpaoI2+YBfZ/CtzsrZIL
PhXIVl4ZSk3/Jx/w+TZ52jQzIzdv2cq6TZzU4jVu7hrYc3LwWXXTKj0CXoOsg4NN
aFGj53oq/Dl3v2wJ89qVSzvDPhJF4VNgxobBncMJC4dSs0QSZkgKxV+oRdoqksIj
SRKqwBC3AR/BCRVaH5EG0mP0/t6PstM9dgnZpAiKl2uDRnHpYjrpuhDz8uM1Y8u6
ElZkDLl+zCijyp5kj4h6m1ij5yn01Rkyw4V0x67928Xp3pgqwSJdVB0aA3zB1+/+
pcTD/LUyj6DN7f25XD9GVZ0QVV5oLdEThhZ8zA1jvRFd6PCVJr/D4gr/0lAKpdj7
AJFtGYpZrZuLru8Rk5VJTTeixdCLqacsDEHx7WZJGeD5SblgNXUdn749RBvCtOaS
0wBlZjIEfmHd2gyCTZWyKN9VrpKRA5ErZCcSI6SemwqLfv3MWfsw2OaLIRTFJbAq
nPxw6Q+XtNf9Nppe/U6RtHTwKWXUzGRjcF1c8Y2L8aeamT+eb0N+42xLUKdvpZ/k
8JHhAdBriGtaT1tPRDUxcuPh85c5c54/6iELznh5izZ1l31t0J2t3cTzB9WUt4OO
vTwKJtBAlTut62v00T2QLRPl5IYnxL+t/mJD9rHRpDMaYb2il6ypm8eXJpOaaS6C
WHuVy0T2Afd5IFVpOpuVwtAlAqslJhs0myeI2EJMcJ1fciTeQoJebQxN0V6qPXhn
Wo04nz7h1OUTvkstn6I1RGkJWSu68PiSvQEirhDvkquU0FMWQW5Wj2bJni8zK1A/
XR5DwfL1WJuBTRJGI05BsuUzPfDxO7pMvM2gnqnzR0tyJnFGT0RD84AHNabW50Xr
kP8U1CwyfjUupB7xDt/FW4k/q3MhNOiSlc5Y/JZmiTiUlb/PWl/WEC3BZ/HXcmWX
9Zg08fRi/X/7eias+OBOWX3tjCKH/TMWRTKozM/RRQ5imgXvbzIC98rsTnANPT8i
ixDfMJwCNJ4EKzIcennqs6OseD8t1k0C4NIuwWFbDJRwS+GlS2jmo4dCM6sJXumX
ndvwYLmqcbExgl19ugSu3vZfXXd8PZLjz4BGNnZt6ta94D5C2pneTnUJipANCNQT
KJCQqvsyxWMMuotV4Kgf+Gqfz16WItgR4NBEktuQmX9gyIoYorsn+pBF5XeJW3oR
r0j/V9OkfU65QCDfMjY3xgqPZa3cOUc14R+gGDLMFDQm4qmzqAUsQ/A48uxHQn43
I+t/XiSwNv+5MH1cSBq1utMjZSDGF/5nK4wCsYDOPHPYc80UA13o7PIJ5hDCWPjD
xtdQktEFqgN+tEPptcSc/1j+smmb9ESapDhzAjnXhfycvrRO6JcZ3hidi3zbyy5t
fqXkGDzNLP3pTXSRurdISKaYhNMl1ijKqFD3juuSpCDK0SUgo0Hj7Gw2wD3IOkAf
AFyE0jGe8bc5Nnzka6uQzT5Ym5ghN9lwo9+VIKu9Dx0JNIl3AAHIW7PNaAuIhohd
bVatpLRqKKrPrPGUxP+6AMAhwKhxAPrXsK3yTGAFy8q4YqtAD+jquWAiB94Yau+l
t/zfDws4cH/j3UByfvSsNt0ZTJyID5+nw/kSc4VmotIM4pUYjE/hr8dkAiarat38
Cf07YyHUOJgU5rtyaVuA54w1CfWRDc5ddy7wjX8Vz+IfQOaqIZDeq0gRRCYLux+z
kDMKcczv50MQTIZCjhC2jIzauw+TsLbcmMuyJWoAK3ocvVIeFsaVgFMIvqKvKvnd
ltK6Pk7OYfizg78U3S3EsDCB4E3FW/6lhPwt9IiCXB2Si+QX1cp1pZB53/OR0hCY
tDA5n7UyBSyixfLndE05UAK1FzfPOGXzse2Va1djbbByGhqZDziq9EYveg25OyVL
GDG6UQewvj3ZzDb7NV21qV3fY3RTv+lD9GucxYDBIEKiZyLiz7tIXJ5DpaBsr6Vb
RHLhD8viDaUVmXL/O+P6MUqy8t77SqU9sGmhx74geAlBHdF0cs7W9piD+XzDvjM1
1cmHY2qpX+eNB0pbzdXSFiVzZHqsxLlxeSZ9ioevya3jgCjnDUoz2GKQbyqR8qZ3
6fRa2sCrlrnih4w6QrPctv0Z7JhTPUSdu3HimLRgYQDBb6O8qIT0xEYK741WHT48
M6BbX4TPSSCPIiRph+iJuHdrXOy5tWTTnScfIQ2I9430ZSI1dao2j3OzKdWUkBMd
6OANlBvq2OSiG1EkbU5hjz4ZxVMlbB+Xr5wj8NjNF4y0Qhjmzs9ih7RurH/bT1CZ
PbSn7Vqy85gV00l73zDbLNELaltA+xbzSkW5vxUDmnfl3J09AUtSZMpzTESwL1rW
dT4fYDEXs0WAHbqF6ZwA7zEpQ0ZN25M3OU6RF6MNOACcbN7LNrWoNEag+wt8obeI
aY5E4Jks43mVXZX9fOBan0hd8YQpXxjUO4V0P70+7ZGHNrLs5Tvug/BsiKj+4jfv
ES00mOI4kF8zREa2llz+YJ29qCQngFp3WDcNKqqNLH9n+n3UFqv5PfHDrlFnUTHC
2crpI1rtRbddtygvwxDQiu5bIWJeC3JAZNjVHWsq9cIRYlGQ1Wjo1UlTVE5yH8r9
9k0Uk0rgvDGmx+7HFsKNKZa85FGriYonkSgdyUvvIPgyd9YpbrurpSTZbk+/hkTh
G1jHpscT4CGYt3bPRG3A9jza3aX4WlU8awKRIF2jZ4kFonyNruO2UKnHq7H7xYgy
DkcPuk6AvjScoZdlXIJgwCXOoUXG2JnVf31rzfKZiumKsuZtdTDS7V1O1rnSpsF/
Wo9tDl9vqY1L+x5q2O930RNLJsah/LWujn88e1MoI/fk/TSP5oW8A8tUEfdDlKZY
dsYruJy2vJ1YE++HwFt8Uf9vY6EA+wj2Rfesv8ecN+zxtJVZtey/LBJzppZ1EJEl
ohTqeVVxg3Am+wGWD0ZUUWBEyNj/qpSv1bQ6fc+cWzJKDbD/QJLNSbs5Nbu8AODC
4DCire8mbs5iSXxOZOJcRH4T8nucI78Ic0v9j9YFSZCxU6QfQ3B2cUCa8+JkynYG
U9607oglg2MXoZJDcRty+AIfirATuz3cvUG0pKRO7RcZ8JDfv278WNoK5ZGvrekE
pQaCqOIBTW6erEpAsltazR3YmHEddERdnK/4KZy1CQpRh1F0BKqSO/XMZVt92xd0
kuS9kFPhhfYwlNXW8FV+Le0dMp8XvW73XtHtxioU9CIXaJKPLbB7451pUkUlX2FS
nNiOt2S0OODqEzfQoTONxtGd1LLputNDc6uszgnpJ8eOL+Cp27G9F526Vm5imCKR
gtyRdWGGhp+fGhPjkimTaJLrE0lwIdAFrWmTgrZ6xgBvjDTR9pfbTyBsOZDWOUwQ
amtjDOmk9DLCOY5GDvjF45SyNw8L8nbuGZT2pdLZJGm3ZEKYLdylZIPhdxekNPHN
Gb012KT3FeEWT0OqvGr8A2XXEhRXlJ9S8Q7eLrlvapqBa6V2NSBry3qmz2W2f3vV
CklNw5HUtptzo1wj1NqNN8i7ZigHVXx7GpxwBxlcEK5Wv5pGo92Bbo/A3H9VEk/K
t/YZhxw3pqB1a7L8sjW+rX9bwHsUZx2fM+z8x4vGK/Dy1yMWp+1BrtKx29NMfag0
GRrgyiqdlhg6o6B0t9I80Qbxp33PyWgmh6w4h95UFRW3tqUvMYLxNRYEuCov+eRN
FQXptRkgxX4wNnDrdqjJrUlORSpCfVv5qIjAXzGyBtqW5eJsjq1vB7HqrqNc8Zc/
41aPIKMRwL+k5KLKOHk9+DvsOlxbxHUAbNcZhQ2TADKNE+uti6UyIKtlkTC3BGmG
8679MZ77PqaA++U1Kmg5p3OG2ND5pakI98CUNp1f6NjwIeuBsmoo4btXZd6EMGU7
1AZr8JQtO7xJhtZKzas6EHj4+NlyCnZNiJVJlahlU4hzl1TMc0wJnFsqPPdFhlxu
QahPwRMzkaZjb+VTwx5n1lR5+zCcEwD3qKWju0HKJcs2eA9Iw0ACkqG7/fzX0XmQ
fbvZgdYvANrEOoMFPqNndYU6KH7ggi8Fgz6GDTVofSYi7Xq8z69euvZGzH7OCuna
4EqY9OjlUM32H5EFnXuQrEPuORkGZ62olBc5mq/zFQj09YUUEgLHhVszAcHjfEuD
NNq6h+EDKEkOG6mDPhk6Q4gNqQR7WlJdLeG6mcWQfzu+cc9MIrCLyHqTStSVG1xN
0IEFW/AVToDWtMhjXjpyNF5tfDjWzX0n7r0MhjIirNb5d21+1aQqRRYoojXIqO4g
qNU2+KaliJK+VauypkfeWU8KZ+U17KW1ocnXs/hcNut7YLb4DYQt0Ly643lmDp/M
sjnHeTuzm7kh+I4m+1QbQDgVxj3Gice/21lvsWNcdWSSv8uQzqxwBi4LY7hNQQ72
LWcW9++gvVcsWDm2/ZWEqCR0MKpadP+JG2QRaVjYCRI+9R/aGA+9Rq2m+YQsl2xM
tcGvDgS/HNibnHO7tSvAiL1RYX8XL+OVdqPy/xYXF6HW43fDIJMGLipGZgDfWfPK
cUD+Oxo3US6QiVQ4+lFevp2XMza84LG1taGnQkxz7v/hglmxMcaop9S2W8iRybwM
Ra9gVLbfaXmJGI6CVMgCWAJxW20AKitUNUZYI3w3Ln3Wx+skqFKom4HzUSwKiH1w
p/itaeZ8mhNhLyn0DecYdTMG33y0lhv9FDs5/kQQw6uyAloKf09YBXVAkpSj4NE0
RIAaaMRl8njv0hdwVRhnKGUZ+fbX1BLyJ+Cot/KghbqXgs8Vyv53emTRCbXpxHo1
VFucZ6yZDfcxyEfYYDASpcT7yIUb3xwLqZdTB8hf7P4645Tl3W6XHbL3EqZ1OrT0
Y7wJglXe/0nawhLgz+F4a0nRBGq7OZ7eAd52cGoJ6dmbR3YzzRivagWh3UwlHLSm
TTumyJQ97BtV1wrndhJHRG3M8SW4IahBWg2/FbJz6/5AUotVwg1i72Q9dlwe9mCy
ORsCa4tWeqeJiZWT3FCxinSNdqeRaAnzSjlijFnPk+21DJIwFh/wEViwUxJ+iSef
a7ZsU46GqDU/RX2xjo5j4AVjXjAkFningyrfvMsT/wcEhk9a6QuKyPVhMPt+ziRt
loZDKOsAzqfJgnnWPYDXjqoswUos33KJ8tSPQdcos/C2616sUtIf0VEJ/ipcQd0Q
GHE4eclJzhXsYq4/dWdwC0nyBy1qni+GEJ09Sqgv1URwWGbcTSZnxnGHLqmT0xpD
5s6bmtaiOJD83iOO8LoMMTX+ZaLFa2oux1Em+zhvpAGyYVbiyiOomjiYYFL1RBrp
emQlEUe8cr1Kwfpv27Qn4xsJyonhzebLcBn8Jftreo9QeE3fUvnIu8nNzqWl1ZG2
SKXoPQIgNKfWHVOnRNl+0NfKIM9oBohJn0ZsVPZzUg4xPdJSTMnamcGb/xCL2IBX
cvxbEgoOFSEGV26PSNp4fez+gZN27QwoCgtLl596Cd8EiiHFLqHP4Gam2xmc37Rn
onkq5iwY+X5JKi0HZ99p2zVaB6FOLYIeYXdgnjyqC3ahL4Rv+1BV0tqM7jP1gEL8
4ygHrrWUn1pdQ0bpmsVtD70a5p5XAIDtxZe7FXcmb20VkafZmMbodvnqA1XIZxUH
JHi+0Mjybh4ftRAS/Ce+5ybF6VQs+om3630rvJKajp7VSdMmc5ZpyoUM+wyX22cy
+41QXOo3FSu8ore41Z3U98k9BAqwdT9t9mXqPLUNxxoW0cM9Fqy1feFm6q39tGdx
iZztuKZ3BCtKAoUsJ6j8WZG4qzRv5bo3MF/CrPDY5TaaSFU+ZCtvx+vEP3YUeE0s
9tS5ylmNORvHzA0SvU9E1kiXl/Fym7kL5P6ed1Q0Ws+pZIDVs0qhLbNj+qcvJrAr
A7VUtRyFRM+BRgvhOTuJLuwMaQRnC8+d7aq+4txm3dUQpf9FRUYxs+AnvbOl7Tr3
fkn0KTv0jo/RU8IM4F0So/PzRPYgvqzNAK7+LsZDkcbtFhFM/IVCWBM/RiNlbHTg
U9hGwza6JgBQYxd5gLYFQTWnlXuvdElSW1nFbxlNoDXYMC8eZzzeUCQWDeAZ7pMK
XCBIJIq/Xylr/TUb9uarlG7fbWv03I8sA7/PMnAbnzb7/8ncKMmiZGAfPoyt34NO
cJbeCm5EqGZc+ZdPBeMxH70+T23gSB5V8IWB093CO9mjCTNYElc1yoisV1moCbGc
Anq0P9F7PrzetoIIr/po4OKRaaoFTA7TqmuVrFp8cCBWIkLXty3Xv/3Cc+QmSHDg
vIwb6BdbG1ud0PSVz7y4x9pS75r5OSjPFeb0Ionw2rqb7ZXggwCNFY5hbz8hboO4
LUNuk4xzspJOq163Vum0wLNviiv7fDSZ/fHWq5k+N16AvBOhbFnScQQ/vluYt11C
DDQu7N0h5AOkj/fAHwrHusyu1CKl98iAlNgJr4u4oefg/kiV74w9vvtpByMqOk/3
txtzec7e/yE5uForYu0SLBmlKwcPnUbhBFKjXhq1BTHnlmtHxUAldH8r7N+X8P/d
qwEldqBAyfnZdqq+7367r7Zcf9L6rx86gxLs/Bvttt7mVJjRehdaObJ3EvX26Cz+
1hUOO+2WWf56B/zqMqxahfnDMXJLY644yghEcLwgdH1AvoMmpsJJdkiRaqF0vhtO
kStrBTDhpFnlyIHqy1cnBvZ4eBGwJf+0wls121IIh21F1jSyqmHuh9pczilPlktE
rTMYiyTfE7cowzcrvutgZQrQOAWhXpAHjlHUICo6/BjCO3N3GNaS4bWAs1VdpwVU
kZCbBx/RM51g8A2fGEC/xepp6nSD6YAmCqcLdzOGpmmZOlWRFjuoCkVATbZntxVQ
zAZjhnvU7u3bUQ5Vwul95yhZUKYQ2lMnf6+RvolsmddMbhO4e2PS+pLbMArwAb/W
F9DhIUnbSerNw7BwNkd3WDI9Kijbh8RNOCt9Uhk08i3rAkEEBJsNtwZ4B0YPdEJS
uJX2GEBGaX/0A6UKy66+HrTYtY5XiiJMRjYN/71XaQfJAvjJECkV49lbkHADHtuT
C0v2eLrw5gKH4c82eHORqy2yZPtVTnUs8CbPiMHrB2omSxZCvEn8nrqNzqpnlQ7K
w2aqRfAePUV8pa5Shlgh8N6EZD0P0yL8+8n3no+2H46q4fft0UF3bjO0KMP//zSv
QUT5N7eF6pZwMYtRbYkza9NxIuIhZx48tgjczuijRQd+1KAfmEJoYffaU4koaCXE
en/3ts7L22rEYtzNP0eb6UxQBrbg1upeNvITff+CaRgvTYQnbr3m7L1mckQzT5pW
VLCOlXRTHVDWVLVtJdxUmyNbMzLNRjKq08zXCuT9tQue9UXLMi70S1b/2o5cf+Ud
aJsQdgshECGOczG9nreJECrPuVSvFhEjOQ/YqB/DHbXIKJcseqtei76h3+OzpSeT
oqSZVffQQy9tQCIjTB0T7mkAp9XuM+CgbRvNfLu1nDBgvuYHBu83+fHjyUezFAlZ
zG5dvghIUaxyh5ah45lrXOUqTuwjpPqyK/77uPLjfBUyXu8pPZu8JX8JmdWBNQq5
baL390dtkKotiBG/MldredmPECKXDCL8FVLkMBj+/9lEx6VDOZJ1JBzPVDyt7FMT
TyjtrqGdKmlHaeL19qmrxjykYVkc2Xi7T5x9bM58W2fWEM5k270crJEdqBvIcaHr
vyzex0XSq2ga1DvAqoUUqm2pK7Caww9FucOYb15GfqrATzmNN4GjSffjeQZgWRVy
9XNF2Ur9blQRRTVZHnpzGOF/6Vh4vxCd4CH4unIC6zjjE89L7Nqi6dk23qpujpfJ
1Jen4EPoAaueU9XEwMoYnG0hUS87B3lGP2OswtoUv5ul+PiU7jwP54ZMBjJcuh+T
yYyKhhqoXCdHUg7hyExjrOr0xA+uEXmOXc0RBjwWK3D2eQsy1vprUwmopXRUEBnO
ks/jhGBfg4ynUHW3gqct6WCEGJe/3QXAM25vp9TIwxDkPQzT8RKQ227cwB9X1JKg
0n4ogH6HAOHIWw9BnygyHDOsqScldRQly6wi1IgkTROR67+XJnC2YK8lyQh62hDS
9h7UwF5/klsDKLJzLW9AzaI4S2jcTatfn0TF8c9U688LjZ8pjA1IlprQG6cTqu3M
TebK0w3zKjN6+htk9xfPmiiD2dWufK07WxYic6oL8jeQyaxI+yoUJYypR2dWO9ZX
aHkCKnd7FVmiFzfazvsZ4eQZhIIGN5/QsLG0JPTk8eEOjpJI3pMtOUCxZPZvcIko
HudZoOIrcnnNCr4CBhTUx4e7oUlDkcgxAYw9C93o4Dff4aIx/7A00CFHFziiyUay
2RMm658snOSOLiZhpPF40E+jDyCqtd5ENlIPIAIoZcOQMceQHBhtIP+kPB2EVBVv
VFrurXngBu/dc2EATLvcWCBYXM7OOaCWOsVvJ13mHJCo6QKlW+Huw1EN6MRt5vIx
WhvIipFMeMw29bPO7qbNiJfwQYfWP4nVLqHjt15aKmUtMh0ZX36vg87a3qnp2M3e
tMvSUBKlui8YHYpQyX4RELFpC6Sk29E/ubiia6e31ZndwgFm2TPF79VB0oDHzmUn
eSQZpuGcaJ5w8inH7YcuUXTdk5DkEyyV8aI8r8fkCIATusPo6YsOL4F4+efXoO5D
x/4//6d6f65fyOhE0wjNlfWMEgfHgiXJxcAp1FxIEGlahVDZihVkB1SRh9sBEF9d
2ObmN38Yu4Shkhm41bKIQZCgplHLoPG+QUrqIqqQaAPzcv41V8nlsVFYvGglO3VV
UpqY6aQALw2bgGSgARX/ptUCj8CFT9t1amWLM5IHdmUDc9rJTMOm1qa03EV/C0Rk
Iivb3cLqVKWQD7kuC/VSQtDSMu16+6xeWE9Gjk941rFQk5qvRC+ci+vP6wPr61oZ
3DXFxzD0qpOB4EKvDgGcuoWfWDGKFWl6SHWVOuXcthF4xc7tJLjrD2/QhvWwVdQD
pF41jAQ5o6qlBFMSZ40ExnLmgzS5Xak29+uCQ7XYfSPW/7OyEUb7RHiXuTof6ApP
8RfZUh9uiTXn/OtoOXOUMxaBjGYWFQaWDjWTJGEaFiJcRxl8l22hYSeRm25cOnjD
q2eHh+a9sk4HmNs17cRtH+8KJD/2VlM4HEBTypRB/qdbrcDhgJk0BBZTNLydeKlv
9+He/htupEkf/W75vwDnmcYCHny0XTg9IvbAOZVWD7N+3dLedr5OZ+ZsKOGGCfnL
H0Lxl3gwUvruyR5cpul6Im1ptIKLZBQ2BCYGzizm80ct/uGJHXGzPr7JNgKd1n/4
HN4bkEfXHQMLUQtKuksu33HBkJHZjrDSikQdC0xUYsEfi38CFiBZcn590AyevCeO
Jn0y1MxVgDhj6dQ6h/T67pfufzVzrMlFcCV1Vysm1MR/KbPYedt9l/adjJoSb4cQ
LHjOK8XA/COYUaOIQqRH9Tu2jgF3A876m8JcINezUz37MItMZ0dnMSpgqmyYlz1L
ZUMmDsHm9F99zM5H+ST0YBnCR2aw2FZuzj/xn8RQ1YVxeBJXFfXmU7dzS06oASVV
orMnCRuAI/gEsX6313yhcf+TCVoHpnW2SBwd8ijc1/VPU/A4/QVYbESeF92fjJgK
b1KhZ2kYQxNTcl4NBqFjJvARgZch1Wmvhk/XRF7pEZvOJg7gT3FpyNHVcd6aqrYR
VlgAwReATEDEnpsofEwX25WkB/5t9rp7Yh1Kj6YXm8TTU7bUVh8nPWOISsMk7eW6
B0dsGj8S1V9cEGJPRNI/4rwB1+hSqWzgXd9WajL0I6dFUgC7YZDU8nEoRESz3NgV
lZH79BxGCDbKnabGQt5g58vAxoYrFiGHSpfcc+emB7ApPuLLRbI1eYhE2G27e1Qb
Y+M2xefxBlokbmsG17iw6SExLNyhrMCQTwwYvkRzE2z1oSY/ct0+Zl2AFM3RskiE
hCnY9slJrGhnH4zwX9jP+WF3a/WSV2FqPnTnFm4Hp6l0IPvLAbsK9OCbFSjM516z
B56P1UR6avNEH2FuqZrbvxcF0DWkF1zK+scLdfWzpT8fiAL22/Fy/2BQipWv+nlD
E9KToYjIVajPO4mLUQuxv/etidzKkCEr5K+DOvYOZqs49h/8YwBOOzxQEdrkeqpp
BnDJJBkDvriW6d0zfvRs8DcwcIuEdzqr1GgHPWcm4WtO0fzz3V2w4y6auhKNHr/+
FAc9Z9LIVRy9tS1e8o8hw5neVVBeeUG5SwWFQQ2tnDZrZzJI3o5SbDZoB+PfJIAa
o7R78WZ5qiepI62vOCSgxZJG39oLnyBP9SWL653Y87Bu6fh3C5Md2qixvvmJmNKP
aEcgrmm98fgX8zYsr6uMwcZjVTihcFMqLHrh+1mrnmHZMSlcZatTgad5e5+mZU6Y
RdU5ktL4lN5UNj0xIMBV/caQW0BMLqOECo5eNYQM4tUhqnUtM7XQyG6JZ1BWo5W5
yJDJ1vlwukyQLmwsi6Fd13C6PW1It4XlrViciRsMAqQ4Gs22IDCNSDgzbFs3/BUZ
5mCN3bxpiOJUU80EXa8+eEJxAHjeqq/4+OZEECmqDiQHh4nTWmNl7ZhLeiEfrxQo
2mAD8eKFvMEUehMtHdDJsR5ToEo0uCmHUJaTknRLWm1f1PBoFCAQUb0wj+iqTfaT
g/uXe5EsjWD7xj3HgpRjeSf45mwCIz/lkddcsaWXff5AuuNNIpUh8Fz/aE54397p
E45XMXysEQYp/xrPwo110qgJrr6JiGi/HSE4qs3sYJgx6ITqZ0jH5xh0CShTLtur
8KDqey9m9zvmX+vWjDWpdVUD4hbk6XDQEnNvky0YKTxcvTwrSvj7bjtmIt4vU4XU
M7rp+3y5/G5P8dnWJz8+trcRck2nBtdDbesGOiojdIJYNxjwYMPaRjJp9TQu5Tdp
+zMrfbCaNmpUW+c91908XyBBkydz935Eh4SyOvkAdBmoVaAMrRzstxFlI852gyyt
/XioeREp6757SRk90gTWojLNJYv/jKxvujcud6WDBykLejQC4EVXR1c01Wi3DrMm
WsoWd4EI4j7zdUqdRy1hEEZhQd/qRQyp8sT7SfuDMr1RnV95TV1V9ExczyWvdD35
KIFzsgiFSfeypkh2/uFCoh/u9afYN5E1DYW3QqSd5jh9mR0nnEHS+8rt90r19EDm
vZCLvfEUhrrNkw4UHqnTI0NBVZ8zAlvYXP5p9nyDVj34D/Ag6oJhjFjTN/Lo7NDr
+WZhzSRB+5w+vCAV6SQhrcst5HwcvsUXwRnn2ft3zNu+8dCeV76hmLgA0pISyukr
seT7WkI7gu3WTJ6Go8k3V1OwleADxoYgKfU70/3C0jK2DH04ziuMYC97qRrigKrf
mGwkTvInvtziMMKM1x76mQ7C+xWv4n9gW+fda6GsX9vV4nEM1K8pD+s2BBfXwJvc
M3Ikccdpc5o0W9OHBNrASkqyvvM/Ho5yhWdqgKUEEFQAnZN3LjBBR8kcAO/35M7q
Z2GgNm00nLNCyCH6myBB7XRMbSgy0K7LCdYWjYqG3wx+U5hGkT2jcDsXi8XGe1wV
OUdF9GGF3M9obANTM8GuB+z2PuwTLhWafb62V9K2lENv93m7FkDqM8E79/99b24B
PfVSUNHPqcj460k+mK+Dzw37yby9TMdiokw0LfLi17uzgtIs+fKpewd/F9dDnY8X
459dMdFL2KbD/4rsGmuSJhBL1wnMdTgwlD/qxVQLidbSbUIomezn8RkXqxKRJn+K
bBz6QqcExTb1Jm2nW+aZ0/+u6ACRaR6sDjnWTL8SycTo0a5T+P3HyhDzAE7ntvYm
JkyIp5TgEuAeDrppWrjVOetQjEOXkTp5/XqigLiv1Stiswhu8z/gHO23wlesAWxM
P+6ZE0iYWYP2LbJ0H1c6jhAYJKDzO9dcu8RoZmcuAGmwFT6QRtGqfjUqphX04O7v
UmoTSvv+ASX6yvRWV6S0m2WmYJM5mbOlNHSWpGV8p9ODN4sMcEjZfVpPY8OLxEPR
zaX6hRNhhPVzYrrStia+apthen/u7Yk33X8RYpOuhH872qS+sPulOW53Mh1ORFWc
wY1qzRdO9ZrQOEsnDnB87NylT6IQYabaMAc1qjqd3j1spQXhN7uSfBvh7lyC15RA
+k4pNqPDdpFD2EKdgb/UMW9ghuTsmE+7/Ejr7zPSdnuFujwhlo9QqFPc/YioSRGP
6xJJO2jyQT7aII5PNObiWr5/2wkn23IsKJ7FFuXFr6O/xDX3hkhDMm5UKMG/315z
WIUszA+ciVM6c7rgqBlsy0dpA6z/KOElb58nYwqL2d/SQ0O7GibLb+ix8MqtIZbH
dUyldzPNElzV/17NZqXc5w7qlOkMtrHdvZjl3LxXclUsgIaOzoARvh+N0RThVZWm
jtqE/zcp9fz5hd+X9YzU8zl357ZcwP5e7D9gR2PKSKsjRxuQ1o00TsA0PwkjnevZ
0Ls9LVmEz766FxuKwNMMlnNu1OC2P8E4QZ9Z/ZZTl+BBLcV+neZtJT/R1Oxcpo3w
UMpPbZZ89p7MgV+ENq8PJpKQWB1aGDMdQt5bY1hteeuFmwwuhr7gLoUKoZ/C/Y2t
OTuKd+e/HOzsrhS5JOccb5yUN/lzov+guprSd8RqdJN87N4u/21ATUNwytK1UjeG
fX2uFfMWzJ2zCPLnGWNsaYl0aREN89kc6mOluQTkohtz5IhLCidfZeYkf48z2VzH
0HNpAC6SCuCVNkRQb3FQ2PI1GO27cAfBqPCJkORV86EyMnZCYATYHDRrWBW/ZvjJ
LxWd5JIYOjLkRgzu2t0VyVi1AZzbCPAhJ0CmzQdbwaJv7PAj7I7jioEDPq0QApdZ
HHPey0+Yqsivu2lU+rfyRPWVw8bsxwM9Ww6m29bXL2Fvb9uic+8hxYnNwDzYWyKG
xYxdV1s6bnMqM01eeLXwiVDr0qSdbAoFhhsDvjgULxfiVnMM6GZY4ypuGFViJXpn
bo34VDzSDgXFp/QG1dKZAhonKdjQi+GVvQuFWK7At0fN/5xepldKXKpp1ww0kzXQ
ci3ZBukUXBX0dxd3fQd7Sl0/wPxKzNDVphIHTrdECJfRgWxRXRy3xuw/pWddLQeC
XsKwUfrx8UPHxQjNs4PLopf5z7Irn+Td1TEobDs/6ASVvAH3Rx9PcULNfQdLwUbG
xaK4qw6GvUrfJiW7eNJGgX8p4mHiEb+RUCi6mbMzoflxCYErIGtE51KLMovFpQqU
K1jcmBuxQYdS/SzVWcez4Zg6EOOYSgBU5NXqM53iNfHfoYZt53Umg367UtI1yqDF
Oj1TbFVev4jco9bnywdZx5Huc4YMV5tBmQDuhr6acj50oaryvYuE66xj/0WlKXU/
RHN3KTBKqFPtSZylojWaH+TWQZj8VhEVZAjRHStsndLZe7zO1+z/xgf4FGv1oYhO
ZyD83U5mQ2J9RCvAOaDgY+50Q6/qJ+IKA4Kk5Iy2zuQ3TtcwvWhJBaGOazZ8E0VT
+wTqPuhuspLTiQUnzwlNOocZ4g2MLi9i069D5Xdtt0zLcKZ7Exd1PWWI0LVobZ1y
4IH1GL7gDd7L8zX+iObBvz5Bhfk1bdBHWyGGH+3+dJCqy5opUwnZJQO9QfXvAbtj
h3p4nhATkoa5j4pXWrz/4+72QwmjQpLj6w7ej49ALXNjGX3srRPg2SYt7XQJkU9k
xqvFIJeKZM6VVeVlzrITg6gTLzOMQul5u0XGT6LSBCr68rCZmv/kVQOJcqJ3oV0V
kaORJPBh9exsr86JFJZdlESSPWN1td9Z7w9Z4ElvRK1L0DOXznq/i9fi23EAEQ5X
l4cHiyDlDfbmRXMZcrv+areuOxdQRj0NtDG/OHyjKh7fpme3lwlZxPfr9xUpzm5o
m5+JtgM0Gg7dz1PCeGlIdZ+H5fmiVTRYHTwxBiA6fJxAl0AOi4/igf2bEqzvSaxa
Zlyvxm+uVNJPz/pUbb+6PQa/epio3yKI71NMQqZ7lxHXWjWwsCre+uiW6Qru15+z
4pm8NtemUsNGclb+o2Krj9XEndodq4qVjH+njszYzdaBtBVg7xYbDHUutXMB4BEM
wB1KqVsBfBNJwEWiFhpl99F/qmUu6Rp+9R8bvqX7Btkf/ewndYYeMus/1+IRi28C
wN2EAPKmelZ6AHLxXOW6Ku5YDXwNbnA9kFg+EGe8Qi2QrA7SeVKDeVLh24FK3uoA
drm5Y8xyN3o55FRatDUJzDa+wjQ8z2Pkk/TznNJWPRal0jbSbxsXslQghfHY/uFR
OtHFBxXchzkcKmISiyxn/6y549sS+dh7qAmyylfTFYU6uPWjU51xeobsXpUhtB+n
uEEY1gjDg8Jazl47Jzm8gNKEq9I2yLQX9CIEaG27VuUV9uB+47HXfaUVeRnosrtz
T/myc1p8wxpsrUtJZurxHRiPf8f3KtckJlkNNHiVxF3XWSmQuiwpgMo5L2svaMRx
qzbS9H2RqT2RLx6S3aD10oVctarigiZ25yjArKsoJrRowOGkPCEXrgBy1oEk6/vu
jtKMOY0jbZ/5bunxaWkxLso2HKL9CfrQJ5IhOc/hXUXW3RY9ngf7muXSs6pRvmSo
uiSghsa7bx8N/Xd7xYmmphM+wxUQ5Mmv8F3NtBEVT6Dby0ew6FGZrhZZwvP9c8lc
3MFOoPJjLux6Ujij4XJk70a5eHadzBAOuQdax/6fdBmhqJ3q1A42MTRAAkSCnf2C
OXINQUgnP3gb34x1EqanAoslENbFy901OfMEa1J9117SO+9++jszc/uSMgmfHjDF
F/WHjZLRfS5ttuq9Q7Xgb9Ucgi65bi7ZLGHLuQjMLvpKFAbYp0bm7zmcGw6Dt7C2
LXilB1xUQODv4nptq5ANNu+Ss9gU378vACLMruESbg+PHz0R/+Pjj1koSHhF9k3m
9ZhsUoRemeqRZaRxshhUJUwI2BE8eqBpooV6PUpm+zy95C/bilmnAK8sEMoXI7vz
ueifZNvwHnFF7JcpJqMN1PPTWp+pFZzkPhGaAW3uzin4kwd47dSambPjGkpyMirD
ooyNH2wuF0pHo9T8mThThFN3o3DAQ8X2ySPtrRJT5dFIpuYHx8mtBugDAxqekrxq
Kw3d5ia1asnaiMX1vCSi1MxEcCV8cteGrg/eRinA2jAR73YUWOsAz2ffCQfss1BP
RBHjFIGWolsta7mEQGmHVhMTCn5mVwMoxWNrRqzgQ9+8bWRP7ZENO3mrPg2BDPAa
1PjswjrStbSMh+r7/ze6U3OYCw/rEIYZohLvERysvLfTvSajPF0MtiIujl8tlZuF
v9Zlrv8ej3j8AM05/6W0vtF47Sx2TAE6ZQ4qmSCV/hMxz1Rf9kTkFvCE7K/alt3b
HSn3UoCgvdDSyhh65aHLYtYKC2w941gbnOU72yV6Fn2ylAAg0Dt/WNqY45tHusze
YC2kP6RRPRgtL6E7tcoq1wzsx1ekFcA8U/TYIpLRoJk1UjkRd04wAL0qFtnp1z9O
iCpxW47Gfku4YI3jLLnLW+mw9Yz4b7CV9tS442DwbgwYvTtuG6LDZpVB8ZxlxOJh
8yYPuA4yuNnm/L9+1LqrD+zNDGC/FDBkRPFuhGURXguIyxB6ru9a7FFnV7N6mTBu
xfty5ZceuXzIS284tk/W1XA7bEVrgG1cnPJvXLea0YvzHyIcSwOXjJRYR4m/1xD2
Bln3kVRoKFCUuG8fgaMz3KBSERvns3RrMGq98b7DtptZTzg54yF5H0wcRkOLpeL+
2D9RfU0PM1Cqiv6sFyHt6HraPai8z7FUkBBS4a7zi1BO9nYnHUpXyFaOBX2LyE5l
jxnvj0+oDe4LwW3s774pAFM1GUINKuzkG+LdFCEZi3XU4oCOqRWLA+l/tTiWYXhg
gwV/VrLyGYcfiYuQ8hjw3Vuw4P8Nr5WiG8W2JhhtRpB2nUNGrUhRU4UOMCc3u+Wl
OpvI7PX4j71LpSKzJXDOFMaCOTETM/Lh14cgC36ZCcYWcBoCwKUnSaq43UU3AVwk
361FbDdTCfrC17e5llMgsVS353l/+cf6l26mB8HflYP6fW9oGjhM9opAhepwPPMB
Y1DUCMvmZ19qoCZUAn6AohgMUrqeKp6KdBQeYYmd2EkOV8FJplcY3JajkYXJkwkf
hMT/T7rbeJhr2AetGnIgxJ5tMrBcZht39aPrIROHF8IJ+gFokmZV2VTfvuSNOWhc
rv/zSv7p82cSM3MeizvN4Ilei7I8PqMFvcPJ7B2qt3UDnOxiKciJI5awUg9A4Uus
5m+cCA4eS+96qpGjl3BvhLbTJU/cLqi2hpCEhrIwWQ4fpHNOsHa/pL2MMVrWFmAe
uPoPBrB+efH+sl5Q1aHVG8eabkbK929UGoMtyaFFF7UdnsrzKfnttnOOMRRmnz5b
PPge3y5mCdi0LFgBse0U/G7yavG+KA3rvO68imO7JcwkLaoLQeDuqYRFHhxgChZ+
j67G1vgIuPx215SjkLAW2fClqcLKFlqfECUXv2YxzelYilhPIrqYmYEqe1dtcYDv
ElBHYuqQHRx1TjAPpFXt+IOpzTcD1EtjRc/RfJNGU7Wh6HL3Ndkpe+yb1FcXB0lk
Mz4b+X/LQO61vbLjcqxOLQMIvRS2JD1PjVYVvw1FBP26HwUB+5A8ut8Z7Qoone20
wZ6zEihE0vaY95zTvsAYlNjB5l04uH5357ElkAuJgWInmHdTznVmdox3kyJlC4Xy
/q9gKNDbH9gQROfMDUenGiY0cUfU+WXcvHrc7eoPN7yGkubKvSk+BIkHTqcUTfFB
VTb9zzicNsjoGWRcvjn1wKycfsy2oJuZ8bM/IbMw7lkCqNslYA8HgH04pLG/wtG0
PBS+7v2YuscD/6qSdMpGrbG0zE45Myg1AMGGMZ88hqz46tJnSocv4N2ILCgML6lf
bzBqpBy8a9aTRlsxdoF4bxLR9rzs1i3Vr0IG8/jVicS4PT7oZuUOTUZ1T76YVzkA
EAch1gMYQ93IgbUuamwDb9egV/QLRVIoh9oKbxrChuCw7BIfMI8US2waIoECOcmm
K2j29sLoKNFvm4oUsDbBFP2CPq4yBOsecUIv7kdmLC51cgFOc1KAEJRUATSkgqXt
MrVH5RZoVh0WtEXWbfQcd8qJgjQp/3g0m4ctH1AFAfIhWKx7+kFFxg5pZHU2KoeQ
qjJ0br+VGtQ2LxVP71jKPQeju7wvw2bby1RwvGPVdRUO070v63CGMFsErTFApFI5
ASEM8ld2uVstaYnFtWpQtEYRhv+BMxs2KqjuA4Z3+rVfKPTUBj3F+f4kk8K5nzr9
VmGE5yVTA0OmXwkM1qpbd+q5/afUkw6bYZd1QaQ83HzOEZ3sxSGLpqBGQs1nGoPh
RBZ7BEdhgR24tCHC5tSpNbaW7vc0vw8Dm/8BI+w7dVppq3e83BuRAvicPyrjZ32j
iKkWYdk32ofpg2zwXbYEAZCyPuwg20+JWHukJ/RbpOIMWvrEwlkP2EG3jVLlH+3J
8B1x1y/VxDU6MqhWX1a1xAIP9F+f1x9/MkRAgQ1t7il6GaqqKjbxSmxX7t5n6uHf
kIlTjyx0uwS8rT8RSxtYwGZf6YEsomo1KAA483pyTtk918Ujtsse3Qq6HK20q0ej
FtoS0u6Ksz0SCUb3C6UZOViAeTOeOexAkDH+JbwNzODxWCiSsa81h0kuMvXH6bCr
DCP3S8cKE6yWKZ1Ut0StpeBgSydCe/hcTrzlxQSUFLD60+YGBBxC4RK+IxzSrEh9
eaOXaVwWRq3WzXi+0qKpFt9lwOZFR7ZbC5xDZgw7xwl0A2hyGaDkSyEw7vTNv2UF
UXj5ju+avA7CH8OEpMDcDVMs97KlhDDG3DR5sEX9RNAvDkH9NwVeiMISgcAHftNR
kmx16xnpGTCA87+yJ94w5eczN1ANM2I7Yk1LneYSiKA64psaeY6wsrKp/SpMvTT9
tc0QICrqyWJZa5VQ4rkhoH6iBYOUflZXrH7ceeoucphnN3lryFVj5wRrV6S+rs58
JdQxXBT6NTYONNkNHm13vwUXq+Ca4vjxRTEA5ajZku5LStMFkdBVUa4jSzSV7oQW
8HpZFKkhxmj0uz8Td0aDWN9Wq9bB7XGnFnk0BsJw5dz1jj3AUUvG8cJrs3UsBttG
9zP2NGoIvYg9dl+ZNpriqVYsxia9xFW0g73ihn3X5O3d2RDYSs/hhtpjdZNsazZd
cQXb6oSvIbfee8hUlK/ETaXv3jdDyeLcKa3iQFHexOj9t5qHCbwX1i0YdOCKgyh4
CKJ5dvCNC+uA2k5D9R51PeuZt4tmg/qMXP9pOaRI+W1IihrwCQmos3GuFcrIVVQZ
Cz6WdQMB7o3AIh4QNbb2VC6osmNzl31pHr2bLFKQiC5T+yXIGyfmLGfWcC+K0VRU
lJYWNYQOBzi3vpLrYYOfiR9zlwvM4TNdpFoOPaCOk2meGvXR3Bzc6tN0lrHGIGmh
sPFS5bxS4k+MKBjIirS3UffL67QEBIK3M3KdZfkTgnie9qUcM6OUa2CAXWqFXDIW
LbOH1ZROwMtkxUC5EboGCRcpUbZZoYFMGLtv8U7qtDaKuiHX2wRAV96gET3xWwDB
GRK9DmzuIlXOaHuC7xAgmWnlKkhIB5Nv0YmK/YtGuwJ7wXQRLBkRzgmA0ziWltOy
UBoKiP4fBr0K0DA0JGkhL2NVqHqXTzS0PCaea4wm0Wg720+mJhGeCirKTxm3UmiO
bRjANdTJHvrgS+BuaVsA5L+VHdA0jVehogfU01lDJDp99Y6fsszxtAg8nN45Od3p
0fMi6yimyKLbZj8TSrXfznfKdkSQZH2y/iWvsYotEdZNRjuU+ArUjnCn8L6n4xNz
k/mbx5PlvznIZt8VYNQ7UP/mfVpdCkOUeS/DNd8iKKJ9jd1Ea8Yr90oADS4dZhTb
/sRDTwO+G9InCGIFVw4hUHPZOrvy8oHbNauHjxr43XHi9n0Bm+k5XDp4VSM2Qok8
BmPSge96HYFBUcBKRpSB6V0+N1qJEa7A5c8unO37QHW/3eyZadhOaLoo3pE62Uvv
pAxcnCrSuBQpvzIV2cN3Nq12bacP8sQ6XmBwT9IJqo4/nLZh4o+PqpN7jchuj4d7
ODNNbbl3nx7vhzQYVd6OPbD5AlbTwiasxmtuv4fjnvpvOtHjGW0D2W2WMxp/A0fd
mFzbeH/uUhWSxfgISmww4irtj6OGvtZZPWiT/W17Obg9X9dCtklSh0O50JxsZxxd
/85dWxZGTmVLyao7pCNl5ySV6VANFHvRnGZ26jU9cb5bhnOYXyTSB/t0UXG1G5jw
TbWxiTixtQUMK3pr1uk9KEtWrFr/MrCJfuFqF5YC+DLtqibO6DfJpYiaS2bFYfBH
vK1d0FkLOItVOO3A3qLDKSnn0JFZneqCEV7udiAkPIG6gGrloCocLiLciOjDC8Wf
te3ZqG7XCn3cmoW+Sn+jHlB10AvlT49nuvmujRgKPSOUhrL2rqxV2pm8xkuUFEFY
UX3GSf5mxJF//c2okT+LeA3DQzKwAcdAG7QqApWab1yaDNG51TwGoNAV5aVvLvLc
jIT6Cuetxk3z90j4L6UJ3Le/ju9GNy67w3ksKzt345EUjSPm+IjoPzsYZKOqgz4h
okxfY4sJNkH8XUQjr/CRDBiQ5f2LpGbklVKWht02ooSQpnM6EGVXApwEFjH/ZtLa
1cYk6JxkUT8vRL1XvSfKzbA6JD0gQJro4jF8xWOoCkQ9CjKnrOhdCvzZM2ih5vr6
1tMGooekyp8MlbHNeRQq4TKsHXvNezFNajAZNclliiPf7RjH6V4DDzyLjZfI7L3w
BtMsJMJMXrM1aPC9vtzsF2N+YfY6x+eQdpoVklYpnnjqo1JuT0HGc03EOieG2rbw
PiAzgK+7nJqOKgxBqHfkFI7JoYW67w9zqEGluh7aiPa2em0pnURnyLFkIzWLdOKt
0X3nB9cgM2ZKo+se7Fp5P0owabbzVhXESk/DnErKA9Fqtt0685duqiodeyGrXY6J
aeBzLqpQyuY4cUy6JO8klEI+J4xj5hFEOzGUbp2N9RamZl9HFhIm+fbvcq6yTf0N
APyC0+r3ICaFSB0lETsHLqGLTdvRiIqy6nZtoeH3wU+oT4IHJYCHuanArBUO4GAW
I5zsQDwD7TEk3Xlq84yhSM+t/zXivvuPJtNRKhiPXpGsq2WRdSEFIp9wZ3eZZaSX
15bnqEqvq/YefglFLQSJOSdez67C7LJ/XVsbhbrpC3dXSGissACkVMlYHJUmqYVX
mKTxAz9wGsslmd7hZok6GsFI1zUbNvd+QqZifAzHxXMFGCvn6EHDQC7+5jPh7GnQ
he2i513K/z4bQkRXParI0aouqSAUlkN2UjzoYTw9N7bbRe9TOkOPLX9WR03oPOSj
g4ajNb0nYFTeDNYnZEpiIkVYam2kFBXyHfF9qqpfsvOrYKGMr1NU3tIQfwNDLCP3
C30L9F7xJEP7pKuk59coysiq80caks/+Mb+fkc7j/+iB1b2MKpDcKdpiziS3Q2ai
FXriR3WolpKRBqyITyY29dL+yQTUq9zgJFTbUrmAkDdND3icyz7XQ8SycyzPpc6A
8gxAH4ztsjkJldfF11PtVhITAUE6jgBnGdCklD3j+E59FAFzFG/LZ83XWCNSzIMv
PlWwWmshBbqi4s9BJpF6Yuqs05xsLGoUEQ9zRZAibD8VQakbpb/ipx3F4B1WAx3l
1rPNJJTUCAPqeG1mZNuAAGbFs62XAxuKHfeiY0wbqwAY114zXD9Z5Eizy4AI2z5A
cywTiufyYNsrtua0xS6leYeVh+NkH3AqscVL3KGViS87tXcjwbrtp8s+NKGR2smG
XQS+NuhySf6LqdvSygh7Nwvlp8tdm3Um2ALElm4gFunDmjO/f3KC7BAPv9YowjuU
59hJUFUYtrb/uObCHT0lTAUiwikqo2MRPvUo1dne+x4X2MhBtVuO59MfK3SBN5mC
Q6acbhR08PhR/LXB85YNP2qHcCnnwMdULd5tN2QvK35gVGfqLISO/vUrLIygkkuv
PsMilLTi9ijUQzcC3nuBmV6G/X6MOjAlJvHm7mdxXv1LuWR5uVaGSW6U60xkRSaH
1N79bbmc90RiRkLwl/jg9ZrNbJ/pYVZJx2fUzErkNhtMesd/PBHQPOyGzpUhsnxo
Kkgc93RMoEJSCfoa0dWxWPLcYaUv73k0rvzhg6YLavqptiHjgsercclhriMIrol1
WxIuLTJxKuGrEjzXs4H4uSnbje0um0RyUj6Mk5ovlz9df9lZmDLO3oh6jCoSHA3L
YtDjOWLGeQiQfYd6GKpO/xUGC9S84w8M0m6uQQO6wcWZCGP7zjR2LVsuojSLjmHN
DsrOfZP53qveM1e0rhGbrHGOgyFIPvzYL4C461O6UquseXZzQoI5bV6C1YQt2DNB
C/QE2bMUNtNVVz3UdgCoWATHerXkxKkHF33Xd+Re5VyBKSDi+SHksBh8Yxb48a0z
w4KnGceNIlWK5Z84iL4KpcSbktYz5km+IT9DrBTh1lyFOLKEtTzxj6VC6Z4Blnsb
vsTeRk5ZqDfe1FM5kR4G0zu86yTTw32Db47g9tBHsYC+ekgBlhDa/oQ7MhF6J8Df
bDRbtpM5+0gxLJ21CIFPaqW91o0yeepFc7L4WFP0v0d9uprI5YKqpWKHaLskaRv0
8/eOwjuw/REdQkA3kyEcrrqH55HwIck2dazj69dN2sshRfZfs9uGzGb2aLAee6Pp
7JnVZKYXLVHf1fRHLRhUis6n4EnX7CbEDnsMDBMKGcR3KqUNeXbI9faf6nj5eBeu
VRiz2ngHfCYyKh3ufdkxzbQVFMtbM245ZIHJAWu84TlS6FRoK4ueSp9FYYFnVYL+
ZBqCv8jDeu0QhTlD7L+w4mqT4v3d1HvH3YlDNOxqUln4TWO5hIXhn7qAiCwC9U3g
U9dEgKFtY6yO9cBjQQVs+IMoaxWmLbeM0Qokkl5MYlXWT7TELl/A4WCTMIGMFdv3
qCRxEkDMBpm4s9Q7imSE457E2QFhyQRul7dskLIZVeSnRGWexk0O4mxZ+PqgeDha
MGWxYm3goMzymXdGGPDGwc+dweSa1fSq4RF3lv8XvY74fp8soX62x30HmZ+MUzwX
H3qSqDQ13XN2ki8UpF61WWGcaKw5Zb7kUWAZ0hbKVJRL06gAykRWupuqILzXf9Oq
64siiIJdtg7a0YLVDlpFlbK4veu5ZpY4hjkWtuQ8I15kyj5sa0Wno7mnkh1qevnD
QT+ng3Hned3nsW+GYvh2zDgN4BLmTubqFeMJQv02rX3+lbIeQmuDIa4NQWXUSKf4
rv/EzW4yVk22Lxu9yiXJfZlr7l1vmfK9id4h2DOdqPveCcWyNbdQIYUQIlK4HTLs
I6pLM/QXsAmsMekEHnih7dXhby5du/p7pXEnYVg6jfZCKPPvWPKnlYG6Wj/F3miJ
HtzAyvmBAY5U4XCfyk/p+leP7JsAU4yQ0F+qCCbiOgIyxgg8khxv6eCtGoZ2/r7t
M6CyHB5eSKAEikladMx879YfD779Rujlr5yMMVXumNhXjBXq+SsikKbsKzA1Sbjk
YIAY+KDahi7zc9Jt0TdmAMMH9a7x9wnjc6UTarAdv7i3kWbBIt9jsQzctPFQWRqP
koCc67BNmXLQR4eUK+F9UFsZsctekWT3olaZP8ViYLUAL5MSNCTvRFWjKQDPk5lV
ctzWqzKDSGuKjMgHLMnWqsttBdFc79rLhI1T+0YbIYlVMHaPjKTsJXIYjVZwW/bW
tltNSphfeTdbohwWQFnBwJnMvfqHDnp4oXsPdnkZupa9My2IsXP3OJYXECiKug/u
S0PgvXsP+wnIvyu2b9SjhgntrZHh+F0ouBAjMLdsrXBoaKmacv/VREfiLTcd+eIU
bXVvgKJSWYwNMwIpSo5ZPGaXeB05CDTuQhsWKF6Mf+rKwBK8iccXtNHCuT5kH3aD
7Zj95z2FIu4jjtLzaenw9b1obcJMNDvO0cIvMJByiQdbtDUzrB52V75eXCxySzKM
pGI5UOdfYa9yybrg4puzmxDP4G0HQ2M8A73xoX/3h19aKvLxySxUu6ffuYQtyFIr
8vQ8avAWBM7NafQkiSrtNTUJQgn13XxqLkHLTjNiQm4AzJSw9MYiYXQw4h4ud4XL
v/d2d3CvNwLjxSFLcqRvIm3rAdv29xz4qciqM0bDZ/InkMe0L9vo2OkbtK9mbu2N
bQarerCoLyuww7vaXslrlQ8jeJ6r2P0kZtn+unlWaF7SvhYrDs+EeQStdfWmV4/3
XdImg54joOrj7WectHQskt2nklCbQjLmowTANyWSoOC5MJ5Xs/FBJSfEkPSUjUhg
pyf77HQTulO2o+YuiIiYhSSOdddI0SF4DytQ3oN4vBIMyxa9x02fJqsXPLxeGUOn
3Hg7woaAeit6DWsyC8VD48auMVS+PoVn4TWpuGX8lqOAnqWm2d7J16zQ2UcPaWEE
OAk4pj+LVyo26QMNPdplNCieU/dCH9qDSsKRr3W3EHyDjPXP+nLgm+bBRUzxqWLR
ZNSEsh9W8ee9rd6jL64miLBHrkj3ACupEo/ZEa4zPwHEthpooXbyxb5WaFLCoS43
TNjxZhXu4ZgCVlc2ewi8GxDTLZHiJfVb3+0NYwc5JOqH8xNp8Hkszpy/X7/tHTy5
k5uJ4YOQg7zn4yup369s5IhCDmBxTu5OV0f3M2Q7rDqem4vxzIJLLPaj7NRcKFGT
L3QChw9kFdwALlDLpr4WpPX2wm+jPANYJANEvZVWYsTLYXKjNGpGtoZx84SyPktL
hC8OhxlCFhT1htU+tGt9/E/LCC94Vwhk89pM6cUrbN9fsi30FJUHzOe7iuSabY7J
0u6RnFWNnJM0FsYCkHzryYUYJKugEEQUq2IvS+d0PTDigFi+VYnyIi93Kvvse6/Y
ddWdU4OwCXPiru+NEU5CHCLqcjROeA4b3mWHxMZDYv1nLax2Mp4/BJq/8owgGf9R
k412WQkNQv3BZm0pFqpAN4Lxew/3kV+Bl6al27yiJDUREJ7hE6J72fBnOwz4UL9Q
yowaFh3UpeDKdBPsw/5WHOmgtQjpQxZ9yezRvay5+MRNGHpuWOi3NZjb8wXKtmYS
SaC5ekZ0Vhjs4+RniwJ1rWA1JQu+czyhS8MZiDbemGEg+UEfJm5bofEjX6PpdJNz
+xzWfjkxdekxDEfgomjwifi8A79MlYynyg2frKf4UZhEdjucW1ubrGHoThH0HnG3
ckXnZDCvceFWC0D35di/ZUy1XTUqtg1m9KkT+ct3xNbWYn6NCrJl8dRwelDnOa12
/DgWPxzssPzjj1KU+UkpE21NhKRwWVG9tyQsDg/NZAiRMoqnm3YtUcdlfss8hT5e
Ojy+gfswVfM3mboXzDFW8RH7recWmiB+SZAV02fpIGwqvYKpPdpvEXBh/5BMRp+R
RCEQBZE2qjoBKrMOApm/KHQeSukAELGWpZ9lwo1hK9mX+3JDSuH/dSPE6kdsMYdv
iF5jZ+vdQxqUgUfKpJ1CFXljBX3kKuKp5rpSVceP4YmnLELCOyCa2nG7pG2gN18c
q8IvJaeEM08snAi1pCy4Bc+qbAoOp27NGWQPZ6GPyDpi+P22tkz/BWxb7foG+QxL
s6h1aFCh1QCcpkURiTyPAHCli6c8i2uvHPn5AvTLGCNVcZGsRDyJOy1LTa7ClF9L
hyAK2AIFgBXCJREn2CTOCF85L80Eih+asNBVmxKBL9PrNYAPnnmanKyeW3SDC9es
Bw5dRNnyTO93uRkHtwkLKaCmC+aAsA0Mf/4/Ag3XLdBWYqQFFKnP1fqSQ7cUsnry
YdaZ0LdBAtrg6lQ5Ql96yS6wUw4YTLtgEL0JW49K7Epn2hSR3TVmIH2YlnToa00i
FtdqGjtjZzpmfGRVMnZWvcnxvjr9NIBG4FeexhTHctcwrRPMt9Cc09lLnTufgh8g
GyBb5xn6s16MnAm393jPB4ity1MnktKFbiUucQQQy0c0eWboR27SVzGJKoQ7hr/g
s//wTNL5BHHpX3bWWmDxi/lndTwSJgdnY32OntufSAmlmWUFa2lgxkxk+JyrmIjP
SDJIxlqprSDKawI3PSWSoJcMsIndnS7zCuj6bQR0L3ag/PPyqTYMDJ57pha76a9V
Y81DVHcMSRdhCsbdDq4h08wBEiEpHKY57OK20JWcalah5MO6kWSP/nhX+Le14Cxu
AyX5PosYmTAzHyJDd6vdxX2SOgjTF16hhjSwMfCzsZG6F9uHRpf+bckMDw3jpVC9
ztYI4/hv+NtW9ENwWf+QC3LzenltjVCDg2e9Hqnirlg3ICGLSszqdd2vjvC6i26o
6qFnX2Eh+zV4EaFpi1L9Ou4b06XjPZBwj6zfxJjkZSDyJzJ1wZlLG4g5A1QtTF94
zJHs5hTmgqA9PP8Kfv61PFzANihsyysmX7y01Xej+e7flm+EMFcOifG2gJHGwP5E
uobBYJOPyA1hiPovhjFAYWEB+WUHxEHY2erVAuVIvg+YW4lE4KuttwEAbZqPR0zd
LDazIbBdBuekzUGIDgRcqCne2minYZFnXR65V1YsOjewdQq6+c83i+TFslG/56fp
xI5KHTk8UoziFt0GuMUjFpCc2Nt7WfMyAeZnxSQyzR5sDIGLjuGoDI61I+0fM72s
xYavDPLg3O48SZyxwdc/nh2lAYsdMg2VJ69R3glle+oYyJYdkYWqYsFECpsguglz
lWZ+B4uhDsSIz7autlLVx6dXWDBJxjsCG+hFWmk46Rj6I7KbdAgPBiXjzLHo28Wa
zcI+ll2wQUCqyVn9Hk9W6vLfs3tUXKn8qXUuXY+eHAgZIokEn9NdMavzR+ZAAayG
Z18G3zSGQmWkhQvBuxInWNndIRY2t8hvxpCiA+rxgLWCauzS8JiAE1foyt0HZPe+
JzUlypqbntnww9BP6aUT0rkKnH9QscQ1iCZHR2A6hv4FM1swLicythUMQcBVBRg5
EM3llE1b6uVTNt1oecSY5J6rNOyt3eKFh3SE437s4eDOzdObLq2uBgTFoiEJxQGl
m2A/uC5J7K4bKAk1pEPhxDfQPAh7g3fNFrpG6IAjfl4ImwUe20IgwZvVvIxQthNZ
zHFCEC4g/DcEakGskO3yjomMz/4vkficpAIjcZB5818aY7qltce26JoEcQaK0quD
amJ8tHS1y3A+UcLNDbR4To4QYJ0QQzy4FGxjPrtgCZwAR/XWVR4Xn6ZCP1c4yvd4
BMlG3zfQNw5QYRErF8Lu7qIqVTT+NxF7oRfOHPIrc5K2yuBvMeAf3BpX0W5Z1DBi
KxT3IkqCubktVABxibwTgPHbYDwbWUe3BfXeuCHOz4WXAe0TGDStAx4P959vPddn
aygiGlRVzIcmk3062mFyNGgaoGpiZZas3IcbdEV/wWyFfKCXh4z4gvTOryBFNbHp
Fg5eOl5DqbYFRbJtAlxA+HrBdzJUTT8aINsJVhdyTQ3rulVU2SNIpRYVQV1HLOtD
3Q0I0hWdEXf1ssxBJJQBp2I2LDMoONwO0+rlmFuzCisf7hwUEvbGda5FUL8pJ/j9
F90EszQZcWCCZxPXbiZYzZbs0nD+mTc1QlCCtkjBf4RSXkYpc7lyvpH639EIvFRV
m6UPtPuqifHjAImNnnbKIVBoBz0NphFlSiAgxqeq8f1+RF4TbLtxj2PgQRjJG8F3
HwYH2YlKCW13vDkZGkkk2ljf8O/2ATFFW5JJCAcpTF9NFCP5OZVN8/+20rwbgRC2
YL+CsBNUPNFDkahX9DQ3Zd05mzjLgIrmdXQHI+fimMGaK7/O0Qlau7qoMhn1tmgH
XpPCW7VwHVB6CDDKbvjFowZiFPCmWCFM3b3/Zjd+ym1ca5kDLDTYbjfaaSQSt8OZ
uGw2t+cx3xER8z1Ucc03sZFNosddLd8pnol74KsIc6Vl7h+8FAUB1XEMbCedhXsS
wJ1vWnriJiicUoi3at9TfxWbbsgzhudHdY9HFNEaPZ2fOpZ2p4zg8ck/rbslwERl
N85mcjWFuEcsyjEIcVZe1MV5DZYVE5oKvorj4hKKD9f/I5n9ZWnhfWGwI6YcMatr
rlLHLVxFFmayAeBqx91ALhVwWyvHCcgVcFEaQXYs/ShKbs/xnHeLDorVSgaYo7XF
/Qr3xAvLd0l8RC7MA026Q8XGZbecdeIm15rcQ9wWCv2Q6ooC+7nr+sPpZ8ychYvN
Cvxr+jH1Iy6exksEingog43VcuxvK3+a3qSXifK3aVTs/Hdtk/tQrJMFRSqLTz5u
f5INd0R+D7aRvU49xxUC2dCx/dI/tAqM3oI8+Mh984rrEWHhh/9GX43Itl18fiN1
3d5PKO1iFVB+5TVfPgqzsxXNMF7YGnS6tPbfg1TXuVzDy1KQ1ddcAnOGy3yjGFTI
VMbASioyHp+JTBc7XummPYU6D7h0rTTcJKD+GPSrowpj0mncZYnr74LmoXy/Gljt
keYsAjyNsALHy38nCHB3YOz/sNTYexdmR0kyowLRP454lHep2rrgxYA5Di+et+RN
4iml6L0YRUAcRCpNzxAIdr12WN6hqhIvdYA/pnmqH623qN/FqT4T4aqaSuSue6GX
3KDjXdi0XDMkwaMXP8EBqv6XRck7WEGrsZnRJjj7BQ+PV66io2QOkAEcAlowHclk
B1nv74CsvelkeBK1Aqgp8OY04Q9S7o5n8PAqjXoq2HBUY4fHt+tF7bAexiYQCwnv
zv7JOuSdjeoqDC+Fg+0hBf8w5EymAGkcCG9Om5hbbEubkSvWmv5HgyZiN3RQllwA
I4osDatMXcNjKyBQOAhJmT+UzL/Za3R7y6AeQ3aKaWE6OogCc54iMz6ix0uJHJqe
7naXpZ/OYZWxG/FLrBd67aaet0F7rYuRSIE6Jt2WPp+rrKrVTGeO0NLeTmh9tFZ1
XLIAac//fqtvEswOodd9D11HSQmIeZwgd77yfupEI49WUwKrdT0ETyaDqxZ5jciP
9x60PLrlfiSpR4hFZz7pNLoOsj+RrUxUfY/PfVpGsuCHeAZz13TaaHz4YJnb8eeL
ClawqEGkoDKmSF71aNwHqZLPmqGhD5Ah29b/iGsqcnQzXa+Nl7XBwN9aw314mxVI
G64GUXQVOvlGrYP0QoUxYoJQYgQnzZ0Qyt+js+JoVQmNv6P2VHVXjvywoKu7R7gN
4B/sf3K4KpF2fxyUxzsW7rWYNLizxPq/LDnvbeMHZzWV30b5kQ8Y1TSWccu32Vnh
8QRLvHgOF3mRazSBGKG5NVBUJZylAV4RJrRq7BaIlIPZg8JtS9rQ9MC1RlTp7PsI
pdQ6vT08TspaPtODbaVJkcCvOTrl8XZLVvyeT/Pg9vJ0EqHJ/Rpwjy+nnJ+JjiKz
EIBjxNb2pVmU0GWrceacubBXE2WK8HCKnWRs0d+7xlPJmTTmG0Ep2neOt/2sZo8x
Tawa5cr111cuuQ2jF2vEmLuyjVasPAH1l3xsWjSb8eWZgp5HOnJmC3eycwCxVEXB
T3yCPH4J9nx1U8uYg3kHBEIjDSOvN677Wkqroj4Cxu4r2h5PfLQjpfKWC9QfCynL
OAhhltktd8lq8/QnXfgGMPVSjGanoOxcsdsHebTZwUMdp7e/zJ/Vyi+l6H4Y4V9E
0kQyV60oI/1Pcevd1doSEuP3xqILS8prlhfHDhwRSrfCHyPikVQrZOF2lxMtXiDM
vK3UyVezupkCmAwcjHZR4saxS1QiTgARgMh7Yh2BnN9yCz2DG1Ve3hLXuiNTJMoe
nwHVh6D0DKZ2NSyahbOa40gy5uPrzm+WTdPFxHp7rtXhLvQF1DSJ4KW3sO1jTqLf
yRcjEadCI1pqp/PN2BMWsnUruZsN3lFKNKefoc6kzy7zsavxstfiOQMq6zaUjCyV
byNPbbYcgGAE6PMK96BLrRHz42rHjB0S/t+SGoOarePPXzc/B6ijnRea0gD37L8h
1U616Zk8QuaoeZOyGsOXAuCQVCWC9o2ba/RA9M8jmVW3jk3xM5TNapVOkdM/u2IV
THr6PGrBhiRhEQba97Dei0XyjfEpm6BSeR+Ngw9kdUCZWBfR5GCSMf650fLAyYCg
/V04T3CnOKguJ/EBAOSSk1T1P+q1lcW7GISqQiioCg4kUuPthn9UqKxMCq47ndK1
QEHMIMjazz4paGJFjpKu7fIUPKl3rb1PdopDgSp76GCHest099a0hrWI7xz6qLtv
8efbHvrvTgeZCVzCN0Q/GLVBcpnElISWQeTsMeKp1qlwDieAZAKRTBmuuoPDlWfv
vJBgiOUwjQkZrVPEMr8yAujuzi+eUfcjxoleKaQ7yAvXsCpJSuj1BYDiOZIXWg7a
IJc0RkUpnBbZSZZ2mDATGV/AoYwQH3nswgFi/7laKdJKzMGbWnX3TplWMWQmH5Nh
JjhOdDqClpa9MuJ12EPbYhmRe8kscro34JdKvY/ueLp2c+XeVYFqCJtAvq2Bi5rC
uROQDOdIUig1Q4u/Q9CtHH+hCyQy4VnGGQ9ahrzDWby1mm+2hlV1zeyurKrUmmbw
Dixmz7+deuO0Ad/k5tIn8UMK9090QwjsqpDMeuy0gxbxOpDSYVI+9JT73B1fBgen
ZYEcwE7AQc+brfBrPf1x5OgPFmbPrG91bPHvZxQOrSH+NdAKmCByV4O0foD73meJ
CP0l+xZ6dEFZHB13SpPYkPixAau9Hv0MHvysznyHrwH+TsWuJxBMadrjY+fLaUZZ
gbMRvi/5M6M6W1ZZ+xU5GduxvMsX71YSuHnEhvGxgk8wBWhfQKmhMdnMI5mvNsWM
vI9eoaE6ejHAWvPBfoBEzRMl9RBf2NLoLIyYb1M3iOe7Y6R32+hHnbaCygEMFRCS
oSpWzaq2D7LqDJkQd32ijGVC7wRJoNC5CVU0QB0X4F/x1pKHIueH9EV/aaAnJ5qW
Ey5KdZkWK5MmM2cvVzC2CcMaHyGwGmOBx7UyAUPqZKWdI0z+eY78mj8FfD1xbAjm
NBjbZtb6lS8CfJIl0BhA+8lKzwJ2a2zqE60diiphCBYKMY2MZ2tXTG4NssC13xsw
nHaF5eZpmXPan8kYN1ctG8nkuiXK+1hy5jyrHrZ6WIdjbony790mVyvhY7Scsq9E
90x9U/P9qepaZsUHzRy5r1f+tZGJF+A+TMjVH/gcF7STx52YbsuhawG6h4vab+XN
rHzbQcUD3qqmyJNP0InZHPT3NBMJP9S7hyO7IWt8YDQRJF8E/DVv4V2ojUrISqcY
qRKE78aCsk66sYZiHjWHEcLRXtB41AjxW3kgjdzkstses+AlQdq0y0QjQt1FnvHy
dlkhWSmDKfNKnGOaCV9oGkJKAAlIGcEyKJmOhdj0e5nfLt4xbmPK6tcxc68KBc+N
sGB/fBKhb53vs/JRjXRUhgoEnu7auYW+AsMKB3+3EDS/g4XLISvfWFGoCAl3CCPF
MZ2PBxLa460+MI2umENjhL9uQ1SLC5dlYnKnlgRL6gIHqvcW8rq4mOEsJJ6oYkXs
Qy/wJjSLeFSRL7yhWg9tGJ+St22EkGIzldmz81SBxEn3knFYHU+lgTwTYkOGK/GS
PNJGlJ3WfZMea/3uGMFtJS1cEM5Y30XuBZAJ2nvE2FbhK2qLNhwXwVPbtgH9x3Yn
Ha1SxWRE8LMZGo0zmY7MClnWMJ+YX0mZAdS0nVmty3fMSzPgRREGBMq/4xiLQmc3
0UrD9xW9so6MLPVhvjUtqWoWf7zcNqlwjnd/EytSHu9U1gNQJKPXznCbfdM6UjOu
v8bTQFNdo5SGLSNJkbKmkGFXkOReOu7M6XZpQvSbMgyYC4Yn9PDRtuT6YztIfsds
/Y6fUsuP1yi48GZUOm27TshQb/VjR3fKeJiwRn/0kOr6xkbxB9N1sRVLLI9ni+Un
67SCG+1HRqTFKT2jWJfAnlbcZzRbM4ereUsS82tohSoFxpcro17tpsLkLMVOqHcN
tk3czlQAF8ztFHfNq04KEpeEHpeb+ifDR9+C8FlIjvqLADRP4c2VfHa6pZRiTdTP
w826JXXb1LAd5BUFcNbreJn/khQAVckogxGdw+03nDHX8/VV5OBTEMaMl1cqm+CU
YXI9J+Sqdslu3P6mhMojZWGXPdZMA56i5XT5fjdz3xhPi0BA//hIHWSj/g1+rbpa
SDQkjJWHv21cNVZYV2KLD2EnjLKNIfN8d+zxAdDT9Bg0zycUONpvzb3DsdKwCp7c
aQfMEirUpIWuC8ybXJAr89whhYxCzumUk4vnSVEmIoumcVRSK8pRxjLdY9J2vGGB
2TyIEJrJX3HK6cNW4uK7X2lWWi25H2k8gcwufsMgZzl+NTeKpUG0TcxrIBOHuCmp
0AhHn/9VVO6DURF8BbGTzpgRXyZOYzDJkArGSUd6BxgxXdJlODRa6zOKW17/uJ6c
AA3r2R9Uvp/F3Q6GBZfldio5ABkkf8oFKlqKgrDUZa8VRBCqWJBTxIyjwoD6AdpL
CYe9d+tI9tErdWGiQ7U59jpxmnH6+1jjErVXM28avkTCrANOQcb0pnBaO3rWQdf3
jgaB87oKQCA8Gf8mncSl1ERtAuo7qNVgW/DiM3jVNNfR1LbxcwIRqsDuKDsCgJcf
ZrV2+iQRGUqPpyXMOYL9KfIc97ggdye8mfdnqT1qA/au7dW3OKbpO09SyJTl1Y9g
aKCks5ynpeK5bbK8xRjGediTaDi3af/oPTfrqesHQPkf8a5ba5JQ++jH1pfXAei2
bq3DP1vb3FK+5YxpQBu/ZQEbANrGM3UskwXM/si54ZLWPPGs0biImv0sznai79nZ
ezXqOrbL2t8SaTGTjxCkhuTjllo9seHIVrWE5aYllJ1jXgCZhCjvupMbQLxYDyEF
G+MmrtTtT3/MPkqkQfEM5ZtOKq1RrIzBj3rghktbuMXK4uax5u/1TVL51AyiTArZ
oHQP3DV3Ajaol89x3N+IOE5hnssJhnIFEawnOR4cBa7Eqcu2zF++yLdhx63GySrs
2TUKXYZyW1S0fvZMQjR1Z5ITNvlwvf65ldvBkF+qyqQvOvH6yqVl7+9NRSsN5D36
DpvtdQ16gCU/aSiRAeE8yEB1w9qnSQ/nNS1CS6fG0QBa5K3NnQFvaso4Tpk8Kkn3
oakh3ZVEVGIfkVLHXk8tUuVPytw7leF+2DP8iS5reSQamRPZFIcD3KqRg4Wgejqm
Gbs99tFE5yxqXRW6XyrioW9KRbaPEtwuUVaZ7NpPZaZrUMch9weJJuBegVgIhfMu
s+P/7uWwIsBecLA7hCmI9JwVf+/jGTzSAcrM0+hPYBXJVzMojWHAc4BQdwU9WxKK
id4qf3xxiXg4bY6+Q06vJZERl3NxKHTdx1ZJyEXGZ8VM/ehQImX7VEC8VhmClgS0
+lNJnaH7o9JoMrma0Uo6n/xOVQeWWyZLvBe/ebFoUxBfLA7336m88EOXc6yCKtII
+kZygrmTOxRdS/5QiRfE9nIAuzD+tQYNcSADPUw34lxorW7c/jXF/3yMKHnS7vnl
ws1NwZzW7RHbQ6YYIQgG4mCV38Ay5YqJx/MF9gdeild4TiRoha1DD0m5vltRXQ1O
1X4jqviWFk4cK+mw4vkNEA7voWowIxsjcaQJA+Tum4aWJaE26VpvTCzO+wbCq977
gF6fJX1KR30ql8JrKwnTrbZFBYf1ZnIA0c05EZgFYThM5AGXOjXI85/TWdraNOX1
B9i4CYBQNNNF7nBOKMqUoIOONWYQmLkNlWYqdZ44cv4XaR1x0jO4xe3tvkN/hg+V
bTUyJQI+XbIwu5QgzaJ13DyuTvJjeVEV+1ecQa0FudzWKGgTCVlv+ctm/WnNLJ8U
Rl7h2wqPX2xHlggdwPWSY9haA9BezkqkNR1tDkhaBj9tovvNTOqoaojN9G97qWXz
C48FzbNQqiDkoiwiQpcUZDkCfT02Scm3JQMaaUnUFGXThEfZnJ2N2NdSC2Seqtir
HEsBrXAoA4emfNZxpX2B25Afd0tJe0dgliBHnsgLrc5XiYIIcISk1kM5+mHnNPMm
kdA/Pw+1kU//Ct2qw7xSSS4BC2A1EM9kUN4156bw7iABmWXBFBpDxU1ykc2Z3p9Z
kstFUx9WkrYyXTazQe283wNUb+NQWm+8f4IzmZuXNuFyUNV11xVMlu8p18DJADuk
ntafi+DeTNq34YXLjGOHh9VGYGRfXV7kET8ZF3iF6kily++C3MnDS8ahf5szWK0O
oGvsqea8prD7uiS4x0xY1D5ZGIbutAVOHczuyNttr+adoj2EarBW6Ld9PAlRd8oh
Vy0AntHY7mhImA8WgURSTXQ1ei487dcU1322PZ5GlRxgSP+aaJo3lRwOfbK1iVu8
oZZlBmgX0Y2bNyp+5McH012H/5JHnklrqIYnwahwVOZiSZvBdIXr5RnLtQ/Dtp5G
2I0AMPdzTs5mNVmbKkAlG+o58YmdLKoinivqXFvZ4AKKaZZ3zrbUe7qnPp+nbuLM
npx1l5izorhqQkK3ZOakgoi1k4euRMvmKuk2mdc3OYZ3yS+NrZuSfeNFM+yu1sDP
LtDy715keJJ8xQXs+YkL+W5t0T+2rq9qDm0c9GRNuIiTlbSkdZ7pR5f4Td+vA46c
+aQNSNxSOgHwkUM1pMGuCEw2aHTS8HGs1ACWQZXj37itJSfYmD9EDPEYgNbio+AF
TCNDyqfRAB+spf0R2HV+faz8j8bYzryNpvAnUhK5pUu3skTqnB3oX9Udv+MU53lw
c/qGaBl0e1mX3AfMjsnuJxz0Eb5PEPNfObQeaGG7ZZGkVVbZ9QR8c+pU4nBjCKE4
DkwfG9N4YwkPOcp6GzBAKl4FHspHk0n6f9t8YSR/39HWL/lBM/B+hLcCx2M88fkk
DCJ7CHZeVb/BySoL5zkyKPLyYfUr763m4u51PMw/iY26TspXMpz0/K3MfV2Q2NKp
KVfOJmAnLMJyLxOV8XEzwiahPG7HJR3KFR1Vk9s+K5SSPRMQ/G8f7RDa27rcAjvR
dRwwod6Pbbi4O1Oq1qigyrkaX+tT8vMKDo73Df/aWFixFw6Dyyf+pUvp6tEWJ+WH
O0Mmvv73/veyCgHkfubJ6OVzL/JvkhfVQzdcv/tXXvgJyFHL/HiZVIndoHbNpe1N
fbQW2lzcZHjS9YFsR8Iy+Akt095Es2OK+9fwv1XiQU8jqIc2wyiGQRoorgNQF4ux
jJNXlwogvfAY5DGW7mTctCguaJoWfsgfPIdp1WCHZ5zvuAp6i/GPl215mi9khse2
Wj1FEeK3xV4b0h4tv9ZtkDBZndHXkBCpvn96nSJJz/ffHIe1UqjVV5bki9TtT5u6
QWupDXnpMZCtVUj+8Abf6c500khy7WRkxufyjvVBieIAeX8wrNF3mB08rxu81HfE
VHoyre4J8zUPPkqQBIfWDCXqjxndCM2yWht5x0zIqe+NPEGMgn3+9T+IULZVXaKv
h1iOZxx0XfEi+tlHFV6IsAcQ8rD+3ppa/M/O+8sCRuKch6bHztEhrQzQ+3qem5HR
7odovj+eLMw/Ypd6G/tIEqKYghd0trg4lKtohvPQ8KMP6V0AGQ2rqh+0bDoeADBR
h7hSM99lvGAmmEujGERGKKuBbQZPBRVisrnNBkcPKFy1t2PubUL1UJOcz0PUd/7s
nNfi/N3Rr8odrhSIgci63HzXqRciMrUj6ayft1PL8dlG17rXRXWNy4yA4fJ1qkGI
VH4qpq+s/FBO6V65M8i0QHZju0dQWWzvMvNn99kohQoaLTvuPwIUiRc4/aD9wtn8
prV+iMDahD8VLvhVsGoazBiD30DLmILkDkWWUyl4dJdXucMH/8aVA+OPzOuziPg/
jcAr65wqLumAPLK8yPu5DQrBe3v8x//H7Tr5ckEXUQyYCfFe+rfev3oytyzuZI6r
Qlp0AMBY9NonkV8mBFmoTH1wkqV6tgEAqjrtgGksmmTXc97R7+RkeOzMScEVEPgW
/EwCVH6MLuXu29cyckYMZRciEI5qDJoTBwNrzzo67YdFbFv9FGhkoqTcftjqe5i2
XL/CDx7t0QVT48CfUJLxlKNrweQIrGH8zFC4hnWliOZv6t5SC7jrZw46mWP+j7q5
6KSy7+/rW8zlyxQrQUzqxYfVCpzsl8SmakcqF324WKUlGT6bc7UK2IWqP/Znazwq
dFwGSlMLM94I3EUY7eAoNxbX807nAY51T4a4iSClwydGOLTlabex4vaOiWgerl4w
wjGfipVQk0vC92wACyydTBT7VEqndL3q/O10tgIyT138B7LvGplkrwDZhX0Rb8yT
oOr9fI5Prnb6fOkjdux4q1xeE9+X1IAD6eK7I4LD+5ilLo2leWFXQC+HJla5h+9P
uRI7T0VtUsZhokaGv1lsSTht35KZfMiwxZ96V5EwUiMwbpszPuz4QjuWvcaDxl85
t6B/bAFuD7DlJIZDM6hQl3472rd4q5GUgysyKb/xr90rDc5uHeegtiJ8VOecL5fN
vxv2Wo9SK5KcDGJxT2VC4ZyVsWxNtEvKw2MDXdOK9+9GBpQWOdbzAMoCg4DjdKrF
KSDOvQKqzXRbOD6FXb/Q532hqRKzqqVPAVEpvRtfzTIv7PdCWMHnKfOROJXIc4Fu
AXRrFbCDglhHtLz134oViOIvRV4q3wzAKvz5gxFLTKddYAUtXbexXw1muF6voMjf
ROjofSMint2oPIka4mUdjw3VY8Gy7vzVsXgP8hTcz3VG/xMebxieaMszOIflfp/Y
L4+wc2K52gTHs+KVvn8eVF+KphZeFhUBJU7SIdvnCFxcMzRY5LU+13gzPpt7lOil
bZOzkcEL16/U1AShd8kgz2Qua5qeg7hgcWfoMLEy6zW4aUAzaBsQrR0fPnTzNHbD
kydKH4np0Rc6vyUgGImW8ff+I2jv4kTI6Qd+DR7s4RpxXLrczOVS07qOrY+T5Rc8
cDqE5ZXMY/dNK0n2lBlfB2o+iHQsyanh6JSdGev59W3O1+pq1VF3hTkkmZR9kXQZ
xSCqela/W7+Bg1bCAH21zhocI3rNyXM7nkYn7ItIOtiv5k20FKczZYq0ExDKXLas
TuoPQelCP7XYLdfgwdjKueE4MfoYPJ94h1fqmgl7U1C7uZ/kYkB/qXV47osdVe6g
P+QrJKvoX8g5uNgiCIoJEgA7QWF7eFN8BR3Jmpk6kV2g+OFGETXM+0tzbdi/hvm1
fkuhB+Cl7amLcm8gOe/095seRxCMuP+a1JL1E+Gmq5azb3ocNx0/oUML4Kghksyi
1gXZEjHcHmlPKGNYcp2kAjqt6pLbhAtPjuNLYPhsGy3Yr/Wx5A66tQWJftrP0q6f
CcfqCrkLJhXZ5Vj7yVOHX1qOQR0lrpDc2Zdyw3Lu7HHXjulCJKu03ElF9dEk9RHW
3D2Xakr4FYV4QcqmpJTCSykXi5QJlCpGq1dUzpYBV4QVDEKPNNCy2hPQ2t88NmXS
tdDHJQGt41KUMXAmeeErL5/eD8vtcfiiDjGXdhDK8EIqWtVYklZbBege0ySDSZzs
TWvn7ey04CHUKokOSX6CbrrZucXUBRHpY2j0YOVct50ArWYfiiXNodaab9TrV+kU
x9nlwLasJHDAX9g7IEymyPxen9ePP/BrmmFXcHMYlaP0xi6R9WtgXhdUnPPtN3Xw
In257cTWRizUIpl6wMC95YWScnPpXeYV8aqcInDPi8KiOOhB6PAuRwpBAuTAFisc
iUy5KZts5/0UNWS70G62ku2Dch52SQ95rhiAcAuvOvRlKnBwvy3PPlKPxMkplCNo
rPhn+kxMY0cussAsrT6RSEeDQALKYnffyxHAN+ktBkA0WqwRKX0UCIx2rEm64iE4
WHlPwqLvfmH5EHwV0lhjpCqqEThtRWgU9aoZVz2k7Lm60d90g/OBNUlNwZNQL0EV
5dLzHUYdMLP5hAHWJXgK2YjzBJ5Q5KxmyyfRunR3SKmhurfROeVyjw3U670MTZuf
pR3VqY5Kkvn87zXThcUwLRS1vdD7TKWc2bBtMuWV6eXRXCtTHncYxa5ZCs3bqmvg
1I1GPL9GbV4g0+7bkTXIewM0V215DLnLJOydVh9V0Du7xecITsRfu1Bu3TKKO8Lo
g+DPGmno6WAhpw7oQHsW4rxbE0RPmE0gtv4FPG1JtyLuEB0FebpEsePHTuN9StP8
wA3dkAdvZCK6QWLHmZFyqrHTyFaY/+b8y19wdVRkOXjgeVyQMcRhyVqspp82D1o+
5YoaJ5AZTYBO7Wod2Urb/tO34L9czC/iiTSBSpr+FwXikhpUfA2nyOaiL8I5lTnb
1I6n9gtVHDbX1MBQqwprrTjhJOmVzhmWq6VNHtTnVkY78FJZsazys6wrlW2VtZ5y
jKsUUz543cqjngNzT1WVV0qudNpq8g8iLVTs/3DqICBKRrqIOmy8z65RmcW2MnZW
Xt/8nOjVbyIXK3Jgl9/mnEa2TIx5NG7E7Rlfzo0t95E50m3PSYBpDqGfrxveu75A
xH4J/E42vVzMgmwM1XLd56IISNIbz6hipi1vN+KktnBqs9ajUhEVOM6puxisoDVD
EzabKHYCCub/nMZerlVD3/N0YgM1xtB+0zTQ5+DXrRUF9Tn3Xche1cJ7O8zf1yib
Vo2nvW6wAvAZl2rXwKNBt7oACIa2BDAECj+deXiqLkLT2qqiOj0zuKSBd8gvBjD2
zX/DlLGblZxv6ilVFMVKurkZpFnTR7hdskZZvSJ7F4F9ZzIM701hn6fvRm0onnX0
44kQt8tP8PDtgdXEx2ARtZTTpaElyZsj42y0YBywGLagGq+F9asYT6Zl4fNMfrZ/
QBcnqJlCJCGB7gm7RFX+TkRIQbqbN9b37CNJB1COLGtX5rXagHlfMNnE8MMvI79h
YCfP4EkusJt8AHGQFmvE5pEvH5PRuuCTrFjdQe6qNGlCW6P8vXBCRBS7PjCj3yUM
d3+JkqrHbsAWmXmf28a1RxG7iFRCab48mdh7Qa/3o3sUVGECbwbXiPX30uLGeEU3
Y6N02ARf6H3/eaKwnI4+IYgrBIlNB9YzStCt4nklQ6s94ZB/nuQZ4Eb//qSy9sWd
0SMddAkf6qqhMuUiFVEqqrL/yZmPkdRPQvhqO9gbjzQREHOhJzOOzIkaY5k6/Ds9
ubzkx2RbQ/ZGPm/BqvmR/Q+XRyyNU+5JB9ZVDIR3hTlolQU2mL2i23CMS8j/iAby
Gabtgl5pk48Y1lD9ewKgEMz+8BSPjqrybQ0/oAZPC4qw+Vf+/P9DRZD/XCITHryU
p7tICpHnriyd8CdBts1mfJ9eN5Lvbk/+n6N84U82KJP9TElDoIRPSvhDNgDe2WC6
5AA7nsZMDDchmVyrX96csSS2KeNZZrsWT85/10HcRI8ZFJKHNC9E/dtYgmRM3URC
j1VPhnpYuhWKcgSEGJiyKjUM198Y+Zj2JH90JSRtQS9O/ekSBiYwi8ak6gQo6PEO
61ve9Fiy7C/qsSwVLxHkxFU6Js3TZuuQT0855R7CfAqJgZ4BD3hD0dQaSgfNGayY
NGBh9jx/uPf+W0g8asTadcni1DPuaWampum17CV5rHYUsCwY6tnwn7AD0Evp8ajf
Nhkubm2dg4mYr3zXRkXzfZqbQqBCiCfC1WqmziTb8YLTFmVeMEnCzOtJjMYo4ydh
E+281bQ46HkmX+8dqrfiLssdsABvh5zp+7MIC1yFCJV0xoQFo8K16EpoOcrphl9e
GR2slKyB6vHbWQTHYHwSlHW73x1I7FGOX4VdOGmPR4QzeGlzGs6mAxk8DfD39f7g
6ijf01f3NlV9an1fqIkYQN5syOUINOGO25fmIcqOkE2BbmO/NQY+cTUIdhP4B9XZ
YhS08ycmHQtB7CPb7FacxVOWYyondC/QTRHuuooT8/vthjWzlqCDoUjdx1qY4lBG
H5AKuDHbcBtqNodxVs1pMXFICwLOHTO2hdbBfJVTuVrZwD19I9F49jw+WtmW0qcc
/9bHfCPkziwS+jIInexKpzcQiuMypjw7tqinDxfr9kxa8Y/Cvb+GEHiEsUgcHI0d
FRG5NeRGlWfGt5gMlbf00Y5ACMVNxG5r9CvsgFwXLetyGhWCSXx1EUK2F1mUCqUO
Uf+wwGlp7kxqPkvszJ1UkO9tpiNF/oXw2v2FUgJCDFgY2viwbsHRq4kQuhuwgLQH
pcnQRK50MwFNT1ghMm6iLxx4uLbQbXs/WQxtsu953yJUfdGCIrCMFRQI+6bPq8pL
QJDh7t875C8xijb5Y6rqyfvqPm+RAWeSC6zDCS5Afe4npN+CIGSqOMmKfV6Xzpvz
WhhQ/X7q/kOT6CwdClMKvPxCNXQjGd5Cs9Hzix4VkF+EJ4A7W81htfsk+cjjBYQe
YGPakjTZ2+E2oPz6D0h6YkzHNNCT32Iup8BQ8AgILDW9aLG1AGHlLZC7VkJeOYnr
8WLEMwJtegvi8RULvbKg/gXKuwI+G60T3WhT+VsqwczD4GYVvPAdcg0QNCIcpIh/
awV06qcf9jnnyWWv1uN5iYEZ+Cozmy14ONCOXdJwQnQ/sGSMM8zYyngH3strRUPW
P3prhFdHujjJBfP9EDG+nNx8Inqfidx2lW4f4OxaPfeuH5TQv1pe6lv6h40XpU++
MBiOzUCRxeXhxCzsImNRPU9ZPZU51GaqhR3ClFJ8wpZA1Q7Ttr7mPocviiHJqZDg
0ToWpWrZD4UXOrCOutSCiHXAOIWGzWmEaBcSHl6Bj0/Xra755nCBc/Cf4fYxs0Zn
5oVxdKd+M/dWQMzV9aFzIRUTOFhoqJqttmn5Wrgpp8soSzJekZ9v0KbQumLvCxZy
IL4PP3OE584PuFi/tHNMmkD5Uv/f3Ai3Ht+cK+rdyVQKOzL5ZkKpRHTRqkLikiRa
8F/pbbQzlaCpoMAHiZRBJl5gi/m10zEf2Mah3C3m5epMrsrB8RLNW4sRx37N85EJ
iPWzfzVTlFghrOYhOu+U9q3qXvEtaRhs6j6EkwWJBjTsU2LWsM3dQDyesXiz5GK7
F9z+cB2gZnqNnj/8b9FJQmfKjyv6lpZsw6HOkO+sfFglyPLHv6pm9pPWiEa/AFcv
/Y4qqDQGBFbPgA8+XhaxRv8aOZso0j66IjmgFF2zNgzDCTeQw/Ax3G9Aq0zKzRv6
r8N+B2XMPLx9iiQTcnMo+2noIWiYTswo/+QrQgxFbqU0/CCXhi4mTMCXJ3TUeg82
LeEzVq+ZOngygeybB53u6qiM3B+VIYibdec6CHnzVc2ZM8vPw/l6VYklls+W0yj6
YwTOozKpQi+PUFKsHTSnhQB1uPyGeUYTwSuuzQICBNxPr8+GkHTdzztC1xOjy9k/
ho9PzOYa9NOWsLxRfUN+tPs2wVuBDcjhKAYRF06vUa0vQ15Hmua+OvyXU7TZQOkd
tznFe4KsnPP+ZiKmItXoM+PFjgaYbYr3NbP8R9aX38QJJulEuRGvVkE4yHE9FmhQ
lMExo5oVH9o6tj2BSm74UnUU1vF9AeclRQlDdp9mISfD9/edwcfXS+CAUfYJK3nO
DENrQRVeV0xWcQmUviyhbIwP+5hknyA8XbsVCHZwc39t8Wt/O/NoMjOc91vemI6i
uxYmpMCgBknEI9lHVGSjf8V2Ld3gPZjVrUc46pVVDbr54+Fx5QM18RlpvoAGvrQ9
sI42aGs4qO7x3kkBRq/3xRA5qyqixntLisrh3H3MiaRKAtFEr2K9QKmt3wkbXCuz
+Wud+q0DBTNAtPb1d2XF6VuCp9LG64OXnrCtBlipxZ29Y3P8PxGyeHASjarnpftC
Z1529j1xCsQdgX6wU/5v4HYP7mVhtmUyOmF2aGsfs6TF25QTTMiluA1js1NyhZms
FgETrFz08+NP+rL+npdMhHpVGkvGVvG1PzYVS93/lIhJv+YgE+3LgJIdYtT2yOH1
+cFhsNZLhl8sudISyLZj7XD0kDTXYj7cX+IW9Rzv7fgTyeewIYyEICEvUDbZFMKu
94j+nBeJhNxNIW9If9ZhxZSOysxnu3ezhhYzrSj8OegizKiooGA6MEWdNjM0XQCB
jvhaU+SiiNYSw03HV9a+SmWB4sbBszJmZwPzkU+l9YbgCdMFZSk3vVKXkHAcYLcR
Kq0D4htl2CbdLcaeEWdtjGqxj7sk4+y6lBlps1j5B+IW1KU3DZFf/i3XqfqRdv+E
pSrzyx1mrOOI+VSxkloBLFcfNp04JMdzbyLpohqU6QAF0zlArv+5cMK5PkMN5bjT
Hy6NXnNcvy9yXb81EHcJY9FPPARYYdUVVbYLyONkhceCU39u3pmoWmCTe3dbh/aU
wbItCjcm0c3YDyAau5/NlekDkQDs3vmox/jt7YKLLAwWyVQ5LdJqUwtHS7uQj9jR
TP+bncT7XGg49kA16qPU5ovCT4/xv7dUOk84hvIX70bHKm+y3qWt1ZdahdDpnuF+
XWbnBmSxPbMwZe4r6NTWtyCuhbFyqJeik1OBpXXgMeUiRWm6N2L9chqOTLitnEm4
xqr0NWSbBA4Ia2tsNEI4Eg23JmDwF9Y1wFnrHMwWxYnkVhIRaMhHLqYC3t3e9/3t
K98tPpZE8u5529ya3iQsBas8saa7EWeayaJQCAuwgykiJMqUccT/vudqxaoj0ztq
4m6rxbj2fOX43JF2dA7XpL35uLXjdYEQeAm03/XZdW9KKanZavmBXV/UxBS1U8OT
czm3w2M8GBh5EoesvGT6GKQ3YZUQofjlCnrwfXj3ZaRDEU+Vbnhx/7qxtOFtR0D4
QiX/KAefywa1bEP56JZVvlq4Ngb4bMFU73aqWPhzW/6emEacq2PSMl2fUpCeC8me
g72Y1nUHDMl+jonu4b2aRuE7bTF25IdtuR5vt8JKYjDSO3XsOi/eqhd07sL2fcwm
CMOEMqzLLZQeHLiY3SHGAMAVYrlgW6CMBjO3mlxDGHjx6lI3tcGKZozo98u0sZhl
DRENqHFMTsoYqXPdePHgnTwwvu3s6iQZCDLhHGTAQHSbhCihtwQa/1gku9rG0CHQ
83tZPRLtPMDZVaZPgmJKpz/o735idNlNhUQ02h039uEg3QrsY8udxG0r3eIUb6J7
5pIgT0CJG26iFPfte6hmucRsfODct8jsL3pqLezgYtFhk/SewNP1uDtVWer7p1EG
7q+lReSReWW6uSrw559Fg9dPCxD/nt0BdqPXQ5YI8yaZmKVsf3xV7HF40Ge+YJ4A
/NxZzgtrMfF7txt+CH6NDUEWpAlUkKA+DXrv/vsgXPD9CXwfLn2qAdFkzonkCkZp
Nn2/R+66LMdNrkTxEeNSUoNnKk5cL/qaTGbHMwcIHN0//xIrstE2HVYBl/TDCQrv
m9Z0rqngPqbQUi8KzxobTFi5w2M7CVAAQDwHOcrPFek4BscfRy4I933zvQErayqS
YvuNnCiqzi4ezLrBbRVHQaWSq7iwJeaYrbLPEtvj8+aytPK2hHvaCK69ggJBjy9x
Vj5gWidvsIhFsA9X7b9l8PoorC8DpU2Op5SLTLBDpLcJM5KdFau9YsEG1igs4LPa
LaPSQzsYYtPlq1kiAGas5gmkGsG0EoUoFUoJNA9RV2tUtgY75NYLRvn9eh5XaSqa
PvY61OVv6xkwfEdidoAYsdrSgChDlhN7bjeyZ6mdtia3FIzD0+3+y9B80jgwwTZV
TuFcRWf9bf9VksFkbUhz7YRa8hTBUwqowLuqjeFzOJ7k3I8ePORX+yoH5aXJU0OQ
DyOnoRSw6hMbAEHvf5LKCbdTMhXUOn6Oiwd0yZfqrenKMMNTQfB07IA1mN/j/S6G
xPmNwyAotfuBrDf+ayu8t/qMUzLJQZulml5COS8KVwj86c9mOvbvJRZrbfpC4wvd
CAkEU2C79bkC6v4e5yTVvP/B6GndlKs2HIQ/W+gsbIgbDtzZXDutRet/Bg4sjSlt
pDa5JKWQbCb3rXwG2FjG0gYuDuuiTls1EIG+9Gc5El/KZXBRwa63LmVKfIOXaODT
2PqsKOdxkQSDr9hdgSKlc8zvLfTg9PE+A0aOuLykXPsqZT/B93/J5/HCLcS9HNR3
6CuixkEKoNcqEd1ixYSTO0yOc4fEn6iMvuHtSXhdFqAoM6hFKQ0mdOOsUCaALyw5
wkiRc8BkmE10Ftk1uD5FocJfSi7thKJu6Q09f9CWM5UuidyFPxdhHJDZ0bRb/Epe
chLvHxN3qUZT8a+OiKFi1yedrcAqIdJnyTwBXHek8/VB4UPUSnyngNdpWqDIz6Cj
pxXBWhdz4opVbXMAbQCkJ+ek4X3TH9p2DEn0R+0BS8X/lr/yxdcBgrnxPx5TkREf
1krMrkp+Nxkx7JiEaQA9hOAv9Kotutd6qm3b2Wbzahg07Bge4FYLb75B9LenQJFC
8bcqKeUdEyLKBs9HZfnBzHX2WwdGaK3RPt56LhPZKiati86JyBjeY6pTh0MVciAh
EBqilUINsWAV7rOudYiaJHy4fpzpqQVGo85MP6sD+Vb2oClJyZNqegAe+BsTgmiM
Kcv22u+RHQj/xBg6Bfsb8hPRk/wmC8A9iOf+YIkDd7i+NFktoCA7HTJSq2dNGiLp
E5gBJxvYmq9Ldu+1n0wMaFvQcemgUuMemGB+aXdv2CBfz7Nf8/nuoeRbgTVTt2pY
0vXG/nd0zL52M8gxYr8w+sSbJKHQjMhnXZL7NTwd6WsbekYUiEKjxhIEXip05qOu
mP1rB2ktPZi7vU9DCBIX58vRyVZ7ULtlRJEsPRUdCDj8lnuvDTSCke70dStIcbxW
uSF/u2EZ9b8mN7WxVeUuNPk8Ccgo2nxezb3rC9b2KnjDiTwoBgigUqjic2Bqpaow
xtej47m2V4R6R61n+hK63r4a8xd44PescwUZihwUznd4Fi2sZS4Mu4vB7bPQRwnj
VzKjV1A23dQGRJa3wEtuSUSsNiJ8xyRV5lty9HBfxtBjQYX3vXOgSWAgiWfCoB36
cCFwBcQ42fF4s2t7zflMYwksIN9ypHa0xhaqtB0GkHf8imxvCWNukxXBdhNMf7nO
r1ZWfLWGoC6SSIGJZ3lUCtWw2M82JS/jHAT0p7USB2RX//WnuEguJKKuXigd1vGU
Ge2w2cNmWmWRpSEf/ILx3T3d4daAbemyiAssxr8sfWCPcRcTXZcFBSsVzM2R+RIP
30f0BkI7WDLWujG+jpA/Y5DITjMf7lWf4Za5s+zlkQA37YbmZ9VSae1HKTu33xNo
OZfcRwFYz02bpkJDV0bsQ7X2AXnD9XJJYN+XeP58WOKGGqkGay3TWzfnjZG3JtgO
6olN0KAnNjv6DhRAil8BPxxtR70tN0KzrKEnXXa53MHoVEc8+ehZ2lzsOTI/pkzk
K4MVOe7j74CgUMlRl0w0URmqYuuvJzoLiYj0g5SnKIhsnr1pHS0wLr2aDpzePgUh
m4YUIQkzV9Ip3cfONxsfZnBkPWRRojTTeag9fim6wDGKa7lsW7mSGOl4HBr1hIZQ
EApacoiubM7xs0cHfXI+sj88UbuXIB8saPnn6BKgaDuDLJzPflTZ9A3hevWn6ret
KFOnVKK9tAVKSeZHg2THLh/tWJ/8uUtYnrgIWCSMzv2cjZ+Ht+ta3qmQpnT+6+Uc
rcT6idL9axS1xuZoFvqBPaj1oS4rElRJJetaLhqlm9yKU7RzbGLCvyZvadFf+ceE
ZQ+PNaVJeZU3lAceGh1v+e5CcQrBqvG/6yNKPMg2dnCW+8YVIdEb0HQlnbwehQqC
wPB5Ns4+DtPSg2QjJdmZRXXAGG8lX9tc6WHbFAXUuCorIptHeuUdBOLJX/LQMixm
dMBT93XbfFteZlRauQXPPhlwMcKmzwOtsUTg0Ygvmf9Gnfxr18yoxcTaSBSZ9cxv
2V9BBy2CLvzYDnHcaRj9Uqyx39V4by00VwLn9BtAQYkygdOKf7U0cl+cNPVuAS38
xJ9hyQ+FkZJiPDUPEBzw8iun57jtcMNEMpRLIT5tqFmIARCMriGuWcHTh7IHd9at
JbzQo2RnYrsB2/HUMSiRfzaB4mUaimPH3uFUWzIeHWrtczT+h9vdPYhcLs8HiPx1
IvnG4sMTHuHiMCG6RYeqivWTxd7hzxMpgmZht2d5kimvQ6OSGShvgpSRks7dDitm
6Tpochi7ncxH6vqrxeCOl1Gna9fxC2AGDPNW+WRrfig8/YLRAAXkc5w3215ed7Yt
+wYJlt+RFkyuU+s7F9h45F/xsaCQKSUnzIMwfahfN7/tRlRGAOQrn/qFDkjGna/D
ZjQt98FhpTf2i9CupBlbriZPzzXA/KT2tUVsQA/NyzJYr+20awPwtmFfEGbZ/BQn
tGQyJQQC9vbvCGzXOTP5iQteypNWlG1IwxyL01FZTGyZSLn9HS+Gs0yuUwODqWTm
5sZPQg3fzVBJQNprW0KixyuJJ3TQ0wrtMhXMSFODLEhnZZLw6SQ/+04pBGNJACTt
Bvz66iX4rxTzJ4d/De8KaqPKMl3aoVt4JPF0vqVawh7FMs1LQUlI/nBImEkbUmtg
3JkpUOwzY2dYlIKhIv0ucqkF8x/wv0atDmWLTJ7kHmvkScdlW9N34hbnhxfh6K+k
W9nELP6KKCAviedTil/1gTa//TPSjZK/WiHTQKiIWBO/YXc+pMVd0WnXPcpTf4Zb
sm/WliYVK+Wn4zIvtX/BQEuh0K2m7mXo6Mn9Dm10ynikGEQadFQu5q1/owgXD/R1
6xermsGp7pA2KnWHQBEHSR2LBTrsQSVCAOsp2gnBv35tMd5s0W+JpVPsaMl7zWGL
nzqW/QHktnhUr43l65n/3o07TAOEADC+HBlxKSVfedmotoRPlJR5MHTvLjaa8XpN
KCZ+LzyTqEZXp2lmtgG7dNbgJZCJ+jUry8VwwxHfKlB+FqUVe6nsJKEjds9Y8NGn
DObtBzADjqHmPOSl8MGqBZ0HA7ThvFHgNRZtTfrhLiy5kkUEpK3mK36rNRB+wyiW
Gq2ievQ1uxVkOIhZM94tM6woQyPLwZdUIlOQ3vzkfFS0rrRcJO0OGOIK8zX/fbee
rgKYyqqtU0xNIPzu9bNrgqliGbvwS06+bT+pEJ7ohYHwp2QW1V/KqAODLE07VTpS
mOW/plOqnutHAFwaRnbeR+8Rmg375IOxu3k4YcYl0XXjajxtFuhIwOBeszrORPdh
A3chBEhzkiIO/caCDdZjly8455Ng6Vn6vaew671CvY7C6LotUToKBkdHX2Y7YLy7
ts9MqcaZEnOMnEqrgFjXeKO/zPAtFmo/Gjk6J63/i9qi1cdxdx1cmbQdVPToYe/R
MoHv2C+Bjc1qh4PSaOo+QJa9MOSfnpdDVeRSmABkKWadE26hnL5Eb40YwUs0ZclG
PM9TwsCWtF4v5XLUYjxbl2Bs2tPMq5kn0ONRxLyjsd2LSLI8X3xw9vogPPq/DShL
JN2I26zCg1krGJL7jF1Fb8vH3Zyr1l5X2eRh9EWEZu1DZY2E6342/5aNeAdacBy5
HWA0R+HGmBKG8lDIFExQxg7jN6fSTPDI18qAg8kWDbqTRsPfDE9OAgMyuDTnj74r
Ir7ucLMlBbA2v5GXKHvs+qbkoxsTJ6WgcxnEv7wqbpeVlk8x92vqJfiYag1bGoLl
aoHWfJYOXM2AV1uesUASnV11rfUQEMHbItH3teTaD9IhJfNsiQ4Ysj7RWbgo4yDX
R+JWRaqt6UwqrRwvJ3ADF56fp+LCOVBycBikVXJ5yoGvL6p2pW3FGW+2KCkinl/b
WdnOb6fU0Wt07buUTviG9csU86CzMn1crlFSoZqKOlSg/oAxqSePW1E+MtYNKDE+
vAneM6yi06yUHX/lFC7V4fGldZI5P+JtCqMB4CGC3yIX+sX4DMOkdlUSn/dQX/X9
kUgziqJuOVAH/qFqwsNPLaceyfHKuZwyxDaHng6EI4eN6H3vzk5uZU4mNppNCAfq
QR2w7/AjS2u7W/9LyRmwFUE9Du/yUH4TCDIF4tVp2270d6MD6l5jWQzHqArR82zh
VxzXpiZiQsa1Ja/k6x6C2SniKJAnVgVod8c/PB8ypj3qp27BD8mft7IZEkpY0OLc
DGNWt+XFg6mtzQNeCLTTFko1+ga4bmANgA8hKY6xd9FoJ+ciUyEYxKYUhwM2PFOx
wZ9382jJifGJ5geQoDq5K8fdwyML131Y8/V7zRJYSqvMZLrYBmM/hOm4NeLWGwgj
nmuy4rWczq3vcTeiFr1QPa4s16m3pvQM1tur1B88ceJC7QRAiWA6BGdtJHRrM4VQ
VnGlVXCph6Kmj82N8dAtV99QdQlWYRhoZ96qfPjZM9p0yoBY6cElvmssDnXZd86k
0uITHO3rkNKz0AZ8HzU/QoSNkbN2iu8LGIh/qNLuceM09Yh/Sax1hzIWVbV1cIUT
97Nh/o5/vpDoTClqkYkB7GEzWU4JfLb20CRj/jVdF3+F6Yga2MKX5HpXJftxU9S1
xzCkZEPFjSadC15JjMrlt9zoit20EUev9tpNJLY/dn18Dn+V82v4z4EVICiAVYwF
Wx1JJY0YSKd8FYy5gojzLzPAacuk1nNRibM/AqxPR3xeiFi8ghX8yyd3IWr4dzIl
vBrv+l6kByEnU3H+qYHj2brc1LCqjLCUdmDjbtAWVRI+iMOJ+9vcscDoDm0xRLNF
oDCAE8+o1EmEptQcWdUcuS8vpYIqcx5WaZzs3Sps+l8nlHN5hbOBr+e4Ou0hhknr
IEWeHTogkI58b8qORE35UrMArq/9ChYZdpe/G0BUqzNACZCj5qIhc94Ik+QYvI2V
8kc7HIJJAppNopgYV79KTOiM6OcWhK07G/Sjsr2b8GK3mO8A/ze44kOyDw3Oyjq4
krC17Z5+6T3J322+Dn17pTm3+sGK17xVfHFAsXW/qEBPq4pPi0PFQ1oJhJwjX13t
9pizY+jLmjFoGnlgAb5r3FOj31HUGBIHkVTyH752VwOJV/FUA3OMlS4CL7l/vxwM
RASh3v0AKkjki+O8RHFsuVdMT/tChOpbh2QYxPsYgCfiFKpWRLBj9wdes1fB2TJD
uQyLMny2UZRJ1HinnLXssEabJJbzDJrH2tg0ekLcra9lBOfvyTEsApu2DIhcMdRr
3M1UuMkN6wBGp0rJa+7Da3tsPBqU7zCi+4N8UZNb/yvbHQLgXBrABARC4AqMq2cK
T25UcT4G3orp0O5Z3rP/xKs59suFnul4zCnCImsR+RrWPWhqhyDX4fYaktjC5A+K
CJDJ19/oIU8HZVEmPdQn6jdVgiKdf/JzKWdwIlJ7G8qtTWLkKyv9UZEvk74IxJSa
xb1Ppo41jLhRHb1vD7+hW22iPx6LDzUo1Z69NEqjvCIWuhnbm1WDfZUl87RsxQim
GVPPUskbxK0l+qqdmfhkwpNe7qc7ClTez9nmFMRbh7drc5DQyt9AV7IRlYBWkT06
aqLYE6KbKNvXwtQTE34tAiMUdpJGPzGs74w3FLaYQEc/k85mOAfTxhnr8NlYTj/0
98C2/NYZJvMxCzFCWOYeXKY1A9BMu23a2Ui/nj9mBdrDLeptSrXT+i6i2guztlLJ
HaV7NeFOuDQqIi9ke+vWeiHcd4U8HR/vvNVg0XU1xzIVIfruiw6GVm7F5ziFHBuy
OmDpgJnH/x/EuNo/fPqDLsl0lro8fJr/fInI9aSdG3/Qwp7SX4wHOdfzWjQwG3BC
6CM/777kfoDvWvuum6WDvRcrz1JzhOU2VSnllbJXmZXQoClUyEGPesFgIezhL+Hx
jAILVJ0wWSsCq1tP5RggsfrCdbu2g0T3ggdu7PkIYuuX6O07EsxM/XJxzBy3LWLG
wvhZJ0Z4J6XgjUJR7RukRGGH7jRUmWM+mbTdTeLe2eMfZwsyc5gbbSx12PGsnCuh
XDmGrzzm6UUz51IfozWohxdKjK1nW1Jq8SQ6k2WCBVeD6CvELNAPEn+FMh2sivPj
35wCmVByeRV6S7h5nItAFG4neqMkkKOF1Lqe4zZqKz5rky6KYmkGxpDNweTTf13n
S/psH36SJIEIuPgj134cJ2GGcCIUmWD9ckm2BPgASJG8zpVrZHfodvvNR/YO4r8b
mLV/S7Sbk4fy7EbX+nhdTPcEeIIFF4PYiRl15+nP6OauaTxrqGtFBZBuE5Wejwg/
88iRcChvLdL28fJT0k+t6sFHYeLfKs9Pk+Xl0lZULxw39oBz/VSw7pMMveaG4q1b
POO+632Eh3NKA/kdkBnonBcoRGBsoc7/kMW5Ce2dxgJTfSfkh3bpLeFHECI6LOHZ
0Y2YLtSvaqr9orQGEMdUsp0Ggj/aq1g5Mqx0tespj/Cdg/g0m8Os+s2pRVrDgcfh
wQdEdn8ZqdO5LddEhYs2X0uqSnebW7uWFExV1GdkO3q+qU0Fwzv7rnnYO0n3WSWO
57vD+0e9GeK0MShyfIvPCOel+ah5caE6C63ybbfxFfiPa57nRg0i6ob6NMEf4RFk
8E6R9q6/XWJ8EYUKTQRwwIseYocc0IAPrnd9T/WYNdEUX7F0kIRTvdOFyTs3aYtB
Mv5I2oiWjDkOQfgcX8Y4n/Lk8zahqr0N3Al51Q53BycRsnlGv2W0nYKU3gQ58zew
mmeFAR0al2BfetjXvvMuGTZgmq3lVQyQHCOZLY4O7t7C7SW96VHgBdt/d8ivZhGN
Igm/RWFysuPeH8Ha28Fz72nsveGNHyM+lz8o7bQTMxzpXZN/SRZEUPLulS10ZFaI
47M0bow0S2gzOwEfIZ2L4xCkKRnT0SyJSpoNmBkWcCj3lAvdwRSeumdRvQGVt1re
psSQuU9DAK3+222isqtYbte595yIWnnCQZ7AvcKMXqtb9ucX0YNehnQ5A7n/lOau
i8PbnbgUZY3/CBczdS68xBy4tDk+3Y0o8Uck3LG4Ax273spZAVqCtTXYvxfhXbpb
5rrTGM6MuOPerXICQG1X7VJ4ogBCyCUOt20UOg3hQiior5wlmgi/VZFPlXDsl3zA
dFEL43whNwGQeGoPO+IzxAO2Ynisg8GooiFF83LbqbQ3ntCGsT76/J0zkLMjjB2t
hFbep+VtOPTnxAZb2/34USsMcqyuhGmkvQO4B+QKmsi4CidpNyfz7IXQHdTYLnhw
dI8H6irGK2Xgw0qWgchPhF7Y0TFnwTjgmQwhQIsHeGEi2bO244cMbouyXMO3g81w
uw77bUBRp+aDMw9Ptd8Uq06c1vMJn1KNPT1oxPcED9/paUUratYdqo+th3FlmQax
Pop2h5Fo7MqWBpjidmnjcar2DfP0U39J+bLpSwt9+iC8QpeGSISOSSCRc5KQuLvi
erCZTExs7DxVPQzy/1GrYVjcKmiQqCm41JJo8ChfnWPzj7AH2VnUDeDIm2gPDP4S
pgE5/bQKFHIAI3POG29qnt5YcKmZLDXrsDb7rYTaJgimMOmV85VxsQUexNLRtssV
TWbpjQpJGSmyAgM00apWBLyve3NXGm6Lb6yFiUi2OQDugNf2RVyLucoTKHOYv+lR
4L892+CA1uV0oaLNUYYW6tCDC6kOMzM6OV/VOxxKq/xX1Q8hQMSpQudEHbdWQG9A
P9jZ2SOfIj69E+w7MrrhNOmAxQJkXm4JHpuf4vJG2abxVcpkqCPqv7kzAi5D2bJO
qr8vhlS52bLzyvVzlMc7xETMsxhj9O3GDJlSwYo6ubq8wwkgY80fYFJVnW+ZFGZW
liz/ModnmFBcGdjMgar3L27BsgEA3zEzz5DQqXWz+gBjlyPqt1yx42bFwHPlw3A3
t8dvh5BbaL2qQ11iTfn0DO1/fjjdpvWPX88+v/+JbmnYgnPVPY715B5yOS4ngMfK
82Bc89Mkxe4aZP/SoK2dbc44uffFkUaPPjv2PRqqAlW7jqFjWU7XtUCTnzURmbWK
0ZxSol7mnRKOFyrAjqBgxQqEwIvyHrxvsasFGynTTZHauhPC/nVaGDZQno496E5p
8aAvlFrRwU0LBihfeiIxQLjlGWJp8IqG+/pvbjEVlNUmLpnPH50An0vuV4RxxJJK
sSeN0TW5QYP3gLyXhymW54KNrjAKf1I+FP94dvMwrfbjYQ6YJmf3mCWMZCa1zL9h
DR3gF6tavi5ntjfQ/ac61Z4L84vu7R7oWHlXLtPBc9uhvnc3B/DIQVBAFoKv8D+c
1lRCuHSCxvFMGqz+uzwHLTrWdLiVOu6mm4SNuZL9ceCT4BzkGSMvqiEW21IzF+kb
CcG3DhdOthBbsUX5aCvsTj8vJGQtbhJnPGD/YM9IGNz2c2cxqbnLa6tnmGWFa2vC
uLzG3GBzX8hwxbReTAjqDrt30q8muQN2Tah6/OgjBvwdPZjQAFUY6ktNGYK4M6pE
0AFe/IKsKsOF8Y2tF1fWM3Ep1MHvFoHq/LrIPonIeWnAJWqoV2tAjSfZ0c70erZH
GQa8wh83k2YrMY/NyefR9UckBdTr88Vc3cBn1k5CS1yNlwhFwWLHtMfTYQkVapNh
RYkM8grTVsySG+NQQ1muh1WIsrfOtaSgQ/mIwwbNcUEJHeIw2sQGC2yXcJu6hMhb
qcfaiFPne14re0NGwkYmJKlDk5I3zYQ2pjWlOxZVDt1CcmFDP23/gj4EOM1vq9E0
5HG/nowtaEumVo5yQNF06PoxbjMDxjEC+BYx3L8M0B0V39wmezA66jwz6alfuT1Z
PQWs7gV9osmPtT/H3fiACOx3c96KpwAMLMBWoNtcrSMTuBfa65oudfEP5uF0Yxjn
VI1iJA/znLFRGIEbpzzHwR84IB0WMtjEn/9pUjzycex75726tJfkhgSizj8DCOAg
B9oyNNeCKZoMI/9u770rBRvpcFHpS5rEahe+k49Y8rO0pAfJtXWrq9jMWbv0+8ZI
BlIUXRYFnny1kYE2ev2Ebjcmp+H4Xk1Ugknu0YWIz5wlFFPIi5+yIf11IyXTB4yG
f0FYDTUQCrudLABDHbnBxhr6e41h9Pw28x3HlZ3dyNFKq3igbbg+BYNQssmJLXqD
PAay03SnR3wnIL99v1R/6Kpo4bMrdstBSSvnuvaUxr2XoQ+otK5Nzbuw7ThvboQT
XQI+PvhykWxmrc4LOcDQ4nMtYahd3bsnpD2YDxIhWUVBAURirKcl+wyRYQ8sIgfm
nbJ/u8G3tK3JNH+zUU2pTGPba8Z6sjDI0t9jQPXAGYd/VmAiE2ohA6eJnukQw4KS
tDpNQ2GD4YDRxDoC9BQ306bHGeTIxVnWWJ7D5vKzt0Go3tLrHwwyCFI2H//oOitq
/4iXi0GlD8cY2eQ8sWIUhRw8u0gxmB06+aj8GEc7qaxUzd3B8R6TmDq958eUU7+V
oUzBwqIj7DocxbmliYRod6+WHaiU8vp7MpMN2rU2gFk/d1I84WwWJSrggulmxUvf
eOshUTkf0nc03V+e0im4Vo1UzZS6y415MNww4nEz3VCLiiUSTAKkLHYzamfoG/7Z
TZhCs34noYc1MtOYRjeiQarRASOPWMAeA6nOYCgz4LJOyP5EH1UWsJ6Epf1WeNOn
+Gbo7qRSJ0CPv+72prbrcdEj7q3FUJ/Wpo2JnwX7np5o3lKynK5cJD7mnuRIPk3K
aXp4D33kohoWOXzVg+aFtLfEq/eNiGM0UYJPm8U8+aAgAJ9ZKJU4yuua3bB6RsJr
HwyY606EbIHYnLYBLD189MJi+da7CF/D5zruEA0zigjBiuwJGTfkCXejWbRjadnK
KaP9VD5V+xfpiYDsnQUESlm2+Wahuvt9BgPk2Ih4V32lAJceDW373GBjmIeV4hI7
iMUZUT93GRLcuywUe27lQJFduuvapTNXM6fUKI+d99nH5p/2gQK6nPMzxM6S5veL
Ete2u2eQIS5KsjlvqD49VI7O4ALgLUbixFCjsuOJbQy6IOEr5N8mX1hKPUphSKxU
H+6Q0ff8LoTqQJFcBc6Q2de5wAgg4FNa8CaX4+YKKtxC0BC5QYZY3Tr+EcfAtZSV
j566Fwhu05JC9fa171Rcj3uPAgXiBzKllEnzGnwlyIcbsjfI1kF80a45/NUEi/Mv
zxuXGfWjVLmxXN/uW9daT2BuKCuZo3/mO2zsD3uxKvOOaYsfctNwL53IgTt2+CEQ
Gq4d47MoH2qxFMNSisTbh6821ukv0RWsC81V4WXywvcefyG53zIFpsFKxa3kmbl7
gLxb70iSELI0TAdMt2NMY231d9pI6Tq9gXlcnJouL+nHEb1HvRJ1eU8O6LQ/jfv9
q1NC/Q6oLbHgK8vLwzT4fB+KV0KK05OC4KdJlkTf9lvIiKUOlv1AAVZgKqiAchhx
WrPAEATsIVnZZ0PzdIcu5DbQD62o5QfTFqRl1UE41Bo7+TQXpiEjJ4iTjn6f5PV0
xqTR+hn/9Koo7ZMxtI1qyZR7Vg5HdGLucuyabELJiLBUTqrDyC14NEla0IvsR0FZ
GkKkQ0l/UR+POIvQ/BqYb/nhnn5u0e2F2E/pRVqsG+Ss3hftDtWldCkdBwHQTXLF
a25Nb4tFkJuFeRS0v2c5yqlM0NI0Eon99RJ7mxk+KPtKWvMYSmQw2jBz+k85OUP6
yrFOzSO9BHblxaaLXO8h2Iovz77xJKMozORL7vSRjADmqozn/TgXENw3sCNN/e9x
ForB1lSzAgjY9OdTCBof9QUiVV6FbkmihsSKxOr+TafTRau9NmV2dTIBzshAkN71
xotSvEZzhirZnODBSym/5qSPzCwuDjKrgOjLosztFNxTq7k6pz+uYPVh2voojFit
atwF4c2PzSwhCbFGXF686JJPSJljsadc0RoGIfX5H2fDNpOhQf4hVKNnUyExcSn0
+gjfKsIPuPMuBudG8SpIKqTR4YCPrmpfBaRS0uQF7uH7ZOLA7+Lz+1+FozGCaCF5
rZNDYq4Ez229ZWi68S4lL4zH1HXA8FJzuvK+zMF7/eHY12LUSK3kbRY6LWvqb3Bn
dC4sntb8m2pPB6exYd5dzacJRBkKTqbi8+v14Awttt6EXIqJ70bLasNgmzVsNbqN
604heluMgdNhJepoQI5tcbfRUJw+iJzkNetLgwGZ1nPq9eQw8YLMgpYrScRgxaga
C9aa7QugdkCh/b05K7Aa5kVP3L8GISnvm8DYjvf2kRkGk5Jk7WkrSaO4SZRFuOKL
ZyizP+iT6iKRhmSy2HydyEV9oZlOSZXMRkiEtNux20wlJBmBDzqh6aibCFq4ZB0l
3fMIMtYOLBKxlZ2xYDD1Ziga9ZTDzxlCSYDHKOf2mtcQelXshees16i/qcEj8Js7
/aHnDmdRNWhJtiAuytogrOmWLWRRpkVtoRYnB7kinsOSAjlsBfbqF7ECGhohW8yK
1yJRzfHjenyaLqT4/WBc1FJzgtq4XSmt1iSRpo/m/4Y8N2hhi5H7djgZhyep68AU
zO2GXOBLuTc8re++24r13miBMQX6ERNJlVCWDmHs8/2ittekD+Wr0YoWRMC5onS8
YxmZMNc9sdOe09XahkYj6DVuCFDBom3/I28VrdVyuktWeW1nmhCktXw8sE5yL/dz
Hxj13n1l++JRTOpNGJJH0R9F7ZXazLp9FTf5mKzZt96GtXqiFgepkFybIBbzRxrY
HbnC79HPmReMJXVv7Nt0rxaHRKYcHHrYlwVHd6QFYL0Y18zwyOknfKsHOD2PAsXN
/7DqA8mVqDmvHNrLdrOCD9e3OiakgJjoA8/ddojfAJNrRq5CW+DqPZsCHpQCAuZx
nhHNEDrVHQfiFjG9asbh52SRoGyn+dioxSOdqz1sIxicV2UWSoSuBmNji5vspzZG
XsFEGVjnksnykkTXJWvWQXsJK4ZyKiZ8cmDDbgM8J4zsJH2EtARSQ+GfQjbUFfk6
y3EmaRasYTMaDpnebvdJQtMloij4t4bBd+zfAbs4jBmzpX9MqydN77TKVtN/niI3
9e+bkdUhLvLQbO9FigSyDdEWzZ8eqK4W+qGoc5XgAoWu1QeCjr0xxL/oqG5W2WO9
ClkJT8BhcA2M8zhQJU8q/t5BM4wT/4U7eiGbVnOVwJ9KgxxSS//ONUYzOnr7RWbL
d+JYvSrvm7lYSn+JFePugIFnFlvn0lGh2WOl+oc38coa42QCI2Ea3fj5hUiFd4Dl
Tj9FbYQL1TAmggi9SMNHmo+ysRI7co89IOp9eHGClE4O3VOw7tD860PiipXjfR89
8tdyXzNAAdc1fInGjOjtZtRA6z9SOTG2tSAbujCwWHlmK3ek2Nxw1Q9EkP/50XQM
iWWKf7CeEEf78ONinWaoT7y0azeJggVw8+Xbyjhic8DcO7IzyJWo3rUT37nu8blh
8HN8/qs1LaStttWksJNLVE4z78voHeMGfFn1hIBLkPxIrNOE+Xjg2Nc4+Aj2WMTG
G7wtjx1DXvScflJcRWVfk4D9b9V8DYaNo8hBnVVpdxEqlOIQYViYZkPyxsD8CK2k
ANGfgz1gO/hhkj1JuqePLB3Makk6EGyhTboXoH5jFZX3UV2YLCKrNrmIjkTWk33H
S2tSUCyCQJImj9pn+DIYWazLEwWOC1ErsOn53sQGy3/hu2drTW8NWbWdsBFQ91mO
JDPhhyZUg3wOU0JtfZfwFmyrR+GjQQgbH5XsF6kczL2R6+U0Dc14KTPN0+6jB3zI
3fXUqyXnLQbxLALmuk1XfQ0Olk406fG2OuSo/GUo+xtPNsl7+xckSlggVwjrM0D7
tEdN18cGoJUWndIm5053oi343ELFGuEsNKrvU+RvZo3kt3RuuGu5PFtAFc9Orfol
4fkRcqK1QDBphYwHwIV3jwZq8mPAblqp6Ye8uxSANY3fFd4Qk5S1e/JfqtJF2JaC
1bXVponFokyWWSyJFGtTsgw1L2VxRLg2EhSUtO1z6DIn893ETEjWLKbbQgtN9b6w
wNfuJd8wj+S8ebESjlAKk1rAxqbxMeJrRWX+ZwlCB+kUrrX7nHQEpniqZmBVJevq
KGUSERxCyrUS1ekhvwcQMLhJ6w05du3KAYP2H78xtU+iavj52P+P7VnZoCd0CAbo
ktS8B00R+IxK3dCtyWSo32r+l34fcfiVUuGsyMB1mEvbhkXOl5KchnoL7Tey6DOL
iCcV6BreG3ZHKoGpgGADJT81fxuKCDuzx1xGg/bpYSiv23R9BzQeGU3uMm4Z/dkH
8EIeyxyYUP8jiqkoWgUJld5v2UXM6EqkUHswGNcQT+exi/+DN7vC5WjoajNaB2YF
lzI9XoaYYh66Jn9FAUUl6AFwDfC7MaBuO2BCx9+ElhkMrPpystFMPfrUJln8XBQI
Hco9+aZw44HFRs8PZjQMnoPdGVm5ealbe0paAms4C+2Ml96wTIZdyBEqp+PYmBc2
wMxHoWE/2ovcB9EX8FLQgzb8iN6vrcuMBW9MyEf79pAktwQbh16gO91aEyVEnMHJ
8YjDOrkPb31sbrPVJiUY5I8u9RtjkiGado0PVqPY10BFs1iUsAE6QSwwxk6p42uY
djCOuyDGU2V9KMIaHHMTWvmRLiVb4wjRP5ww9DZ8DtOlwTty11C+tDlW/KhI1Fpq
gbtUixd33js35tZZ8t6dAeO7iLFTrHrVc3SgNNvprDGCT6MbnknQdTboBE5GcWZM
G/3OwMJ3S5KibzmmaS77QZmsj1g5XIShr0ob4NuFAauDHXOw5HUPG0Px0DED1cmn
lL43hroug8uULgaJPJhA//X9M2FDqiAYaEfyxA9U7C+p5VuMPkfjHm74RN8MN9Ic
KcyZsGb0iT0ylXds4FS6ZGNFa3ncwRLK2CRnT8Pg1Es69xdMeyEBqe83u2RJmot+
yEK+Gr/Ew75kN7kvzbOyshY6AymJwMgmISxcRnFo/SY/03QdRuyZS2u/zCtr/w5C
SXPgViXwTmVE5OszBSPsEqMYOEIcLTzhclZfJorgBq1Zr6aJHyXD4nKTE0zi17FM
DQZrdpOQ5TnoWK2I69hWN85hXWSAxy0Bxn6dqWgP1ZAGWGFzYzWJuzoT8UVUsTyS
nZzwL/UekZbEA+Qs2XbBAFnhzrJsSULwAse5IRVCVkrnTXLqcBhuDbAKNBl5qC/I
1mADM6WPLwxtR0Ew0LKDmJ1DJPB6oEwv4VmbMyCmcj23WtZmCfUb55DVloQZJNBT
83pk97dfs09CK4XugX2YJWhyJJ6qTdQ+sPFSIkYv9ThYjjqfodL/mCUYz3dV3+ra
w5fauJ/tac60vg4Qq30bbu70syZBU5I20q9OT1+/8rxJLyM+aObcpceJT06i3Scl
xGmwylTN/qB5nFBH547P+UWuARNs9WkhBp/IfnlesYa/qGzJe+HErzctATfTzZ+h
bl29+YZ5XSCvf5nT13MVWcmr8qfkbqexxeQxz1i6BtDTPvCulvEDdinLYvhkc99N
LaN2MLPrcpV67cB7Kpcv/j7Kxa+sexVeoTH78/MWsnPaY1yICWGDYfjF8cRykrcL
h3f361c94Vhui6muBztVsjMEgV0cdNWq/Wx9Ye+7kVKEuiTTHOC28q0+igW86yQ3
/D0XSCrBbZfWQi1yEp6f4f04D5nZJYBObJrOIfHQ+dGU5nAXhq5DudhYSwYwcVk1
v2o/3XmprKOg8Nq0GPU8jWaqnd/KykdaRagCYYRiQqlJmFD+6CdfCtYrfoxvz+LC
rbOHNdQ/liTbVkfYcouahLWD5yjm7vnIZ02SxQx10sUpO8NAzYC9GMAMHgh79ioN
WxNys0QsoYxu0w2xX4Va0fzb7/T6OPBj1bEPxyND+lDHFUr6SlP5DoXTRSv9vamM
6vwJcRHU5CDdHbkkd4iEb0nir9DhY4ax9pFrN1EjmMZONHTEK5Ar1L6IWhRSPtsa
ZbQ2zyj2UR0bBBR+Gz0HoZ3fPpaZa+WmgbZ/wP2QuSrFTAZpQ5dMAeCsCiM0XlZ/
18Q5B0gu4JFLSDzjJK659RDXDLLqkShXr1JhJH0ES2OwpsARFHJVXMPErMlk0Bwm
thl0ZuLPDPZDyUsJJSiOB5cStchgrDuvPDEy/AcZQUHkiLB+5RTVMmk3Uo1IOpDD
D84rZLeLiTBtNZgOL0Q3aCqnI5lTqcFm4jHckNC7a5Gs6mwjoIhnCHh6CIdzn44R
JQvfbBdM9Zvjuo5h0/jzeUkTF8tyohAhxLIO0jvloIs7Km11GmAyaWkDX715ZbdQ
/7D4kN3ENkXGqJ4neBOslV7GZv6jbvs6QHg8K1clkYfa0Qwnl38qE9JT0t88qjfa
XwnZOetorr5roknFy/EuxGz08hLEAMGRsI0D/+/lrg8M9oVRevNOBxvFgvSDdNUP
/WtQktqHfGXDPMYcEUyzSGIPcbU946MC7GNADvaIrfXgtfcTeRzt71FKVqIZ5eeM
HRygE2D3XyxpK5vsM66NspHpba0u5IxiZrUfu14atVwWHwYqWbMIz1ww0jOIS+Pd
EVTgak3XxWoU32u3VXr6DN4SHMOz/kHGx3jqgM/m7a1PAN33NBD2iU2KnYN/l3bF
HgAILpz8XMU/vRP32Yzsfg0M25iDLoaLxuxvMuUTv+23ts2Qn6FrchYWv5k4XRwn
LrOTVdkwPhFg8Hjhv+4p2GXu7TjeoHxGNgygNMJfbA2TwDI9jomuaGH6e0YXVEIH
+zYXiRTo/KM5AkxCJwj29cXoKz9SAh85r+JFDnhIGscIokaGDfQtoSwAQDDWIXVn
RtOLWql/irYpjbD5HLfHGqZtFzAZSMoqFBK27KC610o/qYEdVogWCN+aZKNjhsGt
27jRa2/r5uQG5ZgejanPcYyh7ZRikLTliVrM9axhQ0hmbNCK0cLjz0a0yCuJOX+G
kcoJRFt5kEmcLf/aOFbK7ZmqkjauYkjVDpajxBAvNS3JhdU6ed1RXheOIUcqxZb7
Jvy0cwP6gXyGIJWUuYMn0fpQYPQrA7AjqKSDmsb26guVQeazQ103n7FAqttNoxaq
JRciAJ2XHD0OgtBICKrTnph3h9V/fPGS+FjfTLDjbVJxrSvGlbtj+h5ZBU/9qerw
eTqGgpBK3MHKZ5qHLI6cpA1EOEz2yVGkjwQ9rwXqHvOzYQXOs65c1Z339L1dybFs
pMLddnLT684ANmEs20YY4ItdzerNvTOkemT3I5qIiMJqXXAgwBnN5X+BkbhRjhPA
NqirVaIdVo2pv5KlYuRv7J9mQ11lFSSdnREPWek3BJVqGDBlhJyu0jn4+3yQm6E4
y3Ces7n4F/DBlygpduVV+q4Dj0DVzon9ibhJnC10ZxxA+UAKLWJcYsPIUQkF/Y6F
CVOWDR5LURCrsiGXavfZDskePEtdQ+GjGry0M7rKZ7YyzMeKIL32sIbz+AAd3pOt
SPWGRC4DxhEOILyDEBoRRRnAnBAP6AO91PLKObTzMhcvc4VHl2Cz6xW8K43QNlBR
hI08B+5r93GlUBSL5Tv8+mC/C6ZUzOl/OljErM/lG2qbv9PmH9CeXpFQJ0iohKJO
7helM6UgNBMlpcCC3MSttlhexlVBf/RZ9D/3SOxXWgRXW4VH4uXe5E1iyMrtDbeg
IAI671YuCOhMJrJgyTHTSob/01UaeernDa5DnRnfxHU5N8drEd55T1o6kW6wGF2j
zwe8dErWgtN7RmjdvxyRD2t5B0NLfaU+O1pRkIf8ellz3mluhZcqOOOLWvFCLNIm
EAZuDBzvVobAen8dRKe5GtSJ5sGxt3VFpVPeiP7e4GaZbLIueJNMEbQMiWX7bbu0
So7F4Ii3iET3kqUr6Xk9yiqUsV92UzP+/QlcWjKLy083XKdbNbfB27u6U0TPpqcN
ghHE7U1UnEK3FsmYjU2qflgf2/ytyrJ2/D5t+AzeAL959eE2JmrjNI7XvuyeyeQx
DJFQX0yvzG66aXH0fk/vAkOi7ynsr7y6TpoYzvIVE+wfMBiDOwvZiZub0mpUhNwt
YJ4y+a6fuFyeHiqZ8PKDf+uMtbTEN5zrHxXNKwUfcDIF5Xf24PXuURvTRL3vFheM
57tuQSuTKDzWrNfIhcU5hU4QdpvBM30PUJCbFAPNU/Fk8Nvw7opj3NEkPjm6+ShD
GdPsqAXKCQZ14TJ3sWYMqPQ8h+RllfzmTZ/TrAnCPACtj1MhnJHAI43xEB5aaWRD
V+JWu252iwJvpjAbYbh1H1BuP46vHwh+US+xiyp+u5pWanSDSygcscJ/Z45pyvqI
OiaSQBoYWAV2DiPORTnFlcN9N7b4RUnvtzaDVtrfG4tTVnwrObERio8Ce1Ou580H
zJ3OTrXf4VNqbEhI2V61shGL+Gr9Syj9SWQ+rs3NK6kpjKSLSwzIER2cRkiyqMx+
nW32fIX0xhkLfB+wJFMJJVVWgF8CTvQnuvmyjXFrn3D7smglkM/jK8DL+PaROXqv
Ud+PGWXRhsUI/1hRNmxF6g2XoYyuWhOYn0asmc0fApGGjbaFYqkMd7l2funZsDyD
qM8cuvBjB/lzXXMHyWAkjRomJD3cNMcN4hZQPqUJd6YwsJFSI2/VI15XdeSWK5SU
PuQdGDR+H8X4Jb5tSEoQGrm3+h6vHHdE1yiWA8JHxUF+RJhTCFypRJaCgVupijbY
ZI/zg3maT4tx3KvX1E6Q91EN3HTfH7LHwhPiVtKrkSOfI4zhw9G+UdnRKy6hvZQh
j5LtkVJlUbp1irPMG6H/Y62i2C91MFE+9QNzeNjPlMTYt4Cp57nQ8jYJ9ueoH4uu
ZSdCejud9eUWTzDGKB+o+215ciR+NDE8uBUB/NOp3qq7RG+VEMpk/t7PwpBbm+4x
DWU7jNM/q1d8iitlKjPIr/1YB3t6gujAAG2jy2aqZ5kyocu0hdYvIIuSGcoXfaq6
uG9aKdDp6gohocOrXQywzjKLEvbYZqXemONIGcUvVozCl6EE/K61pntkvlhzRJZ6
pv2D4x3B6xF1U86sA61pT9oVGAXV9KZJlXrdxtfQCm4oknsPZAEoZ3XLn4VxEaIp
/RNc/JJLHagvnRw8o4jBwXVPpcKy6eFlMhCDEloOkgUBS0XGGIzXDWnNkJI/keFZ
I6RzhOtW6mEwHWx0E3gfwNrpDTKErErgWuUz0oD1RVhnKHdme+xf0g/s3EKm/j0A
nKOl5B+pPyfzJhfwWDdUCAxDmeYG8qweWquzrinf6lkZtbXiEniwo6Op2AbrfFem
rzJSgPhxd/w/p9Sbw9uRfS6ng4V02LCGjEG39oyfRLUV0YUQsu++JWeb8RNTph0o
VOmb8DlMtFAdxOnC12xtVhP+dhHfZB2W06P2TKjnF0CVKb2Pr4XcrFK1Nlmrn/VK
pg4V0G/0sRm/9nIhgk4lbqcuhGsk2bZ3nXHHC7VXx8sP76E/+pcnaKfHFISpgOpf
fosPXlNe598WX5oknSm3GZSSNx9HZooF3wVKumCYslmyNxT+yvp9c1xhcUI1EqaE
dLtUcSstAkicjQO5ww6dPPXPmTkmRfnXDjfMlg0dLFfFDA9/RK7uv2g0QwNl4StN
ryvV1xbTYz8M7LcxDOGGcp8eq5C9AxQ0jjOJWN0EbOq3by38vwC7IsyXfrus+vz8
8XRbnCHBK9ahN3L7q7N6RgHwCR4gAfZUlGO6FyzaiqbmhG/VV/xxN9qel4EvBcf0
qa3W7V3/vMOvmf+FvkGH1/o5F7gLaUV4aOVS2pxphrqYCphWxvBFcG2SZQIdrFtU
Zr45P9Ejqf/099bxsbsYToQJzGDyjTShgoPWFsdJOroMYHgTuh1uNCWePtqReHmG
Br3YwCI/mIgD/R0OY+HhuvpTS49zHl9cVR2c0ULTCqpQ1lVjJiB4ZGXmhHcqL1iB
+uqlKCY1cMPdGLVYshJuXRBYlu0xcw+8S6GNXBsZKPn9X9Im1aYz+289F0Cg6Mza
JwMKcrQn5YyHNyogdnEB7JH/wd5D7v85UFEZtqq1KOlj+9taneDhdgU03RJ5HXBg
5AKj7ODvfZEsopyU7ce+GGC+KONIw3FWP84JCQnmlaap6kdcfNKcLmxBPFuXpJS0
ws1ya71DUrBfR3FYT5A3LLskotVKUmgAF8VxNSjD1etnyHrpO4qS5gseBe8bbXcr
6RhoY+tWKbQWdKUlTlgwaLnZR07pbmjNdzyTp91uxJYjlF4qgKE5qN+ot6UhQqoo
NuMhqEEyaIR3baqTGwy++bRSEUMFQYVU6KTPE1u1vJlSqARMTofnOb88S06zyUxW
o236PwXOWmteU3t922mhHoCByhW0Zfblfsvf6Kq+0oEi/nzJwsg2hzwnHUn8HF7I
K+r/rVl1uGlLBa8MH2t36ib9aYQ3RBC8TqylCBnki2W+g6j/AdU10cY2utMPLgC9
8VEobWHGB4rCUX4Xwkbb8w2HK5huPRknXDSEP564HTGdPfprvR8tjk97h5aRp6ou
8rzDLRfoYX2eX7k+ln1BGZabgbyDFKir3wxKuruQhc08bFrgeU6oRu9W5bkiYLqR
ZCt4GiTfP7/5eFiYaAYLp6aEbm1Wo68uE0iseeHE/uOymQfjyc0WM45jIQnH26+i
hLN6gvXF1iRz1B/ADHzI7A2zKum+1SFeoos6eKQYuMhbduBc1Rs1yYXN8PUP3HM9
qcuIPlyHrExWNf3kfsJ6uaAUU8kpBka6PGiQ3cpfPH5KZIpdhffvPHbaILObnAI8
G1gs/PjuIkyktMXu4djw42PjVTZd51mWT7gkKSUKpwECcRRmQV10MNLKA+utFTSV
kJQqbybZl7jaihwDVeU2JEf7HO9UptVm4Ph770bLc7IEoDmxScwI4Q2n2UVnMD1/
/vY/3RtM1b4qOLZTPQ4y4qTD3Ues07/cXlBaDEATue2E4X9LDkKkAj+jB4oI1CrX
knnLNiJjz8vj56H1374+vyxYZyxX+FTc0URAy7j1Hos5LhQYmXHzizrL8pj2k90n
5KRBlU2JpLqpROlVRYPaxQDWHoy2S8o7GfYdjg44Y9yEtmJJlbOQJSJLzmTlhFIv
LefkJNmHv6YhGvQFLJruGCw1R8pgCopEGwCCuIaatcOOS73lnzOnZtOiaMBlLLvi
mRIteikijrLmpaxRjwKPJHK/sh7WVuTAK/9AQz9Sc5xDzrx/FaK3COGX6B+T337t
WnHFbxMOALzuYQzh7sQL0oH1ydiXg15II+3drMKFh/gqmh8MWb9srSSd5T5Pdkzj
SE5e320LtBcO1IZe0hsoRfdhTTgbC0erXvE9+LABj+YFp6hNIQvaSPrVFScrChDr
9JFwVzW8E3mhP8JKvB0VAdE0/3bsl8YxMjIwLr5R+Knw9MeP1hWNLywL57WNFTzz
ZNnAgZrJdT5uqvmt9VNuzfD0wref0jtn4f71NAEBmdXjafTwFSP8nyT56fjHBT0l
70HEpGrx6b33n3wcGGoC1ZG+7ZSCWtKL9pkpNvhlKx+lkQuJWJ9z3RVcUVD5TQMO
i0gUQvbBl6klKTWB754YrhGhKqZ3lk+F2kFZam8f+XwRP61ds2GbuR4y2c3AyFqB
RjD47xr4KOwAKFiJj1LuMDjpkpS68oqCHUTM+oaAza2rYW83CrJYkKhAW19s3Bhb
Yh5HzbZKXumLNzXCE2X4fqPVL8/iYOLioT5JSGutOA5z+0ZuaXasijjkBpp2lmfm
kjwktZeh9b3iqDz+OHnV/eFzHEd6mh6UkVLZb2sxzG33OczJ8CYJInJeKZXv6pMF
5WtHPviDNmjiai5ZP74d73Zmk0IwFDHuNvtAfhepJwacMAlHEdI510pvIog4R9F4
oy5T/DEsYqPLgteEPeyTViuoBn4hcnuMAHHLCq5h3UGZyhrnoWnCQiekZVsZn3zS
5q1uveh6w7Lh1tgGktpAFq2IshqR3eU30tFFFBZFo7qZETkeoWMFHicXnjgljZGc
AXZeDm1TnuR/6uj2zznQ1lLLGDKLd4czPzwlION7E/+zYHTDBTh90WRuPsU4t0S/
9d2dQv9FH5qf1qs7f45nyW2/N0oO50u0JLrVTvJ9hEFhqPi4xNrk24F2bUA7clOR
iZ9/1TPT4yaW/WT/ZYrgyPOjckt0h8uwHDpRWsl97IdkBKuyH3d5cADyrryF4VvI
1wMgiELYA9wiKKZ/4vGX0oNUt8+dDEqkKdvP7einkWrAxikHHz6YaRdgBg8nCyXt
YWdY+XGC2F9JNfVa1vmynbLVmzBtKCCBW5Vojifo1qGEGJZI3miWFh3KIHAmcy0D
nLWKgR4bv5BUlYlrSE5GKKavnzkgONL1vrjrh71hRqXEg0O4mG5GMsZL/T2VLRYf
slI97gQe3qOwxvO4R703rImdlQmMFUND6BPRIBAtg/dlwV9Vy6opygcpDyXwbjJu
GPBPeoVfj5CCUWWIA5pPo1l3p1i3/RzQZnB7Dr60i+9cwIpjT/QvPYp0gjkEuTJc
hF2JpOf1v/Yt8SUToBycihoi7MPDiE39mHj7WUt0l5FWU0jWi9dmS2QpkTHloTwf
cNldlCIMK+5AHEdp2h2X5Dd/N9m1CWQzjo5ajG59JlKPK2fSa1TjGpauFzy/4GoB
6lybsOaMSFcgA4aTUL0gz60fuv29soRPPaUK4c1XW9CnXgzGDHMDqdd+9M2LJrZQ
9XV+gU3BIjE3j6v6uyHY2/y9JWC1mbu1H1ldpGQRRwGSVL2dZPaZ7VxRUlew43/q
3qmMa1iUEu3OgZD0bxS/mVYpwA+a1CMtCKkWXvsk2jhx35aVj5tIVxDjv8969MNR
RM3g1BHKAam4f0eNY2KNUT1AX1nLLRjufI3Gqyj5cgaJz8Vm/nJtdAGRmbeTXHx/
QU/o9b2ifgAt97oIMLYemQZA/dwOIumPVs+Jaw39a3eTuclI29oeNJwY6vG2R6BX
h6QZ6XER2zRsqmwqmFEeR42XvBzqQEjdV4opVTThD3fI/11h0rAshjVHrbD+0Sg2
/Ka4w17zawPwO/uIP2jFdMkt/g9dNJmr8T5f8YOjfuAuWRLnP2UjoCRzsqQttIOe
84y6N+9ZH5TvD8ntyjQfF031cQxfT0+WkJp8mstJGZIB0GQ8GL2VTbpfXaSKPHfC
yneBm+dbJMtBEThRbDQeOalQ6rq2aaMdar+fRcZ2qxRiJ6fPF2ogFpDhkidbLJRU
8Px2qGHiwG88tw26yMWktqFEzDxS6KSfo6jyhMJiWiJDZ+mp6XMqaT3Ly8b5vo1Z
bCsSAYQQCwOE66d7U9W93ynADq0r3BCk4s4nJFI8mwK+DXqiX5LBG/KN2eXXt8H4
YRS08YQfnc/ZTQJRBA5U3JT1P0bnADQXZCTgCwtog10bomPryzruW/7hD4FgrSQA
ek/A7RfQkVnMgIO3FCfLuPZCVKhmvO1kK/KVt6SJS6mBGO2nxF2LBWwz67n5P7Fd
I0V49Ei/LQI7uzxmmHw1lZV7hzcNIcFxAXswZP5d3cEqtr4ZkfskNDA0Up2vcZLE
7eTgmphDYPq9h65oRgbYB+QGoMprBEPkkMkPPKnC3vQyHk0TJZEYwmNh4CQpJGKk
bEfyUvhYOLKfux9iafe1OeoZLHoNahp2xIB7OsFwCsOR3TzutQtjRWa7nd2Obcoq
d2wz91/GIvngSzpwZZ4WdA5yllXZCHf8Ns8iw48hGClv5bQbmWyND5lOwcSjMK+n
ydtcpjsOsFT+Ox4OvZO5NC1HeYTOntLq06INx2Bx4h+W2cEld7Mx8rFxHjaBn7fd
Gf1aB+QEqRciQPyrvRN9/9iFVfipt+Afuc+2uDGabuDnjIw83RCIJ/d22bP4Bma+
mWBa4GIlfSXun1y7EapEQLn4MdXADDi57nfVWPg7WbULEYDd6DNAtJ9YHNGaEM1Y
ntkr+B33SjHYTEY75dLdcgVm85CioqipnSxksXQeIFH/2u835DPlgvpenMz5BsuG
r30gA2w3H9zKds8uiFafZISablqAbi3svdHygbPPpd28/MsZAC2jU0bqaqqokwPZ
AQmc4JtZObaB7NgsmGB1iym2XzV55acGOGoXQaehm7pKcXduzyhu1KAqiLO/S+Z8
7h4N25VsuuJ6D2bOqMsVFNpAp6RFGZYpBctBkgQhM7Ai+Sza8/BZrhXcpuF3HheN
Rlfta9qqpUBHztMQWDiePSTQ4srY6808vKqYys8ACmR1+oB2PuBgm/3n46uzuVob
gizKRMi4KP6E/48BVF7bvp0UccggbcUkAico+b7Tj1Oc774t30DeGwbyNAWBYywB
N1u+xyXFp3Ea5K0nfqEXYij1p4DU5vJNiw/n9XrpUWzMjfyieQPLGeFR+EdQ+onj
KIOXMQzSafftPdKROhTo8PHDzjHAJNLMBHLfJCPX8SYDJ6lXhsLd4HU36W9z+kJZ
xAgHZQ+lsC9hbJQnq+NWwAi3sQsXsZZvGZknRYZpBFXTg5HqWkYKs7OMKyEXsoxj
OeDYBcbDb+b/SjmFqMTZ3zbpucIB2HDuF8avJsL8xCdzErEJXojXvxxnmXR3H/1Y
cGgBQgz988VYTeKn92TgdaHdwNebDeNqgyLWheYU2bhLrQfbcRL4sTwvBWyOfSvD
cYEQXHFpda/LcxNU+A7jnV7ZGxr+yHJY8dnvRKlKkW+WYibj2mGdo9kfz4JRuRZT
/RmZtO7WnWngVl37EROvJushbSVhTsn5VzQoYfXo4IRnv1gK7LezM9EB1y/8V+fa
KYW/tbfGWUCFS7hraCUuwdpQqqDNySFTaHsTacow6eGh7PQ0Of1PLgrDSNY8vgup
t+Qjxk7tVhL+/+Xd+cwo9qJXTXi7wBpSUt9nlHJJ0hOGh95vOUmrBWIZPNvkgIS1
1pNlBgbw5wDyiBGz4H3sY+iBtvK3AE3VnNs/FhHzMfgi7+l48rj0Ikvs38+Xsjvm
uSNwU3OSytZSDHfUjitQOdIVRkLi8abSOZ/FLbB7u1h6d9N3GzGkKsFBjHhVpZs0
YIZ3w2y7CB9Rt3hbIi79Uz+dTQY8GuC6sgXFUEZ+QnHtBckLriS5H7R2wOBvYC5p
CwZihpr916L1Y061+OSnbLYfxcfyGOPLw1VI1RLlUXBTIXDiQZPN5c71LvuQEy7p
6TWREyQxEVggiaUS05h3YTDXzOiTLAotoztc/fcKDd9nWxA/6gCNza6zW/LdTy1y
07vccuATUKqgcyqkCm+iB5QJT0xDSeB9BUVPr79+CCPZaa4zlS4lX5FxWAaFOP6E
VG4tdtDYbD4qE7vd+xnA+cel2oaW0+6EY5mujxYHwtVHXX/UbOl1oKSAuq+o9UwI
cPw4lG+KLNRQ4mVM4ROqlN5atT9t9zzy+OxW7hFLXrCXwkIMCGk2qqIuFGwunBzg
6pxJhL0ow4Mj5yoKQcMZiTxtbB/wpGU2wHhrbsk6C9HuMLH8V+oGnw7yRvo0vMyP
j6f+8/WLdtneoCGgjGmllPZGqy34cRCqafzgdqokcn2EXPApPUNukN41skeA7lnZ
7hJ6Q6Ag4zrcmMAxU4Yxa+MVzjq9zb9OJtVEnYAcgdIoPJvi1D5AUsCFtTmpzFoH
hK0YV+TeB11ZXMN60n+eENykK+0126Q9AiI5ogK5nSJDaIYNWlqrhSyageIzKSIf
IbGVPARnOu+BkVm8IxHF6MZq7zr2DkYT+9FZYYwBX/riwm59+Rhsp0fKU4xvBS6u
y+wzDXkywnA0b/4bfj/kYdFdLJakrmwOA93ihLzsLgn/xY18Lm5OdmHkKuKCeJuk
spLWBeo82T0lV/y363GBXxHjFcrPzHPjJvr4LzusiT5NXxmWdGI+/e0uTHv3i7P4
fmGx/liYk0YPeLWOia2uHeaTpjRIoF+/cN815t5w6kEdQ8cp/WlvtjYeRgpv3WMN
cnHDTxRMMZX3qIK9SbJBXGaI/GaS52V/SjAEIqDPfFeIrrhoKZLRrkB1KF+RlrRg
D6tnhOgwBrNSWKjLN8TInf3gY/GAb+NnbQUC1dyAJxCZGn9jhV0HVj9qmZ7PPwKx
IDG0ffwJuYm69cliG0EjDy2uX+dNv6C7lqswKEkwwfsqTdFD/8yxQMQ/yd1bg9bm
XG5ke9ri3m+KSinIL3avColVdaPPWMoCgHZQvAdeaEKpL4SQhlADoTFAqY61S+hh
aXKDbFlmwL8KyPyoWGxOxNmyoPXjZGN89/0hQnO18/Qdn7oZ5pZEkGmkvWnIszUQ
HYTSCNRdPE/6YvT6bS1uLJTpnBjhRrWVOnUf5GV/8uT0CmzOvmR+ovJ8u6kYa7OE
yxKHwujRb9sfhxIqN8vLTV3tpHwRW/0B6LC5UdGIHw+9wTn8VynMT1VaLkSYZUXH
A//Ox24D5r4Rk5uhP8c8YL7RRr8xVzDT+QJseaknBADDRgyIw/X7tSogxFuoXp4R
pMNa5whDaDNToM1oE81E7x9UKgW/XLtjt4eX/W3e1MY3HVYgFOEHYBf6pTEivepF
DiPjoZBKph1YRjb8X0VSKQcvX1BAoez5sL/4uuA9YtUKeRStoD1qNSET+M9oGnGy
Wx6BLgpEI4JigmUqxQwV2RQF1We4D56sxpJwv3frveAiiC0iAhbWKLsET1QeGyFE
jKNdjZLNuiSfRTQJz9BmWnycAwk7YvfOzh3h1NPcdOtx5L8Pb+nm4Qi7XDPrnl/Q
ZgdnFBvEXuptIvk85yKIFyfLtUUOae3ekSlI9AmHJNTp5Y9wAQ25hBCOMiHKwZA3
Piakrk+951O9SbDwW3KdBz27lpwUNqU3igUpAOvjfR1c1NtuQqt2TCdGg7HTVdeS
jvOaYLoukGnsRFJxHrPIqNrfV9Szq7Jseo+GfX4gnx/asXBg5r2gBmwtc7K1A3Vz
5SOUhBL3z1lE+rkflYRD/XluhzDxaMFyjSbypuPSUMlfGZaZM3dd6eBTVDfgbV0O
+zfYU47ru47+taQCB2Qu8NwaPOpN+3334k6nMMqsQecT2wE9Eog51F12vhBetuLH
0krjb3TPtpAtPryZdvl9B9KAgUiRU+ltKtXtH6xAKyy6CeOOWuMU42tMEUYL9kbf
KeduttyAMv13kDVhG4Q5uJO9NMtegc4I7NIB8zmiv5aFvolBrrzmFpJdOEh1W0nw
66TPAS/Tb2vbWcYFipoIJGjgo8YvyG7u1T5TsZhfvGYV8t90M4zs8+3ZXPuNTh2/
iICtpQRrgqws2qHXzAXCOWvbDIlj4gi/WfQ9nzNRY05q2F3EZwTTE8AFnQ7gtFTR
0ics7OtwI0ueM7zf8UPDoK2C4ecMFKITUXNmAzNyRK+1NQpgIYUXaopX93kK6DIn
YqeQwrtrGAqUi4smkmqjfCZKDpnPOpGLEqRRssj4u2c7r9o7Io18uWr6ZuSB0ttM
Q3+EgmIJmYZfcXUFHYC1fthN4njS0WB/fzCuYm9PHNaT59D7ZMM9Rik+wpdrOXRj
04YKrcVmlF6+9cEKu9o95JdwSl/QWv8dw1r4ezs91XgHXrj73QVpoldYMD1zvmqV
ZFtt1R55czIJaxCfajFBYnomuNHldbxJWHCrhi3/a4IutZ2PtsZDvQ/PwhCKfx2l
rLoWPwDQwct02/ROxzLgzceiyosbNCrFKme4ocib7o8Ma3NNs1CS91whArfIrxKW
akEBeclJvSIqteER4NIqerFuAYciCGM2pniJjwmXQ/PEKjbMYUl3L3xO7UljRcT8
ziOAUfNQ2i6LtiC27kXrG+Uitl13GpppQzxD5QN0UlgrEBECfUpPpAigJoghgY/k
M1uP+UHywygsRhFkJg3OLMvs9EBI4wyeyZfwggj5fsVyGWtTklIw1n+ZNcTAIbU6
1HXPKfZCTrAJa3KqPtzUsSFqF5DS/3my5zqIzhZsLsRCWpEFDVinbn0bTIV7DI9X
OV2aRBU6kSYLbzjM/lbK4Zzgqjv/jBc6yo6q0OznyH6oZEqF1VDgRiVc80b+Mhss
ScJLMST+iwAuBaD1PsIZrkVC9WQhkmGXi55lqLj2ksP6FCcF00CS5BVHqrLbsjYT
kyHk9HsRqEK1Zx8vKSN2kgkVDfU4vhWU1KfHQHQa/kL3qWuNOKdUrUGmDy2+LL4i
NDNwAECCys/kPehFHPzWqMdC+6lsZgIXaj4bv9flkCJWQ37Pq16nqVGF6dzI0u5/
ToaWZKBZG3IYvMn/blF3RgFdiRzzE9szbMgT9ES7AHkTDHQHWh2FAVPJ6NzDKjo2
A6ZpW8l0r8Zl+sq6gX1IdaleQIyY23rfVKLOr4GzVdZtVnttjVCbFJffzilaxZdG
r/SlDJ+qWycJkyxrnOpFj7MlL42y2ZajxLHGyTqxeDkvcghvdZtTx6FCCywSp893
pZIG2OR8SKyFeG2m4etoOp0UlGZ5cCdLuSQuWVwh0cw9gTPULaR5WNi7AHz04xUl
y/gD1MwDLSBXFMT89crnMm2UU77jeUVMab6iv1iLusHxDGIPGwOFhXz83DesSmQp
cBSYWZyD8F7rQabD5El+I/R63OJ54h+3cWSppcWBR+jd7u1JC+x2nNX06nSq9BUs
TstBCsjPGMOrj/9HJhvQy2kWSfk3t7ANoJVierk3gF2boRMpufDCqALLiUyDK3qy
nZ2s8XCklf4USMIK8ck+oOLXn1iw4bGxNNiSc4pxT1g2p/QQtsVcV7K5wXOxKiUS
t5WQn2dYMXPJlOw3sb36lmgorJl0E8Tpa5UHuuOWcx8hC3AOtYWYD1FP5TOc+6lo
hWz5z/nkYJGH8zwHHZQAMKtn29EAM64bhWQz4tbcHdqoMJbZ5teZDzsA1Rmy8ArZ
x1XAP5O9ilvmIdoebkDYO1aDHbPGF0+N+SHGCsOKc4k6PsZ2t6JnXEcXclpqo4G/
jmFVNyXp+rxB4TzM8Xnjenappj3Jz9wF2patjdLHQ9a56IvJfxTwMzHfaTCFkhg0
s+8GccTTHa41rsRHjXhnykmE9dRE4VCMuTt0GpRTHwYD1djeivz4estStJgvngug
ZRpI7vX3hJHPgNIZvds7MXz8YjRtyitb2kUFhmjaoTGaCO1T8p+tjpCwzPwG98Fi
MQ0rcq5izmIg7wOhUe9egWWjya4qxStGUZ/6+33APK0KAsWBlTJ9nH6MMGGORYyy
Vlnl+HPO7e7fIRSz1aqLqYHELQBFjSf+eq6tPvILAHlbW1nE15J1hStVBEtD9xq9
LmzHXqXYY3etfL4Cv1BOjoBt5KgvY+qfRsUFQ+NleAl3b5RHQ3krULojoCxQlnko
JcCRUVYtZckwoF+x4+2U+xx4V9JoncPwz6mSTb1pxgwwlpz7SIccRZdqAfjygt7b
pY+IFYZvJIFmYeNoWILlqYJa15ak1yJrI3qdpYVS7LVDai4MrkbzQEvAMV8TI9aJ
pUQ0TvBBGxao7P7bBB838Uawh8Pv0c5mrO4076fmT9iqIZvKugvqENDZA3XPAawg
Mm4mYOpPQK1NfaewwMnsG3Z5JGptKQdAC3KKG7BkXbwwRyg61nFXJZK+w7ZgCUyw
yamSUar47x5Nb7aImG2EzoEqBXUCXDtEGD5CQWa8eZ2lAwcYJL4WY3i5FwYE4E8P
0sy/fifJflxRndi1eZWV6zKOEmUZ84VqodUUxTKnDfW0nWAcAsiqTK25M6er4gZK
XS9BtlVHSjPKXpYJzOgA1XoqsThWhZ4tc3RwNIbZEG0vaX0sqWkGDyUgnMPtLHiQ
Jeb3aR3yHYfoakuiI0Z2znJ/OUpaLf6y8bD+SKeZL6tIf5JDlJZ2plA9ytzvhfvp
EH85LJ2uuwKTVLByR9cEBLOpQqrjYkCwRux4d2kVQKQGUsV/7FAIM82SAWxiA+2p
LcpeANGhC7nEp8z38tpUvRUOacYdvHeEikXC1owCuMUNV7fnUPzin/f/DG/Nl9bE
sfgSz+PiYKgVNnhG8grBvYGUwGbvz9r0jcmK8OxIH6nVIAqluTSNQ0fDn1zDQNdC
JcsXamqD5Fo38MKU1hwn79CEt1XCJH85aq1BC/S0ZcgximFHop+sTo7LQKn4sAbt
/gyTJmCGdNuN3CPIgAru5u0AQ9BxAW5G3MxEqmLWEs1dpGvHaWdGLjXoow9iyW8X
/JFSSZXPOezlF/VarG0VvYiazEId4vtpFH0lG9ehvQVtBaL5VHGWrOsOuNw6ze/j
DFkOLARZPxMowSGhN7BmEvFRDAx5tE4J4KvXXzSWXcwE7BQ1BRxpqojjwYUoHT+F
6cssfhPjF1rt11DXxziUnga21l+cQwQN/2GT4yqa5pLEysSoYXI3yPUjiDJfRd4f
efkQcQWER+20guexAB/noM1+cNqaLkbGve39IR/31evQCQNkwaXtk4MPb+cYXOro
MGm8w48mAZP3NNA+Wa1SNUywRufnvunXSFYRzon6LE2kSOeT6W5ZCC8+z9duKptV
Zlaweha4vhXjOluyJyiKY8/DRr3rqwD4qnUPRVNXB3PHOwX7rfXkhe0NzN+S9rVZ
iKJRiqsd/vJ35JEei7xRWxgJpYb8hBaxgkthmNEQH0G3LcdwRsndUxO7tqI1tS8S
qpP9hoojxGi56dfAUDFCTq/vRdVKuMHrfKWQwwGoIrSmRlOwrzO7Ac3bWHoMAAsv
8UwqRfr5TpTAolQuedNPUOpSJgGFwMZVHCSJInHb/onlEdb+HU+vEUqcnWy3EY7B
+GMQb0LEJxvdZ4W5hstIiKYWz7zjs6tSl8RYvvDrloMeLKQ8H7VOeovfryeCRTZI
GxMo9vProNU7n2AiT+Ds9MFJkwL+3rAGXnDwMIITp6t8lBAb6nS2XqZEhxjgzXMA
UjyT5oI9ClBajSR3qrgCmMsScKZcISa3SLOIPc4t8XIAlY8ydlNwM80jaA8T6gSU
cTPIXlaH8hN8kvAYWLGUzmxkSxmwa9mODEcLLvXK6poK8/5gq3UzJ3Ie3aF9zVGK
QRjVTtyXcs0hTxUPu9yIxJUXquNjv1MRhTOnFuMUOrRPyrDM2pkVsIEW9HMUEVaK
Gj/CNxCPjqzCeM+iK+eukTAYnWdHP9/SeZ8NhgTfvGwnFYV/K1BqHfqCzNjHW5FX
vAufODmJ/P4bAUhZ17Pwbae0+xZxgQbKHMTFIXHctNq1Ke1kEniD2ZR0UgMkXFua
42IJN2hpaJi9K2CtVyJJe3ROX4bbIocehTzT5Wbfg1t1hSXsDECS9DOMK+/kK9yR
Lmq7eQGQZqOa4Y2zCCCEXmXWbFoiyt0WPjvC6kecAng5bplkFUATeNAcJqFTV/Y4
Iv3zUNw4MoQ5+6vrPXUkSK2wyLn2iVGGvT4Yeq/bxfEPZcjzW9KjeZv22ztnewsO
VTqr6e7zcCYZ3xq/LHR6mNlRSriG5qG4Gt6fUhawtgUwYl4iV2CfDRWty+M+Rvfm
9MCQ+3fE5LzcCHFNDf2SAhY8iaGwoIbebAh+LKsfX2JeOKn29OE/IOH7M699TaE+
frUZgnVkAsy45KFQ5S8VX4kGwGK0EvLZf9TcNVUWtMTS4SszBKWc0vesIFocyg/V
pQVgeKKECiCPD+YJGsb2hG53KXQlU3Ee+P7Qbd5vcVV1fR+STVsBUsFJiWxqj3pI
j5XQMye/M63YTFnLdi+R1fmM55CZdAGb8Yg2VZLUevPo4eGrJzTB4T0dVhEBjquT
wVnQKEuVlsAx5YxqEoOTZqs2qZhDs4NsapI3agbHunL/e2H2yl4wzcpP7PX/BMaf
TkG8il55dbPH8YBdTwHTBlYcYqO/inUhvwiO5GnW6t/EYx1fCAW34cN1mAHFzBQs
pWoUFxaB5BhS/tQ5j4apjspqaoVLLjf4pfImnsm/ckeXU6xCryLH/d6hPpT1KqJ/
yZ2EZXPDBJ0c5RxJHIUKkAzXWwoXYtVMu+HcXh5fThh2xQiW5yZ/RhV1Ub90Mp+w
O6zVIjO3EP77v7/9W9IRX18aGBHSjuc+Ysiz46bdn953G4/TN0vTPwrViM3MUJY0
g7wmraNUxco81Xmj0G+rxWEQUcpTmFe75JOYBxIrdglEPqYX4e8ABH8R6nCFJyFZ
tYrzq5napcaaJJENNZ/jRViW46YbxypuHeh4ZiZN8ak678rlPU3FAFyg067eERVj
prhNEVPa0lZIcB8iDbJpdEf61ffBktCBNUZfL9Gvqmb+O/53MrnbgfslvRWtUbks
+9SxGMX0Uvum563bub5L4EewjEAeCMnqgagurJc2S/DMalqklC9t7c6MOKHIzcII
soAtEEAuJi4BJ05hNXc3Oyi8+hSmtFEPLdtJUG88bm0d4HzQi8c9WpgKJnMAKrpH
ORUX+UA++XV4U17fguDZHgjVP/mJzlHYR+g9W9d+PvFghA4Ke7nMzF8p/lyk/AeP
YQhudFrPBpovfs2nRQVFIEaCP66P9XjE7oBhfXona57l26ipskvQMeoGLXmnCTOt
4VD79uxix9myU6NhpSNBGAEMJa8nGGEW5IO5Srq8Raqc85fE4zZcaJzmryxEHv+9
+4eAK0zGzv9qcfcgF+t+2pYqGGX1itFtvmYnoUC1CpShIk7Ll2zVudFm4W5nKSRp
ydhAdgQg9v40tAYB7zLG9dmaJA9vvqegFpFy1q7jCLCrMccXih08m6BSIuTeFHLD
Qy9KOruNWmQe/Jq3rQDrSU873dhf1qGVCHJtdepGayk6LVeFxCYqx56Xqyl8N9hV
Ce3a+tZlFzqp3BriH6erfSmUmlY885BIn7gCCRlMSLaduIw4Izxrz8yg9RYGX8A4
+V7aBYBvxp888otBA7RCW/41/ZPBecXqOBSc8HVPSP89xZl1w0/k/55Fme+D3Cub
rfbSu/BJ10OsIdwnGfqjeobbjEWQQsJ4b02VAnwY2LiPk7AOxyXQL9KLfxrPNOre
hiZhFYqACaNbHWkFVSOy+iOc0gcd8kUq9/pa4ZX4sSW0XmJMzoG2ba0p1G48IWP5
cABqeavvs0qHab4BFpXN8EVkFz5QzxWxiP1RTkBO3a4FQ7LKnPnFp/YLM2h6IXMm
pucOQMNsFzuqWn1wuUTG4UzOX8CAXHphXsu+S8geobeC96nnBTcb0w4G2sIxPCQ9
s4RDLtit8cIJ49wcVU8KDfj4jmczqNOBBZqK5TFG/Y0c3cmS2o8UR7jL1iOIT2I/
04Yt3fuNz8pv6FSjAKxcl6XD5RP5ngheiTZqq0XB+fHHBzxL+Q5QCSGPizv878ca
pb2BbJtEDtqw1AFanQax2Ufio6HsqBXCNN2Zp/JLGA0WhQNqxnhGmtmInzS559f/
k5iRFdsowlz28N9o/krQadWjvpDU8EHpUzBlAUeeCYPMcuHabOwRFFozOOAtUqWi
zFBu2o7ompXbD2seG5OyUcNl1xHn1l9dMvWEbw0l6nLIGs8N7gy93B1SFaeG5Zni
scsz+0CdjTr+qT5eWqYSYMG6ljBOWZNgHbrW4JyM2p7ZZk4aqMfuBlK+XMtsqTTv
/sleVdGnfRu15WjevzTPKQ+yiR905YfVuOZoY8xAstnBNwh5uBnYlG3ZyJv1ojaU
HiqpCWMB9fze2iIM+fJlnAxVPsQEHutooGf/sPc7pPf2ob1u1qat/TFNksm6Zrui
BXS1OeHulOLT4Yy9aSMVpQ6rLtRNYgQ9PokUwCX6DmZwfXiCdzFPD8vEWgvhgcWv
yxNWMNpQL0FHvTrBcOjZPFOflVhUEdpULv812ZdeofBBhvIGFDSYF8QL33FYtVOL
eqanmt1JqlikA3brHE5RmTxh7z/lv06ZW8HLBTJGKKeEB1cbJua2zsfGxrklyBFD
KiuLVWOPjRAB2yOOUPC5jIl261kF7zlx/TC9zZhNH/F8J9NzSdYDXm0zRwk/n57k
LMSH5iNsl10r90GFedPYYwTfGLtRSSAeoz9EMQJOowkuoTMOsXXtl/RGN9PcRLR2
M0wsUiPyWzEUJj/llfnIRkwOzElb+c8TX/CiDz6GIc5U8ck7GxWO75FwXx1ZnGP9
fdeBw6Gq0hlNIlr3ZwtuE+Fqoi2kIsRV0qKKNgrqyL8BLWIrDomCQ3/zPqBHi5HK
wFx/fR7bDsI6XLlI5id650laTiD6GKk036S7Lx3aA+3tkH6YCv/prklom7svF6Ln
NN15qVYfVOBgi9Lnxl2DY9pWa8Fh1UzExu4y/L2TjO1NpNucBp0z5PuCfIo6SAVc
RryChC11zRDuvd6BCDdvf5Rr/9IQjPHEc6UVaLdQT5PseQYc6ZktdqJtWXcXz+hh
z/EJg0z6w8GlS8jrb/au/FOULaI1y47cqjPwUEMFHIg8iO0Yh9OInHxcJL0zXyj0
j7QQPU0FkhzazHjIS7ZwMvu8CwEPqKg35QznNWWZImwxg52FJ/TKjDPFGg0kX5yG
eL4nKPxbHwlGweDNZEum/9UHRq044H2jxIZHrEI+RZn7ioAKIstzTwZ69sghOcFB
zgI9vVjpUySdlr7UVOmzgL6b05actIzV7q3liIuDdAzyQb+qzB1NSME5UIEYGt7q
NiJEaOJRErd2zK76G0/8SSK2jrfkV85oWtrSacNviJo9DBZXS2CXwPK/oM8buL5o
r7KANMa0xvVU6LHwLVYacI+lsfRkEp1g9nsSAMPkQuu1G6dSV3z5I4rMrhk4Pi5E
8xlBcLYbBvsS5iInU9IXUlEERFOA+4S4UgnvWrjlm10b5/boZoAe6n9iiCiCQnQu
ksYUkdmpKn9Y/H/Zs6tZcpsOaWaJdeq4KHM02/g4h19Kwv1x7V2frDnGrsl4v0yi
We8fgQ0VO0lbQTr0BiKhoUb/Q5ujv+YNu6ZVOihWpP9Uv6/SsGbzmchFy4RVhZ5N
f/jFucm+96CqbXwqgzwueRTsS3HbR01zqwllbjmD3rZ3ts18J+Zuoqs706g+VPil
m7RPWoyvrvB05+LyuHugvL8igXU9cDxLFNSNh8CcK3EtBv1Fth/pSlXh7yvWSMyF
Eu9N9kbEACOXpuizo2Yvb0o+bXmOGGtiMi4vp1Sr9zxjQrJv3fTSRrakou/4FrHH
sx5nC30Yz1PoJQSB4BSz2IT9Ngw/WbX/B3yI4lbwiCp4jQ9oxC/3RFlHzhSRGR6q
VsTKdSwjnSF0hQyPtQsJLpUqg+nC5uu2cdtamkL6HYn+JHj+kzknfrAfe4tajm4T
4a4iH4xCZsDScMve3ntgtH3107pYy/iaF2S1P+D60tfquU0ErJ6+YB7U4geJXH/R
U3KK/O2z1vsdVWyjh5BhkrHb5f32b2SYDbVTIXJW1BDlAn5aWes14k862SAvgcYs
NkR/6s0kgG3JL2MarCUdmIDoUFaUjRPHQXuO7/ai4MjzLc4abLBSTZxjjogm7qJW
sNTFTbXThj0luifLPF/+V4ONvZPU+FeoIx7FaJGieVE6x+mJ6PFIJcu5bAEvX/cF
V+zOwLGo/JqSfGSwZyi472Vah48AQt0wF0iMO8O/q2CSd6tO3KVLf92brKybkpBS
M+kv7zvlYq+2a8PzMncw5kST6Mc0zgdj1O95JJDwsnow6OFUdHbv7VaonhS9HENG
omFt9lNU/pphJDxw8GaMrz7fSY9p4ADyZw4oPHrVH3fCTaz2ICEMYvVJesGBqiur
PxL/qRVI9EhIf2tpAGP9o9uPvZ1WQkPazOs/VRY08B5bCDs8SCiCXCthrQEjHNPl
x9QXRR+r+tnTiU2Oao7oX2atxPtALl9orWUFxcxcFDyCpcCReap2gc2Ygmb/a+nI
LeFhw06bHciYcEbk30WM0EV6K/3GpLwisX+qtNM0xMnGDP7tMs3YNzn6loxHZPqu
/ijfYbiZsgsieuQXucore3EvJcsLcxXHIrqs8mbWhEKXM1MJKDEyfhIPKTJViVl5
x/ZnXwP0PEwky+b1fBpV9cGPin5GF5oJHuQ1lyGFPM4OEvKH/eMYgJmR2JDppFjk
cGnH/vp4np3/uViVbxMU79yyNrgVhw7EGlbuzz40d42RqaWBbiSpOy/laJeU4ahn
n6HSWJxLt65PFjkQiS6f7Fynoif8BJfmwrRa9feZrkGn/ICodbYXRDFwQp7moJ6T
BdGP/mS0HGRAE+e3s1w5Z5deF9G+K8yCkV2rFugq2xyaHIuyoBP/OqrUVe+jyyZO
21O/ZqUwozas3RpzcY4kasrSf0fyLw4HnbweAqFJEGdaWa9fAHDtTGUEdno7fF+g
o2t4pSm4rRInpRUW9UtxQHdsSiWIl8MVaJHHWBfVtxOFXnVcRLrgEpKEIe37+03P
IpHy8l8JdNA7Y4E/ye7lVNq1jDPvPBBkco+jvjoSCRCWkTopO9ukJpoduaSUJ+vt
8bc0/gK2/ut+pysBqmA/1h2MtNZAMliU+F38uI+HQVzUbsPthW0eRc/WULHp0OLj
pCT/v3hPLkIxeRvpyLwnmvUd5cAhoXTRO+iZ+FFXCq3e/mZw/7qWpbcetd392PoP
IVx5rgoa3KXmNKR1bfBxAe8tzJCA6QO69ButnmILBuh78iA4pZxRMP97jzzchbeR
HxjvgO2x8DiFuuVMSxdvJj81f3uKS0zFxFzE2k65Ie0o0Um8T4O4IgMXZlsuggq2
fNAGhUCak/3h8XRAuB9YAXNhIy8hx9gc46tZgXknl0YrEyIrTxvSg6Y4PSvLBtRK
x6dVrVXu/0RB2bjYMMvlfCemMNrLLixtv+FyPDuKlr+cb13+95G0rlz+fKii9Upn
J5oG2hpd0iXsNEmNrhql5Poc5TjsvssYAT/iXVldHLwgp+N+georQRIZQ9VvcNXf
K5aAuzf9sy7ZXrW2CinjvdwvzYIIg9WByT3XjOJCfp5NXfyIVs7uJ+q6aNTiun9v
fy4WkxW3LDrZk4nPN1e0uz9F34h4NLHT/xBFg7Sy7+7xOfYNebQcoRv+TMT6QlqC
3FKTs8zCA8boR5wVcmShfnYKO9D0NCVIfq6xb9ug2gZqghmhcB8TCAte4j5Il42Y
0k8dLdwQ8VP3Rf5dnqB+eHZNQR3wx/BkIzGzkOT8TkXk5OhgzBIaMz01Y3qn7M1U
labYInMCNyfsliBrKuM8G6yU5c1Y5XXehtFucC4cT0nmhO/CyGEkZ9SQYqWn2Ppo
l4sGMQr2QGogGkgq1OZVVjiIqLMwb+K5qXPRe4ucpGOWldZaS6VPp9T7YOrm3jgC
9ZKdezV1Iv0cBUAInAWtBEbibyxHf8D3ya4yywFGWh3F09O4EBmUL2mz3X3nYTh+
Dtge83BHeEUoECWT2MojsOl41wqJS7DYFFCoDWC+pfi4PYD/9y+Ttr7CN3TlXDh/
/vaSySRD8UOn2Ocg65rgJh2zoswbWY3n6eeDB9js6n0XIE9cvIyEuaIVGZh6gSrP
SDfs4c6O9JVAA7pvjcrg9mkbiVl8j10kQnExOy/I2Hu3EkAlRkyp12m2fKU/YyIc
ZIQyeTMF8FfOTAASqcjd2lJp+Rha34QW6Po3yWfm1iagxn5uR5Fy+RMsES3lhVaQ
1rcdyrHH+iVDvgm9ks4S0sbVByuOVy5t3+KmIhHl6wiYJIRfl7Rrk5CtN0P+3NNb
rviSzKe1EKHj2OilR/AFM0e9zhqf1YPs8QC32ImcF6r8E+3Kn4X9hN9vP4bRofLh
m2nnrjPa8NRokDPZB5e7TVxaFhguGgfbHeiTWtOQmF2406NH5wyjEaSkq5tjaaQz
VLhhrnRsTtuETozpooUURDMKSr2ZTipqL1yznFsk5zW0/28Aer+V3NmWDg76iUCZ
b4BCbIUxQogT5rTK7tNqx8bjdtV6oxDCowhWkaMZmWWd6qq+DQFSlkDRfOw1Qg7i
poXJDojoCUhRor7KRAHKJOZMBasaSSSTgFSLcdaP4qlLHnnD+SoQgbWXEA0M9p55
4vWBKghSqatvJb1HTba/RZygrSG4m/oFjLgIeAc1kKkIbAi1Gjw5OpljA6WfpT5b
LTNqNS4JFXOxEpOgyPFyxvaJi0tJMHpz1Amy0DQXpJKhwnjFpJW5Vg/NhsYpG3cA
XVULsouJ8ZyWpebQsGRnzU79GX7GwZSg1tJuc14QMCHVfyGawL/X2WIqpbYghyi0
jkEW3+IvH4yvaB2AoCh35JVgdcw3fNWTvExtEi/GlBdMGfFymGpDPHsUmrrdEdyc
sEKW4LhrFcjKB+htx+PK6W+1IQINPL+3f8mRens1f2esDzpaJqMd4vvdPrtQIBKc
+0QAFKOYL93JCoytx1uhTs3BK2IMSdAbgDq95sAwvuY5jUvoDv14bU7U7P5yV95t
SNXUGorBbUKXDfnqVYDhP8i99L5SO1sgTyPrzE0Sq78aPZPwMMB5QhnRSjkrGT2v
9L8PsW4Er6tTEzx4WlWYKUP1km/5oZN3Gq6Kr4RCGwL6UeIaubRI+8ak9BKH2xxk
5v8N3ra8EinJ2tfZ7125WzRmyuMzUrm1Y3vnhwGuLZwdeNHV6spJVP2yVTselAUK
+iUVjbQY4DCGT3bkbgNdge9yQQU5LWQyBQVT6I0zSTdLAkwqvLqyfclBsKN9GuHk
u1Zl175bNXsC+fsjV1ry12rj5kcF0cmKtFrDKcSvh8pVJiS11VmA4hAGqjfGQFOk
CscueadzZmA00ZWYXpHu3yOZv9TQ7+av2QudMy46mXIo2Fmfuu8RQj9RIwrCCak8
Z6397SFNs6PQPXYAefZh0uP+d7g/STiS7iLrq2mH9rTJIWLZTpFPxpJCQsd8qszb
2qeH8OSy6ux52P4+CPCIRuNMzGApqjf9XYH74AhtmnLUPwOgKDUbz31aREvVuRPq
MC6mL1NTUOho8K/ULox2cC5EtmlI2Wk6LnyjC1wEHSPyUcKxwwTkcaS0mE3zGcuS
rOsy2YMC95XER7vm+tmlBnrawErSyngaWSBO6c3aDEmvGurKEaOPrdFVNIC7kFKU
ghW3w00/5Wa/S3+MpyWWJuBACVTu2AA/gXrAbgZabeuY2Yl1vsy+cFVvsoUqlaDw
IcYwApOPeKPBSloM7kd9Mo6B75PuI77Dg3b5MIAdTGn704sSsNmwDcfHDi/iIjsQ
YJiTyUlNDOu26sfColxLmFmguA3kPyev2uwvQ1TwOTKYdA/TPFZwzzJdsd/zDlZ4
xe65UR2dUeVivSy91hktiLimhZH+yViMKdgObanDgmywDRnoMFGMEAbs7dRI26ga
bWs+jYh2xEFbW2qQb84miilDpZbMPJeWOlpdrKMJ9N3hJmije0A0y9pBOsbdh8aH
98bdBrs9ILGuybOdDCw0W2qYmH+z1E0rVAHIZtFD/23zacljqc2SEUFzVwyh15lZ
O0j+2aC647np0wJqdrTUMD0NYVbaNDmNpRkMDUqO1wXvNr/SbQJa0Y1w7l8zFz4u
YngD5db0Tm0LYGpFU1v1WN+NjQy4xJaMsL63CQZVU5k7/fIfzc2zelBa1pLMTGsz
/iTXpm6V7gjQU8s6qN/r2Hp2pVY1dk1fDtzntJ/vkzXmSENm7NPf7RX/hG7slZV4
g0RkhcO83Jksy3ctvkBftd8u/p1qXDAjmsuvXUPhplXOt3xCVz1oLJ9PMx7FeB7d
e+UtDtf1fx7dlRnbH1TbPdmODrhyQHhnC4fZ8LiynglKyG3+IazIcffJHDD2Xl+d
JWuP5s1YxCZc5nTP5u6DjdI6wyCSckxtSMnCJlK61ZoByMJG5+ALvzwgO1jozVMw
OBW6Luaa/jp341fET/ocnFs+kV8K+j8MIe3l32v2pP+g8hNyNPFQH8EsdCw1Oq38
Ls+H1Yx1Vq11CPu+rlDeHLEjaA77mbRnccgczZM4Q7j1KUssnpajG5lDEqoULEW0
qarTyGth2XBH9CBR8uvIC/gyhOcpQWSicCqhdhVvGFzzqmBzqaTsXE3HGZfMXv8m
V9NEX1JWvr2czDrCmIbDoxoH9DL8V7K0peIJhk2a7L7B911YCK+drNPiJ/sAxhI/
b1DVdeyo23oRuhwa+bYvBLrKu6fu0KgAPFKxkTsGjCwLDU7RZlxQT2UdV0t2Hx+C
uiMEaRwb9OzXRvCEbA1EYcg/dgKcJi2CwQrH5O+gppDmkGorPtec2n50HhEUxnja
zACcEAUy+gy1AX4qXZztk00u99v+nj4SdozoohXQzgTnDtBWO+ixMCIBY24HNQaq
LucsmV6JltS38FiQXQS4sJ9xwAkxvjJglElyv+BdtaCcFTpAmieJjdyT8EJHJNYO
T0Ax2Cc1iZUbmgHvZe/xw4U/PbEFUuKznBc2HzsWV2yGkUdw2nB+a5kUZfzQaoDJ
SS4tNupTErWYSmujDwL5qzT1OBuxs8BOij0AZtR1ZBID2zL5Eh/+1uTRr4tmgAF5
yyuEZYKlS+oDkJ11JNQVMd+/ZAuY+HSghiMWq5mYWaOuyCgU3OUPr8N+28B+E9fd
lsP5l56IQZ59+jTGbqvXFWGbxpvQSGRlC5gWKF2OELJGCGTocyj6nxGZNw0LNkWO
ygRmJJ+CwaR6uNs3bwTiFAFSgAzKntmDIlnRt7VflnG2vgOSigaMvG4PcSJRvF19
FUahyGJx556ZSP8LVRHZ+LQDtOFkkHAw9+sPu4gT+zy9mKZ3EKyqMD7kxNj3x5O3
RKrXMh16H88viUIUWuUUOCxhn4Y+dCD2BxIelLy0e0cDjgmkDhaYh1NkBiPxLaWL
p8PVj+9oVs/MIEUwT53Z8YJEGSiJQMvadkhWVochs8x4Mi4SFVsqh558lf5Fmh7V
a8jBYl2Hh5qk0JMDDDIWSuRFv3YVaH/BgQ1dGoy+l9M0CJ1K7Rlp1Z3Nq2ba40wh
m9hODP53eKcrpGPYHnx8P6FtF7OA9L0DewwxG9yQ/8brxqGc0/6BLcrDE/M0dTjb
QL7U9pdRaesNc4yWqCIf0bQ5L/Hr0d4RSIp20onif9OnjQHi2OXks6901VYFBHYW
j+JObA554o7s/R5GN2x4A02LdNjR0PBzTLELmADe55s5IWoLn4o6FBoUlN4VNCr0
r327cxSLWdwFQ0F4BuuU01t7iVnpx48wRL13+FqqQvskqn0Fcz6CaLwWdDTbYJC4
K9VeZKbT6wYBYCjBlWHHY88GOWoHgxGBSN6zWICrI5dGMeXXHXgbgmSh2xPtPCoN
s9rMo6igxiySc78NZIVLlU+KltIuSd+nLR8RZ4WjQNO1niTFQE0EwORC1wgDvB7R
AivzMCSrW/yJd/qJqdQ7yTmAeiYAVSO4sWhDlEM6RqaeSYMaZvM5oEfBfr6yk1j9
Xm3ROdq3tbD8EHSpORSMmArlh+GM5KvoYMPWCT/qarPwTYM3dZEzRdn7Jtr7KYor
sH671ov/ezKlTqh8W+p1WuZJ822SCJTGtijlL6ifO8etANs3kk456aex0tapfOkZ
Tx0VTv8TNulZtdaYLZD1EN3Ynmzgm+X5ns1euHjtdR3Bp2Dpb2CD7dLdI6Ez/gY8
fYcZclFTHlnEpARlYZniBd6gXxwFqgjqhq+ftQ7uhaYR4EaGRb2vA8Hlcvc6sKdj
CE3sRvqS7MuHMQk4+wa0svHumEO/dGmQpi+tyux7AACig8KsjoB9OOAB9h3re0Rm
JH+vLYnnJ2mYCszRqsbojGNpupDYOTlhvTsYWcIRqGQQj2jUJbf1HoWC0BjIUmVH
A5tczpwsYhJuuh2CdKpqTIoig8uMlhVkL2myYoDb6BlRgBxw/BLG35Ltt3frWhuS
wreJJgUmGJaP7GHspLdPMGlNLQoBKUxPziftjRgeII1T415VI7RpLBtCC/yaoDJ5
gsUXhqOBmkOuR16FGe4uiiM3ZTYzBH7OMwOjHMpJ7MF6y2lyLKfvWtAJL0VMMj9m
NWI3oqqn6O55/squE2VmQEzlsjoAqBDcFNBTM32D4cu9bDwTa1pTTO0dD5W/NiZs
1zT9FDuG+V+pWuxykBHKdJfx08C5pXTjWyVGEJZlaQvQ3sjVVibXlCIRK1z/RtCn
2yDcy97qY8j1igG7tXauYcR1ae0OqyCk6PzAn6OeqZ3fbBWcP+Xe592OUThUiSIe
hwPuIm4ADR43Ft2XoSi3FQXyOfdCO2q2QDx+sdUnQR2czyN13NNntoxDD9gMe/VI
cECFeVVqs63/+jCcJL+M2xQLmQ7uMIrvH6vQvn/uv5393YsbKymNKwMtN8PYY7ZN
DExgbXmtUz0Wr6JvIQpQjA7PL/unebYBlwTr1bX0aTcCsMYF9SSB+F8JE7qObLHz
Uy+fzesbHDVNnp5Y65wkguiVbFueru/Gc0nepylDGTR+Vq+F3DT3M3MxxOvOcQVo
GDLwkIvUU6v+F+x+3zBtv+wuGhoTxxH47z6Z3xnrXQX32DvhenpXt7xCG1mj3v2s
7B/Pf9H+ZaGItwLrhUuA98OdVhcZxLlyHhaOKR0T6EEOCaV+rY0T3Pm5uIf+4WQZ
1Hj00MiTWLjIOo7d6yVgVbmr9Qp/OeieUkM5OoRp0hsyg5dKxcEGuJw+WWsHJqxY
Gl4wnWoVFQI4+kDK0ZljHNRGuJSIM7NZJaula81lr0HdxWA2H//h5phuAi099wPN
XVItih4p6ZhmlMEHWGgIhJ+bM7p4P5+r6MMIPII5hauY9bbqdEVe+D8uxNNusSw4
aXiIrBHNAkMq8w+uzHfZWdFhP4JbyC9WTh3icR8ET+qVuOrySd8pKiAySgBVSU5m
7Z1TazfggvHhpplzn+95Jxb/50thjRBnKP+IQtSRo9wMkI0Si8qlzPvcZp4H9/k2
ajPUhux5sGxbv4Z18dS4nWIC4pbfzwSrHBzI3eHpBywHSzdZV8B9VjUCRMkc1p4M
P5SQWGxHGPK0jnbCmJThKLWOKRR7kSTOKgrpfa/8KH4txyZWPNiUL52JN1e6ZEu+
txt6UhxiRSbU5cBRjk4MepzeAMMFowyO74/92bFHPI36HUuWAv9XW/3LM0sGwxX5
ZhRlCIS5sEgUzZ7q2cXP/Dz8ujbHt2FmoJROv7Wm62GtnM0x8IksvmkZZxMUTdMW
OFIiDXHLleyRJ8ATWnFkG4U5MWyxYcomJG42MimXeCfzhNnV9KH8oublA00gJ8jM
h2tdl5ptmvFPaDz3HZWc6R/4wWdcZh2eSR7cnZEMU2L+QO0671owS6NNbMLpsnaE
PILZyphmJpe7FA7zmM0fuNKAu7XOYG3o5e6St4qLM6/AQ/tMB/wZSFSDeflsHMbM
PYjWL2CZwRt2RnfGhD4PtYrEJgnBPVTUIn9BSl9EQwMDUo0aUsiJeT7etyxr8Z5B
s0hlsumZPwksaTOZ73lOe2ZKGPsFHG0jKjFSesJl/MoUwtPv7DHSXTRhTkCzoVng
I9iVCK8n4C/EQU23o/gcizAjVmpLDEa7FO33zf7UdEEKr2vI09FrQwfWaaBfqpk6
hdhH23wLoyUlO+K0r13AFdC9eUlo2DsjaB+VOjkiWprg4+uz6NRzKf/y06fpBZyC
ayNAvIdmSj/91n3bM9ziz84t8jZOEENd1tiWy057gYth/y3wLfGmVLV4WWQbAG8a
qmDxC+IveFL7OHpl229ofI/nQoYfGRe7dCCgJcFGZZXbov/aCDUqav7RWK52uGV4
EsisW89IcaAGgwovmLds8rm1viWB4HZgXCYEecjRyo3Z/Tt9q084nWm/YtoHP6ye
3QLL2F+3Hu2/4104yvIVAnBYoAwot3gw2y3M3ZrEMWplRzl2aqucZJSGRby8yjzz
QLci+TaHZZHDTcZdcwHQMNWhlkpH/wmyNV1KB7JcNbXjsNIpl6OYRaoEtMQozlNF
wxP1Ej0B9TcWnPNL9lNC/8BnXCm0TPp/h2y8GKRhqeI6347X4fXy41OAL4A8wcYa
CuQlE4L6CBMYVwFTgl9YcBO1KIvgAiVyESpHdejpV3Kj060MzYMaXEYpbFP6UoNu
WBIsVrgwhU3p7tvolO2zBEMgHiacgjrddeF85sZhNe9X1SUI2sgVNHMGmDiXDDUw
jGVWqlVcykaOwKyT2Ty4fDuvRxfxLUmlYBeayg+jPLmC7vRSduQaau9gF8dHXXrj
ORWx8DwTjyUGKhpHxW9iKAglr/qnCuPk/lf8kBwKN1v9zYbKVLRYDXejuelcwwvC
5UVkNhhgmfs+rjQhFTl0j1wm5mE7xbzaddkxAFcrfCP1JCytj5C1UeWQk40ReS5Z
lvxtEcaoGCGB4gpcedkmiEljNcvtLMTKJIB8qY0P1nExs0mVGzW2zfpGB84Ataqu
7Gjt1SzEla+noUODM7jVad8tJYh8iN8W0NKGm6VOX7C2RWqrI9PHzV9kaAvAsEVZ
43slxel3f4/AszvHyTyn9AbGRtLoDO2OQFxtbfaI4lqm+70rDcGaGlOiJVhY/RQB
2R72vbNf7suBZLPUy8Ow3jqzOgIQnsyCh5WcMOp9gszjg06VuddOOx9+RWLWLXl6
SpeDDhG7/vcZa2iMUBmlkq61Rz5+3IERDGf20XQCn7YOxJW5KKipDwz20ZrdAvl6
QyFqd7H2pRe/RCilFqzbBERNqwHitTd6k3qmOujASV59zrdAvxBBM+b7GzvCjvfB
lGCk/gekVexJDdT0EjE7dZKTZW8ILfJrouXTu0LyDfsjveTvHzqLtKYk+f7Rt4Fz
H6sZns2VGqvYPC9Cgr2HuDXO8gdOhvKTycpFgXwPYh9p7dL1S7Y2Dg3Hc9JhCBcp
JCf7Oh91ORGYPcV8WOaoWzRn6EOrlZZMCuL52QCw1WjXZgED4Hpbv6u65kklBDr4
HnVuzvTQxG9QGVTMMUm6kQhoX4CL4mQlH6ViFZLIWjjS7Xz88+Ioc1GubPNyDKB+
cGlNWOoz9QKikC1tOpxxQlj4itjuvudOnffDuCqzCRPok0qcn6R1JM9IBbY33JNC
1+MHk9STYiRQtxet+PekahUVPdgHub62WQFjC8suBi++XdvJTUMW+QdNy/jG02Nb
MYFRNR6jCvI3UHxW2Q/IoXLUEADVpaBlkTK8RcFx1a4PvEJaX3Ukfqgx3tHV6u/3
PY/GRSBEjknHmck3LrezVJmIKihffpk94jq+5f8DiohOIBmMtjtAg2rLLLxF5Sza
36BbtxQs1Nixf8+ZVxZ7BdkFUOC7c5TuyqM4UsH5acSaYHSiTGg01RdHIBeZtyRx
CucZfz2LrtaiQmzRDBLVgAvizMfp39N4nLW+iZ84wt5YpJGfaHI+yBlzGsifshgR
qvIt9XsvSdlstqDdWBbbEEu5XBg7UJ12+ylbPLdH5VhPpWlqjA7z0rECm4aPNMWh
ZARvIHzFCHYwoFntk/SSB1YEndgbfdwRS//tam5sR92ZWXRYeEBwJc7/n63JHlHs
gSGaogJslvZhgHE/Xg2aVjpFwTnUznfO5Y1m+Bq65qCOKRnVjr690kgIccNotMBf
t/vJSpa4PjO6a79F8viBhDcvILY/HFE6I3irWahHexDvytu2mjQgfhfsxY0mxBDW
FVJpICrNIq9YuM4Q1oWj2zN2Wj436NxxR3bqF7JHfAiUJfpZfv/v6vTPUMsPd6gr
kzbduSjq+0jqIfdLSNhlUik6fzU95YSliGZuwZ8vRg2I8147k8tKr2pyVtoVCMck
gsMA0PvHsvPeVDjlaP0sk8YmoCHXajuv4Qs3b4l2uIZiKgolRDEBOYantteTGnSW
NMd8Jagn1CWfwHk23VE1EJVRX6CPd5S9QeUm8kNh0maNfNiYqrlCz8H/tUBMuZ1G
NqJRmzZupQOl1DWUq3+gkpsNup0LU0Mu+Xnzx/lteGxGXJVUI03RHPtU980oGxqi
xs3G+lZCFDPBUGGzlLPNpPIcOKhGKgjJs2mZAYg0OX4vDl3wa98CY5RO50aZsNkH
fZB0axhsxERV8rg9JBxuOK9yRAH+P+/6inDwJK3UPU+rnNLrM3SbABQFRYOK6NWV
LUVDLRxFhlxjDj6uc8EFFGB9gUUQmR2EZ1z8Z+ENKARzo00lOjJtUOg67zzkZTz1
4z0KEIXQceQ+XlFp8l0eKpPmo6Mby5WCpYZs1za5tESBd+50It6s5HEAgmIOheN0
GnC3di/E37sv1nYsVhU9MwDelaMyPHWkkbjZcRWjJ8lcjupVx7tOQ7Ij3wjLsRA+
CA7E/Lkrv9NjxFZ1eKM3ssAPG6z+zvicxn3uXhHctGxti9j06UW4KdJA8NmG9P7x
EOc5N9Sk+PnwuWRMbjAjaDmgsyZSe0Pl3jv4cLcbT8joM8687WvDWWDMMybGmpOT
L4rwuSj/Gf/47UuagnIfSXkFQi56AzROVmN4hoOxYaToSqcieg2vRcdExZzcojIn
hBUvuBFjSZoIG5Bl+f9oEpVU9Pb/rJ7cuPm9/Yjl3Ub0fWPQxYel+IWIo+TvTTSF
GPZk9DpTOSfnl1HtSeejWI2dKTF9wsVs5fdMCuPwpGv29sdIdM26tt00k333FoVR
yPHfdt9DqFE8NzsTSXdupLB/HcTo+bAHJZZm3qYFvdaEupDuOP/9UvHGyR4MR77m
toyO3fbd20RhPPKhCiJeWm4SMuoUIpew0HOu5fwm8nUrAhtA2ESvq6bJkAxtLrea
5vGhOQhFyCxWQ6VqIHsNA6r1u6PiGAjdcbsu1H/Fma74Un12J/PYoseetfqYxWQB
ndsHXCImC7YJIYE95UuY5rXYRvJsUPaeLEnRQrxziD3qd3vbG0v/eSakA8GOJlxt
NNkoiioO6sgGt2bHiB9egT4rj8AD8pt4SCL2UVw4wOtP83R6wYlRaM3EvoavVVht
MO5Wu5RvEOvOmStJs3RE82TEAohjDkaP7ki1000kncchQ3X9Ug8ND2F9blbZoCh5
hStRPtYAH4XIY93G1XO7fMjQswp5Ut+s7C5PWrboCbXP2f8woz8JS4RHmJFK4WUZ
eSIqemuQQB9cfxhZRvvjmqeJ6JcIhpA/nbg6uGKhRv+cjr8/CxB7f9oIlVXpG2+i
ZxFloAU3jvQvGOfoKPBdfCMUmbGNfPzgIpv48wEnM5AR9ee0LymZlnXnZqoyZCY1
HC6n5Wzv/8rJNkhkJ4LGdvZdkoZsP63uXavtN73ePN9exG/2sf799340f0gPsDjr
n1DemW1aHvjPNSRc0Az+j3qq3Yvh9v2Y0I/PwgiCYCaiOGGSACsAXe5ZDFRxIay1
0ls+A3HlXdx7ASAz4TegXivI3FHKDAvIp6mByngsZpblIUaSxcB758V+7Pw6BbNa
hN8SghRwOTwlj3xWcZvYdQZkC9vLMaKcQjVnyiu0CyQ91wFzP3DMk10+sa8XRZ01
qVGSsWkmGRHPOAVW4R4GPgLVeh8XHfJWFGtSa/iP0qj4GxLUfyj6Ag/3VnO2AfkY
/6sHLGoGJzsLYKOCYkT83qnIcEGvfi1ToPDmSAgJGU58LJtq6s0akCok4Y25jSDy
zMr76Iy3fEzUNaBaiFxvRhRTOyuP00CfFjelnScwLbaOH6S4wlNeDVGrpBn0cMqD
+zZcm9VAzoggac+7vKkx9NwmKuT7da+5qUtFSKSH55LNg9f8eF1iaogQjw2bLz+f
TgvDvxdWIBUa/at8KjsnvDE7fHXIrX9nFgAsjRWR9/8s/ginm7hMZwpl736sDMOw
7IijMMRGMowMcVxJ0SjEOlv0oYNDTuenvCfsaI3rs3R8UNUsLmx393trcJEra0Xv
R9fBzaSVMEsVJ8/vRdtjuXg+15x7eyxNB7Zi6prFtFDDSl4u1kK4H+YfCcY3KYGz
Qbe28ZVOWhksAbfiD8x6D3NgR9VseDDWsW7db9jHtd9C0BAd3TVs36meryVO4hQj
CUtAAYkv69MWAk+OiUrsqQGAzqhMUEusnAFZq9piGrsEcWFYdvPUG1ureiRn7u3Y
zptTZRaKwwf20YT5uXICkE3kNmsucWKBeQFht5mu9JYdVVEvNH2hYKIF5J75DNe/
US7BRPLtvMr3hI+6Vw49OjCEXi/ePOUkRPE9L5tBk9hHuZHZCDM2sUwrPQsA7h0b
zDg50WpZ36nbK4q9xPmMR7wbnQ5612tjcks/lF9Yj4Ump17WoM5ia+UtIgqOvkZB
arrCQ7zesfD4r3qYsqbdu5XSZsvwp4D6Povxt3M2n7dBRGD9zD6WYO3QafZVd+r+
mhaXs8hkmK68k9ax08G79I8+2LDE+RDskxJHlVH9f0wCKzpTI7VJbz7TMdfE2DbU
ptV3q+Ts1hm/mJTjuMOFpyJtkbyxr8p0fgHrPejIoNKdsFfEexsNPeRPn7WADZfU
IOqlOHddoGKWR1apcBp/dHyU41cVvwZFXr/5B/Qb/5eny+zD9wwIpS5kpZnEmUmm
CD70llhr+J0ydNC2p03mGQUlE9IgTse+8rrY1m862v78k8bocLgcaRtBPJOjJvrK
oYpnciREXPYpYWdDSrcn3sUucmzXu/sjk01cWNfoDij9wI5NIQc4P/ohZzobrrWZ
4qSfnF6tyMzuIpsZX4jlw+RDgSx7mJkbEBvZ9zah9InHBDhVIEF0nOpY9Kj8rIFe
iScbwZY4A8FgXTGRoqLbB/Dx0jc/alJGgmIdlgrlpleWyZ77xukDmhRzEdc047XU
6v0pfwGN6gQqeX7l42z9jpRdrWSWtJqutB9igsZgu5yTPWU/ITBEfxm2guYUiwUP
vN5TH8G1YsmevnJbbZycFL4UiBg+Gyb2UwRSc3Oh1uSH9NC1jYno1kKxERsc6OV9
tFDRCRWeMAc8yYHZOygsDuVr6vc6lrp9WKF3slRE25fqQeCL2aMgsBfj5AtaV6bB
EYLt+uX/mTDCPv/i3TbBsCGy0t573WQAlaGfqlJT5pxxUYo6JsqMOhIhe7/+txOY
2/UsBV9CSUzf3l1ZOtsgIWckqfbr8X2abiGe1RvW9IpBb4QzMSaokENCKhJo9ZqE
LPjZCR7ELZN+P+73ERL4hLwvgvTcaGt6C/YvBcTwhplKRHjVcJZo+N0w6nLBmWwe
BmTSP5SfE5ylneRn8TTLe++eat/tAbYLq74mTUbYOQ2dHrCmix1Gj1pI1hBMlE7q
9M/wpBKKWrurOWwnA5/UEdc0s2y8nN4V0sRmAmi+M0fevmDQduBL+rqyohh6lJ/Y
MOdJ70BKZSFPEMX3hbRCuMC0AmeS1TQc8XwBh0QgOKhKJ3EUnqH0qphMWfm5l13S
uRlyHo4aZe8afCUC81vEtKJxsBLUN9zp+6FQ1zxq5TgUBESat/WOaw7SkR18miLG
P7DHylzgOR//RJjdJWCVJhqCIB1IjIlCrhBBH2v9f3218JRW1BrrYm4xB/Mu2Ydm
XFftYzANYwscxlEXtBHkX0uRYF89t6ZCYEhJF0p/2ZF7b6fURxyfhFZ8ifd0YxOy
LG/YHn5tt3/+piGTWqk5PdFSXmEgc2U2L3CcXCoviRJ+ft5hpGFT0lyKfQawv9HD
6nI3bhfmxFcOpRke1+2xnaeu9U9ssnrtPeRPEI50Pk/KgAWtznrULL3nkmS4tT0+
OlOqFjsdIRTNDbOsFH8wFiUAPTxw4/Nb6Sc7bKU4pxF90IO/rGCOfW3yOSYg4iU2
HEKDJfUaBUnvcYTwt3xv4tGu1eK4PAOqsE1fUmI+XFN2jCrsLnujJYaF5r7LL2K3
dQwYfY5u7+1CxiJukLmJwTdMG1iQxL+fpohrDSMGH41pupAIQKe3ng2sb3nxdYs5
AkiZXBTGGBZbSpxhOuEkq5N3Rj2PQv5mrVNzhRaFuuNh6h/YQMRGrlYQtaPJYGdw
lbf3mPxAr88SEpgHdG3uHHXsw60TLY8LKDbBSgnkPwxLBEIkaB79Pjc/WaQcEQzS
sMTPKm6ooJof4zLt6LCjGFVJA4zpKN9s1WDy4UF0svCuMUlGM/mwptbULmsyohUp
5tDqEH585ZgQ1GNUhyxEBY5jmI/aDxVcdPwox/bHaFMzO47LoL6/cuYJ3IIDQsBT
7HHLY3tA+Er6LksGJb2URy3J82ewNCGHqe+1hjmvoTnQNvBZPv/5vsiKubOK2uqu
IhajIfZoWgRl3JA2lzcY/CxFoGEY16KvCh5ObXztjhfd6lm/lRkq5yTvFI3bI7pd
L16LmHX202HrWClAqF3vzrPX9e19bN9zGlnWnufNGhGS7eUFzh6sNZTMYYOMBZBW
6hp+euDb1oEvCOEd+uWjacf7Qc5NkCiQZT6uNYm8QyNYkpUli4x0fXm695FkdQYG
0yOqTV0BPMmX0uxhxDieMeP4D7eE/gmoNrvYS2NtqQrBSlceiivP6tbVJbKU08Xc
X23VaSgATMIdUUt7DRsf/FHGCEpTqrdfIMMcSdCTl+IzKzrQwzEARKZAYKSVinMP
5ltAAUJAHdAvB3/I2152ewJITYiqhP+vFR1tXdImffOOBYU9xwdKjBI+AZiTvPUF
9zqS3CCVS689WE1hqmChIpGo4Kp7KQ6+nH2BmA/35oASuAeCzriDZv/FDlAt3rE+
zBvjzBlN2QHDDjC9JdDNQvg99O0IqsBoYe9F1Xu/8SJZ49cjRlLdNiqRsfJDZ8t5
wWbAApXXAbXdtvi/sJxHd50auRQXG+GqC9Ni32fRPUwPCo4r8blB+GXCloLNxWfZ
O3ZWAKAvRCZsn4ze8ffufaT2U64DkewIVC4AynY1OdN3qEto9FIw/gr4G9+xQQZd
E4XuUSlyQzl6zk15+q/7jLEkUF78hpLbQPx1HCyUEQ/G9TAVPepofuFQEOph3H10
umMf+qS2tSuw3X9AsZm8ehhT6i9rr20zz1l2lIo0tFW7QRsKXGngatMOuDLXAZzM
hulM3wjkViDQePRUkz/1ypIZoBxahJS0lyj+WTQJl30xaZQvrJ1Tm1e4CZK20bnE
61DbnbTT7pUQtpTrTuMxl2aeq5kpfa3SK6LYY4F8mGgrDvOElfeykdxhRmjL/cs/
e9jUi48jwZaDwnMGAB7n2BdNkra4Ux24RQav3NaDqzQ4LclabXGT44BtlQubiQJU
I5S+zO3wFHEKzlAZPh/8Ju85X6dGMRhXNqkZ31jZBDUzUNYx+FBW7rKi05EDBoYu
BDxtFezz0MONWgz3w9FQvdPZMllr0+HdkvPAUuWrPqDmN9CX1WO0GyIvRsM0Q+ja
0P9n2fLh3JaCWVgod+j/P3eB1LC8iNKKhkfaTBfPmlHPYGgOGM0aCU6fAVqQ8T5q
JJUQ5FGSxzL0Tf9OYPflwVDDE0RVXZntewDClfD6Y/7zRNYk5UsT5qDjgPxjY0xe
XH+32nHmvU3yTExtIQdnZcKNtCtmrUz0ceOKDLKSjMand1/ITGvkQkqaYh8OL+Y2
Q7RSTklSyBFtyk0ewRDqdTUWcAJLqrU2pAj8BR0RvaoWRLr2Bz1o2akPuChU8VvW
9C6CgaMMfrgUk+8BGSeT6q+KhjfQDLFk13n4kAqq4TaXfO5j6ncCEBJ7vT6XLAHO
3O+RQX0z5cnmbG/q3qnnH73tBME8PC/L2kt4WwtJwO7utNzz5l/HQWkARFJKxiEE
HoSsTX0YE5kVMBYQ56AaD2Q8k7z65NafTsEOKivSMOoFfrAT+TL3b/5Fpv665Zn2
QdApZOiGg+Eyo5S3Lrfc13baTP2O7wH11yvBnxkZQLE0ZEKFJJY2IUIRaEDZgNOq
UbVdJjaacKNeDFI3PYbymRrkj3nLDKLNnQ1N3u0cce6YH0hM6g5B5m/HrEX7L1Bx
ViKa3SrdtwCFX85bTGVxWKSZx0s2PQAfculErWBLGqhGiPegyzVBl017c9pIQiSp
VL7LCMdMQHtW8VomjqqlPa1UOwT10RixNfPsM45/Jj9E9+4LFmUPTK2JX4Q4cfsb
XMih+RCfpVGry5krFx4VYpC7lAr7b8G4eUbZJwNoe/t80UukoWgeBMYepd8mBc0j
qYl6OO8Z+cKuaTsRMfB5Zkf9Xkt69LHy7mwQaNRN7HD22/cwWt5wgd1qeJ71NbA/
+Et0TkELvdpGfGHfMt4L++rseNpkZPWmXWPsXp3/i/RUZhmiyHn+oeT4+U0wYOCo
C7U8CDyx6e28R4s0wA4UmNiu4wzAyC09yj5JeC7ChiinsUMnagUxAskmSWM5Vw8c
MJ/s3WL+VxGjIhGTmDxpv7mG/lixqEHUsQ5lyisfbVro+w329lHbfdB8a2UABv4c
eIkT5/0jXwPhzYQe7VJhGn5dNtvd18tevXuwE6sfDeMJSbyxoyO90Aw6oOoC4nsE
gfjcRXDD1HXlC5e7je+JJi7C7WbMEhDB2oPP2yDMw8AFSJM4B4cRSZjhp2pD7Ed1
xMxzVZEPAvFgTJc2sAefq0cLX0/NTAK8jQ1JrtrqY1ZQmkxKeN/tzbmV0cWDo+lk
pP/Z/mTm+t3GXEVvbwR2qqtTDIn2x60Wpq4Ng1d8uQ70O93AM7nc8yXcurQgNHwN
6kI7DDFCzW2dd7B6TMMKjdQHzNL3ahbujhe+Uei+r6KohHgGLOH9xGhePAaFJ+tE
DbeaYVBcfjm4UqCfL+Ywfw5pXom7qy+5xJ3mPxAb91Fcr3zjEjhadHuoR5oiRWG5
OGFjiIW67G/2DImgy+VQuU9kUfhNtRlKhG/vtoxKua6LglJlLDTi04ewYUJeqXUn
n1g0+YhBlBiIm0Ffy7/ozX8Mkfbw+qEvV0mEU88fF3Y7I7bU1YyUyry8j20BNOdx
3vrvLmohLkhVallKJq36zp022uoMypI3HY/hXEil/yO/Wxk+FQfkySmAD2TPZ6E7
lSCgKUwFNU1YsNLIFu4rQNEkY2qhexWtvUBAqKgL4sOC4n7z8CReBvewdiviayAR
9hF9ji+J6Woyl8x/lBDlZDCoivEUuAiWudAywIxGqM2ltER4GI+lYyOmE3pd+uNt
782WsNN9pKy8aFGJHVSHGQPiEreezGvTngjf5UuKdL4tX2lAhugHG2qZgSWI3yKI
gg3poqqUbiiE6732SVypI9x+rPllFZ5dkKMQp+4+JqWMkqTc00tCqKdJo2lgG9pR
EvBPd+VAywDnfeGP2r0GOPFCugFqdpFDDoP2bLAkKp/tPBdKxi6iJ/bpBX70V+/1
jW1HKCxhh6Kg9ny9QgwDsstjkGV6Om7TWj3G3au+uQ0IjKCAo7rkdwVzGrhvOUBD
T2pViJy1ULe+Bb2bOuWAPWcLKMlj+M45G3cbil+AMZkfpqtsKUwJftR9t/S0N/Zq
XjB0Y47qoWZB5WCJ2R30P+4NldtcRGpakLsHKSoJqcoOKOBA2i4fygwCvysjB508
1fF7k6woBJpbCxAFioXKVDp4vvfsNAeWdBzaGzWHbp173KVFgBbz7j5p359Pi+Eh
TQFJvb+BDejej0Q1HbAHGM69cdTLnrk8FIv1vtsYu6K75VQcv6ejK338blKM5aBZ
M77oXYIKubeb+5JoV8t3/NfapvMUARlzoyI9w+x6/Xz7Jqy4oQ+kWpZpRGZgCGdy
PoyzgkjwQkFjcP1HfEALdp+uwxuGj1yxkWVQVhMxcms9wqXcKK1q8utxWyDKn2f3
PK44HZlPW17siq6qGeK+XcqjnHiDb13GSB29Y7XZZdHXc/6FJaj/ixGA2AFuDi9H
/uM+El0znQLmaZIZUct/2xYvSKFUjd/fQGiSwG7eSAtmHmPOl2s0CPNCdyBQqdao
3jkm9ggwWj97HkUHQGRLMe2FqZiODztTSDLxl0g7SeFz05jJGW6jbToHItCY20yw
bZf297QscmquKDnkhFG2qePNa8OErjeGNUIQJlVzMkH8nxvH8S3eWPTGtxa01Gfj
JqJOr0mFNNPO4IutT83EpSFHEPNtKR9UPM6lKhbVLCD0NqUTZtNA4spsbwZfvlt3
5/JDe63QPfoG0sW9LMwMMg85z1EB25AdreCxkU6YAatdzH01RwySy1AzUSo96Hq8
IHVD7C2zP4i2QJCbE9shXDoIvdG4LACA4V+FSTmNuisnDqjRZdpGaUwtatujC2bW
RD42TpjnKlW9KyWRizgaH/eUbNrc5WBQ17nUXCXQz743HmaxMjpw60iMSoH6Yg5k
Jt5WaotimI394EAVYnSkdxvaB/UO88FuKK8BkSl3cdsIJLwQCHPo+D3PlyO3Zs+i
CCTCrJ7DwKANRrFLsJr+O8XqTjtXVssuBdOdNiQ/Gh0mLG3oKdRD6zMlTprAKQSk
VHAN/KdiSsvZRJgKm0dxEznYTNfBBl1oe03XmD7FaPmVjP/YbOe42bvI/4CnMSNR
lxEd6qMPUGfo7U0x+p6Ukn40jA8WuG9YlTcZ2+vRVy2z84TPDKlBrJCPDvhwjlhM
bQHFDaRx0r1U48cOQwJNLs2vgyo39mnn8XUgYQsMvpMuQEcAJiVovtHUjEdXKkTS
7OlowOfj/fhNa3m/HPxk8/QJguif2Nb2/7kxw7Az5nvOuI0hVa6lvTfGcOFG4yhj
Qo+z1Rv/WFs3LaYe3XIfyDsKGCRPF7GCqN/XAjx3Cfp+l4Pocanmu/m1gNcWqKAO
O+zb5PigyxCU908N/V6QdPoh3WkSM954d+Bb1v0x5DC/B7J2y2dDGlNifSXHtClg
DQJ3po1mOjYk1K+pmmjPWa5Ur/BRVYVi6G6Cgb08Sx0tRk4GWIbh0igSp31dkGue
ecUaBgNqbAtvbvWlKcXiJ2IKKSceMdzlWnXzSuGQwsBjE+5o6jOG5t9uDevjJOQb
LoaKEI5NHunfPg8dN+pvzbm4AyqqswXbZTOUcq1pkQPwK2vsjU1WsGL8kbmbCjvS
SMV0C/RaU5Y4WACq8CQHqCoCmGU+kUyaXGzyrg8jdnaWzYJjyXRz+WY2pcZ0nJMd
tgWHYmF5dClpXcWe+gRGlffsRFCS76xcidj2CEi8nzzcZv9ZSTWs+i0yUL9mSzqH
OO7o4NiQbVsgl+8oyMDz75Zkg/garwjWmVyCaJYGx7vwMW0ykkdFGVn1mesgT4w9
ZPht7DPNJrKTeHIbbBAYJvprTJhompYi5VkiwVju4GzwysdrNgsR1fw7uOVXrQB1
KKM4fHn3chut3rAY5lnewrnby9lgnNpFymwg1QwbddCwWHnQChRo5oE3vKyo+HfV
Yi74e2WBwmzekFDtKjesypvryBPAM0ynQ7P87oDo7//O4U/0X9d4tp8zv+FE7HvS
0gqIGdvTBOCEY+ED1vYs4Wc/69n1m3Tdtw5kBeNreJPiuSxjg8BiU7m19E1IFV5R
CS1ph5vpfk5Gaq0a7qm2ReuLQ2KyE9oxBSQHdwWg8LdcWcWznwlOXpgOVXG4MtS5
QYXGxD7SAvpRiUxPPSrjt5u6vO5P0tIrixM14IsUhlma3pQX6flzisC11t5pwJtf
sXj3XjvkOmCsnZaZ0y5oKtTVOIAgGdN/t5F/mdpGMLJt3hDQZXTyb4+3T/irkEu7
pXIbAwkQEhUe3ptJpjvJxk4ghItzqc7WKdv8sXqBwSxkQlXvkf74bI4Go0SmKndc
je4fDcV0V6fI8zBtnOEDN58XpBjxqFzwSmSdsXq83kB1mLXTPXyCMKIk9EW/6tiR
4U0bQFt4YVGDSJFynEyecCIlbHBQeJzd98/bBRi/LYxhS8igVlWQBBieokC+GJSa
da6tylQuYii+qUQm2B1GgArGUtzpIPdPoy8c5CC72UOsnjFCsjFkM/r71dNC2ZLz
sXOXm8MkZ8gwlw4si4BlS5i7D6zJeN77IaXoTHbrXVunkdXBI8URECFjV5Y/Ipy+
UytmrGFX4aklkyIOPakl264/BBzv3eNijd6B5yGE+1tDokEPNuSFAO6JwoAh/yEB
aXJydXcVBdIyB12jFy/LhRm+pa9eqts3jgxKE+153SYFouQTYT5Pkv9xVo3GA5VD
k2MyZMlIWtSa5cHWqTBA6uUuNef4wYgi0WsDsslMPTWceDAEwTkRhx/JVeg8HaxY
EHudGZrpXaazWUa36Jz+Z3DNEbLL/BDWNqX88ixUSjm9HLRmNBD650z7SfXksXYN
8rrwmOZrbnWthtsXB8vZIqD31Uv0ZmuxilXvkGJ3XCH07RceiYUPZUumzjpD9Urq
PTXXVxwFP/fdWz5m8cb5gCdDbrNlu5DQpLzQ7Wqrr/PPTXo2rTuV5xI6K31SjbdA
bS6due9Px+4NmK+VxjmOMMyI1RVoVn/CDfaCQpsyEfJVxnGjEdsyNh4jTXf7N4WG
3+0ulUHSDkkO/3iBy1SnNokKpf5074ClV2skFYK+TvgyGdZJs2cFxHZwIadf50VH
Qs+5nU8OASiU2uoLMww6F9muJuzZV0ZluwpCiceorfqJw2D2txrtnih/HB9tX0WP
d+xGoK553wgkw8F6mnhGAqw16oKvV3MGwZFutolfVuqjJUB25FJNwxB4FIvvY7LO
U0uwm00rWSBfTJw1UD+zbOCqRrZIIXEKdGvUoWgIaMXsVbT3qa/KIEEhEE5IxRDB
qytJhpFvUrMCYbk/6P9ZSZqCq00q764An4sHKo4ya5CEpo7F2qJbnivwghXw5iim
+eNA3MDN1otOdSRIzwhoNo6lR7QlOkB8VqnpovPtP063Z4VSHJ0/wWF8zja+pVaZ
Q3SrBGpm86aGj2ZaEkqcp4rYMcE72GSelcVNiflAJhHukLD86oXi+u4Tzbe+gJiA
pQoRsgdoAAmyaP4OP3fljTUxRu/hTE3LlQdS6luBGGeZzVH+CPRWN+96YuJ5HVOf
PBwd6btrXKDeGBl1kW01uQeiqiz/NA2lhCnhvIRqCR2emDDL3fjsj8wgI2bfoOPz
rfQidzb63Gxksab2t9Dd0NXsGDwkBYpdEdyXCMqUC9399BbhHJuko+A0y2rvokbE
eyXDkRno8cZsYh1s9fY4s64bDmnmajN7AL2KHLUmONjamv3a6uzYt6Z1vnh+jhJR
CJjtKoIYeaT9woLLNH9IWVdtNF0FlORU0f+8GxyTDN4oSz6ha7RQN9pAvpazi7Xl
8FkHghl40r9iPljLbSlZzMfacYZV2ygqMRgnSm0+EIEmVh03+kpjEHqZ+Gzkbvo0
Y9gzS1M8nxQN7qn9ibwI7P/QzFvoJpvbyERe2J0FJiEuMr4Lm3dzjeNwXhLBWR+v
Y3K8zwJbSZaDLJM4cw4dN0meLEkNVq3wWg0Cbn3ZVGQ8OWRl5NcmvHAa8DTyO+Xb
csWbPi4qFbJll9uVfekhZvtqi7a5Je5Hl//VgHNPansKDoIQjC21Vym2J2dzFjdJ
LcgAX5rNufphqe2l8yYnw5/NCYWPsKtB1OJsRiPNQSZFilR8xmPNQutquxV3XjoY
vPMlV8vCwY4aL+TSlKGUX5EVpWjMRAqH61dUEuPjkOUkfu2JSAiFHPn8vnubW7Bo
cLBRAuuyGr0RTbKOKa7/Ndg49cM+LS42MSgaULc20NA9y6TzI69OGOeTZREvehNj
dNZFL+uAOxlSekj8s4/vAg6oQHKS7FcMYD6IBrQgwndmIEagubhNm927OcjzStV7
HpFq8xQdwW4ArNiTwDGKA+3c2STNOm5ut71g2wXdEEaXAu4BMp+jiJTZODFg/lsy
k2zmWByXgTc632tsQYVfyM1jD+KR9Eapwm1tjz/Ge+zqUJYH9gQq0UNkIG/ozXzm
bxveGVS3Bzth0TUwapSNKaoSgrhbKhM8Ek8plDuHPWmNKsrkh7M+I4laiScRk0Aq
USyM6yDO9vMWO3TyaDIGcz970zT9AJUhLvAX9rOwXE1VrZU/PjOFdPftzeAr0X1N
h5Y8rWIQcTrjMd116GjT0XpmEZ2Fs8KHxxeOB83PYiiE+5NlYIDU5NPa+FrgqPnx
PxC348L4O5oi0d/SkyieHZIOnTdaRkPrBGLSq+t/unY6zlGITE2plOuHSsmvW/AS
KNRl652WXHcyOtKkNdjv5gWbZaavC+I6sBdIAwc9fzRREqLkanLf4xB2qHoxbkFu
yx+T5+klI7QHFHZX7s+zTFxcd9OyMF/2vwYE6Midz3CTL89fZqeu0NWhf6ha/Yyy
pbl5fL25+fjRPFHTPaaUAKL/fHUUF6TKrSQAeTfC/w1IovzCpLEqEVZb0FSfAf5n
//0UssYfVaFlcrQ7dF3XaGGKQmDJcxgv1k78icu06R5kCOdT/xmVGy4MSjXy/Nfy
x6uHjWM+ZYzgkB7KrCDUMvYnTxkCV28p/rcB3FFt9x5MjJf1mq5n/UKE237Kd62t
/SMjBcgaHcLuEGna2UMg38B1sEQ7BsaQcIAxvNkQSh6gNpYnqt8/eTgM75pV0rpT
iOcEdxNd8WQMbvJfTTqDtoD1kfkjuGxOt7uF2A33DELAw5Ss7gy9bfB+DmNdx3vj
tQ3F16mgT59y8/ILNE5dtA9dNvOO+7vDndGJmUb3SyAZTnpoyNngyX11zS64TgZI
KThFAcVIVEnUDMEIWjTgvptNu5FBd4GyEtgB9EKzli9rTiFYSwPL42uowtwpJk57
b0vAp3amd1LeJUw+WCe7/PiyrypKReS6ZrtWsp3aVH+G9Na2QAgj8b4gcGkbSWrb
7u74G36uSGuXZ+GlA7t8xKWqfy0lizNYoZEZ0Snz1WSAULp9ZieNjZcsVn+U9/8s
BCNb0uZeTTO4hf3KPBD34ZnXZunOuhrKIkwndj7E7msiDR9FrX9fK4w25m83FIyl
tE2TFWELn+3t1p3fDNK/VMRJhiRmJLEJDDpXRdXd4BztTT5TA+3G4HGgfxvDWeOz
4waQ3xkVQ/gZ03ab2g0PEqoGlUMjY/sX/ziA9IPHGymmKvOqViEqk6jbPY++AAWN
KL+nJbl27G4RqFW4Mk7bmdH4wozEOuqrGCQV6MeFaKMPzOCjnG35y3v0zPa0I7aB
+suMkH3FoNldx+ssN95XooX8CzNbG9ba1Oj38WuuKV7Eh9nUpAYrdgrunDZTNqOk
t/4+r+jP16MqbYg82cXSgGchWXOPxQaO5owaG9HKh8J5fItJT6fECvsxxFh3N5Ka
om4s7oWfifktQ2WQL7kpnsze8iDNFm+i7AmMDsxjDYFiLPpUOFby5Bop+atiOJl0
LEKlp0bM7Jp+H6HAKFQMHtMhNVp0GJCUmU7Lfck6kAkiFodRiNKy78gtvUolyxNx
Fz4jDGt+pa5wSrrUuSOj7F124ZOxRFCECc5TuwXjAS9QL06p82Ad+xYpJCmqVf90
/NvohtdOg8Hlc6chUG6KHeZgXz29XtBTNcrNUBWG5OrpE0rvbGkJ2qepJ5oMVIRs
qy4M/iSO7IX59i4R8lfDar4IfSyzMn0dvn8PWEGxj/iv4MZ5gnyqmbJcManvo6BB
aFsUVzyxQM4zDzB+soqqP8d1oCLvbhQQ+TXb61p3PJinBIliVH1o9cXh7tZyvy3i
PMmsuo0J85w3T2rHPSaQkHcxVvd7tVOs/soqLhhBCU9PmuA9SI/AYFtFj/yVcbDx
uL2MyQaMywCpAZs8IO657sSZUmYA5TVL2VWx+naPXf4kV94VHS+LEowybVJW4ch0
kVnlesG5gBNLNt+VbVRSVapDoqeX4A9zqmBZD18Bfsd4M92bRw7SDpGr+Dyze+TK
PefSOy4kd1e+JYf9Nr/fKxTqKgAOUsDXZ54Tc2yrTdErvXCvHmMoDE2s7j4Gat8I
vBDXNyL3/1qu5rzcg8brGVwFvJyfCmhHNfmKfnLZMHaLddIuhFrA7gtXXP6FLyDP
QZDLCUmUu0bYTVXric09WMm0vyttYp6JYF3xaN8SspU1IWvQ3KAOdJwaUFBMVBH6
TBqT+d6ykpezztbu1Isw7HFrQXxM+N7uXjsyrnguYpwt78jhcPi/3xxK5V1e2fwP
J46zkx4MdYz2+/NP+r4ZRvz0uiFLE7oaKtNeUZzVMI6ixl47lhGNfvsphxnFvWe9
lokqGzg6JQDjPkRFL3+nWDJ59uhU5t+M4FAIoRFLxHxeBDT7lGtfXv24BwfM8FMD
bEmLLwqqkKuGnZ9I7yE0gWTWEjTFZzc3oynTwLWGSPqIUckSqfAB/kB+emFFFrcc
6DxgwrSCZlTj00iIDTUJqY8AKTMBZNLgEswNwJBn24YaNHhL9D2s4nIZnN0u00Hr
Zh0z4NcWQa65IL3F6+llpfbjJpLcoC5+yvXBzzEGWwsrA06Gt0ZFK7jI6CU0h346
gJnbEKzNP5C4AT+VjKilxVGA3S7ekkOLF/JFgllB3gC9OUXoGNVogx9qOQxqPISf
P0bPUcVQMEOdq8QGOJvX19aCLycizVZHzqqWWRDKHe7jvnhPxnudH0AfGt4qKr+E
g0emSGntFrzfj9S7iQMG9MJbQJVotPEo99mJYzBTEVzLNZS+isaBlB3ncvp9P+59
MvG7hnL4S1HXO+yTyJY5UFSWE7CgcLtE49m1a+RAZFwVPLjfe9Jxyhr4osrm1yA9
3tkyX+jNKlXgkTC44wTOrMSWqcfJ24wDpuHTH/qyjK0Rw6EbVkfSYM+bWtCvGSJO
FM3HEprwqNVi0Uo9YnFuKrLnzX7N+RpEjB1M8v0V19pBhkZDgyqaBgBsvI/vVQKo
xuyC0GIGF6Bdx88gteznN2oHDiEZpOQKQbPNjouVyFhXm4KekFzCOA7d8OJCuBOp
jpeoXGrlvuyNDfSvMg8pa8OWKkyLEYQUbn2lB0r1RMtJRn1QBUvR234IIOyL35Hm
OUtWdJer7IAGIVGleo1nJirSy3Y1Om9rMIwr2vCV3LyJDeLR+ect1bsB/8WK0+AU
qcfrKh18K9AkUtLmLybpITmuxPb935oLN+nOJ0u9TNePzb0er5KfTNZVq7y+I2xy
Xo6VfkmtGmU1KXN4lZIR4GowNi5BKG5jmZc9RQJEd8CsXmq1b8wHtSPmg3SVhtNZ
vDOOdhhlZv1PlgTQR+U74ZPbq5eOsg/1UYUbl5mKj+ZohULWrowWYHZJcZPltZA1
rO9zBy64PgpoAGGJ3cDTHANEotyuK6t3/uBxnvMKAt2BbbYZ6eiBSuxoQHHhHP7n
1PPbX4RGKFVruKpSUHJlKepxraEg6LSOwJzjOFyL+ivc3o+3CvVNu/m+tl7upTSk
xDmrtPsKM3iANzPTcTfSo9cmUpRvH9mx4r8f2MrKhkpOLtM/vQ71Gm7vtaqTkeTy
ErwdInFIUZtTiE/GpQUoxXXeP0b2qWD44K8feGW35VWn2Q2WpnuxPL1ycnEAtfrs
kva2xixyUHtf3Y7nnPO1NWq+ozudvt7yf0y4wcx8AavpOH/cek6Pm4zjLFr3t/JU
3FKLB8EDVNEQw1wEJsbQMkgOgx5425OzL42pAV5B7hgFeJcq+SXZo89mftb3Xvso
Yw0jNMP597IjA05R7hVSdcGgCxmqnTIBG0L5mxwosAcTGs3qKr2aMDBWMEtGsHQ2
o4FRtkPm2iUA/6ujKAqqymvczNG8HA1LbFNIDO6+5ZSu4iJCWuJ1o7B4zv4ORi1k
eDVLd5WXQSvIyhEa+CWX1X4cPcA785YuvlaGZE9fAgSHZ7s8mJ+AkIKlnRNl4WSg
9jFVvV14eh+U0T6coE8zCdXUxBuOV1AD8yR8YstaNeA9/H9Y3UFi/Z8HXX3wOPEl
nQ0J8870Wm+V1Z0/yhERxF7YJa4Je3M4Yky5+CyhqtS9HYO4crFndjT6nm7P/O0K
Pmq60ye3LtxtmGAu8XXrcwZAvx8f7G905WQ0dujYgKwbjCuKU4nXwDsFx82jqPMU
rC2iRyqgN0llp9JRyJxhQxrUl4icyFD6WJNpmaJgsCazYFIWhR0WFW9QyaIHYzbk
qKZ51Tf+hxFFaSd5fuRTZPq2lnbNQ42svatLcVnHOLdFIlTp18u/fgakNJN9M2fv
39Qi84LSucSEJHaEwQhBcYa20eOb6ZO3RjmRuHq1S9FLl/R3bOgjTwNwkV4+BHDB
DpruMaz6sd3n4dMGex10s6jOMMmmh4aew2ew/eNMptJt7EH1HesD93f5v5xml9fl
Wl+2ujsH44qoRRrSaB/oUIKanf2NA0ShGa2fJ3XeSBpfH6aOeT1ogy45gX1lXmDj
0/ZZfA2CGAeZlToxxTFnk6sfOjuMyIZ4JnkEkX5bD0NWywLOnldRJLLjVTw2uRI9
lZcpATHLP9UREid84KsPoEv+XpK++Bnpuz7PNZTLTx7GmkDlyJSKSPvoOq/HcVBZ
beBzdVbvMf99rE38us1T37yOZEv7FkLTnkCJskPg5TJwcGl/EvxiFoxPUGEv8Zy0
HsykxrwYX6eLDHUxBkOG6oycED21Rt5zIfjnWtEhT/KYlIknEb/hQkcSXAoz13LV
i44tdZYn9tcWyLZNTqbJuQdqpmgxPEMsLmg53EdONdR9Z6Qp779tAok64oEpgrJc
zyurJAhAVJyla+cWUvSvrNv723w2WDKfR/EQE7ubAy16HkgAXllxAIj+5EppPY1m
zxyJiTPWd7xmuLxeJyEtCfThsFEZdCmvugwmjT58+bq7jGQPlm0kka7NnreDv/3w
cRGNFP5T/CFJWNyQDLH1cXvAKTDKiVrL+A0/D1+12TO2G5P2MRmK25GwK2BXcfsi
08PmUfwEh9hX+oQNZeAReZV3UQYdZu0CfJB2UsBx8jTcwheVoxfEwa1w3OuIZFUh
dk/8AaRd3GjbMgHmWE5KihAT9pFR8e9QDQWizVfMw42CYpsQyAK9YYFlvIflGQ9g
WiN3e0orkGBXngyANDUVDG9yhJYh9D65VH5C4SwF0/VcKdKEMlg+xsFwD9nIYGaP
MwVnpGs+0K88D8wtw+O3/k03X/8Ojy89VOWX3uHqJdFWC1sfQ4QADcyDFhzUrYox
mqaj7WUNaDZ67MwBzmaA9bGc9gOY1t5Ibi6/MyPDwRq8DlFHFreoGNrLAYKi0upc
gYzgrvppIIBTNEsncnpUf/OeGI7R8aDCY2bMxxSjmXCJwI65WAgI0o+28IUy43Fq
w+dPxokxzSdiRnnDSCK8+TGd9T1amrPr2/rpvLjHhQR9Q2l3KHOmv7IjJ3VAavRG
1nha0aAO87YlQWKfIOwjyT/akt/CTvIOR3tT2HgqKrJMPFPl/SWnRZ0d8LyMqbFi
Q0aM6Ex5Cbm4neJvIxyDwp55pP/8SgffIdPNcbNQtg55MYIzs9e17i4jt+6FpxMc
GH+wm+NIBZuq3TB+ItY2nJMLDSlCYjBvRJUErTMYL31oBOxbBpdWNQ4u2XzUJH41
2jpNJx7d1V8sGkDpeNBIN7WQExeLlHhOke0Od/w5eOXL2I/gLs1Fl8xAzyv5KDtq
6SOIxz3yhizwemTJuMEr7NNQq6RC+cvEyQxzy5N7AMFerqtiL63wHr8o3x2IAwwT
nAMuZDFPJ52nmV1D+ciJu3IL/ds9QTs9no+Pg3l6RYUnsqEBj75/HfYMElXPkw5J
4Z5y/XKrvE68QwotMBITbG6IiKuCV59eS6YMAu0Mb2QSNylzethaDAxRG+oQH9rW
wuVsX1+jXLNFr6gfsbRg8DkQ8THtu4zBdd9W8iqjQczDJ3FdAfMiM4kWFMXTrlLW
Wl/r0sVNLhfxYArwvc/+HwFgy0EVM5Cp0JWE2mFYE+dk7hkCkky9XTeUNYSrAwR4
PUBR1wmn2pMh/c6SnuBq4jFW1VdTD/QqTApEDQLhCbB2hIM7iTChlDpcN0dpdrt/
G2D2xYnuEO5ioRdduVPYFtKu2+xQjCPlAoXkNtgHHWBC6DXL0vixy0sbLtEr7+T3
cOZZmxXBIUTfSZ71ECqVx3eWWNhike8glKi8QJf0j1aY+l1ERiglAsmkwe4gQmHI
9yC65fVSeWk7qbsIA051Hj7mifgPYMH+Uhj2nMjRZDJJ0q5fH408G3W1TmtBaSJN
Eq9Xcrym9ewIIN24TGigZbTn4P5oPFACUXpr2APAqGNowLaI5P+yp4431FDuFy0+
nWLCPSGFPYBUjgoo7o0yq0X/fteiZHnqBsyhLnr1D//qvdS4lv9FTj4c61LQRbpE
ARmpChqpJjpy1t/cNVYP8ix5EB5MSfw8L921t8lBls1nWkqDFGFoWx8owuhyaAPn
9SV4I86zy4TZ5uZBPNS7203eBTbv02HZqzGP9F8DjX1UMqXmC95R60UeSqzjNkND
Y139/3C0U9xo3oTYMxWIZKTQYl8fASER2PNRydI8ALYJ4XsnZoW3DQL7MIHrPA8z
6D8D6JyGO1IctZeW4R9ztbu474520Z8p3OL25KPwsxPJYlEkGBUm6Bkka8PUGEU8
Yy/BgOAtAkgkn1Tt00gkD8J+uLeEEalOcIaelMDzAEgahD47fdjRK6Ow2rIFttuG
cqEcpNAjiPMLwKs61/UvQLzaCqem8VfkPuYWnhp8Vz5mDRmJSSaym7Qu1nxMIp5R
qJqHlTr7E4kn30G0Sd/vEoumz27fhouvZc6m3r40DJmlUxXyTChp4LSqtWgRZEmf
XjOeZGTlQjkTcrkpeOXvGwQGAsrXEAZ9EpGvWlgtO2RpOMMWH6rVjuMwjUENa/xe
HnW3gw5IAkO/Dme8PjRvSXdcyNzf+ox+I93dlhEt71OHQullxYWM+IY59ujXf7jS
3WHNVm/n4oWmByL5s/wOPjWWzFWWuARSfWRqSshJhq8bJ6fgqy4JCZz4JcM/md4U
SD6b+zjIVv1tkHrwajAT5qIFiiJz+emp3Pmtbj42cZAvePoPaF5j7XDh3Yxn7cBH
jNJS052XjPNerzSyKgdlJTLJiqk9BRMOd7yXY7TeFv5QbX20BvN8klzTgnQKpePt
xsloGJi1GNNHTtdMMtPA5bjMd89K5wLcOepMq8yQeA7kYTVtSaWLkVy+hxcxQAGx
ScqzsKbC4Ju5iajAhsN39+7rBS4nPK6kIhvuj3WM3TvU4JAOCEv6wBIMCmwO9o/x
Gl3APNt7io7TePst1lgRYPZwbU6zJKD+G3cA7AaYBr9Qv7pFyy9yOEVw7dBBwL20
vQVS0+IHXdaNsfbUzWd1r8Ex5VGSdThN83Scxbs8Zq8BOac594c8YuPzkvczKsv8
AuO/5NaBE0/TQGl8kftUFTawrXgw+BsZ/mcOZ55wg7YEzjNTh7gef5OprG8LM+ek
+NSwPbc+YZK7JnRUAzMKf0Qw5AKz86792XCX7gCRk3AvaeKxeg3LiTVcQJya1atw
kdifxHW6JeD2awxocoyrDI/vtflQao94rYhq8WVlYVzgogRy05+R5TPoWrF6zPro
Vkatf4qbIj8i9KY8sNvPINE/3fm/vSsiUcUa5FeP1Mm8sVkCYneT688AwChXH/nx
d+re3HarhYZouEnp3KD2TKSBTlMrjiDohuQR0I7cvF03djSbj7MtbSOCDBkHxtkR
our++NzdMHuKHmBSelNvUhsOBEc38BPfrdAuryp//U4OFqctAroM38cuB09Sr4uX
NitE8k+rN065KqgWT7C1xpVd3oPSkBwwwvf/djV+PvjkLEJ0jXDPFuB2PNE4rZed
ME1U9N2jMWMxYqarUrIY3TErXoCQOXz1LeMw6wDG7KDcczKjYd2ZehB0CxJWvBhY
PMfL8QQFFgQxihGgmivu2ysEiC1rCkgoF3sgwrvjOm3ZQReWcBbT3X7/Qys4nCTk
XEFFtz60emltRGt9WXQorEvYdUUiFSi0sGwMXCqbePi6u5mNcSEtppbWKUA5uy0U
jsgBJ50tmeuKDuALJbz8egHuG1gSQ7e+yjhviryCLNicMKGuq/jkAiczeRkKWkoQ
IpU1USws11Aw2YFHVnnegUn9+wlVdWl8/gX/JzcYB033kwnmIgTOm9zYPW+X35uH
TlEC5/YVF652P76gqr6I9aqFbmmI4McF1htrEsFyvapFUndNnuOUFQ5Vo95w+Aks
CHCuVHu7OFH8cwfiOjUC2wkXyNU5ReLF/6oUMilhP9jZ7DuVuTDQuuUQlPu1+x1o
8GEmaQsuIICEUomwqM0IEpRl9DAKfRbWNcQgKuLOAmQ1pywMOZWz8MnrqnHILRlL
5xMA0UO1IwZl8MBDze2XyjcLWdRIb891UQHfdcEttiy8MImfKFNCuqIDbVBGgi1K
MgSnZ/WDha52vB3g8BEmS98r2SDgwdH2lkvgajEcU7fbNmHnA2napTQhA2y3WgmH
hJKsHxrexX2hSIL+YC/1A5XpYAgUzi2nlPHvQuuRpRl0Z7FkNvmcut5cDT6gFb2U
dXLKCS9uzDhTG24Bd6JBjEjrtC/RhwXFJ9h71VtjweY9bx9PkSJujRcP7GoXkqgi
1VzPPdIu3kzScddeOwngth6b/mM1Wza44H9RKGQwoBhOCSYeE7K/7Vh9j/si7FuK
FL7TGEAJH5vxGD+ZZayfTfXgghKqnsy42sWACuI7qgVpqy6oNs6gdxGdoGVgGsMM
/QKEP0ue5JcusaoEKakDdgqxEL2dmNaBxdrtzersjJXo8Ekgpm44PzOhKOTCw9Pw
jJ1wBpdajoqB1yS13sonFknrWN2aMHcfymD9JbbOD554pGTvrFp6QBJYVWIZnzGt
fM90tcrBBa5IleG9CPkTS8b7SlxCPq/yZuQzeVJwOxW/ifxhaAFONex38XizIQRv
jQvuv/JXlG0/fM40tSuS/WTQXJC9X9pwJbHE7NgGISXR+cNx1j/HkjKQBi5SXudH
h2UPGgW9Z/fPY5PqkGBLcMX2Ms8Cbkl2vKijXvVGonUtVxIxtOFn5gO0/bDqFkrE
Io1wgGjNNVzDTOGqKh4FwWp1Lzv4OPa3cz6ndJAG8QNV1nSZXdYv1chlCZOXtfA2
ohK/W6FMCyBvjSAmv3hAHNPPc90AiytFDgER+8oI1pB5B2bBt62k7qUFTSNFqgRt
87ASSr0ZB+LDEKWECpic17z0NenqH6HsP07bFujnqQ0OJLUGZPH+zEwjCBADPgwp
hbdzSXjqM9HJbc0gqKtF9ty4oNCIJ3B2TmetSjMWOuMeyGlQNcvrIG/eDIbbCsG+
QWXz19hK1eYpd04mJrB1AitKt7e8P3duyVdCWvZXgXCX1i7HVvuPwGcNO0QXkEE1
uqouBSqdQpxyl39gGa4ALrrpOZRlyODb1xvAjmOhkzHyvp3NSFn7Niacow6jrrQ/
uBEaFAaD6z/lzA/nZx96As+tySYkhajUGGStrlfN6ChFMKCwvSW6SZvthaWKJqh4
fLOYFw61zcEs9zIBI9dD3DA6VueIblOFN6xs+Cz8G+7vp5u7SPha2n1vNi/qy4jD
rH6UABlu2uzrc30+qQuPeuY05LLBFd7ONgHKpW4jTRpcNyHXPtfc+Xdg8tj8S7FW
PIVDxDl+EdZksk9KZCFE/ZSBMaLXR+kT8OX6RkwApvPEOo33iqZ7kjTijwqt24Oi
1C5AfUZzY0+rOzC6+IXobJ/PnQXAuXT+H+0gFWD0+/x4mkNGS3VcRLXp2g3LZ4X+
YooWkOAiVQu9sb4UA4+TM+peWldeeHpA2w1eRrnniMOHm5IDf8VVot/t1qH5jJps
Vokzw+M+W/squR4YOOWUnJU3tTdXBWtaIUa6FGzWhEpxjHATvW8K+LyKcV6Dhfm5
V36p9S43zP89QbG+N8lfwcWLb4sfu6y10b3zuNDEiGeVOsMldjjbf4n/vPWTf2Ot
bDqyXwxRqhhXi4t/9OARE0w+ge7+XRe5QF/A8qSmEceCRSNQj/2vTuctzNPYliZ5
Ow51BBKPKFQTq3CTbEQB7tYH3HIp+l0fCx0OVHc1rjkwLt6RJUpkjJEQOg8yASWO
OlS+Z91DA/ICibkj3qzRhX5YvyyqbAH7G0BljbFiLUXlOT+Zu0HVAUTnEHL3gjtL
KU5eh3fWM+I8cezDneAEP1n2q+38G1BjySxJPYX7wtsCIFH3k07fHPHvsAfGGUA9
t5FFQf0+dJ3L4bR1Bj1d3jMNO9ok0xMg1wzTFrL5UWpnFTcnhNti4x+rf8TcF5D0
5utnYdwfm/ufzcbdO3BW8DproYwLj7b/4XT9khl7oACXgNZFlDUSyVNlL7eA1C2s
iLq6JHz16G1IkezLiswq4y5YmGDyvSa3PuO1Mz77KKoujq5kQwe4FADcSGNLsVcO
A3T0HMz87I/6vj5qtpivJqmCy4JSrL6wb1eFl7EehV/FvOs52ysS5+HscSwqsiw9
zUv2/xQ2i0VoVul9IZI1Y8ZT7p0rZmXJSfh3nbrwW8/JCjKTyO6lWkkvycci08Re
nVqOkCOV8WHks0y54SUkP8yCO9+WZYs86emcGFF1thmtZwlijt0IdGw18VbIAzXl
VFXQdHLSmqS8YXdiRyu3mBLXSPkmjwPnXykB1a+c4IoT5dtZavm8LEPrJ62G/6eP
rtF3EAxn6PeiM0UAjpNcIzzvaPa+zExq+njyR5FvdLb6lI8CdbSEngDLLYAphpRH
tE3rVR/mkXqWwDC5Pni0soYN0RDKkoGBOuiFlY6SDO4TuOWA/PCTpClPR9oHxnfF
YLrJgQpWiZPE4awahIM46PC6P3umiEn+5IowJWceOaaFLPS/rNLZD+GPB6MOGjDz
aEszpGaLS5JiX/i0jn56LKE5eFidAD2odK7FBfOpUO6hkqCwDDwuhmsUCu+d1SYS
YI4O2oXQRU4SOHITsprm9MpWcaRNfwDgwFI5JZspvrrpo3ShDROhkjwukMn4hgQ5
bKRVJEYX05Xub9IoOHVL3UnMp5R9fb45JpYcTnP4QSxtoEyAcX8W8hqhZJT7QnwW
bdQXjRY0DpJAiSVvE10bwoeiC8BhpHQhBd/8cyXQZMoiZpuVcWvcLTz5mpv0smme
pE6cBz3zWnqISCIjhPa78WWfaV2SbtyOGMPB7cfMyynBHrB3bP1VBJAviEp+4//u
+TDuf0PO0Nx5HV62wjnIXV3i7eQfHqRO8hVxJJ9ldN/4DoywjRvYyGhMkIbllQsD
fBr1F0MQCy+Lw8ncg75EGSwktkOg/S/Qq1xUAJC1s8BRVGb+ExZSTuFZZihlRcGD
Aqk0ob0ZYqFHy67m/E2dZ6QAk5uLXkxY6/ntPDi98ToRWkQGso5MF/iBJcN/YZIh
cbGrtuPxHt3rGAn6pKfKihzb0D0Vy6ty3eFeOu0P0YdtBiOZG96DeKHzHbYmvEAR
r2gLdqMd8CikTp6rBTPkr21IiZlsqPGv65RzLLwSDjKMS/GSRfAAz/aT4Ios4WfP
toeYbHO8bW4G9F+Y/dvxAnCe9Yx/fT3WH6T4QvLrIc4wKu41eD90wt9/R1LuLLeD
6qao1QVkx4u3qyDyw+oEpL/lzfNf67H16XMGG1rk2OMJ+ZMMMArccr/DPmnBHOLe
8usTjSW0eaA1Mvkn5MGTTg12RZUVcRzTJzyEH8moYCmVdUjvOKMaaAUht7gLhqda
4EhSbrCsD9LIbQj8kB/Wg1+6cZPL69pDXMWebxOWVIi2cBjhWoUeZJSz3yRI2gmk
4O4zT6yadPbwPjtW5lnV9QxWxVDzXeBz4x5w0JIBrVgpIHdV2BLraeq4oFSZu4Nv
PaTLVLjbhgvVWVi4/HPWkz6CxFiaBdU7mV6mKTSpS1hmf7F3CdmAfbHBXId9Na/C
rBFGItYvebGRfVnzgMMWNWssamzFXu0U71xb8ayaHPIw2OmHcUZ+Nmu3xjqBYTSd
VT8DL7rHRXowyntmHC1MjtTAmqqp3vGx0dj0hve210RWwFmvqvY39+kbhw9jqGRs
X5VQbYi8DyFOF0GaqZ/3rtRpdkAgRDFTnOUtLwk3RqKuxeF2xSNzQYsjCTRrePsD
LcRP2GGzDN5BRdMW2IRwZAuHIssHCRw8GCGPtBYIDyiPVm/qegKa4ORcBzSBajeJ
UuRMPLeApf6CBPJlrXnFUhLlOOC5nSLFSRQjV4t/My9uTD/i5lcqzEagoG3KVlMq
TYawVt1JXjp7cezTdbJtVEJD87J5b2JeF2DdqLe31LCX6/Bnt5vFgdca7Tf1J+l1
IQMLm44EgIF62u1t3sCuZVaGQFpvs5hIEjUDbVl1BRumv7jQ7fv/x60eVGZ2jZL9
wyhaajblq2Y9PmY0S9i5pzBRbeMfDLUYhuvy8dPUU3bPTrDJ63OE7qD1PhxN1bot
xptU1vMf166iM4atagsOltivJu7zX9PpF3zJe0RTli2GOhAE7MbwRQY7X1acx0WJ
gyEAU8KTctUMh+eZsU2rMfzWBv+YrbSE3nm/2Lfe9eezKsohvcpelS9NfzFjz00N
EJwH6oDUIGOAyomdGvB7djEkvacdyRNtdYBJES3kBHcXkqZW1qRqiLgTfGkohSzZ
49P1qfe+Ta8uztHUrQsMB7uFKnmpOQaqXwKXcryY4bmtu1ZcqLXJ1dscYndRs12p
LVnqYmHjr9c3t7k76J/O+SgS2lCDlyICpeMU8qiNyuXheenZWm1uhOK4Fhpe6hqn
TyMvsmad1wtEQfCEk6o7NmSMYSQXIZGnFHDteHvWeawXiCSfUlwAOAtC8YFiG1FI
3UDq1xL3uexazfFZQMHYACuimAZqFnaHHkzlI4itogI9MRoxKgMEnoYmCWShjrsp
VJozz1nQktFiRNILMr3yYIf0403lPavjANZoY1h6it8mX8xzfr1NrmcRBLX9fF6a
z+S/t9T92L4xJqeGKovBKfw9R7a0iQ1236CpiFGNjGTRKa/aIZPD9i36kUJWchLJ
zHsIjKNRl6XgeKkvULO9u33tJTMWZw3y/ZWogLU9skZRKXo9kobMwR9T2/ijZoSj
Xv6dqCPKvt4+uJO8+yAwTZCLMTiI5wGXrBx1n4gxgImYV3zYC/z8FP9JihNhn32r
uVWfu0KEGXr2vR9ezQdhaIsQudGRYB1nCBWSn5cclQ4GT/g0d8mNcg9Dk0IdrRy0
H7KEj41zk+x+VTOOVzSOHI/+f5NouSWajYaBFNdtudcUwexZ9/QzHBijXueYnmVe
zirDVVuL/w9lUHUVECt5ZZPaX2DbJJcocClfBpKtF/OmBmK7OKNq4yT7xPsD9UUq
LO2aGVTf1Hp0uUUmMLDxUdT6MKfsrHi+mZZ4pceFkDEVy7sJXe0Q4sP8RXi8VIl2
02ZHdSiX54WzhIit3/lDLZWnk5H/jcSAuQUjeiFUzRwpsapHCfYOxPDWRXyK9xid
tFSIZdxPwm2/BMqRTBZSHkYJy4WDDRE1ci4SfadMwIZ9BG/i3xLxGb1B+XFOtK5v
hiL6LBVfpgsV8wpTO/M4BmxuFCAHzN1yNDXN6+4UaxNSIHStWMgHHwh/w3FqsaE9
1uAsxxvkxHpvnJMHJhGDcjIFZ1p2GhomsWSgA0qBiQm0t5GCYp64+JnGucxqOKN4
clk9m/xCS45/SZNJCilfIORzZMg0BrxDTCpf62XocfihENo7bbkrBOETj5uobLFt
l1eDQsnbTFi7OrXt8l9H9+QsrU7pBqsID93RkMuP+oetZ6AzMyQ9LpOcyFmCOZdV
Dmil6Eq+LhBVlEHzA8e2FSuakJ2rPRFUl+BPFB3nk7YD0z3VplNimCI9ZYT/Q7TY
/Mi21EM4h0bsRgltvY2jNy/S8oJmVjbRxJFoNfIXZiF3yKhXloh4RHDdlXnlqAym
ukiGyiDY6O5BdYsKn6ijmr62pH7DinFOpbBAzHexFRBPwQJbWHmAq/Kx8LS5/bZR
Jv+BjzAm0FMgLjLEKLhf+gyozaftJCATDzYTqnRU35rflgrRKpf246q+/XpQF2WK
1OHemE/ea/mP/bqFBtagKF4QJ9+Yo1JnmWsS1wifkPBqLxfMMiqtv9NKvfYrJtuF
90mCIkkIldxgrw8WBG7nje9mDVeUXxfbtgGLUYkjC4+Lw7R5itw1JQ5VOPsEXTJi
4ml8qC0iJoEy17r88BK/i1zcUab4OIfa1oetDTprT22QEVaLaaAM0d5y/1Tmes9Z
+joAUzhrezj5gSqlRJH9scrYTJNSbWNtCQ/k2rRdqHYaQsQXDVgUJHl2Lsus38VE
z2smJMMtL1EL4223xm6Ky0Bof/P4k+V6LojiqC3l2f3Hp5txaxthwk39+3iUyhai
ueuTHFTBdwlmZoWI5j/7tbzYHXY/ZS+vAHj1voFFWTn9bUtmjMMhXNRR0ZX0bBtT
z90xYD5Hz0X5S9JmZ/GMJBFLnJDuIiJ169IHI91H+09lMSE7SbcW5omAdizz/y0Q
223rcHqja649xQqslccssTK8OrApbkYFoVJjhpZwvhYNmZc0UlGBAU4HmuV8z9r4
y0LI+Nrv3ZvpSeWD86dp98f23TvxIA6/s/Wq4/UXCb51DYyaXWJDEDQxliNt2fso
KJLGypvbzOFwzNxh9Kiw9F0pbzUc6zStOr1I4TkmAFO7XQYyThYGLveGbCWQ2pY2
ZZX+O/dAdo0RcUddu8Y1+ZXNwMnFU0wVkmc5AZWx/76kqTny2199Ke1QUzTpqiFy
frLACsKTjhOSqL/SaSsWV2qoiZQVDPce5/UVcRPAU6PszhUOWfDk4HpSG4tqmaZ7
MtPsQOwAoVoMOcoQM89e8LjE0zOuJ1mYw8KC2dvxG3o9Oq8/Tkwe2CKOQbvQ95Q1
CTdsVT9PqHAY5F+XDo5CaE+SUhG0aJzRZMliYvTdtQQs2Fgj3oAU/6thkO+5pvJc
jQTrfKWQqOoSAxG/kD8LmAuSVNxSt9UaT4GxWF2JK4+Z2TMMfHcU3RIFZSKZR1Sh
f0IsAHLBoH0wihCFfAooG9v53TjHyHPRDIRMPrMc+3SElKMsc+6+vdjkwz9a1t3a
cRp2vh4GatAwfrj+xOUw2sjY3RUoCZLNuzeeRM8QDuQw+Ke/03XxFGVr/zOW53qD
pQBW6dSzSj1WeFYdnANl9KpljHgkQ7WbH5piJfdZKQEZihWqKtCT9Bi53WdDwbN3
nvanzdcUY2evsqUeTp8lsHHi+fzBTjLN+7icBdwvHL0dIbcWcZxtDeegYQZJnUZF
wl8CrnG05eSUkXKtvP4tMGootiu9F5UkCiWptf9ry32X6Jn6Q9pDw2vlCiYyzJd4
g1JbJ3ubHCmRDk+UMKHqQMAaVrDJJEHU3K9lkVp6/yBq/L/HVrnvIbf9dsrqa4aA
26qYczfzShmDoq3gh0jS0lDN4tS4CDv04AotICbAc3Y2BTovgPYhkvKAJ6S5AVYw
YnyPwQyj64GD7MKTUqs1/JowCEz8LiwdA7JvgmAp4cpP6kBZ+GJ/1YaYOAW+U1Ym
ecLdvEAoSCxliocBoRwPZSBnQAqTGvzS5EEWbWYYfEcTWWemrR7uqeeReQhUeTSh
FkSwLmvr/PNqUSo46hkPcu7jmIbsW7p0ABOs0dAaq5xQgw3OxDuSt4SRnTRFBw0k
JLZEjpNWqqqBH/hl0vPZi6f1wW1UoeHXtFsl3TZvJiMZ2lIWe90QN+mRcBpKayKU
FwtMB0zIuL7ppOfrucmUUgOOD+ObeHxo+WJCpouu796psMQpMZ8zT2w+LbAKrr6u
kcrbQoTjrZ8DqB/8oZWV4etfLqEmP6IXqXB70DLY2pNccf3PLh5PPNo7Jcfq95Pu
NR7kLR1OPANhK2fdLq7a3NVteChmrC4A7lZH5WvsXKBw2uv/SKpGYUAMdoY6VEY7
ZiuZ26Za33Y2OgsJ/eUouNqTxsLScE9QgunVhBzYQqxImF64WbG8NlnyaQ57bHtf
3U6orYzKSPbovXVMcIw/he3fYAoG0qC/pFXRi2GvGLE2whFi/V2v9XnhSAfo7Yf5
Umc9V55mBDbgmSrQwbJoRIQk/dmvjgmKRuNU6Antr7YzgWIltf4waFKdA5QYIbC+
hu1Jmdja7EjWESJd+PBgBG2bJLN6jSZUVU+/XLkzsJXMS3tna3t5mfjryQInDYtd
mhpSPniqOKEYalWL3jpZ0jfzzuGB3uvIQgFp/6PIS9SP+7158cnR3f5qQ83c8TME
11Odmz5s5IJ4XxdzcfFtddvcOw79P1t9iodUGvnroMLdOvJQhYPQq2o2WZi3SYB5
DDY+dUPwaygU82eqQdDQRsO+QyvknvZU1qDSmMa6IkECe63kYUKiLg7gINGvBY4+
r3h2wdm0Z2xpaVV/8S/GAxa5lP07VcSUfZ1Xs6YdeYS5MX86vpbGkEobGwhsYFUE
O3jL6H2jgiWlEen8D4Tkb2xY0gHQDx/hoTcbzRfeyKUIx0ZFRkQ7+UPw2lnqE+op
1opR6GSh3g8ljbpuNKlgs3SQjpYNupavj5wXnDQEaMS7Jg6WeiDOXt9WbGba8MiB
uGRQibOqAo1rYV9B9Pfcl+v3NWzbOpuf3xtuwnIWflUtWskRi7TmTbCZ/8ZFQM5y
mYn4GnnCIpvYek2b6yx6ulfXZszZLp7nn+EnLss5pjPu/M3/zWvLrSVC/lqYjx1s
vKxzcikPO9ghMmD3ziqB3dizGLSdSVAuZGAB3AGAXZYvFKDAxEgINuqqrNyX9GdD
0ZJkR829oWWRQbWn6ay6Zl7m33AGa9HuU3+SYiHFVavIbJNyOxgSRMLMizzo9jzh
3p2esBtPMrOyrmnZPlnRKycJ+z2IBH3Y0OP7+uQmS6hQbJQcG58M3WsYdz0Gdm/3
U7P6+3wvZfyPAdh1zRBqNqzO4M3G21cn2pHinbs1NTsNnsPKvTZkKvsagp6E4Vou
u59ASPDxuVOgrvcoxnL0R0XcJSnW5vilgbx/QBUjcN9XvAg2KKVGPmnVyS50rWQL
wvbuRsC1LaWolidYJVPHB49elIHKjXc/1MK8zraRPCOdhYg6qh7Tc3z6bXjC0jNo
m5Emya3x+Gp0yvGn6uEXzeKlm1b8R6jzq5RQes9FMAokKyfzQOOpAyX/l4fxi0bg
BTRamM9lpwQUmBv40vzjMATXNj6mlwV20UzLIVTB8tXJhoj6Jg7lbYMT51uPgfnm
uOeCyOE3kEyFj1nLdMBBfVYmZ5sF/ZzrB5ZjmDwWxMvzv+kCZiQESZdo3PLfIL1z
BHHeFDAc1oKwI9e3VK/vec+VF1IH7SK8kOOrIk54QsNj1NExvEJKclAYjVGnf7SU
EfFIlEO22yOWrDrogzrvrssPsRU6Vbm/War7SvvW5LLvRv9rMGSdjDzdHUpqTS29
m2ehEAPUIzRD26Pt6twT+xSUJp9SlfdBZR0Txreo3RvDwGnwbMrlqSEmx05w00OM
j9wRFZlPWCnFNP3mJl0fOvogp+E0oQoUHzdcttaH0TSQOmdZYDGpZQutC4kIJT5L
jnEB3JokaQjT3i5z7bW79NtMeEksrkOFNi9DWA0C/DiPFrlUpfrHRneu80MS4Qn5
3Mht7eN5J1o80ItXa2REOJwdCNwHbslhIypcdTUw2I6DIoWsLb6mZKWyv7VcIh/T
NO35gk3nCGrPgKGCfbLXtSrMxABZaDW3+/MYFTyJUg6doWKigDSoPS7fVV5icm15
v/AQuqisYq/Da8EFKtoawytk7l+FEdAB6ivSBDOGVI2yNCzgIF3XxKstOmp9iE7r
XgvH8UffJDr38UfqU9b7CK3kfF53eRJCKN93CPBZJivooeroBvVkoNz4kigcdYy8
8h+6fYE6GnIRUcBNEGd01EhS5zxZ+QCHuDEPfybnEc3+puuMUPVFiF4MMGHcdbrc
x1J89xz3dQBVi8ezbBvRuvoEs0+3tW4g4UYOI8CjGEWUyeGcv77gxEHxMZG2ozDo
KX7RcoMEtg8cjBiZt9VaeIfPtuC265vHMMwkywxg+5N8fn6ltd8n94ROhM5KXcPQ
qJLsxXTPaeFYiUr+XKAiaxSOhsPmEOon13+W+lr0SjTmKrrgVrFZZ7HWjWXkPY7Z
c6iq7+dRTRIcxQE6vTM+lrtl02Cu+twMicYfPhjuP8bojzrAMJcPzJXEKkaxu9iT
9oLcfjjZA5OKd17RK5rRDic8Qqk6Wzc4OQD9TO1m0KjiZG2Tb5Y3ek+WtNpK6P9K
VXycvmpN6s5n3lnkxyfmJ+SwCD4ZWMm0mb0kz/aMs0aakLcq+18UbWq39X3HJjG8
Gy+viMPIx3Hcj/Ptf/qknOCNaKNg2BMNBJt2b8YV7F7CRwuqy4HbTxiwjs4Y5A2x
K1I2IKX0fI74XQz9gv1Qmzhz7guZTE5Sj/mZPmZ9RhD6R+nF+l6S1xLSav+HVgLH
A1zEsM8mFqwHv9YqkR/E1ngOmokwy+IqHd/bYJNGewhG+og3wSKjCBgNBYlClYC/
Fq2CbJjWuoCENSJ6d9xoDTLFLR6+6Ydciq5xJ1qoEC+yIfPr+Ckzb1dKaZB+JmLE
4clD3TcOi9VI+hsFyICvFcSIDgCGePFBPyJhu9bpSALYiyfCZbxha92uXf0Xmwwt
Us/liZqL4rTFmuuNY0l5+QGFJ5iax26fupBdJA6v38wt+hC2qoI68PAzlz0Nywoi
nAJgx02P8mvcKBq/h6Qw1g9ZuZTEVOHiMO8xqG1n6MDBCjglAvCUbTUCTSufwaiH
mv9zFYrQu81o1Apg4iAtRCWjZis0N6aqCt1hLhlss9HaxKdQ0BwCSLEkJIRD/j2z
qmVtKPEktw4tpJlEBNebTbd8cct0SMt9LvWbQULSoTEebYI/Hph9qhjoIphs4ncy
bvTwnztvT8Ex0DlJ4Ls3X/qvbwCNlzPSYZ7Jx9hwf36pjw1leBKiEJqLYN09GcFv
WV8FTTJVYwR9MTSarADZeq6qWN7UGWyn7yXCMUQIrUKac5RXcvinT99kBhnTtwaq
o5NRC/ISs3yQcrV98afwiHJxny4vaPb86JimLvyIBpt/CyjeQggCpw6sM2GdxvFr
KRNqfbVtIXxVpYoOK+sEq7pqLNy01eZU9+kqWmHOF287CRMyD0K1RUf6RRGNEJUp
A+Cxs/mC+POgW4q8EZ6ScafhCudzqU/kSpRXvHwh184UK99a10b+VPWNXsh2+QnV
TF32Hgwuh8rT0K5kP6WWWFCJ49Kc94TiCjQPDdNeX+69cavR0s0tj0KnNHUwhbgI
QE3wPaVd3TShZR4tCA/x+ii+y1tmf6refUWVw2qR0tKuMcQPtG/h0FiM4mlAuhL1
7Hzy3QIys9w+23biCtvOZNWS0yfd1CYxXSsTftDpFnIs3a7CeqjBhSnGwW7Rdcbq
F7U7Z0UgWw28gLzaGCIXwAaKWI0BfccVrS1dQY7RNtXLvwoqKnqvoC+f3+vAME/h
g/3rrFNxuroWx13KpnZbv+CuMvoDjyEwfxbnrHpR+3+Y9Lfz8Hkm+iT3iRNI6RjH
u+GVBt91VlQEU0Z97xYrOMFYoutTHcdJVY0a3gCsjhzdxJV4urF1BfThu0y3HRZC
8zDWtwZioTcPaMLkoCHE7S0Oxd6DkpFJTR91op8aipVy/rck2CGsQgRncfgyX6QO
4EtsJVoBoje+swQyhVP/yHlDdQOG3X/ed287xLQqFAcOTSHv57LmTrxjiI3LDKOV
XdlrqvFzIXbx00ml/EvIR8ecZhk48V4UYdjn30edy+S0Nv1+dfmW71ZP3IwtytXG
QzrAezVHfX9V+b44PxTawU+LZjuE/R5L5jK1I2JzVjWdIJ9nD1nimKzwNWhUhpLt
QuaEafg5FwsF79kw7p5d5UlvSwcQ96mF7W9BBRcXaYGwtHyAkXaQLl3DASnn8sbf
1IY/vI00+/Nxdzrqm4OjuK6xlrghh3wSjulCBlMq1VPx7gSB6QEt7cKGBaLLfthI
6PNkRyEB6Rz6aesXeClgp+ZhQRllEKdUhVuSesscGnZJa169hMC4/lhvef4vF9b6
aZg69SeQ+KUo3NfqaD2gcAryPbrgxNqgtZrFWpc+QMwwbZA/vnP1b5VzSHAtjUi3
XjXgkLZp9obgcQytAZe3JielPosdl8lcpq7ud/zD1LDCPngyZR9Zp6q+5jn7NgQa
mN0pLxP+MJZi095TJnHl0ceEYZStwp7botRcGznHFe3h9iJ/vLadaqpcsYN6nf1N
Y1i8xE3EeWFfk+gKeIh4dLzTIB7J4GNnTV5UHGa/ktas+YKv1Lm26dP6chyaeS9n
SR+DGLqeeY9PoObIfJwG+eSNx4ePcgiQQDIDWieq28/2n6i1JPTnizNwcM8jvWgm
aNd7k0FnxXtnQrBVOQdJMdL8CWSiZNHUdMNPo/PT6fVycT2jjm40BCS5LF1nFgwU
I95ze+2Ln9gst+/+YtO2H3aJTCAeEomqdX9jvB60++tFuiRx9o4JfC8FARX5+UEy
nMxL95Hk0ulyz9gYACmYW7gj18I8Eo2jlNw1aEy65ac+2IM4KrOj5+AxVwC6T0MF
jK5hHHooSwxKGDuh2F7/qPGZMfqm848E/bmDtqx2wjDlpeO2MSIllPeGbUOfDLmg
sLcD/ojagT0tDC2iZWQQhIU8W77EcwdrA4KA267sV603T5FqduRGBDZaC1Z4MLDi
VkD5pPXXsGnhF7gzjXPiFZIr1Wpt4RNmeNjw3y6nl+VQd8zxped/1RUTLJXppTNy
FoDNikTyjDFwpS47SGWnyugrfxI7tw+kGuxWJd6owfuXxok9pu5/QDHvOhQb4qKV
HuP/j+EVBhTcTVkln+PrkuJYji+sAInCX1IUWa8WzwSKwGtlYoC7zfKc17q0/bkH
f6TihBQUgTOkN74Z5feVN2iAkLeD7eMUzd6eDrTMxTDRQTkaTUMNiwPOaGg2NsMd
R0rTIvaEg1esSTTbr/AwbPC/SXdnEQ2aF/nNPT0a9BtLJEeh0+iL3tBMKtTsZBK0
bCBvcdz/xAnPBXlI6M9umN4PZqRNNm2ycE3+Nbii2pp9qn078tMD97YdwKRoM9tE
AinSKh3pdxrBbgfUt7N2I2WVzk6+AYdO3zi0Aqm3bWFq6dHj3LOdcu9rB4wKhhj1
0WfPNsMNi2SV7+cvN09XtdnmsiJGadc4C3HMlVD1DgrJr8Hut9mRqWk2SGb+8BwA
1IIxxmYi7fdDOCqw2LI05xzYN6fdjB6L4RUrLsnE38V4GC5P63dicD0IPlM9HqW+
HwUOGEGjf6lYGvitfRKCbTRkZpACDP+o3BMfWJejISFLQU2VXC0YFp+ezI+iyT2E
E06z6TPU+06Eo88LFQMkfHcn3B9EM6E/IOeqSqFmNUFBYgDp03VBHrUGpNEz5ByM
GSgOy49jpA8JWz6hF/RU2XKhTd2cX8x4s1zX0noww+RQQslKDk7pK2u8i2yxgE4u
5q7LwFFxI6jCp9dZ5osCwbebTHADwM831l8v++BO8l+yMiTnr2pki6/dtuRb/V+1
Hy0Op3coUH+jB2VmbbTh09xYAA91JJNFeuWC3nNNbAaFB/RKH0RmO1jp3tW105gq
7iD0u446faIZ7rboKH9zityq+SV5xcZTSOyUgMqHxnihwu+mEFwl1WXdRSG+KeFx
8wMB3lMlCdPx2Q7xqO3tKXFPwcBwrRBMRXW3gRMDRKIDRSDHfNWJhxVUSZ7yy9+d
F1np4T392bGpj/2vEmJ8tdhI0PC1DSC2lA6sJRgLFP2QAgABRLe/t88yH5JrflpB
mVostGH/RcCNi7jtYt8Zp2iZG7be95ePeRdoBA5MO+GAerPTItMDeDVqxbWQFrDt
q3WOcTLBqGx4ePMVYrcSWwuYx2etxMZTfxuXsEZxuCBQx0JJdbPDtjV088rV56m0
678yTvYn7DBgVtp9kp4JNvqMlbjo7HvLCpa24mzpJAmp0mygkxVqbTJHkkA1Q7Ky
21Hcx6kSC9KSflqHB2ZbpWdxzTf6nbFKH+JQ7Mgu+JLMYkpKqCtouMLmUZinwpUc
0otrTyGj4rVaWEA0LIRda2uniyMg1AygncIPNaWF36xCnCodwaRnWilNjjkIpp0X
3O0JesYMOhAS34U/ksl911t8wz76IzSS5MDlH5Mawa53xsiRdbIbyOSEjvnvPrp0
niD4tSyQZNq4i/uo1Ewc1AGPke7n63qkqVbI6dq090T3wAy8qgDOCpqNAwKHFrRY
ymzehUZ7MiAEXMfSruIUfJv6eqk14OgjjXIpzcdv3l90CLdPu1sNVZJyvv7VE+VU
5lFI+lQ+eQaYJQayFi8Nesv32h/HUKxOzMOkFJ2HQG79jOh8HONeit+LC2Q/nm57
AhCdsD76zKX9b8LfXgGFnFGwp4PeozLt4/3cMFHwLP4xRdLm+7UPz5YepPLCY3Vj
1IWua1OP+Rp1tFbZoCsNzhpZTI0kys9aHSSprn4tj1s2Alw70hwiG/fc2IanN965
3sGj1Ph9Sc+QUi23QP1sdengfftO1QVkNLUwlicWr8kCNqJNoxUdI3q18vlu4M+I
XBwGdRt0lLKzt2ZP+T8XoeI+PUMugzELexABUFhxF1eDKWiCegnrCjMESXyUMU9n
WHPLfbE9joGPmSBr0UCrSYBWkKq6MbelXkdKf5xTB1h076O2ultE7RXl70xHdOa2
czzjPyx8GRvmnJClPimKB18pj4RVk9s2CHrhosPew5M3+nj+q+gQsMlO8/auX8pD
8vx3s3Mps6sOxNNjTcwetyKJK5geo/XhlYE5OIZ9inzFXZw3AVpz7EqWmec61BXO
wf4UZNf6b9Ly2SUUjzlNVeS+zBUeong48oRgnhL40Nwuw9J+Cx0sF6XyPhBDkGFB
+oVVmxlnBApkXZkyh3/jmO3DvHTYrTkgjB2O3URxA4aLPVIpHUSXui2gPk3mRaew
5kvv+b1mzoGoL4wKzi+sE0VjRgbc/krJXfLnWCF4n7Rm6KKYGXRnTO/BtJ43dXng
S71VBde1dlRzSYScZu6iW/xYRigDktuFO0b9yDtpcnuvIKQyEE90rzdiGZSKe3h5
+zGyT1kfb/uIckq8h0G/hHz9TAgGuzDIv2GBwNHNwolSPMR9VnDvUc5DVjWWFulx
YHJebiCNZ+gy0X/WvCyNkVHZNrKO94/bkFdRtF5V/vVQgPe5eprxAHICEeFP6PeK
gdreLL+fbK6uBOxNrD9OQ1t0LOLRoyJUOEH8voj4U+SHF0182VqY38R47za4A7cE
7vvaBpErFWzziMLax21AC5D4wNLrQDm7QNb3WH3Cv4CyZOogyMN/cNVVZkixwwKP
j69Am718W0VBSgmm6FjAD/5bqh1NUiolf3QxXL3hYndkT9W2v0cVpCPExOabnp4g
mr44KSSFxUZ1/gjuTOsKl7GBUrgsbQEnx8Ld2nPygqbDlh/Rxj/BYsRGRqrWgUiY
1rn2cHH6BaABBpynl/pVT8B4Qbsho9wkLBqjmSaH0XUgg/X0XsvaLxhCNpjOXZOA
NlLLcePq0546p81r6x4bg9mqXfApm8/iGcDB3j8hZWqsosgyRZP1WFpSxsTJ44IK
JsTnOi/RXnDN93g1bS4YiWuyvZljZILoASqrzgPHtgK2Qn7nmooe72KN432Vkx5v
mSnoSov4KJSRoSHgzCmf7A9q3Tk3ToUCtHAJFqA+T61/5jNXruRp6G8Cj9v/yAp2
Jpz6oA79B9SNThQAToQ8Qcc6z4YUkwdE+mSCcqcLjZBM8Zv6e5AnkgICVA5nCSQh
esuMilpuRfiQupRXYTBnaZF/7AGon347/LYJEqfcrpFxKS6Jx79Cn5EPwTI0ScJm
dlhGxqVj68rKpMG2YrordTHBUh1zwP0o7ZLHBxC2AJfL2tKGgdTI7XSkQZH60Ubs
BYHxxx84aGukfxOORAUQq5O9A05tUoPBw9LOG15u5O/cJlPuDbQLix0viW+0gNgT
vnzVsMHat4xViesrv3/MAkDOf3MCDpkP/ofF4sQyV5D8zviHKVacuXuYwfCDdo3T
o5hxXRrlb1ThHKLF64egMpaNukdt3e/xEtaPDfh8kERLv+0+Ni9SmGHYW3sJIqDk
MpFgirGXPTjz9vymM7BFWhL1lVZ+DNyTszPjjmkFfxy4ruIBr0NN+BB1xskNbI03
oqgzGtGcKI6wasFkdN6RlaIgwSInkcKhM3MMefCeOm7+X9lupz3WQDJX2A5cVrOz
Sz+SeFkBxWFcn3SyprmpgfKWv1JuVKLSVGSncp7DCebKEkqISqWzd5HbTRqqvXUC
/ak+QxNUIFOfx1jMA3tO3GLr1+ImhTUm5x3MrJsLd5ILhTGspHFdTmPOeNqpRiEb
fVZ+zWMd2zzAsZPjzPXhLOPat/pBIQurjjWgE1giT8/WJpqmiihFcK8y1wyeM3SB
TTDO1axneus4uC0GxP4ZjArBhusTpXUG7j/9BoDM+jQu6Tuubur/wBCtkMD/1WYZ
3AHkxmMZSHQUNKzXpklWLz3E85cXWZKmLsyBnA1sV9k09yjULvFnrXpt7oWvTRXP
8NTQwHUHyMhd3gyooYTxNxf5QRVyMCMShLfTPpCdDszbQEQmohN/twkjF9Se/OL2
wLvAmxrRV+UQjyjq2sYSRqXEE+Dux3KsD9NGYIhT4ENG6r2AfbV84C2BujH3aDfB
pGB3vD2uYshGmFgSg50Kt1Gb3h/WtUi5iVEaW2/uadYTFRaJot8TLVXjeRERihU4
6f0gnuOFis/Icch7us4YfVaxGL39TpmXtgFPJVMno0sCD0gKuya0NzMCmgXMtYvm
HnUPdk+jTZJs4HW2ES/BW7FK1o7JHYwqWZUW7HNXKVTOlgoi96e8r2PCga/4Dx9l
x9nM3IgkzUQx5vwbLkhdJTcBR/29eBsluLsWmW/deMAYGJ13GfRzoKNWUW3jZ77D
ZSh88y9UAkc7jRp6qCSBZ35N8a2Uf3ewLjosaHg8Deqx2Wlp5XFTaaJlONzjizBs
UE2aeJdFMAagR+Mygn+L/wKCuZ3kKkSB89XHLiTKMzHIdQtI2bX77GaBilY81EgY
w8tLPgIzw1XolAu2PWJGNGRY+OOmraneCoRLw+DFi3TeUXxz/t0oZ7eDVHlSbMcj
B0e76X2rapa7H1ctt5JkvsgJY0yCaT7PJuE7XW4dzZiTwkYI33KCEO8t13+puAwr
QN1usYic0YEbwkw+1JgGqJwnv+fD5kSpsHDMK/5142yz/esPQbAsxP3WuFU+OEgR
L5+l1X9ICPylJzp0R1jfWwH37W2+f/9tgGyBejTmTkmSHHLYaeszI8uycF1zuqXB
fayLginpC9IrtcH+aS8mrZsDrT+tlS/27wo+K2AVhfLxAFlbyP9YXqCrq7tB1dvL
kkr8KQK5YRsthpD2qaZxMRXOVlg7962gKcZSFd4C+wXENIQaorsKyyWlqTKFEQb/
pwpzvTLUQGpqCDrpO8ZGCAAm3+uraeGU/Sd49IagG3djAOIY69Whx7+egpslFBuZ
6VntxfN/GoKlgD4o2NEuu2oDF4w3F08K0zVrWonZnGGE6pxQ/7LsbQT+GU0yF23i
4VTiuaqRcLl9RXDr49tSyC33Kq1OlfVWvxtA82avsr1GxWn5A8oJl7gF5irz73sM
OdZClVjnZlJ/Enys7klz2xDfBM329bpCF4FpI8MveptjV4moC3An8QotlD5cJpQC
0v3vt1A32cSzo7eVUYMx/rkqq9zZpr6HMvOy+ieNfE+5xTOEOtrVHM/XneattsTy
97yBCguQ0TxEyeTBnhyjzywmRStnjNIc1ShBqZVeCW5/hvHtcFdANH+CmzttRy82
/Zk0JdSPP/fgOoJ7tmlIqcf+XBxqTmQxz089OlqCg1NX9glY86Px3xJ3D+VrE5lU
eqqvHGiJE/T58n2BZBXeEGLsIfZ04RWuotbDrBdrGcYBj4/nKRPux0b+S1TI0DNO
ayg6rLODbTqbX8HwFBN3Z18EQMcUjTbe2pDBDB8Loiy3hFSH4EnKfRhnjxSXOpQ5
4fLW3lXIhHT9kYlgtB+Naka23aPLr6QcWMkoJbp3+aiceTxxGkMkhoQCif9P7DNz
HZA85ZyK7m15CuEb1fNOeiq/gccLMx9noQW8nv1TkaMCyeAaoqGsVfYJWRZwUrle
GEV1JyI/7vJPQM05Jf/cQkgQ1pL1cJaQASF89QUEc6eRJ1a/VhFTmzjDrIsIZc59
s38mLZn42NLb5yltPE2ywKHY+Ej/rxR4X7+rwXWKRVGiloR1jeKf5OJuM4Ct+dQ1
/OHjV/3WS3EfTCkoCvT6jSEMzVgVBbAQxOJemWhNIFEAza7hf7/Sf06GKl+doZ0/
B0cnAQvSjn9b8NF/qpkUu0xmZ9y1lP8tHtHouIIcQeVOe946jsEp7+pLp0ygTL4D
G39+7xTZXdkq00EajHEh0YOnmn97z4mI29EkBEBFffxu7tsen+HbBsbMqRcnNqSB
2r9s/B5KFMmX8J30PK/WwHRG8q2FHnZLb9DD5RjtuypvxuCDhCLoiD2ngMxNRLaE
4poeXy+5By5rjTlnTbmxchsdv+xASUrogC/TDiiW1H/6rFqqCe7TFG81MUmPncVH
Uf6c9mxqCmkof4/NcRZAu/e2Cx9gJkxcbl1zQYpu4JdI5DLRjPmf7OZC7oeqzzXa
ofZyGuRBdK6VXOPZ9zcBN9FSBuDtfExuQpywoivgfkxx0ypHgFwlh3mz8IhgqCDq
Vlbcnohm0hGR7Tk/r1NWJBODZ1JRzQ179SRjHDA04vsAQ+2ErOegGaPZQIpY6kaQ
cVGd7DlJ/R7ic1y8hZ5KCi3yKJn4Hm4wObMmIinrYR6RLHsW3691umYz88UQ1Pmb
BrupS3NafXdKMjgS3xYxfLq7QsamzTzauYciWpZjkObySVqbc7rXtnyOG+QwhTLf
kA8psH7KdIrSbxZWGeELrniGOr4F2Q5EbkUe1Y1MBNR3SWTRjfQKpufelWyDE4t9
gjueTtz8Mr7XYBzI9CcCHljmi7C911CpIInr9xFgJowCuJ6R+xQMWASTOKm6i/PA
PxiPm3lmR9Rbm2I7VX6pCz9Xnov6x2+VnLmD9JU6ipOKCG60imZdlbmfC0rC7gNh
gBB7TfhAjynGgIHdlEOhJekseSovr0+vs7VskhjEsS7vpL2UTXgLZcAXvAzkIytB
jOw8nj0MG3F8a+GDjJ0XZO13XpGmIg2YmH9tWF9ius2VzQ2uDXqPVYuK+kz8bC/4
O8XhPuAPZd8fWBX0njssteclzqbmz1civlS+Qcd4nQUQbiN2Mfpef3c3CbMiFoOb
4JtUo44cH95DyCusg1pTAUIuuT7+oF6tfZsjVYvo7NAehpOaqT/NBUFBREH93YAr
LcBTQxGTu4gEvW3VYJ51qZlg/B1L0K/IJV8FTnIyuVJXaUTBi6GY3AreqDZBOotN
X5XN/t+22bzqROv1sKOXBUj02HmYtp2KU/t1OSFd9YQ2aAko7J7pLdM/U4eqVI3P
QG40LLFfIc66ZVDcNmKbTxYK5ji/yrtu67DQocBDxB0Uhp+7M45UTxEbEunmTl7M
+3CFfRjYF0BJS4kyPMj0Vt5QhxanmpfXY/Q33A4btJqvSAcGPEPB++iVd2n4QKTJ
dyDLHoNG1FlGd2LutzBgPPnBqZpoyB0NyyxAky/HFrI47IavSuZfaOF4pwyyncRe
risSPEeGRB6mUeLhygeI/Q7l4VvoJKbiuzuvTVDulzLyes5jML9ArrbXI4TZqNKW
mrajPr82TUg/7vst9Sek0tF6PtfOxKvjerprSH0whL2NB65KxH5/5HhjX9qNiF1m
WlQ0YW5omIoRaWHvAtWmH0fuHm7lxUVhylczEaXt/Gd2PzPMhdw9oQYi6PnrNhFG
P/khNS9BWS7XOuwNWGzU4qhzisucZnVZxQ6N4tJyXpxMytmNqJYH+NWesrX0D0QB
kFG2BCOpIr5XP5y0ISGvF1ai+nrbyLvkWFw73fNA7xq0RD+1nudcxS3Xbba14V7U
kbx7an2VHBFQXo5dzpJvQzWOBmj0POf7O1XZ3yiys71GeDSqYEuXrjlTJx7Ih0Im
Y4fB46Nz4PX5sBA2Fwg3u73VSsqIlq08eY+4kylyLEy1fBIekLN1746wSEI0kjM5
Fghe7ASK1VFMvrfXvpToa73dovbj+yD+DWVfHi764rTXt97EB0142DEeJHnkRyBu
U8tVFGYuRppjNHtzUVMrjrsRmIapcR/upyRpR8GnyDKDiS7rq++VXFjX1LtdLIE2
GokiIoOAH5Y6pmGf2bzAAGmafxr5JUQbtUxrAzehyeMf5K7hfyZMHnKKXgFbsNvY
uZJaS8rvkpw/owvY4NokpZ3K6wXhK6CqwGLDYzGmBWN3Q24tHtz1IsfhlYv4fSI2
FyVk6Ap9ObyK7/YrX0jblDMRKcE5le8v8gE16zSar1YiiMN2XR/2QynXmkXWLd0g
f5X2zZG6yVBuPzWYWhZ6g6dKjanS00zcDLhTB4wMFE/pfMSmBB8Pq87tqH02xX7I
RMEzPnSpH20VYLegJ3ddxaU1R0QM6H9nEpt0op48N6UyVzTqzouGPFp6InysnlXU
O4AneKG9GhbSswCPFd2TDVwGZphWSHsFboHBlhllxI0DSsTteYKvJgJ2ZAHE/owW
gwqcrZXKozcitpcmKCbjSR86Vpx016pURFS2aHf1QWy21dcs5T4HdOUaYrRnO1+/
gbrtqzcqo3YB8YCY+ijs6sCpbFw4RjqHwH+/L5gtllSyg3fp+XTfLM9ZcNLU3TgW
n9GgfcmBtFVo2pA6ao+KjYeTJWJ7j3hzxF1La3Ao9x2VgVb/8pfX0c7h+D7L7me4
JTcVQS+UBOZBPu2MZPL6kgjHGAXzA09d/y17+GMfKfx3Ki/y2iCG4mYrYbnC2jM8
Ov55nveUPjQeqLNsmC5XiBwkSfKLV9JaV4bZkTz7rKOVZiW8z5FWnayrtJLy0dgH
Hu6ERRJIYKOmV7naj/kcYSLybB08SB+f2yOG6QrFjDK6xoMddiK94XjPzYRfRHDn
Ze+A+sztsaciO3ZHeJvgGzYPjlA2VVdp0aZg3gnFCo/ln3VvoDrnLRoZTNOlZI86
Q8EzaRrudoHkURsx0/aKp9WE6dTHUI/BG6pRE7aENLUrg29OslqtZSuiQLIXft+L
gEFDhl55Qaf0l6cMbataucMZJ9rH25s/Pwc6nWplg+y0zuRhYB7VK1Tiphgrkx0O
C0MNsDPfMrEZXODIyuf1sJh9xSxDwBJtE9iKcDXo1ekuOGB5a1EAfIK3g8ZMsPnx
TWbTDXf07a8jlJIkGmBT0pBtVzEQzHnOJgLwYLuAIaMMvHjrSFdC5sx5qpWHsEE/
UKH8Pol1S7Obwn/lbWs+0kzNepS7X5MkX9fROzQ0LJ6bfgHEWtcxpVhYSmmb2Go8
YyrGK8UFa+a6ZI1UmE6wK2EhOMYGmFXGGY8pRgt2S8TMegcTNqSRadVlYzxTpzSp
fLdb2gVlP7c1OWqxuJN7HX62yKNPX3f6l8ysF0ILDODXrWCNUao7nAsnsrFlGKBv
YYPV9dWdqpHHHMZpnxSVk3NKk1HUhadJ0buoXZs2jU71fy6l8+S4jbfVv1Ghl8RT
i9yASqsb9ScIbz4d63922qLJRrTOQUoNHjca8VWirfZK6cLSvJ6660GFboXmUHnA
uSjpzmQgz8qPoXhHQVO64UTM6bSoUY3v/0x1IZcy/VsGjid8+EaabvZo/DmQYuwU
JiPbCUO7OCRQJ3hvIstbpYJpnLbVi7Hs2Xl1z1CN7Mxs5mrT/G4Kszr1sqXwJGoW
nikl4tPhlgAZSDfpy5TspimEBS/WWj9WMKDioZ2PndR6ZBdid1eLKzJ9i3KPrFNw
De56vdXymGKAgLa41jymajV+3YfyFMQIfcAv9hgScED3RJm4vRSYrN08wmMcC5au
2krQ8jyyhX3WNYyKWc/LYKNqm6Q/EhmWTm2urAlPJFV2EWMKwvBHvfkh7VBdE6Ki
lAeSDfAh3zK8jkCus18bz4bbjyoE4D05X7paauJadsckS3X4m65CwZhl4MMUsLT7
KS40gIF+jN2beg1R70qW42F3/IM3toHSuCo8sRdeWe15dOPbLMT3p2w8RrcF00Ad
/cHIgImFl74CzPCHA5juBwgoRVjCNeKA/elDhNHG36WveiwSZUeKs5EcVRsCuhuk
eKpRc2xWH0tqMBwC0Z5ajxCnAqRf3Y+z+4kCgpsvvju7S/RYxaVYuOeckwLqfLIz
ldza8PlIsgyv+ORuZPlTJas6inB3jjATwW07HFnV9T7tf81txSYJX+GHj0NqVvS9
gzc1mXvCWcCiJqwe159gz5K2TQy2xvWPZBob8aBJBjjIhaN5zNFXuQscQAJJjoo1
IoNae96O5+Qg7fzuHXdPXiZnTGR1YsSBpsNax1CtNR82gZ/K+QC59D5HpuvtZqCM
0jXPMOzSdqi8hXZUr7yyh78kkbXObSbJQVDVgfGY6cHphr9bSySKXgSsXzIkFUKH
jGRhMgY+OH4n3JisYLxwR/EJqX3Mc/FGQPgH3hg5wUIn5qtet35Z2LOvQFkTedJS
b+RU4slPd68weLmq9zL0gNwHGTLKyYoSkGh6aMrsXhEPTS5mRVWVKghqV4KhYOPk
MCYvqbahHboRfGtQCGXr81pR/r/VOb2o3e0Gc8z13OEc5SzgPjPLfSTBVzfDPtex
RPSld00hf5UZgNkqAh0F27xKZ9gSUYNsnYbV8wN93Feb9PkHR2Ri+7vxcRFDc2uL
6oXpCqvv29jn79+POYWpp+HDL2+mfjehg4K/0R1YQSmAvqKTo2UCYAjf8/Gx0LM4
aBEPtoIv5AG6+AfyIEazSgEekd1VJI+witEFuguMrHhEQIyU+/K/pyl3Ui/JvXUx
ttPMlggg3Kj7CDV5lV9KWcFSYJ9r/7sFPWasbx2W6Y+//EMrAXIVEdK/2lTcdz6E
Ko0P3XZJ0JjvwMj9UdSUVIFOhHOKhz5ITzOLh42cipMqWxiuQyGS81U8dXvqk/se
hCaXPyua/p9ol4qAxT3V7WUH6wcafuyJ3d9y5pLHz2accXr8ZmMGUyOu/SMythcv
tXPy6hlgKMeFKQ+f+Gat5kLebeYcuUdNbWvFMLiG0O3muIWLHEJUJkg9BpmqS+kF
f6JD4l93lwplN3lnPa6naa3ZfANQjDsUKnDTSQ1+tiZ+r62aK9FUbLANaSotZH2M
xmuVDK8up9uEemY+s19B9G1IHTyqtyBA6akBvP+NCKuEi5YZ6DVsoM2AQGvdYxW1
MVbIxSizArfxghuazZUzA0I/etef9Y9Q8MYlzkQLsf0dzJxvupgqAsE3FPch7lxM
aPy1K9A9RjAVQPF3pCc2+nyxiHsZEhtb7Mw2sIJzGXNRDbCaLZipbG80mCzpNwO5
MuOZCwNNedu1M9XXsQaV0Kef7E2+xhHRKQlOfEeDV57sx+4YAZMrTwBX+wc/d/NR
m+SV2sqnlrsJ4qkuCw2CwY6RTfhdgPCtTPxiC62GKTMDHwInTk2o+MTiaSAyIzSs
Ri1z/YsM+HWGco5/owyU+MZq+EGP1I9OSd9JX7iamXyaC/BSSUg2QvyCrSxbv0ve
1gZx+wJWGhX9sdGjggc19BaNIQHtoCDa9RRv0Kv1ZL08SHRQw3bJ8gb9cfxukdfV
PXxFyJ/YWu13wMPorPc2JtHl4ERxPxMGynN2uNZS/lj518y8gA+Vvs1cEgu51yyY
oH0L5rqY9ByPnguio4j5zfkZw2FgYlEvDgjGNjb30bNy9wFzjPNk4H4KpzmPVUie
nSz+aYfIIthppWeQwyhXSYp861Sn2omEB8WzE37VdLrZYBD0Fmq3/5TT6k/cC0CT
GHeGlQOi6/s3rycmF+vwtgx4rhgY8IYHvMKNZO3Fju2uF4TgEshwHMPMY2nsyf49
nV+4e6yvLJj7K4PbZ1+N0d7kGpf8L6WSNKMc8NNQ1lnct25FHF2/P7mGSaYxx6ia
BjHDrOZe2V1P5u6a3/G13BUCXQVOkkcDT6HAM9GoayT3XGlEpogYOdLnPpEr8tr1
ATpBxEaSMcE8yCmyMfAUiVuyOKXtgUxExvr99Bou607488ad4X3tPlGEM0uvxQeM
LZ7a28z4Vyrjs0qMcTU8qyR0PBT/7pTK8clUHPM72dmGP321S5VZKgZmJ09xSUKJ
swaCbjWBQpcg37DdB4mtJ2bk27MlYdZDkg7Y0sj69G77lkgS02KqzbULLqs2WdqT
mdap4cVf3ubonJyE+QoBqEfDWBuxrVdYilqi4GQ9ajhiCcP30tW+fJgFgihW02GK
tITBTaV9V90n8zVnG9weNkRjyGPkbLA35wsJUAbaRiPXd3mCKhCj1JB9XBge7Oq2
58QVubW+9jN6dSEDp6xE8LugEQJxBD00RML+9p4XnafXeLPqz7cSt6AFOF4ygaiH
1eg13DKqER2iVOvKZxGLzrRUyDqA5meVPG/pejQylqroSs0cgfnAfRKzRz0xoxs8
o3SZnPbmD/EthVRTXrKYijmxBiVV/fdDR9rf0Y8UwquPmFEkwZkeu1e3TKZfVhHX
8U5s/Z3wgySXmS9GtX83jnNPw4dYGSvOV1WLdsk/YisyjwoQrbJZVJn+2hg+2M0u
ElHOZahB+mf+muXJTNEy2byqJJwDm6lMSE4tcunn7jwZL2yEJlZ82EsCUf78HMqS
R147Ss4qZ5nYw4K37z0bw75NZPnkqX/MtDix+A8oi7yaFiz92qJEGVhBToA1QDnO
5g2B4ja3jNVPzFv2V33jyAYH7AGd2pGex6wzVBRdXpjq1JBFBs4odKdjICXD35Ma
ITaj7brDpa9ZRLlmAOmFFas+/GygyjqrErugnzotTF9KXR/UT4ywySHnbA/CUKcg
Isw8GpxrsPz9yha0jc6S2LltlyAglaj2ZoECjxnkoNA1i+tbed3cNelfMUoRbpFI
l6/KsNN1yZMKNAHunjltnAig/coAP648kA9v91lW6X6D/J7FFBgT4APDgwHA+hXr
gX3MzaeZuhyanOX+N3WtZFp9GB/egGR+JLqBbiMA901HgQsl0llg59GWdfwnA8j7
ib7wAbM8zN4ATsIn6PsAJP0/QL6uLr13YX8WzFN1k0MyFcOJBjXCQxAK6WuO/ruL
jaz3AcHN2D7Q6hJC8nEki4uUldqdFv1euNRaVINDIfKGQ0hgpXZex9CG95b3UMvF
krr/SIfvsqAOZEqLhs6DS9DcbsF4pnhEBQIgE+4NKc+JIXO7dhq3uR/900lwLE5j
S8YAY++VAB67rHcGvYJGSdgLhjy1F1tMJaaJ3OlsD0Ru7M0rtANqksNagS28Iot3
oa6zIYFAzzcXwXCOofODABbHUw86eACaV0JVFvp2NJM+jD0PkClgo45djiTRnVGB
lQTsE2XzyUS73uZ2U7BcYVuVAe0KbwMomYxqa9cbWJR8Jrn/WC5VMKYLg60xYkbn
ZhxxWYgbIR0dILIcdLeHrDvfQE5RuA9Hg3cPZHTHdBI2AkTnwQFYKfFFifpSyugF
cBzI6E13fKoBB8rpJNm02RuRK05BLs8OJRrMlrxa7bh5ahvcZyej/nIk1quDtChK
Yu3Fz855lPp7jUbCWzjkAtZ/rPfOwuA7w9178K+uGfHihVmwC+aTnwMU43aYZS7Z
btB9SowbVrexRIZcDNE+TsxdnJ6WHwOJwTfdECjX/FkJYqtqg4tY72TtCaQcvTGi
0Qw6Gnu32m7Jrgc0PClGsqF1vhQuQ+P82RifKkitqp34lgcDegeB9ERLReDMcXO2
xi6m0imlHRvQ077Gzzrqyu/4UDbNxiCY9Q4i5vUdoi+BKMDu3+1X4MM7TjIc2XVP
DVIucB+cbt/y57QcW28r5S3Wzs8uWb8btqAeephGo8VgsiAiqMOAsKz+GEBCjD3Z
ou8jJF1PZMIUzTSl1si4A+jeBwo1iPPOx8gcO+YSD8fKTidPtvtMHqbE1D2o4bhN
U3CuPWeRetS8g2ODtR11wa56nMdlJ339KDpP6dQkelu/3FlAGyaYyIJw1awd/Rcr
iNA6Hr/gdfGI4mqzutbXP8UYLvoMUpfybJ8FsYvpFLGbl9nDQVzML5rF2251xvcN
6BU9moJy+MLZcgaLawjPwaxbug4zyJF1LNhQGBh7ZWGtigNju8UWeXj1PJyuh5Nj
WJVt6eggr2V3ye3XOGwxWcOxwtWxAe6Prg+MoVV8ladu0J541DDaK84EFTCaoy1F
r2MecByNauWjYvWU4HehIBzUX+yZTo/mdj7rDQG9NFTtC1nLNPUkx4joyLb3p6W8
+iLbxsB75nm/WGwcjZrsblv5+rwG8OdcF8Yqrwm0uSZjZjrm2H4VSMOded7bnV1C
R2BewZq6N++OZnHzgPreU51SBhdYimUiU9+pDbWnrlA3lVc+JezmtA7BZM3EpEaa
O0cb4cgSflfX/eYV7F7FPGhcCsdRvcA3xY0TjLRokEkTh5SwIJFMKyohshSqMDHM
f2y9ZTaUe+ET35kR+9Qh/KaSZMcvWPXFLmHdaPbUduBDN+Ur9KW79nPB+A+kOxoe
0HiI+9eWTK5df5RQ/bB/6FxBz/a/Xkfo3ZYbRn53EP/idzFkh2SIuwFPNuJzmcjq
48rGB67xoC/T0aFhAhf2pxFKvHxUxZVGHOKcNisTvmJ+QksW2ZQn6QvXsqpZlt06
/v6UCbYddOlgff17TkakDN8FyljpqqejP0Zq20R730OuwbfMKfOEODA4Wrt2lFB6
lupphzV0fgoWKkn4McmB4CTzphR+0Bty5rTDHlHO4U5yKlAu9NPn7OJBRXqln0JE
hnzNNKLUWfiC1G0G9wUXuGKuSYVFbmIReBYpG+v0KW/DQAry4iSKOa2/+g6RpYAX
Ja/vLnHZ9t56hGaFtI/Zyizx+ZG8fxJvVc45jLKq8KjIQ/fUksCLCRQlG9QZh0NI
uhPXHoRNlGyseSxyad3So5RW5EJ6SSN58wRa8ii8HOvO07iX2lU78DK2hXlxmkSW
ZUf+toIuOgZz7/vW7MZIqT6sY5YdTFq7WuPLneIpI3bNv/g0pNgUUmw+muMhS4LR
c6huxOFVJGhsjKxq9Zom59x1C0/Wo3ifm9hAnK0GVz6NIr2aK83gRAdl2oOdOyN2
suSEIlmJwtjBHWHVNJmtMX0PDCoy4UYqDU6shpJIk+GFAk+TCHcZ4gHsqiH/Y9jw
AC0N0JZq3WDcU45gmfULdLKM2S9l5/FzWO0i39Ihx8P0SidNz2n3s9grhVY2fwMg
JVaaOjTfjgEw+79HzJws2oCu1PlV4SwTHFis9glaZmF2Cxx0G/h3qBkYFRsHAShh
yUfC3xc8qypprf19S5y8YZOx2YtARoXPowi/h/jDHMDVa/qdMrOCPu1h9ozP5N/U
Z+JTVqWHkTEK7RAEcw4eZdIh5ozZn1B0KBccO4Y87v+v1/g+4UIGdMOHIpUGWc1V
ov8KElvm+hje2wfrE85xknZedb1ukkYWMDdykrPRIvp3510gGIx1wRHf+y2BN6mN
6ovLYWuvJBML11bMAlQroLYlbSzEBIoTcj0C6qV3/FSt/vSN0t7vtGFpABqA7UIv
PCvRCGx63VxN8AEJO3adQuXN4ktXj1xGYdWfdCnsrvYtwC3MAHEIkmKbZWd6CAtZ
j2Uw0L5nB6HJOXE6GjqurnVb7LIk9y+Ap8Hw7n1PhhURGSic/Fw/Fr/pC1LbLoqM
4SzjVdSG+cT7FJCaD/rnYpftJQWBA9auDQKiT3sfuCEAQHZcDubvPcwl8E3WEHDk
hekMlSRFR6uBSv/sT3LZslIAxzAljCHT5x9Ns3CFecBtvFKdofxoiwQ4enNCp6gY
3dY17vI2OQd6/cc4r6f1Mu2/jtRBgfRa2JGBkRq9sO4qExxeAXFNMWaNFRgqWWhO
00xBYweJrWRuQnrl3FJL9IO/tg1yccXeOJrvZWif8WElakQOHghkN+bs3Dl9U30Q
2FvnSNBh3Wv3MmJWyG6iPXB1DUCIE+nVTzFvKmYQZX+hXIiIucNq1G+1K7v1qxvg
Kq7152aNm27dPl9FEzbuzC5Giku9LL6YPDzkzQANTNgHyvrJl0WO1ZWO3xnXRa+M
eQL3uwuI0HyVQK7vMxRa6zZ0saxx5Mj+mqCyaXNnSRmuujuOWRZtCGg+LnzQrKJI
EKCTT6lygh1LBMQDYOr4B5eUkdiBfJa4RrLmqdeWTqDHPGWv5ygdkGNDoi2IEC/7
ttgRwXmlFSUcFgal+5DjwAB1PAw9HmtLivp5ZkJzbEyS2zXQiBTRkP4JAXk78pbb
iZfr1LDPf0o3BY54zrOXjei1ozJj5w2Ab/iM3UiKmd/37YYTsjnrgPTUwnAVo9S5
E/E2+xQT4eWlkGicUd3VLaclxpGsOvxAoyVzy0M7jJQQV8YxavQSR+RZDTSv97Wk
egQy0f+xUaIjm2SBep52IzvZKuDtOb3pcdNJgWCPbAn7MjXQsZafaR4gUYJ85opY
s8HKcz9HEJeVwUMdXgGx4v0Qo7V7MyKXkFkd2eRLJcTbvTafEMkNduBSTTG3kxF9
p8nwO8OZZGncTO6xQuT1YS3LEC9dnMQfgfhk8sad4EdAZ06aRMcs47EurlMN0Yrc
qUKnRm/HS7SQjZcXHIrAFGyjSelCno1X3S++vNDQej7nyVGCHAiKz2fC7EVBr1H5
agrgpOcHfhOt+MJx2i8EDTvmyj3BIEGa3PA0TvAE10e1dORrR7ERSW9rdz3NA9eS
Gnm3rB/V6VaslUgN1cPXw5T/dPxVRMx+mXEJT9m7uLu0t9+ouMdz57OKXj/++X1Y
tewv95uxi371i96qFaRexdWgQRNChLUiJGzW+xFsNZQ/0u0rXlC/3KZXgvTgVlu4
9WtIoxcTWvtLsLrtZYT1VqXChyU9FOtV+202Ae65+DpQcGaGJlAd24Ek9MQkb1Hr
/YlbVdnGThr6K5WAXkjUMyRjfeIhK3PsJheWjxIiIJGE+XW1i/9d1PJuO0nyCCko
pyC2n9UX4NEDb+C412VsVT1q3qmnwBPlRx/YA3MOuNTZrPmmO7BlWeaV+JHkOWDy
EHdlP4DyE6GDyVn1UyRuRtN7Rd5XkuNeBuA4q5BRuRq6fiCByW/YwlcGcPdYON4y
pp67KrmsfERlgJxB+Sh35mQITiopXWFg1FxNeOTCq7TXavmB67TAS22WcWkzc3vb
LZ7gFlQoh3Jl505BaT/Skh8xjJNUGnXSYxsfUA1yl4ObKcQi7naWWXe3d/iryHSP
mjSrausWc8+W4EXsJfdydeS8MIWhdm7zWeziWS5106lgm2Q2ANVjYnviXSy+6UZz
pee31AXVUm4C/NapHGhT/d3S8Od+KQ3SbxwKQxj7czRwXAOHnG/5K2Tr80FHKzdh
FM5f3cWiDPJLIIMoimCSJfSsspoujEfJ9zgNX22cNbUIERd4DTrTaZhoyTnG6p4H
wNl9Y2TsfvzjaP5Q7Qohb1Yxnsq+lURuKB/nek/qYNxYvHrBzQ0MrClOQgt/5z0+
gJ0YKmGLIkiVmAA+7e4ybL1yDbEbpViTxxg33cLWHO94rZT6gBW5i7zhWfX3G4lB
f2EdNFJft+fGenHtVy7Ozkz+1RJlk5AwSK8SNxKl9UX35Y8CiPoypi+rx0o+l76y
eSy34Gpw/sUVfsE+zvY53G3Z0rZlGKMasgd8Tl+5Ofjtq0YDPI3LZj22p1LxgaUy
u8B5+eliUoj7Bdk+8VvM35RYMiHKm3cKpvfJMaYNsM/TaqlxGXNUXHv5ho076uED
m9nRmyJZifZ1O7YyD6XtsN+KZNFTsDzlt47PyARXfNRTRHzoAMOgjLJ6wZ3UZJOD
79w8K1R+zaqcV8hSPqIkgz+DGAmANTHmeYSU3Tu4pieBtMQbcyOiRCRDEr173s4R
23wIQkSG5svqB+wMknRZ9CK7wIB5jkSJvqE1/1EtIS7kN+7r/k5ddIB5+pmgJET9
UCnRCK8zm3E1gN31An3u0WA5aKAf6ZHx6+YdXfP+w98sgTHJERk0Yy3TCFWraDw1
CI1V/X3JwoKsaOgfKgY+1gBTSPHH2+nasdDN9TEIrPa869OBW0ZHOSKD94MWTZ+s
BoONXiSAnKAIe94O0MuxtPjZYlyVir9FS8Xc+qnrPkIVy5HlO0oZepPAFQSny4Ml
rn+BFuhPwFQ4suGL0LiFpIosMkMU8r8kPPnEwLatGJ8oNp2nNUN3MgZDczubGg/q
Tkfvzoi8Urf157p3ONGAWM/4E/f0D6ytJpZcFHhQ9d8jyQ7gGnFLJrY6+k56kOkn
Kvj70aEJQ1kprBum3A0PVNmnIsgQVhHT4HqVQfFOzV5xbmCmFQ/uKtPATHZnUc7p
3zVTV1ZkvYpxCNUN7dv1i4v8pBrI/rIYhlApCF3dAk5bm6Y2IvzzXnRlidrehBj7
D7brjuvHaM9fwbpGgQpTEwZL3BJMfetbUicmyPmQX9q+LkuOHdXJ6KpvfPuOXNZk
AXLubuC5vgZqw8FeI5Q0bvMwa3jbuOIm7YvuR3cEvoUyD8GAi5WHqUfUvpgQ82qX
lrSFEI7QzaQwVd1TOHSMWd6CeBw6CgrO2nonRRRjgC2GMxbeJthMVJWsYfYc93g/
7qB2lycRWTwwWxJgcU+2Deou930zkWJP3Ap1JhDtHKzOJ0AY7mJWWu/QJGVS/BcX
6amvRUdZnXjtrEX5hSr+4dV0RCVOqmJjpe7DPFCg5OGARVNJAAgX74cz42H2S/S1
xV5xqoB1lbM30I2rWQybbMBUM8KpQP8dlORUgwCPP6VVcErQsVmfcymCrZUCQvyZ
2EJQiJNznzc8D7X7YMdP0o073fQsZhXg1AzgXkeIR2vOqtqHsi0zDB0U+6NM1+9o
bWSdglT9yS2n6zOdaHz2KqsntVA7th4r4Rl/SAZwVV+VLazHM5NyRsSmXHh1Edm+
XgOeVobRsD11Fg5LbjGWppYzEZjF9YNDSJdLFmpfQvgPxrne7qOajvISMqYPJPKC
QKI07ZSWdsJVR9jMewYbt5EPJbBTQQL+5liF0LTGWuzfV1rw7Fk6tW7Tn5ifm7yL
Ri4Obpt5av+1TLTdFxVUYXqkWvu53yGU4PD2L34ynwwODPS2wKinuOqiOZvjRD4a
m0sxJPyl53T6F3xXV+ehY4Uhk22WHeMt6PuvCwscs0H5ZfBJSdvwXgf7XIJpThTg
XKgupi9VlYesIdpgHgDtlg6CFqbzKrUWRoAecBbjNi6/ExOiAlkfMrRxsKW30gUh
WuZlS8m/vOjqF/8oUSmjMqR9Qf7g4RlQ8JTecuTSsM1N1ZxwvDRoM0H9UX5MsJf4
jbUlzEZkhrR+mf7VEn+iGipPYu6nESvm3FzwnY1qft7XsO5KohxAgLLgfoQMdhGG
XQOsYplsxEgjfPIi1LK9bIrUHMnCpSf0rCuVVzkRZe+qzTsegLUZtd8eEytWUvPg
qrevaWBDCBzi+Ba/g0dGmIuVjV8CiO3EwqLMeZ/taCLbH2M7nry8cnGFnCFdjQUO
Idj25Y3SmnmM/S15XZ13c1Mwny3xCTiClrpJfmBxoQJsQvkzYyHwq8AlNwWPVaEu
l67YRW9lQ/7GHU3yk7SCNzkYxNn1TG2iSeABZEURuJVTVScU/qzmdlf4A0IDQEat
vzXlwShyiBd2P53T6+7AxLNusVoCpgN0viyqSBD+z8YoQh3MdNeNnizEXHdSUOuI
FJa08Z8dv6GbflEFVwPNUFAbTgqoa1mfzEecNbnAtylRMqyGHNcVKd4ytt457vm3
ihUyU7Gn+PLYqhnn174E/EFAx6H1a1Y+s3aIx/TW3pEE1GflibIjPvC3vlLxDa4q
nblG0hOll/toEEi3syyn58Z8K7LWd3lMQZ5rWy3COT86xL03HJXRA1HyinfbU0Tb
vynClPLo9IhIZJL/fRSM3EtmMQQVaXr/Zyyk9w+bWOXaehlbZY7oHG09/iTmffpl
45ZaE03gCqoxdzE8kpJ9F4SLf8IZB2m+LFW7S5pJzy1Xub3GONeXMO+cypwgp8B3
v2+ADJw83w/thp0CF+ZHLy2PpB6iCg1YGpxQzhTTbv4xRe6APR84HQowP9etSviK
Mz6PG0nymkN11sO9No8btKodXesxJ4OS59rUL2kPlCtOx+IZAwjv+qX04rMc2y7m
1J7+c7s47nRjg9i40kgfQb0pUX4ANWdOS2maQcElHk4XVa7twUrTnbE0M4szyAMK
uoKXYnarLrKW1TLui1oeDKaEJPG1R9aq+YsctYBH4TO1utuDj3XFBVJ/WMh/omiu
+lL0G6tdepy6h8NOtpcQcxSsqsQLuCu1j+kddVpa33vTnNitA/pbXQFbZH+eUevC
O1ZdPiaCio37gmCKGmTuW6O8Fu7pfya5/HJfDnleE7MtRuYTlkSn2yF9umKTqQRw
I7lBu/2vr7EBA6T6B5BTHwUWmvg/dZJ6dHuxAkVGA0LB27uQg8x/ALk/IfBGdnhd
4KwQ59Qf5CBH4lQAO8HPgRx5yLK2ImOVU52OlTd/KMbmz6SosT1crPZpEEcroabX
HYjCqOZ7PupTgdNKB3UUba4iW//B9hRP/9sr2f7I9+HT6Veuill1RyLDtReXPCGl
Ot/CUyouugDL4RPnVL3ny4NQpx3HzcYllhFOrXDnLVMc1HLSzITUE8akAJsFPZlN
iAaYow9YDhLrlxabLe9Ru3k2ntC4hvrZ2y1vsRndu3388wOePMSpBy1gafgQn1hG
+K1P2FZDPJM07Tir85D3SyxVZh3WmZLfKq7jJdVWrTrt52Wsde42bT0uwT6wYwcm
7etws/XRbYAG2w26eRaR5+1/eDZtAE3/NX+2O+rTOAmG5piXRAOMDcvA325L29P6
RyVTjMMxuMoBJYrDPUh1LbguW+PZBWzzrGzd3V9WC3DiITETK4X3Mpdp0UuVlBFg
orWAbMLh7YULpzz8bxgKS7G9HZkaafofb9QdIR+sD307eO5lz+ziJBLdPp3tA51/
2fhk4hSiGopwpDs/TcvcSUxlrqEVn2pdx0DJM2eLhuyE47Seav63ZtgQ72knIdBX
9NEAeNpGXQ0y5CjYqrKrAA89K1HIZnbZaI9IIDFDIswHah/coinPJ7vSB87/PZXS
5sLfuUaCBMXCs/WJRkXPQVFiWDqIqYWd9O2dnTxcb76rQQU2yRGEGbwwzNcMNz5d
KOlqexB8R52BUCKTqSZzHOUvzg75dtdlc2tBH+idUgasUSHC+0RE/9zPXRCVnCk5
AtiVPaH6Jhob5EEaXe7K3v7I0TycnFlRmhkbzNPgqYBdoBn60O6FuGS65go7/GOK
zJoXNCFhpsOQyTzKpp291iouLiFKnF04WFgPmlCYiWbikqaX/0ti0WBBJJOMAiAw
GGkboqzk2Ik1nrzMoNKiq6NiR/8/Q4II+HmZZmDqBi/2Qh1LnUVhxosGq30U/qVi
ymJG9fK4wJ1boTVG4kzg61QOwP52Njg7VKjk+NV+t9i4db21KFBB/xK4VaBnLpi7
n2Qo1bR8HjzFaaSNs5ue2Q5wpKEm6abvBSfzjwluXgduv5rdVVf8N4W6ggo/lZD9
+t2P4QpJ/uGcnsqUuVSPO5MGVEzvtDg/zXwnr2KwR4l2QQYN0OefPltL16I6+Rqk
crKglz4NM5xeARultVi0krUwjrUQn6cQny+3QwBARVn5voL2wVIdou0E2RwSbCIX
Fdz2l1bthstsqSO55LtJ4t437BBgdbyyz/yMn9dtvPFvKpTUF9o/U1eZAt3rZowa
4ahqGC39YmTqst1iKo6V2l4M62rOH7YJRbU0f40owcRR2P5w+Pbu4jqYCKJBv03e
uPAFI1t/YcpbVaP5rjHokJqEkOYWxbcQUjUas9nNE19p0pa9Mh0CiRHCzjFCybwN
leLdgjIjsAof5rauDGC3HpANaiXmZ1YeptK1qWgjIKH0Qh2VRIvpWe2SsOD/FTbS
CBShzi3sh2t+PQx5r9fe0wbupJsuvrfXbWnhjUDmsXFVbGohpAdFeKkHNV/LXFqv
Z+A3T6Mt2n29Jz+8MZCzU4M4yFyaTcBwpPcDdeHV/U/7BpkLeI/VzuVkAMYlYTOc
HlEWe2WrFM2O8/nTw53cxHAjF/Ng0pO51gygkm2sH4QAGVgKKPEYJA01r5eIrsIG
DO81z9GLPOT+gdT58T/hlN8G+4qiB9Q+04QfAs4CJgTzkwP6sndqQHAYy0sC3Ylh
vKmC4ui33iDBe5Hosq64/5gSkVjk0KdhBkALso8GH+YuqPAfpBPlvnvjv3qcH7m6
66HjPtdgEq6pigOoBqfv0NBOZl9no0xGrHxzq1sxPabYTrQcv4aQKMtAOnBM9upU
vSCf/fdaLlIPKJJxJ5WZIot3jXgmmBuX72MnhQkHRyLh96BZCsipo9zubOJFafZj
j5n4YbUUFF13eotOMhy6uRzDsFCkxaVl75Z/+9ilJUx3YWmLlfLAobLx/7ACLilY
/kaRZp171h7hc8XpE57YqskzXs3yj6BCeD+AmCngxjqAVDb2zPaASPrMwz7GgP0D
h9sOtYrxRXCuCD3u2XQ6h90nN6AuIab6MaT1prQu7Y7PTCuHtjcCbF0vwAV5Er1M
JJ4b2dRXxLoVlFLZ5EK20KbAJDGX01qo+1cjE6Z/ofWrHmcmnmcc/iX7D89gO3Y5
2RNZvwX7dcliDjnrsPSM2S18EA9GWOwUEUv6LpaCIjU3V/O+xCP15ToXg/9+BqR9
t7GwCc6wzDu3pbpruD3OGbSQ8yywXNSCQF0ATkS6j8Z9tiJPlCYTD7qdXwRPq9Xm
xD4MLe66lM/5R/ZY3HYcTOrhRpgEX/+p3OKKAwUEa6PWS602ymcz8cGRTpr5PBLA
vtzkt9u8uhxrRAT+Pm2wej/ftj+g9S79VHLq9Qd9vuTC2tAFK1K3FTwwW2IVDeuM
i6GHaNw8dT2RFeONZ5IBHmEHX4CTk8sa+myN2XKCz33TOruoF/ctO5WoQiZdIvNh
0KZ0atRLSRFxMPoFZMpbtyU9IweO5JC+ocopPtCx+kur9zYml1NrnCD07Zp9nM92
yoSEHcxSC9LHEHcduDtKjZX+0kxOgRno5Lf6WjrZkzSN4BThA3ZI4YWLIbPqRbU+
utss0dscmF2X5x+keavAUfe4NMIMNmkH6Tvd/jPoDr7qSxe1r2isyr1mmwaJU64K
LMuMEtZ2RRliXR3Ng0Dp9etb6oBirLKfeOPE2O9qm2lXk5CFEVXnktxxamV2UWMX
Wa10IzMylVOkrTr6FaNCioc9OweL5uJrwEH4JqJABeoBPCyN27B/LZhIG6fnJRFf
mXMD0hL4bVV+sxydRqgewEH8BsNfOIUFdcNi83Zbz8ZKDIVyglD5hYY8Scan1AIF
7T3IPJz99gsnaK772wpyU6vgQAFDyv6owsozXsXi7krhqG3pbvkuMN8UE+5xHzHK
yds0AJiH16mYTc5p3zsMOAJf2S3AcQ0SaFbLslCbMlVNnnSRblWnqH1b9Pukk5gi
5f6Lg3PEN5xZJ4HL1brPXr44pwrOzsegT4+uCk7TQNGzsgYrv7nHGVSnsDRtPig8
azGeYEuzFbGOj9f5m6XjfZdpluc4NWBwLfsTNg9E59wPNr0gWRHtuXA2rusl7SvU
fX/lwY6UTQw3/R+N2hebBLxs8J8zmXmj/15HorusLxmGp2PqO5e/iso+0xDD7401
Yn3oYNBvsgVoMiTKKqpDkPeFi4RcuKzRMO9s38dAhwHXItgZe8ZlVxmCj6q1eqcU
wIzLLgjLNdbQP1YKaNEqbbwiik0Ct1r4nNqPEY+XkanZ0JYmU7asU3JC8570t+3+
IGV6ZaPAx0xfK0K27oRuYjLzVh0AucwLYZw1lqnbH91jd0o+TWzcRR5HJeIu2s8x
DaAJFIjqytP1gfg9kVGTLAxWMnqwbj2jPTq/SSzsMINK9c9VLrtJ/xQiN80ey/tC
fkbDVBzlKodxg/ZEdcct8n9tp4jLTXQYN3YqRh7T4Rjc0v1XfIMFMPltFVKDNOrP
f5VAXzUrG2w0B1tUKU+vcUsqWQ1dA1l6h1UCHg0tOe/jd+RcaQlb+vAGEwVZPPQ4
meHmTG3iyl85bl7UnVziMDyi6ME83kQ4cZy2rO3XmXhIu2E9IfR3wz1yKKQXDhmc
6bdsKn8RCocFl9rG1aApNRSESqvjGkqlASVjPfVRpzl6FYzQZAed949ITx0EQbQz
qI1glofMmwozRuZbKSLmgZp3++liF0l88Z5tvVEUjQEPzd4Pb2kmhyAiFxFp0Zad
fxltypW2OCmEHIdXGT2fm5PxvYkQ1Y+LKC5kl56rrXc/bvh/V2mGtIVvZCvaEG5u
djUCzFu8WQdAzonUpdlG+i5p8s+Een12A3sehUYcgOS09z1mnTbKeHLnoHUmDJfi
FafQYYkuipYU7CUpkyffszAU6+lsssrbABycoSnvHPMHj7kQt9Zk5REsG3BAiCBW
YqpkHcSoa5NYPP+r8gEglb+bUm81i+jv2h25npfBuBbTwb9v0ZhTb+hFltrwBM4p
v3C9BgYHGPXVA6lxQGHyhmEdGDN+KJxKO+bRe7dzI/bIJzOj14Tq9UdrGfjkvmM0
lb1au0OCQ+sjPUOKB0GV2/xM3mrWBuYcsdwqBLfTFVfKwRfEdYtpImc2kCI9VLik
oyN4zK/I0zAAn3EkDKeRGjxmbe2U0g3D0aGGCJvgn8LvaSOXZOLZItq89S6J5D0q
yp+1wK+350KoVwE8Aggb75Xec8i/+6/r9nGhlNkdswoQcew1CnksdBq79zVqEYi9
SQSJhHqSRsCNGVTVRHke95ciqYqOdLkZe5hVigg9BtYSNayFPz2HUtD4Iqe6IPSS
c/iDtP5y0RVUmjpCOBLNHo2iedBCz7e+4qJgzttK+nnOsFpArqMtzmKCIQGG3ZOm
OEEZxiyeDX49ekKGa3E0WcVsqb03a6WJ8OdJCzgDUD5zE5LlzWIpmwxpDiESBt2Y
88hY64pFJwZDwSxUXawVu8H1bnwdNZi+6u4RoTvymWDH4WB39MtF2W74zxl/OEsF
xUOe1J5J8wx38yCrQ9BEO8N0Wik6xJxmrK1iIsAlRsuACqXep5wH/JLw0Ndq+G+R
HL2JIR9Bf45b0v5XYnBAswNJrUuLv+y17aNPeD+CnN4IbU1sYpcAEP1l+BzmYgo8
PQo7surJ6UHpUgTFSiJ+hFYgx1sA8bgYqHE6qvA0ZmBGrYf/w6B3pNgfUktniPfG
b6LKCqLAu/qCADzyhnkaI/G/EG9EVGCriJX/GsvUN0UakYNl3DbuzPDaTud2P9DI
PA7WISKQ1FYFa9aE05imBdjnIBxyQoy7LwWG2DeGXIeinstAdXMXcc2Tq7PjwrzJ
JZ7f1O2EKmgrVLYr9w7j1jYA+YUGDiqXfC8t8M4aeWnp+O+rzyIDEMbFSJI726Vz
0IdYHp/xCrmOIvXzQlyp4sQLRqroav4Eex9QvjCbdvOXmzl1hKYy0pSJzA4DB+e/
8Sw0sbQwNl3ZYHsZW/IJKoxSrtS22LuWn69IhrWi5D4VDmVEnciJC2rjt4YurNit
I4YZTWdmfM1NwGDHxjztz6wDrpIeqPMNeFdCQEmfhUyA6gMcg2N2oh3GFUfHYq7t
fWOQauwqEBlllhfU7E26FnoSig3Zf0wf+2XUPNRznUzwHXP7FJjdIhh/+kLbOFiI
LuGex0ORdeWWcdrqp7fMHgLokN8U/P6wNapYG4n/o3FAP92h6816aCI84VShTMFV
PvowHvE1IhcRTn/htDLpMPBtknfIEpuv9AXBcnRJP/DU/nDFNvPNQ81r2a8K2V/e
GvOv2I77r3dGr6oWX8Xex4yUTWvUiXzFUmzEc1Y/PsGfHlzjG/RElR/8f8tEpsQp
e8QDvApJiRCYfIdAgdDJ/B6CeppQ1j+c91r5y6TvjAkHlsO+5+VsV5I/XVngwdTl
LKooZ2S2fU2y8uTWthNzhZYPTEZFdgkJfPxAMbxKQQJodKLSl3Wc7xrgF57nhrWb
XAjiz6fOy8S0fpq93t0K3Cc6Y7M6mD33+F4BWAM7lWGzofAihzatUDN8Qqx6/gk2
gJV0XTwOX8wLk9PiY52G/HfwqDh4Lz02nvbeI6EIfD8IKyl0nrQ+7kINCsHZ6Kbu
5KdOV0/8PdDmsxUmSoNFNx2VEkDQn2vsbZwV/1lNb3RlJbZdhNfx5e+NgYhwOw1p
Irh0KhYoygkCY2SHtLkuC+nbskWX8QHwdCYijk912Kb35QO3kGqBW8+VkzyE35dB
9xPv6pcuEP4NtRk5SXaq4v76gSKQEf6xOEhyRVxPbui2ZKQvwaBCcU9fIbna5RHY
T89Vk644UgSEVYFHBWcD+q/hFyr5fCmmCBbKaz/zuRjEWcUlvMFdA3sf25eFBf+F
hMwhwicKwFj19P8N4sH5CugKxHuEuXgarx9L8koVhsrBpFE+x4uB50kqJBO0j/Ak
0+unzmfnN/VPclubdPRgavpQLnjaQO0PtdNuxc+aWzg+a4vmMjhzHdfWtuMx0LbP
e/mSoLzBGctD6uXgn5X7eTVQX14qCmGOHOoORLG70LHObTbec5zfVgC78m24x6uU
iC29ZtflWZvpP39tV7w6t0Qj8TWmdlzB4a9PhYR0frHnLquIQVOto4vT0IC2MrkN
PSLoOtz6DHxbDbZtaABTm/cnmfFXn6yDa4jf4BMFv9bwkTRUKBYDZv8nAriEDy+5
8M70swtwL2WNe33VFnEz6HmB9qS64Zc6TrDpLIJEDfxIudzAbxZlQg2yIe/LL0xu
vGZxzPO7K6L72Cp98y/zRpo5RNwN5trYBzrNbp1JvmPcBoufxoLwxwhrsNLI52Py
opdr1Vff/4/HJ84k8kpkmWm/9UEJrS8bfuwkQXPVn0ORPqy2YIvieIA2w2pkVl7s
U9p53sNHMdpR7ft09xYUZOhLK1ZDZzgxBmqVh4A7gkd0wpkFD9VZY0ve3a20RoJd
47T9cNjHCFmw9oYY/2mavn/Nd4oU6TCgxOeyykbelfpzaevYt9rnNzNXcMR6daVX
hXt7m79zynJOnxVF4p6sRVUaZ0EufbNzNc+AJ0MtWjsZjrFzrO0t+RBYV/zO82Ee
FIDRK5+is2w6ISPGye4PAappwV3HJSYErYH2SoV7YqTMcRWMbjKEvcQUwWJmVY/+
V+aJpSnxxgLXPbu12IH+XvUaVL6/1EWBm31W7C8Erh94SXgz9hT7dkU7BKqNAMM8
RDwUU/e7WihZeICHeGVB27e8T+hPyM8fVNyrDdf5QLmiJswS+8Oz84uExl1Z931f
l6HsMCfLDDRJJe7Du91YDZrGxDpYjCPVcSGZhIS6vqMNZmgHh9y61Ejaq+/e/obu
IIiJqPMltA+wh22LHQMr9wr3jN/Hs+G/j18TTKk1C5FBsHwdTypvBV2qGI5uUKVu
mWf2+amJeMxPf6pJQMd7Ni7L6nr2cG1RiPKtx0qNyxaxl96u1TVrjuPsibYXb4r4
dNmhotEHWTSoRsFYtlAiqTRs2uy0Wb3acjQBi9mLJPwLv3dVtXR22YctbmtbLNJA
oYnpmIh2fyBxY33dF21IZ9hoT4a6XNP4LM0zcIck/94pnML3O9Zl5ZiZXMPVvx1w
LyHi4v1RVtelxwS1r/4YBw0wjw+FUzmZ4n/JTL+xAed/++gnZi8RVCd2RPkZe5gq
oV9QlLjbQmzs8/B2f/RE8g9ati6x2qnZfpck5FXu00ynG7Ah6EfvEtaGwrRNtq+7
4BvuYbV7iOlESu4QhMnxwo/GEqkRQwrcFx5kqtTCgwJ3MvlwEQuOI6NCkWh9pGEy
zFGuQTkHU5UmhVk1enxG6NoZHh869SfnD9luVmXS9LmE1XC2Tv+wyEfDvytMACHO
sl4PBprWpqH7XOSt4NJVRO7tnNZYOer0wvsPArhdn6Cx4hI6XQG35InefV/trftR
hmGnVkyQQvvCAwl5imTWXodbnnpBjlymcM84FLSeeEcLS1R6B7kO6WZ0ecizKfGC
6lpAc9a77Udyq8AzR7HgzLdM3gJXqEPPgEWklK9WUBZ22/9Uksg2jQC4VYZejcgi
fShGCeHcvTFJdPAnegtgOYNMopoEKOenOmgo6vlsjLlUORHHVgYj8vKLF75x0M3W
Kyw/Q9GjddVE+YzwIh+rqaRPeK84xKTqDcRpYmBc+h7DjNg7+UlJeHDL4SHuWsZr
nuZGd8ztSrpPZfXgpDMT0xnS9a0Lu/oJW1husRyH4xfD6Vwvp+0vsRTM/5OC3EEz
M8BCecq+rsr+IubkaGW55q5+7zgHxaR51H4oLrG/pdNvo2onO/7h2C/PJAIWkx4v
Hhn9kXTBM4KdJPftgUNqJizI4jZY8jIbrLEEkzTPJIGr5gYcblsVRyT3CbiTBs4A
ve9V6EwBpWR81tAwzXVbVS1LFWnpJs86aP/sAHzJsnJZU6bQsurB63oaxMjlhluk
ExqaveYvM+LHHyhXNLrp0qhbkO/96Z1X6+gmkcBzT7O0T32yEjeTgUSTXURD4sYJ
8Aw6Zmw9pLBF+nJGnyO6Xq38ODXYAD2Uk9/vBw54uLToBrYTvF0ch8rHBcRIazxb
jT2NKS43zRGZWF6skJgvOD5TMXPJ1cguR7PL8TLuoPF/5y8t+IMA/T3kUWHKgbLf
9plhJrnxnsGhJTt4mhF6FXAUXVLj5+Z/ORRYOomX2Av+JAZcMA5xcs+I5xbhQewA
lBox3z1FKzU+H+ZKo4zj1sR754VWnmHiN/yb7Cw8PSSoWPiKX2F9Mtg7ogbE1Lrq
0XqvwSs3wfw3UjgeYTrCQ/t9mNXNeKmXO9lbM8ODaQhh8goMfcpaXNtNHdQOuM5U
IVCpmbQBPWwiyXdmkLYnWf690peew9c8FO/DhcPbQfe4FW0HFbQi+GjT0LmyIqE7
VFeRuxOG9xdhXFfNleitj4MeDX4OdGlSDzRBUHx5oVsvbUYQAjBz1Y8R2brXIgLg
1PWDFM7HDti7yaozEEnVZd3n6xvzvdLU/wD2gVeAc/5n2egIfHviVwh+C+nNr8mE
iPV/2tPjeMVTmlUc9mx8PxM1mHbp41pWpy7GAHmFH7MTlzr+GwbdG+mfixpYwEIT
Wukp8w71x71+vxQEf1oK+amBNI4EgjJFuRepWzkRB8a01fvFHB+AYVfufllg449O
Zwt7U6/sn1pkHneIaqqG9mLlheSAOMSd7Y1Fr9a1weyIrV4qXxT3uUCmsVEOWlAw
/qJ0SQNZNULZmOCIRBEtpeJ7kE2Z/84G2I5FDQkrVRPa5Iv6hl4FwFbgpg5DCKaJ
oFBJ2MFOfMnLpwsnz9WQ7aCvhsbkP32vOcVFasz4ClCHmfK6T5EIraCB3ozHwAS4
8YMWa4QUtK6+OqyGmOGtJor3A6zvVhhGachOw1NLBvcRH8Rbhh52AmrFJcj1Uejb
FEri7eaTr/qg1tIX06bFK1g0xP9QUxxBc+5aQTuF4ZuDNc1Y5FzTwmnA4R2Py/PM
Xt6DshlJwYodduRnIrITRWzZpGIj/DH9eD9NKnbSmyuFjSq+8G2oMKDaPX4BYmSr
OgQ+nRahVvXpMdo443yGS3AikmZnQfd06rZsnn2IbWSpjA53blfL0Myi0qb9XKJ3
6Y1FeQh7L9mlioZpDIBN3iB+vj4em4tfTL8B2rNEF+NBK6NpfSMYWz2iCbrPfCDF
sVEPrpp3vx34fXW0Gc2SWgcSfZ+/jQoW15kpMWamU5NfbVAYFQEcJlrTlEk7sYZA
3VBOo/qeqxXgHiAE4j3FpBMRbarzZl3wg4ZaRAvT8vltpuLEbiM37ccAtd3nfrAD
xWX69iDodw1TwgVlcMWjsjVeKIROjj+vgchkL90iDfty8UkX15yeGPdzqJpHi7rn
INaHQ9LMbL3RMLuQsKYU77vfxYPPsu/Im0oy4Ml/39ZytUCCL0mtzA3Vja6DaugJ
xkFMfmDClHUvF+fQWEN5iL059JHrOXi/jXTeAYtQ7dDOQGKsY1KVHeYf1Z2XSxdi
fQLh/V5h4KgWvqTfUUMTgHiBZczB6xwQoiufFJoeGtXKVdPExCKwFN/GP0/MFL4j
HQIgV3DqZF4PFVMhyouKfJzZOHqfkWPCN8kbQTiRN3daeHTidKOmzXkAILyr7PVD
7J1OEMcsxXm7yLN21hvMgee1uehIXUh9YxxQPXKl80SzsQEebS0hh4/0mkH/DfZG
oj1jENEluZRVGWGt+JcnP5ZujDs9NSwHrycsVQFA89g9EDvpDkZbvM6j3rFfMOYA
Yhp6pP+HoPstGC+QQj3En4OlUM3MFnnA63JGElekuvNyRsb26YXTK9HbVvY38eM6
2wEYZztpwRWqeZX8dSkVPQbx5iS4lXFqwb7u94ee9f5MrAkgIT/MuRVz1biZu6C7
BCr78BrlzXJ+ohV0p1+AMTDY8YheDbWMkDu1iiNAjqRmd2KzxXZ+uIaJlXvneBnx
Ma9gLE5wQMsZu8VowlMk2wJvi9dehRv0EoNfgRgwSO8PcBSK4k32Eqf7iP84rdVO
MblUmmznLATHSsJB41EiMO3GD444B+UoTkiY4h2umjeTzLvIRrX3SSyhDTHDnrwK
oBZUda/IZS81wEoEfF2mTXa3kVRF1qfVSaEXyn+zpeTIenJfzSmP99JeDg15i5B5
E2GMZ5nfCYxUfxULKMQXUGXqlBBh7r9svLONNsBtQXWnyKUvaBoeVJpBYyfNNEhh
+QzhKWBeJ6DVkYLPem3okOW50D1+zdCQ20BJ2H0uzFZEcIc3U1hlip5xDI5Pg57u
UfAkPzyCb8LVkclduWb30cvrGWKTPvGR5LvAmN1YAhDKO/ed4XdR/5fxzqsMvAmc
zsnhsnRBhhj+5HKXleByh6AMuXosSOVFctKnzwXX9CepZL1HCizSe7eM9bRFCpna
3zOPRU1YL5p+I43P24P4GSiTCqYw0+KbzdbdErGSiSGgOQ5qG4dfghb8wBYFZwaF
2ASidP5YA4Vq/5TC9bsOouOe31VLcjm2h4qxWYV+1iWn2+SnrqQbRV+oR0AaFXPb
9hT8n7opoIjxGxfE7qhxth4rfsIWXC90Faxw0OjIpZym0hnU5XeDgwE/nuINHoDF
eEnQr50hzNegzjB4ZCEK1uqnmNJzPHMhEutoynbu55fI/kgSrUdD3ekP+FgQ5GLn
avAKgh9h8BWV3fgeuyZOm9nBBnf6LHW47thvgwwAK3usNSxW4FVev028Vyg4PNYm
7ZQD9DP4MvkDPiGdEi5zrFlJCz7FV22MS6T9XNbrJMq8v5HqCa8zqmSn9p5QPez6
6huziEVzmvbZ9VFbPdcPVoF/zLTDO/b1O19OKdkxlegU2OJSz8aKXCKRIH+oLhne
TenrC+WxLMmvfJZ/9/6C2/GLAMuQ5HOEusuilwTQ6jv2dGLkiqFnHb6BBJkohm5f
jYi5eICYO++ZLmDX7VZ4nHSofeviq1NglKLERQshu+sOZes2RjLJZgcdW+0HTjXX
ZGJaoHQjJdsWA7pQDDTa+4XxIJCCrSqBSKhDW1Kc4fPMbDEnb/jnBD1TPstJcGu0
4661BHJvhXKU/f4bFmNROIuq8ZGs9yuFzCyipK6Ct0QAXfwrj1C/H317r1UnI7vh
sWIHfkHy7xbEh8ZoTwmyGRFxB8l0TgPRQovXVriNE6ZiBZKoHysTenbTu/cWsm8u
IqxsgHYfDYyFxDVvu4FkbovGcUqdAeJzLqY7K1Q4YwBLgOVdAOYHgCBfm2mSRy0q
8AKpdtyqCGprNEHxG8rmuDP+vS+C+Ks9bE+YrEV2NQ+qzjsn831FPB40gIfAC8oM
aw/NNpo+sxBmHtRiNGRTuWTjHfaYW802ZxwxfDWEZjDTM8P/oEwCNwMGenIpbcmd
oRhQ3FZ4M0/lRkxgsxUX0DYaTP0J0G3mqVMwqc+YBon0S1l3WDbPnwMODBiOm3YN
UFamlelr4A2IjJSCwTdBNqKzTJrdkFc/zDKzodcTC/QYG3PazLyJTf4LVef0u7Mj
inOdyCTumU3Bn6LJehqSOiy/CAgKeTv33aAk1wZg0m6PPSV95eTm7F40LYP4IbBy
wtZdwHMMWWxr3hJr71CzA4IC/FZ2ewzsdCX5PfQJlSRzUVY4sPRNNMXrvno/+ONd
xZUMK1cwkar6zZmeCaetPL0keG5IpiAh8+tf+4H4zSszu/rN5v34yPVMfJAeH1KT
ns9xw/pJF8dxQ6J0lm7xHGuxzCi4nfwy5dglSSnwlIxqI+9QggNsqNjqSNqVbpEh
I50Bu+Wxzpx3ygCYFnYesdI7ZwwvjHaJPbim2+DN4PIgthKTbTZOrNN142y3Q/4W
36O1GQtL1dNBUb8aFUFjNXlXkP1qoizOqRj6pWMKwPpBYZrbtVTk6Rr2h6JB78RI
KyDU98iM7I1T1cxWHelpSbp4bKc+uFqaR2WVJBJLu7sERLzz5uHhC33jAHlIOE5v
lAWcOZYbNFmFoEcoJDUNAqJDbfg3YDYdLAYGSjCl0QvptKw1xTBji9epqnWh6u94
1U1W1XSIG/4NmUiVLqX04nn7CF7F0Zu38t5o4rV4rhuS0XcwY71XuLbvyKcIG2Rl
eVGBTpnloDwDlc+xO821eg7AMaKFT0QqLD1Kq0kfMDVJgRsfeTirGbVy5lptpMu2
sOyTNQVUHGwbJAYMkiULIYPLxetmcd+UHkOW1wG+h/j97Ni+/p/0N1ncjVqHlf2o
NgCM1u1LKj68Gt3b9I4jVtnBBQVbMumzyFXgZRIqLLDS6a+7SUfozolqzBzIDO1p
Vy0Bcx3IFi/P/A8yOcp6ktqy27KTGGH7laAi21VjVD3Quz61rTZK5/2DBRzyzhmR
6D/E2SPDMUp6dDcY7K94VScS19qKhqiUBgqv9yxBntbQFaELUDRIVBvEMKDzsncX
/FRgFZN2fDUFDqRMd5hfJ/cS3+IK1pEeYd/4Utzhd2+FLRlkXxPBaEsvwtg1GnSE
d8xDcLPbJ4X5C+NTGlWdlOXGW4i+6gA6j/r1Uynz6UrV0T95kuwHf4UEag9CLxvK
ipdejrN1f+iW1YE+Of3nsnYR46jenKhG0r7DkSj2SkKwoaQaBkIzViuMKv3jZy44
L2YwWIZPu070ddoO1ldMIQ99ZYKk6pqgZ+fyfseSDoGV9dk6Wv2ZePalnBmWsBMK
+tdLIrvfJeiYX3JPmf0uTWUm6vVWJffBcuTOjEccDtA6q010nibNEN4QRIOVD9VS
ldYi3nt1VD4mnVYxBeElz2SrtqFFhw4ZRZSUA5CnFugkmmDvg29O8Eh9hfPXv8Dj
e/QL23/5A/wNXTk0kwh8mtpz29a+/KzEr2Jv0oh/5kbA/c/WYn0/GPy8uEzcjytL
nDfwSIZSL4PWAVej3fLMtZGzqJLrzktA0Sh9Z4Qx/VW3Nbhh92uTReA5IpRsI8Mm
gQVU+S7ck6+o3iOrAxXq6xNYZQUZZRBU4w/oJEbVyo8IEpV3HdqY25U2k9qarnNr
29OK+FDd0dWJMBx5tBQHCOlYeBer1jkRvr4vtZrnrAd8Rn0gaTyY9JNaY5wZqZJM
/LSbHxtOh+wMeDhRJkQ29pPQ0T+Q50/6WJhcg3TyGOgG7U4I6TN+TrsOxhgk2cfm
35NPgnwamiyHzefSDpDInEjR+2rApe1W9j3puoVwShjDu65RbdbPrF7zZ9YRu/a6
IP87skEXKUED5ryM16KT7+phZ4bKYL3xKihxrryfddS3YOpeYIk/YPMiy8eug7fX
bvjT8hFhw7rvnX0woSzzfc+KWuXWYMvh/DRJk7fYto8Oqf3p3XKFA/vtjai8Sf3P
aHo12KTxGiGlRUJFh2dJnh4YmhJandN1qnaW9rjyzdw/5+e1CpUufjFYWsV/bgX2
0CpTmiuyMV0jERSA/Yvf2Jk0dBWqCIlt/yOUfoPQV38XGNSRhla9VOOHI2AKBy84
2KUcSKcR+6T7AjUgvDJGHp3KHVklY/5UI1rgVCdiTBGXho5x9ltQuxNv7eixXA7B
JB5l27QShL2hQNc1jkYPnRz4MDkaPqzBn6rTiPJ6V2FHnH0WauvCj5zq2/PVu7v/
r1driA33PdtWCcnbs6g5Mc8q5ORA6GbqKKw+baNK7EOwxFkfpDtzpoHvfZJWbcGu
NFj4DIhfUBooTl8QKCT85laKUiyx8ljbUjatxEe3dqiGCPRzcGrj0k/tIEOmvWv7
nX2N76cP24CdPK/+H3AhceiLPG0rD8vLe+u6Tig9Kq2qSUlr+g+H7GbiSRUcwH2x
LyvWr3j6nfwFTvSKpgzREaT0j3FCs3TOXo23rLytOGvpC5DTYs/DyyUnXKLwg2NV
AqZcqc1NtUs1KLV3CO5fA9bWGY1uI3jfO+t3XVf3X0TsDTCa1f4xqflIoV87eo06
839TMphcUIWDAfgAhvYyVDAHT2c6/H0KDaK6I6XqVrH4mVLvnoVplmO5ikjLxLyU
5VPw3X8yyhAKCEeIrJbDgEkZPTopKiLJxBMk/8lEUEL6aN2GjHCH8I9v34eHegv6
H5QepsC9vwQZpHnnYehFpeNbj7IJx/NDZJic+ikhDK6Fh9PXSeGSOjOFOno1i6ZV
c+Jttxne8QnxAFEY52UPJ8AyNKV/KlmfouKjeCv96R6XY+GRyBw/mMf6VeyKANUE
w8nAZxElYp8zQ/UYBvwGH1UtpC2xDQ/ITTp4lzgt4l5Wrw7hbufm5wUujXTprAzJ
WL+P22lf6o3I+wwS9JWVtESBJrChypzGXU1pc/2T7w/+sLUVyECuyF6edVIHfh4q
Zl5NDsw76xC/aGn0Z9ls16BDlgWH9ACvcDfVW3Mk1rcsh+U7FN6Wu9TK0qyz7m3W
Ke5DmyO8sB3iFbGun5lrAp4EqDylztXwp+Xwe2Y33ah0DFxlxBVICwcvg5mkottD
ngZWG7zPAiEJrqAdsBpxL4xnwJHhIgqez4LZjsZHymLNFwzybVmiuA6TFGJN/62u
ueqzQKe1BWvqJyY7DtL/s2peShxqIZCJkmBVMMszbatJyqRk0LkxyMj/R7M14UGw
1wfumKQhtYr7zNn7BZXm63XAP1xr2+mmXTstUZoO50pX51N2Poo8i9H1Qk38MrSG
AELvJty6WRERhS0V2AH2eWkF7qcnHmH+eS1kN99NZIG9RVkVyVEFr6bTx0w7vShT
G1MFMJ7AXrR7ks6uMgE/1QzB/NezEI3ZYZG2FfyJ/uzbtprY7YtpnotpvxiwXmiG
oG8GRavNPGQujuKaS2hqo3gSzEuhYCuob43Wmh0xneO4gKGPYIVN6z6Q1AzaXJkL
DcV0pa2M6MZIyBQgYwJ6CGJlYg2SQtZb6WV4PCrBrrqrpFnZ8tMyHPmBM978JyCc
Lo6OkShMp3HxXsSKGV/+0/AQTfCZqGCSR+2/Fi+uLYC4Rehd3xF0YUolQddDR5/5
emM8CqqgVl/GC2ph07UKI4h3QJBBPNpxBTX7PhTWQC04Zwq+uwmewx4M4HabyPbD
mwdaKJwj4DV6xTjGo0ymqnn/7AywCvCLI2+auRAFuC0GVN2JtadtuPn8dkI1FNeP
Kup20XbqBoIQquH/XBslesL2/2nq1U6rbhgZ7bCEM6EVL3BCLOXaRtFEFILXvT7W
CV6qDwwy1qO0+6zFXYtgipoD/WyM0v5XvoYBjVLFOcFF79mRWBbl4XBPAh7hmLlX
gFc/A5Sh1498CYYUQH8udAwg626HChjGnuinAqklhZsjAM0R5JiTrCOZCjWsQw0D
388SzpWSBpAWV93U3kTwM0G/4tohX0uChELIMRm/fyaY/km7MGOq0UJobYjMG0AL
oydSpwWlRdMd0kwuRa7ArHFCpxUAiKI8pw6NVgDNBLaFxHVUA0+i2NzXsv5zFW1F
WvkEMhZVInd0+gqV+RqvwwenIjERoB0F/oa/1TQ6JhuzPWuLtLQ993bjeq+XMyaG
GPFA2AQRZ5p5d1Dh+1XxL138g/5azc3mezrzM29MGE5NLifnavb9YMQF/MqouUt/
hqmFgM1lcguaacsI2RsUVRFOtBPoZPIHNslvganC+8SRU3WxzpDf4O+Dt4C88vlM
OmoR34xZibtL9QzphaYEs/yTPG9VpvYa3pmNRAwPDO1iBi4axK9aBYDI4G3E+Are
GU6QANLsJVtadQn1w9vWFzhbToCHjf6VelFYe8dk0587Kbd64PAerREy55BNqcRt
ZA5eXIeQh+8rNzxpe9+zoPHc8ngJ2B+i8a2CkJ7jz8i/Zf2IWU01zsL5nrBV0lvB
M8qBApReOSp/BMmhT2SuceOekWn8YQSOjDPgEGCo3X/uWzYZduXmXqMQbN6GPfHf
u/nX52v/Ei9RWZbLOQXRBZmVF7dbw851YI+Xu9e498yGOkVsF5QaUaVJP3lZf8PM
dDm+bTjU4pHOJDDCh+cvYPhcj/tWlj83haSrmXHWXvwxEj8inh5CiI8TSR1wtd5m
WuyvJPIjPBe42/IILRt4vbIsjzoXWbZEHa3GHaKJbkWOpDTHjo06e3rrkBgO19za
LPdvNthriaBlGlNaxOuVNk8e+Pk1OY975cp/HYhCUhHVJLoZbpRvKI9g+I9w7D1P
95sWGjys4JWcI6nOwnifZY9PXxQRA0RCJPydeuoMDVBIQGxZGeZookkyJuJxSX+V
AbAsqzjq76U5kwDyy0CXygdNWYYGTKlT/ULY9hYBxl1sRpJBbsBml5NoSv/9k7Sn
r4x8mOWDTUxO96V1psjgkgGVkONBlw3KTqnec0wZVPr0hQA+D4Wos77SbuMrefRz
kY/L7J6Kzmp7Hzy5Wd3vwbrDFyQ31P4/aglPl17/BJxMHUqOiRvthj/sOdJ7dY3n
XqpCrfV+iZrkoYKRZ4slearX1XUa1W8gMduIYjZuoXKb2K5tTU2UNT9snPWWLHnV
72SYGNRdRd7gPwBJgiDNaGSAGw422SnUIVlYxfmIrb6CQtPkQf+zNoAvrnNHusAu
XyIk1EikXNmSF+Fz9KSD4qJeNtvWdSNJvhBPU80asJloS20tYcu5eK++pSHei26Z
xx+ewEZCT9sPgG0EuxOWyRTqsFz9KUXMw6ZUQTcyZhUbANgNFzZQROBOsV+7pa9o
VV0+eYh3kBKV34CaVFC3sZXQczThq/YcKp/ORwMk6xvMkz8VHqWxTGHzlMVvk+ly
/dSxtYXz2bQNvukqfuX5bctGrPhsszfJBhUEkTuROE9hJ1mts5NQt8ADZ6J0rIKT
ddSDqgDep4FwUqEFfynNw9k/pJ5Oc0Sx+SlSaKIiH669DZKo2CcNsZuEth2XeUPM
gZqh9se+epZIxI9vCmhkpPHjR9PB4PYgt7+vqtdwVCw9qqYGkrfkdLQYEDFLginp
VblevWpkjgL/SzgGNWGOl+rmPySqv9TeB/azzYuCbf6IDDD/VIdei6XSK+fz6qtS
SouG5S4EMz7Mi9tiuXTXAZqWcFLL8h5NYP409HS4H1MSlT3kvEmnFHb3fqcN1m45
Ro3QytryF8nOOKiMICvmAZ35j7zxEZVMkwPHCxcsmTb0NvamWpliOEi/H5oQ1MA6
I1OhVlu5T+9qpQdTmGg/pCCgpwVwWEAJQtW0MUK+Ey76wcYeRfIslUUN4kSy0HXh
Z2M2Yw0fFXbbdogoD3W1Xb8gpYx5lU3EHQzz/yMTP55AEeJmkpmLF2UNQJ2IBKCy
uRozjDMoobzfTA34jUUzjChIzMIy2kztlE96IQIci0rP+PlXsOHdKhCuASBcHcSc
5V7ytwmuIUWcQeXhl4urkiZ0OZwkDLLOAF0mVYHl12TLa17VcbwX5tSsubp1SdGQ
Layj1P2YKdHQDVfmkGOsA//zxOlF2xLiez+3xvygd/dYKWG8z35R1B3JrFlLk3ya
xe1645klbA0qHvOUZ8ECjLXqpqk9DNazSq4kL7DZH6JlKTxQoMrK80OLl/37qVsk
gt603U9nB0k4+Vni0VwnymkhP1Pfi2iVjcaGUmcUizAiJ5sTclZ51MN+2ONJQIeo
EYBOKYW3rRbaMxcEsipX/ff6Op9v2PRS7neiB/380SIuAxoFmDnumIrfXhvGymuV
mY+EBGJcnP0DGJjW3Meg8I0XNExeIg3J35rREo/7qKxyOcPMgS6WPnSqZIQWows1
+THNowXV0hzKWvAmlEZVpp3m+jo+U5jqZjULSJVnoHHZGLwArDW5iBfd8irhQkyL
kqeRpT9zGQCa1/dShTMsc/vAcL8elHm92wIQGIRc2E1yrVIcgDZZGcOmTJw+XUKM
+KIODgyiVcT/ojWKZCQH0r6rORN+bCPJiiOap+X/UsRGhnxEidgSSaxtRTCJG8vr
WZzDwF7JkDaZ2sJDLbglrSPuNdDhvbB/c/rhYSknDeLoVdJjQuhRUJ+0vdYclu8r
M+iJW1JYIfV/qDYP3S5JZtVwoCby/+y1RFhu65yPpXizet1NcztVe0XkE1RxptUg
wNtRVp7/7im6o0MQ0jhC4gtDReThPkQuN1o3An+FIjvsyb9/ek+/Y5P1gyIR4UH8
sbKDoUNV9hhkV69xNa5e9biNaAWFdJ6icIy+PZtnlgSKvh1ahV2rII9q+djBDmXd
gbCH/nV4KzYkcNQqZccTMVuHzjwWPsMAtBPJrEef/0y0SRPht0By7DPioPm3vSkI
3cE3POl7KwF+0EkIXeSesNlebHPVBbHN7qVdPVsAWxdaU4GsvZXW7VHQWbfvI1Z1
Iaz3OAEdY4lovYusDp+lR2xzirTB8V1utTmbzcTzpjT8MRrC4woRmmR5p3ZuMweQ
K9M6ZeTXV9bduqNNjt9j9s9ATXSJF/EkFrjeF0nQFuLHXiieQJFBNp2TJPTI0Am7
8BjiaQU7HlN7wxPjnujjVyLSYutvN8Bo3xUsMYCGcUSaGGEelvxdRih49k4T1OH6
D6k869bj26Q1t1tbwxuHPHDzrn1VDXw/MzmNHJwche7Q5gpfjsqmoGwxLzetlNCC
SA1jqp6KlbVN/7OD1FLlp8Adecm/o15GsYvQpIGuLOmGX7f3DPd2VxzA03SlRbj6
JBhJG7fvaM8b/yZEWtYIqTouq0Xy0n4H1YJ1OtPCNho3YuanR41MArImpaMcic3s
js+Qsm1QfzPRW8c92G3ot+r3SwEz6uMjxpbUDBn2G1oWPM4Voev16/7vUu+KlLHu
JCWsxNDsxOF0Bf8kZ/OeI1a/n4tQ2h4IfO4Pvhx7KMvD3BLzlEFmivuEAAUdnLf7
ftS7P9yJkn9rdVXG5MiIzOIs3SWF5imPUr88r7tDstxLca1lObKQbSwdVVzzCOV+
MWgO4zONYMWly5n5rKj1HkYszFgeIru+xyR/d7jO3pu++LOmFijrrqiQPkL4p0nj
YBa/LlvySYLYrKxO7q2Tzpp5XiQusr3tSd8hNAxblZGNIfO+jmPiN06c3+G6hkVI
PSsrJ2ZUk6j9fouUXJEaCts32O6IBkvOa6dGw+JDR6voCbiH3KLSyy1440bWEe4x
ScQ/uQg7YOMO8qHtQ/H+w6tjng8R/2qUYo8bstNMXe2LQmYrabVqEisI5pZ9g25x
7WktfbKclLMSi0U07QxBxePzlt2hwIDy5M4TBK6CvcShEa0IRgQSjHkHlvgindUF
llL3QfexvoKmHfaDstmCjjHdBxz8w4gg/2w7h00aJApjHhkzh87fubio9b1UErVo
nrmZxeA8/QFRvtd527ZASy2JqvXM/JH4rQYpjVuvrc/mpt/boLQOjFt24tOrnRAg
tPZV0yai/zr6LubkvfOhKwvyJCzvtNd7cn+zyniV3DOlal1abtU8QuG9tnZhm2Jo
zaF2YPO/rB0dZRZVOFgrS8Ws//H9WCRmOLCxenQRi/jYhUfnP7oIZO/Shbej+LWy
WbBhUnA6zJ56sheLw+JnCKDuNqZCE7LRkMfy4SmGO6sZ4yjYWoZAZG+23UoVP89G
hHPgCrBs7catXF7GqHuoLDL7nVg8SqjdwgZjuniq2Rl3oq1KRjV9ynfdAvbnal3W
s6tJdUdAZbO4mSC9ayQk1pJO7d0tJlphXXQI1wrjXZ9VbmP2RZ0xj1cahE0WNzMU
Qgu8HFHRSB+B0fKxePNl0hMtjI2M3zrB+V+spV2DoK9DfgtPIvExGy2t5vMBPECG
SXp+PwD+TVndg5Lf7wPSxEBg1muWeeNRp3Fn4/Hv1ps1CsjybvWB/0XnFDwbt6Ti
VNU8SEuduR7Z68gNZwps4Bsylu/Zn40h4jjnQOVHkWZW03aQNUQQ9iTIXvjHRmZS
f1kCvVKHSJDtjN2/PJribuw1LFLpJCZ4CKmODNypDTQu07CfmR/chYVc+gYsZgqy
qQXPWQAyPdZG1lzkSYun7KD2hMY+DAx6ZrWIGC7F47QveXdz9QwKt882RQlvNnG6
18R9HbRQP+QkYNbHkuyoteVe6V8AQ9VBeDLflm5DmhPOrxOGzJJ0G2ntkycqlSMD
Jw/K7Ml5DrVU0PPnOrwCL0wLJUWuZPihx2q+XJjgJOyI18Fl/X2CR1EzWyUNI8pE
3bERxCKrQ7Stwz+1yiMtuUvsxvmRzz3BB/cA1lRPBT0C6grTa1lwkUNhgNUM4w+7
uLAGwbeBn9sfgrj459Xghj+WVgcM7edKsiRhjiY48dwhghjQrxEprRImM4ndBSWY
PMNR1hEUcXiRKCpAfnSHzfOWb65OPlbxek/u9qXoDErVS9PATqqOsXsM9zCfiW+R
5aAkULQeT9HxB4Vnzz3MlY84U0ULplj7xR7ouTUjxZmKD+9dPueavXSHaf64ba3c
EdVwSvAb38NYzvXrHDecTohPA8APE5ObsArac8SAFkT1/XMG2tSqLpcEhYs2g3Xg
0XnZLPGiOvk5oM6cP7n3C74R6jBfmx321lcIdQ0hjy+SteDgCAVl2zRmi45wJJ0I
dkRB3Sdw407u3Sikw7nFGjFZEzrU6KZqDsEgqMpOtQE/BSsr93j/cZzPEUtzR+lv
8rPe5k3k5dZwl8P4lJSaonhh8QvuT9lBG9QcItp3nTsv/YBgd/Amft8lZyAW1x7w
ZI5AHrECVXP+KqaT97b3ooIhDFKfLWBn4lwn6rXbMwTGUZ9B/lqOj3sVhoUO4YMR
bPPUeC+Q6SwUuVg1NHPlAzX5mA+aLrHlG8CVllY8/TDTlSClMBV6gSSJZ4DoM+2w
lZLSFy3mwNtC7nx4AK98tVhFpRTOKPYnuK3+Gq91tcpuLYJee1mTKZ5DVb+siKMO
i2Aj5ZFrJDGeZczTx4q06sWsxlHCt9WPHanrgTcmXK+7J3W0T3q6PruJBv+YOSai
VyFZONeYo/QW+UyPCmlB/RpXT6IW0UHtdGq9boFEZSkEXseEFF6J4t6AnxiC1xwX
TIq2/LICzxe9yd4/jVQo1snUaIJOGNHp0lwtyyTmUCRtmQWYczWuwAcU/YMhH4aC
HD2vN7MbhgxIm8pfSBR0yANqREHn3NbpQ4pMlCb2EEv8nJaBRD1gf6Qb8dxs35MH
F7Sb1nJQZncC9uH0lUYDmTCut9cc3agiCafIE5hXeXgjgsscWHO1KSt1mnei0jI/
TKvIP9SB7hXJRe5v9qonSZe26LuDoCgJzbGmwJj6BXGTDRccsK+LC2g+eTb+uYQ+
DnsK8fMj5E69IdjS8XpXzqq2bYjbRQDcAFla03KlNjzaiVXsssTNoP37C+de+hfQ
Pe6laOV1qS53FWGJdWOjJaJ25QMGq9FvFVvaYcsL4bFyiou+S4d5hsKyvVbqR/tP
5h8jnGC7+tC7aUx4Q8pEayeD4nGho5LeI3HUjZ/ZFMoPUq0K3TJrlf6VfvdMbh0y
im3MTCbzkb/1f1W13qcbfw9kXjWGyY1selu2IltSTAXSoNZq6RbpT7Zqzk3JnPuY
PHd0CCeRZpd9Ronb+rGDgxXwC8ns3qysHSGMlViSaeBvt1f1z6NoC9bvVrlPkDME
pC2u02rf3cwdtkRI2+iOHskru7enDxnYoFpKm1+k1rj2kTNO//PJ6385Q0JLBa5J
PYnCjxDhI+CgVAUEEgr4PObXN12qE0gKHTeE0t/XWrGNjcMV2e/Jbp1we7qUBdVX
d5vhc2T4VRub0/FhIOHTocwiV38eYWhpGAStMJ+F5g920F5pWXSrYTWgE1YBfi+k
qg6yydV/gCVBjBxr5riPfxcEcFQnA1XifCWPM7IZX3EOMergat74LaYZ9tAFI8F+
53cIPtSlChMh7e6OSBHtghh6s749FsKzxwzwFrJIB4f5ehVabm6YTakfYWSmvTRM
7tTONOxrL7gFazrcmV7B801PQejYppHJK3iaJ6uwZWuLeS/o9hcP71QK8OEopvPk
qi8eW/aBZBjWEnq3ABqIBoZtahlKX45wOu5hdLQGiZVTTC5hjc9otOUKO1dt9vGl
EWU9YVk0dljtO7pMcbIeIp7J4SDA60w2XcXLj1PPARxdjHVPFgzzIf+Z8jrAUY0M
otVUn+jQrsUec8Pzsip16UyozQ9NQpImWRVEL5jrSmgxSza1kkuMF5jwmLXgFBE4
owp+RyYUFS5bIIIfg876o7P9jBgEkY6g+kM2VcY3b5kttK1kUBiOPy7gys+yR3gn
1/EzrXd10SFQgNfaEnfBe9TXaFVMLnXWqOzTHpTA4HEz2B+7F7XxM4W4JF9V/+MX
73sudyKv+NQfW20HATM0mSRrrx/eLviyGgzu9l13nOe3ltIjN0mQVWqNTEHEEjNn
zDzWRzsa5SGBNAB82VCUMw6kwu2A5ftW7d8YN5LUyxdh9MlrmewnMu5+tqp9kYWu
367wj6A4W6LzJmp57MIcoup/wBrTpb+pYguCG5CxBawNm/YvFri+UWHy6qPt8RRF
c82NwkQi0quOcBj3Qo1CwTg2R42d7fvQLxlkiunl0t4FkaKOMIg5zHA8SEGqASdy
901bqZxNltRkNehoqjCBEJjAl463xZf4czxmd8/73CDvwp8TAUCEtBMxxttKMK1l
ZDhqV97xURZ0WgTQOB13DuHIfmSIzWKPAilRElfuunVO10sOHB877jg2gpqGjQPE
GO4l7ptWElsWIzG6ahfYi5UjeOk5jjYPfJzSrTw8ufqNyqJ0q9abX3Cjmz/pTOqC
s9BEf/jMknr7lmP0LjD/dbFhsmpLAN3vPqIAr5cbJahKueL+GCiDK4CY60+CoSSu
ekxfSgD0qy7OEZPNLMQPzebn2QuBmkXEZVcwwJcFF5ghgLBUC6R7vN4BkAjXWU/F
wp5T322/ScT7dB1xJ9GtyeivZcDqcbPrAjI3ICAeD6ETMXTEXqylrnDm2+Qkl2bV
5FWRjGUn9YryDvB/7OxT/YefmyE5c8vUFHg6hGvA4UuvOPSSN0MB+q5BNliFBTuh
k9j5kuxV1Ys8lL8WNH82LZPuiyCfy22NuhRYH/keg0o9UYOb5VFX2IPymp4zDoab
TyaNn97xg4sY0TyBuFGBA9EEzRYYRbXtvkMwtadrDTmnCx4c242mIWVDSTaX3rXg
3zUwRvy7Rqv+nK9DMbkLk2rOXsv8XiJIKpafchA3iikxFWD83mmoXUYk1P/0KN/t
imLckSfgMsHb0ylI6PZOEF9CS7IEcpmX3XQtJEq1lF7ScS+BCHLTdJiv8YvjUxjZ
HgW9iJdk0myxBLjJdutkv8K3U8btGDz9vX9wW+iQStFFeVjaY8k8X+rez2FrEDqT
gQT7iRIfx0rkzzkXFhY6A2DGhfVG07gOusCjjaDlAkRpdoWeb3RL3vmmAqrxu1Vp
J/eWgeJJVB3gczJ3q3qIKemcrviLKzvmXEiRmS6JLKEHRebpEAYypfkHbvFj2z9I
3lgDbnq9D5v8dxDWUBE5nebUuYPzyjiWFtbXXrEgzPz1vCFXFUJ+wfuo+scnu+S6
Ck32FSUYqZ/A/0Y2b2elHLSfaqFIV3QZZIGt//MPsrTszpBCdVAb3OZsOHvwgyK0
lk9BWmJE/Mz1ul04zzSNfZum2IWvpLS2n8EjDhCnQ9YT4Pmpqtd2m9qFb9mHaf4w
xp0UZJETUQjAZHcR0yw3QT2mlCeU1mJxlGyN446f4pbz7H7eOAjybAKt+xltC4hw
QnTkgo+csyuU/wPAAQY+bVIDHY4EWSsUwJyarXhc9c+NOPx17Kp8WoG7HVDPOaVh
5OXvV82AEM6H1P2K8RDgEesMELt8fMLEGeAXpONvJAkRXZui6r3TlWXZq7qJdk6a
FBSDwqkiRtoi7N8MYmcHe9bwoMEUqP0CKwcN11YmsPZpYqT3mjhiLc8fP4QNS+hy
jV83LNcupFS5XSJXcBah3TAbkixPlYzGXYvq950NXGM70clODfsNhEJaxtygQHKL
XX6X2PidxjsKlbZwxrWQ0hcRMyHV+Jr+jCjm4y7xHX7/T50sPW8mzn5rrsd6hx14
NwGeWr5A3TXtdmxS6XOKa0t86D9Vl3VB/0GI35wYe6swQ+z4x+Zr4qUmWt/8Tzvv
PSMW/0lh1QJ49asVpOdz9pDdk4kGFaCm3dNoqvpH2Zr8qelSqCabx2tZSQoD9NEn
9CVXV3pnOIrvPjLYQHjjQD23zj7hy7PJfHMktS4eQAwkky6FguYsV3bavgxwHJHR
62/9W4tfB2tHnZGDbv1tyDG8L9XmBz6XMZxYAK07uIcOk7ItgMFb8ZQ9CGXmavAG
y1tvZkNBoxydXmg269P4cwY9jGkSxMqybw3nYXsFTUpNf+MgvDpXGmCXlg8W99Of
k06xB3q7G2RsbMuMFkU9Dx0yLpy7sX61S+esdDnHh21Rk0asCkzM/hpMF3u6sx+Y
dLjGIEhte7FcW8PzG4eH3+afH8JrXtvf0aJe9GMGL24ZVn6X2NfrX8ywD6OW2XZc
WBoDi0czDv/BTYXoQp0BB7/Irfkw0KUbRuTA0hoEf3ZpI/+i5p16jdUfRzOjO7As
PBuPnQPVhWBK9djmLuDc8vmaiUbw0e89anx/zsEDAsYpNa/Am232GkB8AiGiINT2
O9uEzSoGLTfi/2i+X2qq+htoU6JaoLqJM4qbyIPz4rQT6LEU5V05hT7uaBAC9q/E
1/OcUiNuRprV7oLc35bBbdoZRrfRTnQl+x5hf9V+gbHTMhKbBSXYqWZYDvQ7FS9L
xVzowmjt1zCiwsW+4v1T3uA5COwes5U5tmU6jEjpw4+f6RS6a368E2vBzrNXIBwl
xL8ODYv8cE+vtj+oIkgp+2kCgK+UBmXjNZX+k1psid1YKIdDz8HoORWXFlgPMH0I
T1qUnLbAHZyA4VSqLpwXsmTttueAMVKvv8MfANKL+MWtSoBwuWkPIIADSuR82fgy
DJ05QHf/Rt5R18Gr5pnmz+0N/eimxslCfjta3k26PC07uyzqlz+4VqdRODDqejM4
+BWB69hJEbx9WJ4q1dXU0psWf9llptdIHcoqQiBxGRBr66icF1PKkZ/wu8kx6aVA
6QoIYg2gkQfrF3lMmw3e92JLB/YiORVedfz7lFGCcsMc1ibGhVXm4alJxyoysmok
TlyXcoBg7Tt+83LSzH7HEC/R6UUygXTKzwu/1Um7bzE0E2UqDTrYMmhiOhTHXBta
/fJqBdPSX2ThHpgzsUwwyqy+32ZKCWPbYnifRFA+nYDv00Sdeot8V8gSWGCoQAEu
ZYJeW2Ic78bIpPykwsvL4CzmJIBnUhDMx9lMZauvu6rNlbkOpaTFZILwAcrztTfl
XaPjBAMlohj0XY/x0ny+tGeEmJhUxMVEHXhUr28s/X/XYRc1SdnMZuLBDdZzxDUN
+qT5KM+/cjMKDhTwD9m6RBlYsYYzmKwtuZMjHE7dPjgvG6XHDkYC2EcVJxd0j8EW
IQ58Uxs+ae6P+lg6V4SP47qKR/EZD5mS9LNM/zn27ryDjipkYFbGTvz7HcLmO9cd
MCpWi+b//K01hd+pWKyreejFNQjPWXBL0M0iyxHq71TlfWMKLkO6FfdJmKhpfMXa
bev8qreyaKKdOwhTRo9hE+aACD8mGG9NAq2f+Y52DOyZYf/vw0M1boHs9jMcjstp
adIG+E2P4OD/vlKw+HAaJ1n6sM9PREI68yRKHDgu0JhugMPkfOTcByFHCfBNXgGC
x8oQn5Xl2SGzcc7v2J1NM3nzUF6bQMPgWVJjQClV1MpkVlGoOVBYga3HScfhE+TA
5shCLUFh8l2zUaYxgkX/otKqpsEVCR9djyFQlAcvdKyMV7rswJ7qpEoJmlA0khP+
/IiDL1euHHhS5b4x3mEzEJQUQpEraJBf51LcLAjZoWmTmSfp6uVij3TGPBQynZ0z
0/DGKc+UMBgX8TD1hLV6L3W+fkvB9HmuAwM5ubhCFmNDILrOm/jlokBerTLG2jVo
Ighm9GpwP+OgkhmwGohftnp95XKF1lt0pOGGpOqM5Lo1uZweXkURADNRgWfHCHAx
yQ8wltJl3tP8voIt2a0BXKUQuxr3HlSKUINC77pPRi/zakx39MxK/iE5Vb1krYAF
HOGNfVTQFq184xtF0K6uYmMdAPKpHbKAP03m9soDnG7HBeuyllYK6LzkXjpXFr+Z
U5wavAC6dIC51LYOxy/ZkL2xwKoVXYgS6H+XWLmNRRWYGJXp+nZRGEZO/K6ocCwG
Qr1D18pAIhlnawf/OBWpWYzmP+ii0tjTFxBf0x/srtOQEloGL1Ps0bC7+h4XgjCs
X17qfJXdHcHE+jemk+fw9dATDH/QaCxodHxy+OP4HtUo90GtxkeBDsQ52/+IQ3yP
3hoft5KCQT0tl58owMXLARBBGa63f9z7VgfUNTbFg6t848zMTNFk25LxGbsBYweZ
fTfwZ0/rdYRPOhl2whl8Z/hgzMvobjj2J32nl97E7htwx9Lj18AApttmx+TVxJA7
21DQBNh0tD8oRbRMFdZXkvY4c5zIUkR4q89rfcXLua6Dk6x8tr4dd29FL9XfRR2d
ZgIWMn82GHUr5dwSo+JBtn5p4oMdsN0KCGRkt26DDtu+4fRkLFYXYr1SWnsehNE+
dCyLJl//PgMSzlPgPIFnu8y9Myth0LdFLxLsczd7gSFcuyP3VOjHJpqVnbXojJY/
Y17hy/IkVYuaOR2EWCINSJU59qyxsHRpoQ1+1HssAs+imHC47a5ZMBgeKaB2PVDq
R+svAkimRTTwnHxXoawtXLckjCG/tIfVvspJWLeJbV3NP1gsg3o5+9j4WfNS2ir7
/kdQV+v3Rya/tZCG40OevoCTESgNwOri8gaa5PJepARs5BZzGhAmvoE9agGPO+FP
r2353s6hb2A8uEAsMf1YpsI7kpbJmFBpz81e9zBTe8GVO+L6/dqbKGcxUiPRW83F
HIDxrI/CsZDAjEAgWtWDid5gn8I70LegFOjgG/Cyb9bysCHOw8KSN00i8OJgkYLB
c/RsypFsIAB7Fy+1qDRro606eRzXTqkH1K7+4ztB1BZLnJMUq3RjQAP/pbU1cz11
7CKDMadcNGrjlJeDNlJ3N/sMvh7f6UdYE/yLDHgq/WCVXtmWEqfGo7esnsTLkE+Q
Yl7ih7GqNcUlLwKHgsRO/G3deQpmbpM4bB+i8QRvrSlKLUr3sbwqaYNuAttdsT4L
7woUYtH4CmB4ogDZJoIijLWW/TIze/QVBvoHHy5HFeDvf3XiofBaWrEOy4kZtCK6
qAMf1IgMqXY3XFGhSeDXOsNBauptN9u3zFEhevS2sXURVxLushbZxrQyADUh/MrV
+66R6CoW8AK94oM9+Su3jo7PQNJPDqiVCby6veVLDvZ9aYiM/BKYeLYbDiLYwHLU
QNP3DWdICtZFeqh7o7KvBNsFE9lg2CeFG1lZh58iLHyYuttyeo31kJaMib8J3XwF
n3Rx35r8wPMFHRfJdhfy7GZsBFlTutZwIMhiUpriqSotbQUpoUNNitzKJSGSYQdT
qMmHmk9qHuKhL6jiMtodnemhlM8+4ibmGdDmMvfI/1CkPEh3WFiQFcGM8R2GDrUy
QYjpB4vpf5K8DlU4RBGzgx9OB3Nwlu6ytxxpSkw8WbrmZa6IeYyHKwudXQXYUMaW
YAvDgOY9rrpo2/bldMUpVri9Y9FAmdixr4oEPfKKwIor5ieDgcu3RR6MdSTedOdh
8YoQ4RZNsjMkZ+Cuuo2htBcreA46tF3WKZuKUD+LZkvXzn0ByTiJ1KVmR8B8v/2w
Gqdopmay9mY5KWl2ANnRW099geTdiS1KDfXnkmvA69KnCc+VMZw+R6HMi/GS7lm9
DQmR+jbQ8SPriPkNLe5zDBMviOAwGfYxNg685SKfuUkJcqcYukVOsQ8aUq26WveK
eUvbG4fqNziV2mBHnPF5lyLTz4gZf5d6pMh7CIPhD0lmkDDcoN+Io5jS5Q/EB61K
BcFNMm7wulVVQs8CZp+e4SX6kiIo0kmZe21TxWoNYRZlK7wPlbR34upoFaMQFm1X
DaqmRRij43fLTsCfdgkaJNUqpP1/zXAEPy7yeRavxbQvfx0mzyPHBo1sby5txbTu
SutJKkeR035VwDT3YFbw3lLnUdt+4LOeReKB48btEoG1+YryTTBncObB5PFQnrVW
8LFUado9BqhjlvQ9eekI09YhJRVK+v9s+E1iUPEUMBGgOkE4d/T/Spp8cm0YLvfm
FpxG+Zc6K9Q4zdLC65Jp0vlh/7r4yn/5xLN1zEiB55ij6LtzPPqaxYE881ai0Btp
PyII4Mk0lIoNrB7qHWZoNvIc4y7CPr348+UTK81Ah/7ZcuK6nvPSLaevFqEPpYzf
dfed7iJ8FP/i0cPs1bqCUsMkndOy+P2PTjwrPttjNtsQRTsT+K4awiUQfBihDq0i
rFt2vN4vimlVWqwjmQYfpqLWBweZM4dNU7QKEHVGDiJkMJ647DCw6WWHoVZpmpsC
1bGI9m7++W9mP504bvnhYgE4Io4ziq4aazsG6QxeyzjXfpl8qergndwknf5G+JbO
++rgYHZxFO1Ra33nqWn31/sCxB0nUJdUcFPJEC+ztUaKC4nEu/qz0q0s6qyo1tL5
RgbReSkucmFXkDbCVw0xGBYiHlz0yy+HRlrzHa34NiiodxBNDiMEJOLxnDA+F1IL
VoSyELLwBfPyhyTakPy779s6PoNWd1I5TFOXIKHrSpBM9Axc8eUUgoHMXaxpL+5F
xyx8+s4Rif6PVeN7eVC5W8PRyoI7hy2mOqBnzGfJzUEniFDFdqaMbJmEmuekrkd4
xvKckfYmqB9BtOLSf7wlcznw1SbPbokpRLP9+FX9LRgSJmpDOKLEpijpbmgeHa1K
AlTNUcNtHaR31deuDgFy79ORVKQ2vP8LJ/NimCM251STunsKf19r4HH53/afgCqq
jusoLTmEhzZDPVE6+jTL9WSlCjZyaFqKOpk1cl+6a0VZk9QKoqhNNLdLAQCw9T7v
8Ia4l3Yl7TG+W8NTSZ9kRd5d/ysf7cr+pI0j9Qhw3tj3DIXRMmvub8r6BL2pnM9t
DnWJ6Gue7tdgnu+Brf1tfBcViKYGMc8upymh9Bnfe3vHrWBVrn2c183E39quJfeG
/EJIEgKySR2deP6RNVP4+rXCOItYp1E3/uIKj5nLHto6YP/OQDEydrKYMq4OxX4L
b+QuibSLOQ55O7WZHze99kk1bUgZ3Qs0Vh/Nx6IT5kqlc81656+oDZbwhb1lGyhg
tG4ZoHLs7J3GGkY0+NAh0b7Vhcjkx5YSTNV/d5FrEgf88HLOQuBD4ToDtfOUk2zM
/dZE1CWZPrIGV1rgkxBsmOQ7OeAkLtoestTnQum5Ho5VhZE1883Qmq9L82CESWDT
60KPq/TDoBTewf7TNK1i9a7y/giRfI1KahT9k1a8Ez8cWIgmwiQeJ+b3a3V4Pjqw
0VPhYGu8VMWfCTixoU44LAcz1hGdQbs+NGcUcBiJWSWGyoxlQ0EwEGXkRjgfh/Gg
Zgw0dqnt4SvEMY5TBM3q5bsg6EcQjtq6GrfQ+WO0WBGsKnjsccPxddyuoSkTcsN7
GQexgrBsTc73OskQp5D5xVB0Mo+N8MurCxi9ClHFcKjQafLLMVS4KZOcWotcvu+/
CidL4RDayV3+m6i42umxdd6xHC7rV13QTRJa17avVztXFXYCTeleFskStBNjkejV
3bweActQM/YAeBIVKshecgYNVR8/pm63apmxiFlNMHz2/RUtSyFP1kbYqgW/Ooag
Hj8BO+vW1u6THIYe/aA8LDxocv2FuIm4fHUc3nGqAPoD44BcAcFb46RdZYZSksjq
aItMANqxMhjq4WvLJsvbVoPWuIo3LuhqYEHueoXrrAdXCzyaRr52T14m7MLjRSAW
1BzpxJUt78Ppn26xDnezYnKXHHUCuUE9dL2BLEGscK9vy9mgtyMxBeBTDD0atB7h
9USRuUjbqs5ux0ccNdfMoD6aNgnQ/0uZcIiaK+Ys6nFLVfUQ4velKbgVZhl1coNt
BP9cMuBDwEKgIP7bwbMRt/aX2yzHO0zQZx8i8l1X65D0lXQxDMjpsdb8Jj46vC47
HVPKbOU9qzB20UrCR/VHA1WFzBr/k9rrZEQUVq3im3l/4dP3btgX6voD8L4nKbtb
Km73bvdNTRkZkdM55DtkhUU1Kl8Pb9QFV9/A2YT07M8cQuZeBj9ATecdFma45ZRf
6vAicFXp+558kjPWToENnMLoYwqiH5C0UWo1uxTOaV3H/BmWUVtaOnhbXUpT6lxR
103ZfYo3qq2hsfY7Z/xtVVVoqLko73SgZQ/YABirLyB+HA6NI4OV3MOe5l+SjafH
XcQHVlBauo0OoFLs+WauWQAvOEUQbnRAaRezcSNZP3PxbGqc/QcOjpzz4qz5M5i8
+/9JytaL8I15iFljzsqbRYQdYXZcsg0fqjgXU3p6uZlrlBd6l0wZ3q5uN/CoTxX3
h8nSuyP4i2cIu3pCS7WLkGGQ2zY+OAoXUBMJoo3HXhJMHgo/nasbazCYfCiK9o2p
4A0MnEPiOD2X4ueEJTiLyRZ+RYs2qe+/YrAqsIBnG56CtHuITMOHtl268HSN3k5O
FOYzB/UKvwaKzEtAa0WqJ9hGPbt2Vep+0JkvuUabTKptPm796biqlVRl8sVoHO4x
wchwbtbZvhOPYD2tB+24OuL/bn3xnd4UWjLn+QxwOnHkCqvXx6OSlBqKSXGdbzer
s6aqDdbVoK1tBpCJIO+JB2fkvUDLsRxD64m7B6JwzuptOfRhshnXtsfsda55zqgQ
+agw8IVxyUjJpSc9JQJDDq5tgtCm6dm1L+QNH00nqHril5yPNFASo+8vebBWdvqc
CD0z1NqRpPpP3RlIkn/W8zf9k9zYptHdbZ9CrWr2gzWBPHW8HMsBe2Mhy/IROKY8
nLwby9ur2MtOIFDN2MVrOls2QPVEbYJdPfHZW26Hqo6TFqEp5cR+BtF2iOL8u6tW
wrkzyXpphvXeb6EPDGRfuxCNWSjayQA75lc2wtIApWnNOSuSVnaUBNGZv2QcOlFt
tJcDsn04TayOFB3Cpm9Dve0hONG98zyWrCP1R9CJmNweK/DBnhUyJOMxs/Ufqb/B
llZaVYv89+LmcWKav9Fm6zyIS7RnGM/OVIE+QJbeSSF3d9DFcIgAKsUQOZCL/Uyo
z3nA4uCVzMOGH+bALBCtjdm7lmWH1RP5YlifOmuIs0AeSqIrRJpuftnFtn9c5HSu
jt29NEc6+uZJv7F/SkcL+/RLnKKrtMosu5lbtfKMvvOmBy9KaxDPV2UCOuMF7YKu
5J9nm/4jql4B/Bir9Pyff4XynJHgMuXOyfW4BxTutP+ZqHpO6/ckMQoiNl8ppXuJ
s/fWtu6i3srGe/nWMVFUlWF2Bm3zGQkXRcGJ1IPxqRYYMVBLSmQzeaZDKqIZXXiV
YZOcS4l6wL32kon1t5bmIAAO8f+wg5FUVY9mHSv2XayUzEQiiMS+N69VjhIXqsIB
ei7HOTk1m6UcE+hE3qROvZStby6Z+WCv7v8YAn0YQdKsfze8cvfxjk0opHKqtpgz
XxSlkVs/dUdRehjOA4HYkswNF7wGUUpKt8ZbHogn57HUORLqOcfHkrirPJv2Pn81
UJ847oeSN/BBvxm6S1bhpruwaheNgaOCOjqoNs23iAy+L8ZLpZ4pmKRcNezZ993/
UR31K7R/wnLisSO39WIZ5+ztPL914UypfUy3cyh/nkCRrMY46GyDVCkHzF0lTAsq
Kedu4cG5wuabS6grMcajs69HTXkax7+LV3vTMK/cbfjsU3ZWzd02dsgKFakW9OPO
7Zinko+xiYCtC+dJCz7UX+8pP4vxCPdIzv+CJLRMiJzzxjeeZmBUJdp0afoi0hA5
1Nv542JMy+DV/FgvwS3lrznNprxMU8FuIcYoH5JLCJDTsHjjlv202UK98arptFnJ
cqy0OrEx+sxSSuaPAeoneQxr0C/pwquYW3YPCxRfVs4Ewdl0k3f+AZZW0Dy1rJme
ltJL4jnUHVs4X5+QNOEac8dXtch7ZF3iqfA6oPPR6RcyWe4rE/au/bd3LF9qVXcV
UihkccF3pRuNtEGLfrMDa1btd6zMic6LU+r9raeTibItaRsMJ/TPB2inh/vguZd6
vTe7nsHZlfGDvqyJCKcOhxT7USEllT4LGrUbppdWIZAI/tcABInNzr0ntcJBYcPG
MV8yuBpMDBe3EVx261MX5jCxDAZ2gzXsbOE8DEmu8UJ6XbLR69EI/lVQ1iIOE6bF
DlyXYRbTe60isFxGArZLdZgtLQi1H1MJ7J5/OR5ub6U4bH31IJqIbpvQZtkD2My8
pzSKKoI6mWFFCAisanbtsyJoyl38un1AHNU0jW/n3vlUmt/YMy/h3YbtEdQTDxE6
57dQZzyNOEMXw29geTCIlYJgi+3aH/eB0kF0NmYhosxRtGHimacqRq75Nxzk6vPZ
V5AQRsG5HblBNq+uAkcztm9+weL8LMfEKU0LylpkNKdwJ0nQAia5choW+X3IokiP
plAh/YPPy6tb1AnWmRpDvTHCjtCn4m6uJl56Uc76DthBB0zDtycvDAlqbk2YGRtD
3Gi8tcZi3kcvN4FXs8ktfQ2fnEeJrPqQKhTs3oKOfQhv+b9uwFaoimesrOevR4rs
SWhTxEDChB3yC7YhWgBl/8Rl9KqzjLgZ06h/G7QBKXtpPHHRmm1MeXzLYeifTlww
UY2osg+eyqD49aTFSCRtB17E0ktAuU/gNaX/lJpqU/kvDIqcgQ0ILwtheN271pc4
fkxshpr0xmMjRqfyeMN8EdtAVsxMqBJ/G18JXTWPWOdeFmsylmlXnyX+w0ckHbF7
mFUGUlBe61f6i6+bai6RiDPHebWs/REoDMZZTNgUoOKMgu1bbb6ArnbBbKvnHNDq
o0TFZlwv5VVh/sKnFlmZM5S+hDyHuVV2Phup2a9S4DoRe66KAzaaVRHCpnyFl/dq
rDUNptzUnvYXS14LUtFTUTw2Xu1zNKQdN9zFJiIy9vlHanRmVZIsBKYiOT4eiD6f
4y0DE8uZP/VRcJJeAVjNR2EqztHBh/wol2pORaHS2+g+i2Uwo4mxhdqhYTffQJAt
EP1VLSUfdqz7wo82uJLjesbry4n/htnn9O07s2QP8CBz53W/7NQHFtMwG6QOpOzh
VPUhI8ZqI6iIapgx1DzeHamzBew2XZsK/v59vavtMCsmiOcn5gW39F4E1tMn99GD
roziVDv/rRh7256alZJLmorsuEX0hY5XpIbtcuRTD1M0xElhIveEzJXeydHlWhFX
f19RLAAa1cv0LCw/m2mzL/EAl0ROX3VL7dOe9UaFyaQkv+kI8pkHWYrOirZ1MPVU
ISalbvqz3wXiMSwK4LGTP0HV5smnPgsDde6cm1f5bJeIdGMUmZYAtW8uh+jL/XtG
sKMIS4VsXD576ix294fUisY51gVqzCxTuqbiUJfCqq4oKYGXMGsLKXO9j9lAd4yO
hSy83IrDa9Qz+uLKISGZgelcv+NKMS9WezvIKtMpReyneInNg1dOwsiFjqzr2lih
PJRoO7IaUa7UuT01mOsEf3FH2HTJCv1WjIoWeTiv0FCE80oRfOcW5tDYiq5n+ZQB
LLgR8KM4xk7CPeF4GpYAWOJAxF/IVrIlmGKsUw5HxL2as5cL/JgDfELdGuvgg57O
bkEBzYBBH/QLXtMEu5icYn6fGKqb0CRIYlBvPhHsjxwKn1JKONt+1+e7hKdNE+SZ
wQtDKmiaLdVIcIOnEQtCHSDtrbJWc1AMbBIh+Jq7yEcBaGFgm3xEuxOpOn+aywcV
3nknGR4I5CxaXRCMP+UogFGBk3i3nNlmzxSGgtGHW7UlbHJkJ7SnMy3BGq2rE2uI
TNYGB72m/3HMPe2oMBmvTS0FmMy9cafI9HQom5b8jpieOFoNPAmmFMY5wdOQFQIc
y2wqCk08iaO+jEC0P89KGl4+B8/CVgsXifAKoT1ygcQliqytATIYRDpUKpyQazJh
t+ETQkYk60fwfQhOIIchpRTsZxAFr5jXDqWvWzv88fHN3jSK2Xma1N9OwgmXAeuH
d7zD0WwsHqFryPfKfOn7NUlb3zVj4pVd9BRzrc5p6gJgwWW7ug/MpfldaHbwZ+JN
Dpm76MZH5eYWbN+lRzI8w+4xKlYsnt9W72PftJqzIPU2kCDH2mP7SO5MftT+t9VB
dTmbtDpgcJbGAX7QeJW9xubJTsrXmjkT4DVPG9SagP0uwUYT7WaeptjLuI8TWDv8
S10Sd89Y07OIs3et7ooezHfpb365UDAK+hLlkv02VnphXuvcrlwYL9E7TyYVZR4J
DgrjnLzMj9VFhpIdXrmk2qfkljzp9haVZHCijotnsT/+iXmklOhpII783mPdwVHN
jBfLDSyZ3RwrYLOQ4uhbIIPQpT6yunL+ET52uBfYByXrJ4dzZwEUKvh8qBKWrN72
fVq+doKjHwyxbEvhbzuO3EjuyKz0O0ESVLLX/UZG8hxHJ14QE+gAZllmEonRaSeV
BoVbvMv9ZSzEQnzt10EdzgeTw55CmR/qfXkm/v0YMHSnDKc3KeNqZsAUoRyQdv+p
YR/3AiJEXwi4sNYzKMnCl2PcIWHMuImsDkeoCQqVMjyZ7sxL3KsY3YgTidOReKAu
0ZpVJsfhhOJoiw67sI2K2+u3lE1InVGLn+eVF9W68JLHEbu6WLnZMWQfsNxSDDm+
fnYWdzl5e+8XWp89nOCvviAr8HszRUZUGAKGF8fNmUslqj5/v+Drj+cxFTHeRQxD
f7X9GB2K8xTqP5YrNhYQFQIjASx+xkITsV3RFv5dxnRV3BRN2im9J8Qvxt3EdsRR
g2as+q1QbsXxNcWRKuAUwuX9/T2oKfzKNoPY1wQZ8miyjn0ulilA3BGRV5vQz2Gr
0stJTU5bUd3OPxseFhwvIx5IDBw7YG+EHVBaNTpAwRbFHaYQ+8At88DlD0oqlEKI
NW8wmnfRvBO+6PaGV9Xa+EnJyxEG9Nb+QCWFy/R+pVL+oZKnDIaZf2+bX+l+IzbY
/m6znAb8xlfszyrlYeSCTT5ABCu2HlreV4lju5vr6xNCeituGOMAWSzQYThBtOgY
vnepmPriZAHNMh0Qd5Aw75CGoPKDOJTEk/s9wCmqsr9pjD04SNFXYIeUT2U0x5MT
A7QmHBEoygmGFTGLmcHlGm3IsMUa53LDpma/4oCXpJGS01F744fGktsWC06m6c0q
zIpV3PF5E67yRfJ+PTrH+w/J1tnGTW8IEg1r1TKMcZB1HCMpyr76I7kXU/yJoVoT
eBOJ6ws9n6UxP9mtGrlTZK///r2aw15h64bizYyb4UXlbk+tAGsqMuQiJsTzCSwN
1EvcZU3N7QWN7vJy2EUzCYSF2AqK4DATfN7go1BeOGy/wqX3K7aXuf8yA94L8VlE
gWxW7ofWW4O0w4jciUDCaEHOcTPvrKVlLoR+ah/3R/B2NFMFvcGlEGOmDK0BEQ52
8tfl0CtrsRKq5h8CKiX2ywY94FC6zTXlnq4+AJmQbFwtfRkc24XfAOWYuQESYNdp
xel7kYfvMNmJpPVcqkkMSTYdffcWL7AI4b0QtNcSUcLPhBMB0wNL9nYfLedgSU59
nvNcSFnvKASbl8f48PEk8c22JXy+rFYg4JZHR/4OFCGAyARQoQsXbDMQg9IdQ7Ft
h6tB2A5Bv5ht7IEXmPHxpW405r1vjhBPt3uwnHG15OUW05iVSSK2GZzvtDPX3TM9
QhaEMeqwwGUkUlEyrpdvLP5MW3KPzztrFkaLszWWSeex4ul9nz7YeFoujnyOECnO
4FqEfd7bH2UR+2IxZrTAFGhksrXtTCpz4pOoXpFA8kseOrnb9syYpB+QwWXay3zi
UmNbZKuNYUpoveQpzkYxK8m9f+LBKD550acu8x9frLBNEyFWNo4rVgNyvVAkBtl8
i+VD03eUXMAyQbisTUcSzP32Nc6gGgTaVDycw8Djm5mGD48bYMeaYqB0lvzmZTEb
1B4N4Ozcqv44yIs1E+EyFSSlS0ZDjxyxWcq8e4idcwbYm34Lbu0HBguTtEaaxtNG
suL3IMjzdWtYgyjBMoDEz0U6t16TM31RXIzP7Ylg+3EW+tctt2iWIwXQ2kNkTR1B
kGCKzblPWo3HsK5wW60/0gwjmGvIEKPANJvjsS+qJWyDxoNZ/fxEhSVK9glXgLEP
Hu25TwdQNigSgZMSX8K6w+aqsuwCaLknNdr97hQ87gNFy7ldzRxp5kZtwNIuw9JF
C+TF/aozlrZFiyZg5sXH8ByTrXYB8N8rL+QvEBCHCpNB8LaC4UiyLSQShW7DNogZ
N/Rq2YBlIlfu7YDbcqQkgXMD36BQwsJFfJO5FsCtZuJecjvWrYfPZmlWmhSdjGLO
IaJRZlI/O0BMFvUJN7OBBZ/NMd1oTQNPy01fzYPe+qIIe6C6NY0NGPam1Ng3v78O
eDve1XLfA0Y/fXDnIk+AAmN8wrT5FsHVVSMxX1XXKyPls9ti5ByBV5OywVa3kT7K
enc8yWoPN6o0xHwXW2bkX/3jIhVwQQfA2UPAw2FHG9we1CTgSEIniOstvOR8otjN
nsFLuSSpDsQNFKZJLATbwQ4n5d3IzuMmMOrUvLq4Jbws/q0lODQKBssyn48guf/Y
xgT/yfd80gwCWED46oVdBrTu24TZBcEFcrgMGOMnciGFby6f1VKbF+sMfgQoX6zp
eSp8wSfpgEKVPrWmKA1+APm5DM4HUzxCTfc2CunyT1esV6SAru9BJPWakd65X42K
Ywxd4Yc6nX7PAFNurbIiajvnsGvu9I4EkxnpzPTgAd63k+jsMa2j3nhDelyvlHAm
xx+6CGM1nDCI54CllHQxzFHJVdFcFbq18jKv3i06CZjHciUVSwEczst/GbLOKXJa
Mmpx3cSqMTyHVW8VQb6rO2jqtiF7QIDtKkI/bBb0zoae8iZtd/vf+lQ8nl/xGLXl
qT/egHUXg5RIGK1k1NQrlO7DtZs1Y1fEPqWFyo4L1OCCAgF/Sl+qk3fEUPvW3SFg
mnEcNdD+itTzmA3rMCoxD4N6GwPyv63QNj5QkGO5IOBQgq4hUAG8pAvF5eTZ0n8g
s7BWRbbUCX6nkmi17hRQW59esnXZenzAAYLb6f4NOmz9tg4Cpq0TuvagaGZg0SPu
GhOeRpvqvT7IE/gTFo0ruLU5z1vY2haMWZDlhYY0xrRmuxhgmXwsJ7xPx5Fg/Ktq
2VRsIj6CF+jogeVzt7gqAfmBQsNrK1QFdLIjYL/7IVzj8C6QL3VYx3W5BP226rmD
6byEG65/IxWZ0umrTr4QshAUUygsNWyOU0sSN07oIjJ8FkkbEie6Bf/0E1y3biVU
XK7uDFpTC2mBuht9fQmggW2/xS2sjA+qzV7DZyaFFF9D5gTeFp94QCVuIySmHpmS
xncg3ItnWGRHYm3sXY+vqVsz9pu7q3DfOdQi/2Zun5s3FMjt4cAGOsC8ems5ueUZ
/zET/hqbbYfBN/aqjeZ7jdBiIUj/czpXdhO2rMr/Lpnix2D4rdErbsYh+SCfVpHe
gOifhw4bz+2ef7E5qGflrjOo3iKjizFow6mx+ITMcEHIZXLTZNdvSuC7mdUhvh2l
QmtjFtbmAdx8Sk5Rp41A4qdfSna1yh7FTxZuFokSPQ9QgLmgTNtCKgLqEmMM/fpp
znsygdTnMZEi+lPZfSNxjY/28tRxpgKvvSNp3cTwelgznW9YVdi7y8Q4jh+xiB4K
CJ8rIoi/x1sWhYJYk3dcnNAcXiCM47OiXfDoMmu1YbAzzhccQfPm2mqfslzpbKmA
bGmob3MHzdaYCX/XUIVPDhMrw45SdMXIc65MH1mF8HgeY9MTQnlXaZsW4r2m5o+H
oBbTS4ipr9hjs0UuZP9IMucKUATDzg9zPOSQXkXBcW3GuFx38JmkEigp30c845AC
Tqlv13rbwVn/6g+mYCCMO1dqkC08gSP+2aKeR88cEzFiFZ5i5XKC5MgAfZQbVj00
DPuxGbB0nxm/4ERy0nD8BNsjoMgWe234AxsdMfq9NH1EhcWKeze8E/++kMrdSk3i
XE+23mSemgcRwHGOAlDgf4/J6gi8wRB/zJa0xS1dtpw0flQq+D2VyoZCj8EwrruE
X/DfDmAeXOQX2aDUG4a6QnGmT9MbKuxMHo72dgfjlPlillhE/c1njaxDx8EXlhUo
Pw2IAmhDe7KZ87jdjoA21QhzDJ2QUVBy6ofItZjKSpRqpfhQRpJAH/pJ7tFDGWqu
tJlla8b42HbkZxBO6TmWo8X7YgHyPlUC5JzJDOUzD4P7+TQDep6v0GOFHdYEDWLM
j2jnQLMC0NdkYKHD+G/Tik5QLgs8F+0E0jerKggHE8+mrbKWGOxo+1c3UWchKCPT
sIGKKnGV70Od0CZNz3h4fkiLE41pB3U8mapRW0RFyvMej915rZ+wf1DOL4fo6W1f
6T/2Lg/xfJxehQidjP8hrEZP/Nyey1cV49dS1ov2fjZ4xY2EtMT1VAyt/ABBgrM0
PGZIgtVt03naC0j33FuNML5yA40sMUsHiQ/iLYdmFdP3/1oUavbRb15JmRmzMEme
7Jp+bpNHiPK7xzC20RoIqcQVfmFRAEZOJWIi+CwVuA2XkeUsuV3dLSU07GWyuxZy
m+WEopPFuUX1UZZDZOF/3wWecjB6ZQcsDeKFoYjxSvfSrI/OusVayzUAEfaOoWOB
JN12Gfzxm1QhdPx3ZL6AK7QB44eVrLUW09osEcqAOGEAChRKKSiY310R3nAu3/Bd
2ZxqIjqkB4TXp1IQKxmsvKO192v3keSeAPRvDKh3eAi4WYDQUZE3j3/S2gzLPIML
nk+B2h6OYoQYsAhONsxblXG/Flqy3+yoSZIEagLUzJOjnf5367efIPPb5B1nQpoS
jibkFby09SCYEnHpIVNOmLA/pqtuWV2fJV1vzef3xLMTX+pi9TbSunUfhg9xy3jG
Jk23ehwRKnRpcIwjc7GqbfBIRftfxA1ZBbLDoyURqVOF+6DOjVsNetjnS4EK/i0O
8N6d2ZkuF85CoWQCS3WOvcPhEN2V2epvVQsBjYPuqhv+QVSwn9iADJ8W+2MtHv07
CRtDYYJ58isIFS7y5fnsRNtYcFZSijuEXVvrWhb29diClLvIXt8E+77DrRmv1+Wm
JbN1wdiPX0U+guCixGwAMrljNB/Cmwy2zK+28qtObzg8QLJGoeVWyW4cXyOP9Qjw
fUCOhsxOrNupMJN+orSb41d9cfRo5B+0W/jOjjThr1aCzGN/du7JjVA7DrHlvdwW
IhX2qYXT2/agRclMXiRErhREK/g5jqvBObbtfqBoyNzCZO5RAIn2g0p7DYFzdSIV
vTx54O66QXHRdv/A3/aSx3FLp0xAZn5PoIjVFzPhF1GCCVdGcBbUCF6IKOCkmvpw
d3qKBD47gRkHlUuPE2uyhNL6MJXaH8bRaRvjM5UVrBig/JQLbN4XCJgscA6XGicO
jXAMc6Vs6Aw1jYDcTXnOIPV1IzGG5DQ6ZvfKntnV0RFYDqobzLIRPxGgk+q+1uNh
BNORLRcvy/WQOUSRkZOUmiLy4rBALVcpbjv8qZPvVgVP+E8fK6mlTI/okHC/O4In
y047v/+Q5jYtCjs8eQjgIu/4EhQUpgkSzP7ko1iZntmZQrGZxZe25VUv9+KVI+JG
g7s2GaEsWgnqUCDgj8hR6nCEb0+hzHWAlthniqmPi8fKc17+ac40WfmrrLS1TZfN
hs6FrN1ckLySXLq7aDwNkhapvEOc1ukqyjDVCLz9SjRf0DLC6fSN1ufpL9rgVk2S
s5aaQ/leCW27jlNMl9KYpY1XRJZBY7KlFK3YPkPMPp0AYLEye90hoJ51XjuQ715t
fT3DrCOZPipou1fGzobXzvWT2NJ3kuIpEJnjiPxugy9cvefrSToMUruTIFHuwzHS
p6KucLKdVXdezWkpg1ygVTanTO3dCu+S9JH96tvYPm76N/SRVlgXKCK8qDMNVoRz
G1q6eh7FohkBAXY8H7VHwHwmsZfRDxD9sln/lSq2IgSAWk4HfZuGU92GuzIVb59C
bAHnYD8kVgAqirj8tbPe45npFYpwc8vRSHoHWhqddOw/ZoYaVnpqUQFvG/bKv5HT
TpycXUHZN16fLVPei0XvDkbvTLNQ+iv/CMOGkzTJmgyn7TdlWQ3EQ3DTVpfVsdzU
+LfDpnwDHfTMWFwKSDPGE+GEtOiZbk+S+k3S/66fMG/PdkSxEO3iwZPsR5ovlNOl
4IsYcPEDHC2OJWncsM8UYIdUb4hkZTbQZPuSSr4P/fdQnPmILWkJkLuZW3q7w9fu
JaDT7F86huOHKk2gVCt8vrsWHSBST1q3BDa+3Rj0p5Uw25gWyFsC4vvXIHQJEECC
kl7k310lLHGo2e/5DqibXBDSKzB83DcH9jhRHfSiNq7ZklrAi+pJyhml1gzRvvZp
j46PPfLhVPVm/CjL8kKxCC5zSdGMP2dpxyto7CjwFLwO34dF3mn/Bg5hQenxxnVg
MAXCeANmRXUU09Z0h3UJUl6+Um05gRr4JiNsafAEJHPhHu77BOWTFLL2C/CD/eUv
bJZMPQlqqaPPnN1Snq74Q5pTg7EJQX8DzMrUtuadf/ItijxsJcvTdIhdwIiKlhtd
R7eCK0SgyXY1thBrg4Ktshr2nWFR3Ow0AfPb+ozt4s9vorxWBfBgB8EesQYlgbqi
A7a7KYCCVYLuaPYwq18as7hiF5AwqrtwPm4n2y09+fWPD7v4ncsPY/3xzrIrgPfS
4kNEJcS260p/IaGiskFNvXPvb/KJFs5IQqtwviXDFZlqmBMklUyc8NNDtxGXQQfu
Pjg5lgk/BnnE6c0KU4EFXL4mMau8ZM3d4m2HBLBClwMSXzNT6bUz3HWz5VWQtbji
C4bAyXiekA5gp9l9+GBfTgwTNRws9Kmspid5agjvK7uyUIsv5RHdBl/+FCa7fS2H
de1TltsrDIa0x5mRN9iWBVlLlqTe9GI6cM66P63w8XJeWcnZMRhgBqyVSVLW8KBV
3x+B1dkdR7MxB0Ly1eywV0IfIJZVrzS8AO2Fo5u73qr0jdWKKoYdY//goxcKMmaH
OH4a9rYFtiXvLQ9goNCCc4sIXZSgZ59/QQs4GUk3y0nZBEqLOoYBmhwLcr9TtTJm
B678fBySip3nZrd7bAaygvzLk84JanTQ1YW1FeFO+2hRC9rYyPT/2/yDyYpycI2o
RF8t5NAHZ8o3VPrzKGsU2Zs6u6NU2EqaIi+KtpIiGIRdSKuiaYeeFkHHA+QccpeM
g3QbBb1kdU0FM/L6q+nh9bBjJgNaeAw5gICETUN364X8YXQtD/D3P/rBXJ+G7Ehg
A/8WgbKSggaHY0zhIG12AyIFjU2t4Mt4o9wL1rBRqV8uYVRTA8ax02M1F97t4kf7
8cD+XQdVUc4GVuX63t2my+wuzGdiZOTknS4U8yWHd8YD1TtJ9g545J8oqteTFgQP
wHCgi6DR9wukY2cuUJ2/4oP7nGtt700DEvl9qJNd/hNTUvyHkOZk655g0+daymBo
xrHeEmRcC/94M0ve8jhUZpgIu6ksSMY5C3HMOfxFIQWEiAMjtEwQ7a8WQ+OIHJPO
yzlYt2SBg6UBdYPnBTINhkX6+vDQwWSVKBcHQUj52Qzu+UYcU6JRRnTQS90AQL+C
2LCFYHKV54KrA8dSukrg0rMZzQXtfAkL0OFRFPqLc0z3O5K0Qq8C+glWJzNkmfFV
E7KdxiGuzx+gYFZdSI++66kgVm4AU46mLHcKh1pgGK9oW4pon5VynIvCoQNlhHQB
32QspUiwYy3alQl6lKSB6gffdftuPHMSM26FdmZsLxA8rUtZUIXz0C6bo6Dk4KOT
ODfjptuzchMflnhhdhNntZj5fCf2dT5+FjFEVu6tsHb8I6i1nO8dgaKnIf3vkfCy
f1l5d3bf4sN1DbMbFIClEfLUkZKYKWnyjNNViZYjzLyhsSJBxf9o4WWSvLyRo66z
ZjxVHoPgzljKFShkYlni9NN6KsHOKSOwYJXe95LxlpBC7fmKbrfUDFpQ47IbdC7T
Gk0uHaGGs5tynMbS2H39c4vULxlOdU6pqemCxmbeUOPkvrG+tw8gZwxe0kr71+RZ
PUQQYFyIkRDNuh0hoK7gee2lBg5J+TpV0nWITucBkmQx6YdNwsPjTvTzHWj2tPj7
kLGoyzZogI8OcbqYczEL9gQ68knUrYhXC6T4AZxQW4W4ophBOOIX4V2kmJkDSutr
tcMrh7X9VjDW8qr61nqMRmS1gbAU4DEeWPjsoI203aYNKvD6P78PeCgmNNNXxZRi
vIroqf1PpIdwfXqp1F4reMWNL31kp/n54fZndyKIx2hcNdSA38TyZJ24cMjxT1L7
zdPNUYvW1W6Aaue03yvHhzbSd0vTsL88p7UASSFebJDujqDruu2v6txsIzpwC/ZM
QyqRRooo1vmMzTLeycmuq5fbBH1N9BHjiq2Ses6Xk9gNnubfm21cTs2hcDc8VeG4
Fq2OOBCCzEyC0YjR/Wvx7gYN9HYGen1CNCQl+dWclEfzhzbQzBw++TCagfUa3/Ll
n74XRYT4NO+2fhfkvdBd36t2uRn5WJL7tEN7mHRZKBjUij6YjfOXgB5Xhp3Uzqr9
WujKPhWJbSJxpniqjz5w9RB/kN5DVGG/jXNU8TEIUFyVGKhHe7eqbemgxxA74fgJ
K6u/D2zQfGi/Vn6cR2eQnc771LfGJ2vXUZ4VHcE3G+tG6G+kfytI3GAKdg53rM1/
H+hZqx1d/gZGtiLyiCPzIh6aoFLAbDrw52hWh7ESn1utoB+mLkp8Sc7S6kzF8dVr
awPgLE26MdTvmplSbeNjZ4BGDOrZJCYfe8DLdEHOrCXbQxDBnIWs4Gw5XfXla75b
uZYK+L+Q3Ud9YsTsg+wNuWvKpYEZhohHRhf5s++tjv8M5f5NzvYK/nFQByQ7E4Am
y3p/3MaqIdFdMThFQcQJVypCkng+OhteTAXA3VdaC02hOxQvx0tC7o40Rx7rI1YN
Q2aKTte0AADn2h2uTsyEPMt5LrwekQdU6dgYZO+5h+sghJJRtSRAhS10tzSXQDrd
iO4NFdH2pEOlpw3A/ZAdGRmBwo+YG5HzkQVsphoHjaVi/RQSpq4+TFYspYyBrNfW
FucE9gHP38j11X4oV6Qj+Hi0NYXUL2seX04MMEfnQvwZGm8gd/TxfR4kPMBOi6iC
5XpleJKxejs6wxBcwqJnhnx9cWf/uAhvOgqCraW2vczZ4r5mwX2UUVO10aCDNOt8
l+tqcWxHHLdatewpzifZiLAANH7mi62/ik9jD9eg8zSzVNpxBI0iIZHQJDTsEOmH
o/gbM1lpVjfUeZB+kwvCj4QiQ5saGgMg2OcxiA9e438XDE/YdTtx+kPMgPudr+Pg
HoOL1AWOF9CTB/mThETov5XEC/Iizder8CqIN2p0A8KGtasC1Kt5ungh24/7n+nI
5H4di/uD0JZRs2i+us41472+7YX5CiYBOj8Op2cP8v0iBSaDEufs0WtaZIs0ABPI
Wg3rtb0nydY9AVElheQnaAoU0HQ+APp9SlADGuoQjtqGDSTIpfMRmQn46kHD99c6
YQ1ascIyBtIIdL/Kh8JmYBvoEbNc+q/GzNevxItLThQcDVF5OcNhOS3pxZlWsXgQ
lnCf90yhPrKqmiHwE5GDkvG++pnRI1XUexcq0T+c3jpf1QR+bP70C2/UZSXkKI8l
FjpuMD2Vhqi54USKz8lqDICuhE2OOOcT4lnABXLJsdibBP66aJMugKf7Nf/aGv+x
Uo14EaNWnKEdWYs6A7nkZ0wpBT42nhTSo8sq9gw3+7/LRnGrTuBwhvE2nIlj3wvo
WDcnNxCSwBCw7KlxmIjoL+4Z58WUH8HD7Ti4GR/LUGjwiEtZuW8SdLXxXbPqmhPR
CCppm4/gB2vLrmKyLH1ysheLGg8Pnu8NY9ai/WMPpjnWWef2Uko8QZIZZMeAaDOE
yTfPUAp/d4AhRXS3GuhzD6hTTSI2SnbLwLkwgywqB2zZl77eGsmG5ipKWx782mVP
9KgbXvLw8h/lmFefzDdKEpQdysNX8kJ9sHGIG42uXT1UULnqY/SrK+UiutzstJlf
slRsA6goV5JaqdnXHjXi75jvakWCNnAF61IWmtSHAdtvuhIMnDd+hTh00ZrP0+J1
kF7RhxQUhZaZJ3KmQEXk4F4HmAeMrutGq/sQAaZ59aK2M1leSslDIVGRAkuSOKw+
bLt9O2YlwIOFk86LvAwVRc6KaNrxRLZ7XmJNj7t4Yw8IqX1jyPFvnojWM/sUxYMj
f12r/L8gNAzt+TQ7B2s2OZrj7rT6gkEuVfCTEvE+DsdBaLQnVjyzt32D2QsK5avs
qlvG/qUD3D8y2K9QMAr47rh6FTkmV1PdGYH5SV0azx31qpxIydq5sIDXKGvaDK5f
fSvJukwKpR73I6Xc4Z3sWvwoHt0RJN18KLOdzpZxR8u5CujD4ebE6ttCgl9p/sVF
tsAmRiheZGynC8vozrkD71rwpG6ClLWtWknIAS99I5wEuDEOcBU799RJP/NwulYd
xlw5L1xiiy3Mgh/b/5NXX4Bm8PtHFS1mo/blDSYlfh2wWIZhZ51xa9vfpQkvK0BE
AtUdfwMnUgvZKa8slRVX6ZWDYF9tW8OVTZXxnmBO5iufd19Saq0AGZZC2EMAfr5p
xGn51Y6s5oAclC7y3lALIKXHaFHOa7dHcF/A7qoKHwJw2q//GKT2Nzs3VTu7oA6W
Dm+2WwpaGKEg0oKV2mvEHisjwhHpsvwGTlqkfOXE08KKx/8jH5a2bCKvmPjWVnAS
SN3CfnePiK5vcaHq/DCF7nj1DmqKydrE7TB2oMp37Hd+qLchrzU9y+W2Xr3+OT7z
JE8KIwC7K5ASXyVJZlZxriEIKLophH/eOfeUzsJe/pjlSoJE6Y1C4EFcCNkTNU0u
7chsnknNTJZY1DjqRsFOkjL8fgcGcNX7whJUXKeyQPFBuqKvOWOwd26WEcl6wVv+
LWtRpPtB0FyFMw7WjeJ7Kf+2hcB7npWjZKhSy50YROC6aTktoZllg3LFl/6nOGsu
6RYlX498AJWuRdW6CAojz/T1SZgfktEyh0Sj2Yc8KyjZ3NrfoiDkoFsjKgcCLtFw
5eIlhvG0aMvuKnAqcOQEXUB9isFr+3dQ683vDEDBod2zvbd5CdPKrk7L2BjE8+FH
2BNN9TuB+sOYxuLpJux0nKc0YiZqVmPAESAXm82RoG5U+tznZIgbnKZiLrDyqbov
4lNmWn9VZZR6fWgUmxjz9bwI9JL8ycdYgomN2aMAHhrRLdP71QCM0d0yV0nGEJKS
43JhYIdYRHhzqHY/w1B+6+wziaKL35RxtvrFRLD4zJhHV8WdOgN1+RVlkfF0GMXr
ng8IaI/uBicacmRaOosx1VtmfWYsIySpZ3UeGW82XVnqyvLyvg28Np9a+CPdyLLq
x4ygvi3Bh/X0t2/gkrpq13btO7TGZQ9zkdoCh7S0Oga7otbC3anaBy8b5QlxJSJ3
/tE7YbfEgujYnb42hgCVVghlK2raHQESECXG5bJlA+1JnwvvPxnih8TBKqBNgKEE
HheOASeLmGI4RfRNWjg1sjk+AHcM7Dz34bZmXPB/ZVSjXPxlrTcbE4Q1KIbKp6W+
kbCoCurqvvvR0QLJBkBnjY1T+xmbEs3gI7W/MucMAUnM6dDRIYVk1Vg4GjjrrMvg
xBlQlC79ARx7wxMEfYsIeCP87DTmshU6YXEqwotoCGVe7s1sKk4Da9yIHjCqE3Ro
xlMV21gGCqzSuFmzYSlbswRlAVJb8W17q5ExNm8a6I0uouhP7b9EMvWWW5vgZQIr
rhPRqTl7QK5ru58+1BkN3g/qFcxZpln7he6uKr6dOhMJcqaLCvwR1AxaGLOq662c
U8ymizF1xeTMw+aAajBhsK9v6Jq545XqY6lxxRKpFuunwdi4246ynihumppQ/PzO
8bcab603lZ2jv2maQGlvZ5Ln00UkIwu+9b5zKTZVm/fyDxsfNFUpV3hWXS/O7hHC
lMr8Tp4tDwrTWnSPLO+TjolZZ8R0CkQMXDIqLoOnZMI6zssFsV31GyOFn3mRhwyY
r8ufXX8AUrjK4sdniv3xDZVpkq42Vo3k4A+U0wOvWn/1lpcq++mtusPwG31hsSqc
X+UhxHQDW/8HealwX4g7iDRy/FRpSgXS0Kc+SZC6hg/0fglY67B4wKC4gl06frAK
9efvpuz2yjd2/YIF4aPnfvb/gHH+8Urm8F2Jq9fdexL61K3JynVlKbQ3rwAkAYiP
H+BZOY1j9qmpeSfoDHkD5Tiz++7lgp8DHeKWMB4So7lDk7rF3+pCvJ/Zr/AqB33K
YXb5jnxtvi/VNcusq7b6b6NIqyt0qcV80zgbAtOqVdAr4sXcbknyn1yT1eIm+sGD
RHx09jTnc87tHc8JVTU2La+cmhtAFyb+hBuw/HwIJoLc0/7oAo7pFNjYzmcN6/ZQ
aUZa38rI9oyhwS0yOoZRfNnfZo+RUODgFqxMLdONAxZ6jEurR8gqNgkciT7LbY12
+/Ml26In7gsRdrAWMuT4xCsUOcAMROIjBrKhj/X7+9ghp/qj6GTAh0KngSleYEa7
gFim0f6G+S4NLoSUtU8xQbvnjFco9vaEDNeH0EqgBOBV8mwTZ8htN7oNgmh7xgkz
7ZqvLTEzrAD8KqWHdpnshVwAT7OiFmXL2vz7k/10CmP9Er9D8ZGA2VA0hmtwonYX
5/Fz8jbGdo5LwtnlZNwvXWKwOIU43Lc9cFp2QzeqT6u+IOASk8sSnsR84GLnxxPQ
pXETPBCfi4o++IXTZifU9YtUCABm1kQw2HLUP0ywNn7/GfxrZgqjEwc9fEJgD/dG
jKCHzMZ6K9dYChQwRATOp4G9LovWCE90Ev7BsYojWO3XHTowN0QA806Howxh0bVc
Fxb7k2XPzm2cIM5MTFRor/9X9sLJvwta/WFYymv68nt9+/Hjhzq3zrso+OpOrJcR
/fSg2iNpuaSfDwQxVCleOpighLaR5mrJqNhrvJC1NxXVZx+oNEMipetqWhYD4dpk
ZrFIRBXrMzAmVW6HdM491cz8FCOv/vLLhlZZNQuxbE6Zdg/6BEIHOWxA2F92v9n9
OvFWNqMfjv828s3/znVdSICgw9tHWJV/Kuxjl9PT2W70kBaCkEgiuOGEE166edrS
1ZNBeW3dzl4S1KhduQH2bhYHB0SN6zSqa6KmUks+smpbhC5fPT8DXgClftZd/Wph
pbJimDCpbnBAYRtVM9dcwRhSTluCl4TJSfUbynCzxXkVdRAfDqzPhaJTgaAyiBHR
ZxvBjak8YRCutfsKE3ygKjhTEp2iQbI3TfK/9DtiFaJNThFtx/UwEACphQu7p/Hq
VgxfdA6UFTu+C43LKQkBDYxYfL8nfNo06aqyutIKheYvLkbqtTYKITScHgit5heu
YmpoPlSON3vxLxTUkhlapJn0eyYW+RQ0hPUXUYdU5escViCj5ZgW0pJuujskTvpg
GYpx0gdH9uI0kbSPhQKRwmn21X0Pf2PgUUUEvPjJuNaPGQXLe6UL5CRO4u2Hi4CD
5R6Xipr7yTVmFGfms2dBPOvnC9CLZTfiQOButbfABWjOcW46uW9v4aB1RweJx97Y
DhG+t/GHbihHLzc7SxV6+thdS13Ta5RgAMcodHti58V62cxTqBk/H54gWpOukZjX
r36RHw9z9mQBUPTz4hhvDeEkpjVCeYZZV1YPND97Y4NHlJlbKmqdB1K7Eww2FdiH
6p+fAV9aJBEJkBKqKmdZeYK+X4E7lE85Te9x1p5CxqmG2nW9s80IRiiUHi3E3QwD
Kp/u/x4CQYYXghDXZyNGXgedT7tvk/x8OMBjNaeaggGbnPe5ApPmqWiNn3uK6Bok
HbnOgAayRbOpoi8RTt+bcb2Xjt7SqbWTeAa54ypJqm+tGZJTFAL56315xpYNTcIg
UN/TO+wxTTodpHLs9WxHLmTn2oyhn9xGJnc9uyUK18NHl+7WiVwkEHsR2WAjf1JD
eJJGfuD5p8U+DqvXC9baq1b420nru5usALboOYn736afuv1Y9jebDe5kL6uxOhvP
j/jXkLV2f79+gVKBEDCtFUgLMqRUEmMZr8O5NumAUIwSUI5JKa/Bhwvx5X2HYNOQ
Qio8GYuBTllMM8REISyympHtQTRf2zEnJ0UBJLff1TVNCqXM0aXJfEum2eDW+Puj
TQ80tk6vWzUL+5X/xAZKvxUlODKx3bcKfgohi8EcIcBSQ68FqwjTcwl1frx3ckKG
9hgImQBCepAzCyPpUSQKhg+m+CL62+82w3vZlSGkZcAmcBEPgxxc7GSpteofQRXJ
sH9UcJqnpHa83pInkGQ13ZouliDNk1Krsz1GRFqn/jL0z4syTVgRRX3HR5a1n30c
+MEHKuWrfsccm8beRG9voq5txMMOyCoWAV6PIG69Li6ZG2SICaZW+0moL34yfNzF
goBBtfCzvVPbM2+hmlcAYs2eWKL5BrgafFH2U4C0q9Unb8vs9Y3i7l2iGzrlR3g5
O9NuizVKj4etnvAlqk9vcTH93oqWOLWfcKeGkG3C5IQawRZcL0kjdEtlmhPxwnFW
G/+18tkTPmoNmps0X40y9ZAyL/39iaccFEKdy+/O+bAQ9Jh9iFKyUJsNGkVb2xC4
jvLU8aQtXCxaPGmx7axpdM4kdvMQULZsawrbbF3vl0rnrk/OGQBy/yiuBybO/Qvk
cPkJvQZgxNPVd2nhUE3CHDkFR/xFZdfN1W1QfYc0af9sR3IQDFb7JmDsO7kt00y+
IuAbRfrkQwyY1gcEM+Xy0uabPwOEfKhA5Vne/VcYd22dIQs16RLlCBqf4ION+uqV
qKMMorBAHBPidLYH9gi6swSrMEfwxdVHGXEnn4TjUdvmyvWUrxht/AfLbfWZdXAE
0rt/BCIxg0Qe+D+ftIcBrX52u6u2ez/zdIIGrAWiqPOjvthIXAsu82Lfe3kGJtmN
pqr0lUrTYwITLseBZv70MME/zAp1MpkSdwkqHtOK88WzwjN2IB+V/FxRv2ladz2j
AHls0E6rjfvN0f1LXUKkReYxcGw5Vvqld27w8i5+ZGnaECfrjCW8H/sTl7zQ1jTf
P6KuJTPEupVIj3CAZi2TNt4/OO1e5Nh7fBen5ZiKu4gwEeL2hq1RqSlFbHtoDoSP
VzZqBYu1UCVoXCI4y6lcKNKBux2zTCU/wh7Ms/MeKEoRXp8BaxRF/MQ4Hfq8Zvtq
1JxO4g46kPVDew3L+5+/qN/N1WLBFm5xLqxkrV7Ec5U3/53l3niXw2UF+VlWUUuI
RS6+WUFJ9YHr5SW5xZKpqqd8N8yVwyQo9LchmHoAcGRBlB4A4xf1uBQW6/VsBy6t
zYU2kd1yX7cQwK+ZdvbTjp/yYZdrPDRwosGpObdhlwOdSWhFus6N8rffPulHDqb8
lehZGQyqz7u35pbwU8xYhH+SkZOraVgo4z0ov8RAq5r8CrDrL4k6U8/dYOyuYs4s
960z682//izdpcMceKUATIM9BUel0HiZ2PEC2YYiVSijEn/1RGg0tiuCqhMMEEIR
EsTeC7AUTQZV3JRbK7+OsnDde2ifolA+iv92rSJ1iN/3NwGO2YA79GMApLXwCfqq
Aoaw+pIqjuL2dyOOhKHU/cznb4RMcgQr7yxAqY9z6XCUpH0Ty6ZhJqZ4Pg7wv5ld
hzYNeBWTYr7KMvg/Zj8rOXo5cJ29HEr28mB8xx2AnCmQv8itcoek9eGCcjRaK7wG
NJ8FECx7snRGo9n6shsbJykiT0u5jPlXBZRmSA4iEBGGD+gNByO/wCfIb6c0Ed/p
JPbaZr8tcZI2CKz6StLnKMvkAv/bJO4EmPPszN7UkpEHjgCqvHwbmxvSJz+RJcuN
rjFMYsP9/N9leGIgbDw1yh9ow7Z/UPOB1HUsuCDbcP3UW06J5bXDIf0QxQ2PgCJ+
Kic7eQFLI3jd2B0fxLoJ+KDgd3GEcUM2lkvBezZhdTxSoNRQBBRtW0xHM9vXgF1i
84VmiBvBlqCtS0FbLVZoTqbhXAgKv5OZe/lSo495mHMvojvNM89zDwF0VaE9Jc4y
1cNgABVetw/31uu07h9zJyxItKIASXwEeDZYo4Dz7wiQUGhCW0WxTVYC+y/tM+90
iKp72BjJlO7ubEsaHMFrNHITChb1U9WrfqZb6ZMNPYOCV5l6OFvN0J+LLQR2Mifn
Nkk8yKBJtXLhOBWYOCRmgLrxjauUlbSVbUQ7eAMM5TaKngaYQzr+zPuKYDq3MXM4
t0LUT15xkbzQi5J9hwmnaufnI+SUY+cHwWvAPei2qJ2xFREvk+5uyUPM9bwgiXZS
JJC2e9yU57XXv/cLnNf0FuyrjVOwbvKaU2lYXyVcQbWzTym/sd8VftIAp/V66aXd
x2z/U9eE994Ob8P0esWF+cREmID4NdneqV0A8BrvK6/iY7F6kD8KjFXtMkzpw4GG
ulaKQ1gLppr/QYX8lmjoBEryPAJ1F9Kv8piGcNX5YcoHcvZzmUxa5J7KNPt2BzNE
xq5DInyOz3Wakx+cfMTQUSMBYWhtyn/VW+MvWwfr46OZ917+ywy1COgUTvzzXF0N
MQdlNZE4j/dTGmCSOhP9YbXvgr6eb4qKpbOGGDh1Nw3IlMPex+RkoBGGS8pVji+G
BiEI7GswS755IPETELnNPDkWb3l0z8U2Cvp7KMhqaPtt0iTKD4q6VzWv5mwyGWnT
9qTz1SMMVrhtgPcqRw5pxkwXqJ76AgkIlWEnIqTIFi3xnLjMYGqnWSpHB19DCX+V
4ZgeibyRninkCAHfnSOuXnlDf1FVMMH8C0ZzildCQc/T0yd8qmbG5XSCR0JcdF0/
lRHhubD9xJgBOy1N6HcWQrsrBV7AgBogp+yktC+0Vnb0q8YfCJd6qG973ZKr76/j
UWd3W47GQq64epGRYjdtHfLjPF/wcnhExv+Wv17ROVwBZshlte79uv6GX+tIocYA
evC3EANfmiqyclEdn/xUAjfvHLGB5ZkQncjfr5KPxdbjmjjK1KmuZyOUE9MLzB2Y
Qk86MD8L6qNekZp9tE79lCAxBLIg3pkZcBTTEbqb/BYLCk3QJeGoQ33eEDrrW/11
2OunaPsD9ljCHDvqygSxUJlQYjlqpjYiP996/R30Y83W35d71VaYT/KTCrEhD0v2
5OaPD7LYliLKpwmvT1P3RCGD41GJkYAtyDPi1mxNEdzLZXnMo947gAKsrm6/SOLY
MAqOqMc0M3lLo1LghKev2CKYVgW4AoLLPnWkWW00GrJ/UnJPNIezI/xOZJztaL09
LdMFnKiQ8piaQ7GJFMJkz9KbraFZFGuKbcqu4sarcwUjQnXNP6r80cx6ye76fOmg
2GoNbag8Ld7mxTwZ/CSeTRbIqbaBbQaVxaP0QIUID5wB1bce/3OhUQq6Xl3x1a+N
ohA82qBLH8w9TjKUlJXRDB4KZ39RsZlRVkehQQwr1NRd6EJKSjpL3CiEJNiAwuwD
g97xzQsGx2V2s0BVCKD+mlciLScCVrKunLJxRxdsP3noxpYpv6ci8WNX8rGmloi8
HFUGOZhawTpa/jPjbZ2+i22bccTK7b153wpMb6EhmoNimief3qw8XbieSgivDhfb
79G5i2CNBBsl3uMM9i652fCnhSq7w2QvsDplCADqImvbVcj1tJvyIefXOsGdWU4g
0eW8kRWi+4IvLKNa8Kq53AZ/UTnUhzocaw1hpaE6c1CDIKAGpyZ+3VJgkFHcxz2k
dNxvZqPdvvmyv6FJta2SPs8/SlxcADHfyILby7yCWlsws90fAbyEFAkt0eMD0HE6
3E8sU7GCJgnn+P7h4OF5CDa9HFwTO7sc0/f4tLw0CaW+jZxV8mx5SCgc5vI6+qiK
ehwT0SMWj/jNpCy6CCdZPinYCOXbVcPrmseUqDx9kJKsJfZlx5nghvsqpthBp1sV
bYHx5EVlyiJj+3yCH/cCGu+FNRDfCmz4YjSqiRMEfLn1iUNu3ChlYJx37d66YG/7
h0plnvAMFedUJORQ8bgQWV4IH15BCNbVkuBN4kXVuHxYp4v+/PYWwxAvhZQj1IR/
VqlECznAhaRLgMlHfzkEj7pvn9KnMo6QNJ1OonTUGNfo5phOi9iFVS0wGXDTmssI
KYCoLg2Wvka3HlT2Vy3qe6VQamw7nReseG9UTkfheq0H36uMp3CIUgRB82SE138k
A8qAOYufUutmimr/LbWB4EK3xhK9FFzfTtHDMEwUBrciPf0VVSPFJh8lE1XaZOtc
/nDvakZcf2BhNqzf1T30mytTXrgoa0O5yEVofGeUnba0W9yu3a+MhhJHtFdD2KSf
7Vp/pU1fItkVoh3m4RXk5Bp7WgIjo+Np8cUPMA9RJNPRPBQRLuC74X3yE5T5bsrg
QhqwNJizl1djTsLlGmc3ziw8SWFdMnH5J3ko6PJxYFTAy3bEDJMlTyKQ3F1QT/4i
uJjyGD5V7kbmfO/STzpgaZ5e94ZYsrySAc3WGenxntuK22jALBf0fURWYl7162gv
rR15knjXVMo4QOs0v9q0V1V//w/5psqdl1RmJNN8bOvsJwopfjLnsYNmrgCFl8VC
cgnQeElTsJVGUwlKxBvukTibDzw0/kANp+6QyG7Q47MEmpYmtvuJagSVoiZnk3lv
PuvI0W+MuVF/wcr8UtZYxw+JQO9cImskk/cuvMSZHpoByEFZq5ECuiAY6bvStTpf
rvcR01StjHQU68cUmvO8bZeSA+qYlcSDFlaz2K/TjjDi/7IeLsSHS4ovYeob7QQC
BkAeFCbb2D3ysDJjlhHvHf7uQ75TYTYKkLQeJl0Q1MIFMWxDdsQaKo+pQ1Y/6D8X
RevvirL1/MQsVg7jyrV8jwic5C9d3i7IQEk6E65e9ZNmV7p4Jtro82wnhSe+/aLM
nHFErSQQmP5Z26l5NubC5iVWLIUbx9oG9T/jREewxbnoC7FYBjGPyY1M68JOLOoy
g5KFWJgjojemvri/wGeUdUE1Mn4byTIbxW0g7YEuZGbgTneeYciCYpGA4wqfdHjR
unLaCsjBHLwvwjf9VcBb6wwslLKPdfqxiCGynfau2b5o6HXd7OjWEh/mNyky5fxY
dikkv+568l+6QaL3pXgUQfmCw7sbp0nlQ/UWQGqP787RbFCZt0zixX07EYXMVJI4
QNftzLQEn0RM5o2Vh1E9hb6iXyRZijoKvT8+nLLQQgMQtO+pELunUyaQBvZUDI1J
x2bRHAdW2LE7+Tk5kDOdLr3kLbvr93g3GWz4muh5IXbSaTP7no9S1dWMubxraMDk
SUe//9QRqpRPOJglqpxPicCCq+HCHLSTST+Ht5QvKNQhOTp5SkrA7PfuxLFgXN8R
e2yHHpA1eXLJSBMZaTC7WN9tMaDoniSYDFLm/0Ku8sBu1y2iVA06AlU/W3opbpjx
iLZKKJZRP9g42TNB0WfkbYPd7HrSfepVBSIgtKrRGqxgn7DEZlielHIG1tWHvTor
J9G8ScmM+vwYYW90XUEVPCRvj917WQi2z+xLktyYdn85/Qr2PtRPjLvEvmsWT7/v
qfm5s2a0CNJclwEuyByUFuqmQq/5qj5O4NZNXzXZsbWpA/NCfprV2UFgQO+Qs+Jl
6c/e7hGK/reH6+QZ/7XDQma1aPNeKEZ5Yc/LimkqWUHoT/jn/FyYGonbFVCVpLtY
YeEUhwPwAgoyVEXhQUm6J2TVGXVCJzN/usYbBUcwdDw2Y71NjSHQn9Q9htvjIvf6
wo27KZ7yZjfuoe/cpd6ge5KSqBDCswc4v1s5s9k2IanWVfHS5GkT3PhvLcGb2jkI
e9oIhiU3ZHfCZtITsCk/zuWsJ+Pbp0KKr2a4RQXlHHwMFFppwfkHxpSkcx8z9mRQ
LYWROtPVYvCMJtSgLzrYSMg9MdtIQGSetG7g4KfNgjhr2J+B5kLhKunTPRJ6PpVU
c19i5YWjJSHsacYDAr6PYlnmdP9pdsP7pGnn1VWgefhFlsBBf6RA9hM+Kb34stsk
2svhaxrRV0XOSlkZbaFrxPMn8UdgevSI30SOIrPeVwfQebBJmkCib3GP7GkXoPOz
yNPR5hP3vVrHbfKkmEyvmwd7dUTPZlvr6NBLOGTl/1FPIF8+o0sj7KNeTFmtiiyS
L/MqRzyL0dpW6bY6mki1YOOgAGCrfAYlbjaofVwgl1GhOjgdthW7rc/sMPBD4PT4
FgBqn179gkikStjj3LiNowUfc00oIqZqlgb2KDrV7YKIXlWErGm+XYzvzat/9dRV
P4LqNAx40tuO2x9nBQHx9IytWLM8nwg3mYU5W18FoLhz2lQOl5s7f+AfjJ+XEMeH
3yVb3kXSbZ8qvLatpcKHTqN2hIzRkGFdHTTmcqJwMDWpOkurVEF5ZJXOcr7GK0WX
AIsHYAWRIM863NCRFOrn9+3Pm1M1WL9iyAAnNBWT0rhIGtI6VftFnh1ZjFbY6ZWB
afPiBYxM8TG1ESXUqZeNoboZk+6BMIR955FBp6QGNIGLikGKZMYqsayWwpdNjK2z
xAJM3YzONJFmz+ru0rSCcgtY+X/3GNg6YqiMu1HKZTyyvt6SVKIVsDpiQ38hbcoM
8pK1QAc8RyRAAWemVzShSRJVj7NGau/dBKDGqJgyyOwumUrOdFENLBqK1NBs3426
MyCrLRzv6Zce3k1tMcA1PPG/emVM4ZAj6M73ZcP4eIQSEzy20llMKaRUI8Ah4Vix
P5EsUstndlteG7Uco+fDsYe/VxX5Nfc99sy7N16/7hPuGkLvLhHSG4VH5hV2R/lH
1otjEPQeIxi1vJpclRZ8Qu5prDppOC/IMHPEPCTYV7NTN1OYQJhRXBgMFTZhq+vk
ATe9Pdya7mS1/LqLuOXqwmKj/ExusqpWozIYx7OcUNpdT7baCs/ACM3ReVozyxSy
l3dqHsgqeDAUNeYtbaCTroPL8aTQKAfEIUveGy14kmcM5wWRAuIc+gAJzz2rXlgx
QFIWtesw1eOtHgl5x13yuXIVRlnJFGakXwdoX/h2BcRkYlYQiokxCyA/wzWSS48d
YVBXvOln8x6ys89Xpg4WGDz+kFqY86SoIGjMq3Qu2YcPx0eh73F0CVKUPjhNgS5o
VNeewv/MyY7j6pURN84+KFSa1PC1fmO7+mfRkLMVfvjY46jbx50KfP2y9WMAMPXO
4/cVGmw/KXoWdAlAB+hQP+ByGegoRJFoNGLoWdo5xBJ6XryjIYoMDGSf+BCOYpzq
hMFxUn7sayJx6Bi8pA6AlE853OqvC0qU3xx0ZWvbKGTLg3h6ggbNIf/6e7YinVN+
QLHCrdDFrffBD5YoErm3Xgy/jaWETvsfXIcEaP5IHPnqk4Pl4iwInYtJCLf2C/I8
hV0oZCNc7lyFnAI3xa4CKw6vUXerCPXpPkYPkkUO6KBYnmGqAvWxFc8rG7xnQKz0
8tLb8xDKYlYRpbS2cuXqKHBaegFMaYcCnn4ADW8vfU3g5FqKoUv3/ZT/6Tvu2iBk
lf7852WvOdhdAVUrbNkgckueEkEsLnJwyOc8zJNQ65ouYS9s80jMlLSVK2IbFYPS
gTtVc01yV5Tw/l6M/jvIl0pe0N78v6341FomKCdxBfG1aoGWJKZqvog77NdacSeb
2ITvin0UMA66f9Tf3FoRpOovz54APs+5W4T7AytmwsXNY8qbdfhV7+NWaV69saLn
AJXf2ZgFWoaMYCl/5MGa8VMP0mJFxSgIjyfCrNW05rbM97SGkowGL0w6tSsXXdkw
iOfYKmBJZPpLT8cdlJmLDWeLn/ZcPq23oEql3r5dV6i44v85vaBJocVVnSk31TQQ
7/+Ih6CZzL12uJfrQobtwONeEbyB5LWBx3R6Ci3Xu8uNrPAxMQcmnv4/ckRxEvuP
WYBX5KBxho37V7OB/a5fJWhyVAiyYQJlN3p+fdEO9qDflp3WQmN12IcBicis91wa
l51j2RG7pUpn0y9ESFJYkL8Uk3Yw6os0C77FVJ3UWorD2ICw0bLJE76H9w0uruiZ
Yk2qr1Womt7/C2toW/3t/7HZJn6HJnBPm/2M2Ljyx8XbiOSkQC/NIVORxeUP7+a0
eL94b3LjquiEKhvRGu1HDIuZ9ymAlUQ37nSi/BCkx0stDM8w5y/uoamhwo5f0zM0
6ohibofn8Xnrq6+lLp6UcDGZpeykWhM6XAcTTsDCMJK0LDKcIwVHoLC30N4i8oWh
SYDykBgmgqqRDG7SWIqCNOUkYITO5zBzVwc2Omhkza4yhEkR5HrhzdWnY+nabEu+
GRBYz8/g6mMLzSVya9j0SCmuQX5SWV2B004i9sWCBkhBd5Ank6oWjK4mkyd6eD2r
9g1Ax2mDQ3ma1+f0VZwFksOFW24jDIuZdfKTKWR26rqH/PFEnpXom3fCc2LE4VDf
nYXPqOL5dYj1SCePf0w8onxc9Tw9LhKSq++xSqQadtdKTD5fCV/MHBW6kWWZi6D6
87MbDTwAJu8pvvC7FeAPsLJD+fTgFndguSiBcF8WoTtXNWKh7ze9wH/7g9Ybq7tM
3YSzGeW3KwWGL8hBONplgEHIuyrY5nduzQRx5eGoeQHaCRwTSyjPWdSPeoibrKYw
wwhNby4L2EHXLOscO/2x0Y3mI8BFrefn3uLgeIU/bibKQ9E1EWCi+oAkRWgMObYZ
e4WT0lwwOyE43BBi3tSvWIypJLMuUWBkeMMUol3GrfXzLTsvqX9EYes6TOefIAze
cWgNZ6u6TUwgBy4zVW8UJ/cjJz1yZmc82qpca8jM1sHEiGqlY4DRaClhpg/6gCKI
auYKc3jratMVYGyCDr4fmIE1FeaIGIjqcbR3tR18p5ZLyUiNXbcuRYoRgqYzVdJN
Y4zlUw+Duu74K7gEcMXDNqIw/BKWK/wWAcLhWKDra+7VA2WBPFoWDIPeikTApBxx
au4IA4TR0sLl/aX6hwoAXDRlkRu4v9raEXWREjSMmH9cGKMCnANmRSlfPEBALpAD
JnkoVCc1Dn1Oxc54AP0uyPDbAGIdYX4oqFR2JeojsBImHpwtjSEecwLu5xJPNUqq
NWHUsFN1HO41bMw4KxOiNeOLaomomhrwRHG8XwmKxJrhHBkbROfItKsFUnsEqIF/
rcBUopTEIgI3TwbGRD8zoRwzAAaxGM5+ZLzTqvTiivs5QIVBP9ijzXnMLFgUsB+i
4VPAYsx16cQ+GSVV+75i7QNhzw0Q8Iu72EUIDm09lXbV2HFfTqtmTcucjCc9xdhz
vDzoJ3SXAEaImk/DMGEXR/ZoOdongMycNFYUxS/wLxgbYfq/r3MX6wevwRWYZZ06
KwgY203dRG2ikYaNtufB5MIXETriz7yEP6FIDSsZQisZzEFVmeoBDQARn4MKXs2e
3R260aHFM+4MtUidyD8TCb+NzTjzTdnmrGQaVByjtoU1eB22ChcBO1uHW1GqjNWT
k6sUR4d1RRlfb306ID9cxhSQip738wqJb3wuSvxpNYwSRslwZf6g5inMzCFuVTA8
CfKyqW14/poam+rGju/PRvc69elo/QTpRvheQeh9FGBa7QBHQFipb1e0E3KyvMKZ
fL1XxHkBQCyJxUYJfLsUrD59WYPDo1nTwqHh2wo2N2C3A9QkwSjMNhH15gpdplgw
iaTKkQFAPpizQ5Sutrtta9Gqx0umVWcIJ8eN0Z91X9+4ylakc3Gl7Xqjl1o8hSY/
aaCA69Mzt/FYdri31IMmlWLn9vbWH/d1YpIxaMe+rW5w14cnwevH0T5MTLSttgsC
CuzeihCS2UPbUcnnP407u8sMtiTi4eznfrYKvSQfeuMNLN4djqY3TwLUbejP50qH
v0+dOjgYzZNn+0iMr8rwxdIUxRiMXleVq/cIsHpt65VPycokVRr8WwqXRpdYkj2V
oFdWfyXd9fSgXTntNhIl1j8bGyjcE0HxhJjXNhfT1MkG2IC/ao4p9Da4SGUXnNfv
I4ccqE2Pwzngl7veP7xecDMRRC/7M+pbNAJ3lDEuBnZLz0kiVIr1fIT65gGqkYtC
bBZZ4RErjBzGZi/4yPa0BH15Hb4gTQiD9YPumKBKIXdkpqlaptjaPk+/kgIK2out
f2Z7Gw4EhI3XIgYx7CHIWbsVNmEy1LQXdNe5MbOPQ+ojnH8yXWJJx/ZIAZ3nHc38
185iKyibrMDFkUbz3a3Eb7RlFmkZG4wIP2WoHanwZF76c6ey/byDM1/ZAU7B7CUd
jpWyDEYY77+wdKP9MoyyjcMCq2lFigktZvUcktdJVWGfnXMhW7BMCZda/uYMesYu
5tGp+pNBUKUs9mkeMoA27Lb8AcRu0Fwda92Qt9p8ZjnAsgLIOD0/JEQzfhxPQ6GB
jfOh6Biw0UKDG9Q+N9Glpo8eAfyi2LfA+3xO3Fw8GQiTqSgfLN1bWIN4jTB7Trid
ttjYeQ1mJgBj5aIm1ZgtCFGmWbRlJAWAH9inutlsXJ0AuzjY9T8htojxJNSlrQn2
t7ZKmc8pu3M3W3Z6SlIgH041pywyWdEQfV/eL4yiMfwYT1jGDs1tef8o2lvTJME5
ME66I9loTrHtj2W/duzGdSxVy8OVr9FBaOZDtpUQI0Szu86/x75/3ee31If3uiRf
PEfF7+EueYSPgO0yTXGKLlLNNvdwy7xustqTkFFZiElM7UZiplif4li/0bjFdj21
1HqQ68Wm9kx5MYSMz3An+2VCNs3r8GZdYkO4WXRkJRv5wJUkUO0xwVXQwVgwtpdq
sarM8gcDH6Zrudy2ZdeLZz+yOHaG52fk8Uc3Vofe54wslsBipJXuIFgAybisIav2
LXSystJTmCClq3hZoh2jQWmH8bR5sme5zlTmTNtIeEEIpABzbyO/CgVXQkKOOAWH
TCC3VhiSF3Kx6raFmvTqeaV6hdhNyLP6A1k9/n3AtbvDceNtdtjENbcXCzFywrr5
LdS78y7fBW733nNFXXykMlS8W4NCgJFv8SrZklnR4uGISjj3WxJRGWHb6/BC/jfG
xk2w2xc2bV7DJEjh/ynXX+g4mPufWAZzBvDdgZUeC8s8i6ZK2CQcO81VjgeA4Guw
wuXnCu4W6BN9tVCSRGrbi53PyPHQjeqG3p3AE9aaaC+RV6n35tjSL1BTUUZZqk9E
M2YgP8zlor3M/cDOiR2pxdRVnwwQKV32PllUYKCOijZUw5HLv0FZhWvvlonlbJeR
hQ6gsJDOvQrbQQWAGYV5oQ60wZxlpsNPcuFxgNw1oCPGz+G72Lxv5Ik5kc+6+6QH
b4wbLVdFz2qBS1k3Ot+qPq2oeDwKVv7BF8F0vXcTIq8DIFxs6mrtpHmgY/B0FF/3
76h9FOP5MqrClIeVcz/HPrM7vK73EW1FMT/Psz3KuvJX+FejZeNexH7NZQ1cNtSu
Ex41Yly83B1CSTOKtpWPvYoq2RVrr7FZ+u3jqGvkj9AEg8tQk1ZjEsco8uLskdo3
nx5vqLSOmOTD3PwiWjIsBm68b7/Aab7+d0NXpezphGOG7sFWFBkRQY/EXGCYVcnO
XBHsD987f4M3YbR7YqAFH0pzBnq9ObhqM6jeMcpS/Jf4IfLPz1cWuPXR71DOo4yj
hV5ufPoeqFl/EDiSbkwta8UNrdRRQy3vCtpvzTywzxkpiX1LofbkgesSG/UUPpHQ
0T0rArHydRWDQ9Fy/KO0Q0j5nQBE6nEIIFClEau91hQgGCmxXVfigTxS3LvxwpFY
InHb4Z45+jYW/PyhDvEJ+Ty7N8guTQgg1+BMLVbIxjJgngc6OQCeh0TyboZseKxD
bhxuX8fnSzvBf/Xmv+k25j7YBN/J4NJ/rTqWiRCLUAhDrioPQoIyZ0deZvuieJKa
gEVoto3WEOg8JNGj/ot4llErsHIID4feUvYn00GqyB0GwdZ6ivetCTr4JPlHzzUY
uf0OaJ6KmhODlD3b/Nx4uqD1AE33ymVxsKeD07fnL7XxKWpCy/7I+XopFqbkKPuC
pWUYXbLsr2ySSkKdn8dTOYkFBbrtmicXmQuo+VXdBRH+P119kPY3MsEdspVBzi0V
cpNcQ5EKHTEljXIvzuoqUqOEmWCx+XkEmYsA+Ii7vEgjf6SmdcOHugTBdh3wlUjT
3APsSYxg+UWObsWCmh/JFIsXxYv+qzrZFI1XZ3eVsTg3won1XagJifPSBxFd6Vfy
vOEClQCGbsBh2zFjxDA/zbGmAp2x1lRHZjg43AJrArJR/iCDPavml4XS7oDylN8N
rhHKF4N3Xq6+3KoxkDu71m77Plr4micfA79TjpEMMt7fdORgayZk8sjwdCnDaftU
16kC4GbOVL40m0fO/xulKceoufOFwwV1u9g7/iXRzDWzPXcJo487PbHE3rTGVvF0
uPmge5B+Q5iS/Q8NFJ2/Fz4XtO3x/xtEwAGOrBo9EYajkwZ8/qNzEbKLQKqpFaMI
LFNLeCHxE6hbLaf9nGnLy7oRfcE70wn18zVdHWnH4qOBn87GRYzqBxxlpy5y6dKi
jSBqGpkAhZRAlckn/1XM5zTeIcnlu3fzF2kalZrWKF0+X5tq6Wn7xJt1r4u0Ed3D
wNwguxhVMPOx7QkEsKiMRWgyDnZIpvi5j6vNV9pnuwzVJ/iWFRXeVG8LNlJCRrN9
198r2CzxvirQJ9qjj0kph3kPBSH8xSQzwzYRZl6oq7cncbjbC6ByobcSTjLAdeih
EAcXcmHB97cbknpRxU6a5xWpfxru1Eaa5wzwA4kwtZ6MOLDfywWmM6dLR0UGdxkD
bRVGA309bFFLiP8S0+eYMR5WvW5bOIswE2RvKhKNcZSTu4jxNsta7TYXQgI+6FRv
qDV+Z6a+bzaSjEZcFInfvp+te5M73UlMRZYmPlSkoc/HyTVKXtIIVyoE1Hf2IlUO
N3ejeWGNzUZsO4AXO2PRMSe6QV7QLoMM9UUbtnZbDiWJtk8eLfpiRMhCZZGWM5/q
J0XCPPjJS19AoEBQX+M2o6mSLyHFAqkNWt2YuwUo1Rab6qS8eFGt/fZk/+gTc5O8
y1F++WKN4/+1ARSC6Vp5ZSpHpvWSbIJqTPW5WcvDU7H8ex3t2EODzizgorgIFTT6
nTgPpiFpf794Bb0YP7Pitg+Xm4XEZmDbBAH+DwvW7Q6XJAuRJ9luP9zmc+lZnkCw
daP1xUNS34+mVwMzQP5nJx+IgdllC4DJ8XDQ4yL/lELEq7QHsMoqFl/ObYkZG3AE
XacOIIW/SyGPM9IW7uI7I6jywmfRt0bNYkzlAdaYVfCeFF+CrMR3In8dhZUebZqJ
Xx12PyN3Zv4F+T3vuKwcXIlrxCZCeSvGffxcnevdagX+H7VjJmBjVKDvu9XA93nj
EpnPwWThyxh/YoYmZ+xK0xPGg0U22us3YYiCVMqWdA8nkzVV/VSFHbcaLBa4oVbD
qdS7cTkGnMwX9noVLPmdUDQHNU/CRy9kSOi93SGGGdz4rqWFDElrXVS6B5mDLsAv
jgqPSNbEcL+InGclAMBGChbuwCQfONp1QaDMweOgEt7syEzlosbmbjSFgBaMSmsi
vBVFXt2+DWPspbx4yHRLZuAc/Au6KIUQPf+m6C4ut2mZuWi53PHvbxM7pX5dTjZ1
OVrTDrurM7MVadt7EeJ9ILtKZb+s3NlJ1nlzpYprDjpW7mYa7Kp+ty18NzdmK7Ys
XR45QQK/zJDm+IAd4u/jKVhfZ8uX1MscIx1HA1IN/sk6/B7fGO6Je382bE/wu7JQ
5SR68tpIQh9kSGDpcLfQ8XNYTsOm9V+SNwzqvzCA9iEp7zqW6QqKZ2KHWXUufVqv
pXW/wNCTQgizrhNjstHYfZBi76ZYFWK2jWq2eBzcWEROKbuGNtb1uI9+a/IJydXN
N+1Bi5u1Vq6Im0S6swHv3ycwWSdImnAQ2QZ3rBCZ4em18/nW0EUB/qcFUmJVDGht
c5i3prbhslq+LwlWIE5+Yiixj+lfc8OHO1GCTmcz4Qib0WqSlGSnJh6xwT2rpAZx
AJYA3F1P7u5E5atHMabgq1GKswNFUoZC86QRHeGcbUqK0s8osD9+ohtbPkO5kl0U
Rl54LdWs607lze/b8wEhg3oAtAmhOW8CJfdwKIfK173ffUIgWMjwIb010wkeg7cV
qDSdQA2eCARxCRqgNEzwY/oqvfTHJ6S1jK96UpmSP1NdJuhYsjbvNa9wzfgguzAS
ajLt/e+WRqxVkHE7b3xhfdJoJPvYCiPKHKOgdGeO7G+PUGFVzOm/orN6kTU/A7+o
0F1rcr0OMoZ0zWxHJn+ruo2gZbA0/zIU3S+VX5al6QMKiVllveG9JsTwe9clQd3M
Kucu0hc2U/I/iE4LAQwwxVQGSwSQwf33Jn8jYaxp+gFJ96v5SqqyEJVaiQ/RD/cn
YnvFNUKzey+G5D66eAhOZ/usG08OQ7Yukor+Sd35Dba0rhbcLO3mrGH5Oag2q4sy
NO+52XfCcxmntaoZW1CaOVs4RF1B9Gn44X/Ch87+3RszgOSRrheXqVWhgSE5Efp6
ZfLoglU0eIuM/qBlIFHQanQAHy0XpRFCII4lC6I5kSoToRD/kvZsM48CN4bYs1f0
JiQmxZHxUVUyjKZVHWfjO2qykHeBqdyYuRBxfuhzB1dp0yCOkLba/1cBJFdzjdDe
F/HFrwO8oaB9CzHK184BGelY7X8inAdZapCCNAdWvgz+CPHYORsYgO3yT7PD4VIz
i6VOxXm0gZqr/LtQz1KdbElWezgFBADmR04QYEy8FtXawHgcFAxmZkGVyxwF9nxB
UpPEl2sRbQKBLuFRd+b59F5AwRl9np2Dnn7pTM6c2QitHS3OrXp6soxknODgjrI5
JrVQO1hbasoj9QD8AqoL9To7Naa8IRm2NTzV2ZQdLfX8HqpuPchypsavdeV0Eju2
sGsxtBJAd5bCr1qpT1O5evw1C3cRIbxTTvTo5dkbX+ZmuVgdjFt0+DKeOPcDgR1p
doKimOWWO/2kR3xT6uUFglQJdoaSDkjx/24PrHZHpHOnPOi5eROHzC39Hz+F7ldR
yq1UaViGU33BGE9OGjNLl5nP6OUb/cLQ8ck37rRmMFbTMOgBaIZrj6wz2IMlQTqK
YI5JuJqvXwxHVhaO9zRO4M3gp/dd2VnuysVoCOPKbE1H/AyHqw+lrXHGmQKoJEC4
itMNdYv/hXOP7vZbTmLqdaVoTWRDQVZKCpc2JdtTvpbvZj8B5i3bKe2EtYpH8BzF
76EYFjxgK3s+GAcP5yZOUhK2mCeMUu1GDB6P0sFaedLBsx7J6QevE9phpUPRtw4a
f4asB1ag0TyskHGcxwTgaXhK/mIfNz/FdAuqKFclZEMiptm8jjfBqniXUp0lsMnt
coDcgL+L/fAC94KpLw0uuqKP0/IL4Fvkw2PfnCTQFHaWv/YvPMGvI17yuPvkWOmY
7/eFc0zqhNK66USzRZxYV4DVBdRwD8RjeFZzRgwkF+nJL838VUIz+k3PtpwpZWfg
r/lF+9BUn07CsPT5IFRn5mHx+CggLq5kOoR50U20KIvz6lZTv9SnVWPaVwB5sXCm
4EEoWkC+dK3JijNdp8uLqf3dE1KH9EN0ybGHkE1kGanjzJQd84ZwzQj+SYW1UmyH
XrNBlZfyQ71LXQexxkNbbSGx1jaZQKOAgwUlU97oVl4SQ+YSd8kFr/ESDsWZa2ve
RptI1Fw0khBi/3RMAmQrhVUQTaUzl5PVkuafOuzFNwdMVGbfKbxhqt+9ucg/t6Kn
nSDs/XgV0YlWHLUh5mekP1AB0xgAhiihU6q5wW6QAVa5r/j+lT2DNoo8PJsloJgg
LqCQ/lH6Ky5TiYbQdzkrzDvRYr0tUdCK6X+wDZIkQOpnaY1mibJAgPKcdTlaW0Yj
D6IBqTPwtM4O5oRmoau9i19sC2VofYOmaq7SCH7XEw9HqQnXlk5cjOYNnT8sDV6r
iBLmJPuBaHJPefvkf+uM1Cg/j0UOrWQQ7IDZtomo+fSw+yX4aHXjR+Kp0YnPoYw7
E1yGIF10FnhSWrn1NjeAAWQU8ubc1oOE7+YaCiwzJsOASrVAp8Fqnq655VPxfuWL
oPVoGsU0WvK5YzSlY5REAtujag5QmMrfAm2pKDLgRa4b04ROHwGP827o2FUpTx+w
YJ64jbVskLf+X9P2pnUTQvcMBRPm4gakw3kQCll28xaBUA06Mmq0iHDK4mlw3hy2
hau5Yem9DJSN7t7+m5Zp4ZaiuBltWHfNw9246TnNoSoJoaS/DsgMDhSeM2DS2DMh
qUfqF7Q/8rm+Yc9EqWl60CLHxPLgj9jTbrC3IL/4leh65STVkbi9wErdcz/3nmEO
XnKuJqvFnqovLAbPqiSRrdIH4vsJ60nWsJ9QoPYJI6lTJA3JtjnQKkWhW7DwNtb2
Pn+NdtZg3hCjfF7PzTCedtTDLjpE4sEowJBxyKw1QdEnBHu5cMCv3PTLxgeQ3qYr
FX/93qaGRIHPJIrOEaT+DnnDRXoHNQaughaff8rMUSZyjOObxSQJ0FWMZbw8mbOv
xmMsRYjh+6/GTm9ZkFAhZZTQEpL1eGRAi3jpGLRunyqNU9nXvTQKyfjd2pfOxYgB
rawlfY0hnhCNOmajq/32H0ApXWdW+kotByo9Jyhb+w9iM/ww1vSji9UYwsApeWl0
cMaSKSQkZ4QlXzTykLCCEiXrDZyxHaGLYwa/6Iep3SacLHTWtywkyEjk3zL7X30E
q22zbnVvqBQm1JPvikxL3V+FZo/p8h7YRoeNKnoKIR8J0PULwkn20ahZ4IZs5YhS
etboXtKUHx4fY8Z/sLa34CSUElOea4eDaYnFja4IOU0wVP8FKn0fNB772yXh6A5v
ctZcEQghagX7AQ+B6jx43SLLve7H6wOMypN7MIp4Oa19KJcUdHhH01LvMVR5jCCk
9OIY44m3aIdR1pcocxEeo46jLX8aP64Bw9WYqpSSQduYP8OtiLvZxfz8mV4tQnGt
TEAGwE8qivVx07HfVQ03dDd8kJcSULa4oRl/AC0jbYM2k3BxKP9rHV/F5H/fg6hz
mJ0Y3f4xP6NDsSGieea/o16DoU/4GfCA+ZA6KGxDBhmYdLvuxGk7UfOULCv4Go0n
pz1GyagEPyQGsmo5bneEqnZDsuQkfwr7wcwZku/kae3J2SQy+uwV3dfSKCLzedp2
DT7zCADtYSy6f2sXEGIASx+gFjhTC9gmj5KFh2eizr6KV5IwQ/kKjSHoWDSUwYmV
/JPkCS9mWBI4YHmPFq57pD041almjamNge4mZ8lQOPoSmwdrvQn8r3tV7hg3YKxD
8FyoeHtW5T01Xp2uKUE4tBaRUO4vPcnN0qmqQVFzlhySg6LEO8Sl7TbqkqS38hrr
h3l71NC79ak73mS6WxstnsRlQh8+jDI06Ic0txBpkMVUzrCBO3WTnpS4mPBGOe47
CzVGU9I7mTlNt9dwvjhfUffFhglf++IK73vnRhaa90n3MMMZeDPMbWDyG3tRpGrZ
OnrJu2H3J7eNUk4UmJtW+4ufEhQS3UTSb3yiojmDRrIveAZb0eRdRfn8S1fQVfm6
+eNJiiQ07HYzC8xT0zspa3tyjbRsDRfKO+vx6yAVf48XZjwGPKGxLTL5/xF4ieTd
vxAIQ1UKQoon55lwLyFxwH/0zRmBEmGid3bowBWhRMiCeMuW/HWInIem2hKiSxzf
rGaP2aeOWdt3G7GjnNEPZbPFqcvNhdI29XuwPc99j/PzGP3Ke5GAoUvxScepnyjg
lYHokojB7yuQFBU4Um6LIsUs9G0w2p+VHsmTVsOhqp+vWyrJyEyCPxeyhW6PQ86L
H0k4R7OQU/v51vfbcvEbt8TnQdCShHhvw/nAa+z0BnBX0i2OTJ/AjlZ/Q0XCttAJ
KESF3Njp9DKPBDRvGpm9toWxdpvNLuWWCoqRN+g6VGht5/xF8TF7a4sKYhXd22W2
l9UTXgEQQlxYrGn7ArhyjyVSUmdt6ODgGwqyvG/vosgYfPJd+4JazInrR3Sdt1VA
+4+YZnQZCocGJJpTDSjGukARAc3hrR+JaSquN80e9NLtj6uo5s2XrxTqohyFfj4c
vjnTLM9yOv6IgZS6rO9M8zBx25bKa79L1oV2WI2dQI0lb3Go4i3pWqC7Ykw91Jwa
UJIazTEjvaPQ5uRtxfz+sm7oOKRA0QpDggBsOrg7OqRXwOYXCaa3cnOvgzfKEtO5
0h7XNSPO+TxSTfjNDC4d64kcVySS7baxRqMjuULbWUWV/0+zTmRvPN9+JPWK8J/N
St4xip+mlu8Txw5R71kXoNfqg7g1x5RLficzXkv7VPvuNXOlcAJj48tlzF8p7Mcf
j+e4a1BquqehPi3gzSwhW1KYfABdHZB0nILVN7VrODcxU3s/egD1xEZXCDNpplK1
bbIX3J3eYVimsYMkaEmfG1GjaIAljyxQesdij/7XXshkXBAUCU2sOevRsmHljmOE
p25LGdzXbsRk/JBU2MB+9yuGWItYpTJ+9865+tJNFDf9SqgQk6GWzaHNMVaZlY47
wEDvxiKzFDaeA9CxwjDrcvR+NHTNb97t+/tN9TrbNDr+DJJQd1BWjJtQnDXwn34E
yRhhMDwpk+2kNrCd5wChunySnzzvYVBDblnUd1eB1ujJAMrpw3UD70tfBJmBjhCs
QkF31G39DGFEW8sCXLj0pPkwgqbWaMuwKxsLe4AGJV//kuRSV86AJppIJAHZZ/7s
SJDTZZGGOcFTomD9tblKYWKGU6ybqFjLi/rq28ZXasuf1tbX2bHMTqTvfFSZKySr
QX3fEUyo2PYNuKyuL/KC7CWVTUjogAcGmF5hAThuTC5i2Y2A9ONbb7mgF0siXCBv
SKM/wXirXSpckK9tbCJEc3CXmCH30CXaebS+ZymTu94tfEcAm8T8u2p8kX8hPaqq
ZlEgoHglM+2gj0p3di1skRLnSiGXImqicqLOwJ40ICCYyOV/DBhf84fkQ6nvr0+Y
Bubhy8kV0334/wUdAt5UE8L7Lqm7ge7JCT8BHLJNxFLvoYQAFSU1KOT/OFBKO9wV
vZuEZnj0rs0R5tVWm8zpACR7wJ2YfsskyQmOoSLUx71RWu1Bp2lK5ugTmBeAJpkx
KH077isS4GB+xemIhQWYZ5w8eqhGT8gZT0qhUYpEdebWNVqwmuSKe6dopk+KRH87
isPdhia0VRrz7+F2YJFagRYBBJRtFH0DbPlm6+N6ebTseAiilkEvisnySTxHEQHF
+feVcquXWm9zOFynfsYeOYWsKDh3Wbz8ve8NqOrIRLAMOmtb4Zlyd7nguna1SE/V
klQW6IKPanQzcyeog3eOZ0MXhTJQP1KocooQ8P4BS32NexN2u1N894UsrSVeFWOu
etH92/Jci+Ee3hBNOdnP/cgtAKBxGHKuMZwUISPh5nmBfeELkW8LXDPHYKBcoklB
JyBKRn270f8FpIO+opsIxigluAPOY27I5IgqI3eUrosy+NoSbesg5rXnwFL2yE9q
S8+LHk6YiEciDkKZDv4jkJXM1LypYhORfZN6nCiSxm9OCPDFeUzpGtXXzFr+jaPI
n5ILG9TrKxUtF4D/ESKT3mOs4/bigBSkqVYlHV+4xAApN6TCUQgPyJQ36rI5TgcX
9Cj7nVYsikoMdtvNWoN4Ow3n2LLXGkcP0Qcmh59w5d92Gg15wj3C7BCwxXvEoH9m
t0ch2RKcoyDJxU7Cyh38VPDwo5Yk4DVM9BBFzQqOE85nGDgLXjseMhyTxQ83WMaK
VQOooyMhsqJPj2mlO1mro0Hl8uORFdd/VHbJQd3ma6HLs5pG79d6wWf7LsOFQuLu
Z3TLfXPEB6hnGah/fs8/WuIvHu1titxxA1c/YS6hEqRI6lFlEU16iXD1JPl3nOrW
j0OZIFgiYVFU0hHsYPpwwiddfy9Mq9+bRCzzRk0TsrqWrgZ5IQtKQdc4hMglpZBs
9exTIeu2qRi88iHETgw2skA4Ssra2d12oZvw2gG6Xllnt9l+4jgcuRqrZFO6XC2K
K+G2KShnwWpVJuCYUGdmB921RySEoFxiQmnoK4+JHSMTT1wmsFz+GQbeR19U11mP
TW3padwFmAW2qeOM0UKsbCJkbhqW9AL9a8ZatCbSK5EsysUfpGgvLFZHHBZvsK+6
AsORU7nmwH8KwOGO+7kz5S9yV/hMbU/m392KplDlr2HTVZD9XHA3WRpnXVoviBPg
QrqhaNnnE6XNliooUskOKu7pgXLg6DFGj5EHlFz6cUoDClxnhnS7mK1JrQ8iA4dn
0DByPoeLWh7WpCRLYZ68+FuNWCuMCUlxL4U3xKhD1ZksTywETGXZwfTuk8/lARHX
VFvePCDqGxQifHIgouXDin3uUDspgiZorqV2R5AezrLQ5qUwwgwwGEpksrPcNrja
cBieBax5PZpqmsrXfkk1VZBiLvHp6eSHklZrB1Uw+rZayXVZgMUI6+txxD/IGYKh
jui4R/rMBsT5R5AB1x8RX6IpyXvccg3VjBSXzFXWRIQCvscGUs8X01pPP4H7LMty
dhexlGM2smYJ0N3z/kfjaq7IN6Xe5iNg+uC4VGsgFUt+Knx69EECkexIKLd8uIVd
YuCqnJHzMKGmkUnJPpFnBAwGy+F0rufAXaS8mMULM6C0kyzQ7AFmhJbxFtWGdJd2
Wi/+tnC+RAqutdgmPMx4uraY8R79Oh3y2Blj5yCKIUI2yhogGT2XefwYrXkqngMt
TlIR/y5nNoeu6C8O/1UNSqHWytheaTBjEDUqX8qPe4UIuVA31NthFUmyo5qFQRaj
ogKb4Q6ur2yrWjA5IcnGnnwdrpASYv9MY4XKXdQdkjEF7UQcO/ENFBaHxxwt48V7
qn3x53XoRsfekYNHOHb3sduNE0buXt0u6GDvsNspnU+H1vnLPNZLY/E2Sy/4PSog
EqCctLazwT1L8JdkdUz1ARpREAEWtjJwaMKYBYz+L3yRVlR7lBPpABIs1jGZXcEz
0C/amWTZHLbk5k+PyTGAdni9u36Joe54R95atkTEuYXfq97wAAhqzQb5UI7UGhyp
OOA/fOG5a+6idWLPPOFRl2eBl3rAr9TXTNC4U3rOgex5lesfcZ9ce3zKUSWhNjCl
/zSS36Bel8iS82WONT73EYc2Q4QO01N2PtZ4+9vT2fHuGkgULOBk4SOM9uIfD7Hm
lSyWQoRuhO5jDaQyMTz+lFFtyLbljdkpo6OT5GWPQlSrOXC66UiPtN/wZNhnLC8j
Dgr3w/q0LS2QdLRsJPIGrTUt36J23O6g/VR4BlIThn+tGnHiY4yOSWkFSU0O6ULh
5CS7neQA+RFZz0Lmq7wsggwQOdBD8hU1gRaIpXGb8cYvgHC/Roe5cOUGhkazemZy
N1E5OauEmQF3P/vwbyfaAwxunjuemJEnhHIchz8QTE4Yq1z64q6RznIqAZ4WgnPC
+I65zPzRN8mt/oKnD51eDm4j0z5KADHn9+OY+wCIJNlfi7Q1bpJwnQQVHxK9IbIX
cHvHMGL3rH3ez93q8Gk4yWs0WbE2Zqspo6y+qvd4qHF7JZF2pTqQgwv5QHRWoGDH
ZnnRXjMeq9AhPztZIzFJuDyYVHGy3xr9D4UULM+Zsmcn50CjAAchqPfmcnJzW4GI
uW8X90YgD3fGqfpVlGX45P05Dd+rf3Oo/r9Iek4cnu2KvG1GgK5FAYKWqU49/2Vu
sGEDanlOHomMiR8E+yr8udoW3wr1aU9k0kuG5jC3tod1H3Jz/XcF4x5khgXipSWC
G0UOyfk/9MVtntsRVRHmqKNChorMzGl1V7YPvFOO4dJpXrsPBolrN1+/ixOeXd79
zZHdavCgABapkE6iP6vxAV/QVfWJQaF+Zz50hOcwS2KTOjsG3meWbkqL2vqpsGEj
gNFk5jvHQcaiFZVHvVtD2075ThGcG53oeYDpgGBHn8b84U+n5sOhLgN7xUI36FuX
BzLVgYsOYfcmsPXX2a1pfms+NViN2ruAaEpwMs+2KVoW2mpNAppsamCKCE1nMbbi
FLpa9ojqULrKjJnVCGobE/hld+AMXo3ADoZuzYiLe6Ajoduw/lkl/0fm30Y3ZfCy
vynmyIzYYcndcxoWsnaUPBfNMUdk4up/CntfKCkB5Mqf9oFzQF5QJaN43EQ7KC9Z
SL/57UBE2u7Wj4APAKkGmd0BBJcewm4f4E7CUwMQNpzzGPKE5Ox+pPYUI//jXGdv
LwzzhbBiPdYrS6wOo09MTCfMH5Yn2zZD/KFYtZaiMpr9v12ZaufSrO4Uy9W73XT6
p0TsJNjnfmAc6IaMXaYSdyp5bAR6q/Yvb6oO58uFyN8FMFjMaqlWKKT+yiA5uVaI
QbWIzx8CPc0b1tAtiP3y2uuVACZxg8dxPjf0dVynk+oXZQ/0mqR4FFDS8ZiEX2tR
bGvelxM+BArE419lPusyPhRmb5piQLAikktOj9AroN8w0Gs20CkAx7gI7IZJgdA5
x19lw5RrpIJCj3e78qpFlaDAN5NdlEMX8sqwcbs9F+4g9v0qvqLwbLR5YxNhcUCN
vLgMC4UcPDQjT5obtIXGm4CX5mcdTkwCSETrNBpWB+ADco0DV6Fkh/HloeROz0Zl
erL3NiffPuPn7PgqEeC9gFfKHO2MYruAotmSX/ksz4lvQd/i0KCtxFKMAn3gK5mJ
uMEkujxui7AtnQnMuUEkfZkjwfF3yYspNX4aEI/iSPoRBzWmBRYX+DTGfizSkI1k
V/7J3U+gUhl798UFB62DBKNTp3gzN+6yUTR9U6QP5X8z44+CCVSWSQuFnrtOdIPX
9VpwBxwkCCBC7t3R8UzDh3LpWZ8bgZPMzIKr494lV2riS5GlTjYF9oGmUMBcjIxS
q4QxI+2yaIkyD3LPFXTqgzC7OmURTvl0ANzTRIqyQWse639zPTlIF0I332tghcQX
igNM09HCUjlP9cEbTBmzv+UXNucWkgXAt91EbxX7tf6dJAxL55UyBquO5zZwr8kS
TYkd8k7gVZ40USlwGTtowOG16J2SzpjrYjndJOnozUkrgK7Onc6qqL8LnY4REtDB
KpWhLG46cPT+6AkfCXKefW0iZPSk73vkAOjkcidnKMm4mtCsPbW/MXIAcgxprtuD
6qwsM7Q9OBscmKLdJf8ms30Hrz1DenFiFFBK7Oqxl75KlTDLndPrA5KYDsx0rZ0w
macZF2T82WaCD867swWuYV1BAIXcJKPxlEWOSnZESLsuykMUu2yV7WCtrtr/8bYH
+hNvvna+pltmdRRdpZypsnj3Yw/b2Z1mCAxkd06idYuwzdUDd/HJDO5V58+8SAkx
j8OZTXZJ6FLpCBgQbys5KJmsNd9F8u8nryDqhTIZKQ6R327hpcCHzalsl3W4vu+Q
1V8UHNJeBztZw9H85fnx6t/LJD+525WYjBBGCzTexeFI/1PWgxz1cgTM6rZuOh4d
Zyv6JD99ZfyC1FWfAbxRY18bcVI742v4sw0MCibFIaa9VrXph/UpN3xvAfxRoJh5
Jwh8VpA7pkJKbEkdjByVw/FP+j5hdhcwPfWsv6nP5M+fDouUP4tEdf1+vtyz3RGS
yutBE1fRinybA0FMoZ7v4tLDew5K102lsAMi8dmcHVpbfeeLc4Wv9Y7Zj8W/UBfI
03+muECgsH2Au9dLY2pNNY8+7ijDeXVuFsCp4YMDFP+7kBGDlquawr6LWZ3qSgdP
ZR5cKG9ocTekq5Inc9Gw/r+/Sgbl7AyhkAah+V5+RE2x3UvF+RWIP/chocyGahz3
ZktGNetdoOZRu5TCIqEoiDjSNSsykRnBEeYhbvVb++JS/+HN0uExESTAcbbSYNFj
CQZoZNcFcmQQvpoq+M7S2fvxNLas3MYFiG2BkYLwuh0WKEb2t3Z7ZYL4BPQ6TatB
pG27FBn+3G151HNSaROBZB31UPnSJucCdeM2MJGbyAFu4KodCZyygRgxP8XC8AUt
pp4F2SD+/vzdQvUx1xgBDEKrFCToyAJDFHcnLal9TL9+8YtD/F0b8lhL4kNjsgbA
c9bQos5WWUH523JYNaKLu2GUdxMmNly7a8r/ycYH9vvWqsYVfFsaiRf5gFwEVyqt
FFvl1WHH9gy20eTyUvmtwV69z5njKU6Jm5yc0xj6n2wPuSloeuBHf5JGcmLwY5v8
Yu4lhchSht0j8hAWxkdRgOh5rF015gOysVIL/UvXr393m7m18FzBu+uL3oj+uUKK
m4AURvgAOp3UuzDNG4AuULUsBUWN5u6WW5EYyC5oXxIFZL5Jmrrn4MARwdbM/cDJ
1GQrerwjWkGE+4geXdL+r0InBr+sE+wQR9u5K3rn8+UFVL+SrGWMm31/etmwqZOw
vk7l7QsoLfYAyxRO97hf/gOeNHYImUXqJukPPyQ9cd3HLgZOrEzYUYoJK/buLOtu
w4k+LKMyb5WC+Cv2lPkRW/h8iLCArw+zlONjY6qGWgkdvpDwzpiBK+U3nlxdo1rs
9tuyyWziX0/u/YWy9IG6MFIvmKbqhFsS+Yp7cMO3uTtA3u35oYSgy3pFQw8gF4HA
z8JXK/lAtXhubd2BQCcnELvxThQk6i95vpeXCStDVKVExIZaOsZltQIueWuOmBpo
nMyHndsZ0tiziZ2Q25bqAGff7IOr4PXLSqkB171L7arwOhsjgyoa7t5nwzuMgVKB
1xvsfuaD4M2hcrh1+E6E4fMnJ+vU3urP0as5gIyR8AZIgFx7uBodYzdApZSScHCc
2beVmeZzycLYedbEHQQoG2TJ6NfdC8Py9MHu3KzEBPwpuweqlx30E6Wy5dmt7oHC
ApYxeEAo1/4NS6uYGrXzHvKAKHfWeeuetumHgbp5TDwYL/DCL5/iXQBUy+MVkqNk
/9J4Bs04iYLe5fijC4oar/rDlp5yAM7bW7EtO5dL3ANUtKV8dZ2BwDsZKdQgJi3o
nTgkF6b52uiwP8argRV/ciDqtZ9I9xd9MKImOkvrerOs58P1f+uKQ5H5W+XnGKPW
yjm+9b3KWmlcFQYxPvqy5ipAqHbEq0CjomnOzsZRhAbPSa2dNgj/Ks2Ru3+uL+jz
O2F6RmtbeZNnw/8smJOiNhqKDMzKCIFeTEYXWA1wohAWCK0Gpl4bPI5D9YHtDAfg
18Z03gr9W/g7s8D6Bb0ISWGgnsL5xdVAlXdbCqn3BXRu0tx/ppvVAKd2PUD9LZKI
IIJBAa4itDc6srfaMOfhkXLuhNfhd1jK2UJvcfKxIaLt48asiY4bMQQuFonwdG5g
05tgnPQf+dVU5mn1PwngwxBqXq/lrGdBfmhl4m34LT0hKLrg/Cxgp7YR8VwgTTX2
/TAMivD7AXMD1xSujhVReHltwVjgs0SEiBgJNgEptEQmUqAjUS4+fban7JN/fZhd
CjZ2ZWXYRnVeVyiO3SmCzYBFNSusUHKyk5+aSPBszC7VYk4wdoamNSieo9sqLfoX
3RPHNnG4HJEvRLYp4jJaCOjcubnf2O39MOytfPlVLa4cjN4We/+b3E62+TRVKkGH
IXT4nfOsQByP/1krpe9tV00/lbHJ1VOWUbImxFPGdsMLpihbKiWCCB/SwA0CcpS4
dC62ZaTghdQnbK9Qr0CYl6GRYGQYfPH7NgyAyBT10gFyvRpZeXXgGf58tlhcqLa0
jMIt9RQNwnw50WLYjvdtX0W2U0rE4FA/Ob891zP1uENZEf5PBtBIHm8juSmwQ8TW
3WVBE2i67rdps2L1qpzirQjXMCO4sC54oZVFgP8qq81eBeX7BCW+8qIootHWLqlg
9P3b/LdhEV1AHd58dG/5n47nln9s85Y2vYM+SB57TQ7v2LTPAHwSQmiMRfao+Ynx
65sQ/G46BIFppTWEUDBQmohe9SZmSU6baBkbjJs9qxJ01xSlirBDwalW/9LCEWyY
WM8vTTdD61Nf6CoHBvKrRPb7Orw3//opVF4t5aen9AasAR2HtIianJrU+ED3HYtO
lzmscZO++xB/32oxNozCKY1XRZCbM50AgAV+HiBCwCr4gmnEdty3sAeVMWC/L1+Z
QXnRohJ4ANRuJnKlXaArjqrQ1CqEIzfRHa+N/1OEYBBqN95jH//om7LVGnUgR5NE
ww/4JGWmlcYIEA+ULUbMLjFTPCcGrEyrJALZp1frUPbF96t1+lXQeU0/t2agDGYh
xcVa2oULw/tPPlxtt4JcO2kQmyuAWjzHic18fIDfCycv+LUyNguxGtn/lBBcxEEZ
2jzSajweOIXhxzruVZX1fDqVpPTWrNIX+4Qp1lgn7+up9GLaQvmnj0usjr5xB8G5
tuU5kIOqoYETQUiIPwTrDmXNXDkni08GOHpnyUwBVQzcNbny92NoNlnT91LwFE1O
n9y+kHRH/eZJ8VDr/r94YYIlxzYAnozADBal3ZQ9TNf88kZeXBNytYyo5IqLB49F
GQogSG6cSLQwqh9uYhe+4WEN/WguWbQhvbSeWMYSwrFTbijvHmMOed0nz5K2Kzud
vy2WLxlMmAre2QitBbeNItbwfqn2SCHR5ahkXMBv4erTMWR4OV1XU1vZOZz85LiX
TNqcAq+BREvWa+zlYb0cJi2eeaE2ly1QXgPjW6eBrQkLbf/Inoa+XTo4aeU/ll9W
3QhX4+U/tBqrTQ2PFHAcj/A+s0qK38J21Hwntbm+HBRu1X/w17P9ZjdoaZaYN5Bp
nsfU7AEzvEQlN+5YoQIw4ndAnE5wqAewKt+OaceSVMLB2dWV/ZC9IrzRC5GBKmxN
pdRP+AagyQbwuUTlAElrZDhpHRM8i5yqqpnEKo+wwTcBvkaBFK0lMkevIRslp5Xs
1o5coOZoecg3SusqBCxA+Ibuhi5ho/tnuODDxd9c8FylW/dyIyJXlh2ajf+nluI0
aKf9XvOX/KUwizHtVLLQZKW8lwKwgn+n9pLF1zd/O9S3qhyZgNxqqmxopA4ZlAxB
VEPJTGB3JbKRBm0/aUe1Nq9jrcq0PxsLsegK3e1PdC98KxZ8fLnONz49O49E0kfQ
Se0e2DLT4F1YFMg5B8gEkTRwEKhA+MAx+SuZimwB6z6s2xYP+w+/VkK0esktrpQP
Ms9/itj8y5lKSbCx+GgrxBNCXVPsJwiyRYCv9tHrGu3L8J5L4RuggrBiCloG4C/W
kzbJgK4/wUZyL1kbI47YPiTLi8A5Ub11QyoMcM8tJk+y1TN8R9qYZQudHJletVuq
GPO3L7kFWyOLvhlrnPi6sNjz4S77KPVOd8+A7ylkOmbW5HZWxI/OJdWPm09LZ9iG
1mGtN1RvkSXIp9DkHRvi/7lLr0zukiwiwUMcu6ydOcy/UOgwvMbjHBlvd9b3HzPy
S6mUHHUNhyLC+HLkaC4VqAApBzPl99+E4lEvMaT5rLFSPSBjWuquC8OwtFN/Hjpk
FXqQkw4yofEpfn5maXRNePPuMgDv6ffFDxMsIyri+hoRIYYOp1di5tonDfT3NIWX
p9/ni3iDMllwz4vvdLe00EA7+rMkewM+3r0yn++ljMDLelKO0Wb6JArUXI/vYz2e
vi0CpWI97QZ2nNY0zTGJQgfpGcBasUB1Z6m+2BjAFSe7MUGVlTrNDxDi+vx/rkjv
B73gSurvWqO6IArZRRW6nfKWZ9v6NInCi+KFQSfpI6B4X/cXH+TxcpBVs2PKdepd
FNJpYF35t5nCg56DB6psB2CeeHo+JMwzmXIKbSIXAEJ2wEurUvcr+kGwl0AgVWIu
LAM9WbHDdsiwN7r5g2BSM21c/NK0Gu4zdSy9sisUB6amu+i0D/XCGiUV7rvblsMm
pEOGeCA3HzLxSpm5vpFVxsJPhFPpxD3q9c1r9nSRM3pCBh7eTvt99gv2trTZgsZ0
RArFeG7JiWHmIjJR6BOMOjC77CJ/a7eUuwZq7DBYx0e9kdE/ONX4J5emSHe0MY9G
NMGppr9vHUe6dF7xolMTCMlB6RwrnFZ4FpZyHVxUFMV5nvVwt3Xej0tbwrxnVz1w
upHRUTEGE1gQOKHLftEF+4eaRoBBaIvBh7GQ12u1rsySN2NoWhu1Ua/erIM8OJgE
Ir/ML/0k5iofyc31aNmbAe7tziE5xK6g8t13zPlvF5BPnuz8WDMDdNftTW1r+RfH
f5sH5xG84KicYyYicRLwkF7RyiKFQCn0t93ydTdkfzzMFbbl7P8oMWz7wYt0L3v6
yvCz1tKrIJSpPzjTp7OaZRQur/toOb9WHaVeNlRI6a7t3P2JaRNklzGsSYcp9T7l
gsRV8BaRixBtqI7YW/I+VEvD7D3vogYgjaLEGZTZTMgRNUbIsXmWDAGp9LhsKyfb
zooRU0n31Nmum5w5+PNGVjkkbbLfsd9PLpbVAlXGenewhYnVXPgCQmlS0Fmtl76x
cEbaMmrSp81l4MEHXvAREne5Dr1Eb2g4Rkk3C1RVH/SaLT57RX/xV0Xcn0UXoGVa
nepCQLP1Tuxz0l11xxL732TurWJwo6kAgINCN8y6J42lSPPTTJ3Z+BK14VKH+unk
9gdQj8Q4epAb3NP/q6WtXjzFAoJwcC4Focf5h+WIxOCQkVJkma6ydVs9YVd5C8g6
W+x9s4wLoVuvFoogZ82lGOz05MFm3azp19p7buFNMPvuRJZU6XSuIhn7xBw2Pufw
8um52gGnYASI+WGdCJJ1abUDBSHM13kT2+GuBcDaQp8H9DDkYLTnvTbwWwRZheNX
yVKHTRkkeUE/tAp4XwKcrOXqjWW2/AeMUo+tWf4JZq+fiz8r7RgazKKmX6XJgicN
2KQjEZ4E6oGrQMw/RNoR38pcN+H48PMdkyfjIs+XipiY9YRXIgcvATFtyHuCMnWy
lYoWZoPEciejEiYYE13fZ1y43JNk5nwmoE3x/OR55kXJZ5V6aJ9OlZ3jQ+gGtUMt
T7YVXfXpADaxScMpOGuk/qBsUh1aeHBa+l61EUlehxKb64rhKSczlP0Pdu8ba2+z
FxWydCtxK1w8332xEJx1HOjNvxagp/RMvDFbFwFK0kxUM8E1U/84BWTABqT88Pt1
m+HpzpscY2fxSvYuICQPeyXrCPw5oyGeRhnR4Nu0EjhqFxbaYgZ3rG1lrgg5/OLN
ywnJaqBIIE471Fs0nRajSxmHuMYmaZICp7AZ5/S349MC+L1x9Ywb/0Ww9BiZqZnc
OOKa6OdHhP3TlR2J6N/YNv447qkdvslg5alW/YjWn7vAs36h39z8D1V8Ey39QqbG
MrmWwlygJHwWBODuJyFang8tvio+7bYn5dUVRvrYYIntTsXoI1RTr2obpq78SMC3
O1rid/EzAeOkXen5DxIpcUoluylnqfmAskRMVINUtOCF+fRQduRDCdqo2oWzeM8D
nWAt05iw9PbjBQvV8JX5Re9G75hRBcurQT3FQbFvYLQW6NDZZ4sfFFAdhdAqCeK5
SFYRbgYtlVkZrK5gNtWxW4guh4LcF4xp5d39eUJVtP+bEXBYDEGSSj5/hHRzmWpq
ExE8cewIlPAk3AP7D0Jija1tBQaSP8Cn1PsYluItckD9fRoaXuVWGcsxdY/EGE5s
KDaKvBZ/9Xj5z7yMLdYd1WSid5Jhhk9frnX1ylbuHWiE3Z8HEi8cGAxtX9zK+yVz
eK4Vf+DtP6HOXkjoVrcskZouBITX6yVvq5vJsUgztOuI+CdMlGSlMwkAAY1Vu8jM
Z5YJajvkYol6q86kU5NLUdYNxvWCYjIAk/4577ZPt5YhxT7j7yTv2rTDww0vSd+F
+7NsOxMjHcRlv3Gb6BnzItpcBxuF7mzbFV3xhUe6MM/bP4Wi6NdKjPdnSJjlDCkA
pGYzRxOxa5/bwY8bFkTarfDziaNgHngZOQIi6VMr0RjROwFfyooVTCi4GvzSeTYB
OYwDjA9TrN9Xe5hcHokqsUilBcwLfOsUw88v2gXcbuLeKWHjXyO6eRYxnNTjOh8w
h9uwuP+24pGkmoODpiCrQJ7QXu5gU+6rhS7T5AzNNwOJL77nk8XvZrxnAi8zU/Ep
uitdDTPf5NNMaXNoybD56VSDHn5n3o5jc6vOIcwlQXLd9iR87lfk5/s7056vnscP
9npFv3JA4aFXIM8HrC0NOhEaXtfE/zjqTJjuwwvqOErL4A5YqaXP74b780wuAfyT
hIElE4bO89zf5E2d36QhT7CfNCVw9jw+Ya1LIQd/K//Rx4nnW4anTaYvOOG1oozk
7M5xKcmuDm1/VUNE60sOlawrQTq1TvwJZ81HDnsKIFJSbCU9w06wJtALooDF+xBU
RKT9X6YlN0tYUI2LswtF4LROdFkTryexbMvQGGFEoWbUTZt7pQ6/ZFB8ZOA3AqWJ
HgNFf938dHkOqSBjf8qu6lcaay9sAoFehMaXqY32N6M4KIGWue6LQu3avHsf663j
fJN9K5EqVOwU1B8Vm/IUE0tu+VPyjwXeSeiLGLW/IUcEcAxnmHHSpvRgj4vCVJ/x
ZXJlWX2q1VXAfhkbd7TQtvrzd6hVLF6Aug3bq6xykCv4nKgWM6b/L5a8B7P5T+fc
mnExsC+8I82/UNwcQGPmcy9h95Fn4k/1zyDO5zH2NXzY4nTPBSJXmUBjok9D8PJ3
oI1uqejQQb71JpmA6mQGoxEpgmkyqLJ2o3/kRFfHWliOw+qvY7ZvJAyk3FmUm0eI
4w5Jwl9z1v1xgQJX0L2pqGpK30GvjUcbTYD8S9Wt9wGMAEjxZONzljZOSct21m2H
o2Ccuagblvp5ltq0G2Ps8ADA+FoNRLjek+hOgm0YDvxm5mc7Vuv5re0iRZZN8e24
5IXdKCEEkn2konbdVvW8HIGCNYUgb2qKlNzYAEDkr3kdaaEYFv6sgYTKu334/pP8
wgFBRvQAlfEAF18a+sBW4G5L0/BG75QXTW5uTV1L6w7iJJ/XBicZK4CF08eGiHIC
iB3EypoRvIWZ/eTdpOBRLhESaKZiNaUnc1eTJJeRQIQH86vb9f2C6+/TLDA+N/3G
fFJyxpmakXTtoN6i9dQFIeuwd/Eeoq4gyhf2+qJCxZZ53J9g9twsEc6N0Sdy8AvF
hrBgMiZUCKtAa0h6lDlyctCixIET4vEGze4d5wZRl/nF1SpUIwykLGQZGysS57Fk
xqLR5RdQ7Lm03fVMl3xnTUaA/SMbafnFTl1yydexaBiDNDXJ7N01+9HVi8F4ZoMx
xZ+OfQFIq5TT5jn3rjouyH2WUkt+lCZicgva5IcopoHtf35C+RMoBpchQI8Jgfn1
Qalol5UOSqFkNG8Gm9j14qlJCPkJMhAegVvvTi9u8XEKRHGvQXNAk4MvqlDoSd6K
bDd0/RnWgXyUlmNUYyoC6g1pOXscdhg/zUGVbn4e3oxkSscgCsVC1Nt+7mBWf7Ey
ud/ZLvgn4ZYnBdthcn2V3kDPWR75bNYNHchKj7qeMntOobTlVn0Ux/Jee5zSkjVp
ovD3KHM39LtuKjT0InfQFN8b+QeOctR6HWH9Q8xtao9jPCaUXEfUoF/UGF7EeoD1
wb1XuLDXWxy8aLsTc2NI4dZyIX7ArW2iDsO/xAWhCM3ENCjZfAS7RZbSCm8DJL6w
m/pLY9RyitlQ75vSrxNwdme45sQf0S59RgWRkXxnGNrXYrLMHe4Sn33tGO3FpJ2Q
XFHnoFJePIi4qhzu/MxLzr6oxFZaCjnapVFBiYKUmowpS6rT54+jveGNeen3sdMe
9mGCxx4HyNBWOsGX2Z7RPX2yhL67ronZSX6rRLB1utRC7xEZJ1gzIwF7DrxCPluR
UZIPHaXbvp2upeoTFjdw/pyHLbvmxqmGqW2n1RaWo3AtZAlEuCFX7MDxv4yGuNB4
IFbrEGnCIF3rgQPqdH/d5a8B4Gq/9/J0rn10V07j0x3oHYJI1UnDVZbq15yCXeBx
fLtn+165T04z1AM5E1CFnZ5TEtxiQDTeOBcf4EEj6bJpXEYkKWb1z1A0UAb76jDA
Amc8fOLR1W2AJbaB4f3I5rdX7bEfHprd7RQm+amlq5BBNZd8bzqqQa+DpyrCtuiS
iaK0nE8oQ+gtLOM3Vrb1kKracLcA51muxOtFVIQsNV5r2dEGCpBHFZyjbLHkV4SY
jilX8NhZwJ7qSLn82O8Ck5TRbL7i3fOznjOcaIo+UAcAnFULqzxqIjcG1JVUFuc6
vJEhiJB7i8MXlrRQ+VaHOpDnQ9Gyxfx6d971pBkoSu1Mjet8JCNd/lUAlXC9YuYL
rxrVGHzxiN9C6KSfXyXcno5LZfZ+0xNtwDqEqd+smuqMWI6kA+kC5VREK4S9feOI
TpZ+BNrBSmSQeLhIHACcGp+N6h+ug/BfaS7l0hXMm7Cvjs/a8zbWhPLGQmqsg0O6
PZ9y+7TQyghM5J4RGdj1Jy4s5jLNWCG6fRM9RL7VN2soaHifgcpihwWg5pfx9Aft
gjyLJZmHo2xKvfxZH9dr3jd8xkcUFBa4dUmtoD0mtaA7eOk1tc2Esj86YkxviM7G
aQxLXtPK/IKoeyeZUWMbNzPScm9wSSphAoVVuLldcuBOhA16bKiAo4jeIlYNYxzF
ceKVoGloaRzFmjPsXF2eZIxg534zu2wHq+A0dd9Eh5rQtUFRjTtfCH9W9ULo03PE
io8hv/cGjel+JOPhi6ePLyGA97pMlVzkQu3QdYm7h6Du/eB31+WPdwyV8j9IEsn/
CVoUH0/qbd/kYkcDhA6w4VLHZJmaxxFksLtaRBDfJ3a+9aCR5Mko7XSuqMg6TMco
KY7v9kWFL6e3rdyMeDOBSfn3kwjVbWmbYN3Qqe+WPl3vVSYL+NEGEc63PeftriNe
ftEKCMX6jD2p0KBADRWOVrZSHXwR4HuFdBZiFgbdhbRKoUU376mVoukoy6hAAwx7
LDDc2Rom+KLcEb79C9jZD9+sqP14JhgGpe0GhgsIADDCtJpPzKwqpcMvNGpqpU5O
YsbWjJcw6736mTW6XZtoBll5/vbBMbXaWlfNum1GFbSXlJzKDwFQ0D253RHqfn9+
3hIx35bYaC/ELYL1FWub8jvQBxxLD3+f8i2iZbHPNNBIHoq2LFdZXlcMKj67AQiJ
GnTW2sBY7Pq+4BPOFMaSI7FevPG3nE0zilVqwBRBfiIFCrAeZemJUT+1PwP79o/3
wMiTJg5/wjS0QqrRjA3q5weWYkAviSUeS80nPwrYTn7ic+ppF74Q8gCgJDcfXiE8
Oom5JTmoPMazUt9eNe1ZjKftxeUA+28UxV5IxzXrhGmnvbLbFZzqBBAzSRQFmeKz
uiXE2dME4q6EPtU2vP4R9aXluC5U61CQDO9ZvPbKvAvW6VqDe2eAOo8eqyKD20fP
DKuzMAXX9Js+dbVN0ytT+OdKlW4hI3U8FcF6heN+TbeUjR3RULllPbjsDTXLkNpv
gvHsSPY3vn6aIp3YojswgGGp+qy7rJhUb6bUB8fCFr+hRn9U0mCxERstTBwG5Tuc
6i6ANgvYSgkKk18jhNAN8wuxQDIE9Q3cvuuw6nHAplwbHX8NQorbcS/uLO2YfiIa
zpX+JhtpT7iRLpWTT+/YXaE5hSmt8kCX/48fn/ivRSnMwlnTPeLncoIiN45ZBYJ3
Fv2xtvJBckOLRFyv7Jj44Ng/EtzLCA1PZGzh34nd96ay6c6z1WMG0jeABP5yKOKN
dC86OlBnPxwyWoXTeSdXhmeihzUlEBOM90DjjD9Z1CQv0Kl5Qt+bwkUczGPscQMX
vK5ZfNQlE7Z57lP4hyFV2XBnAYkPiRp9lfs4oOd4VDqtxnf+FKPGJog6MLGFnfBG
66XlQKRkYhS4JGNKsQUImFhLoVvLUjyt6Bbi3jwq8RZGKyfK97d4EU/XGk5FJAaz
Fy5bnqkPPIAQuaaxS8HhC+WBOPuGuB3Mb8NCzQ0QWNJcIM6yEwcfflL0NbppmYK6
v6Pv1FGYSJGTVq0l/XG/mw2KJdgHtJrLhAIkQXEDVF7pTePLMUCie0/+sdjnFjtv
xqNlJeTxtzrFTfIz9z1gsJLMFC/QzSxFmLwP6AlkBxT1Gazvhn0+czAAnUOw7kDJ
R3ZIR0z5A7RqNmcoit//BoZ3ZIAUmygMjzVJi+PIUKor9MbDpWAQavWBsYhMO2JB
3r9h0pFibpG4qGdRVvYGEzeMnpoX88vWImaPJP8GxlrXcGft9nSvzuAtrRw7AYiS
5ygxLLNvsm8kS0NepqztAimXx6dPmp5DOpBuZ3CUyFEEz9oyZf/13f1oIWQtcKaQ
085krVkkjiZxxZSKqtN4ZPrdH04F17iHASeOxuBL6kVmilvkbzYDqF/zUSLZiESx
DpIG7L59CKq+4ehHn4P3AuluzlN8vTH9StvBp9B8Rjf/iUqSO1Ku7XweaIV9Z980
ExhA2yNcLtQfSiZxHqbB2xEXhbySEY0xpAjW4rSyoXKFcCFP3sbgsj1OB/R3SFad
BHSfjn+ucNOX5pUA3/eh/wyiVgj0udTEPIocFplWmBKcY/3o1/Jf55VOkr6poqtW
IJEiRLQ/qZohVPU2iiZoZMtZ8CKl7aIC4JAiFr0u6SV0ozDdqRTTZSbW1B3Rk7fp
125AntC93Lve6EOu6cFGOLd5y+ZOpOA3/XpVni+DIE7jWL6XZygLXELp1njMn6NE
SYiXihO6CzNvcK+VEbe11KigycTDRXFIkj9xPvKYMq/ypfI+RnFATlmXhG3uFkIM
EGH3/5gMLcUysAb1SIWzCiUTT5B3D0QFnrkqvw9mB29JiGm/kKAQ94U004bI+Yww
RfZlgZmZTi7veVP7/TRsoocZaB3pgzwZRRpYwEBhSdsFZjthJzz6h55X46wTCOYQ
Pjbomdc2hJ3lNY/2Qc+TkVy1Uruvv0jK5lcPvZ2F3On7p5HO4TIV7rKDx349RzuA
Yzx4ejJs30Q+VcNVSy7ye3El0tW6zZEPR9uX+CBOrTWyRWhRA1P+7pMmQKTE0zVU
tQ0oNb3ntKuHmIaAipqmKqNoSXhoGkNML8NigMXAzaNTlM6QV0zfn1aTEUVWgdkD
g0Xo20Y7G9/tUET7x3101/v5KhHAZcJHqwjFrNvG85pyQFbt2TMZd09Xi4nZULq+
ywoJviI7oIYaC0GUz+2nYEg4T3tNEE1sk2i10jaODVgRal4Tp2z503/lgpBXUtuz
zVxopFj2I0y8vbPCcrN1J01imd1rUg7mUlfLWBUYh2T6DuXblEdkfvDdMm4DGxoS
fvC36sff0mzOOMHpcz4PfNWKt+mcVKmcE/nZNFDageTUolgIG5s7XaTkvYhHivJs
kC94szMFg7gMqIMiMk0i+IcHJNChKUBB0eIADdqoKVpcNkAkxA7Znfj7ZQMvjChE
PxbzHgnfAYKqzj+7r4xlNC1w+1NWxIshN1zb2JLJpeJsmd5hFbByfhyrZAS3cVyF
IQ2wxI+sEgveh3bRF6EyNtqGCM5K9SEf+UBRSq9fuxcGsfyKa+AuXn2vk7SCxeaN
CzP7Re/3hO13SLLahVjWz91oHhQBZPfiZzRzZ590WbAFYgSdjUBP21S8Fp/QaS9N
iZym/5d1ol/I0QS00DQl9tfafxFIACUH5bJlV1JlHP1uOIx2aY9kyoE92Y75ZEfz
bDMU9KIXYIqhWfFyirCi17+QEp/HNejRdCNoijyo8zf22Z2oNwuSFJiaRaCgi4zD
b20W6rr0x8gu31uq1xIUYSGQbVuA4tdRqhxXJONBZ0QVMVxdKKUOWYQRRRPM0EYq
rrWIgmDWvXi441cfOBsaGpyj/Qv9gLterre3qODPYfRKe3Uo7gSqm87W7cuS8l/P
TmlxgaLv/N+ZuudyvuI7f2qM6xsLAhGVjUpL/d5p3UvAk51HYlg3LlfkBjhNf+bE
MxHk1UDVFdVp+/LrmN0QSkplwfBlj5/1hnyL7xuLQajJAIK9kO72s7BKspIC7+87
FPOXNTpYcXx3lZmBJqao/89NDbRcsednQH+qOQpGxDvCgOb6Xn7eGXV2qqwsKJ12
nkB+TIhkJehlxtTybpym7pUGpmswy0hcxdZaqLGXf42p85hSnQufegrcuzQRlEXi
XNpupNWLxa7H8idzMNTK55NBMQyDnnqBnJY4BQlJiW4jwNBwD0StIJAmTvdzDh0B
t1qDbke3YxSzEV1kQZCA0ZamsR70Rfiahxq1NFifYB/KT4+62U+t6ywgFyEPbJ2C
eutfh9HULcMRdQ0mWAR4dVWsHB09snDshubEjS5GDkOxrb2Wmu+gHrDN0ZfUOspG
QtfrOlcOUuo6CG2Rj3Qy1jcq6u82J7dtpomsxjuK4kJ7WQsejo/3Ok/fkd9pNf0C
jtGD/9JBsi9qBYAiIoLeaO2aMqAar0f/7YKOPeXn8MPTfmk4jDjp99QurMbGGTbp
mMzRVyBbO6ZG5LqxM8NhO/mgCMD5luWCQd73nDnHtiPk66b8Nkx7BAhWWqXqQDdn
dGub4R6ae/R20Qth3N8kwCVSAZ2yddr2Kvy23kX4B41d1Usb+LRIYrRemHcdzzpD
ZyMf5zT7F7Osc6Ovl8/FKa85F0t0h0QFzTQWZ4hHKLLL00eSTLa5mRrWZamfAtzU
io4GW6MFTFAeG++pkGpUzMVD4LDR/3sBZkelUuq8MHzHF+vvPIklu/WvdMDUAyTG
YTKJUsBTsjcJBW+XY6ylK5k90+gRMZyXYIAgvJCtOn9ze0wZm4LaL5Oo2yKcBcND
e9zafE/TX3Hk1tkLkEQb2UsRF2trTyJHZIo2+nNfXC2hxqPxXM9iE/AAwKNfsE0W
Kivoympr0BbOU8QYsu0kFzmZNy5EiCXnkSdBkIBNZSa2SgVRkBrUp5ncSmBxzU2X
I5cZMUkgmmLQkgh9CSHIqkgcN44pR0HfMkFkUuR2aEJsDzALL4bkS+xKu4NksF2O
yQ0mKpPjpM5lAwB/qhN+O7oSptj2vPBpzRvjWANIJGnCLZkFW7Mq9plsSdXLFDRV
uxCh9dsiq4Zm0mKS7/H7zD8oc8N1bts9tebGsCmssPrCo3LQah0iPeV9sk2FMAR4
mJUWJ9DekuffM1N1kGt/N9UQtDTFI5L6j5GRqbpP4x0ykR5N5wbGwGYXdDkjYt/W
xYjYbE6C3N7n+ckkyUzyri70Flozt32bV4Aphm/Nv9wS3N705u7jo4RkMVF0bfEl
FI3DK9ZAS4OseD8SuAGmO834NOFXCdAJOlolYjV2qteijACXoGUrb4mGhZSmqIMb
lWbukZo3PDpH63u3TqPALCBHMRsPX5pDtpFMBIi24McJDMGelH3F0s2Bx1LhgWyg
F6bWoO/tMqNRxSUpEgnJGhklNop0FB9+nIfhrB+MDEJnV8XvvuElUWEQ3QjulmgS
TistCM5tQysnHVnKQs8Vo0i5E1DNPSMat+SZ6/JBsVj+CNtyKe2mHUwlcB+XMjnq
8ZD14DghF0/e0ba8RVDaYrKmgfrBxMrWIJqrEgJ4ggl9YI85kXAD2Tw1/tEzm51Q
eC3L3mBNlJ0sT+crQu61ul7lSeD9uG6I5ebXSHtNT0mLkKCQMnZuOTOYSWbVcCTF
xtg7cIKfftXX8UVTjEh5JGRyToDbD1W7CR6C12xaVzq7qSjej23dJiQHuwKy65wu
WXZsByHpbtZES3vcwZt9UWXgaiodA8nFtGnfZImeT1kDaRvuOSCP67Qg3ueu7YKP
du4oppcJPKZjTSLsUyfTigd/bG77BjW/SPqvzpGUShdCc1NdowzbFhuARYhAS/W1
Pyai/NdGc5efVJUB49a0iGX1JzcQfGagmn1pCirF87kEO6XY5SWWON+g81ymVdAk
Ujnl1QhUi8LjcLK+KmDA+e71SH/hIpyAr4Ze9bMLTLu3cBA69EtGl0CS4Qg+Gepe
Gl0LZJRiQwKlH3RmP3dpH79ueJumuablMP969xrpaogDIampU53gG4k1fI0C8ypC
qOqDQ3flaUFeiwWMkNMUM9LL8kCIolGfrxCqHV6iyj4q9bTHfSbd8RtnVoGHx8PE
YCNffxyQUqHAVWopVrhVJ3V1T76ZicYomkEO6roWwQDxXSjKs5hvluxWxPMEeoal
JxaFFQ5CUepXH9M/Isph5M2fgrYBg/2im4hdUYodMKxihTSE4qMuWceZ2uQ7iew0
GzIg+00XzXq0seqrS675agybG4W+a4SJ8pI4HtcEUcdKOP9Xnqop3DB8+ZGzxHkA
T8cxHt5T72HqIbgv5GlXIp80cLraeKvXZcExslMXSUwnP+opi0wMGs2osIVLb4rG
GdG2UUGtuTCmrLXpgt2toVMRFpdk074AW6LfuT9pTEEvHVBiRjhc05GGvVDSAtuR
L6WFncanXKK+9WJjwCRcBHnpkUXnzVjmPj0ltEPRO0RbaIJHWWgfNbd8zXJqTRiV
t3EqaPPj3lP0nD7jjwRoHkQSwBOR5NoUYs9bLCbmeToMCQ4JiGIq2it3gn7XYkGA
fYNj328z/URegQRsZx/BUY36FF/yBnssjw4Jvs23m4IRN6czNlWAOXWcCWQoQa2s
/00nm3BPWHiRZYTrZbfRPwOSEluF5vuSTFBk8sBZckY96a6HIXg58ZSp1hyFRTY+
lQrT0G84nVBayd4tOpm+56i7Au6ggC98R2O8k6xePO0OWOKSElSLEO+pDjMMmttI
09m1NQwSn8pKYHwjQMNW56JiL7us+B040GWSzSDk99kpC1Kw2P3juxZy71pb1Fb6
Wu1Se1B2r2NcclPj9TUmbQH9eCBFgMQyZaPD/LglQhh30wRQqbEMoAuTwMgrb5vo
jbI+RskzZzwRmw01DbXv/UHk6NWu5Ne/pfg0mPaNc2kA0ABCWj3uHYPsckkPmych
E2utfn7Eahq+lqSDXeyWSWQMc+DQ06+mcx2VuOUII7rPSdJ1TDOKzQQ7tjQaBfg7
dYUT+7Em0GMNrC4KRGAXWTNNFm0/N0jK57lwyGpOzKDCuVJZKFdgoEXq+C6T1sBt
hAYSPe/xt6wGqEHjflHGVk5WWAt6KIwG77bBye4FV+YqRHQx50plBd0uKFxFEBWc
Hy8aaLAkNbK2ukB437YsAIBTTpIJZZfcwyL0mLGUU2q1iNSJPvAHApr4doAT5ttt
87px6nWzgcBJ7sEa/CR4ZM3T/1a8KM9qlalt+Yf61c24jncHPgfSNLzSy4ucebQ0
sLRhzWY2oJLPzVCSW1eWCLBGaYWpTF/2QAWQYOMn3w5yRIMzNvde9HkKS7T27tB5
Zuynlf5yNQndPI3wuAQFsKih+V1N8zHXObU/wZEembGRXfDpmyMiTfEgvYHEWEtZ
kyECX7Clg7/AWrVmV5+G0IVzkx0ICl0NarRT1qi2UQ4aW/OgmuLGkrjV6d+SRPn7
NUgRVsOCrik2ukyl57uoMptNxSvAbOXsvBcnC7ZlAEpkRZqS0eLjIyWZ9steE5Vw
9Hpe5SxigcyO6bobmdzfe7qjdBEA4T7r00i64AL09PXWjp96QIbddiDdw4xmpqrB
GgmDhv/hlT9CmmTmFDqEWZjeKs0JK+MuenKZeBNGWHqD5OUTBpdR6R58blUDEGBL
oY4lKX1IgpPf6WMIdWsaFJ089Dlb6KRJi9sXQhiyY7cYdt4O6EyZxKMEbi4ztpb5
rV6gOCJ6u2/Yxpk9pU72P0c0h+8IJrMK0vWHr6Lf2JSEioRuBqK8XHkS/gprlunE
L0dMEMKhVnbXjZX66lyqKuPESa2CIqWX8guqNtpfG4C71c7PQ5VgmQkakLFDjmtx
Ul7aFyDP/n6vmOJp3GL/+qMX4Agh5pLM+wJ34/PVKlDEeMVYOn5eRgHytS+iOc/o
Pp63/QX73Z3bYefjA9lDH2qvAIv+SUM5viwgLysnGiYxI3ZNsj6Ocwxy0oWX03+O
eOfmX6Xj+s0AZPsSbSxZ/zmt8U0vQ98x2KFazrvCbvuDKWYLtAUzDXoV9sPwkvts
CgzQgOALbPM9pCpoNTRR2ZqbhbzWWqyo4Tz1sapAm3GTsvnE39ocKNXZpRl+oSnl
TzmFEb5s9tbIVY5ZFziO7SmpDx+YJBSo4RztE1eB9QvlxAzYpUsQlkdVWRTRz5fQ
loZ/405HqgQiPZ5qTHUpEtMG0K/+7svYrYPgR6lVho50IQB/OUBAG1mNr8k96qHG
BA4dwh/ALmly/Q2QqbYsC2I7QVvgj6Rq0FkmhWXtYNjp4r/jASC564YPiCr5zAIa
HLF7EM8b72EAN21aOlQ3A82n/q6EaZURKh1QJ7deBiXBJ4NlcYRlEVbnezorbnkM
nZAQ1FXpph2eiT7mZ/WXDzl82C6Kbu2V3PO3iGHv1YY8Yhdn1OKmA6aoc6eUbK0S
QvaGTxvZuUn4eQyNIBUF/lfy1KlgfViEVyELSrkZ9/hbQCsTLPFt8HS0Bo5K+Zub
g8Bs9Z9Y3Nu6DlGg2nSRVTkhtKYqLPsfoNkHQpwB8nlRSpC05GX6z3vXij/vUSID
kwuRstGyUCgLrGkZPVPsqQFTKgfNI1x2aGVcDUDEfr5CNeepGWisG3HK0DwydaJT
9gZkY2DL5/30m3V45OsHZ7apqCt1TWwXpymoKtjY5ZHTsXVpf+kaf8yskEc2bSnp
LWyTb1kqgziKWA7gH03GlbuLYAY2orlg4Xn7wWDalVMWS9BcOJ6Comt+RDBuhG5R
7WO0ugRR9/fybuaEf8vErhzc6CtySsWI2kliYeEtFT5cl8pg/S60RPyhUc+CAy+S
z/c++BsTGsC37XjGTMcxcmAvwWtMEvAKlJsY+lcegTb9qCRby9VXICbWGt8T6siQ
7mkzOKxQI3FBFiv7G95ooQTDSLretE79quZDujH2UkQdOiITGK6TQOoubOiVSseS
hzGhvvJan0GR2xzjrduNk7ZxRiQuSE3Av5oTJe/GOFXv6+qnN+mFD+A1UHo8mSOn
nUMI5qLfv7bT7Vemet+m7LfPD+P7VFa+Cs1t80oHpMJpKcFb9Z7CDVZp+i2FOoz/
+zx3nw6s5V3F456eOyTg6hxKskwq3AW7mNKCtjj9zj4aMHYU39z+vAPEfxUiFwgV
ho6blnct8TLcSaQDXjmrREMocD+zzeMKKEH66B/giOAVMaYR2G/k49EuPY4YKasB
QuSDtR+EtHyYY1mKOa9yl8ZF8xs9sgXPLw4JVAVZZiusB5oqy18EtqqJsuDZc9Gg
wiZh+z9uuy3O2yxNBOVOiBC/iYmLTtv25cIGKo5mOMvzF16XauTIqb6ANLhmVYZ4
WPLgr/Z6NKB5ncUGFEPYgP4itjpCJyHrFbEVia7iKr/w0r4gACxE0vf3Sj6uOnw6
8pcElJkb0yZbLCJSxMaxvFXar7ykiuR1BZi5GlZh90R9xVCYK/2X0jaJWRFKnPo3
N8pVMZc/KpJiArZ1NgtozCrD4xUkTN5djYlJKfC+pEhn97IrOfVvwH2uRu2iq2aZ
BMZvtf8t6SDrpifASEwswRX4UhhwNmXi+T3lQ2rm0n9RJaM+EyR02Hs4cDsTMPNe
Ok4iqAQy4pFYhg/Lb48T69f7k77uFW9gml/WSDst2ktmyHM/ergxl6yPR/k4qg9H
wsvsfBhoLPRMfGRL9IeyBcKDgRdcD6rxznpG0vuQd+lXbIVkOPOaMjvwZpo6JSXp
NBsS4cmwWZaU19rILJ+cUn74D1BfK8s7R77k8hr7oNLu3j006cV8/TUJRi7yTHjW
YE7VeyBp0uTYWqk5MxOIDoICyAuJ7o2DO/STS23Z6GY9ZwijWfGCfzlDtcjcI/Gj
Pi41BxfMRV8V3l/JAA34KR//QPZFMbnqZeCVHkhyieov33pKAT8WKYZ3YgsSH4sv
b73h9+A8ZGqnFNaQCa5/ycSdpc+Z8meg1HTtTFJ/1W8bBQkAZMYH6xlhEQLr5hBK
PGOLwxsrzIG6yukT4zJW3/Q83JXO2Cc7hBKykkiB2JGbanOJ4TTO7Xu+hGnsSN3C
3CSu7WDA9vXMyNYCsrdj+k6Hike9VCsKXBt0c7IS6Ad44C4Dauoa7UMLxo12vwb3
pXMVDnCfy31dG23rk3XmT9iYjqHSvukJyZPUWUcSGBtV8SYdXx9t5lXbto8tlhKy
K+ncE7ZcOUhI9NyzUMOutmcJACCI2oh/PUFGhEfBRituPbN0nCmB3ko/zTZWY0yc
j3p4xXt3HX/K8m0uw8RdE5uqavTwzACE4/z2Sk2s7GP1Qq+I28JIV1Djwdr7/t4r
IIV9OzSijEwL2/FN8tYn8ZW11D0Fj0qMOhiH3df3qVILMkuTbf6nzTCdEV0vN6Gi
J7ETQOeii6ndXKL7EK6QV3sGi6j3x93gf5ONnRjEPmXOlWRy4BTXT4s0wn5Pio00
qspIy552GbpsY0Uh5uuJ8RXWCaZwJBtF9bSmoYf3MlKjjqkS4pRwJ+/S59E7xrwI
+cuw6qSaCqvTKehokfpjp/79NcpUib0ebBf+IVP3isfJ3pVLxSoQ5Bj/huYWTGqr
GoDbuj/Ic03VMrTjX0+cDpUcYZGmZlWOOzRnfo5pcyTF9YYxJQYps3Tyk9LOgeSc
/kZe10m8j6+qv9aBZcCiwfoorfSCv6plWP4KydsCL061HyTV1QgkiQvTQKPRpfpC
tWCpWq2JAjWYkzCK5Xf5zak23JlIFLboiUzH0vyWTHyHMw3KTdU6TgQMlY6nCfBR
y1sxAMymxwE12y/lWul7+PecH1vs8pcvcXx9n1PSDFKg83iGi8EeN7TsBEUXrnFF
zQwhKKoILmjoL6zLkl5EivaSOBITdWJZE06Pt023l58hwBVAQ51+EoVr7csx5Ebe
KYAYgGLGcAspr7vvnKP328WoKYPyamBkisOZ5ru1JRseLAjI4MwWfuOeGKL/GHUJ
wwhIVavLMzszxFVy4HluOQldur+pTwmu5IenkiqB975djCeO5aM73k4mEuYlS4ip
LmSu0bCiCcnQkTa+Buk3WD1JHAlX9aSD6++E1d+ph9TPZ+/02MIDES57MBONrxpi
tiYRa45GVNRAYupSZ90v4WPJoWDmXig0SqkU5BsYITIW5fQ1n7tkdc7ypmyB9KQW
ZCM5DB9REcLR52PkZ1Cu2HC3AvGl98IQQ2Tkud4IhfHb9/Drcm489NTZ0g5xFX7o
PtSqi8Y8xMRhBuHzFdpRUJlw3aKPcogRJXzdlyAvZHTwkMARFGVxLaA4EDWHWy4E
otaM75mcIaHJ3GTzpbWNCl62IHb1pQN890frIhHfPMYtrnvTx/lo3oRrS4P+ethd
NXFg/Glv2xQzTzVNWrFO62qoF29xeUfqHvtDMbDJsXh4oDkucQH6UfbJcb2hkiLf
a57F5bUP8F+L2/QnldISfo6UCdLDyzU5xZM03RyUjGL0Uy8OWaFc1TDIdc51b1NR
Mxtao5fQOGcRi6lgmvloeSCxeuXWbN36uEzUEXiOxpNeGTFLfPpzGuAQ44agJRk2
RYgp3x6Kkg9u6cqY5jesHG5IbH/CySpHaHowRKXDpzdq2OxOQwGaNm6XMYi3W/0F
+dYbe4Vax86kHpToDUXZ1/d94P7G8rrQpA6T3Ms8eJl26xAkDd9C7z01kR7wtaMo
zWumUj08Ko/WBQ5hrYE45kKjiTecjoyOAIYfldqKVBpXvbMqO1g7NaZxCfUw/UQZ
e8FIm6RN+j2bJym1ccIC04k3oRwjmDXARazds3Bh2H5Du53+/qhibZGnVp2+eSOj
a1KBw1U+o6ZLYQpewiJLQ3CfN09fpAaSCdcXbrTNpSOofAsV1lpV86sWZxL+N9DO
HO2KFYMPT9ZB6kEFxOWTn5fRWvNwuh5bH8tZWBwv0NnwRhJ08OgL4OLSIbrNHK4L
5q+UgRdEbD5W02WGPr+Vo6U/5qoqF0NIVWKR/vCsBNiWD9SXvhg6bvyllKmts/4B
E8XXvbnluLR3JdY1/UPp74YOtFqeRPTEPBrRBfn9yC3eKBlzO+waV3sqOb83BfI5
XfKaGdtbCiP5SH9PhWcgp8aXBCyRVpX5dGI3Dyjd3FPkDWanvtoir9mIQmRjz9BI
sUeDadA9EjLNQFDtYtRtThlxRqFuuMOwccjcX1gVlX2f6dOyQydBqhSAxh2ISA++
Ki/4amSAi2ZhtQvgA2C1DEm4L7fXIwteDKlbi5NM6ffnyz2Lb58x/PFGfyzUjNvz
PzoneDFbbSLGQS4yaRhN1e8PjmSppRniqBSgAyR1Obu/PxNeTOiXo8riSwraHJCR
SxJq6aLPzbYJ1Q6lcRyoBkg6gVJu2M18rP6JHGswwkGKJGkaV7CIr3fbuaASS7do
B64ZvasPPO+KxlCwD2+8KhCcz/CpRi/uMjglhhRxTQJKvnQMh7DPKQEodg3WJmOv
pb2zuUkxH7PfXTItet0UcbQ3V6dwnQWOGNsfOFWmdIiPqni778z4ri3ihnLfg9bo
MbXdijIeW18KzZETRKbLm7CZQIo7wYcGAMCgbgoi6KEjk2M7q53VqZLdrjMLcxHt
2sTDUVKlQPxK57eBkvkOZPdvhHvsgReRMoPCPL2w+Q4uPxoWurVsYq+3/gOJmZfB
jo0DpnGepBvT5YGTkbG1y6p2YTjQiJ/7qDFyFnjSQ1YctEy9PrcQjVYx6iZNsftN
1ZHEhbGoJfYNKOYtppzJ2LfwjsO02FghzRShuKUkFff4VYcrxJXcQ7XnwIO8drRM
TlxvapPid5E90KOJLlnol5qM3JGubFUrLOQqiyOnIfRJi8gObstFcxlsHyTVOIsz
+L1UJ3f3Y+QDmlrMRLfctfCB6LByzCINhPwOuTokMmEr53zKK8Wg2pLcgEMserc/
mOl6+b08lfVhoxLpsnEH40hqs1OMz+Lo3PoHMBO5pFTkPSTH3A/WGEh/I5o+GrGa
41XuJ7yK6HXn9nzkDZ9kXpPCxbeDFP+Yui+3vKTX/dTUIMqUfjC0lFxKTHD2EXrM
q+a50uQ4s03Tn7vbfcUxIBESti3sk84grQC7/ExqVUwqu02YziBk1Asn4Wr5N67U
KEoBtxo/auCQRD5MuCvc/v6JM4z0ooDkx8kEFTpXmZj+RBjgM8I6U2kOn9y5cpw6
G6shWHmj23XOUQg4uOWDFxOlqjbo/7s/AFbk/JVOitODH9+bWEzSSCaCUikEGtH0
vvqCPUuyKg7Goyy9gEaCMWXZT0YmdpuZ8M+yX54S/OttVpz/KsTxiNlFONXX5zb/
eu7IXHS7CxaiQ92nZp4SOC3rjU93UO1cwlKEsfH3OKBbgqBhFL+tWh0Dbj/+M0Lp
tuFvxIZpv1xXQYEXT77mk6HQ/046G3Zw1uNtjZHNMoQlIWIgQO7Xu+yBO5pX2eqj
P5SD3QK470lKn6lIGru3qFvZ01+pvj88qRT1gfNTHysf6r3pBuZZZcOFHc0N49MR
LPj87sk4BCYWDrkc6vNOFFnqshD3zHvWMxhKWtwBxUA/YmHqxxvzKFxQgvubC9+6
wFyTUFxuFrGRMzbcTzJeo+v38IsGJHyDWTb9ngck3MbAG4sfo+yhU86KWBxU5t0/
xFfU9wxQn2iq3dftmMerHab2Oakq/1ypokZYjpNzUyKyUVqrDY9Owr0s6Wv2oMcJ
A/ISS222MjrxMJxxCsqsA6pxXa/jOZQgsuXVuHx/AusioQdJbWD00Kct6dxmENIx
wWDikjsiwXe9W0krLfgCt1PiIzbvl6Z0BuUV9R/EdPq9FeTL6/V1bM0Pg7nDAl0E
OUzLW8d/OMof+0coCfB4md43Z/r3jyEQuXTLf0PvGrSB5orhvb1CSAMwvVBxiMFl
9j321Cx7tfS5A2moKpFwPg5772Zdh4FLBbc4FGxCrVxPyOfuRAJxUMEGMwy2bIN0
Xfsr3A0wHNCwYd2UeQjg0dEyHUr0E5drncw2+Lv557zFmpSrhLuvb8W9lsZ1So7H
9ZMOfrODEzhwcxSfzl294xxPLp5VDw/ZXGOwVsnN19eqEaeK0GsvDiZP5RHxebIN
5h1RKnHfHZf++dvbXox3pcE64VF4cn5x8UvQuDB9VTirGBGU54c8Dc51SUTCuoFb
5ZoU/foGcghQfsgfXb5fx+mtiUH6MLV2R6H5UJuEDhEGCoChQolJiC8wcgqs4Aqy
WDFtQa/xQBEEYhSLWMvVRjjK8sDJ2qAFd+XXNxfZ0Nn2TVohlzhsYHn15+YNFHoX
HYWVqwO9r6P/WLICGwubdP9Z3i7gg1PxnE+abwiHczu4TIxT4fA57i+GoAUuLjKV
/4h0ydvucy4mbzImqI3f9NsrSXFn8GJ1k4EZeNMc7GKc8uabP4W2Vc0iDWcGFL0N
wxRekcwWILKU6dO6exOcWwlcNTc4wu3KS8H9kPQkyQ4//RP1QKqksP+xsGM6BVtX
CIy1SUiI4ymtG45hTKn4dUVXrc6OjlTaFMRtgmuDSI9PMHj9VVElIBbH1yhdsxZz
5caPHkUaJVRlkt1sMFKF3nTdvlm3hQqaQDB/nCits7+Ft6I3lk6ovGdUD2GOosIV
/8+QHQ3BabpHPr0NOezGXDuWb1AQjJp8+tJqdnnO4qwy4NWviiC55EeI0zB3zH24
/swpw1VXv5Boa70dxwryzmxTMAGKURYgwXRVX01322E3qKwmPND7hAJHHZ12a1Jm
j9ElmtWnxlJs1YwoCwCxZmoC7QUSqPTmb34HDoiIq4YYyFQrH7C7EjpxcaTesLBi
N7FNrA5LZHjiPAfabchTT5nkNugOkDqJidKLtrv8mLDDk//zeNj6+RBoRlp+ORcc
GFRypV+bmWVviELs6W/bHf5+HlQTV0ZgdnVE5H9nxbBID0FbokgEMkaIKRilwg5b
jBNAB1I0ES3kPEPHZOvaIpaD/LGrJRDag+JabNzAF4Tv2Dczqd3xMzkFIriWAvMR
yY/ZCZIjuzz6DnE7TnFEvbWDhS217SIBGY5Os/3elV+k5WJvHpLkemFfOMwvpcFu
DBZ4eql3uoEi1WWQ8Va2x/3AK8aWeJFL+rj1Giy0H5qRLUZoO4Tmq/rWZRItaql8
GTmugEiWQj09jX67XMwQjz8Ot90rzeaWFb+i66tLSlsvRsoMMksjJGUh281F3vlB
e/jWmOtoWbDKw8Skez74GzY8D6M2bNF7qyVn513vL6NUB+zd9Z4QhCLZdqLLSr27
P18ew8Vsy1tB041PrjzGJuZsM55SpaUPESpFF05C2ZzCEy19GJFa6/QSVAe0aIjA
4fbsecXnP7dUOojmg3sD0mRr0JuhM+Tz8/j7voWH51D0CmuditEvakcBzmxMvdXE
dMcbznfY4w0VElvDmin2T7BVErWvT5XIVduegKvKP41CNRgpJf8tlYI0La9UBC24
JD0G4VE4I8a30sw+TCFoK6K0myKfpeJ4QtzqMq3aLTkRu4QSv8eTnn0kbQYlhUat
GDCc5fnJoXtS4A53zT5xcPStPwJSCanaF/m5A3B1F2Sda1mXrhUUnf9iF8HgOERZ
YUPqd28EusbaIuzXfpbg8atr+n7ou9OhYKMwq9iDDmKmQjfxpCjPE3MExCZRFxFA
ko+KxNX46ltN2UyM+AdcjeDyPAlsEe0peN34o8DA3B9F9podsKjztA41hP8UpRx1
19aCQMiYjpGCrSmO6pDRJ0TKecBQD+tUeRpa4GX6t0nQ6wdPJNS6DA+Dm7mo2HZV
ryurYqyjlKlpHeourXrMksZCO3MS1cxn0UXDMJ6VbtKtYoq4lTUAHseJImlzivRS
H1O5pUMAOrOIjwhxrLw5mOgx8gssShMRfipDshZ/iWmfR5sxI9pvCY6fQcAuHDrF
0WadV6OmrViCFVewoqLwIylCezj74I7Xueg2mC2DJAToVJDSAcLZ32YOd6o4b1wK
N9YJqYZglC4rNHpFsFGzRZWWYJEbLsA6YMDcPSjoDUG4afXXo8KuDda8k6a4WnXE
47PQLQPW2cu43ZwzXVEgGeMSYikEPSoc8b8Sc07ropIG93A92/Ov6JT3FOoqvuoJ
kMmuWOaT4IIXy9ZzoKbyMGctgAdlW8ZjiXyZwZWVVBJcRLzN5VIyK/4t9fnzJjU3
8w7Ls5ALDf2nY/0bvHm5TwL1jweTWOUAbGSLeisbWzjykp3CdFm7M6GHi4LG+wP/
YR6UzHd8yYKFdtb3BfxjRo9rd0UBm2VhmPgNU+v2LDaoSahamn5vTbIbXl9ZAxIv
RKj1PYcOL9CEXzatMs/ApB553JGXJzQSit1MfR0LpR3T0Mq+DdMMVeZawVdtlv8g
eSUNN8O4eUpr1oiuOOf3iCyFK7mE2txEJZ7AFzuYAPQP6VC7oUt4jCHm8w0qSYDt
XNyCqC0/Z6HXTNX847xbvCUcAwXlf1Bynvzq4ollgWtj0KCTzj80gLijths1Wr1r
/f9x4mqGyhoN67CwR1SrVzkp+vU2hufsSAg2rOGzzWzU98ulf84edGyVZ43JX+7I
FGEb2SvKFIJzRlhJgdM7AzPS2+OkYLGf1dpc0YplGIxGINGtz460Tw8ZBMmvx55N
FUQJHIZcCEOLxmkkSD4QGr1QCjVVbux773YVJv0udQnLMqnA+ENtSBzALdG1io+k
faOe/1+UYpKpoeDwl/JkrSMq3By8cJ9WgySlBrqpQfybyDsZSINWmPTG3hh0+Lue
MHYdfXX0uanWu0E/2Um51Veoltn+MOGzbsYyhgG1G/ptoonHB8KucuSGmT80/tnT
azyPwIGlV5RX7RWDbpO18SrXBp4VQ2ykHRdYdS19jMkaT8EwRUCXWMxLQ6+1iHNO
m7tq877wYCQ0i4T1mT3hgZicR43jbpMtNmhPLaYHhubmdjvFiLXWN/6nfHOUMMp8
2p/Ax3pppLlAQ3ZlmMT2pmK4tZDYxZ+I98Mw51FBPZd6GmRLcYQxBsMGj09JGSQF
ENeUqofxv4uZgatMlCzSYzbipMH0QHxZHpedu+NUuNnqK2pWaWsfzeQCUzt5zfJq
qRasfjS1hR0klvJbc/c6AxVPSrzR9GmsWfhhbu/hybOaj/SwKgxZLqGvHLHDn0FN
VNJO9juBKpK+VQOKzrp/Bpg26duYpvtA1ecpphQmE+I4gk8fBWwMsQajFbukb015
j37nRsVlK/WK87jdSP+hd0lrYWW6IENAYRWSmlx2kcKh6VLHH009lE4edYk0IkOV
OnNad5eTnVLnESHuh34b6XFiH4t6RWEWx6QMgFnxjo13RXesBLSkJ3D3GMJGa58X
05kTaUNfFehNvqbnu+6OFOOsJPKehdi9v5Q2NOgkUrWf9H++mywBSg9aO06B7Hh5
/DJ8zC8POUfSeyxf28/iPkLNan4Thc/V5Hi05WxzJBOfYuv/ohB/zAlgV6NIgL6/
Tec4qMkTxEeRJM5Hv9H4ZJScMa/6WQM+j+iNV1j88faNbtZOuC280vBodn6AC629
QWP/CEWgFRHuHwrDlXBTlEB6AXDGpiq1o72DefGMt0HDdXz2lJXIVySQHeZrIUnr
fl31zgyAnGV/8ND6vZzDWGLuzNxE2d3uVeNO7KQ6Qfka1V7tdlg0/zZwsPGGKv5f
Y2HJqq2Sx+oRs4aM+Vj6ZtMt70yH8OOHvj9GTWjgIVGFI6q7XFCD8ALtbMfzV547
pZ0dr5wKhe1pmarSyQVmMN8Pafmvf8Pu6rrw1YrbYF8ZVi0pdR3CHsEuST/stNjO
w0euGEd9+Xu3sSUvmR/t/GOZseSNF8/l5BsZ6EZHe0fstKrz7FnhC+R3NT9DA0tb
FGha1o06yO/JSKVeyP5ndn0pSSfu0yyq5DMMpWoWwCFemrthKngfSQe+qaZCzEt5
U0mWOwWVHuiMbCUSyDBTOajbw6T8rIM1b3VRPq/k/pBoX/EtWaPlpRyB7gKsk5ln
HjX8zcyCixaIcabnVLL/PnrPzxytpIlfQZ8KXKKtZtsmKo7VzhqEAbZHG59w5gDY
iyofTZD0YE5xWqQnT8ZP6n8mqCyDNMjM04RREEJDjAwvG6mmr4tnRKUybv4cnml6
j5R9dER5nEDT7G3Vhf34gGCN8pLbmVr9oSHLe6F+vEQaHSrIn9/pCqsNlKvUwDQt
nYFx55ab7KzdjPB0WdC+x5haH4npEX86ynPCFZSRxZoJdc7XJ5JLav+Nx5sZAZT0
/F0zD7+S9JR9ub4Fy6/Gp2elClAFO1mHKRS1HPZdj9q9xVh82gbySoCYMA6bgidP
aVtNvThNnpld1ptSDhILVEM80E7nYwX33lH4F5rqH54HEWSpHIyNpYku6qfoxKjo
9apXzUANT5IcCxQE7RrNTO9rjOYk8SV1uavVAP9UNDX2hipF1ZtFF7dA0R4EpFy7
4VbjU5XwosttXP4YfTpghaV7HkhKQmcv/MW9XGjaU54uDSvpNACpxT5iQo1J6TTM
mDLUXuJwa/MqMWR0t0eDJmXnSYNBBFuEkNHHQ10iA/ITHis4Ifax8IKEFZLKlp5p
4eru6HHhaVqAbc+s6AkKypDyS/gqRGwyFWwPqBxpv/ErphUEnV6a0C4vpc6R7Hku
pCp/ABRXZyvKbi5hmu3UGPI83cyC1JPqAGRnE/VED6PKU8JMGG4BTpVaG7KpmvQm
rDnVLMClK0jyJSMrZiB6YxWtx66HqMF0Wcj+7Z0QUIEKPgw5TLkJ0Pq+UDRWVSPK
4ruU7bdCMD226Th7q/qffUi9ODvt3QmZsFQ185G9XCFgR36/xghzHsvLGkd8Tky4
Yvc5Hn+tNk0o+C3wJhQ0NglxHtJqFRNh1C+jzlQNAS0weK/8JIvUg0zgm/8yruP8
Cril6hVy+rqCDAG8rX45hSbNG4Qg9g2PO/a70Xc38xuEG9zn9SURk/OUJavUbf22
/PBo3OIF8Z+CtU6gHobACqQK0NFrNzPxWQOKZ44TQsldovf8eulFAeEKKXpd6Q7q
9hhmb12SJcsOsnhJeO/gQeIoV7mNKv3qTpdvAUJoX+8e6TuSpijFVoQFd5U5FGp8
go8+5yVMuA1ogTNdM7jXOrTG5Mu5HVryZ7WrxHn3uq9mke5sCzerxGeRw3M7wmZ8
EcdU7egEiirRCDQ/UJ9qJ2l9MvJgVebcMzZ0ehX+2dGvDJrKnMiD61BTVBM08l3d
nCtnDJfsOsUXSGsv6s+nYhQBGn2C4S7bkmnrJJVl+ZmTgUQ7JgTJBc3ptlBmkVlW
r9mTKSr+8jD5oiv/RpJ62/SNdGwh51SfiezKUi/bAfPdx3wkiIuQVwC0AjO/wNyj
auzK8GofjCUoRU7mxkGuRZfQSdLajtesd4puUXz/CTESLuccavSWPeyy1abdcQ0O
6aJlcf1/2ya6+hmGaXlRerqoojev0OaMoOOxiX6HqXzu4IA/7BnChtLyk/M6Vw4Z
ioG0/FM5g1o6qt/Jpq3AByO9HPCbgoAr2Wp59bgvrunOXyysVt2Z+MBEKx5uax1Z
Wif5V/ARE4eFH1D0AZT33ZwjNc5pQ7xvI4K7QSV3ZDIQoB1ZD5fMIENJ4F7k0KML
6HbEPOW5Zj3LYHmt+/HlqiLKbn7fN9+/V6ZaTBiVjGAJZc/J0v02H/qSaP79Tpph
HZlL7iRni80C49kIvZclFfVIYZLkXMmmUEbyIANNC088MBkXVeyj7a4iyd9aoP57
8orJQbWskTFX5bJehdPqr0Q2kBzOar9uJaOHbhqfMIxnn8XTP2y37TSD8fTW6wP5
LPlBaHGAePd/FDBhHnVVp1jdjxNnFo3+MwVGgkFYTAloCvrXH+gFjlMdM2A6nkv9
dIXOdNrTpqkRHvE9vwRBBYsQavhZgZkHAdP5dGAXXCRjwxQPE14wucJr5SxIsDr/
RMnAhLFDJ5xGFisKbTuISBhP1RryP5QPrAhTB/T7q16nAAsPatNa51WnVyOZQziG
ryOCUBWc/slz1+I4bKhLTAMJmnX97PIZL+PyXefSqYphpOdKt40+oNjOdFubqYzT
MC3pqoo6YvWmcMzZGbC8c4+frIeHufLWo2MyViJN6rDogcJulA3m3Qne9Au+Exc0
34T7VmwZPCUVRqH2RVLZvkq395lyraWjzQBuYAg8MGupqgB+WqzjnbqoM+oZ6Vul
tZ5OoEVM3aFCNU6msNKshHpBpddT231tCsG+eyjD0TMUoJDNiHngpGR+XRfbs2Ol
DhIMZXF7duLaY6ihxWqeezswhsiT4+3iLa+0xdtHBU12snh0RDiMf/4XO79MC90E
QkW5vddYzkLyJc+CZfLOPptNx2q4sV+V+g1ZRcY2+r+rbZU8FxXyp0cVU291Z+hd
kMNI0AcCG9bDymYHNRPYHnBfF5ekwJTboaQJttStliawMP4JS+7GKirUTb+YxONo
pPxkREaeszGKG9Sqk91hu1DV7gI3+cQGJZ6Un8xBTw91TZXgjXooOvakenBtY+r5
QqcBbHR9biqc6QOjNRFaXtmbQ7ICGS4OUCvHkpJdFphQFtxad2A/mPNQP/2Nf1bo
YMMD+rt8W69JZ4iFtBThGLmwAjws42cKVdAAAxyYesJenFhKxORUU/9wDtmLhiYl
1ogDXA8ea7F06KRLzO55dcImF8eCRKnSaHq/iTmLcmSgt8lta14sbFpWR4JWlBjC
h/+kPTs6i2nWScW9M5WJV94W5sJOzW9AaGwYSV15qTpkdWm7dP+peYrfPGGbrB6S
tAsh7Yn5lWS7AFCl7kQZ83jtadu2irnumXSH4tkZ5rBDIW9ATTWvD2NGSHFpKicd
Oml91UR5El7P5jWXSTNlEaRbSboypeAFu2zt57rEFmRPAqMWrhDvQ9jeYmJ1of/m
IIM1fJLCFjdpoJuzIHNQ5JlGW+7d04wTtmC+/0m9WZMtKqe1oTv5oiHOin9Po4VF
STSv4JJy8I7Kdk5bhuDz+sy2y6RXDoq+cWnuuOe9k9253wBqLXlH/KlDWUo32ENp
jhI9Ifm2GbI/YCAlIBrZZo/mkfqkwYkv7aC0iwjBB92TwNv9RPBbyAgYg+AxiDI5
5F4lHeKrKNKFIuozm4bZnrdY8pNX3wCXGTLj8GNbXGa9KPw1iyqHlqUL5n97qOBf
9O9vjnYsNQfXamUHl7PnrqnxTIFSid4Qt91Gbel57BK9nA/Xj9LHwt/wr1KNkWoQ
1rQi5ekffQnJqZ6chp5FFrOBDNGfdp4EOFM+yqbTlc1pjWVxB+ZsF5GlBIG3Ufwp
l8b5eYxLUVZpCIsbkyVWp/sUNrwz7lPsF5Ut4jEDq4m+dDrDK9WdKoiWyc+4vS9Q
3l+8C726N96IoivoTFWhkEOUjNL8torMI6+DAWtXN3krVeeH6GBR2BX6VWiezxE3
+AbUNOGni473xi0AfILwvVV7YqFwkb0MWo6tDx2pWI8uTvCHzSdytLptd/dV04i4
sELzeobJpItm0gSxydL7S/gWUgBmwSYYM/qkkMlu+eK/xIIl2m1NrjnoPUzt4tNS
r8aebwMNZvI1xqdAnwUtWXPncYrst31PK6XJeu1nOVmCLbP5mCVD9XlQgcQXDjeV
rS7pE7MCW8qrdKA5pS0B+ixk0P9q0PL4bdeK/XspaBINAjWRhv/XIzeRZ+goG+o6
orxzeNQaUlKCjKwf7WLbS+sqclt6Y2Dsm0OKwrDoY6bURy9hHmsBuQPEagm8SRKF
0tEr1nA+Cqo9bApdZpJeHS9nXFk9UCWGsSXsRd7YdhQManA5ssltSdijjSiYGxwq
2BeZpMY19g9EhwFyui2LYjHyCPypO6mrMGzw2TOBcqf3qce4ZV2C8cTDnUr3nZWZ
p1CrdQ+xh8KNA97Lef21YvMOU5d2SdF8bCZis8qyiTPWsFvR6q05o0e1sgKhh1In
vv2ncB2/enfTzQwKKHp80IQ1aaalRM6a29hyGf8eTipdPGeKmkih8cZ3hoegtj0v
y9EHaxQQpr/sfP/9N8lGB+HnpHgl+m0fWIygTerYhT1yi4VB1DO1+hg8JzeTtgIk
9OxfbUAmBePx26L6yAlXTdzzEU4o1aM7hMdhqCJu3UpUuHdwJu9XGItWjB1ZdTHZ
iz6CumQ3Y3n1bP71gGuQCfehzbL5ZfPJn0ttR7Xv1vo8jMUv38kDOvTCNrrfo+kA
dIOCfzCAA9knU31RAoXVamv6pWjKaQMNB7aUNpH9Ky32m1eDzzsnL08mCPdmWPKr
ELMolt/O2pEA12iWhukSg/vBJcMq3kbmCSC9BpbTQcEdfqYG7EXLcJ1nGBrPMtQY
NN9v+DymhXUVo1dpZm11X8iLWbVvCbTC0xwYQE0/om0Z1hrR4XsqJc5YgwDBFbub
ZYfNNYdcAwQHL7UiQO7X6KTY+AmmuW5M7hC7K88SzmICcIuAGD1Er0Tp28PyIsT0
IQ33T/5ogTanGqPF/20X5KRJb0ijA4ICGxkreGmHWHEcYbPgTr9FOn9VlfdM1ErR
V6719xVIqSCfdjIvZDR8Vtt13vGvYOZqEuZTeCEi0F+p/K5fcUwWnuvEOhpVoEqS
FskxHxubxAoAo9U1Rvv3UQeqfErDzeRSE1J7cp8KDfjPVfMidTOXWE7W3TJz763+
JsVe3BNHfOKo/Q9WM0J3JWw6G0H2ZFZDyGEA45whIbbxgexkddggRiFa7/a/dndC
fnPXgmZSjsWzAtslXaJ2XDoJ8VIEJqqKOXx49AcxpZbqXdmWuWdUTBx7Asg9OEx7
m/pBT57T8cThSMLbC95s04knCI8BrD1h6l93+rv1AZeeYreX/Pfwle1QOjWVIfuu
2OUZ28TXe67aWv4dTBru9ydewODUY587mVCm2n2uWx9h80pq3rJAPf1bl0xATc3U
llPjxf5kVr6hHf1rzQyDliGPpTRRjHG2eBxZYEVN5Z8xa3Oy3DQlYh9bZpyRb8if
NF/rqipqalR1vSNMtkLXftWJhXpXxxYfddP/kh6EljmaOOfIRSnc3gGne4BaWQQF
25nBt+zoMe5rjiEfDEApMxaVgnaBDDTySs4yhyfaRGXckVh/AOjykHufpw3rqahF
WlVsIsJWE4F2+KNMy2g7U6FXlWGPALKQcLDzB6QZZ6jcZ42Ww53NoIGgNFLpmMS+
vI/CqE0OiIq48MdnnGCyilWiZ/dGSOqbIdWvGSxh7Y8k75lY7eA6KtMVOR9dSqbV
PcSzW6S1IrUAenlyAAzX6JNocXWuEjCimOi2fRs464eheTm3U29k6U7Pi3lsw/Gc
ta+zQgsfVrzhwkNDWbgSpjMiY2JxmZU6BLBTCOG905uVlaTD3jmecoPpSthtgbMc
Q06FRA8LNbzvsNw3VGbzvzpnpQLcqQaSSPjNtLbTk4/I5t2HIm/KcaTh+rhnbJBK
qViL+Pa6Ej9VJ0uof1GVqFyjdXcoVUYMjQebFQQqA/l52cMFAJbU6cPpDTHhFLDK
9ShKi6PJqGxF/wXEvQwfJmlmJZbdFRqRwwwcAmRCCxYx2lUfPQ+h0abprIDt4eR0
8i6r4vo9YcIQl+WcBxEf8RHbvjU/378Wz9YnsQRQn9q7fhuSM7THEGjkmjRzHNfZ
3Z/85iRoMjvggodmD53L2WAU55/JyVOM/AAXEPYCvQe7o4Fh25MjxNeaSKiJLY9g
OJyJpL7HHblykcB1VJA8/OtY3qbeqI27qBpJ0hKGoWGMxeGgD/pD4HSvBH2Dn752
fUmNY8MMunPqemEXnpOPAPAorOVdre2sdHbW6bG6aW+q9LTe7ozT8zFU/2ao0w3c
ktBD3wTJkPLFVhUME0Tle7w8AKD7LuIlwehpP4pHkb8R/61XpEZfv+BvCZ5dy3Od
NjfpbEWtegBASgKJUQcbhJAXOYJwUY4YZJi5GUvoITNLue3+Pr0M6mthUT/MdpkI
KbX6eG+FAO/hW/d/EQRUYd+u1rlBodPcyXASZRMl3M1e7hnpiaY3pU+hD1G5JpOi
5PxubIsxWgwRzZpHZGiB1Beb/O+K9zOdu1fkVhHwpF0HiKuxlrCE2rHyBYbtztlW
uirTEicMLHZyNLtTf+a975niupfrvQzIy9EoUJLTS9MorZiY0i+mBf4ScPfHpEFn
BozDJRHVw3elasxKj6XM9hWeiUIOGwFp4pjTzVEB2TjUaeZoah43nGuCB6YrHZrm
jAeneb6fQYtMTyYtava50Lezm/WKNzXwZA4fWP68bVk8K2HAeMpuYHGcQlzXi4GN
5xf3Zjs8GqYiXjkioL6CYU6OWow+7EvrfF/qLiaiR3Z3YBO54CPmfnmvrK7ff3m/
twdIh6g3pF2eAWscABzaU/0sJ/In0jMxnXuBuYQwLLvttp+L2o6/hQ1izZU5QoxM
lmlkV2VPRt0NAQPCtmLU9nBpZq4KbUSoOKYsTVT9tyqyF7gDnQ1hVVCe2vh8pBOO
RrnzgdZG7hiU6cV8KUm0dYItqwUcKl84LN6xKfsX8huuJUmMng4nhHnICdFIU0CU
ru/kikWdfeHid6miSfmXAW8ys7eYBnxTXsTTV8apvA4JChmGIrletUgBCx5XsFsz
PGl6hmRhzPpKkcpse7d01qKxpgqs/ec8FTg68x9ffUFseFDoaIfk2HgIQ1x9RYkr
d5111NNfErYMFGVaHhjuEWN8TH3ttFs2WesOL1XGd198mT5hmX6QSwkKPpdrbvE4
PfAHpk0KDP5JasbCts5K2Zz1IZnMRg3rLEcxJzQSM5xkuAvFY5+ztjhlwF+8cc9e
V+J/e323Z3NqNIrA5ddOZM0PWQN6RojSsfpo5KPu5wZADOfJ8v1ai4DIPs7CbCqd
DdzudBwSIQE/1XYiDP29e3Uha8al6PWXAz7xco04ASBir+sNDjPB/Fo9D1Xk0Qqs
q2ISz7nU50pc8Y4AVsfjaKV8ZcJtZnJTbyK3c1PKGGgi2mjV1TM0ywYkZWfWzrI1
mErLGk7DxH2GWT77S+8I/Tc+7B/IRYLKfCBP3raGyGqfSAtRWzV9w3EpwtvunTKh
TqdP/qYD59UShg3uNm6eEDEBKdSVkjfGPiE7UsDFDE/oPikn+1a3SLy6IMYrCz1n
yD5CG4ahoxR/9BTc6cJC6wA/hidZu7kwYlOZLHq2AvibXAaapibH0NV6mT5H9tTx
I9HWhZnk7BjsEBzejzwL/MqQCrUu2Px/MOWbdVC3dIduLBRkoISiptS28OiGd3oe
VijLlUEC/3yUjiaeFmVrWG1gYzKT8kP9IOqLNXbV+RyhrEVLWfjU2p08fKdDGsZ2
AZ0C86SFZXA2K8+uLLPdgwgj5yevLu/qBbkxXkoZtI/I2LvQfXLav08dyftwzCnj
V1w+9XiUamTqecQwqhuy3uVI++8gCBsHCQyKTQQp9WcvZqAcVJNqXXNVi05xB7fE
nzf4966umiez6MzPsnUY4lyAafF2bWFCXjEZR8FxmaAV30So4M7M+rnX11js4uoa
RP0xQlNtHBc706f448yAmg1QvwVICn7ag0bT1M51z4Iq9zDnhqCVRPz6+kp01jXJ
tZ6iv1zLBHX9gqqg4Sa33d+r5zwHZ0tRptxzEHGtGW5oeeHUqhsHe9cym37txwmZ
f7Te7cHRB7Gm/4OwwuYVwKWSho44BiM6RgJURQ6G7I1xBUYx2t+2IWG6O4q4LjEn
IR6zR5JSbwEQ0lcsegc5lw1vTsfRnL+NQ/Kk58wmDonhqWNPkagOhEI6Y903slut
EgBQuOnissiFKivlfCGC7mK+5CJs09Pssf14NfP6WGzopG/Xu8SdwfOhzePOtuBy
6zAB8ammnHo+baK+Rl7hyBCge/7BDy8PdCX7WW7EWNjgVsiJwiGnjVjm6X1XW2gv
5IUkyIwTsIWbJmWX6ITI38l4s6YUr3qRFKHouFyoWy9sQRm9CmFHCzuGFuQYHM0o
ZIvlHPD/RiZklzJSQhxtVWlStIquRUQeP3lxblyTYHld/qvciwSJxKXgycDsPDAr
EaS6zGVrV4jg9g9Q/ZighX3AI32ItA0kL79en1PBWkueAQb9KPijX/4Yzm5rTtZL
5sJBZeEjDeLJvKz3ujg6o2iDCjhLWrz4NYNtTEGLnlaTsEa6iewj47PAjPEJQC9p
eVoXLLqA0sS34R/4tQVjATBce3b/1ocJ6ye9rx/JEMDUQAwXcSWxAw5njtAZ6vMB
dvpCg5xppKvQ0hj/UpxUlWeEyA6l7JzzniD6Ejjyf2sb3q2LbHe+WXRfe+MV/TRr
yq7molloDavoGbwhn4qLOEVEfnj8g9qxOgGVk77T4A04xmhiiSfLH5bDDLVgPmz9
UzZgqs9hsDXVzxGPjDu17UtQa9yIGSfD8jm8w5vHrnVlWwpTdfgDa7GO7aMiVuOu
THhB2PHgTHqvd2V1/aWlVnN0ha9ZiK2BXPJfw3uehLKF2xGcKjsn+EkIdn2Rspwc
wX9f/mn5z8YsOna1pAaTmEqOve6mG1j1gkTBxpd8QRxcPq4s0dzRmQNdndOtJcL4
S8FEgrRO9LTDb4njYJINtsY2tuMZE6a6WzOsZUDhZ2naKXZHduuDpdwvdjsvGu1V
17mK7/+6Y+fa6cyJXyFofWnFOoQoSOkRq/uZlhRLog7q9pnFOZA80A8XqfesCXZn
Q8IaQqk9h3vrvaQh5eCvnHI3YOXAukpWHfqKM5IgbQRmF7+YoY1WZgQLtQxkW2gJ
5exWVPEsuMvsm+ePWFdfXmlNyhA23O12COpEh2SqlgZoVgQa4H4rGbtpUOoq2a6P
VpN1k3N9WRJXLgJCn425nwD2gz436NA/0l9+/aDAqZu3t3Xg0hopIPTRq97GEdJM
usTwA4a6bxCsPOBmUHs2BqW2ou+Xcq2JubTckPfwqgT3mzpFf86pvUeRvvyFO3Fj
a/iHJj62Bp5PSDxVNMfTBfgLPeyY4frUomczIlUJiGPxmhiUzaPe3/O5DmW5GV7Q
v65OVeWXgZX6rFSDXNqzUbQoM1UxrAaM34psPOt4Vg4hH0psgJigrnteM+yry8YW
A383qMapPSjURWQfmCBbW7ztHQgCQnccFrNAL2gYCIrOsh4utuHaYdhCAug/upJK
+jANQ3KGlQmvOL4pcYoE6Ci+lvxdpGzEaG769Exj2c59bAfT2FggVxdGcXeqmauZ
9fDWoSvwLze5zYbT9fpegBc0HhI5nrxEGc2N1Bo2CeZVwOT/kG1BxSHpfdMcokaj
QfyhPoyl8XwaTLR8rpC1izRK4ObdufQj6wdpOApscEdoz2Eif2wuPHHD9xpCXFps
bLYyctJb4LUlTCeaNkWcG2JNWtuuEwDe1w6ODZyRYCzxVg1ft4KIGf1VrGrxjgex
HmH4mTjm2o4bgBogF38Gg6Bv2mnMYIRXK2LDc8XP40iiH8oRQKysouQCPi+8D4eR
EnzyaUTI248LZFI292HrYVNKY/zVFsXf5G/ozaheNRyF8PNfyJlnxOLKh3hyZPzx
Zd+RoKaCHYDATH5M/mI19li/xySuKlbrxgG3rxisWynnCMcgr055LjQepSYDDK8s
kIRvxOgn86MjYh22AHqDY22so320w5Z6IOH1HMpeeFw/hh7sRObUGK1qK+eIIaSe
5Gu7MF7dO6osbtVG49PBTT+HH5nW/6lWCJAoydYug1IBEkdB5VoRBBZDs2KJGEkO
/ibvU99tiwbtzh0Xno4thDaQAj56K0Cw5+mymbZyYyU+OhF18HHzQyaGJC/4bMjJ
OHC3D8iEIjIzZPLK9Sf61DwfC75zClDh1q6a3SupHdrndvwhBvnf9Mlko9QgjLnz
X/NF8sSXcAYLpmqD19RiYSNn189coJj3cEYsMnc58Ns+41LjsFvQqqnk1SJi9HD1
QQkhhmileP9zpgS6o7v0zwuL4BGrPVRym2bHVn9B1BgeRWDv4jF6m3NjL5gwe/8l
WAuLIwAoBqCCL/qMJySLAuWDzf9EpFu0XGkEAazD8oxYJ+j3gxJ/B1n0dSE9qnDX
2qu2P0BtEJKyps/PE8e+ARm/3YpjZTEei7CqCikIGJw+5VgXmD06u22I1DBKx52T
a+KJBdUpal6SlYHh98lxVr6ECdF50jK5FPDue7lZgK7h8hlgCkXZAoZ495QhAa3K
Y3W+LeI/h5AwFLwY7bP4B90OvuWtVuYt7R4/B0HYoHc3OzgtA4EBeJ3MLAAMVicq
cj6LaXesBHvzUFWVZ/JS/RBr6bRPgEi03ZAStThxk5DGaqGE5Y6JyoUsVW8em7FZ
JIeSLbEex5g28C/3ccWL32dB1sapUO6e4BTIeSEbrpmb6/xw3QWyGe41ufJUR176
aBSgBkvH9VHezsw7MOVCLuAKYAWyu8dYRSTyPI3pCYTQUmilcEbVyUVgMPvkWuHm
vszW7sdQ6OZafatoO4Rhdci3N9ltYVxDs6eOoAG1vVVP+tvpVCd6W9UaBgBLf98J
8E09firFtUj9AgKFaoPMq8f9svHdCURAyl1fZH5mphvb5zT8w0ni6zxq9tn3kw/n
B2VGAEUNfKd685VE+d4J9HgN5FZXh9MCu0gascQ3KXRX8cNI8OtZ4clcnG4ATQfN
T/nc16YEhhhUW1rdxKvUkW29Fcy8AhnT/4ul2aq59XGrk8wze9V6a7g+ISPIpE1I
XswlFHo5XwApLM32PywVh/F6pVgl/ab9yEdMwK5ARshH3af6w4RHkl6tjh85QZmp
LJLJJTJAudGqDdaQgwkhovL51fSDtVfSR12x7mV3YgtKmZa/GZrF4vsoKFfy6I8V
P++B+CkeBaV/yyEbHhcwFWnwcPQ3SQZiBjQwf5yln947M6Pq8TOwFhhEDh3XFf9h
fEXng7yIA4AizAUh20a4SL0TB6SEIqOLZDCvXXQi6nJPFwDGKT28zM6l/eSAKoLI
fWom5tDiwu6H9j71K4PWsD1U1pGhl7E3F7/P/kdX1yrUR8oMyjZISLyp7yElDCAc
0oFxPs3fn5zK2m+jfUQrZ2vEVDiIQ4SW86a3Ou/74IwO/mjpvqtmu9faPqbbgn4B
EINF7lZPgOqcvianbna/hAK+8b4EMiYGMji9yxJPkCQuMkM9lAihYdvesE1g9Z+a
PTG8LUVk+k2ysGIrr4WIx1GInYM1Pm/EwaLa/M0uwvoZiG2VJiwdcwITsqyMt3/G
1J72DWp9jlaTQ4sC3tpu/S9kxIe7QrrilJ4xB6DCcYZtSr1fdNcQnWeC0Jsqb3R6
lXbG4Z0JsrwFp+tcx8RR2+BhTzAt2s2Jw6BNOdopo93XXPWlT/5ExHYYYMNt/zVn
g9JERcwyKz4KvyTAdWMjUtK2iXgs3aKfHrpOjhX/QYK6BNeoza1iMwlyC0hZFDaS
Bktik1AADj7UfAIWIfImQLfEUZBSFoVOZN2N/zVZA+aOEpzhCl4AYzMF5phjdiMd
b5CaAtfmJFt/yWz5WnpJJ3RUsuj+W+EQqK9X7E4D+dCfRPlN/Rt1l0zr8VTOe3nR
wcyFB8FK0eFpfpfFOBLJZ5pHFoQ3ZvIgmAwLPh5mX7IU/hp0WBfXuS7Dm7A6YxKf
6kBrp8Hv0CIUu9bJmew46Q4Eil9z3vlIW58U/TlMooZdsUkR9f1PspH6yig9s8fV
+9kKwE3MQfULZFLmbVyr+yX6x++C+bowjZWG5IPExMI5g/TnTfFWMet7pGJiwBjx
nLZyj6nKehBeqTUjoptkDT9snjbpHlQNi2/yLjY/pGnKLF6gEB18iFS0xiqRJLlq
+JUystaONIUm9m8o6D4ejxEETTQTPqd3oXi9jriYxeyNPiSuDVrpUMygB4JMj981
7GMO6yRj5oaCJxo3282z+d9soWjo7PAYVSchxDz4eIYj3aQyJk057qM4OyBu5v6N
JTivNhrtiFoBZwXQHEPlIFmXaT84JPnrR1VKTEv675xuyfs5mph4A2wh9Aj8zB9Y
2H0g/y+Ly+MTu+0jVQKxPNyQsbumwFMUlddxj+rgWiwu6x3JRWcnGzEfFpP7Kj0b
cCGNFLpZBzOOZCgYmBX31lFrUo4W6BuAxFqCAS3rUlPvC0xgiXGl/L7mmNf/6qa0
ruHaCXuHlwqJ9UOZoyMjSNLPoGwjlxltiWeoHt3ZnkZhNbXuT6ozp6h+E6uhfRjF
6O7cwP0JpuzEqBHV5RcNFqrt5irtdfdwXrCRnketne4g+4TRao96v8+5abHaSGpx
ur9u3GVo4x1gtt4aIOIdOQ1WWRtr6TW61paw4So82AQwNdKDSQI6TuxNpcoN0wj/
ve7i12rFYZKARjANB6R9zLNtFDJHVkyHn1BBzdYbZCefKhIyWF+uvS1d3y0a/gsl
HPgV2r9NidA0PRlgmVZGXzvI6nZTUqsPCfZNc/Z4Uhc/RYXuTxLKkv8rWQcCPgK1
+Bgbu2dfa+FnFl2wSGU/MfUVJoVCxycZ8xRwsNN5ET7vxSEIPyBT8GwlYXM0jvob
oEjjzkAIgHX34YeBIS146qAUVIqkedYH1/T9HDWtUKgn2ogmErd8sZQ19J78ybCG
ZIxPoQHEKZdzU7q3L0DlndkQ7qo5EAFs1jF3ptm7mjBHPdKgK10cFe/WdXW6M2lD
uqa6n6hbYo1i+erLRCGV5Rbf/4Z7loGrO2AkeYdLlsxXWQLU2Tz6H2G6muFNNUcA
bABVOi7DhwtN89Lvyfmg32IrMAudLx+ID0ALHO7pqKk1C7ju0TigiTOuXf9BkRtj
Bx/kebYcCD9L1ie5qIzZGCcLrCA4M6Qiw1ZV01owEmiPj/q5KDWT0H7NtnzmLSon
RvneONvcmWKPDjf3GRikvSt77/WLm/PnEwimxr1jCp0b2YMAwYR+C2ObCi2d2CsH
UO0MWO/z5m3F99/nHog1yqTBrIFwcftniI1ZjQHoHZevA8ugtOoNdLe9RsE7B9GH
/2IS9MXXOVxnLBmchphNc8HDXpYQ0CbHLeScTi73A5LirUbtO8hyxkOdcZeWtjgc
DFs8VHxsY4rkWf0iYS0F7lUrxnRJRyrweV9NckSUgkTjl/twFZfFWfbvvuVHO7xV
f/xUX+5CJWQd5KEWFBmYZd+CMzHQkYT19qCbKm4RLO1ZePJm3Z6gMYfKA0lwpeuz
FjCJ8zAJBq9clr6oooJV6SdbNxIYkiuBO7j16Go3GkEifP9cHk1JEw2/J9Sj1nPW
hmYvOpndFtnq3SK0pWoef81v+cdNf6QWrVFRTjqCuL3ErtGQqbqeb76m5fe56Hem
43zgB9goYBrioHWP0iWe4amP9NGQ82NJvAi/gDKjsQI/s8c1CPccVoZMgx13h0PY
grsHLf6ivuszZ5BT0eh/InKcbY0smxkyHWHQofABuh8JE713+6MckFvgzLB4y/is
UMIKuLg8wTLH2a5tur+GrviatZ9KY484DgjL+jMOu3RfW82kGIFt/tDSI//Nguw4
KY7PttPlWeNXUZ/HYSh3EkES8DP2UNaHrM93qhnJHY0HB4k/d8Ukc3tsWsMvxqD+
2NwBXfQI/L2wmRxhfquoNtyyoGhdc8Ek+lXwc10EXH2iESAXVHnDKwyXMW2+1VB/
6IHFUm6gVh9bOyDMDL7fkeel1mVgLQyBul74yjEsxKKgAVPoVLleMXs6u7/tm/i3
QWtzX0NxJ4ZWB4NeBWfJB2D21w4WLCpqJVRDzupTZVkX9Jtdhz9ntudi4mEjT7Ea
zQW5nQQjxEN7eVtLUNSltPN747GDHe4KfWJNuXqMM5zBTg0oBiP8GXg/SiSLh9ol
jyumZLLbqXxOOY6IWgU+03cvShy0fMa3IEIjhNmMt8gHLz4aFOuLF4CvD8Dw18G1
0Qw3/EyFyrJ0E5YlGv/yMvJl24Qo/j/Ew7daPGEBpvrszCeVRdkw4Kijkghp8vyX
eqQufTzI7KUt5Jbl1d0pulgU+4N8X7V+HT2d+RvEh4DD2Q/xgz5tIipT0G+4R8wK
QXqIn0Kzg8VQOoesV2XVR2otP7Ngp9Yc/nZX7wqYolGscawRolqLb0+XZ8L/0RPw
9NV2EYjD/TMzb5RwW5KcjYXntp0r8ifYP2t7rUQxZw2ni7XtIk0RUsj9mxxiIIo3
W9nst5WDL/Gst6linzIDIJa1k9RysjqOS6XGWSbt29W8VRp2xD2I95Fxg5+qJHp9
UbjS2R0OEkX/Fz8IvTg3ve6nA+vR2dBSJ5WrhmAd2MmmQ8zcrdXgxQc01C/Ty4ia
FQm2ZfRgxWpzIi0f7SrQbea1wd55J+sgTfXPYdQ1cF7vpOMYE56z6kPKZkkLfjkY
2eTTVsPl7yT3l/DHN+h/NscIzU+PR9rzwBk+xVaClaYwPCBj4JUIwkweJl7sm2/Y
iJpImuCta1nz8agoRLoS6Ong7aYqxhaO7kJuzd5HsCOMdINiCxoO+px7RpzjOEAK
hFL3YEIpJMPvPJmQjOlb0ezt5TfuxNykpQ0BNuPkQUY76MnG6yMSSdKr8bt5+b9x
qKG3lSOECZcNWMs8iyo6eYtWjjHyZPD2Ax7SvO3qcQWqeS6f6jfeKZTrTPX9WPKJ
5UqJgzfqWVUbqPJoj7JcyBsxZDh6jZwgwR2PERRtyWIzLx4IRxeyR9FbguHmpHSn
dxXv8v345y4C/qAMRDjf6R1K4uGXc8Pip+FKzkaKRfwCW5FICpyR25f/aHm/G+U5
Vrt9UjgZ1VYs9T+EKQAi0lOYdx8m8n5439ZXOK+P3sP6f7KgVlJ0oNRV7gX90PbS
kUuTLnLoA888hxpRhpKtWvr2Fy/VN7BmJm6TZIJCUq3ONJs0q5A6RxqTOuL7i8ML
H+Z0g0jS5z6GfByCa9SDWLXwjiuIWgIyCLfLHPYrq3frBMUfTAT68Tzp4AuyC0C6
XNXddWmEYPLXa4nHq3P46oeG4pBIqaiWD0KG5q+sn6Winxi5sMFMqxxGGDG+2fpA
lspUfA5cipnQsr0YaksLTHweE46OwXTUlMVP1o5ZJ7b+f0agcMq+Hv/Ra4FOlsTx
HkAGcAUtx5tobd0jgSuyKYeiXjstquYqTw3oWIp+f228GUeWORXTHvk0nBjo6pbs
VET9BeOnekb+LFcyFjxkGjYtn0vPgu9H3cx/Nuc3loM+KXbN0wr2GkiMjRXXApSp
4GJg4ZlfPR+9ydMtZVQKZWk/s8CPtG99u5RTfmgkPCUIa0sJnbkmSSzAgTrlcd+x
snEBH6r11n1C1prwA/gF3oQAPmcDMZTRZtdjD/SgZek2VVOkV3+Vyoa/vx7Yejca
FZfOg/LWPk5vztI8xqMiSqhCvj2AkLTk/3f/y3gkvFCS5a6nj4m3IyU+i4CiqTTI
J8CjQg7A/Otdd6mHqvf9myQZK1wFLe3wU2mTdxMOZ34hht3KzuVERgbOQpPtSYEr
NQZ48TJeAiZ+X4f0drnlWte5kCtAPhOAPtuhX7jt5HsEu4SqWw6LwYgMM/dY1SJI
drCXOdCG5NTEAUqUj53xCKdfHf/0uUDLu7MhHIZbWmmKQXJdgVDILIoW+VUS8BAe
gXT2sLg0N5FrkeC7J2eVn6qLlQmfans5aXdH84QpOfutuhf5wpNhYyKjuf9SKd1W
Rm6SFyueEYttIk/TnEJ6wyuCk9EP+oKUFWVNmIiKLlvvow1g+m+fTd4L+Riq4mw5
MgXpM/2RNQijVvxbtkuErvIvMwlt9VopfVZEfraU33VYr7RbLrcJikHkjXdrInc3
5r1KJLNh2GkrIwl8lv3WgpmpbMz8FrkpDAxTJEeiNI4Y/rL7Xl2cHyZ1lJrhXtAT
bxvVHxZ08hv59N114EPlqmnYnianuBRpvBCQ6FxugVgtjbuNWhAfC+ZtDlSlqHJY
lbKN/qMpOdWi3G/G6GpQBN6za66AHTygec7BVqircll1ThjCenGosQKtTjmekZvb
kIa8nUbc7nZ71BAb/uMG473ujp0UPpresBZ2NAUteDECSlXMrPwjvCor/KxgzmxT
SfDQL4USKE7/D0tZPJzm3cbJ4f0SV5yHF4jr8ieAUEuranYoluo2EjVAjxFVrfAH
c4HGYPkmZQi66kj3YV6EbeQm06cZeoMC5MUVO37Ku62VN7IS2Zoxe0S2Y6DLBLt7
nzbdZKzsXr43YustP+5XnBMpgCm09QH65DlHdOBodWt5YAXmDIqLEtT8Mt3p4jHh
2QiPT0nsyjlqZITWG84GsSFp+wrA9Ywpi/HxdLd1HXYR2slRT7MurqjvMTJE9fAV
DltwKDZt/NlDngBI/D8F7o9EV9G3aabidYsxAe5QU1kglWin4E/34p5Z4YQ7AvHq
G2dgX1E+V6fYaPVXIhIqHWci3MVk0iZxJrSMdKgGo5Q5H0yz7o1+sBnZsS/VkBhF
odnbxvLESSLpx4VaregyCJMb1BGkWlEQqKW8wRiMDjy6er7Qw8docz5q93b0IQ+u
AZVnv9yUOwhGmuYw676n3bXdE2NITkW8JNdbcK2pSbSEl6fhEPdvaAOvz2pVWtrG
WLorhPHfddvqr/nuob+wCCnaR9eifHYaOFjqq4VDHpNneZPDzf+1lScCuDM3EsjB
O9brtlRLxzJX5SO3sLEtzUi20NoCMQgDnrdXztZ2WgqNGqadR8cLhbzPBAC2ug+t
oUbcWkwvza+WH9awpqK01c72lAKwcZlohpJiN9xXXbJ3O24+06cMnVyhcmNVvivu
hQOBPBjl9rMkdytH6mqYcjrhLFxUlq5FkauZZISkW2bRDsAr+YN9IJJuJoujce7H
sQvRZcfnytv5OZcZXXzA1UCX7D09pJB6jx5+s6i0PEphklLScSUVmIf5zz4KiKJc
eOD3IlS8qMThwbSiyO3clTyS0aVxZ5pqzvVWm+zs5sm4YobgyAil/q57YCidgCuy
3nSLdybqgitPMkj5kDxJq/sFsQ+VZM7J6VPfr1SGzgBLhEfU7UD1jEtV0ge6uJbg
JB/nuwmLkuHexECGeKK1Mj/vNQAH+GVQP0BBRxbi5t1TxHKo8x9LhPx4QsJWRLFW
jTq2SzIhvZRH+ViqEeI7amUkjFfJ30adNDg0UpUcrlbPuUQUUQrPM/4SfDPxrnKA
TEzZ4Bjv+eI89KYOMQnwyEjRbvX88FxMMAluhCBhCKYLFSNL9FVK3P3AdeES8Lpp
xoqbP/E5xp4CxOe3CG6ybkFdGfo8MMVFqBMgEVuPtE04nU6OwQO3NNyfHgTviisY
YGbMhHpxiiwjIfbGxzXODZT7rMO1ElSnCcS50UnIw+9s+79q/XWT7f4V+X7BUIqH
wkyfJQ0lb/3gbO2exoHguYQOMJ7szS6B8PheW28kYL7zCH6o4CFFTSY9a6NDLiL2
A+YFwRhuc7a0UqJXxkHRiqO07H8/yxG0nWv10uIQuG6TJ94pgH33USwG+DovNFey
uRnsdt0alE8Pp45q8rIDLStXlNd+pZlTWNP8ckZg+JCNLmxP2EHF2WIXXEzPZgcA
C19EfvBAlihz1Iit0X57TYIueFrwy/JD0Q3XYelCjYSks31TvrOPbkDsKnGm7Fge
ychFPboIQB1e7qM3Yxug+tnyM1WMiXe5J0iyAPrCfsBkiFOhha3oj1d09EoveyhE
0764LT/4I9mVUz5kHqr/WxrcF+3VaDQ/18ExIn5xfpjAlc51/CeD6GVq1wdrXsgG
D/VSeTDaaYSKHplpe6rH6HWxOGvxbgVDtAw1fM0rHTajKSgoOyPjlc/ePLN+Etin
ENFzWYpLdp22MeWVuW7Ypmt/xLUhmILJR0SgKdqEL00ZWedu3IZP9pQFUD5CQ1LY
zB93SoYXzGBWvUkvFvpU9W6qKuoxO8hs7T2Xrk7lBeaMH0nGPwMiD9VpF81jOEln
tlkojyAt3Ja/egGA34xnihFz1VZuwGwr6PefP/cSfl8bM3csolaLjy2vVe8YN7jq
MRj+2mex17b4BUt5Qg2dlTfBcb94ubq2LOYmvjjBWokC5CagZxbyhpK1fzoiqN17
uom1UMCu59a6nbXq+6obuKpjZuQ/Q7CzjfNe4P1suN/KwyAwKND/8+lsItXzcVNo
03hNWTix8Ga9/fk+gLw42sveJBrYxCpQXPa6Y0Qj1TjVOPyLpmebG1OVVkhXH1bl
AUJm6XW8RwCcXoUoWTQESTjb+N60eAHiRzmFAzCzgiRNg8wtKFbgQlMT5ZZRzcGX
6TKXBytyZDb3s5HKHKSS3MJZZHdzbTuUHA2RyfZY/lN1MZsasHhLqxJjyZz8vPqe
bC8zJkoHFaVp1LKKISwMOhhv9LRz8udTIYON/m1jEUzfX9owhDGpE8FI8V4PQX4G
pi+k+AKdKYyOQrti0IL3pIBbbJBX9rjYLBzXTEwrvfYA/umh1FYFqjXq27+I4GE6
G2HPPMKfwfuZi0UoefPE95+LmcGQspUMfgGBXipasghOzI1RtCpheBXi+GDNF9ue
9ysDKRLryN1cmkxVeVlgS3UU5ywOpA62FxhcAGal5sEvYpKwFyo7nVVtG0h4W1XZ
FZvEy0UhUn6r6z5WEuH2VcD8XKqfqHdIOa+MyD9VFZZjBzYzKzTPvKPMx2Q04HIy
A5ByQMXMyo1EPYJNmDNNOOmvVIyYNMJZJeUey3yiuo0D1prpDpYGotCx12COK3Dg
4Qw0/x11o6uENtnTsIqSwRyAUee4mLkM11CcSvIBHVZpwYDYB8wz1oA+K93TzvWI
RcvJIRdayZlU4nqIWRWFdc6Q+vQPYz0sUwKqpy/RDMzrwQnKa84laTXY1deiHT0F
SknMcDFE8XAtKmSSi+7IJ3A+O5998eFa1mJKLgpCdPBEuuB9KdGXOOMJNesRQSfZ
1TCNNuBUPKh3ZQ3DapM2j9b+h8dmd9poHq8ILYw9ndmblFcW+uaiF+VVeu5RQCLQ
Zg7TpJyBc9uj8yXDgrTiZ7eX4FYQGf6lGDmKo62v5E3bDKUG7F5Rvdm95BX9XOQm
yBoHCoIswJDFu46o6XSF9vo1RNhCkrUID3o07XB644xPJXSd/Z5JURvpBKRf8MQY
v2WmIaURchCVl1yUIkIALaFbWR/UVskIwJPrrBGmVtN/ywCaTvy2bhyePnVVzmkv
FomyT1vt54lUsb4n4Ew3n539v1zOfT0FT8M5nga4Ejnt39kSDztQCHrmnxkohgIY
HSHJS/bVGx+yxcd5b0FdSrYMDbjTK3lWSKk3U6IEQulM5vPEJDalFxaR24rdcG1C
PuACjWHfl6mCJeGznwripysyp49hbp9TSQVCqnA2pIvxBpEisq+VVzeSkeyktg9s
p6z5jeXZqsVBTyMBXvDeiva7k7auirfkfb64ZRjWmi81F422D31ttQee3WCfE+tE
+jFQUOKejTlsKILjV8SIExi/5EeIEEYmfrJBjTLoxtPNRR98OQj1cgG25l2o9fyd
FTfm0ty+ELmyCgTYQbuks0FXtQPWrLw0UPIcZ8JUlUKoF5Jt5SJpwSYhukyFxDhn
cp1ZED5GvTpL1BgiBq5MAtoRAlmQJSkgZH5GSePFQkx9zYjdlEBbeKvFJqaB5m+q
W3jW5z7dPeCyk9/5VhwhLY/0p6PhDHEdz7lfwacZKMo7qGWQiXZqMMjvRinXS7Gz
JXpxQO4q/uJhexR3ThFF56Gj7t1Pa5RyPDzh72bAzcbzDO8VwSyUcOAQeyLjdPjg
MR3kJ7oDtFu4BsVuvo2P4HiHDPe8X9oPBa5acRpsorAXDsh2NMVd846XTFQMiZDB
iMoM1cnX71A1C6Htmz22/xjZFOaNrlqSjsyesWc8tEaA9yFxWR+fKSfvxcqJ33np
81O7QOL45XZ0YOOSF37ThJnNpDpv+sb2BFRfZ6WCLHQA95bUxAQHvWABl1cNGsry
v3iYObnXK2tgxMFJATty6/cH167qQ5/e5P+luNm+vMUW6j2gZ3QOBreqVs2VBj+W
P8LL/hfx8v74L/B+aOxz2I3YWwOP4L+yD5X91Sfg8/+QijdO4npt9NSYyOP4582K
da1WQEEKWqxUjE6NJp9zlToH5BhxzACRyHlK/A94YrG+MYfg8o+wHJoAY8AmQkWR
ZYjmR7rA8sFhFoLSzmPlnhr+p043SuDa1rPLkWqz5b51HXgiffkK9slXSnZbnTtK
7CMXTKLVtHg3n4dW+CdEijZCu9L89C1TzqCrkfcmB/bCToviztqnb398hvzW1AOw
iTrXOpXMZt7U76oGrGZNqkc1fbWyDCn+f7k/sOIr9Jwayys3PJPMeMC1p0nphrdv
DG/9VrB++G8qdES4agOLpZ4bdYHxdEXitycJBCU9bpsSRmfmWMhHZ136vQcZZZVZ
Uj8v1OAHtR1iNpuvkciFTe6zIYnft3aif9Y97Tl69WtdcgHRVv3WlsEVllJkv5O9
EfHqwrgaeBci43u+fvwvZodd6QThamLXUcApKzRXD5dN7ylPqzmXGzjST98Vfnez
NbycQgB4P0zcbUaIu6NS2+izD0vMWmqrWtaIwVgFktrZngVmGgtGq8P/BhWl+v+Y
8QUa/5qvNWBVMEV7VVaNLrh+U3mihkfS/TpI/GH0GH8s2vh0+jMBnA7VH5lWSToI
G023U5n8zuh2ccUIBWZsxPLDS9nFtnUr3sl+tRrQEPSG9nWYkLODyEjgpIzKjaU4
EkgVqyRNW4itZLLqSV5ajBSydSMnWgX+wTxBK8jAQSbts0SYocjyB3a+lsbUDAHI
6GaBkbGRnH/uuY+bZLNzYDiZjo9nxgnHGGd95v3JyEczZgrCsAQophafGrq/zo12
SWfMJg8ARIRbfsh3rV+CoTvMZr7uA1i0Qkqs0zU17ti0go4LesLHfK0+t0PIjV9a
I6tWmSZon/NiGAfakVYnblsx6GhE+VGg+xHbTYJ1WsCbyc4NsvbX9yfwWZRQQCrE
deiFMJjSa59vHbrGbTTRbWS0gtvRRRLidreP/TEd1hUuSIgoMJFa2ptkw7WZst7B
FP0ulYsjz5HVV9DdBv23BzT0UTXAoIyqRk3uobDyIZNX3Vybeh32dUUTty7cOzkU
+9dJKJvU5oJY7oZ5SGh/RmFE3U8kWUOsfVByLEWI4psBjmXwVnVEP0elwNyYC+xK
EgLSS/hJbS90lRh2E/F5xopcgTF7s4R88hMwV4jQAmebn21EY2OY5BNg9g/2WrEY
WCdSs5UBWS85yjS/K7Gqzklu+SF8CHBblQTVHAeKyjGlH6nvIiC/heaJniP0GFUy
yHy0auic2D16Yg8Yr9wpDx+tFVwpEwB3g69A05W/RIId1/jQIJQEeVpHMBKpm+Sq
9SmuQJV7+4H1oDuZi60q9aUR8pNcY9ZOlDJCUzBk1aGU5MqFpWlSgQo7ZZY0Psw8
kQgSgNVaznZXIXlycGlWAxM/AR/qj+jLQ/BUXCcw6BmHmxb5ve/CtWoDbW2JgHTa
vwYf9FyTPzmVHK5XMjKhIueXW+tsSejs8iWiJfF1iaaEqv+vKbFjdyJZEf1401NF
pyf5CAWg7swuCQPGokDeUUIRmOQPN9BODJ26CUe6MbiRG8obYXA4mA4oQJOSUQlb
koqU+ytQwrSHQ86mk44I6GZKy77WAc49y2A406M3iOMT6B71pJYGshkkx4wremXw
1IJY+3VyJ1NZgUZ/aabxBxAYe7ULsC7D5VJigVhHNOqV18LY5UA+lmEtUltcO3UW
mDCyEPfmMylPU836/yiF4kHa6mSvrWGtKXZkD2KgB9AB5M5onXvppUndjUmaWUqM
is8rL6/TgqovDyQdgjtPGMCHG1TY2zC3gqHi1r4J02kZEedPPas7IHkWWvibjTty
ZUq+93QyTZwq3KzVMP1kazosz3whalNiPs7bvyNun+tcV5VyZeO9vFXN5OjYPM+/
X96zC04q3ZsfBvbaHpLDmWeyTYqHdrrVsZyBum4UJ+LelVGbg/WAKoOgTADlbiA5
VtP4na3Mk3ZpkB2EiANnbWElyuTt5x9wiXVk6LkH8TR7P437coVBk90sJHmdjQh0
7GbKbdJAJx79J70gOD6yU6MzswI7BdeZT8W7LsMOWxIlDR8XAajnefMgzSFpgWLv
zwVZ/lt+Ol+pNSr9S98nTQSJIMpPERdUIauMIqQXyUYeDcitJ777DKUjxVn9CSzU
4qNol8ddsxUez9NxvFwaPZMPjY2EspwQX1y7TY3HnttIzQea39eSgnnv8uCWroaH
8ZcNuZ+dUyHI8LpE4DplSo0YBHdzcsBxf9OL0BIba6Nq1Xdzc3xm7vwVgo6sI/lj
I6vxuvecIcSyodkIcYxAbauR6b4JsQEzsQ/GmD6jZJ/oQXDwZZSuKLucPCliWaXY
+BKAJaX6MeILFsTVogdzulWQO8P4ixT/F3xLyHBGk0RliBLk0MklLo99SWFpRgWk
CHuw6kzwR5Y618gJNWxYHXIesAUkJqv+7xSPs1gM55n6AUYfwRbsOgRlQRRBjqsI
aJzo+N9m/1EGSiYVLMxH8g68Q0v/hB8VoyERVAbWVU4zlmB8j3LbXM5X8h1Uy7qw
PdTD43ipjheKXSmldSbBMFagdaNn3KyaYNLgvHj3Fl9OG/woBxI8FC6kBrYfcgcp
90hDgQJl2+rQiMkcW4xbTWZo+DXNiqz+EuXLRIJwqAHNum8DxxfU8jaz2HtUiHbI
/4CC8P3uTB/pf98yG+B243Yh2y3orNJEbldtEnoD3dXn1jKWxDv/q5RitcBOrX+D
otNcvaEE6mI+Ad/2TKAcPK2BrVXVNb1uJ5byYBlthk0jlrZo+4Kr88siJjESK/W9
QOZU/G+65/fuiLGeeTy/v29mhMbfIdlIMqcR9SEVF+Mig/M7I5sLwWuyncw7v/qp
OKBMKm4SmzAzc8xPFyd8XfjeXa4NTOLrZBRmdIjz89AUglxvCuSaahVa0mRotagD
MOpoR3QwfAOp+ZAFZii9nWUiQ24HMsyVPq7FOHk/bIZNiaQQPWuwZcqz1iBIU+Tf
WE9hNlzf2mXM30MnNEajyg8Q7UYbvJeWRFVsfE7hXj5MpoV7AYsa3lVlupkMo46D
/eB/VejYbs7WVHLng717hNQRqUtDS3FoZC9DKkbY421uZt+HV4Eb0q2qHeP1oyrp
oUFFchicygISlnvL72pDF6t3l3Fu+cfaEeFvmO0X+4d4HC4lDBRdMm3HGn91Sy2R
QoTxCFSn17dNQHfSWrPiXPHjHMfH65x39fb29/yZBp03xdf0lLC9dNtglLrWHJiN
TlY0e0GHWEpEYZXb7a7YzSStryOOCBZqUrV/ZEevmBhlnVKyTnGKclX9GhGISOtO
dJvDbG7D+aIFyZSlgNjK5lTM+k4Yf7EHemJTuMHZjr/hBpvCue+kCIFl4Pwk9Oxa
tV3yMrRe0ONcz3RXHUnFo0ohrTcqYe00l8Na4NQ1L985HLcgWtiSdDBsd6ovXWk1
XXQFMzsjAaiayfR/o8ViNVKgvgFFlbZ85fxomunx2q31WFRNMxJWXkPCn3bO/9wj
ROTjKZhayKbxN5osroWyV0Y0zMa76lDsMKFYlXjCgnKGLw/Sm4a3bgqY8XwJBgWu
cHT09Xgj+s1/MVhbWcFSXktIx3YvS+jQaL8E1cOWs2IseuPoND8HDVTENLCunUMW
ftVQCO+IvAT0uBwKY1ZYcnuTg4lnPGunSG/q8vlv6TxZWWsJNBm7Xyf2ezeDkIlG
KcCpDrrZ+VGWqSGBWS3wqgeXYygEY6rC/66NZA2Pa/uxl39eMiXXSk7pS8ib7hO5
MpxlKZ/fX1XW5+aqA3EE+iQJbVu9y88wG8H9GFoL2eDk1sCxmB2SAC3QVLZlAqnL
88E1H1KGRsywnPAcIzwvlEhtbneFDkNCDbTECPwOLOxpP4LbrqYJ1hkvwYYl1aLM
VwvETjD5xKZvLmvvCa9ZuUMxvU0x1GbQv/Y6J/RqpstheCUpFf5bdG5tO5Z66rAb
3Z9g9rNrQtW/gVQHOovinGvFOLuJVO+nKw8A7nOyTCAybkkcAfE10hz69baf9aRF
C5M4vQC0A+jFm3UQ8grTtf0CoUY/Z8Kh2jTlQM/d8qDRLH6VZESTeRN2rHSlphHj
Hgv/9R2kuDh6y6L/65casHBIIkoqoSUTTpMVZfpHPz1elFajlnC5g/6kzRL03Oyh
4PfG7pz1gQjrmhaOGh+y5gB9gdzAz20BVfAjOFDp7TqlQY92AXxUwrLk2/+KAKrX
KZE23AxFYFApXe5mu2aDj3Mh7dls1zv3B3Yirs3TyhxQjYnfCVhM48p91/czmsb6
xvLzo9T5Xa0uMEFLYP8IbK4D9BkwuAQljSWLv+au29laLl+FzViSM+FdP7PwrtVt
w5RqIccVq/ibAmRTBy2aSYZ6SjfFIO8ImLZhyIs/YlSVHB7wHZQjKm3CUAhDzJlP
7JIz8hOhOnY6nsjBYXVIaTlKBfmG55xbr8VLapzPw2WSKpWp9V81jYH0kWIWYo2e
wm2xQ0GEisGvtcUtDuZlpgNO3v7cAtIkd22dZnWgINIxkMPRi32OMS/Gsso3+Kzx
46kcPCGUEI9hFckaqXCsTgHNY8SRnLiNmhh4I0RZQMmStPYd9aUVPDGej1Gpj5J0
nvpF/7P2DS5Uflr5LkXQmuxA8VGnX9KJNpEERRUnUnP0qp51YGT01ko9aQCTcY9o
uzMmYUO4yY9U2y142HjgtGSJtlHFr3pnqlja0ZLESxVHMPCbfkJeSRJOriGVrmah
l5wTjauQzQ7WaMA0n3ByjGKIVCvPTbi3QpnoofoPIRt5fy+hpxp47Br6VeP6Iza0
0FqT5K8rXF0WHvTsJZyCLIUNH+Fops69Yerj+2iAnIml7cEIZR/j/4XmsRk3XyCJ
Gaa5Yft5pi+u5HoCX1yx9LyfprP3ejdufKxoW8bpiOEsHOFAEQVtMRrGjxLPHDuf
1NPvZNCYWAN+r5LbLMO0KoMT4Br9rg5fG/ocU/HV1soHJ+oDsFQW2kfmiDGrpSFn
vpYMi50xh0A8w+gTkfNnLDZ37pnvBX0UREnhjpN/XdivpZb9MTiMYszhcMZS4fpU
wfj8G6WhXcW6x6oYBn04VjepgL7BurlFi8YrwM+XoEoyJq8KjP9DhguxhTXbjF2s
RhZiOyQtQ8aJ2VL+Ccy8E+zwbpIiECzcW0vu5MoROT68LgroyZwbtYpnl6DnajbT
c6YA+vMtpQGkmK0c14lrzzBqvhi6j1j/tOWYNg5Eh2P/AoH+3MbTpgqAZud1ukTP
WHGh7gPW2YuVf6NC+iFEV/K9XJLaY9a/RiXN0OKq9VyCoIF7lZJHKJw7RCKbje0X
UI+NyIeQtNMCGkmVfUfQEy2mWaH7906iDNjeU4a0uM+tkRVkGZYTkvwDCbUN/kGl
5356gMFgu5EpaHzjqMFldH10uTPDKNG2B+THrdHOeQyFVCPnJCuFyYKcVrI0EnrB
xBK1fi2IE/WydDn1SggxBzWef3LZ+1t/+dJA3xyjU5eBtACR/87rRx0Ti7LOtojl
5pxa4lN4a/0kecgDWc6w7pusvQjbuln+6ancKOJl/+aok+edkHePKz26mYpQpC34
C7mj/nck9iQaik13UbziSJiSUSfQAaC1dI08aeegUEOOzg1UDdqZ0LaA8eqi5wti
O1VgYJBnoSNHqK4KYSGAK8K36wV80EUofP+blViSEjeeNX++8ZJkR+8nLuDx+iPU
80WHQge1q/S5bY/fSZ49aouFOrjgvmRs9kelyguA6RU5DZ+I5RoOdRBef1FeUIwm
bBlYuSFQSTugMerDkr5yO3SrVwt4PDSescil8Yr2i0Vcu7tUDcvfyNfjRTGMZO2Z
X9BOfRDqlCX97eNVRptLCRwPAhKxqJzZZ/LbKTeucZ0OFa3icO40gudSp6+CUYeE
vLv1Ra32Cxc1EAQ5NBidEI+QaePfy6nOnQP/tJQuDLxn3Fm+g6dV5Jlu3Mi4jyIc
omXqBURYrsUb0+gTkpXRND5PpzmBlo0BmSRzZ0ixj7ckawxRO995dDJ6OdUqgf4A
bdJFd/WCWTzLrgt48pjz7T7oyNjHDgyDjrqy0CoRwIuPDKDVB3H3LBotZM9SlTSo
qnahLwuBQxyD/8ArvA4q+/SEf3Oc+qafNDLRL0TBeTBAjpwRxO0JE60lqYnDNYEF
CiBBzS0OxtrirqVhqnUPNebUypi5QA8uCGRIctgUc2DlxYhP3GiDvYFMOaMuDbmg
ngPKzcpgtvigiM+DBThlY5kxIE2zpWUsZAdNglca1tgeO4xt27ZhAUnHyM/oQLkA
dik35vM5GL2DuERePC6CMOOBr+Fn9iaeFROZzTN+d9IWjZtF2OxJJoA1jJbH7v5j
bThUO1NA/Y8fAUALmxKeu65RlCy8YoQYN3U7awtS2jGoW+CXhI3BNOiRyugzC9yK
js2Cl8yxCa4+foZTwXOf6aOiYe439zwuEnUtd9r48432JubgACjApKgJd30Z/47G
Rsv6KvqnZ6bQaKTpI1NGdziRrywuwm7arrbLQVqRRvRAc9MyJDGigH1tU8oyyEpp
6IBD/vxfBw6BAQHbJDMM/R1QCN4i6Vrxm2YOFYlU8AMRLk3dNFdijt6xXyrPkXN/
/xrYoNW7M0hoLkSBvxL25SfqyJ75g0vsGHJUMQy6U68PP2Rqv91U3xbZfhW95RzS
fuEBioHgURmiZNcI2GfSe192+Y+9R4EFDIr1hlz2nAPvaHMst4h/7jN5zeqllqfg
m9W7+8Idn/4145D+KkjxQJhouoL6orlqdIcWwGd5M6ph9A1L1FjmNxlRoK3R9NeW
SPIUZhAwQXcTMFk8RFgnj5OS9s1OMk3660QZE7nCMDm82MhKmsPknDtXH9dAHhEF
GARZFIB1OZBoowE8kva9fUo+uCSkVASe75+Xy2+FqcHyyTlIMYE/AbMSz0XFMclR
vyOc2NilaHA+2NJ7FVKJ5Ge+AYHmqmmOxwx8xlB1V22iC736ORbVDcgKhQeA2oxd
91IeohLTpnPVbQ4g//wnWscdVOQ2cvRhxTx4PHRT+VN/+X7EAZt4xPK9e/yaIsIj
6Hmqhwls8PdKkiADSqVh343O+apUJe+fooy7IEf9EvJGh73iChacJpdGvPmx57FI
Uhcj9zviRm3me26vkrzTpOUUkerP7fr18K/oi6CQAO4JEP5hYMO+T5CEqTBHR0Eb
K7PquWU4eEPcTe5pRpxXmdtTi+SqmlZeyhwRgb2YoK9Jzyo8Ds35SyflRehqILwJ
6VItFnRYAYBGyhjqEYUP83OfXtGjgb2imnZPFVlpvaOtbcqh1rgHshbTH+HRJFwD
vM5PWnE0rmhq1dwmEBA4CqAi1gBuEmwj7mQ9oXjxP8QkcjF8qJ9RpWZsIue53Vol
AiT6nmx+yVs3EWdKnq5HoQcBfYD7p2xQAarS0ARtQcRBPuWEopNE8S5F+pvR84J6
gL9expdlUfMdHXUGHgLDrAQJ0mtdzgUytptLHQTMg+6IaDd4XMTjkIsMjO/5WnMY
Ax08isnhCS8TjUBMic9SZkwoagT5UWYODJoSLf05S4b1BDAobkyOd2SWf7xlc9vM
QgT0lWeWi06A4jHNCroXmJpz2IttWG6eOaWswjsNzO8ZHz6TenVqOSrV/wULqC/X
6KUXPWhNV/P2rMhFQSyIpDIEjY9xMwKehRpGAS9jtuJa8chcDDnkHDJeehfN9rcs
ONbKeJn4FB0dFEW9z1cMaJagdlXYjhJlqEr09TgyV9E9435qfIVviDlu0LIy0pD7
UjBZ4EOgjHfIe0zHMwgBjVOrXjMukIBs268NEYGmg8wlWzq/g45JF9M66vDX089R
aFNcMGXvzj01WH1xPMRQLCgtfGU8PGlYCzXKap5R+YQf+vpNeXnTP6ugFb9RGR3M
EqsxgFN00s5uGBhx5gVMjaImQpIju6h4P8OH+FN8tJuhpBriFMIdkWDK0nwW1aNJ
OMVEyyD1f7DUMId+LLmh4H+S3YHfPX6UGpy7KVtpPV6OPsSvS51sWzjQfyBqw3BJ
G+CQtNKE2X+gwmyDR/a3v3E+5QJJVLkBG5uFjdYo3Oid9IyNZhYoa3M5vJcrd3ts
n6fXWNemdgvaPxVmWsGGyl7USM1mNAsIy37sMAeitBFQBfvYEPCkyVcVjL1YrHnU
IA5CR11FQzNgvypc5RZxab8padjoMtV802zIdC4A7sPQVWAEp919cSYRMVwWMdRw
NZu6/+0HGdcCaMwIjBaBSP8Wt1ZmcxS7glZj8D3BXxIc1QwDtvDIWtYzRt66gZ9/
Wf93c+cermpfocmwYW0eKXpldDr1+aAVoBnTRAR8PIq47tYaGkiDaHUybe84W5AZ
Mc6wK5wcBWeo2P6P2KWzXXI+Tw8OLMBXNGZCYwVFeGy3QBUg7YH7c+a50ryD7zjH
TngG3DFjRs6Px1SlUpWApEP44l1WlbelWbASbC4XH3F2/wYLGdFacB1OJu1/ZBlT
/drpCnF0wrDyR/59xY0VQA0gtqXK3iKCzrkd/3hdaxil9nEYs8qdP0mVxs11mhm/
pdBK0UTaHAMgjrdVdgAJX2JGHIRJ+KLNHxZMmkF/f2KGWI9/HIhjQTMkIaIOELYv
bXICrrKtQXHfVv2wA3eEOlX3UqJvpJ/wXmeJzUKlblfFERD8TWXJizreJMAfj06q
qu8NawvQ7lwI2meMM9x95diBqcmoP3iQuOsoSci20TIUlqzYGawDD3wSGaI5g0ZC
zjYBiQy7yFi4rPGUbkFD1zMltErKaiioUwlkCpS2UIUqM/nt2UFKu/itWyhemfhV
Sq/BinaCk6x1muF5iPxixpPhyYVyjK8q2KPGXhH4wPayX8TC8SNXIdbjojQJTrnh
Nap9lioH7LzcajuDIO2z+qv93dZRTens1vvMd1ZlCK7vMtiFq+uzve0zgCqSYQ7K
ky2paotM1C8JPk2JCIyVghBSio9Wrj5WpVul8+/v2TZ7ZnZQ7WrGajJZ+pSFNTH5
dQxUHyEXByYeOIlmIF0s5PHSp30fMWjy6+gPdcAnd9q9EimgTSjcRqgGMZyKjMPi
j57Pjn+KYVZRJolm8aCBpVsJi0CeFGG8R7Jhp2D6AAUrBtQWHE9VdP3IAVMKFl9B
C9wJ6maGA13GB3FTCubmw7KrqDXgSNyFHBGPhUMMs1BqNjnr14Lrya+TyfKL8SC+
Ux33aFQk/JU32ik8xKtxDN3IRuqmD226QVJ3N+TRz3RxuybPCtUMA8RGVl7Vuuv3
MSLVqGt5yswtkOErbZREdwHeLzbdOVtUaGCj1Y08kvd1X8wDrsmR/rPrknJZmC6N
fLB6Oli8qadkfLAYJR5Xt9ZG6cNCL2zLuPeqLnSEbY0y2vJMu6qWZ0lsbEyrc5xH
62zcvLFwMDgdQLliCu2i0fgho3BMoPpsogvzHU/NY4SgpvmZB68Fd3t+I2ZDtO8W
L4wHuZRS0G+OLK55ktTus0WHgTsTN4NrQxeBq61KaPjwPCzEk/BCZym15i+xOd8K
Dl3lmqQADEDuo4HYSEYoNwkyktzkmZxZ0EC4AeCeAx/qQCElmIv4OYFe0ZYO95Lg
/L6I7gDpTC3PaKXwv8ztMc8s5mQSYYAcxPckcC2/ew1DBHokGRf9Q9K09rzYrm52
k7UgBdG/hlL5YlU6BdCUwVdmc3wnjh6vSNWBo5ZYYY57Tnduf3oW8Tt5DLa9HnYI
As1Ktgi+G1tim1S+aP6LuNAV+hkW3dD4JQUSyQUlRDdHP72pYfj6YP+VABN6lhia
lUcSvhsaLsg/xfxSuyf/bGNWHg5MeLqR7aUcrYK2UzwCmNCMo1yUqPwJV4BfhwgB
EYVBgeGuQP/XQkgCK0tNSUT8IwTIsGc8t7qna8MnCz+cfhmtzwYUABA9aPrNUIUX
aIO1i7Jl2FEncdt+7Di1p0PmDf1XGJksQgeREG72NxLogeM0YltRm8KmfV2TslgB
W43l0djHNFwy8bZzQkOJdJJtozDb5/G67ElH1EBUGgr+KBn6bM/nyuajiNu776Cx
e7xTxgq43JhXyNN/n7Rv+3BDwLoTLIbIF3S6hnbhtqq4qf2oRIDi77YtbuNIzFAx
YAixyWwNC8oPH2dZJe96Sb2RmXIBmbU7fhjZSO5BEZfqXgq6ZHlGDeW8fjjy6PCZ
vIBcYnC3E5U/ixBWGgJjmltObcAliSQzrBPrism/fyCB1vJb0MR0OMVcD7l9oyc6
v4S1DHx7hkB4qiansprqRgmOgLfTht0nCJrOzozGr8F1ZEfuvkSKAectBSdpMfag
CxCHKVlsn/Ionc7yq1Zc7C6BiLVy/EtcrP9aKUaM56/0ThMmgs/i3zF1d55MUP19
aMzFq4V8C+brK4vrrj+Vo9HJmbp2VLC/JziPf+vTFUPHXjMxg+0EjOI5kPPYUYtz
hlwkBDuWs/HCiy3AJLhWR0qK0l7CKmurDUmHiWW7+kpJczJL3OEQb2ueiqW7xQd9
FudS9mKCmOD8TQ1SI+T+geNIjQeusDJU6ZcaL2GnrTKjZQrlnJDoycMkMwIkhDx+
o2RDJrXGPITSzZ22m8ckFCUAwzrkImID96DEu25tVnbjobnzu2Md6Nu1kUdQlAjS
gFexr6s7O4+AJPS2lLyk93Uk0DT2u6uoAYpxlDn2uyPlqkHqK18IM0BFnEhYwNWb
r16PnOlBGvZGSf7WCs6njvWPd889DUHx2C4ar539+g+Xqf2WAdHaVaWT1G+QZjTC
q5XShRrgxrOdfPXWVOXUWl/EG3YrkT+/7MMMn1xEe4GoXPdj2ybRiN73n1cALQVn
Q5OPWXuDwRxQ0e1Ho7YWYRGv4M3x3NPhD9m6jgwiRjK0Ja/sfVMTWlsxYvMA/nAW
BHKhIb8Y+B3LfG/VH/vfOY6oisxM1nrFdEaBGWwSSqjXrZo1HY4CnK0xCUz8kHRB
lyDdyTgjhgxYvHJKXSE7O5cjQkdsdEAkWRdJ4WVq5AR6vXzusqcP/rWG/8MfEL8P
VmTk8oxQti3AzGslRm38Dqn2zL4f5BsgkiGlN+ib4G0u36bUDuZxflogoRA3i9Bm
4euxTT+BXnLb4P/T9l1x2Fe6953M5eJfrf3WJB6Trvrapr0tb6xg1NARGKfyKnkn
E26i+z0EwKC5SToycSe1U4VU4AawPbuUQVUM70qfwZM1C2VsI8xKjOgYK+STey6Z
iNFA8h+fph+gCwNlPx2CdxTxR6+1xSOOLg2n2L8KwnLGX7vP+uixHn684bcqFEVe
mRbRwefSZ1mVm905vQDPYUEg0dOTRMfEXBkY3i5jLqSHaOlqVF9yuMie9yA8grSC
ETp7fFZmLjSn26VkAiB7b06oUbp2YuIavufSazLO7LaxGnMj2wehuGczIZ9Mz4Bc
FM1S1kw4D2c+6Uh4JTt3IWCP0mb9oD9suwWc5wNhxfnXqaYJzVzzRcZg43V0H84W
rzc0VRq+MF05a7PDMHy+Fo+XhwSeRHKQjFCKTg2/DTjH3mjZqFYU0y/5KZ5EDm9r
hW8dAuIxggJsaTyK41YuVjplssXyEcxJSd4RuWDS/R2BNviLA8UDCQUmxDnUDYhm
RnbEBaFFno58Y/pOoOSstcP6EMrteZnWz8+xi9y+Ll77Wxn+hapSHCS8Xi9jlrnc
OtFtN+f4cL/JBVGSEM0RBeYF+y7AJqMVXByUNQ/8Fvlz/nkl1ZfvseKC6Ru95XW2
r43WgFs7HBWpVSRxX4yjcdynB2KghxwMEnrZNOuDEcJ6oWYb27Z2/QaQzbnwr26o
VpziDo3Agk4NaZizCYBxtOOd7rvHiWMBSs1e6JtjuVrl9FZM3EXq77GHk1P2sy0L
ZTFb1PTmmnso4EheoflQ/omEG4/GGYFXVrxTY3Oj81E7apXleMULK48Ik8xc2q6j
w9Nl1NCs65c1+oAEOfHLsxB24MMaUur5pIIlBmZqcERwJOBSKYD7ILJN1eDmHw6m
ImMtm/AW+6n+7djsjGLIFNiQIwqKr95T8TgwEDPQToL0jssm3qOix46O8q0t3eq2
DjN9HGEjzBZC+08tQvQ+n9W+ChUpxa4RbxU3g6eFH5BqIS+aEC1hwmvOuOyFbwge
r2/Ibqnx5VTy5/IxJOcH/YGE3HobDpoY4k4nAyHKQh76btXI882lQKsmCyKq+GIz
JisTVcWS97s9l/utEBA/uHeXUxfzH3yHAimhJ50n7/8Wd8TNG+Nmod9j9NiF8Li9
546q8HBJYS7PYaaPO4DlBIddp07Wq+PPdgCqh34UBiuG5FqWVP+pk5pstt2gmcsR
TYnDv2ggRS5lLj+wIvWynVM8smRKe0iwA8AmusDCxZO0oMs98ytuMln8vE+holOX
YoejLaUUpjxl113DfWqLK2FmwYvEG6m8iJLu26cy9Z8n60cMgm5Zmfl4OWGDb8WB
ggL8IPJkrjRim8+wYVbGBCE9n+EQr1LmYknMSKS3JoTjryD2KilrzCSzJEvLxEPD
40WP8BaLWQZm5pjev8o5VAEjRZYJZLnQQ+2AfMRx7hCFIS29G90uT//LdjLDhHXM
vv7g1RH82JGog7CbubHe3qmAuL9dfX8a6CoaqtfPMNQZPQbXJJytjvm2ZuEXya+k
oWMnmTpVPVyMGPzHVN3zV33P9iMM0vL8N2fBrOGSMTx5bzb4eWRM2SZ+MoYLMaaq
dSa65xJTuuWJ6UT6kRCdYvlLD/Seilht7jSdiwRoH+tyo9QYLi/U7emEuhn5FG9f
96n57Gh+J8BhVYtnu0Yg6r1X2+mNkXZZp0yvN1n7MWqD2YDnhnFdNAWB/1pD1pDG
6e61hP25RfiPrXwiouy/Q2BUSfv0/m5wIp54FIYxIC0nJasdNyP9ryVrZbrvE2Ur
nI/iQNj8Vqf4YqFluWRw0ChSVYMcfV+oYQvnqiaFEGAIERp4+J3ItDZIAc9Z4L1V
ozvgcS5y+7BYuZoGpyjY8ouVNXz6jJgng+NS9wv5WhOvWAECOeA/LPw0F03ZoamQ
Zw90iRaJGuquEWmJHPh5IOJ6gZVK19ZidX0/WlW4c3RK7x9Xn2/83OeT6ZGOLSkU
CaIcgFhb0DIm1mEgmUf78TXmHMsGNL5DVy1SS6btsU+vBiBFTeYxoarHq0JQxX8s
b+n55HTso+acIjox3QBqAqGoMf2UDJlG4+H+nJ461/4dkI8xvExW9B5MjQgnSAUI
biyvvvOpPXCZYoRzlC39tC8dOqoINw+1Smdc6Yo38bBiba95Y2GYyZoTyH7LHjUE
eNOPwH5pLOMnJFRB/7rnFIAReU+68z4RKwVXAwN4xQe6dmsEI0V7su+Gzt9c8dgP
TLH/hMBUfKMjwusjjZoSeejbraVQPYSkS8slCzl4K3Nq5BG4xXNa8a9v9U1Kuq1L
d4cGGrsPu0w7clqqLDXqDVNniHNOFESCfVcuV19sXvmoneXDoRrKiftFfOM+P8b9
b5hek/pVpJb8W2874G4GxH6gaYUGAzzv3c6D2iCFghccBRs5GPX7IYH4VlmZC3mH
IfvVlcRMutdhpDohsSXuDiIhD8XNQMrjrsHx2E1I7njHaCncsaNYDjRk6jnhVpFT
zKJrGStn5/A2EfT5GilUOzr/LDShuhMJqSnCG+lb6YOOgfg7jbNvNHxdh8Tbuenh
QkBWlARVNQqiKXZ0N5YnlrtaXK73j01WroQBwvV/UBg5ODyfUnEToTGVkyBTrigt
Qt0r3j2sJGd9lLoPB/Ein7HprxHniDXOJ/u9n/Nq6KNkuNgQxsUjIhbV8Z45bFkS
eQoYg7lWflQrvY8KZmck+aUpi/AqhEWLMpZzrgr87cZ7P+TOnuxozCf8M973bhax
6BIWm+4vqBohhrriogkQTNfOkyAKTqPOPC9685xLSOPNhOox8P/ANzDatY8lEmHu
xupVyKW+4sWdZHt51hZJFufQO3OMeK+GDt+myzdh+YKt5HYbirgrb0emTKe5Nshc
+A1SoEMYfy2LyJ+gEKvdLjs2VAKKNui4KUnNcd1C65UxxgbaR55mdAnY30SgQujT
DGT7Xrud5RT2T0pcZRd26+ZDob8hA9BVZ1xBvsHtRo/W3kEe6nkMslzmvH6EXRkv
fGB+LMDimxNkr3B/zHTQg2hQB+3zmsc8SDgym7P+2Ciex8CNluplmAv0C8migKDy
A3t5WjumoMv31omBRtAOpS/JZwTAecWJ3W3YEZmKvSb+4N+qZBoND6AT1Pco/TUJ
AKF3CQoUQpM9YwUSWJtuBqoJgeKmvCHldIBH63BaK51520O63VJoLongUgt6afFt
HtkKCc6/wz5iNoGhfFbfggQie0yEk0VuAD+XxVd4mNBcI9yV6GN1pb06xaNlj9/c
Y7TTF4WI8aI8HK/NOAUdbT56H9NNFKZCzMe4L9qTyS5a5o7X05guwj0WfAkVwCfS
GF1Vk3RmoHwYytAXo6R76uHHodl4+lwQNqm8f4I5CfYntifvZHWTPSbhSISyUSnr
SZ/KcEYhtPRMnVNWiNjL8SMexsFl45Q4zVTSUHgFrEk0S1W0koTPy1NtGcrGZPmX
tSRrwi6m6PRFslai1QvR2pSPAI4fCox/Vzt89mYlqncLmRI3RpabplA6JMJ5G2SR
DYjuhXHqJsg6AZ9kI0BahrPFmkHZFIrXIoS9r8Kh+f4mz0P9PkwkEi39vFd99OdJ
AVofcS34WuTEKXbdDiB70jmni+A7E9hQI6jpr1psUux0TEWrbDqPXZW3T4yZj21E
OXY4Ne/15ETnH1/DfQg0kBvAmfumNcQKaeEqIGNe+fg3FIqVNUjiXXwZgGYh+rRA
k9F9zFTkr5b4ZfR1DM9UzuRsqZ8mEKFZwOYv301PBrev3H7eyGzTKmUpFxc90YG/
l7lAl2+gOaSi2Q6QkdxwBKK/5NEW1xjpj+Rkghr+5kMvJOH+JbAw2QIYLe0ug9MK
9d/8SLYD4lU/B9tp2BcS0Y0aMxKs5G9EuQM4jr3klZVEhsk+15csyLgs4Le+crq2
fRO/m+1tPj+dIx8apAwzP/CQHtKftMgpTENA8bcFU7Np4cvIzt6xV674vGj+a1j4
JkH9yX11nmnrY1QdeVOaqt58CMp5Qmg6/L2RSRvyuBpwvW8ZbyAnUNJ9pZtXQvEK
Q3DMJgxnl1AT2q+GYpCvHY8tY5MPNFEOyHDI+36sOAGCs/xyth1vVGGVbG7EZXAr
bzKFz2Ll+hPgkLxTaDGwXPRfjKIqMxkKP6+UYhJ1ZYEQnbjuZXIzfDQNF835wyXG
KUxI3QrjiOzQCjweTcwB7c4jw5Wc8KFbCTw1U/ReaOihkMoCVEfmudpy2HFS9Umi
ayPtifAqBUqODh9VTk2+kCR0GQJ5jGCohPkifHjxf33BqnzHMcZGjzADODEaVO7F
vxzV8mOSuK9rqwkUlOPPRF4Z+1PinP2orydTrRLZ14NOLmLVbWaI9Z9S7OfWMzP4
Vf9poG9CQz5aRgYHSnCvnU259iVA2b1uZZQehQ4zCndSXuThGfILsp2oovDE9GUC
eHqLX3UGJ7wbJEep2O0F7E7idN68Y98hMl64XSxXAVeALAe9vQSgRmOzV5YZzQ3G
+Gd7itR5vTZWhYH/CdZdAdl1oJcayX4d5EQpglKiy5+7rUYaFMG9J4FjBqzw0lQJ
tF8cHCt69po2bjR/N9sJ8BzUPUqMjZH9xMUjMfXngLab4lmIgY4GO3i7qITevRSQ
IIHmp/tkM9CwurBigKuPkxvIlItL0rYEZsobVaHHGiTYjjqatzjdyZ7hlQ32oEqP
oTwXkmbolRiE5nKtBX30VqXE2yaNKrTNh9cefIhGV7sufIFtTDSzSzxBnK3I6xA/
oFRLqZvLEdDHMx4148tAUFT7I5gQ7TTf5LO1VpAq/fe1sU7E+MDNvWI91+7dutLR
M/G5XGsA4PIITgxQl5ZHMjZIho7CgSwccC355ZajMvhLfot9FiXgPACrkvWrjZvR
A+sQO+rzshNFw6Jh5Z3LvpxYps4UWiTqsybaRZA7UsoLYig0fF+Fptj0/5v8y1yD
T71K0FdR/v0+HsxW2y6584AH1Mk9Ksj2ukcrLRJbJT4BnN75JejMpJShO4e8j9u+
h8yIoJwvxm81PYruTviyC/xfTL5EwcUBf4yYCygvpkJ4GbTw/8bJx3pr9gORk6wy
fViWoUikDGRkXvd+F2JQfO3aZWlBmwq0YQ02H9hKqa7jWJHLn8Y0chGrgs5uOqgP
wv8u7RyPFtApyF4E82K/5JpjJZ5D5rvJ87j0/PhbAZbNyZRec0PpT5gFnJJj3nfM
q+gU2nsneOPn28IDvX/o84g3WNRUI5nKZoA+PsMoa2dJnyyJYYS/rJyoJD+Ue7f+
FeAUDXD5/tlohfF3x5NG2C4wGY8xZarcIYhzhnt1ZR3COUI+38HOqYXvcr1Xg1Nr
4sV51oBz9o3FVN/Cqpa0uJUMNChUOyfqRf1QjtKzFfBKcx07h0uZa8OKVyoDAts0
Y+CSscftOZ2x7PaHu8Ok2deaPOjUBbI0CtXJn4eFOFhEAd+B5WbNqx3EG5fdvQIQ
Kh8+5Yy8U9GYPb5MOhcTQ0kKis1DYSDiR8QUz1VufNgx6J3YQO/4tNecfWlSjezL
PrIHNySIGrZQ/8NxC2mv2xN2pSGgqV/LBlr4i9yVXBisyDMCC/VYMTQE1GVQ4Cvf
O4dv9GW0EiNfk/GCfne78rUAGwYzHNfRXdZUZvPkpY1hHblEh2Lce81mEjSDebyw
a9RE+uFXAzRm4YSzUYBpFG+kqwCoSKnPQjZsTQqL6ROcFyMiiktav10rQT4H8MwE
1+m0rEYMrQVmQdR6kwD85LF3/2FDSH/3zlNDe+/JYqFh/rBvQuZ3KbhV9x4FBxVm
xI9Lu3WWyIUJLAc6IoclpOJOl4ivri1L9X9+GwtvPWaLChK6Iz3mGwc/iRf4tn3q
bp0vSzCjI8t7TuqR+KPwJEIEAUm5ULir4etyFOuWGStlWuTMlxlDAkKMtwx5v5iW
WArjCFkC1j3BnBjNGLWvse/Uc6eF8p1EKXlb30sMGuzbnAqj7oRKrbtkbB022l6j
qhOsw9VKAekwSdrb0gRrNd+/Hff5uRyFp6qr8Ydm65z3nxNbB5pFNEfpFnvs053V
L2GxIGrNniE5n1YW89oABDjaw1xToEB0S0BBTTT6vVRxIztliq08A//ql5OgPXXo
w2ZJX0c4NZ7mlhH+nVVlS49Ld2SzZJughUs+eeMHB8FSrQQ3sPdTI5TysQZjm1AY
wobx+IE38g3G7NeaF2UCS23ee7t/PYhRYWuKrItUAEz//g9X3Iwp02Tyd25JMVx2
aTeVMP7+GOG2rui/JuOaEWTMRGGYCmgZbo9y5wpf9au8dckWSCxOyh75JcFmYn0b
HDp6uY7tXJUPvSydUAAMid++7aovU8pbaTJlSgIEdRysexR73GpBB8QRa+aM/qKA
5B1rI2sMv+i9YZTPWxv87XOqNhZTjYtFnwRUtX1FW5sl6HVbIVUNuB07HUiwDUvK
il1Ra+Y2NA3jx2PtfYv/ALap+6ZuOWXzj6Rz0remXbNG7lHjPo4noQFfqqgHtxXY
3XZ3SwyPZIOi/dbkgp6cxaxkKJaMIwyxdHw8QHjll4GmiN+5VF51HQYQLquB0u+1
+aRSusXumH3s3nrsepmUw204Wodazjs3xLALqMwDrScpFNMZT/CoLY09zzUqxNFX
dYj0OuDVASK8ZOskTg8G8PeS/ZFE1uRLBUQ2otr2cuUET4C3jL8Fm3YQjBcPKUPW
Kv0j6J1iG/VVMCUNveyGctF/8SqBr1fgk942J14N29kn+A20WhbHVHkf88xtlZsd
q7TBvs3CDJHLuYvhAAAMS6rIdc2rhHEZFTDLQuT45upCeU9mjKDusGU9yXCYjl8N
MhpCmYlsVZACljoL+CazAiCdJJRHO7putNZvi8F2C9opzbPwlguHr3B6PPk/IRhU
Bmp2Wt8IT/LWPvceqRX4q9PvPFVihcsSaM6QspPN2zak1VXjVIwnsTSWfInlYZAz
p09f8FPKNNoKxVND82TO2ejotEIZbauoDVpHyrm8p27CJIIUGocirvNIf3e7VCda
DEndZ9zQb2J/PrCfoMJP24BXJyQnLJDbntyUCElUT7VqD8u5j7rqQ4R/bcvp2Byb
mCoA2URr1IIfNchf2KXfUF0sxIRmmpJdLo6m7ocRDWG4ZbLwX4KY03WiJvYc8oqi
TUPZdgkG9lV77d7DNOwlv4JbHGawmzztwM/78PJ5LYhoofTVHQOtw7znEphxt3ic
F7dyg51h+t1kopZFYTAVgXAGWUYOgIopE4cbAH3NeDXLNn9vjkDwg5r6mj92A1DD
rDfGykWJOhTcQ+Qq+ahGPZ1pBudPVimMdASxvwNLAPOQM+Z/Yxg5+/E/nifkqYVM
YwWgPooo+akurJeJLtgjdW165q0k7p/EP+IiD75OqIRzGMg/NGxQiac4mGVENdKq
zw591UUoWm/WtyW355xxTEEfnmA95vrZO663MrNBmn84E3Gbn/+rkZM7+IVS5Crh
ryZn888iAwORk3yQbk5Dk1L3TPvNQk/gVUuPigqCdS8bTbKoUU6qLB/S/3lQVI9L
fnzfT7LfG9BMQR+HZuzuGzkR+CmklJMBNg0F9vyTlhpRoXz2pp1bvDASQNhTirOi
/FfaTmwuBGn4K0yeQq/LBK5fwZXnw0na54q4bq2P80V+I8u9SWRiwt8XYFEplBur
mRx0vq7irAoAIQYBg7UzePyBjRGqaAqu/2a0qBvYMxkRFVjxTnXrhklTH1037sY7
Zm9AlqyedaGDm2n85kgYG/3w3ZkZEuLS+P8MwdA++lljap2EjCFGGPqw1a/1JmtL
ATwcnCuon37012YovjIcYAyww52jPTtSoaUB3p9plAKZK/xX8m82pYmos6fOlwHB
/owdsST/0P24ZxWYBqzfR2y9X5sgt8rRFD5bizv4qScg9r3BN6NxzrqQX/qNQoBi
je0TmGbIKoypOX7bb2t6z3b8JGGtFGVfu6kFpmLyHrJTZbcPzyHleyDfsSjdLnRQ
gBHYjLJuHuRIKlak1QpgG4oceQgsYxv4KlpP6EwuGDRULy7q6Dam7HQHOaMPfA9s
j25n+Kig8TGEzdjqbTjjHEngP4vPEvJ1x98obZUyLfH9rhvWbgf5q96e154aPsRO
xUnH4v20gNljbBWX+BQlEJX/8qLoj7rsGT450PEcHDkjs9iU78uay1wOhAW7wsh7
fkHdg1Ll8uYqJpNrqXKBVrdAAQnT8GjM45vzLS4Irud2WppPg125hm2r7O/gwjbz
g3gLzw8u6nAbWJcgfI3iB5X4JW6RoReIOP54KHEbfqptRDeJXsSsZZw+/1g6iw5G
N/MPZJC7uVOG3/8+c7/4pGITFM6n8SqBd9coE0lqxJ2Vpo3tYAhMVOkq0zyuIUZG
sE9TKVnj4whQvXfcSUXOnOeSCLRuCmOWAe40Pwwna/9at8wQSwyEVFD/ur+RpIFW
WuLjDZK2AbS2xOv75vFv01l6QeVsCrpHGmLoEm+Y7LcYCuJm7mvRedSJP1QhGMEd
SPJ0RfvIHxKb29WhhJ6Ja+Fpa1Hn8/a3+1BsKy0MI7I34HeHLTSup3Nt7Trf21fb
JJF77Ivh6lwbtsH5hZZEIuoh5E/HLFJem5xFiFgh/mNKubNJ4tyyNoLbG5pxz3wQ
/9Argl5lKTRpOviI7s6WXStP82ilAZ8AVdn5tWeBcE0upfwBXlfXID4s5vAFBk4M
YalUSuz69wFZH+vc6L6TftWuXGkoTysn7OHW/E8gL40LjV0QDqg544K3iSj9gFe+
0/pEbV6BXzSn0nhfsj8t6CYKp1DZYQ+Z3PNiV6QmNBV3+bBkxQ3rUYOJ7KFAuVhM
N5mJbre7BHxd3WIhbf0E95LXoZizCZMk4LZUvNy9vyhVX+KKByILS7wSwTFCfG5U
7fRdJ+Ol9m0NTHtWL2ZfBn7xhH/cVnOp3TcIjfS1iv0w+ePthwV3w2Vi1lLActlJ
jKecI6EQ9tbEIHxHcWXxep3jL4RLdqLWNsC9MpRdSX+UdyPQst4mukOuE+k42jVz
k4JG9Z1Hw3DcrBS7UZ94P87PzbvqKJpiqFeKVwQ+9BtVSG3GrLlcwPiewxjTxzmz
0TUAIxysEftFIYRZJ1IGl1/ZnhcAbEjUGUAR0G6nYcWG1nMNftbQuinikWmKcnz7
0rOSIoJ4GRIJpbX5dvHwc9nNhT0IlLd0VXlK+jwjioxuP9lwbhmHxz/Z55Apyli4
6B7giSrBi5jYBiespjcG0ZPmdZVsuEYcnYrYxS12D7408xQALLJ6f4OTc9n2dY4v
KtD2TRAS4iDVcaE3WCrANeZyy4++FevXE1Ush5LiadZwU6DSjLhw1ouaL0tTa8i2
3kwhBHnMPs0L1Bmnp5w30dpvy4qhe5pl8Rp+hhduQ0AdZUugqpI+yvFDcOiHSZKg
xjFCzGXcc4KRDzHPIv4HahyjAVFHPDQxwhdAkCHrin1xm729nAkGVQ/2DBx7ZX/q
Dv67PAItNANjSm/eFE3XW1TNoLc3QvtPHSKbUDxt68CzE0nX7M4iqlGfi1DQSVLR
45cv6I0La+inZSmMYU8z5ZvQT4QGBLXeym9RLB4gHBKdlYAAFbjis/Ax7h0MmIjV
0a+SVOfNkrt2PcqDOekd9qcPfA+tVzE/rruDbbY72f9RcpTbqbwaQfoooppdAG8A
jfQFx+jYnB2zgcyu56F3S1d+YqnoAfASvAUlnUCq30JPf+6TaOnsVjUKHO31+Bh2
FrEYVJfK7kE3bz3wEfAZ1NH1cKw9U4OiRohWm2IoCyq4AUIKuaE2Bb39497hS6ID
KHc5CRQ/YZ5dMUXQccFa+YD9byWcGxPQP3KYSbtzGoNTWUUYJNLlJ2fyP5gxQO2N
VQJhKHpKxkDfmYaM13Xy23KOTgC4TphFRDhRdLzIouzkmsxhv0izBQhjgJMa4/LM
rTvbWXSKaBWHgyTnT650e4GkYZmzo8ZZi953QiMgauIoejxvbheGbwM20alTa4bp
+MMMG90EKlgUUcY1Ke10E7CxlSQtBrl1czjFsiI+a12TJOBjo+BkjHA20/f9kos5
mD8Uwac0V75BXzs9vmsyAL2g+ougQiaGTrjZKEQqgdLUEiGdLDlBmAzhfdLchOnK
amQ+5hAbLcz5tSUh2oyiIJtgWI2nMtI71Ckpelw3nk1QW8T54onOk22X+Nw0ptOg
Gj8Ef1KdE+gtGlJt7ktWt6vjah1GU0axvQcMH8jWZS1kv6KRYWmWjasz3gI2Nisc
iH6dVoVb0+cgPZdmpY3+eIsNOGq3f1dF12qYvp5X9f+GAmO+tI+IXq5uYtWB0fSl
R0CLdMYqcb/qRhNFjBwdS8GugmL3KKv5sXmRCRmZ2Ms/SAd3So3Z4uYhIRCrQW3A
AqpD/W3/cs0w56ImIyb7sitg5utUWbTko1hPkgrnlcflyeVxakoLTAZmmyNShWgC
IGx5hdxiAGcmw5VqfCseezktjRFFDtOJITB2WfeGx6oCIMxc8Wg3ZDJHoGlXHVBt
O6W9H4B9LS+1N1X/EjMSZTtftFi/iJiQ5k95lEZMUl/aEHroNScdCrK8M5PS1xJ8
U2zYRMBs19l3ml27DqmQ53k4gZgKOCCmQBVfmGVQiCzHRylGjpb4G6byFgZcLD2j
T/n3WG9wpoLEyiRAiPttiSseXjdDVQCvmV/aC+UyNDcS/koGTMIUX4I6ioOUwtgt
hPWBkSVg/Xt3pb/X3rxVIUSyZFKkSB9gIvA6lGSiKmOT0BJui6OlbeFzN8RFrz3z
0eutGLafZUjQQ+tpS6dPqTJgEeaTgfJ8+6z/fYcYSFc3hwm3NhaPDTrJWU9KhLpb
6Ic21UJHXFzts0kn32uiqtqz2JvJIOxbKXcRGEF2RMiSkt0lCKnc7SAUbz9OLisq
O9QtbtniUuciUWoZHltT+0YICp/oc9Qbx0HX3HJA45zLr5YTry2Z0UJjwnuvBxPW
d/yRj/Fy9Ob93cimk+A5uHaWb3woeQoiieeJxLtJbIgyF/VHbowT+ZdPSm1mieCu
1t+6WH8OkUMBSsz/hlzDHPFGkO8ePZrf3pp1ZW2SM//x8x/yah5LFMvqe/w4Gq/C
uhVS0J4HRMQC3j03L0QEYYEulSfGiAQTzvpVs2jklgFNK6uPvkzvLRtWJXEcYj8+
pmHi35uZB5G4e3CFgSyE7ZAqpPRLGar8SXXXoKjQB37xALOKiqq0+KOqbl4qVwoV
jMa9dU7U4ECqTZQqQq7/IFjpBV46T1K6ZshHNn4Q6tnZtIZlFd7ycb9DCyYrChpm
HJTbQSPTFVL6esTv91W/7ogEr1xOjKlddwWzQMLiU2ehsY0ahZwyF0VYntyqHTir
PnyUtZMyACy60JBMPtK7dwnkl67OrMQjQ5J8SwmVz3zG5zBcAuY8Eq9smG5UcwuU
W3Ntm46ddUn5WemV5g0Rrf8PfGxHFAFqqV6m3Ho0l2dP2DsnDPFBNGYqM1nPStXH
5nnpbrIxRecGqHogTiv2DVyPEdPROVUc5V4NBprLfahFyUWumH+wEvUuMTQSgQ7L
hPFY3wI/oVPQ8abbJu5IEclqyNoasoE7Xto4noE+rRmmGY00nNaCfJrbii5vRp19
0oIIahE/ym50v6CWHbxZbtzw/+zyOCmCsLl1wPBM3zysr6gMn0qfZLk8L1aLTJKi
wKtT+dPdc2vo7InIvs10pZUoADuwsWt7Sws5XzRs2WnpSiXPguh1t3zvwdlZD0C/
5yNy/2Opt23qLZJHVqLcqHfc+mAEo086oDduJN+IcndKk4KcuKrqQ9fBXjfqZnEl
kpCiSvpzalWJj6Afiq6c3OSqUQus/d01lwDBBjuiZYF/zfBWNbS8gRHX0jm0ER6q
44stxDpot1l1nVtICbGJTnhZW8XsGB3SIwPBEg6Y0l5jkXgsBYo/w3oZAyvz7Nru
Fpt/i5y+qBZw+FtBJHxvuC7wedALPMGoNnqb381azEMD+ndfPz38J1anJA0OXPw3
cH7LLs9bH7oPlkH/s5lLKw1FD6FCiCUbImHJs9MHniMtR1E1xDa6505h93bJf1r6
d+8QzXjEFno8FfQmAe3c8KbKn2GOHk4tqxRVX3B5vt5pbcP90BxCwjwHel0fWimn
kz/n+CReDYOAqSB7E2laxaoRqGgQ2yF/hTY6hSnwdl0wH8eRsSvYIVDWNZzG/RKE
HVaD/8t/YYUd7FvgTmddeHJ6VYjAbhXeusUJD1AdRL3vCKZevEAM4xXcKUsi2urt
2uKk1CgLq5U5X3JFWrRwDU7SiaPS7OFHFR97/f/g4GDwiHtTAaXsPP7whM0wsI9/
5q0Qe5I/DIzfGddz9GfgLXAzSgacflXql4xbG2W7FnZPNFqF8PBE/750DYUUu0z2
CjDILp760KyS2FaOXVvJK6hMLfxrfLy6JA0SPZnChP6lZI9wocxzJ0vnWkNjcvAk
sRl8uS8eZf56IFWCM+B9bTCrl69tWHkCrONzS98lE2fT3vWqOFFP44JHyjhs33/v
cCUF6bPNpsi67hlllTjAlzliU1rzP+a3YAcqhXBwzuclk+GN7uQ4UYzC72u1fhZy
lw9JKCAOt5vkpjZbaG9uVcbzG/mzidEPdMBSwRwJqhTx+wImgQl0qfcecL5NFh5w
bHzXowU7F8bbezz9NlDh4kh8qdrYxAdzwLZYCEHy0vXaMNR/6cgmxBERa9/K6nBW
d1MPUVCUNj8mm+yDqMlZ1Myp1YKKOCrfyU1ou2cu3M6mve1sEmLIL8LBC+9Di6kW
tDiFVz3n7ny7NcM4WLhZ5dbKlY7dGqFZPU9F5jmdFsqUY6mT9CS+DSM28sOmj/qx
+gkpwOQOVcLDmMJu5/RxgbpKiF2SLJqqlDosZdNls/yJZIHSp4rLupbfHJGXG55O
oUqro7DunjwGpl9BrpeJxe4oL1IYuJvPBaUNbnDiFpiIyf1vkbVSS9QZkUtf9kui
E4W51/pUEBllKsNR7vDNC/9T155iHKu18ziC1t6sH1Yopyzy1bqHxw2Z8OIFSjM8
yVraqd4V75Isy2YjTEMOAIlJl63byalQxU7AmLdO+C7m9xkFQdah5qDlbINtsuld
U+aaSRENEnItPUiBN6PeLZL7mIFr69OR/ki4jsqfFTeVT5NUOXZCUcVc4m3mp55T
XVbWfccjstC8J0MHwCiHZ2426fB2V0ikfXwDBurewlpWNaZnIGggVcDWc16SLHSo
leBq+dIEau27B4O6egDV38IiGRFONRiJSf/I9bIyAkluvRTqHakW+0c+ZYV8/q7W
nyc8F2A6WGnBCaIfSGufokuoKxLaVGRFNFVWN+7hmIqeNRB+dc6+TQ02lt3+W1dq
KO8dcHirZc1kjq87hTuR1pcQoSVcAkyZv1/+8F8BqFwbILprz5ySoIr9bFtD/b4S
YQ3rTzFnjbVjKZf6JbUGxCk8+s2QRLkh/KEB1TwM8dG1STnuAXPQzy93TqvGlEa1
wU2co6RmPIfiUqo+YcZ0AK8E/BcfsPA9xV6rQGC/kJSKVD/4IQwrq+wA1KNId12M
Y8g0kA89D4L0iTvEeFkgZhuX148qKi9dxvjM4Yq7qzVabXmviCrKkD5uRiD0S5qT
Lfke02j2KpUb8DIBamP+MGPw1snII0HChdLHjxXekQWkwGSq4QaBynSN2jGyea82
rPbe2ZDZRkQhfqGVZbS+GzAHe/IXv+gud7ZmIhxB8W5HVKLlz9nIYoIKW2do5AA4
hXYCQ9CspMbggVeBKgAdnTrGwRTjEKuFch7iQODkEAY2v0TbBWLTCEqRrR4xw2RL
WnAA8+nwd7Rl64tr1u+4FyZyz9a7foPcw+BofPrzuq936W98mgM8urdHNE19x6d7
HBbm92jWjMaK4ZKVhbxtXEjGtaeAJqreCjuwE6AM+HSY90k8TLileSkWh3LaXdB7
02Dk30BYYC+OXgPEwaZ7m/f3PV1VHAgNs3lzOcaucs/lyqlRmBuYXrGAkFnOwjLj
KkWwpp/CHQ7g4VGHlT/9JAqs+4HHARIKZZSLuMWzkhIL0ABCUqKwYXMX4/W+oJYm
e8qn5rBhRB/+tPQG9d9GE6ndiY3uNEgnwd3vkoEY9eH1rbYdp+j+yoYxZZKph2Cs
2/g1e/GjS/5J+fE4uJWPyh9sgk7O/nihw/pdcAnzeEOTuFj6IphxkioVCJgqFc9y
KDjOed8wx7fl3aLP1u+E2nO9Qqdv1Wad1rRQp/jVp3oVxkbIGWsjjuYaK1GE5Fub
xOZeyZdFCTtl4tEayBRXupLlty9As09ZXqh8IuwkdLqAA/NNJ2ukv3XnheQFrldw
tuM5tPt5Jadpkw8rjH3qWGOEsNYXHVHXACqF2vFD7v2uAkN8uHz6ozLdL5xEvKwe
AkM0CVsWrQiDRatjxwdD5dhbS5OiJWc2qkPnMhDr8Bnh6QOCY668LQZR0BeqWJzf
5+XiMUBapEVNT/trsAhMPemWgd7+uIvawj6bkMw58ENBTyXeuuEBhMyDUG4u2VC7
4G+k+VUpmiKVqbJF/5AX7ECRiVNYbjy60XxGSOnrxIq49XWSXP/gE5GSt/S4vt5n
mM4MICDqBCv4OvXWVM9Puip5A4azaaqL/GYbseiShLOzF78PXrRccoj1jFBii09c
aa75cFZY4WWTZiTVyQSCaL9H9XmaDLi3bYXOxPj7rNwCk4qt1THAWnbLuSOVM575
6myHqFxR/h37zqQHMM4hurwAP1m6mXYt308xxf04kN2I9xOYZJpaZL1vIGyJ0tXN
e+U+cehOuy7TCA0rhvT+lHC7S/F9b2Qq+gQRYFIOjl/8T44cL1zVinKtABvBFf6M
X5iTE6QO6DCOvw1x2hnh8GoVcS+aKACFEbUyl5RYE5bMDSS2oW7A9Z7LEDnx+d1b
en79zgvuL3SBHNCr43yhWoDkahNKSv5tPFHopzC8b1FSdEeklLisnQ3E+6W1JwmA
1pRfqFH6GpvSBDS90AhoDQM1F+Euzpv3BHZCTONM8b3jrtRv6GGKrlcn+dwSOXKp
mLq7toGhpMgu0qu4QTNvkZZDJfVWdIQddMQZ4UxYeuqgHkVBTj/WnHe+NNy1At79
lNV/Xa7u/6OhjIbxocF7jiCb0jHD7fEhEPb7XPt1tEA5tixrUqai6EX73Ejwk6U9
qtyOiZvn2JkpNN/Gr5gt5TAPROxWzB/Od5JiWqXPkJKkglTnOjXWeldiVT1oHD5c
7IS5POlhShVOrLl8EKfS8C9Gt+xDjeus3aTmEazuz9XEjOfSHOdVeob1231Aw4NU
0ZPkvtTiI9mH46l9dHd+EVeYui1XT7hgbsXdRtjwvko2QoJbFIbZNFNpvtW7NPuX
sT5kQNHeUdpSj2iNAZUcQEpl9LOYpR2fQdgXsKU2kE8HPhDy3Y8SnVnc+9s2bHOQ
0iJ74/JO3GAdU0dKq6717eoEN9+lpk3guys3vsbgAHWpomztoA+U0ti9arS6ECwE
mBq2J84S0CvUQYPxpjq7qRPCIaGPWVp+SSn9FdZwAtzPGmgoBCfkvWwStoYlDWxD
5XxTs43W1/8cHQwL+4DzWGllB+iQVxYnqyhNbYrfdqsS0WwJ2p9RyMwqn9ussGj5
L0f9+oZNZ5EvM4brAKsHq8W4vMERaMNud/fueUDSmVR6SpyRetuTCYJIxm0CxWCl
e9cu6p0utoHBu0llaXwO1TnpQnOvLhr74h6JJa34Cn0W9e9ZhC1JfZDMk+6sk7W9
owWppCjZgq1sNbCjb4/4t/PSODDijBuJc7XyuRa21OiX6kZPzOjBt2MnyAaw73t1
AfECURYgTcQTdBpgIx2RWHu952+xYR2D2oBQwiuWZRHhEpBEkK996wJLzffq1KoI
2PJmvcx7ZXOA/fw9DU3mLew80D9PGPPmheXA+FXqb5GX6fdcu/Am0J6T1NheVqv/
PgF6KHyR2epTazlPh1uAtJH2ZctbEYM6phKvANY7xkkgqAtv/bxKcd7sWI+SVQUh
oCa8joovCAV8XaA/a9ofTK0lWGVuSVs1GQPQ9uRzlYjZXqePrI3JUFgrfxm5tdXM
EqHZiKilstIy0b1J/krKWuq/hgizou6714WdNKTav8di9QjF/XkZW40RoLOPjUNv
sLGakqV/IEttUmjaOPf6K25+WkHFLwcz9OCvtQVABpYtAathF2wAgTeeOZwtFVL9
j69ZW853a4U1UdpW0aVeCS5AoG8xzt9K+bPY9weJk40w100O4fNZplKdoYfoZF4M
DNSt3NqAX27aeMf2acqXVBgUG0YW0lB+S1+SI3VqIe2Is/sFd8uz5pfgAm2u5YKZ
XU2vDWeHkraAxjX/gkjgAWmIYE27SK+Ova/a7HY/JMiX98ylyRz78PeZKuiUDXpt
UOD/k9TGQHyox8r8EKkg9EoaSaGtcQdvjx7l67mbBrF1H7CNBcIzXjCmxcWxMAXf
a1yJ23d2ZTFuEtYyfETqwHFDHj3kwbZeDBlAXS1aE0ZSF9nX4ykgCwrEc4vVuSxT
/rTVQp/eyHd9rdVTn16bzPQMEobTXjgOqznurcfcv/eMP0qqwEIbvxVf6Wkehop3
Ao5t7MmMz3P+iAYscOz776HFHWljY/U+eC/VaytdstWr64TtHYXxOjOmLBjzEBmV
5jZ4xHlU3OGT1gDIxncVKdtvJLfBh9Kp5oCu7r8pD1S2PGGFQ+rGzyZ0k7skkDZw
YINYSY5y5bDTblC9kjJJvVK0ERKNUZAVJ+YFZLVX0+DGr8xdEN1YvgYn/1p56BdZ
hEFckLtYJZ8iI+4HIO5GXINuvo1jqI5JUgBLIlIbeamrfwK5r9k+ivdo+IaZa2G7
SmWvaqf/prq3grlPamVk8J+SBqFYQE4jhtqk9R6zjJfkheuBYfWLTQy8oaw8Oaef
/ap+qFtUp1103fTSyEqLeLxuwji7pfzuJGZrxkFJBbaDqhXxhLfDh0F/5Qc/oomF
CnzZFEZimQDlY8W+VDH3PUqYpVmR9Q5H/NK/IIN14Lv1xWLNavT4jh8ExPuqyaak
o56u15nFTRLP3HvYJjsyiJ7YysJjDcgvTg7uBtfmG3uvhcHxMblRiC4eH0hV2xQt
grk+qC/qkM9rep5tAWHc0zcMSiIYO2MYOyM/hQFG+tv6XwKHtRVxbK7jUno/R7YY
L6Pnnwpl+sJ4Lsb1XH/F3/1SwJDWLqhcT9rjBljav5tOJelAQ7XLAs3BnmP1+4Rd
PRKIH+20AS3GeOUfjxp48uH67G5dbud652noWM4o2BtGu2CgUo/pTuZFnWxIblL0
dzQrP0UpnmG4HfdR2eGyk+eV+/XFbHbimg4I9bkVBqZ6YnwzPxzeqY0ns3y2Df1B
yu78ZUvXA0db9TWV8Kpumh7inXph7XqyF4khhF1VcnEiFDyMRwd6E13mHzWBYJMF
CB/8qSYFREfEGATb3N/9grJQVXYHMqpZqfaI5VOK1QPZ9xsWEkqv9DuAtD4AVyjH
DShRKQjY714K9M/04YWOEF1NYk4jxVCw2wCIZwSrFiutnY8pnbK4k204g/4ZxC0s
lubQBXD/HgbOWNPVNGV0A7JuFjFvU2IDS7fhA5HGD6D10regu5YAfIW1Ls4Q0Tkm
dJXxqeQqInimdiVDQSFQciYVvdaGIJjcBHi7e7GUw/NlJhKHgEIxsfvxJNzcqcKi
ea2RaJ4Bs7hI3TJdKE7ZsgpHyKSDwD9dAfFBxaXyPlqXo36jSkR5doVccAyd+DQv
/w5or8v5YH17qq37hdLECtuxkcMKftqBtAL3mqnPbrY2bLNjn+IuY9JR/LNyPqmH
sqqZoB+xxgxHUMt2ZDbCHjdCLjTdk5NN7oare3JhXzztvpA3gdwW8+b5G9goXDO1
vcB83xeHmMHDPYSHqTJrljaBl2S2YjQ64u7nknT/rnSlDsf/wICtUhNlG4lXKyAe
6mFqObvomD/cvyW6PnrmildP0aiIrQROB5DZygdNS6NhA3LdZBq/aiCc2VQcliM5
6wkvL6wFLOJwtkAY9U8Ec0LZ7TIBSLmQGmOnLl+IkxetPy+Ks7bzE+5KMdCSp0mq
bEjI0oKq1qENEA7seDKklj2bfh06R/krdXQTX8r3m1/sVU3/gcNE9RX9riPTWS+w
Z3ynTDkfL9PcQRvbwWMSo9sMuE56W0EBautxgUCfdEpvsNOG+OFd5gTo7qXuG/8b
sxQ3NI71p/4DrNiM2Gp3lvVtyVn0udLhc9LTYx0+G8UjymOSNY3flfBbXUmwBj57
P6wiv+EIhqq8+yaARftWVJaWSQoSuhgC7gEFOr4l7Fyb1qK2GvBd2MKX5uQcYTPX
EYib6v3AwvxYkk0cheysurKjxO+1hL3tFIclrLydhqM+9hhMQSvteVtM5+R3mYZj
ryF/7vL2YbM3Ei2yTWLDPAevV0lSP70fGaWTBLEDLFWGoQqMpVPacyxEBwWV8BAc
f+Q1yx/9R+l7pYJcotp57me/fopKbVraz3u70u2XLN0kCi/AyhPvoVWABlWr0EkR
Iua+s6sSI0jmswGWfgbi4ldO9k4I7bliZIlfPIgA4npdmnOFOKsSicp7z/zO8IPR
+kOTChWVA6b0JyewydNHeuudilQEWG6vV1B13ZQKRFx2aDiKBUzkAda3S1P/XCMg
0Pc8UhC/4Fm2mZjt8ejqOHpCGSQeGAd6bvvG5WiI75vK66AXtj/krJKRqSgnBP9e
DdtSR3xArH8yNQzwaLogTFWmb/ik5gpnZx/rMKpYYJnit9/ltXf3B3L2+wvOklbq
13dXs5UVWGGYEkSCNliXEHR5aTedXOfIoeMZNTBynboKEyulNHwwclqXvvxySwZQ
HEXBRW4ORUtFuuoTPu+Z/7R18zA6Rypje98jdiNqg+YJoi+3ex6ucqIOCA1n7En8
9rPbTUun3ond6q9whuzjLx7GKgsJRe9nCR9eNhXYzqiROLm4nYgQA+XTmE7+b24T
xtOv/UwWL4FWNHQ9pXVH9gwncPleixN7HI/HaTf+wKvBW4MInUrrt++hin7c4dus
QtRDCWCDTJunojAumH5j6oW16fIa+4Dr/PxiqUnYspi0QIsRd8jgJZTTep4LI5xg
RYH2Sjw/hsizocIkpyDXskfSsGgDQFlKCMozmeKjz+aCOUnMCkEG+aJ4DC4uxTNL
Afad4hjKfjJgQnJ+lq8gBzk48TQH8hDoyNdZcP2XxXcfe+2DeOKcSkwIxxGJ6wNf
NEiTHXRsPZYXB8qeMOfn/EOakLrBnRyJ2MGdD72MnfIl8FIXycqzZ9eWUTYPaEf+
XaIZ5gvmbj6oVd9NH63EALGnv2fWVvjxZOr1SHyXBdu+HNm4Nyk5CLun0WVxSq/p
4EBWveSd4AqCi356ysZxxwBxh5JiSa419xVhLxMqLyC/sHUx7axIHyNYOtL8gsuF
xwRPmk4pyb1XByLZbDDGH24FgCkp86/nQucMIs703SKAxKgxbxczQojwx6yNnbCL
O1zHDtZZtlr+CIgLwyNpCzSGnUPxCTHmizzC5XwPBcbbgknZn2jOyftacK4tegnz
ueeNMfzFmWUt1ppXidXLk2CDIjeupkNO0/SauWsuMAWMe/xzj/YOL9zZQN5sr8TG
yeAAO7wUi5GkBlw7jKxzMbDtZGHJiKYctzMBVRkBIe98j9gP8fo/f4vygm1ZNU4A
cvPlGrFEufV6whyjF2ABFtHxZrBycUbFWMHEbwhAV0b72yIzU47wCQLcQ1GcoEo3
m441MCR6lfn+1Fj8PwQcpDwlw7siAgbUFNd6dXXdrGCzkhToqIW+NLMlxb4vYACG
1iTMLkz6giiME5kfrfvnNIPYOdsHDkPmjA5R+Ds10zlWok2njOUXwnc32zsM+ing
LRLJSedJBDDIwzQNFMKn4pCHKWpejbYhKflU18Q+Ci1jLPSYdHuKBBh8h9OxVizl
DYony4n1CgIZdHhW19ECPDC11EnV/cRx0x+ubBmvMlB4jcoNx05SW9TyzQay50VM
OF/p6r1EgCL9cTsT87MMbbkxaW2o5QUkLLyMhpKj67dwVB6cp5JakRqTV7OIVhyv
FeDVvWN7u17UIYpibIOkJ0UOdZfPm1srXbscuyrEn2dpshq5JD6CnNR0ij99Od9o
Vt/zheZx+POu3QAwK9rXIQTqEKwP8pJhdJFF5v5SlL+S1a1OGvDnXVNpzzgY1xEV
NxKB7Ww0oikLvFJcJ/7KDAdkZPGynhOez4bIyPua9DsVLj4pz45LmV4+GDjST6t1
yZCR3RfvXVVj41Je+E7LkekRLBUl/7fCen+eHVqM8saET/vJdMsNJpLzm9cMEfuo
p/LcLvrAhL4atQFLRuyzrWAMUPRZ1BawMbR39VhOKWycjRwtpilI8EwZxPEPYlVt
hb5xZwlaMI+TrWi5vPcH9xdZseGls0SlPS5S4LTtRXdplNEUnPn9hl49jsHP/l01
I9Uu/tizPV1isO+1Tfbc8ALXM9UoHNgdNPCQ76D+dl/omtYD/RSy4ianCAU6P33p
UjVLFHI2NkrQYCVIsM1O3oxNkB/GzISBIcPntu1RrhpuFxD4qnyqo7QeA2cxXYCI
6GEz3rdiYCe2sTguOdaZ0eYIRtiJGo1/KgwEa6jIYLxpLKxVsEWseBUczXhv0KPA
mUe3dzDCHnr+K89fQVBNAfjTude9uWZNMwyFJJ4MS25FDdtSQgsFLFA1TAB5UFBd
1ulhoUhUjFI8UqWy4aR9RtngBcjsgtErDhAY97awCOU6dlbJ/AjmgnhaGXwOa4Q8
n9hL8aFVpIcP+QLxZpdOWvADe9FyK2Gmx/tlZCJvXOMx9R9h+0WZlHg5+mKXQVub
tmDF61BuHaTR0mA6Odv/AzhnZ3dxLctDIxpo0awudYuqopzutUzgsKiENRHxch9k
SfsLKi72bZs/fLNjU6ZaJko97hFcyuwCGXcfHqrpYW4vi4niQAeBObLwFzqR66Pz
5T4nkVL6GiVAxb2zz6D9dtA6/YAwjfOV+Y24u0OuswdTjlMjwr3edY8wMSVxBvRB
MXjDEog9OqsqajFNqbv6i94F/tsLkz8oTqaRrkC9XER22dURci69KtQ7aT8tEVX1
3tt9LbsSFOBgpngdV52foigxts9TyeWMSlmqyL1tQt/EaPfsb4dQSyFbb+bmB+WU
k+HE+NYcssAgfoZ308K7mXPmBHtu0jOafK2MaC67HnwkszdL6bzD3JY6aBrY4OFL
FbXl5kN71Cr/9zfRS7ent4az7JQ5NX9ZoFNFd9EOe2gRqPFFJGHEFM0mV5ug9qe9
hqLVHrdzXXoj6JdGA8lPf2urc5yAUKNleo+qvpQpQyIPvVXwhHMr17TgvxLzwmh2
KreE3puvSQFTz08FUn1hFrKMa5bJ5Wo6PrLbZut/k3yPTcpWqUEO0CU8DV9VeBnH
ECOxaHfRIqR23KOAVFz3tt6nn6xWhyi6u6W59FNGcQ3FCQ2DEPvuuAiCPiz1FQ9x
nQNxLng6HgrRKXlnev5IeCIQDkIwyudcwlKyiM87XDml5Fo9fHV8/OjfsHF3+d6V
febvHHgBYhxNxC/qCUAwC3RgHFMFHc2AkIIxo7zdd7vdL7cAjxTz7hCGepe6UnEB
3wn3lPZYhMMiDRZX1ZE7fsneYcz4yoxbgVrqq0CAA0uX9emuPZLGX1ScSNs5A4ee
nMhxVaHVVnUnnrqrNNBU7OojtycDtEkso/Nuu/9s1JURuNqoKbtLxq9Z26d1lRxT
6yFd6bLB7LXoSGTu177e043FL4MTQMkp96mMuT51mHgDUw7d1tiyQJd66stFsIza
JBSCsT9UoR9t7b0xUO2akhJqYiktsv9x0KRxtWfBtvpThNOKIvVUpqajRg1ctPhG
Hd6AzSyk21cEmp+VrjYgdPSne5Gw5++zud+NDrQ3YXoEPLU0ZVP8E8FrJUidl1VS
8lhQvi6eePJcwuXE0fyU/gqBNT0pmQy3iDHVtcVgUho58ITAMvoRZAOIqCughIZm
ih68hVW8y8tivS1HKOy/I39fpiRGHrcronTwF1gM/CpNWqfUPRKxcCzj4Xjv3qb/
eHEVr7RQe+9c5lXbySiyYwfmGDqUNCFr1LazUD41ngUwOAplSq5O0qNynCZyiXSY
gGkmdI3rW3pSPqYpYAaV5dQxtpi+OG8JZqOLrNd0Vzxer3obFB1VgtYP3/lVQ2Ro
Afhnr0oucoTGmvo8qGmUxYoyn8E9M+Ld+sA6Q6+xHOgL3vz6615t/KIewDPpxfDt
paBbLgZQu7gMilHoLh3PuagnCYPIRiqpFHARtZ4nRZrpdj2TBLKDpwCzUAghvl2m
G8YHO9hgi06MxpRIsbABAVv9tdYtUic/OKsqSEjcLSXQHzhdJ4PJlLAqfjmZL5NL
khf4dGBMlNl5DWNKSQsLcYmic8nqmcM7ETOdlcdyiWORjRCYfqODcBdswhmSR2Em
HSPfJleF3EM1QwNcAO7UEZ4oZGAYM07r6MywP9UG0dsPOkRQBewHQone2V4s9ctS
QR0j9Cx6Ccjpz47pbjNO23mICLyfhdvVeTurFs10cUZXFgap7Lq6K1HSkz+RijT4
NCx17x7Hfq81SirP0sGCTtJOslxtcdG3gcOFqbrEOFS+9QyHDHp4KhhTrtjfLmk4
8ivoqR8xalUhEthzeCQSkmwdBB9PL4CmIdeAaFICDPhVFnII5QjHiDtZBlfii5Jt
9COsP0K8kiX30MG0cR9IOvjab7qLYTPZuMJDgbTmk3/L6HIORs4z+cjX9VY+P/v9
iJ956Oi2N7xl4RxKoordbxWoYGUv5C/U09uwm+XrNXc+5kTBA4JHDQGnptPpM4CZ
mtQfXCoFMKdSIBhJSv925VKTE8yvLlyorfrdFj6vcZxhYLIgHDbFSGkf/QSkc4jM
CODVUt/ziCK6LiOqBm6f/z11I8t43UcPyqYTrW+fXn85XzTuhR1AKbmy7G7T4A8H
IQgPgULoCD/GrPWdslEdqdMnGBPwPh/GCBAkqqS2uejK5H87rCUXH2LWhvnNp/Ch
CW6YypUSsxHXtjAKQ0+R5ooeTwkRDBH84bvQr0Yu54T44Sw0ygy1vkw1oYOwOVW9
3EZSaNEaiGpUYoHSoT0HVsE64LfLuwc++PvWx2n2KMPN5XO2jAghLK7rJ6pOd3fb
VBuSAi1//rJO62KKM1dAmdEdonu+dJXpTIfirtxID/rNloDt1vBLT2PsraclQ4ln
7etnzwz1VwRcSMbarEUjOmEjZRN+5CYjs8bvWoHVkUEezmLNW1ZC21H20n4w2ZCF
581vkRL27gn5sSlDd7QMeOTAt/bYelGp72y9b3CynBXbc8EymHWe+7ZOJHfsLsxR
FM2PkGcTyyuwSk9nzMEjf3JgAwbF9qYRJ6MmGOqfvA/lNo53Z5beuqAcIFX7L375
VV6spkInM3AgTzXG8lCpdQ93g/YXWQI8DnFR4TkoUKV6v4fkvSqsFDPlSalyFaCL
sUcamDeFjkF96pPIKW4/Z1SrfBRtFKVq+NyZYmmcSqRmB2/tawa3z/cr00tPrCXs
TVJJ013R7tGHeo3rB8FdXxZ8gsJW83tBOnJYbqZI8Mxcp5rVP5WukXhF8KcrqqpQ
BMI5j+ER2Ko/lm40tR5bZx5oJbA0tEVxpElxtOFAwVdNSb7qI0UL7CXY9pnwaYfW
J4EdyNmkzbMQdxU6TmaNDbrJWgGBkEHh+25GEHPnp3gbW8zxOFMzzprPB7FkE+w5
2plfiEvQKDIveeP+jvxdswLPV/uFvpvXtkFfcyGZRhx6omsTc2Ze2ONrdL01Shm7
eW8dgU2/rE0jjTY4aEEriAQt6cBgi1wxzoJwfwHTGOwUQdAROUi5z/fRIqR+TGqS
K8euiscFKjzCS0Ic6IWxuadNaO7FIOBJ1tU8Q9FSCOB0iubLweU+bi88VJROlsXz
clhBlY8KoWAEY3UIuyK3FE59PA/XLoihQv7PMDYTqt2U467z3doljOgzYuqLVQDE
dKzTKwk8/BQYrZQeNVe0pKFzLoiKVvXdMog1YJ1YSx4K9WnHKL0DmR+GYOR4YyTU
jeCW/Vfzzv0Sm6kdPGdpWd0FC6LzKFp1eXxUOABL9UfBhv0p9o31RbYeP+DUQo4G
6YqcLwQe3RoxYcfEWSJkxKIZFHtXdUuBZLOCCQ+jT/Nkq5FzeMVix9Tsjc1zJ5Wg
5UHzRUF/SH4laHJmxi35Eltv7PFlG+V2oQRS4tTUJcM7+T0sJZj2yO41unt75twJ
+DlGUTppE+tDfSz1SNOKSTECD/hhylbYR+u+oRWFLhKE2hUjr6c+aDx4Fhe1y/SM
7QVJNB9rIKxM4QxjreR+EZySHHu9xtVW43pu2kaqiihD58a9pSk1yt9r7eO0jPIs
msEW4b/QJEUU5I2RVMIK/m3eiQElSqv3zCcXsPI6qXLAAYR0TCOR4t8TPpc1P+4l
PSaFy2RZg/Xgg2M/nLoGaH2HBxi/Ej0W5Zou6V8w568wz+ov9o+s62soD8MJQpTI
97akJia9fr3E232Dc1+EdrnO8EWTtq4H1IZtIy8CcVsPH1HKHLrcV/WwRf9017NL
0FHlyKtY4A8ldCTEf0LI3o+u7dbtsO/6kCAVStgaNMGtDTIR0BEddyrT/H4l4juT
fMfGXxzJifyUz43kiP40qN5SAmNFjvCChkLH28zXkUajs7XfMLGT4eBvOkoEMdtU
otM5+dCrr6r/Ec/MSdj+35FetDhrukZ7NLJixV6R2MB61ZFSBp7LrgKZVii3DAxN
eHPQF2YunOVmLykJTteScJzrPznSSLqzGJo0LC/uXBLYCI1oEVCLDuwCyljw+iqw
ffrna1mDGH+aWJOnbM0NwlLXU737E+Xhq7CSg+S6c4SUMfHwVBqxsLEk8ft14g49
S55Vg5ROQPaStp5kg5+I4uewoGNhJXelop4WAcpFqRTDChoPIfTFmbb+raml19iv
4HLUAZRYnRyrjr+Kpt387acJoykN/57n5oobD7xricG+VR1XSu9lIV2vDx+X9RoD
SIcLNaBu9LnF/1Oc8sLgQT8RGZJiata++HVmuzVT26QNlwVs63SSe7rvbgZGDezi
m75vmIo8zq7mZOBY1ynMFSWr+GNBEBtoqBajKytW7dW7rvHXP4R+AIfGwm6/thlq
R3+1RjPwaPg0xuNwGVVWzGvPb7hu6MbM3LzAdifFyFCB8HLn5UJzCZ0HLhar23xd
O+0GWrA4tI3YDHWRxyVoitI5Zvlq/Rmw/Vw4euu0ee9IrX14HHR2PmktplYDY95z
FKHPRhZZ1gcEYIr2EPzyTtKA9yXTt2pJxixjLXy11q0wOJcDuz6v/qDQBw24k+ZV
AAp2bzkf/BgtW0nKQ2vNKVp36om/4mcWdqDgMGw9I1/kNOUY9e1BnxruUlWIzU1l
y893Nbldnk8pe8D4hNFjIXqquRTg00UXV54I4StSLYsCZUzHIacfMti9S2ltKRyT
hgLjddmbiqleH5MyVJ6qfPdy6DaE7AvQf2Xo5i/EyMBAUaAM/HDbAq/YM/+azJde
FUiPoTQapb/WlsFSlthIcXj0+vs5ZyWnIl3m+KiPoILRkgVhBBU7pHt0PjgfOFrs
Iu1cUmzJLIe1j00zlmmAK9clkzd2FGy76gowjV4XpSjgJFmO3Yr8qDgu1yu7RdtO
6Ds79kT4fTiSine3NLQ1Hnqxbwe1eWIXfEQaJxmXC2u+qp4Vc0l6UIjCG7J4C9lo
LRhleDd4C6CN+NwR70o+T+R4v9thCKhvagiZGS6s17wfKhGJ1kO3Axy5TJWKsPQ5
BQrTM7l6XYcTle8KAUD1pZ1VnePo7d2iqMX7Goe0GXvZGEa8jWUNFoClqaBXRG0d
4EcCjqNgbvzdQ0/GQ18lZa4YBxcWVA8XPYL9JsLEMbSORkvc6weJJIX/IL8lJvRE
UUe1MdaaGiNmog2V6PQToxngt7csnlqeGGOvuvwZBGldBubKACTTWRKqszZHkurI
jJuVno8WaX7WoIBGrRrSLWFJC6/SF/jn5iAj/Rl0ysKpSZjeuBBNPCyQhl1U0N0e
Ne3/DCtk6YSZ9Zb8WEVYysX+gWTdHD9cbrQqbeigT3F+LUuS+/oA+ghZ+DFjpvmk
cSs78E+cTXyVaolrctckYJbBqlceEcE6smZsrPJvbg+jLB/+g/Oa+hPvvrhIJKKR
5dSnqFV1zg9mQOel7CC8QGHEEGgQH/EAdhVe7GHgV7KYb/7M4P3RVt+eHJr1jC4v
m2rTd7Y0U1OUu4oPWmDX3a7cHTugtrWJhjEIqA498p+WV2bHB9/8ZmCpJvFfrx3D
q+lacgd44K95oUzWWNbIEqv77vlcRt6FkHwzsEcvrdpJ3YNnYUr4MbOZN1bxWBnA
DZersiIuZH3RNgHzKg23O4kXNeKHzmcRuYZrqYtjmPlWbPtZRQFlbUB1LxyCYk9g
vd0rSUNEE5kbQaA3BjqnKTebRcIiTr20EYyrajtoSrIV7FNzzeJJbHt6IlYhki+x
6iDFm7elHFn+cqeUBPbLawHiBmYB/UxSc/hW+/LmqDak9gpeqVQZWbrVu+1IJftX
ABL0NlwiTs76fPt+YSptQkZu/nR37zhq1wfI08FTeZklQyK8HbNzslxjax0f2xE8
SLPgCn7yb/f/PuICELhJJqv9dhtLAe1EvEsCZYz3jmJKSZMu+R9OMfg7tqvlgt5I
naxX19zimawJSM/pQCEo8YEWUZGolr7hoVB6hn5+lq1/ZJ0nCDoVvonYkWp9gILJ
5mfMvO6haHgHHHYpVnuvRrjhDzg/TlsRykEf0TTS2hEmMObYrBIESFtP/yv29BNx
rE/4iQvr55ygbvRkm0obKCpGRN7yUSqcRsBRX2U1sJimetEw55EGpWAuUm6FEhQv
Ent1RdJaOq4FitJvtxZ10Pi4ht2NBc7cbCp/JS6yufl8G7q+jIEBV8ba/qg4phYT
wYrCp/TLTtM0F6M65Ao2XLH9IqnZ4Q24nrgvsZYDx/Gkf7sQz0uKXUbF/0QKQUqA
1tAaLKbjJd6jITDsUEto62wF/VkTuK1JitIiSBF1FK0WfHdoj99xH8SN7y6tBFFn
+G4RqylUXKGVmTVKu30LvsM4RBq6yV+9IhKjDFs5CXI3qJJC4qXWyPxM9ap4I2vJ
iyg4Jj37kcUNX70kATjiJnYjGGQ2f+hGjaUA85W4dMqTjPqmyvKxgLelYXsvw2nD
5YNklF24qPcLwrXH22VlIg7Hnrh4sXPFPH3BRVtZrSggqDxLch89cPJYaQGl214h
tQgrv3wAsaQBLyFrwCpSGpGJOfsmsgUvBJWdu8nq5lPsnpYms5xyEnkYW31uXIhs
EK3aRRJCLc/o4eXQB4R77WVhEDk8Tsj4TV6ItJw454ibBMqRRWswTmlx/kbqCkCn
s0Cz5mmm7UeAVBneCUFf5mQ8y1Ffq6K1fQ0dYxLr3kBqClxQr16F46WdDQwt5kFy
gtUgt5yWmbueW0R4DWRx/0sX47ngDCBTaZHso9JYTBtvcytyTmYiMA4FhOoZS0a4
js2YUjBKbDf+03/SujiEA6lJqEcn+ZoewhOREsVgNi2BBgoJ40lPiS5qpWA4tCgi
pypgJppWLmFrmIvFnYgrp9Aor65k5VREGHpDEFjoiLDUX+G7VSleK0huPpRMNnfc
MaqFAjxgUqhqhNfzf0HOlMi2nr299FOdT5oO9j35+GpiXw7WB6StDqE4J47+Iepf
PlZA+vwZ6J3ICZuU7spb+pPAYXiWw/7GaYrFF2KM2anC/Sr5QJmgT1EQj3Wn70NB
ayv+4WudrisYEssMpquvsVSdp0uNWqu9hseKq78AvBmRqtyRdWYnW7/ZFmYBB2Hp
5E8bGUhc7tOpzdj1csYHhVkVEnSJxpUS8N5+P16Q/ITYq4huvYOycmFsFQkgVxUS
LfRp/L6RosrKktwchWeFK/pHwxiFsE1Nmo/apMT6G132TN9SGCWH+AoJlqkEScJD
ERvyuuWDc3+eX2guxWZ0tBsv4AHmPosAoSk7tPBUgHjrY/c5Rl707sZAIf1Hrpnr
oxh+QayVJsVnVyxJoGrpvQbSOR56gDC5mPosb79oKwTJo4p9pHF5egcOVBz0J5Nn
ia1NS9HSxIaJf5/H16jDkXDR8qz1Om1cpkhMrE95V9r7qM33zEOE2Ddm6a5uyI5v
IXSHyb2snkZG1rlS6oN7PrTal/S4xw4L4ZKmGWwpEFdqlDuZDaZkHGhkIp2KTVE2
M5WHCRDOiiOzTLHco4SSnUsY6CwRDoWV9hpTs5bR4u9f35/7dDFhp+Zc15ACYMZa
jvyS/MbJBYH3KVlwwVsKbCgNxKKuRCyN6PAFhyPXgrgE/JvGg44QLYwzhurEerkT
6EswKlq1wFvpHpnAQm+AWTWF98AIHHVjvfJimpf34L1iGM9JOrCdvUwBq88J3hl7
+e0oqbUXzwZb+STBcmu5GWtY3eNVubHuvxLoQQxx1V8r/75qBnI24F4wNPe357z4
PdRC5uEeg5f4jkdXDTSPIvKBA0vdgj/Z9QxbhnelChl4AlRvzEwQxL9L1B6rOjcf
pQqk0ru0sfW2I+ITWI+XTiMV+PNhqx7CQUwbRLi2u3kZ9qd50nJKyiojGCV+fG5w
5b1DNLB19k8+ZRpFhLHW0rGmKIFDuoARghf53NzDKm1VJaVRrUTNJIn3WaUA48pS
3pHhCEei/2CUd5/cflkkVT17SlmnYok/LwOdWHP1Wp/L86edgqs0erhvp1mGWrZf
qxgbI+O/fzc+eDsHJiofVtuhs/RjUaNOF7N7Bjw12tUszX0JhavH5eETxYqTW/5p
2HjTycj3e/6Bx/Jheo/o8vLSlSEZGMJQC9GETPmL70WlooGxOXYseCavLlMRc9y6
wpzfyrEsjZloGNmYrmeNz5idhmaX28Ruk1eEQ9SlkYPzlz8B1YxeV4MgKPfA2wwe
EKN7k7xjWKzvKFEuBdA1OLPZSzSeXXDwkbjufQKodNUAII059agJJAKGhjMyfPHU
tBQ4yyLMH33hTaPhOgu3wZMN69w3Ij9LAzDwJZAQlg+w7dZqwk1g0MwV2AL7vQuR
R72x8wrIeKpgQ4XquEUeRGxRHrykDI5RgJPD0+bR8XCHJwnRim6cU30irMOTPzUQ
bUGcaOZhRq66GaKJBMxCkK/dsCDo3MNeERoYnYzQKrXFFnHM2lXKAhxP3AANEXNH
fA9LjZJ+FPKZ3bomgz1wt8QwIyAvCf1zOOh2hg1qgGJbKMAHPuAKMSiWEbeQsWfQ
OcjGvvSfJUNVO3mhc7gLq647qXbI0SJ1SGZw45oCVhI9X0Uzh21m1lLt5DQQIfjY
1kzjozoK2AC4Q/jXm7EC+aqg/jThV40MgZncU9PgWQI4aMff4TmvlC+b0qanoPWY
Ov7mlSdjXqUXVSet1X5sp/GXEL0KzUvEi11VnOQnxxIaTzSUUtJR/eU3EFr1nS3K
megyQUxOEdJGBPPtOVKcDSMDjiOqMg2z7cJulNUzCcQWkTVIPzdV0jIWOzoBMssi
pfhnLacBadzQxCFGZLLgy/Vp12VY/4/hjmV0caXrXlGCPkcxWbbOQZGcThkBPRUQ
6Ax/GvZ9QBLDwRVZstPlGd/K3WL7Ga//mnwHWXeu6lVUCxgSjtUpzSNaQCSs5iw9
4wy4Ll+4z1Mgw1NDQmQJcrUzGi6Gng/QTy27EviDueB6k0hpJ3IGUnB1PbE4VgYa
PvhpnESylMQ6LRcqr5xh6iFoZKwV0PvP6G7sYXGquJOuhRFEEmRbF4sR2pvE4M1l
LtDlxrpVW6sabFaG/ERPrM3Qk6JTs9U9yKKnxegOJO3UVzXrlJAYGXy+CNisDudE
cKHhz1ijE1cIQAxOVfQvHY2hDH0w3Y8/vxaWF9741fDlAlJJ2MJNc+9dwg2CSbj4
5lpEmtINbYP+BnvGAnjKCp6AlUwnwpEb8Q0SiowOSCy+lbHofcB9Gp8cV7b0XXtm
x65g42ezNxXz65M0vkDNtwplwFAIAd+S11nFwWTkl/Lp28nCmDV/6GbHwuO+AWdf
Kfnpq7vBm8DygV4DgQ7JUl5SKHh+zGB2jNpCSsHbxlHX10Qn63W0PutOpVSsnCG6
81ahWh+Gh5hDc1Hl+hEfdVi3wsFV62eYElCgy8OJpPwBS631nLvG8CZ0osAs2B9m
U1WTaSBVsUz/eUJ8T8yF9Z/laaO8efKHYWILGHSIC0ACBb3hKhqQ2J8rqEkv161T
W4oEiMAQXwmXgaP0OTHa1DPQwPcPNVB3ibNUkXwGThK8C/qeEuOjQWQgHh3hYrPD
OV2MWLYHu27KrPDFPBHNB2EL/PytQfTuNroATlD+nh+LbLGVAzUU7+kY8slVyipr
jUJSOv9qzrH2tEfb3pQwqwF7RWYCJNy7zF2fFyL/L0SBNfJD+AFlGlshmwtRY4cq
eNAxlhETAv+hItrwHWUtmMYAmqYb1sET9wsa/G1/UYiH48RjC4fehqvU/fC0XDfg
RIMhhi2STCcGvSYc+iHHnMrgorJ/fV++eNPuX2slpVo9GpIrLkbAS+q688JY383V
gcZcUY9+v4/8sL4MUU8qS9QD9CiX8Rn3g0FbMKfLoxpbZTJ6g2uwGAZ+A7AG4Mid
GNjg+tTvNXlA/v6wBIGs3T2NpAyLSiNPEJ48SzS/Mg3cbbqa7ZTQD157dU1jYKEn
q0FOmJh89bUNYuE76BPn+k+Cyy6UFoePnkMYkZImHjte+7pZ5F5tAdjPHeVxcf2e
P5MGs/+yKvVYDICT3Xg1/gjlhRAf+iZMngP/yAFd19pcEY4dvRbj2fFIsH9oIzY8
Dkp4eDxOUI7SDr82zLDfYH5uRCNB65tAuej+2sJV87tnSRVU602qRBNGCpRTDkk1
BU689BR+4AdntJHiEXwAIQ3L+JumiZvNHN3cfE4S4cpLJKHW7f1A8SYFy3wuZkoQ
VUPioEWc+K4S97SxdY7VEn/TPv0ceDICrb37dzBM7t6ef0tYgJb+v4t6qflj1CZo
RBdR5H9Du4Ua30y3fvpCQ9ZesPzp50cIoGhdYmskBBNhsVhBcmKy0BaaHApV/JB8
R9vmLHSAcIe9ChmiEKOCw97Y2NfZ/eX332ALrT7fVpHivGsA9mMWBYJzZREtMGli
z4z+Vz+okh582HzZPRVUpq693MbYrFYuvkGjspIQNaIP0gmUdgYki75QLhrzOw+0
Jwdneepk0Cjo5I6xC9N1q+jBASSPEIwNbco7GJzHbCfoExJZnX4BIAu++ZOGvayQ
4jgElEYfae9T1dzcVylgq4NBZds1L/ABfVmvrTN7YE2H8u4mo8EcV99ljhCf9rlZ
L2B0wpD1kmT/+0HttQhDKDc1haaWU6GnLYIibhHm9ryydN+S9ntYwt9y75HlKkWv
zeh/tgCW/RpvjQdWuI4VwYemMV3f4G2+Pm8njRojPgAlVDSKfUJa05+or7Mxg6Rs
CD0cEKcaH449A88kx9NDPQY54ltFLMBRf9N7hgq5oOMSyZ9ROx5aFn2q5PiBTbow
aj1pphGy2FaDMiZi5doHpt4Y0JRnDXKUoPZOKgRbsG6JDNxgtYMtYdllbsGKyuil
XB6KbZCqjyUCNQocS6dVugNsakYOUPC8mten6APKajc9WZKmmC1OQDuS5EkpGi0M
bOrj/Hp+vr+RKcHjIoE/BDNuOR9qUIdjWUSEDl2tzWUt3kkLKaLb4CqJoLTiACWk
FD/4YVyMhIAW3R0MrtOFSKDJB6Q2yCRQmtX5HmEIk+2yH1W0dlLqjAmHDMQS2U39
IR1nr2vU1rH0FQqXuX6szdjtfSAn7oV4/pMmzixypMFuXAMsI4LNsWHBuh5msM0z
gjHYgAirUtbNiYVMzJjbOhC8huJMlrbbUWwhVGpzasllWN9VCNfTsy8+ROPwND4v
8X2ag/6FovOpG9K38utsEzngZm109U8E60j16g55wz23QMDNViZAxXBmJvDXzuM1
sSotNaDXlliNh5H8yq8aruF8T7ox4mu2pVUKAZvhqfQyDKmsMNPYdJMuSsf3YwjF
5OkchyWintuBs9J3MoaNFOTHkyCOemzQtDnSjMZSyM4csWRwTIrYaJ97nde2e2ss
9bZ0wjty67sVnzisNlfkdlE0QRvjoPJdus291KEJufYRpcw3RT74sfoC4NW8SXeO
qkDlRbVc0+g/LG10RPywZ+tCYQPAca+DaFMCtCVkz04h+pgoQezY9fRLPpv52xIQ
VZK6Scj4SFyNrvvV/swEP0TYWRm5b1Un1FSvrvzd1Xw4xiLLda/iq/IXza+/EZ9J
9f1W2l5SJsBqNvBa+a5rt8yxhWu8fziMnWTVVxJ0RuyQ04nqMspv+qEZ4imCh7iQ
8U3Etgvc8+cg1i6mGZTCMR0KCizaFEjSsNJkmtvYJVJDWiON8/rPiHQzJGDU6FVe
8RIvNiqtLGqUza6PukAtkvvOnNZYbdd4iGByCmPDDmgtcj5uDqKcMkeuIx5EbCwh
ud+VRjLeegyfMe29+5LADzFbH9c5mFsIJauTNOn1pLC3QWufXmJt6D4mWXkla3xN
JP1mrWPIaYqZ5ydw+TAWSaPh3nyLYUrQf9gOzk/RDO2jcJIkGAmtfilnVN5Y7ukM
ukPWZHa/cki1GD9xSRCCekdWL+UhzPuENafWGedQzvVWOscvxIDArnvGNm8IrDHM
cMFIxbjnjPO75Fcvzj/rn20uY4P9u4yZuL2ut+AFAIUGPBw3CjMrHHrL7R8poy9e
sFj4siZHz/WELMjhETSYoElmZvyjwYdpiKMg7Nb/MSNG1UL/yQoh7aHhrzryE04D
B0S5RWyUR6qF1a6pLkCsZqqhgR0cdKoZgE/QZQ/JQB4WFj6fqj+mjaq9aImMfE5o
WD0KwGt26B5Vqzt2UMEXnJjoaH0/qZOEpdr2317nLQdln2PlTpE1znW8GYYQtLqt
W5aohvPYvrLfhgRzafOxnajEUdtc4NmPZqwJf1FzVSAgFuAGM3d3XAd9SPH38lZx
USppY2XlxgFDzcQMflKJzdNFkQj/jwto3FgmHiWnI4haaeHfzBEvXgEbxMeYx4ZP
xfekiQSn13ihAUtPOB4iio/y4igZAvMlHTjI3wrJSSKhCgg4hTjp0L26FCqD3LPq
GHmWbJ8qvJrwYiKEtPCTqcCBvnMiZYQ7AFWT91NqXgBvHbHido3ivhrmD7CT2bIj
QgFJVREBLoVFqf/CNH5gCjPRmYx0gqL9SR59RxqLr9ojFGcoa3qi5oUw3qu8UKD9
uKXcjXcaDC9NhJuD/MuygfHPpKyqjj6ZU8RcL11KHknuNbqN8xlwSat+/+yXAig3
2bKEH1nqootsgMx7C+6kzlfi3zd4HkiVdlsB0aRVFuFsP9Z1+X2XHOJFT7JP5Kz5
BvbxAvzvw/iMnzhxPlK6ad3EPDI5qXAsAR4XtJIRIoZaZEceZlTqtmtfbs5CrzdV
PerCe8sfFopPRHcYqZFE5w3/SAKdXsBi4whrqDKwy/pwiGORNMfB3f84b9HtIzbw
noPdqhMlxc3anl7mFTKRJeJ3WwbogMUF3mIboUmKA5yytJ4Az+1rZUVwz5jm337v
BeqMo3Uw5b5DxyXSX6Rz+fvGXFLhcy2/H+lSXmZkYru5bkfg2E9UV2rFjOik+3Fq
XHZhAZHRKV7eoZDD2lt/eG17a1IHoHHOmdtlPpS1+yS4Va67mSRdm2ulghvfPbQD
Oop9Ks6ymxiIQIQeAnxBK608K+p3cs+KxsAXcwXt7SuSpOpYS4E6lppbocCqVvD4
eryKOZXyPNgyWvXysl4QlUoujo/HJ6ozzzXIacH8yXXkEcwPD+/nhmm+g1YiqkXZ
8aU1Q4MVY/3LgD/oC71gknHSdhFlYc9lZeD39tEGsLflvkljvcTaCcBqXAZn297V
CHX3XkVXXkmudpsIKjQPC1DQFjkQaWx3PnXEFdcohJ5RUxGg3S2djrqRVAmgCDp9
0OR1LN4+IQP4fL+pQulCL2unUccUPpOGJpTDRgJdhwzphA4Ke2F/CsrD+UKnyC/m
Z9oUy1PdZDYO8DKmVgRDCLaRM7oQSY/UdlATPS8gUuYcH5WstjJ5D9Tn3Wb8oEER
TlOqxlv8OprEVtWtSwpJeU6Ok84RLQhSvoWNk8xvrRNIt6zM9AMeYuq4SKITxy1H
NmlhAUhJb3TjzxYoaYrrasP8awXNADDV4UwkLNH7FeT0ZcIuj0d6kMK2lzs5cROH
Qj89XzSR4s1zk07V5vP8s6VAh2oWupYF608IUV4b5VGei67TYG9ytqYKhtGmoOq/
1HnjHVF+LRQDmakR6iSdL5oEcfmgZd824NIo4otIBMqW8P5W4tN1Izggvfr2OZ0C
FXF/5wcy/9IgtSsP1s/6A75HujIA0REGL3Jqd/Q2KbsC6uCGhs8pHdb5gOf9UvrJ
U1L3DJrlADeXAyuqcR6S1C+HxdWsT2ZMjrWIe8AbPeqshIOgjmPHLeF1T3zyq0RO
6IUFHiXW4dBmV+Gd4A8rS0/XeXqAHOCtKBLW29BTYM9ABctEofRudJp/yWsUUJoa
aqCTEJ9LBQ9fuIhogXV5EGzQ+iplTY0P09L3KBsJzucffndaNthIW3D4Zgw2HFPr
k4ko9R87bMmaoTUmdnYvQBLKhUaCOxb7iMu/Cwqij4Bqqp4x9+QGOHfjnyTP5frU
qtYFKyQj8y5wL1q2Gi5DNjpPR/K8+Rx00X82iPPrc91d3dVKbtjXti9VSkg/UeO8
Cy42jZ4Tb1uvdJRZIgEkUO8l7J4rerIYjOltmAxLlS+MuGGp15MAxBCIRNVg9mn4
+de1tqFq+l63W5wzb3KDxD/6n6uowWuzQabaSB+7hD1HMkXAV/BIik+KxecmZgwc
wV31hj6d+I9iWDf0SUW2XLpXu+hj683H+pfNnxeoMpOCSXgBx7XRuJhJf4djHv0V
xMaC/PNV6so9Xhwt2frgKuRgOvoTQnEt5s0h3k0JOgkviEx7t0Xs9woAEyBHangS
PI3Bjue77MYP+MzZxAT0yZ2fYgmSBZ/bAiA5HSz1QsbWJkWOrqwo91lmusMDZdWl
Z1WHuj1kJhyLk3f3GoX8Wwu9+w3tvsmkk3LjftuwPhtb9F/hZDPOSPGz5aviTNZl
2yOhMagiYswvu1LpgYPXHmm224mRPnIImC/ztFgCGMtwhCU8TFl8NxGTBLNyLrSF
DHnAWMqDmRSPNkxE6xCKcNiogEH+nAFZzadJWJvUXNlSP3tgAlk3O5MMyEyN59R5
WgQoUUxohoKOBaqg/OhC0mm9wniJddtQWkPQHJQ3EM7ZySvz2f/0MlFvRWDaqMhZ
K+JpJ7hGzvDTpa90e8PdI20DSmvOp8n/NChuwERJbwjJpHoGe+HnwjsCYadp9qe+
5X/CfX3MXPH6pFG+TZov7E31KPcIx7Uthz5Z6GwOvLoVaRv7+bdShY1QR0HJWO8u
Iu0nuFamRro9TovonFJvXa8RtwhcgVNpRnVtr/Org7MZ5bZn0njxhW5J5jziPaNc
H09e3xwCDU05Qvm8v/1Gl4dZ/GlaDZApQ51KHamcUE3MTOX8oFbtl7/8XJoTYCPD
2h8NkDss38W/6CM5ToRgcBJ+84YdgtergdstZsoal6uNVr8abRjO6ZCMQCdBoIgU
sr3eF8TVuL3Fif3T9wBAQ76gpAoJT9ULSqIFbttvVPxekyx0ZrOnDbmGsV8mPotn
me57ojFRRrlupr8KSc+P8L0aLZwk+ogtiSwxVoz8ZJlk1HPNF85w88xfAzSr0UX4
7Uk58/mngCNLKG9XwoEpUoYzaA9KtIHfyaZ53a6iLbpn30kQsMNp3X0ieIk4Nftq
oiJyp9O2RKFF/whjutnTSV9HDHVBCzwECb8qITHKMukT+CRE2Q4D4DXCh3n5F6BC
hptmVSKBujbaYUPMux0TwwsSGZRNRZTM41lg6ATFZtAxCfIu2/7oty7l/SrtjgF/
hgPk/Zqc5sD4rFuywaGsuk/za1Hm4OLSHO1WX9RACE5bVj971rFphkULNESEkQkK
AWi2stF4IFw1qpPFVCRPjw5vn4Ih32bmtf5CBc2zJveQbzviGCI0HWHy1HHTM93g
kGgvBVk65EMfnXsht2GyFmX9UhJjtVWlBwRenowZiKFTx41ofvYJQ8F1ia2+RUKv
xNRPoqltnPnh4WTr8nsN8jVXgPTqq0uwMQd/go5mLwZS21b2+HFhye1YapF9cxB5
Oezem5xnuY8KYxdT8fXxEpjMdXLPhecBDYHprVoMTSrKQ/OhmNaI4csIikaW9r8k
pMDyeX1ybujG8qT0F5qAIV+uvrLQOl0Ef0n6BSwUtuiWA20kCTUrY/Oe8V5gz71a
PNdpwhPBzByQpWot8Vw7g0RvCo0WVPhDD9Jhky46wsnWGE5nZlxQqMcvdr5Ml4wX
wxuRW+wQCEaWbNYflWo39w9ualSeNZLY5VSWqLeR31ZIOqY8vHeiQOwnDTVbZT0a
bK1lOa5rNGWjukcWtq33rvw+6oKuV0AKzka4V0erUnBAXOWi4R33UkYzsnkbdkC4
6SvvlqawPRl3kAAPC3fbQFOQj5ZoALdjai9JBVnAOU8X0pTKAa+8ZZpKZDKgz4fG
/wbOxEvbsmTwxxL0/EyU2+p0heVKOAbTg+9K5LQlqhIAtVR8KnqtjAe2ZerFyYbV
En6rdZDtDfSbrygZdlVCjpIH/pWB9/Osb2AJdf5yeuAN045QW8pBt+f1o3fpD+Ov
y1YWoC8RIiLNfIfKe0HA27XD1FRWlRhuxkOlVSswsQ0FV/iWnO8y6pTwGfkYsU3R
4qhts8eX6Bjl7n5uqMI2Yhqcq5BS7kUE7ibmQc5V2PuDi3mxQ9Y2m/h+OU/2vTDr
J5bdOBkY31ZzZuAaR2T/xURFAVdb3YGPvy+dvS73So30IrPPCSvkgPxzpQw8nGVS
7IseC/5etSeDM3Psg/WKQvkrDw6gF0VW8tEMFU+Il/woEy3cXIfMRpIR/+XK9LOb
zYguidgu9IH9kt8C1WL12xjYV5myTBvEjeyBNw++LZ9fprbxtqrBT4TXPVz4DbO3
szsSM2b8DgJ1PWXZVXKUcfH/ouPeEjAoMz6QxumrELONUkhByk1SB0gvW3rORL5P
NW9SgNRJS14SabWHYTq7NiwifhJvsd2YmxFgR0wVBt2dlkE7WK+Jc5uVr4qIygJe
z05ciYOasZPNN31lhuu0rWcJvT6TxKhpr4eXCg5is4bu6XFuENmqtLvYigjfKBmT
UyW/PCeqonsiAwieLAZCMLL9g0rmguiO2gOcpUNpgPuoLZb/pxJAL6qORF2uIFZo
7vBPxbBWgaCM4VzKwPO3++t6Sg2B+7PYc/PUSI6QO/Jcl+z+pMocJz47wAnLLcwD
ih6LkJHGQltmNsy42qKozMvt78WPrWWfjnLkjSv+DRy0cN7yOwnWpEbObRBQJ9D5
KsO5nfn36mk5Mo64djkCZcYe3bKJZ14vBL+/1RK8DI5kYCxn0AtxOmQEtDDZDW+X
HLSCCEiVokyNrMV9N7msUmARaGMfPF/yN0QaqLE0db13ICHCMyxEoK2KNzP+Rahr
/NIfyUZxdDVeaaWlcUZDM20UegLj0XExIKMeeB1BDaI3KOxuU/loTIsqTCamHAte
iutHv5Ezv6Swtl2iPsfcCpPhfkSIHm5DBoBA7OMUFwjgvJqAfY5iXzRtrCMJYolO
b0VryWF/4XRfcDXLSz99T2TmzLo/ouxGZgScyTF0Am6+8Ek8JuEpMggjUP0WXrcN
99GUGeEfE0/t9V+V/dV04bMi3BSaqY6Up4yDmKK4zjsahxcCuhYhcJVGZ2c8Hmug
0frCjwLiv8Su4o5Zfc+SE3HI4tvwRFEv6P6rNcI6q6Ci0G9fkGI1BFqYQKEMhITx
+zKBOBZe6jGMIqjatC72Wr+7AwCZxYbvBSk4t84atpa46+urtDnL9rPiuZpqXvsa
SHzoeoXQTWf1Lpa54AfHYPvK4MP84R7s9nupHZjCeIjVsJcGC/9ZXj/P5NRRe4hA
cLOE86OGUW6NEZi4b15IlP3cuLTpURfkXXG4zTRQ4qGoJykeqwnH2liPlDQSLe8P
TmSixXL8AgOTlRcc9o9rN6zsVAC7eREEJepiS+0IXEay8GYWLJDOdUBei7pbtgic
oPP5xiFM3ET5Ztmb6CZJsIvUBsqnYFhTtd/tu592UDTwLehWeBT3hR2NysHVUzIr
CvSkiNs2ACGZLvONqXfFKFKTSFRYOpbVsiVQJuWYgrFLGH8EpFk/iA9HJ77fYiWt
asqiU3y5xpYcqgATwk23kKMguvRUXv9MYamU/Uz/VpaheM6IX9MYOca0edACtnlN
v7jsjcsusbwy8FbCb0tzQEV8dO/npIYAJWh/8RIolsyDsZ5JbLODne/Iu00quNo8
NY9Rw814CPk3SqnzSf9JQFSF5EJM1FH4M7uPG27ZwjUHDpfJqnJrmmREgtwSmjTj
NqYdKwYcDXL2c+sbh5iYK0MakqoGjKmPMpV9IJoaxkdTa5E7rwBJUUie7AJzwJXv
fZYmZisyKbb0VSjo2u+9EM7pQHv4QqhndJ095b4H1Nnauj5W59TpaX3d0OuAk9XK
Sg+6MoN8L/ZBvs8d+kRgftsxzHvsyI4lKVGLceItsSLm0By4wckGLdyNxLXIPygP
u3D5TotjD9HjaYn0FWRAmKf8Sj6ShyleFHbO7evU9+9f4xTLd0QFj/oajfCnRRqv
zyVkq7LF9fod1QeI+f86vrbE4ybMGLBEoh+QlX8sM7Cga6YYazRZkPLCtvxgIEn8
RSUtTQYlTkP7Q4yeBe273qljHoVJtt5ejLXFHFGZqnUXQtUZuAPsN63trx4mDIMj
h+ZnFpKYUd0ArqB1LeZMFbTrXhoIEkt7GPVtJNH/XHdRmEz3VkJYQEdtW6Bqr3oF
bLfIXWjznf30Zqz9rGi1YsWhEZ5vC8hL5KHHqoSJRcBY0B292Ql4Jz6JjzEkYIXc
D0z9Yhf2ayFVzciKUwzyPqh6sKybuF04yG+qXx0wy7BLwXYV2RCJArshlYXMK/qT
EZgR7dlv7p9QueQRciU9Q+sdWsoNi8o6TxzwAYqQ//GD5oOaLbYNcF1WA4WRn9/V
WhFHtu3VIGhrh0i6mzj5bDfkI/ihrlf/4Bg5tk5jUHIpK49iXcjDXWp+U/BtXdnk
sUxF06NMbgw7NhuDMW/KCulTl5rNGwzA3DHZ3d0xFyRa8L1UxWM3hk9k/wDlFFLj
VidfXt8o5EgsvBfGcjfciiZjnN9gqfjIi7k4e1ip4RHVSWtS1sAm3SQcDXz546us
ZIbwvfJqVWRonApvYOvQkZjK6AeZPZ73th73FkVKPKlgTCe3ZeBKOLMuYEWNxqn2
mnpu/9C1Ft2cpzyDzRUsc21mXRGJl9FtFz2eIX18dC0c8/Xz2A7WujtWEdSq7dxI
yztEK5XG1EDTbI9fT7nujgvvxW6ARO5ChFRdRIAcxWM3UZTOM69aqjA08ZZCosiV
/4+SIZixjqBP3cd6JmyB+eTnFt3hUELXfnR5EWx+L/Oll3eBXCFAJa/8XYDSXEHL
34Zi38nPIvEXfQ7dkVSajiC5wDMYsEUgh1DXM+DNIzV5xPwwKxJpnaoQNc1aqhKH
oaCFVh3pWwK/CGBOlMSKMnzxko667UvuQm8wB7oj2hZ39p5ZStMoY54ljq46+0+Z
QwB81SSy5MdIOcLFqE6uzA+i7n7lvpJLCHUWv2RII9cxFAjqXoEUUdehyNmOWW2G
T4sQyOGN0revjRX9gTJ9AW91wItD57CoiWjssUOd125+uf0VU+Syu9C4nn5PjCc7
GqEHXOQUV3UMf6JK5Yh8W36pEhyJ2IiDd4ObGsXfZn/86Z6qPdbWfXzI7tjsmfqQ
BgSh835Ds3eFXBbIf1ze/cqOzzGf4y+w3JhhuYc32q06VCm1szo2ZvzMcL4qnQ1m
icNId3VVojvEYyDHveKHZHOX9FGemU2lP9dyuJso+b/pMZ5CxCo+Ob5BkUKdDUC7
SfRUIi5nOFhPB3YaV5QZ4eM0lAOT/wfnMb9wQQ+cX9hcuFBVxg+7JMlIWm8sJIhf
7TIbN5ZqzpVgfJr4NTz6ko5StJdUh9+5DEvd3DDpPtNREMVGOTMsHN+mKgJ40sRV
w0ezYSxANKqfBLM6Yavx7AcQ4P8aA1yytFqkqU5UR+z+qNhuWAaaq7ir34+aQ2U0
4cxXmOnP8viB1ZMUqsIxgVr2pWV3unZ9BfGzKe4fJQy2KjK03YEBrUnDOsYbTMl5
dUDqIzFZzsYPIYarceHFv04fwHS44tWLct9T7mY+Fo99XnuwykM539P9RGEO+ktE
DVG9yZIqVbwRWesO0M/gkj5kvpbAXQuc6IyeTc47WqqtTPNO7HhoShpqXirCjck3
pPJgZcAoDaLKi7nYwyX0T4EKtFvBiQB1TXihDexDmlacDcPk8ZbNcz4E2ZTSH0eO
bLW00jVybQtPgdPbAYr4IpKQMOyuN1VQArHoZmGorLj3eSrjM7YJ1nMZymNB3VW/
rdVyFkJX0UEZjgirVTe0vdvF2YNQAkEKiE84DQJSjKFUuzkmip3wis4HxP8j/s7J
x6xoU1o2NgtOjDT9f/TalFRxg4tbV+rLHpEz+rgySUx7x1ZSO10VtpL44iCkLsjU
bfknqt/VXN++NGmIfyOZVlPhnG+3T9zPjf7drQ9PaGssPHotLcAQuJFIB15tEeuF
XbIGrd7JF/zKN2/Fz4L3Nzv2KyQEabFEsib05K056rwoyZGUNhA+NQLN4iYhRzQ/
eJd7p/ETaNCPivEk6z8dXLdrjtEx0HSMjRgTlQNTVqFXNm72A6zPO7OFv6Wp05vi
KPSn/fwI4Gj2RHPba0E7AQ76dv0tTvEvKp1dazMj4OcDX882JU6jJpUhOPzrbqgG
KoLziGnnmZZYNcQH9hNpHJ13uUQ+nGAQanpnf76yzr+FbmDXLTt34oqpDTUdhi7S
HwNtCS129NnjLR0y1rjmIE4uuP+zWyf/KyWmeWfA9ZFjPFcOtmckNEQNaDqQRdEt
ANopiKl5V/iZ6hNaumUgKJUeQy9TCSGU+ILD96mPiJLRcknC1/AEsTDJ6HGK2ZET
P+4/9YV5vAIiPeWLFrZkScgr33KeSbBDJBF/qEVdOEbNAGWDwLEH3VIn6JnlZIUV
uVvnCK4U8d484TmzFT8zGDIewF7NGl4ShLGvswE1NvW47nlQq0uYGbQ3URyYBXhz
RU/kdZZqZvve7D5QYd3AueQ648KqdGeQwpNnb0O84Cl7U84fCxetukWwZWUCDbX+
Ofjfh/r9J2c45LfT1e09t8mDCiduEMyZYdXMWYasq0ZxMlxgaasfYeT8SRddFvRb
EI2J+3Cz6JYVp637muCXP/dfBeAeg/vHSeaT8yI+kZwyC4euvhWV7ft4Hds/VGeT
5n5pjHTQElP7MWUtmJ1AHdDxmorfx2zj0AUGmvjLtG7WqwCZHeGSAWDWxzdKR+zt
wmmd2C5TzZjF3uJi6HBI5FRISdoorZwa7RTlXR7tzqqqTfSb5kWy4w4a2jCQjlCc
tm7r3xRhTYf8IKJ4sLjxASqJTmLSOIQeARYkqljJoldafKTeEzHlNbgVfiLK/CZQ
p6SAGdBp2rDjV+24hFi/F09EQCS9u34hAbKMuGSUgcLhgvxXXpnb+lG5jqHnnET1
+UFxh1PpJpwuoaJuYrxKCGy0+DXRXpM7Mt3fkfYXm9j+6HIAyl4qOQa3Udyp+IXv
6vALxjF0pLlLhIicn08uLdI97HjtbP+0UmrkmG1BATh+n+47ZcBOD6Hf9hPfja5Z
nATY3fpuShwBH4kLBqEfq+qbYGQGcpk2S830vC3BAtcI0diMBV+gWzMy9saqhUH+
Gl4avNKV0eHNZvxAG3d4Fn3K2DgcfVugLqmhNfNkRsBTYPF4o8BUjmazhZDKxDD0
arhJx0Hj7SKfe8N56d/lZvQdADgJ/4NEAtKr8TIueUiHt7AhKf32Tcy4YmrYl8/b
gLiDQhQEyeqkcNkhTLMkC1maSprsrwg/x1R9m3ZvuteXnLzys1izwrep+4XtHd0X
Dg8OdO+/IuB77RmlFY0OkqcsQ7YMZmcgS8LkLsCxBvRBP/WQnfNZYg3/uBFX9XrT
EX74TfU0x7IPkldkG3E31VczIzqFKuk8bF+B49M4xBK+yJ0lDoQ9PM4upL+jz8Tz
UPd/yySzkPBYmoYdnWkS/RbxghSCc2nUnFTV2NpcPtpXu2vn9zC0n3stEney1f2q
MDwoj/rEvL4+sKIr0wZFVbz6iQ5I0Qgv/4Ynm6nxYS9PJzVX+l5LHq5IgxPcD3UM
luXynvpcHPUH0BO44iBaqJFz7tHi745ML/xi5jOMgzHKz6+dcWy5wtB9AXFtCNJj
tNUSfAYZeL3CcY+WwoFScZcw33VkQ6yhZyYSEaFJEe7IKEuVZnt/QZFLorhfncsf
d68wtf7oQnP+WmcQd2XxbLAnGWgZi5tTQoVHKQaxSzLbq0XkwDOjmpPOfpJObXBg
AujB7IY7a+241qX3whQVlME1yRmcgX2L247Tgo5fXyeyUsRzdwS1Q+c/CXi+7ocF
eJsqhjuhNPYZuHZ3bnFLKuXYLIceD/Ucekv/y22LK3wu2w7nDU6vijDurTtGrLDZ
YjZfbDAX0voQ4H2UMobyWgdN0eZhsjBwb2Ly5oSrCWNKB7wOYxlepAYHNhQyMFIp
OxfHw5mw+H2tbHKUK+WpAhkl41P7+JRZbdf0HLyDE1Mj8b97cCwkHKSsf8sMPOnS
4dOuhSmHC/Wi4yRYg9Ggf6PEP15tL4kUSF0hsHz+MFyeS7HWPPNYtgIyX4mByWEr
U21yZxJy1UesWBc6sFNh5hhqz4g1rZaq/1MLZcPCT0zUBZRhdvSdPreHYFIiGO6i
NKzyWRoMns5mK2M0ov4oKEYxXk2duFnw+i/mehlCNNcO/CatVke3Y0dFk+DgBrse
OdL9X6EXYMPBrKrTiTyh1lqZuJdkJO4NvLwl3v7ceq4NTR7upwSv1GAUkYzuX0pf
LUGinC01I3Yj6lr8eGHaLjsqNl398ANj685B08tpMJND+XdEmiedqC7U7gtetUoa
5ctUC3RKCKSfWBEL07BTTsyERTfNFyDfOCA/k6LKZtJ6fJT4MZ1Q6vAbT3MhYKor
vF52BfzycoN/iwkgtd1+CYKx2jOWJtkjltwakoZatw+iyPUcE9EDkxW7i35ehLae
lHT7+w2I8UAbAtubxTupMn/CrLCy584A4Heo8N73wqS3YQJKQgWumeUaHdKgfk1S
9+cCTBJt815Ao+R7JiGy17CdgiAhtasjFTHZyMxR3BuVBl4d3FsYOG8jLY0zwXJI
5Ga2NcRpQ6jxOw2uvykWEn6rpeWMZN5HfSRd3NF+//G/rV0zIBMYCqqfjYzdgwMn
I8SstTFxN+EjGkinrDOTgTTEh3B3224GXqX2LVhakK2NcEdUo6M0GkIc8cPAmhvI
0KNqEwOyukpwe44eqw0CyL7Wi4lECw7vXmmISCS+fUKJ2eeFrOqXRn+lHeLESccR
10p7Dr4wUmHN80HWpn1vfewqXnzoR+fiY4Mu5rYyZc7GOlWDhCFLD6Xl4lR2iZYi
27FmA3xH3D4zxeevOb7patZQQMX6sSFb0e4FPrx1W0/bzZUxisZf/KFyYgswhRIs
QZSmciQD3RBv8+/+NUbisd4w4pDWS7GY/4cmox3i8W6LjsZkGUMFDD8b2D9E+bd2
oTyBgTOHnlDtY7AJbiSTYcdzW7A7/cwASrgzWh4E2PY8CvmJJJ4eBhsK9VjuPJb/
IFzm11lFT9A+R7PxKIyk/DmoaeD69Cur01gv4nq4IyBm7t4mJCQ6GKPaP/8TxozW
lQ1bYSNzvEIy0cIhhGL5Yk41vog5b1AjpfSIxBX4XOfw/w7GaeY8wiRetm38iNmf
0RtxIuUy5wEOCUgI4sEUQmYixU2kWS9ZRDCRXEDU/nyUDLCvq485/aFvZ936Mr4u
c/cR1YwIo8v8hjs5NGPr7gEfL0qRTcHlHTdTEk0eCordL7WDnipnvmiU2dN+sSoR
u6q0VqWxQSygNP5iAlxwuzjqxDYWQQbVyTs7rCKRD0aE7zw99JYAAu5wYCmKw7+k
UEbvWXjKJYrzL8EnDDhQTTHHJvgsJbczedm/MQRgAQFW4QJSbleIgauyUdh5t5lo
UznafNrxehIIdbJL7BsIbl39t2jqytoZGXvXc+DYrxhwwFq/kSj/lnLa9fGigGF1
kDVUlk+R8Mq8yjd2LPwleD0x2DUIr1hecEt4EEqVBhwWGJcYHnkUgh6mhW1fqSXY
pMbf/S6RQgSaq4ZC9T5GkgrRWmbS67cRNGA6A9aG++4JnA0gJOlRczX4rBk0VsGu
/+k2ieMf/p9JpMp/cI19Tg0gpq+5p9Kh5FbVrXzONS7bas4m+F4xUxbsUrHKJHHE
dCHTxXxvaQo54wjJT89dHScvggd1uFQ+YbUDsinISmtdYAsmNJB0QPkGzd2mxJAJ
fAJcpV8SPkXR2I2Q55GlHD0IuQ4vvf4lYNDSoS6JZYomFCsvwCP1pMDLl60iLYvv
1j+hvciJUd4ZxiXib3OKnACxIx7QU6FD+mj9YKdVr+4F2HULEKas7v/dEUdUKvIJ
kYZfDhE6smM5Ss9N6SohUB/MEqG84RqFzjG8Npe5S55ZzluH1ni0PARQniG4XMa7
CNtt2L21WVRFKL2yYG+WRoejPTBQIL9sgnxI17f4qDcvxo4TG9u/ZheCARVlqPQc
liECp2R8vlhg2tMNLOJM4M8ZHhUlO993Gxk4QnvJPj2n+2JP0gFwcEh8AoyJpCwe
A4GWzMqz9mSLzpMv6F5ScSwHZN/uzrR8Zi07P407T8DDXn4spoX980LOAlyJhrnk
L3J0Hbj7BX2bJl6hSAXIDXuSnEUuRG+/M2UfzSuICfRdU0u/eRLwT7Cj1ISAEFo8
Z1G4Z2fkTAIgHY0GvhtZGw7P9yG7WZoOeHUdz2X/H+MmoRJOEUxbFhBURVm+do2P
PZQPZ2zLtRc01ZhcV2kZY8LIwgusq1G2MiKCY+CqGddspp3bu7wogML4LZmiFu/0
trOEPEbMWyBK+WCG/HDIP5Lqyk1rMOCH78q1RcqUxZEFlEVvUiVGQE30NYl+h29K
MbFpPjmiYWSMu/uBznD5+WxGD9jN99onAQuzlHwN3i+cvU9x54fUqGt1SgpaJwWB
Ee39sO74S5iU3FHqLP9tUzAz2gxwev0Q2NYZpyeLuH5CquIRx06cYbIJ7eeIffTv
BSk5WXf0SEhc58ZO2d/crBoUWnG8m57eiczm2JxPv+YKXHArDOacOo16b7/CpYSO
0wDGR9rvS+dkckpgmn5xXYJEX3tjNxenLBxdU9/Kdcn3R66raCbSOG9DEFGBNRi7
EZZsl8WMtYNlRuFKTXPjeuip2ZoAyghi9UwYooInwI0ZS5QNJXn1v5eFR3t9m3WN
wMyqIVwUR4kTLrtyVUmj+WTYkJoa1BSfVNNzha3DKbwW1TDXX+uXSZo4fjLXXMHo
9/AIQGqBv8SRTcoXfxyYv+J1n1bftcZPXR1ZLf733dcgIN/tlxr0VJ4W1iHO8paN
H3yMtBVdB/jyYvyKLZiIV1H60Ags5derCtytcDTiXVrxCBLGu8jPbPhAd3Pz+o16
exy+V/g65u4cg5yWd3vYEOfVZdo3170QJWYf2tVsoLwVamJXXOR1+a+R1ZVpcYif
Qde5MFfodEYBF2hfpp/zfJQJLfsLDTZ/rSkOO4LfYBa3iq9jdX2ZpBC38xb71kTA
pRntxhNibsL3gXp/fpt5AJ5AMeX+1q0vSby6A6Xl6yEZUHL/Hqi9JdVeQVnhcRE6
XboJ+UcA1fRZmF79xozIlCwkzYmebv3rXfea09ACqLbr7p3MzlUIKkCerYD9qPwY
7FYGcI3mH6fMYXEJJu22EEM5OglbOIn4bEZPIzyTuxSHewp3agfAtdeoZLmMXeTN
SGA2hy7LeGyJlHjorxZPnAdqpnIgBI0orlB4cXL4tDHOkn2AcaaFR0S0rb938HHQ
ruG+Z2a2MkFUkx7hgJI61b3Mn7BrHLECI2KmPPFuDrKB+ulSda62s1ilzdP2itqu
4nkzPGGinfh+sn+93JF6RmIXH9c3PjADxwUPh3ggFvv3ZqSb1ZndzPXUhHtSkLmx
V6zB9eEwYwWcsmfDoWZX6zttGyEC8aO6EC8wkDUG+RZ6m5/gJEF6l9+ZGTjUglsO
ot3bVBmTzKNAUrQXnLZzjjHUOa7efYUih44Wfur9o6uJ9r9UnZj9c70vDc5OtWwk
KQudG7giOBviPX3z7W5LiFpU+xbm9GDM5KWUt37w7MG0D5yWo78R5/HSQtYRrIOh
9rBlWf7dH78VJMAKd4VP/uw9pTqwO1L9OTSku0igMyLQn7SWN5h73jjcIkjzswFQ
hnZZU487+EzagNPexIlCaTOwMiwgQKlaaY3VKMatGyV7mAByIKliifIlmwcRyEr9
AaeEY5xo8fXt6cG8rVVD7PYyZO0mXaXne1RqZvzhsaTU9Subcxdb6HcOggFeuMqB
WriFH23ThyBRzHB0NuhxkIssqCRKE8GQOLn1XUamd7z0OeZYrKsPfmxLFKbwB+oP
YlSPetPl2hvQ1JD5tSWny8NI5Oh+Y0k48WnIvo/tF2sTTCLVkWLlTrhip2SGUbv3
DeR0eOAWhZxVXHFDbq9tx5j117jwEST8HW2uGi/U2kzNgDG9gk4qdTaBmHauMBoG
GsVJdL/BXduFUJ3jABdIRqCaK0XdLSR+wUJgTLggPlJ6YakjZJ37rHjoYFO+HQoo
IdV5/u6CKEpYwPIIYx7Ll4JASGUAypv+xj2uUl4eH5XvVk+hIygxGaPcHngHUQo1
1sjLqaT4ED2yZSl5BTDUxeZCXRuzlxszagrVhR0hHEG8RN8U0d98SlBkub4/a6iI
QrDYPsDpVknt1AVZCWYahTDjTXNVRMu1U67sycUx91A/ALkpqqHkSFAoy2oXTTqa
nRn/nSIvm4b6i3p5aQRaWpvBwfguDB2tATrQ1AERkf163MLQpvyyyCSVLooHEk9B
Tdev1YXez37AIqILNgSZyY5VBXBSWhPrCdF27NITxMtezNhVjk6HDaGerYNb3IsI
lJ2/HDdT6l+xV+WukfndEM8PvP2o6My+TsxJDbPzFsVqj/X1cfn+xfno8ngMEcLl
0h1FzNREPshx/Y38su5pd6sVl5p60u2i7v0KuszdXxgN/1BM/XTFs5lO60H88T+m
YwRmwRJctMwWKQJ3UyZiprnxg1PTqGSKaHRxnLaINOm7k/tYRVm6WK3nI6SToOua
1aYEJAB7ujan6wG0R98Ss7ms9IgqesPf6JWRV9WIELzBNwuT2a3WkjVDwb5PmxLw
IH1ebqquBSyBJua0rCzu/w1+uQXB6c884T9qDpWJzYp+WdvBIrSbDGJi8Pxi7wsD
XFiYis3Pmg9atZph9friNBfkiLp9hjmQowPsHUXh5ytapdVdtEqNitkbil/RKxop
NvKueypq6ULvhuPFXUJxRXKHDPV3l9W4CQci4eZuuGpzViobTRotZBr2IWMk+ufK
lfpyONq0OlEz0Y/cvSupTcZCQUMut1YSIhdAV8vGApkiY0n/tmDwNmfbJPmJNV4k
ufzfSTYDuO98vecxp2ak13roo8JPE/Zr3fUQgvpbKCmaw+cn6YXpSOMmixGLalR4
yX8qY4Fo+PY5kJHf1Y/DGrWT0S75gdIdUVsrTiPMaA9B5V6WYMG+/Z0svhRaBvQR
28uYou8gMUyKLJgGsPYOYL1KrWyC6eLTFpfVo9T+zx50w7yen2SA/0jyDeSF+t7i
QKWW2nSUj4YIKEZ2mietnEsDxpTJ3dLGhT2gl63jOLAg6ILyc5C5k/wr67fFOg5O
dUG3wCoSgucNCXO91uCMMd4Lum09zNInTCv2+mh8hXzRHlLtAAEL2qIOGrI/w3ye
kaSqMdK7gtSk+FzVzZubjmJAOgzkQLPnPWM/+sOkIjsd7DJRZq24XmKqD9lcX+in
4M4Agggf6EXC0PIvPwuepVWUKAt0P8t+l4iiPxqHHBUnC7CS4+lBenvKCjWHRzLn
RogxUDRp2QuAVLupNlTPSBXo3+GZ4FWackvXBT110bxiF+skRyNsAJV9DAKeFga8
e6+ogjAXrvd/m5xrUUYZkdO4VGE5wIEWrDuenh3CXWFDf0YwNGniJX1SPD3QdzbQ
aCamCX0brkuvli/JoTNpMS4mCn0ey6G5RZ4PGKDj3aG/r5nyH9rHnwdwlRrtDvXx
vJ39t10FP/Xt1zScJ1yHlo39cxKfV6o9gm8unenzzPvr4OJr0gTzJpR7evoqAvLW
z/BLTBiKrjQF2uMa1CF9g2lAFlyTeP+hoQgclXvJNZl5igXskNR+zPiR3klwqw+Y
A/8ir0fnzNTVwu9c30X2so+a28CIJtz1Wo1VUoysZZHat8Rbj7AqKbXELqvLQxBA
tmC3YhclgjTr+WicU43nnjJHAwjB3odjgozDoVwzX8wh1J96dgiKOgTr4vNqZ6V/
eSiKwEUn6xiaF8Cuc3/I+HKdfXxps8y1Uwviln6mSzdBKi0LT18u5Ul7Q83LSN3c
axfYswpSxNOpvle9ZOk+SmdjzGCyav0ZAc36bJF3LhOIn+do4rIM8O5O7PXcbKLE
g360FJc/TRv13u6drk3w2qI4Y6I6Ls2u1n8JFokJyzKoECiUMkaR+SGYyxKM0sn0
puybpiw/83Zynn0IVuOU84d3hc5QEXbs8f1XvzWTQWouhZ+faz2kqKOcecMlIk2e
PYe4UKQ84II/H5NEyMn9HIs6H8gvgDr0eM/CSYAgBL9WudgAHk+Jdwcx6JaHrdat
Nm7gCfgB6BdXzYpu+39IIgVMyjjzMudtdnyi6yOKFHK4V+8RZ895kiwCQQiKcc68
XemUb5R/kM+KobYdOIrX5WC3PftvStiW4VV99iEFt1Cgj2IfC5wAJUjfIZ5Y/lGQ
lGNOuspKbjE17hmpfo7KcuQLtAqlOexx69lMEOxkpijzkk0xwc4XHzkDQdo3sVe8
GNCftkuXsuMdw/NFk5dCdlI/gC9rKxEbkeDQ5j9bmwBQVYdJrNZUTXKh3a0/ezJv
alnBGA+57Vc3kSOy0dTfQm0X7DH3eqpowp07iw1BjbhOvneSwb6qnPNQR/9p4mKp
LuMNQzH4bZ8cDf+s7J5xQYY6I60cXa6Fu1IEQCeMXdOsRVjleoUVYBha3EIO1GQy
w8h6wsV/l6119SjY6m9dZD9F53aK76hqriaPpgRRL44/MG5VjucXaNAd7e5ufYBF
yyFPG98mqgiLJQzD47B6VnLqbglnGsmZG33edxqe3UN2uWTcM1cuD4n84LRfvYdJ
K1Dut72UryVl0fQcxRWFUB/78qxjmzDgAdtYdVdcfZtM+t50NzlXtDCzmD5tK+hd
QaGpcwb7Nn9QJpWI9yDBaMGdZLiYF4Vyk0FH0w8sH8C2kRs6dUDgwUwHO0aPdhH1
A9k5VbdXUUI6JOiz0zFN4RYiXBzxhCoJbVjHmyn39yqLmTnltDpkzlsUBCqGrCpn
uKUja+XhRza8pfaUiWVtcdeII1JrQm1aUxrPza7/PihjT9XqT6L3mkOsoCtxDHUa
9Lmrpr6hO8pU9CFQfimzJGfUbH3k2gzM16PRyP+vBs0lEPo7cXG76qWTruI3iVyS
DodXE+j9OAd5L8lnFZQ9puvw+2ZrWMnIoYykBuz+RXSSIQ9QAVvJ76WgzkdIej5G
MlirG5JtSj1SQT+gBaQwVr5OInLMjo32L4EJ8LZpWvfZbALEm9Y1CFyQ1VeK84zK
dOvEIdm15XvmiQnQjAWF/T3Ksk3vI3cQ2HcKgEu4IIqzHtV84mN2gTlzqiuP9OBt
sfXuHAKROaMWrK0IG3BRdNYW/ch2j6Q+/mQmgLh+fRx9vi3of0aLlyFaMhjyzMps
1T5oYtL19Cj3REnAjhdMXo3uyV8Ec55uv60BlbM3rvCbPLxAKKl5m+4ErGyFDweA
4wU+77ATm9u0ZvrlN1MpLeKVfYG/d0xiUmUMkL5v72npwb+h7LjGSj6Jha0q3NSO
yttI8Xz/G9myv+zJzECHtgwX9wcXRvFpAh1UcM+CNDqlPrdmiER6FkD+v4/JJQ2c
n5j5zxvf+oRGCPj/BhTY926SrUGJIXtopR7f/Wadm5NHJZQxe+IbkZfW+PMRk3nq
4nLL2uju9I0SnwC575g2aCxXCJstmMCxrk9KO1bHFcPPz+cmMOUX0MLuH2+zcd0t
9C/J4OoZwZe5KMuSswNmAhXQOUHJMIBfHzG7pJE9RDYemjL0+G592Pqb0yw3UaSq
Y5/CGpMghDAStqDuXfJ+4n5VcZSQ9XtwWTWePSybF616pP74WZ2RU0ntqIM3PQ6A
h96eWR6iTVEyxl4jBUlsHXuDp3sUZ3m6Yw6efHuVSm2uaBMZXYUWHPSo3qd6/aDi
DjZvemk3nMCa3u48npnbPViutPDzmUtPdaVu+OhPzZQOkiJnK+c7olp68PIN43b7
dyXYFmcQt/Vfk6iseNm1lcCkGpW22242o0b0tvhtHQ6KILINamGbsry6xYh989qN
8uEj2+q9X91C2YNhBTbrj/IhMXIibi8Zi9P/Ikip0mpYT3Ift3C/Qg1C4b5SXG/Q
QZCgqidazuCNbOzcBu2RW80xq+zFG7Y9nndMxP7sI08KkzUmzxumr0rF2+oy249z
shEazLnZOVFgYPTy12qEYruTeC45AKXO/nVJqhS/jB65TYVeej8NJ79wOMh9a2ip
vYmyjewZ7LV4e3Y6p8HIwugWgo2rIXManFtBMkOkFsJZcqMC+eXb6zzX0iv8/wsd
HnNB1gIJvcbjT+bMHO5ceRS/UhgfwSWBiHU5uqsQdQZ/kTrPFvLcmbMjJROS0YoN
EmBsrRmQ2jJGSyelgGz8h6ZKkEn83voZHrv9FGPJmMP7pCvYWt5CE1QCkcLnX4Ek
s5f2CE0kH2/XrFVE1biQf8DRLeJ5f2E2GymLLB7+/60CnVoaJDtmIQYqY6b0vMII
CNYRuasY0/J0GTjRR8kAUzmjS6kUdGIrWH51ApKFXy3yMZEWbfwqK2r6aOIdIvVW
tvG8JlFW7bO2fI6BFq0/sE+JOUeL43K1ssySuGcBWBtgm5ELlOFs14jM3tqsaik8
sD616DNN7ne92KI1f2EC3U1EfNhgE0oHj4o/IJP3wjjj3ffe1IHnLa1fhnYfMW5b
eLVjERBQWyIJNin/z3GBvqH4bvTggYYSyXHq6Iozg/zHYwg29kExUG+CTGYC97nK
TwinKIa2Qi9qPopvn8ITw2sQ3IpEkx4P9ck/NmvYR4xsktEv5U/9/7/sxYXujbh5
dkFDvbJr1dyF1O0Y59uhXjhfAEBZyTvQ2azodwTbir87hmbipgjsXUwWFcQmwM81
zPuXfgpnTGzapMXbPea7GFADCl8/g8w0rehWMxeZdEGp37xXppuepKBmCsJ0wmv1
VoKe5nsie+APdws2fc21n2/cfL9o4EbO4hQ9sGtGrxkNPrabAMY1ywJlndtOD5rM
93c5pijdjpaaG1uhG5VC2dYQSQGDz5xeXjanbkjCbdqTjCOWY9VQ27kZXt/DH0iB
UJv5OK9Fg5HcO+hz/lsVb2sVu4qFgRZmN6gv6F9GllcZ2BfbO9cvZo987Hm3yaf3
G9qYZsJDfoXUo3kCRdLNDUg2gVrUSAMb9il3y8EqfMjwQVpEsl7F5l0YsyqVsgTA
ZK8zyHckBMNHWvwV3dcQAL4Q8lS8wHNp8/H2PuHtLiVPN50AeE8+oPqcdoJ0gK4p
q3zZTXQgf929a4/D5JaYzbOeZG9R+HwrZtw+b0td82oQE349ROK52+OwqKRcMxnb
Lk7FU5laiu4i6ELjMtZxZAQx0vXkOeOpGB0LKFEGIavZleizKgFPqy7jbfbpyCYB
gRUzmYavmrJ1eJJwrFnCkR8zcTUhxgtYX2kB5AkFQ6KuAcc78ZvGzsVBe2btPOgb
4DMmkj310k9OauhN/KiGUOgR3fq69xcDieQGVTC9/mmq4A7l6r+RM8AXUauhnnwO
4sI+itcw5rsIZFPECDxzJ+PAoeW+R2TZgNmKuGnRQMJiBNeW3lSteMpQ2vPcJcjT
SkMRoWxh78S9CZexRd+SuGSGBwyU4IOy9My3HKzBqzE3UWDAI/OSDMNwnhCjcNgM
J9BcbXf8wsr5Fq5g4y9JvGU0YPsuYYrH2XofgEW6eaP9pbuw6fsbvrnSK/fNUEj+
w3sr1vu4+0Df7t72Unh3Kk9ajrH1X/B7GCfz1jxA11zUzeUOI0ubVHu/9mvAqRW9
7xq+bIUgr44MqbRVlG4UEGzoRC6hDSnNN76NASkKBW76NJyWLfhmdJ/YbPfSUR/P
OYCHIkPBu/8jQk3Q0nSvKr4e4rNlKj2OUC8DsJNMyy3AH6Zq9mXaQLmcuQGStIbV
GIh0pv9po94BzdEx4sUqT6uOkKQVAkmvlUoWQOIg7KuKT/iLVL4Irj41JwsUF3w7
15Bp+/vIqdxNq/nKR7dq/EZYjAyoCDX3SZrxL0KGOEA4IZkcVTl4xUfwDcTFxvwn
HblLeprMpSMgHQhv+HllkxoUzJnrvlv7XfmLLhiu5EhEr0EQn1ozrWYrfs19lGNv
RpHcMkmfMR74T8Vi+kgyOW1E6A/AH+ml3xSPz4LZorrKfGlT255w3uLJwbZzFbbZ
B472zxsG4+HzXe2eKxwzo9LtvqqxlUGYtWYMHUOqbZM4KfhxLmRQKBrHEDRJl9u+
fnyhESVyyfUUmVLxWafVU0bZHr6kqjVDPBSZzmZHnon/Bu++JSnMAmxv4t4PS91Z
QDoZ2aHPWoVAqxk2iCUHt/bRCKTuv9vB4SL92ckOjcXnrXTDtgs/LmVQr3AEB2yg
BgyuFcO+ltUfGfafAXGXYrG5nutNmQZ/rU3vvBzZ/6tIJux3pf1WLe6T2kwyw15A
xZbT9ty8TKqGMPPE+faRNxG6XXDgkLbyDmK14FDLo+bAVecpKUdLkNAPdmpI0mWb
h6Ypmaf3IZ84xx1MYY5t6DiTs7Hwnj0AqM2ez03j/T6uug4yy/PsibWRL4xZ9faQ
84iaOeUUe+2hhaEKApNIpJEQgyzHWQQLHcWD8m7+qxyHDUzK6fiDHUJlobcMDvjh
cwpiYwfnRYYgpRcfO7bkIJLeTFXRFM1WePrv91K4/MuyDADaKBxlxXtg1rOIpj9o
/DE1pYELnAgLRISAY9wovY06nughZ7qAZVIWiqXSizNDCu5Trid/bkvRkZl9vGxS
+9WYWOnK5rA4hLAe/WRZON40u2RuX5dqAPsa/AR/2WzRwVJcqQT/zcKS5pdwhcmP
OKtNn5QgHu07al5dk2FE+AJ3j/N7eeFhbn1iGb0PmbRnQs4F0QKF9lUh3BW6FjDC
/Z1etSuD1SxkOHeLhi1VjP1uSGfw2oMXcn6oVNm1Y4p8IbPRsJ/eqY9FQq3ZojIo
FaBwpLBki8olpDEZ6v/K2J1NtlKMog5+XxPJBwNlycDoqYPy5Nkc6UJiVZJB0SZV
52q9B10h40D+U3q+CORCpBgRMYdqCgFx0TboFy+KsmfBNSvgqyieQzKoEhm5L9bH
hMtLj6pOo6J9UZroIJwuz8haX3uH5cML1Jr1QHm+sYc4JCGvruz1yIPr/114R+xj
DO1c+OA9VgD/9ZQ28ARYMcyGd53NGoO6fGFo2OVzloQDv3o7Ux250OlM6GfL7Vyi
cWJhorbe2eisc7qxSLUdTcjPXNA7AY3pDhuTxFpzmws4S+rZ2mTtR+tXz9JevEQR
a7xfRFQ6Ckk8pS/F4fQZ7ehM0iRfXysetDBf9vbj7vwV+YdSdRqzII/SjU4yrnSq
dcwfkesoR1zlXeTlfq+KDRYrBW120cvLQBjg/lhV+eIUVfpGhUbtfWo2Oo+7v6ZW
aSkYuP/2hBpBXNAXzOyBO46wsMkEyqfTRpGTdwwE7TWsJ2d/7fzjKJ6KKs3hHDbl
EAAHzn5Sj5kQHP2hlf3CXD2Cfd+sLfq/KSHaNwC/p/uRJOAVrTD0W9wmxkSEfHxO
vwjqoguaA7BJ8BqA5GGKraguFiQeQgsWKQWXJLuoAMGEnUVcF1B/iQM6iol4cyTU
OGROoAS0y4/w4MBVY67I850OlIQDGKVIgOAtpSR2gutREE3vWug1ER2ccFpkYTYL
diS4ei2RTau/qvF4TNYvrE/kLUpkPH4p0OUZV3ggyNG0mfRL4w/kOqdA6+dmtUws
Pf5Lq1F9bcllRRFD5qL7UerGDO+/cjPLLl773rA74YMbZ74gujvkeiMliJ1zVr/E
bOg5Duxzc7yt9UYTYTYDY8cFl/4ShnyMwsYAFQwpimZS1BQW0saNa6MVTYLvJaxl
vq+HADmXGDAspaIGvuTVDif92pcecA5F0kIQ+gMVr4kMlsm3O95dib0uxYUVXJT5
d2Pmuk5Tnsc/4q/NYkrj6WBdhzHHeyktT+ohlFsvpW6IYDCBtuSG+F8tDVL/R1K6
fm4QXVU2KYNkNkxkQflY2ExZifDvl/7EwG6hMfepP6S+0pg+xlO7XPjB29nksEIh
I6hLMLhUGf6s2u/T28TMRqukhRVCT7rkkRHERmtBkFC6S13ijbOD2vEoe1Fe0XxT
FhHaVc1Ih5Na6gi9rMtGoGP6wkFR9nX3UHotBBLAnStY8r32Zj+T4JGB6A3+NKPR
dAyvYl6LUcS+PqabaHskqeSsbakTEI/mqto9Ia0xZLOgJhBETgyR8euEWwpyRr7R
9LHs7ILWINUyw3Sy5ZUqFALXR0gtO/Wv5kts97QXeaFdKn4A1Ait1EkRsxmGmQEy
vuyi3AnGj3xKXdIixI42U5dBLB+sPfYIUTuk7MipzPIHB0gWUDmdHxahQMNTR4Qo
vHjemoUkR+TIxfTtZa5sUWrDJjkKCf3nzGuVepBd3BwXiqL3I6aAx3jJE0KoHjVl
gdTqOZB1rgwAA4UvuPt2FA95hoWLwB9ppH6zg1/diwwUJ9CXWckHz7OMdw+Kq0OB
oKv1JLE1hV6QxKgJvDIe7s5VCbZSttxyZXCzCazS1cI2t4cpvzC48UNa8clQqrNC
N8AKFXy0sRAAE0Q+vn1QD8ZMgLYuEP9iE7s6c+uEhvDDf93zDztt6MlyTJOfBdBN
scwLOREDN584WUD2QGkNd9XeqHvbw1UtS49NZpspUE0GCLETnHeg6QpCZSvhnTZj
c/if6JtLnXJyNSkv21Zoia3TABJxJ8ivCLK2hQi5klguqKEl0iElOphlkMXaCvLL
pHhHa+VqlTB0N/lbIlArZYyuS7z0dQSi7dqjocOOw287qPvOSx3s+vhYtCmMP2KC
zeZsseJ0XAbN0lf8uQmopHXFPnbtom2+SgEkzP/w14z8W8o1nquf6MhtDKcDFqLm
0onuKp4VMS/TWpClF/MIswgMW29d80Px7GK/WT/MB6ciuDMqMcbHROQWKa6PUH1p
xbKnKp+gzvoq2z+Wpq/qrGVRavut809Hn8oC196rJ9Q5u1SmKLvKRGO/GppdXasr
MS/JoJghl16xC3jsyl093mnnji2vfC62cdv49LE+wiQjgSc2DhNw6LbTCaivTkFR
QMOCAo29QQcCE2gvD8xJSarovoBEp218sYHbDyge70g6gjRAZLdU5zUWAmCNIyrl
E67GWkezzCjBc8JMVsgnS1AZl4rREi57OcvJaN707VYR8bwMw01k+KDFjrxlSQwU
lDuLMIVSrk1UseaJ/+0iYfCUmFqKr0z7UFzQGIM66qDDp1obkUaHroTp87NsgpM+
0es1ulr/Y2VoAld6h/7uuWAQ1A3r3bKS2OLhxvA7S7UxABTHRjSSNS6BTnuuSsjQ
KQgou8P2Ap/fm8k89m8wBF7jzpq7TNPxwyuf9l4uU+paf6TnXwjf8Z+UYjxWAyJe
DYyiomWMxyUh0X6ozsEVSV2sZyZlEBn29/3/tSRhzB/72E2NTe98T1yJsyQI23bc
i7/m+WumJtLRYO2dxoU2sPMd8SnV5oQ6bgoevfBF/C7BCp7G/ys7r3wCwhPF+iPu
pX/fdwpz06YKJyCOb9X6kaqsqA676V+EO3mZMMfY0LclgwwpZf7vhDXXg2k0IOQA
B2gjZ9QDm9EvPKMkCtv70lrXT23P4Tq6ewWtdZD/azqorbjT/CmjQ3u3chrpiyky
gNsdWJfQYfjW8W6N/OSjX+88mbfeWqbiFuiUcMT0sJoD3wlIfi6IuKZWmtniNCvg
8/kPbvWA7oANJGk71NSix6YfLr8rHJY1x41Nu7dNY48e01AWloCbgkwpgK4WEX8J
gDCdIGNwp5xCncJRorNGUXFV7OyzAYVm7bt8Xz84mppM3Rv97MTxfrMM6+rmhA7l
NvjcAfNsUGbeJW8m4269tvdiQSyO3zgLBTuowAelLKREA1Tqr4PMpskjb9Nix2hH
nKFPTdWdNWQpGI+pISvtBvKPLvgYlWNcRRA8uTluw0E0BFzRZynZLej9fSjiTQ2Z
hcpkrHMDhY7u7gm1/6xMYSEr4XVIdmiw8EnWjS8SBSuD5p8qWEcP4DGIW6tX73Bo
PNDwxqzjlRYY+uGnuYPqzkfiOT+kxMts8TLwfxC9Y8OKYuy1iv4OMEqqUVgA961Z
BXas7hwN425ehtGzkzFhmb7wTbTXS5TjmyR2l4TMIZw8AcT66vwc0ZES0jHRLlpt
sByYVmUtB6TZJDoavdS+LYbOAnS6Z8J/9DR22QOeMlx2C1jOWL1CgIQYCZbXcFeq
B1GdttaiaWrXiUEAD8cm1aWVHxhuzgjJg017kCTUFOCycemjeSOLPvm2FfR9BPtI
eGI12RqVNItexXX2CV/8FQ7PSOJikLrkb4Bbc2JE7sGAUa8H7Mt/7FLLrKNMCmXl
nID0lbu7KU3kYlekkgI86fWiq6W4/UtuOYVB8w5Y2DfvlhW9Cy+FEjLjW14BtyzE
qW+0NmizndfyQBXOzEdvT+CdhmJ/4M5w0PkMdnf7Ude/NVcbY0UGqJkKekuNypRG
O8hcTNTOjcrTH1NgjYvd4bzO6pypXi05xVX4vJWvU9IQ40vvmQ3RUSw68ThxQL0n
U0cwi7T/hf0UeJ9NV+l0iBXgq201YfL6uaXbRMGz7x7W2O2hIJl8onQCr/WjKJS6
r5lOmAzOj8sjpHV1LqgS6xK77shpSrHDz65KCKjkx1YQLOPwMf0wC2YaO6tAld3q
OLHnahNQtRk4wxmy4glysLQmpImfWouU5L03B5FWCGgXzP+0izWl6w2qosHf4j4z
2QaydqQVMOxAjiQMgPiWKkdXu7OEEp1yc3znXnyd+62Wwl4FBXkN/jTe3jAcYnRH
oHKcPingTZHpvUkRsVR6KQPOth8kBlFFRISxsh/4xxRLgy5Gyrj1AnnYPWautPUi
nkAL8u3YLmXumT+sb6nL+DvQS9eoEdcnWdo2iVfAzwy5dghrQz0JXCYyWzRV72Oz
hMkSgBfSxl3PQSq+riN39saKhyGBXvuPJUZQ7H6tzQhsmRr8Op0rs2tjGuF6y8U0
+qXxDbHsjXwEr1usLbCZmVINK6xH8jGJ6qQiLh8LLkixvZ/2eEW9BulYpuBJqi38
poSBkblCRq++M4139giyxzLr4wltlOCh53wl9zEX1TI6RFoLfm40vPfLMFqJuyeF
/IFLOE+YhfBg/HZALyMoOY05pe/IR3avrEyYh9GX/RzSQLm06NzXDmVD5MAATkWC
T+ToIEzXqZQqaWmlmwCXAerT/ChkaGASCXiRn3S5LWqjIoGJXWSxwktWqAJLbQpj
3C8AbBds/zPv6WR6CGpeGWyNtO9Mieiptz8f8HUNF4utFKWNG+oWbJE9pihChaTT
J5j2VuJqF5lAWHtFjJeg0gtNvmFwy9191vzcoTYzRHq9vZjdpDr60mKjGGCnjqW7
xCoI4pabL8bZ+mz8LQUmfsCGZSzeXjfP+7ArCz3OA3HsyLHbKi+bFZEt2OEh/9Ci
v17dgXeH6nvjkq/u6JqPNUOQvZOIRMLXfO4FOPnQGU/7fdux9DU0YnEw/P5bB3d7
zsBNBG/jHq5vZQwOKo8vtqCp9NGApieuhcERc0vbQqvkBRe+bpAkDp/cCORO52fC
sKhqiekgMZnm7QcaWrqvysZpq/BDeR2mtoz1IzLWMNiAC0VklcbKYsEeKmI2RckT
qSjvdtLdZIqstdIYTREq0DejeXFpg6FZ0txlmcCbr0i9B83U8bplLcQHEcUn8kKY
MP1gDBcjxvxzlBqmBIJk8hDKY65QD32uTQFGFgI9TtYgx7jBs3FQ30UwT69ohr7c
hYUqf4GmLyiMOFxQ3TOEkv/GXvXm3pNudu8GSebZ/hTRo/Mx+55bWrimU8r9eHQ0
mcfjfN1LcEYoWGzFE4Px+CBRDN/+6CDNW2oEm37463afao86aBdhAk9gK6aIMvfN
v9qtT/ocGP249JgXrKFeHU+mWdqGhCFSlsaWw6olfOVmz5i33wGBL5TQ9kSAwSJ4
2wAmIMJe1uFAs0BRgK0uvY0/kEliGsk9XSt/74Etj6wekUI9BrGj9YdomMMDZFCh
vqBUhaCy1d0XpeyAfg6odAHMvsG1eIrePmOlEM8KFNV8EwsN/Dql6tnZOeyzc0IQ
QUgICQW0ihZsGtBJku4TuWGWvX0Vzus+smZKi3ZkhIbh9J88hE6TfpiswL6orcBN
Q0T2O8uP/61iZBRthBkQTETXlyMNqz/NPxXMaCm0gYq4oYvulk2LlVwFAUEjCcH7
cQ9skDndEQWM7L6Vw6VL507msgtWc9Td98/yX1Neotpzbq9YYqXG9sFdUVrNmEPD
OWBeyJqbRR79vvH6H5qgdZEMcUGEHIJF3dgw5qPDyxd9QsSqv+K2ZUHM+d/e1JyK
6sDOcXvM3uJBshLDIItULuVeaBcZvEC7Ya2nNpUU3z0FBY+meeHHmDA6vHjMEQrL
YOdI/kO7bqulyqx07bDuQXel9n7PGKNBh/NlknFCTZjJKbluDx3nhWSyhhOZ2w13
iFiAwZSQLBZ66bMlBw0wW+N9k1fqVOm3ObIYZ/NOB/WlRODGWeLoR1E+kqAeogOD
TRI9fZs9B+uRf8yRfSnUys5rxM5BC9QK8oyf4LUtlSzcOVCgrXKzD5p47wmziwG+
6N9naibIXK4gQnnxgLMPErQ2qHxigV1YUdWxOoTUC2UIdojBAL0P9Zed0g1iX9Bv
v7ojaL+92r0bWvLENIOYrhahqLPthJYhmF2X7d24uXEjm51aPhVw3tDo4mtYg7QP
24kTxOMeEwyL8eJXNJ7xgTf19F2wAaBE3ORwG5JpWcg9/7v6ijF9jDmTBMRkoA96
r2/wj3vy1QmrRpnnWVXqlntb2jBS0TOwjn1AxaHrbpjcT7E2JcyQjYEmynMAV8OG
oiGhZo2UM6L50cW8ghGfUT7HgRVU6xTWSrsUb+86qjBQILvq37g2TXnT9sRjaB7q
txUwo8RmF3he2T9vWMAThOQjVIWyNmvG/l21X5Cal7m5z9Ck5TWQjr5qypYGiE14
hhXg9Sr6Oqo3ja5IF3AjjGXvthB6f3cXCnw4SPXVqVYmcnfI9Tbss9WmV4DaDPQ7
Z3GLKqGMyJOp5QM1mJ//NGAGugP+jk1Xs9XoQV3/JbS1zsxD+6h18C4yGJ8tWBms
sG0uL0kS80Y9DJ2P0VKlrgSKdgKfvSM9yzKclY9pnhAsUp+PMIVmDYJRjdsIA+YJ
DaycQmTUM58W54VYOvphSYzfMVjeiP/BkJWmvU6FNuEdoztFc2CHcN4YVODgZcm1
oWQNooY8Gy81aaJuHAlGvaooBFmemG35kJTTBym/77tJgF2j0TLBqYPOKQrWnOd6
Dv0Q/4msIRIuLFJRKkEsfTtOZIo8SwuzOCoP2J6HfcXrLsLhe4PNP4DFmrXpsiGW
9D9bEjHm9jmO65Hw0Xg2qKDADd5f+lSSsl8/55EujvClLp9F4HOLFmVzONkrxEVU
Ac6L5MrJzk2re4PK4AnU8XgKEZWeBqzZcF6Sr/jBmgcm4fE07WNtINXFa34XBMZ5
rdQnWxCwsG2MLXqAh+z790YLLlgdXLyvCdcJzAKyTEbQsttYGz3KTXGBE/FC9mn5
/v29MCa6udPK1RJUT05q802q022azG+dvPgZuxs9DuNI8HFjVNnvuvjAos4uwH6/
Eckk6sNfPiOztr8+xe7j2dtA7A9wWS4KB5sY7KRmy98C2dNHsA/Gfw79Gryw1coi
vd5n0b9bVp8r3KT3bOMDSwDbxjQ2+Oo8uRAaPXSCAaY8/6yqy5TUe6Alw43Eyhkp
sdb7+80uX1LWdOUpRKT++7EFOKlbmOKVI+Y9gqYrCJBtWXEBZH2Dkbdcljh1+Tm+
+sSyN3MAx+V/JNh1bjXUEXiXYX6ptHtuAhuJiYWzMZAAIayAjtM913nLmobSnUqP
e62fWrmBhukf5R7+5K0z1jTT7qI5aVfluvoOpJSFbNB2+TH2yhNxs8IoKv3zVu8s
xBOPeHpLc8+VugBW9dv9/fAlkhQmqo44nZqnqtc59rvdt4SHqa6fpKV7Yd51q4hI
/MqFqBTUKLoSflDmPfFN3OBBvzPD/h27GwGQN7zE3Zhs3CDhypu+cakpmZvAXBQs
TrEEE+rh6YbfbcZl0wfcJXUWGxNTkb5XldjcAwlcy4QqA3+DnaUkM6y59+6sNEcA
GBVHVM0CxDBXdVqS3pjXXjJ03EAfFjP96b4uYKo2hSpzsTo7OHQt5JA/TjjaRXiJ
SmBjC5rW9NDupDsBMIVqc/hvrPu4cYJWvTbrgkRah/L1lsRNMfqO0ue5EnnHBwiw
CU8mjXQMk/1eoTZV1oFz/pwmIlDht63ss4aBZco4l5ypENaW5aAF7R+GRSzzURHx
p1ircvHArIM9lR3Kf/THLEA8eApEH11H9ZaaVuC32rYrBDyIIlB2T+BWMmCesAdl
YbL0VILrmJ7OXU0dhsqU4UT59urkBJiTRn/CK5nx4gyZCgpQkVyCpWy5m7cRQwHO
D9AKUjyUGnQEPPE7Lbrthy3t0GHlcqMCrQoKrGAeODA+lP6LwzBuBTJAOObja/kN
7nSQcz+IEF8GXfOhyUtnbFU+onrVt2mk1m3Y7G/sWDyc/rLymB4cNzjiAj3SLweW
Bvem7pu5cc4WHvKpuSQTD096VOhpWQdTVVI0r9BGCUobkJlNuXA+vVMUwGRHFlui
WgO7+GoOq6o17DLGngz+ScjSXg4esoJ1Rd5AXEuoxqdV7aDJPvCDqlcNpUiwL2AJ
7dODYX1ocCdDUgvAt2jEFFL7rkrx48w/D+mLADTYYX54GIz5W1wnyJHIt27WEUMI
6mnv0Ai7vjyuJE8VDi6LrSIc0QUyCN9E88GHCVpDRHSnow+T/BaljTii5Cr8Bui3
FarnX3+1EjuEKIuEtUWkXrVAc1BdG64pShHeB0rA6yvW7TXovTAERkFAk6yQtAfm
6wfXLihpJkQlddYigp/NbStfARrZmePLrjiDvuLuc3CU3g81EGUDx+aDjyqwZyQX
H6zZmGYT/7A0Fmj26lwR7N6ChQ+QwxYMFOEvGosgzN2Nec8cF7y+EIKVtvUQ61iU
OBAAM4KYMxvvhF1RGb028TEN2lISaSPvVu55inGHSp2bN6IcprSYnN0bRzanXW82
tgx4HfpfNw+BfNHZ42wtFAFdMrr8KHGLG+Dl/vQGSesl20EkwBHZ2VfZPnvZkUwN
xIxGHFa/glPu9EEJOUCbY3KH9SClzVo28WrpZCTLRc6rWV+kD7Tr+OjXgPGLdS1B
CTsEQq5ZoUWq7+Ks5rnhvGTrXTmMzxt6Um38GUgKTfXJdnre9jKFPKv0wABPyxDl
SEErJUpSGCgCyHp+VgFSHOtJxfIqKZZeHVJwZAsFYfbzMLLR9DwfkI+0cnv4492f
gPuAuTL10EEylWEV27kQHLNCz6oB4ddMpaPjzV9A8I44Gwd3cRWyyeVYwQ2D06Wf
GFZRwtV3I1vGd5aLEzThsdOBVxYrrK71Inw/vZ5t65DFGDRj7h9ZYm5u3nuCvSWL
ALoYuJW+/7TOFc5zYYros855nTO94s2NH4P7lT/bAC7wnGLteD22xxLZoCWj9QNS
9kTtDF709fhNmlOXZt5TKFpEd7K+c7ynDO6XWyA8jAlUAtBLSffIz4VG3rvEZR+x
zwF0i3jI6S1uii9Qqv/Bx6TgY+vTvKCfJ6VZ/TsG5UOVN/WTRZ9lLrKFrwZZAvpa
owuf4Us0XmHBXrjd3yMDLjG5GZMTJXTEFVFfFU29e0yhgIVCLd/tOZBHk1EYyWql
YYZScr/382ZjJ8l9vTyYzq00hFyywi2mKKO5Ut/3bNNCnX+1yEbEWfxbDiLYcPLT
7bd5YUTUepSXxmIvTyULa1S7k2jNCoWboHqnMS6KMSopf4Dcf+gfGOhGF8KUjJs7
GM++0YZZBtQnavPWzLW5nGgQLPJt6KTo+/U3Tzvf4GLa6p0fvOM6YjqvTgLr6/Qi
ZR2H5uX4r6Z4HmWgWsOc3JOI4NwuSEf8GRLAcRbwPz+bu6zL8zOLK8B1pS3Qtt5F
Qh9htdAtA7Dd7myM8Lpulv3JJmSvI2gsf1QFtyEtYbArzl+UE3LO31LNyKeD5rc0
FjNm51gpcuIeJEtKMK76VutVrbsSGo+sReK8/YHnCBya4C/6Ccl2uEro6GdgQKzk
CQtyHOPdI9tKnqJE1HUoPIrgBmWNhmAgigzGP5+uyegrChB92yC7wkcrJqRQh8dS
aqcVTXhoobYhpj1hyTHbw1L+0ZhQ2igjYXs3Yp+IgVuJPBur2WTEQ7jMpDTBue9n
sqgJib47MDO3hpxyl1C28XzZJ0LQlg6QehFaOGbLTZZHSKh4ix+6B4/UNTJLLrGl
itxvEYBClWn2uvl327TXaMiiPn9JNiQmmcFLUSxgv9Z5pS9ixbwNZlOT6STq0stW
fGIGhxyXaDTM/v0sTZoNZSHlmBp4P2wyLnD3+HTL3SiGQa79GlIttWQ3PkaXONHv
E7EXNH+QBeZ22QyAzEJq0ZjpWndXt4fN2pC5Kc6nJYPbp3wjMiXLUOfaAkPXPeUn
9QpafSa2sSu/cwTJ4mLAnEsX38Fkop6waAwc63jAtxDUis2bXravJbxUVmZUDf//
kKl7ZjMbCJrEOJOEtSO8qXwHhu8K6xoskOrdT8RJYnIL/pcpSAnEPLHb1tl5i9lP
gUyGNfOU1Ylq4xMYrvK4Ki/9N4DeBrkgfdsI1wJ8d8h9Hzlvee+9nwLi1qOq9yV7
xUUTP18IJ0IGoSJko8YbChe18mnZzNOvZWB5eruSPWA3Y8EM9L1nsmugp0i5X169
jq3KDljej6NA4p029/EXHMNhP3IdyUblMiwZ7sYMi2BYMntJwpWxLFGI0Tm26jtN
UwHxXSv1TAYBQU5njhRP7ZDEIfHO3ECz6xHq1AyCVyRVcoIOzMIVbRiVCX1QKBld
S5K1u0uuJYoU7Vah7gwErTbwBcWGm1m/BKAg9CTVBrogwWCOS9iZ9uasxxxcS1y7
KzgzzK+/EMWyYJh24C7TXSq5DOM2Lba135/nfJHa+XLQsONRstZU8WCNNzRvBYaJ
oSlfdBYZNUAEgP/y9hDXzr+/Q5upOVQV8gmNIMujz30UcA8lvicbS1nQcbC47u2C
HmWkBZ0W7VC1+xI/AU2ufTXpkefwJiYO2Xs0Mdd1Vzz38R25vX2AWv3SiqWqHPjO
qDtCF/OMRNaBTp6x/T7Alex5Yl0x+wYERLUq+GFKIHuLFmN9NQ3sVP12uCbR9/oH
i47sklZSvYUljTpF5MuQ6wVrgJKJHgpCgLC4ZRd1Ud3R27fqN7eEHNoiO5gRzTB2
zJ5EOQqpQi2kCFkfYi1hOTggGSEsY/88+pTOMTtLjRF8KXcqnt1M0EvA1PUdaqem
D4P9xJkwTr2Sj87uiVr4PLtUzW38qBW8PZ/XHMji8cMfYNH5OHyIrhBVEaokdpD/
315AN72sW0ywETeldXSP15O9HtFGZoU+tvjRg+E6PU1W3sYCAF96XO5jUfyxw0au
tkE2hJ5MHAskS2eU7GBBt6uMkPCtcyxVDhqj2H2KTJR15tuCg+ZkcBTW4vvTGJ3n
H0EZFiId18xwxaOMarPXwaGAXxZNWWX1orkOE2Kbx4tjEzWQJlituZEnbSFAERxO
zEGI0xO1T6iHM+1cWAz4BmWsXseY0FGDb3MxwD9p13gDRQmG58Myl24HcPDy533M
Vrp5zo3sI1garZ7tBmh83aZO/gqNq44773oN4a+OnDNGYW45Lpp0bGEHHbm14pqR
BrdVjtaxXYDC3oalXx0rD5HoP7OhR2qlDrU1um3JxCtYD662JWUBbYQPWa4CNzEe
uEIB/8JZWckQiKeR+IgyVzbMueIM5dNPWlySLWN4fzttFCyUHV+SE1TbmMN1Omuz
qpTtQVrFHIFnnZ68wmSyzN2uvayIHkcH4kBnB2MUh0BAKKcwdetOvXp/68fqd3dt
hG1UifdFZBhUGVdBmA85+67fAVBwSEr5oGp0fjFTMlGYdywdPH4UZkCy4kgUgRXE
qVmhRKhANT8QJjmH1wXIQPfMOfhNRhpGUDMJAy/nbp9auhTcYO+SMebFRkYE/+kB
qQb8gaP/C489MKpC0UV9weBS18g58X482hmwVTSKtxtzdEvAtSuV+rQ1dkomd75z
laqYbjR+lZRG6GHdODvHGUKc00Evo9yEC7ceZKo5+p42ZSnF7ja9CeiIaLjxyT9i
Ww+fvye+ATF7yfyIxCFPkOBc0sLpWPZniiqzDEYhmPNV7rDY9hcy2ugGrEngmrAI
Ukp1okJaMiJFsClk4VYU2Ykr5bkPAqgMwCrpvzC5K027gOpr6x6M6O4WTm7fTE6s
R8eH+t1/Y0V7F/Vj9o2E+a5ndU0terV9zavjytYmd+QQ8DOEOFR6X+uWkp82VVz9
lZlZgI5+xV26BiJoeeXiCyaEzRZie60CUobsjgJbs/bLYQf68oZYp0/lVGX8sxnW
dL7nDP5Xb24/Wt7eI7EutUX6TebvGdAltR+5hIhYYTYwRnYlILDH+LE5jHXieJwG
lF7cRSwEIU1YxqyxjC3niZ4ajDBbH38qNDr6P7z+h7G1zp7OC/PXkwDZrtQXgI5r
vqQZd1RAW4ly+dMuNtQA0LF6/qMgqnR4Zgp0e+lYtwf7sTanX5WgRh7wzGbCzrJF
4/VGcLFJrM22dAIWQH+w/ipMzAyayvoSVaRnpvZXCjftZ9Q6pXu2wj+Y1fHS2Lt9
b7KDo5cKdhOy/vxjVhMqezkX+qKtdMUM5OF8dT4lB9AEqUcUN46nOHz2/EIng7Gg
wC6N5b/KULWXyvtGO3E6tIpyYpM0YICBMrW2ptWLr9iZsN1p1GHdo3qEDo5zCPU9
+Uh1lIGyObx7ebOvd+454Do+xr7kAdirMWeoP2jpVAw9cispgEAf5R4fSVV2Dk4l
f5DE/yM6epr3R6bVAWDD9g9RAMe7zne28IDVb4KnY3uCp5SklvFyrqAFpLpn/LQJ
tnUmb4h6g5jvN7ggqJ9IHMkJX8eKbfaWUQpN2E5QxhDs0f+T1isuW9MDm/G+7lM2
89hklExp107WDcrQ6Arb3edCGxfhEdoavINCKUc+CnLzhRRLe313ORlDck3j0e77
YpSOoG8Zs6x68f5Z9faA7pGsUmU8XeZt3N6eUFqGJJndOU8P/78hVPxB3kQHqfe+
bxbi3DJymMCd/Yls95ZEZ7HMFp4mNXUS1CZX4lsbOHctvFyhMpJbw8kWQsfkHsNB
NLws1qqxXcQw6/ufDwnbGGQNwq2pa7gZbf5kwu9Vt37jwF6kZrhVnXeEWsK/aguB
gE3CqyKj5Xa9s+XDDMgh2iUxriaXiDWPTZNzv+fK+VsL2DNsKtHGOah6Cuwbfr0J
ugErOGtgYCTswHKs/ljZmgH0L4MsQ5K+PkCE01TJjWcjxzwL8rmpN2+NPeaJfrbq
uDOtCrCnRcLNz0AaqW8hR7vrF5UcDWQGMCuIr4/Q1j0gtzNtOOh6zErd46N8K5EQ
X3ip7yn67mw4a4CmLTMRDrdoT2IWLkr9Z+zQ5t8scnTkE7wnFGkNQoaUqR1uEqfH
Hkj9jMUD2884zU0WTQlC4dz0Km7u2Ax2Sln1ArEGqj8/SfrVNr1Lg5tfGBBee64D
ZSx527rfmcdevyLiBtU1LKLNqIIKkaFl/yZlMBR/zzZApdKq/26kusC3lX9MBIxs
TndVqrI2Of9fHPc4w0hSx1EtRXBVHse2CtaFm3poQMN1Fpqhza025wwto8qnOzhx
AXRqoCoSR61XhPdDegg4plk0Rk38XjbqU7CHcONfYWQxXoLFcBBCtcGcx6Og6ps+
fa6joEmV4VBZ4aWatwuujPMxPPh853RrtC016cOTAJdwJPWfk0Ry907wepIe7eKw
SSVGsvRYrUwQ0BhwL2RFDXuQEBtx5cloFR5WZT33SnuyJTnaIHWPQH9pz72MEkCu
wocLGnS3PoCk7gxWSzPVFbxMmvqZrPDmHCzDmF3Oe+6ktMD6UI3HcrIpR0Aya3wL
V0u5cg287RxJK/GFJMmwIa8LotdDpMLvRwnOjpbqn5sqhQPDnuKUh0Nu0PrGf+qo
90hWDDzHwcKAmsZRSFTZ81vWhAlk/a2qsVbfNyOcut7qQ9K9m33xnx+vVF2aX1lj
76vn+MpBSHbPeEyy7nSNAKWNEJq/JyUXvWJDcLPDQy3tbqeKkUlCkr6aYeNda478
hKTtTk6GTbYDg8umk4BM4L5VaSZK1HifRNmLivDb5hPbH2a0EKY56zJRFKWw1z1u
GeNLcwZJPx1eoTiSxjIhyogd3KKm/ta+SdEpnRs+VDh970SBSna+lZcjj47FZmpf
Kn9Egmc/jfuZSrfuXHsRHS5wLhflOWPFl0mRYQ2XWz2GpmuSUtw+TpJgwehaTsUI
1Z6m0L/GIqjSQCyPmNsil+jMmHRmB3QV0L6kXuC9Rjh8sql/4I8jmPHdrufd0Nl+
1RXM+1Lb72tOtX0X5n3hBOOQkN/Y4HsUSPIWrmZcYNYvOq64hnD0l+QQmnMCu6MW
w77ppA+37oXK1vRU5S1dM+YAT8oIOU7MvHILygfRdFzZULpqLi24LdNe/qu67wld
u/jQreGpYp1PKRHK93hlNbJ5ygCwg3hWNOkhpgW0FiNL4H8P5fg2vZiNzje+puv8
snyA5/Oz6HR40UJGgN3nNLeWeyszfOFtCaEKf3MbUC6F+ipEFs4BErkonAyV7iti
ZtVY/+tkFL2dtCk5Rxn7yzGi+fRFd4nEmdzNE0Bn+M2Pqvd2TBMhNG5ZBZvBe6ub
eA4w5DbJzZSEelF9/t3sA4t1zIEobATUq0h76lQkgUuqrY7XYN2TVXY8j72buDkF
KuRfaMNLItguVC8ITieomnD6Til+S2O75gGYonC4bN9iODujv59utvvm92f9C41Z
Rj++M/wjWuEJIldlFFll8t4yuPzIZAaxJh4XN/YV4zslWL7q34pFMJ90lOV2TRsB
qdfab0SF7PVWKatO58QMWWAMWwvZC6cCRSOzcoPH6DITVyUghsJ7/RlGifPkY5fZ
jWvBa64oYgZnIMvkVD0f2FXduYKkyrHswhxL4DS5BD7YvlvgdotYIeGC3G1knJyd
Cv2dhfJidesE7Mai3e4Hb/PM1wZ0Qu534t7Oz1UwU4VcEBnTWrWpOqIz5vkdHkeX
vxIdrgd1jZ0ilneYDoTkrRrqJ0ACls31LnXVROZGSGWw3L54Q1W03sj+349cwsT9
fqCxf491h8OzvfdwEt0MbZwbm0HHFEGueSiMUBzN+eJAeE+95Wrr3+dW1+9vqe9x
gUAopULOq0/yWQdwXR/Z2wWj9gIBBLNKkIWgpcAtwMooDdkF69KzGAvrot3LILXd
ldN+TTXq2BMTkwSzi5on2WRDcb0pJWky7ftVSAqu6EiYdMSrNRLem2jZYuO4gQrw
HNa1ee2blPxrjST9MnYB1WLRaKczB4p+AdLcjtNYrmDgIFC6UWGd+mCWRIGZzfxK
kodsWYpZXk+FYXHzf6zPfBXDVTjobyTksO8UQ0yHSNQyIkYmNuDe11FgC06EJHfJ
+Os3MocaGg4af23I/In/k1bcg+yRTMxUQ/tf0SkRLrKquDqch8vnYtaPoRier6Fo
N63G1aokyAg0sUyk5OSArDu9yj5N8i18P8LYlfZbdjPQK1CIVojorbLUXhIePbUz
X+LfTxJYePhfw7eiDAZJrhnbsmJcC5hYl9sqEYEWMu04C7hKsgSr94bpqSnrSAHO
YUmkMGrRImt4vqVX841vMMKeInH3S0cq9faheWYKDITP/Y7LmSTxFhCeQ1qakP63
Z5kiLIuw+VtiBEa3QSvQdTZR/YAq3lVtjIEO049aaLyFoFBr18BgdPt9cV3MEYbZ
+nwv4PSJXfSP7q3lprAzda2pLjU6RD04Zc/ZQbdXZFdHOwWXc4RXqPV636jyM+S7
jBS59hXPKrJNN2DDYwOyhmNYTeVbxpieEKiyeHAKZ096/PpTRDdygwAN13wtz9bW
DLTRQN2ur1bukmS/RLg0ptAIb/pgOWhvT7+WwRVgBVXoaKkDY/L8d4Ylq91rwBtd
QJ+mfKii7EqIwI6EtD9E7mgGdOPjurTs+8msvW3JHLP4YOfLwv0uBH9oH08gcB9F
TiL/2n3Ctsze28SqHdPvWoxAKZ2xDX/upbTUbTpPTV4ptsUgFeB/tnM7AE+DFzVt
VRvEtPd0tVCH+sEzOgxxujcEwuI2XIEHALrKXHBySp3Wdca0KlTM+Gzh9Ew1Bu+g
0tfpnZXn0yn3b/pVhnrZfwEcCrwC1vlyyaBY60b0vG9OWe+vGY0uEb5Dhoe4K+gb
SjUSwzogkGi0GY63hNmeqMIYVcLuxW/6Mpuz11cMWmNqDYbAPJFUjbp/PcpTcde/
OGZ90Zv6vANo13pLPxQKV+KpEmCvA3X6ZO3xSezY2BdwCAuKwTwPW6+27KveMq3d
9suuVAPAcArXS+h/jhf4q8ElPBukWhsv4zbO9FQTfnjJSfKHptAJ29Jer6Q+0uTY
QabB7MiRXEwKDhZk3wzNskMny43t8709e7GmVa/mlmRyPCoyu/XHuTTWM0PVXikk
QMiBcTjRnufz23P4J8aUDq2UT5VOJ6YNLI6aHx8hQxfzTIoItsvLWXm+WAh2MjEg
Vnhz/oDkXERDfKx/u4aV5E2o0Op90j/j9YFrD0KaQ50b/1wjJ+E9gaWkXlAOIFkP
4SeMaWz8rbpDctBaGhb4qzuU8Nd2EnnviIeJ+Ace7ALcpL/uuP2vhxkP21IY2JtB
b4nbCVbjU7KVmqJcIeSm7oAPrsjtWhhAe5DIDTbRB2PXSiLBxV0tNCxZ2OmdeWF4
GFw7G21o3uQ0lVC8Og1zKnxGKhmvm3BYfWa2XcsEwlGUFCSqk5XF4Ne0nzcJgkXT
gdOxUhkE+9joXbTDEBrh3Yl0NjScc+LwXzeSx6sCGkU1/V4joZHxMIfzSqb5ZNch
kOU0N2OhRWemosspE50votmPhMGEhmln8PhZrTQz0fmHoTdmQS4GB5MG58TXUwtI
TirSOvk/d8mZbOo4y7rIT1hsEsBuAUvPzmcazlBc8KcyOQIMYWQGIyfKchYT7G2R
dT+EVWlvm7szbsboxm3jWXXVuaKBLg8F2BVvue9wtm+Rt2UvxN7gS6OdWdACIhas
GdnAC29vktjvzA8IOl/8tGZoJmd4UHkymNp8w+bzOPtvAQSRKbF5Qq6GIVoudqym
ywDRMI58T/x4aWeL56Nu28hJ1ZVuBcZZVJCxrH/I58EER+njALtjqLI+CGnyO+LK
xKdmx2Q37pWAzA1lpeawru1llMt7Wr5aGBkjWEIQMmRLN4t0ZFKOnFfGxjcZg4Gz
rwemxoux0xngXnqAZL6gvc+T5LaFeDXYDRWzCEARjBOQltPh7bmpfD86AOocOVrY
gKET2gCmorjMl/Fu11ywTabATr1p9vTypqNy/sTykku3wND3Y1KIg5/8w0O4G9jW
rWkMxdrjfohJReaJS0ihqVngXNbBwBQO5gfU4zgHXWxatKDg6+LbCODtHfCLq0v+
mxn3SRsSMBJM6/488x/lvi4l0lb9iC0tHMKK6x7il6/hCkv9ytUumzwvkgMRijYm
eDcwg8waSMk7W4/re/UReL3cCA/8BEHrFcoFhCoP28wfIa6N4oYYpb1eunRtbmd6
UVV/vTqElr2Bjb5STJOxJli1vBa83zgcQeLhvTSVlRUroBfFJBLspodFCRjcxPFs
k2otC+uT/PClQxM/lgFoUgUyj9/d8Vh37PMUxugrY6T7jJjYAaiRZ+SzITZ8Va0X
JaTo/D76e3I2cE1dR75mHt1AgIo0ttQic9f3u9abN/xKwt2xs3ksIQ5qRjHQ2we4
Y7DsKDmz/Kl3/jxqPCPopHBSZRlHwGePheFTLkm6yU+thCjgDVr0n0DLDZMlugU+
dCLR+FxpDuvJJj4HjmTgBrtGgTf2DLrJwUaIxSRMr2IVX/0muor8x3jSJ5E2yu8G
kgJYmyRhOWOe7SKTB3nrrY3SlM/KHrAQqY1fKCpZB+ckLxbxmkObAvKe5V0UR6zf
zrijvEPtDw5w6UjLQIcx5Ss+quZ3dgvw+KcB5fMp91LiYrHc/x1TOxGm6BNdAMQ5
F+RwDNz9kpS8vZkrube5Oq+bLLPzWOGr/EuEAiIs2wugGEi22TiFGVZU76vGVsPl
DOqmqSpMi3H32JcUGoNJbzF4zAKBVl16OZ9PsvOD2LItxP9lCx6nJFBjI6Au5I+o
vofpmRboptnheVAhlOQmPNHz8MSecIaolZfmpnzLntYjRE15LV6q1EsNuyA0AHPs
8+bKbUusXS9J85pYtVxz4LwWgg1aPQIrV/4Ri/aCHEBLPVjd4ucUIgPYGyO13DVQ
y7Mz6PopBbvqKL9VPWKIGdfcqbvR6gTsufb9RGD/7q0ZaCsMUjrYy/j5Q9Qs3xHJ
b0OTMFcvMCm8dpv9pjqiALR4FzGbaRN9zyujMMqdM+cEIMgGL79grEXlTg2Vsc/L
m6fl/P0ukAoaqFMQVw92TrdH7KObFvYTODzClF03KbsqxGjN5UA/hjcHQqn2K162
sjl8yOP253f+HF5TgW0ayM8Sv9cJ2VSZ82+Lnr1P2guhd+abwdQ8qNncUU9HCkJf
GLlQ6GvEhll/3XQ3tloJxNlg+pcRCUfETJqzLl57IY02Cj6qh9E0ij7v2U76ecFb
gqs4K/+DkT4Hrcfxj5jWfTQgUbL8iKQMeQxjobJBvd6cC6COTt3FzgiCtxXhhxjJ
nvMq7Ub0+ZEoSxQd8AxoszpWZJJQB6fWvDPx8pWshJOHSpfi/efPdonWBasloejA
C/FLwAn3HT8yu+FbvUWZG8jgBb5nZd3GvS4f46/iOSF8Vto1UaJ6Blak+H7EIc9X
1FzeAHmcdcvw0raFZkbrZS70ieyXAzP0gfEa0khCiMPA+PzmMtZSSJjseYcdUhry
BhT6yaLQjiUV11J1GYZmi/BNo2Q4bF9zgmnp+41zcJwPSW0SmOYUxiLOUTIyzw6n
xVeOwdV48BIbFzfjf+SxNcRB5B8+8oPpoXoUOW1pRHiJsXPWJ6sKnVpwbp9oFhYY
QSw5TGq1pIDOKzYphFsAyChaL7P3TH8GDmYwvisTpMtXEa4UoF4jXFXZ8wXsea51
609hHIuE3EBvgZeCpihfxXPQWrIqYdh7vDaG1XNSQ+ia9B0YEW0KbLoJRPy+BCKY
Z32kFevXXwiQm0eryuYzTWhjxc5NscMmt66ymZU8fVsjeZ0xLvp3Jtxn4LW0C4QN
xXri+r9uBuT5JcVVQxLfyEmClrqvtFQNYA+3wpIve+ESQDS9+uUw0qTfL/KaQyrU
wFJbqf/Hx8N3R+AgWYJbTuWINff8b3QEi0XLELf7pscD2mVDixeKZNvBL42sb8Rd
HhfWQWXBlQf1kLAbvor6kxQp+44TKgiUluxVbWlSArNyH0GNbrPlMCAplqUaa6gu
MGo2BoF99pT3ofDVY2xwFAzmLjeKaI9uOJ9/syhSyocE8wlfANv1RuEaaQO0bDVx
+j6JFGry4QkUOZ0HomIbi3DFWo24erX1tWQFRRISvASYhVExZwssjYMTgWFp71KB
ac0sCri26KVBGm2GOECRNNA2AlkOL+GnzIltxXbv/irVIQetyoQSMlZzxknstFh1
p6Pb4gUxDVA/QDC+BdSV5HuUpntWQ5KWaLssyj6pR+9WjIJHBLXWFjs+jNhfii2A
WuZf+hpaqtbyEvPAn5gnE9naa+K9asiPr8zcqFJSXDCQ0c/Wk0VJvwzrL07a0+1k
dLM+y49CeoHAi7psnxK5gq38/ANK+JVB+CuEYd5Gio9BhxOhRf5ImvVF2tYRZn73
guDUIBuBcAo2Mmqu9IAcUuT4eNUGfmHeyzyUW1+xULXYW7BR1MeDiFRzf+8Kjb3B
IA4zwjoSeQKnmkwK2mAy3BPw4JPn+yO1f51+Tg9TRH5OYtWRDudr2xrPjrRrzkws
pfX9iJqv02CVRDnlnxN4O3HflDaX/zgJngnkdE6etxM5ymSeqHJAuzSelPUdU/pw
3zzzWZLOKqPRRC2hz2kHuOjEhIc7qLycZjR7AMk2fUqVrA07sh1vVMqr5/sPj4Lt
Hp3urnfpF3ssvnNq4b4PODq30KHVdmj7/WT5QkDI1FPMLEZS6rEpzsdAfrAY4pVh
M9GeHLlHggVUzSEjEMejImJ0/Vg5s4oiYXd0QGj/iL9VG8PkRsdW3SNdnaWqqLuu
KtyyRDT4axGh4qzj4QPjK0Jr1dzsdE2BjGgcgswogWHtU1n5NiyG283cFUpigF38
7Nwj6DeN6vjVRhUdDqd5AiXbwYrioDYcDy8doKHL18FeJlOxOSa406bZdUSStEkP
Mc4anKpEPXg4GCI7ezX02DG/T5vZFS0K2b/hAa3rAC/zKBKEoXwHfuChUEMYatFp
aAd9iDMEYxPXex3+NbOBqFgcXzTLtkyJ/TWZCx+3/UfudjVe2PE8tI+uGvn0Dd9r
n3NxK0NlXUMjdvn6Gs8EhjFZqJbha+TRTBuE+nWhcgZ6s1ew2QDLbjn3R/KH2sf1
4w74euJp3m9g/zyXqNuheESICnNCo6ErZleg3O8nKFXmHL2d1luCTjywkN6uOr9J
INg02J++6XzVq2vOWkpMf8wNzeKoVo8Ltu8qy9o/b8z2+4NHq2FzdvqFusuL0RfW
JxNjRjBwILRdEudfEw3hBEVDk41grJarDz2iEtVr12iOWFjBR7AJdjeE7+Vj385/
jdRvwOaPIDcTFmJx8LDiBYUyLGIo+GZ7Tw9dV6So99HiBviF/p+UXmz/Kod1GSYW
k9qYQ8++mwr/ay1E6GruVmVq+95/BtKkyTLKN8q2CxPavDDmvWW8lgqPodCgzdra
34626wkwZFaqSxUE91Af5w/xIZu8cNYTmnJUmhE5Vkdr/oDalwlDEEFTh4f6bMAn
FHSSD3APz6egMnlkO10Edf1alpxeP+5VMRxjOwylgVeBTWZlRt7kHhiLRY2dlsMH
32YQwENc+7iY/reFMKgkwKcc0g7PhMe9urKa2XFE8pSktW50xFWhH9aNqU+6s7e/
b2TQ5AP2cT5pDpk33kQr527cYVryygI9ZUYaq1HCZehQOw5zumBcssAXBO/a7evd
cXLXkKmoWWwMM7ID0nt5dTTEGGONY0Ynty0iSgEM+SUz+yXNMR1jlkEubTgipXKU
l4Er5fmLxhUtGzDUY4EtmrRjVU+Psv3s1jvhSUp6UMqplVB62Z5Gf1a5udZDyNNa
9xZJDNSJkqzKVzUlI35ikuacDOVXYCzbE0XmOEPqFniZOdpbseS4UWSRoJpkxBO7
80y2dFiX53ANMdc47TWUL+7OHXm+Q5D+GHPBvpCxpCdXI3dqGMP50Wh9ozU3I0m4
dI69HMRPaJP1Ily2UWDvlErbxSzI+5o4CrP45KnS0nJvWxBswFj/hejjmMsMGZv9
MO6DguXAt52rw9boMaB7WrrSp9qUSz3RHPaFBOYgFedRQ1uWAfWyuXrwVif6Vd2K
jtef9E4n4CYDKFuanWIslkbBi3E3uw2wtR+E9cgH9ZrpCmYBWkoGIpOM1fXAgdTG
VJKCPxNCg7k/hVTw0u1RQ455E1aLZnjULAKiUnXoOid2rnxEpxJUAT5j9nekO+Gy
9BBAvDM99lksrba0N43597OQG5YVhbecK2JRWzVqjqqLUaOQ1YHGUDlI23BJfDCW
Hels5+44lhMJnyHMQKmUczvzrv9zuAUSNQBPPr0lNMD81BPLx79RQcP6cT6mFHZp
W4jL8Ymi5gfOEGY9yeG4td3vU3w1wdX3wFJWqvg4G0/yUSnTOzDmAPpR5zgyfba0
4e02Ff7qR3MoCU8kCXOyl+owOSf51uHdQPPpUUZuDxPCZEu1N6ib98QUKWWXA0KO
iNyqn22fpqxNhXeLb+LTxe3pU5XuKADfyfZFz5Y+LcAMZuCZCJz0fw8f0BGrjDdu
FWTd3AsNhE8D//30tlrC1PZ0LO+IWaoKJlmfflS4ONJ0koFpyJ/wX/iCoWPgYEQg
psI4LVg4NBXpTazhcopsagfQspO4CuUvyx/6kKzglGNtBDsHG/JmFVGRwHdR/Y3B
4ndl6iJZb2Bdc6NIp/yIMFMntrG8dYVUh+/FhbRjYmRPCkPrKQbazx3B2uk0VnSt
zJ6aQVUTYjWOwq23R0zU1TYZiYukZljTVAP+w9cOOrpMMwRCMhU8ldYU2XVT8Kye
T4ICaEPPWnpbQGj18CpLcEdBA885T6mE9V1gJw4U7GMhpszb9ZcV1uDX8V1yWFxK
/rzjA6FH1WjRuXgGlmI8icefZwCF97weMoNGvoOPVQr5AaGOX9130SAh/Zyr2Z4L
pqWZlsP1qdMv3U9sHeOLieTBdyAduAv/RbtzvtaoaP1vggxrby+RXq5v4ZIfRJwN
tj8jSMUqqga/d82qS7/sRNObLPtIzinGH5aYPZR7WOBbK7YyWhjbgkMvD3BTzRon
GXtqS5dppKFkpZn//m61sVX3rH7jZZ+ELL+R70qx/mtcuk1OZueg127lGp5lXNFA
1NT8K0ijh7jWpOOFO9j5TvIroSNCthpUNvtjUIux39uTTfNCWrxV7TamYl91uHK7
q1PA7xkKvapntFlDD5XecxCH6x/bTPA95dy+guNdIPgY3sUS/lUkzYgAbsudG7nl
sFPgLNCk+OiTqCLggvtGtwThIodlpc59cE/pRt7WO4+kw1wVEJziJh+XegkaP76s
VOfQyQ1ivWjnLQmnI9xHdI1ufYgY26ARIaH+0d8s4bkl0lxZy+eO9bWJs0VQUbx6
IjVyMTsOZoP3ztkWvGwNl+2dZibyXBDv1mcvtyJv3y+GXa4Bf49wMjjGK75qAVHA
OiLCxbA0/pg4yoBJHXQamaQoyfFGFBZryVE+R3HLhQXRFhq2OUAGC4wOKdINA78L
11fLZqrbrbMHYbGVkWVNcp9RgNRYWxyy/pMb/TwvOVkWfXxF2nHgeTsYcAt+fiaG
+zSSVvmogsyPtZ4Kuz11msywVAglivIoNVEUb/hXTbIHiILFw4LAJ+repNpD/v6C
UiP/wJnG1HFksOkAkzoX9BeiNOb1aMwJf4qQO012Qq0jdWQ2MRWyvtzqvR2LSPXI
/WZk/P/gUW2mBK7hM1JGhxmEbD8Vx8Pf5hyIvoRbbkn7+mp+ntdWif+H+dCs7oZk
3qZnqIUMe1h7Qycu7NLHIW1U16f0DHszJALKz/cR+1aggKPLOaW8g4kksdDRii73
tXdNzfwjHkm+kOBkvKO7ekwoJiaUBNC71K5wUtY1O6ksgWOgiiGmR2d8BZOpZLM7
dvSN9qYOjaDCeNa9HfanIpyWGg16wIpHCoe3rbYMdX0ipQNf5fyYpNfazEoUVJ9E
a5gHwFpH/VvjG2IMWDJ87Pu9aiVgSeEgVzxi21JtVHHo8Xc92ZL+NwcwgpmiTJhE
gGLQFGotWUykz3tns3o5PfEA7xNkmv7C1rEORj3pZT4B3GuqUMDFPbjWOw32DUoB
PAbpTYt5GcflI6FF2DEVvGisxhQ77Y9U4dd4SmGGLMnpMt4/1aZofSuQrdhRZtXc
LZHY48sete6vrGtJpdQEFGP6GOjYN6reggAhMKZtUT8ISP2ZDib6Lk786/0iLgfi
YEenW4UnV2KkXC5tc6gZZ+ytJI5an96wSyjTKzAF9Py+3KLBJdkli1oEg/uLwDe8
bFKhJSiRwv8nIaQbEbAS/trIrrLXjU3k82/UzUOriw8Ka51GPTfuH6Vo2w14CDxR
43gHZY1dKQgj6L2USD5CJ7vcxGZxDsEeXmWdEjjvbmFd7KTE6K/Zkgc9e1/1Dcd/
TGDg6RsrPQTAzAp8JI15n01Wdm+TIcaFeXAcvXifKcNnNv1xOS5kPyW47ZzxIcjE
Feu0SRatG9HPPmb44frTQcG0CwLJzmqOR0PtAkn1ft0BjFgW16RSXYHzACtWSo+y
BqlgSD2rXpwf1tTEK0PwK9DsjtBeCEAKLW1HZhopXyl/Kb6k6awK/YuXuF8c6Wde
cc6CQku+GAYyNawTpnOA7OswCFzm4q7xdEG+EkFBHV2vm6Nzj7Q3H6caZexjoJJF
ejnJs+hCkdTolWRrLiM2OZNgyfovfoYTrK35wxbylCrg4r7nKq7mBB91RTrWYYrh
C59tThN1yFlMyyzx+wGDudgB0UuoVMZp6TLN0TR5vGtvkF+/WEUVlfZksypGVjSn
l/czUqJeJtb6+5TzyYnDPTH6ltpzV7QgWqNFwX0DKBtpBkNDnAq2ZqTSmrCHgufy
KGTqLcBPUZBveahNh8A/fq9Lmkol2pZtLUtwyFUlfX1kginLbsG94IqBCKT8SDzh
76ghOq/YtD/yNuYl32IzBqlO9P0/dAkhl8VXQ5AFbhwPnxnNeLaFYXLduCrG3dSS
BWP9zD0qoZwV63T7Smo5Y+gfkCArkCUIncjd4x9YbepDWsU7cCOcYjbQjHV+Taga
ms9KM9KlEpxYcubunbpVIUvuFoLuHZBFjQqIEVZ1odowltXIG59BfSSiytt+DrL7
+DChqVHuLfI19RxGKhO2FgWGpXz/30o3CYs6EU9mWQA9BlmdmqVbGPh5OHyeBCKm
cg7E21rHkKroDFWIWFAac/qnXBZmc9egXsOs94+VRch512dvpGX2sjI/oL9cwVHQ
MbLua1EBBZa+ehrDlGVWylSLFsQ6iqKeRUbWywnryerbI5//miY9jNlt+DP9Yw6P
5bYcVZqj4DpfJexi40P/DAQNa5akrmiSr6+Q3we+UwU6tX431bM5zwM/xuudaxxI
xu/xy3JbAKCR7d01snbd0HYu7BaFK1/2RLxMPl/pCqM9Y/Rny7I6yItLro/z58Qb
1Oc5LMywNgxCLF7B+EDUD7qBTo22JN2vT2+t5zDwFLyquw7bJTfIKSGban1f3MFU
CjVlIo1xQzMO4hn2R3F9b06VZBm93bpbdS/SM/MXutHjtwuIletmkJPgxDGdXWPf
6mD87bM96nvsLDNG7X6L/s/+BoQPyxSKyvvy19vzl8oecKoEyC4gG5FtvJuEwy0X
LX6ab79ISDnb/pCRwh/AjUEzY89SvL2MEovvd/ehChJeWm2IJw1VKXJB+EQ/ho0b
g4HVokcmsZX1LvHqeAmnQ+eaPzKS09fbVUxEOI5Ybt/XEYL3UJVz3Hc7Rq2F4bYh
WtbBfGLq5hStwaJVEhuEUq61lTMk+D3VJ91caGl/wQrb87DrGRly87F7jH4vozKf
bBbeR7/9jyNva423kZ+yCCOS9Zhwi18jusQ8ZsMFP/8RJm5/WV5U2JEEba9PHmIx
YB69/BIk01ccuhXpwrhmUSAGcH5zEdZa+IFnt3DaMLads6Z/kffHwNlmiJ/2jDMu
y3WXlwov9HqUOaRIZrNknNuFUWnKxITGy2eQGcMxLgvhCeF2HTXMkW6d7HpYc6p4
89OODZkj4gIpgiYND24aTzEuPcx4ElACqKHBNZOsUgSkS2NfbctP6F0C6V/1FUk2
fV4ab5/bpE+cLHc+wV5bJD6Z2cc3JpAiAiN/Pr1znnpKjwMJLtUC5JEMDRZQeQ+5
b0mxJlCnhSh0BIS/j78634J7ZUM///UgKj9IaeVnJSnVwK9n6TxVwVPl4579txUQ
aPpde6Iws4ui46s2TK3DtLafKKQw+BoGjH/hRoJbxOaPMsprFNlM7LEvk2dLpNk8
HP9AUsNVKF9xrKJHk4NNIScc3piM+Ze8/mYASJuEqvbdwjLHFpfwYBrx8S+yPNF+
msNarDKuvhBV8f+yVNmI46ayVW89iJyPPn2CdIk8oQqgdQl+SMUZJSXTnH2Ky6QP
y0/bvjOMmkoaa+AV0xhoT9jmY15apIkdjV0BQA/CZvFjEQFSlUJ/JIq46zGGUjKQ
6gJSTxArfYA2cpD08E5fC2GvhfFdGgzWhnKaWkT/jcD1EF9/gv10QJrdPKnp46r/
2eQLjY2dWTgy+HFn6gEgCcwvJMjrB+frReSzyMdaGKIgJ4Vvlcn3/IdHXJj4qKT+
UPdvYGVG3+Lqe/5HIQYmqnaKXc3wHLnyJk6mKSHO0Xfvu1jKATvu1CyeKsTfvd4+
mB9wRU5iHlraoiavt0oGJNBVDzRZfy8Vz2UBIrPdqXtqWrWLS8U/VtLAWpRbI0Zf
oGNOOk728UavPynxHU+dexJnbdsNvIrFN26LwGU8ke9P4O9L4FrA9LJbb6N06VVi
p4KV14MaQ7pA0TkxUyC3CdVNYv7OMY3d0TL70vPXZzwBPb3hSXiZsRogzkfKasUz
PSPKTEeZlkTf7F3MLWWB9Z5iLTUnQVkRhdLfhKX2kRXTW3/UROqCI6NEmTAqDzJ8
DHhr+fl+M1+wh1tTImvUlVc0Hl2V4NxVjlvXCIaa8ZbRA1Hde6vAsv5mw4WZ4Z5f
2drdMokU5zbCix/qy9j9+YoKEW2Fqq7zaT1zWrDNwm5K2O0Si7CUyCNCeTr/3j89
HfkAOtIpVUNjL9EgjQXnodEhHbpjIauRFAvN6i4duCP7qBL9rsOoezQEcMC8qGWI
DsfB0fjogdRhfn6jNPna4NayqNRqzxButiC9LeHXRXUMoeTHmPpMkmhH2UbXcCQ0
OCwZwBrKsJmaG9hJAKSz4gq8iIP/S0JI2JkUHgCAsOw8S83vm/m0/ZLf27DQ7P/V
n6BRmhViRTLG9XOnkbK6A//kGs6NRpHbMhReL/4Tpz+fSl8l48zsYYdPLFYn+AXt
ey/5FOmjO7SKco91sZED57OGNT2th4xa+xg4Speb6Hlhac7yAUaqmo2ABC1eNrW/
R5rtFFvllDb8UE1t8O7+5snp15E7FBDlxvsuTwxoO9hR1tt4ykj9z0+w7qdET+LZ
dEDO05CcHlRNrAyBHrOa3d84rs4h+CORlrGqBCyyCnBZkE9UJWKwNIKHXwPN2RyL
NyOXOdpQT5FoDEm+yc33TFf58aGNYr79sqAPgVuHdop4HUUGKUoRzU90zgF2Bpwm
26X4+Bb9f6zKUnSABvTpQWMlQm75+95tIR6FKJpU78PrXzNg2IOHX7F4ggW12xPi
1DpMmRO8HXBjsNpKn29yD3dOOTpcBwPE3bldkZCKn1VRpblo6engyiFXJpK82WPS
pB4VY2amf/Sykh9CzEOCLCZ7nUJxn6ecqCh2f92MOLYm+hyWqPYLrNgOaerdMGQ3
j4d+EgvQYDUAHU1LOenD8Lsxy5OCkXcXuLkTHQLSFk8fbFO5ToGszDKJonWamrBq
iO568cnog18k0YObh6QQ9VD6TXnOI/scZPATSa9cSfVFPLLjOZbLVkbnSulnpbmC
jbQpL/KQ5egZFqCWEMAD0ns7YG6HNHzjcoG4LTRftHxssg1EvNhHwl56CHJcvsd2
/iDvDyRY7DD9Uv8w5f/hYwhAbqn4N15aArcGCxHtCxJ7wM+a/PtDsRVftDqbLMRh
ZbWAsONk9icsg0M9pyh/9Yq52n6zp58jqyfJLppkaXjIW0O4IDkbi/G3Z3vig/yr
fse87jm3TCCYLZJ85em0Y7sX+SOrRAyFAyVNdcWV8mmsiHr2VlT5N4cbTZ3DUM0F
TvQESpwhCNtKLxgGVAJBt8lJ0WfpIb1KZAtyKrinkVcZsAMgNC9lSeIbdxUtowt1
4PerXYjIFv//BBFqlmzjwLcy3uh4ZA1n0gOKVF5OCZ5ooyXvQJY0kbKvvLnxxz22
jGKccgqtUlm3Oh3N/wErOuWpnlsRV/wsk9j3bYB83Xed3l+rp6GgqTqyNxfRzmzM
582Ygun57q2Tu+HzKhEmmMEYeTUVrPlYEqKMC0o4cnsBZdckqjP4Ol+az/1QHwuJ
85iqAFwk7JFSnejdvbp/tdz/Ze9TU+zf/7fkm3rhufT81Z7kSRlE4WDH74zUlPko
6Jj6kg4/PYq5jELExOJeECYPujeERJKBTEChxVxFtE63ZesW/cHYAt+VYzOxoWLT
Z0imrvE0yzLJWt+sW76pKYhOC8v0PxFXiSsaPYrAiFrO2+7l0fKM/F2y7VOFtQWA
0glvCuf3UMA08edUBcP3l6LOtteIKXadaaXCEm7+O+EDAkSv9xVjaSEiEEeWmpVP
mEup1CHRFjAAGoGo1CYF6U6twjtFj3fLKVIStS3Hu9tttqY8SxBiIAchq7JiTu48
oSW4ilXJYkpuJeLFoAbK4R73YiFuxh1mM0rfuRcicZ5WLUs9RUiA0m8irozpK5Ne
IMldV7bjmPWNsUcuqJJpC9w6qVK1wNQw60V83u9ODb21QqXqeCYL8+IAOtVEyj2B
O6vKAUgmGjKqeAUne/MvMFz6bLKIBiYE7haJbpBHhP0mgYJJEeBIVegeUQySY5wj
Y6ez+b6uy3Vmt4eOmVgMddL+qXZiw0lRZg7BxUFgEoUniDb+zW0abzMnaRR7GfVw
ZJKJRIGE92AEWXhD28jXkCL2pMIrZakx8GDJsMZIUQJSwrRVgl28do3PxXKl5LZ/
osUXFQrJLykPtVBj5riez28EOtZDtwUZ4D9AN7IOikaRMIuJ9Ddmm7NmiYafCrE3
hTdzAk8YylbPcRAJQX/XrVrdcfXKlGNq1L/fm8jklmJmH1YdS+I5V8l6UajJ/2wB
d5MXZ5DCdEQ7VwtUl3pdTW69O7umWOV6fJ/GqhXAhuP6ZBjsM/uJrdJaHvHT+3HR
6ykTc60N9hV65hJtkZNa316dlNbqqFawxH9AzEbF3G9RU1AzSYIY3rK0VFSK4r8X
mx/DbphdEdLbPNEuLyQxmUbGQ8HHz3WLaCntlNgGf//8se3tVnQUh5OEcPAz+c/d
zJ6HCgYGgsw/k2TbtPpo3dnu0sJ8a3hV1ENshveaxOswXyO5XaGXGr1xQAvNz/pb
FUDSIOaTjkoVvEkA4XtLtwnV3rXaKxSAd75bc1ATuh6Jf9rFWp6aLyKBXhkW3hlI
OVvmQkAM/hIu9ol9TS8NHg7XS+73CtgH/A0Vt+QT/MXppw842e1J9H7UnWYdj+M1
EOsxAUB+bcaKyhzZWgfbbpcUSYVXjuT4IW3Bs2N712Nbr6K7/c5v6exAjOxB/1M9
v2C+CMPFAb6Hc20x3x6panakyqFPjTPnBsYl1eQo/gdb63hLj3zuL9NDOaDVZDig
ZQZ3VvLQupAxPwFUDH+B14t3URYdDIWUEMX7wkgfaxSBVJa0fp5XRz86dzo1pZzi
SKHyrD7Y3QyOn9XpKc2DGEN5MczzxkCo17IEsOuVdt7ut47EplMnft7pRAjcDIiL
k/lzYQZxL5prn91D4m40mWbfNnsaWsJTY29YFF0LQdmh3E99mxVJSMMORYfwUgio
tjiZbjwO0kv/p6YvlGfRa9qXJBg7JJ9/5k3HqUD+cEbslZbVYVlSY7+FmhxZngbr
cep3LcspUowkIlMPbI22f7cqIGS5kd/OjKHwM43aMvohXKxPMfVI6jkreOrUNM8G
UPN8KmwOqlT36tWbNQU+Xa/glc/WqcK6E7RJq9AA1nnCz/Qi4ODtcrJSsppd3v0B
qT4JdoAOTpi2XMCPbqs7jP1DzYaP4p+h25qmJ+G58RPtRzVXvMTBn2kl3VeTjBSi
zFSePm/xer+auCPa0wYlGCC45SCShjxe+oyEhDR071MTnM+4cCH2U2jQYAvbcvT0
XmEv2DhO9CTIqLW+G4PgqOqvVk0p0Hm5HuRjDyawRoPW/xGumvY58zxfry2+Akc4
S191G6PR2psSOmlJSOjMW0tZ5aDBkXX1/xA/ziI+L4noVgNBLXU+yw/eAw+p0YoH
5Zin72cu5dCT9htsWyk+qGpZC99+7W+nc9UlYJeOHmRS51VhP4KcWgn74NAW5Dwk
N3FHqqcJmNUF99Myms7Oi4zpitWgw+P6W3W2WBYnepEQyo2XU7IsCys3Z3XyASjl
XGx+n3vSXcmVg6wOa61r/dck0vBVbjmVNbPMTbvNrxDFdSQKzK02bb0A3V/zOygo
jGCWtjPmJxZBiAls7/Q5dR9Yoo+lSnryC9nUWYVBUGC1OB09TNvnCXZP2w/yVC1A
JirzzF5oNoGEGy9rZOGhRrDONVDt0ySGwz/cpawWvmvJqzAGcv4mcTLnVJgwKfft
l5gUyW/lLSsrHRgzKM6yxVQJk4M1s7LugBgN6wNatD/np3lhnqpGL7KU4VXzE+H5
SbWMjYRXf6XaQ2cFeYMsFjmGvLU5cZBPF3tYwfAwnqIDuRIh+A1EwFoKOxnBvbc8
a9uGoMlOxaI5XEhbX+xy71LWd5O0PNvpxsmgk0/5Xx+/kY8aAWoXfEy9SxS3fBTL
Eo3CzYIU1S/C/YDfsd5E92vn85Z2CxniCN2z6m9TisGPuji6H160E8alAPdebHS9
UiofGv3U3OJQGO/G+eGiDqtGzZjSWIeS9xRYbt1klnoFPk+EzZPe2fJgpouEOeN3
bVW8uB6ZxKMG8A42m1nXdQxkCPUFHep1lC3XyyljR/qsKFQR44hHGWEpj5Qn9r5P
bvNjDnAguCHXIuPr9/7y9uFp7czXsjPHATATjT7uWwDsIwsnnzUnqbA/yHTQWHnw
rPa6xzAUhcTCyoCoNd608vV/1pLkvHeyIpsx/xuNQoMKfQKjq+BNXvIPCSBBbhqe
0kIkdzFc3t8niZt/U4UhWRIisHDTJF+haNpCRrxf5F2+y3r4h2/4bhGwed+C+baA
HhSYN2AHuZRKCCqfEAxlm+ZhD9JmYL5+ITx21ulE/mb6tKoMjro6yRC3iKi3XzgZ
G+Lpd0mr3SeUpQB9b6Qny2ix5YSBxxBBO+aE4Nl+B2HHVOPJ9w4mMSGQOZW7jI+M
m8hN2dSsJHdyVf073NDBXcmIX5Wv36jrifj0US2pq4MHLzVazWiRQya/efpblPC/
LfKnjk6peuCrWCfhEX28KoPjY3sbvifzX3oWmVYW83a2Nz/5lDtOo9V1UApu/z2Q
ics9P2X62iLdCTNF+a/OcmR4d9/iggdXIM35iCwgGVbidf4527muX1u5d2+JgUzi
hf5rhi7WFTM4/OikwLuu+yYHMh9w3MLxL5gwyDoValET3unXWAuxVrySRB+2f6Pv
PVSQ2RnYXtOTMwKcLvjCMhM3qtmojRJdbaQVYOkamdKZ/gGaRl5NeRwclGxOJuTK
HJ2pOsTrgn15m0a2C2E7fPXerlfZYDXPC2dbfNbm1D6rdum6LZiW06EK1ZGpHjFR
W73lc2eXNkuwUbcABz5U93BCGp5eTX+0wLgQG2Hb3yyFFZSKXMAGChzs4q+qiekw
tMecXDZY2PKKebjGiQx6mpqbjKD/44SvQ6zYDhclynPM93pi9OI20SQet+J9Mm89
BQZYmCTswGurap7WNMj9n+0eRaf4dGfNl7kSFQ5LUxdvE96heuBaTi0lsmsCgKL5
CQP75udSO1J9L65XW7BCmyGasrK6r4K9rGQx409Qzjz+eycet2b/NkJbCvXbn5Z4
LQSgTl72lNMlLgHyNeJiCAMqWVCgbn4jIR7MMNY+ekYjfsqmxxtJo07Lu45qi7sy
rKQKWjT7PNccZHHtxs7eFoDRmCUTGtfecA1LWffS/o0QVOwsf5SPz8GJJttCGr7p
d/A10+h59aka0bw3c/wu1skCoQx+w4IMMKkZrN7t26cHX6tBAm95d7c+uycRL0N4
I0tY1BhE+OIeDqD9ar5/u0MTKXHm5HtsrPjVeTfti12MqrIs/lLQ6DYhEE+6Rbmx
SHox1N/jGCN7fFMWXt+5nuZ1p5l6ToZPiiDqJEBBWaMpgdj3xSCt/mHc2B/otRPC
EhHGEnCPKL5yUgfot5D5V5A+jcRuWefLdtjhUCoozhG9LXZDWEQvTtLzIhaWedgQ
l/OKZLuvjWp1R+B6F5fnuaRK/Agk1FBf6dz/CVnBjAbF7nyyMgcZwef1sehKcFM4
n217/TTU3nhFLcvbkki7zzV5JWByNOeZREUpEyoKGaKM7udOYL1OvmwzERVAI9JQ
7GHWOwWVAwtiwiUCTUKiY1hWKmvKhtv1Y8AE0BRaRWwPpwcoMa7FHBd3WwrvXecV
IVKKlk0MQ9zEDnPK5VJFiRdOgWqV9fGBAp9vp0BXA1EzD8i433qdlQwJhVBSDM1f
CXpB+FdZqhnjmB6UkF+RBj0wyfYsYVxw9SFIqAOQOgUWbySByWpDJNcC56Y410c7
Q3tumef+C1AmUE+CDF2HeLZ+zJQecCvPYQkImH/mJT0FijcZIQ5gcpWm5VeYKNbA
xLVUes8Hp10xpudMhDMdgLe/1wXMyn1RJVgC8N8HwvNjHE91tIBhM2LqG6zsij0Q
f/EPvekrf5Wwy6vunAP5T/rew9onk3ELIlBSDjBb4Le6CUdt/3mnJDOluyeKvpj6
VhVsfdcFPrCX7rfnjywOQ4Kvvc/I5xpBDQpOXMttjaOFYiw33V6J7NOFHcHuV5u6
YJnrC4mb4M2r5C7iQ/0wN20mcToJtkYh3z+WHDXNKcSs1BTo0CptwT0XLSQJQI0S
PgcJX88fX9QuqB4bRDhCvpBFXvMYw3miHr2jNb8PxRZk88R9yP+wiadXdbDLjD+E
s0wpPy0y4qYs28JITlIvrLGDe/SrNYa/sqNn81wL6LNNWtdVFXnLQMAnQXarwqpU
omwhzBzSb2hdkdjBtENhf3jd6E7U6j8gj9xSJxeA9xCUcvafaPB3MHrQ11dJHtDl
GgyANy4AbHicC3qJzhsEEabBE5J6nxW79LBYJ+86bZyGE04yHP229/We84ONSpKu
1b+GN+gkc4lDSAwKrqgtruIK50pirT94Lb0Qq6gwjk4J4dRPVBjdGGtbQxC1VK7l
xUQLsmTbwzfWzQb1lwWQam6fI4EqohZfCKaNOy7zQqq8TtbpZsXbGN5gO0FFblmV
q/o/2HGAKc+WJyeQpl6gv6tMRENu7QaFYIVmcp9yqscrLZFFPLJH9Fe1qnVwUVJl
JedTvLAtilxtCrhSoiguWZpvQOOoplPBy8o3xrUach5RHBkqQb580BFIe+RJbAIX
opStox25j1qJMpUQs3uQ9zpb15ibCS2ImlkPZP+OpTyjKxyvqpV7JBtxftpCpyR9
s00ZeltYjQllmWHss9M7e8n6ebt2X9nIQBbQNjCN88jIRswZ482Kqz8lc1+9L1jq
ecVwHy0RDSPghPX8YNMrzRuRri6J4IKaFW1pcIj1U0vc35O/iSrnTgddOpDxTw6u
4BibXkhodmYJlaobfpkux7CyHrGO3c97GVr0waOLEfMZ7vtat+hHLmBDlLTVrhz1
HkngaO42yJDtEsPlm4eDMUdKJmuR+uxrilVlgnhkeVrZA5SCR+TMWPbRFLuj0DMK
gfVb0qNa+y/SpQROGsVLb6hdB2MPSZZX9gHV1NOcPdJVONhX1RTFpr1iELhBizBT
EB2u6+9C/IGDG2G7YMEVaRRzGTWr0AMftp+M8SIlvp1AusXp1F0yLR1S+3186ddH
qcbJLju6sQYDWVb6wqA5YMGIoVgYWh33flhZVGyFs2A6sOU31q8VqW5uZFp9P1Ku
82RtsEJRC05ZHkLSa1B34hPtp1Qco95o69x0KIrHChTgLTgQXi5z9XZ1J8BVMXUo
J5gjmAgt/U8uDmyqtOt5eewqGRBBOn5+/AOgA9vPNAI0Y+SUrmI547MJcstpxMCp
1NVJx9aiUPAcMcfjYwKT/TflMJBXAMapY+Tn91FbfS9hmELuSLQTYnKNM941E8h0
4bn3LySTbLFTTctEDRcxa9nJXcBARnXFN26kPy3M1iiagn6oR9fd9sAqnNXNyyRe
4b8jwE56TFrUhxEflPlxQ1BymepuW59bBMBAiGZry56djcwKSeGx1ZUJdf3lVb7b
3AU75ogMb8akxChdgAEFw7PcwdEwEIOpd6nhqQ9DwmH85Qu/J5oIXnlFWclX9ORu
OWbByPp26TQt8nuuBAHVrUwUNhZGuBTVtsUFZ8nN98dpjm7wEi5zcULy5NQJpAH7
9uJvKbKEeInx8R2CKUC1ZWbY3omH+ukcT7U4o2eRMK2fEHJgQUa22Qd41a/y6tAH
xMWfXNkmrYnm54+LAR87ony7pq+Gz/cy3fyasL1mpWA8RLy9NUxiOzjNutcsY3IP
hMbpxUSdffa0OuHRHPnKovtQ4PtkuUSPsPjq102t/UzZae+kp3DmJ75MBjVHNVzB
TGBd43SOjpj57sjaeJgizMRLu5WgQtknU2eEwvt0o9cydMIp/q91NSnvsAFA/4Q3
t5rtpzeP2sVShehWJI24bcFN9G2cjSGP9SB+4y143Ooqo8yQqkigghbOckVJDc77
KBfzsCo85Xl3fv5Q1R/dQyyUPhvszONe0TPMwNoR5IfZI23eRxZCFPQnP+LNsltX
Vqxy2xAc1wIm6owfc0206EkkjwgzTI3AC6yHVQSTwLBHmKKetuWnhypVkPVCeiZg
G4zLk7QKXYKnu1a10JABt0S6Vo1wnkGYjAj132vvx8fXD4vosIbHFUX9CRK1bcp6
lQCT6ZwnAkBf9pZ0lhMnMJySdXVBLkX9/wwHscfYy+tkJuPEJcHsBh4jOuyw7Zw2
pOCpTS9qyAKetNxrVKikotprTgA7FIDJp9kJhKzW25Z35R0JaAau0eVlkyg0tkHE
Z9sOdsWtc7UI/hw/ejSU95rGnHZ40E42+pfzWiehaRTKVZjvY7czugfYRf1h7gtD
8+KAtA92MdUtG/L6h7DFLelPqJ+OF4/K7Sk2gwf0ijZ8wBf2De+MbpYFCV9u6t3Y
qlJjkAkne1dwXeKfFLRK8PkoAI7xmHBYcgPYHj9UJFeLj+u45bQQ0hAKSlZS8XNf
9v4Pl5NP5hp3SzXdqQsxA/KIHbJ+IzRGo757j7pYjyyBdoSp4H7o/t/KFILgtN6O
Eh6HZsTdR8RlQZ2hRfYkH5rot6YXK4QtuIRX7yT4HOhNW+EcTmxPp0B+CdUfXuQ4
+vlHc13zAq9ZwRk1TU+3U/CFf4MEEpOWcbrJO/c1mpCcQVNPfJAY+IQ1Q0974Awx
GCDNnmdF2d9M9W908GNpokGfhAV3qq2XDAHARJnFIuD2o6uwt9Nlaescfv3fA6Ge
hnJ7BjV4tZQqmC3EoUy4iaOowWGnYrpYm05hSdkKXdV7h/SFpU9TKnILhymv5jxF
pW5nJv0VkLxz0lWoHBW/i4y0XGTTXXwRJh2r7TSdlHm5dfxY0uEkESixrpP7I2t/
e8LfSGEwy1cyKI1WuHqVliyvM4OeEhJQrdyjdt0Q0hgv+AZY33W7oyMD3/zGcMQI
RMbltn4e9WofhiwjV3F29lzIu06d29LOwwANDbRefWvNhIemchjFJEZHSg+biHsq
Y3kQZy0U6ZYYzE1CXXC9cw7ohhhtHj6G7P45zKEYwggk55YOYxl19ZBgvNhGpYEO
Ub+SUAWWNIh+ozhhYxgdS5cRNiPBrhU7QXOfQ7vS4yiD96FMmh/S+6usRt4VQ1je
1eUH87bmJIr28Wy+Oy5nQKdDFxTASP64K3h9N7ueSOh7QbHrbAE7tl7CVx8NUxd+
t07bpgxfbhXZTzhJYifTFZV5CrnQeKLvfS5DUO2J3gZE1w1BaucqG+tNkkooX+5J
yEctKMTzXn7npT3q3JNdq0NhFBMfYybrIEAI+0ZAs5AGVd27uD9qoJhS4V9T56b4
d72y0/qHtqzY4+4d6CpgPnJwenEmDhUXrvahhrb6azknLLnwavUVmQ8Cm+UDS5d4
QN3W7/Cyc+nkQA8FqTjWab1fUv59hGyC+3s7J90vjruYjqYJ7Dj4lGG4WUA2jReZ
2jN8VWXA6p2/PwKvw1ome+Af4r3i97Ydq1XiV9hfH1le0ZM6xA0o+ngvzAgHcz0a
HhJXaXQKrOowgB+urjnO5UbOC1zeiZDHzi7WnwUgHnpNC2+A0ge397A1DjsRzcqZ
/lIFm8exlJ6+XU76rKpXwOgihr0HL0mkVzE9CbfZtHpUkLKhABaUdQczOkKkyEUX
CA9iODnE3hHSVNJr8jvPvzk3LPt2hmPmNHBozoeOXQgEim57kbmX/ncX/WfUc3VB
Ek6t2/s4p6n7HJ0oVYksVhqscruIKbkMQNMhw6lQSJULnApVXByomRkQ46YhmSYA
dZtQ6K2VHptCh3V+Yl2ujvN/uRjsDlUx5MbDtM03XHguOQg3OifYmN6ISj9y8PnL
kvAobdNdF1+D4SiowHcwaNqysosaNxOImgni7DuYnBLVYmRYxIzHa7nkz4R9Zxur
s18fJwvgxvpTCjiJ781H6XzZ7rtb98soRprHeW/Y+gmyrRvtyv6U2DFWe/CezBnP
pYeqS54MdWlFBHUTt2zI9Z3z3WKSwuRUf/41rqSKO0U3+Dwh52q1NF3PuhtcxoDf
plhmO/lOIYcv/gOt0snrlaHtwdoqQuWkBuIvleUanF/zdjAejv1UKrChspIQ6V6l
JYoJYmEvy4NcvCRdiLC+nYH8v42KLestY4t/p8+5QSW0iqF4qVldM+nJB2TVio+C
nf5NEs+FI5SWCJhdHwTBWLamn6GHxbYcQnlE/aRBMSxL98eT/2P5SNBRQ3ap6bEG
eiBPhfoxSi84kNeppHUIs4MkrqDCbhGUZCI61uEAf/XySWhNp5j9mVig/un+B/eO
lihqS5z4XcM0lcf4dmfigChP8PUMy3XSrBg8WLQP3p3v+xnys4GqIYCIWyvhKKYp
Ls3zS0A74jDkKf4MYtVxOd4v1QzNQJmL0L2FOdD/IEq8kC9MTVXynSZKFais7acK
fxfDcLbKX0U6cegpcqZoblxQ843xo7QRas1mCMZkzkC4l7vwvRcX5l9kAVDFXq1L
xBi1W73X5WCXV0Pg+0YwMfkZuBpgJ45rnvLXp96HJAWJV/QEy1ZYg/v2jyYOxCDh
k5GYHLGHdiKw5lu+ufOpmM96GEJonj8gv3PVz9yL1wSWKerEm/CdscWyki8F/IBI
xwzbBxV3N4HEfG38DKV9M5tN3lGyLuqKde/RgmJISyyM5wx4SbsoZa/9/mg8dlzo
bGV+h1MO4rAZOB8HjwWP1dB/AQS0rofJjjv+6Ql6OarNXAmp3UdVlIQ4iaNmClMI
zXfu12eDP1lF111ExXLMLlBV6x1Uwqe+Mp38ZpjWHwhXVaef2xXz2YfaWRdfMGDF
+jiueNQhcOhsso8p1C6y3clhcwbHhGcrD4qcwePbGTEvzg05b55YbI3paJB6jEtR
t8rrfhBkCDR8d6jH4EvDLlLpc9UWsa8ad8AzkjozErlBOsCeMitlGfucIAmesRyk
RhS1A9eh8AoY47nB5iiooE2VWe8iRtTzra7aspXnIPrNlkuSTLplXBZNzctsZj47
xFJG/1qYxInxjxxFBpLKCQMxLiO7xTaFEiAHk1CTZKgwRVWVkacYX28gXKx3yBvx
bowA7mCNiB5AUDDLRwsBsZqnD5E9nya8XeMm340csn5t/jx5H99420meUyfZQmhE
G3QBpn5UQE78v0Lkp0BO2ZFPB5jbcdqksSqJtPWpFsqcQBs3KFl8KLoKgJrhbKXy
+JVCe9sgHunDh5maUEjI2rrtd8SZh2HJWPOP3mOqG27LYj5kduMuECnq8I5hXfsx
Mo0KwxuLDBAllt8P3g27Q+PTgUnOzkkAzJMebspmsTbuZudYLmzV31xg+kn37/Zt
Jl9H8qATxMgRFcHO6Cdwg5To3GKngJV1/Ach2u5Ioi3eOg/+nWwJxPIxtUyhVOMg
o/05cLs9TijrMDf69fCX6kwplsZ1p9u5Tw017csxmKI2gfattFhXMUSlVwPEnCYn
CEabaFrXOnEmpgJx4XWpy3srUPbiAPnTlcbxzONHI4HdcaDo62u+4x8thrd+TEuR
3nZ6HJsTQpGHsfxbqNBfgF3uFaMkz9dqzMl6MJb+omySduBEPb9zdAu52wdg1vyQ
xdZLgyMVUh0Dl+PpNcWjb47fcJ1peYt88xz34XvkyA1BS5hinS4hsXcdkY4mK/Rb
amYjcUTk3+IExY1d35ypLi6ivSqmigGjiQeFsHgLjJ3P4bl+GRO+MZb7/Gh63KjH
nhrCHH/UxN1yVc0uKLx4FVBkk/kw1paA+uVB1+RBmnkwFSwYgT2UbQ+3/29rFqZs
KhFbtdatBS6RZ2wpf1n6fcuN99buDBYOLOBhkdvZQp9bISuBntFpuIoGJCKQe+MM
/4EzFqw0Q5Uver0hAxrfh1ZmDRKoYCaLwnQLzzYuBN53tw/lb0ImB9FRR7U4e96g
PjQBcyY62/Y8/eRAxcuh4ecvHvTy1iFBTw7MKBwSjHJh8iaJ2Zk5FWZ4GCK7JZpp
pHiqzUTnQbS2FlL2dexFvylpRBGOs9wGjRxgCoGQSaG2Csnpew3iWVleaZQQVpTE
nUVP+s2CLAbZPSAQ4guQ/8cQuOJPzaa2q/muCtxvd3M6W9J/xw5UAsU8JTY25dld
HwLsYb0A14X4LMqpcgNLX033g6nn8NdmX+tbhbLMRhE5lhgipOqsKQevZFEvP0ch
FbOYCmJpu4g92734SxX4fP48AzfCjONo/l+d4anKAngtivpiptjdtNMtNxXoWzYI
h+w9mLTFAhlDPcbl+P2HTQAXPqo6A9oYyAWi99opEc5CQJCFKlFQHbxhS/sRMcVJ
TzpDhPUVUeUb/STXS13LwzysADOHajy4CXk1I0zrfBriKgmfkekXjBE9sB1CVOZw
5gRIgBlDaSH+JgNUBeAzovhw+X/2IcBZblYkS6iTxcz3XJby+LdJuS/KuDaHX861
mOiRi5RyyQwhQrT5UxFvER9y9TIaE97inXoIOO2Hf9MJTEe/QgYNjV9Q9NOLTK2Z
oSlKS55ul+KnD8ejIuKNL1+3Nor4aZ1krFi2KHG8yhGxjiZ88xx23fMfUZPryPe1
WQ0qnJFF0RA9PWB89yuojeiDSQIhGwIVzh18RbQnY8DSfpC2GtpeYDvQhGfRbJGJ
+cv+wZ7UFM/ejMmjupXa9QvZPslVEtAuRCIMTTgwWkCieA/JDRLee3Y38y2Dig2B
4g2k/1f++s0vgZpMpFtEG3rqZYCN9e2IFai21LWN+s8vH5+FfPpyMqPF26ZNDng0
ljZljylDUzJdXbGWdYNMIxScGFQ0vp9Kl5L5uHDs4exSGyDF/QzpFNh6i6rlwXZ6
UYedhulYhDCUYXPPzD/RvNfb6cKvapnPDIsf8U0UH25AqEVt9ymFQPKlll0BMut2
k3N/fY47qBrgbRsDLQ0zp/hZnmUDIqm59unqbnRoQZAkJX4OwR79YyiYpCb4+fbK
3CQUH+HBuAvIdYqac7vyQloTQ0r7PK5SveVcy3+aPUCmXXQsGuE6jyqUz1A89CsE
03QvhYzE2GqAzJvayjiGkyOPBOskxD9xOQh36zgK7SoXsA5IVyuGb0v4vDeSRRLq
IykhO0aXaVnfcDaM+QUq6kgBY9HL87xEz4UHmc9qICYdItlms5K6q9YLUCN5OKiK
y7x8/n6QA8ZacgPAmApmEUuqQGxPXJ76oBlUSehL/3CeLZHVDc1/1DC9yidb50oW
7ZB4W5I22GCMXvUcQ1s3mRwk1NHPlQihdSc3Rwm342l1E7FFrVXnT8cpRc1AI8sQ
2i5gijF1pN2b6Bkt6+DCt1QA7lWtwjjyV30MOUveDvzOx4pz6MhHF6wdZJDKiQKa
u2JFqJLFVlbsTHetiKfKXdsdciEVz2PNKXyVqwvbkPA6Q+fdX1+7IJqYI3DUz9oH
8ENqhaZdarvvh2Q/MDpRSx0sJGxXvYZi9x2ThJSrasdAQ/+bdEnRY35m2RY5F4tM
iHK0niP+7m+JqYGT0Kyk3OOTDNR1NwY/YC+/isQMMjXrih0aTGDVWPoit0D9JxOf
1ffowOAe1xITyyNz+Or2Um9NcvrsyD6bNR3+G94UR/dl47/h+OTp9JBXenhOgMzL
IOaT8w4s603+87T8EHn5PawCuUVDMi15E+ZohBzY8aO6mNgCbrpbwO3P2/Tyeq7z
UEBgeDzmPUETqoxSHdMAFSmXwlgYq2AAfcAClc9ZU9tdaaC0AB4FvffCGf+7kUkk
ER8EBW9LLfSvt+bdBoX7eSZhqKOGJCj3AJMFZsfWDC/9eMv0JR3Mwo8i4taBecNx
Kc61UHfVUoQT2mAI3nAYHHuNo2gHm9bagyroEc21SxfpgnutR+nNZLHC9ZJyVJhG
+73cMK0UnpZaBovrtBJKwavwgSoWT2WaBYDl8bduRwmwmBJnp2yEgeRX9oXIA6nN
SM7SrHiZbaS+45BtcsAT0IHbg+1Ut2YdEnmzF96IbjoZXGARraCUVULN/nGRXubN
jexaW1rVUqdSkR99Ln6XCeimAey2v02FyjfwPPiKcF7F0pO3Nd0cJBvzNSQaV/u6
IzWHw/XpR1dnfAW3aRgIWtBYF00GFwQrok4Z7Xzi/PAOs0odTELWLhc50I4+I7fn
bdb53OO68ZBve9z/snyHyp4+0h91YoU3ItbkY+kUn1TxqzzL6BkdpKt9vhbw0EXh
C8s8CRCCx2Q0o1BXwKTroz9p9XuL0cDUFJ1OXlSlyslDrs+hWiiIue+lUmLBD9yQ
DEHZXuBv2ScWEHtM7IBGKtfwRcJOzz7P/ydw0ANoBJ1hFdyClLZGNjgKyaJEUac3
tG9NSyw3fHQ9rlW1uU3vASsPJPQJ27ZqlCBgYSsaUk0gGUuvKTpmZ3Jm0xWokXJm
NYeeaTApIVnUhK+LW/7vi+BvUSabRoAKPWboSdVdKHil9mIaOAlGQ91qQQ6cU4bf
hk/jc/+erlAqo1HHCnpQWu4BFL7nKOyIQwr2sdlCPTZJET/AHkOJhax2wRGPw/4+
5nFvyoI7KxvbufKq8CpNTF/DQVCPLY8LJCcQXoagqscv6sTL8+v4/NqnbVvc2X2/
5g23DsU4KvybJlHsRI224HzrSUNeFHsCiyzKmXgcYYx2zt4wjHrTj329zfyZ8VJH
cAE0WSRfxrT0HMPG5VdHBnepbl0HMHm5tLOT2BkCu1pwbR7T05mlFF2dfxIq3t+r
E+zDVTXDLwPGkN+oNdP3ELMkflXvV/mE1YC4wbhuHRGbojxRtsTckOe6ABortK7b
MhAF1V0y+b7CpwM1OZLKVyiT9iZamZP7KbBNrTeQCX97P5quGm1YqLTpu2KQqonD
H6vSWkBrSUraYDVZbwFT1KmN8RwBCS6JMEz1uivebkSVFhswZdRA2I+S5MTNVUOx
m/TzV+FtAtCWIABp+M5Qdu/kge7ziZf+pYP+QheQQRa+LUVzKDh0PB3zbo9nF/ip
6gL1fJp6x6wdWH7gU28/PFgd2aLTBTEJKJH8EQgbH1Ojd6SFwHRiy2hllOKu5ZCN
PYMDr57g+3ANIpCO2lRbJXWutVJ7fMDn9erDB0k36ROftWQHdpSzaUbcWmTMLJjU
RjUW+hbb5FrVPwLSKC4CDje6Yp6lafpX9Pc8ApfgrSg/mJZGWhUoL9TEMCln2jNC
UrtlKFuonhRRNSXNSPA5X8ac1ZTxOFmDJY+y13jZocjS6r0N27BLkt/2oK7aCnzW
UDBUP1mlM6Z4ocusVRcFUjtXRBnjV8NSoBZ/8g+ODm15UnuhiExj7/qPQCGNtKsh
Qrr2NbZHtIKQrEUsh9heizWJar/lrRqDl5lEJsilocyA7nHTW99SOKE0oddo7nGk
+dfVAclTI2ykcn11ayEhzZoJWNOnpFmnTnRevZSRRFRgUNyvBOWDPzjvRg4TfJrA
hFvGsOH86EW9nUYc73jorLC88xm/Jk44RiijWzABrg+xp+8JOIEmAdIpAAG2a4As
793/NwzFKUGPH/+Tg7YZ4XSk+ubxofxA7PUAzz/FQc/EhPFtnNdwUXj+CsIYvd5W
W1smSXOIS3dEpxggVOT9H7UtBs7qmGeL4wn1NH26+lTP0dYoh7GODhELDOuystDC
FMQiUZnpPhT/O3BWNm0SiD7vvKnMHCt60D80eSzNaz7t9h/MVumq2WmPC4n4WQYU
j8hFX2+J9mDz8r6ZsjkqS0mvcXtRVT0JREhoxUkIJr0f7THT+DOnkRWdPcYK1aDN
LuIC+Iw7BVMXFxOesphpEyoyifRVgPaL8O/XR4u24b6Y5oQoUB5eiWjABSEBb+23
uc3mt4A2yhXwHTy3lvwlH1RZx98gn5tf6KUQXvgxK2RRAYzpMGfVztsc0SJZAFoq
K+gEUTgzxJKjzKsn0BN6Tt2fbshdVHyOF2dOelQvJ3sf2NYt1UVaVLC9pnL9YPU3
/C/DdbTDuwcye05BIk4N26CDntz173S+iCrEDvCaTXGUPq0G+ggSMLKsjuStwTNJ
trJ3Et1eSJn15IhyWD+PZ52F24bRnXysIU/alnz4ZTDNEqlKU4uwdQjWe2ijw9DL
MTUEUuMbXNCFVJZlclwhuWOcd0oNBNAe+Yr4eRRYDzAaxGwBhUagl8hBXOzxmyY+
NNR6p7ajqIyT6UKuN3cO8y4ns65WGXw3KwRSjrBwFVmUpatlRs/C/dwwOjpATUK1
JtucXbf56UOMt4JxuQOALAinEhhW93g6fPcngcZbfdG1tPCc4ymww4t0q37tkJm9
sH2Q8j1Wspmcf1QewaLhcTFxEnseC4WOTb8yhIO1R6n+DWE1ODZN0nJy0wtWN4mZ
Mbh2+3N2N1QN3jV//QOKw7ffV5wvl3LkKuHuxguOICj4WK0u7sxJI0Pf+yy3B1WZ
WVzulGkRaO17fdo+0zxHEw3AWnUzA+7Rshh7JzSDHz8v9X/s5GP/zWfQKAcR8u22
Am6BM6z2/kML8rYTNcmM8sVvlN0Kw1xRMj8V4r6fZn7TwSgSB8WT/HGrcYAC+73d
OEwdjanX1dfdDosqWVDqs3eh5hw1zuVdUjF6+IvOwtGSRBkya1SELzB03ik1epMB
A9vvUQK7exMJkwdjv4ZUa6qAf1CumMFCrcHcCu5Ke0QIW40J4guC9Que3Qw9X5Zl
cGjc+B4LnrBFl3pI+Ws87eTj+/q3X9OCzJSXZAa2VVEkhLn8yaOFEcEas+glAnm6
zvq+cXFK2E6PXMkUmmEO4vSzvYe+qk00whI7l+n15n+cU15aPSB4HEy+min0RTeI
FZd98WleYxurBm/G01zI5hnFXkhLGtUKUOAgNSUH9a3keB9F/vjeb54tK6wGvWRt
BaC4c14ewkW0hesmavhixSst+vTT6UdJcyCGhRdTC4wNyh0VPL+FcC81WzJnzRP5
ze+61IQ3N7QhKO6X2QfMAWPE01DKf19TsRXxEJnAzKuqCILWstfoqcP3MGOUNyoD
7ixEMTxscnqis6rfc8Kla3Zu2Sqhaergmm3Z8aWqO0VGXFevX5k4rCncP47qN7eD
jSGrAMiC74Dxme7bzFunXi9Bs3UAx1crvv2LFN8qLyslEzESR1YDTcTF2FKOaO0j
KQvC/SCMOa9BbJAJNkohQl//Q1ZKSQIaRQe5QFRRGyH9xFje/ekWLTzS+HotsozP
+bQM8M/6ChTFe6jmvCiC1h/IYhst74cYvCzj8yNYWa/GYvQBrNEgnTaQGgJ1djWL
PepSzp1szmzU9qhJT0PVFadA1t4XonzrXI61UA4SgpuhueAzm9byRI3b5Rx1SKkg
Any+jind7ILTKndFIswZG1X165EFAJRoysZL2pf/p6uAv9FlP56dlHuMdFUkQ6wi
DGK1otal6sa/+5zIRk2k+bZr1sBUV8Yz4vJ7lq2MZxhbh1KexJKlChBJHYwRnAbj
RJ+bANaor4Ga0M7UmugUAQxNp/OhvOMerudWbOBJwzyE+VrkgnQ5Cyc3BG2ONnir
oGjTqQ6HT+ElN2raoAU0ZzKexXr+N7hTkKVg5W+/JD1i4o88QsJZOmOjuUNhVnQB
8G/iVuum27Q2eyU8kKIPgmdnOe7Mbfd+PNy5Z4UQzL3lOmo+FXD2E5DSWZw2LvQp
1UZUlQ+4ljs9quJTqztvg83f717ibglWcG//BpBjup1uQglgqiQwJoYUDVHGHYvA
zEPXGJRTtpP5nV062GTH730LGpKZvATsuh3kLt8cqwhJ3D4oHS54BbyQCkiLSFVB
wU7BUNvCuCDjddVC1TMRtrLhz8qXJ4mnH/FFwagxWFF3Ae6/xh4qA2Zg684a9VrX
XhfEl01x8iVH8I65aUlBYN+xwNOp0yDM1aLLUe470Lvmnx9Gavs7CfKQLTqm8T3K
3pfScvis7z6hEqoNuIA3a+XO10olp5GVjJHXnDmjDwQBB85Omi5+kWT7zUEwyCOv
7KAgs+INvh5uRF1lULULMcTeO0lAj12eedyLkJfFFJtpsLFu+4fc5I1iIJYrUqi4
AnrdIx6S/AxsZ5LdoMHYkrOlH9/rC7E/8XkT116MJfW2qA5cBQCjCdNFYPPRlz+v
Fa3DnvWuJDh6IpNx96QwP/o789ZQHWRmC8KdylyIME61DFRjHdtU+hUB1fHperxb
yjIX8qY2fcple6Lskcg8JeoAg+0dNepBcqFC2/HNX/wo+ecgvq0FO1YbDTS2uOwf
zFoso2OC3CQsACGud8rG37ezyYuUwHmZVsnNKbiJbueRsdTsUdJF+ldBGMd7ImfF
LlXfZjWy+guKKs5X5OhboTG1E3mt553yc6Ua1evt/OaICrlDTDl3LWF2+qzrSUgH
JGVx84XLD4HXJincQJXON3C5fZoSQ9MAf0GShuoAkntJphh43kLPAhGoK19bp/T+
SBqgvVdwjyy4OmPu6w72+J2VmIZhTvyVxEXyA3djxZwv9K7pYQ22P3ouCCXvX5C5
bjg4x+1uRHS53oW9XyqAJKSf4VydgHOch7Vv01L4up/2SvNTO2TXm+xhq1owTMeM
lSKTo6LlmmBnlhk25TazI40ZtbMnZdDl37M921JDW4TipWxyf1dgfoCfH0/87zZQ
rsjUdGeTM8OtM125WSL3WiTikDzCGCKghGkX/J3r4oHx9vq47zhBuU/8XKn/bOu1
aPK9fyIP2Gv3opvqMMV0nKMMfSmVYaLNYzpizmNMEX7zpPzM50Gc4AGDKon5nsoQ
m/M6J8tgjWLgMBkSSuy9vVEFRmfF3fRYOek4MK9EV7pROcj0gPFS2OBHntZQTOm0
lZ8TtOTtqE8nmiAX7VTa5ebLxJ6lztGtK+tOqK8/LKhG0A7jXK2Ipz1MvO2EK5OI
rv5jYhJkWsacAB52vWwmYMHm2FLmamXlrTvNs+GMwVk+CByLqIUUYLENUYo63lDo
wKEMb59M3XJfom3XpT/AouryOW6ErwRT0fW3f9Hle5yfDhNatWPR3fLrXbyIyC+Y
YffbdWkl3INOCZX8r+fENDm3e72Kex7xJL+aAtJNFaTziHYdYRh+OFQIWlkzro29
qHfdCwDDcO2WcRfHae4CXB04IatZPgbgZchsGP0IIoNWERSxnVc0gJ5kK85gXg1G
CSioJ9MHPOREDAFWCURgkC+pSAyMtKUoj5i+q3yL36KUhvdyEj5azZyZrP7n3UZ0
JvQq+QcNKKtPazWM4i/SDCHUy6E2tKtMZ5IBMstPoldePgBVIqr0fi03oREiEqX3
EKqckvRUhhPsHOxih605fg8h8NUNl0u0qtSbiUGrMoYtjEgbeOqvNm52IXGzk5Oa
DYelbusTOUULN5eM0V+PGt60iKW0qwjPQ/tdhqdVC5FLq8ydhog6azvp2C3OR2BC
MaPRJO4cfXk7wTRWzZ/iq5vws7p+YXe4LkyK/IeeOUw/tqwp/iT06ktF1V1VA93A
GLZsIoHbc/bC6xpqwyKyzBccYAynLPABTukPCla5rI8lz6mtj2j0Cv78kiP3+cbc
Emlxbb7OQqQKDA3eW7GZzcgwgJy4r4FXGN3MnwTi2xYh3Ssp/FRLiLFL9JkwsIJk
8UKdX1JZ/MW86+gQfagHbaW0YUBY1xkR+QOZB+Wrc1pYu4A58ZwqEdALUZxeiyTh
Ts6gaE8KGOfMjfPL6l9owjE+ZrJYiSBd5a5rrb3swrjo8z0+YpPqsgoAiBzKLDrY
dLG53D3F5pb4JPJ+Jlt5bpc9mbgAtOphMrDVYlMhoZQahdu4eICdRRKHt6v5VG8x
KK6dsVdvmMrMUvbgzVxl2CWrKZwtUcv03BKU3f7C3q3Beaju1OiTTcfTidsS/IKf
m/KkMB+PN7JQB6xcbjx6CLgt/qWuIFrP1aCvIq6fNfZmgnsmZXRr3PELSxHkoGGR
FOHAqWFL8ulNXuM5jmBYIonXZf1Cp7He1XB4D3aWTBWtyhBMx8Z389aAoR9d7CB7
QQPCgWelOj9Uglz8rPMjmOVzk4VJoxhXlZjw7BLQMlFKSK5tbr83DbUG4SXeDrLk
YukuWUsH2Ssw0cZqKkFeGs3rUu26SkhdY0WfEaFbfyREuZLHtG5mfjmZNgL7u+VO
uDeBirFj1GwZOpuDJ03Wt3Mx+w3DLYF4GRWVoj1NrxbKnp9Hmw6mng5HiW19Hw77
6EP4b9dXzSI53T4shlOsXOFD+LHQkOhm/dsyueLgQQODIo+lI+ohkb98Ky6b4j8k
Jq1f+LPfxv/WaYfXx0Kgbio5PxQ4gFx+cXxYZNzwYrleBRgk/73Ov8cu6R6NL8N5
JlUKffjfQB5Py0PCgVI+I+Y4Pr+nV+hFIfV0eNXABUdRPS69IzIFokqhJQAcraLm
8sHbbFIC1Ywb6wG3CUPmKc3oqePbK4+gefqcdDGpKFwTXoXQ8c2i7TvFfVZcz1jO
/ubICf5+n2jLNEb+H4xi3o3fIDmtuiJ/fpP9xPNWydZ2QhbhZMtIl7ZfmsNiZ8mX
WaufUAlwpG7+tOz7vltj1legj1v0Fjcom8wwKgwlF1ozyUB2SGLCpskWPh+Gm6kR
cMo9mF5g21UKp2kpWDxkosZDN+2p63eq86Idtb9+/9KMHHPi+rxN/llsQrlgMftm
VhhqDIc/SP2auo/1zo0duoIBYYdrnHJf+JbLDRklJDhssQUkUARk19BMdaBglRxj
xPo9gbq8Usr6ZcLqLh7qQvppU2nhxxrqILo3NflWd1wq+wAw/9RmWeIpGh7cG4ch
0prOQ1IaFgUKd0DXTsVTjE4FMhcH+bxXNEAC/BW9TGYDfJPIQ5MZ/uCHSwL6MBN9
+XoiptVz2NKQyvSj2Nyr6pN1cCBmrKSsA27T5A101bbZOfeNwXxUhfvYIW8+ftmh
RL/J15P4nEvI5F2xDWMe6nSRYjzT0O/7WU5zQuElrTuUikvyIk+81OuYeHuGHdKK
4Owmz2MAYocHSYQTxRYVMSLZQnP+e4en9ALQ8lVNU1aTzpDjI0HKyiIRjLfPLq2R
PkD7XswZV4JuGAjJpJte6tP6ETHC2kfPUgzylhw3Vz9eK8y1oEPefhnvfvj/BQvP
ExH3buNBlWGhOAQ+/xVwwi/QdGax2O8B7h83bkd7ZICm5O4p060kVvexc7/RpaFA
ySJbLbP/zyHNKp73MqmeVeoETB20u7UargZJt4vVfhwhQdk0G1/eUCLT/eUqZ6Ji
QcUcwrKpiyxm9xFznbUyZqH8dQQEURptJ+A5/cNiQtPijU9vOzACIhLp2E1NnyUN
5L9rEk3Idheoty4enyGWWomJ/JVmDk4C2fY1BCbSv1by5NNBBme1JXBJelfgymDz
LUD7dxj10BHVqzQ1U8TQYhc2W4px+X1eymlxgqSBkanKCen0hw99h6/Fgo6k0Jr8
BBN0CrouqRjxuOHL7ORMEKxnqDbmJS7EWU17aL3did+3iUcN58jXPkTeP/dtqkC7
iZf+mIU94Iikgj65OcPYGX6irYX0hLm0S84YY5OVT27kVWDCUvKXSNGW825dpbfj
Ll6pFjWGbYVriKngogT/LdrlM8EVjqUmNAouESu1fKLjtuBNUuV6J42u0k3B73qk
dVYfHupwCowt1RUmwhywhB8pNF3fvFgDo3cHT44PXgd7LvyJeUVrugfqShK8evCy
H3doH70EvIH8xv3CLJfAFYNeQIeIAiphzzngTzMcivUkDPpRv6yFFG+HpTqNKN6+
k7PzkKFnm61gXUcWhWcFoiVuPltZP5wbEBk7d2z+wQPSqawmuuEWPPZdID9qCAAu
O+cSceMwVLo+k9N5H4zGbd63zqwl9kDeWX/+xA7hAsC5iqWHI2wkHlFyVW+4qzEh
2Vjs/NwF8b3kM9wihsVSwykLFh0i9yewMFvkDy0xQGN9DNNpQXcdeTpGmR7l82Xc
aEJOvex0IEHryNXlcO7gXmbABNDhpZglY30AZPPQY48JPGuMAIeStByuu9VgGuD5
k9j3dYa+VoNEWygRu9Nf278kVh3uhpfnI0UqohCxNp2QXAQbbF7dUqXHhn08opdz
0rqK5/SsH7nVbTN7KeFeXirpHdLJMdBZj5ZENeE1gxTC4/54gv1Tzk7PsKWsEMAc
0wogyPQa6Qn/lfRjrgPta6ePY+lH2pZmPOYWvB2AhEK9pyYJNk4VdMO8240kkwxZ
GnWhd+2wwxPo+jrDnDaotZCnHPLWNscJc4v9wAJL5TfEpf15emjiQ22x5lw+L/X6
VE7WDMOo6XP3izctYFazMqvoC+Olsc1IgLqrlts8os4V/qZBbPeC38ZvpJxQIQRd
zWPheQ3pNeN8i+o4TKhIm8ANmQ9127uvfj9hA0FUCvmVeA/lNBqSxJUzLZA5YT3R
jh4LGENPPrhnZUVXKm+pAaiBAJyW62mIZjMpuDLwPJmTwYTjAjHOu879FdOZjZ11
ZatZKBw1oz/XttEqnpLCn1b8LzBSeIta47lRuDAzEIEwbuew8B/zDKW5LFf7hY3+
raLtExbRoTGvKLAFglYZKBhAAwJgbO6rAGjXy3eTKF3cHJLNOz7LLL8U62QPGCoO
ioZnTp4cB2QF+ytxK9OopVoMF929nZBbjBuNZbKEbXzgKf19HEEDz+N6qYafopLF
htjwiw04hQpfjBTmgDZS6lP6W/FuRPgMI7wQYd3kA0irhj7KizAuYPZg1rfcfAUk
GGqs3hedSrsxpsGe9Zg0AzjCg0nxuRi0A0OIki9Wyzp25V+EfYuxPCBSo/lEeWQZ
aj0HnJU4dgNDIrUrJFhK71v2hpmXAS7bD9Kmldr3+jZ0PCn9EQu+ZyzJ8wVEAbsz
cwEFAgSoJx8JL8FsEfIURMXYNN/k0dpfBTfoMyGHBKHpJnNbYXQF75dTtteU40BX
FAtqKZ0xDyAZhlH9hF00RW9dr+oqAT7PScE7MjtQ5NcEDCiYe6g/WFaXbOcLiHLn
qmFn74AewgP4OI3Y6DcqgpHY9PgFBL6n51+TQF+ZK39cr3eepFAhNL77JQw7QQKX
befCInGAa8iLUDY4c01UECE2ChkfsRh2Xt5IYlCN+GwQs+kix1sU2BGvV8212ZZa
OgU5HyMsDKV4pFmU3AsRPyVbFY0g7SJCcYyyUt3tN7cwuRI22Tspe7I0wuLa0pdm
ObQ6osW9bmwRhGnWFYJ6YBhLne2WfGSeKYyfAnATAklpD7nw7vVHORrXh2xYNT0T
mH+XI03Jmgcbpi4Yq4wOCAXeRbgWffm95rtunPlphM0hGU8/bgSc9eV1RnI/Wb08
fkA4VnvnECg2H2xgK52AbsCdp/sHltCvAv5IIKTRjj+1LOKxV/tXaMjpCa0Wog9f
I4sKG7GXwK34nUMw16NicP2QR1Xra+ziCEDoamShDsImY1Y2dzJ8UQpoY02dkgYF
V9nTSWCKkNXDlds0Pm3/nljCN0xUb8/VLXRjLpmYK2iUs7EHU+yQWwTs/oJRKUMx
cjDnT5PJNm/ioWuCK9VnSURMN3ru09eIpMmvz+HggbDLmsndGmDjzsSrZ5v1LR5P
4m8sBm1o5ohRe+G0o6tFDKm7VSWYuuRL6qbuZRwiNFjVE4s1PO2XW2GVcE1g/gVS
CYlQLWXQ92e/EONieU/IqwV7oM1+VztxEUTQMJ4CngP2KRm9ZuTzO/ntE8uuFPat
gKeMZPUvl/5iYGM2OUKNbXdHTM/LE64QNA+zCpZ1RtZQZLQfQ0AcjilHAwQ4CmV6
baXYdNif/AzzMeliLn1WIqDP71rg42C86aZewmInhPcILkoCPCj+IDu9a/5ZH6KH
CnJ1eqQvr+t1z07cW/mfzCG9mcu4HrjsX9BZMa0IrBKE8np3XboTFTVjxQe6VzI7
1Pbv9MOI94L5xOJlYGdK5jFe748aGGHF8+T8W5v5NMBZogKhggGexbOwyn14lr23
2GV+MTQaS4IL+Nl4zhPS22bS/ljxMUQkR7wb2ftShaindTuMGmL3nzju9iA+WwGd
QAknkbaNdgCoDp1igw6JOFnPuEcdiWHcayd8SMOPjNPqnm2tEUVapa30Le5BJDD+
ePRe6E0jvM3clXS4gwf8bQXVDYmqz6vpLM1iX5ZFrc8kYrTFLs0yhyvzcUFeHVe/
PKlJFlN6lF2TYH9vC609hEH/SmOGgKrFjc4a/xm1+W1v1gsjplbATSP3xooMQLW2
BaMrOCk4zKfMxjFDRoTnUbu74PZRQ+YUbRtSxRVgvA1vSv9OppYuiulz2060+lye
0S28M4KNWA90h3M7MZTQYM6ws8ycGjJRIHz7VlouEOMUKWezW9/VsGp6XbT0Me/w
30gP80/bOO8WGaDoAcq8v1R4Fo8A9Amop2q0H06YIPQDCFyKJUCK12T5A/bQ2mkP
eDsNcUJWhhGeVmgDPxsbVaqZQ/WTPxRNMgfK2XWjmfyeRWKUIA6vKIgFTZ585M7C
nxhF+b/DhdMVd9tG0IIbvHqwblselPCVj+J2OOCfoe84mKP8M8XnCOXQjsbZGMWy
pKuS2DzNx7xVMlk0nVnjdDHtXqyYR3LUa6BfZgQEKjOf0n7ooifzJ3tSJq8S7j1V
+Aw4kR1KtrWDrtwzj5Lkn3C1iD976NPU/uwFmMra7sK2zXxPitvHwecS0Uy2cRLZ
6mXB8zKUznGLfKHEMak4GWk+rwWMRMCt7QkxfHqQlViSUNknOeQsQfwWl9NDZJfl
2sXYfFfH4fINfnRJ4zjWhPEoRqA3rQPBMKloRzogm4z+mumcI5HM6iJciswhTzPN
o9Gig0bqcwf0PGZkObXTfuCRcklK6JQ8mX4QEB5jX0FB/hKNtHdY4sGCC4U2d3Os
lsJKJ+uXLIu+ApXpdKED0pUCGNozme0LvIFrfAAwXbi0RnuPPjMdnrGWSTgv7aTT
MuktC5mxM8x3ksXE7WmQ77Y+oZ5R2G1L1btjaMu8n7sPc+zhwZBzI+fmIuzjlKQ8
S+k0umeJ32dq3AC11j2dt14J7ei1c214tJb6Nw4CDs5tx4fcvBnvk7bFTVNQE4lu
7M1CaCQW61MebGPc5z9EOB+wIzDJnU6Ak5pUMSRFoBDEdrZr+BS64w9mbFMrQoD2
UZesSuXbCk4vlIwtQ5QMM56rm2QZUtvuSsg1W0a5bIzsfmNeH+PFmn8y/ThEI/7R
nBWuJaPUphQPvrzbfthiTF0GgOPGaB8OSmTRwzNameuCRT3eGC0Kgm1sjA9LfVOw
XL3nuWrGKO7XultvHBHpXPDRN5d6WsQGwdEXFqAH1C2qDUcd1sSCIv6ZkLW4byCp
rgzyhv0irEwsN/ylUuwRbSryjE3PjKuoAXV0Nsec3/Wm6ieG0XuTsqkLJChI6R8k
8nMK5jAzw9QPferF9PMtEpI4HG/XHvDP3FcVd1SgswIxEWCUJpaARIwn0QR0sR6V
WlUtjLy0Jrg5LT/ADhhpSk9svHQA0KY56qyyk9RaEeBENbuNU74us4SJKtRuOFtd
Dxvc+w/SgQRCtzSBfkzsnkcEXUoV//WmbQEb0db5A/dWciBFpQqIz64cUFSEa1dX
Hr2T4P/eZXAtLz7i0N5DbDFJTWCiM9tATHzAGO3EzcalQksqDrArrYtV4cVTEuu5
92Dvjr4+IBcwRa5BcaiuSwJjF4t4pB3vrEJgP3lPM3a3T1OdRFl6io7GDfAvhJnB
9gXxSoWn8m9IVeLq5eodMWZ1o4GrhCDCvO6ALGsNs7nOz5RsB0RnYgvdjzSOVWBl
jQxv3tgcb3LpHoxV7U5ExcXzl/931vWVf5XVKWJSTv8XCeFixKayojaZElG2+yIH
PbHJtsAfu5nweumSwqdDkUsrQttSMd7057Gl5WpplmxFdgxGcUcRtDMk94QLfQi9
PoQdkrO41sj1mx/nkGYpBdjiPOhfLHQ7GtdKhU4xK3AViXmLQl7mIkg3Kxw/bCyX
lH5Ue1sZm+SNGap/tk1nqJbWWsjJtoiduZAfvUTy5RxsZPbJaJ5UsrKywArSkRJW
cu6AkTZIoL3zhp94uCyZfqRCwd6EGJhSUjm0MyfeLpdumkZwOyXcp9oE+wiWIOm6
Q34NcfJ43sm8OlQH0L9ap6O4SplsfukDo6QR+ujhNBNJYFjPbYgMHFXsQu2VO2Ct
E899O7XGMFp5KvHfOnAbGXyX87REmw5Qtq642ij4rBgSwVKuaE2I83N6ElotMdJM
j0wfkj64GK2IpYhq5MtBZN1CwLKjqFL1Ak9qLZnFDZj0EOXfR6HQUI/2XHfhILIC
g8v639EO3qArDxZz4ZvGJQakyhDIsG5yfkIokf/8QU0JSEvQnXeOAWcW4qg00Rvd
yxbGYoTy33wH/H3O+Emtf8JHQoE8mTg71qXf6lUunw6+vnVeAVM/XA+uBgJTPatv
V+vkt8rCU0UyKRHYOKxtn+xaOKu5ZnFJcMcmLe5Oxb/vA3oHByeF60bH7XtynHJI
ptsRjz2EwTyMY97DfmtJMX4cqb+OjxyCjdCvkkT5WtkVi9QZL9KalxpwfDfKz0LK
nVia7Xm2vn/vVUfh1hvTsHaK6QpQSfRFxS8SCq4kinvqmvDuT4Fifx/3McD1YWxx
q3CFb7klcxgSiSBzBnCvdWVRZ8qadgcTmN5dv/v+ZG0E3srO92Y6MNVsUvc9B2C1
M4PdBtF2Y5yZs0G5trhKgeA5Ewf7xmh45IhnWkFCjN3/2vWSIXnosNglZYNfon3R
+T7ALClIoCMDreTyQZuFNOLIYD6O1+mtuJMUEZHJrL3woVBg2RURsDngWtcFJBbw
4/WLteTrcCGd6Xb1rUcGHei3YghcbHLQwioR8hAKfDGEtab7fXddIKdQ4X4prFmY
wyJKbg7DSUl61Qo+ZRztNh0aHLMmNBZz5bimawVRafwZM5YQOBU7butpoJeY4tIU
Qj1wRdjJLsQZbXgA1TTUFlBXiiHcQGTRjDMEEiAah+5fnMGGtLRMsYWaB8xVhT9B
tuWtBjUUgBsXc92L+GEibrsTkXn0zmBO9kg2QuoSDRGO0mQYdBdRw+4LWJsndYlB
3OMVWedvnLLGz5Mq4v0rmT4SSamrrSL9IStvPFzLpbI7HZ7P6IzRrPumbE0F+zDC
eVqaEs0Y/H7whflWfsGOrRlOh7grweBDDuIae9sViGodLn2tedJFWBdSdG5u1fqC
TAeJk5i/4hleNIF0c7BuQDJZIkpprraAyoCEGaZivdhxA+SLtZZd4RSoCNNogSIG
7jAcN9bIu+d2lv9DQcpKb4UQ3N56jLrAf7Yn9QbpljRUvV098dTRZ9QgrmSDIcu1
GT8B6PJ7ja36Op7AI37X3Qwsz4ygQY4gzbXQjHy380X7KRuNb7Snys/xy2w2+Srj
BMNBI7oicVl9AwOL2Fdc7x0Bay18946rcd85lRE8t2ODwM8uCrYfemqrNAHvSEMS
yZ7XFTSa1qHtaUkjJlquSluB5lB/pAlTUUoKPfwFXTjuH24EZ/A6NWGylypLCE6S
VAfW3ioWHDdSk5XZ/5ta5MGNQ+xbNOsHtsJZ/oEK3gtnxF7wKhRGj1gwLO4QQvIA
wJQ3CB5limx8AI+lCA0A3ukiMT3Z+gyr5TjswPCNr+3UnPI4ZTfN5lWTg7WR8PAg
fNRECiPDPqJ2fpGRK3kMkQv14V2/l85wXos4HrEZbVeq+7jHvZCL6QikudQqwGMm
QX/KrDEiHEsRYnM2SosMssEnQEDgoqn0Yv6reNqFh2Aq9TnDVK5IPKtrjmpnykxe
J/JHOvOj8nvrk54E40TII/38aAZavg/ruH7PlIDp6xznHT9TA5paaq315LX6wiC9
s/IrEBCdk5msABHjikyqsTPazt3ABkLPyxWP/ZxaY/4LYd/vJ6KcqBlykAIgV9Dy
P/eKcSE5eIyXEQPI6KM2mt/ZD0c3isw7flIzhLCwavpITO33tcUdy+cMcgtuU6lP
hefPKhKLkmY4NR3F4lKbwB6aGcO9JRRA2v1SMwXnXzfri9ghNjkqhO8gsWmjYUdJ
5u+8adYizVD/pITthw4v+btlhsh68fHzMO6T8DQCsRbxMeYFs6fAYFBnpcgNmtGG
1ShQVVVJbXpMHi7I+ShZT97cMAPeHQ3fNq/7pEEtwTkujSMb28bxXiLwObDXXM2d
WnyGTiesExZULHJHA9w3kNxR4i7Zz5MKlnO7bL7Mrg34/n/Zf5ZE4DRNoakXpwoF
sRbXjIMOMfw6Lk823+T5QsOBwor9bdO4PKuxdPTiX/fpCgWdbaH+K1O1OYU6gDt+
DE2ZzzZ5EyW4VxK2dEC0KhVY8B8g6u5AJGGCIKQCoYRpIqsoZ8+H8M7uMJ7lFQin
iZhpLGkcPvj3edlcK3kTGF0PVdD25ynz8itXMjAkERtJeMc55CHLoe7ULU0zKvg4
S5DDyQY2F2XmqEGNDTpxIkyxSnvsXKCaJYWdmnAjQl2RaGCD0/Bb2Oeul3e8mT7f
dByKwzrCaNWkeI/Y7QFwOCkVqyRtezCaOURFFQXufPu6XAb4KXwwHCvTUOhqaQfJ
WDVjXgCrdW6g2bsEKJFHD8yZ25OS7QDanvP6vFYmdJr50acfz7y1YN7dnEt6SKh0
1zpvXmze/ih3Ce4uWdvz9QDwHyHf5hS6K2r4XFFh8yga0/UO3p1vHokVbuDkRXef
VQeqLyTZrFpX9Er9jjhJqX9lHXhndoTkCuY/SG89qN0SY+dpAnrsrU1AHnQPdv5G
voCs6Ve/Cc6jE5fmsxYKLGAEQrK7oh0seNGR5ndhnd2bRhhUOrKO0FukfNM4lEs/
z1ofVCwUFgIQcsx3qpzEv5OgClMnxGv6rXLwyndpVoFSy/c6Wj9NSBqIjkDMNRCO
TyIOQ5PoUFLnJ1LoXHO83XVYL4IL+TIENV1wTDuPWvw4hfol4gi+yMbkrPScUXcE
16hvkOBybqdaBMl+8I7FgtyMycpTnNgLbehQRBtonvX6Qs9juCMm0sh1oRQYKON0
o2wZ78WSWeWdCEONd2uChxBRr7po3ZEo53lYU3gU9O1wSPAE23Ksh+sebDDv7qnp
8E1kberE45LlSTyguGyEiFk7TUiO/lx7i93uNS5IlTgobCN2/1pLRbRASsB/hN2o
M/xtbq2gGKdSseipqJO7ql8hr1Z1jPXPG2sf/eAgwDMZM+hmtjSmsupunsxUAEzd
7zdmOGdaHAQ1x018NPO9YNqOU+xFyRSSTnl4QZFLWa4TkPEcor8yA6DjIyNqVTAe
bq2SNJce3aCh7Ucnc/k8IEHrMI2IXQ68ehH+RXF/sqHIi1PJBG/JyloJKLoIzgFF
gghGD0X/S6/N5kLgjh8a/l791DZaxATJDRoArQazUXqkImy8a/K9i2P7Ff8FRjR7
P/+y4tYdpsmNVEt0PqDcgnzSlJVBqxUwY1Pgxn/JrEUUDgQuvkucf4bImtgx6fZv
S0R7A6+b4xZfCPZdtgFcm+Vck/bKSX7xmtkDqsLczyZ4EEnAGDdSeLljEm2SPqOW
wr101aziJQvmoeTx4nCNhU2vziNOKYkgkqR4VyR3/oIgfOiHonBKLQ1INf4W4aGJ
f1Tr8VylBsCvNZxmXq550NeyQ7F6wrs3f44DpiGwuUISarh4eiSHq3T8POeEJHrj
ZSJoSBX5nG+Njlgaw7COr+MTAXRtijZbm28truCTUSuMkZ2pFfqvpszCQDLzR3ey
KTHXg/QF4l72taT498Yw2t9AhWePipQbWyL9bed1hU9QxgcwjzK45h1xYJ/NvBgh
vumgt1KZ2m6wzhf00idBpRYzRdm5DkuncEiV7fBR5QXqxdHrRDtABDOzzBeqt7a7
1V0PSagsv1dPekcGxyP3WevySOJk4lGLqON2/dIdNNvt6a2cJBHkaWOWc5lt2wYa
ki0M8QGnK96Jai+STg9beQ+uRqjq19VkzcWfyb2U/gdebJonuKDvCyP3CN3bcmls
o27QQGUyPZjV04+ls935HIlsXnr+lovbfmcz2iBU6wDzx/2LsXdEhX8p+jBIZn3H
JZvCeHSljO42X+Q2vXlByiJnjTg7JRZxSikYpDA/5TXlTOPpCubQByD4ROvxrPZI
939NFKcwUxmtYyMusMhU387N13OD44HRM9i8RRRVMGrLVXWXAtMHmkx+U5wR3l83
SqraxjVXjJKYGXqINgx5spAOgaMNA5fukFnEhEMWfLbmMgtqbizNMjWe4u3r90EY
DMb3UxtEadwYUIpZDwxzCupOSqoVrVwk2GpUI8GsAOce7/q6v+Kk0UdgCw9aePTH
g16bD/0yarwQjV+oAr/JkKxqPm5QKXvXjE9CofyUAtjE5zU82tBrDzuJZw5ySzdA
evbjsgKfnITFpSLT/2pNqZM641ADMRzDj9kLg5ivKSftVwhfMh5TMd0I9zczjM/y
lCrRVkRLciENhz86NQhQ+VfeUMxwyDnojsmfZAZGBgJndGmD2waR33+ztP6HONIk
HlRiwNBJg4RyshsXKG9LLw8iHgOWyhgfSoPLdNKn3lf3+orhkMUOdZvbNMHnh0Ub
qGh7pGk4YtmCbb5LfatAI0iTvvAFgjFmlN2fVxenvqnyMWfjkyfly5WBeahPQPzf
JZQ5t9+f0GBnUcF9rarqFADbvjm95eyEy+GpPnvPaEDiU5MyCGG8G8urS0l9q+6l
LeWiRa6jrMliUU5s8oliclfOSgvU1/1pPPFH4CYExoiPTe9IDNwhinayv/VdPgmG
cWt/G03jUyDOkzoI1Y4dusf/1KDgJ+Fbk+fLbFAriCtfzybMh+fec+wALGK2D8PH
cK3tyb4pKuotGekkt9U5DseSlJUX7K9mUKpabq/QDud4hvgVx1wsI4dSz0eKQuvs
J5Vs+3S1E3bFeoAeZ7sqAdBuvH6WCFbxuH3MhFeKIu3uZ5gI7CWb4cq9z31b+pL7
12mMzL2oph1rNqGswbwCKkXMK4EmSsCagiPKXBgDOkXq1mxhR4NPO3MxA5K6WjEq
dvpE7Cg6YF5buNyXSuS7ve/UK/7z45IVfzkd8W2kysCphn6vGgiBlWdDkSUHi+Bo
1vMwZXQvGpfpQAY8VvDNEDj9yGGaPFlxhcy7mhjsxxC9B2fSO4fM/jxWM8uX/2dB
6AHHXP9Elij+070mUn2hwegMfFZhUiyfvXAFM+UlNAC+L9Q0DX6KSfqOxQFhYzEY
x9PZd/5qEex7KWf8Ep7QOjGbJmH5lzJ1I18OhEdsfTV6VpjggQc8miw4vtHeg7Ox
aybZDV+NDHHf15EoKMYIew7UZPZxoh4TrPDPu3tCMHR+8oFlB4wTbDwSOgQULE7t
lcg9dXm/S4e6U0edm/COqAelVDpwa++41rcOoJfdVxs/LN1nbNjGrOK6lCuhT+Ll
zamMQkdkSZqVGD+J7eKY2zgWXPTLNn+PphofRdsl4NYBnWKR8ylBVydgS2XFZ/j0
wlhiJgV0cHAp0jHZimXb0JgmbNy2syYv9LJH2lPCBThQ/AEkp+mxLcdNKi7GxTFh
k5HuAcGm45L9Qkw6KMSZsrqVm0BP2AP6AgSsXcLQrRqVgDWaHQROUibr/oVBma7+
65vJ/lj4DM//xPDrmSKgyJ7HkSrrbNhsLxu31PNOSK7OJYG2ChbmzQ/z4vPvdQXz
CwkkJ05eeX+OuY6Le8OxSDSF5tAPL6KudbvuV4GWpH4D5m6+44pHsKWtBJ6H21GR
SM3S0hgWxAJWj66X1UdoQMlA8Xb+i0fqYyEPLqeINBRIRMhpCZGbBdlq0eu71ZvK
nWke8yHrjj5ESQKw5fj3fVrip8ZRo+qdZ1U0sI0oeXbsggT+DnB144a4Np6uDIKO
JVYrO0vv9cmOlgqTfyTT2BOWNkZd7va0k4SF1ypqPQ2tyIV333Wr5hqijvSARwGD
tJv7MNnLiDEqIgzFqwJxTVV5Bhf8Vu/Rqb8QGdolGVlo2r5qMRX+BmQoXpRNrTK9
cFUgWWDs2oYBHe+E1oEbopVP+ussLxJxqShlW3Vp/FHnSUmA5jBSd+slB71XbtVu
qrgJA+0ydPGoETj3iTMosqkyPS6pPw5+k6ghCsuvB8HYKadY8mzCk/YizH1mFEru
Dxvlfbf7AaUXh2K9AsrNFdfD9rG5TpcesLDLanhCezfaESZFTqpatOa6pOXWyC9D
eASXMD+XgOkRX7N+E6h+mIhLsvayS1Bq2iEGyaYO0HTFO2mkk2yjejFxfzUY3mTJ
KYKyX1NppKli2CwtKivJjcrCWiKvTLJ297Zdo8HZnfa0LrD2bXBdI6Rih1mXVcbb
rvSGt0LsOqR8e5EjUs1/8blsyES1tWLKp17afLwYMPx8/lEOr140fX97Zqk8YfZL
Ss35pFq9VN8oP+IUVxoLNkzODp/0ZSV6XFuX6Fox23RRSU5zPjN3dAijjEwDxOny
zU7dgCuT+fdCMXrHHGFDPvjaduzuhxbw45lhU81Wrqnm+2PVwULbZXAhCi+lQX3f
1Prtdgd121VrRu+xUkMpqNH0ygZgqkHmEC78Pq+QDE3Zsg/V3hnwmig+lDSyYZ4D
aP7F463X/DEHgcB+klC1tlj2G/U6VU57/9JdPRhal0bMpTRQaxFhlqHxwh3fB5Zk
yU5iOBbdrq6Kfqlh5ATS9QS3npwcBTvegCi4TMfSjsjT2X5DW7D4bVnxr3U7+6TO
9f8mFO3cQeNVTShB4eQtaiEWNAVe5l5/q34u7lI5K26Pqoid7Wb614qm6lmaOcPz
c2sQaCnlFVOC6kDeherY94AVgcTvCpJaRXau+0sBtHr2SCaSjkLZu9mWFFxJNESy
MTkeB5An+rFgsRH9RRgtJf1KUJ6RAEX4Hl018ZHSQkDn4pPwQRHUj+1Z8Vi3h6bY
U3jpCjfkdA7mHHWJ1rfzprF82KWK5pbkKeEfRsUbcrMkOqPMtnH25gaofL+9fO00
VIqNQ6aoWvg6d14wC1wLrGoya97vbtY76nhf0QcOoBWQtUHjPeOt01mB9cYcfLMt
2kYiZYEBiFlv71abADrAr0klan4yqRsV7U3CPg01mpH62JnadcEb1acCZCDjV3FP
DQNGSr4Wjq2S30iQ/k0bvcc1kaYecZS6jHQXq2dxTpIHSxo8E262oMlIb8Ns9Sa6
bqnzi/0opXiDqPg+kPKj86uyLl27kFlRydMctX8NWy00EU4ii71TeFSLbC7hSMhZ
qW+uUsZMnr8LvQ3w+gKedY1XurEE6fTUH8mdRQ4pJLY0NrnmnIj/gjZcZPAY/see
2VYLbiwap6x5QVkrtzSVvYGB6/hH7x6scoHppIRGU0c/6vgy+h5zr4waED86cFZ2
EtBrKu5xbFuGw0iba2su7NCLnrKtzNkO3NZ6U1pIR1XzVCfhfmE427kgGNeCurNo
giVtzvosuVdKznTKKkc19Wwt6cCY3Io6ac3ZT0pCSBj6D+2tjnAJqSps6z9fVZ9C
8fPeFYM7XbkpFTHlHlTXuGvMMGqnVBuUKSJIHXodXkcIjnN8Zdv6CN8YsmvOcvzU
PUn5IXQYexSs4lBA4IzKkxnBMXK7wy2Xwg1A51hFLTonn9n4eXYfrWsr6BZdpAwZ
Vs9JkTfbzff6xY5ioGmQFC+dOavNY+tsOdCd/s4+6Xm9eaDB6P1eDRDjTjALUhAB
4p+SFJaCaNE7dP1c2IUheyn7WbADP3YCJy+95WYyYVpViPfbiJqvdD1QsGtDQ5y/
IzhYZlJFPruD2JDoIWbvpWvRpWQP7bG+SBlElSUY4zZwHFwHAPN7j249u/nq8c/Q
KvKfdNDGQdEuXBWtR7vWP5UXBMLj2tJ5/HIGR5CzXhoPzcb7RX6Ls6E92Y8VXZU6
N5DWFKZoPv3okmS9AkdsaYfP9o5cMPVAVWxtXEm1TyITi4yFjqDFux9EMXWIXnxV
PAJRJJRCQ6ATSXAUn+pLRUmM/Fhor/D84UJZVIAEqmJ6KgJUp+xbnmOnMx/o/0kz
714any6LmqDQR+s06+aqHRfqDZYT+hnNzS9rosVVsnCyR1uQaYS3XHyrgFZ1jjWL
UoNmoefhLsFM2d2YbSzyLNKP1X3dmo4OC87U8GdcxT6cBsDp2aBJ7UGVI9YtFkrU
oW7vBfCTSug3OoPiiZH/53IzKdzQ/LLe18ST6BFVj6HuIx5dunyydWw+qdBuRRku
QUvJpP5TaU8tM819NctrNMjvyo1G3WTPL7EY+oVX+dDdGBTeeHLOGI1eAMgCgfxF
vifOH01Xvhe7OU7xUVVA6YK3pXEMu2RKmn+FHF+ptEjX1E5j+52OpjIDPgksfBt/
lMCGEO5Ybfw+Qfs+/flbCn/OhUwrNt2+bEKBjUpARnFHF8eGe4A/ISK7TIJBr2vd
PRes1LdEkHfEe2Ojtk0ewytK2yIjOjDJTpJFgpYWp1XTbk93gzLSn14krrVX+TcV
hpjsb/XkrOOMj4AMVsFZxJGI0v7KVpv0OBPUTtSqfZ6EmraHQmn7VjCcO6NOWXqV
aCLnIup4bEqaWKNMiIrthypUVguNX2J3ShSbOndSRi7Q9OlOnwKDP1CnLt/Kt/1M
x/vDFUgkYixnrFvi842Vs1ofCayhmkbHCI/vMlgJztNXtoJm+izxtK6rkgG0LQ/1
UjpbOv3sL8UbiSbFdikwKrcnlZwMhPakLRYXN1rkIV6cVE0wLXTcfx8knH+tChWR
MeozykbCvgp2QhjlYg9vk6aOB15fW2C6T44Nh/SlOsx/RYRImUALJd7y9i0gVpbd
VDXHMMJLQ90azMUHPiOjjafqZsPoJmBUzcofLJvJEt/WCLHQuscsd+5uaLTCWE3r
dwuwgiOG5yNIGkgBicG8+2svASMapzfo+SBs73fkyfNxg7mXDrQoICOZ183osZY4
u0dh3wDYYjH+eWS+aa6TXJYFSyuZq7U0iqs5mBjsjGh65asOSf0/d2cYrNTmaqcB
kutyddvZd2iXoxwWRh8hsUoyezpN6FyA94Blqgz2DCn73TMC5X+TIWNb+y+zyF1C
85KtsQgNS3nyXosT3FxKf29y/dFKezyjbpDnc6elaR8v0Wao2c2n/IErUXsj8eKl
yxdySgYUzTVFhB9YmWWGB3PhGanH39u420MRFnIFKiXCFvf4h8dbm4Xhar6gK6gS
X1xBWyu/rWdxWd9OowR/nYqPfPpApZlxkWtcC//oTBdZX5SE/FOAck+/G+3c4wUY
Z9hK7ETaOQUeYv5oNPL9JG6BdqGRXbFZeVWJb/QeXktY0JE3HhMtnfwdP4/T6E1t
OLi3guGVCiuSauRPeQQB/ofZSHGPdccHXVAcMoO3bgEQV0ZHJuX55RSBoNCQ39WZ
TBPeWWIeiAe9EopF4zu830xEjiCe6/DfGCuChPQMpwJ4jnVsc6c8i0PljxJ+tzPz
/gvGjVqeF+RyyrK1PvT/tEc7jaCxG8aW1iuDvjHpz2JwqfzoHjVL6tMWZKzewadh
VFiOKFqcjuVg8KAtXcAGCEDCcDfMkseYDj4aEvSLYiIf3OfyB5I3NPUqGPDt7qlS
kL9EN5GDw0AY+MbVwNHHa0BSpgGW4ezLivzPlAYQn1uT8UYvhQwK6R7Qs3oQY4SB
AawFxIfTkGMSNRA3KIA/2bG8PBamaSaxYf/axu7aKDhuAy/dajXBXSpt7ySHQD6U
OLZ/6m3/wd1d3e7cRJQnQ8lpmMe9Bxzkx/X0AyMs1MZYLuugockgZXvHQaKGcrVN
646HXqlMXDcavdtGOEDuwdCPnQ8DYWO1OhYSThxnfsljs+HI9LaZiPM/ypTbcsIL
JbVyzuBj4nS+T+zVO24d2Y587iNVTOCAfsuk8JWI5Nn6LYbu4n9ZKtvA3ID0ud7p
Y00b2sUss+ElOVKeHOVPYzYjhrn0hcctrwbFd7/rvgqFuWyvNV9hkQZz4Witn7y4
1h/x2gLhy39vQu+r2+jAVWI7ld8FStB0DhHMSHMdQRU75492uTVIhtgi8/Za6CE/
o4AkGKn3GaMmc5SXha/UDCk5+dN4Pj8/3aQ6vBOzWXMc6zyoynEp03bxdmIe8C/X
zT2RiNPJclnruclRXDj7Z4OxNUwwFnRyTd824/JTiBylwRY02K3sURVN1WXHMevg
Vmnmy7YJrjSy7dNkwsYEmoQ0TSz5/ifDbNDPzoN8HZAaoV8mc4mjmFbhJTED2qzM
8Ez+4AI99x21ynQBnrKgYhgnu3BRhhYZmJNQO13lfBiCgVs5Ujw9SN9LB6h8rW3p
7XX1WFSCrfp0iUmdx4Vn8DUdwqVKQpTrGUi5EIS4ftD7K1wqHubKhie+Iprp9bz7
KWUSZw9AJVscvFJG4w8o5CLJQryNaJWfHjSpRNEUEqwe6Mz0vhf4hvfJqXjiE+/e
35T4s3jmdJ/0HBrmSNxL/BTELeGa7XSdECEjLdXxIDipkUcb1lauJZbPTIcBN+vG
/nVPR3VY9Srw2NhgKLEK9d8jx3CUFzy/QH2t4G+uvr6JK+dkVCMzA/x4lk7I4Nx8
Udgc1gx7wLl0WtTzATGpskSpgX7/dejLAYmEDEnvBlIojmtR3dKzTFa91O3TraZL
gIO4B0+AbIxDSCLwP/4wBOHw/ANmR3PY3DUYPakx3K/wdmCq4Nj1X5V3q15T60iv
0xSj6iJa+V/8dCAc8AJM4INQ3UtcdX7jCu1ciPME92RQm6e+Cq96ZzpaHJJ1bI/F
6yTnSBapY357XpuS7f4UcgmaTyclQFOEbDuRhVgTAdBcwRDChAfldSTF6C4CEcbi
eU+HhbEAa0qy7J7kXlYsW/7ISRFYf2qNfKpGeVLh70g/t0CMvHsGXorx9dvQY09Q
R5h0xi/Fu6bGSQfn/kBNgNVJQA5MUL/ktNo0QW0ssyP1ZePTq/yowX/Xliisbiiq
4gFaDgp28FRiVeXV25IQwp5qVU8YpBQD/y9l/GsS993pqfGlbEHIng+nERmveHlZ
dlCmxNSnbEeMy4o5wOQUJg/joAYLncTKnk9K+8OheTfh5oxQhoS5FpcbtSsOiwHW
lQjfDJU2sfE0yBINO374rHGN2vF/mlc06IP+nxQxIOfelbObXOWSXLMIOiV4UXaq
c5zAarsLl6EA2MBiYsAKgxJQN+I/RkfWs55KvuPjURHMmG45YCotn2fAb5+vvVEq
OzAPPS0+3GJDWZbYnwo/LGpMOGiLdQ6MHj5LedjwH2WsOORJtAU0bfKSZA2GrOVz
hG8MibhWiXRa9BnsRSwS/pXf5CcD4H0F8nuQnlpvnY5zWcY/Gi2+GcqTquWvtG/H
rTZtEEGMESTkCDeuI/FJ0iGnLAq4NZPi5uSQ0yeSrQVyQMRHnMsaaaT2aZAcV80q
mj0+gbQo9tO6twykeljKrzeKLSA2Ig3SLtokTajFfMZs6OxCBi9eLRi0Hqm7I/AG
EJIg0hTA6kk4Mz4vBLYwmvQnWAF7xSEidknMsyxbgShZrViqJQzNTl2hGAeopLaW
bLrXNNDEFjn21L6M2LGeL0NiNbdflfmeP+qcUi3ur2+MsV156AayAhbnwMw0J+JW
k1evch+yUcIC2nHeuQ2lebnchEQ3zmjk3V7kCkzSOMilWTEqCEuf6T3AFHgK4hqk
p9EcHe4YA28ycJLUPGdUaIKPzThYZAw56hxitgW+EvIlV0gPxEB0IjwxrK6FM6cG
ADIifnWIuaMhsS1wvTkdKCzXahgGXQQlDUKs8vJrQgaHEX+r26WYTIncg1WQN6Dl
/OTcoZKuLwGqMq2MxMWK+/Mb96zBPwNU42LLTuz3x81baZ0aUyQmwIqJCLW0g5p+
+t6lbvZjaFFr8PAVdVBBYjVuwtz1x3v//mGXedJuuAzl36H+BfkXI6TguAzmXVhI
jGn4I+ntIWqufI5Riw4O2AxnC7YvaVZqayr76cYhdeas27FvN1x6REfa3VPk4Jdp
vuensyH9S9aWCgSjU86tj+jS8wElIXEdSanYOaArzAOvIBGIfxl5ukmOPXPiBJ8G
2L+ywNBzn8DrFVOs6PjLbqzufzR2f9Qxd+85HAb2FfcMiefEt00Blg2QxONu+30R
pTw46L6Z+6PEEr1V6v0ogp5YT7ubjrAXHCWgF1pmZ7jeG65uvhWzhfbldyC7m8nK
pX3FQ68ezn/JvhC7+6CjvlITrPgvxiwHDAkWARwUGYV7QK67F0AAm7gkeS9ZjkKD
xT0zRmzJDZQFTOM80o+YXETHvVjaHIPYJOpWSJVELJTyT4Qkr6gkG5tP569itUj5
bF6XjpKgNziw6Zu/81qjqrQrwCXnrwyks481MrOrtrTwnvFUdrEXvn+hkSuYkj1P
FhE01bllEhSr7kyw0y/mpWJWIinTtNHBbi56tZQvhYhJeUsYw3ZlzbNEJGf5ITY6
ojS8C+mWFU10ZBH7rYL558pN7+8YK0mZoSPoechnWq52m7fRq+vXNwj45ogFsmWD
9MaCv8bs7HY2afGyt4A8TfdH1flEA2wRGhFnwmlRHZ3h1zRTPO2AfBdRkZQStuiW
Yd3QjPCKVWMPJomvg7tpuOEmNqonRgnI/0vLumxm9tXt7A1yp0clfokN45rexoYW
Ot82OJEadV3yIb8Fx+KksWbfypcwXDhUXv4r0eiAiI4+qpkW/m8pkIFRWDYf0Wtg
3JXEkxahZePucLFz2XTxxHkskNICQFLb+B8Va+F0Q2eyUKin1nd1aXfaGHkhDU2H
bph5XsdrR9gkAcnNfpzplyNeXHTF9rM42y0gAHUqCew9RBBDLjLJA+V6HRAu3R58
8ts0fzldkYtaHfiqkRJjzzu5NaFG0/jq2yMrTN+9eYnWBabVe7rej0CmG935pOcQ
GDYDweQQhVlUhoLk9mlS+B6I5YknFAfvQWjRdoCUsr313muYnUVVQmzIWUH6dHWj
GJl072nqRAlTghtFXrLAdu4XWpzXOlJDO2uxzprFuN31EIOuEfv4oGTl+868rmCm
jpL/PxHyK01i5Vt+EEKhA9SKrop3JuuCnewkOF7ADPdKiFnGmD5Ds8GROQte9BXc
UiHqpuTCNKYF2T2CXbCSYkliYw4O2gbZZHnIkgpOkDrKTrl8DX5kCVaWZYbzUmhj
qbKdDD16feOfXIMo/aePKeYTQfTPPeLaEScgMQgnMKD2aV/dGnMgaMDdIaeYhpk9
z46BNka7vGlCfAOT+2P8uIZoMYSgkTPxytcS97LCIw9TfSCEe/EptfbozjA3mud3
HWcLBdvOXhI8QnsvGxUe4qterlsHl+YIOGXd5agNY/k1Ti9KmKDruQeJRkAF6pkK
nayg2+8QSLPkqBcXJysavqt6YDyRtpmTu0WaSbf6mhOLBmw2iqCFzgdTr0hgSpPD
fyy1v1QE6MIbrvmwFpq+1VrQf46DrFBmalfteC5UFP4xC96O07mShmwjVa1XgOX2
wAYlbWhnQpsJOAL3oDLCe6sWlp1WvPDV8zmhRLbxmatPCd8/aRXZIgIcBm3uM1li
5D6jzl14//Vh4oyMuomSPIlGZjictvlzS0VHDdn/uJ/K3hyZU97C1HbwUyc+Lv7W
KOj0Cl85PmPDn5UZUthCqMWufcnjv1K+m4IkBbrwJ0oLxKG0Ydg7MGGJ4Mq0hBSA
ZCKP6wj6pryg4XQcLcg3L0GUvALzoI0pOI0YZbzZqoXy6VVe0PPFEgmvsIgXKNgb
qGUep8CDl/ZmwYebsUVhkFwa1RcB1SG+XKLmUYyb/an/0d16pQIomtvXnW7RPdSW
rYIATvifI5U9o/3CVRTkpntKJMO1zDhbjOclMIAs+hjmencA5KzImPlJdX7Zv60L
183glOzImo21ftf1Bv/cl7ZTlc1QWwQTuZFV6eD6X2r9MkQdtd5OyASCrwCpyPSm
7EdojziK2H4Ha0ZoG7Qp14TxDEkSUkLP1NEypKh6+euFlSZFqJMX4NyZB8GHhnUu
diqF5FaUB1cHDxzbZK5HGOZqWWAbRZoEqBQScbe6XMuA7Rpu8235/MKUkwBPM5kj
sD94vsJVSheq71Doie2C2gAA9SV1jm9LHbvFk5Rw0MmbELFdUf8fZl+G7rTUJ7JC
CB5iXXmWcbOA3PkYwHtpCeaccaanp2KqTyQ36BMyT13kCVtJxF54cnvz/M6I9rsA
GSGc0KKSxM191kyjAdGt/9CUasXvfoKwC9Qz5n8W663dvUleDLYm9csojzTu7vyF
7bUf4DwQNWZMST/9gJRZKx1qSmkJHI0NKanPPY4x85D6QgOahlEU3LqSqTuL0bbf
MUsjKEL4SKS1t+Hd1onZ3HK/9dUPsDdta8/pCNgpHiOTlZOSnfkXabT/Qhwtrx+2
VZE1F1SMO2Z0kEef1nEE8Qs5dQEBbusxzD3XPrQDzXHOgsFK8dESHnXzNxcpsGjn
iHfsHd5cPUEZ2zX+Ymnnm6DffYdht1QIHNg4LB1sruxm3hwjcnfvCo+9ZwtnpUuT
z4YDi9ez5mqujtnGV0A9MD/fb0fa9w319Ym2KzLHZjP7JnZjjK/XA7DyyhUuW7jV
Dxa0iH8MpeAk62dVq2tiJeBjFaHFRHZEqefvrtL7w76JvG/+C1kkbyK4nzpWrcqy
fQy5CgjD/Cgca0Gbm6xtE55xOrB0C0Jph2b5qXSCPyHJcMfwIl3WSxSMCqpPJi3o
ToBvGk3Nn74P35GBnoLNr02cv4jrXD6qw7XwhLJ8oOQgLY/NFXTlleJ2h2gTtwsC
4Y8VoTYVcULxakvquySrmwoysjd4hBmZ7T07A5ZTanc67Lea2yjtpF/5fSWeu4oX
zS0WB//7htk33GH+B/BXWvq/7vxFmYIzGiOcXgUVX+MwBcRrpsQ9EmLUJ7zxFYrB
qwjGWg4yEKqBAXvFYWpAmLhOaK0rgokUETOHGB0+SdiP8VCIk+3P+nknI134f/JF
IIRqClEANS7cWdVhP56CIUfrwbYeuSpjOUQg1TaB5rsn+xMjGUmdE7HKlS+vF0Tm
Je8agqKVuuLCJt6MMEFAts7/cl7TtqPVDB6x0wBFD8A+bCdzPIG622RJ3JU4CDtS
dRecOJn24vBBphP0hseRy0J/eA9qVBMBlc2XlIZs1UHAG8LoUMOiNQvmEIGSvJrQ
192XE72jKqVEycKDN9/mRkzC8TgJbq6n64r8x+CayXz0P8kXDbRmjKECKAUV62TL
NezyHDy14GNd03DTslaPHR/kVLnRo5djx7gZlh5qd+51imT+f+MUsbpsnMk8YABl
26tAIVkNS52wgCuqdE3nYN0L1vwPeYWHwJapa3tcvf7kZ9PCYBtmZU/8VXeVDahz
x6H/VvivMvj7nagcHI45Gc07YO9W02IWCSq7nIQFS0gqlNpwYF+onfQ+rCK+RuFL
6vjGEbx5xs8CycHr5zr50rQxx+LeGRu/2PNb7QZpDM9NhYeIEl3o8+70dQLIpk32
XaYjoTNNqcmy7Um9cdBCa82vRNSxT7J3KoZAK0P4fzHjSJnly8G9WwRtmY6jS9Kb
86Pp2wKYawm1EnkN6cULNg/pZQLjtaxuuOLYXRpYPmLWjoKHriZ+Z5g2qQlRYK9+
BQ6gRzQa30OV75jnjU/dAOa0CuVMj4lj4ltvN6l7ktGuI1mL/tng0KipURZGTJit
sa/2n7SIwEPMXs7fa3LghOcnEN5elxigDPLX/UC9CEcGtoElCi0iaTwyHl8FfZLd
aJqctTjpzvMbNor7EifrkUiBJBbdneAND3FZS6h5wQpE+0lv+ta3q3jnDPy2BzvK
abfjYyaw3quU/xeWaAsoLracgUAC+bk4TOZDc4fduZi0dAs1NxvhEMLQ/PK5x6iH
60A1OZWviTbG/TsUrdrr9z/TuXQTlNfXQnaJPoIu0K2PiXEWSP/Kb5Zr5n6191Ll
rayu8CXtDSLceTDIKe2s+OXF7AO3uSKvMx3V9nvLSOSEpFT4N61lHU7lOy56xYOf
yrlRufxxM1MKuyaKxf78deAdHI6cSiUlJWzPCPrpSAaSwgKAaloT+TSUK/iU9Qh9
qmm6ioPI5z8iyTOMWTzUwhp6FpYQEyNnypPOHdbaGryYThhhnglXsisHd4Agcg8q
/8tIzdUeHzpzbjRZwNCNdmMusdfOQJ2uYlsV8NmYmQPr71KGjhR8Td7LSP6gEwj8
QsrOaB3aBEyJRHacKdk0xG7pF3rGv35LEMCHcuzidKpmSFDNNBkixRlK1SI6ez54
M91BEFf93dl76kc8zHpVzT7v99RRhg0TMAXnK/GWkL+vOQ1dcmieGSLA+075dMJv
KBjWLPehGZVIWqtUSYHMJh4y9sgBuZ3SLaz7tYCBNw/WDpersz3HhJjYX0c1pqFB
zIXa3Qj9JMTCQ11LrqFNjAZLZmirz1ut89c7SsWNPgOuQD1AQcX/T7sgYVn7/xQO
YT7dBISVbq9TujGQUcrp3wWC1y7H6s0aIcXIELJdPLCbkEFHF0G9oRLvlf3bUIkM
7G00K/rO5rZloJYC4j9KhwGolxYnoqAug+OgfWwwcKJeiiwvMHTOZ/JEG2eA1u2O
12xyVJlMkQQP9HVzUyW63tetRyYqM/duYtRoVS1ekJll0zbIRKReosz0FHtJI/ra
IEOfgis0PsdlR4pjkiOTwnbRKluqvesF9RtCn8CpSYsvE5+jJxf/Ycr+r5eYSdlv
1zKksejWNOFEdysXrK81mfLTT9LBa/IDj+07MC0shBDseJzEpMKEzVAhbwlkRzL1
P7UrYPZGtvOGOjQvzPk9quoNqP2SMddziAowUEdhBe9PCKn1/CjOiojWlmKXdYcw
RoDqPtvZRY0WJJvmR99vwRzsqcGWOD6A3cF+W548N+Y1mp9brYH79WHffumHcUOk
nCYbPUXZZi2vF/tvlum+ylRoBYb0PHGbtNMh0U/NyyKEwj8GiuV9tJtTfhwEwIbn
qAj93zu8lEH4Ghm4/qxhPp+T3fRYOHu9ez1jUB3rJmKANSm4UwRK+R6lp6FA5nob
+sVokBmossRUnCGfLAYofLXNqQTNCGtIMHiRcoshKqeC/LmXSCIPfvVfE/AdrrgK
pUoaW4k3J7RoIsX2kKsvxTAYMvls80irY+BYw+QRJ5r1NBTot4sQESSCZWOXMraV
eZiDfnApSISW2U0IezHNxoPiJ4NtIYusLLevXbpdRXTny+ix5LPx3LzUjJ1v7/jV
A97+8Tg7jG+IaVPltzWjRkk51y/Md9361Yrf41nx1wRYtAdk8nSxENK309diZoVb
oRDPaL02HRZS3QdnBrPGmHtkg9EXZ62kRAxprK2urRxnFMLeEd/OJ3cdYGX+VnSm
5KP23sYwqu95eaNrnlZt/S2+49v99PFKMaRAd0X9PogWfmvrSRUMcNhVk2bM/Ig8
EI50J682KnrNeE80W7GFd4TginpYuCxB6WfiJQPeBFSk/9bCEc0AYLhxBV8tHbhO
1LULjbZvxSTMo1Q08uYl1v81c6CFL7OqusKr6ek066jxpjWg2jpOjC5LgvJevMbB
YivoWABzWyNAi4+XFVL/q9FwURceeYU5boGaTYMaUs2Ee8rmktGHvmtz0+CBur+s
PITta3zJJt6INvSB3kEr9TRvE9SKp8eSupRUx3oQkmj/yUTwLlqyalKHnqnZ4Aeo
n7vKugYdupe4oIDQ7aXVBKvuVU1uRCBFjcgpgt9sEq3S6c6qNPWR7JKVqHTa1jzH
12bPD5kZFrZ1ShjD9XB05G6uNEncXYslLQ4QSS4gnQC8CXglszKq+nHUiKMrwTWX
5+5RZ/vQFCeiv/8NMcJcDp6JXZ0guWY4sg03ft1QhluGNt+rDHurOl1JTrdE7IEC
yvJ8i1N4u6t+nLbVK9kdqZVlPDPKzTt6nAsy6RcR4JuICisvpsbjcYrDCs4wu15m
AJrqbe2RampNYYZqfW9VrzWTNXHClvgWzSTM+hu0h3h/g6pdeawmPRWY8ZwfpwqB
RyAbiT3spJfA2ECf0nD6Vs+Nb2x2sXqUz5dXbsAVUhbXRtcsLJR3/ax2WiDyLUCZ
q8w862K0RL3+b/m7ApYNX5oNnFGhEFsi7UMz30InwM6dcLdtR6XE+j5XHUC2p1Hf
e9DKYAzfsKjjPlLQHZBddu+Bp4SEpZEX4UlSeyfy5/4NtPvedWB6CD8DFxNaEyER
bA8t1xh2hVWHzM7IXlqYpIw4GsspTcsFFvO9PeLx+YgzjLS/l7QHklpjfLSdyIP5
L0EB0+U2j+3gIlWeSeVll379kF44jCnFlj5QCHAqqdbYYGnlrUwRH+dJbzXyafwe
tnXZmcpSgV3wuMCiYJmWFIutQeN74f93jt8eWNJDaLYo0BiNhEmoKp1bxAEUby3l
Wq6BBjAqkS1ZLs9FTBCy6H57bZ4lIE244BY7fLwElmrI2lKZyhkOQ6R9+YzSdPVT
y70VhehA68MNOefRslE7xtd2DYAaASr0wNOpgIQtaMxMxm91MBbfRYpRRV77JcnB
sZp+IiF1FhZnmVx6yX0nIOW0RfEcfhZKKZfVv+wlbp4GsauCExVNcLx+caUu+hY0
a7sQ1OrOxUIAcCv449DCqq556UvA84lfHpMatb98WItEbp7hhL44M3qnb6tdQWNi
BOnSgjK5cNDoh5EEEpAk4Iu8/SKHYLCB0UWL05Lb+ncWvmtlJ4Z1ooB/bOR1lHhf
21b/A52jabZLQIpJ3oYBaq/wjrtZ6Z5/FYu0j7RZ8yACT1ft6tFFc8miFqUN+BQt
BKg3cm7tyeFGrmtB4DJTM98xHhYlftC5gUkaL5TnyyFsvMHvMkSx+v257k2DAGuo
Ejv9BAo9HW0HO1bGOsRmPcpa669mpu9uU+lkmBhXFNyEI84ePagXVuoY17DEQ/uU
7PlEYsygDkkYB1WfU/GhdQfgKMsxNJhtbd9RRFyPWVwE4O+poTlUWAsEVfvc1QGg
OkTV6FeGQQM8Y8ojKCSregk4f7U81Qe5pb6fjsqP+nZjd0G333JnbXpvYVZDyxH9
cRuZwFdxBuc4f+NGpCMpxCalopZedClPqKt6sT2z8A3lmQ3OOiigNGsSwjk4LthY
bJZFFsg/A1ltpCh67+ioQcFy5t1FwOF9Is/qY0N0ujBAteK5eqVEBTPcioPNFTYY
IGhkY5jRveMtt6S0rcjBGA4BWyq3KBGyWZDZ3KdSaS4vn4QdzTh6CJj7OPen9xFh
4y9jFkgkIIy8Cn8UEC7LwnITSlVHAc+dhvK68nIkCT5Cjoe+VY5J18Urbdjd/I2k
q0AgpIpWbvPkrnz1oRSLN0ddf4v4Y1TYJxGpc/qw/2/+8nxz8N8eRX+1LumKLy7m
PQt01vE+sZhUQDJR47BgzWWUcYVBOYJYHzZ25By2w72rE3aqTnTArb1kmwKx6Z1l
UI1fCZMEWcCbMfpnClUBe2BX7qpwo9kIxUURGlGXtUSiIoeroFFaC0lmNcQ2hKLi
n4jBOcVltWqB1w3EVqln6Tt8+IZxU6Pp2Yc8VuwXQRU8m+b2wNJCaU4f+AA3//B4
seYa8BTZKHkqo5bfjL2zYlS5jG9ht5vysTVH4TshX8u+mflppNySrAjoja1znE4e
19OZovCG4jXsHtqRKx3/PTYu5dveeaWohMP5pD4P0favcStOQ2t/Xl3eTpf/WSCd
SYBKIq5kjoedWWiG0GK++bNW6SGpD6hIav4jpyYiIw0x7P6NhRuIChjOo02E0Cj/
gk4h5Mxlcya2NehkZXX20asmd0Izt/onOu2OQN+CusObanpCMJIUO+FznAV4YF3Y
mwSS86+GxluRFfngdcJM82Xu5JhI6s7OrBLFbFHxsLkVg8R2HXgWIr1rkMgIYApJ
bS+fvm5LO4zcfziU78ZjB7p3T8NNpwRu7fc0LJhOM/epMSF3uO0Hr4Vgc/Yu7oZx
6TYGuzRWoZ46Eac6g4qsviiqVhD+yOCzsQ+scJVgQNIXdS3sPVb3zbceYXCrx5pK
6hH8I3+3ruPIOKHMinIX5TNxomCI9WcnltcarUblEyOyW0unrK9sV9corNx/ZOgB
o1rviy2jgGhWeaxXxMUatJSu2AWK/UzcYE5TKbAMG2h8zcSSCBH9CtagwCqA+Kgl
j+WrLG9Xc/no/MZGqf92NXMeslDioPyj9ESS0jqaW5yKIP5i2Bf33vulWDmrfIz1
zCPR5BUNCpuu88ZbEYcOIdrvuAwA1YN7rQR0d2XtvxS2aaYdQHpzIH550nakngTt
rflYJmudkOAEQf1YDxu+jUi5oyXZw1zWlGzW18/jZH01IhvZYewCNWUkluBQ5hcC
oMDOXBbu51779QmhO39ykjf+si03vgMA6LhDp/iNgTgW/ycFLcZJ6lhB4wL8DgbB
jJ38txe6W/Ptozfdd7K3lNtn5tN6Q9x6a7lBhielPE21bBSvg1ZHs4ZPWEQ3q9Jm
YrbixWyopn6EcKwWO/lGbIl2xswCmuX6nJrzV5+6xvyUP+Sw9fR7X8UOcoNxJqwA
b3B8FXF2LjJqQNUP9M5e9Fuw8waVCxy/bfFUIPEjYXqb7kZESLVC565oVxJXp2Ve
WpyyOi6a0y0TSkELCKSNicdIHmn2cmYNZVjvgAIJPp3jXrrvRfeX38/I9X57fbtw
iVUZtaBx1uUizKSjDd8OS+LPF8kcvy6Ua9/NjxnfOskLwxy0p27osIBhyLdrDs/s
JF3fFIcjF/pT2S4OjIV6IzgNbMEAuqfd1lrCIO7e18CWTH1x7tx321oIn9SkHIbR
fCDaLkKlJdMGakNrAGv83S84H6csq1537ONtbGBy7d4tYqWyk5AEBT0PkmJJyUqR
O9MgRz5fDUv9ssLbRV8JB0nwbUNJXK/m1VjCIqF2xfq+51yWOx+/V9nSPTDjORht
rN74wiKfR4nzCAKHdcI6pG9sHx1zUWpcZIljq8urFcPPl0+Gw/p+h+W1u9DHuy9S
eG0mgEdCVHrepDhKTa8szNoNc8E3gDjNfHy6MYMkjc5OhOP6/i3ba3Wh/OWUAIT4
QmeElv5nWlFCHIV18xv638Vqbk8x8Oar+xpxVEiNL/eWCK/k3OX3/twHsCUUroBD
oKGgKVIr6rsiNjjB39raZoYvXg9Kmo93atqhSQCt9OhUJlPbzwLWjwiukp/BRsbF
w5IMESJIZ/chBaMnMM+pLBDh++fLBDa6c8YVgtXYIMrT3J9v7IxUlaCxrRkPbbdW
2BG2dRz7n5dcKDXW1a/awceGiBe/Wvk/rHbooqPzbsBe8jX9X8p3kv50LkVCw/8o
uFMq8azFJJMnXDkDuEwnIf0s3pt8DKXeIPQmJFvba2gsGwy8wQDzMic4cMPtqsx5
D6P+t1UkWQheizcrQIYd7LPTFpEdiDApQAxRCEarySGYRNebvlO+v7QH3B3V+TMl
eRHtrWFsfaPSvBNJTl8oib01jweWjJy1P93qIi7XFAgSX1r3voKYAjHEt2C/HqT4
jMzR6xVMaa5QE0u01WJsTdDeD/ZmtaVgP+EOnmrReOC6LRyKumw6YPcolquj+sw2
gfLmp5B3jPlWKut4pt7ysHpCklfNa6nxkmXMcvOAXI13l8YG8I9ZONnKQnNS6Euw
fvL3y3rIdJnmcBWuuGCAymMTlTzYlz4yPPTv0EGbaK2FMCguLwZdR6Jbj+0Ur58S
JhLJJ2Anv8Gv8NIfHWRj+EFDnAyQcwjWOVFR6hLBfF7o3Bw6hxaVqyx2WQ9KdGoX
En5SFwB1LVUVEFIi23aXVC/w1S/VgbOQw+c4rk8Xu+UWMhNfK3P/AuMIEPWvhJ27
89AdhqjK0aw109yfxAlh40CrpBP/vI2NZEsjK2l0dwUqK2NSubbT1lHxKhMpSGOz
zf7KnUS0AHXfNWLXF4I1VUqu0itsP122YbHcwMjJoPK/LMRbNLAG4N2B2TJhZyMt
tp3/e6XirvfGsQWCtVZfwf3Kq0oUO5DXDAf2yvaM7lbEkFwgsfzfJOF9hJ3LWyLZ
MA/R3Zo36+fgBr9ZjuLBs5OPq61ILREnVGj/dVIeZ1fWCI7Fy1ZkgP2Gvj9fjDCb
P+9uwPI5D1whQSh1b5ThOKgKzf/k5ghbA8stKQ3j4HObJzdTDl+6mtaTHIKBlKNf
0OMeq2l068x6lGY1h2Y/X2d1jV5KrfDfOyXIBbDfEQ5JlO9+E++8ZzqYNcZB2h4b
T4VgKHeV8RullXaqESkezFw2QhSlTFxmCONj2VVESuFRk8JaAzapJr2mfeskKt6f
XuR3N524FzJX9cP9WZwTdJ9/M+XOzFqsaF2x/xauMxgZigPtAFOgR84Eii/vRA3J
qG5vu8MtMqca1ZRCFSk7TwZSv0tDi5ex5d5EpWTrHBq/o4m7bCTZH7AKGGbz2LG3
nJ4Atjzxl3pfFj9HPMpJ3Co18rvYRbJDHhlHaL0fInmOqWL9TohH1vMuCSSet8k/
rqvuKAiyKivjnQIdQUPtaQeDaI/dZQTg5xURRRso/l82etDOZc0lJdsd+6Pm8nMC
W8ilkr1e9yC6BD//ia9pF0ciiqk8B6MEwo83dbN3th+Qc+udKvXjgB5fI4spJ9d4
Yv6u7PFdqqiLm9TggkdfkRThG9oqNBIPPmmZEQa7p2Eoy5RNIGY8WJ6dGDz99GAD
9M9Qr+KlL/6Lf86Ki13l465ugm7fjZxc8aJHBeipTXAkkiGkUVSL8Qrf1UhymPMe
IYPmWTvzAAVVxFWAmQ9MZJPZvhjQ9eRlM/MeFayKi3Go0Lbbrxa2XqJuEwHr26/Q
0GlBv8+bJ6zBkaAOsJ2X2BxeabRHu5OU3SRK35pAo0bFKziqXbz0SEAkOHx7DzCr
lgppO2ipJ6UiLn0PUEjWQWdEZg0CTgoL+urqGKkDVTVihXpAAC92JOkvGksNd8ri
P2vD/blykGnquanLb6UO6vVnU84ocSV+eHKaQDa4KAA/zkH/xet4XCnO3P6x+Z/n
P7pvo9z+/e7rVxQXHY/Tm1/LSar+pq8MOlSe7wQeCW9mSh+36WAu2P9UmgI0X6F7
TvDF0M5vIq47nA6+mW9Rmz0DmwFaB/f6Q+X4QX9Kl2bEjfu6xgWHB8DXQP9OeaCm
eNKR15uqiS1LEUEGvDI1vJf/3Ae0sVMC/8ccGoj6LVM5JQLTJOpb/um81e4RvX0y
uzcVGQNpYCwI/ij5AEWciTt2TUpvZxz07dXF2Oqs2lqhxMfeJcjFau/1LaRWH/Fd
oglKxmeIdcE0kxJvBcSMs4k9yG9op9UdQ3qSSaBHRltbXyAK0ZZjD7cto1Gb4fi1
egLGAWhmZ1Lp1OnPJ0d12CRPb9zNiqwVc1kOEdk5+Zt2RvTRNrQ9zHSAg1Gr752a
B2FJrzqP/ksz/kI8BBFRXQxtB7f5IB5jTCZn0Z/806ECIG9vF5CJ7F1TDDg2yjtt
/bUmmQPSvySEArnZn8BHzdNDBT9WBAo0WP+QMfCncH4WIh1gIPMnZ/M+VfwsbSD9
RN2lYxffe51dcS2+4s6Fe/wG5y+t8+CBmt9a3kUwO8VAJgKbW6dBsn3xl2vcAYKL
vPzySIdLkrCaYQ21ZZ51+udy5pmSeUMHyoIzKTIJJSNIuH8ZrknWtIlymj46YMCg
qfmsGuQxgXyuEHtTVMhuxOKVSy5WVt2gk/83FsJY3mhS0GW0o8yIIM2hUkS/hqfQ
eb2yW3kyZ8bciCzKRr88Pf3H1t6NwyMekOREJt0UMVQeWaHKjr/I/evCnH4ii6Cz
KfW3THwkxMFQeyMyJhmcBwA8MV0zgjkFQB5jnm5T+WwmmOd2Kg+gxgBc4YEnhNl7
PKzf1s8suh514D7D1UrKVPklJ2ZWQbmWT14wMEYF2uNcpQoW2ls52OhSGipcW/Z7
j8pVTT0qtA7w7kisXX8aHiEsvfZPuCGpEz6pcZKrm2xi3Seh49OivZX9oSKMebHQ
TMG8kQChm9+c3xSDPWghS1+9HxkPO2xAnmEMy0hlXriRoIhR+2VHZkwCEbdfGWx9
gu0hVIUYoLq+bsWzt06S0Utla+xvr0EKEhnoNGB4idiiXmO2qJHijnmibbgLXlIF
BH0f2WdNE0UmLrBEgV7qGRhNcWDQAfHXQR7lEpZs+CSpYVj6eNWNBCmwPxExEXVM
oVR55KxqCJ6ve+1Isfwy6Q8bLP6S17NUdMLa7QLil52fWlOjNrdFcguAxaXSQY1j
LID8dNauMYSeLOmOpHOH03Rws3355hqRpD9xD5V1s4RXDmukM2/umAwLZZKF8EGZ
ReWpSPlVQReWLriHLNu8PCjmi8PL79MJWCeFdJRTcDbK5eatS/yaid80CcI/3BxT
QE+vOWlL+qlj1LnRNgS+CoLhmEyT4rKKlIp6vTCBb98d/MPXLasieLkl5kTxEDMW
+ZFIXmlKyDwVZ4cLWa+xEnChacev+RJpPGHu6mJHSCdks3QO77ThfQFAGc296Iji
hUsBeWSODQ3bwsgiK9A0qqynYD1RjLPZfldhWf/9QTUDjrz8yBMhJn5opnR3oAtX
MJ6B41A/3+LkBnM1DazeF900ll+aBrL9xyHe2zu072T3BJvu5KcadU6NmQWXXXiG
ztw4ZqtfsNO4zl3yOn4xvVxrK7iLw2C034Fm6tCY4mCiWP954ZKRcdRyesICkqUy
ZZIPAv1DGltlM2tIZtSg2I3g0kwqJ7k1D/Y6k4U44DCxQgOn6EYQ5rb2S3UL5wLg
+BYB1UuppQoUyFU0JQRJk0sMRNiFI61pLpTJkQrVNRGcTDAg+K0tePeDUUI187hK
ceinizX9LoJkLh+dhoWocsvaR0wq7P9hBMPesXOeuzz2CoOEMJFlCsnrA/lm3ZBj
eMqOh0juATWnvI0zWMsbdPVYne3iEKDPbcL8wRUm0jBrnF2G76lt9mqhaKklwvoR
TaLyEGBw1I6qjwui/H9hJqmfVZZB8miFQXYWywUXDZyuLc5XUMPyy3G223Y5oUg9
uEv90lhz8p5Aaw7zP7FFct8BOzCbwLkQm9hniEjmUTs6itatRXxiBynmBhCthk7g
Z3Pr5+h3woFwGa7YFNG193lQI3aXxkbTP1ALcw7VY3+ue4hfEoN9EqgTc5AEKXNB
ZYwqX2X1JAuxfLW6aTjOu62c+W+jwPevDt7TghbcKP/Sihlo953+giJDOLEByR0F
sD+D2KNTwQDL6S+y5Ow/JLMKvmwDnYSkLom+8QU29RFfeaCulVD3aGnCUAPbpOi3
4cGNrpm5SmF2V6bnXl5Y1VlWvpR2T9tI/TGsUUkMYwqquyv0FU9hW7SDD7cTV/Lh
Xu2nuPbxjP7KhrAyRuiVSgn9DCHG11i/e3rGqABCUTryaQD/JpxojjpO+6bLhmUu
9mfchVNiUvLUaaBWV09zsF6VIfKcJYlLdEHbAXVYmLVxAIpg5l6pPQEcnLPUHVH5
WMSXKGZENFf0Tr4nqvba5sjKkl81lgsbCQ+lSwHFyrLpClhmoCPdWVyVJ6N1Jqbk
Bl//OXW97ahacXuc/pRxntIfSK5z8EQXgUOAXuwqs1gSXqcCeQavnUM2M9ClM53s
n7yimGYw6JuCqmHd1gzebdgd0s2IsJmWQgXJbScg61yvTPpZEEiYuKnbJ1DF1vYH
vtpUaZcHdgCTNyqfqKWYFKBezCZoW4hl3+Q7Z18JywxHSN94i5MCp5peeGQTr4QR
2hyjjICBq7EzBvC5pRRtzXJGB6J8eMfHsWkqsTrgwXDIBNY5h65I8qMJpek0FubW
9HAy4tkCPnXCg+1P8dgEQvL8/oYRMnyeTNv9axMd358P1iHuaBUOE+B5/ZFcQwRm
xsCf2lN/CPuACXCH5wY81tjdysZTRY3EopMrhikwlKqdtrgP6boEwvQ1h6jOjL1c
Lb4gDstFsTGCef3qeG5wS+vrxIhQzqmCEIZvmDTfErfJH1rFNpZhC6V8Mm1TXoBa
5utES91Wsip9903ASOQzsHIAcMuZXZAXNZoIc1e1AqQfgP0jLuaw8tiSrl3iJF63
emT8DzE1fPsyNyrBxVNr4Wf9o7AFYwh7LIPw/3ESYOBMuTPvr2Qi2PJfJ8aImVbd
IZxnu2kFTN/sg1fauSPC2E7GCqZs6FYTWDWRmPiK6P/nnJTcX8tk3yIOnr+D6OCx
vclNqdWCRy9SC+6a0JDwCKyWg5XgoXypby3+kgMfBSfYlU8bkF10QUVXMLGnFvNb
Pm1GjGScbv+K55eXX4Dgwa9ZkG/IUCTNolnoi6WT0oXrXMbChmPWEEx+RCXPa3Lj
rFtVhRbKeE6QZncbK3TqcHiXGIhFcLopITGMGH2ZdIBvwZPyOu0VQ7MVlMblIGOP
z0fNuoqXXx3p8CBeLej8c/lBGAAsMtsQg9A/+0Cv+X/3R4pnhhddouZu6mnbkHTm
MsJUKtNd14aWGIFm3OY+XVLihz+5XpFCqcUqGwxhoA+ZeefYEMj+ENkFwyhtP9Am
IpIm87U2mhsGT+iqT02Ct58IkkHLiCNSXEGppUpTZL0zQI48JHxbD4mwWSdLgjv7
sSAddit88dj71xCjzud79tg79Em1Q7cC/b33ulRjAaEAw3Z4mbAONp7+PynmRDha
mnLVt6jhBOIV//vRA4q38fs0mZHUZVMOQb6nMq2i90k4qAQjxK9Zw91KbI7G1pou
2PTzgffDC8LF6sL0BtwaAh9pSuz2TDEJ4WTHYg2rfjAY3541HpOa1gb7DON/H9sy
cVInH4Qlw9PH34D6nB1yf5whT2jhw7xGh6D12TUxxQpbVzd2Y1g71OULz53QoIov
qe6MWw2kIAKQ58X1k53/ycq9rBIY6WHRTDrOC10Ya6unKmmXtRfL7ceXnWsEqdMR
KwI8LS6VYYNJNprG6G0sCPuc9zf9cUhe9LPI0mv2Z1mEMT5p1j8lLJVBOdgRIp1+
Op9RvugWM8eCSwLv8y1KGk1OBQ9sFi1i+SQImUqcBsdvyGxU7bL9FK/FD5ay2P8N
BsX86zkSfZEEBX25/lXRmXeEC84QwS4RKeaOWdZjAuW8jtmtd/bFdCcvnzo6pABM
tr9becJ1vXRBoJSjVG3Klodk7ERpcXI7NF+uG1s2X5JnqD+Z97R83uuG1lUJC1G4
pVcmbTUMX1B4oE6cRS/hvQ+AZF1Yjg8l1dDyVBg0+DCndbPfysxm1mp3R8SsK3Ej
dniRtjZGa9UNpeppZa5VvUe9TSAUx1MMA1bLOw7n0968glsXf3sgWSD7xl5eY/xd
pR1qCKE0Pv0jManK+9Jn8z3b+dqrI9For1G6DJRS2VsVwujob0t3hfEwjipE43oe
xdVM6GY6rSH4eYliehCjz+UwXqM5d5x60MnfrnAtSDDMJW7jJdzH9dKK0EqQAg2X
KwAn3XDbuEN7AcqL1PHbzL88t/aEsOOLgGxO6fG/Xhb8A4RFkr6qj2VcAE0r+Zd3
dpbjdePMZwGKjzcaIrLRJ3kk17X1fIPkwk7fd8MjG0to9DebgxQ4/AMgE/RnRbr9
iKCgLtraxZrBOckGPhiIpf/InhZhJJMnnD1Ax0/qOM+MiCiou3+Xl5fLA9u+eUFl
8KMy/tfh+3zenQAXXid2upn2xxftbY+HthAdwFu53gbnmP2UiQpYvYI5aiGS3F9I
YXsRzMgoVpJ2OEPLii73MaW0aVu349IkpUbYPEfewR7KbUEFpIJh+PqynauDHdGU
tEE9MwQwIQPUw1u3+4/WN8MoewXSNbQn6UMotjozCxVvNCBEODOhJJPexsyQFMoD
OM2PaDtb3D/f4/bkLE2aAuhiR/ZDGqzCocgBQHYwgmj/UQ4yvwD8lAP/ifQ5/fkl
ZvbSoPNQCa7rXVEgqAC/sP88uZrUlJub0jPa0vbdUJaAY6A3hCOYOr2ICXz8sMgx
vc+4TK/c3Uz/Y1cu+SbGk3NETQ+oYuEvQFYTwbqkuIvHFJs7WQcseuQcIvgnaJ3f
zgxhVc+B07HdBlJBTudZXnLzSh6tuwqXBlPHUbgJblxGGS3t7bb1/cZtlndetJ9N
dNxdLVxm+hJWcYmpmwgEAjIMkWJDbwrhcAajVhjtOeW7TuNJUtEHvRov0F5JKTg7
zZMf61RAdoD+UH+rREruWEFRvYIJLeSoJs9SLJvaHT5+vWfQF4XdbZzXyrymO4E1
kagMlT2ebqOclZ49eoyCCYVKIUyZM7l+UgCIyjmnRCQHBILjotGc74Rq4XWs1dGh
LuoT2AFunnBFKZppSHgyACz5z0GanIY+lWAeZAxNu3hvCWtM9uR3Ykr5STE9ng4a
x9e1bhfbZBRBsE+J1VNg5lgXVBFWevhik1IdIsC6qQXxvWeRYHWpEyUBIpcZaXlP
ENS0BlzmwvmB1I9PrPQeHbP7lJ8cSqgolGvcAAp5PetS/XHQCr/CecKBeEpJJfrb
T7ofLokktJq8yqr8MWECoUY6Q7KOIKpPhEAUAXWER9vP1nDirexE1zkYtmzE/m/O
4hWuqcZHx9hZWxJ9UDl4fZMn84BFPy3peuGrgOuFeLjYY3N8hUl3vxZBp5Z7dHtl
CVi+IqTWVL7hrVQ0Lo/FAFhaIs1v1vdAYxT9u083KBSzY65Xa0AM71d+SWq35Y1X
X4/pZpj1mNUml2OgXVzvBFfn35Du2rZnTOj1s9RM2DHVF9jG+c0CSt2kfiWqmI3G
joKEpfMHBPQtTYgTWEpEaqwlKIRn8Nfhh6jqnRipDC+um45cytzHLDJgY+Gtj2BQ
GdD72+cqQVjtGBSkN0u/7rT3U3sq00EkgRQiK2QJB9mbZbWg/AOFg1Sflc4jUXO8
lXpG8eXGMJiN8SPx5bbJbsvFaOG/KjYZ/BKhbRrp48yHHRNCy8ed0bHrMrwKtiDg
Fqzdl7Lmo+Q9kh4yDf6m/G+Mx+mQi4G+usy3lwH34kFXi76Z2TQk0+hPO0GbFXgh
s9BRPdrGp2441QEfjRc0Q3oxsyp5BrS3UMRAaNbOG3Vj+486h0Gr3zRuDoCF/UeM
NchIXginKyi9/ACFJj6yvOgQIkJ+el9P5BHU5J+dPo6psQZahG9eC8/z7wVqwTKD
XtgZK3GXEXN7qr6zG8HTk+t+LxBuCBaNgXrqw6phphVyrwMaJQWAmx+1Nn2H6Plg
wVbPji/qdEBa1w0CMVlxtuYUbBjQjEmCemPkv+MSrwEfKXz38WBC6wjMt/dANZC+
oKSN1xzEaUZU8ZDHZcroDki9V6Ugax51x6OM+HvAkwetGoRq4ilO7Ns3/n3IEuzx
ToiSVPwR15LlHwJXZ9aR9SJHis9xWOlA4jI7moxqosRU20tJm7Nh+OVl/Qqv3zAn
sAqXHzjuHdvl2n+///g+dmxE/S9VjRqI6qaFxy9xh+nsST/XjhtmSAJjwfQxTxR2
AzrWhBKDX8cJMSX54mf/kCcaTSSNP1JCl3H/GfXq4RWiJ0bf+geueL5Kx7cmM1O/
j4A0QL2pA4xUri4BFKXB4hMKuSbXWT9HHljHhJ0Wb0qOQXSApDsjUKIx3b7/2SmR
uqzPAbt22W8enZEE2MA/55S1mrGm9IWOH+Hud4lUbOIQOjL6kfLHC2elweEcGFlB
ciJ341eofl/BZ3l15UWKmPxNpF9GUEpmngQ1Ou9eEW7CyVQ/t92wEQS91NHY0/1x
jY0/UemnHiHfvPJpEWSbWKdPZy8offH2EZU6ymXGlboBlvqzCzCAJUJVfDkHf2Ev
Bcuh3jjDNUZdj9c9RqJtmRA0YnJQhWUJA9Dsj8u8+n87oYOQ1dIIx03qQB+EVqgZ
wLiGIWGp1e07l0LGzsEzlTgFxSID3T4XvkOp/3oBP3lKPRNSHF3cC2HSGE4cSTlH
9wsJT/gqI2B73EXH4B2CtaiXay8ISXACAtnvX7/qNq8/9CJmEUzNBE1tUYYKs5w0
hor8/B+Vzq/xNJvGYHkfFld/PIT/wqo6jDj23AvqxqfgeZ6BPsPMP+9qPiGPjdzu
MpzcHMkiQ5fid9H8ST59Id7eSPkvgWxc1XIIlSFrTXYH16SSQj/yvh7WOEDbnzww
7xwzgT4QWVepyf01WJxwudSxCjveJl/cPM8GdVjkyiSYAXdcKCLcQgfVfbKQ0m4h
8WIeKoiQu0DVKeXyf7orwPnVAqeklkItxK+6Zx/iBXN92vAyIjJYoDICAwvBmxC7
6JdYnuPfZN3SUyy99L+wnd6PB2QOeHlVMR6q/RGSsLybfL/vj8c0Xai2oF0QkVGr
3efxIXqmqQbQSHfBqkUiyjwKqds8RuQufO+yKn2149zi2PoayhMK2CA2AbEhihrc
fUZjnauo/MIRPSO0yITjkeoRXlM/nTBbaH/ZL2hRaeEUwRsOpgLSRXFhCVX/TmQc
jsnzF4Leyuzar4Ym9oCiq02uFVVL9ZI9c8ic/5gBZjJG3HGm9+bvch5mV7CjuhJR
+SGtx6YxQ02L5/2/iF9PFvpTkjkirqKnv8nxtKEpvYAPPdnrh3e0Re32EdgAZuWF
gzU3/t7OTdlHhQ1AtFJdVdeolQRWC23u8VftTwpHA+c2ATpjVTm2WU8Vdc0uKZ3T
i0+rmGb3IVtahmgBYXBapyU5aPHFfzlM28QtIgWz2/ZG/ggnUuyObSMxJNJH3IwB
ZrFzIzApU/9vRZ94rxnOIcUDN2MMhrDT4BItJr8mi/f5YDlGvxhFMt7ujdD4uwtw
oLc1++gdcyPya+e02kDBgHeQxcLCUtjLMH+KNVFfONjSRjsOwHyHLe6A1/Ce2WW5
hEEQtdKFIiMnQuynlkM7pQigpXpkZl/iN9I/QUGQ760edWnnVmOrDu5N01xI+gD3
msYXP2RqWry/8T+cCS5XljsipFObYnnOrNaqeBpY+qbxykhwhU2nAwoAxEH3ZLnA
gj5MhvA2A3egDHyHZ6mmHoTj309GRxZ1XHVhJ9brg0NjhXHflRcpGqGqR+QzoxTN
bEmmqfV1nROy1VYpwz9vwHjniYu5bAsUStzvRDYCmncK0qkXXoNEpGoakVKRqJGG
/5Rb0lUtT2ESJp3O4vEtP4LmVALUhNQh0rjT89KZssHdeta0E/4VBNEMooQX+RBI
JUe4VzgXex3Gb1y9qtpHPHHirphgJi1KvnU1AhiLaS88IguWrT/AG/Atyp8MUdYe
AnomL7GNNb2PjrLoV5mkto2MBlbt8ls0TDjnHq+dYJeLisTjOPLbRsdVf0G1PtEA
ss1+GhtYa6h5/LedFXNZ7kxxPHm0uH0BxMX/b+bqdjfvJDnIgD8QEYfyVs8cwZY2
SbaQ/r/moS0nlMTDg82s4VCHueWEaSipV3tok4EDoYebPaIgGOjYHGd+Fct+RhlH
q8raALfxq2ifLu7OhfGYp3B23Sy5abQdVphy9d/OPUxF2knAsxS53mMev3wNsFbP
zwQqtF6G/ZNTyc4hYSocU1xvTM4u8DaTG4SwUL5+yP1sWviHCGqpv4SDYJityw+G
R6sVBePtxsj8O9Det4uWpSufxiAPfDJrocRuQHseUVwc25giWAe2uVkmayrJsLh2
3b7hkPHA796qQ66T0sy5Iztfy3DLQ0ByMVts+1JfHMfQyogtHhNPjHjq1kO9kudX
jwSqME2wUGcZS2+sFpTBM6lKWesxadtS06j9kI3ZjbYXNr6LhBm50yuHt36o6fOp
F8OrI8CQy5dzlOn42oMZhKh5UtT/+RVo0RJAsS4IIsb+azrXnUC6F1u7IClib81S
5ocQWhc3HgqMv5EmZiQ2CbNGKKTRzXDZAeI/m39L1l/HWk7bwfVm9bxMyqld9mDg
Bw1Es7Z2a7k0gLTYDbiBj/QJh2mz+GsTkrsS5PRujaAHo/r3OJKIvAcMvWK9dR/S
hHZ7bavIa1YvtHL8jMpjdt54+8ZUiEAzqkqnIcCwljAqxCNzU0NYk/C4OjATkt5K
gRMCcXQW2ET0FT6ldxUQ2DefnsUOTM24NuNSgo25j4tb86hK6ZlnhLxOtx8KFKnY
r9nQ0jF6+5iRoO56oLt/3V5EklmR6S/cH0XHPp/7UQCCkuhJXeemfrOWrRUJiq1M
hZZp1DMPTVIvq0FmqrcXmDoFKAoHUAw3uzesr129a+xKQLVGPdw5bODy/zfIXCIg
KwlI64DxnBT8iUew7l+0x9zyM7dkfnKCHYBvFcyVN5906vB/gAC6/DpZ/6ilRY1o
sbuB+kjK8WJTBLanNPEZMOgsTNQyKZBk/TTa2/4Gk5Ot1gTvFMA2eg24ChTZdmOx
aqlH0NHE4RjPoIiTmqM1GeWOY+haKrAT/3GqDLaylsTXsiBwr17ZWiI5CRZp5d1M
WHw3qgK1gh8Scdcj/5KZoZ9eVZLde3onpat5KZCOj0GTEyRtfS99yGDTdstjfYon
AfZ+T37QxcDjBevR6MHBw6cOelIEjwYwXae12PYqMdXqnxQ1sC+GrSUOg2ja0w7V
Xh4yalnDBBRfGzj7SfTqBKJqBvAJ8AA6bFA61t6r8ETW/komK9hZPAu5nZKEEbr3
BJTRefz5YPg09oWqrWhsG2f9RPuwtcYohfy21V8N28R2KH6vheXNDQ4MxCRwYsux
Glvy7BYHziGSSDpQgpmCNeM/pt9GZu0YHmhcDbhpOnwuFKlAcE+NDknvgqntCFJD
/tdVa0a4A1J7Rt8ehPSaNphXuaiT6vvbf1Smr9iV510jTu8f+gxbTmRGPn8ZS/Zb
dNXphMzKbsup/QLlpscRv7C+gw/8A4Oz0SxcqwFBKMHp3ouUIDUwOUjUxL5qWlI2
NCTCsA9WXU2qQ93C8U2CBwlFUo4qF1MOFlVVFS0KvgqvzPvwcpKAOX0dOFpgwrVb
XJewqwrc1L0XkI22rZ8UtpPmgjvsmNX3n/Q5LspDhA+6mMonN+toUqK7knFbuCFp
TJJi1gVfmxfVn/+WD0S7UIqZ4plTUHJ+8s+jlgXoP/mn7ihEqCLdkh5V1fUkZUk+
Rtie2AiN8YWZKi6JMbaP5aGzgw4IoNM3ObOLdVEqXQuYQHO5BNHAFrbvkddxzv7i
F/+1Mm+wt0f6lwfkkKqQNAyA1e0tIlBsaxuyGM6o6XK20TJh1iLtZy6xXhVeXRXF
x7UfFHDgZ+X6m7aVy3n5Amky5QrD2IZ39R1++dylo8TJLLkVqOIIlzthHEGaMh/c
vzTUirza4YxVA8tcvSmo7d8b/IpIFvaaK9YILFGzrhGHwA5wReHv0HX6Ajguvsuy
p513UySMiPuJ/eB4Uuo7IuV1/mtxW1sAYabCKXF/+RoMIBbo4JtDNn8Z7aB05GYe
6RDpjgUR2GBAH/o/6pCk1m+mVdE3iwAUw+Sj71dGc7LtJPO6sL9aIzFtQHb5io51
vYqU285pt9yPEX7Ht1SucZ/9gZxMgiaXYOcg4SmRxgkF7kqeO2Um0eowbR6nosWI
23gxhdTbqh/h2rhvBdg7mgiH4RWO4EpsWvNNXwTWlfnbOLfAh1cRoe+kBeRBpOOW
4bGjUiQzl2q+dYfOrPBdOM93vQQL8J6OtXEGVhEwJCZg8v4DeObN0KvGRJu8ulrw
li8/mVZv73t68WWfsQKB0MSM6cX/vlHqdFc6LuVkl0yLeXgiS0+n9m8W7DCCkFwu
jJKns7meZ+gCK9y9wfxKFA8xtSPxS4Mfs9dYV9v97SBi7l/idMzn0WznGpMJwsMS
27D0vOUtJ4w++Oaa748m+zFWOT3D4IuV8iRDsoKhXaxkANhbdzorpHu4nj26A7IC
usfUYlA2PScbexoe+DKK5EZ4zS6hzpVgAqGSy4m7U6RdGlej5itpDeJoNq5E0EIg
LcnojB0ahzAa5nhYgTDUZEomFNt4lALr2cEsZX8hqDFftaWlSCR77FtGhnlNtHrz
LlZUloWY4OmBmjKnsPxkv1kHiBgAbwzPkuRmT4TkNX+ttt/WZE4p5osdRSRx4+PO
OHHTz7JtR7mtAC4vB6T/Yh/D+FU1OWXOMYNIWJtUciJbWGETNNOC+VGIxtt/d41q
vHHU3Pi7jUJodDsou5A8nNK/qpnVwVZfRVqeH+Y8pz97jCEp953umGXwBob8a2Pq
SStA5kuW0pTr7+FZO8Szo63/HsQEOF7mX07rzz2uAz9aIE/hZHiTHlPQKHJkoSY0
wQnYbj6GiYahoQQZ26jxPVGDXzq5b6lHgJ96L8darzjvROt0XUDbuFHVYThBoVdk
u8MP+M2lj0zq5TlrJ4tLt1hA5JZMUNfaboH7u9gpRuMK0NUZgHrf2BLuq4V7lMnV
/QGlyQB22iN8f6Yuh7ZfGoErl13UsfqLiEKKtGgCH8139qSw2yrTxy+8cT9lHtyA
DgMxYqUAg3l68QBnWF8QbFIEWdTfN0Gv7b5R7kjIxyxfl1dPKfB8cTp9jMy7Vu+4
oPC8gIu+Ft+oA+W0lJgONFV2+X7y8qWk0qXYONMeIBxQO2r11Aey1yddgmERKVNa
RR3GZuBlsHfQVfjnnSOX49FZ2F7ASqVj/h8k4BhcvL2FDj9vWwELvCRf6sfDmks6
Jp710skMt0+jAI8Lp6SaeVt/FrA2iEtYWJX6i07DiNfuUdU6oAFhsNI20tTxryHd
LaToagZAfN1+jZrqCxeXubSIpnBN7+R1dmCr+YHVOZ6NxjI3Jsqbjir9l0pT9sNi
pdGawfEF2OoW/9/u/iZ0QK/5CTXIZFPsEv6d/Sz6ZG2lad+qj7mY8vf5n1XsiAXH
VbVmO2f6Ae/dVERlu+OG7aGhkF2xNkE5lsJVJDIuGBK/V2rdzObtguw5MovVGNJJ
gq3mYD8s6cUy4y4eAPw8AxTIXH9RGWSs92x7N5kXewrV76dsEz8W0CQP4ToJQVSO
OySvDKDBTxpoRkCao9rFILtt5JuU1ju7UMPWvfBJqgBGhsebtZ18zYFdJ/iYGAkN
+yQTGAVEWve0DU/8pE8SJEY6gX9Avj5+8fWC2wE+e9NgVJ8sx0NgF/qhbERjJg1p
H90k4IlAfa7yqII+xPGSBpL784BlVV9dNYPg+ZqbJA6r3iPH1Ovk/jFY5YzFEPF5
yuuS/S56/zwfIml2HSo9CkYfnGEijgZpzVRqoVB1dwh1V4esb5S12nv+iHB7X99Y
LbXQgEcS0/eE2OFmwxLIT9SnwDc15wuaaDPo6MWy68CWGA90g5sz1mJP2aryEt1V
BJPr8l1VcDCtjkHSt4bVfLyFR7cNGUZTsfKvTLmOxK5svZhmYsRMS+Npt44Ed25o
4IPQNQlXJ3YRTwxsUWH2wWl5OadKLoY/eRtIKKCv4elMkcIbQwXZa920t2WSg1vH
HPonZ4vpbks9xN9LyMUtreH2pTFB+xND+r0GNHvMNUAkEV8H7wNc6WkBf4uZZ2Tc
Fb56i755xjB7bOiNWoZHRcn6ScVlVcI36J9xLW1jLYej8jsMi9PaStCjpZ5uZT0d
Ltjo++ZKyRgsM0ubHH5phF4fIKOKRQy2DXDq8nySeXf+P8oXD5ynFPTiCvzIUSS7
9PwlixWV98oueuhTE/iaU0pMWfA8xbn26iEf2vSn5ZYKmOSLvASMi29ocT7SnPnH
V6ryT/uVP4+PODt9g5QVRu9z0XLv2KwXk8rrUQ1uof6BBQm9PCmv9frG9Wns72pw
LYeIyxaccCsuSMMwMiKm/2zBcm6wApk2WFeOE3tHdON58Fd69JDXEEMJqF/aZfA7
GYS6jNQ6ALKXtAnpfSMOg5pahsbOqCvcWCMSRBuy+bFYAhWRe1wiN91Sv5kkrcxJ
oRyN/FHmU0EF6ImVYc0sr5Fke0sEfYsGdT2F4WwvvaG7ZFh9Kn0Vp3UcpI12egbQ
44Kd+O4fr5AlFUh3c75HpR2tQ76isYrkyIaqlL3Ntd7wVRhxv5mJHlL0dsu8Z8J6
G489vmRP3yTVvLdMti46WrH21kFWNwaqL6Jg8VR6Ia1k1kKqRnlh/xEDEarqlnO7
pgmfJaREgnTv+gBue5dICyNqfRE6C/pTRaiQIee2xVyjap3UXJW63C7eH0c2F6yE
razovztQ8pJh7X5XQ13nrVfrZkQo/H5Z3PMx/FdEGBZkogv7zCjgs/il2fB+0AC9
rehDeLx0DkoWSnxtQXn80J7C8Ij4I/yRU7kB6HNEScjCnqZzhcW5My68knt7DoU9
c45k7E/PnPI7YM0tbfQ6jAYsL7LzCYTxUdHHhI9WasE333MXb/m+H6c/z/yUnZLO
Fo6P+SpGnDgKD+HSJNWbTx1Wz814tXVtFOrSbDl2HB+uC83xqyAsSBr11a/JxQoc
H0OaTU8uSV60jg9OArLeoUAdeQ5J194FNN9WVVtjhoXfxMyghf5Y4CXeDaaeGu8y
TQ8g73N/LfXSlBRvN7zxKU0pLcW0MGJoGLfb5dws6vUWop0tnfNHEs2LBJgZudF5
LIvSSVKJ3DR8nWvlUkdYguvGt73Q+RyrHkvv88iF7iCWUHOZJRDPOhV74kz941Yq
Br5L36U331dQQ6aUG6y1Zj2n6zoR9t1TskeT429G5od44E5LL329Gwcl6D46XisH
gXuu8lfKGl6Yn+kMIkBhKGEjTiMSVBFV+HHUUDukiQjlENB9bUidveDvU40ocd0r
o/JXIS2OZb2Gp72VH4jjWmZ/Rvx5ulXdEywuvsNr9fJ40fiSk5VVPGMZEqA0TWFL
txOFjF6jbPEL2p693TddFiMLXAagF1PcTSWN7oZ9oejE2C4Kh6tkiyUI2CfdhJ0k
a59ZC+H4/zjNy/Ezs4d6VPewhBIG0e5iWUW9DI+jMNgV5ACpmTKXqpcjrbm5eNAE
Glg7sEMvD+hinbv0TANlllfKCwt8P+393XnEDTI/0OMg9/1kEtNj/OIvSTOLSKzS
iIkH4juZp7JO/R3GAKu/yJi8BDxYHlvM517E+s2k9dqtsS7naBfc7m17LHMrLAqy
zGgbp0uzYAeCGORWHpIKcufdw9DtrrQU3ZBNOohc5CCo6qIJTF6Gn9fa+JEgITF9
HrWJCkBh25VGmQjGyVAj9a1wcDfZFjuYrCnR9pLlHSUurUkbF8lSsfoOY1v+H9qX
n2Iczogzzs3cGIgitVHTOfhvzSjfq8LhonCQuaB8izp671mK+s1lcjMt/kWf7WCN
xu2Cr2owGji7EMOaJrlPmvxHBegCNMOfCfn3/sJW98K/GstDhAzCn17K5Z8y4ovw
savEt1PeEPuAZtw9H48YSgA7Ip+yPcOr5ErAPOzUcBGFsX3qxPRkDmV+7cr7EQjP
JQ0QJTGCeJrrDxlqW4ckxbyfiDx7K7m5zMX1UVjm9Am5qRlH/MdslXdlIYTL3H3w
//VYZw1tqgfAEcW3m6jHI/sL0YCpjVHut7Gd3tbTpqMeiD3Yd/utdT0vA14bfWwJ
aigq+7dC7gMr1XTOfYE4Fhyre6zhoXwmCakP52LxAhRt9aifsBZfD3rE/LJYURky
+ykLqqMAxv4R+uzEjhZi5W7Xn/vUcCHb5Ts9nhERdc0RA++jMtU7t3j+dmSAkgjI
HxyaAf7uGmOicQhxp6UzMgzAdmgY+1nd9D/6MlKGdKhSmRS1kiDEH9tyaovzgB6p
eEJl4MrMOCIdAxlcVLz2Wa3MBoi8NrrnwlAKeYycPOV/RlHrlEdsrawCWL0g6s4V
Q1JAO3cl1HVGDvyuM6Cr+wYfulBirQr0uUQ66zcpi/pKgXShlgiJ7tVUoyvwoFXO
ssZ0/6FBRqJT21C2Y6hyvBioSSdol70ccIboBQR1mYrQyrPm9qJIz0HzmNrSPNLX
9zOVACYTUTqoOge52zwJ4IV9w5zI6O7nDMcUKcYrhZBQOZBtFs7C225VpfO+Q8GZ
3trnKBFykGGyCFUoTSRwg0MCpA+E228BmtJHSxzbiAKDitE/pfbVUMEnI252QkGJ
1/VCraBixeI2BP0qtzjLQaNuesSsAYTdrnGEo67Wz/FSWb8nHWp5U60BIIfrh3VM
PP6LW/Y7jtlEBSdMyblLDrvam5H5pB12FtSSY7QyM5QWNcUnFs4Hbw9WOdMPWoz8
zKCBIPRyv9QJVhjtr2hHjB+zYNF56LyIMX3pbpM7PGnSXRMGJW1Nx1scgDVdMEGp
G/zYOIPe/ZGtlGqhhtRtXwEO2sybYa4kuPyeFndGWEzWWcG6qUvh5bOmOLmaIaMS
zPBhP+IukibnNPyhY2JmqJbwn/DhqNDPt6oG9t84BE/Ij58HaBydWIGmaU3YQ1vE
9pHq8e3cNA/lBNgMf6ME7y/91wir0PStBGMofMzg1HIeGS62SVWWGaD95PXWOvfY
Q+WLXgsSbPehe1sdABI6+/JZv/7+lGkv9oT41rbkeFsRYg3lWumauxP2tekn/ux1
EVZEtlvl0mH+Omwv7Z0YsOFxKXBAg3VyA5dfryg33SdPpY/qMugz2KmtGnm/0nFc
xUSDM/MBBobZfeS+LT0wTTxxLsWYr7AKzNzR5uaL2AWZyajmq1FOnMZM61zF0wb4
JuwcNzlqucFLmCIhoyZ6tQFTFS390p5sacgAc6gTDxTKmsXpUY0nFxFzZkhZBFZp
iV9LieK8YRThzv2h9en60J4QQYb+iyoga3I9lVnqQTtWxJzv4B3004zFiDfcKPMt
PICg2sjkR9d4Vshh/nG16JLX2vnIk+AMPGM25eE7w+0L/aXWciCl/sfA+BxjGtc8
xBy4RipfGBDWTYtM7F13KYxOJRo01nXmhsToBKiSIh3zOhn7/Cnsx+UOQFNs+yIu
MELBs1dDrf3v6QGxeG8jPTUvcJ12YnPyrUp95RPc8nDYRREJpH2UW5gR5PLqHDzk
7v/pWdaSXOdbvldQSUUH2RfByQMbH+kpYXnu3hIRXlZn8cBAoBevtr636zqT7Nl3
/eUMui+j2VJjPSfc5lOquhcWUY1KW5Ia+qRtM6w79PWkb8BjtOx17t6j6OSFpvlb
JlS0pJlH+rdz4TftwFbWl7v9UK8/krNlmXXp5Qe2XBYMMRdEkxeF1TQWaMUBE/3G
3IEVVqptD3cxhVE09zj9Yo0UIa64RTy/i0ewElHoccPtNNt8jQLZ19nCkyiygFja
RHnsVK8EyHIcdsH6MnI89faxM4VQ1sTqXBSw5+7xwBxlgFH5sytMj3INYypCILcn
snFlcO99FCknWGK2F1JddwEzMQb3C3xskxhcSOq9J+frIRcJSTO3MKQkQkp//e8v
vSlZL4hD9PCZqWyFNPTBBK1zIB5b3l39V/xviDSWCkAyrZi/56g/R1XH35MGXGK8
ax5IZkVw3XKkAw6gJWJ8RSNnmgjNHEvVTU8B1tRM66wDWIoyxtklt23MCeN4rX/B
aGne5Kw+/hJsscQShO9reWboBdOGmBS/RT3+ziZW+o1SJxvzwuxJSPoezkaetx25
BrGxTfJFE4oAn7An4Ajrm8kXHOBiQxdY/sD8BT+GZYKVXsb5z/Arpl6LvhilGRkR
UnZrTU3phbM8D7GWt99Bn0RNYsSbb4MSeFbCr+maF3jSPjJ9LjgucIBUQ3gSKqjq
pmUFiEELRl39IuL48tkRszRcghPFdfMFSy1VebF9KQY9b+p+H6zQvF3ask8nx2aO
w1cy8WScbpR567RbYFlu/LKEzkET80aF64h4Cf08DpY+u4HuiHkOFzxZXE14HLiy
LXAl5iaqKFZIWI/G1QLSgvj62t83FqXi2eCU1UqSQyfpYsYqWgvAOpyax+3dPavN
oX8eqYLCb7dqRYA9uDFKEXTGnIJbvxOyOGgx6LQVT73artCjdQFISbmkTuoppICB
PWl6Tzv3toTYrq9+xlUnkYtjafZG32h2Cw+pPwpYpkW43Kv1sRwXBSYQVXoCLNyZ
ZuKXyaXLkx+BPTG0vvZvWQKs98S/t4d3i2CQ8JrE4AuR3jZgP3T1IUm5FofAyedX
DPcI3hR5+9/lr4L2J/Y37KLD64UiBssaElVSC33ef6UwxHts2JB5aMEA9MhXR+7Z
Ry9X3r4Lh92lZwVfnURB/fkLGMnJM+T6STqDA1DCbnf1t9wEpnORgxD+c9mKnXqI
KfG1zPAt3Y0sMD0P/O0oom+ci+SGPF7ojQuvrIUc4iK74Yrr1QFYvtnN5P4cyGz0
0IQVZ9P9PGGgahBc+rSrJahKx/RbkmWK5kmif1QO3UL+qUnWZVoeapUeG4Ur9Ipo
JLFS0D9vGrzVJNmgT6P4uJmZ0ZdYJ3tr9UJvy9u5F0EW6ltCO0t8kp16yWp/93X6
jdw8f+5imh/w9pr26kiZi5OWbYk5OEovgslo435ce6huIDAi4C4nCqQXI7Tz3LIg
yXMIruhrrH+PyRiIK9M5hFR/eKqaiBbwE5KMAo2AJv81Q0baGDqLznro1mvy3pHO
LKusmGcPJ/10H9KcqIPcQGw6sAEjJWaEzBF5ssyU6HRaK2K0KKN5RwPzUHKOhQfI
oREjzbfWGsrYuh55ymRmLNEwVAEn8yi4LMyqN6jOszqiThk0sDmR1G1QLHmkNE/m
0QfNDqsusqahfQwyjucDctcFxWiPHWWpouY0o3EIgl2KGehatj86ie3YTDV+Decc
LPEDzWgYZhF/A2t1NU5HiVeCUSqJFGKEtGm79bgfIcRy2KdW+ovXoDQIsEkXXF+K
UBeQtBD6DoaJgdh++4hrgEew8t6mP3YopyiS8RtFcfxwXWyGgMPLiFiOFDqFv3vp
GPUaN/elTHBwEvpwnkiGgPdxqRUdbW2078INWRDfJ6rVMknz29SvBzj0NOzImdJX
pGy5x7efz23oYZQBcjKEdF/m/MmCP49SF8ENuGjDZuhLL8YvJRU4zq9/tWqEywmy
xj6ZQfn/YNHZcweUy578NI8fZFOBLZw3B5eAEn05wHjWsmXegOO1BYJoIiu0IoVS
LxpcesMX3D1G92iIfp4MZlKVsGYljY03qw4b0caCoqeyu9JLb2e2hsj05UsceoK2
AaIhiy1NOQBr5tmYX9/RPBS2jkGafvQywYz/Q5yE9v2Z3AXryMsvX6J9bn38R/SO
l4wNGCvnH4eRmpp/aoxONc0DDOTQuqZmnazpg0+R7lwqekou8IzfzNLRXxr3dQUN
cdcZJsbgwuUUZtptvIPAX5jZUVxtzlD11nda2zmdvEtpzYwrrnd3pUoemJAQ3eDs
aR9AdBHtwYZdjv/bvgfjkmQSADlTKmPCVAUCwAvxQlMZLurkbr5mGHQPh9xuBV4S
Qd1GH7yCm7vGT/7bOHgm8toNR9MvFr8D16aoG3jKGW/vzZ3f4hNokBB2teU9MIcp
Ltfz30p5At/f8KP9ofJnQdRMt1iDqDrgwiGW6mZfBqWCz34Vh+VXnB1qstbefh99
+YqDZsaH4XS03CRyfgxcr2anG6HnCGBTIiSstPc+yy49pu5zKhY2VLu7xCwbbYs1
eewTrEXR/gCL3by+oJmmtzuIzfMKxOpxElrQ7dzxD9Z7vvgHCxcjfuT/zwaE2ZsQ
SWryYa+Dt5JfiClGnjN7kX2gNT2sIOXPdZsksWfHFLTAePNF18gftYcJJWlDP7fr
T2norWNNAIjhOJc1ipdA0eV4xMjM1Rc+fYb1ZdP3o1At1aDJ2Fu+Qclxui//aUpN
3/72BdgLUSPXXFB5Vgl0NYy7GPITnfdT2Rn9hIM5Z0w1lGRGguKcyDr9/fF587tE
Y8dMFooGVZzopn7RCkS64pPynupzV9zyJPhVrOxg1wRG0MyPjVc6jc3Fiz4Xopqj
9v/S8EnJDG/F19P9Rm9xZMQb4/XnLCpGbk5/Kcx8A/9EiC8Am3Lg7m8LYzj2bW1Q
dgd9hbmEOGdlWhEnDN1GtuBVeHo5wa/kwZFUGijl9BnavHkf2NMb4FPL9Q+OV94m
t5IbBUU1+RMgx45rLJruJuvUgzcQ2VUiWiCe386AViugx9oMSpynFG+17Lbb/qa7
CtcpHaBJUk0lu1Zxz8az0L70N/FMzNydLw5oWOGUiyhOwiTTA+M84FCPorE1Hn8s
ASbcE0JOvwu+r2rimRBPmgw/PChoAgmQLD1+q31IM/K+aajC4uM8rSA8/EGyN2bf
t42Q18LMoB0LYzjIq8rQRDlmxcBe56IaGyty3rvMvGgC/81Fr9JYtV9SKAyPRgOv
7pL/JK1oG0fhBZ593t73aMSy+mnUTird8ZsNTR+1T3NBXORg76J8ZmJ25FkRUfy0
UzDEwq6XlMd258i+bD51EaK1b0bv4zAciGePEvS3hQtLOJdvx4wzW1wNjonDypJQ
Fbqa98+rGGRiIr8Tsg6rqfQ6ZMB9YyKRysKEYtYCQkP6peTXb+7HsfGwri0ruqJP
J/qdd7gix4vsqzT6fOcALhvWHHwHqej62lYfmMbQvlbpx9v4Jy+bIcBUUlNqR32x
cWKYOEPcOeTVKeKkTsTZQih1neAu9ydHkvuyu+Fo2fMHScm4Az1kXpkIsbCJ8YzU
+XDIl/DC8nGFcYPCCmupOkGVjf59aJGmmu7X7sSjyJzX7w2vDiCBIkcPwO/Dvg5K
bTx9SadKkk3WfB1IYU5qUnrCpTV06iDevZivARQ8lRA8jEguBV2LinsKhk9vcbE7
5eUG05P7b8jZCa1fdx5VmUam4ZimtEkmK94UpyE9GgYgs1ADmVHHAgZG3vpsXQtd
vPsTvumVO2yTbdQR7EyBH4D9kw9AD2AvZ9AsZsLtFDafWQ01x6E6Z8NscxxQGLbU
qRi/ZEtKUzeyz/KKdhrER/7F2qN0VdD1zwH3E2HKe1smuunHv4XkZ5ioIbVEgLoW
rhcrnqWrovQg7ZGvQTB5FqHDQeBe4SlGrpCvfJtEk/EKQL8CfJwxD4MjIinF+0Sa
D3wP5sY4Hvdz9Jw4/NejHEYMJ5Y81FEODYL+E2qnKdm9V0BIgKbDMNcYthXnfMCA
VtzFtXj2SkS0HPLmibugp0zrRcVCH2HmOysCrnLTt2DcuHiflFWIL2qz3vwxsFMR
TWMX+lEuiNRevodECvXNncaXHHEmnYnC7jtmMshrGZ490YoNm2VI19vhIM6adPCM
lddzHLImxiAjF1OfSibmHfZ7/0giCU/4M5rtvJyv0aGf1RDBTG/wlTioU2kSslrT
pJPVqIqXSK7vRUtumzYEMcZNeSv8F2CA1/+7Gzin/tH423LRVF9GBQvNZ+mj/Jmg
rbfb6pcvtT0Rhbje5O5o0a7PBM/XnCUDfH8+Zf/czhZeKyf87G8GO31ujX4JBcO6
p/05ncFVYQ6t6QPy5J9Uwc6C8nE994owxdUAb3Im8oaUo4E8rujnqKUOCAD1m/4N
pSVoratj3EL7m3AGRh8n8S0IEJRNt3U62ZEXlH/Y909cU19UjAJfnMjvqRua6DzH
wkjajhmLJ4Lf8AziGKfjYZqtGnVQS31lClSP+f/QGk0dfzVxEGtKf0Rudfa5WPiw
0ly/4NCwAmKjgqfC9hIWD8OPfvx5dMAPb0Hg7vqjzSLCSsb7efNcCm9mrUOhK/ZY
KfLCOeJRMSnk0/1z7AOap+2KZMO38qhGyhqIZ/QloFdjBnA8vtlPmeZMwOtIZe7W
2sPc5rpodqWp5NUjQegN3gKOFiAOtTCBX+kbU49EZc1TaX63bwOHTNnIolaa39xm
I6eSPyOX7vgxzc68iE/2wDYHoWr5GNdlPsBgu+4tXpheTwYo0aotTcShptwYwTIf
B+QciAf6VzA0w1im35I4MY/GN2E9GEAuvRZZ1qYjPa+MED4bbB25woaz82HnSFZg
TFWLY3XdpJ/QMg3WgzwWyHUF+ZyOjc83gu2hQeCTm94qfv84lqQmft9JrCyGjO5f
81HtB+KUvr9FUkYTPLSwg/R74VaPgTJZOy8LDtOhhsrIlZRaEpMQp898Dn8+NXhZ
5JUk7ab4AJrRdPiwiw5BFr0mZByszzimmz46CoEicv1QKjftdbsgPMke9r3AFz4K
N0h2Mb4z5ejqDa1n3Ds4s34fp/JIKX0UGBeWF9t5w/rbz+h8H1K0Kmf0EfZqKzRM
kAJXpWnXCd37+WxGLvQUq6Vt8Y++lnEaUCjq0lhI6VKE6UEeTPN4mzo5mNVNhaZH
AyOhE0eh/MLa/Y+gjoZxWcl7uRAHugHIuHA7ffOuHeOPI9JOlDwxZ32q1ZfJonfH
/FCnKJ825AC7sc5cxFaJO9vN0qQpSYGCK/KVxnGCeAAPDf0regupi7URDmiFWW5i
iqSWg3bqDVtqjQPLUxr2ypf7nl/lxcUX96ywrROYK5//Ke5T3Zi+JAXZqhY/fOsq
EG0auKNUveCLx+lY/R62l6hz7FH+xkeUQqFey3XZi9janjJkTdui3QnOGI1F11Il
pk9Px97bvw5TkviAHM6KhzhBDmp/vQd3ycN8ft1HYXVg2wB7bZ4drJJ0HbcyU4rk
LiAVr8L1zZ6v6mkcqAVFaLJEJBw4L8u2miBuMsVU0vQgN6Yyo1mwDCqSgYXefqch
s6plWBTsaeDFw2fJy2CwIqMRd1BBFZzh5jAMz2467JJfZpo2oFNDCR1qIxobWeco
ZtnvFAjDc/O50mlEid8LFKNCWoyQb8BYg9QEoR1izbHPIW12Y9N/GlXhScxYg5TV
EyZT0mpXpr9y6M7oE9swF2I2h4tOuUDvY7ghm8z91Rak4GQsBtEfpKV38fLdoZvJ
3kYBxZyJa0gRZDxMghdpJsvoaTBBQZdfquSvHM+YhRQHNfDYDHKpPdcAtGBbVrx9
IXN0BDl/hR0ndCIr+MqzB4ocxqQvt2PkNsT8PoJxXLVGEU3c+iOMTMuPdjJMX13C
24Sqq6V81ssIt29WjgOs1dPlxQTN5QThJtZ3tjn0Z+dFbpYyn0QkXAELQHrZiRnl
awFd4hyH75siaD0jsZFdgE0/P7kVqqjc12Eac9Wc+plZ0vuM47mTLK0sZ//XgSOy
NCiuxeUDPULe/SiEXDtEJUmvFp+GW/jnodgrkeVUUIjPvnbpKZYBZGdYMgB6p4cD
amHojO4R+AW7emrzk5GbVY9DtGAVtrIUiariaoiJD/qa+sFCVZXJ+JxYop+s4p9F
/QumrrIzFA6NBA2ww197mUX+BfyXHjQHnWj+HU9nA7pxeKx8HEjci5GSq+XjtFYh
9b4qgr0xZNpt4T0FVH9khN8SWCdERnkIHyAsQh3YEjBe4N4sbtFgN/c4yeRANFxU
a9BAY/5Rwp7/VDRMd64LwReIE9uVdpzzMtQ2onJIBH/CGGevzppGGDXJ/52RVmHD
x03luOjG3Nd+RHAX8n07elQn1KhUa4aqIwpZ75dA72cvRIDTrsQMADiNE46nM6cI
IwJqnuj36W8SMI6Yt3hnKnTcBc7/qQhad9lVqjA5hzDn4k9R770HvySbLRi9P2Oc
yNbubMFG3U4FK+cViSvcPEbUaVGTz6IDspphBfgRoX2UP4rSos1QVRZearLYjyfH
Y0k3Oyu40NsQT7UuqS+/vb6XVbIPf35p8RbkKFSgiYicapqLh2/QtzcguuiP+ajt
3fwlZjeLJTnaRlozeOYqxWlMryMmR1xqm9bpvm/xK3IIdxG1q6b5LwaJdnV/AmW9
a8aPwOc0r9azQOwuzvzwIDK272qQHRj2OQAV7ph+DHZ7+7NDRcMlq22MeOih0Q/s
Ef9uPnwMUCRo/U6hk4Ly9578CRKkk9IreCSxCUF0FShtdxjaNW32tKm3Ob2tKIjl
0yAr4i5Txmn57nyD3twmr+YqtYYhNoTMsQVhmxLcoj0g0+sksOoGoneC8kZMt2EK
ivDWbyDtJt/q7hK2JIgGGp0NqeS0zMbUG0E0GwsP6GQDMRnnsVFVFhMF/8vG8z8R
of2B5rf4eyykH1JrBufrmGlZOsfeSbedDUCJxlxO2OIIGV6aM28IsTYeNfrdQsr5
SzVGgCv2qGr50sY4Ff/CeIS2UgjlPbzS9t2lVyZCjmWGbsbsx6A7O3tV9305WWxH
kTRnUhl+nrZVh74+yQOkhuFM7xQuB2njxPdEa7XW+w9YZutUMCZgdkFNuHa3V4dY
MlGukYq1q1+pgP/+KrOuiGoLqJ0F+8nQhIOufGroavDC/kO+gFxEa1tKnQbd2bqw
mzzcUJZ9yw+w7kYXphINmPwfCEDOz8yIqDAbIZw24uaJQf7hyI7syOwZEO5KbQ8K
GGa4DB16qMGrf0i1zcNOqXhnpMpqVtSMJELMQYNDYAz6Zie7fImUMpe7N8FFDkAX
CsoAX+EtQQ/PT5M916xHoVIRmjLXS6LI+ovISP9kcYI4MmPhkxRtbR5en8kGwaV9
oW9W2UzbFKqzwBAijHhV5dEBxH2rQk6v9hcEg+O+81IWaUTA6hymMPq8hwZRHio+
uNKK8RXp8S7+rBZxgyPYxcRd0W6K8pDJXbK2PLsUhGtNhP1WB/VWs6e6Gi6PKv9D
ncEf3UA423LdavhsT9enxve6fFCqpWnHheyn2XrANtMW5JxK5NJTTMWWNNaa7cJi
eMLIZ/LWv8VeOlvV3OCbh1Cs1XyBcBHnPcxW8CDkCiopkKTWuRQjKS72bnNPMrtC
WPec6HX5JVZJTnA6WGexphFb4DPTtgQhEeLjxxqrKUeR2FH/Hvxiwc0qjorB0vbL
8brq6vnEaPhuvJzgOB2fBWoBbYErsQofP/GlEZ4qWO137c8L0kGMWwyG24vlSLmm
7P50kp1N9SyaCj0kBd6Nb0qhX3trhYghrYFAt8pu9u+UilZo6aIFcstF+IFA3wEN
8CAxjbhMsXUicp5WXwW9PyeV6swt9/n0Yj6vwFUFeUjgzFyUn/TRrL4/p3oai5ZP
wWYyINy1k2kje3Nn7+xqPXCq2NejQZsgLFVnwsrq/Nktj0mXshdwEdaMAg3Gdrim
9fYFBKjATguLpPzzATiBJYLgA0crM9ELYuf4CsNinPxaxdGIaeaxzsKSwVkc71+w
uEwUaOv6gBD7oiB2XZoRBanP5DkezrNtXpYjMvbpH9hnn5OoGY/FdRMfC64rdvHU
Ar2lLaOtbAUe1LFy/aUr9y1wy8xZHTzEFbC9d+ZN7NIePSb+I4gZDpVSpEpepXFF
hvFsCvwYbxVanivGVlzcligS/GQY+zF1K8V88DJIsTRpY7tMAcsoKMuHrlGRldFL
7VwAH1BvpdK5fIZ7yv1/bQi5ZMNpKlHqo/MxvvhqGaGC7wkV6GkmWhX4Uq9dUPya
pm8DvkeHPp5DovZVWSZGLwsxw4N2cizmHDY1afS5BMVm/6DLHzto/UujZ9nbf5B5
RHvrocjE7r5hcB4sBe8Vzwgc2Z5WBnFdQSRAM2cKpLMy8o12JlQ2XnGkLTy3nHNe
A3rX4SZvmpusF1JYiJJzh8pSeO7MvO38/rYmiuF7bLykQSR6G2psJumccfvNMOpB
rUGggOc8kU5z6XVrkR03cyqeZtpH7UNglECV5747dgnoHtVBGkQSAUD2V05FaM7V
fczuZQAQRyE6/or/RgEm1n3axVqikBA30j2pfb7krd1cwV9vdKX7N0dURFsjLOZV
/ytRoNZIFCM0A9M14mVGnMr7NKE1CSpONHzR6QSMNgtwPzp4IskUZ2Dwj7O3nTvy
tA8dfGh2PMcENOBmAGD8vF0pcah5YZYufOBiHzHFRqaYAQ2JJwg6Aqne967btI/p
Dw68jr0oVRix5FjgxrlP5CSQECXTOv/fkgkIft5n2cOVTJMOLbMQAUOHeB5UL1hN
wFCu8UYqa9UpDwPhT8x12KWPN1UkThGC1ySSMwlFEIXBDhqkGy52s5iI2mXchn02
zebG1fxUzJUUtDZJoslbXHOflUGrsQ9Hs/X+uCKxOWuRCxB1BABgGTuy/J9JKc3g
u1D2Hv0jlu3yWZ4P95aRin4HH0jEtoY09iLMb1KyKVr/EQ2pqeFP61sQbyRhNJ0S
+KaNJDR3PkuoIJsZGLzRx+d+mw5sq6T87diZCIiHq7LTDKBOnD/Nh0BbgBn4UZf1
iGe8JNhAY/1nGKLRXtEZqc1OX/aJNHBcEH3Irht7xXiQm9UsW9X8iajy3fZK4VGQ
Rydj7jrP3j3rabpBG4xP1IWSvcb4vnZB688WpdpQHbQKnxmBlWMUhiebBn9ezYX9
D2xH5KfmjfSA/UUuHihWHmOxSDrWCEEbVDHAwFRHx04G+hGGDA6Cof/0Gw/KoDpx
feZwYF/RfUivmhdo4DYG0TphCwYqUDaCK9h27epLDJZ3X2++ClPFvBHt1SWkKRU4
+0bcgGpabnBaNYAIwHXT0RzaROS+7TmwrzguLSw/SSuoqCBVB0WcIhljiyoc15yA
GBco+sBjtlciOIRdKxs0jIRn/Z3RZwEwVuQDfw2E0c65I1vcxj4bJLTjvGe0ZlOI
8YKbD8/6dxqTfBiasKkBIm2xfMXt3BI9jDI5ztlBmWGcSmxOP0blqzBR3JRC5f46
iLwmGsyn5iGDguW1vMKAyrC2+9Q/QGjfU0FARCPYwRnq7KuE7U4oTN6aZhpJAKsv
I9PNTABhzKRFr6Nhnxd5LwV7HLCYXevgXHGp1dK6AQj6iGHX2YyRs1+4A2XtSB9e
iy2jTu1n748uR70qgBkPqtKlMLZT7pwIKCobNXFyybSXNdOqSnHs65CHNKHkcfED
pouX3rY8Y7LSZeZZ5yRI9PFWAr830NqdFjfFo/RAK6AzlXOTYViK69AOoGTxLbFk
EF27mVeXnofmLI7tAAtLG1aaPHxTtoMv3qqC0rZZJ+RG6vNnpQIBQw8TTU2sGLYd
Nghy4SfQweme93+saXqHlPHFIb8xMPokJFPE3/7byasvBojirwLME2xOhjGqcWYp
BKo7Z9vBmcLm2YZCXS7H7j2MMHuQAxMmk0R9mexUOPc5vgM/qQitBvyetCTq46GQ
uX3gPZRLX7SP5yTduqOUnFsRGnRTB/k6vsHUq524+ckWtv/8hCzx2v/keEgskEva
J4rBbnLArtLwEIRs7IXqTDNZrdAl1ZPZfYclq2TOkCwLHL0YVAuCypWb1gKbggIh
5IvWXD8w2rnbYzlTUbD7QaPvcEJIh/feHWM0Q4QuNLwlJ5yEiNBt1HgHuoke2aS9
VeyuM0z9zLjPR3fOn+3+MB8iqhCN9l6oSi0qSHs/u+KdDDiROnM39a5NpdimSCTN
KFcxuuaWawomgQbe7MVoZ+uJ62EluYX26Wgm/8ABU7F0TAmEHwK6wNFlLymwZxM4
fSdJSrlApK8czoAKVTJHp7Hc9CBVy6pfkg9uxKNDkEbzRQkVxw/uiIjTQjkXx5ay
KiHNSnzdzGrg/IMeRHkqtCmpw1LxB4eBe5s6ZGpwCMVigkziV0eQ3thajOTH6uXX
EiHynzkKZ5hN5EtvNv8GLTfvCKbV/fsD9OY3ocTQC1MuaxeUAUPu6Qwzj45eTJaI
pFNB4FYDBz4uPLVf7l6Wze/J2mnmxAtrysJ4JYvi1xzk5NF7932P6k/X4tqd1rUD
HjjO9G4PJ0AOIlJGKhnZpXzzRB/RbRy05hgxkewY5Tce2Co9qebaBOU76lNhJZaS
kBJ5ANQWimL7NGayDwb93L3l+kMow7uNqivT1adtFZUPN/EtprhDZTR97ag88YZj
JEj4xp+mLzaC5JAU+YDz2rBoYYFe+u6am9o2tm5+EIZrvmMmRYHsse+Zvw/7UJIY
TqG4RTbEDoX8W8/JRW+ibCgSprgZHH6LbkVmzi3b5d2SXyP1r6LG7A/rYYHf0qhp
cyhR84YcUpeF0ZRnyYsfutIhrSMjHnL4FnzBaOirUbhZfSEfs45iEI+D+bIbHgIp
WXyr3HIz9SWD8Jbx4ovZRkcdwUE01wgm/w26m+e1iGwUTC8GBnK9to2nPvvqlgSo
+7FNd3l80xC12fhXLCOGxEEw92R25oqbLifX/fAtfP4AVB12xs8q/dnO3d6GE5Ep
WAC243wXKl+1tMJ26uHBoIzP1OFAtSSZwY+62XMNKhrkXhUFKykVs9mqfFFaq0IA
RUGNrUI4QAYKeVHvxf+1YIUXMUjPd+mvsGPxDV8EcaZ3L/FdW8WazZgGIqyTFqOU
nrky/+mJTSjARxA+c7r+yoh8HkDjqRfdfOXRRBsFbklg6EfXuSwuUZlRVr2BIsCk
/CJK+OazTcafSN4aDB+NH/YpSr14iPp17tJW4oqIEfAD8ArZ0St6glJQHa5qxkb9
DFNX4M7qP0swzfmgcPM5zz/IZz4zCdGX9031BVq1jcdJCpY5WPiKVWKx8P39uenx
e9uTnnmF0K2edGP1iSIYQRScwJLm2HOGUAuZ8MnPh+HTaOPkYP6t8ondKdUSuNQ3
zfjuKpC0kjT+/cHGBPEwkvxnQiL68ydqjzlEh6yhwzwjXY21l5dg/DH3zd9A/+49
4SGoeN+wNHXyMk1w/n3Fj3XTcbwtugsGFf3eSLlFj0qxEAPP8wBPczSQ2GyOZ6L7
6AZ9chZMg2UHKcxjGaDaknXPis8jadbHilNgr2QjkFVg8hm3Br77cUkDU6/4Zza8
iF76kZauZ6vIS3EnjF01iC0JsLlhDXWfZg3uEWhaATob/KZ7aT3J+gRXY+Bw1Ex4
8/NcJ+Lj2B4TD035CQPL2RnYQR6ZULgt6OSr83F5mSB2BqhFc7jeYAkkvB7vockK
sM+I7NK6eRrInltnWpHFsgpFyv8qd7NVTEWVQNajfAUGOJKcpSGCZFTxhDv0TdPM
shRHjIBQzAUmEsh1CqMTpeY+cDTjxU7ZNCALPYK3qRZbRqCScLIp4Jc+8WqsHykN
K3GSpqG/ZmylfLkWEBD/ed5cv2GjsQRIC9fUyd9Bu+LdHvTCFZXHg2PE+nhfT71v
H6vCDTEfNrfesxg+KhdMtcqzruz/o978CKhlPPghR75Z155lEMDVxhdWphLssVa9
cdaoCn2tIFS+dfK5JUXFRTSKOXFIrSQ6/v2FOf33E4VuoyG8bp5rjOa1MhHy5/f3
H5vwVSxLt2NkuL+R3B40qdmtSVDPh3+zalh2f8T51tt8sb+UWEizDKS0b8wuhxUI
uIw03oz6P9QIepy0LO19NBL4fxmG9Awb01eXvhydSdVOK/Uga7AfqK7ieE0TZWxr
ZTqb03XrJ9xrPe+tzl1PZo5sv0zMt3s2Tzhxcq8AKebAkw3hQtDZq8TvOObHOUsi
EZD4unXbGhDIhpbqyxyIyoTlThrg/2FChywEINRDS/4OqdTrz6HBTZn2u43q3DSX
W1qQB9klAuDaS5mFuwe5804vIcxPqm3dwd4faz+lyv+YYlqXE7ZJR6nHdui0HSWk
M5tHETLMXzoZSp9/7Pray3J9qeppcUGyOj9uhKQHWBjbOAVoLIDkMNrSw5e19K79
wpPSiT84gwIkCwgxR4mBBCWDg6UXeQqEhZ6WjLTk1g9qdESmt0hmgh3k8fRrctyQ
hPEHk1k10STXQNSUbQ4NwDJSMzLkisxC5bvQUsWzquqErmvEOD3sfkVStLo1sp9P
zKndCJBOzf3TkZHXHBgYFfhcupkzIH57UOWMhixxL4F60gobUjNQ40u49JUTsWw6
I6WsyH/b3FbsMfz1uL3B+owL3TYUP2L0FGv6ukdIVheVWz4Tgiw0NTemg0+NIhbx
Xdp3yYaPX+iX0/NQAX1xKlF9QYlUtCVzSTT05Q6T8qA+5vRCjOWcsjeshjltVHxx
HdEojmzTNplbU3ux4UMiY6wnZ5ynv06Y0veqz2HsXb3DmKtpqrFOnBZit6n/Szt6
RqgUuH4OxxHbQlHR5TXDVh6E2NAxLnvggnqqEorqy6JXct5OB9NbYX2evtEbWXbH
NuN7SVgSYJbpqFZmNEXeALhLjVjkw8U41NlXtq9K1uDf7zJQ7c39wV/oY3X5WOuT
PlPKAWWhqiUcHMLkYpsn00tMfhOJBIctJ6BWw7U2EYSeifMAMLHIKR3CrCSBxLry
zFCRTy3GNas3JuS8WcjQOIOkkM8f24zQHVNQ0kjBXOXsZkMMsrle3onAtl09e7YF
3lpuWDqcCzoLzA11iqt6XryUECCVTkC3IYxh4S/ymd87EO653XGENeCGi6hsyHm+
Umq3xQCBLq3pP+TllYaJswv+dVrbBrdWW50DjAS79YZl0E5SG8mWC7WzDiNrnTzL
Gm3z2mBf+AgbjiwAUQJHifJSgL+lNoh8rEb1FiLS3WT85ZgmOFWRLBC/O6BFsda/
JZqegfnjIQLFsa5d2JfWH5B7QK/gkH9CLtAyHr6FHoehFFq0kzvIfCMqtgkeRxMU
lwVD0+b8TeejHCKCaeDcTPCN5D9/CstoAbCsLvlUAL8Y3l1Sg5c2GLjJ1R6FUA9g
bGorQzcowrAsk6vLlQT2lQzrQFggfmJKgjqpNoUgVdM7rVDbZqQTetM+H/cptJ5P
WoZsidTOd5ADzx1HU8ldX2c4Z5OImupzy5Ibuyz8AoJ8J4XRzs3Nlanuhn8b7TIn
fjSexj9qPHhuMqhKqy2ZzmJ6YGFtfQ6Lkwpj3W5DFoDzIVnKa/ctXOfygE3n+FPV
EdlyzHoO3lK0c7QOmoQTBRP1YjQbQkTRHEoFsGCUu57ycp9dIZhQBLac/1vvaeGo
YU/jKODcXp3tDvod9rLN4ckhCcXTckMz73KFw9Y78gbfamPTPi3iMY2rZs5+aP0b
QNMfNw/jIFPtIO7bGqOSrO/3dt/wVhghs6snFo+HRWWMLTwLt2+lvkselOgLwEOG
8PhGiCzljRmiZk6Vm5kzZW8hAv9nbfkp+4G5UIaOSyw9M0URzCt9RiNJ6sIspECa
sd2lMU0u2SPxkxkvBHtYPi/hVPAY6qRKeLi3RjytOwpH98/YNRpa7cYK+rvCBF4H
4L0qP02Ja8Eg5iQzAPEFJLBhAQihCDPODMlCj8tcapM6vzdo7DFMJqQ7Gm9Qm7pF
4EAsQFlqt7IvOr4AExzc6EHy3BBmRsaVlzYgF/6obJTPvxJvJRXp38I5LFQ6CbVj
ltGP3aw859Er2cazWwd9RXrIgPRSrihR8GU/HASbf1HwG0Z8ZHLrPm3W2/FUO0jR
HQUat1v2q2KELZUEIdY/Xm3YTkAJ2hScyItXimCbs6T82kBm6F8RaxddXbBFBg+v
ZxH6ZaRo5o8LeB8tlBOqC6fwfIETmHjNbduIoruRB9H2C886GBHq36kBKTT1nlSE
w29A4iz2LXwYoX7RcJfV5+g9cDX6cxJJ/LuqK3rf3zqqMOdufG/yuNhRORtZXpyn
HkfhnjFCavV9XlHU7J4Y73aNY0Q2gWwBhzOy1xuxD6dsCPXPFVtF+SYdoo2uT7ev
feX9C65av9V5hJ/QuQThgUPUdA27IC84H7DYQLJOv91s/cMMVaAy45X4oDSmL6Zt
Iiu03j67+reHplfzNML/SSQdETf+59yMe+KiTTfB1jFPReZGlUtCp9M2rzwAjBi2
X1o7qZWsilo7eNBZV4EKiJzvC+76WrfJbXi43DfNIoinRJqU/unPDmhcuQ0C5wOv
vHclvxeAa5B+75Xa12staHxHMqp7A67wuoIDcE8Mz4WuX2SXZNayk9aPsXWMyWC3
kS1IOlfT89if9K9faNgAOPwtpP5HJKnY28ZLI8QnThlhIoD9ePtt6w1XdH9QwzTD
4/QIM01NtT0YhxypsHTQRDI4RB+3R0cw5hoM09HpTRWSBuTsdQgzvSYUVx5I9HV4
w8FElxwepAKktFVqINJQDNnLeLm39GL5Ny33QrqxgGykzpqR5LcR7vYAoBqp0nw1
RmaV1PpIzENhDVJnB0Uy5btVPWPIdvgJqzZVDfpnqaEbK+jCddVsl4yC8jVHvk3n
CDG5Y3PmBHvQok6J0uQZcBD/XQHh2imUCzWi6P8NfO7KVXAHR/TX3AE0Oz/exc98
CueOuvg4+TUPV3wH6TlpHX6eafCUd39fRfIyed2LxG3LTzhag4SCLbzYS+vNNqB8
5aV3AdSJsRC4GvrW9WO0e6PyOiB7NAY+Gvduff8oisIXfxyviNL7LgcGCC6cenpG
lDGrPEjWsVAgFwFP2rqIAHGoLljf3Tuyl4LWZoB0FY92H+FD3O+JSZLpoWPtOMVI
ym/T/+oYjbKXGXV6E8HQMCycG8RzBOMMEivVzDZMx/kuS2287MyS6E77pV6Uw3Fg
YxwP3ESG+Vxh8zu6qa5VIAamqLr+bP6lahsPUsh6AT2SJ6/MSdhWYOJxz0f8mCmC
kXHY3t8ArjMLgwg1IY6oKiSEUdC5vRDZJY8PyYTYI1FnvkVMshS0MLLIN6WTzgIW
yOF5izWp6gd+B0wgWRSr8RPgJDnfeFGZBlro21/p5/aueAOz/C3CXiFen74HWcGO
ER3OCWuF0nqP6XYHAFzq0QY2oRL8yrqInnDw4I0DzeaoVF6JrmsvEKrH4ZsjYNyn
f8wVOvLfi2Bj8JUzXooTJFJL1HsyAlpDmcx6y+Ssv9QWy/O3AZna3G1dDt0O28Aj
eTdStqb0uzAQN+MXZJ+fSuaHpXgmIIznFyeFx5gTPahPLLq1pvTcx3n7tyH0USyw
DUwbDd8QkRQo8XFXuithm3tzGJfsWo6zpXLPxkjGySCjySNuLEId8vrE59BTg1gq
bGryn06BJTI7ldP+mDYo62WN+ZIzv/wY1JDP1trFGPyYx7vyTs6Od0z5dndFTUQy
7hFcZHHEGUekTlLLueOxFsTjW/xpSZN9fZGaxy+CauS+WOeOhyHcclqWPOU27fdt
xDxqgEwQTuHGYph9y4ntoXYeixC8P4y7MojLHCOGEqfSN6aPzcKOae+zebKYHar6
oALFABaT/b+oYd5HL6kLQqe9WphhnY3I8biJ7eIUr71KjJPswQs/NGImTgk5ObGb
jBnzn3J5r3kghuRS4MnoL19z8kYHUrWqJvKXRBzGUP7ZMCOi/9JgZBif/H2sxIgR
txSfQxjsreKhFBq8WITadFNggrpEaUowrOqH6q/6lhNFpt4ka0QhFtj0jTkbS3NG
zVcun01YA4PuJ22SEPUcR67UIRSAUemuISdDaSrDpUqxdidGiTj7+VH65XBk82Qv
8Lu6QSx7axbV/rw5f2w1o8dj1CLzPaGkB5ypn64mbDmiHafSuuwns13TKqpr8em8
arZay4NuLtZxutwjuShXCVvlnqliwG8aELnj3DttWkN9HzTnL2mHHEdKb8nXO3/M
un4IQk4yIg1gugGfAH0hqpSSVUnfXMlVsWWHPG97uZ3WDPfMRx67EJozsXUu6TWU
B2oULfOVFF4G+XE8eQNbmXgWY5vmbtxKcBs38vmfETjcjH+qye02dxhXjO8cuD7H
ZbTx3jZn89ylJfw5qk0yMMINubCP1furQQSaqfGXr/PJfOMeN9kke01FGqbNDru1
YUCfGT2rKF2tUF7Hd5LzoyUynubeNgDNQNKuizIezh4cW7LX/Rq/JQqm/2toL7lp
t8fanFY0Q26vfXKmYWDjaeZ9+82SgRlJqpHsGp2LmwarG9gHldKCp2VUKK+wwDen
fJ9VNG+DZ2+eQ1/bF8haz3wXWRn//GjBdzy126BDgRir+IF4qdQuDgNGn+xcXW2/
0epKcc8+WaZOaJenAj0AagMYReV/YTy87m+fgfzNJSyX+8WtD8gjQ7bMCNImnSBk
OXspGoI3nd9/GJ7F6+TQrwT1DXese82GYbVlOT5CBkgSt7Gdi6ZsQJ+0FrKS1GE3
8Eeu2j9IQAhrqBDl8X70yDYmHKlSHoReud+cuVKyvtf423vFaVNpmp3ay9X0ICE+
m6G+U3P9Qbyr4GY8N8oH6t7zaza75uM3zDzpQzfBKtnq9fgWWY3y4zTewn6Fb3gV
2axMHSFYtkgcBJOepL3ngbdC2+LKH3r2YYk8H5WKSDy0e9+Fha8CVyFw0Y4BNW1y
tj4Cu2VycPVwWg84JSppoqXQuON+LdnNtNvJsyRCO5aYLiHWzkGZ3ZA5JY/YHJwv
DIiwqQd1ajE01Cjn8hwPLSKQi/1Sro8QkjmLCEMQcnfSeixhGtny03fW8aSaDbZX
mPKSqd6NpxZ8ROb7kRbVphunTcsmiZsxU90kJetikddtwrfRRaNX6E5cLrkCP60f
chkGw6ylVIu407H1bpWeosk6rLfyjwvsC0ez/c8JfvLVki0C1r1cyVJwTTmEvb6Q
vpUrYUy8tmDFEGakjZr6ZrvUCCk/Xth3+tKsOO33rZ31kSOV0PWjEPIYJLLiylAf
aIclGVTLEn61PkS4eMA11WvMqjh79SjoSAb/BE2jg3vqM28tC0IL3mit1iWavzy2
ZmpIb3znbiOVbbGkXwhZaxoAuI3Spy6TED2OoSlc5qny3HF6efVYt88wUvQUo91e
z2yAb0vvWuXeO49R+mT17CCj6J8X2qBjDOk2eeyl43GzrjR/urgFwX/Qy1D6BmfQ
EviFad+u8BfWAa9UA83T8zg9HoIaIulo62iwQrJBSrTdpW9dXgEcTAo+6epA9lu6
FltKOE28XLIgnnUY1bkT0PlstY2Hw+Pf//itVnm74Vs9z6Uzwjzvphz20JwMY3fE
ULEm3iXVWvemOjGmzt0lZpAfa2g5x2+2KSZ7zNHzOprc2GsZ1hyVW+3/ixhObUDO
XHhwaT2r/rjK+uuHIA4q4KYGYxieBgs1ZeaGjtrYggJ/xyfQGGa7rKXgj8RnXV0G
/SWJdKk1nI3VE9Z7/juypwwXcvSehV7zRKAOqzCIpNztgzWjnwneL7Lk4PyPT5J8
smDOumidnispC9IDvcaPVWPeHjHY+/JB2Vq5mp2HochUuNvoMZvrb2nNTdPL8+2B
b0CjJkrqnFOLlbql9WcLjR5OoYdjTZwp/itOtzaZJXMzeREinisd1/DVSGgD+l58
9y9g+uonCZzYOvt8+ytxMyil/eCsnhruQ9JCbEhrb0qAyUvIz7axlx61ojyJDQdC
p5JsUL6m5CsfHFXE6Oazf1zhQ41/cTUr2Ir4H6v+uqmxnCFFMFcSixU7njBXqvfl
S1TurVLpoI+DBMzdz+tVxKjDwPgVVuqaWD/yMIRmZIjoSo57BF2b93x7N6iYKajB
O2nnCkdcsPa9aqtaDKv5EsComylkAofbtf7IXj9b8E8joqBinaJ6vtDRF8Eu9iVX
7GH6VapyHXKQsnFpfHn7rTa7Lu84J14qxVUvt2FiCTsMPKaFPuRSl0MfzXR7UIrP
T4oWMqujx6obbDNXiT1ad1pbcO3iRhdyIS+T++RfJGECEr8a158SAPbQlQFw/dot
JvKUkM0o1suVj+SfTcWtUlZ4f/TpmTXeoVWU2Na3hoc+AXI9+nobCOhqK0MCxcaA
WbX40t59IkbaTo8/8P/b1u/lNjcPD4X9qet0LF5wNoP6fFc1rPMnPcOP8jed9k0H
9X8uBU0Mu4/bab6933YOJhaP+vzLOGctqhi1Hv5rFvqZmZQWVw/I2pqT47iLJAvy
3cO9w+r7JvuKMA5Nypl1wTEkRexlWajou5yPhjyUx2ay2EukyFvnC7242Ar8IBLT
VT1m7riL4/Z5CmGSgYhI4b93MjZlmRCGP/qV12jjv1AzcFBM+oFH9h3BAYiHMioA
5G6nEkyrperhiAFLr68bK63zopDSuky/ULxO+zLaSUYgWCzycoH/xrWIV3vOU60D
K965c5ZgX9QvGUylH46HDilQfD+8E2i++eoXCSz95dyIdpNRu0ZWFAwLcmLwVsjq
4ws5MzUns12QzT1BSyEKc0T8S9Gk59K3/L1FHEFOr4gsUvjlDQJPoNnl1N9vD7Dw
w9gHjkbIVxeU/GHFThuiuOFy8MuhVYtb9FoQ+nXpL53nAZ2xQ5xgVLoEzDo4rgOo
jPO4ocK6RksXxZudsZzlZVcSsRva07mw+ZFYgrr09R3yN0bOmfbZ8vRy67uTKZTZ
YCP9wbvzJq/3ECmotpYsnin4fmYY2CDiPlBfo+v524fhoTCUPZ0e1LAM8TeRAj9w
o5A/isd8scAOCqmPfjOH9h/hMUlw3l3aYF7sibNBwjHgqf5VGd8LTA5DGrEiH4aY
jg+ZSUbgZr7IJqd5UqSwC+mYW8u6wdPahP2wng5pVZwZFKzbfKqcj6NxUAi3rjGx
eetv1Kt6s8zfytS5hX439FDGqxAKVDtbwhE/NiLx+eyCT6WCHnfB7J3lUrZnMeYf
JTVi3cIA0OYc1or17KVrnJJfrlhNwgEGDSIHJJvXPfgYk5rj8TNHhRcmgl8N2e3D
r8/dwJKfy9wINZoqURdHiR/RIF/Uui/f/4smRT8j6J+1D6Y3aXRH9q9FXE3NVymx
IFbhQ0WY/KuUN+KNHiNLt5jCHCctKtKEv/KVvPTm3jbvJUTngXpsdgrYqCTkHTOy
qBHB7NJQ1KXmNRo7A1GfvYWErwRkIKbk9zZl7xViRhVPUuhYkoFy9IXPrqcHZ52f
A7WJaK4Mb/eJtpB5trtkBwqwyaPr5Zb+1fcOkApGVOP79xnHbfCxsTKlC2rJIY3J
eFN6De1jhWkJlJWtyBSt0TpQN1ZCEoYZ1sSnhP7eVgQAnR9X4BH5G1rF117iJAz1
a0k3THTWSKbYLOAaAttyJZSowbsONWr4oJVt7226pxUVg5Fhk1aZs2yJKcmK7ou7
U0nQ+YKPv/bzPWkLiApItRatxX8Sng4dcOoJRzHI9GnZT7nmJz6LPvLT2KeobG7/
K51ESqQxo2UR+IedDSLTgpuCzxjWhKlKe1h8HF1A2PANMoG+WKhzF7fyZLQcZosY
3z3Nl4d594f3gxra/HiaWunVRBpQkyBhSSHvLCeGhOp/F10ULKSBbw9EpNnLoQ+C
eScP6MgD+2QL5A8R+6VvBAKScJ2q4NZC2lOtdL1C/xbEAquAs+EKucPcRcTOvIc+
BmQtKHvdtikrT4rLtL9P+ICzxeiwHy9q5owbYG9NxtnY8cRZZBtNjWQt3JV3tM4P
fNL+KDWGrnVoKGkx0PTS5H7nqOSdd8CuS7L9fPxebBLAlr79+0modG1act/fI1lU
kYxUXWl42CXm7EeAPKLBJK+U0Q0RqZ3rlYXla45HX1A1PAnSQoiOb6cwIpoDJbXY
ej6ZpnGososE7rMXQAo99vAq+u0H5jQXjgv6/fvvHgJFGasyZ83xjwKEqgL++9qX
TZgku8dvUwG70mfN57a98ztelg/tq+YwuCFJakO8gqsyqsDC0QP27jkM5hvQdwDf
KiPEGqzldG4Zi5sLdCKUIhMp54s16u9MDr9Q4n+U9S/SlK/+sIRYriJBz6OsBqXP
YpMz8TynyGY8BEMNnobyAYv3L4MFg4K9iyoJc1KLvmQhtjK4LzpwgCcQKe1UFVbe
pvqEpEgnuO7Cmd4tabFMku82ingZBht2D/ezI6zhCAglZqB4HyAF7t8abiavoTjI
CsbALoZQv1VSj7dQp6TfjrD8+nxC7ysiHYsw4iKQRy4jvxN7kEQVVJfZTtjC7WBA
YC7vcA8TONflzDcVYSNnrB7aAMqn1O9gdkGEAMuPyTxSRBadhiNGCw4tgaohiIJX
AxwwvmfHEeaISnvLswfPfnHGSCKRXVz0oi8O9YUBquQYhoo3pea3VA/fE9R6g1e9
7Y+wQhaM65acGBMXMkrR3/DwVzBdX13F6RvUk/7szJYn9OOfXK+W2BGjMflpPIfE
L8nueZapdZo7jiiVjSSmhO224TzUpUTwMd3F5spLow8e5r2H7hL7KrWB6tF7esZm
YYXTPmgl9EARiU7HREi/T+vkuzaddg5E8v+niKZs6ZQ3yJmoNTJqSAQFayggzXi+
A6PM1fHSHOSWfFmPwldDI0YqG9JEbH1TVp1SJJWzcDam69nVABXSIjWauuqpc1oA
IEjX6VtNt+XXB386wQrmnVqt3YrI11BYdfsqpecAYF0voZ2UPvqRROj6T9eKFZhG
6f5K6m8N9+Wjneb8d8iYxMZyeAImmFTCxPzLGbCbdrYzA/V+XCeLwZN1fGBJer9D
CDj5M8JL/NZ34GaW9Gi73fsha2zJu5rlxQdlXWKaHccBnorh+SUTbxvb8pxdPBW6
EeoJ10c86PqQOOuaO7V+QpC8cuKIl+IbngtzqfZiSNlNVuxZ8sUcfRVfWF6MMoOR
ZOkr1yIUtywLaR65Sw+W22TvlqRwRgkHyJFLIpLww8oqeM3SUL57YC0qic/EQxjb
t6MC1RY4I/7smBLNPWuHym9hgSeJQTA0tnXy+TUFXsLM0oxAQ6JJUmDWyd+B2wu4
k79KpDi+0VQt4mO0QASiA+Hn1faXjUxgoeNyBxt+XRsnhHJHYjKInHnAGR9XKwfZ
BLlwIAzYtW1ys9l+WYC0RPmW7vk7CzQzfcFlG+JdzGU0RHRM4VrWywDdGXJK2M01
zguoOiJdIHUCJMBwe/IrKQ61jUTouNsaMorVCHTAWMksrzpB/E6Yg3yNH64cjx0y
TkxF+dkxtp4RedOzur7LtWGWSeAPo/0Nw7//jin2/LDxooqZpS0AAiwyJd1mMu6L
hZOD+frayv24BmD4EWmoMzi93kwHY7gcFIfa+9/ls7tlHst4ALNHj+6fNfKFHkcO
Ke73CbnzRPkjmeyAKNufn9b93es2N3C2O9s0P1DjOjvLZtzvU3fIujumfWoy66gf
cDxpZdr8T2AXyy7poIAkG/NvzaLnkK4sf7tXNl9CPSbp+ZuQ7ri1X+EY7cAYtUIq
Z1RBioRdjlE44luly0p9l6dWGmllD9p6dOCV+KwwooaWzo09BPg+mziTT+sa4Eie
3J9zHkPog/Kp5luOFEUHSV41475RoM/8l4wg6JSwdnxu0EztYR+z9ao9GZJ/rSgH
XGmoqxX4VPCXEqDN/b3Ik78z1vTNaOm3zOhgEfM4TlBA1G6T+b3feuZNOHcSkRNh
ZymFtBMMX+0Okvyew32YLiOMi8uFmyZPXlx4+t2+0vJX/xMGLKf8/rpZZfwMQmkI
SEZjYQ6wpFGVgr4Pi2ZkQmNwN7Q529eQ9/fGhA3MxkrvfOFRCfokuBjslbIgptlH
sxB4kh3bNcEtiLvJV1DeC0w9nsVZDlRwQgnPri2ZRPthK5VeIfF185c/CGtH8Q9T
HOgIo28MLOzLWkm7vdeJ+xLDm1Q2R538l26hQVbkj5ZYCSQzTjEPn6zym9ahDX2u
Jg0aDJ+/nZAZDdFaS7xq2IOg4DyrNG6tculrChwcChAtNl4W7FpgEV43P5zbb72s
3dmoIwJZpfOmkpPuF7RC0yFoPAuhDMGPHNCPo6KPaac2mIKvPUuXufkagPsGL/7+
gw64/BaeiYP8G1rIbV3P4Jj67dQUdAr9Crwd7TYNhv9mmpsU6IOVTj7n2strBYrk
uwot0WvdMrlt9AIWVnqFi7V9WSuMoTuqEZkwXDBR0zo0IExvtEYTNNbptbC4MONa
+lxt0dlV6MwBt3hX/AVMATtKDcfTUK8/E16vOtKaVn4rXYUuudFUG5W2AIyM1c6d
l0Z6M8vtuFvtjSxfIUGMO18Ue5wsqAeA8DDu/5s/eKVBorfrdwjAoDPklNsvnRvj
BRMwVosJ4Bcsi4qFRiOgVAKjQ1yq0clcslKZXW3DsouhkNoW+IK1QP+SVcr9MCKG
Jd/d4NebVXk+bqkT/25CyChynbUUHuIn7R0+j/Sit9FH1eo4uFpRqEm/KCHnKkvo
wBAZCl8vKQGMnO+VVpPHmDTxaRQPLHVSUL9ReIKkUBFu0JJXz1XwGWH0bXmN4btA
QW2CTyEMZQwF6AzFIQ+f6N/PCRB05bRtsy5nOsqwCTmnxRs/X0swALA6n3FA4pRn
0JhFysgjgprDpEBUvovaFCbxl4gV13tZUaBInjq78ohBmJ2UHY4SHa7CLY1aQqAz
yqJZLFTM4pU2tegcQfuF/oEk00lCAE4N308U/P/zJtB+qsK9Fz9FAZMMuy35hJm9
jIJfddPBUKqU/Kp2V1fZF45oAwFA4K40nIye3apozyKbGawcoxAWcLwvHzCUzDe5
wOWj5derpXp83ioNPGIo/vkpt2aKg2oMUkacpXTWUmAv6DuayHmgpk2Km7W8HMIb
WfjTvpdTch3ugU8MRcSDMUQUOdzBxFEm0WNURykifpzbB6MJ84K9rQFPDgpbfpVw
Ib6zUUtJZweEliIkykTX6MEedddbnRpBWXMzYkJr6V86irB+oQYjeC9ZLYnG/+Fi
Lx1dCcNVRF6o5nxZC2IsUPTvYrM8BkP8+hEXuOzyUJFyFKMHVhd7+kXUDVBeDOum
/+gKai6mmGsSpvhFi2Hx5Iu7ZM7UKvPY0pgU2CSK9KxbSa2TRQWDD/YNmM+NYRC4
DmfCNuKUYMOplCn5NBVA+He5aNn2AWkF02VwRkM0ETR1+i/3b29NkIrF7nP+zKsy
Ykrp26tzg6/r440VUffU8ilawKR7wR0/frag3nZ6DleBdyVgw597xc2Vgcjj/pST
BgWhgnnFFRMOX/nAJiWapE639oi6KgjHkSCDARyM6Vu69AqBsocQ/ze7hs4mwYVO
1gYxcF3oUOZcXdub9xLcvIVJbw0OGk6eS947BS6jvUm5SWZkfcYYu7l4yBrooYsr
vxp1xnD9naYhYjX9etWCT74OWfpLLq5KFC87Uy+YIN6ZhZ7RXGhYLIwfJsrEbj3C
Ihv0DaFcDDcvlWudQHV6rDe+g8CHdLC9xAfXcgFqks15RroBmKcxETAATLbxS5Od
tJsLks1KPSZLmBFD2pqXhCL5eb4uiDgZo3IVLuo4bYWvm7Ct0sAIRa8ydMwWu/Vv
RG5RIYpO1V+I+hlKscK/Dp5hZkB+La+QSTw8UwVaTA/33RXUd2Hc9f8lqKKdb3yk
lV5iPvgo4QppkLvNnpr8gY0DDmaZfuDwFdg426o+mHrFtZ57jN8oRaPgeAR6f95w
qCy1CmadQI3mnBuKu9edN5cJsYqEs0P7VgDsXPXsKBoryH4EznWMcU2laSssGOqQ
Em7BntrqTkbDoMm0ylGX+7rFuEGGN3GkrZtutsSgVw39uKOlWVleM8LGRMCFHXtn
f7y4TxvyJECD3nuh2D0KxCLeVKLa0SJA6yOmsqzkyMLdiDSdUd3shvyN6s9u90g3
XIBtA3pojg1Qo4EX7mOSHsXtqb1hGpB+FlzL0im7ggX94Y7ZxTciyybJMKEUK92f
VmtBF0YRk2Ep7ivgjWvk/pZ6zUkjva5l9RFSaM/VazHUJIUSY9WgzHrmPXR0lI9/
11S6QVSB+dUjIxf/iD2YiftsVqU/YGXUw7BUXnwHlfksW/8xGNai7thoQaVSIBLf
lmmLvNW//gw1NpJCVKBrySaTptDtLcewZry6ay57E3OfTrXy1k8yW2STULDNMBrk
gXyIt7aWuFZtVFOOtG6Nf5OrXQkrAFw1P4S5QGuNSWpzs0Xe72Wk2v1dqTlbyWLe
vMwwAi6TNzdwVTiK/pgIMRBZ2S4awHs7k+41l0Kd2gN2zf0sAIe+AE1USHDnsGt1
5DIfWfvAPsc3JLKmBgwJymYKfs/EYHsTd4Q4IWwp7Ga3C2CekRtYr2/AVmajw1Xc
x/6tPBR8ShW77uz9fw3bRnB0iwU+f2RjLwGXF4rfhS39rFJlIrikGMBiBoDw154n
YorQwLyXpWCIfn5Lqz1cxOlizUA3h6D9bNjIZkl5/ga8JcvZ70gGw62RBMPbHP8I
er8rPloNhtGkKfJxISgYGT8fU0xG1z7sOgSCC3LpMjl0hWma4QHSHDMyhKeww2Iq
0h8JMyzjidX4zZVv0zrn3tmhQ499BaypQWGj+b1oeF7wf++VUSd3AqAu8M9RzVJo
Hdtkyp8Jl2tLmmtt9VpLqdBhuCHt6m+Tar7mnJzt+1SLCptjiVjv83dQZppdhomO
HW4bYdGCdwIpGcB5z4hidYM0CpLIgC7HbyqXl6jZLF/Ylr1lnqtXrXkecbDON386
Jvddu2D8nQGUa201Q4C6YyYTHYNHru4ktt/+JvKmIEYaAERry0eKF4nC+voPobKt
4T+Xl0dNmObred8iYm/L8D+KcPoNMbAvQ5V0Vm99AjnXWMZkLUXpCtolXA0ThZ1L
YJaUyBOWC5XsUg8wOc8RubUClZ7g+Lq4GT0WyvI0R7SFBc1RTyqaIJXHGNbHqI4U
v8L46C/15rCBq7akKs05ImN1JsMqlAgj1quzogeCn80suXSUpgGYX7R2FoKgKjhh
IcBZK9lS7KT+eQTP+pKOPz+4gbQi1pAVZsVW9aC8oaekJRkUuz7op09lAcKzeX7j
JP7IUqdwfkGcpKTg+tIswQI7aCXHKF7887Etqtuf+B6C2nlgQnX4DLtb4fKmLunG
tBK8U8ZuQlroU95SaRznnw9rwxo7Dy55qibD7Y3uu57j+Q1G3Wu2k7JEFpk0pqso
y+UTYTvcLL5UANnQaPWqdkYoqeEOrXiC0GDXq2lTZv3prvZcEjF3hpVl/hCy7SH2
gmrIPuR4dor0z667D7+oPfH1aXkFXNaQ/WeJjZlqSDNyMw+vn/a+VYC8I2AQmmDF
NCVZrEU9VfKyrkPtO9OT5u8uPttFwM0SIBoojBXq079WdCtGqwrlYv/qnu5CZXOK
oDcCG+SKsNwjcWiwZNcMcV3fJHYkBZ3VePHpFzx6I25penfK8Hq48lfjhkrU2ZTS
zZWeknkQnkOTFX5x4HPDvfhTxTjrIFegqEFlLaeHO+u/9FVU99ybsuvtC6lKnU5/
xLPJcDi6RVjr2oGskgL/F08lRNBeJ7IECO2jBA6vchBc+BWsJ6iiUCxSbQNh1VpV
MZD3E9AtU3glwZfNj5q9ByMmsLIDtbJlzu1E26dRHzP+FiT/vkyAT/c4/Ay5pvp5
iVKPTqGNnAPCHzX/Ex2VFYW9QDsSyGsyhwlmtUfWxLFfR8CwZ4D53dmBN/MjqJCs
rQ8IE5klSGpFs4xCXtp5nlwj0YYqcSNpRYNmFPnI5YS792QOmg4t0HpNjwW8at1i
25gbRGanHBUyUtyr2OU63Z3oWZwWt2HyDjc3IlgGae/eiJ77CJzHxCKxRLT2VZen
58XZgca3J402Q+TnkGiiXd0f7cfofqjaquSmzOr2KtRkJ7Edmt2X8pxXjqeSnjR9
KU7B2qcx3pZAxK4gtZe4VJqFnTDhHNg7CG4N0vtJ3Tffb1g78B1oGN0ZiubmlxFG
ueSf3YzAOL+F217DKrTMSKEZCoQRxbPPZRrxRrGhal6aYQ7s86L+moOFZSr7J+PN
64YSLhc7v8LnWtuZ+kRyWgbHWsFtO6eYNKoWGp3/KrRb+e4ng3fz6L0KUWn4xkq8
M7p8NyxjGH5FAfvI/GAEKqqFG2jx6yVoaWwnVhO73H6iLzU7Z1HRInCyfHjB3Kg1
VCnmeoomfbXcWw+pu6rZiQ9MInINO/0uRAJYtc1WXEtO7U2tGaS9lXQbAizehxOS
KWDWjf1kISNojjir7/tgq40y0RJuI4nXiLCwDeozgxpX9nsc1+oTgJ3z7ydQi6iE
XBPcDEwLfRLOx4N58gC+IEG1gUTpPa1WhJU+st4gocBbon4OCq4jmO4xGBb/KuRY
dLh0AmC81UFi5+j4dx4F0fCfTmld0mh8lkJIJXySmFF2Jifebgl5+CcFpvBuuJ6C
4kA+6ltt5LQIbY7Vk5xbC5Xlkb/lahM2aQ/IxpMYk4MTBPVpGSuOPoTWRAvjDJfV
mW8zXtndpGAAF3rcPE99CAqfMTQSSX2RO2OBuIregLayu9J2IaVVvvq59CXT87rF
l4AE5dAFEVmrdLtFx9TotyovpmSe5EwKxpMIflYeQjBfm65PHYMJ7CdAZmCROKJd
7cL+oQbeNei92A6/O4j1IY+tFJ0yaSGNPrka6MMHZstm7x1NtjFYCxaLCi/DKx3M
HxLpMZtQ2mijiLB7FMVrh2F84f64wJg6cAoaaGxMjyZa2c30RrP4PUXqNGY9JNB4
UkYiOJVhT+cRAB+wAtBHINHFVD0oclsCgO0YZDk9EzmyTXYUmV/IVPmifH2k38ia
1OiPoe2YxwfrndWh4iy/wQ1P0vFVCdRyDVrTQG81Fr0sXrsDgDMUub7HE9prMtD5
o3v+My0zmWFAopXrByrAkCdydYvMABSPAVd6PmZSKAHgytP0lsrT6c3f3x+M2gN3
vrv2Ux3AAwVzg1nJL5Y5r0gy5TYoQaDilZc6pzRnAyfDRz3rCSYrDKVSgB2gWPoQ
cmrjmYcrJQi2Se+CKQkketOK1FR5y8JCyAvW71F47jskr+pfn1WqWrrtLrSTBPwx
vqdlSff3MtnIT9h6BdoxwUQPtyCCRl/4micN49fLs1hvSrV/ekIddMK2pXl+hzAw
xBtrYGcThU+Lm0Nz5Mk1SJ5sEfocFpxsmgxpMj0bwyMLQFveChykrxEdz7oquKSK
9syVMc4J5MeJ37iimx67gV0PHaKwCptE0TiOlZwsHo4wJsg1GhDZVW102Jgqmwsu
iY7T4W79c8r5e1C2gyuBer8IBp32GJcwkiGUlWNUcFZ9TnFd646Zd5ADH3JPEfYD
I2Qqorvv/+ZyuumQQkljG4nCEbu18GZXR+ppzRXB662t1s9QpqyTyFauTvjKjb9h
s4fZPiZggX32iLYjh3oKfHU5u6lg5TN9Fqa3j0XAfU3IOe3mDE/K3JkGpR1cpHlb
vR8aAe/7gfFaapOQzodc/lxiifZvDnLOOZiB8beAS4Vj+BiHEPHasSjP7U9pI8sN
u60BqLTR4n7/8SS6zT1KxUwKaNX7J1p3jQ2ds3Lk841hL55Sit3JcWsh6N2wOjeh
VY8LZqnbjfTH6A9VjKjxMhpSxXSoqZwhQuhjLG1ZbNkPqX4Hg3pEbJgd6YRfILZp
l3ZksN+UJGIRl9aiQPdGkMb5W9JxClDYFIW1ZAc6C+4UMuMsR+Sg4dknn5PhjqnB
2iIWmtOHvuuOvA2vLSy0Kiv1tfaCTurKUyEr60f3azEM7U0dBN94roq4LLH+Wf8X
sm2+d95mD9B89qZN9YbkUarETHfxP6Y6MsaaF6ro/PyeRQu1tmHC4CUawLMzyriB
HT6FqXiMW4VMZhf+an89Q23WGb78gKcQECzO3oIHlGNRSvYcTu6wCWcQCfRORZqw
0l1poT3Qsjm/Q2dwNC8GzDwQhdMsf1Xl/+67c9Lr9yNk256kPPKPWHLgsE15yKrM
A77cIbNDTES5wZOItcY0Wy6Dw+YNLzjrmX8Jn6cORjHgYCLyK57ExDjx7paw+GnA
Ton+gYMMNY/U4cTZ/6KVPZUCqE+eivA5eFtmHKYUo5p9yDf0Dr4KY28MrhEiGi77
JVZUMTjc88D/vzCw2SsnkLBxUTtwXKFI4rl70kJH5APYEiPZvepPMVOtiOz8Y0Xh
fknIzH8pGdzbEm4l36UeGyDfWTI/ycGbD8PyL8lu9VCZ8YJHdZIQYYCP1zsOAPYa
nWy+YZlxAegF6JfoSk5KZl3LxpvhY/9KaODU6RP/l3AEQQk7v8clENqcjl9Wz/5C
aFSigYYusTBwFzis+KSoeZz3J0uS76Zvvi4+lVQZmmRa/6Yt/sS7sCRsRGfdS6Q6
RPQtX5HZTQ0ctEp2TPHTMdVicvMeyGfxHhEGFwUuoS8LUmm+jyMC2v7JWppcRwPG
RfaasJQeWAYVfaO5viN0VEFUodGwJYPjQ5T3970v3nTvKmtxAP+S+x/Gc97nIad6
IZjkFHg+UCC4Y242Iy242sPTLXUUFZ2bICdlS/xSuA0LBuc3/1SUaVUEXf4GjY85
6h3yrouP85D4ejgvT6FBRTpBugKG5Li9lxziAbBXmtMZddqym5N/SHJSo9/Hu9He
iSXIo4MgRSpcL62sw6cvIF9GKhaITCXGXLdfS/1FSwVARSAuvftM6Ch2joQV2cV/
rfC7uN2ZuHz3Q4Ke/23IXd59s6uZa+AcxViY0afEnBnrMlmwDBnPSKvSyXQgd7rX
cYKKX6clMjK9A1K24rWfI/SWVSlKi2X0ehW2UBfQz7efRZSkax53+mi1w/GcrAfY
KsdPjWlGcBkWOlyJgKxv1DrrtVyFisjFGAkvnbclk7sqTJAHIzQmdekWukwRAg/w
jHoK1TIskpc+kETEd41fpenhqWR9NQ/u1bIy7SNhB2qWysCIm4cgg/MbAb+2F/L0
va3xYJKYjTiCsR/JuEGzLHjv5cT1Zs7Meaoz00mw4i4zuOx6Cg/MYUqRnxYChjGs
bN0euyyMqXG35pCLwgDGpJsrTcgZsWj/stvn1EhfSE5PML5SsCKCmrcUbti/YCvr
6xoJzs0IN9RAO1ilcguhWQHZthJ08b4gLLeN6pqzpCk1tmdCRkTXnlAHQURFnnk6
WMRVnq+qTSHr0wvrAsliasKRCCcCd+bkwsNBaiumWJ7cJ4Qg2th9hGCJopxKHMmf
UdZOCWNudl3ziDI7zLsuwQpSUE8Eip0QW9qxHFzR+swwiy9jLa6RYIva4gAsO8Fj
Y/amjMMaF0O9IICYsP3dCUd2MQPn+OITC+vbfzFDMulULU6hXZ+IGL4GzBFcwoub
AE5pDRvAFFcF7lyFLL7jafP/oJiNe/onLQ0XW76JJipxswg22OnQeXw/AHHIz5vm
vGtS+4byACgOe2S6fz5We11+jgDJhZJRjSb9Na0gbXCl2Jdh2tr0qdS1S/Ti91zu
qEoYcroQfGQb0xxgq37/2AR4eXtyqiM8B4eDpTUB1RAP06FDuYPi/kx8/7sEtKWa
qaZUxLzp94e6WypryfQGgedFhWBQqIlDnjfm+X2ktGMxXOXqyXqAzBv1D+b0ivxR
/i/wjZyRzepg27x+cjRU3j63x8ylX49328PmE8OE0HeqHm5bSHad4qUi9J7kZraz
vx4M4H1Da8O5HznCDlkvyLI8UPKibwKRaSR3JNn2XeBMgJVvoB3myprxib2X0Khi
12Ax3LUy1HXTRFha7TzaG6TEZs77jTKXABYycu0QwSCpyG/XchcQyay3EJGYGZy7
Dk7oWCCe0fzmx26Mj6oC3jNoiQh8likSO1+pcJv8l2K2Fs82EDrdmhjkVnXhq2xI
pSpbe4Y5+pGiLwFCP2GOmKlb2DpOMuEAFpBGSsyHyZgK7TeQ6iND4W9g6kLjZEap
KfaWLr0RxAk77wmMImEX0sF7sivDpD0iQuXvhrlxlXIDUaKHPlm1ARsn98Dujx36
H9RD2doeb9gcE2kyUjfyI38A+5mB7Iua70MXTF776NXiUUXftJXy9DZIE4ToJfdJ
X33ZFObrjM+iCLu+lTfxAHqRDUywEOYZYuneufdQ/7x2N+S5u/2iB8lIEmP7C4KE
FwROL6ekIPYaDyLS/7CwbxzXDiFFTjAK67MNH4M8gWyOGqb9+KVW3LqSstNkI7I7
SRrH+XEunrS4BD/TknqRj5Ry4lLqeay+SmCeLrV0zIS91cBjcORcQsQFGTNhQr/n
LVcxeH8vRXQovC5EpdhnYzwit6UuuMVSD3EINQlEorZLPshyvQnGGokDqV7Spb9R
VkcJAmUESRa6QVmZqeSoMCTnG7zH1jXw3Gx41Cz7ljj9ADeU66oZ7HCOz0ZNydBl
bGz5W3OclV1QmifJXZqSUzLnWknjHB12hY31Y+WQ6cILBa9t7oLuFOVmMN2DlDL8
qL08O7GLfXRoB7akHV+fY7Wt6WgPVOLZZuVlFYJg9r8GIVG1Oh2/DO1HQAZKnZgp
VBBryuMDv6o6NWnOOyE0TYnXg4u4U/es6U5xZufFjFZFosj2YR3wlFU+k3jZjwH/
kwPHZ+JY7Iv/NMB3cTxf/pyn2tmcEEciwI0N0hV0WXw2u4Yy+Udr2jJu2sRLzruk
bloNx0V8Xn42o79PhM5G2MPaNYC3Vjegh+3YdKICPe1VQy8GXNzGttHnWhgd03m9
Q2QEmtNqHo3HC4m6XwVgYZnjyHbMzNwqJhu+UOxFcFCHce8n3RedS/GVfS6ohphJ
7WpJ85P2nXNv2GwMfZ/iJ8fiwWz7dgfrr8JOs+006j9sdbuBkvuFh/yHrJFehs+R
H0myYdl6knZ33k3q3uEEoFvy5E0W1gjfRksNbOSdqfOeIBBimhOnYBVYlrg02bSc
//x/h8WZv8AKZFenS5AwUGiFg9u0ta0TceZtgz1SA10TQJ+18uu34QfWxyIewtSG
eAFJ6qX1h3UR9mAIMDJ4v/6rGbHato31BpJG2RzgEeLbA1EKfpgB7EPyhme7iCBW
mefbJ8FncHHnwyqlfaQiRjbentCHPEJVnNU6aHOQtDtlQGItGXH/amcBEiKBkhJe
RRtuOcvE6HbjTeCvEKE+qUZir4z6XcMXHTpjOGW/z4dtTB718Bx8oBF4+Y8qV6v0
MSL0JXptEjfWGk+ooublu0eC7RRyLTvrmv2Fdzx6S4eRh+GaLMMHL/npgw3Ck6pc
BQP2qQfxTwYKVKt3/EX4tjY13XH+60hq/zl2ojPQJY1wnuTGJr0vP3/PD3Pc0LMy
ol0eoGqITF4v5dihWvgLoWiA0sQTQ7WFtFx56ayS4n3tCTPdfUXghgJa+L/ZHBFD
JlK0WQVqKhfuonTnLu4CJWO4rNLPQtwuBMyaMgPSObHl+c15WsYNLid6o32/QM36
MM6a+4UPvDZYKzDODpv09gDL+mPWKdG8Rk2l1pp/Spctf3k1+Q0eAxYPmUPh7kZm
mxQTlYz5q8JSMeXWEGQXpMJLfvVvCmXeusqp/5cY+U+6OvOXBOP5pVaib0Wqz+b7
fO2KhYEEWvfRtxCJsQfdnS+K+paY04v2tmPZXLIq76quoT9bHfBiXqLzdILBgFTV
cb9HV56JrABO2imgVGlkTT2VW47wfNUog6azXpwtOrJqqQ3hl35QVkruZW55So76
3csE2tUQVoqIwukxu5sZ/shkldFWpmJL6le2nilr0ZJ299BlqxDX/KFEK0YSJwvh
aOls9iMTHL1tnjT/ctSgrFT/m3yfdbndmx06GlGto9WUOi7fvueKQU4bREmvwEre
sj9BlmI3vyTQx0hKfsc2Pf4Fb0RlkzIbuh0pQDz5L3N+Nf6Oyg6tL34uvWbAa9fM
9crMzxkCDL5ndeO7TAXU6ZKHpX1dy0cbvfzst6PtOuLmq8PErKAYgqqkPU8IxFy9
33huZFBQck/zIxFuC6bLgHHU/AzOywoFVcoCOGT/G1lFMI4Q8AHI5RhA3Rt5+NgH
EYL1P87opSJzVJoFcvWspnUDOHYWcc9uq2xd4fVeBlnVJ0DaouB+7BRaf/2LEM/D
U/+K1goNstpr7/FCmqZiN305QULfPAo0RCwYbinhiZ+8XNOGVi75wHgPE0ECkcle
E8dg422gywsY142TcbnFxDEBRvqLTEMOXDgcuBTuhF+JBvkOXNGSFUpFzn2MyGmt
8GQaJs5fXojGvfGDMEcSoZizTATiTwmsglVB6/rdAROAbxgfxS032JFoNK7wRWDi
KfIKaUwJU4TMyUNFAVTPq0zROvlSijWVWY9QzOFypv3Yzr9CMB6MVXOFQszFyMzM
Kn7ZBGD/UkIlXhkTcjUC9g1Eo8ZAQM8oUBP16iL8FyHtt2X9MquqyXghK73eTlOV
HH4sUtqiKSwwfOU6crDMy4L4oRWt2rO3yeGc+7LfUZARX2D6uNciQeWO57Hmimi8
W/bpKTTl5M1pFmHhPMUPuCy++bSA6M24sSPWN9MEAj5Liyq6dBi/BcY2SXVh3UcH
zokzPlkvrI12uFK3Y5dhVEeQ9vMgTitfJxetRpCVOaiX0g2F7cMJCsmnA0KzUM/F
g9kWEQR4NIVFddG+Dri7675GThqxmZHrBEsiiclJPfwEMZsoHnEQq1z6x9otYdIk
o7BDoadUXaqYjlveEjfFbfBYLvxFf2FiZFJGtS9FmrM5ReVBkepjvIpeWGWKicVt
aTebBnQPcZvfgool7LT8cgCVLLksgc26teU4UUOiy6TjPAQTt+MDwlwP2ED7jtA6
VDASk0pWg7wX+0yp5eUyxbKOiPZ2iYt4emqN4zmNP2Z9xSbeG3U02xUr8KIMCuHn
d6BRnbnQit8hA/59BEHGY/AtlOGRO6l5rD+GEm9fCdML6dS+00ZImbZycsi0+nMg
9jczEtMxjf1YzTprBpii9AU7WXG0INkfVe7tyWYQNOdt7l/dJh638i5Q7bjcMRIV
dcvmlA9fP5OVY3ys01A/2wcd5u08k3fLH4ZoEWIJXP9frbtzlTG0c5/kaSSNDfSu
pYpQMsg4xjhT1mWPbTsKZul/Oyi09rhB7yEIzKCiaBu0lBAT9YjPT8lhTKmm5hFj
/9GgWRxh+6oHgJM01901kmuDA5yXAnSStJ1UV25D+cSjIDv4X+wQJxpuvYvI8KCu
flSBl5Lir7dR4bZOVnwBHJBfWM5DAkozZ4BOEdEQ0cQTpZVLFm6bBAig6yrlvqEO
hE3E9r4suUpQ3y+BZcqgHVpPUPEajLzZfz21PuZaoIIy/5lgB74zlx+t+YNCrJNT
Jpvh+2a8T2uQ5ZxmAqQr3DouIxzK9EJJ0lz6w2fM9iiTJBv8qh3SBXFsecWbEcHe
/jv/z5sjwaeHFdMK5hUs8I0ArRsFL3+fOxe64MFf0MOQ7cqtSrMyvRe++xJ5SKh8
f/lmL7PdtPl46hBoUf43HTwKspDpOwS8QBr2D1tpDxpGPWPFsvAVHVNedZ1Ru7c4
xBK3ye+e25OWHXA1lr51ZXCVanzY725RGlfwzkJjUnqnBAfvem4DcFab6V1uKa/4
C774XqK6KWqB4KryEBDVNnwcrUIIkFYNPKXKKAOCMLKkhtFqUYaoEwGUVhrJOM8m
NTtMmdrTpS/PO3PTK+62Ay4rG1HajUJpjc3FUbbHSVaXT/NbAOBQKzb1o6O/joLq
GDOaIkkK9kfM6wZctDvzoWOiPWOp3guD+aSjDWPsHL6cEccx+/6LCUuNtf+hYxXb
RdkyNjLNOkVJ6hgrUI2Kog6cgJVkLnJIKONGNnvAAmbr2+I/9d/B6g+DqomrSHeV
QxeIGpzN4sOkK3i8DguXlKzKq+XWK0W70ZW901uxRZy6nZJx5qZWjS8/DRszudnm
S67RC3C8k4fPMzLvtk1O48v+McJH96R13LgQ6fU8V9X1hOD64eq575UCKSK6M9t+
iRdeVtK+7p0/TWX7PDPI9QhgluKiHjY2X+fBGdkpOxu2NISPurOoyTponbEVyftN
T8OX6DZFqmkCoNC7yA8RBlipOIxbB8I+T5hagPk3Lloxt6ULD3pt8lsqlWSmkvbj
Rvp0ij16JIud1oOZMTQYXRxB2OXktin523faHBaaz5tFHX4PwQ2J2A/Ghgnmj/JT
321OLNodp9CSkIrYVvuaFfbBJdFd+76Wg26HJhrZ4bknnn3wdRMGGSC6lF2/yFYF
H3/NDBqhFrlTts4GWvFXMY65MVFZ8cjwh+HHiPiSAujCJopiJd3WphdabHaPuTcK
VV8vE6fv1YTbROrLazl5TcnJGmC9eIFdFIuGhH9kflNNOp3JlV3aGNWWiJVIGrr2
RZVju3c+ri56cj72ad631I4crvFa7FgV2tgksgmg4B+YRpa3b6E5NHqLFTNZ0mtr
71edJnSWRPsVtiKybSHLqcls1+nz0gkGamxjSxI2tQyJ2bSwtgoRpTW4eiXOaEY2
i/IilMZPHQWgE/MdNfjyTW52R6TVwsVDYBEPXOfZw2ZBuT+XT6yihdqXziP5KH1T
bNtfU6nolW9FrEbPMLCfD2lyU9PuysDiZ2dpO8ikjKshaC9m6R53fSdwvK2BCcJl
QiBskR7q3hMIRDfBEELqXl3Ed1vrTw9236lFL0lwJ3SvqWeSqREAhaHf9MI1BmNB
TYqyL3/ciZssJvNExhbRQ5c5GzqMmpHIRnRVPMYwFwlRupDJDxMNDF47PXoUpItH
TTH/twp4H2CWfhrkoqBSulTy30eREpy9W9cjPO8cWoAo2rUuP1CE7L6F2Pz7tNFU
wZKI6DRrgQBlkwKeoV8c9HNa3s0MWZVb0sOi/vI24bpYeN/e/LI8YsGefLEK98ZB
ex4m4KrtIAD07LvO54XVse6HHkicvfImH6gyG0PTBbpNofs473W3jWYy+ApUrndB
+2aWXY0m7J2qmeDN6/k2AdkSOdwrOPItzgaLZNk0oTAaK0pZk2CYJHk5XJWrn99x
L9sgvEmCm6BxFJeaGcWXBCN3Bi9geSlQYu7LfHFyGC1tnvVtJ5ABOwOn+79KrBeD
/JUWZj3uF7RWowlO3bvrk7YuXP79lvC+RUX8LFGcsyB+LMKJ9fdfFSQntLX8FaVf
18WTIlY/5VhwGmel6GWcfo6C0g9rAsrAbXQtQQ0HjtHGua1fxUo7+WWMGLeRqYQY
e41o/bgOj+RxqV66gHM0UoYUNp0NOK3izyounRNASjrXzfKcZsMYpa526ztyC6Ab
8FzI1EMgdV5lvetlLafZnhgK7UJZgXw2nmLDrj4KBveCPi9FA+M9BHbk6+Nt1d48
9m00I3AqxrprhW1i4Vf+9mhqEPA9/DAo+Hhl33+9iRYahNEpwB+LRgrdr5WpbRL6
xz1G7UQuLmGkoZh+TWyOcf4YrX84K6mIK5JIJ7L0R4TBR7rDY1CaS6LPbJdxmtOU
hXorUbiMMHKylHLMao9fdPusnbdp0ciWUAxHHkPgt3A+ZEIr+MEfN9ydngWX8Waz
BQ8r6i83LSx+O+DIkmi6Z1Q8jVT7dpB51NJA3+tWR6BkD6q8uCSAIy5ro+5qN6ea
cpjIaSUGbmQjVvmQUBXVBhLOp8anojmWoPhhglm4w4CecKDX7HuTu/+RH3mgzEYH
Q2OSY1U7Cy5Bj//5AXrb9tKM3A7xlKCjWoGzXsLrWgJ937qzuhNIyChaDIPQyCvI
kuQjveMHvT9PYlaZqWViDjXzAi1WU5g6Y0R5X44AVNtiQHyUr4/8FG8vpWNBEpW5
l1MMJGHF8L16F0Nbhr27UoxrDwzHpZP+YiZV2HP6Y8r6NfJvLUa90Jj24pK2CmHk
zltjkasVOxr3smUpsgOw70sb5Y8+OLsxyafVmXpgxmQq+556ly9VAP9kxStPdqmf
oFCpIYRpMEiiqH2p84pFIsf2XEcwzjyI7EncRkg3umCPVXqxlFrCwRdjhx9RUcNb
tShOoJ4L8ysG7LXPghUTHau73Z+xQys/GrpJzycY0zqYZIm9Xo88rO/C9nzkXAZM
PhNaG1wvnyasfklwTaAzNnhsvY7FVeNEwx2dYU3EfdCh683666ZWG6waVXzSIRlh
ngx74ANE3SbFR0ezZlNgxxhMc3qQ0aoY6oq8MBoPsG2tC9jswAI2kmAbrmNnLESB
6ODX2JVNuD9oEU43oqtCBSPSAboTaQ7sN+f1kCsLKnXUKlwooTRuBxlGtySZnIWE
fbw67AM7m1JfIBISr+/hB8uwcx/zeT3RW6agf7RenHkGFuPD71ICqUdn36BNHogF
N7DlSYZWDkF//3XmYV3cE69QeiOzK/3/rZsl8iPAdu5LP9/orccL8ChJo8+hQ6OO
s+GX0KGMEqMCpNynv2l92ED1eekyd93JyOvEh0iVfN9sa6txevvbffKPmGoiGD27
raUqHnWtfWRG9t2gspTn9X7vjlbwvSnrn2Jf56Cm58YVy+B21w4wuX+z/lgv6e27
wqMiIXSoP09MfFkLx12LmqBgf5CuwnNLDFJyuaHCaHIrIRqyTtb1IIcdEOsvA+td
yLOZjXS4JtXrmaPsFG17lkerhzmcn7guwqmI5LLCjgwSHCnYOm8IYcLhLHv9yCVM
HmVle90qBobJKyZJ/wm7gkOl6XbijQwa9x0rDzfDWaK6HLiUnvSomh/IE3j4iBrL
UhwwtKSZGSpuu0SV8KIV9bKDTEOptZ8HbZY0Qhd/TKU4NGFlyoHsN734u5OrSI8K
McpcoK7JghRHIc8JI2kkmzgqraU9a1Tc8wDX7iTh7NicfI9PhtVdi2arSnVu7AXX
xHx3VYhYZrGmRuTyfaBEH58TLibh8TI+ibgQ0szKF3tKFbAQJtapOy2ppE6YyN1T
z0ZfAvSq/B361fvO3JrRUCvB7C8WKOvHVTiTRm+rmw+2ZXBMENcXYa8MCkadNs1k
DHHTLYeSsBhWUPYCR/qX1ebjN/uRxjyjGdvynXVXumO2snNaLDX9YUYEsMgKJ0K7
Ku9QB/HSVbsSFd1Z+yJ0UYMz+tNFwfeOn0GOF8NgmWKo+cgO6OSgrOvVaZZrh/ip
Hu0q7muLV0v8sduu99ieaPbsxkA8ekOJo+VQ4/voiyoR8zpX3ViYCLfC389Sn/Qv
oBgb2iCKKxtn7mO6bDnlskfyBrOOXGt9113ZyODw622R7DHQoXOXd4+rYHvzIlBa
AQ19hQUZDOM79WfJsEuSSm5QwOG4hM147p1ZpvCCVur9saPlXvhutF5RGktdPZAl
g2ygMuyjqtfQP6Q9GnGNaaRftljfyz0oh1kuSObNdmt1HF3yp2O58NJpfsHgeak3
53kdqXni6mfmgu2DHVXd8+eeb+9pB6b8rmNGX56D6TiSn4rFIOetXF+bZ9kG0viq
5BY4ci4+bdgBBteJ0WeLO8XFGo5hVldUktqCn/4nV2SFxpIfeiBnOUOaJPpaKCp/
Xt1bMDGFrXWs8J9E2Ryj7LUqx/ROoKYh+EAi63Dh54+E1d3dCQ7jkvUaKgfnzrCf
S3/6Q3SY4pmhFHDoLEDFbZNg2aacLAokUpCckifoc2UtaHZhrpMN8hlUaSYUxLrq
ol9egE5cdwrV1JfJhyPQlXNUlAxh5AKe6VeVIjV5fIss5hhFBGKcTOT2NfRBKNLa
4vJ8qWsgxJcd2pIv0KWkLsnwDHwW1wJcQFdGD3H+ehJBpudtwi2MziVSm2oYip0A
5S49qiZh+qrb/OsLFKJG1xo2QPBrFG/oZYLouZ807qgj5tv1wEiP4pIZ7/NzmroJ
HVDa7i5U4JJUSdQ6chNgT/SLNmj2+tQn71t6dtlE3v6PwSwVUqnut/mSg6oQXUve
nLOIQftM8Zd4B8XW28ihwHnDrIx4pqg8XBGCerIddHVKon+Zyh7/VaKeImvQHl6T
114arBaHn58/SNJQTZtQOhyFNdJl/MvVj3kdRT4qhmuXP5UQ/tIImCVTzmreuKXF
L6lFsZkclmHovjxdKpX2WjHNfrRwfTr251fTcSadXMCqdmdps4lZLmUSa7bbh5qu
U10C3HgSMb2D96vrDqNkagdTXz3Cw6kI+omn5c2OCQFRdwejcjaoLV/TgHBL1lXw
KKVvkVj/i/ZHo6CuwvyC4avJaNrxuaTvIFoT+p8a2prrTZzNc4HP4cw4p8GeBjWu
H0d5krj0PGHko07a6VrfTHaOp0NIuQ+q5N+3WQjYg3RYdZaaYc4zBxV0Hf8shNC9
1PT/bg3mTFXA8+rhW5dvNgNlfrwRx6h7KfD+EMDmiRtdTp6bLfA1yI1MdUGNB0Cu
AUIdGVz8exPN/mxy72hbocZFQUSydFs2TzUwLa7EPOkslLNw/YgfnLdscQcUQkn2
SSxC80r1wXxy1mIrgfFM05vw+CgY0JIC5AIOqNsZ98Yf14801RGszzNxPvRyqqqp
NC0J6K2SI2qa7xqG9SaZWl2VFccXta2BYyqvWHXPOH9hxIg642f5rqLkAmxWNnwZ
T7Xb3WmMNDDPIpT/BWkJWMiIsMtzUQ9szWwM3y4gufR1bwUBNEwsRkx8eao3gkAz
VzDgnSgBkDAPiwfRcRGPgvopAEZ2MmnYZhjbeyyFODajJy/lQKJuF12g2YfWZWjU
u6B8o8TAqUu83yAgN87rKqfIGoPcyUHvVBsMVKZ2nzVrlkKSl9Lq0rgBYTEQqZJn
HE6yOvNj81Mv/kCESxcWILQwwOiceFP/LwvKQOpBbeVHlhgG2MAuy8k5MBYIjStb
s6HaFOkAneVNnyja9l+4nFCvt3rQqNEyYekARLRgdXNqvtgVm1hJcoWupMeZLXjY
iBkn9meIfdQHKB3vFsHkTpjnatF7qn+UVnZ8ruWzr3RiVmwKepFX+EJUTlyrWGz0
o+e3oAAT0nl0mHfPV/naxS1DCdVkiusl5EJXLL1fqFI5cmaKBxHYH0wc2nifExMQ
v31FIGEzXv3GNvmSAUaCN3//hr7lU4buCm3RW1NkCfj53VbIWXU7Us9Ktfvlg7jb
avTZYrihLsFKB3E+1dfm7dcHQCzP6+b4sET3xFd8s1bAPWo5chcV/2+bK1qT2P5X
vmqY1rWuqig7FudfavD05eKfgiyjy8M2XepoDDsejQ5aZYiqQ99uM3YGXRhUdl6e
Iy0iNrWsTrYHK1HAvmM6PxZ0s4CDTZaE8A/PV+p1KEdBN/KGuDy6phVeJXvjeJTe
qgN47ZX96bkW6j/lTSlF1THzcchsrQNGPX5usVKpVXN9TDYIcdDETN07ZuJPPh0e
zOyVjbloA6eGHiVnwiM6vEw4Hz+ELD52kdkUSv1UC2CXC0xBWwNlLsgn8PDQQSJJ
ZngN94crklxz8qYjg5wEaQ1NLJKDv6Kn4lEhlgGo+nxcODdUnoFdG+AOV5Y9KTXL
X5zv/i+b/ZBl6OoG+6i6SAS1l18zedze8XY4Khm0ZTyhLoEebMoO7I+ahLi/jwgt
/al6K362Pgmgipx8wGJ3lkXB5plUbgCvtmcmVw4nCrTIAQ5JjXsYTTU9rJjMy7Gh
6XXv6foomC1XXv5sZIm+vIF4vo1Yp9CUz3yWU0gkIDBZAlEVdVCkkV+OC+QMWfeN
/6xBIXKIUJiAwM3Awb1Ncy25xLzK0UvW8aHhkbkaKvBw3D2ioHl6kKEsMR0tWn21
5N4YFhe9127kotY5l/gS8fac12jp8EkWdAQr7RQIpKQ+g6GEj2SXKC4V0XUG5tjc
j3q/S3qkIzXIyepVdlC1GkUuk8/v3VddA3OB990QepW5+s3ISURZcUD7Ob2esIZu
aheICYAL7tHdA0qQ9WkbqMPFnVbeslgBK6DScIGQaeegX1Jg+knm9ttg8+TYA+xG
b3Gh0yc9onbrwEHRAWNQBBIoKHoYRUQndM8a6ey0WBBdpZsCWjXoGrAIsAb9UrdZ
biYE5Cr2kXMEU6VB0K6ALySAiyvVHgct7YsjnrKJ3SiJxeuDAiGOvdNfZmyu/5V+
RSyi2L77Ox1hYg505Qdq69xFsI/su0eSaJ+ucljOJ2MqZpOms5/zdCtpqeqkj3Jc
NU7jnlQC7/Q0YBuqGD/q4GsxRL0Blrb8pNrt5lcdz8HcfJdKkMRA1Dbhy53MKiD5
sqjmkt8tZ0lxCWe9Alm7iOPKiQL5zg/3tzS2iktUjTUFpAtFmW4gPy1PQ0Kv7vnN
c5rU2/7Vw6i5HtcWCCqPnbFjn6eAAsmdTROYJxAzMmWeIVvqw02bAY2MUiieIqwh
LBAbgieHOShkaqk1eL0a/s5AFK5WqpPvJnDmUshBLOjX7svvW+vOSiEGuaRKNhF6
Ua0CVDEuZ7pwg2Avx6AxAarl3QHG9Y2KxrFRzsiz7NzearkrK3hB3dh0kwOId/l7
I3ObgaGlvjy0FsICdcwgDZTO8ghGGf9TQ6FCjrFtRvhdFJxPHQ0rQgdckHCpabys
CNjie3oX7ckrs2BvpKv5+ktAwjTPVTL4PT8G4dtCFsclYjB7ujRvIlRm4OgKLYkn
XR0PTxbXbExBhaZMU78ICyqa+FBrP0CMAOISsBiNA5IKN5d8zw4lhLf/0uSofdDm
w0MZ+LWRNzvgXBOdZsPg8xDegyVdxsui52zFkztonZ9iQd7PTbPrZYcAEnDYaV1H
aAFGLhiSzNlKZdTlMxop30al0qMD5VEusXE4C61n9YSOrnNd6zYt7aLkOG8IjRNH
X4wg2GJ9hpRHGtIg1AydHe0sbITa6IRlwKwRt1sERl8hXRmq7mikB3pgZFgLElu0
p7M2RLNxsAmdElBgyhj/l8XV+do1rio27bmjiGOOiskvbzxISv+twpk3UccgUZgT
L+/a/OuEP9H/PKEVUrR80lKCxj5voyr70Gk5VRr7nVGYDgdpQsm5SjILjkpBBlaU
sp+1UdK4pdFLWJFsewrW+iN8lOmolnAqryd+VCDoZmEBqHEeWf+ayEhAepaicwpV
pM6O7to2RqQmVvI2AUJ54qcJ7Q315OPrVLFilpAFP+bKeUwJ6IXVr/o/j9AnGZGQ
keRuCYMtzMKReKfJ5Cx8EJMLN7IBs6K6Ee//MDaGNz2s0wyE0NKpTfyPiOcyvrUy
foEZ2j3Ls+LTFVGPUmUtL7FM2aZacw6ucBXlYykdJkngFz0MA9aRKqSbDBOkyouD
VrjmAaoIoyZnto8yHh6vSpY14v4+54QPcM7CeQa0wPo8eZWvuxvReUIsP7boNphI
mhXbAPJUsf8ejPlyE/T8LlaIvUbFgFKVhCs+ZuNKtTaEzN7FqfHH9d10o7F2Tli1
KEDGEJZ+TVZ61KtjP1u0zvVBCs7kYXubs+ITpYtizQAOHcnHQC8rJFykdNCRJQIM
4WHt8Vv3aARlHDk0BzZ6EFg9lIMtOLeI8SFdnI70BAmWgHtvTCsfnr/81Ahx11CI
/3S0ArVGBJ4y0mPQ5FlJ0txhNB/HTZtikqEi522rApoK87hsNlxf9LRHFXX3MO31
194v5447d+Quf8FfrNLJFkdJ3WAcl64sw7+2jIkxH1nZQREmxyCQoJFYN90zccM3
vItVICv6l+JOigiNBTGK3/lLVmfgKAiwW89pY3XJCdjGvIyi07zRMxTwMfaPvotL
ZPTSlEaYRYxQQo8WV3tuilrSo3avSgK62Fr9IUbwmPjxh19EZdhRTGO1VQ5cPq65
nbx6lyiIpdri6/WdTO9lPLG0GWPHf7fFj9i1XJFa5+qaArEInI08cdbZo0JuC6Nf
Ih+hQOXQBZ5wJ4GWm2YIJc+5+cex9XeLOYzdlsXhvK5IPj0xfAL2IUhx9Onm1vxy
8mhPzxZLtmXgZcJzVYb/PPctJj7j2m/tMAIalfU0H38JfTm1fWQR5UoFPVPAL2ZV
JLiog82UE0+Hg4vfmvK1WaX5bSdV4qFeG1+6ORzFl5NaQJX+mPbkykYuSUpMMvPR
Z3sZBEcpxDRpXgRu8/KyR4vSerTqNcdzTOV30Y6WWZdaQLR4ZDIo7jQJJa9gSCFq
S92MQM64c37U2OBtXarE5XdWyNlECiCaAdBUBvG5A+i4lz4F3UjFSvpB9y+7/nEv
QZlUzzqZYt6kJwRdOCdW4mDgCgE7C15Ra6Fkqbit/RYN+ic+O0ugd3vCpomQJxEZ
grz3slCTQsRO2QkY6sjls57PPLpbCM7xgxY0MJXPef816N7OWwEBi2QBlYE8OrPl
iAkvm/4YU3iP+Kos44/tSCzQlypNRYVQrBGH9YlB0Vek88Dl6JyWPXIGDlM4aqBn
yAd78F9QcntQIyWXsSFR6eOzF7/+lYT24cChmNGpD8Cm+uP8vd6eLyY1nVX/xbg7
wo+aD5nI+qqewApFJM+Nezm3cRxAHGLCs4ThON9uY8Cbm/aZ0NpqmAPYRAroWcno
Q2XBppXadxrmCLuGZKeOaupBX6+E14OfaWDoUq54WHSfE1bv4PthpbEqf/khqj+M
LUIgzOaKjaMxXMuu1tnbkkF7ffHYXu3plJAdtDmDz1C2fbIL7jOA8/ZbKx1mu5Cm
rY0++lpKQZsguD6Y3KO8zHAYfYeciQjWe4yn0XOjEJZhFAQfi4uNOYkqshcUm4H5
w5AWq/wIjx/Ok8JPIEo8Vfc9OhQeAv11BBsIQrk6pjEUskPiLqNM1dhM+K65Vj22
rLJQSrQPp8vLd/dpBiiacSEfDL8/VUINadwYeULsdg521kF4u6N6KiZ2+jMXxlhg
/vQVnc58588NjHwzwuALaWASk9Bmp9gFCu27MRy/hUBTYhtkto/8RLvQ5uAio0eV
K5OzFNO629REbvzggTzGxubHhINLJHXs0faOVfS4dySh04aVfxadB4TzSYTh+cYM
IKGa+yq48ngbep6OHJRZmpS2BL/tQc4eRdzti61zHd5yMKFvSMDLuqIclzGCt9/X
juFBREmBova/wp5zSVN6MH0guZ8+lDqMdofvH6fApiYCBC2dlwLZXPPQv5E1+AF8
xM9Lxsn7Fqz4zALBFl2geZfaLmpAhnWQLM026ukoGfKG1t+4+prrgWd/yPx2I3NN
as9HWDD1yGCEtFKWlW3P6jeo9iXkrsHsXXA6JgW7M9xNWG5C7nXVxHe81WPuxkZC
wrFr3OiyrgbhtYQAQFd+Zs3FBOBCjjr5IvbPgGuDQTodS+Dp49j/aYHoI3doh9YQ
Y6zQEm4OMNTL3+LKFmtT4LHQc+T6UaB6gIMDlDqYd3IkcDv8ZbXaf4lE/XE0DZdo
s6dHHBBKOKOnP4EoX85akS4WOrSQWqlKLLMbkbT+7Lb5Re1J+Lsrw9MYQwTB2ohV
7+zh3ut2vCNXD/L8VbklX53anlBnqSy3yys+Zox80JMBNeVk4wt2VtQbWdvmGkdT
q9enaPXH4eFNpyc/E61y3gAubVRC03xdWcjxUSiAH6ldFYYKNqGJyzpEo5F2dwcg
w+N8C//YwYWN9T148NUxX9e4WIT7if1k+67BcxXj5qize22JRq/jrij3548UzrxT
AmRzRV7wsjHcDwZGaPl5lFqUlC50xJQ58YcM4LY8jeH2j32GKW6zW+uY39auaZcw
0VY8yKshbZ08IEIkVv6nHv+atgKeWAKTIcPOshWKjJ0XO2YUl/z1vgCo6Y6bkxdR
LSDGqhxSjsy7oAnKaMvoK6LtqY0a9uBcR1bP+YO9YuGF9ax3I2xtvpLhzgDjcCbe
uWM+o6nM8aPt5c49WoD0JrE4rNJeAS72faeKPt9cW69GWmseyXpYlkTjfOvk7QuE
lS12FAs32HTKkwiD1gWqLZYihWZFQJ39RhM2VJz7eAs3fTb3+w0Wu2axzM5Cqxgi
gK4YdF4grtUg0X7MyqJOOQayx5eTau45jQL8xvwxI5ghplS79l3WLydJ+op2/K9A
+IntgCvjkJ/GulQL1JVSVDCciZU0k+gEzqTiR6ioJX34wqD71aKLs3XSeWIgRy0T
UFQ+cPKUSkRteugmYAgKaACOkCspgdRrVImWf9qgx+1l74SrWuUAWzUYFbDGe1sa
JFkn4uHBrB2ZnoFTbKX6R60HIsZhQO0jRLPFQ1ey+KYIO08Adn0EbtthTSJGs1cR
10F4QJuKZm5mNOE4OjkwCKC76c5VBDVlXqgmv8f1jma7VtemJ40KOrtaLTQHm7Es
u0/4SjdeymJbAu2Rj556LZ+YhvsnAktfmoRlUeeklKF3qHy8ATz+CIxOlRHmIQY4
2tmaoOldy84lTvoL47IpnVFxP8NaPbRusvMF4Ysw9lN/4rMj84OiC3h/gPLbkh9o
gLTXVYbReDTfgAQtQh8KONtoE2wpDQTVW82OAsFEtQq4zdpX13Fp7oJvrrV4Am8X
ZTDjYx74oNj8VzAFbngOGqOVWl0ARP7vBMjmJoRFhWpr0lfpPBIXr5p4hvhQ+vJn
H+mVx22rM1rIJUObAO2yQE5GloGAFeYjN2OyrzxcVOrXrrTXIeL2Dx1jPrNg3rPF
l0wfKyreB9bJtV8ZWYMM9Zu0qZ9lQ+aMtWMAJ71MZeD4FZj4RzIp7K7JaCM2tVTo
RUY+On2Mg1P5N3uKXtZF4UOhhjffajaR5ctSA7LUQNkvdm2NuTmAQS3Inio5CEXy
lT5TePjw43Wdp3M2AgwKhsP7mTq5NwGmoAZPOa/DHKhNzIrPrAWAgID8HGrIaLP1
a2sb8FvFzdR3SYIgSpruGBDAxcW7TNn4oMBQzc977w+PkWmyHZ4nAx0+5yJmdNet
eArmkJwk5mQj5KfqIkQa0TuQbu9co7V9/XZlWJCOcgBcTpsUSIhCL5RK8av+OAdY
mS4p+lfNDAwSn/yjxZhbv34lhATZZONsV7OEblk77zRm+gtW8U485dttU1sE1EMo
FayX/5Cm0vjm1eZugeqHVUlP4BhEfgAzuGNJxVYoA9mgOagS3qy8rXJ5B0I2+Gac
qRJERt32dEysh1ZJ25b/OLxWaoDsDHDSmVdUmDZ+jfpWJ8vpGM33YHcRsL4qnC68
q+8rh9C7IgZevwBKpBanpYc3qyn98vVEt9hooKSaJN1Xl/AkkyTe9GQJAFF7rhX+
Xa/riQSOT8F0hnM+sM3cFsTL8dsZy2yQbJkA8N6YuIzo1n6N+aI4mLz7mgDl8BGq
fNLgIZmwdAgPxmU8e1nHClxsEng+PZ5P81oWtB/xCdpfFcND/pCRdjswFW72xb1r
Q5p7hOXUG7InLEsa0azGq8igY6/6VNFBqJR+mOe8hTB1uIdFuf+4vzKVao5yzEsD
LDarCL+NQFqZ03Ri9zS0fjxLp3I2AhRxpeWrvMoWIJ2s60Vn3NPih1Hhq4iez5kY
XEngPN0F3xU2ufSnZ7S0x0eM6czMT9P5f5LR/lQ6AT8+XVXK0SgSdKIwH+qiPFLF
lWcYk5xeSs3ucQs41Sljk+2H5MbF353HMdoYjQFBakKsVn7VIgzVyN14YWCS9nZ5
xBBfI4vVHqo0G3xFkyFjJ9ZE+TM/kTi8cp7ng+w7JzFMoeoSus2N2IF/iygrjl/I
nduAhTGIGG25l4kn7nZWRSH8VZR+fgmMd2Ql560QVWm41LAwmUnUkBL9wTntoejg
CDEa8FnkdjcJdELm1uyaU9y8N9YCGqNcEiaY+ku5oZft0jccZCZ5c/lTOJWm2G9U
bTp2eJAsffgmczhPLfhZdnRPfc2AqOnrL66aJLRhkSG14ynd9ORxj9f9H3mj1I7y
tCJN/Q0KK2zQXYbEG/QwE4UvidFfrevs/W9fibgh5FTUrQ8c4wNtjQ3+7kAnXfVH
HARxlc1cCzGi/Dk3iF3XmSHHU89ulodAYTYjtrisgmxPYhp4HPknp+Wn7Kup6a1i
DOhp3TRekmW5hngii6aTXVU78zBge6fAu5yeAMlcVxrnYvRVSrkxRB/Qde25uywQ
vfMLEKDDEmge5rtUevpf87AddnxDGKonuhEgRFRL4eK2HwWLaQVV8LA3rFQxbmmP
xuSMnAOcwz6xC4f+Er4G17H46+AuotctNrvAf6v4FXgm4pIgu0HqMuoq4MNO8Iff
LY+o3hw0RKipCvnMbIKbQwmbEG2zjUA6ZnMvA1q+0DH4Cy4qkN4cr9+mRkhKHCWm
4MtM2k/lG7erYtSOUC2MyQBvQQ9GrQUuDyKVj9jWxmWxMI0b875z58fLnDz0QCPo
q2dAX1e2okMM3f1tLclYtfaRYmHjxTSgo9MXY+p3D073YiRXEIP0gZlkXR8JIVR2
Cdz929xlrnWF4tqDHvWoLA+GQ76m3uKkJu/x0FQ2MCth6wH5me2ZuASVt1DK1VJD
Aq1QGxhq9KFnVr+U+8LxoOulFxsEV9QHokY627tTdugTKNXdPhLsH0ji9qvCg48O
vwAQpI35iJ6qj1BO9otXcWbejZuv3P2N3AI/FJZzvbK9UaURnXLjPLFHZb0rXNIt
N4VGgDdln2MgEmBCjQZTmOxHZfGGHh0QsxgiROlIU1Aiv0q5rWxCaMEaatccd+rp
2U+3WN9n+mM3wvbmqpvO7jnMV8/8ZFaxgG2H5U22yNGowvgKkC8oZviPddGJbKRn
FYSK7NBxggSr3Mf3FhiHNfcv/02XmfAgMl+T/AlmPtNQJ1vzuXcPiVGMXplf54ny
wx3Gb/TF/KOPf+2p1mwluxr/fOSXie3tXzK4zRQqDytPFy7d23zfB9b62rjYFTna
FrI1oMxlHAJWh12Cp0ExfcPJuweFs6qXMgJutkF1hMnLG+CmdKgzaCBO6jo1w00k
8fHZgMq6rCBLoW2PnAPC/RGyGfgk+pw4oYsScQiCvwL41+ecuK19i66KEBcqV+91
FAm30KN4WZC0l2PIFRS2abtpb8LneOGC2G3r2sYdKMJE9nE/OTELvRRYt7/WzK/k
LMPlhPGbHOWheL3yYaXbeJFTX54hIDIkIire5P05445BhQCSPf44aNhFZWctCOD9
IaaiYkeDwANNnCiObphR5bEyxPr095dW7cEDG9QbAwz26tvd2dxE/WhsU9CBgzEL
m7gQyzrbcfOTfdcn2fA9d9nyxR45nSY2pSAnKQ/2Df9GURsnepttMokIR82oRHoQ
38CpC6HtVVZ1BKmNJM+19YzZAkUyIuC0DL+GSmLEvvZy98xcYrujLGfVtX39K6uV
CLjaUhzJ9Yq6EknSAvBZVj4SMKL/LBf9mbhHjXbcl8HLiNG4MxeR9zZeoynsnU+/
+/hT6fAZuei2ptRxyaeFG1dg77tHByXBPFrUjz5KeBHoYo2mj3dCacMp4M9AHb3y
9JYxN7JI37C02qRBTaOt54VcYVk1qBsfml1wrz8NlyMMKZjYpls8WneWNcqezW8D
SMwtgzviz89FU/HZG/w6skgsAKK0HMrN3qe6xKlWnazAGj2bbcUZJ0LnTRXTGghg
q3Wc5Unj42IQ0YW+VK2RKJVuvrzQcXa5Ajf47Nr6zZs8SgJTQE6MOE/sBBEaucv8
5T8Z8KOs+gwzGDLuH7LQndnesfq0FcEWM67DN9PVEqd6eT3aPkHeSaTTCpsqJ4G2
9AgNFtYlERpTmtvVrEqypS8WeX3stz0WsepToSrI7ui6e0ZRqz/O7zlG2dQ90u+D
1fyNL+ut8gmmDUD32mTpp205xM2Ys1ul4Ds3xbkC65FqA4X7jVm5ddVDs6taLohe
/7uEennAc8lIR5Yo8yjRvRwt2TtH25ugSB9JOcWEtRolG91xdTgeLvnhFMXxWSci
vqHG1kid09PqAAToMuO0h0Bj2yUll98nwb45vmSLrn+cQ3binaT44kG+826xvLST
/etNdmFuxv7hDAirxDvTUaBg9OzmK0RTBNlqPzShgm3F5Pq29iQv9NkA+pJgeaAm
+lcEjrL2OW8kn8rsIqNmAESBp9u/wMBRT6yb0alyXtR36z+ThsAYiwjKtt6dRVVi
+yeZ8oEFiFv6c9QFg3489v2ASq3ix+RBQrmsBeHPiRM2D5fi4KxKutRL07IKMb+K
g2t3bXKsP+utYbngqmw454Gro8gtNjjgH88EWvq/oBC4rhYGotNekqPxeLM7EEYV
qd/r7FGClB1klRuvqBGP+80VI8G1PfeiRQw7xekk9A5IZL8huYMDUty9IZphlxGK
FksWu5vYkejmVRqYqPVbvj5y2qFYf+JxFdiIaUIyoXP9dk35kyhnmH1Avt3aMdS+
0kfXGLZ1P6Y8dlvrJ3gXqodrEDu6rJ9dx/W4gPJuWgXgWtbobfGWULGDyDyg/t7Y
BVaQmzUHdJE+JxpUUuZCz3kF65uZFEnIaAQUNQ694Lhh3UNX1tbveTwl5iZcehmu
Crc6J+khr9O3fliC7KW7R+zly2X+rhhYYRjUqZokVdCl+ukzkDmH/Tt3zWPCxOVA
qiE6NJPgYI+0vrEsKtGkTsv8pQvZVFR4Zvc8PWvCvpJXww7tGWL4Ul914alhAK2f
G+cdYbwzl/n4N1KoK4AkfcuQuKXS774/gFNa5574YPxJdOQRBo84SverY28HgQ7k
ySLBIYUCnMY1tJMfsVFUJmSgzyJ8SVmlQIW5PTuqnk31lRTzkXQRVTzVnt0ySJ8i
WZeyorU27LpDaMJbsMdSJqiv4QnkllDPQH5onPv8UR3Oeq8aByyQ/4nKObsNDqF0
OMC81FC/ztB8k/nIDwEOp22xSg5ydM9Awt3QHiY18zpThA6yWVU/GyDHMvbXx2bN
WJnCNd6MXyPPYstQhRyLc8TYkBqZInfSpA2YqlU+7CeSuDc/Ba0/mw9S0w/ffbnC
36sCOSB/4xrk40q7wqEmxxv2g3iurrv2a5AqHx2SaYVwfr5GSaUHIYQjBM6Ee6l/
Yb2EbzJen9/Jg5LpQEE1489Dg7ARMdOgnwLKZk8gwxx8tv01rpSWibaHZ8p8wcUO
Han13zCBB/CX+T4LahQQdJeZqlSvq4kwZYEywSdX7jO2xvtzW8PpK4WHwyWiwhsb
WPLBk4lqkVf2c7QZa9x8S5yiwlRYFdNhXmBANHbEfUfd93Ztf/Yq0kq5F3/6jvEB
TdDOn99+BnT4DOv5DfA0AjcCXkQ8lsm433a9LUbqbo3KpTPw4lGZRVBv6SPjZr8y
R2jKlVF2U0TXHBt7nfevtwgoSyocUKxePq8b39ngZduXHTZleBgZJfaN8rde01x4
zYARgspNh4VxVLu2tky1I52akSuwkW64CDSQgcfEzJy9vnPkhgAAghYRCKNsbqYi
e7H38T+PHeJY/MR4FY0QHM6syjOdXHJDo6iAdSPE959vx82Bd9LM9MMwxA3SOyeo
q+32/a+2JApGnr02EfzUwTCpvDvMeF06FFoFj2PpQpB8GmW+oKf3vgQSnPNvkTs2
rSskWsSM615e4wm+6A4O+Vpee1yuhpaYnpYs1rbuR+qb/IVkfnhXWtBh6OZLGB7t
2uB4BvUQUA3mmDeygZgD29g/m342uBC+dFd1TFoUIYsUzIREi/s78X56L9LAZY0u
IrwMYh6eVp5lrs+BqMsEzKB1EleDU5pXqJaRxUE7iM4h8oWh1EO4vuRbAalL5PbX
KZeOyo8Z35p6gBUXZK8+X0GHbIiLiiXB+UvGA3di3F12KVkcs4zleIUB8J/PurlM
f68sUFbGcL0zOUuklW+Aw2FW9vWF3UnXonc30uMZspoNa/oiyJdOj+a6NrNDGAEt
2U26wkwjkusX7ehFwppl06hHjTcjXkX9wuInNdfolN6B0ChOzXSam8qqrO/7ddvr
BIY+s70jeuCadfL1RQ+c/sJm9XdC+pLGjTGDg8snbkqoRXxb3erbb/D9C4L7ge71
vuXDFOe3iU2I/O8FPNjdL3/nlcromDA99UE8r7ot0EbIrmtfPpi6G5Ox2U90ONne
ko1owjcWZPK7f42MVjheC9RqhusSFZqKP4VtR+gHDJyFWQGg82M6GE6kEOJeJhfu
aKw+qzuhpHD2mba3k8BQiFYqM6uYB9HWoU8OCd0Lc74ffHKp3I3bht9PcdRAapt3
T+ofhfyxmSyiG/WwUtLEm2U5onwtFW/hTfizjvhJIbZb4ydcVe5+sbH36PudRoCE
q9/3hwKtqq1JMN7XN0vVe7pN64jQuFM+AUfOxG345oW5FJ88k6IUW8/Z8Ihth22R
cwU+1Us0Qj/hylt0VpcbtRaJst80yjz07hrVM7KkKQ43oLp9xk1EYdbz1n9yyre+
UCEgrfqnuKj7r/84VG4RIdQcxAZB4IT5A2bqCtcBFQRKXX1BBjwJAQCp6TpgseRB
av+Ad/nW2T5oMpSD4Y34K7EOphFcFsvsuE21dPsC3lj7xSJlAvXpy1+dyuVGwdDH
kKW/caKTjJcTmFNoXKiwb2WI4Yt92WLGe6w9JN6uq0nkLgW317X4V+DrChl0W69X
Fpm/Xwj920nBOG+wGilH3AzWj95z1kEARKp4fyu5l/cl/VreSiam+hhcvxmt053w
7lVFZhKo1VgQiuq+cPA5DObNSpNPzpNJUUe7BTIB30YxKIWAFStpCvbfqiAG0jVn
361QTEcGSWFt+Q3Znr/9rEZGEIOibP1eXzrmSRqZJ2EWygjTdH6SMTPolQYtu9xO
sbDmEnUbvqsEsX4esf1BTCerFeCatOWlx9SO5XlRfn2Ovkltu72wJ9Scd34cKeBf
p3q08D0dp2n6VdcDY4PUtXwoD9qbGoSZTyUbwdqur0q856TUlOEoE6Fm65+1hbU6
CehlG0wk105J5VoYM3XwLN6rXgOx/2j+x7MkOaDKnBUXwgk6exr50R/eiWiXb/tL
NNwzopgrpp5k1SI07oshY57xsW/9bjsM69QQ1T6eyQzfWXo0/eLeKK0/CzJHRIFz
DGlejEEJ6sFrZ/tum7SKgeVuTvri8oUBXPBUYjmMzBo6xGgNqJmFJdbaiD6whfdp
NNx8YXB53N1zeyjSfYXhe1mHEIMALzToZe+oMMzv0PZa+etnznK3S7dHa5PGddGS
xMJiWK9bUelfOZEeXerQthzoJ1h66VRJs8AjE1L7NGoD5/kLwGI7s1pYeLzMUFAR
eEnTYekSSyEazRLE/byzQgT5EopVNjAHSn+ixAbCaIiuoaUBik373sVZS4HCwARN
1hQvDDcjr2iqTKW0bblUe8vCT+m4JLguolPDFA30ssDAAx4/5iJ447xoAR6ovc17
P2wYBd6mQ2iFNmh9Ux3qitVDbKVDt/wrelJS4IlcG6qtyW+SVHaqSwKaHwqysDzA
COYEkrUFITgTKQrLOPWHGOMXnGzqxmFIk+ATHh5Cd6xNgdUnv5tj58ghDeX9l6EJ
ZtDMjHusnvi0d3DWrZZ/YOPkwzWZR8OR8kf/1fy/pmuCZ+WRkjbxixc7rpH0MR9p
+eUOEqDEfcKp7Ctrufak7uUcRW4OXO0NCQq66QMa9oT8Sf50SAgMma1KeIIHT8VE
XLOcuf31Q0t8cjFav6BIb8y81FRpdIp7Y6YYTc+5O1yVzL42BGojmZEWdITsZhT/
hc1Oh6PIhJoXbRadqT+9kqJ5+gEty61NfA6eiXUO+JDquihZAWvWDeiDzDF0ITZR
+hC5FSmnj/54hox47xDAZe5s2pUXYiuTvFwSxpAWnNtIZsO5NNgTSLVXAXO/rbnc
Yxeecsyf51Qry9LWVHRas9sjxESKkzWjnCZAM6oL3dQm/Bxw8Rj5SSjImUVLnCVn
XZxZFbOKSjKiNjia6/yECPnr9M6QSiNYNu2CY4b8wII4tHjJem0U1FGQh7lH4k1n
bfGarFBDHDHMoUYjxAkAXUWCzkg4UPp//V0MGcajEkkLeS/Xyzkgd3ouL0w1Xjwd
ZIOhwVkusgAx0PYJaFeY58gn3PXBYigGI862OUEXBDVG4tdgo3RJxL0lfVr62F+M
RLBGok46ZenXxGrwRXq63yN3kYhH4ASL0W7IC5EhH4H/hrDgWnQyv9OkTkHh/wNk
Z2S76TbxlRvYpqCQXoh48fZkaL28CN5k8spU+UqaL0Mg8Yf0p1fUuH73PPnJzIRc
AU3CghnHQBMr++qZVCsGXj+7sjgust2HEe+f5cwnEPPWsjBo8ZzfMeHih5Adcrwa
CLJSFvcFRTGiYPi2LUII/pO5avm6jjIL95idMUjfA1z3Udy4DVPT3LAlHDR/MBIn
XQXAXOQwGrPUC5XTjtqt9T8JWBrgW9pSxZPZjX5VpbBkDN4gFql5Fi+Vv7xu6bmH
3IWMMNCKq0vViJv9SXKYUJJSmzKdZ+TVlGurOPN+a+b+D70N5H89qdGQBN4XzZE4
cYKKRbiHxEhakpvGf4KA0qdBFixaTEM+f00m9sSHNleiFR0OH9thmIysjmPrCdC5
HN4zde3oW+PsLqh6IwNNEDJvAe9xJFYicOeTKfKGzbKzWlRCUT+CzE57R8e78Vj+
kesc4sfg/4MfZ1hjWF1Wtsyrco0+zl1q2sVISuwwnL86laVlfect5GnHYw4Pxixu
sSUS+HQEXRYf4XrnPrQYX/KunxxPD7QjAMDnps6NysU8jFn0NIohfbBzva/cMO9F
DhQCV79ronpOtKmya0hTXxSzCLFBbdZmuVYK8itL9Ay+NPIojlIy5h2Jr2UXEhYz
VRi1ykwwCUU+uDiO1oh9oRcmOHVU/C0j++VHbi8lY2kRgLa20bIFrvMTV+nhqGj3
0r2dqB9mz/kYd/9lPbInhbmueL3Me9fM6njswMrYzUflGgMmi/HkX9+1TAEFyd/n
FBYHA1QA2Xd/7I8ghnVYAxV24rrF03I26V3azDJ25tgmqVFcs0QJ8YNGfo8P+H91
eP2McrAdauZxyP0XrlM/ingXYOYyApUv0Xb+XuWOMBaWGaGXjRqVqsyFzAkbbS+s
E1712w1Mqpo3iNWAVAg6uKPxOU8/4Z2PtPmRGmtAp1FxbKX9Xj0eFVrNKRGCGArD
i5A2KvcW0JL+OdafaJfCmBPs771RIYo8POLlNEK8aM5VAJBHpnTWZnFHsil56DD2
xyBOqAQj/Xz/7j8TpX8AE1CkrwGXVA+MM6FvZsBGuS9ahjKSMx76k6DeUOhvZsu6
tXtxVSPQbf+/oCBDKra2Baew5aprfUsJZibL/cbTcjH0nHb0hAfBBj9TKmU3PEAC
dQeF7c+LPjXs3GUuMvWYQIPR9ODozCRnDpsP8HnUwpO474l8uCW3izRcCsWE2sg4
x78jglQQxWhOnxJwyzZt3Jf7XK3asKhd1ZA+7wIdVZ5Q4feA83r4dTl6xVEIYYRf
zBIBEj/ab4VI0kD7b/e0LlwuuOBDmUw3E7S13au0njiOUBolhDZ9HNd/dGA8yopo
XeWKQvQc/ksczMoV+V6cLbWWfAgKFxlD3x0rcP2FuEegr+kO5P6MtZiAbXK6VrC2
DVgs7zCBtMzCxBr2licdepC8ccFfOMdXUXkS9tagI6dFeZYlzbcvqKAr55ncukkR
RLAPO6i/KsyBzH18LQ8jEpAUGqapFhNbpbhpEFPUInEiK0MWYQM1xjSUBdlRe+s2
5uNqimsLH3B0ddgS7a/6rQOpeEUDlVLFkbLGHdKfRwS6NZh/ld67pvsfcBt48wfz
K83YF0yEsrpN2vaqjJcpelrbnjAI+VUxZ8Svhw/EjL2QGMBff1qINUrGPch7m+iv
vz3jMfsTx+bou03LAPxnvqhJRkCRVdrM1EeC9GI9UPmOanM6/mCo+hBYAwKPtGFf
4hzTBDzoQ0dUgSj53QizzXKVq0kkrH8iZVoU8YJi2ybUmL4NhfizrlEHdV8tO4hU
YiyYWX3wzrhLYvuFhmCoY+gTWzCfw5ftpAuXBxqwOxWAQhMKULl8bUuVghuu9cRx
uSFTqXu9Qfjx3+qGYXLAUXVl25NVPqbog/mx0+oWHeSGy/tKNSDWMXtp/V+PORkV
HYHdli4fpi4deKIDztO1dngWz6vHIvF9iGeJdMRHCWJIIBVmSDAJugKWaKk25NhS
TkprYQoL7blkmCmHrazJ1NdjnbzoeknD3QH0lB+lxFjq+nwMrODE9GCDVK9Tfwnr
hpxNwd04e5dsV5WZ71UTBQTre7EqnHndjXx5gvP1HhWb5KIDtcpxdmvgTZ7H7aIM
/fN44iEO52KRVU5w24/1Kc3uSWRUhH8CsheMWohnyK8Tki3+uAMP6PJ9Ojk6tNmp
gjogx6WN1sJiowWB9fxiHYP/3VTMjnaBp6XJyY8J8tvO2St48HyPPGKHX3r7mta3
sdEEKCi5wK5J2ymEMnYYjOYhbj8Hxkia7ELgcto0M7+gsmI8ANfsLKKExEtuUnhX
dSfse6GNDm94oooZtCw5VkFBtM9YNDNVmZpL0PsjSESOuka8Nu1T7U52q84nmY2N
jBV1Ck1wyT1p1q1btEGTP8PLCaQo/79I0n4j/MC84+fS0acE8EGphNx+C+oFHEcP
QZrRJf0qZx0P0iWFvh3pEdZTBPwW+QbB4S5tSlcetTTh88+EkjQWbD3TxYihD4JI
RVUmdaffJyqw8A0yDnzbp054R7nVsFYGyQJltxKD4K/gq0OXMeqhaObiTWn1qvaE
kOPef/m93icbly7MJsaKxvMLaRmqwZwxrBhpk7XAiSQ3eXtMK+4g7rAkG0knWTxe
e55taSrd5QPcN5LZD0dVam7Y1e5ALWScvDGNZnUiu1DKI1NqKGWi82WjDn/gEiPd
RhvbQNteLqEfxaq7Ty0G9LfLRPfvoMzGbFs6GvYQ96jR/3v8Weuovmyl+B4+j6jS
0FK13FRhmHE/sFWRjluAmhxVBx551LjctC23tBl4dyrqA9Z1RFsSkT8DZugjC/6x
i70ldZa7PmbThPnTjRiZtZoRxwiodMAPh7h9dW5M6ssjr59GI6i8Ae8e0crEAFtF
aYoCCju5x9PX8RlNM36Zqgo9f/jCnWshi4W0RU4CAP5otb4VCSweMvIbzbGWvJau
Ji7IacbUSd+u7szEhpLNeq92WzNYL4Zdv56JkJGn219FPZOZHC65aZB4hKkuvvzP
VW1xv7RGOkJ7EYq7zSLkkrUwJ0b0PMHiqY4aCDLiOgRm2cF33nN0XSQ2HjKs3h/y
p3+4fM3CRbYyXr19CDDwWQZLaaz3s4ScBmk4ldHhv8d+nVJXtGk/6g9S2DMrTjMJ
WZF0PTIW8IB+9GZfZ2TdmWyAwcruBHaxRx01NtODDYWSHN4sMLaly5Pm45Sq8L06
3UAkgM4YcXqZPDDpEhOskMknP0Kl63yQkxSGbbtOR8NO1203r0oMr+9RXl+AYmCi
7uD5T7xwnilwUT3ScP/csvVA7w4tPAj7GPrLA5z7aR0BDPhA+PPZ4S6hBOvdCv9m
Tps4aAbl57whlerFswf1fTxdLfbxrVGL+6yA1YIJ1g52bKF6G0u7AEaWFSzNG94X
rxvE7Sj7yUVtJITea4w3cBEgNARzPzqtVTflCsvsqSn/IZvKQJ06XhWcWwwKGhVh
TsuDJuhoK3W7LY8kI2HiBk0X2OdLKnr2p/p8LaKo+MwA1bFeKoLnzqPSlvfopLhh
mgYnpjzDtSFl612aIzzZ3M8k+VqYutvo/3oCPTYq8qxAXweVoLC6+oG4PVbSYbnu
hlDsMQvFLOIexXx6gDgezSM47hmyzPIQHkESsxyTH2zj9FFj1Hy46r1w1d9xdz/p
zOjhs2bZjjc5yqhQwk4cfFD5R4GMb0wXzv8TaRP7QwPFlBOZbhaTSgjOB2wxlFVL
yKJ+nlMO+wgF5SdHbPlO8TDv5CM7qwdvBJhsSErlj4YNsQkN7lTt2fgxCWnKk1DV
wiLc0dhtcxvVU7Dce4NgJ6bHITq+LxLg5s3dgMcBxgyM/zrkX9tIsRPEDmqiGR40
j0hH5F27vg9mkDG72rDeaZNOEhkPIQ35DZdcntWhL+Hhpcmd4VScReXuvPo6BgJ1
/JY5xJZQ0OT+NLu5ElhZM6+vagtVURp0UucjuEqucPTocbvsS+dZiJpZ7yQ3N/k4
NyomxFYY01BB+BV16XUFA8xvBEumbltzuHh2KYrvIfItaW7zTMsRrBtvq/mdxnDN
EWCnttOGNtLPD+Xh3PaIE/ObRepAh8DFh3uzAb4DXYI60QC/HsYNEU01THUBwVmu
l5Pxglh/kaoc+4DvTs3r7YS1LxSXoJc8YASALg8JgYiAphwcSSN7ezDpeTMrLK23
VkRSw3AnpcUtJXa3l3bdKo+cLYEUVuwE0ZsBczWY9el2C21HazEXlYKCQTL/NZqO
XBIeFRnch8BzX9LM3CCKXi3YXTeJYhuqDnIHwoqImDYNjoTjnr9kzp+w8Is+pVtu
//3UdJlRnNnt+GSoSA09OEp+8R7uqF4ak/YClgoG0MuttgXzW9UoNXMEENseQ2kI
/DlP3U+xZGTHPMfSpf/jhm3MPFk6lx64fhxRrikA6XEhXOdvZZexdWPXvWXHxyvp
9Go74oiGAWsLz/DDD6p3uivsabomOZIygogK1D7+N7uj+6de+0n284W015TzaraZ
eQO/E+5oZDSseZKxEV4F+m/BAT/JkOkwN4ZUL8JZ6saIOFSTpHWUvccBis+kjsG/
LUx1+yNATPTfPyJARghgEOHmzww3+7NFNQG0ksm7ySM10u81bu2/a08L1pQVmiSE
bedfOIXPZc27emqqUH9YQN0v68Y0lCPiZQXZcAnr7n9WYO9NQvckPj8ykvCqDIAr
LXHctOmU31+KjaoD9MF5oOr9MjUdZtvIY9hTTaOZpE6+X+t2ul6G6seVhWoz3Kqg
g9QK6Tw+rdhoX1YTYHEt6luaYBcKpY3P4TWWqUnK5Pir7rNtxeV8vyu0HL4glFrM
DmFxRgltkH2TEj8fc7d5hYb/0H0IsmWYozeTK/F3tVUMM6CPEhWURKWmCYKYNk/1
6SnviJGUNefONJwIXWryhHX0TunO9TAP8FPj5VFwTkjjBe4Dxw0NQ/nhYYL8wDYp
N5LWKbi/OiBAoa26RcKXrJNS132UYQw4UG3uH/6/NkTyTV7UPIkOE6e3ZyfThSHH
2JQTGfhY8cWS4y2aZokuEKD56AkNcw8qZclr4nCDLPt4Q0sSzJMDXXhulDd8QgHA
2Aqm7ueYY/6Cld9k7PIEEcv1cOi+On4rRZ8MhHujy5RHtopBOqs28b+hDfwiqm81
wagFn//5Y+PT+ZjTXo4FzXpEqDC8GogkHLKo3jQkST6apn+kfPG4km4ddnVMu85B
oA5wP8oVqYKI0o0ne5qH5jFtzS42aSjstBn2bPrqPMuPZzgQ5ukgLw4RANhBXcYM
IDWyDncnjTVlVD4yp2Fz58/dKpPG2P4eipRljTgmHjVebomaZbzDt1O9gOhVK0nI
GOoEt3e9y+CDZvnwccCDc5xScv8R0dVl4L3HypOnrcfMvhjrjFVplofGPoTOjIn+
7RvOSSiqSiQ7FUoYCr2bGtRvoZfr1YB6hUNSL4g9pEoKP1qFZuMTND3OClSjXI5d
XUcXMUSy7QqAiM/KQAxofxfE93YJPLHAB0zjmOMruISY/B5lyV4zZ33iOvFe6o5R
HaVR26PB1cQy8EPp6x9YzwCw7CzjVApENTb7vS4tLpRcs+70udiMG8qU45l/tCm+
egSqa8RqRElCTqwiT2hrKHciigztjppvlf6cmufgS4fmQQ3m7K8zwla2Zh8nqKLy
c33GBk9ZaToOTpIRDeOpCCvIADObepUknXOhysD14MO0LwTymkYN1TGM051k3CwN
RkmLy8E3cSjygi8fCRU36Wezmd1Po3O8CG50aBLtGxG9Bk3yIxnD8hH3DAWPCEzy
9xjVJH78UIjgdASFUh3upicPW6S6jCnh+SHIM/3bFqQqo0JLMWlq15RqYEGEzLvV
4QOYOIWE/V0HuQIOR6bvoVPK1/5DDN77+BQwdw+DUeEP7EhuNgYZ45fLUzdrUZG2
vfYOcYe908pnUDW5h0e/rB1hN1LdN0jjG2JhZIvY7bgkfXQY+6K841QRSPwn/E+x
EmUGLLpjQMs2zlg22Jl8ssQ8FlZqRGah/iuwXHjt482kTqWQBKDdbuof0zvzfV/M
tmIa+NMTUot8QMjrTK7GDl+9wCdZw8wOhsigOVZT3fn+KjnK9bS/CZEJycGv5Tkf
L/ynCpI4J3NEyzqcN71ZBNw0evFdI0eaMS3LKq7UVxiDgoPupOiTBIIPo/NcVc73
X32VYSgNW4U3qs7V5vPl/XISdmlJza0Kheom3dz3e8JyCjLwx/W+EuKq+R+ufrTz
kPDNq0GW6A2VtRtraXry8ZMa1t4lO3Nat7uivjfFyRLKZWN25nwIYMBnfvZLEmCO
vObAQpWAmAfU+kwvRhxxEcD57CajfSqTYKp2HSFd2jjtco/7NtgQsyGTH7izkJou
+nBEaUw5lxH07KXttF5eGCNIla4ZK8lIrW7zDOomhp4guBjAZeStvrxg8isUza/3
oSIeiyTUbYz9qaIdPtSWoE8RbhiHBccxn2LzYZxW/EOYPnAYVR5ssZtz4KWDZSkf
m47Rp4DR8A9Tv5Dm3fV9QyILkTU+cmA0hy7LJXnsItoD4E0oiIDHoaSHstYr5/O1
8EEtDNS8JJsiYQatnMD8taHT9HWj5B9zcuU+3/mg0y+BuJ5G0F/wgfsE0HbMcRhw
T42D1KR6CD9SCR/NVoJZHFf3qGxgXt7zP3AldvdW4vxQDNdXQjty3G/UXJTkCvsX
1FRpVNeHW72o5m2cEz4FrSaDoUyMdJBQI0MGAaqdCyjBBF4zmWy2h12DHpYIYntY
uOdvztuGdgS6u7In1lEmp7YSPM/114O7UycXh1kPfifEjoS2/MHvmwXWc5JmCpmy
+P1/SxbVOKp+aaCYuBmW+x9FoDqKgWtg9tuOE+pQQS1+tCrsNd5LLxDxeg9Hbz+J
HVmaknsMjCIr0rbTNK97h96AEu88gEt1zsx4gzx8dtyC5/6ST6xYfpi+6Fh2OWm3
CpcftujObvFDyq0mM+FFZR41LX9sGDnlQcdb5spIUoQVRgnUyiuVHIycDgKlDiOD
8mtmVvarYUmc7F5jqSXMx8T/q2kYvjNUI/SoUTxzFP4J1hD/lwqu/YJ3txjw7wYN
UsdTnzbztRW8Pxu8dOhGLbDAwK0johV6hzlVhvnsWhNL8Qalxi6UbQp3yFLhc5RF
eBN6wJ0wAgvNycmhUsXt60dpPpYo9wmzibyx1VanavNeLfPIlHatnUJ6NhCoXn+Q
dMLBysvcD+bSmG8OKQbDrtDzLTH4zJ7JZOpdPjncZP28t3tXP0rf3KMUR+4TxwU8
3U69goBwudGGyLyyZiv7dLuiaGiWUOdUg3prFsf3vRGrh3WCec81diHp1ee3xRAT
B5sYVEySkPaeOi6IFLVVUAyOy7lpC0z6NsMF7sJ/v7qb8ElGqaQv+y0IILZSThz8
SmXWOQBpqPWp3SgRJJr4B4h2nrNAXzKdaLVjT8qAYG1+P5bqK0qYInNmojs9Xnpw
rg6SqBAnCd6uzNzRcj5vMmthzK4rOS+1ZIyWxO222T0OkyeP/9RcHcBH6nE7nlDv
kqAXnu+U33mhGPiqadjga0rhu1Nmpn0xLd93CAjsUYlFX7TyXrxDFs5jBbgPe+dS
lBUpBmkhAaCdkupzPAwymREnlidYkt3e6DiQTkzHij+IFE2RXkfLP3mykIhj/rlq
IlDTF7KfR8H/gZtE9F6i1QRSy3Z+74YM7mBPTeQ5tszo2Y4uSXYuj/913HOXp2FJ
atp/rlH/QcgfF8FQrEiaToRrUd85aWwQIf9pHyrBT/976pT/BK7BiBV506H7Uohi
LT2zVnwB9kq4kmeeUDiJXbpwoiwd4O+XT5jv0v+s2cIbZJmBUdKoCxqntEcj3xua
NC3Gmy65vYRpyr0YXAFCiGspCbpM4+vFEVL+YmqNrhnsv35yuKHd/ksUQCfaHbN8
OYG7sYhzYBBM7Ro1KptgcLBFq0MkJuxVXiKKpS3QpmQmlSjrgPJDPpMm9hxi6plr
CnAgD4hCS3x2bJh+1f57QQXzjJKkfXtWp5DgPIdpjlX/CyJlLpTaFiuGUqEDV0Yj
EDZFV6w4ANYwT7rErE+cG361JhZ7kt7sSJk2+jjhmu8OHqX30Ag5V51ZQaEsf984
8bW6ZsgwIOAS/s0dfffZGmqXxusfguqFhm3SkftLzsVPvJoKwlphSk+jwJdIzUWo
BNrD1uoFJHMLSd4BVEQKTmoGs7xm1niieWxYhYXjgZ5bbjsv0etZFbFNjM+oBbXV
vTyVeODIUltLUpoQjrw5PUoBwESMrZ6vvANx2jR8oUlxL4a9ritVmajA297ZgPoq
c0Vy8biQtoqnYnwx09uWGT0IRMKdTK8UxxipUo4YQCUACrrkSESkIBj+O3jCDP8Z
1bkLMPyEePYGt1QfJtKdG0+9x2onTLBEJh+6JNCPTfxQJYui0xuMwhCYU2RdaU/h
XjuMRV3wnToyQ3Rm/cpTecdw95l3GlYNIoxVYZttBSBab0auUi6Koll7QHg97CGC
PnAA3UyvVO93UW6hj84G2SAEYvYncSRB19i334LaodBQBbEHGw+GcuSHbbLJctzl
fNsNkAzzAVM6l18hk7ZTn70gW3YB288mKWwvN1qVUIK3xe9gFacANIIEsfUqGfpH
zWayRzXu4pzRrv2pb+bQtxUlotMXwWcpQ/ALdmxmw60iu5tW6RLzb4Io1AWctCgW
TZvf0fnmuCxImU64Kzo11PfhFEDSk1QXAgzqBe+Yqvp02B2CzEes/hpPav34XuRB
3BqyhCZfl7GuTcON9TP9Mff1vjWzGAGNflBGCaupO1mDORP2fojzUNq7sHyYr6Jt
Ga8nv25rSLYI+yetkAQXfmU5Qtv1LQNJyUJCB5t/RqWgxcRJt7cv5w5kxkqZG/4F
DZpSkJB8Mm7/nK4OCcB+ZFGdjYS3okQutj0F2c3n9Vyln8EuVKXshXqMjBLBthq7
MyjKJ1OmpNKOebHeb9y9VRWupPs3oBvYT+wdR6c2bo4F424kkNEDOREZHfs3kfrC
wpzJNf6zBP+C1kFqbGaj1pIIWEU0noxWpX+ylePqQFq9kwUhXHm8cQncE84oxuLx
FGFwn+baZGhSeYlCWkKA08Llt2gR7YBSqbPCJHMsnuwzEGK+GGzBuDyOqyUZoNNb
ahDmJ7g5SC2PzOo40uars3oHqmjUJYW6ZBrRTF0AaPeZBNuDSgEtGch8XAMifq5Q
h3ctwSJutA+MxFQalLLO26DyVTb9Uvcuq52b5pUwhPaxMS6pVjx7yPYHWpdwf8WO
I8wzeacXVt273DfH+ZvEz8TdL3bl3T/yQCjUSDzMq2/3qxPU5zqQI3VeRZOTHgwQ
N/wjRlzOnkqNDdg9/HPvkCXM9YFmFEbXV++GFz4ioAdrjnmwbG3Z7D5ZtZd3P+sf
8mrTorQ1edzxlYugqfaMstn9TcVP62PzI2vt+S1JBEg+7EztSf6zhSDZeEYQ55TU
KCZygM+C4eau3DLss+3lWT7Xj4Hsgn/qWUNE3u6CeFdfCi0uLeMMu9lOsAUfNSu5
UzKEkx8jVoSftExLlTh+NLWvjUzcRt5Gfr31y6vEeM+//FckQ5y0Rn105LkdBrL0
4hty8lOHVD7tx4EpysVqB+1QzbCg/9wyAt5IRsyg4/24Ai0xeW7zR7fgHcMEHYKH
WGS6Ukkg9lIDXDp3JkDERtVb+JyRw0HxmFFA72LD6FTgm/QJmU0XfWWzk8KvysZN
ywey25Hsi4py9zY+Po271oT8huiPE8p/6660RqHDopnGVzZ+tR3cZZoFH1Xdv8el
gp81ABTP6pLIBbtV9pqNBT90gm7akvvB7pONKJc6Y7GqPm5fleKAlRFIxVnD/hh4
3QI4VWp2CTRCU/GQJUcrcpY2ekZItoiCsvStnr8Fltq0zGzDHlZ5xiKCdCtR0Dqa
rmYaZWHrjTmAdOmNa2C1q1YlVMmsTrZf6Jcvi5dt2xC5iPnsGyeVYINZr3GFOZIS
dDumSp+YzJzFussF7nfYM6UuzyfQ2GM5hrudjnRLZqyGt65j4QMrg92ARHuWIv+H
1vx5yV8T8aa7FdfF5iHZXvm9zlfra4zLT4qbgNd3ohlvSjz9cmnk1Ce7b6mKEaPa
JNOMHeexXPw96mvmPMN0tPwKVgksP3KV8M+nbiSVCnJOpOfZ2kZZ3NRISAeAKZR9
Tci+JyDC2UDykjuH4SDS+hRPY+2LRgm1yz1wXZ7ABgPkp3Co7KHITHeNfiy2rE5J
4xE1t2dUtO2mS07vGSSHdf2mDHuwzk0LeP6EesAPuSPNVTro1uR4OQ071Vyl5RVV
3FPk8sat82mNNGfz+K8Qsgbipj2YEtfoAVe9Fbaqgz19ZwwfdyMF4g5gGLVPfSKb
kubaa7HtIBkZuiq6POK+muTgAinrUFsRvE9PcD3ZQoR9qr8SOwuyYFz9G4awWgjC
nrqc+DBXEYpuRxnnSbfP/kyPS6xcj+PlRVO6HMODNqcvnB1M3tBhNs+as80CdGiB
y4vJkeA/NBEpbzSMYNaqX9dpo5lnx+OI+x1Z0OqekMw2RNwlOKMdfp4bLw6zCDcU
Xj8XimHlLGESFI311S3r+5D95f/8pD/YzaeDOkduwDvbJkLCox5cT71xl30uZoW7
c7N9em+hJJReB/pHJSEgRkHgLBaJcQWeGpQxLT7z+eJEt+fMhBI4yHfHiVuk1Ie4
wItlUTJXvJvA63XHL33xnF2CBOLMdJEScbJfJPhTrYBPJglPU4k6UKAclm0+IvAT
2uR6asjGLB0tV9pTj3LC97V4gTpuah0425hDyMP2Gq2KEsOFg84D7SFlMZJCgKMz
nvtP57lALNdREgajjkRBpPm2XgyCXwSKrQ/wlD//JGj6IQbbHAuEDMCI/QP+194S
EB0LeXjPSdaV3GkWJN2rnW81g/7SHOLqvUaFo6FVtIQLDznMcZ4wyFltRblXvvmr
UnYaol/JiC5BxeLA1z/KHMYObcv+jTsC/8ozoz9eL69AtuYf1RaAO8hj8y8MxWVu
/tCTqS9tm0xxBXSwBv4UtlCgZ1JUxrbO+h73tKfwoRpkvTWEyg84a6ejcXPGdcVr
oSspq0zPBHL1zxVcOc4LsJ2RSP0NXt9WfcFm05+8rOU56MpOKFUXt594iAdPrJyz
pqlss2yczlFVqwF6HTCjuSk5Vb9A2oXJU1uUtr3rf6wH7VnwBDafQE77LFQQeNUA
XNXNsRFt6luTEd+fT+6giXzsZUZ/ENXVs5Zcn1/26tHADgiPgbWPuG+YGv25RJEQ
9M6UOvUSj0MAqmDhLtGuRA1H7aG/Jpa5pV55HcIVWsEo107LDrsWSZSemtuzwCvQ
klNs8d9XTC3cPPrIUmjoosx8VVzC5u7frEURpmF5xvQeHLZn5/vpqm4CiChxl7+A
QoTJqDx/w5f8eVV3+4C6am9v9pL6+/mwSLo+xNh6CQCHiOr5ZPdybLe0CW/CHTSa
YrskcKk5t0XT4aQuexStoiidaSaMFXoCRihC3/wwGC16KEWCtizWDEYTnbAHJwV+
tVgqzVBhUmU7pnQfkz6YhjfVusBoordZ2xcmqjWtGbIXCWQz8TZ1ZD2Ap0NWTYuO
9Qq5Tnzd+9+5P1l1nJu5OElkoKz8Xd0ax4kB1UO289ksd8Fwdew9qg3HFEy/Z2TU
5zHy+MjvE2GPKGZi1lilPgwm8rW9ct+nj1SatX2Jy71I6YLhohVfe4fWlt0qewWi
hIWYjIxZqr9ANEw3yIcUDSBdxYgeXP0XjM9GRsLYMrt9HspXa/qUiz9Rl+HUGXu6
eAp8tCyDHrsNkbW05xTwy35NkrlYKbYMw3maF8JbSEsy1IYsm8xIGJB1imGMvaC/
2CiUha9sp4dekYDbalPWH0cT6oU8l4cnCVdZDpP9ZO/K7Gx2Rekm7WDfNzH9hOua
iZxUXkfsIOxqzvrX+KAEAf8FHhnX74ySfi9RD+SyUn4hFg+w8f18QrDFyCDXJdYc
2xnHkvtfS+jK78174uEUJcLoff92w1h8oYEi5Ga9ZkCKQI01OuTrdwy4v/6+7X8e
NinCbND1TIEfSm3KaN6iFx6oxbCo4KBUtETTZ5wfU/3jweCeFzsmm+kQQ4eW04pH
9JOh0FJr+/PIhXcMreprLTzqQl8GbToJzMQFJvt+CqxRL4wt9F8BuW06uVdt32ku
0SxtCPaH78lywSDSaTnE7zbBDM/+RP1xXqJ1ich7lxDRi8GwI9NPydsfb+Y7JeHy
Z7NuLC8I9ho2GekQ4aAY5yGF71csTd5LMofqO0Dac3CNz6/+AdmIJdLNUhMtmTKh
vC5vE5KF/WZYsNWFz6NoC3t3w1ByCEY0tOYkmWAX/1VFazkN8iLryEqv2vFcCaLN
eLpVbJrR+oc8i09e/f9G19HY3s+qv/7ID0mKC3i6foXlNGB5pkOraI3wQTwTzUec
fNQRuV22bdn0e6PoJAaoCjC0WAzQTk/9NAJfFPUSktUstp9W4QwJBOQnxoVHj2O/
DhFgDA6LtlWl/f+lEdYG+Wc/cYwwnpDRR2kWnl4aWbgjYFet5763qDbtP0ElsqS5
HAaWccWu/rkBEFwK8zIDKq5V/YywOE7W4J1ChzfZ+1E0rUrYe/32DdccqRTlW4Ox
OsfUclr8MYSHfNX1EB/4ODDv3YFOj6PE1LoMI4z3H1oODxhFRbhx6dV4f0InT1uY
dT2cpST20HfeT4ByYm3GAJJ3mZFpA3Rp7n2sNWHOoNNatGPnHQb27gJlJ8GDKiu7
hYipznomTPV1tydwJOKbFaPd+zaI8DgkvJTVMLpgztezb20EVYwjrcpahOHhhQN+
QX1Ugjexo2NvGQL4Vpf91S0VkdWE6A4UeM7XtwaogShD1JDsxe1UxXo9M/2DkxsT
TsHCzad7a49nTWgUp9CUunZosMgvKtX+DcbuXYw1LIbTTeDC3+KoG9i+mmIOZ5S8
v+hqOutUP3ZFOzUN+Eg7HxlGqSZu1RfWLmdSCLtyQ4BHkwa5/u0osDzYDE5lRgK5
x3RXbOjUT5xqKsXxxGg4gZIDbvY2cCVe2J8Ct/Oc0f/yLRp/lw4GSiqH0PdF5ov9
rsLy1QD33mkJh3N9UdvaUuUZ4W9aS1bo9pnW6PhSybLxtH9oLGIvhI6ml3EpG/mO
4fPfua8or+8wQEH3qLX+rKLCXpX2CeSJM6iWxF85jkLuOizCklV0HKNlF1YslLnX
mUn/dNRg3MO7f0anrwUmo9oiX5d0Ha9GoyOdXfRZ/Pkb74z/0t/mFz8Jtb1WenD0
wy6IDj159AJKQx1ZwhN1ik8Ti+9nXdNmBOj+XgHB1qAYws2Dg1Gkw4lAOg5vyLNp
IWHtO8zxekF2QRkpp/nw0yBHqm8rZO3SG5PMGMUrsN7MFhnYT5lGhSYyK9fGl3mt
6VocTwtmX5mOkwFUuV3fWGADN5g6zVAdXpsQl1xFxais8VCx+J+1MT1nbKY4foG4
CbgbBdZ+rE8Ra19VlW1rRA6dYCpH9ZqfUeGlSe2z/MMGqFN4H/YBvdS2P+66EFsl
6m7g9zDtLJ5S8XuycnIHVh7202rAJVNllGdSZlsfkintvGK6zbVRq69bWr90FdOe
5s5U7XHb/6hDWM2Al43RfxukYi/pneD4qe4RC0B20P173+sa5xHawlazf/jVffk0
S18Sh/6VZWlIDhhXN8fIrmPssBZtBID3ZYz4Yn58XO0F4kaL8mzAQHDgv0ZCaKGs
jA+WGfE4SrPrKw+AJplIZUAPGq/VOxC8IgG4fZFyG81Xl1+rLdJtucDnQKy2CbCr
SnPpw7nXdstz6hrWXHv7rxlA5/o8/oDCYcSDyYh7IMHOqtjG+cRZ92GqMA8atGW0
L98F4507uwGNI95/opBET9tdEyW2fKN5f1IwArHqe+McLcR9vGLi+H3l6qvmJy67
H/ycYnl8gj3g9Mz7EnKKl+go8xOCQ1zHFifoplLxekoUButgyACOxSriQXmtMLe0
lkYd9ix5qSiXZTUjREN2cwt/EzbtITMt8yVh/UtUpSJ//csmD/1YNB+VS0CiRynh
ncsQvvfOjl+LOlu3PWSQ8/CLQonsRN0Cuc0lrKf4a2rU13Xm5WoYauAsWItLXRNX
o4lqPYRI7mAOdhsFIOJjN5qtFpCMV+xaIPR3LZhvCODLjXydLKzaY9MD5xtSHmAR
FkA3kSeD8AQs6IHJBld+slvhXDqDCCLxTMSFSxzWI2q71BfNhxOPVUV00gNtxE5x
OBjAlvC1w4LsVxbVy7m5sPoYL6wPn6myljI2PO2pxpEwqrQCNUJmDYojqzUXvs5R
x7YIHwR8UZEKuEfS7bVTcefcjbCbv3TSR44vqswpoGfwwVki5/EOSskGlT8xySA2
Ra8aiupPxyfG02MyWfHPj/6EAfw8sm11nx5SBA+kcL664U6q9EmEUTwD1h225g+j
0dIkFTfcSVHJ4sCk5liE7SOxM2WDCDsooifi9HEr7Wt4a7+J3UlBS8U0rmgM4i5J
cgaPOAxPfU/hsQk2dFBKoiXP9S/dHaHBhZlRdppbfBya5picxeUMkptN6g+AdSZr
gDRu/oED/OmDCvzmeIH+Ah/PFTUNB2G+LBAWwAnIR1lewUfXOTom4HFE0LVkVxqk
0wFXjkjIgswtcGykdUdSAfsH/Hx+96NoHZ+qzKdvpS7NmuKGyVmwOS3oeyJNAiI9
QJngl+g2oJASvgjPkNFRp2qwe3N+PyJmbn4cUUttLdd6uOr3AvYWbfwr5MeMr9Zw
qPN9pVcvHzZm3/rlyH4zQ1+Fd5z519hg5ojGee8/NfanMS9+B2N4lPDzwCFtUNOT
nW+TzoAAApIYyWt2sI4vU2zGuJAOgYb7AmszHghL87TsdTlHu/T3zVuzNu4GGpjJ
0V1E2ejWXIQuWa1PEo3HqUjCi9hV7pVawqUgAvwzpg8bw1401wypFL5rH5DCNv6J
TzW0KX8kOlPZiQfI7C8wtozA43TEesJWg8EfEJBqrOIFd6Giro2kwEhsLR7Khl82
DG3zdzIO8XqwKFBVZdy+5Rap2oSUp5yUWoZ0h05mHDsdMtH8O7Zmz+zBmUSB3hj6
+5ifbyTiJJEhfN61EKvHX3wmpHy/3HqYK6ef2V9ielqqgYd02rcXQ10T5RX6E1Rr
BsM000nCkON/KRuIXliPC/yAw6urWJXLUpatUdk+iHuJGpIBTsz2GbbkSmH42Kon
nZe+S8z9RtqIO/W5uemg21oZjVCTmFWlX7c8nFflVBP/gz3OrwUKQWY9aahUouN6
uBJH4R6J0wG9Mm8Zs4fZ5DPspFz6f7n+MKyhiH3x/hD1aGt0S2f0C5RaFYFtal1q
fs4lmFV8W/OTo5kxZeVOwd2hdstHf49XMWyPheU36E26e0lomSzg3DI6Dilvee7r
KLNwajvi+iDYI1FHhZ0MHxCPTR2N+d/5MCBkoxec9HT72ykpz/PrGW0rQF0QkuFq
C3OtyyY9rMuhh212DEJf2VkmQlvv9JbCoMsJylUe/KZ5E8zwxPArp+Pq7cQIaznI
QU3rkOGZkpP6lkKQUipMih3M83bp1XytuCSg7kdUWgO/CSjOuaSnbYtJzcT6q1+b
2KbjcemKb4O1Q03n2tQw47xNrsUCp968TeGSjOemhk9+uYP3aJnVVj9COFIKm28l
I+4g50Q+OpxboIRZN7j3OAr44zXwENl0LfJFDMl7v39ns/02jIeNn1HhKFdkKdB7
hf4yDgc23AVKrVkob6JveVRUrPQe8bp2+LeXuEeDjSBmwUbz2zlR7xrTWXhwELOi
Hy3KOGUnMFB8iqIhtlw0BdqOpcgjRXcy3pH71FyuTHYe3DjIx1mdYIBpMwSI6DOX
hCgxWNFxja0jxbkoaYDALO953pASXNI5MCThpmDiPNfQ2HQDOYGqcHVZ65pHyLcq
0WwukDpet4ewMBpkWtIBxOzY+A/HYGamnbmfOMw0bT/ia0t176xVMSA3Q8tzTzOE
zMcAiW04sFEl+3qOvd4uLKVa8kEyWOaaT8QGI5SQtAF6JBxdf0sytHwtX0WT5qIG
Xs1kWAiyO6BhbPelW943yYe+YlZtMXh8XPzVh1/Kmox2htCZQ3nF1rJ2NqE7bMHO
ywI8YTA2GPCADreB38t/Qr13THZdS26XddwhUwVZUv1R4h2ypwBW8Nwhovmxr0ix
2yVOH7nRurpejxgb13IV1deHTBwsOnilFT9kIcOSsJbMg3AES7GnBvPniOHWmLS+
lo/wMlVdPaLoPAwhiO9oAp4tUzsY3rILHgZPieLYmZ/kqqgVrC43MVnR0Y+DE2wG
ctp3rEup5pEd5XvQ+oQkLPx68kdiko9egcXFD7OOSD0iDWvcfLpUm0BW0d8RZ3ji
+ob+wp8EIATv9JEqvr4l4ncvFPoEk+fTalf7yRG372qXBZ5d0hds5/M5/u1OHVub
psrIvXfwHjNalrrRyOuJTFZVhg+iggrSMK+MbO5UwRIdRIdMzgIe84E/btWDiFoD
PQUmtWHm3oX6+BIdJqXWzek1HTctJi6S4jwbuZb4rxyZQG+TMF5qgDdtQ4lqChE1
gozKWfmq+gI3OESebsOEiPRI1dvOpdFG0KM0VGujh54hHfIfmrIUj3M8kuG5YXVR
JJWDCT9qoDPyDOujKQsme72B+yLGULuZNMIu6sgiUpZHVAGPSM12oODfnfNpjFI3
ra49OZ9HrKoEE/Jk4cwXcQ0ws60VWZJsC3z+YWHvB6d6qGUausP8BM59lT1TkHn1
BJj9uilSmiuILSw7rfsQJYBg+tKzxEzkK4f/RdAOKy07zDd/5JNyjCWpdPsaGd5g
170OpdTS1/ihETyAd1bsrEZheZ8Y9LLHM0aXcXg+O5+urYyENGVC0k8TgNHqNwKg
H8vGDFB2L66IIlociRQ/qQOeFNWScvpcPCFpedrjXAFm+sy33xhm5XCHd9Fh1KsW
vo0nutD+QsuW/YzaAy0VXkz/T3oELxEhPbH4DXDa4n/CR8K4A8wH0CwbWTrhDrOw
27lM+m3o5dNASZK6ZYFiKygisZSgDy2SjqkBwK+S4R9kWuhZfWZ2GyMsXUtwVT4r
4ZtuLnHs77qsK2sF2A/LI7IS/d6qvSncLNzllE0kWFNbWqubBx+2IVOhtjXQ/U7d
QVn6ScSG2bdjd/EKXrNlG4VaU5dwogY4PnlVLlR2R8xHnq1X8ACShrOcoL9TgF50
OY2oamn2KYjzs6E9s1Kqc78enMzofALke3UIl/yC/j+1EH2FSS5HH0dMga+4QKil
A2ycGZEdK/9WEPxciR7UBpUFBrsKnsFnCOo72jfNeFeOKh+PxDWgFtvfpGTEQMHE
pdqLFt8gnbelFtFTrh51iH/eZcaJwqeBUuhbn7jERHxp4EMER1P/c1c5dUBVOdyF
qw1y4pbQi4gQGwxyJSB7/VB/Og81naGu2EP+xAH2thTd+lqEkNuZc4hWWGHuskkR
rQ0VEHfxoIhNQ/URVsgKKqfeTRHrVsSf7yZF0J4RnWRwG5Fk1GBC4OXtJdabX89D
340LFQWiVc++yCh18BeEWa1+ncbqyrK1dCTtlw9FjUx3Sw42DgmMlsq4VuqTfybn
BosBv7tN7xGxMU3HS22RUHFjNDT3NFIsIvnKj0aOYkzZ9FE0P9LrWfF74v+TcM98
z100tJLhPxcAAYeVL4lmtybj2QCHN8uwLYvnHuVQ1QEOJ+lypnOBRk7S1QRxOVb0
4FMx2+YTBLp7DG30lZpzfO39cS8Dsbpa5f33q/ECSl7YDTFaPuWpvNBed+kuWHPp
eZ9OiaWQ+VscMpOrjtlVH3OIPTHtPqiLfSIOD3LfZXybnTDP4HVrY4t3BBe3lWvz
cBQYvS8DF33VJA1F95zEtCheT3PzmSWg3ExUlXq0g3GOvLl/WhctO2qZFDGIZyPE
zwPr58g6GGp7BsXSZkb9G8m4zJsXe/L/UF+OdOONs0S6kkfm6Bqd34A6DmbAd4X/
Tv8TAoYTiOCSf95ARXiLZmvWmwvmOHK9FkmSuIH/EPKfQ8lC+tKLX7PZyJ5FBcGs
khJqvz0fas2g9JqxHoc/OaNG2RMQA+1HM8rEKOgSPbpdytezoZL8rtjvVmBIS4Tf
QUn7gKA703h3w8tQ0XnHDdXt1JtV9W7gfAjyzA5dS85GTRdC2AmzapGcUIwH4WCI
aJtUFUsmLLK9QtEVHOCYq6CV7sbV6Q+cMrPPI2aZW7uPwevrC7QdgdEhG0sGaPd6
dSl+uqgvqRYU6ZeajaOisdEUs8iYOtv1hKhRM305/GxCIxaD8y3DnaSfPea/dzfO
sml7KpEREMLY9bKTNvRpJhmNw8tkTFsSqp+bohXE6XR6ltRsg1gAb+vUr5KWWOxa
4HiaQ08CdbIf+aWyk773pa8Mdk8E2otbtAYn2ZX6549ELreAoOhHAfrnOkxfiOLv
/1MT+LgJZlGMwms2TFxJ4YHeG3HxJk2t9yuSbBlhDrHFIEgXenatEWz0wipVStxQ
25zskBR0Tqtaag6Zn4TFuCnrgI4bPMqCNgW7GTPF3biC5nblKkp1UYuIR+bHwzZc
RL1rGtLduEn2pHp81c+o3o2D96xaGQ2jx1T0Dr4VRWRNHwcc1SforeMUC8aCN1SU
aBNu18QU/M5TUnsKXfK1kctYbwzUd3m3Jpf/1bcFVL6wDO5lW+vnUsCJiXcmT/3E
aEOQnRYYhIhD4v0a/eriVSwGAMbDYV+YBsL2eNhWgNvt6ipGuwzreG+gdZTjVBYn
cmHb8HwblNbGHnDxwrSVfLyHDKqejjvKni9ho5/vyQetg7qUMF37j3lIcNwTCKef
IdrwWSYi4Q17jlR9orYVJy59r8Kc+YAqI66zV5fvP1gt3lcQHDmxB72bC6AJ6Exy
BAJfmO9wd6vsGLzdeVjpJ7Waszn8Xg50qmYRBhXtbc99m1J6vpdMaOvH102hh5dk
B97EcJ+pVfNy5hYdeKA3tm2LtWNi4HFhI83uguDRekOmdoghilFo2ePQFdw9GB+Y
htm3IHeGGbHDRc02iaS4bQZZmWYsZjmxVrCHqN4d55AQM1fJrWes7YNrJDyM0LxL
7/gnVhcmuTO0qOjWQRAZ/antGXVTCzglc3ljWJybDwJTkK5qih4vgGXsgc87ZZs2
kRs5U77FFsQgGIN75HavSloalCkXK81kAwfVXTH+v5vDrsb5DQpzrEbXKmYL3Tm6
UP6sywanV/hIA9e+JWrBsJr2e4jFf8FlTHtnktOzucVhKoKYvuSRvELy/afMZFAe
mmIBZNUWMe8EfAzgQtCHIgfHMYwsLTySjvVN4bx1gL+DuEiuJqypXOefVwXp0BRB
rmHx3150nfDLYJHxSEisC8NfswCA/XEGDHssyH3WqieYcABl6rrtBzUL7tDdcbbR
/T7dKEmGaa1katvXChz8C55guYTz7fSdHNFMnQ9q+MdLn4bkmf6JjM+O3eCDrfQd
GyIxcx/fx00Jdh5JbNMNWcYevAHgWKmoqbzsTVUlKywvTsluqxxcjHfh0hSgRwqA
7ng4xAwAYzWKl290/i1txhZf6LnHjFx6K+x5buBVAflx29LZU0a0Mbxizq7GIsGq
3k4BRtPHXbnwHhIEeFSvhkWJaKjWmF+gbEIJsmV0e9MRdYO4lJ2iVe/raAZ8Gmmi
hVe7nWtEvpUznvMIB0zDulYsPz09BZftIo6vDFLEDlQUpsOtkgD2UkSZb8oxfkHa
j4BO40UH6IhlCBg8fNZ4zm2YpwMqOd/M+ae/VyLoKDNQBGVH1ZZhitgO5kvIk2ZY
ZlVGLj4IgWCO+IOXH30Qf+VoI5IGj8AcdBj61sfCywQ5ZKqzDmWEycu+/yvkee/9
8PWlUPZwBCytqGkeWzGOIiycZC46UM/qMa5QGe46Ffwj9nLaqRNPaR6eB3IMCHwN
9nDzObYHBitlOobwNHb015CRkuhP/SZT+SYDL7ZrMEbCCYoTbaZd17fsMsJF8wXw
dGrK9V8H2YPR078LKOvqrsRHb6vUJvmVcVhh4iR1tKRpU0/ZRbtLsInuz5DVnYn3
l3jH7Tc8Nuf2eSbubBjgYwy9XT8ghUbwqyapo2L7qHhCIQ9fSMxr74NvEszdoTKr
/8NuB2KkXXomtxi1SthfMxfci02ADxSYAOzOQNtBPGYq9SFT6LYu9tGivTk+y57l
jk+lCydkM0rHp9hpfvQj1LWBtNjAGpBe6bojpHgBLmCquZ//Xaxv+WiHkdvBzEb6
gXztcQdoHhiZqEd515gygWHZz2uShmTVkayLmdv/XlEZTK7BKGlp8Xh1V81Z6wL8
uU4OwNdCedNaioQRW5/k+2R2dJ3E+sQYX8J61SH3h1Fdsz+FrsSWC+GsOjgpi/YM
HcTxqxS37eltu7xr6MK1n0nnyHr4cGT9zfaxiD+b9NpJOpwSYTecZOKEvU6LbNv3
5b/p9VkdzPhAlaAKmwXLv7KiIoQURuzcfrE+gg3B6ex7fNl837wsn4JMSJHKSVyY
/+jUY8VUlJAzx1cKlbFB5lXqsgYlLs5xOTToD6UvLh8Y46dEyDviJ0UKM8oaDGzh
dVKffuO5Kny/CcVmAsjSsZTufuDIZCiSA47HrXfyuBQB/2ovJjp+Qr502Nq18BTf
Q1HJH3vvEhHg1ce8ZqNfnkqA1TwXgnOpv37YU9ZjPgthnPxOHUPwAiY/sO9kxThh
ZaDfXQV7nddfg7u+KYG66N//gFaDfS/yK6BFMTCCoRmkYSH+Pv5fYwTKRGu+Ho1+
7FDr6u9SlNTA3jvCh7WEj+Lt7AtuH9YfgXJEZHJwMvq5injQMg0jp3dfUc/WxHBD
sdyA5ruKqmTSyxKaXef1ZhJVtRM9dl5tYu8iHP8rhmUW1NL0+iDCTZs82ajRu6Bv
/0i7Ska6L8B+vsLrEQP6UVvaO9pBNYFoUkZw6iAy/1U5WRXQ94l9i9heUGfZyH0D
pnI2KLopfqnfMCordw8LinecYXzA0idLFLz6MdXCnSJjWnH3pusRNJCTcs3EsLN3
U0d4uWlTt8wY4/bDU4oRJvnHUf2Bx+qJhpDXZZimtfT5CUqbk5P0XS4EWQ0YaNW+
3fWC3Ua58eliVObtFUj5PM9GJXWNsdMRcJN+oznFhMOwFEc9FwqzwylQuNES7ba5
7kebUbpGhTKsQHeAkGidjRHfqDgcEAECD9Vib+5tPRozBdrnlbIzGbZxzL5ffb3g
7V8HoygLj6IxFK/TDCfRdtqt4m4pYjeBnKWgBPzpwiNjsSkzh65xh4EyXgQL40rH
TT0rzGGlvkPTdCFIPJiiZfUlsQl2hRWpOOzN4b+1yO6Gg7NkW9zkrnnW9O0W5fAX
uuJAMyYJO9NJyj16Env/VFpjFDXXeNsMu967zYTgIMwUUCGxalrebZg3LnuRcrJB
2Ke+yMWvjNcqD1EZRvWiCE0lgQEZNNUENH3Sa4uKVJza2Ky4yqAsVQJtQijxWa28
IJLPWFc+oa8Y4m6nH3lSR4Cosy7sn0cmfQJ6fGAkWbImIPE2zBW/FvqK/QIO7+2B
IzTCZbyTRFAYmTs7jX5a9v8VpeyusLS/uKhlby58VHZzRnZe3d0/OTk0++WICHLv
SKNfqbrBwwYR7dM10cs+kU/Zl1R7sYfsGQX5+BMs61VfeY0nbp9GTx5mG8TU1BZy
TrI/rnmeFMYUe/DgIIZpt/BRfPe7pqSt4Gl5qe/ikMRT46gc5ExFe/kQBNoJLmBg
lIZHgckRO+gk6kvMpb5ZMcMEuRZYPX2Xb8jJI/65VLh6UVNxFNgY1pmIv3RNQ1jp
eiXcalRat6ByF8DP/H6St9qO7gZp1PwDVCaFDEktxbdvxC9Y/rr0T21yXtg+Qyjm
z0GSd7zPiCKQ2rv8H2wlIlqHKqI7QRMe/j82MAQ7CmUwTscKPgnZb6XaPziZS+Wb
uTHBmxNQyHA3K+iczXVGOt6GnF4isguPBOR8hqj/9HDf6BCR7lVfqmYguWhk3Eoj
eQQyApjmspi6IuJj3/orpBdF4wN9J/39R/wdgLLaas7Zyll8DRrr6QVqSGkXuZAZ
K4jMNslf8QMH7/jQjXw6fnvUO87D++XlM9ArxyFbDAYJzjXgHDixxm8kixw3cdjO
XhYrn3/zGiv90Gn+kSGBJ4qpTWo/uXUS5iAyj1eiR/78EI2Y7MZoz/Mm9sbwqL6W
/JetrnxhjJLKLuE1Wb6jDZ+Oj2Rx2+2x8m4ymSDNswp04d0BDC7kUe0qdQNRQwtJ
F9dmt+AfxkVXK0kkijIij2DRYW9zFFUp0W612b9A7ddsaYhkNe6+Geee4KzGN9xe
knms1NuapglB04X+e1W5FP2QhQdLGdQG8ZT0SfDlPT1xEr8n6pOxTEQjExl7tscF
KVmPQcLCcy9hEdAktyQsM6uCgPvGQ+qad0xmsLyN4+vf4agA74S/o9e5u9uelkwQ
2a4/nqHMRUo564KbsMcVvkPABSSn4mMc7cpTDjMPovZN/DzQuVnEpdx0hy5Z0w6Y
BZqHJAtTaerJI7IbjAXL17KXXy7nTuBRI3oPh14YyZEVoLFAjOc7oYDxz/3CQaRx
0XUnPckg/LQgxrAs4bNi3Nggcp+X9HNMhTJauWdc/WPwkOgJJ4GaL8D0WkG0kaEB
0XsamD8PHjmzpPso2/2ZYQdTNUaW5MQTqCXq0uvGu0bvtdmJbtODfeBnWph8nV7G
+W/gjrprYIPjDIW/d9mOdnpDa2u5Wb7KlW181JrtCd7i8wW2KKmyiyhX3Zxn9hA/
JeZrWM3LW7je7z7rD8IyJcgimc7ti4mFjHE/l0ZuvwkyatTDrWJ9Pxp2sWdg9gIa
AWcxMg9dbvY4gN7wtk7TCHR9sfx/Zs8XdWmg4idu4GUKP1oTi+Adgs/84cj0v1NY
3JJDPnKbqqvLanHd0DFfCQLQWtQzF2cX4vNXykBvYb3R7GQBc98pSlfPQa+1b2GL
XK7BhsLd0bp/Knnc9B3THQLIKGKhgks/aXD9Xa0VPMA738ZG045pEH0g/jUsN5Fo
ooZMWAYFWGvZ5k507Ik9H0grcMfXNLCf51WBbp+k9J1bDX3g8aqDk1633HznoR6g
4lzomX02aoG4JamwKp0duz+yKaiQHvbMrL2pa1ihIc9YIT8Geso3DvIWs0zS4d2U
Ti1tlGBrwYuRKZVSnKLqmQnB9mMXH9NJ3yBZ34IWhm/gcwWo8wFTqnc9Fk78LkYa
Ym5Yj/VoqEu1tLniHW1SuN3JkDJ/aUbWbNtz81CZ/yIPw0VlEv1qazr3yAcK8n+l
5uTbemj8pn4JM5v2B5+58PDgkK2xSUsp1odq1OSY7zeXXBx3N6KM1KZX/eZsV2dO
jv6omnvkKwi8dQlsCUmcgic8e/QtTlr93TjMxRSssXIjS/GIj1P92e3DYxktI/uv
L090vU8vyq9spguzGb+Ak/r3u45fsFPGi300GITqKeI58RJMD/rfsy2C4W/Gu7er
ZFjUKmtLPOFkYv8KhNOH1GbJ1saosuHjT34mhMVvIVVQsopPzGNzHpFy902EwqU5
3aAi1522JhQex6OiPYYHHPH0e1sDY9oQQmyyajgXj95vXOrPSW8fOkVZWq815BqI
alIo3tuyAe37f2nFDra06CS/hV6sBw/brlFt7sfkj+IKu376c0KvERGP7WGwVvmO
bobERoXMokNAxBiScOyMW/li63Ham6kD5PJm9GpNDDiHwph2SMWBEiR/VUKDLQPA
POakSZpDwXfewFJEEtVa52ZQAwiJxCOy6wKcOMiTZ5ZrOpRY+u2MwFF57cbu4afH
5YKHaffv5Ue8qrugJp1cmLZMwUe32dAE0ZTiyIqme0expNQLfbSUPOJQ6cdFSA+X
FLP0BFwwuymEPFkaTN4ZHJw1XboeogU4cfZHvWqWJNTZcX8NbcMbAfNrvS+L2/ww
17TPQJSMyA0aYykZz16tyZwcmwgNobUwXWQXcrRSKpxyJPbjDEq/l0yS8B7nvN+V
M5bkUgjYfRYgae9SNvT0F5Mvj95Nurjb5aLVmPGExY1+Xiv4tBeaXgrmVlvHKYAg
4geSCuohCuUw750KJR1i3Sy4Cw4lZqUb+5iE+DFD97sqwFAMlxIzz5UwaMqm4nYV
OPkdcCMckiHeJauGDkDOu92BKD2z2L60Kqs9xLvPCsy21nLkidEpPBTU8sgr/ZcU
kNhPPBBhS9k41/6Ekn4Dw0Ofu7HcHCio9EQzB1BCy0J9RXu3qVQ10UDMunHgMK4b
meDBOF/4KVFrSFtFfQIMWvzaOonhGt2SaqLky1UCfsGP3Tj0Um9v1PUud0xmC2y5
JYjsI/BPtgmOteY30KFIjE7IJPeRb0/IhKzkz2owlKIZ1I31NSBGhfFatiseo/mp
AN4p2crqyIzGKoZ8sZhKrWKDWj8UGPHVpRoo4lcuohg7tesLgxKVoeQ2w5G56iYM
nOirhdASAzWRD/7lpZrVTMVbaU9+ozNR8x27l0Ms77MFmOaR2/dCe/XBN2Tun1/g
S70WQ5bsHruNXJ2GNGtqNO8OU2H6IoB/Z81hDu60026QocqjFnG25Xbk580AOw1c
Gr2kQ/soGg5tdrNYYSgmy/m7xp/bBzwWna+JO+RwavCsptVbWPgOXW9uHYiKbUyC
dm2h8OhFRNKIsVhZ/HzJajiZqV/3KsvZmCGVNofifhkikGpqVKYP8Bl3OiLUxTCg
tIU3dTnEYBk6LK2dksA8HOs6mTVoX4KCTJutcsYUh/1+k5MGQY9502dbq3CttWf7
KxncTx9i/y1lhvyafi9xO8k4P0n5PgFyDr+RzjHA5az4UU5sg3Sb6gl5tKe+/H7N
G/T+Mjl/wEZDU7EqfPX3aeKWCD7lRxzW00kcMPSwskNU3owZAoIUMg25j4ROxzzX
GBekPE0F/FJCFcHsXv7J4ZVhCXN8zI9PteWyff2sP7H7/7CL0QlOhdVGhf3Zdpje
lo+s7I4sYxgBKJni2sE57hTb1ngcbVHUpDXd+5y9Ppw32Nka0DmO6rIa3o0qqftG
D/BQv54061JHWaGIBMuLquUea+0OBMMOaNlpHeqE5djZdbDbASVjMeFDhTEWEcV1
Q5VSnSK8/SinCvuVPiWvpmm6TOPhoDZXPjGBxTjdXmD/W+xpYrpl9S7soupBLv34
ZHr/ItuVnRQzRlc/az90dtpIienYeIVgdZkkzAsX3Fz5np2j8r2lHCqA+RMH/BgN
HfoSEQC0QJbyCOceSIfRmacSpiF/iqxL40bHDINwQwFh/S9yzfk/BeNBFStiF7Ln
54qg02LoSrIO/5TYxyYZyNrG6NXI5ru4Qf5RQnnb+O7AZtkvJEALRndsjhRExmka
ufXaalyYrvSMnpLUezhsAJzP0Wvngg0YMD+4m5R69pQtfq3iyqznPxiK48Rellx0
/66jXJb9p/Qxsp5fjce1MKz2342Dj3BZ9aegmEl0o8J++Z3ivOkqiBw6YV4tf1X8
nXfZe10bGOAQm7QWRw57Ym1XoCgdWAsyHCLmkWvSUceaHNKQB7YdcH6vQP8BzYP9
7PeErsmQOTTQZ9zkcUMuVNC+vtSgmtVZjhAq1Jb94EmCRGKSDvOhBKNUKrlnHibM
X40PNHaZLtlmE+CUPJGKQBCEekpYBzcWLYAeOwdrsR7Vcnh+s8q3OmP5Yn8xzwe6
RErH9fKkcekN7eayLrfucgcV96RKn1DovmH46ZNvRxL1xWYFEx7ghon3qsgtlD8k
np85Yms+ap+HL+/4ddRaq0/H4KdkByVWxV0d7KkZGo1u7ggchOf9VwEmpicvKmIU
b3N51nuP1RnedNBvoSUh7X/knkwIHnGxKk9/c836P6NSwcMV8rktshlAVD03M7V8
kMhkeNmLUuRdmV6HVv3VU/vbDnaBA+j5IkTgmKNIvKh5jOxvVtJZ7+xbrr5RRGr2
1m2XuW8J0dZKJt8l5DpaAm07d1a0HnWehQW5UCyAc31CC7oll8U0XACsHMBBhvEt
1WlaoJGug/sogJLxSNm0SlzFIIIWCTjS/38GS9RkiVTBvCSwrUuThSOYsxd4c9BQ
cV2rDlhX79nIk0wzZhSGo5BgwckoMYoZaqisuKKmfiLtayhQGboQRc5kk523JYmm
/eHfB/cNPgE5CZCXmrdnS+fNfChuBD0oWXRFfPzpGLWbZMwsRyb/10rgNOw+SIwH
CPUuBL/f+YGWKX3xEhTxp+Ss2puMhSeHuOFzNABIavANYEKZ3KCXjahwi21q5/yw
2RAKm0FMkIr26soaPaqWqh2xgWJd3VYp0Ej/oeuKwxC3IJ6yYHdOnMbgbYM7impY
K+/fpcMi9f+EEmCb3ODaoARCDOhl8PNsE5NhAsC1mbnjUCBQPbYnZkBB7H+vQGO1
bNzHYYjj6wwv8RV2veUFRgBz4f2pXMy7ykrfTKYtPmhCOGYs4Yc3SsFUS11uIQzT
ZUKeYGmp2iNzMSPP+CaiKMZvTTf6ttHGK7Vk6yTmn826lVA2KINyKllurG+WkSO/
FxTA0ZTU3mJLZOImeqXYkwmo7QOOfOl4aOEv+d8Dh/xGrZ8BtT/9jMC2vPoLAUaI
HOVrwqbGdIohgWPIeGZ9VZvMSjhB0Ugnq14HW/fIr0VysWMKMcuXMT/djU1up5j9
/CMfRllqsgmnFpWXVp8dO/I7lblSxkR2V3TTWVB3FzQAzntAYALUOt1yRjN0p5Bm
49u1IdoN3JGWQ5VSecE4+QGhY8GXUbEdXOGqG5ZfdKQ0ETYrw8vKCo1lgsNvaHiS
yfGqm7jstDnARt3axivvcZoerU3DhsPIhfRKO0aGxtjEZqEn+S6JpRRviGT+DFo4
oPcvSHCf6v6iQWJmPEvSaxVFzkFIduKhHEDBzOeFIdayNvjLPD8+kPAN7PXY8Nab
K8c0M8IX2mSP7f2MWvQYYHU689ab/a9HvWduPOLsXgzQK6v4poXXFSxjQ4RgQevB
RUduIStUpvxz77oQLfQeu7sBvohSQPKUejZ9BSVa/2E2reagHfCTmpqis+P0KuBE
Ppmxpz4DNxo8NCJgI86GLlDYX9mjygzg6nyNFoEzSOMYjzuUO0y8M1bY1rAFVGgw
Xzf1poZ2PJWDjTphBBR7l8+mlhGC6rpMKnR1Oecc5OdGIjX7EC3AKp2RsL+EjMNf
1816A3hy1HCrH8sEX6Flc8b6K1M62rOBTSSFXNyKEUPnh8CjHydTb/oe6a1NkF0N
rDdhy4ikIPhDZsrpDpzoPj0Lp9WL1ovqLYLflk0pLNuEss0HhPZQ0oulwbEEZRO1
rdXL1xklPMhoMYPXQ3xvLIDp0GJzPEuoDvH6saE65vccgmEGxeF2W2dO41zAM2ZZ
M0Z1OW2R6fMoaQ9+DgKD07O1+4rciHkmKPy8tvyt/C5BeBjJ5WjEVcSNGN2Gz+Vw
7nDd23UVz8we/v9B9nB4DPOGpYgFnAAlyFWDl3yUeT2L4kf0A7LByJ10BTSObN2p
8fE+C9SWGu9V8SGf6hY4EZTOEVBtRkuymIMJ4JlQQScDZ9Y/XcMFUjy1r3216Oih
M61ZZiW3Si1Q9y8MoCfRHJHyhqcSvNEbzLvi6b0AMpYMV4uT6VQ7pWniGfTvv8jX
8ClRGjtHlyn6lFGoAw/tc9oGQOBmcc/+YitlssjM6j8IKLda5i8VJnpoy8OM07hd
h+SjgtMn6DS/4xbPyvdtKvFKM99XSowQisMELfWz8MRyEDNFFis3xMx2e4TtcqSK
42m5HwEBqQhJsvqXBy4+8S7Qq8HaiCh8BvGxcLriFELNruQ6AVKBI566Qn0W3E46
109cC3SZ0PSY8hlZeDAQzXRSPyImvcmcobeUWf/f/oxfVXXeigsI8EaymlHpE7a5
b6eNKSO2MKoe6lt4gOYkyMy1uDB4VO1YUslvuik1mNoV2D+aAvVaqMdyx/gpxyhL
GHIk16nXLnw6nuC5J2OppnP6DfjqlWVozCVJhfbCWIec4owpwI/ZT1a6EfQxW/wJ
VMFlEnuWcuYXXoKbveC5W8LegRSX/jZGHvFJWiCgROUT9y3e+4s7rxYmFj49jGFT
C1ZyPytrj/SQquiiJ3YKBT+5ACWtec0yYw5OYk+o4fwi8RboUFq6+GyqYAHsGG7W
MH91qEMMiZo32YMW/hQCM+2LmXBVXSWfEFCfOtgGGduIuwY9Q+rqxmqA6+z6NyMn
EOCBkccHwXUyEGHm3wVEXsMSJuWIQobtDR5jIM8qcA1yMM0THk1l5GrRu6jp9crH
oFNmqxyPctnB5xPoETQaP7qvYikgceGhwCEDXZ+R3sA7+zaBTCKTIG8WHlyhkTSI
o5A5EaeYvWfGM8p8KwVRpU3+0Xp4a23jDZ2SkPsQhfIhHlUT8kayLkDSnd3C3pLJ
cUCwepl1FObLeWDXH4A3Ko8mmrmz2nCjsArSl3L6U1mZrPSOXUj/Lh1rAXPPa5fI
pPO24d4z7dAmeKicJWpJA58cLXcS21DWUMVroCF12aPGjgINYucUK6Uf5mD4gUHX
WqKBQPj1h7r1W17uCiVNTBgM0dJnexm63KDDwab4lR01QtPMQ4R9WMaInmWD7GJ9
Vs9HjxaFd4m9LXwLjoOGEd/jGU8WndZgkMo+rBC3l6cvcfoawa4m0TF7tTpJQejf
yrwaCZt8VGM51KSEm6bA/4WzJdMiWezG4Emhufwi1usxkTF+jwGTm79eJmvbC2d6
ugtqSYwiDjHyGM6r1sCUO8sZoO3fMM66f8d/YLh4EGujyFHoQeilxBq0j/84wO3H
GCmdenQtABZxHtMnayIK+2ds7MzhlHfdd36u7x78fTsRjNCFkT99H4BFdnVwBK5A
uOrp4tQOtKwfOMiXyUhyCp2CkLHNfArUBASDxxLRf+7187BKtGuiS4zX8ihE40Sg
b0aMtlBH26tkTSFQoKnR/ow44MGRLKiEq50pxrcDDE+C9JvARBEriSnvLcG5Y/96
gGAIh1avgM4J0z9fWUv1rsywfxQge6qWr3upSn9Bv2yPPgs8S1yM/FJdYMnafVFS
O64qb4NRmrWtNV3cLohTmPhsrQ/HutcG1tyjeWkD+XMxzOOxJW2NEUWtkd8NNPAJ
php9ztPw71SB6DkjJ61hoGBD36nY393wZxnksSo53csPrUeyJrFvm1+aPTRF8XEk
VHDhhI3kSfQgvbiJdpQoQAq8FoP3pU7XmT3z+O/IWyieQ6C635rZJ4Ey56ISzh85
b8ne4NfSW7UGKKolcHYYosOt4unDbDwv5dxCOE0b7GxbIqIbAHjRiXlNckpMNFBe
kpIQUdnhfMdTF5D+X8mO6mYQtzC3RHuLbE/Hoike1QbUBA5zfDp9mP8HMScskvq8
S0J2G/vea1bncnZM1cySCeFV8LoeFvA5VxJXLS+eW7HC+cLxmLs2RJMjxsgNvETa
sdwK1yKMkuDNLEBbS5lLOFG1zADArv3x3sdxZkCxcFMGcMmM7LOCNRN9jAWiQdmO
rqdQQBwN5G7ToHdA+3YowzYbzenfdZEHBSpW1H4SZvrlIAaMGkmvItrEhRxCYO3m
S+kM0tbA0/gobGvdonwg3KXZIyVrNjvUQdPsjXWwPfiblrBvFcIZXp04D0pvn++/
z5ddn6oVAV3XY4mnNBk0BiN3OeEXz7rKROZWrAl8QCFxZ/susyAhvdHiV7MzXk9u
H5sRzosOnfeg0nKhmDK5WyQ05/l5LA7vdjTn5nr5TofgISQIy+I+OWtc+X2alQCK
cHtoW17bg8o8TMvN2ptDues9Xyt/xhLRWaNhqiAYNJvXl0LVF+2Hy4dnWe/T4/wT
+AyI/E0C761XOkRqqkWlR/hckc4aehHVhD6DD04TXay+owcAkmW1AnVMCRhEf7eL
Lu0uUNPwHnV6SwQ8PypPTHE+o8+I+wByymsQMPlT65SIjROEsmd6q7IZag4LWy/u
l3RPbs4pwSCQgpCN+M8DzFRzS3/20LQUFPCGY3h/WaIhRww+X5somY9ozSBU5MmR
jSZYZVqH0w0EDNuZ/Mz3cLIZzWw1ejMFmSoTlizgX3GuQ0KOeg0WwQfckPG5Rx/V
r0n3jn7Z1T0BV1DAfvEQlwFzbkSxFazexnAUiMcoASCZBbTwD6xJkE/EcuYapkQS
FExoTTESNFSPHqhBC7NPXJ6bmtlXhU7LSQltIXVPRRCNyRlxUXDGYVUgZwFxto1Q
9Ls7UKeIFqrF/SXL1EfdAXFY1xuzvdvdHNvTQh3wRsXZygg83xD0iw5L/LJXIjJ7
KXsQsKao2F2F6K2EVGsj8K8ncw7KUp2M1Dn1OBbQxd2+zH6JRIDjBw01Usi9o+N/
8KE/AF4kc477Agvxq6FV1T9kQiWwF1Qrru+3uhu56DIId0nrx1aQYRizRGTdtlgC
KIy5rl6UW7Ad9opwPIY7Gs/KReydQ8nhHP55PVnhDTeIIhtFEEHvUVToihPwOXW/
NkyeOOLgQdE9ZV9rc5EoZYeCIddoueOw3Z9OU2VYEJXiVeXZ7hBKww8ymouAtXul
+mfXLB2nGX3sELSqDzvIXDhUxXeeA87LCN6eziO986bhNXQkZuMUwPlNSIra5Sse
Vee4XrBfgpl3pG38L0q+pITXqM3oqHtHhhQMyMnJ3JBqfWQrS+q4Rnacxsd1wQQD
iRWfC8BfO9d278guK4rOvMDeEl5O6H8D8naVdXqwNxWwR6QwLpBK086KLPgtLErs
fUmB5cZfU/d4cf0fM9ffI6A7GlHdDC7+NWsxE4ujnjdi1K2TbyzTbGushGAiMGGb
Ep979EprezX7Ajb14XvFTWKfpi89+0G/JvgHJ0YLMNc3WkJ8yQHERVNQy82lRth+
4sTRPWMRXpTrdtFSiyVehO73kxax1nekNNwPJF3L9d3OvF4tqD5h5GLIKh8afhs7
7aUGrvBV05tFG0dpVeUZaUafE1rCyEEvqlTJLhYlO0+0NXM2uiw66g7pZaUyHx+0
kOT9EcM6qvDq0pPgwgGd7a2Kqew8OVUdCqpxgn+bWuNc4IFqEz3hPt9DCUKAPjis
5WhooyEkwzmy1IJOKlv26rp+Dp1ZPDi9RuTD4OjnvKpq4xGSwEeAfc/cpd8jfnJX
iAnTuNJneRUhroGR54LnlL2tgAI/sFgPAfil5KB+BXtylo8PV3+9FfNU/3Qj+9Do
33TJj+LbjPBOgxrpDrdTp54Stu9jxXDWfYL9BsWuSu+Y0leiDOyvDc2ifnEOG0px
8AT6XJs3XuYfddf1V1EstO24VwA/tKhp3WX/zVYOA7k1D+J5dclNbY2Ou4dwrOTr
KjFtr660BMBSZGt7+9sB6SnyZIpjFvKARWUJ2f/1573Do+RUXFWPaTjoVLWG8cBC
8bBXeiSdGHF2FgAY+dVOPBEftTOSnXGgDgZY4BT2fliSpMt0MugOjyKMxJ79k8lE
lxyutrNojcImiZDDkxo10F74Ky3GpcBYXqPywE9/54/+cqSw1Iu0iAUy3XMxWOio
Ez5ua61PutYpDRquxlc+FYPId26l8NbdwUc95Nejpyg6wm40acWLNjXfWmpvy8zE
uZmiCloyqJ9fNuQxnsYfhzdzJAcd+vXRRm51xvNKITXR0LpEXdkVRrHbSSSWdHxm
SsUeYUQVY6U+2kmMa/yEw8IXKeQM7TWRjB8fdjq4H5lzfZIJTvhU6qwpHdPM9ZiJ
uyISls/XPvMPjMldlAWQtObDB8EQ1piJhBX+WXmQinuQXaOoi7WpSjzT6T9q9yM/
bfedWcPgzyZ2PaSwEx8L3yk2s33x8hDTVDQ7zWnicOzn/vNiaf3Sq66PD99lXIaW
y3RHLjw5ULBlWrGleB7rTTpTcjfXO2+cY0OU0KPRV1UHSk/MT6A/F79nmNMOJzM3
MyAof9+p0kFEIiZvb0nqXme3YxgsiqTVK86lWCWFs31rcmpCjx3E1ojYkcNBS39c
523771NIoqW+JcrfhNA35O1d02gyEbMLK+5M9gHWz8SEG0rZg50qUFMYqwsp7cOz
UTggdNgD7acLHwq34mtcCIiQ9VqYkegzuhMBAuPHzYxJuPdkSL6YOv28Eam+6mt0
tJk1Sl7Wdk1NXgBayHA/p6qTsqeadG0Zmt22ULr0ChWtEY17zmE3+gZTLEaDl6hH
a0qQq+LJlRjLr39JUopfPRoe+bKhFswv7V6w/L3Rf0nymqGkzTWVoLz5CuMyb/+p
4aA6PjRFxq+4vnZhumUN3SC0x5Ea5UPjLqQY/lWayDoCRmTrxW4UVoBfeU2f8pLt
76kMuh7J7qgZqIanmEGXvIKRWyfPPDVbjbs8Q0KJQrmbZ2xLO7s40YDkWlTXOtdr
YP2Sqb0F77X0NsKTrr79gfQ4cD04CgvuA8w3B2OWMLA9itZihf4gXNN7+PXBrqaM
fXlVFV7jLxjg/vMLa8q9lZUuMrNhblSjrg/REdw7+X7ry5ySRkdEhaPImzuUAeyA
p6IY1JZGkRXWS6IyQEe++ebw6MKb0Wk3906uNRO6p1IhF73JCbo071mOeevKOMTl
6BSp4ajNc0baFOEgHh2G8isw65DnFg/K7m/74JaKdvhoWRFwknzOQw2G36SHT862
pbE3dkHVb1Ah8itvtWqPZWV/ZLPVTiULN8Z+HtugODFuJsUAqJjlgxpcfG2zkI77
TwradYZ/zn3rQhlNYgOgfAukMOI3dceakoBNaPhEFc5BioaNA9kDgOl7/EQG6vGo
Kl0ToStFMRULVpMVYlIz1qminyd4uGLKMLMDp42LdZemHapE29ML6qqd0uPOBTH2
3f+rB6fw/sdweq7bKaLqfiGMt0Qaj/QNRlOqB9Hm2y7f8teCH8AyzsOJP95/tlSK
WNsdjct82QdgBrdUmg7WHnzaTGWt1OXkux+UB3YfzU+EKppsqVUcoANLnuyDQD10
wkBlpSvMno0EY6C6w1NapuBSWThWJleCfoabT3b5rWPQSZPpq8+A/RACs4v5Yi3s
dTdeeL6no9yig+HCHs+tz9QDkcsW5he32vPo0hUKgbY1Xlc3kM/PBZ+qgHoh13Q2
fMIOura6rZOoO8oG98vFdyKdPM4kIHZFMIjonCt0xRcDr5gC2beS3mVUO+WmvXp6
jXvVDoDiaIzwBK9aXuWAFswsxmtctM03lbg0CdbUdMSdfU+iB3ZQ7m2CmPnqRN22
Yl6G3/AZC4OiTkt8Wi4sCfYpAKIarqSGOD8EHFXu2BLE56RE/fYIlnmS6AjvNvI7
zoCnHa74jhWPK0oHwtb5GsD3djGxWra9niPbYJXSbsTHhJLgV111iJhxkoiTpmLG
cRn4vvEe7b/+zmGHoogdzf3RF+yurwX4aHelnS3CMZ9MU+cJmQw3c3AMsfg65pvG
NF0MFnV623EkdOpZsO7IDUE6U/xFB3RWGDmCuXG7l/CRQQYFIFEvaSt6K/0ijeai
moBnQ8or0rmMyquBWEM96tGGkMP8U8mCMQI18mgiq4l/wObAMQuxLq7Bue4CVz5Q
E7EM0sCvxVXZD3aoNPEydM7S++uvxePtHCvJRTyp6ET+vEmye5AB12LEXmLATIjr
fzv/mROFACqQj3qqJGyw8ZtlDbDNItkQErcTTmMuL541RmT4PUfy8wX8HnxfYwA/
Xg5ECHxJUtFrLTYiWx16PxbGjTl910Fk0nJkbBzWeP5HO6UAz/cXuaSDSLFOpCcz
iStEv89WzDJiAq1uRAdDiVoRjI5N1K5F9x9dWEfFXzxiV3/x88pxZ6uLv4qlnOra
n8WKurq9ZarGIQROp6tjVsBAyPItj7ZEhdVkXvnXKTSakPbx2QrYM60mNgjo6WOB
RcENC5NJSm6yx/NWrc37tvtqErn+XrfMD745ci97o2CN/6NBEZifR9v5rQA0Mt3h
Szn6ALR9Z3u+5ZetotpZc8J/hMVNPn+I9wzwVR4A2oSPYgyXeA0Xeg7zno4j6IBz
vNTcNoK1HgKObVuOsrCB9YBjKBbk5dGoJDaSG9SLjZt3JTdV5Rwq1Y1KOCnzlmyY
wZh5WrISv8HB0CyeOuzo+f48+ZJ0Wo/wTr0Ab7PXQBtDgMfTqPaC0ez7x3U0IKDs
GGCCP1EEsLe4b0zMncd2FRagTgSpm6u7AXpxzEiGm6kZ42mRadohWgAnIHhumGp3
U66LXtvUDq2GVWriuQ6nZx7aiaHJSMnuvT66IMjnFu/8+l+IPL5EjLrEghW+VgBK
psPHMbvFq5Wj7Fr4L+M65u54xlXoXOmKVcAYKxlpw/wHYReZf0tn4LGS96RsisrQ
SQ1uaKiMFknQnLrJ8Te4DYNRUNWJqnsKJjJ42n/jYIgfqXr+6K1O946Fo+iUBcXR
nCY0MIDkNB43gzN83fHBAijGrg+NjWSry5p+9N282+uUema3acKIaczyp0MyaNQx
/UV6AkvBi+EZs1vYpo7Cj9r8MeuEOlH2CrryQTqZWFlk7haOSmqlOebg20WZjyj/
RmtFL4+d5Wt2468fM974OUEmus96zhMCpsXqm1WBJxUJOqjcx+5zthML6qCZ0k6z
4InvilItly6/YIiwieGlLkOTcQI6rz4bSHNUQ+xYHfmLA+6gTSPePhSWXzkZI4xD
XaYRDIJXvFLXzTo1rceAVGX4DMZuq05deYscSmwDeUBlES84ythdZ2rE4oiAPdt7
YoOdagscuX87I43Lq+ITpmQIaj/MSECpmrkwA2iQAdMxBiiCX9rxbeyAB5al4pNa
5tF69opP/YzYH6ObS4FeFRtNLhXcOrGRX4TMT18bR72OTNT9qkO8cTGfwk/ubW8d
2kgQJM03+Q+HtdIgOSIXNNrMpYObZP1v/duLpygie+vQW6kQXR3rcNzkf77Ojk0B
pbker2DElvotYiNIvwFxTaJnLFbR6GI4p9GihpsEYkM1P2hF/mqfGwBbUkI9CLKt
EtVHjnWYp1uPT48O6p99y4QEbnJn7fauVNN7UUogI5JFUU5diYVTWE0kf98MwQwC
MRtZdNi5OdLjiNRGoi2ct03xs2fApnbuyzy+mVzYik5sPGwQSBFdYwdrCxY0flFE
/G5BceUTs6V1XFGGdqJu1fVW/IfuuiGQXtogWOAdizTweMvTbE8NrThSfXqZ0nyi
Do7Ly7B4lBRm6tN8Biuy80QTfvyfig2Brrcb5fzLosYYtKOJuqTIlrBmqNypOBdR
O12oWg0NbI0GGgWqmDtc2uTGNhOiCyl45aFkV1Je5hc5q10LpYANsU2ETsVtFy/3
N9xe9w6Gj9mqm5LZaTDjbO93D269+n5MyTng+sI2m3ln/Zd59bpl447a2jBID9nF
CMN1nDOlKa0ablDJCA1xJEdwzxL9b83pqN6ow3xa70WFvMY/8oMkrQEuPhLqLc5r
WpkJhACQsUGQrM1l6F2Wxb3eLSMg+zGtS2JgQZfgABaNSzi/1VgxHX8TWN9+BPa1
xf9Apz/Yb8FtOdwDVrw6D2qu2Mkgf8mKdSKh3BmrVJv2VL09XhrL2txVg+wq3Pcv
yWtd55O0tdIVrSUxj0dxNMW+M06tJGaaO/OJCJyApRgy2RBOiVDKmLvzXbH0iGPJ
1SNXQAafRSjkW1bBISYdmBBcZeBITDz+kPP4wadZymFX08RLAbOuSfhUMUkWX1ni
+uXC4rMHuw7M3IBFF6NCJlIpIiHtFry3pusc507QayiGMa+HeWsjLxutHV4Fkhuo
84XMjbTqVJuwmZnv39TEdb4p3Vv7I1iEfPXDbEBLyI/sQhvjvLj907OFximJZUx/
7eKnycPeh6SX/o9TNB5ZBsy61mWSrK5V7m3jS8BUeUNTBKavepTZuwCkR9d5/s3e
891nq8Vk4Jd+OulhtQN7mMuVA8vMyDISaX5sxXhWutD2Mdlu2ErZ03SOEQKwzQNF
Wh/pU9KHkGadBWPfcVsYpIoS78LciFzJgTlVT42ydfiYpVUZ9vzOjYhE8QTaqILr
thqmjNfBSEHnW7SqMvgLG0GQNrp+TJXDqaaXR3NrrqylMYAOXDkpzjnL5UiZE2AA
J9tXHZEjUWwN0viaz1gmyxS7ol4cTW7XFccY2DkR25LdRlzEHvJa5V/SKHXL/a+/
wXEe3cWLe2Tg7GntCLgRmw4Dmf06jnevJ6+TRWPJnZmotWTzkkxPjLkjYGXGYew8
uhEnE/v46t8SJ/qbdCm6lfPVPGUEocE0W3SMTmIvPqB25+WKnpeMQ6vPRoLZ8bst
7bpHyCo2Qx5wNWLuZG8E3ft1DkQykM/nf2TccvkOFr0+C8QBb0hV6tY9bGlqAiUv
JNfmdDT64clp0Zoh5sTfG2aMjmcrlf8WUo/HlC5OJKZ4eGbKMFct9DZH/xJgPJ1I
+Ii3Q70yA0gWShEvrnHLaPTdj2WhEAhTcNfr3cVfzlfXOquuSAHHZW/ekZ4dSfWS
Ls9bLi7SUPi/r02RV+v2Ud4GJMOJJv7KNIep98YMid0kvYJw9AgB+CYZgeo4VCo8
ZGK4uHN0ymHQXotc6xLMVggZGa/1zE1WQDDdo9bhG1CrrOhvMPsao5U7UqTsqzBE
XMcufM48sVy5DF4ZdA2Fu7BrV4xxP5P43egSPye7ErOxEViZVXluFq7q/2HYhXng
2Y8/DVQNamDBA2b+kLvg3UpcO4iHGBCi+hp/FBJ7QcJUGOTlSzbXGcA/vEf5WYb/
0Tchix996s/BMNw+GJFVfDdM6BF60NBIhyTIrsVeiTH6V/5GrtzK0gMq5VTAkuaE
8bC/caBaOVUtT0kWus9zx6av7O5utJd2yyk3X3lfjAmAzKSq3E58ZyaF3PifDdEv
dXiroc2VDwpYdSGnNgWGdZ8tls8TZWiuw9sMkk3ze0Hscn/8hNvrvGT8/SjljHSY
K0CQFfPcwUE9V1hks7w5ivRi7dhsuNV8wpcpoIb6TfSMNTslwog8OhYOm8pKkOkY
zq70H5jZ6jIlmHhIU1fkXN6sLAL1MjNPCzwiCRmujk12h+beYpXbfLN0VPaPUSyf
y4epCpJfpvB/3BUsbPWVG+8DtHpN+pPJnyb1MYpe6ij7qf2ZxXE/ZFCEEpzhZnfS
9DqdXcRPqSnNwldeaWub6/myJRU+6IUHaLXRLu9HN6hsMSxk6maiNxlQgMSeAW/L
OVBFNW9I8YDGgSGSvljA3o3S47ZaTycvDAQisXoZCEzzI9Af03dISEyYEvAf/mX0
eqtIrAzkxuDZOyFK0E9r1r7b9nnUrfVWloxOmZqMQqvEYLz6N10SRNjWwThpmMwv
ntRwZ0bBAcCpQTq471/qANUizU1jCfUHTwvQTnq0k1CY5AW++O65QiGJ1oOQl6FM
F0weAcWfuD9wiwYY6f4qz9+jxIJ/7rYmKF+eY0LOsps9pTGEQT1wEnX9RiryHbDH
4WCHL5Hhpbjgd6wcjMqRtOuuj4OCBIzoPsBRuT1PKRCoBnJyS+vioRy5h8OZ2R8i
6y+cWX8EW+ZOnu5ajJ8o7VocEsSfW2zneH2GSnWITZKpog2XRE+nksl8a8PBKbN7
psXbpj5VhQ1KDlPIGMnzaWIubxbjKFx9RiwsPHrbKyM586YSg09LAe9+wRrVqHan
NI9R5pPG3OGy/bBsWbo+a07O1xzG8rECJLASRS2y6Vb0Qzq1Gx5brrcSn2kyTt7L
8MmLqOb8uWtMVceXhsO2dH5SqF/gSxiWCpGV7Bgw6xyfAGS2MdEGuZd8uR4nAPib
17ER7RRXSP0P4F1nfsXiwjgIxTMlzukM/1/wmrUtY0FMyawvfxTw9lRIp0o1fqEd
+foameZ510S+7UK75BaUxzNo0iug9NZt7S1kMEUK+UeJOQUSHYCGF/1BrsNR1sOK
D06JUlkpnFATlnA9IgEbRT835bQw2Kr8Epg0yZSZG6MN84lFINEZeYd2LROOW5Uk
ZQ6VM5XzlxxXh3goLk3pSyU/OD7wBTde7mNXDM2STYvmqh4gOaYb42lLrb5cOB4Y
MiPadmwVmYIhxJjHRNw5V9UyR8uR3FMknTkQegTNzL4i9f0AeYmysWG8NVPli8Fy
Lbu5xas44NWH6+PsG9/XeGAVgb/RI4bYPwDilBGoaZRI4TC1IZklu+AFh57Mqmj+
nnKDSd72o9CcQD9bFe41GvFb+maG4xxduOJxp2iWmLi7N5z7Ffli5D9ctyANFKzz
qKrd924UoTwaYv3kagGeij+jo8ATMHej0YthMmvfZ2vnSoqjrU0Uy953cddkvz+o
vUtZSZXdzICnuouKzIc5Rr/MHc4+VoUOuHGUZ32ZMIPx8HCurOyOrIrqxs5xGsC4
UxJetoAQiqwy4VZeVenMqmwVSOtRw2NDpk/LxUwyjBUp5mhZ3lXrcNFOgkPlT3RM
rdoI+1o7yZNip6QJvJca10pqzP+C7yfdr8BWGgwR1azdhuX6mFBwCkAp6Cc2rIL4
ZAT82dCNeIt8vkmxPLQ5CLtc+A8mlwgEWaYPHMeLv3fStY28DR1Fj0T6KkL1t2mE
a7PEq5hQj/z5Z5J7MhLKEChbU9Aax3fleIDyoBmzB1gitVPzDxypFSGkQrmnnTN1
GB++d58yL02BvmeURkYa9vzE0AFpfNbqDf+8O7JinhXHexsFGOugB0TodA4QzGp8
2U5J6nWqECQbhag3Rag1HuNNRM5f+4qOuzVHoey1rKe4BqKwVRH4D9mScIYQ5+wY
GA1iZ/RCFmGVkrP6Bv2EnvK3SWchBBsTelcEmgPY5V6Sn/U0nVR+BOyKz+E4SE0S
K4Ve/D1glOkHTRnf2TQas73lbksT0k4jh3yENytCiDAoEOOkta+k/lpV8wZ2Py5l
8PVMd7q6daSG4VUHuWf0345Xi6zw6dxFtCMczmsrYvYTZhoTqNLioBj9iqfjEqLu
8VbaJQu5Xui53XmHMnrOumf++f+QcL0dEJjXpO5EPQZoN/tYdG52BmrqXzWOZozl
RFFFxEflvdfJFxTWWMYWMo5Ecdos2FGoy/TehtoUY5+RQ0VcNCJ3IBUPfB1sgp7B
kaEEqva5xX0E1Bqfzy2kcF0kfSQz6twjP+h+scqpmnZuY+ZgHGAfkGOrHBy6r32L
PA6cUm9Zh+r30EdXmBKsC7JEfbfOAHE/GesCu9/djLF7AUBR5Hss4IGyrrbn368L
fgva/w0ynTjZGKJf1xWFbljd6AT5r8rFm4E0kYHvdAlBAIpwAeg8v7mdbjp4RRuf
0l7NqnsiJhY6tD1/yiNDEc3Fi/m4LDVUDYgps5A3agKSFhxqrCpmnYGRGXCN/Q3O
/45UUU1dsDDSUR6WuDxP5v58sUZnDCKgCkQhmZLZ2p7NLkDELyPWLEsLB49Q4xgv
fUdzOVBJRSHsgtKtbGZCcQU7alnZf1lDefBTSPp5DCgZK6CZCvsuVgkRo4+kohab
wVHGRJiJl1JPz90viHAl64TSuSxcdy8rgclebsqD2t4JMWJvSb4ewQlc/I91l0Nh
l0HjeCfpkKHnA0ROmkJJZH1P2QvFOLSBeUYotQrxeFWuJjfg1lIEPPzSTx5yoj2g
cmv2TVt3bobKAqKADicdeIZkTnDtVM1LJpCGme5EVcx0ZaDFiIgdBaJRjyXqF9zf
YpLz4nYrFZDVkNh6fneOD/5iEbL9VskJ1txsNc4TZZFubQl2+MJim8p1WeoqQOlL
lEThOiugCo45HPx0b5YnwjzOFEyrU95hr2UHiD1UvmfPEOHszoglMP76NySdsGy5
ubpMJjQuiMcnbBW4Po2Mlsz2cK/apbFx7/xoaOarrkJvjhN4GJj6SugMR8f7O1+a
SozANShIF4ahy2cZxF0P/xYa+6wzjNJJNu/YGe7C9nXyuOUjuTlL3fX/aHBfaFtv
fSdOeiOpToynJKMI5rASFXE4rMdMuFwGtef9eOtnO1H/qRToiFIX6I4jHpjdgYit
3ojuJ2oScePiZWlSqyDyu0yQplXS02N5vlgORpaLXPsh5Pq+C0zqfvj5ne/9dOSU
6tTV8uaDZ5k9xzbJPj7oY7fSEMEwszUpYhHgwUNGE0DpjYRYvNNCX898SyD2wgoz
RueUxhCagX2T+XkVlNTYNvr95oIWyxaKO4sEsvNg9AZ2VlEaPaUrCREZaZsxAEZc
wxlbFSUnM2hsgV9NpT0dhIXJrivT+S7/u4kYgJTvwwU1JTlEk/E1bqY5LVPBCojK
kX/Y/N+0fAeNNmgjN8w2kuTb1QbyAIPTXWkdBcSWWUZWBvSzFUOv7SNlY81PDRB6
6D4W25G356DECYFjjNX+Wai4tDbNzk1Z5xXLhVF9kKkzTdnrXnaYZw9ALkuL3xUO
NYYSgQrJ238QPVBjDWPADVlF9DUTabsZppzt6lPPz9mEzvghep0RhIFA/mRFbN0F
GQDcRzQf6SFzgCQAlNt0XQIDRTYh3AOijpVrfDQfTk3XOk1pxL5sgfsCGNNCiFa/
Wm1N9J6kBZhxlDviEgNYKsw59jIesB0dTLUwUMcc2DAKR8AAXx2UoKaoN3llRkjo
9r/MDy1oLtGDW+/QjEGqOerx/4RhVIogB6CPyehHuJ1aekr0fA2bUjLCZMSdiF7S
1RxnXj3R7dddLWxQV5NfXC9jX4Pd5iibpo2S/ruEXLA/rP1IAR54Sujyl1uZBRTm
PY18Tvq9UmXrDxxxMVoyScBJayEzHrBgrG46BNWCPXAV2jncnZ81JsJh7mJ1Z+kR
qgaQgszFCsUBX1+/kKOR161sEphFtZlHY1wsTxit5csnfZCiegMOAcInqRZtwr8q
3ZA8maGzGqqxKpPNUyBn/Nwv6nk7AzI9h/c+orumUi4uqdy326+TF5DplVp5Elo6
/R3FBfmX0gWpR6fDzrr/T0TOIOsajlTEBosNYD1uEt9sZRYbKsYbJdjtYETs0dOE
veeSfscFogixd4zRLN3ieZnNK5f19GeSJKQAo6g1qyI6Hnpopn/nDXrbJR4B3eSH
5IH1wuwwYtI2YYispEisGeN64ivnqwk9+VEz5lE900s993D0eTOnm5QIgYoU7YaG
0NaEKpOo8clk7Vmrj3yufaDLojWgrwKmUpFDkV8dWK5WPbZTvkt465dREU5m2AYY
HMbZVlXoI+ObMfa/Tv9KiGZps5P9Cq2xuWIAa58VkjMFjMnvkaxirEUeLkjL8q4s
rQ1wTUaeIfofjXQ6Pwxcrl5SOaUz21RcrQqgUKu7d89fISWkHOkAgly23kV0iB50
m6t++30D4P2uEJmJcS2ICFfG7ukp06VuhonDX0d/2SUgFzPa0wwJh57i2yFaLmfh
W21iDi0o5QN14ZiHSQ73gXMS1E4TOg8pIO3/+n0z3CVAa3eG9bybF/1d42a4qlgX
yB+NJszfpk7kwSddYBDFubqMrPTkz8SUFYv6XZP7HoPH84KLcZfTnx4gQEWgJCUB
AAZL8uPcydmcMdcQn4ktpO+CH3BGftL3J4hCHO6Gx20YmCjG5hsH6zxiLPWiOe54
nRe2d+mLQ7NWwsTdZzSyOV1AhzSNG+1g4lMdDD3Rx6oRuzn8cXLQ24+7lYUnzrNw
Lh4809BUwtgARUNWtK87BbP4g2B94kH0tKOB/3vnoqJ9HMF35trVE1MO01dB9zBe
9BQ/XgShjF3qQxWTj4KOzzNBVE/k9jHRMoDE1hKtW4DBc+3nTgG6QNywWd6KCIta
Dn252PjKDySJKZ+nr+2f1lFGvQuaYdvPEMYpUhV8YgN9ezil3dbL5GA3bARBxqjV
fJ8EqgtXLnD1hX9ZYK0atXVqk8FfLZqcQ9vVCdnUB1DvLwswLjsBt/vfAdt9z+gX
Ce8BC30sZFdyvWvxGwVW9kzGaC5L+yya5zdBawCDKPiDQrlyvGAmpEASJnao+xGK
tCPy3eNzQZNFeJG/KWfKKFqxROGtLR41SrakMoP8JRmnWWTUo8FnLnvtC5HdPCfw
7TQwh8buktLxBnkI6QqkvY5sVxM4mU77i2nyPA0fTofsUzOPL21ND455rzVJfbKW
3W3KxphmOCRQ8R7or7QvCsIZ98bGdekvxZVPu/Alixxhx2QoEcYoYqf6xcB5G9Fe
vHTaCADxdD99DQbwsFuOjC+RzCThtUjBUtvXlFQCmMlbBLPEXHcRtrpR1ERSQVIN
iPbv8AFE7f7JI0zJPmkCUAsNaftT2ZeH3etc9HT01KGDdUQCOT27fM+MJDEjAoNz
RBdWw096LKJ6Ddnf3jK/7XgEHj5Ogl5nD71kCH7iaCUfmN6Gd8R20euQh6/RTgPi
3fWUjac5iiyQy9gD2RrIACNmb8wrt+YYroGi92pALOSBs9WoZb9FFARgVYO1AWOD
OE1X3IViZT1yyw/yhPFhpYn4wdeToth+ZuQfP0kmc2Lo5UzFcQL8sfx50LP14EBW
NGGBrVT5IbZD1grU65GERG3gZMp9m17Et3QoxqTs8tze01arThTLR64FT7helAsA
YLrjN4R5g1GPlMSUfcfVOfsNk9qw2Vpng3GsC0/sy+wCl3mBzwJ08sWAkNpA00l1
WMm9Su4Cvj1knc+xW07HYrDmH70QvYNX5ROj8CydB1U/OJ4BuOJJ7K8qgRZC1Ymw
dho7aO0CH6eZvwzaARmBDE0BuX9xkzlJFIwN9EFjapuLg2cv6L/m31OpUAr9b3Jd
mShyiBMgAqGX6jIbqxr+66isFhxz54kdWvLd7FXINN7uUo8hmqwypYPQLAxbk2J4
erORv4wE496kEB++LYMc5+zpljZ/YsJxzJIpqFCzoKf5fuq2OX7KLeIyDv3fanTc
6cZy4DdsfoWefMn8HogehM5BcUggodZQVMhJMPE+TCUMLLALa6mi1u7fpZj9Dkpp
u1g38nt+3PVnqodNCxFlK87+Dnp3sT5rauTOvSDtohqNGYg55LsfLokzQskSXTLo
hF1QPYKc9UA+J637vpQ0GgspVXh6xTq5silGPuhgzupqtG/XXIAjtSCKsrCJpnax
uRCCv4dZZ2E4UYuOhoWWd/wHrqTpOvTulkM6XtLWk2BYA25Eah8t8bi60ZTUdAJX
bxGJGLC1A0WlloRN/9gQ5qOdlEhIN1tlgB/PbJYsjBmyQRqzyImQgb2JxPqmldtg
/kaPF1px+GEYsrAXoPpzI3BWRCJSC1NLEtdui1STZtGEQanYdo1cRc1qgxyf1Xgy
RTlGyimiY1gLnd9J/yIr0UWy3tvJHF9jUwGh7B6QYZkl+whe+SqETB1D2vW3yaRq
m0tzBFp193gRGYopfNyvDdgngf64iVDLQYqa0tJaWwoT3H9mmxGtmbysTgKUTfiI
EoUgm8x9PeWR4ry0hylB4k6eVRQWop4MJ+NJVo41jo2FzkE7iLDZ57CnueiekoMt
BIpTuXi68oV/U4WS9LJBgkvNyP41EtUAgJcPHzbEYiKY/t4RBPaZq995ZlLl6UMZ
mRuCVDTFiFmAiG2WlG98VgfI+Hor7rd4TI2gl792xiFlBttC9p7f84ctUtuBXnLv
78oJ3IZamwiNnD4TDeNlyRkyWAb8BkzFN/x6K3ZlviLjT57IM5rVciCzXpeqNOJu
yE9cOdhU6oVDEnRrmzk+TFuteCZPXCgMlvZTOsEL/5vBvL/82YzJ1ogIJoim+SWn
DEAPyL+CWClR1lM8ETpoJKtVc5gedI8QR3P5Sk/DxWLYJ/GyVSaDEnRn03I3CMMM
M0X1Cr4gaVz3lz8SMgwdMo/hwD7311wYacZYrQnmDylXJmQAPF3GdQnHnO/9S+Gd
xGDCxreYx6DQ2pfR1BTFnhEkiJlg9W4nKxzekGDx13cDHZtdbnObF8We9+kMVmA1
Rgp8uuyWWBNapuP78T3IJaCWvmmLaUKh5h/Su4Jn/VLaJ+Nee0n9hKynlX6OrogI
tYyeJCTdLs5LWTxim5negqOAthmafH+7M2WyHSOkVhzoZHELBgqIVot4dJvidKOQ
5+KlgPjdKTaG69tCeleEM8P61AqCWWDYxfPQrIojWnHAQwMs8AhPYs0jxOcTocA6
dCZqQiiAOdSLXvSIoycOUVuE5j4gzMgeO43zCWMxH49w8WZPCv6M/4WFoFV9lCTx
KdEjpLBDiFsD6TAqCefDudWq1Ehg1itCG3FTAp11ugCckddcRQtCQIkEJTp08aoU
jVpwy2RT7G9Up7m4HhNCFoo7G341tgGQzZqS7T5ZqM8eMRlquiVmJ+1O2ndBB4XP
99OUCqPuzjT8FerJN1XkpYROmbuckRu4MYTw8EjMQ+Md4KLVbb/YNeNfuipde9fh
kZUSCgTgs1Dlj0+xJVC+mmORbbRxll3YXzsn8dPioMMzSmC1xK5Fz1DeNbKy9JkM
i+o5NqqOVgx3ruDjL98T+lkxTJPY4liDC75//zfWIJvBFfbCP/ETIFQjMcU+A0W4
xPcDloab1IFUS+wW1874sd82lqEQ8zPtRiZqRBgE+BhfdzenqGEncv/ShkjJeOBi
tqocfAi2ExqKkj2j4N8DPDvDtthEDcaUwKVgwqlCCE5PuPmLZrs/oHYLv32Uz2SQ
czu1PJ3KB1SiDNQ7c/QLkmpFPIV7EUsskIrD/oe3KNO2hZAFWPJC+Di5ZEjz+a32
PQWRA3dDNBHn3yGTwLhD9/rVlZYghSY0tgk5XggGGBQJxzwbFs/fjY6Bf+B7XoTP
FU2bH6osAz/noYqMBVF1kVzomgNw0sN198eWjLEqhqLKyX72YeZ+k/uwsI0crMOD
K+6nkTeOIWiFNdzVRs+Bt0kioH+MPJPVLmFBcyiiR6EzvnpEstWdKWba3ovRaRgD
7hTWkbYZTsYyNFhcl8KyBxgtLfrJrdmN9H6KJKJBgV90kIp7Yq1F8nWalCqyVriZ
AGbMrZniPgUI+7qZS/fts5/6yfDSjNahQoL6FdTaFe22FflKsctKES+jga06ufR3
kX7UPYB1S1llI8lCBPg8dlp83a3pXJQtZ2Tp1GvoxgvMyWfuKtPa7MPsOZq2ySEx
SPqo9RfKCgOYYM+Rtsxa881DgupPkXz7D26VVdVWusAy2anhQRlQiO0mXIqjcGm1
5HBj5eBIClwb1yl2lgKIO+GvwSPbPkzi+9ilKiDwgRUmuJkp+uTAc0MKIMr844Th
y+yAjKnx7DyuMKwSIrO6Oh3Gna4ZcFUTdwjBh3JV2zT8Rw2D5S3MMBD95914Gazd
TpvBFvoRBvNuWMkgCmRJIX1hIZBuyGkpSIuI4OvXn0TVy/ThQ/j4WFcWNjrJHenf
+dDOkhBUI0KZ00EoUsOmX4S8bLYamUhkmI1uedsOEK5MFMG3JnfaQuJvYELJGOnI
0xhvA/SjadlkU4WAusJHGp59/PXeSz9qiyH08ZZPcXDBSsTa0k1S48Ge1eMowjLr
xcoRahMKl2DMae5dELR0VJA5wUEYpe5mUDwfKUxnfMu0X5LEJjKhavYBDtp0Lh76
vSNpni0yVN6bHetRfKBQ6ewWEnwA6a7a0UOMwHLex05Hh4xxch8ExwUHvPzOBgmq
wnK8BUGmACnWFA4xXP3/fsoN/EvbIBlcw+Pb837qwhR0L3U8M6+zB+Pg2+R+eG/d
2KIR0fOt5gJykM3Q1RgiEbP/xXaLzQMY2hwcTJNzOp2YXwMb1ygA3BQNtgdHIvGH
OWUhAP+odEt9N8eIv4YFsjz63MZtPeoJZ2qzYWEjcGKn0lDQYGSCZKqUvXIAHYnl
dYSj+WdMGjkTZMVUAbgb0a+nklgePfux8VUvC6NgYat5ddoJ3oL7XR5evhMRAhpS
OC+5kOHcuih3veALhpajeEgR8jgpvBu/mZHniUrzsBsjSP9b5OtWC7+oHK6+zbjv
h1f5hVXZ4F+tOgVoTZObdx7Cc/PESe8CM3WXacXTdMI3viKALPsy/yu8p8A9TdaL
BP8cBsWE5RgfhqGyArBn/AuSJcyb+JbSUB3PYQHymt6OL5lEs+Gg61KR1CM2E9B7
HEcdgNtyHhe5uO/EKdrZt+W3TF+25WT99f6Srv2a0UZULDv8EVxvFq9yaT/BCc/U
zpbgrr1spunvT5r8iGSsS4PnHT9HpV8g+HXj0hzqppVoMiISDN7H+aGz9rXHywt5
03uGOP6da6XXBzMQpnJ+fbpliA51fF/X/XyWhHquCKVtSigf213vOMuERnKCpcSY
3CBui4hTQRdxhjFQG6zq3Xz7gF+RpP0UImfUzstCcTKFb44pbWg71fEv5d+pb2bV
UvxXgQiZHRu0KjpM0L7xMJisAM/JJcfJj09l7xFlDbBwz3PEIa7FSjFngjZU1qCJ
3OThfrluxq7fgbA4vTMB0GA7zr21/gbCzSxaBhRANo9jEfdKAeNudK+mPjtKC27k
Rlg0R9qrl5wXvKrHAu6Y1x4qB6fuUb4pWw7AnlpobAe0huwmsW09nIxohefgS+2x
v8AVwPPpPtMtvk7MqsTvg2J7aa9GpCMiVbxET2XndVhFxlYF/HQKUL4qwRM9gfKa
l9mCPThgGgyHI1fnDm1FlCvS7SWsdSFmiZXEyoqfHt2P5fjkGzXE0CuKl1/59YHI
1se/x5/jLEPmgkdlbzj4rSotvCiDMh2iGQwOZIoT07ipJC3pamrxgGNOrFOJvTRU
ksRS3p0dxY2XrCYVCO/iWi6pmH1qeQE6H7nWk5t6oD1LzUh3ytdRFrqZsk+UiFgO
H9AM6w9Jd+aFi0yGC9eBgwSGHMBPBk1mGD3Qm0PW3NY9jmTz5da1ZgA6evkT7I/W
YGjdAySXjU2lssstEs2VhEwht3hsk7CpWHqhdwkRtDQQFMGJY0tA44E4XoK2/zIp
Ja+igrNyQJHZo0k5EMy9rmgsFdt17MLyOxAe+GVfEaE2cx3jyKhw/HN6ECfYw6Sx
aLHvMzb5EFS1MApXy/XUTD6cLX4kF3ySNunJs7haPMEX/S1ZjIcEoalTz0F400DT
d5pwUUQvujlAHu+HCMSTnf1beSu8yqduu2CfTk/oSOQmI0wF/9wyMYSPFwVlF+qf
diOCXKPk+N0h13onX/JhorAyPIyEomyZ7fdYOHXd2cArFAxRoY3GzKsmdlj1mL2s
saNthRzg8adHCD3tqKXwr3NSZcJXJqdScXDGs4/LqpSKRFRlSu5i0LSM13+bLJ6Z
4jKlLoQmXtm6zhKh+ZJ2YVitcIX4xCfimwGcQcPugQl4tZ9R+SJU2JT2Q4bP/pyE
WOFwB6PfzNCl4Wa3YTTJCaNY5eLMELXyVOvLO9HcBvnXzXuqF2NJac7IYN7pJtPm
tMN8vDO4mQGHA22Fytji1balkOFqxCundYUNvMGGePcFUgTnLgefwtkNwSEnexQD
0GPHFdxjtGJbcrToLJwKfonTrWLYiavs8Ou+rbp+DD9O1I9DP3VYlbhmnVESRi8y
LuJGE9Q+NmYppr3ETsZy7HfxDtka60Mc2uh2VkDY7AQryxrDHTy07rJZsfjjf5D8
xW3jSH8DD20ayZ0epCtPS2E0JveFsRTZT2xHYdzQiZO991OryGo+pfOBdCfi6HSk
5nLhrIL+0YnXfEgOs7eGJ6dvAvZ4baJPJdzwLpjKMkY98aL+YQ2INRwlr04nEcX6
BWX1nC3WVHHhKtEHZCy07dRm422BRAni+Wrlks8dXC4yxPhSQfn3zGXIB4lPg4Ba
THzgajGD1FDcvmblh60pZbi2Pvg954VRbFu8z72x+daiMTRDK9oOR582RQyN1wsF
khc+sLzPwO1F+NLZz0tn2QxJevWc78zDhdyRMFt9+z+oB5sDkXQIeXKJfPkjTc48
2V+tdviMp0OsTMzCu3rfefxD7TugN6+haM1GnW6GBBPQMF0iWkxBMUyjJcN06laj
k7FHf83ikdxOu/PL7f/5UE6rGIoe00YZOrytp5vxH/DEHk9PuApvo57BZ88e9I9+
RKPnAOrBshwB2lEidW55O4uEEuLa1fiREwMGWZk96MjUYG0MPXMsXlqWvoFJmAO7
1xr6JP++CQx3sHS1iF0PUazMDZ7WiNHz2Y2DjyLfbBnhRJAuVA0t8eYVRX8xtqkh
RBD1kNCssFh5cgy7tOSOv6C9JuWztZPTViT0pkAaDFU0EqlSFLzupP3C8IAqamCt
VBNAN7wLiqNMbdJOHd3PP2S/mc+4pVc7ycsH7/0ISe+CfQs5fxlAbMSuPiQbzSe/
LQwZnft6VEWlP1uRsU4AMvb9W172W84sImLYGUmLvESpXM1KkdZuFPev7Qx0W5t4
kRsQUugOHbr3+yvHnantVcVttk5pIGZUZAg4zGymWJ0JfY4cfVLtqjvjYEP29jnJ
9+fLVnBcwfhkgqrhSnreMYiyaoEDdYQWF5IDFMUPRxbRlDKtcHtslJeIwdsupT8O
TEolj7Q6wBPqRuAUoIdhRSGeKPbruRmjEEuqH3dQ0C5KWC8kvEcj3Ukk7YnnPZpz
0cXcy7kyVZDUuExvW48ZH5tBEmobIORSwjjSZWZLKqvhCrsFStf8NyKKeRZEsIGJ
xx5HFOq7LrQnjpKXTtaBmxcSTH/5C4bpU/rnvL8MuDz3REMbQr5Gws7jlF79z5XQ
neV/YFWMBFyi6D/BP40oD8ohsgiSsdPbgItyDMFas0sqs4Nwy2iGl2kk6xCMt5Z4
5r+/i4VGKoqzeBuS4duce1XLHGU95LqYkIrb/LUTVlVr9A9yxqFCbjanUh0VQxPl
y8yDWFryeW6OX4jdOARqR7Yqi0JX4fFisj4306qTeEjWR4N/GgC58618A0sGf3FU
kP0GmHSOx7tCAUSLufjFKutOxPqOzkxp86WVKM7gQp3LDswAthrqr8eqmiz21xpi
QwdEAB9NvRKrW7zPQ86aF4CFTk5NVFTqVV5lx06lC8JVOk2GgweRhsUB3J5ujAfk
ix/4nl5nImOiuQax4SIvxuP1GaCcEnjPkzV7A8o78wUiITra5hYeFEmAzf/73XmZ
y1KTEDuhoR/wNQRUnTl6aCCJkxxRMODdWyqsW+Fx+7OTAgOOEki1SzCvYhryXB1N
LZ6PVoy1VbFWNfSe2XuvefvMVOgPAvjXGbJxNe+q+YNPCNG74JLz1QCqTaxWzH5X
FzeD7zJ1FmmkUPVvsyLaFjkFnjgwTlDpADgKBY4nz+x/4lwlbbPUwUlkGMjh1bOP
wGvNKZFnIckJbqphKhw3ytp0L6U1q1xAW2YAatN9pAiKdldLdYoNC09tk2EZedbR
Bt3Ls2FkcgGYKjis5Unmjj8cEt20PpV+8KUHg999vux0VnQBbmD2s3QGgSTnx/LI
ep+ELy7IaPN3hFeEU54VkgCEuuuZn3k2QfXbmkZDc7DOZnlUpHWafVUC6fzq1DQW
nRIV1uTmjBFwzt01r7njKjX9pHjo+i7RIOJl9vb1tzsUSiLYcuQTG3y0HoakJQXH
kwPJNH6de4ZjfZ/W9ftRlPMgbuRXhmlckC3mGh9gDpKQvh4y7QITk+5ReBztLYIl
kiNR03O7PNpIHvDXHOjhGYwyBApxgQGCQFIlaiDqntfrZlVD3VT1BrI6k+bnR6n1
HPI9n7DwRwrohXJfW1sAsaKlLQ0RXxDTab6lVf2wYfPZO0Vb3VvquRmpOVig+vj6
5dQHxA3T9YywwPY5t349G9V0Gbeu2jG6nbum4khon1LQz7IV+6E+PR6b+Rsb6y0D
t7SWdYheImX0VGlDYDYsiDnTohAXtVFkgquujv5BOCBgTpDZ+Bi0zdfYQmn7OGn7
GRdh8/MigRON8ECl4JfT6aXH3RnlpzlHg6nTm8VcZ8Mtkhm+OEZeQIKbbPCigxvm
V5Bn7AHYBSKl90i+MR09dZgNHw3OUiXX9EqOrAdE/ebefPpYYCl1QfZxvUHWDAGo
yN6gCItHY9bejg7EUkQZbHdaXn28c+Xp189dXc/Q8sfW7MlI7oOv+u6hfMbIeveb
+wDk9lpLOM6VfDZ2DfWE8KWXYrhA/UEcw2+BGFaj41e1Xgtx7J553YlJxGzULiG3
YxXmAV5DY21EyseN9Vu5BTo+oP0QBYH03Ov9O4mS3Anmf/TiINDlfcJOnQfKfBlv
iXFo0Nmmrb72G4hlOBKrulST1AsZ22y+hbEDUBK3iD74aiFyh+ixVg8L1zQeq95k
PiPTC9PODCpMnUnSKnIJtNhE/MyBjwstzBXdaJO0NxhP4uxNbt0t3l5AZIZcbthY
Iko3WMeXQBwEMY1XZ6kOzKzDFtLQxmN+gCUlYRQ3batDSkOy+S3YevNAb6ae6eOU
xfEU9a5IfnXjhVToIksZ0v+t75gi+hSLDTrubJdWa79oX1+aN56CRIvQ+f2xxSOQ
W91K8wGYIScFJiCMVcqAiQ3JXSBT0p0hy0g8u5Z2xrmgox1HqzitVoV3zQEWkvB0
8LAQtYdLtp1LLWbW8s3lS8P5KDDF3ITp8TX9aFeAyFvlXrJ6PtB6kcOxtGIq00Oe
TPwFlaf5IHL9gnW1cfAT69rHyl/XcwHoOc2UPKGCqM3YEhGBGY3c3IpEmkTys79H
Jz7dgykOWggGdSjotfIsN5FLlm1g2f0OPgkYQ82PT4iTBcnuaXm04qpi2EqKsd7/
BTnbmfzpxveZbOx2y6UJ7jtJRc3WcPNVyruw45kePP4+c9a/BCQnOsQSzHhiALbf
ssi39ObuL1Gnz7Xm2dmGHVydFg080sAm7RwGxVQMy12Q1aLbZJ34RS5TxJOG+gr2
FBFrVKC5aWfizx2C1Z+HX02VzH9bD1P5f/kt48iz001M9AYlghjLn3bW6ox8qarE
HATcK3H0/wdf+FdKAgy1yo8laXr3PsZgT38eK0bwShLujd7Y+/Gcl9qYapeLMuXY
+tenapGx/Xq3r3nnHgnaQt20p1fQmiuHVqr1jO9/SRCN1A74qGbMmWv9XkXK3ppo
Sb1zEhxpIPuKbWv/9BntF1qaeTluxvRcsgif82NiqUm+zvKiSeqmE4YJqJzUembL
ZQTaVEISdHjvTY0FfaWYCVN8s76inww5yBp15H/4M69Cd5SYo+AK7+bKalAI2EHq
zorEZv+y+Ohx4KzPT1YN9ATJgzb7FPiwf2OvFa6HnWVw08emGoULuLtQyCleVJfH
YDdprueGHC4KRndwQ4//sGSO+0pC8/2f+Ex/HX4566OFPYeCp7vjNr7rNr0mnVbJ
s9cLA49E3neAy5gHzbQX1qNjdbXMyz/CIhi2SOrNfHkBpulDosKKyMU54TCMCwGa
jXy6Mqz3lW/vF7pEgWEn2fvNkP8DN4VELlPsS+KUEt0/rVvBrLTi0/8c81O+Ti8J
Tm8xNvDxmCOhifyRutxIsSD0nRm7qTBSw8J3Jzsg/jWw2ez0WRWMhivMgvYIZ8CP
qV36VlnbaWN1cHSyDwRDtdGCtL109udq5GJ8v/XkjKkagDIEmA1YjgmxQfuwi/9b
G5AVvainQTC4PDvDvRhfzJFae4Zz3y3wqNceOuZk6pV0GD0Ek2GX/4b5xEdLUzVF
Bk+14fim7H3MRBII21AmJVoSlhntWha4Tk+sMEdCEM9CUuBFAwOSXJEMryUXWy7J
k2hqklmd1c8j8hVBuQoQbik0nfWBH87AQI0kT36T5HE15WjNIBWj7SEhqRd8GCSP
a3s17gFPtE9vQL2Y45lUc0uPOVcfFwxY3a0dhJA79lAGXdd+Uk9NaabYIF5YgFZZ
lCvIL+YtfJzDzfoMH8y7pjcuYR/j25NT5fuCF2lI0YVp9f7zI06QDlpB76S6dUTr
/NwMF0nvqOxKZFI+ANRjeGJ+jWD6LrnapYNrfDOJ/D4WscPk/3i8iMyc61/WhcVg
Of2UE+prisXWRX8soyFFTZiRFKTO1go8Md6rmt0IzWw/QhnzRHau0drZyWwf5xQU
EiAjHP24fBSilp4ORiur3DKFLNNg62w1ngDhyZ5qmGGfoq1ihE+Fchh1KOd5iWms
kAtV4wIcWvwLMIUlVLsoaixrh9kxYYSbB5OiCTErafQ0ljE2k2wPuZBxnwhcCvSh
c3BCweLq4OcO1R7XMqrEE8HMtu2eW3JHd2AHs2L9qnEcLPfx9ZiNa1NqKo0d7oFk
Rn+0bM7HusbMZ7Y9Ywd8zRwyRcCW7WvZGc1unxTWxFuNxzj928Dkp1yF99ls/s7U
mvn0djEa7WWGlgnsKuphubu4iAnQSYrSAByE5oD0JqZlJf3/jHsclSWHow8LJ3VT
vMNB5s1VcDex85hGrsfPsf5McqeEykFyqlmJhcGor14RA1r+wqOpzy3q6S8enXXw
QRuZAMFJ+YU/3DHiGSfXpw4CXMPySrW9Ei6rnBHgMB7QYWpoPfD/G/3CNkgeUu0Q
80Iyep2JOQz+037TDCPv9PmWU8DBYcCaBQyNvXcoOFrBZetm25qfX3hnCHlOdGPa
L4j2v3CuotY5m59BdI3Wbo+XADNbAmewpCgCEAolIqp7HgmM4P2J6O94q/PBdngU
K7jP1AhMULd986n0ZK7ibeDNtd4PP1E/LDg0t9m3fnaxojECOx7rTZYkMwIvlxTE
iVxqGpCemzv6D5av78gucsW2qfA9pLrbufgCs2YtEW4k5nAJPv8jFbxbSEDfKjX5
AoecZv1af5XWmQbBHTX18HZkuqQjOEK/XJuRB2UBp83otx4/B0uIwoyVBdoISirz
fYWd4H8ikKBlmy6+qI5JITEsu8+FwwRoMJzAWK1RVxXACaalXrZbMyzO91HwbLek
JZXSWF9vG5iwzQo/G99fZxEQIvuk48A0ubXizAByXEX6/BZthKfPJ9N/VnhZctek
S6ZCsOA3VGVzSf5ZAQ8M8BKJeyx7uiZT7CkHvDryWVrLIfivwFgUK5Xuu1NOE+Eu
a+2yfwzQYRUiXbd/2IyTKTHl/T7tSzjxEeSyM19dRMHo12qeWhksKZNSOHx2AlIi
V6uoaIU/AVmuYLCTY1LgQyEiBkQhzWQKmOOiDaHokzL6sJAZOZZtdBttkFAvs+VX
aMHaCtzWShaJ6phHw0SmVTrIVAfYLF7KqdcTdIGPk4XVc1FDNMeKqDAN91ULJ5eq
ZKoeG8l74zYw1dk0izbNbh2wbySot5uMJra183tZA1iZodZ5NhXQ/9IXxPZPqQ2G
AuNrecQUZocgb1ABMqde6Fqk+0WHfR5zCf/WFT7swqVUliAOFfXCtsVYycLb94mV
SqYLSbMKynMDiYHjQPQsdLI1D+mWN2REsygULQ8q2ZsGubCey+GnZiRwt8GHVC9m
N2mf8zvcSrQplldImFokHkutwsV1JSW626SJY9dPoYonHsEhOvMHjx4zkP7Td+mW
gh7TQn7lQCif9wJ7fa2qnLlfhgF6XZsUqE9CWh0PvR/sysFHpx9kU9hpRcrPvspc
JjnL5pCX6CZ11q5LpokiI4CkqOfgJlKmd8EMcZMaxQKlnDwgpPfvJC9g9ECH3akz
XdrcHt+vy0DtoHrIEBXFngUigeIKRXoxxBVuAcrY3u6WfwkUUotIuJegBeuFMwWB
pK/ZcitWHQjd27pminSunLGlvrWSLW+3jmRAYMTOlwkmZpFqwnVGOhm+TXA9yUep
sA41F4gg09Wb8fXDPJrWXBjyWsiAYPdCZKoycI4yUwW9OguMp/3au6mYSkp+spYU
zWxBW8vqniP2eLgndE+TB+6W3EQwZhg6Lm8hnusvi162fzGNEGsKf+bhN0Km/D1m
cHRxq+xUwBnbT2sDngik/rH8ih1kIX/8HdSxDbTvxHRfqOA6XaDTXAcAcijxbMLf
Kxpui1Lao61pIgjAzi0LCCeLT14+wIhhR9iTmGeuwm8f5viea3/WnhYjBkTu0S+4
lB78AYHxWB8h1GWuaumHRUxlRJhL+A5gXJfn7d/L+aw5YPfLTxFQ9eAluarWAs+w
0/WbPrRiCVTq+F/0IKHfvHuPHZVlmNOKyA5fB474R28NGeVhOnpVnPGfwTxCEr1L
Mdjm6X7XxzSbd6A5Zc8nbXur0UkD357vWgfRL18my6llwvl7xBKQbVnFZDg+sNhR
2gir8rPF28/PCAwWGmMz5DbWN80vdmDhkmbEegaTSgaCM/lpVZj6UWpil80tHa1i
TD3HwrwWGvnl45H2nkKFqWKnul5osiijb0sU8Yy/cIiFl4PX05qnNIIPlsDvPk68
3pRzdyjidhitLOJ4AU24U5ltjfVA47746pz/ZqD1rhA9RgY5QPzhRpPp3NSqqbag
QyXOMFPmIMpJjM5bD+o0/E+7f5mIUQR4OhI1NSz+t+/VIV944Lf7gGdBkbRDPwMp
ZvGWrlMxN1yGI1oy0OQcZvdXivsE6qt+HYHU76w9MTau92wxw60F+vHXbm/gfIoD
1irlI0n4XZWTE0TUgEuw7QnsolyUA347HLeJhOQNq+o1l1war6hwEzCLN0QNzXyl
UyLPfbShQpb26snVHFcARKwDQP49+CiTCXU6lIpYtvj9ph4tb4Xyq2OUPGqSDGH2
n1Vh73/n2l9OGGH3QvWIfLiqKlQD+3A7dmi+IntpsZaqIkg/Q7aMIoDVDVDjeSbX
yNmaGoLSiYjrHB3bl6fxiwx8Y2RIvN3wMttJwr2z8GRHzxUt9f49Xg5edG4ekDo+
+nxGujKTh1Ou4CLAEvP+pS2qJACBvYUf1TJzxS34LDhT+mmX6EPsm9SnCTSRlUy7
hf+osVLpUSc7B0z84ayHqCOwPTaWXpF8c+khY/MtTkox32aERAZmVoTtKOgTjiy8
k/tAkKWCfvSsy6/XOix3s6+A6qG2Q1YzOYJlPtczZ2Gu3bIFsS6qm1aoOvRFW9IS
scEeNfNgweZumWo0I6o1aZ2Twq1QLKAXRR3G/wxhQ4dNrcQgDXHpd0jeyTaRH5ge
q62y1Tw4EPMz1coKAoPlTnFderEyXiS1mOB0DEUeT1gSJGeJ/S/vh0s8A1e4QVn/
T2aLpfd7lojTpN2JDP8opeI6r2qkV3HgDClz3bJYNK+3SVHv8exE9BDzFPRzEzNZ
q5wA5b7QfDiu5vo29Zx+ENNfSDWDLhwsGpNF9G7MpzF4HRK/Pr+neDDYHY5wblaq
JA0xU1/2+L09mbNaxxRVSzONNihUaqxynhS3eamJl1f9CLGKaYHFhMbQH3iqVAAN
sebzTbiqunQsWbnNiocF/+UqfOC1cajaZdG4aSbBNWzaeSgnHS3fJ6YH9JfC2gX1
a2uuVu2DajebK8KZlSxCr9yFYEvRGi012NplDSG/QmAUPK0uUiPd8Fd1gUui5h58
HIWVvZTZG39k/Bv4lWcvWO4ajpb4wqx2lBaOo2/6kmjjhTaHulovP82gzzM03A0K
9sPJB5YWEkdSI8g3Tn8tn67Q+vHITgJ9cn6BK/iKrdQlT1rrtMWkLwMS5LNR+ewb
Ti+t6PiCc/UgtKvI5tRY1JfywBqrkT7IiaqiyjUHOzofaxPKGoiaINvtFVvajF8n
C3HFqLLdGztj/SDQ33//TiNcrA3mvelfN7cICAoMgTh/z1wXOITJbq4L6FvyOQky
tOj5BdqW1moUx+1TCsW5fnOP66AcqiMEa9+BXAKcd8ZMBdcVTyMaG9kdzDPV08hY
w1NGqFIFCSQ5K0crlD8SoYOsUEF2ZaCU7AqkPFXBkYEN2LI2o5351+qS/A5CFz1H
M4MlAIZv2iMXA9thZg6TvqHUDw9Jrb2OH9kjZi3A0sxoH346UO6TrznhFGZ/U63s
lv9eFQWnq2fywaSZVtthKCba6Jakwul0WZCkTFaBiMtUOKChSRSQh47fy2Em0VNw
BfDO1RYo2pzwV71YPDX6MCBVjUXEp9xZ3LiT74x+38YvBAPN8YgLP73E0pU5MDk7
JL0Z+CMT1UTsLqk6yhBfZUGTIYXDbTp8LCgfsk/WNC60icD6z+LxUyt1W6H/2ryT
Ba0AIGQGZWlwGxYZiQGyYAdTqUmDLYs7H/VjxJIzB9K8vUmIiih8HHtMlzTlmpKL
c/UVjXaAlynyk3OJVFXJMCS6hdMdIiV+0zQFgX0xuVFsKgOuWF4za1nHxCWmziIf
DD9/yQq7JgoTqAGX1ZyY0rVr61Z7nJvybNzGFJMQb57WOPEZmLisEc+shshL0vju
P0HaguBWFuKTIg928kgEdLjOhFR5oaJREsmW9UfuFYW0J21xjxo5MekPx4uBJHOD
6HcYlfhjAo53ZJziwCw9kC8zjJHro9K0QhSPs282Q9OmpEmy2SWz5l4XCndWdnfl
nyqw5ZeFHRRb8dn4csaIV7M4TsnzxeOGTjnVIxvRIrHWnbyUmNSyCfScbW10ada5
CRqQRn5inbu1/4vOJiOcUYBIrFO0+BCyJWUdY+a+Ag6lBV0F3H5Kk5SAXk0FMiB+
PuA4qm02srAMqLzPGeRQArK1ldA1FAyfFg4JF3vfqsfCmnxX1mHgEQwFLT8rkGEy
CDnpDFfyeqcVEnn5hBlLeRjdNu3iYnXNQZCmTpymeHfBYuEb85LQPuT/nc3rz1IL
E4JOhhti5o7NBcCgTUz+rUhv8QRwk2M7hWstV0WbmJeurCX1o58DC4/qn6IYl7Oa
5KJEEWeVjDfWg9eTa0ziqkqpKHW0UMy/ewUxV9PoBDW88NgyiPJszT3zh6OCnhq2
+1GsXSH6lpdsZUtQGdpc+DyNLAvcv7b6xNcr5tdsRmeho+nYR6uujICdMLhYqeWc
1Z+l09MalsvhPj8rAasdpYt12de3UfSCpa4eDYYn7aB4NaXRF2M03PqWQKXgOmb5
75SiJA+ukfc/poOQ/XomckGP89mOvsgm4mUcOH6lsFhIo11YaDbZe7O7E+C3ZVMy
CxzdrzqaXGpwopyqIjFVKzMJ1VHZjctw3S0Z0AaH3usFtOZEEXQM+cRMsNZsEx5V
iuqoZDmG6ia9hvmPNOSH21R2RXt1D0n3XHOgB1M1iBZMMynCXrOrV7YwmsvOw0UD
jGlqE2ni45Vf0YteFAOk08g0DKS+faMDLDuJOYhAiBO1Sq/RKA6XAhw6HwsdXO8I
c7aVGejqLasL3ngFaUc0a1PeEI9bBMA+ueRzzTLQpizWGjeftLt9Zqo/6I2C0ZeN
zhq+McAPVIlzbRrEy1qzH9QVAFLC3RCi6FB+HF0f5PvzKmMDsi28wn4n+gviZ9en
6UBX5CACQ4Z3RUCpq4Awy4cLthXfU2SuXfxypPFaDvjkeh/zaHQnci3f/7qjEVbC
kd70bD2veOa8hY6a/mZg+yKsA+SpEqIznfSXkprUkd7v/y7EVCDzrxy+jHPhpFb+
CaTbyKhs4TD962Qgnn+7lGRjb5jlYDmtbKA7xc/8SWcvC8jpll0QuMuSBpNgUb+I
aVeehvQDbDkzQBxvH8a/uBYuwvU1P9WATfgRf8HffAtzcSt3/r5coW3dmwgtBx1D
j7y9CqDQUi5nsYlGtRlqMqghqXBVGR2AL1KywRTyAkek7e5uU2MjNrC2/W5s+3/L
eCF5Ve780yi9TQS1WjwJ7Q7+dH2ojCxFqZv3c5Mu8zxd6T6AhMxWbSdMrvoKU3WU
H4O06m5nVFIpsv+v4kEIQdhHx19dU2rf4aTUHkOg32NZZGLLe9mEgAUB50T5Aw/8
PJ5jD4780Rk/C3ZYGbJnLsZthJln4iAZyJB9kpixWBYiRMBzGS7RROORbOevGrLD
HkpreGovbjiMgn/t2SyHjdf74YHABaLiXZM6smbwVRtqDmfAcgUaXJXAYSVWRiup
fXwhnxdCwUhH57ODHXLnCs0lISTISz/DAzbCg5cpnrqquqANVJ5p8jxOdas/tIBC
8RS88C5Mtyt+omCCEauc9jhyXLc0qk9VgSCUo32jwbtnLDjhDaoGxDsGkIdjMUvy
ESl1DGCPaeT+l17hB2KxAA5yxvboW2cQWzyzffl8Q7XG7W7YELL13cuyC5qBQ1Gc
rjAvzAhApJ+5SyigmqTFzieRMymNuotnl+yyXVT7svLwWA/5PV49+/1F/8QmDFvB
W4q0kZKSn8NiHStC0j0TDgXgOjscnwrofwyW6zheGDOWt2FOG0UbxBLjeH4/lorH
pGrCDObGBpOcweaTR5d7AjB8JkBfpAeWjR5lTe5j9TM1sRJtxAu5dgbAhKRke1eA
Rj4+HnSbFef5pk3TXUgmHlSapE45ElGx3KplJ10W0VEJwghbHuUpUpA8uNUMriR6
6EXJBG3vUHpenz8d63olS1Nkix0aWf6JWk2LxnSvH3eg/nVoZpW/Lw+e0kaib3pB
tGS/XIJhecz+swaKtjDFhMtVNOdOJc1qlzvBvz+8RL0alX9atgC5RHl7dOua2zRq
iYWr8K0cocFa3Vv1qSC8UOFr0atQ5sApt+mO9+9fJNjAkdLs/gsLjg3OvnIjtf7j
4BxyKBDorv7oNy5M2zBNIHcYEg+gjBcoxMixSQbJgfjuZ0MatzTs5wZr3aa/3Xsi
48KoxgU4gP3t3+G7RSwSUm/kZZCCXfijnuGgqPY2pBK3jJJPPsBz50GhL5w0aNV3
Or5HYOI91/kPBWePyN+D20h0BenCkicT2a8/msRi5uzO7zZ/3B/0A63Q4xecOzhT
T/I2qH6z/4ZuSYELFhRcCfZLpAEnaII7gmMUzoeu6yP0MdayEvgkkoSlGGDG2Ipz
jYZp8H0Nflb8+nbB4bnFW3NT6eS2UiqZ3u4bH2udLBEnPG21mxnbd8Jy/JshTX47
xKSbo09SKsC8kx7gNYnduqa0bgorjTIo/xe4Cjkvj7m43hRXJ8ViF0+nsxWSN7LK
67C0NLJKbPeoYQMScbh7BGZGwLZ0PYCZkGllS9+uDDXSp11Mp+moNaD8T1/2AvHh
nlxEbykzvAx4IWuCWG6nnFMPlveaimydPTVhENEJAXyy/gs+wo4xheVhsC7wfCIl
G87lR1gIcrc70DmrErwU4jOFVnEshWgj7bheebcUABzy4M3SxF9OdghKQMwqGuDp
alrmEtwoqDV+pyV1/jIShpoOyFE7xInyoFHpS+pLPGqsjbmbE5MUl85tDLVSYDu5
4CDkDugqOPzd+wpkqi6tJ+QA3bf1KO+M3j6lZr8/yrKkr5Y837jhpxRp6hCPlaxv
gh3IeXH9icTvcjW6GAFAh6hLHs68Anw4nGWNym27LrOU5Ny9GKXaxVpbnv3RIXoX
KgQ03k9DIbrHnpINgBfk3o662hgpy+tcmwaLs/QPbhjENdc7S2KZGi9nfUDRY692
TtS17mkzxBfxdwiQQXWv7vDS34sVD2pI/1MCRVmfbQQ0Zx6B/ERLS7RoUF4MizlZ
jUJV3xzU2c2FzUHMHNAE6Zs5iBkuS0i8IyuX6N8v8RDbW2A0xRcySHfJuCIwUxMi
/rVGiAp3PLGB8h+brvCWWuWuZBU/4JJvf1xJmK3ZMKuluM7m2PLkwzAwG/9MJqMS
i2z4gnndz0vTAWnoKp1cPd87rOVp2UlnTZUI6pgyHUTR3aIPsAUPQUNIghHjfm4F
cUcN8YhGFupomuSDJkO8jGajZMdKsu3dhvr68ql1zGSWdHu5O8b1+V9e7OafVXoT
MhDFcz2BnBqRw6yeOEERy1cxyOb21Eq4604eWDloww3cFyTMhQHkH0xf/4Dt0jDV
+cORRRoIWOl7nGRTsV++Rjgo4894o6OBn7fxoWZ7cfGNnktXdMu6xOfT4ltgQURT
MY8bgCsarhoxNHK3I+vOiFSIanm9eCdTJfV6Wt5H6pslW30UedbbWdYyRqYUnmlx
itp7ljbzNtnodyYVj8kfti/NPHjr5yFmFely/OcsAgP3oMaJdxcx/VBgWMVjY56I
gnENvKSCuFHfB5qm04jf0anX6mvCE07ZuSisxceEAcANHXcK9r6x51Zn/RM67JQJ
CawMQti3uzssc+D8QHXHDWqZw6qIms94T/7njvryggj0AIkXK58m7I2KKzTNlFW4
9F9IdY++F7G9O3YePBxHp1LzHMQUY9FsEloXknOwdv3IpYu+pqf6wLm/D2vmg3Cb
5lDXl9lc4Kn0OlvUpX1/o+gPc775RGExWu2qQzRcyHjbLQmtzdYKsiwkBoeSD67a
qqjj/5K7pqkC6ghHcCwkOBu0oZgmf1RXb9DEld481XlrQanLb1RyOyAoMHKUOjXz
k3k8xuEiDKLrFpV/2IRD1UUOyw/XUDlNM2RwyhCJQLBViMHF6L8f2kVDz/ZOvuRn
LzHn2zjTl0SE4pO03SvOoDULcIF9LEYheArRZ4xe6U8CDik6R8kOH+bDxg5dOlKs
JL4SLKZTq4PitaqxtVsys0OHOpBXlBUNI7fxvJRrnO2Adjh2qnuS9UXj54NzMQiD
VFp+FGQQMenvlocbiVPAZkDOwgALufnpS8xaCcizw8aUQrF/FYJOJkVt44DTQqLk
cIdg5grIJD7dOQg1eEnc1b8IjedD2LwrhGVWXDI11KKzDeJOYlHiBKPOTo8yPrwT
kswuGyDIeT+E5xBh2bWcDULG1NQIQRzLb/Bufbw3ZNUmVuNcx4h2bMbuiAp9y42/
8c4htrrzXnG/sPZUt8TuT1DuHX0sJ4LBXPIKW8Ttd8+AC4VJrzY/yg2kgbOQ6dIz
M8k98o2B+M48GZcFqcpRl4CX6/VtRFG1WQpazL33g2YhVZrgBbK7GiBNB09VnBcy
ePewVtfCXMt8F8oWCjaogSkv9iB6hR27VxCoLDvsvPOFkqZPliPP5ccI70BpUlJs
vfzBdR8dOLVN9YNCEegoN+2oA0KQYnjAlWssAAGUmiYqqV9cI/QvRNU0ZXvFmkQ/
I1u/2Xro3HzYup6CuM0GQ+u9icYHcUBPGMcP4Lv6ioZFMnBJtGtw3DGgl2ZEQYS2
KVncf7FvTOMGFKQMYCeuPrLkc7RFU2kNNCIKn9TSbXtH+oB0gr0O+DMkIfWdCcc1
fhrCgypQDe1FUHNE/VZJ05OpBNz/h746gsN4MPx7h+QpNSHTzR9saGudIVkzBh0x
KvZdFYEr3us4xdhNzzZcvFUOCS17/QNVPeSs/Emzzy2K3XHYesKxjZEaJlL+7Phg
ZipD3ziuGsbTl75I41zMWi6kWVkV2s+GU6yLimD6yXi4TRA0mILuZqlpg1D59qmb
FSyisv5uZHJZIvMRaH3/dKWWvTF/nQHhEWa1JLFNs9SbCGmhKI6wud1TFQW7RR8+
ognOehfHLBEym43EoLWaqNWxGk8dnYs+fWhJ9JSk7QiXH6O1KPPlkhGuRDaDKVy1
le2vnuplt2nQjEQ6DToahDXhhmbdMKl8LNXGk3R/w6COnrmYs6D17iTOWcmX+wSy
VtB6ctJRSpGZ/3cgX0T6yH7kGyE9bbl8zMZZiUJQwY44vijJ9n5Jy7PKWzh344ci
eQO4b9Ay7/U1iEh7HLDvW8aaWTWRcrUK27reKE7fa+JM5a6BhD82uZVix85ucRj+
sAjmsoppKvFUy3wsKeWV43I21o+/PXOI12wB1XjMpwzeWDFDPdxVC+deIx216Df8
dbm4/cCuyQad2vDsqEgVSh+fG/ivjNaBvFFBJL70+HVsZbN17AMK0kr7XjLAP1RH
ZYVnZQ7dtvypNcNkXQj9//wtTKsosiEwwfavYns+EsEgXtBPeMUvcnMyVteZMk8/
RZq1fTdYwblXdTcQ19DeC+NSFOccvQbJlOFGrLeaQGUsXWDWfEY/WN+30f1Cu/wR
S/K62rDj4bivu2dfJAsuLNI0fY3d1x4vR8UtgAN6sTrIkA5hm+NGzJfEzRksDUQJ
+wkU+NjsPr7CYpwXZ3YBGo1ihigmVqgvo+n3wyWZE2nTjmfyMzlRghoPlimy/OhK
cm+/iRXQyyw4NLAtcGTEBaHSCdlJpmypvi3MXCzO4sU9WqDY0lM2H+39dU2d1X4z
0g41MWoJYXpC6hbQakdLV7oqyYipKhsE7R2h1UMF8BU0ZcoAYG6gm+Bshe15nw2R
5YiklyO2wrFIFkhjneC9JpydgVYojs8sqrn7RlbP87Lq2ZynD5DMB+RrnvXDPBpP
QP313r0+AzKT4tDRNtfMZWPq0s5wUEg9gzmV3s6FX9krizMcvZmisGSBnmV3KYS0
7AFw7zdT6Bx023DiAzXHUxUSkAmy1BFhx7p8DXknQHhYjZVEfqTyXZ46FxSCAT6t
+NqDbOHBRJhWJTy4MDbIFiok+BcCOwv/QuBZD85bcQb5IwNEVdtRzXdQo/OY4asP
YVJgjG/kunRo4OKxDaDImyNhHRJf1GqtIDKxYzY1fnvpcJCAsnRfIZ8dSpFFqnxr
LBe1MUqQlaieViGiIuSW/XHNVX3uaGP64/McWegF9UNmJ7FJLgxBKT3p4/8I9Boh
BjONIxPfcIxlVESvpPwN+w98G5XB+e10bGYe2z4XS2d7DO2Tu1utsgwdBj/R1Gz5
srtmhhCjJZl1GJAJUe1YjFSQQTh4v5hnRBF9zfNUY3xUfI2IviNnLL3wEolmKv8Y
rxFEas73QXaRNPbNgG9KHDDEESrViFneVZ/g55JtVKzoZV+Rcu8QLWKEmKbrPbSq
2bQQCt24I7YIhLQFFSSRAveUmDL79GRNjlrptOrOHq3Bsx1xiOcGFn0oAQUPx2Fn
ba1vSOuR+nlav9VXCvlFqj90fCCBjfXwPLtT3Uq/2qWdBQamLMt3JIESAR4p9qAU
oYZ29u3JVGmvfNQuL6IwkmDj4BjrhbAp0mLWTJHI9Tk3Kj1Yfip5htn56xoggDT9
U1h3+dx6avh7b7iaWPJC/6c/CWNuZLCf2b8Mg/lWhxLb3xger2AcV5lD0UJwrhzp
yaRDO9Zd6EtNP7UfP9+jAsn/5dZg0iAVe5nWoVHFfRirOAoJ9QCj/afuu9Tushhh
3d2UZ79W0rtaxzTSoVmeB7U9A5Hr0snBcovN34vPDoZO2VxXzy7grdinCwLqEUN8
C1qODI/waGBv5PJEGgbQR3JFQYjvCbbZoUjJNvVSmh5ak7y3NPydpl+QwCbrUG0u
Z86L4E5T2JtwZjGYo+uhU8+19ZI3MQhWIeIBjuEy0vOMSGI9OVbcfnEDm/0o2Sb2
MGD75tSod4D5P2NbKvycgqzazg+fHmf22piXaF+ROPHp3glIDJdLNXZtmgT2nw0t
HERXn6InjcM9JHxlxfFPTfR2mqGwt4A4witWN42NS5hgQX5O3luXONlhuuCdOTn4
cfX3GqyJo/ii19U01BlOERKjoxa7qZgUy2MYGz6NlhU3VXmBunIU3ICzEN9xj1pN
1bfYclo51lidTliuF8b0uPuW4S6YpSVWp8kAaDzEPHLl/3ohQNbhBEx1v6OHpuCL
Iefcw619d2u1xz1+2OqNY5NzM0lD4ltqxwi/LDey/YLv5ZruV8wubVGw8TDZ5G0w
qdXTc4n9+khxxshA4x1wRQ/EfkYAR+Uv6CxhjxfbK0z0LEzGgKwCTjX4OZt4kFp1
IFUoJzbM6niGzOa1dTTkpMrbRslQzUUrsla/BXHSDYydD4dm9iCb9n2kpe+UoA6o
dp0sNaOzR4Q/qAPbYvM6MyP9p/CntRVqIGVRKdsjsNLmieaEyxTVe5XCHm0v/Rvl
vdLmB2O5ZEa0el0xGVXtxksxsEpo1gcgU6Nec5f8YfkuEIa45O6/QP0QGALYqjO3
MOd6Z1Ob0YcpIiaYqrzODD+YcKeTZ36AbrebZdM57RgbpaygX6mdcQvTBQOl1P9d
NqkinkTYYr1WawyUvKSFOhk7PhUNLKjFRZqIuy8HmptS3qxELfuuoDdD2CkSOhyt
QtMeEnqgD49vZQq9og6Crij+h8VRGGQ3jjaUpW51hIZk6Nrx2YDhbfLoQjvli3ZS
ugKdxPk54c6s3Is0af2CesThvwnA4ug9R9xz7z029MEyE+gAGe1/pfDxD/T6YcV9
eROz4qSzR8wFWe2AuY6UXMfkltCDUPzR5mUHsY0a2OOqta1ifMLRGB3tpVij8loH
j5L9XXTbageliMjc/FM3ytYRtdQqJ/qcZpLltUvfuTvfgGbq4iK8jWpRM05346T9
7JiCbkiyPsQ6HzGAfoUUXXMic4NbnWYEJH9Nez5eBGR+FBvRJW3yUptvQ6Xz0KrJ
TwcuS8dJlzK9Oc3WrChrZ94SvTd8sJ6svCRX1opiKmNcZHLmNCfFLZbYQo+uj7iY
2Rocn+N16ggZHkGpb2ddm+rz3zxQ41xDQClwHP4i98tbMROuJK9iUC62hKjVbikI
Ke0hHnPtzpHeZjYxoGLkOMGQxL4SvSeVwxA0JTw84HpsHPB6hruAz1arGHnKeMTk
YAw9YlFRWIpSGxT4CeSKjFPaTcF4gL/IDDF6+ka8KPeNeOF32bonw9Pu2na9Pj5N
1CvBLdxL+jK1MVpCUMETE9k62nrswsBOXSt9K/89bXzfyygXdAlB7Pxi6r5fI6Dc
rJG6n9BvJawlcGyY4Ax3F4AzAkCKe+BWZ3UoWzLPL/g7xWsE2mqLZjNtjljzE9YE
MATlHyVVMmJfjXvHAw94c53uvu3zKIASgdlPqNLSY94FzcRst1H8qjeQJOr2QSiq
qhh6Dng+bWEVqdBvVgGeOFYw+CfRuxJB9ZKubBuulCxqwkx+i5941YqnVMU6UTiX
Adh0WfQL/V0XH0BPD9QW1Q8W+u/kQD5yVhkyhEU6L4bMqUWoCHIQYanMFeAsX1vH
2ioc723Xg7VfRoN/IC100rOhNJekeUwoB5j6j7ViTxICJD1P7zAbKkcgKztP1X2E
Hh+2kIJJvuaMbvVZRFLtlDU1POAQ1M1OzJd4k4GCtXavZPm7Dfx/zHQwiGzXZpX7
avW3GUQOxclg40AoGqg4nK1HN4g2xoxA+PC03yj1IdpfwYiChLEen3xcWPP5TlA0
xgSdcXdJLS7wqcBrUiFdiOVc87FqcL+emr9blBJ6SPxXd+G65Oqu+8fLEOmLSO0O
CSv6PBHKS66mwEBk/ZLMsJB97w3ILvOdmNjBkI0F+d/C+SdnDxtxAmEwHGulBjFS
jQrxUJ+88kmpVZpaP4plkexMM2CPVW3HF5kxZh8U2XpUZfQG0HQBZXZ+/i8hbjYD
7gh6d47MTlGA0QXhGQdoPW4MOMUXmRHhBUpPZw6Dhp7XUf7CUPqQovVbHSM7Fjc1
2uUXRldAUU3Lrebx+twyqDAZt06/7ZX8+NHlxEj3YcS0vHTS7DJKpR5J7YLOGqfE
5cIcGbgvMW5UGrpfBbsTaZ1Sje9GT4SUkcSsKfMgkaAOYX2aYLkL0xwUd3BadI7/
27GwDxYUbvDwECNvfJ8GDgeS8HSov7keaXhnEt4s17qZHQeEVTY4gmC5+woZ3+gU
6Z9sIEFw9hCQ2Kcv915VzfBzuz3o/569G6S37bIqs304Xg8Y3m4UO2VXNZZNhsVV
vTiIOXNwcXgzU68Vge4V+E6I9I48GVmWPgfafy2TcG8rTcrnNjsawX9CgPxe0OHQ
S8bVLG1GYyExdltWS/ZA+7RcJ2a/74blEWPIzWiop0nq5feJZCx+jEdKkktTZq9s
7tcf4jqBVt/8RltjW2COULhDmZA5cFyvU09fmdwZixpWBwaHfTXZQb8DbaqCzF65
eY7OLX9FBBzYYIOFUiqjiWX+zEF+dfGcpY3zJNPUWBiXrhNeuDsNQWJfSFQSVPaE
93hdOd3emW+h2tDsg50P3LC5Q/vSErZM6rGuxsIJF8h1FvYUi5JJYebS/cDfNB1y
d2v033WYDVOWnn4pVEksw1Ehq2muNhFUqtLUb+zNJ2O2JXh4gqzek0EjR68ciGwo
AkfedEHqITwcOtTeZZqKf7oCmrcob2Cm0/IwcZDReJsQtQTnDrvAo/inWvadQLTS
Vmn3hbIvsHdja3nicFJ0nqSlgqfxa9sb+1h5yg87zhqQ4ZSQiaH2nRMSw9jwAD3T
DVrHJpbbiSQNBaAevWRiASdvN6Varm4zeluNjHFbV2QDW7iXb2XFhasWnPm2gmR5
CaDZ0ke9DPboAjlIFwR2MkfcgMiNz9OIpySinHMALJfIqCfIAbzQUoEtrUBzd4L/
PsX+WuxkZDYdMToocOS0gxf98eNhBgmZd1x0XDXrnL9pzdjxqxK4RE6zJAbz3ryX
7hid5mQKRNl1NBD4KYrrDunOhQVZEjbJb+5xBBz9ROKBVb+GO4FTJ9BybRbrz3p/
YLQ8sGtmYr6JnHFZep6oPBF86LAOU8T/BiEtflUTimqrlZD6zupsClV5RT0LTYsc
ql1PiDlCDZDYXxw/wIdqbv7qBAzj6IrmEpVidlfG3s1xlsPJ4TVAreDhhfvJN7Z3
RmoTQnLbr2BZOJmoTRgF6LFOJB6pLQChYMIxywRj9EodIo+7HzN9hf9IztSrO6LW
KrwS5XCMkJUn94Z7mvlzFpLJtuhw/Yp2SRJV+HqrJs6VWpEWPsi64MWGIMpV/02l
GFPRXNhtHeHlsNbWK+kqKM+wjTmI1L78Sclv56vDmveX+8o6/ejdjOugxZYa/yCH
KjyeapgiYWSOOuY14hdsMmQ6j2hZo9on8AGqSFMtxiUHbz+B+GfoCT45amp8hJw2
GMH97/yudOAStTY5DqItk70WOxgjp/g8QeN/odGlkZ1Hy1nMTOIPqx7qHWF4+ayZ
VQv7ysbMg+x6NcfszxJnyCGoH6IPiYkga+44AttM9YKXKgkHes+SGQUXNxjjw7RB
oZQMJblOwc/dMds30RyWjH1A+bgTAU8Fr9TB1d60RtXV/BESd4ofErs0WWSQLlEL
WPANeE0jKDbHV3rK8bEZbU7Ix8sKUucM85TUxiDlzzG2/jyqe9dmI4fdpQ8VkvaA
GDiGbyfSE2MbYGhHqNG7uMB1VDh9kiLyu8G0TK96DY3QNIdNYPG5MTziL6H1m3B/
8iA7bcUOU9Ou6KYGO9FEvehpaWYdR+PE0S5jOy9kfMvFcVEUYRHxm2NKEvAGXzQ5
P255A9h2fto3l6A9m1Xk4gjR85hT2eIvKae9kporVZTdBKfhrbLGNjYUPlQDCl8D
Ty9YziEIGGTfXMien+K6CQqh0pJaqI6UR2RN3XprmtVqlJFsua/8TokaqaZ7aS3n
RypfSLdnUqHq/+PxxCt5dktXIDA3rMrS++jxMwL7SBIhzcw4JPcd8hpda9f0bVO1
3LXuZQQvzW5sYjLpqXVnNzwdaIsdG7w9YJYiYWX+SDUQH6+DdiDKkNtwyt+Okd/v
27xBiNNGYZrh/aB+/SivYGmCMBYRyb01NITcdMn1jjXQhopm4RGI88RuGixHfv/z
lZzApsTZO7zob5t4gp2Im6T4g8szSX0tOqM36q2MrHyHknNoMCjsoyWxMHm1jhsK
8ts0afn9pOWcxhfNJE/mmv5zyNC7yqZTKZWcb+4WFyUAts2MbFMCTLhQAw7Q8vY7
Wky9GyrtNE70QziTeeHnrtbaDwXchjfW1NjiDr2ucdLoe5qbj1GHJoAP3FRc10bt
tKqZp4OiCnGve+ZaJrAdskPXxE6wEpNuIuQGJVCmWGL0T25hLH8yhuqf/ZwH30SH
p2VOAa1f517CPG4fuyUlEqBxStKq/txHVtk4iJlynn5+ZpxBwR6tkYL+OsbLIpLK
ZBm17PyQ8rlDeDw7ZOjX3fOwxIcaX5XbrUWmcmaGlFPzjeb+q/cmTEFUgQ9d5a7/
gDtwCNvBclHGVAv8QL/yvCdcOCSGGO1MiIJ15MkDFKhvjgUaYRSORTuToABSbcbM
ETBMyDMlhl0jMJ9Y4v/AWZQrGvMo8M8Y3xEi9OSF2M74y2gwA/Ci0PVZkCjecBRz
mbPv2uhkJahYhcfH/h+BbijcNkStevHMZb0Hpp2T+90TJ3VQWXNDKhyue0Mb4mGs
qCg63Lr/1TepxB28v1UQVViLhmPY0yYfOt5RSeNagwuVpZB1HZqZUotwaQeMjpZR
UXsBZD80o3JBaI343rQPtBJs/2S02rspjMFL9ujvBkc3+O92KEzpLVsrI5hvntEe
Vzu2/XxKsBiSjHVL4FqAbsEH54NhiBwRYQisA5wTd5i1mYhSDUnIx7URqw/EKGFS
tpK0HSHwfFPVVitJAoHNwDu7vlkXzTWZzHnEshQ+fpUCR+uflF4ZTOE2rqzlDZtO
+4ZACr12ZcshVvoqXKVFMmLDYlAolBIi9u/0rELG7AtnKs2HTnOHAyG12mq3gsyn
MG2gtVLnt5BAGBFErtGIUtHVqx1KtbGf+ayVbJRbUFxREW5JQKS4BI0g7pJsP3a8
uz58NgWI6q3MRzLdr2If9MDQM7qrav0LFT+R2y1H2GociqY2dhQPW8uy8BlYf7PH
wC1B9PKcV5SSFkgfWgxAxHecnsW8C78alevqvyc8fRstmaPvMQUrOgrg23kyJy7w
YBeSa/zks+Gr34C2DN5q5wfsV4GSmhwLWUssJ6vQJ6wwYvWXTSq8pK9NhsoC6+z1
aem5IiEzfSJZdztnSizVTBwPanPoGc/69EMMIhqqMnBHZ2GnyoRxNuaJprWBoFc8
BNMXfTWuo2yIRML2g/Ui9MV0btaeDE5gDJCZxJp8YWhgNndy554fwLy7ZwT99cj/
J4PERudGRmIFDoDS0B3XckFsmfn33UlYOUUfOJJBmT/KJboAH0aN1LKotpTYPXY6
Q16GRRdgcK+VTDhbWkU77WTdTp3D4NyllWfhfHU3aKHO7C4FKshW8BNls5eyuziv
fiKHmSomWPwQNWaXLZgVxlK+SmTuNhzGYoNbZjObfKC/tuNtuoEnc1FjV62S7gHt
UnafBuGel0PqiZ5LvQB05Y5FTIQMNXoLb3lo5TX+bIQPgZyqsXGKzMZkjD4idbzR
JhrTrwtAjwGen035js5h2V623tEJLX5+SHA1vM+IjnMm+H2Me4ZvDmm2Z5SUVaBZ
1fkRXk+aRNhsq8PYPXvIJTbAUKvTu64wKURTAon4TcdHb4qBrQEDsywrT5fLqP4g
5UG3DP8VyHARidEYVA7gwap9Ek9ONxKodA73l2hZSp+92V3D2Vo14XI4EPKzlcz5
+9CFcQY3xLXZaYN5GhxYX0GSW49J6MDhouDZkSoKIe2Gp0njceoz6lncEpyyr1Nw
1g5N2CEhbEmy11T6PzBzbeoZ9j4xw0BGCHBxyTM7FbvFI8LM5YmswSNWyLxRFmqs
C0CEm4phfyQ4+sG2yh8XSifoc4WMafm2nYSn9Af+0P0xa2F5m7H40DP83UklG2Hs
G/NSpmBICo1ggCELur4WfSBkQ8LEChZx0fraGZdDZjhsmtVOQ4Z0j/8ahMHusizH
576PTJ0U8BIz1nK3mI1MGdS6g+3qtvUP1VWyq36h3ggF8MXvr7wnE82rRbIQTEzM
4JGLjv46sIZKrKbQ1M+PpKY8VMFzIdTPv3E/3NNKZZpz+WbjEp/6ZVsRJ0FY7pwO
jvbffN0OOLiFBHgkxNGt0t0aRB6ITT/N/C+/Jtv4WrVMU39KSpXyPZxEK6OlLpsO
WfKy2ugIzzun+qQ8yEeEh0mhixt+QYEI6lwvOOoWzelGvqWjvVMGZ44/O08L2CAy
eziBswnOMyrLKIJjsKtpkBvX5PbwWDnBSOYD5zAORbQBehjoIVtgDzSoif5HbRl/
AifsWqDQGn7EJGDsr9GB7do3LZ02fwkBXRjo6VOwjkcFA+T57a5skWfM9HGAIgkn
wNNz1lecSOy0oXIM7bLhoYz7XBC3n92FXs8k3Sdefj76pq34sysmiQb6gNuSjkfN
Eb2jMboM6kOYq9pJvVPecJ15BYxR+T8BVBqH9NmiGkOJkngKdL94+NxhQgge69yT
g+rDxlVRxkMvFLvsgRWs9cefGQcPRedIazRLru09jBU3Eb2HN3GF+98PzizWePfN
fa/uyEIzv1PqU4m5sB+mA60UDSTqvmWkkWiEKBOHAmesUXIkLuy8t7ZFK0o6u9cs
J5Vzs0e6lXPnDrC0K5Rn89Z0NalW5F2QYwrdkWoZT7Tjsob9ACrof0GXBYdIrsif
IgeudxM1vNoF23XEWVkwkbqUpRLDzt5r8brHXDXKu6in8FnMK/MVu63D7nLHxQEV
RFQjgNf3lvfj3LHO4yLU/q2oPaOvtmfaV2Hj1xC0bhvYUwIbMixHnlfM2FnHzzNS
3zareQnEMukYsep6XVmkS3y/xXnzK3V0GjRR1LtPGIuVkVf5+tI+lIV2I+b/IKiH
V+J9iJCT8HV/CzG885zZ1uIbCjdt76k3RzARCglRwEIBGVQERFX2CROv+fYstkqU
Dg84jPq3bxJVQI8IhSppHOytUZW6IRUuXURG4TYB0fWIB6AurJF5U7+h/xuiV7XC
RVvOK2cj+AMss6VmY+IWmFo+YiugnWE8nQBvQZTep44X7WK9iQlkWWiQ667IzZl2
QxR2hrnHPKcPAzp7qOKHYXVb5Yly0K+5Qj8gCHMrTu1B8noaPoZ3BwBid0KPaagx
CT/hQEGyw6gkzUQTCm3EPCT4aJWhpwfR9HE+DQoorhu8S0bmSrBEdHBzimi2sgXX
SWhvMzsp6+FLjMz5FdN3YcOZGIgzvyo2gB+DzgSvCKDITN+hzEf4GqrGK1JthjAG
K/ULN4JFxeGH776oOG0biPy1yAzNHrj4OmKVJIAVUSSEOyaU4OaAF95eNDOOIEhd
5V+UQxjmeNRcBLHc6j8f9P7rtyCExr/NVR7R5Dj4DFTMeNMyokcBglxIF0O/oALX
eNZ7yufoGGTN0A+ehnmrRAlpN+nHgpxKxva8nl0eoBxZ9huZglyWQuW5o9KJMVyN
lBM1J0VcapmavbI5iVnkAIh3blgueKh/vVcS5GftLyAKadzoLgLQyjbOgz5VM2ui
GH9bl4avCUaWCE6j2pGdqc8XN5bzczmsJY8c738i1DGFCJfHdpo9E2/ZAT5q0kXM
m5FEMcjL2vUQCy1dkm64Xw215nvu6icccXCrWL7dwVqOzq2qRDdeynyO4Bux6cyk
S5gODS0lZVXK+Bjf14wdK6Fitx6GY2UkT6Xaw20iUdFh7ohjK9DD3YU7CfaFqevF
G6oN5ea9O63tqdJsZNF3JEkpZiM5m27lq9km4uBj9ubU0YhehG1b7WSm1ebJvaIw
cp6PSatV+M5AzzlwT902g3IoguvMZadWwjQFLj1COije7VhUHeXM07QpGvs1KEA8
xfjn9NEOBLftoTozLGktyfDCr/suhsbwd9Wde66k326Rci3ZTFlRu9j7TEwSIAim
jgaYP7IBMS7/ZdV6nZNR1boFDVOeRPpVA+aGh7QbLAfpKv6xcrWVM1EASJoZNnJm
F7E8UlhuwIe5qi5xW0uKfwqr6yYqCVuLrL0ZNs2SxPN1fQ4CAg+M374vTDCPkCeu
uKgRw8WTuLXtp4VBKYZzOc+ujHYsLOoKMEy9hoL79qaW4RgN/e1BqS1y59q9eGgW
XqeDBKmY/0IJKPxdpQ+5Vmri84LasxRTHCaaYC4tmSVVpQ0GYKgU/m0Ewx+BoVCH
5ZzhmnMfgnNoJj/JhOSdeO0SeB5rQK+9KHLn4QwYzMYROMXYnTb1HR8ikex5vp/L
8UpQ2FJ5yyEAm7kHhTR/qAA1bLIFZSduFlH39Xm7J2XHxiunMpRnyC6/KqbetOKo
v+BiBlC6H5Oba469plSgEPveQjKLBEacEyRuMgFeVR5U4mC8n3RUPNhxjZCP++Ew
F3Bw/P1D0cDH3vHLYGg0MGUPuwADDf2F4bf6+efJVZvxXYZV9x6jK4dIrlvKrqSZ
8hnloKdrtyYHllm1cP1hwODONA7/eXYvUvh6ZAIfAy25RPV5E/ycIRuF/GqnvScU
8tiSBq4/Ievo8on3hcwOOtw0ih0gCQVxY0s89B0E68fhhI9oDrX/lFIbRHkvc8OA
2R9oljpNxrPApEdpkoqifmFdFH3hEBx7fjaUvCfvw/Chpf82SEr7g+f5BJogQayn
MdFOwAN2n3qE0Jhj2MWWchm+kAOY2jN6Ne05HJJMKgUv0kPR6QgL8c5FCU1miHEE
iimngabWNtJKDjDnE82c5LEE3xGNnUzkz4zZ0igCsJe4VWLyx/NxD0MAecQPxZ92
G306ja8nBKu+Je4pECRitqxzE4k05mR43QsSmGShoQGRIou9mQM+SY43ZvkxSoci
frXmvf6r28CMwjSrxXBUaRJAcFrGy9hZ7iXMI6AqfdZ+Adsn0X+i+P8H1WJYuWIq
6oamOrtcFx5UKb84KBiZXjKSdyj57k+nZ250sugK5xj1TedAffWsphlG2GcAnAIx
9uI2GM4fP+JtQeVHRX4wAlLnvQaSHuCb4XamJ33VdULU/LVyJ0vphhesqAV6wOma
I5XxIlr3p9FvVBW1Ivx9HPPan5NpKYe2qUFVhtqgOtKpPlkUm9nzyazHmzSAS721
Ojv06VKC84JhzGZuDC+LGqjB6+79CuuaqlBh2Q8/O9IJ5W6oeB1pHTKeaYxHJcay
/TUn62h4a6KXd0x/ksmqvkMbfWfdP31cHvVM/yQFyKFbAEIzqOrpExvNT7VISZJ8
r2iqNhYFZ6pMS5YUTsApGuXCKKFZzdZbjNEZxM0z028JVtYUW79bRCL7CApogh8n
u3tRLTnSVh3IY1BYr6tchAbkiMqm3Qg4ixS9DSmlnpdqWro3M2/sZhHw6ltxdnnL
RSdygm/Fp6qIBoSy8cOqB4Juxhr61rbQrc/nN2lJx2YIa15Vbi+DriKU//hqAsp3
c0VaOLy6NuGgHco+uzrqqkq1ZVyZ8oJnjN3jws6noxGG0VyBzclHOXy18FHOl/Mi
5cydK3qfhAHhqxia1tBb0roSPIqLSRyKW5AFH4Mis02/Md5ViOR1crS9lQLVr1Kk
q/NUS1ScEXDgDVHwE+8hMY9z+dnMotJO1kJHjfmnW+p0Pti6OwOIS5Cg+8E+rDv7
0iWjbRE3SzOO06obIiPGKEVLlw9nSWBWuptau9nitOuH8J0DVVLpnp0/L7O46uDp
yvIAihG4428MGaRnbBqEF72T/HVMcUw0OJdp+BtUyZpj6BAywhVNaFT6cpvXZcEk
9D3iJoGz1eSqVE7O8DRwnextoY9PzR3OjYM2ygAgJDEMnjeV9+4625AR3XEFMXrw
KOBvbz2lmMx9PHzi+iTB7XtYjzMvtUb0ZadkIORtjFYUJLkHxwGXET96bYeMB7Lt
VtPZWdRvdM/jaHpRcQTqAISyVY3xFey3W87RvB2Mc+UfWSF7POqUbrmuMITu3BiB
I2I0ZNZuIfZdlfQlMlGzIvi+UB/iLu6DgNFxk5g875AXoFyd+wFz4aW3HsOjKrDf
vssmtlOn6toQXa7to9Bf0Y+9NFVecKLx6YKMH/XaFdBnyAKV3W7UFbpc3ddNXhj0
bPqgtIeR8TVSqYW955+10ra/Tgplk7/Naf0Wg63UT65h+N2AC/hk2YHiFUQQi/mC
vHNYlKlGsES0u2ygAlXPZ/BBq9tXtCOuZ7WhRzFN2vSbs55lNRdD1MJvuU44kTGr
zwFbqQfILDITcR50Ghe+33BAiF46pBl1NUGuwR6VTbgKOnZnDAumXLjXHJrcfzh1
Nf0n2WZyKBTmXKSIy3nqZ7a4ycE5UMVRv4xlagNb01xl/Dim3zL8E/vGoX51M0Uo
GPP5y9tQfnzfhpM8AB6mngNmmxhrGnMXy6XRZa231IA8f69jY5TAILeQjKSOMhLh
Q725umo0jMf+DDOaOptF1WQt1334R7jw4W4CFZ0yLEM3owNN7KgYQs2loDdS+tdJ
dF84bs+t4ANK+mooP/zHc36K21Aalfpz44Nyzse9liKx+0rBeOjV7xMboXfQvdpb
0RAsrPjYa041LqWcWPPY1e3phT8F45O1Bu1Rxow6FCpstUKqrgbusUT84uY4tzuW
MVthNq8bmi2DN/ZtEJYQ4OjUAo3+nGWFFuXQY514aK6Y/52hU6k59eClwruONwZ0
+FeljC6TUuQlaF8zQ3uK808YkVo6LNa/lZXgl6mcjcQbwU4OwJ20xzEo1pmYsyoG
bt9bLT/dTKDm9xhGNRb5NX45/HxMQO+hkY0ntnsrewN8kaAAExWzHq0vne75tlrQ
QPNkNPvnKHSu4IGBrVB8uObRzz+OppBSZwBKRkRnb6p+A5TRSj1cwQtZPUt2x3St
OP1+1wZxt4hS/smLdxKLhdHdXI4mZuannA3Wo+DvV0OmKpqGWqbcWzzENNun5f9f
DRIQDwVWZy971/UMBt1Whljh9HRmuu3SE4maCKPv2eMHZoFHPFIt74fwXzpcuRE/
nif88OBGdHYyzOe3otiwtoglX7mQcWQLfOUbe7y+8pyxhAoFDRZraSwT6w0A4jnK
/Nr18QrP7eepgKHVAjQL3U0CsU+P9da3K07gVgimuLk6KhVpice7tSuXWmPqoNi4
blEkW+8Vnj5NEhUYzlwoPJvQEy7geZmZQe8rnlvXarv8p916K2E7T1Q/a7B1SCB1
3TOwGeFAwkqZ8i5fwURsxqIyrb63OpfKzHSjtqvDgqa+Fe4xOJuaixRJ1owbtT3O
2LowpzZ0kIST8vNOvR8aGP6EYV8daWhbBiWo4i1XfOar+k2zTtmqwqR44Q0NxkCS
mj6Yi5gXvaHxXgW2cen4RhrcaR8O/bHKwx/V2wuxgQ7cbmZBYk5VSHGE+wi5zjF4
pVFunO+s6JcqVrhzGErwYLdrWMwLpiZ1W26TvQmJKDaidTo+5v7NgfUFLAmkG2YC
dno2Op8rqScwunODZe4Fi5cHgQtmZXQFCqOs4h4bm4iAlanl8MlbVQq8DZjAkKUb
jle6aXZb/VHVeQPNKd/6EXDPPB4WCm1KhDjr51l20Pw5STkTNaMasFtnz8fm4z3R
Z7/MdN+oxIEDq2toW4zaldTVpL3oYy21Tp8Smzj1kOkHf1RYozjkRastp91dU0LP
IO3ONQC1lGP0Qs2i/LFwiY4KqP8PGBwj5hV+u1u+EfjM5lKiAfW0jwcH0IXrC7NT
KZ/ceVhCOqK2CaYRRF2RKzNYDr6oBoxGE0QMt7q6uatjpZg2N7FU4FVqpZagCU5U
q0B8wL/IefgfYpKQie5Z12R5WHSELH9T30JPEkEjefS74WiBhjQrhfqdX3uSAjVP
cAKv86omHlkgaRN0Jfgqllnhcmz8mVLW6gqBGs+JVkO7r0AMvFyyPcoVWNZxlQmG
sR3GGHIUJKphNS59CPTqqOOQWAh+k5Kgs9rBMUUH376PFI13kOvSUsEqbEBRl4Zx
i7bmkWXYOYWpzN2dAKuVx6bWVJ0BXkFSuoxJg22r8N9N3l/Sqfslly4LepiooCb1
8AoQCR8f4rngTbcNyanFZTyyRhxa8t2huk9XaGVyWCZGmOHrqnz1CiQEwvfwj9sO
s73ttqk1qka6AInlUoJm3+IPFbXcBru9UXl3brqRDLsjEHDpVmlYSUSg5XRPs9SA
6O8I0LpmX3K5QDujRG9bqvTtiVKHgX5/+ygLfhjfbl3hN5QsEgWVvy4jqEExoxin
q84DWE8wsxyl+l6jUokYLjK/+N46Rx7pQdK8/oLpUHsFrB9HfkSTsZUREv6kpuw9
sGVEOBO17Rh8ZUfo1CACLdcYzGz/ER1EulKGnE3YXFIfa2xQScQVGbe98ckcXGOz
Ic5wRoK6WSxGogN0CJXrv6upS7hnFbM7BSHGfXFdSKldes4PSqAwCqLqVM5GpHVj
4uycCVBxfZabiyUFbjAutq2UXqhH0TlAziXUyVP5WkmSqHkebEqycW5UMvWfFjeo
UPbz2mcyTwIelDwwAUcfI4lqP1hkrwBNlRxU9htCwAsPx58F9M8eYXqgG2Wydg4k
UTvLX5r8pj/jbi24zi1ybH0DBGK62ik5iAPF71yg8YbbPpIuijXWj1Je1k6JeOgN
k1zXxqIU6qBxkmvUs8IyILDJcb6qlnpDjxQTPrj07VIdFCaI8O6nPuxlvXykuaJ6
+q0fxKsETnwVNzmbiPjC61T67JCDWk3j80G6EjP/PzpH1F1M5OUclsvKIZCb8mND
SBdS9Aa9RQ8D/s+W/7KxJ9dWHD4RJQ21IMvpjSoRi0b9ej+XooQxgzs/gDu1KAts
ub1bD7jNSCbpB721GXO8F230kP+eeFlf5QCX1z9UvkhyKfpDKp2AIUKRZLnLK8Bg
pCvy14ezppKKuT5zrBz52dqjzLZ8th+oKAny0pLJfJRqTwEICKXsxxQQ2GrefVSf
EcexUaIFSmVRQXinDB4GwO+RyWxv+2s1mJzsb/8Rs2rOfcFPVv/O+4TcBBnlt41Q
cHMw5mB/do5F21pAOunav5GwPG+VdKmAGsOfeAS4/IY4FpWeBTp2GxBWDJ+6jPVk
QqkEikGmsyCJv471qAxmUYJZ0luvN5gVjEh8z/Rb3HS8ZDu3814hxk7M468WusPV
HQaewU7f7MHFGg5X3Oo+xf5ZOeL19oFs3t+EJMoyaa4/U1ieaoZFCX1DE7eYgic4
XFdXyDagMqhOdaiGYsLItJkfV9/TpJhTD1GRvz4pmTibk+W8ewaLo6BEeqIqj8rG
i8NMyMNvXS8LXBTwQvvGwobGa1eDTnxxnLcdD5UkxkvMrO+FhdU6z1n8yXbFFMB2
3VAEsCqOYITfdQx2lBVSyhRZntD2bgWHMcX66GfQTAfFCPMmnLSza+eg+1vlITDH
SRmBFnLw9U5BixcObk3LeYrSWecVaGapvCj/nOsFvlfU8KMM+PYuem29Orkcct1q
XjQlVAunwFhdHbGU0ghn7z+qX1nIcNIl9jCAYqyFW+tq6blhjGenwIv7dsnAUH1o
8/HvqFR+SXq8TGhRQ0NVCIMGrXJGMVGCM780OrVIgIQmn4VI0zwHFnIhvZnihF24
x0CaMmgAEqwZoOQ0s1uuN3FP8wZY0caKuiDZlcTkqNZCicOJG018G9r4TTyL/cuW
B+stOySd97T10cuVzymr0PRwl2wqX9KJkvAzKlXSE+AcjFHcGp/C1CD3i3jnOY72
4yS8gUXpBGZlLmGdSWKE6YRzJijU14pdo9RvgQPyR2MoZOE8mmZasPotWaaopqDv
q517tTs8fq/15Y960qa8v6WfhSzsES2kSn7223/qxVMK8XKeZ954qVVwRE3/YkGF
N8PrV/JVuKJdjT0Bw+ZwHAI8gcqftpFcC+iQtESjO7ixSJJxPOa7WKN2dKTFwm1b
wqs33uwPUbi6GZk8xbvGAIp6xaJov/e6rPnPKV0hba5qQcMNVdUm+vjTc1aVAooW
/osWOW3bqXuWfdq/5xXq5jneZtHp0PUhv0ZSDTWqe06gEMhsVl5c4LCHk04E3pBT
P65DzDE9iBNNBbzbOw2DVMrdZWJQt+r/9OPZerZD6AlHYq6onRtS04pgsj2Zd/Fr
FVUkyi51fL7tkILtL9E22rgO8ZHSBIAcVfzLW1mURdWvYEk8TqPfRWNKKJcvlZ+F
Iyd/amMbnxqniN0KfUceZL3yCHuoPZcSswga+ox+J/EfW3sWWGphrMuOyrVe7kPb
QfH6sI2UqVZO0e+nJSPjy1ajjtwaeYfC+sF4+AN76hFbuGsbp6sfG/WtvIxV7WR4
u7ZLVSZo29T/bM+OMxCEG4x3pExKVOLNFbBrdbzrfzOboewqQzLC2WNHTVHUTiK5
0SxiOiD+Kcau7Oy5ieWU87jeytvveO04wh+E5DLwKPdUtMt0ZBJ7gqhMyEEXl2GH
9KObvwvupMd4E7kXqPwoMqTy2OVBlZL9ad5dN2YNe5SepYXcnokZmEPmDGF2vsPw
jHB6pXtuB0KugpIz/BTTCN0b2uk02bqMfegwKuOUvhhuqzdCAnrS1FomTi+EKpI5
ljsH/mkkidmXBy6uDEuZBDlrrCkXvnuZGkV2IDH4hG5vSvpRVqgDlsuAVGRR3zk9
umFCaGtoRa+eNCOYRmUoIc0RwTOwMe5JhcXtFlH0cFKh4QPUGTD0Qdzt+pLxuUR+
coNJCq6YrlIghBkS6hVNmJo61uc12ZOqlgGss71913jCApo6HqeG7l//aGB4zRqx
x1eZomksLjP2D0X40oORBA7XvK8SEwY0N8gdbUQT1E/+ejIFc+gTk+I+Az8jPAfx
YEo6yLF/kMXQDXtsmWiylHniJaNrAnKRg2ZJ2/lvAPekh7yCuWgAz1bQknSBHk39
tReVynJ18FnjrB1zT9JVp5hzqXjJ2CUgZywfTPBNgAZ2KU/c2YXGx6vUDv3X01na
sEcX70nztpHnC2Rq9coOAi3PACd/MXp4P+JZtF7Z7yNzdBShVgW//t/50HJGOjmR
/YLMGSUQN/BICnieSiIVlfBEN2z/WLJ9tjx8wHkmrzC2aHx1iUCWje23gEhL/dJq
2uUXLX0NGplhmjB8Q2ojlopg5G7NVaHyKAlZxyxcXFy0AYQ+AlIClBLMKVbUlMjE
+sqwu5sO40Y+rj89PTAPCgGoJcuz1clHZC5/cev/sYnE0AcPoxmmnJs9aLTcYjBg
t+PvJPGkE9XsFskNXEqEYtNzJOvE976XnI5KUUgxe6spxoaukMpDto9l5U42hYbU
4/VXiBd3Ut+v/gaJXxq1ggq+fmYSCE2eHBV6bH8dsXoRXNjl1jQw+mqIj5fXAKO8
G+dwCGjHACfr7mWQuFUjB3TQERv56eDdAsl5mio0XItnSphlgy4/ZxMXNiZwmiBM
o7LAS5ieGAVe4ktPLwMte265A/NIwD7iTbY6TkcpDsPWeqDGDEYWqM4aSRC1/UFX
t8EsWFeyN01UrPX51/RwLrFIfqXsAaHi63VaJZQakw8bdOBJWjzHEyDgXZhBFQmR
TVMzMca9i97pFRTT1XfzWLUu1okgiLk0pxbSdwfQmU+noiBdK1kw5uuns1nFP17A
wX05j3/kNMce3k/8k7622vaNNtXpwtJODQET9pYYF2t27IUWaU80qtwmt1blulKi
rlSoeEUtlVPS9pubaXpX/VMwcX/hKLQ+uOCu9+uBEEytNL6+uiWXXPz70P3BGSLG
8qM/gXgQMc7haNNwL8XvZoYpq0YCU1AQ0d7tC29QoyIxUiK0sxcL3AyuSS/w6LZQ
AM9NplptQIWCwpy2o05IKT55XBsqA5Ggj0hyGuqVSwYAW45wTmsYho7uc+xtMTfi
lAFKB+beH6CjnotAgf7rg41On3QWCz6KqszYyEnIYRDrn69+2v8xyAhTpz65Z03u
xPXjgnMSLjQgLQ0rdQDFCIW5JwoOB3mQyg3W107YU+u+HTG5BuZMHZofpamQ+/6K
3Jb4X0XgtV5ItN0Iud3OLjAVgphXV7ujncmgORGFQKGtkIFpv2iW+f8tHVXuVgMr
IERAmrX9EmMBP/iHYR09QDSS+5tkjw2+nt1XJof/FmyuOK/WALgjzBzuzN0SFRy3
VgRfM63b7PF8LOzBZKh0xNFWaT9l0+Cy2Vdw8TxCuJHArSiwyUyZVAkqyRa1qVd2
bsHa2q71u/vuKiecACQolxRzbqJnK1jBkIAQHmER7u8f+fYPY21dkDWzphqG/wly
btVE9tjKHdae2C3D4GGIqqZvj7pOb+HMirKUdCo5sh6KynlRApkXRaOR7btNrsJu
ugnICiC9en1e/py8WBNG9EHStsERJtgKQJTZHBXrprV/nsjj/tYq118BaKV1P4gm
AUvFNluHHvTieCI4XvUz4P2wu62VfobcPZTD4y6ozgMDSyApY9V8xKL0eU+ogqm6
aL5Jq1qABRil0mCcZmXHUB1RLUSGiiK02bSNomixzDji85upoeSUBUwaxze72i0e
qgrLk1xAjkoMmCbop+2tpto6fZmHe7HRDwuvzPI2245IJmL/Dhsgj4a3WijxKXEt
6P68pNph9bO8xAc+R6wglWk2fECrkAPvokLWNhc1uJGm1/ufLmWhsUSUtIWHl4lJ
xmH6S6oMrbVDOH3vWTJIj/kNx4MOJrFYlkaNUp+j7JV9K4ODhASJkzOSHhPtELph
NOf/qbesokubKH18WAZ0ckP0thIUbDnAGkMU4dAPLisvVxvo7AyN2svDVoMxHjwV
v30zUOzixcdI/wSslqhF4p456vvXTS7cH5q0XpqPvwj0Xk/EyukA/W6gg6YdqnSP
AJN75iwbEMJTs1DdA3iUs/zNYh4BNkYoLNnX4vI3pEXNUTRXEk6C2DqfI/DOYQw1
0TBJo0ZXUxZ1/pNvDTdHHQqHUfv69TPqSIk6M2gKjy2aOk8LQ0W+4zJt6NBlnozA
J1v85TmDPopbOO3t1rCl+MpMmukCeQtzaQ0Rdizp+ZQ8eJ04DUSY7fXCwkYJ/HOj
9ekKL6ZZKVESx4elVKYhLqJtU/oxr1tKOCJ5HArOv2ePsqpF75BkfD2kUlDMNkIY
bq1vdKS3O9arP0ISZ5FQy8JQbaSi7rrx660kO+oMuxdoCP1B9BPcpq2ad2HFsOVZ
HnchS2qzEI0vpehkEWgKDJu0qjtzslN39BNcyWjnze1U29T03arOhjrE2ai5+oD3
7tCa43XKwHiwpjk5uPmlInwgRNgGQgwYAaUGcBPbxAiqhpvs1xMly0c21zAi7oO2
b/TSsE7rvBajgQ7M8WFl0tk3sylcstR7OtdHVzQNXf3qMmRt6o0yYyU0B4ic+2g2
TnxwqQMZl7zTCOvbmUM851OuYvkiEOyzbCWU+iILRmlbnen7J6i5D5JVIl/vM9i3
FsunAX8M9bkLLLse6EbhtRcVFVsoxWUKLTjbesTKz5Hfb/681Hwh6AcGLDJyVBLh
vESA3dAXCTYZJjUVQ/Q6N+8NqT4dH2tr1ivlMn1Qir9dgJexa6iSHRUaAsBTr3sF
4xSX/2opAYpi7IUGY9jNxNsG/PVYC7ViUcqrGpV4vl6CgHomCQ4Fk5YHFjw94mBO
WXEn+KdCjzNX5t0NPaw+58ct/awfZ+bBDcKEj3wVGe0TUmjK7iwxk3W+37OUvykr
9RRf5a+9t+sMseQrlIyDvkDca30sQB6Oyuf5gzsuvViufqElxLCbQhDDKpAFlSOH
tgs2olasC80jyvzcAZfeqF8E2CcdEfwWAWqzves05rdh7TwGX4sc8dY+VnX63X40
vKeBUjHO/KQA/0foaw6IpBsK5BBVzpvRl16bhJP6ulNUmeiHqQjT6ZR3SE8me9/2
KSFd2EH2TBzynvC8GY1jj9Q+8zixzrHOb8vVf9DNrPgo8acOByC8Agnyz6IK2tOG
D66M4Z7l8IQdaSrJHJf8owLMDZcZ2+BBAEheO+1DRDcupaZCXyUsJD3vkQyufbBv
sw4UvU1Bh+TeG1/ynsDZMxSRn3RE2CxI7R0+nyDjDK7dNerBXRaHmJY+/Qd8PjlV
6OfWN1ZjzI5J/w3n9CHXJejt7lYNQEAsDeKKw4kbIMN0cEsDUsbnE9cysc3GJjGh
qVNVDQAwCsN2/YTOQ5taz1fbGGo1pjibqrSe44nV07GLNbnzp+hz7LQ8IQhdYk9H
RZrDTqFcUEX4ALPGgF4PhobJIdX+kfHGZy1jfXSrQNFek6xp0Rsmsi8wrbdYtC6W
gsarNv5mjWc8DDP9LpZ+BabwsyzXaPQYlobOfxjOlklnxS04lbqgkdtOH6sxapOu
Bp21AvYpaqgq5rTHXxr9v73iuRULqvZqGzInMDu/hiqZlz9Im9Qkq+Wy2K+MgFUF
7zjVsmewT+x+ZwsNTTLzjsCsK3FPzwVq67wF6cQICi/vqC0nR/pnfJ697LfoiO57
VwGDXMhfXoQRGjx+KDY19efyT8vbf/beuuftQofaa3aIkJyQELC9puYGn8ylzEvH
NA9+yv+kXC9WZokfd1/jMLaRDYKpvzRzBv21R0D+4MKVHDTUjWKl48Gz3j3PfYD5
iIRv9Qhy/JR4kwcxMh/7MhLR7oON/8NcLKkhr4cgqktPBej9lKsfhP9W4OxLdFWz
91SbnX+zumH6q2gewlWmb7kZD+fbFytZsh9qYKvJUkGyeQhu6X9CFbBGKTLHKZh+
FrzKfEJvkyhptzxF90Lpr3prFVVqJ6iAkogT2w0iY8DXm8L5ViQKrkBpc99iEakV
FZaso6vvKFClc8YL5JXx6CjrzaCiG7ThqoFTAI6jOtJqcfZTXpw+NCdSBv2UfNjA
8rMWYA47geTdfQZ6nj/LlF5mEDXuOQH8WIkwg0vPLV/fCaamXRwxAedCTVBftQMB
Fo8M7BmnyfQGCIOpwQiPyFKuoqYScs246DxlhaILROKqSryvJIG97J1Op+ztLiKe
Y3FuCuVTUaNpNV/+uHszu32afrz7Y/vnexF80iSL5Yq6AL3dFUaMYpJB1XLkjuLu
9sh16FJpQN+hizfhwS34FzxfiPFW8zZIu4o6C5yJOrc+g5PKiIJv6p7zIAYRbWca
krK2aa4toKRHaJlppnur2wlZfVfckGJOPJLuNIDOXlraIu3mVkxkHrsoRYP8eUQk
uBlWxxCOeG4s7EMiL0qm9FgneOQOwfYRf+Vr6rKzufpQSH7mO5Q/mloxUCOQnI8B
hDEqTjxP4o4/9GOWTVcsa3p7XaYsibJukKrpYJcc09hr9EqDocgStwXAQku9JTT7
R8cwvVgq5Z0mncwqKrNfgs9ccMqdysWxVIKwSjR1AHxByias+NnCEBQKfZDX6Kup
AL6qtMr5mkxxhUGiOiAfy2zbuJ0Zm6KSdj5CI539UHx2J4z51YQd5Cct7a3vivJN
0mH4kxox2aSU02qvkRKB7nAINo3J5o78mkGXSFVEtOg4oUkWSK8Z3kkBktGqLCIf
2Tb1MhybGtdszwhbFU2+riNpab+vHj75FoQ1TUQqiJQLZuc819ALRHp+W4GgRLJQ
9nLMLNwZtUSBquJNth2EiKCLgtCJql1dtnTB6Qqx9pKToi4ZfmpQS67vfNqjw7NE
praI9NZ3w6C/fj3mbg7rWosiZwNnPB03SE9knmBeHne95I2ul3XS8l8P8VleHhl0
V7NFNN5JonEFEdURKKKtR54HTx6sP+P4gen2aXy2/6NXJsO14wCyjrxrMZjglNqv
UFS7ENGamECEa1DVHw2AuEO/sLQGOywMLQ3q3HoDxhZOpPdO6bOTPAhgQ8Q+56bs
FblMwe9w6s9x3GE9Ah/89west5A87rTF4rwa+DgIEXNeFeUHrPw43VVPab3wClN4
NzJmJgY6Cy3Bsfj9EfU2oYCtk0jg0xZovrvVyr8VuovAfclniM8Tmm2ClHRpakqY
Z+pnK3uvI7Q8ljzpBhiV+sb4+nxcNJ43C34bigjizba4PLUr6UMtxJvQ6PBa4ejL
MV6JGn/e1m/ScrXlmHqXUZhevVrmnXy5lWRQUOMO8OpFNdQfPvpEHBW9jSF86erM
2rKiazTe1jUhhHlSzHufOb4b2b/75LGt9cd6vK85Tvh4T2kMRBMUOG4z1E6QApUa
zmLX/tfdDnFhPBQcXx3xWTtCnFrU2GSp2MYWUfQAbA4zELVhWa4UNDljl1AyCetL
48D6fJZ5UeaHsE4B1cFxkvR/0+awNjxRPDkqepFzIvX0fs2QxvG4YoerTskX0Zeb
iHCRxriyu6+ICIj2SC4k0cHa/3bhm1FsNi8BxtDzPR+sAMYbyvj+h3FKxVwsKjIR
JIfLtszvdJPTkVJEGKf6c6rs2xcKgidG9mcVCn60V9SUG5CS1t021lMEYrw7qIst
s7/ALOSjJqi4QYqRA5JZeaM6T6NQH2jr18B8aHqVWVjpLe3EocwjcpJUuxb6uxZ9
nKhnCQKrYioa5QmyhM8NPO9pfFih9UoTaCstTUZuOZA1WUSA4Aua+TmEOhYXiMdq
Oj+A6I8CIENzCbV/+WxiYSXiIIuuTzSaaCUv6rQkz13Mo8ubQJvDDHM1XXolkV3r
oNwOGU1yOdP+CPYpiW8JId1KmlSv660Ri8cBAXRVGyzOk2jbhTmLSXmDhbnT+nt3
4CVhs9oSgFtkw5plzL5il1GCzqmFz2hUnWb4Qk5OikIm5U9n1UleWKi5w7rq0zTe
ts0zxqX6xqlfo2yjsFBdUZ3IJ5/Q7hrSZAi5jGRUT6s4lhP2q5NvPHO4sL1srfJp
3jFb+okZIrftVjX3AL2wp3dkz4eOuhcra6gdAffreK8lfp7JQakOrlhlVxASBTtZ
T4ZwLYMm9nlIho+jxBnFVcbDpxSkqxG7hdmxOhviLgDZ5cQ9E0nc0NcTFk4lxq5V
QMCS1oC67cNAXjQ3HM9z3VGGZPbdc+QdCg9LmuyZff45m9z9iZphyKpV5WcIC+ne
7PGROvxcshwxNSCVTouxsjMOlaqOFY9Pzib/Wqu58wTdIIb+B2aVGd7zCqTpYx29
n3cap/+TJ55ApvoygsYOJMrvI/WToyzoIIbekrPYllaomwHnPgbId3+nAoZM5SmP
bgfo0Gt6MWEQtYITr1SlpWFLJd0aczo/Z4M/sm1K1FjD6e5foTxFO1AJrMWpPnsA
krlhBKP8kNlQyqZQaxaCkyVkb/PazR+dCfIWnZ2rE1UEBP/FewKCAp+zkxan9Ns7
JhNbhQE3bEinAfkEiEDPO+SJVhi5FWXop38QkGMJbDjFoZDIeVJHfFkpQoWuNLql
Rb4Luec7O9b8ajNg/yGotInOL0gEl871iwesmEN7TGg2WN/nDVZYJ40HlygKWZmm
td8+h+F1q9aV/86Hhg9YeFUBvRFL+mDcRK4dwwLwTZ+Mzz6Z2JkBMVY/116Lm94b
OGtiM65mBL7ZwzxFN2ZsrZP6ISv/bqaBohrdI2SfOh7bEsNAKrbnLXrJPjIzTe54
2uLVdyN8GN+4JFxCctcyMbph8xWtSPsBFgvFCSgVjaQxSl400r3BiNtcR4DgsNim
CK3VYyF/Bfuz7eB3HEc1ddQp20W72hfPjvHJdNwVZTTafttHj/MGIhGGyBsgy8Cd
o7xkPlt9M4VFkeaG9sZa7gXVXyUDkaZXXAf2GooWte1xsAqdvI+m7zbvD4qU6Dee
U/HNgYJWKSPifqQMqd9pylSGOIeAv7JoSC2FCptN36YHLbwQzxGr2jgXsa10I5UR
U9lRU9BW5sk6fIfnbAAECqLnMQMlad2xGVmVQKwSOpXVVf25Y/7xQ2xRuggUQZgo
QImRJsC1jvFx7rXBdS/pxG26wXU1fdiHyKKTyREPFmTQKXDf9u3VzJiSE3JikYxq
e7ZzihQ0bVzkBLvQFNVrADnroZHbMCSs9XjuMYzLOaekZ60uZeH2QyX79fcvTrbj
JLZ5cvbYUBmR473XXnvl4AgSAHVzzt4xppexPQV6nZt/GrxW3BygZLH2MPUs5orI
BJoeYipejNgLW55djCrjM8DP/+Y9Vo50+L95vWW6XNGnBy85tkqXH6geQfsuuR2b
zBrljVrhn1d6sX4sUmOpPlUecpCabLTKohpz07AVhmGPxQ9LHA94VcgpMIp3PZFF
SgX/pBXjRGBE0wcs2X9tqGmqHxjRJeTU8g5lGVk4nbipD+LO75dKvp4654tv0Nni
D5XurQRL6f8S5Ewg45fq2UEiFH1L1BQ0uY5wmNCZ4C7fc/iI4PkS+VvtwgCnG6qW
Nu3nXY5MlMApZa6VSKcNJBMQUgEL28yODPlfsZFLfpQ19I1YaB2aJvqISGAHgc/+
0bZCWPI7hxVpnZa3ru/q62Lv4XOfymjQMST1wydbeuDvFa48xnSmCgKJCnNVn3Ce
h69qezwqeHgdDPJzyv1Dfwujuz/leZY+hEQQJ1KRQF7k3apJW1IEpHfRfJQKlqAW
3dyhbZqnkVrMS90fZ+zGN+XtQZHxhKhtPB+G4kev/LFj4aUinIzWy+zGNROTeWfO
oAP2LsrrGS2n2KX9uustXUxIhrYbYGnT+DdNLcxWKtM/sixpAi6kbW/oNy5qt6+n
Ty5NAJMs3PhRgYpxy5/pvEmJ5U7Ou7G2Pj+p/SOemWcD3Qk0lt6CPnB9QvpiL1dp
Y6VCH5FLMIVYhK3nPPHnVnQfMg+qpz53MKajCMPHidtHjaVWjMEPXkVDWXnAlk63
pARu6P8yMCZv4VqgeWn499yVo+ztLokY9AkYYxMPJVQcyb18zhmfNKKH5zincjVW
a5v2FlX3WPSKzN63dXLv5rI+88MvHkU6WQbrABRngtgmNtjMN1dTLyJ4sGQB9YFq
7vvhVBkdkTJwTrwsaYkfk2VG0gf4t0Je7gVx8vS8+579UADdkgxiZgXPaU/1tvNh
bqWYWRWSsLhsWQ+hLpca14sglTEAt0kAYtyl7ndnwQ5IQJei7pX8TXnDKdkw6Gb9
EolTE9+z+rdrFU8jC/6MgSpJJhpErMiGhMMndnkBoQuxBflraVCKanMU3yqKPU6F
8AagbGDmhSBJh43AF3ep0qjdDQhKT0EMj9wRM7OqKfi4L4wSEY90mZGEkafjZfUd
JoEAZ7tDu3St9Jh2EtgcFUwfEhFBdIx0qzIMC/Bv/rhSCBeombK+6NYcCYbewiCW
NarS/TMVDidyoLnIERSCN/hhL8s/fJ5HExhFqE0HHTSSftp9ATkjZlXEhKrFalbj
n/4Yr4ylmkPyNUEtCrq7Ivevmp5iczCr154grPcO3Sfdq4zqhSCK8DYdE1q0/Ngz
euS+UJwDiGLZPmUsLFfLxhOO5zTJW4hMtY2KSUM2SFK9ft8G42cgfVxLgNkjGkDM
rDt30o8VSlsOtjpXkEOzqI/ul0daRBM3PwVWWcILXnqvvGJzJCgUmTmq5DPO4QWN
xFbmFI85O81gLDRmriht0u8/CBHzA0myfuvMtEzjgaG8LNHbCVp08Gz3j+D4ygmX
C8eEbmtAyvIxXGVhagPtPCO97JL5tBF4iigU+5DyCgd8eB4O9pae75j31xXtFLVl
ECcbGq+7ivwVSX/VpDs327B1gj8Bx7aIvlsbZUxvYNbsuTNVblKLqnmRkrs4Q+YY
wB0qHKnxhOHnUB/c5Hr6KiSHY7x54M/4yLgASwEWsGy7q/45IcVhqJ1ME8dofMMC
ajggvaqYvS1aiCrMzRspGISB+EPqUApuBoJbYaCWG/v4Yd++0rm3JgCEnCT+tvPu
PKw1iI3FMYdpUAsmrWDOQnggg6s1sroVKZlyrH+Bwg6pnRSpzfPBnZs1WD0BY6Rl
0Mkcq8HSowt0gi+xYVd8Z3zy1Ir+Z/YR/K54xFQhrs96IK1+ejUk5eLIDNPI81yl
RZHWbV8jfe/8ZQVt/1bjIaBYr+mnqW9LrdH++E7QO4ZGTjFcGxbFb4MqEpanpHqA
f7A8x8/sGg6r/Kt2I7fEB5YRQRhuOByRQjzVGEZwxzB/AxOH3fffyXVwAqUnrz6W
HyValjcDBMMeyuUKfZZvcqtCLYA2UgSyAPTLW1ej6QKC093gnSCBScWXFgXt8aZN
0yZjiMe3fLX4jp20wtQ48K9rvHit82eq7Yzjzswff2uvBwwwIuVaqIEMnZHaQTv7
8gXfdCchRoXyR8VqJBPBw6vYrydilPoWwpJ2RkJsG6M5R0NVK1sj2d3d6Aam/2ad
IJfPP1yUsUB8s03ypVIp7w8LP17dDjlKVdsan6MAGmeHlJbLkELVgV8yWFT1bxjp
nfp9MHFHLpCnQn/pWkpKjIF30IORXGh2TXa9MegdosUkblPtjaidRGO0EC6OpXOa
1hGtWbFQd/urflC8wEXde+qxC3l3qKnq1yY3iycMmIJeu6UOkadyE6p65jyXabkb
lhhabwbjDt3gwX3pGQqYE2abWA+RpXBGI4HFAPGLpmuzhtnZK5jJ7uizWO8ZOROo
lleACi2iPyvsIg5n0DBv1vX/UR5iOrSTiFi6SFnGoMhU5BlEaRAYfZvnWB+2Smu4
LrjhUw3ttZW+meahrpxCwSaqFXzD1hC7ikOc2zVqiN4WZJzbZl/ELncViqUnEW4E
+bfzFQYCGjWUdiRII5d+lwcplrLtC3iGgNq9Dn/2aDPWD1keg2tHJRBNpNjUVLVR
9CpNkLcKiTlEL1XeXfaTFIT+3fxNlRJ/tbS0bUTzBctDiXC/5EdaCQpwMj1Wr6Ai
waGA5l6xQ3qIdWdPJsELzBnZmby3P4zmamOjL4ORcBKNtKxNkir/mn80MJVQlZM3
Nf5W0ipHNpp7WgCJUXA/C0lUYXKNPbcWDdzhxZshIDGVm1AIM0mcKQ/Xkte/qPSK
ElKCSu5KhbxAWuy2yapcE0drKKzvpqpdIryD28rKOQgL04yPFfX49J4UI0/y2DfK
E9wBYSoMPCJXysBfButCNYKE5cC7k5P2ndYSBfmpK16dkcjQM9Agd+PMoJ3qdvM0
6HL310Vry9tLFz7zGOtMa3NLkJUk9H4wwokzvHMKV2DoiFSVUTarx8KYZsLhpcID
RKP7AJhNPXQ/D6tuHWtIyAiooq8W14slklsgI6Ywscbbt77Z2sVDe9IqJJmJ7i5r
o9s6GuRHnRO1wzMKg3zQocAiozFLzHkTIin/ca9G2J4JykSO7d136id6s29Q+X1j
NpZ8Zza2iWj38ET8wLyf+ZSEvVZYcKeWx1QFbF/Yxt41qnYOPU+3o7F+xna06mtp
YQoaFr1NPj/DbmQZp8qWHqsqsVp0MUFwDFpEltFxfiv6DZsLMW6Ssp/51XXCffhm
weuZniRzJbk9tqYmEt7J9+9D6UqGMnjZFWVlhbHN0yp48HaoYDH7mKODA7wg/Yez
Ej5xwyakOF5MTS8ehZoCnUEtl1NS0DkUyD1yVpyL5VsGcKa5g9HjhjSFUkrFs5/D
ZS/yj+wmw0R0XbmEdpXWRyEg7pnbwW/1AweeTo/HDUcd51UMsDbZGSiawsCF6GK1
tQGGOyV66Zs5ha9NJSzYG2PeItlcUf747Atb8SgWCtLQzUwS5rHuOl2SbhxRHv+E
jazRDcR/JCIEicdt5V5bETJKPZ+0UE4OxZuSAwWZhRVXehTYG2O7lc9RNN0fFn4B
9fpdf4j5SNhMdIOzsKymdf0P1FaOgP20VTOHVIJ70DDdU3ObfllaeZHQskpLDd2F
eogwwWgqI6D+fhniS1Eo7PDZjceK1GhOHPdn5LV90VwT1ykrNjp5caHK28rPTq0b
8uPIl+HVf7AzYfPSUYWPkqZtXT9RQnxpZNrYKyxHhJjfBxrsLjLtA+SyyJcwkAzF
lOzRBd5FmwDurGWBaMcqOiHGLKrylCVDE9cjFZAAm4kGnrOvqEm8whGrWFjmJkUg
saBPDDvoZ89iCOWyA//h1tnDUzr1luHqoEZxpd8GMOoLLQZEZwT2eIjP5Qp5XCNf
XnjbdWbRt6TE35tfh1FI75EF4845t0wUWB2Z0DG2gfGrN6n5vDp5FuO9RV+TDTqE
afFZSw/OTH3Iee+CT4bCjYQYoNZ6cigizsGvpqMPqJSuKNKJwJ+8cdyhxexWAn7F
NglRrrUuk4ESwllfJtO7Zm3ZIgD8IAacs8VKCgOes5WbM22NVZDA76Dd5VaoyiP5
Jeq/K28N6fRyM1A/CMCWRoqPMCLtQCCXlu8QH+L62iLjPIC/OqqAhCvS41aVpgc4
HLROWeH+c5YvtBdNuQiRemvn9+1CT05lro5/Z4wI0+IpWtZer2ZRLMRyFr6ROnJW
VhrSiBPocuPREXOxMOJYoGcSKMf7S1i5XIeVl4IWLWMZKbqzwJ77tCIJnKZb4RIi
Qere087Q5JFUVl+fH7MBlY3BTCr0LWnqhH80b/jEY6PypjuviBiIPkuBiVrFZrWT
6h7GRA3SxUbJzsWBz7+tx0f0tmvpWpnpfQeMB47a1cghvdX9MZIpltkkTI/8QP+9
RcW+kc4XOfZurEnwcQfITcH621fKtK0qXnf3CZ8x1WThfOGlSR9mAVHizhKosYDa
0NKJxlfE7DbcQ75MimRPonREZUTYAKyYGmOLadDowinIaDeltGm1qZWRtz9mvHHp
ibscqQj1o57CUk702YZKeDzKEcwEcDdJ5aLIbeY5nzvHQH9Pqu22lI/j1Xo/jlt9
EV5gozqosNJ/OEe59pXHZZBsnc3liUwRNGJKIkXeEj+MGYpdYQp/Bma3C3p8UXC3
+DqLdH8izNdGWYh0z/+IziEd6MOv8/av8y7QUR2/WGCTA3CVRLFdLYVhnnCzF4Ze
HjBAbHghQX8Kt91p9d514GgIAiWBZoVi2IwV4sP+VsTV86ws6IDLVv0A1O3wzcV/
OxDf+LWk88GeSw2FcdkUZOzT7HPkLGTsIHIMRgsm8YprqJR6oVyUeIXvS/1c+I8f
V1lMbolSPXp5Ew+hm5zCs4tv7hrEKTDLhOF/w+twFQCXchnz92dGS7lanpapeaRb
BeIntp7PLtX7eMsHyF/xDx46HpDhJusDzd45UMJLEzWrVJ7gwW4EUAI1KcZwHMRv
CzaAazXqnbpgAB9Tc0zr+cpiN5hY8z3SiFaQsjGRutShbKOfuwymTPjlKGCpqwRr
ENVn5IeNTvgWkNZhjX5HffgHSz+NgITPPSBWXEfm4RdGRUtqhTxPi/SBTKqI6o/a
U0UC6VlCyD/MwNOqRoZHN7ivTg7Rmx7NLcwiQM1BJFHXaAFTWy4RmkuuUkqEq9/l
FzQFFmSb3DftqMcKY7xTyAVsPte9T5uKto4Vsj2+MEp0i7R2Tj/N5hBF60yGY2j0
BAgtxVjPu8sdpAcZ02n2PF++PmuYlHR4PZfxldKT3ziT7KYlIzgK7ccYhmehTiYI
IdvV+xsWVVhq8Qf76ykx7n+ThJeqISF1p7HTX6ZHYkROWawieV/ZcWXtah2lhsFq
e9qh9JKX6ul9SVIcdVwH+6i4injr6eFmIh1hmCYB7dIaIdILNw07UXCEdW8CUVJU
kR8lLe8UueMabZYDDPsJRgod840/UqML3bZxUlJCd9Y8b5eoN5EnNueO16582Cvm
Q5t2Xic6X+aFWpw/l4/DaFfr8pDRdKnqHBnUE3x92b5hHB/AD6/DL6vxTfNoicDu
nHp2RIrShFgMNmeoZslKAT0VnsKb5aaS38gaAh7i6I71bWuWsL1cBkPuktbs1qm3
VQHVzW4GCv6BettfER8/ddi4UViGdAfazX94AEsPzjfWu5dbDV+SnE4cwAj6Pw6b
VCOakLj/Lj/cIdFc8qlpaSqn/VZNQZhmls4Gf1xT6q+SRalIdaxwzWi5HL49yfXT
r+j8YPLP02i8jdM/MVFzcjeX9KJApHiMt3eDZLGXNL8cYjaM9+7RsyMzcehRUOeY
ax9MqBpPJaT3BHpJleIkA6jy6PiisLBXqY3gOR5Df0uAY2Jzkx1AUNOBe/B7MBT4
K/Lso+MVnK8VXqQNRwphE+SJE5hkSsI70IsGPB5zQrPG4U1/KFHSqxVBMi4MxodC
OJ4hf22CciXvmpDViwhx/DDHS5V9RSuEsxSYgwSyX6ZBBFiSX16bLYGj4gpCUnww
QOj2xtL/kKqelGv4d3KaYWdHMkhweUn4XUrVFByfeSG73Fs6IlDUd9mR2pbjcJBz
93ZyGhlnwabaoxqkmImT9Xypzb+Q9a8Vb1yYaZNx3iBgCAvhBPrAfVBmT/Y/oiek
ppPS9y45b+7fcBM8irlaxO0gziPZdBHwVp+I0jTbZXGUK6TMyO6C9r5s+36aEtKE
EoHe1wsNpvJVus8Bi9jYK7jXcoucP0iQj15rjXBc5TvNc9baW75GkJiLkCZvEXr1
vBg/wxi0Jrv79JpFMh2R9oVgjlWvSlt3BfMe+cu75gkn3+kYc6eRvwDTZT7Skbnc
vidNLracgZbcY9aGbzsgPyfAStuwc5QNuOHRdDFLy362Fc9HyC43UX2Sl2R8GEAs
7cjsFGZLlHdSpXcdCcjRGNQpe9g82t2B4xywpALPwaW5wDOLfDMs5VxWTIlK1bdX
es4KFxx5x59q/87mgia9IW0NY6jBKlD+dyEeP0tXXA+qOAc+GhjELyPtQ9WcRSfi
1mVXxjrZyEWB7b1s87bhTMdXqH1C6+MoUaCh1rYkaC8ilJE0EqxcHV+19Y5HMF+o
pyfJkr4D/e5QaehMNw/uB4bIE8yspyZTJX8uQ3RyLm9X1GDAab5Zs6/KMzmrArlW
5n9IGCtl7BSuLp0XGZZLdFJ/iLsexEEdaPGYqIxWo5Hea9EXf0LQIytTidWMoNpq
1YaJNViAH7UtGEDorrkHxJTng3cQnCIyEmdToFHjXAHKwMiYyZMuX0iBD2pWJE6u
aPQmWCi75z0yR1MqlZex0hb6eQsXhdYLO7br+MGuL3zD5uxK82KTA0cuTgtu7fc5
jB/fu2Wt47bS0eANs3ps0NTR42hoGRtL8FbPxW9hXWXDrCQdByasL2PxyjcJM9QR
KYnm/Ckin4yUTt07FrVMbwEHs/HMtBIzD4wrDbk47nOu6zv1tauahwmgJIpspCPE
ZTyjzglE9fMhyQAEn2p1224LJyqNgs3NY1NreIwrS6OYIGB/cI1Sa6MaYoKgXL2I
moY2IowZcQzyiSkkz4VcGKFD7vdHoiSjVOjJOZI/3f91fd6iHP7kqxMebMmzxTlQ
hBtP4S6gE1Pslja4Ruo1lTB+f/LR2QqRu6QISHFY28dHDcDXQPJeWrkz2MFoOH4/
cmrsaSXq2lXxY7KK+RbQCY8VAa16bgUm/8jPhWQIUfEsK0U2LVKKsnIhr/OwUr3o
wnh93IR1ttBfJY/73/C6jPnpBvWjLOFPSEno+xM6yHTrtVgAXlu0OYGuPsItoyXK
h54yGTRKsKR12KM2ilLCLNZc1i+v6e6MRz67S2+BxyapCXyJ9HkI+aYulFINk1GB
/BRthEit6CbenypI7k1mAjTvxdR6awu5R21RS4B/HNfB/ias7xFKFKPZTmL4zpzC
/U7ApJdd7Llk9jhWM0d5E6zRFdsRUPjxYohHGfj+8xPVSfypSfRDAcvNR8O/wIuH
fX+zJxkre+ygwWfR7dn0jlhHlbAiYUam5KJIUAGI39Q/HoEAtzqyZ4wytkCB1rFN
Eee6KayQdeWV5TS3U8f2smeo6yWd3ONtfmZ2wuP+FCPHt3Q9vSqu+rPjxxj925H2
AKEj3B2oVjKPsPIWKPwq++GyqM9MFz2WHk6rEBfGC+fIMfcHx2fP+nVffAJaalIf
cGVcotReav3buV8qiSFyp33BuBong1ECFtOTXwga2TYbPRAfcW6QyOi/a9s1KXL9
3VqWyyeeZHRNYrB+rgaK3gz3QUkvyAomlNscbqSmnWR5CldUUjdmsxD30yQAP0tI
av7bsLtDLTjOItiV9BlXrDhh24UeCHo7otuMIXOjlILpu0+P/OSz2FiQzmrDmfo7
pGRZ6oHHB79FVKdo9PlwSINz6wlYNjwXyveGobbm6tm9HyGZYEB06VutcSc0XJhS
hedrxv0e2teWSeuL9mVYlnTax9kUUh7So8BuvJbOD6K/OcJ/y23CRkU8ItQfQPHv
Ut/96YODA/XENPH4PXIQIkdR53+5HLfa9v07GDtUvYkTfPgpNtr2Oh5bpnFW3mDz
/KKPvQ/QnCc0k0ZcGmz2uO8SH2+VQ0aS5+MTEeufI+jc8cs5BRd66z3BgFuNEAHz
l6+WM59pbgOZ028c2f35HIP5AYgXfHf5ybd9okAMruOaW/XtQJ6K0OF6fsi+vb+E
Ec8KbthYT4xJji1DQViNrAlu+SeF6265VoE6uWbkE8Dg7NXqP3HrTP55Ovn12m0D
vntbfcq2v3dgqrJC9NdzvfmOy+hK1qnF7c7w6Hfv5RiBHkAHOLD/Pckqd7Xj0bdT
BGiQcbu1WpEydKhAG++pM/3KXo0gG9VMmIz8/nVVxLy2QRI8YGGzFQbGO3R5bhBV
UWPLaUmrAfxWHQbPgBn7/8MrFkozTuYH0+lmeNwu7Ojkq6NwUkP8+s/8Vq2WXzgU
tyaEE2+TSZxAwry5O+RyDfgE416kExiGKhm9WSSUI4HirQlrctdufcbWNQ0woTdm
p/pe+HJuT5DBV3qKRfKEvUhfjPxH5IWxarU0lQ/guuSf0i1o7GmJHFyjrVHkkHPd
iS+x2BTwW7ZtiRqdrY7/gtRJuWsH0MXlFFYpHiJV2xZ1+hv0YVWc8a29FvUo6cBr
IPV3bKL/vAGCWzDrbwPKTbqgCj3z6xk2KPzTTW7YRY45i+S+MX5ybaj8Iyb1OPkg
bThuAMXvcLtwVM0BfIQlyB/mOniero+hUScKqqKzkiBH984r254Vk+ZWhf+NGItX
TLbyIyVFVeRTuZC52D/LlVQkgQMwOUyD1VEikelXe09x3SIErQ6zYIhqaB8JH9N5
QEwWu9fxGdRQdDX2QXfHpykvLmGTin2JUoJxjKqPUtliGh4zq4c3rwp6BVxRRF4y
6SkwJNzUOymqIieP6bOf9EQgCFf8dhrwEzGcX9h+J1B1PUpB44GwbzFMz5Imvfm4
UDNb6I0Gx0zoqLOibO/AR1mlxp1ILK5f3XM2zLBWbxSQz1HaMgth2rd/DZVFD+oI
D+TdLaz9MCKV2vKBV5pzmgsgFWj2zd4TVP2vZIFUXnjwYeOChzlKXbVf3ub5IZbl
vAZZOXM7bwNJZNGdf7epBEZxRUD9fc11Jiz37YSx+y5BxyCa34TY8g5bQlukx7C+
QEEkTg/2VeLG89kqtaJPeINywokmCk4ykG5DcYOJcaT4e3aBeyV0LUAQg4FiMs8H
isI+GyL8FLQRjuFW3uiOeNfWzleeeUr66rUlKAJPIL0VG5nGCGNjG3mSvmyr5Ycm
ZpcoSDbJU4MCJzeDAUauLpQGC6tgn70+i8Xo+jK3zX0ZZUog74aMCV0CIP3KCO+9
oWgzwbBqjxLzVIMVAWhg6M588Yr3YbMDPeLTnHPthtihl5nZUpLn/fDHTEQ9ykM3
DmyplJzeZN6BvldvhcmERnVkh+QPB3x75dyW6gscFMvsyW2GF47CiQm8hG9c/u15
OgBfN4iQl+2wfbGlo/EjKoh37BN8lCeydEkTGK4Rv2TcUwduH9A+zp6awmulmUN2
uAgISFhyhToPbUgpvvTKsfMeE4YbXjZH/tKE9v+6/Xsa0tnN2UxiU1lmEL6k1OOh
cA14u1N0iPchbMnowu47b1BJ6Gz+QRfdzJJhS2kxXLAf5l4gLnLPKQfC16ouag8/
yp2mh3DcveL69CNfip4goxyk1RSeE3Jt9zofNqaT1xI1Z3xUHZMEXD7TJlH/jN8O
3AzG7287E4CvWLjUZswaQoJqEhRtex4yRKGk5qVsKvez0CC28Hq18NmbOppUbEr4
iR7lrpT9GvpvLbAPMhZBhFu6Pj9J5N7UkrQ6GI6jfxl22jjo8EAnUNTOXcIKPqt5
ufstGYkIMVhf1WJ4mw9FJkD8QyL4Bi6tZIrRN0B4xFSEY5QBNS7CUnROzuek/NGn
rP3Cz96UhYQNCx4ig+QfDgoc3W9rkJQUePsG7DJk1Vh6C53f280FOX0YLkX7su6x
yTCYSlfGlhuh1gg7kS13xNfspflxnn9ug7TwmIFidXfpECXSq0zMC3NJuHqJ2lc0
QxnwDecZoEGyHCyzcdprUfKnNcrTt3+5ElQnK1l0x+wzoQjlS7naG0EVapXvi3gj
4XoIl2jIQE4BjIypu9+iab1aMxXFbTenFMOr0+zlWpVthLqW0UOmC4Skkuvi/Vf/
X/WECgMKyEyhqTso2aXkuHc3TPsqpvTSotRonNchWaHXJa/JzsHjO0z/X/DTd7ni
94zSVBjESJLvzBsJGjWicW6nhAbXRDLDSzGiUqh1PkJh89wKwaXK2+8qVxU8zOmW
gtRtLj5JJgkjUBB70s0R5O8lku8uFHRDCXVgI8wvm0OF6PcvB6tNjr7iZIQiOx6g
INO9kRUv6F3ShkmAvJhjMhP6beMN0fcCmFJTgMB/muQC2FOOAca6xrZYq1gXFjpk
s1FFo7uOx933y9gfNyfmbsNWWmlItjG5eGieHUEGjNRX9SMk0PESG7yGSt//mExs
44/aZOjeaNxUozMDG9ATIrZbDcgmRUtpiT9eogGk819MoDg0PYSVhlqWOt32DHdh
CF71F6HylCVwEH/7hVnyYxzrbk2Mg/FQg7ApP9ItZG3aUZRcPW/irhZTWzwbwrIg
PR70z5HCUFX0Xpbj1tNGQYvemsRoyJhOzL/07FXn7IMAx+cyXK3mEv8tSD+Ygb2h
GWkvqyoDvERfmnFkFT5DQp3b8EZOoU6ShGHvFbkcAEYzDLVAR7vhOvuO2QMRXIRM
UKsa/NPWbAyyp99kcdjQGBMTxf8gOY3WFWrAW5qydSS1SurYNExL+tEVkX+lZ61u
/jcBIIR5k3TvyO+omIgjSClXRj9GT0ffwodYEsNBQz0xG5bm0eArlrbd9Q7EDGvA
siMM3WTEAXVdQ8MQH7yWfi3Pur0jZtq5MO7G3pwN32zIcjl0MbLW+PZLOIc8iOxo
Yro31mVLHC0uvtDsZhsrCNJpeUdzEr/RsllQ82ryeNy5MHT/l2I9LW2okZrK1ARH
qisAh4C84EPysZ9wakOsrOB7VV9A/BkLIE0YwT9IAi0kcJL8xFMOR6RSzVn+FLVy
OQ734/V9C+RX4FUj8MflTo4GXu6AL77NqxT7142+x8dMFOLm45GKQEqJx9SXczRc
ZPJWs2eG2VMuE9WMfV3xQmvtiv4HU06okPVLQwXFDOcW6rEElPOREt1jGyXZygR5
8XHv5Mg9EcfxHAoW52yF+dX5My8oy1iaJV+hfyG5n1RwuWPOpsTshy0jBBbjfKUD
OXhuIHbKNoiDQ6Dr3rkk7YXwq8FPJaQPiV4MnrV+h/CTLnIWP1eyuQD/FjkvB2nx
fSY2tbNRy7S3UqyTClBTdcTVsDAlBA3ZL/2BioJKdordZK7mcqIoduCQGwZytWGB
sSXIK3/Lmg/1pVM/c8kL9gnQXB+QuD/l7Kk/XMlt+Mq8Yf4PI5gReGa6vbjjabuu
ZltxSQl0hbmKeeK8DV2qJnyqfIH0LXs/7aud3qs8ptuFHUrMFNwSx+uTrPEgHOPV
P4zamfQWeBLqChMLaQkRwUqGSo3K0pq6FCnnM7wiLLCCjzX5UBjbbH9Al21I64Cw
6+X9cz5c3Aapj5OSBg+VvXcmGUGjylyb94siAi5fDO8Hmsi+xOK97PxrXsYtQTSV
1tKxQ45PDwDoOJghQ9ZoKcfd3zzFdlm8oiPhtvi8JWdOtVKnj3jttGw57n9TrcJ2
iLdl2+s/S5G34SJs4AIhuC88IGoBhsRnKRHiP1WeE96QbUppxxPN5afYDhOxh6EQ
xgPCdB37s4nqWbPeXDTiVdAJIT5Xbkdtqe6D7lyXXbpjWYr9n1JGpbWhjjvc0T25
O6B8O+gCcR6PhWYG2qe5GsQOQLPYtdsbkhrcQt1OFBYJBH12iN/L1hB0s/JAjxzF
55l3s6LFu1LZ9qB3Bl683NcEy0FQfDfAxSxenDtYxPSlZ8jbnLTkOxGjFYs9oueg
PYpIGJuFoIVMty15CJZTRbJOgzHRvyEElgh/1scamr/6Krk7E2KFqtIIYSIESRrg
U0AC8EgfQGkRbC/AutqLTgpY1lufdp4si6ABjFrkgMGCi/JG0xgRmRyciKa79Ell
VwDNvQ5qhZ2K1lYnia5esluHdAJbKoUhtr/+WPgM2qavDaW/Gl+JazULemLK1lVC
ZcWowqyjBoGL3jGPi4PPdhfAqileXZYWkqgfmACFV9vZNFcIA8KeO8YttV4unRGn
i8+Y7xNzRmHTnK4HeDAyJ6i3stoosUYhE6kZY51TH8QX9s+KZbXDQvNyXtSsloNR
YihpCeL3pRTay2MB/Lx31ji/1/3ezBnuHVitJ1jufECgmEMKUg4lODuTPOaVLUlZ
XpsgzlvMPHGrjuxY5YZi3VCb+sSLifrdASeih8rKj91de1nNqtREr5ithnIVuHbB
4yOJZtHwXUZ40i+irjjjqeoNek4K12BhPeuc+aqNS56cy0tZH8Lauvt0PGn5T+Y0
jSbTbSzAQ5xU5yRpe3FW+0xi5Sf9Q0XS/CELGWliBvvchNxl7KWATPiDchlkzL1P
eSUnVM8bc+N3PUgBNO0zit9oLIm90sreONt3tH4IoRJH3GtUBbIAQrcIlvl8tb3R
aw2GGBzi0lA0OVhaCfvzg+tGAUboXVLeEm/bxHGKMQIoCM4pBNpiNmiAGey55vkp
Ki8l/xiQrMbutpL2LBra11AxKw+TVujLXbl+2bW8EeT3h3zfIsDmE9ZWkOLGBkS6
MzWC04Sg1uq30CXLmrkEpiT4lWG3rSJV3kmQRbGqjfLLLQN98P5yIm7YZ0c6kVzU
DopKSp+bzX8D4H4omUFcij+YdHhTWOrvhAvBjXLA41kUYEKHoneVrxzfpqyWV1VU
NFnSWqZ6FMrv7bmag6eeDhyFdI1Wz694OTY3OYi7wtMiHoF9nQk2yfu3Ax3UCbWV
M3PXBqpoG4MfF5aMM3unBZvj7CrIoOeAVQhLgs73/xY0zfZ27qfxbgaScGvMQhok
v/Y+AzpoH3GjfrB7c/01w8pbaw+77pIv1JRqEFgVnWvDABA8IFeKg5/lHnT35H/V
BqnNvO4rUDlBKjRW/JreXPoerDqUacDX6bC4fqVMz2aKrMVDCgeqCAIW1x1M9mHE
15OhiLSPe156NtlH5DuK+ewbQy4dw3UWAQHJAkbs3Nsy7lH2CxBTbz+8sAoBUzdk
8VzLxS0KXn1BHrGpABaKPKU+P46RibtVhtEvjcoIhwX8wtwBC9rQHErjTkzSz0Lg
BewGnX+1l7fxH620m+axrLk8JNeVjAjYZsoGJGkuXcV2aE7rQaEiWVLxVQB9+aiv
BvQaeulfu+PjF2S9NroqFjxZRHPXkQa88GIrfet98YJMAskuz0zreidtHKnK6SoS
yOvZAf1Vwn/jWrL5C51X7ZZB94+j0qPhavrzoSjc52Z1+3Oy9YsCMvKbF7kMS/4Y
y04bkVG0oqgo5YBo+azJhSSBkbFZ5/sgxT4h22qV5bwV95EmyccuDymJmPSC9dB+
3eB/9hGP8awrHbFUzKB8JWFR+GB9GZwtdUQ+qmCKxINGYwDZ7PLokjGyIR8q9KS0
cmwyA3oW+TIy/iMQIuYs4M5hZEMOEe2qA3eaL7cG5Pi9fXT51LPYoWTqlv5JDMkd
7JdZmUpTyylbjwaJTOIBWAkHjGVGs9HdlIimxNvYKMO2jNKAxxnVd0Nzby8DQ9Dw
3gOrWROyUcXKVYOcEVjK1FN/LAoWMRkOyQEOHkwz1i1wsCd/Nrnx9IuBv4dfhyCR
NtvEEU555Dp9wguF9oe4mEHG2uebL9Lmki7RgezUkyxe20xjU3d/PNWoCNCt0nVT
zIjbPErbMYM2sSI8d6o1CxYWtjAatRV7lFW3xQw4lB0g3KcNgtFiGQZM/XoYkDFK
NSFc2oSNbzF3LDC2VBtaqz/aYDBbUe0o3YgxyhxZpBdIwgwS5IAximubid4LvRvw
Lh51gEEgAMLSIV5P7flyk3IRIDSdMeQGXwqjkoyNTDdJ5zP+iyx4K42YChu7Ec4e
4sII6UJWX+fcuC2fxpBWw54FrZBvYrzH2hnDWIxWdhYwaiPR0E6Co3ZoDM5RmgH5
okVGa0nPMANg3nO0HgmaPqsZ6u7ozglMigFEeo0wwHjjtlFPr5AdZdB/vIMHglHC
9CCA01FKsQlFEKIl0iy/ovqSeKnL4lNGHKDqU7P7sows6V98zGC7ZLx0+IzJ+aBC
H0VzE8yJYRXZtwf6r4aqnUVp4WTaf88wNvCwiEbFn5RpCMS1wcrboZSBF71g+Owm
ednC7FEz7pBOa//ktQUIDQOuQ4eX49MwYpcUL/kU/krNdCSiq95Kz2CF7+ggvsxi
dGBGN8U4aCPJIXOpZsnIHlxHEcez27pLIEFxgUUaNAVWx0Zrhj3BV2Lip/pZaUJn
xj7AyqDm2d6m2MFSDt4ye5KlxriI4g4eKdPyuw5sBBnv+EEZ1Pp0WZfTgKLtBD/C
k/NG3ByVmtJ+ACCNYv5QmxpUBZc6EfN0XSSwCO+FlgoOGfrgH5d3ohjSjjdX1CDN
hhONjSiiOV9UypfqlryPKptbZzVFiWt7yaQsXuBr6H/84xEYinIgkFlcZ+UESTMl
pCi8Z5fq2v9oTmjU6CjtlXHCYaH0PJeyRqZDxKYE1OTNIfZuGsrlJlN+GhsHhI0x
c3ScvNVnm9V9IIpu/1yk61nPoCUT7nJILtE5tKXmtk2HTBVblnOnmL4kaMMn+XLx
TMhNhvuGwbho8cleUaxwmtpzScuPzSNJpocbxyGp8WlDhHp/nsGr7CXudgsnfrIG
Whypj3vIZPuzdQitooTKu7S20Rt4UClLi4V52qVLrHgJv6OM63Ma6U6eLBsToOCr
UDbFWdKkNWeTDOt/pUzaAmKEiheA5WdUiSv6QCPUO3yjZATYFuZI1s6+WK8DphiG
NYu94Dgps3S64eT5OrUVEaFPaxbZc6FGFVAR86CXOsvtbz1nWgfruYzilNqVbN/C
bPa6GyuiqrXoEauXzvRemIqrP9YfT1UzfS2Uq5UeHMWbqfcJZG7am0s6DFhWWlFT
d0Mfz3rd+rxlqRdxvu+k1AxQ5EZ0ohWPUOPKra0U5sczvX+MZdIQX6M0PBCfVtZY
qnBcbEDT3KnzxMnRJ8TR1urLC7vaUHMzOG0B/Jl63dJsv4xwPZm5cjqD73BoLAoG
HSt+L/jjJCAQEdAb+QwODi922TCPnteZ2CMO+QG8WZ5oAnaQAO6H4aJmCAsvRnvP
Om/QUTN6DldmsSHI6mQLFlwjU+ZX62Tjr5pepBdJGhmTgFVGeJvFFiN8FjrXEle0
ctrBfkpYqnr3RPRtE0zwNKxUoOoa9WcQPeoz3GkceCNb2RLYup443I9aW3+xqcB6
IECp8V3MBXrN1gEenV09723ysLnSBDvbHYqQFr+kQi20l7Ldl9epIcMvqXeJbSen
Df0rv8d6c31XE1N23ycFdqlyV/qxMq+w1jSOR/w8p2AvGS1ykbax8OJG+HmJx0Nc
Ku2GC49ak8/sea4hdBHEB8VvOIX0553NsI/swEloLiw1Gy8IcZSFAPm7/8W8qmOO
1Jzo08kkIK6g8v2l/V1ukkAMo55tGOb5wRQpcGWHYfC38hSUFEC7EzkkwoYEReHz
9xcEgxqoUb5rT5+yaRmJbuUM6M5Z2LxTQYW0m50CmkCHGpVhiRRBZtenI9eraPh6
WKbS0PMhspkK0wJ66Klc2jsDEYqf/vdKiYl3FiJi573I6N85yN/druA+19CZ4/Bv
gqyG5IMpUJ++w8srl32yypTxsPLta6uvefC8XO2OMDDmct8tz4hGYfdpgBMFYnO+
6j1zuvzN95utlJPH9BddVCkWf73MFTrl0dFuQYGwDPq3ig09VM4w5Q3tRGdAbmo4
JTk2WipEeez8hzpsxpL/6WIAG27LSuqljUl8+GhsI1h0fVBDRN7n8JsKbRoK/d+w
ATtVPcQjrT0HwBqWSNRt3h2LMdj7jOo8uAAEiq+UMn3tElPqhAF+eNpPgzu/Y6RV
6A4gCKNGeic5akp6VCV+u3iDzTx65euHH+OdNkne6r4q1ziKxSS9mjpOnN/jnwYG
pHO0qDQHTh1yHzZj/W24YERD8patpnoZHzdPUAPd8xI0KT51ku6QR+WWHUnz7FRv
IBLUE7ebKcHlpBoPBBDHwX8Wfl3n2udAPzXE863CIsVG+qSslf+JbNcHOewp26W9
2zbfAJeIv1ySrHjVqi3JISsEukdwF3VmlfQ9E+kIodf7Ui5cJHG8bWH356Ikfk+N
caXgLYpSAw3AmPfITWmcw9Yt1fA+Pd8vKAPwWhVM9/QmZVbwtPbx/fAM2nc05jjJ
+uC8PT0oRmQo39NS0r5I1QdH+DcNbSAwa3fkvrWW0Ih+lxcgGsotBcHHkTZotpfh
fL+b0UjgwZCeEF3uzOLkjjYyc8uGz7wEwAiRKNMpql0iTzjrrkjhApuKSBrbXN8x
vugma9hkOUOMVTr/q77Eegx3sCL3Bwqgx9xGe9G3SFGKt/FUy/UkLSLHJxkv8k4D
GzaxGz4xKEkyYPlHRjDH4Am1uztdI+k2n2DirM+fHYxcVoYS4wYvE7Wh5e5ZBl7R
1dx8X+tjqW6sy+2GbqjiXzuCOJM1HOHVDCA1Ax6HHjlDDisZAiVFosQgqmBFlGcC
7H0j+alfrKho6SUjbbogDrql9riKItpa+/jh+F7C6uilpTNDyq3zKLSQFyLI6oWY
4EuB0b5S4pfzDvmn0ZDa/oagSYEeGU1QztOCyby1sg1rzN/lLvOCTxD31FPIz1Hq
z3nUV3HJQAeJSy2qUug6f+8JBxIrkWY1FRxoKqJHM07bHzJEV+HMTtD/ahGaNXMh
l4JFCyib27D3fEBEkgEk+7qdzNmCI88//a+uq+q1bwbLyhk1Lk2or7jAk/ANfnDF
AZFBHhihMOfusD9S6HJ645ArK4BF3LyiY7+vJauPCofc7vFmS89Wa4KVI2P6lbxf
2z4wIV+HfkGUr3chw0QVyBefHKKMs5wPWR+5OtYWolU9R3lfd9l2cIOmEQA2+gDW
aEEFYzexywlKQUcwiFDGaSbJXJ8mjxIeC+QHxtWdEo7UExbItvqrfpusKYcBJjYp
jbGIZiY9ZqquIpvKG6r1EDAkNJyKPwjVPZ2zUjyqtuP902Bb+RhvjX2pjTpE0/MA
5jrcfOypM0Q+QKA1Kq+2UMvWTFkYs5NYs9a/mlYMsSZSQjBVhWO2uqFlv7RBsfXf
B70NpsZ0T2soea+p+LehNrK4pWmhY9YOl4720zRa5IfXG+xueDJWtiHujZ9QKhqU
bFc9WbwZHc4VnTnloycBDQWrvuVqoDzH1T53NhIHUDk3xjtAXnAKYUXbTIEkNcGS
WCPRbD3DFcncnq6ymDzj0+9PB9mZKwQH49Tmk8gEcE6sanxqUwuCbwyIeAB57Oih
LLgb3IHJQRinAxhNUjCSCmrgsx02KCdpOJbFDFLkjJYbaPproe42VUdX2qLc2mnA
xoCpmgdvCauC/DXmaUXRfpVlhxe1np5Zgm5y7nZa1SEF9tHocN13jBGIFbkAhCsW
13FdZXJbqNEPCwkyXCcMTQU1+/DDtNw3qxKYPf6u1WvJL7ZnqcNgi8ETBV+u8b91
xd7idEc6aCPYqX3d9LlAUFvyqRIUrRUfjgWDccrB0wVkks5nfmVFQ0Edta4dN/no
LNZJPKWlJXtU2lv34hSVVKIJyTf3M8seMOCgCSjpTK2gGRPF3kqY+5hnXDywFXR8
tcPMLBVcxdRcPlsBtoDcXjZkvmTyVU6Zx8I9m591zLGanKN6ntvrk8dwbS4Mo0/s
LjTSjIUpYaJIbW/C9cdLgnDnBO5aVQHovSz2RWWSDtqD3dvZ0frLepga/83h8Hw5
M8tu6TCtLwrFAwElt0Nvn4b2qkNb9Lfg7E3346Unv2xajlA7HQS+7HwInpebjfRl
LT+feRrsD5B8uGDyOi/m09cAv8G/WDuStXNrFoSH6PHI5XoML3mjh0ALHMOJnuqD
p6z2sjcs3FXRiLsFoVS+Clpl6neFrMCmCPxi9HExxfkJTBx1yOTn6/tHgliDCmY+
D8ZHgRRVE7cmV5w2JLpxPB6QRJkGkxMkChUfGTqIGJ6NOzxrJ+Qp4qtzP+TFzwjS
j84CoOpjTJkIP3mcNDKfR7BTlLGpCN4Xmbsjzxvwhieg92XR195C8ifrlCGpKMuY
5uykV2cPOFcqBi0Yi8FDl9INgt6V/k/sXAPuoGuV4GeZYDxL03Vcc+YCVdFJKWVp
5WHD2F89GGe0IzaiH/vUQ9bAEmXNX6Crxkk7oWCxnI/mHt08WRFXkVoNIMFH/+Np
kSOQAM94d2brQSQIMSzmy6QN54Cfp24eoCa1HNPEzh4Qo/C+Bdo6EU0Wim4vQkvY
BYRYQLdaXZzI6wGMJpXMKsFx+aDx+SlR1lvNEluktcJZfoTx15ITClzKCoxaxgHo
NsQg/JcZl5zZwxygNxwKqejVI4K7HDyUCHnCiv8PS/HfCouKwKKdoWaPmhy+ZK/K
xgZUPp6hnmeV555p4THFDtAFha/77UepWqSdfKuFsJkfLMq95TSwHEafcp+4HMCA
FnuaNpY1f5JMss4RQwJx0OsKqfZpPQPQt12LY1CW5yTIRsicNlZvo0oS5Tip6xJ9
qKg1+NTnO/lolLOIboysgYkSNkW+QqsquvK7PkIrGI8Wymc+78/Mr7KUKRV9ZZtW
e/N8KTnwf7W7PCf2lytrRAxnE3Nr66gfYI4x77htz8uzjmICZLh17Vz711NoJLb1
OLV240Nr8r22NTSgBi55TdxbWXts9wwNeUAbJE0J1FRR/dbwnWQCuJulFQIEl28A
+vnirRy6Mke5LM4b08ZTJ8LycAKsNGpZVPwt/DjsofESY/avoCEJnDyd2bZT1F4U
uUUNYsaHzVNARj5n9jSUTEUXIaVj8XvQ7a4H5hysfgrmjChEqjsrg3lI3bTSDqnO
epF+ubUJ/DkcYNd2988PiHMUfMre6jij/3M9BgPkC7lvSRID8m8/s+l7lI+f1xum
cpyYNcdQSAZsgjXAFpHQXmh5AZxoUFvxF+AceZ0Ph+DFOUTJRdhD0CmboWfjM5s4
HiKBdu73GMSfU8jbbmjdWStvaS4NSecMSPzeUBN3uHRpcxCgyVcbaN5C+xmC+6+5
r3DYRyCM4i1EiRt7FB2wpvXlTu9ox/umVWkrSvUtBua8cly9Do2cHR1j+lqkap2A
SMoGVlqJKKIvmsmbZDhYEYXqnJus4n3SJQ1aRUohDlpN0NrRfXatlQNgxKr9Z/bs
hAubFymC+UZo4D8bSonsv0bZaa4btpTW5UAf19jA42P/2MYayJRYqyAWp5e0HF+c
h+KDaMWVhg7Y/z8r3u+afDN9PIJrDsKidP6x8LK6TOIZbdTEFiR2jKDQmxS1HwwO
OyoKbX4//N/A5hpl64nljGFa9yZr9Bse6b4eMPEyDTVm6Yp61syeXJ37gnmi6BNn
T/XwbNzwwIJ8I0OgLj0kev/UsRrgmUqbBxOOvkJxiiH3HnXCsebA/613DJ1/VbI5
9LAtApxm86JF+z19NsE2T4aP+d2RMECnDkvz5ThPq3R0mhU9npSKLazFnv8G5Q2Z
kOt3guOZ1z8opMSkIhytvgVokRmg6e/LdOZkTkWgVSX+kzksAKIsBDG0lPvgG9aN
JA9zDa6FiG8Upbo9X+rUL2POFV0dd7xMhf/ZBcnEe1MdGlBP0FDx3+pgHv4e9RZu
F2F3aTJ2NKtTewjKIUouFS5MryLQn0Aq/bJ5qAnnQXo8XUfgNOrfAccC3YQsoroH
geJxYQhEBH3h+1JIHz8FaBaXVpSV9M3zBYn2gn+doTF2qexAkJ+ksH/uRmMbNr/m
xn73kAvv3TZMEWRn1n7B12j3w1dHuc7b9LMsr0d+KhMMEa2bOSzSpY8+5DKI6coc
WDuSe2SBaVmxeh7zVI/ggqx5yS/QsIO6Z+XqV6uIfR355QAoO4aXrCLD7PA1pdpQ
ciIJSIbqQo7c8lW3PmYPrKlopYWbcwtiuqGM5uxFBLZEiEeGKI94p5YgfuI+M3i9
8iRaczvkUJ+Wx+ax3j4sO8EckS4PKjtcgBf6B3lFgjDeIiIFnsZZ25zV9Qvp1LVo
Eg2BEbZvMOpPJivxCBb1ifNg+tMx+tc5K8dj/6maoYXLQg0Yk6vVbOtWRZ7mM1lz
mlTnW2TE7tjtSX1cgtnkKL4E69j12Ct5yRffI7en0Z2fAU5sJaLfQve6Dx2wVkxY
z5HVxKad6mvKVjvB/Q0rKc3DnUD9Up/ucxNmNtpSu+TEJbOmHMIGHZPySNzdcuvl
iplkyj2n5pi/AlAkXZbAKlfGvHjRRXsmvH87sdU9mAkvtfePVeWdjWBI0MaqIuto
e053CGo8qI2Jd4FGwIRShLB720f+FuLPTlFmcYkC++rrapvgs73GxzEnFje/Ofxf
/2lKhyrD7qirFOyheKDwO/Y8XXzA84QQG6KSL9YUNfMY0+jdMAccTg15G0lw4hw6
U8mYW7eRn0EPDI0hAlgTFD7s3erjhdsaeikpI5K1Vcs5kU3RfCEi1TAtbjnVhAis
x7/nU3Lqjvl6gLO59sXSJG3hy0OEGj5aZOFafT0/bJwBRnv9b3MnkHOVWeRj4BSu
XddvNEH5qLBdde7GSto8LeumlCuGzn4HwMFL/OmRH4bXIIuNpWGwSl6ke/0l5GNT
Dj4vByxfbaH6PhR8vtayR5OYW7RLhepGfuBzj/Ae3xEovJSIMqo3ZFpMmT1US5w/
AbHmuhnABl2lwvBaSUAlJIuO4bUZhIDQzU5cUUs+Dpfypww9y/1oAgTjpeOsY8+e
cPjRNdd6xj7I/Ki135aWXlxgf94aMcACPUREWaUFvm4xl42ac05x90ML68MA6Th9
vQwyZ4+wUlkYC28SCGa0MpCNpTWrMFHRRpZtAk8DUCxaXYXLmC/+chZ6qxKkNW88
NFYWpydMwf7IEYqrwOR6rW8TSU/hvAJkhb7fpvecS4QSZivBy+hUW3YSwJ2GLaWD
LM/f/U/YNy5In8WAYDe+OLTNqUy+POG4YKb96zmxySRT5NUHPobDlRlq35qYJYeV
BURduZ8ACCgzQelSmgjvg4t+1ri7KtxDSAhVqWcPnT9mXcJHwmtEfRiwIHNfiCru
qgppdZpKV0SXFgpMzu/TcxLgAZNpvcKWuaB9hHz7YpaDIXfCVM4IhVzOjs2WHuvB
umQYuh1bxaUtJUxtXu/LcyJ5rqY84IrKMSEmwk3ZMdb2EFljc7nnMMj+L/yu5sKz
ZlJVPQBF6d4yxIkSz7ML975DxN4/GxUzg4obTzowoUxa5+tr+x/mXZNvlnq6x3s8
N+91rTjHrFMBtRb2JHVYXgXlsuWQnex90jSY5xRHrgLZ0XBwu/2lU6QP2yQRxnGG
NbuYjEW1aOVDb8GB3gDuqY5TkAo1USGNLOtBwgwm36va5dOu6UzYrhCjhFL3aBVH
dThIHln15SXYPBP19yYWv495yQrvsKtkUp199SoCYnjPuF57fWLcg7I2FRZtuMct
SCz4fATi3kx2hO+kB+L9o3AXOik+VcL7XsZm7siNMAXUOqYE+lbIeXFvQha9QCd+
7h0uXr/psACG38VeBxWF/lheFuJpInzT1TVKa1Uszp536+SRcpGOW/rvaPfbcZVs
Vpl14yhAgiYkLj1MkGzxGphRbZubq/XRxvT6X4De4wckN7rfpgWkUZ2B3qopnUcT
TS0nwvbiE2OyAGcBZQJFCN3smA7HwCo219cZ5ajuQG6gdCF+cz7TcvowReJrhdF4
UdMwvKmfduVpPW2Rur4z3LXvUQzQquiJshkNUR1ZkyqEBpvqPWmE9MauVmSTMhFu
2AGnI2wz7QEZ7rvGHX+2J0fbHy6/iwpcgfCfZFtpLoaIrV/LHS055/3+nAZkPhDU
uPJVYtTh4RUeljoxGaBYjB1UWsRDYadEoaN8cViU3WCSRmzEM/Jdkj+F2L4QhdnY
f31kIBlZwHa7a/7ONVxPppx+WvnQK1ye1o3ON6renIxKojDAPS3/UHcrE/8yxh+f
Mun7Obb9SvGA9vgkOIAVvWCBWEncjaR1Dj6OMk6irNFpTk/F66wzOBmh/7b0362Y
Gu3O+tH+HWwh7QqIc7JvUUJkmxYpjv6xLdD2PlWQ/lCAii1CDFDBcwuI5aPF+U6D
S9x1gixEuXFw0eDr0vp2TZV66IzVGPDVmZV7Dg6W8pocUG3Lbj3Q6jEAqKfb9M4k
wHdngiPe7H+bIPYDFLdm7ShEwrqsoG7eifLZ1Mnm0PhQ1MReFQ1+acSyrxCiKcLT
giSjEe4p16V+7EfUyLcPBnahju2B2qMJ8QtNrxNCOtpwpOvqSMxovPOmw3Hfk3DY
WOa8XI2MihuQN7YRnydgrcM34Dsdlv/BW9f8V3z2wn1h/aCOM14KqR7Vda7NJx6q
yaqiTso+1hQvOfQ+nsbnCWLlBA4EdI2QU2Y259KwJT6aWsfawUoVbY6ao8GqWSGp
D1727jsFKrVXFwo16tm9vfdBf/d+xhiVTkmcIf073NCYgbBM7gjks4sTf6C4E9UO
8Kum1gMHHiXqBLzS37jkswbwgmFZcZNyx2TssCDXXpq5vJxRNQ2R+ERnsCbG4HUW
fvzsBoH8jI3EFQyQ1uoekouKYhtogsEm+WeKXU2XEZnXKhjvac1U2Y8KijddDtCu
nf8RTUsQB9BptLDYJYHOmYNxgo2HE9+Eb21qiqvHlVnqmAS7mVtPoet34xYjnaD9
qactW4Bp6p6QvFV+PEtYzZvHHQ0CaDRlFKvNlFh5AuDnS0w+RKG1pzptoJZ9j/V/
VaDj9S+VdeSoKPnaNTrSxKHkYcxAF8BZ9L7Pka/BxXiimatvz7bjY0hGT4jgScu9
w57wqi9W2WeVD4CIqGKi3g1e+yl6R7ZjOIHzBvV77OzMa8zbdTjHqQ1xIqrfZyI/
QEMpNcITBywPsKjc25yQ6N/2+ACUXH3cpwVxn3ctvaqI7zJWZ/O0Y/TB7UWeXtVd
ZV1755B7HKPvfoaveR4zBneKxFO5xRtoUl6BzbQdkUobRVRYk+/DGvWvbsJPVuIU
Igl9qlh5qprE1WylOo1Ka9iJklOzQh5LY06PHnasO3PhhrKGnbuxraT1FZluKSXj
3VL+p8zZSVSy3qTf/nzfRSpTZrBAWFuZuRWIhAhRnweAJAQv6Mq2cHDdwMJEgTZc
jeQ22tWEJ3Rhj6yVRVebvfifDGF5y0sSRwdxXb76G1aBRknqoiQ+v5ThBh6ScoPj
PtgE34zIXVF58FeuOFgr9l8itwQ1jcNtUPGryBGGft+0gOfaT7F6VkEgPle+rS6p
bozNpyIYVFr4qcEvISdM1DcT9ej2QgGDsEiCUUGO54IFIDy2bAQ9nKAsh4OVdUex
UapgcOX3HJTAMZ15y7Aj9vSNCGYoMvhc8UAxNCy7cwNtixvCD8+pkX+1MWSRASYV
Ym1FEQXTY4PnW0Qi9IYBdHkP3Y+6rOC53k9TIiClXi/PtOZc5yOA08dtH3OlnFRi
jfhpefnv9yi+lrPyLxtspQ5BJ2yjX2B6hUmKHkTdTs3DdSTgT8Noc2VHztrqQ8s7
j9gnHPI0+KD81IVd9M18etrUFX2QypUQc0WEp9Awnbn+5Ub/S8Ws8snlPjb84izi
2bIML8lFeSa0sEdbTnaV78+VfYU8LG1HpUCQIdLcPt+vQkiTX5Dt02kah1x2Mvty
aNhD7AYAx8w6luXA/m3Bqu7QgQTrOJsjoOQi1WeGuTd7H31Up1X+iKdc/MNikgH1
wxLVQH3DEdbZXRudJFqMyVS4jnMEJeLNyKEuJ1D/sX6Pc4FWclu03el79+wJswSS
w+9yH/YBcOP7GGeiawY0ZKhkappe5IiGqrFDSMXhVKHOpC/9TU2VMW06WugHpt+H
mi3a/w68dLvgTkECz15Xp6co3ZzmIDmCDc6+NTzpz6q8l4L+qvHwSomD/5D1+Tfj
3wvTp3qkmJFCiJWjFNEQH+lyReZS5oCdCHfphuiRL8+M0mQaydaww5L+ytC8r93B
ZAfR7dzUrs01DkJwa7TLyqQZ+nciUR9n57l7GMtYlpVNj3JCTfZhF68Que2LrQGJ
+yZZhvdPbphmxSxJlJPQAheOLedDTo0jTH4Zi9DJOBbklVOwAdKi+YbiT2f2PYCg
bvS6qDd2LvCdVU1gPDfvdDAwLjj1YzKeOGvlw5BzaxDJ7J1c0n3YIIJU21xnySzF
Mufzm/tAa4ihDAWROyHXyDapXy37732InexcmB96xbC3rDyfVj+C6H4v/YNsj63I
Dr4TjlW0XOCBs3fggh+eflRH+J+kBBcd2BLsjf4sroo34pJlP/gMr3m//H++DYQ3
gv7ayW6SYIGh8CEAvloQSkeTb0EBItraJPea6K/CI2cRIPSnbsoWp3DIXM6HXfMu
yA9/5kvGXth9e2Q1V/bNTMcrxVq1OuTekMzyegwmT57ba4zF4ZWwXBf9jhrYWIf3
6TSIx1McgcKWE40fhnKiTjybxWPZHBMj91cctmef3tzNouQgEYza0voEP8rktVPf
I2856BEIkSYAJ4ta3JAy7dmjA3Z2aAww85i+/EguKQkYqCd9td1T2LLXhgQCqtOZ
EHpHXiZcAjJSbW3z1HgtNnAogScYM8DtgPuqF/rro4J168uBooUQJfyB4BeFvhqe
VVN8PhhEZ2369O4Ldakna1IfZEQsSlIyYAsB7X2C71ANNhU6tFp+vzqlqhcVlGjA
LmliLPk9KeJZErGYe3ckKn73RAosSoZ8bFpi7hi6RDpi86XIFIpw8ooHutbAzEbS
KM/2rYtLMNTwYZNl9HGFKySWNwxYDdZwTI6/3KcsyYCtXga3iGaSzm0jilHshXPu
4DCoILzsMFz5XVhLyMUyKjJ1lS3GYCJw5hQt15DSFnSvn2rdaPDjVEMB4BfdZ71t
xX4bbiuZOBvPUhpFEOhcazntwxVdEXt2LKSbU/YcjHNDAAH55eyTGysqqE1Lmwg4
wntY6n7yWvJDSy/rInXD+2Dll6C90g940a6TZXgNXlN0qA+s3VjWuVVJp3HoJpaU
eDxR6D4YtOMEgOkLOzNK41kVcn6tXPDcJ2CZoziUgz3XZC8c+bxzJcG5x3KB0H04
4ZRAFx2YWctDYWkdIhnRadlthGdi84891FwahTMH6qITYTbx6Q/60otvevw1HdIt
gdIt4ybdqx1l9uSSge7BULUiEjGzFaZim2lpv4R084ZNE/utbypkbFk9MJB1RiN4
GyufXxSo5YnMg4v6YQwUs77VQKbb7koNRygP7Eg9cgndCZIG8iQKVXP4BAyngs3t
pJq48xLC92sWSWNvpJBfYRirKuoCvB2ggRtqTsdBS6cjiSlJNYnYMi2ulrev7RDA
mxf/JsNLTtsnefvZI1BHxGBeSXBuy/jgvjp7WBxkpBm55RNocafH1vg44XotIfjB
zWD1IXT1ggNzP5X1SJdVfLjs0T9ejo5ArnaleIvbPqPGiM1KFiR0KKLocebiqXGt
mJDvsN8s+P/0JrKQJRKObuFkpb6OJTbxyrv3vC6ItXbav7+Plod3pB8WN2fbARiF
/UMGimVIVOJnGyY7Dp/mBVw91MRnd+OOOR4tABHnmyQ7raYiQU+ZJM3W3AXyvecd
I4/U/4s6J99ZNHXIO2Fww8nCq4tGk/5CkvoyxrcEa2oXloQV+3AiDE/++WOmPJPa
f2jDfeyJ7M1Z7hgL0lDfZrPNZp6zRKCxrpqRvGZDs9DElGq8ug9jwwJUvxQt91YZ
sN50DXLVam6lgqcISy2GN5p5GIghHFVQFkKRZk8PmGtVeRrqHVB9i6yyhSpqakKc
4l9MGetgdlXOo72vxZKO574Kyk1PxCeZcdbApIUQ9tzdx42K5921WHf/XY7V5bdO
8Hryxf/rfw4C27UmmdNNuxPOaZYg4cMFQlVtzvrd6lc005iVlxQO4qU4EeMQOe2u
nrhRGweZ0Zk0Ul7X8Erw1s6dPisGiRPQeWVHDjr/RcmmZAT4T1Ueyr9Iqp8SLFjL
bW06RCl33XZk27mY5xks6jd9LbDiAAwIQaCRIUkVPhRrrOJFnq8RMO5KiVAvpJrF
rmn4VdT0JGkFbwwJDdCVLHmrDMI0OsAoVJ/FX61PgYa8ngHKj+TJt3feWfbXfqO4
QAf0xKuc4o0p8YInN2/MsZM0dbZ/uIqDxUK6AYL0ZTW7LHUm1Ma6qXutnZkrwexD
FubmPEg/bidTyPrVWJVDDYBpGB/HbcJzu6ah8zlDwYksrHd0Vv9MVv6yRV56+f3/
IT3tbUowlNiOfHwTBApBBmUXUATrVsNtGCy+LP8OzUUo+2CTB+m0n0f/nU3Y6B5F
1rsPW8gzT3wST4+Op8/FdrwUpxOf1U8O9i75IA1AikX4mjtV/7QO58BqNCnABbjC
8ztjhlSfpZzf4dCCf7YMhs2dz1//TFTY+6+aPigqbZHx2rwsxZzSglpCTACQVSGs
tAWw/JuQICENoRq1BBFS/YJf1nxiZr6mOT+OXF+Ukw2rFtM8UHnFg2HE60hwwSyD
w/yBAUmHvksN39mElkkSg2lgYjH+iddvbNCbDTZIkahAJsBdIsiqGAXwtGwA/Ojf
WRXXe6ShfDyHRNwNFxTueXB5scPs70amruRKg7eI0zRNxEjJWHV/SAgDbV3h5F06
ZQuaj0JiPI6iAvjP2uf3TGsR3tvkTQpqiD0KjMW9HnLSqSBWS7Lv/UjybBjUeH3w
AO4LpCHxunpcHpW9rHZtNb1jZKsT7DSKor+bwUnz8cTw3Sb0jUI2ubE0GXOmKQ3e
/kfrLccNozyYPwTQUfMVNDyaR2Qwf411z33zZ8tYYj+jUz1hl7453cznCrI4f/Ot
cpw6EWxEhdItS1saC3MdpYWc4Jk4aU5Rv1VKHVeYgkY9Q5mIwaa7T2Q3hIOuWNVI
b4pV5j4yF0MIeTLly3DLaT7wK+djL14LWLTaoJf7tAQJlK+NivPUsbo6FnwKtaGo
Q05kOORmAEXX9n9HpkPW1P2dUxq+bTTrmu3rSNbU+DMlrFDeNgG2VbyOzEr8AbjX
5KXzNJYkXbSIKhTzO2X58lKANG3tXYeQhHxGNbyOMvGxew6c1nCnGUWBjf+DZa8i
8Em1vonmNRDMTgJ+/8eh+D1f5pr51fsj/hbIV6jx0ao4WolyvdmUllb8ozIoiI++
WWy4edIy+iGwR7FcRLEAYY0OAxNdoTF7WGSxkGt2fBYxNKkew2BhDROrmLeasd8n
zynJA3uzhU7Eua1w8VGiB9TkCXIiTFAqSRyKYoN0dsoArIm0w8qHPWynpEjLFuXN
wbIlzln2JzhZIkhWF6mDraQU49VEfdxtarh3P2pCg4c58YtKShpO5hNkHb5oVHCa
TfKbdQzxAI+fM0lzxDmdInws8G6Lgr/mDjwefezpbPiYERdYYUOnS6FH5cBBvYnG
guXgNNpU3ULLG2eqcjFDLCMzsGj/8cEz+1JOVCAtBomKV7/OR14nxgyqy4mKPo6x
PEZVBcxWiVqX7Gb3AnEHzoCYJkhsM8m23amECs/WwM+zCzifsYMswkuHlwTxY/kL
WamNPeE56UFutLDJU8di9K3/xeQSrK5lVggm5bugCOAtqTNK1EanufItopVOdrjJ
LG44cAtbZ/ciFl7f91YM80xCkx+Ev+gumSS/6wuR2q9c/kUKOZgFAupHPH0yCMRR
VWGVfb+LaaZ7FBHVaRNjjsRGjAg5qwASKUQlYIkvFtaJ+ysb2IGVCbmfwFMth8k3
ZOyYZJd72CaOnrEbvSxN+7ClC0aTH4XnXxlkOEJX0QDDBp+FfnAZLyUYd+pdVt8x
rpgzmgC9E5GrjI7Fzy00eKVIMaiTPa5mmxfSKCTcf2sMOiUn3F865EErF4lNR+Rq
XfOcskSihJROU58QQKy8Or3D7kiG5U+YL+CkCY+ZNS0DxL54F84hYE+tPRlWap45
WvOyMRC2H4jyWtPGx1PDiUzGPesT3MpfvBES6iagfcaQnoK2xVloyrKoNX2x+Yet
V3YlaMOPP65sdwW4ttW2qju7lvKPyElBTPMJkPZmD6eaCwrYccJ984dgGJ1FlSue
ephdDKEekgLi3oJ8/eN/fdkurOZ/XIPEapzIUsSGRk6os8RxoS+dHsB2yEYe+0lY
jdX/zY41Baf0zmetdpw6WMBVtV3Nl5ttmRPznPkbZAWR2I9xFH5MVB/DPxu+j3MB
cewncGriImn+FIHmNMZ78d8buq94tyve0p4Mv2NKAVh1NbCzmTwBdW5Ws22WBUSI
yHtiGIe+Npg6JL4scYqfnnIMBwKxCsyqHV2dxu8QW04Xxp/T8m+jqaAc+DxY3wfW
nJ0Q6JEFiim6uvOiXjDH6pipEvhYMgY51z9OReRnXmbzANdRrWPRf/95c/GTy5I5
rboafYQGU11dY7rizlWA0VC8ZatRX44vq+MNY8g3K+9yRAoW37vQQM8H9FtXNRY7
AprWIlOPByDEJJ2fXgRWcM5Z+8JuNo2XLBEByCarB2Oop5x7piz6j+6/OUCJZjQV
K2Fx5XyMOOWea9YWVKfhxvItfhTP1noV5pXLADEolwRm3JJNPKaeeC01Fr7Jg5rn
BTqjxF5I+Y7281sp1V1vxMgKSc2hW3ZrQH/z/A7+rx6ykmtIpkJIHap7KC4HEJHV
zu+qHtZ/fpe8r24bet1ksAWkQVNH/xDxWOnljOmxLI4oDfbz/1dB/xCDmLF/hLtc
KTSxOEWxe7vfCqn27eMLLDfIf+5jqEIHbO2yUxqCzbQWZbHjY0ueZKBoI+F1Cmm6
zOrHNCmS2EPQhhiNAif/xt4T8YCMrZUixNtvbA5dWucaHk0U/nN/1h8kUCeF89eb
4Ds6aBxWDADMLCwYuGdFcr3ocGB+stq7d0b2VxK1EMUzAX61PTP/vwrOD9kNluYi
rLPZhDvVziCR8yRDl5FKKanv798TEJrp3Z1jHi8lEaL4CQFDC52a4Lj4opnP7KnT
otuXi2XrVCXKj6/HW4hhDiKTK/CRNUVmWKQa65kV7ZHSWnFxZT7EHYFgauW+HTBs
U4fQUlOI3Q+CR8r8llMgo8dWXr3OzfswpUqMxal67KZmDGk5VNm+4n5/22ikcpHv
sO00S0GHqNPdtgxrZi1GS/Z0na62rXVDX9jxubVYgiDIkNJ+XLg0X32TTeXDJG/m
sp3x1COlSM40euFTQ2jyhgO7BM0iMZczKZhcOfama43b5Nkeuy9H6mrmiME5arrv
GXYXKaGEH4REckLzl5uR3fI2wOHsLfH2UhpnBX9gvrRKl8fxQ09TBZQJeyllwyv6
y8pHW3dAhFQWb6z3lqQe8BbI2IdSzSwAuKmASOp0fzG8ypvIKdNds6nwltNBSOUC
yVGMAbgXNBVFofJNwXZzuz1WrPzBfqTaggKlFgu/nvaqV+Yfjb0DsGMDCStaPxXG
EE1VlEQkGfSrZHyg3LdclxhIoc1wHCti8XkWvKEEQqBtjC/iLv9OVrA5+uFz9Tub
gRKLpW1pWc3Z9viMOiIXipHjM6b9sdZj4lzUi6iqXqoRbebClBJ5hEJwK9yrk69/
5BMtxjFrs2UrS1TCeC/TAoHvmLhGSHzpebqwzjwGzrd9vDRcUePsN+qZirIX7Igy
MvElhBMVF25k+gg5dsF2D06n/Peg1nGY/WCjd8myDMAPIlVJ+20PuKRP6+tgX+rX
SW1UvOZuk8Z7c0xBk31tJvN+ktZExWSkNtl/kFiTLUO5qi21g/VjAqnPP10Y94Zn
afrCK66GtydSKxVJV3wrtTTHaUFO6vwacrYwuaMJcV3CRnPTDL7BcDw6QnMRTDgi
ElBrfYcpE+kgyZ8AASDnAZHHX58766b7ZPy9gxiCiPYMKMfvJWZiYa8cJtgBkt/u
7d9BHHfVgWPs0SKpl9wrmyUzAh6gT17X6NFFQuIewvZmobOJrLk/Kx5/Geq3H5rh
tmHLYi/c+u7tzcrz7bwIKIWwTVunHs6UhpyvjplCqIbWSL/37kKAhUrD/0bmSaDT
GQ/syqxpFEdgYrp+26I1/vuv5Ms0PDVRgNx9Tm3Aif9lKqkX8byyFjbYJCB+zSs7
pj+Ll/zM2rg1y4zBODSzzGktxzMbKovkVjBShR/4Uoq/T2OtqMVYfrYNHMoveTMF
x+IzR6rDY5La1hmdi3l4Etp8Jr2Fsgxk8jzcIV7inNqAeAqqnplbrF4aqT06x/L3
DIFFG0CNLb3iGLw7nl+j0LuAO5eMQRXY+zDv1tPdScuOc4rnJ4rV03NvAQ8XANRZ
Hz8G6dsddXUd5L2V4oDTcemp7NljF8Bk4wHf0ZNuwpUVWiz8x5/aIPqEZb11PhS3
GtcIiEu+/H2K6mA5nectCI3livJ6T9YIibJ4gRA8uqMfbZxedr9Z5+doSWfm/LL4
ye/sC5+KW+FBfsMQ9NGJuGotwJOABTEomzGADUQwbIPzBlXs/emSJ47sLr1O81SM
cAMHDQYdBMaAnVQi1IoD0qhzHlG+Gy+8bL3DK7eIho0wkqdZUK1yHTfokRX3ApaW
km+u25KlkM6HquDPAtumsA2vbiI77I2V/Tkt10LX+MvInpzhkXJSKcw7STMD3nst
uVpOlXoi6IX/uwQj4KAp+A4Le4kKOtMUhQsdwKBfaHrHCA38kx2fLi+fmNw6bHw8
iXQIz8N/AKt4NydGB+FpTlTEojUM869iJinZVIvUna1ISyraa+hzdtDfGBc1Lq6D
USiU+VZtipi7mpHEWU+q4KmTt9NfM1EqVxOKNgBZvaUVu/gB9lYOd4VofamQD1JC
wuRicNM4bGl6Cgmg+UmaZQMBGEZ2cMWJ1EAOftYvbqsunpp+ZwpV+rXmMgVf/3YX
Mh3UkTBtrOY2K+xspNwrt2zMakxTaI2jOkCkdGwZpfW4UK+akZzs527e29aBTBeU
GG3r8pT/1exaERv50puI7weHDTfv0bCAnBh51t3afLcwFp7vZa66esqyhFxafby6
UUHM1Rz9fXJyaKcLnVHd3VVhW10vn/5+a1GXL7mSP8Aiw5xg8ENa09p18RQtdZ23
N7XoFUcutSG9C8gz8rfAClbfJRrJeEzf80Mjbsc72QpyL5sWw2sez7+9y5dT2RCI
KdrIBZlvNu5oscSRpzQ4juiwP8NbxNot6+TebHUmFOcTS9G6gUpcdInCRbU+EeXb
sijjmT6afpJhO2jZmCVur62Y/g3OFlI3hna7LWs8eWKv1eZh4QMy+/8kOFzd6FF/
c4nH/BXk3V/tYHFWPciKdF6dQTSexp/cdmUi4CKZJmsG7woBF/o+j4X04wDwG6Ng
2JuyygRHWzy0tv5Z9OupYRFhQkmtw0fjaD8kdYUut3uQsNpVx1sTwuW9PmZsiGpd
xiOC9MjJBkGpfvgLii/JprbBt35JmBaUbjqETiEKM5wd1JCWmUBHLuTSXX8O1Rfd
+KinC5vght5LKA+moC4brd34XYyKpa0n6tzGW9DnJm4LaDMm3bsFOEDtfgyZ0JDG
fntaurseFdJMAz+5FShJwvx3/MOLA1dvAcwPhQ2p7qqK6QNvEd0rENDmj7lcMMWX
/kPX1J7VbR3sypIPbq0Yt5J7C/ZnLXPDdgIRytvmg91GAkaY7T6HMTB7bLqiLo2g
X1lzODjBnzlUil5j9yH0CBAS0sAdujeSXT83uPSWToKb3lzcI8Qvk5JETFbwEcO0
PX7gNsy3mwII3Gwe1CytUOrwWbG3KCVgEUEELkZBOFZRLQcUb4SJpS12Nz+sKJX7
2MPu9Ovwsm1oNHwCC//G8MNcg5bhvF1bRLDmj3u+1ljX+PTFCb0+j5xnH96qO/jC
dUV0gVXXxdboQUxHQWdy1OXkjeaGl/Se3LLII2w8HFiSSRUZdwNMAsqzGVvuo6jN
/L2tyVqVjQvTbcRGJWclyDYPP/iythNnjjl97sly9dQy3OIuC0vpauv36nF89YB0
ogoTaQ+Sy5lkxR5K2QHB4kfwDNdo8jg9wHXYVVirABJ0HcfmE+57uugGRS7YkVCN
2rWcYn6Z+yX76eWWAtumYbu1vDK2+X2gV5a8Jt4XpiqHGUcFP333Z1lfSQtxthMY
CJv4CJWDwvVILXE/vRvcdOIvVSXRMrA+HZu12s3F4Xqm2WaWUKLg/FxWsL19hCH5
uwTnpb9pp6PdkL8hheK/hwAdKEMbUpuH0BS3w17wJhjQ+7Nf2obJkCXEkoYGHC7o
HssCpOr8xDj5hiitRqSeySXToqr9L1BQLJPhcM+ohMLHvPOLum0f6dTJXOpD+Ftp
9frIjHhX6/bh4+C7m+Ssp1Rt/MD8qqnWRazeeuZj1jJPRpap103BaGsAW3ozVvh9
eYu1ANwkercrGxuondHEAFDWMj8E8Px3h6PhxXMp9WkfjJjzIvHWPDhjVMeBtAIe
AfBJ4pdv1ZoB2ODAboroITprSxmZs9nqOrIz6hvz9Lzgs7PM8KU5/xq+NIe9cBkY
hRkuLIFkVOXSFldvIyVNWRqHZpIkF6jMcUdJy1KAUnxgeQN5Ir1tCxSpxWNdXnOq
j1UCamQ8nMZKSPkO4CiJ/KYjVrNyUw2fD/kGHFZFoMH730Md1+TBcIYA8A7HtI+W
36I0rQxjM3atvq6uNN5hRhMcGrytLMuN+4CjMqeGYu/Jwc6ik8dbefmiWNP3XuGb
xyCzUvKaXUipClljeHKzNoG7we0Ha9z7V51Y977kC29jTZQ9Nz6oOBP/B0UkhBN6
K0cl77rxWPSSaSbrPegNDytl6YUFal+5tEJpPLcTqfhi2oC3+VE49jSAInPVlh/4
VggoUoYwpfzMdlXdxiw0g7e1ulrhErh8hDinAoxnWopQOtsCGYfRe0fOjNHW56AE
gjVvtL49aX4kt6kZwr3oZ0O5XcRJ0R6CGECKVsSCitpCDTO0JUpzM49nxJ3U7LXc
4qeSG/rjF9UUXx2+c/p7LBHTHvb4GGErmeAibNFPtcH8OXeNFcGo2PJWAS2vl/zv
BdcQ1YxLFiJt8k5ddEHrczoQ+WGmaAhLif7vuL7vyj4Yj6tyRk3xsqPE3rNl0rjo
5gkDHTPCcWYVATy1QdI7GVFMiNsWi5wvvV7trtqB0B7yNvI2xQ5surC/yieb1fd6
k+zcn09YErhv8fn3ggn+1RjP1NsI5UPt3To11iC3IXq6n3Z9yUMG6m1gMw4ViIJa
qcqnFlyMntJ0fhIJZAh0CO3wqapQy31o+MH9pb3zUw8bJQ04jkFfCIs5HD5aKLrv
iYUiZJ11H5SxbsrSF0yziSiiJpjfTT1z/NtLcyMQN8GIoJ1z9sDmtJf4HpRHfzez
Bb0Yyt5n8vjLgt1c1L8PgB/Lu16IllLz3Gx2qxOI/rjLdAgvHyQns8XwSHKijzKa
gsPbsSBRVv2o/Uj0gd5CdAICNsgP7wy8t3t8vAujevjgvsl/5KewiXzjPKy2QFJW
hj2j1wtOw7Dz8/Xezq8rEnFUaL3ZZeFiKwrSubCWzlmZUsn2JoHvyCTMNfGFXw/A
3pr+Au5QvSHSoDm7mGB6WfrIXx8ToY60APmSCHulwIxMCXRvJe4FlVa3IsvSHqeu
qhyplpx2NBQBY7gHUVh7I0bX7v18UWK4NGVMHq2dDkaX9VPhBHjkdqDpYiq+d3sD
q+2RoCzy1xweZe3G6zals2YvEhBunU82VMAAc5sASMY42gyeiXRlrF9DE9PZ1O41
YuhN3ub3x8cMdZRDYf88F+d0BIwbjmJ1yBX0RDSafEZS36dkeR8aOx8QNzwFlUY+
GfCpzg/0Sly1DbIsswvA2UNRAq8U6cDWCXg6GLwiS/hm4LpgVobk7Mzwh2mFoYBG
8BRYPRLpvUY4YcVgs/7q/l2AaoPIOTr5Q6ucrOdOUHtck0arS6clHfbKtyYDhniU
l5HcWZ0uGx2MFphgZjWOv2RpCLaqcA09JkwTTA8AL3PvWqpsbHKkNKf0RN/9uMzK
JnjSm37O/97JYhwkoY4plo+QPzFHYv9BIJFg2GEwXqoRPJUblb5RIgJXmNxbDfkS
iZJeZmCo44NCJ4pfgYpDZlLJWkuzxD/47/0tbN/GIjneGDyq2F3pIpZOIUssX9Sf
l4w/4u92JvexpVoQaISSGFh+23xkWSWzy3ppG1Y1vvtNNaBSyE4uV/6RZ+93vJuT
SHerto82ZMADBYO7hhaEBVSrNIN7/kyiw7msypuyWmohMwiBAnxUlJFR2ZBLoCmc
6g4PKzurxT74V2yKEOxbMe3cZzlQulnRYO8ek+LtJT65BPTavY4L9IEAnEUeIaxs
IpCp4B6KGoAtiYyox08wo0xTG32l5ZjhqlkU8g/Cw0h5cC3IDa4RAMQSJ2XTlmhf
tTqDQvgMxtUeiCPcmnfsZ/3NqT/CKlCU4oX+zE5WjZ+MzIPvaQbBYC/GV4zGlUUu
7TdWaDD2v43dJKOHqyC3p5Dh1gUB2gS4iQtY7mpEX7UyTpw4UdTopuKDXuUovKY9
l8pHiJPNua0bHH36SR5ZlJtLcVwv6pd0ujH31kOhZ3/PQsugu+4LaTlbKBCS9sDP
lM2zB/Vch35FXxIDipb/KfWt9Oz1kQ8I3htHCbtr6Cmc0SgPcdnJVkX2yh4ceMTz
jMR6ltql6oc3muLN3Dq6ntICn4pnzbfcP+C1+XGuia1LPXrHfq6097sKUdnkJ4Q5
4HQwrHA9Abeo4CSVc3TQQ8iHyjJKl/LbYpc4sQf80SYpjZAgkds5opY6fX5icm0D
EcaoiAtb9tdhk/wpebvTV2mM6be0EZ5Tz325ZDIom2NY6zoD1DULT8dg15lZcpaB
W+55N4DXnJwLvZMjc74h3H55hCNo/PekK6x1FdpU8WxjfmQZXbPrfixxtB0U1EGR
UyXj6vA408qWLs+coiCvmInHiMRWVTLia9/quRnHXmvb5iZlK1+9hLHnYg9ipy/b
2Yc+Fjkdm3Ws+6V2z4YlFeEWVHSHr5nZjFtEDwomKu5aWOGpL38z9jJs3eA+p5Xv
Kz1ydjpfT55bf7v6DfCy4zit5I2h3Ost9CTC1D7d6rFCq5pxGwxJi/eFJrMtmr1o
9c+3OSesvmsuCJ7pUpwS21ps7hYojLEKqKwmBfGkXaIyM8bJSxyiXvqichpLLgEq
kEVHsRuvV+AfJvv5zRqrW3U6x8joYwFnusMepDcoKNh6v4m9pd11x1nQ7nFkATCm
NZA0TJU6VXGNzA55KaM+Wib1TFwg2S9lO4+OP5VHywb73e7ulz59uQb4wQwlWGMd
fl0R+s/ISJvrwBsuuNdIrqkcAzZsB/Da75/hgKiVfS62DwISJG2UBf4J1ybjMep0
QdACcmTX9Nusv0TBzgCNMoj6FqWW+ljHPyT0sLwC5+qnyFnobpGnjAnfQDg4+BhY
mrKDVBhG72o5fXa14l/bMXD/vM3fWgBNXvd7lISmcQ+RYifF/vbs0b1zHS6jXyxh
mhhWdhPpDPey4fNP9GuB6c8cCOufSvzZqhi95VNLhZMy4Eh/J5Bf9r+lCjLpHKDv
Zs/omMLO0VKzsn7Dyg94/O+QKb59ew4cDW5LRRPQ2HGxHwmaHcrH0Ym4qqHUfMta
Z1q0kTlExTpPKpmciOLrAff6CsrV4FPKjB99CgEfBEUh1SMSDsqgUmTNvNNy6oxw
c/4D4WN+eoDpq/Y+GA+71HHLnA74sWbCN3C8o9QjKpyC9WE5yTvrcoIncsYBkJpq
YRCp+Q+LnydkLr+JBcR0ZoazBwRGlM1XPSzv7fQyBH8dw7FbGCvHIvFZSlZUGoep
2FU+B8CZONKiNf2xF6IglPmI7hVnH+t1JtVpO5Me35XQlSZLI9DouKqBCngXcfea
TewsIAQyGJL1f+XQkTVn1BIAgNSmurZuYvI1mFK9glRZ7+KFP0AEGHkx/kNTH1d/
XOz09XnjIWyZYsJqp4zsHehiIAh0zqwdPP04sRNGlMJWwzWHGniBsL87g58rUH13
QZSv2tAAnQyKFRr6R49U8A9skQ5X+DQQfq3wz9ZcRp5Z02rC5UHGzo4f5gIEuEth
xamkPPoaH+nO6wG/vpBcNE5NTOq1zEmY/V+5p/99WKWdcKRXS0WO4YDwClNFWSMR
zXAPKwkg8egTmFyvdhtGdA43dvNQLJoeEc8iQiEvP7omRDY6DBt/SPqDlWzIWdkg
pxghhkIAERAmuzBS8lvEDR5fjbNT2nozenVWJAlTpskV38sq9a5qqtilbUqp6ewi
EXUwky3XppyDCqQya+hMgye+4WA238u5yJF61wBCtYgXA4L0E97a5KhMujMWOSTs
AQT0cgWzD6cxRVQyYqrLaIJM9t7aQpXQzC0BWoUyTEuOQi09ZDxYWeU82mYDT4L0
61lBJDY8eRRYzK1f7liUSAa+F2BfQvy15oUqCQaeb/t9xZDa2kdUgTafnXEQ/cLF
t4RHTOi6dlPIncdntkm70C8BuL7bGjBBVDsEw5NJ2l9QT8s6FcD3HhjF0HcDJVjE
o16K0hDuaCGO7yH5RNkdYq9VkRcaOJH05vPenwn2qeVklIVlDwCzBrxLn/7021Bf
7Lu7MNIHsaGAJCx6LyCePcp4NKtY9OURFa8cCFBQ6eaVFMo09wYcy7/rjoraPlhM
6B52AWJVrKKM0AFSI5T53RdhbwcyJEuhfhMYrqxKnHo6ojwF4wg1rhr2WsraqL9a
1sRD/PX/py+/34SFPaI4jU8P4rR2uFa8ygltaSRkS5DiT4ztEgqQtbUQdwKuUIzF
YwwwRTVoUEiIBjZUyXc3ZfPk5+EuPoJCCrikIO74VEpwRX33dIXHorDa3tRcGgfV
d1pjQLLdu4CoHB9SMhllX40k5FkDPyrbz9md/uSWC+gDuvldj6nri8yBdd8ZxomL
VsYl7dCu58JYDuXz9HnMFEDwgqq1cQGPK9rHIamVy2Vw08slECdIq4+wNYrU3UNg
2+d7EAHIunLhMlBPTjLdff9arYUWYdlywW+mO9taUXTCpGW+/sGsKuYHMrb9d0Ww
rB9pq+bD4P8zUkb0XuUKChqyxPhLhz1E+DFUSU9aJ5V7sqn5UVVFBE6dQteyzvqH
dItLG0FewmvdwO+RFriOlFr6RHyP9TWrv+rbaKbFOR1tt27i9pSnosLZ/ye19UKf
mvpHcVMj0pIQTIb9uQKq9ezKmo8apGaLRs9DvTEdk1ntPGuhUJVxSl8sBIryystT
r4JPunRT/l+aIAtlQgK3IbBQC7UCkaG51lkRg0zKphCHLPVD8slCVHlWZYA60ENq
1rF+e5BlzQ90sghWM0QvUZz7nruhgGkGdk8ZXDgl+Y7IbILTUFTjw159y2UVRORo
5CM1Vn6U3X1NqmLE2hJuOn08snlh24ohmdPV7JwBgQGVhuwAZVaX4Djkuoe5QcfO
LCcSMUA50qNMnjzGBBib0m30gBtrV4nFYgO2a3QIGGdb+hPUc8ArPmulaBzLyZlC
bjcruaivNrNy6+jxcB9Ej/LUjiDGIwR9oxmvTS6HtK+cRoLkvQXG2kQJRkpHNby0
uYUn/1KYf1vq/yYXCH4Mw077GK9mbiiCj0ovCWpUCCNi56p7qv8whLujwYkbMUsk
2V7hewV5TSazAu8qt+tnBwY1wLOcLltYhdLBQAM2DIeiPHo+HIye3sDRxEVhV59r
OiYHF5s0uU48oj/JTIKtIEuw1qQnsT3odb5uDSMDZ5vjgUqdELYUEEyN8WaJAJ5O
dH+zcR1JTyhJw3FnEqEqn/KUnftUm39faID9iymaqBJiteAfRP/aJLCIOCEQmSgE
uq5sEmDPhJv17/ETsR9L3LOxIHo7bV6fj4V8PAMLj6Lc1w5NGzGPT3ws6GVDO/Bg
Ja1yQNYGSNOaaN40IYgMXfC89c+9kEk6aNScx9taU8QqE4DUuMla8F8WJL/jIdln
9YK/pl93ku54ZaeHwO/+7/OPyrDc4hZdzfLZeK2tnsN0yfeoppHqc9lpnUnUzpTP
22kvyk4Z9lOEPidH16tQK+wR4q8dPeP3/MTRWvMyQF437KKHQbgzk5HKXmq5NsL8
a+jT/gzdPoS9v4Q7tkF5itvf35Y7r5Rg3JUo+3++nq5AwoA7Z6aOSMsxxfLMjdxa
U4md79gMinNulCHa5Bb+Lo8dxbNjSGKXqxID+gTPQJbg5v3IBp8NG1J1lVXKo6QX
N6/hKg1iLK7g16Aq+MQ2rJi0SExKW0GbgETckSNCU10Vkr1BS/rwjNqsRf+K0wBG
gbunzfzGB8mpaVvXKACN/xnzbtg1QaIxxUleySEtmPYAf4pxUz71UhAlAvGC/yqP
/4oPwl9p6pgWzBrhLqJ+AeYYyaIkbpES4gx9Jj4RVMoL1x+Ha566xmdMZDt5aiKo
1gh4H/6i7dBHhDSBS/m3K84U46pbMq+2d+Ube3tJmnP9C7cJYZP9w8KIE6xFUVcg
Hkr1W3HcqqOkRrncYUR18yE12k+x1yXutAhTTTtliJV4V/uY9gWoRFMUFBlnvNyl
jDROAmG7JPmKW8q2u0LDfCZD0l5GKKVW5BxbR/vMDb2aRblI91CjRUK9E/OAty8S
fpJxLiDzAdUjP4H2CSUXmDjWTOUNzNWqz2rx78/knyZ2pxORjo25zfQPT83cQ6LB
C3dkSBaA0hhr/rXAR+E1Dpf1BsWTjWd5rhJik44Dkw1gPRdqe3ZP5o1UZ0RBi0yK
FB5GY0+bO2XH23x9OFwIkL4KbvxtxEP45pe7DMB5jbFVpnUx63WhZbburYW6OIBp
/Dlg5pT8ropjPfeLGeCXvuPOmsx11zZhvje5hbgq3+j1nJ1KttNtDsWVq1xRTy2A
0JxnLTFDjlbWto7Ge7jxQqvbeBDr1ZZJHJidfD97Hn/mx8N3a3MrQbos+qCcFJJd
pAGlB7shuqtPLUDO7CDMrPKncOOvgrnYrUOUR1v8EvapmWxQ6AvhQE159hgbfqXL
X02KloVWOjTSFEGMHFonDTJpFYbFJXSKUr7cj0SQ+KQ6PxEJywthm6Im1ChidS9l
Hyc8uyFKTCAZnWVpvHl/OSgwpxDhAXc2PcIJbz3Cw9tsPbfWx34B5AR5CC3Zk0hM
WbN7pYibiuBZwYnS8mItIAnQQM1/CCY94yyABMk2JRew4XvwxRostMqjhsTeem+j
RFjX9LOPo2iRM7IaQK95/NyJ7PK4SCovos1hmO+FSv8sBx74p4t6UBzLlCqTB2R8
sBmczu3gl/exU7EEP3jZ7M+gZD+KO4NbaEMZF08b6/VQ7cyi9YYpLQ7YXpZg2Duk
0hkde9DgDGOosvLhcjvnLrwGcGf9wdNQqZVmMz8lI8x0gfvt6Pre2LQv3cnPmD5c
sRtZzqb+MnXZn0dM/fLBLhr2aq9lqrWtr4KteELl5z1G/cHWrqY9gtbvCt+/3yDc
mRYiayYcOzUpWIg0IatDiFFtvwtSdU85y5P+JsvdM2Hsef++rDiqLuHw7TobOv1U
a3gLiIk3gT6Hu0Uw/PHRDeP9hgpG2AZE25Dm5vZ4hfn+4DwqJA33PFfCoONPrVVd
0idFPrMMrKHODOztuKp95ALmO4nxjsEthOfZNvDnkZZLbsVeZ/gqalLZapBglAsY
dv9kOrRsH8xIvb2fMiZGYpLtO4QtzTZXRffi1txikXcAygfXbhkhKpJGK6Zp66hy
AmBMggCMq3URc/n18/e2BdRSihiaYeafT2RtTXfQ+7S9xV9IjdarlT6vmtiFHMJ2
qc1oyR3x+aavq6e4UapaeGUT/y6OfuSpWwybcCtkL1tom8laI68HyYwr1DnSG+Ux
YHR2zMtDtxFO0BGGVADBjqgIneRtNvlLHGwap0fEWdML7G3hc3ONN2MVXlp/n70O
KSW2eCj26N2n5HqZk8BKXFMEXtdnVnOK027Yj522ntXcBYM3pnx/ik/AKWU1to8w
vVHBgpPUT2COsY4+KvIPheHMMO3wvubEGOwUdqmJEQVlZsGby3O22KcmcEaLsBRA
QtsRRrBgjobwzaNPgdWz9nm1PLdts4h5TDmLeATYeMcRHOyRxB+LYzucXw520eq/
LQwg3RvCGPiqwtoCec2RotYB0K+8OT+89b7npZtaYIe8Fq9TsETq6UmIKEkPIGGk
JusjuXYddNdix2LOYqRm9y2P8oUUyjbBAIkoNdoWk/mW1yGVbixhaKjqKTppgzK1
tmIgrDl/MgsUif1QwZSBjIAKhdl/DMoYh0kYYrEFAyWlw3wCZ2iWI8Fnc3Jn3nLa
5c3TAVw8V3N5vXAfdL7Qya4sggCWfAU0jrxY1XsBCqg9KkPrXG3ToFLtLxOLPMP/
TdEoQnsJ+KCPNpdOyY/NUa2/9IFRtcVMLtI20DToP1nW+FqV7trl1HNPuLAFoskl
J2Vu6oHusmA1+oXlqWYAqXLacMIlX6EONCa6fS28SenNUQUkzyrVr52tp3vdL5sB
5qKMHTHYYB7orEgWPMFEPegJwpIdiSebTHdYPTCYYXVmvQBPsDrb1oI0c24GLZ7L
ZBdlEvtF130hst0n4EuxpU52O/CtbcHS5bJvcr42VkMGzFbsqBvxsSmLOjZFRcov
gHPInwUc2iVDBiYxd2uNYhscc1UZIpjJDOj4ZQP6LBeq5G+vpNIq7bqeS7VbOlum
hiOVq4CfrPZ/wM8p2n6zJK6N8nlSZG9atjgt2FmveO5YPUvmfndNsMX8HkknOIjG
X1bLKxRWSEZIuVivHkeLOhQR2T+3bJFsTC6/9wmWJoVqk8wnU2LW9DT2bnhucoS8
EwF6xLLpfTv0jIWH71WpixfrVR3BXNGxEW4DHDI7PzF0HIb/OaiVzA1KriDfi2r/
b3Zx3WBNcwz5/Pd8PSmOSKQ/0mHRp09ZVplnM4W83EfEMKnFycSkqxn6NP9U/l+f
YLC2X6qddA1ZqQoDE9Ig6cMgaERnsvx1MliFu27KwTBDVgA2uS1MxETidbdRXSk8
SBzPuBuj04aiiceJe0Vksyuq19YmT7gzTR2qHw50dH/ysAMsrk6vkQkoTLHLI8VH
C6WOll2E3HS7Jamo9u/QJvN/J12ObbwLjGrDaUK+jx4DQWMtShQjUNULqMXWNTOQ
X8Izk5LHxc1mWDXYuSGE8Twykg61HFryUBl7qoCssXQNYdOdz1PdgjzgXAiW/PK6
V02rYV4jhTMSp4WgpGq2GUoJzdtYwOLceIkCk0yuZf5hQmYK9B/XJKNnziOEPmRH
7ILkzNjKSJGkpDeFeNwffAlXlSDWGBb4rlYbMBNT9Wk4R/rPa4D1Z8mj6PVa52nk
+U1fAPkL73+AOtNMxza4lK5y52sPeTjzPql0MMjdNJ4Fj3jJ94W2PL4nIEIgugnA
o3JirUydhsonzO0KpAsMHgAUtdM3IDjsv5s4Bu2td3gONlR7qVE455QLpmUBQpkQ
OO645dfggqVltESSrL0CIPwGRs4tiPnaK8sRBMb7kyXA5HbaxpoD4tUnQxTf6Ze7
6XmjWerwaQbrDIz+fxBsh8ari9MKMN1+sGQiMyPnE/30dnJ2NwV7wiB0ARsR09+K
4JxQoGC+sKXJw8RUY2Az99t70xBcEuD3/CdRycRcrFhYo5cIdUN5/RAj+xHf3AEq
SUeuk4pl7aUmhMITzMWJvLi/tYpmCz+VmYfXNE1FHOkGYGl5ypK8jtKzWfY5S45x
JwAQxBjlxOTg9PWz0su+LbuepK0FtNE24fiRiS6fnOImZQngI1qA/ny61q7pbQs5
4a97yM01cnMioaf0Ibseeh6MP1hGaXNZXmNQRtszZu1xiHiUbyRAJSA8dVLoDn04
Vbv7bpulA72QbEF3xEVwVrUxx9yKXwg8CM4N9bN2TgC2gh4lpynpHziKqWazlMN1
snL0JJ/SjoTyLwA60+PlpQULgBMqfYX+zmoRwcyjiJJ9V6VsOwZsqeQOeNcOSWdT
o4dZxckJGnoYKp6WcFszElWUpAYrZRY/XqtqM9M7tzCIxJU19A+geZ8Ox1BmEa+e
Y4rddGlTeESFiHk5f44+RZUdY8jkiSMReIzBT384n1bmgn230NTIBE2f72E1p0l0
5A4ldqla8YdIYNLbjIuML0czf2CNmB2hA8ccp9I0N0rlFgbRytGqo0QsnwDWI2vQ
tV/yTWzEMlak6Ovx5KOWMgRd+b5XZfmfH8q1B2c95rP46kHCJBAmVTlUNft2ZAxr
ZrgwCBDJKNtXyLXGhqLQB+SgsIA6o7TY5lIT6Dwv9+GXjJ97HtHNeW5tMZa3U22d
YN18DitDsi6DyRFM5SScRaI4Sy/Tf7X9db8JVnwBMVMfeHy1QnKcwPKf+48Is3sy
A2pHykwvwbvb9f02YuUvd5AxhYUthsdxFbRUhLBjNIjXFKWxchWvFBpjEm0Cbip4
YPzyuSrshPjQdNsBjfWSMin+QGt/qPBYN4D6BC9OddAMfkIvnG8BaCceWjaT0NSD
2RRiR0+rQn2LZBfRpOTqSe6WVsqx2aysSJv6E4GOXpIuik6rU9L3PRQh/0TLlaUU
J7ZNYhxv1rFAqsBcZmbO4/M81NmPV/VPcDDTO1/FkjKfPVj2vtrbWa2N2Qw13jkS
JZ/VwtK/WJ89tRGreR5jm4N3UG1oQk9gz2hVe+c8P4XQ4HWThfayasTxVjOU3VD3
RuucqRMM8oqmiE8lZ9s7e5zx+Zt9DmmjCkvqxg2D1ixbYhIVchOrRl5JSVZp2UpG
5EHfrged1WXfJAbLvA0Q3MKYUV0m2eaA+dz2tBZ1LgPuEHrxiAM4+/6giZ38NTNf
0zyDPT5wHYPQ1wBP0p1JdVJzj+OC0h95TlVsaDI2dg9MruR2ZgGfYNz+on3EiuWB
QEANEvgezIEiDBEru69+/2xlP6w3h0p0CH2jQSPK6Fx5sL/aLZuwcUZ/+UUsspXR
kT8suo2kA78Y7TJAi1QWlz025mgX3+Exy2K4HAu9JjrldHQT3XguIkmnEi5GuFgz
5H/QTOJT29vsykJByHq1Z2R6zr50dzl4lKDZ+YmTsNZk6as7oUVGPcrjNYykdn6Y
YIspR9mivsZ02TtRNlaoVuvdEso2uGlxfRUcZxpvEEob3HOQz0HgoakiFy+71XQP
jTSRmDtOcD05S3SbReKllcvcHLh/7MxtqKUgj9gB7wKiZjWt/Nn6+uDANOxTAhDc
HhVhuS1xUxskZ38CvgxZle3U6+ip4xyM7y/BGCbn2vMmh2Jhi669U7FVZvEizHhy
jjUm3SCqGx8jMTi8+wZ5qaHPva+cYbg3R2nbAxG5pNEz7GJLI1PMjOCaqDRNlqg0
oegJE2ZHoydStk/8qwcXL5fv0JL/aEVuKnnV6Pp0bNkEAK9r7npDIb7JgSL7mRPn
kdo9iJrVv2+Ex8QE49LObjEqkRRNUJAxNRzUWUoqQU/Yaar3B+2CviTo6cAGeTDM
DCmIy+sFh1jZa7zxcxAaF0zNibF8i6rUFJGVDnmBu4QZ79SPTK9GjixDQMVSKwv2
JBN04HvC8ZRkdAEKf+d4Nqib5fV1aFUNvsqLoT50EEJ1hc5UlVxesZut413KshEo
+o4cHNVL4+C3U4DUOVw/KsiabZxWCKvjNR9JfZeH9PORBjMZWeejDt/321R5xzSw
PYorODCoF17Ivfo9oJjShTdbyl/TEZ2YzmvkmZ6dqzlA6fhzY5vvrE/usH9K36Aa
diomY9RFFpn1L5NNRLBf8iQFJP9+bu+CWBUOfpaG28EnJjHS2SlwqcRzOuUmhPzz
Y5Mz8rXFWE2widNIeHvBOzlyovWRwaJsy52OCy7AdaBJH+4vjJIoXgWOy9oHAQfr
MeAgSMXa0uaI9gkkAWa4AB3l9qpxQ1byzEVKxfKo2jT463rfzcHWICTxTjEzXDZU
OdO8+3NAPISKKKxM1hcjvwPOYJc1tu3S6e9l2AuOb3eCVKyftFt8DPkrnhyxxuAK
jCgPSTb765dpIOP+BAnIzlaSHyGznY+eIaE1+mUF/KFZcuIYiyCJ4MZ/7JhDbcc5
XPpjVmS1KE0vBDo6aYIMNgQBynhilzJ5hJ59VF+DyK10cyPGus6evQThdhM/Qgvu
rztJ/xfjb4tWJdu2fF+zk5W53UCG/iXYRdQXxmF9dkwRiEwcQN2SvgxBYvKGSFxL
uzl6Jm0Tx4eV73pO0m7rhlVoEhtqubcFILJfE6oRJqzUfXlLlc6Im2TKGpndGAg9
wYpL/5G2i2BkPtcXwtADB2i9PPVXMjJK8eOap9nwmxwOwBR/CAckhBtGsu5s7V2T
/YpjXnTqFqvgwJIq0GMwvS8INxX9av56lE7iYzD3W+lkzAHXkPg05ExJ47Jcl+Eg
svKVcqxadjPpPjq2SSfH/8+pFLH3Qo/Ajj/3bpd7HTP2KVburICxCqnXuD83p2HS
EvmagpcfUPuIy4gzXObfx+hAwSH9C5IzulryTtSwE0h3fBAGzuUNKkfan2HeJaA/
avE+H7vb9VWl9Qnf5khb4lVCg9aE0IdQJD7LncKXjOHqdLI/NArewZM+/Ll4+0fJ
sAbTW6mhttPtCCw3PkPwB8UDLyK1xL/yAh+vYyMhH859iIc4FOjxFpbvn36ydgmi
AqnkMaPB2QwXFQszwbReireZMiYU2QByUr5cB99GJ5nJTQPxA5LbWNyaFC4xg1UE
BYizRwIlanvdHgsaVEm+RfCXLRrktNjXdHgAd+o6QfFaVNyOpHhxg851yfU7u6AY
4NiSD6vSE/Y5Tiqjli5bpNjeo7zsJT5sfX43bmljl/mSeFyUtcTXihMaOm3z5vSZ
w8VcxBUzMeWPj3yMxUeGAJ1aWDKF96xSc2/mXSOU5+ig4IbXA7psi89Aspp1cbqH
6deljerDHi/0FjU2HOhkgER10RRdtgEK3SiC6r/dsbdbMSH76Iv2Fc36QnlI0TPn
qOGXFy3BdaIgsg7x9uWIwVLeiAZDMYWyyq4BAs2rVV/DbdTvefehStW59mi1xDxZ
j5t73I1xXcCqMDMctbMz1pZW1g/36o/itlboG4xba6G7O5zJB7HLhmaEoKcdhi6V
GBG0EGZFydxp1kTNmpTyi3RtoHtOR4k8VhuLYmsJFrYg2dRiTWs8+GAniNCNFwcN
/4O5k2awNvNjvpL8rBNaJ1utDz0n4JjXNNd6YATh0jfefLhdlt+wGmo2/ZtnH45/
i0I9P9Az+Sv/T7k5uOwEv2DzMOZC1IeWh0tOBaP0qzSqZbX5pbcnbWbRrJAlg60F
runD4oM1sYOX0BiRZcwIFH7qhWLr64UN9Yo0UjHqu1ihWJzoApiEKt+Sj/05brWw
sXNHsw2WTb7Zyj7Di71XtMzNymDlinD1fdeHGnhYMmLT7nStQgqXrG0cBvKOR454
HZkOhzucki+eZUnOtuSjuHQ0Wfz7qmQuNTE0pybbiIwVlFMJNLjLLVm38Fpqg4qf
fdC3qsPp4VDDLzoQ+Nq8A05yTYaAtxFhmbetVloNqA6LOZBHcZs5vGxLoUlkx8Co
SB5DHcsbxGjWqFsARVaNVzvStluJZ1au9MNP9aAU2QUFnHnlpmjz45WIV8izqpUG
VwFLBvN+ouiIQ1fGoTiXmOzA+ftWG8OwUsMehV9PmdRNOeyd87KDFmua3oI054XL
KPmglf5c9HzwC2fm2qGmWk8MsDwfaJ6HrgT8e65iwFXHatn6xtIdVtPJoqkCirB4
hVN2d+PKFm2eSDlY6gN8Jzx3Z/MrHO6wCJL+lfO+jJzOvnwfRYz3+ZAWh92t5d/K
CZLa6fgS8bBG4Jf4skitB94Ch5BCk+zj0Um0m/Q4gdA3GhMl2LYjSPYciq8LdVSf
hXlNuop+ExNAVnjwBuD+wQK2DHvA17Bgj7+EMHx3q+4dSDHBhdWRSYiaPFtU+m0W
g9r9X+xRZOAV4W/YVcCw/g1hLIJQzkllFftGAaJYZkCQgASW8Htli3ynx8U2tZVN
8fJAgEzHvQvouvUHMlRlYz9V1EpWrs72gCytJp7FD+TAaV+31I5AKpFZQZwTyNGg
RLqcfm+VzQ3ii7/5SXTHLPT+5qaQyCYJpvVaeYKKDmawgoEaCeTRaIGHa/qDBQFZ
lhrVupLCm7DAUhp1uhCb5cSYCF8u83k9qI2ylO6XSCIGqujnKOfDf+bMI4GmxAgU
PPipTxqDVSSYW8ti+aasayJo/Rh11NiYtMcGlKpKSrDK8VkrkvWownBvbxlEmjfb
DlM6dBH4iWwSVwlgN9AD8lJWn5taARFaXq66G53mcvEuj2ynjLW74dbECKiyb/ux
lXjc2uYtEZZ4wFtLleFBjHbcJOW+leZ+J+zJwY62FQ+JHQIlxGLxZP5hN/DhAvn9
hHFsuhaVhlknFzKQL6XsLK3KDtlMT20t9I0qWAX1Al4Xq2e94lv48PQ/BmIbSRVq
ogIsHF7CFLHggV3sXjUiNM0wzn/PeiNjIp2bYqDAilEfmz/8VIoZgEvsORCxDc2l
WHADoNoFKTEL4DqYKW4/owRbbBiBI9ToBjVl+9Zae9CVRLJXt8XggNozdQConx/X
ZRjzazf9/kOQFSiAFsI8tNrCk+p1N6RLLURzkUVydA0HO68RJzBsoYjylEIMOy9n
cw/SXOrgNnDo/DmXiN6tMnwaWtZ4wdCVg59v27iblj/AhbA/UgK0phozGPLKBPVs
GoDokTWlyaWE1zvXUqHzt1WzHd4qlefjaHQ3S/iQ0Rq3DCSXrSIvaKiOuyazDyE+
te5r1HGdMghyT2RyuOHuTvIx9omyV1jbCr60kYORQB4vgeBqBkRFcCq0CMHiNuba
Bp6Fm7/HtkLEiCGYxhKWpYmT8dkvvlsFLqX/bffpQ7dG7MOQCSwTQhTDj6dos4nr
3K6QMND8T1ANTjM7WXgzKR0mhbd4GXje5He6cVYQvtJQEwq3615b9UK74DkHXgVj
HGAHuGvffUKY3HOjKn/s46gqyF466zxNRw6X1f/qTGvdWrWD/uqX/iQoEAkJBiU1
MKaLRB83H/jHkKBvdwir06Y1OkgU8UrDvFsd1vefVnCkvi4wQpz1sXfurnmTGFVq
T3f5qhY9BklU+SjPWv5LOm+/Z+NT5gVQNky5AdRfGa/jfROQPX21c1s9EAffaHEe
aD30NvZsnw0O6pyWi311XWrkxv9UqKx2GfU9UV0p+sLNqayjWG25+vUnYnMtpLdW
BFsBEbTyKQZdgi7IsupwRUM8cPdHshda/Zhu87Zaz3n1B8lLswQKXwZNjdbfYU4T
8AYNPNZP2z39a2zbV1n+RGftLiQYZdFguxG0+iUgdffXQccQls52EOxKjGCsuVbu
/HknLXcyVGtcCEEWQKVgP3vWMFBBu14mReGyEiC5ZeoCxXWzSUVEjT4M9z7VvKeu
7beENGLEgY4K3V9DxhYmpY4fxUxzHKl94b0o44UjvdRj6GB30/iHaWFEU9RpVH4F
a5PQUAb7ymVO4ZIcsLXBsQLoR9m070J6bqYI0UCgFxBUaZYq8dYqsm+/HR8rO0t1
SBcFspKGwojLEraCSA9ZvSuJgntMQ6UZqT6ZMqmn1cbk/WxQnhZ/wDFrlu8DJxvD
mTdvmk/FUzz8tYe3ilLhCdBBKqb+QafqrqVwAmy0dwgRczbluwt06C+7V6zcSoJ/
MPFgaAcZKnD3ma2+aGsv5u0kkHd/wmqMoYEm5box60/Y3wf8ryW5NwX13/CIrCgp
6sez+W+My6GPg4LHaMbo0wusaQuJIzV5uaIaau4AjQTmbot3aPvCR0qhMGdYcrSi
ZBqq5D+DemPLkjJJB+ofAW0YcVGEdg0XMv96+BO263aVIsR/Onx0d98mJGjL1Ejk
0prM56VjMHBnWk+yBjyMDLbt/Obha/mymjMwTtAk9h/4u7lK69JWrBHsGGBwoPa/
JkLRo4ERkqQfXHZDKE7i9pwTJMg8qZv4JGJUTPBXJMywvhdqzVmP0iGpAdticVSm
l93DkULD+p2eYVmdhh1T6sqThH9Ix40xG4/qFy5oDEmnnKZe5Q64fUk/mJM+BqDr
GBD+gbuxmcI+vpaelV7qHhsRnQe8KlS6tyQSLUDQSYY2rg9BNOVa+glgLa3vwhCZ
je7ctDugeMk/E9trwvbozQRNxUAndTaZqCeANayAuSGiMFt3D8h5PwvFMQ1NB9qc
8virJ0O1c8Hp2hJkZH1LTttRcsB/yoBnpkYhVKvFckEOtm9Z8QtKUtDOKN7zntzJ
E+vmrnipgxP1+KwS+F9EhpfeGtBYPfYBEeU7neh5oQaEM4/YThR3N/OCzpIxfrHX
u2Z/VsoBc1b2L96l8xrCpCz7zGEzMw1tryxk96+eFxE/FsvkByWya0i8SU7qUEpQ
15NDo/CdPLwPEGnhRiWximbNo8F5OBXG/vXcupDYUCn+jKS/hX+9sXQEsuu6SPx9
AuBJeLVQPU0sxs7ECOsrsHPA+pfzEgyEna8pUnB4urN9/ULKwbJjuK0xBUURxrzO
FO7b+17gCgXaGDHAxxntUfCmqwkZXSLKXVd4QhDxuFxohTA1FKWKx9I1oHhAQLol
rWPwkrXMsXZFD+12LOrCGiYmYZRJ0B9f0ocax9x8OkPpdjUNoN/8Mmx97iG9U9dE
Xve4+nil6wxrk33/dwMv5Lt1P0n/kwcs/7AGsWTC2YDGxf6LVaaIwDpPxhR2Rjro
uujkYfKYyPFkPT8qtW3VEk6EAscspQGXbO/vt3qpNj8wg+auzM4IZRWzb6tCg5Xw
kgZdLHTl/+xizzXSMOXxQl58LZfot0mFi2i/o7s4+37jy4DTVFYHyuUR8aYGYzyx
YK0rYDj3JsXiJ1OW1tfidDOKc/CVkPK6jBCtp2su++4g1mmCgVM7aF48qnZCQrrS
wf8AcSRoxN6vW9BUC4Ze5rkz3GcIaTxvzsSMkm339zkmJYWWeCNf8WXFcnpz13DE
7FcGEw93wtcnyckg09DNltK/sFodPn1bl9CIyIGwwjMd0BAvhCX0+AtmBWF0qBDB
hb4Szv2NOrPKsZjrsWdVZg0cGepTNG7/ZJ9URFGxciQLNPghOi742MGZtAkJNF3j
lOsRX1myu/iM/ckNHUyxVDKP+AFd/pCoqLK6Fa/+kXKs85i8jKxQomrV4dg3d8F9
ieqJK08U/0kbGLXbberHNdVX7E1WUdUroE9MFm4NHKX4cGzWVt2aCzUCEB1peSAu
3yNbv4TPFTXj7Hswzwxzjv9JVNdKq08qDisThzyjXKE4e4i8RJlJwonO4AfVKQAW
9DEYbjZCqZtpe4SjSssUym0aJKqfWpdUbMHZuJB98aGgGNDsQsxTNeDZLnum/DfR
dALbsnQIetuYiHObFXAUQ7Q8WtVioBGW2L1K8ycsblS6E2IGyJ/khFEf92iwQg8c
OkvPUGn5oFOK8pcZEMptgjA9sAuwminTffjjJylirsc44ixe8EAvNcWlcFABAu5C
eMO9pvIt4AIQfYWrMIJMG8s9Q0uh0df71V7MDEfLYABDMUEUv0WQpmJowFNLKMwY
M4ucXeWHvGxV25fbM/rqvXa9DIlRgj9PXNNQ6448n5kdKE8DDGL3Sc/HWxybT5wY
sheJ6btM9eTcOt0gyyMWhi/Vkfi9QKoz5yHH3069jnluUxVGf7J7Pk8XIAO/7NzY
FP0zJJl1cig56FcpABVBCOeGRoUUcHTSjVI1BzBKEqOBROzuZbHJed8gxCyUSXJD
dn9eifim2aPaPlMRl9V7mu45kZw0O6NLiGA7a2DqH6RD0cUL1CdyYjMKJo1WNq/B
gnOZjQO25S0gykkvAE2dRwht0CAnGgpTypIij9L1S6qn9JzQ2oTafiw+KvzTh1Bx
8XyabHYZGKdFHA88+yDCmSoJcShdW5UA58MzUTvMhhFA4as8NVPC/DR44zUNWTrV
ntqMrqhFOqhy9PyEljTUyNrqY0YploW0FdMgdqn8NsDFYxeUhdUylGTmxRhMymu7
Rlx6ZqvhbFFBRj2x3ln1WzjMm51TRIwQvG/1A2eHD68hLwLOe3Q5kOVEmLmwbwsC
v1hvrBA7OOaFJbvge+Eg+zuG0UU6XVDmAzxJA1EayAysvsMq7odAQx6D+D/xCAP4
WLkCvWKyvg1d7FDEwrwX49qh8gm3YLK2ZVmavTRhtqH6qrW1XeY+dsjEf7J0UOir
acOtoyg+xPAOHxrNTbY1/kGL9DWkqHXKjreXTweJlOSIYSYrv1TiYOxSHDPDtgRe
sqN02/NvPDKjzMd1j7OFb+4bjvpS2NGUY93KYn6XSWWKC9kOOiobWnA4DSv+4uGV
axbfrKXCS5CmKkl/8BtJ8IBsIepsjNE99sKXqePG0Q8vmqsaQlyk5srYv0g10KPK
sCMhLSPBLTdwe02lEmgtCekpJdxcIQlcy9SFl+A5ylNbBibAE7bVHwY/i8XavWuP
B5FaqB7tYDbCqhU/Y6e12jfFoRCmlwRbAnm/mdWFlyw6gqWrG41Woo8RVEN+jLEW
36vBf7MedB1+Z+/YYWXroaRYsf2Of/3mwKbXDuCGuQxwiwJ+pTU3Sl4Riyi11oZZ
OvGw6ED8aiQkf7OK+FBkmVxiEoJCmeafGgESE3Ghc7kFkkVUVStEEShfnVxyU2F5
IjHM9Esb8/ObuK9rmMBXdQBqbMvXQ5dZaN5fzEzPOiFSgeYNL0RicTV4CwTpszJa
nws75anL+sMP45XUZcAfGI5xfTZMqUAlotEBS4tWRm2OeMLSqG2cjVYC2WeC3WIH
QiwSOosGBn0E8Tqx/sOCUo64FAwnAvSJZBX8zAwRdZQ5Jk3hHYkmCdcUFGCVrLhF
Qa1Dhed0xrZXWh7spinqKFOeNYMOVeu317McbBXpiplg8EBuV9lEg+VeqJ3Get5N
PhlAxIozHoT4Eh3s+wf0Xd4UZ6RqietYSJjtLjcnmmEKWDBmTwas+2CxqiXXiQ6+
UIe9CdWkDyK8fboj6hWbxmnDcvxOXOnaRivRaO8eicxRBU7+ZONcd6UH5tVGKOSB
OaN61l0C1FIgX/Q4qUutIh1mCsPDXNjqSEseStbqIuOdGDUzhnFOv0jxuTFzxfg/
b6pmbvYttuUAN8+Bq37rFaqvfKql7nQG6A96KdtzRFBF7iCr01iofmxKXex004tn
rrWlgFF9qo61aLOSa0Zx9lGyn5kQuMXSvsO909YbP0YDUE5GDOKXgkDoHKSO4p0L
7Lz3RJK1NdiGLtCNIXlpzv9cosFIUw016qdcpoSGObGrw3FfgxX2k2loZQtz/YGq
BBjC64VXkiGN6xYqK8lt742SXfvWU+Euf6Gppcw5JWDv5AkTYVqVugl0aDGs4gHk
XSitNLI8vR1mqf9jK2Z9PWtqiouBpP/6SLgANOt+YS+kT4xUTmxaWR635MYUV3bI
PkE8cEkvCgn/UkeRmKD+ZTjuil89y/coHoeu+SfCmYLQLl4/zHZZsTISFVYe2hJl
+DlBMKSvslBdYGOt/ShEaWDPfM4ZWRgSq1Bm299u0c31QgFxLu89BxwYMf601wgA
m47pKh6Rg3ZXX7MgQmRIL74PkLZdZUmU46NXs7X5J/8/GpqipFR6pwZ0M1iV8vdj
vNbK9AGRBRIaYtFGAS1qexu8CBlw1V7kmcP+q1pBONR5aYpyErMKMJOoOS7wDkEJ
+I726+uY9Z9oJdjYq96Tu6odLFMpl3y7v3CGb/ypW30sVjc1OpQySGVX4LdiAhfI
YP/r/hfpVJRMdoz9NH1hQQK2S4X2ZJCSeNVHSUmd9+wISlRuZz6Yn8IAG/f87fMh
4Zo8J2guw3m4FNdhm3g0+q25a2n0bC4FL4q4iETYdhwxRrqZuYdT4Z7U3j1MxyT1
KCCd9C2jTV5JQdGZPmvAPnsgqMoWSrOqbkcy8of2f5H42rls7ZrbmD0KUtyhEd4p
z5HCuO2PUWBX6tW18MmymcsLFJmHpIspq9knJnbjtmrWPyXmUBzDu7zY/zhucdpM
llaLOKPiZtHZkgd2XNmT4fqF8qGAOqEEu1j5IyqwS4hngX03PAIQDiGhjeYSdm/u
zkPpwfwp8AS8MdQiWyK/vW8IMPpZPvcEj+M991Y5w9RMjqTibkuO9R8cLtZECPgA
BsDyoyj6Fn3LlGu2U0/xvoRq5P+6bbeWDFJdSz2i7w0Aa+5Xn0jfePu41H3y/BIW
VJN31a6dti7tHUEpvbjG9N4p+snzi2B2asLJcBPuViCW3n4eZeDnV+hOEl0gzMZG
T0Ncyt9WFPybpT/2TKOxyGXcJ/jYhyHLD+GX8+f9gsEJKCqQGoHfbx8pJ7H/VaQF
Nz0iZdnXIDzEuBj/3nROOJa5ktVuobP6+sFK8Gb8iRdpF/+flIR9r+2zlrvX30t7
vhZb24ppdU6789ExC5HD4UqKEpEc7aCrJPfENxB09kBYnQnres/bbCOkuSe7OrEW
1XnHcOD8Z3GEMicXxILMEzM5mtvGdsmhmZWKV5XEQZ1vjDmfpcasqmsLA/SN2pth
eC0m5CrTCM64DQ0nImH/6aWRa6z2ZqlkU+sCLER9sSRVu3yEZRwCWzmYAV5kWXbl
Y2etEimqh+hur5Gw9foyH51kUMUXxaH515AdIP8SWL1WKtt18xI7C4si71K10R4S
J7N56iHsEzd0Nfn8dsU/OJkzlbkaQSiljZMbIUskmyKuJJyLdaWd41scW8j6HqE6
owGlL/nemxoEpBSsXv6KGYaYajx2PF3E+ziKA9dJNDhgZ38s4uX49CnaH/NLO03p
uXWyU4CnG2n7Pe1+hRdBlEhUJKC7zO1ET37lP5ZcsazFaGBe36iyefHOUsN5jSoL
winYqPFIU4YLDNXM6h3kvF0KoudsQPZ17SKMaeVxKpUuXMySG8Vc7AmBsUNM4BYN
+c+6jn8EpQf2se/koVh9yQ+mF843CyZlHsHkJV5pfztAk2Np8nCwZdTLYpp7ZJ7j
HDWtN6V/ERhwHx2BHbGxwVpBLJeNoMoUjmrfi1DaeJTQLCuESwl0LOksAd0xWa9q
Um8378SCLwbJqOaIaLenJ/3KOu40f5DMrvajHAV2Qx2fpDe6tSyEMUcW7zOjCz1+
uqW8e2MYwIbC9lvhOikePqB6Dlb60msHXExKqLAMVqMavuLsRH2zbUFnmJQtj0ER
42S1lqU9tmmTlbPrgNOCvzJ4hgVYmrjzIQ7oiI/kMsIq8BvuGf+dd9hU5p8FIXUA
FLMZMzFdVj+Wuaplv0r1AUkbGNA+rpFQhHDgY0Do7dZWqOhW0RTrobVPHkPU8tJA
nn+GlOlkpKhGkecWbrgLZzZdNqx7Bke4cqx990vrfJVa1xUISLsN0t9PdRGMFLWk
2FVRlYazkZmBv8p0wjIe37HXcGoO53rEtD0zgB08geicnei381TlZoN/X8AmLdiJ
ytsNBWckaixQOR0Qxu9XbTMEBSR6yn2J3LrvPLLThlBZLXdUu4jalr+nHKUNj6VZ
RNDtZ7m5pc7CsKMZ1hH3ZV77Z+qdj78bix112Uo2+Cks7byMh1sjTv6F71QzDqkc
JoWtu9dEFmEENonrIVD3OvTmTHBnMalht4lSwIJFoNoVbe84n3MrtD6FzBViW4Fo
O7B2NOUYcIn5bp1G7DKP0BDsBnZpQyD40qEc/15KiYGo5Rf68caKseQbGTDi0N4h
zwdZYnteehUhCXucsbpgFvrW090hMqXbcfbF6IZpePnamZNOf7K5j6wp0jA2FGOi
EaWQZOJasI6N/AYJFaSnexDZMS9YuVouDvFyzILkifG+WCnKuy8i5XDxKndHQ6M0
+/ZkEORCvLYbd5EawJDeS41EVZ3W0KkFYrjHsnksBVdLCP0bwnlwVWamQ1K5fxAf
jnCpQDv4a/jZwnitTTESyjv/yVd+42LJ4EKbmOL061+dAgFJjz7VN480QPqAFn2r
SZJ1fgXv0//z4otCJjGBOja6/Vie2i/qLVmJWPv5wx/Sxt5ZAY1cp3f4yXUFgWMt
wzC6WjcRsTBfr8Yf38PKJxXW9OnaAc/Lpv0XtrexOxCnK/hWltywpEFMfPbYiBU9
qWDZGW9T2LR+n9OdFIFtS+RHeea8/EplQcYV+qGT3e2Pq3WtMbVN+eelR445kmPq
QiosZrPQ3S2+L5LZ9bo+talg3U4JNbJ0EmNmphCKU9pGp52UNh20TDAmF7kkjL+Z
jBTYIfN/TuIHTC4nWHCHtMoSCe1d8CJSAi3cbCI8iB7gSAmSEmGNNAfxRSHkodow
fagMzom2yTnwdM4NYA6RnQdmixUmA4rsPhedrcKw1jUo8yj188HXu5HrSC/ZMwJC
7V9d/H4L1C1vmTZwNaN0UClFGR5XQEUJJf1bj2l4fbe5+/O+yXxQRJf9ltC29+Qm
0sYHBf4V8zl/etd+ZUyj7H81gXH62idJ61qA/Bu23/+R4yWcMDKnZOScCC6q5xPo
OduS8LnMQv9JSnaw0xzlV+yrNx7drsElqAqfF1A1mW9JSeP/g3UfpOyF7EgCXd0Y
fedgMqN8wverIJ2cIDCARxYVzVihZyVWrkZoFGzKFMANUV9iE583YrxjjIzlHGyW
ipWwb4bD9qkBn7gD0Qvfh5Yb7xOXzMpUniNLEPbrOQzQ/sgikIgo/Z6il52VBqXt
S1P3mOAdD0nXyL7dFtTnF2s36gi5pas8hRbAro7FglVNoDpivGc5f9oyqYrXdSVx
qIfPEtGdR3ZC16iIjU0wtHHvsXirergph/kfyzrJBZc2Zp0yUSNELzqoDPEe+ta7
G7GFaLWqgHro+RCYz5jpoJcdTDDU2d7rfWcDlELusYB7oLmo2K0k9HxBR3dgdfsP
CDEJ8eSv2+mQ7+82fAHmhBDu4kQH+JdjQYJuxIPcY0IBoE2X9v89fJSZUbyAvHJ8
Nj/8pnpK2tRBIHrjqPwK3w+a3it8T4il+VpK62N0ipXuVFh/x3lq6Ck2N2p9qqo7
n3tdeVVYGI56gVqbjfNh/kPsec2g6BfoRCSNMwAf7+g1aG2YuCY+ycTCbdQ79bvw
xMrZKLkcwvldS4YiaeBBtVAoMz5i+JZ4hfXyAo/X+53OO+nV/MQDQJI/b1D6irIG
Gge2ISRQXoZbdbnT7j+z45UnJh71BWA8YDEAod68jvnvAa0PwcXritA1K0vX5gsT
q3Hg4prKq8c+yhl9E8ZfcsYMf3c9x8HYVRVOjrRALnDK+J/PGvJpFEpjMIgLulwl
pLQdJQUdGRMmq9T3GvRLkFm2DZipHsCtSzMP+GzaatH2/7KwHBDs9mvmImxN/HT6
p57k3bKb/7bEqm4woykrg+I/VkRphVebU1Ia7lay2724jiDy6mlpNm7cfFYj+lfa
ZChk8vUn3kkTnOJpUm9HKDTAx7rGTPNA0PFbZiQR/Jdds3mJ0JCT81sddDZkCfPu
+LIlnY5BhTqzYwc+p55E2XwJPFcZUlWMSQnAitGx2Rwdc87YME4m8NZMeNejVSSA
NfFYr22/GN3m2B4MaKIG8dP1+WKevx7t3lmmI/Xd4g5L/G0j3G9YWozqAFmSeQR5
DQf6IyC4zj9GQ7kNbs327R6pBfnBSl9EgmZmzq4Yl+go93DQUedaBQ81NF/5tDmK
N+Y+hh0KMkI3Hwo+4ZUYBRnI9UVX0kaHb+zO9Z7mrwH/YDFbZkjwy20BOqDXYqWg
xqjycUm8eBZvoSWxGwDiiAl5if7rVgSO7H4JReDgbPnGgbnzyL6gM46sL2hjPbV2
tPczIkDUArONnp5pzpll03TJh7fNXQnEh/bXTn/oTiDyXQdScWdsRLHu4L1OFZzF
uIqAvEu+fqph5BTHFiv3/zKV2pLAFg/Q9hIYyS7LaCkL3CwHXr/TQ2quYmXwWy5Z
fLx2eitCEHMWiuywP3l+YUvDIQ3Uz6nnujq2XjGX71uGxVB8thDKWgTwTV5mLXnT
kRoJpzjqarXHJfLLqP6zPBFTll0Buy5ND9fBJ9FXYhuULLs/HGIZtRL9+xw3orqB
/E18O5lja/mcOl8K+JJdxHHT6I0FASsgBUA1kDeSrKEbmvCidS+iMAscPWULNHPE
x4neBg9Tjjdw++P4LqROJI5jLCDCMKt4mCmuqvKNU1iKaSrUeyYKeLR9MW5CfN/e
Bzr6400GjdKr/PnFBb1dAY8G4fgZThNjkrJYCbHUe+Dyq6q29WJ2VOhi569C0YHN
iS6Uz5EH0CTRP2CPmqccte6Q5zMZ3nRV6o+gqMQlQCQPkmndM5AwkpIuMqkqqUG4
w5mTN/2+N/dBjM0Rv3WwThfAegmPmKAR9Zlb42kkPX22gDwM29ZLYpyO75vl4Zhx
FgVAHmKbp43QcSczxiRNCAQgIRnNdA2dBF6PY5xzmMcsY5nKTkp0QRlCF9AAsN6K
47UKzie4OhBM8XuYjyEjxUVFC1u666WNdAyg2kqx+ySMcISGLUGiUnKbk20gjzDN
2mvZguUQg4jeGZY/g7Gup3kOWEALY/ibrJN40EY6v97Ev2PsqFtVQScFKxBJfdhP
8nIMeDeJ8uXHbC4Yuj2v4IlmfMLlMcSrtqt/zPFcVBEC8K2kpG3YG3vQMCbylvEi
70/KtxQYfnqrWUiBxa/le6Lnw7Lp3//XT1Rf7l4V1zbBkuRbjMyr+f3AZobniox4
ZMknqa7PEm7hPG9rwr21tI2HqAvbv9213JuhjrzLVSd2HrSAOOTVZRP5CCKLDLxP
XlT7gu4qPPJOcVcS4KhsH+WUplh2lHkZpUnCqfD+swtFc2t0qX1YYty1qApHDlYD
Udc3Td50PyZzmlcqb426f1dxqxNHDFKWyDiv4ON5TQnRZqxATB96cRleFvtzz6Z3
N9Hs85TXLBRP67UnY42/G9ssoUgKlLtmQwX90JiTCRxmMGW++rX/fZDQzG1c5/Er
aV8e4XKR4kozTxPULR5/0qnLTUiMpbDTebiC0047/Jl4aBc2wJ8DrbFDpIzeim8P
X2ABMnFNv3aR14n16MwUeYwCGM8+D2WVhRZMO3G+gASGs+2ghxl5KvJNiPXACPFw
536nQwcO2qH/PPng5oq2TJHLbcvpTNAhWsg+hxyl4SW0SRQrccNapvQAMejPh87e
DgU7FhShjTLnNRaEih+HYD9iwbPidZta2RDRi16Jr9v6frEkRg/aR9zF0VtNqBC8
L8ClohF6m6LNQ0/uy7Ol4PPDsE6bk4OahJgU7/QgzBRBVHpYlhchqHlj5IQDIRza
kFSqABUyT6L0a2X50j55iU0el80u093GOwPWI89ecWHSgsDKZKWdAm7VUxuAmH7h
ki8WQg23qyPMRvM6cwrAPWTCfma9dLsZPgDtFgtGigtUgKQqJiGbZZ2VgcPjNYmS
wfSHhD4ZzfB0zbPCCx/Kn/+NVCNIyjEISVC7x42F1RnRftB4k2TfbwDCkBYN6eVx
n7exCDEmE6K6sd8JsWBe1lvBd7A2TsTa0VjqIsSXwoDR5FS11D7WKswawEJyKMH3
MBK8kSY/gvMob4pP5S6vomZs30MCJp8vNKVniO9J06j0293dgqVSPdl5vc5U/0u1
GO7Fqd5ckht6//Xcj5HXJ/K3mg8EnUVAvU7b1gSmsbQmULUiVFa5GBuJRzKDJvIP
3d3bRgxqGqu24ToasnC4Hy2h/StUh0PhfPv6O1SkFKK91XEK4iFKw9ukr65n5tF4
oPDvBRUmVeoE+sdMzQPZjETKFYkUCX4g/InYKW6NZV5yWvAk5yoHnZu0yBw98Sbo
ir9k2NyzI+SfGerWHea9Hnm/h/XRgek2wySi3sj/1x/twi+S2XRqEMikHb5wvlCq
DEa6fxhLkJt/G7lsDR3UpICEajsPO+vubrG4YgI3ocmgZnM+/Pwy+VU67H5rqxPb
lKSdobnhDQ2asla+45+Qeiwbc0evCCt4e2NyRp47tyikgCALRHisULeYk5gmm2Ss
LTrNgFcNo5VmPrpxxsyya9qwYKTdyev/NZR1xenQh999n9aO1jPO6XnVqsehpoKE
+jGhC3x3HCr9Og4D/FwMrT/k8Ac8MtsurddeFH1OMs4sW25XczMa9tNNN7aa1cL1
ivVJPiMLUTy1I4LCVx4P5/jAYtpWkBpXAmgjZ1Ji3nXxx2V88cy4uF/OUdc+Sp3p
iBUkHvo+DyI4kkjoMZFgu1gDwGoza9ZDjLJeq+Cpnzy/7cZpUIeusQq7cRTd6RAk
Y0llbxERIcmk2mBFs24YVhdAVtgRF6yc2DvGIymdSIHpB7wCKsiW9RvxyrOehMjb
3L4MyqYVuo1eydkuEG0FjkqqUSpcPcy3oItGej/jhrCj+HvNmEpSU4XlDwTFhOIW
JwY6YAUe8B7ufdZNoKeu2KKKtpdlJuIWJPOKUiNn+ztaqMnHwFWqJ34ZYPHi03Cp
upq9Q4gy3xAAsblzft3OFTVsgCr1He32qOyTf266W5yENWEylDGVyeuAsABc8nzB
8FdnpxUpi4FGRJUD1ivSrRkB3TaWV81dr4P+I0DpkxX16EHVAkxh3EbaJZ9EiiNV
f97wwiPs20PGcO3/g2KrYiZWkznWBGxXygeuJN41T2cZOBNo11eBRzsem8dDsdNH
0b8dvDtZSSc4oMDm6e9p0kPew39yaTLSqoHgOslYmIz1saHu/efPBhXY+er8LQDA
ima3EsxPr+A4E/XheQV1JBBjFOpmesrSaKNPeqRTNQOS2G0zak5gf1/MZtHmpUba
YBA4g2RUZmcNmIjCL8+Asu5HJ5zOTP5InotCgtfu49aKI/jeQFIjr/2xN66bZiVb
1nY5mIHkSIEY6oAn2rt4JipJ5I3gufbocD8D9XH31+gbWXlH7VBjLj0qhJSnJQ6r
lMHPXQMBjBtePixut3+6nsiq5CI/E8001Ojhr72tSZsL8+x3nIZeFBjdAr3umHEy
148eoNmkAWk2o46E5AgHRJ6nmag4pUnDiWE/Z/C6brs5/+42uJFQTQVg7OQnChMh
bsdeHq8rmaUbx+X+bwVI1BN/SzgxefKpalgSJkCig+cPsouAsfD4YyJWU+S3GTad
ZNPZBHa8xREifQoS/nIFwRbVrFgjdGhgbxh9bfbwpdKhcrcjGoCOo3RUaFoASwLr
Uvr7DRHIQdAn2fxZBwJnV2OR8uKq+k8DxRUjbAn7/NYpPS4J/5UIt22NeaqO0Q6W
k85L+fB9OKWyCeFuIbXDv5mYPQcptpgIg+HqE9ONmQ44zkbWXEGg+Ordbou32FUk
SehZEE+QNuqFisfy6cznM8vieiACIe0p+3Xw0ZiZNKXczQR0g2jhzH3l9/PGQpfw
xYExDyQMbRQjqFCk6HFxOMmSDxOx7Piydn+MTtDGMOI5WooidBlfAu1WNDgzjRgL
mkHts/3ajfmfTq2H2dK+OP0RgjCE4KeC+teqYvM4SKmMGPji/dbAcMypr4KAj11u
LOcAuyPvzUN9NYLPlQH+v7Txen5CyaPQlQDWnCYmVUEOH4WK4E2ehi3ZRC9TIgnT
hls0VaDgOFG/wdjfX4Om1iZkZ0yq4RKjz1lWlfh7IG2UPFFFRr6surRsXbRDnOdy
W85xcB1v0apaBT7CrgTG95mH4ls6YObt3dzpVOw6SEm4yKbjObGdQQTNFo9LlJNV
DikaNBz9RRZgZXeJn+fRmLnPPrkXl/UFnVoYd9mnDNwJ589l97zlfXutvozajma1
1eCIUBOQt5/QKZrHws6ZnAFVw/16tzryUMK6H4oGtqJZaMLVREf/pFQuJKO5THSH
TMXnCdii6dzRvRzIe7JWqZD7zx+0dmoHVu82rT8mOGzl5WW0zzjhP5jyOca0vs0K
5SOUBv4Wf6JtwZ/ay4L/OnDpTaKGhSnIamGga+G3KoigtWYTIn0VUKL77turAPb+
UoJLGlgPv4p6DUj0nTy1XIQnTS1S/Ospk42ItaaCX+kZqcBA/MDFIZ3OGE1i1Fz/
ksX4cZ1upMVqx/ujL1cNWYdzBfQ62zOhYsAjEadhpkurSjFCkwO1d6d0xZZkZ5sD
ZOfy4j3Hs08PatW9H095xgI0v858cvmJjzQW67V6iyTzFQD2NVGOVHik1zHTseTY
DuewIQKnRszDF4zrIz/G7wfV6aPqVGXBn7LPNYnt7tyPXEnTnlyp4fLH8r5jRUeu
bXxcaDnKepZYOvogghP4DeVRufp8OPQQon+Wr7B7Lo2azoow4z9Tf9CbLqZtS8N2
sCFYruOfAe7exciw3Kqej5XrNb34Yg8gBSB1mKtPR3NAZmq9HFZoscGHhV66xW2P
qGnOC7oZACo/oZhnRR+d8XSnK+auBkr52F5TISe9Wa0bpx2bC09embsDnLLYI2HS
kkudIWGCgYLOHPCUz2pc6j0xIjCsN0+gum2eAHd6mEn/fFxDF24AKoGwsFDCKCeh
JM8mBiMcAZzi1vzR9leVhz+1faZ+btkLTUadmpQx1/rsTKFyDMQb71JuT0e+NEvw
08+NtU+/B4PR2VuNA61Yl3+dc6jEOXTyIG9BnoXdr+j5RqCovfUp+kBku61F5zI8
B1BCZt8eSY9gDi+DLROADd/IOKNySpjW++F+tpdYq7da2x+wr2U/mXNZ0KPZxoUc
Nt8dhLEx7pffNd29y0rEKm8KE4ag/apt/JBkaY9avahhg1vKl/EWzCybPIj6sm2+
rL/qXRhmkhn5LaOkML5/PdCRhk4ZxKJpH97jxQyEckC1nuHn/cfpS0BhGglIWLqg
0anqN9gSJWB6B7oac08Cc9VzC6E4JNfj9taoXiabi80uHJMTt0fDs8n1znxO4u0H
jB3QQMCrZcNnxLSuXKDEMCiow57ykfsLAtbnXODql+6/qleudpL+s3Ym3fQM1zZC
gOLP3blc5jPd/QLjpTK1YRTjfWORH5VK/dC0xa9OPoDPyOLJe3XnNsP6jwze5HRr
OEBL+t+F204adGDrP/8llIKqFyodJjBD37BB2cEMeSbLOzm9X1WrYCaiSBkSpyon
NyuBmucRI5dYxRRscEEgl79EpSPOmsXX1+kyfHBw6xtBTcMl13FVfGfxJqpbTFam
MNOVkkfIOFoqxC5zBNjlUcC0hQ7kreHUoW0+WDTnLFs8JRqJOHthMxd66jpe8rg5
a8ePmPoh3zolcelkTiMNF7Vc2ps6+Suyc07hsYhA3g7Plg3BvVWUlYsMFODZhKZv
HvjGwbFJhe3wUG9RvVvH/bis93XObNEshmSbKD+bgoE3Ey72ZT7Rv6AGKpE7mS2d
7AOBNQGlYWjT4rDffAzElmFMghJMUtMWwkSe0idXAQqXQNRONjP6AbTvfVjlnmQn
UQffosIb5mGropHSCTXSzNftOw1VO17jHf/3tO6N9AvnndkjonPZ8Odj1aOaEHeq
vnsXM812cEsu1+QFyE1ge+turZmuigc/1a1fOWTnlw8QYWJQ4l7Ye20eWq86XmdP
NM0VEBPmreyCzvhbpPqFrxO7lXB5bQxiO9P/kl4zZTw8pOMmPROEBTdVoTYX+wwp
JkztG+ZG8TRsklfYKy6R7Ypv/YOvrajiSsw+JKVlSaQjwJXU2M0DpwOGhUvE+amH
jvZTvzrBvSuLGmB12aO0a9vKOgPiKMJy57uApcjnAWB6Blf0qjjQsDQzBAnP1ahb
v2ptD+rER12Gwf8O+VbP1LxRzrWfHzTe5593lqfQR3THcOpitpmPluLoOmlmyJq7
ARAoHLjxe+/iUqfKvbCpXM1xgC24QiZurRgynAqXavaPBYPN5zz0WAatRaQWG1fm
KjI/KYNwgywszWj4bh/3WUmvdTMa1pJgDbK4WAKYErWmsAP7NiW8OvtWjZs3RoGO
h+JjnmdBWHs8OiOdmdDCr0JASzlH+tf3XmqzVvnopI+2/EnADyYQk7mOdExJJrf3
wF/irHXLt2+04xQZN7KH0Z+y4xqKDBPxTfntEnavkuS9JMR6PDcMyM3fcx0Pw/6J
B8rl52OMg7wNAhJe4jgY4a3jldH4pVpO1suZAchb7biqpMN/zQTzXBPTJ58ktfIp
fdqaUQbS83akBGVwk0JHZR9uJ4/1IXJLu3QUBPvubn5X4aiLlHK4fvM0CmfLu3ps
QUTAgXsBzD/h4w1fFoWJAOxOlWzFjsFldS+QlDU/s7kuF2Yp+M9dW8mEaDqVcE93
pCXx40scuKJ3Bs1CvwEWY/sMg1QrYs6eEHXAI8JmCQNhfsVWMCVKnrCOh/XTWmxU
DiGKOPzTs1Cf2hQkxsONjG1ACigYlBza/+fYINrtbngeWTzBOBD3386eBW/QLrVo
XkTF7aIECODqFEXtowsmPxTXy8KGHnwuXXptXYxig7gE3m7KYqTy36/vogAqi+mk
bJaB1a8utXxBVwYjQdi2G+PjikavdMe6EeBQDxkfQXe9OzUHNh42htXy0wDJT7cy
vy4RIlzeWQ4pgktoadFDHE3JblUMPhHuQVJhtK0yQ1UPL33hy0jKtPy/e5jcSW98
eStkSWkbzfiLYv6SJ6+RhCdTiSEdzARR2pTZlA7MCMgFzFUASCWkDMMCmo4+zCvx
wkxV2K9tSb22huw1jwhjIevB8rkm+1Gn8EZ+bjSmUcPd8LoJbEvcw5xNO5CYRT3D
B+jZeHex9mGNi1X5muwDVOLNxdrOUxh7EdnY6+teHrzOchPQcd0P6rQa5s0WdxqJ
8WtTHwBg+6lJHrv+kU1sLconGImlyaUPNGqDqiI2nK4MO0gpYNLiQDRcBrvUXFUn
t1jOAK/blx2Ol/vDOGkp+BNBBud084b4gggIQmnMarOnFB+x4RtYRCVCTALJmzkU
JHOprECUpUeAN9IIB5q2FzZKBm4uIrDbO5IycfqR72ucC909cGrUacm9CGWWxNN6
mKwJmRCu7a0J1HTKfmx2JstPVBJli63EKOYe0nUEWNBsHbyX5lQ7Cbo3Bm4vFT+z
cxIby0hq74D7PXqsjFeiwke8NJym1ipIwys1vv7f0lqvdagO/ciAYuqPezyi+GlT
lQd2gjcH0xxpIxYYlMxsSjHxQD7p4kvaD1MRG46tJozn9kbdn4/zu/R6XRVrgx40
HLRn0rVBtvKDv8elmK81RT+zGoMtjlMsMJ0E0t1Hz21XDoaB1DeAyo3E9ASnNapJ
rVD8qMSTqDflbPuW6309jhP3wjaG5yY3NsyNjcV0NB3QwjCGo3Y5kWmbx4wlGFb6
eIfqdVasKsDfnGtm3z/g6Yn0gciXTdiqe/ENvElvewvKy1tGXFeQUUulbJbjW+zt
oWgy4JNJF1AMShq9pZc79U21o/WvgTG3cykeWZGp/XWjKPt70U7Rv0Id0NKkU2gO
T5oCRKUFWG4hJNq1K5+xRoHHzt0j/o4Is668LYD4wmoQAT19gpkKd85WomYxVcli
ziI+kSB177xzfFow2v5ISpIflgWaMeYx12ITW76VU+Ewva4kxCR/MD/tCDnVTZ+f
H4YiZ9Q4IrwR5xu3pyJr5bdG6OmkqDZMVHa7qCgM4LirhKbacNiOSuVw+Jfezc7B
4cmJt5nh69SvLaXIXq5mopOYyQu09+49sbYvzfOn8BH2/J73xDHyWa47J7BkqLB9
NLATTgwN8qR4NbM9LohFojOO27j05yq+qfo3UYa+NMhxWTAX+y5UKIpkJk7DWC/6
7NXPLEyhj9drcNXti4x2s6gq6IO2yYu/mLkB6G7k+R8i7y4NIIIU6DWuaNLUB1hy
FqtQbYYhAx8eg7S3g7ric80LBjQAdMEq7xiU2TZzPIrEmGjjSEfJAGFydUAYSzGO
DEpPWxlndvpAr71WAGSXHrBNpwMHwvyqoXp6Zc2myjYZzrgBv9Lbkrxgxi4Kgp4i
RzumYCFPQfe1ZVki8FJhbt2ZWdDN4TUUuzFpFYNoKUh+eA0vZ+ftD3DUo1mwpB2m
5VAMzO0qLvVFSeqVEMzXGxvYjMhwkWaPphxSf22ZYnXAVb/2h67QuA/1QyMzPCK5
C+MNjNCvuiqj6Mx8nLfy/T8q8To2x7kfn4HivOYVi/hx46Zw0fXnSJTaM3XPxTjJ
DizBJackfXYDViYcs4spc4GPg4cBYdbsu7sd4I3FDUTeifLY+lZ2VApjEYM8XGCz
mYMVebbZD5waFezpWZlphJyFKRLGrtrOil2nMw6NNGPhAEhyJXVetDTIHKbHG8X+
gqgsM/Z0nX1dUKWIetpTk0YcoCrwNj+A9Jsv65qJGwa3oCGzG0YrGllOLO6lrkBR
bJoOU5694V4aFR32bxBdJA1c3x8/z1guhcVIikaeXr+OtVg09gaBFY706bbmuWzY
E7bouekH/wRJgw9TMFPpquxqJSVWZKywX1umwN+uDy5ALee5Lld8YFJCdywadm5s
ldOYkxnxjdLxST4afgqQCSCkRcILQfXb/ZEuOScX8pZvrYOryE3gHZKF8SI/406J
1wjyiuB1rZR9ek5Cm1bSSX1aikiJw1khme+IUjSaTt/VkqlguJgKBoCOcSk25vTU
h2YFdKhhIWt4oTnpndA3UXtasGMi/0DG93BxZAaY10UvPAhESSZiYT1sKboT7q0Y
6vPT8HNwlqrxlr1jQ6W7CM3o/GhX+hQF7uUiCPOAWIafxZa1J0ng/NZpPTJyQJrE
PziX1MLVkyPuzA6bUfK6N2KZVajRNJ754cppJm7QCKHBbQsxSeQUNrb3aDhGoDll
86ZZAQpR3DduChOW71iqq4GFqGti6KRd0logjPc0Ya2pZq25aIGAMROy4uXjaR2Y
6e28Wa29Qigz0TK+6hYUG/1Zyb+1lsqaq8gJzWeL83+oM1ySjwrwy9xNp7TH5nVU
aUUlp+MCkVyRVYSPCzRI7c91zqkejJrrc9lkOpKImCQVZXavvQVQdL8DwYN7l4ca
sTZjCxHtlXJv1m6brlqtwz/4Ruup+zyHbobI/EPtgx1/En5e1RvIi4CZpF4sM5Kb
ZUYWbU2TKT6M6SM8OSTTLe45y6E6lN4kzjneKrpl6g8fz/nEg4smi4t3Mkuhnks8
WgF7De7TMXBjMMW3AjMZMsWxmRJeWcVKouIlpd3L5knUDecu5EHl3Hc8SaBN1Vix
LDkTKYgtiN7hd9v+t8gUN2gptv+PwT/rDizJV7rdewO369GApVLfg7dHOJhyvbgX
KdvfpglVwpjyu13zF0kN2GKfnD/Har5fKxu1XMcLpgz7V6Zmv1Pzsa57ZKiceesa
KX5LGtqXwwlyKOLrFMNme2RaTYb21uRxbn7gwM7hcYobwbpJTWf8MbKgqYl0khtd
0Jyr1mZ565VMekLc58RhkXPTyoGWuYuxFMRRvhlPk8KG4IJj8wC5FjNRyhXVjGVh
Ka9qLNc38QhsW3cIjMHYvzGcGyZpCmx6LaZnVJDT5/aoHSWwFMIg4KxxUxbBcG9k
/FNvCdwh0Jmwy42jld1JQk69PnJH5Q0pGgz0dEs+GUFmwgScgBMVJzkVODjxdPIX
pBwd+f0MhIREOzVS/3I8YLt1p/hSLIdrlnrArQXDZPzwLI4qJ9unK4gnWYTg7lhP
Y0kIBrNxMVy3fjJqFLEnvJOewGiYZJxtjNHgsnYZxmLMExjF2XjaLuc7FyXDR7F1
IXSr5ppNYCxtcFpls9E5t9p3oFbxS4DIqViMxsNLtcwtNWaDUUlPv6vRpkFJ55SQ
WmTnVF1Y+STdV5xHU/H5+rXLZw5d64tPvpM2lpnhn05j8c6v5tkIkAR02n8hUH0u
IpOKkdb3sy/MQePPJo3IpPmUDCHgSo2saoCZSXxuXBVe4ww5oGJGMgcMz66Tdls9
9mzGMrHApPfuD2hI7v5Wseb440yHVctIvIxV2/kuNqPI177P3xpg5Hb+HQUksgvM
o5BwQtpaOL3vZ5NWwcKKo3TTAoMgJt8l9tl/KhBy39M67gH5+e2wBxsocFsXqHao
vB1jPme46TjAeFU0Qp0mAOq/kukizhud4jvvpUMXTAMQ/JFQPyn1SeGDNeKlvUzH
YfpT9ExnbPme2SYVOw4aXFntra379SbVlLtV8MG7abEbeYYjWJI8RTPjzObaCduo
R6y4DDke68iNHsG184tLIVnrx35VtBkOLLS7PYnMZyanrddbMbADRgrpIFQ9Kz9t
Q2plLfUBCbzzxAFMBx/R6mUseso8zAoQSACKuta1FoOqxMde1hmmnJ46DOLOt1x7
pBYs4q0lNBJGeyCSPosdPcVqsWo5P3EVGH6D0E0mivjFsAag7dluQlIteVDw1nW4
7axygQBdfrP79B9DX6UyMrnTJBz970/gOA35qqcd2jtvS3OIoRJGfJI3t9pHGoIB
hF0L/dfrWCovJ7BM65B71mCv93+JDx+r5jZbizPID9o+MFmmJx/fYt9vNMmrXrne
AXXtzpy8nB/t6nOMbq6fcVyP7goLv+GUI1shGom0bxOozYJ9Gpr6tdDWPYy0T62i
66ZRhECzKVxKy7+UO+IkY+TeW8RAgWjAubKD+7FCFxtn2V4l0V+vDthFAcbUJnh8
Pxo6afK+iAZ5+eVgwiiRWXpNtiqt5mSri78/ScQKzJZbkBExiU+YWL7gRsmR+4uh
DKNFiSSHHrcBIZvw0y2QRcA9hB28WRXLp7QjTHnXZq5Y0d5DqbXFjIpWWD9vChAs
JEAyiuOlW2o70xK2eh5gm83025M2pQofSGctzvp3JHnQEwJIvCVudF7nUm9HOHZI
BFvRbgFRRzBDEUsW7NtTrjmOPLVmtVlZ8MNmzpsI4KNNnAsuKI4vNFJkalQB1NVQ
pGMrvROQwWQp4NG/SpbNeYDIQ8r312UENyxhg6K0T8lDSzHZtnl4kwlcsOhvPpsg
KyQ0HqJtzrVVp/5X01/O5hNNVbKY0MR1ItvHC7ujpABQihTWivomiDl5GfDz6QPi
uy1H4UiOEe0D+x4IGnG4f6yhUOqBVdDTfxR5XBRp/voirTnl5J4yQ22zUb/rjuv7
9GIiDjN5wGKvB2WsnGSkpPM3IaK3le5X4/QJfzGp2MoUqEC+GVg1ZPA70cLMQdmU
J4RQd0WGKPxRn/zbnCgZXxuDx8AU3Pec3AS2RwxIu75qWEVKrPoffAQv4FXjDxqH
9hkj9g4hwqIxaYCUqiizOj8Jh63OvgkTVRvsEjdr8tNb8auaJi7YpgqXJX9/zMCK
IUJzWKQ0FR6uMVVy9oQE+EWDWZ48dbMpNaSTgvZXJAGv6Cy6RRmdueN8PilU4V9o
nthDNejCjsyPfLeo42ShTtl1xLC0YIoeHkCJoAbYRCYHfmMukLGCPCwGe8RZM0tH
uS/L2R570tFYSWIMR6FswCGiDkIZtMldMH1zfWzirs3vDiit7cxoHO571AiIpjnl
Uo09dBcC1DmAvQ2rj/h7NLwRnJxcjiAlUSUDzd4rXbbEpBhcNNBD+5xUSyyCLFp9
i64mfx6va1fHYvDJRjrupkdTT7uIQZPPfYAp+9JxRwQottBByLJ6kR6il3afrvon
BG/lTUEXOc0EuZtsWeg2OLpDCyKs550gojGw3ne5tpGGv7gBtnK7HtFb/2XCcmjr
LOPWwBg9UfN/C0n/ALBRld1y+eujMVVVm8lyw9Z29OM7tpG8/GseOs+6w11p68lk
efl8EirQ5vVt2A+b0joxdE+jdNlRfoO5KlCipzanwaPc4VdTlAi9SZmIqORUrt5y
+arWBVnZLw+fH0zqqlSTc86DXYODtuYKlU7kzuYI3maibZldpCQtADUg4PPHuLGW
zFIGoCGGtAqmsJqLiwn/8Fk78lSl1L0PeUHjtIMv46iDbhyK9xmuWdFf84WAwT0K
CwfQkUUnlW21rD71Ex1uhMJS8n1clP6SNHjip4AWThVdr4TatPDhl4tyvcUsrRjB
/6aDeJgwYle3SVy1kbFHbofb8R0pcR54mUBegUFo5fUU72jQRKoDOrjsDys+Pppq
9bzgWNDNxCJ9PvUCaiNYmeDoZ6FCXG3VaNAR+3eyqC/ENM/mUyt20y0TdoySo6j8
ZnF96E/kVYW+TJa14Z3sgG7/90IpM5I9VyfYXGNGEj7+T5EuLWoGakKLWsttsr0P
KU5lxltvuPamAJsoPcJ1pUoylD/Cr1Fnw/xpLszdBV4chyIGAwoeHoMnVy8sEg6X
vJ1Je4X8Zy4eCRlNdtbYlifCYe/m53j92aURTLtqt8xjMT+3Hz7LgFdBka0oRhy1
kDYRS+TjBNh9E/Fd3kPcvGgeMXmJ6LniFeQkVY+jtKurd+Hb+FiNjC4e55pHqJ55
aJoYj9SzQ58p29zaHXfSVH7ZBX+Rp7Sy+uTvr2jiVmly+EB/Rkz/T9QPhA3tM41A
Gtk7H5c6Q8uhw7CtQJOaHjR7UEN4tg8BkduD6XNEZJKQPJUi3WpzZm7YIZvQEiMV
kZAC0o/p11vfq32TfBekwiCd/xk3oX9yncuzyQE3dJcckFuhb0Zo8sOar9srK79G
FkWtqKgZCDxts9+fbEY/ukFfjAY1Y4nCs3vPBCSZHGhiaNJlKtPNNoEUv66XfV+E
drSHeTvGlS8x9fCiu0ADGnVKbNOdu4S2s/qK8l2qg8Ty0RNcqjNXRs5iRH5NhCk0
hNOJzBAVpWL+phWjj2vuvAsWQqLyHDTc/jF4z3uFttGHy21YgXZvCwCzP2dTnGdi
xiE8mt48Od+uuzE4L3dGgjEc4UQSdnhv+CSz3uk6mkLF8oLagYD2BxXdOB8zPV+I
+aeWN5uIMfr43zuZddi1MFCDLC1wirkeYh3HxJambBpwqN7aQl9tKf7t4JULt21S
IN/olfBz2z9XCJdwSo+fK7ZoIaqsDbEPfRFqR1k8fPOYBd7tPQW4dPoJmilHnKB8
B5UrDSyODYrFdDCOqgoWDC2nABWuE5NIZQn/LM59Stj0eVlXs9jgosFn6vUF+cQ+
JYA4XnGGXtAQPOwtokRyMazIZxEbsoA7ybzpo3RIy+iNZp553QxQvi/CdNxkw8JD
5zgXTeZ9PfIM+JwzBxq2XrlZjgN5AZIyXCvbAM2TJu/CXyUJYiFJW3rHsSAaVoc0
yYYVp7T8Yi8DiHrjk/MqAO1ArgRXaG1imHITOn2J0gdIK0m/z/o3wg4Kn+B/MsNE
49ImeSQfQ4L9g8c4mRXRSYw4njhvuw4wtY6ujp0tLwgFFWP88CiWLcMa85JLuJDf
SCcz5CZUuEdNfQWpIMdNnWJa5FnFpHf1qsn40IvpwRuCEfrA4cDUOnj1OPdH1RoF
2fJv1+cOTa/nO0oL5nI3HL11f9GQPtey6fVPfwL0rWXYEwX4w00muK1UPmKg80FG
0bx48Ap4uXjO5OqTSt/g73hnj98om9GqJfGKLLln7ALGLqmfAhsR8DV1khzCnpUl
BLlzI0T1ZlcoLAGCg4quKXzLHfJq0COOTSAjkwk46WTdR2nWBiO45FCpDNvKUY6/
wQihbengSPxZljebssQbEI151O0E7TGkVtcbsM+CYcqi741ds6WiTAX+bHq0Bwic
3cUkclCiS8Im21RjenFqhXBWM0uaRg/r7W9VV5HUxivmvdUBVBaTc1g/t+szah1g
njc1qsLbTKXtUvm1FDm7ulAx+MlUc46pGZsgeKmwYOSXoejZ7AeDmjOG5OfnCVDH
eArdNy7cJ3XZ9WN+nBXe3RhTg9eWWa1S7zxJyWRK6wBgrYgzheQgmRUcj8Qol1Cd
c/WsY7uThks1Op9rNKqeVD/ODXSVxkjFJmMPNRSQO1lSZ5/RHEUYQC/z43lWegW6
T7ustVJSNE/wj0ng1usNh7mM/PJOh5GhTsXrMH9VYEnW9Btf3ojkYb+f6m7fsBS9
JrYOt/N1MqCG6PpstkmrLFWZ7EyHJ4UWr8E+g6Ro0KHROyuX8zuVJkrlZPwVb35s
00kNo8u3gtYOttAyZDzyPily7qirLOgfWv4Soh1X0CLzYUOKETxBgT5iXALB4pqj
D0uHUgs4Eyaa1UbMZuDElwdoXn7vA4edc69H9V0F76GPIq08iBn2Kbz45dojnsCe
pVwqTavg4aJB2XgFCovSg+nxasKKKHlM3h8Lkt5z3VHAxEyK4ce0gVtoFx7T4oa9
SrXmsI9M5kx68MaOHdy+Zy4+0HTR6SpWgzKFqoBPwXIbmpljEDpWxrYvKTGds5l6
9aG40/W3BlQIdTiZFXUs4Zfv+gMlaLLfcswZ2mCkXPZmyHZuy9nU8HkQfwpC8pI5
3dTN4su3us7IzGBeFzKlC/y3ORObOx8oMr8QsQHd3Ljn/nEIiA8zVpkaPNbmugo9
VfjMW+Zw5RZNL2zd9cqTAYl5iiRH8HDyHf2TvNEKtUok92ArlTw/GS/5YM03CdWh
kb5AdReCz/mpJCSUJhX7M8mBlzaJI7x/Bt8V+VYDIr8MQrp61ehiroQfdJKnQC4Q
jMFAg16GnSGKQePKNaew0XDWLuNQbva1htMUMk1kkNQ0MxQC9DwH1eJxWetlUbfW
EF5iui+J4tqXM3QAtHrPFBDRCjX0nFkPErReQCZzLVnvualLzqfBRY5qFLBj4+nv
zTv1HrzOe9AYVvZMSvXeIaIWjGtX4lm09T0hB25FWTNu0YNEGfA+opW7sck8+DRe
TqkQkr55Rxry4nFtQeyEpbkCgKc9gJ73j/nCxEPGfMojccEBrVp6e7s6G3J8rAEP
QgP6BhcH95dZ7OUszkwImM7xER8opI/ildBoII9mPmT8YLHjFYUm6xYDTc7gbDWl
hR1nxYtzHXsNbjDVu/L+266PyKF0yc218uXb6eCLuePLovDEeNrLUOIwb1LC8sJn
2GQyPBadTspctalYu20/GWaS3ANx7x64bXtGZPVHM42G9R1CcBdsTSdpjY9EgU/v
dt9IVy3d2+gzVN7I4Pkf/jt9itQlyc+47/Ih/T1xVsF2kHKBPuc568WLJXOeoduo
X1m/cVwNM4fnRad2po2SgB3vrUuH5U3M0ydgtWQKu/7ZZwx7/YmyolyNDaIjme2L
ZFsuF9CcULtbzYhjX5AhinJHww23V7foG2LKCkufkHXoEFp3ytX/ScdT8FEa2aDs
P3dvGCZVn/3T0i7RJFaTOKUQZQSJCf5hXJm98anttiU03kgERSS+I+3pDV59Ypuf
s75EfAmqA0ZTzo4Co4CKKbPmMwl5ILCRqWGdxL5eFjDgmryLNdgCX3aGTZSWRy3c
hrgFafl5OaQtcp+2RlSkiMXeT55InznqzNr3ClXhEgOebTFYafMCYiYH1+QTfixH
PE1HfPxCqXhiis4dsN94Jm/gkqJQDmFkjxgLiXL9kFd0SOBtv0vn+Q9+0S51qCt1
y00BYotLneQ183Ml2UgmrJkeSmLkjgUBJyMvfTO0keJ9UybDk5zm7hm1FR9rPwGm
X2hmzGDC94m1FsKm6VgTkVBj1BvuJEOnqMkOu8+ryDWd9BBuUBGTopmt1PQh6Yea
CZ1baK//PJiRcPF/GB7Zm0nE7DuolOurus11EBXK/v0LkpPsOLCHrb2hE3IIixKi
Fl381JjQshqRDMvZMC7hPriEUrRuemnl/GYkaJ4PJe/l8KDwTCE6YU8F1qTSOrXQ
6olbNrDj8VE8y13fmD2ILdGPrxrwzVOo1iJkFnV5059Wcd7eVNQm032wVYd2Cvtd
nGMeduFcQzk2qvynR7uHq4bo9e8erhuEEHxMHbjkyCvAv0w703+CSbfjMN1DY9JX
/mB2+NaeoYakTU3hGg5mxpUcOqtqHCJouQBoWIfWfjW1eo/ntaQmEYJtg3lSnR0R
oU1ud6jmRrZNPynqW2QoVuQRczzFQfydXzzCzzMNy0twgxqnHUU2N70wrUQCfCBw
Nh/+gGb4TSYmsrUnfJdRutUfBVtqaCJpHzWtdLqwxWN5+0fCsq2qMNP43yGzGNWk
kqKyUCrx61L8v520woSYjy9yCcemoZ2k+CUYepOt2Du3+FXZQ8za2MdvbS/vqR8s
Gm8ZrBSGQP2eNw1cNfjbBi0E3XKEClAaCBFaHsHW/yLpAUmwGIbekzJdgE/VdAur
rmTk1pNjBKXzPHjdH1y+NbIjmZnL2cQQ4DevAHkjGYQrrkMYaiq25V23v5LQZ1KO
qPloaWRTU/gWuVrvgNOIIWvdn6n8068uMYEW51qgcVrtecB8CQVL2nrJIdTZwJuz
2GtVx4lZ+ykSkyybi60YEEUWT9iTmZ2RGhDpc5icyf3qOWMCYFRfnNB2ysyj7Gid
NzSUvusMYCUBRbppzTXlGzDvUs1lMHJi5xLMmsaQG1tWZDI7hqwng8yQVhkbUtvJ
5s9ItsJwNOnnMlG4EpFXqpCZa3LT5UIq66ui0oT3bUaZe6kdS4+UhEfH9k+lPf2Q
karCFKgdoNbf/h10yd4fDIeXkSRhgivKi+xJwXtTLfhuozQhC1qRm3Cd4ZdIwBEr
NIR8JCF89BaQ0wAPuYOnt03My+T+Pg+l66HQdXLZVBFNScJv9ErrXWQfQjEvmToH
Rq90mozj6H+HlYgFsRZb+Z6DHN4E4sZHXbeEZTzo9rQZ01j0XpCzd9UtUwY1Nkpu
oZgkmoyvNd2vkIxpkuVKCxzeSiCky6ttX3Na2vhARUsAWfD4v3XqSkivPox9zymB
+ESHAmU0rZQLh9OfEHJkVftc1m1mlkAputTHYYNQlHFkiFArj93WfIuIt3TfBR1h
9TyDzJFTXRMTLEuo5vepm2+CCGX0YQ+Bic4CpGTJmO6yrxbWGy3+1z4fSotsLgM0
optLN+5NW3cc1amWFQacIpK3nKzL9VsDxzFR1I5IEmLOGQ6tPmA9d6UNZZimBuKe
NukyN4SpgDJmlJHA0ruqZ7nJZzPZwxQBc6liK7ajB/JYB/TU3JesT37vNpZkCfl5
kIqnIf70sGh2myUNrvzLwfb+3ZaoF3PInxViJVPiBHtRk+pfTk3e5S8jOQ8YzCTL
Pk7HM7I5cD9q6Zh+c15NHjK4z52sfHyfrRWD4X6QLnn+0Rh0Nmg6oZxIhXeLSBGW
krELmynqJ9pfj0F2TjoiyF5x/PNy7WNF/jLOCvFRNSqZucCY7o7HlNCqxiFR3GmP
e2+OdUb+KMyO0iQr3hBY0/Zoibjwv0YwFAQyG60dFfX1PY9G0XQ6eDAtaAWVPUm8
c+uy6Pt5VKhi70AvBj92Jy7wCACFFD+CGWhdkeJ0y1xhL7n7X1+Um/9P2OD7J14f
o+XN7ahiOflF2ed3HhuNWBJTZD4UkalV2cq6lFYzNPAgsEzQGUSFmLlb8DcV5CMP
MpD3jvUmB93BVCt2LLGP8avARk5QCdsDkzDHyf/0SQYFExplo30fAFrZzoZo6/eL
4LeSNisapLhSLuZ+DbxQOM8xrenoCz0mX8CiTZJU5XrIaL9M1haYMaC+s9iRbL/B
TUQBe4BisQvgHwEvrTl0+KIYVwwIdPrSJI9qfxzvDuR6pd0zcFZYppGGsH/fbDjK
UAocz85hQeoA/UvOmA8xh+PxE6kBa+iwH4fgLK3svKCBhvv6ZTaScb61Ii+IHEGc
l6Llwo9K6GZ620mQUd7Fcqy3upO3SZe1nowcxhg/kTEZ8dSdraB+Hf34WosOru4J
pqHuMT+OPaEA7KdHguDYlkp6phhRHoij6NdWWJmdzZxPum3vzlX5yv7pVB1hU4Al
BZNZBc8UVldXPECycM8BoOzp0ErjbvSfTXMYxievpAIaDBZRMUMNWtImAhW9Lgc6
xAAfXTgUEZ1RY9TGs0ssIfmdFj9lY9kEvoiUAi0HL5e5OO8byVMezHzJqRBvR+Ac
MzSBLPG1tZambGLQ+HfzDIpAHdKw5hd+kv2VQxE9GfAps2mc04w830+AJLxP1u5a
v1y8GU/8cOFQ+YxQ6AcqaCsIVi9gp7zmgCllB5SJm0aNF9CtBtcaXwaQkhOkY0xg
PxqaPEQtprmnaVAZVdN37et22ZxJp3XrWDF9xKcvcY9DkbL1QEvJHY3GInggTgY3
IOZka7PYaTktsDgMcV2dZS6kR+L2RyjBkqogeTVLkGFgJDqpFpxjzIYohHfS7FZ0
ECSc+q5K4HcW6LIEgFVWTeUaP6c1trAflnDHoYBrkpcH7GlH51rIgVFmxw6UUNor
DG8RzACSCdWG10VsAEsQJ48jV+VStEICJeCc/haOwof1CVGL3bDJhzF9T65fMjFM
sCXXpfFI+xtOjZwsx2GSgosci9kMRt1ezfEwxOmxQzyFzaIItCmEoaDP2+92s7N6
0GHG9repo3B62wL9v5mLqGWJq9sYS+40ufklWNTfHfow0zuQyqSr1l3riw2sfxWA
xUAiPpE7UU9ugLvdyovOpBaLJnK+K4eZC1DWvDM8tHWlSYCftYDHbjBaG0U4GrrU
UYoYdVaTqc12HxLntoYipZWgTHhkyeIqHT3F6YhTYzlPWmvIwhngPzBoiovOcyuc
Im++stpxEed/cqzTHwD9+xSzz8+sP684RX5IBRDYxZ8MqPDQLIQGAFxlMpfqOhL6
6H7cE4z/EV7BoxhwtIIxxvR8mCh0s3eCEReBOlFx/7j7xj6DMQFmCBN7ldOs+HCQ
PDZvsUkRvP6f4JF+qx0CSxVmW+Emy3/MB1RBmj6lI0ynrDx5hB4qb6KfXM0JkqAq
1wWfrzTWhIAJfWzbXZDO8EUmIQ0ezmyk7CdxtuxVH1d2ooCSZ3Xi3eowOS+4YeP3
u2vPnzyYWJC2tCEn5P66UviC8Guv7j/C7YfNVc/ZXD0FQWxb84Z3kY9uFBAZXSiJ
KxtjwPg1Ut5BrkNTuuWokblKT/4a1fBdxytB/7dRFwHtpLMxaEbrIAh2BeFHvb+d
p7v9cj5eWKszD5IYYE59D13tYHvi0m0h5aL3Fo+e6B8JEFkFEgP4gKCCM8djUdlB
bWD6DJOWR0XTOD6XeIjblOP3zk7WHzhVdL9miXfTp/5ZVEWSaA4gGIMLgys+VnSB
8J55Yw22/eTmBoVjGnG+p/uZB/5Ly/Rvs/xNl5xuduvUEglyaRFLRcJpcwwX66Aw
jMGoB+zHDfVNHMoAxGaypmXWCvoHhKmgle3v8mhU94YNlFvSGznHo4I9UGDZ/IzI
QBwgA6mS2GQREV+TEozJ+xnjmiXW7TJxBDR7QGiGTV6yFeJEvzQyJ2aoLttNKRhN
O0YyWP9Czs/c2yjyLd9nid8X8Zr5FSLwgEIERttqsxdDNRPrmBs58vWK8b871820
j9IxXvUUF9whjFoVeRd5xE1VrclBLgyHGR1Xajcgy6UT79DZJ49mqTAPFOb1Ijy4
n7mGxQuubmYrkC1r7ZEWPSfAksqaiGulYcEH7Y/MBOsIIMzXE9RmTCsZFjSfm7QZ
WBkDaYyjydCv9+cclJfezjLnH2FBDcsM8l5ybGScGf6o9TOYzupUVE0atxAhkBBz
D/Ert8VunxVex9tGaA9qKxHvymoQ/jXpHF0o9mTcvdqVlMnXmtgDe+Nbv8z9fcwh
mJxk4IkKp5uaMaWtNNepX/5wWsMHy8kW2SuSt592i2RYB8MWrCr/kRv7G2g72l87
XmlcjhCMP1eVVgkqkzRf7t5D2yWEgDnQh29TEfF8A/OJkNyDdcqJ0hnspgVUo4xr
JER+6fgQZvu3HEPz5U1iV5bXCbSsDB7KraRnsHanMRxuyGzsDelCELIky04lobQR
FVQOHXCdcfpaUBok+uYTkPa0BHh2zbqpvFJVlcKhfWBm+lNK5MiLf2ZQOSFYBppd
9oGqkm+s/4IdAQu3lhvKTliTJBAPXigwBx3I/bMwXjPwwtKdmhiWUF6qzLKcsIEe
MSG74GTBhj+wIVEFsgahfcag2y3AbuCsmDu5f5BpmLNZk3mKXjMg6GQ7WjjKfznk
XcsO4KvJ5Ce55MbfbtgCy0EagwTGZ6QgoDurJGLTSyxxqaMXv6irePyK92sOS09H
/hgnrjz28Qys0V/GalFwHm5H+35I70iB0cOBXgpUVwjEq3EpcuCheA3gbfCp8PLF
TbOCAuxM2S+1qFeUPepXfLuphDBsPseXCHunVFsdhGzEc5NUiQM083geFysoHGSt
Ldl1FZ1IX3fn9MlJwH1T8EZDDhPv5bbhTy9ZhqXjDhlF/K0YDE86d9GGJVJLAkW7
V6xsMmpefYzyBIKavHG+tyOspAgtfZT48TR0dbxq2PM1lTYfw3wTVH6ynNLdL7PR
tTsiPvrOO3kYv+m4F4yCc3DrvH3UWtcWBnQBIxaLAIHBZBiW/Xfff4R+BWKyahaS
oKzWPCwbSHcNrIwlcFtPZxypyuFKtbV+9MyJ+xxhrWwbjCd5Ps5l8JU8zDPabA2M
nfoTHj64nIZILuO4bEiZOBTLbel3B+GF3PVstBR/7HHzh/93XGHzGH6yxhNrsyFp
c3DeNuxnHpQbW/vYDlI4W1IVbN4QM0vevQNZ4cMXfi083VPHRHW/Njn4ULYVJ5zq
z37IHgNpN4ioIOxSNqZR6LOQt6fGxpaXfHaEu5ynGCSlgSXtQ56Xyc9uO0B/+6F5
ZNTW5CtvOrTzk65ELhLK3OMNsP3vuKOjK9L7aADJZl2BB27epzCs6Y0DriD7haKr
F/88I19wwGMOpuXyHebgp7FDW2CKvX1DD/wKNnvTpDept6I4XTU5LujEHlL2FpqU
nqFvYoWuxW40VY8xmSRL5z6sM6aPM9xkNkapHssm4KcPJHoTxvG16hmVGZ+ya3Yr
4/+yvKoZWqD3HIlf9Bi77GcLYhXoDdPt8cnkwzULFBAS64+Yty2xsWyDAFeOlPK2
MucUGc3Bj+tRc957WMj2LyfZsRnsV0tbF7zgWybZNw6RGpZR4fJd4VKeWKhj90z0
q3sl7EXliOUFNl94pLHefW4huoW8LCCga+Bp4kSWd5b+nFiaVi3/7olFKu5hZpD5
MBesdsPYdOBidsX2Xy1vpAPI3Xo9H87NqlGKyVJb2HxrWt6EUSQ5VypUMwL7G/IO
NL9bxX2Sf0hCIi/kZApRDFLCfRQucCQ7W2ZyuDpUdqf9iIdyrEOBfVoc6guKog6E
iYcL1M6iKhIg4T8bzD8BiuSfoQkFxqV0SGyaCinSN8dYMrSpPvviDuFdModIYBld
oVFDosIr0Kd3KHM7bl5GqKdVw7DQci3WZBHvwhmogXSDfqrfvDE4+CXTHSzZxh1c
xpBxV/Wl6Qzoc4BsSlZZFSLhmb0UxnEtQMbGCYlrZy4YTlmVruQzsXNaJzlJbTxn
5NTpYw12JKXqcKtU6uaxPsU4mkvGDPO12ghyawjYCJpMOxtneQLH80NUAy7g49MA
2cC/YqvjboGyZ10ooHU37XhoEKmfEmbZ5YRZe23/V4h1XQn8L9uYox3DfYNGGpTO
r9k5vw22/3O9Brk9YK1u1PjdN0WWFx2O94MjZJe1tE3qpIIknZr9fOKUCFuo/BTg
t4h7C2WFDYn4KmC9bASZdarbk1aNRMOyYypPdkrWjI8IVd5iQa+EBCjPneafCyfD
OMbNslJmG77wNxvc8JSyWU4zVYdX6O5n4qTipS+QZ1PZ5qhg5Xbf9Ckh6NSBcDmE
OrDzx9e2E3Ml7FEli3HtCGtHSIY1hccRrCqywhun3mkUbV+2S551QXRw0zUWzJcY
Pc2sQhQYJR+NcIxqPpH0gg8CZOe5BLP1YzyL5NonlW/KlO2c7V3mm5b1hTJaMVFZ
k/ktof1O26ZvTmTSz9S+kj/RsZMcrCOeVzfSpY9LcZu1hWtIlSdaNavhh+CrcmES
qWfizLMcNDd4wLVCp0sTDgbg9F4xBzFerUTKp0hLf9F31byEjFOMTVuFyfJCfQ0D
ACs6cUaF0NyggN9uSIUlLtf9GBcHWkDZjSHj1b6oEa1BnFHD4xr7HyQ2Foghu2cc
2lz289Pc+v70jJJZUnFCFiX+oB3HJrGfUd4UkGBgvvWicPQk3tibDjy0z8gHCb5B
e+8vTk3SJuyAAv7kj+NKeDQF49v/F0xzlcLhk3dUYkYi+i20VMoJ5ISlCp/KOXYX
iqzwIxGDsB6dGV+6UdmElM/EMsNeaEgoQ2MH0emUVZvG6H2xe/ev8C1VIsFIAkMe
65Nf/wt8wZQjtjNqaIBrzk/xNQEP7dHbraHwVqVeSvgCEjzz0ic2AJuui84XJPP4
4gGB0OoyFk/syF/bYDQKIRa+0JycuxTWcOeX2Qv1xOJK99ClP1W7QlcyJ/xQqhgt
/7a526DXJxRQmNXhnB3EpnwFawkJQNBqo6s3W29QnpnrRrRa6W+3OlAG3TRQwCfB
Rxx/UjkUBNG0DEcG5p1Z8akoxGzUnowkycO0UESiw7mX3QvOz4ryUUMI0NyxDfjx
762b5bUuKYkBm97+bsXCv4c9o4x3SP61+Y9sp80H/j5FfvLrRSE0lUryukVU0JxS
oEACpYM8rylCs8vv1ha2rPB+qBgJ3IV4PN64x5xz/qWOuRwSTxWXZwBQiRwdyf5F
TXGYDd4+0OtnxRokAvBRGphkdJ4l+OMU5g/fbksfPkViKf7hgWeRSr+2HczRzgcN
jNDtquMlUrM6nY2ekwRUZFH6/gzFep6mkU9quNnx9FHe4L0Dau8R/bPHF0+tuWu7
tQll1T2gusY84aEmXnYQAxwH29gD20G6j5njDCV5hIe6ieaoc/GD5N1rNCToBYqA
uc6JFLKIYO5kJmA+4SjJFuPAVnfpaR8WBkPKOu1rG+AU21ii7BXZ5MWtd6y9VNS4
WXtt9+jRo6DO1fqDaVdpDajsDdZjLmIj5q+n/pYeXzpbGZrDsswayQxYBn4sgVVT
YumsZHbdkcsadTvRXTEWcd5Jn604/UlNs7t+wjOhMKLyAKFurSM+Qm8pfc+YS0mj
+y8np+OHxSAvqPpty1QeKuBMCm2+PXqFh22GxaBXXvs3qU4gtGvRi0su15Xn1Krh
AcS9x0cqImW9zQlAPrio9F/VCkrKJ37c+A/+nS2D48QZkwI3H+pDdXedRiQibJLA
3CjqJY1vBAAp7t0esXFHpPiaAgTLeccdv8OOXw4iOBIju6E+LLlcLYuWpmWLwDFc
U/raklJcm422RuAOGD+5iBkOD3EK18hvHAjGLBbX+TY/xc5NAKssOZN7bF4p+Y19
9mu1DR8s2v0nQMk2nxlK+qvUJTfj15MMfx+oehr4FayJ/yopyZfHqQPumjKfIX6v
PqYEzjX5Ssowv5sK+eHWKq2ehO9y1VzrQ/lrz1zGIIqV3nNBMXufsE/UsQuxxff9
Rrg8OBaw/10ZGMMARJ46KRY+vB3XgI/xhqBSRx/JLLWuuR4ksZYD7S55iamJyFY1
Xm6oAP1MVuXF4YAu+SxTz9DvI+fjwOxJemyHH3FWQ8a68WWTbt8cEW7WecU7ZVma
L83xQUv+hIJQ4eG2DjrOkwaRQ0nuyWcQAgcLcpiv6OubmXpnQsVp5IZiHkmqZLIu
2Q12U9Uh791/VJAh+a7+LSC6gTr0DniKNZvD1a4NfkIRyO6dFO8hrMNY+DzL4izZ
XAVjXP5XUZ8Yy02E+dKE+LjwEZ72hsw0TIV1P7HsD9q1eCarnvmlGcmpkP1i2Z3I
36Gel1hk7vzEOdUStq+sWQqRl1lTr9hfSuoO2SQHWRJi0BVjqUVmncZs9yYIsTcC
fMlSm4GUgNcUr5AjFTBqqE8BeS3+Az0XtJnbnJK5UltI3JNRP9jrW/WccF0gYGKf
so+v5WHxRn1/WxVfGLK3jJAR3jryaTnY/1TMl7U82KPT0ZLRT6icUBXY+FouqLwp
5rDyPyH7Yqts8Bnd/WnOMpuQQhRZUBmsPqz/DKM6D9V6fRnJ5H4/akUuZ1abMEwL
uHEtzfwcVkK6w4SCPJL549Kcm/KkM60zqvJDwgqZdel7dUsFbYWMKVPhA2w7RV2w
aQbJH5lOIf/5DPXEXzQ5krKgl9DLA8wJiJxMv2wIlC0k9kX5l1i568kKFB7w4VQD
Xc4Btvrh5E+Yr7DoqLE3OJ2bd73LQBoeuOJlxEBZgEA0+90HTtg7aUZmDIsYKH1K
alxXScEVdHcJcWzK53RXKgq3xfq9dxCHOyhaRDQiznwoO2aQe858qkITCWoCIGAD
LC7CeLS6V/QIM4NRSBqTnImm04Deu4oiFwu8HIRSqWB36EiZw6vaY9fGPTf+t79b
n+BJM5vrvdW6Qb8QgmsauWvJ4Y2NE+/JuD+L2Ke8IY+xl5mvjixDYOQbUyt9n0C4
zf1e3soCX+PkUvHTw1hcd+pY0NfiBBTvxjpS5Q9j0lbSOWn9eFikmqfRZymybuL4
usTxHx/L0XwNtD+55jMxkdfNHbwpvDviCkgGQ6atQVsL7mzIm0Mw9veqC3TyKOJG
vs8GfyxafsaAfmClTJARKiDcXve3lo2wdjaQJ6Cu2ASJ1ueHcCCTNejfATkfxupX
DPWApHl+8gpSozjLjVABeTIkBHBpOn6k0L5hczRVwLe9wlXBLB5YM2CiG2I9SpLu
tfwyVqFKkaUtNjoPA+6Lujx7/ZQbccqr3+mDRlCiCDQCCowuML3SDckjbiyx6kN+
UlpcChgXqqoSnIxJN5xgTHAY4JUI66BfFhjGxPklDpOZNnAUsE1TGvY5cQamQn+5
YHVuHq9nNN96hQFc4RVBlfC1jJwgVP6TWbt+qpx1k+/vAbgzThgWLA5631vHQs1y
/Y3XMgan6YJSt3x5W9Nfx+j+Q5yYoPBGThU/P1n7kcMNLPIRwrQwHUEqsela/YR0
xpu4AyEIpWlyDx29e7/Er716gOfa4HBOL0kctm2uNMg/LYtntwLedreE3HikKdKR
unnPKDG7fLNPgJYspo2R8yKNw4QfhHUju/onuYd+lH1ye+B3WzAIDFwZf835ZULc
88Y1ryEky9tGn9qRAgXrhvpZxmLsVo5DBvYYGLRi08tdfWSsQ9VTbB6NMFxo8NdU
ys/cADYzuteM3fUjVg157cplMIaonp8GTQ0h2nikm3kXohMnQ9Xu+ZMDk8Hm1upp
CQMl9sbz+O4PDgP0nv8mQVZgFNe52YFHyGjlUG/w1K0C3w5XsovD0INsLBuLUhun
jd5WN0E+CYoTmHMNnrXpbiTUeRUrNfbBteEkdm4/IASaQQxCWOW5JvyKV4B3VoMN
Vn3H9QB9vwXy5apRZT0Ux5+zKSD1Tpz8EQhRq2DV0n8sFj6npKB7R0nh9ZffEfUx
T38MigP5goDvGd9KHR8GgraxPQS9ZE0kycHJFoa3KasUVYHcmy/xQlSWYfVQzTRY
bsbTeI9x07piiv77rOrkcT2eCUufDj8Xv9Ilj1Z/EFDjQEbEdP7gKHU1VELAICt8
fJkEBZySppOZ5Kz0hMi/D5oDNIG+tKA/A5KV3WBnhEraPy9Z2Ett0AYyz9VQCGoh
z0Hp1wYgyIOmn98xdm7739eQMqZOoTeeoeV6ipDGDLVJ5X4ClCkFd4wFj7/rZEmD
UL8Q3Vtn2YQHO0PSbiqk2CyQrVTqusNyMgbQX4r/58FbQZsqQ23UpTkD/jhFkNaU
q99j1f/TV6cGFWVFDWuwp7Ofa+ZCSo5WhiiRKpsEuhollW6oqHyWtseUillrcc1Q
qsHugjw0kd3F4TmVworCGza/ZHDitqPth4/WHJvkizeTUVyn9wCn8UR9NbQAi32z
E2t8UDXxiP+yoM4RgnyVXF1rpiKpZZ4wBC2+vr/YH5IFzSASH5zTFmOUmyCclIT+
XtGAWj15eRKzKtTlI5gaOQUnzqBA7J5ag2GfsCv//sfJNc9TnTFhi3LUbaPody1d
oPb2+5hSIYhidPJvGms573JIOiD8x0DR/n+jaedErg0o9P/RTEoD+QrcDNwLpUUt
waBRiIpQMnSDiZFhgkzsDR9qNmebYfOwEP1UaH/YiSI7HUTiPunGBNpjiAr/Bxwn
OWNXalCIrNdrVuqnoO5/fPQOB+NBF0r707I2xaHXpoOnYWdirxN08cd/0KVryDFr
oeDhUZr58wp9UyoN2ro6ZuPLnEJQ5O9y1ruL7UIDvrzWNEapoH2zGrFAXyTg4a4+
7zxc/xc4+WKq30HGz08CtwQMAQPBBAZHhim27FPIXmA8q82LEr7UXr4LvzDzOWD3
qrqF5ZWnkKHsUN9mjt484Jrynuw9l0b8NQ9kgx7lH0L3MX8GV6vd9OooJBx/jzFU
ORyviSMHeeYVxN1wZ09MYIm0qI37Cs3LS2AuszM+UP+GDbIC6aJo2r7Xk9DvAoCv
Kb2QEhoAfI6eY5+EXnKydOo7pwt+GjUWfwkYOXRQmHUL2DwSHUDFx7333fg2y7Rv
TP4WgM8VY8tGoj7OpjbrxKpBKihzKIfjDt/2qW2n2FtL5JcFwAWgmcXyb4Y3fMcO
EYg/2cXRhQ4rYOisordS38o2gwVYTkW8sRpARNdr1tb5/K3FwHJ1nUzSLFwFjQ2/
D24kfl4WJM83CNJfpDuP37c+ZwkARpx+2qzwvqFJJkhmzS2C/TJubdD2YuXP7/fj
YpqKsJIjexbunCqVstmgC929blSme8hjU6XDfjIxpb5rwEiD1HA0cidU7aEQIc98
vAYZSrDVEoQYv99CHUnf8cCdU0A3ZNdrivIgoUFdcr/8/5XiX7eM2iLkyF9XVIWk
5NY0pGzfZe7cAIdQqonrEABaFQHO6DlJeI5nDKyXILsj7/FDmW8rMuc0cJIj53NP
KWdDJq21qNQo+cpOA2YG+/7Eh6eNnXl9Bhxk/9taeP+2/wP+xTehNBCofX0VT9lU
uVs6X8hMFtfzzfRN8CZT1cBoSCQFqlT/hXFU/kyujNrs5DJ6ZNywQ0IYi0ZdKM0G
o4AE+QoNt2AyzYYj6R0RExKLgign6VfN4T4toquZHSnL7GuvLbBU8c5gPSndqCsT
4FXy9zxTPbXuslYYSEPRcZXbWXRZ0kKwADEZnivdBQjzVoO7irSFcZtLYN0hCe8n
jWUB4yhzG2EZ9Jt9ltLcrNNYnc4Sc+QcD5ECC70IpnCIuJfc7N+Oaxdmbvz+MZw3
ynVSlMMXhQD4HNyZao6Qz+90eUv1XpDMY6yq1PdD4KrsGtC0WUnxz3Ny7MkoiTSq
6zu+JBQFQ1VyiTRo/OqA74KJpGHIjkV414fedQacrb+vAg9zX9Ieh9LvEUFXAEdi
PX/GshEjWLIlED6boTaUmiE0QVuFNfnByAphwOU1idSUehwBGgV2lklb58y1kL0F
vgwFvBLmEU0kUrVVnaaGMZC4b8x1M0BZ8CikQcWQjDt6qT4z9X5wluOP4scjxdkp
TWpjrqMFcAyE0qt5kkivWQMJyju+GnwJ6DrDLcdxtVPCRScxSV1rDJyweqVbRYeI
fkJaIj4xAjQfagAUpfDP3Q0KrzJES6G0ijyJZ7qriFdiF/ow1qUexlx6r9wlLZXE
QDjI+H5f3iL7UJnHGE+SZ+VenOnTcp0vRDJ+02QrzIbh4tUGtSANxxNvDRoJA+Z8
+R6D7+P1MfMJZXkNBQBQ5rxwEqagqj33MQRxkIcfbUx5h8DujufI4l6PyEyhb4yV
7wWCD5cKzp+84taAD8PicrC/j4jo8wCG8DGeBKnR2q+Y1UdYiabCnLm2hnm+3NEQ
VyI8EZ5tUzn9jzFSxuCJVvWe3k4HTxk6vLc4ib0/6oP5bt2QInSYRLGBDIplxmoL
7KyBlWMkW/3yIqSSG3GePHSGQERLfAyEDt4zRC4ywrV0wpT47wQpEulCV3nRYlBN
zjY+D0cF2SS9E3DdjPNrKt9vzOkT329BA8B1/+wLSHybf9Z+Aw8ksLfArzLL130J
Z9HYGT8EHgWzIP1eYfQhKxRU8fvUcK6mYNBYCAp9Tj05VB+SqFJXK6Npg/MOoxbi
FeALEmBELAkdzO25na6HY4HW4rKCAtEyzaZD2eojCAuatzfy28chiejDWK+64/wH
7ogGATd/tj8Bli40XLBbK7UdvG2Q2OP39ZokCvsg00ibOzGHj2A/PDMv/wpo/SuV
Mu5qCNtAHKgk/E1QAURrYxjNzRqzB4qDo0BEbq06zjcX0bSOnYY+kVJ8+ZQ5uaLL
p7dvrBzQrSFB3cB+vECegnwJz9I3VQP6rX8pLTbDrW2vET5ONlbrkuipZscN1C/8
waVgCmvYNcHWgcfCWxShepl6/HAqBTaWm5cQ8Q0eaF9kmrZ5FccLv0mJaaQh9eXg
FTtfZ6bvShiTUvnnX+WryS65hrPlkdyl2dFTfDQFmVGrhx983VrAtWz/1uNzx8I4
Mgqw3on//oZdrchUP6eWtDG0dzeRjbosx0ULsg8dETpeeKrujYWBDNFoyAwaKwxF
Q4UXUTslDBUNqGtnlSbCU/Gaj4r9NE1Kg4WYcXI+W9TWYbs2A4XXloo0EsE8yi/y
g51SaZ/JuPI7nzRFEcaY2EHUDSX03tR4GvZW9mZnpy119rdT4Fpe6+ZbcaDNFL46
NO/F+lJjbsx8cm2B/akLFM/2vaWMuFPd5lGpTIbAZ4Wpc3L/EJd5TAOl66pnB5uu
wf+rn7Pu0H76QDwk51IylHmd350I54dVl9Fq2uMBzuyfhk3eHM7xgbf0PR6TW4jU
MoonCkolSxst6dnfQMVi8HPDWMCidaPDQ1AhZTODvGGCNwvxQpQA0NUIlZ2lNXZd
YaKdGPemhmB8W3gt/g+5s/wbgw+RE6NLHDZbdJIE6ja+rlyj1JpXwnhbCWEU5QCA
g1GpsQ+eHjaPJ61h6FJ+nN7tqLaWu1CzgLHzUB5RQQuXYlcpi7RIer6XR7lKjoSW
f/kO/5TmToZjcpRcm8YzoI3Cgl/HsYkc+pJxbQRAqRAYHKzh8ezLO8Eua05Nz6c9
WamVgSIXc1E92B4WeLdvPc16Ur5n71H67c2chQSs/3LFJ3jJ6/tlWPFneGflec9E
ei9+TKGYwuO+/AlNPdCW1cr1aaLBFxuyTKPo4Mow8aeOFn49saaYXTVfmIkxrjO/
7q4gMlow8ktXvVbYo0sN8XB3hovjhxcBtuRMvcRhJZkHxQbow7F7FXflD46jrSmZ
E37dgeT8LqtkZc2ZyylhBXFZDvTrWYoRYnLwTlLdKERcyf6rFTJD2HmZM+/3HytY
2qRrneaSFq2i8aqSukNK4NCMyWWAvs8+8I9qlHpZFCvhQzHzTyNhusQx/NKrJGyV
clHpsKDnhxje0khSFt2GliWFwNe/zNWxcunnzOLHLd6mMdBMnr7ckiCbGNb3EcQ7
ZRFjzho6I1babBWDJ4YrdF1cUvt/IwCCjrp5G1wCODOCct2fKPH3aWR8mXztIYGy
mNzQ04cxkpLe8xGE4ydjuANBvkTK4KdhcI6o7zWTxDrHrrqdrY1VhQgnbxj5WW8j
ptw8YDAr+h7uYEE/ooI6+TB4Pt9hufVZJ/RknfAcPwrZQcc15urAvzgmiNB9VfsD
NDsvNrDyRgMij2q2Y2xy04zF02mB3vlkNYEiYl2iL4TKMROWGk3ntOOlnZrtuLwu
vLPRX17huSotFgTlVJPOcf/1mzl041NaTJSzZdTqKQkKqkSjLIpm45/+1HNEnZ+T
yuc3fYuHzSTK1VPyCjDXcHNBpStkV0rpD6wSnyIgUBhcwE7ww07h7rHgZ2ig4s/M
EMGRDEwUCrnzwP10Z2jApDikRatQ6X/oI2Y/Z5p9rnu7acRojSXWh9tdzPuKZNHK
DYm2wRz5Jb0xe1+3SZfi2of4+/ff9VuRdNcIApdcLXyEJj2xOYHdhZLSLxbS8aVj
GCw4ZiyTSBSfeeF/z8W32Y6CrQAPb8G/4ofULNyQcELpDCvpZYhnHBhTgDM2w8gm
FbIEoXpMf/UWUBUwmVV8Q6HIeW6IyUIzbzAW/uOUGYK0c/MKPK89AG/7DQIy+la/
mqbevP7nKW/eJqN4AsiAHUE+RqU577U41MhzHo+xpZSoC0lXxOX3G8UMpz9ma0Il
1vCo3N11MdGrQg0rbqp/HghW/8/aJQDHCnwQKMZXCXXTuS1KssDkbcreFwNx1g7A
jJ85fRajeEl9dJpTQkTiBJPgcxICcu5nyCKeGUtOTPcumj1kq23kkCup+qEB9wR9
snTvLpjVzX768V7+0CzF7XKyXJvFYgXSeJK7VYKr1F/1YjnpK/rE+JGUb98mbVMG
5zBo7vuJUuF2DO0mYk1pMlToYwUEGQtLel9WDxh5sbDrGSvIyQ3+JtkqwnEXZtcH
HFweY4iWRdB4Wo3+85W019icZAFihCuFVXYXDjgkQkfG37FxRkE1wSMOvuL/h+ow
2BzBprrQQhOHrrKwdrEuazp0EyODO+ipxMOHqwXcPwYBn8LBPdJiudaXJjLWSV2b
lnARJavUfHSLdMdx/Iy7BC1jmqkac9ChFYZ7aIFLlrQoTwSoSAcc+DLKDSL+RJxl
vfvEWOpFweHSn9jWEsWbfUkKh8TD4Xe1y1bVeZvSKDGNkgjuR5FpJyFz0cjUWOx0
MamLIk8nCQTOnp3CmHHrHRT1N8v6Kj3LW4cxpCfe8EsI6xw0qJ5f01unOnWXHvd9
I4x5umObi4416XtPUTs1J5Cz6Zeb7goxvjANj/orVxWfj67AwyshYp8ZVVR1OnLc
c9td/KXCad+v0x/+4ysgYAz5+MiPPBWEBUKMhtj2c0KwQIvomU5Rlkph3Ed4DX47
P4oL4oH+7wAdkPT/CLQ4eXUOqAvqbZ3Plao8uUWnQaeMwhEwTbK+1opT8bWARs1z
IW34v4EaDCql0mV/754GzgYMcr7uvy7+wjPwr23NYLq/rI50wX1Kq2WmKfKvYoKo
B7qZHkLR5lvEmGUs7LqdOKbQsjY+QrYUT56vyqqBNuj37M29GQDVfd1z59bUe+qY
B6MDuwpWEBz4hFQB15Q6g++05i1YZdSfLynWBeSHa+GMraAAkni7Wt7NNvhm/vtx
lh1z4nI4Ly9LKTqMBRsdxsJWsz4ykzQDHB4pOq696/DR4hjFV1iKEiP2Jf3J6Pvl
+qh8IHZKVetbBzl/xzw8GOLj/4t6zI8w2NHvPMd+G/XkpwPl3vR8VEXmZmij9Yf4
jMlExROuBkrI+MpPKHty6tzMo5kWnLcUO+wmi11T1DvUO5j7xR7HoByx0wjERCVL
d5TtFgBtQSyBU9hEtmdXPQLnu+th81PaR2elxsbWuW7buNu5m6RyVTKnBCw7rnHH
2WjbaSvU5Fz5tD+CQ+XeDSaQOy/nsGgz56sxfUSDFSVTbWGBoTQv12tvDg8C/k0I
ePNfyv0rr4K/IJ79hT2bCxxqGNnBvMfAIv0Va+sHgrIcphi8DfjCDN5HfQXAls/Y
/eM9pc64SNnxWwVOcae0/+kdTaipMXjCthvsaFsu/dcUoOlFcsG/0C/gI003goX8
V63iaKAjRrFvRsz/R7iqz/6YToGDGIQXRuZXeefOD1ItUh90Jxeb1YfEiMDNJWOo
gqEbiF0XIHOOr8uPktqtZVFHSRM1Mmu9HYdDGpTzqoXe/PSRdH9firm5GCWy37Df
slLwr6domSziKx47Earve7gfQUP3rb4bIRc0Lx45GXcdP7GI8uDBUPCaeqySzVpi
vgmOMHMS/JPGoCc8TcwJSPkn6dHzxa0jyqaSbhQCX0c8BccLaEbTg586geiIhBZN
9WvLgupmDd455WNr2cXxf9+2CdbzY2Q0gW6815aARVwaj/pZrbqajNPOS72H5oo3
I44ECBmma+5pfSKmY5jwNP/kPw0k5x5XKKtVlyEFyXs353QBq1zwvJM8FIGJJ4ci
HPLFGYLLQ/i2xa3etNHMsoYTIWXCYLX0X69SPpaLJAGljGO/rzHpybneQe/xVXl1
IfBAMmaf2sknPYfd0jUu9LZHHlSiGYsfwOhrnmVr0UXhZ38q2pNVmevxmXVNgVNy
syKzsCzK/uHbET6UIy4C3vr/BP8Fc20rEsiMh4+yINt9/gD9CU+b41NcU8mnFImm
OOEpla/Rh8ft6pDi4VpuI6COScVkJ5wuMNq1u10muA57WgjpUlGVqSImecbeDY2p
lGzM3cqkTX5wulK+ajtEZ6Yi4qQYZpi854McgFhW5MHBH9sqzdW68Ht1tg2HXMc+
Ns5ncFeNeesbW5gCvQpejBsFJOeEEF5AON8K6suiH/EvvwIGCkh2X9qLx8Ce7gpu
LsS1m+DNjCr4EaooknoWa5CnVfV5lqS1PalIecNmUZVkfuonnu8e1/9zXfEjBSei
y1ZVrvGk3cEJXnHtSYCy6teKOKoTHkHgZ1qZeCgS7EVtW3xys4IqtyZVdHQdWHTv
62AS00lADs/MECHh25LsZjpJsvrvInzyYQJ9udLPIdEgGukfOR7xO4hSgDLFimSE
z6foNhIf5kNex8+zf3q39IaW47U8ZH3R4UKPC32pPzw74XFJf9Wwk+/LmAdH0iuk
bbsSou4vslq2wMW3L92+MsqENydrrINKxX4/rw4wjmhq/xpJec2Cm+peFvhNTuFP
Dmnm03Rc6mk4VVxHwalUcH74/bOyum9QiQeAl8vh107XwmDHJ4nIlMitI1fPvtwN
EvmMDWye916JnlyGtlR8AnEJlIdn5OIZDmYkzulYpC/v6OMNJfadBWV77LCLyDYF
6+LyHDSVZQ0KfsrcjH56AxY8VJ3zK0nLWH3AaF/xqf7qFUjZS39wLazCVoZ2aF3x
rb+FksvC1dTecbOgJWe+SNNG3ReuJj/UVrF5YrkQn8OjM/kYLGBwonaDCln6kNAd
7nS4g+8UZUscTfGHTtMqRt7NYTbT8A1uocCcdiuHMTB7WzHSsr9djqt3RZGhQxQJ
0CwfUqde6xrY0yhjiAGBuPAfU9oZ4X6c2515lCF8eAuoTNHy0GHaLHv0GlEY/plT
uD7b9p78cGjlpeAUiYFEqcE/IFXbNcDRo0yaG8xJlM3nC/m4c3Rn8qWz3uYWBO1w
0Hi9NpcQuX3Oh5OwVEX+4aYBkk1Tg0fleinoR26BkVqaLU05WYyLtSTL6IwnLYxN
Svyl063k3rGsHBMhANunuPGOTH4xJSptEp2mNpejc269tfEpzGNqzAFecIntfaxb
y3ULUdMfvnQAlysx3yNqjkeLSLJNRTvbh17jGROoODTLtXKahpjpJX2U9OZqJ+vp
PyTClca23tf/QwPy7TxXt/gbaTh1qke7Cxn1PM+33EgjgkWjjzm7wgxT2ntxRLGz
RocMQveVXh0y2vEc6uXA5wAXa2/PGkBl0jb7Wdb2E2hwPvj6hhRbehidPA8cvapa
N5zwUnePdqD+kWp5j3/FY778rY36AKvNf1isD9BlXjyCeMj8Ol4qERzYL2kiGDrD
+jjW8NXhkZuC5WZlEcMDAe0SWejsAew6giM2MFMEEYhvpzid1J56yhUrCgKTljlt
yQy2DSL+GIeuj4yFIlix8BmjwT4qBvpKIciFx1tQG54G0Nno/47RyUf5SkUt0EfL
36arPQ5vP/sx6ejuj71Of9CI4fNTtmJwuBfNBjebI7q5kqU/4BH1TkO7t9UP0iIM
Y27vbBQr8ZhqFBdLsg1w63/ArOQ45R640DVQDJXnEl5HevbwY9d4of4wMaNSJtmU
cq9qTwlHW8T71sQdVyz1boY+N15Z5l+G8TyoYedjhv5iozS+AcOhr/R+zgADi/fY
z4xVcLuKy2774ssYt/lxfRte3w+JssFPqG/MEm4ZTGSTASR9e/51l8XqB8icG7wO
hCHcP9Zo7yKFzSyKQ2Bqn6nuLyNgs0RvljU4sFPe8MeQX84mMkGVuPzGOOO9+CQn
ZXKQdncVSss1b2saGr6zT4wUe6y/9A5KMcVVEKmOANwFDo5c1/Eiu9VVLZy8gm3G
X9czlgPgP/BKGOJWcmXhqjFoqxj/jkisJraljRIPXc6QE3wFa4mXsHEZxrfG0nei
J2ieIuGyl4T0pXndsErfsDrbeN3vC5VX3544mVpTCS3k4qPILP0nAFN+4UPXyeDy
6DbHhXrUn3k7RFV/2yM6D2qQssWVChnYTauLAa8E6Ym5NJJOAoGnKkk0j47CXERV
Ue6dAC8vEe3gCp+OblRWqgIRNgP2hPWciGOfZdhf4RdBeZs/UB/U7Hlf0Ym2Cr2n
Y/14mr5bF2Vwv0OxLe0wrRi7QIMZ0Iba/ehfIFvtEOtEkqV+Etw4yVuC2qBk1aWj
ObHsfsVDg6B9NOnlfuwXTmxR8BYIDVO4QA8nL/2W/FNu6w2/mBI4MGuuEm5SW73j
dLqAub+Ljjrlzc9lCT90bhsfCsvCXBdCoDkNPr7vw5Giupk0/S72k7QEYdjdeCw0
JrRuhbjzcgJ+e1HgBFZ883ZJeQb4eAYc+jxFiDOL4O8V3UPhoIQgrPfOyUxoZ608
SpXZUAho9vvgkgs+0i+V6qyXXST4brSIqd1MyAHItfInw3kPdCayqZQPvzcRfbri
5+t6pHpgFYLXCGkp634izJ4ZyepMCuhryGAuF7aWoOhAVS+BcDf2p5FiwsFj7w68
O8RWzKej1l5QAwF/Ju+BU+tYSW7MJBSVSsJUjEPrfyArvCARhtgsOZw+0+aA/55F
D/46jJP9bCA6dZL56mIqgq6llFw5Q2MJSyXqRoIKw8z9AFbUy+YO6uw22EF5pPVS
5YddrFxaEAvQWqWhpRaPK8rdJSLx7RnZtHEZdTeOVr1jwIfpXXoZ+4n94PTzHvqP
zCUrwWWWlfPJEV4f1t8Yv5s7goG52aXKrIPZ3p4dmToKaB3M8gJNKVx9drIgp/tS
0a/OXSwJwY8OJ2yT975wI2SMa7hYyjUJ5vPEqELKS+eyij51Oeyo6k+kqSLSHIj9
9KRzJI327tWxX4IgMLitMVNFAHfk1Cm70yUlH5fZql5qVft8By9V8GpscMewedpS
w/hFPMvhA9lVQAkoPY5LHfVWHLjhchSE8nMeEdrnR+HpUjHrttHsoK5HSkCJ2Ud9
SkaYBRjASTv280yVDg87YEhFfvy5Wx+f4kevWBWRCVNrpkkVieY3vWliCES7Tpag
d+459MQYvjl9rt5LYH1dFpetcXgdc8jmtSxwq9lFEcMFsn/Qd9Zj2dqzhjsRP0aq
iCO00NU28/urBln47WwHllUseegNK7rNBixdXQz1T9H7xMdEOacqmPQThqKd6zfg
F7rNgITUGVjpsG3NwkCWLTS+pV+BpNoOXfv43buqB0p5nrJxJLgxoOzg7znDT21z
9rFh3cdo+cvkyffXSSVdvIXCkXkOMY3NkSutHZrjwGsMs5WwQAJHF9B2m+6hn7Ym
cQ8FH/Zoq9u1OnQclsC6sy2FWE8t5ROIhXu8+GtZfx0Yed++r7/0ztjjBdFtrKbE
vJ0Rj3ltd+OIiI7QyhPLOvHkL7O6UqcXgOSg+hoRyBBYNPAvYqOjMQF30PcUCJ1M
UIQBAUIwA6nB07GDgngDCd4Yj3s9ERfQRicRzRxUP0rXxZs18+1/3drYcPJ5WDK5
bfuY8mmWPAMEUwj+tPLLeuuQGe0QCx02Ib2+LPTJ6+tzzRtcrMETn4dTHjJtVT/m
9XLPu5ptmHRoXGRpbb4ibiLuLbRE1GDvSKosdDWnYIpfeYgiV7/luk1XipiAjNDJ
b1k2Ut3YhQ4+IrUDmpWqmyvrtLVJ8bxM/7HbK8pCvpOxwvuq8mV7XWeZGPnPh3I6
UAXmaU3NbgmGTUvDjt8hJxvd+qaWDA3M1m9tBztZ5Eko+Plubh8i+EO993IPM8lm
foQukBAr5RYdnp5wsExLkWcay1V9ier4Jb4OI15qqydmJ2G24kXzfpf1OMElCEVA
n7dGo8IMCe9XmyujfZW7qxOMvsi7fy3lU78Xn2chH8aS3JVZKC1Fg9bJ9OR03hlx
Gfyt7OBsPdBZGjEP+Ujq2R8pKt1X8UEvwyOfjYzLLaAfJvOhXJysEoGHeg7i6Ke7
4Ju7rVncw/j9LU6LY9/SNCadiUjbyUps/my+rTAbqRX5WggXnEgXfGKu57SqCC5A
s2jmmjJX/WwSK7/cqnyE8gR/Swc9xNpcUcdiI3yqWCMil0/6B87unVsSCo9wmfij
VWtVyPRwg4zPGZMUMMyUG9Uvq0ELX4fFDdS58JRgBoaOqJesql0RRUK0lS+hx916
r/J6mcRWnCzZ96jFWOWqh+I7Udt9qRww/gjiWrg0UKJhl984AGWtNPQrZFtvj8ov
JEpdk7GUoaXii1NoVXVaaUU8hIDJyuiCKztEFGwCzztMIjKBgkedUUcjZFBDyPiU
Y+sAn7lHUKO66jFyqefJAlpeoUk04kXvCq3WSOq94Y3KJbbnGFEQZK4B25e3/6Eg
bcSDWxdC+f29yzp/TgOVHvoII31kAjnHo4T2FY1+7CeHT+s6gZquGhFUCrFHjw3f
OuWZYnAyV2g6CFJXf9vN3vzgkDEWDO54HHTVqdcBe5b1AcDX+/8uVgE3vqX11bj7
kj3otuGkPZB3GBqM8A3GiMZHdE8QfvWhw93ydvFg7G8B3JDlrAlRqf4bc/WdzK3p
M5PpbtBZspj2fAXTuhcaqQt+HoM7JUA5fsr8ZdFlD6ma+u+I74BHbx5Xy+anl/wH
DUbpG/WSEZt1COVLAUABcOjlCJhTm4BrvN7qOXHnkbCZ/3LOajs+KJwrGFgVwY10
juxDFLqr46ApSeMhWIb7nClMg1dXym8tjbgL0X3n12G9lKY3SRHXAliJIsECAR1O
2px/FY+84GMFq0UkRXhgECJZzZxiakil0rMqFJ5cff1A06JgMCE3o/i+bJYesCX7
BE7I21zWTneK3bl4ZhImaNSRJpzDnqCN0jONxJUnC1XCnrS2V7+gHkOmQPeCvDH0
cxu/jSd5QOSdHNixUUGr1CjbSKzlOmcbOw9MaAa6g6Lt56ONDUOdvFG4jenNg7w9
qexcLz1VgDt0iPeUYpqMSUk7M2z8WqLB5iqbpObvmi0rsLH/xkLlvCSE5qTmAfmp
y5GZOBgC0HH7fkEB3AgM5ZsJsZ00CUOgQ4FkD5qXb7WO1X635q5+TrJOmN0ZSxs1
N/ZEvy/kjUr+GQMfhG+pMyd5Yci3ZfVeF4Bavoc9hg1qa8VaaM4MAi9s7bEojpHj
hv2PPLObL2sBFBKAG96YpjZDJa665LumZi2RLbYzag/JDVF0KY7H9cBOF9cmdW/5
7nAKaz8BxGDbyc3O0kvy24IRNP/8tQFHZUeE8yOVAafTvIgVFK0xQ8zVIB5sm8OF
neNpa18s2CTTYxCtU9ZDlz+n1C2iuarYczemnoJbeKhbz5visi5K5jXfqb8KJpME
ruDbFGOekSSJHxw51tRpbxYhlcyWpHHNEvnTMzsUwOjWVHurkqRlxzJ8QaCNyDSw
gLHG53p8DzPbgaLtaFx0fAvmKuTM+DAq8YScpWjBdItkO/CJ4E0Ycqtn7XejaAw7
TLRkMgI5igf+s/tCYNlsBzIGNJpJpEF2Yz3sIWKUxutQX8AN0rjBc66PjRV7zHCZ
mHpMF2JSx5hFzuwjYuzP1vksBZ8JDSfyfXz96LofcU970ZA1Kab0ZrziGnuRZ2pb
cyHXuKSQgumFGskLb2sqVkFE78IsQITE0Q/6pCL1ljInQihohAlg1Us0ZpXD5HlI
HOxwLSuHB58GaFREU9TT1f3OJfSgEB5+Iw1mYQS/IhggQpYZFSoHYfLGlpPQosRQ
gUNqsYOPgZT420rJGHAq7xjcAxdSqIx7+WASeM+CV/LbCQdswC/lhFpjiCJ9ANGT
4c2vFszz/fEHCGNcGxgszTOjjvqCt+yR8cU7gkKJ2YQy5Ryh7ErqkOY5YR3AgdDf
E++2KbQozssPGIVOwKn1sqSQeNavFE/wig9nBeKuI/jzUUokIexnr9VGwkRvn3im
PyK6fbHAyr6pt2VKpdr+HR0goTXVilkO85hoN6pe5sWQ+7Q6hvigCXuPx6Xbgqd/
azdCr8rh+mt9nXaPOjlKSMBtpkLCrLfKZ92YX7iOz5HXmf8LAxxDNQHNwedgp2zn
Qx+fm7XDV65vsOfkvyC1ZuAR4s/OROcd0vkKfNB65WaYxRyqPiZhVZX27/khZKcu
KSQxrTp8EOiA1FqlLhObaru7Nnp8TAl1H4IGX9RVYXKybyrqziJyuUbrjEMRewrk
EqqVaKM82Rcdhs8KPxpde3u2FnKD+pBu19MDtD4xxqHPsiswmKWkdXiBRNn8HT7S
SPo1u/LO3rIMMOaqoE5nCYgEUp9LlH8WTazG8GXbd0cordP6CUGQmdgPBgtU3fSs
64qR8gIP4bL7a73AyW+S9BYkeIIejtW3rLayXPqkINFW2K/gg56iMUx9mTcX8tt5
7tQks6Ki3kRpDu5S1RsgKCMPo65A9AqbzNxplIvvQ1bCCe60zybVwtzTmo8NdHe2
GT/zRc2/1h32TJc3X5MG5M12FQKQ94s6kWaDquTpJKLXsglKG6jpZd2LJVoNBE0m
NFgmudTNxEQN43TVhm+NhAZkwUyRkIYyzEJV0GCDcNT8Wbya9ZWhJxRbruZ+zsCL
rr2d9enN30ANCe14WuBcB2FVcdfrEpzjUh80+hzi5Wcx32TpsKHrNk1NCgH3n40k
qxI0V45Zo5YDdA/DI6ThZCFjCax+YCrF63naNvUzuI39+35MnIOSIYouvEJrP0B7
tI1oNPOXXAXX2B/cmEmOjp9OX9tk59B7TSY8iPmbjDgInUDXAFdkePRUHrbGpqrg
Uh4QM7jrsvYXq2Z0J4I2Av2KchZv8gC8JnX3sfxuod4012TPhQEMWjv/c4bTCayk
FI3pmHQICqub9LBQX7VcPcEQJUvsD0vlm4NUxYRJvVONOTZMc1nn7upuYHO6dlHM
cCR+UEFpV4UfO3S5+SCBO9Sraaei7oxBXzuylQlZAtdS8eGrZ5hRYxolLfJvdrYR
4S0VZdSpTo+AmWsfdoM2sTjhYYJ4QIf76otXvmdCgy77De2dATUIr3tEPjlPcGkF
xMo4IrYs5okrvXnA3/vupBpm8jY6Z8mNwed9/v4m1c7/XFFjf9nWlGL/SePXAADg
Dr/VTQwdgM8IbCJGj4jfh7JcUs5JEuHwIsEeWR2arSkQ6o8pe7/gffYYh3L5qtCe
UKirjTThtendrr8dnT9aKpKQA7juet6Tf97MxKds7dv8wdR5O298H3MSEisoTpOd
jhauXMUTAoOKgom5qv9/HEwj5ZIBtMPoWBGnVrnyYysaTR2S+SzNGqxp8RMHFKi+
u4aJv4sHG24/5LJNBcNwufxv4fvOMp+jqVxSrFJMddDPJIi6GUjklEjFtH0PC9Y7
es7malBDGMBvV8avl1A9KZyxM8djJzdqGMgedfI9vJSNi094Lg+nDyuTu2OFqn2d
6D7jSGp769GdsFCcRNv1r+QzA/8gSuL1RtLgpn5A21FNWiT3poDhavBxdFo0lPQB
l6uEF41LR3i1dXpJoCKmQvd/ftwXxx1aXPNJjINYC7/VafjKMuXtT7zTZy6tIPQo
SDanMrzCmkrPwHjdUSS03Bq/C4auxt3N1Fc9pH5VRxKKg3GUiaKyE+qZ8L4TVdb3
mRyax+YpKCO4FU4E2VAFzEyhDBfkfovibVrVCEk16RjP4nQihdOq0qDbPZvBAWqM
/qZKZH6wxJghrjZGaqiXZ/RKyYVHE2nASk1NQ3pSaAAclyHELolyzgR+v1ogHMKH
Kwk6CCfbCcjfgGEf/RUynHuGC0hXfKm3HmPBIYLySeIpTB4gzxZFgw0bfwrOS/j/
RMczusD9NdNaWEv2eq16mPNed9PmK8nVjuR5TZLocsVDowLJwlJQTVagADd3Kvho
bDMrLjaIYQ/bYteqJtfjWNPO4gaEiX/X/COzdtm7UXY7aqsW9t3nYhDal/HhsbCo
bGLSWu471HVcveea/iUfShUA8/5Plm2398c9xoHRtQsQKqcNTORhhXKFXlKlJ5f9
0icYkTyFXGlRYTthYcybqR+j47Rmu3NHUtcYZRx57NnI5ErlLfs6sVldZ/K5RuHm
RVp84XRA1Hncn67zVVXrx3SbM5C54tB/naKtXvvIOwygiVolkQAK4wYCD7HVDRRA
EUbGt5g/K82mkZbdG2K3yEBLidEkzNr69ENaymoo9ohJ/9nSdoLMawXG3DLdDp7X
kRirGvbf56lVZosruxmIcc+rNAZ2sY5mD19RrhcwWQoC2u655JZyM5cgCTOrj89r
t8IZq89S7c+SkM72HytRTEikvhZNkp8LoQvBtu1EzGXPwKirY18vGAEG2KQWWpy3
6lQJEpD5oMOPmtpY7rQ8IDcmqEQ0ejxCTEvrzlSwVAse9RgKjMYTGnXEBJI01877
Uzfa0cWBpxuLrOZSDAlcPmq1dVcEeBc3HHreFbWJwwOjRHpy3ZnZLY8ggV9vBs54
2+KCon3ulJl4cVnXftKD5tZscgqSDDE3elxceNdlZTZSnqHqOCMVgFrxMdE+Os34
GNYV6CLz1WmGlbcT6GMfNhGwpurtykZoRowrVC2HAsCLZUyGgIJTEP5RqtDwoxny
j2adcV9tUAIRk6kSPmdlC02djRuquUHLhdmN/35TNHyQvN38U5ouMhv4AGy9q0TF
tr0waFKYfx1qW6UbSDvFbI6J1K3ROUPuXwW966ru6KYoxAnKB2sjzy5QqPJU4tbo
JTgsOXLZRUmY7nvE3YeLuzhq3a44K3xPRexuJlocpm0JDXmktFQEc2BAl9pjgsWt
76vgNOH2KMf7NipSnuA/T4B4z43G3rZKejwFEiedBP1VIpYGmQdNJeLZd7OmZFVe
XScb/a7HCkN9i4Fm5eS1SZikqIND6DnW68h1MHZql2NMQyRhGyre7w8IFrAo0ceW
NpLW0dkln9Y/PMSfFqYHQjAPtgp6WjaEcRhiYK2Hj8pBIvmTLUUfNqJCt0eb2a1O
aj/B8ykvZtfp8563y6bINPhm+CEM6AP/Q2us/jCvqhP0LXE2SMXdk5cgJ2fMJ60o
zS1/csDR1QRRxrXcTboTPamQnztg1MTSSQM7xKajwCXO+cbFYwZFw0pvzeK8nZ9f
5+ykm6f8UdjqrTXY6q7fVNPBdkVApMYok48LwOhWPVlmTg9OL2GfU5rZWvGfYcl9
3W8KyNxV/2RB5ZSuBSOgc3I+aftlB7PTPzDXWf5yRD28Sezc2OlwlDHpNdO8BKhz
ywYLW4aTCBxk6ioSJMfbXmQGBAXnA7ArPBAgB5nEU8m8CCr0WOGS7dj+tGSRB5S+
0sbAMy8DixOpVlxQtgx0fw6xqdkK9Wdl/+/T/JFN0zPDM16L3FIpGp4y+2+WxW0V
C9BeBrAmcw//2X8tiLF+xFO3hqkhpw4jFQBEt4kPrrubdnxgX0PYPEzH5Me/Lknz
7JSQEx/SOwheyEDjTiOG6or2v7rQZiegee2QEmSWYotwvIhuQ8TjkOi9P2u9brYd
MCPTmEygth2CklIs4GBd4Jqt182d+dU7LXgmq+fHD9/1GMxBSTfLo0UlkUk93X9r
K+m6siRK63/BrvaIsUX250Z1sYeaLwRCDfNzBLKTgbImQNMUpjo/uZFXyZ8BKfqK
h5f7+dK9bFiL+r/nS2WnxLoGZKoK3UPEgsbPQDIepA4j0j6QwvZeUHL+MljaSLSz
CfbR0EPib7ojex87Q/rONK2tZTInBM+b7qBPV6i9vE2UJL1VnR3cvoxEDgS49FDY
0PZyfb86KGRVY12gC6oycefQdaCp1IUGPRos0EHgDCecDDPt29x5+o9Ty7evh29K
K/nsbi820VUOSYQjN6Oa9HU9yQjrWElhJZTzXB3XwYKpIb//lsygbh7y7TA2fRA1
WSkBt74Exjm0RD7DaHPXRRU+PY+h2op4DRtlSHVHWst8SJXjWiUA3JvhUWMSYLxt
b1DCrUguNs1GJCUA+i14EU+te/2KJd1kXtuxyu6afuOHgBo5cgRUyhjFzS4HtfEC
WntxgtbzHXVgfcOAe4GeH63VyecKvT4vw8H1I11hAHfCos+E9W0m+rCnEbgQA+2/
NQmjuDFTqfUcit1vuSjwVbz7U+y6hVjrN7WS/hiZ0Q8K1eVuxz0hkCMjUtHVwYhy
RGIN8zt0QhBIboQeg7SHi4vvUqvVid373lv80G3fNIJ5wtzf81z5uRFMU5sIh0fR
cW22UAtf8nd1x/2e8CiVewhgSAa1PjdDAU3eW+aL1xpY/mkYxJd/43TtFXmiIyjL
IxH2W7obJoM0RKCg7nP+kTAXZc5hMidREtuvgv/xo+vN+F1dHF5AAeaFp/FdxtiS
jdB03rZyYoGaWuHznBaTUAGXTIFcCz02MKtytUgn6t6KhGBoeDojzD65Sezn7Jxf
gVL2jN7TtHrJJ17WkCABFZl4uM5ZMuz1sx/lPMu0DcqPxjxjv7SwFlHw8zoBcGxd
NLw6E/uwM9l/Y4G+fJgU8tL8CkyTMO4A4Km270ueYoQz4mvMsnOH8zky/ipW6kv5
YAT9kzaX9lCcCV0WptZU1XSISZ3p8IG+69osyaK6JcSWuaCG82D3Vk7JVEIqlmNs
bUxOGuV2Q+YkJfwxDkVtPEtTGZdleAaB0qq6DqgyzprlcsBK80H6BvJBqKXJRXOS
O/5o8zzAXCOFGNHa2G36JYjV3k9nCKQNtbnCq5rOYioGPY59xIDdNuRd74xVk0Ea
6+Veg6XoLZjdam7LBnmWsQU4H03NMrEC/ZCIAxcM3DvBh/xrN/g1jAIm06wi9fyf
KZleWkayWfBgIUAy7ZK1fWlGj769aovQl0E4ey2P/UVw7ZY29iFcWhs1mfiwEYgK
oCHpWr/dqKZsq2HimheuO5nYYG3GaozbQaAp/efoRMTxICk3dv7edS1Ekz3QX2iM
MJFxqxGIb39WDlN0vl2RFkTPhe4speXIiXhNqWvB+XY0aksKSfF2SgiCzVvV0BEu
3hBpDs6KzdWhYcEdVHuiHwujEwEBRNawqHah+E1NTbyp8rO97W62oYpRxNHJKKvZ
uE+bWTSTzMGBXDBUmO6GEZFtwL4hRrcQiQH0IBHf1FjjvyW0Ip90BfwJ/8v8qMpy
d/L7MA928myeJdKRn4i8PHHkXlNlekHy+2Qv6ebsN7+rA8fqHFqVlmNOrVDz2JJ5
GG6x8Cy90aWawa4kC2o/AVB9OBAqltMrglNIx63GOXukeCa6AwKu4WdkNOJdykTd
EITXT9zRZbzBBsmrLmgSYDOAooSSn6NGjcTk7pfdEa8JDm32ZTbA7V5RhJZkW6/S
IcqTBndQzbp5bLbXw+3ss6HH1i50cKCfJI1W63ALOV2NItgbtBzQf50dqSsqgyCD
nzxpIs0/orkD41RM67hk/LmILGFcMjN3lYhL80eYyi2ZYxMPqi6UsP0Qo0sWSExn
r8INcB56AcmOXHBnC2S82yRiZv9pm+09gJ2ymoVn+gPe2fKEZ+8tiWePsKBzAN/3
tzsBO9NEUGyDqSr0Afh3X+wabmNPazqTtzodHYj1+FRDgkxnLL68zXSxiS168INh
snV7zZ+ymBDn02IIqGr2v77w8H5gw9OBPF208EQvOn3lbou+EDWZoQ6WdLlqQJEw
67MYqI6curRc0iUwlsBFl4cAOgiMMLSacVKzg8bOiIVRqqRoFIMIKvS9LxdVr3ma
+IZ8gc4ZVezLc86zwOPw+ZE0avzXbN2dX7T5ZPfMr6kVN6RO2rgp2zxdKa3g3sig
IFuLPWp1G5iPtTrIxLDi/gDSQ3A64n121/rSiIfEwEiZwqX5On9VssyyM+Kkmpvw
/zl5RGIQ42e4vk0o0tIMYLw2RZtUcXe1X0xY5ra75G9Sa/JzXashl1OA/LNXaCMj
eyCncfivo3iaM9FrR4cyw9a0hwlRGUm7oRIj9pYUMbo9bV9VHL+D77KLTnk8T5kO
6b/UntgF/o4xzxX3FzhKMOjPSu/VNAbWpPGRAz4VLoHWzFTQcuWaNr3L6OG24FIj
wTYTym64jYC9ZHg5B3QAua4qWfB5tD+Z7ebCQL6JXeRMuuGzh1L9Wj2azp03IFpz
OAiWzNTajYmiVgUlqkrORF/Z1fcy+XcO2mpMqB6Cdp+LuAidx8gtoThEXjGi3oz9
Q4qvT8zEGx+DMmfKiMh7PEBuKLYMGaho+Ks2Csvw4HAJfmLHqPoKa2qGeCHqw1dv
b+Zhr1jkb8DmfLjH5WZkUfgduR2r6wRR3+CQdw+U6VHZeZ6WvDKROshtRX766gM6
RMrkf+HAAET9TeNCepUQshhh0GlJOMTRaybFgFKauT6UZfdEmdmTeIJ/Kw5vpmb/
mLJ7x6C4Gyv/yo3aHLTk9ifa+WUWUqiUDwg+CE92i451lmDXXeHEnH1Vvt0TqVdJ
PRugwfHAlLtZZJ3TuU19JeFwXoQawJknnlsNOdr/N+XrS3c1lg608/jxHUMjlRp/
z+qdXN9m3nq+oSgyHykGhpW6w6YzzQiH+kdY8Hpe360TNjpGZMun8vCHfDZXI42Z
jTp9VmyKWzfgaSz8O1MTjBCStGnPOb/SdpLhzpqrmftJvLNgEQZ4ePJg2lx7Dzmg
hLYdmRWH2BvKgrDAjTVfjxxFFKiLZ4DrfRDdqxXP2oFplEl6mfeMzoLgFBvtA2MA
wUgkGf/C6HNCTy+iSx7bwC7bqiRkwS7SamE1oxpcAWhsa/PpYClXuyLQi9/ULXI8
4nDK4rOl5BlrERHNc6uCSRSwdoDRsjrlLCJ1Q++f0VS+tjtHdD8/G3x1TCbZ82MB
AbYVybHrkDMMgQkoxCeMFfaqxIgdpzBap/EKJvdWoW6t5Tlqqct/m6BhMF1vGud6
URkkOV2xeQip/FlVUHX/a/gxTDHMbhYwBCffd/B+qRopIxzlGEVWhQtwGHp/xVST
5moReZV77oXbv3RwsxwqvwE7QqDcKt0Zs/gY51WEZETa+EoZGgvGFXfkmXLG7bK+
FMgGMeC59Z2q4sCWqIUb5i61kpks/A8ZPCN7SZILbYXV1SuIN92feBbH22dFa/jd
cWtsapWlqCI2rrCASFR2QpAc/ujmPMQE+v/PLmYIEL65OaS0AcDHXanDSyVzIHe1
iaaH2g8p4eEYtJiaE8F8hadPh3jO5mlEvqs2J2MjKwY5Rs6eDkhrL3Ib4760cAK6
+XbQ/l9CBx+D8Xe/XR/pCfv8GCBR8pa/hjuxZqfpl+/nzExIMSZdk3yHKfrc2Fra
myWbUP4gbl7GTIMypIwSdMh/bwYVXSbBpxLFbZOvi92+OycrU5W8lJ2euu7psCos
aSS0/BePihkHqx9H57ZS0Rol1obAjDhEoNPB/CugJIPhZsMz50Xky9AzPM+4zYSN
R0ABsNBE9KwoMCrfKpjc+WNkBmjie9k97cBgcaor8YysIqdsIP8FYZmiWAXLsivz
K+IgTvWAKwxVA9290O16FGd52P0UFTGm+ilxxnJ7wfiIAWkJGMCsypiCl1brkH5g
iOXxeUIMuYs7W9z5LzXQynMICvbxwEz2mhkhZB/5z3P9mwLe8zCMZak2Mf6YJ/Bx
Q5lCb2L7M6GzjNwMkR7OE8jltWwCcd30y7ooabWKuvqoxWyJQpHt6Cx7au3JiFM4
+DWjcDEN2lrzK3E7Tz1sQrtb5W+gc+DQfdvnegmVvPAzKw97i42XE7d4MbOpyTAj
b4WYKL31XtaBDJllfWOwVSJNBLuFb3PFoiqzSlj13FAjyT3FMSN+czQEOYgoRSFc
WfVqYxxd4/8esIjMmE0rzIL7IS5537Yayj8G1xyn2Kce7vig4U1n9eyOlgzkTwfl
ekRCOzj5F8NLBRx0cUc9LwcWGZmTPicft/K29T310GRDI6i/QR11lyEaInB0a5RJ
AjqPP7PssDwtUK2eopy5Xgpt4ICTzzICoo7nsGV8W8Z41UJ6EhnD5BGSNo8Sj838
FXY9GfRUHZvbOlD54KdxLl40Yu9nusZHWf04x66Makn9Sm1w0aaxxaRXbL822CnJ
mmt1z9W8p8thXmw2TVrbFT2fe6xKnOhmas3UdAGbDehMZ2Y2o9qOL6UHA9JoVkyy
ikjVDvYk/21W0QOuv+FiZKM0fYFivML2kfGO0qze9n5OjqgWfn9us8k6rQWh274y
KW4GPUbddsGhbQEszAwoMOdtkJN13N8vDXKp8+POJE9UfOJwnGe0XBRTMC07DbZ5
vJ+XOCaSry3seN2PM46BFVBdCa1kYDdBFe9BAHe7uLorm/YBYZ5w0J7Z2bWc2T+2
t1XJ0vVN+rLtoo++84IbKb5cuggLNA42sn9iUP48zBRuG3HEb4VNXeqoVFUL9Bxa
IpGNnojCtNfU9EexdsXEs42tsQvqMtRfl4D4cSxKiz7uL1R0gXqA+sN//EvMlHSY
km5foeTKjLubIHA0gBitRiNO+nsWG2wRa5AtuKoz1IePot+fiM1hahXHyKKFWu93
L8Hzg4Zu+vh22SzNyglYfevgPUeShpFB65uw+4WuRsTSrhFkOis5ZFfhGaF+8KBf
5LY75+nv4YdPsveIRCA/4M/K63ImnqSZMN22mSQRY6ywHST6E2TFrQZ/NAUDizdu
8aPBozH/UWLponOZ6QvWPQMvTxad6LvRZzMyOKiPy6CNRpWcKpkzvgnzVqsXm5uu
IOCW2A/iytVUNtYJBfqixo5zfTqU0QsX162GmwcISN2Cqbz/9p+QoDeOmERgvqtz
XE9ciCiKFwmcvZVnuzljQb6EUsUbGQ9GtBUm+mKM8G4S0zHQ16TXYcVC+8q/fugi
qUBBiKee9Bt83x/i2c1Qicx+ybiDqp/IUFEFgjC11Z/Xyhv5mcJP7X5Hi+NxTRlq
6RY9HJBjnV8mk02/Kvx8i/gfIPw12yGGa+QdUw5I0VciZMaKeEZkbtxq9RVt/SRf
oaU35VoQDASAvAZOPd9HOgvUJbTZoaREkABDYcy5Kd82oidAWQT2um6ABpaWrIFV
0OkuCcLr43pIUKl7Q1SxTXE+F3F8KZxDsnAOr34w/vOYHYvpg+pD/DbCcDHSOnrU
Ub7CDfH7v0R6PmeilWsio+niUr5LVF5W+0y78tsQteomBqMmlqQ0bwIdoyd9XME+
44xjYXenfr7yZ4AJ79Dsp6rOgPuw9dM7nF/BPRt7nNgYSAX+jo1MKhFt9BimMYDm
EjdVszc9Srja5pAgz7RqzKn+/Gj70ar2g4pAQd52TFapR41rP8P9jcPoy6FiqfTg
H8+wK0uC2+7bwp+WRR6Mp3c7S+RDgXCYWU7mRBY+wpiNs/SEUeaDb6xmF6F7QfvA
nFF/gkZ0uTGpXOOaJx5xqWgbfwVVuhzzNiho6TkHC4THmzns+hNlo9iJL3va0ya8
ixElWh4WAC76bWPiu5HeItti2lB0inKuDXhF8K88K7ZTBxuepS1eb+11TLMBkNld
jBEotUYXqXQZr4R2bXWlOwZKkXufaMbfO89UmfTK4CD/JeNpJIDrK5DKl7Vg9IX/
78RCkxqYitrH7l5FiOxlsFpbY6gMk/iDndkBEiLj7d73Xxm/4Vo4jPs40wzEDy6A
mEwclG6q4wPofU/LlFUwjPedzXCHM8Cj2NyeqZJe3MYA5nnaTUVaHYYGTD1cURx9
DXWnStFEnJBGZpJKQ744N1wfJdwLLRyjQQ6BYoI8VhMFPf8zR/KhZ2ay0VlzYV92
8DybOBLdt+JWUMVIulNbuMI5YackxRDykOv+yUAXM5EV764jykS8qdtBqBHBVqEc
o/rDnawSxDcasVvA2w5Cd+s/VGq9MgGi5mtYwthL/lwtFoxfoTepoH4Z5rhnoe6+
kJqW2v+iyVgaxZLLxqehP07EtMjvWDovMQv0zkKtOYX+7Kr3vPMY5lBzDDkMGmpH
7dUWds+sYRUaPob3cLS3ia0x/ZR2k0AWbRkB3mdW5iJE6ZJy2F5N5OnLUIcATZec
yPVNV/n4PX5ARer7MmGPqSs9xFAu/DzeZjgAaCggMbAJb9Ld7INXYsGt1ld7TcVW
9WlSf5Y2DKbHJIgXCp6zGsd9J8MC94/ygV3nYmzjIuhpIXVELfzoDLy3lramfNAQ
XhNWdCfoqTnXS1p7i6Z0DbwwrKkLVeLRgiQBBX1qX3vYtE/8IWXXFFU2CgpCZvaY
a3fEW8aRSqy0kAUa2xCyK4Yjs8XmVG+OfLs3DawRg4vzNAMBylOz7YkZviCYDTpO
iqmaW9an3C+CV4+2Z/3WaQK1n9KTnxaCT8/e5Zbc2uKqlfz8UHn4pOT6HmaPkvmz
ltSGSK5X4rxQTJlFjk2OKTATvboZghcu/XfNNZsgu96WQVl5s+ORaMlSBggwxdoW
vPnW3f5qJOXOXbQRqMl+x62kPYm93ZDaWVhPj/OKZ1XKMo4yHAuQrXIgDQgrM/U8
D34bAtvmxCQHkmv7a338aTGDyDNMrBcV0I3v+kwIikVnt0tqZPRfUWhFqEAoTrBK
IAc0gju2RMR56e8HnAQB1B7uEMEkd3UJ1r8LoghbuSBeIJIzq0ZUNYo58sSec4x6
uLz0h8KFM1P72WLPq+OSbvrNjcdmiN+Z/PCV2YfQkl+2aM1jofmjRtrHZw+xr7Oo
zW/UjT5eeSIiBnTajgqivapTKbqpU6e/2TeuDP92M3cTns/XeHYkFBuOJW03buFw
8zlCKwHBsW6SmEqQvfnaNjzF8KlUc2u046vR7v1+nA/1PGLPbYsr8xkndOkbLdwC
hMhCUqPucmshKz6Ki5CjJ/A9iwSHg0CQJK064NnTLaobo7kpoAZ1RHJsYW6H+xRR
X23wn7Wbr1lOhS3jOSfxzKa/qKCYloS7L9bk3RNc/sxB3j3LKXZoDZn4wQwT1DjS
j3MvExk0pngmKrB5R1W+CdLj1qTG2hA+PohLOGMr1ciXhqMS0FQEh9c9lO0/y+sj
b9YOa5Ov7b/3g3ENFIT9S574iAtdpjxLv5nO90RwCxGiVswr+cAMLviofpCX0JLy
XvgeWDRn0rzVyYu3zKXKZX404lj+QDnOvPp729bHEC5+3rIAst7Jzoz57HYGQRa5
4g89UJE7r3WN2FTxybyHf0bxtBlUK5YfCY7EmuV+ftqat5zJqPReNq13MPRb8fHw
ETJADkXqgGCB17Alqt4cnEy3hINKIx2g4PRAAD3KWgvB49aTEGeVnkXnGkYm9Hfg
i06dWXK9VLPSVM4PB5+jSvYg1U6D9FyzXgkXt/Hns2dluFLENf3XPFTA941mcbbd
NzyyLyi84NWDSvtSnxnBFXiKJv7r9PLh6akGIWtzV9zLe5KMxTLp438eI/XUI03V
2nQSFVmrpbDYh9JiiAzcRJ4z2zrusbMfMjkN8bnJhbWMlguETTiqarkQluYYndPo
2tmt3WdNPsM80K+nN27BMjp8chw5CFUdmXdBfBqmPyj1wNK3CRR6ZgdqYE4PPqmy
tl/IA01cGY+gNTpwM2JV7096NcFn8VykLBwiI9lQaGMc49/yBPE1vIX3qxtVf/fH
DNRMwEzyzVhQpN0w0o+QP6HlQBztoAFnErnt31JtZ76pwyK/Jp90DUq2ftYdj2lz
yxXxlveR84WzeriYe8UZJKdy9lavz3AOWcpoW33F4fT/ADekQBQmrqRb/z1u4fXk
5jMYNG11fc7ZsuRamd8nGafMpW7n9Iq0QfhKD6RwEzMRRO0UjKSGmkdGDsqLs1f3
ZL0TZKFEYljqpI+AmXayYFC5EeSgcJC4nmqHxjCg+joI7QZMgktnk3zPBIKp5ygR
SjUU7eqmmHNPDhIplgM2jxZBNNHJGv/55LDUC5hd3YmTzeqSFJ63kV2kvEXiWAXu
c9wrhZNg6SXJarJHTzAIVrVjl9hgjCGUuY75nR1kj4YlMBk+6KG9SvLzpacykm3X
eSSQmPjh7qK3EmsaRX4w8HMCvc49WlaTEkfQiVdpNZtFcexE9HwJUdtET3tH5wQJ
ptYzBpvbOhLY9g9K6p2s7Rc7mPcIdypoXW3t+a93CgAi18rTJg3yBiOAM7i2Sxpl
7QitgiNRf2ZakDM6mehGWfeceM/DNl5vaUmUMgiFOKM6/B3Fu+FFKnx9swAb6vnq
fAo1Sv3OUOUmOPro3+dyIVzLcSqVOTlTPUZPwBpUR/F09DHt5OpcLc/Jf+DG4UZJ
Nxc/T8LxbmoVUDAFF7P8Aeu7itoSaCbdO4BhB1sinAAW/qhDnL63QyQgOuTw8S5U
iX54SlDi2CFxNPNoNqnfgqpdD9rAPeotS0Zwhlf1r7gUKViBikr0UgY1tGN3DYBK
06rpyfXXVOn7GGv0VSFS7LesmTP7GKOSI3Vd+gmvjQh6sEO60re/UJbNLH5P073L
h6cd++cmsbDSWu63WrW7tIwvljPVZJvV82dKgE/4QRi0i771t3a71MbQzyO/Dytx
7Kbe6rO+v/F/0sJRqFMtVjB+SWmQ1iE8+sjUGnDBvXV1EcnjN8ScUh6JNLffxoM9
U7gsqNW6f3JYWZNrcwvWUXygOkdjsrtmMpWE5jd81NXJcdqQsGjGj5vkMyyhDsQf
5Dwh9GNI4d9v+KAb6E3w3elYjsZ/irk3dR3bbB5tNqSM/Yu6jhMfW6pmCVsavhm0
GMlWlfJqgLDyj5wdNTLPMf4iqiDbkTYs1xs4/WLuNIFJCvvmdC89JrYdtOq3F6EL
wgFsn1ivj6Ce1absbzCptEzhHeyWyJh5YFn5RaQN80d8s2/d9I8FI6I4bqj+4Md6
jPzOlan3zdX5vATlU7M3iRxqrtMssMmj88v6nDsGUERIp3oWhJ/Ew8CJxTHa3Zry
RbuIDAYnV9nTjfkoVj5gCcelx7XvmfsgcK4KkXLHAYU2QpRedsjazcA3b8PM8ksO
LpNEkKyB4NzEk3LORvsaIdrxj8UB7VQeQ1IhtoJNJdPP1NrSJTBtGjWOmxWWg/jY
kXfz6z6+aZwtc21lryiArSU++DPvDeD08xKXhZfs/VATNaBXCaapUnv2vkPW70A6
ijGO5D3U1i/lTH6n7O2Ruax5+2R1L9FLyio8j4pPopx27oEP/h275s59qbZrgERB
ESXxa2lYZsyUKpX3MmcMBiHkZRMNxA/0ZJuqF6xo0LuBqxO7Om9YOt7CvGLcc02R
C6uXlFX9bOp0tAC7EyW1GGiuJlODz3NJM+cjKjbXhgIdPZfGYlAE0ih6F8Cdk7ks
hoFOvpT3zLxk/kkzjxzvIGfHhEvV/ILobEHbPTQVTWWP3Qg+d5UBBn1UyCdxezl3
BAxCdRYOlliizzWYapXsNNs+RhhGL30lTU0Hn6lZI0CrRlhKprWtOldq7vX3Mr0k
sbUkMQl/7B1aCLJ6GhFjZUm3ReXAqmn2ypGtdJfBpjtoLzUde7nViexD05/xA6gr
SeTQIDFYfhlvNT1X8nh1a8INN91OL4m3LD/VNcyBgy/cHzz8qf5Jhbbr+LKP14JH
di0IFlmXcEEMqEfqqNqx/ZQeYW7/S2u/u2ztA89hzeJsb4Lgq8HgaEom5XrqRTX/
1fY33u49Vw2TZ/5EON/q/O9zq5jnZ3Lm/aMfFYxm8b+dyFOKv6b3DvMwFjd/nGYt
v6Za7madeCXaERiWdfdFAjqGWyqr+TxESQ3ASX5V4/bKS+SVHNiFEg1klUJ2ROS1
NUpd1Tr5121D7pzFelhe9WdWFDLPQ7Jq1cZFYPtyoFhnmLs8+u2q6AWyBPOu5m8j
Zf3TeJ511MDTD4oDfvj7HgYpD099ObGqoKlDa4b2znRq4VuOrbNkB3/AE6L+NjZ1
cpzCbwICiMiIOWdeLPn0G5kgr66MAhm8Xy0X8+W4LM+r5O+GjkgKj90orIOTl1Ip
Lp2BGqvdi168Is7/lH/19bn0nQRH0H/IxdQNnNjrJBx6Zg8OdB3LFAOoekailIol
6jEjiyzXuHE2xjtaihBVQ4hbKMCxYqpkG8EjG0ctj6LVMhyuQayiGmRgNrJ+h2lW
WdYqlzqA+m+i3eyuU9a17oNNIKaqRhLZJ98hZPQsyqqm7jRKISHVr9E8OihleExI
BB//J9l7xyNdQlmihrm3Z2sWcj4v/oqmcumgs9t3oN8hhqgBh5IMAh1y+VPaZIs1
ivIdMDALEHiAKlOD0xOsidhZIGfuxv8moXGNmsmLF4AF/UP+ZGCNgV4nN15sOK2g
wLwgv4hnq/co1NoU7bpzfIV2KD2udK3qyLbN91dWLJVVA3pEfONOjpGlaIXFqHLE
exjxWRbLDmMufQWEXacci8YYNpBpk/oosyj6PJI3aLq5GBSa+PvxQR4frdNOrrxA
ouMWqrXNekbou0No5agHajpzV/362GyFoT4I/TMahZC9M8kf1TdlG31o1LURu9Qq
nvf5H1dfvmvQPeyqtWFI95XA1bYCUqzrQJzxghRbDxhQIwWhyHNWpdCsFXZ9h/O7
Gwu8p0Uq7XTgmgNeAP108jWN4lYa7M0lcVfXzHUTnSa5jlCHmnRAlRQLKdUW/ogI
OLzw1apmswAcs4BlJrmH7LwQ8JdVecj+UNSeqEoUepWRBTJdYhXSlq36UDwXVDB/
b85IgcKj1ET351t/KUTaoRyxD4bVxiMe4RltU4AO2OhLz41vdy/GuoN4cDh/Mzh0
xw81gN4/6TILwmAbTjYYI+eQRZlivwkeMdNrM/bjxPvBjtXihxQsJX+slk1tfrka
N04ESL/1UbpGK85d+f1XxNpnMcfUo9UwPPb6MO8cSpxfX21sI6KRH3av5O64DIIl
WJl7hRip/65Xlp8lV/+v1rGW18wTtxfwySJXxxvYRoIQsj4xvBTBApm3tqvE0dns
Yb/dzILJeNK/usVUGV7HMe9HPHt8dzsyKxooRD0wFLuLYT9E3efRGY1TgpNqU6bj
4Nr4So8BTGhzPRAqjFgmhTQHXj5t19mikzQ/SJTdYKy7WjcrBqEl5/1rL4MZ8ty8
O2mldkkgqk9ZnroEZwShYL9pnnFfYdK1qVPqzNhssJ9buVSCpwka+j+x9Eupx64i
k26PEUVXeVVh55nGx+zHMq0Qdab9v5SgdrhED57RgWSxuus08P6u+M4sPmIRXFSu
LWHwsUr2x0BH8RZyJsH/Q0I079dQw2KSP7vegRsAjvS5tGQf22hydh1hapWtdIJS
Dftbf6iwyTaU5buSz7qf6PoB+ws0E/l8QNshb8yV1GToLXMZrXgZBaNr1xxPcpiP
FSv3qzH8wzR9XgwGcNhPimqSez/6HG4wS6gVVWpCa/UGU/9QSq8+1d9VxazshDHQ
T8czlbb0Y50WjZSB5q6WjzG6lBcefIrG0sEHrixgk6PDm03bTByA+NSVnlMKzli5
yW+Enp8gQVI+ErLcgkUPTkaitHr4XjX4DSnc3ODGAtl2CrxzuJVp9ptPzjrebNKr
z9hGu0K/uP9dc5LpUngwga/JwNuXaHUXf+UsHcdYsAT0p+ydZOKTvW95N5M2gvGe
dtb0NnV+axtFu2/RJ/7HERbJcTxjQlxZPUzrGtpGXGcmjCPrxlZKmek62cUCwqEW
cgAa0Ld0MJnXwTaO6jRlkGyNlvL9YUjmmACkbonNjLsi/dX3I9p4nP7g8uVp+QJG
r5waCYSRSgF81xITnKz5KA+zxbVSPB2dE4OmJB0vtcaGmv/ZkOXGTl6d8qUQYZWh
muloXIzfoXTGywi3yhXW1DiVwiu2tYIkXTlV7t8gfsTkibe0VGtffWB0mv0yTqJa
Jn0hjl9lMaNiMHxPPOW6ueA0ntRT0NYOhxGDvWX8IFDmgaj1Rzf6QJj3wuOF5lct
UErEPac6DzJBc8fiMEe3AgIP003P1yEvX2zbeZeoKf7K/hhSwR8vfJcda8HwWnku
XFtG9q7jTOAAaRvOnJ6GOcS/p6JCejVF2zCmVeI7hl59RxqggPjZVEip7ckyaSpn
yJ8jIqrzbnoAJjq/wUFOm7VfKdjPsXhUyQDZS/iTCgVImth+CxLMn3XxrLWUSM93
OFA9j8a3nDhwYbXWzLk/hNHtXWaMDNI0iFPGPTdjuDEH+OmIkVFEoRhBBzIqPSwP
Vkoh03I5tSFJch9I/iSqab2g3fI4lndAByE4QoG3oMKljsLY7HJZ84RPpVW76Gne
qhTSre+kgsGvIu9/wpVlFhzvNsFUYLkMk9LNQETI69OPOV/iLLVUF1BWnNHQeqMu
rJTz6bV6ronI3b4zUF7AJ7B8HM4pwjk22Wn1vbmIn41gbjSzMM0dUS+Fblj7Qs/r
JETqPMD5dp2vPeRYxfWtq36iMFULiVVWHlSbDbTVjRAdjplaEOHepB0nC85wD/9c
QosUFzTQJx16ukwXcXAcUTeObNJvODdnMYv4O1K3qe/8wsOSGLTsE3lc2l3ZBGF9
qL51LgWwfAFa4l50OBOz5Q1HevS7LrWRmVTuYVK3clcua6jguf3bMHr9YM9LBm1Z
AvozTWzIze3RMlu+/IUFNqWhm0cyuJ0JXekCAgDH7zZxzsxLsscomeH0NzkZscbb
4gPo21wlTGsjYOSJqd5LpUeKJGcB+3GVCWPw3df3WeAwC+zwykbBwAxW3HIeQSfe
sOnhD3Hzjzx/kTLmY52IKP/d5prJ32j4ugpNjrFGToe/zK9b9eR/n1aUx5voK/XQ
BY7kuNrDCh+CCDv+u7TGC8SKzvmzbvaP3eP9aGD08X3GgtBfZPYn4AYqawOe82Xq
G3adq1VUksWSicmCBZC9cMeM/BTzQl0uqPuBMfI0IU0SQCKE6URIwO//RxT5cOtK
jM5R+qLROw2DfPbSvUB14RfJuy//T4pAAJWp2+LWWQZ23vMudHfwoZTFxo8B2kel
KNyANQ/jDjhgU5Zu3Sn40X8zaQrVz/M+i0BmTFeRIafreO5/eR71p5JSvHjVxGro
2l59sR+iSgcWKgEeFcaejOcl9kWqcsEiZchnllLQ4Y3up5CIpD2NRhT6rtcBMhJk
67ozYMKtZnyofLVvdEGDt8QSuxABlZpZ9KSrXzR93DLGEnXi1qBS3G10jmPjfL2/
FWwAIDwEVdqfuMXw+xhZkLlJaPADEXxZA/hdwrjN8ml6O8LKdQ/XgD/9tAu26AAz
13I5WHz13E0FKMPxP/wt5Gq+t5m7ARR5Ij2CXkkrC57djWmDjjbApAqPHKZROGjD
x1oPvYh6bkKndvQBc9n2LwMnuCfB2oPp+2Reidwid1gWQmssSD/WYDHnhyX3Mc/F
elx7H/h3FD06+4CnEsxY7fwP7zYLw4Wz5Wx0byuHY7kDbjfqicMyTWu8GQThD/fY
g9DSTvwdL/DTiO2cmOdu2tFkTtB3eQ7rn/dGsSHpwVsvOPFyKfPOM814jAhxO6VX
p65HSnZb7tQA/3Vg6uzkDR5GR9NmlAu0WkT1nTP+ZRbTw/b5R+0Klv83yoXAQk+w
uD6Vh0TxrJVsp6VWdQixyNicg11SjOE55ITXTMseL4ygXdrfivLXbvSusNsZcO+e
nm8ET69nPngP62p1WmaL/p/pDqU8QcovBQnlVI7C3cFtJgNKEMznEy8I6wRDi4pj
fGj+TEkdgf1lhyX/gekd6rBmna2QOgs3gUQAdj0wMlw+WZnHQs/pVO14ULTtFAI/
UUVYzvmAbsAE6DPLDjjdQ4Gg/0XYzfNgGd0SkBZPaaQeOdssaR5CGtCT7FQMyiq9
3IUgno5ctFB9C5OSK1nuXBMLkcapt2lQyjkl+J9Z4HlatrbT0MLTiGohEkEeLGlF
QBARbmcp3G7QiuhJrML7nvAQ6TefkF5/KLccwr5OlX1Q6PRp44S5kq1gq+Y6boAp
UpqPqVmR2u3OVhI/HV2v9vZGk83wkn4J4964LMg8sGN7mQb1zgMQu9k6JuSpVGhJ
jRQmzAaczdUlls3Z+iq1P5nrTZldBY+SuapdP6kHwN+EK8KRgDnY1D++9kvCD9fZ
iEr2DFeRh4SAgvO4WrYle40AERZrZr8+f7XcGiiRQm0stSxAhBgT7QK6hyehM6r0
Zzk6ruMD6jh09aKfuvr3+duxtlCfWrujvqdkvW2ozp99tnY7VWwf+AvVL45otTcw
roMmtmmzGa6+lwx6hkBBYSye5ICeST9yi/omSicPGMAAOD1OCJqzx4QjBfAvMdMn
qtUC56i8T49sYaQxw46GZeC8SxUia17v/Xz6D0zj1wAwAaKQJ2VL2B+f6tWkbI77
2IRX/lF9laYHs8rePIr97id5NBerkUBfVqiJ3F8A6IysFV6sSY9HiyB/jJ41Gy8o
dlTKMolvMeZHx4NTj6Xna0Qb+hZX31spx/ANALuc4Q7F9LxBDxPtQ4Ow0aOgbrHy
iRR+7Spq/YUaKJF8ROc45ydzf1Zg8uvr9LWBB84p6px/99XIDrTS4PAh9CoyYf7f
lvg6O59sijLey5BJgF0BU9bJunzogfFGthyDZWcV3l1nW+CziZ6Kq2+p2aHWHyE8
MZoNk3ezbJI0upFAuTjxFLuDuzrvbZTsFunyGf+hR9c+6sM1S8t4k5Tp28Efit/c
KgU3tsX6WGMFFw29w41rZeeZsdhdQ0KukH+WZVURzZEOcvmhoW4RkLaGqDbnVnZo
4aorm9X3JDjOR8HoQaxyoiVrcpbIsxTWbUtEHgnvRISB9W+cxlvaKz8F9UiIvigh
x5p9MD5ZgCgoAdZskFegYg5wEZ3rBzHdx9iikDAGTh7wKO5bdkAyIqQyIoqaC0Yc
1BoITce38wbgF0FJwUP5LAuEx9uPC7HltrC58MZztqVrhNsQ7XBOkmsX5RUAV32T
nNgQNVoN21/doCKOtfMYDVqx9OlF9sNcBvQ+23eS2v/nlXKsx39bn953eSMjYY50
EtH2bd7yhvwmv7oWhuLMFh34LXzvNx5VkFk2LuB3/YIF7uFxDVAVwKNYvYRIv8tR
hBc7DP+tc6T3U451vZX3BPPKqEOekFzcNBxg8r4JXgESR6q1uTTmfIyJpTvS/kWN
O6nNo5JhStz076stma2GbbPR0QLvE5PLHZDmBni11KbaF7dWbCU2hKEy9NnirLoc
75ADqebaG4J3uUerHQjz5eeYuzsXjEwuuVjE8XauziMHYSIZLUq8DFnD5zucKDLI
f6cUaWhIESdyJSZR7pjNmlZSO9SdGvW9WBgTL5sPRU5TUNwGSAxBZdwUyaND4dK9
7gOhl8mMTAO8liEuBV/wdvdkJezeT+MXAXpHPJzRYdh/M3ZgTp6GIWRwVP3ivse0
kGu70GlHs1PwlBk9PXc/x0kBhASFNeUxfOnsuv9UvIA7YM5hwnHZI+3dcB/wdyeC
XZO2UCDSs9B9MddIS6Mry8iRkw25rZ4TbVjOPbclH7Z7ALZsCPjOEUbcYLjp1BFL
+TpNEHSgH5V7H8BloR3bjaa4or+V4XxMhi+ixoyUJiG4mqChOVJk8AjL5OgJAnWw
PJwwD0mb90FzzTtBe59JvRYeah/73fH0vzQEdIk+2de8tHjxIJFOxuEIIjh8sTR6
Jit4jsT9ZC92LOw3ctUrH/iFsLQ7P78g+62SL+nW2I4+Xp8AInteAy+YhlinmbJh
ksxG82ggCAeHQKWjBOYclhshF13fW3am7daMuP7NDii7LYjnthJZkj9TpO2mvfkc
OjkJ2YBy+QNIQUOkf8YBSnzqRjVDpy8TpLL66H5D2M5c41R0LXp2/kjis7Bbusnp
LfOetXvvqBjGrwc5FuPimoJPHIq46T94S/acjO2dLj52P8pLd8bwfpdDRp3KrNoD
0xjoLvqX9Dfen/Qrb4d/ZwdO5oVHic/9RJoSQmeLVvJroRMD777438PbJOK/uECp
mnkcn1NMf6oWuLs7YwHcRDTXPgbyd4kNISeJ6XrMjlzHqIIS7kdmVWVJj8X4IfBL
lhZteh1LiyIRUy+SUts5PHAX8hQrQ+G562lGZRTdZpLaNmZHpxG8m/rl9ImBaoNM
khMPEOsx/y20vtEm6KyitWr5MZYCVhjQSv6fMM6a523coEdbYt7XpGn/FkHRPKVu
Cu/RWhVWwCQcyPm77BldYd20AtdrIPw7icD5eVXK0nzZHUhz68ZunqTUGlwuWVlu
xo202m1x5WsSGfotJlEVvk8n+OKlMrBmh59JZVJFPIpmkGOD8V4TmzA9ofN2fHX3
bDpU1cpsn59ABR/qfDZbDmdGeoYJOjPadOj/P5g0U56xii6XIsCF0p8WmQje2mTF
q8OyBeKTuYSQkMEQtlP1Ei05Yg833UQmm3/7lwbIHvmMA1X5c75UMStSlV5eWW1m
hU6r1LAiqJSuWcksj8l79/lD6/QzJE7V90j4W8nQrOYEt1HtDu9phezfNyCUCQZm
QbJYFmpahLNhKFiNmHGF6cTJ/O32gacsQR9SDGhnMEI+l8yNl/0+XilIUuwvjBA7
7lsZ/Mp6wqX2eS9GFL0R/DUUQAluMY7+xb/wFQN+qBh1Zq217nfSEN9odS6keJhb
rKiOG7lC6lb4CUYqn3lVfy65W9gGGI6R2Pbgq/TQwyiz8zOrZ5jTpuRbKy93iYjj
HxcMHapjy691QenQRw8tQlgcEOIpnL8V2nXf+cK5LIrjnka2rrlealSk7gnMdVc/
F34TLMVZ5cgYJhhTUKfdo2Mc3o/6QzB5PJfl2wr+1FGesDWNGpjGV+emfPG2ViYe
zTHN+WA6382u838fE6HUb5tW4w4lZuefaSNi1316JS1/BrcaXptdGk2YhUbimL0N
i3zHNRJBP7SNtiS0/WiYtGkEjddDhB7NBUzOk3iR+IklXa8wafX06b7xN4p/v2nz
gXXowimSq6MMPQXuaw1mJXCb4y6JsHw/NwMXFz05V9krccODZhTmc1+p39ndmUAP
hF+Fo5cz8mwlpWeRgJaoPL+zs/IyvA2gUUr7lZm0PsNAsWpTrL1VJsK9H6qCGQsN
tWSTADU8uT69wuCUFHglcEBMLScn8RR0wcGdFh2kV723JjTtMfXbfDq21h1Pg7ps
xBMFJ5ajO/4N7sOr35uNGumjcSti6CUvBMEGdeGAHudear0dMUDHmljEM1+OkE7F
4klgkEj/62g2RUI1ekhpptjRBTuYGPb5QdygZzf3w5ud4zZXt7LtAjJ2aRvQ2CA8
iWpN2W8SKSd9M9LmlTEvn9LukDunWCdjld1JR6cLdyBc8BhjgFBtxsWXo3ggVuhJ
lb8WxCSygYJ9ke97hPxpMoOPc8A3JbFo7Y3f9Tr3Z4WlUsuCoix/QyAOya9+gitO
EZXJD6F0FHsXh79E+z1slZCd9p3Y2eZ3gc2GfVoTs69dwm7q1gKU0Ga9jXTyz26L
ow4rNTcjuAVwW+mAtqPk2sRgFAGh2Kt+QkUaQLg1Pq/RgTphVn1uJCHNZAce0J7u
6rTmv4Az9H5E3dDGJXIREdhK/1lLf8aEgi56Yvs+9uGMMjhuAG8w1WGFfAqrhZUI
gcQnttZu9Ou6EFi/JTS8gWKex0+ohn836rqDnXpFiIX2tO93SwV2SAsLjlxCYhsk
RlqZHLAdkowYvGVgmoO8vQueRaKesDxKok+dBwUz4ZiiFCFjJ3t7LiX5XqJJPllq
5aNG7IsCgKOwgeBygqog8zPS6mPTFdXxM+0K2K4SMEG140e2YyV1iQIKw1Lqwztn
v+9bbP1MCA66x+vr4OIs/Qxc1yQ8JUN/SHJMULnHsjmjUXM111lJzXEfDGdxfR3d
Jbo07qEm8lETtMNr+ACkUg2nm9Ia2ok5VUB/9mVjrF6zLAaZ6NiBEl/u77q0givg
l7WLSM/C2VMEZeLb1AonyEMZ7XiK/mQIcv1FaXVSM6hEFQfAcZC1JNLj+NG3l7kU
M2XNN11MSvgW1HlOadBVYXx3cnvclHLUfIJuFbMg/155cFMEyKbzx67bjpkFSAyq
UIAAHx2sNv2Sl/R2lgDc5MnrkMDILefbZQwG1qmd/252B1+xpKsIGGw2MwLngjKz
Z3+kMeaqabVITN+GHVyTAU95wakSSoZ86HM14tabCQ+lsEYj17ZDg6yVR9MV9K4S
2MTdj/ZCxYh7E7LqTEVwCEaZCYD604QE8ZNRDnxhIAwwqyl5ucJPyhUuUPG7L//k
Eyi7jmXb0r1gLN2QimjN8mbhw8ihd8UKdRunfwsQDfRki/t6nbc51PfouPjkqMXM
nPGFdYink4IQNrHueCh5hkfKKmYKzU3xATE/OHdOl1bQpsDfIF2hvAIM8Je5Q/yc
8lMFf+1OqqV2DFg5DU3R+xdDzvgFw8TcAzZW1rA6i2KF215ulmDRgTwOSJiQTQLZ
4trAWyIrCSn+zwf5QMnlNRzbnrsh24/G9XRefyvJ2RPYi40FJaAuQ8CyqKDUlEF0
Qkz3U/rZl/y+wEzsqzA+6+H89N3xASt7+ySOoKkeRdAm7LkKrmyWhqfhAVxSi8Cl
+4bZfuWzRxD1u91KK9xA1wc6g2BDCQLpWL4Sih6EGOHBvA2MBiZwtLZVOHz7zfWN
t7RT7myaQFudhAYZ8y5HULH3pfvrKXy0TRruZOcIrBWnQtxltoPu5RjUYThS2gIU
hzwlzvmym98GdTN3B3B/E32qqTd9PW9sPzpuz5CSuLCwaPuow0nXe8Gmc4OEwVsH
TdBKdRuiWciHUHaoSJO+jb8oBdQxBF4Gzn7R9sK4eLnLcR0sx9g+4XKXX/OW4H3a
ZZmxTOzGjg36GFO12ABj1OsWsD7X/lEs7Z/+CLUcKMpTxHBQZyAxgJZKhzZ7Fv+4
m1ZmPaVY7g5QIPbdY/gmxUOsKEDxObqKqwimeNMb89A2vL2/9cTvwW0gfp5QtUHs
Nps53gXardN8qlv1aQQpn+QJPHXmHrsgOo7IYObC3HViRW9aw1RNuDvRoQmco6U6
uFLfg2Ir8TqxoEaIY4ivha+/GJ8C6Sn8mVDHGhZZT/5D+Mnv2oe4wDVWfqd0lkar
WzodbxeqQli/3d5+ORWJ8W9gp4MkW9q/tH2Cur/6bPeTtGgrW3o4M2gQXdd2sETy
ecsBufloA68fSzf7WxlIP5wQZ4yU9QnlX66J8PjFTCQco9k4JT3h+2gfZlpzO3ME
tM0Pv8CpnXInVxUk7O+FHmX9J6JVMg4m5NzJO8Y0d/L0/URK27i8zUpE5Z0Hp1kZ
k/1STQYqR2ZjYfaTSxEI8gvQNzbRH0UNglUNXeCio1cFDNp60TVtTMm4tm+ln3lu
3WnkEzeOtlH4OtI16XU1cXKeupcm4Yc5gYmclSPP5iHGgLqo72NNqhRMQz8ukhQd
kHFdHW+GPbkX/80GDmaQWg/1m7F7C3gsS0fauImFQNRUYckUdB2U0QTJFMNkjgwb
8yPkpuAnBYHtqZlmDQjA6tjdLr+giAz588aq8lVViCamDE2WrC+Ux08iB9ZPFFNR
zmOjAZJlw54xroXcfnEbarhMF+JODa2W6kzb6W36XDTZV+Y+TlZr2iJE6t+SIo8G
cIJUtM30RZObszJwlYwA47xQ3kzb6DTb9Gn06Xka1L5t1Ih0kljyUIri9zUF+F7v
/Qe8Unwku/DuqFXisfiJ2H7asKfpmBXviyvDgVmXrFSXNlrzT1a/D45q4vUKR/R0
sm4IUgltRoecXcgotP8noYfcYBXl6jaJJaKYz4oKTInnQBJtgVA/AGvU+wwdKv4y
tJHTxZH8Do/ZIIwBczNNLozcECxQpe26TQLUqjICv866R50yJe7Z+px8hoLPV6e6
x6IRLorWXq8iWEg0bR9YQhfDAO1pz21yvSrUqmXNnMfOG7+bLcTIgup3fl7s8MZk
L8S5Nw6Q+mwY4BWJVnKpt1Os1mSCZc9zlSXFFscixiIR/PP1cpw0a79uCs1WVAYC
w9BbIzeV1haRA7Bwu9RQRVsS4Z0TSR0esvRYe+a0tWDClGi7cKyqE7k6vzN/LvlS
gUixAbOJFIcvIPz4Y+/1yab+uMQn+kXaIKSeYyZOoyxlUbSJzZtUwmtGCvUhSx4M
uHrpxTLn2EHz6p68O0J29ndARhkiBam38dTXhIeamhxjj4tEDHrUujVjkb6Lnidp
tlTUWAue71RA9k5QQHWNggRJLE4mlobKCSQRKiA8ncoSJ7tI7Fc6niHAcrXrWfj8
swp+arj04S/W//VdtR2BhNRy0nKP6Efg+k2iZGgU4Bt0S9yDxbK+dbi/CAlwLAjm
k3cDgXhPonFBMPYQF4A6b85KWo0z6U1KJuD/hYaBItp0KGplCyhLgVklpTr12j73
LVg/7U+/S7nbPPpqhQ6YK3saxmD+dJKWIjBXnRyZeEEA/yHTqQRhe4HNiediV3cY
clwXmZMv2SCq8RhjKq1TZv2nhzzQYctYk+ff7pS4T7xittk5JfRNhG+3tO14Nzz0
HqnVs/r/+4kmIJImKjLWSX/mLm+RmmEwTNeDVY/J3tF/nhmYoVyAYJR628dGCowC
rgvHXljJHjf4VW2fuYFbxpEbqzQ/suayJ9YSco3zsn8kHzV9Ta3+7fFXJ2kQ2n1S
4C/bwebVxKqXgeI0dS5VaEPFnV5ifhSB/Sa1s+sWTW8A7K6WUnq4MaEMGJp4fka+
URm0aUMKvLvmzqtRfw+QnyE2HuVZhZ9ei/C/rmSDg7ToJs/2G2D17VeX9438NEN8
qeTVTrnlFXhcZ1x461ufhNDYtR+W1NK09NE4k2ltum+iyzfuzK9aB9e72SqgKQRE
dflJOADJK3EjVBnOrImhzZom+wVKMVlHTT3aszXW2cJLxJXpof802wI/Zk5nqqlo
5qABJqfsNDARpiBUvp4WGNKnOiFbLu2/mTnXWsC0Q5KaLAFH7RFmRQEyIHnsxTzB
B0fHDna1BU3fG//v3IXhKRis36kdGDrV2D0ROFiF7VYsEvzglwK8HrWyq26kwR6t
cwisOzaRV/thwVraVwDR5tkARXheJ2CZRkmtfsV4sSqodFTpRu7TaEUmkZ5euWvG
0rv624DcCSJU6bBx9ucY2EZntpywpHllckNuV+ufEwAHqCS8xxFrY8p1ZLga8/vB
7FxkFWvptV7OoJWFxqjNvVV4VxPI+uFaxd4hsMhy8enShHLBNWXZ7+e9YjYxhvOX
YH6Y0ipQZpTBs7tnBFh514jZfu29fR3RoZdcrh7BCW7SKwkXfHZLojP9Uk80C8CY
1V385ZWa8q1KBulpbq1EjcgvGQXEqmED+1OhGGTNdzLpB6dEULjSHrNTv3H5xzlm
u7ttDGLP7avUAxb5V1uJOrTEpDephAnLN1FtINziR2zcQI08iSxbvY9u3/XCHGaD
81u2JAI3IsAQyyH1L5ArG7y6Xn4EjywhvAatGqWihTWwz9/56xMKTa2aFmDyqIkd
G7kddD5tDs/dQM1kjqidOfVhUBkdKZrQeckM16onkvFGs5UzbSQUFs6L9zN7ft79
22edzPomNgTm/SpeCScw4uiSIoDuC1mK59KadAkiEfTPPEh/WYPDkNundAlirsvT
I5s8b7XAbGjmmWHoXWPtifFpUMYLDKAIig76Oan7KgWfstPcC/COFhiO/0l2QwvZ
BNqf9O/FfCqiY62Gr2w7JR/qYqalusjPrchVrUQ2gz2GrJVC83c4Lhi+ZBMYXsQQ
1v+7Q9h2eQuTRHthdexWCobw89wJ8nz8MgBvQmGOde5G+bYDaLcio3JDQtnN/4B1
zWi7pNr5PU+BUgNty91JDiEqXw9Ds/ZUWt7l2ELBMHEP+1Ce0WmMhZgbaJ+WyLji
6JDufTdLhELNuJ0YCrAyXoQaOwkgMZYN4H6MC2qPFD6ZuC0RRblygqBTBICo1mer
mWavh3YiS9jTMfpItdszUB9pUrvrqTcgpGQ43/R2g3YvaHOTbESwgHq65FWT/+Vr
X+Zdzzk8EjCa9AtNa58nIsuGhQPQATllIdmne2o4q18YRD6swMf924qfOlJ0GwGI
Bw6rzXRrjEO7KglRvEjV/NQXy4cUmvVv75k5zxQZX/zQJHOxoO0BGGesr642/ECm
5O4J79K60D/uT/PTogeFKrSM45vThSYzpP4feKDHd1pmeo7lNTQC6AgVeAj1LhDX
+Y2ocEPt1BgyBsO/1Z70rtPgwx0LHKkJwS8PXjz8VfEcuu0/8uphsCleFlmA5KD8
sAzn78Bg3Fik296jiDkTyOja+jKZ2rjE3lEnqPVluJTIHyEkxB2UbGD6rEg/owfq
ux81LUO+/MH8Qtk3A5Ik3/HSHrecZJChvRIqL+YbW4g0X6RBkEgU7Zo7Lp6Q/+09
MQf5zgfQybLDPOH3Kw+PKKmMuI/MiqfmwpWJcO0wZsHJ9fY7FUW0o9Aq4nq6sUwD
DjebkNGJdzOL+zttv6pogGuFbQ1oudogHA4ug0ca7fv+U6KPQ2RNVj8eRi2yULjh
YiDFxD9gLGxaGmMTy9Llg2Hf02M96YtxJjBWJCjaGalc7TnIqcq8CMkGLYnb1BaR
dcJ48IcLN6o9cRFAN0RvUAEqIWvPf3dN8YbzW65+qE4wxJ0D2fFz+W8PywRQrbz8
4AVGuqyMA1Aqb75N/ROGioKK624NL5wh1gg2qWftzGOoukfnPzSREFNGjofn29AG
txF8n3hIvx4jjypz/2MsEBJfa77iNFnHU/DCUXRANd62t2ltZBRtonveWlt7NoDn
XbDX0vi6Uubhlpq1BqJSuKih/tCbxKbq8CKK6Q0Pu9UIrDOhCWAgsVQ2pZsypJ93
ETuR54Enkslc6tUDJ22YBLZy/P2PVsP3DxnMkJgbV4e5n4TleosLNYmSmorMtaqX
CWDDbm0+3lL3RLgG0d5fzlk3dMbP5T9v0RSsgNHANZczABlt4tefBD5xd3iC/S2r
doDk56XYgVNphMAVyyF7ZBFSSKWNlW9e1rDIVaUqHlp8WeQ0yWhV5y/f1aSJjmzd
zSlJEd67IQ0WVWdspzwDAxe61Fa/p0IBGBaDAHLhcsy/eunCkW2flSWUCqzW2y7y
e5DMiSApOZuJF+57HrdJnlksiZ9M2Z/SN/mWbJqXVFBpupJ8ZhnxZR8YFqu2hw2q
8QVBQytxqrugEP+kTzWaUkI7JwxSprZNm5HG1HoB0YSa9IhpZOiHGzigAzLXdYmo
OMd3t/6+Eaz2kUqlZisymSWnCJGsFXLuILO+qS7VmLkiyAufbzx2965ew9O8uYCC
beWP9VUHavqVmZvAZttcAc83Pa2OTtoPLPy+XJj7nLCZH+BOTIQj9QqKKSl9wDBT
IQgb+yPzZxPdqKGQkjvfahrma0gOd9UTiaU57Fyziw2/Ng3bOpFAZdd0ZpR88tjh
yAOJbjhk5ybJ+gl3RpZIjnV9dg3zLMPgID5+uXn0P6bPvALBXymIXsnuBOtnWOv6
b5DAt/AJZsKqAj91enuMHpZ+rWTImWwcGmNcOgW3hiV4vlv3pDwqPuxCWJKZ5Ufr
bDI49x/1EGRpdgq7w+2h8WobJdjZNsYOfaOXobH/iUanHhYoHPL5R4t3IfDPi8QN
wV36EaLpSzblb8SK9zaF3XHPM9WoIPkqjSkdS5AfEm767kZPmnNoDuZAcJvPUypO
WQ3xiSvgJ7N6Z4jC+FijBe9TcYdGRgVMFrWVM6enBtIZhcvOxMTrxVRWSc2cDgB5
L5LEx6b0b8zivaOwvkd9sIeV3lLpzjORZ8G1MwFrp9+S2JM+N89GK5wXv2gXOpe4
3stoVP5/EsTwmvM5hPPFtSngjuG86nozzsUkMHQxNLeUTpeODI2JK2lXUWDebLod
PhBjZTIbtpST1PZavtEihYRV0SOkcQU/dIH/xV9QGpgoS8Nt2KuflTaWVO5PklIA
B7muYC2Y/gJG+zEwl0VugCV7sH0YJmIKzRB0KFKyxIt5X3t1ZD3E1g4iDxjtcy8Q
/mW1m9DWAh6AMidIgIeH99iJU3Mt8tH113SRnTbQ6DNac5LDhuU0aLlUORe2D/6g
3kRXYiBE8f4Q1x+MYjQpy5WkkxqniUg5RZMNj7SbewVlwx+3iOqt02XCKVkKOS7o
s3Ks/aEYJNFJKpJFsZMWgN5Zd9ouTt7aUjnxQnX263hLhbwcLhXlJwRw4noUTYYe
RopWAdJV0WDR06hrabPjZSj7cAIgQ1lmxsOyLE4fVy7mgM+hjtd4S6JVP5W9arOY
vN88fWgxfHqOT4mn5LD9S+xNl6sYImtgFZtXHYaT8DUGEMFRNjuSq8xX8qOnQZ0q
r+RgMh8d2GOjbwmUQBzCqCT+DDsmBXlJHSfASFByfniH4fAM42aIssWC3ALVj5BZ
u0DLhpwuwby9+Dl9KD5069+Y1zl/qvtyi3NBCVCPZS2Ud7daDid35TiCIzyxjgOJ
56cwG8ZSD0Iq2B1A8DqynvWFJpHAkzmFqMOiQ7JYP8r15gc45V/PaMay5t9KW+OI
RVlrhhg+qDT75tYzbrx0EI58jhYkJsDI9/2BRq4hmo0SYpAtOqCki1kY1VTGcBwn
hJkU2l93fu+jeGgcQJvkb7xXleclUkf3tlHTecCJbDQ5LpFUdC8g1box0P9H/GSA
tg3AAUUuxcPcJbjZWQUC778YryObpZcaDJKS7X40gww+MR+w+0PlZveJmu5oCqKx
fgya9AtNw+3X99AwUuzWc42thrXqrKD0hv3E4TC+Xwh8HX/DV2YIGfqrUGmMon7A
eyWyE4KXQJ0urFx/PFME0ruofEOUmT9He7H2Um32rPAO9ZGTzc0mWPffNS1bUb08
HJ/dp0xvKZqqTw1faG8lr2vnm0XRx5P1gYvbv4FUQtJb7EQZfm8dU3g6owXa+AS8
f0nO2PEkxEReW6JjsEBOMnsInu/pHc55MLHDg0OqO80QpYhlYluunST25CMhxKr4
oBlQubUb3k3msgKiHhhPTjAjKqjwU5Xod9LIsOVCyhHeNwwlmRb3xETNoZPQHdXK
aOcHhOiLW8GK84gJXldF6/JH37pUQMOPH/cz/V6Xu8lY2Z9RZUt7Gk64ZtrpNu3y
ewiKpKPm2jrYEZUsRpPst0YhIkh7Z2Vuu+ayMH4Q2+KhkaKH5sDmACdkBRxBH2yP
kWiq36kYRuGC/LUV/dWKd2CC/2YdehklbYwHmL/k5WVDLqcLk/PqTne3R+j9pY7i
rfSwlIPxueSmiS6bYx3X0AU9F0j/V6jT5kJ2O5CXl6IXN6YIvZ89/HQe61iunEA5
ETj4FLZXtHl80Mc78zguo6dRotYvQCr2CEWM5NJ6eZs+aAcvWsI/fKnpEOQuuqzA
1OejGsmuquR6B4AUTGo7CWZs1GJAaJ4wRSsCYCCdDqP6ALIEFSnAlfYirf0vRRd4
74QnRe7ahV3Ng724dvqnA3aUaBTvf+QtcMTPL2KNRChzKoZlMRwfEYwUgOMZuycl
5YCn59YxliVhSr0E+zvNgCmIvdT7cVggUG0EiKq2/OzpWMIfQ2BQWQRDx8p17ih+
tECFRjhbiV5Kou3Y7ajMgp+1DSPUMzM2PKra4zL2HF6kEqheoM+FHROOyvm8VmhP
uBZjQBQE6LRvb3tC9VZ2iyGiySR417JbJ56YRziDEp/dVWpzAMI7JuGXwGGz1uIw
O6vO95Sg2ykGuK6bdQecz3TxYtv8Vn6uVOyPzkpHJh1KaXmtP5HVTcC5kYH6XEwP
Ef5vyM3A0HqZO1JfzGAdsT189Hi+70P2FqyKMNqVl3FRK8enuHrWKBtoF7ND2h1H
u//Tp08nc2OvZoYfZEJwZF40ke4lCf+XtKqYAw5RRWK5bsf4lRQC1wJQiG8/9AqH
OG+MzgmIgukilvA8nxCsFJeDNGAzThclSoNMHi+C1cYZgyhLQZU5/n6S2AH4BSDE
MuAtK9czZhnCiCuyUBj4cMkWH/5WIyAPONfEArgpWjYy7wno9Hh5D3hvth5REhfk
2+B7PjK8EZgzGt90U2oIf8Gf4U0+V4TKG8LBWwZa/yzth/w9RtYXMKPCriwmHof+
1yj/cUx9EKtpPvIczRZmRiTivxnNyIdVYOnKmXrwMc6IpXfhbmTiBMea9QcRUVwn
pZ5XLA8hmrhXPurxsYP3CDRgQFWi8LW56b8LRxMyj+/rD5Ck/gp7VcW07JSoW457
6GzcREPWbw9D3v8pw1AIkUruTXJCRwdPJyOH0UPIWwkwtGEA0fgu/69DlLeMrAcU
/rVDD4t3JW4/9OQ5CU2cdsxgnhoZ8e/UW6Wm8N3inQGn3tdT++avZbx9ijkt1XYO
8s/pz/i3/IYJxI2ZrSmGjBdc+71RZAdK7YEdq4MlsUuMar0wjwmNvDvoE9r+aGuq
0Dco6lxh3bDi8RjietXhfenruJgbKCchN5Ku+zhvrn4m8IrTRphDp/K52+3tJUls
opjVznoBspXSHrDpP3vcOVnz6zi36fXoXpCE6VKNJ2NJMR16S7VvgYqcFeZsYN0I
1Z4+ALrNuBcKcs3SsMnZxoSmqNNGBqRMZrmccVyaloH/Y9Jxnr1shc6AQY6r30xj
QaK8G1AoCh7LiyVhhdDa1kGEXCqM6Lkp32NjY0s7WRNN+TuH9tjvIo3AYksU5Lmc
kZEsH2jnHNenpmyzll3ToMOA/kZvbNeANjBg3GcOZxRUh+m+vzZ7+qZo+zIfy6ly
r6u2Q7mztGA3UxxwuGKYoljVxABE6HZmJ4sX16nHXfVEQLaPSuZjvdaP/tzoIxL4
L+zxTAfeeTo998OGHIs40JFUl4OkikVUXGF/RJg+gF006883omqp+ekkv5ws7eVe
aH2yOtw5bJL4GeJmE7pYixl4WGj2WKtCKWbH8WfeYDzsAFTZwaXBhIHSg3WgzUKD
eyB0UKpcdqLFia/PTShQuDqo0Rk8kBS07NxUUGC63yKUfMrd6n4uzjMRUcNjofR5
FzBcjbPoWATTQFcsbf+yAkYlT5TYGAtdhK+HAJd2oGS4HAs70HvYsGj9R/BJJfnZ
Kpesmcv48a2gjpC61IDteu8ULeDkO6YDZHfHxHjfUn95fr5+kGf7Fevr4mYqOWc6
oxBjovFyMZ6dx+SYEvYZ75T2c8wuaXrrJYDhF9D3HzPrQiTmCqQQOmYHpNuVk3O8
+uccP/JEo5oQ3pRBgbZT8ZWwwBgUzexnVanXa51jeKQSHfVrqkRn7qZ7DnHh54Gy
ViptuYr8hh7/sWmBb4nNj1sJDQhGmwBDHw9GNGC7UHGQiIDl2AHeGvB/prERCRso
52cu1AgW4LhRPRxpsISE44ZDB+Q4YYnUkHr9SZpbM+v6VQGmxkTPs/7PvXx5mA16
GaQd3wh9FZ6XGBV7msc+UFq1ow+GtZwiniAdm0r2PqiOfyjBOfuh6cI0mu9t1fXk
EuVr8SFLwTHxW3Ln4n2LIujeNi+XaZ5Y3YOZMOrSGnvXu2tq7r3U/PuWc/3iMt8H
b9HWJ8qjHscslURjyCbT8aAKiXjOpOXgiiRn2ul+cGNe12Ku6atTrNKLfIv+l3Dz
nx7lWQTzs6FWDOLJodP7AQEZ7126dRj3qi3lTjH8IRYTK/koYoPcUYre92Ky4DWj
ftj2lKbTLptJ0Tjf8QwD7bQLx5cKZuifyQqk05UalqnKluABaGu5IrnyKMHGX6Qh
JpDJW/GDT3UQY6YyEUznzgJNzsCBh4w8EhUQ6oileydqKqQp7WaB4OWipcMTgkm7
4Hjivhzh+JieEVKe19kXVQwyjTFajaPtTOD/FEUtDAeZtGL72OkWx31aI5bnIk97
ruWR2B3HccQZovxEkSQ7LiWw/bhqycbO/6ouXvfUsBg51/xO/HHwjOf2rTcCmYl0
rGme4tgWLupXc3Xqga5mvSPROHrNzoBL4msDEB+r39gi6lQR6VdhtGEkScEimSXf
n1+Xto2gDbXNbbc/9M2M9391Muod+t2H5hJBhily1xJARm9HaeINWpEkLJ9PjGkO
sx5vgJVbkz4t+lczZd2QdUglTsekPPDFqcN0XD/DJCUiU46iVDwffrLoRMHkxVdH
Kcql/PEKDsIOUEtNuo6TaRKAogv+XjYEGj0XPh4hTGc66sZ8ap6OVYyQCgsFwziJ
EFRyLpSuySRMu33K/E+a8wipcWwxkW2hsfvTh586Sv+H55fHTlQcnh9T3PUliFcJ
KjVXSEoskuD4lIRckXo8VFvODb7ZpM8bd0w6fmlKpPjVFVlFuE92/1uGNXoYWINg
zXwSvthzOuppURbWB7h4vSKxhrUgX+UVOgtnqJBcl9xu6qrfgT7e2qfF6t2Y9x9Q
cm7Tv3KY2IwSyziDfKwVZQivX0aBh1PR7fWa4vdjgWYUuYA7mxZE/uepn4b4KK+/
+PBmtPZB96pCRP/GrdtVZC+55jDs2IGy6M/EsvhnL5io506BDdc6S1SkW1KZ+OYK
51Ieb30mcPgBRLdTERLCjwCkXN/BK5UVAV61AwWqI/41Vh3kJwZvuBXfHH4uHq0q
R7edBbOL5Mz9/x1VyE8EqmCgYdAPnukWhys7lsTNMtPcKQodevnY/6efvLp5kDvq
Bha6mAroyWTJ1xUM1jcBOfjYfT2hcW3HFM6G1xl0ukx46UkCfvosw1GgVxqp296C
FqjivIxHwhrDufziSFSMYqkrdlQ0tNu9HiboudoxdxtIh8shOysyGQ/HPJqr4cx1
8apX9/wMaCZY7PxzL97l2VkjdRPuU1lrr7iX1HxEL17n5Fi+exYwQ7FIoxIyVSgW
klKX8gSjtc8M5tluk3Ox/PGZvjpKZdTfmaUN/I0THOyJZJ7GZ+QzyAw6mLlpU35S
cyvUDwkoqAKDZgmdBsrL0l9lDoCxMPV5fzCYWJuZscXnJXeLFNYTiHpg94B6KLfR
Z1j0dWMGtCLOU/pbPJCFWgF22I7abvJvtNYK+g+H0GXQ8P1uyzwS03gMayLmgXUf
nS9J19qtcVBzGve9x3XNptJ8ES3P6DeGmv/M/vOR5THyHnY8mhg11o1pGXkwNSxY
gU8ye3qAK5MIbpJBD6mQISkwfbkiqdLirSSV0+fHPEhR1JqrIBQLv5UvXqnrxfzQ
5oMMwxJsI/P6QSE5aFPj+KDOv6O4jU88ch5dFQVKafIfzR/DiwoZwI2HFT3a5J9Z
7TygDGzAhocYPOzDUtujBjcaM7WWUbUX8a+RoI7+ovrcRg/31KSeu5/KS0LgMg+f
5J2dSciKf5No0m+5S0geWC+OlwlsVYbPkLpC2W+Z7tc3ZXORLstiwGsD6z51uDin
jt/aWxQQTGakK+nVebppcZT85H9AHIMeBukpyq6NBmf+M/5cfzUikI5r6MHCeHjX
vAHV/gfN/xYlEbPWGZsIwtMmiNQ8NtOUlNU02sAQdGvts6xSFHk4S+vrLtiosrlM
0Jsh2D+dl0rsH/bG7qwj2D1s32qy0T9/kwo3vdFhbueKCRjwUbGmUF0I1kwNG+iM
QTVg33l9ZCNTlbW99ie31V1R8pvOlLbm/1kBhD6L6yPGgVEVW7Xjx0NTexdgNLa9
BCdVv936DMA/48dOiq9BixUkya2Jd+ObpHNPEiXrU/wm+vEjV88P2htOle5Agwc/
bEknB3AUDMzob4bfCk0NXnWuPkkf0WrEIhAfJqhkv8NhpJMxHxjmnLONAFq95pEh
I/YtzyMEuGpjYBqRPOFxmBSGyOB8QsyScMiH5eZ8wbR7tsaYuNakTl4yTMRz3Ggz
ioDQTi4XcAdb7TaZLYJQNn28RW7MhpqnAgiC6yi3SovHIdo5xrMhZLEvgXIH4Plx
lbyqyxcH8sQV3+3reC2HIN3aOPE1yocuN/pvYXzILdDwqvyJ8ELzOKqSgHJWJJ+D
g2vSdN+DzeptZ1aiqztbhvrXiJKfHIeWOKDBYDXAMYj5TakryzRzU05Kxk/2A4UU
uTetl1N6WyGaimNhQotHpgnDOfqGAnrde/N/UcxHWTH6ER3RYNzfKjMclweE+66G
kzh6rbftnDVsD9LTi3jkEqNenCAaIi+nw2qIzZazuwxvTDNZHmqh+RYGVB6/SjSi
XOPfi/djyt/Mqzkr6B7WyL/x2FDKsjC++QGZ9EIIBNPmuwpNQvIIbXw9/C++aTwf
VMPfY2y2epYt3LgGnZq7On/W2Uj9hGgHy92OlU3CunSMjw1ZqycLO2XwJij/X7ol
SbEMAVC7Qu82aJQh68ioKZriXe2CoSqkpnyaYqll+AVTYweu0VCWF1qGtGFG8Gd3
Dz29T3gkQm7eHGz16yBKsJXwklLoIGRXojbU8RE5zxe91wZv5z4cW1YJH/TMljoP
2LfS9ImH8B0uZs8xaWV+7pPOVf+z2eJ9JwQ/yRkb+9iqubyIZT4MH9j2D9E8LELz
l/gP+FSvSeAFpHTDTpA6gJqfG+9o0YxxHqn1/wpoiqmlyui6nMr9vDsx11xHXQ/8
EEzSTdrV3EIHOs6bs1DCArG7tDN5tHs8ue8uAtLIMZNcWjPPUm02jfL5v3UJfLEx
4IHYhZaf1D84iIFIJp+kiARze0j/2+wFmilDwy9RTvRhO+7FxWwBzmqmjLLyVscb
EmWFtaQc0oLKkN0fn+nOXOhF9/zU0ZGAZDIAwAdALWNseWaVeoJoWibAap096TEx
lLJSvE6t9tqLE8jXa/xy2iLSDn7VIxPZY2pVans+/Kgbx9NrpAKepv9HwHS0FbTc
NSTw3j3LVV07yrqUlnPHa2wvy8fyIArUiHwMBOl388LPsHl9l6568RNsW8WlDMGn
NzimEArk3il4J5WivPe08o8hxLGDXW1gxGVIHONjlBmXGPUSt498xGo1mMGF7fcq
xQNhLp1Ceqk6RwNuyCjf5nx6k/M43ILszM/eHVebQgDcgpu7+ZRetUBXiWaW1+sc
IgyFb1vJMusVqIeButrIzUcU6i1ii/onD8X0pOUvQS5WcyglMGbKeBVs54L1cATs
DVuH3GJ5+0NClrTkixG3p/IXdZvU0GqxbyTG/FkbmbRHpq7v0rC1iir72vnyCxFx
opZXmd3n7KK9UAstZ4R0HTIGmx3nkq5qgdK46NFZsZ+Q710tkRt0+tuivown9WJW
wIfVgz4914xEcdNqIs6NwDSPxMrr1bKsf1CAV87j8zK4lTnsIynNPhzR1+x6TFJO
OT+gGySJaxGMrNwiA3pLRYXlztRWK2LSvyAl1B13hr2C0LQyuU4k62ySmErPPveF
xO8ygNMxD8wM9mNAC/9+CDjhGnRtHFWlCXd30wk44b8uR7HWsS5aEH4D3qIWrlWQ
sUzaiRsJXwPEZOZvrCmb7zsTcrYlFm3iKuyHl/Jy9XcZcyDu+erUbHmAvPwv+MmF
BjUh2qIIB+INT9Qmz70Rso6cYTahkNiD39Uc8SgAv+s8uBclOAUWUv79fgPCLipx
7R1D/SVjCW58VYeJEFG6uZE+RAnLNZOP/dSOVnnD50rotUJoDuaQ8+F9o0uLNNPD
+94u4jv7MWH4T2Gb9oIIQ7YOUB/845GMGb99onvcorgVKzjHInZ7EfHNaKLB1AuU
WDW6Y5N9bVBlyYCMw7O+1I/LlWYxYsMbTIdAjkPDxgpjHUJTPwPWxlIRs8wQ/B6w
XRvHsvJjPh+wi1fmkfBNc81P7Jkwutxabm3UKtS9V3zJVl6fFzViWwL74HbRzZJo
H83INCEe+tE3OpbeZGtdNweImG8kajJjwKti2SHf/qLwoDAgT203M92dtFuKbnTw
E/ngkjg9caif1zEutrOcRw64DLLrfuM6UeNvy2OGZuMoE4T7UHGs/A/JPmq3Alvt
wRhGZHxIFF/fXPPhEvh45V3lj3SyLf0ittx1CRgGyIG/t0sT0NIMAmLLk4wWRjaq
AYv3RbcnsRSdu8pkq4jwiUITMvIzrD1p/OqFEpfDoGtgMTyo1hMHFw9IBaLgjHrA
0J18MhRZVloAGaEs0ESQ82ejrddI4uB43f5/jI6oyghNffH8cDwRRdUrnY8LBPAE
PSF8vPKZQmUcXTGx332rLhWCRaoM9ldqySmD3ewEr3zNmj2s/cGo4rwq45d1/TDL
lTNpz/xB4vgzY2e/NfNogUUU0P03L64LbXhodywmY6N/5M5cUiKw7gaD9DNqxny2
BTXCAoFGRvF986DswsjFPUQXpIt+8dT51XqBbRlosvFdZfOeEB8oPvul/Y4eUXGP
dKwzf7h8V1oT0urMxaHFpqnaUW3PvTqNFyIUxgToaDCBSk29gWy5LK7fU6UYFf0u
BHlQOS28VmhSxleqG0ww1ZkQNMyCtGpxZtAKREdYIHgI8zFvt7fDjxmsPg+RaM90
trC2d6mfjwlXXlaom1P9OAAKmgPD4IxxZKrXlO4GeyWCiGeVF2BqtaQ4hSbO5Fez
mCSUlirqAEIX3ybn8B74XxuU2ZIE4w9JaJYpAIUxWgUag3yNSaP+EBpBMbUDvO2r
DF2GEyRgkbfmK84KAFq/dkv0xv6pF06Yk2V+Sjp1yfD8+y8C5wS59rmulsOF1zHP
/pZ7NT+abXFqhSRbf4y4cVrDL2zjpZDOt9NcFVk5P3hdLjL+OeM3AEpBktg3+eOy
spW6/sMqx5NrDDYLLrJMp6RU6rrIYZNje1cr//AawFYPUWdfPx/v/hvKRUBE7jba
PHvrX3uSZNhDeM/qP+ZGwTYzzB5Dv8/niWki34kkqEoCLwHJ35HDX1dS7AV6Yb3s
GcyBjvEtsvD5BW/bB4nZrXVm+q7Bv/F4XnRRfEvRANLXxElnH8CMeS5sf1abN3IE
Mu1KO8+ds6nCiO4q9kSOp24cf0Bc292lY1lPeLNoH8au7oT7l/y5scxx2ezH7PaJ
u6JLUMV9LRDHi3rMpSdRpcEWEiUFDoTBfxFpUAYehmJDsSJTuweh8f9lL9zFyosh
3NgBHpByRw8m+25/HcSbBlFoRFR//h20VagtWxJl1Wp7t+7trzW3LkZzKBX2+vYu
t0pNCOxh5e/NJ7yv4coGSIm3yAd6+tM6YS9yuJxMs1EGRVRHuS6fpWDDkJFKtUeU
zNcHmdgyCW2AXll3et3IV9AlHvFHobAv1O8gqCHLLr69It0hFloDvNKZXyi+yAmL
78XERVLr8FPuYX2bV9LNeOSwJEONTHhehHgVEzN5Huh+JMizWwxJnk+Dk0NnHxmH
XYpgsIrYyGfGCme9iemv4y/0IgPBfUhqKN4/WWbXMvKGa5bUbhhcJicPwiTbyi3y
tCKYkJWtBenM98T+SpX+pq/pqcXEuia6T0yWdwnPraNf2wF9cMw/IEtWS4XdhlF1
yrgJ/RiaFEudaeK+MvbS4RkAA791Z8cK4Eegd+PG2niIMPsO1dlvbGJ5wdqdYN3m
zKvndJiTa01k9xqO3Zpgj0CKBsu7/QgOLovE4Gjp/QJP0nOXFRizz1qP1j/051+k
OCbTskaMSG9ji+7MN8LSfXZPoMViOq4XElDDykTl49afwaP7IE7rWC64CSD2o5gS
9+pTCS8oMa1CPy8FWRAMnAy1YFlF2Wo49l6FrJ3sI0hxjzdr1CLQNrqJE/u4f9hl
1+eFNIGuDMknTr+O6Dult5smha5EJG3AWpO5d/PF+ejB23Dxopkgpjv3I1JyYOeK
kndhkHjBOCmQ+j0MnDAyRlvU/J6IpG7BAPDotIlGOKiE0Rm4GUVMZO1IYMC/g8iy
MjZ1nV+hd/HGBkiV498A5CZWNwcQI9yc2FIygbVTMJRR1+W5hOpK9QN5mmBPYeZE
2r6Rlep2NeyzxvxTDk7wvzuBBoXQMbPix3SEAMUPAHpDe9wzqwgjhqZPvA3fhT4j
UdOeUhhyeWQb32yKyja9+25Z9DSgLC2VjMP/vBI1upOsAXOUqR4sYUCTUVLRVtEQ
75hmF8d1wXoFc0Pwgfo5aN8X36tSLErutRaJ7HVxh6SDqpTcxBuOzs/Il7x9CeQf
JhtNq2wa9jrS3Rrq6g6taAgbIB2yclFqP5bEI/nkn3wiORPMD8XplbKRieg+pBw+
AWzAMpv6EhGmaA3FyMIJ7zOBNQvfSM4Sx9tW25nGJ87feYbB1X7foRE+3hrwOSTB
zTyJ3wU65ncel+h5Z6PVKyfnkjpuJ0gr4gVHh06p4DFBJm0DM1c7rk3bO9pr2Tzx
c1usTx6Q3jLAHyeH1SFxXmJsxSuZXARMA1mkE55fYryK2l0tx9jUeb8FQ3c0clJE
MCtUYaqY7ImTPqq1WwtfrD/p6VO07BNRzz3RckvHsd5rF1fq3CERRCLS+xh8tXzn
wRZo6UYGO6TrhpcGKej3H9HsUXIvucF3uhJx8XNAfBsdHpMFMhMZPfZ9ndWMDNbV
aKz11hJdsyebcSOZa9hh2fuKgFSJZ02GEQ8X2u8ze76rABkRS2LVsiRenrRS+Fgn
JdDpxz7WqlFzoE6pWMLA9DK64Ilit1b5ZDfzRyKx4ZxO807JswW5OSSgFyI2EBgE
xuQPMFWoxmlkDm04qT6c+u0faRvJhqi7oP4JUh4IYhQHB1xzGhEWeio72hiyxObV
ZLJKyIv93WWd+8a64bXE4yf4DJmbyJ8iF0do53JFMtNhGbRW9YJ3M8tGD3JJe2sA
Li2sq+zzXlf162HQdkPsObkiv19Jafi11CbM4ND4G8XSPQnW7eQ2F7vSipmwIETE
QwSftAUuAI+VFRaiLRStE6feEQ+Yx7Y6jdOqYF4bcdtXLjWxkpgZzcI+JTZqu2Cj
Fc+go/ck4t65tdCu6AclW2WJex2yZ4TUhxwJpIteyYhEtrMJ6qQSdYQth8VzGjCX
xp1YI7EE4GZFjt+mUoGZMwf+5QqUvCQRjJU9Z5DbDPFjsCGUoMEZT1gSdy0YnxnR
onkrGlVYEL+B0bbrfPhN87zGtO5O90gWQw4RRJccGhezKCSk2B+DFoOCDhr5bR6V
QnJG1sbNUlD1kAjCu4d/8O0XfCAC+NNoJhE8W8ZOv+FYbWiARA58/JCMnUmGEIyn
+twcJDbMky5eiaX5Y2Sp5WC/sgSAvwuuaO2ZmaeKXK0ZCFV1NYEBOz4I068ogww9
p6YfPyCOh9t328zhCdH8r/r7igr81shi+lyhEqYuuFTJyrMmb1icTCgqMytIWkjc
a52ucwXvtH2+IkJV7FX8MsAPJDS1jqgJ4OSFpmtwUioCJxakOjiNM5MurOTV0Yvp
NR6jHDjwTlES1UrLBBZZn0Y3Yz3PwZPx8VciJPHdCi2facp2iD3IHvqMPHYasfTy
BbMKvrnTaeZaaO03Qih2kdu0x1m95ibHVSZ7nMOAa2FQBlxMQbWaQ5nv1o4BNy+p
KMbuOP7lycUE9vuMxWAe4J4PULGZ/4+k/YjAyautIDqelvHhTjlySecj0GXmiMRJ
T91tpj8r1sMNK+6EgxuxdbTu8YcCLWUft+/H3pa5Tuat8cFv7GxF432YBkyUobZk
HjnjFW1TKd6NR3auOV3/hROJ5/cVplgI7XF7OIaiEB+g9/B5VkRGCqGtlcexB1ht
E+335jb5PZM3GlY3pRIK2YPjRbiYtdYdcW6rG5xdrRjcKkjPqSRXV/xMi01qJzk1
dEcn2NnVLGw4mom37Gj9ZKfl+MfRcQxTG9H9u0WAm/oKUtTtG5i4ABpGCWHiVPur
USitXYAavksPhrg+AeerlxQIA0Ywrl50ScS+UKBDo9HJGQjxbgbKQrXc5K3sKtbL
132MRH5tjE2f7tWOxDzk0w4Yxcx8nuNKirpU66f230XwgeNq5OTWuJPHaia8cZMv
xZ2RJwFrvJpEsxbo+sJQEXgEHmcEgkmF6GebO4nZ1u2DvL9RfqqBSZC4pNNuN4S4
Op4fz1RaNjpuaPSnXqat0hZ3qf4JG8LH8hoPuCSHCWUVoYfxAGnDhbOuNwyn7n5M
/LipIH5vqusVSTs8MHLET6HxSlxeimE908Tx0ZhkSzVQhWggRe5XSH4D95s5B/OC
mdmD5VK/4fz8hcqpLVH+7C7PEEqu3Fc4y+j9lTHbErg17RZR5UwQlpagx4GU3MxC
vn/XR54pNVZYYbCSR1jSfz529Ajg4FJOibLNvIpEJlv/JoRoocr6JnpDL3bIrSy2
i1MiaonmbVpwAheBZRwtKk51P+8+dcuikCRFtoHkfLopl62nyfeP7/pATyK9SSCR
CV401L6AhySwUfLMg4fAYYBv0fZyUY971BNpgcZUNsdB6fETgXGOZ3klevl5eSSw
7Umi0qTTc5xRz0lCzM3Q4YXg0QhvG8CW0apybVO/eTTxsPVlcAI3S6xK7AlA4oRY
IcWyrpl29vh4DBqETD2ApfEtfNTB3hI9VoZut3T44xViXl/PiqM2vRiuJpt3phG3
LE/CMZRfXTOp60Pnfrc5b1JNyRVeljzj8d0ax6f91NvxE0DunUf0X1qxnJIc25Yc
YQRyhLUp7XziXGFxKfTkHOWuAr/2xgeuPr5e52sIxMhjGAbQYcgCPzEYmdX643Nr
M+A8MzDsFEkkOxX1XY5ulGc69f5pIspxVrqSvrY2MpufiY/5UYl20r8oYXTz7Z/5
cgo8DB5+q3aaLoZ4+KhHHmcat8xDmQGeE4F+5Kigiurl06qfX7Gjie4KTGUVJFEI
4MD2VTiNtUksym8VmyZ9ZtmzjdGq+vZzINAqa8yX1DtLGxfEEoN1sQiL9QCfNyr6
iOyKc0MZJQ3TVxkpBK3NMZhs2hatUb2VeMUmPL9zPYmI12qhk7Ik6PmOs5Um029e
v8Cgrl0sc04WYcyWltpyCEpRdMEoMpsrxHkc49t1sHtdFPLu4QLxF3z1kH34RY5F
JxOokO+bCLN91nLfe/OFp0OpdCPy/Gtt2iYcIhhIkG3FEZ90xhTVJ/XeAuQcea8S
057JEs+lBxahU8+ziMdXspruCsLF0STcPHoNTrO1gIzbEiIabhzGX3ofqJ5Ma7FS
5osQhU3PI6MtRGJfq6lkwIqiNHIvbFFXqKnjGVau7wOSp5HwODPv+50iFPyUx9PR
NPv2jFS0Asi1Uf25lNpgzMSsSLPvqUpURDg/lr+pojzMwp6wdNo6aIociE2gClYt
KKhBTZ1002bGInrd6POgSMhOnuqb48gQkmNjqQOw2UUbAFBrhMFkbI1L+QN9jIl2
+3IdjDm0mQWFpbr6+dMkWS5TUAs9Atf6ImWfxDAUuOVoKXVzZr9RnW2+JJFdDmjJ
h4NHC8NbiYUjLWOiArzAuJZB5O3Gui+439DT/lrVhrqBGZDL/FjcAZ7n+Bc8vI4D
O4/QZNqwMp4HG365tE3UGA2t91TLEWBF6BzOmlbAA4MvrP3iaySUaVtqBnaoQmWr
V09BMVMJeBJxPTMpFt+AWYFY0rS2+ek/CF39sFF/DM+h/4udGN1Yh3HB7mjAQSD7
HS4fKElzibRnlvpOP/Lucy8CkI5mH5adtFwnqtXz30ZyEmqI9Rii70993vG2hDAC
fn+cnRzRD8e4gWMOuPGl8gTdZKb34zgFxOAAIrhkMF3y7in8Ab1g2SISYAuHXWKK
sOotWjbKQub+MjuWNKAvVlV+Z+HQ7wxzLC/VKg1PfZXbTdStHvYU3v1cbHB6lOne
bwnHBvH971gxwWTpO6ZICaMqF6Pq4wAaIE9GNnMBWBdFhrAd7Wfn0q8wISnG7D9A
bT8W2j2NgXq3GTJ+2SCfzWf9DPmrOHQW767IuCOD6BYK7AxyNOZRAPyvwNNLo64i
X4EsKYvlyHVK42OLeWTTHJAm55iI4pW2uwSpgHZPTsNxmHYID9qTldALWerhHoDl
ULJP6SBcOME9ds2ekZbzDVlZFHytjT1tQOVqEH4H2K/eUN9GMYbE9qK7D5xbZpah
pnCWsoyjbJrtedjqMUAXAdLODP28qz3eu5aHf5q5LWJgD8UkCqKFTWcQth/C4dkm
nKsX2SsIk8T8El0b+JmqYSND+syjw9QStMKGbtlVPpWHHAq6f9ms0zeRFIY7HP0s
w6UJV61+3mP+NA2h0pkQ5bPnErDwgq3cJ3MxKmT11ejrdPMvW7QXMmdu5whA+Ozl
YPkF+YZ3hDGwjlW77g+JrlAqTJfkK3l8FmqY3HoTuSRPFyu6/DqCo0mVLB6OuiQy
0B0a0dFruffDatxbEPE4sN4Q0E2F3DQ7YQJ+vYYZwWWionPGMsuBLrjbOrbrjm0w
wPsasIu4sZpc8JzhAysHwNhDA94rJgTqF/rZQ1aA5WAAQXRsuGU8Qxp35VNxxweL
t1r2XgErsJ5PcdgeDLjGe7Fvu1k02CPL0k8U+8QDyur1CDqt7OFaKM6dwaEnlNkW
f9fTQ7r0TukW2Pj/iLaF8XPBkv0jebOogptLbOjaDRUVDIyL6E34PBK5e5nsQmta
trrT7Yu5/mbpFIG1nyEG3e+rszlh43ZjG4J0uDrS+I5z34A6XZRzGVbF8SoYpX9b
cal6rqOsqrtwJTrsniH5jtmXUoBAhfZ5SOvrw4Z3HrKDXwpljTX1kGaCAEO9pYhQ
vs91g7FflhKp8AFPWvdLjpgDezBjpTMHVIkMwPzoIxnj0wjMfNyEQqzL6zYGf2My
xL2y1IZYGm+30Nxtbf7CI6MUF7O6POm50KuQN1DJAkGVpkMs2gtUpM0B4cJq0OsO
cYZtZumU2faqogZYEQbYxDJvmePBF7RNy862zf+cdPsfsy8mkS/ZvViu+4no8moT
8a++9GzkPgHwk68V+SgjyoAsoT0x2SyYwiyL5P5xU6nUa/E3P9gYBjQs6xgVsI/b
ZU7dOtnck6VTbyTfg4NT5BOgq1Y0xYpf0IO60wfP5u51L4x3rniVS4iDoeaONRkT
fyfI75aE763zU/eFkzdc3vmcdcB2Q8KCTom6ZB8kCNCcMMzsMOiTdD2DcyuOwXPb
3wlIir6sdEk78iovJOZgVOAelwl6rGFG78gudWNfEc1+MPN8RG8i59QFSbKtQJCH
lc5uFdLXLq0XrC7Tz/73aihe/ZnlZwJiQ/Lq/7u/5lrTX6Vsmhoa8eK0POwm/QOF
YQhw3AMNH2h/VJ0jHsufgtdBFqhYrjhoaF/AxuOGYzudr8qLTmwKc8de9ASmH8aJ
9SMNd3SUsbHgT4tz0mNd9z4KxX7YwqfZqLDCZSNX1+jRf13NRIpWTFnXycAAdWsF
SM1jfIIiNia0XW13aOuHrFZ5YvR3DMnP74+d9uQ4UH8txkIXWCiQONzV/wGCqCmt
z9AERhZNUOK6S8QskViMr2WHxMEKGoepNQWM06FrvHMLOhW/BVs7HA+e3PXqVpIf
AtQKT3YFbFp7tlQhjLin6Lt+7ZP1T8+i7ftdpmIDG1q9Rp42sBXithWK7uWy+fsA
xsCxEyKi4nAHmoBlXazwgl57vfWgRuK+YcGcmClfqMiL1Q+zG91LoHxYy7oBeLjl
UNRFb4+GkgQjmyowhjw1hi5hhE7ATobon+IlWmKYyKevLJtOBY7i5Up8RwsGobK4
c1jf46wNS2WdbXDqNWMcXbXVsgToMARNHliSG8nvCGxYnmi2mgtEe3l980Z1jtzP
lQULx8rgctWswZB51AhP7H1zwQxOtQqzx42IJQ9/He3hLo/Ncuc+Gd8fpcyCB43O
ta2YEfCa5SwpgUlKYkR15yRKO4YzEfpj7wOYDq3efn8Z0d+U+uehaN6QHm7AKSx3
7F3GhSTWY3TO0oaymO/Vv5HV9ds0HxIJOIGjxT4nXvxres9EEmsFcppMGSdfory4
daFP5k1tXBJudRwc3nifiqMjGgIS3VSUsDHtApY334MPMytM2F0J9J4Y1ujvR/Fb
P7+j+hN0nQCrTFjA2w8zm6yZut5tfwmt1OWyu7PfS4klMNW30iBwVC6O1IKM8wIb
sSozVpuHEoWZyfxwDz+KqdSO02M0v6gBNPSfYwGn/KbAzbtahpgLy5UhjZzhCBak
wpEBB8+eEWG1vzbu6aaecuiGDa/Ep+BTGArwJVgIeIUwzTvW149o9JwkQI9sSIEH
uLl1wHOzhAEpBfbiAiJnmuoFdloj4NT89yMqzjs8iMoELXYCqMVGmugUWl5Rp0BI
lC+3vTrJ3QBd4s9D5nFZtI73gQvdngziFZff/bb8WAr5xallNO8ndhCJJ9X/F8uC
z7dNWDBr5ZqCIpttMagFulyuWi9KtUisFtFr5yNU3NxIkPA1n6UHjSuIvZ6c864K
56NZcZscNCqcicToNR+P53HQA9oKmcx+623OqEos36HyncLqNGCCY66KdpW09KRM
bpW6ln2SchhESI/HPNCyMssTKSQJNQ6xc9/19UJ13r0KOdft7+78uXmDDktFtlTV
cMlzm1/DfCFOmImTlovi5G9DMAgd1Kr7Fka1mZjxfU6VUW2XZwaOyFLLMujcLpqc
VshHU1Z8qMAZRAi2achbgUaATsJyVFo+2FP7bw14O3fVDP97ZJGLd3vgpAoEfqZc
vjD9tl2f/odqZEfdJNm6YfRQyDuYEQ0+DLisISJqKKhrtC8fQ2l6Ve0f8/ssQoEs
Frb2nf2Xgf5miV+I4yuwWMPSpNwaxRa3+jmTqSmlQ28tz9rOuuF+Z2p0EzcYLQ6Q
xbvBBIkF2mmNy3qkL8p6gfI2fI8ULSAy+30Cw8TK+i+xZFy51H+oWT/pC65yuZAz
MjrG9r85AOgU8+cQKreRb/jzeH3DXcipUZuCb9FO3FXzph4qA/yyAWZXB8wdmBVO
QftgoSyqYY1X2vqBBpny4+ZBxcUzbcKIeNHc3AeSK1hoEDbKASWZZfjZqnnfzj8A
vXyd+xUyQkhBbDmc/JvUP3wNjIu8gwpn7vJyPSNLKbNNL1B6wYYILN/LbPtpIcFM
FRQDEvuUBdxrDSS0XHnv0Rwsudzw80t7jInhXvwUVHzI5XAwn8dwYyISwvQ9dRHi
lW51pc8PlDxcYg5BAr9vrYmyfGLgS2OaXe+23c934jwlfNWIv3V/KLHpNmB1BLga
/aOxcg/L1QoKs/rRLJroadMmQdjegE8IkxLoiKt5NnNY1QfxpM+d9Y0ifY7wdSdz
+9X0XQQoKYZoJZfdg2+b7shF/MBbfGTSPd7DYOiv18pJi1sHYjrFj7fvhd5IvpXL
pu3vLa0BteS2iQFngX7p/gi4f0TS3oA0DbqyF8zzpeTF57Y6AkmRBTPWQCbyprW4
D2HF/ecuzbdHOP63bcO2q7WHDdwxZXMLPV6bnnsZqvndN20jJAASzxPotiJ3P+U9
kiU205S4UVqzEcA5nt828WYd2PVhwrf2lzV9ZeYBm9EoS/LG9o7LIFGWWsnUOvDb
xXk2iPZgpV7gBqkxd0RPpdSgSS7vnOpfzfyEdFTHJbwycz6V1dMjDl4Dv51d3xTU
cu2/JExi0cHCAX/7bc8AflEeCI96QnfF086hiO/7QA/YivfxiSSKCIj/IvH5NpoD
v30K/F8dkMlZ34bG9QCI4uSQSp86/gS330NGecTk6Dc/ysdO3gQ4TGpzazHkED/s
1tjvS7zI6jAI8oJS3W00HSbV0GC/f42CNBBYiFJlBQ2r4PuRiaoLOhA8vJbq1//r
30CHUPcpvoWUxF2Pcibwwb16NGw2oBwrM6V4cvHMfaN6QVUnPhSfl/jC06X0NURv
cgRDbea/R+d28p6awobzm/hAAAE49YqoPMRdHIdYXpWEmcCuMH4hv+jFbQtVWW3F
d3lUFoc9Xh8etNV6x4hKyiDp1IEp74oj6W8xga6+ee1EC6lj2NA00vGMnm366aqt
5h0v24YIi9ImVNmyaVJJms9IpBVrle5nhG3TigVGSbRVEn5qElVoohbruKGLhA5v
zPsWFzM5CYFW+KAQDvnVXsDfcM753GERlpQ7JGzsS8l2x+eV5Uk4CH6GlZwz3GCq
+HZV8jUAHiQ2IcYF5VyH9jq+ZpOkMPBhOPeyIE+BYtPUD2K0JwgxmDtk35fssmZi
8U/R6Om0kTO19pvrGbmMjdfTsPgIdSChLBA1bHVJfAim0/Z6ZXYeB6J9PuyDtd4E
5jdHdnsgYr/5/2Yk4rZw1MUAtiPZ+SAvBqHU3kZxQBnOzvq0YvqWpH/9PVaZWmKs
jwFemIZtYCwdqN2fd1lmYfirzikXxugsWuDqEr4HIZw2OCKGoYwMSrvaqxSIP1Zz
cclpNS0Y4PQrNJVgzNdZdC0QmLlJ48CUFPSRSfVOXpi4BCWM5Gv9gikmKmKC17Hp
zex08maFrJi/HbuqgZdF9B+LOGXwCHPIpyadwgQnGw7pEM+1JTbgufwY0jKMhFTL
BSCY3aHwqLvTvmFtCBApFYeih4GETZmvxzPAdHfv1JpfECrn2WDnPhUkQgGx8yyx
efQeVaBfGALdEh9H03XfcOqjJRRp1tE+k+QS4IscS30JrlmZMNv9EAYNyCVyEv1f
ALt+0aXvcSx2pgOipZzaKQxQgMHlZd2tJTNBnRYlFLmXitfra9IPgmJd/Pc7c5fw
EdLU3LQv+RmdolC6SKVoKuQCfkevfRxjefuL4tmG5J0ATmpzP/QXQTmCSYoH5lRw
9e1y9Z+6YHbRpZpCdrTnDCrLt54eyP4LyPziNyWhxUhs9MQp3dmkiWGH5D1/hU8Y
rybi1VwGL5MUNcoHbPYkjj2DyhGh9KF2m+VQtoARfA5lnE3tqbmKhdZ1mtSai4sB
gorkMeCN3B2xQrJJtG6lNrucFlSPZ6r78yfZNZNklr9EQDsf6KrVmEortSai0hO9
P3tsR8LBSu4BVRQFKms+kaWQBfrWLnaKdvkZF9F1mZZq2E4nSZIA0FeSmJUa7fAE
x/WSROK0h6GIIAhi/1G4Dhxr4VHonOzpZ/ee4tT8njjfAVqdSYx13G7Qne3PThzI
E76FAY641FUL+SyQ3TQF7pk/RlFPr3Bwnl6l9OOSUuBw39+oVGDmS16daFx5EK0T
jKVGQd/72zDCEk4fWxsbeEeERvQdOlOjdQli72laC2p+ZSU1uH+8xP08AA7Gdk+A
7H8k/3tOLV5SPGbZu3YSsme3VeqRNwtGkhf3hTyHHRmT2BgKYh01nNcuJ9yA4o4d
rSbK1TeSgj8WnkG4roEN3NgUxmiHK+OY65cQKY+0jqxC6ybFD1meCjOH0hEx2mjp
JZc+9IdAlj/o4NGHZjZUlc07v6XW9YmYgJnD2gKfqcp87f+K8p7M8lmapuzVcvz0
wothJ2Jgha2fHwg/94rec8h54+K2mihnkauZZWs5wR7QC/cza9EheYPhWXrM4gty
MKJLHesmCwKb1l1kzVdVLj+FmooZcsAKfzOTRIIB5QNLd4OfUkaCljzb5ZCuIpsI
9ty70ljsBKRNCWr6wndryQovyTSahIR3KVFEKSati4UqRvvFnPTF4bdUZt3lgNxe
I/WYoQ4SIGho1fgLG7m9bDT1jlWKtsyD8MlCnCXagbXyxf95uFO1qqq8OxWd9X2Q
Ln3uUJIHM6daYwFEsx+SPe13q5+EWcrODmkSLbgU++W1JZFE9vKXp2PjtEJadLKb
5s9K4EjDUXJDZNUfdbMmW7+ymbwh3PpImDJthQ5ySqsBhA7KOqMzLrmybxr/MLdr
mq11cGjP6+7bKXaJtypuXBTcBG9njRQBDmwo+pM+IKrkguZHhX6plLOdngPalclo
kEt25dmKK/gp9hVs+iPWpY0OXpcz4pIxMwX0CDKrsximQKXxDlbye0cWDOJ4xFuR
eJ7E+syM2S+rkqytwWEwIhemcjX5FMazDbxrkeK3b9FtzR/iHsptr2R+FOXw6XNU
Q6zJTzQ2U/zmv9Ma9ZihiL0xWQZpWN2E4qTe5ofGOMb34bMWwY9YjCnIvY4G7Jld
xAp6EmQ8CxQ06Ova3ImIDrP2JnAAegYGIt5OrnefPEB57KeL2ZFYtPrK0yVOPCIy
4cMkXevR0XJewTP/uxVqeFq/HoiyH4ez7nXVYMeX/z3VnnAs5+XcI2XgVNzFS4ji
RkZYBzV0XwihWoUkS1hiZzN0NJXjGlo2Jhp0ODUvHnsMhRQtxuLeCvPcAC9JFMDh
+n743ZsMcBLfbzlWzcB4Kk7JjgjEW0PP1yUy4qoGRo9Q/6J74jAOP/I4kPJ/lP0M
pOkSokVLfOfFZxaMMEk1Th0JDgUrP1fT2wY2V++a2wZKfUN7EprZkyeyS3hkC+KN
6q2CV/EaCEtSwdbJCKAIsH37481HBxxexAmzdOcxugz2B2OlyFl7RFPDBjplAOEk
xX61WUan9NBonT3DuLVc3yM9guiRoNEm1BJ5MkigxXzeM+VaAPtPro+R+YrmLoOk
ID3dyUaSZgSvvGEwrkaMPj4ePGsroN34Ufs7XlxT8NZx4yCY/gM1kMS8eY0C5XoS
JtdNwL0JK3ZPYGkRhywVriJRMh0kgwCiKJWEyeZehXV9sF7tXD+oNQkKyuxev2Cz
K89K9OHd1DiKitDKYJ0QUB/m0QT1/CRKjMrQAGajpTj6kKS3mWSVIq54bpDsl2gY
766Gn9kzVkZZkY+aK3lgMU0/tPtDMbZzHALSzLgUEK0QuPyg+BZBR4DJ266zvv8r
Vo+ln5LU0DyuGGpqKvq6X6m631BVRL42bPMA5T1qhb1ee0x0Hz5fzNgTYw3ErATB
B+J1UeEqLSWf5pPBt+tggnIwTb9tv1v/b1urJChzaz6Rrrjs6zqZlU9S2ZfrdgdC
RVQVpmbkEHUuoKM95jMUfq/m+IYv3my0Db/OoYT08SjZV8UQYtPVje2vCHFf/F9v
jv0Czl5x5/WUvfPPJ+RSWY5Sm2lhvDoPU10xD4/w4R4mIGE/cEaRqWf5ZTomkk5W
57zPb6jRClzzPHmJwHLAGgnmfjhfDUTenkdm/6mS8t7jPaLM0JYrlg9X/ZsEKkIh
uSSMGd7jw3t9bZEvASnn3yvQ6l89gb5uIE7D/NTtQiY+9hpmke7Fb2O4MhK2V0rj
c2bUNvb8hbshOEl7piSsFtOwjh48W4PS9vEcVCc0LjvZhgmsJNKLVSiCpu81if9G
X97qUSrzIYsakTLVvOY0v3VLeDrHTwBnCWiIjwuA/JmlSzke1jI+GPsMrLUfWrSr
uw7R4kohCeiOhev0VU7dU5LjIAHy8a6uedtBAjx81VZ6Hxa/gm/ZD4cuQ/EA4hCO
6YySD8wQVzpXGgesgyg8OrB90Qc07OUqiEUM9LvxaF0ZvSp0wPck1MLXDSPR5ul7
gciduKlln7UsHTf6m90GriOa32nnPC/89h+7cJii2F/yNitOuq1NH2lQDpDcAw4F
7idwdQvdvyJkOliHMHvA8JNyw8xuRy10eRXkHXmN+rsyUYVKd8A79EKP3AygnSWR
W//Z2t+37DyhZ+OARz+0ELkLIzuHF5pC5E6qnK03LZAWPS60hpv0hvDCllVIWLR2
JQjFUsyRlTv7RbKpcsKAY8qd0f4sTukMrhaXJI+/9xT5gu7XPbT+FdZc53wMXNSy
vn100zxJY9C/16bPp3XiqcLSmFUwPuyHz8ZCjz6rZaHYJ5207t1R6yXF81q8MwF+
i6z+lBuyui3+D8C0Apo1v8bKk1p8NrSJGsc2MbyYOqXmpaQ/mtLG7A4XJWYRuX3Q
ykOKW8E9rAHEB+iotLb/8VIB+HxlyAPzCJYRRipI8JkqbUv3JdkY4aOjlh0ehq4B
0I/+JAmCEkGx3nT6z05Vj4G2u57sCngqSw6btr6Fa37ktYiyhJhi8juxqBVbyX/x
eqllEQVxL8ZpAGnh3nB2zItgFRy6bvB8pfWnZ2iYsWLKk2It1v+fIYPBEQRjmnzD
hEWgxi0+rvMTMtat0MMBa3zCRKvNgurExwQgoMj9Af/YUuGEFcM8LLxlhrKbd4rZ
OPL4YkSuhF1visKcRFoLtRUfS8SIS7OIXKyPiowXVDZQWvd+OkE+HYqscnleVy+d
qhyXwgk/rtucs3DHPC/dI7Qa8L1+4pKpYw8bWLuCn77Ge2AfmKEpzpzfuPQ0tQIz
knUdddKxN8kFp8hwn+2w7TymnTGZTQMd3bcIGq/oLZBsuydx7VkqHb/gCLkgbfpt
zwiOD5vFhSZLdCeMurKXvPnEAcHbXruNk99AqO0zuVwJ4roPluSrY7T2RPIj7mtm
Sjsql/uANqETBPK39Um5BWGJxWHepSPuY8gbNkhUnWYC/uhAQDUG79px7zLjb69T
RKWk12RQj0UBGcjYJrvUNROqoyba51Q+QVV2c+KhFwomz4f21ARKZKL0i9j8ePV5
YQhChijJ2UlHZq3qVaUeW0bCy8VmlRVd9SjJOzaNfhPrISBhKyP/0GvTCFwNoGiC
cJYsLvo1RokL37aDvxkfWl30LdX7vGdHtDP1RHuVmMKJvOHo6JOpu2Tl/vWcGHcF
/msJ+l4WnYyJyrJbFnai8YxB7cGzmJTj9C0iQXIn3Z+cs2+NEeebdwby6tig1V54
JBvk5XPy9XjrqyTzwxZ/QRr6t26DcALF+GWuSA6KK5zQhV1bfIZHNSsXynRHgZ+D
6PNPetOOjU0lOJhesx3jaeA9HMyVe9kPN8ofQFmHQ+/nTKt64If0B/7str9hfpJn
dK63hFFteDD4NruGoG9Vqzelt9B+wuCFs8NLzK5X4r9wskA5JPSRJg7p/TDRdFG/
kJu1Q26WpimP2dP3UWwl8knZwgfNmHcmh2PYoTePAOv/yLuaHWqF5X5/xHBMRLCC
EGD3y53f1f04+sbV7h/woQUFwtDwjoY2kxqoUw9ujewdyidF0qSS+eHVrps+hFhm
Zyv/Baui3+Jry6tDq9ZfBImZMvFDq0dvK48HE1IQkJG4vaVa0JisDJewUB/VeSRQ
sP8E5OEMwtmmOD+8CJUzJQKpZ5NzXack5jsLiN44suzcx2Roxke3Ws374iPyrbBp
aeQE8DHwoCp9QxtsusHUS776NTTEE8AXajP+1xgmvGbAYAOxHBilj+NhIne2IZ2w
KncXJlGX8I5qXCafxN/dxUD7a+c6BszbnZHhjAb6q3pS6TThNyRVs5VMAVuwtbfZ
8yHuHryxk1a6leay/EnL1O9cZCH7aa5g3Xu6FHN7gbh0CmmRvP6vXSDEAmVlegbq
xTwvdOQDbYKZJFwkwIk/p5WNHa8G0WxI0tNuKc4AJE09v/cGcbVwe/ZQA1YPVLRO
t+vpUAeILKudPyJn/xMKbIAkIQKpl8SQ7h9QEMdKflHjHi6PWpE6cw9k9o4M/hly
lI8yAle/3QCJzSF+boSaS4hqRwBC4mWadIjglnlpUs+gjSiq/D2qo2r091RO1HFT
03nnudgnEClg/ILM6XgERDquFi1CT30sTGUiQMNg7ZHrFmrr3i1Az3EJFlQLV267
ut8gx4CNH467RJ7odqWDtXXtUW0WGyd6ABA9OFUyiOH9W8pbOfSE1KTM54Cqz6i/
D8X+tqF7ZWOt629KMvnNVLo+5lpevKp0D3Y9Hx6mVkHU+wyihWng2jUkHSm87uXa
Ljw9jqN5+vo3xl71hHwDWPTLjA4MMOlZyJA3qQVSDe7/r6OspsjygUl7ccuo2uQ+
GD55tdw2V5HNGRyAekzAEE0JDips9yHQ5E/9ooJPqyuqu6gsQDHD0fvPdHhGzIhp
G9muGXnuQu/mFH8mzSE6eVYFZzwjGGXS7zOPWArwD1YCam8/EMFd9MCDEqhBkodx
aZumPOuCYieD/+M29TI0k8k21XluBJhkOmwb/NZKajwNZHVhrIP3GAlrwbw4ofFF
/R3U/MrLXtnPMQFplx1En8AAe3T/ry+J5ksqwDSY8loc+7MovupS7rVvkd1kTJ2Q
aFadMUUgUfz0Uie56XHqg9tnFmAwU3ZfD3e1Yny2uWYNwhf0DA5qTWgGS+VfTsmL
SVOHDjuGQlwdHytdg7c5n1dICL7OI98H3ECaYAx0Qrlhk1ktiwerNleY63n1WqvV
PWbzeBh0W6PImTChyn44yf0JgiVbmLqxo1z5a4uofgF+ouNNlI1EX3kVM4SAd7gt
QnEgcK/+8apHBeOxleV0d2ffXfNZnWARIg0nKyL2pytmNw8ax3dBCnxlYSnbiNpE
SzdyULSVF0b5TPAr6yuFFsAz7S0eU/+/WshQ2y8ifZdi1brpGOGatt5GQ9UnIIFR
+xOm4ox9OQQdOPlz91/wx1MPtGEB1DVPaUBc4SAI4OSV4sCvSiHbdeixHdF5darx
qLJSGZDGE6aFnmM/XXuvmuXEmKeNdUJtAGCeKJAAXdIZ28weicZJnmzrRuRD04um
sSAhoumUCpiJDY+CkuSgZDCoJeonKBm2hTn62PZ6Q0vD7ijY7yewi47XW8ywB77g
w6cwx6YOI5eDF7EOUQ/Dj4OTEE6uLAgOMY6IrJu5ylWQlhjh3QSmnmiCg1igaWGU
UhtL67LL7DxWveV/Q6z42hs1SBHxdCkZk7DmbEPw0lJdQXp+l6Q2j4WkT9VHrMFl
bbY7yzXbCWYC14CV9f2+XfIkfMcDvoLgtQq2Vw6j6MVVHQQ4WpMFxe6u8ejioDrC
D4OrqD4J3cyukN0dHU3ojHI+r+O7krWi44GrsmGJiMis8VakJ3CBEqcLpm1lbARb
X4NoUoAd09L9ZaDKt6/HmCBcEDeVvIlSqJTZBnZOymfsI0oJAbnpaWy1KJvk8ml1
kPVDMaYp1Ae17wlPCF/8BXnhKVDXueScSeittYIBan/Ko/7gpvCwRo9MYXyULsCE
+ifA1trGlxhKHceuueIj44fzDv5wa0AXLRx113QwFLwxRX0q+b9ufPon4CPwRkEk
Kms/KYX1wJukYhiSmM4UVGVV0t2USt2wMc0slwjEyxP9zu9uEY6IFVBYbtr7ZWsI
JMGt0DJySckObCpbxfoykM/q51G+UrhJcfdJRU5dnkR9YMAH1C7l+hWJCCWfF65G
tamYfmWcEq2rsW32pVK7pHUvcwBB0WCs9GOvCNfjlQNKDg0L4ZPP+N4G1X2zkK5h
4vRmWZEEuRRn1u7vwO8FmtzELOCE7RJJM8Ymc46oHkcjKr8qxHh3s4pHGoMN0/Vn
B99zBuqxgrDgJqUmoMQ6R8SQzoWgxgRm5bdNfW2rzg5txDfIHLzNqo1Q9VvsSI78
VdNfEoNxJkx69vpCtRuuo8hQpBrps8eUtE68qO7Dg6JNtP8bmYCV8Hx5QJdqSUXz
Idxe/h762N8azLqsc9oFBxQr6nSf4ZxF0qSpXs1+SGwG7cP75BnBK/sPwF3xG0G/
mo00yMyWdP8k9hfYfI/R3L/kINIAwRkycVkziFyz72j5ItcGA5eSq0WKuq/G8TnZ
YJS8YpqcDPbAjfArv6ADF4yD/lKNLzXquR7ZIXhKfmsQxNhl3Zr+KoHd4ei7Ktcm
H6hBEY740LF4IpMePNf7A+RkbMhtIfg3gxe0j3d3Ee6DWg+FQg4p4MA2wXx6zlFj
6I+xXukn6AR5WgCqyFTzHChTpG2kIvR2vZ/+QUh62EC73TTZB34IqGNF75leXdoz
dOOFpTKlA2H0FWJVaQOnls+OXcmp5sau/Ksb+voDA5Vw7hrOIZvxRJZqGSpKhXG8
OAcOYYNhu3ArzbOqaN5xuHo819zrdyYrsR7FYiKwBN8evwkBYhHgoLAAQt25J75i
vrn79TTIYzPzoJW/Vg0hPtGHP2P92qQ/Y5O4f9BV7rupPEkzRhtPw8Bc0BZuIgEB
4EVszuNKMzR/vjIvcKHyYoTEtPskj5WTaj2inGEh/Ah2JCwxyBqRNc9WAx1FqHT4
kFv9rBgNrnocxz2MF2EqVunr9cufr7AJEWdqlj9VpdymHErC+QvlE7qJxvC9GjAY
Ft3FErs9rowqdlH1mpXEd0C6KTJUDqpCLFDusrU3LJuSoy7KZoAtJh2FVmdDuyed
Scs/B7pG1PGjCNFepqRAYMseIZkQWNRhrC2VZT9Lp1gFS82xjTx8DixOKCqyfhe0
MrniFrzbXJ1zRxYXlNHxwwkS9T1mgO0ApoAqEKS3l8HMaavYnkj7fBrnE4pyQbL5
DWSF6aWgKfYKtNIhaLSvvPb4xbxK3ovdhCYrg70o9LBqeczXQ7RCxnoQKfFY9OKq
Uxt5+ZdcdWyMHZTEBIRK8UMr6lAGs+As+zBI1xQsDkNlXwbeGPYDqG1tCyEfd7CD
4WCtYbdKntN0EAXwLuZLHiwMYAlEyYW8y6pi99d5LlVK0eYYcUk9/4FMRKzhWUll
jhzP2NhMk6MPpv2xm2xj/xZg2BpZVlXcksCbpr4t9FLJzzQ/cWyG9mFsYX5ZTuAJ
XhUVZAj9Y+SZVS/1kWI1Vicf217632bJdN4n8XOwXAKQ4Vww0UlKlKE6yN84NUZP
S8E7vI//cpoVisTYQ1dhZh1Kc97BG1KZE8SlTIr9J2Cta2wVMsZnEKhprRfgoTre
fNOoD5Emon/UHIKlNJK7GfubnqpepOfrIg8FKbX2Qp7VTMKu9z9jxlWvXVzqGBa8
HX+ChdGhkseZrMA2ayMWXMDxkZMi+QdoxHTOWNMgHgWTknmUVJFiPdTpdj33l0KO
/Lz9F8BjjaYhbwUkMuFwNNwt+sagl4ND5thItegvwfZ2rvHsSIJTRwVQBVgL0eqx
wE7rVbjsKWnnfsvuhJ4HbFvYnn+y5Ph66kg9z+FykO2+z0oJOghfYST3MofQajp6
hcMlxIvBP/TCfX7qnzsKunsYR84l69jG9h0meoJGkrhSBN7d7I7FB1CZ25ynB74y
FUGwdeCT45+wV8EsOZfHsOD4uQYlwH7mnOIfUf1kJQmlRi/LRhOsZkyH2vY5IzLs
+wGfjnDSjIG/AWDd1recgG9nsHR3DZyx3SGkGcxWplZxI3MaH42Ynh2ChF2bZFRP
BakZZuJWcXW6eARTveRIzBJBMBFEKyq6a4EEGl7pPYSQfptyL/SEvZ1EwVYGxcXS
i4tW+nQ0/oBIz1PiGpdTyQ2x3epXTfIBYrvHCcSwmOucCX/uey9qHwtoBGK1yJHF
5cqMLTKuPSmcY7uYv+3AVQ31lN0oFssxZDgDX69pyWiPQ0MN1d0qMQ2/gRmOgLpA
NLZgWj4maN23gY08+5oW5d/LTHmGGA/HNX5dOOFRxrbZtt92D+Ki3hwgUx3ORpWc
5bdGZBDnI28kYjGQsJbfUqllSBvO8BbLh1S0Zq+MuEIZR7CBLRy4XjaJFsVvK5ul
bIPgoqXFrrNqEUaDZqIiNzr4vgpRAuEwJcroOT44w1IOvR01aW+mLwlJMVrKKwMz
uRupr41wNLREWeYKE3nQZ5gzHhNecD7gQmL8F1MvumpWhiKXVjj+JPfXhaSKKcI4
7QIC/aOKZ+KGBQFxzA/a+iKLYjP0xW90yA7vVEyHGlw9Otl/RyEJxQo3S5/8Nr2A
L31tQhQ+BuOde+LwzEziK65mqWwgs8sHabGH5L+/lXK2V8lO8MTcom2fa27on3db
k4WZ2Ykz/Ujjx6uQRBQbwEjJS9IlEm1WGiMhqRDEh0nZTyoo20l5uDjm7vBbfNgt
L7Jhlv83fjfs/tp5xp3382cI2kP/xkuZel/75j/bWs7QO9i1xSxjcNWnzhjeXsOF
mchxcqxZzoSqekv2gSxVK2pbshYgkqBx6uAfSy4nW8GlNr0F+5XhDGPpj/vScXsk
xYbgYVGf0p22CFCS0MkXBLg3jd8wJBHTe2OyE9G4SFKbgNZqYrLtRb7h07TWC5QN
t68xwnxkuNWbBkYUe2lMOB42FI4F8vaVIiRGScl/EPt+R6gxrvsboEsbQIb4eppp
CVBHmZmkZNMDyfYjARMmGuMrDhZWa6pAKtrK4TEoFxvQNE3/tZAnGu2OVFS3xlXv
xlScMpG8zGf3OtViS6eyMHZChwz3EZP0PloK2sT8AkUvsMU2aMegoQQ39Wfbpn9J
C7ltyJ8+7O4q7hnyRs6O4iGUlE1IDVjYh85QdrDG47BjAcpLuvNSsLoiowmBAivN
LftrEiCsFN6Qxvkysmg9ChJfW+ThdYkPCDPhi2l6QoJTRuiZL6L9qQxZiCVV+NGW
ahf8VoudR9X+1yDX77AQK9F9LL76TYxxhRa0OCobQcTPNGYGQ2Q/tO4PnKVJbXL6
645EWoVsiE8HYxV3gZ/LpROBb7yhL55Hp2RU/9+MM8iTdjBzvuHBA/1U2UKAKFMg
UyROhiBnO6K1WsqJ1eEpqkBMOFxusw/pryCEAuoitM8mgg2YZStV2lokiGgrrYcc
9Z5Q+2fYEe3LW6m2mawn+oYM8OLmO+5FRhwf8IcLR2kbnF6J0M9JjvaoHo5ib8wz
C9eBeorqjv1SeM+5kt0Q+9mfdJst+j2VlTR/qfpXhZQ7rNQma1kT572yvAHuRbtq
Cx5AGMOgaKdDdU9xqXr5Lt3AVREmrM9sm2mM9JKJurhPJ8KIoNsSXStRO5aJJF1k
yylXXwg3B0LRydQ9bgfL0HuSF1QaKCi3+yhwGCoh1hIFb7j9DhW7nqiDuqXIscK9
zu6B8FDZJgMvUvzN54ce0jyHXRgtFgfHEEruorkv+W41IT4PaBf5o93DPtf4bzkC
UEJVeNAJ1/ACT0S6FhndryXBonapz896WJD3T4B4IUEKdDKCAf+YqhqpWE9for9O
Sh5WLLxGX20KG3Y+mTC/1HotxylD/QiwOEKq9lWeo5Zm+ToeH3klsZIfp/mUzkqw
GniGiuNOfRE+fMDgIYho7T/RSmqK64qX4DwO4ObplrjxB9K7HsIEqfPGuHRkXmDK
XNOrdC7H6e1jCvPZFvypxmT43tSk4IQz6MBjVTzGxeLIh64jJ7RSQzwiQDOB2dsf
Qopji/bAW26cNL4jX1/3w5tRsHD8o8sP11eGheufyKPCkWq1rKkza4JiuJCwYsTF
QnbUqJmr1GqTvRADV3Z6sjoCLiG8ZY3uQVViAgMhFUKZ+dOckFMBc1SbPzMdwXVj
0HBuvGAsxnVZqpbCX6YSGxONylgzTQ642wmaADouGZvQ96H1+7lhMt0BeaW41EnU
2OQ8UdUzvagLdEbSPoygZhnvXjlsfiNl0PY2Oxm6USjMpfRDeHKATewj3Q8kkNFv
7clAFXxXNDJZvwEqgfn4+D08CQlFp5TlutvYHM/cnnpZklGzyc9QOTAQH6pV9mX5
C2LhreWDbB9CHYF7UWXOzKlw8oF0Xnk0JeULNrvWXWHm7H/fFQFeakv31+kJe9a5
THhq99aik2xX8emkLMD5HpE7ONRngo/kxT7YcAyNXxpgE55LNKHKtiSS3zvij49e
U4DrKFdeZYnCtJguYwR4x2WEjXEwbOKrwAY8vMtqt4sWhNC9FoDbVxQCc9W+l2++
t6fBQjjukswQ66YIwAWdZGBdpohNGU86dUHk44ocCQud2mHELjuzVxUGVfx1dN/9
1Ra13kGc3ebuhbwZlvP7EDpd0+Q/IoEVbvWsnGKwU7MPFHd9LEHTGhbUYoUxRKVN
9DdgyU/viNLxxNgdMCNcqKoimgi/J4vc6rNU5F1lqCTEo73xvseEUDyULz982HTQ
D4qntrotgN+Ajexi6aT8JAUGMlCnirPok67B/WfRd3TbYDzkU2gwxJpCBbdjSJmL
CCYdZWisgvrotrOTbD7LITq4DTfCRFHFlvzqqAorT1s4rSo2eDItbrRn1ifWUh64
Ie/A002ddR432EtYVLbKGLMvBzk8SCm+TZsuCQeZa4qaPts1xWxnhsLDv/yGuLWw
FxLkqBtPmp4uDM+fr/uDh8bQkis6CTCqcb+dl4Nnxy+hGmjZbvDs8lPBCSsA+P2r
P6sEbaQdY6axgzn5j917EKaduU7Ig3vMqSIm8HpFLvHmlLAFE70tnBWW2mj4Wljw
J8klaDREGYAUOKRGLjRNG6tCoUJtLxuQ7Xmhkw3uoAU86zZ4/WuW9qVwa4FhgmzP
S0z5Db+jL9H/ZpHfKb1EGNWMvGeGGAE0VNdXWZz37Z6fJuXW+xaDUJ4hC/R1P759
p+drHlmzcq5z4V3vbvDvwQzsW+h3t8lCwHuTiRYqqLigdMkONSFWycdFAuYTR0p5
9GC6kG+eLNR/GNDQLZe/pZ0XaUd5Umd2uiwPehC0tcrlXb0jetdt03oahSoRhanX
EY944f3knKS0sDBeGSKKAhaGB9UqMSOf33R81GU74+8mtEQgLEnbnDJ1Lgo6bKp/
nqx717LtUD4iNTbcFqsmZSdfvPQMCD4J6enBUW8X7lQS42v2UznDgpex5P2ysQXe
g0w34ressj3KD7SK8M0X3COXH3wLmd2VpqUzHJk6r2gpCQbJBOCK7iHCKmpUdbwC
JRO2QHKfrv8XQmSVzrSfJ/CR5xIpMuAousbZzq/LvghBeC7R0wje6FUnpOucZD7Y
xltPzI1/nQOdSyH3xQfsiRMCAjHok/f8W700M6lQpL93kao8JvhiKRyZGtIDCC6y
3GAFaB5q5kjSkRIg6SMa8OXKWZ48RyWmbMgdsVAG0oTBsDBlg1NJhLHLLP2IH9pl
XGEseexWe17AjIV8L/Zjf6s6S93/NoXqmqfOOfoHZlcZwq7l8QBmEnBqTCnNxHpB
glRBLAV4s/ZIHATGceJbp2ZxJkB0h/legf4m3VGXHbgaz6tVvSbPMb5QJCKvqQ0h
2H475iyT4uZJuecLvlmhsAPpAoLMutITIKhY6vQuTBRgPKu/kLYOC8Oy0vtC52kk
ofPfBgFQNuA5e2tQdPYqYsglJyErNeTNHADUCHuZaqi0W3fGljWfYFdNjjhU9CuL
mLrLRAvBh0FT0JWnSFlTadd3BLhn3h5y1wP+EiH9AgkKH1mBO7qnyQ6mrRncAgTe
XaRllzcJo07S7RseNek46GAlfcB2IFbFy1Tba7ISHf0xDuzEkLtGRPyjEiaNQCVS
rtZVHRTUzXp8AC8Hq8c5vWH2oWfyS2jJIo7KGbpZ5qMKdypDSt9z1A0qDiw2vD9e
oJBijqP3MDvH3bgSiNWYf4i4TKKZJpa+OKg3lvMd6KRHOf0GaC/xQNQVPUE2kMOK
3YcUOTKJGyhGlW6kuXSTFcGsw+sfLwaIRoHE0UzSXXnFNhzcmelPr+HR6WGGz4vS
8xUhcoOja9GlfVhj2KkGW61J3UWe8uHuLl5F0aXDwvSVZgqwyhOexNHqfNbLs57n
EA8kpVxyy3k3Adv5A0JRucU1MjX63cSTEaQHGqfPmTgbsDtDsVvvZLiw3XoMZLUs
irG9tCRK88SzSTNPAwf+dij23KkyBlxqjh5IlwdLlrnOjlTvIVYB4mDQHN1x0K/K
+7ogf3PBSTN2U8iP4kk0H+Z18k9dZb47bt2ot31FV7HzgCllhUpO9HQJgKPfvEju
YJtbaxYK6d5IdkLiej4mNqbqDOlUukI0DMmIl1tBy0PCXxV2EPVwPrKumse63Yy6
ySyAQ1mMM2/nO/pUcHS7rVpDFMlF4gCX6wK5VO/+v7GAruOTwDCf1aEq9viPlaAH
r0Dpb0HtKGMnnVMRJjok4Nw/VDB8WpPtcPH2BAWB0PAZeKqrY48u1CSNve0ES25q
OzKmSPNqymqHJNoNBeFeFpVS4bpT7KAkiQPpO/4q0MlE2OZdfhjXUJWrm7Rcvs1X
q6FmTccVKe51BJiKcF5cDfJXFdvjWIffhHT8V6zGJADyn7geUKiA9iJjaWQJgzNi
BzYVHkc931qh8ynJ4kzIMmdBFtsYlaJatWCh6jFVwWiV4Mh/rmn6sYlDPje1rzHw
x3JYvig1ZPepMkNe3/hxiLA2YlZC5Q/x1I2u7/sPZeA8Zwv/pWNWyA4/XuZ8aT2v
10RQdynBhQ5mwMJhoxdlA/cogm5C3p89BiIDTwV0QYp3REVhZQmjKqfF5boh3TB8
9M/dGK/VpuzW6s8AvrfdKruJRW3KVEakYVoZzBuYETcyUXftmHkcVV6lIydgZOoa
OgydHKT2YMRKwR/pluSMUyY+MfY9awR88lzeLVceQ1HW/DZbduWaT++MM7HlXkpf
NtMsnnPkx6AiE/0s5NvetmOl7iPQWeWtelppCiXdj4aAIcxll37AJn5Ed7Fe4V0L
EYo3nDmVDhaaFQLpTLbcRTGglZZL7jmrUw7r3ISwr8iTXOyjXJ1x4tf2ddQBxyQf
RuphxNEvkNNEx28C87qXIzCiWfqWXqWcQAXa4tDC/v76OvJit9yth3MErYUyAFcH
Rvd/gr/3MOBXyOJVPukcTl0Pzpzb9WYtzWABhkNjubVqbDEfS2xFjmI7zLfgMqKA
CP9vl9pM2UQHS3XHuP4lPhafVqjbkBxTKbE82LdFZhV9WCkaydSXW7IPfdtApurO
B6YjQl2vufJbHp4NE8bJZmQbeevwj4cI0pXzHsh9ccH2O5zGkr+3sLQMw8/VWcrt
FE/RKAOXuWColBIHUPFF/RNf8+vDAS0F/2UAw15P9xY3WKc+iU9mSghFaj0yZd03
z+q1J1tVj9ODacaj43lp0dO/dPgvDimpS9q/1sry++3/FMEUNHL8PS0a+0L4ejQI
NbDgCcaPqFUx40j9+bboZb/1a6tG7Mb4viRsewErefryfiS3rL+n6IXzqiPIr/WQ
4Dqe3BqXc2HYkYXJ3yn51QncPnSePpanDjdE+O0F6rZ5Go9JIel2+C3zpbntywtb
pfgLbJLelsI7+qa44LchHHe/sX9qZ/JzDTocllOFQG7iJHhmc43uWIeKwC0JfiKn
abq9vHhmo3B1ggqie8nyPBipP/3bvW9wozZ4AVPmIgy1xc0VpZElRT8KfoeMyGKq
O1Zf7o3nqlocN4Lldus5g/UoEzxA2nvL2F/yy8UYJXiXgiyEFgoCrlg2LamqTG5z
OvzWNFKJ1jDp0e7EyZD5s2hbDm2FhKxfYP6xOP2PbdmCHR15NCNsJQqQMCRy7zev
rcyc3q5nJpfWI/n8/1+ZPKNdVKLgyS/YOSjUMe95g+wXvDRd6iYWmjq+pXXQF36F
0k/I3hy/l5M49NP6lt1N/8QerNZlIh7L0HsYTa+nKqVm5jwvqjOMFVME2faYXGnA
8e00nQaJvu+djj149Pbr+JRWPxOy9JYfw/3GjNh8c3vGEIM5DXutE/V7ra4kF3CV
JRqTfas2nud11CIwrzHdEmIIEyPvuA6rEs89w2LoOJfO2oe01HkBH56pVyUl+2au
ITKB9ymsrZnC2a089hPBm+KS77jzksMP8/frWFbHiPJJ+PWqOOTfiTsvwUf3KHhz
adzNXn3Xw8xKKrmzqJl3qGrKxdYhlV+BXdZsvH0qXUEEn9UL995z/srjnwEgPAdP
DIlv1VHNbaDxqwwBTRowqiZLz8+OLmZ3IrU++IYUeGF/B6UKurbb/naYcKqY68C5
lafdagm1QE374ZmD7PIWL1bfNUZcB3KrTCAXGqKg7/cmonIqXNexA1SvQOcJFsrE
Xj0T7lHdKZPNaTM3Out+AiqhUTsnLwFXrZ4oDXJSHGiN4+AH4bkeQZYBzD8YvnVN
DYNQzeNyKQP5z4M1xC1w0tbytObVwj5rxS8UrQvDxt1WktucCScw4qjQKEj+cdnx
zi2vrm3qk/HWUt9kq+o7EI9eVk9hgoQshzyWBkLehED4t4i9FwGW3qCltP1uflut
lYRkAyiF77e6YtM3Wu/Ox6zcfoLjKYJXlWk3aVXWirZXTN9WJKrveU1jfpMRmW1e
vdxYayWepJBjUzjRfXPBlU2vXblA2YZWMyCdiQjjlVcmri2u9t1qVWqvUm0VYOY3
ERmnwgCZZJaAHiab2mmMe13f/v50p/uFCFLz49CuClCGyRriNxR+5Cfe8S4rZL/4
X/qQrEmB2iF3b/SmFY/6EY1VsYwvlkYx8TjC/dTig7NkdnGX0ujkTNl3TSJzzt2U
NTKSz/AVyhz3+yRIsSBY9m53TLp949Suos49RNDNmKOxuvFj/9+/MsV9rT3w4/mW
aCuPveGgYdt7k7qIyorqxzHbz7i7x9v/hJPAfTth57hoUBlISPzryPrRrYyLcsoT
lFrAXe/5LZ66BJOH3vgmP3AGt9qaAMBcu+fJQSu13Lzv0D4bbf3dr2eJDWixbWxY
QY4OFrmiPNufTwaMk+u+S+QRD2o6DiUEwvMCDJ+sXDAxbCIW0s2m1LmI2LXLQ/9g
wxmv87R89eD+CaSpgkzdZkKct58VMwS5kr/JO0sbOSEG6UaU1NbeA/UbxIqI6YYt
gtlZ0daVeD4qF5ezT1dNse2qV44iUgz8CoDsaEL4L9SOhPI8okPPVfwNQybABUK/
WvEcoJ97tYyFqgpW2CRm9TOVowlengn9CjrBUGS3nQp15EuxQzAN7Q+alGHEgefN
Sk/eVYAN+LBWJMM/iyobSGfbboB0obHmr28+6FmOGD9JGZ/l9IjtNl1+LGB6ftLT
PsXh7PQFYo4HoYbGrFZ/4/r3pDUvrxhzNvAjmBTJPNzlIpCsgZx+6Ob3X7fMMBQR
0g8W7XUiiQMWN3zhMuuJn6LgbIyqEBnAmgwkcFzCjdE1ooEJcgRLps36JZJYu1Ck
dn40vD0L03yUs9Zd28KjRaqwKq0d5PiGQ5zRA+oqPpbII42vd1fEwNwdyfJ+yaTL
z94Osulx1FHZHqT48OogVKWW2Tsw/FIhaRJ5uVcCtcM4FhTfijqrtGVXMDckiTpW
F+D4TLXs6/mzwRJprpdD0+3FzfdESEuwPi7cDV8jkAtbY2QuEgCItCGhjcY//YWa
Hg+gBfiPue+XgD7VzVx8V97wxEhIzvQHaTsuc/VcyIFQwfOiZUodAQq4jKdANBf/
Szlx3V7OC7fHoR24SwnqQjQA7ix7mi6u2z1J6t4E4zDhNoxI2EAt65KyO1InrfFg
cM14AErXUA2HBhJ7PaTuhLJaV0kJvnOl4qiAKIrsr0mIKjXiwqBpSwYjHIQnx+vn
NDzT9DQ70wY/PPpfYS8G2ESi8xKuAC+wAfKnlk6LlB4inicSgu/sK6ynZ2h2u9xc
Y+yt9pTV05nOzx1Z7Izn5N2qfak2iTtW4hTkNOTw6tuUncZGzD9DflbpHaDLceGp
GXNrmeueWgL6KVeziO/Wm/elWQLc0zkG/DTc+gQWE1Lu7LeGwW4v5sIZ6q4snrbD
hkN1aXP8yjf3T5jwRRb/JD1TAC9yAycdHMKSW5aIW+0nQNCruFHrNqHCQNWku2R/
nECYnBqOd/7VB/zaqXP5sei3GIcffz4S3R/jekqjxuQdr7BM4r1yQ/Z9OGV9fCj/
P2TNJ7qcPXu/r+yygX3DSnKQUgSqY27OOVOxuc02GVmP7Y6201+61SWeCwjEAnhZ
8wnsHKZ9PJdptfHFrFcoaz7LFaSWnae9wzSLRfkpioTDz0mqTIA2t63zU29V+L/a
WyDElXG6seIwObA7vdMSnpIv1tFErXU+3WLeBPa0Y5aTx7JCNdnm9duJZmsHLys8
tGtgs2eyllOZourAR2Hw6eA8KgE7cpoKJQG+VHek6IqHW1Pn+UQzr/2OKv2qTQAF
x9y1XPc0ccbm4YvVasvm4Acnpepi/zXLBHWnthRQZzRnX9yJx4ktU/9oVizkitt3
+X8357khj6+9TbBELImupe3BrECuH3R8AM96flcch5CztggPpJeFc2dJ3borehwc
oVT9Atnhmszf+aOHAOnZMUsb4jkY9tdhbWLZp1wGQYtLkxtA7DP2srk4QlQXHlYY
lME3+gxsDHpyAcmN9PA75mcXCBi/wZcAaSmq9/iSLDsWcPshDr4hCZMtKkbvG29f
vgdoQ/oxJ25TmOb9sW7ctLcWdDAACGEHUgtjUqVsHcziHRz/Gxk0wYSSotI0P8y9
YC01iKnm58NTyB+eXjndgxrE+varnixQKv6El7QbjGEP10qPfUL27pRW3HJdSlTJ
Y9CgGbnzrFe2M6sdrPlG0GDVj4X9xFkYc4+xOnONUjNY+v1Z5g5g5j2lER2EbQkj
tfcVRxltScbdgTy3RQRxBtYmZCy0vbFC2cx77ZMWugSJ+SBKV9Uwl5ygK8t949Ro
x/kZBtNehxFJPhTrVPZvuYSafiu2PlSkhet1XlXAy0gvXPNxW2dIFo/BViokOaXl
Pj/VqUM+nRrwRen44DgAMqL+ncMfSk+/nwAORbgUq7CTz4zWzOBxdjmG43JlgarY
kQcOWt396gPdQGVD4eAKG6jccxLlo/bQ73mretF8wLS3rK+6E259/U6Batk+FB4W
4wfpLwAg70K2SJwZCkcfb0jTlM+pDV2mDaJ5WSNtFxyC7VtK4HKYTidF+uf7mLot
rSU8f/RcPN7TuioAUbbPYbPxWbzIGS8udhjq2wmaxkvrNTGXfbKWgm6WF5rNDpX0
D9q7TbtaKWkn4g6G84A6m2ua9cinDgLUZOUDneHNF2dEBbkz4AdpxtPWKCJyG+vx
qEpzWVkwKPxFmEVklz/uF0TwoqwMa0h8i8fRSfJnhPVlaJnHOny/8BygBpt/1BeI
FXzAYXtbw/oYt45KdhSEASRzAPESvjL78AZ2vQSjaIQJRsaon2YH1DLQ42K0y9Cl
mT29kK6hLqbv9MapZpAaJ/QxlW96FdLmg1DnDYcxqgZPM4tAg7StU7btWauiTTX8
ZdzyGf4hgYGzMK2kSju5nIdI/uUiWhMThZ/0Z0QcZx/t0RGyNQ18jSshVFKhIPbP
qW1dnvQUjXu10nr/E2dA9LFH+K6LyOSj5O7Xl2f4oZF/RCVEZfZyiWlI+o3XVTA9
KWQX26luxfB1hIs5Ot9I/WckHD239ELl7h5gL/4dqGVRcWTfbucYM/no9rwdwkQ8
AKBWmb2Q9km6z3W6JPy4zbnHyH1+SQrYSVMGmJWerXsxxWhJESPkaI0A7gWepnUM
rnUXO7cBQnJK9C449kQY8Eo2kHAob+vqkCzKVEPwiNODqabbdzNKemmuhrHgEThF
u40WRlDx/s7JMKzXHbiEa1TjtaPq2faQ8EcJjdKDHHxlmyyX6u6s4YXy1aZm5ixB
fJAs9cGZ1rer21mUrMuToLPbExNz1HH/uRVEWlxVJjUDInFdbrYr3fKzMNPYFi/6
c3wbk3WtQUiqoGy4tx8aNLhBSKrjGbjDY7xe4n3MRodnOTmQE4lgmsuoYS1i1+A5
m1DxbfE9MmuUw7GvRPHr2u9w1gX5OqG8CUjylrmXpOtpFPpoqdcJGetDHF9kBsPI
bYFQBEKpcUtQysJ+gVGSrsF12zv7y4rqo58ahDEmxxsCTjA3N5uBwetuFRXJKULE
xcm3rM23bC8W5/q/0jGCZt58qwKikn6TS5SkFpKRjKJ/kyEe0oAuNbJvKSUZyEsr
CZ665LhN8eL8b4HkCDbZZXGr2kaJmVucBJ61y5A7D+Ro+HhKkClCszL85bCskZga
si/aCogRxkObDJFDQg4X7N8wlzWnzvduFHQhxrLDcDi8aXtm0TlB3YTxpCYV2tm3
W3xztvdsMITGJZS7LrvuY9ODdrY3vLzFhAawDYfhaREzOOT+SFuhZcRBqZbrPlAS
D9fECzBMZyVaZOUf3IETiBGGivvHJksCvPWf7hJ1rYdRlonfFILOgaxJ0zyIxvo4
JsqDALblJp+Wm/6IlL8MRQ13mfQ1ZQSzGA8D2t/CvlH8INb9uJz6gcfDPMRcTLYH
qX2SQLgFpFU2oqmbYczaDRxJWe9jYxAISvNUXVEk43m0brWoC1STO7Y87G7GNdPl
CMDPgxEiHy+o2ISC/8fhXaFKaIttDNfaDwfKSn2H0IcYrLkukQcUCNo6ChEHgaiu
Dvs3L7JmmT/3Ne5NHqAZWQPGmmmIVRfUtwJc7FDfYpqRg6EjGoAaZVqv/TWUblFf
57YR4fdmJD3Z11Tlk6ptsVVziBqumcUiGC8hrxTd6WbydsRpsjLRgwu05h652IOD
wOA97eJVX+Kfv6f9IdOHxqPm34sx3DeNtpHMYJgXSeVha1XYwwgzYlKLAd1/QjNB
kdLGpz0vtjiPcER6SUdAMkk4sS+/2o6oc2/XuSJryBC0Ib/vlmyJGGkwKB506an0
p1bnTEhoWx2Kwm3OAgnrcMKhBkEmk4uFeJa7dYkfJH7VUKV3R4Y2qzelPCf3CXdk
WZJGqIP+DwKdnb/8mRknkHrjepI6jr2aKT1dSr7VuOxVVVekouYL+OuSA/4TN0aL
G2B0NbWbp/eCmJ3P2RlAV0V/NBkdOpLoBjzyItd0/BSKLfv8UUGAorjgh07KVPK8
WoM6DYvdleMDCq4dUQGnJ/ntmey1Yp9jWv/ilP9E4Pp3PNw+ddwaj4awAuVeqcsV
gh5T49/fWPqfRLogdvsr0cpdQw/2CmrGdDoNIuCj4VoM59N7a5O7qgksLApdilz2
Se8rndcKiBNH5F1ztwspF7toRs4hIFUN9rIVD611UkvEsthfeNV2btWrUSxnZZBj
DzAJCy4ZkV5gW9yaInJbTupT+EPXqTbBSosPFHv1mRbkxEhkBmZg6yYHi58Ro/sR
xbt9/DIFxWXPzTdBuhQwnonv5JmFsL+jTbRHoRYIP5wriQYtwuUaUOS8q1v6WkQb
JV3dZgoxVfFrTFZXhaTURKM+jU45oYa1UKZqPUQcVyFQxMOkfHYCS0L8qqYpRG2V
8Cd6j9PjFS8VKVKfhZwn5beXq7JUSAD/dSP7EWJ+dkSFKpJKXxEEyJB9nxwXS5Nr
EJQA42tGVgcJpL0QHJLr/c0p1b36xU0BlUPMcG97A0AXtVUuY7vW9DPVuGjBmCPq
jXqx767v47jqkP/rk9kjbifecKmt2tDUJVjSFfutI01YgBAz7Jl9DPqpw59Opqcq
wMiF7iwiaJlPKMVXFON4q4lOoM2Y9ZZCVdVWMzNdN3wc7mAtwnAaZrjSwgLx/uNd
M/DUgqdNRpBHVnPUv+JQLQsJCqCX+D/haSfG0Vyuz30WL/dYgQ1ujUW4wa22oqvi
cE1dWHBelDm0fPsoP2wZmtKjqxyVwHkJWp/LM+0bKftAyla9zjJPSQtgqwsa64wC
iPffovEajwgxseoFyYPeok3bDoCgEOHnlMZaBOTNBdf+yl0k13jGONeXVVXCs6cO
tv1MydVp0Sz26zlS+D3TaMl0C4iB72onNMwXf4s5HiN5NgPnz5o34aUzrSefzqOO
bJBN60FoKMr1Z0PWb7hyWB9PmAFk2o8x7ZnPpT4HECqZIKQPXtdbseBvfklxzeum
SY/QBpiGfXPP+926uolPFxdP6QZf2exg0ow65k8+4B3mahTSliUOGifF5CcXL70D
1uaNLpuxnjOnfGuzK3FaWkkYurQ2UNy8JBR84e4HGrdRKciUP1rlRU0VzMALk061
gk9pYb09RUSMZ25j2/mS9qPkrwH5yBF2VgneIR6r8RQV0MZRJNNIUl4wKB7mmJt1
qUVOTrseJhfaC5pfjECrT8TYv208gpk2LQSQUibI7O82/QQykFV+wiweFwKdBRVo
vxDC9pWW7TBHy6O1L+EeNldBZMZaKucUJc3StfbfGOgYwupmDSBK/WnJPpIo+9Uo
2FS9yiFHLfBzZw+RPRuw0mOw0MdAmGMoSfnl35uu8ZZO7vsIYcLle/a8vz60PwUR
5wuuUxk5g3TqswPeVuABNWuRmVZAK1QyHCuv83e8Es3q5amNabyH8M8Ya0eC5t9V
4noSfGNp24YzMKc9W/xT0Ympa605q4MUG0bSHM3JAR2pAXvMvy7rfMrProaHlIzG
GTCVhjIEto7xvVx1PFqsgHmw50pfMucbFAMp0nEGgMii9A7i8ssjQPmISO8aZWKI
Ld+mr//V7FaGc7ZvZSNuABdoigdDzTLysikIv5EScQDdl6mDFd6O8d7Tr1OQC24J
I2eh0YwX86c4p6NlYGVHB88WvFwRRpRyk8Po2AXvIdy0WKbGMPEbDww+Q4Vt7zsq
z5O49xQxJPwrD5BE7VKPrQvUJ86l1bLditZ4Th71sq70x4Ro91rpqdr8ytPDTlMr
5NnhgbfncP5/5ZVja6cDx+r4HZgpOPwson3NFasKkzC6texwMq2esArIT6ZXEean
03xpNpaBxSY1UvY56o+kA3MMNEYAZz0CQVuLCdBKJkHwbw4vdRMkzAMi6HYFE0cH
IeqiZIkdUue2Gxm8KsqkuMjH/dqxs9aAAEHlaaEltoXsBz7TE5aX9goYI8a9t1iP
hGthRxcF8DWo6CM1PjPlo4HlsO5tpQ810fMijW2tJqdZBmpwFrRY02Y6N70sKoVr
+zTaWqJf6o/mBCwPn08GW0nbvHEy5JstT41n7Z8L0q4pa7emCObJ97ggP3PR0YAB
rkve96AOcnXCT/taNz3Mb1/PDSyOJVDF5pIua4iNtPPHzxnO2fWVGvK/sepkBoEd
PWMUi6oOFLxYzmj+xUSjTYbbeZcv2ov0LtOiZCDbxVOjngyIE8I5KCjSMe2XUKY3
vXALRmlOmu0ytrC2Jz6afbKp7ILhgGrVxGycRWNfK2VJ+dnIaDCNEzeg8dytX21w
C5dXFXOEcrJjSnEFhVAU2BYd9E3cT17a8TskiAR+9DkSfumqcxCuKzoXcrMcy5Fs
za5W5Gm0HAyF4Vf3q9ku7mrk+cCgNmfAnBNQsw6M+UIPm1uBMhZXW1ohgB7KtEhO
ItoOjpeP5P52fEQhALQvZqVDYFtxi/ypOzDyExZ2GQwDr1EN84qoNqCC1vi8aQjZ
h+U4cKj15m5k7hSfVz1Z/F1Z/36GR80u27mrAhtNw1V3eyAMVNdeDrjp/EblyzCd
EEewUYll/foAuAjl6/c08K7K8MnvQ/iUG8m2LtFLvElXn6hWT8JcrSdeHYIIialx
ZXRzU0w/s8rzozkBxwWzlA6jXqjtVob0XHcxr9628YPi9AbUIYrG+F1EWt1z63o6
xarwIRZBUUNhQQNwaKODSCl+k+g2kIWig7CxZPot2ccBVfnvPKNg/andrsEBxmkR
5LME58qK+FtbHXA+SXxG/r661gnVvvCVxwz4QJktkPz/lWdzpMC0O+e7nH3HET0B
HjZmwPqF4qz0I5wcI41lG1uBe/rrcsFVEoqiu2YJJ1HlEJtGJyw31Fr80tTEzkHu
0iry+QOn22iJXAjrkq01umfWZemK3E60aeB69ao2cF4NWH4fSPGy5VRt6frXm+yD
Ul8MGv5VvDSjrCQ0ATMHyVRgWA3FFov024m4As2s9MFzvcxhNpW3pQnLoVP/ms2Q
/5yW8UeoOTUpZ+IWB/3v1uMUG4sMovg/1YcEzdoNz2zTGvOmDMGeuYHmimhXzQg0
n5w96Rv5vRY5+ZPr/1PB2HnstJ8lcZuXSAxPrCieQYcBOLLafjFzaQbWwysI7mFu
hKEprLHjlg96zMf0Bse2zAk9dN/Fpi0uGeauUusaKGIKLPF7Xvgw2OgK6YV2KEFc
8OzEybhHNvFIilIiupeIYfz9UYgd104cTkigI8iVmxU1S22Lbxh3dBmafUKwfHOs
Kt4Ki3E6pcDPz0MHvZ1WvumYnS8gEI+GSVJ3mv6Te1f9/V0KAfx7FvT7W32yh4JM
ipbaB3oWdC0wl18m8SpRmVG/MteYpt8riN6EiTcYVnawDPMIW0ApGmzl2AiVf/RB
LEKUHh8IOxDdeBfBIdH5mvpt+r5ieJCVLu+9Pm4TbHKhoDxdPpNSpH1AvX4M+mUN
Uo6YFW0B1tZA6ZbwatVrrIItTeYoobG7dIQiPldR0IdU6q7F7NIJENElf9Cg5HIY
3eYZcq3MsUuioM0v9gkoFE0dmLXTB/I9eLjqQCXl1rhKhaPkYhdJlD+HTPr0s55M
F8Ahov2DMpnbXhP64EG1CtDEciVZZe3Njl46I2TT6XyZ+6WAfsCxCHwKiQNkcg/H
0gxw9kw4pthrwGPSvBre1WcVe7C/Cgpocsup8GRvBEomPMoG4FrEs0QZcla2yYnw
gVNPNI7XivyAOFLgR5xbgC1rdHsEhsiaHxFYevNleBnwr+zyHtMaznyyKwWKOa9Y
oBxocUS/4xKCtIZu/RR3tR873zds1DB3YTbNHRudwBNW0ZaZYaiAyDLIATUMjoR6
0D0fcHfZtzUXojJP0Cc2Lap7X3WhM4XQYq3o6qfUZmvEdm1C2C47d5NxKy8IXo/b
OuH7vmioOpinK2GEc5oZ8O5VbLF6voQCJWMGq3VeY05iaPjO3MuUp9i8LSXsXcsy
7125djZIY5428799+K18UKHL7DcWfL+qnLTJrJV663W0lzrS4k9jdI0ked1sC32L
j6+ZvnxQKVzEbthvglKVDTuPstHl9uNnPOL2UnocFxEmrSbwxjKmBknwqEGjoDtb
ZJZSwCJlIPObckGbzsKQsirAOmmtQSbg9FbTSBY9ZQ1t8mGUyk0ghqT+f/61Bvyo
hIlT+lhHPeAbwWZxjeiV6P7h0RCPz8+wb5+s80NVjBkKPB81fCQlPJEbCaQlF4HU
wifxx95aCYbDsAVn4mzRNk7QmhfMEdhhrjxFgcrRvqhF3zHlOe7Kmkw7LpYulLYr
sVuxAkbZygFYuIuOl+AdfzUhQNjFcI0LyXuN3PSYu1DS/q7zlXqBrqF86xCeX+qN
zTIDn9Eb/hOmF8tAQ/BiBo46GSAZKJcOS/KN1D3HTncNo5pjyHdjtLzcbWXiSQwo
dj37KIuUmB1FQL2O7rPsG+JaRMx/fQeiClvlk/7FX8ZtuVsY8FJLgkpzaFqoeXLV
ND8yvtDeEAIPNkC4V4qxAnFmZihOlG/+xve5tm19fQDnftZ+kJFMzbXMEBWRjI9o
uSRU5C5wUccz9wqoi2CtRu14oxNG1VgrDlKJ//MvOt+Ood+UJp5rCU7Xw8xQjXTG
lDXb2DMOeORU+eV2gOSvRSqoM/9Gjk5qPbwPBcdOPD8M4g1E1kFkfJaL6bJ+gX/j
kgImslQo+6azrktrJWzPoN3wQEnoSHrIE2suna9xOwyxz0S0vP4VQPhZ+i3s71rA
3zH33FBaoikMWHlOPVyFSkbk8uwHNwY9TDL3D/kn22/UNgHRGKBN6P1kcQacIS8S
LTUSctcBgFwEsxPtMId4LnwyKZkoNv6eYQUhEkG/ygtzkRTVCsKkarnwBNq4lOSY
6QbYVfp0mvSSY+26Rg3D8zACtoUpq1Stky5foZ3IcG19XcI2y8Oc+Ze/fyw13Jc0
pFQCt/3LsWp09CiUVF1xlJUjI8+DK14ltZ3i7A0UtkvuxGYvkDnK5+udkG86vhkM
KW3HRW5AFisi7C12h8j6oGmDTGqheuXRwaIX4jytstrKUAxU+VwcRT6n3PtdYfmX
K/9d5XAsC7mTFp3NIRCI0X7VPC+VZieidD4Cf50t/PWcsfJ8tpB2uNXZ82Br1/bM
Qpp8DyVBHLD2ChXKbRY6EQKLZE6aSjrTrS6FGSuEnOeArELzWyV8wtcDsL8ipVjm
bDbAI/MDjCMRia4OFMJihHNiu451FeArG1N39pXQ4z4SWY8O+LSfT7ACcs4LYw8u
6n382UExPH+2KLjKKOcIexpMwlxHBevAfMVfPOivqwpuQGA+suL7EMEbZ7j69zT3
V4iHMuIi3d7prig3uGYgeqpF3fbAp05Nxrw0lEUrOMFwZBnLrCudBexlDh78EUg1
JCOpc+ap4vkNg9niQRc+oeoZcOU+UepHuu4JiiIjuChsJY6IuWqs99e05dYLsGNi
TxSFLQt3/Fi5uSx039cASUZ1r9O23lIZvthlpyIQ9ryhE5IWDXkg0Tuqy3T0HSHM
zJ5eO8M2OO0orIdMBQcUSjvpfie46jwHztFR697fq96HUvo4kk/0nr8YT/xOtpJU
YseQjBrL6DViYhde6CtKwvmgKpdOAKmAIssH3cwfo4Q8Lu5Lh2b2L+U9dpXD4TOv
m8HmnNWQ45MOATilMTOP8f9aFi7nuKKimEExUsmUP8C3Jk1k17emwC4b+idTyj7/
u2UskIpvBf+wiZ5qzx8PfJXvb95YX9lZ2nZSPDEYPWLLGlZjjwrb1cwL+N0E4OSL
T3aJ1+j9e53f1ZHD2gchOQV15TkKzHxuGwRdnW8gYZEnN1KZnbKShYoQ6TGQj11n
KBeOYi1BkVuLMZTP2SeCEWMxK9f3bRj4ApqKtrgsz7o+nRanTuk7UCALEgYwAr1g
asaXw64VvUqhW3cBZxdGceKZ7aPw25P25zClpUxZ1sssz0SgGt3reiqGkfbM7NZZ
ZFjZZ56plJJd/vyAlk78BvSjnHGwYlgvx+a870PtWCqdrUX2NZImQSyL4s5nxW2D
+OYn6fJDnEYly6whta4Tn9lRk+Bibj1BU+4S4iZtm4t+/exFTODW09zQ5xPB+t1f
kMbI8AQLQZSnlwsnDqr082XOmEMUoR4+TgnUAahJdaW6Lg5l6hPfc41vtxRzisp3
HzNN1m+wWc1OXDb+5ueIpyu6ppnXT3cMtzw0gfHFB/gDIJ2w4xkGfxqKJ/zgxZU7
64VTwnZMid0mf38VI+tFQCGMS4EiV4bLg2TvE1UBaVu4JyS33eI15ZfLSFIKhzaR
FjIqrLzx/u87845dCsmMAW3nfztGudNwu1HyBD4SfUe1AOVSCWo8cYdGnFEadIB3
BbLnoL1HEWgfUcqYxhDNYs/7J8zPr2nAh1JsjvZRvuOjvNx+VV4sXpTiZ28y5kRG
z+0U3VgtVj645AXx5ZOCN5MXnSHT77yXsVQXTXlweOWrajabkjihEs8f+9FQfL39
xARnjx/30mzb0PgQ2osAAgh3GM/HEmeCcEwGvWOZeu/thC6Mag6Q2zJooxAtRSgT
oPu50YVBO1KkRhQ5GG6WheUKJL8P1U8g/rVdNIoFv6CQ+12BRMDoQtsDg1BR8qj2
EStYggYPA2YESf7mizIk7opemWmyY+8IvKA8MOaGWni1VKFUV+VEXOF7BIljTfsm
wQHLYbFAO9U5tKBKX4GtzhBmcooZGmAXPD84vrh2M29niJR8jMGSStAqwY8IZkr6
MtZT2MEWoLT9+lS+UX1yyush+NKtcxiWuExDe9Iy0gKDYoMY0hYXwbYmWkxS02F0
3onvwStVJ9qdCtDeglF4CzuaNdCnxeAHU7RZXvqs9uQbnPRAZdfM0yxRieUN3Zu0
ANJSAv5IOvOqoGzg53SZH9SRTcC2mhu7NrBN5z6Gc23y08bXp5IzJIf95tkNwXNv
n6hM0avKeCd1Kvjcc3FwhBejiaWnW8vh6RnPaJG5M5btYvCLUoN6OXTGFHxqgPSC
LCUn3GM8BZlFhJKzLZB/4rdxZflc4+vnxPw9oTZH9FTYK/Jqgvlp26kToZzF9O8/
YKDqOSCFYLC7nIFbo4yAN6N2otH88kyDUpLaxFO9xhRrdKXWq/cjvOq+nnspJg15
3h9jFlthJyftgmNQb2fkrvlI18mvKYa3Wlkzm21h/yWSk/TOQ8AZY2y5cA3mpYl6
kV5OBTloFbcb+JWDZJkhrkszxUlpRTl62b9AKIauTUupKtGhOxLOBrx1kItaNms5
KA5y+FJl0pwSOf8JcfWjDuBbhhbb/5iHD/BiA2zxjDFd9S8rtG5qt+ouIQV8s9jP
yHFM2Ms+ZQHZEf34Gg9O+JVa5OxyfQquTD3nVkSNVcaSU1ZkIoIBM9Gv9T6f6HIM
Jx8wCZVZvpqKNlPlYBp7oLa8CKEoBeS+603S+TNivbDvy6+mqOmTXnDJmR8s3hK/
VrpXhg2MtT2tEDvG0nehobgDRRpv78G5kYUP5p197JXCx4Gzz1ulo5WP9s/Cnz6V
MZ2Zr+SLcrTvTrlYHvp+yzHl/iQK21zmoNE5K9hH2WOHcHX2jVg1Lz2+9GcH5Egx
44Lxi1Mil1TRVbqyjebcPDnKoTNr05PBim7IicJCyYBWJxUNZxyP8jvEnN0afXkR
nXP5K0zV1fuvC72w0HYZbkvUySLQTUDUm4AZssxXCWkgcqMfR/mTZFI63rvPjypt
DAzYMLaGSj9BkMxPTsuCLMcDrBr1a+a948SQXyUibjSJEAXY0n/YONRjdCT0Yq3S
Dg0HT1pE8cmqmmocH+pymoIzHdM84KVpcG38lykc1/Dg9u8ZGIMXWo6D5jdB8cXK
mGNC6y4EzkjEySUyM1uzwlWpiwGhgXGmwAHprb/EoxHcb2720AMeDtYvAJqSH94l
E0QyR7IeiyvkfJA0XNC4oVoD4jqF/EEAhhjIV565qrtbin+69FkMh53zNTbQRCqs
Pk+CjctcjWxd64wdDWF14KFWjE4FpnRJGPAb1ttNj05Q1fQDhHRVMcwH648SrzCR
kZaWkIF0K2smFcJHWVK3vyolE4DF8+5Rg4qIAHSLVmZqSjiqznZlHQ3oQ4YWAD34
v1gzIhK4/QfFhA1jmJTl8HpjXZY4ph77h43EHrwRJ7tMXG0mZdtNW6V3SF9mHquH
ZnYqjHQkZecEVPlkiqxKoFsr+13dMAGw863mPNKjzG4wzXV7jCbho2imVhNvQDoK
mhndhX68FYJ1kywN4wD+h6tUhQ4yd8wjaIWHqkMpF75JMZanLQTRCif+m1QWJOTZ
aRmpM0+q/AdyLT6jD5WxiJNCY731UHlEUNwRzFdVQD0K6Bnm5kJk7MS+Di9/IZy1
1TKkMoVLlB7Pk5Wjb/Hcam3jdsKr/fQd8MSsufSru4Tc/5FrkyoXEWW6swP56qoR
xFv5YJon3yDfpU8nNHY0OfRAKYy93lBvbESzX4S6nc+392WU6Wf4bqVo5FsSzdya
/qFxS/nl/dI/gzVXQYysZXlWmUCCJivwq0PTVUnP8Zf3oWp1TMMaSXKULhyBts2w
VKvP3gkRPZjkmYPePQRr8jop0/vI8N/pGJrSm5WnO7D1+HMvfEX9Px1+6pXg4sZS
hS53Me8h0qVODciLq8KTFEiPi1dTg2VDZkAmvjXlswLcBy1FxB/y6YUxB/sMIuAJ
psf1l305EvHmOb410bZ4Zzags22vk+RuTCigxj2vK5oDy2xSTcftXIi9Ee7QFgBs
efyn/CoU/DMZXEex5bECnY5on6WQZZZrIbLsNJ8wWBvsoyA8iJ8antkiSDN272G1
9NVcGcac2mTt+6mQ2MrwxlY8NRrfKL4mz6/memXUERYkMY/n9N/ZK9OpfXfqpPZl
eYj1pHH+8ab55yyEL5MVbjMr/fjoAZoy+ud1kSEMC9w1SN1P3oLGnWZGyX1C662G
MALK4CylHFo2YjCIRehuADGt0Lx1oXzthwrazCI1jb70ArKIv7r+pSDJ/U8liEnG
XZUf05CLJvwOR4UTGpGHVaCbRLTIQ9E/dk0XPUWb/OocKBa4MVmdDQwIlAmU/jDK
hku8Ehk8/+HXDnxInEPAhiQIoT7DuyKGjGtVlFHq9mJBXNB7VaSjeKYBxxnYilQx
RbxDyy085y6ImPqBqidxf9gx6yokHfMh3WeksXEfmZme8E2IHU40qgY5NEBq9ksS
pT8Kf1sApP6IMzc5PevOWyuiT7EUMwXDl24HLuI8InnEWrthA7FhGuU0gH+nbglR
1gSZK06hqn6vfYtHEnP9Kjw1/cYoAv9ka/l8wjJ+3Tj69UpvYf8+wXcFKcXh8uLn
IEptBGGITxtLawWfkXUAVFCwBx1GxaCAnEhzSxS+np5qLYi92njddB9CoZHEdJaA
thFZ0vD5M++TBswiWjcKQ8uRB/LGavYqyvI7VG0mOk/VNsROiZvdF2YXMWBmQaKq
lO8oJA4F+D3EfnkBrZXN12i63cpkbM+P6W/IPC3ANDNbZ/89NcUyHrQkwc/tly8f
nl2+RlCGnN7Z2dKq7H3zilU8NkkwLe2PShQj7EFN5fR7MZET9/kSnYrgIks1Mkih
+kWMjmdXNRKOVDIltqlrEHpdWEmu5sCOOQPRBbcmatIJuav64ARqx6H1l+iSCPA2
NYxG5v1n7CC+0lXcbWIWXKph5JnwF5zCSkC9I5dTBYxfQWoAc9L1MNJYYbrPCPvH
D10EPQYWNwGgXF57Oj/x5NUQVFcrG4Gu5fpLmV1+XPrUivurqpS/u8JPJEwdhm8g
NZGZJuMzNfRRJgdm9TONIKmRZc0XhpO0NtGJRaBadBbOxS7PXSTHvnzYqz7OG9+4
THuEdUkz8Zu8u1GujM+5S2b1N9OviohsrhQd6CzcXjbgDFBJwVyyz201dvrlE2Ve
g8dtqE9RV7+YBSlsH+ZeJjKlwrtstT/6oUInKXu5SgyF2/IWW/tkn+PjWCOpH2er
96dbmpzpqs2/RCGQxFY89xKn1q7a34ED/u080iIxfyLxOC4Mcp9SmrQ/tbMcHEiV
I2wyFQT4ZfaEe9SjXQ0SHZ0w/bIUQ55w9Lgn5OhyEkTyThRcTKTBi+KnVC/7BBf1
H5a17TpobBe9KB7LAlkDvkIilaKC6Xa8HXqcwBlOG16bsLHROU7fBaTGhVln/R7A
3om/V1B7DM2vlm3tLd9NiWbhWOzqnionWegwhNFOOvCODIvUz+uXxdFtem+3+n/2
CRh08fnETKJUC/+6RBA2uWgJnqVYZeXCw+OguwNxgl7HEqH+D5x0FUp2obMyMxjd
BDaP7SbDOYonqhjBi0+3/Ltm0V9ge8zQjkAh3euAET2HDsPpMH+oHPXDkAkR3fT2
R2CIOnzuMO0FgueCg3nJctlVKcAifMYXMX7l3QAska/YMCQxLtIGlrzbk9RhjQja
4+vDcXD+n9UOYlyzHDFuaqjJpxFNQ4c+QL0jDb5AoDkEjVHyD85np8ADTuLnnc0B
xpVZdR7m6qxzTC8XMZ02W+lu+fDJ3gLaWx1tix10gjwS5bxQdE3wtAxGDRAyHMVa
U6c/iemgS3MkdyTwZfBCyL2hDLf/3GZ1hbCpZrvlKoznHPX0NpEO9xEeYIvjQHcg
1uIddr2h/K54AD3T9UxeEoQxr6VmmwlV6wzY75g1x6dN+DDmedTc6L7FaVQiLLN4
pOXWhvooMPhiCHRXAY6v4SZzvzaJ3mumaki0VhN3+ieREw8nTIX5+mdi/StcPY9k
TlL0aTaZN/q/LIOdIbkfk5hCvc97IhHLuFybb/A0OAkgZV69PPz4rivHWXwPUCDY
hvO75Cq0WNoeXExaZkjw8Hi3reC2xhIixXAVBjiQuux+P5DHFLpeAJDhyf/+NI0A
jdH2Hvx9dWwyyVIA0Vx2jHUpuOd7YXLof8L4BDV4kNkZDUfx34pwDekMQ4UYFT7A
S9W9HUiRNqqjGaPja8udRwxcaeRCrSUTlZdXZ+gLE9FmlnMBHjGPc6cJX0bYdH1+
BgPiccbYRsZZJesP1h/MqNJm+1jBqUmfDEPpDQQgNBlQTT7Za2UNwi5OigcIaJZH
bxc7NOf44U2YR5CCQYtGxrkfmuxHHLVYVW2Klonai1NRYeIs7EF3vSRs3BJLYlMZ
3ufvfK9mRlkfKdYsRd4WfI7gHP1ylrkL9wOFtmw9uKLAyMBkjIHTBN9b6pHpqtt6
0+MKSa5am9cTet7lGmNqRWW0/Dl6blSFlUE5lB1twtHmA/HQ03BSeNuhn13GuALu
zKx3r+rq4lhnB+nBVtDy6BIuJ5MVJKJa9BvTgszEVILPkkGWADeYRra4RN+SOVD9
+pJxRig4toI6nv0crq181Iqf/u7/5l/Ko4sP5iXaUOgzXtmInsYkp21bvGUq3A4a
sbE9K+EgsTUAujGxFUKV44V1d2ns2B8DlLa7eiMIVmgNMXjCtXY5rYuLPTI4XeRw
93NrjD7PasqzejBM47UXxOcVYrK4cHq/SO2XC9yX932jjkUj4ci/5KfflEaExDUV
Ey7oISx2tHMYf1iIDLsbIinHzyO+5UR0jPT86BGK1udKUG9K6cfdj5cyR4LBFu4Z
QVoqfrtyc+5cGfHlC7xZD5clphRorqVvKHA451LRD5Bs0N47bgT2bXWoGi03pdM+
9LyEU3fyHNJZELecxTKntRjGPsix/MWAooNxSRCrLJfOZyOnUJh72RNr6KHWDChL
51fs2l3Mx2yAOzqfWFp0Xldrhtzyu2rrV6kg/9QSc9IRAJz9oYwouVgUu+bn4sr7
nCwNV9nWQg4mpESH41x+wr1qS70+lEk/S0PLsmfGZAjhHudAOCryli1AG0hbWaaz
tZ1wX5sV9qYe6PCUMZ2oNM1eyl9TCnF2BgOnHraA9yxV6GMwHzGE0i3HxFlVc3sc
B8twrdly3F10ATQNtArAcdJbQre5J+8D4GLgxCyZStfOe7zUtJJk/n3le1wWVhEX
ORrikvdg0GzZA+7sFgWwcrCbm0LavbvRXQ/RxB+jmY5NEPARf8jWeroBazDC7cet
PkGwWCorLtLzrQ7wU9mRqJiJvA+LBf1JaiigbNZKl+gOFW6WFy6sJncGV9VR3P3r
mVf44CsMfurcoWKoMDDKIICyskur9kjfT8NlXEx2/XZoj33it1K8sih8/tjqx+9n
iP0xS1RfZpINuq812bHs5+vR02FDmj2xAcSHc9H1WNTYliunReI09Y5z4vBiH7Kj
Dt2td21RYdYpnMzpUox75wXN8awkeqtqKKtE4fE5683ZSU2aRitojkqHGCBFF9SH
CL4ddwrYz1fa4ahVL4ZqP2hBk6hSnpifSG3Z7dKrdpUT8bB6us7UIpHF6At+ezb8
RPlgT+aVWs9DIG7uzHb8CgcdJGlfrKwzEzUiPlaWuKUPCk5qn78XwzDABMVkP8av
Lx/0InFubTMmV4Mdcr0JsgUq9FiyVFJ4VHotgDBqrmsTiVFaSqm+janMSHKGhb5Y
idNwVx7N//qjcnfccKlfl6A0gc31aR+6BwSSF5+O3HTG15Ip+bOysWcS4swldJLU
f0S4+3ZgbLLVpj2l7uUYcFTqWAYXYDoIiC1fGE0kfgWajADT+U/6rB1iV2oAAY2S
/YvF1JS0gldkafbAXp7ceKn0p/ZhWL222fngwvZpRx+c6vf3hzE3urOS06irtW6Y
7F01j5yGQUKDOLLt0jNC+T62f8+0c9nCWhL68pvIxw/yj7HXGioB9R/VcYVd+tbV
SWejSrIuvUR6tN58IipQOtF7r2fKYOQ0nN8EIfneD9oXfNK8Y9E25xqsOTJnNrBs
Glo1dCp6JPhDnngCjO/DTZppp0JYkxTNQwrul/9fIfErhkSi0K5fwb+SvSpNxgF+
/B1dqmM/tvZedBovHo1Rj3YihaYG0yaGdLR218YaO9BS+hxTaZckZis+402pFRl6
5fmlWfvRwTFuwBVOeXgc4cyJzCh4gHVwxuV4/T2LiVyXx4GMFzwK4/kuxfQOYUiN
CvHtugZs/p821sAJGlMob8LkFheLHP/EQNCh07tNv8VsGTJd8e6mscOb6yblO31J
0gTyCOlEmc4Ou2s7e993QcBvjbjKn99PPCPTm107RlGFvuCXf/pBHHNa6PGdqt0i
GRn7CHr8fA9HxPE9/sgTvDkN14iXwv3jguiT91XlltCxVEVwCDYPD8l7Hdqp8gW9
zIXA/9OIRljFEMKPJA0aL18fvrzunqM06fHaTLhTkYw+08plisBlA1kAkdhzv1bE
XgnWHX9RftCttzsIQW3+HjYF2TrHsp1ro3ckaGGgCMzg6o8i4GdIgMCuIiNLR4+v
xZnTtmniF9GoNFFPYvKBY48J8YZweNJspQYRuMhEYsxuH0rQUcLbhDfemyLJPOYr
Zg16RwJ3eNZDccj/w7/2BVrPB6GAosbPSMsmdpLstsFEqt5LChGdnd3O5D6K2BS6
jRFiAMBemkFrZGkt+1DbCFAs6TLiNSa8DXdCSv6OKaHJHyJCsA6l+SozUwQwQI8T
zSBjs62pam5T4AsUjEq2z8TktMY8dT6i4KpEid60rFL82d4ZT7HPXKmavcDl/A0t
OAZjoeXZ6dVkhL2+Q0i+tWR0HE4D941bPDKUlRsQBMFeFI+1n0n2llV3p90wh10h
MoYHdRgNAZaYxePcF73m/7gq5s+mPpWdZ8ezD6GukeM7KdM7LyjmY6ndsLA3mNaL
KTz+fjB3sfPNyYMdNRP6+PYjHnHBJ0TW/D8GrI4hq2hC7QbFRRQBBSMGND6OC3mO
I3heZTgyaDH0qPHhN6ejMrByLlzRb/CJUXwtfHTkvWrLaR3RDZvJLIg+W9xeIFeq
QyaE37I8WZ9phMDUrGyUN5uh+xbq37Zzk191dh861Z91UVdd2mYAA9fsvX7uhC7J
wXqCsT+zd2HPCdPid30eywWeUh//Eeg3Q+UMyX+/1g5IcXHPhrSUdKpOxZJ9R5Of
hAkZ5EWg2M5viM+WJvYd5eYf6ZSSI6y9bFGeG0bekFGzv7kqNm8wv6sJvGk/SeaX
eqFiwB9bf77JNsZxbawdBRsbSpmmPA24LULt6Ygjh2pb0Vze+2jujXgU89HST6eM
WMARqMa3kxvib82WLrpL1Ug/FUtJAT52wQjq3a8WYWkfkvYze4HT65eyyR4fGOZ4
0PG72LhWDXryjYU1b9qxyYxTPTSYoA3ZM8jX4xJ1Uxpi5WlN+ZsyCx331FoFn9jS
TWmEnIa2z4RpHgqL5MWSvndTHc+CaPY8bYerv5u0SOTJDAizpSjHtd9rpuV+grG8
736i8F/yQnl9ty6kscklRBFAc+ywXFVm9gMjf+Y8sdSHMp243QfNFQ8cbZA3ck4M
p75R33WTuYnoMFAM/nkOWcXFXGqFRfx7LKUaklPzJRQgZnUeSmtHAPx2bzyrbgG0
jNqWH1XHiFury8Q3CKUK4MaP/mWlRePZhYfYus0dxBpiRx4AYp+OIwBG2L+mvdxh
xRODyFO9qUENJjgicBb1WXzT5qlwJqfhVdrZN1xmU2Qihs7AhK1fL4/lyOzX3VZy
+5rVEly7619WLHVH9i5TXrtVgHt++yKL1o7slh88ZoKWJXr4hoi/xL02FBkCjBkz
CbetQwWrrU2Y0Hb6W8O5sSdH63Rfp9gq/OLLSvd6gqL9009Ko7sVnpF4UayxwzMh
RWOTSdY60zYo5BOG4h+lwKPj/0vC/z9vREMIER2FYXgLSMGYM1bhFrgegYnI8ZCf
tDg1vgNE1R+FckJ26+CmCB+5fjJSqY3VENPFe3DqSP5L1O2+GqsYmgSpOkavSQsB
4eLFXL2dPXsQbZ2kfHi47sQf8XmTAfoej204pfScSKoW2LbrbBUU9rqk5FeGHDzk
/Av2GsXZsINM/H0PPPQVKqKnxu6zP1OzAGC+Y2rXOBXMa98gbgJ3SSWZlwV7ds8w
y3qJq/gWi6CC7mrraDeg0xDh8cqNJsTR10w6YNo/pLrsO91ENk4JG9PTv8VnnkQC
nTOTIknqRaN6MaNWbc1U/VlyqeouEw/WWGusGRJvSnGbVpw9cZTMLp9gig/UxNyb
57CMLZVHnybQesvRLN4DTk64ebkBYPHgU3R/4d7oibWd3DEOwaxfsy5rkyZbEjsN
OynzPO5Gp76cF7TlRpYRYIE5VTs3IAw9UtHhLHk0XbCqwiIS+t3tIi+ZmOJqKc9m
4hg4/VW0hdi++5yUFFSsgH6Pz8pPk96tJwNDd64jVLywSqnycv88phbufYlc1V29
hlhgpyP8tAEHnKnr8Ft9DtcPmuwgypva/wmrj51jQ46yI3krHWJAjGDyEd/Hz+wI
zqGIkFL7BHkdK+AG7t4Gva6KG6PCR+igv80Q5BnDea6EOkwuOseoBjVF7dCJq4nY
egiwr1bMyZPT14Ja7np8il1y3b1Fyja16Kk83L0A5mWMvUlcE9R3/DWeRQUZhI1P
/GpN26KJMiHT8El8rl9WEUm8ZKZAbA0j+Pb/clcuPEZsuej92ve1+TlPSaD39MPa
/cionHe4aSOLgMGc0YvkPQLHJDTKhDTF2KsLgdhbLfcubiEBsDKwJrICwMRqqhOM
vBdxdKQPCa2QpYCYjqra6MjLDbD4UzgZabRCFSWY5XVxuEygfsHTOMJzcGCYdM1H
7j2BcKmzry8SGv3j+7eLJRDUOSCSaKvJBSMl4TDqEW884Zn98hc142pRI1CAkblT
9FdGUZ48wK/79PzfrdORJsRXq2Tqp8FUnvVrZ9lT282ZuYYWMUh4fYREX70LeBJk
xzBkrHehAA9tFC+2yjucMK0/IRhjQVaSJjSWtUv46shUHqXYOGONJ8GXSIsIsh6O
wZn2t7hKb4HjpFF1F12TedIaiot2vblq+MDz4BqQjgxna804Y0j9mxh3YyF+DMyU
/iE/JPLoZbAs0V8hRjAyWng1skxj29WJ3QhPKtnpHa9L4iuDJYeiEIDlVMwbjmUx
ETYJVg3+VjvGM4qsSbf5znyzR5Z/c2o82lp3Z6ya8zmjh+7RITWsDisyic06VRSm
96fnPXsidHMdM1ixMfEs63KqWCKBE0XsRXYdxsubRAslj+L/3+RJYCtD41KH1823
s/GPGIavY1uY5MnF3PHXqYdCqLWcFra4bpf2JktfSqCDfV/dHMYbfVHPoC6QZQOn
U5jLDKLAmGb7DBjZa/zORECIEYi6VmMNwIhZXdwtNw3qmqUTmjNAY47+x0slziXw
sbjblDuQV+ciouL18U/K+j3eQTgsTgyzpVKNI+V9vefbSgjR81cTkvE7q1H3N44B
B02w0mehs80GweB6ZOq1qyDJSgE4KTe0/NSAoL99mWwN8NenAMkXG88nY1X96JmI
Mdfn14G+AXJi+2KxiR+wkYq4SMFqgon9sH9rgHD5VZ7fhQFcJlsKNo+7ajjgPP5S
oJJUh2MwSBAYXx0fgo9ySp50nCZy7WjJH8nKzKVAejS+MXw5o7O4s8Wv53yufwNJ
QYtpnxGkucOjJ9DuB9ojxnZ/DQrtReEfOFp44XuQ5LyXwa2mp/3SdKFTG6axrLaz
UP8jXx0uk0GdBmABz+cW81clW9tFaI+AQHzeIaMB1ChOPVNMdRJnjwCbW/gW3vvP
HYQzqSKUXJ+D875V3lri0w4dUNJ6iVc5kif/fijYGZ1jbiYMj+U9soR1TS39VB33
ealM8ySe9dN9TzQOXyp8bKbNKlxjd9Q0Cnu4/VXg5qod0DOSw+0Qe62Qna87tGM5
VTIxqm84XkmnAfsw5Vbgi/k7tbysmG7C3lwqQeo5WCgLCSqM7JeFueRgAIwdVyuC
fogVa48t351ZZXDIqDeVubXMMWz3ZQy6B6D5hhaqATpxxbL5fKQTnoCu45fUrR7b
ftQrwJinelbLghL5B72LE+O7sTyYSKtUXYl7Tc33WM9OnkZxnyDG0PL1zvhhGXHa
42/oiGWhXBRB/cUkot1ZZscAlaTs7JvV6R1fyfbOB7NftNFjhes7JCJBIBrWwVDh
zVzoVwUOgQTIuFgFEYN3LwNMeNJ+j0WBR9F9v3DwY1eBX/MPnr0CNaCKMBC67qYS
7Z1SK4Eyi601nqGc41trnk/uY3pATg6QkrAVNx3AcxNrtlzq1NWw5U+lpdCtQgSH
V8miJ7u9isZ6cTokASiVdik3M2wHOekBOQloqJxu4u06WKtw4i8dxp4BjxSOuA0P
W2U23YT3s/C7mtju0Y8Dq+cBwCQMYeBSLQ2d3JZ//Rekttma1OxV9Cug0/WfchqE
XLa3ftPrrOY0JXnNqfQfutWdIirJYKvjW6JQRzU9kmXg4rP9RO+hkVOQ7I8CJ5qq
Y/6IDtbNqyU2LjWobQFAF+E89C5KLyhdoXLKPhRiv9hjlPYL5E8EfD/yMfL2jIG2
HNB7iq9WdAiFPHuWKaVZ/h/0Z/MkctPViX64QrBtTSjKQuqPMvryZh2WCklV8E+T
KQVatpo/+9DyejwOHJvifadN9q1TUliKyMk5MxVInk7z4Co8PC1yPbiEyfeEQ/ld
LSj5KQlnqNhR1p02A9BlHbHzMdq19L3nqZTMvl6zYwpM+OVE0ZQsBCi45GBs5jqJ
2S63bsKNfJz7p333HX8EyEIUWJbrOK9X6h2pIfClSExEKc1KrgzWcuJWRgwRNaOu
XA3JqAdmFIF5vD8pWeZUSnjNul0ugYm1yznnqxhssfBdXGY9s/s/LlPoGqi2oXSQ
iybkya6ZqYwxlgjPwHR609927rMcfDUBC9rviVPO9RDNnyTxNIyIRUsot8UjXk22
oeFv7cYeB95y7p/Od2KTEB2f4GAMH6bCLjGau+sJuAaq3SkmYSppS5fQW06CiJ1o
Ajtt69berlO61/AbMmH8iWbnvY156UeqGHsmLcYqKP110tMBySLu/sEgp2FQpXgy
6xasaI4SzYpn0iAKtCCPUkhhapfY1J2GKQeAyZe24B3qSJzdK5uxuQ4tMW65nxUW
McQFpAAKT/GYHjLTn86hSO4Zo1lL71k23ScaWuQkZyICVO2xHU1gYyLTIcpES0A1
0JxtQR22E7xUXCVDvPzLBvumVn7HkDmmY0VM7lZQohRFTkeiEXJ70OB71ZEP2nyN
X3dqOiYnDhuG0BLSYbbWP0bQ2b+KD4hRZzFgUzVJdKGqxlnvpsPwQLXZhxFfJmCK
BThPWKRRB+ImOwKiZsWZaznnBiLKLW1/cHP6ZdUKTmS53zgS3zNzFIJTH+22ntes
8ax9QVEit24iiTuufrDrNWU5L4ZV755ue1UEbJWeK7a2m2rYiyf8SUbrfFSbCgxO
BVFcDIHaB/dXTswLrQGIDG4mZKq5cnKGmDcFEm2XRP7YI0DX8hB6Tosggfbqb6NK
wwRJM3jVrCG8GSgpXptTkS/Rr0Q8rATNTp6b8otwQfIPow9xxYfgrCnKtIt4/svv
K6Ui3W4NzD7Krub8/74uEyf2MMV5EmzMS71iEfRHL0K/4Rzo/PXT06z3YY6LDab7
GHlbnOCoMtIN+C2VkjZy885GIuiZQ+Cg914E2lvef5dm3MfnX6ZKYHi7FlpU3vOC
v9FjHDaMHz+05Y7OPzIsWpAHX70jEg2BI9tyT2oECHOIk6cPbwZfVz8qUar3SiBE
HJshRdiOmi3aKTMSOLp1z+6FgnSXk+RCFDY/8Xju51CQ9Fo64lDRCy/QN7ggX+YI
BYeOaahkIV2QZitIClwY4tOUIlI5D21MXlaYIwzKcxOhMZMKSNx+KOhoWHiqKsd7
loTee+HG8vkWJY36PztEOXkYmc18q+Y8tMrQUU5k+r1pDcl0tgB9wgU2nUNpx7vw
cPkS6H+uqxGB6ydMgyvqY/csOqOqJoB0NOqJT8rCjZc8KFvNJ7f65gaxR+GC0Be+
cOJSJehLzZLeAsGkq+bZOneheXnn7OqZ7O/KYYanWvuGe1jN5uQ4t4VaShIgw/mK
ZG3MbpNZhI/eInBc5radq7G+Wim0tEBRUx40sUpzMyiDkkqvrF7/T9IMCvwgT8cl
ryyK300X96vrLjFMfB0LKvD2sUeVam8Ab3hI5NiayObrCRCrMnrN5p3g5Ddque+e
JY7y1G1gFi0n/bVP2AGg2lHgAp1MUjeZkKFwIRlmB5Is+Teg+nptbEvSJR951kqo
COvIX+i8FOqlhp1ae9vsvBwtxJSA+iAu3Hu/coxZg9Rc16Lf/nQbCFHRPq5x/W5i
hVqhYBYMaaOFtSttngvAv7OSN1ZaLsnkiJ9THMiH1B5v3v0ZMm7ECcS6xu0aLCN4
gKP+7LSpaluhum5JNhOjmQ6hC8A3E86ROH4VZMbNblxFukvfC0UedAYwx3ePKMEu
EHir3Y5HWn0YTBs3oPh/wGtUNIlgeImQ/gwoA2Fs8JL74qtnhsJ/l8kIq2RYf0d2
I2M1Tc791M5eS02j0ubUNCO4LloQXibeI7QUaq+N9CMSgqBBRXhKAuxK6KgWXWzP
i/8kKNTx1cdV87umrNEjYR7BQaBQf/rufQhznhA9Ls6PFQLiPiTqHB5jLoaiAQnX
Z5rEfpmJujLSxOB3sKN4/Znvpr5MlbsKEg1xL8ZL7EHHc64NF+no5C7Wr1fqr/Uu
1I40i/+sLVAuSbppQOHoDqTESvHQ9/YoWq3wdPIX0KrDUDU64sOReiqaIgPVo4zX
9RRnW8sN+nGzP6nlt0Rs8Xw/+W5/KvG+gJYKTtrRo7YkLGj8f+GhqMJtPaoOSQGW
ksQZ3qw4ZkTqoim50tGnE8HhoJYXfmFhUSFZF5FrSVFlTYm1t0TXUI3ZHrpy4XWb
LcHG9xS29JGZeAqrAxEYLH4BnZpawO8n3+iLoirSofLpVyty02mZ1PdWFmNfvrld
a1nTREpfE91VsfyVjMZE5EZS98oJMEj42LKkpG0AaUSJOONSlJPsx9LmFqMGj6i3
KtEU+o1c7h9fAWivROI2L8dVSKvpIdLvA1A3cnSFS1Kg7uojnZg9DJfLSEG322GJ
jykSP4/vrrSA2h+xVC2VCHRgZZZeiqXJO1/BUqu5mbtaQcjCib8ot5g27auNJjAx
auI3XlcAADIlmPagrg8TpfImwv6dwkzcfsXkwofYtFlwvdIG2nEnrOpg8tG79c73
cirq+BGHCwxaERyIn1A/dgwbEl0BHSa/o6NABcU6BBsWob7EwYUPfHuHPdS2HqCm
hn278dGz0Z/5XlSE/qOXHEHrh2MfvfeHYWrr8i18ZPT9dhduJPodlAZ2/+DWiD4Y
qDSCQB3VksuGBpYngbcd4Nexqed0wxsSUZFe01eHdw90TlVYe8hO1oYGx1WFcm/3
xV6aELM9OH1/oE7CnozeEjzV28rQq3nHpp+alfEX/NdodXvGK3w9qQCETsOLJ1xH
yh2hSa5aomQJxniatm+3KpjgfpcLlrW0V2zYVYR7J3AgNS5++zx0iqSQJLpsNe/O
mhGgLnu9LszQkheq+a5eaXeDEOYgKTwd0YE2fXICabvzD18pTL49E8rocLslebeU
CJYl2Abbz0zB9foDqP7y77DIN83+StCxrciti8s1S18ymfXz5Xy8hH4iEjaOw5EL
hLqEWyfTp3/+BvYME22FcjGFn7bs9LMGaQkrQRCgtpKoxIUzIhtQwutwCRVRWQ+j
B7oUG2fTavBMV2csGAiY/C5+ugPNRyaAFzAPPuDDlSM+8YFPrZyqSo5yVcS3fk+G
q6w67WIveoTwMvvNIfFXeovQYaKjSe5JACP61ZWhm/7PRlfJ6alqSSc8ux1xA6PW
1KivX/1ry7t4JIqchxmnCsd8U9Jprobq0Hw1adKvB1l85FOGi8gUQZSgXCoMAI3B
otdw99kJ8bvnwhr1QPBKY6Uc1uaOq4Faxi5zd+I4pIOrD+4IFenYKLHCv9+1915U
cNl7Rn0xu/fwqCAXIQ4eVdYQWTxyly9jcOLXOVGm1K660hGqYHhTLGLMAH4MiREy
ewrZsp1CBO0RN7iWDdRjUXS5gPuprAwDwUJg0N/ESZ/VVwLWI/Ln43fZPzOLAT68
7nnMvlTK0+IIoa+5pC9iQMXLeYCR6lzEApFh45yEV8uO4dinepkKEE4Bew+lqHAe
t/YPZrqX7tujh6VR+WAyz37OegEdceIRg/+zIXqk3FzVWqRwMDGoFRjhyiwrRRfL
APw8cwvRwIZ7O8m0v0dQuBxNvDFrFnKIY4ZzJfWNEHff3Ah0qx0wP8UXzOua5LsB
ay82g9PasxuE1Zokl0gVxvHbeY4r+NEv7o7VIcnqqBf08w9mUjSMdSTv0LUhgKoO
ANqODPfBjotPItPubNTYh7x8YLgFaph59N+T6n9+N8SmFayc4HT5THHKmW/J8HTT
ML35M+e119A1P+Ln5hDK4OZU+kI7JIte7BT4IjXaEFnLIs95ERpGhHSA0yM7kKHs
De1TysSeIiZ/6CY9eKn90BILLVG+5HwCCa3vIQYmtpDK8boWZDF3n7Qc7imZ/uIW
y4+EmNMni6v0X1nHv0clEi/uYt42OUGePfavy1hPw9a93vRXvBslT2K9pjBoWm/I
cCKRCaJv1GBg2hAldpkVWTWhWSMcgygCns7yBv4c8waLqaKP4XJu2ASmdV6oZOUA
sQOThh0LB/yTvMdixDdEHEct73uzDMOEPnbhGfdq26SMWpoMz6iK3sjGF74ldx26
97hY0HUFOkfOuwUivO83lDZi1+tnxPUrKqNRGb3ZFhxaVVW9Bxu4K9FCAYfkOryD
9azKaXX7rCFusP2V5KtQzXs3U0g0cIlww/uF/UAVdJmIyIKwsLsu/CCSwnQ3Tght
m97AAi0FuEhIPKHolWIzC2w/uq1n5Idp0BzLqYIUSNFS0vvtfUJ9baBcw8qaH2AF
1mW5KcLGPV7MdMIHnbJctDMMgMVelQt+EJUmCq/LwY+DFsEl38OIgeGZjJa9q2+U
MdjvuyA9OqhHHKCDIDre6k9e1wrfMdrvdU3LckcTFz5boVVyXOt/QLd52jtsU8CA
uRs3D4thZJzlDssJZmtF0/lNdom6RlabZTRtBqU2E75db33zQdmQyuMat4nFsZIS
h2/Q0C9ylKmooKQW+xkNzuf25v7bcHHuUX3X4vPheTkvhsai6442ZNDQFHfXcvsK
39wV9cjss7nVv54KkCXbOt+hr2kM1K6+wWA+//iO3UYMzd3ME0FeuQOzear9rTFS
OUGhghefKw/wL0ketbZ83zRoGwAqe/oUjLOH48BdVRzggef6u6f3+CHxD03cuRO0
dohNvoMpWKSpOrMrjfbhGCAeggLHSCk9QTtydKVSue7Om95IASs3DVjPQfZB8J2A
HnhE4tXTppYgh//ByH6i8Lv8pZJV9G16tBS2eKXx7+Q/Vyv5ZByyel8MomLLNIaV
LBWDEG/S24BsSl1VmMV2k4w5dHPt4+3Nb7bEsK67lkWQgu3MMxT/sQQOYLYV593h
1pC0pq/XtC0TDOle1f0ZhgTOsfhXZHWDxtNdLpcFzDBB19UB8owgylsRD0eod3KA
BKbtY0OIlC5JMX/oZ1hve6ENi060E66+D291chhcj7iVTYcd0s934d4JMMrldI4L
tLgoO4WQwMz9W/Fhf5QuQduH2i449Dlro4W+KqFyx5mZjfitQ0ZqUVWWTbuj+Bdu
HzWjQuaL6lzA4rHSBgiwJsu8bex3Y5Onh7swjHUxXJp+ntorl7tmIHLYff8D0n7Y
cAxtWNTWKVBuLdRjGjz6aubswHhXVQ1PiWgbFGnU7rE6731F2QeMwllp8nOiogDc
LcojV36v+U9A/RKTcWUF2EUu7J3hHeRlU5zbgkIlaGes1jqkEn/kyZipcmVxHzXU
Zmo++U0wS/maniWZNn4C8sAOzWkv9gA6d6/4vLLwCC+Jl1niJP+2JHaZdvyk/4v9
RJEaYxygYjMetyzS9nM+PTgjBIi/cLX/poiE7iH9Q6etI+AfroiW+kno3E2ozAsE
aW7rYW2MAJ+Q7AdERYeXMF72RlcdyoN87zXQ6DsMBxg1kiBTNWHj2/SEsc+npuFf
Cv1By7nkGFf85FWcTFhf000+/cBnkA9jmm2+uNd4Z6oKWSPnIdkrE1ps9/t1Do7b
7chyKiRCoZMeaeRSEkNPooUsUJUn/rBHRSZhXvFdcG18PI0CsdiKHzVpxvmoehSC
3/lhEvlxREs60xi6CtgYegjqoXIZMCgebckmmuoUXnAwAPzAsV1sj/er9vqX7kPz
2oCx6YZsqoT4PA5kURc3K6DxaBgLnIZ4qLh7sLmwbUqG72dS0uIWU12zkIGbQdTJ
DJyOWeeIS+tqUtWCfgYyb9q5fsXy7zmSlAe85OQ0aTEYg49sREe/N3RCKLlyvNNs
o1NLlviZfWFYMDIVmmtMTVMQczW0lWB6n7PNkKwY5uHgOxvSas9UzM5pzwiAdOhE
eGQIqLJ0tjQFLd1sz9Y313k1QjUhZa/4i8Vdfch954TAXnCeZ163Y3LIEqzFMRIP
wV8JxY5/j0oYxX4dWbCYwqjEvYRS3uzXF3CofN8JaxkrdhYL7pMf+ODzjFGvpilO
sA2Irke88tSe9/20hb/nne6PpPhP/vdrkUjBoJI/zSPrijAM1jVzI7fiUdBYBk1F
nwjw66qzoAHB2PRnqGapeElnmKt35Os/GnQJGHtSRKif0l6cQGHJNWrQ0sODuw1T
ZXiE9CQNNL41VTuYpbGps6ZFIA35737znW85d4O95HEjBvOeUKHLfANCcPvz84sv
QbDfcrMG526fOhrmRLLWNWr9XFdzHpSv/vggH6L/ObdqYGcGXzJp26HnZq6LnpjO
2hWMYXrVxFeKLUj7oAQd9Jk74X1BPSNaklkyCZX8fjrA2yq945ejnD+MYhW8EZjw
dExFc+biyWlW3CgzF1/MO5j2whELSAMuMxrI7wDpnWyPimEJY4zYifiuYfvfNJEW
itX70RGULsMLcciGiGrnRsh3vAU6GhA6Xc5k1kVc1Ty0lSo65MEOelfH344rb5Vr
fFC9cKZHvXULtkIeVt0bUe9rbLHDZuOcRDDRrmVWXws0oIPXSLQduam6PB6lOla9
pGwelcGlfxeX81fY7c19QSr18LX6L/87/6q3U72/xF8bE5SKA8MLqafmfQt8HeBy
Cb25FUbxkzlqTTpUvRJgUii7kTf6ntv28K69i4FxNpYH5vPHHU5Znh6TplB62hJ6
QnWsqc1r3RfiMkPQvwjyzBCGx8gMJUmHNrL0h3gdoAR7bLF6QJOhnQEerZR1a+n/
Gcv/gWqpdrh5gg+vwcURLoRWPA5f8aqJ8GD8wXEJskc5OdCRv7zxp5ipsZMibV4B
OqVFTkg2EWWzVQ5NCnfYSrld7oEzyi5aIAEAuW3Exx7QyFowHvv/doNgB42Y1rfH
PS2DSUL6pV+oFP+7QYgSIeWf+CIZsoLJ6+JI9UFZby5zVOlLt7yoB6bsvUsDhbj5
owaqEALMWo0W9ZM3mRx2NdXt77lPDIH5vCMBc9NMI5xxjekoAtaqEhAqOvITzvDp
/pFhGP1hhsbjXDPZ17Ftlc+rsZm4ylWnolYBF96wVTrKaKywUeSbVE59iOk6Q+SQ
s6RghJb9kvhba+Aw1JTWAJh+h0IDgvWT7lFT0Bf9CBqfF0733WFnngGeOeQ/lkmG
AhsT3sCSScLspHHV7mZeobkjSn/TSgXUSpkkMTvK0LpuTWWzIgEsRFNC2Gz7kJa2
H1oh+jR6jCnmIfKocJ1a/fNEOcWGY7OLhLCFxQA3iudQZ8NHMMjbRXUq9/ttSwNR
ye2S1wSjY+y32UCsfdqvxb5v1V6JvVL7rdnhG4N1Cr/JzhcuT8KtKZwZEtVq15iY
nFitRM6N1hxmWvaObf2F43MdRsKOZ9RIKfcKkvnNGan1Clm+ZWqgS3zihUGkVCUD
s7zQloSjd8Xjvhks7C+HCWwCx7o+ftmQq+CwmhrwUAyv9Wf71aBWXdxBEYIvAECo
Zg1naSliQ6Ko6VsOOhZfhI5ROgbw8En1yXlM0ZPLaon+LGCEy8QNw3B7sHpTGdyS
2nUxx47GOsZM0evsTe45bvRvOxvVweGWSOsqwTupnch6Q/28E9VREoZS+P4eqwy1
COLAyEoubQnl2yF+VtAsxFZFVXbIKKbL678GUyIOUhZI3QuFYlHlHiQMtqdmHN/w
pRSJstnXPFAgKOKSvF9uiqltWUwMwMGnKGIQBOdsIlGgTB9iPPH6NPyEd5NiRR/y
ZYKz0yY1awE4/aMfgFv62WvPQvvo6N7j1rMDWLfTkfk5TbashMOBFgmBzpSPmFYn
FWfoLn/lprerPECioBO0tivo6cJjlTZ0ukBO0K8ulpjQBeIDM2gWSuL0IR9hO7M6
b4i729XKcDSoXt0gs8UIpXpr2GKMvBvjpNgCAjLbi1D/MEN7UVM40mYKNONtoJNs
PLALBvKXRoI90hTJEaJS/QqiIOgtaCi954m7wJiLicpvdrProkkSe/P+8d2CB/+w
4QWCcyPC/q2XQCdHbg2LqXnRvtyNdYklssSlj9cMsf3tPohhlc0owKJSjQ22BYWT
iinY+jfXKJicOcQfxKHvjmWm2JiW3N8yCDKoq6YhPQGAB2ii6DIHkrUom0lh9/RV
U0MRjJ+zLjFFSUkt87GN4f73DapB0ZLTMFn7x0oG8KoXuvncSVzSmeQH4g1eZ0Qs
HiIBaRIgCeArCPtgH3SYlbG45jQhFU85nxzcxSmk+UsijxfXDuak+eDm+z0C3HsW
aV/6Juajj4PYWrt16JTt7CSWVlami/9QzRohf747IA3yFQuNzTU4aOP/U6NZTl9I
YnihJgVvQq2j21d4wOe/bH4MJxF0jJT7VwtmWR7GXrJl8n9f6imdRNkH8Y/z4e8m
JfyFTShKMeOmdW12gpc3gtP/rfmQbhZTQprVLeBHfU3uB8GGi/bx7mdIBWmbxwbX
pUJEb2oTeoFc6xYSytjz849QXUFBm5unRrYDGVnroON1ETwsh3Q5t/8zSEH+M+Yg
uLKAp7DOf/TzLkshi5jltkCBTm23K7N75TXPJ8BRBsVL3U7dGwjQNVQ1pTmbwy/I
7OUBx1K8nsVkLnVDdHvvKNoz32GBViOy+Qw5yq4nDGERJcekk4Pf8nzKf4C9u5+2
QwxafNAra57SxUJUdhCicdzr4NnmJeigrT6dEM1HUzgsovWWwXV7r4rP6MxgZrLk
lh+2QZNmI6cRI5QfryNHhmuZdBZF3tilFcqz8pA2Fs8JkCwkAlKfwna9xxwpuOnm
d94Cn7O2M8HPj3U+8ioUO6FNfl1+K1TwuVAJaOzlSnZeTS9AOID06ArKpDz7RSqD
jyIi6o62Z/mwQEA27JGd6CrXLH7dRyve0oLnTl81TB/m+x1dFj1zFXb5wRab+NiM
xnxIazsoIG3V49Y63D/OkkYCX7Xlvj3u5euW/5jBrt9xpwx0Qltey5POVwmtYCnM
RtpIu46rykXIX38WAUlhNeJI9nmcLxug06u99VcBjCSvd6JhM+Hq256Ob+XoSksE
mbWjISRjHOm/f27PNLLAuHdgPJD0710F8ZmLyJ5qQZJrO96yxKy874mJ3zAsvz3I
M1oKKjhnV3aZ55RwMo8gOFx9m1TnFrt4LDIW0wYbX3/vyQh9zmbuok2vEoWX+fJW
XNvFgy5+vcO4jPtsPIAj58bf0SPelyVBcXfFQUV86N64rFIXcqhSfUGNcJqDap+f
BBOHxW4Mf2ecNH9BcfbzApjPHBAWGLPEF/2ARXo3rlAyvdBzCP3ddnkzyQGik8dv
RTGtxYRwyM0Gj4Dw4JZnxil0+4qFJOkxqPFYLnJvZ6onZM+sTmaPD2mhbCN/b8Pl
E8IYOXoHwy5NDv5cqnxHeZMp/3gh2PKM51J6j5MMWytrl7qcKdw9dLnTmMtS5Mek
+UFIDfut1XQKMdtK8yNc/2hzSZUrn9Zm1ePkUNvB/2Vth64uUop9/LK9jY7NLHs/
c48/kt0D5AV/C3ofXiBG1Ja0VGj6F5Dvl0tNWDe/SpmJokq6dl7Wk5Op43UIIhV8
69gt8dhGc0vIGr6LNjV22aiKX51blfr06lnB95Hl8FoL7rVqw69OUxl7fimcvpra
mMjd+pmkBI6sZC1+P4wmbzn5jpDj2qmwBusnFjEOFB5Db94r+YroU4MWdPhJ0aaS
2RXxmxcUjBkafj3nA3gYQTUW3pOnBA99lbf3J1X+ajzM3KsvGIgZAcxuO60OzkLI
gCnfU37Lxy327ej31Q602Nefxi1w2gqmn7SP7Fh45zVX1TSiCLFtybP1egoeY4ND
/BhW9ZEdE8W228DVf87lhkLYCke9jlJsZ8Um5spPNBeNFDVASk83I0d9loQztLsC
wLBt+MMuKxKKhgcDZSGMr4+hjfRY4EesMnaTMCdKnbuzLz9Wkg9HgyFNDGmAs5d6
MjSXeQJTRi8+37BW0eAsGIA9RFR6A4jA1Zu6fVdAHxvQ+bXSS4u1JFZU9JmmHtI8
aBts6e+NUjUVZdLaQpHdhq9loZx7otDHNZ79eZfmlt7eoAHFijGaVLZ1wxjMIRa0
WAgqXZHgnsm5XhqQAudaMcPDuPrgYqLncaX7RonuYjBiYkRnRyj4cHaD3MXO3pC1
dn5p0KWDnPZkKHib0CovT9QNqwOCWUW0X8cDNh7P6pvfllyxiWrOZX+axloOUgC9
EJQcDYi+qqgP+Jc8nLU45Ogs5ZkfA6SfWKQivW5eJQzUw3lCRJEnzvmx9ivQzC8L
CGUOGiOzFYLX+JYujc5uGcKiVKa23stPmHjCtSDY1zhBITbOP3w9kbifSjO6Eoab
uRD4kCEn6qWsddWSs8X6VS6PIhdTm/raEz/rLcCY3oP0rbDIPj4hLlwvrOYG1M9Z
iKz2ZXVITSuAA6XbUaFU76HK8m4erCKv5RJhgjEjmCMK3XbAHUpN4WgsCRCyoePU
sPh9iCCXehdT5CKXKhC2BtS0+KN9t/BdSAaLAcInMuslHKS7SbIJk3SAKsw7BtL4
9ctaUa1mZIOzZz8fBfPVD8PUzrvGDypzjlKHzcpY7e8VKQ8/cT2alhrzaJ+W/r8t
gsLrhnml5dPJGdxFx8Ix5Vm+RtjYrVj0/IjSDKCZOOfB2fcJTgzd/bKZgup0sGn6
UR+doAAOMcGGDTIS/ruqheFVXsIEiKesV/o/zNr83yflp74WEjm3uOc9K3JiBpqN
3yyoBL6fs7sp5GKBnOlhDv2IutmBjMNov4n3APSvQsGBfqjUQMBb9+wAkrCEaADk
V5oNctu+k8jHQm75TzCOouSE08mNW6o739wYXCiVWgMnR0Z8CHo1GO1ifnP30/cL
aGRb0Vq3QyQfpPE5ba4HB6pTXgZA0zSwoHUWwNphVc+1gzzesYyyOkpfLOVB5jfX
8IE+j+wLHQqKD5OjG/ezqK4vpGO6eSEaPUPcYAIuyEAnwTuaMcmj3s20pWgrUD1Y
N3uYj1tFfjwokboSGO2DFVNo9QIhuqYIjViNz9Zd/lXqGBzm3q1cuAzJCneCmcB9
OfsfVoXUGPbNUpBGaCd+bqlmKriVfSQZVV7zzqyFlm8wpsVWieEor1eE7FldMWCr
0vU92tm1wktHjsXGq9BagsSBGLy9SCZKPbjVzuQMDZXKP6tERdvWKrTEFj5/3zxh
TRWOrC7Fr4bI0gCCb55aG/t5XyuBs/V3vZD25RCOmsUPLbrIfCB3H4RIn33Nicij
uvcPBDPf715LidYpM6XQhcV+jYXdg4x97BIeDOgDJCpu94rQG+buxnTaCKaNwmGB
izw3OFtpJuVm3eG7pzlMJ6cVj7pp83DJgM2K5+VmhC8mT5uUdxVea0yfx7LO6nwP
AG6WQ4U5xkV9IXWdpPZWvRtmMb3btIRkm6vJNxSPnWAA6zOeaMlsSy8mRcyGOIk7
mqSwuNSZ2EEtmi4LRGVOkIWxI/uLbAVc0uyHOZMTuSPZ9n+G5ZNGUCh59zXj41nB
w2QTJ+zi6SrPZ77BSx/RKiU/YMZdh7qhu3jqkDPCh3wiQV4ckhIFeVL115y9zBPG
ius0rFlJTZRA1zWRD9q3NeRCp1k0kmwrAYW1zSE0dLZy9KEwkqOLKJOgBMmxHEOt
2UcIHsNvf6CuRYpRINRVjMtlo+GkC281w9pnpJi6jgkjEyLnQmsi9xVO1bvExZx8
Pyfub8vfhPyz9X8rEhNWrEczEMhDTmnABoit1GZzgyMrBSmNL1emq317X2tMsUd1
h9CC4V8Ux9ehVNZE6CGc8jutPe7n2ToVrlsV7BqXLx+l7k3EwIbgLY75k2smg7aB
B8fI7NlGdzZ1KIA9vl+L4g9B8oOThAApZVznoAeS7Q+ZWqqLTTh7uHG/QVxhJPji
dnedr31TVua87pJis2DImIgHj4d5SrWMycKf7B7ehcbtrXvHQUmArDu/b8dYTLF9
/HYUDLHFdZ+qOgRY+VC+1zZxaOLupJr+nJ6AhhaRa29d+rInNOX5qEeYP6nEuyyo
kwnc/HL67apM+aAqv3A2+GHcgRe5KUmw4UCEaPQhlxBoKctqHFzxdhPJenJ5pz5+
jJiyf1DsC3MJ9JQytK2JvcWf38q9oAbLmepYUqR9+em4r4X/Z50fyRZe5JtXLZOl
AdUUesnUT0XyIvydZPXRb/cWZYZV/SShH13BR6Ch4L+xwls0JmCv2Wr0jqtqHHiO
XatS6j0AY+rnfw7lkJsyXWkGVAqyWPK5IdUv9gZGtIhbjhtwU275XhvsSWFPdheH
yqUmJmOXO2HsBihwbv3Zx+466c1ZRmu+muibFpiwB8f58bBJdCR8vGr7egToGRML
0dtmd64h4cOdoMcAx2edtvswFY15REG/YtZ232RvNtopwLkMvZh3o0XCSKe3ZKXY
yDhhJRNa1AGrZS7Rz/LXk2BnQeKuHqbCj8dCTrZJOayIDAL1yuxz9L2ocJHEGR1F
3grtN/pKLiVQwWwIV9Yfpyvj5rjNKCSk3+HkpqczVF5S0SPOUqetF5ciP2L3f8hZ
R8Y1gZPaD2ah4Sxi965am/xLYar1CVcHUKsurcQc2+nRX19rDlk7hIfNZ4Y5eWF3
B0YXH2luhnQylaaq0eT0GooczvnH0G/5yNRQYVwtUUtysUWR2LFvKhh29QQPENXN
FhfeGr07eI+0ED/tq7xcY+cXVvobp5aaI7QL1edOjlaIdUyFuPZq7YIk7bMEymWn
N9mvAlI0iKyejQ0GlBF8rbYlvlMgsxvv7viViYRSzdCHUduTBIr57J9aFZ5Kt93O
gdOfSTLArzl+T5UkSQi6futFz9NWwdXWQt5HOP5xYVaHoCPRzuLLyfswBmNirWTQ
LHw8zb9zi0MN16zmEhUSLtyrufStf8PsDrNlm3rpvatfS/8BLVWuuLTQk0Q1DvsC
iT5FPqlSY4FfDiOzOtH40nFfqtoyUt9V1ntSNrhDHfrCcREY9I0RjtXigxCxX90R
6MhHOnSZtAZq4mzyFu3974qKiceVvAd+Ql6ciVtpUJGnGLLycUG+QaLbF2P0KrQg
cHVwr+BESLLJcHGrprPGe4RV3NB2+6hAkfNtAg4DgFP4q1mjd7WoZZiN0YH3yP+n
lvROR+9cFCL9oHTShXSZk2HuSzeKQsizFSyTaExZbN05Q3rDxE/9akBJ284zRJi3
PgGxImWmlL+9REukPCpv3MmLXFra1iBtZKSD4Y2ceRl3zA3o2u0aBxKU8q2vVRJs
kMXfTJDOWymj0qg6zcOQ5PP9TR1s0AJIr+KnAeXfs2/WUdpRRkjMdyP1Nu5sNm7b
vusTIW1BLb0xM7jfe5iaU7RT7Q0f+usGMa2EoWHxuFuOVV/rqoaJPtwVQhVJOqPG
VG1bygBXKm/wCOR6U64jLtB2dj35aqXzrfutra5WFoj2JmStOnZHpDoA+k+FpD1T
hAMKT8UYylZsalNubCFAZnHqAaVFa80rGlxwl+k8rUTxsJllH4X4ywRqTHtakV6Q
MZQKTKffVstleHRH5Sw+zt0Kf/mwl2VJUX+u5G4ObB9mRMgYQWNSqvCSqXzH7GCL
IqVCErH7x3EvYWKDXAx2IrV/xYjHY5dg85yQS49tURGoFagdnXq4b974DsTNPsKB
v/9k9ctL0J4ggPhzmsZ+VwLqP/jolZv+A5+nsmszsub7tU0mB1EZORyxtRw5vTqQ
arRjwup3w0MDlaVYsTMQEEs47MQsCSZKh4meImF/UzyyRc+/9g1pHS1lmKhSokiB
IxJNq+QOwd+GYX0H7wZh3+780bybD5ptC72zE/knNQbFcsT8XgM8DUE7awajX2yW
qwZf4BoiFFsZ9XnBfsoSor9LyrPcWh3A/0bTNVPsIEbaMRl9//DwMMt81GGoDkOq
eQvdpt00DWGY5L/ErockJh1K1S5F1TDUIrWPa7166NmG6bsvVgVOmQPcoraTSAMO
YTPWSjbXDMiBN3yWCOIYH78HMW9K4ngMjuwqOl6VDUEtyJVYGTpW3L2CcJdf0o9x
UpHlOdd7sNvflunpYU0O8KNoMoVjBlwOmdKRJmjvbzTwGiF1gdVcEKyfJYL347WK
0Bpk1AKNFrVWPItSd+rs7LKIFXcxrFSjJ6qfZLJHmqqCFcyIy9Zn+Io4uGBV9L9U
5aQIvDGLJLQt2mOpG0QJugZy7fzlYgQPBZmHBDxvEMg+TLdJmwELoJkiS4DKMYq8
5PjdN1FjwcajrIkr5dLhstaXJYCS95yfJ9IiogJiGJDGyDtWZ2WYTtqSdL89cEcJ
RMYxGtxVa12wVj4fZvt3I3yFD/S1s7m/zoILhVFmaU6vn4OEc1l+lkQal5LEZQ0I
tpUS29mtomgsmoKe8tWrrsGxiZUBLcGXEBWrOvcsPFnXpRD1w4wL+EKRfE0zG1Hc
Zaxbe7LphsiK42MARxwOV+ccKk5CvJ7NIiBexBZaUcCeIdaopj5U7ID9IrKQqZOO
tVJhDf1L8sY4SKbYHYeNnvdCxxE+Eubu3guCRwKz4g53w/gNTnIdovxtXK5ErPUM
LyftQmJUkUnwjCwkoHneWy0Ni0M6g9uqezY6tt1P5lANm0y7MMXfj0MvqpsKFqgF
x+CbSr6R8EFr1aPZ0+A2JJjZyqRMEmjWPfHyjgVWFMkKWEDNsn+w+YRiDx/OLUY8
GswbC+/PBCaS0aDM6fv1wmk0EQO5BprPLuvj/lLCNkbi9liFmRQ3L8jR5axezPY1
skfUVOOmvdYCK6Cgq0GAAeR519TJSUbVA4GQ5xNYmFrfVcwwppywIRc2r5HXBjK7
sQ2vfYIREoHoiVAD+vkTPRP67/ifPS9++A7TfyyNvTqWzYJTa5RhUr6aFNxq0Ljx
iLFP1yBdiQPNzJ0LEnJ2Ndf1GEBEH1dk4LId9dZ2Gkhza9Z4P4+9zbzEJdgm2TMM
xBQRYnkoaklGAmElryvsh/UqMKvFWUeAJyiDhpFvEzvH9LW7LAQZWmeU44qqgdrB
+amqqH0AYa6zrSeVvyqnCGnkuObfwV7gfea3h8K+ZinzrcJTt9Lb4h1x83Ye8WBI
CAErF2iRi34otEWcqRqHxGm4ufgOwoRe/vmnVScBU0uyxRd5abzyY2QRKMi+mfoa
AMJLjqe8oZ9I0nAavoSOKiz31YmRVCAKQXspX5wSe3vj7dJm71L1gk0S0ARXOhPR
KmFqFbkuJ9Q5aUPQ0vH+lPHoEzE24KQeOdGRlnH4nFI4hY9RD/mDV1GTnO8e6xHE
ljUn+N0nYzYMpz1P5aW3lHYTNn5NOs+fKc+2HnMp391QCD17cDk1Z9wGgDwV2aZb
7QnIPEsFtTm8xUgrwAHTcV0eYr4ASnXBNQXuaFPSMqpRjW5MGLcALcD7YwCglBZ9
cm4ntJ/FyBTlQTK9RmdIZLOliMhHv7uXsjLd3RZsc1MwVDVglPtU2Mxj4L96xBHy
9WInM1BDAz/V4Jl7v0VuvCnn5jMo0EemB9cy7kB/QGFRknS4nCehl3DbmRRRM/mp
KF8CcHaTrmVFE5Ruwk/VoocHaWoGOtsi/dw+EtqCjr9CYvIBLz3EWAh5wLcDzUfz
PeGnYFBKFeF1B1LuCk8PMABkEFTBkZShgi4uJo3sinrxdXb66HFltDaRR8iAmysH
2UuC46YlH7ThsKFTFBtA4ZZBYuvn0b3jcGOv8htiRvZUzIZkGcYmQ9TtLYiwj5AM
qufAYLiRgEgD4CufvBsBdX3WETCifqcaTX4biE/uUSmijMlN05QHl7AsnYIi2GQZ
xg514Yh6o4l5KDK3Xo7zp6IB4s6xFryHQU+UHbDVUvH65AcLyAj6Yb3M7Uo9gIU+
VEM3ah36VUSzLzYeZOB4u5IqUeiLzmbFVPnfK8STCJvX0ziyQ7oJX2K2AR4gUbJk
2dNJ97GuBcsp4iNuS6GqZiVJ5Ao6DvCmN9VzYVR7NwMD9kDTLaBIRaMUDEXAxts4
+EFQ16oH9ykK/6JlZj1JRVTOOon+3HbBgUov/AAlwSDK2N0wXOKIJ1cm2OuVRVlZ
HPn+n1soiHbFpJN13L0IkzaUcOtptrnxvJliB9/tH7rPViDpUq9CRY+WFngfS4xG
Np5+MxG8JTNzi4qPq/eQq9XWEbI2rb46ZVF4jMaLJ6TDWVbaPH0PtH7MuYE3MkwA
8J2QZ/j2UNcPdWjT/6pdQgfdeHFZO/wWzoZwsJS/BaRVUrKWOewpqvpdLGTwe6c0
LNKrfCg5dAvDPq818hQC3yKq94WcKh4WPLeTV2GbbHdV3W6AjqVzezZSNaCuaOB4
iFIH1adiCS944OBQSKKhSHatKdOGqHdF2GPslPvYgBN3qz47ZKJkvhY3Uo8CzTrf
2gQ6H9kCycSC1lsvsF2e1WlqSZa04WH7b8HtsmaPTetx9BvbbleFczHVuPRcV8g1
ifqEril8/6T/jsRvMDVjPDi1ZX1IC8JOHgrUagdiAOy8eofrMZm3vwDpiy2YPowV
GhZ0Pz8iY+10e44fJu9wBMZREzDM5s8AA9dh8vgQF0sXa0za8f3EGQBFpmsF+o4b
t2u2qZXN7trjst6rJg2UaDdt9X5OY8uud870xY/f5DjVNZiIc4u3qgMMlry3wYLq
SIdHGlCEMHIhS7PQGYBHhqsJdTp30jpSmo2Hy84Hz87+cV938xzNERc3OlkaY1EE
NtSBd+IyiSjYWGdXM+aRqr5gAa2vzFUcNkcuqAQ4Qrxre8p9+HmCZhXVX2gKVJlg
VNsWZnPyLkunvM7QlfSSWxQcKajoF8WRWm/DCOqaPPDI2ifViEbqqX3mYmN/XQWj
yie7/0CToPely6/TlhrDyg08KnoFxln1BBeVtc1zYoFTUZ1QU1XMmo2of12xP58W
20lDO2M5SMF7u4yR9ZGD7Exh1D4VMtdCJ0mWVJsU067uuCMS5lzxtWnua0TGYAhy
y5QhY1dSLUlCmZE23bEl83A9AFuBfxfONsnTe7piicL2nm/S9IsYqv4bezYRDJgA
Odtp+GxwRg+vwQdJfFCLHtaa7ZxfnjQ+rw0+DuDHmfhGIYqy3zSXMpzdLe+EdP1A
c0zU3cYc4VJh7szU2l+u1pdG3MmUVNnrhRFpAy29+aRHhRELvM8RrvKB/c8bbdIQ
wwIQC4d3/g+5jpXyOJlvvxH7Rdv6L8Dc7hOALF+WPKKSmD/F7bHVeGfY67W2k3OK
NGwOxXys7HMk2fCQPiNiNm6OJMG6iu4onzmDuljscf9gH+JOXm4Sunp0iRyve54C
B2lMwQDous3A1VqWvCsrm4PIik0rQ4/rCALmt3kAHzzoNzLQieOP4sv77rIqA6BJ
5Al+RlqD9TAqW9+KXZ3y6pA1nPVr7q4ptQP387soWysAaD0dziberR37phLans0I
iiFz9TDsjKck6YLhCcTNLroPeIcV9OuIYOXfDEnMBTmI5Qh+RYY4mcvbjvhR+zaH
owqEGKk3BU6IVi7K/YOpe3oNAj5AHdYd1JyZn55AVJ/lueMIiAyhUxfRKEV1IqyS
VY2SiXMMF6S/pKYlL7rKxihI3MVLwBolq6i0LeDKadAaps4ykJJqGjiSgYpFB9bW
k8i/jGYlIXg0UNyledyubeiwrJfziE1hvPOAAyn3P2Be+LmxqtEAdIPRcbkyxwB5
yb5jFOEZ041NoEvkQSnOQyx8bzPoeCJeGjNGoFw/52t2j9iH0ftUQrwroILvS8Ce
FuSd116AdRlmtXaK5YD9XgWIj7wZtHDOiJ9MlCCaxZUpHZ07SCLEM0/qG3zSiF3X
pRZ9XZ1uBwgJg78bV6Nt2MjH8ZD6V77I9Iak+46XCFGZ+vPrunoc/o/Cx9hKK08K
zuqhR6UAqusbeRbV6fkGKVypQpla0i68rYaRSl0gNq2hIDom0iDbscVbi3+ThlGm
6WNXeXfP7fPmhdG4HpOn74AN56QHzeV+nd3Q6gon/4qag4H3s1zYocxQ90w0C4Rc
IDZLRRqR6SKBG5iViixRoXQx8xifSMMAxT6DS6ZUTsmhA0qQH6YiRIEMKQwWeCi3
whR3iI0dwXGA4KQQ13xuMRnC3KokXBSYhV3i0DGajN/1jS+e+s2bQYH60h9rOPTP
RnwUEMjBXlOljnG1bz77fikxoPgkXiY21ZtHbD4wf1j7hhmDutybvcLk7WY+Ei/A
u3ZfcwBo7bdrh0HhWI9hEPDh+pSNJDC4rGEMM+Etd62bXL/QCLvHQsrnaDv0/cNY
vXNCDOqotgtlymNrC0DxNyj1FQ/yerPoM4mgYXPNCaloHWgG3U84ZW5GHosXzeul
J1PyoC6ObSoZExo44JsHxJ3YgfAKr8RdZvA8GVfacqBtysz0JiJBDx+xCjhVrIuc
FciGEXMuW9g4dU9jfRTXju8CbvCe/2aJ8cOKTP4QA5pKiX+VJRemnVuC5nVas90C
8e7HEA0ciQtGprGwzzVg3dcwcJgv1qVkM8wUbNlcoLN9OI99H3WCEVMLKoxS9aof
rsOI9Uqih4QWQBQDsIeBa28EaK9vycjOIx3oLnpI4X158a3GLbgEIGFrJfAEofo7
eRqXBYNv6C2GQNxH852XXkZ7aYn6cRCJAC8AHtbYjGP9bq+rghJmlvNXdqvyalj/
M7Y4fDdUxhxBncF/5Z4jyzttku2kh+5nh+mlPLISPRBSW7rys6oloh4kWOsEtaaF
58OPLSuwDbfyamXFPkVO9B69WHdtdG6+TaNPGCmTRRrCXVxgb+DWCgxwP85dQHc8
67QdXhA3pCza3QXUlB6BquZa0wi2Ch1EfL/u16k33881Q/FvXoNz52MMvThmf4nI
FRL/lBpwWyPtpVHqBsainArUCbEPZ2ZnUdYh1XDRjeGbS00JkueTYMMJD1pAhhk6
0UweEz6+2F2mafNyj/xyDYTtOVUclKCKFzAJF2eO8y/mifN2bLaqopO4q/HbLM1f
untCbRPSYqaTz7TcMnupJ290QlNWdFiPqjdLWB+k5+bKIYy16jgiHmUsxxOxk8ay
WUj2LMShVarouE9CbHWyweoyjb+QpPUKhkJhr9MwJNOB871Kjc3nGHbUTR9wJfNn
LcVqghdW3otJoXVcp6hPDWT1N+qc2fOL64IIViJ6BxOr6dBSGEUSIwF7X5aXrFQI
ODhbr+X8h34PwqTu0iG4Er+i/xMBw23GO4/dHtav618Yxx33r69Vpe8SqGykB9jT
7Cixq4dhIlW9rVAS6VIpN0CK/dRvxCjEbdshGhysW0YfR2QN99HjGnnlEkZi1M8j
bjGjGrEijymVoIBFcZqZDVbwcPc7ddSREk1MrxvUQU/IOTeVLpIqMZ6hnyv0TeGb
U+wxX571jO7Sstm8b+hI50zBfRm0vkH46jbooLBgmf/7O9cXtJ0gYauOgkRDvXSX
0/IiYRUejXPxwXie1I+6SepmcS4J6YRvuX/seXHxEyMbYkgjXS10/Bb+0S3yj/id
F19k/nsnfTDnIivkqNbUAPFcWGSb5bJHTO9cdbiqnJaWFXAEmGbN+jAWgEGaJ/h+
Oqrz/Cjq/fMnq+gugZV/tJiiyIH7vd081kS0onEdzNLkGpX21T9jY3HiSSvb/AoK
5fBpIGBvZLuJFLnK2Sj6qZdgdlx8KLUxOXDc6vV03iO0AxVaxuPkjnrl6cnkuDYB
5f8GFATdbCUXEwr6BTrd2Cdx6sVA/ufpzb+MtDGdrUhyaS3lVCTzhWbrrrGPtl/t
JlMcwHqFPWcCsq9yADhCZpJtAMqtDQvgDJu6YBF8r9NewcUSIz/CQSvNtTRtYden
wv3kbqcGjwQ+vnZ7Qu0wsjiz9aSMJBAnoiwQJrXqTvl60uJbXmQA3/YWopQFlsVo
YfwpeCOihASFn4S0q8QtvzjwCAs2sah6Mj1s99NImyKfBQj/3IrntgHNNmrxnDOJ
bCqdslxQ9w9Rvj42qSUOEzk/E4V4YpBf/7ukBesRkI75+ctr7GX8H+RqV7saxsHO
UmjAgNpV4tUXs0n/hQC2x83VbPfD+LLeYpxiKvMpMH0y71XFtxsI10oGJW/ewQxl
RTgPnfhkKlhShJZshOE/sMwga3loDyDJ+T3Jk6hB1Cz+QqEuvqHKyc+vzo+8wqrW
5vI01LVZv2GP7Yt6ho5Rvju29ssb6aAe68JjQOpiGjxHU+UWGGKJ04ZmrDrAf6f9
+Es4vxVzKbQh+Hz4wrw6JgtyyDKnOL4QjiivPJq0CSrcmDnYAF+HPSdYhQAcQU1k
fP0yJ5FknmY1VzZxBK0WMhu39F4HoGZhEzbmTlHoSF1tRcZ9MaLoRsDD9FWW0jCd
UCijI9Nf7LGcISvFxPl+qlLw3B7cw0fdvdHnO0/PrAW9RioluBuYD4zcIB2lV8SB
7ZNXXOvX9EuJPDyjllXrW1ug1JB1JWvGr/cVWSkzqCbgnnv6ueQe+A9pYxC3EKHL
y5huLupSxFAZbMnEjHGcRO1Qx5UwYsZw7LvVgvXo8oE/Svhxkpp3IX3NQwrM7hzk
NNlehUBOf9/LI04S5Hu2f6QRgb+xyKSmAWMoqMekju9vygyWXGqFdoAE2AoQ03jU
zTydSkn81cFkCef7E6VY4yWMtteLvtOr/Xq7IfsUtnFtmvxBtDrbfq1dMEJaJEke
m8Oyb+wPvwQG6WEaFrCFrwY1mFmYrFnnCs8BYTQiswzzZ13BczreqoACxJ2RZqy7
ifu4U928fZzwkMqa7plItA0fz15JxLGBhl5EViwjFIfnlr9JnywBmuEyJ/QEjw4V
fJYj/p2EeVrJn6RU0SM+kC7QB++EFTjs8GNVQ9G6j4yq653N/8CZZQMVlJRXoAHl
jjVthImCmMmQQ0kbTv8rtGm8anbHkHcmqsG/UisO6RUra+XFZ+BXYVparuHG7Gw2
QUz4lJCbuToPCZtkBe0NQpEINVN3qYjIf+J5iio5PrnQgjvB3xoUWuR1c6bFdgt3
fFvJO187RXPxkBTjArzehiR5ncBSJIPNh7pKwRHMiMWPWXN+CIAOGr18u2zDRHAj
Vk6uPJ72zWg/cJ6rJCpdL0/fm+AgGGgouf5sl8/7mRSS2c0Xdi33x3fCwIMF+HDv
aku3OyiunHlOO3aadfBaYrZrpNOdAWsoLJSEUwW2TGE0iR1/5Rb6VLnzMmMeHlsS
lzRgqazjVfRsNeD2dAETECBgJvMu0UFCZFvExzfNAkzoXGh+3v+irmF0VUG/tWmC
Nqhrq258MN0R11TEZQeCAdBE5bC2SSwflRA5wL11ENG44yDFFbxbkwvWJru4IRGf
qwSN2Xu/a275vM+tdaiefnbNRHNGQi+tSn/+wsofDdeeCw95c7IJKQieNXPhpqgC
HK6+Kfovg6YUfN9oZsXMXQsvZ2jGBBL30QD9PgB+p3jNIJ7Y5uiYkPo6Uz8yGjjI
X+wfZymWE2Vs7KkBwzlV2VJr8elZvOxPdFfQ3WGF586E5MCROakoezuR8TKv+oDx
XJ8hvV5bArUEZYyyfRULVmqBf9oQ6yziwJD2eVjLJy7zJ3OWEDxRJFz4Krj74kl1
73D9zJbvnLOCutGU6TKc3H7hM/XE3324I5NHjxesRjC/kFpzRt4Ra+YM8wxi+jtj
WmRqyTjd2T6HUJvEQZtdLZ2MOIpgv+Cg9PjRPMjsIxMB59JP0mDgpB+JJJYJ5Xmo
d/xdziPNTlEs3Ouym0pkJDVGOVsxluD7P2Hv4hgKYPjV8/0W+7GTiwiZqVD9l0bJ
Sp1Oh9LhpK6L2vPceUED+RgrlSomaa9EMCzAchECHYOaFsQcZqQSAlEs9wxItnrA
p+ka+gzPpO/DxV2TVkeo2LhaFa/e0Uep/C6VqpKk252CLylQ6HCap1nQFXTzgwyE
6hIGSp2BAcaP4jGG3bq0MDph77h3jfGAAKZlIEq20Sfl36ZFlMp4/1Cqe7QJJ+dk
8HMUzPDKQF+rqq8UZiSgEzSldD+KbEV6OaxpZO+Yqfpy0t/U+b6+EXgNnW1ZpqOk
yXOeqAoaP8DGAmE+ElLEqypHnS3KB3Nb7ley/gW5tA6ezqzXE86s2gAx+5zT8BTR
Ya9dj4WZoVoGyrVOrrXAZdFMQfifFrpsL/ep5QL7g87pp0vZeZ39aJQVnhsYA3oV
Dn9B+wvLbnMHEmwwyvcb597u1VufB81AFASiDzIfsbtDAxUT4LRoTjm8OjYW0bIP
M7wcE9RVvlbuW8s+oRO9MCKAnY2X3zYBKjiONCNj16/aOcThLvDIuPkcb6uP4Fq8
cZfEbDWl9svnaFFZ727bbZ0mGOBEY1rdt+a9KsdirqhvWYQhMhNd0x+LpR47vtW3
TNdsNm37be2oVCoejtYoUPCWi08dMrKKLNhxD7CAW78oYWHwJ4agqFCfyp/ucjiJ
cUwLEP4/xqI/q+EgDnv6WG5qW82qP8bfsqCyOo9Dx42ipKU8DzRaqOI8lxbXzhme
s7kG+lrrru/I1Rg4T+QM2gUylUOSDccRHRcbmKR+PH9dpH5xIby6l/OY6i+SFyWd
9gIUjQDktjtlkF/nwQ/b42ZG2mM4R2JD0wv34CI66YbYv/8IcK3KDRC504s4Xtcy
Jtx9oQdc8FbT7FnkhcduqQWFW8gegVJtJqZBdeTCpxepAzFF0ZmxuOU6uYLy104l
neyV652984z4GXPrsy/FusnBDuDP928X+E+r0KXI7ffeLsYynm3wgouWGaMHUamz
ZeIfoVGQ3CYeH+CXep6PwP+cbuXhrG7iIICjhOGxWm6q/RSwChPMiHrv2Dzw3mCk
9fOa59rESAMJ8KAWYOEAJt681FiA804fHBOTi37bmIZ4KQKamx832xG5XsjFSX4v
DGaUjQ1uBDhYE8bqaechGSs1qcoXTpRHAQP7sKbIrrQBwXVojUxl1WuOvF+Pgoo/
DfImE2xlaBFGvqt92vrC+xhYxJdqL5/l4g5ARQWj8B9/0ZXlZE6nimyN81gH40Qz
UDq+Wnl1scogCiBKgLKPH0d4WSm9mbdYXWUIERmvS2BFaB9KTy9Cp9YrkCqhfOCp
wnsttqi7wyp459v8aWj0Yj2pdw4fUB+WjYPIhX2WpeXsYiyegUia1w1bk3zw9nqQ
IjX0MLGvlAprz7to9y12LzvyUbTdxJuDgUO00n7q1PvuRV6RwUfPhE+mJdpgdJvB
pU4btc4U1vi+3600sIbXo6ou4ef2TaD4rFKdZLefzwfU5UJs8DfSdTDlpWhsoUQM
aT/6ekWM9ZVI/8cpLAiQCUVxd6zA5seD5gOCFcWaFpdjkhauVHf7WfTUKtvl8PgJ
SoPuObuhsnV5p2UqqDbJ5m2vMn5HTX/F8n9t8K8WpXeTyts1BsXvaAjSWo2q189Z
pT0Al5m2Y2XEswGInuziUypiiaPia6M46UB6sSKFnzhQE6oe9rc6sBHVxfyJgtlK
MCKSsFMeFrhnKvgZ2Dzwu94taWO5Ci8nHXhyETK3k76c58b43KhIQNscjpXiYoYU
hCRLFLmUT0chTqdmkslQ3XBneyvcZM9eADOf0CF6eIwkrhae74H44MeYuAwpLMAu
a2xTxyDoaKhwXseohKHf2Q2d04DCFjRB47+2SFNQMraRoLPDb0i8pxvBeqYLUfqu
m/WzbTiQXZjJTDMOMafUPIBDC8zW2pwtNXJNQg7qse4R/za41A+xs7r6uLbJHGkw
TqwcccIdUL+eUXpVIjnrI2GHCH1BFpprgGoT5hvFf8NqFws9M0pt/QbtdLlA8bsc
K66V5FEjOrddFDmPbQXIiXht3ll/2CZwiZ3fTzBEtHqW+qlXbPqoHr9TOW1GMki1
xHi9SznAc70tDldQkVa75YnKOHxVBrb90bGHvpdLHaSs3nWFEaeTjp1o6J0ARg/k
XY2B6pyReuoQSQmchIK9R9TeMPo4WyMnmBbcdcMeclA4vfQmBi5Ox8PWe9FimLjq
9yeNvouWUkkDZIsebCMS3DQqlMIXcMOb8mp/JxH1cZuDTvE0uMnY/hjnLvool+w0
/5UW8NLmlL2K4iSXYlJNIykKFK5VNPq7xUPI8YK4JSZk8xlY3bt3YVrVyDIfNwTo
XG7bfFk99JtVikjcLWnp3YdLGT4lwZhasBJ/lly1cH2QMdYf69W+YoCMCH2j+lcQ
mDezxvl7AVQOdVlDnyoae/rOLEg7GgqZZraWcklrEHAKZExZE32HZAoAuG8XvRlt
LLQmIpumJ6Hav68Y7h2V6NKV2VZdQ5s3QZ0fVT+1ADMT61fXzCgZjaDETpMrQAPM
7e1Ngl4ovsY1vRoPIlTjTCqBgAVq7WTt+mJ2BqVI7Kd4mFgEt9L0YYmchW2VWRgd
CSMgrOoTPXnwWlQIIAG8SrdxW3VEVNJNGdS/JsbvixjDQLV2YM72Rh4e0YfpyCMY
1IWrYZDzAxYNrebcEXmaqbwmJQVXvsRGEdrcsggkQoijZUJqVu2n2XO+tdBpH12+
zQoUud9NtQAUFd8p/RfxDwnLlSW5z63AszyQYcvUKjcY8dUL9ZUjPiFmmmpsG/cZ
h7Bh09CtMr5jSYHnRUH3oQudl8OTbDAvslKIMu10potWLPkrZl6udqa7aKyd7LoN
7Qm5ZUNttXd2HHa5oko4u3QYiGYxZjQKf5Sfuf087SMzKzFNpnL51szIJKerNeK0
zU3tJ8zv+Rfcb99FHwfcrPqkz28xKY6DhxlbziRj5qbyKfGzk6vdlY/PAWIa2m2Q
OPrEcMSRUnbxULZ7/fyes1BUbsHrpS70Ii+an4ifh/aQDZyQM38tzN55ro+7QqCo
xJce8F23JV2/Jg/76SQepCiyw03Edg+57Cx8W/0gJPy9SYPPVifH+SoqoS/xjDKa
t2l74YpGsEJlY/a7BHF48lVU0Mlfe0rmbjupZZERRsrNx2XIO5v6ekF4+LJ0YdaQ
jXRgqZsMWC10P55yc+RCi/3mDWb5EI2bpDK6apnGlCn3ijJZ0nNsr5A851AVC7Cj
pR0I5sHvMSCb0uGJ3+FpzOfieKOuV3tBzjMR/klVvX+DVany3lVSkuptCqCuUYoR
LurWWfk4z0mhDfMIsNCzI17wHA79wsYG1u53W1FLbMF1cpsn5q1doLskT5wP8Sgi
WRdWNNefdyT5BD9CqBvhVCf0RPzkl4Ratsg0+4PGLckx8mxYs61hW03SnOt15RNw
tkerNgK0sIXg4OYUnAXooSV0dxRJqnGqs/tU0OQa8cZANwWQsocjjH9rfHMhVTQY
IDv2o9Ss6rNP1b830lQmrdl8UNEGT2Zn5AoqNcAlO+8p+4buq3P9AOWRvdIbCNu2
tjdt6Ps20V39/rll/mze7ejfC/Ub8zVXZaM6Ai5tVIy1Eq1CaqbjILZYKpxvDYXt
8mUcHo2G4oU9Lb7GZeB/krZPHar9BtpBQJlAzLMW7HFuPcEB073GwPfiOTsaG76s
PiFYjL8ZhQChiCcJD8dsrkIDWxgk11a+WY5lhMIv2m7R4KhGe/gWEeXjhMXEvMPq
WKsiG+CVNEDpK+itlXs6lCvIGXUoY/adjJL8WnEKa1Mt2vWk5sLk7Vhj6q35+66T
FK+Jlkqn9mjfaGB/iUOVBCx7qP8AiiRO8Qoacy9RRUeqKkNvWeiiyDTb+DMJap8m
XtyZsbwMvvBZnDDzqirdhfGHbpsTn8raaYBAjTwXbIy6ymWQkL2TcrHgbNyKI3rf
pEDoAP4zdkQoQHIqDQr6hAC02KhQKfqbKYYALObilzxmJgeIGevSTwkT01Tjz3Xw
cdpCEL3Tv7jg2EPa8pfpyJqf3njwO91cJg5lk7H6PsofvDbh6vXpv43Vl6oAcRDX
MWYegFApIa/qhwsQ93KhXKo9DD06eI3u04EHjeN+bsN0pgpKywfvRCq/CaoC/6CM
Ss0JVuxqo+x6h+HfnzdNil0W1qHB7kTlmBcditPtAp6pBgnYLPCjvB/UZQnq2WpC
GFJ4BOrRfRgyJY5xDLOSIzQuQZam9dGerZJKxqixKjkmyUc91sZhUAfKeT2yCI9b
dHNssP1qfp6ICld4POzw6sX2mhZv9baSgo+uHUG11f/2SJLACnlpyDoN26jpb/4S
MppTbrg1dsX88aDXdKN9oNxGM/S0R07NEdfKOFk99LOQOjzhebMVxb6BqefPlh7o
5uALf10uzzjJ7JBgF8pFmon6dSzRIsjxNkGQESEojnVq3GyNyQEtXktHIYYyzrcY
WrPGkqlxhkMXyITFZzrtNYwRCpU4eQ4U0TV+/bkUpxOaQnepnP9YoMRfwRm07Sv8
IFzprTTMnbKmAuGKTimwFOvb/EQefAtyWKgp+V29Sr7Ff3xTAIB6n8IRuMXEv3nZ
T9fKzmo2LnizBCBo28hJ7fxFwUMLc3QDuV5C8PPAYbYWDG8YslIFYK0rf8Rn1nzB
D+p2w40lqxXY2pmqwFO8kBP3hiphs+T9pRDrPPKaTGeXO/35iNztCuzqMceHdDOb
heyoIcOMUEkJrkKFCXtgLbTd2JVCaX/lGFPHMA4D53uY8QBZfPSXHUDm5SKz2HEt
/9E4AQ3knDqhxrvsz31kX0YlJCjY/dRjnLYhjhfy0WLw6BXkxhoVrzfPShXKfahI
X2mmzGsEdhDl+9lkY94wd1Z2lkjiWv2cdbIoWk4n+o1n9FOx2dm+vBkXLDuLx5Wm
lwbZIRHY1rn/KDJUvdlqCZE4IH0Ijw2VZS7X9lwNHeosGPFjx8TEo1ipAUQ3j4bq
dsi/H0uBdW5Ntfytv9d9j9mImg290t2hWsuuyYzLXL4umvozlNT8yKnYdogu4nsy
KhC+3MBzux9G1WkbQEuo4bpWhntqvcCN/DPk49VuaHcZqbSUiPEZQH6nrKxv/cBQ
Ju20p8cMDtO8ruo9E/eMklx2MDeePjeB3lQqZm0zs3cpRESyoS8TmKkincG6eNbo
VJOiGyDpTYPBOl+GQVoNAm86sOz/DNSAEmVxo362OJVAs6mhtX8d7/jqkzBc0waJ
H85LFKMcclZ/ZOWGYU9mtssOpnJvrlNjaBEuwxi17H6vv3afcg5+afHVaNuejmUk
q2B4+PsUfRwjvKN5zPELODvdTErIlqi1lkoKqX4g352/PicAQi4Q/GcOeMf9+Jwd
nT9oC45p0/u7WtyscgH0MfmbvRfIvfs2ZfHgcVRgeBS6CwedLmbYAlotqu8h3obX
c61PUtUJo8RCWLfBNO62pFnPuAuUF2sPzzGpyP/xfOi07d36DLRnqr5CiWLtXNqJ
ogOZXM/ZUElJUvD6AFbrmonnD7BmvjNNJapMs+0da5NaNZbxaOsYi7GLr0SrYMf3
e/ZUgobD6Fgztc86e/X3uu16thmyTw7fW/GwdBQ92cNEN6ZQSrs6NsdP9MkrKynk
YzhssmwEW0P9czQh+7TbtX9Z1Yf6mJVNjgZytaUS2THFYy/KxdGjKTgJRjxTDij4
DV0TOMuI6Agr64lty26kfMP4wsjk7TCvJfDkvBxL6MrzAf6iCrK/uOimm6KnPWcV
Tj8zVRMwE1DTnHJMh4TGdlqrE9gAIt7cPKNJATOLUB3JH8z+zV6k1hMU5D7alHuN
4XTXYHwduyymHNcnpzJJDRM2lMmN26CZQJ5XDH69S55yn6HoneeIUEGKyS+xh/HA
a5zdqY//u/u4hEuHcLNngh21ndbQlDJz9fdELuFSxIYFqspMaAw59wEOpd3U89LK
26aj67GcOoHSvt89RPJ7rAvninI7A8meaRo/axGXSlVFEYsuLG3to7BJvflxMcIJ
is10w6pLIdnMseZcznPad9e9Gsc9rlszZk5/UwbIuJrgrNQRrsMuEWvdpbYehquo
UKiPqVuUxSuRAI407RIB8Gd02IuJjXQhnvNXqCZFGVh00Jei96Sti1AGNCnVtY83
4C7580yEjhB6b5mbV6HFs3e/p+NkOoH6RKhAYgdOkm/avspJxmjNKgTAK1FRCj6T
rqE2Ji6GIwOIYIw2aOsR/nwIGL2ucPVi4YKRDF3q9F8Fg0cWJG+GYuZCYcnzcM2C
iNPMYIAunP9GO+oov5DjN8+FSwtbJMT2dNhUQQokzyf5QsY+L7bKj8Xx+Tb6Hx/Y
VSZmzMr4I6WIIvSrRRUwFxMzjEt/ECHewuMVS8cOvaRT9OjY8iPRyMTmzBLH7S+7
CBWhTpOAE0PYFMV9duCkgnfTMbvFdp8wg8kCI7o2GCwh/ATeZH9c/K1Mv/nbRyZO
SdCG2n+Up2Q2eZhjkx3ystu93XP6iNwz/BtXHfutPPidDoElmKzMhy3ld0A6CFdQ
NI8YPZcMEc6DPajlYRnth9/2dINDNm5xE0VvY/AdNQcbOdl1O0mwXRVKuBSgL+7S
Bi4yse3Bxi4Q8po/SYHP1nXtRzVKislL6QeUU2/axrEmy3+gVfLh/KmMTRNoGQB2
FplEs0/gF1EBI8acG+mJ6yQtB2bc/ApvjXOP0wE0Zlm0o4LK4i6ncBiqFjc7p5hp
caQXX1Omg+jxuQovX4M9v6aqc73bWsNcZ7VGEfli037LL52Zs2yGSqORpQ+hqArm
N2PfRusLCVBw8NdmO4c0dYa2Nxa82TWInSuwNWzXHOje0FrojOaexXQKxR8lRgZB
Us/jqfBohvawMXPGHd89SgvHlx7/b4KcMxknYtsMtYmkLhEAf6Xf3Y/FZCQQ2CHk
Rrx/JOmZ43JLP+DAh+iHtn3hiFD/qqbRDouEsMVLb3B2haW3jajC2VTcZTlnFKNB
nvzaNz+EqOJCQEVDkpbK1Ep3S7c+nqslzsEigLWbZnAos+ioEL93kBs3I+NIxn4Q
JQEpVXgCyiygEXxvxUuY2NewxBO6SZQH3SMpIEYqT5XCnyC5qoWK/vciLdhRaCiL
4XPX6Wh4PLpUnO1RWPj1JjMd/+NQH0IRoEbZjPMobfM2nFN7WHMCaNX5Vkey0lVz
u+vPQs43VKEBAg0X+tihsD3NpQK/SJVB8Ed7xndzYC132vQ0Y19Pp1QDugFtaxll
xrfw2tbE5oz9k9NJnMzwlnU0SaLxyKHDovKBzPRd30TiO2WR3ON4hzqQciQweC2k
vzBoDwadWSeAUzH8G5IA74wub87Y3ClTL8sItZ+pM1ShJRn/gmo1XvtiAm7vjJah
6ItXYTG3vqCdQX8j5IE3AvQSjrZib8PYTBX9KZNWROggXhexeDebBFAL73CG/KW5
klT3o4q8raONFMFdtRtF6+2JtRelS/cR7QDs4xAZeXvetbQyP6iuujwqMPwxggF/
CzKuqntnM+XH+RYz0o1Xx+8aO9Qi991bLlukkE/LSPhBwATGN1M8Iy4teHqTn96W
aNMpqsQc1KsWgER2d02eMzYO5LJGjUYhSByZtj5D/QUGF55A4C8ubEjFjFfY2pLL
XpjIRGam1A15KhMWjGNxoW9qNmO57JRj60b02H90JSz3UQG9vzPF3Sj9Ly8gyBlH
4KyFXoDi8GIZ6YLN7uUNMXmcUHFaqxZ6QF1QP9+9tLCQd4pN7X+jNFljEawrOei4
xNa4qsX27Q0dm1P90UeLOgKCNqHQf0q5xmxHQ+qVY5NwTA+Vam0zvLRgemRHsw0L
QBgQQc3ekYwhAiaxinV7bKfaKAeZInZYDf+OEioDdWB4g+m2DwmKfJH6DAbsNjXI
w9kZA198w8GcU0DeobbLV0cYUfFqD9JZMiezimMEPxXWqgwVlKfKE0pjusZhF5f3
t3nLminYERxM+Iw9Fc+NEQXsdBZrCZu1tUjvbQX1qMBbDlEPVCfqAvTxzpnmmYdb
UltNUmOAPyceLUVPHqawOY0Pq+4fzNSml7eTNFRdp+Kxmb8pZDdVEPrlvWINeARP
YRbXm/q9Tw4ckMGIT0DbN5XQiRUHst1xElZEcrJURS9Qn5ZY302hNmSLLSfCsf48
dRqDiuYKezOmw/Gg+FJUKIE50T+pYzmBfJFJ98YIBontUgpgcbFGB5qUtOp0qihw
rFm+kpIhvOcR6NbBL80JXfquIZZok24+olPryKmqNY6eW3PFHT/CUbKRoVXMia7e
J2Vv6VCWBKsFeLEg3UXLqLBwjBFha9rV8Lfa6nbMKzS5IT49XTFX47Ys6lI36oD5
7aabHtk4aJR7xG61/ibstBDooxk3yiwRl778L6z2MKM6PWOqunYaixU268Lf2vyq
0+pCC16iBi1G2VrgWimWVAtA8aDw0fleoI3gQjrXjEUn7yp3J27Bp3m3JkfH9coR
3rhdePrwlyBO684oomCXZULk4GBnsoQZDP69TgEIRjW1i2MQzGpKD5i1VNoQRoYy
r4g77EXB3IbQwIPdaKuj8ae0L35d/QBE4YnVJPDYOsQuwiTITuuLLOXzAd19bG99
wWpj+6JOycU4D5JUimFIU8bZJkvkOHqUGP37DAdQeDdD4MLm4ZKa9IJAWrwz/NRY
C2wMoPlEmqQzw5vCGipEF8WIFmPbHxIm5WyuYHDflQikzBW+jubN4JHEMQw0+WUw
79ZAHJa9q5HX2PGSJ71czfQrqPLfmSRLH92lkiqroA+xtAH4Ria2ZjHBAL2Q57/H
QZj2nEnDQ92BDWN/0aDkz5hzmRdccYjv040VrBuqZ3gohIFCiLnwBqCyK1i/6XDP
DyNG1DjSdaJbuq10G+rR0gTbMkkO4G66G56NqBMY8LczWc6RZPS4ierfLWk7CuMb
4TGdMT5rVg/dZc8i6eoAHcfIUaGdQUKu8yVcbWvR71VwLyaqMkCGcBVT3hIPL0KV
2tpRLEAGvw/08JHHkS3KPfCuMSS0ZdcPFv3XfWhx26K8EV/DisMvjCDsajjf+c0y
KZLOx6ZhH2iqiOU2Aa/rHzQDkB6B8ymypigMvfxAcjrptHBjfqtlV3wmJhZJ1EJv
gnVk8ManPrLy14zkbWLNMvzvdSSo+kN5PH/CYM9xlZXGM2W25rAKljhIFIDqwvhp
9F2zfn0JG46BjFOJp4Bn4IFxC21BPcRXWqE08k0qk/z8lO0zeCkutarl/gV0G1Ep
bcrKUMYrP/Ae3vYimAYfKQTR1ayNTwWQwIAwvm5NQAPLmuA0v64zbISlhoI3q/yD
XwUngWccZMo56fCIrBMoe07SL9+47lPLSx85HQlrIgPTPoiHO8OTKOUhwR86vtJn
1lXEI4pidmRPghdUfm2EwjFDfZ0BvIh0SzXS9UJRqq+nSCvssIgJyFpVebe+R+X4
l6QORcZO3ZWEwUSZGEjANlkI6IH+XSDru4gftKwtkXvVBHNx0cAOBu2U5SpCnmO+
eDYTRHPtQAsntGcJ883EZCggRSb/7VIjhQKV0+ojlbKjDyy/K6gDG8kqIFSTTGoC
MBJaR3lq8rw4AksYtKV/k2IUfJkro+TU4E7Bj3XDvEoDg/ZdLJlygUU3V7NWAp//
wx50+E91uuUuRXXpPyG/BwkduS+/5au1TgHuT/cQHZ/hRPNrhglNAuhOtH6qmEcR
J/GOI0updDvPH8TH7nUEAtgGUnAhlqsjj+gUx3EvaTii5QgSUIpiDRqz+LqIpsj5
uhWe7biOtFj2x9jcHKLf2aP6IVIoehLokQmR0HEzEXDxuxdGD9rrkjLs4q2D116c
rtVYhMlPWuw0jGuFCuxsAMYJjH/qtFSH+by2FFBiBJR9BVsXQnFH/TjlWe4KyJVj
vQrHB+QHTpbMCdVkfU4I26WvmWCRLpbsJcP+VE1uexC8dCGf3WGni+ONze9lTeOA
VyBwOleTM0SLtwuL1/FCurb2xlRCljBAJBxpRb3IiRfmwoGmzRq61o4Wn88nCim8
gtnOZkms0BY7YFasge51HSuPP9WezthcK4A5tUoBcK+LC9xk5SfF8rhYPAuvdBHg
+go4hEiwFJIWszIIiIuXakY8u/1AYEkvDKtaYdopWYNNVVah1j6SblCYhwxyWS/i
M3bfPmuwtuaHdf7uvrmao+Fef0MMW6Wxfqif9XMA/xCHDMh3XOcwjaiyuA8/lkvp
WghxRPXSY0Z6QpIDjdQ9aKY4wG1T/nfMmEd3K7XYE9PyAIH7gY52oLBE9U/D6cGy
TNpcCyvyT84FDlOnwTfuzD4XbSlqYXJ0i68Xfi+EBU9I8W3tZgOGCLVa6y48TH2p
WUkiPaJbMUsLpDqpGpm2UlRqI6bSMfEKjXYKpBzu5SLMfU7GNY/9hyoxC8CgTPnv
BJm3gm5KS5iB38GvnvK0bq6GzXBPfb9LLNEZXr1gLsAwprPxpU5q4Pzq6V8u0n7a
zsMd1DNblRk1DzFAdiwEq7/5w6CgeR5np3kH+q7PZUBGEEpMZAMJtGRf687d5yBK
6CQLGIEoajbVeBb4T4g/lKxKRIEkIxCm3tM8D292jfMTrSF71HJsUQMmmmoccG93
WqtAcvD1e12eZe1z2Unm583aEwROBKl5gcj8aS0yjiN3R2PelIAm/S1dvanFdI7R
54/avp7mmi9YWAh/LlZ+kpm8OTplfETkJSAHB7I318nI5L4N8EyVJe9tVyRfRrB0
viq4uWXVXUKhN6FybI9a5+9y3QJbeGBw/69s2hY+1Ux+1kojT0t222Hq9CTZPfUZ
0Lyh63yBtPIMwtJWdYwSLq2ovjgHQa6B60xM2EtKvXUAYwxlOqFavXMxBBYyozH8
+BXRjTG0kxI0a3YmeeTlsyfrKsajqIGhzeilHcMvXlTYXrTNr2WJE60cCYX7SX4E
4VPlmAoh5BCfj609yFAMKzZLmZ6vZ6qFCZSKutzx7Ec0eAqsC+VVvgbBl0ZpzSi1
a+b1f0DViQGxBQ7MRewavu4lQSbRwTqaYml8ls/D/Biw1hT1ThJlSdbxqhmh3ddU
d8OKvDrQ26ibSxqbQfCSwn7EX6gi68yXl9SL5+UsMSxD00dLhg7J2Iw5Ddoz40Bv
eYNPSXaRR8kG/RWHF+MC0Fi+CCzx7n85/6/k4se13tMUIoOxOgq/asTapcHVzAY3
G4KuwZHwtBRsQ5k6wgUHTZXxt0gN4CFKMQ0WOqrx7XQGj0WTxerVtRjje2To80c0
Av5mx/gM6OaeirHLoeRAUm+8Efp3BYwJTSsK+FRUqsDlx/MbX1FB+X01Wi4Z3A74
Fc6oLvxLr9VYnomVGTgiL3xjMwwtsGbf+7jmStfcmeHD81Y4JRzXd33wHU8QHV6e
XZ2q1744rzkz7zO3ZQI5Tjj5i6/Ee3VkBihCVYr60roWaxks98nNtwO/IWLJbJwb
Y9kwY0TxKDmai6MBEKItO1SaCd43TJ8o0DXyG/oL6oSRJWe00oF+sYTDmiFhmb0T
VzDVhDOIC6T0R8zRyU2wamqFjRLvsJkt1H+kTsOTWgV7a5a4yPsblp1miaTGkSXF
aOaCCt+lCBFeyPFxM6wWbOq+Ccnn6Yg77nNHNzHa1wyPVgdkXLuHHyfNG6l85nqc
X09n5EGHEVnWHBQxMxdB1ERmsfdLVoxJwLMJWmeJTMTo/8MT6KSZhDythyVuqawk
QEA+kAENhhso1lQrC6xQOOZctK+bT4dJYhe5VTiamEv20z08CrnQXFAA+8aXYIx1
ijI8nM5u1Or2M6LowMMOVo1WojpUvok9RC5u+Wh2dmx82LbTi2ao5d8qnGT6pS7P
1ONFJIxmaEisc+goRVZKJe5AIfXVTd1Qjk9yfcrcjsFMnDPC89IerowC+pun1nE4
7L/7Nrafd1mLvRI8r25LwcFfLTu2V5NdtGUP/cbcX5WcjZD+djhPPGzFZIGdhc++
sqdcf5bQH/IN9vWq96l2V09zcVWPmweKrSg/ntx5ZD6z2oMYKbHiH+qokuswNs+n
ZMwrGGkS7o0s43Wdxmqp5Bv7q0Gol/QDn1DEqczAJBTlEHUuIIZus2iuQpzfWNvq
2vp3CRBVcnPFglS0myrzXPe7VRGZ6ZKRvCFymt3oBCgy7eRmtFn1uL2KIVCNgqwh
ypJdaw1KMd42w3ptiPfTRyUcyNtW0vZewAO++JKjdQXCRXUNeCZufA4sPYn69vaT
u6JbiXK+Np0+VzfMlJiUex9+D5PAVIMPhVdRE5dyYGR9nAPNYa8cIlxd5pQN6hrE
8JT5Wf0vu/D8Tp/91Sss36S2jX5284RZCYsSdSwBJ/M71nPpZDJTJJqjbndtIngj
fbWag3a5VfYNTBcmErlLMvHYShIpNcWJYPhO5aIWg5eXy6zh5z6zImA1xNTzSUVy
CZJBJXEJt4KiuOnRynLucpyfbffX2hDIfeAMdfOgrXPT8L0tiLyI4A6tZc6zAEv/
j+ho+7y6d55piUwWkGoP3wGNYOZwoI+nw6C3apS3ouPQMg+pnLF02N7JyXa22Wv7
xRGnT0EzX6igXeH0ss4ZtryfhORQlK0HGoeTE7Y5AHmtbTWCwgyFlhHqlBZwOoS6
axyBAOhWQor2PnDPf+MtGl0VrsfDaBwI2a6SK9G3+W1eDMNCpgGfoOYi9i1jHUyB
2U4zn0zchOaQVOuNZ/2QRL2isI8yv7b2DSnTJVSjcYoSt7ivbH/DFZosIz6zll95
08q6fTQUY8T5MQWsRzvuksurUI1iadSVNvkKclCosRBiMGcyIA8TGXQreftbdb/i
zjF4HN1qZ/cUfKbwFZLCglgudLIcZbv/jC8huWJsJjd3CWcyURLfkwWhMTIHp0HY
MLMgXNLQtwldmTRn46rG+Xarht487ravgblI0RWBdQi0R9KIjaBt7e6LRp/1zmlg
dIuMiJ8z/sqwLCy3HsuEuLLiLLgv1TLnNJN4Zgpfw73ekyvpq840+NtLrLeCuhHA
7sngjoenOM31GKcfAY7C+yXoS/cdwWHWuDsb0SJ76qlizBqB5zaIoW6g8rZoCGWE
XeG/d545gxy4SG4EAhsURwB5OxNTUUGlA9TXWLq9A340gfQoRiT1vQDwhyDKeajW
n6tNUSKhKA5IROVVBp//eBkbUz0VMkSonWwzhblKDZ8POcHbhGFZOjlpYJYHyzeT
QDs2VGO/rybY6tOac1fPCaY7hBL0Dk8I/7Vi+9CuUiUg6NzYIuRWSSlnn6kMYvPN
j+QNJdnxw4Nbjw0aNERHmW+UXYjPKH8R9VrJZsysIS1dlL/dzuZQwcgTAmGsN+xC
ClfXTnF0nkOmKbYtpte6KiY4aKY40zcZtcRQOmFP60qUrYClKO1jtjxTP/QgDkeb
UsWti2nfPDDFub9OceYRKOmoplfikWl1Scz3pnYe9IbqmrJBH01qhw+Lr212U5Lu
yQAZxpn50XtXbw8OPQezJ/KGq/dtkNrTA53ZafM5NNBB5AvRNAf8hOT3W4o1jFRt
AL6P5Cvle6+0Y/AT4qo+Kkq3R2ZVxrzp2zcZpu0oEsFH0XxPdv9ox/nolfLiyGYb
gnCHsfpKhPHXjTMaIi06gSu/ggGzJoKhmmKlZ7zymMxQoX0bEzbIo9aSuEz8Y6kC
FNEvZxdSr1/Ylr+u4onZWJuki6JnbWZZm/emvfqv75m8jl+g2xRKJfrHbaWIMR7q
PqDaL7sembnMP/moXWQKO/N/JMnYrGLTeR73vyNtEQkq01aGiCQ0tVNQyFi8oX3b
eoOCffVqB2HOf3xmYN1otzvY/iuciVNW+Hhw0LCYaK+Lnf4ZShyq4d54o+UcVDjV
GwL7A5cV/hWkA0T97gxzPHufDIklmz7XpxW+WfqE28IzFjlanKFx42oNXa0mIptL
YDpR3rCXol/BIWCCGBNkLChYFcSpXgUYZQV20RBCgYR9JP2BkmjjAvG8+d+HkFOb
rWbxYmJQ9CuEWK7XZzcsDFNXSyDTwzGis/CuCibQN2LX25BG0jE0lRaQ6ahUES+B
ASGox27cyFk6BA9n+ThSNa/TJ/vLLwGexF0ePagi+TLKS7M2HCrfnJ5pol/rj+PZ
DmPUDyVqeEvygCfaCnzd/zFWxRepXS/pK9FCQhFVuhWLiWnRbtO0/ilB1ARQZcYe
a5/xUK3LgbqWZq2rT68NtgThA3PVPr17vXuVG9Dn9h13V2/F6vrjrRW6xd/37vP0
HF/vKx6HBzqKJL5tjdKD90VZjVrtX6SCdRA/L1NJryocMtWiXeTOmyzK2EVPomIT
W6jGDFo5xNFJ7auJWExOg9j7bvHegUaGEfNUtuKTXzMIpEQsFgYawDQTWkmGIpYL
UdST1bw4OkXEVzQvmWafkGZKUelP9TZBb9XwQAoifHWDaO2RTCCjGTPA+rhCkBDS
6BxvcWL1CQdbmca5kK4iqGQcENJfUw5B4jixD/kQk+MBrbsEqy3A5piWDprbgCeP
8b5Er4g8xa8olzx0P4uud41S0vDdQkFn5hO715JpjaVgS9UDT+zjRwhrYfCuswJ5
OhZppigLaw35Iystaetqahao8UiGwPeiBZ0GeGcySydfbq3YrsKnwwJMBJPC8anY
eoHAayIZEsbEvJcOW/cmno0VFLQJ+VhS7Zt5xMqqt9Do2pBEYVXmWH7B0ZdwsyEz
vBm6XQ2Ib/rnIRDJPq6BJJOkma1OpFMmLlSFj8N+sbkC+G3Qq3iCfygu7PR0+oJ2
7YrT2XA7WKJQoCglYKcw3qbt9rDy8tyFuTl+jFx/h/KAysv5jsYd0Slof+livAhj
YJiGY6Pr0OqItCWtJmEYZtA39ejDSbEbSS7sYdJfaVCd+uxlb+ewWpQoqJMbTnS2
fU/hu34aelSHrHlMJdCNY/0rPrg04HNafWnCP0VBV/ymRRTVsRKl0kzBZUKj5OAU
KuGbsNQl+GXxeiZhpa84DLPoUIr/ZE6NMdQkPMklFj3FU3G70G412ieCiq62TkRL
RygA2lusFLeB1FlLY5cdPsSzkZdFpa7XpmYwBKNJ+0MhfDK3ZiXu5xhxg9JsCD5C
ogsXp0KgzQy5HEzd/NeKQIXn52OVq6/yGgnaf0P98gQgbbJLdSIPm0mB9jdg0zFs
xjWoe9kKq3FZBE+t74B4OZZSKSXOO8jq/i53cqitIxZmDzZyIASQrxtcw9jlEmIv
wvgNOHLoZXwBCkn2b637OwEIhpBctyV1huXzBAivvkT0RgmiruHkzLc/gX/C8YTs
Sgoz0Ph9ams9g1ruH31VNUmGxLUwBx5ogL2/qR0zQ8+x1sw57XoLhKyvw3HBxEN4
sgYZsez+7y0/eXnUoKyfe5KHfjHY6Vj/CR5ykk7od4yvTIFL+sxNmKNU5JzY1s+s
oL/riFn91X1jRfmsFA4+i2fG47qyY4LtIFUolZTf9/802KUgHoq57GEj4y6aT9qd
WGOM4+5kSg5Aqox5EHzqh5uBjSpy42pppMtM3extejG5JH1v/L39c36pTECkT+Di
FOyduDQLgh2W0aYwqnOZO8w7rIdKgj8pqbhk0etrojId6Fp7BB/WPkES7ZT+LJJM
ctoA3uRriFnr0TsyeVQE7zTOU6fcKmUHJt//gBaN+dGw9rca12Tq8iI7pGgJnt2F
SmYu9Nh2bGSBnGxaPJ1coym3gEQE/jHMZiBiJ/qIlLr68XLtk3vmIfE4skvtxOzx
+eV5c8npPFnvoWVDfIJXk6rMohTAnb+3dKO7CkHBhxiUxhp/DvcnhdyeJla2ALbm
YU5B67HFgnCq3sv6VZVduLBVLd7VKAg10mPUgxtQpTv0JAeV9He7wDKLrBImKPWI
lI87JcIlyvWw1R/rnuGHUx2J9QZJQ+FVCFSB3DJtW5/dcEzPDbi7aLBqaZX5u7+x
COET9KEf+3f2/FlwyzMHiLtasO40Avic2PVtJLRdnUZbhjwthsAyXDnw+XRtd0MO
XLdCd5otvho6jnyC8o+fDzicWfq9NbtyPXte7EWKM+4pBjavI3HNweEkyHfhysa9
Qj3OS9YkYnL+9+bXjuZnX0/wtfNMReAC1E+ae48mALii9dqNEa3tjekeYAf2SL+Y
U0FJGWOa0F19grX9D48Sy2/qvgN8FGAfzkKr8Y/qEXY/+epcJB/TNk/fKpwLuVvm
5nGkvdT/LHcHrXKnSaR/9xNKqWJkVNKiPTo4rvV9T9awGBVXm1R5aMKPv0xVESbP
3/G5CULnNxs4hyYF2JqhTvGiAPhtp0ylEuPLriseVVH7ytO75X0Ud2E3SXZJ83uB
2J3QdcKDCVW3zkVqpeHPthS5EDVL4pbcdYuGPBJcSX0cacURiGbrnM6KrBk9/HC/
uNgdZmt1ioK+f44v7v5DqrW052QVssKgGPCbkKwg86zMZ67nQD7z6zSec9kJZjLz
06eO/Jiuv0gMxKME2oX0DhYeb2uff/IDgvqdGKc/PELoEhC6BvrACyWqEP8k77Of
XQ4AhLh53vTuoFn7Nr2+xRIF/V5duWgGC7gaTt4O6s35FXKdtXn73ZwDTAj2+Nsr
fC8t0r3G0QGnVuUC/t0tFmEudyn6doKthdA+4SAr0B8j51If0GSJJhnZJ9fA3XpL
R7+m41p7WvT492JrXtfPSQ4FAA57oRIntm75C/RdcpmmNLmNmz7wmQNgzJ4bFvpx
u6vxmTYAeXY2xde2mY1F6lBg7KphDsz2cJl7Kzy99dD1qfN0Zfd6Jr9KB3QmfJz5
43Cqi0s6GvUxwd48f3o40vkFqKOGGxtvDFRDXcUTUj6tb6kXoswJzRnVGDutwwej
fXviEsAKnCZXgFnWSkeyPXcAZ4fRa8fu9a475u074vWURynE/zTqCwPQAHBOdxUN
469BQOUkD9KZ5rTggnHsaO3sl8aEnIguyQ/FAKbxdhtQK+GCBtcuctJtGIzwQkZV
kXTmFAKDjitG/OxDByPzcNn0bHKGYc4yiAMmGjxbCGGoqGktlBZOmPHsO4nw+PrN
cAdfwLAUwksMpNmJSEk7IOQ9yD/sErxHQFemYkXWKH0gRmi08PDqFMIScBsYkBVS
d6UUkSdH6per+Pqaoi1H8hD+mw1DhP+Y0hLosWsNn+qt0znYbN7+TzeDXd4xbKFM
zauIzsyyDqY0cVUib6leixYSHuV9FlKQwfKWUrIabyPEw6we28N92BEYwfTfKzC4
Tt+PPEICgGQ3BI3fJylj1g94FMDsdNhC9fNebR0swiNGKlwg851k2S3/WsGpzyow
ES6/H3VUZPLYYfLDTSe5l0Ev6tbMeN/0SizoTjwP+Ag1PunsPBx371Di6EzJChNO
FYJvYQTzbY8/YTsxAgitD7lyoQ+CPEw3BX+zdT9+thF4Duht3GfOJiRD9KHyF7Dd
RhyBC5JWkrPU3owTZrLVBpjW1S7TnAkaH6J9x1dvVR/+yG0a5B9MGOmWWVLQuWol
ry8aviVWlI7XrL7YD2V1DBYKseDj12/LgiME7aoEBs6lkp+bsrC1PM7kJfaC4ifN
IlDWQ3CbH/tqZULS6XymbaJ6tvrJQF/H8S4BK2K/W07lerZA/L8/fdTNO/yNnFYb
lRGd0K5TtiwYvJ3a6/WGEfgXgnDvUHFJkjDbB3iWJk9Ls2jNYWHPFZRKtzVP7SL6
2MhFhlt9185xeVi3iMIWvamjmGCGNzrRpUir5zFcM8GE39eSPhsnItDSzQFX3CQa
oza49xhJXVyb5MDlcUjzoSzORmx395j9gxJDocYZ7oWs1hbzeBwQlxS4xSttmY7v
+Oi1TNsS5NbMokRRAxQVaBpxjch98leB8HVokV10c8NXLirXpr9kesQG+fXwC6FS
Hu3KXGg8w+3B+5W1z3uRowL8X6asUAGCm117Ml9tGYzRBYnj0/a8ZPQf+LFBM2Vo
cANE9HSMebdPoz1PMOLNWmF4YJkyhwrtFKTQl1Ur4tOJyLodV0AmGVwCDZRHXi97
veyR7t8Ktj6LWtIZ0cAker7lNYBHewcivV/xb9+SDscBZAUnDj5b6boFez/PSXEZ
yRNg7j9da8KoJwbAUg34/a4zx2cGxJokvoNS8vf3zKQXOUYNWrE6E6Oh693xiZfp
y7GJEqG6yG8GLglOYJdpRWUT6cFUX9LOkRCZrNGuq/yDR5HxFt/j0vZwQD/YFsyh
GM5p2AqSEkZr9w71NNOKo9KrmNcX4T4Az9YgNdR45DHpigJR7tOnfbuM9eItP3AQ
ZnPMa+uPDax/OqMmODPwAEhdNyJ8Hr6UCC4jeuaEHtTPPLeoo9qOUIp48K1YfxgK
V2PlqJ2X0Y3Vn9nZJ68N+Y1UPVYcFPEczeg0qneDEBHRGD2IUxyS5WPX3vMATu6G
ZPy/Gs6hhK7cqH0iXOCGWPLjYpAPxJz/rwguV6BS/tTphhUHL3gBPocAS8+ZNZUo
9lGPuHVWQ7tDUZ4gl604l29DHt+DlTSYOA4oFPT1u5YSAeHFfpgmint3qgHhGCQe
rVQb6x0nPzVgGTV8oPNcDZhECw/RCUHaV8vsuDZ1IOE1QSmLeDhHtRVtmEEliRTt
pkceZGMUmXuOtfWZQoKkNe14w3+U8Q7l3czgY9DrtHNIQ1Z01fmKd4k5b7eVQIhw
0uxQm1YOCON5hqHh8qJQiQIJj9vlIUAHxk2BJAWY44qWCDERSdYE+DS4qx9R2fHl
YHR8qj6+V5QOgSQsJB23MZ/dQjid0W1sWScbuvtWYtJTrU3Ky/1L1xgmv08xRFHy
uLFjpsBvqfHIfhFpL2jgsq5dcQvmKr++oh0Apjg3rKO46AtC7IzhnQDpxAiFUHlV
hjhMJnyNnD65Sq2GzicxBEWKrGHWnvrTKbmVuMLECxRJ30+mZknQJuYQUxycvNy8
pSQlyDa5p2YdnDj6ITF8FdWeI72pWJbdJ+fkwYIbwQmfA3LogR0ihuHjurR1Rb52
zR9chHkheC2xuzTuT/GNfswDJXf3z7fXjjg1PsDD4Pd/Gwscd3KMp5TPdIrDDs2W
XQrnawhDAMlrcesx3ens8O4LtdjUvugX6Lyr7R5zvQpS6ClAlxU5cR6cfbuILNeP
wSF7moSNHIVBU6e4Ppqtu5s7mn91upQaabCYmSYdI+ZWbIVwIgF41STiNsCnivHT
UawQ61nC2iHWxWjswpFNkUDI47hmieI8GfiZ7xDe099xJBBApqf/vk94eKVLTyIp
byRo7/shtaIA4lKHX/q7/ddvGi7Ex3yd2Je66Jhni+kq84jsn4q7XFwKtm4wDyOD
SpL4y0eKWBxT4rfGKXGB5LfTlQgrrV14OHcSCyvlkaXXWdt34k6gGeLvxOYdA0lu
ePVfF2t7ZDofg/15Cjxuj6beZ4D3ZCujT18zLHmS/bQowPPk1NVlA3XDZzV2M5JB
LZ5ns3XqGClY3A3fWEXHrYrzaAZEtq8uvYsQkb5H+KozNM6WxttJ5mdoHgihfsoE
EZ5AteprskxQilxLEkf78evQ+MKbMZ6dpQMWth9b5NMBpguDMqNFSeXPYpfz4vfL
+z/xx/JLV5rbQAD8StICtoUuEWs2UsSoBIsdKqd6SaA2UfghdZ8MyCwKaSuOPGXL
/V7bX45AAKqJZPrNd5O0UsayaXWv5KAzCB2d0SMGq2MdVZVlajoxAXeN9G3/4gxf
ECR2n/KtIut5qO7G+3DyIe7wCgCNznA246XmWYugxRvq9INzcywO2/DEwqYCj3VV
6CqvNVg2IquOYQmIoEYy3YifHayAiTDyz1yZ23wI1ASdVf+6mWNIJOyagOmpS1Sm
Uyzq6aAZ5sKTYF78GwDUqfGPy3znj/bD2XdnzOyHk+gHsdl1gwCjwusUJ4oF8tFw
wA0h3yLm0Eabn8ZxjO01kZuFimtf9zVIs6CCLBQzJi8Hq9n2lTyaHGaFyJ7tGMPU
hFkIjvDXte3J4W7RFr0ftzIxc481yFjw1lQT3/86fwuT1M5IN6wgEHTaYijfXQvy
6H3FFpbJ3MhGS7ky7ztJLr/Eo1yZuvZKhpqyGgigYGexrCnN3f/p4/xTh7LoXKb5
6vf2G4B6p64U3FYYzqwc+r2bWvE3hkL22u73+tOrkx82rb7D8egT9tu4UmMBktwz
UXYgTfo+ZF141CrN+5IQBlA/snFwGGBdoWYLJM35lKCWn9HuRqKoB/FjX8u7l3nK
ajCXWY5IPMiCSXMUE3lcBSw291L/cBgSUfjVd+TdwEoIhk/U/vafuUl1H1MQO246
s8qPk9KLtFPKI3YIQC9t5H+x7/ad6dfJ4unrFhWU2+tmuSiyXl7fWRw1t8k9pnJY
cYFUUdeY2YsRSEvE4HywdrfuRM906fWGaRMMifO/crQ0ny1MuhIQBVD6TJZIElc0
QCIxw7vHKPe22annyBwtes/XiQoadgTi+9scucRG/mRk5MN1BaxrKAZEuD8YtA/V
sUcVyqKHGaOS7AMq/M+nnr69LNdzw2S6JkfGjBI+bvR7l62dRf9dstZnSqoYSdub
J+85OjHNIwxfUCk3j3JhCQ3zF8NJQdW8nJIPbY2tHN2UHzbY3XZMDgmuALyhyj1s
bXCl2q0yJfVoNAFG7CLMvd1VPfvtAJATUnu6Ln8x+w66+xDSzmlFYCHPXpH7z+UG
1HV2u9Wq5XiHmbd8UT13XuHHtEz4O9KKj5joRBgyNKiXGkQ0Y/zB+gMgWqtePa1b
nMph9lBbyJTRrS/U5BHCV4hEU7gMAs5f437qaQ1n6NhT3s8KWkcDbGH1HUEJZeZW
baVUdmt/K+NBhDduZZjP1iRk7/9T5qobY+hCg9Nd3vefJE/Oqw5iBX3RUeSB6Nf1
oVS3Ojyo2/0REEIdqLaKRvJFq4tZ9D8M8swvop5MOE6KfeulpOWh7JMG1+3sxiKw
Yh4WqppD4IZFWEJ9ABsGMlyRS5y7s1b/IHlQJOwdyvp9X/1RrFkxgAa1GzLfTFTx
H/VWwzHQKlWCN1fZmlASWHRO2PR7OpqaT0I4/rBac2GE1H4WcHhdkwBiT0KU+8Qq
cT8J9EJpIHuKBTgZJhk3n1jDVmKqwNh6ELyUmiTf6zHrcHPJMpYss4ekASe4fufy
QnXLlWiwmRtS6AKelAJQd4hXRo0E/eVkSZKuGU6GW/Zy4L7903DJN37NPT5OE+Da
ts8lR1Ghj9zHuCheJ6eRSQaEm8FRMncwMyvK9YiD2oLZpXDMuMkzc26EWq+ntZ1l
LS0sgtKDBaXg1OS+tlUdcWKiM8Il4vTwEf/F/7V5jjB0YsvFPx8Y3M1CVOAP5Tf9
Bl3VYHcIXsz3jt1ekrHR47qotvXbk9TqINe5zO1lzME9pdTPvpF+6JnJiGf4UeeB
UOagVORw8bHHJ8y7qPMrPdb5o5BxsyK7FXn0k4zVwTLAvAKpNh4ojhW7F0eI8zhN
JBLJYMIKTmLRzJV7JQs29cizQD77p1vJVIkxT+DtI4WUWCcKfrWzYrSkbeO90Aw0
wgWT2Q8tG1a9eObnTUEZkn3spYX3JrvFNGDciglL9XezP/OJonlDge/LdpGku3HW
KtDYflFiSWR0PpyWpZVUBxOkkgjiSigqOn4SpKYwMYGS/QG5+BiCmo1xZ51f0a7y
cQgIx2UvM6m9ADOGhx7G3bC7gJ1h+vgHdOOMLgLjUrY8XgV5TCbjbGZa2n0oZwUc
iVNOE09Fpd6YFNmjR6ycQ0T/4xVSkEFWkypp0hqBjOmf1q+i0AByp5BCusAQmlGw
0TilKwSncmOG95Hmmma93mQllEr48QigCNsEalHVmSQogd6FA4jj9oboskbXqXIS
iSOyH8L/RMyIk7KyVTQZzuVhidH3iDB2K9xeMdhE7WOLIqwoLKPE4G25RNam+99v
ZGjOBOwaJCjap6RoQB9ff4jEN/R4nygBpMp8ILOttAVqngLBx3+u+k7OoJ/vVp3s
qyFMGD65UNWNqipksDdaWyPR1C4nYJvu+H5HK8iv2IvdN1F4vVehN4DiMRwspJfq
9jJ1/4/m3bqplVrLFbHwEUw17nWhnUim81Q3LE1AneMIO6SKfLDrploi/5t8v5ay
snuMeieXZUG86MD/BNxzaYktViL37BJivvCTok1akbCUUb/OzLHgZGWhyQhOaaoQ
/wXQ547vBH4cUKGIQMoLbDHK1Szg93Q15ofJNvz+i3tY5DMDPDHMG51pB5LQW8v5
fFLamBaqjyePejdsIyKIEUW5u76gef2ukV/RRdrjhu0Fzr2wpSwzSOlaSrsMpKvL
mcmla58wdnwK+pQhczjqtF/1hvEJjXlMDEv/mE5nuY1/GKPuE3zBZZF5qmngeaTj
PAzTKC4FoGCRnhqTSQAQWx2bPvly2KpI1/QPTjcErh8Tf0sn5yYO5LvVe83eoPVE
KB6kXMM7z6hDXgr2t8GvrIAwocRLZ87lI+oTc1Bn+Sm2ao/UrXqNP2tHa8ooE4nF
jTY2JUuCjwLWzwTHJq0YkgdRexHzJvGUgQxqau/PSawLuzJ8kNV9YkXB9enb0REz
Ali1AnOweM0nkKNKe8y6C0MDV+B3ycan0vFXYGopy/Mns3LwduRRHDuu3pSX1LMv
0qiDgJH8JcxD8iHXpnOjmMhvDYZK18LWCdwEB+RuIkRyJPsnMu5QbV1VOZIgOk/p
dVTIxXDyLRVtwywVCTzuU5tw2Y3dSEXCHU2uQOVgORk/RUT4QPEV7sTDA2ZvSP6A
tpzJQ4CaWqhMONohXr+opCOitjjPY7dTshRFmrHAHY6Ume5wA8mgk1A+VIpH6CMW
E6LZkVVS5Hu8eTjj4HpYKY+UGSicGTvMnh5wXOvXy5Zf/iP91FejYaIpsHdWzZvs
J+rMM0Y55OaKyo/2UwPvTtRfzrpV8MICoIrcO1xQKjmdCRA2GmM/kv3mZvjLXHQ3
u+UN1+f6wplxI0nmppQCkGjaUS3QmCiutU7fzd0SS0JQnLMq7qn1s6umHRndPWX1
qg8sFwrfsHSMiPLdV2zcr68zUgxuGFGotud6SyWC17CXcyfu3tWiD3JCYUqGrFlC
EP39RssSl/igsb/zQ1YIgSU/mGjyMO3k6K86XVeItfOSM6rn1d9aMVNbrsgp7ssk
9OV7EE5BG0NxS8L1FG5XGO8ZTXQ7myC8ULodBrliJqu5aBqXP1Yi7bsRXlcfJWxp
vMVghfi5yzrlNoZYDEvkVVl6tMPy/rztpSC9ltsSfCKsZzybbwfWdL46O9PmWn+l
fbVo9YdNZ+BhCStVBf/MjxbPBsR3i2b6Elp8xIibztMHT9e6GZlNNFSUEYJhS7YZ
OuhZqkACx8eMpGYXDlGMf/DjFnfSy31H01m2DMzicHhJpPJ495yiDcpwQHmR/TCI
esy+0YZoUwu6FFLCRmpuU5comr2HI+p5NP2vFlCzioZGEBQzICbqm4baw/xF61PL
xQ8vKSeoI+0uYv4PO+PDatsIj6KgdSRBgxBXJLP9FMt1dkUbPfxAFANT46JOhCGA
xEYpJXzr04V9YCbjE2S4DIE+2Pzfm7aQwsAX0wpLfsuSA4kekqmg5xo6VTojzpcy
3aIditSbSNMPzI7Kcshkk9cqo8eXzwhmvh2vwt7Ho5g5bInSEQi+Lfe+uTZK4ATn
5ZmfZRcgZLdvBmGUEMI62yxm8W0XWZVbsQA3mZykW9FUGyNc67O1ZkNe4QH+J4tV
uIpyeEf8B1krsu+v71680AYL2eAQ/2KoouGl3f0KhmFOfgAtv4OqZMJopVTAU/fZ
y9zSDshOpQi+tGxuMo6BvymY2ANiD/KmphWoCSnpDe1DaHgLNCCDywyLlxVnhhvS
sHBSGKqNuRgsDesVrYwQp2d+LptWQTPmeTb295CPf3QctVrJbFrhvZJc+MVCG0/n
a3InVirpIbvUx0rU5PzygqNy00VaVXDwH7ZD4t/Vis8U+x/3ITuCCsu2amHym7vL
hgdFPKrvwq0DleIe5Sw1PawaDBs6XqyPtEQ0sZPJukH8Dx7FBQRK4m8+Rs9bvwNp
sKCH14eZB8qtPn0VAhJkAuI4ZYk/3jdEeJ/6gth35+aRordopVfA04xWK6L4Ts4A
Eg2srxl0GOknD1fahKM0m9nJU28ZvNflD+4feKOqr9yZbSE3EZ8D8yQQSJSuY4mJ
+z+vdmpr3DNgtV38u5vuVVo8A/Z8SmZjAZxm7zaK7U4i0j3ay8IiLH9ww1duy/j4
H08FgSky4WiV0hVyHSqRlYruPP/BbthSPFdTrFbRD9u+2zQ66OzSSDfXo14K2XNj
Cw58M25w0NTtLtkQvTFJt45MKbu/aqrgoLeOpdpM8AUcQWst7RjohkFtLPoS0NBN
MbIY6BVytPGUIfgRiq/KeX+ENyF/XM3Uxh4Was3Y4oYxXFhdwp0R3lyUs9cVO0xy
8CYPfL1BvvUcDNbRopRIJwb+ZmmUA8Mce6IuhCbrwupxHe4hi6FcQ/jEIS7n/tn6
HUEtCrMJBj70+7nWY0/D2u1tAKnG/WvAL2v2QXsLTxtc2Zt1YnhOEjx5OY9o8o82
1hqpBvizILUybGpzLJUVb8LYpwBPpITa2YYu4R4F+jnwEDgTOBwuahuL4Xyz1Xrp
qYM/XX01PDUdQsGtdqunJCHwbHYB6BoAoOmG45VjtaZyjn1LPIWIDqoMdhKX5weS
Alwp/AT6+Atccby+hTh0l4Au01fr3Bo9ZDtrlvvnnzPzAVThmGEJ4gwhVZhD14lm
9ennkrUsqj8iLG7AI6Y4mVoptcwH38njbtKO0V7ExHD9vdoFr5Yi1/6YL0xdKzt1
2002o/4wYptNPGGDIGJ9Y0ZLqxJUL07L3MzkAbtj9XUx+4LreYCoY7ZXlk/+GCaB
UUs4s+fyfWMsirMSim70yaMUAgO713GeJHhSQhwukZdcCD6xuFVDEuQbjhxo4gDZ
Ob8tf8QzfBUZ2Fm0txF17p/k10D6IBnx5OKphCDjUG0M7wQtgNat0tx34hp/12UR
aYxhu8g38CHkmVzDKo/b7J+9fLMoFG0a1bGEaCeAeiRm4u5XtMujYlOaS6nlKpZv
XYK4WSPDvQIdEMrTIdFRsKW91k4YXdZCc7mN20xXaeTnTXt6bFD72QqmLlPY5lnM
v9v+IiEsfpyRua8yEh4YwBETOhxh03W535adMOEy6rGRDLbNBgyZ+EMMr1AkYcSE
HmUMS09Ad22YtHwwqsO0x1tBjwuovD1hnJKuyZ7YtoNHDWl3PZQA56cq0MoH0IXh
b8dbqi05RH505FJm/CauqPM0/i3kCYu25B7oDXNmh31W6F5BtTtGkLclIF0Do5Yp
syyR5mLf1VfV0cr85YeSluYOz+L390mY8bYaBw3Lqzfl/dpzOLOoWAZiJHuBBgaV
AmDDtVVfTCy2UMe3qPF9hJ7GtLDlQGdQAPEmeCVJVOrWaMR8HxDcCEruxzQDmjL9
yKF1VjJOibx2Imo3JPp+lM9YsbeRPByw/w0ahkfghM9LTx4oViYhJ5s/bxsm7o+l
ZlLI7gKhsbeM++T0FlIiuPy+qT86FN0p0LMKH7UgLXfEo2chyxx2lzTbFtkp514c
WFVBRcp87SBEHjXYX2Acs+oLpwBEfL+HDHeMtvQpfigzbd7FvT5cm9bSNFKtDzjA
7QA/C6yTezwky5xXo7C+l/UuUvZVs6QYXjE1l9RpRtoabX2ZYDxjOQhgmwtcETSP
1/C3KWjFuTBTdtCSLvJJ+y+nE+GbEpKPUzYzZBcFv0VTG0LJA3ctuFNbPnQzLy/6
UvUsr7PfisgEzedqWKZ6CZTlqEzxwa4A/uafMsIf4z89R+ztxxwC5o7D+mrOvA/H
yj88OKvqAgkzaGKqhWuq1NO2hjcwgEJNDaW/qscVvA9jFNCRYMQlzhiyexpbnVPi
Jt8/IMszvcazMT32QBlrygM5nvPSuPOwZNW3K9mxDNhZY/wJ5oMefIbk1eaXHt9Z
1DXgc3wBPZ4JR26IjIriV7NiSC1D82/a+tGvRIQREcwNGdR/18VkIT/ngwbyhToG
RszIOZrWWe0pqB8lyUlAVJ4Ufy16fSFqGxmVv9LTf9iuwnIgyR86i2CAeatY+FA/
dtQh6bEu/tDt29c4h0h7LMbo1M76CHiyCLdvnlXyVYoL1S/42LXkDxfWxsyz/VGh
yJNvFAnUcA9THIrtr5cu17rPnmvCX7tp3bPrErLIO5NmQKvtLKSRBcEeCU5kUEJK
kbwtTYtEy4ePy6o2nYcGjXfkah/n0CEuM7fkDFXu6Yxbv+iGUthxztfjmVDIoT8d
BCrBChXp3EldxTHK0D+TLbonyGBvVQ9pV2o6lb+/4v9UT4sFMsQh+ZSrYVb4pIJJ
nShHlvJoXDiIq+QPq8qzQuHItvkhdermOV8C3Nz1wXy5ZtzKiSwQBOhPGNFVZMe6
G4cVSgUTR4qHXXdGrb8djwrFghSqESW1DeMS4/xfQOPnqs2U+uwDrhpn/sDGnouV
pBrEjM023I1tDr0f7AsucySRX+deqQ7zTvhZDbSgsxMZAd4PFUqzsoMz4/SLq0BL
Zr21JMoYB+Teo+P2E7SyTCKkmZR9m1KjIFlz6EuyZQqVWYhscdlOZlUxRT5DBxPb
8q4+A+TUHJVWbOgvmfRIqvxI9CCy+NCvZdeuLKfqrvcSf1doxup+AN29ycDJ2rLh
jyPB/m1cRk92TNQd6y6UmJoyaFP6Hf+wFCVZQgHTdgf1PTe7VuCDEbMCL7eylUCD
xvm0qOU5sTZ/fRxTjf6tMd6/vWhN5HQkaxqq/95gjaXHRZVCLhgCGZbAIcYytH9B
+vxgoswRZawF90G9GMzGy5UHc2k9FhP7nJ7QGgfWnjz3F/BEE8Sy0TgSKhP29yZB
ey4Qj5VIU0rMFpj49yedQYpYYPdsIjwyuuwpT7blGhiuKhoQIb665sQy8OjMLar6
inyXnpgQb9NBwnmtOpn23/lC215UDOlExTrwECXyDB0Ws5QUWGdpwBedEo/9ATfS
UYPKn1FDv9wb4JZQg+T2Fn74jUk0TZm64WOvHcZzrf3Iw+CcigfUNhTj/TK8uLEv
URcotLdVGiIAXaSo/fkXNHV4ia7U8Z69GJ5pTAYVEv704Dj9B0nQbxJjSnkotvXv
6tE53GDYtozWwuIxEt8p4xVl27CDd2v7lm7oYjj/4PRxLTPxTOme0jrM/CfYRgJg
qZFipMYnZceEDBs9KZVeO/UQBf6byu4PVF4L3vM/9INmHSZNCzlUEMSIv19wu4Wl
s6u8C71VRkZIaubYMCX3doyc6SY5U6lifMjPS4wgaSwBV/4Fr+D/f/JIN6vqQh1L
qe3Hvv7yrXCqykQqWY6AkOqQUmAvt3rExUF1lXgPkIe6fvaB83PToTznwkidJXkh
FMtSQL6pzv7x/q6PIe2ce51jM/SY5EhuyUJbcGimEo6+FIrCIWmsoH1nPCOCH0az
J745K88FR4Falb3ipsGMvFpbOy+f/iRraX9DxMBWh0IpMrRwYOGL3/kcg5ylmdKV
PGY/2Nr+YqSD4PD6FD2ZSSh4awgG4B/doFlNDdpOoGxbu3ZZGoPx1nRFA5Sw9ZUd
gxnIvzqr0u/M2nK1NyK0Qguwb5Kz9wm88db8ruGLep1lHASkmJQ8/7WzNvNU1V86
THpPNsoTamxLpY3bHpkVC/vs+FtDtspUhWvgtM6guGXlz1JpgHks2sKN80EsPuca
Kyi5DnXcPjcJORY+N+O8dTt1Gw82rSU74wTlHqJsX/6mBN4awpKgs2jOCMIeB225
7lukdpzoONDI3SEDYPlRfEGfud8qLcw0jg2vzKkIJaxdvpuW0LohdycUfZjKyiv7
J52TOJ361HXVIu3hiofjT2yu6cQqN8RURNzJLbY8tyhTwqZa1ui9shwy7C3Tbg/N
bKROKTefcSoAtz1UKHhb534euuq0izUKvNjQXkylTs0xl4mZBaIYgKeLAfgKj7XR
6rj4/F7ENWnlXFKnu4ZbDuYxH05FoU3GozRiDVP5bRlPtUf/1u2eUDWdmRM21Ycf
Ww6j7yKkQKVxwk24Mme6NuFl7ccslXMHgbTKWvix7HwrB4V7VSzQLgx7qYiG5PfY
DNiwoJNhFGjZsDOhDv1JtP5bKNXijyVnfkQverZ3a19aon//Ld6n9SB45zEvLksB
zxtsnVi2/3/tYWzkeKONUkRBVFPsWy1Gxuyk9WcyG6pRxeQZ0346mWm+hn81gC2i
BL3wCfQDC/stt6EfvGYpp5Ik/p4YSV+CuwXUF4j4XCqsNZ94BDYui3vG4Xundokx
rBZcagiwchM/bA4kjOKuQXMPrhiukb19L/ufSP2e2zg4zqPw6OWktHc4axDARY8u
ZXo/L4kD1MF9NfgMsJZz4HBxySzHj13jtE+7NGUjJOhgb4BDDCYo3Y3WqJIjfFzV
4unEJIdmAUyc1leTO0gld6NiO3OwDD1PpLqs6EHylI3s5h0zsTkB/P/RYqDB1mwC
ysErmDpspEVFeQMls5QYfQjkgGnpxl+v8yznvI3RUlFWahPxiVu5iMxoQ3EW3grb
gm4pLqEh6O6rxVd39VM4dUOGgXbsBLwF6XrNL5tEaRI5e3Man3efK5Sv46G9yyPR
imy6z+jHg+G1XVvpeTOkvpchK/unleLHTtP6tLup/Op8/Rcc5cJzyWjWAraIUaJj
PdE4IEisXmUKzMnjxsyELriE3Nxp8H6gt95znjpLyAsZUeahDc5RF4tku1hkk1aa
6Ht9hCrg7jqs0mSm7uV/2sAG10cKgxi7gAsMj1l/Q9RRJ7B7F8tIQByLsbfBi3Q4
hUM+bVHIWglOMB6mijepCR8aCC7j87+YDqVM9rGYO8oL+IdvhfM3vVDge1UX1lG5
/PA9utlAHF0icYYlB31puw35HTTp6Rbzui6dk+ZpShJ9a/gdr6h3el2MebAASEZz
v1hCe4nms9mzEaQeLOse5/klyvWHJ4Loz4za+ENTnipmBpcb9RVCBDU+64VNGx7m
5I7RuMIt9emhlY5ueyAX8lVFtkk1imOkEEwvJU9XIm382ot+ZWdktReoypdCoPq2
zQbpI/pQVwpLG0DGXMqHLCR+F2OfHH1g/V3/DRJXWtMoHNe8eKipQJFCardlH5Kx
UFtDLVz9U/3OG3b0/dxhoWUXATe6qRV8SSeTbqUNHavl5MOcMtpdMKEzGMo9UCot
AIN02x5LtoHrB9z8QSScPqFGLnDxzGr848ccX8ycFYcF1w3DqfC9IkJ+9CQ+1FSX
3xgRQm2MLpyezB/4JHG1jDJ6SGvn/2+zkd8pcPsGf2Jok+pE+0wVpTlIaPDeO8Bk
SvU5zdo63HDAsJjGxBzzDWH76gFWNfTz9KD6g88O/QbABt1rmvNa+EgOxDnJL4R0
sCJW5FsBrpIZp6o/Yp+5j1/sL3gPlQV9GBcUi9ZYBNLsmR4/RrxY03XCsTLkiRbG
kjG4JX/jJ1qLMQidpiR93dyE+IltWziqAg/F74xFDIIhSXagGkhc/DaVvbD6Obet
7ll+CwoMUcBxKjB7yv9NWN6Zw3voBTQ+mNfJ6hQLQSopiIZp7gWL3d56yMHnFYxJ
nhVlgP0BZc8/ifVhQoMtG9WRLzf4fLAN9QD1dmsZxGfZ0LkdRoyrJ1iL8llPgna1
5voD3wsEF24NuFsZOLLx7KHiIssHzrnxMw7K9bDtbARBW33SpUnWIKUFKzSTsEvk
Zt+HpjACn/XgMpjr7jmmcgAV+js5iyzYtWXwcPUkZd5TqfgBens2mQJeUE52cP0S
IxcC0dfzK7DP0LDt6MZVpuyZMTJrAszocrVUYjzyXbBxwudnNp0MbUkovxpFbGE8
PexBwjuhuplE/EuAgLRuHUV3Xn3woWy/EPPSdqkyoOui1ad6DCrEwEJo/9RBfe53
EkSMGDPS7aYEX6gBLJpJ3QrprBl/JlqWTyZiSn0o7tMSW+XC7K2dV2nvA+Z8Tgve
bhAzci7L1JaFGfuB9/CT2AI6e7BTO0Xbz2QyHB+YTK7JFiGFRL73IoeInbLRN5Vr
2wUyb9FyRxG0w1ekM368mslNygxfHd+few+cnPMgV+VjZAYfdZfyEhKi0A8YXW2S
LLyGoZlr7oPkw9ammukeFbTMM8+OgNjz930nqLbBa5WF3l175VtGK8bKRYdS1tDB
cYZLoH0r+BHKpCiQ4Ue4qi2KU1tm8uCzdOaoj+b7wXIznlZpxbHZ9iv2FxhRBInk
1LXBwPMVl5I4d5LO2WviqzekdK6Ez/3v3zAoPBM9/eWulESyKr4g6dFD+pdIRU3H
J8sJ82R8xVzMvE9x/qTbCnO2nM5ZVOtFyHNXrbgpBo0cDWxYoqsNjxQ+is3qLklH
Xl1nss11HMtkYy+FqIcuuj3pQbj6WalCXEGZ4iTg7PCdoqEhfpNtly8B36JANtFe
EeNDhPf+2Hkgdf98kZKM4ppcoHojE1J3o/UxsxDl1cYEKgpQQ6P2ru082eK4vMSD
fyC8GzfGfV7CxEipYCbdYZZj7Zk6k94e/FEOYOTMjeO0M/d5/qS/0QdmejdckP9a
ybTlkyLUqCnWlWfkn9S3eQpP7Te6MRuaCSkvCJ/eWMApNOWLisOW+Pl1Nz6XS6/W
77Rd+uoVpFxTlvwOhq7lsBlLlP4ru/L2jIjTteQo1h74zGwQystB+7Wco0GVvqub
hV1X+gnO8yJCXqOt7sQ0h+EOOF8FCUOJVafYSXI30Xo33M1iOzmBZNoqxLUjBmAj
6s/VgXLv4807/EifU/xa0lNYa59wVcKzkUFEUjmNXHEqmXvvEBvLrjkjKB0p5ral
oivyVZO1aoK2wKcWDWVam0Mu6eJGou+aMBEby+InTL29Z0qLe8vzhgJwXx8WMa7U
H7Uty2jAPlKLVLszWSLrSJsbrr0Iwz0Q/qKPvPYu2e5ISLKLTqRGMCv5FaMj4W1T
H49K/2aVqxj43aSlWW4Fwo48uf6XP+OqKBXb5vaoNbQmbde1iam4N/icxH9DDGGE
8D4aaANSRvRl78k/EGN5KB77bv7xXBtDvb2Y+2J48w/2VV1GLBSRpREm8ZB/wWPC
qG2sqTWK9rTp+K+c2tv5iajH+lNgIBbRcSLRU5FUTRAtydmnvJH74PaEeNOgX4Pv
w+jjo3zjI9W0YRLieIk7Lm7ykRz15IFgQwwQmTOfGGEU2jtkBunjzW0d7IVKJKaK
8Gt8WAhvgosDRfRKk5BZadtv2EdebcqVELCiHi79iu2EMG1GQ6fS4KG1rVqWzs8p
sehdmANhuFq3EAn6mQOY2CDlEqHSL6IG5mO8Pez+4TEnZ1EZi3s29ym2i188HNYz
x0m7rO9n4+nztTDZ0HpPpkh76RVdSqqdDxsTcvlb7641MLHQDfVV7Wp/JDO/l9CX
V2cd16d5Q/BNjyEqzyDjfApSxmqvVrwtMdo++MgTGqk9kdj+QUhhdl0AzVhwrAa0
81LoTX63ka2dvJOktKwVrD1TJclgcqf7nMPhui+c4hGuwFGMyCcWHhQr5LlfgCni
HF08bkscYDgVhxBAfo/X3jF50VOYO5VbISj/Y1ty+x+1FebgzJ8q67Gh/pDM/CMq
A2Ux1t4X7kLTmTP+LErpNHWFWzkoO9cyOBmo24dh/pJtP/BN9Oj+GIg1bNaTbXHW
eTO55Frus2V0JRChgKeP7rFl9AwF+vCy67qhSgd7v3MPeMoMH1D41pU7HznDINNC
BNK9aZgTOF/o9SfFTfgAqVQnFoFgzv9KISLThQakwqAGzKVrN8KRKdL6+Yqf8BYm
DBrVsXxqUCGxePejml+BZdWlriN7Io+Zp/4NM1jUW1SskX5amBtPeu/7s98aOJuC
elC5Ele9v6GaaD2rGUc4cID1IKTKKVgfp7mnRUKVRyeQPCDLPnt5iaf4QklmyO0l
Xuqik+qrBfwFf3YBTsx1wUwcEwQs/kqqOtyMDYhibwEVsQt4xjp5YRY76KXxytf6
ftyyFhbxWWzNA/tXwRWqHLjwTFYPahCBix2T8DRJiv5h2oaHUEbcQJlIlVW1jQKf
R68NaP+IFX0W4vryY2lWZ4H0HNJbx3yRMnrhYbpwCi8JJWjzUXEgGRCuLKc20ISC
806FiHf0cDrAmXavIO6W5EA2VKi0y3bpcAz8NJ+uf8eAjrt3FJtKtZiV7ToSHFYz
UeUa6Vhd40Fo5kRr94bOEuBatCMWECNuLG+/Bfnpcmw3syFIvf/t1CZnZ5IRoMey
ZG3/98W+K1L6giGxy0+dHtrT0Yn8Pv7LdrEt8o342sybXXFOPN+SpNjufaM5jh4v
56w2D+n20Q8SfxC44jv3pjI3eKN8+rw/5CnNe2gbcEbegXeKnbHSYKLdATJ76x9j
9O8poh162/NXAzuPvG7BIApqNTuOi6wzqvOPtlsp+RdpAReVKqxgsQ4DtOh0ezo1
dP8c+Ll3TP/lvfhNMJsyEFf7NTdnINBFRw3PK1unKicWbEWP5gtHCNVii/BMboAH
f1X8sj6HsOVO6RZg5Cvc6do7R3H5KhWoYskpVHPwkzAqlU8b/M/qRLbADKMDJ6av
jrbnIZG04u8uvpxc6C8rZv0Tb270k7pZMh03y9z5WJrYrvTX0uO1tLkwarAg0/JT
AVtj09254USnNDW7LxITKuqaQjSa1X70kswZ76Qst8Wp0dJ9iYQcgU9T0g6uE8Ry
HgjUQ+IHVkTbW2T5wifVAFbgv4fPtTTHUEPSZ5lB5/FnU5rduHkUkVBtEbbPv3z1
/ItB3qMnOusyUts7Z8lh8OCq9MenEODQ+Mlk5t6s+w16gfvNB7h0q6AIW6aDJzR5
MRt+pKJo8c4Rac9lKvawsvx742YWqOY3ZeMBcNcydftCeGThbdI5HVQ8UdvHrmJl
Njv4qBYorKfvVXlcQY0c30mrVUj1f+SL3vtkHqkn/OaemT0UKevBZ7inn4BjbtBI
u9bqoX18mGZixQI2Aa8MgM47rP/fpYvGgu1mRHdPkV6q1emKXoTpHE+0nhKosmhg
M0VTG0E91YKLwBSVclwE/To7GF+jWfnCzH9tYYYdjxshjl4cnmaIAay0mIq0iVKW
stwiXKO0Z5kE/8BABd/RdNioIj/DT7p2M30ZCugxJlZpFVzQytesRyOAuKCeGMm1
4uKLVi4ryZBhGbEe7TsV1Wy9NKND6T6oHwwv6R7ORVUdky/gnxsnSCuaxf8pwxWU
SmlZQnNt1Q5ijvnX+uJi5J6+tN0SKaedVACE0bqznX5myoxfxAuEQOLH6r1lVWMs
z/L73GuacnysJ2L3nTjXcC2BD7mlbXMPcePQUenG5uHrxw1lFUJHMyAFLYiWlYSc
L8ZOcJFD5/2KFm4eTmw6prHDYWEwrhVs5xPGbAZHBFqu2AGeS0Bzq7IYmz4LTgUI
D32mlLLK6V/rg6U9A1YbYnyw4G9z22ozOEdXVtB4Qj8EGuBktCbhLwkK5KitvbOq
aD4Ddq7qoGqnNthuk7+jSoK2EDSyv5jOnXnD4Zbr9fbW8YpsXgf+Zi7Mk0Eu/cPR
amI7OYeKLajLqWbD6ZUE1FmlmUrhoGsU4q1J6eRND/pv8DTAQRjCgIx1zhNr88CF
psNaZ6920d9Cd6j9+4zi3I4GvTM0qCeUE52dqsWCJhWG/cdytGcjRuDoFnWLjX3w
npsKq2Cdk0GfdGjVj7hSciitrlpG+ffhuNAwwbWdBlavj4VX1zB8CIRJLLMYdOOK
bUcZMawWFAB5rQEHuAJhgCMgcNZjCR7Wrg0zjFDI0UR33k3CXXqRtfPpWEQlDk3h
1RjeDDdgw5G9Hy6rmqtXeM5J26vldYaOZZ73KAImpOiscZFbdaXkCympnB5VJSNH
WpsHwwfALWGoJihjXF5O1n9+gM/1iJBmMRMl2gftjkEtmg1JxberPFoIgxKwUuFm
c5KLz98ugcQC35lE3NA2FLuQxsqUN4aUllZS2QYf+xuUMK9aTSUsUJFUOHr4yEnI
M3D2EFfKDVVSgDNuo4YgXJbkO/ZpCc9SgCmms8bvJryhJXCxLC2A6dPBzDOm3N3i
Q22V9ScHHkLmSfmXQ+PUSjmWm9k1brRMyHYiSw0cTcd3zQ6MyBLmxbBxYgC/KPMU
dAI6T0QWWZg1FqCmg6jD1z86USrYtXZxeRMP0SzqqW8WaMHWcUe3120qSgT2O2Y7
DVuc4VT77An81tVKx2b1wXNx9Y2bbhW1cwe98CZTEQ55jy4syxDqx9c3V/Fist1h
x+u3hxbF2a9dVteGlJ6MnFAe/VMjefwxuTvQqtfqqGZmoxK8ZWjkyLgtylrpO8Vy
SqYrixIOnIZO7/N46dojlF/QTs//1xmXDppQ8fvksFnqSqa1HQa0ZJ52yOwWCCDy
lifFpenc/Ex5sZEQnhmNZGcPRaNQwDX02i95c0O1RtNl07DvzEWucyz5aLtu8732
ME1mscuCQST+4a17SgE4b69FTNBvOTZIfWDu9SxPw6nuRqFkNJwoglXgxBuE6nGw
rpOxERHmrylnGn+/A+GB7wEciUCZP1RO4NsGyuOQaq2Wx9haJZYv+4hKysx3D6Kn
iMqFzoGVYQsMdOiftgci7ax9BxiGwl6l+ti8WMgnP3dFzoOil16bNU4YiRWVEV0t
kn1AKNG+l4GZ0rFwfKfPnsmyjHa3iHMTR3xpocW3ikp2ixwbAIYZ+Xvmf5K6odSB
9/dxHuz36kxaPkugTaLcvGDygSDZGiMtTMua2hVgkDraj45cUCz1/mUbS+26p65Z
/dpFSP8lS8CqjMVanj4Aj7/7ybwBQF48thtghXr/2zIr5tl2RzldpiRzfrba+sJQ
EeMhpqehFqeMvEABq87Z62bBmqj1We0if4XPgQl/V8VAxCKX7XG4U+DNrXzk6oYW
PSE2kgiKT10CNPNcRwd2UnZMEGw5/y6Q8bU4JcugxXjLEk22HQ9zCixkPiBCvxFI
re5XUCHVc/+LhL8uceeagnyCXuj2bdqtc8eU5i8ZY5p4Frb1UY8Au0Nakpn5Tjo7
T8sIWRYCmpu2aBzJBbEFBW2NRDlOD/Th5A1dv2qvMIWush/8bmjv/a1Wtgphb0rs
li5WpN5+tHXu9Fpf6pT0qQQcvV878Ut+drgmYA55LF4knAvGWzN9YeOoSbw5l6yj
CIaZxHCoECsdbJfrrjGBvEq7uOG5PxV6HG5y/93L2+4TPR2wc1Cbv8uJyUMmPxeN
hVou/fsUKALUVTz/wrXVfOUelRmxP5DcMVu6bCu3vhpCimmbO2W38n/098QS/cG/
Qr2Uy4u3gUigbR9ptbRUdnBHTx1tqQweZjvumfmiu79Z1ZVX5rq27/uBeFdOIblH
LYjv/EPeMoHgbCpkXMEr2vB/FvvYvwwqabOZ0soZgB9tbVdOQFH/UID0HQS5PKgQ
rG5FrF2p0vBSibACLekHUfjZWc5W47cf8TaqdiKlDBq5fo2tkZ3Ze7LrnqBP8pk7
tL5TeFvCgMRC0RxzMwEWqS0BScKmTcv+oCaxmvRCCZWMvjwoalJI+fbgKoo7i4Vz
U77apNyQVV5t2z7BLLjGYTVhqgQ1vUO1KXHv+GNaYqIkvspE/oiM+GSxI38p7EI+
DBzLNl6r8u35xZ5/Vh5YUugA9RJNQTPO12WfQkxGttG6lS2HJiFSGk76QQ4n7g5s
yw94XdXq5MN94XU2yiyc5bWywVfswGpjOVfpLYd1CVVORukY/bTbrFpVw9Tr+Knj
IdkoSVaLklWwUR7XniMtVp7vJoapwTe5m+fYsU6SL/DplI4YGw6kwqDBCfqb+33j
deegpU7Y7A2HgazTESqLqP6gD/hXzh9gmPDQUrXNwpG13nYDESGLFtKsgj1fQh6h
o3XUpZ63z7HLc/NVQhHZ4GE014ynRcTpfiMmErVBXBBGke8HUJstoZruEnPX2Uv1
35cYS9Bd94fic1f8UabcJz15Z663/0MmWQoeRReI/1MxzFtBINKaz6tAd8W9Kuh4
epdspZnp5DBoAxbLZkTTKQhGlILuZRrxsZNjAA3bSBW5U+R92Wc74AlI9ERh3oee
60NqaKlPxc+Qw6u4mUAiKakR3jW8td3yCxCBHX3Ke5NlFw0DohLZS7ryIJSFpflO
UMDpzg6cvzECQDAjTsitqhAJnwuEUETRIUcfAfM4M2eOxerJGxs6ln3G4m0OLoXj
ZKJ0oOHV7fDpzBW+9lVYZC6PHGujdKdLc8Cg+Fi4B+ShNmTC6jdlQ+xiuVx4RkxC
1hMb2/oODcm42Mp2uanAanAFe0qWllnI2Khrts/qvNr1Fg3JeJiNUJ3P4szuywQA
nrK+40ElBmitwnVzSV3dUCbYLuasu9xtuUxDiaAWqxGtUBHKdTPz+57iweXjsyPz
ykVkMqeZcxcyw3LOgMgH/FkVeSgCvNBgvdCXZqZZGq7ziy1QryrAkBMGnHUwkdmm
zDS7J9Mkm0cTMIzi5wK9kBzVYTYJvcsCQJhICEHGnvF+awhnx+agMYkeuaoXdhEc
V5VSZQoDIkIKhCI2RK26/n9A6pYnM7/lIr0rmQfTK0WDc0t07cwzFszyk8zqmfIJ
U3KYDuXPtvZBpNsySdlGPLpsVL06+qWTV3CzB4YhMs6UzCYvRAdxqo9Z4sgbVrCJ
RrMwmB8wAMh4mIFiSftgYcKRFzKBfunJMvX36YaRB7Hwj32oWNo1lVWSRpCBEoOg
aSKI4Mrk74eSZd2gQFfH6SDtDDObuBK7XNjovNNqzWntx+6v/rM7SrEw5YYmN2Hd
qh0qDILdBporRweWQ7yPna+2H8X9drABQ3gkGeD6dI5ekfgAdcexzPfPnRFpfZh9
1OQgjXnS6WJ2ATfSYb9ut4bYdrq+BnMS5i7qMSa3agTEvKTyLnQXCFvxx9WNsebE
v7EoB729zDwWBY12u4St77IQMl5OGjBjdFbFFnxnSwVBAd/93q3itDPi/BHCGryX
Ahz2TjrmdWiyBLAmThRmAxvygOmGtiIwU9KedzGMIwgZVF9ZCHdUMrkYBa6oe6hd
a0WL1sWYilLGUWDrjawJs5JpG/KN0QDxASAHd49fsv8ep4dwUzxexRYqfVXaioVJ
z9XzdKfFCehUtwW8bb9rSfADH0r9O2k7qkJgeIqk9HBsquInQjbGvaTDXq1YNskt
1JVMJOvSlYWJn53pQgbDtHejj2xP0oYbms8ILqxLMsvFnWJrp8APv0ij9QXYtFwh
Yawe9QTRj1SEVXNjo5rGr7gIibSXcMNnruWq4P3ktxJPoIEzmuSz0JX9+MojgcD4
DNi5IynQEbzdokjuo7VWA4oIEixuizcQogGVwgqqgV1Xy59eXn7qCB5gr6d17h4w
na4vCftoqNg8VtzQ1urpRD64hjYKsJ8DRUduLP2baHu73CZWMvKm63nWtSTx1ciC
6rn9kGeFlHwk1jf12J3M69tVWgSzgNqoMfjWmMeGU5MPrOfTP4hTZyKS+r+zt989
s36aBFM1ak2teBU0AlmXGB4evRwwsWvOyH53REma3qPzai/LF045EzUFeccybrtr
7tmx3rpFTFXTPu2TuixmRkv0ItdXrCFcK5Qcr7OtTSwOdEZEpWPh5mVxPimSw0/t
1R0YxUYXNIFMfkSA6x9ldYO/F8188IYa+ChCI3C8hbEStOQgLGK05iu3IyKXTjEL
sYozyrN2ZGzxIXrbSX5Ty/B/RpHFU2YNCw6QhYAdpMQ+UAGuVJmJfVabdbxROuxP
lD3Y5RQYiupd37Hn0WezBGdfJK93dNAmc8Of5Z1Fcd+BrJFwzHmAR/46sL2skG3/
HIuP9HFbbikLYGOnJwWIgHdrF+ye66+QbIXasIHwYtGj+Fo+BcdOxE5KbKXn4vsw
OduStpn857yvQ6sdBlVmBEAunmLfz4dQPBtNWMnd2agDXKlM7JqEEX39aS4xEIfX
SRP7Loy5k65mel7BAFmqDCpoSOyzeCqsiTPHPg/JuCCw4ZHLgH9Kr/tbbc/GTeiD
GKEUGgnQH7wIaswsHlTq2zo02M/5HOuBW6nuC6AcvXRezeHt/M2iTf6e+vuo2q4s
a5kUwARGkHxskBOyHURznO1m2EItiQaz9d2dM8K00IkSM13aH2ttTAiDsLZdjjhB
3c7RM8lFjdw4ZsWmscQBpmhHKI+8UNR6nmRQoolz0jUJQbZebBDhOFXFqjt622NQ
Zj4e0ZJTNPmMNFSvSMrVcsArzxDzL2vhP+Oq3ddyCitm5xBijLTGyDB8YF6d7F39
CuKVwvkVsx9E9pi6nJtYiCMouRGaq0IQ5fn/cM0Cjz51XlBOL6x/mz3AuMXQjqKJ
82etB+PJvooxkzqeZ4VeILyH0pXXkmJ97t242ZIrV03c3+o0KohqKViTIg+IKlsC
/aII2w+XzdlEJVeB1nC71U+kH+9dLok+1Fg7DzKLHhfW5hduGFHnD+GhiCSOzLbE
73TF+H/3szzVhxGXEJOpDMASqnyS0rV5mIEXYQLONGunRs7KizKdFyxVI7zPCH6L
hmOUAL7Fvn5+GKUV/yjHcSw6ZleCsJhfuNvkamedXlvrzSUu8GpfSmXuzLLa6viq
q/b5Bxn08Aa20sk4w1HjGjz340GA4LSAaIKqp+T79aB9jm/Ps5kVQjm6OQL8Yn6Y
FOHYsq2Sa/SRu2MVr9oITrcCpC2MxOm6+vwR0L9K9oxmKEGjJAWpe+OfQy7LK1yl
91owjqKIlglkc8u9qRqWKkdKhInXa9FQGf8g6X0IDtKqI7JKyqblgC4BwVwf20+s
fZY8qkdsNXBOqgQRciAJeXJ8KIewKTKDqm1/pxTcaMAP4xq8rrn4Jgj1Ql/AaeUT
Upr1quhd+lOFuvIlhXbYoAMiSeW02PLeS2h01wfuzdibqfLJ2wU50w/h2ONqoKeM
xT8Qikg+8w86b/aPvXPP1/LXzMGsd3Xvy9xolBTL//9VQJQelwM/GD3iP5DusaIX
qqBoPMCeJy15xFXaZGbZ6vSpHHJKNvaFNXiqDD7aFr9Bd1ILzsq2hIbOgZUljB+n
8J2GtJ7AHOCe9Bvj94Nz90kuTVuzUmZhRY3xVjaMXYf9UwN6JLy2CY2BsmJAK15N
JLPdsciEXaE7u3iy5aA7er0yVFpbiGPFFfLXQy65jda6lmtuHQ2H/q+uUbv5usNr
gnwSQSMvrD5sdur0PsUFvRuQUtjTX3vgncKF98KuQmVMIuDh8JX9Xw3PxH87WeSk
EQlfXfRHX2TZRG6gcz6r9y+mES2h/5yCx/erhb4bHXw/IRqDoCg2TvPCRD0LBLFB
Z4/M8GaYsaRv4c4uPTQtpG7N5y4PLpjvVcXIsmxrfN+c/OyTsi1aQTqND62+w9JU
P8d3sC0ojb6Qt3jz9jYfwVSGY4RvcVEGLcIiSweVCf+a6+ISjk3vD710rYQDaLT1
bLIVGv2/Cl2MC/5ZJplaEwXjn7PXYAmqAfz1w4QZAfdb/MykDj5ecRcREVyhPBAj
9VMrtCjUfXHtKvuhVa0oPjTfw97W5bmb9QI8hrqCrizHmSMOs8ZL2fnF0uRJe1iT
6Ex0DKhMTRKt4quCQV2trWxf5bvUBIFKafLs63kFEG1t84K3bUS/erU28SZIcMSm
1VF9LWxTKWshDeZAFEXRCYkwvmXDwG6nRs8efA7YPyk0ux/6vq8VoOEhGwzcDFmk
Qgekzwhut5FWtElMG4X0CaFQYSpkqiZqsXbY4BrhZ2tznIhLs7hxVjmX6tNB4fSq
D0o96uTJ/E/gTnCR+t81mD9BafPQ2VOL8JzM9gVsZSTFBuj4eCnRTI1lPcFKQooY
1w9a8g+QCpoEserEHtzplyGzM8j9Fb5fujHJi18UBndINzrBxLm64iszUq284wW4
63yO0++2XRWsI4BC/o06wArVOJivlmy4vv/CEGtLM6im9sIW54GLAw8pHOG4ynD2
d5s0DKGSRS2iti+/65yFReQ9jacHOZa3QBqAa1wK4VyA/7iROW0Se4JgtUmDA6mL
h7E01C4ipk8IEjzDSIPX8Le2L8jRVrei2d8xakOltmicHLSv4mh7aSEYNI8g5uk4
A9JefLeQvIpu1Ufq4J1MCGdcz51gIJxtfOaEb4IYTSRaasuG4811Si2ZDBHKEKt1
O9eYzRwhEL475B0+KisN+ANMDUDdp/+Xsa97Vw9obbWZQwJ8+V8JnRxlya0XGEEm
jKvgHJn2Vomn3ZR2Y1DqjZGEo16G+BIV6SvxhikT9MHMe8xIanRtJlxN8QC29/Ps
2TGaFo/P+HRL2J7FH/Eakt1lyEZzONQBGS07OECEaYZ7kea+5qcHSScuOJDHjODR
PQUHT/pwz06Tbieym090i9gR9DAi19ArfTvQ3jki7PlMYPUwkOuDA0wFe9GFaBY/
LvMTP7PvGVb0EyGmMKL56WaNbdwCHFwD8Z+KfoYaMkzXtyc0YLleZZnatSZQZ43V
l4AxDYpGVLQ4voQQDvwrocbXHcbl9U8dKKe3i4EGLrEyO5Vqnx94GClLjjC6/PWs
6+o9JRnyyLE6P2P9L/Nz3TZpV0EHSfMjiJ1jHPP7K/coeg8ScdwAkiVl3HoDvGkV
CRrNDYZ9kMqukYXNYLYKI+p9QxWzFZSmR79Sq2k4iofiE1ty9smuLhtxpJND1ZiF
X+ileGTuZaEzRcqrHhJBk7s2W2Jt5/HQN9B6Mezfyu09syuedaWsfuXqxBoWZEnv
EOK9ujL5Bj5jRnJXScPRnSEWmqO1IFSmhLjtnrvxlDpaYpIbRCVL0QRKKTKkWPnq
y35xePgb2RW2AtNMe/lZkVXKw0TMBdl/RfO5O4jbrPsj6FUU4Ql8EBYBWLfmMTrd
Ze7W8kUKSu8UqBeFCSA/WURUH809sGhhf2hkDAuv1/ZVJ56r+xuKGlsKniLHhe4B
OtGm2DyS9Nx0hhqBuPaHUFGKqIjhaOh/WK/3T2Ba7a3hDdwtL8b4PQVf+r6ixkXw
vI+H535sqCtLtsro/hsJMghL8M7E4fBCReh6iyd65KMASheEl2HPhisMDm3Q//bP
lXjoo1WxmbXTeagT2qRFfbHnQxQH4E3hUJut3rPw3q44G/qcuy7p4WIM3EsnNn9I
7QWx+WWRz84eABnN0/W6fdIG7TjsI5GvvZDgV/rqNNZDixLVxM5+QhwWDtkR2y8+
dJjr1rfSBeKdv2LRp6NyQiNEFz1MB5EY+iNn6kvW9LSZDZonf8DuE9iJaDE3Tj5i
ByBZH2fLEzLiggUOPpcrh8/0iy/y6TQDicQFayoTvRfWKGID/nXJfrspZzA6+Qyb
OAJH4VUHd8KDR99rd1DfE+bL03xO0Z3u9uGlwJ1+6xi93YohIRcTmv2zVkH8uD8s
ZnCqLW6I8j+Pj9d6vYKxtQNK+qcDV+aTdIsruGOo4C9QqoxS0uzNPOIS7leTOmJS
ZuuBJo1P92nlp36GVBOV5S+djeN/hJpsnaUhlbp85nlSRftfR3PWZD30DGngTUGQ
E8P2MrtgqrlhUcs0HnpZYTVrSH7Lt5FUXXiiuN5zubIhsTj8OmWVjb2hXaqA+4Tl
9rZ8uC4PcAyaHSumlpRueC+iVUyNAxTi6TAhwey5NU2MzqVgMzQYw2SBJMWp0iMp
bA+arpiWVR14+2fT+9jKhQrNGHFGIWmgY2jBsy3NkRCPVg+oIbr1Qj9kyEuP28vO
qF/HuIluM2nItnUJJtVNyYZytYzqssgxYCziOLg+E4p4ZFQ6HbM8AMdn3o516Q3U
q5ij93swKJcXaKUhmwPjfSxm7Rv8kWQW/IIgZoPKI/ZI+2Czd/RUkvG6q4ZaF6Z5
KSjpArX4viCvula8bwI9yXbn+ljox5gkYe7b41aHqyhpjcNvJ4t0qWmLmjRjDG0h
Dlvy/QNkKt0SYWQkONnBikvDZkLBlK6zb9WY/Hktul7zvy+ukmXxzV0XsbLB8j6L
GSBp1oF1x9qsP341ozFZXHi6Rp3Jxhv2Wp1zULJBSsDmGZBEqNcEQ4jMX0AnjD75
6dqjMsp4vRjQUjvvvr9c52ktAz4Bp/fm+s1CR824MdGT4Ku+btGrukl8D4vNrgB8
AB5KsrotnM1aZaZanDme0rw8vxPimLRkH6/SivyGmtcsZvoayByon7llbjWsOKzx
bvzgew+8kfiRnO7K7/QWHqw39V4YghlhyKNXAd7aXVRQJv2QHpYF/ARqUm1h1mrQ
OltdZx2PDB8GMQu39N6eB6R3ZY+nefitMywipPlI7SoKRmUBY9CjYoTIvqm7E3Lm
y93iN2JIQRLbD6jZ5IKKfWWdrSbEaOsrWfPt6yW1+BY9n/OkDxUWkcGHw7z2kNxu
FxwzS3dGbHFC0/UgrLmOCqIbPg9lp6nqDWVUI5rdRrHViKke2hfo4lioTGlLfOZO
y/ubjszrHKAqibKYJ8wn0wVO+Xw3R+Ph18tt0fBumfdFSeAvL1Q9Ci8q0CkLeyM1
B86I3wOLqxoWhrz+SCO3u9lLxgaf2NJj4V5l4JdK+83AP1ylMQPZwdxymGE6BVrG
AfiWDSHvtyoWnfjrP1gn6q90GmoZ6wQlKgmv/NPz4AI2KH0KPCaaq8fisFYzGy+S
HKm5DYgSrZgyfrfgSe2VskF92XL4m7OvoOs9/yHys6Qiogq2CrFlaZUoYj2c/hSL
ory9b0YIa3D88kIJ/J+UV1w50SeiRXilq4W5dZ/zIJlXIqcGdxp7OC6YxqSx4CLw
sclnfZ4fTh7WqqYGjqAh9pF3oUGiuaMsThbrogHufkRO34ESHOn2XYT9xe9VLQig
h7zsnbmQxkRT6vctaUAfkc+rMrtWXieaGwtaj0WArcMwKYwnyrDBlj8ZJADXR0gg
86qkbDyQDjRhfDSVVvqnnxPhuEraMKrFcU2x28pQkzUv8YFPoCHmKhfIKVnbrFLW
Zau3yyE1W12hpyUA6OkeUtPl93VpL0rqBb5H6ujPe9CVTFzMlgjZkCDw3xXnmXkv
M8QNrIsp6w3SDMr436bW9+eWK5J8+Gbn7CXYDYEKkNCq359Jwwc1XiZj0xUj6VOd
6QjMwtL7cn0hbS4VKOAPQI+W9be+UQRFTUUs/QXc3K87rRQdEYryBFkhzirRTJu/
2y0qIBzGg6BqEoGXI8+28mDCLne0oDpMN8dyvKY0SRIY4CMtL0/ta6AeZ8QbADbS
gj+AzyKKvlLy+VJxyqbLbkgzM+e79mcaOsJrgXAiwEMg1CEMrkEMdn+8HD+fYRW5
tusDcMgu+TFoOYQO55Wwsq3fA0KPO3P7HZWfIC9WF3A3d9rBE0jbsGkfIMtppa2b
j98XR6sk5ruU/aGp64tycnFqA1DC7YksZMkPiZ4jmYJKiUC24rN+yLoO7wu67+DQ
3Zd4rdsuVasIoeGNNUfWMR5HxXmSqTYCFaPHDLY1zPmegozgbFN38/23KUSAU2Ux
UCWBcKOONbiPJWLL1VrtVvOn2+CUFVXec2fjhp3rrmbqYoslZNtozDgJwPDa3+5c
vrNKvzj2w6wSBFE2iqkmX5bR3PmScmfIcKTcBhMAXPj+EQq196beRTg5vUqP3uBP
fTZnujDThDl8YXuKAK/yTBP9DsI8OqwblZM3Q4onUD8lGJUNCVyJssFRmGvMclaW
rHEEF5eATLYAUXp+qmkdJfUuxnEMPZu3T+lumLQNMh1ZnQX8do4VqaZiuUxOFefF
0+xzXdiuubolKzOHdMVPrL2y3CNgWn1VPpSXnb9s1jNJrubovm8fzT7KxgODsTcc
3effcfte5d5LlE/W1+WeCv38dRH/ZjuJwJZlBZZoly+D/00PNVQoSsOjT7xxtD0A
SN0Jeb5/4qZCXbEnpf28M+xeRfjoYMHfR1D8SaRhHe2JI9g5UrD7spgk7sVRXZCD
FDhrJksMemnYFjXrwIJfs0itcN5gYrp2oWyOXjXPXXA0wECe+0YxjpLZgDr+T6RJ
pbjITrZV6VI/CNAMamXHgfZMO/L/4HXuwiaY/REUXzpBboc2a6qCzJQzIWSnk8Q6
S67xNtBHCwo86q0rZsXgdVtJN+ng3IiQZtvjMiO6Ziw9sVzi1xyEVFavEdJVQ5WF
2ufybjr7xul3lHH+7Z5NUFSSpqcB/i16sz/dm6/yTaMQxCtXwJ4HvPX5xLRoHDtB
Zww5ev9Z+xdmEmXWH6jcu3Zf38nG1liDyeSDZDRYFH8qkcxR8TFuCusyzVLzY/99
ne+nU4KDLJu1De84BkYVn/RtW7YdaNXi2Y4g1+1MOUYtRiuXKRUDyiyehpp7Nxh0
RacQ8lJbgBn3YABnKmboVkx4zkQkPdkL60nrXTj5yiD1mCSzC/VkB+yfXCRoV9O/
11jGRA9ZhSBkVMt4j0gW77JY3mlk9NRmLvtjLNPzNqNk27EatagbkWMk58lTLVX+
YQog42ffr6APowK/0JltniR9BtZi0SqPyUmsN7b8EunYC6vo4A8VS+7AMw9h9sOb
21AKW98W2KMFaayC29EYr3dp5r3E8BbIOLFfnD2b1XOzNsZj+1nakB2KxyRjlwHw
Am2+KKiO/+iqf0SvxvgwKJVZNf3YfdlkEPAjmi5GpnX+OeDx8c1BIzxD1juiBtzp
QZXXlauADV1BHGL34SGFMTZgFwkimtD7F0AXIt12Jc5FpO7Dr13rv1JgTe4ykpRP
EAYx+CKOYnLm0Cn7JR6MlPWKeZX+CpfGvPhurVyNKKK6lOXC5JOTiGUrY5Czkf5B
ZQ321xuD1xgN+/no5PyPqHv1mjUv/Yxd374DajTpEMU4ZRph+t6bqW1MSHQiwEnc
4m0cZBlYju/HO1nj7mcd1J3m5fpnA9L9DoWKbq0qDoX9703/PG/W0UodGuDu6ow1
sq4vePKK8N1aNgLmwGCpOsuKgWh9753AQfe4r7j06oHzEbFUKRiXEZRpEjVsyvnJ
/gLlCWKmF0rP2PT6BU28Aj6jwj3M0BSStJ7FIYmqcnLDfZRdde3rSMgs2ZL+3pfs
kHUyEYq1dk2y+6+H+q1lrcyNx0UwmXbidOqWhXD78mTsTaRvFLjQ+z7ZKTwjK0OG
1U3wRfWLoaYABV16cIxGXYjFGmHo+DBglXwaTQvKw5CUvJB421rXraXfE/fBVb0v
z1qU0vU4V1zVPZzp1k6tky+yDCBYkTAGMhiCmmUtsFxY22QpvHWRt17/e31hsfIf
GMSw5neeZKPnLQKzwGZOJpjc5wg+YURzeGXqiyYKuHTplP4JTmOAs66x3BsVdzHJ
WKKaSUulm07C6Z8MBYNwfdA5dzVSSO5OdXloYbuZ6KsPobxrjjlKzN3ESxDJfNxJ
PEZNhlJ3H0QdoUTDD4acHR5yJaqdIe6HFVcIyR7L6PFqSP4ZFTgQbFGxr7CUFSt6
K+D9GHR+0ye0+eFGqReRgwSZhAlJDhxgez63yoYtZ8IA6F58e00+32ETX6Rg1jCg
MepxtjtR9qGG6ikHlaaumJcJBpRb2PqaO79CGQGovFo/PRQWpMblCHw1/GDsiuws
sncV5c9HGJUIRAOywoQb9DJ7EqyyivMLk7daffTEermVPDbKCv73qwK8M7t7kmgL
kO3/r0jzPKB9AMHeTGmugi0QyZEhXUfY2asNBYsacZrEcR1yGjpoCTm/9s5OQGyJ
AZiENeU4Y4CWQy5bPRKDcwruHd4F/UoQUPTdKclAdHzicLGkzOyH76HWuK9W2XkF
fuTZ8CBkp+//qEMUtKzOUcYEtCBlPel0velah4SUvBbCPIhIjgjzxoGOv7aIC/ZX
F4LXnoWNGMYk8ne4S9lTHlE7xvO1UHJRBeHnWWYbimtDgm2qk2BR03Y8wpHFqPEd
w9DGDRuemlOd3zwwcv7I238xlIJ6Q5XG/esKpi1kWMczhAFZijjBbdxrgHpazuoq
ypaNeImK9W4CzAueNFGDFlleOufSCMpYlrtNwTKLQgFuNVMiTRv7YDIh0s1ShyfJ
N0cBedu5mzBsA1IlX46myPzdIIVknpPstIzVB9maJ2Sozis5LDNQ0yJinP5LLpFF
zYmFYzog4fw4adOyjban9B3yb+8YDNHj/dUUUX6+gu1R3gBFayPihx9WIvikyjgk
O6skSRiBJcR2ounNPDXy1rIgLHW5LMeS2Da9/ynULVpTbDvlXPS6MHDtK2HJWONE
R51uABhjc6Ths57vAXynYaAjDrPOXgqv8+bPiTlQKUfoMN08AuBzjTezodwI4WFN
a5gMx+aRND9sAUGPHSUW9TWrYs0P1nrArRhNnxyZVxG5tTo1rMbRc1+qL+BWbs1L
zdrXiH7CniHg0vBo1Ns/nBZxegCeo0QUkCxrPKCPxndwVrZg+31ICogcao7Ijqc7
A8tVYWbzfpCompBp55RDbt0kaXuy+Ms5xZ4b7qPFZq/WHCeOC3OP12R+2za9EI0P
I4AZhugpc/Sz93epxyf9RhwR1wGDNNgiEfsVLG8In6iIfhc15B3unx76uUuQjJB4
8FxhSZbvJhHmU75eljL1Uyn9VZg3zKBXx8Kqm5cd7MrGiaHWqeslX43ZAKLK0iwY
dcTXn8hoeBCzIa1kYOR1LnKpMYk+FsAP6pS/sZTyEefXyKtRnB2yDztX4ZBNZ2TV
3jHSuK6cgSAKq51vxkBfLBtfBJhfh5OMul/OrYxNw3ijEJ0/E9JugBvmPFUE539L
1hVicToZG6IsPcXpLDN/jwM0Oj2bNqkFNX2SRE5MtCGYikJdAA1h4POLrnwgiSBa
aLCjUtiyQqeIa8hzGNZvGQhxXjQdR+bsMM0m3xR2XSfhgj3QkWQk1EIzXAMJNhnU
ukd/ZMy+AygbQFvJvkLSQIniEU556vXkjh/GWtBmnjS/N4YvrPNcyjJCOq+vrUKU
WRehw+PVW8fSgaimZh0GndcQ4cwqbR+mKMN2rYVgwfbX9ISd486q1uTNyYiLQJOP
UfBp9rGrkEcwtRNUAf0wmvgLgkkC4YthlvuiB5TWNa5mm8JS03K+v/4vj4BDB8kO
i9UhqmW4VUX7GnPDCkXXv6m5Kbc0Ryc1SPNHjcEJ/iUTivuQKacHQkZmdjc5yI5H
tF7BWcaufdGBq+tlpOBfN5R2Gp2lsF0x2FfeWVKgzzvNpMgTNoREcGYaKZKpZEWP
N/jdz+qLw8pmRm7UpFX+rl7q0PcP3a5Emki5VJSP8E+LyAcFvzGhmFq/NxsPySTc
fyKwPTwH5Si4JWWRQCbfgzLB/gayJgk7sDa67VwqJp1FRCEsz0C9iR+tipQO3l/w
3ChM8bGU3KpcdaYpxRdew66ygLd0tlvlBAWVp15AQ5KhLb1DEtRuyJQg91btiL1b
fpBIqssTEPwav/GUeATQ1GV54KfDb/gjkUwlK/Z/+OEsIWCfd/9boGeX+4o9ixYK
kDZ480L1SCHTwvjW/7BRgwB9A1NkxETlrQzh98rgEdBNWmo9AF4+KJuwlaQ77PBT
IzFAh3vv7UvfJe6HO4w0IIJEc5yFBzoTA+nq4Y557JaGxyPPFJhpyDMSMuBeLv2X
m+vCHfUfWSxCInv5sxRqubrm0jCVMMUj/BkacOEdUlyddrBeeaPqfb2Cgz/03JCc
cmw5HE1gAx70IIr7T+1kZ6RPUt+Lj0XQXiFKdov7XlOx0NU1fSP0/HMcFSN7oYxq
14Tu7Gs4dLpQWceSf608eB6EJx8d7simSwOCulo97TeQ8JCmYWmwfqpsrbjgIiCP
iopFXNSik+ah1sGOhgFLtorhx9kz5nNl5fddS7fcjm7Stz+MNuVzGmanO6CVVr85
oJUqDzPdAmOixbR/DWJFdwD8kUL04PnGU7l4AWC7+g93HTNH0i9RKVwXYJP0r2G3
BTRqiqU+2pm2gfP2WR/40P4cq2fG9DRGKyq4Wa0ehZM6iC8bGaojNsn28ZIQAT+V
WG1/VdH0vQIMCeMNRrjzv4q4L9DbrxbWC9gcj92U10SFQ+cLxWXLzBAjwa7aJ69f
JN5xn7yVg+nm4q+Md5swDtru7rB79Jg85Tf1kwFfDfbxTbtdgScjU4XDampUYMml
F66yZ7nY+EV+cfR2Cb0LI3sorRsSUdz84KtRpL/UzYw5Df3opn9zozthMEesggGv
0oecQnXpTFwDAbkEQ/7xd4r4yyyW0rCeGIoCnJtFH2++PEPkWTqZuBcQwhaA/Sin
PFsFkceCElwGSFP8LjdiFTndXzowJV1aeCrQMkGHL3wVZUYi4EIu4HzQz12RAqaE
U4pv3JcWKam+jocysklFqAtxxXFO2CgykNb1j/w8Wv65SwqxHT3iGd3XL38rBejV
1P/1kIlvpaff+ZwTapjlbmbMpgF1nX5kuJk+SUFji3f299SUm/tgeUGqtz8kC2kP
30kHx/N1oqWW1lLidBqZtgsomzcV7p9cxz3pO1sejMTa6cPBCklC5sZj3qwW4M0/
lUR4yz5Iyz7KOHusSbdsaOwZ6tccIRPOibxoJzdIvpDPjDt3875DN3ycz+ueDoAD
XyCLtGdD6HiBaFmvySU5Tc3ncWebS1OuFLoUMx608GvdnCdH/HLuCnkujp7GQ3LG
yaxJzA++vEjdguixeuHiUemh9+HgVNYpJ2sXMDjs+hyn0ChsA5kY8C+T0bIi6hIE
JHyTDewxD3yY75p7VQi/05+22jz88DJUjxxx9B7hhjBhP/27/vDKTkKGy9T1h3Yh
899kbMpp2Kxl199ju6YHGT0SYo0sppAOfG4Y0YWT2Tv1lQmWOwIq5689BKeAeB27
igPwRfYvs3OUUwVWPFnNNxpGJF2mDDNOfSrQ8tm0fD+F0C/PMRyGgzEoBQKiQVDu
SVvQoqJgcMcJ/aQWhpQtAurRSF6GizxN1+J7SJX0fGQo4XEjI5RuBaFvAlPgJN+L
Igq9zr8LhZ5JtWaluuSUu+zaX65Tc4TbGlQ4YXdR6BiFxu2r4OwRBlbVgUUQyD+4
dhhpRFOBV6UKnnN0PDxfMMKMxQgAh+cE3VsAwkueXCzchh7/HpWgp3ocFtAYPKgb
aXvedvD5Qd8emaYoU2niu//wsM1sRtDmeEhOehDctQNKD+fpDu6sXPudC70j4ZI5
Akq4EcICohwZZk5LJaRr/P5ILjbqMegzKq2NtByJktOtZkyEyyJqyK+Crz2QaAv7
RMnsY+giDPrNitnPYPpyI1+jP0R+w4d8Y1BZZOoK07SMgWbaHH02Jx9rkO9HzeAY
RCumT+O2GjkiWJRrg3Syn0S/fMngFxw1eNCqr92WPaxaJiDtGF/zqJTyzrrvU2rR
g3v0w09r8lkhkHEPIV20VTVS7+Mut54j74IFValV0IwFrR6ob3mT9N0Qb1lNZbWz
8banhlsOerAxMsRFj7Xec0mMYfob6MucAuP9owQOOK/ro6QSGVZpaV+0A5cbk8Py
tab2FVfURiDMInrC8xC37bnZfLkIkaQfSK543WeNFhumJrnDVl93Yx/F7pPW2Lf/
6UVJFEENYU/RXoBF0Sx7OuT3oOkc1grpLAaZwYY30WP79pfMZcnD+pvbi9Uhm7pk
l4lmUlKH7on4LCzool9eh4TrR68HVuwRT86fRQn+7ibwJJwSbI43b6Hwwe3MxHNx
Pnuseuhdi/e/qeDN246S1bZdYR6gvuWXsu0bG1ycz1dT3JQ5aZ9cCQnUgJcqeZT3
Jup5ZCYRbGpnYXcRRD40oVYWDxpHMe5W25Uy5iGXR34Yk1gdBGH30DL7NQR/hjaq
rWoOoYpZLCi1jIX39Z1NCRx009UZ63njuQ+BW8molcc87PYJwswMvTeFfC2zkFGx
PH9ou0M9Coexbhl88Mq9J1cCRLT9Qog7nSfNJMiA6Tt4Dqh+BW037L2GuC+1FPDG
qP1y0L1zFzy2kIfEyt7xegN5xJHYDSRaoeZqWx+eJh0ZrR+mcIaIorGzpcIawrN7
GMxlnZ4YFgmUwNwYYT85ldX3Fc/9d2su97JZODr01xN1LvUParA5Aaq3JZD1d0J5
A4FLXx8PsI7UlcEKQEl5pKeAZ2V1zgViAmGejlFiviBTcwzFr2v83wiLnL95E55Y
Z6XhqVb4DZGIIrmxSAq2yCKL1evIqHhgPOzatd3E81KmRxvAIM9vuypl06nyaPM5
cqk6gxUj2qHF06cGnZXN49a22honhN1cTqKknh6gG2mYzuwOxtPIeBf3DJ4w75Jf
f47KWFj3czGknWuB4p26qXEHacoCVgv23WwgcmYHCd8uznN1JyE69jzdXq+qR0e7
MD9DyXkW43ZvUBAZDhF/BrATryqUkmm50rF1knvmRlh5ZH5ZJYm24O5ax4M3l1J5
zEQHWV78gzJVPhpIAdBGtZNE+EBw9Qo3dKGV4wMU82IsTcXqhaNpnLYLJ7c386uQ
bOEOqOgZCCTwssYdrTqKgaIZPSfTBkN1CQEbj/4xqGIPlV5T1HhvllHfURcQXtzn
aN5tYhvldOdHmWT7XqLYz2Adpxv4aoYoEiFId3kebHsgxU6QiMnACnaLJkfcywqo
45pXtChfFAkaWrE17SfkpGXNbxsimPVM/4RmecYyLqyC8rYbssOFMpCCuODePMPZ
F0GQY8P70EZTHHy13+97ZNwLsru2W417FxiwrATx4DwSRTzGRewFC+1gjjp4QSn1
d0flF+VGvy3jLd7PLVOTbm10w4KkicESm0b9FdpmKx4SmeCMBGorTHBOAMM1/0uh
BSEsGG9qawvLv8RrnNHXfHSEumrIJVjWR4J1n/px2OZ2BwEHepXh0ire7g3h4gA6
AeaxhznuzDBf+yoByGIzbhUUQlOjO9xt8AEl/PPAevjKIw/S75iH1nQYM5zj1+c7
W/mxdTzJbwfcaTPZ/gKxA+vyAcGjol3dlwEFXPJo7gThFKo9ciLr00jooDo9sOYK
yRqCj6v0Cq5dc+ot/mSd8vObmcWzoLVmfiNTyuU0hL+pVvsXodwr/d99n4lxQZzi
1RHcBx5WcDXXUJzzXkRtiGmw0NLx3GhwhMWtIXn2B17zR8zub8GqEyKHzxVdPym3
xAJ67TUyuzD3SFH+Vvvv5yrF47PVKaSBu19qOJg3dyYQcwMnFcy0ebjYKLG60z1h
Qggjk8RdF6SgLIpzGC0WgrSZY4vDAvU0vDP5oMi3tn/PqolQi0Viax59ZSlEs/4I
XGiZ7Vz9rAV9XUkpckGEQ2mU0OInvvOJZxrWjtxGf35jDsO+1iYXFOQxMkzNBnT0
ECs27M64MttQgEftaZrwaRL0ENfFHiT1tAL00CYZAQe4RJzI8pVwDVfg1aLOPtOh
AkP22pkKjYc7/0BJgGLWNIs4FIh36gUT0oPaaTy6uWqCCPmeH27/AosTYhAsYVHH
ELSJraQSxjJABC/C2nLL1SuO5djK4CCjo08Bi9vvXIVpIh8HkvZ1zaPsugPlExPg
uYtUTxa6lhC6cCNgEg8pws160aXKwVtaW8pcK1B6/dayA3IoFNcLO2DROXH8R6pq
tffG0zbLm1Zr+T2sp9y9L5pNqWSFxpUhm6qnJINQp5o4p0mvy0kBkLAYBxnWmPFj
c/pINP4YWq/evvgLTq3VUWriEXbJfukp4y4nindLEVG1dZ8yIkVEaBjoHpqyFxPB
GUCcqSkiqrVnq+8/FycK5vDMyKYZig6BBtqcmFMpuWCG08GcakS3+UkMHKTA801O
y3aacLaa/qW27Egnyn8tXMQhugT/xXJGkLe87ismcELBgNHLWI6G8ZKyIJeduj93
LQkXHeCY552IL/Be1uDArB9mZK3SZhMlVkVbM9WtVG8A0g0ygDrf7Xu1pS5GuaYm
yjh+Tzi7bpT7TBn9bw7Jh03/aVKDDIa21sONXi+ghD8l2SYilUf5sXXIJ/RGXI0J
6CpFieJbjrRjOR20WTantpG8kW0L1+Nof0ecPFvbeM5QFfd3t9NY4M52wr341tkb
qYC9M/upBtNq2kWIolhjlCCJHyjdeAMsPsVatA0zsAerFXCV8PKli0SltstoUMuQ
KCoGdSaV4nEwoA6W9/VH65FOXbUIqZq3j7S/5w0Ther9w6fZdGb/0b0jtIrtRkO6
lyo7ISeqSy3IzJaDBWxtvzH2n14IISoiN0kiQ2+3t/sMbjX72R8GkxtQS5Y7nOjV
g8VIM0ShXQOVwm76ABf00YlikCEa6Xg56+iWWMGXZIoqs5rC+dVuHKj4Y/n3pwc5
0vtDA4ys5jVoupJ0Yxs263pnxT3Xv5sXQpnJ6eudGIEV6+VQLzRVlk1To3WzOgBM
8a2wtkYO9QtYh9BuNS7fr0jncypcgIkvLmleMR+YLNwHdA6g8EzpuxEIZTlyxCqB
jgXpL4bic1jB0K9djQurqkiALc19XYupazfkttbBFOGqCnuly6TTWP6rChZpQrkf
TEahB8MQ7lgiKG59MawXyZPPe4BGoKs38zQbqDO2NSfp+aRUleWGQOzk9pm1UtEC
h3xAZ7kT2kdp34Dw+qbo/+r4rzh6Vn6tvw9N1Hu6KUH8j5IrKEwRPnl/21hRiwpa
wrOYa9nxRyfT1lYFuGttLW03v6awCnfaBPlzGWSLJQbKVXJEZ100yc2LDULT5kPM
fDSzuoOaBhVVW2QxHkf3XScvsLqETOp19FnmAS3r4Caat6t6BKV9kCeoBrdA/MOQ
6nHeqFIjpwfMziHT277dJlW8w5fEkK14i669mi9G3IDjeKfED/16Hm+oHDJhsSYv
mzzLc4Z9ZNP6lgHwpZA/Y/zgCE9WcRkEzt/qlBThMlrMijc0TqiYZRQp9u+nFMu9
3BrmCYAfWGS5lhUTUyTogZVBRpJirE8uL5z5/WkVcOLeMj/HjhJ7rWsPFUVhNGkN
o+B9GooN0RG54N3SaffRw7JMoN15e7ModIk30kbqNeegIv0PKyaylODNnKorw5Mo
iJGKQasiFl+Zvd99eyWV4PJUmMv/nXoEV+sFITZlsaRWHsyBm63J2LvukRCxbaJk
bqHdrf5my5ewtNvedU+ZPzOEi++blhU76mLEkmpA5WIPpl93r+FouBoy3NHZTgib
HqTLoxEJCqJfOYDNz7HTRfflrSubiW1fV98jNrZITXStkXtrlZOOU9kWTGWo2rZa
989A9EbtNSnTyqDKwB2oV+HMK9Qg6WXiXaFshqeFmqW1Ub+sHWPj1Ha7xhNtVwUD
kYeur/GaFwB5fgdqxi/4Z9BrXxUBHUvFqw/Wf51O6js2ufMK5uts3YzBx5fb9Tj/
8nHmRjU9EMUnh3OpOXD+aQHNmdT2kGpWkA9PTC0g787S7vdPBk4I/sfZv4kGIKLM
YE/1jD5WgtalHz9y+ZMS8+JqyCGYIu5oOvd1c9QBNq2PR+JdPIB3zHnEGJNaOUfw
TTiCElx0h5TGhPSxLAEFN/w6oi7zd7xPHEWm5RFqbJmd07L/cnUn6gE7CcqJ0/Qf
VZY4pEdbqxTDWma2Y0OyEnqUXOL4zpqyTQdridVzO/+1bGO1ZyFI6nrRqFYTLl4y
PjK1Mug5kXGJ7ZXVFZSxIn/DOUFfkPrvNOGh5/GiClj35kWVDWkZ1RPVzzqEqmY2
cK1CkxwREFXPSppRVA7bEcqG9rC4A26y15JonkoIQxM8f5V5I+2n0GaC7WIfxGZf
DDT6QFu6NvI1/VWuFipVg9C2XyTriqBs7aamGSl8u/KiyArCaNZT4lAdNC+xAk9b
Jlprmvp1BqzH3T6OUOoEWPfQI2N/PpXTAyXTk0cbOVZIKikhIPRdkNi7AXppibMd
LmDXzenn+A5+Se5zgbsCrQUixGDcT/neBNSWk79BdNhC+P3Zc8I3axHaHw8JPqwu
sgjl5LwWGMC5b90QleVoXh13lxhq57H88u0wB+OUXOY1tIyFUN+ki+PSeXJDhCb/
s/IaHDlfHMNTkg11aaW8rY4GcQbRHM9hM5ely9z7xvz+Bj9Rb+T/QnNkgCOX8YrR
kydDAnlZmRY+TTO3q4bgd+QNorYcgm5qUxuQSrnsLo3ZbBYiDQnGhhXVRC0lzU85
LYRLnIcBUF5XUW9u3G/RvMxb6evD76mm9X7Oc9onZ7ZMJWzqOyWQAfhHf6EkQiey
QCtfmT/KJBcLJq3eOv0qqsoNI8JLXWSysPaEMTqccWmDvyH+Kg5I4xODQMh6yNsB
bme6ngX6P9+wHxLBSIQkfPE3eZEHMKqrJEHaOzSgiPAL9HeDU0gk7JDUotvcigLx
fhK1rlY5Db9jBYEtJyxxhnFw5wQ7FYXv8Wit9c+fCoT0sAPjuLefDl8/HVX4gEgn
sMU49uEmrL/TItn7UgH/BzZ8/vhs89egAwFIhPDl2GE21TU/U7nc3y4QxebbtnhD
C3c1mwYCkDApDK1fJU2PBeqeiVwov0xk5nl39m2pqOgXQXmpWwfQaTUCMOTiukKY
W2eSIkPlScQod1IAujul+Lz+yeLIsbn/VkGoxAOHUlGyHUX6bP4r8gj7m7Hi7How
JYRtix2wg78iWeXsvmetSz/GIYeafR9jL19xlWt/hapOof22//hMrQJYhmM492//
IMTwWIw1Ua24Y7y5pRuvUYTk1HM9Ogb9uHrdTqzv+Qt1rFv89a0hADeZK/zs44yg
XecYWcm1yNG0QfYPpjeoeeYn99/+OzuJ19xAULl+BZP76zU4VjSRB2eT+ujw+BkE
ArgYeeSLuujdn5GO+GB+wgiOPAu5r/b4Za6xOjOaIjC9p8zV4oaO/hnK58ySSptC
pJrvbvRu0Z9crXUmaKVUDZuRrz3kYItLxR3D5OqHWOARbEQ7bxpfPMBQ8qeimVOi
atmUnO9vNw9vU+8B4FJ8Hxu+63QpFUw/qDOodXlmn1hflYgkHbK32YmZxf41kSml
NekgBs+JAd34ESZnF/gM1MwPHSQ27yIyg4FolZL/afN5g02yxWhPmn7B3DX//N51
ocoytrKCJh0Pz9ZTWCFe2sIny3jovLR/qfviuG2nZwZ+O6RYc6rRIIe6Ze3cmwtx
pBI9Ly4wCpp1rpm7RrrjHbH/gtZn+zU+Bo97eULLzMUJNzyZFJ/sNDRWvvA0nLdg
6yU30gV4+uVl0UKoq3b8lQ+aFgDlXK4RW1jRh/eyndMtl6f3sjJR+RYlyQEMn+Ff
Co6XFcKKxumtFYCx1uBKROLTcYFHb8Ybv50GByHhwGoqTmLAxDd7iHLQhgD/AcX8
nFr0m3jcVf8EYBe8rWpqd3k+XDTMMEQbnsc5WQP5JepX87n+cIwP1qJx9rc7Xn9X
RY0FcVp0A3JOisCyPdXtvzWX6rmYnQz5Wjqp0SUrNwNll4/AWtZbPB3VklxbwAAY
WiXqVg74J2zrBssPdo33W0bXbyXACxpzGK7q47hdGEPw1Yh/HlgbWqyjLPUaGK5P
bRoF/0AshZ8MCSvE62ftGTysX1Wt0Bo3wNoacQ8YBrLaWnG0fw4+4VXTYHifHlLR
GvcH4l5TUJ+om0HeYkwVgIzfZHrgy55TRJlNT9rkKhBIKBPohLrLmGmUt0jsLWdO
YxWMPSHaUpPx+HFQWD3BV6RAHW/iKDUrRmV/QFLXonBYJnrVzRTRQCW2euO84/VN
1gH/cYy/f1NNNYAZ3VC9eat/Qigqx03e9zeudoN4lkaoh2l+hHyTuaoNxds6Mm/n
0WKRa37+olsYJU2rD2FeB/ynjxJG9ffawajoIOiKXeiPiG2ju5GC75BwlohAmSJu
Z1IiFGlUZ/RQS0t8uhSBGhR8ZORxrF/xxJ6esOUYJqpbTbN/oIrsP4aZ1Rx97Kdq
lyAnQRVvSCCF8egeL6iquxN6WntL/nOSdJM/hSHpuUVwiiunpKuTQ9/mYpgtTe/k
AGcKwXI5Xb6r7pW2N6feLYOL53HeBqRZr5tjcUJtpEyIOWYDN1evWzDJSMwfHO/2
4tEnAQqvA0hfT1dAESlsuzZWalEfpUPdYQ1Ix6BOvapOcBTS15KN/BlSYabAaX8v
2aM/Lvyg/nr6MtDR7elB0kyikFdtG7VTsQSkwb1MmnKzN9MIqXBaZMhYCYrdz1+n
GoydPgRqA02xOvE9TlJHwG2PuSG2l8+IFwQMUvDfo1sF8dV5Tpt3FTltmkEe+65D
lgpcKgRi3SmoCtAQ2zLQBRRpSmyvXEqX2DJeE88a+JbdYRu5GbRTXrziT9LyqEgj
McTS9a3aKeqV9lQf0pEhgoWsei1cnaokWtSfgjvvo5rCcRj5uWkmEe1L74F9J35y
7XXiVev/ERFa9HLBoLStuIPHmBlT9A+bJBpPi6gsAFgPaYFM7PweUBbsvqwtOFSC
R8Gx9kuq/SQQzb8KAyxDeS3pZOCo8HD33huEX/INrbQQ5C6SZWuAqFYsqOp/bcBw
L2MZ5ZoGEFVXzim65yaPuRCx7vY3DbHo4DoNP8M8iCNGMdxWFB+MSSx4NDJJS49q
10s0cWUvkGA3ysnN7FCczh0Ygr+7jdqLvORdd6j8SCJVC3FIadDkxdu11zxKdV0g
b9vdxBUaswaPDPUIvSNTt5mov01V8gcBNG4LS5Jm5fMgS3723An5bz3RP0UfWg/U
hftMjUA0q+f+lobFp9aEzGJM9S4PNpPYBgvrOtpeaiPBGygPYa7nlFjY9ai2bFMm
ca/6pX8OqChuI0dESDcKWqilcvaKV1Jourun504vvTmrlm6y5p5pPLV45Z02h9Mq
K9m4i+XVQStR1Ej51WJkjy59v7WxEqzVmw7TlO3EVXGSKPNcPO2gJJB7En7180w6
68lcL6I/KVD713HavRO30ozf/+uoUIrahdB+VHDn56SC6EdDGIAmtsdjorcgBaIc
/QqXK0+irRXg7h1C5vJLqfvPmnV3zgqYxVjEAcsqHC7b+AnzLynDiRUpCWzPzRxe
yeJsJPsn9UQ0Q940f7oauJgm7AJz/x1u8M1gzoUyF9OAYXEw0PJ3uBVx0rac3E4T
Pf9BJ/scJqdrbKsmj5OjVXHzvv8YNMLmSUl63CGD1xd57NOTBkaguwUzZVSzV/vP
TJo/XaGBKuvNGfR3aqpcO2PiuuGcmP5+w2YMZ/ivB56KWfghmkHnT4V2Sl0IBqNL
HHRJxAWIG/ufA8KGwr0MtBYHrvSlAIyXH5S6hjl7febsaqOqJWx532tfIZyp/Gog
3TLLr3WvwQPr97NHRUIDv8/YMFGRe6yMBxdp9tJGn3/HFriibctm0vzTS4/xT/we
Y4Jkt9FLZJu0edYuGcpLRpoLItyXNPn6ALVwgoOL9a4E/vzG0QbrONfA5HQD3LPk
lW184T7u5ivvZmbxWUSoOM2eVl1leT9koPfX3igZAP7o41dZki15g1Y66/JOGuJb
03FBLfdcDI6f9HtUXjNK8BO/X5KCd6ZPjELa6MxMo/Dq9Wm62gCRfbzlIzYTqw1r
ocIN8MzS0Ow6LdMcPZl4OxQFRByzli+D5OFVY3v7UGFH6RlTUnmrV1Vn3ltFfK8G
Xk6qWLsy076Ifn1PkPk1GvGUiLMOLvZW6Ke9jwbtlDLo2DiOB3mvfiU8meHqJF6Z
eUo8jS8aXnG6iRA1gBlFNKs1ZKHRdxV3MWlQ050CdUQPgxbog7PnqcfMOftmGCk5
iB7XXlwqcQcTo8qRXI/lNz6jc4VHtClpuWoTBQ3yx1sxlQrRb3wpNJBhiG88Pwqm
cAegnPUMTxSlAesoUHLQbveXqpPkW+wfcx905Oqf45TTN5q/l8Ssujb5msJwmDzs
pMgQDtnN+8bKYFXtDzuiaVBSp/j9M9Jdz/I4/KGlSIxCJf2zWiv1N8b/fHECa02g
x7cvE9WZ6XzraNJugk/sAS6CUDiPrEptDdoEo7KSPNuKal+My6tJ8EbK9XkUu0Jo
2e2Nnn8TG/XLATVVyIiwX+vHJhvZKE8O75p07TQ+Dj9z4vNFNSCO1wnsWkvAueJa
9kpi50M05RuVSdHfC/NEseNcX1aKUPcIs1ZKJ/SRzDLlODmikET+6b1hhblnOdnO
iDoPUwFoSGH5DShmFSyFMeaeFvVyK9/ksI3Arnwj1F8AuInPTTz5enTTSpQ3TxHF
nrxK8aMCsvtci1OgOpCqfyUCKTUmMAAiIzu2169DWhZ27oqJ6Xj/hXRYJTRLSNZf
htBT0T7EJ7DNQG9xZB/tMnKfAmea3sdqpQler/MQRY7oF3n8bwoyrgUxCVyX14QM
8HkAqvCxJZA5/X3AWedLgWfHPqypfehhIEHG+KBrnucFVRYONhImJRUgwZZ2wWz4
iROPumDxIbvKh3GllQVf43n4C91tDBus83Zyo6JJaW5KshSC3neApw+mQLfbO4Gd
m5txfycDA5DIwgga3wfNaqUWckR4cCTc3UG+PtG3mmczmyql6UNzdwfrewS3+sjk
HVgksMbKdcnW1sRwMuyIKdh2rpJSqeuAdjZ/PBFB90YipjHr9Q39gIPWGuuPSPPa
VeJdiW4e7f83737ykIZDkYvgzizNB4Thmu5pBL2nc+itEcQCk3CJ1IStljV7K9/S
r6jfTcZDPfloWPatyjra0XeqcIB9gLqHXOByOBZIRjIbMLThBGrVyZ4slDOBGnds
tMNc3xBvf7QIu2UNAvzXEHSOay7s9vl3VyVLIzEWt1ZlUx6ume+B1PGY8G5UvrxP
Fc/+9ONpvIOK60TWbvwHX2k7vMuOa5jyWakymGs1jitA2rDrpv8HzaCQ3fJzX+z9
1cmgBdeyKC+fgWleFGjZUpuVJSkhwrHciCJ4koXNPEgGjhZiGv5BHOqJeyZT6f94
+PJoGD+JEIrAZ1fWjAfcTyVqaLuXPAxhQaMeD2g9fM1ytCFRRAA6isfjLgD8FTgP
1daO6951Fteowln1C6eSFJwbXgapIl+q34t1mv+/QHMs2MkdbCrq+luhAU0z7W+d
DG+xQjUsFkcHmzm0wpSnHUKITTQvElMK+37Pg8XTmwI3NUW8eXUOipEZ7/I42YDJ
/kQpi/4WkvXz8EFNmaYkNe/Ep3dxKTswCqYOocfNKzyNNSiMsjkw/L/tQ60rqAdz
P3ML0oFdJolyOPE84vf3QKQK4BrJ2WirYQjELkGwCRACEeSJk7Q7cm/sTFblXLe+
rGD2yorrJAIaMG1Lqdd9+3wobVvnWjEiRU5m+76Q2zZI25a/7KW8a1lE2PYMiFXD
OYHvrPmU+8EauqciATe5nqCsho7pu16tfLGZZF7CkqTAdU9aQx4EV9wft4lteJY7
P3onxBlyeOthjW7jnVvkaJn5BkHc5PBckaPPC5Dc2UGoSEd2ja5qfBuwelpwKoEi
BNU23+n1/zOuZ6JkNB7hL+VAZU3IhDrLMhgmSn+CvY9AQBq7POCmhaZ65b4Cxu6N
Z7H6Dnsd+Cy9hW5tH1ajMHjQeaOk8tyPUxwhZBeI9s7ZUSrweowdEOSsoSvnN2ma
NxWU2kJx0SrOjmcyTJA5VC1UbIQI1iVUul/hOcyYicUBWGNR/wLskp9jX3W4NtA5
ZeRnYua7n55LSfVZiy5lBLDDQdjkBhlbdjVDTBXz8OU2/JwlZNJ0/M3k0h6byPhU
bXpYHLMICJk/ZpCLysVx4neULOpDJcbn0JtiywgGP2T2NoFemZlUJWS1BJ3P6Bl4
5Z6tXDKQbkfarap2rGYd+M05B/b2KhHudJq6n7/Q5Mn0tI6ZR4e+OQjtHO8uOo4x
Qn3nh/Z6L0z0QrOTe9q1sT2cZFue8Vg2D8ckUP6GjmIDm0mB8ZlqHBdSFPh2Ih4g
5ighFHjWy0kmbJNsZ/nfEJReS8Esbou7RPMPOG85iUkXMbXh9NLipQ7PLKBv3P7O
jxwh4tN0T348BqUOfR4Z8l460YsGRg7FR4rtQeY3YVfCB3EyOTwAldKES6d80H69
aRRghz4NWkjSuMS/lJkIEQNyI5YEXERGwT1+bj7pN3IPpElglpsGbsje6dmKD4vX
vE656GtSjBscrDf1brb9Xq+4zv9tbGYz6aU5ZqGvP9jLxplgz6v0WrtbmUnHiqYM
/BdxB7cLaF9TzZ8rGou4nOriKpEoOeHPBsnQ9jv/450fBwxU3lXiob02P9+uJ9jm
S/zcxdG38QEHbjp1DaEbvwOoefdwZ2E/g4oh4EFJJEsVRU70MC+H1wSIUqjit5Lk
tL2byuDH23H+w4awa5dUrRg3w/KE89sMRg2Pc4qTDyIiCMPFelD3o900SvXBjI1J
HEdwM+FuhE7U3g2V++wPzDRYWkj+auC1H4RbJzyy7qxmNSFxYFeTAnxd8WBKs2ev
TEKFd0RBm6vR5SnbLZKJmqbCPlm4VWAeG7MhR0ZTZORj14f01MB2Pmhhn1an5AtJ
BYX2XlJzg9Vj1+ju2wvEGs0FBRcymw5c6VP2lfe1+jJgi+tKA1TLkYim7DvjsRfV
xhIBayoCUyLd16lKbRmfG5A3oulojubr8OaBbnS4XRz82uk7c8o6MY76I/VJO5pI
oiDMDzSkYkjpPl2KPN5OsRrLPgEPS5yIW15TDihoAcbwoClONkO6D3awGgpharCP
oleQpixc4iO6Q5ZSRo8Wlr/3c7I6J7JlWOYlh88BL1ngQdd1M9bkg308FUoLkI3i
kwVYrDCU0AYadCsj0PQQ9GEAnu+RXid9f0N7T/X43WBFFplbNzkW/OsNevFODxUB
JkuunBj/bYQ0iY5Hw9/A1DK8DWkTJSKVuilJ6cWI+jlVzSrT5qSlV0hgFER7FgP7
WLWJ6WqA4Xmtki2gcf9iUB4/EtbqLnHvSy8YlzZTZePfJURYgU5fI0JC0/4hALDD
f1bCEaKVNZw+VQAtQm6cZGBQpEt0nAwiHU0OXAwqIrWFeXZKOhfNNI6jNgE7iwhh
QyEt5OTtONQhO7ayr7B97N3jVtFTWC1d9zslAw8NO/eATbugAosIiUSuyyfty00s
CZjHGEZ0uTgDK1hxkvpjFOkP4IW/WdTRSkPZX0Oz7ekVWwHH7nva9MRUKTOfeaEf
1djvYBuwJV3ym5fWcsoge4MYPtsykhToNj4cRhN6S8lKME3fsqGWuHcfBcZU7UMG
j6otCXvpEHyaPDGGNNuxwedCRrvSz7CLIxiiCf2I8fjDXlazStoXMluvMSt9FGSb
Yx7pJUgjs6VT0Hj5xRXbjBubS7dybg2TQnHE8UrjUiu1aJ5IG5Z+NntANw7N7sZm
jB2+j6yF9JCQ3g0254Vb6fcy38NTUu/R3ZGLTesxfJeDaBpsUvDy0Ut3J5uwFnCh
Tnx1SKy6/CwiWEsQBOGTc9rjYNIgXE3VU0IczVIfysjhuMb1N5neGTNQl2ajT5nj
QiqU1EzIg4FyglNbfraU0TgFzFulHbuYVaRqO30DJzf9ip5NggMgevbHyDmvvnYJ
AFeTTzefeq4gjnVCj0njimi3iq1deIR93iJlTSsoZDkZQvlt7iLVOy/DJT6e4I/Q
s0YZuNgczTSdnzcDgbKTn9B/PBVxVIgcbXmu58SaDL387kivrXHx0bsEVwaqRPU/
BoReCNQw8KZqEKtFGNyICyQXMm0UKYKWRZKiJ3yUOAiO2tVLd6jlBU50whZPq9cg
NWxNK79bNExnH6vUnEYWH//rVn3+aSzuDakHIQb5zKFYhSkL9CgjP1B9Kxdzg3cZ
mCRDoSzx9rFTBGOznqCVFGMwjIep5e3qOnMa4b626IFI0NUrKhVJy8oaB3LWw5WL
nXzNrSRa4fIBUIyAvd2BhlItJ06eFOjLLd1QASvSPhbyZQBsdCvPmODiTEEXJk9s
jpt84+05gZ/6803NwWg7HrVM2cmswgcQHbBNE/D4palcAJxaMdb87YV23TIDWtJ3
2yqlZPHMXv5C7sBhm6gjdD/d3y+A3MkJO7Jx1ktryZxVdnhQCdzbpKoMLcvW4UEy
tcstCtDplWNWY2maOewxueEa4m2kAF2Yirld2vPCmGWkQVVtzzNz4vR46Fx5WkC5
u4n34EPjID3E2SzMtUCXo3vs0qGM2kBPbYoFPCfhDphsC60o/xqXpjPGq2YsKb4v
4N4MjWWC3Nf0NbDfHGroHr5QCnHyz2FJBosGFt+tB4pBgBzrVZQZUa/jnJbDYKo5
pOVncAvA784nQJDTaiQ6+fJSsOjrDc77hvIJLkX9mgms7z3NsO8Z3pR1RotApKga
Yo/oukS3MLhLlomR1DxfDPk8pf5idaoOTHgy0aYkvAwZ9gVTowrvi9IclS6X/uQ7
3NX1PCTMg/Mluu9b4WTBn67jijSNduJV6k+A1gGNYE2QNAMIrTa8NgK3Rr7aNPuh
LBb2Znj54PcWi+GYj06kQn0L3GcsKU1twdxT8lbAlDbpiftHKMSS9VJwB0pfaCK7
Pn39//NVkIy2VsNyTA0ODFVY3LZ3w6ssiGePiP439TYQ0HvbCnhc5tN3LxrmRfw4
YtTAbuCJ6v9iWW16ybQ49Q1Ndld14eWRo3VHOyB1dj/uE2nEPPA1R/gj+vk3MX/I
V+BQj+gFg2gOTvN3S9jo38HmzQDAfKtDJWEYuk3r6RV/8S+siNUV7Px/pVpLyERY
h+iheTNAy9ZnaZTGyScGsbSI6YwyA7e7tHM15+W/oePLFhpSl71jazQxJ90BLqsD
6wxGQAHweZZOyH7h/oQR3zoGaWQvN+A78q2c1NFQCqPZ39dCJVT1yuDo7uyxgYN3
8+iENSXmymjWqYTnV8CLI/2nYt52c+JQNEcMc4bxgu/ByyFXSYfzoWYmyn9dgh0H
RlmuPUnXnYHI1TXoMhsgGkmyVDAVAfYzjMY5n6tFQNAEFuFB5GJS1oRgvw/Gb7h7
h/jdK9RFnhdG4iK0jj4USgq5HIfhwJ1gsgRjR+mwtim3Aj00cJHy0ZVpas+WoqBx
AuON2kSLYDlVPRZhwfI5YSSASpIlWvZbPRD+OLssrjFmool4sM8U+u3RGIG1vBQR
EDBLpi0ZoSb2PExKTW279zT+cvoeaVkVtocP8jVDja1Pw4qevT9ocaS14uqkn7KM
uMJLMrIxjId/PSeGps6bzJch/TqRq5c9nv1gkZ7sbpyqyJAQta+03ywurdd9F9qU
HA7RpSlwq0dsQkMgeUmGN813vigvvg0S4880NVwQkZhTBnVAuIVl7ZDPn54aF2oI
1F94VQMIcd01//0Jx2GGOh96T/K6eZf/CHBdPnlas6tHBnek2piOcE2JY+bhtupk
avzCq5BGW1tODVgLMB7tCJYyu9hc4KTMCofWj2LY40oBo2TDs5LlByb9mXM0h/fE
5D53F8LLAT8K2fK1dYnyj2WlHYc0K83i9KSFEMTG5XFIM/HLH5q+0PUlT2iyFf/s
3Zv7NsYlk0m3Hv0m4r/AWN7Ispldjwx7/M8S6fyk0YySBu2OfZZAFseZdnt5xxrt
leKLzbRQwt3j5l4+01zbNcvBllPK8TJD+Y4xA8Sh5y/TyTtNAffX/Br1pF6IpjT9
ys92DPBHj4Jhzdy/aqbzBti1NzzBAzG5alvrV4M7hHTS0VZeNh0QfiNwfEdTaAj5
bvA8o7UWdNXHWrAgJLU+TqyUcBgJlRa43yOS4xUxsq568M4ZmiS/5bNoKLaGhB9a
OaJ5Hx7vrPd8vzLY+2M3coJqkGH+RgksjwoIwhyeB3LLXhrtF++pQQwv0xb6qjpY
LClSPpkeI+hB5MHZkKm1GqXb5PbAP/bqMLoqJ3VklvBmZbJN1AVfuGSn2ZTUCXhG
9e5Y+urDySQPoHLCm0oJV1fLk/X7kYiSygORyXEzji19p36eLpm3MfPvq5m7PcQl
fI7roFpZOcPtHlsoG3h69K0D/GfWonK74P6LOGRI+n1WVnihT21POPqBwUzbI3Vf
k70ubE8mZPUmpj9w0f70SlKeQrrpllE2d1ZFL3y0mf4Ci3iN3W4QEjRe7UktGOqs
0pQrHHQ8ZT7L60x49AoM8LQROs7Y+OdL/3r31TheMOEuqBXuNtrUVq7nzzLVkwkb
KrJSX1CqfbsfG7JJT9eZ0wgHFND+YXQILGQCT36hf4DY2P788C8l7p0wuq6Y5JFn
exmkQ4egO7RpcN7/uGMXAd93PxxE4K81S6BYWPcOwVuLFJ4qjZLroqwSWBV7yyjy
vjY3kS+05FVeaSrMADt60u3LteYx+OMdUYE4agB2w3kg/kMs/F1lQJVQH+0camc8
N8Vub3nIqORSzAyL9rf+OXYkkWhismKuTlt+BOjeqYspdPAKdUBggzrRKnjAh64Y
bXyEo4cRzsnDa4vzR7THh0zgK36JvfNCGAEzST6qosVS/0offLy6TVrJo2y4D4/R
AZ81msUgNTIx8Gb54rhjKEaTMDmhz1VDhwsUo7GgTBlcmK7wrLQYQG0vFjZUsbBI
qCqPWl14kuTI3WmHfa0fDvylS2tl9UYDewU8zsYdzfGrWxmG1Zvn3646TmMmmPrJ
r3TC8toV9j/RtiUkdpJdykREXpSx84MbHZN47fjJWFxy6rfkGZaAQoNFqDvCPY4s
IQle9m1vIXIjT0qMJPdxx95iX+s1ghp1r8s1KiYwbAg2Bnm0cmtF7gyL3yi1ej60
DNjwMWyDLVRzNDVsnLZCPtmoiSqmSc8VZRIFUiN9MOCD3WtchfRBlT8IkV1a/7Ac
Ethvt/89rES1GVk7jITdh3qLv3yp9mvFJ7NPbkFo98qRE3kf2/mmSEXV7Wdf0lot
w2Sc4NOsAPqZKCrvvogGSx366GRB3DU83DS3ETfXvedpk6uMZrztLwvl8IfZldrU
C8ZMBnFYBmGls8vOZi7LorL8BIyYGWNfa7ysNHcQtWCKEzoA12Nad8WXbT/YE9oY
SRVMuqGk0g+Zh1i/wu1FEzLeRTlSATgaDpWkEq4s9JDG72UDUhk78as+7Y29spsH
Yqg7CEd5rMBYR3YssGcfp+ckSWtacHjMYQWZdB9bW/s4QvgEdZ0ukKyIn9VqrIh2
tesgPvPchL9zQ5E2nIkG00THql1Bdqm/vmLS5BrX4H+JnXPXTmvBU8vccUhbuLZR
2OaCh3aAWc+ZpVdIwtbHRt9o3Xe/9isRaZznwuCZp7X2MuEGWxvWRwEk5dOz3cLD
HJZJGDLWnflyehz8Psf9z4eMXCwCpxssPuIOZ86TNhMq9zgiCgYK+l0LisRyUtNe
f4GUjPT34ZXFD6LU7WYg+I59axP1oaDa9MQJxo9c878Mbyw3PWDRoXReqzJzWZF6
Dn/CoASVXkNLI3M1zeSz9nrVvYm7TUrDME31JX7GXJraH1xrGKDSxiVz0f56o2pq
p/a52su4InpW5aBU6n3JEikRH/S/VVodWgnp8Rh/Tl/ddbP1T5Io7bweBOnQ2lS5
RV0+ErHVksmLV7XLzno13xTqxuTmVvccj3KRQpc+iZSZQV7QqlbajItb3UDQ10Hn
mWL/ionbA9nNtq7UbRguJqmKXdqHDbZlJcwhvJVqJxwRCIM7A+Mdvdp1iSRML27F
rwflxMJK2VVdMFmSK917RrDaBQhom7iO7vaFyzVjmqxneic/MbnqfPwRwx9s8od7
M2zsBBljJujesXPuWuALc2v0X3Etbc86meVO2cgU0yzSiO3IaLMTVDRjaUTI70I8
b1M4WM5P4Kwd+RcRWlRYIOyZz16JdkSjFrbOUtYVcNs+D+ZyQm6D5tO7oVWCvqK7
gAMGUtudVDU6GJUWIR//+z8365x1j4v5MoWaGf6emYx6g4ObCkyQnh+ZpSgnyeAA
OlOF04REkdReeGGDDQDN38CC2TqaIWf1KajmlxPj5E33hW4hY9t49/ZK9XpDsudy
E+WXq5QyhGPGU2gDNPGiX4HjFYr0KCOvxn9JQ7foe0CJUXWl933Kx/y0KHRUcqvR
FYIjywLmVnE5Gf+i8rPw+h7lMBP3l5UE/KkPZD9ndRuNQ/yTGvgseEDj8reRvyiq
hS55CkVSb+U3Z2mxniMnoXEheJercSXvlKulixFu6MOi0AjkkKq656M+LGVr5Q2y
mBnV/thbO7y5F7B1fztONvPSZ5WAZxSd2cuHnGdQ9VGNy2M/kEruEeW5UN64rxLX
1qMUeZfj83GwG4SQChQqFyNlChVTffWSVyEOk53PTwRf5Oy++JEO/694/7QjlrhV
xhaaBmpDdVvcn86QaSsqYGSyYGbWiw720tRpk4NaiLFumGoqgC0cVsh9JEF0XL+f
OMt/vDR3s8QNlW3fj8XcEJwjwmfRjspG2RTUDkELWch6fK21zdj1JbeboNbq68PV
5a37qDZ5M2lO2uAe/2BJYUfEKIhNuJ6mOqWNPRfE6vg9hW9nUv85nGTl/MWxY/zN
4ZaP8Jnia37zVhk8Ik3mkULpBPtoUvVkSXzZQBnmjrOBf9amVfYUwcT9I5Fh/WMD
rU6bfuQFJrnquO56yjBovmSxl+ssb8tltB4VSjsPvnd1ULAuJ3VEPDiUvyjINGZP
JhukbXNki+r+UzCed/ZaxHzOyFzGcabcYRQY8HqXFSSfHtz8+dF7mpYRkdsM7lXW
JKhfVdWtoUHLhG5HELDvX22ZFpMjcqcPWc39+p+O/l628twmaoJpYoYBOzH/s4/k
BDreKVrZDtYyL9E5R5oOl/Qr16jzYA1U47zH2II2iB4I0LqwAo2mOoUcC2tuKcCB
bMboZaYMPCcZuqHNSw+XYOJ+TC7yIcVgUgs1xe4kE3oIEhjWqksOogm9J4ApT6DN
rs3flRLkx6icjvOjM6XhuZXnK6pHYUi6qwb+mrcqRK9Nk4QXAQfy1nXqDtLuftzK
XHHkMEFcsHiTM6YzrB7NJGy00VugJmeCLSXZyN1c6+kMofQg5QhwORZVghZpP7EZ
FYdtEg9nilTZU0eq0xRJNv1F1gw64IaL23oBc0lGdfzTORkYUNnL8UqP8IKSbIuH
7W7ZybRKxgErr42QysZ/WwF/N45/5FSnYsL0mki8j2/l8iydppMlpDRJxyVaxnb6
ZWJtSDLuuwAG7Qwvf3EPIrthIM6HdBx0Xm+Wrr/TOmroPFuPuJlLTBrp2xlYIBvE
hxAx1FKq4QMgJHhjCTwnAwzExESz86zaufA1b+DcR6PZw92i3+mdZ99h/YS5+UQv
pvTb4ufkHOSugvFIM8Jpjq9TPHcTSsCRfzgzfiLZO4FC6rT9TGoiw+GovTopZnKE
IMNEjuEtpxqTETkJLJ9S0ZADObqLGLP7qOycT8W4w9MrQ2az8951soSI2bshhUOV
1MtC8Jhwe7Z0cfET9c0o+ER6G15XPdshCQadu8cf4Yh2qi1wdWFbq0wFuKevReJ8
MsLZP3dAhJgQGh6cG57mM3KX7ZR0uNlEd3jYoYkXxWKEP7SDfZHUulpDKrsdAgFs
thSXTspgMpFa5sLGSwf/O8XYwS7wqesccMyl9TX+QVE5BwBAr31FFJZR43LnX5Ne
pNNpyz2qdGl5EpUmhjqhsnNcF+wHZvdzSk7qdzr88ErlpN5IXxvmfUm2n5vBReyq
wclhCO4YgtSxWEOfQSn7CytkeepeseqYbbp5WOQAvWvU7hlZEWMmN8Rkrfm0sCoQ
5JMsgsuYgvzMKBWFfCh0xfIK7T8eB/ab8FmlG/u83uXn+59cUFDernu7SJDzBICf
jNQSvxnOZhtIBMABEnivDLmQWYQtkY49bbD4l9r2V6bomCvXOGSIBcM3B18RTXq1
OPoqilGaB6zdFt4NEpEwbQcESugqOpF6U3o5JDyRoz2oWOFqw4nhdn625i0jRG6z
eOy/ncEZ+rfdi+iOwtbm5vk3IFzv1UXcAUNrYe9Kq1zq2+AztfiLOkxQqaSl2QC8
X6LrMT5nrBu7s8c7/uyRwD0DDQ5Gz6A3TL73Rg+5A3aQQvdaDZZMWKo0pImg9/j+
lAhIPSTFxeOvDAQocgMJgM79zMAmEKz5O/0WXpnSCG9LcZuzaILWRhXJ8p1D9bu1
jSeOanXt62HP9l7yEydwwMfxTrXTHqPLd7jDEe7J/xIkxHyTNrOFwiVTEYBhjNtP
FEAKzdaEY27LUsGK0WO5/TZLY6FiYXAvb9QA3vbQY93dfDHK5fEiW9/Pj5qLijcT
OgTy+b7x36wMeomlmKQEzAfKHDBsc5leZGPDAjAxIY4wpMipyjgH1ZbA1/RZBBr5
Ha0qzsvXZTCaZ+qT4iz38ADrVKo6jIs9mZfaDOS+6HjAd7nM+FzAvh+qEVSRuuRm
gwF4mGjtzuYoChv6UG+Mv6w4j/hk8ol3QbswEC4EuBttH6dBnVt0wCgWX/J6WeLe
8P3MwSMN161rXNcvOUzL0E5/nrAcXiE7FIB58wG+3Uk76+YQkUAw3jASEqJYYZfJ
l0RYm2Jv+F3KY6acd39yqUMpF69DJamS7JK7NTp0jUppDHZNLOjmR7qAtLqNYyBD
Jk0YuViDQ1/h4tisF27apzMudA2GuTIAG79FoN7CKmXmoR3tTSsTUa9IqnX1gqdF
nKj3vJwuLclPx1y6AUTIC5TUA/8PacE/NXS1s9gsltRAIECLF5kBYmUYgH1RKsoV
juKJwz/bTWmNfn2qQCMAbaKih+QbttjPyOlr7Wx892qZ/XHuAA4vTjTSJZnVghHZ
T3XrigYj6OKSQ9KDHJZ2gbPhXf/5yrvUIybhyehH1oIA9M7/6CXaIoEVx0BhKOjD
XL8qaabYR27bMDwb2k6VPgzRUfPlIu/EbJqqPnCXBeWhaZBgAuf4cAWXRxTH7yhy
b+rWu5Mj7dxuVpvDpexbOfTsYhw+oUUFMY/gQfZ6dNoFOS6x988Pp1GbuvMaaknm
fQZWZq4KsQoWpp3uXA1uCXYeS/nOEFfASKmWkpJhM24rqjCiGXUxW06YWRraZWOQ
FQWYNO/9AGcVT8X8Pybo4tv3P+lQxlcO7fouUS1y4FuaB65AnY5vfjd9A3XO+lgX
DoH8VYuQ7wBCnl7us0bSrTbwAwwo/+YL4w33Xg+tyurO/P8owU+q0q5g81VYCuTa
pTMXTsASfhnlolTVx5TIKACaotx6E3Aif7IAJcqLDBusVxD/cTybkDW6yZggsuIa
YA3jZkE4NUba0KsNSajcRjiJAUesSFB4o/bMgepbwX0uxcwtOF49uRWUaB1DEHGV
KS4MqPbazUXEhxhHsw7gXsPMCq3K13Wh4ZmSLvhFwS3IuXcWvXHtDgR8u+sXMVPD
Jc9KzHTIFigovd/Xux9RtuJXeRbBIaEuPxU8QRB/tjkUqs7nKyw3Y0JcNFOJFIdX
Zm0fe1eGp+bCbRVulD7Z2FPXjumObLc6nlCy/mC3MTwLUxEvI/2I1qFeCQstsQ0z
Z5TxIgdfi6OOdlOGK8Jt1yhZ9VcYRP7NnZLlvfEVMi6PAhmmrP4HaaOO0/F/y2rK
wMwPVEdntApDH4I26WrPfHB+qc5j1HZ+Ig2zS+P4A9QjSTWaHqVgpYaNLn0SvKej
+8hSWq0a4Y/buV4TlMcg65PWmL5Fn0ZBP1jCz87th5RfOHQAnG5FIFrNbERwkgcG
Lx7NOlIMZS2x7kqig3nLgzQaRqyE+n2I573NhH174d7106aytHG0+wll0YTICXsM
YbRkqBm5JLIpW0zt0VdHpUMhyKpomObUv6htCq09HR2Mc1UA2Ry+YC7DJctqYRhJ
Bh7Ltj/MSpqjQKKr4LNerucIxYdNZ5edMzh3k39zEXTFfPhwVvNLLv0aJcq+NVQn
8VLxCDM0mWAATPj/47Mi0vgFZvypCWvY5MGd2gt7OBFCZnaGkUTFrJ9C+/8BSeq2
FgTmzKtWoxP2f6xQ6g/utSlg87BKJBSNskEZyFWQkbHr+dnrUdGb0SWsiMd8aMsW
cjsAHU4xHqoTjwJK8o20EJiP1c4SlPF1cBsZ51oSYzgp8B8pwpm1ztA+8JHHkBwB
evgkyT3YtplCbehHYiabXgmuBX/l48GYMp0GUgKfn4X6qL5dc2WoVmpRGTHWWgBN
ag0yOWkOtpHOQJoYfRlss4jfGulgZwQtKPcptWiDcjBER01C/stXcmzgqVVNQr78
mulhGTXe7Wf9qFDAVseZpbccbe4vThvmBGrS4mOhjJv5HmLwyviIWeHsEseaRDO4
KISdWJHGDCFf3u2teTz0LWL/Fktg0sAJbAnCVtz5Y4M5ohIz8SLMmkzcEe+QcZ+E
iJglOboyAadb2V7WJ9SfmgrfjQFk38K+FVVTGml1JSqOR3/DZLwH4fHcLcD9kMAT
jk+DhjBQLePqaOLn/5ylbKGivtqnsg9rMjYbok6x+nMbMtDfdH+n5lg5SG51CjrC
nRRjb7bI0fbtZz3a4PcmqGXMG2DvcL2d2D7BzOJgSBPzMs7wOVN88KOhOYPwcHiv
zvQuHAiuYW5raMxwVUg4eXMWKmYUtmdcXW+KkT9zyaNJd7ffcc9TitXhcwfVRiNa
Na6SwmT67D6YMTYlCev9dg05CVc8uOivn5pvJCdiQ3f3+4iDW5UEXkPuzZZxU14J
9hXJQmrVaViB9wE/wrqQz7aimo9rlXkItWfkedkswpssZVD0WUMRhPirTwsPmsDf
uOe+CNujavSSMdFvT1OHV5HJmsjrY9/BTkiYzxflQVdOH48mqLxNTLCUoEte+5tp
16q3NRj2K4OwGX0TWsSWThbcMT6pdSb0PwFbALRLI4S4MUIf4aZzlT0uEOLJrlk/
E8aPKpue5GhnaPSSjAMiK6wXmOESzk2uQthc/M11yo9EwwqO1HmGUUqLux9B8pfq
rZsT0lncqml8h6AaDnrnp22TDUouC3EQ294Dowy2uBxzcsvYiShI84WN7yVUD1ZY
TwkosrDpRRH8QidGJfHoYg4LdxFJfJg8+sT02MfFZPUAXUHqKRVltylI7UH8xeJY
/PebUsWcyrBjCyxLEPzKS9RgpD8xOjyAkwKa77EpRgRu15VTsrLeq9e2bUKgufqo
Ih2XS0kFC8G2WDFu4Ilqf3d0EOOQS75D5b9Nf1OXJhNKtRQtZInjlY1+7IhLZJrc
tPbvHE2i/Xio3PFc/9iPtHHHD1EN8n0BXi2qOR5YbqoiFe4cYge6cEXMKk5IpjHh
ypCX0/HschMky5PScGpWWM/WrmPgXdbAC4wjvA4CnKtr1Jtp3v4tHkSIPHYqPQ+8
D+2gzSTgSoSep3Big39vsMePKKcsu2AOLmfmsA6aS1D13hCgbPBj2kpLl47A8dQr
gV8UXZ/2zVfD+GxyD6vwUfqEYseSf7NPETJM1mpIPhXcF06QQ0WbOIpmtjXSDhYX
Y2BQfkat6bqSXXX8yZ24NKHlK+AcvdvKPd98zhdsWWdkB76UixrrTOp6p6isP+ZY
LQI2AUF0KzAg0MfAmplAmvrkIu03ars3uZ4yhBmrtcY216ns80lE21XU7MxOn77w
Yx4GYRT1+qk1kH++OO6MO+96+jz5s/U1bC/+rXoTU7SOD2vgm6ivd7ya9BZws/Qo
4uqfqvzu7M27FCqf80qPfI+uXw0QHB4JARgh+i1TP7P2rkCrI41xF+NiVdV6vPo6
evh55olFTxoY1CDVTYuqAf/yCv4reQ78IgN8hE3/tbo17fPV7IuyMxA2JtvK1yp8
N4cx+Wt0mCs4986xoMlSQ5WxU8zPigZy5n7TMY09Vw7I97mM/ZaKquh8lul7zbEA
iw5spDskB/N0S4s1EumHgvzsGDfq0W7vb9hcdx3ujjnOPa7C4I7rDqPdFvuf7zkf
hDlhoYnId2VYDUC3j/c9jxXQZZg+VorucZyeu6s+gNlIgtzDVyWiTRs4NsdwYklQ
VzeWcvZKdaRGPpqPh5zr7UH5MqMnlJ3CindFQOJcZVLzmLwIvevmknNwHRctvBGX
NP2LOPJMLXWrK4zvDcAMPqf/EZpO+DWNtY7cVkDzeZlCWxxcNXuJXtZtTIOpaaGT
UtTSTQZTVvqPQZEijAIQFDKVyI/X/CaOKddiiU9AX+jXRbZB7VF32JGk39CcO0xF
wQs0y+CK/D+xH9opxj2KZ5O5/IH0eWaWi1ooqSCBEizlgPq4bAVZQ5xmpal3lTnO
j+PZ8Z/XDbgcdAIc6G0VmGFxu51K2/IN22e4QJoFM0hovc/uVb8dgN5SlzoYLLlS
O/9wCB7WP4B9YqitIIyom0LK9w5/Fq5Z5LVuU8NAoKeYRWKuzOkXkaIQsr3lK1Sx
qUgP/lJc+iibDOgN9IBGgNnO+ZHEcjGFbLyGlo0Y8J4XHape4DrNk7u6IgUTHsXD
IXLg/4hprta7kODmx86rghQZD7vTZvAGjuNapnqYUWk6cxAUmZf0dfyjUwA5nzU2
9rXRdHU1nGvCL8bC7OXgujPzu4nGAsCZOHMIT8nBfYicpXAaum6EoDBqMpY3kOK8
/dAGlk2iDWb/LmUdJCGfmipzS1ZShuIVuNx16psvoANh7OdnYy+1GNNOyXxy6v1K
Flwrecq7mbCC5w6T4F27hLAhbPJWYazpAEU7tHM6LWGw4kyYZ6WvBJGTo/Bw7rP5
91nQR+cQNiZPsPZERI+i0LIgGsbJycHr1+q5YCst3j8ZLxOmmE5DBESyea4+SJ0q
4zssHrO7m6hyexwwZJWwQPal3Wf8xq/KAJfnnqnfY3kCI0LYbr4TzTrRKGJjhKk8
2ijpsLSv8nCRbsFbcloJ1yzsdHhzHmIyTRbP1I6vVaLy7U4k7yPUn5qekxYjV7M4
/Px342qaW8j1k3Cen4dVieAawwllRFmJyKvquo8ikzt3TR/d844tPcPi+6CVTrYW
1ro7YHNaCutEImdglAaeN0/oPe45N8KaAzLzhQ+bCCeD44Ab8KzFq2VWEfqTi01j
KtM4jN95s6JMQUd1L3L0VKbFsIyIQNHmu8yncsamvjaGOZx+lgBCk1jq9w88/ZNR
UGRTDxdTr8hYMNdKxZZHKRHE1OhMLrQje+GLvkrmuuXMGgVJkKw7UVo+YHY7EZ1O
6Wt57LDZwR4xXVkq5LCoNRzvBV5mgVwM6kUNaRSKNdErAGECpXtt/Ephh/xBvkvf
sIjivzK1CM2ciDbxVNOUKpDVkOHwB+w0QcWnI7sSFhi5zbWy/AIxMXJMmXHdfB8r
xi1OXYYsb1l8vX3RiUtsvtYeVBRBY2E1Y6ykIcS6oM8scYWLzfVfz04eZkS79DyZ
+hRJEOBqnwXfpQzKBfygSeXG1/XOdRG3oOFRV/fRDAPxgDJ+vOItcerAOmJZF9G2
TWIffoyyOWzP2AbhQP8XZGIlKQU2aWYaz9gz3EnzfQRmZLu5CfhQi8w0KznoByib
gmrLlnc78tXLLMMd3dICLvPI4DNeAg5vRRU32v7i/TDB/wzcGXD1WO4A14Y1kA/R
qhZ20m+bMxWMJv1w1uKp1NFsPjIhr4RAl5m03wzP4GTQ93nLY20OFc2OmBY+5pb2
QI6vjJCfjVqz8eN4msGq/+Lgm8hubAliwlETEHPE6hOoMR7bwiTxtbCUqSa5MgiP
YPz4ILO9Vxl70Go79882J5u3QdYhtceBPXRes373fYCC9YM9rVbrWHjeD3TSfPpD
99ajPNn9s9Omi6M4iG7HRecyJI/1IHdqIyLWPRcegh+FCjRiS8FcmOw3OQb4q96W
7GGU1T2Aase/dAbwgvhxRYPZyoBTQ+o+vEy48+XLkd4wzbn2JmKco5BSO41XjtKo
wZIARXSeiJoM2uoSty5/aIYWPdDofHGYJWdCNH4gZLf2y1VWEtDpH2oAbLWTt5LD
7TJn95QQ1D7juEQGUC6phGty1nDolQjcDAgMZ9SQdHDGwCjp/wIMm5CxBbbTWP8M
G6Kq36MD1Nn53xuYcS6yfLv3502zQWmiLwamtTH+6mrlfoqZy8n1gZjXiN3Qu043
tvXzslnIHji/ZiNoBhi+9LhM0OkdaBEPgO1Yak23Y0+kqtEan//ghOKDMfewj9lJ
InugYRfZpP1pJH1YNufhEccguoa2Pj/Bax5MOXna26m6AsEHGq9t6FT9fqbR8dDV
Hj9jqH7BwzO3ZcJozvygcAbaYYFTJBCYShYOJYNTne1YQkN4mcb9ng+MqAC4iWpT
cCA22UccApGU+64TXdxIC3RSvbLq1bMDCGhsjseKZmFqEWInIwtc6/lQ2TNVmggJ
HHjMngibmw0IXoCVUpTv4zm6KYQO6LXelpTbQ/apD3Ggs6wZ12+KDa14BAuPPYaW
KdYcKUYlhml05FGzQH6345BVrYjwcjP+r6Y9PJJKeQC6DOI5hATzeY/q4WsRfGpM
mFCu8QIFO6RNdrMF4c4uvkS9G5+xhvIX8mj9A7r9mbplk/Lzwv58+6e05ZXI1thu
Y/qNGDfeo9tB9QWAGgGC04uX9XCgXjSXoJ0OZ+xfc++W67xfl1cZRZykHTc1t7Ft
AhZbrJLLP9Xcn1knsyZJzUMsVAbxoYaX0YJxOlzZM0l+/hhuyAtBS3/W6xvSPHSD
wNIILiD6a57GmDhjrFO0uRMn3kyFUjyauyV3Po/c29qkBfJ/76ZBQXsVQEnGp0cr
SmW4H5kuKElYsX1/MQ50yzeXXhGy2LTLa/2D4VCoy2hAGEyLpwEc8j4DIuHtmuK2
Dm0MUbVHh72p+N0FmbLkCAwsmwcNRZtiv2jjc5yU6DbsK/oIMcjX4KothaEXsXJF
U281LGVnwTft42O4+RRF09QSZtdSxhC8d6ilXhCqIf1HNPmC+ueN1JTG9KVxTE3r
aoQ3ZaBT6XGMINdFbcKW00DEv9gVV+WTOjBoXody/if3CRxWgUORpVOXY9LZz6mX
bma1QsKnN01hD1vSXrziPM+jpjqMlgGOtj160tb7EaSOjNNKOVP6PbodyqNS9bDT
yIcvwym8qBM+ULwmgIEz2yN0gwiapWgJ1sJHGHbx7GnEx3GEjE4q2gnm4VzlPcbR
mhwLVSKbmQDeoAjSLduCQas5w9W4VvmrndVvlE5b9qkP/UnyvVQCVW/6lQTvKcOG
nrU+3ac1yI/5wZ6ymi42AnpauBO4IOQWp5ybi9IEIXhQ/FO4fK6tjf+l8BNTDiaA
vJxPO20E6jxYAj1C3a/J4LQndntCAkUQCUEgHD8jbV9h7YV1vTX8GLE3yaTHg+MZ
I/5+LmwmxvEGzkqicMWHe0H9yiefOipFMN+28L4hizJ26nlYOUOqrKR2Ey9ZKvao
fEynB7NUFotDdtU/FtVJzb0BVv42NJFCycWeVahVs1ISt8nxAp7BBN472NfDTCh4
9+wzqe4c6JfjHkBJlpPGph/UyisKK4jeyq0Smqg11rWdnG4lseSBXZsqHm+0u0Wa
vD3M+G1Cpg5KyI4K006hgJ1Ik0B4t6sZeQ9037JBBeNFEASvObOtGbkmSOeaJw7I
JeTYLEI4N3vvna6gleOwFQjEBeuSW0rm6hwq/wqJEonb4gRJD595xEHVc5htv8yQ
K7QPatkqahLrkl9tO55VmvEOhThTkOwplH5CgqUt8CvNpMao45zBrrzVXZi+EWSK
hJ34SBIrkNQL2Rzlf9V1f6P2mxuuVcElfNO3KN6IPdfDJk8gyVn+gkAddKmArtjZ
5RZtsTjOBjBZZ7b0VY9veL9yzxX0T+ZNGPRSX9mebZqjzw3uQpmSBtBsKIB4ipu0
RcoO9EQFLtj61H6g/FoYwIg0nhqvSDPgIc+cGDMDgAbfKw53LRnxzYBK2XHVis4H
CsmUpsdFKCzG3w0T/MHUynBSwgQzNTlROMdveQ6WwH0Rdw2hRLfrUxylU9SrLwAN
094yC6+GEdZxV0WIPYJOntokFXx+mkAbxamWhI3h9DF8RpxRu8vrzvxX+ksGyanr
5HToZMZc6e6Au8UexkNqrpIpgN5bW3TsuEeK0cRNU+jBf6PjuUNe51l/BTBy8fP0
Xq+EtfwHntM+BinAJJk6erGJ0+H7Y5MoHbKM1PW6AcmxEuXuzaZACWH1fjSRKZ/C
Gc4QDjs9VGgA/QFzLPGlWASVt03bwzxu9qBsuidkS8D11Ko2uQ2s3LAP6nyoD8LN
NLyCFAZBG1Th1PeJN/pnH/aIgnJIaDE8Z/nERySnZjkHfOd6PeT0a2dokMvuOLVn
3YYiYkSGMtcTeOvsnZ9e+/QPTzr1sGadTqZ6w5SwqJv0MEXRXKC4WkkZro4URJJk
zNtBhTQ0OuDeVGvJDcVhldUr6Jz0FvVEEm3X7RTu4IgF2lyisTOWiXF8WIH78YVd
1CCkuNNIwKlM6Iiewr/63CMvo2QW65+QDUSW+fv+ldhwlvYJ9eHtrh8ql0nghwjG
GDSSh6yFrveFXud8AOfo0izHf+Mr/aoylCaM3ZB4lm8CQtPAYEG1EtlTI8I8NYHG
TELgXl6yZQ+YZp3WXyFJg4ggovGV5WU7iw21mrk6o3aOfeYJJr+6gtj1lGZbbRyD
oA57SXiYwkW1ymDNblwYLrJ0XFCOuwhNoH52rz8VKlW3e2MJWweGbHU++u23oM1w
efJVu1w5t1LOQJPigZ0W2XQjNpRuVJBkRAGJ/s/Bi/FUCNdpiBcDNqn/P/We1jbD
ipa4BUj8VDwRR+lvG/9al0ykGUyFj4+gQ/llfzZP4NcC42bCv7oyE2PZSvJEZ04J
A4AnOo/Y4WiYwPHufBGnbfvefMkVDER310VeUY3PYGAyaaZ1cZZNIYp7mbE7SYV6
4pRf/Yi28HY+FSq1ZcfMHJh+LQkOZVMmuroAxdET47neHj5exfa1XecoxeX88Xfb
72vKOqNZCZjs5i+bQrx6IkAy0jJ3PVquJIJdglRw4CO9kdnelwp/qrd9fqSI+QOp
3fx0AgGemAqfs6WxiENeww0l8cAQpzZWFDS0aEe+mfOqt0W8vYTcmXRHdveFcn9u
2ZhXiUQbXRgwpvCtkYYpc0VzHBUNDf2fvFf5XcSb6ok5mWYIU6VAIQuuof88gwjf
RlZovR7I1fDEGT51qF1SpBtAd2M4H7Hp9A5R2mYI+pcv2gnp1xXvjE418cXvzyZq
SASn/RdvI0zvF6x2Xoqw9IpL6x+nyLACe+7R+GoLhYTsIf3SkTIksW0wemFBMbxV
4xLp6EMylfTeKGs+LrNB2EJc+W95obORStIGUHLjtn2Y0sH+p5QbXxU2NpQzUP36
OB3URdZq4Ty7zWYt0Vgn6eu3cyojHpF8EUnCaAROZ5YwF5FJO8MXf5ZF349G/OcV
wD4HMYePBmRhCD9hQh10Nv4OO/tjtUSfPfP+bY3HSGTDY7ZMiEoUklIBUgj+Fahw
wckCybhEBR+OF9QZGwfDbFPPsVj/j1xBCDGxZ0WquaKKviegSz6TikZ3PQyAx5h5
ZLS26VB9uiKIyH81+2RGnpDqpic01yPVEjg/Tms7mMuUMr1sh1E5TaLAHypvlpvO
tguqXsTlonQvYzcXJ1AHSJc7QRtnxBQbXScihEByhaPqkA94o/p1+Bj3XUboz/bM
4q0G6akuZ5fnziOqyQo5Lg70JXssudurEDN1esWWlkaUcAlGx6L3RjURww39Mb2d
Dmv359Me5ktn8S0IijSKikaDgwWSYAjkR02nJ1VPE+b+8jGNeZl9Sy849QHKm0DE
kQpxnn0GE7Mg8AOu0L41TdOjWm0C/SvJHGgREf8B4Zc0mVy1+7tIn6J49pWRb5L9
TKniOA67JdZ3VKirBrwI3jEtrsxMQgo7jkY1PMGuRCLskInzwrix+vOkeQRyLki1
aAaBqZXCq1NFiUAWR6YXB8ZdsP3FuLwIsc51HWYmH+uDJ4RQqWjX3wwsViFCDWtz
2ITNzqkck2oOXu1dB0NS92etD1vhSpRt9v2Kt/sfqW/GTXWdWgd2MhUfE8ink1Uc
yDjLgXwKAqIva/VnlSTABoAbGUQQVPCzuVh7YAzm8SpTLSJCDsub76N4QXnOqGUm
yv4TBF5ZSZ4qzfyevKSWeTRPWos24lrRAMk/IrPHlSZUtGHhEuOLuKRvSfv/XJLk
mgFukfdDCNMa9JD3mDoLXjP8N/jYzdNqfNuXv2yIBlrUefSj6E0VCRMBureHR5/0
oT3zuzbKQLvRAACzvmlXj3DngpTO3n/HVeJi5geag3PH34G2UKPefecRfgeLOnaa
s0qGTdgLkiA+6+dZMJZegQTpM6w6piPD3XPguuFhv7dhH+UGC99pBrJv30LD8y1f
RpX+bH1gR9HN+znQc773tPI9zNd9Cs1t9akCsq+VF/1e3zzepoKfI4+E+bLnDj6b
UNIp+TfDI4HZ4LQA2CVRgXhUrD2te3CaFVluxM4VUXF8tjAUT4d/jhQxtlf/uLyN
Txx6WeGbdHTs6E9JLeXijwOG3HeYo4lvdRj3090R1gFe0LhYno1UPFuVDIwyMTKq
/MyHmldxzfqdjan9/qAshzwe+4n0Y8eyU52yiWDGyOCjypDp/JiZmOgyBAA+ljDD
/ZSotcE5TPjyJ//CUmp1WYsBgXo/PguRM78TMggnvcnL2IFDKar1ElSNxW2rhgnX
MVeW9wP4iVYwZ5Wp1t8GhNBEVjQcEmkwJWbdaaifmAibY5tvvNPBCrDfLIycNEQz
f3D0tOg6brse/qWKmND/nrzvv1JZXWkqM65GAbTkH/qq1Kgmdpk11dyrOY0Y2M7G
Hd8EvN7NAsq3hB90itPcmRlSFUw5g8ZAqgKL7pPo/Kvcdd6twyFITwUfgh+zcSbp
fjRTydtS8QbjR0xNBLU/rfV4oS0ssBED9W7d5RYIxLi2/qtDPCrrv0jNmVGjlrgw
ydFWYED7IKaHG7dVaEdayPJ5tqFGRNq/KPiE6LaSVZm1o0lplG80TcFukdZXLjBJ
Lyjmmd6TKI2D70T370eW3eTkwwkwa8r1/DOur2rPUsceViI/p5TGE7PCHiMA83TB
7Cx73ahi8UwjnWbQcu4bAIhi+2WX9oBdt+1aTIJr6Lf/GpKLs3QUs7/TXbbWNLTa
D2xSsSXAZLvMV+teH+RMoHKXujpPfKVob5+6plW/ekQcbzjU9NeY9O7k6ebWSR6K
4FGw7pAYoHAiioNZkIyXofswXApUK2x+Kf835+Ihhj1FIcRUdpvaswZ6aCgiwrt3
U86xBPruc4tEQpflBTmR3m39FiLRQ4x229B8f3rSN/31wyvoVajX3TZ9uEN9RVrL
nFYLKYBOGjQnh3kC1Thr7tP0tptb4dft5wpcAV+EYwAo99c0EaW2YR4quATcpdj5
bciSLYQzHiZ1Z6ZotYERKOAmqjou0Dm2ISpNCTw9lz1Fj3lsqbCamLjDaDnBUkC5
gqqkqnfx8zO3cmvW0gFNBGVkQtd1AiKkIQsy4uMVqLWxNwDO2mDEVSRfouKgSDXp
Aef6lyuTzYnfS377IV/O/sPDPL2re5YWaMTQnGBfC+nXcNf0r1TCuMN3Awe8rMGn
fbRMbX2NHKLxC4NjCuyxuuZZbESor+wz9ocfekzbMfhzV7wC2Hu5BRJG6JUVan5y
atHV21UYUlgbDLGU8qRC0jmMxqJlJq/R9MbObBO2GhSSrqizEmdML9+WlE8VRQU8
iftv85GdSR0nWa9lr9IkoXYSnwWTYefCgJ5XIuEJ5ve5owjU783CKbcC/zchnyFJ
zsH3P1MueeyFgvaIZ0DrLQt/cMu9aJdBSN1i6nrXZcLdUdnTqpRCXNA4COMMxllH
1RfgIOnAyh/kxZNzaE9+SHLHzVi5RrmRWrHHbxQHesxAk06mAMSiZXcynyrPUlry
GqbUXBBJoA54ej9QhuXgBGsKjup+JG3kGBRvvPC/Y5zCWJ+cSHoCgb+dZtTgaC2Y
V84P4fFqpMS0B65g4LOE8uucA1mhZGCKjFTD3kfBG/ybsoFU91dFCLt1nxKxg7xB
fom6aGFIP3P7dWDZDK57McE9YrPU/kS+SsLhPxqhM4DrX2GTNsXsisuIs6izm3xh
64LhIEdhk0zdqKWTXZtixZqTBpVyhDZ5HjkX0lJPeYDHKyyjfqJfCSfpSvQYzyKm
j3gDqio3Aq+yZboHn29Obdx+Fia6pdV8tCNV4xqW+v3aVOEUDMeKzLwDhHPaIwhm
XmLn7RaKqz/7Es5w70AyvyEKcZh2zV5iukNtUT4a26ePVRReiXFb6nEqfH5CzMfC
h1JnAMulch3T91lUXSC2ZFRTG3Bo5MSBg7DRHslmOTEdp8NskX0JMF4DwUW6pGe/
eznB2oO10ASY6uVBjnUwnQfWwsNr4sPcqH+lgZml8AaXo1weFs0ib2cOYxIEtVPv
hNujgHyLd77RbdwEYeJUwnwL+vlNlHkAhm9LcVg5gfEVprE/KGxjvaoQ0sfj9YYB
KDPnR1j7tGvd0JwV7Hbq5hF9m873jvAONSEnuoJ1gdA91ddKUdpwfZZcXvifAYL6
iqvqSU5CHgFwy3dXuqXGLXAlE7pQrNWs8kslPR6ez5q6g19Y3GOIlomEWtiQJQB7
3ZDXgc0jgM6OLGtBBhCXhGd3FBbhtIYQEGVYxUoIWfkYxjroOfGcDXSGS0Phwfz8
PTAsS0T8XZSaVinr9R19up5FcOt+1A5aPPj2ViP9riTgzow1s3cNgweCRR4v+qiB
uFD1BQ3KvNfCWEcn+mVqUb0RmkmyWCU4RCT8LPUq1fAbLHuFussneQcPs4yl5qXA
QanOVB6hsIWW11zu93I4DIDvRnes0xIwfOZG1rzHSrMxB2Hb2lc88+ggNyTXAqOA
gyQtA7atW7Ff7pzEopNlR9VRJPwWzv8xwdoykSFrZK0JxpMjMok21vja2+4aOl7v
hsZfdzG9zcXcASvW00HF4+4JTEgIjCF1vRG/bM/7PfXJwoy8pqW12OjU3DHx+KeX
yHygWigsEDHyIxpjXL8Sx9Jnfw6V2lS9ghccro4HE6/iTidapZYXoClHsG+J6txr
J313H6UEQ1dMpiPurXbXEq2PirhGhH7m8Nx4dehKLoP67lIbq/iNMWWmpQsbAIkR
hL8MYoiVXFOEfWC6myttrznuB6RinhstsESHPzVy95wqe06vwac1ecFiTOMoUiBq
g/3BwjNmFacyElxNXgksWsrfvfEOt0mtY4yo9ACRtQbT5RXx/NjGBoLDBIr7JIcc
o6tN5ZM93RMYHS61qDXW4mjEzLqozsknV1pKZz4Hjk5UKEnuSQe55t1zdWgw/Ofp
PMuonfOFTMDfzwTJtb0H9lXTQMDB6hbGn1HuqRPA8thCkJC3LubLwXv1WUG+VclL
ozE8oCWCcBxyeOUh1nBnzLFF7nBDjrj4U913LMWt08285UXEZQ3bihFIplr0hpI9
Az3jy8tJE690gi/IeLxdNatUnYFKjB94gf0hX9UBMJ3l4LQI32sjKmTcrC31dCjN
AXCpUd+YlkfEy/Vzojj7999tLuas1bLs+FdKDwTv+lcV4Oj7cMXeDVUx43Czl8QV
7Jfut+dCV2eUrwSA5peXN1lorRhsDzJS7OcYPWryzU/awcH2SWJ/ENkcT2vlQfXr
qz1t6t/EdA26CSVgQJE4SG7L9hPYoMl8uw33h4j0VAwkt0q34c026Wyc6Wcl+V8n
16c5Yw6tZilTEiPSMjWmuDtd1iHsilFRry0Fx8Jpe99qQ7k118SZ53Ol9TBsXOpn
xMiZldaHfa4MELBOcitHLcFcS9U+PwzZL4fYVtosF5KVQYZQ1E1yyMGcM8nhp+bE
2ZGO6jwHeqUE1oJw//SrRW5c+qGr5oZnsAXEtK7j8K995tjn2nWdxxDJTHfzOjky
yrd7ZMgsZpkq9UrzoD6OQWounUq9p74hbFQ0z94m6lEYE61cwrZRqmfhYqAc3ZH9
7ZEnoiWjXZQa/hGiGdTsNrwsWnK3M4uRIZ/0kdVCHYVXaGWkeAyO6bzPX54+lh4p
rs9guVlsVQHYCzc0C9KbFTIcRSozxwsSp6h0dCZK4Eb7zK5dWIR9XizxDQokTnPx
f/vEL6HYjc4GoUVYCOvC5wITVyJrssN91Tgz1nyaYbhEVW22VGK+yWkTnb2pECQb
71zr/pdVbLoHUMzTZBFgIl0JyVtyWVDeTPQlq4BzU72oXLBb2eEZUHXDG+W9W67V
v1OeP31Q7cl8RntVwBNESsr5SrMoEYWYDc7rg7hqWYiJJg2B/i3LyhhGjt71FSAn
NLa24Tb24iB/nQla0YCtg7QRuhoQPuSLRVy/qD4vteW/GAvA0HEAFiSjbjmuWLsJ
rP5a23QxcMDZ4+5XiSM+bIqcZuRVLhnRxNrV1N52KpTeLn6dNa5eDPbmUl03cYxw
PvLkxbaGjFdeEBv38fRpN+c5PkEEAYYh66LOKrvN/ZJ3/pvRHSGDqN2s1bPhDWgt
SO/KRp1CooHyVxvTAQKrCSv+AjGxeOy19DqWkM6PL+kQfOmq1zq+O/ZEHmGLpLqY
EgWjuegc1YrDfVJhwNk97nOb6P3POSNCXXNTd7YlCmj/lU0v6HVT8vkdr89PJwaG
S0O3jMohJ/jR3SkZvSQ9WvgcJTrheSsIuPw88rFE2Nzv1fLeqgcdqNgzA9//Cfzk
ZRjkZEb7xjmEuBKsASNuNWbo0W+pYQFl4gB0sZqz4RlmCRcyZY+YES6l6M89ZjWk
2KH8yJyte4UFQ1KHiQzF7+1Mtz5wb/IMaNwcDGIPU80BzkKhe7axKlDDMNxcanr+
wfiJEMHBkq5dVzwSepDSEwqqUscJWl3s+f+xXhc4QKAdiSNojZ6ZB/UY0rB4bNgd
dLGmgMCyb4KTFmE7HGAu8kbUR0vjNi5RjK1uQZEBTSxkucTBnayzXQRahZjMVo8J
YNAn5UHDkOyOZr6UQzaxG37CkY3Ai5Yt6Gms9kCpYRq0wBTUFIP8F5uzFbh95WwQ
gQ63H65VXEvgMhktXDsGKM9CWE2tyXcQRGa6VWLbeRhov3qEJi4XWGpi/AF434jX
v7dbIbylLt1jaY90HLxqgTt/n5AkdO7u8M019rx+dPkkNt+PNGC6XCCopO6ecF5f
qicnPyPCHkg7cFQMQOmkbUD5A8zzF4+dPbKQZVWJRT3hV1XXPVF0hRV4U4f/riJI
mjtzRhDX53V1BChGQjo1QkfPtNgGM48kLI5DtpYoa5F3P7pTpqrRbsKuZMfWI+l8
3DO91VxWwo8gvlik2Bs+JIhM0/njlV4t27kaptjVoaFeXnXBU9fodeRNnhDxEQUR
Cn8Gsulx7k7GidppkqpZqbAtPvW3puMbsHjIjpfmK752hUNPZmkfDrHpc9Uzrebw
8BG6EW7IcNI4krOPc9F0hiIwLQG5vVhNvzN4h0Bz7PKHNOaP46b7+/1zn0wdkk6T
ckaC6LrsYFh+gVUoPEt5V6ZXtRgjJUP68DHk6UqwpWKiW5ZwZMg6+aoSjEms/bCE
gs5pdn7dHfD7eVOK2vVuHs1xHW94ZIfVFHMAXsm3c71jRdWDVa0mB9fyE5uXW9Yn
ZpSeJs2qK4539bSUxT1addnRzOy0OPPNRvlC0NymQhRNtFxt4Z2HARMxr0ffAepj
ZpkoJqy2B7rtcMkdJdxcWnf5i6tE+NGlCAtQa/VNWGpC53nK/pkBjHzVKz32M9ao
PtNQpfgMBNgd/WMWy24pOeZ9tOAllOGS0AOjFJxCYXZqJ2Q4lmcdXxtS3I02doDe
HUFylDuMwIDtYQSllRcuXEmWuUF+Jk1vHgKUoWZFZ8HjpJns2Cg6AjogfKyC50rM
qiXAPh1uHQ6Z3MO6siVVjtNZTtelYBjPFVXDBiGh3HGaX6pcvmAzu8IDU77MrpII
7Qh+6Nb6maKW5qQOtA8PLOEGJBjXWAtJvmgh/VM+T6MhnAHn1Sh5nhS2+RC1q/Ze
WB9AM5yOLJ4fsrLe9I0Pivl3HjkG1/KoJwJut3KBjh+j0r0Z02y1G6mePGWJPKWg
t76vcvYmUa0T4jMBmiVM8mhm43gVa+MQYsuhavZ/OAGbdppogNTrTX7ME2oLe98U
fBSQZyXSNYf5Z2iEUtMhOpAVWZmewt+gSF2lHvBJV40bTrlTEF0n0GrJ4d/HjGFw
qvQotBTumqbfHUa3nCKphgp5h8pQu9eK+CGcKN95uKj7xeR2hI3F0lRxO+N+cXcF
Txvs15SexsFNAkL51UtijboSgW4x113nz8NXbDwxP5GTzveFiM1p0vUNNn3Rf327
LIjgQSjz3FnQ3ForDGmP6HyHf/F40S515ezIbOlZHLxVum730X61kh++PmKBy0YT
OlFau4SzrqrxtQmKqm3EOvvtx/66A3Yv2c+pW+q9DX0hGlJ6AekYqzUUfV3HyWWG
Nt5m6icjDrYscNyrYNBG6bVWhblUkNHyZAnuaODg+sHSdYgKEpGsH0iDbO+5ai87
v2kgOzukBqekFLU8fNejyAo5tHVnFXMsiKFQloGZucLUp5wjlqE+jF+gREKBFViL
9QSWA/6XVDa8jbCLfT/iY2oJ/QJOUhW8ROfR6hDuxINJgPzescgFfPXOrBx9ZbvD
8S53ix5sxhEnFvcEbu0MstTKoN1LKKOJMh22ugJv5B1p81m++JTho0RtGTOJPn15
OPNpOyCm2xTZoXw7smGxXx/W71LZNerMWSlBLCxlY7z38lgCwq8fBRb1gXBF0HNS
atSvdPpC6y7TJ01Tud4/h5qzu73sHeG6MOyoPu97T+JJElj5ksxSA0hl5P5f85Cs
huIKQaUMa2jlBRV6gEixTO/LWI3WvQVuWPQY90gbV7CUeSb5xLKgkT6vHxwDm/VG
Npjd0vnDDFsrV3AeGNKFerfTzq6WFUVNTPp2OljR0phw6PNQMRJvOQqVSLFuqavk
C/3XOJ4jpmuesrWac1ZjzMiDz6yQYm8nvb6Y94kr4ndbVAF0kAbdtb5DpERoTvli
fjVxrL16dA5+NfdSGJZlAOwEORz6DIfu7QG5XFo7pQI3iUAm2hWxfj1QrI2oq6HY
c6iWAgMwNe+FT3pq3m/2lMtcb0FCp2sC1EyVJ2LcMAFKps26+Rs1MG1zSgmCMOcQ
hIGkspdEK+K5afeQgEIPrlxrKyowDrH1PZkeOa0TXLbuX2jyTfTfkk+4+cUGwpAK
MKDCbGoZeuWbVuj+P+YTHoT0FBf+y9+Ek/PILqm3AvNTioy5E5igr2oRVANbmwuh
Xc3124iJPJmc6bXfPSug02iKFgxVETeXYe1WxcGfc1eMxLimYy79+/EKrlOsslZH
bw2J7mTYcbWvfdBxIjb8PFYEH9v7E/7BPnmdzuDCg7bB3anCjyrG0nNNm0sZHyRI
1UgdTh9UEyY/V8uJ8+cmDsbNq34gyKy5YxWeCqJnLWpQ5HnLv22eQ1kbtMF6cNxG
8v3sEenYdRykZ5mq5ZmRtF18RwNKzXt7TkxAzVzuG7GuA3qeN9epvnriexPNWWS4
XvaN/x0o7/SGk3/yEbgUpvoYJvmf8IevRlROhNAtZaSAVvHj2a6DyLhu0t5JBS/v
aOflezbhIrNd8c1NF+C3hsAUi5DtrsqknYqWVPnWczmNZfjs3B6IiVU4YvGLNGSz
wkoVFCn0o/scs5pcvi2pUH1jCgmoTKly4ykb9Yyn7biwjcPKZr7LfJW8fJLbQ2zw
o5x3tz9HILT271rXmrgI661vZrWM7Rg2vROadnW3QgJXoIZl2+remVA0cMrmx4yy
jE3aFs84G5JHmGQLRLpehfEsZnbRL1WYe4LF41trCxHVYUQvYzMOonBJF7bC5y5R
xlyU70IU0SO5PoGY1Pq7CVlfBk/0y97N5Z5YgmGVA5B3e+8LIU2WpI8/SPKRSPP4
DWhj+knZ63NjGJBi293GFezBg6sD0pXjiIZWzpyN5uzYPCGy5tocoGbCO005BA1I
HSUVR5lh4d3PhTK4hnJRTt+rRc2qsjSTmBwZzLdcnDYymM3pI7ZhKD7t9slynWka
JFKgf/trCwQyNMwRqxu4oOCFwaMRdLwNtvkbUNkSp4DFmwQbuPA23L413M5QfB4k
nMpskH7/vlipl9GaXws3kxdQpAhCuAZ/kij5IlSSTQOz7CDCUVGsYd6ghG1pec5h
4XFv1TM8pmubAM6KQIWcQHJEicLR2ZB7Zzjm75RhY4k3LBI1FzJ4XOXQx7/Gcy0P
WL0cT4823GQ2Xbr5xhNxhkXB2K21Ju65O1U04yDiqK7fMwnraF/ETBUU532r2p1O
4ZJOhqg4WTMSlBUrkbPBa9AfZIIQxw6AwpX8gWSQNOUA9D3t7wAJlZ0kz0xPxkzT
uJkonIPtgmGr0e20Ho06cdOnikZTQ4qHrvTQBUWf4WbpCdnc+6CGgSdLh4oXyi5r
8bgUV4q7dF0pIg+7hQM58ENFRjpSk6Bql/c/GFq4bAQRFO6Vf4D5LRmdR4BLOvdI
lYqw9kHXmd/50Un0CRpiHkqll+TPMa9B2htgo2e7l37VoCDTQZ7MVGOdBhd7+oeG
30EJ0P5IIe9KLaDe9Wj04UCTe1pKkR1g7za2yIGNqh3MgBXxQj6TrKNqhUHJg35Q
bjbIzcjQOMFWDWjIJAwxFeIHRtXhIEX/fTIUQ+eqyl+LRZslo7GdT0jeaX0KoKWG
ZT0J+UFW4p3VdFHrGEEegMVAHA5ZYu1lGBF0/twJ2V8vw8R31yrKy4eJ7Mlrb2ht
UyEr5nBa4OXa2w+dLmGeToJ6bBLyY56IAxcZAGKpJ1esNRLz0MgwEdTITa40D1E1
n2sBveScXsUOkY91B7+Svy8IiNquf+bGU6RbnzFLOqgJmV0rsTs7eW0lvA7ONVCv
EV7haNKjKwErSeBNL0vPodC4o7+mbjXWS72ssi/oG9s+rInB+J/Xjsq7vwxtTugr
+dGGFI030Hop3dlIR+b20QGhI48mmUFg7YUL4BQv5FOXkAGNz6CiXizIAitMqFcJ
iNgw3Kro71ZJQULgGu2dW2L7BOKxKDxwL8PPCIP0DgqRhREyngUIf+u2e+kwYh+L
YWJT70LZQYb+u0Jaw6TaTZ4MpA996kSrt+OhNSos/XX1eCMd3GVGsU2+FZslDmBV
xx5Jp0Az9gXN4etIaxMedItKhZXwoQuuqaRQxEBcImv1VWwgQZZXKAoMr+z7miOz
PVksOwRGcIzGC4xyaBQKWlV1ek6Ch+oHoAOrLvKzWhxmQ/Ju8jwCRn2VwRCcNrk0
ZSdhSyBkGmvx6kkDnbi/JDgddQuut88B4/axD5JcAyLLMWsQ6xZzRu/ShbnBHjWQ
ydRCZXLzLqAB6DrlxCkaIZZ5ZWwAza5vP3DXLPd0JRoD+r7C5uZqJtmMPTvabuU+
edxEZbhHXg6HfXYFy3iTtUsxj4O7QGGbs9nDKXDQipUjeNJAUo/ML3g1zkbNvm+K
lxZ95s3oxfA0eP9gSBg8JJTfowWbTc9Z3XRqO38ZueJ+SPQzmGkmZc5g3TdvdTN5
RtlfD0sldXDLrADhixja7tpi4IZ9W/JAdZg9npjbDJLFU6msg3aYibDH4ChRe0aP
1xjDhbOVyUvzeE5pNwBmboUgccYG5VbPIwElyNIfB1fdCSWto4Xldft5cKF2+du8
+vS8j/OJXQGLyMq5em0xLV8IN2k7XBsz9erBhRUFSSNVCMdxjOsVkqn8WFyckMXn
asf41NB2MAKmGFRPBZERBsfD7rjqjGnuiBP/gsyTNbd3BTPgidqW2UwTpZl0qO+y
M/9tox/1yALn5cIlUxh/rf9zmc8Q0P7D/Sp3dOr6JpsMR4EzWKUChmYOs+OegBiH
4CurGuUkc+9CaPJ56sNLRjqEGO0aF89Z1oSOumzuy05k4Z90uAknKR0NIuveGMBw
JvQle1tQAVdZkrJqHdJ4BL5JYVGR5X/L7dYgY+n5YvPGSBbBAGx4pOzezqxN5/De
IwfTaerZUsMkWHQYD6uFSRj14fOeMsVhPyXWwXemmuXpUzE3HMf58x1iiXZQ9oBr
Jxydfn9WICGxwz4UeaWVUOvF98nH6bAnoVhibYz3J2RMqSOkH88/jdIBY4p/WrYQ
9AMDiUHXkF1Y0Pvk23ZIkr/+Tfr+gMG+6dr6ZrbAX5R7Cmzk5Oc5abysNgXSukQ9
Duc0cpl5C54rWUuWIinxqF/wBgsCsTqbB/c1zf7bJ/vUrgzuwYJn1mZz6H2lXaPe
JACYe/p6xAgJ6IPRujfJC3YTDoAXpRc1YZqSuDiXSpQprEnugv25mM2yFCqMj3ia
3Dw8RbI+3KmRyYb9nxTucKOQNMWDQF8NuF4n4hNwN8onCvi7vawM09sGFilPbdD2
zbPE2FGmiiYzr1jXYrY8hCxe1ayGEhkXg2EZ5Lt7JBsMNfGCH/WjlM3Dhw1P2tHm
sADsHnLtw9ypB2eZ/LZkb7cTRbAmdAbDKcuJ9mq1qdiGrUo+1vYX+aBAEuTiR/Uh
fifSiUWALaEb1lTvm7LOrTOJCTts6E+yGfW3TeK5BNU64CvnNbm4lCymiG2nsItT
DI0QCBd5iM3Z1hjsNjBST7oePT3c/6fQYN6x49H1uaNnTt4tUoQWGrWl031ijeEl
ZsGMMql+LUKxQoZsY9hojd+hN9n6oDRrN12y1iL5e7K1GXwxRDI6NonPpLNksTzI
37LrbaqpYGbY1LgaJ+N7KNiK8DKXyAY17rRMLLAS/gmLbSv1jmucLroldJ8r4tJV
dS1jOIKktJhkzom3dLeRlC85j4y+tM8owADmNRY+vU+/tmjOzJ6pq3c3X+BBS67O
W9EFM7ntYGVtADDNYSLFRJK+RHq/Mqex96L6UADiNwV4fgJg7lAu8gUTRC5vRqwp
D4xiDRli8oHDttLcPjNVrLWzav4txAZFeIVx2sN3u93ABDYDvvfoYQwPQGP8u2bV
IvWQA36Hpgot83v3SmyeitkUd5XddMEa7OTwYMJLZOyqK0GH6FsL/cFLzXWArV6d
K2bzvkM0v6QSULhgaRyJl6WNbVPW6XIXwxcH+OvZzI1Pv/CliBqga1slNxTZcxq0
phKIQtk5P0lNYfU5clgtNPt1wiooZe/qHK3GS4Ttc3IV2O39IHpUNI+bHJwxDz6S
cffAoMJXpoq3K/afd+kj0Psy8rRR/C/3vyM4VEeEvVp8VqBw77/T+mhQGXV9nkiv
r72pL4VKE7zxxJTlVmOgMekLTYajJhTg2zvLacVFQmrc9t9WNUvOcHHM/chPV0xM
HTsNMsnyrtSy0x0fnFz5V3jy+FaPVUUbcld8rNT6Tb5DPrzNHD1lqH9vAyZneCu/
i8mrqrFBrEJWJkbYgcrfqgTat5Fh+jZl6fXofujxxq0FO4q1QVF3WB1TXs6bI8mM
zXH3OALLUOh6sfZf/zYiW8zMrWcgtdn+v0GmOW0dQXkSZvYs1HKksR2iF0jzCuPq
QEkInXEVmEdUQhBex167oMAlpgpsxT2mnwvtGO0G0mm7s5IVTyGcG7adntxzDjDv
NqmpFbWssOx/PhOrWLM7cijrYmtqx/JkOMOhM9jHDR2hzq18feihj/nHqwBZhOeK
HhQcbi3/tgYm0KZNRYY0To1Al2KfuUmW2R0Bkzt4Dk0yz/qkbr+LD3G6UdZCLt86
wkawZViIviWFE+raG09E/MpFpjrtdL98/yO58ksEUIMHFAK56/UoALJ7b5eIdImX
fheOEF3LHYjV7ro7ZgnBOZyFdf71TfZ1kMLcxZY1bvekPy6QKHx2sl9PMaUpaB3F
PNeJD43r/S9nQODbcYwRqTJvSBK8YY/Y1hFSBQIKHpYnhJ7q+o5F7kZvSMDVq2qz
OipgkgbpmaNvYPwKezPY/uGWqxE1pLE+B4x/MlH59Wws+NtZt7rg1GOqInr+mXb+
uIs6TgjF5FQwTNZtDtKLe/qtTbZ8tmjtjbunjvvz4mrcMGv5lHx/8ZhdQcRBW2Vz
k+hszERqpha0l+tkzrkhATN+dQ9YNlHjVKswLej9X8CrfIasAB87mXz4/lkuDeYQ
etMfUNrhX9/IGGcZJxCOTqxht7+ZTH9j0DmPPw5gUTNHsjTGvdiWgl8nlXEY5Phm
91L2Drnpy5iebkFGpEqbovhvmS4B0K0Os4hBnVoHQC8HTygIkS2PvYItcYb5gqMD
445xzGYqaJyG3X54I1zfd39NpDOl8VDbZGFWbMNM0p4KErHgXc8gX+rpd6RZxBZd
6wXT9xXM5jRPANcGHI8zMo9gQSa06/JXdTZ5tAgvu0zSDYQuHmDBP2duCl+7mhBF
/aw52sQ1SFnm5AV4fTBva0uH1OMGwyP9TS1iGdeh12QDgasgllHNpRPaijSwE1sT
rjJ3WRDqfceVWoqK1khYDLU/GQyNFNAL77je1vXK5oR6GpzmQGIr3J+JfKjnh1Vg
/nac/L0O+R1kKmt6u4EGLK4elRvqfraC0/lKskoXuvlB52JKibQoguQKKPM6mU5U
1ytzB4+cwL2pdzSLP7JDOnIfbe2psVpa8inxiV6YBbpdTfiit40FwciyQEgDG8bT
FDyGqkEEcZiooyce4o3K8aVZE6phAKgkpc0ZdYT7eVjaZG9Z/KtXsZPRgGS87OYo
oLOxX/bxEoi+q/tBzf6vfwWgawJYiYKYXYo5y5r/K9zUpAPwOciLCefzKO1A2fv4
IgRS3gTOwMP0R9wi34h6vLZMWei8wNo7vMSR9LKLFFHZ+bLXj3/JvVMuhHNZDUge
BAm53cyF2Jxc+PKviAUJpjuzOws6ljO2mDH7J/RGXa+6iItQGxsykSq+xxyn7CAS
5twvN5z1hsybh9ASXlyRPqyRet2I84gJBCN/CHjOBq5kay9NJrlIkzeyljsPWtnr
toSJs5dIGojPwfZ8VcpisCc8lQngq1h98xjxmo+8v9vekmG96PNkyD1Hk9PcEd5R
5kJlC2NRUMr7hGE+a5j/fiE9FtYTzsOw8hlxSGDlsjur8nUZgQBRgxHafFgl9rJF
liM0nyRvVT36tTvV6FgDyEL5Yi+EkZ9fkfjiRxTzhmibRKxyS/uKARh7QjqZX57W
1whzTTL/s9xeNW5meBlZH3p7NtZVRnNsg/AmKwpvJfXr9Ye9R2imGiLiVZpW18BD
sxdYP5qO1pVFWCZeZqd/JURqbyL/UR9G51BKIWwWvaMS78k+zh8QZNrBk4MHuQU+
s7oliMr1acPYsHfIGVc+x40noKxq5fdn59d/HQhcRVHgm/nf27BCB9HkhUwgzpti
rWPnJPumlRZ93gJcGqXJaz49BVgitEdW4htL0xh8HYZovO/E+N6GHD9Ah4Z9ArXs
0kdSPpiZOGy4ReJFh1qUBM6K6OMX9iOG5Gq7xsxG7p90DmH3yqIHzWN888pat1qC
pm0sHQk1EFrbeHow4OgKkpefVmcpk3ay6ZcPQJKkmxDFtgRsO8SNhwyknn8d32av
PCV4DUmKkqyv1uI4vPQfIrjsuCV8brZVWuO5vhnfHCw9A1NavyqI01B4gW4UaDZf
1/7Gs5qlyByJLM5VMKiy0d8UsYiqJjAViwjCS3mE8Ig5DhsBBvSSvvehhVGnoTT3
O/E4TtdBL1x7zZmQ3AsZYRwfObjvyVCzXEUJ/0FXuFpTcnjWYKV8l8lonDAQFgXH
Jyq4r8SiexTzyalJHo4QAnDc5Nhf7/lSP+3IMOQ8FCSu2niL/bqinrdmA6PBuFzo
wyIRvHiyvNGJDWj8otyGRCO3u7722z+XHaefs3byQ6Yas1XQ1TcNQJ2pvCl141ye
CIs19Bj4lE6ll/RRAFrq0O4g5Wp5wj5FWAN4Y2+qPb5Hays/qjvTaOukfwk6PrUo
mmkxYjvqOY+4OHko1GzkyjtUTMinkIeCP0d2SoOZYETj+YQZBL78kscFZO3UPYmT
PasbfKX/19EmG8Ejw/yqFawTZ2K9sryGABKBCg30gGHx3veC7x76QQ+V+JFQLSis
qWquSKAoIcVmT+urTa1GX9NQhY0hwsl/2q4nH7jVjKJCKrX5w6BCI10+ncq5FtMo
UXElnUOnKJ3/gKu1v6KzJJ1o88caYkP1nldMylFEd9BT83s+fttzb9HlkRrh3mwj
cYpdG8y4V/Uh787l0FW3IoBzNNrl+9u5sMt6xEw7mPGdsFtWBI6PgE6nNpHL3qL3
bUArHa4k+GisTTefwClhQkcvQBMW3uOpRHYh3baMSPMWXyshqqyJg4KBD6+/XQZd
dv09UdhMYM36RY5SlU5JKGmDCLKj9nWKisXx+ptiDVWeA752NKUeHz30j8ggfoLy
wcFRFfZ0FoWknPojDvGTyJfsQqx22dRIiizVsxI7PemTQSYKmZKKb5OQQQ98OVe8
k+xeyBmPPHz//GFhwaT2uoAJ3TtI4sXJmG/ZpofEcKmmdAgXOmYGDoD797HhY6O5
Z+8HwGbterBQwK/dpOSRJeRpMCr6Sk4078oAB+svjSdBa7Uu6NPYxAvFVOcKSpiq
KttyUs5QV3/5/SqSGqUZ/500ZbuGkWpA2n0rLlqlLihROlXVOBRgiLSUYnlo2/+Z
DnfpG1ay85RzQo7kBhzl6P/UVguwfUD9RzB9WxQdih9xAFThI70m6HBQwRqzwFgs
/DKSe17P7FklVQ9laOx0xjdqT5ybKiVBSHUwC5TMbezZFO+B1yjUQR6xG+E5TZFZ
teIiZj378Tc9a43IIAXQ6cGhBZVjFGVAhiOjGeH4RR6sAjgRFjmiSHWM/yr3kZVU
a8GhYsjxPl7NygNStkZFhQ0e6EOTlA3yw4xpoXWHjy0Q3fLr0pFRaPvX2tv3I8It
m5GhgYAK7LfgOydTfTJrbPu/zwPpYCYioGP4gzbNBti10T/12K1huvjqDpKR4TBb
R1eKu+sknsaXyw8XU9IPGQE9Srz/lRwWS2QNCs3FH0cPF9gDYe70EjrFXjUEa2Tu
tsxHU0vTjEC7+5c8Q3OffEd4700xLQZpKLxCJJntEBB4XO7/Ofyx7+rpg3TLuKzo
2ElvWD3YTOXHzbygpg4VCD/H9EhZ57CyiPa8Om9gKFACPC+mKOhmvQWeZzz5X3+4
iUZFALb9m9UAs4BJ65tem5OX7KAzHaegYgAqa4bdDx1XTFgMiEIql8NTOYIgQFOq
XE45C/u3rrl++PJrX0189/INIwvjt7dtuLHc/FwfOX6sBhg+ChoCYkrZTv0zeCq2
7Xc42zck4tuwi+pot9b3b3iIgFgwk+98yJACc+780tpLgdV+tfweCdnDNfW5FQwm
fHdG55UN1V7aRG97vtUaSzSE8ozwXsFNMA154HOTswIhhXQt8O41P2LrqWVQKAxB
Wd3lhlAkFr3PGV2OH87ZkBdvib3bRE7tNhsdqnTmVXO+87Tyhin9FMqDGcTvO5Tq
IReOvLEm9fumjMb+o3o30VO19aYYmZng7DEVCU85bsNpizOHo/9tM82YRYoIb3Y+
41KbC3NqTsxZgsXxrFxsl/5/IDB13xz6UbCAqdqfQ119FpI+DeIDJsEg2tTlrLZv
LNKL1pRrOorQONo/BsEe7uLrGm+WQFAyihHSKgtBowkK8wzIDt2N5uzvzYqnojWp
Og8QmAXzRpMip84ophaO/0lojem2SLbwIIHP1E7z3IchCUUCkLfM/pU0RTjRlwb6
3q6jV/GX4+vQnLuNsZRY+WGPcnKKPMX0mO4nzblfXvD+e/Ezx3PHJMq96c+xKwlK
AZ5wa9AZOiLOLfw6Unzgj44VhBiWndWze0jYn+WiAZmxMOBJLrU2GoFw3qyHnF6a
K4wu7F1xUEfiDyMAlvdu+Fc5ViXU3enH9aOPekpFdXvjz2bNf09pEl+ajKaF0MTl
h6dEcRVH9S7iobmX0xTYjdqp6+H9vFoXu1ZDPqg5QFQ+z+sjUgP3d3f4Gw4dM7SH
D3hGYghXhu5VYqKFXAhbBWwqEZoFo3yD6FkyJTq0c2YZ4oRpKNeCBE6lSYCPJycq
b5W5yXXDqkO0zhVmIt9eAPWq365Vo81JtPD03cwWQa1s9RQ9VmQKOHU4h5j938hm
zZF9q44v4XQbP3HZ1u5Qx9PU6AOhWgK9xCKNg6IsJfCGX9xgw9JtdE0RGplBnwH5
4QGYGdi2NnfTnoEaT9EIWlYe1+19MHmnuya+0KozHE5lP+IyUOqgWc2XAznPOGaS
RYzbedH3ewQoJ0rRnsPkaeWg3lkvyLf59yuwd9lfwtj70pi8OpnNYFOv9c6ECnu9
JRy4uzMxNLdD/AMYHw6enRsPM54Q2aIoVxGVkHADlunefSpCM4LaIUZDXkPpwXZe
CG+Tb0DKVKB+Kc218D650Rh6vGzDPPEoNIItviyea1qXliPdFmAPNF0r9Md4Ei5E
Mb0wtMHlOLPrmOw2pOze5/44KEyKAPMPKkQMi4w4Oa+PMZONiXMK3HZY4E3Ss50K
+FLMUx3qIxegEhOSmB+WFo3t+9ILwoc6EPngCMRQoqhdnvAWxWEBMQfsVxN7iwg5
bHgW6TSQHTKhT057vw5DzvdtcyRxzkWUJZ7lp1Ss20Fkuz9j2NFdM7A6MEnUm6oe
0GaHKctPFimOrmmcqLGk/PRAvHG/6BE4uwMbunCkKdwdWOaTLokCXeLfxPYy6AAy
E5p0omER7xWvu+DaiOGlOd58UxgULb6wmwxr8B59sCTpDByP8Hj0/xIytg8gDvZb
sJjhFP1O+/MvhCDeFiubkiy1B+WOvBeAqvl36iDxPknwD6cnDx9r1IaYK5bSaxv2
Fq0irDO1x8Vcsk0isiDjZShnhrIrqYw2f1iz3vfmcPxYscwjb9zK27ed/f3cti8a
XBbQq8cbXQgrKbCuLYLBIDBmOZ8tlfziDZWE3DTSU2TdWYJs7KWWf5LlXyusRufZ
f1fUpemURTliB026dbl4lp1YUNgy5YN1XCRW3c6+SKn23LUTD522cLdToivfXGHE
HUKr4t6D6aWXtH77Q/+t7Oh49D5QmW7cGjIlrr2gRXZtkV/uLOkUuuUMu6BP+rsR
j6vansBr0PWbhA2mL402Fn2YHzVo+Sk0BhqGU60ApwV7X4SPwCuLtIbX402NY3Ba
9IS60hXvnkvre+XMn4y+EDEWjzwhzYekQQp1XowMvRz6fu2oHzO5MQ1my3yI2k4f
VC4k8OkIRCsx7g9ek1jwFA2Jra9pBARR+ZdToaLyU5DNMS4fJz71S3UHNln5FxnA
U0envMkiBvny4GCCex7mKzd3EQLm8GaLW97X8Vd9OgslbDFP+3x0enV+UgVFNrSW
P5qFtV4URtAkf6oIjzPEa/qak6doskjnc9h68ic2yU4/G9YP/PbnqSCy/qXJCYho
uqNJKfPBjc5WnrcoQKrpghkz62rpj0N+sQlKVnUi5thU5ROSKEOVj1dIxkwiF+Ol
6CoApHyDFtgL7fO5UtgdhnxS10dxgUTuBHzoWicwKl2hXsxHswWdyLasaO5hfRjQ
f6QHQBWWr0qq1v/Ri8uRcCfIjuU+SPvopuvJLmCOJCDwEg2oozNNc6ac4LIhdJnS
nX5bzLbQCl/EmeV9DhuYYNs/5vPftg1v2F0rDS2yOCPpIMX+ySzM2NZJdXAkG6ez
qvwT6ix6VdslB1LuGOIFtlKSfM5YWx3O0idiMVBH2cnr1xyFs0gBwkFnoeViwSLP
ndYK0yqdECU8Mydt1nWw6Yi0Uk9nM/3uy3CXSVkBYYkLR3lc5abHjIwL2FhJxE7f
/m1RLab4s7jjmzt+5ctxQhAKJyPOuS8s6dU9KyVN7x/R/1zTtTXRMdWkweTvJW6c
L+gFVBqCpa6tAf7TB3EvuQF+pSEuUQ3eUefOh5zEVl2zq9hu6K/kw/Ob8QM/Z2iE
w+ekQf+qJc6exbMJwhK1xXTxKAWB7OdgGf3JAQk0o96z8+inShYDa1pQRYdhhwoI
F8loDeUXWA+IPJOTNbk3kWE3aVkt5AnPiW5JM0+0Da/z1gd1n3Sr1avgktGWlAM8
+Yrf4MgUplzZjJghVWPYdyD7NvckR9ZZ4UVDW2FiUMa/muap1KZGj6Bk3OiQP7eK
tpOYBlqbWKb/5RZUoqKWa+WEUplM5RidIXS6kxujyPcA6vMfPcwmb3TFlL7Vpf/C
zFDzqt3CADw9xY57bSm5BuovyVCdk0AEQv0TTv8JLbiObnKKPx4lrwlW8bPM+rEE
bsSEOX1nMvPIlc1Q+Rkaqvj5qh5xTmrFtbE2uu5eFFRM9G3l03l+o+RQJeH6SPr2
4J5uj+G2YneiVVsi6IYlJHcrkpyQxGaTxu4Bh6v+L+FaM2OjsP7D9ccN/EEQ850Z
dXC/fXldPlRngpcdam0bfOJxiwLfzlpNht5oGH1syOrDqf2SrZBmfWKQQchDH8i/
118QOCg2JcYm2mjBA50kwyVsodVtsie2NfTIdEmwf/2nLiMyql4R4b0EP6YDGEIg
1VLBhT3KD2yK8Z3q29EslStGj8jkBopTDRXRD0sm0jilglDrp37HwBBHA6MT858T
gwsxeCYSkadRldfE0PqOXDdViruezoaXJHUeHXW975W2ju3ZgSy/lOYHqUzX5UUR
6LxvSfsLrubpcDKJ1Q5gFeXioQwfFiiOMo0QGrGossS5uBFw43DcJWe5xJ4LW66K
8Ativ/9Kbrp62iBNV5qpAiuL2LqFRJObtNxBzohFWujN6aAGDl1CydOK/yWGKqjV
gnQRcUYdbgIoW3dacazhcufP8vtRO2btJHtPd586rC3gxitaHI3lPecrgVRWPhAR
8zP3NPjH3+jgVOOSr+JOG+mNMS4m8ncSfpu9LWrBHUkIuRHtRK+QEbZ5qrEGYdE1
tFAmvTm1Qiw8AOBi8BaXX1Vw3H7C+IgP9JdcDwnpzUDvRoxXOjT+WPV8JZOF+A3P
641tlhEF+PIXUQ1U/9yxVgp5yS5GG3OskuB6c89O2PeDK8CFi4/L4NKGL/HbxbOb
EqR3sFU3votLTct//mfu4bKV3sQWRoz0dZGuONxR9L5Xygr3a/fDvZXNni58xOBG
yB7u/LrehhAdiatjC45Qdsquiy03wiHz+WfUSq3Mi/o//LxI3/RaFrq5FAJd6pkI
3QWj+GnTglCAtug6FRI6jghQ53tWd/UrpbnhMRYyKh9GbUz2/qAeCT17prLx/O7c
gsRSkkVr+Nh/rxV3651C1VgqPv72tDcsxxAsvXdhi0knnBznlMnHVjvCBOTbG/yV
kftu0YeRfOSusjmpUz/zVKqZBG14xks6U10uOvUnbda2FLbvlNrMhGXueMygr008
2gscQh0mVmiKqMRWX5lFNOBOJPdfgQ0PbC0OkGuz2WUFbzdoehm+7TW6Am3eu+W8
Np/oFDPJpM6q3TVYRi1QvURxBOunkNMomZ5BR1pal5E1CGMYu//xqyPfY6yUh0tX
A95ypgXFOLasvMUMIPd7uJ1xAb3FHuhGvz0x7J73mf7k1glZbp2Ahtx4vsGBZ5gL
QKJehCRTDYIAYc3le2PfC7939JuDPecQ84AgqCu+gyIDMJi2JMq+PWfmS0ZEfVKO
eIlgtXcrxuESmjKtvBYLFQFnPXjMOuzJJ4qva64kbp199ephj2JNI3Na8BWhKhdY
R2VJ9j5uVmvQce0am50MOvXBLSbPDb6gA/MgbDJ+yLj5UMiSh3M3Kelz5A/bD6Fd
tfTggtjdnlZUmhJbqfh8y6AbA0FqoLF4kOGglf+LmmihXmTffbfeacAEKHY+jEHR
Vr+kNyQH368/G7Iv5vQs8XiTrnVAlQweyPsdgpTHanofGEISuBlDQTYnNBH+YaEg
laoQbWX0vJWhRKoPEx+oIb1jBVpt/av6HqFpjfiVZwq+gedSD0RX7a7ADWAGZ57j
oLh5WoV1JzkIzJHisNH1Qg5vzFYpwNrhU39evS+u8ZZywzg3XwIrLVx6FSPFyKDE
Pfpt5MwGlTNLBATsFcZuc9WT3rL3IjvBmGEMlLIjDlsnZbINmReggIj648qYrDOF
3tTgoCj54cQKdwD/SF3c5cNpcFhaJwCt/gqovUHsnt4p6Aws4YAAwg0ww9uCqbZR
VR7lI2dhvdhHGbJQcfBwWfloJk/NQETVxzC3OrdwoHphwu/aV7hWgkoM8jlNLNG7
5xWtpsPdMj9Qlw46M4xMPBGULv391ZN/jVr//PQJaRV1XdupRLwYZIvM9RQWljwZ
16LNe3DrLwSau3JaXgHyvRtFVwB2PEMjulEOssOhGqZIADz4PIBipfGAv1ybF6Jt
Pr27WlYmtXYLlRbyMZwzIsYMU+hDnEAZW4FpMY4K9nErC/0b2Y3LsFZbU9WqVNha
9V4aUyiCwrgEW1dW0tSdWT7Gke/4P+c/vLlOuP5/szBU9MZQhEk6/NJwRXmUlek3
h46xMGcMoKLSavcml0x1wiRyZZzmWfhJutzxc2UKLNfnQGHMRpvX/auJM++jlmWT
5PgBEgGl0KehkZmG6NehK0DVtXvlrQ/j1Cg5vBPCCqh6LNqTHQE/8mxSpzYKUxYB
GMxoQ3RmoPuAxS7sOv35kGuHnEUCqgjmot+bsgSLFSp+MdLejxrxw28PwbAZ7l+i
okfK1o4lCx7grM7UsA8rjtnLArFPyQ3krPnVK4/uAFBHd5isYIJv0wbjIJ8iVtzd
WoJ7ct7jX2dvjS9eGyY4ffEjPlZew6cBhgefrr6KWvT4WqFztRpHkw5sLb1EEAA8
oydIu5KMqq9tPXv4JPPNFFUxxl00wXDEb6luLtL1pE1s34AXn24FzxOSfgh6ouIB
4H00qYUBKvaaJiawZAXEcV+dN6s/E0dXoZ4OarQZNYryQU5oOX58nbRz734sPa4e
P3b/Iealy7mMhwyu5nnmOZJOAvJDTm4xC2VaPd2rf9plpbMk2R494t7jWkDqKHGX
DrK7LKFvC5Y/X4V7VDNjLhcs/GrAB91w73vkibuG4N/2Ev/bnPS8kAFDH60AManh
np5bPxk7I6nnqMtlhHDfAMU+IPG3h14BgfatwH4e4XMEdtz6Fai1ZJTqRyHfiEHx
2MskQY1wA1RVPNMm4dpOssngfG+aD3Jpa+Axk6vJfvvEYphQxmyQ7P/V5cr7rLla
Y6PE8faFrVu5kV0IMd2dv+DZxz2KVO0e5neClFqjH3TXmkju30pBfqWQXznVuRyy
clZPo/lAVC/D4lSz5xZGJUgVRR0Be7HdwoHzkl8DqXupzf8F4eMYcJAqcl097ALI
FWmtSDJIyraOGruX+TohPgU1sMr8Dr6f2Vclukt3FrZuA/I8kNl4FrhOqLRk5BnJ
bTqu/NZFUVLdvcpcEFd7WcRWJEdJ01gdQzHKfy5Oi+WvfJ3uJwbj0yM579QpRKXr
cxHw8BdO+pwYflYiPAzlPRC+jZmiWIk1Ip8DulbULkQ8LdFkcQl2dAzfM23kW6oN
7D5kpjs5gVf6DiEfNF8aErz4FzGVhAwglCkW9ncqpxagqSKlOJ3hfes/Jjmjy7bd
Kae524vQNuSTzdMT2xieueaPS3CZq4E3R7pwNcLXfFNtoKZwEk63/ER2qwAwlZL+
nkSkN6ErKxCMONqht9jwpjKSGlCuX0zGJPCI6f1ZWFV1AJVODQfywkbsJ33b5BwA
6n1K8CljDx+GI/9uIILo+89dQcvIHrW5aRU2eBKX2VbUtk2zsSwwZOYWznfjB2pP
Tk8BZm6d4fhT25KE3c0H9RpYoB7mj+sc7u3osGKbgX6Y+1w8TwrmEYxlXJUN6w2S
eIDnRuwyrlKSwspwK9Z++eKUJx9vpqqYWs1RO4fr3hA/zrdB4c9uKxQLoqxmhZmY
iZvwIk42vRvYZNOLCI7h2xpVhz+0cDOXcGVlTJXCXWQ6jDTrASuRXx0JPlkMjkAF
WHldtr7hUw0hNnyg90TRB6+Za+8DSLLc108NZJDjA9PHhaNJHC30RFOoA3gavUJx
zUF/3SvFUm/e80T787SXAtKEo2fk7H3bLm/TMzPM8r9q/Y7svnXD+y/Qwt7006gI
PTzYEDdtfVmBKY1/mie/TSad4OwG6Kbkt10ktUoJ1qjxZ0amzVSB0So/Ph5ADYQc
4SBclsXJZdXnZMXoa8YQxBGI02doVnubSZv4BppsBv/slVDgSqe9qx5DdmcPdATg
IwBHFjrn4nCFIcRd1IlJW+kwwP5Nz4mnm2xxLUCKhR42HhY+qlGZtP5ie9Ps6D0M
lYDl9ClrZVOXYdhukyYGev2QiTjHLySxBpyA2f+bKNYd1Fb/oEyztIeE4XGc+ob6
B3h7u9icuagQb3Qvk595+rWLoLPDvwy5EOELi+HNNy0ZW48+R8hhh85MOhkn5dSC
VuX9N0vjkfkOTIdhoVNA9sRaVQPkNVuPtCDGD7M5ZoTbeKgHSrZQ4Xzvh05GeOEo
uPajUmv1h2dUUw8mtNylG0WG4BWxlx2k+/8vgn6tkraH7fpq2xuhRujCwyB2Z76q
rkaHO3kfBnncFbXLlPXEXIevwcViP1kJ/NMB+PKs0ibqgpOdWJagtCiHBPkPpm3+
imSPOobOSjLivsf98e2YSXSLEhznYso5Dz+TIcsSahzgA/GCXb2t3nn6Hk5oWqg4
178VVZhEZHod9rbLHnc7TZtdD/JdgDdO3fMvhsn0bMMQtxxk5KijY4IRATeEfG8V
HQbU2EjpRx4EIG1SYJGbECYjArpr4aI1d244iPl3zrFb5+J8kAHmDuHvOelrQ2o9
BI4n04e7CKV5JzachIVYPG9Z3J3gKmxubeiUVOVIxlVl6Ai1vwT5HqX72amPb4G5
xzskBs+sL6MmuhjR6Xz9JcALlOpCRqwWgHAfh9JoqG2146n0eMuJScQdGrq1us5K
tXg6wLCfy6eCDTN4JquApyyKVkiR9mmACsBJOuB/yGSULD90Vtukm4a1ivJg8i/k
jarxOwQU5V8b3U2g2yswA24Axx9O8n71iFEMYyod2sN8m19LYTJA0xma/f9duIDx
gkydUFxIpiix3Sz+WWPNXNJRmela2fAXDbSIfZiPOoZWcvf911v0hE7VDQtogl4x
HGcTj+cjzLIIld46FMv3bEWY07bUOtrBUZykyucek+eJkRVqZnacONiHkOVqRpGE
9yf6bSPsNSYygvnx59yYxg5M4Kbu+ML3xAf7qgUPdJlKGzDsBCZLqa5AfCvfiITp
ym2F1us2KkVrwyu+5Nz5/UBwY/U3ZsGGPnYP7JANAbZiT400p079tFBQSFe4ShQ5
Q8gJz5HgaUV45xu1ui97pvRZNTozsOwEJ1gKp/7kTFnuSyBDtuhIdJswgagY9Ap2
GH7nYDl8rlNaRSkRPSndJ5jMV5kUWcbvPlveq27KOnjU1PSDoNDUcEzqyemnsTbi
XQERBg5p2lL4NWBuJ+2/bqgxu5Y0BeaXWCOJaV44UvPGenHwuuVUQdaEBzQYHhU8
uoeqFm/7R41pA0EH766aPw0vFyyfQtRRqdnyL4NPyiERp+4/m86ro4mExKt1Equ0
3bqRjtZD/aYeZSltMqtnR7/zz3IM5ig/DG4AYmQO46vHMVMUQFvzhp802DLB+sLx
ll7/yEF2KDuv1qlBzrFC2BFWst1qQUieB7qY4U07J2a42zK/2iCG4H9kWP7MKeCk
60HMBamU2ToKf6hHVPkbEl9mBoarYkMlUTlancyqXrjRkenIa4+1IRhczlSgSiiw
Rt1w+LmcgPFkFogA/hMJAEU7tsW+16qtkWjfSCAeKOdVv7BECRaBzbE0Pi/rnYqR
UwtzhzvSgpq3WQgqFqTJ/NNpxA/4hdS8HQ/3q+1l4GxlYPMd7sEbSRbpKgFnBnLk
HOqMaJpiy9fd21QMtsiwoPZjFGJwcTHJ2l+x215dJDRnyjVDncLcWoJikj5XFfK+
+rAwi133pHAMOjvzawErsfZPNH0THJD747Z78MnQ3z2PEtZ7UCmpSqmhbQlFn4RY
vqmRXorvUzC2OQmoctZJjDCTZygaQKAqBWrmamR3kN5G3jk2ZHhiNO/YfVXJZ3Ki
l9KXWQMH5SgKZHSOvcApAsSOaVsKPS19JfQj8kEVnmR/FZaKEHn8McZ47qDUll7R
JMBZZV93I64wbSQmZ8ouiR3+zmobWwPPzS2+pS+Cdg+PHKIQ3qCOZZxNIszNRDzd
AYeQKT8y712W8gG5GDAhH1XrEQOi/Tdjn7IEaJCBeQU6a13b/nRx+YoMZiyARMqP
1GUO/KgnDokls5gYpnVvc8lOXEbTx/b84xRyz/z7YVuPwoX/EXbQPljFBzl5MUEI
Ho1xWeFvzJT9TasmVkN3FOOIjFo2f2CpzO5OPycoTBtDe/z1lrzhT7MnrjLkdodr
ZgWmbE+v/338mISuXQWwgCwMR/Bdsf5bLmc1odjV9RCqKN4JlHhIWZMALVjEDnej
9a0KdGUnjygKbeQxRr0SH+yu5YQJ0rebHHKI5It7sUUQZAd1rTsLc5NWXp+V9qPi
NBnon3wjqP0QxjgU5r/sZKrcpYaXgU/pQhHF+H4NnLFm7lxz1wwJMXay5OfimhET
JEwZD2q83q9Kg+kR2TeR0j6WK3JBtPf6/OrOIgutMWJjK+upgwB/31lubb7nI1L3
GEOwO1IKEWcPXbfMhza5ndeYi4PKBKupdTnTn9iIc6v25h9DIE/XP3iKDkFI/dl0
bbGEZ+fFG7N5SoJwAoC8NvnYhiWcXPUdmwA5LqZ4GyZxocS4eRbZeqTqgPKt3RfY
eQMrW+DHGbR0fpE40gC9RnUYGKiJq24Ex8NDuUyYXvD7No+3jBV2bHMsBQi63Nqj
70Qdc/K+LVNhUAULznJzxlxXfQLbdhtnuLFIuAkwArJH/uIMSJb3QFwnOw1HyA6q
1GsCuQD8qoTLp1a1R5NYDuvFrV1cF5/EsKTEGPvPVQaVhKMF0CuXzjInViZSKs4j
uDKwSqhpcRW3ZPCtIkL7uSOKPdTGhI/kwtG7nv0iilbpAiEAQ51fzX3KUdHXbd2G
DOrpSr59jQWRJAJ3ltgU5fn2a964YsN1zx6PDuvnwAhJj/yKamWiZHm6j8KiW2gb
uE9hzPbT7skFuyDzRUPyFvBJlnzPx8wy5AtTS71v0UCe7pUM6mCFymtmgNKuUgpW
iSlClgihO8Ad0QBs7nG4dUAOXugi8b/0XtOJUXYCKP7OCgKHJXy/iw8Kb0ix8oz4
tfUpQiCWxh/YvxMum++wU/uVQgjWijMSkETVJ9EbEeO1ze3eICa6x8nTBeNItIdd
0rtv0s+S7dRFZLK70/Ij/6m6/P6V+OF6g+8pm47/ZLpyg3dMUWrwBnKwMaDbSGMc
qAygyR0tsR50DVLjfba6oJ5ELXsZu+lGxS4jJf6oE6KIzJLVtzSaZY2aU9vo/Ei8
qkFGUgEfif6GuZ2sZhStATkq07eMqSUEF8KzQBlwuHYkfsWh1orHzHXTK9Zydamy
mfIvZGhxoW48KnaZcV+Pd+jXHoOFhB/Ul0JpYeifR64ZmIgtEfxlT9U9ng1q/45Z
Hr5DxjC/AGUwU/bkC1PJtlWQpx2NrhtOuTfINs2tdTS7gHHW9LLwO2ggxF0euOZn
1QfzpmdrWtHXWSdc7HeAgVq3HyeM+HI+I798M+FJEAL2l/WuLnhWanE+bpUc6rLL
IBEbdQLSORfycT+hFE2s3FeGy1CeMQgP5p5sqtHV6XoMn9mU5eqBuIVRn6W5b/pc
MV52phbSxo2NewXSYdeEGvZFOSntH9WPuMtqTj7Ja9KAsq701BQyyg4xYIbDv5KM
QulIFx05h0UIZ+H3Q5K9NXevkOsn2rdeo1BRO681S6SzVNWAS7lKy0BTYdWr3xav
KsbJMJpaBKXUBfBKT/8OmHaxEaGdFZtWiluJUnt+aYjRxZszm/nc5nQBdoYxyW8I
tMI0fPCbSYL2LjE2HxJRlO4LECw9A7TXRnWYNJBXcwTeXexssTBRTlVqweOGfmyu
cF7USsQRCuOQDst8xxdw27jy10wRyesRVHzgsXox2acLasFxVQHNiVtuc2rbosEN
lmw/nWvr71LDT6mk7fieiWFpHRVX4DOFxcve7VY+dwD64crVbC1/fAZJIKhwY7AR
lAb932QXgK0IwgbrQckk2nARJ/7LvXWSwvh6zrttKOtERekc/qOcaAGNKsMkIdua
+RbDT4kWvvBvFB6RlT0XlI9a2I5ChBafOLQihj7gBZ9Epm4oV8tt7oVLrBfP4zn4
z2nH4aY+JtBHLn+oD6zpf8+ocCk1Q/1xc5WlVlnhvO75f+AXRcevyYRZH29gmbC6
r+jCYDPWfTYM2D+kXDKZB00tta8Swn2sdCJSmM1xKZwVN6RRpw6siWhy3X+GyMVG
Zq9EoNrwF8mAOuKBtgI5ekKpqJfYnCX1J17GMhT1UQeThkqRvs/dO7Ivt/0g5RFN
JZ5O/FbPZ8sD3vvRYGxUMuewVTqwkjLm0ZMHdPcTXT+tNk68Em10pHMByvLvdSuB
aSyQK8TnnIKWdNfuJfmiqbqmnCxhKSU4X+gUpWNO4gMrsCoduKdocS/0Ek5wiNJE
z+Dti3MdBH8DxoBMla3xSF6mzKgnVIQd9y9f5Wi1GP91ZzObwePdZJdTCD99Fu2p
ahAeshpnrMaQ0awAh97I3YPKqZ/h+P8IsnGqGNARH8KVM2BSGNpga1c/wDZoSm9N
tfS6ZxmA2JQEH2Vid3LCCOVLzeCYuyL3iwHoL2fq/l9xgt1GkOBcBVd0R76ebQUd
hAiUWNeSTN0URtJjB8onD3qTE7F/5elsrhxU0QHIJc2y9ABnemseXPl+dVnuXRCD
HKI8TbPQmnwds/zT5etymezpEY+GSpfZvo1rHmKvZ5XdElOLwN86ULz3BZNaEFsM
9HUVrY9JIVzTWLellG4HlhYg2YEkXalOREIkcvSvcpI5NSoZ6tU4wGSDBwmUknzz
pDT55R1ICPspqtV6KoTy0Qe34GRB78fjot/I3XDz8Wi+d6M5JUoLRPTpHtJUdxY/
gDtR3/swXFxEFcJE+5Iu2xi5FgO1Qvq5wGY+L+72F1n88ekzOHYDKxXgM79J/hxZ
CE9KBNs/8f2t1FMcDCVIKDe2+kqjYRzhH3PcFKV0Q11PlSG3w+tcTunI3aHD+CkN
v06TC2leFuIzX7qcr1zzLKRmTlbU29O0EvagtSWtzbpVQt/1RlJXvxkPgGj4SEN3
k+RCI8H+oWUOlFOxdn9v1E1k4JHcVuKPCOnKg9fGIGAyVlxQ9e3XToE/6cfVOXuj
T8F0itce3ujiuCL2vMD4r9brL8zE5K/GWcg4aTQtmL3H/6t6aRFuseY0afKaR29m
a72uhjmqJEGTmXwNDZWsol+rtB9fib012sNjPuHew4VW9ivn4PJUKKwPtSCkb8pY
hl/B+KWMweDGboIqF2UUL4XLjO8wxFFRmbalyCTeRLTEtW9d8qKTAe50T27z7hSh
PeBAYkz7iS5jwDHaxnRRZRBUXyq2Xen9sVcyFv7qaY7UaJXgjejMWvHCzXHY3qoI
5ZPdGEOqQ12tjE4tL0BZxRzonQMufgUAAybGElivRZQxrQuh0ztpuYL4k+D6sJj0
GrGfQZKM9EzQfnVgm3S3ZrZMW8jwB1KHBgv8SwG3CasZPcMzj+RwqI1OqasyFbAW
Jl6a3foMwoV5U0BYDBM5lN/Y1bgnyEnxoRG8o9lCPSTtzZnOoycW3wgQCET+kJlK
eYb8uvBNhCWhfDljoxjQ4E/QUBgotnoEk8wYH6bJgla7yVlc28H5GS5wra0Zn/dY
e/PXgw6RjSNUGGBULg5JjEywHgVDUKwr3e2bKpzc0hPxW+5FRi/GUqzrNPYHfTHA
dWVXivzHXaVZLpoO8oQ1TYJ27ZcoTi8PCCMzUDPd2I4O1aVnXZGpY3wSJ/fvGb/7
rjk4zjH9gFyd7oZkysF0u03ARgMLBZDUaIVyavw0TQISe7iVzwCATlGTI+zBLMNb
WyCyO8NIjFJcQD3OiALfVYDn2G1XBMMWRvISDj9mWSzMdIMJO/qfXL40tDWtPhJk
ehSU1/cfp0pfDtvARWh7H5GArP7iCyC6KROXCm0hSz4PHF9kLe9l/p+zZDvYsWhW
0pvwVXI/ttZvql/Kgwd6OXBTmfe+T6PbRH+YN6L7763PqWGydHKHh1+3L6lI0vnL
k1ai88JKk9iC3HtFqL6en3+TzzGjFSj3MKo03byvSU+V3+X+o/MQKVRu5hEt3cmG
S/oPVFq43fB81uryA2dTy8zrOEw5XBm6npt8uqe436eNIAphsBuox5WSYCPA36Iw
M7RZaUYU4J6Waa/DgZiKgyAcpa2jrmf+ERHA31WFSTC/XWKqSbei1V2m9PmjheJw
8JoIJhpnxRX5+BdshOsGoCoU4v5yupvI7uGZQlxbbTanCE3utqyT6lyHvSahIymG
/ZH3AzQj8xdoxnTmc8FQ8nrOr4mu36nd9jukdkmPMx5OwFmLCX8I0e0FhmzUfr0B
ct6EmZjC5ZuMsfpLayBdx2bh1qzXvhTtSJE+gqXrYiuomLg6XZdr1tDIgNGCtZgr
ZNS3JQ0m+ru9ArQAL7AyjwRu9UbMiMagKNnQ1YiL0UGMfaV+vJW34rOvGmInDyrk
EEicmxohuOTN5l52q4DzyL8cwHX6zHlIZi6YJAEp4ytxC9OmOcZojxvVZ7RlabRK
vdJkaDNMQGicGOOwvbLbhbkBkrLtUB67rtSt/aeMtJDkCMO+87Sn9WtIMQVnIkP6
GNsqGvcckc01i1UWc9bYk7IlHZSbEGXCsNuVDunwisB2n8VCCoZyQDUpkgB5ml7O
P+NmwMAlJNOSWG4UkmonGtC6+f7BLapxqLtRppMsYgcxl+o0CrS2qo15BdFgUc1W
d9RWbOSEJWrOzHcvm26UFuqy/XNFyIY89XyxFP4Y6CCcMTWVUnyNznsTVs3dJAz0
DD/vCy1B6ics3ZhEedXauzR2gQ5MscCoscfXpb/XVOZwlfJJC+ZdUZnuS+PnKrHY
W49CPTMm8bw5z+LNN53sSOxOm5vnH13YUKid6WliBiDT9sXOX6IoZ3XmS/wjxeKu
gEL6CXPXaj+uUnLkYdkgOKNX4pQ7O1jgaKb+KvGsJ4Pn1IhUwuz6mMHyDg2ER5fj
DzkulufICyflnvXt0pLk65UOo709Oz9er0Den6BBLIZ1hAVwH2jlk5cymJrJvxPq
SEeOAJyx4jyZSp3Cs/qA1BXioepIigwLBZ+Fbmanz/anneFzTzlKGfd0iqBmwLjW
wJJli4Il/NBDTmHBnN0O+rr3LDvVgVRPFCGNs8KUnuGE3diVrYCIzI+jAh2YDpy9
PaUZk8dbBDD5nRJm3UNH9RmiyJBSQwB/+DXq0amFRjO+EDlKnp3k31BwKeSLp53A
GCtvUfS3RNN2wH1gIzC+QIBS25Gp9fWqRODmZmGenlxBbVTU1WMm4wfaLGC6YVDA
3MMmHSGwO8sER3aA9po06IVPL4gehSIAhX2Zp7Ju12lihy2eeW9j/FMr+id8Ba9k
zz5wu3mvnXYOI26xUZ1OT8xKsaD7qzn5s/zTFy+xlzSZ2zKi72zNa5EodUbWQt6t
IezMTCBp5UZoTfpeFnmtGYbIfUANFkwYJVkVGZOFZhRZ3O64Txhwij/5Odgn0f1P
1ClRjmHyjHpHnVnWGEoX/sBunUooG0T/KFJl+k61J7V9uX5uPfB1elB8IUi2zw+i
TElhpdlGh5DE9e75mxqRpVG0J0I0r+NYW3i7pT+XHz7hXpzeYM6vX1BggqsUmFyz
kj9H5osBEy/JjoEv2x5IRVMBg6Y91lv4Fd939wDeMKcFDLDKz6HvhJKcdZ4yZqlj
S4PYAmdozttXTlk2qMlZL8D40EAeu3jDlIfbVnkHjTvO0vKR7N6qUxOj5RDYZg2y
YMIF7yFhdrPVXbrMkTVKBZ4EfXiZfV7gjnBKt/hXGgIix1qYTdUgMJe7XNFMHSSw
38bCKgIjappp02zh9SdJCfRaH5S+eQGygjfXlxINji13CzBmHVHe8zTk5+D9GYb7
PYuRk57ZlXg/nIsxwmb/zTH8Q72NlgNI2qIWI3Qb+Gd7D+YaW5WrDDrbevJ0fSv0
vTNAxuDNOPoSDNuR+sna48SLi+KZ7e0/Ly1/gY4Bj1RQsc06ApnuJum7OOoxOO2s
e2FAHIJxvH2ysFze/WDVHB/McZEWphIEg7F0woX2I6WorgobplpG2VCYpAYgHNoH
OkPe67B8MeBnsNquAaRfVw+Tjs9Bri3F50qYKF9LM3Tu0NA6fpny5RZkNRR7r1hM
GJ5I+154uyl+xPzMG4c/9CSWGRQI2CADbYgro7jviAxaT+kS0w399/M7S5BBCa9i
KHcto8Vt2i6xEnOh7noFpmczNFij1cC+8adeYnYKwXU/AHClwTpSs4RJBisPXdRc
4bft59hC3tIn2dmynSv7vKindfQswK3bdKCpbjQWj6qRzZBzcpsMw9uaKai2u6dJ
nkvi3AAjyEisBx2kGTgQAP6fm3KzUadGuSaJby+sFRdYUeH3m34BwAtIKmr/8oXa
lJUbOQ3M8xEzcvGHgdq5h2kKApUn+72PiTBECTf96T3tGD3z92HnPEmomTEYzkdk
djbXd0t+ZXsTanoXbS3J5U3vOO0ye5Gq2Ra49fsea3oFPUu5gJCN5CKolMqseXZm
oqOTuJAJ3rj+5NY3hyJM9A3vZjy6yn70mbSP/6ZS+dzDDdfbHT38zzuHq/JrmB9c
r6NqfVCyWdQoW8ts9adRA+zEtONuSCuJlp/cskd3kqMUD2hCvbOY0cJWY0tGE5US
O6N1TUs72yfVoMPS7BnLOuzlTVYZSQu6IMu+h3HsbsZ2jYvz3GmBUjVM0ONYN9kf
dGW2ejpic7CSwpjyLYoDl7haZpHdmsbS1UP+gHBENfm6HBut/bXyVo1Dq+HZw5jW
ePoap1bT9Qb6XxluTIOmD9Mfu7wmXAdV9Bs6ookeCOVuG5AijINtDzrN/v+PH9m+
haOh8+zU6VRv6zQ5UdZczRjvQ9Xdz33t429NHmXj75Yjm50fSrmNothNsf34Mn8b
o4dEm3w/wr9a35Cfu2srWOqnEVN9xlSbbMRrUThbV6XBo3lD/hO4Sxy9cXTl3nxg
BJqo/2SkdYkdyTVF3PwDZRQep6YdhcHs17MtxoQWSqMu4ZIFN8hdKf8Z03kufK96
8V57d60je4kYm8X3lGAytYQ4zoyfl9//8biFvo712lnCZSe5jlC3hfvhgRlaaPck
MszjkL8XPbcmTTPCoUFQVLRNzsrRQsNtF1/wxcRV5Smjeqx+NmhaID8VWln9QQb1
gwaPCES1F876YuUlm5zZRell8Q3q4BxmWKa/Yp/FcRiw2Vr3dtAswxIDQbqfbCl3
5sOwn14Np/HsBqz+EV4G85qYzkhLCKS/y0BM62j0MEURQALkhYGtunvN/x5MWwz1
n6TLo6+Te7bKmQVY3EBu0LrSWTa42eIcZx7lGFMOY0pycE7XPtxpy+z5Qxg/rm0q
jXKiiTcAhabygXFQCiwxmVDHQbCP1xyRaKyXQpDaSXRRoSo4z5Pl1AgpTgqWijDL
PRP1jtbLq7Hgb+cYxdBwMkgqLP+jNQD1AsVNMdj6HXt7Gz7HVH269QLEbMIQPjY4
pBhQcRT9vjjyY0eFsMq25XJosRvJ6obuHLTwUHr2hCq4af1lSSXzsjNEEE0g06Ep
jgx0FkEbdq+tySNScgQ0ghV3LCZw5vtBhacU+jRXdWMtS6hWEAv/M/EvG0l1Plgb
NnO25iWxi0aTXSlrSpBNrDe1PxW5cBxVXiqLARqXHbE+MHyhzmhDa4IOWszNwoOo
LbqnsFQJuxCnVc9i3C9SgAsOaULitKwSx3Y8S6xpDuY+B5mFVmCMeZHNq2Cd3q9U
4jxTv563c58AJVU8zTbVhlpjFDJ4QclcGNLkTCXoOnN1Vgp/uU/JMLz7ozFeNWSn
/2nc8ekZq7ligAzihvgm0tTNfxD7pvde+6IckRLi0glTqCny/xikH83K1o7wM5mT
qE/h/32Y2yZZv+Nf4WHQxUr7tr238FxniTLrWvYdd+ddWRhSP1IJ/DfYii9kcs75
t7jhxwZnAlVQqJIaU9hJ4W41JpXANTPbYfSZg+Se0Ez+m4iT336BHoGqws/N1mWH
TVu4hV+VQZ4W8NZ7SHuoeEipsGbBJVctkm4OANQ4cmMR5qlfjUDh8E838cAmZ1NY
xh0VG0atj807ZDKqczivv/kMBUR5zVAJUwqCM78mT+pYRuh3dVjRTsFLSW/CCCfQ
6ipBq+hVniJaX1d6wzNLjW1XyxXI3ceGv7VGEcJW72nlSetLj+0UmefKJDWiNsmV
Kh8dBsMJr/wGqEPMn9iXcvAQf0B5pF3lcAfCoQQLcD6XaDUIc8fiSpRBL9Ihxy4J
P7+uuVNDO5R+fElSVmZJ0LiQyLf/8HHJhyKHGmZrw3eAtGmP2hvIfbx0jUevAYvT
6tA2sjXQ6xNQE4KSD/tQTMZVMTeBifTPUIhVQkVZmL9t8f0Tj9aI8PJSJAluhgOr
Cy8iuI+LzdD8zJF59RRRLDuFoJ6HENQy2J3A2AL6iSJX3QI/66CBKSpUgfig+SJL
VNfkrQ5Dhzu1L6B16mamE/LDfOJpMmOQJuh7CKaBGzFkYZ//+iwh1kzbcWv6tKlV
R1Osfh6X8IgmVPSnJpZ1+0r9ijqsurdEL9osAS+JDA20rmDTAFOHs+R5szp/bAO9
70r7Ag/6WpEDYj61HWsEui8ISwA5WAlGEBs0BviXq+u2VoZsIN+tlhrUw3ifsqR0
bi402GGnyL8DxyUidpwqj5otuvtOhCBq3drVKZEqK80C0XBbv6Ybacuo+prpWfAa
AGRYsxHW3W3rPL4QbqBeF29Tb7J/GVJsqH/rXuPjxW/yXYaFIZNV5kmU8NBaXwIe
BaFsspPy6cnLMVAwlr+d51TBAfas2nAP5qwu0yTatLnrFlmaDStQA7w0WoJM+C8D
3daXiI15/OMEic9kOVBdyfdJiaYFb5wc/hsPqlV9IG0CYJjIAKhvUcOjrFoG1yEL
WOQOAR4KvGzU/Ep6LxqM5HeuGPDo3NnbmAtEIZvma6l/VXa/U+bMFYTrdRB0hROu
IRwu1fIC8RqOGkK8NOYSGFbVtGop71v2JeSJKVwGqLc5FEGFa7PQnnFc+SlYyxb7
f+PzQLL0wpbU8tb60ABS5TiqlCL0oi+FN9JM8Uw/yJ6cMUiwOzTo6lnnROjuknlD
oi1/Be69XorOE2/0hYUVx/v63W9BKn/hnAZCIHi+bGHITiFrMlnDuHwM0WHdp11m
ilfpa6EddqaU1wEiznXqJilnrxV0zEw35zdhPpHDkLdd4N59CzHf2ciGM+OEG1au
mVxndbK2oDgDZbMkv0WPhkg+QzOsej7dTxalVVYrOpanjyicS+nwtJDpcmfXv4AI
UozCb+s3OP3/3+Rw+on8+i9V89ctonQnXmVvRagvNNVUGmpKev6t8D04OC0TIUyA
ZaYQCYLVSCUoxiqAa6x8kdUMomU+jRNyV6ZGN6P91NOkUzCLGIGoimw1tg14Ql6b
WZv6TgvWYC4Hauc/P3fcGWjpwfS95JtWy2Y4M1sgrvszR8fv3XEe90bVpMSdemAl
K1JGunb4lbEkD3fKhXNjz4ZiP3645ZOeQdzijKRC64H8jfSUuj+UdwcvyGpWp6/c
dOtsakfeeKi9GNbHLYKmWNEB/F/LSuyNFZf2Snlh3DZzf8uMHakBagr5sBVxb8Vs
5x9Wlgt9ACUH2ubMwPtIVRfoSSt5NLUHUvSVCqm0aJl+4ASjg2KUZGDB6Da+pqQD
YZ/5udPqvIaks8Y5xhFKjzEpBFphJOB+3hLdV8LpvZ4RsEExYhyAFIk5iSwEWYk4
JTzAlmCwVE+lFy5tCIT3FCmRj+0O/G+BCGVQ7H7W/UxE2q1sFrkHELw4kqxawR8I
WWlZtLKhIqiHNV0vFGvsuu697oHV4E8aoVJfyYYNkRuFJ3Yu/pzDy6ysPT/58EtP
gXOgYU9Qd/9JHDd5husuoo5gUOu9ee+UjpvpR9kXXGbdjDHfV6trprm/5kE06+Z1
IFt11qyDJASsHDhm885eUZwRxkNgwU/AZQH8CkuG8bF5rIg2Z3Y5zCVUYH5ZOwOd
HVGUmDp34MQ3vfFBZEZcv37230CjAa2dCtRzM49x/qawPAJNvcRH6gf3Lec1f45Y
jMLPocxrT0pVwi5SDLvwr1s+Zf5nfWUONMpQvsU/2E/FRUYHZbDwTVNTbftqzXE7
JxldLEWOgFP7SEZPAvaqv0DtssGI9tZjYZZibFQGj/CF+FEaDUiwN+P/h0HFQtLk
5rXArTtla8aXj6hIOs9BJd+jWcxkbKFhyPVsusn2p/ieeaR+HwITxAz7yDK4RRGS
WTlS2gcvmsa2KvL6jCM08WpXa86AEEsLYNBz4ITZsZB6+Kst64TwOOVqLUWrik+r
f+UT+cwy+6hwx0wS3f1lAIp+qliGcFLlQxOCRhdixk1x2edlA1L18YZAFj3oeXhP
XMTqNq5kBMsQw7mXLhokcXVXIHyQjE16a/su+q2UCt1C+RfiGgD8lqJfuolaxCgn
Ber3V8Z+yP5SAi3/n36n8bvZ4gBG9kS5brH2hiEmxtwzPWYIUrg90dpVLUm74rjy
Gw/SJtZRHCxvHjHkIkqvEJbdrF0xrv0irNQIRzCGFwcDccZVsskdtUvwXAJCyD9z
i559o5FgQVxn/Krm9OO55wES2BERQbwYnk58GCCAFqDQ8/ebQK0Qq8X3/9Rrzgfi
NzM83VQArfvkVExKmdn0Shfk8JnZl5erGxPyb+HMFXj8+8MKjHKvUgWo/ibL04DN
4wMPSfMIDwulDdoM5GEnY8ebM1ZUuc3x/Bu8QzbdbNj0E93m7+6iWeUDbFqqRytK
4DgkBQxRMHArMj5gbOB5Os6TQrBXKbbkwUY9bo/kO2vsoysV1b+IEc/STzPzNXhs
Cskyqxu7m74pvOx87lXartfFKKIl60HsI36NzofNiaUPMo0n5nAPVFlaGK6P8XE/
bg5Q0gDKB6U94GmTylWmlM+lYWJku1CtufXCjn6ZVrcOLYhnS1ifN+zbh1jgYMyd
WosV5DzV5df0lz2buUhm4jeBVdurjIIoTuSlhyS2OSzisjvuNb4iJYFf4QwegHms
9LJmiqrYyFxCzbZa7DRYX9dEhmgGWCBbnFXOpdqrXYUrVb39n3+cApObw89lyYdb
eev6dPWjGEYh10mMrxkzTN/w8Jcrh+H3LOtopXH76uyz8m9qOAHZsGCWCNwZgwi8
YrpAxxfo74XSRorNoBN+haOXlGc6JJWXCVnr5aJWX6lkmD0kE8Kdyvm6+7Ha4As/
Kf0e+u+Pv3LlX4mUsJDF7BAOKMQSnsklaGUoEE/0QofMGYUWX8PDO5cvt8aOQK9K
a+ckTnJN2abqZ2z/+VkJEQ8BMfClGs+rpkFVlqQG1UybXFgRSbRHu4R3hU30AgcN
V7qDr9bCUERWrCo1nUgskVLRwKHk2fvEyYL9DutnXPJwggfg1CA6ldUqHScRr3/5
wFL1qmXgxBICatFZ9vX/g0j5TActZIomQfoe92rSezGTNF2umMqOD1AW4/7jcVSE
FYLRR2vZ1o3XruPNi2ELq56h8ya/ow4GXcGfkhPvhbTCGMgezKQH8+8sWQmcx4EB
zvXX0uqIvVGR1e5kJPl5LL09LWKunWfdgMwX2vvwTBpPRtarzzk+bMc+U7Z//I/u
9iA55xo5mXdPp5A70LDZKfxH9U11bfkcuVfehbzpETekDV3FTXD9posbLI2YHFVU
jzvVberoE7WTSXO6hR42N8/xtDavfGt5c/JHWBWLl3ref5xNq6t6rKY+ZdRcGz8x
9XoBzI0z5cldVuORvooemAYXtmoY1vwxYIUg3lfO1Oj+/nLCTWhDlUxx7QNmuopM
qpru+vmJsL3/cn1MAXYnYpVozpVQ+uOgCTMRU92KTm26awW34PY88WdEqOylBk6I
Y8f2YL1fVd49dhA0UqWcX9KpAks6q42D3hBSRnI12saci8M2adAirMuTvi3y3J4R
p0Z3vDkBLofen+8hJ5g3MnSJHV2Yi0kUl3iyQnHxMFDM/FeXI0YpG+JkYGRJJSx+
p2izeQ/KXktvQOzjUHB/BMfD5wW66cFvT3XkUWclsvhR3qUWoM1wJtnrxKqQswOy
2A5lceA5tIV5mFB3TUu69jXnPunQM/NI5ZmNX2xWUBQNLA3iIaItpFUwwDzjQGV4
O/RwI/leHSt4JjrDDq9ZejqI8F9DfnmiyDd9g6/Ygad1UuX+G8Xrnotm5VJKPPBt
1e6M7O38hKC9NrD8lt6B8dJrO98W+4bDGtXehRica0LONPFeA4SCOvjSDaM6/6wo
OEMMjYUWNnTe/mnWXYkRS1TaaV1V8k2kFYZFvsybcQZd/PR03n4d24U3bGBqlb57
ZLgC2ZPr/7irRsWasMS9pHsgInYCgd+gz2YGeX3BNYxSMlKlycvxK2zan4vVhSKf
NawYBTVocN8kUQGy03gfOLB+czM6ZFTrnk8iv+n4G4ol3AaxO4DJ0j3VXPc+DPeL
B7hrsXWSTrZZid+o90egEXl1/KjI+B5TvtJ61F3cHsxXWxKjCyHs7NVn3mRy2DD6
bho9saolpFS71/e94UhuVc2sUYp+JdMqwsEb63zWhzbgq7RQXqrxQCDNs6/DzO4R
LDYLpnXysUV204NnygErud3J3eVOIzf9N0f0Qb2B9qhc/5E1UvBcf2d1om6HenQZ
q7+Y1KexlmXW/iCxbULrPbef+xfYfpzE/Nof/M46/2irmFSEVad1YjO4wfKfnmlz
BDNOr3xaPb+0tJFhjUrtl10iCu1CIqeJvDlr4xLy07Cz05N87++lgy6HRsAjQz1r
6EFlyVWgp3AonuzNUemrLG1nMZVkSIo/NCYOJMk5PrxJFkjhggSz97JIiZH0ip9X
hG7da/Xw8vRyoiKM7Lt9VHJFehVtd9KeYwyPH57C97QCqMX5cEquMNsCZ1haQGer
06Gmz7EBbcfaj7Ef2DRu+oGXLffbOf2+nx+LiqCkz3pmvFEDS7z8PNReZFagXjiO
c7KprfnlNqPvcFip213vV4gyofLk7Yq9b4GqyZg1JGWWqeZ8Jxgihg5ZiMCNtfFa
PDu13R1c3dQ/6bHK4yTrEc89W+zVqYBPp3khmwcnVhfNKWXxzjyMqSB7Jy39L1Es
juwD1rKxebcPHfgfNN/LXVUeudLhBbMpTuHgBq9jKz1xfEGZOhJ4Hw5lrZ/Q7Uo/
B82XXt11XFdVx74/Bh9agFLGlJTZFZOdwdUtYaqnmmDqQYgHkjw9ZMSHZ8L2jmBl
W8EOX0aFpIvNQtV7wlbt3nstcb4hfoT684SS+ryXvk0rzxZePwSE1xAkyodndNOc
7vwety3wuauuBY40OLEwDSD5CRVzpbOUD1tmfWHPCuyjJgM+rEHvScqrGY/qKkHS
DKgcCjjoGoj42i7h5HwKi3oo9X5C5NiYYgLKGKwYuIuyKO/9vBvXt3LhzTe5Q9mw
73mxWar88bvm5YwPDhqDsBU41by+l0YdJ+cj/3pDNMaNb5g+HZFpeg9Ft2aGkCC0
gB6FpdVnYdNIdit8ArSY1SoF72EOyxGhf+y/lEUP5je09bxWUISWP2kz4GAYUNk5
HRxlZaUneCQxnIYJnSVSg2Lvg+gbSJGP7SlBiVZG2Mr2h8kzsjTs+Hv4k28vfVui
ugXhXjBw3GM5hxZE73vW2uL0jIRJJKRK43ErXe2UV4MgpBD495W2HN8AHi9EJ2tq
j/IkpOFoKNbWEincjwxm6hWHXCB8+6JKg8jVMwoAbo+GH0L0C6r296vBpa5fuw9Z
vYJwHgHXFIH03OxC6YnZbZoqQ9VTdex0MKfHW76aDjfoHzieY3nN0FYSCmGumd+p
nw1bnLybtnvspqU4P+l/v8aJuJJtb68fsIYiqLi+s/npsN8ZvNQofcAD+yVTdEdb
gBqW297lGFnMbD9t+HomFxSfRnpSwuLV8Mxe98FoGr0ludnthRW3z7d3IvOG7PJO
+NM+dVSHroF1kXnZY17heoFDaQ5YtgKZoofdPVpojCjbjIzsUQ8tVVmFZFdMVXrC
Lz5Le5Bb9B+rMvsjeimol5xgawHKCtAMtLX2iAUfyeSHwC0AEkU9vnSWtlHk++sO
Ewsh/ScdOTtRDeW2uS4s5nX9cSS2cd2OXwFR+MjHzkzupq+8xSRf6bAwBquK1dC3
dz86Pl8fa7udEBSSdAOL4LttPsqpt0Cxn/8E/UyJLTmtagkDwUnk2NL+9xB1nVRZ
RRSCKy6FMco/ZQuUxcKx8+PObYNWaJnaSZwVlhLBRig3p3emhNKT6ucTEKYjBo2J
NocCqbElhQTUOk5sRj9MdfhtngF3+O2Aqwqr6bfm9KP2+kouAK0BicMYwTex1TpV
JlyMx+R+np0cpJ7TyIWyHL36+PnIokEqjoqfZ98zP8gC77cNwlnHmbjEo7zjRKGV
mHoFzKdbOdJ0ggsvPKa/h0K6sEHYMsuCVxBOygYhmFpkv2bvuDf4284kGkDEhq1u
i1qyFlZGh3mom563sQ85j7+0pbMTbrrTlltmhiDbYwW3YUL7HpMA+AO1q2gboKO8
+7wGABBLhUahHHQ28hZPbD+NG2yauR42I6QozSFr6Nv6lU+AQ6H3nvEueW7i2hx8
DDyx+Bl40dtXcVRJjLQ20i8HX4GM88aZdbjedPdYGlwjOm7buJtqCiBGjo4Rxw53
jV76o4XSdtAQeOnxnljF524erDgcJusGQg4FTBpdc6OiSMOf8nYW8NOkeetqHdjr
Soa+Tk2c0Y0911rURrgDCVWPSYCkCsrPgWqYJlUbfdk9YSl8Vd3uerz5pqnuSWuM
7pY1pNj2qvaSs8DcJUSc4u9MgKq3P6Q+IMAgPxQLDfzVdDscDE7JmYlTBqQTIbEB
yLZhD4d4eFo8ZDm/kC0v7OAJUjT0Tm8ji6ypCRsbSF56xjguSRIARePsKyzK2PyD
m9MzaNMQp6KmkJHOHFejPORytor1fdpBnvchOXsvqMJApik/N964/AmcHskSU1FG
F802obFUkyVqGXklVnmQn3Azk77n/hWbmjFhNA8UPZx4TBlVdQcKOrOKJGnRlCjp
VJrRgnMu/DOjrSdpKbFnoc5lsg6RIAiqiPsPWzwwo0Ic8BzujdRt+Yau18CMwsjh
ZaINP9Fz22acv6Jcs6BJgU0VDpmWFqKtJANqe0H64Oi1NTBUghD3y3AfC8Oo6MlK
mX4FBoLqwo+o5WPfyAjm2C4a0xb2zNm9MYkq10Nc3VWfk4Ukgo6nk2N6vlf1nvBQ
YuhguJN4Npaj1tzqkeWKvbh8SNeqM09MZ5844EJQILXDgXXM7QPIY+WedCPl+c3o
Ao8Pb+vc7Dc4/rfJWWXsP/Otv3DFvpmVYK0rsOtyaDB+rCjTmetC70JOXtqKzDy2
FG1PdPCzX3+s00h9BqOOIZCw9yVzc63Que8dEaMIvkfsi3IfdJN9zVenvYsp0kbM
nhWyfAb9PmP5lwv3zGvQMXjV2zyLN3n6cfgwXvj35jmjxCHUeM8IWWUQBb0d7bwO
ST7JD+roxNGT3ZZoEuzXybvsLUheU6wqmBg21pI7U5DkG26DH9WpZXBhIPQXYuZw
/0/0hf59eGfF35tnvUMNcZGC614RTqdNGNJGfFFsVgBSQqCZJCQK+3HWnnI/BdoT
0WsBb2yU/LfrV03O0ElHrZ5HeuXFCzzqXHMpzSkGIUZmUjRLA1k7KZCo4iGuWmyt
YexCw1iucWF9yZ0tziS1rTLOGc7V1czWrDFBXrY82Zs2vZtCBUmH1e/b6gWYiYSQ
dTHACGFmFFwWOCJfzMf+7Q/3fqqRO9gTP9p2YQNJBT344jvug9HKzdZHjguBws6b
1oiE68lk2goMJx/RmgjYJ8Riw7w0I7bQO7/kDeVnD8xM6idg7IphbDzIeHS3QSUC
zOvTPVEr1wMlRHL9Hg0t2M/rqhnL6DuyAFoPo9QOrmHFAagsL/zk8XtBn2Qt349E
HyafzxJJpEDrOGoL2Bl1JNfZUUC1A89GoUUe/tOVANUYpPTKo9X78H91da/KncPr
eyWpwjsYT6cWINy14jnMGGBtF9OzBvjBNBkXDwot4MGaYMiOpPJmaYZtvmbPs0CW
hBN4c8RwPLDJj3pXkezx+LyLGMflZSWzNZuCqLnPBcf/vHM7doTpdOOK2DsrfLst
Hl+vNiQwFj7IGLiHFfPQloCn+ggP5n+acorMS/HHrfuwZK3xXUCo2m3JG8TvL191
JPXMoBLSKfol6ZF6ZB4er7px6bUwIElxCIe1LeXfY37WuFFhJ3N3vDgRI0FG7eCR
msTmLcHI8+LoVygkuyQ3+xOWiUnMtOOfqJtm1/E8duHFREOTUQKu10Xx16iTjZLR
j8h2UVAfXpizqHG8lp2EMMpuq88/XPKTq6rMNJmIwbZ/jcCOE3VX+36SqpJw3L9P
1cfft72ab98Lb2qDX07wKSMa195eRqN4ncDBV3WIDnxMkWO+XAYdAQGETDR9g0vN
5kJgC9g09+XZ62HnreOflxmOKIBzacMgWgKxQVdJwdSM3xKsqJIzM8wYE1SdBYl2
acmgNGw6ApI2MPwAQKhlfUuipsDwpKXt34J/jwNJt/FGc1iBRYLkEDhhnr5ZKS2a
1XhRIT3zFVzn2iPCQUfwDVmDxgERQJYO6yNdPQZccf/xU2w25Pu6ARLR7Gl9Ad5D
SgOaX/zvP4MnKjQQgUF8TiQ0shS18aO8HA1tzUfk4aSQvhpZDywY/sKSOCC5XHXI
mlt/aDxOlZvWe3+La06GAaR0gLNuqFg92TnIKLHElS3g+aohSKS3IIkD/twvLVrR
LO0YrR6L4mfSiFMhl79K+sB5KPyIdDaGzBdTltnoNdL0hOtVgYgnkWVQpsbrs9Bu
sec8kVGzrxAP4juuCO/yDAlpibEe2IcLWLo80v+wwIHl5ZP0l7+fEi67on+1qbWG
iSp5gA3B2QC1oHEPl/uAFQ7DQWwyqndSlNofe6HsuGBM8e478uwy82Yyd9ETogr7
2hpX43tyiQj8zXrQvt68DmiNBTNsMD3YKMno2ZJuICNRVqIyrBo+JcMG72w7RXxu
ICCwWeAfsvhEObCHcRJqlV6xRO2yAHMI1xtlg1o7q2LnkaoM5dxDdwB1rcb1G12y
NkSxivWgc/CULyQkhhvNMC3sttHvc/Abhnk5lKxfTSmoyuQ0yme/W2GpEBZxgM6L
xxRrD7WPvZs3YQ6u8/frC/aembvEdpIZIDgpIoiPCOCc6tM7/x3OBfLmY7rmJ+qb
nIfEVYLkaKtj9h8zS6gfyHuc1xx5Ukni7wxUQhHsE8foAX32r7l/hYdn1JOPsjbh
cwbHvPH4H3rwvfCUygebgkThAZASfUQPNaGhRvXGFgh3Quk+FEimyEd54jMf3Hc5
BkHR9VIXdrirrr2sVwBiHZ0KaFSA9c3XXMO7c6zdTUHx1GKtoGibfAkr8nYDvTXj
dx16c2G38ICTvpSZL2U+B5YEgialblv28VvLyvwLiimnzTOSHAQAAuWDQ+gCDmj5
+Jdjnjs8EJqytZvTyOhI7Ms8QdujTwRGgpKSHfXVUQNN15GkoPeUnrWabP/CGuWS
Omz5EZXRgmcYc2oN+9Zl9V4VKcUVIkfKFi/WZQQPc4GWBcOGfPAnI385FWDWZkUl
B7xj+eZ8dxwcnUD0tuv3naUXOEAJg2SkJR8gVqXe4O9TIwUPXdkCOAuaLvVuYPoH
So/25o9y4DUR7z3RUThGShNIo820hsZk53omOW61ksqzQU/rkGXVeoHe6vtYxR4r
QJWypBzdQUtu2Fec6g37t/LcrJOuQ3wba/dp9f2m9aoTqdAizLsElfgK23jE5bDV
IFlfqtLa/ZtJshbUp0UhzwtuPP3o9cR83bEnVNWQwgkNPO+pen63WurG7ZXHm7Bh
rD2g8+p9BMxPhwWAOMU5br2fh3LwRGEzqiDlb8vFGHFR4q9aemcXCdgCWlrXiyJ8
vZIwVOSlkx6554pRk6x3rXa7aRdIYIgP7dgxgwZeTZtw/+OlSpuANmMmndAp7tmU
C2Wkr5GLUJhKpha9z8dRfgxcMGwgkEtoI2X6LkE10wmHJ8sv486R5WpobI+FSzU3
xyUQeOVSmxgR5x12dbqeLRyWVWCHlVesybMUuI5Q4ZBDy5CTYw81uDxxhx3rcQ0c
vY/lmtHkW9z41CNvBX65nSP4InRuV4j8OCKbedLJU4zf9iOKzVEE3OTHvKmGvbqK
I35zueThcnCJdH3Zegtv7czXevl+T6Ct/cKq2VZEBm1kpxw0/9EaTi1LDStxBL1L
mm1GavqeDxq9UIEO8YtETx3un/yN8QZUueOqvPGbg79kVZXbFaJTtF5POToSAxBd
lny6tHPhPKL2F7OyRUqSuamgHrn6ez/MX+lZHAEhE4JrjWzXA1GvruRD9m5oCycU
ylz7FJjtpy8RFXfXWLooZkknpOsv/PT5AXlq1nxOzJciyw3mz/PUOAM94vTrSGoY
Ugb5zwkaoe4B5tWygCrunmZYMdmknJugTeBUyA9+vl+nR3vX+3Ecd2P05xYI5WlP
CZgVA2gR1nWcrEMU0x3bBmF/KC7gJJguufug4rgtzKPyZaAuQVfGKczDrCRSo09D
IeEIlC7REWtk/R5DMF9qbEsjr73241pZbfyHJkO8fVNGZ5gNFh6ZeMsf1unzzZPs
wVyZdb/fTcsfwCrLcl654SiRYpicqV+bFKdCIOnTLmbN3XXTaA33zV5sHxyKWong
CLiK4GPVR/BD4du3uBVBNsC/VzgqdwrS+g6A5uiosejuYq9CPyjkT7+0ITOTBsWA
gbrRVT33DMB7qlOiBFR7Pa1clIkIk2XM/JRjbB1v+rU2PXpwoJyps19fBdAeqxs5
vbEg5jtORZTJBWcSSiRR5pi1hXVVC7ZHXPM7mmA38EHekm6qFDJy4Fq5enn/F8Oj
6rbGfKy82XRMhnrZyZMpKYeFxI1HkuzGAG4oV2UML9E32LEiSXmvNKWEQEmLwjdd
Eh0H0aayqW0p2jOO/ZV7v2mh7ikZUe+EaELeHreHPoG3VIioPGVHs6GlxBIRQBKE
RpJ2Jpgv7zZTo8eMAk27evsbyF3rf+YJP9hCBocys7xxNx0S8wpJ7Qhv+1xMMMEn
84GBdeh8LEKeUsMGhxsNWwMThAF/k49WX1HRmzZWDjG9wknIjfcuRqQhk7HeSe4P
Y3/wdAZIfoB7GhV0NiyTKh/jlBsmJfWgR6lvPLqbjbiyEIcc1iIIIS+JmpOCjbyF
Zq9ZyjY6MuZIMtEpchCkSjHEpdDFXRY2RcNhltsqQ+vaa/jvir2iwoX5gANZfGfN
BOje2Y2lPKh+qHITSM6XQzhfEvvsBmXqoa12UhyaPCUSa14N2u6QxrLzY7q8gJfw
ooptfMoMy8VLspi78dVUlxYb6umRi48CpH58l7L20/xjvEgol/eZ7JZsUDkNmcKd
8QJcS36fjeqvaImxDohfjXqVOEhMbFq16/Q4s8hzN/aU0q3SGVVkBIHGd4ZdHSQv
AvOa4/Uc6HZNMjD8GMb4gtFiRo/xrmUhZ4pZHYd1kxnqSnpQq0DQggNZxLM74DAW
mcvX+OreXLC8JT0bUhVMErEywDUc/p0aEu6QW972MFgS8TZ8SVgEP24oL1psLU4v
1zCBpLjTCtpmxoXzY/4fBl5lyyASw28moQSmowwnbEWr1Vdjza3fLY7ciYe+obek
inG8dony6ck+Fz7AH17dqRMA2gycsJUpwUWQk8jK/v0TDaPIINUIajcRSGI4XHEf
TY6iKf42wEJnsdQCydhAJfhklFEbaxt7+OZQ1mW7HscgEdjPyeDud6+e0xlI873W
ZDFt/0cFE2OAkPG9ebCY//+OX5CVBqP41b4fYIB8KxaC9msCUMLglZofvUy5TbtQ
TnOSq97Kn+LwIU5fCoc5GPLwmoN5PKbG5W0FPhs4I5/2lnnMaQt5sJrfAmke9vJr
deir9Ywmc1xHFlZps6AcKN2qak1CVCkShJkCV0EZhNHaBKjYMsYW6D8AkNoTuK/O
zg6eTxareYIUpZb2ejH/0ORRga8jClZZSOnUHxh/3b/MA+0atBtO1xw01mAebP6v
pI1wCRjMY6Dsbr4qG6zGPzW00e5MYi2DhdWe65BWWFn279gprr9RwPrVVmP1fYgi
xncUyvLIy/jbPjSjwCoeunIkBgon+5WStfN9MI8719Ou6jnh6cXDiT5Ocj9zsL+N
6a4F5Wze7o9HuxGOa2RIhLNz1Fu8TDY/hMMWuVaySlfY/rHBfnoqlHzTaKN+asK9
HarwfDIT4V8HoDjuNDr5mOXPn0K5ot8tDFCAA8P2WFtLgyMvayyjIaCl9a/R1k/b
FVoB4fOFMPnilze0vTOE0u7uOvj2yEW+2J4MQ5zHCNzgp+AhJMKZWhy4Xf9bchPx
tmEVknoAosKfl9tRRv3m6MfcF5JY5hUSqUwk9+jh5KVWMb9L/anKA0GtkYsg3YGL
X2I2YfEgaQEghwxLAR/34s7vNTw5OehlXQQJOooLAi7n77Xoiqe4lSDIAye1XoQc
zIjvifItWcoyqx9vZ/obpsNcXYPO91ThfVZ1RdCsKWl57eHvKPaRLmV5VMnph1n1
fINAIA29OXbS5aRdfF8t4FuTF2EC2/vjDxbmnB+oi3XnfUoliM32noo4acqolS0a
lhNKZOu7Mu8kiStVuK2HsGC/Snpqa7o4lnmFqBe0I4qJZdie12Ug6v4UkPu/I3HS
g94faKaA3H4uElyb/OWEaC9Le38rNrBAhHoQee5ZNyGefgkQpo1KlsQfgzNa9q/C
mmsDBTwWyYkdVd+WUckjEQ4uNFyJHMK9qc1lScE5VgDyf6QQJiez6HI5/sYeOj/R
Wwvzjh338dY1/bKc+n94eArmdUtrzB/OGa7kT9xBUL8KTYTnx/82G4o/LOyG1Lwl
T+Todxq0ByG/OPxWywPRdENP+7GG5F0sdcRiqTleEHY2ORUfOhmNVQLrvCq85937
voiV44TPEYMBb+D9U/vuOHYohnuHgqNtDVDNHRcGebjrJesHA/2iXfoUoDarcxIR
f6NlfyEoI0NovKcC+jI2HxWdzry39/rcgrd57qazQ6abAjIXWKzKQd0TiGIKQBC8
HBbsNkCjfaE7NF9t2hhX5dpJdWgvm30BUEyP3P1vBmXDNl1HvRyO5QN55ueapIYy
OnPNZyr9XIezjr5xvaeGwMusw6gNbjCfS4MK2lYBFOXhf30dx795zJjSqZk4zpYu
5EOIASfG52T13qd/7YXOZg7kRWkUjR5LQYWDuGyG4bo1RXNWHNvVWKCx1gO2om82
rP4aH5FuiSuPz+427XdxJ30vtSgKVcLJLg/ZgvmwnKA6+rNytEz8SWXYtuADKGyS
BJ51As9QQJHuiFhjS7Xh0/9ZXR43Chme6gdKE68SmDc9/nCRIzdxcyy/pXARk02L
u7mgWRziSPUMtbIJCvHbifQsgbUyS9SsnLuyex0DrNaJ+CVli0oSFwxp+XOMc58x
aJxyYYsKYBAhsqCcalgm/v82PH+VorLCZLJbyrA2zHuwjL20LjVT1XAM8EetzdhD
a9iqB78UeyDl5bzQ+RYeFRJi/1PEPlK3bgbYEjCwv8dce3/NMp1d8Hv9Xwil9hhH
Jo1QPVqG+Pkbs1CwQ0X9YZPDNi8bPYmO22oWZOnNuYfnduCjeVkYIGxPmJd5UBg+
apDv1FAx8gbnxrhUDbjEv+iEvSUvTYkpVy/hHhhmsNywXSQEhq3wGi2A6TSk8htn
GatOVYLqoitJWEoccrN0khoLEbU0knJ9pEcN1lvFBfRJb6UMApgjTV+dEslU2Xha
e6STeiNBV1HQc/hfEFSFjVY516YTpzXeO3jZ0u+4fftc3DRR9AkmdBJIDrWI9e4b
kECdO1hTBk/NlOLZPR2ONkh2VxnLpe4kj04b8Qdr0QnXph2x6CZyy/s+ZLacDcHq
j5bCQopUZZVClJ9qqgFPpfL7Jf+UtfQehGUOJZ/wKUaNLDOxfl1+qv15GbjpCovd
ZdHm0mCcTRXwwh4UZL/vRq4XmdB06qGFtGjF0niQzuLPqYH7a/cxO3XAO0OqrKh3
VgNcymj1bcKTf1SDU6kQL09QeSdymJgezWvlnErUfMFuCu3b8aapwpB9NxoL1A3T
ToZbmnqfkI1qZL2V6P5OWOMIEniIMExZHN4dmGS3h8G3FvmnkUA/t+9XhyUTDQel
gqEE1v5K/ViKBAhgjBoFCAg6d5saFV4ONAZuQ3xYIqPoY2NUFyU4ivSPvjJ6OGGF
Gkmu3PVCf/pA9RJvnMV4E5PNU7cRK3hCqxDkdodkViXtm3LfH39oV/lC2wwNTA7N
iEVsbbulkPRLDsDRqHKgkYVX30Q35IVaqUN5i0ntzE/+qvBW37NWOybO0VvsaZkz
YyG2sCbSkJ9WClee9/58CsZcp3jdfYxD60l+EJiUP9D0viiPBOKT3PdbKex4kIK+
eghvgEvRBP6FUF9WmpQSZvVwUdeAzydoDzgEzVeFGGO2HKCD095aCsPUl9JOsEHe
geTNBJ4DSGnlHTrkUahTVXcO9qNE0OyikvnQ9cQr1bSrJVqklnTRaWCkbRjBMXY9
hb4FSNqsotT9lXa6ql2NZCIgJ+1LXNRAmvm5cJ2F0i1Ipm+KIbW9Oj45Izy2+58p
h/wS3jslTZpCy7ydCmgErBQcX/xPLuEguJzhCr4Z7oxZO/fWZ9y5l3Kpsj3ZMGVx
SZGKHDYwK793wbKiNF6nHdfKKk1jbo//BunE/4Ics9nXSkiZ4i1piDVmKOwRyDwA
kpO7hhKQKjeBSkln20A4mbFbbpEJlQSTxm9q3APVFSJcgORtyW9lnRwvIJI2msZ7
QHNDJphxz8rRXIG8uYvEa8vumgort7FqnaeKNMTShO7jFPrVd/h5alkA8bMUXAOc
FwzhT0SchoeMLJYRM15v6/AuJGS9XGP3n3IEUyRQrLgZckR92dfpUTH47RoRTWiW
N0EhmNxz+g/coSybR4SY6cKi4U6XJTG6gnF792/048c44EXtlFiQvB6iyVZG00B5
CsCGbPdrOuxtGh6//1wO3nCgOBQgkfUdXWs4QykcyS/DovDE6PWd9RsoTg5AhwSx
N65kqGfB8MQ/H/8cppOeO394sfYNKujgDnUZzdO3ewT/HIoCE54XP+voNL4XeI0J
4B5ui3Wpm4gkvW16iPAKMt+Lk0yGZ2mCmT0nVa+7POmXhk9HXjEy8NPNmZufa8wW
psYIRCtF6XkhHxHbbPvOpkMe9RIyamNBoZbL+TC0XEOKuDkhQu1pKF3FwH7YFr8O
D4ig8bQ/mpyXj5sLlQ0GhCgqG3hJ7m9dkxoJb/70S26tnAPvtAal/vkFswg29jyQ
Gz0PzkSV29DwQ8A9OhsgjuyLa9kqjsZDEqso5Rsnu6NjKzsRhpwWrmWqdoX0V7V6
Zb1+iD/ZBcP3Wxwh3kRWaY6GDdyewafFhV0moZJDOA6pjM+FTH88xNjepxsg00G+
/e0mP7S+CFVOIu+M+g58o702YL2LnLqT0Bgjzejb03cZbB6oTALE90awc2RspfVr
yYdL4lZG0ryyRANqmaE17BDV9ja5Q6icEd88vfV+iPfrlPRt5qgF+YfqIyCsQ5yq
JSwKPR4NlI4UeaB73aIqz/67Z3ESTfcGOEOlStXG5L1lNfkF6LIyjUlk1QVWrF14
vxSeAI8T3imrjdlEPFwNRKHELbKCgYadq3IRwIU8joBZMLHCV3RaXfBRP1mTgWsw
8yqKY89EwFg2z/JUBSPBiYrgt933O71tKbTmPlRPx5ED/PqYfl7Y9lnYiJrf2Ro7
eHMkEJErHdBcqD729McfnugDFZMdZDEJ3+y8NOZFOjoaB89EbosM6tnWHgTWoPzy
Ddp3DBZ4o/Pmh3uUwr63ju8ypblWkUpMo26CwriSjI0duZcGgWHDVHz67Ko4w2sw
+7RA7WuQF27QqyDK2iu6M8Ta/FBLwrFXM64KxAA8P3ShFoMWkImVtF2rBze5RPAt
YD1hMWSA8Z967diUAcTvuKkWzCYhmY2fg3SpJYgIlJqey3Qpoj8Rr/PncHGI0M9D
Kg+P8pef7rlfAH518et3HmFsPhtgfDQtxH1A3YNemF/4wAyA2W1phUTC8t/N7L/b
agYtm3BUoLmn+GCbKjNZdAk1KIBXHHnCjDSTTwspGvZGnVjc1p3Czj/iMH7BcfNz
0Az9KqrjcJZqj1z2kK/Us/ozxlixS+CFAaAhQySCJD2suAFAvFSyicIc/1RZAnRR
zzRqRgScPNucLxIrcjVrwYkziebk9rymM0mo76A14k80/PjLJ7A9SifIQsa+IgLH
IXcB3eQ/H11hQRlGRDV3+yPwij68+PJi2gc7HrmmcjBIAK+Eyb7Iatp2FYoCkees
lcDZGhNQldm8GSXyf5w320qaIRCHj+qXKqF04YlTv9UNblj/ODQw9Wkp+R+nC361
3Zg16GMvGCAJe22x2wwaLUPtXe+P2qBvSak3HEAgxPmVOLgScPDFYar4tMbDgG8i
Axub0I89cXlAmbZFFVupLLyib5vUcRNAk31orLmSZUKQeHZxgX+UtIedXd3RRfkw
rNfGl3JNJJwtwKEWbqIgcyetA4PsmVIblCQz78NevH4VhXIi4B6LVffGab9RdI/T
yiUamqY2kOmrr+DnGZf6PO9G8Dd8Jbz6aeJlN3t1cwjB/ViODm1USGjwXixBJ+Sj
JZozkSUSF++mBj2CKx12deI7enbn/lZOhMM8kjUtYhZ/CphZ8t+WvstSbUFnawmq
/cAIgcmPrz0tx6q/ZkpKS1kbBEzd/uk/um8Y4LLGhphVqFzsyM1otN5jDNxAnH4w
8A1AtU+x62kvFOEKQvriVe26ClA4JVwR+MYs1QDh0jtUEJ5X5njFj3XduMFlQiMe
Sr4Emf+xxmHgqSe1IbT11WkBbjHbT7vEel6GMkoT+p0/frQFkNilXdcE1vJr4631
ArVbLiJru+rsDePh8CsHFIljRTZlF7o4Qgwpfnw8oSABIsYrbuYCPHHde2wFWcye
pmYfwuyouKMEwMy3A1pLMo2qUCau2p2hTCbuTtK4/+iYUPaysvxOidmJghyJ1W7g
fk2vLk3hvbDiDpBZgSHpWSyELxarst4yLAAVnfCWnjN9LHN/95ewXYtJtiow4x61
ZofW4/QvLeQsMfaNQiNjugquWcxX5JzoIj29Frl79Mgfrj7iRmEOnbQRC5M/Izjt
Vg40MfGcqlOMZANqoPiPoAsNAeF8/HnsnbI/1nqUH8r0LmEIDwZtGE/ktLGwttkq
jRoP8PflnJaRCvb/mlB1O16co1TvTqSy0F1IiIjqePoIRqzWMUmkMfQ+8V14PkkG
7nJIyu8Kkt8WKr4D+98sp64K/aGwA5vDUqs6LRgnP89yy6F6JNJM7O17Ia/D3wXF
ssg0SPy+v7zMOO6rA7Ov/Obusn3KN78bjfrVa3yq8zU+QQoOMM6Tq0wJw6GCmeBK
IJf1ualPWawhOhmePJKVJEv7hJvK+6So5Bq3enmxkjVjMg4zJR/0VMf7sZxioxT/
VexA383/xCzTJJsqzEk/wCu2ToPXgob3JjedQOXsooYdi5HSs00QJj1/iDfu2UCI
UyOj3lx7BhvrWOuXeXEQn1OK/JmIPhuYjQ9isNe//M7bq/MSS+Qx9YDgdIS0hr1L
b+6LPksLW5MsS2XPVC4la+CFurPJLwXuV9O+g3ocfcNiiP6P/icZeB8GGA/BQ339
nxg4AOl8+DPEbUiYJaHJnlkp4Zq87UzRE6pmkEzwthmIGHYqcCslyrWorgavEyLu
7yjmAWXfy2KdZnEoYqiu0BssxxfQdV42BnNAI0cPIMVUdmmb26uC8eJwcUvP8LXk
DwIuV9RKWIHtM/3T6bdUHupLDrlimsU3ZNVhWE6MLks8Nz2mbRX+p+twtiaXufR1
m4bSiJK8rcicU4dyuaYChUiqYLqW4GIpQdCyojoDGFqRtVDGBbdlfoY4aKwCylkK
7m6s7bHqkLShvOWWDx7ApLPb6fNeOjhTRJ9gifAgCwgARrDf0qRihxcAbIWplOO3
3X17xOrvE1D8eXNvG3dhyBxgwoql89mj3tVuHbuFq1AA5Y3b7J8fVBa446jM95s+
UL9x+UYf4p6cmha3B2VSXMHm9EV7x2ZEZ4rX9eGV2MuIU+uInjZZrJDxgGBTsZWO
PsuJFIulzvOvcYhVb5Em3KfkYN23xdoS9nh5EsqL7iTY9eaCfx8x6yxFg0JIE+L5
ypjJLo1UYNum3RmK9Y5ekVnWqm7xlLC6/tcZep1PqUeTWjeeEhvBYcdFK9mgrkLl
YhEPERvmkuZotr0sonHlmERp+xQg8DuON2Zgr4oQ7J3N77YmZhufcKU8TAQeWpWD
Ibdb7kexo75OiU3aMh5V7XSk6BrU6+HWi+Dv6D2ov1cmDDtQFbTqw+/FK9g1Pldi
Xttae9G371/7ZE8mBlf5Fhi1du4mBRy4ou9um8Hcr/x93C6D1LFggHGWa9VEDE78
mMgowZh9TpD/b4UmP9xjsrPPaYu2jlkiXY3cQIu68HqVOOEzxeQo0CpaUyI7nnjN
fVSYD8yKwdzSIn1aLuw4pUsIxojxvZmxMqs6y9JSe+REbl0OCFGEMovwdBs7LJev
CSSjXWJ6RKskOw7/s/4kJKkqdn6jtwEvYUvMzQaS5zZ03BuYZQ5Z9e6Icf13Q1JL
eO5cmINVfvhXE5CtEOU52N6FwOYM27REUZ09If4s6udlaC2JDhQYD3I+t32VUrTJ
IKmi1zr2g70wxhyg+yn9DUey7ZmCfFgb9Q3/O7gddvEW8ujFxmFUhCdnjTyUElUT
ZnTgwQbRHCV3/HZ+sz0EIwk3KxIB7lYFYYsJ9nC8rTS9r8TZnXHlMh0KD4XUgKhV
GiKVnFeg5r+NDcULP3g8Ui5iaXBp1Nn0HuVJUmSCnZLo39ts137TNbKHnLr18miF
7/QhHvTV4flc4IO3Lj2ylb3XmcnRESBFBPLP0yTHMaaF8t0f42gzrPSfbGt9bKIY
Jl3ZYNi3B/eEQP2ZAsnHuQTdHtvBnktXdB2dpGL0YSWucocPUd+JWXz+4wOxaPur
k0tHgjytS4+MGDHcf7e1rZTl+k5jZzonp7B9Zq76R9brLrNjPfMgrvWETWm5XQ2G
7mttVLc53gSlAmNw5H8+2TtclrgwMBF2qTdp9N3YCfUY7Iml2MhexgoBh9WVmaW1
AymNQxcrPYbZFw5w8/VbJ/sl6k/C1R6x6PjIAGmQnf+h4gCjaPwIjhApiR780+WA
BVm+QtShmTRZiu5OBJxW/8Hrm393t8jbhygkwgu7L0dmF1qn+FmPrqp0TRn8O4n2
3Rs0dgHlw96yjtZ/IazwNQevP582a200INMDHMXMKvv2VChV/gvi1Bvflsa3kUcG
UaxtH4xDGSWy6DWR0RNgHGwcXJ0UJlRRrCKeNRInRQ1Js+AiCDVntH+d5MnHdaP5
i+u+fvObM0MZf0xpLHh/E7gbdgjh/c7LvOIIx0VDB9WtyFxbiQIZl4subqNyxz27
cZutJA9puTeptKnrcZFJtm+VhtRoUBU681sllG2ERKL79ArK/7rk+gkSxikOXide
DVLCissoJTeKr7SLCE5XwWh+xuNkTHG1cPeFA9lxpnoHT22lu0sHfxaWLD5BFiLV
ly7TYb29eHyO15VvZbdMkvpIZGt1zD4+lvTSjvSNKOoxYnG/MREU1NGfKeM0e96Z
4We+OBeD5CbFEcJ+WX2TzzdARLZlGHCpPT4Lu1bjvEElDRu4ViNhGjmk1Y2faS71
NmbC1ouGHIThszACz/T8iLWLnL9VFuEO3sn/m5vu6cWnx9e6dU1VN3cE4RLZBkd9
7I3jFX9pBU+4sqATWw7IPA1qXCL4vt1Lp+pNUQEulufjPsx9hserKZcGzbALOzR8
Sk/3JQmdjli4ToXqUAy2HVhjBM5fjJ/rsa/uEAayFrnZZUFYITLQf/08kvh7JqF/
jp1hKIiy+rp1VvQg6qCCM8GzBcS5UxFbNrc7N+QYvD9ViMzwe8agsB//m6MDAS9l
i5vtImNosZs6hP3Yiwh/jY1MZFWPI00oMFLP+RfsKeyFXDePPXy8nq6hTHFfD1hY
lzo/B4TlYY9E9Opw4sea622QDWD7PSwenooWpTY2dv+vPlE69iJAtdssweSRWXGn
mOUVD+Kcu2HZ8n2C7DJ1z4cAu27vfO1aVI833RcpaKDiafmMHyb4Tger0H3kRBUk
NI2+w9pav+OcqdV9h5WS9TI03rBMBRkwBU72+ZCiBPyJeyd9UVgx0Uh0XEBKgvYb
2iuxd/i8WCyI9DXdguQ5/Cgiu344qDhyzUJpJsdE9c3CxYQ6KZibQSaj1wSvfEZ3
6Jikqm8nJ3VYTQGgd1+cYAJkUeSQFYfjRFg/z9McEj/JqX644GfJihfS5J6Kc7gD
rdZML5W8FzgHojJgRwhAxwPpD+T0eWd0a/m5ThwwoO/iny9WglBteaY6jQKIhvub
0/GWXkUGL7SWPcGaI+8aZmBwvnGPgdNF6M6rTDbn9WUJOclQCrEgsZjdCCwvOS88
U5Md0evbaOpGMUd0o0qx7gCxtLZJr7UFdYZjApsVUTxCc3Oc0sd+zGwmjK2mTVuG
L7MrIXg2tSDZgDAHbjY+we3gr0bhRenj0bfZBsngUz5SSmRj1hI6XtB2pzwmgafq
q0SkXX5CUdAtDSOHohn0Hm1tJZITQ0C68BQ9KYttoAhI/ViwfwZxNI4DrGhakx2M
jL80AZtGQaD31fppytPqM5zTcR5NIt1DEDA6L1kYyRq0sXP4v29mK3dS+j8LSNcv
IjkCinYNP50ArL5yT24K0JIVCBEBvb8EFt7fs3YHd4LnbQQ+JTKUcIUWcP7LmJT+
Kxe+BRZeZq6yf4zs9Y31LhgOTj8QbvOxYNBfYrSShOdUxQ4U8tLgK0Stw6WeugCy
KCccXxLeNf0eZHnpj9IKvPDR0485PFzJ+DBjZwNJcGKbwlf/TeXzVsEyYPdTfxLc
qu8/kqSrzDIcSvG+By9o/Md24sH4wCK6E6ONPSOYNP65eB339EuyPDRLu0to21xI
frRTf8UfLTKSCc9qSQgY0RMCWONpMIqcUYOmUENYL2sLNva1GTeENRnybz/l1kzh
3BsQJb9xxknXd6zrKH0rTXwtyD/ursrKFcLCqnWyFtpsae1RSejRZ/Yz7cpZQug0
VEGGp/5ESerh9wfTbOI9sQ8vFdNV6bdiD6S+QtglQC0vFvZZnwEG3mWziRp3V4rt
oq1VP+GpbBLyyxvu/eoa3VZyK94zShhx8gvXNwroEhz+n90MN+2HWPBypumYvw/S
uiVN0QltMiP5fAdjM5PEXSb/kLdRB1JEQF0oY/gRYUL47uN14/0x6hqzSunz1fGX
dS4dVWGMg1YHs/tif+/o8WYhvUg4M0OjuNN92WEoBgDsVTHk10k25cyZrEDGGLGL
K95J1NA8h73B7hB9oRssF1IeUjpOpIloIUVVLKvh8Ct9PoWDcY8D5r1jmP64oBiK
InWbhZxPrVmRNOA5ciV2JNAODPzrjUUmJdn57yqIlVZS9SVylrN90OxbYRXeMRBy
wOdy0wvgIWaLgOGwYWZOPmBWi3qjTDL3JCNc870444ztj2kuLCFNYyOsrLKSgivs
PSgzJj6AmTww/WJPaR61o30tFwxZrRYadem5DTTl27exg5dL9RsKGCMpm9BpCs0o
H1i5bqQ2ih24X57fbScF7gBfws2IyV3XAka47EKPuhyyVTOQjGon5fEOxoymo4rI
adD0WZvlEpyu6fH9AMT6iLxLway+wXXL80B+NftiwSsvvmintzMNH75Wo2mUvQvI
2SlRn4k8uEMHlcoZR58LiCa08KGi/YGBP3VbBZfifGVOD/JbQiJANn1GgGdpXhlp
3Jl7sgzEcb2hXHXiK1ijDX0KYw7tLoHysbm/mF9zhlGmKEER51zsmm0W1MmMy1oM
ELfcI23NI7iptRIjN4bBn1BgewQQvR+ArYWjSxSLdrWk7VgqvfsiAFXdX73RiWP6
ly1kFOZnVAjPFy6bEsC5voxJIdh1zYj9q1AzlZNc7bqtiI4O0JjWXFBhr0AOVIx0
ebxMOUK1+AHGX82H+Fsbr+5jPPu6tF6yoQL6KGqFeZnjwukVmBCMVNzXNwU0FqE/
yR4ATFDBhCkZ+88YNo2gBy4rrftumDGlagyOJTClQZA2s61tWsOL3BBpSALouGpZ
wDaO+Le/0uc+pA1PoRC4KBBAfiFvXaZoG+IGRJISVySZ+C0Ee+EN3/CHru6aEBiF
oZ470wHCsG0WFWWSnK+ObI0Nd42diZgFnOCMNjab9oWbAQQWogAqLYvjdl75faUX
exSj1thcfshxwt7IyJfhS5QpvCCP5ZCCHyLX8LsiEG9YV1xcy8ccW/FrrJbiM3ow
adeWF8z+uXhgUXFetDYkR1R6NK4HQ2tepCKoVeihLe2mDPrjQA+RlOW7X7yoYxqj
kXDFEYXPpQZX3+1Q/TLeH8XowqT9bMDRK3NexbuiEyLkrtVnKSnPvEvZ/AW6bY8T
7Nq1MXs/qJgQHbC7eLN8aQimGMgixxMT8pS0wxlPv6O0vcvfTLRJSNvDk/gmdqQI
LGU4o/YTyN1v99Wdaa1I05dLW/KO3FEEEdBxeO9nyvGwpY7qeDsL3XmxARTzr8zd
zoVqDuDJMK+83i+ONU8k9lk4/yi2NKUdrZsEsLK7viPru50Tr9O041YUMSNre6x9
nkKCwMePL2+loOCteFcHbT7O+JFjDTiji2WL0rlgJqryaxdS55cwx0+45m5iHHtr
SH5si8urloeAxqcWtLIZS0NpdeuplTDeN6wZSTG/Tvvsr/4w8qx4f1s+C1X3KX4i
0qx8MkZJfXbq3ftq1m/90mjUSf1Ln0Nu3YAZz++YjnWI7FBXNBifrWOU+P78ioqT
Yb2iFSTzrgAvD5c8ojJaKH0CFDXwiFWjOYpbudDOZlTpQF2TelOuTQnYKqLN9T3t
BU9mM8TNabeZsBtanSYpoBybJJJ6pxzRAt2qPpSU0BcVKcaGXZSx2Gl8/D1TI7Gc
0NfatqYXOsDZvgwoe6lbn65g1PeJXqGzvCIXpaR3J+1C8K6N1JuaD4p7DaRtmiSg
iQ1f6fQXiCqdhl7sEd6Dfh+sF49J+A51QpGCNTRd1Zoi7cwEHfkZZ0pn3au17x/f
2P+T/YwtC/rJrG8my2CzcZmJ9HgGc+6HqaMV4JixHRTouMpE6v9WxZjNXqKTKwiw
XcgXB6VgD7mxEhk8nMlVEWvXQjmlEmcF/WCL0kfdj4CCxrUTky5mLUCJUulLDg6E
v8MQZSR0y0yZOwtg+evrf3oSPMUvxxxSI4hHlT2WuA6720ysHf9ACLEC5AICEMkF
689DO8YBrWCUU4S7Gnjb4b+BuHTFuZMm0ryR2q4hNLnlmPKJgWCpqsXI2r9mnSeY
1+lM4rWMmK2TUCBU4WqEDVJydnmQT9FTEHBOETz8BoXoGNnyWH5+rbZaDg66ji6L
0udYdXSUD1YTsG/JUKMyVDu0qoa0gfz6ic1Ua+XTtTKzCVdFPP/BZ2xhkmbCCwKI
FLML7sGK44FpSjTqwZkIIT+MC+vDc0oDfwDL+8JTrbS1u9/gM68XPBE8vMXzV4UG
Iti4xbtv/v2PLIGuKT6P26O84xFNKfMhrJ1mVrh4Z1lz5hHkuwogIicE+Ep/T7ld
c4JkUs4U8KHsbQ1jQ8ayYiXkJmK0WuP0lL/BpXSkzwv9IxunAKx4RPSYKRj98fvu
hUphOvkd1hOCprKUHKf+I68BKqesiji8LefIFYlbk0VoR9jAyS1D+EBm2TDhkjtq
1Zab0CuxiayjlI7tjRauHoPHOo1oLQhyOkxfabYTkjfbHC2BvWu08P8X5yLc4pEh
2aep2/hb0JC8nfI96hAFtCSLNi0Iw2S/QNVEWFmG0toSewqkLYvm0W9c17vMfQfe
1MNljfdxPddK8apgMSt9vPMmL1/+PH0I+BclpMSsUnJiuRGBG2tqnEgP6FbbW0pL
kWBpAzdhbGadvUDQFZMWFalxBXOB4UilPhoQrNy1q4T6cbLjebauxbDOcmqZ38cu
4Dobfb767Jzwps9ZZFUOGiLB1xCqs5OIXlSPNCNCJv1uFXzfZM5rBbyWzaO/5BXM
erMKe93jhZ1euvZfHFTLJT3PdQHeocjXM89Kn6SVUboWzn2p+02ZOZmuZ1b8Ed11
SNXIfPbJxScG3h2ZmCK77bzJeWD9Fki2Bc22FKIRifOo9JYHlbDTeCXDH1wGZg52
5koulgYBwpEi/uh9Mr1JNc1+LCkUC+qytykhdLnS1trGZvyj5up5GVvMchEva7uJ
7Qunc8QcBOusAupRxN6t5UVviMRivbueBjEtA2xk7fIie36BTHGjZXIpM4/4Tueq
ES0DgxG8P3TFcmYdsFB0CZ6o2bATC0v8mNLgrJaYs2poXp5Kusz/3s/gqmZOQ3Lb
4VowNHwxqvD6Rfu+vtL2PS77ljSpB3RPv+0hbonjd+YK2giLFz3OAef8kVzPVm4z
VWsn1XESqK8PqsTJ97b33apTrGktItY5TSohsQciN0XCudJJjzRSscR0gY4vcsl0
7xojCi8gH/cXv5yAXTIRexxnd6YdN0Edbry/CH9Z5fZKXPU2TlaPWBDKR2qF2nrm
fdzYTycQX+l/3THMzX/zPhEaqi0N/AdQpfIfTjzpO0RgaATfxHUZmC7rp0RisksG
Ks/b8JqdG6S5bNISg4VNcyjsJmjgD9WSRcwAAMFTuXOYwa50jO0RRBA4vfiPtNJw
+vcc6bkIFvULU42ZD3jT8eZlf6T1TTesmm/UOY2+tzl7wMdyCJMNHTVWCoviXPcV
q9rlEuo2dl/yoDokEfwizQUdzEL+FD5WXVGniLGvLa+QUzDT9YNs6GaC9Gsk1SFr
oJUtnDs/u/4vznL2YQ+htaqIWZzq6e5vl501xWVFTbZwmIzBaO4GxMb5FccVEpLB
CPn6QwTwbcWmKGI/NCFqhtQQsHUIjVLXkiQBJi4C8m0yrYxYlOovgoGE5yN7elNp
gHov7f3cHvNBAlv46aBTpoL1MfVanlH5NWoSKYG8msDuOt2PaxNLxJb3BOTLxnDf
hCb1uwA3zNsYDeDBPg7VUsmCK34PwOHr+S+WEbiSVlOtyKsn7cSfccroqw4B1gVb
xhW6cFyZbroZww9J0wHu/1XzKuPtm7eFGyA1XHeFrwKjKt5U9iMteN6S2119KxrC
PEM34c75EFUYQ0Mr/lrR78rxqGJ/DRZxGFdPr3l6zmCFQdjzhS67ugBIKiNpDTk8
i0A+8JIbsOMZhAhL4OIY4dLGNHrgaSKhjXpOnfQc6g63XrcJEEe16mzCpMWxqf/y
oQB4xRf9qKfFjWfUAUXBsJQgm5Bl1bxkpQuxlvx7iIMESnVXPd4P1nEL9A2FgVq7
nf9b5p7sSkfs0R2MQnUUt1W1/6MV+XvBehwV+ORgqJPPat1SKQ6Im+wZC8Rk1VPv
9bGYLgAnnPi9mLHFKGjYJGJy6wpmlib50P9FU6GtxGhpsKMab+3Q4575ENTxcZ7n
yRknDTqjL5U6JQiP1SnijeKKhe/n9zxw4TPgHQEgCqXoui0/LClEF+LzfX90x6Ig
jvGYC9ecvw0oa8RjN96ENAhDiL0O+9o547SRVhEimY81JtbATCcKLDMZHco6pXuS
NVJdvsfnBqDlHn4oz2Oxk24Ov9AX3+z0rZd8Q4L+QsqAnbU9UloE5RFhzxlcv+06
Y9FobBOSaSwksNxGI3OvlLzkwc1r29LOP50cVJBNl8p+eL1Y00F8Ls/OC/g+W9NO
eHeXmW2pvWtrd4F0u3HTlCA7edMcaIm7VlUTn7Ek/EG24re5E0mxf28IIz+wMyPR
Mde6JtbUo5Fm/XjraiHq0wWF3IWj0FhcVaxUzoR/4yt1tjkhFdseCfEZ1HwdG9mr
r9q7XYFCT5Rg7a3MAJq4U4U0bU7tLW7jMVw6HJGpeGG8ce6yUmPmHKggGgzD++S0
Ppbgk1aT/y9YjClNbAjiyWZk3KIcI4eXKf95TRVq6kQYVrHkbcCEUMGieyI00NNX
r6HKXUcvokav7Fmfh35iaIYQ8cWSUo3K+s4Io6+dvrsdyu1BanAArZf//9JJ0DwB
FKQK2Ym+Kvz6O254CPF8UkIKp2VgJlxhogTqR9bot/nlBgbWFSWSQQEqz3XS08ig
RbPp1EGBbI7m+HfD2ZlolkPB50qhWhIyAnduETTMNay7qn/QVsVsBYKVVQ+ZDjcz
ebBsHAdXar1V3nzzMCWwWkPS5eH/9wj1yNs4nysEKOBrowcTTjorxvL/pZbYjQos
xfC3c/AM6MpZqOjxBQ+BDzoeofE/n1tE3RYOTk71MT+BKn/HS7/0jV5hIWwatLFt
I62S3FZppfv32pj5wrmeB2U2BPx0CKjQT9sBbAHIKYpI7dVovupT023D5roiNSbp
ppsmj8zeNS6/lqtvPKbKaEf66aPaklwfL/kHx6z5AiGG8lOvVla+BFV3e4M7cIOA
GdKSQn4EFW8+TgW1ezIM5nITcEu3bmvjRFN45Uk9364AdWuEhdKW9GKU9qEHB46s
p5ZkE+lBNbwPUbwcE9tfoKxgnbj6NF53hGyZKWyiWqzx1RSv3YdhNoh5I0fy73eh
Z4+dHdZaiv714zze24KFxPxPjAIyxS6R3LaNEhQDih/OxbwiCYHDGv0GdzMKgxMv
NMiC/vpgOO4KlIKcG1pKcCd1S6sH9dYWQ1l5B20alpnDtxm82gZ1/b6iXNFPh9rS
FFkER1bZp+BG4qqStDaWv97412q5aK0b7i7QN90iFe8pIFLaUOIB50Nw9yLgt5t6
vJcROoBaWy/Ai4oOouX+MM6aWI+TIUSKxiYiR5HQBOHSlD29IEf2VGcOG/yiQ88K
qyAQQ3CrpQWcX+hov5ZNe+xOII9q1mX81w76og9Pv9yq8q6k3CswANV1jreNn4QK
+fL5u7Ah95UuRtX1GRD3ySwTCirzna2KTTqRpirFjj120VutK1A/M+iCaJyCBPYu
Jl+ecBkopowBew+ykUEn0e8hZhiu4ovehWNDOQqiYIFgu411gA4JNYe5AwoSmbtf
08hdZKuVxjFW5d6RMRltxs7XclQwNiJA0aab94m9zRFSf5rzZq+UPwBjBTX17vmr
f/GvYBAlnxkmIuSaRqsLf8UGSAgmtDhruU6HOPZ6uYulbFbpYgvO02LmvSCi0CVe
2zWkc+xmC77pPqsXxr/Rl6f75Y/eprEhiEO8eoKbFE6LPYYwN6b6vQtS292eNhWy
6m45Cck9IN5Q44MFP7DDWTXKiFdCxRhOxm38gYxL16kUjyT2StFFoMOjUoI4XqaS
OCWIIawmyf4pOOVxt5HvanpRW8omPVNR25HCBsosUzciY9emN57DBpsfEUG4C4Ce
e33nLa92OW4PMI0jKdwaosJi0eIZT11NIbhd2yRbcCRI8wu8mjWkN9Lneb9qagVl
K5Kxla/j9s0tkNk5BRUi/1rIzANW+MXqVJ223fsEStQyhDPEOjzP3sbRJrmHOQkh
v/M1gDsReX8YiZgZtTO5BihA/Z+XLFdmPYCi+h9mEbiMYD6fn9tPtvH83wHjWsCx
cAj+9X8kjLYwlint1d+K7nTFzjE4I4SHE+h5K8Eh8l/3lsuYiPCKvfTmMBumPAY0
dltNlvJch+BlJKHGfRpPIuVFdUpPc/LW537Ljdg6izX16yPMSSd65U+9CLdxk2Nj
ApSCNW1REqKdW9khH22AQSAXcnXGinmMSrtsNgEr+wHLe7tKZEpe4kwwZsZz15W+
sKhDK1MbDvjV56rYE7lDua+h3GDbAv85aGtB3sujKpHqayvsByBZZNwqf/bhhzOQ
jNXltK4X5gAu66bPUbV5NdHNwPM+x3yzT5yM2uji3Lg+wka4skoD3/q09w0bRMXA
IlETMMTpWDy8CVOREDnKKOwKYPswkQGiueEq/FDanTrugJsY0h6zwbZh4cbt2hb3
zz/b/cvR4cyk+Y9JilWCN6EbKEiPyQ+1KiBFR8LyKw0YaqyNWeL2KAdmph+dWHLe
uV+ctYjYa+pb5ATkGjDZQ54XZhSOvh+a8H3xJWrEs9DxwNMUMcG9iV1bRKDp74Ja
T/OwKY29x9g8qvFgs2oNfebR7dQ1VoupyMPHK/O83yuRUtHKl91pFppfAEmZM1Yv
5eKTfA/U/x7vY9Lfa61SnrCYBedmHdcaQAPYA8sIZE7rkKtCLjAgZm6D4AkZYHl6
EuXqJmRi+N2GFyvg8T7Ercqv6CS+omxa6QFQ810LwqkKnnkInKxQk0Pv1zZhibXz
00HHvOcrgppfjrR/3+jdKzC6lcPu3Uact3vJpbDuTlVA9RVyfh7LoNwYsvSw9H7I
AwIsFMdrdMyX2q4dYF6M08ht2VgqquTvPa3NduoLZKUON8pkeCZchRXTUySvaxlr
+29tokBZZ8CrHdZnKY3UnuprEGRe/sM4QboAAgLBEVXPKeCbcKU9KaCzvNbytEx7
8t6jJ0sSHsgVzA1+NynQsgRKC3nipdfCasRU2dgfGnnS2M4IpmBnmeL+Gy5KKXx6
lvb0XYjMSF9L8fVUTgck74uUjbCujSMuUbhUlX1ix+iQ9PgrDRezoajY739FuGLz
lQOQjRtRy4at1PVD7AoYLbTxa1v9MfGK7mMn4zpAExOqKs5f1LWB0VtnNaBwvrgh
UYVsp0pHweb3U8dvx5aG/dER2ad++tkFCi7v4ntrrk0x8kclBNVaxkKKFJ4MXrZJ
U1Bcu4ORRW1eKTm1jV5RGUE/XrB1c3GJFuv+SGZFHs7KI3l2DRRWqbniTvasz/VM
u9lapxhXHSIpxDumf0RtP3fb2/FGhb4A3/D7JyzWzODomhiB/baU5gHvWzpJSv3O
bN2VLE3yFINbt3VEAxdeZ57C7T26ByqneYuIT5pXnFSeD569jfK5Eb9GL2/KFcBf
d52ljLoyU2LeAunooQ37HpDHRZR457pvUzOQW4bdtuYRjM0E6j76vjPA+6pKh98v
33waYqp2sE9OPfmqg2gwlgoo4ha5Hg8e+xIRbnrasNFmGBMx5lKt6MoX/2AOAF0x
vAciveAwzIuY8lQnFL1rn5fhYQq+xjCOn5A3eW6Mm/Q4Bdw/fPTwh9z6xZNXT2Nw
4aT7L21kSnu9FxJ/mNaxc8J9fMJlBLgNubd+dbqFY2+ayFZ7qNFCBVpkBTA4wguT
QTosCDJ3AydRFWVPoOeftrk8YSQCZ2DGbERQn1whUcKA/qlhF0T5GgJst40FdqJj
VxwlkybWcNVhz5qu/71R0nmhpkd6GEtCbgXkj6H3hFoagERWIHS3O7T9ebS3TJ76
8tDLnwbSa/qdjyZhvy0i1VqbxBQYuyTgZ+8F2wm5K4F+JK5yy6IyycrsBVNeuKoD
wZtFGkge+H29fbb6gCym1XjOjYv7jPEZesV0XL6UZXzomgP25CMwKA4Yrx8qehbU
w+MR1refWachLwY6lVs8F2ENgKAwfHBV+eiAMTNct1L3/l9v2UcTdBkvoGFpFNEE
K3hn+E0eUnoNIkADbK9wIykABA63opy1U2+DpMCempwzzWDiCxOD24Rr5y1Na1ZK
mNcp5rfQogF9qNHeElxfM1JSBgUMn7oMpUMXWysDdOE7mukzF4RRmpaoAiBu5Mwp
Y+F7l2g2tBgwnfPgCEziYKc6xNi8+c+KSHMfomqySNNakna4tN+TwpygZXqPXles
fwjEssbsRkQZuWQddRhiZE4mO+I/AM8D/D3nESyYNSYdy5BB298K+dGYpEjwJqrr
hKuRP6N+TJBzmhoswnweoaY9W/GD3stjtfPYWS7jH7P0twCKCkKeQ9C42i4OBVRg
m6yK7+nfQdoDCg1ubUl/iXe3u0qeGRo25m1FfgqIsRo8yw3RGyxo2h86SCi4N6dg
mLpf/718R2ddX+ajvTB8Okc9uh3Cnu/31gEw18x8SAec7kfQtUxwxOipvEb45VkL
5MzZ+/FjmCdvjTwXxrWdQFTfsMKnFarHhcflqHu5c7zP6bRuuU1LpsK5F8WcGyPT
bAyyiW7L5WnouHRSOfzBfF4b7dIgiIwbGX1j67s4U0acpNmIlk6WlDY9UO//io7T
/2dgl1M5rtzTo/KGvP+Or0vjkubYk7DEFUrBSzssgils8iNPi6zurhGC/w4SH7lB
+lHKGyZoPfy2HhfowAbPiudL/4nsJFGazCiCaK3PF+psbUUTXRjrdHbe9ikb2cND
AdipG87+JUruxfZKZBE2Tccb8M3DM16ZzXgHLkNG5kCo8Id5PX2ZVZW5fW41HT0T
4VL+QhM7rYWKsefOJ8D7wPuPuAdeY+0YGyBLhe9ZEAjPn6AI4kB+NxTkRCbjoRN0
+BJ4HK5VjQi5+gdor1Mg0zgUFscYpaPtJSaKT5PJ0t8GS5YdXNNkVz5TEXx0CJeT
jiLSftIvlsfTX96RgrtngmUUB7RJ9r49sPWCJRgwSW8VwjpkeBCLZCGkFgP2hjjX
Tg4PyrY3hZJRgM2V6jPvQ6Q6dbvwHo9i0PLRynz0tn6WGST0C6XjNrS/m9wVI3iY
7zc78eG5vJQmTShq76N/eMGXnwnsBPMtWss3SZCrwczNgnbzMrV2bk+D1MYD02AB
k7srh9ZPX/iwHfkmejrDDg69xz+x4OP3wasggADRL1W2lV0UP0yt4Qq1uFArjqLC
Q6grpvwOFjhdbPSe0/MqCOjnHmD1YIJyJzX7CHVDqpj7FJgi64xpgjgA1uLO6/aj
ISVyHpTo93+a2bTWL+RckODX2bSb0/ENnU3raK5dqMbv8kex4R0fLIirv76JhtDm
TMBl3d0A+ZtflsFzvG/69ORblsEfTlNGLM6pC8QCQvd55eXNFAK2uslPKqXUHK/6
lOc/Y//ujjbYXYb/m7ztv0ipCEQts5xVbjDXZi1vM0WO5FRz+Zf9NSd4iAm5OZqO
qYllH1Il3UKheBw1ztI9TrMhKMTZynKfUU2Nijr0VayUkT2+E25aEZuGeDNHAGyS
4P+udfILOx5ixsVva4JQWeshL2G8T6gj40SRLmX+UuTiyH4di8cFh2dxm6DZoRGo
PjO2mifX1pPhjhT3jprnHoVpEaT5qNaJjarjpJF2xNP1b92j9Qfr6uiZs/Ox/bu4
1Ea6ZnxcydlO8R85dFPQjDLkxf5b+SGg8iIEmHNuGNfczkMzwuZcjaza49ljHjv0
CBUCmnbVZcmfY2EI3s5MilL5tnhC08dacOMQ/0duoY77+Y5mlNw235BMs8uymKnu
O1vwqtcBhzsgzbqMIyw3T5frjVil6Z0HY2UeFmynjccDKTej+0yhFLwe0ZbMuMdq
nej33cLBGyJMVmzCviM8n6Kq6xpCozXr5zdAsmIgI76frX5UmgW3uPaOmbDI71bO
7nMHacJK1D+99dZtK9uBsiwGRvtw+DVIGOJUKMs4dh14dzjVvydHqw890Ll3UCMc
YOwi/1I6QnhCTNxPQWIF2Z37nGcmUANt8YlBzIs97FJ+ckER9TeSaZNY+7p4JCTr
PX0YZ3MajB73b6zCWt/ZN1DbRsC2ukKMtjCnaxPSOg8W2laFG5k2CmE/JGCrU+jk
27huQd0XpzRdxdSrhqtP6UdECxMJim7h5Sb2oO0v5trDtQILr8w2qksyx5azmGIm
VLBBZxR3CupWq3g0CZb3MksjmSvZBdzjMxatf/0FiN2H5wmhpC82NffYpJgc9vWv
0Hiw4Zt6HDZACKRuYTjja7/yZexdUBamN76jyU3anDbGpWkIV2eIj9ycM3XXbEDL
bJpK8cjqoypE4L97G7CQqu5asMtQJm11KfhyEuW9TqUV09AanUIbYg0P6gCHmYWo
7Dn/uFi6ordix8CHvX/JwbvnmsIDUZAGkSFRPC7NIXkHERtN36aImiWXszuPDXpV
0GLuclLbPQlglUHg6bGWP5TLutSyHfgdJImGrEoHBOkznBtWaQWERrUS1PEV4oW9
D/4nEb7Lg5RD41Vgr3HvEDIOPAFjHtCVAQxycy2plwUL/ao4PjAXLaqt3F7U1Ijg
yboWVeNLiC2JNEmKjcaLjsj108MpL/Auys/MkYKx8KSbxe3v42P94965uzwX9646
k4UzgD+lK/N9Co9a5ElPKVBkIq7DvRu+jL0RBMq2Iqt7Ovsg9TvQZmR0aMcntS6A
hseXBZ28YF1V/2ffs+3D4E+TQVf5jWYgTMEsXzjdhU7AoiTntRkmIG9H5+SlYfPT
LGPeRz+h00iSX3YaDsof0fFdyoTaOheXs4Q0QbUnA1bJls4mox4twpYlu3EB7YmJ
ht1sqOuL65Br2IcvtTFGaTFvXkD73V+KwxjmGW6B8rz7Ax8p4Q72w7hCiqsw28YT
SSJfMWegxL8MVD/G7xDemC4jD0IiZxYTvFOBU49pauBeS9lVAL8BiKAUOjYYlumL
dg6IKFvKP+dlvb4KzyHBCtFIo3YZOqSc+ZNbXEwip+CW2/+pVcNd3DRAnZUcrunG
D6uyVszMScMTfZhVAjcs+ul4Pr8ps/fUCrlgFqVCqNcubrGlnBIFf5TeWMksZqwb
xx+AqVGYYIA7DPTLT3pZpuiw8xJAoe3W2HlUllIP/39tP8X5zsM8+Yta1srlDw7j
keG/HIMHqxIDQOvIooaGDBpNJOHEXGLX4bbIxnpQhR8g7E+q0mc3w9G82aAaorPe
LayA3tDQHdxTa+jDNRuAr0U06bB+n34Z/mNbx4yb84Yw/1NSzMBX0bHJ+RwsRvKD
cneYlX4kUfcfr5DRIqhoSe5iz+cRBGqS0eVjgvyETSr17qiOddhT0phdT8GNqWdE
qiGNzZrDRuE2AEQaxUyNixD9G4Xs5EcI6jaG7NOykugj7yuozFji1m7a+kI958kn
7XLUf9SjFplTdymK0rBg2bWZqdKBwU6VUA2PQCtp9lmwzr6afnSsrmYNbJD7GaPw
Xr/ydwCKCI9CarlLewxw1fZgktvPP57l4BPTY0Vfkhtl18risNP2L8IbIb0/cXvN
AU0dDkh2uHgBc1LWiM77oKJkSATR/ICSNtHOrh1z+W54v/gTNeGc2x/VXZNX1U5F
9mTBSS3qSVnr/lW2Sjnys01Jbgwxsj4qjni5E4tn4K86yTbMHsqvhQg6tfs/u8KV
QmLmy+mfRlWaN0lfEgEBbAsHRFh36i8PiDjd0z/ucsanzvreUSGKEHs+DlKJY/LS
NHoC+dJAHfoYbTQR/YAIWT8kqqzKpU7eZRt+e9vVx/uSYIFuk8ygnrK/a6BPifW0
gQYCn6PPcH2bYY5mWwyq71fMWmP60pvPKWjA/it3IbkL6sA7vP01YpNn679e5Cg0
6Ac6cii2W9oMTmatp2VA3ZyxbpoVwLud85w/a7vmiz2vz/w91ZXIF9iLfsBxTp22
HJ/u+BnfKGK3iFw4vGkH0ZBdb8Wj2Bxdh+wlUBMk8PmtadB0YiKO3XkWG2gwa8EP
Ft4omZ8Ejjipi972Fl6K4JIfcgZRG8fcyET9gPR5VpfGYgTfXby+/7KQAZs4lkEW
1SnMrvllIVqmI+zxfG6Omr2WEr3QWM+UDN9dId7by7S3X4YlTTf2UWIC3a45DBxC
Y5H+w2fp6KJGNxTaSbgr0JI12UL37VO4Hax52nNF9GyKQGORDPssg0yIEe/Wj5Jh
Qn0qDZCCU0yedYoQVHEVeRrXtD8gZLpBnDn46DP/1wovymGePcHvgxii3UxubE9r
WQ5thxwvF+kno/nKb/kCxWJBItZfOznTUERMOW9ly/6kxgte4j5ZABKbcQfmtm96
jqRgOU343OHStdXVfmTRx35yWMoMWoYreorsk0s3TGusisebe4+ixf9YgL4PzYBE
sl3zaefqinnOmPEVQv6pt/DdMEr/mdry8esr8lBfvELonKxOkBLOhoxI7iNsD6oU
pCOzDAo0RMewoZzapeq0Toa5qoltXumx0dR41lqn19pIXzOnYZNOWdYQdup14zix
quPHXBsw5F+mXcndrqfjgtB+fy1Ebro+QDsLEgRse5pdMnX7MGsZLyzwQ1ZQ3klN
wQB/G2zBZe+8/dr32Ar+q48/3KRtyiGGtfLgXczlRYmZbaXUEKniF8Vbfk9Rlejr
e8kK2QcpeHyYW6eGSiWlKYd9GXDBiEajM0P5I4rW/IscGbp6/kn8XTp1W9oN84af
oCfE9Q+6bJ8VamAI9U3jftzTnRIG0XfiRo59gSC19smEbQVxN5SxbnkuQdplFxmr
YAcYQ25T65rAL5BIByCKBVe+oTXXH3OV6KoSkJL7VuTu7Dr4wiz6zVCuMS9gnqlc
soDNtMTqShtGOfEIyrIf0+BJi8kr8QPvt0NJ4nVoURHLIdxMkZdPZTzdx7LiYsgb
7Qrx0Z6WY13yRHJCtW7rg8NjOeePCZL/+HQ9/jD229AYnC5vryoqXbDfmftm+AsL
/rAa9949XvTzY9PhBujTbXtM06UIQNn9DuE06IGzTG7+MuaJ4YhbrUuDLiQKSQwM
zVQuF+o5KTn+6oTqyy5+pJXotGRM/YQOX5d8I9yaC/rKKrChAGLKhd89kETtVTcB
PfUdfE7P/FzLyYSgIHM1AqxwGNLugieolsqqwialNB9PbIxLI4T0C0/MywD+OixP
IUvSRY8mOJI8B0CRvfxh0sdd0ycsJ2H8r+00fZYoIt3niBDvsXz4i+FMSXTX6AKn
GarFe7gOitEVctg2Rd43J/IP4H/F9/ALPr/sTdjQHw3S6XfsI7zwhMx33qaUgTSt
4mJ4pPgFgIzIwx81rFeY5JwHZOvehSGqYCWe2PXes7u+w3hWHCxDS8EmF2shQSDi
mgRyBCynHIR9/gHUtmJTcm+ZBx9bsyK2Hw3h4xSeVbcMi9BJLNN0IQNH8GfJXku5
1LOvsuCApwfNe1/HspyeB3JdS9ti8zjXuYTVS7zoa46wdufio3Qvjxpx2gv+hOM3
tlws1hEhGYt8eep8h7f8YYob6EMIq1LbB7gnFnYSjrnKUk7YDwaziPXYzEeVV7cf
1HDTs/Nf8l0St07p3tE94t9PaB2MJWsYNec9+/USBUpoNOi9zKCvdN56pyR8IHIG
9q9xZ+IOppi900+P8aTmL5fx9qNjxXOnwyzDiX5lf6tA09LJqBYdZeYzONzKbtwb
aLU9dh3xfPxaQ5EC7VsYHM7HXWUnlbtw/KQ9YXWmdoCb5NkekQyokHGa7SZFmL5Z
CoYiHeivRdfbji2E5jB8jNANxQ2DcCzEv5/1wrWGKN1r600iZvVL9sX61aN33tQN
mSAOgLMZuuSq9Ufh0YtqcF0i6fZEWJz6184BdoAqI4zeVhUz7qqezfkdtvBHfALi
bHH0gnH9abNXYX5E2DnQ7mzLDww4eD1yrB0/bwnKvjbHUY/nVgRr+wGWFCQ4Apla
kr2N5vAdUQWaaqV13duaq0YMKabQWyv0d+6RAS95pBwYNskxe+vK56DaXJn5S4DB
F8SkvhyNq4XW+75pD+AqQa0WpbDnMY2nv7Z0hXpIz7D0vEeU5XC4aYoEXls3otaf
igGySDlbgPhK9KclI0wB9UeUFfLJmVlI5+fO19eBZ7IUP3aJMQRM/uqd4fns9TYK
6JV2sFfABNDBqt8hXeJZ/gkUDwref68ApOEDobNOpWII7zkBZH+tnBAw0CcoUiSB
4lj1MheyZmYA/uGXOS1lf9GBSadpbAHJDYwYQaTEdnY4kN5zaYwjDaDx0TLbBIci
ZqfUsQHyDcr3UHakplskHSiP453OIh4SHvtHKwZ4vnVoUrwRESG713Kp7xoyE60q
dHeGYpALavZMGhFmZjuWAnR98j0Otm90AOH0pMcVqiTXj714KQ26E0BF3rcCxes+
TLfp33emHTnlBNUyizB7sl/NcBwcg6EQXXN3Akb2DMHdIbZfTUoGEYJj3Pnxi8qu
JsErypa3Q+jPjtT1X7t8YK21Ap2TzPg4W9JvoR/yaklWBL0xMOyQ78A+y/SDuvns
27digZaCw8jU1sWcTUAx3/CLOuYT6vTknZTweg7DAVPoaIPZz5X0n1EieOWF1i37
G2Q8j1t3vGuAHqeJpKYpWOZX2kOIBwxPRLEH02O+RPwrjE7lLxPZ0f7vWwOHpe+a
ies0yaBSmegwdl3JkeXh9RWn7d5nzU4w4UsmR1Nt73Sf3dBwy4+oQiC8+/vPxK89
xF0nUNrsMrcWiYeyfkY+KNzBgNQUQ69wB7ZJXkqT8eqIAQJLxEC5XYnA5UYNOlzM
Hx5nZIAH1lXuVdemOKjDH9lLjFD71ekwgIdGW2dwu+hecZQFGdKtcSC1fVf2Iw+h
J7IWp+sOT+1RVyyw9NS//NpRoPWPl+MYhB2m2hkBLjYLtlqCeSaQHdesoj8viDfh
tJVPm178bI0SqxbjJbp+fG9+SAvue5gxjh3Gi81vzISsSaiidqdnqs9ROr315RNF
cHXounD8lp/AchoPlJT/wDolmR1wp6vnmvux5Mr89+Yz2wT2ulPdDGAl+JP4hBTC
Fo+eJaXFGsRp0gYEaNScOiycgELWEsfDJgDZiLazmYeFKDiktyMpge4miZ0gilXI
wf6nRyX+qeKqlNnRuvmxPWCZ2q0ypuhBzHXfcPEvwDAfmkDByPrje1Az5aLYaPTB
0SZmAiUksGC4HHj7zuwtKVLyByl4XtLHWkHdQWMzA5a7N0eIPBjdr12HsTaFPmFi
4VG3dPSSC5YFR9QGvIc7aP+GzBIbtMwoOc5e65xzUe9YhuB+KCXsDfkzXEkFWNol
TD+tZZFbIdCQ/Em4nzIQ/sYaMg6Aqs+dWpkir+75zMoQ2GHSq8B7+swi3fQ7fhz1
p/oVRJk6EHUfzxfWwYf2HwSBLVZiIYa6s9QLPgVyV3YDAeiXEuBwpLHslod82apx
zr/hkLiAhLEjzB/duATO2gkIjI61H6jkP5uRAmjcibL7stb7yOpyOReHVTw8j/uF
kvkrAxOFx9Qw7NA0IpSPB9KXCX7Y/UhT5eGXJpXsjuq+KMnRGoZPKtGshH1pCN2R
Aw8w9iBcJCLeSgtza8C/DRpJ8z6C/mkTvkgCKTiRdOMUe6vXzs9lEFit4AIiKGr8
FzzLmI/R9umdfQF0NRZ2gdhtVxMPVKh1BdhC1RK5LaWJDDOBu+GlSUhPvp2mXQLU
ODGve0PyI7feIXSh00g/iZvO8vUPZy13Dxxlo7VClIlDgDXBzHgqeboGzz9Iue3b
4QMkLV/3T40FyO4GypsqGP/rRoyh5ndH5Qz26+MBPDWuCGFB4203LTCwQyS2MTiQ
S+N1ApBx01InOiZ0lWfVw7ILLAnIayelc2fj+CG6LrkuK1F9OQuWpk5FDwVAZVmB
cKZ4gMgRn+Nbg5519pFPX77B/icOKFmu6Ehb2EX/DAKIXHG9z1/EPtQ2mmMtwcp8
IeNEnqnTjjpU5yN13gdUYA4bOlH4ub7xSBhBOTvp2fDCrD4vY7kvezioWuT+rieZ
herppNn+yBSwrvPLScu/fvNbktNiFGHbsPSViLj539pYG+RbWYptU2KMdTTxOB38
UkAb6LSg/vERRri073LpwCkiey7Jmaf8lvk9xBjZerHJ1xgMbRQsH6mKCqDRJASd
TqgpLCmwg+trKv7d1oFeMBZdS+rzi9/74pF6meQCgXHa3WEsK7B1sd8j57sp4S+q
wETPFKLACf7jdm2npC9rK49xG8cb+cbnS7CTmHlCL7Ft05spoOq5v7IBMehKFMyj
8i6qyKO4hkqX3zD2MdAYC7lHQAEn0vACPDHT+/m1LG2SL+jtXiCmkDhWQu+6CYim
ccWiBwZamYEbkHMRVi2ykHFDM7GNaVIU2P8Kwx02u7TkeFHZHiMJID6fysVGhDnD
QgFws9EYgjZJwiNT4edukfL8Sr7CwARCHfxZ2uItQ2upFLvgGQ64i7UIq5OcT40h
8G3mcJcoNz/lVVF003Ioc64WtHEggIx7QSUdADBtsn1WXAe4gS8n63lZrIwBu0he
/mDserlfX0M7RChSAAxcqnGWnsD3x90tyKm2qdKV6VSq4WZ3NLrbnTXGNfKdKXWO
XLjBRituis6bLLLgGlzaDRY4ZOUbjM+SvKdToYhoezGtokzVBcUCwUmsB1hLXtPh
RlJfubCI2o9ks/o4vN+Y+xCPtqZkaSFcuOR1EHV0Idq5iW0NuxmfyPTctV+Oxyr5
gAaZfOIbFCbOeCGbMyD4YExaV59D0OHHOrWVe0UqPklZ8GTMZzJGI5Uxbs606Xd0
cBOm97euGcMLw+5Y6FMIvM4lzMjX+EBv/4syYc2SUzSy9v8StB2ECb41rJacGsbq
trGVog14NhX2XErE/AoLxCv0lN60e06agQie+NBtZrA+hCjcsogncJYB+VAQ8OWr
mHRLWvoSlYI8GvPsDDUCum8+qRVv/mpDWg1Cy3fkQRpwOO6w1/b/bZrcBLlNCLGT
oF0Q4wGZ6aZCYS3gye8dpyCIv6oWtO2+W7RvJBU/SnVD8Zjc81gllH/vmjIJF+Sq
wrMKyCYrqsy/L4B/koD/GPWiScAKSrdkSf09KDdJv5HByrpYZVcL3WZI6w7rGwBf
Eo2G7O4ichgROdOToEncDux9Sx9aFKioP4UiUoRz9GdCA4Y4z3IOy/D1dyygNfmQ
RdiuBbZcaQnm5GpIdOcOl0qTe8Cl1OYHfy/0+pQS+ZU3zf7bUTmuiI7eWl3K0eCX
m/PjJWa5bBY25mAWvVgHoNeNK6HUrRLq3nu6Z+hohl1th5fwGB7+otph5T3ns1Nu
Fdz/t99+nn8XzcqYu2KogKNg0WTnF7nRtivcQScj7tgtCH1hUfUqmP6tLjS8O7ff
thOxXRK1IZZfwwUOl2INvR+FMvDBiS2YH8axGKBQ1vZoL2E3EUdrYUiGaXmVlI0T
9B7dcyvIQqp7sQwct0YY9Ki+qZks2ilAgmnitZBnyUcAy/pry2buGg1JwD84vWVn
unNMlE4pk4HfXVtc/fjp17cpYxbTEkjwwHpuQpaao3LsDcyG5AEXGfb7Vd5NJvcd
KvoCYN928waNQqGwTNUkBu/ZOrsDqfW8mKSQSFG2XLANz+p51dx4rRdzNIjKH0ct
VGAhr7oDib7xQv6zLSISFm9/eoNhqweAU4V02EJwswrYhyMxkSJ5bgfp0jY4wD3e
9N7+hPJNvHnHITVof9KhIUIZj+wm9beZ0HHslaeu4DzPanX6+HAjqQCzeDIIdS0n
mUAaXa3eLm88IOzBJTXB9DChIim+rS7vu82qtCW6qjM4HAaJ0QkajWExWXHcsNJ4
CL/UvqfnLTccMTnnh6LfzKbSQwrW6NZETr17UX4zqd/VXAC1eQcmxwOZiVhdHadV
YoNIw89AZuGk3qT3nl+23mcsohWXCDZ6Y5OJ0kPxtjwtztsUC0DChslK9PSTVFI1
uGeQi+AJK8P8UpvVcjlo3gW3azE/TpqH8ie4TKJD4MIk43+Wo9jzoqGeMU3xHAUn
fSDayIaz3FpTRVBHKFh1jzE0ExjMmFfkiu9Qi1q1G0RXAoVX1y+HI3PvlZsHFqgi
TFrPJK0NUmVP2ZD+FZXgeACg6RYZK+QRX8naZmbmdHn0yDS8uMdHJOiH21bBm2BW
Y10Vrx8WMrS6b3/5VBP+zPLWIWlK1qZqWFxqBiwzzqP+rtg4ZMCkr40msikhGLow
90zjpQqKVxpO6mSq1XM0yaGugH2LxAcLxTKj534wdu96xLHWUqaO2vOu+uhLUSTT
dKjeoH6SMsnqieHH396WqspzpHQwjYJnTkHAqtUwvNBpOeZ4sRoQzrL8LSe3Vcv/
sQ+IevTAmQjBWi46ZwqglF9nQ2Nii64vc2gsfuAG6scYFM8+x0eqphi1xG2jN0yr
nHCaQm/2U8yCSb2XLVbZSP/Yn/RGiYfI+hs/wFfa/jcanDbYle6Zk2L77T8xpuMS
IURrCF0QlqjaVZrs3YBlIglPaAVR/i+qcOmo/Y9mGdLZRHc/D+cTHmEY0dPKV+d9
hDQnfTQT5pzRMvULCVrZMWi7BRLpjxGem3z2uwOG5ZoZzapal4KY+wz8h/JCu/HS
OUwHcAJHlKhDd52Is5Od9MPYyXcm2UbpkzsNoSzmN0MBtIqE/3fnnjAw12i2KKtA
skKvW1e98ybVqINwLyWfKY98f6AF0elpOds0ulpSaiViM/kJgmtMbxDbyY+IDa7Q
wKtVioMhKX+nXA1U2UK8A0z9mlYDgti8YCc4Oy48VfkvEc5LUm9xg9zZvzyRjpRi
8G+B2nSqPN1FW+SFPEovE7JVDa16tlRN7871zl+E4Ud90YWQ/pA2mFaQhWfTqEG3
ITBiu7KFqW9QX6yKwOoMdwayTABPbCffjV8hSmZ0Afby0SqT5aE7QQ8S7RYLg5OJ
+7zYT/4MGJANC+jg8ARt8gyglUYf2sRIrcegCW8EBjjlS7lyP84h4SgZtkj9W2Os
PHLr64k0jn5vt4geMdOFa3YjtE4LU/Y24et2xoe2PkJVAUoAa4g3lC9sR3I5UPom
50/2HSCyUvySN2jH7dfdqk6BjKMAqt4rt8iEJAaNSpE9egLH7VKfZ/ifmUO6vzvj
Gf7oCk0rPwIR4uPP+3rYRB1pUMI3oJmcqfhUFPQufv+TWj9Oe6Uq7xpVRe07nAd+
v1mP+q7xYQ6CL7nm9heW/GUICTVtM4T/kzQJ/msJQ7vKu04z2Fo3C7ofcfDHPTrF
r3phCjxSuy4zYnYtV4EWlYpsuvIKb5HU6Iw1lddpNs1dYnijg95RaCjdMkeEW9ge
wN484vb/UelsgO0gQFYHpUpFXI4//7ySfVtkXJhUX8pRfEjlm1E9eI5XVpoZdXuL
MYqh1aD8HE/j4xZD5EW9MtB8AXX4ql7DY23xjGy1LzVVva3+MvP/LMAJQnmRoox2
mJirFN5Mf30h4PFZ3F3mwdA1TsWf0cI2MS5NcR16/4fOMuEyLNCvzq5dfRcuUqp+
ugFk54qewrqVsyXZNhw6O4rD4NwEznqHqV9xWNrMqRGzRsU6x91Iwf07ywDgY5ZB
1LHD5yQUEXe0RHZq2VqD5NPTgIrHVrQ/QG9ncjX639MhIXHCMktCl+zl3Vafg7xL
cd37ofj4fC46NaP1HrjRmDHoC5Zl3C6BWYnmj6ufDTz0Ey+zPFQsTpWg1b4dLx+R
5xxtOCohsFet89P+ge0+tXDxmXr9bB5HzMcKoml55IRxY863+KcJBPF29da6Jn6z
u2HBjSauVoeM3TmgCOzM0wYhjzg/HhAO1x+WSha1QYi932ZQtBe+NKLfY8aQPSM/
E+LgQUsNzGwAEXqlcCAL1Sgf+EzTj/BPf/ctXyB9q1BZDJy6afbj/+0ng13koAae
0FsNx8DSAVvcaTJPATZelccMZ2k0pjvM2mBY8lkDcsr+OB2s7qeZW98uwnvnoetP
rcm+LdE2He+sSylM85N9X64v7T+XPsj9XDVlp+wB37eM8XaHQiosD+RMwjE2Fp5L
XuiJQDDLaRaPuAF7VTKKxjbPIYiaLibvmJh/ofRvPDqPAZxkH0rTAkH2cFDsUUJ8
zRuvpkPlEB3SdjMRb3hiRLhinCQnHuMCLziT6Heq0yg5dUoUlrmIElkPUDmPd/x1
ehYC1Ooi9r8BTxUQ+lyw28Bwl66S5MV7MHOIDAeTpXbzciBsXhRzpLiWIUSp2SYm
kKHjaZpmizklZJPWlYTFzMjp2tz+EOLjEpYNlhVHpv994qMJFuqfXCkhpqQH9AVR
n+Pf0UNNqND7dT4+TLkAIVwiQP2exgn1opBCUHPujW8IUycTaKlFIdonJ4MHpZ3j
KMh3+YdSHBDdk89Uj+Lm4h0YDFGtxF5Ut0/GjUe5qh2RsqKEpgYu/Ply/OcZZWkh
YvjfXXouT/Qr7d1EQ5MSX0BtpTFKc3u5iCMaeRT0aueUzlDiwcX9oxdhor86SF1B
nIr9re/9MslCI722G6iMAQ5Yi2MxLqX8QHcMKstEpFMY1iOlWGls+vkgRxBDNjs9
GrK7hFcjHMF9ZQxdxTh0MhAXfws6nZLahVk1dUuZ4YbEkHyDfmoJH/+lQ/Q8wnlV
uCWjt+VYvZ7H/XpK10oKNnnRXAibGKhhebHdslfK+4MJKTkRjOzzdr/XcKF54Znt
W7Pz8qgW3OIzM35sqFTUlqiZhAlzhYVFhmZrCUFP0H33+OT3dHt5jRRGSs2Ak51x
6JBLCUsKa4Zd/elP+L1r0MSHqMRHI/Id3TFRFoKqy41xHgljOUq8UStAJgroQyL+
qKyJ0rav6+Mh7S7gu6YchaaGb9IYpaNUsvG3sZWgWBu63KUNMr39PQqP8KPGhS9i
63LfYMACtFTHUOBCLgSDi+RUjTfaZCcKecwwDC9g4yPi45+2wmrmjzpAccq8p9qm
0OuQXNM31nP8UQfSBf75VOKNLcXQgoL3MOyA+HAVGjqf1Q2Bws2Zb2plp9VIRODh
b3ejMgJIfSVJrij05l6cBiYcD7nBpkdiL7eOgx3aRiufNAFOBldN98jZiQ7Vy2TQ
he2SgC9ZXuEYn/qozxvhs6J7uWmMULVmtrbe0ad0dS1VY9nJMNZFHTB69kIGjyUI
D+4bTsGSNqtE+pMewMkVm2z7o26L/3QMv63VVZvYoAnVaoqqksAzf0BPG4jr6UnU
dGZs/nPrjook1RUbRgbOy7vsVaGTn1e9HuiNDLpX0P9lejSWpM7HzO0e+dBgzU7O
wQZcqh4Gyjxywv2ywl5I1O8OYop6SjOtxd+3yp0ojPy8jEvT2KfwQdSS1YHkELL5
RdUIigQNa1rSgVRKcgDWNazoAcZ8hW3IbZUmMpyuLkhBSsd/bzraqNQ1ZtnGtWUr
Uiv1llzACCcH77SuE1xEzvPHfjF+hFFp86UZ9dWA8dlCpLA2KqHPIJrD/j9+t0l3
zMtZDZENwPtgHD0qD2hdok8e5C1EvuxAkgrPQ/RhyquDvUo/yIeck+KH4fvtqkxu
w7brsnYOuugAtJAU4bcr/ToZTkEDCmWalbeEZJc9fxP2388RpIY+nhZczqyLQY4P
9xn53A4+VhrRO4rQM7QsvY2XixfCn/cEeJ35JATRl79SQCXYbd5r7wgHsWrOCPeM
xK47zhsNEVEHdF0TjBebmp4q9QAq8cVLV+afeAD2U915p51stq5f/asOvdYCm76i
bkfkylL7r3U1RnoAtcfGmsm3Bpi1k2Krbganvq+lo77QlJOOgtyiPeDg7q1kw6YX
NL2eLsA7+g4VQAyij98LojMFvVF3SNR9wOecYBKnKwF/QkbdEFgBn+KVZ7Xap+nQ
hiN/Q0bvWsE531DB/hppZuDciqCC/tQke7DCIW0LcC0ORvRKk8U6PD96NrkXQbO/
AVtM0n+RrrC3+yr84OdDDpjx0rsiilDO7fxAWG5DexqCCQdHX+aMTdbkzc1Zk5II
r6I8QUZtjrJs/jzoS9/WioBB9kTyDURPo8Ai/dlbIa1AdBwoEbdiJReLjpAFqBMf
7vuWy8dIyfSHBRH090Lq+7fO97Kqr8u8HkJKtOT6IuoKPYJa3aD2bqEWoS10LFPH
LhP0wOA5oL27aT6L30+ydlZwmUNmJAnc1W0xdo0lTjFziDPokkuK17xVYF5iFHc3
3YWftXZy2ORqTZKZq/S3j/uz3Ivv1sN5q1R44t5Q58qesr1Y16y3kbVuz9JXoYF4
ZIuj6FFef54JnKCeOJOnURC0it+iPyTuDYNZLeJjDu2MsAl7APGvzN5xxYtcMj/B
3tFHKnEXEuXleW+NQVmp9dYCA8PObmxG5AcrtlKqSN9kCfxWFD/N0F6OwAffvqRC
7HVHvo0sEIaX6JSyNyoJvJfCXTHLOePHATKwoT/rOy5R7odqnKGdZaObOyENW+s5
QvWXGy6Uuvl0WcNs9MgQtTRjU3TDVrDMN+NHuYJDWwU1WESwe+gvpaAlBCinZgOk
IKas3piLjtvM2EXki6wM8ZwuXR3i//cpW+SB56pM+FcC5mrjTp3UUCQfLxIBOkGd
55fHDcylYovBSBpxWDKWhIK93ZG2PZR1i5LbupeiXw7PiP2+zam3jHm/06i+fto7
i2Ll9TqLrJ1FYcV6k/DCm1HOt7XtbTTOt4gijovD6D2xe6n3AlFq/FAQnWwX6EFF
N1VejN9fJYFMHrIiXwRMsUw8RsGUBNqwMHaFYCluQyswUnI4dIpvm69gmnm35j/N
AIOF7/IpNXJmZrJxcQTXc6Emol//iTy08x6rPp5Vmj38u7h4frIWyC5wELgGfhGg
bqXt8vIsItesC54E4se+7OiIeieJ2D0fvURseqNYBcL3zeJDHHH9C484pP5x1YFh
smsZPRZBDJrnK8yeNzTFx4+1qOGDk7oCvyoOfJU8jwkxKm+FmXRtBgJBWROHF+aV
AYiCMU0ER/cyXmfRFeulM+GmNOz9jz1llD3UotOoxvuWjlNNDhs7dG09bpD/ZuMY
fRkizXrbnLsBXT3a2ABb4ny4DPwYtgG8Qo5fb9NugjwJLaO/3o6A6cLJoNBuOnud
nerGwlQQmU3uXDvRx8cxmwMbJje9OHS2v4jMRq4ZfVZWanCK3+DTwIHw0tAqs4Nk
aViI0Q3ppDLm3F3FM/TGXva0tYBTeWz2bCGob/6C53DRI3oLqnUauIhPJI0pmno1
ACcAFAYWpngxvSV0WfFZCHyVPiFIIPQznOiw7xBA3Za96np0pPe2nmmHoP54Fhzh
4MMeVV7Xbb4GmScas79ERAuc08Sl+AkVUWWdvyTE3NPT0vcdFKcrmTfe3Z3eya8n
1PXRxq7Y6ZK2aEGHlJSjBDqZhh7Q8TS4KO0TzTVmhUuBHK7Dkz0wcr5G0mvfz9Z9
u1Tq+Fa+juVdaQsvUnHUdtw1Qj3B4UTl53InhVaJj5lhxqJY36cbqxqPrPZQUU2p
o9HAZDZDPABhUcZgNvQrqRyADbuJ0dq0MxS/n1VOlfYmBZ71Eo/vxesDz57hCXkA
gWW9EYFTHytzKXMZmXOv3sh1oNLIE3lPVnl8tNcVAJpJg7wUU9jTjqgCl3jbuIiB
NITZMlrYEtM3cijWAvEWLHPotJEVR9FDqYZ2ANZEiiNjYSIrYFKfkRcYoThQBMlG
1O4PDVTYWypt4RyzJ7eGyw9RIfcAyhP2YJ7/1ktGDfmk20KXRgqQXWGnYoi4H1XZ
UDUvtluZVFgBXpaFDk3m6XtkSEJNVPpFBJSTwcZxWq5V21fMhHh+EZZuSPAtaNuN
lAinf4X8qdyQkY1XY0bYJdFaQxgRsdXJ04qpC6iZ7Ju43RdYIuvecPXfsVQijbPt
QmYyH/kzznTGtWBBMVVHGfJdJWDNCNjtF87IU+WEhAuvnjR4dK2fKOxg8livP72C
C6m/0Oe+rgyHc4w5zh/72mmboxDEk+du7gOHbHQSjukn5Zr406Cn1RddTTO0liD9
PRg33WgqqZ8viTpxNFWGuBEMSHPN/OQFOxeSpZB1dg2wBcGyunCtPucGP6UJ+Z0H
25KpKOaiVzSe5PRZXWTkUyweqeUIm7GZbBrVDQkuJ4eYt5bAyhmMAmim05g9pQ4Y
Z6O0KlSiJ6rQMKI3QMZuwR1jU723mPubYLDQPZmyiGGouepyPqeHYWz9WKaxA2pF
NJm6Ex1dpMpuXv4hi+biZDQZeTNV9ocvQAAgzeABgLMEJ9binmAhK9IYgMi2D6Wr
0cdIqJ9p7LxYa88JSDYRWLM19DFd7TmvBCCIPOV1Of4r0/FrTsxdab/oAJQqrEju
6aCtuvRDFRARFwmHxbqjpK/o/n3B9vMpjgWF+DvXYSGCQxC7Ng47s3trVWIvmIT0
xNIIUkA7D71nNtCMHGkH4Wgbt8SicPvnL9Obnz2CP3D317y4bcZtefp4s2QI8RJP
QFWshFttVh8B2IzUeBEbaX60308Zt9LoKDgTuOtpWq/6Hm2sFVO+ak2gzPt8voUO
w3YjaRYQGi86t2aApzhcU/5AAstFS16gWM7ymWn5AT2A5+DJixVEW922UtQlMSrr
vtOe/+ke2CQ8faiOSKJb7W6lChidS9sIXcmcgxX1OVTtr5ah69zLZHJ3puypS7vK
Nl00CLJyrfID97Cyrnt7aPSj2k1vvd5HZRYtGrUB3ZUcMQdG4guAw+fQZg/iKrXj
+vXoVcumOhBt5W9xd/NpLwHP/dmNFD5GaAQJSMdhW9ikkpG4UHGCrF8/rRHrKVHO
2w8lFsBVlgfvmWkRToTT1oe7ckbUdqCp0qGkICi/dDWOFy8QgAHFc6/wpJQ5FLsE
WLnU3nQGO0thBu6u1rWs8eEEkSmG2Uv/hkNbLZELGfLnY4aOSiFuy1XrjSTuGcgX
n82Ou/yHPxpT6vEyZhPyOAFKTDxsiPdkW+JLCV6uOqEVECI+mejmIjqO59xM7xxC
dqnc3hLtdf1pWVZhUbxQ0MEJW6Uhaw328c7qh7d3GiHdLiVK+QpgTlN5eK5OLmgZ
inJ505Muhh94WuYEtkAfQ62UZTvrDNGTEyfUEkj0KBtiwGHomGrFvWSPILP8xWG5
e7V6cb1LNukyppSXUcrKgTBIe5uPZ3wXmUgp33hbxi98+Nwby/SFVINO0ATuOySP
/+wweXvmCNiZh3Xb67SPBBqz2j0cf0L2TdJUnRcnZCyNT60y8wrxbWExLe5YHAvt
PpNG6W2UZAZ02R2lyGfFcLFBjMw7WeSFZb7IsfV/7C/khNEYmbo3+X410pHgSS4N
Izx3wZpjil3JcuxElSpwaVma8/tbb9o8lrh8mdQQl3FylqQAtqy8MlVR3/fJFVCO
y3dF0lW1O26BXIzE79Jnxm9D/6dyZfNHjV4eFF+zQPR9cGrAhZHFpr+t2NNcnclA
THpr/FMsg2MFKhIc6uK4cwhnwtyDM3RVg6wbSB3kknGMKe4uWWmNCi/DmsmprKzY
k/D+NIiKq1O5oMf0awbW08A2IrNsiOkMNozGlv1tcckZV03EJ5dq248j36XnSpxu
rsQHn28efYIN/VTt04ZenIHblwjJXBoYgizWD/KTdI+/1Ovsu0/BeJBMR1BDEmnT
enjnq+Zrzt7nOayNJAjePrM2zGybW0nJL/vTVDUa94ttQuaf1aOBGE9adhoznVe9
T8chkZezxphDC5Wk/JGZsJ03Dck2wP+P5gSIdIYnlUjpCOYYRN9mJ3ba85SqdpRf
XSE5QjzU2kKBcAKGaSrIhzgLGVKqsyqzGLqKgC1sKi0TcgEwyjiDeVbrzItSNKyG
KAtnbpZrw6bBPeolfjfT3ufE7EfJawUtd7StcDTxQaCRv6D2SL1b1o6OgQYR+YAB
IGXPRioyhI0BzkJKRpmPDynGeyUvLEykIXihoYL9zDCHYTpN+dupMghsLhIc6D/t
Mp3+NJVvkc+FOu3hrhOWND1X3JEO9tqne7Cx00o1qVg7ADVZNr3MYkpkp3QkzG3Z
dUChQNBSNW00i5MBCwN0dgeYH+O28oFtQbDFWB3KvdPqDiaC2PJu+ymuKb/CCtFO
BzWjCj1szedojRByRZzQJwg/7CUU5Ip8qy+U0hTEQLRr+xbsaoCvAxDHxoJq2sGO
BlcJGFLrhC1JxQiMdZPzxlBecAqno75q4ildngDRdQ2JRPlLl0mjQmomQRPKB606
4vr5kh9Z0++Araw7QAXNyNGU08fNhiSzi/1xMvxaWUDuz7VS5Ro/z0NlRJA7LpR1
Pn/EuTHq3Lb6iEijAhdoJmLpRnoOhvs2ZCfnkZ93cWdEsnQT0OY3yySn3xNrCsH/
WO9mI47owvZ2lia8ZZ1iih4ck80Yr4KFfY1tfoDmhBy1KJfAZD0uSJVyaADD0b1L
YCVpUuvUzGkUOy6wuitT8QuSuxEWnbdQY0skaMpUxGa7opoff/NM/hmpIWyPdQq5
QQqgrl6uGoRD3QWdQoKak1L1SrwpdzIyUj4sHMxZT61aEe+3or0/OHclinP25nw/
Od5fT+tbhFlUk0VyF8Cvp90HpMPozXhYb+o6oJde8W6WC55o73mWpniu6geeswsI
IftbHo+ASSKKrLsuZ6z5PClOe7v1IMrVYneGCQov8f1RVfdOtwnCJtm1aMhglrNr
iZVb0qmqp7cHFr25/UzhlDO/tfrISu7CvyVPWzWtCRg/0co6aWEmZEo0VU7djpOM
OCsuRNDpy1cJAqDEA0xBPCI8Y+/cnJSAGtjlFRWYcN5Ds7z016QFirjBmPKv42yv
6eomyqyv2bqL2QQQZBXI48wRH5frST93vx+9N7c4tDW2eS5Ltt+8R2sTuCtW1yCM
2+f7ChANzT9qrTMOUEGw85AeZgUe06O+F5wO9iOqRW+JwVi/tE42MXNwblvmjQHT
iseu8DyqEF4tZ2uknn+GajWKQP7P5su8CS7VEPSW4AoN8kl/ug9Ux7Qw/fip0ZHP
/GXE/yANIYSzxDUpozIbhsbi6zg4rEqiboSJ5fmxRIdZH6+OBkbpvFFLmSweSAyv
w39O6zM+vYeGWVYn5ir9DamcobDzRd2da7VCk6nTxWMCYj6qsUce8ZCsVrd7XNfA
VSwUGRrmx+7Zo9ad+gwN6mmkcaBEpJ17tbwhSe8W5hveiKAvnqHFBFGLSJDsSCvp
eQovlqvQqrOoY/A+/qlIZdyC1b84qPQuvWa8CY5S7lZJkneNSkpV1ckbS65Awii5
soidslJeM2akRUuAZI5wVFjZEL++aOsSPqXWhM7saC+O+JxlVyTkky5UWdNkJQPF
/Epq6XDoDPTB2lWTm4AdQOQfbPRgx6TTj0IhgfHe6joBQeF3CAxPJQOAl0n2LY0G
2QnV56rR/gtv3h/sACiR305iVOaHITdxZxBhRpPYLpGMHO+iO1g9TgQYjoNPhewU
vSWPXmhwI/vYlsqpqpqFp56FsZ2/9mm13FiTTh8VCE/GFDD6XyZIsui02nM1yAB/
57EvegmCKax7O6j6fZ+RQpQCSrspF9TyS1zR1emEz7MH7HoJfy0s7aCfdlvNJxjR
jLdYTi6TUfFJydPyK6ICBEtk/FtSPnkxUb+dSUvOukosn3f0RcWuqGF3PdjkdGTW
AUj2wzUpdW7rFRoLtBtB8mQ/WdrCE5zcXVqehQyZRiGPXPirsBtnDOFcHRJIei+e
LcoF/9gt0YdB8jWpews8QDHwynbsBKjPku5ijaYtuBqdClvmbuhfMK4BL0Xx+oGW
Kcih8rb4lehZF6o14vzzosPyS7cm4+Ch9ndLHv+ohDRBttx+VdEIQM+mgoYZF7KA
LLwI1jpJSRKevaV0zQ0uAnOOHu5EFii4kYtXFPPm4lq2coqQ58qVXwKWDrDutXVt
a4/AdBGhICDXw3DAXLIVvtofmrR50g1TE39phQp/kVzuBaO3EXxPEAesiKYui2yR
dgG9W8JzODPDUMLoFt5W5Qgu0GuCJf05pd2RiBDq7G66YsnRllbnXqEzqO+/0KI4
GngcJMVfTQ66wh0uolPogsnDGFuu1L1EomUzlK2yuG1NZZySCPcLZ/TYzBewoKRW
KkxWlNwfRj8MdA8rBZBk1HYa/5i2W22p7VgHjhMcRdjH5BmghpUYWfngrmkHzQ38
kI0nVSxKddQkQxRs7BHVg2PjBYOxAX/klXc0YwDkyWUBeH9Ig8KIF2LS60luHKKQ
lBs0Lw4L03MK1pVT5BQp7J12VKrFnyLI5jmz5h2eGpntzrro8BrUfYfVCILZ3rD4
X7brufllQaZiRQ37IFVUnG3JDnUC2HWFvu1bBpYzhzp2KVAYkIF2Ls0q1hdDyWtu
d0Yg/DuU4jlmSxQxujDs4a1p/8AEhuWUUCAwKlnQeTOXEvMx87rKPis9Uvu3SMbt
avz2diVTdppKGCdH1apqJmYt36Eg09WfFxeZKKQa0LmehEj0k2wolNI9uBo4HI0U
kSExlAMry0W3AhTV+3y9+OFsC2UsLpd4D8xVEu3a/Q2XgK2q854XCng5JRSOg1U6
SIDLVhlkyVwXDcUe/cwI4OQqyUJfNCsfBezpd0z+KOToY86uatA4xHwPbaL+i9Ou
fv2e8VTpW9edChiVhp36hPuxB+V6hygG8kz9AuoZyW5GAyybj0QCZfxXxTBsEony
GrEew0ggrc6dmh/LE9LvMJMB91xAc3i7ao591nMtxDykByd8+Yc/A8HPqIf0v0Mw
eCsi0+F4TSDTftU+ry9nSzcfyC0v4fYVwUsIUJMDB9fpQFlm9NI01+CoBzalRAqk
WV60A7FMvQk301BkfXpwtD9W3+0qD5n3CBC4Vvams1mlCDvnuRryPqra3vDT5FXr
CRd8OXFmD1cKVXe6HO/c/p4xcNtzfGcYTxu941OAZ6DDCyqXFqvxVxMsbn5NboMY
xjHmratqF9ueIJQG1LLYXqY/j/NuhSx3s0DwNxx3Y3uFMHjiD8qPwMD6hqL4fV25
5HmAZW5BFBq55eOC3KulAXbI3q+qTp3uGG/I6pIMDED5OclkDWk5/QdDtznAI44p
gd/roDFJL0quUNpHCN3FHiUPIxSjlkmiEaI1agsY7whtGv/P1WT8UPkxt/aOYqDJ
E/B2Q6k5LhxLnVTpXW3hK4BiX0urZdzx08cs/pOWB/4z802FQfSp6Yb2HgFhXNbv
hjCyrSc3rk0SqVfKJ5F5tOGrp37T28tnGTQvlHNEK6aqdhG8J4U68PPpageTcZP/
W/xU0SpuLaTAx4LfslGdyoGLli6j8TQVOGmyLG/jGUe0XeNaCra4eO5giQjdGTUG
IPv1eM+AkkrgGgdWnlgs+bv3lqbq76AcbcDNjNEavN2pT3or4O1cjL9xK0CEm1wJ
AL9CJHT4zK7iElxSHW2nBSAiBzud3E/wh7U2o6zi7IZ6kRyEQ3/RjuFFqfzNf9+C
RZ67UPNSJfjuibksXFa3YhAkHZ7Wbm4QQX+DBSIZnWhhjbEZQFSFQaHCE+mw3wMb
CHz6XbTdJZiRFGBVqQZc80yBB+vtPI4Eo/Tyrn5iCXC0lPaE+co1OnjBrvg3zVWE
I6WEmBFR1BUZ4gAQcgXS2LTjdkgdQEONXboHfTT5UiqFO1c0xsfuakj/m6PwkOMe
sh1LxPrJ9XWb7MxgTLpzSR0M6Tn/P6xfCOjNqYl5aJ9qQR2ekURzokXUT/fjNSzb
50xtSTI1d5rMjF9keXl7UXGVwaPzetqJpJ86opm68zcbLMiNlBKCvgmXmljGeU+N
9Z6c365V0Lh5RfECho0OTz6gnnqnsksP2YrDp1s/xsqUXDXw6qFRIFvxI10ixeGu
MbUteTfSgiCGaBYee/c/Qhbq72GOU8WvejLJb85Y167RFvMgQdHus/7GaAy4ooWA
V3ckqUPE0bHfj1veprY/nur4cOUjjRczzmqQS0v/pnbxHR8uVqmS3IhGFZlWteBt
y0KbftQ16qqNzYSCWprbxXu/YVsfC8jOnXtpR8hrwTrJFdqxp+Iq2XCAw5wrYf0Z
LU4EIX5KxqxXUsDmhKDlT6OTrBUWLnVv8hJwUlp4Un6YKaTQseZg7effy5H/fptj
KbUFb5XKE2k/o2xZL7lhfcXcI7asdzqh98Ws4ILfQ93U6a33J9u+8Jz9gDR8Aoi8
7yWQBvpmi8yCEQQKC9kM+NmXACHVUxL2Rz4r5PuIuUacActiXSeKFe2F3AOm70bc
LL3Bj+lyOleAB8C32lkFdE3SYG/dvoxYuoQhBtO5szMFhI9A9k12o4PZz14UnEuS
GZ5eEXxM7yN6g88LKjCpFOJYckAxR4rFh7Fm539xJwBAjIwQGHlqfOac36KGhkc8
q5BTQv2PKkiLdUFS9WDD7S2QMQUpkUtUXs8pRXBk/bMJYPjL6Q9alqIQB7FIee2B
+QBJk4VkgCm9z3uquVItvLvGfzjPFFgY0P0gOXc0HByDzN+eHPEZ7sABrbAchHlW
TcM7ZX2joqYrdz+5sFFwV7ovM8DeFKFKeWUkiikXfs4ruPsifJ5JOkiPCiAB5d/z
3DZ3eT40Uj4rLS74/MlPoQgChjzaqsSAKyriaumaP/DqfXWxyIPsGkHENxe8NhHw
0WU2w//rXvBiTktdTutDndOKWhwOhRSRtUqadDzpDeH4XKvrCwtm1j6RFHxdtAo9
CCZsukrvyjxntK3riEnUTcHSDEcOKKG1hOQTrM1ZocxJ6Afm9j27KLqmb18waXKe
If3UEnksiWwRIyjN6NELUZ6b66INO2M+Kl0H8lYIqdMCHwJmnvhQm8kYCEbzlvZ/
omqF5aa8VsObOonu7JUoS2B6F+CDaaYg2AFsKVWIy+Tqxc4ZN5bWrAmqBZas710d
pL20sg0e1il52haWQLpd13FSN/h55Xx7iVwSZTER50EQdxevuApdCTM6zhXdr8MQ
H5qWFh6CUIgsCVQ+GHo7iTLL9OSPLj0HigvGxqnnKNJMm+fC1G7vR6SLeAV7q3Md
w0A+zrckdraLWVkEQnE/lBVvMbmlkdsPmWil3tXKTKqQgSxDhTOeHRIq4aahFthT
rfXezUEAiR/EIq1lAvKKqkB3hB5XA8OHEmPYWExCaWUBBLlodoGAGoNTMl26q8Ky
1wZgbkwRRHVuhN21MTVCtjM0BV0gSanc11wmYqgU39J1iwXQWkMQ3vKTEndsKdHq
AtZyYCLGU9v6cquZDgCEdzd89cxu3U1tZb21c6tnSNACR1WPlAttz0hCDUdKTzJd
Y7udp+nTXFYggRgQ4ALW8wpS5mo7Pp6dV/jsxaciALkqrvFgBw4Uu3KEiyIqXhzb
IUatdmrhFK8fTi9lq8u1SMPEUC9PWB4TgZUvZoioY65Q/p9b12zbOGovPxXpvvBv
ykRFzmT++CiM21msK4dRpY6ZctDFN5I7I7aU8TXSB5cpEwGhX5kqCZds6S5C+k6e
ihiBcBmzIC4auQ6BoLJK2vbSUal7QCZuD8TxAhNuFaFk/VkLP07b/bVvorspGLFr
aAItd3PRQ/lprul1CFgAE9j5fHQH4f5tNgFZXLj6n+iYq/8RL0QeL7WX0wVf9cJ4
D6zKD4NPQcwqsB06I4RMtvm8HAya/Az5X3q5rpXQhFVdtsIP5r4pf3xCtWS4R15N
IRHvGpiLJl34d4CuDx0VsBMcrEapK5VHXshnpM09icRc5optE6fJeycGY/t1ZBZT
3FxJUR29dyX4RJGnBbQycJj62y0DuFH0hYCvLCzXNsrlZzdfE+uqXTMvujWC7eR+
nVzmy7XKpGd82YXe+RfGOfiXqApKdE4lTofK/Q9c5rlY4cdPl7mQ/lklyZpBq53/
59PS5GELOZPfm5ltzpnJJCaRhM6XIiDfN05bgSTLO4xsuMnK8w80DL1aFi8jA854
sQD8wNt+uy4uSgAM2MYdcovDeHmbK5xdm38pcaIbrXSYwAGhUXvxbYX1RgtW9RL/
yvooeA54kMgi1y8QK6T+cw0S9ztdj83lCNF/NE8kwl1946pdPLsdNraTcER2MWmX
sVidhK1iwQjhYMt8Z28ZnJtHtgKZNxnuH2gIaW1Cz8u7F7V1au3kWlNTFlPZgRB2
k3fe8uoEw+DsiyPh2c37OYwmitRSSSuD9ewWkJc3zUdk+Tv9jtF0lorRAaXENgeK
cDN7/G415KZGPfyWRffCtT954PyqwU0R0r6IqdGoiV0qTfvk4+Xd1G2eq0jf8iTG
UzcBUgXZ0wwEe5bjRPPbiU2CGuMtfibvwZ+qTXRBwUreu1f4rIKIA+D6uYJ9m7+H
3ObtGbn/v75eRUGfROD6W+t4KJ0C0grX0N7KAmq54gP16EuU/ov6yorifybeZxfD
jGD9oSpy3TbVLzxkBf3aQbEStwvTpk8qM1gU5lGbi3YhFkyDWbO9KVcwRUf27UP/
uVf6kvogbiNVUcakqcPuk3wyWbbyAqo32DruIHhWoAOAse+ZOh3HDvNWUhKBWz6w
wjPyQubzBiGAui/8VjINLvTiyOGEAjDh0JL0OgqqeZ78PxltRg6/jUBzNa/Iasxm
J58tokdoJACdMdTW4WvnNZ8NE5JBxowbraBUeNTEY+2u9enFdol/rwdw6XY4BPZH
F+rZDAxxivGKJGvkAYOdhHvnxbm01v/RZX0+PrUrua1E7RXwDXX1FE7Jq/3mHjO9
LBgwxiYRMRT6+RZ9q6zdcz+F2HMGnOf81bBrVb+FHIdrm2oOpv5gb1kjBZ3B7esE
1BezVT42vEbIj0WDYM1z15ATkxv3UNJEUshO83dPl6yCQcR4zUDeuHVWq5bIAGaP
izJZDdY6g/xzTDh+7EbesLAhXWwQWiZzjUO7Ck8ZV/LnxBQyOIV1cTtb5oc2sfzN
Iouud0H1/YqMnxGIeCzv7WQ6Y1dRTkdfwBrP51P0Bv9ZDO0BIA0vyTXjeY1PzNKQ
eKzYLgZmmhej9aVZ9fGYO0+kuJ2oGUGGbhfPaM23dVZBznfFuoki0ko5upTrxPNU
T1ouDIUbL2v3PZQSWJ3vLd9d2rficgNn6CCPLlTQNLuxqv/qdc/hsJzPEipFV7Ll
vneb5U6E1HVoPwq7zmYrTyc9F42cU8yJVsUI2isRyeds3LDdFavfXFEyw1sDO4nz
hXDMQWTH6Z8r3waFwcuSJbzD+cVLflUKQYDOB3RjWJwhYPYZFGP+8Vg7kngNZxpL
bZCHVFoe10G1PJQ4CvGbnjWff7P+2YwbVb0SBG6qeZ2umOl2SiwTv/f5ZOwHHIFA
7cNgbN0eaXlbt564KhZtr4aVTKxqOkEtbeLxVYgZ9udsOYyYfouZ7doIy80E6y3C
Kc9jm5jPXAas0Sv8Y+UIAUhFJGaR2JLGmm3166h//adF5MeVVCviJyJouoelRGrs
ftB2VveExzq1EDreQFjGp683T7XaT2r9tW3SrmatXpTu5IY7MKMM7Pfb51GKu7bj
5kAx9xNX3Q7K+1NId+gDmkwp93L45FQoLJnW6m55xMf+UjV6bgSOgFSaEN2bB2px
23NbNrd/k+ApY39plKJ+nv1KX7tY9Eeh4lmHjWuExVlOsu/WwOq/vrVTqcw/kLxI
ISS1MCSNCPBgGlr7JqeBWAgcdN1h0NWZYTlcL/mWUWANqnpWKU3BJBXR6/lNI0qY
REIpsIRcBBmSok074eOCscicZFrkva8VFzEiUQ43IO0b0DJoiizqSqWm4CEwuptC
0RDigUQ0lD+iBt4oaQyD9qF96NetExTYsC39rEw449eQBO0XrroiSU4QYbHF0OK8
mTHlNAKrt3OqxWJuaiMLqOz1QjRdEvx3SqNXbrvTsAfTQ282dnm8+USDKvyVEoWl
kBsftTgTNTLqPMBH3+LZMc3CctU6tgHFBzQrUc5Nd4KBdwVS5WHtwyOT1GsXq3Oz
IlKOxQixtFcJz0u9J+kns4U8qUb8FVTQ7lgnK0mdIYFjIzyx/+KukXDTpvloBQby
hjcpmnjAiQ5eWJHAYLKUUlpw8HRw1Kq2ybfydXLNXW8Fu/UFfO8prR8X8D0oWvIq
bSBpj8jawHeE1pkGcQ62QK998Jo5P0bCSldVT1VaEazdqJsYOhn3H14MVZq5KdfD
2G4H55g//A7dopA7sMeyCLPOfDxkLle+EafkyYPM254dj1jBbFPxu8QGZKRyLiez
YAtwHLVL6CONvPYtV5yR1ZaeqPZbeXCbpdY92Hti9ZQHUzBvAAUsVgCkrcs/1rXI
QRkBOTkEdd6cO461vTgv5q3yEDPQbJZ1NG1Fu+Ry+H90PkypvkmTMDqpWnhsry7N
G3BbUuLYjFkRlm7iFanM+nkJdAb0cE3BcVIND5jHE6wE3n3oIGWSrND7QPRl30fe
cWHnq9851y0wAulXuWdVeAxnsW0JDb7W6lg3SSJXVGFXZC4SuegoZkdZfa7CTR/2
dicrDASG7O52eheRnBjKcMRR+whsSWuSGY+Y8SqUt9Qasu7oZUp1pE4MqYz9YZ7Q
xg0bb8soyNBN8UsL8YDJXOu5j/ADxKYzVCwqIsEAK8PWOzFc9csJtlxO0i7YBe5F
305Z8aXABmrDEpOlJgcFDTm8kHMrq3RsZe3kIblrOTqzYPOAY6zy6QhwedLHtA0+
Y5dRxYJaJt6wkKK3wWJx6V3Q0whmArMGgiJzJ1VvBhgzcVLHf6tkaxxkOiGwUMj5
vHPnYZ+AEg5qB6IJHcPh1Scx/5XU0HxlNAR4ewJx9dpQdMejD8FvjHHTdYdYOVK5
un3JNhKjrpq+p8nbSg9cTVkqjDuilSBVF3CtQMR+Ghq9eOO4bdP22ZA0H3q02I1Z
RRV5jSu+CKll1dmEnPw3UbV9F/vlQBEV9FiPP0wW4hbjRrMSw/hrb0sIiZAE+7fT
lGWqTeGmAJqvUmcBVwdpNid2txnezTMHRn22bHQ2NfNOdtKauFU0My22vHRS5TSL
mOcVWLNRQjt01lR1PVd/CV9hwskaVdePW7Lzh+QmjZH5adaatsEsHCSwth5xpO/L
oeit4ylogwB9ZrTspCgzsR+Dn+K3Y0ZbThOedxttpXm8lm6hHJdp+LLPtFktm+kp
YXJh/Fnnyrbaqj9bqGjGmGj/oahfyO8u89zd0//XywtKK0p0iqal817RRQo5GGoB
pDCnAxYL94uAlUKyY9fEwQZTJswWvGnGoMjylb7SSlltJl0fez0B1qbbQsIs0jXm
LNtAKiR5YGYWliLnBqFaXC69CDlePDwR0iKne3vqKmaW4UmR3MHhsqPIVO0uzsZ1
bFftpB+sF+C6gp/SWAeDtPDlCVFV0jgxIEldW4/I1BvIHgn9nT4zBFhj8dzgtVEK
84ZV54/j2lnDP6PQ9+beoHt0eGQtPpEyQuLSxUllhIwqduX4iYTzHQvEqm7Gd238
BE8TQzdCjbqKQ0FuVFTxWZ3lv9OzbI0xBsjORiCiGuW06VoXLRIejW2sdMvbeXpZ
U49P2UitCZttFfRP41CHfzxXykydTmrB6DftOKXFtD+TrOgCoGGqRm5kXZ1ubFWQ
r6AORwd89Sreh4suS6tIA32Hm0J93LXDN50wFOjO7J5irtoqFqZ3BK7nrazdTZeF
kVRziNj8oJijvxOwelkW5Hf2kq93ciFFu+YfwgsZt+C73RR4b9fjW28fOGNDU6LY
GpbGHP/vKRMVMxtA7CIlVPUlZa00raMyagi+VNIVMXfehWuD+ZratLUXtWK3rAwF
MYO39Fb7XHyTCo/SKCIusGLXqXD87znzOLZE0iVqlUiCNKuy+NAbKTk+J+/vjNPR
it4zSvD3NfmoAaS62u4ocupAy0P8Pu2/qK2BXtianPZ/UbgNV42m9D8XNS8BcVo+
MiIZ+YOtexMIQRmSxW0jXZTW8+AaURNY4ugttYgsooZ9POGZUAhiAFh7xUFODP//
ojnlIN8sPvVSt1eJQhlZ3zWR3Gj0z4zgZtQwKOMnZmi9GVg2zqPwcdpVAw1K4TZb
QgI9YnjDSw58XuD43q2lSrcg38gPvgAINVN5ka3USJg0o3tdYF6wEuz8Unzg7v1v
qI6WES7RuZdDKIuhd54FNs2ima/r6p5UAY06PDrvLj5NwW2J3Jf5/JHDA/PFp0sp
iHvagJBtXx2TWOa5jQiBa9RoGowVKIjceAGUTpNxVAwpEbdJv4PCFwOMb5o30L1p
GY8rg/5gtE52rdrx5jkqAqz1QknKEVPUIdEiDdSJ5Dal7IU/hNur1VCd09kAG4qO
lwk7dxzTOjg8BULy55IJ1T1Pis6YK6erqJfElt1+eEGBPLoBnXOcYmYFo0RPKdQ2
eUIra8kfpoeMKUgBcvSMxQn4OigziKtxSBkFzR3UjJeeEXkLElsy5Y4lEvs+DLVY
cQPEGvXqT8gwK7gT2uhmlYtR9mwIblUoXWkiAdv5TgMMknkJcQ/fvd0RlYFfnru0
3yNGVBe/RlyGxkMxMqDTo1x7TSb6CvohzaMVNe0BOLRxaQIesJjEQmcRjVfnO/bq
jdE9YqlY3R+5uXGL6kMEdJJPxrXy5MSUTmrXEUwmMPDqLJJ71D50wOlvQJxO2n8B
nSAUtyTtSzGI4X9A5XpgyaL6wPoSCDZiennIIpzfpWq5g/7RN+S+wZk7bMehlq5w
+kpsRHMLrnJDb+MBsUy3Z+pWI1iGCW35dxjBnfBkX9L442RMYOPHEQ2pPN5WgSRK
0wMxy07JmUcz9IVTtG2CX9IzoDIDAyKbYYQH3JjDgV1ZYXLF84oOkCDguig6qME1
eSyvV3gENMbWu5Z7XPdWrK4BmhrzLFD8TkK4hqh43PbQ/DohSi+Z7alAUKvqx8Js
5qeEcjmw9FdyHQmWcBhE8tA6ZeVjNsRi43EBypMSwYS4F2yTFjteXajcde2xZx7Y
zjzNLR4S3LCTIhQtiyNyZEQZVuEpWHV9T8MVhA49LrL5nfpd+2WW7KPHXQaGteVC
hHpVjHXi7d+a/bYApdYx2vrhKIE9Tye6NS2+aOF8uUeMF/O+aiiRq9lJ8T82V+KC
6HY4J2jziiRr3nprcHA/bk0jsJIRRS5XsKqhak9MnxgKUWVV9qePGEVV964vM5qh
nkKyX5JViJlF6sfQvMliRvHcEeGzDOGNieVNRBjWwqPw7TYS8JLxn6mSjnmWl+zN
7+u73Oe2ez47rx0j3hPrLLtUbk8nI5/qqGzy/VEd7jq3utiNMwoxq9SnJrebDqCE
lR2MpCHjuwuG6GXZjmtdzmYOJ5hBlwdVe6/9+lHg+m6mPbIbE2uP4Ig7y4bHMUUz
GIGshszdJft7DRo+qeHhYrP1xcroOuzWkvxtqSqK2oGHbAk6pi4C2Jk5XWln1iSx
B66AOO29gQg6pKTx6KdLunQsBlnG8ocUzAvUf3gCUfAkNgW1mv0w55LewFoA2iyB
6lOI7Qro5k5tr3ZWh8dxcL9S1pREGGdr3K5QReznsQVpHKB1cq4gW8bV1TdiVQ66
kw6zlIn8nc/gC986G/DfOYbf7auigz5LsetJzAB1flomqfj+ghyEdlVInjhgMv5d
9V9AxV4FquX4FAMpinrOmYhdr1c79hneUsxioHYbUm28TjxzzAsBhMuOcUqKvtdH
GlzCUEiN6hqKKaSbfmsETXjNJo2Ch3W5AEcQyQ3HIIiK38keVqv7MJAijvyzqJaU
krwPCeNz/qUgk01lyNI9ls9qj7t4HOdqiQfROR6xgjOJ5qp0xT768oIKD4RTMt2g
E3tIu5ZJpjnhrbZMMB13VJjWSfyBnKVWrHAySbbDLCYorqPEcfeG9f4fvxm44Tit
lAsCApEU7xHhOlG476CB/Lu6PpMDrtq1j9G+yizTgtnC4GXH6++f36MtSfkarKpY
mn0NoiJJjTpgm9A0MYyh/gwK83GKpRW7yvEoxYobgnW9eJHJOdcbRzN1wep3UqV0
lfeENfiaRBIppxP2TfOJxa2/LX7FmVZnJaMZwBZeIiNqsWXDZTPdFml1DZc5+mDL
BJL50+FVOnv18pQ0dvIkqq3WQAb91FQA9QHkbnwm5nZ4NmzjfdGRczFrEiGMz+1N
fG2cx2DipEs4jmAS1QUG3JGVkOc8Ad6udVTaISvB5EoN+ZAgEl1SpraOzXpImeEt
Z4p7Gt93y9YvK8w4fm4/Sym5rNbmDcrFm9EC4YSKecG8CfIsQSCot/nI41SyuLmu
Ywqc9F8P5KPdXOKuihfhKCesCQLdiddZrMIEB+kSCfDUj/criWWXt1t7Nhmronbk
B08Qv70uCanyULNa9byC4SEZk3n9qUadLJDGY6VMxvqhH5LXoJJk973mWDOJrm7b
dpxiPLtAqzGSPzHPfB8QpjUxq7sxCYjVfandk48TCVtXhj4cUn0n9uCadHlU/l6x
UY4vBhZyw1DOM+YBJilpj+PYmmwSQTfO5gjqbeO4AelGHYttFo/OY9TiZM8S7oIG
WsHxmEMn2lSDjRH7B+7N32L7NmlYP2A6rXJbHXXiGIoBnqGHVtkPfunsg/bVHr+d
Eji7XTRRzh9XHJPidnS8Ws8t4hB2p+v+0KjwvfG9HvZNjjCLF2ECisB4b2cI073z
DQGRrnYZDs6588OYg2DjxRVgP5wbBuFhuxNAi3PCHB1I8vzeY2TYtP+clbZKPTYh
JwA7UprOMfP1YfZ9e8x/bTsTCqX9mTxNKchhtK1w3hUXCEsF7nM7pt0ba5QfX04W
k8CIB9fEQ48bFFWwl+No7Pq0Xo99Swsy6TWsu+FOpvQPI8VUU2TBsTFtwYCMPPk/
gszLFEnZNhlHxZVcnVgnRG6S2bFEjpkzUG1Dvgvz6y/biGQBhaPcoBKPJJWL2wdh
wWgeYw6ESsPXIQDwRsS1V6ztacEdMNHoNSVviyjK0aiseS9Tv7lZfagqZlyQex2x
3vey+/WcEvIEz2s7/PfDbezo5bmeBYGPx8pFjQLeXagfL+lwLhz8OeqPhCyJZGA0
T+IxaC0PKTjnTM7LvPsb8lBWRzcausIfaTSVVonIlMnQdDad+EiF9G7KdDNPKx4G
41FuDGDiYq7/MzrJuVGcmMhn/Nu4rrOgFcXvWQjHt3Xo+EWFhQm44XEtaB1MCVjR
5hmG1Wsz+lQFttiKVZwbA9nhIhWWo21kiCXXzFpTgQI2Ol1qIPHKUI0cqf2qk9Ao
YvnnU5oDA08MEhc8yUr8P0cpjuo3GeZ61VGJKugPWeojJdTvJn5AthkMxY324Vvw
gUcqyjDIU8xGRu6mLqhv4qe7tId0y+xv4yXC5rU/lt/CAEgs8LMdK1grnMa6qjfT
t3imaJmhEoUSM+ag8rT7BJ5kB9Bk/86bpTQ4pVo5HRQOnsj6FU68oJ0dJRCOI1fN
Qc8jY73UKY6GBGpqgcjnC9skb8UT7JTmjhSwmfGrt+suvtW7znYbHjPBdh1Ha9qY
ZsFT0RzVEhtqpt8qh2PP9uksSa5tbsiUQwW+ZQYjSkZbGXUJNLVQuqFhB5BY9lJ/
8k1pBxyKM/Z/x3NE2QGLvY9HfMqffWZpUmt6MhlV8oMQ/6s7BXaLcfrsuHW8u2OF
C97FHO9iNCrpTUjFlg/VFbpCad5yGyCbbp44UHRepDEVROZf1JifnvS+V6Ude5yV
mKbtkIbAJq3KGHWCYxqKr2pjxObHer4OMxM8pyEqPQj03xxYH19YaP/To6YPo02q
HXlitllJBG/Q88hedculcTOCg5ER7ajn4s510TIxZLxN04GNNsvnrBsx2uw9lDrd
YokHLGh8HDGsavgFatozU33uXXfaYUv6YVoOeybIPkw7Agx/HCNdS2IzYwF0JWlR
ns6quRbsd1Mp29DjNQu6N2j1EZ2kgQHlQLRnMZz7qpcdDmZeNATRSwdMKizPG8LO
0IwHLbpThBKPXL3qYhjWHT9IQBY6J1unlEmidq9V7RuCxW12eI+nXetKtn5we9N9
6mRogBm7EL8ueNRf2hlTTs5li0YvaYMEHIYPliVGCmxTNj9YskKGKga+giWi10A1
YRC3GUEA8uMtu/zz1t5gNzEBdYJ+FgOOT8lf3145qPsX2OzWjhjrYHQEHw6rJxj+
uAn9+RSR7uo5H72hUNLSILhcf7igONdh7egtopZvkouvwrcxnyl/y5t7/ZHCp53O
4gxTxPVq0gZT4r5/DhVFsKi4UOBlstOnI/yq+s2zUGkD0dUDwHbquaT8vGfaPEG/
J4hXSXYnOC7T97tDdygteoRWWZVEEklLj8RVwnylTBmz3TUUBLlDD9+fRqpfb9xx
Vg8/g5biHpDxDhBuPKD41fUYBmKq+HEKgMCzSELPOMCDf/+dn9KWeRNfdoCOcWV2
FfisOqX0V00txTnXIyuXIzopaR2bFX0+rDCakd5OC9n9DnEaeBFgBR+ZObPp9LkC
o8kTsM5XpTr+uwn9EULpW8JSZgjVXpbUHEghLflcQf8neWw4NMiEa/VSKgc1ksNV
FeESS8igkG4eYCfjFHIq2zYhhu5ZHCSxW49qxKwJ5eQrKE5+hUR6vvAl2e+EN1RC
JEE2TUjDWIf/6mBp29+vpj1EqrxGrfEP/r22UZcwpE2hawn84Xx7n0a6ZtvuUlsG
J1flV4acXGJU8Z0bTaBXm9hiC6tuIlf5VGw4zsWcqhiT6rkj+fnlXgMU6GYDH14H
+k7mFblzfDHYDGDAm9rYP4q3rz5qNSJrs0UhQ6FakTUPz5Hr3vBL2dP1dsI0FEHE
61j2cvBfTo0Lp1n2VlSib5Qctn54whWrrYJpdWFuzH+X73+bLlSXIXObjrT9Wz58
BY0ay5olyu6IkbWVGnHDCz9t5wWBaBvB1k2iKihIP7LR9mqAkr7LwnVhkZNRt6rW
V7erDA/Um6Yb3OkF2kAv2jFMk9qnrY2E2L45RktONzIpGCysRUIyiaX+eiUh8afG
gk/P9rTD334BHfUI77s5QmJQwmR+yez+GwZVnevOb+hI2p5rIgXprcUeFlnYGge5
06WLCCNRm7BF7lzAS+zBBAonTfxaetZU/bdL7Cj5NYTsPHa+yP1OuSZPP+aydJQ7
JoJzL45/D8rVnoBgbpDZDC34xKv5oMbPhSzl3IHmGq/JhQY4ijconeRyh13W0Ox7
j5FWxzBnzWfFlr83DQg3bFph7Pzwv30MIQMlNxEkO9/miiEN3nwHtWqbOVG66qDO
ppHdwoYdri1ECi9p8Jx1rEDxfRxOIJo/1lrRqPM31xOBdvkX3V74voiN/fqa/8uO
chHExcubVa0uKL7OUDy9gJz1MfOshFM8Ah+goOMzpMPg11uhlzw25JC4V4S5T8P6
QtIVU3yg8Zvl4RSehj8YEAwOifmQHbimVaubEVTikOVGizNSmn8cofITmYscBjAq
QLI/OdvELH/BeivXxFCD2yz4LksaTI0khQlILimIcNedC1hliC6i+DuyVbGqzqte
or3QnIAnVBIwlqxUVvHcoEvOf3vQyNpb4ifaTI2aJ0kSRa4ipF0SBj6MnriiSTpH
XC6m8ae86OqB5K6ZbzC4NxIOT5E0ytQU5Li/FQqi70yaQU3gSnfgo3ILfZt6hnNk
MlUBWHjTe6TT1/iIVPD+xVy1eTbhrPBo4TdiqAKiBbqk/aQda2D4tM4iPr/AXUeE
pRBFIt86g5hI/7kN0h0Zc4AfP8s7MTWy2G1DopJYJ9cg1YbggnZzxyCYVXudrkpa
V0Di6rAUGUZLc2Q/fGuOQXoS5lV2YH+VGE6JCv++p6ICAhWs7PFDdSdZQjYtgflu
9QxOXYMuqEyAnP0JsVRN0OpOfUGjLI2V2riZuBw3E4wlReCVm/iglJeaKjdy/3HN
2O9lsh0SX+3RM2tQwPMLzzJf0kQk1VvwY1uGM/jyOWBAviMH432Db57T4q0vSFii
PhU2fNcI1kTSThU0nXEVojWNN9ocbaVBEUQQO9PMnHLAjgJ9c3O72i8TEzB6s6Os
TTHKQDvcjFMpRu7Zvej6fH5+z6JmmGGHxbr1l6YIKeRnODSHgI1WLjdw6VrLclCW
AgMksE3lOxjLBmUAWHuB01Vn5Hm7CUiRUh6urrAdrqX3IEVF8w1mjGL+DGNZ9Jf/
mCwrbBzCiLSuzYUm+i0KnnaDNrOjcQKvIMYcn2V0y2u0BOFfZkvEFSihEM1ZZmou
gamqjz8llpr0iYDofLckW3JWgzVqgfFNpdRLVIVl9gpsf3pqLZBfa7aU7DUEAhCq
le8efTTaUKerq4wf8oveDQg73RRyMAPEOQmAfUlona6SNkYnLVC4/QzR1UVpc61o
TBsF28o9Dw+9YT6oS5YX9plUQQOc84uI3NkHvjSRjOq88gmjj1VFEoLllbPd7cx0
TmqYuXiWMas28oVzQI2Pj6tThQauV/+0oprcHJ0L6ijgIcwzs49SNdwXsxpG2OhY
hDRTMhzQZveR4lmzid0pEe2bK9toWNEwPanw9VLMDcokwgzVClS06IgEZZ0m/83+
9mlV6VM65eLt9D9ypXRNziS6hpg3xQxiG91JsfagVaqZ6SOm1UTPnLtwbXtqeqMk
nDOfZWZvPKU0yYCXat+SoAPCHxPGujhfPanRAnVuKcrptHzXVR1Ul1Svv16gdmqN
Rruzv1idJ4vjqTg4+9s6xUqaSjc9QQtdcdvdJZeUA598bY4p5ElH47M4uiHWjeNh
hQbpmXjM4IUNf+x+SPFjP65vm2mlGczkBf+rjvATokuKSxsErEFN3JjwkndUVaEv
vUgtPnBCwVXnTF79jc92Zc5vJIA4GAv32qqfGmbIX/2DtM1/wYvX0qVoAHeTlrea
VDB8kVu6yjrF0OazDfgNZVKwWYB5eCWvSBqF7H4fABjAwhu6+xEZ6FW6VOVzpEA1
E5rvWRki2wG6FCwwJXBm08IkG5oYA0j+l/THo7kjxS6bzyiuU7NFzmHj6a/3EqDl
mpU+kqIiol+KuaSv1jE49YPiGtueDuwNkI0Vu58p7v6Bc+pBsdsxcqY7XdDb2IGJ
AHCPjljtKZP/iidBzoSuPPlu142ZwFIRnVrDcVSi0ti8vz1Ew3Rf8HIuXLsE5TiB
SUp1Y4S0PFRuJXRV9oNg/AtzJBvECxVlyzj7Mf7FQQFajZkM7Znrx5SJs4pQxTV6
daCTOkHum01lTSaxfkJHSbnsLi7oEgNocshTmhWnf+qfaooh1RixUNtAs63eofNA
AujWMMlTgp716qmZOQT++v3qbCRqT8zQ5m6DCOvvsE+d8DujusfLB/RUyGwSBGW9
qeFyUdH2ocobHX81IV8ox2Isg4wVhfUD9wwNoWuH11tGnSSf2ZNhkLMb37ZXbGKj
NIFJuUBZZmCSrLtMNJtcvd7ECTUy+89JbaKMNOQN7H7aQA75HHA8D3Vk363Kpk7R
ZVeUFfelzlNXeQsYyFpfPgSd4CIBn25+pyytmBTtRu0YrXfDfKRh7M+QIy7hsuqZ
8KhaegbAxKzVmSqTljj9JUapo9Gqt1k+tXuUWb1a3GFJdxmAFIFbVyTJZKwtn/Pk
2zw2g3St23UIKZxpfHbrbptXxbW6xG0tgjbJxH43fkG1ifI+WGZCrPa8ENtPIWzU
oaghO3C0SK0KiGiwBx7UdwCEVZ8dVG++MBSYg2zGgVkkwkiqmjKpKzTPR+yc6TQ9
ZPAQcbB/jabvxfFjv00bg8PdO9+XN9aospIiHCuLX/gBTN0vl+XgYnwrX7ncG1Qm
NfFwjnwajWG8/S5QCMH7O49Bx7Xaq+uL9OzSnVywqw9yWP7piSpq6cQtw4iTXPEt
yfbrH/koxLTiL30D92WqHc1ueXD0xDuyzgtRrmoA5gi8gr8KgFaaU8sNIEahWKka
3fLmAT2DBD8nKY/aD9EI36NyywsTQaa6kj83sJL0Vl17Z452pADwuwQenFuRgw1+
LTI11oIF8syMEuHFzW7fJRnPWY5kNGcNxBLFfbpxbSDo3iqbrC6RNlFTtFF/ER+d
u95cYklq3+bckHIbqoOgu4x0R4CQOaiSKdIhKYbUVnhPw0hCizhWPGeKHkX4qrlE
sVOhVbxM6M5TfF1XbhdeTm/oIrDKaNIZHysjczqlKNH3MrHnx4vs++1gRd25abGm
gyMDY5L5FOelxH41UiExlheoOdpc0FD2FqCZPEvOyEDCaqTZJ7p8ZaX9FLaDSdIo
YCy+CdXGReIrN6spITWVXWfyxM6ahb0weZN1RDdCnTlr/Rp+0FCjWZNBnET/G3DC
m41M/vPbgF8A7wHtnY19D70j8lDIOnxebGpur2YT6PLwc5Xx5IT1mBJ5XyUv5u3d
kfOlyTQl9/gnSQ+pAGiMk8EMhG3pWRCklYuG8ngCRUZeN98yjmMdjcl6WFFxqqXn
HGj2FtLyRnUw060/AoEzfW+5LVaxHSyp4pQpBhGVR+cwmq7v9p8u6+DI8/hqVg7c
OcvzNKhpq3XQp5Ctde2PmW6QNoH8tXqoxYi4vQZfOzTy+ruoKebE8Am83HGfzxHo
oK/1avB/uS+ccUjBXodKnK1576ssFpgvmze1ceu9S993Fpst48blPYzo1wrM79GB
SSPgr6N069IuNPDhZkuQ40CeVD1OtqsHf3D1n2RgJTMZVwPMYOO3iP3ImFUCffwG
2hd86pxn3JYvoqTEvgT4iiLqNDyQfO99Hg2TG91KpHkWEuve1dWHmLeabBjWPt8+
XPSwbcb5EHRnxVcIZ5XxBGJqDQqyU9HTlAjrsuNmiMD4MuOvr6EPy2tNVEGu/LBH
Sa1wRo+u0QVscb/VnwftlIZeK1VmYFBTAHdLJwPhKEQXmd6mANQebmRE4BdVEEPu
DBU1GwhS5yGP949Jh9gp7vLSjwjnkSX3Z1f/rOot9YLZwchPEPrKvF2BewKR4Z5S
v2oulkB64iiR/h/ZKdewX/iPLXMRjRQSheuszs19rdv1SzHfbgnd5IeOsbRCdiG0
iX1RjPoWP1C5NVAn2NqlJBiYKdGvzWsNq7OPBEAU7YkssrdsGITJTakLjGcwPcmL
3L/lC30K+9uCyd9cjgvCRNo4D9zuZgOiaIpx6yGFm3ol/tUquQnazzjFTWicihxr
al9YqVnTWrOTIdGKYSeCirS7SjMzvVF3PMJJvBCsWGkmcr0pTaNeyS0wNq/pm246
/sI23BAEpa+2/dAyB5QjOSxKpjZ5MwD0gMtztiVrX+ost3T07YxevrxNs9QWvAmJ
t0N2c2M1Y2AZ7UdwWcoqnzysI1XRAfL9TG/XuokEfolc+/ut/WfZvVnW0ppIkV9x
AUUzq+opb26AbFhxE1DSlzshnGx/bJ0fnHQh9Sr+sRY6d7jXkxJymVh4V541dGeE
1wp0I5MHL3DpE/lSY5H4dxjbGZIMvHEcgtXMHNsl0L/e8tcj4SvP6cAMbvihoCyp
CS+wVvCKPgPxv1p2pTcQEb1vaJa2nOHLfWJPB6f9kf6UQ4oMxwqP34bIYYLwvUGH
eTZwcKBy9fR6N4UNZgh4GzLC4cZ8SpoBzf4Um++GJKvZEjJh9CeJREm1Vh54ckgq
Dww2CORK9UK+NLRT5eq27rCxJGSqAXJ6lbPinyEXkpWV4ZaK3WufV7w/rnhQUOOD
aMaRbyeSQaTzgBdRk8vxOAiDnjbIehszg79B/s16hqStAaa4BYv+YFIHCSr+qErM
coWfyIw079ZBrmBGj+qOpe65RnCbw0yb+dFXieBX7EW1fT8lIAdYBqseta7JxTq8
fSiH0jxbG9LthFBkPN71cHRtw0AM1dsgj9Xj7d0OdJ8ngeOdi6bf9x55oBT/Spte
nijxMcD3h+IwRWTMve+XXhmIyB/XH8xDOja8qa7K/c2+nkM8vMflhEei5A84AWln
7TzebedOwPtXXB2PY1wf8LFSaDEryKKaE8JK1e+v3UjokTnV/eopLvP61FyjWb1d
td4ItR4IbROYKUK4pVU9aTremCQac954lVZOhekTqaGI7GsRCdWpOeAKJ5CYllr9
UsLxigAgU+BG62ZFOpwV6wm5eX+KkC2/mNzHhcpuIHE5y3BhckzDcI2amAS+yj59
9RjYlhMaPGBk3+4dklDxwK+mCZLNebdEQoqqBWJvEnonwauInRnDIJHMZAuqlsP6
l9XpHoe2OBZk+bSpu4kNc8WTY9tytN33pKS/kqNN6i5EDVRoBPkGQmp2n0/O1mh3
gaCPFKx8+2AWeUzNoNFaK+780jazGoAmrqP2qr+WJHffQcM3BC0JKiIK/wVH77oa
DVmDeanM8rfYgYUrbRRtenVGYu/7S09zQqn056GbYx3mV2PB7+WTjvxT8e/37AfI
NqDdGhNTR8/H7tUNGevlQC0xecL/Rrd8Fs7Wu9SPcX6SGCws1DyA1+P3KAovT36n
g1/IDFP1fnz5hG9W80zTRh08OC2IJS9NLTKHZxbfVKo9BjG4cZdENF9QP7exxIF5
vsSWBksV6k0G8UL9LrDy/Xyvh/rtNsEeffgmYW0zNWspmpkVnmYx2gwuC/URfdXI
b3rS3HI1qipGtEZHw89QI28DeMi5HUzRUSpGNwkPNExkc9veO022jH/GO6IE2m6L
WQF0ZsK3mAZkPndge+577FrXItwDO2no+/PjnGCkB7qUv/r2E5EVo+O2Hq5J78Zx
CnPdjCiU5IlMc20jFnHQG5xxqJh9PJvGArJHTAtq7slq1UwvHBvHBqPqBulTwb0s
z+6Mjz/o3cYRnhZn2mySzOFXLCsTZLnGJXh66kzS96uEk4LCORjmt0IBkPUOiqQF
WrBAk/GwHgJXKFHI2n8jM9FL9M+qIMXWa0DVFMEDcOrvZuGfGvsxBVh61m1BIjz6
fUFMcKT0ppvtRjvCBuL/F1NVkSWNCcHsDYFJHWftBjlsrDNeUjM5CUDFVYMlSqHH
oUbPRajvjdoHV8DhUTXCCl9dA+y3PlSRRc6s09rzQ/ABm6HZmRqyfKYuV5g0R5kx
w4WstrK0oIk2KMPWg5aeVYhrOP8B+VPV5S06XSZKNFp1oSra2j7MDuRXq20a2Uyb
8OQ4+F+WxtNoL4LUhKWrhDmrO9yWbsSPUUVHV0UfZ9LdS/NP9K8lWX/3sAHSVhaP
ZI/vG8xJJgKoOYkzb/em90Cksd7aSA4STANq25i/I5/OgajQqCfp1BAlkdAlNuDz
cXU4ywNEz10PydCQAzE+lZk3P1POwwGdpKATUs3GbKprsNKGLwqaO3P5WWF/yYMT
/Ku7S8Zzx0q79wb3P16bcDW+jWg0mx4ILbMjYHXAAtzSojKu+EqxRUuqRqUYHBj9
in/EaNTCTVDadFN81UbiOqyXPZZt/7CpKg7SmTX+cG/+VDJW/Mj3dcSj97lNdTZF
cswlo/EBTvVV5AFpbaNMgXjUmmwLIwen1JncfrW3gah18Vn7H1pbh8/iltlc7/tO
Np28cRnyRRRZss99gUj1wM0gjZoPwK56jjZaJQPGMBVBpgGwnZLve1NRJwPuiIZy
hBgC1930Oeb32EgiGPbEsHtxjWxj2XN3X6n5waEQlgubS/4/hgh+Hk3p4gv7WnJD
gXqNBWEd8jwgg7fA/Yy0ZNX7SmTWJlz12FCGbJKP0Uj9Cidh1GMAgymV2YftgMr9
yzwyVllYPc1i45Mw69VdUhB4qKrGkU+0MzvmDIiivhtVJG6fEovdpXRo5NhAoqWg
9qv2YxHLH/z6Lqqgeee/O7/lcTrpgEwmXrtPsIezJiHbh6l5Qu1jyKZJK0eVDtd3
jdI2dKZbesDbl7IL1df7wn5uJ29JX8xILC5hdz4roV6M48yz5MHXaTLIDfn3aEe9
/2AAAYScl4VgWTn9D2hGx0iLzdgWnWmrqHWioV/0q5VMfaFmHlF5VltX/BmHGvNN
31lpZRtPLAzYJlvCAVCSNo/ZhdMlEtWkTmHKFd+VFEuMpbJyhNKbH0MIS568Ic1N
ienQ1HFEgCIpNb0li6x8LqmMXstX17rm6nHt3cCw2otf6fsBxkwyesK6Xv04P+JC
7exXC4xyB0y7rbmXWOlJYQYzfJXVhWhIkTvm4BS1DidpmV5XjF+M908IbrTGe/YA
Ji0g00Yr70gUdptp+AQAINzw5BKUJOsuTQTJFVIN/dxR5Zb/q1+e/4MAb2zBAGPr
JunzEHAsWyCUHrIv42vinOODmS7eOUv/iT0hjbZaGKXPuGwzze0juZb8N3zzlN+l
+GR7WFjZgNRca5cD3KQ5B43xUBHr2yz5GtgvZcYVix44OKSuHXoVG4c4FQHof4yS
MnsWKIsjaURdg2RWr7YiaAdGeXO+WMURoP1AFppZWgdrC/0c4hoOmsG9C68aJUKH
zMKjuoDQ7aWs9B/MKcytJ76oK5oAwL+GkHLYfTVqaexXVclMta7Qkhc2iF36yXNJ
pK4QmriZWY7ijFLit93atRddPloL8TVM3Z+F6vmifKhPBmnSAalXXqhqtad+YKCN
S+/9DmFUGUT65Mx8XZ6TQVTIRa3mn5NAY7d2bjiA5/asykKld1cpmkhW5zcCLtmv
Ul6K1u0uOBU/IvETy5yreRQqnfigpf+TLP86dz4xuBpQCM4nsYtihfjxcPaypXMI
VwGH7EjaLE4Zi/DzMjayALPCaZ7U59TBLaGQxjP1ZXneXxPTq1qbORTnFKjew8je
ZIs6etO3r58FsbX56iyLnuS+RQAyqlLD+Dp32y6rLqa/oKcvGy/+Yo4+lLFRALBy
58Yc9SZRlfTnxadVA49uqpyz4fxtprJZPiibV7spj6G88odLAbdbRW2MkoVZSZC5
Ug97Uo6XLqQphPjFkP+4TxFg6MRqOxfQU/UieQ/+jr2c6xXoJOUay86ARcMmivFy
bEXneyYZxStYlFG/LTFItUM9/fKfVvUbV791vZwIJbOLFRUQ5JPXfjEpm6BfFxgS
trBfPep7+0ldYuiLehPo/Dp0GuxVmHxhFbbzYY7S2ikHiFKJ9V7K6+Yj3v5zo20r
gYx2BGetOcJz09mwkVOsMBxX4BjCyfZJojRAQ64pyB5Yx3ZpZXltinh4fvombE7d
K9t4/IOmuZSu9mpw2cKtBOWXJdPDPikrXXe+skxIsKjDf6d98bVt6xbSKsPYhLe3
Um9fRxkZcBbIGcs7RyaeJjwgI1SDOtxKp+leIjVE1jMsyytKJ4w97Rp8es9sehOe
ZMhctsJqQQwnHvvrFuVuTsTqzYXGInUvb20JxZ4HtzFQ07ajd/ye6VqBPEgQqt6d
QpIPC3JXkAF9edqAfa/ZzCha6bvI4njFCrvEYOtrsKzgKGgIyYezI/52tJT1Arj3
BNlXautu+u1poOf9khoedO4brlxLJf2VAlj4vE8phniAtM6D87xs7L6Qlaaze1oA
8+rcjlmEwVkw2hPmE0VzhgHBYTD7cfjuOXAokTXns8gSwb87Ni4XOaskTodIlCxg
JFVjY8adJ4rAym9VA/JubI225tG3epCqcknLC8JO1SjKmWgEOlKh5QlLQd/wR4jz
mu8p2VvVz0TnVpkhoDaaf4EpAiOb7UOgODh9OyejepDR784l1zyCgN3zVLPgnPJS
Y/xrkPIF+0fDlul/1TZldcCnhQWnw1lXl9QHF5ed2PmGv0QtTPxb9REgXAnuzhkL
Lf5/TFJIhT+8Jsj3Nc32I2u/1AkCPmMvoG42h2wJoNFnCA94mTfsb0Phz0r6d4/+
HzMhHhYrr7Cj7EIuaG24tGQ1fkBahMp6Zg+2ty+xgyIUkew35dNeHm4B+k/CbnAK
s4rRI/Y+iM5Rj6RPiEUo2Ho6hjXj6R/5fYwmzH7+hGfkwH55+S/JE27pQ9rHFEVF
+3xtdHx+EueJuDEVlPAyMgGYNgPh4cj6CyPRzhXQRi5WzGyDbT95VPWMqVgEW134
LeMS7CuLB3+YTlexgiYr16cJngmZH1GHI2zzU/HGMAvoQE03HuGewKV1qCYwQmvk
8InaQ2Xm75iOA0WiUKnc0WyptzAI/rhe7XLAYqJjcxPqtK3UPk4cY3qvF9m9yb9q
JFLIJcxsZabUvp7K6BYs1BxwwQaT5NBCJB53QkCnqSdBZwtjflATBbFjhrClYEid
Ncv+dS89dxwS4wzaWepqf5klCcEQqac4FgPiv17zBWVdBnHotvUx/+tVkVGQl2tq
xUTAb+0lNByExS3VlbMo6pzyIn5CiNNijUGmq+Hzl2RYu3SCJy8wER7ZuK2ZG6mh
Vrfffv2e/t4Fw/TG+4dEOKXDcEhN0KNv46Qfepi6ymDRlNW9USt++cSF7kNH3vLA
J9TbIyS3sKB3UFy7xl5U90Cgia/xP8h7jzBv2BkbGKTJNBdM0WUT4HTfeMD5vOpl
I80LgiZm0Fuiy1aGfIYSLdX/0VxtfefErvwG5pJx2VZ6uZEF2+upZxlO01n0Tfx9
p/YlyRSytZYVAD0yx3l7/B5HzL4zI4GSiG3KDZfVQqVEJ24nm4u79996N9WDagJQ
OJ9AJm3fsVY8xrJPNJGpVYXNqhVgC0I2iTpV33Sw7f9TNizpUyO7IVFAv4sjIyNt
2zn67G0LN07sU88OlzuqPSD9sXQiCIdycbS5E+eXrehkwLIfwNNlyeTxyshs44NT
N8X051WWb2jnPFIqNzOunYx2PYI1+JegzSFjTVn3GlgOcyEfnjX1fVSV/Eq0qEqJ
8vUZFJyQZs2CSpAFxQVvxiUpA6TZu9TloHsVcw8vSIOeH26iVKVV0l9gzJGjmrvO
kRnXeSZPXNhUYCpT4KwlP/OKV2dxybQLO2IYuuV7ZIdF9OHpayN19IBmBVBTjpKb
gM2VK/PIgsJ3pDbZ/qUFDxlIZZzSlThrSNJjrJlTujkAyVqAmqlyyf5++CS88RzS
v5r0gjyBaxqkuOOUpQdKBRlfwXso54j2vXLmMfFlUibVF44zzqOdi2h6MvRfBozL
OhVnyABBFMSasUrxZ2CzGQVjIs+0q8dgHFkYoMtJbA/HHTPy6YiNChtUFsfbbp0S
orWh2v0aHiFBhSQu83UXNp14L+zZY9Kes8fIbhprRmxBhGombqVPWoP2f7oJkiAb
ztiVcyZEWm79PojpLdBVWVb8/tqYpZy384b5T7BknWYfLCDuXBZ7LS+cLy0oyWtt
JXwmTpgyxcW0rh850w3sZul2naGkxfQJMArJj4AGqCCGLYX4ke/pXxHJCWXQcbma
yC0GkUipZrQi1aChvuf46u8gszXtmeULIl4rOYgU/kCI3hE4AvVTrjvvnHb8GrGH
M7J6e73Tpyli5UChsb1Qx3v3L3cpIV0R3V+qWHida/Gw5xmsONLkf51PM4fCt4Fo
rIbPkOgEbrVUEp2qUOj+y54/XmcPrYx3zkrHhAqSwJnOdpZcT7v70VubltlujLQC
ylNLsVoka1wXaKK+20CxFaymHeZTt3QbkXEVSVXdx2KfHOW5L/NaESXSnhWjDaGo
yBxU9BbCd1BboBpZPS5DPKlGHv60JmBJYZ2zrpRIeWSJQr0reIXHzzxVWz9i3hwZ
iVTr1n/wNWAWx00604qzltDD3edkzfUiG54Uac0sGXMHe0YRmpANt5eGO/+C6x/H
+sIEyP6Rz2s8jnp48++2gksnSqgVe2+2K/K135GCkiEcPGqErZBxTf1IHe5H1xJ6
zcBWU24OERRgmE/Gdpuk/ldTY3fsZGGNioqz0H67rwB/TU2zi1FKDTxUI3wAOXSU
7C0a+g1bsebdwLpNDDjKQ7VM12/2yCi2d6fQBCB1vu//cYVi++5MZpwQdL7NbVWw
4vYHq+bKzAnPQZOQ0wSDBbHlmOKhu/koYav3OT3M/WtitlIAfZJlX+22MyJg7vTW
dBxJPBeYZBLK39ImolLx4Vmap56abk02taW0bZcEcyVKvhciVnRM2R8KKXwZLPgU
iIga+/42pWEf0aKesW2mEs3bJMUNjKffICgrJo6ZJ/Q4mdFKIjKV5l7twuPvpld8
YbVt+/8BkboHJ5lDs0YtM9qOuQ174DAJs7ZAY5UBXFp0THwfYr5uNBgbtmpI5KtS
POaOOTah0Xhn/SI2FlFcZKq9Egx11go4wCgBDC6iroo8djTGrlDHYx3RrOk3z46V
j/kZq4wg8KpkfkeQrFKXZS2XE4liMb5s9o86bLmpa9hvgtST6nZHFV6O/86mC0n6
VmFJU6uDssM8XXJvt7yEJjvYo8ghwcKc525gpnagzgF2+m5FTIQqTO5QsdxHdTMq
3O/T072CK57ag3Mgn2M1g8SGyDN76+dXcQVyDRZE6HtLEv1NmOJkvhgnKZ7AGbVN
Jz94dAydbR+IFWydn3fP9YhGYfLCypuqHiwvOHQTePa+nTyHybYlsaWCRV+c/nn2
Rcl1+HV4/GcLxYom+/fT3gmVWrbNcG37xHVnH6kANi35NG6BvZDPsMctCkDKuWck
eP6DTy73A3wQ3JFNfN5G0aG7xRuSSk35inQq6Q7UeZ/0bqBN8Z5Md7BXpvmM+ND1
TIpg5v2z1T6Y/brZ9NAlZdLKBScUvVQY4HCw6JiarB4Tk0q/xDLlbjcPxr+X6XaD
brpdN4M2yhFhh8mNywV3ppZCeimHyeuWBCpmg75Zbj+lpQCtZRpvVGIg8igHFtC9
p+mPSIugVbKk1yvSKcP+nXcW7+IxuKabCixAuecaNKJ3CA4EC2P4gnM2uMNisqOO
yaGPl2nzmcgXMwqnPc4RKBQvcGxwqffTem5MZhyv69ZpUNyBtxIEABt+YcAqiz2G
3alcW3nursCxr6ZyibKKADVf0iSMkpoCUqBS7z9HIb90xoFtvGaM+pBwFbw+Ggs4
MHBO+WIMXVxBdZmsqp890wAIFuOX8qk/X41D24JSzKtp3BIfqeojj0O4NbkCm/hk
Tt42/7dj8mItt8ULvoIMI8WTKO9gGnbnlTLkrRGWBe9JsIMliKVYjqIUc3pgYu1O
g9jaacGfYK8JnzzqRkxqvPLluppgvYb+IuBMPFzelbaLhQ+PnobxZ/FicVbRLMdg
zGfYysimnEkOIq0jSbQ6z/S5XqIIgonYDust2d21RlrRe3K3kN28C79EWw7Df39X
IUF0sM6AhshBpj3lVVnrhHNcbUqia/pgfTnpSJVI59nCnXIvWbpaTkQSfKYDcJ+M
/psFVDqxHd29PMl2f9VAwjA3brmxmd9gGZy7+NBkXIDzqZZaP9vy85nIiPAxk9kw
T2e/pl1rcmbO4GYetL2At8EC8Ia5Wwrc2tSYS0gmKyHUHrUyCo07r7pu3sfeFPbu
MiwWGp2umnUaYVsW4TDRD4ZW9jmvleTdWTjSEzI6ZeJuR+onNpI+RqrUQqh891xV
9g02cKHAKK7wqrVNqC0iO/B9xfetiaokate+mfvY1/VHa6OHPMvTAjtRHk+mzmYo
hncDemKbSlPFVbz4y2+t2tPscLPFi1isXzO8pyBDdkKYHLTc3hE2ODjJDMNyYsRs
7dE1xdMGsTrSntQo0NNJRCAKBgbFGKFF8jddirIxgbLsVAYcWaDh1P+EiZ04wkoR
7rbveeZpaG3jhe01Yci/N/6+TaThHvfwY6rRIBTjOOR4gOxrhkBNzPzk2kwI2VVZ
Qax/HMB5S9L1yt6kDV0UA7w4fAykQTi2D+30DhwcubSMqlAwYCUNEx4hn6QPHEKf
104BntR6ztLJYi/GMXhxvBw2mACIvRFPrHhkWnQKyaVLLS1DXaW08zwzi9xgh0Fa
9fpoIiqkaYh3jI+aLOlYf7i0q9XG4Nm3bpNgUGOMIqaEG6ZGFImbMyaNXRGbfYHj
LMS1ZloKY+q+awi5dzKtnu4eeNU901lTvjHNO0H6WRfv09aowb+C5hxUubcQ8wB3
beKfYMVOsDoZzTeG3ThYWMcyM5wx9kcygzNtzrBjGOFrHIvdZHorfAW5kxWjeUKq
w6UtvGqLujihMuGmHXQWNQr7UT9N2o8/B/0C96a2K3MRtVDmxIqZWD4XuN7RLE4x
z8IceeQU3OOnnP2xM8901k3GoXsW+8AIrW83kpl43equJqDFgobNIE++umpBrlY6
0hv5VhaBiS50hrO0vHbdVvwFs8kY2r+loBO7lTem3SacCE3BZoZw7+NzJghI7pZA
0ZGSsueAULUIQ/Yw42kMxBN5I67XKHBDoPnuX63KQnbWGFRJacMzcVKm6qdxWy7R
z+8p/IIn9gweS6vMLnyBrudUZblOkgok8XvjI/k9wCQqdhuf9349HLlSq6Y5RUsM
WJY9qz8QtKrGFrpy/km6Pw2FZneMEJBGA80jw1uAH+ECMsMJ8DHprpGpIgndynjP
GZc1JH3gmQE48g2/bslJd4uyRVZlfJRn+9uGy7QXsLbCXg6rbXfeN7jbqKBec0Ga
uGQGD1umtwiGAOBHoMMAZhKPt4zWqTasmIXDvUtP+R3SLBlrwg6SwrnCI9g4B5sg
aeaKPWijU+zUr5AAZ8FaQi83SKzK/UHjrlKcuMYq7YuVdEDKSrB4lrdbMw/9X7qc
NsK2zj9vhRG8TmGcOR8+okvuooPT9iZeskDf9IkFuHO8LNYAJG0yhWk67IJkXMvd
KiX1W/hPkTVY2azoY4IN+R0fA9H/t0ApcK3wtPNG1WBvwIKmPPOJ9O/pg7nWqsDs
XxrnQaRgPEI1eUQYWCArvKemNvNo9vI6nHpT92QWynOVJX0ad4vbKnYLHykme6I3
z/HFLHWDxvYQHqpI8+YM9spEahkv0TI8WtZK+YGksvRtRLJggptiOgWtiCtr019n
f6/5zSqE6ZRZtIr+Gjm9vwUfd0I2WprgHHKO57gLgHjDtKagjI41bkkomkRSV8RZ
hZWN9CmI8a5lCdHQpjmBBhY/Cel8swQikl1kDOodVpfzo/Z7vgGUvXDp6S00Zk+Q
TUe5sTszxPtxFBcoKuRDR5WZGoUfDBwoHsbpzOcC5ayp7Cx0gVO3VAVCza3AeU18
NJ1PcFK5829m+BneGgGLt1W+l0HwNIsJHCJjSJ3m3rD9d6DSkzkpdjhL17fj5mEv
HVj/zr5u3XONlyzneQ6+F0ln9+MINsU3kwJAhkiBobkvFEDJsPmMGgdjr6waSJoe
9g81JAPBRBn7CKNHbXg6BF/xD7ecSvokXyQWr3VelEG20IdTgdFL+4D4CHB1WgxT
bsHCuI3GSBxJ7jEJ1/rkeGHN2XwX1ycPCUOpqT2yk2bewB7+jYie/THGS0ZII5bd
mPnan+7VvkV9zoi20AjeT9ryVDfY+mLtN90s5X18G97zjjYZ8n8Rq7AyuS9EZ3Wl
U6vue8TZaJrs4yLQUyv0JNqHGhvvBCwjORbqctiaxgeG+BLwUQkOwNmF/2I6bnAc
EApbu1ED0og/OY4HMpV9Mum65/3PloEK2sBCPCNCCSNrGcImkcPLBnZpHS57erOX
bXE+a3B5va03JaYMA4/C8smybqwcRwI2ikCo0RFfY7vjGrL4mQ4HfcbxRUOn83iE
ZTNIEZessfG9HbTc34nUlhqG/X71oJdK8i+MzKqcfSaaXa29D5TRzrMq/9X4Y//q
5J/M6M0YEqWcKR4YmEJPsOIPgAFOLfKEHmf1/QzpbgcIUHCNOWOMMy2o5YDlZbo0
7OrqOJJkKUJ1qZ1mxM3svlRkfWN5Qquq4ywpqkw9wmkIOnDflvCYd67/UJXpoPYm
OmDg7frooBKEBHwkwuMO87eLXx38N0PaTYI4rM4iCWKJlIAK2ylT5Fz/rwybTGy4
7x8/1FxSY1txjcNj0UGf0ZaulwBCclIxSYf6RqDLwv5CQAtX+mFoMPEVSn5YZ0WV
M01xqgSxwQr5c8gmvTKxg0RMkSt3FiAYH9g+JMjT30XcLwVKJrul1av1nsAeUErB
diqBwlBL1FMTtBmxS+KsJf54sXAg4K+b51nTpwFe1a58jskwlfyH+xFtzoKSuQNz
oWBZxTLuMlfftqgA4XJp1J0TNZg0iWfXM+VEM7F/GZz96KuWB+GKA1n55CqC51aD
bIuN6uu7i2cFjdiKYQhWk3fFroKVVijmrmg9oHCYDBfL3mFwwA2eJGZ834bs/Ftx
HIYgcHqVCZxcCfsfAyuMm/M985baykxAvQ7nXExPSWeXd0pq0IXSq/zAP+pOj/vx
bg/pMvUsVw5m4WlPMJ4FUB8nA6T2jQeIjzpr+7C8fnCefxNRHIs7yOooh4riQPiF
4KC+RUF2oVEhC/LyhSpp4BoQmDsci1csoEtYagMe3c0Qjr6yI2mcRPR8nofxxJaV
9M6o4GOGlfmcChTGnhiL5TFGuba3F9shPg4WkZ7onsraepIwg0NPbGqDrg5CaXnT
ywLkaPo8JVTGShBJggu1rVCdwXztyv5fvw8GzszwphRYbfg5V1fCZN9c5T9Cm7bV
S+k0c7VyOF5g3RK0U+5zDUL+yRIclud9/JLN/yH7FBbIBB7j0MV19XvuBxfSJFiD
QREC89yJ9y9BjCbQJTAilCEWxMgwYu65EBoByPUDU4L7YX4PKzhkEPKV2NfewKfe
OHFUJWN/vasElMeX7/c6sW4M9llHRgR9DsHBsfF8GdT5qGc3PtiLfY5n6M0gTDl2
Blz/czgRsS8V5+StxDG2IhGy6nlXufh8aTOcMKz5kl1u1SlTMghM8JUg7e+vNWCf
TvgVWRlBP0pFf4aHYR2Fdpnq80rRoRWM7drGWUzhZFpxgw9xprdtZYcym1JMCt5a
7udiepIzqjeRDE8Ul0V4EZIYl+j18niiic6DauwjVWuEf3KhXvy1/0vCFwtSPnGH
7x04zJAkhAWlpamcOC/ssMvCCf1Xye36ek3ppsB12ijAt1twDvk74Zz8KnjmAj+w
SdWxrbkbnN/Hi9SDzGyb5bSlMRNUDnZforIHM+b7lQrIqswxi0mLzhZIBYiXMwGk
AHUFCCAp+1RuWkZcze1egDUVXKwOfYfVpMhxEihmHaDFjjfkKpB/LgAbrHtoJ1ae
sFBqLODlKctp1PGHnhhv9x+4iJO6ewZ7MjDUDc7nD7rKOtvU6wkkkoe+o/rQR7qF
IbKvKFw4HM1mCwCS9T3GFuHTWuMEYgd/Hn9GUwlB6xgpwCCFDdhHYj7CvBul1DC1
2k8U8wOaXo/ux8ZGtmGKybiw7jdkVxDqcbKCf/R7coKlASGdvHLPV/hQMv2w31NL
HwJrdJwHK4bbLruT6edbHqRFko93JBwLIqvHeynXQHqVLj1Y3hsjI0gl2ISIE7g1
Rgz98l/WYumS1c+yv/NzQw8xnBcu1Oz2dBmoI7xvSroPQPU23aGVxzHWfr/HWeCR
Bri69MexBsj1Sxb1eBYO+kHCyDfj/h0RZ6fPiMuWzQksgN3r1BJqRDo37Ysx3y7A
VvQoAkyf71aKdlm1RkH4rpe9k1CkwjimhcLVTargUrJCWtqXu0lPHl/x2q3l9O5M
tpvorD1FrPQJV8E6K8YNpIEeqXrfWTZHkwTBNbxp0mCveQ1XqCScRiBHJbNmnD0q
SRyy9HTcOcfvktpaNVlom7zYlDZga8Z+8Lj0MRiM8gE43e6CrTM+29gQ07+gD/IE
orgW4EoDT4SMWly5fTR0FTBnb52wWcPCGKdyfLSBYr8/r9aE7kpqBp/G77PjnNYy
8vRHtXjEArnEhLUWxLn4WrcY0XKDKm3lzGXamGfrZyxWStl9/ambPWyIjZyzbxtk
4GFhqc5DxNkl/ZJ7vYDxFJfbbHgn0qkwOodwi2PIBAjV5vPREkFVN50YVLP3ZuY2
4scfQYZvDNENMpoqO6cJLmA5bQZzAdBmIjuLxu73iYQ3GGTEArwNGx1lIRRZ2LRA
jQnbsGs8l3fLgzVQeDQy2r2qmEsgc1+t1y9fhrdf2ccg6f3YBs8BCqeyvigMP/+n
8trf0nxPuEqNDjmtH/1SLLvgTtU0e95CW2F7QpFmHosPdoK4IoH4L4RPIdHiPKTY
dzVco93sjtX3YRU6t1uFJlW0ivAPh/DdIJA1ipNO6ifnSNfgveMPCD0kXfRCZ7TP
yrzH/Ox57T4J7gAgGBoQhxllUMx/VtlT68wRD++FmEK62l3Rdevh0ygC3XUmSI+6
iIbhhYDLKybkoKZYChEadkNjoPuYVKL+93f/vHOZfWRQ1wIljCNl719s8wzf/eWi
eQaAdcovRADVLi0RE2/kj0HlLGuJqJ0jJv2lQZvmB+6eokId7PylPLo0SSUKms9h
iUzJsWfbq2R3RzrNM+7y0FiZ1D7hS+gvZ9RNqHRhcb8eJoDu1iab2NhKRmCN4/2L
0L9QkfNT7jdhCXQJRCr6ZgZZgOvfWqMcY+E6tfgn6nON2lFo2vkmYcmwFPYj4egB
TwJTJQnibuTYHAqbACzHYiTQdtYvMT3an1gXeUUSHB9y1XuBYF1uDu/flE0qvqLB
pzUMah69uVOCGeHyn0RJfObQm5e0RshORqtbViHop2olyuQJpOuQOUccwSjj2wro
i/RxwayNCkGJyxJ2mhrv78/y14doBxeyYey0ULf8UTEnyAOSUojaqgdzHNZrUSSQ
I/xKG5mx1NjzM8BykH0CgTc5oKTuFLYxGEIxO8InZeI6Prud8FZ+bHCptYeja9Th
4wZWEU1trayxitQos/fldugdu9brmSPbcshi1HkOzVJoRmCcSjfQYuOeiDCoFg2K
BVcc5DFmspaBQXsOcqmHLbd8nNjCiyM8ubVzsgrPwAQHGmxOd3gKX2oDcy4VM3CQ
WkGuASysWOR6iuwmi0xSYRHL+n7u+nBXzmb+Ci4z7lv3CFXtyhHBlRSobNrZGt+n
m5YbVyUpaNCVD7avk4ogjAAAGBSMlVyvkOaYNVsx5rns/EElrLqq3FsxtnnpcwrS
g9v9UHfvsSersnwv8WBxYYJcDrMKAGIperwE53C/S4LjI+tWUSOE7A5vEDYWXSPP
qUx4fVSbQln8qASJtKPqxg/lMwygvDn7b6ARYOgKBf8X24PgmJN21TuzSkZcYU73
X8Ytb0Up04UlD4/YdszmAFrLJo/Zki7xI/TSrONG/r8ewDjmrKukUg6CbbQgG/Rq
80Y8EAuKHCuM09onR/Y+NXFQMNk35Mte+nlOXpR6k7/LyA98nmip5SBorQWpwubJ
vSVw8bohCsV8aviukLhY828OZWVl2Jzjk5/ThBdXmisXdw/PzSP/kqvTNEVQub4K
NlHbRql3yJRTCh4r+McQ4HoeDSyEV3MVuDmOMEDKm9U588CKHqSmfm63epLoyG/P
FMBFreQo8IG5X2GjE/1JaAc2VLz16flYx79COeKjg6mHtPT5X6kipXSVSpohCIbj
4IGhTDBApl8v9+5wmi5pGBr0l5jqN/YLdQxns6fM7r0y+rqHUc6d1akpu18/CRfk
R+wRmdX1L2jbOCwQG+s26dRMYUZkHWcqffEtee2sQ5QLHTIx+64qqc9SuCsZWTVn
NGN+bo6h4XSBctlQIJ95Y/rwYnVIkXRuWxnoyLxEuC8Ci/qvmq772XaImOJyW/3e
1MYdaWkDrcat9rc1pQbxuayU7iWXZG+yVS7hzX8quIcXSIGgbJbDy8WwHCkQRmD1
mvmA4s8caIusmnTJfj3SRiRpQSk6a/zfVYspEvTou464ieh9BKhWgPLnEoVdT2bV
SbdbCUJ7YnGw0HfyaHlMuWjS7K2KiXiWYO0BFwUx4f1sFgrvP64U2x10QwpYWH2/
6JjC+IQYTl/Onwxrwn9oJV5zo0bbGVmu7dOUQSL60gWDZgVVPyFSoJo0+qW8LmL7
Q641zc+Ukec75LmzX7PCzjZaw8Zp/3YnGcxuNkNKiSuOXxPoFJ7UWobYJ9IfwJwe
+Wk+q+e6XoSJfJbbvoOaS+xmkyzVJNYjwUsNltX1dORBlKfr53PTczANbOJAuf7e
EJBrObEOjihSgBLyFeRUwyzrDgygdGPiY4PYVgm827M3DAgdB1xiLuGjzgtTpVw6
YiQ2eLv84TpQ4zj/RNrsODwRLjLi4PRxrP1OGb60GgI1SVM5It6dTJpDNo+Npq6Y
tj0YghuJAhBzycR1Bcw9chZdx9/Jh5i/AuC/ypAkUhZKQwxPXQ5HjXVD5efKKUwH
d1W2T04qUR+TIYIlFEmS7+ktB8VJ8mW6vUnTnJgTn82Ih/kOy2XKDA74CJTX7kZq
hDoKG7p08QR0SQe9v9jk3Wj1+pE2ZKh+2dxM7XD5/TVjiCX4p779ajrV+UaZpkdx
LbaQ6eubxLXu88usMcttC8M29FIOWWpn93nc5BQVAjiVCKw57rJVhgBY/i9tm3A2
UsH8zWZ4PavprgDE8h/C8BNAi6rvWAJJ8uRREAZZ1zj0qs1NX46ViXyfUELEd8Jy
xs+PcVMXxGzn1qhPnAOc1KVqgxx7iaKsRQZwpzaAjKnNVwYvfowDjMuucr7knNCq
CXOkNTkPiSdmEZ0oxmMk/3krSc63JPPq0GtFUXFiphgfDKUt9qHnIpxAaNvsRvdj
6TlORmZ4Gd7SaiGLohkX6YGtRlDtmgb8LdMpTSqHtgZcFQTBLQ/Xb3VwddVhT65h
3kzC4s06e48mpnk6XSaL+jaHGXTwHPIFx+Gq29rFSTzT/nGClkFsSfO820iPr23V
lGlS6rNJKWTu0JcIxuPMYuB4tzmcj/Xm3SE3inASx5itTD0Jo+6x+1Ii0Q19uRWp
j/7RQDIefONv4PbRz2Q+jgEstxrkVZRE6oeeRmWBcU0mQEwKItVthI2q4J0Mr1r+
NLusujZD6qWUc/yeZyILnRt1Ut1I22+mo2XKXv8+ZPrywHSCNhxn6sTnGTI4kvaX
kIE8aIfuin/GitcvbklGpN91pCyfRhhJCq7uD93IuDQ44kaoK2Yo3Uu7TLZzal8V
lSP4JEqh6l/kS2kDrziIVh40V3oXV1sUYUklyyUEDvTVzB5JvCbEbyHunGcSs8Df
nc6IM2SHgmJk7tlbv+lsPZ1hjzxtDd+isLc7RwBok/TF4OssKR1dVQI7qQab8y4x
7QaagiYUuyBaCFkotg16sLwxoEoghC+F6Fwt1sdgRFzx8jrod6d/3A1kcjBWWm/T
bDkMxmLHJNwh/AJdXLMaPpWnvfHYnapTCYl04pRSPur39Ae1ccLQK8Wfkasb77ui
qMpjPC0Ph59JoB+bFzNHQnyPZ85ZwTjWxgcjfBsd4d+jpsozKyJxZ7Y1Sel3abw6
x8Ft27yr8LVtII7abRQfANn6rUYmFKAG30WYKbOOsH3h3eF7FPKHqPKjUXI+9/gp
pavBQi4OybDtgLLlu08iT/Wwmpj5zAHUdpP0SKDik+pdSg9N1PasMXFITTz4tEMd
RggqKpOe/s0TFwYhXOFyIQIf4waOQ9UIAO4iKT/9+eqE3hdfSnIa9fj/Z7R+QBAg
2vUIh5/Ewzso9UPHjaHiShuTMbXyjGbQTZ3Cvlz5zK5prVlj6OEgLWz4PQOVjdtG
6gxY7iljgCerTsov7ZSK9DITDgyU4BmYT2+oL8JcNT5whz0qLY7Ot3j48/iIXrcg
Etx4vpitoIDTvYE/NNf3CZle7zO7Oz5iDLXIOxjVKDUERJXBq6tQpQUmIcX4ar5q
3JzPpFmMPkm+Y33oo8eMBhm6iweFnwa2pQyeYrninNiEItGsAYpfOP6dWWP0L8OU
JCpNCw5Br4boVTDpZiWYf86Tqgrr45kY2C+B1VSIDr2xjpsz8E/jZTsurG6pCUjz
5ifl5uvk9Anrj4fjImqQfNu3kqbjkpeoYxgj73uW0sENVyG+GIO4oz3byWDiBqsx
hdIgWPgoM9qfA+KY7VyjadB35AIcF97JZU95nXhA9GKpGouAjOtvhKKkPTY+hiUy
vQoMHHRytlFPROnredxeGR2rls0EgJ58u/od/O8SCJVMa8kNJig8VC2YSUXXrEzn
EXHAqFgQBwCnF+gYbMPrgDVjFEBL3MjKBNBifUzh0nb+JQ+PkKQa05gA4S6dKKMW
Nc9HB0m/77IOIC+jQl43G/mPw9KoFOHlHLGIDlpPNaHpNvz46J8ivDJdENtuWYph
S12N9I8erdDteabWEOkIi2+udWeFYp2UPRsBzj5v0rMkZt9EQWX5ZyWx87S7bVDd
8LhKoDp+Q5aJy/H60CFUhNe9eM8TJe8Qko5vq5rOxYKRmrPF2QQ5HhtbFb6al3ZY
PT+9bNLNVV6azlXvfW21cL/4swCFsqq0q4J7rDFjqAev0Ldfssav8Wx7YKAPdF+x
GF9sDOQMVFNsyNiOjQjVloee/DzSusa++fMdtoU4p6RT5jI7eXHRRdm/wI866Ipc
RvWgdFCpFEHesxqas0HH8DAdkNkGqlQ1xOwyJfH2DqnY5X+3jk2CKMbV3V0tnLSz
+Sz9pqD95oFk2Td1TuBbxqe9y8oXxHev7/H133q9CrG0jGABAz8/ldKxcNECOJYK
LrrVbSFITPunVBkAHLx8Q5nPaYz5g+y3MNln+/yYMGHKnM/rWgMWvwx8ariQQMXG
4c2ixxrgLkqDrUbuWBrX+bKaOUaGzjcMB21YJyVAfnpr9AOOK/Mnaz4a5/9hOIgb
Zb8f7x+9crCkuYnViBt90de1AU5BGLjOh9FFxBZauvp5RpNgpsaOUm34imbBgiB4
yp0d0jS+5peb6S1EcuIhcHd//82nP9Tx2cnAn0b6nYnDoTySnqkioaGBgYuqzpDL
4l0D26R8GTlrmxGIfIkG1+69e7GOlr8/4xnZ8BtEwuVzb8NnSvnSF7fu2m9I8JqT
Wwc5V0e6VmDfZEiZRVoBkTFElOiwHUZMX7QCmlR5l7prYzdI/LJpjIP0thZ6Rx4F
XOwWhMQHGjhEJgUJWDFMxXks2p2xSuVblFmMAQ+zScNSh3TOIwl3OMBUr5K+uxsL
u+FLh9e8UglchldZcPmOadkDm2cW+lCunq9qOPp5v9itF1f/0tuyzrJ3uMz5V54/
LA7SIJxaAoJkdMjd8uRAEsU1KcGfW1qk0g3VLDrKfr1sD9RTtAfW2h5E52WuVxYY
Mvph2bVxN/ueP7R45dAAoM3G6TVS1Rs49S3n8QmNWRVh1WU2ZkI1hPg9m6Ch9dAw
6tno/nqABkIhPi/UY8D98RFeZ2KC0Z9N+tLEGL/QGAxMwAAhYDRoJ0lDDZQ6ELFT
UAjdCU/7zg+1vf1TA2tQTA31z7toXAfc/sgHq4U8o+MhRCHGE/aMxCtzBkMCZw+D
Q+1H5Wtx05+Z8PK/OS/ayRpPw1EN8Qx8m6WZoDwoxzXOvGtbdhsRymJm0nZUFjnT
uNDJUOv9+J7I8oVrIeDZd9lv1z5PZgnvbTC+pr5ucqoAbH9GTOE/4qzOCAjq2wsB
N0CS8oFt6Gly67/Iuu3On9OcGJxL1vx+wjr4n4KF2oF74TuXFpE/v3D6Iubhiq+v
xihSAol1WQQWm/JZ+jPgB3AzXcQMKmFGR+tqKsBOgdmv1aC81zGhkJN4P3sU6pCA
VefX5Soo2oIYM8OP1rF7wRG/cFZsVrXxPfqCWMVnuVSv2Os56VUbH1Ck5YH5gQSP
npGZJS3oLJVl01tUvlZZh3ZMwyjosnzJGxkg8Nmi2vxp4Lcxga4IiZURuANO1zLY
GYiA0V307286LRp5QWNNJiOmb+PKYfGld0Qd/LeEXb4i8kP6PFVmiepyvpDw1YSp
28jP/ahGNbVgdBtVZdXngRgwHc3N4B4TqgMmrBgWnGBmpFyvh524pZz0z54JzDOl
TzbDgAiHwZZjMMXTgzjhuOnCBEWnBMjapFqs9HYxzg13byfeZdldfs0dtVietAtY
P8pjLzV0CtOJJKoWH/hBEMGE/rxEZPJU3Oc/xLNRz5H3uwh3Mz54OntRwZLmTQXo
/7CnhvzvmjGIvQGQV5onjgrjlnuzsxuTuGi9GfsSyKNw8UemH2r4Ax0QprMdWTcA
pqn6yttkFfLJ4bIHVjlUcncngdUOcUWiKmSj6WnlJ3+rTIzLe8IHJrMfcnP43QK8
munnVXjPGFZuwuKZI5UzbPqG9poHWM0AOk3io82E6Y7xz2jZHD3x7VSQ5zsevNix
ZDHhKlR5HwnVZSwH9fXbehSaa9A1SHdWnluUT1qei0O1wenXKzweIMX7Fuk83xTM
ZmaFhJCAfwjup7gZEzSx+k+TKUPvCUZetKdmus6xk0ftnTpX7NHjsD2Y9LjXT2nn
uQJNj71gKxKASzn5u0V88T0doHr//GA1/B6HhgDPsBF5YuMNlo23oX3OJz46oyFW
5X935kYVp/y05WBB+YfFbiFdDs7oaXiJL2vVJkxef5BAmhv2qc4UIsXonocsk+l8
xpqmHWWzT7MeTBTx+Bn9yQhssf4tAqDVY6RQChQe5UPiT0VphE3u47rcVmUcjqrj
nNyhaoWF1sT/Q3DfW7HIxnFzQ01EG5IDaQpxaNlhhbIhLSsTc20j6MhTwptkugNI
q/gAM8dESaS0Eu/4MguXoSfKHdg9zRoNjpzHrPNZ9lrZem4PZrHFbLWWduXI4gqS
zNsgQP6Ovjf+41frdfjXOe4y7s+QJ6ltL6pjA8RGJK2Z9HBm/iNSXSPPj7aeObQK
F8/Rdwmtct4sTATj/6WjRY3N84TecvED0GnJmQpg9i9ZTCkYRTmPn5vxxb+34zvr
BeYPTU56uL1FIWdAILJIZIfKlpJqz/Dg+z0agkZPCQ40iHXhsnz+wGOxc75MbR9Q
5ckyi9cjmBGObi9m3nHqTKCgzNA4W0/zh+FSSgxxtPVBitp7Su5eJgbC74Bj9YcU
c9XXtCkZWNAD1v28Kd8lsiXcqLBVABWKOcfCHb1HGEUaK1l1QM3qmc6TXVijkZP6
bcU5UnShbx7Yi5TYCTK9KKVguXwSxWex7ZAjJwZzFIHl+Ss7zixLzwiREG+T1vPt
zOu5tN9Q0csELS2xW9JAWE5s/mpbQvWj4QCF/Q9/ZdRCjS5n6krmbLj+uJG/LTzf
QNfsF4vGVP1IVxL3VAA+FPfyDrafK2kJLUPy8QPpqs7VbTtKgly+GPLpjm66mYS3
vttt0BBPIAlnM7sEn8GbJrQegOnszUkBlvPpVsiMw1V76JnuyAPAWpRFh+/Ro8wU
HzbJofKGJWVTa5nF0pEHTlGxxGvbO3g5GpCPmvuzp2w0nX4jv/KXtZHpBEz8VVDH
TKpKZlQpEtBVby0hD4LLj0WlwOJm5oSoGpAe2CBJizGSkrsuh4FQZsssuy08/3Mw
ffNUYViPGK1lHh9RRwrq/BkB4kF69dJdhUbgmKbUCk89+g53u8qyi9t8KM/rAKP2
F2lkGK1ImEXYFsRljiiWCQOre+z6+35iG78xJmv1Umq0jebPMk3GWxdNHL9TvL5n
+gV4AuQFvFh/phmuSbLmrZ4seADYfLFMTA+kv4Zw6zhjQ/e7pzNgJbpRTlgUMiGA
fv+ALf0dBtaqyWtCmlDzwIaRYdZXPN2iGu0wLuMzKEvC69XCHDbcE7H8xIyNeT9e
/zYCCVrbZSoa+OcCvuEgbkOiv0Ch2FLKqoIyw2th8NGh5qRcTx2MEQTm/wUMAPZ9
TljOZXciJypZ9pardPz1Y8It9yd+oGQY9d3Lv9t1lM2h8zb8Tq7jDxfVEImWB0Od
qB1DtTNlkVPM0VWRSZCgIno3MO2FStF4ZhweBgu7hrLeRdm7U/2tlydrlxHJBgnQ
S1et0clgWrJuLHeXbqj6iY0qigICSGry6+x2vLUN/5kUbFSdBieSwMFTB5DCIQsb
S2cdLydQxbqoY4IqoKMbt7CHn9FiJ6IYveX4ClwbFrbZ1DHC1IjZGf/H71+YO8tE
in4bG8gwM5O3N/b6BcAzbA3y0g4IL+PY09Db+sfRzGdLPQcH12vi1ILXj+OeR8fT
wW0ZBcPmtdHX27e17E0XwzqyEm7FlECc6eA5TukMbmj1y1tWLjmdi/1g5mFTe6C3
Lm6qDkItPtMhW7lAluuPVTWW0hHAsJJZsHEW9QJJAuRCKIufqxcV62WGkuZzJyhC
8HgBcja9AsbAom64JkeGB1fXRowg02tvoKE4FD5PBqFdiwXkjY5SvFS/2WuRX/C+
oOQ0y08elG25yMcLkUa313hiLnGkd8ufmOXasZTiq4VvFLFGKYfnyOn5N9p+S++k
da3Ro+w1PftGW+p6jxOPkJ5mTufe9bY3PCqgw1LAeZAzDGGEdOJm/uqoYvEEZYzE
fw+FIo7A1gD3xuozoB6hZT7cU6iLBAzDW3f/Atxdf1iFUT4vG1d/1I8Y+NG4H2Oh
YnR1uOkRBRiUP+X+cb9+51qEN31+v0oX8v4TAhGZQK6aIeyl2OfWdnWIlYflwtn5
3fcd8XwUEtHVVtO5rWDDJUm9Brp6Rsl9mFL190DGpsKvC1TUj6KMhS52DyilyghM
0OEUHCNcbYCwm0gsRoQklX+H2ZiMXTEV88o/AiO8aPwSrO3ROKMsrgGaMykvamUq
cBvlQ3ERhAqC6+nSyvNYBSryFFbvZIxc90xoUw/oOnsF1d0cASq///CsSi12lATv
oXxnFqTLlbUSgbffJQheV7yWhgk1ug2tWyTxc/g2DA6gWPvQHcLRW0KTX7/ti9OZ
hiutwOxOJNZvzm/v1PPyhSMvD5RQw4F1/9tKYn2X7m73L/AD6G6rWLAd3fp4HTMX
0tvTf3L0hDJOaldmp3dgEVqP88QCg/18XSxetuOuuHOL4SvPtsLuPy+ct6SJ737f
OS8PJCFbPFecdHkJbcfmogIR7uACE6GhcuXG7YD+ms7CzINMv0LR01deix+FGpV1
W73I6IHJ8RLvm+KaYhsU+43yhLlp/qYfNfNw5SyjFzlezcX1U5zXgdyTPeb86koN
+E7wV3+MCDeVmEtcvMTupwD72STnFXWVh5PhLjnLrraeNBCQ+cs+BVfZk6CH4S7z
kzXeuamjShzIabh8hz/djnky3+KZ4c5mwz2cFFM8WYFLgUFDIJGjd14AbunVkZss
cZjMNuQFdeevYZSNjtwHtj10tUnwgsIBg+zVRM1E+46dt2m6MW7NT5KZL2xXSxLe
/4a4VmQAwxHib/fILg2O/eK04fH1ah5mtfHAr48PiqbZorgdq/4kWWvRi59DAruW
8kWAhl9GC2rronIizgd6NWp/i9BnFTE0AX02e9OwybmbSel6lQlwKCEDnudBpVVF
34QasgeSkZaC+9UGv9DNqchkOT96W6WioQim0MMv2awk/ESQsxw8XesScnYEnyjl
ML2IzJj1tfuIkCWqppIu5SCVJXew9Kcsi88885ODo0hKdVokS4GU5d6snHyPEFxq
tvcAajVeIk4RJ1h4+bVxk4yaXMh3iLHq6UeM/tWNnJbmEPsoqLpp+vauLequgL2l
V1qMUcNlGREqRhoOV0DR0v4bVH+4JC+tfnSY3PS2cEyvfmpf1OO9oJ71SOnEke0A
IY50sV/a5Y7EyrzP3L1pSHCywmIaUd+A0b5te/JCRjAreByPpyCI3Je4zTP7onl8
yd5690//jKNMejyVNvlUUC2n1TMeqVqE2LR6/7m5TfZY97SarAXhx00l/gWmcBXO
Gbmk/8zZMOmA8QboP717q+6wTyAH3hy2DO7PGzie3J7TSN4dHAfvanE0Tlql8kXE
ZNX0aCcMt1WNeGS0eI0ieWTlnGRn9L7EuykD/BmW2iDv6NYrfVCLNQQbtgcHxYOy
tEu858yLZrVDbPzCT+il4oIVBWjS1+gTat8yNP6JSLv9iMFvxoNXQZujJJ84/CM4
EY3XrjD1hFfhl4iJo65oTBF2N3Lkb0rkUUPEJw0+vE3chl0BjThPQv24pxIsCfRp
//SjEKVltV6ihJzF8BNsMficNz5NKR1y/VC2fMovVgL+wcKAPDRtt7l0DuGs513c
f8RLHwjYZHZh5X6Rpo0F/oQeUDgjjJ5ue8Ct8V2HrBhhE96O39IbNrdgcIrj4VMC
if6blXHmM7LUqfDPG1OxqaNyjqAG66v+0Ng7bdVMeVTRh8ljlHJAaoP273eK3LQ0
PnE36WSC/NxhXPWLY2izLm5hcxWax/FtTuyRPWSTXuXxx3xKBz9yvwm7azAuImSG
KNIkrY17KBkmgCJEBch+cr47jymu71lhsl+iwULXa/w37HgRjJcPmAP1nwTiuMP8
sLfJODYiKZz2yo9ih6GNpOSOqzdNfZtp+JvhTK+1n852+1yGWff35CT3saK+0wED
YLuflelELrKky+qf2qDwu9KIAJFqPKH9oeQIuY/VMKz/yGaqKdctu7MVZcvGnYcT
kLI1DxbGqqsqh0llciSQz7AZpyReBXH6z8HCcACoONk6PFBDpDhJky8Afu+nlt0B
jHMNMhPYEPk6uDWUM1p4WC1RNXjThJMTfStTY4Z8viZNbHZnbyAz2hS7oi9CBi7y
1zRCnyl/LhNgOodEfh6c70LqEvIudoEw3O8HG4Vrsp/PxNbSs5akHv5+rDRvIXZl
DT9Lvuu739OibNF4vPsrUriDgv+kwYWAWaPYrTDtLyohF+YLyiFGXppKK66TEqsB
twRhgWmDwf7zJtHTJQnMIDFgpCbrxCDYkFM4CTSOgxB35SrUBr7ViEa56fZaETTU
SstOXb5DcRV0/6Tk3YNlKOnZ173l/4x//qWDAWMFgqRMKpIpXFPQUTrmBtsQ3kKt
w0JZskwlj6C/ywLlMKcSN0xEm2mg41FFbjdOJi1OO5gCNki0ZLx185VfJXfiLZYH
u5V/ChJo4l7uH6bqieBVANgRn/E6AIyyC0LWKlNTJw74hQ+Ogt1WgZSVGQjaDkO4
cYBTx9EPhEE99ON1p1rq8+3Cp7IRx8Y47d3cgWGgj4q326UYfYUK7UbAHkvrI4S6
Hm5stUKlvXrf5IBjfLOkvKqaVAtJRZ9BEEhFCxLTi5HFccnb3uKtkW/IPRFgijC0
9ZVt3nEQfkuFntxUk2TC8bLUJAtdBjq8tmWBh35GHoOMRFxPpf1z2mQQHOjfQR+N
Kn+zSY2nPnXjXl1XmhN9FrneweJRiwPjTKfkTkWbcR2UI5djjy3zm0V8Wj7+vUSR
spPIkdT54LUJuVI6HQqmIZEohlqYCAEWR1iMkFPrOAvSNpjNlKdcrue17BHTRGS8
jEny9AKRK+H64NxbCBu+DZxPDvZHolH7i1/by1vUmDGl7f4bCCjoqs9OQDrVfTaz
t5m3Jgu8mbME+LTOawTkOlsS7JJGbSMSZ2eyKxuxwOYYx/B+HrGzMLKteKe+xFiU
X3AYceXeLc9MAjGs58ZnuIhebNoyKHXNe1719qFdclveTaEV1/+0yLJGQsmw+m3S
XkLurRVx1YmzjhjT35sTaBCwdMtYlH14ecajNNDwILwLO3OMf5idIFmBN6g3Etlh
Fr0q/dZisE6bi+mScs6tXBVIFx/HYsg07dR/mfGs2Cr5f5Gtcb2A0uic+MbWiT0c
rHCsue9JiPhPwnMePzkJ/xYysV2SnV3kS1idKv5+iAD92SKsCqbd25N4jGMX3ivO
JA82qJskrHuJyjW/ISkksi1Cw5PcYWRvndeRwCaPo4MEGSQOdvgGe25Aj2/rK0m1
gBdsOroWsfC3NCH4+erpvFDjD7kJH+de1iz50BIdFGtXURihTk8sDR+Qyy6Jwh5k
hHFBHcAum3HehY5DA4VAqfftOoDNxlcQ3VZVsYWxT7HMxzvYRPoFRn5OZH69l90S
V27pV32NWGeGqD1DGxWUbOvHgpvnMVkMRlaUDqtnE+IK2ZUZmdsOdT1hIU2eIjl5
81oRaa3Er3S54w0Cr0/yqZNPhJHsLYGe361HepHfgQVgJBOfAbNjJMSLlH0Uq70R
TOtm5VOags6p1GvE1kMM/AdbtLjk28bF1YNL+EpXj93EfoKZOghToYBZ5b9J/US6
QQ+kexeGynAreSzjg+jRcG+s4ahyDk70rM40ibj0bivGGb8TO2OProrhkILuFJSK
NPhDZ8APxPXB1/vnctRMG2GMvexCg8a/Hq6vz4xcpgghYLadqrFePjcG5jenM1eI
sTkOpHOiH3j438KySiuLVT+drXgOQiDQ0mYCRUEplRjvBMYUvzEBzXJJQyEw4tRc
8v+H4QS8A2LCgcE9AJAlQWfZwQ8xO/e7OEq8lWpG4YBrfjJ1vTnR5DbXqDyUWl30
rRJFmeQp1Ioj19kfnp14bItDmnDr8xH9m5W+7NNDJM4FkBApXWoewxpoliomMd1v
ikIc2S5vaGS35ekp7VVzwdsETr1IhK32nHVRbxEQivhWPxUtp+KHkylHn9nxGP7/
EWvEKOI+FcW9UBMGHsMQi5tgca1rN9sP6Q25nrmBNndgX/akZzoez0yI2s3REbIP
fyq5KkE+RgZR0mBj7mukA9uRo5eOkOp10JM8ZF6/+/XmWhlMj3WY6S39E7nxGQWn
ACj+fpzQhFezTm7yLSztcz2MB942flMH0jg/nmx1/D8qvkxn6Z+/TuiBWW/Q8ftd
4CvSWPwGyoSD/aBI8KsTXaQdln14XhUGzXvsO1V5qHD9EH0fWg9oDM5K9jNMERPy
63nuM8BJUIYKvWFRkQluNfd6BMYAHdNTrghDe1gWo92d/v0U1KdeB5kLkz8AuzIU
37tlIMp2WXDgeo4KNvry+Z2v8g74NLGuJXtBm+VL6weB8kyWnBw5AoXdH2ZIIdFK
q4lti3GI5Hn1WolAcQpeS+3GpB23NOiwaR6XLK9mwekCKOWSUITkamP9njpjCXHZ
3ytkEDyt/8YYPGsUtJnvbaQ15yzbHiYBaGHmrZ2TrGB11zPOUH9OrhYQCQlzd40h
FR+9okfol6se5klK7p5vZsX7arcBSHgdX1FB2tXyfu/wc20IWXmwzWjCwgTnBZxI
joVRLRQP2fNc3FecvunrFnrmWiMx5GW+w9ukJBv0gxzO5kR+LfIyj3IaXrBJ2FnY
sE/ixxRsOgOUGiGbJLsN7v5YLAYuPEZO33WJQEgfbJF7UYHn0cvRMABoRJokE0af
YtCEGuSGUSjno0o5nT2EiOPxU+w2v/gBx7bKUniB3q0pZCV9RadnioQIu9ueWQrR
JinL7rtzCuWsUhjsUJQC8dQuA5hxYs1hQcnx/b8xJNeFoBWGRnaLj6Hcp8a8b0Vc
BFhQ0izE7SSiYr3ugQBg7BFYGYYTREvseGmSr6aYhnlDP3tfbKoXN732c6OzWXeQ
BAjwTpfwQMpeHU0lWV5IPxDpBENpEAKApu4HVabw1tY3MCG7VFhxTwTL5Zb+8AAi
18aSyB3TN0NtHoO5Itlj9YDpqE0Bqp1DZiUgyntZbWlB1OcsSBaP6E7veqmdyM6+
Pg9l+Mvl2o3pyHpY2y7xndjBDa9esxeAMJlujAHKvYV1boC4ZXBMkhl+DSBfjl2q
J8cgW1Cb0SXfoJXiC43ZBG2KtQYct49aG1xtFmLwkW13Q7Vo2Hfjpk7yD6AV8IV0
DPQkCVnaSEGXIGDewbvBda0OFglqEXnnImqGToECEVECMZ9SuAGEe7EgR6oHGW5A
v77axot80cDZUj/mGRD4/cJgregPWGOi1XoXgkeP8BjSKp/3SKetGiqZl4iD4ExA
MHmo/q6ESzAsnSIBrpe8f9O5E9lcmXqInKrbJwTX0MpdnD2H1vEq4xU7TJhvueZ4
klqQ+8nBqiKV9cPCufGZ00eW9BhdnTI6H20/962rvXIoyzkk/S1eLKz0+IRwUcao
0H3WchhD008G0wG7VVOU/Vdg8poGnMvOHW7z9DwwWT46l+M/dfOnIrUOhB60mjvw
60QncyLpFrVSXpO52FLmYULLdsIkp76/7LaLs00SteHu3GvhWsb+dzlJu0D2Gmaj
s+/DamZ+9e9KOtb9Qm3cESKlSUIIjWNDvUHzusR4hpyiKQGwdZHGLXKOAfUTkIa5
UrfM+0LqGj53tMN540sdW+JPq9IMVMO/PLrbHfm9YhmrLsU8AKBJZL57urGDHSwb
qaE4wFJm1mmSHB85znBASt1jmiQYdEal5Tlkp1nJbRRslRpvQ/RzsnlifVzG7Bhw
N4yjRQcw+hhqp9jk5T1FhPEciIhga5Zrl0hpi6knHIQgfPl1VpsB1wYa/Sw27Fms
dZmEtEo2Jnbf7EtPXNmq9x+hYBw5/Vzeuk8Fj9irqTCNaLf78tk8zu32Mh3ahgHa
PFgToZQAainRi6xsoKMRsvGJLn+dzyHj+QTxWyu8gBK1CT55UO3WWofRpV3AuEe0
t8MJvURr4LmK1rbqQ1q8BqPJlFSl4M9S0ZDXuswv5PyxN/m/GqobmYzkvYXnjVmm
1CF4+W+sHTJPHTxLLfyF5Kp4zFu+KeKctdkm5MVNBI5BjOD876VMDQ9wrwSqI6QU
si15PmciJ4If3uiJUYzCvqDAAintBWEtbk5DGIoJeE5Pq5rDluWVrJ7UCc0B0pm4
lOF2XatZMnHk4D6qcp0q03m2qnGPuw0F9EVHXOpuHYUJu7SVegGK24A4Bk85lSBj
jQFkKKdWiadrZ7uXRfNWBvghdI+4SQ0sV0uhbmlsJNAj+eNe1D4lQDeyYlRBE2P+
q9q92OGzY7ueX3Ih92r5W3rBU0nAR/A0ZQyj/tLuOCzsAZMkscFCwqmdA6JeSuz8
R1N23OY9ZzRROdrmkBOhjljW2nYGJQHFRCHM6mnkmGQLnnoZwv3dExQc9t3EX2Fg
QXkPwpNXQZGPZz4RtYjrjNGmvT8VbDVby5tW+UTIWDs5Tgew6YnvgmGctalK1wfR
hXNt+UJri7/8fElMYCwymPf4WHj3+OAhDh0GcBxlBy+Eybl21lSxGkU6MUqlwAah
ODMgufsEEh+m8vy1Di7Bm/EOvAeFbsU6C6f1m/009jGBJLipgUTpnNQ1pYtkyIgO
QsTkXafGyA3ug9PdGK+mQtlAlo50LKBf1UQ7SgGDQQSxYUpYTsRvVQoSUb7J0dVg
6Yi2j5yXj+gVJKxn/WuGg3erq+Sxt7jfkS3SB5rXRkGcFOieaQ/yhW4HLT4H+KYB
034/sw3arfprczaCDZwjhegBTwz7opcsQo2Ayz2mNgNtacvQ9/4LSU50ky7Ul1oH
xWtqQdpTY2Vj9zbD00g0f4MGYmCge75SfoVNc6vBRvtouVLxtXpVx7Xtaf/Tft39
2dyPGKgGOvl0RREwsScNsWc4CYef1oTvylyiRngIWYYQArp8hQYhvpbTSX+X0kaH
zt7T1ZbrWwEOoZWCSUg70wxdN/jYYccUyICV+LVKI651eDOBAuIbmAFfkDT55cmm
H+GXxp2024ZI1s9CFk2/N2gomQdXFm742uaFxaFr8TcecQABo+4G8MXbJActKkrK
8uxUZ8OfP31BN9B4TjVAR+kbmNNDNn98a/5pxgQGYOppoehknZ1Fimr4zDLlYLFe
YoK/IuzPt6owPXEKk9kMDu94PMSh/yqD8nIVCHYgcXQOURn2zAYFOqbiNPSSFTiq
vserc2IJaspw3wYptx/ZJ/YPPymWwu3QzTBqp7kdmGtjZXgBkKvwgmF8bcgOIJfq
scxy5putixbkL3k3PUDVRAik0tW6ZDOiIyv3uoDzFO0OzxHEYl5dPeiale+btb1w
JKgTHLDOZH/Q/BU1ny4/nz3QyEgjlajnPK1I7ia7K/+EIzYLAarFWYlTztWfyVc2
BzZZtbSgYSOdEPLs9npAjMQPH58VMsc0LVUQSkxgC0DRGyTZ9CTc5zjMV2C2/x/M
9FSp6Wkd+sn8fMns3EYxXP+G2qNUk471ZbpyMa2uvBFKE7DdQDPq2VA3vZr4sCeD
bZA15FfIwD46fKobGYUpBUhbckGcOkZB0tt03GA/ZAkVOgfvJfBaMNevRKJIIUBP
auc9vWYPhW5MYd+q6tmGAUHGgfLHS85Sy/TRof9GTqc1yaRCn8JIGogBRMMj7V3Y
HziLeSEhbIY1GsvR/2khtPPljFha62x4lyh7V3aTV+FhknMvbsaZW2kv2PzGqN5O
Gglm+e4gJE2rQKQKRrUVJ2oabmAQ3GSZ9nw0xSV6NM1gekH4voWNM4r13GfYLc3n
Q8EgjKi2V5RvJb5TEBNGLKEAcrXMVn4/T0mOvZreUxs+TFsJgARKxnxcgoRuPB54
S69aDVeGBRX/DRZjMig+G1h+LbwL9xlEfAVTF6jaAOdhXBxhERKsTdkg9vIC51Xs
fkSE129/8g2gHFdiw6BTl3l1E3zRQJYNovtdbNudFvyhfvXfHg7hILfm5XzgphuB
41fzO/DZ3RdJG9lmmhilUc8m2dI6joW4JgM5Pvw+0J0GL0VB/mF5kFKXL3iDQivk
+qR7RigBYTDIh/XpstJJB/lCXHTaSpjfAM8t/QOt+dI7vxWUZzJK9hNXFq96+5xS
KLczNGJ5TIFb7x11LG7RDfEIM0kGrk8zRI8fRvUW4jwBf9oWuCsJto0naIs9p3XH
7jmm24ov6wR+dvJyk6vyp6W3HYwVl2GjS6xSdKHuDBRvA43ssEJpHoxVK1HkHHF/
RynNKP0SNNxi1X0tfE1S6ZUZu97Wa4yNZurYOKcR4s9ShSDk4q8iPRqet3StoxBH
32i8Ut4xCbx9Ho/OaenEtBb8Y1OhWwzH5izZ2oClimcihrSlqCJyVEnbcEy9Fm//
3Fi009aDuEuHNyjthtgtOuaSLWjbYGkmYQ8S8nI8cg8fxaKyqDMFGOKDolQYhZN3
avzZ9WtQUbclMRPLK74uFgQYs99roMZaPohCZ4TObN7dLAkZiUSTR3PQRQ0cwGzY
p/RjZbBmkhn5TqwbQz5qckSOQp7qmOMML5swF7Da0QQY/DQ/skEcQtmNix3WKd48
ayrfRf4hFuJK+yT0Wfgy8CBnkKzpuIu0RxxnrRip670F+I2E0xASlwTHy7S0+opg
NIYjBl1jej//B/W45yb8wokt2lMr9+GIZ8TaMrNuEMSXwjxDxwSbyUIsOQ6JuLxL
feieTXXShNks6l0idFuD7L9eUYPHDDoywHfHH5sDC6+5Sk4wIdKlXxekqzxfiK4U
NftwaL1/MMeu9atiuWdfhIosH/LAP7jwXjseS2uAcc/MhC8OxmtIZSuJDqdII+SV
86Tlq8Fy8wSyZevW0+ei4FFey1WzLP5SmHr1fAd5JD5NYL/YJNGL79FWIxqD3NMg
/Y4e6Frsgy4c1wCUQKZKnP28mHw2oBtVBTXs2YN++VshbS+UN8cfBUgC8b0jFfnn
gDTftjrq03gBe7zaQBWrKHm+NbyA4Bk8gV21X2TZVSBpb4JboAdHKC4uHJ/a62tt
zUS6LN3fwpMgyO1r8ltBLsh6SfDP9DxNogIOf0L8U+NCWj1QA0GUVbTyuIOWU6ib
LHY0UVl8jcAGPa9iwxr2FFbnEXe9zWMiHK9OIdYFoIcYzs/9lb7F9rjjkrckQ5DC
JJAkoo5LCEucRqI1QN64ko9S2N/nXZr9+fabgbbVUoWeYzjmoVXOvZdIPTdTbxL+
MMFOCmmleR5WemAd4QoRFN8DqTpK9pSYPOVOa8v4SGlgU3GZLxM2aZZZJiIJKPOd
ii1TRJNn1PoGgAyn6s94O+qS1HGpTNBUCjx5qoJEv1YYAqT+CtVjxNjyifJX9gR/
PDnWDQutXbkvdY/CZsixMCwYpDPzLMWxffLI0KFzu15R9YaHaMkuhc0lOGPdhMLT
lQ9PZ/Ya1dfucoelXzl+SDjdAYsOcy++Umn+KGh61OgY2WvfyeKyzhePvoVPSP4x
Lq0AQkPboxewcba01iKGRcTu6//aoS/pfLyjoTAtSWsuCibCNPkJ1h2p6vksdkej
agPKjdTh5Ab3I7MGiQySG5z1n3s9MbaozbYXrafuBF/4hhs/VOhjMGi96vewJnim
7lcjQpsukEzVnnpuXciGHntACFMB71sisaq/oTZz9Q1uO7tXvLaf0vzZfYlYWgSh
WNAVMtBlid7nVf7yGyciJekdn3lfgSVxk9el8v+abXoT+Y4b7dGes4WXbgtF6BP2
f3Sb9D5WASXRyHQoSNokn1EfQ79qlEjDq98K34K6xjQaVL1bt8WHFV5aC4DVKGtH
SYym+s34T7cbgJt98JOJo8OsLXlOCWpcnY1aM0fmUYJAJbpWoHgxcCxy6GmN8A5V
HesPH6MTx2naWCxEhd72TcGPgamgGGOkI4W/QrjEAQRHsfikJW0fnTryMpq/pSPh
1xIp1rUok6L8DDmmkKmH08fp0uibFr7cd6sPfZXFrLHGP1kEJt+Rluu9j/DlILO4
X4WQw9zn1twmDb4UI5mYV/QyNfR33rtAPBWElUN/bRKMFrs6GzJLXMaUVmrQVuQb
55qvB6GfCs9OO4fmoDOXKGBodLPwYUztBLEUzOza/dFkNjv1LTYu9MVqbmNxQnSU
xGgZaqS54yBLJx+LO96oONRoNkPJVxebja1hbnlCrC1JRwcE9y3lt/kfw884NJvp
TOxLIN6Lsv21iwvufu2sl9kB5kffPED6M6JT5ewgQUO7HKJBVeBJiyjlG7XSp7Kd
ch7B5R9d8nqWGZo3YB6HYvmwH8jViepW0HEIDk2Gl4k4BRFi2ZZreBKxjym3NXhN
bot3i7Q3zCzP4PqGwkoiu63/sTlUMrD/HPyv1oa82GHsGxyhL31aITuR0oGVh6xR
2BhUE7mwQUbk+7U0ej7qxOKAVB3RJEx69v8b6ifgN/ldZ20FLVvjK6l4L9o9UBUs
cQQ7RzY2OqZcdTyjbXpV8uQZg1yk3m615ugvTpvux2bPyn5hdw2/1YHhViDi4ndH
6b/4IM2pwDVfTVsVUaReiYg1DyPVbhiJC+sNTZ6SLTHwtcvUa4/ewGpDeKSUb/+v
j8PrRFDXx+G3//pe41LRdej2udiVvanDZwAS0hSF6moMqZqtDa/YjWxuHvNz90MO
ou8TXXffxe7d9VssP6pI7bhp2tD0QaztzIpmlStso/q8BRx68fgmtypCErXOddJB
0ScYBRLHhxBd6QlIpZ7Co0axJFo183dEgyiv4mPOp1xJP4dt3zaqy4hSHPS5/yxM
2tO0actT7X1vU7TWi8ij8nDcBU5CQfetI2gEkywpmjNz6FXO9DsvuACr+pHKeEPk
fZwvfYbXqxVzDOdqVxkmJJpVd2yipLGQDc5eE3Z1mv9SH4wQ++KbbIK/6e7Ekdkq
b2l3550fHqhlxUOR4tAPvD1l78DjSiDdbvxpxg5XOefiUlIeaws/QjEUi0zXtztA
JczZW0Afii3PC04PBnAPWtbaZNFltO4k6kwD4AGl19UzWPye5VmljDdH9nhAGMw8
F3xXr3/futdxEFnEkHcU4giSSoU0iORHvxdiwZ2/wWM9RJYKQJrD6RbsssdlGjZq
o+gnkPou87mMOMG2Js9AWFizL+LeHuO6B90QfIPoxUgGrmSRVfwy1oaAkUH44eVJ
VgqO3SxY+MIUpoRhMHSXzv/Ksc1/mX1DOE7nSoRgDZ4X6bjnDY9OUiIG5HAGwo+C
7dUXdEF8LClsHWdVaTpNUqwIZQcLi0kuqfly8tIZWer3NdYmmSbaKzDu+RLe6IVs
LBhrkYQJKhLqZ4J1bUWQ8w4nltJluW01wtk7qQMU9FZOfzk+XNDjyUx/RMHWLTjI
q1xypo//J60YGehgtjzo+oaiqtreYdSQAEzrui2gfAjxzt/EIAxLzxIFX4EIPqXn
rV6cog/UjDODna0JyO2ZGMYTQgqszw4hB4oAcbbtQZk1vnDCXOYnChmf1w5VmKOs
hrBA1ibGTiJtSNR5Omgi8tAVUxc6xl2wX4iNYEdofvpO0nxgGD//2Zy/78A8eyCa
Yi5Y6YQvPxvD/3nRsERgY7X6cUW1HeHEsV1P1gRKWzwdjWcm1Apq4YXFrdkNgEfI
XGdCpaMgDlpf+YPZRZ9LDZJomCqEAYZCdTVxIC/SKQrFQKEBewf7AwnSGgMOWgrf
DnjNPOD56/iiu5Ppie/xs1brxdB+wDaGOR+VWy8phBS4DcomdeH1Upr8KNucC/nV
pU1N23WKJWDvtYSACuALTDFi0228bkeeLMEsFf4u2FRryeu9Uoy/AmfPwG4P2pDS
4IKGv0uM0bNV3YLnKqn3ASTCOwlCrcTg31vtvc7TsS4J1yR/WqeAV47zteuJp9Hr
wGejSPi6mRZklEdPLRSc4Ryg63ltL9wgfUvipolzC2P3i+VaNvHw1X191O9oBs4y
s7Rx3gQC6SiMhB7rRDsvuM2J4mtFbDIpWYvqrzyH9PK/kZB5HgwmAzISXvwUhh2i
E41hDdR1LBmmk0sQIL/0H+HYugG/2sf0t6EwbhQK/eMnt9SToVPyoh6Ds4SriWSt
6h7R9ofNTDxPJpStVD22GYFmgdXeuaP7KkR0ArBXS+SlX9bRZNXAhX8w7ed18C4p
qZwRBuf0Dvg3KvbEQskfhxYNcCnaqIy9RcgjCbLn093ks+sYcevXxzDkuR6kqcST
LCqpvddrwCYpx3JzVZVLoGN73vEPVkxq+06rpYQQAWmNjSNXO9o2Asx7bJaX8oNX
10N0UAD9YFh3Nh7/p0Zq3UwnFfM9hA/h7t1TwCHuy+/ahT5waEqarBojSy9Ek+KC
3GEE5pdAJ4+NoNAuuymVvXX5PACVjzPlEH4BcSlalZkpI02OVDvWG85FCvH3bY/1
lJiyp5iazJKQw+I96oUwiQtKZfQRbU495t13tLaBv7A6ivdmjQooNu0TN6/JSGqo
T1I8I0NaXkd6eSptRRezk8pD264+VJ9/imiGAtzn3GTfXIxSU3CktWkzEi0Oj/XL
z2qHmjSsGovKl3dQpd8NHvaqOK7kEnwTSlGy49TNA2I69mMCBYAl7sS4ZpXhLvJ6
TtI6vjmLqtohXzyKz/9chfTfifmbB0Evbj/D+aJUWIs/svz4vWoMvp0GLwSJjFVw
67MIAUJvjhD6MQ1PVZBnMo6aYnbpADZ4ivYJneaBbYn5AseaDsvAeTmXrSrIvdOW
MY/EBULmigKlVV51tiAmVPY24E/3A35fx0sdJqsRjjgOmdeQZh1R+mKzcd4xnF8u
jiKG7hawSh3djqN5HhUYc5J3nKTWrU3bCaN6GUTLWoWnZ90aTUQy5EnPuXxhIUSa
ULb4vaASGLybNLk0nT46SyC3mUmA2cq5A9dPkNx8nGgGLEF33mOhOZFI2FfiBbzY
Q4Lq7Abtq0h1steEJbUhYjEzcwLBDph4YPbMsD+c84CdZnIP5xsbC+7elCgXo8jq
tJBvpgb2mCN1w0/zy0CEzS++SAQweyRIGbRyBi4MLtOwQeyQii5ecGtoLuUdtbIQ
0BTlWMIZi6g/SgQjDhH9MZrWiagguGmLNOuZcr9OWF94EjNQYfkS9EMY0ZqAJLEQ
IGiC7/94m9mepCrgrku87ir7qcXK3Gtvh0s5x6xaTnlyId8vuKC0RsIMCla08303
rHIb0BlzHIIpFdmIyI0mnSmBZwl+aDj76CEgN07mzS5Vwqgwa+8Huo5rv8uvf5cT
VC2K2L4ub6sYQWRnv8cFDMauUyxnDEmXax1r6pGW1Tza29bwefQKoWMU5opM1DMw
q2M5ra9eDCeygumA/4SGV5A7EWbFxr1mw/7akzoz02zoX6ENE5aJnhLhIQpPyZQg
tfVfrxBun+U6+L38vwkeyij8BmJprS8rHRNcoR+TORuKuvTSzpJFSaZrG2br0Cn6
j7yVtAcnEqIImmoNoa1tRQE3JbkQM30qWkcQcNNWSBqZxMIJiBw84GJdQ+VR4FT4
fT9XReQZS056Cwb/fug4ELfQ4TgLaNrDbQQp2uLOBmAg2fJzH16KEetGRNFMMiL/
+V6FuWwv93bU4eAUrL6WZx0C/hajDJCP2nYLAOq4hWQWfzzS5JVvaG3qqM3FxgZ/
Yc6Flwp0aR2yqsqI6Rmgd9Y8xaOIIRlTr11/P62FndwGqe0fm+xOCARxjK1mKaN4
hnPKMRvqkiQ+H+9jMBolPQ21e8rAx7Z0daHAYEv07rW1b4Vqz+7fUwyzxn2V0rHx
lZ5JEg1VkRmUERHtv0+OUJ2+qXDATaPZe3iO18kxWqStM61YDu7EX5A3TyUtxot2
e+prPHNOZmGQkDNzGiJrE5t7lBazvjRwPoi6Z9mjuTxH4RW9xTUK5ZleBqRvBQnx
Pk40dgSGnwDTkfldBCFq3eTzyB6xj/Ax7ucFoO+W5QwrQbga3c4S7fmDJ9fv3VVt
cf6CRGJZ9OEooSOFbBIQEyp5WRkJNWg5NU06+I/1/qY9rXXw9o1KQ966Bk1/ldSx
skwzP8+6g7Jc7SKPAlTNpJSi9D2MdtDGoT5SmHF78Y4JwXr2p4dP9Nb4RzzaFgoH
dNA+bQGVt5eID1o+UvVXDwLU/+pFsi5WGDQCz8bplvFBuXcMd8FNJjD5SqQJLBl+
+2Y317p2ZvdvVbIArR7UxUeFC63Eo6SamoQrW6XHCKc51gmJrxYx7TSVbrpXLSNN
nP94pBg8vGWJEc83zoC/0H/TwA33Mth/4ARhB1Chmd+TP/hO6I0qD9NtS3P9+udT
oJExr6DfKSdrxMVzvaRypkOIUJoLsqEzD0wcn2Xwm9d3OWU2YUuhXLRMgz1FvPXE
XSezOfZkmVQtJgbdJ32UjbNZnLjUlHDvrlohd/H0XsX7egTZdr1yMapbe12iDjqp
OVb5EXh+xGEsnr78CYCy7/uJuTckXG+XRfUaQPOM8dmUaJ4iNez7xsiMhlH0azYF
CgL93aFkt6Kq8qiSDeUj6O1DgzbikE1I4sHBE5KllAATzS+XSmy1KT8epdEldFr3
dQEh6TZ9mYro9zHMiRc7FEooUgBa5WVJfnZb/EDVB4YJDB61+Zw2XgBlDivC99Hc
Wg1mJ0DlOslTpAoNS7tui8wGVfxe9VfD4+YfgwXAa5Q3EksLguRciQEBq22JDkLa
Z7+yzBCvB8Zmg4l0WJlU4sU8G9eziQp6D0VM08UpKsScG02dySkS4eJd1iLxckv9
nYGKHY+aeMoubNszZyybu6VZ8HwBRLxTEdegp1/RBO8VrARgZg/JcSFzfhg/F5qS
GvwOaMZ2g34kD5bOOabVVEajsgmjxRT/9kaQe2/1ac+wg/CRofxUmHIh2VH8uPp5
5YbqEEg3OfIjITfUzYsiNggS+NDCXTJXcauyAzVheRHLbQML3Blb7zwtVgiOlRHQ
dLqBovJEHuGsaheQ4zZ6zNK5JbMGWxgQ6TeF1HvI8y5tSBa5mqh+5vATA6CJkjPb
dyUrXPrSHVTeQA/2hlK/EC5YBKTQiRZsZchgnNnLoTgh0OgDkHXASvloEZ6HgepU
lHT8qJUDEEd/p2PqE4v3qXAxWXS+IhfTdcnudbT/QpuXWjD95Q8D4hiyiXU3pcpg
8xEChfnU/d0TeAnU2NK1ZTqvS1AL3j0Y5Ekn4HLNnGCyG53d5U5rXWvfKho5kyZe
YlgacIwQxgUpV4nLBp1FHIQ50ig+TvVhSQiRayP+tEL0uVIMuHuR6TPZ7t+U2Wuf
fUca52GuSsn2TRPGlVtFswAd7HINxfQnC1zdI09e8+xIP1n4uxFK9S1edXC6w2ay
WTzLF4Q9pLx7Fo6NSMSwqNALbvbii9XBPCMnYUNpFRmp7WUTPGym+TfEcJpbNd0P
EEPaLYVfWikIsbtLkLh31dEdR1OSIkIn9KMM5sSG1anAgVQ/+7G6085qn/KjfQ8G
5yw/mvlvTVpmhi5K4lDytWXnS1K0JDgC2LryM+brqnF9T0RwE9OY/eeHuQv28Uz5
7MjkvqS5GUtnA4zjBL0HLJHnYPuFnSiZ3BGD+WYJ8xQofiTZA/BSy3p4sCH6rWld
bZd0rNQ6F6piNzlHKELzsCAKJ6b9bc9yy6A2KBnJDPPekAo7WSjpT464BkNYjzTU
tj0pl6DUm2V3ai2o21UmvEi0pPfHtI25OX7JrcAUH9HNnt0uN6U1pS0DR17cA0+o
tVajRzNyA8HYjtae7pHtUvE2qFHr/uQIq4fsHex70mI9wKIuEaFv+Rezu83DdIHI
nJGIVlEs7KIMCsuZm23EDp8d55E/Rnq9SVyRLTdh64qFcwBsBUwND+XvBuI1e8R3
BvSs23vp6zDy3Zim7McJEisyukJyaUb7Lll7hO5oV0bJEuYX/54ebhqni+J1Y590
8D8e4f1UTNQws7/FLpGQwBQL4wjrsJ/+irTyecASg+ivImeYJQgGe58vdGSjylLC
4sLy453Ony2Nj8vTpqWgVj7ufI5N1S+fA69YZJlaYlW9HrncQddSBSkZU+PA+IIn
s+hSmuco1mYso/5kfSI5Lre74h5r4zrrITtMfLNVAF+Iu70zaq0uV0E2FajebfRI
3GF/yXzqL1DeOrIxGxlr006L5q0I4AHeYp/53GZnzfARSOmnh/xF5PvHMfTlBdHK
pJ+hWFML/E9wt9XgkMAr7PAJlPzQWo0TTeHTq1kNRnXoWti2mvf9wWetrqw0+AeX
1kZzD8O7/pFyzujX9SfiFFxul9aXUMuA1WooGTL0lbZjRmFs1YtgFUn+bNVjcoOo
7aJfaAbmwKEmcFuhJ88DrRFMy6qT1VlUN2FP+Vu/GmtdyDFdOMvBNXxtgy2TOiAb
eUDuh/n8l2hSFLX5W2TraM4K4bE1Ut8/kpwnloXPmkPg2Qq41bmIdlZcyMJyua37
4lVMUbgekzh40xYnLpkO12t5ygy3A4104Ghj/5Wf+vCC+XpQEYTUIMRq+/4Ix7HR
tDxiLAV4CLReMgrU7vdEQMVk3PCZy1tCpr6XtCKdNKnqoyMSYFu+pwcOyEsm5Y/i
GQIUvN8QUBQipkh1UzoFwmytpN5npvwBZMiin2bmI/kfOl0+B9Kmc3ZvnMzFylwv
E+804bq16r6KFUeFRvKxTqEK3Hq58DP1RrB+3HK5ZruTQM2SUPFzX5hgUybYz0ra
9xNsteHn7w+XG1jDJD257RlUK+WWhTEeuWjyGvGidoLa7mkusI+p85Hf0AJKQqxv
74p5HL7v/EMO9zkAT3m9ggPvqKT44HrSuuIZ//jndczdRH9J6yZGvhDS2T2iepxF
ikouPPNzlRBulUupUNTWAJ6Fv7zKGoPMHLXCToxVJf9AvFiF8nsJRx1CDVKzDieL
TZCEBdKTMaZ/5CcHeU69iFnb+OjdxQTxT+FcnTQFpjuVS39Gtny13Vt1HHAYK+5v
ttfzegpJOMS0MGkGdJu6yUeh1YQX6ABMRNlKgaNjbd72vQfBMWKsmlF0FsDYxc7f
gv/9zUX069LT635WhOekk6ApX882Sn5vbiMIuUfion5uLFSuOzxtHFzQo4wxKw2B
bQofj5nibmlATziuaYnxQLizt3GMNsPGBiknEz/YQsdxK38fajy2cf64gWOmtQcv
yBUn+GhptFEEpUVOwc3pTzEgdcaLH4cuZGZkHIiyG557QPkj8Ez1fMDiLksMfiaO
7V4i016ZqRl/SzGbLhwPGV7F8Hhunvh0yQiDd4Cykq7b7R4P1uk1Rscjq5zgT9wi
YjL2c9yQljSbcewNSa0dwE/zg33SCp/3NJHD2m5IOVMzvsSVfQJAfSc/NI42njHg
xCN8JjIcTgBsvv4N6pcQX41TEUbeUOe9wCuLBo0HLgWZqV/hkfoCWJ810UtnIk++
bKMZ7cu7m/BFOFMJL0Quc+oRlAiqwZmnr5RiJ6PzAR2IgAldnnTkPsbY+bzJ62aA
TMyj5klVuULMAqrlSWAq/5J6hNuyX68f6dWZx8XHaJhaeRi/vgFfI4i8Fl1rAGMX
isL9zI1dII/4qqOw0lhnUzPKj5v+HFvRSwlRKtyZquuRFA5+s+/j+g2a21uYwDqE
o5F+p82urITXUi6UKBPKFvn3QNRkfFI+sb2PlnDNOOo6rmFlG38xzzjsiWaYus1R
VawJ5VHkKrc6yGbRiI5x8fUqT+jCcfQrSBxpLan5kH0W1M2RWjby9crzBi9O2xdZ
a+3/23MKS30WIjIMVvmF41gGIN+2VyW/9gRHgXMVxb4snxsuVInxnDA+5nKqjJqt
8laNmqSD1xe0YZuc7wdmCOmHWCzXwyHqc5RFo9oCpOBN/ql1nwpZ27ZHuRpSxFrm
SDkC2NBL4Kn9rVgKFc0FyWQa6HhnktR23+j42RoR8OyWxCKo4FnGky20YOF9Sdu6
LrqC1Pp+jjHL6s2D9alnVRGffsBI16oMotjdv43NuyZiahxJTGAqWm2F4LxiNO62
JDfreg7P2t7BzhNTQMUOVesYnpvgNNcWPaahfHlhlTBYHn12R1AXaHIIk/2kcZ6/
FyB3F8psbtBYDucESw1Yw57lc7G48fsc/+SeQcCRH0742TiyZw/Qb12P4aB1maAN
wiPbG42I/+umudPufAenfCj3HwfOTFHd9wMYaiBH+PrpdLgK1ynPp/gW2mXhZmWj
xsrMmzU18ljWT1SRG06H13SEl8T7HBrjENTZI7nVG5gE97ZAdPzfzpNCCY8ikMh0
czw3/+DeDjgPhtz0nmyYLIzd/S3uv84cGXdj97xgeM7EGiz0ExdjAsN0CctgzWlr
OXmZFvF1GDAkVSS0D/D9vH+PL04wEYM13zpyy2JxfTiZoiJuB/0jNWDz5A5li6G4
12FghWG008OzEJvrJZ7DOO0EmVKSe/qZG49A6iNpEBjyRPPPkBNtCoqANPKkkCL5
sDyzZ7SJ72/bbacufDbqYwRUkXTnZZMvRwcn3qlCY1oKgKQlB/xdDYX/2tgp+zTG
FEH2B7/LezpSV0zWMRbu6r2Dy1yNlUbALUYVcun0bE3ZcqBNXU9r+p2ECdlFk1wz
gwNT2XDwjmqjazDiUGA4ixYlRD8Ts6O3S7sEqnNogh6wHvv2D62rnoAP2MIOTLO8
/OjfBXfxq+TgkRp5y27JA8HWFxf0u50ctC3nEJS4Gh5ZMZEvquTuYquRTV7p8X6K
aGJ+BXKIHEOtZb9JjVT3/Zv4zNmDBEJyhfYdkctAKKms/c4MjaI8uxOCdl6ZtPnU
Xd8knQk8d8I7Dl8WAlMAR6nH1pR2++Lay2ZTiZKtq9JqWU6ukEvSpepfzwHWVFJk
mNRreVzS5yIZ4R5Z8vu2rlan4pPj5s49W8Eky8g5AYbrZiwtpn1hFT7jj02MF06e
/VZ94pOLGKba1sVyiPMx+mqb/4KnCj065iC1mXxrSCeiGNwVr32D+uWEYBrpD9e/
vVQrHsZ2zUb2y2MPLPrQmF0GY9uAaGBaoB8ZISAgTWzJCXQcRn0xKACI4n62mTeu
XfhqF2XfZkFb1j4LHK0QKHEQhV6LgVDg9MJo3eKTCOCstsF/EfzHAxhG1gXU7UgW
zpEckgx1GzujH+GYjtD4/RciyLzasLyNqFpUVMpH/CKc6991ZeF/xNugxlkKNIZ3
EqJW2QZ0qKj4WyiaCnhGcJ36f4ouqtwFgQQCweF05b/ZS1sZgzuVhaVoFaG06iIe
FNteCM+chx26A8nO890jQtD29Kd2WpYYTRqbd6C47vz4TBHs2coySjgPjQQl3MnS
wQeQGkVz8muVRD/3sz/4UcqxnnfyiIQhxxORJjly0upV1CyH8iEioteN0I2Dre66
dQpJIqgMK6f//JmeIdSBB9DNphAMYo4/wv5Vfdep/xxV4qkCJ5Ffd00mruw5Xdcd
YqKAHu9DfwUm3M2uNq2mu1lyYUms9dRfNIGD/TblyKKuIr01cjsEboF76U/DPqB+
FFBovqLcOOFRHEIZ/GDT3gc/x5jSTJU4mwsdluftYOdR95HYEZv6tml09h3pssST
bPTejpj1xNFqpc+b0zHglcrOOvhkSCZLpMorxPB6a1OGm2gTt87D/NkqHtyYkm9X
ilLNC+gM6/TqALKqOE/DUpNqpB8CacHaW/Eub39jnAn0I+6Rjji6GR0L+Oj0EwTc
ARjeE4NHbOCzY3p14mwn4tZkBMHbigX+X3zLAQPk+bTR4BDElsBPt1pzsH0jykAv
54H/VLEwpyI8t3GoJ4CvEa4ddb/IQxuo8A5Ae7CpOuG9vPwR9MMMgCMVpm6NwRlb
6Gb3MCmq8xFpJZ3ljl515QqUAELXql186WBv1KxOeU6304C//CxI8qNUzfBDd+RK
m2WzONKLP7XOeUW7pfKKIgryR3YjDFYpNnbjR8MDxKrVJ78N03+lLRvFEYxUn6Ic
W+T6+XTRos1efiE9NhnsaNslyIiocC+Jw6MFtrsoT68ONmFH5fze7DhqCNZ+F0AT
LgiuRhxeS2miSMyMyOnEIDaYVh1ldMDrAiBaEEd0q+58zq6b1eg2I0o28zjgOHsl
7nVFWF64JJJFP4OYHZ+9ss6xw3LsjmFq4muXLR/vHF5KZA47q/hKNtMSo3QI74mc
97F0OI/hAZR2hfHM68bxHWVJX0quznJWhW6XO304AtVUVu4FBxnCRkAJgIO80VHy
uKlHnPQIorrnBcCl+nPjo2/xQeV5wC8MP8JrDiPdl+vnrH5lZCZqPwTjmfO9lBue
yfJ4r8iE48FW+h9/TQZqXAo/OrMdPAQdFU7zxErwsqzJR3XCldHmdxIqxtEZfvKm
7bTFoSiIxvUmuVaBnPdQmHHP0T2E5h+w3dMNgu6FBsRP0w4MPrETvyLrT/H58bgs
OkhgJurd6+S+/ddR86HHxQSEYktcHsM8a49Li7jb3RmYAhnqNqOlzW4qrOf22l7Z
nkwrA60+csVZBlfPLI6g0kejXygZZJ+3lHzF2w6zDK6KGExY+uMlRzkP8akTfQa3
MB5u4/YjTPkN/e41PoD4WMu/OphjqqTHWezxSb1/q7LOHrlKvsQooEPyyyIMFl3Y
czD61ywo6AaTSsJQWZQMT2I+30LdBb9SR56bAKvzopvX4cRemgQNWHYWTmKRleBn
WAVEleIKVBR/p8oOV2as+otr+OTZ5JwuA3ows8LXmLf6W0VFPXMIFpqlJAV7cQIb
aLyoDt8TFy284fd2YWxYcD9OxUK8w5Tks+G6e5ywqYCqFrmcdeqFCjxlmvKAg9Ml
qUIiGIj8EKbXoUER3VBCHLgMlpQFNpXGQ9mCKJDsX8i98aiaHzk2bIzIq7YN8iIu
ER52PESHSufBWzC4Y8uzp9pPBjgy5wEX9q5wgBJNlO5G2tFaNxqA5degS+g2fqfe
NehnCkjbwavW1eNUY6a/Ck4MxtbDLJS3zrlXHbvao6O7Jg5cZbBzvwZUtZhl2lWI
5t9Mhk7m00xG0iQnrqpVN2G0mV5UdP1dndKZEUE8KmBjy9r5ifkU5KyZCGYYDZWW
PaGzamlSXdKHGr1jvXrv0kuBdAR5PkM09zMJqlyexkRtPRNWyr58z+zewPkIgpmJ
danG7cv6ZNTblVtdR+wIPewics9oHX3RN6gyy9gre4DyVP79JHlAYBLm+UJLTTN/
Z1ry74jSern4PrV3W8hLBmeyUewMHq+jBqcwIKRp+ED8QkPIa/dMSmHQOVR+ITjG
bCrUe1ukPTpTWYSN7kjsdZmhwsUvQ9KgYdCgoLzjyNQo66vFeWJv4YHhPQPfS1hC
RTNQsKOKRALZhb8biKw+8JvPDjIZhgQZhXNSGlekg68MhJc8SdoleWP2rDftyfkJ
9lmg6lmPQ1wjfngaTHNQTWrn4B6VIqRUu90EFmXF+DEVFS7zDGx0AGiivNxTwU9O
KgatQBbFQacJ+4uAX5vQ8WUYd8SQqQcVkqiYmDrAX117iJAIxCp5Oh5WO2GpDqjH
YDsC+tb6KymGtsOfRZHPgmsH5GRCJDTgmJz6ral6vmaHDZR8GqTj4lewncs8JhDL
GWoFbtf7RoSrL8xuxzZif6WyoeYE7cs+0oVNPvY9XLmM9+DGnX5g8XJduN87ihnU
lEL1IGgSoOPbTBO4AEtlkNd8dMKnza/FBBHw3avuD4W7yPBdD+2tYg9Ng0Xgci2V
lyoVPUrNEQriBBH+ZYStBl7B+yzqpXRz6ZvsNVNlpeCzs9XumRP4ZlRqlafBTEVv
pHzsCNPc/QBd8980F2dFQ50XE15pot54/wsu2i++b/V1Zjpa8kLwbd2h2wuCfjBA
jdLZ3X/86qv5XHi6ftj2/KqqiRPks3c6Oq0JKxLvpCkFDbRnU8ewylWE9hZ95opf
iPUTmmQ1PGHSng5dFae2w0BD0fAJwC2JhcsLKI2MVfhQoflrH7OgWNxwxM3TDRBC
53mOLAEsMMP/GNmjxZ18iOjgUYM9d7v+NaJ5hIbL61h/6TfZms5uDwuqBWv7eSlO
yW/lVCwHno7RK+IqoUU/nPM17FVIrSjOEPCSv4BAgyq4CsHba5jaj+ucpXa+chKb
1i82VeCiVLoP7fcAENY6+bOpMhZJ9HwxKSlAYkNIlwgRegTSRhFxOwCM1zz21+db
02k/SYITTM+T4g5haE7eQ0pIF9wtFPJyWX/kYOckVlaLK/ywErwsSQYWJ5ZgrSA6
xcy4Dmas5/8GvX7MGWWPXdazMN/8oB4LncumOZY76jdOaxQEXOpz/bPrDGk626bE
4N8EoIuNyRM+fDUhOFq87N+QCy6/Bc9b9h6zyiDV1w7KznPJj+vh6ATY2g8gPhai
p9+sjGM499ejam8qX3eG4ZzHHwUCyq543A9ROrXjD5BQ7clYfSibY9GYTb0IFkLo
Vv1Mmbkw/5F4qXOI606g4WXF8RtUH8fEICjAd12Ukwf01KZV1/YC2p5zx4Wgs7z3
VQOuDORVQC5z3Qn1kHUybl3xYZByy/ZsB04r8qdqKcYyxgEpzT8G1v3uxoAMyAsh
xwanczorq11uwr2RZ6yIOn1JMfY9HI9EEpZ48B5Wf/V6vq+PVRk+UCs1HTV63HMd
bhismB1flrcejZKTBKGyI1CcS2b8L4DIPVcMQeYFFGEJ4qEh10WB2JEXcJkxRt6r
SnkgY4EG4tETJKBS27sU2B1S7s6pPkiEikp2Hw2zCNZn6lQS/Lv6Upi1C2rtKGiR
QPQ6c9B2o33DvqosKUl2/88wDMQ0qWWAHUaD06e6zfO4lAguz0gJVMtKnYzt+oR0
AI3sNOSZNc6wWJkl4a33S8cEJEg31fclTF4WKq+e0o8Xnc26yCPrH1zGloThTxkJ
M/B+NyjR7pjiLdhe7U5HxuRX0193dJl+pT+10ZcrBpwcpZdo2ivHA41WmVU6nTHj
8FlUC3TTbOv55PJhaArDfdvbuQXigH+JJGDEjzD+GPJ8ozAvFaAs5ceLcEakcDUh
yffuPpj0tjbrnRr4fECJlXQz2MS9vlHBfMBg7OiTg3sBn/KjBiW4Yah78j8pU22o
im7QpVC8DTUkAG0ebwkfpZSfshnS4DkIERtexPCX0054qy9JOzmCkKyubGxNl6aJ
fOj5SdfyYiBgyJjyhu7+S5cIbxua66b6OS+Rlp4YLlwWXWCD+zb9ppkfOz6aLV47
5FdeRaUhwYsiV1qSo/NrpprS81YeQKOZwnhIttz/3Mq9mOAFaQ5FlREHx2QCwYMF
Se0RH/k4YRYXBy8FGtAbk3Gwleb8CphPqSAiYGYP656e96kyQIpZdIVcQbSGcWzU
rNbaQVjFcHrfbXZ/VOOAQWjIFoHNiYHBeQzC/n7OlgYYCGx2aj9W4tIsSj8xTVOZ
cdrkNQY6pnWchLNxvZjULE8KJcdIo87Dh6d+AdNzdeX9Gv7hRBsSBzcRUnnwyOgd
yxuQyV7rwwQVGDGdVQaGw5IB6N5xPL+Zosip2yRzQJROIxZEEwrqucQTyacneP9P
+poFiGzNB6PdL0zEqu4vyK1BrBNcgbQliCsedQAwcABNqUmKYtB/qUxq4fpi772F
JPm+NhMMsWM6Scb9ckogFcidMDBbJxta8i/hMRBhJEKO7yQqPLREOrUTpLGWSWzh
S1zs2gaw1/UBOc+1fbbdN/jbwDq7mYYEFdApPX8fubYygraNCWsXz8lG72qN53Oa
qUZtKuBxERftGFjYWWiK16kaqQsc50jgK0YTrDJXeMhVu5+TzvclsWe0Mcxd6ly/
jiydPGgKc/mxpS2iXV9hUE71bH2XETPvpHmtDbqIj7JiJyilOB4j+i3V8+iTghJw
Nv5ThYRtgbNGU0NpfkPfW5iUu2e36aaz010sXmiKM+nGA/TDZjaB7yA79xK/IaKG
XEzXMUYcZXdxKrkC+iFKzY9y8dm8rvt+FALFNhqh5WDJmB8tFRZtnfgzwCjfI1x8
IalIFqN8pFs/Ok+wDUTQGybWTXuwNNo4yNH33+opycvb6unWaKGlcA5N7urzK9Cg
22xeNUJYzU5zO4AD8V4wJmzVAzruetVAWzwUvRvk+5ubX9amHmXaiJ/+p8lAZ98a
ft433QHGb6wxqe4TQKfyPAQ2YBRnTfghSigRHj7QXABV+6RHwkpLfByxZm0vf+Hm
+MZt6ans9JN2WUYUfxwXDBHrg/X8sl8KPKnCxHQLbapy3v2gUz2A+1uNiQgVTv14
NnzNuuts4J1SwR+sZBe2NmIkahrE+VSwb7JICTMaMdwPpMPNtV3R577y4Kmv5H99
62P27eJd4yF5wPKO4dTrSA4x8QxTB+Dr8dz7lCHaWAbdQk1Dytna1WQruiQKG2nT
Djnn9ohX4QvYje3NCfgeKIhR/0KiDCUoxwa7W7eyoFBqxrvI2CYDPIQiPcjYq6tB
hGEBx7nR7GMKhjaoXh2ud7bBArSydkj6cLVYv7YkNfNRthIciQbV7D9i1haL4Cva
V4mxKMJkOdJxIQgAOz0pXwlb6QsSB99fIxRsn0PONKIDG9GoI1R75qH2geetQF7Y
J99GqBEHa5+FX0vL5wKmBqms/VX8asQzvWssJpyAGkNLVqZTkFmklV8ccTWQuX80
oHKGgD7rLn9zupJCc2rDFc/P61Qv/KnESC+N1et8tSfpotJOupg1IoRcLDx/JCgL
1i/e8x+RZ7BFpp79AL5Qai9SwKV4oB1foDCXG9ZtXUEMcte+UlEm0zIjCMzXa7UN
GaNwbUVw9HbV0f/a8U6t4BHSTyXmc3bfkEoVx9XqQ/O/EQJr/tkMiIyiMqRkbt08
GGxJIll0jco99YdrERA6RtOf2wGqzSbov0/JY1Q1ID48spGjeAygcBKvIQ0onSQB
xKZ63PZ2IxXsRm4I/nWGRlprZGcMZMKxIobKx1KUAAy+n9F/c7E7mWYi9P1u6ENy
8T066qiEoGyxy/DG65Xale9ixW24MoZLWQmwbG/fcHKA6hgtnvYL2OFFCoKlYygM
XyAdPlo2+AquqSHv9+iIy9Q8RmRzLRqB42Yp3PW2+mmBTFPOVmP2OnjQzFfwmBWK
JztEg0ZFgDH/Tl6i0flbiDuc3gqemVXqqxYsSMZphUFFcy7aAu2HHJBTusaxcNc0
1lEMFcv3Ay96cMlOBdsbIn6LFG3B1pUMR878rhYAJqHXhUi6gmP5qOkBNJRa++1D
5DQG8yFiIOFbpfjwBwa58uWrJOdGB3Yu/YQztM+KxNKrL3TjYqcEbe+ZtyK9dqpw
ydozgkwcWBJMoRgQljWo0say0q/xGhBTvJcuNx8udX/Pmvo2CuI5pMMjJ7rFlprK
L6TntvTfsdIagGX5DOqECiQGKKuGsvVZv/B0s/PSvXkH3WIa5yUmzpY/G0QC25dd
WkbmHzErmR/+F5ydHuqi6ZJzJCXNpZOBSNohTCbj2yvKASbo2UDmeNmzxIejnZsm
GcawK71IlJiKqbSg21bbKv4zp2o1PrhrkIHR3UygALKeZBU789m/PT+0lNDCyYJU
Sl2mm2mIOj7YFo4N5VzcyTlzoJO/4uD//8eRi809XgHrTxmO+yzpdoFxQ2xlLXkF
qjidtmuWhgvc07Z88cM1KzZbLPG6y2DkCAk0eA1Jq9NAmeTGiNE1PN/p2R2tm38L
zX/FM2aiIk9SKRygMu72C/3j3hm2nxtwSyUyE8yXiC766OvvHjPVnDbEsqawofBw
uQU8NNMhMdvXaZ0wNxWq9bdDbzoPWNIHVyesa9gTHnATw7vKkbYSmB/0zBwt5y2t
IRh0PydFKlzzR/A+6ucXoTNmWXgNUiEeiW06IHpBZ8/UpBKf+I6lN9LV0hihiFma
AcU027jiGkqTXaFs1WJy8IhhyyCXyySIOvyTZmYK/TCwhATQNOTqAmhXHCBv2MYN
MIml4QgXkUr/EN9SNT7ghkqgT0VHwiasendKpDXpbv4pk+5KBjECpK8YY0bJWSm1
4pv+eFNaIuhQ9TI47ujBti6w441XbBSn5L0z7OQ00XC3Kc2nKNRqFSUvWwxwnWFK
rVtIBF1zsdKtPLdoS4KSqudGNvrqXR78fqoyjOkthSy8XBPIxmJwBQ2nsKEYdoub
8x6TfEjB6fXjpji/KI9eaY7YoRjoOgI6ki84R63Nfh6FTlJWodasti6vOevgqFz0
lndfw1/25ukAxmDQ8m+Z9rkEe38nOxjoNlNq1Jb4GV+0lTPs3Mhg1K4McTMSAddQ
YlKa+iUbRYW/U3BeGiHkDOwqd7QTIHVxbHTOQnvUmO0Z56mHko8aXsPV4xrqqI0j
LobDft6z/t75Al0wqVd7qKOWQtVE3aROTbrDsNNqJZsZ8EXOoQGYoxh19M/lGIVJ
ZoBC6DPMg0xlaOkYaGgV9Nmav5Kyw7KS6l58xPcMGE1575WjfxExlENqMvUJ7XFk
DoChW/p+pSAPiFCLNi7l1Ag24Xo/5B5Uj4jQ4mCWqiqxOeQhIUv20f4li9e5HOZA
3JljcQfeE3eUz02OLosQ9Lw3y3MWM/qf/Nt2KFuekVWOmvfF9bCvLj0dE9UoMTQf
4wwOmp8WdT9RvfYAWRxKmB6c4FcgVnB/Y1RBJTdaqljRaDxvYVHsQ8BlD4sETRDB
8yGeRQu+m/49KA4XJ6CYJlx6MUOx6ieXy15196rHusYqbzKfSWMBMy9zt2tcXYEU
Wyy0jSKga3+JV+xmSqp61PW2ZgNY/MpfVPRITJ0zTvGR1/LY4eDcNarTIe5hBrtx
6IFY52XbOFhKMYj0thY1zkU2N6fU+udoNMIwiine13CZ6BL+57tcZT+TtFBQF8Gd
7Io4H84tJ+zLgq9u9ELcZg4utZVe5xQ12G8ZezMmvxgXw6//b7oS5ZAYFeKjDp+c
wVxI6U+VLc/43xwBFL8Fgu/0xLeHq0IFV8NxPd9F+3lcxeWmVw2NZNoh7vEXJoB8
lUfXgHBciMxxSwbR0ZzpYOx2YZpjl0r+/6pz+349R1Pd1byJb1H4LWEO2oN7M6TT
jhextk9UXu0zgoC37h0IfkIvtByFrjFz14UXzWKL0cyRY/Tbh9ih8MFbt/u3ZBY9
D/B0N3kLn+QvzpRAOb5tQlBFgAm/HG1lCWycy0IPNm+9k4cAwV6QDiodP6P9UqNW
XKJ46auQqxcLQMBzHauMsJZAX8r4bnmy2ov4BgJrA965cUVrNV+PMsR0tXIjvX5I
WdylOTBD92XoDCpGutdU4OJbi6PyWuttFBVCDsiwCgEfxFncEe8V9Af6k+YxVBQc
z9iF1r9G9esd7b8zCmi1xz+oRMcYPqlJE1v4k8OhexHlt0oH1PFo+DOTh6udOTtv
qNt/4v42kaOiF9o4vrJCz1wu6LA4Rt1O+b/bUcwFOK4gNVxaSw9LUzOiivYlbcf4
JHioNog1X1LZ2nNCuu1WRd2leDInsE5agaHl0X9RyGnJIBaqPZdcSjPEcbj4LSpG
xsCfoMWbja0S3pc9FhaZ1FNOXDg86EeSOhaEAiDyoLFdeDYuJ2xFWLeLdsBz09ho
KHfZdlrLv/NYK/gOJ1n4V7+rJqgAOM+KKWUPaovBY8QSUnr5JWL9jqNgI4Ms4/o5
jKoh7UKhgteniNkWoQq+2nC9VtpCtOyxFaWueLbzir2Or1ur3w8VSX2A7qtqg+td
pDV/Rk1jXB49RgzcGARR53TQyC+g3c+QjWfnkEvMDius1yqd+njv6eRXkqKVpanH
GCNsxCyB5WX745g1yNigPHVr/PcHxr79eafW5BtcsBnjLQE44Yprcac45Tq31jsq
7svSLgiYZgZa7owKka5kGKDeShWACS6wU9CzyRx4KDkf3LthcmlX/qWuCwzF+DSz
YzokimDNOjMYYrTyxDNdX6o24ULC4Q3fn8jSO/PKF8r+uLGpFwMZRs36lYh72EBg
4uFIYxX3DobHjcuucl+m6mDtC6jB23PaDNhXP8wuc67/T/tP8/KXnLVkFgRYP7pW
DDrK2txakOwanKVzxud6zqklas039edfWoF0pD6iZquJujFKTNtiPlIXd27DVIo4
MEcDnWFLDHsP8yTPOew3kEe9p0akCG6oNxeli0knDrA5Qu0srcWH5+w/RAEwbah8
gxO6xl8J7vC+5DGdjXsuuyKY2oRsrs01fQVsdrCM/o+NiIT0GqQ6XP8fA4vZ815G
UY71hd/rKHv6cJ2c7pvaVvkOLRVUuRNu+/Idj/NA0f8UXfG/j0S92nYM26riLA0w
mwIJMsFqamxSz2eghtabupeXajmyrRNqkpFX/Sk7Yk9wBQ/qEOilLFhPCW3tr7Hi
TmEAozPlH6cnzd6XngtBjbsvXN+sqRaxSZE8wTQ3L/ZCsCkinWuDMiihPhLytXeS
NOKI2JLOFDdSBkAu/kmewev5vH9OORjcTpAPLLwkI1pQpEOpPN0xWKLPEm5B6zXo
xtElIOl7wC6b8yWCMmjcferDyIRKTsW5sDu6EtY2bfARI48fD26FqVgB0EBC1vhI
uxAiovEX22OxIgqvrtgiM0+tIvMXdRaTLUECKM6gDoYg/1U2jqNaKJZcLF62/tZK
F76IlraFztw7GjGTw3nzaT62Ol+UsP3wDi3esyFbGxQ+XUZCK2nMPeCKHOHpkhhQ
Vhd3CjcH2x06DT69RDnL/u6wejp+2Mch8P+JSqYh+y//QZB5THXShZGPFdWQlcSQ
x1qQISOM1hrIbucAgB1Xumwja499mSQzu5B+SD9zZVqVsNZeNR+c4S6qvlPQ2VzJ
tGJy4bMhHmn+IzpKr/JfJweB4pkcCdcxAEzeFT2Bh2oaHKWE/PnEyYbHCQ034Cmo
twKb7ADIkETk7un+6P/y0HqrfN1G05YIOQPD2BZuSJgymjzraaXU1ek8aIhA/97t
zoVEsMkAv/L2ZxGBBNTfo9Ncvhz+yt3QtnBpmQx5SLPhsLJeRlbuSty72VslC4cA
98eyNK6oeCNq/EkKpUBL76yE2aqebxr+Gf90BhctF9p5y6YjURArO4h52xwOLTn8
fR3W4sH9DJHYYxVdtuyDujhQdsKl5IvnMwXUdWfFbb5GCDGlmQnUDizdiI/O9ap1
kJlHf7NJf8A0oTIdZR1fqzrmp1SQ6Zp8c9KPIDaabPj8uFHxKPBLndlGHulwgzRr
i3mb7PhyHeEqlZ8MCk+wdaGJCYNsA9iCQyeFs6TWe+AeBonGjO7148uj4FIvcA9b
8tIceK9hKXCA6DcPXr/KB6xwrCbNMgJMTYETJZPKLglzzTaWJ3EpNLrrmvGeZq9M
HS8TfsHhieSeAh/TudDqV6nOp3MT78hPOCG+ZfEB3AqNH2sq6GYqx5cCz5HwKjjq
Sc38/K3LLcaZG8SgmeAXJF1lY9VAjPA3k5pW66WeZFd37JqBGVnMr7v3CbOeS/CG
XeYJ3mx/aotH5vO/o9TgpkR7WDg4o9j1IsYWEGYfo0soY5BDlb6O1V+scxXKF9BD
x1BFwGgBj2D89qsuXTX+ZuGoz9akR+nJSICqpDxZ5PeqEd0KbgfY3qvzoWLtkNyR
HPe15NBcXqjoQk8y6UMKJXVrpHzFft7yYCiFPSOH7o9JqifUWEfzHe7zAOkiFYps
JZMpIZSH59d2utb2UtJN9HecXC6D3VKvZKtSIM8kmgFSOBvjHO7adg/ttLUQIJfJ
9YlEKtyp0Aue7COmyGrZ3x0ZlboRpVyWRn/euF5EUXLJh70iTWWbOEPIMjI1FwN+
lIiC8K8gDrE55MkW/dWcOoMZ4EC/vx/9qXmfCo4WdGmp4oekIj50TUSCGtL4v1+B
S97Ee6o68oNM9w91+PEVkeWBMZQNmOXpOwRZbA9bd9Cw3GaMtUfjWCnetwB9swjK
nKoRDU624CGZEfAdD+nigYzB5BHBK+0iQMC+oviaMqEsdXvBmQVJnUwTXeeJqvih
2Y5xItJ0gBCXSSxh4BQKETeC5SW0xGQuIwzZD0yITOMpD6cg+M/u+Z/lC7XL2HHS
jJAtXajZG0hguOlRjopZppOnWyJFH6B6TaN920az7i9/vJ/FlL/ePClxwHIgmwIy
wB3wtP6VL5QKPDzu8v8sR+6P0DqacEUCCJfUYvYEoCQ8gVkvkoQj6wzUm075cuyE
pGLy7bVz51feKDM/K5hellZzZmcy2bsgENxLJhz9WPWW6C8OCm63CdsdLNZySe9m
elMhY079stBZOx2nsoeUmvN58jC+nOF7nm9FsOIkR0SN2URJ8NzuZsGOEcVLDmMS
wnglFDpf62s0PCljwOKKfms2mr1LOFCDWKRYM1P/4y9oK+bLymM9Egw5GJg0K+qP
JAWr7qfsPM3AQ2vsIv37WUPbY8OcyTtQVCDkYQsQR+TJLXA1LbWI54WQ6Z/QYi+U
QUDNWlOBjnfyDmBySAFAJLO4/VuL6soERQ9lI9Ha0tn7XZVPV/cxa8keLmj58DRC
S+4xJVJu6J3WJOzQNpjQHbPtEVui2O1Fy9dv7MS+5HMg/uY5pqY7/ch6fyFlKNqP
ohP67z+fxFj5ttQCwsWBcBrSglL0khhs5fp7pBzcKhseKEsKmp135dI/aTBkzxV9
cpustaxnC5z47us+0u3cytUwSeF4J7JLFLeiZ9h1ki0Uq2LUK0nlTuGOnqvBVbLT
Jm/mi4+nkf9a47TaqDCEKYRjAjQ7/gWPF0d/jpEPOupkOEkiNqdlKc1aHLEJvbm/
/UMZ7kXBPzAjLZNAsK9lSYfdrYKlCbopSfN1SWfrfILtwtx3P1MQOlAXDCpsV+g6
hlxeGR3cOd4BaySpcOPR+WASiftE7V2hPne0jAvOI0Jf93dJ3hwW24i3hvKGsRXq
J7WYByExQkZHtaVyL2UjJafffRQSbmOEKFUCjFiO+xGAw/uQXx50ESboNUZf/91K
flkaMfTtLU3MuriwuOw+HV0mvupFRiddH6xXYLkUY9EIpq/t0T0Qi2TlfmULeuFq
+uYnUTMwQreqnaZGu5cMj541kAUYd79mRNRkVg2b4scWOSOV8dqkGOjOLgDiiAUr
9XLUvqtohelpoBSYIbR3Hs77CJIbVfPC2k7kJt2bIbM1PQI0AsMpws3rOA0DT2Wt
6UhYus4+jXwOlac6ynSCUBTiBhVLrbVYofZBsRMsNp7ZQgDr1XknVkCoP41CWBWq
ScccJ9R6gx2GpxD8648fMIAc8PNTQurvEC3dnIXOdWU4Ntww6dgIvMaxZya6i5QR
px/iP8rdCYQTfllsPJHuMdy8/EEC9dRYk9h7N/4XOhdj/HJFEtOlmeXB7VL7Krea
6DjxPPk0hpHUuPYCMVkvKRURS9Z+X6ZiQm2Cw9owh076cv6rvcnmkZyx3Rnyz8Y5
Bh95SSjrg8Ogx2p49se4mN13/FjBWs5UV01SsO4mFbYjW7DqwC7KLjWJkgLF/Q39
5JabAgMl/qbRa0rmcy+zHOPyerJytOn5pfomCEBpQapuxdBIgLIpa+N2UULddv71
f6OIIi+VeTzmzSDtxNcgGGEb0iKPPzl7mDdcTD6sSkXqGqEkginapuZuJnZaCZJJ
r+vQXaEVMAbs9AsPMeXTvnXeL5fpJTf65zr7J4wdNOKgXJz6Mz4BCkWmwLxWkHQ4
Daho0wHv5liYHI1w6hGxWGXmVbe+HDUt4pJjoI9HjBArqBC1/LK0sT17mqXmTGDH
U8OnEZWgoEXD28hRdjwwEw2J3vwO39ZD5fkBUAQ1Ly7yLTDcZSD3ykiIieVdYOgV
AQ483MwFbvZ137DD2vWn153dTPlM6o+IlTTlS7IjbewzPuZoWd43R40WyjPl1sFC
Dy4D3B7KXSTiMkL2EZitfEr1IYfWVUltEoaCDPoFddIPatdcbVlz65M0JcifjEBw
G41gunuZrxucfvsA3deGPyhQq3XXvEWqt1F+xumrJbbvGrbLgYRNJ/ttiPwsBKAC
kqP9rKpzcVwxhNjLSIZFOIk1PYY/jBehjCs/K5MT7AT5CNYwmR7+DGO3j6VOZQ0s
MnsFR2It0Dt+Yc6I9shXJ/wHMykDWqCdgfKjatt5VAcvgPVhvCz0K/Yre3r9Sw2G
FXWMCJtvhPBfO++fsgNx0kRFIRHDenvSVgwxAflibLpR3uQGt/kXTh9SzZ2V0S9n
jFD9oVdYSGvD+w/sT2vKMw7dSbv6xr6DyYk6P+BRW66O4tFO01/s07fZ2uyBXNLj
4U1lSN0XEJzdT8D/TAnJybhykTmDLSPSZ5PiNUk79mv89y3I7he2ReyW+QRq5xXt
o/N3fzZOqZWjgqfESzmFsJgjwIeYAUiSY+cubxS/DWgvofdqlVCFdX16tcQJ8rHE
/EOlnezQJEG8kFCqnPBP2lupgAbzpdeN515W09iFXQsMRMJxTR4q4kvI/6APru6n
/i23002Dta4QbjayecRPcIpYOzNXchRtolnqdR/lqkMZMNVrzzooORdlSVHHT4RI
9+X5c3UwnMGlT2e/DwBmbn5qtUeaE2BLL4uhiEiBXW5kZwOivJMdlRJGM/hJVRSs
1T/NW/so42YtuVWvGX67g/+IQMRjVlMBS9GFEiNxqlkRgRj5Zmyc+9fvi2LBaFnv
/kVGwznbkuIQT6G/xD3N8s6gVVkqUZk6avEfFKfdU03KjLeEW25x13zeHmdi/yju
XjJzsRXSRGZTIa5YqO92qtRC31GjZzukYQ0dk6YT6sGtutkN+2lKigKI7RCcK5FJ
/02ZpcRIYZIgB+RmwyHa601lGPLusbm3uwo1G5fLBfYBSYQd0IhITjDrmHaZzzRT
ncqIHK6kFuhn8Zl3XB6lqlvfcFWBhDoiGd00iNyQGKgbPsDlFO3+ypO8xL6F49yS
80j9jBf+12wgfPA0x/TU1eOsOCjVjEaq2wxBOisG3vDfqTMNjNlpndLJQWOXSGcV
zz9c/1adu7v6iqH8e+gE0Fy461qExfM2rOvptfUJMylK3Lj71UeO+qMfUG9o9gUR
hriBpiVOHKddjZhrpiwZzy79au0LMge+PLWcK94V8MYfMM6uQTap9AZq+/dCimqN
Tzk0+CfTkCITpVeDt6QugiISwSO4TA4FeTf9GYVEMW82FCCtbgbglS+KBD20wsmH
q27td2/hRrAotSQE5vTTTey1RX7/o8nHEbr4DS4PDwrL3Bn2gLUGyUzDvqdbHGo8
Ydwmmbwbg9Hlusl7gKkrQuFaFDN2a5CXhM/9z4EFSIMPpqhO79ppLo+cZg4zJ7NS
azkVA1q4TNAc5uB2rjEJwNl9Lqe6y4q2zshw5dHOzDAn5L7XsTPszPssDzUvhuNL
/RyAF8DSzVNSeYePt4cqfapEtbumgLrEBB6BJY00hLzPqOG+CkOcddH+4ZGtRON7
8OS3TYU6x/wupXntpmJ3dW+bS/fy9M1Onb8T3/LGYX6/8BF0P4szKYcb+AgkiT64
CNToj9f7oB76WnmfIhM1E0fdsN0W11/TlvnO3rLOowlqucGHhMFMehyvMh53T5TB
PKMzr4z2LmF/d7MNTdpI90NDTzcvaNRzdZs/eFVOBa5idLIkKUx+awL1IFBjkTs5
WlVF6hL3WGshn8+uOgzLMmZ/WyX1VPQduXYkio/vS48tnyk8NmpAapJdU+nCwKg/
hxbA/htwhw+ooKpgW9oUlz01YWw40DgRTQOVjhcsh7JpgNGO+MgV/T7vyNhCKBoJ
IR+xcORfO1+y+t4OlI+B3xXv2Wf63nkx9PqSWRKCO0YvGFyxPl6dbEYKNsEr99tN
7H4twM5W7a6yyC8fHt/JRI9cK4fo08mwa/s2CvszTxroxv5PrOeg1IzgK8UTgl0T
YUGZzd1BkGB48+CzokF2TLn11yQ3cHNwl0x2vMV9lRrRKAhWD2DUtffNXdzaGdK+
cUfuuDxneJCQNbb6rft/Km9pSs/z9qoY9Prtlnk6zjyeGYEiy8Z+WeM89d+JUqrX
i05/+zBxnpY+sio0c4iXnJyel4l4GZbpkH/sd5wHpzaaa0i4BmYa9YLshxsR+GWe
9nEZ5iq8W9i6104+MXvn7P+gQpMtZT0ygVDsySU32BvduVLD4X5yfulMUi/m6cpC
Iyy9I/g2SDhbRAozpGpMfHpGwFx8LWjcTBDhx/IvsvWZuAM49xDPz5LP/XNJ2EHV
lSocgwHkxzCBWuqJhtciU86zTTNj6r8LpeGEfYlGyYyt6W6Sba7wW4G9bUcRzWzy
EKfF32DTbzRlQiAiGL/GJyYstU3XDyX6SjfxdFtpVtTGa3+F88JTSaa9jGfmI876
/zc9KaPX6/Lf8woWo6dFY+hnNdVuIVJYDv5SEUka1olXy1NJBoPx9OnwNNwfOng8
GpgnTp+cXOZh7WgHJLUhxTn2NtzxLt6VP/3dwg3WvXF4PT33ciuisUN7RQWg60Qq
R6gyVM1mZOjAa83i9ItolnmB8ITZ/oz5CHE9hIXWtHkRJVN4JxrcjfEa29MTaZpX
LGmaIdODG7lokXGmqu6/c2FM8ySmvPWGo0gdhao8XUThxGs5lTPyMkCULszTsJB0
AC7ZjShFqsLtk0o3tFJCFNxdIJyY4nJ5Ibm3kF+DVEY1D64TF2ENQdK64eBAa0Dr
3Z56aYFRA+j+K4tHyxrPGpWLksc1+eInLKU2EMDEchM6BFIf7v6TfYgXSD2qkC2a
V+pI62yZZfoTXr0EhCJpRZDIabCCrVnDexCJkGHNzKKNCXpFDOVCSyrY0lmdD7hF
KwY8l0GTkTrD34/nRMtRnPeHxZnmGilRN+sgFzHWp7QboVsYVh74v+R56dtZEvAQ
uMJ4ckZJZt/BHlcB3iTqkzo1cbiiKcU/EqFXZ93QZ3lQIrhgMgd2bTg7MB1mbGAB
AgFZ+qhkOzJcF1nqz+OkH70g/QHhD2HE95BjXtngxzj7wZODdbhjt18AaFt6IUqv
V2+B5UAmp00fatzmbGj4xWoWUAiZ0faO7xZU5o5eNjyQBvGF7egj5bZnkcYyKpc0
1cKCnKOFYcJYSQPfy7eSHdYV8ommfRA+W+chlgzcku04WpUAQqHQ7YoVuN3/3MW9
x16lMQoloDmdscQTOCxl27xW8rQnfNLSSYYo9WS65VenF0f1x8k65Lfk9Mwnvxyk
2hObH7pGGyxPciXCG9DllS4HLEIM2Jv+n1q0a+rsTPforu6XUIUt4JIhV4vcMJfE
+WjITJRylTG3+jG5PM/e47/XB5Awn+18XxstbfYsgsbSm8O6s4L9kl0ueU4NSKel
6JuEA43sPuCIutbYXxzgtmUcLzfuwv28yGrfAUMHYRRP3j1xaOiZWKdW5OYrg55h
kdiU9gyJw4cxirAvR2657v0/4is+WWw5mpXcfv4Tnbdu1ouZZfkL3vGf8NEd/UbL
TVtYskvmCsmYPJP3L5YrRel2+ZaG7dyUmJ/WzZuKyXRRb4y01f6FC6E747SnnHsw
+vBB3u3zZJKtwyvVUdkmzSHtPIBZrBGX1J6u/1b0GNf2Vo5IKvEDG2b4Q1ILk3lk
+Y8PtRTh4nLdzA0e+EUX7z1zasjubELm5JmPqgSzemKC0XMjA1+LSYJkxkYmLjG/
JAs1mTYyuvZVP8AYRZ4kuoNughXu8owcRlJazRuR35yZShkYZWmj9yyjIcsKIxbY
RRqrwNDyPyPDT/z4/gvL03B/eb+OjCizs24kAyJpXKC6UL3tcXro7JM7/SHfFrzK
RFsh2LvHt5/CmRznwG7ArCiTv2yPohET7tQjWQpaJPpinyLLzJkoXHWUAKHvKROQ
Bc0ZNSfsYzXshTHq3elqMDtJVEVBlUUW6hziS/uA/Hg2f1RH4Gb6W9PvtXzMJjNO
8jwoSSzj028b3ZLFSGVxUdhJKV7n05PbRsxxo8UlvQCj6+6iO2Cq3HSyR1Y1++D3
V3x3p36CqNEEezTIW/RCG1qpfmZumO6SQ1IVJKPb6nzKNhbY4tyhBddmjiDFKwaJ
eCNaaWF/fahQO2Rt5Mu8OPl3QBLB/aBHMlWWKzblGJ2rcFiAnFkjMGJJA/lehDSI
G065E08p65K88m4o9dX/JQ2+0NRCsy/GChwTaxQ0Q8DL7duDZB8SL4bCA2umPZzg
xAUevv7M61QGRt6yaUxJscrqTHGtKHs8W87VCBp0upT7p+G+U5dcKNJ8NytX6ikq
s8Bd4beZ+mU3WINp3bGJpHCobAsfyetIwNtBpZL7Ztkvlx2w0ZtnGzbR7PmpdHki
OeHT5WJzTSD1FCTMc5BMSYlvpMMKjdrT7gjC9gjFgmrKkxu3YHQg1yt9riSsviKq
RKWUIxFxFHnp4zxr/1v8l9/K+oCf/qn5hp2rKqO5sVtPXWrNA3/lwE+IPFUN90oS
R1nSNPdMYX6PTAxvuJ9fe9bXIIcacaW/9bHfAuP6Btyrje28EJ4U11g9xpz8AP3+
34AKvICkbIhcH5ps8wQWdko77ggOSvz8VQCGs0au6S5BkbLKaA7/034ZNXJjvuZK
5cBukcS1yc02Aeu0PObF2a/AhSI2fvkNC2SxL5n5LNrNqkt7Kzs3TsLJ5eaU3fUe
v0/w7Tjp09NiMdQui0cmv8cEQwuUj/7Hg4fxoXiSyt9mdlrhMcreku7QDkPEpLmw
92Ha5RVOqJxNm/vddrocE927RltX0sR87wPdd6pcKxau2pVoJ7heglPfIkAp6vi/
G4u3olZo/0enVKHivouJ7Nk+MEaZaVFmJaraPSvQlPbBCPILVFP1wHto6dz9W4IX
sbEDRtYpwm97sugB7jp6U5inrv9mlu9R4QkHXY9rxJlZHpD0/+3UYDYaYPwgIo2I
57ZPXp+VuRumvUpx0gW8zTfBpcGRRUDSVjUEPFRdhHRb9xPDO+RgLXYQ5/vf1OPG
r9w0oEZkHUnkXsV8iiy8SWdFqKxlTkj0a6OK62iXKqS5ZH1qi6uHwZKmiLlLSYgd
ucRczNOcZCvjYSFRqcH3bCfVRcsQte7ldJPTG1FVK/g6Io5hEovFvNPis/8j/sud
J3k7STS06AIaPQgWabbDkpUBgH8VKUnc7n0Fv5IjKbHh/4RmRNfqHU47UA8tLniC
gbabnx84tgfd79jAf/rScFYITWhV/kmyHejCYEFfuUI2rJ1FNw3jC36fV3Af1tvp
b4Vq5ed0MH9dl+alYUg1WEifYbTGe90aY1BGZ8bG6h6592m9BTZUYIIzsbtb4+yz
kp6o4eDL1L7plMwgsZAmo2eL+nZ2FqsjZOyWu4bJvSg44qlZkaT2CI5p6l7celsE
irA8UgtURSsdVj2TODIG6N3PnF4WjB8lbYQaKT1/Xy8xEWYlEhBn2p0bdUaRqzYB
m2i2ghhq6yJ48ZTqAj08FlYQaFvbAq56xJ7PCdhOaZW4W1knXH79t0YRqqDl3iJY
eZV8inen30OxHBtXtLQ8OZyK6EOJaXSKpZkKnPqzgdiX/63h4DUEQhpa/3WJYeGv
fSvJ9JoR7H7kP3PBwtXWhc+cGT2nStdnH+RsIYDFMBEUunGMjM1Hy8cHINiE1dd6
n1+ZAeO4uxgOcwembpoIvfR6sffGYINrX8maxQFMfH9QCUsCIbuuLtuNhx2tUez3
DwgWzg0cqW1QtvCQGsr5h8aiU3SROsGy9EoUcomZcs3oLS33o66DdE1MVaMN0UQa
9LrUrnmrAoKdUFAVqT1EuWGZpAnWLy2lXmG+2Na/0QSOuWXKjAsRRh3OoFYvFH8k
r6rV7UCH1yZt/M2yl+VP10muX+paa1Sz8Y+i1jTDMR6gchCzGvBIB32/4pmo6QSJ
uJcTPDt9PlqejUMOMhifJk6ypoRmL1dhF4RNzb9NPksbEIctLA0PpKNeXCIjav9G
fjzsMEYes/cCLdowfu3WdOzzmH6JixhQGXV4RBSyuZfWnDxhOWL1hUWqdYiqF5/d
884Zi1AAn6D7bxnVLYqRzYAn07sHqcSSy1Gs44OmXTABD1jS6JaOYO6V7SAEp1Q0
E0h7q18iFXS77gFFF1N1S2n4MtipYOYWkvNUTaNXBg1rhPKGMRmVURebbvHVCY5J
whjwGG+DHfemDPaPa6MC8/dk5RnV+xX+skKvgiXHaU1vMK15ITJ9lRRy75BF/woY
tdJJH6gr56cd7l5/VaG0izc/fvToPVy0yrvs+5cX7d5LdqOPPW2+h73C9/OhBAB5
uyorg6pKMtKluuN8NFhvqRBqFTWo8nIPsa5dakvikn3Sgr6ync9mjIJgYXkxQ88z
JAkeU1up+iAet+GyQYxVMmPHWfFWqrtongg8jPyTRa8h3w4DL34xTUVCZ79N0zy6
kCkvVJ0lsj5LRgiKpEDnJG7dG1m05ry9zuiRtDgz2jR2znclskEYg9ZcHYnqFxZQ
GxY+uP9NU5Mp5yk8TVeqVssYR6Rkl98LHKned2+jJpmcYVQdLYF2kWzMjkbn3zLk
We7Rx4Lf1CJb6tBqqOmKuzXQbBY3RzW2fcQfv14+qjWWBmi/WlvkkSaJzyNe4DXl
euaKrxFUzc3u9cuZTWWFgcjS7ZmiOPxUnF/nmYXzuIXFxOXYSIxzuUJdL9az4tZ7
k+QiXEAtcuBWHYm5Iiepv8F4GIx4QMOBYXjkQAhDoLNgYC8O4rtl1m54ogWpUHcf
wY+gJ3arjws4GxwsxA7IL07qCZdz7sUUVf/uEi+/Xvaeq1fFhiRs231Lri3i/rIM
GDrFOBC/kAb+pV+7ldIbVXHp0uOmHOuSplLn+mOtT8pTtYn1e/Uaw2kWmNy8nUNl
52Zeoct4knt8w4pE222UB0f2ExifwAlJOZa9iibiwjofqpZJ/C9LKJdfEi+bpS3a
XCUAH03ngHsLhAo0MCFYQ1Le6kpYcAikC95eePnmMD1y9kKPSH/OiJKgPj4oCCPF
zHKB2KprqRt+TcjKVCk7D5gj3X4CJ7PYeq7bnVT4i3DREyi4y4H2Jzu7UXaZ4/ge
/4iRPh1ppBR1I/5t6HxTRV07pfosRrkGNhXoRrFGS8BvOKk3ZKHTqEeSbScfE3sB
dsKi3bPahZEyV7ZvurrZRgTVNbZiUj6i4DIXQRvfIJ0yzmSebpZE+rCkZrd9eEpx
v1VySHnpirJqToBhLQXgVRnxIUWAN85SthjXq0pBKuqNgQmskp01Hr2gqPvMqkx3
4quDTRs84t/GLyeju3Xw+SkGXB9txH40d8nbsuO5Ak6aGPgusUXFFSGh912x5Jpz
UcOntnrJ8KiviMiERpBYMbPYQoqxYkpcCFK9IpmXo/NkDnAQO0EFFIVfSq6vdje8
MZfdZpcv1ICpgxhb7mQCdTAGixCYqHAqM/VSR1m5NBz0Gt/BAeHcKQdTN1dSE5+i
xk890UWhJeTCYTtACd9Apcxu2dtW6YZb3jb0dBv764mKllBWPvdtylFn2JW84Hht
XIUbMUDLpOd7ryxSF99Ocpg7gXyPBqLn426DKqr373ks2eWvi3nR1og8qMbhB8gv
wzZGeLHr/SGPU5EkRoRsmxzLTUE+bvp5owE6+MezoolnV4fhc7c+zjRntr369WOZ
JHHTFsZa7NYpOzkGKWHAdjYNu6nPd4Xk81j5q/CUQ62WpZRxYcRCSBYtCChWg99N
WZFr31yGXrM9HhB04ghTTShUeHxOlbtU2pG+DDhUBG6x8+QTO3F/NIw8qrK/4kbY
QVOFkCaUpKi+0OqstWw9WRNsLPxghj5KEradfPAxq2NU98kkq4R08dslB7zl2qgj
xeQ8917fEC8OTzlIzeWXPb6yT8tJvwNTf7sJQoAD+Ju0diJx8YcLtmZYp1NHVtFY
9D2h2dAsryg7sIDtDuq7VhzPp4S8dzIJgo5lJnaZ48V8QD7oadNjOYiWcDsyw3he
8Qt1PcciZXtAOEQPrd3BWoVyvfM3qwo3Mr9AtN2968EeYaTSLC/W7f1mc4IO6Kwu
oMW8GkvRupLGPu3UPUJSNjPX9IyBq0nQdF3i/0RfOltIQx4L1K/nbNEi9Jm0jaoi
dkFNKBYVAuOM1J0URwbwFIik2w6t6BdVzRaDsHXROp6pn5qL+JWlPvtEfnUSGI3m
qpTHrUkFMSPLDuAZm/EEYQ/TEPkXDDGcvCV4daTfuKiurFEreKaTle8m34eq2c5Q
fAOKLio6SYaZnkPPZOldvdIRzSB6RXjJT7tslgMpVYPu0bN1PrMCePwjXBcr4kUb
5rsm4a6SiQVxB5OMqHuHQfbGwSngw/THt4yoUGSSCcEIOtwffR1xcI7ydGND3ZfT
T9cEpjde8H6EjquHE/AK6r0gBx7hKp/Syj7T3yegBmcQdgZQX2jdsgcYQekZUGNo
gIfNKbEh+TyHaXfKBFFKqDQMJSOMlhDnsbS2YnQbHamnBwmfFBB7vRDQPIQt/XNc
S6mCH3cv1lCP3tFWm1JPquTTnRVm/0ep/NjSbGZ8X3urBeJjg/SopKKLoSpyk+br
lVf5fMHcF7bBBex9/D4GWCQEcw2bsXVF1IvvFoKAFz3dtrNYo2fLD/ubA6IcnXfq
vfc0+Phdjs9E4yRtTUx9Z/8DSILEjGkvBXgHy4NKMfWbcszqWklSTYg5vOgUC1Hm
JsgaPRY5BCPcJ73eJBle+/CTwB80cc95HVWI6aFN1I1Wl2zhidjYuhAmzMLhmei3
/m1QG+CWKBZaVGkaqa2w6kuMW1duYeavEktRbXOtpuxNlPGCnzf33GX6ouhz4a7q
6vBg38ahU46Iy+Lr7dyxFJ0QiQgn+osRIKeHtdsrjzFvfNijPd5kPIJk5QhqL8dg
QDQFq/lCTNHeftX2KMVNxIDOhWwEZ3pv9TTFxE/PASwNHCFYX4erk0aUIyoX/ewm
Fw+TaKOSAeQehT5TDDSY0B69UUHBkZbmiqiCtBxqTilR3fXG1Su1GfH0TIfwIJ0I
5y+aywQdSne4o0k4rP2u8qAPZrVlnhY/STvXnKsuKDb1yAGkNC8X/jbj9mLCHeji
HgK9x65okTsCTrXhisS1QOmIC5N6qTsVlpKkYYerVzT1BCsEnAYcbymCTEY+0Pk+
v1q9tDOF6KIQOKtCwSNsPrEAoCYh2cW3uycill3yEMupF/30c/zpgswDzeqJhHuT
SsVdDX1aG4DyQ1OqBcg+MleJoRZcZa3oearczDHLgv08oid6Vm3S2IglHsAbO+bx
+Ayw/4cc58ScMxGXAaZUlL0+mi6sK755k4sdcXI4BeoFVd+4vrDdndp/k7UKM2y+
VZCUH3D39rdt+Ti6vu2B628j3swWuXmj8NEl/UC+AlPoG/DXnxA3mOpmTYJrQRO4
Ox/MsCxuUo61ycrJPXObXrd6/mEo1tn8qWkYkqZk28Lteu0uzTBlPSvNj3NBVidO
Km8rX4AphRXPxOhoXemvliKMAdTRShNEnRJhzlm0kSe7ZkfyOQA2OaafiTc0CIu7
IL00yw2dOKVjDaWeUaTvQvvVeqAgodSAgSpUQAKa+7Pmblyy/TjFBNl6YAxVdF1U
z/fvwH1oNy14nE+emF9Cb2D68RbjARzO1mkvh8mTQfoM3OssqK00PxiqtztSmUDG
dD8kKFMFF8ZkBNfxCP0uFjhXyOaFol92rjtcs2m3gB9hf6NwO2J1Ss/KElAX9F6l
89q6QI95kAfrAVgylaU17TExm4zPVTO5YHh1O0gsBWsM8VVQdmFjS9zXh0G2Ru2S
OMHKTgmDwasLtksip2awEzqdTtvGPTF6GIkADmRsIUoYcfOmzwwCn4uk/I43zveY
X5txOsZfe7DtKprVpq5OKpl2yfr3w8EJEeA1Ni0R05gEOrLvmiqt8gjy+qng1hSs
KFLHAPyh2l7VTK8Ujs7PqUeaSmc8Sju9JTxM6H9Z+baN+jiDAyOPaPt1xSHMHt4I
cNXr7/BQ2wMCe/42vRx34o5/jQ88RMQPTh9nO9ie+ZlK/9JB9DmwriVKX7TNpim1
anhks95QT8qktiyT8A+7SXg295aeA87UiYw6M4rWQfIyBriauEC3HNdR+pDzm3q7
4151d9XnQKNsRO5PynE4UPRwIBqyaRO02gaIv+tXHTtpY+Ew70J9tFMvJdJ8Kb+O
wWGVJ7Fspra+xsVYjcBQF8lKeKcWgliXGMYtIHyw79IqBo8VzhFxQjvn93RDHFyq
HT4DYUqo0QFCn/itlnQEoBME1ciAHUs/wzgDXRC05Vz2dL/z/aHL1W8YnMnF4jYv
O7hOmEXQHV9aU8c7/Im5T/B14tLpvZvpXZf8JUFobOMSHPkc9jiPKSHYr2BG5uiu
oc4Q8UrZlkZ9G6d9fyLDQuZCb4Ld0d7GCCXldy5FrqRnNL9IqHHS2mb77y0xb87Y
B5148fMXw3HGqTn3KIraEXqhcP0VRaKWnBinbvu7B20FzTYgvsWVm5hVPZugP2ya
se8lF4bqlsR69yqV4NVcH3fkCDbY6snwYgKhBAC2rVHqjw1GK/amcQzR6wwMeDbZ
jYbW2a20fumsjr119dCyWM6MghWC+L4Be86+F2pRIPfmGx08FPYNS7/JVcPNh/yz
yLQf/PWRpt+c0gSzVxk3ZfoXk0dEv1R5WbGDxqEr+I0j6btRFbDEZ3PegWojwTID
zaS3/NhXBMPRPCaqcrGYd9VR/oY18/sDBgTkIT+xwqXhR897+1PIUHA4uJKSZy3O
S6KZhrcqzh+KFL0dZYvFkCQiQLd7PNh5WHnatuzAq4wvXqdQv3z/7w6ENdh7XlsV
lPfLfvUdRrnfstvm5SChf1leehG9zyZUexgZJf97qZsR7e3QZv+aKz/N0B5RU3iG
WghOg/Ky3M2aVLP7R24VZMRig8RuLXBKNn6VgdsuLscctOw4lCaIlCzhFd8blK7I
EV/08UzMjPvEaoxjhYOTPr0WBA8esuBdaw96NBymaAxBtk7uOkeMmAteiTeBJLJL
0/6bDiMfT4SxxkA8jfukqnJVMlqZjRnwg7r8uLAmvSFIU3vt0UOBvGOmV6N22D5e
+9uThRJ33aiPu6+/rlxvh5D3JIQiDNtM6GD2w2tLc2o4CK0hmngy1n6EI4NTjh+h
kxzQAkGZT942C64NRY7/mOalO5JAIhlXQJBx1yKkOfQEAo7XZfo57MvIUdCoZlQl
8/NO5Ps84MbMGk/fuZjF+pUCa3eONvjTv76QCVWJxav5slSpZlD9Gk9I2p0ldHV3
0Tm/Inf3wBGjqRf+DrRODU7CVAtVmua1YRzbVkf76NjQauPPaW6okFYiMXBuc914
iqlyqpjDzaerf463AEZt/WDKgMnZDeT8yNW2oeQ/gzsPBpQ7gMs5IImNh9ki2paa
jf4pHWHvmX3ow5g14SJxyQqQ/Pl81G/aqPWeR2aoxdm6lHe2cR2k/tBFt2BZ8l79
ZghoccbUxE6xvveRYpHsfW81UNUmBvhJ3BbpsjEQ37+csqKktSeit7X1RDA1onjC
wAErFV/L4+dVouOZr+1Ou5cWGjfMGErXKuj7Y3d7pxjMwTUsEZHkNbTX6rHKjnpp
1pHv+V21yVtR64Boebf4Ih7waOuo36EV/qji8rPdBUbm9lI4vjjowHpDTl7pbsRi
b+C+wta9xqnxEA59GbmjH93wgnpp3gVjc2dow6wDkAUGOu4EggSpkQZxyIic3kTH
sAbTTydPf2hfWb6sCXUfuJur8WFT65Wwhf+Vyy7hWWZGiSep+s99C0MnBUB1myrZ
EKu1rq7qGPlERp7M0wydYymhgmjzlAI5WPWv4QMaYnPcG3axgr3Zt/JVc5MZ8Gc5
lwwshKYWM0O7qSQmhn9AxK0pClo2Ks4S4ullbIEqRoFpHCNEOxhsmLh/3oJGIcZ6
3F4Co/muSlTM+nB8a2G5dGBpu1UyzLaFy2WnnIdqc9WZk61jQi/vTeMDETJ/ndnd
dEqIaUiFCVKpcsBOyVd5j5YzT5pJ07AS7+3uHuzBAwAEXR5fM/E2JJJXMOMsEhg4
Q6+3LRmrL/fwcvAgZyQ5yvPll5Aews76OJ+OQLc+TVgENQx+OCi3/ljYl0nLmTEw
5pj6/8Er3RDQXixEgwvYuO3HZ7Ylq0+LdzF1aRPrtQN6feF96unGe84x31TceNQ6
Gap/eCfF0xqz/nyzpYiP80fjytWquVOe9C7gl4u8VVnRTINULMC9BKgTeZLTHbTw
qa95ifjR+rPZioTMJb0BBxCZQDm9IUMcjungoYjTUwoBk8qwLKWbmN3vU1X8K6AN
R9zOBZEdK5HqwXmvBciQ5Nx7f0HikQpOnzP3Of5RCHAK3M/FO06DMP4XaMapuCR9
Q1bdluqwOI5uhep4Ggu03HKSXpMq9kDA0jalbtfuYaf3DFwWspXp0NYdDmwkKsMp
DeXjtAH4HT6vZw0r9S2XNmjt80C5Vjcis/s3f1Em54hinBkA6CG/ebPWuUUnO4WT
clRdAiEKZ9tT015ph6uSLN0ff2Mghex6A5z/QAbFCqayT/tfsqQ7B9Rqt3SqRbsk
kE6ATRmg85/g53BRCSadt+bouhzTftT8aRgnBktzq2cjJOU1AZnARP3WdohU1tSW
2kFb1pQDVsA6MpYQN1htVSBqkdL9SuQzMNCQBrYX9upu/3Q3dwIxMcfisVH+gvYM
o+0ZGHsr4FIgZyRuQWd8EGDqaWAIJWCZmroxf9PlDVny91amzMcTAgxTp6r95/Jk
cQJKlyqTuZm/EXXKxaH04XDLY+KNzIBt0T/HxfKgegq509u5V2FNrd+u/lf1G8h1
2aGXniNeSay6/mdRoNbYPbciOxv31xb2m5CpWpWjUfPVQrmBUUvme4WgDU9ZO6ra
WsjzQHBUFLn7PBFpkRpoAyzXPIvMkOslK7GRebVhDpKJlGjyalJxep1pTGq4xttI
sC7B5pEwfVKzDRq2nnh6LdJPZelXgbOcppuuOMqIsuIO+3Wt9vyRkppftzp4nCwd
RuqS/7QB/cmWWScpG5M1zLziNdxiiqOMI9+rbi/7zFkYt5LF2ZESZ0ziNO2tCBV8
kUpAxt7cYquHjPeuZHiIGyaPzw9BhGPNWCGMwAsKDN+iyjTqVWQxx/7a88S9XEtd
VLLxxDsbGRN4E8NF6vJfHa910q5rahuYCSW9FdPB3aTUkbYH1+NEITxt3wLZZetW
Fz1+R5xZzAhqVHFxL80mus/TCX0j/Nn1vXBQPg4rHBIhOSZnpFZdaGSwC4n00fR9
B4/SwUFkvYXdAW/YLSc0ifgv0CbWiv/mx7Iick/eRcnVbzuwc4UPhjcxMxatVaf9
4uKRXfhNRd26ue5o5Blz15rUq73zWHSP3LoAZpf8mpJ51GNknOwDpF7n3x2nCxMm
V7/XAPErhhojLcQ4Nz2eGsp9Os7j7KjUuwiuz+SDZ9DmX9X9lb36AFcGZAZU6lBD
6RahASXp5WXb+nis6sob0fvebzYOkEuMD5NVjnjPVIo8DanxbAeVm5lM8adR8Ahb
6m7xJfGvql3NDqlitlLe8aOOwPTvA67mc35a89fk048HjAc8sMaIzUF53OzKSvpu
VsE3pQaUL2GU+DVcJercWW4zs896m4+xeJvDYTypdPNSvi/wHVcmn0trwKe9bazj
5+0Z+1Mjd+GDI526v/9jAV7h4x425e5EbJNt38DBpbryK4OKF6jlinLkMY5GLQIX
qsUygF7xSL40ShzBFd32R4/eJbd2SsmJJ/Gcsu56SkWLj2XL8TYmMLyO9YDw/aGM
DLQiV6eA1D2sOnw4Eju+f+s28JLEwrpobkjjYaihfsdDHcp6mDjJvbLOFYfB+u6I
vIOHAyeTksA8vc8vVp0h8wQeDHSlMuDr0rUatY2ei3qEHFikrAqFahcAzrkWVhWJ
0dWe1OCkV/DTubnL1Twxom/377tfsxrVO1tdwj8wnOXje7d8nj8O5doFxE5oJL3K
zJA8Xe0HHVyokFYnLEQ1QQZWRPxBloptLvz50hRLbtqFW0KjgEhL8jV6mvficwTC
mJ5TWNsjsQJZ45Wwv7pSop02MBQIQngnclVPg+g0F/Z/lOO8ljqTOpQWhMcync7W
pOvuAaYHbiDJMXOrex4pDzjbugbMblUpzV11lBPoQy77I/prbrgwY4ZW7bxLWt2T
dHLyfTVazeHqR75ZztgnHDeXI/uWRmUWrekdv6DjseY9l0WU45//IDn4XyjUbg+O
2xyR4dTy48fcyVhD54/+Gejm7WW9+yLfvaeTlk6LoijlQOJfNBGRaFRL5E+g3ZPd
6ZEfJo+y2M0F8CVI1sxhVrHVeWrLRdjtEadwGwHbiuv98YNyHTykmTnY+i2TFD8Z
JsCeJ/OJMOIT61Y7yDwVt7/MXZXcsxriskkZgGnesBgdSKoLSpBdYoDTyBhbWeov
U+1pedhNM8AwwQ7AgTNxosWeWs8E/36S3ACnsRetI3D9N4/VYcgdu8eKQGVqt+pi
HY0iPRM99P4Z9g6J6k69hM5Yuw9celfkTw+2IoOLUowu/Cp4hJaN8Jg0v/sek8m8
gJxYEoAKH1ltOQO2zhFaOXwolHCN79Mdeh7Mtxs2c9RegSP6kqdGnroZJMGnFKqi
fT6vlh0Y5NkGzebERii427JpC1eGDxeBe3tMyHb0zZgSUN8Rm2TRZ7ImbCE2TMBN
YAx/tqjzOBze0nziGnm+9BWP+1lTUMHgd+nW4D1csOZO3vE8BOoIXovojQDRCsyB
A8A7hBTES33KIeAoYkzzU2rZzoYiDnoDw1UsFFzKW2CYtwBUE43Oa1lv59X1ByiV
qeoxVMjJ2GYQkf68rlNjzN4zimCOzKaV2XihpHr8BPb/9wOuhypzExHlqdwMiw6D
5VhXuOTdK2AYkargSQkN5C7PC9HApyCsK9fAWDsY0gSjAutimzlwkYBbOHPJD8UC
dZqD0ODqOrh3OWpezlmVa7rDD7Was0BrkWsbq+dZ/K5rfblBcMXvZT4UmyzGOyB0
2rR59aHnonAUto7YB5YZOBoUQ9Y/P+WdYIGLXaeZ9x4hCgEsnxS4Kdup1eshfSLu
s+sR1Al099JjKfrarGJ8tLXnvtqG2my8l5VM7r59Ermt//VB8bmyJYrm5SA7G01t
vMsD82fbH9XG2Ly/Hbry79LC0EaXRDjnEDw6pbOQuAdvmKaJz6CaGpgLiCIGX8bR
+XsheJLDC+DPq6h1LJBdTJdW1QbxsSoakG97winvNy740YO6d6OilLjCRiA7NxUP
shGv5Mnl6mg41NknlNSn6N+KB/oTV9C4UHwJYAwsrWcoTsFjMIl0Lj1r4i/LNGGv
+x5d86KeAwnFQsd564vkQEKNhAEr4Gf9IXIfASSKTxm6UtcDb3RKlcn35BqINvsa
b4MI3+k6zDq67L848UTBPp+XqX9st/+lMcHJzJREHoFLYVvziTK0Trpbyk3L1P+x
VSfVFC7TQakWqPLKQjZ/5n2yq3tAcvo0qvkABOqJ+41x7fGmzNSP2RU40uwx2ekD
4j2iIJlF6UOtRjMXczH2S0sy4zetuD0fg7EBJgTYpu8nDATv7NlqPrbdU1yqTLZx
+hEOyRSmpb/nvHLhbgluJXofPPaKas01rXPZDxbb7NnfPVrDBOZRnx/une/EFvIx
DfOErj0//ivwUYZX1prV99xpzqRvg/2JIykLPdgsbrfy/qv29PB345TrYboAgEoK
oSUFMqjAnfhVkPjVpengAg41gMkCh1BPvKpvMvNHPE36gRFfZ+WoJWg7dCexGISc
h7lGaKky3a5+T34/ZVaEjGUPxPQvA7V8AckWN8h7l8ZS+Y9d/+gkJCu9oYLgnzJ5
oBUFlwuuQYqohd4yg7/DdSAz7u0n2L/1ypY2NJDArGpMyN4V6B3zvgqSN4UTh6/t
vRyoWlotvEvLCng6ZDfmRcgIY556appZwlIrzKkBW5/Ss4uzS+9sJRu4S/18PQQl
WVDrnJ/NAlUMju0kNHo9HfP0nXfzsiPB8GP1jqO4UnpBCc1MM9R0KTV2A39gVLGT
2kyJeld7xYcF+5xds3Z+DJDKmglMpTE29YedZT7/viCTTYGgF7RGFo3fl0fCDSK0
duSfOq8l8ApHWxRTTHAgOj0iShxv4GlB+YZUE1HIjh6kS0tJNN+8eSuZ7ICZnvuD
ezTVdC9nqwTXPaTPbLQdBKPF4BWKDcAWHS/GX57YTufgSUNANlKKLWX3jUb+gJT+
5kH/w7i8gOcflaM9mX8tCIfVZaflFipxEI7EGWqnUUpLy6J6bWawiY+Yelcp58Kg
j0RaQ0wOGDoYrxl6106b+a2ef1ATA18vHsGxI5l8nC26hTNpGg47OHM1RY5Ni5fZ
ianSIsRgm0C0FRvmgLTm10Fp2bTmS33Ha1SJEX+RArtwnRgTzF7zIC5pCg/5PwPP
TKI8kWCYt3lKvchtaQqAj9Oq6dDxcveVdJMC//ObDyMb220c416TLDWU60td3z/c
uD8wbdjfwoBs9Q1caSlqw1sx7HUbe3HpYjKNj3xV1KJxkEowgK7fcHI9k1jpFWIP
katspZqLhVzDrEhbPPYVyGSJdvxjrJgGyejk9fNT1EwJH77IU/5w0IRyYV2sEQ15
0grfRm2HDZiKeq0AwINXgSt9O0dxy2BLPu2KJVYx6pPIle2hqD5wChshQtY56gbX
1TxJ4Q+80qR2KBYJex/KlLaE3OnpVam+F2recvrD9dVCscWcM/4vHK90Nj7Fwy64
O1VwHYKkgrqx1Ijj4Y5sT6tszh6WSTSrppoH2+17z4u3JsBPzRVnAwIxxRdgwwiG
OKH+UcS5PkVsNgZWDfQaW45TrrPgkgJkk9XsUcblmJEIlyOjyW5XVdbtcHeNEv5O
L4eJBLFgIWMCf7Z6r5vlmh9o4We4jh3vM5Na6j1Ukbq7fXXNjvQBbzsZomql+dpd
g3v1BXFJNg+P/7LJ9FOCNeDuX4IAvlfYIN9V2d02fErMNzLpg+TMbemUJJ+1mv4k
7WlyefnWqtUfKujQL1YOBkF5OFH8EQhYGhtE7QRPzMtiT3w0M/hc0QXQuV31imay
fWMXKM/l05rwDEjzQ2eBXPL8m11YXCd+ILcHJgeYbY4rk6uR0tnU/L9J4+2HYotM
8Ca1RNGIagFNqBfuHp+75pfh9k3YP8mY/sPOfpVwXMeQ3+tNCiE327G69qLJP01k
mq0SPNC82G/eAzsZTsMmXtpyf6FQEo886aEQ9PeB402V3NfuzqAV/ISdm+/bN3n4
aEZgZ6vOtsVMoniyxgiD4fh4wNvBXTUTQAvrH0aZ9WZObJJg6IUOBAS8c5VK1jUo
NiGSyrNp7wfaQL4hCBerucvmtDqhCBKNnXcGflKRMAh3vxEw7XeEr4E0dZjuW+Ub
+iwD4sA0FGTiyZJpr+YDoctD0Q/2/S3QF3dmi4UVFkNWvJVzwwXXwy3JuALCcnGb
WAfFSb5k1JQAn3me863ekT2Wl3ShQUrfTNwOq+D6ELGQH5394+S8NwOm8eR9x2CX
w/XXSDN4ysl+rCqkX/Ut2a1huxZ9Kc63eCJVmXyex4qatrKt5baXkltvOHSI/G4b
97kzflxmp2B8Zz++GkJamU8EVveG2BvfidfrNGMUM1DpfsV2kj/kApIW+8k2ofpL
O0rAo9oNFeBxJwMx8uY4iZ3JxXspkcz5ZPlwUTtoS8m6z5PY1XBnJ/IvLc54K2+P
Th/Gl2HyofY77V7ZIE2dD+qWkVCdFsWRBXjcJwKAd45feVHlA+hoS+72I9AOHblq
aWmv9R4PEtfGzP4BFXXtoKi/WsDhp/STdpF0EPuQEC4icKPshyRmwo+S0G5HnwNq
1xpK3DhgT4RXS3mhllxKnuE36pUq3PNAjMPROF/A7ejGOxP3CSOeFcTXaOWvGxHR
0qqae8b/X11f3NkubyWK62GwO9skIePoHT/wXQrLznNhGUTCu42atSTPnXhYRxUe
JWZLtPUw0rGYmepvxfuGWABP4aqw+u060DdU/R5dQ2KGuN5atOD88K+YiIRMHFta
3vRbD9qp/iUcsyPnnQlVU5dkn0eT+6szvXs0cQOKxGzaoEJMueYrR+kmofYirF6o
W6te4bSEYo4APAjoJh4qeVKAIxHDOdvZuym28hEL3NMYriAF5z/kCrAQMykv9nb8
t5YIMt+x1A4Z5GETajZSX/AR4U2QfZsUDyqNI51IIhqRYGLvaRx5D3LhKfskrmi5
y4M5PRpIIgsq3AX/Vn7H9uHkixDO8wxB9RsX4QZNh7FsyM2uzwqZFNqeso9UyueT
/PhNxRIC8ixKucnb9zowTaRCSTa9cUW9roPabi01htUWfh9c2JXkgxbjKju8yQpr
oaHHY60vVH0WP2K+dFpa0VHXFHEyGF5C+CBb0NogrD3ojzF1sXkDpAfwf+Y0urhj
PVlKoAipQU016Rx9saBWfllkAD88i3tYfqBzDt5YmR6zvLxl7mEmjV+a69q6Weat
4jxqhFsT0/D94PiyraD0HyzXTS04RtxA1yNvZM9pe4siIMqWuSmT++/0oFm0GLek
HtiBNwq3sUgczvvITIhc9YA00kHlZZT3PO4pew7d0XGTUVmSwW3VfQVIzqC1pwpL
e01zgQ7lyqYPE7ADyUzACcSYMKz1LxkmiWFNUiDknFJaonm+o91Y8zgBrbvRSqbi
bknKJRUAYFpbx2eJ0LHWNcJr53OcqYJytgnRfuoScUaKrvNaCPrHatQdTe+HzyXB
Vn9rRPwBadqk1BLgIjs8DKG/smsXUAQ/wYd3IC+kHBQaHjlEvv1YGJU1NmLvWgn2
H3KMfGQ6DPg0yr6L2J0JeayvN9KJqhrtQ+LoCbIeXjp40M72K+Yjhi+hXir8mmi4
rB2eOrATsVqZNdD5DKou+MhkDtJqarpXsBko7XmWs240U8mX9RalEcINhYbf3sjA
9B65E6lzLsb7PdLVz8Da+Mh6KuSsCXwpW+61B8HzEGoRzdpSwWO6DkmKUnhcwVGE
3Aiehzrp3vSIFuxvk47j8DaNYTaHbA3A56vcm6MFagTFjttx0f4qUjjsbKT2VCC3
B3+ZL8pvef8FMVD4nHBPCBGUoi+dlDa4WXb6zW/qqEOAAF1CerxT10fdBlrxY8+P
+QMWX2WuFDbb37PmtdnoOCKSfsbNMZXeW2a2CxL7oPMMdoXGq/Z8xl3kFgnkV/sC
Aq2Y1aIevJbYYRBNTjmitE0DAQfPRh/T9NGEdG95SMIzH8w8Kct2dSWZnZFkvoTs
M+pOYnPoKrHaLGNGdPsurR6PED6h50ePclNqQ9baDZz5RSXSHY+H7W8FB+MjO0Mv
Uz0tkBtA8/asOmIJYBzCxsbYuYXGu25Ul+ZhGbed69/h9TJ1+fumsffNFNFeuR7p
QwZ/TsMpf1dCTWscwQrzmx9tzr2GcQzcG8rBR9tBRahU2zhylG+Z+kb7HfU5Uq1o
ljkJS2jkkSEe3QaG1dFdxjIPDwh0/VwSIbjfhmrGd+R02cZYBSXxBCE57fbaBuoP
ffRaqaclJehaH34x5eAGEjB9fDPgj6JwWI0d2FN1NE2x/zLXYTUM+z0XwKQCzFz1
xGAnuavDij3RaJDomUVshB+2Jnlwp0ORXzTT3lshZzCdRXqSHZST07eR/S8V6be9
jX7UYTBf5ttaHsQi7jPMSIBVDUEnoZ+3jTEGDJoM0EhtMVg1L5GXfYzqxohUw/gk
50WT5qCN8KizVwGAjvw16QpQewKGBcRXw5l8s+2y3kCLafNG5oBwno/QpoUXNynl
paeStEy/JzsCqSxA4YReVtaaMQW9TSGXfUeS/K1HiCOrb7W6dHnEascIEJIwQpG1
mx+jqwtV7eXvvF2ADg0ZTQPSxQP+gpIQs9+IgKcSsexk7E042gWkffxiXW+hYsAG
pOYZnwyVTEm23oDPyvK77dF6rrOqbhGiqMV4bkW2z5kWSeGagREYtHbPV2hc12b0
G/O+KFB8YxAVIzC+T8+fwk5tiJw9ljTSC5+o4FxGaXMyd9cCZMrpkN5Xdn3aBjL6
t969m4EZ/KmCo2Kggmghr3o9MLzo9rrQVeFIfDEaxUljKg1ztX6MGgLJfnYUkXDB
KtLuOGG/xpSfI0Z/fesN9ug9J3k4JoqgXRvCVBJgaGuj/zZ3sfyg2rqLRwHEIh1T
6gF4D+icKsk1KEK8qbTeYUQILA1yBT+bOBTepykoIxv0y1l8pIRcW5gWIptEDmA2
AEkkZtARC9jYHpqM85uPmNMpm3ib2hRecJkLr4G1pj++3orLWsLR8l9cQ4uZT96v
Egz7PJ0/f2F3jUwrw1kY+lcbzn+er/aST1GzL1RCemFQCeSu3Wx/hyMFNltZRSci
7W1pCQZFIxn2ta3eTxe4n4XwZFnmyfp/zZfTR/80heeP2P4ny7qshiVea0a2SM7G
8QAhX98XYWubw60n/ZOmwy4XfnXNfb7E/fRVGHqftygKVreTH6p09Ch/oKfd46O1
zUp+GLhdn04Jk7tnl8Ez58cmSAo22/ms9c54lev1X/pthVypEQnIdWBUADt11v1L
OZapyiXAYzYUUqF7b739w3t0PWQ6E1mQqw6vC6eilOb0tZ3yjbctYAsU6KMXwRjN
6e6/ZQDYA/tj1mvloI7KphLJlN8x1bAVQ+YFhrKV5yuWTXPc5KhccYzWdvEqr1zG
ncCy7WMV5geUQ/c1v3R2Khyt4wwmNOABai2xc6FPMjwwYc2JXYXZQr3xq50c4N96
wncmQZS/j3kkQiuhkTgJgElIfZ3s8RQb1KjVaDURDDTDGbwVcoV+SWdS07FNcw3x
lteUiz6/GDHFqFelhdcwm+OouPesRjI0o+2mk3wjI3s8GGQnGRunKfEsoxSMl4aq
Vr+k45+PR0l+fovsmoqwxFKIFFoYpYBwjaaHW2TbhTiZ4Ai5tbIN3wsBjckrj8CJ
/wo0KhXnDEy2aVih3eH/y2drYQgJiccLNleK+mEUQuPief4UnDySyxVfaPV2hvef
DO7sCix3NN9MPStvgxemYjWanDId8cn+0U20skIU/Ke0K5rT0TkicEncPkd5Wmf9
VI3lV67dkGQbtiFCCBRINOy4VWaqh8I2BG8I+0w2RdAUBmCqwnYal9DvTxFklOnA
RdTwZvjvd870pp47v2FB8xKsC2IOPdHMcPR7Z8zoucxnz2/R7NxNzTEK7PiU8M8L
0vs0bRjvw29DAaDlacuJ+dgg7H69Otrjv1/wkbuMimTJep+/uQfCSMq+M6wJ94uA
YmCEV6A/8VhI4wH57kQf63as8LNRqZB1FdCJyoekPud5wn+acvLbjMRGyAChPfZT
Mz9jcbK5vCJCxdko0j1e0zGAb0xhy4cCNNsxvXO9yKQqdgF49bi4SZu8b84aK7lf
w9XMk9MeCyEKnRwqh1592GdAA7UDaqMXapVve9gsi/5yyMXIBcwJmK+yGptdip5e
xwDGW9xJ6IOxkuE6bPREFcXzW33H/T/k3MhHh1cwSZlUrMykVUfhVdj7ECRvEH26
ssnS7KzKJLrKrdCcuYxYwocZmTtRONBRzpxIoVf52CBVLwPd02tXB1P8dviVEKUE
SOBIYyp42rZf6OqewXmK8ZKFnOx1BRMHvBqygWuQoKviT0OKfY1cMX6fZzr4bGXE
CFSmK66cmDsSWa5kopEQNAzGz6v8Mt4fXh2fKLiU7XN3RteGHkuxF/Y5SDmMWqv1
vozqv6mIB5aSzDJHIIILJxO5tRiAjWoCzamlhKI51ErG1y2fJWT0qdnamHCe9G/I
bglog13bfXelNYFXj320xvjPqmegfqrnhNclvqCVx7DB2nZkQ1JO4rB4EkV4Qofp
oLx04W5vVwF+XSsw1Tj1d4IWH3G+JXQOHJh+tTLr5i6NRFv6CCtVnL5szbE2ZZss
GTIzokEYoy6PimaTlAn1SdENlbWF9a15BLhvF5lcV7Hoh7qHtutq/ZuMztnRmBa5
SYSNqELJZR5f9nM8WiC+sT1heaYtkWjlpWUgNzdFEGfJFW7DiY2lKSIwRqbJam/A
GQp/TXNGsFiLVAJm8gjT8Oc77dC/aV1KNNYDMpAwSwMza+m8S+JKJjt/XGZjR3Ij
94rt52SjBgwZH7hRBXBkeAHXQA1vak7m+WE7eAriEglvEIKc6IxcSp37qS0qC+12
lgCtafDpFGZ2yGUf/UPisnNqxkXvOm3ookbDqWDMVkVo7Mmlu1nxr1dXQ9vMG2yj
4jQuPUtmKnzxKwKpjjPwRm1Yye+OgwNkR+spx+Y2+Z/QHxfQ4IZMKbVebzrve37A
vrgtVo6SNAtqHBKfRNkblHJ/K0Y4kA1CPtaH+VSv/LnTBiLsb/tXY4TA+OLhb/hg
mBZ01AJTRS9h41YV9dlNo0yc7UrMVlceTtZhzWDWS3B5slGntS8MyBIM2ow9ffyw
ebMnCX5RvPEAh7rxpaqmdgSEBKQybbGPOebN9tFh5ZobN/auD3DbhIH2x4iUpppG
chC7F6KxYOkOJTVhEyoCaOlM88rQAc6oai95V13LFekZ4wT++VUqYhpBUYunySrb
jG9LI4XKXRoHLjW3vgkPSILk+4d5MuYK6A/prn43L9Y07orMF1UigAx5BsuYT/hb
Ghh36nYybNdQEk6x5mxTnAh+c4Dxwmj2AczE71ydGo8Qabk0QtcJgjBswvwN9oOJ
2V9ZZKhXmC7wzciPa8ex1P4EhXjO9+jcxftMAgyDQeRdiK0hiTmI2gRMx90E40cT
iuZh5O/IgirVf0bvJMyDtwDWEa4dJ8Vg5HjS1CaQyEeZneCoO91ZycBwIZiZ3ND0
nbel8GlsO+TV01hNWRQJ2Z85zY+RjZaiktHEv2V7l8ao/lAq7P6Zng+7qhcsENxz
LsYelVZ2TjCbeVS9FOm2CgOk+6PreGB4ZwlVPHi/ULaAtvDu470LIMQG/5I/EVox
Ricz2eXPTVQDLYy/bzx5cnwva7Ew9elX4muUEMpp8BawOePSX65o5lT0yWA42YVR
353LpJwYFEAUBnj2qAtzeK/A2hq4k+9uPQDiXkM4lHXDeJb3w22WbbSkrVWoJ7nC
zdd7KVrtouS9DtyeoheTtjN/UOcF1D5Cvvd/pliZAW0Avf/7JGiKT7aCn8FfCWGM
uXQ6+rHzH/GZfys2/NjWYjQ+zVU0kHFLtxfyv42QkE/YSE40r6HRPkY5B6sxzVJf
ekl0X93NHtffnBnutXBzAeYYsfBMvmuSYllatiy5NwEG0kCf8kV3i8C1FvRGX0dp
Fzk6fqr+WXsE69MZJQRC6OpYs/uvPPCne9gh4W+DArDcUPiJuE853CQgKV9TqZKP
9ivM5A9dySiqDg91orooFcExgXM61dMzzGaL4eTSwylCk4JCWvdhwu8lNGB4tP1H
u1FanPxaWh/HayFXnoiIrUo0l/8PNa+M1HDTCq/A1WvtExj5LRAtGHqC3rQmrHu2
P/NKL3A5fJSg1ZDMFuFu3JkVyIWYKsmm/eneifeUoZ6fS0bPVgJZk241HkBbXzOG
gxBVvReqZ0Eq8vs1wwsnSMQqUs7Lu3WM+Fa4IsevN7SFhvZEmA96tWbjp5l+Uuc/
sfT5MXE9ktZ6gxvVONOQRwdEk29PHztMg4/pStH/1MvDkIU0E8SM6IK3eRnoC246
HBNBDLon5i768tOGUsccgPGDtSRYkI3DyBMfj0m4aLrtES3rw68LNgzG/1IgqYS5
G+TrHjQAmLbCMR7lLfuosdx5Y4JucDaUCnq0YPgKJvkK+nQisbGBV7tHcxqSUAfn
4OOSC8EBEfoGhyqS/x5EURU+GNCbtQzjpLP8+p8eFfDeu4O575EEMS8RTohK4Yoz
wI7VxMa3X1/6LefuVguvvEejPAgRuK4GXkR9TePSQDgm5tjugcxFuDTbM9zYWueD
FtC+nAZq64TfgeSTW98g1qVlLTWppdgqxNeiSYVHjwrFNWWq1cU8Bhxn7fJDWRx7
e3/tAdiuPkzLPlmTjnUclNzQ32OGAQhAB+qNEgPVJM/hk3u847B4txQb0vQQTJdK
fyQljw3dKH1Y/nT733mw6dJkhx4rbU1qT40OfVKF2an4zVhO6QIbQJhdundje90V
JuYKVyF8vSGWGDh4DD+1VbfnYw9hrNB9XHainNEdKEvFQQcAWL9Oud8BElm84Br0
xARwcIwDrYNTVOCN+fM/TWGqXwO9pGa8blwqHFE8kdrpoiCwTO63Ar8jY7wBIKkm
Kh1OZ5GC1C3oBeAwDV87SjPJViNZxK0UInz29DNKNroMfafnL/aQYAp6jlCOLNoU
X0UsuJNBBG9PJmfymSVjWU6kKqmfidRtRWH22iERIRUR0jq/ausrFB9Bdk6iarsJ
znZX90oTChawzf4HwF9X7Vj/3gXnwO6tAE//SwfPSz48UMONkKOg4R+iNjqMJsIv
ZgWoUDdZB/iBev50Vt2KfKHZj72//4z9+WiMbrTcKgym2X6kJ0lkENJBBzqOX8m5
7J9AZEQ45PkNvwCGFnGsJ2qN6WtpXYoC6Y5RoEEKdlBAsyKO1tmlG29I9wH6F7lJ
UruzFQC3VYerE7JnZUDMHvgHHB3evbB5S4LcDOGBDrOdonxWmj7wIbYYptA6hJOx
jIU15IEYzxPawMS7qbbu5pHH/nt4z21E6mzSXL6nbS91CXuVJLUCF0CmUEDNbPIr
5wt2gfoeOgtEo5Kn+Bk6TpBm5334zJuVqkNCl5SeQz5BmKluonO3BY9/73QuH6Zp
Vr6PCamjVv8emf4V+9H87yYoPxFqNAnDGdcePqa+btgEKqMW9NSJGqINhC7BE2Hj
bdGyl1UmlQK74UN5+5OZGakjal88uBsBNiKYNt1fIQ8JD8d1x4fdvWuMSRrOEDwv
tWx/7lWmyaGEt8mwm70VX8sGpaNbJNquk0uj27nAFZGireXXn/oKmO/LTl4XZez5
YpOCN1S1Tk/YJpm5kOF9LrTQRpv5X8lLBOh5Yh0nA6wpyLQUALAW4fJLXMfmgvWk
3L1k42VMZaXFggctNRBd9Al4YuYzMrK9UcASxY6M7zVBSIlpGCTJlEY4/+a/p/ps
qOYtrY2jNcb1DSNHHnvgeKsoxJLTeP57eHRHeuzlrAeI0Gtv/+yFmt3DtTe4URhy
S7ZI9H9Xl33rWScjqYHUW14FVPMJfE+RgApjz8ppnmW1Eg0egXZEfIRtdRLSWB9G
Fq/EhxFACpyExeA7vrzbqfM+jyEmgBdePlczI+FaX+WZTgXijt1r5rEsDVoh82H/
Ps9lzW5NgmBo71HwACXwsu47XwhU2MOuBmsMp/q48SRDAQGdAbfCZbHBUUHAb6/f
L+DfKbJyzkBhUxiJnggPMNaLUuHxRzFq8LUv8RKGfPRIsbzZFj4CDSlOLYMtXwnY
IeUd97zwFzcQ9KNe6rwAgc10ER/nC9+7Q8giaBqxZ3x5cgSOUcadl6gcXJurccdn
wKbkCznO9xnZ87s0uy3bHYoUb43KfCDvZT9x/T5ExNrP1JtH8CrQo/vewMH//RhF
AMBF0NSMC4JCsTc1rEy7/Xwz+Bz2T0wiwlsfwW0/ygY9oU7/dqXLN28rhuhV+A66
dZxfJXwEWRMYY/pGnJeYZSBv4KGAszgKM4L+cYd/3t8EoM/boYx+thZEwiXGjo9r
6rkAar4lx1F8fv5awtfk2Da7bJtnuOdgisdK1c4bR1TVu83FWuq8dxxBzZpz0EZP
XC2PzOF2cB38C7iRHlw28bzbf+bMbYa6SUPYjTKnUUAs5GWC9EvI3OOHlwuuQRLz
tpVAU18RvXc53KUTelvmNcmX+G74h5YCty+bUT+xinCOuTY2TxPcOZr8Ohq72RDO
shBmwVxbE+863wKO/cYv6+iNEkw+9D9A9tDFntvy8ZVftyR4sg+p5L7z+rH2+jE6
hy6m5BIdOsNyTvTftaTfOzz61XddDPH2J6xwYT/1e4ChqLISXEeNkOnWF2fiDj6w
PPDQ9+eBEtECFX6e1iGFiKoyQZt9pr8kQZifzAIM1pwF+ommlQexQrtotJWEEknk
RSTZHC6dV3C2+10ous7r+jleK381kfl7ugwbJI7/+fZJW8kUg2IfElcJgoVqY4e8
WZkY8xXAJySo58UjVa1Hrk/E9KUjvz0QmVho58S8yhpX6DEdO/0InbCggrYYlT07
mVWuOPTiT0bKRwYE3nkyyl3tBqGpnPlGTjC4g8XoRw7V8VAyhznExWmUjycrV9+0
usjny9WcLMCIiYr2ewJP7xV9jBcvQJ6Oj/ry7afxefyUgaAToMoU1yFPAqvzdl/9
nvcxBRes6oqmqNN9dEM2k5Y/pEZKFx4muCiVsFVc40SzRvK4jibUbPy2srOa29d9
y8RvJXwZeejDcOU9MsLkrhGxnxN0dFV4D3IX1WRWbfZPlD+2m9JljxVm3z6A1w4y
rN6pSOpRSLTb/YtQXCxBUD3GVqY4fQEhPHFHYWjuORaNzDnRbrChgNAIlBzlkyOn
sL9fEUw4UxXbNJp3DQ8AlFlK9DLokXI2GgN0SDr9Ln6cpz6BvYZ+vANcorRzlE/h
ZX/jEe8KuHo35TMWXSFfxxC0izGBA0tUbtZDkYx04172uI4n1SCsg6wAdHLuyGIh
5vaIt9zvJhBRAHK/TYpUw9X3j4TUfA0EPoHKv0/c4zYCNJyWS3nO1k/kaq1+ED3S
F3lQkA+d8PSW+NuwOnuh7iQfV3xwGVuKZlCTa9Bwmct4m/nzfmwFcsg7hngJ7p3F
0m41k6CACtotgS+gToIVZRDqZ1Wrz1PgE1j9zxZQ+YH/CISSrisoWj/joFcSuVvb
XIA039ruGnljx113Xst3UX9WDsBh6nlpeuFERBN8haoUrBIl8NZEsskB3+SfgCy2
eO9I79HjTpvR37ojFyInvaJSPDmgWSkfVrhDwvIDL6MdYerJ4fJRW0b/qFcXBfY6
rxeWR+/6HjpYSoqU/4ZXIC5/44qdODhjFANT6936jxI/+QHTOCY+tL/x3YY3wmrD
KCc53yv+FhHq2TgXdUaWsxhT0dhLLeIKsW5lhoTuyC/u7JTuRMpIkoXV9AbuzxuV
lvsqn2NJullIeCoL5zvJQXx4Wc7sqhf8VglQjz3MKw5pSf+Nj/0QxO47ZMxOegJT
smnNGKWSXpDifiE+L+vWBpQG/+YX+tA1rMKwKgKu5QdOYCEpQBgDurW3smAHStje
9j88b5fvGsf7PUHQg9FZ86HazgKlVePclIHp8iD+XdJ+R6Mp/flY147O9qWGxIyo
eu+/oZ+MGicwNlfkhquGXE2YQGy2auAQL7zO146XxbZFC0UJtSg0hp8zyqa7O0tI
B99ubsr/sl/n50cAOLEPbjFHxa09KWQMfZxuzD4Bq7bMH0nG/CzCOM7zLb/K8vVW
f9PD9E6GIeygz09EniZrzDbXIWa31iZvPmFUnwXtp+NsXWyN1fgNhuFKQCc1JbmB
ZQW7TuM4E0lkSJ6NiNtWFrBQYROcQ72ENV+9MJDgkrdHZ42cXt2mEt/8Mn6cLUp7
hEQH0cqrSMt1wwYYHXZq6dZJYopgmJyy5rPqaGfUksP9Iah8NVsp2MZ5MfMLoTV9
l7A9osfGspn+CCZ+LW4KmSz+MM2XpC7cgg15Gfttpa65hGPx9KZRLlOzwqWNZoBK
6LtMxYBb2Vqb7pTA0qocdE8W5VC15o3dIYfWn0NaYxZuS65UwVrZUGJQEoKd5yez
nRcEcMod4AkF/KeIuehZxnXWYyCv1neURKiaJuxHpIMbBg3OmHkeE6BDwh0VzmiM
sJF0zL10VGKAARK8uthkqjgpI9LkEFlT4VWtat++KOFZzwvDudf7m9Fiaw5pufuM
5hycBcZM5PyzH/NPBtLqL4gNzt9n2NkL2JhL/NJEnhbVtmTrXbuT8aZNgYNUikLT
6j9izCj54+wrNsJ/X077N9ExFcA3PGa1gqp7YFWsQmKLpqDJ7GyTTWxG0dkdd4Ea
Ns+qTLeJzq3qddnpXdGWT3W6bKWNUAfsecEka6rIk7oCbH98Koz+Tf6h59uiDs0C
DyDyPQA3Xn4t54BCiP9ktbGrXnvNIWeyT2zYMAr8qt96GRRVbwLXazeo3VzdEJao
nSUaORdczS7UQ0RYknLJ3dye5iqGSN5uP6FtWkgDSamB3RrxgdD71EYmS640RjFp
NiZnDFf+ynJF2NKgmCyZHBqwlrLDRkf9Zyj/Ewe0D7X+KrYwc8bXzGBMnXJTMTNP
yrEjpvs7NaxhEgKc09DUqn3JGqd9gdhNCKDFHeXozgt38RLgN7qZWTfNtX0DwgzZ
gQdzzm2dw3wpXXgHN9db/XmZkC490JMukHZQ6fnRyjC4xlzCQiK28PSN/ixAq5fp
d3DMzRI/8L9AmY4ITtm9VW+PcqJ7ee6oOzg+pkl5cmr/lF2qtrYZ6k2WdgXXrMfy
sxavIAXRMoAMCEsZetPkBVa5xEeX53SqZrG1X57TgT5cQdMjqA1Ssx9OxYB8Fd/m
I4g6XiUV8cESN7hCTfFWCL9WQA3lLOK5DOUG7Am/aEKuas1CjoRwuCFncB67DQJZ
Q2fIF9m3HIXherOrAIVcSn2qNE5iACSJwq2RNS4XgGotQelVAO1KVMQXK6v/qQTI
YpRRlHuF2HwoIcMnLKvPT0ZndHrT12eWyJKYvEROipuXA+eYsJUufO4c5sDZkL+T
e/TpE55ZEgCqmxRc/96T9X4XQysIdCf5ySE41ltWp7fnqaWkej1F1CaoXwxIVGiw
n0lv4rd+PTkQ3D2rnJsiiEwE8ZR7jUDAtNVUf4Vh5PC8hfVqNpCzUZC5TH3piyXn
yiRFffTkE+87y4fAUqrsPGtWk6Jx26KWuW8hjSZ80xLiMYZTkaqduaCUc1NMqtu3
zEVqGJH7fu+niERD2vbL8JNpC8eSlM2FCzgMO08TFdaeZS4kaLA26uglunoDA+nI
VaZ6PxUkFOCgYjh/ZgzUmauHBpN9pvMtqFjttaKaYbc29ogu0ZPpDJ7zgdTDZEH6
kF6+LDmEfuvWNTxDdMKoi1YXY3cGeE5ZXdGFbTuEffytZ+pCU+dDqnEiJ2G5UdI+
9LlnyaAJr3b5o3KuxGkpDHWwmGU6mslOAora2ImwYGjs4oNrPxOQ06b2KIkZKyvW
ps2Q46zdSlFfqFoG4/E6Pwc51MpjcXzLJlXUkaoBzQiOvr3qZWVU9nm1DLQaG6Te
T9EYluyWFuGwJaI5ipW5gBkkzBFA1rXPnSes6fFM8F5zLdy1gndxNFpPnZf0hZyX
ORbISwPBfHz6fhN464VIGgPEMCi7fSHd4GPwKojfC2chtEATRHghqlpyWCBO4VTp
51v0bEo7w0qI7i1k+j2XCY6T8Gi9qHqmR6rerEj8xw4JIB6Mqb+pQUB35yRzRH23
TuYG56IzCbYVJ65JEifEEOzrI695RbcToKY4qyNcn+qdoyHJRCDQrsOPC18sSy1N
8jQPXBASbK18dZ7YyuJmOyeFraRyD8bXfzmHIUPcXH/2X6yvPMPP+XuxznHNsQbA
fJxp9vn0G+vb0fokOAjwalZh0lldI9UjmyNhakWvReZLWb7ltsSw0tcMfzFBan6b
eJu8Ogakdqy1e6aAODwHAbmDiNbHazDuT2X84EiQBiVpJXeTLdWUqEvoOqqSuaj1
rvqerS4Ff1t00nhCrab18Kzuq+Y70PdNNyKkUiOA3lPFJQA/axdBFwyGyzsW6yne
5uXZTSXQCpLhTTaENbSswanVs+LHMbcTdieSVyVskljYM9ShIgaTEfJDia4wq/4x
ukEUVeYY+gYQVKi626Umo79JaxOL5USQ/+FXGSBof105XLV3/PQXyIUzHs6qRvJ6
jmXAdyJxWo4GnU490ppn/YplNXdT48PjOMzp3HTOmty9EWtBf2JFOzh9552igr4P
UiKCxIrbi+Pd6ybsvXjwyIFIf61CiWYB8dVn4BOIl+whaHTMQJY0Zl5pKzwQXiR9
/CuKh376T2p9Uv8z8vubbM4lcWkCFYi9JQIoeCS3kqhP31ZAmekS7Xk7hBW20v+C
vRglt8l15qM+jzNVEvVX1NBVHpUiM4gtb6uvJWVMWLXEPaIb2489Pr0BzEZxBrVt
ufMlN3uE6SUytPAvr2P4n3vConMYdlF7B0FixMerABi35WRz/7sCMzXWtQwbvvzd
eofb1vBPA7xlT18tQV4WTrk2MyWXn/+HLz4sacY8zgV2H5J2xsEuaqkjRZL17vXO
oRIdNZjp1VupRPcPrcYqHBH4qPKe/jZq97kwv7AFEhsHGxKRC2E6sKIraqxmTd1s
HYyMS6A6fwCVro8IHgm5snRojLDjSpawqKb02AYCV6Xy9sKgmAs/tNL9eqb0JL72
BN12fnuE/+tmY3+cizGK6GMBSfu2s1AbbGubjytzcmdodjQc5d6Zcfqd2CAykMbn
mjbLWvZKA40h3CSHren5ZiOim9nfOFGX1Yek+7DMCAoKa2YRrLwjZeolibXsM6su
uiJ5faWrIe2DfVKrIcxZbasxtrObiIrCwtBCnshY7u4KR45CNtqLBgcsBhNXqNeU
bT6orY/3lzyeTpOjexqeDFQ4zDXhmfnMI5tj5wkMoES0g2knPEbUAgpIZxS1XRhN
pdka5li655s7l9X/uDC8wP4SKVZjATLFmUG2n/VRskGfMGoI4Srjp3YmfBqr7t8w
/o2gWP3AeyZmV6OvqxfioI74lbFPoTabY66ClpAMT1tpJ48IeTIb2Pqb22AEtsYr
6R4T4btERxr3BSDuTznBZsb1bc2FYhS+xaXEYOao56IMm8phKTCbomsC9AVh5pfD
+YB0N7Gs5MGoUKrNLAeyPlJ6jn0WsNs3VM/0NN/z59yLhSSSv1tWBd7MUUXM5F9P
FxL8wYEEl1rAkPtPfqSgIbobDtt87S+9qTZcFFnIiSXIf2Vq/vl5Ps6RKJK3zMbq
Wv3mPYTZFh9bqcCv6ICWrcpM9jYPhiP8hiuACupVD69K2F5pdXxg3VvFo9gsv2Yt
dUJ69AmAv7k2EBJQu9sGKvC8Kts5sdgKfcrX4XFz6jOy8jHUVuVe5qF6wOyU76oh
Bx0nOHyb6RtKPpKHzU3H9dlQbIzNTkplgn2fKu92vuorOIROsBa6On3iY059bcok
rX4C3K/okx2RoJrgnmtfmMzZ3Mzsulmpu2VmslojyMzz/3nlxnCbhjrNQarLvg4t
8s4Wj+Y5DHDqT6V0D5bWKjrtfuVt1wFM/sHYo1+F8hQBjZyb18fZs2aszcoz41wl
nVhQoUz+aP5kDLrnCeMvW/iITmPBxf+V/l/VEVmm1yojDWX37vvZ+3Y8sxaaT1S+
lP5k9gk4qiTYSr7utXD0T7vYB+dbCUyP2d1aVVSeNfxVptZTFIrDwoVlzzj2frer
/0CZdUc3+YcJ/uAq0H+iALErTBmM493yf1R6KnNEiC5SP+MwdPcMEGzFqyPR7vsp
q9+31sRNj1ZAZ7afR/Bbc/++1NiupJdmKCHdwPv0xEQvI19W0TScwivyd9IybMtL
mwewkFnup3C7kqR3obVdMkWEiMwzz0Sugf4hzYpeTMRtWSgLZrrFfesMPdn4Wwt2
Vu0W8aa84796lvdtRE/bkTxZ/dj8CaNeJ5/rLn6cevfyX5JYttWIEaNd0iM9WOOc
VqpmTLalvhVnlfMNGuWOcgYO0Q0/NX8evDXUGKFl7k66+z9Y8RrmYc0XSxGncHUv
biMJNnQStWYUPeNcDGte7XuciFLJO3mMrqRs6E+w+KdX7TtxeAyv8wMssvDyQU0h
W+gwVOVDEh3422FKzzmCFAduMElcUvaphZ+6uSvlFbx6EH31+J4M9vOQkEVT9VcF
AGBrH+dKMm1+fUs+qDLDb8ipQQU6o6QTJBn5mYAb7nTuq3wYB+6TpKHLUkc1AvXY
V9znmgY2mAHLzOSGsTgt4yLq8UqjKZIXEfTDz2pL/tpDelzPPzmFVH4QtnMvN3xZ
xvnBG51NQIIXKJ1HNv04C820swY+dj3HOBUBIQH57zvZ0H02oNuC+Z/Bi8E6PaPR
2w9/3/9Uxok9oSsIS1dSo0aHiUnqFogN6SfqGGyFi0T8ujNJF/j3J1UMJh0HgM/8
XaacXH55QLErygv/txBkKXdhxxAd9QZa6PBOy6xBg5AAkqI1CI2A9ozikGc7XSUQ
2yrDM/04uPIHOV095NpQc03ZBVyHNxvDHBapLXKDsdV0kpgx5DS3+NzlqpJmu+ul
vUvJyEWOV3rzNVMKQf7iVAMEOKLs+L4RMhHI4zakLaiHyseKD0pTc+WfWHPfaZUX
ANOTX+vzk44JFxggy8hgRvEKbOmdTrQ+d7sIG0inbBq867fVFznfLcY8eYaBLgMS
Ssh1jpAdNz/5W6z1MGDVYgWg9+ZDGTeIuc9/S7Mutp0RCEIIFHsJGqP1QHqOCZmy
sVyzelBqdBEwi3Ac3P4D1I0wTd92mjxJovcCd/fJiGn1UnyCItL7XsUZ61tgJ6j4
hef5jJEfFQWG+minjeBL6oNVOrhLPAwKef25i8TzQsDErZsGoCwcK0PKCP5ZQgBO
mxMV2dnFm3l9gtykUN1CQGgDxiq/Q+4j3WbsFrkKUamIhu55saS2xxf2EAtQ4o3R
KOKtXuqy4ueS5pVj+TY0Qxub4/VnL7TdZUy1jf3hQ9lTaB/BanLvcZ29sAx7elkh
9pvIcES94oXzEopUpzdp1py6Emz0Ilflomm5Mqla0Ona84mS/NZdKttvnhXGB0LW
GIh5zkkmbq011jKvSFXms1ybEX7VAB/arMootyxhduAqjXKDNCx7RjxCgbslQ1zd
0wqt6kB8j62Ay3JG9OeMiOSTN3rs4hx1dvT3rqf3vVkAK8OVixfmS1NORHN0azgG
jtV/igG90lEwxn4e0nSYDRsGc7G5JjjnccMHTzuEG/wjt0MMREufPSrf4hEXn0Bi
fPi9m/sQCrllQVtHgQhLrCIezh5Ldw08Vnvay5pCJWq5CmhhUnXvg7sQTKsxFlI6
HYy/g0HnhNx5bRruWb0biR6pxWg858J2voxlv/sazuqVcmphbC3T+mP4InYu4/Xv
WybIJS0UWGcAPixrJfWoezZFei9oaB6LpxQZJrsZt8PLe20YqvnC511WCn7hlUOX
SjPw3E1WpwFCVB5YUk8zCeX+lWssAE2OQ1AoNMNl3CERq/arWrCilu6kJ61HCAQH
vs0rV9q9Ey8AEOy/XZ7vvfmn07nnFHA0OsbxtG7TJl6y73dxVB1ysyuwgNikRw5H
fg7XXCyzPD/gjjpOv68osvMZgo+6UUuT4iHjvUL5Tp1e6fSFsXyrSwFJ1p5stCMd
ViF+PrB/ryHIorougklcMOQigd8hxEisuUgGgo/nr/A3Cmw8oDDlEbBRSqrDsobR
v9mKw1l0pB5V3td/gc0eLvhkd0C8RLNd91o/qq753NbMJN8bxTr4edsqc95DO/rh
eFpvgmRA734CRrX+Q32FCavMYihmHp+2fFAS1E0hEyWMHicJbWb8WrRfgjMxwrh1
MJGz1dJzXT0k+3DdtC+CbvQV/hA+AclBb+4PvEss9WSwoTLXJq7R3nqN6D59rnls
I+bps4ML0923eTR/miUREifIR5IMQwSEybxcx5fny9sNbGHXwHbE1m8Zf8Fuh41S
5A7QyLEzqSb1AJl4ZFxCAvQRgWvEZFNmJVhRHTNHzaRGgKO80je1O63/z5R8/Sfh
DVW1d0JQNGMk6xXcbtsPK50e9N7Q+IfePdaLlPzKbvfoCAONhoGMJXDeZxao3pQk
7JglapoIeZjUGEL+mO5B5v/hhgwmJfBEJRtXoTv+qOWfIUDYnMeszJk1S9bBYYne
Z6wlaYKu08tFEINX5WbXhYXpcG6wOLaEd0dy73/Z6GI/eKtL5aIVqcB7sYnrU1CZ
ivxqxRKNZl/fk+WTqSxmzA9CbxfhGaJeOlus/LiV2nRB186nY/vTbQcnZu74rArs
OMA0YAVEBm2NUynZp378wfJvq4vMwKw0rn5MdL55K/YfQDkGcjqrpftAiXNfizK2
34PM8wb/b9Bgp0fGPL0W2bbU9tQu34DgMNMJ6IwupN1fATzNKfQYvS9tleLKIb8i
20fjnXN3DdGbY+HJ6SMkQtBFN7QsUTHbgbHDp11jZYtLEeGfvN4ib6aotTF3bkRN
p5HySaZP6Stxwa8+2qmFNlMGiHUAY68gu1mEkQA/DW9dTN/USyypdzRv9Kx0RPOb
GstWFzzNjmeyKrmC6f9k+RBSC7pPh8ea4fqojgo4Le9meSWcZZuHUDY3Vgy9nSNF
sSCIPYVQAx1dwDTov9qOtgQayR/bIl2kqgZU/V4GsEYMFlxqTMSr+1sYHQpOE4Jk
0bM/YZLKbCQc26V8PwaPRDvVJL+BUf2MzMXo8NPXU6bJ/ZVouk4O7F+vV+2mpV8z
FJwJlxmiTn30COUQW7z6jL/d913/L16KTA4GZeCRyTfXa1/fyfVPXskgMaeM5trH
94BAFwd5MI6B6UO7NMQH9kMzVr+c3GXygE0YVO+oj1tHivceVp5x9BGeKhIdCp/R
vdCSJ6XCYlpgfdTn3HR7skoDdaOz2Lq0vtZXolEQbdM/fv1ChhS4/ESBM0GCrEKo
NPOtUKZUdg8iq9qJBf5Md3jFogzqqne7EQ6y3OsC6gJPheP0w8UDaDAKZyirAqAX
hbObtrKgllxtcebhlGhahAxIB17r/ocTWyKx+uHZwp3Iy/X40JRAs3S1piBlp0rP
0ngryYZiBG1AxVlksUq2R5ge6nNV7YFKCSdsgnEj+bD1aIw8CcEucTde0OiD3Og5
X/BbkjICHjL84JIOaDqRKGOYJElbU1GIELaVwR+TpzCLNq/KyKzw25GQ40JDtK9j
fCLsub0PNvw3vPTGF/BwkUMgghR9CX7SFFv45HBezhvKBnTb5Df/jyEJNP1reElw
Sh9KjwGgRpFyEpdp79D4yu6Ipl4ALlO71Fzk8aza6G+tp9c2vg2SAqI3wrag+TmC
/Ka9JeEvq4s/TsEMjCr4By5FaFUsVZbOSlsLwpdWHHDLj6jiKSJUyth1I3TSx4Rs
vC7zR0NEuQu7JJ4Q+SKdu0rAXWJ42WKHlrQ56xlU1Fuc0tCXEQYul2M3WVx7K4iA
Vc0RleQBPQVr+LxGEapxVxsB3P+qZPN/ZiYvLUd+0KBi63aR1Z+l15HjIIVRBi+m
zojP2TnKDuzad4deLE8JgZAxtWJMayLwVyA1F00M/diCPj8ZgVI7hACUGdxKsSGs
znsznt1tLnq1cjg1VIeNw8zr9v68qck7B0q1en+1oR8HD0pmezdiykSfo7NuiTZQ
Ej61ExHO7vbwJRi7xo9XIgD4hs8PQnp9o0MC007ABQd37pTfzRRfzKXFYDPpALaB
HbGHSvo14mLDsHEh9Xl+aTWH3boQx89FNSTlFutqeUBFKo3fGuuOjufDIp3On8Fc
MawEu6KajGGYCeLtWKNGTiCj2Ift4/nm+9xPSUgd0FfEQIDsonaedn3ky67MeZk9
aR1Kii0us/ZLdDsVWS3f1PYu/F1a/mDXTSagSSsS+lxx8y/LKK243hJCQjdauU9R
+qJCIT4Ila1VgD6EmWbeGnMkN6bI2V2X7VjrrLrFcQ/e7h1V/COPEDb9k+TlBSkt
K/ENffhXo341g1R0H58bZEQ+JXkb8u1kuSY5gqfk0VT+QsgkHVwzz5A1OIJnMtQd
GoHTyggQSWT3Hn+oiXpBP1V5pettlBAMgFsTZ18eqMrdV0UdMuriPvK0zrkq62k3
RnCFQoZbbA4rJMj4DHKuVP4r57HrR8SRE1HkZ/Gzgh/cie33M8K1VFM41gPrYcy0
sptaPZxViNq95RIMTPjBVd5bGtU4HCz2dR4P7EYcowse5hsg+CQaSy9KiJVk5MQj
XRDswkIKxO57rdM7QbqjQINivlTklVutn/VERdi9Ao7wUSgyH2adiqUHs2fXWA4J
JS7fmGKIwztJkhV1tob/5ruxVIk3ClXB5F0cgsOV5O7hQ/S/5doTgqba5UlEIz+a
7vhpmYDTbZZXjUp/B7akYGc2volMkw3CI0IuH4lUqQe2PSmxdP99dKoYvnYINuz6
VkpZUrXxGFfvYVGSDgT0hYcAMoSTtUg+Xekr5zU24F+uZM01uufoY6QUaMf24Sg6
Io7Yx1vZfXqApRhwOiPfoV3f2qJHmV1hYwYQIFpKZE3GbqU485bCIwostmBgHz7o
vnGzm/GLhW6BphvAj0qKcuQtqaV67jmvX76+uLm9GvxjunBjbhG+KvBd1CtpurM+
7zDtByPKEF9DHf/EX/nD2sghFWRiMTs6Q0MBCUztAtY+PkLiA8I5rUrncNafnkp9
i3cTHr53Tj5iBq3dxtjzqhwHebb2q9GkjpXo1aG2wNDVUIkxypyOValVb5y/ZCYW
kJkw55NZxv63iMGq26RLvS1DXNM/7AD6ie119emyzj7qLWi6WZwjQBsu3VqXb/ou
fjFTptZRaZiOmLm7qM9AGSD9pPM9X6OunvMVdei4p1W0pAYbY6ixm3j+W6T22BnM
x9QO9M1rxOqMWB1+0R1IMDHml9h/aa+liDmvH0X8B/TOLcy6HtYBVmb6YWiNERUF
FGzYkycpJZDglGlCSpuSyFiYfkuEgx9soNDZ7w46cfSQQtGOMe5th6ldP8jYaxQm
PZ+O+I2wk45ivnUQwF5JMFfNxDPdn6SoAWu6F4LdiQyO0SnLnpzFElzvaFUYJPvA
2Cl89aeZMGFPba1ucgxL0SRnwMDMWFiXmIHiqHQ0e7HsSIa4aJYwf44Za//XdQhx
hykRUyv+aDvwl/Yoz4qq8kN5QLrGdN1/RHRzAfrpOpnbKwUJdy33T2NxJigJNyEw
TumlmuyYAAwQOvPk8xCxo3iZkhaKCdK5yTshamlyO604DJXC80HrwsMTi9CZMkkH
qccL84sHGtLvfG5xLWyTlAAORAWyHA3amLr70Fv3Crjg917mcKcuWzccN1E4fF27
AZ8H3hZqQN/AGypJwrzM9iOmlU2jE58gi48t8B8MO0uAXQU3pXwEh/tj/ylsCP0B
PNoYM7THrdYOh8EivX/Utfql7fDy3jB8uy+LXaUsc47uPuKwHyB3OdBdSsBi8mUh
y3Jo7oCKSGpd1gPJ1t0YX1CLRwUizcxrBs+3Aq8PvZVCZiG4HsabweH1+Bw7nYhl
6Nvrwnk2fYdZuWsmd3ngI8SbbdY/1T5LkFsIt+4pusxFkCYknCy9JHxiQvPXgFvJ
0OgZEfxu0PT8mv43qUEhOwLbN9HK8XBUzMc0I6EkyoXBkGGtacoWcRmrSBzK8KWW
cmr+a3XtkQ69nCorGiNUAVy4I1MhqXHiwaud7Q3rIOV2EwRUMj9Bzv8B0RkvCYMK
uMgqF1rw7eP3iX8JCPnWmBYj8IhCsYMua7ZnnPel0vnb/p+TyP3GkeUXnv/9ziz1
sRyfepGbaMwQ2/Ky5iyt2Uo616SrkvL6DCDKPbXE/2ByFszlDkKVjv8ChsKFg3pa
RzbM3IPdkR5eOoohRF0YAHjq4y2Wiq+s8NVtWeEbZCe67u+8fwVaEPutueEuNgB/
kAisc/LrbxU4Ul2e4AMZjLX/ebP6NITLjQcF335m3PopcdxGCPfc972tvlC4jd3R
kt5oWh0v1WBs32BaCsy516rlYSzfxYdgmqpxt0WwQDUwk5sAv9b7PpaYFH+dgy3Y
lRkYtG+P95WO1Jfzmrdt/5g/HSL9FwpAz/U8IATCfzSLJ9q6ShxS5ToRUiT9f7fa
X5VhvcynTvg1OYcguTvE98OrvShJa0nCE+XHwtRZd1vKozewd2NEi2m3Tc2tn21S
pmeSzdzNptiWAhfus0ljV7lDtNyKU0RJ+Q5t8uieXuTA2ZKp7pbNllFwuketyjiC
uJrWMEn8ZYruOR5hYMymSuEOERC0JD9Uck7dfINT7uEIrhNCX9LYZjqY267a0Yjy
qLEGEwUXMoqcbAyR9pc/YsmIyJKl0fnPcURYHYuPwbneGArZjabencti37rvH7Kp
HabyP3AyL7w47YMv4wXNLQNswicvPo+YfzonkIFYCrOhw+ReilPtP4BCnHlfU0is
/Qv1CkQ9YtO59rvRZYxIBrldag0Cyojty9N5n6k7ik5kY6KLd7n9/HkTXJmh1INL
ytxh7UIfoTJfoKEgYqk0jpoAqT+9mreEwqm2ES+J3VxYQC7Rxz/8FuxZo0g3eKo+
q6fgMOaa2ar/AhRS/8eK0d6UYX+uNvALZ1CzrBhxDNH19pLoRG4rOG0qqHqe0n+3
1NqKhWjaTE+H6amaI5j5gbEEgGp8dcZd/fqQwWfqJIhy2G3MZJQwGTko0TJfWc1O
XlAHx0AVz7ePjy21ngYYv54ln6DBFCX4sNK39EL79yqmbOV858neJZTLX4rGgf59
AMdNswEwDWYmpfHfJwfi9WncuCT8RxhtlNpOW2RsSSEUJXrpM/pquOqlquttKzAz
B41aXbXP6+vQJ2DqYLAMr8bqTnpCeQRzGYQyoBf88bU54+hvMZgxUQ3PyZoWc0EK
BDmsCDdELtyCDDXp1mJZEhnQS9PVQZxmIdu+iYrNkid3yBQWaU+CH6Kw2kA9Z7HW
VdlvCJnRWTkZ5sOXUWL3PHqUPLSXVhwIyfvTqU/5FmElpGN8nWwZITEol23bDl3v
oDykSoIdvCWulgXX8EXc8k4ExeEmUK/WW066RiAxPkK6qrO68hH9hdWSkxijniR1
PdgFC6ijXz1M5EGbyN6dxWm4XtHFSIwHXtXttwt11R734TkCw34+JFzi/k95ZywO
T7R5raBa6WPUknczgDXTJIDGBbJrh7+U+Z+RVRnyudZWmnMWLyz9SFj8+c7Q7Oj4
6kmQT1Y/H4RFL1OttREnkBLKrlaKz2OfxjJ6PfWi390/1gTBZcG/gUVBkTl67oLo
Y4iUZG4ebhBfmnA0FufY7QXXQKPWs0RhazdWaowqhtQOxFZqpZ2C5DrC1PrqJTx7
GNutb39V/VPxr94IvUeGgHkBrMDds6ssCJUA49Ow/my7cjJNvJNAZD49q1iky/VE
aQsOBLOfyvSOLSKSAlX+p6VcU/QSmTrJyBUZ3D7QUESP1LvNsG+Kb8MJ2LjhzxbE
XAbTjsmteXwjiu2tWQ/pts6nK0Ir7jvD+bDQQhONMNUHHgbUWG0gF1POt8e3va1C
qPN9qEg6DXMBKf+oQja3Z45gaoysu4SPWlvf4JyGBv0Qrip0IbeN8gVsw+pbFJA+
nafacvcrzWp/oNAUntPzIXW2Ui/IAuZyQtPx+aThX2uXL9FFqXR8r241kwedH8NK
UHq+PrCrAcv9kylhpjo7fAmgv96wJcmTk/ZvLQiGScb2Gd5dkU6Hbd4TmaxqKlmn
S/4y+ZM3IIotEhCRQJfu8J9R1GVbSTPXEq8rUwjCPrDGqM1H+FMOvcb08wrv4jzV
RhYDpIvD1SFCl6D2ZPRH5qUlbgfZPXjpXD/BUxzR6kp9nZyV3o57VcQWKVLRI3GD
CFqCT9CnrVhOXyTM+uTkeRG2V1NDf5OiSmSHdLT/omwUriA/XjTS4iNCsPbA6FDE
6DVFOSagb+uK01ZehAuxwAVWtiasfE9ThvVWiGHNDrZBULtPjuaGfsf7TOzai31U
xRZzNHtobEAqrg1RrEVYJlJE4S5vX/X6/ifMoitntg0ayWNEDaeA3Rnk8qc8uZ4q
Jt7TZkNIa6lUyKcfBeYz9RZW9B7n+8SuswHvSopoaQZr3hTCwgObL4M42o+7zzC+
xb3PXiXTD+QOODLs+Lp5RzS93ZyNCRiufkULp0j73gu2cvEOLfCFKQFz3aExhBxr
KCiV2/7lLbkcpHyIprytmQEHK+BcgAGrbdOTBjJDZB2ZyPCrghX4UCVqc6l6izg9
xdQTA+LozqJyU9tyNMpmq4YWYr8tYLT9z2WhkV4/vmiPRG291Yr2nKY8S9VmUKw4
yftjdn0Mqg2F18nfG4cBbPlvDyMzBBja6JgwpfkehJYtO+1rsBgafAFFE0dGfMqj
Iyrxol5Nmlc6ds0e2GPv3picV2vi2Nrtjg0LIrjzC0iiuPCHFdPhxJqwqWg3AZFp
7FP07mfLriLoQFWKuVotXxKdaLHCealBgj4F4lZmZxW3G0XlFqf6kMyDHJZy5Uol
UulkzmnKKgpEiemcTlWVpNgfvq5favgU+JNOjE2vmVBA5lORLmfbgPbr7OhZhXci
gJpqjNKAat7LLKh7iHH+Jgq0GSuQpKJOu4Y7f8a4k8Lff1oXn8iBKm6K7o9mwgyj
fO3YO00swDNlYQpLs0rHG0pT3SsUjbIptkPhGJ9V/rj38Sw9uSwzkwt0Q+k+2RfR
BIARhEGiwYWjGrhm+QHGLmmuPvtvWnyHTI9LAqBu+y8Sg1KlLYKg7MMjRbH3fR9Z
QSwzQXxxPKzFJf3megA2IpoUiCnB0nrw57gH65q1xtvEDnLK8hGKZ2QxysP1c1N1
NpqPJc1HIMeSrQJ05pWNaXJ1P1Z5pQxvPbxRDhptYaUtBsjkACmPRg3279kdFCU/
CHA7szRQ5+V95tX0DELNGX7LBxHm9kS/d+YNBWhWJyaB/kCP7zsS+U/SACGLhLVt
bpk0F0yhw46N5SWd6klomaOvfXldykLWJd0dLT+c3JJjinPdJcqCmbj2jKHLLkw4
R0GLY5fRRfc2ADiyxdb5v1u6SYS4isp/gpev9Z6QD3jiEx3hL+4+nzZ1P4OTmLu8
wxvRVqb7qnk+GYz2RGn5kzfdGNFQtgXaA5shIOSLRYyAWOGclJryCKDOz08SPmQw
L4kN1Uuk5V6d+MT5lHi54TjfAIqnMT9g2p3aGpKcyu3omRLb+18vhb10Xu/y6RIY
W9cmZAc89G8etPtWz29AJRvGOR0/045RVs2MvaC/tEVnYGV2h9YmFfDCHUIstuO9
p8MMeiOoYX6xZM/edX8dwphBGTkliz9TzaBDmhASwn1JKv/Sy3XoWHduS66mkWNL
xvmJEVZ7YBa8n3WZ5kmtMrxAA05VJiuOTEDG6SJrAyEtOrXwldswZGaDDIv0EoJ4
QHF45Fn4q2INWYd3OhEfmLuGliRFc911sMOa+o9E4ZB+LRB/O1ltWxY2J0nDfpqC
1XxadU6+tKTSp0ZMW6pbCxyGFsH9odzAaO29jruLgyToDq0Did2wufFRNjHUDZMc
B04iDt41krcICBUu77ZvHc5LxQjIcetmeQyJdfWpuVodCxk67XVxBli1iwvVCHDl
n0FfrCana6pyt2VEp3M2B0DEsF73tbJMRXO71uJYxJDzdYFTshJcMF9OAAdBRI8I
iEC3b8+y/UAg/8Of0bNJYTkb4KHdsD0OECm0QcCS1slCEzlUumukmXNCMb6DPFi+
zrXG7JlvCTmkU42IC1O/W3ElPVDy0LuODcnHhQs72NZSeDHxbhgpcfuADHkxJmq/
7qTGLCAi1Kav+G7ZgyBj3hb3o6MINO4mvZqhIMbsQixrC24t83gdGSQyLlOlmuKL
icwauuOvUh0pBR94rkkCygi7PWabQAb+//Co7HAyDoaxEjwRqe/Qoc/1S3+lq/0I
yr0WEcNPxGbYYt1Nmgq7iVlsuDyjlr4obCCfXQ7lMTkgf2ld9GRvW1l1HiWeYvGS
uodYqtAN8xKdEElReNM9PZ2HSxA9NbTf1Sh4coOaR3fcaR//BVlK4xMPvE0axulo
BfGeQJdejAzJphmUDS9fejOlMAhSYHCqs7h/X8Pi5dOF8cAn78YjlimzHgwqLmK4
hY3tMNbyciz5V8ch+oNyU7cTjYHAXGcL+G1Ym7DNB2GvCAKglMw/AmHgAHlJ0MIk
OeW9PKv7yhqPbdFQRWohTeewM4OA0iuhBri330ViFyDnjSidlkHvdthu/5NwfqYF
V8vN7oYRqntOxX6pQ+2DM+LKLd/2XhDu/KUPTjK0bKPYzJ7+5MQHlz4FhJBcD599
dfgdYJSwQKdjE2zCdBCSxrohk0NvQkHxJf83vDjIGk22sSBiA+TBQbpSvcjCIK4p
lDA4/GEAOO966lxGuJFgw/NG65ow4XaFyfgIm6RzJE5uu7V9g8LE5CCZyz2dIr98
/U+oE2pOBqE7jV7ls1rZLk15MCPccovBnZozTSsqcV52i3QODFCStDgvnODmIcbf
98syCqmspxvz2lwR0rvwhzBf/w9ZK0ujnpkD+5Y+h0vBHU8hrcE5NHNDIPg7dJsA
y1B1ptax1xX5QnwMY1bFS3hVMYJuckHnzxcAn/gHFHkwHOxupGfIXCN3POjL9Odb
bNiyYzlEgkQmtMYbklMx8+qHWhThFAEuvWyWUaIhKevpGY7paFSepQvG3kiBYRjo
3kfWPv7SDqV1YJLjE86Z7T0AGQuEk3JmTvt1KR8YIM61EPZc8rQbMzawB647otoo
ghs/rO/1Ne/Tsp8BXWWk00B8CFzXp86wbyIr3qP2q7cd5QgDM34yD0+kZJRkYRSo
lWziIByN8Nq8w0bKcK3KxkjMPueVVuVljpZ46kNtmQW39ZvyR55SvSsHm7vBYLPu
DfRXPU/P2IHrnixNl+GPrt/p3rsw7cX+xBPN3LBTo5u8stQG/xyAI47sjmVqBnBX
083XvESuJ3qYT7ru9lidjKQZ+dtsvXUUryXUBah7XIGwVrXe6ZT9oGi+Y9vKa82M
vKyYCQKWTQ7X8UOQYFFCgF0eCsGmaSSucCEmwxxCmx5QRFGD1CSWTKTLN5s6gRsB
LmpiCGt0ZKLSXznSXmeOBm4YX52uZ0TAXY3VSeoNdkJ7bT+Bk6qFdbbHSqg4Gwj4
bLthLVu9VrFAR2cs1thL15khzRbJUrl+5QyCM50SBgCH7HcEyfK3AUr8jKBo8SSL
SkD0m/pc5WSBZLKiUerRuxybiUOo9hH5MiDjy+dAPDQqTM5Yv17bJv+MXwCRFX8G
02PcbXMHww2uXaWMTRe3KEFAXd/s9DO2V4JMIiU5fiZQCWUT5yvQW6/Eys7SmsH8
0lmYr7uwsrQFo3XTUvfhXLt9x99q4YyBYFRCX8/s2w4lGp3RvLBhwskFNGA0MDVD
ET5Rx3njRLq796X6aDlKVZ+9FtF8bhjiMiwkMjkbBE6O17K2YLXKF0nbOh2Fe7iu
hlKGJcFNPLHyTeudC/W/m4byCBUf9MnS0WL7Y4j/7bJZogalaYsMbjJ3I8TNgukk
h+PdGpfVZjyMb7CCDzjTRIA38ELe8BspLBYzggKGMsDWn9AQ1ddqRCNR5bV0Xr2u
mhUatq7AJmDoVmJNDE26JW69S/3AzAZggzQFdfn+J0gdpEdAxlnMcOLl2gg9F2Qn
JUwUmtR8VTNWx3F9ouIl6NmD560vN5sEZ/J37kZt4ulhL/3Cn90lIUeXgJd3nhrs
0x0tYHVlyTgkdoAjwV27Tn3y8J3pyvJzt36on99d9BT1dXdpfVcZ3ztXFkO0A8r8
f8l7FWJl8OHf/6D8As/l4vsv9bDpPAnKwuMj4Tggko277Ni3WT9uD427K6cCpd3r
bZJEXaEOOqI9yfSlXotsTjHLAVNfWfn/mBmVhWPQeRwh8AnrztHEjn+S9UYFqzHd
hz5WSKyQ6rJXRZp2kk1rEEDKSHQHJOYrpCM0fqnAq3AikQpXuFpW0QNIufdtRlS5
r8esQ+favrDapFhEvtr08fhbjvGQq9bt0l7qhro0L/X52ZVpgqNvLp0DU9g9+Zco
25cPmoC/wXuYKCb15cY5l28UKs8ueDWxywTxEtno5MaXbBLbt5c6e2hOS3KYZrqZ
jiZ7kwNs1GNoe6oCwBKcmGbwaqp8EKfJZDl+v6YF7LrAsgNdNEkdG8Kor8BARXa7
OfomBZnft9XxbdRPBzjWj7eHwwRNHuZuKTq+T4uUKEq4tbwf3khrkchScdBf9hqN
+5E73+l4VCs6lYyOpuVs9z0K4i6p2pDeX7TP2GhKmiTKZwaqgrvZK4xCiAJPVgnw
nGHBbgyVEXdUbXVGSjUOQycabOvpICHzT9TSyW9cKhXzXrn5mhwqsFMxDmLgom42
WJR5YraTZbFq+V5dy5LAY2dN+Nk413pNjNPKDuxG2t8FDAnUK8CuUV3Xha1qCar5
DogOVm8ZaFjDGU3B6JSUc568dyXU9NCvrYZPgGS7c9Y00OV3oEvofOsFkF+V2z/X
xVllteRsEPYjqFhcud48JQCBVHS6r7B6EJriEMrQf2L6bOFl1vGU7XameBDxSgle
4vOkTmChZ6Ra6yHiT4AsTAOz62w2Kvqu9RekfATAcismT9Lbq4iva5qotjXP0MED
biFgYpm5YPqOtTBv9hpb3fRS4/smZrJLfZAM6L1NUc+D1Zhl9Cuk7pSHwiU9QP6f
xyBa+keE+nksGtseTkENRcfhgZdI5bhN2U4fYm1Ri86qsV61doZ7y9LGxHlYkGzJ
GpFNcotFk6uKQOpjA7FJx22e3tLcwTYIfvEHjATQt4Uy8YNPrEhSKOAVJYVHZ0vI
U6xaOqX7NWnNmFRCoLWZ93jxKIjplyJZeFDfzJH47EKSKE1OXD521nOene77Rw2o
lOKNZWjJNE/PhJyE3DcdVTKttIzokZOcx1TaD1sF2PP18QeN0bktPDdZJEYK67HJ
Y7z00A2OaFzu8vPADpkNRRIdsGXSiBy1Nn3MDM8q0+/jXGZqt5btKoqEm/vC6lL6
zjdRbIIt5ItWFA0WAizNzEEpvc/kuP9+bU8TCVYurX9OSR11jMV1xFv5NFDKS1QF
qqz3ZIN72cxwJh2oREmsZoxyXOmIIF0EhS4qOp5ms/nHC8axVTbmjY0G7SJAQat6
rsFzwR1IXj7PTJfiZ5K43v7b2KaLentxDl9qWWQDGTK4fXPDQQD9YFiAosS8L8HI
XF+uUvvFp2tRSxkBYQkwlKxwS/KgVSgq4jUyEBpcerEdQd9eYaR/NXtRBD9PWE7s
zeKJ0Pu61rMotWLENjrIaDnBJ+l4NnzAIa3FUjDJkuET5zaQVnpSCo5LYeJlou86
w256894xHxy2ADaevO0tTJyOPK61nGihOQZKAnvvWuvkUNCe7DXNMrZLTFDcZn04
d2PIrB2T0wuq2Q2qrfoVTmMfVG0lg8L/NCIh17PhWtXoCMt229p3OVSqU77Cx8Pw
TIoOfg3968ntkoGX9Gnc8Z3QEMZ12YrxMqWKp1rTkRa22C2MK9C8YiOj17eznoEw
3nfQuz34zh5jqzErTL6NyTvr0mN0gOVmsjLQCj3rwBUK4mPbIuUmdbI0hSuoeUF4
hCUX2OFlScB7JJRpsZoRsHEuAJB2s7i6B75jaAggROQwjxshLeXLtuREGMP98hqa
1REcpsR8u4mEAAnnZZMMmVUrLbuzsL0IyIPNtAkHXde9hgL30VSZO/qFWGtSK1vb
nziUG7kCIkrctPuRVH7Ykj0iozhUqeDJkRdgJxuGqAcfmFZgGi4uKO8hG/yd6YQ+
GGrIAOstT0wBY1qeFCDYRfrWkkNGbKbDbU5faIjP/hOavWAxY5VrhrSjq6BIWZvm
R8yv+WT4VCKB0aeHabfQjElQWJwJlKJK1A3LGpmWHVvgBqRR6c/FYydF00nWNJg8
7EnYFclhJW9E8pZ8hkGtOerk4wtHb8DCo5FsfimWT+aNob9cOjC1jIL0XVrBp8jJ
KMlrZCDix0KIs90r2lML5OGP+S2hIDC9C72R2odNJMa4QDWysI6V+XKScFzoaMAl
6e2FBxp2ICsRqihiDI1Fsn+5XVmYWY1ig7xwZp0iK2wHp65YuZbMKBCIAsTEKeAs
kVPapQXjYFZf/KtEvZ1wBdDgL33Fg505V3ZMulv9X5lWNm4t65Eb7s4muyUeus5h
JLN3s3IBtdwOCEPS6lGVhd33IX4FVvsK8THMMhjiJiUkXTGT0LvpXwARO9N/vGTc
ixBSi7YT7SkDZKN6AYXEDFsTqoapHLsIcRS/C01aIywooWyXZZSyUcG1a+LthGJm
P7xUG1TVbc72yvhIMdU38MYXke+mw/Mr/rriZZCSoOl6qWF8c16m0K/iFm8KP+BX
MmTQzzwt8XbD0AAgeGx+jtAvMQh8bbPdByXUGm72vJmbRbTaNFvmSTRJtMMbXguG
Cg8to5ok68tJmmf6bpeUvVuheqj36VXqvkluL4MQOQ9AAynBQHClFYD2A3pQEPgy
DJqFuNdwETjffvwCgY3Zd5Dd0U/+V3oAcbDlSV+VEKA8DahJcztV8KxHSV3Hf4bE
5A7ehlZKRv0ORZVea4NlLhFpi4s4BcuN0I8uvTIy57QdBnQbpuiavZbRg5AAV3HR
Afzek6kLrNO0wh5+RYBM7mQrp0/9A86vG2BsAg5foI1ovK9HBIEgHHlybcIAfqhn
RsxPx8WQ9M0JWgmJVP0JTa0QMYUw4dnJDC5xdoyjHGBJs9U89TE2cnt97jPS2RAl
xKT5QE/7JKMvVLoi0/Tq/QIbxnak2qP72G5rXbRktL9CFhH+SNtbIr6djyM9ue3F
4ianm0Do6ONQPYuQK71MG404kLBiWRJ9S+lhg7o5X4JtNl3bx8P9doP2KzzNXBRs
l++1jIapKJDtp77XrHEJz5nBf9GvjmHCSbkCaQ2Yhu/UYIoWRFVjJpCl5LuwG1gh
sdajVsz+ZcoXpTVYPbhjUdqtFt3UYQJcBIEFkK+zCnolitljB1w0F0WcQBHiLq2K
BuUDhLuoc+VfdeQoo8j1hNf+5lROluynAk1fsYQquN/B9oIb4cG7R01mM92Xl0Lw
XVeqiMqbDj0BLK0f3S8zENXzB5BdHgIb0x0nb03X5wRRGQuZsiPqaAVLDnBHvZrt
Rp+0diYoREb+4gS7sK3RI69TgXZpQkCmkAR4GS45jSjEBVVn8YJbpkvIyuvKQcVx
Fv6ob2StoT1/23NBZZUsYoAiKap2Mv5b59VpKNM0u85YudonOWdju1tM6qzNqRI/
ciahN6JS3YguGY/ILKnG+kE9WNNs5XJpSLhW4aDOfz+85GH5XY+BAEV74T+w2nhO
z+3SSTIctAbPklZhg6wQgaMo/No0YL05qm/PM3c7ikRC5Coii/lnZDg24JGG5L0I
oZo81eTDLJfoMwyQxb3N6taS+m8gvM2CQH1AoaopqqT3ELtUt49Cwph+gaUHKAxF
XIkzN6OFFgn1vgGU3rjeT9dwgntX7i7PO7yMRMPa1KiIn+N7LbZKH5kirETsvyPm
/kWITA6R7/OaGFVb0CQP8AHsE+m+qSf++i6iVp3hfOzlz46VPLZhRDSeYKP/qPzF
x8yfqXOngzpHLjvdkQ9rbnvp3an2JVnRBvHECgl4/G+L4Ov3JsP0xCshQipDx7sC
Phws+IW1JDvFdblli3LNPnd4pHWcqTogKjEmHi/Q1YVvxmj3jUEMwAB9Be3zcKWv
6MxE5IRMlKMmKnVN3cnBCqwnFowLS2eLLj1qdM3YSDd+9wmSqFk1ooFH0JEzZI7L
9TrB9tsQAXVVqe0+IieA76i/PX+FRw9b/Ej4qX/j63RiQeOuETIyn2hZads/Z/zv
6mbS482JZrEBILi7PEGFJrvTv6D9lSyxKYbDuQJlt965XCs5exxlI/Q3hMxcNylO
XJUxRnkX1FOUZvVQP8Otn+5moZOW/5QrL6+QPK2dEFSV64BVmBf4Y+mD1WaAkrD6
LjXcU/0gvqx0HgKRdhZ1BYabikp8F99xhzR/FNGkoYkqDUZKJhqvvZShX7OWyC0i
SjXo8o2yagyGMx8pk0FQyy/W5Uje6zNlgLIv6W0XfkHNrTFutSbz3IXVhjD8bABu
+UOTul/j9a1KhuCLZonTkCPoyl8hI4BN5SdzhN3hnodIIe+sjLH5Qz9fntMiTDV8
Vc7S2Y0VAnR/9tj4lXGnRUDLAMeakiaWjuxlTYoseC0PQ/gplWdL6UHcfyx72tki
J/ZCkKaTP+nFf6prnz/oBkD5KrEOIvwXTXP4F7qsJREyWfuGT3RP0YrNyU7IT7iI
MvTTUoW3x65xFXrys48OO5MKUCSI2Y7Xgv766xFzQ9da5UW7CSwbqWDjEeJFDwb4
VaW5n3P/SrvuCqvnxfvElnuurAU6LOfZbLzZyrntoKJ2YN9XFNS8rUUxjOXYJAmP
E9aVI1XoAYGSp+mN+Bgs+y/s/6A60x+PntwHRUE4SrTtWCttLsEYYKJ4I8JpUgtL
42pNg9UWok7lrv+L5sTCXkVjeWZcjv/ZeKfPJoXobwkjRFzgKoh8aysV06nstUeG
2WXFZGfjjAyT4+9KxTnx9dH2qcRGjbkxsn91q2GnCSIQcMUk18ebcLXYgdXglknW
CClYHnkFnKm5/L2DPZeKF1ibQH6rXmCgIzjhw7OdeReHGCMev8L1LXWeOcIYO1+u
XVeS2PnKSTKxXgRktIKYAWWk4U2CKLHP7IU6RoFHC6PDSzS3e3LH4yixP+q5rN9N
AzHzqDVQ2YTMFb00Pc2JHCYkv7gV4lUTJQoh27OygB7Yk3CLqqyMzgbR43L8WvoG
DNlPGWTzf5onWk6NNoq0SE4HoY0kkQr+yTZ/zQeeR80Vm6UhR+KjuCd9Bjq1T3yK
iymte0krOQooKFH+aQDdvrGWGfKBKm7gMZgglqbQ5ABmzHmZQVBUEPnbYDXLmYHb
PhfEplLYGVVTRp0y5DWJedHS/cx1EsB80trPX0aVbS74mO+jRTZWOFwOExtoNz/1
bs8W+LGiJTQ+GguhCj7akOZZebVMBCQJv0cZ6f4pIWSg9LrGrJDOxuDY5r0CWhBK
IGMsyEiDIWnCQHEGqnmoHLpGD3NqSnAzjt46RihT+4Yj4sS3gHI/S6gzhSmEGAwR
OEy0iu2wrwqQg9lLbSzaSbZXrvySGaQ8iVLKjyofedRTdCAaMrYz4QZtRk8Kt6wY
o3pZ9K7sO/CThYn9I8zCpCEILkXGtAMk4JV9Xnnhdl6FkS/KY7BLyE6vh5qzcI5k
rXMlfR9lz1/L5SS/1ale5YurocRAX7pA5pA7JXpKYHZ1BBwip4LmrFMM5YqGVdbv
SKDw7lvqApH/26v1hPOLG5vS7bqvwfScSJukT4mFL0//xy1szy6bzZUiOzaJ4dF8
8t7CGKYOAJl3IRneZELOtPmHGK0hKRzTTol4Ax34zit1Ct9KFB5bVuuNCsiAAi9+
1wfNKCtGJh/bdTymgoreNTsDynGCXLlP1gp5A5x8OdFhWTdboxBUvQL9tdvBcaj2
ZiWuld3vwswtcryVXHTTYSuJ5+8E+4iFq/DJOScyArEGjemlzqtRzsMRCvk4h5oJ
ra5a3I6OXBzc77vIU7E2Xwzlz+vmt9TdvGiBe1d3QvBPKN/FeubRnG3R17JaW1Sm
BpKPjQgqCHILV8R/9xZ/dAgHbZ+d8v8er6Ir9xFoTcXVPGC/owgLwxfJMZj75YB8
xDkMbzaYASqBR9mokL72rJ8M5v8w5y3I6+LM4gcymiQ6ggfVJ6Ua7swf7U2Mo4k6
uLsP0AvbcEInn2qc+fKEbVWRELaXqldC8EpuWXU5XIWmm8o9xpiSJ2jMnM9KZ3de
NDmYzgnpFh4iIpIpw7tjJ4ODNZGgRvrvdhYzSZi8x9GJh4fJkHSv5aK1FCLORcXi
fG7PDn8Z0Yy0iXU53OuIkQ0XJN7vkUIUfN5pTYADBIKf8SzJ7LG7xjxSDrPMhvLy
TKwHlKX8A3AESEe7JgOrHgpGeM0xyEoBbnVav2ikQqdXtp02AGVb8XdJZqy0fLGq
CQtzNPukZO6Vxly5e7iUW8XSzGEHbhcUuw7hzD7QCFEFIVz56Xf1xiZTja0Y/CCx
IR3E36WSuL9rn5dmhk9CkDalK4GCk9GhuCsR4YFClWUJ3xNMCu05FHB0rFOSbiNI
ZhWILC8P94YasxAauzz0y3YKo3gMLK4VlkFP42QpiO8M4X95k/cJNHX9xDvoEtA3
x5pru6dpah1fb4i/2Ha+wDSBJC2woAMz/47/gHs4mZ1YwXPPeOkNO90R3902E3gO
lTf5frFh21ZpziYf89/MFbH3w5lTqx0H38nbyTG1macRxpKK8DNf0rYw/es2bRb1
2RV3YNvQW8IK+Q3OVmS7hLUZoQPk3GBqXP2/+UrbQRpnxso5zb41gaL9HGDGszq7
jpnMjTLdJONwUINllN4tPv5weXOjZtwvCk6p7BkIPWw53QokCIwycKUV0dP3NNfM
fVivVZBUQs1qau5a43wIw0sj6uRR3+AUUngB1nvCeUzhVlzuOTFg68RjmDOzc4ts
lS0m4jDIU+2SwUc276zApdit+33XaA/SoSghjnT9aVH/HihYNftj5u6S5wOJb+wx
YZCz01Qqs2aElZdk5K57h0NI1qIeC2LECaoLgmbR8paBAp1NPJFE/lN5ig5zGukP
kW+YnxEJ00M4GWH4erTD1bIpeJ1VqsmSr7+Bo3TFF1kTbloyKrb2+ySZ07d++orl
2B4ewG4EpbPVo9APQF6Bo12lQP5a1BCtKxhiPB4zKgtWbuB0yfLZaYqfjN9s4ZrD
jKElO0wxb6YMjSmEWV2rcAat6l38ERgmJFhWKcfchN12KKfdrGMICBb127Zt3Ucp
ZxtA1dDsD0XPr35vq1pWSxs4d+0hPiWF62po/mhrvHisc0U8C1GuT+4GVtjgidul
iEq4Bq3i/wJmblLUpn7CgpyUv/sDgBmsWcS78nHAhJ+Xh9pdlX4IbzNGa+m6qJVI
g3TwpWPFK+UIA9788dvOPZrtNlhELD22bS3jjDSOvS6eP2zyqDMQqrIgRuLJum84
/OyD1xi8or5hmXxTbjq9r4lFIcWLJbrHKkKIu9fZaIuaO9yzSmQlWU+W/rNrwryI
6Fc5hRv2Jpg+QNS6hD34jQFDYu4X2H0tfTC6M2xMmz3JWxtxcP6c0FzRtsHkUXlB
3qFJsD7XVw6gjb0JqzjnCTyBosaqdUidYdtV9KvbrzbNl0F9NsOm8nsbCV3Cv24E
9lOIcaRhfOMycHz2rSWyumU8FLa+CZDcdxQpckQPHVckhuSbRDOJN9i+N2yfAdCv
/8X3TEWNkc4mwFn+40a4+/pLPu0ANI2FrPOKpNe0oO2UldFWnWVgbEIg0nyEHP+I
VX1Nm9F50AXHGeJJiWMgJukymDnFUS08hvgF//rSo5QP2lwFpHokcYVRQkl3bXTr
2MaJrdHmAy9vokkotwfp4IYAUeBilTUWu21DoBUCmidrsiQ+Y9+vZUDjb91T6Cao
i7eWQA0PvzcUu3Ncu0+bj/v6ROJFlfaTYjGfgK4+396fAE6EHQjq9QbRd/87vQ2g
AFb1gXNXCmzp7Bq++6ZELVWuw6ywt8A+zZzO89rPrcWw4b5eUuXj8b7zuOssFV72
gWgWJGv49AbFXuAdWJKTmfyXcq01gk0jYFhrtb9WkU8oOWRBPYuR7SjbpBfYWrg/
XW4wgb4DYhhTnbumr0nJRd1ZeBSI4L9ERaZJhsJVPy6MdvqDEVn/6xi0nK9fnjrK
4JfbVBoNBLbLx1Jk157thmXDstTeQzc5S9FcGy7GRd/nGxASEhsz+wZpByH5+TsM
YscIxFf/4UvHu+Nm2+bekmNRElVxEBkK5EnU8GF6WBPP3uWlIMdPw4sM7VIzb9jq
cqD7mz+Yt3eKefvEz6UsBSr2DTDGd9mJ2U42uZwJQPoNyFT0ldLmXpdfkxfIgR0K
CEo5PJst7WaZPWSKtgUJSbWp9nZHLYIVYog66XbECY/pdgotcKgBiVxmgu9UFo3d
tcErmhmNckvDtwEeHpHij70FZHQgPCY7vvte8Tnu2wKtaTYL4gAIJ34FIdWovrqJ
BSs6bTg8sUV3wEyvTd64T30gdZOnZMcimrKYQDbBKm56Nxd/BHbjnfxUfVmNQl0H
JexdCQuuVOOvbaglKaZCk+EU8VMMjkY3e2lmtyQ5WNezlkCyc5AHUs2Qf0Cw3ARn
k5UW7pcuZmq2dIlG3cx5/75rZ/QdgjTVlUQcNFv1uy1JRa3nk5FmiVTUXjvFVzVU
GevbzCcRyU23ffyNOQhfW4V8pU9D52pdZtL0jeEEGnTG/3l+MdC2XTVLvO92+5/I
7Y9kZALi4RJJi9Gdoh+LCJo5Gox/PxU5rMSqJh2RKutO35E2npWF0j8CiHUqRd0n
kmPpCwAQUwlBtqF7faMWe/N6u4CDDXHIe+sIOuHBB8hVVEC/4Sd8oNmlSkWBkadx
nunNvC5xit+ZjqTICZidpafEhMk6E1GXQyMAk+o7sQE3pEbKqqao310/7vdG76kd
HsiBDk+bMtFnKK0GmB6t2knbXsOjl1NztSWvGDYkoyJ4w9B5jDYEymr+ctYao+PS
FyrwaTLDUlQUjAGwfE7vERSumlmQEQ4zU5bjF1Xtzm23/4GCmsIaeD09zr+ln1ao
U6G7Oa1Q43b37HC/GIy5aH+F6KysTg8+2D0um67yOKu9gKh2L8K2UG4H9oo4u5Np
/LtrxnWR1WcIBaXg0I8ehcyzve/d6BoPWd/BLI33P2opeb0+ypKw5V2bB8hf37vQ
Ni/Cc3dWXHPdPUkYi5kZjrUPHgufrFPTI+iQLaS5XnijwegxJ0tZj9OX+gA7g9Xx
JirVGsyWCuduGkFHwcVF1slNtM+88YqPeHr0g6zcMGpqChNqwVJhUZfhFd2vsj+V
zv7j6ANbgXc3Pj9C42GuYE1B0So0dmeL1EkHacdkrTcm5FqrYeaoDLPB0heXKrnk
GNzqwB46//JIA640T4pQOzH742KgthCKJBzhpS23uQLdksznyWZdP9WxitLCOPnD
uVbsGf1GmtmpkjKGZETKVNPX/cGuXbVp9WzZ0SMb5EfsWEv524zAEWNUnaSDJ9TL
NB4D+NnFhbJHVYz7q9uQCJ611QYRmigLqe4vUu1XytWl/aOnayVD/O3wlDy9D3sM
C534YbnUaSMbRC0ryg362s9h1CBO2RWonzQj2Ol/MgCkrIFOWdvkjpUT7oNqcJ9j
kIrKsfRrOZ16BVpGJn4fiKQ+fk0Zm5z/1itMa6B1Y5J2zFyVFd/6Kp0sCzfgPRPc
/04V4wypR9Wjq6B5lcGiLuLcYOJP/GQVTwD9kzojU6MfFCS2Gfu/CzxuHpcjYUkG
V2JFoy7Pm8uzzUbNbcS4VYGiayRrP5lSdAVqjne3cyGjU0cA+E49aVIgyvUwW60D
vQso3GDSfvqFXwGLLAsJgigZVUzu9CqvVAGRqikg4pEmKqpFPkyEy0/5kjSgS5im
XCAiN+yPVGgag6h2XmB5xYKj+ien27ZdZK08QWTr2KncQPu3VTzqgeCV2Kmutv2W
nub7ruuyB6uytE+svR3/teqHkciktaxwtnAcrT+V0Yj9tT1zxHNNqwoKBCBD5umd
71jiW/gy4Uq162oxRnHQD1pgfSjE3DsJ59kNGnD+V3AqP1OygE1xLg6zDn9g0O7g
bt7LDopkPKXM3UGplj60UDQNtlYlNQ4YZQ6H6xXV5c9VX/tKudZYF9PTzCMOFvJW
YcPNNYf2FRdMT2rEbnaZBKzPrD5CTZMg5fHDbYtF3JllCQB2NLG8uf6MuoFYRRBr
U9o4RS6SZhbx6bLCnZ0LVPEtkJuprqo2Bm11aIL3VPZAkEqpaAP7n8k0NLGGdQYL
agBS1QXO6Brxo2XdrJcOc9T0MNn30Z5ixFwZr6aXJGNTUbSeROcGRbko5GR9XyDO
nIwku4mBoKWRwv7BXT5ERCh8Fv7b8hqw4k9C3H9OrFMNessBuhdn2LpFU/A6NCjS
8U+BTNpEE2Fqbro97Y2dz5DQSw/Qgi5/+rdUm8H1ugQWYz52p9Q3JghW2aApBvMh
bYuSLpMMV9IQIRyrGcht93lPQW6T6vkCTRjdd7IITsNKwHOhFYrSPpMFGJvAXQ/I
qG126Xgx5PVpzd7AivInV1eTLGoxKcroGaeFdQgzNsvrWxKKEU4of9ixhVAto2zm
gGnTg3JawkAg1P9CD2prKwQBAS7utbzwcgAWmAwH+dLurGzWf6vRu7Qdi8VA+w5n
y/lySQhZzZRpip4dLX0yw0DNNj0FvbchDR4nnIP22Ij2AbTS+sTH28LuaCK7zC6p
YeegoOzswHNTEPAo33vBiFIwCZHdUB76MoyeBGVNNC9gpRzFnEUzkEEnHbXjfixn
ev2sdjbHVQ1T0Wf61oJoI63XsDNVDHYGu0Sx4HLEvD4Sy4rOXwpOX+Uhuhv3S9tu
g5mymNQklVtYs35JmFq3HcaYb8LuGP4D2yCh3U8PSPx+pOS9D0qFcz43y7mq1pPk
N3D7K1bqVc2xVpSzaZ/6YuhaGln4vzbOoBBvKAc6NQ9/3E6Qlq1hYcH/OfO6XV4G
q2Abw3nNr4VHfjfHsCn0S+1/WL5BdmMsUzyDfu32O/V3rfzPRe46JKwAzbmPWMnY
NvxvT7vDTh1NRo6pOQaAF//NM6p+bP30XHBfVHCzQQH8E4/PB/oS8TGub67CsfMd
JX8krFPtEYwMyGJRO7Kv0/rdp9u6WuCq5ANF2tlBFoOKSnpvWPu2qZRV5nUyF42Q
KOES9Ea9ix1lu8CG+fAhPMuZZniMsBBRU3utoeIgdcjyLMml395HSu+mgKbaiG4E
Q80M4jS/ICf0Sad49eyBGLsIZCv29HGZorh3DBBl9r31Hs2K09JLe5mIlJ4Y03d1
RHcHtxlic3kNpXwGKUtfQ3jBCvD/Hrp6eByrbn9nARc6sofwwicaq3RkMO+4D3R/
K65WX+1oPSWLtbXfDH/jDwTogqHmTJBWFv+ZfT3Gh91LGqeiuxz84XHs4X35lGw9
sKB5sdDhRVbYjPnz0hWsI2+0to3jhEfEHYc/eAmoP+Cj92eFr3Nq3LqcdXqfyRES
oHhrafO2dE3dyMIYGj/2wiT8baEQAPU0BQFUg7hlrOtPJLUrVPoX2gU9gquxIKr8
2M6MLGMCwmpi8GZ2v6sGWg2I4VGaniZ1nY7+8yS0C7CE15M8djOvtXiVUvmIz6m9
6Q89bAHimacrYH3vc2MzTqmtHIAV9P2pNoIYOlGaxtGuoVPFWBnqK4RoeShYpHg+
LU3fcsbZMuDVI8j2bqSOWEkY+JuqjwF7ThqzIB3PcEJbG4jZPEMjY7VmlIYPrzr6
zajWdYjeIloh9Vl/n0NjdTPqcmeaN18HFPgxNEjwmygvoiYAhQPQxGwYkYnMQux7
SfRIx0iHP3jN+wvZaAikLnReixgv+qW629BMfw1hpzwAkZWTYC2jeONlPS4NvCBv
l03AA9C0q/gymx70O7kwNuud+ijqoPhMXysL2ZnaLCGr+65aFAUomlHzNiCHKXwQ
DteKNSLMqOL+QawSh+1iMZy5AXDQQCVLNhPoPeac0UsfjRx1CuFGge1TP4Rb33cZ
+A2Fqg1UTYUTpA0g8R55HsM9n8QIMeKx4c6cOmj39km8zMrCwoSOjHySMn+D2QuL
y7vM6bf2IQJlr1hTOt7CSs3fjxOSCoI4eLeqWJFpgE9aWI6W2TkCuBRIJN3KLWOf
PShpPtv12SEZvTeAprI0ZNITGcO80glQpXvCR/+F5/gC4CJA7luDBYKQC/tQgP7L
4dCc/Y2eiUyVvcaV3finudaF/WXPUPw+bqz89sYHVDGVRt4hjXIzHEYP2tMOyCgL
c3DEGDlPzRsdQsitkhL+n39MCkFoGQ/WrQQFPkjSn3vxjcvNfqlZhHp+w202IWAd
M5QvYqoMMXRsQpUPVKH/A7dKg8DIffSUw9IPH9vjSj8ujbtZFWazViPVFAT+Ug5k
Z8sg9WQo2hrVLH40rO+A9ZVsOTZ5dhJr9OqOeKzmunhZCpsbU/f+TtiyN/1nuVMM
Mv9CElsCLn9BbcVLM6r8KNs/O/k/FyXZ6JiFonZPaYqIHI3VLU7r04dlwfrXzX4h
/4n44l5BKECoaYpgnGmkCVmFuFA2Eie0LJ2JdwkWQD+gm4wg9ygr7uEMAofuGWYH
UUofosjndfK+/rkzbPg3jNgKEW8vhlC4ons3yUASvKN+P24OflTx2ozNJgm7uBsR
UOmCw9T6LJGvgVyIwKm+bhKj4mhrG2wUunxaBVYHzxQKHb9ouUxrITPqCFxHksG7
yun5r9EGtlBmGhLp3QSLC9iSAFoRl57gbAc/j4WHqSq5SW6jgpAAOE9HJN8Tb19S
+P8v2AjuY1yst+eVOefSGq0phTEVghiq5/MJwjgRP4nofIlUwgdTcTPbxOG2tRhV
Yhn9S9xaEGmQgY0jJDOU+D3x0SrbU6G9EWgv7daOmHVg7Dr7NFiFwO9N0vJI6gKF
Qnfs0+Cx/q/OQRPHYJ92HKIu/vHgyCP2Gx6Ia7u9y2BFYRQ0HvDTuVZIaUHsr17Q
R5UyvX7NvdR3KXTqhNb6osbofEKaH6xUd56ysF2WdTwvpzoIBkHwfjBSscSFE5Hl
lnoo5OeQ3kMCQrwsHOnuIfM3PxiTHyltsifyZvm3w+6dPDEP9C0ry9bUBkpwAbmI
npA7dwAntGkUH/mjdnQDTjqQIqWRT6jEN9FbmgVy+k7RIiLMnmiJu2sP8Sf3AEVn
9G28xI5mHmZFLL755RVcrEqA4feQ3uTVY7QU7B3E1VhyqgXhS2/YXVmKUak1gK4d
hfQZ0IYXAOCYwqFmVgmeIXBnPwjZ0IXIllm4ZJL36wWI/8PruYRoWOHNuBUmqKht
RrvWkjbEbGETX+vzC7qwgTYPGsCjaLElSrgRD7J3ZygOrOhCRZ1R8YurjZUyvdBt
HCBDHUbsawq23Ke5S8QZqJTiPPxuHUKRuToxOZvD1fr5os21GM2yq+h4n6MbS/Z3
eQl10rt2+JEuXchPJUJBrsnzRadqBG04d08CQ7uiE3Mq64CXXOqAteIAWOCqjBkS
iUVVVUI4Q4RJQyuLvOdqnWun+M/Ts8U5D4MT+E3YVaz0QyC7zV03Og5TvvdekeGP
lKAYg/AjoWsGCjBQSzNhqa9gF3Pi/cPmOhwgklBkCcITsuu4EiKn/QVMOfCEBSu4
sOf+lYP4US1ZYdoerL+3libErKgLfKm6XsLeN32XGlXbgBLqr14XAUztfV4rsQOK
r7BoquUuBvuX4wjwbrA5hJrrADe33SdVObs4+FfON0moQV7IYVy+2/Q1mRoGf4tL
01fFMxlzoYR9mv2e6iAA5en1/u0cQfPiMHrf7iA+NCNXCppB09Cjb6EBN3q0eRzL
NyiAHoFm7/SqTWc1QxTqALmr6dd/8BLQ0eSa0nZO7jM4SuAJO0R2okJeYGTCfUmk
1MYEBP8dfr3X2AXblOeb9pf5WQzaJ5SmF6/1X93OZJniJftOjwBcOPBEB38rWBw2
X+kF7xjvND2R5BJ5pTGlC1doji+6Dj8sq5xmvM4zw86IkTm/cA1NSDkEhOij9b4N
wJAK/v0eCAL4HjtYP+xJCUx1ZJSmCLsrCeR95TgUkxOidyohYSOOvDW4ZIABFdOp
jw6XkQAVNo2UIVCS0fqRfcO6xRohfls2K3kAwoRDX0BIZ2xzqbvi3AlRvxQKv5n5
GX0nk5mcgPJRT59MkakCvHcAVW/Df8zoNTsnI3jTm32ouAuHfL4Pzikh6E4U2/Mk
M54U2ljcakwGT2CeUG9CqkmQ1mSqnHmboILATF6inv1b59K/wcHJ63LR055G4jzR
b8aymhr1e39X9W6fTOLZxHr87sthD9vnuSMpcTmpZRnkZIFesdz0QdACICyPJ5NI
jaSEccVX9NpPT+XIQRtheuEvqwzCutux7I8D4M+m3R2TzFeYCSeMBwn6H9/DLKYW
2czppBdz2TTX6YIJgTgjeosLvVwY9vCYBJJqbzHpmz9HyHkpnA2gpLaZU8K0g1En
PCM4MUElVvESXZXen04WW3+ww1FubMHf7uVU/WtgIZhZZ/hF6Mtec7gm2EijkgfI
dShi9uZTho57Sf+I4qZCGpqvmSSMKeTceyRKoyvVhLXmBjRJzBLamFVnV46sN0mO
kELt5pWc6nPsyrBQVxuFRxbtb6PLAYxIc++tO8wfy4cyhXAm27Bq8AOlHm2LHbfr
/mMiHYSso5Cvt8i6ODeNMpKdkIV+ShYu5nk/B/vtkiEeY95q2g1EuzV5e8n2ASSm
37yDj1fG/oh3XHmCssnE0egshs/hVsVThwnSIJBrBM0ERpB8Is1CE8v+4iiRImnk
5dDwOLyG+xH2RJOFvQA+6KmxCPU29ikSugPlWhOL/O5Njo1W5DYgMHk8PT5Yno0M
sOMDp3Df+0DRyrI1/47N7vBrAKm4YVDkQSFV3NTjfgyuyMf5dsXMVYq9ZPiKWW/n
2/a3USGH6hZ9kEkyNUrg6ghrT8Q5wetleYnt9oRYTdNOKFsl9Ab9WH2+tInIke7D
BiFvAmsLTSOr975BTlWUHr1mCs7rpnd3msD4FClXPwkD/LQRgESR8Fn9ff3JraaJ
jeFwAd0MMLkkuXObFLqOwsHuBaHe5WxlJveD0yhQEb7tr/fyXQHaRH8tQKpYSHz2
OtZmvDlw8WPxDn5Qk9qHfGbNZk4UklQ9KR26vFG/bhhGs4kdmvx+OKwfbphCd31C
wx85JWGAtT+KsKAxf8MpmeLt5g8wcG974I5leGooZeAXCIVeXTzPT9zvVmaKasIL
/0yhhnlFCUSWPccINsakLac3CDouDIWEk9x7M3gRG9R2KERR2IFRd3pO9NXHdpj7
hNcmypzs9m6DruULCOx7TI7US63siXCxuCc91GYi5zAihfkuQKWKPFkuiDT42oDr
+Mn1q71gKINtqutQRxTk90EEUY3QUOri8lsJGcGmr+ef1u8T5ICzxXEwUTQKSMM9
NuRuDoYSI+06Fnvp8d9AC/h3FP7OkT33o6at4w3rRr/KbWarqdWvZLrQrBryqXSP
wUgESpD9qch4HauFCVGldBVWd5oqq6gk9dBTkXscv5op2dpd0Hgipotx+zIDO2AC
F/qW6UI/JsjqvCDY+Ar6mF6AoqgrvFbEoqOgxNQCewWl0gMREjqaFE2XCtFjbNHW
KvQvdVHQsHZjHVrVf6qQKFhM7AuD/rr5Jwc1rrNGp7OP61uk9c+bJ2oBRpdoXanY
6S2iX4b4Z3X5WsgthHtbblLUeTXsG6PW3rbUzGn5tb7BrxW5wreMidhgWgqIcZJA
q28h6rDrdpt324TmCFX8MPbRWhCue0NDhMsqUsVzAO8aWnY9Vsqc/rCv2Gux/4IS
24Hit2GPOlUHuJaLfAhJahkg4wnpUDqK2MtkixTQ9b7rH7u0F6hA1lcopvrqxbOJ
O0l3MlqLJT7VTcfyKHW4YHNRYfUGhLdfuv7NNfaMFyg73Z3nb3ahIPJRUh8jGc92
KhyFZqPNtr81eUc7l7uvifJ6OHJdNV5mMTGOEKOP3Kxbji5YdcQL5lgonS7AIZbj
8nnxyBTfDgu3oM7IxTi+T2KUtAG/VU7SOabvbFCXUFLJJfL0cnFLuSJrb6iHlBCN
ZKs1t/WRkjs1Gx0dMNZy/8A9+e5+8l0n+FB/PdAOrlJScbTFw7K5ceEv9L2VwigG
76Vkb0a6Mh195Z4BLUEtekg3gKhNARhF43iUtZFDhnylqE94J7611QPWEMwA58aO
eFl8s0qZx6E0KPc+jFBNEcoaIAZ9uxseQTmfLkVBM4rBXatcfDH1EytLV/n9nTKU
a6RNm9V0R5MTpwfbN3G1lYzE46gIwEZ2aWhkzWV0QF0++H155kNBdKgAhPEPmX77
eR2bwiX5NHGEBPml+4NYe4jghB+q1b1nMuYNydnIF5lQ43qsZE+7Lapvqp3Kf57H
0WQ3hAy4VfmSx8oC0oprAx5850Qv/gtFdUqrTkbUT2Mrsoaheu/7TUtr7tyuo5F2
6UkF2tf6Pz9vAF6YySYturXpMCUMX/j5gBdAWXmT3/YwQw9QTIoK4aT+cJR7R4d5
felts6in8YwL6Zpv75AE3rhv5ifV7wAa4koygYD/fP2bsos0x/c0Wpr8jn4Fh4EW
jpIieC5yNz5NztLKS/7VVby5eTNQyzaIvBLOIxnftniAJzcri4y8Wvs9PyR1jHqS
wwTP3ir/XJ8vaFpLQ/eujJEPylfrSP+IU2uxx9OPAPlfVWc/xr0S4ZqN5HSxBtZ/
uCO4G12dbO40raART00rjaA5GcJe9/19j9NIuC9enRuNsPEjgIbLAoTs9TarKd2c
9Hbp19zHfRVuvY+NqdOlewiqXG4TZZHMyVYKLGuAWAMNY/TKoi+NKwaMqGVqWjx6
J82GQtXV9IEST9U+ZKiHLw+BKnPq8NuI3vFy5noCUOoD0PSJNuWLlC+V7ap82hAJ
Dk195/yl+ItwhJZI+nd1Y5txGVk2zyHnUw3jtab8eGasHMMqylvs31nilfWozrla
Yi2QcXEYDOOzNfrJsstXEIhkf+aciMM6eIbW8og06tBR4HhnBip/jZuv/01kZ2BN
8eJDoY/I5jyd4UFst8f8FgNmsE/jkZw4BJMq82xA2LmXg7K5BUhf6QDzrf4jj3de
VLOl6SvwxBKMhfhpCtoTicZuFBNJhGzsHeSbtUX9O7sSRfGh9uFT280aatQ7kSCw
Vt8X5L9201HwIryJr0qA9brERnKCrmbKZomy3fgwmMCX02F1BpVx6j/t/Tnpl0We
UGU/hQA+Duvrzt5IGWZOVl3TvfEExbNqqYUeQaDy9MSDSJUyBl82qdENIbkwk/GC
v3+oS3LemhxUcPC+SFAhSQfydwztLE0ZC6FyoZm8BcYxQp+KIiIFknPWrz4lJnP9
zrKXnaax8bf5DbgGCCiokbNTpezS5T95v2ouk3ztt7pJDX8A469V2FQX7kOMeUFo
7VrsJJ5Ege+x0r5550pxZ4jn58E2WFYr83A4z2Hg4H0PS6FqEKE4AfBOy9zS5Fcf
8cZS0Twi3pbfI/ZVrezdNzY+C+e++h+Lo2RFwpYhL/errEEuCpUkJ3RZtxx1BGRx
TGWQ2Snsvb/0m+EtV3svMDB5GWPB3hpbNFtt07Ii2+8fpThmHLd1YgDNVojBVPLn
b9Ijb4olem93M8ts/9VG8Dgi9Uw6Ry1RAAMAcIpAGeKGXMcriq7zkIS+GjFloort
lKJa5/dnIgbtS83IhLn6t1aD/8HTnBd+TI+OZO5aRBOuVto709o4aqSgJKQHZlfH
bcRwixNHayeUET9ywsSBTrVyfobypWJhJK+MqWCM9YGDphc8UWosibxQBjhYmKO5
0dp9oz37KYpnpDPh6mJcJ4KQh9Hg43NsmGFUlOgU1NVT0KS3RE2Ti7+7o4rqeqvP
MsOqng2GG0AkXCW8wAjIkaRDvNIhK8CHWFj7fq6R8gbBzXZm0dDmyIaB3ohtBk4k
fqCDkRK83wkhCtsawh9Izbe7fP5ge944m+8H+sYjdIlMalQdrCMuiT4pOmR4n9vh
k4kd7rJd8FqMsCd4c3Rx5AF+yEAjCj0gnCQINKwQ9+pF/VX5a3JvL7E1Hj2TGYjl
vmWij+F+z0+2txoM6iHo6Wz+aa9LxumBmaWh4F3nizsSMOcOaQTsJsDkiRhaCg/l
vlHMis3r78HkSzgb8WLxnWpJHrUX3ByTkO8hgX489Znp41CF4l39IEPeUt9TGVHr
hnWC1jiffdVP/R0239/igjuwEW+NUhdqI1DI8u1tEtlLZH/6Mn/fNmqK/JWtpMGb
y8EOoixlB1kI0szSN9mM9BmxmFUE+/BMGDW7hx3UffawInZXMVG1sFc1jkkQFZeC
XA5Ezb6A1kGWGim4EmBI/A5qpvFLR93Npt8KzG7HoQ3bS1NJwuPP2hkH4LTJaj9o
5JlcR8tFi07Z9MJEKmfyq5gY8n7JNRnB2UNptMjwyXMfQ+wPTEJCbbAr2ejX960h
1QNvk9YoEu20+Tko6ereFY4XWIK+jSmrFtuKP/bLwFOg+2HJIyRr2tMyj8Gi0x+k
Ha57322ZW/EZIzizUPw5Bx1BIiZL+Kr7tCRtJy33xg1aURLZyTYVUMiNv1/v71OK
KupoZ/BTdUbIds+PRrP8TjfI+bAjkyqUF6spA/WNQdDeagmTWDyLNzXqEQqIGT2T
K9tadPmgVYcRjjkuD7l6hodt5hmkc1XDLHeOEWx+CNzXtlnJSHqF5fSShSPg59ty
j7UJwLZM1JZtiX2jNZxbmFe61YU77w6P/wCGbkmW1DL7IYiP+blrWSCeaFkHzqSc
1kS+iahpA7bjT6k3XjrZdY0p4BG3AlMb0l4bWwdKOTeDwfxIO2/hPWEo2oLHnc+U
AxPTx+zcWyyrAUskMndDYKhNRhTZHw1XUZ/v4FnuvC/1xKkOpznKS3vUk99uWEbS
RSnoAOg7Qt0m3NlhyhGBpIcpaONgED9gd3Tq7fZ2VsrWzp8nUvWghzPH/L7vXJey
TeijS7Eu9reQz9dlRJmW2MTC+IrqBs9xfRKixmfySfUPMRuG6iOSmXMgKxItHW/v
QuzIv5qU53P9CeazOda+kxCWXZpI7xstFyWEfBmA8hhXShJTjJ8jc/ONfL0hWQvh
QjYjqrOGHAuonWITrLi+YcN26oQJHUe7w6hT8FK9NqCV4uVpC+TAzu5ahFQMUuek
wun8UGpxCWrtghI1kdIX48HstwLgJzyqMrxmNDWLS6J2BBZB92dvMOITgewZUsKg
YNhPkB0wkM5Gb8k4ACANjXmohbirzssuXX7vhIUEFjt36/AQmTjExzubhvEE85dr
xNqcG9Nn+PHSIXWU5SnX4q6y5HerVtzTm+uDv4sao8BlqbICu6Rq2THTcD7gUWg3
LXtYmv6bbXuJFfYTter/NoG9xjSqB1agSrQzT9/zjl384dSi/xaVskbSe8tuEEFf
f74xsyuQVGSEJLBTY3AKfsLuMv9mNEe1jS26B0TYa6D3mf9wUEdWPTTLBLa5xAbu
dG8dkOPDJgWT1unJjnQKSrL+0fw1k1jk1UVNU4hVdYXEfMyuyL9hijzNimJj4TjJ
T/rFyoH5VEJ0rrbPzLDKGG6bCK4wYZd9UVjkhA5+aVUCjNdZxPGja/sZQgWS9ED7
NmaSeU29wejTHU1lJQ/f7rdD1WATpWkeD06MWe2Mr5EfTib3n08kN2PATFw/FBNa
AYNCg4eJrm3GxuxcOLU7+6sbHb1ZX2HUs5IJ6mCXcB/MWrhM65aUVAMC7jFN5NPj
p00p5gfHsYLcRxbT1q1n7sOF0ZscKvPVLOvncLu+wTX5xFX3TB/a4SZsNHAVWdVX
sea+pl3yPU2xCEurNWfNQ/iBqufbHrN6rMj2zYs47x4Dk24NS+SyGKiWH+7R9soo
c5IddKctEaq9FqdlgwTbe873N3P2kQTgbU50++nsKqCykOh3cklvx/mwlxWwpMu2
f/Byq3C1xIzusJYjBWKOAbVeTAIIOUX/lXUB18aM7zoc7CUJT+nHoM8QE/MSoP37
u0qH8va6uAn0NAQ1+TMD7DMM8CTDFHKKMUWuLrVhaUMtzPbPBpRbdGymaYRIKDMV
N4pielcgSEfW+pXZfjJkhPYOLbm1zgUTiNArnWpJaO6uJPnSrOJgPfC9Fxjw72/7
sHm0bpBX7VgYjhmoYHYs8+MQZKjMj+Xwj0ae/VNLtsHJoqoL6C3SfZpj1kUb/SIZ
b/EdFQDMeo182a1cNudb4UxVz56YR8IYM+EcB+qh/Lk6WdpM5l/GnnFi88KD64kZ
h/xpMDHTDRUuKri5gq6D7kr4lJR3ufo+vb7Mp/Zo+JrNJvRXrNZ31ZhDDQjCs8HJ
IrkzQS0eF911aWxwPWr+n5N4gHufGhb5pj/I4Z+b3/5lzjUIVkAtD1PxjbRBK+D/
EKgLb9t9xJQgEAVIUqBKzRNxvuJkB2PtUBBf650Gs/jybJBfYij4lg7msPEIGpri
f8uAkWafS13DlpfFTWhxw+WlsmTnOA2547pWC+iyr3/WMr2BSE9do6uMhaoNceLO
YKPZurVrTsiWUvzZ5WDnSF0zCaV8lzp8ICqkdsx6gcksgE4jgIOH58kDT5d0F1rs
nDNQTU4dCM4nMO0ONoFqaqVViOd+ILtmMKoKphvEyuqpE1rwf+Et/uEXkh1xGGXq
e+3qvqwKmLdpsm3VDiE7mDifiQ3VMGCId90kEF7Ot4tIKGxdT6SZ5iDekzfdNMN/
uEC/i8tuBwAAHHIJtoSAsCZS4lwzVjU19ekTWtlOuIGo9VqD6s9208V87dfqGtM1
YvqN4BSKle/Rb6r16H+u3OmjN4tTVxdrrq5O05RyI483ip2g6O0nAvNao1rAJvA8
a3cOaVw8xqCSm2OCnv3yyOC74viwYC7Okn4z3s0dfHpaj/aKeZY3hOHopPkFEiTe
x6VkXnVI8fZ4zF9eCbklBWoO6v/w9oUyKB+0OF+aVmj1cc9YmFwATvyQK51IWaJF
lfmqLpY+OnNaF6QY5CDQhC1HHjXexR9Pw8EYRWI4ilt6asebBXh5evM5w+hyAhgS
khHrCvYUOPBrK7lAEjUNReSdJY6QqWYxu6oFWUdIismxcUoVAQQ4VImg3iUIql+j
T2LqAGyKihQ0wmMM7JSTdsOzl0pO8TPEAngKG1d7RvvqHPuC9su4Q9p9efVl85OH
fw377yAmjS+a7Ikl+NFvFRTAC3u5Of2Gsit50aQXILmynoDWpVQ7mH63+ijm1nT5
y4WvTa43i2pVFUKl0+2UAMx3S3ltdnzqBhbP9VrG3ZePkBSmdfxokuuHQpDGjvwP
zyiu4WxSjY8NzD606D51rH9aTPEJiBwL8tlRfNUBDN+FpdBis71CxrQf6MRKnphR
DNAKgE4blKBHsyVdMTZpBKASA1aIEvNXVBFlb0/KFO0c1PWXm2rcUdCUJZ6YiuUS
VAQGq+al806WnGKJInHhBKAMMeb0zu1HaTnMxWIYbxkdNzRC3G+7mAIsaBVwZehw
kdyfMm6gqj/qGcEjMim0vVAUERYsGitaxaQoE1i0DQmxnir4exK5vyuz+z4HBP3v
8UvykwWAjJdDXtby0F/jymG4JA8LtVFNYI4WBhXDnecvJuySlkEE2yZ0bRkQtQKo
FF3kh8g/ypmHu1E4UxdhF9KEcgYu+A3Cl92oSBmy/gXhvf09Y7xXSL7DTQP98clM
Ga5r3QD5TF/7Lsjct7eHYVycKVedXdoKykk+WEwaskhfUPx3RDog/wL4hIcjcufQ
/yJrP2MHuhiEvAg99Zd2UVcp2v82dfRCdcQQmY83ae/guYrtW8Rojg2LMmsbfqB/
lTCPu1gntIs/StEC9RI+N4vfC7xmFBUwH4mRDYBA47VOQhUHq09ljK28ezpVDVZT
C+Dcg1QncAQX3JV8YfqcI4a7RI5KiM/aDphsEtdNMeUWv5i5Lm/D6cvKTY/Dbims
d123u9JWtsz1xogNsqK/nHYK0uidjJnwJSndMAXbpEUQTPQkxw6YWmZWCRjZj8kJ
WQxwM/iU+94aW5qWb3PTthH5nMA03VFAbcyFvWQPMaOrO8RGNV1g3ttGKM36eUJu
OhflAqGTlzpJ6tHxyL7CnG8TcWeFMpxCIf+A2wauYI0tF6J4G8a6Byfd6VPd0Kpo
65vvJMBqkciw2Pt30D/5RxMlWv1U9Jsx8Gqf2dyRjf4bnYy+Ut50VE7SITnzKooq
6QDo1x24yPJuZ4hhaUDI9MtWCiVxOw5sjs76DQPwPdMQ3u0tRCgmm0A8BOiumhL4
UdY5FiIojtEDh3uDBCmUFWhB0QMLvtkdYbLvP5P6tSVRe+V3Sn3A9zVpCLAypVhI
fQhzm88XmeeeyCbRcnyjtS2+zbbzh+Xd0RiA26JlFiZ1MMMc9hUCcrC9YmoHtac9
uqjVg85CW3XkNCSS5FAlAzXzCPvsO5dnouScQWsChJucMhm4DwZO35pzAhPUggLH
JGLGYvcHck7FGj96yvHuL1/tcB3JWzBMjiz61t+pqgizGsAdoHCB0iEGIDgk2N+a
/geyigpYqC4AHz+BzQC+DQDCa6SFYfb6kY/4oPdYGZHoJAhknyc2kh/CEirVP0ES
QZwztf9V0bxynpGCTGPjo7aiDI9Voc61ldgr18B+ZMfRnA+4Lm3YRSj4OQA1mdi2
+BQANJkR2r7ghWIz40KhbEPhX1BgH3ppkFxgZllWdNvNxUgisnVbL6iF9fBoZx6N
BeVx8eA3xYc0cWQsJ8StynRbxVBegvlL/9y57d1TMcJkoz9KqqT+Bpz2mMc5lad8
K94MoSyUYn5cU5yPzo73H9pY06edhSUWn49PdEkieh8h76yEt+4lAHjot0Af9TMp
MTSDipDThJRBVp5e2RwLxN87onF8FQLCozN/RI2IDuGuaF0dmFnZ+6H88L6B00x0
371a5WatTrBpSrma9mGmvTmZtC/InteMkJ9fU7mDousSBLwu7BBCgbPYJMgo3GEN
cGKdE/VEiWMCu6xfDXSPgEnDUawyH8FsoZN1tcDsQyv3YlyaIckatr6XIKQLrrPS
9PolR0rbJ4FgMArjR0bYG2uWiQgfQaPYMGRFrlug+V3oMzNuf1sho3Y3RVKV1XJx
slknQDzadiuqhYqg+l/DlzCmoF5RNfSzQg+LO6KHPA1xZVPFPc3/ljocJ77ZN7gz
SiyYDmwygl06EO+80L86tPW8J4dM36ICUFkl8pa53g1wYwbAO2AejG938sTDEK7i
CQiZSWMZJ+gSrfpjHmBMw3prlQHdDfOxyCDNTeHH+OH1J89NBOWKW9KQg/69Bj9Y
fVZZxUkp36mvArgQPm0c426JCoby8fx0LOFPWnJThdA9is99xVX8AmJuOK40Y/Qm
I7UWQWYldQPiLf1GZ3XlovlLIJpqAjPoQDRupm1woA7GHe8+PkdDsstwYog1vFiX
XX8uDFknZC5ZDh6dEQh0v4KwQg5kS/ohoL0xotGZ1BI1BLgstocTZToAACzL+Afz
PTFGSgj0RNsR3R4192saCMGCwkO6yOB07cOxY8wGhDIILJfc9eeWlCyn1YykS42z
BywiQ4q/TKp4ry55ZtHq8cEr2Y+GidBksVwb/8XJRqV36u9g/DTgDnbsKzTMnhlo
1yrk2q/sO4XJtfevByKoP9Ha0ROoe2+pPI6SymN1daxOCRtcN037hLT0xd8NC0ul
TufU001nYqC713lp6Q5VqcTCynjwoNozONO0BlefO6MYQJHESkqspM9aoFIy/vAs
PMurTk8zJCwC0DUyZVgJqrw8rfN24C5YW3OCsN1qXk/WAIkXWugadkSMlZO6cFZT
EVM/vAsS8Oy3j26w4Ufuz7cD52he39QifN7ObzcaXLY4CYEyxDCrMWTM0IigTXTG
xC6/B4DlYfiw3EfoBzpxOnQpLPPeT+PvDY/es7ubzeW36TFafzKZNnofEJ+jBokI
fcQ9FAKHV4Ox2PVWdFrc50i6MRFDMC1xdb+pGkM6I1n46CGklE9hFOfziE6/+tMA
7n6GXomR21qsfG7QaXDxP5gxQY2yqJqBQiKwWiCA0hJ32vtYT6ccU1FU6G5MpP+r
fTcNDj8L699gld84qBNMeuM8TgpM34ynL3HoTBgCZG6mMAq/Z3lsoJoXgN0ZjNFb
3mS3l8k21sbAfizAJN9d26XqKsvw0FBb/JuHMbwy53DjbtrWMpQAh9hzb+FbBdSF
jOOc9U1F6/U0yDE+N2X+Xg410WwHCpX9jS0+MKwuimylyd4u6h3nHQBtb3jMHxvS
G2Qgnh6Uw7mtorSo59zaMEmBlb/C7ivfWrmE1TxuYUoET8OBDONWE61reG1q5nvI
SY03sZ12Y12S4o1kAiP8chAw9hGV+OXgrhRQu3xH0fcJSCBAnGt4WeEoGkSC8DC8
OA0UuDGYRIrTAlGKvSuftbaBSt9WTVrKgsiNGGwiIFRgAnlOV1EtFDjI7KC6a1tW
C2HegWB9Kaznk+OttRknSsMux8uIY7vKSI18O+XnI/fqieB9utRmo5fyFg6AaBOf
rySQZCifDrhGhSKd1aPtMqmBZWzlTRQVehVEYU3PKrNik0h4LweD6dtpkQ02uYug
Spu+Mb5SGXranxAsI3WGnW7botYuAALPsxWMYtdPJt8TjVhRaOD0XVO0gfa96Elr
6J8Gmls9RK1wK/Vx9JcG6udsZyRamkEB4Yr2YfenrIyI4dvlJdGgyIYOT2BcVrgC
D9fqxhRjYzmpk40Mr+cLZBPhiTJzSL3cRxvm7g75dpS2zL7/djia//2QQb+THXl+
/AHA5KrSlfVCS1O7jHrMc0TDFI0gxULcewOAqqxvLRTiXwbAO4lv5pd2JkLm4z6D
TTfT8xd4YAQ4oNMSTHqmRaMYI76wNO7XDC2S7FsRAhpbuUoY3PmbXr8s/szZITcI
pA2FaGGiNq8tnAqPq0BSU0JfzAMCk0dAygyO/XV2Wqcbo5tbFg27cxURkr9NsyTB
px9itaRtjhRS+N0txYgOc3HfK6gkx6CAVWtTeY6DSbAJUX2K9pkJ7arEGCAqYGsm
zg+yOLB88nXr06/yEIbl41KP1kNAWv88h0eZwQ0HN5lFvJoMmnnNfvuJ0hZQ64L3
uW10D5MIABoWu7bEKzTFXY9bmGhEoIVXDq5Z/RczhajyCptDXKZ515BrSRGpmq05
CvHyfTlgD1QGnZFZr0R0xT2HW/vsoS/9x4dvkgOd4Po77SF6dV995cs3qlDe6cjA
srTd7MxBwaJC8hjq79csFLC5gnhcEXLg0ymQ3nzchhM6IpXOluMMyVAWuBKuPVxW
7db/7XRiZP63TH3/a+mh84DJSsVTUvkRJpXA1BzYSOOPN9PJJUkTe9DJjmTJz5+2
i15C3mb51dW+LC3+qsI0I+VzdoOsTqEhP3TDdHRGctOGpgNIQCPseWNG91xcM6io
z1g5mdlFQuZqqVhK/nEwmC+/apJ6uBhgbD/Mid4tGU9Hrkla2cxqcgATuehnywph
MyYwhuae+7zRMoQcnxaC0mf68FjXhxFkXziIXaj5930l5cpvlbl+bT3j2CIULebQ
SugzM3b1ck5TAYD+DYyVnPLEmaG6ZKnz6AdGRpVsHdW/sETZ3TC0cCPCgqtIJoXi
TPhefgXiLCn8a6y346d2eM5Xjc/01C2d5CWhWLgWnXX17hBYOMFfXapIgbqAOqIh
YkcW3q+38OGuZg1xzMxvH14iUQukpE/bc9gRieQ5OfitRtx3CDzdkDIf85f32hyh
KFCWzgUpRkIWma64Ltd8YI/vZzM0PruZSi9jA6zgKZHchUk7bnnNkppz5PsgtAHu
bCGP0+++Gh3EizdtKe2mTFdXUR6TICo+tdcMYvfKlX6lVXthRJWxbTFM8EGHfHEx
mpDoRfr+05NQij8OdY3LcO8sDLI50kdKy4phNUqYo6kRGcVPiC2a/RL+ox9cIqD/
R1qd+QoDRybLbz8ilj3CO+0uTxsOhTOePR+cFWmEL6qUICKuLjVcH6JXDdYLW+Rd
M896R1KiGRPiZbZBzPa+1LrNHDwk4kNbJhJDmt/oF18TBEynZr4rlKWX3Rbbq2I4
zEvZJTHi1IExeXe1NizWOcVND2REIpX36X0WoK5el8yz7EGm17OvQheXs0RAwkUU
uP4bmRrf++lhg0ryM4Lw0vZmDjI8UO57UJT35nwedU1Fjs1xRqMvRAWNFqHCb5wL
SVdAzk4XOsGFlP7Qa+FTDSe5RX8Yihcx5dZY0oZg15pHJ35/hWjbOb9cVXUF/unG
uqpCHQsDw3OctGYI3NqzPCnHQzppdqbVgcuFFIfCK78OHcsdN+yaCKLTGcwcP7sZ
fPjFc8JReTPV9uk+rbME2Wzwk+UnwjOa3y1aa4yuL2KyDQa2zq8bvl4ocbApj865
5kY3e4iBWrSwlyLQcbu5z8nSEhnho0th4bMNrW/zS9rE/PWXxpyvoG3r6KLxFL5w
JKp0MYDMxzR0Pbdj4CrYeK+4JyofNwSrWcop8OT2LsJjRwd212bujws874FZfO5+
KisdLG5c+cfUQTyz+RCiVJdySus911KMK4tMw/bLCqVCM+vHhqGWF8MWqmuefN0I
5IR1nRosdcdes8pu82Vxq6ScCGnCZGtwE5AAvctletUuwigASKOnUcXZJ/2qTgcF
7RZm07O90UPrzt4nCC7QEDCNV9jOKGbpk9ie35dHZ3vn8Df1yB/e4ws2dMdrz+hk
pR/zjjmxlJgDY87I9riowv4CGD+ZbPl2by2n2W4JxyeWvbQNXF+7FwVQPJjSRu+G
g3G1X/Q1HGYl0iV9WgIgHHam81PcJlKGAj+mZY8lRJ6t2bjUwqZyeqzF99kfzD5d
gCVvbDu14fWCDbHTzQVFOgIu8wiKRCAy2RK4/kNqpwAvU7o2XFo0I20KYX/OIi4u
XBcUbTDue17cHDkI4m8ljNFrQByLVnTVNxpKz1e6ptcsW0MDg5fQOgtCdRuQoaEL
rrVkCXU92x7SrIuVDk6hLs1ltCrtT6vUrPtifV4y2NLGNMxyQmannRjOw24nIFzS
kIBZ6/4b7pT2YN8WFPqoPc2XZiluGW+HZuhBnfQdn65rOoys363ZRVAId/gJl1aG
LjEZ0SEpU3JdjtE3dq4u5j6e/of/9W45kXSQzhXhD08OKoTK9mxyv9MDFejeu8P1
1lsW75kdoAFsB/HuCjmk7mGPkTfQ5OlJVEITreD+H0VgN3+1eBvz1ngI3fEgAWms
SuScDBbWhloPxqYwFj3fLasy6L11zop3UNGk0C2e1L9EQzshj8JMjQzPrz6+C7/I
sWn/VlZFUEI7uXNoeByrMDZzP3U68vMkYte0wAWNlQr4LHEuX1qgBOgr6TTGuldV
Ki2eBStOhljQxPqqXEk0DYpuyOaNA9WMJScfURNU5/bloLDZ/38BI6mpHJXtbA0y
764fsog1kd037I7/hQtbrASlEM/N7qGez4LlzgZXw/agq7SZoy/UVnMeTGtEfxvr
UYrTXrMxipUBRo5eA5Dq51QSX9V+y7OR9FTQp22o401qKSk2RYipW3/+e1OsfqTh
wY8HHHp9cIkDrHCNdlGe/38tw/RAwdmCTSnI0lu8ZuXNZLBveBnrmaYl48rHe4Kz
6dJBc0G/KbBsejPDsKiBDnmqCYL8yCmk99zUotJrdSjXC8Epx5m8Y11hkE01tqjr
Wv3eSQkwCkZrdHlVwerJGRd6wC5LYh3c9JPFC+5dRhlbdVuiVrD1DWekHQr9aZjZ
WJc7TEtRS+I3UsQhU8+Bav+eizC3bU5qzzNGOan2He9brvnzlmdukfAZ5tl2orm6
Ekh17BS/fUCd1ntteQk8ZBuuMBmqPfOghqs0C7X/dZEa3HRXPD5OfziuYCpxZzui
5JBBZPO4dcHDwpDtjk4jE2Ecs/J+Ndrwz/4DXi0kOOrHu6hrjrGuQSvvSRCj8nny
zVC3TSZfrwLYQhZlyZsyTSHxGwTBJmTQq6YQeUMDxiHYkf9xy/Qo2Rc7lpY7h5xx
kbCctj+fxAHVz6GuFVWrL1Gl+AMokeMivVJsfBcoyB9nF2CzcS+c8rI83by8/q54
1wHRgN5ntBIEwZqkD6gqldfzrat7LuJmwSjmOjntB2b+nd7BDYyiEMhgDruJ9DUu
y5Ipez085jWe05jU5lDnt4kS8ZERlQ4i1EG6IyHCt1wRKEjgv6ux1TvI9X9aXg8L
FsN1n8G6evKRp+Rig3rTpT1ZKc4hzA0PmHEGzqnu8rLIqONNjSrAXZDPcd/lcnK4
Cb+qZ2ykaIWjJC0eHt1uM5Ppl+KxslTNQp47jefRZlBr0Fp4HfZh/kROCcEcCqcE
+r7bgNTYHAhOOKB5gd1ggkUnwbuB/TSa9AWo8u6KbNZLFcV5WcLoKkxMAn04xP8D
1Z7UxbAFIMWidJZHQgXyjWCHPvYzTxpnOV74ThZ1N+KECZl63ooEOVX/HpV2V2kx
ajt4w+Z60voQKFq4g4kHiITrH/Uf2OA+8EKFhwp8vcLwUgjYZvTmGXjSsIsYy3uN
nqkcySMesfkULOmfL5usoZruh97qmfZroz4Mu4BE89Ovqw1SwAoAibSlAkx+ldWd
c1D3Z4ErtPrEHmeb9DrjVMdxhMr4QL36xYl1JorifGYQWFiSRSduLa7C0qUruKaO
xNIfw5O3/G00jDO3iF/Vs7CR44q9pjKey7Es6HbHQ7G7NWh65FlmNREVDhXwYpcD
YX9XQGZc/mwrz4WZQSfYibyRcL2I5ZKr6lM6hCEX9YM7r2XLY2g+Uc1cnGolCqPI
xl4mjwlcGPDsfJvhPJaPvnz4atPyvmhtFS4EJpBqinX7XHe0EvIQ1IfBY8RICGMr
x8lj7lTr67E2LFa+EPjw4xqr0pi4zyhkFYLezggHrmFyHsw0EEOCusZDLj86H/f7
XvqIowhqD5pOetilnMQ77bMDCpb3tuwAjNnyRIwsiTrS3xnDTB/ZGzWZGbFjNsmJ
PfG88NclIyqReevVgPFMErZabcQSATrVCpWwKD0TyLTZyntCRaS3TOwYvAAXk85d
ylX6LqV0oxpdW2G/atE+aPkjujK43+7hbuFQDuTKYHaxMlTUsVhdBZpxMjQSshZ7
dlwNCoLsFG3wfFVknEHfInDHdJOrf61WXtCYEyqgX+yHEbGWsvFw9xmU/adCMd32
wiH6h1xP2KBZ7kMw/FIIAv/ZjAIoZgLoAVkRfFgCayU6D14267rdor6/+ncRCyTE
lgsyjS56JuVGLoCFz3ArX7a4/nOkJm7H4pQJ1Srz5eXMUC5gH2MPRYI//NN+PGyn
3AXsBQuvQ+pZdLNtaJld0QcX4LYynSQaqXRWM6Pg6tfI3+Shtj6u+xvmznnodRIN
VQTU+BMDOKkEDLf5PDkLb1cieDA1lMk1A5aE8YwHWZ8UDEcNv3ElyspfsaBW3j5T
gt9484WbKbHquPZYeXk/WRPim2jL8oj4PSOHHnNRlZhUNRqwcf9v/3jnNcacNcQo
tqRczCW/ufW++6mG3JaBPJqBmiSW3+B9UgvVK4Loti+2JrRhfNvpARPN5lDXAWux
6RX4AfGzVVV622tBSsy6bKq5C5PvG370WAHCNC1x4X5MRLPzSV6+Tng9mNHfG/wY
fSioetPAyTIvnrGVH/A2uch3S48DjM5rG6LAE7v4Oul9uUJ6DwL5FHPaQjkBteLn
4r4sL4/+0XZqAkkzq5mLxbBclnp7eylSV1qdc7WC5ZMsmj3n3OXwhtJ2OgFsaerU
HUFf1QSz9qm+7RBEeu6WLEGbuPHyhPOurz4Q6uRn9lk9sTAgGRsfjNSVVZp3UGz3
/wW5RQXI3t/lUaQGuiPEk0tC6P2VwgtSCnSYwobzKUe0F6ZGd9aDZmoT1YZ+aObS
aoRGSwhLVfxXXR/vgA4542bob1KyoTX9I0NJ4nwv37SaB/hoUoQexkzt+Lso8nUK
6D0WT/HERpM9SZqFAobbyZJXd8RSuFPJZK0lPeVj+WYzo/PuUaiQY3exU/z62mze
IXb1okNIrXFn9dtMRMqgGw4W6IsPeruR67cmmevjJNg3cc5giNqnjgJBaCl4ofUg
Ia9s80qiDQR6qdDpYXqeL9o5oFlzh9uAak5toVK3Cqh+BpomhhQp14Mokk9IJbbv
4mOERm64fzH8CHBDRrtYVtaz1L+Nkp7vxZg1EpG4Bjva70tAUbSZ2Tmz1Oa2X4yp
jRnoxrkJ5LnrJjBFm3cHInm9sR1HNSciLoN1eyO8Yc7QvjvbXPPwbW1tGB/7Zf42
BgvnGRpNHrymjVFvB6yctpZYnuI2I5vzO9MjoVv6Jxk/XY7QwU0SXypZGDtkx21N
faQMMkJfRdeMmw/7heiZKDUpDcTQQ/FX72wVqn83lW2wsnt2/DLxvYBhN/XkbbrT
+cgNSyltIxzV4v1UeuPwGA/3K//9CdHUToy0gbQJPn5KCV4yUOvYbSu7YNShiB21
fzcez3qZAGmIPVtMmv9g2TnRO+Kdo/usBFl/YnekjM5Wq+3R807xFBfmxPVNnkYf
9jPcCCh2Nf+mZvek6j64yxiYHanwlhRyDw2bOgoOnaNfrLxiUAthOr6gLaCaNhl7
NgxDiLJwdImPsd4cttvQ23XPJGyVdffuo2CFWrd+kCZoeSYND2cvW06YLq6GUJDf
kEEh0iwPU/QD+zLvaC5oh2PArdvUfZ4Zuc29NNyEePHbrpXtTBoPCJzEFNa4bYmB
KqJ0R5MLCJQneWtb1cI6L1HNLrqusB2jtJAunx9jA0bojWL8woQj5JUWxiVo3YIO
dob2EjaCDfnH1TvSqUlOAnoCszhfojMjP2eewr6KRicRoDTl9/uajEwzED35Y1ep
2LScMgXUj0xmkL39AmTPfhtn9A3cJVSujQ6JOxBE3s36RlMA3DLQ9ArSO6B94qBg
safa5e3rSg9UVjXufu6KLPbEwTgPB4CJ02EchwzyW2Rgd/6VUWg8Q9V4h/HlEQ8q
Q2WVwfMwrboHPUKYjUgUHiKY3dh8UG5AppBGfODbvYkw2eQk/mIZM0N7zPgGQ3hw
RAGaH4rBew+5fscP0B0MT09CvPojBRgaOeABSb8yzrBDfR01kNnrPFqEHLcbrmm8
oG8lbP8Gyh79iBKo/XDnuVo3pf3SwUxXejG3yq15M60/NetXX+JWVrqA72zD+7ig
Bg5ZgwH9UMDxxB2CASapoogtPFivI0L8eDhGqHNQXoukOglAEbbWypQPOwaCFwyv
MRo5UGUqRuL6I5ppMC4sn14n21bAFTGnkYzBo1v12gHcup9zKzhKPlSQlboleXnn
EM9B8Jh4glddBqqVef2iYZfarKjE62NWVGc+0tOIvlQWdZkgXgVZij3tlsPwWIdc
ZSW/XKxs+MCyA2goJVbeI2wen596z2dfDva59qQOEWUAc4SB19rMzdMzgbf7gwQd
oSpZiwmHvQ54bjK1G6hIzBhyfrTxxF+9gJ7H0jRUppiDifYdY6n1mYNO967QJU6D
58EjLE2m0MJT9LH46tlPS7KWAn72Mhv9eU/Ql0W8/1Iy6en3Ep/iM51WEOoyRVmr
GIvvWCJpuIncRTCrJdxUUuC0pbD5EeLrlMR4Ggo3dOhoUzLMoItju1l/DihPQ7Ug
JmeQXYlSzqEUD5cEYAxK8rcuny/y38lPtCN2mkdkjfXQL3r5I9Tg3Zhjlg1AVmxN
uzVLby2BDjVUGP/siBfd2zfFlrSM+VH3fDZH295hqon2ZoRzb/NstoewgDeFK/6S
2T6UjmO+OUtDn9Uz8R8VRXs2hwGRpfGC6MsiUpJnFavB1ZRGqt2Oo5N39c0eb1Ts
4ue72a9B1FIYs33MHDmmRzlL+wJDuprmCe+p9qBGm0oQ+MgOJKM/nGxKQQtm//ia
r3HxO6rS9vo7gCa8ffQbpO++vyQnxCjJsThjQi9ilTjS+pV4Z51AfJt+KRWLWLV8
QUGkf4xNmUxDgF9Qm6Thg+JMnf+vvWGZttuUpweGqGu4Td7Rp0aLvqA4+xnWbinH
0blxcecp8vFa4xBJ1YkUJLtun6beLA6S+lInHVjTb2OFDvRLzJOXVIF9rnOeiMh1
vip0UgIBC0GPzinsayXvQWj59c0hwV5mteUmeZsj8u9xDVt2B2gIgKDFFG8l8V+V
qsb/e94DoprQLwK53tVDMD/OMepwiQCWEEZNxWUbkY5636kV8qIXr+BxaI+vkkq1
qcnUmeILcovqpgfkz/pashlVGqK5yR5Nas8gPXWmW0OwSrhFun0dM5ICj969tIOC
xBHk+Pw8igfmca5jx2HGMjxhsElvL6gMvg1K/0IO4aQJLcawkWjSt2WHb/z8oQfx
r1CsbqfzvA567UUOmeb+jTLg2Yt3B3dMjTRd3dkkDs9peWlW91qqpGWF6ei4cOs3
NuUjF3n/qDyBW3vZmm4oBJ4JII0+0UtXgF4ITULMQhOlENMp0+nvgITrltlbXj3I
L/aAg51gK+4F6IMTEUEZNjBt7/OcUHJe4avGlFcQXoicHr0ZEWImIX/ZRfGoSmVQ
AQsGm8jwMkOP4OW5ev28E2LkHThv6ipl5F+rKLyEn7A62C7pgoIZIAIjB+c1f71c
ubZb79E/5ixyhG343QvLC4jchgwwSqm8MklGbPPixYJhLxJ/9FOW31daMH2qdW3A
sDn2jRGpiMYW+ZTSodnRSjz3r29V97pQRK5CLX530nfo2tfbEoe1pr4f2XLQOta1
fgTT+0B+kam24dJGWteBMvhLQqcx8K85qC70lAGZ/8VyuHAKpbpB0VuaXHLbAMKT
RvXIATBXA/nz4F4tBPd1sTQoHlY7Nbl29PHByXS7OdgzuZHStZxGgj+L9OEBfT2e
htaR+kR7QKOKlsxS9AvZJ5ZIVMV+T4GjPvoCXi8do9aQdTUYk6AUjx7Iim0gKUda
MqXesli3+QcQGUHwsoqktPbDRGYYmkPRvIrxMaHGK/df2rhO0TxbQJjWuCa2n1U2
ADRx5fjOvQcO49iolGvq2iqQcw7sdpMjHulJ3RaypSrxd1McnL7zvcz4E2z1oYq+
R/wRUEz9qKp4M8tXoYrodqfPLjWff1xYvmHHTAtQNYPucNdA7N3ATFri5PxiBxS2
lVyePAIgpDqFLsg/lS2XTTg3/SjflHrpE8WPjFFfNrAKdzKKctOGlkQpGXev4Hk3
/t2XCvHeD3lkY9gxo2cpH4t4cFnxnKRpnoEUiC1BkwDb/cbSZDtTevEKOLVCburl
uk3VUwbQzBfIz9Aqqji4hjNlcS7dlyd19vx3oLLjHAijNaRMWEX9zlg7txDRQOnH
l4RQAU8jPFi3kfdG8VpsDAG3GBHUcoXbvC4d73OXrotZPHO0ruHy7Wc98uTNB6XA
7AnTAZ6ggceDfOaGOivCEYGQok+Fa+erqDIg/GuynWEJlGsKlaWWPZXRfByipzYp
F9VNMgKxFAXKT6hI9z1tXfZhcLGxoSo51Lb6VtdET5vPGWIYm6v9TJku/p9Ff7/X
RKL+oBrkxL6x8qVcv4xbpxMJEFD0nhw9mJ3ZgmpXHs/NPlp4sl9RTYOZOW42nQLf
97tnhyCVPKpOkuWsXDySLFb/quehgiuHo/m4fI3XbImfZkxEV8iYQ1bMu89EXoI+
/wPGLr6gxqS1V8MrEWjNYxK7MnywvRJ0Rimd4QuxH0x42dCn11mRBAzGOvYkx+4q
GPetmdsW/zjTO3ZMYzWL1JEZG3QcpWnetPJ/HmQwmgCK8ZuQXm/p63bJ0ADEb9WQ
/VWrES5tBBzDqwEetBgdXjycFKAw+Hg+k2JyU6SPQGVJfNmNeN7H6I5oeDvAOArA
1vHulzCwV+RppT0P5iv4S5CrNOUcf2LDEjiyNzHqJxnulZIn0EwOJC9FWWy5cq6A
+ZjFvXI3YVVb6FqO8Mwf2gcXDLuRZ+NP2zYHyy3VK9csS0oDa/lBsYuXOR+ov8AJ
l4OkIm7X936uNoJLkioL881r5R6j3c3FsYdM9DnhzpnJ07dXeIiV8VuD0upO09xA
TNt5/OFi3VrWWH3nl56J+cj7n/I3Nqu1l6VyRTavlaS51UKzNanr5bJyPKuNA2Ow
7itkq90BJ4CyR0BKAgBQ9mCdNV3sr+jMFy2ilxmz2iJhbiqOrS9CCTb7puSMp9Ll
9GIvI0kPDCTeaiVkLkBQ5vfgeKhxlWXoSDgJzNT1wyegWY2FBtEj3hzCD15v20gE
n/vYiVXGIWTeLzOp9zeGuVc7+N8NmORHlprDTPFZJnZPip8+zJ3smECZ4qeUMNm3
eWnnUARluyR1nfP0xq5usBqj7qQfbGSZCNylhwavnTSjG9fRi7/aqGLA/BUMtxvg
xyoeTEdYdlmHrk9v1RxdCoMRw6lyn9RGuB7NkLiUuq2c9/XaFXMGt3Mq7XAjpK7g
U3fzbjy9iO1LJIfF9m8RjsaXANYDoS7SzQwTLwEgQjEV/8C5OLBDBTh0lkCcs0+9
WiC11bl+mpWBBRcqNY616AM5hSVcxos9McnwINHv+1yKhdCUocJnQihmDIMNMSQu
jFQ2YfrqjX+OedDBBY1ODb63xmsmYJ1994TTwGWmpI1F6FhLeFl7j7aF//pydGQq
n2zSeEfslj1IVIDdUWaOZwtTOnrLSAWqRWFUWsAxRbEMsnlGeVNT2ltDisEE+D3d
o0+1giRCJqJjUj19Yl2T/jzG+wAM2AM2AMkst92oMEA6gbZSXiEF3XxPPkuWLg0A
6cmIqb9QuSOjG0IVALMDUyU0OenK7nzngAYcx9c/sB0mPK2eIV5OeHf67clre4Z4
+gYRg0NLr4pO/vHKYFgzzBwhjAH9C3SFU7t1kiMa8zqe8Rtz/hiweWam5zqY+cFB
ZowPTF4vOVdA4W8rKNDi9DlbfuqM3cQHCb9RoUKm6TN0X2k0TjX7Jl4nW/9FRlt8
yVRPK5kUGM/0of3R7pRbvzK1Rh3Fg2QOWQksNctRuUo43q+bCmCzQfXzVG5O748z
sDwwBSWAHWOB2qhCx+eWpVKjmt60opxVXLeOA0Mtr51L0iB9SaJWnuz0tXrMnJLC
w+3VE3yO6R3S7hzJRBgVvTWoEy1WUP5vUFWGmFqROacr0hKJBKWcezCb8AqrepRQ
EBGkZFLbCIAZ7yEeHoZ1+qH5UYRmoUBPoOc0Q4kvKRjTNVzFcmruyg5eNYM1toHA
kVJizh6UnMwi3yxX5fJ4V1TdyWvKoYzQxQBSgUtpNY6FcSzf8G2a5IHRkLvHeyAe
A0QF5cqgYJdbwj+0duShdW+rxqhJuC1waJ4UEh4Cf1DptT1fAvEONNeLTWJxLvQ+
nH2t3dEYfBJKz66Mf7OElQhco8c3/44NtV8VW3ZhOCYz0gBR/DXvHzwQuD0Ty+k8
xt1Fq3FD0RLc0qFiV3OI1XY9g4ZLeCJHYsjJk8HfU5ULZWyJSCktcRTSr0PW1pH9
Z6DERNPxw2cRYgq29vmByZLwvS2wtXAKG7H+qT/gBxu6hzPAMfvMzyj7HJQdMgr8
F+mP52fEeiowoM1/Xf0cEQDuV0wBQyk5Ju7aSz3e+HQY6Bj3tqQoHVj4poJ/axUm
s2tSFs2YEybrp2yhRK5HIxa2xx5AmPfka0jfBQozEMc96Mabcf0Tmex19tQGy0+3
luMjye21xNxBd7LdPKsNLZe2HFXzyBdR76hMx6+oZr2imndwJaDfcHYBFeBwEObR
rF8gFT4zo4KEiECAa/J2dxWPVrh/y6hajirbijFa+qCMaqt2Juzk35wD6/gOAVYH
p6SA9piLqLjJ3Rf1jCHfXnM56DYkvo9KTbITmTTq66sw2U8z24qkQLuuuN1k7sZr
oYSUx8Ic5RyqeVxkr5jfT8V/Ck8SwEeeQfYAZC/IJnOz/0jKkrPEPnHJFcGD0c6q
u5ni9TX9SVm4LcJ8YUuHZCH0KuIiNr3+ejhDWq/ktt2ZXQk6J4d0zmyFGoIO052C
t99Tk3uwI7aE6ttjBFeYHy5WxbL0XiQy6aHxylN5Q0Ev+Ax0XfjGbIKALzisvk+r
OQe0JukaCQk5j1YklteMLbIzR2SnXsWJ1h+GEoRqrljie6tbs731ceBnqRXUAFbT
epYlUQuwBLI+KQuu1CUu4ur+o5/k/UW5Tcy5N9bJQK6HEgP9EcN5AkPV02tTHsxe
Tb2wuicsdCJkZrPWec+oxp4TBAft6VyOMV1ce88Olmk5YFFNkfyuw0Hi9gcZc5xT
2tp6MW57A436FvBqEscOxomGgyDBJHt6O/zdfFbL7o94zopgoNdxJJdyoKLFvAWh
5zkcBJUmGzpezha/TJwolesRDvSag7+qGIADjapyaMjN2TH5fEu9QN/cbK1TrjZC
FUpRIXihJfDPvMGUOJ38omND5tSkGEKjWBWTfJj3/MV/8wxvQaIC5e0ggD/FTFzu
sliKoGnVKytSVmkQ6uPZdzC/J9VhPkawKBd2oIgQAXkh82lpd/yDBiwk7Z+Nc0bD
i3hlCMfz5z+L01yjalZGKwqPo5RapgQnnboA+1ljMx6b9q/LtshmtHGkrP7cNA7i
PF1wrVZNnSW1uzrasBccsV+wbEQ5dBF1RMzodxVVo2rvwuovg281N0EGWRyBFQNp
weR9nnoIu/Rqhfk5wHozhcZ+Ca3n09Josd564/xlzsr9o1IyaLuiL+U3olCBss/8
e1NJmC+qLA6bmqblPK0GSjuFjZzl8BUqmgAf5tIeuVzQ614bIMvPvUYZsCfJuQve
q7KybEO6A2+SHz+kv+4AeiL/U08PFYTbSwvXUcD2rCgwoe1PWLo76OO3KPCzB+mS
x+9eZckf8Y4EZYuiakbqN4mjWb6sAowjBZK74Y42MOCqmWnJ9rpBmKaTS/wt/kn7
3YyzKbkiylufdzAYg4RsYLXu98Vf9mWgXPAEjmRXOdV/ut/b90kdx2mc3k76AdHC
tQRN5qsQZOdUEUqp7B+B6PT9I0nhyUOz75Kn6a7XN1Q2HyGxcj2JdSv5gH9seJpo
ueJiZKkEkONraYNTaNs75xGMf5Mx83bKoWBsle32Bf7pz1aBlboKZxEKID5CC3j5
kWIc0KFyeMmxmHVw1PncbQHp4/IRjbuQ0LD+FZKhIE4yzJK1xxA1yuZX2g5Emguf
C1K5H+2UkfleiC7M2NvQdoW0O2nJLe0OvNdPAwHzOHWizJHcsYD/V0dbLrliWR6l
cdtHXFXeSVoZIdlDyp4deuCYz3jvpbkr8Bz3dVkuayAAmpf0mQhLaqTiS0VfRBzB
lLYpeIiup4DkMjT4ALAjAFZgq7U2qKDbSItL3m5DHdojbQlGAi9pACApgDw2RMXt
HclV9gWJqnTMuvxErD1M3XS+tsM2QQywyMOcpRxSBfGg2NTZpEkaKbGLgq2IrhKs
GBN4s1Mekmmv4pjRnT4hC+UeZWhWnSUIxJU+u1rBTZmvo4ZKNhRx+KIBC8H9HtvK
Zm5yUpQ7rrkVj8F2RmGDPF9CvwPnenEhGGdsdsQndTcSavsfWmEMEAuWSFqurob4
j2xP99PI8Kz5r1L7xQQb+3qdhjsyGCjZPdKiL9uWKHF3EgO9pN0Jbtkv0zqrreqL
nzcBrvRzwZ+cSN/lGEbZxQBlKEqnGa4JWqSrnbQBa/JMWpylU0FA/j0CTEKhQBPI
9m99EFYKveo+4zxPkrsBMJ1UiIVHHVxabHD2PvDspsUNXNtErjrViv8XK3Z51KnV
wW2RSgvcG8dl2uFYgqmrZSU3A67nTHMq+Z69MsLZtIY45UZVJAl/4wgvEw/EAoyz
yor2vGmPIaN+wzZunzoN/7EznvOuTcumWbOC/P197IJZ3pGcDyPXe9VCfcKpLNaR
aCJVGyTCmVKuL3SvR3ylqFKAdeepEUzfvDFsBcJkYKMtTnj3jflDbEBvSKZzhEnR
rSdoK3G+t5s7AXXK2tE7olyb7MAagyoypAS4QELnMZbtDHxSEoan45rw4li9FrfL
aINxQFtqvFNCc6rmg5dy0ip0aK052woWGPwIyfcNX3+mI04wfZSLN29kyJrAL2rN
67va0WU7jJ+ArYP0Rqy+hxif9m/cR/sH9dZXW0SeBqDX7QSharduJsvmt0lHH0DE
jOnDcmnt45rRB/auUOOVrLenWP2nAj2XxnivJn0uyGDBgrFpyAgk303t0rA8NKu3
BBkeUEZaI/gBDlDunZkndy0auzHMINkQiQCronGeqHpudLeYVKTNG/0uHq/qLPr1
RkzsujVc/bgoJYhHJnxhI1M03dw/apPN2Y/a5jTZ/ZD/RILV9st30124QlEHhLSM
lOc5NC3KJOfIMjtXB29CIqlVLgUG73ijw3NJRXWHOOz6KUkS85lkijTb/6LDQxeW
yBRSnkIMiwWsq4sa2vJrvxkAN5GVRPdZkwQcJ7OQpLIYOJoS4UZHJemRTB8+txVF
8wM8yUkJSGxwq7MgSCIG6YYX9r0nPQXG+XtLBBxAv0Ko/drNQE/Ec6gPFPA3SePV
UjrPthBa7muduKsRCqlACzmr5zXbd8KBx/XNqSwXQjFplRLkBngczccb3EcUEVqX
SBb6cz61chlDv5fD7se8V45auKcoD7Q+Xky4lgqO0znII9qK5R/Htmy8EmmAqypX
FnL6Z5TcZhUmHDDbYbg2bqTdf/bnZqcdpzLYeIv6ulreLH+1AytjOKpEjm96uxwF
QYbFxBdh9ELQD+0ScRRyuPefp1AC+s6iCYJ27bulEHFc/UQvx1DGuxy4fCDMCK+H
pRQRbVLj3FUioubobjOl/SQpp1/cqjhuQUdt8pxsyyajQzBVVOS+fowpM2lQqNX4
mKcnrJS5p80KfK+mlzjZpzFfUBmNzWYydMGtKAPZqOhE8cnrX7gvKm3xsZLHHqT5
lFbgkxQdZIa5fwQgCkUKWL6Mngtnf3eiep8MebmTALT/SO8M/kcHw5HWC2K9fDWf
t9JzWuAptKBAjehdLk/4iY9hXumpC5AZKVY4a6nvop3D3QFxnb1ZkvTTKTf0vw4V
VSawBwO+OQc7V2BDBEgjpX0/cGyrhhu1T3Fl9Pz6IVIOg9h5N4FwJw7WVstqKB3n
ef0W7TynMDTvukP9iB2HVt2d/CB0w6seTal5rbcmaBtfAuwp+viXC6qhhB2Ev03D
sSsC6WIPqbT+d6jOIw5ecuHUf7mQZRX+DYL+a4mlImPe6HJguI4RYB9B+lzI/9WO
gEHzY0vH9nbUPLWb9f02zm13Dh0CupVCTVu6uiRMIaFwswisxn2mj4nDugFdhYua
TWV+8f+ixbkjlVtpQyMMP7RTIHi4LGm5BecIyVDc/AFc+Dl3V/kCunqNtGOzucLF
0PlvD6bFTCtbJfn50zZ1jbURBy7iG0JJqjjjGr0JY9AiE4gdx9aqmLkGFlb9Y0kX
oQlnBG0ZOaWKfNmzc4i7EAhdkoJSGnyMRMTBNWyafDBlYoamlcy9I6lgb86dBw9H
Wx1jZoaM6t9sqGl6zKpxy+5dj/hvRX9MgM9vHnPkCyEl2YsfcuRJbL+xjgWCSeec
R/xBwBoJcQMG949h/N84cSdin/hEwqqEf8WWl3XiWOaFx2kpU5j122InEz+QrOS8
j+PoMYC5V4UK+GPqoukxEQPnE63aL6z9Uf4TeEj84bFe4BVp2R92V2OY18Ox6150
m7QJvNh+q2XaSve/m644nzPzcq5LhqL89PoiLUgbWSUcHITD6NfrRPPHKhtK9q2R
9rKBvf1nxn+WDrGLvucIIKCxCMZeP4wz8G9F09ZlWDYLaEqjLZqyRtTYoyOKW3IG
2TgC04vaOh3avtmj5iZ3kfSes/L0j+oo6IGzEqikSq5y5uD8k0O705UJd1Uv8jW7
2Fx2rDAS5Jv9LCkjnekZKcJLaC7V2kWKu7RDAOdbzV6aB+iqriLLG5Onmku1rQMg
pLIhWW4Q/wCqOJR/JLj89/9pQOOOuhg3uzc4eE6iMevj1E/wIBvJAibkcb9KN5yF
N6o18Xz8jndRYM8F0LGfKbb9RcRbkGQ4MdyMZ5OSIZViQweaxmopsTBNJ2RFbVs3
CHlRSoOv8O2TU+ffG/0AyKagmB2CBhbNRQQ5lr1jexHAuODFAKuR8bsdnjPgFCuZ
s+JI9kg4ALoYPA0zxNzFqKJ+Cq17lBbjt/BLcVP970Ne9icN0xpafW02QBJD5kvY
Ofp93XGMEQjreNlPHrwX0g33E/Bdckytgc7HhTNeuarX3axTSu2lFkf23o3Z9xPF
zQLuWecY4VyO0hr+gRcPWJPYS2h6HrsjYrcBJZ5SGJjzcJLafnJzyEJn+D+eiVuS
CWJqk9jNO0ttkXNs00qzwxXZHdul/063J2yYt6yxNScJzfpKtyYElFwG07iVs4YM
3RE/DJqOw9YXvTH482GcgmQmKL89bZF+w9UYJGc9WDx2l+HtCQgHQRsNDC5KSakG
sUyZ0hdzPsYEVwv7FO76tRLnWGspwseUGhBugKiFFg7J+zFIQP0MM6+G4t/lHX7F
NgznHgNHCNGuOPXaOvTen6+jTiYRmPzu07Wn9/cwcoZsHuTs9fywDiCKV2LifJ2u
7MgT1e8RWKp9WdAg4U7KUfzm61wSYketf9FlHWXxA9lTsYRgTt4yVYtlzZdKMaXm
H4fmmRYL8AM3M2A/qoFus8J4dMfiRbETNFObOmBFK15fgUOntpQLq0eE31xgpCYq
pf0rg3HzeoRph/WvocHoH6SisqV8f77GZQAQ2kLTXqFgvNvg9kYjgdqfRD4yDuet
hb9kIDzdtzuD27JUj1Khnzs2kZ7tQKhZ48uX3yROyNIKfwVecvj89V/POU43qcNT
YWbQsQBiV5xc/AWjh3iHIiZePMRVZeGRaRiVbdQbW/8B6wDqWRrSN/UAUIQ+sejp
CUjN0NqyjfnsanLDk7Oabmj/D0JhCoGZV3CiQ3r22yFfHzTWateqLlu1GaBRdoG2
ZDvIe050jua+IXonV5dn2k3rpMNZm0dyDuek3h9Z4XxnxcbVbQmMvGEUBzPzCxBy
+7cwA1qfGcjZa5XEBAuTYIl2NfvnYiW5bVpkPYsRWApHntRluxXUGjX30qd3DKTI
mSu4lUT2G2ZdEIEBpPbYoPL0kmEml/XJ1iuCCo+k2WX5yrQae0KRwkWKr5GDM9hK
LbOqBm7EDnXfaXBhLeVLWxA0OuZkx7TXnZiAf5d2wl7861Jtl0so1klScOp/3FsK
dK7YhTB60eP3HONnYQbSkheSwVpRJFm10IUkwaUpY7USqZBwRmjBOgcx42LkuEuN
xvTTWlGsHcMZ+N+97VUOZR/bWBK1AEDRlYgFVHmBRnVTc1eYfQ8Q/kTZQYeBZoeI
UabcpZ+kITThaggC6n9IetZ0YmgZ27HBoQwx8mCnoaBdoP5ECOGfaQv3NRP1Qxh3
yNiSnpRooMhj8KIdvHFkhDt4CiACqacDvvK0CVKHtFA6BnooRiZ81Z6A6UBYhEg9
aHRbDQFFfvUK6TZDrJHDzkUKRWYyoKYtXDxFC/q8KuBBXzBT98IRtJelyq1WEOXR
CxyAXYeX9hOtkQVoiBRR/3E4PKTcEb6L201VnPah78XhLE4KEtOL6Zffg060qetn
ZmV2PB+3AeHOWUe3cwHIL27ekb9FAt+3B/i1Iqqvy2mWvRf1NZPZDKsDw9eZrSQU
afR0TLisvmn6fCCLhBFHj8D7B8qrX7o1SmChzTyFcOOYUrUuV6eQ+VltAHWIhetf
WlBxjMHg6fCs4QRe/GLeqnH6SIZTNX/f8GvetqXvzpMVjgnXVcR4DAyQeemQl3+0
ZDHEgj0IKWhieXK1OEAOnWz6l20qZVaZ8MQWhEoxqrQBhm3XPjdVOFqRczjG88L2
VhHe8iVHSA3gvF0jfYkduwj9Xt7nusgsVORGbtrRZU7ujWQPG5LjsL10EFXr/7RL
FEjqvARN4Eu/bDQOB86TsRPzuMWgH/hqjWxjBHVlEpQIClPwWkfWjB8KDxTEUptA
ROl80cTYVl+/o8o+gO4XV1DAesVS4xCyUUsbwXOHi2bNVdUv/CwsCVJgcqpFkJOk
FkrD3yL5TIG41SJfXLiijhr+jWtNZjZoGMqkibmhgjzoBy+H6jYOW31NGZlHrzPw
cgbq9mROyzGHAoCOTrp9ApcjXUeh/cXCkKkDudjDYA1SPuAMT+fh3SEP7lfm0uvW
nj7s2GafGviLsSrIgSh9Gm4EJAQ+Pv3tGsJ7kJwOh8VVX5yNRFk0TTP5FytFHCjA
HrhqzWyQycKVNKeyS3NHdTZb5S+CPdGccP/KNl0NMAU7Oh53XKnvNyU0aqArE2Rd
EVZEV2aF8PrvTgworYXe2EDn/r6r6TuK7YwD0AlCOhcVYx8uP1/OPP+/5Z+n204f
LQr4w5Z4CMhn4YGc+TJ4FGnsPjuXbGui5fmN+sSpBpuOJAKjsb0Zw7RNLSTyR6oH
wYnQLuL17iTtx4q4Yiz+5R7alG1k0DdBpSEbmBUOy4tuE7OYRF6tgQ5tbQpIKncV
9Rf6nk8LEp9T5lfdYrCNd9Aidp9P5aDO57w/Y1Vu+LJrS1OV2kUEyzTXEY3DpDWM
GAFczfyfAN/Q2xbQ3TaTTmx4+rJQ0LWcd7nbrbvCQGKhe7P1393VEvNFc2s9YHoq
c8KpwB1yrG2R0sG8UardtCQtrcX/p0dWklSpxC8OOZzOZLLU/celZY10Sb5AaHYX
bok/U7c2P6TMHZSd9aNr65bORsxf18/bIG8q6LtKAg+3tPoO2dudedAQfKyQrLgQ
M2ppskEQ3ZMltO44Pj/vkkxEVhjHYaKx+cA/7zQiFVqHA4jHYerheYb4rS6LqEgL
1yFJu1YyVAuxZF+8ex0MOqsekg+8y4YhPXvBBBoDiLSXZ8d8OUFg993ElNNG/MBC
m+xt+CsFN4O5MSu5ImAKLeWyv3XPrSPNWYqWjYuYnCso6JVBFINGEPEX96oJA8Cf
yjfkQGx/iiKoRMviP3Qa2KS4TIaYKV53qrqGfMmayQp1TqQ+/uGxCsbhWydfJ0Kt
qe9ec51OpwLvM74iYtfZrcoUYjK1l/o4BqGVYopo8Ax2jk4uVvCyIWac6+KHCHrb
bMkcKTI6UOSgsdjswieaH9WEIoqyfSQSFOFIG99MbNprGKR0tFQHP09x2WRAtM1v
qWrN3tR7VEkgBFx3v5+rd6/MeFISwyeVKhKsgjiiy8brxsV64LpOVV5T0VZrSnVc
ZtLkzaNbUoOdqIHh3yZGsF6oFTdoPXyFxvVTAGlBmzPwKB9eAO08e/aPgrawsLlP
VxhwJJlZNBFJnq6MpL4W7jwrFp3kmZuSXbRqn7UvxHEBTw02loBeFnETcyLFinmv
GP/SR/DBYTwk/aaLUuEnhc3sc3PDk2/DeK1QPStfCsq9rOHqPNE79/p9Vl6pAzVZ
xHPvcsSYx6KfANDpmBkdzVaTBHFUX/LG3U+cgJZz1hTOe3cXw9yZ7Ik8yaIRVW4a
q9P+3cCvuD+bqiZYL30GrMOsbM5mMdv0EQilwxtWjNF2eNjskf2y7mKcMTjkAnpM
EyX0QauGn20PdCjxIoJhWpXCeLnWhSX5/AcUW+x6Q2PjYunniuuqtBH0PQGbDpdK
AO0EiGYgVWQkFmtON+k7pdEdt7nZrV7o11tf+CdkvRYJRg9t8k7WreSmUzitt+1O
2JRJxt1YU/uIyVSvyM5Tucocuw1EtHO1z44ITHKKVT44KXOmNRRjZX/O5AtsnCFm
14FwchdgDsvDe1aCd966qdxuQWg0eco7z/OZI2POaXtYfLfTrqAthbbSlJVMe+oS
fgkRLrv5k9AwcBQd5YDidXk74xqzQ/acyOMw5ZHr1F1DBqznDcUEcp4fTfhtE/fR
NFh8P400UpTD6RmUIITPbDmL0Y5UMZrSp3LehbGqJaftV+1EzAWiSJk3ZAB0+rB+
8a67zcnpuEtMN5QlClWo6uWbSlub8lHdNuSmW4I1dyn57x/VXpxBV9EdfJ0wKt5B
te4zuIcZIL+i6wUZMJj4G+RbbKvdpkYkyDfDoKNKdBfgyV9gs4t+qZbG4qFj4gkp
6+t/tcPE77HT+dF6Dj06QgRZi2FsheuMlwTqKHEg6BL+ZFPc+xl36YIQCiYS/8/e
nCxK08NAcCs3mptwZXE9RGZMeOfekufXCgHW9mNIw/Q/bqQTyqXshGMh6RYzfJr6
R88rjB47pPfOeJVUP0BHBk4do9MXs5tJ1Q74F4bJ+nxFjQxqXPsFhoH9G5oxjQ8q
7wK+SFylk2Ksj1njD6kAf2j1IAiyF6ZJvgMnRmE+JKiZhx63oK2EF8aXCAO3J4JT
RtPMSeYtMWcPw6VUhnERFVQeMTHMDU6nd3REO/TjjdcB3JFlbyCPlwktAsWZo0EK
LzgxczXHnUeIHJC44wIITdOHfGzuV4OaM51Sc8UiOBdV+gcmSiLqnOqJ7w9tW6f8
KIrpW2YmZEH1ZZI6o8pLfms7ufjIS62AVxtwzx+oC9kX/N+vZa5XlPOVu0PjWrcI
Wwdu0OJT8KFcjC15LwQTx7zSDwcn8uAcOifiiJ4AUAqz/cWFcjqSZszhKXw4Hu6v
vbqhdvJ8Bahm7luFOEijgsrRUfFBYcNs3wxZu4vUTDKq5ejyYosgULEE9B7ie0vX
XXY5KAlnX7RU3WO3b6O9U+XorYeBqSxdvRoCKkOn/MHeFR4JAoHg+KAShji/McNd
hxlH7hpxiAcDXpXWHw155E+T2BQ5AXEegz7y6ovxu5V57KCSWMepSqTOi4Xxervi
D4XWO8Ef7uS9cJNCkGyjSo0Pf0W5RvnO5PD6cYK9YdRu7OjgVBPBawAal9j2E9+o
nUjq+mL0sUzyTSwIReCi0qqGnwBLmXKVtXM3BxGJagyHue3kwq0DNsUes5pybx2z
JbOWhaCUmxs1tsT0MngqkWGEMqGe4Kz68bmDfZr0CMbW4sCf5uqqr5arq2Z5tnwB
4Sy3GGNN74tlvduR7J+VY5wcMV3huyk17MRiLfj8zh0utzLB9t+mUthw0dotjMpZ
snieFymHrcUdi9UdjZluO/z5AXElApYwUzQcdQbt7auuLfLb3uvESGr2LvBk01oo
2uMSp+AdY0DX5G2VRGdD55ku7g98lXPvlp2Vlvrp8KhiLu0uzaQwFldQPt/nWICY
fTa2aKGmf7dI+nqEUkh+a4PBD01feBz+mLbh2J2r1Jj4VrW+V7FAhg5+gaLu3XfM
xdVXu/Gc0V2LCCyfyzIcj3HzftaKyXpIgi4Ua5AFOIK9lfCt0Qduu5ekMVXc0FB0
+CHtEWOY6bthxJdAM42t6btaNXyC6LMltFge2TFbVKPlKXJr4roMdX4TyESU66pf
p4vmF87/QDj/4bhu2lVnL569hUNUZRwC8r+5pG7OJ4qBoDdKEvLPGlASD95LvIRw
7bhpjtNNIlAWzrl8T8FZ9DC5pYXv1/rVNSPrjy2CYRFL30+4zVB09u2MpXzxg0Gk
8CI/tQV/uBAkz4gR56n+lzOLB9RE6dur29cKBFziMaubcFkKh8OIGfHEM5DLr4K0
W7obyWR3giAOQqY0Rbcv+aHql12FbGCf4EhXh+NATQCD5fr+EUVrgpyATk5HvWu3
136rsF47P5czcWSH0qqm4988LlK1dTWjxzCEUIkRD9tE5enNCOhl/kyjvSUe+oL4
RCn3xkzFy0Ig+XmtXyG7R2KmKWDKVli80htAxETakcPDBzkpGxN/jGaSoSn+QfSV
buYuVk7bBKLE7Na5nWJOCGXQw7gX4GwPqhfTZEbCQF8+pveGwhUvLJakBNhpYYAo
AcninyBKJoAAGp++0iF8665j3C2woqb0ZB/5/X40np21bDLPuAM7RL6HSuxZ3nQ1
BdMf+Nrm++gdwMpYT/K2Asml4OxHq1xMu/8yuo401D8ueEXz6bDx2CJpYX8+Tn1x
dLwIoaOjcJlIAYWZz46thHHpVlvD3CG+kw7T/VT5D3rQgIZeveIIPspORbsZuRji
2p8gRoUN6XyEkCiak6B1FvyomzG8xvMvVAuUuDdikNEQ2d7/z+I9YmH3BR2DpuRb
+lcfwSomlBnnHvLurBiBSBd9c0L5r094/2CzyRvS+t0pRowdxlf0g9p+9Q6tV+Dk
mv2nHetSzsWQqj98Z9abPseiN4B6rVGJfyZt4m7dV6NcrG2T0psZpwdBokX9ECAz
vgEx+k74kh5wpactG6RL5K3hipsWz+yEhdlEILe/rMIGod2mZh2SUF6oM4Qgh+uJ
fBZfykqNC1JJLFJGXnxfhw6zHPYL4aVgq62RcNLIKuZvgWUrxeyb12+RFdysiCMw
SJ3bHt3PTBGKL34Kn+EBadr48rp52D9IQ052GX+uqg7Uyhf82p91Xe+lGfeoJtRM
Ziq585fiAjhiMgyzhyPIlbXUcXbLNhUPuA7dLGNUHwNMLh97RWc5ZLlVBTs96HeK
BH31HON/5v0aeEFbgExsOkplwhH3TVxR2PxNzpXNYgiMijeqUxZ29sm6Zt1aX7JF
ZdGTAha05+Xkj7U0PwyNMiRPoeNNYM3f0NRs/Ujrfb2ig/EqjxsKo+7SgNtalTga
vevdKFHHY8WV/EFUOfUuw41pv1Vrvh6m4JEkWGAy/wZ5XxFZpe+o4PwbLBnO0kGI
+LHbnxCiodRvRGzB3kHBJMMx/PAwBFlJEml4pJnSDrcaVIdYkBXc9Mqf/Vch8E4O
cenC5eWDizYmlrkMH3392ZZ88vpceD8jYUSXHJ5ml+3QT/Z53Btuf9mWF7wFyuY3
ddAWQNuzz/Jqw7OA1CxG8ify2e7saY0DxOrXtQU/tPsbRJ0uds/3ARq37ZQZ8Bxp
8pKLgZOmNQPF3t198oFxRPzmVgAwM70OFhhVefdcKvUipMsIDqjygsxToEfKeINI
rhBIHmZ9kKwp7nvV4t+DzPgnPCnhUOgavJaJkUAHQHskOiRXgXaNUQS4ur3EM+l2
qGGCMBQ8XCXap1OGBJtma03zx00ZH+Bjm18o3yEEiVp8nsRBaNgdHXl2i3DjnWFx
YH76vmuZCH5eMfOYpvrVALWMl/18tyEjyUDnu7haZkfEik9L/YBoqseaD7tjrZAr
4C37HhaSJKLdlxdJG0kXrGuEJlyGrnLitoMmR9QiR/RYZsMDUsFODMsp7p4tgN4K
DFWUsJFNNS/Z6cIxhFZYHalRHqPPGvs8vbnV3y5dGNA8f+Pou92dul0vxjydOa21
IS9laiUn0IDuYLlJZghALMZNL8TjYwoare2O5NzekSoYx4MEsDondjXdSiRwPaBf
LToCu9lId3s3FClx/tUd1vgVfmZkvOYz29DLPyoVWn9c2DzbVgKTeLvKciTOwH42
r8AN50i0Pxsj1edJnhM5bAxK9lwDEXKAL7aeoO9v2vK5WVA32aN/PZ2LQq4PgHpd
QYWJ/v+ex9V2JIegQL0DP4o4fycAUelP5fyngzGK+wCsZ4nqVAk71Yf1TLDblRKh
wy/qqLj6nJQXPQWEBVc/ZRIwqCJs+SiB24YfpntW6q3ab2K2BTXjoiuKbPppL1la
XNTHG5kDcfPOKX9pbhWqktIJ1rFPWm9dEOahNd4cR95bGzgrNfbAkqlR/wvGuk3W
67fg5mWmu7I3JAdVneULw1kCrFvRHyEhLJGUx4ys1n4I+hKyLng2AvwO0w5uQ/GC
EzArHGO8cdm7Efw22Y/qYJBa3cSMd7RLwrjcLd323yiy1AqkdSJX8awhbFT14M2n
/06MpFAnRpLIiiL6DSkPX1V2LhjiVoxPZyzwP5S+OS7fKz8eZBOYDYwuYd9QOmPq
V6SBNk1xTZpi7y0ZRMTJMN1uHOKznARM3hrsxH9cCj48ReUu1Y8dwusZpNmdOMrA
8H4b7Q8smNJPLrkVrBuW/3WpbOWnR5B8X3vzYUE57JehXiFlIRpkX++ep8dZzlc4
lMh9zXlm7eSmjGOeC22ETEhqFdhnixqmjfkJRSnBdmqnM1DrTIgxhRR0f3OMKbPe
zSOUaED+sKgmkLL0NvCVZPGu96RnZzjyX56AVWnj8T3k6sl7Likqi4BN9yZKPUvP
pkEl5rjHGcwCpdaiJHZ+6IgnccB8eVmfASvu1LRJvPqKXqCSbCfLrdfHhNEHrzht
YF+sYEs6PDOuWdinT9FnW3uGw+xipzD8lauKwJkWPg8FFny692QOqELVVBiD2C8P
pPn0ojimHt341nbF3gyDsLmjTnHwvPhJ3Gzo9KKRmA3kggxj3Txn5hhjlZ+n9YRS
8U2G2qJbfnkQHOUq3jHtz12i5mALa/yRcmpQ25TEiL6N2GkI//vTHkwVeEg/8+vf
ZUxWtYxW8iYgdg+BQ4CvpvjbggP0SmO94csA3sNk9S1fj3msDLzfoNZcujKuOTaa
Ux/lGcwb4W6kk2NWhky13TlH2HUpF5GWWtIigEj4OY7Ewsunxc+7ook0/cUqnbGb
BHxdSgnUmirE1Jkfr+bRc9sSXtDrBkOfD8WqdBUhY221FY2k3C5R2n54elc0tfIQ
jq+7nl1ekT4iks0SOOD6T4vI/17W/tno2J4sD7395X+KbBMjFfCypCmpaiJYy5UQ
e2dVuJh3wsyblTMa8bgvE/EcnYfEKFnBzrUUs1RSv4dNnqZKG6O9/2DXs3WBMQXT
WZDMYYQVl4/WEcOlwgzfX9qD74hM8MzoryXSxasHu9+pF9TYviK6gZI1se3mj1gl
Rox2kFRzVRmOnSCOb/exCZwOtjCbNQuWC5w1Wjvsqu7R6tx8TwK+0OJFYHsUAFpg
P+dozHbJF/XytPEUsgn4YM5ytv/4iPUXBATifKLLqogDhwYX9TG27LTeDLDp9yO9
T60ktQ5R+UlEJZaG2pltVad+3Wkh9KS40ByEoC3GRkPhga5+VuJ81oZMasFc2ghW
UG/PRntaiR40xEpO6u9Cred7kUHdYXCoYZsAmuMWJFfe3GJEw9xhxUHbdQt/+ufi
jNCbKnj2t42pJD4hOAjC5T7oZ/qQ6SbszLJ3Z+aWs+eLfc3lnRsidMzHVkNE5pE7
NLRja8Wee7xjMvmWxUa1L4H0r78bLJ7w3dAk+HxOWctlaG5sgtEpnzic+XpOZg57
7X7m3KOTWw1Kzjw55A9Js7kENV+3B3tiCcimuKpnVaGkdqNl/hOH6DCv+rifANT5
NW0+gzp2fX1gMjBKhdcS70PlT+Ur/ibI5of4j2+VksSB6GHmWcIz2gJRJhvcKmPu
5BLXw7oim5TMDuQoUMSdNVZCUSKRDvP/leBOPi7J6XrEbsVCnjPUjBuwwmzSFfyi
cPiFrLh5/O/SK6pSCFk1qgbJKIjqO7vgO0LmDcAMzyg0gideJyM4ExIyk1CkoW6N
nKZFPnIa8rFtjMm2ZhJCtHWoip5VWqd3ERQKlLoBS3j9updo+//kMT0DhRRS5GHy
8IPhL1cYRgCuU+mgxO1ZBe3IGk48Be8e2XMucSbzb2ftM6Qank/0do3XnJ0WRrxu
YA2zIrgoVZrU/0bk7W+3bcUngtHjhnpx9Or8grn/BtklyKqDWBQOz0cAqZr28+Da
3YOA1JQKD/XNn/XTNZzjmA+F0dRT0HSi8E43eT7xJJWl6cfSlyqT4FKXDrVLmuG2
dqN49bl9//x5y+WTPk1j5GHksKXsuQErRfSJyYuZ4+ci57qYu4oZculUvPZ+Tx46
WUlWE0b4SKkBsUsVLLJ1M+cUA1Awt+euVmJIEIKaHqgPw39vDTm0mKQxwJbBkk4M
X7LX26/PKcWibUF3fq0JXq6WFnhDIIMVp7TUZl9+8dypbEnt9+95m/BYXfpY7yOV
4Ra69kZCPuVWaSfaiX0L7YbGdh59AMCs1H7gpxiBN01vecQvemYvJOUMxqTyWYMh
w/ZDBrxWIEC6tWjBRUMrEMDdV6wuBkqylSKL6wLpO0ijzU08ZO/HIQMrvyKqJf6d
5HrDhtpFQYQjxZsqbHPGQcaeIs15tZw2zg9hYRwFJ50IkVIZ1Fc+JJXiwl387vAi
Jde7ARXttajj1jeVA/0xVj7H1ZnkhYcE6IeOEj6O2KEtKAs7AgESQElY5IOaVVjC
8JyogeTa0vgGyNjS+zuafZedm6ADiy9X7+9opNp+o0cjYfdhVpi+7Y7htSsoR2pJ
NXGdYEZOkjETd4TVlRA32s7geDyH11jMkJO5pAOKwkm1rgXtKmrbSWJiUSlKt/1c
PF1F818fCq3J1w9eF5TGf3p1uFEiXIMgTNBZ4yaGVAFB2wVqjjFklefHSAviIA/g
ZXcxdA4mtsQCkDL/1kaB0gjK3o5Z4C9NNElKDyNtZ+I639XMbnO49JAwEP1ixYQv
0iqnl5EkZd6TkEqKLIeQmxjoQg0nGrpoo7N7/03Jrq8IQDpaS+l8x7k4of24luAi
UM4wdxHqJSSCfD1Xj5bN63his9nX/IKLaZzwdoO+6R/NrXoPDKunDsvyrOKD4Mdf
/CeGumJxIMGfLpzPg6qeDDU5aZIMOBssk2ZX0/Yu9EkSIxLfJjA7MIQ2zR5M93jg
gAgx5Hdv8GvsZDcBcv4v85PGHyUjhEo2gsVKAaTXnyUJ4p0jdB0pSAA09U5szYHw
O1JmIxaSPLKrU9Komps/PeTwhzkAax4VYs+LMUdd90vi9dcXwga+Hc5yARzSJgYl
OYmnutizYwMDpjtmuRO1alqNXKJnkInzmfbeCiCZLqtk6NYJUD+gkEEwQveNBcf4
/Lq/epl5LZTX0AGgaUzqiX2HAcXmDWtIJ673IasyONm5UxC2BA6JQAHm0EoPDKuG
G9dx8KLUNvmkF9nj1XAt3wCYcMyqJ1pzBY2xcI7O+h3BpaBVbY3O+gA1dcSwRykV
72t/TCXaTOeUo6r85KbsPE2gPOF0j0mqAqMuggRhMTkmgkx3jQ8wrEpClc+lmCOQ
xmd/tMN80dM/LTMnzBx3FQh+y7b3oCldP+X0HvGzXrMg6fP9NOMwGw5w5ozOaDw7
zyto5CcrCl8ipuaIW0aI1mEUGhLBaV+RFNcM9Ls/Qu7jQ2JvC3fHEAUX0LMW2zhr
dgU/1c3bh3t0pWBrih5fetq7TZR+nb04ImfPOYA4iwVIx0UE45HVvcspb1pECPks
Zgz0CDDms7CXHDPFiJAlQNq1bNR1p0p6HZMD693H3ZmEvvU5o3luBHpZM6Ml1Q1k
LmuOkQvXUUbwkzu1efGXBxXkxsdV8gz0JxKWSmdy1g/iy+hGRd03Q/v0W9OT1oEe
NVW3X8bsehVBP108Cj3lzS/1iOR8XPNM6w4GBi6atuNanvytyQRru5pr41mr5oS4
fzrHL5idSlUIcS3QlXIqkgu6Hm8uGbKASIwEQDn/h2j6kTQCvxOfnbPZ69Bbt886
tQ1QxjSCep+0U8STjgqnO/q3rGQaDLObMbdXByN2nmUZO5o9cKCo9Te0u8RB2Xtb
O95l/TpSQXHwn4axOCu0mNBCaNXk8v3DcS+wZy4cKwGd1Ui8kQJyDMl+fMU2lyE1
wB6uU5xi0zBmgyhYkvNfuQ/ytNiGOOUjraSSlSUZ0enzHwSDLrN5VZs+Wov9S1iE
LHA2oKogywjfEHoxgyXedFfbB1mfHRznfOC97O1tlbwNS5ydocFoYPjeNjozgu3X
vyRiGmZSaCbim/vkVCTWzP+K82E6TutZovm6GBPT+vw6xY5TNqu2s05rIFQ87p/D
fTj0IgpytZaoW4NimfVPDRwvN04vQUFjCznfAQAGm4s1VxkYpHYuTpKaWrEbjWLL
hvyL4Sjjr6IctEdEoreptdu0MUbwr+zNA2+92f25lffFQD6Wuobo148CzF9ljMeP
RLxNOiESzQpuKtsI49y3yurfCM1Ftvl0g0eIyqZ2O9fbNU2MHFk5pHpgcR1E/wQ6
XeKcCQMIxlhVd9cHCPkQYdHXaGVeAAuquMfk6EGy24s7UhG82Gk5UYgMZQ4f8dlJ
NCI3wTf0KDvap4npPrEjWZahkYng9oQgiaLIRTO8HS/rNzaIAi6nI+H8ApIYn4xE
SkIiSBVoNz9AKrR0HAzWfSiuNhkGHyTBOrVEyk4We9Bh20Qae0v6q9xHq0/IbMC5
Q2Iemf1+aEpxCQIFk70EdQQcG7VzxhHJympaALmYe5ZHlTdkMYxDhBFv1Q3ydPMk
6d8NmkekR7tI0ISfNlnPFDI75wp2boslpyXXxV6wrhCYBmOGDF9Jn3suKKcWQUMa
askC5aB2FVIxKRT4EAHRpcd/8ZESAKDSu2+KmpPLGmoCPCQrdZNziiEfXP9pX1dg
ZfzkhVxzTXaDZ73gpr1V1EjGTp1SEB+oNX1Q44lzvrLpjEkt2FckfSp90il6wJrU
NSPko2N61udcuPkAHtUNrqRFB4YGfLI2LyEs+zeD3zCia87aQ5V4b7AWGP8C5r2o
u4EyKw/jYMhH4XGlxsTI4FhqEi+/McL1Y3eKDXitP4LTpED8kGwH22D5zCuhgZQ+
jH2LglqhYcT1Nqg82iIWjivx1k6B6CMv9T3kBWVk1CI1Ve8T41mP7KYCqj290vhQ
JiR7XFa2/N78MYX3H5b7fbZX64Q1G1vbzrChouGCaBjzovlARPNxLT6mnC4+81n5
xSDZICpuXDfpigdb92fvATT5F/GtibY7HApJsmjZvsznaTRHjSGYQRpCC7FjqnB9
Eud4hEmuhv5sniCGCYSWG7a+eTryxUbCspwHAylr8UuxdiIpOLnZJt7fi38T69mr
mU8Pduulk8Q6ZEkVaeoCHYcr0y4XV6EcOVyElxkvVMZxIJZE68Tamki/qzPFW3Xx
bEJ3dS3Bc1apAhu23mZOUsQ/iVXW71deNuGusUz8DxirU30ftU9lGGDQXxm61qYS
m1jIu97YAJp310QElUEOU2MCaC8VDSq8/xqgIEXMpXHq8hFXx+j3K7ERGkZmnFZf
qH3ttAwGM2HqVSDNVWVIQlN84CdnYPW6XH5zmC7iSG9QlQ1AsZQcGqXQaPV52i3e
GWe5oYS3Cgh4TbjxYZYePYmpDHGVxaPed0qBXyfzHG5x56Dzb+U59UqPhOUaxEkq
wg4SEPiNGZ6tkejDpY3d3G/Nx8Har8fLZoJE+Z0+FsJfiOvM4e5MrC1QsQrKokRC
kPnrIBW5XEOdgGNmkjn+lv0MepindhANC0hpfrrcdoqyJjAletlim7fn8IxBTIzm
N1ZDcxz7oklUQZCPXoI2GADkD+J/92jGs45cq8eS2ZQuuMkm3ibuaTwfFD493USW
NxE91S524DASXrk+2ijVzpcPkmIVHtKjzfphpNN0WzxwBcTVnlCa8/DXecAxMlom
TqIidL/gTfIRFhTsrfdMcvP12cxmWkh68nLSheNvl0C41S12bMFHZbsW79AQk0sv
aZJnogU6IpJco/3mWs5Fd12bfm8FDGz6LMTPv0AvmHqQDo066+ZEpT5Nqc6sJ5YW
XA+Rs6mQHhdgcmXdz+3fSEuSytdy9BSEMupNbFzzDNxCgREp7MMJdT5HkhM5v/4Y
ytbs9KuHFC3XWXH84FFnZWXjh4xUQxowDa6tQ29JkfRswKAUZYFIwgfU0RBYuIOJ
Xb0Jsu4tWIJ28idf+IAM9CKraNsjhTSHcyndYT52I/KXUO7x40ZQbUMqH5EjS6ra
GWKssEky1iT2WT/tvlhp6AAUklmwiV9yJIMnKggxGfUc+D7eJdvQhPqtG76O1RfP
SO9LdaWvLUc68jJjh/10sr7VE4n5OlWVhtA7544P2V7Wpx6NMk6ousPFeDbaIiE9
4tXWsd6aH6Fm74O9XDXHGDvQCB4fc/A6rm09I1WgXaxLbAdXvpaROods72fgLnK8
BAOU+pG5PCEcgDwKBvG9Yx+2o2Tfd5Wnopvqe3B4WbytFQrwSSxdyC3xv0/fLiay
HlmkZycNVkdWw6bS8qNbvHsFT9l20Rih5QIqq/7NEWPOeyD2eP3rrV8DANkvLcoi
8zYY005OZO89i5uw4t1JrMP7om9aMmNXk5vWnDWCcvc8AiA+bji7GMnch1VyledU
p480DGeSZqUYhgtRzzNWPurPogDbLW5XCu5H5Nvm96UprX6/w7V4vHFNK7mILvvM
pOPLCAtpyJKf78fzuumrxip2X0ZJRnBvYUDoDgCl1dXx5UZEP0Q7lkB6yEpu11TK
2+f1XB/OT0kJ0knMKzDcDF2+kZ4L0CxXSXRCmkuAV1J3NRfchLZuC8Wz2aiK9N5p
MuW9kyna75RDrMowiYaU5qeg86a1yGjJBb17CXO5qdDcvwFymF9Igz4mwkoZfAL5
bQGmjxyZIF88YWfX6kFKXBEc8S6YFMoYXH4nOdn43nLQY4oelpqs2jsjqavFDE9x
D56Yn88czM5KPqJ58KfLloGEzBdXHdRfLyDIAy/nmJN+jMP0PydlB0vxAWJhJenU
6xRCIgR86QP7NotlxAwncPmxQMBuGzaI1NDzV9fkm0y8CMtxszX/3YaSFK9ti+mt
uLmnpOxCJ2lFo8GvHc8AA09+eBcrJV6CoMkged8kOUydRByVEyvduHY+E4AH+SwO
LZn7liFQxmlXi9TOA4sTSOCDymPzizxQ575hQWndNVjY7J50OKRgAHtgXbMRdYgh
IXhc7t3vamTJ2PS7lzYuVKV+4zQGlUu5O5G9B56l+dEFnjtWKJNrDlSWINI3SOtE
l8kEGYpw/dJ/DPwlcVHLififa+9Qr2g221Xp5O79zRnIQKaAA7D7WgreQp+Tmegm
gumb4LBwVYOzii3CrM0y5T7EuPXWEQ2VUEKmO6n7b88vhsoeb0BxZvaImGTp8xfz
GlUkYcMT+BOgM5KOrpfYxWlKdqLQo5Mo8+qn5jkLl2SyfhhEDWcyakxaZwUigTRM
0pFIdSEeonAHtFrUCdIkh+YzAKm2wdaTr8BRi/c9H4eTMz9peK6PAw/I61w9iXak
pGV2OlnRowykEJN4WEBT0x+964+dYkEcqXuN9LNyjh44pdS7AF8X5AzncGsW1s/k
f7bJnAMD5XDnxg0RalgEPbVI5JxrHp18UfEa9XLRvKch8Lhf2LMMLoT/mk2Xiuwo
6jukU6TfGXNhDeCjBPrK8TnfsyQUmlfGdOG5OOUl5oZtM6u8pD/GpQ9FN7Q1Zlsr
C73nnEkzK+Hae6AFb/Fc/4qZOMqWZo0HNEtVYQtFgPuEuJHDx4MSf8TouHy1L8Vd
atOO++qtvM0NdQeqzrT7a78hgClTBIb0lJUNyIISFy8taKhYivHPDYn38YONIFLZ
3M1RP1qSwkTGIbvoPS6iU4/wYsuFIKRjlMX+E8SLfJ3RmbQcX7wNpAjjqRETPSlu
FqGYuM6dE9sO1I/DEwGjyXBCdUjmrs6Gdha/twJI6sV6p2QA25zCV9ED1NqbkJQ4
7if1ANFwqaOkraggC5akfgiL76mgMrxtxi0ZKrQ8LmdlrDV1JS0Mhk0x4tKD+AjM
kKlKR8oxK1rngq4Hp7SKirvRDufhdXkpW5JlWZ0rGehTEWyb2p/nQveNt6OAQUyq
DV1yJax2Jf4S+ovrFzb3iZWgvF7f42MH4F2d8Ep/9NGyLMrqGw79nSd2HOiVCs/C
8qn++D8nZoWG9pZ00tpXK8OgWuJLkKPCCvX1rQhbie/4Xytc1rUeiD7O4H9u0igT
7LYkLpwM7NhJhZwcnhuj4uplYu7XLWA9tblWpZ3MrIa0KqGFTz1oMlP+/cpgr4Wu
8XsaICvereSCg/ed7LFaB/lfj6KpnhoTlsZCM+Ojf5FdOIFAjOGwG5zR7YABYFKS
XpmxwPpr4TCVZ4fIBv3O/G6wnxFCxgz6a5YRdoc+As59BKCExZ6EkYBUZd6ws4ni
DqvAUW5vc9Af/5W0WU+T9b6kIVAt/2Mf8dTntcgBRJNTat7hQhA5Zf5u9lkclot2
TBEGiTRmgrOnuXUk4GDyMIkRlk6hmo7qtUS7ErHst2IkYS7VdF2qaCSXXLVKwIgx
IFRJlwgmsNzHK7gqrtfYZ0dOz3tYC5D1SLn6P46plwi3yBIiRd7TOSJlPGUWq/Dz
LOBw4E3v/4wCUpph6JYc2/dnzi0pNcMeTcMmJJ/FD7/ZAvNUszZH9K0ZToFCtj8c
dNi78sX12YZg0LewJQXuqOjPNyfMx99YIk0Z0T4PfNUGYl+bW4DffautFfu3jUry
TtxKxAqYiFIFwvb2xdO/u+wEalYUYAEJzSsD9qludquaD2z/EVLDW6x/cdVardap
eRF71VZJGmNdADxO79YmJgqj3WNrFEE+8yX3v4xL/se+EvDPpZO7EET90gLeptU1
2yiad9bqu2XiwXBROQJpu6kF7RnoaySeqleQUN+1dRqq/ZBWvZxM9OLAWVtT2D54
JrrwOdURfBBDClgfV9N3KJFsl9iO30TQmH1MHw4uDMIUujkJvUz8UGbJPTNxfBCu
XmwNxOJ1ASWNe7EcIjjipZlZjbiVFOpOSb0rlsUuuuX3/KFnI0uFnIKX1Rc5IbNG
5Bw2zV/e49jzbBqFRvmycTyEj1IRFiqOhRs/2iV7VUxHpSo2merquXD1henqbk/2
R4DQFvumEExwcjaVGHwjsr3C0DR1H/eV2jzpB8XEptPG1X3wc3Wx38/k6/XBHEzc
nJMvYxXgtvg84iL4fOpkewQcRLxEktxJHbXjsAN/SepORxbV8xNICwvPfZQ6pCqg
DkayLqxSvdYiXloPzUig7IEK58JRn+Dqy0wVpqpRXGXrEGHoSV8WR9w20rxHLq+b
WvLxjonKXFW4ONAUnEiLUBm/Lm8UOx3y5ekmAcqU1k8HlMYEBbNaWZDcTowrJ4Dx
OYIUB0zzIyi0kHbc3hf9AvB619aV8wRM8cN5Jz473t3rvDgtJPOujjgw9Yvdmiv8
3beBO8hsr/QjCwvY89Q/zVQjhxPZoOk+cukWSROhFZ7qlPiGop4lR2voHAltwtAK
pn6jkm8YLT4NQc7Vcpi+Kxg8lUgqvUU4sFYWLKSaH93GQwWscV6DbuF39ts8eIN+
3mnJ8iYxW8KMbNQlRIzj7alx2/YSKzVM2uBdBO2hrWfic+kpU1CfGW65TMRGMYvH
FRarPGGW+KdZWH6SfBRyxst6oqxMvSj33QRLErRemX/6QXGfhODMxmBnZYukfV3t
h/by9eRj/r7lMdrcoYQUtR86GlehYnCaxVPlHkLdZW90cviTFw3q5ru1sHAV2fhP
OTCyl+mpl4gjseXDKsyMdxEotVm4CaMPpzl/lJmYu2dJeqdB+A8prTDr0PVt90E3
wbEhz8Yq/ZMmKRMki2MZRLB9fruLR5Tqy3mUXV8wzHMYNBC0eT3lEMywFqQIqLFp
OlcNuLghEdLe39uXwl4DKHvE90dJwlc0KrKIp69Auy8JzXXHZbFpE4wSN1SWmRA3
2TKzUnkNiYVRLJDxsu5jFZAMXxCdqyxPnvBgsX1jwuuU3pSBQPcMAY4WyE1PwzOG
B77dFX0WqEPwozVCIgP4xtMYhnoAZ+artebTTay9mE+//KlHRejDRCcqCOocvSE1
KmSUjiFkTLIZ0aLXvPcaeYPbh4dVvnpPC6clv6ahcxlS9MFfgBURYIV80gIlXwJu
IpZnR4d3VKd+h8yioxIqD00nzN+mnlXd5rIrEY+fHyBBIlZvFt4XRbVBNJDvky4j
IhrSv1kWJ4I/pERM/Wn5R3H9RXYbbLYZO3xtt/MJK7tM6HO/c22kZatFSPdo6lB/
y2aD5shDq8UO4msp/jfAqssr5HKr9ndqUNnE33Q74/XFpkOVVe7NeC5GiFKR41vO
ig80svn+clQ7AY8wTcb56ycVYBpTLnzCdWcX55eLWiWB8lhe17o9VKZ4Pw4pxecq
rQPYqCnTRm2gcd0jjutwGdWW3Eve31xfYV4iic1aoxyr6GbbPbC3VvR85gPssQO9
5EcWDeB1RJzOB8/G2HFRHuJWjozq5AF2IblWQB+zX0H1/NRUwrRd65NwKYIgyTEF
zJAXPDsC48NoKjk6Bfif46Zy+jUucBHACP6BQe/l+tRmcmpBJ6jheRUW79TRN4yI
dE7AYc5KoSq37eJtVTZ83SDBKiSRFAZqwzbqsmr2yicbfCagIY99KyvWNJ/hXmQb
Y3u3CDP5WFno6JKkPGU26nel/0cIL2x6z7EQUs4V9yBoMt/cSlVTHGQwZvKEVvvj
8eqkH9IEB0YKkIwz/RjMO5oaRNJ8yGkz3N6acLllagkWT0WowljTgXLyFzBZuonv
AO+UPWyeybaPKVdNUwOOt2BGFfpoT2A8WFFOEn+ukC7VczYAIW/mN98154X+paSc
aGWIacXQ+OHtZlGgr4s64Bl03bIJ5Z0TsGrp1ipjdT9kX4he6CDp8uzEM82AUyCu
LeRBP05KEc1mkELp2F9rRTPKEfs89OW1C54zNmjHQEShWndiOOX2L7VTCCa9ccyA
HLIOYpjrUo4fQGMNGgdpsWGT8l7jtNXPZ3Wzts7LyQmroKv2JEbOugXbVMPNBvp9
udf+L0CsHYpqHYds4V6mNcGCFUhf0BLEkeBsqTb+xtuHHLpHC7VSN7Wcq50b+bxw
ZF5xgUe3OKvx4guQEmOtuTuhbIJhJwAvvoJkGsG9APikGweDnem5oi/o+izgA2QJ
z3W+hmbSD09D87pdrc6RVlt2p2NGti8FEmANTB0Bn6u9DSnMS3r86i7WF4Cd4gl2
w5kYHd1MhSYQgCWA2lSTR6z1/GxBVbHwz7UgrJOltz3DiG4gz2lU+4EBdxnTYKmz
oGclsu9v5lYRqlmfJ+K5B7yNi/ikvQf3ifjIEq4JkRCS1axZ7xGPnfrmTn9WZKQC
z8d+B80sRYaVZ0hktgZk6ZOW2AvTdWSkOTmGBwNcRvK8LkEdNAoQviiM1w4vA1Q6
fvBzds9ri3EouMJUSmG3Sy54KGWKLPpYOd/XXcLPrm0fgTX7+nLTvjInP9SMlWIo
du4HtTru2GGgg39Ll7kt6fKQmus5kiZPD81cAX3ERf1vAjJE0R2G8yr8h0oTAe5O
LeCl11nanOIhJLFac2BHVsoZq8Ro3ZgwdTtOH84Vl5bJb4bsv+ZA76owm3pSohJZ
1P5cVqhSNszC/5iotSUN0yWnjyxxYiWfSBleW0gCpid6a395kgQjw0+rbo168gsf
ws5Q98Uig7USwpIPiOBKZaqrp0ww97LC2TVjdQJb4jH5DSmW0biKIy106s/vaiIJ
plfYLgbVVKi1FmjsFIYTm6aqUawr72e+Q18Q22gXYcP/G7Xn9ZF7l4ST3JFIO1fE
bt3e1PF5NX2Idz7kalUK1vuVFILpIzV56MuGxMKwLQeEixO/5Gmwpssxh78l14Tv
5Hnq7bhjbVG4qzfz8OfACrKer7HWnqpc1MyYoc93GptMjjfO0V8F3sa0sXAMQ9l6
GRQAHV6osR0G64RBTO7cmIH4NPu4dIaWf7hvExcGGSGYssEHvM2fRJlCSMv7V39R
eHibHeT2itNKl1LF4k6AwK0F/BTnLd1Be2+K7PxrRKl5EX9aFxE0VKHNAvIXIpAu
O6hTvE+n1sk/+79BgJV//AkxTG1fDw8xTgSGMOAVaSk9lDttJqHLJfSq+VEkhT7r
BP8ebxeoJ3ESPkzFsfpsW3+PwTuDWLN6aeTognqqL9GdMLOS4qCpDmGyh+DB+IEX
UFw4ebKlcMstxQDVzjmhwuQiCC/g1/kvM26OhQwoL4xgZxhdQ+qx7LBBDK1olgqJ
44UhDYn47GGbYOrGcFKJTtSohKFl6MVVFkrqKtDNDnrWMZhbSCH765pTtT1nakwA
i3horcq4g1K3HRTka7sWg0cUnvzCophIdMSLokIeYfx9eD6Cu5GAO4vhq9gr4Zhj
Ba0rQ7WLuY7XrowFZzOjc9rlbxqZiERwaw17PBVb1XXdr519KPKHDSlxs0JHIAiz
JyR6Um2WOXmi+3fWq6is7qzEX9bGbylnqsXz7dwVECs41YU/v6OXqbb5Vzqat3rh
hCTZnc5FJEeFFnnWhuOOEF+cJpY0/tlua+ZwflvbHiLOMBtszcxDLtzpDJVK0wgA
JMaETLDHT7VvAI3nylv0u/RJ6VEZx+aZDssCg7jAuYkyALNsSqP7l0M+eV5ciipm
R2HDcAddSsOKiDZjnysR8e2Xd1ZCgxd9F5yU6mdzB6b3+7IKKaGXaeG/SPHHQFIL
wJk2tMUIlnSKnIc8CeK3vZp5sM/oUMNDLwUU00+ns3uCNx8+fqRr9rvX56zW1Y1j
4Hw0kDqolJQDm8O4bXKci0a5XXqAkQlQzE+z6MdRf9p6EY0TTABg9a/RB3eKfCYc
BCyNNdxWsDfzC8Dd4U8JP1hE2LAWhhCIgevkut2a9z5QSIkmuHDrGe0w62yVHndV
t4bn5CLfpAWtwEUVAWILPah6kxIVThgjyCROY52Q3Wj9YjJJK38mPQR1gpqKbwQZ
Tn4qB2I/wNc039I2ViUGmNm0+e3TcQMgBuhWS+MHWzcuYIQoeXaWjmrMYt/qGIzp
DelbfT3P4xompU7lvzLHhWuBwB63SObkkQgTnWfymzM2c8Le6h20PHQJk6e6t7qK
kkfZ8olnX2RYRSm75bxU2q56UJZ4RJD8O4wYJuYNdHVWIlZkA+lUsFCRv2rDgCBV
CoxCXvMB4EMrMXMUk6aWWN9VmmC+DOBerrEz01HvfnISEYK8bwY8Q0Vd56V0Qe8S
9rxlboxW7dnzTUoV+wEOfsgOD3XmAsBTqZj/AGYFsH1jwp4kjpqKMaDQb/XCctNe
OL3E1YMi3fxEFiYFYrTJYqZYwPtUEzMdmiJzd3F/nQPCtUBoGIA1BtsiAFi5j5Xb
lLpLCy1f8I8emjYtfVjvSgshVJatbGbpVSn1ZLud1cFYiVGW/VuER8GLCdWd5E4n
kfShJVL83qZhxeGIqY+cDrd0NMCMwRWffioVUnPpTxwDz09fB/K67Vy56sx/vsk2
uuV/URnR+b3JQ+ye/0sSA2RnCzTAl+A3cPbEbtvvCe0sVm60Qln82ZJvcGMFrR8Q
9/BDfReflp6v5bfB3GCPfdmlQ8ROVibi7JWOwgSkOn7t19Teac0PIt6RLEkhzFa2
Rh4/1nLPFV58OmDyT1IqDTkNQeDdvWVCsxrOxLkE53U/KCn7b+MRY1OGh6lxF4uj
yZmuJNIjezkZ9guWPrbBbvnsKXFX8AOY93La0Wv/Vow75bWt7Hoe54HoS/fPRdzA
8ls8G8Y3TSy78sIPoLE77tSo2+Im9w86ODC8fNq7O3I0BhMr7l0bShPFwPEXVXHq
7AhdeB22hRQacxirxm6vaqLz1v2qiLvCVbnHX2PbxncpVZr4Yx3FIEte4PEpEAs7
Es4Re7czsQInz5HnebJKOUhCk0RMLMfFFRRA6NASvhmzenyp9sQCVyU/KugAMwnX
aIogcF6eqkEm4/nFIGmLC2c6tFSSsknpOtT7J7flDhsVv5AnJeeBBOvDxQm83iq0
XUIaJY+K2CfEq9K0HWpzuXM9rY9JlYNB7sawU6Bwy6iAkTcMY9N6rm2gBmCEeGH3
3a6H9cJUqzieuWPGHVxXkPMbMBytJ4RccdcbTpWV7Q0PYbxnUpnaWy1XiTwqaFZW
dzHTAwHlRKYqo0LNh6pnNMpH/G3Qglv/Z8QQ9KUpTCJUAoVVXAQ2HvvaVS6D60hS
wkHw5IHviHe0bB+M2ogWZ+gEItsTZ/9s/sz/PX8r9wqiEs6Y8yreoNevbbtpzVZR
1G8IFj6gHpo6ZqaeU/hwDzZcNqGd1iHjT7XplTerNBftEtniihjH1PbZQrSUf9F2
t7hJTkKKXxoAJ+qSWaNCCRWKCw5qMfekRS/oP2PpgxHyCH80Nkx+byqJh9ZLTs9L
hRKLJPjOjaSSI6/ivTs7P+IXXdwpkIHrZL+wmpa2Oye6i2MMKcpgBQSsUMWC/i4/
eguQS7kDT1/ZcdjZXWR63CCxVxHH6BBNiEW4vmafqfMu2yldNxqK1wHR86yLz6k7
8+whyifIRBdYyhMkfs4PqiHqIlXqPNyseHLntkRjZ/v98WYswVWdHLa3alx5xRKe
1lH1xU6nVVCxh5vheH2vqgMrUW2nF/UDPgiiSHvGzKCH0lNMQi9oDUtBIH2vTLsI
3ifLe5hAoPsBWMrtO7Uy9xIEKxGDbMZhZ/NVggxL5y3sGFSOYOKNV5SjtDkIfRhB
MPpUH+w7Lll8T2b+Esqyk2u/D1949FziTvLZ12EBi8qjr1Qqs2QKd5XcJs5egYac
HPNcHDrkyTO+EY3DUYlHJSBszPksgu0aqvEGEwcpAS8gGk5N0h8c+o0GXqbTu0xX
WN1yvyOu06uCP5gZHk9smdY2i9hSvYTTv/T+t1mFhktJEnQSvNRtjpEcNyGlDMZO
aLqlnDyJ+XUzuMho90jbqRVIBzRZnIIgsiEHC4dVLdCjpwnvcsbFGS4OdDf4gM7C
jXmd9FjzWhF/EMyUuQEMbcTkKYZEXdxcOYSvt9M0fTv0udNrL6btWOITjy4WcGAi
EooSc2/57n8+Ih1MeBTK2obIN3lrjn43z8l7nQ5ZIjGIb6s6UK4T94+kH3jSP5zy
qf1XX2tx8iTRLEOCSMIz7gfgxKqt4oa2K9Pqo2yBjUCDPzg3joGuk4u7BGwPV65J
yP85HzBZ+6n6CUOIhAbF0PGRavdHdG6lEMwHMUEtbZpKFUMbkWvPQHTou8GDvFHY
8ib35RNHKuTfiJLxP1PUgzYMmbw7pR7LR6m3Ed6yZXB18nbMroWA/Lx4KH7xqfwY
Xgw4eo/vN4adAcaJS6IuojNFYLYWcoJ73BFjFn7CoPqRXE3m7A4Y11Qs2/KcjPZJ
yfeYkgWBggT3yEz2rq4qgunn6G4rjnMSHnuS91BRVzU+kLQ46ah3rukZXR3aZe4d
RbUWn3wklAAmUPI9ZZPabz0aXEgFXEoYOUKccfI8G/Ol/vxD0dNcRAeMZZZeWFHt
hw7sYvH5UvWEZeY3PSdCKRZbtnTDHIO2amcOuApvn8rlU2dRTYm9li3Kj2A0U3Zi
vggzaQsON+RYME24SHLQ/rpaknS10MzvO1ilNr+P1Bid9d+rm23k5aAu4QCguGuF
S16m1ogynC7TWi8g6aZMMDodKlET6EAzsCSwLcSXQ7uFyz6qye6t2hhlgW0OUs3Z
DfF4P6kM2j4jBA0HkKtzS55fBvuBlGIMAQ/SkT2Ec2J8DatDHgyxjujZThj3Ovsf
vTQeArdARdva270Bh23PGFUaPnjcC+kgq77gNe0jQTZCJh79OxUmhSXwydHnzl+W
WxspKLCe4bkpiSTWH3WPDAzbY2C5C3xBxNWd65/PO9lqQDf8+UtCY5OKINPPcY0F
v9HSgZdafPwbqF9DLqYq4eM5rHjv0mCB1m/udly1D3pkcOD8HHa4GUBw/VwwoDqO
rJw20CO9V96otM6FhnYYyfrwO8i7pASmloYi7aY6YJUGLjaZANhjdeoxyXkQCoGP
2SmILptpuhnIL2h8OIFWqN+bW264R08zJBz33OghAGP6/wn749yddeEBr2h1snBi
hslZ4S8r5p6WXAuUX+MAWiQ6U7UqjX9fyrk5cERO38HyPkiwbpMC1HFTBsglD8Fl
OFbr7epM2NQObsT+vT5hO3fPRSPkg0b+rV4Meb4WPUKIT/wCJcSCJ5h6coRrOW30
1dcSg8F20hosqm5WOdNqf86EaS3UtkiIocZD5VkRc3L/2L3sHf9imNzelU74vUad
CkdIhSmEYckudDkL8V5Og3KWnM97kpn6Z6Qg3p8sPI1/PsXzupxcORFmMuF5EFe/
BA/zZ1bAXK7f5Z6ZI4ys0LbE675BJU7zcka+DwKyAotqFM4fUAczD9tBrx8GzSHv
YP3Hb/aM/8grqWQYgX5NSCcKvP4QxlnZ12sSoC3AIPsJSpFQmoCHYU62s5HHNRu0
bGs6uaN5FDqsHdM1unvEJQUcqWt6K75/AQ3lM44BXytXASp+R2lnRowVq+QQoPi1
zAPgUxNEuQ5sRjVkXjT8H+aJeT44H4szW3UKneId3NthvEV7oOPztQS3esQRsb7d
ELPaBZqqPSSg5jFGmi6keNapD2S7HG40zv162dUt+6/VV9avy/4Jt6Z4Kw9NpMJY
iYgmbK3qg22nmVIQHP0dt/YPUlziXM/IAGKL4O3ClldxnL4hBE4ndifEyT/nacN4
BImdlR2tsHPDuSeytX1BLvvhtvZP5ti0Srhzb+ApZaWhp1vyFAsv8bcVE3RAGP/n
5IYllcAOtz5B1y7+VAMmCu/RdASQxCAnCl6BkPPUEIE/SpBX/n39G98HkYyhkal5
YwLufIHs4cvmgmiNRj1jH+Tq2tvb3/q0as32xJU0YizLk27VuErg8ZYXeCHfG7kT
hFk79cFV6vJQ78EbkGtfSgUn1XCt/qXoLcOMPlth3R2kRJ03dR6F0r3W0NzVji2p
TZIJvoAjFoePUXeML2nDd6UZdaWiuB2X8mJPrl9P5HKLlbaKwhWglgAojqZ5D0Um
pimxOBm77eUKhVAkjUzbcpsr73klGnjOjCad2fJfKXQroFzF15iPVJ3JdANQVppK
LDcikTau+3Y1vln1O+uJlRUzBO69Nrf4Bd+Dj0iBBI3kltw3jlg72ouBCuPr4cP6
iYVhaW+022kg8DYH041LSS2vwq3GYijMagCn1UPwi2NCPePU/kle/KtioA2go+bY
8tFN6SgWaUBxMa5r0viuSxQet8R2Dk3FnZMw22GBpcMWuuiHgWmIwZ33mZsmRQvi
2LYmqkzay5fkTEewW2ASM4W9bgMpcuR6XDeEaKkqlesVZLeNU2tuyY1OTX4qY3MI
tHDLXP0W1Nxo63Hgc32rAmSFmY72Fygfh8rf8w9gll00f9w9RCNmujCRHoWDAU1s
kMh1BBdNUY3VjH0FtDDl2CcorfA2lShD9YokPY+moQ9zXrOgudyTNHdfci7pYnPB
1D9EB6t+CxciCgpHw8DhY7mVPSMjt/+XSFIZyuR/xV53S2aPgjfiThHRwgKw7hpk
knovPM87uzZjkBQGu1vYZAuw1TBb2n1B2zwtVg6RnillDc6SodvBSaaQX0HdqW/d
6YpqVv265QTX6/4/jp82PpNF2bCZJcFslJHmbXuJmclE7OMggbznhpP47242y+Ec
woy8Y3e+B7aYbJ5Ppni/unwj3JQSsv6guwFcaOxCm1NeX+7JdEQD3E/5goxlr8MB
EJ/2TugY02jiwqv1TTvP7vJjriXoLwJDD2JC7KGB+Gxe4cVFPQghMrQea7Qwkxj+
KiBq6jIIDHv6JcN4xDwvFsh7ePvaXC8WShRa/xAy2i8htI/csMjo07HVq8ER4+YW
pPzSPhagGizZuvwOSm9CCqomfZOVZqekJKh5NhmiLQIedgT4RJumiibiaL9BXybq
zmSJqz+gv0bWX89+tzwvXk01SYq4mrhscDlFvICQAoTzGHsIJrmDgEjds1T/wdNc
1Yp143gIfWVnG1St8QsdVZ6BVsDXxHP9c3a/BGzyBkO1zD937c0BKehSb3eLK8F/
Jt/KGAW1vjanq9xiUaAPCt6MNNEd28EnYNbehUnRYuUd1gK+WJfFE1k+D9d0Yp47
KnDcH0ZFKNWEjouV4Em3C+Yyt9Ige5gQ1q0e/DlbEHm8V3v3Oi6o00jB5finDLi7
yTJFNuocUoKtA7kj1Jj5XrtQHRIdwG6kO1qvYUAkNxCHjoEYWt+9oNGa7gS2hcxI
7xT4B2yhLeAmCFLralAcmI0goq2ijcdrsrrmredP5Vvy3hZfZ4MaXMNH0JeOWtN3
oYXCh3WaK/UuHM7m9OQvOwsd9p5gGpy1/Fqbi8lJAIENhoipDd9K1d5ui+kgbuIq
uTvfROsO1MRAUyJ9S6QusfDsWphTia9MreIp7LYYMPE9B62vIoxhSbUZS3ZUQKZQ
XLvlAhdLh1SMR6fNoB8C9v5fGDIhgNk832Mw+t+uiRd/ysIOrPbu6GdF6dAQ2ugt
m0RESa7dgCC/FxtfpqrnYHc6RjK4eG5iIYOMqTUWnW/QJtsBhlrbhGRHQAND/wox
dg6B8mXI3YHjjbhTGeWibzN67iIDz3YD9tQxyDRuY1vfcyjyQChqf+D7igf3kFX9
p1gpHX6CTva2uwx7c0cz3B3mqv6DTEl+JLYFigGD9hQcNHAXPzB0/u2s+hWsO/Lr
icHKiszeaCf7MkkHSq6FtL3etpXRAbxqqRFJCkm3thwPv5nCn8THCNbl44c7iV6H
aY231Dcg+Hlx8nHq7mOhzN4bgKeKUL3XcRaz1/cVGT1ML0MY+TiXgc+VPo4fETJl
7bqpX8DThnnJsoWJYkiJcS0+NDire314RjGAHp6G0KRIo96QvNBoBrfVLXV/YR5T
pseDFE5UsVor8y3JlALrQwNh8lwVMt+Pc/yUnyB5t2ae4EP1w0fsgiUzMw+Hp+iJ
XDCTbfL/iwYd+FBnTHnY17PLK6nX7s4DBsCzFWGSBG33zGc0iRsX6tQgpfqy8wFc
S98S4Fi2MfhGpMgSp5jQJ0yjn1Ha5dkfAHqFCmvAx6Qsx+eOO16Zx17soywOckjC
UsyIFetWHSaYIY+nHgaUg4HhLgIFGrzbQKB/dtYtRuXTlg9u1UFURPseCu9/T4M3
g3D1/kQBsAJ6tlMHb4J2pA/lTEKkrwAC++AwAqp3zw5KVwWKDcMRRu62uI6XnH7Y
3Hqg/M94Js1wPl675UL6Yb/lOLGiHyeeCKgDzxSs/FV04LfUXF1QPrKQ3DfDKFZF
cYihCSbqW0rDix/PPddaUhSWu2JZfVwYHecWDj24Fg/Z+fSQ27y1HdcSFEps8vaD
Ox6SJj4Uh1DhGS/GYfacBO0/TIUlqNZNxwSlxNCSTZZk2zfdsgN/YpMsIG/ROKrA
xlgQQgiVXLbmTr2oUvOsrx+Ym3JCT5wvUKTrdgwehSzf4u9MilIfFlhlkGBWzWxC
sQ5cXgr62cpVUzRtn9GiEnYDCU3kBVaRBLuReajDGDQhsYLYdeEnrgNRt87vtusl
OuhQKUZ7kUzLTP9jugSjXYEXZrhpYQ5Lh90Mj96wUBNd/Vp5XkLLro5/U8q8YVgS
OjmQ1I49yeQySD1HN3Cp8EpK8RHcq5W4YGg5gI9mEyZvCqu2uQ0XoPPJ+kPcsMbG
ONTm24njvABwjEiNv1003+PHpGsMOvW6VZf1VnB0WDMJxStume4PbZ2QMdBJYWeo
X48CHoVMqZMiMF8oddXVLnb+9kcdSHlpLX9q7r/wURr8IPOJSlWlyirxFB7FLAMD
FCy0f/kGpXWkQkBV+gAgtLJTCXjenO0gQ0jxHmmuf8WqET2lKoBsBqUup+ZlgQBP
EjzOfzyi4+qCMet7qWVIEpTC5lrbS7IQAEuAAIf6KPCjwjqgDIAN7wmrmqDCC/TI
2OiJv6PKI7WIOV9UivIYWvYxNagxBmTL+Zp9hZWkJeUjJbgr1h5bAs104bTBmzz3
c0rPHlQkMmXSTsP5RdvvZaWFFoxs7hLxtr/y2LxmPpWchX/mahbaw7Sh3KuMFc6g
wLBqzBYWNKIi5zLK5un+MgTqVp422rNyIWHuqmrDJN2ceLWfh4Z6xdmQJVqyd0zw
hSLMspbNU5rNqnxZHoz6hOB37mHPD+A+1doCRGa08gRy1i8PiKj4Zb6/JLB6bIFN
g1jWyOnUMKS3qORzwvAPL/meAvQb7VHWMQodmMQTu42cOx7QL9YIsfQh80WPoXzf
gAA8yClY2osKLWO3GvwzZGHZJTbZldb7iIKbzOyyUr6aIRf6gQDw4s7K23grwHKs
DqvUg3NvCqI5Uo00S0K+Cb+QKh2fqhxzY2FMTmtkqiJGfj/iKgKG2x93kmpxKoCo
94JojP1bbZE8b6bZYZwAjwssZtb32fWErNFUIN7LrnR+RbHy4GgDYSn8fWMQ3WJB
x+ygIJmxGPVCveg1si5Lje8SxLm1gBJe5UekpVwAM7JwXTYdMEUezHPglSt4pDHN
UAaJRkPbBkIb6bGYyJ+w+CoSDmLTDEK4M0US2Kf0MwS7IRbWgn75wlw2/0MWAD+j
+M9FeaVjE1FfDiBxDVsIXm1ai+o5DBhp9yMALdO9cW/lfMiEznLqxpUyz7BO+hjr
XylXUI54K5MvQ2fPl8tDPftcE4h+71unZlx6Ugr943AQ300p/KSccBpFMXZsUGeG
EFoINJFB8yRIcHjwzxKu/VRCYhr3tG7llhrrQicnBwWThPt3CX6C3HO0w3F1t62q
qTdlyX97ZmxKuF6Fu5D6WCYi0eRY8ky4+8m0aFQczzL2iYcjnYVRJUydZ8x1YFqR
hFtKn8LCGlQXw37ySTT+ENk0rMa6QBWYKrPNuylx99VGA9a+RqBmM2E/2eY3ekSF
/tyW6AXDfZ36eJKkxRFytjtCMnYubaNdT6Sn7U514UoRwbYLCU1+QRqiNJrJa9yV
IzLBdbHoQMeddY1dJaJOrhYCP3LAhBDOVGkGvAChGGAUzmxCdNDbWbb/QxpLjY+e
RZ+mTzJLf3k8hRxbXBBRjh4JFpK9EnQA5LEvio6E4vJ4+jobRtHSXCdg4KXNqaVY
eJpOpUPMmT363Vvc/Lw9tEdNqjOc0TLijEjOYGk9U+0ICONbHWuvRak1Ai8dRAj6
kmxPCovIOgIpJ9vK2LusJBOqMOZcLA/s2hPWmg3wIwRT/KR0dvHCnQfxFeP3btgr
zl2wvTdq4tz+BL+PASxTMPLheEnQ+arBKtTw2SBafmIQfc2QG6t1EwyRvg61VM6v
36+Iq+KPqh4r//B/ZUyyQ1XO4HHoSAcmeGOKLULhCKmbpZMECpuPw9VpE3/HgWdA
THSH027bONexziQg0zySoqPbnnu4X4Wdq9x06ikRsaJRd8nn0fVB66hEDai+OfjC
KZ0fqLOPE1GkQcXkViAATbuD3YxiLxUnPqLa2OqXt/MKYyqE/fJMAbYgaAmDMsfL
gSR+iPSOnLKtevleHwrTvsQv/RlnJmkgKFfHF/JyM3Ue+mnmPfgelrEA0Lv5+/rq
w5O/5WVu7PQhZM61xIlz51UPiCXj7txZMxbi9Oz+2RXKdj3ghEmry/X8ie2mfsDf
w3O27kCjkot+LyxMKerrLg2sZbm+iwq+4oG3UGRDRa/zFl0tmwenmQJvqwfHRqdP
B/1Gd19o41KIFyZTzPCnaiKppZDb2BJGsuNmZb1anZfagS3F3qijNWrPqOhxqddo
OAj1He1V7GzEV5ic1/CzaUUHpsYzVLMonL1saoSJ9t6Qga2O0lxlEBZIwbXF0DPe
vfup74Q1DQOti+7iXhiXV0AsIjmk6Lys5c8JFdkFr7x684BaNP9VgDJYIXF1Q1hX
lOpQkTusiXbllJ09h+PI3DdFOf4UoYvUHRQpB/2wekYDrUz0RSd0qQ0X240zo+MF
IQ1y6wfMJP8ckSHGTDSSuurtJXqcuVMcLu9S/+jmwqS7GHKFI7k97iudj7Mtzt8f
TT2M+clTGUPnbSWO9ctm31VAQdKNEEIi4va77Tb7VO1VrkcH0cg0dPgdsVlKWU19
OORGV0YN9A1yF0xmPBdypE8uQRevWWdpKupXkE9Qwp26cdJz3UUclj4T3oS07GWM
8+7crJG+B882VIfhvoxbXnmMfgm0gXhgkffjFlXz17jH0zHD/+j+foSd1sgjz4oS
uZASqFHsXKyDzvEvue/1frUpsom9QEs864wus52aG/CYhI3xDREDZqm0me6+W+jJ
JR3SJGQpinPfegaTpuZZ2wgBYGigzU32h7R8yZHYXWODtzlXhrx+MwNpqBGSkeen
+6T/TF0van2MPTsWiiMDLj9oWak9NAMob8BGosvJP5d5uYx2j0EJZYCpiA0maIOm
78bn6n/JV/7pK8yUWSUO/DypFl0XbOHB3ciPPRTulEFHRJH/XQCYYvuETjhSABTm
Hnz/fPPPtJ9YuhgQtmNV5oJLczcK3vISGdikzl2hYZIIOtf28FG2uoQtdRF2fNjO
waB6fqnWZQn4dd9Vs9sgqfmFsl9pww4QL2qpzC2tZR1cMGQyUYlbk24QCS05aG1q
U0VrpSCfcJInWprm6bbYn0F/yLK9t0ryIlWpK8f9ySAIQOVagK2hZmQ6HwOL+0/Q
AjmYfAyw/G++hUdJ6xLm9jP75YyC938KIPQtHE1MdDmTC5otfoUmP68aburRvP/D
T71CceXyOuDRslPiFu7VTNxbXWhGJbJTI9S7SM185yzk6lF61BwX5qsqNnSN0Q1q
FT3lKLyOTc4A3T5OxmvIPr/btZlJD90nhF7FPl0Q/uOyxKWcrn7iUB/5iT4H+afm
6jVbIm18dHDAmIUiZZxwZdTLpCraLUDacf975/vjGtuQ4x8DT8KCIrmNlF5hrZ/H
F+XaMk4Kd+zojvJSwLrnnzeM2dvRXm7wwR2zggOIIopxySzGVt4+tmTVyX43h1DY
Al3u8NaUFRbJd01XpcJFe0LcjtKei4yBtsDBcFRDZrQAY7ZmuxeHU7Rgf8gyEYYT
o880BCWlSsYVQL7Bs51/rSl/7KiWv/+ZQfSOgx9HLMJptb9OtLCe97juii9wmND2
xuTSPjgxbPHAoTg8yxetAokuw8P75ZxGDBEJuCCXTKLeqpIWOkEaKkXRvQrIHTux
GR2zbDIKtZeiY/onIgutZ6VXzIWoPu/cYJtXnJKJdMP0qEyoTIWjGeWO17xq0nrj
XGFssiWSEgmn+u6h3VSQ/oWUE6mkP/mLLtkuREqm07cWwVde3iSXLj5Mx5K+ZGSF
/vUM+g5KXMUK2m68A/CHYgm6KsDfQm+vIDHQzxKkaWWP+b+YdtfNLI7jfWldo4f3
9FGfisLQ6zjaiyl0D6d0ComgB0Jnqr83/1E+mPYVxorxWBMQeFFDC2gYZKS+7E1x
Kq+uXI1Jk62pRUh9R1rVo109OH1mbXKggrVbjivQZj+ZOuq7QzTmHNnjs2qb2MND
618nZn5LCRHx259KTMTmSzagp6+soazmFVfncftkdDoc+pFRN/dubGGlFAYY41oJ
KoAOz5PqF09tM3/aGBYlHgjUfA+vTgxkAzhJ1oGd/dklPhssQPBOEJO9Qr3UJ+Tp
xZsmBhX6j2VsmCckAvIFJZbujx2TfSqaeLsae0ZoGcLf8XeR7ZcF14CmzMLlI8jz
T/5eDF3xwWqwDcfxAuMiFr0X9KK7XeQWYpFaNdLw1AGbl9Dy6/EORRU3+ycd4TUK
8bH/YNMstGKAsYd2oTgOWGIeQNlu74W8SjhXPB/P7iuVv4cEbvl73y3+SgUUSFaz
rUzDSL94XVgCiJFMw3V3p44k1b4J4tGEEuQaoW2DLM9A2pl4ySfNwFjTynlapoRU
Rx0vLTRWxY9OVt3N4SaSoGo5Uatikls3SA8VOkYEVPFu4syT+C4LINMPmpicKii4
GhWHdmhFVgI7nnHMYS89dGDnNW3OCCQ7Q+14h+MnFg7bUyfRU7Y9/t0N0Gl8lJgU
TUvdCRwaG58p0tbrRGo80KmNiQtT5bZTTMtAHG2xTEYShJed0cKhGjtN3zyFnie0
L8bEuAZsDoV1DDBMsoIJbZ5XV/ioUNsB0+/PRhxjod7ST7EY8RXgq7U/DMh2Qrok
+MWqWaioDEz/psIYDfh3nTbgbnP9n8P+QpqFWc0Ija8eR1DL7JCVGnajdq78C5CE
qMYid3bOOVY0DxjdMwqOq+CZKJRWOhiDoFSJdyNOPXDPkjxNaErNuxp9gW7idK3o
oNQ1r7E/S5dn5zlwt9DPgxJaC2H2fcsfr1Cb9lW7hZVASIuy7ZPEQH6H564kN/Pf
GPCbVMQw2F+mTCLXrCQeovAzI4+PU5lo2PfY1TMqa7AXgxSqkx0AJBxs+72HW4eT
GtENYsDjGiHvEqBzmURYFq4gBaa5lEeoU4p1U4MjIf5m97GGGnDMNih7tfYWy/PZ
9vUXDv1U4N4YX6KPUBzG6MjJ/L/ClMT2fEE2J2fUmPrTueHMEho9txIiGDJmfsp6
FkHc48VwTcO/3aycmKJh63NG6xT1iYE6SuuZWsb5K+Qh2JE3qiRIsbpkTpcG8i4F
qIWnWr2V60m12Hj++E6GZr8cABCpd5r/hbZrookoUWeyCOOgc54WtDDSI0KT1sO9
hKIZ0bu42ALmH/MKbAqjvWViyJ8e2dgK26N/C4SN7nVwCtxxeEE1jhjkjuYxHe97
V6AKYwhyC+9HDyzg8EgVhaIId8215osuUedZD4U8PApOiZg3CAcCTvlCzA1kOTEZ
LqOVcYpicxkm6plUzWr2/TV2pPFegr1oeDNEBesidbxoTGd1iHu6CNhqAeNNnbzI
I4Q7bgwzXb+4yW0aNIIEH+xE/oV+/Qza65TVMdtFQIfjxiiIDJVjcaygHd9Pt6dD
3POJpALdwB6QfqrA2O3ta/gJNL24vU6ukd1Hrg8yAdHbachpWew42eyASqVO4yU5
D6RlvCna7srF10820iY67SkOUUBQ4Ih8/i6/rKYud4xmnVLyQ5YRCvKwiKMDKGDp
TkDTwcRW5hIiosei09AtgdYGMEqy+lY55rW9/u5QxnEl6GEiV8V+Ih647wEvjVUw
+L3MC6wsMOk0to3/Rg9vgiLCZtPriwEKCScfketivhcvtALLh2/5c1e+GkfjcmpX
7kqmTsRj5sG8KCAeQkoHyM4U6hMQoLUkJbBEwwTceQimD12vboH3E6xT4cpTsE+v
BVzTPSMRGYCLq1a5+fHifVQH1acarC+67iHNDjvjWFnLEufleLMtyxAkN9rgVyoB
S4yW6hvOTKnfghOhTvkg8QsnuMZiRB1jEKLWA3s+kfJQcYBCF1hhgH/E6iCv/CWO
gx8FXtPP2bhSyPSNGQT4ndH3UBtY/qa5sY0/ac5cKkLCNILz2nm42+dOC0MzRsWw
BiJjq94ySdUuIFjycmWSVsBGtztCIHakN1+MAhAWUuIIJBzI3jsusMBNCXfJ1VTn
O/lI5C4gqtpekJQC07x+5aY+E9K3DuyrN8G2i0gQFDxW9U6SNftmDpOMI+oFL40f
1qh3+L07UeQz63NkdnEVfEDp1zXXplcG+Iin0K0UbZaxieaAT57GGdWqog2kRb7o
cM69gJX1Knmy5Y70yqMVQsoSotfldOcjOgykH393x2dFQ7ZK75ZJP+vSVysDI8dR
8YenSR6YgftDvkdAg3NPybvtj+Mr6/74F4er11DxaJNpPPyHsMRNhEPSJn+xIW3+
teag3pXfsY93D4FqUJ9DRdNjrqgTPAduAxDnPvwKDc6gCZ60z+z6xgNZwK8bo/+P
fiMBE55KSiOLkxmZpbr2hpwnkc01oUfObPjGkfsEEx6Jm+aHKWVFjdCgqZF6XbMh
GIwuS4uvWGdyMJCjzBG0qe14qNB+LTVuRUFTzD6U6g7ia1WZP1RF2ESM2gX1jEP7
3LNldPuXS7wB5VTcCxUXaPYxFx/MPkfktwwk8Pbdj4Bm7aBEBrsHm5Fw1lwksy9o
V8jN0PbQuLAgRqn5NRboYGb8qprVV3rsFZGTjeoh6RK6Q+hTve9oSAttl5caeMWc
11tlZN+zxqG0OzUohyPyeU5bP/6lH5g78XcEVJ+sEwaIvSF+LBLQ4K58ap0RASvB
y4CQ25YEdxivg4Qp/lQxO/L+uzOIF1hhGxNu+G6Ag+qjrnM+XCaRgkJQ3Nf4eoWc
PyslVK1dNmPdtV1Y0LMeUvEwn3Mtl+WhZzFX1NtvoW3gE1SM1BDfzVqIfb/Te9rv
DVWjA5W69gQFBR33pY3TvZ0RrQZAf1bJX2WMJkcH50VToRDdfZWx5yl+EzJirHuh
HJ0hUkX6Fc7py7h93beVXM5IhXb7VTc9NGADMGV5Tc8vPBMykT6bI1Qplytbmjgq
bDWShTdv6DZ86w/LUT+moIab83c9SNWB8OykW6NxQNPN7zWVCl5Aw8FjMWkWoRg9
Bk4wbTqHaGUyObUKI15Get00DymBYXmGaR6fLrlUoBi1uZ0M8uy/5qj6dFApUTyK
FAiI+sEtscZ6Eid4N3DO2jcZcFlmQXPABH20C8F3jLIlhNKOAmkgUXnP1OInyz04
rDm+27a7TMTh+JwbfTyLQFjep4Xk776rr9cLGiOBJzTSrIZ7mPq0BoHBivHF8qB8
5+Wlmdb+GBlfvaWZYLGtAdeYuu5rJlmk+wUXQgj1nxj+CY6eij8Mc+MLwugAMID0
Dy1QVXA4IFTKKUAh+1dLweuhOX+uVYh/CWiQTur4jI1PFYX69pQ/4AJElVOcAvRy
preIDwLV/TZ++o0abNeynZYHC4tdsSyEJYjF5PtBvoUReVuk4xeniFsB0m5ySF8a
2IfogPyYTe+7H0IL5n0A2CHuk1JFPc93heJLTLXQnVKE83jFPxofNOObJAvPmnzm
aa9ry7Aj2zXuRNJMhBFlZT0w6EarNUEy24f+R1Pu9b18SKGoxnF7CylGp2YjCsxA
9/NKvrjWQalJxG/VeHb5xbvmz7h/Sk8kM5Yx3+a/Is28Uo3rl1s2m/iY2/3CC/MV
o6epWps0iHRjo3IKrBMO1ZdT1tgWlpLoTkK299ezJesb/8y/ZASyAa7Bz8UCQS2A
o/ZRV5qVMJNeRBTO2G3bFwg0G4XZXak3rO0en1YtaBZOLthPhkKUHpl+yNa5oZwH
xpYoKGZNpv6BzAPu0gzKV2ILo7j8WZMXwIpTAvsXN4dGPDj1a/F+a7tBOyjILNOS
XeXYWqcDtrLH+MbQPRCFXOsezRxMR2W9y4XqrP+8slC+j3vsjvQZW05u2Gqb8+kk
YRQFgHyhR3k+IxnBNATgsAxXMojhJlXsUzeLjEi9UeB6TGgWbZbp2hzfdNuP2tYj
IkK++V0qIgy++cg0qb16wxXDmVvkL3Zj4I8hyqsOuKZuBv9J6hqL5XOBly+CpjGC
+uy11ePPCfk63YoChb8AhniS0vVG+i8pGtgwkLeEPabA1JHmjAUqlykhYwPES/a1
6LDUQGlfIcjlP5+xRA2TBjbRfr3/c+0BRSYnVWQhyoc2RJRmhCL4/aNulOsuJ5+g
i0ByVKne9ToCnxYNdJJfXs542YGYM6CIP6kE+CFky2fGVMio5VfRYhIBsz6uZ11F
//bGbKFsbWYCBDjVsXNEnH/al/RfdtA1vuA61OyGSWmHWqkKmc0GTIQce6hA+q85
c7MeODXaZp1Ph1QJm4TIt4yxC3Ycx9Uaf1kw8r/tWCACvbN02omgFeqxJIfIP4b+
Bxo+yQNnxjpNIvzdzNO2mcxnkc2wLV/amTV9+JF8yBg5/0PPEpbUVS1fMid48nsx
JjYGtB+atZFwCoWs6xGmNwfzzBzWMOgvTBqgJYAYoBIttXnlGPUi0zINcJAsK+29
cY0CFLepGAqw6F7gtcdEpBGWT5rq42Wbp6lRYq4PYhtBsiVgd6C7hLe9jwd+cURO
CQMhXXwhc/AvV0TuOgfn4ouaG0yj4meaqrCQmdq8bCvnrJ2hC9hdXdHzZZfaCTh3
D1Dd2hNkR4XmXLzaPyuxCrXW5gUuf5lob46mUYj5KyqXmZNulEvzdxa8mNOcArmY
Joug7i7BgWyIg1+fH5lWGlyd70VUkGHc80Vu1x13EB3ouvWH3uJprPDxzGm9Psmn
w/c5u0Rt2z1PVBJaS3xSxeGIbQ3fjf/subG0qsdzUbvHszhnX5FLC6W7Nr2+OOhO
pcZtdxcxmTHNoqEwvC1xeXkmmw2Mqq5yG0VzUlsRbfCKhYnpLiKiDZzO1sTvcAog
qXFUTgodrb4GEmW4MHr84tBeHkWLShE7sUgxvl4H647qnzkGrtZ/IbboDmaf/oj3
Zx3XrqmhkOdcSt9tUdAWOimtk3gpAFmIMqF+ujJAx5bIQen9a+DMB46PMATbz/CD
PspxSnoaN3YCSKjviJtB8pY/UQ7iH0YNrwyeSjWRYbra9KsgwlAfSaUUUY+9g+sJ
vwx8vuq40gaB5tK1ctrV8pyab64CjTsGahw38CSPB1twlnuDliH5sW0k6Mb3GNAT
tcajnoQfwbEXp1LdUC8cHQhUQ+XnGDBPiVcBgTICw/8lGR3aN7YQ99YbKWFc6Mgj
9u3HUeD0yBVIoSiF/5V6Wa1WX66aF3JF+9ocoSrhVK+4/wgf76SsB62M8/tiIepN
A/TGaN/ZMhA+QOAKo0wuBcodaL4cHLez9nMhD5abLzYbfQ0J4rdx909EyF2fbOcj
NP4xyldXkVEqmma/mkwFt1uCRO1B0xR/YkL3sEq67BA3XUb6mBEwRofq8qw2LXya
PpZ7YNNvu8yeIbd0Rubdzgm1RD8nb6PyyOrOgLZaGZBHCRMYve3srNM/+Yw1FQ33
xHYQycY0Am66YG5282h6Bx758sBjP7gtccfub2u0861BnPC2z9e0rOqSqq076Ten
R4B8I39IwgsbwjZE1llNVmecbpYNKmlTgJzh1oNZuW9grcuj4M1tQexzu1kaGVrR
ZAbdF8BGow0ZI19GlrsMcke4RSvzenX18pqp+nxjcUD4PHWgzG9espfUg1JNXGy0
7y1UsFWVvoPP/67VNDIIkdGzRmCxRWswsghO0DcLMBqxlF+Vh262OSUfPpj2CSIE
YPztjBpcvkaOIwranbElvhwehW3e61H7Cs5UgRxvE5kBuqGcBuNsIsa/KwrYji0M
7SPh+g5XidwaYLPJbz6rJtsB7U/9nTzp/WFkhgcKLcGPkKg+mlByUuAcKEsQrlze
h+PHvEEFbU7eUFMalubG4YcoWqnZAclS8QSYyQdS8y93b8iV6bEmvtH/pzhHvNEb
awdBkdi5jRDbqUmhz65qzCzEUrEKn1Z7QaXTX9lW+rh71ehH7suqScfxNKbda/35
MGIkQ59D04S2a0rquLiupCn1/bApJo71Qey+I3jc8GNhSw2DBl+gu4mcjBCRnCxA
Ryhpzud/goLo+qcJ1SkDzbLJCqwzGKf03qRUD1VqQfXCNNyjfdjFwMqbqw6TbnqH
/YXyAjjWyQopDGFK2fJcowlM/NZoq2o5preoDF4BEDo4rZBaP7R9lyOiszWt0UhU
1TjcECtRZZdBl/ePTbGYR9qUckHcdxOv/5TVdBujGe2E1Sv9/GeOzLhT9tj8B4xL
Lzr6KNsKx2p6FHnoc7shr2VuOjGMhMkA5dEj8KKWuuVdmlBGXVye7Uf19gVV8lxW
ugm3jnlcb4MagRl6yDom3EyrsBukMOxF6qTsO+cTu/SsEjDJco/QDd/KwhyIg1/t
WjsRMAO0ngib+ZWz0vx4nt/h/hDOaeC6/6ohSeIXYwYrHhBSHTBZM3nqFesEM87D
DRahL0ssKwrdDrdCA+exXcPDBYU+2R/1m0P14+y9mwgeluhYrl7CUusdpADdr8wD
igRaFm5BzYRZDcGVs1RkgM1qk0MSTz6mTejQ9dDxuO+VwIjqaoJa1MlD5ebqNdcO
D1xfp0MXADMjITyP7k3eGL05JHANem7TW5AJDTnq31OzqtuanfhfRFrYtjLYCqlg
WBAPzOrJT4ncdtmz/b0fT4zaXG6YHUwINeZ5Hb0CxCIFOmenTROUHqm+zc5q05rE
Y7J7RCyepclkO9hI8iSihKRYxzhi0rQiuCg0bj+8oKwVkdS0PxQMXrnMsS1/IZwn
IbrZI84bbANxEiK41mhF8tUH12VcAlVFtsjBv5o5+eePBkyiQWn0pXU2td8+iLR0
mI9a/jjwyFAKXEbOquOhMH4Cbkl4hl0ARVxfQVwT8gmGWzX5SEJff+AYLbzfTwRC
JX1hmaiIEdkoXdnGlQ3JBpk4xqZLQj21Jq9cerN17XxB5aZEvcVolkKfY/Voq29q
A+0rjCNEayR389QwAbDWgvgCT3nHFueFFKdT/lGdwpHYRPlSoI4K7X+C3F7CHVtg
yx2W+eddRH+zvsCUbPEiZEEr1JKdLfI066ULIpewYKsZPj0f37R12fe7FWttgr+t
cUlIJSiDMEp41H9NiIYE/oow/ZELYEGPv3VH7EUr/O0h2UaqFwDxm+jMNdOlOW93
e7Bwv4m0MhuQhQKhVdOy6eXsdYm7zIyOlauSAWJvQE5NmRVLF6I6WnO1s3VG80B9
C/5Vc8r5rCxCxxUagNFd2hnNduIatVBknsXy3lbLRzc1yfF0oBN0nrvQ4QPLJP9o
gZSM3d+osSTGlyc4O3QrvtasMgRThLB/lesOBpvwy4Wpu3S4h3g0oPLPPXKClb81
XIwJ16LXyyfuZ1WdzqySclK0Y5WaeHQ0YoZeYNjyIoYAoxXZOkYEhwpHnUmGmwsr
pqp0gXP/l3NHaZuDfkv0WPXIP89YU6L/qYyvLee6ZX1G3pegjzFQKqbpLzz/qa37
4fvoqNxxkXx1RwEYclt2RpArZ+xvyLLPq24/X32V+vPmuRiaBMRgM8xt4hYFzB+q
aTHR/aMkj2F9CzUvUFztNJFV0gyuR5kzruNezkiXrTlve5nuXQwe2NP7yBriP8wG
lhMVRiDszj0tLcAAmy0UUe/8qPu8nZ/l0jzL9xhxeZ9NZkWXdscZb+U6fR57JtGZ
VQYXUjILkDLdTqKfpFDGOlMe+HZIqZxXAGGpjvzDKMARSDPVz4ymE+YYyz/9IIu7
DMVJ/y5jILyOWgXF4aDQHFwHxd2V3e8hqNfMa/vLc2sP7lwY7lTo3WK9tp75ptVJ
EbhFTczFUw6SjE61sq6Civc1MoCZ8bctZBedz/5vGh8arEk/UB8BUTTA7D2khq0X
/WYOucjGkY8OheMleP2QdGhnVcKqDDWG/Eyvbd2gc0RjPa5lsnA32wtOQAGVYSoB
TTtDOcskG4w9CMR9rc8PJDPXZDFxrRfzrZtJ5dSQqkP1cKQ7dSzg8YPWlSLtSk0P
j1+mnQkz1i1cUzVzCbnZ7lYEZsuanbaMjc9+5z1AO2qoE1Ck1YJz/DZMStGHYIlh
xMRygvdybDgWn41kLW+5OsAFdYeuSCMJKTYDzF2duPRgUoRQn6E6onL+bUX1N6T6
82hnhXnff+13N7RaFfmt2F9voqxAGz/UlpCDN+N6DvwCEMWHMd2ARnUyP7Fs6MpS
LAE9wW5PffOc8+i5WDzZa9X0oesQBD1gw/G3picuIYJ5u5ajURILyZk0UAsM8pO2
uOG9y7NhPNeWjOIrkSIVzg5FS6ZOPfZzxWX2zGebFES2BfI/QcyENgLIqNF3nHmG
F+2hs7OJ1M1rj99oDl+7bK6SYsLRhl4TC4dUHeRkCL5FfxvRERbyvfY1FV9+wdOZ
udUNleUsuS5kcC7qpgTDQ5/wZmkVEWkWKRmGrUthmzbzh4Tkhh8GTgdKnlIGcGP4
vX+lLrZnWNRGFTtGkpXBwWz/K4PTVhqIteorzuTB0UYEyRuUdWGkBqCAaqwAC1IC
A4zXGukUAL2ZQ2b6S01nMMXjJpwaPP2wj0OdUoeUeOP/Fi6HYT0/FEDZll0U8V7+
Nw9KwCNmrZu2VdgoLxBjZYvgTu9NrSto8eJaqe3D6e1TWmx3i7Z2VMD1SzHix8nQ
wqGBYuohsNvA613dnshAR7f9qNE+McXstFAtzjyLKuq/2fMUnB4Eb+97dmYHgnP8
vHL6oXIkw0U+KSC+IPC9HrB6hu8pDQ3ojOZTlOqcFlTxRl/TKkCx350wgbQCmM2p
wFdWyFL1wgw6/pE7WjPK2uRJZ3hJwzd2/ttS/jrTvdGEX5H/jWUGpLjCAq+Xdv5v
99ksWU3kZZ4YZrdw2wyoBkkMBa1lfs/ivMW++hmxWWEw2+s+UY32zD376tZYK3b/
2JAhdnxyARTrkMpsuhC+14+B9wjvoSuIkhrSshpJXQ1NvpX3+JQ/o103mWk3++V1
e1KGLox7AWKaGUI1n7UEs3PlAKRukRgPx86aTal047Vw1Cmfu1HbmSGhAc6tyGKI
o5+bSRLPLIG5hPEQ3FgdLjB20UNq8lsIqwLD0N4y2pBzrfx1Lgs4nc4pzfaQMuBG
tPCNgOTvGLrbryYp573IxpzP+9Ewwq2No86TaK63Xxs4yPUEC28RfbAsGFwYTcQY
AH1zsYV4iqzQgdFmVSyjrnVVYO3mbWSV/LAsuHpeKSfkZyu8/hy6nEN59nR1sGFS
9BiwlVvJKKdeqIuA92+4uqGezRINp9zC8ljw2x0sc6RJOt3IhcdFVg2PEdO1uxJT
0RCLrWmhblqLqv2PiyTChirqAJPNT0FfHBgWL0xQm46FR537LkdkyvY95dmYEsJX
CecRqbf96wRZUWBtNe/e3Jj5i2uH7G540VhD6ASTZtsbZ9tDrqIoDiM7of9s/lYx
dmMJwe/rldWlZa86xytoy+jN2TeX8mAPCLpaHt8gAt8EooPeEir0lyq8XOyWnKkv
8x8UWmCpD1RQDcCuTyCLMhbDqdByOqiAHTrtYp1VmdLvMA0wQmp6CyKzZcwvthfu
pquEGS+KQrqldm6/icQ/TEp1r/lGlG6BOwflqTj9e72HfgLRz05jfOm+znGFv3P7
VO0c0QWKXQB6srKu4xjZP902B2U3HhdNsprbVmCudKhY/lKDcIEvLBX57HMrJQ46
vRaJJxKTOqwpOrnv70KmGXDCUgY63vXfkqdtns2j3o11m3I6tpiC8saEOjCqfuoG
0UU5yR7kAtZ+Bj4lqkaI7J7szoWXWrX96rPewz6D8SJTzQQHb99mJnD8XWZjUosQ
lTqeOg4uiaAnZ6wpde7Cdrrpq0jMQubn08sSHsEyfmgHc49onxsZmLpBHqoil1/K
IhwRaXvB5ofXychWuRPZLhyz/a/8Fn3trXRHaCEPiap+F854l/SncVBriZm9ULl3
oCy8eccgsQUMtw8a8yC2312Exn3vSm38R5vLywNtVWtHpHFji8H4anvi+HKKS+bU
W1PBop44cfkfUYVX3WxN6mzCi6cOIW+meCPCDuZ+BxQ+ohc65P2d/U3LMENH+/Hp
jUwZ6oeiBIzI+hgwvOn5ajy7nrv/gPW5MvabpKZUbT8kvxwLJ46WdLGjboLVF5hR
ArwhDM+nCRYYXC/09i0YnF1I5HXzwfrk3GJbULr3JrRKNN2jCFUcs7tAynuhd9P9
0mjds2sA5BjdsDTn5ohlKK2yq4VR4jAaP+Wdeu78JBgvW766po0F1SJRyKiq25tw
eJVHb1EPs5X54RBhmLZSUI+g5h8UY+JMg/98FJ8S3beH1dRdbuIVj4GZlsXhzy+9
VCUHoJHRVROpvclvCYVQshthpV1qbzVj51zLzU98JSPj6Kbw0ah/VctW39st4JKd
CdftIVVsCHpBXeFTOj0Rd0upJVud8PkGlQcU7E1XbZ+DKnSwxVXwUup4z9xDeBlk
O9kxbN94J0pqI8srPpNhqmmfDQy8PpasBL0KMYzNkEZPgRJQnaR8zBsouxZZL/kR
UEzJwdjGkCDdiH//VTpzfF3B57fZAPRUY1ZC3fN6+m0g1fPSngCyjCmtI0va/n3X
qTbBnh03O3bpZ7URX++BF51X5xlYb5mSGixkhnuXlO5zouumU7s6UMjHgZAnhjhk
1GBqvdTgwN98VzT4MnXvBwMYdMCt5hskge9hMAK1530aUQ6DlmBQe6B7EEPSyrxj
vw1gu6JZsqM87jO9s919KGoLY4JS5hYXueWlY2/we+wCHS8YcYGhcnoQD3ffiIOZ
42kE56Q85oxLdAnWw06yMXPQYeZarwVCKwgHx/87txim3J4URU2CSjDOuJoe1i1M
whRwXujdHVTPTDU6KI+wzX+ijQz+8Nqitv9LVRDSuPvB9YTR2W/PZSL6TSgosTD0
gxp2VH2Uf285jP3GEvxWio98ZZ2whjqN2ukTwRx7lO9nCmZHI+3lA9jQ35K/tixx
9iE6SYl8yC4sAwG93bKHH4pbMhnTwpS7K8g4VcQPNHXo+eP6wKSBL6opxbOfsLAp
VpRcw28fG6zghVcH+9yNcOWDm+u9pF+vRBzcSkAnq3YO3KDDZPPimZtugJQerZWr
+98MzLFKVJx3yQXVmqU3khtILDAuESate33/F9mHR9vD2n6Sx80TW8C/9vQ45nck
TgjCaEGuQvCNyErc3wyAA5Bg6SP4GNK9uUM8ghQQ4b0KYifm5fAUxDG+4z2joGXf
2YVmZ4TdhwvxeCKL+rT4r8vZXCAPCCQwA6ioGErj1jVgrhKnoffdHLP7QBtvTjEn
7kAUDnw6DWEBrsuBH43phMZCPp6DzEFNvqIirpNVSpuXjzghMv9IXmey4DUpMX2g
YHM9/AUqQmmGzmOsuztETsCX9JVuyn/cd5HPh3j7iGIOd+XrMNYkJmNAx2tS5P9D
YGCePEq9ePkI6hauXAvt47XTWLgx5PCuOYSz9fu4KPfQAecDV1qtWpx0843nUgyU
13LOudJkQdlLJ7yU0yq47yFL0i8d1qR8z5Uzmt9+8t175x0lzI3k5rnEapu/ezJP
YUOHTEmmtousInXv/oEZREUT6rxrJHJe2h3a50q4Kto5+7BmPWLl5EkchNNOLSXX
dKbjyz4vlXvEWlWRDMJl1IJCFeWDHA6W3rFsmv0ztEoAqbXprP9Ip19R2ZPfn8dh
0AgcBz6cIrse7bkGIiI3ElTNpqWNUiNqYBrzNEgdesSAuULFl0cwZugZdF7qJPWK
GYzgDFkNZvYFOgpYLSO2x90+XNA/McCOo4YaI3vEFXga/WZ1+Lyc3ONopSeIo5vb
THgTnmsPOEnTNWWsz4LnRNpRkV7vexwnij7IJCNADQ3sHLqXeum2rxOPl6CiZcQa
k4OuoFQF/J6xUfwd5M2jaOJi5A2rfjpPNqCK75E6JS/FEOKH4ze74lIfF/tiBHwV
iZmmqZXbIRZ6JqwcFTE2ylm01ZnC9PQEtUC3rKeiBxCtZuMXu6a5R7aQYAO/5TWW
Bm8Y0o3L36E+RPocoh0X/PUrNGcmcnglWKN17i9zZA5QGZJRamgrLFa+XUBXHrdq
EokjkcqbbFV9V+eGgqw8NtyAWTq/fJJNWYx6Pk+c72pVmPdSWHkpUqtAK4d2DtZ0
WpxIxPI9r8VTmFdsPliA4qQq1wvmjGVTWVcjgLUyGY94Nls2fuw8qhDWkEcfmP8c
Fs/zUlM6+wexR/6yCL0oPZEi5cho/uvOuJZGMOeL4Hc59p6R4Q6eLzCPcInULK3e
X3Q4VDVB9xhwb3w8MDzXDIzUB86XTGgwHtMzJC8d0dsJ6ktSDX52z3x0o6Iu+ECh
wgYzjRfhYBfoMtlQlPbHGgqHSuhYihFVp4Y0Q8+Eret4q0q4WJOLULQ+Bh9c9QlC
fSCJxVrZknsMRzwLJ0mzSH1df/nIyJTlhl1IukO6w5MW1f0cgJRxsp3cj4Bx74hq
GtMVmdoF3R+xRZnNHAjSPz9vqsH8OMpDLVw/JcJb54K3DVr5u+LW4EqTjXqTODkn
r+CoGb71wbKJf8BnF4FUB96YfqHe6Jf+P/lC4K4wdiemxa65uW5tn5u8f7fA2U6w
Z1zbZlgPZ4M8cbGhpmmC0+CPVdBuPIufZ+VPFipv3CAWqJtI5cFbuTLill7SW1jH
Rkq3jfwAFY3fdLSlZ7448eQbuHhKN6xZ/cJ+lHnGX0UfW+MVyqi4SpquwCcma4HW
6NY03M2sH7HorOyO02BGsV2IG+A6fknkLec9L3rUKt1JftAbnDi7pNZVkfPYSNrt
PoYo55eE5p6mqUU6jh/fsbjrwITPmZo6jM/m+kaVF/K9UdaGdXQ7t8gfQ30XlC0f
N4uU2GqiulroBgT1ZZONBMBci9zlhIOQYFj1VMYkY7z983zHwxrFUq8GOp6qhasF
qlSsi4YPPLO7HDBNda2CRreSMfyisMPzYGslZxtRBhZSZ0r9iEjhKQguZHydxV8W
A+rGsKG5p4wNJEi5gkhnraeMhrG25rqXKTDVinHwSVquL3oVz4HbJxEjEspCzpzT
fehhQjpP6M+GgSAyUZnXzQQXvDz7dAzIKIDRqXv89w9P96hG4aLLcejXd1SABaT0
7L+Gc+tWOcAM6HlZYT8mHUCFJNp3qoiKKnpQxA0Z2lM0WBjvJNbyHDTWgUCSGu2M
tez28+pcy/zIexascxEq6HgRFJlmubr9xqRm+bqp6BufHjNTi5AS7Ja4nGgjbzLK
E6nD8ooE7W1TXz2GjspUDWcyBTs3m/Y9gOmBL7JcLbE3tXuIbOYQ0R5pHZ9mfI1q
7/ABnuqKjjn0h3hENZO7aNMEz5KyVfMmr5eiC04wTcOIa56BPMrJSzTk2m50B4/Q
QmHI8Ov41bnXlEkp3nUKxVAh6t2/VRswXpN/ffdjo/dooYD55UYOGioML/JTuFaP
c9vvJm68gD1oeugDHPiph3gkjPbPIgUmbnotYEvtl3mZ9G6nObAFDBu2UohLEb+I
sk2iHY3YSnrAk+YzjAHqYqtbL/IvRgDiI8mWj7kSEKUbs9LcHNyyi9s2vHJxpz7F
AUdow7s0Nx/WmIg1xW76xE+2kKppBCpxsEkdq01iNlWGNyAGEyzhTzI1Oqq5f2f/
v4Umx6BJ4PrYDGw72g9xGd/u88P+lNPmwwj/LTAJfVYt+st0Jv1rug614Iu3dydA
zkDhjwnBCBNJyfBhrd6ilZqS4BjVctOWA/58lGc3aNbS73plW4Zt9xjDFR+knBkY
p/cMin/eHqbVS28HhatSBQ0q5MnQaShQgOvFLophJKXAq5C+louuAxa+i9lyBzKz
GhzQ17F7wfQP0apSu0fQxq/r9nIQsQZFXBDpZMYiY+tRjs8wWcGuLNbO+LEgQyUU
pnYzpswVTpjguc1wIfZPA0R0ioTkR/yWcErZMzdszM3XvnKXAT7EXTCxjs38hqe/
8n8SZrAvuINTxJuAGiQzYgIa5ldSJp5gWwmnv3QV8QvnIHxPA19AOuVIlKpZp/E+
By0veM4Hs98CmTIAkPUQ03o2gp0FVl5YqrN11JxKmQBQc1xOQshCyH4Pk3orMtPH
4rq21nV1hAZ6lQFX/lren2s+XcSIcPbIcWHpk4Rt4zDKHlVO3e6lWVUWnj5F/LiZ
rT4iSxd8F99KHAZaA6TaukXbJmAevVSCCrYqA2LSdcdQLGn3MTeTTByYM9wvHtV/
SADTmkP+RvWCZhhkEV9KpP5R2JJpTJpOiMVTifi7cG6xCN5/sNiWj2fU4uWTFBo3
XgoH/qinwDsvWSFcYCaRZoaSV3wVyMU7rF1j1VzBjx/MZGmbLbwD0gCGHauZVnJN
MBDGiBp5PV4B0c67sMsDkqddOSSjWTJ308vn83uK0lXeligcEajxI+PeU2gsJNM9
p//rmcotH/GsZ9mFQJPSvRK/DqTKUNWY4qFKbSoFGEv2F5A1eOLocnPXYa3vaK/O
AZIgyhU2CHlucv2hjGwwMLu/sDwcqELPFoJYbgstz+DyRpkHwbW2ZQLVKZ03M4mh
p5I+CkK+OHm6jZTTC2qbA5CsxTBrKqpUTQZJcPl5k46KKEP/D7+oD5CgwQ3TN/XM
b8qqNqR62PMVrF9QHVEDz1Em98av3YMFQBfDr7BBwErvqZgxD4ZTc1pAPzo+UbMI
NjpHU0PrUFmPeGuNJWfYvxv7d4eQMzxGzsBMFeZ+o/Gc+Y8xMBWyrbQ48Pgf02OB
1hrYAM4xcwq6k0l6tijYlCybIT5ihRX3xzR2uy69wXUVfkovQzv0mBQLkvro+3Xw
ax3XDhn4zWSU931L8zN3wEdyKNAEzvXMhcX1K7qkWumsehF0vNTORuLHB/pzXrLL
4rZ8+VpWdA7zaWJBxU67eAkJl70z+aDkXEGQSCrP5qkWt91Z2aIt737yEcloEMkU
ELKEtD7+0JEbvOvEL3Wk6C4wA6bBllkw/FHOYN+4E/NZlUpJ/trd8Q5YgxdFGznz
/6/hAlagfFg/jYAC7nHVU7ngQr9xRXX6AlAsoNfV0A/ZdIUO+Bxpu3anMXuTqcCo
s+4Lxgd2eJyZxQDgwb/ut9ZRu9HaYbkrm8+JLGJ+6e2b0WsT/qjJVvZ/sb+gWfRW
JqnLOROaA2BtA6ETZaeXYH/8gapK4kSGmHGzWvlO6kXqWzvc6R+yRhDnRwUd/GO3
rknk9cclCdyoBMfHlQcp2ZTCAStqabJjulvAqcMBjbE7j0LJm3gRQOg7ip7DOAL9
SR6ccXys4Jtag87MqPUBTDJo/flObJ0kKV5PX03KoU6Uo4zt51YtlyNUiStEXHAJ
LQTPE31qWThtgofxj+3SUeY2JriYi/TLOS30yXgm5xQNFBejIrgrOOX71EoU30ow
a2dvH4WI1bZwBqZVfOKxv+tcjQ2eJv4FpeAIzZbjZZZ2EQwO2q2HUOSEoAleIH1B
AxBgaTB1nC9ue2haZI/fsk7kODg6n78drC35kvNC4wps6e4rAIREvAGrg1ln96Rf
d1R4VhllZyo0zLq/PsvTdY+/07hmqJF5ugEVTXCmG0B/c0GYdiq1FpFZ+egY0Kj1
Kg4RReG9uxRrZbFyWxvXcgxOR4WiLmO1iUZGwNBD5NGcGfnxGGBYdaweYNYTUWI8
J+SD7SOmvjZKDwPyXly8E9YmE7jxiMzm4O8/4lN/zwAQHYXWmh6/vkpVEpwi20EW
XtN93dcklNU8ZKxVkcmn7ErYsIf9L2xs0BxoObsrBWDdHAQhTUMXeB99QevDjDP0
y9zCgUc+mDJBWPrH4PLBOqjA0NigEvJVvc2r1Laa3DGyFbA/aaxsiUiH9XwZKKZz
/FKWqLdAsVChN5n05oY9KnMTH9i57q8Qn4sz9p8pj1npLAg5TqX9aNhk9bLcbKG3
+Bqc45ZMESupMpLV7vCbk2v0SiOT0rjO6f8QcOquK9FZCsNlokLC0tQrGQ+rUv2Z
UQgdDgkb4x0DK9EtwAaf5dmla9cA9/RNh2X5aHFNYCt6tMeY+ckO92ecgmyIWKr6
rAv20cQ6jqP9OkqySih9FmN0LWBwfYj/vPw8jFUqGVN0AP1/78TCvaIfGzLSCwaB
zJhRCFLtgb1i6njjEgF+LE0I2alMKQIuNooD+2m8pDQUj6zCcCnxy8AAYQNdpS2/
QXjfNLjAdu0uzXvhWe5blI5GTi6PMEyXqmb2HMH4CW4esmkSDSmRJgm+YnaN72Xh
iErmFanvI7E/KwVog3a+fatzQ1qd6KzN2tlaMLXwfdUP3rjCIfxn5VGiaPs2rPiX
an8hcq1V5Jm45U7L5lD5mvCw6F5KsZFDRJqhGMIBg2NrIhTHp7R7ko5ipOlPBLKT
jog8WqYDnzcKxHNyxTbX8lVzRhiYjzZK0gbqHTtyDPweCJ50WNIrnqkHIgHFfQv3
alEvixgNdk9ntfrtxtYx/SVGuvQAD/P/kkONpehkl+JPrSj6Y9MGsxAWwIIUU1Tx
Fj2sfGFwA5eOU+o5ArqVgGJQPu5TeJ3sciMMKe3jf9oMUT9BQxtspKYkhIQ1xWeb
Lyf3QwyB+i5+yHVGdP2xLhsYSz9OlONjxKBD86c2mfTnaqzY5lLWAaPqjVN3eKuJ
vNxNhKbDxGj5FdWOJeuUmqMnTHfj9g6iilJ3dfD/z6q/22npDFzRr2MrLbF6GSDK
B8OxpsLcktPsLyizZT0LENQRYsSb+9mSgdPZDcsLtIEcC2L2kEvZ3dypVFzMkFu2
PB1GQAgW+WRbEk2pJee8gfrWkWd68YJ0HMluPaq1onD/aLEaC1KigG4xZOAv5IXb
jjznKNyT0RR/9aGjMguIPp7r2ptyv+vtzHN+6LAGvMfbK/8qGSRHk+OOmtQphpEG
/Z/pKbROS7v2rqQN6pm7/zMq8UWBwsXRRWIyoWKSPUL/5HxBlgr9UjtyBEmznTlf
cyeoBt8qHY/3olYA69LNqo3foo7d84b74gIlYr7kk+irOyo1V30n/EEuhMeIeF+o
lQ/jprrpMLPR7V3YVEBsvvQYrn7RSXOvT3qgSJIXITpmzXX8kWBBoVAcSztap++j
RYZN1NHB57EDNsdE+8O/P39gBe0Ge9/SPtl6DiuoT61+o7M1aqf7YFcDSjqGv2Go
T+nv2wAmMqy+FXLvLSxugro9ZPeH6ZWVb75WqMnvzwOKsou6BWNZhTPLjyHpVkyA
hbibIHtFFjz3aBhgSULvd5nYeQeNnSKxsJAkOOM+jgTw5O6txyn1RUcVw9xhh4+x
JP8eMtnzfWf3qPhWCqF+TzVPhDMvdKTCAD3cqTPd7rfbfasQP4JHSuCuTtcvq8BT
foNK3HDL+LxNU19qLjAjK68vTc0aNzMOuhfrU03Y7r2zpVhbu32G5RWVYf9JjaqN
3/9Llv+iBzMXJxbH1htQ2uBHCJf2Crm8WUvcIpArcjLrzzeE1UmcFOEjl3rN4GUk
GWmwY3SRFDft0kx/2fj68R6U1Fd/tmEdrIaItkpThurR8wyXJ+5vbn6w3zSCF72e
uGf3IGB+XZZt2P9QNxjknvJ3DqG1SmXOa/9qoAXvPMruI+S691ORmihRjp79aRIb
T01/PofCjRkKsBQ5EB2m1bsaujbv5pVsUAACOAk5NUnRxCiFAs71aLmFCWWkXJwl
uE5Bn4nkKvBJBFMMBe4Wg2BmOJSS4XQmFX5BsTc8ObyBPc4c0jbp3Q4scRAz0JQz
mOsERCIMM94SPTh0zSUn1MeANZp17iyfwD7a9qPFRqtqQNPZYXSGEDGs5JYZojB9
9mIb/bNvuWWw8jI1PWi/Cbi16K0ZWiIs3ec4PDW9DhbOxs/gPg/hoNm33qDF8Fj3
ahUVDp6gy1e0+LGvsyl//h9q1PPcd7GW2MrLvHRjXj6gUmSfhc44FW6TJegSdRN6
APtJNLf2nATAm+95ONQalXEJhEHhrf0pkiiuxHlGYpHVxTsb6vpiVdFaM1E7Pbeg
j9zgYhCdPVD4Ynyf/3tJ5LcnodrA8hA1gW0+wtYmm+BIUBw0rS9LyzjENucWwa5i
SnlKGYd59g6BM3w7D7Cex01KLL47q2ZHYJAITrSMmJVIQfIyfFs8EUUmXLzOkanO
FgGt2CD9AptJxlqD0kyNH9ub/3SrzDtLT9krGIendgAEZe2IVFUUKqO7R358frn7
fyFoIZmRn8Bz6YKYPIcUFwSYKKvF3x7V5fNJUBFP0LoH30z/Jtv53St5K60jjnbp
ygjSVKn4jkrHV8VKVbxdvkFFxUG+xYC36dCRRW5IgDUhegbZzXmMIEQZ+yPo40sa
FnIL+8rAiZ9JK0pIlitWPRw6bBAigh+t8PTbg6FFuZ9ScdhWeVQIvoPo14DNa45h
RKxKlBR6D1VwtGbQW5Q7RKnsYRAItxIWrfebSrV/JvL1XtKkDek9M5LTKatrMamr
oTjAs6NIVU3j4rUERLxlfaGqwSZBt/yXLN0u9D8KW7pOWgojx4FEP3BE1bNlPtIS
d0Hk31v1/qYo3KeyrWCDhR6XF7vka5ma5lrIm/+aftQjPnUNj30HuQWs3QG2GO0l
rnGxCly9Kc04fFc31Z9vL3f24ND2HKyLwibXLp9E0QnlnKZTj6vGRTMbm1HcFPwz
NK+SJDnoI6UEQD9F7RKhsJ/Nok6s7oRdjcS4Yk6KZA3vfaHfaJJoIV82hBmf+TFr
IMBWilI2hBoTgO0lsdWJllvXze39K41PlMnqVzXW333Oi5iY/XWPmJ0zSpAjpmYe
QkEXY3rNos1/TGBjPAJ4zQBWJJmzfmyeX2b/84XRVS+/cXr9HAa3sObrpA1M8cac
sM95G1c047RmX2wCsgQJ2cfpjOcY5w1nM1OW8mw31l9lhED40h7fB4m2SoPCo0ID
Tf8cscd/2e2kcELoJI1HZ1X4blsPEUuDmDb3HjqZGVPOn2ppAtp4IRGq4ts5oMHS
V1iJ7DKd1T8pZFjXQqzzGH/OfYaTEKx27mvfLKt7nVD63SdmGgmAg0S1qgHHaRC2
AFBwvvITtOw896qUIZySjUVKyI14s2jubH7MxPlAqQQl8qCAk2Inu4FOGyUnmrqJ
SbPpnCBsbfrOMOWmf6n5z6JMpAadyZ2VmhFQ5uIG3CFWdEGaRooScyZzTlSfIvB3
wjGr5JP5cTuzkQAf0EmgiqwiWJ6CBeyjSLUPTERF2cD9wmWyzHYZKJOdetgRKP9n
fYR31hv9tXbAByoMxImgskxpNrtTbDfkTjg95uvd2eKAGqqDtNTYBfJ3PJliPbVy
xssNDNjbdTlbeFSh6r7j7V8sZwlwqiSCzDPqmimXRq7pd0q+ZsfK7KR5ngri7bqI
/whY00Url+p6zNGFtF8KUlAJ8ZxCEoprVWWHJSfvSnkq3I/IRIzNKG3/m3+A23ED
k0MvmLTgeav1vmSWMIyt9G/As+NuZG6B5S28gf+FAzongBTO4xV5q6jzLbrbSHoI
aXWj6Ya1xQGs6o4B8GijdjrMygcgtWmH9IQkVrbrVf1PfF9a8PMek7zeRIFyfK6o
kAS9VYm4cbPe/gFl8yZofAKVcO6FSnv8cL0Dy7umjsJO3Mvbs7Zr7eexh6HDgf9S
C/cVe7W20lgOdc7RhRkrwva98S7EycjKyOaT2yD8+nCy1P64wc7CGTKdy5o/e0r0
WSGCUElV08h6Y3WP+XnBSXLtP6Or4BO+hvLAokxABBVy9tBgavkOiK00EUlIVh2h
aWsn+S179H28nRZHxJpNGmzIkaeN3SbMzPpOMRGsLKF7VK15jhf1qehymk2avaSj
RJMTGBVI7mNo3TyiZFLlC9ilHEJonhRe1TnA6eVxCoOeVBYgGSTuiuHjSivpyErB
jxOESXxgp4gDLd0zm0qni6p0yziy1lQ1KLk2eBd/sQDNFSzukCgHHm/3iQlwGfyc
WDVVwtJdrEZNrzwGVzFlJUMofxGetna3d+9pAcqOwWy9JE9sHjPfPkYA7anCxQp6
GvVryc/B++D/KpUEVclDqGvcLrB9PH3o9Bk+eHW/kBgTLhoUB7kIaa15uBPi4jIX
iMpIDC6BDuiId3HGvZhPPQzESw8ktQetLTgTIHyevzal11SW6E1hWPtZzr2d6Scw
Ay2cBtYDNZVQyq6Qm/ao5tmVkjXw7WhW2B+Zk+vuLsqMlbizrOEjymcIhetpEmVk
2mpeI8na/UhowqGpRI6FyNBlZC1AAa+dofxciOWi1Q7s1ImwdciYbG4zfSOcygWS
LuqGeY1Mx/o+8EsGSM3K1Z1GfeegQ4JsKfJDBf09oqcgAwGe/2JnGKDyPm1MEu6o
HNe79+nCuryLKqq87n5Zt5GlaTQWy90yrXQGUCcABRCZntKsXezDHC2SD92kQTHg
D2apTbxpHnxQ+ywrqfguZ6Ovx+8lE6HDsOyncrfdLAIw7U8ppcUi0zHfsmS44NZw
H8OJiLOMacQD3SWOnZKwFxPACBypuolsAlGyR3R0V6eAuh7+6uknZ9M5vh8ddyDU
6wdm5JSPnZ43hSRexgnGpMd8J8EcXhTSYc2LQY6Rf2yLZvnjrwTnahizYH5WsXSU
ojgG8eGGb8LcHYc9e8tV7RbhW/wqL2iaCzqbNuq6ZBQbB9aE9u2MHBC0+W0VHoyb
0q2bLirGF/KB8KMQnVB7bsjKMQ6nVKmFouNpomMH359cwYOOPMpNhmwlczsnB0yt
XRoGyW+MMBgI+ui8sTED/fxQWQ7DVJXQzPgcwJSZCYKg7ITrwfNY+KzDznTRbxg4
TdErJJdvAKsFttcEVMGp4fufXYEL/13XDTq/3oAMSrtV0RIXp1D1l4fRQCvgyY5d
Aof4+Xy4RfA74n9JsD0qXNTAvjc1tX40z4RCrJfhP5sGTOGRs+JICrC5cd3gA0tR
Twp/MRMkyBZlKQsnFoT2dqmOeh23LhmdI8seNCWvGNUj+j4W3QByWJm5UUeSjy4u
YaLQWQtxAbLrXp2BIibY9ktz7cBPcg0bmqEtjqPswarfGkYvOVWvBdq1CRvLESJR
dzyBYwQCP/ZXFjEHLiQV4IuxPAwBAIUq1Dm5RTt+8tvDEhPIuy5svD1pDRboqEOf
4UiO+Jl6IVcF44eRbyeWAwzdPFT5z1XqOq3OWcGyJESf2ZUTReX/eQwft8Ki6kMn
pGF+YgPcSGe3lcpIgf7MSApxW9nq9sLk8s2wi1o96xRAilwf8SmBUYkXF0jxceoL
lY/3RXKPkYBmP9CkGwzvyZ1sT1dluD7EsfaPAguwFpECqNrGiZElkCfKRCY0MSr0
wSI600Yv8sQoR343Jt7kTvuKRH6XA8Wb868p6NDnhAWPOxR/gH888yrFMAB0TJCv
I/3rEDcTaOAepjzdJEbxru8xc/Sa/CsIFIbZDf7dBLO7mbhlqtqU09olswFZAGFx
is/iyV7aSlqC82D62/eJbfsD9Olf5MQMyBqqxgWkigCih7NkbtkNrRTOTA38VkQq
iuCvGYM0JkiMRb8DL+mR6mDhdt7gA95zZMhreIeN0Q9hnmK9OJsG5IcvBCoxp8of
dH2pisVO8ElV+wCM3TicCSqYIJKPTuauVPz5wJqqkgVZJakQ416h/FPXXNAR5I46
8jlPLsbdkGJdAZxHd0aD7Ev70EA4jBZerpzcFenBOL6GNwCtlsGyO5UxFBAyqJm0
T+k5CtW1uIleeULD7xLBSUk2xMMR/Sv/qH6rRWxw3NOMCODzKz3skj38zInS657K
IxCPQg1ryEBh1yPjU8TVzZWBFBIu+4etb9CNlGpJyMBGGGYBbgbpKEvzxmY3q3lr
KOQ97IdK5TT3vZE5R1S7v1IgTaqwO9mfqVWmA+w/v/WAM+zRahJhEcKZL1SEfEfo
mas4X7lEY5Iyh0uNx/giHH+vLFmXaNMXI7trLyf7KGwTE1ADwMhIMfvzUdzZrphU
90C7PXtD8QG73rpq/V/3WWOTN4bj52/fSA9zpmKVytQm0Dpaw5PvXmgXu9CRoDWO
VCUCnWQcuYMWfD3KIN/1sBWA+ygjUBzBufkEsrNHU23Pu6tYS1fqkpkFmUv2L8Iz
DpuZb1USmEh3lJV30jjRIAymDcaF9BIKqTJH9E09l2W/xGrHRn+2+Y9Q7nq1Ibs4
E0Lrc1ej1D9kARJZ1lVKSQHha0ClRqLfBxhYPkmt2MnelyOAcB09MLMrkXGp0ezy
AqwNxJk4mgwi8uF9eOD3OBLEO6Ps7Pj5Lw4gqxncpEK+KCTvwPi5qzfuGQuf7QVL
oAcrL/M+ifoXXPE+1X92lLgUIOZkUtrg5vDm9W31cTFM86NlqjBF/vsNctb64IDm
5N6P6ghnf6Bqhrv7C1QtWjaBkLY1t06ThJ2Wg/szp1LXdzn93nVSz9qYmLJwhRft
fL5Ze4SMEM88K0hVyd+3jecD38YE0HzN9aqaPKukuVdcAmrDZumMzsnQMoqURxAg
zy2G+v+HR5neyzTarZxzx+eJULOmxft9MP25BbNpKqiY/WD5kBBAG3FSp/+Gq+at
6bitqKBXTU8SL4TeP70ctUeqe5UvcKWnaVOgM03R3XdNO/kIs9+auczpIhCo0+Oo
Pc+TcMcGWIWmSLYsEpbj89C9hbAnZB02njURyQEzY00KQeBznIt8I7CpvH1Y0SkQ
MoZ5wya/e0/uO3qHofwTbl2nBvoA9iDGwojH8a/fPKixEDlS83/3v3urVRV5Bcxw
glvfW8QF3QaS71OlMJFRWP7pbRSpoaezTtegSszB1ECmPXSdJpUx1T7Yhik7IMCz
DDC/Gsclq/w+JP/gpelN7u/jjYX5SXQLbfgLzR89pPUX4uPjEpKucagsYwRIAkvb
zE+K8PhiTOiK1FBhf5y90w6SO9Z+/Lf770Vkrip5iasj73hHqhSjk4xtjfLeL7J0
nOZ+BdXh5AuPIEgyz4/NBeQqYjm3TCGhC1tj740P0guIrqQbumvf7kk76EBWW1dW
w5u+Uw9ieNEYBCtHCeaEGahpsVRbdiUhj35NGey1AJX+F/3VaR7ekcdJBMe77yrm
QoMYXlAmWVL3aDEwH+C95h6lpQQUjbTgXO8PElvF+VySap/MdAmxt3RasbDdmZ1m
wpw7n6qPM12cD7z4VUy2bIhJbhuy5mI8ujyRiznCPPqg2HxMrPRBlsgOxtVyfHfr
GDEo7L4fFpCOS/5hCQJ7ZoYRLVMcnL0+X8ek9JQM+PZrzUIit6Hoe+1UnD1UZ5tM
mLX+FmZE3DHED2cI5KhCjEeopaIwmWzCHOsKgtbvCs6uLzLfDAeSLd2HhAnhk5Qd
JGou4lQ1GykDpF5plfPUY5rCatafmwoK/M4gKw1n1ZI4k+nD9wydv2/nMdYhhCef
VuW2I6WE8rJtSZGzSR5pwuo1X2fTK5579NcGrubek6KxwwGuNPrxi1OhSLsqsCTA
OyuxOH5OX1FCKBGCF+V4BiUdbsz3MZYh2Gi0Xgy7COnyLuyurejjwszB3L2Z8IgE
VcrlNj/ytUeyl1rqdRx73gUr//CNAyOWqqnhncWs+yrQWWxd404BaVsU6DdxJoSu
2YukKsO1tY3/tiRitAyV3ahHdwgvlQLen+2pzgx5VdcKphXYgWQTzyZ3FZaW2Kad
iz7LqNwT9JBn1xxtm7YThQWN1Re/Ql65stnjMGfpjR8+z1cFnrlMW25apo0vYwl8
5M5efBaDmqfRtNTkpDZMr9tCUJOo42gHQReuG5D1WiQxf7naYe6TzdyaX65C8tPm
EzrQ2cN/EUbArM45NroNFMEoovMgJFByz1ZjnM5rDkGm5P/Q5baRY7+loRiZy9eA
87113v9Dn9hFbDgZW7I+lBqSqaji9bd5GayMshcqCiK70SrFWrB9morsw86zxZj6
Pls5ujTq6zi73h+CmSDnx+6GLeCphyb1Cq7SHwkKDBNELi83PrcvZuV7G/hLq/0T
zVZYbsrd4l6x8Y61wGuXqCjr7punCMZVywC7U9+6U6b59oO6X6UnSHPpl84r1ECJ
OiDar8Mopa+vgWal3sG/sr4P5+Ht3Yzc8/x/yJwSHosUOL2PquxZevhScb+5Pd4k
f5tsgpeBJT1lgl8kS4heFXmQoZRYKmIMYkDD+smbutkiqLIB9n/5cN8v9qCYVXph
RmjWf1Sqbadl62Hxlmbk4xHT1cQnoc/dlE/wjFq1t6j5Wf8KzdK4v28iFY6PcejQ
yT7zb66oP3Dt2/MlHt22LZD8PaNLur1tn56ELVFiqeNm+NDB8YCMgJ6USdNi9/sa
nkjwOH9lzSRHEOaE9sYIrlOIGQKzS7wTJVHmqxXNrk0sLMpMvNYJsAPQgtOsuXqT
KtvhlEtIBGvRLhHCXQJcpw1zxUtqTJlRhCu8WWskIMGarbiQSol3XKqIgN7Q7F8s
3q5H9MzmRPHFqK2NFIHbbfKjftbUM3wvnyaRg3vOEbBhicF8vyMM2g9TZqk5Vwjg
IEfM+ekeU4R7qXn8HSWF68xESYlORwjUekqwWyk1zC4cghX8Y/ZNVycYgOmFvqz8
D00mWawMTa3B90N7jNbCvbcDN6UziLvnKTwGNa60Tof5zi3p6rjv2a9ViAQH/IK1
VzNZIvanU6sVdO2nrW+9iCNNQLRdtU1oTHls+GxXm6dIr6KXjSuVDhovV+sv1eaX
VSdpX6rlNuZe2l6OyWP6IOKjxn4AccWKlt9MQZ8UQ8KY/VkIT3hxw8O1wh6YjHzw
olUBKy3h6pfmmZZT70R0vHgGhFdXjJ0Hx5wXrmlMCMaYG+01jP7CiGYRHhpZnDpi
fsBdfL/rKqfGnPypTSn0e04T7aYg0UIXVvb7hqTfH39j8jUq8Hn0CeZITEH5hTLT
Izm6Y3Ak+zb6sBVlFs5kv8wG9BKS9SMymqoFKb0GlP97rkQ7rGyIXvqmW8+UtLvT
V1IUzYSqLzDFUI0D2BW3A02FA1kh097GbotrAw18cQdyeAoCtvf3mptsHlJx/eZ0
0BJI0BZke8P47j2VKhgwa6au5zmx/vflVHzXGjtv8/wkTUBe9b+7MEE4+nOpuRmU
0kHDciLVdQismLAqlXvGC03OsdXZDjoQ2ogdQxJ9mIyUDL33yrQuT6trjDY7gGIs
gtHQXqaaybxxFhRMJXKnyrKcAwLi7itakOHPbx8p7HX0u63VcVEijPkMS56efpsA
8crromlthRafs+U3jraxmPDt6+cvopGExvYlww2n4XPTOMiyovP46VrFuaMXcK6h
cvG2MAX+DN/Djmt9f3F6TS0v56H70zqmGI/pMqmJ81ev8R+6bfsQZVwcfAaQfoLF
xW7s0ApDxOpgkxt6rQMFV5EUMFljKsWIUb+rvmtk/wS3+JVsKGlcTDJ5uCTcxRwy
dBp5opU6F9Xltisc353iviJeTZvS81ZCIRZIjFVJkME3EwzhIn25iMOsiM1v818E
7EdwXh6HvfQBLY3vcnONIHxD7VT25Lr9wH99fL/lPHIVMY3tQTmeqIF8Rwl4tzaM
33xFh0Iihlf8bdO9iFhAsvueDuB3Y2CLvWEDAl/yeV1Zza4nbcZuPis2TPj+4k4e
DVVpwv/4cNie34vEyxIpm8ecXLdn3uvtR1Zi0f42yBTTqTu9FXhaX6TSbIoLGkJe
JpDEAg4mkN16GWvEvKiOkw7/nHCux/DFaPmE6zMdEAqRbfVTaCo6ixqXf92qjkWO
pW/JtrlEQv3+gcXh+7WPm5rSLHByoeysrRkpP8CfP3ntWCHwE7Z7d7Kar2dHYq/a
FCES4uACtD4mt6uVa4rZPEOWgpbwfrDO1E359YoimDhVGJ+rG1fkmJwNK+cMVUJ+
4lYMoQBCsdMawecFiv3E26c+WO+leeCqsNtai3QHsSGNFD6rgY47fBPYI3qd3EYu
o3WaRy57WhNL3P5lqYUi9Y+/5GMMV0yEOI/ykJtFfGZafYRS2wCS1qLRkc0oWpM5
m4AomKQi5l0gfGW9kIndj44lX1ml453reAnb9TgGwbkorPWqoxcRzqyGnTMnZ72M
Cxr2k2pWIEGpXI6IsXHEaUpAJ1+khikY6G3df8ogar+SAOLyncUJNbi+bp9l2Xw0
MhOJMD1glYwXHPKeiJtb+DdxzYFkD4yDQlb9JOJ7Q2lmALtXXC9voQSlHPe2NVNY
t1J8cJgTRP/JGXyq4xw3cq76h8ERgBZAGuXi4OEah4H+MS6aOQfj/LyB2SfSW22J
62q5iQC2l/7BVRI0uW29liD1V+S6E6hLTqiyZvGSIQf5CuHOs30oTnCN+UERRsYl
X75hslDssFsiuKbvCKgqpBStbZAZgjgjx3O8jpYH9gLunfAE9zyUTbbNeSUuHSIe
kizLwvGNnK7plblG5XF5b6XngqOf+GI0xLuhbfGPpIBx4DJq1cvlRoBNILTXi02C
/UL8OaidiMhzaQBdr8XNc1UV/DQyP4erQ+Gl6vzmjoL8jMS+Pa5Yu3Pb9in07GBp
3bL5jbCkL+tZq7lIxuU0KJd9sAyimjtewPCDxOhp4w/QgFxcUHfhq7jwRs53/mzj
2qrkfdB/hii3ZhPHxsthsrkH8lggQJsivRA+njGmYAK0UBxLNOwVT+WXIFV3czaC
EE9Fs2WkBueK247nKeRDkFkATPSJ/PtNoklVs1wMt/8gcBO1y0usiXf58Hse8iqH
2MpK9KKIAnEczI9x2CF1kdXIhgWp4VPxp9u1b32PsUIrGweyTbI8JPZzGdq7auGl
1iHQs+CPiOgCK20P51B6+Py5gHe3cSnBI7WK+YcOKGandlvw4S4SYDJze3pV2N+k
lj9rS9sFyNa7YG/TaBo9OEaQSbEJlpWgvMRh4A3heAVUmyIwacz98Q5Wm6GsRiPf
aLreLmFZQTYWVa3CKyWcOalzrYRfVK2qnU9xP21ldd1N75FhDXt/pAG4LaHAZn00
4AOKyg8m/K5J1vDk8qQippQozgmc4K/oC9qLCnbuhabnDRLBBOQlMfCG8R5yIq2z
nHWjsFSFvuWSeWgxrtBJiFpiJ42YPi0RAjXmIpUEx2GaSNGyDeyZe+h7UvY4ZubR
mg5ePBHyTyky9rleYqjnbdGpYqWPGyf7QiRGMD4sE5Qiyv+hllvsRj4Tfzh+UNAc
f2YLKWLTTh4TQo04rSaP3FVWVMn/c74DN/xqdTNV6ZVMr2dN1NTP+LILNIlK6rLl
GbzkR7jXReZGKZK+wB0gAQ6Kwlhu0mTdYU8grUfIp9sbK0EGZrkn4v2Vm24OPgoa
q4PaBPjTb5jgt9ND7eQh3MJumb9yq5HMxZ4N8yGmHYwJg2lZz7w8WhADSG6p610L
l9l8VZoBiZsGEnEnI2wiKVcjCBGmokbJ05+U5znxkjlkWVSliwNOcprawImEQQMe
juiV6e41tBIx98fMJsL8d7Gzu25K0PxJLNlTthRwEZWMF5kqWMZxdx71dh5Trqq2
dcVPJYM7zwhHsZIHhO7mvYz0ezUkwyXyWQfSCTlizRrwk3k2EsjPLifgkyFZ27Zt
W8mTz6tcnaQz5NS0cqXtTyrdydK/QNL91t1eLqMydoQ1qF2Tr0Bmop5c4anQ3nfH
8gvSctyuMQN5uZAKkR4yFtvJZKonJhxVGUNoDIvAdaZHYhiLKkZs73oKZpYozRg/
UeBhsvzfjRjn73E4fFZNNmYP8ul9GAk1FremdUGT60l+jIUBUCAzJ/raQ1hpAaDt
PgwniynZSda87/vWuE0HhfFfnSzfWFCDMF9cO7QRNvN9Zk6NVgD4+SDSyI+wHBVC
oLLRBKK3AmkhFr2Iq1XtKDAJ1C7wTYDYXAN/5LmWey9/gEC2KmvtZjVDSJYGasgN
jnj41tX4TpFp14Mdbpjdp4JuUkbkNWRXxUzVwkvFlVGl+R42PW3XvD9i4qu8iSA5
qWThA0F7xxGX8jXA3XHxd8xyBbZAWFZl8W/wZfbsBwJKNQXcB8JL24EpSUc7oMVI
ibhRUoCOuGqtou525GpLC2Zy8puvCIMLiksXwbRP/fjo/V0HCv6xj2qC5hcFNzuk
nPdS5Ufp64CcI5k5XUguQyyQVpHdgAWTDqKmyS/jZLZqToZ2yYopRTB4BjDpp+V+
gh95mp1HQj8l8QsxrcENV+VfZ2QMizj0ugcQeYqVWI3qU+C7w36xLWYsahROUmoY
FpsiB9YEZkyacwVJJ1+VzwCWVAHpGI7ybqKr9DjMY/PG/i59RhNq4VDadKrIyhSh
6b7TgkcJ2Kd+ZwOaxJbusiApE1HVmfvuYDuJmtm8Te7FSbSEnrmIpU3aLezDOPfS
MqWW6aV9tHRzBgg1PwQc0U5qO74TmnKvuV8SjJnNTmNcfs4D2qYFzqzkJ0qcE4JK
Xy3nnBsqzHaUHlkOpLpb4BfiXaqCyiiVYn1NdIrr6JphxGRrDZ/0SNgHnXH8kpzb
9jxqyCK2ZeMRO8BdV/YmGz7Up2aFs8boPXHrr5zVoOEKiM3kftskyibcP3w9Ifg4
8v1hJNMWQXleuJOEpvJUb4o9T2H1yb7anSseQc7Zn4L/zzkjJ9//z5F71++0T3/4
TVKJC/BlYzCwGSfQINPuG45MBBwME1tOtoiEp0ONKxB0/7lIn9BtSrZCrdDilzC2
w0dFRbh5dqf83WEhHQ15N+aAYgHrx5Uxmlkuznfdlkpc6m2Ah7DtZC519GhU9Ups
IEbBY9/IrvYHMCfEXD4R3N7Ej7TX2676kCTvTvwWoFfoCN3uKVF84MdFtEZM1w6H
bkbYKNRsO+ZuK7sA6BeoaFEpD3j3nE+xiJfmM5MNEqURns3S2s3GfeZXpSQswHRr
SMunz3PzrtG59svJ3LEspDn+ndljvT26VMFm2xuYJj1xoD2neYgbsbkIQtjdPdHX
DyQrJr7TPxv+z/W5c6g99Ikb3h7PN1jBJtbp4S9+ayICVLRVZvyz9RHZV5ezQK2a
aRs8HHt9ujrTReeOSExSYUEdTDwLZK3ZcvxLoNS82Dp55AkvHrxHhlHI5dIaCdar
F3Dm8bAi7Na77JCGQ9doQsUiHYTO88P29977e5TjGJ+/DZQrJxtkMX0QjTjODKLa
LPrFHdxK7yNlr9r+wn3/ObJeG5v1vFHoEuFmvjnNe7uPSF6sMM6lZWC01Eb5bLka
BJScLqC5LBzS84F8Volp3Rm8qrKdNjNYc6g7kmOwp58RAm7uF4Zy+cSWJ/ycis3x
9LN13MqDfddMVs7n7MeiNOmbs0ZxruPcLRq02OG4/8XvJKrDdBljmUsbhPmc/mTG
dIcXOqyuKGeSRdThu8yl3MGg7fXYzwQJgDNK63zmSsEe8M8eE97nS0wfove4ZTZc
uM6G058FPgOfE4MyDObL3bNcPcicXvFYnWtg7/MSYuNW9O77hQn6EHAnzmS/ZyFa
OKTSoXHItfIM6mkIdHThUe+YyiH4pzVfAWLgnmgwTDn860Vf0Y73t4LDoNWDsIJq
Hr4/8LjnEOJkrkm10ZXsJ6a06PLcIlNxbQ1a4bkkHDGK//ROaWyAP/TjfsRmBQX/
y8gDjvH5xKwHEmI7eDuxBGEGy/HcgJz07QqA+adxgFQYjwuY4rUQzc+tAK1CHPWT
SGkCqvVDb3i/8LhRzKOqGpBQqNgpH9i7ulbmdgtQxtbGBk6vMnrADFIQ48QuqhNL
yWPxqoufq9mg0I10iVLcXsuyVXPTBXFVPVjV6t6rK3cEu3migO0bQaiuSp2Rw/uc
JBGQcuproaHTRNRNWLWlIuJR3yjm3j1BkD9Ur/h6eETEVzylPtMAZKDutgOmn/XT
HbfVmabJsitqWys9/+60ujbVWrYJlGegdMojR2Rw+pe+brottNBsqRjOy668dRJA
ciy75zLS6nMR3rSoIibQQT7isxJN/e5Qc+xfuxj4VI2GfG/vF5iuX4LUAOM/UxfI
2P2MnReEwKGxBGC07IbgqkJBKH4fJKXLWDAXEDFMVsUeiE4braOq0am2JvuO6ld7
p0S6GPfHVTULjKGyema+hfTxGMRmBq7nN0RE8Oh0EgdvtX3WQh9CBmB+PxGpxxaP
En+F3VVx//XWNi9ux07SGRdtSy5JvacSJOu4DvlsbpfhuhW7ZtYe4iLKV+8lwKpP
gANwb3Ac2LlmDRdmzMYUbbkctPQerg4NUr42zqmYHSsuxkJcr0+X9NbgFCBCfSD6
w2JIa/iMzJ6OObMKqQWJIDKZS3mlAlJGxW0rW6ui0mnH090IFALF3dfI3RN0E3o1
OU6ko8ArkMwwWS2sU2MIIyA0ZF4lCNdzYRDBUeYMQsB1s5dLt+pf0lma8BjALgkG
vXcKf8/02Ul2fMoljWs/pC34Db2JAEr4lopm51tqJDlNi5PUXAojsOAaOMSSmhs1
EbGwa8yx/YfgiLwR3rH4DC9UnkANYa5r+iZV6w066JteTOEW+EaLsQY+FBpBUKx2
nI+6bbxrrqk7UkfIu1+wn4ykH0AnKxQAClI2nlZOr9cRrpZtV13TcB6k0aPvxbIU
bFxwLT2CdeZilaPH8PIAF2jcoUv637HIdsbLTRuWXWYldxPAqJrjsHFmFHW4j1L6
7drstpPzFy2Vh63dgezeWNE60IuDW1duFXilwM+77t57ocO4dhi6su6hfokhv7Uv
07SrBb93rZVjKglXssr+KTJNiaw1g4DZzED9GUk/z7aGvuwGOvU1W/u6OLfT+LCA
CqplLoso0rmhEB/6OypoHyZ7HKfiSOHQJRbv7Kv+OTbvwfq4rCWPICxJc5hHt7j5
4RCUzvz6nHlWp4+Cxanad+3psfjmYA55Vo3r+k5u0aUwYA8Vkq6d6pMiapoDudki
KYZxw0LdFQovUf0XUy64xxpPlYj9zZ1b1UP7TZzGBssXo+QXAFHswSlJ5wwKtdcz
lVf+Cyg7VLYgqVEAKfvCUWWxf2A4eu6CDre7nRVC9tHJ0lPZ3EMWPQLIf9gQa3M0
wc45Nr6JOPlry47SaJBlCOrG5fVKJD3DBIooIfEgNumFavj5qSjQLdert55pEys2
NBYSM7mMJ3hLk3ZMKbwrSHpWMc/HBPIaC8fVQbEdFqEkSTLsefIJE2XKgCRIkx8B
ryF7+ltNB9Z2iBFq8DII4USMi1YrfrDAhClOa0A7Bxbj/ttN4zB8tgB7UB5LPvRn
VyFoJVXU4ICTnlndowIO7s2JTup3U04a6yf/45lypRPvhOA/kFYdMuGVnkVhIRJG
Ec7m2dAgjhdvHf9Lg7ffDDDexcD5nnnAk8zFRVuArC2BSxErV57YzHPRmRJ7q908
wcbSuznYCijO8uZzRLWw3tiWyqqsn8/q5MEiBkjoBtjG1jUo4Rot//i6rDpwmDZC
HNWWzkJrozbUQJq8UCyHc/Yim5oNIAlI3KLZTQd9L5TNIRs/xXkDisZJ5AVsZpbK
6ySrsZDoE7yMCJrHM9iCXSyz7C+3BwTCuRK+ceGkcmAZjZcjTi38H+o11pK2t0r+
Zy5Y5e29u/Z44mXW/NZSC6Y6tDJfhhoA5QeLh+Bvidq+SkpG+/V5+rMLADwLDWIf
Y/dOJ1ztGLiD1WXIF5SoWfFJAygavOkCUXtyfy1MzXypZLWoetCqB7q2QEiKhYq8
0FO9W0T/ZWieu+CIgx5iPZjgduI2xxw5UpaarE7Mg336praJTKi3xmD+kZrNuHnu
efrKI3bUOIAYJCYyReL5CdvPvYnDaGO+mzSpdrvTWjiQKsMCGxNGmC/800nw+j5Z
EdgsxaZ1yQCnp3t0OfHAiyVm7O7qZ8NQQXJPByIVomnoBW1YsgOhuwRHBrMDhYmx
S1vUj8Oul79Yd7LVSOjU4ub7hdbIXbRs1Nm+40PUuxjr6Q5IFPwnFyI1oumcP7sd
he4z32va2j/jYDc0bEno380MYm4eHiSM4LSQpzWc8TGCS3lvrVu2fNEQBnSUrcUf
AKsGZ/E6JTI1+Bke7h/I0RYI+ExtpqDVd33XRJf1K7mxvflnNWmLXAvCa9SbyXpx
xh0RXyJaRdn8rKfBdxkFwUln4NsQUzj/4rc9Y9mr9YQpOYykfQ7udwf18dQvVB6F
b6Qw4pLFzIbnBTrrlkrCGeT0wKaN0Znq9H97zqpCJXtNEFgxyRIybHvGavzGt2Ot
wTprNkMRlc5yFY5igaTYFSVcSEZ1ABOSGKLq7qfzL3SA606QketHZdSHPMKohlCX
dbuPLqFf1mfuxrksb8ko+GqXukugw0o/evcbXREKEfr105eClLhNROd/cqE19XYS
SkkkXoV16861lXDU1X/P/1fK265fuy1TA/I72Zjm/nJgi7qIL6AO8kTUudNF6EmS
yFZ57Hj1zuAB8qyIn2H8PFWzoQtvU4WGQ6GMSZqIM6VI/Xf7+h2hM741dTZXvmGv
4NFGqJGltIZTThY8C+0lypRjMw20FtXfMeRam2vwT85gnMTMYwkqTOtdltQt2ebI
LLvi/3MB3+pcoYcwA56dkAjZ94Hl83rGTdabjx3heLLUOWf8gZA70G50JrVSoenC
WAxmPedWkhcBwK/W7t91Gp45D8UY1BP+9h0XHrjuPNMRCA4z1W2SW4H75x0oJqaO
/d6Ki00fApJjBlZqSksrH9/j+YQDWcP2qZD800EGCdwYORfWrwgNW7+dXB2CSLKt
4MXurCbxMyJlhH5oh6gug2+Ld2/edAwK3PntUwTUu9Luwe3JrwguyIO7PcqJQLQk
wnuuk/WyKvpOzLGHzrxAikiGE+ljJXN/eCWLRNGQjvtOUiDAC5cIvDRQd0dSDV0/
3lmhKpfq7SNZ/MUo090cMXZYj8Uh4ygZH/i8unKKga7KCKw0ovmEZdUOgDiSmr2r
2iEL6w6GHctKAsJ+5abzfYQhXZQO8pJw2TMtKyHrcEs8IvuXNKA7zie9Lqx8DqSh
W/4oql5nh3QG0jtafoJNw51pwSNPYgWhMQH/QP4+mttV8v2VTzhAJf6VuVytMrTF
jqInZ1iOju3df8QYFXTi9YYanr8XFL2sdDRCOIyC3dEmhVo/NpvAD0mV6novDKgg
kgOs6St57w64YW4foHNDdCqTjTa69tnuWvBYiZhoMmxupytlQgH6/+8oR1+tBclM
7JckeF2apIZXasenjvUMxLtMJdii+XIFA7PMZrV+A/1gttJ453RVwKLgdgr9oni/
wf0Icr74yD9sc/hRCKQhOJiwVLtyV2qhOWBBmXcS21QVpRcO8+D9ssSkceHilI2b
2bH6MF70Q8nlVioLieweqLXpwOOeh01s0L+dhpb4NaKD5alsHIpez8vqWWPWGDqB
aG3OXb5sJ9xxULcMfQWjKCVXDKQMiUij9xJCy7dUFDMuHqdVJ03TAgjnn/oIYlwb
meM2Spt/z8yBsw3eKZcgvjvvJ/gS1AfVqe4P92cHIcCoF6opghm6Jqxv5IFgM1Vd
Elbl3hQk9Spu5qh8D/C4IhuXb/PqfnoONOOkyhqelpen2RhVdI1ixzMJckqrS7xX
FNdzN16zcylWnw+dcJuj3MrAJPwRkJTCgcgEZv0gcSsNqU0YzgaAiQydUoo2eenE
pNYC/R+ljlnQVC+yiFvov1RdCz7l0cd0n2o5Hz6CAweU807KfEv5oyoesWVCy+06
Npar7WwxgYree0e3XhqwtrEC3zT4TFRLzXVzMrhnF+emRCxgy2xSqP70NwrVI46W
MCZBix8+9Ijeww252v9GDkelXPgVoTpkRQ/E1uzt0EquVQpd6kdZZ2JFYP7+jTdF
+lmrEd+u8lEuWbWlJ9wONP+VzQgpfMGnbApjJU3G2XQRsxYrldboUyXpx5kr+FI9
HCqFKDo4i6hcxsMndt3Cdi0NdUv/sMzEA8dOSneI2Jgg7GOac6caSYYAxEFjfYGn
z3q5Lxnf9OEuY/6yQNDtsJ+932cEUQ0zvX6pyhWXp0TWXe0+7swAmGbdue/ulwyM
hER0qNcWBoR8GSxiKSOUxv4qzX/fhmy6jyiFNhMegQbVhRjmrhImdyig5kkqOBBt
mWtDF5InaSrv79TJkNQ21Ek+4oth72vUQ2smzBFML+uFRyIzQuV6YfkSW12K3HY9
jyOExEHj0qszDxRSflfJnjcrKLZzyrdDi5tjnMmQVKrs5ZVOoN4DrQrhJ6itaceR
ea2xPtE+U1tuUaaoEs9s8AVGKR9rbu5TT5CXQZfa8ccpEYMRSoTnbu9HIgVDXbXa
yB/GCl172i5Tv+Xm+EhC+ZmLvv9I4nqx6TLA8XkOdZZ5CyaUVrBJPht1jaTtxzDh
gjdKV+zfPBLMXRj8k/ZFFKELUyQ+FMea4Cup9gkbG+exzeOHIFSbRXOxhzkudL/F
cXN0420eV+9PHQYHZRhUjzPz+tJPhtmqhBnIy1ysVDkyFTgxGcUv3thn+ApC2qMY
kOEuEFV4SjNuZte0/9cqFp0ntD4I0c3J/OtVC2DRtWQNaP/bRpnInOdRyjxNJ5cX
58u7HFa65GxHY5/wQZiarZpKhmHVY99Q1waejv4dfEZKOPfXgZGytPmiu5yzcfJ7
VPkC029RFMvbthyOMG7CkcNpWpJYPgSM7R35I/trYLHdCe7Ap/1rBrqKz2P8H9Jd
wQFlbjFsPq+l6kdGVy+5j3/jXC0ci1l7qTvASz2IPTWXtgMKbwPrj/qCL5Yo0R9x
PvB3n6xtmunaWmFeB7QVFknwFnl6S2xIOYmAy1LIl4j7Ne70fu4z2aIJQqnHFCCB
nlwjOSPRWN/QsVca8jGP6kaLxY70pZtsnHP8owMAHB7d67pYYeYUi0H4S3dDYqrs
tO0RgCQykOmSuMlBWJ9PBbvT/cOUFBcM1I/sUbV5Z9PN+EFKhJwWPVIDmJ0JAKGh
LD8FsiL4hEWLPO0UlMxdSRD67fJiuSnJL30eaeBZkuulUZGWydoxtXExu23MGVDz
+xRegR2JV/yltqUNAMdk4Cqf2jcw0Ju1VcKfCpIT/Rfyc0xqE5rWBAweit3iqolX
J2iIOh9mbbeRd7yc4muW4+PY8giQKv9N1JOTaiFsNQxkG2Wae3WJ0z4uyeOnuDhU
fiO1UpXaDGQaCYLt9ouf3cBVUdMEkDUxb4c2thBGJb65GeLtcU4yCxqz8vsEEdkc
qxWuKJPJA9LtSGInLZcOhCTF+KgKbqv9Kh/fIQwIz4nvSxdeb6dALwGGDqCyLTzd
8nQvoVjp0XTGo6esWAG6DeY0EHAQG63W00EQtuKPHGIOJkRY4nFv1HWAuSNEiFAP
Iz3PgjRDvXzDoYIx58p2mGDOjBL9enOBMDniaKeA06FWlwU1cC848o2exggj2qbB
QkEHWef4MRyekliWt3Ha9+hYcH54pz7tYQiZte7Fgl39/4BXiGkcwVwZNaPM5WR9
5+ReVisYotUvnp+8KV0y00+ZQeqO56YH7wV/b+7C74HAHn/+8orCl4shd6z4aOAH
PTi4x5n2YijfuxAsD9JPQezuS9EkOlVcCaPbA4wyr6vIc5s0ycfAkKaTUCb8Koq8
y4y0dFeo1EJ1F28iruPTMK0VNmBNofKyXr6HP6eLDpvFhqsenwaxgrfgEVxzISq+
91nEvr10WTI64Jhp/ZN5Eve8ZaB/cxZoZ7MyyphQjy96fTklSvbsZW++GxgZUGjj
pgj3Mr2T7nMfPo0A4Nw+T8nlaAwxMFvXD7JhtodeBaVzvKMq0h8czjx5GzyWMwLm
sO11wcvXV6uCsCSp2N16RwjMcXKvFHZCI+EvzYxkWcpLaMCLUAH7fgSyl+anNHM7
vvXe+juHNYENmNV6Lpzhfs5oo3vcaeKQ8IB1fSlfu4NouHYRcaevYFCDuhzzrPjB
w+O1+GX70Y2OKEusPmH3WRC4RZZ7kwLIU4iTOHHmUmItUInnCViWjhB0yDeddN5R
UjZBWQll4MZKdBMg0LU9LKVSgvHvwIIjFTttR8a4jgOIIm4JSaOdV6MhPO4F7cLy
ojhw3Gh3EQL25aX53/9uQFu/HR6AmHdbSrgLyIUz/nZexo/K35RdiFaV8/U7LwiG
sNm5qJHw+XAmsgPANR4BaMY7hRoNvjvLJJ+JKsSJcqPRcAqL9ZsDplHLSlC10/EZ
uE+/doTbmkSKmXwD5yBESWzKJTr/agydUxIoMrzSp+uSMz+7Owqyvgv2ujSMjcS5
gca/eYY1UKBqiXLJETDfrv6CX0Ub4IhcV3xYJr04wnT7dAtDd1xyx6l7Xe97ctGu
gZRStSYgqMTivKNjNfYvk0h16e87vJABw+Ojt8o5dbD6c0RPJ5037WFHcW0Wume3
9hJq2pmkt7mu6fK1XU2RU3SPZRzMTOtrBMo5QuAkaxqp8WfvGj/RHYkTPgumLCbW
jEsjb/GdJrkGLRk+DfFK3e+B8MK8kK5YEIsg3nR5SxKu/+JWvsIJt3FbOJiWL4YV
/XEGFCpCvnOfMUU7BR8TFBmJV8uS4008SX9rAJgS2JhiL8g8D+4SsIjX1gOSuJJo
TzV2LGxnAvzsnf7e0nLTT+GecBIIOm3UfVO4/5hJ3qwYyej6xslJcNkjkxFZ7ZnJ
Y5zliZCp8roFFfrqjYw7d6nC3XUCaJnVhdrtl2PBo0QmOiOeTTBkAoSmuZFXacOP
7pY/v+n+uO7RaneB4A4alFJo+sxdIFskSIAOKKuygtvzSyNXzpKo87IBhc4AgHmc
zjDVL9v3rJ5cycR5JeWtR7lqT5r5J4eCjdRYTAEEGkapqDcta3u+ogaF2igClZPc
cHS4W4FbDfXypoVhYDgvjtL0sxe6diaIa4Urprv59yGJ0/Rb6rF1cXmojSR0Ejqx
Q+Cp7Jy0gTyPCCOGJ/Ec8/RmUWgAcZaEJYVmYpcrmKhiEk2gNKqpiLIATIxRG7Is
y/b9N7My+VJZGuOiBLyYBsd+lSalD5dGckpQZFSVd89uDHpDmiyYxiAyIaMN5vxh
8dbxoQNOkm/dklCKmeEjuN1bDpZpyt5r+l3Ygn4I9CPbFWQ73h3KsZPkDP6uSAwW
9giHbyT+yPN0ltyFzy8tUExAKQFT8crHZ0haY7JRQjSFVwgv3KB6m/GB4JslnXBQ
vztiTSUcAiBT67geSyZYGmeFxJpuovEeKO1B7AzL6GxE2ZLCzxHNmPyRJwkZv1id
sCzuCmZM/w5GeyjUMCXBD1pJNiW5cJFAeVKpiU732r7jzT3wi9NHNhDtnZwC7WqI
c734qZOS6AmVEe4rUT9t7YPXBvGtxOs6AGCkp/FJ+5AbSVt4IwzPY+Vhgc87nblS
iW4pPj49HhxK7cq6Kh+K5FLnAODr2C+JYdRi/55+4jvW5o3HqdfkeH7PYT5CxX4S
5ZaeZRonXt3KUkZEbjl8enQJJbGMcKlFPw9Ah4nPGSqyzECNQv6jMUs5rNYMQZbg
759RjIj8UHnlk/5UYzwVXVRvp8t05UPKA7ikwqkNKM2z6f0z4Xvh0iU5VzEuKPF1
fBNWn6uCm7cQK208LuCXTKJuzKAKVqNpjfoboy44Nl8WUVrJmprEirR0f8HjckFa
ROctj4EXuqwU9/a69AL8lMDxIjVC6OgI/bXU15Lc6LXmqcGHeJu2ybDb9hq8HOlR
SwgSe98a1d1j3/d37tI8lr5k2zStALZTDgF3bfgsUwoQtk4v1aQvLN371aqZsUZp
ihnbztqcViiJe2r/8Z9tp9qnIlpCbxuaKbrtjNYeyxwaBlxEcD3FQdNCV9EfPC2P
/md7DUMp2pJ2MC78Di4Q6TGbamqpNzuhN+3zF6reCyGwWaRYQB05qre0ynIH9cV1
T2ixqoY499HAjqUYKVulMxzEzMQG2UQTHw6kYKE7KMIt9XFZlpcerey20BT5Hrm6
fEwyU1ET4CBFEd9Ohzza3Fu1MbOzOOV/NaMHxMq9SWwg/7JPOAm5M7xEne4+Cfpc
utReNpaIJU/PC9Zq9DsPmM3wM+RdiOQrbtJ5FBpDWDoOgm2FCXODzM/XPB2ugz2V
x5gXZnhk/tZYpIhm5duAfxpAQBOof0h1APd/yD1Jad8Ji3osd9o1GOmSJKcIl2wl
cOsqJk06KaqmDU6COMKvLvNdqzE/LRzLPjI1nsV3pYR2hsLw5JXxQk17aa8JdQeA
7cEMep2pJIhCz/lY4lDQQ7QvnGmCl4LFkV2MiQ6xIBFTLF53lVKgWGsWTpuT/W9g
hkc2CK7FltZk9ESKq4YD4D7mYXFEhnwqNGNC9JGH0yfvs/HbwGvD5BRY5sbfXxpK
ly+yPA9ATIGVYMiVYoCDIubixMglyTgzjadsBLJqUwfeHU83aXYv047PL4UmfUxb
CsHrlAC2mOxlKk02bMJ13i3eH8sF7XLvNmo6JFwiMQYAx2c04MiOi9BAd9n4pBCJ
214wlLB9J7CExawgg3tJfgYqLID/n5nJUzRk37KPIHbYnW+9mNu3bTmZj3TISwia
zgN6fbr0zk7RfqopW5deWdUmz5C21DrpnBXqM2RMD9GTQBPy4iY63lM+T/36D7Al
0RfW0IPhlN2F4UTQrFKX6FOCSNehi+ULY5xX+tpRzV34tt3unntoIF27dsK2UsuP
iDCNNgR/UoDb0IYZWwqCulCvq7vuyqySY47FZiy6ppwop6hwRr0W2wADH+lSnu+M
NFFqPBlM4p/Ti+qJHShzuB9LjJ0dLb/o/XwippHvWw+Uv98HG7EpXbDHS6u9W9L4
8K++er7YUAzOAu7fnY/ZruLIc8KZi4rT9vYpbhe4mAPWG0ZZ4qNKOenuKiWQOQ3f
z0DLwJpNUGM6wt3piTCO/hlvnnzF/eEbGi1J50AUpsQk0jDlPpR+Jgwct8V4Jq8I
C3IwbKec/D4Bu4N4sU45Vobb1opgmuMcAXL/FFvw2gTOasMiV3oJBC+dOOykRpOT
P2ySmMZoPys8KUfiZ3Ccsow/PXShHODAU2jGY4ZdyqfvtkbXiiUDLdC39x0oVJtl
wDOV0qj93qG3F+SGGJQPWwjI879Vqm3qFs1uSIc7Qj/jLQBOIu5Rh032eSt5XSOO
uVYXfF6xzDXwIotB6/88XYFi2RyhIwXWxE1ET5UGCAqsfRzi//dxuMBx6xPzm7OD
p5pxggAN7atMiFJfFo+oGckQMT8/P6CscSZUBuxNYPZ9XcJSC1hhleggzZ6EhUAN
MCW57IagnFHD+p6XD94oJn4fLzrReLCTi+uZkt9E1awOEq8mEl0Nw/jiZCJz5XH5
Q4zs42s4VGgCBnp9HPNnjaftbpEruJe0rryzEXqx4yfczvIifSC7js5JUQlQ0a4u
k1ARGKbvMKfm8FOUWS/lxv0fF5oyGb1drDlNh30ViUgHmIEL0MWlqjwLCwnTB+sI
tA6Tq+/leiwkJJZO/bhsRUJBk2sYzd/xC+AS9e6WfWH39xr3g+zAF+8aAhLdRIlh
JrMhqpthap9umLOUN2lod7hfs6MEq91zE4n82KGrA8eDNDVVlxL8NPY3W1vg5Qm6
Xpd2JALFB7hU6Bbose5XBPBIRA9w5pyboTYbyAdbRVq5FSyCy3uLVLws4nKrRbvK
t+He7jk3gpoVowtv2uLPY94eq5rtHPLddenH0Qvb6eWLxtRzs2DMYNAyRFB+ncBc
8mONFyaUzKIumeaOr4tdd0I0huFJlcEL3hsyxkDxpLj/kcB11fElLCpgbBRUktF0
bSDOZpv2g5MpZYfYCmsU95IxAnWVNgO0Yn7PCwkr0c/8F47KuZvkPHh3LI8jRO7M
KsxtJ5+8M4MlV6cMGOiaARnBVOdUw/7aZTU04loq2bhCo90aKkbeShImv5E6XqNo
dsc14V6OaUpAZL9QVgUmEkmUxMJ5t6SIw5642WyjbrULbmh3eY3S+UgwPzJ/o42M
j25mbJXwk4xVqT3Vx2cK6NjiiCTZAO1GHZmRedo7LIzmcVqxjgoh/sjAmEwY8Mhg
WXGYCvQYqMpf46IlSrwYNfqAlTg2H7JW3xmBw4FarBNow0ScX4OsmogZZx8cnjc+
XA34S9CyeWjZWeuXwMlf1SlaBm2jb7+Kv1OdoiYy6Rzw7RVgy4SWOMfQ/sh4ljHB
4BG9siot+sfFZS7WK2W8nkC7f6dAJQjdTHhBgLfDc9lgs+8FgfqiNOzQbkbpyqqq
3QIAqI8RXDVkzRFILNFJ/CrDDLZpxEFZ3xAFdW7hXBiAmndSOAMG4goXdt+PXzBU
XA3Ne91+M4M1R3gsUCs/Qas9SZCLvJ2F6EGQ/pFcQiTANlEK7ZkDdrg6ji2Htj5j
N+HX1Kugg0MrQ2n8h9dmzl1w4gp36eSp4z/OjR3bQCDEAST4e0BxeGqpSdz5UvKd
9qc6H2BMwJuR0juevew/HphxIxPEMXgs0NtZNKTyq1AOcSsXZWGZ50B8VpkRnpst
LwtVfZ2WIoC/II88g3NP+qdxJN7e2qBWOW+thoWZLvwF6970DXioNhhZn9RwK2m2
ay2QqJNrdwmHuxUULwiK7U1eSFhsjcbRCo/urGIXtYZ4Gu41G2ZY0w5bvKQQS8nn
0MCH6F4iYN73jvrD3CmDWtkrgEbo4twTb61uTCdoES7XwH9lPHcSXkZ+Fqf8ViUY
F/YFfGNLAAjhpM7zFmwTIT9+cVgj+KggRJPjKZdGl0WNYIXdIcti5I6RcGU5Njdr
4ZPBP+V/PwnBIZ389fsdSxYtERY8r/X8OOyoMuil8CVwf4kB2IIz31zYxf6aj2ns
LGiTxg8xvLB0tCwL5VAmerLlUXAG0rESVE72sMxCDGYrp1iqTTnlT9tWAnztgq5e
aGzg/S30OPqCvIAD+ECXtP5WE8s0KM1ZLTC6A/RPPOu1sEwmTRnYWXcQpy9q5nDg
2S2Vq3lsMDYfr54uSzYGoJWpfmtoEuMqwC1PVqXocyAeg4N8NSwnSaK8T7YlNS3j
Jzni3KuOtYiR0vLMSNokZjZwQTc6/nnns1CuXTxuybQxE6cID7ODcYwBe1c3xV+A
q6pkBeQaWoNI27W5JhV06XTlL1/fZuCTlUwOR1tq+6rPs5mAzzKPewp4wQmPqV8j
qYEXI7SZVbLfnpLd9mTN1ue3O/WD6B2pCmfebp82hruhY73BT8hwjiLu5Q+WPZPg
A9bnTrMcMmu8lplSFCuwN/pP20ewTRnh1yBlNfr62Y355ZelBMhzrTIlNmW0Pe1U
OvaFM+a2CZ3JO+XUvppeYDSfcP5aDMTCUkiX2jCdhwXbVoy3FFjnhS0PmYsd8izd
1XVOz58xxzZDgfrpjcl+hc5BnyT5SJlUdZoyYN5Zl/WWJfUX1jFnM24De0oXJ+3V
37Fhl3e1Qyf3i9AbJWfrD1lUXH1EJEhQmH3eBx8ZBv2scKGb797EJZ7v3Lpgo6ZR
H5iBZDpwsXBSPwEWJ9CwYSRt/Ex8b8ptEeD73A9SDp2xhlghMjL4qZAjmjI934Oc
Lys0GI9/Y+w6AUQEXXSH0OY2G22XsK6V8KqmqSC4X/G1Napt9hEus99XdUnFP3dy
1+AdqRE1Hy/Z4Jda83eeMLYemCuH00WWjUGQsOmP38kW0gAXDPMOahzCJVGOXXS1
Jb/vte2bhSyMUjru6N8fqra/jfVg2xkAmF/nXhlKcJmPhwobi2/qkjFhCJgJ0RB+
9AI5hqhRG4shp5Q95HWv4VUUfsj9ezID/iM+latK3APcojsemEEoQ+dadCerhFTD
629+l1ODRRnzODecWgAx7OfHohtuFxU9l5Kj/qW/S+CfY7f0Nv5sMwxXhed6szqq
RNX0sNCWnTgh/g+CtjmklIbKxHXwFTFoGwHpeJM8D0uDdJcj9evQkiQoduWn3GX2
iDHzO4E5rrMqA2we97uGbXPBuFOkxF+adl6U1c0NC172NA6lmwCjmVbRj8e/pYIS
av/kAqrGkkaxl8ty2uYKa7Y6kwSDruW58nPKstnTb3zb+Ai/VVuRGng1qehby9xX
lbBuloE7sHyod8ZDi4YTkRtJ2UXFhnIGxC4HzZwpsDPJJrYcgcJYY9NErZXkvXwU
cfQybK/lJt7rkteteVEmlMpFvAcqF/VrLpuEBod1GAAeHZlmjD3xsme+igYS7je3
DovOB8KOuTveN9bCuNcBtKLakYp1WJ2yxlxGLFA1jsvLsr5kFpZV9c7GZcf/ND/W
6O4+/Us48b0r7wRB+CcAYDphqjg4X7+rVWQeBnx3AOULAsYOr3TM8dYM0NDHxUgi
mBZoRcxFljrteArCnJje2OJgg53WdFe8ed7e73jDZWIUmsw9ebpXO3z8ytY85mfB
JGexEvIdoy/awxC3+08RG3YtuiXyDuXh3ZXagjl1JkydHKs0ujzkUbYB8Iu3fEJr
0rJzuPPO1SDU45Lnroo6vpAoAL0oYvGNKZqpuLmggQ3aHyXQGyYvlTCMVcApT2z4
DUVMKEk8Ngtucu+udSNyfgXWRL6HudlH0UVzJbqTm0sHnu2yBcIz/W06Qz8SS6Qu
+++lEtbALKKGjpeA3KL77cIX94w6j005e6Dz6m/aKUD0RJ9ZjvgfKeEO12zglwsW
ni3GV5nrachQZRsbF0TWSy98eqPgAlF1WiqORtalyeX1zT4XwoVHofoy8mWY4+qj
2gO/n9uCMhzHASYv55Spx+prWCpBXOpulPHfvrHEpcAqfqaoa3JWp1VnT8hAduRu
35QJYmx8EqPu+jyJojmQgH/v/x7Hv1/jI6ON965jYnlA5wC4o+yk3hPT5gcUS/hO
CKURcaEC6Nc+O4LY4bmAN2Nl6RInvxLXAWLuKzuZa+xDdyUkWXiOox61twziWEHr
lV1sdy4AAvgBK+rIJ49YuOECpacFRGuzE/PJls51/7rmw168cFBxJVADoRGByGUL
3n74foy5lT/6/fk8H0/3xOrR6OueALoiWNA+fMAaY3Srry6ycGV47KbqufY+4MLl
vbBtxFf+ezZdLsr9RJh5yedKA2aOux2wlrPqcjhPKFtLS/f1DQ9QctPZUrlXFhJe
OOGRVowjG9k67kZHDasQ9MTq3XfE/KLCOPsxDSXJrJl5YQ0ONlJoZL+j9ZdspRfQ
+QcXNh6ixmVvs/ARR4ZHz0i6Qc6bcpEhCgrlS04dCm6wl9XC9k5ls7cBZy2c31c+
wowy+sLG5+uOcSt6iRUssvHo/m2gLUfArdInbJqL+5D42OOwQ7Dp0uDILf1HHBqL
i7B80t8a+sMSphqeNeMsJIKoibJ/Z5K3zeDOrt+SAZclVydfsj9053SF60kikq7L
ijSj085ATOPeiScjANEV03+wI0wfiXjwy53bZ+SbK/mYPcc2X18wJTuj6aSuYqQf
bwm5kJpgql5DAFPxHIGUzdI+Fg8rE4tGFZ42PGim1kWEHGUv/boeqjuaFzCF7G4V
3K5oA8oe9CR+OyMbjstHlvyoosSmEZg2q/qE80gxQMSItuA42M45qA4t4GttAh1w
lz8s/sxadekmXFNI/LPd8kUAkOT3Tjd5fPrc9eElCDJv9IS7X8Wnluk8vm4IbwBb
CkO8qwvX5r1d9V6M62SFH20pXkI79JWluVUOwgYG3oLsYgquoFkbw0FBCWWiFPyw
PTQRuw76ToxwdLK5bZfn15KmsH1Il5efYreSDfPx64PbL9RB1bLtRxmPSRhEoAWC
ANiQgMKfvEY2a/rvvZf00GXlvIUet6Bzn7YFzic7EGPw2y9vAaLw0Vb37o7Dccsr
NUG3F4yOkL5tOB7HRx6mMrrPGVPa/a0qHECi4XLNuK++CSqEona7feBgvlCkMukb
Z1fUhkzv8OB8ODvJTwiQrt9FDeVP4jXc9S9UOxdriVDTmP+P7yCA6HhnLwKdUd5R
MGQySTQP2fTUiA9Plp06ZZhHHSruZBsaClWEg4BksOywFKRdZzxw5RogRWZ6t4mz
f411tQAOPQbq7e6Ms6hlhRKVFkHZTn8JC4bHpLNLVEE76XC7XwN24bKIaJyhOoJe
dmUKPOjPjXjlGzKDYQlIj3KMbddhBqxcLg/fOamdZSGGgW/2HkEAKWNOU7WfakuD
mABqocgL9XoOvkzgYIxYZbaHDFcYvo/rBDTL6L15pL1VamxtvrSBXHeYLk+i2gyi
4gEXC3YYDLBTnTJRUqOTAQFGb8nh0aqvbCQgXcqJ1jGfZkl6sEsfzUPQv9NXAT+S
93bTTMcLeGEQ9ULgJV8b9CREYpOYzZ0tni9UFABTFU41wRHiwTtTU1slo3pwxATf
TltZvubCIzt4jy9VMhLuOF/s/LLdlziMWwN/A6RVu8bR4qhEwr6ZjirGkb/g9efH
HbIfOckAhR6aL6Qjl/mYKXmKUDRmKSZg+E25Qcpc8qVX6EqRwIMyMBJbpH+LYYNi
OnmvexD44y7FsYEp/CWeMr4CTt5w4psbanQR+JDztpkMjfcN6VC5/3J2PWtp8N38
chquLGJkDvRkdZAw4J2VD2hVQHBLi2p5Y5WXiNbzraVNwRK3iuJ/qsnAIX//f5Zp
ZyTsrMKkUMRgqfZcVXZT+l+dcAK2ebF9TdOMLw0eKffDncwIiy6DTMBkdmwV8eIR
p4HOBOz97ox3n03bufnNOuik5MyX65q8ecAnaZeeB42HgZWIgTPRMDxthPdtyMSe
Lan24hO/R2rslhrJnBYL/ow4h1/IMUwof5JfyXIHJiDXDAkoVQhqyQ2vgEXKczEB
e4dpqfEj18d2nYtTtxo36m1SzUDke20NfWTVXAYLCmK1E4EvOUabGUxfMyEWCvid
r2QhvFbWY6muUqDxoCWCal77bYOKXfegct3Dm3h40jia1TsJfi1ZIccvlZwzYSf9
huFjq7ydaF99fR22ke3I6Qjg0YbV+cRrIZ9/Somt9IMBHTxbMzw91LAZvpmLzmNM
aHb9zfkPcAQPaW4GfPFbVL95gmS5qoE+0CHEK8ObLUoVtD6Hd0fKmUi6AlwYr708
4iQM5cWaV4SaHfyCIrKtTG5ViV/uB9jbGid/0huODlyiMU6Q29ztYSGCwlopc9h2
BbGAgqXIhjNC8R3tSBgSh3npTG/V6UyzHe2OO8Jcyj+thUHl7+BaL6EPhjIJ6uWL
IoLR/VMrN77p9E9GnrmdEELj24jfbOmJ62yTU7L3M0N7anmoafkDQHXly+jHme87
aS0HCidlfDwBexjIBk7UYbkUon2ZCAMfUHZuTRcqRncTFAWD1mYUpikV8kHgbRfp
P/VWUHgLx8St2PQz5rhTvXLPRvTXwT/ysa3EsNxkRM06cFLErA0mW1APOBE76WQO
JEFJwMbyk4kvvFeV8z3x+Npjegl8zqelek77800/JlZUyNRz5e88SW7L9C231iZu
aBGXaLEL2GY8pV63ncKe2WLFkF3JpJrNW2N6P9Nz15KPSPS8SNdpf/OTth/slHcc
CVi5NX654Ws7zci5BmRCJ0AYtWz6xw0KkRX8piTKy8i+GZqb51ZxUGTZlMyQHdMl
weR8PFORknlGKZEcF8Q5hr06rRtEyMDXu1tAF4hSQi6hQFMtJ+EW8NJ1dpAWmBfx
iKAQR4Jm+wDwrX+kn/vdjWM8I5FZFzsoffnyxzFsORLwadGmF8i8q1eqXAPbasun
OS4hy1fDsfSDXBV0wkXTEB2ns6mYkzr5v6S9UhbE5F7M05J8WwedlcI1m0MahhyZ
GWmuXpi004UCOqTCIYSFWjCSmi83DQAFiCZRgUoGInTlGa+wLzTAoHxI9lJSXl8h
A5e6lQ75ETMAcFrz+zho0JWJbScTFvWZeV5tDElN7kyL22deFg4eo5OREyu/wQ1Y
UFPQA8MwGN+ILuxqHWm5+N6wb8SiZW9X5KW75KToQQIVjRdB3N5zi3W35lvC9VWT
eCnZKjabQabWQ0yx6su4bGSalYYXzSAZYUYH0N6JpJgXDEvwfaipyCTMU/0HYJxI
2EibMok04YokdFAxgOMOj4+E3hW2CEB4kyZ0hSukRvqpPVNgne/yNBMGgKtyfy96
/3yE2Pv6M+vQB60Pj1ah1UrdcP9DJQqOGk5eiOxA3h3v4a+7urVwq3IS79PDORN1
UdyZ4R7aG6AxTeyclbnYGH8omf1+vTALS7KDXUCwxqWFomR+0H2sbDKhQQt2gBBG
DuonV0bkq48YJvOXxj+XTTj9ui78e71E1lWaeuzn7X7Ed+/Oty9U9OVRkTeqdWRR
GrPn3ZzBxdlwitR3GTNCpSlXqN3BA3vVyGeTSXC5fonaIK6rVjWjDqS1Xqqp8IGR
zOZmKbHKoobKsyyJTou3Vp+z7DIGe83tOvmXi9jpOWSWNpgXu/+2lezixt7+n2N+
9sHdqjcHLdVh2yOH1EkwLCTlpk2tT8lVA6M58DSjIqTYvmciDIRWn9vnLWWXDtnP
h3ppn+Ndi8KBL80Bcy2Fx8Uf+77wgVA5EFWR9DcyjdSNtJLKHf6Z13F56/eaifYE
w/KgSkE9VajT9y3LplOODrsMyfDCbw7x/4Kc6zNum5kfLMENU9OHe3XcRb0YU0QI
eRSWV5VAykiegLQnAZQ5McI5xttZVkzE9id0uiXkgR4qq73iQB733+BxrrWHlMvV
HyHXyqgEJhpuiWu3MCUgnQil4mbF9T2xkSamxVPAihNl2m/NR0BGu2b17Zd4xX4q
EzlzVKnaVSwOS8hvC4Yi7R2uom9HGUSxsjoOP2TER7XmUi9wdAqwa0LEYs7L2Sxy
uovaVB6KQw/Nvz1qwFkAKUuUnWzQS67ywMhVbUypX9aLQBS8cngB5k6MReBe1fIG
Kmq6CsjwDglZvMpLSWd+7n+bOTqBqaChJRqP7jWtuEqcK/pqPoeZLHKI1Pb1hovA
L5uX4uwUp2f7VuHho9pxJyNQ68EQNodXjMlioZavMu22tr7i+tLXrZaX39XdjtzE
wyja/hT+Cun4zZks5VJacvqBB1RCRcWDK7wMur83a5DVzn0E7FxRwWGMJSbE6jNc
igki4B9abxnVoAvBSWgqATbwdtk0+wYGGoHMeVwaBR5MQ8KAyuTVyXJnYMIpqxkE
wYo3sXgB5WbcB4k46K65NCZZwC21fsY8WQUrufk+l7p18+dun7VN2WsixKZZnOkL
XcsNJSJJrZaKCncnlGhfvMm/HP88XLfVA+5bqVvXlOr+/ckbymxtpuKS5Ed1zCrm
24YS/tQgJW9mF0huFUBZEcGEb40RGN467PshtQs50C4Hx8nyHjGzIdGaS2JYM1Lb
UEf7zO1LbnKr/ZSvyVE2g46AMTLBpClbeZ34H9WKIpb86AXCxo+w+TYOHNhNHG41
7SYiZaTvonATLwshAs3eSE3Q39qXakFZro/8wz9cbfAMKOYUGSAdllEqVXynSOmZ
bvJt+AlkfOkvoRPtRqGlFZdiwvrCMjwlOHubdBNBlDvtwHxFlZ9G83pGlFN7t2dT
fsWQNM6Lxmdb0qs4P+pOYZh69Nn+K7HLSVnITr2la0JHvTnmhiKGjN7hrQ4G/KDu
da+dW2AoR1NWOnZid4NShmXJzs7gGCQI8VhVTOlWc9cIpNYmPPk41/TqOzsQe68J
ryA8W7Tiae89A4/wZK3lFS92npBXx14jy0CJPJGBLJJL4mouzxwns9Ely5jMWvku
8obpYdJZukdo8OmFdudiv0DTudMlFhG7W4QxKU0p5HQm1x0EmOihJTmKT4YC3RdE
n3p5hU9N4DbdLMzkiksUzAEmXGt+UW9zzHkttegLPrzUnkMy33kmm2b3GdchgHUE
amBoNqQtByVzPEqwCr9Tx2guaZyXoN9NSFkX691g75jVvnFnVVXa8YRVKUy+U0bq
EHXHaDAtVuKVqEBzWulvjKGsAwlTrxXZu+1480CCtXSJA01KCx3zLigNUVaJGaoC
xlNNm+WIgm4uxlM8wQb+WVQEy6+HiycbXr5iLcF5PEE4Gsr7XGlT66xhXFB9wSoy
pBj6srVHCSQpmJ7lOPVkes6ID+jg8nUwLIVXk4n4Zrvij0bsuT9IZGN7R09FJHh2
SdF/vxxuem0301ouvo9ecog1bnpcYDOcPxnuILrTqSPKNAZMnsPBL2CUbhtaaqNT
PXHbqHZuN0qyhfvcaIidiqtWWXDEkCuNKbA0kNkG3FQ66RJoV84GBSIiNFTuK0nQ
0g6wQdT2OObaPEHOhu9+7AAHqJSsoiQ6sAmYrIk/73qDhiXoc3/dRzi6FHpMWfmt
WXB63NqG6N50sEh3OYVMsdelTSG4cNW8uOhh49VG/dNvvUs+z/oegu5CE9p/XIy7
B3xl2cL+AsfA/UrzjZNA7J2U8nxo3Br6Tejrqle6EqrQYp27BQ8boD3/Gs7HBVJH
8GetvcCrDTmf9jeBIAsanZSKydX1iDWHOP6Dt0D0jNTZ/7gXwB/RDFVQDTG1EWbN
gjNOgw6iZ2UlBrcFsEbbm86utyjLyyd43xVGTnqBE280Q5yRdKPSYt3kI7POh9sb
HF/x4m8vAe5YP2bZYNgx3AUvovkaDunUGSeXsZLpBn9FPQJsDsV/1l7+Cyw0a3iF
Hl899e5w6eacnWxqc28qdRYsOcQNMWpJqmz9fxKpHVrihbAHIrHFV20ocPT/sDab
3OI8+l/Y441fsM4lENhtt41LYy0dflqSQv69XG8lJwZu9geFAK8q/xGhA3p4k+92
1FckG+je2e1vTEBJ0LiWRAGmQjqs7SQCxvVmoY4r621VMPleKW8S4TM9GONwP9of
JiZiMe8rYGIR2baNIN6c2s/9KC3TbiToftCcvWT7fhhPMYwCZ2BXNGD63Z1K2NI3
n19Fo3zOJIdHTFwcTa3iNMnyf3iKV5SDMM/s28rXtU8P7VeFz/U5KbeEIzri3/tE
lGbLNLNEMTK6TNdkOUPcZOQR11QRltG32roVtukal1Wg0YHtJdCZ+o50LUyCvVOs
O10NkJZhyB6wZms8O7tvSEWS/IaRqmMAyX5FvHL+COUwODnv4Y8T7fPrg2iS5t1d
VXsHS08chSIjwMgCnb93JBLMVFzvjGPDOguoTPTGpfA72JpTKjd3DXZPqPjvD4Bl
hd8f0JmaqNQ3V2t8dJapsz18v+MEV4ISGbB7HOxDGQu08w+2GSTS32lOV8jeMNA/
S1L1Fsz9d85UAM87MKuQirJpqK7tKgCmR4i4Cc8EDZBrs5/HNbdCe72U6F8qLpoT
tXb9IE1r3GUIGFVPMjd+mwjLOQw0kKWCV6R6blKzemGkoOd/X5FgwQ2M0TbHpudX
0ppuA0NI+NI2dT6z9xl5QgrX7O069HpxrsiKi5npib+5U9MQXlf1KcnTQX8kdjHF
9OXPkiqddeVpAP5j5YlP82mtyYfyXe+IGf3C8takjsgD3ehDHbewz+KlA8+R0bSj
fWiYJtqYZOj7uNLbqgYRFPM/rm+ogoljxNzHxm+s7xW870B2bH4QfIAyBKDn/qJ6
9kzZ80x5ncfgpSmWkQbjDL/dCupia0JuiLPk48reDfLroM2Noc7Hx1rdXDha1pX8
VS4prxlpkSLlga1IXHo7uGqDKDcKgkHIswr0jQH2Gl4aTqytxCNwArpfCA1fI35O
ZaCLowvt9UxNSEFLIiyhpK+hOueCe/OrV3O4cj2YCEXf1S67LWJWCd38n27N7nLA
OZ/sSlU94rHxjbdaVcueyKR4ZMEEzPuffKfKSTiJFw3pjQU5PGw6K5D8rdmg6RvA
DD0hp5GkfhOQJAxfBWkQjYICPe8NPrtS2eOJATuEI8OcsHmFY7+9KIbC6nZpVZl6
WCnB8cJhyAeNhjdTZjeTYxtoNUvW5MI1wTP31k1x9Ad5xSoGKPY1Acneg1OfZudM
mAhuz7Ltps0q3YsOzV4mCL9p4Z25JgwfnzxMfl76/tR9/2HBJoBzOI9tLJWw0o7p
I/1G4aTL2vqmIasbpH0Sxd1S/m9v7oGkzl/IQnWdxNRDtJETcY7WvliYYX29mFu7
YKI1FmaObWJ4eUqQR1mR9umQCDRx+lgpzREjQbu84BHWjPbnmFZTiFP45mWqMfzI
l9aLmrhvTeB8PcLAw7ectmnkkg/FKjln6MKdmQJ2QXRHaEqjhjqhqo4XdP6kBcVc
IMqX0oznwpnWxTKhg13/eord7x1hjdlV9mhtG01UXbcgDZ90pxXBn60ScX5okdZX
Ze5v6XQujuu9KUd+Lm3tUw6+wdB4rDHHRsah4foI91cGizskOHk9I5ejLbHPJY/h
dWXT1nvI+PY0MIa/7YIoO9dR43o2teJyfhN92/vKeKr6Qz/ec8HOnpH6p/qU4wxG
+CjrSmCjpbWNcxAopZ8p+A71jIQcYsBTEwls+A7Utbmt4BML8uEU4zOXoVtbl8FY
1NTVHFzpTWYwgY4+rS7Q0I3nEAwS1b7QF7oe+BTLayhiejR7WRrv2IPUWnkU0ZI6
wIIWeysjmZqUSWvTuTaXduFuqq9OvKUfQ5j5M3J9cZBpzLVJpuYrkjv7Aaml/wgP
JTK+XBn1iorknD62P731Ea6nKfcp6JiH2MfshEaTHyHFtMCMB/FwV8PnbPvKQAc2
0z4a6Wq3UTH3u7J9NNRcVei2oNGc+nUU3CPZBgzh0awD5gpKuKE3H36hCobNOkS0
7h+Xnu/D+wzQ1DQhIkL+N9/NOaFzn8x0cq2lnyIg4sHzXAnMWym73evPfoCMhixu
hyL65aLigqoPCC+xtbaFhK9YqHoSFc77xe0kt+CSlH1FdBv7+KlXb55GUR3QO/CK
KxHmL7ax0F8cTrVi54to5+EcyJfSPMNfBzw0BwUMF9de8uqJqN9iCGsMk1mJtbOh
FWxOsYXvYzzKYxx0MEDnd+FXtqM+gYBnAQZYfVaxicwF8v3WHrpfsFBKvA/O9/nc
htNu8PJ/8zIpek6hKmLILA4tTQxW7XWda0VakdHnF4n9pVUF/lo+44cdSAhoYIRm
pEk3UoCsvBaCBmHipOR8GYAMw3sH2RmVmz5Qtp6semDVUJNkbxpfmJYyH+71fWmf
h/h6wtjD2Nv6x4IE539d5pCI62dLG3R3NO1AwcoiUItpeVndHDXNPU6xhZZXKf3k
MfYUIzjKHMFyDR4Y9FdcIkFlzmL5FfWXOMMD3w6twiQwxvAs9yDw6SCG3VMvY0Wp
UPVtJqnsudD5NxJ2zo5cO/Ud249xJTpvsAZbbkD43CoG25PMjvpGkHZxyLCG2xa5
vXXBRCwOepn35oyIo4PDn/bcEbZwMSIxyV5mq+zl45qg/680GDQTc8dPZZMWw/v/
8n4rSHQNJ6NKUsVRQ0oyHapr700KtaeC3hT8lIzr+72ZKQDZqrniCppgqMBXtB55
oDxwPVF5lY57AzWMZ9HPMGYy4hfqdHf10Q0hr7cab8qpWNejNg3qgEvDPUSTL72d
r7iJ1LMlMqX/12uaB8GzT6+yak79R6ozuSjT01mNPN1AnO+fpFaSLd4RtviebFis
ARjv2s6XWjDLxcckSO3oqltvDh3jBHbRwnGZ7UaNJY6mnobZruUEagSeNvwrWIdu
BkGdNiHGNy5b6HB29MbeKSliE/sGGeGcCAHb1D2bSyhQystbYKI4IQ+hlONBcCGK
mPXCICC3dt7FgOBLIOLcPxnfprlmtoTcgXFi66T+WuZnBEObg+iavPq1IrW5IAAH
nEXIifvjlRYRgIixBguUEg3Mu53IDfpWWjUNgyMXwFVjo3IWJ1m0oiHnm7YJC7lt
nT6e1QbyMeZcOpVsCB/YFWZm9PoyPSIZhhdGyPiCm1POqT8yA9oCyEsx/4GG0uqM
Jemh1/wbPKGxAzzvUp3sXL2UwMXbIob2a5FYsOGXZ5VhK77PlnsNfDiZo2ohGJwu
gzYqrlm8dnfCGINmK7P776XsVauUJNCojNuyERPco06hr9tQp3BoypDoINzs3q7O
saT0+xiVRY70gtMyIBuYHOTo8xK9VFux0feQ/sQeGkuS3HqIdq0yb/tXaqzSscGi
2j/o0ZbZGkNwn2eQRfRbSze/tjSGgiAoaNV4f/gyp90g9bksfdZivKL2elCB5kZB
T1CV8OFrtdrnAdWrunfZXjr8N0MCbDyzeemwJg+bJu6dLuGkJpNdNWTEoyj+6vmt
YCpFKlY1FNr9iXc3WFrgJ+bREt313OCFAHGrDBNfji3p5Kl7sem6/T3VTEvXs9RA
UULF2ih05PR6UFJBEhOQyWJ8YXYwKOLMt3DJp8d5Fky2QrDzGvEeonvWLjy3ehgX
2+OtxANzhVTHfVEljsAUeVYM2qieiXivl8pBErGnc9eNokPaEexfxifmvPzqNh14
Ux3TY5IFW+xoBgIpbewGsnSGGOCZh9LcGi+cr/nCZ345HYlaYtj+L3dtS/qpeDvm
Gm7zxP91I3Y1RJXnPdvAre7qFD54xLsf7FXPGWAwyKqmsldWJGEK6qN5/wnH+Dpn
tB0gsaHFFmyMXBj1MvCEb5MB44L/i7leYGjPtPN2unPyok9/aiWLDgdpoJaR4Iso
RL3N1JSacCeUJ7i+xniVzD39dwmc+anC6WAeeKcOIscIQ9iSlQXaphElTKajnoQD
Av3ZO+xm2mnppfj588W2kysBYQrYi04hQgpf+jBIlP04ceJJnh1YfSHVT+91RVtp
0WgYAQcTWaHsRm8rWwdtkNvPMUbYRz4tP1palMSONF4Q/31eo1Zg/WQSdfcCZc01
vxmk9dc+McJBfrKBnkcW3mE1IwGzxESGBMKcHTdOJ5jBNsKxgFvuv//mGXrFYc6A
RGbGYBH0AlWqkvw9Nrrqne3s/W0gKfnpGvsC4lv+9Y2C988ppCJGBvNKZaKSO3pH
Cy0EeVmmayztSa0S1Zm0le0r0tg7COtVc4H3jxTXimTVDczMBK0+VEUNKw2+sJR4
pP+fIpEuALRGSfRFqAuAvCG70H9tW+y5hZ7ZkT1k9PMNH5yxHI3o0BfynoBLbUKI
etS3hcNGajTva1TWLaLqmNgZvs51TPiMDgM6+K4DFRtPxrxBP0UjD6nQr691Qa1E
zMX0j+nPI+w8r9yf7fnd35mcmAn/YDDDoMEH6AimkS/F9e81AlPU7qNLXuNGkfm6
CwtiYBHydGtT7jzst08FKvupsNXDco6/akjsqYS1AmN5AIqa0Pf/3jOl3+55kXAH
2rWAYNd+/uWnu4CqWf7iEs2esqZCaMmyDqXKkL9eMsx5nI+1esJQOh6DYQlETkTX
PzIxk8B1g6iNmc1sjaxwDbkjtoSjb7mtnKcH4eLlOPIIY1HvOaqXcpzzoFuVLymP
vPAMityBhYVwyPYc9aAPfo5bRcuZS/dxuwqX+mwCbFZvmqQNjHooch6S3WEsuRdt
1XRlbdQKvOB78f/g248C8uRFejcCv+g6f6fkYndyboVp4cL9LPXkK2Il+3b8EhFh
0tDruYcjodTLRbuo5JSoGuHvL1U/zEIRlXEgL/ioqtRST6fO+159sa+iKdhMX88S
3K7P6SVveDJDWXrmgvpEbhW5ZUE566UE+h4x83X/2OWAM7wDOyty2GI5KBdnaE6o
HLkqNIrVENGWd+jFQs/WtZStX/BjzXi8jsJhVD388/eq/HLY2LHvdESNYHQks3Fu
dlYn/u0c8NgjWiNKNKS3I3Sg+OPCCNbhijvyygP3CHMdLG3X1568ZCqdQf4jvRxL
+V5KqmOoA1Pu6WmY1BzVzhaWVoWqWnwe8QkQ3Fg5L0yzvFGbokjArOouDh0m+E3k
o+vxEqrjhxvRMRMCSRwjPRFXAs18/GXebO0mckDP41NCJE8JelMmLJLRSeqhxdyc
kyUkgVch7heiI/Z7g3SNYgWUi6kYid9xE7Ijn8n9lX4TOBv+lnmxVAEMIKtnTDd+
7iZwXWismBfDF1tnKh7VJFxRJKr9+wxJV6TVTXMzb6evAyySrI00y6WNJgYoj9XC
7ube1uILvGGnuzEjUftZWcajmpyP6+nziPhlkOIYxjbK9tngS4Ttmk7sDM1qBbIn
9JOP50rBQzei+y+TY1Hquq75EcVAeH9tlWaq7ITh7tWXofhLEsKGB3ykCC9DwQbd
7THAIn6A4pilAI9EhrPzwghoiNZF8peDyd2EWPeTMrKVowdp66uwr12p8keua+sH
3QkU81CQ/HR0l4rSnJ7dq2SpQFFkatC+2rh2+cYD61bp/qHLDBx9tl3SNzBj50rS
OI53EwgHdPpBEvaL47N4t3iX2fqLl7KRvnCUs5NXJwMBnVr1zKv22vNWr8owvn21
YvhqT/07S9DXtrpGLlWZbZvYyWoN3xhNWS48oPdlpvPb9aNBang6GnVOThUZI+F6
VLHi8jRyo4cXedcGIEg0hY+OAnpHUON7aap14tS0MXrn++HuLF5U/NrTKl4WFh2M
KgYMlbMsOWI+DdhE51nypVayPYJs96xDrrcKVQv56e0Ej6IJA7Fhz8qbDOSz7RuO
LNbxsrRmitxHgqwPIR8GOw5uPBA29Dpe0t5aZRY/vbIWO5AjCb30GNQLKxCMZKTL
OdsBck8u2WbvySclhgDeI5sXMvu/Xt3h1ptWV87/qnWoF5P+C8hdBZdBcqmhqepF
zziOycV7ZbxNk+retVSHd5rDBibrsbNfC+uzghwDEOFjC1q+56+v0av85wFfw00T
zJYKkNtA0oRcWX3PbKN5TP+D1MCFYdla1rhV4ccxwq5li4as9hOC9dgGiNL9FcN3
IaaOdagzUjp/eLrbJSjOKSe0YHTC2WPXIf/BSm/MZLmy28SnOUAOjY2WPgDMYIoJ
dgBB7WpsH+uPvhpkahF3MS5HaWMpBBtqoplb0DCOAAaLP3qsMZM8t+sb42Y//sP+
mdZAWS9TX+EKawHjo5jNudgNr+cQLxRgsDIemB3xOouWLpxZQDkL+laLQluIJaCz
BsgLKHi4ZlnBxw0Abp4XmCHa4H/wFIPOtVuvyDTQLZxQoi3HwUPzPv/Vdyn56RGW
pTWf15Qo5JrJVx/86Dp++13wDSUgAh6W9EgH6cJo6pNmTiyYkwRsp8nHcgaY6Zsl
gkz0cZbTfTRY+9VnKMRqvRB/mRqn5uD96+g8MMRI45yJfSZz9vNR0Yb9zSVg7jOe
T6P0/vNfoVilYYVcDnaHyJCgGKCpspoNKcoqWeuA9u982Y9nYJsU4KmnlaBY2aUT
wBkY5zylPK462tdMSDzBKUneWtwV1Fo6AwwQELuAFT7nt1sSJNw2tGXeHBUMpORt
u00iDSP+EaU3uU73v5ezhGcePrfYc70WeQ/SEKGbFRH7tcMN9feL6urTG8lfdDGM
HGEpCqw6eON7fSAo1HCzbz2tQ5RQJlvG20TIEQI346SaX2wPOW8pgUOXeWjeqqOo
ij7xVfUdKDDmtJEdwFfeKAg+P34/ktkm5FwQnV6OM6SFs0uJHbxkEKHnRkFShRKy
PGt1Qbsozdi5AtFmT4wsEpBGC1B6b4euiqx4XowqCah7s+gnFU0s+me4ye3sCATY
oa62ZFlJPupWVeXm5nRYZyFEJrUmU59PIzAV20+iqUWuaHmZu7cD3HkvvYjK08Gn
osI1IuZUDGNyLPxYkWnxxx72GA+NcGmS9g8oBKpTAxgN3Fdstrt9plc8NW2Xm96B
jxPTyAwcPokK2QyudXXUo0HFYlX0saMDj/ZnH08+EtEQLX/oqZlSHiWbTLZVakCm
nMXajnpOe25+VAUanSna5lFwg/VbFDUvdKjsN6TN/F9i4eLnOlW8cSpRdifszAhO
JE9ZsWiLsUuxZ+/yqkNFGNf3rtfD8Iwuu0K7qT++ZsqktmbdZIScM2qDXy7vLLFA
3EAln7t9NrKTKVKKgGTmDfZXey3wHse4ZRcfNKyo9fJr8rreSm4KCOam1/fzuS1o
4IN5t+5fuaQOIQcYuk5IwkUU6ayo/KHx/thMTKcZ5JkvBK5iq+3ay7h/yFJCFvpE
K3D38ZVFeis6BPKA3rIOqpT5OCocRkHd8ldzVM5cCRJBgMO5LFy+cgo3RCwDJ8rn
YIrwXnO/S7QmDMIrSQREQF0Q4jikS0GLowkT5kOhLHHAbl/XzkCiNEPcl3I0dzUL
m54hz5D6VFdlV2R1jQ+UsbtGMMZU8CGaok5YhzSq4g1Ne62sEnRXlWcP08NDHhSm
wwyCbvKbbYIg5WSRH/312GjAd5Hc0ZuWY2DEwtslPkTGi5qUpjnBEX3kfvh5tlV0
zclsjQjAEKP79XBOU2bysCYPCwXt3vY0dmNgNYN7KHO5C0MNnUIQnrAQPXiy9dt1
CVbKvQzWOPKkLYTkEU4LtwKwqNFeEWPbPz1QcxOO9pzc1kBIKU8QnkBwl/RrbBSF
9Rdz/0d8lElfhWcTEXqgyp5Mt/9rMeoH7n5WNl4nYs4ClEWTkSYIg5N9z4RSiiKC
pOP8SXpMr3IYxsbaGLw2bjR4GjNi/RGRNugIUndV8JBnII8huHfQ1mMtzGWYQkyO
4zD3w94h1aSujYfpF+B6puPMJ8AP8i0O5DlPIFnCXRh+XvM9kJa8hDD/YLV/1FnT
A0RN+iJjJ45bYLC/Uglx1ZBNIOM0yHB0Mw45kYcxAwH42vBIGcZZ3yyIyJdBBvY+
x6CyGfurDFoEZKiLkLbcK73YTjXv5h0AR6rXJ6wZygwYndU7/e4vyXCk1dDx9Y5W
b3edJ2XTmd1L/PLfnSFLhOIn+P79eml55g8ha1UvwEwWMrv0De+JcbD5cK4EdgbN
lhL7XBJ1V4M+srpg+NNnjM41uTkJX/dkT+efeXb0ioC4fMLzC28F22LNkQhHoIET
BczomiF5zucXsL9Opa9573jS/7adW2IwFz9E0pVvhkU1I4+V0YBSX8+5qwW/sMad
NS334/srcwi4J9ZGpr5NbD9vqUj1xFjfeaPof4+r60e6gxehkiBS9/ROxUVLijlf
UEk84Hi4CzV9hHTnM96ubAQV8Fw6qLDtvlbC/BvYGX+FlWzvm6WRAdYrbvvN1PlA
+om5HBXfPP6AyVPnDhhcxCdrzIgiKBdBJt9C5uBPkAiORjYcOJTBH9HAR4w2ElQ1
es8a3mxyXi7FzINfLpQDos2sGjRWygqTKRZh5FVh5c2C0Mk/zkDSIzkc5beu64Hi
AzKV4LaFglN+4swX5dU7HdpAWZBRirjiZbi2M//lWl2rZD2MS0Vh4B2lEN8dn7FY
qaF5H+7a4YH97ELejnQCv0fF4mscaIKDZ/7WzE/Xb34twmBcyMGCZQALUA6fb5cN
mYB2TZKNYWE6S4dA0ZGKr4aJT5T3HvhpjwKapehUpOpYCwpecZ6fIqETivpd67LY
YBc2AUI4Fa+7yr8/Du94VwZL0aeG/bbYifnjIXvZhQ3Uy2ctS+Jd0ppx6A8+qUU4
CJBKm//s62LhpV45z9Zd+JNgzl//oEJwIN8l5+pVh3TCe0ojyB5LWyILIEWv5YgB
aPC4Vz5SpxvHRvxzWXZm4hn9JjDR+EzntU3iyeqNtVViBJTaGXkks4r6M1muzzuG
4dqFSVYtCZw0JP9Nb/+5cdvcem0ilKVlBi/0RrkUDeunInFe9G3TnWI4QySPC3sQ
MUiSUeAJT4qgpbeH25Iy1M99zkQO0n5KC7lsRKL2HAlfnvwgF/paGvQO/+XuFgDb
oWL+ZpV5NHklgQhwets9qZRwRRwdtr8n4n99L4MaQmz3v20dvTo14ip+jYofU99d
oYCZ5mCfJ2EMjaCVgMbyMsg3fUQtx6I3IHfwACYIE2rPvGLOpFUyAyL539ses+sV
/+1rvzreDbBtMgdJ5w7GLoXob0OuXMH3cTVgkHVSkPhdaL6M8DXnl2EmmAl6Mb6O
jid0SUDoEu6pDlNvwQ0M5MIh/9ycaC233f1/F7XWkiKwN115EwQCrHVO/qvoRNuQ
VmqSn0OauWID6FkdtwiYexHt57gEF4TDQUhlhnQnJa0SAgiwFN+ZtSn8sE9hN+no
krEzSHv+eVkCxIVDB5oWC4HZxreTYqbMrSXGnQxpYrhNXrchltbASFvXkoeKoyxR
fPPkqeJbAeS57b+xtSMAd8EsbPu1jQpUkQIanynjAuAj9v1kKCLyslCFCg7wmTI5
Pb7GUcBt4Nk/xm5Z1H1hx0jfrQk2GOWZrsZCCH184mUB8FelJKE/Im8Dsl2yKABv
1aHPJpLPo7RUZ3oAhPWTOsWxyWfPcrF1y5qqXyJbhCMIse3M748eXw+wXjaxkqW6
4OLRAykRdR9NNSnDkD+owMEtsEyrgK9UNz/pvsvYqhDeYkrUe/XRvfIyTfqLDqOD
9OsH66pdk9PpH//UfFf9DFRpdnys2sqoJIFrVqPuBr9IrxOwkNSWwSd78HhDMX6E
HZ7eNIv0LITnuIGnryLDcQgglTICsXTA9uZB821jStJUxA5BS2CZDPBL0YNvBKLH
mD4t8hxpFSSESgGIJXpV/2CJUxPl0YUvNwO0DeEw2p1bOHWUqssLL6WkhZb+g42o
xRwe7oT6+ZYc7Lr/HgDQbAq97fNQV3MZYvOzifArXzq/gzAyQtOoO98udKvtfGV8
Axrhg3XfsF4emSBzhqX2eEcmRnqL6vJ+hWrdGG6cCmyvPRhoq4ckwV4XnOuFyV9G
fXok0rrNERXuKFcozC4fqprnwtqG16mYlpUHs1wNTFch7mEQC6PrcmhtthovCORv
vcMweAWw0CTq8LPQjzU78xM7qAFQguXV4CKWMoWri/k3vUQln8uc+aUjn9jC4kd1
CT9pCvxtMq0HkyDxDScaSQwWK95X8Obxii+EI00CXT/u/+l0SWdHgNd9U3GBWJuF
+i4vsyYInYFYpS5XsD2IYpXve37V+gnJ0rVb538f1AQgb6mto16tzOGsghcn1I8r
hJ2KyszTRvT/SUH5Sz5xe9hdt+5SKFI1jd+7NmGgloE+KOuzbHoV+jzQZPb19tGh
gFgZgfRy00k3T9yu+1gGbp+zxLoTUjNrf3C8KEGzTeaRAw58dcgR4ImTyaae9Kad
gKTaJQa0vsvqCTiQimjwTC/7cddpNXrt+LF5PxO/IOZlO7Spon9bTPunPVbtJv1j
1Yns+u9UdSGcZgbOrISEqC12oVDjYkvbudABefQyK2VsOytLGrfAaA+kZFaoVpn5
vI/70CgfnHq+1XwVA6ApcYNvd6qW3DNoZyUI0jLHkg0GNlKON8Z0kUaUR79iO2N8
b/qz+4Dazc8E85fUz9zXqaqLk+IcRDGaylhwvNrGJofEOScUJyGYj3+0Mjl/y+gj
7peMx8juCZEwbKK3TNDHXSa1XMU8+Vmg5OpCPUUWg/ZPyiLlotNr04tIez+3qux/
MhM2OmZ2O8rej1MaA4pBarySm9St7kgn0FPqVGKgPbCVcxp5ZeJ1gqgXkzPbwJSQ
sPLzfbXazwFZ6mTEN7qeza2EnHp9+5R+xv4Yjzc68jc7zZuyDlXkjYfkU2f61azT
cS/HH0X+zmXzarrNsdNodVzlDARubmd2uyz+DTQhExVQ75+eZEnWKbqq6hjrmqtu
bA4+x+H326sSgigI4irMB3hcdSlCF7R1/cFBaB1f3Ph7gnrFOR81hpb/fEU4pNrB
XHq7ANb3Ql9VzQwxEvt6g47Nyta9VZrKg7uaOZTMyc4X8L9BX8atLlP65FbLyGTa
DZJsscYHy81GrXTjYPEcxp8ieLWW9tsHkrD7v5LkKoLZyp6iL5gt96JZE+dK2DXZ
4+EeC2EmO2/RsBNkr+SG6mUt+AeJGcmDh/Pnn1phQ6gzgHQIjPc0dnSFd7k2Kg2N
A10WcZCygvug6qPcH1gBUZTADcFQh0eXBJrfzEmBi1MwPmnqS1Givzg4wBOk4byY
FBUyv0xJKLTWPxGquoCkbQI/vRaywnVsWaciJN0QLvOUTFRiNPdlGUP0xLdFhTv2
SbnHG4yAto3y7POOWMXskbiG4TpYK8cwoVKBau8EVIEGlZeV9yxwLZcQAZBOBeCP
ZbA6Ym6mBN68lTHwywk6AXCJN1g7JEMbUEWVpKDKvKn/rAhVmBfgEHeoQlEnRhkp
4+zGm8rRwJx9MeIkKqV5yVBX/v+dFZPNah+REFGJeWda+pcaB/cewdDGl4d0qnwh
Drwja90FwVJUsfCsoFC8ZBgGPGhlLot/7sTSKsl9nY/e+KHlpPj8+xZYmbBddaVp
noE2v40FRuZWjsBqTHmezgpDJhmKLGLAjKmPjnQkKeUala9b21+SCK9D+ZnB1FFt
F8w8NgJgUMChcYKebb1kCYQnTtyE3SB3dyLvpfn8dNVb3qAISfi51vOGRi401qMl
fdxbDwXhJUteD+4fgIEJpW4BS0vWWsbf/DKvH2X1/Bo/TkFtbhNj4UnDph5rSsCF
b7En5RpIg5yykCvMQDe1HQGdyZRwIDdr3RuLGMssVS46DaM80Josu+4ZAJG3y0wa
yAOmfp5d362264/L56Wx/frM2HZtws8bHeyycakm/tzNtTaZdL5KH65/QbLgYPPT
mZ0WOg3Alwhe9Fo4+XR2vdG+t2N1E9P9mYS/AtCFrzjr2PD4MC9l6H3m79ct8MPt
8FdwbUrSoyqwdvTwHOvL4pAJzR/Nm/jSVY9Aj5u3+UFcgC5C//MH2bGvMl0NbdPS
/jJXouTk58kgP4Q6J+2Iw/ygrWFopaTQlQn67Vnza6fcQlj/7ymYWdsXGz4FtA/0
szPK+RYUE9/tBgQEZcCjwyE8AsWZZuER/rvbTTNF9IGIczwae2JA37ixVF7W7GiC
h0kArqraz0MQdXYxhdX2LHN4WIymvJXnHe2E6NpmyF03IjzLViyYQjBuUWI8IzXT
2apjDpii3uEXQ63b4oVvjXigj+mWcG0m9jUeqasH2jIxeKxBn9M53kdT63uyRgXm
nUTa9PbCfly8TXcMWh127dT2BZSPt6ENUuAWIWUxCFI991oG4uQ4lD82HLjamrLO
PgWhp05kv5Rn4nCDQqMgaE5NwTWOWferdmnpSTZFPTw13MSf089hcWxqviZdnWAq
pg2D/KXAu7ymI0N6aZOcVJgsivgxzTn9xANQ8TfKrct3N37iofqQ+yZC6GTKQXX6
l7DeuNmxvlymSZQzBxsV/7rXzrj02gXbvH/lKC6Gm6As043KVqU3UBw78vwCZsiC
JTvYtWL5x97CVbYfSoDC0EKCrtDwTGyXN1/Hs1lbkNDgnS5gMEPfdeiRY3bDcxyl
8sb1NvOWvGcO4umDhwG1S5R8ihhiMuBkH/7dJElg1WMyKWXOfTQ7rTxVCC5+vG28
rP7TCfvnB2rXN6SZxcgc5wZf5ItmuBfTNTbeP3lk1k19FueHyJytxBiWMUf2SNAf
duBB0Ls5GoetkWCr2R6uqruoGUI0HdMywjUwxfGDgIRgs3etk2XrxNJL8iTjKNHE
OBSljcNL589vkfxq8QifuduNGqdGSDVXiZxoCsKS6GYdIGGShONCbB08E3iKkhji
ELMtpcccn8nge4AN3lzc8MDe5+X0fFwkeUtcuUSJxP5nWhh3+9GkEQBMH+zD+Nsg
74Uof+xbtb+6on6SDLownm4HXe8865f2BCoOPwLf3NIzfBc5fBbz0gF21pQiuqMW
I9wW/24ND12SQFNdLAgVZSO1GkRvmHB8VHh7jDjRCF9qtwWtUV24b8ZAP8ZeW+9s
CObizDlAe3m17jp7GGtcpOD/TrIbV3/1NC4GiY3kdKHqhJTjozIXs/Z7WGWg5dql
4GhNJivmpdsQsJQA4sWQCBjCbYX5qwRmpvYTA1M5LDhKQ8uS8F6L4BsBM4+gjwzd
u0oLpgehzcCPljO87ZUO9pHNOOPvFEEphmdk7p2VwBhBP2RCwsUm0eLL9NSWdECZ
sexRRw/ZsXZr7ZfP9h72EkkvOXggtIF4fX29EUNswFH7I5N/4+I7wOpZcmjYPJ5F
UYrBhzxX1WS6b6P/VT2HYMaqq3RboQZhS21zpz0mDQ7GLITmEhGiDSIS3UKXf4MU
aTbim3HHZl6PrnW+6Y4PoFz+SusGPS5tUedkPA5HDiiPlIY3LIaXHKbz9R2Tsz4x
ilul8nDB574bE4HBRTTV5oqjwWeJGoJ5Lyhp2eoHaaR0GfYpwYreTpUEZ8rr+sAV
6iLLr9L83+UMYOfPo1ZW9J1MvJDJLX0pzkmaN2p1gTSJY4hNRK4wefs56uV4xqLJ
VTU/uzjfR0xPB0VfQxMvZ5/Yzhw5HHX3sFD1H/oNRoppB0hbEzvbFkqhMFFOoQlc
XV5Zj+g9YhRFaG6s0GuFZOwVOS2ElLu1cniVdvYl+PC0PwpcXK90/5UGMGwoXmzU
pDBy+F9DVkEXr6FfIZmVcGLdcNZJTtZEt5h55etkE0IHXdq3fOk9x/IEPBQmo1fy
9aeXr2R045MumrfMXWO+8JMtGcEydiIrDyXzL1jNyzCYp/M4V4spwmXzu8D63/wT
lStIveHXUwVPaZVv/pMeH3Yr1BqnIvcaLwjhdU4AuzDSVlgRdrrR+6nwNn5t8oqm
G4c6CklGN7oQD/j0LcAsus6oZxi7LVfxxmVNVSOreADWS8uxFA9qp6f+ZCVwvSfY
48Qn5O1IXANguL4yPfzoqikGxOyi3eo72A9gyjqDamBYE+DB6e0QbdwRyvM/hqkV
DvPqwsn/Y76TsseLNTUolUH42U7T2FeRWiJU39QHpKvbsARh+BRSkf8O2sFoDUTX
FPd2LSci7h92/RMrTnkHlcIEot4Aq7NkDtNcRpvn02boCbTYEvWwFaZ/r+foReTY
+gfBxRvboTAk8Y1eSWaw/3Dg++gk0/dSW3UE7+6eEbkoA++/sebYzaG31yFe8JRb
4coZsRGpzCenuA2kYG8G0C8752KGMKfh1ZpMLAxHxIQrOYqsefhIpZnSoy3LpGzM
QZuSpdsWNYnfJzgK5RFiSS/+EpuLwxJhZD03nZs3EzYfgtxx/m6T1QXKnQmJdUkd
A6FC5jy0pZy8f2vhxSBhFbdqyPTtIabHurwcehB5ZaFiJnaIdgeCzH2jhJxis/SE
NHqx92wnKv7V4iiWoe0nyBQ8xN5edG4nh9Rr5AVlOk1kL/rYhnNryRzgLyl+rNYE
74M5exXckyXIsaabv7BlprzIgT+LO3koO9ePhz1fGK8ctxhWDZslnoOVNh078N92
rCLvItlHY7xYWJa2//8YWHil7vQaUoGw7AGF48xFY5Gz8N4WBI2JRGRPI9i0kQzt
wIOgi14zECX5YMNQFbl15enVuOyMKuEjwSUm0sR7ozJOvWIzCPcWJTPhLnwiNe72
j+rpzOo09J4GD5mCpdy8RrHq5cERZiBHfLNUJdwWVbzYpouD9kw2NuCUGptBESP4
MENebiyWKgcchd79Vub25VE9RU1HKcwNEFNdyExZea7lOnZI6ziZNSCXixfXexBb
ajT7qdfUgKTf3hvxnFUo+YoOyPMS9faBkpgcCbGbkhOlU3Ig7pDQHSago8LFXrlX
88FEh6i5em/tnddpIm18as3AOWijSdjCTQpHtjfj3riDfynpROms0rbIlBspBNmp
En4HUfXS635Kf157h2Tdjzs4m/xVTj+0lnLT07sSacCxqG9Rww23uX/pa84zUaF1
l3Hd7Vwx52q/xiMTINWqzkMRuS5bCbWS5ip5aJrg7yzioZfWylTDWXaE+SL8wSUU
r8gtp6pw+yMLuujQv1ZjYVXgRZkWgO2XJkDz/fMCD3x97Eytl3t+Sw//F+QRibRN
iwZp2tWSfHWzKhSZg145sIkCZXfcdeNwTRS2X22tlEsi7qPlLghKZclmaRUb+U5C
BifYQ3/bMdb3sTXBLiNZfHmwxCg+2asMwfajgOW+4YKphQ0jad+wGXA2yHbUsLCx
8SlRaj+NrjSjcOtleHye1/E0jQVwOX4MIcjIVpREv+C2Gb+VZapEKFB7wGV9LpHw
7/xf5+DvEnq+hwormldfSctvS9aQ/hyZlqT26P0tmP4SKTlIunGE9UoeRelYY4yo
MRDxmKZalxTQXTYX7ZmkKqts9MSU+kQHtx5+ND6xjhAovn26flRUkOFwyDfAYXDl
6Ip3snRNglXgQK/MiD/Q0ERWJniEjVjCzbm7wLh3/O4nUGvGw9xXOatGQOXlOD/e
LEQlfQyOht8dv93dS1EP0nMfFzqcvUdRKpuTKRE/YtFUH77VWiCFyKLVGsxbkJJQ
chLiYO/rQs0m1gDtxgWbOU5CVnwDseqBe67GVUOsZYnFEXvpQbuWFqDkvLcg09p0
WTD7Pgm22Gt0ZgpTlWhhlr8OTnJoVEL8nzPhJ9kzFdlbJL3KLJxQ1X+DbgD2ED3T
OXFRjRl42aQ+20XFoQDk6XAGar1CXNX3XZ4ECsVREG22L7O0XYSrvfYFdCKqoZK1
eRudoEvB4rI1TTkzcE8URJMnt5b7nfunk2mLiz0MLrxLFzWi3IpAyD0abF/EJoTA
zuKpx8JpB6SXdp7Wg5sAFLUxVgTqTTGcTFyI7hZhS/VMm4F8AB5CmqM1b9xozwyc
6TvMZK7GAceCRc2SyvJlW2HvlCqGXTJTeojS09cYFRBw4D61IZUCrK+EbqFMhzLB
uPwtnT3XZVOQq6jdu9oU+GFHOaT0wnS43jA6cuzUWIf1YGDkPineQ7SEWYwnszY6
5nP0BGMr3NQBu5BheC78mU5D2pxw+n08tJwumhmJRshVLouDyCOqvNO+HlnYQpOW
R4GmesSEynbEbDo5W+pcn+ZTkVoWWExHWWk4j4x1a3V1FJS0d10gCfzkOGaxVjD7
q8P+iZdjhBSI6bUa/7gN6RcoVIu3N1yEdCbCxVkkIhWsUS/8kMuM0yJ2FnpnvlKV
0icEm/o0i2TYR7tTOl4qUXUvn45ttZnVeTX+ld5/l3Nvh/c4L/ESnXftCj1Fezdg
uVR/VuHBtiXeGd3TMn5cq9O92QPPet0xMeFYD/el2aCOM1XiqWccP7o2fO4ey1po
ht6yhOS0jCSEiAL+vci6d+bwJaDTEenYUQXqWPiLx/eeMO7f8baiveZ8PcMHr1um
HUZ8wHNIrOBzpiVBnZgupUh+sDpzn0Lg+d60/JobDn8t2jJwqDUiopLS2avhwibt
JYu6Vxuv8VX4BjyNvTVjXjhBRIXrHbbM0t/rXd2ELLwOimKR8Et5i6YS6jYeeRtN
xzY2MWdVosAeJYZlM3Bo6e8At98OayRrP9eNhMAM9VYhLlQl8ZYRZ8wAVqhs3T6e
y4wYY1+b6G95dh9Xp4K+HmjEIIGUMaM3HSBNaPZ54zofHAnS1BqjXGTbXNXyQxvX
chWpQhT44ooKQaui+1yVRHDlRulUxUqqdyoczX68XU1yO9TGTScxycas1aXnTiEh
7AK1hLPDVUP6yE9m2S7jsD1mEpm7aTCDevTCSaFsnXKxCcKiQ8BwLWw0SYBZ5EH6
pSX+oTY7zx8ZWE0eapQ1X6UpDL540LtWV2IQbskSXPS2qn/E9aet+/BbRO8CMSvg
Nf6QW69oefigMyLB+XtLZkv+qOg6L2O3NHaWcenr3k1qeNN4fZ2hkdN0jZdHGnQw
ysM+VeE41kEuZeIynABiTdLQAHmzmcsAOSv7YLSF1fOk2aBoK9BZWfrGP+KUi4pU
Kb7CSpmUli4jD/rqe4EGlMYFWN5vBTmn2JmWeUtAQUjopWfZKcsnOsiAn0IDF5BY
Mn0wCizniN/fDrNb9D/od37Epw0WdGMat0moNOsys2jARaHonK1iK9BuFCKbcyL0
cQuF+aNgKkdd3sV25VCcWo5SgmkgSb9wyEs5mSrLWWLf/5O/LOHYprCD2XXKM7/n
IYazLwBqUwMw3PUfb3Ni6MnUGTDLpd9z6VlfCFBKbtCkU/jyk3zHX0usUi/3JD5D
VWkIYrgJgnBBpUIzwFf+8VnyyZ3lnKby6N4zw9geQD5plCTPPNXRPa/6pqTinVFw
pMFfCt+nL/tYeT11mAKPYpMTaXt12imrrzWGlsoPz9dk2Yi/cWXPhoLvELWGZ7oD
zB4hE+45g0iyQBYLv+3SKarkWKlf92vIoEZq1A8yQyNRSMuu5G9anGHxhoPJxShh
jJ61HqqDWYwiWCLb+4aDVoMdua5kPf7qexaPVe3VjbWhvi3i+HtM+ctWeKqhF3ar
BPcm2TieG85Rmtdw4Q7K4bHCOR9uaSjmC4WrAuwnoVfRRTG/jJhk2+38xgNjjzM/
WSL/hgWIijzERGEsW5G0mG5PXUCQaBFwQ9XqCCxheYAbR82mdEb2SfoY0G/2mhNT
plgSflQrJz5Xqu2BbhYYdaCfijrfs2CkCkHvc/z8mPY000soRpqVa9ejKOd6g0/C
ONuoesTx0A9EnVAJX1v3NA9duuk1W6p0IMDz2Dg67a+zPGbfdyJYFv0eUmXsbrSO
NpeJLd2QtdypbmeJ/SU5u76813TYTh6tpeMH9glwEh4bWbJWouW3bRP4SQrnkUCj
71W/BG51kgYKy+BHOD4GSEWJqeiXKO/QyP5/ftC6w4yyKwHykqvdJxG0Sgj/grLg
MggnbIUy47KKhcIQwWlVjtoveVYAAZkEmnv7fys0GN+f9xe1WfbJ4G7mm90lqy00
4wlzcz6RyuvKTk1h8Anes5rzjH2jdM+PC/xraqoI80s2sxiYoB9uzSqWvgYw9Bc3
6kzJBDrrkhP053UQ79PEWRWzASsfDzVIHHX0yqlVEkOKIzOr7Nq9V2cOsrvxBGi5
IqShMRX1b2THaYplS4bg6AkyxhgFSW5HtXDhgL+tThLeMsVkpveiiNmp6ndL4vli
z9oi8qT40G19yKyMLMikbk+gkeVRD3E/rdxDYQ/E4W6p8c2x6VeQR9EnlDY/usld
ORezCPIauaVJGQJVm+jbeqplqudVpoqmW0jrUs0GQNh8yIqq0RaCvZFG8VzdGGXN
6WYhVdQ6SLiHBhpTmR5CT7r94waWQjwcgbcfNJ1eG+teiMolildIKRW9zDd+P7iw
Et9cLiOVcXAlYlmXKIAwqSG/wTm2fdwQfebc+f/9GT4lPsetUj2TDKN9CaSwPpLe
rdxoPetnuzg9a9wU2FyF75FJPjbhNPBE8bl4RzBuTkxQFpAwiK1UnqBjhyzP24Oa
EzL49vVSVYefSmKKLVKmCqw0WPxQd/2cMoFyU7pjBq8xvYMXPX3AlIzm5uOda2Qk
s/osMtUjmDHID29FExJ0Bjtyd+A/5J9DPJMqWt04pTRTQiqw5ZldYWonsi9jaEoS
y66O/xsK6qjBBYaSbRTN2/YliMl5ZhQswwIPnqkgQyNtb8A+W5MaCZJNqo4wFg0m
NMe7D6dZJoijrtBM8hCLIk4xcU2EU8o/FATpzkkBtvUXa5DJkD8qYxsSEOD/vChd
yDB47ktzI2F74kmlBTbjT4mxiJCgPdrkd4VALQxQHY4BZBSfp8IwRh84t4WljI33
b4jNOnSECmrt2gfpJ8HfUg1WmUXWIhpYIsN57aUIxXRED+OQo1KNaeU0UY/T2kOn
7ety6WkJMO9UNVHOP+374uwaNjTMMxztds1hy1K2XD5bnyj2bh0Hi234R6Z7wlzg
jBM16uEQPg6HssvbwDzRrk/RWtudXlnCq415C71n+J68U/K3cJP6hHP+vJmoDqQS
UqJstYqnqno0+87Sm5tW5m5Z6Y5bbDB7Lko3ISk+a4SMr3GIB1ru+gl2mht/uoAi
O/PUlIMJ3rBZ2FkiGKhD9pdH9DLEzn9VVk9KbDj8eu8BEBFQa6iz5snZ7AgZuutM
Vq5mj7iv7w3P6PsXuhpT1CG8oQz3zPj1fJpCYly2XGoCRwCv20PuAtvG4nxz2LEw
51trTD7sGSMKqTpsZ+OdZ7Wx4AiZy7Bb+54LsQoH9wIoDffhaCfe5DWNho8dGRg5
tDcTlY3+ee5lUIWyGxJfjPADtVDEXPo+lJYxnJebzywMpQ4CBVumTSYjGsKz/Nkf
ScG7zTqYaPvSJN9DEjIxzXPn2sKVJpafs3Hg8krYDPAwJ0De9sN4/y/tfikt3BqT
fQ1lbXB+a4PYNoCZyRJxq0BQPwjtDwUOId7Z9nsXTg3ltfm0LjIJasTsv2W01nXE
VHyTQYJ/iAR6YkKgcSXqW2SHtgMnN0xlzfc/MlLMFPm15rI9D4xhPUSXRCaRYaHS
+IjphKsESPCQrlNSoxg+y5woRkyjLWfgWNgRABWCMuG/25PZk1Pb9ikL2zXF7jFl
GF9KOAAtI6NEXQqPtzJAb4VmBGBBy7mVR/d05Ot+WqO5fIvzHtQgjn/nSVkdPSQz
lyc4A0Ga/DEywM3lxGDHrsLN3GC/Ykm6256RwPmX2wZwML0iUMfKVR6WoceTICaS
ML3A0Q59NmWNcaFI1RecGMvRCo0UGH/DKlkWR+aooEj8eSygvTxnBP1eEtSIbPOE
18D4CgqJi2PeBB7BqBU1b8o5ro4XLdh1A39O3viLQXAgdG4Ji1PXeQ391M3YReAk
xTEsstT3HQJVCcvKpDqGkP3yHDzOMgkEKve1o/M/LdBPa38koQ2+Urw9wOWXBsXR
HjVpTb1epGh6vdzbyAri9LkHN7XFYQGPAXIh0AI0Hl1wzEayHEjrit7R2uu6mB1Y
50UnSpB3IA3WkZsgYQ325hOOMFmmYxZoQQ+YEnhvhPtXC/UINtMVZj4/H8hietcI
myMf0Yb9NXzQpwzPLvc/4CM/+JXmiizcaGyC3Qbol7lxjaZhh2XjejPWAku7Te1Q
eVhDOb05JWXqdvCH3RBSkGpplgl9nvw4am4Hy6Aj325suejWvb5NJaoVfDI2B66U
eN6LBIfT+WG60eJ0dRYOQhCQRlCmntDJcCNVNsr0eE+kC7ypLHyT/CKGDWpYOur3
4hNp+QAJrX1vZp1Zp9dbzArEKjFPZAsf5vYo2hCAFJwn4UnxOJF1OzSCHccDEAVZ
tanCGEtgoyxb7yZO4AheiYP9OuANoSSo4U+g083j54uE4R938pjYxFWcrruroM8v
zBQVsJ4Y8CTEboKRRoxQOUwDByrCatpKI5O8BKc7Wr0qczd9f1qWuVW+GGUm3Cy/
7TbB6Zw7rPUk0xBUyyWyPotSPQAA36f2N0I5+RmgY89ohXPkfb+N7Q3R1e9xp2cW
Rg/re9CNyGL8U7t9WsSGi/cQ2VKr/yiztW0GBIMlMR7Ve3lCf7Tp7fZcUHJ9DaMu
2ePKGG3AblDh/RwqGoCSPkP1Sq284OAza/Ib63lNqY4QyJzxIeTiGmuqi8Rjwswm
1kEdbNTfkV30qLfNHXfCfFTspGNIUy+3X/CufvZVyhV7VUqpk8iNJSf8SI5/Hs2J
pBRv3/nr99qonNvGGOTK1ABDH22CZAS2FlYwulkAmRfIhX62o1fZJvFkGsFqX+IN
kl6e04N8W95NBWd0FdK5CarULU3PPah86aakM/S8hO20LqklneHNqZCGBWgKPAbP
jcfXpuJ9aiuCFblLKiuIbKpeu2YzZBKn2A/kI7ZFnwHk8e3N5JTyb4I+kCf1bNz/
OzBJ+f0iC67f157rq4Ly2YVTbyfSEhvKtwheVsHC7B7Y9VqJVcFLWAg0KcSzSZ5p
sCiFxflMQlDmQrg4vWKxFn16qZamXBf5gexlG7+fYvZFexiabiiqlHnso/vNwo4j
P+yNu90Cqgk8PdSs/k0O0P95WO8/RMfEkv7KpXpu6mS7oxMx+WuSpaTk1xyoslR2
4ffpvLd5tAAhnL2Z/84zZef/3Q0OgGx+9GYamMbAA5ebjqJw3Pore1AqloqyC9si
NZjTBjX2puJyati81vEUcOJ6RIDuI1XSFoPSB641/JrGzww9xwwR0b7a98ld8rpB
zZkMkIKyWg3fydhJlcgKD4nNnAC3nGMuudOPDCU+mjaPxftA8khylAHmLQ9Zqfcj
tDy9Oe6pOumigXkS59QtBeJPaCDNSiWeN1ipAnpSC3TH8CTy2yW5iqXlTK6+yL8H
Kfekaz5Er15ZO5L4wljehoS9XxTTzJMLV18qt/JDGWi182EMUZ2aBscFgM6jUeGq
Z82LR7lgwu5cMDfNALwiaP+twuejvx2CCMx+jOGvYVY4f+GmkOtw4zD4X10LgwC+
ijPYETSNq36wfsHxyAzEyl4AcWZjDbDHMvITeluaCJ3iMQOgfHIEw0sZMpME/EDM
tqFMmSDI478sIz9MqgAMnSN4scpUIsUo7Z+5WUVNgUCUtKL3wrpkXVNgM4J9zbwn
PryyZJMZUjnai4JrNIwbmpR73oCtqvtGgD9tju8tftI0Pgdw+mDWrdV0XRDGuGzP
ATvgZPDM0UJWs+qwct74GmGgnMOA00TbqmRBp8//sySbW0u0eT+8LNV37h59sj5c
CNby1pZ/vNqlCMNbb+/7MRntYrgs6yK0E2a+01kxjDYiYGc8Y78YWYXN0rsi6vbK
mn9VESDi4Nw2jjPHURKVL0vNKp2W2SWhomxZHGs9NGZSvxJIAoTN59nCEnNJRSyo
HjWU2R4HBiUwbblGzPElw0YlkG3huUD3N4jtTI5ca/7y98RmCzt0TD2t45FSs1h2
/1bP69xNcJCLdH2cC9lRyrbG0BCwrNQjx+BdaZUZVLtELvJaPFZPeipCgUIU9/eO
orPd9nFzeAwzoU2s3L4DY+tc2VfWbspAWDKzoQ13iktEWopVYHpZvEdDFh/61lSG
bPO3orxiP6pTwW3wNHStT1rJ7VZJD/soxJD09+9Z7NO9/6HqKjGVnvkvz2Fk3oPp
ttbJGhsHPkbpwHYjBL3FOWbhfyNERsPTBsW1eVtwJl6990v2JrhgNWxhO50WXnxs
KDluhFxUUXPzjrZuxnu+1tbxI/j4Szcatb2ypu+iWFjrEmwZRUWB0KfTrvCEz9yc
1QQt2Xbq00z+/WQQoFx5mfz/oFGkx79aCIpoDxsSdDqjghVFlm7cdjLmZdeEakio
z3u7jypA7afeeZSrrQ2s89qCr1Pi4yYPJKSvrQ1e/Ft0KWsDAER/JwNLZRb2YU+8
XLRaRjmOsx/bhkSTltxw0Dks6DrGJNJwIIGOXi5HJFRRvaTTiKsIXN7BK93X5c2f
zgj7Tyj3j5YptHFk2E/6/Hv47RqsDrSEfw33rNkd7qo/bdR1vIVAy0Dgn0gS7lZJ
WG+jNul9OOzcEGZQLRgndP2gfSkZnaUBQP3Fi5gfU0NFfgLq0co2KNVycOXYzUwe
7ff0vTEEdONGx+T6YdITus1rLD/zes51KkvZWTd7Zhuvs2JL62FE7aC8ZIUBXm2q
Hf75ATsF8nHu5z1ro4AmymSi91wkzZI4x/+ykirUhV/hqhp13E0Hf2+ZdoMYmB0t
gWYOlnmAtXwiTWryUe5jIxCqLNZeBt0jDDssSlMbQc7W0kgluQv0uyQrujcCD0iA
vGXk/RuITRglB9cTDr+068o7PNt1Sj04eGg2Oj147UZcU3e3OJ7sx42zIQtKGHQs
MqByIVOiJZbbAdA2biC9wrRBYe0XNZQ5OToMWGBuhL1CWxR7nJ8y3sc+X5VpnXwx
NWdyPZx0zCve3LEuPAUm03XShqtdRNTG03OWBnkvfHyfbr4Vly5yu9gGa4bkqSMF
tetfpIXaiZT39l6RcSeP0c2hLYHkp6pz+1oOxuZwIM12An8DaxVp03Da+aEEAyCa
PZLmbq5T9LPmheJnOc19PYvvMsULHed546adjlbcgALuVSc4A8Dnjt0+ZW6Tmdsa
QAPkNNyaN4tCmF0sVySP1PxSJ2L+6tuUt0GgCaaMZRq+Yd2D6k6ob1oH/zsIdl83
1RXABqjBFDS3kWZe/yEGZouTn7+VIfmNUEV7T3qbrvhWAL1uZOEakbGfw+xP1pz/
swbuH4Nc4gizBoSrUF297clvnHoS3DA7i8CryPvB3/ZRgVTbXLjAFaN9LWYG+Jro
B7/2wUX1WN9k1bZzVbUAYJeltQlPqqPgSQ3MtOiJJx5y26ov/shd9WnEItRGaVH9
avZyOfoixcYAw83fwyx6llMbyT665QyoPocSTlo6ZM6bL1ovefm79jezDBtWWWGP
M+vVt4NyY7PoU1aANPz43FH9Zrp0Rd75CMOXYU+vN7vVL/y/BrlGPRalYLwM6Uq3
K4Rrvyt6QzLnvePNBQHVqqu3y+sgb1xODHmgZ3H421PSldbnIpOufOTSFUrmu3Vb
JpWUsl6I5S4K8cmAXwPbL2gCGms7Bx4hutpUUqV3mxyQcOszTFooqB/fLqrIMeE+
gLUI9Ro+suJy23LAWtSF/tE9lkfXiI9XAVgo3J/UsOFIRvIRraz0vVlU+TRlK1qa
45v7gCjFMktyUV1tpje0YWGiy3IMiyxeR2xLBnv2fgythr0v5WiPg24JkC2POXsO
FscsQPNE/tidkQZnuBVoiSmKeCxzMrDgNEU93eqM4QryKi4klKM2IkSRrIX9wu3z
JKDgfNelfc6ZKcf3pv7Qlx+zDdysPP3DmeepSLDKBIet+5ShlvC9MVX/HQ8v83zU
QN9sDYbwaKx620FSZ9bxVFvBK66/QV7I+ybXPwQ9yQh5c361ihteObsmUm+i0uRf
ZogSI3sVYIrij+x8B6+xGaDDWd0gGL2C5RHp8K6qzVLezEOwquPTftgXZ2yiW01G
ofQKbGp3Ry4FMT1UtjiQf2sX+IgRpd0LIwiJNft7kljs8xZZ/6HlGg+wzPbdUxgm
toUqI9JehfHREO2a9xWLLKfYooFMnq1QwM+Zm4PX9UtQhIMzPE+izxenoXqAphAF
n/Bb3TYbl60j4SBF0Gh3KBLjnvf+RZWQsr5EYEZqlrOObSajUYjBrbSsC5azHhD8
/jq0ZxS2I2Fpt6CKvCx+cIDr6bjT2wMJwAF9QuMuCDN1PrffdHDAQNb+hMZYKN+F
e8Sq3GSql9O+ekX10MX+ILz0fuUG0PFLBDIY9GnjMmvgsKsfa+DOYiVcAOWx/4iA
w+2tWrEq0c4n65BPqhkl1i1HPsKMbwLidY7phT6TewjfeHDHvKHjClySxe+RXzOD
XarrVvz9aylhO7qZRByrRuxFIbZMgBqXFgpLaeJcNGflkT6GmVouPjTq+BAh5bJ+
HUWaLSj6wqBv+oer7oKYTQcYuDj8j+/TwM9mmOfAxVzT6EPSbinlccMY2/JJ+RCq
3pKGzJYsBklyeG81yS3Z9jYUrMcw544+g5z+V6AD0aHfJqB9R7W59mO/nQMAeSvB
oQFt+Lpv/i3avdkZIDOOcaGkGyOZHHdxkUX+u/9+SjUIzQSYk21qQ5ODnq1DVKm1
MgcVlYlbUPZW+u6rLZgH/srIvbVa4YAqeKTJvpY3sU+yBR2RB7fJEcY3+RQefvqK
9EyRGOebZiEA1ba1UpVlGuYGxN4M9BGlqdIiG7/oSG+nENivqUPOVg5fmiFrIGdo
V5t9EEqWtFxwUPt6Gv5bklgUXC30bwnTEZ44YqTfwvDXQ9GnlX1GDH9PLLxpbAjL
YXAjd/Kgdz1UbZwIQ+6plc5IuJIelnd8E553nU2huqFB7pShJr0y5v+sM+SJXNmS
DgFqMMMiPdJpAg4iL9f3kAYM22M/vBNuKJ3kdTOMcZxF7MQfbNHK/u/1Q8LQ81eg
PXy3GQQ+ZRPvlPXlcNd0QXoZqf1m11qGZug7Rvk00aT1dkXOrwzb3iuqCagtDyLG
JfWYghOaqBbK2xnTYn7l/pmK/QGoI2HnWqhBf+ntJkLKOsXFQACt30S4M4UmwG8B
m/6GLKw3K+dQhahjms4mRF4cBPoNE6mm9qQoHAX/RcXcsHAKuly4qGQsRojCRh7u
qPLdcL7asnOKEh2TtwUXN1HUKjHDEGwq2ZhCnNkoq7sj48lCEuWR2fK3LNPmbYjR
NsTFHzTUq1/4far9UHiZ8NuFJPtr57Qss/XBWCur578YtJmwmWvCFxmSKPLTru1Q
KKvOs9sxsI3HNnpRuHI+IK6TfeDmtjwmybNQ4IBvoCbd0YSdwBNM7ClrLmn9cheX
zDkRNd/gVlO1sDZKj2Ui1A99NSlBhv7pNo1thgCiLp3JvcQvUhnRNNVgFeZycYkf
3kYW48uD+159Ic62U9GcWc98jp73e/LO+hRQQwXTL1kWn6i84+QvqV3WIC+MbAO1
AomNQa0rWZ73TdkWYljvIEOAqz6CG7rULklSQULW5UNjoVSzxbvygTmYW1WwFYtR
p2juQO+xK0BNitIX2RGVKuCqwfkiRSwhK8tVToGgszGRpmRxWlRdop0orRcATpE2
SRLTVv4MFYgwX2HFtkEKh3ZU9fJKF1cphU8rCa0qvwm7zc2PBqGrJXE8D+7MmqFR
qkyMd7AL7HLuVdAOCL2JfqirCPbTqjSaBuQ1pXAyyQstkPDFEe4dOso3eA+KGBgY
X2uZaPHDBmMDS94TMqXJJdNhHt/Hm/QXFSTJaEuaXmk993qhKfkcu64Lr5Y194S6
fF3ZsAG2uF6oTodWr0j9BnW7lDsmckwxOXqzY1SMLJmIDn0u0bDlm9pqNr4swiBE
kIRfLcW0SdYNaeq6K3veTlFG2fbaErISdILeIuowdaV1RyBJyiPGyQnal+bi4XFG
qokhp/1slVLWH902QSjQ+5OINbLhbAxQOkSK/66p7TsWcBmzt+pt0hAXiguR3U1c
3jE+spQKcCamVj2OuzpNRkhlEqO9GM8KKaZd6ConGC5f7i8tm1vQ8TPIOSDTSNHv
l8ofNrmfcNLQCWUjLdsJNyVOR0ohlT4kTMN92B6Swy56tOiGCbzXejgLYqonbeuj
wJ5jTLLLTKswcE06rFurjKjLyah2TNVEpmti4L+99eg8SsiLkyWM0LRpEy5tG0Dr
AV6yfWrJQvln/c9+R1ycGLJpINRKFP2qZuM7uBAYK48W4dF4S4aLBqPe1mfXGgcZ
ntbk/8dAcngj+apxkgY8R5qO85hjaW9URpd7v7/ZecAAQvPFz8qb9DHRJ9M62fCz
P4tKqoo/nqtqHY3I7Gs0NHGjTErp6DPQF9dG7b/ItLt13SCc4uscgguAlD/6uMuz
sRbUmZKLLRgUISodC0df4VGVl0j0+ts7Okt8GSG8S2r+g5u/mvqDGlxwg8JL9em0
kE4htOgKmh9G9goPpqXNV9hceyRiMVfouVPPhDKLO2eB0bj6ux2xt86Z5hJlwWce
ZRtO9kFt4wLPl5dRrQ+w73QOaA6pxYF+H2iCv46NQhc7+n4jGi16O8VHoOTitPTo
uADPokjF/HkctHC622zGrpstsJWZO+NFXqfLAsBMKCyCTmxTrl3ZS0f0F0xsJFva
8MzozFscSyaXUwsGjxRyAFXKZOR2LE3m7KMEjnnnhr6kIWUXcrbmxJ4PJmiEMVHE
qFZa9tY6KnAfN2eDftheAlvydcWPwZ+DH13UAa5NRZO1p1LRDFrPms9vaZV5FePu
AkntmYaMD4t+Uq2bj1TK6ESc/PcfN+j6IEvnEUKlxIYZOvFdyLLitiVMSB4x5Jci
uCLP51PcF3/wnC9PyzdDSsC3VcX1tlkT4deyThRpav0BH7TPVN/Thy9yI7zppwDU
uMRXcZ7Yf1/4A2zvSAp6PhCn8WdlkK+nOabBbAKYMQx6lP7XioZGFIInN9OYSU01
5HQWDQrRcwbL4toiJTUCLAsAi/0beNluCVWOrlGoYk+Ca+ypooPQIGl/GnagVmmY
F0hBom09EiNeXWCHOP4x+i0WZvJoy9yFfYrAiirbLlXPUB6oN/F+V+gDoCjqfCsX
A7RPKlvMq6cHJwX6dkb2GnSkxB+lRIaDqjZtyFEYpuF4HAD1OTSI/lunlDnlvinn
giC8/PJ4m/flHApqIAHWLM2SWrSvNlYXK/jto+JofFI1Jato9zDISp5QS8nkTgbH
Kn9zA6346QAKulj6R9Pdj4FrYxjU2kAZ23lO9ZihX7DIBpz50mVfqGfdnYp+s1ZO
uVyn9DqaFmEWxnBgiY0w4G2ahyCd4lpahp3DkhlHoFiwx2qAIiWewn4escFy+68Q
YjdLEB/UoBdp20/LA2ZEKnFwNMuiYA3CEeSuqv17Cp2ZoFYrZFG6o1KX519R99EI
q4fgEih+Mng1jQTJ+klLhTe/WozMF179DDdyE0/MKweeIF6Zdes2NDf+pNQP9rgw
5CMUmqXHkx/f9F2Zjh/xvn6OmyoM063qoGyGny5m2KQ35uiB657/wZjGmrlxiGWq
DAcBlh1mheKFj2VQUVUpa6kALeNLQyZCCk4oA2LyhczTklU96xE5CSR5j8lYMUg+
q8EDB7HoyfqMP7faFYdCC0JuGtY4nmEYiRtW5/UsWpxwl5mG58oiRXlZ6HNZBlcS
TuYyzyYE+bdfnVfC2AlLBRP9aynTVtbkoV1CD1IMpHZC3J0ZgHy5fy220NVX1cj/
i/wrEIZrMWVLpQbIwtfI/5SJ7DFJB/XtMaG8zGWgEmFi6QlJtZciETMmNIyWV43n
aIV+ma8HHuknRrIpflYXwoyUxdSLGlsRXtib+rRdZCaEsbEGiVkoKBpm9CJdlDJN
THssLVG8OJ4h+XSEdM2jdZbpC+CZJiQbgy59DV4cyG7DimeO3wVIXbu0gvRcmYNh
B8xSlYkHN4eZzMtdQM+P6wD872gAGBMVA70vCKhlx0ZQ55SXcWrd/oTT5UGpe5n6
QxjTQfW73UCu1vm/kAtziNtYT/YdCmbM+AU+h9xbxmzWbwuB30scMevS4eb4hF7k
bWKpKYBQrU41bu7buUwhmtZrMc4CIp0CfxuNCNiMoQxq2f0pVPQGjUbyE3mebtOR
LCuS2yM49UwSXYaKyfcR425NJPesLygjPFVeXb9L1ZuuJiX1Bq01swVzpYc+QMn5
B3Dx3xX5qYXnREG4PRj3MXxWJHAwkOQn/7Zmy+SGkculvM3S6KX+mBnNWUec1Bti
u16KRHeyXGMmh1wGlNl+y9bwm8Xw20lYZx6a5dAFzd8bdpisH6NY4VezbWbD02tv
WablxdyFjWX21taxd6g2Ijf7gwXK56+iMGmckuWBN45waOXhGF927L1RLRMoPMn0
40Li2P/Tk9BXgg/9hvR83I2kWNavA4892szxmhXRkCAyb6+GSdyCIE35rux6wJIN
vRA8SGNe+i3YROK0DXi9fQxVeFY/N299GkL8HPsU0g/RvDxwAbydcNZjjhuI2f7y
uzrvbHdK/jPRJpybESZ6S9Izojp+DJv5yLVd5JlmuELvYyBps/VHjJOJsn+C7FNs
+a1DySAYaBmRlsboE1LCYQw4uaiPbFMWpjmp4EFJbuHRx3hGl6og69HHma6axCWr
Ow5GQs3JNhUsKWSkK9w1Vmaq7mfvyOui9ckibYCDaopWtOL+jHzm+ySVICJxpDVD
mEeBU/k4/a248rHpLhp8lXr6i6c+//s4sz+RvjWKaaow1oN0cC2e/QXiJ7Wb5EQX
9ezyx0d5Qkj6K2kbWWCm4BqiffoJNHLSODA1u6GontYI33uUVDMOb561OE27sr/b
rh1Ee2RBrrgId++BY2kzqKUhLkpaPVdm/2wfIgAkzOElBdgrwOHo/8ZT4SHYZjMT
4LL8TAsvwv1rvxTmxs1Z7Ij5dDtDabCgiV3L1tNUsEcoULfyyxgqsQEvjfDpJh9y
1TDUgMRXT5jhftXxyXScym9/TxpF+upodi7p0U859yFoFU2LbOXK5tkNzZ/oeIti
IRLEE3Gkcy2ydVAJfbZpzez78HAAhm6AXbpXzzrnGTRIb2y0C69oLfSJG9AHO8vP
/tQR1sbJTmuHsbJct0TkimUwx3HpqtC5jvBoUpcLXrn9hvPV6wiUpzUiArPEu88U
OksmbspNDhre7HmcHUjW5s4b0EPeKiN8KZRMtTUQqb8z0jyDylNt4ZFJw/jd/Bs0
Xsa97uj2NM5XARrKW4IMMtQf38iN6LB4XWvwJ7b0YoeSU1W4a+UPMpwAIcDlwl0J
ftOe6V2nh28X2UPFw0iRnhVvMVqYVcxonra3XI9vKdnze4gK2LwpKzb5qjunJbrw
3x0NvQOyYedkX2Pt0wpby9apItVewihYUp+rpyeZpjylerlHPqWSF93c0D9MDx3L
/Uk4DTwlSX2UYpyAgWCX2NYl8P5v51RmA2CljaLjhm4yq0bLqpAPB/icocu/EydQ
ZQYk6WTCL43Ewo3wYnlZgTrnApuewLGeBRhgtWI+lhipL/hSKm7JvXNUZt6UD+2B
t4LqUcIHuu/1oHryZunOOtzOAub2bVZdX3lbDLk2edMRNNpfk9CFw7ETv5gbNWKP
7aoIG/7Fe4DRPlii1d4F54BuxLxUKjj4nxhutqwu1+TVkmApzKkzVqOAaiGLkng9
NCOmwLInynZrNdiULGBvBHvElSJF3A7fk23NEg+mvpW1AUCx8gRsd4m5bb+6XH0z
J9TfrojJJXkKy3jXmzeuuPvbeEU0v+dPgo4wVVu9fvJqAe3TgH/9THYHFmQu914F
LqXN+Jva4qJVGpB8EmyijTGUruAPBsBsVssgM2t42wCcsnZMOAUWOivQm0Trl3wO
gaH+c/Da6b+dFEhDZGRIq9dstm+lwnlGnYdpFlGY6brR1MtHxPn5I45vyfFVaqxX
SUyKFu7Ljn+C8bPWUO49IjO4Tqoe3Y3CZzRYts76PVwC/0WH7hawaCww8yUdgXsp
Ue0l3pKV9Xj+mZ2+tZ7zoP9z6UgKvP6DJM5GoO1vzhTB1a7HKon81KoxqNoDKBPm
03iKYQYjR3i4NmaEZlWyeasxGakrg4dGrhSJ5p4J1/Hkc/aTNJ0BFidHyzanW/Py
sNm2/m60JCN+hdPCGrudJp68AOJZBdWH620jzfd795fsMVtnnH4l/w+1sRxk6ZnZ
g5mCN5GlGGNHTh0KUXr7vOl32H9WvlUR1hVXP12adfxBEaZDyEN5y6MbTs2+y8iy
iFaqFZRiJryeiCDrNIcj9rtSA+TBZuUfRRM8SKn97Lpl4OxcU6bxouMclMyLi/hJ
MB24M/6CJBiMYmwChtBe561tCYZJLAAxoOoIa1bt7T2KgRZ3zK3StVdB41yLBV1B
nEJ/saO9Jq60SKHKSY8EOVSzncBvFR2W+rpjylTyEAphnudHk3wjt7xdbvc2Erh/
c0kuPvQ2TSHGMxDf+WrXDkTdJgCH+KBZJuX5ftAW3uvHuYxCxldx5Xr6xEzhLeG3
eR8wO8G0i/9R0iwGI/L7xbBpi1q/7XQV3Dm3rGz4vTG+rQkmp1UAmxH2B9PjWfnD
BXnb6hjpQ46JYe9yJ5fvgxgjXl9fFsYfG0MPHkkasrELrd8K551kNv9JZYIzpM4V
s3D7/lYl+0gK809UX3FGNFNmAUxZvCnC31WrSEcyos5fHpvLTkJhdO2New/i2vRa
FpZlLe65X5+nYDbT6SGo/Q3RFr4npiL2qYWbetD5UaPt8G/XfXf2aB9SjZ7h4wvd
lhVSljy/YKCgy/0nWrP+E7GN4z6bNQQpo0vHV6Wx/O0LDOIsIYz78mHn6T1VGwDd
aJwUl2XP6p1AWMMwP8q4F6Agw9g0k5FuyusUabQpbnUD+kXbodBi9ZrM/7eisG0J
KWfyseO1i3xTgmnaYYriBmn45uZ4OlnWkC+k/7jN5qJx9KyqdwlODN8rh3z4N/5b
rQ9BHmX6OV5Dew3JB5BTipdF7SkThwuYyVdHqtXzuUBBadjyPMp+jRqyOqG5JS1j
oaBxBunnq1+5pRN+32RsXmvc76rQPgqcYVZ5xuO91RKcCv+pavoNKQVI12Bo4yUg
2XVSe34KCL/Yl0s7xG47sPi9oY/YCs0StvZpyyxKIvSva6svlid5mcn7ILrozKTG
A2YdE6TUHQKShdZmXKu25ahMQF6kg+ATjC40KgU8W+5r2J4Cevmbt7+syJICyMXr
wTqvVaTjO0x7r6VQZu13kQNMwVwQWFRp0Fzp/aBLIblxqA+2vN76Sl3/v8R4Rj46
9HlRgQYauY32eo/BjSXlTi0Yf1Hv/bzuDcrtTCA4+oAD18niAiOOPkmYjVq0plgm
pwV74V20CQHSuj8VOEZlKHTHwIiL/6s7RHIL9p9OX3HuL3jWnq8dLx1cg6HeBAS6
hOYenW4riJUHqMCp2lA+q2KndVKCkQYyQtwkP6+cM/S35eMXIafmrhpGGOz+wAAO
WpanjPCZAepFs3CQuOQhU0Po65syL0CO2t7RiR5gXfQNxZeKx0XgZG26BJrtoNv5
ksAJrgVXp0i5+ixFK1O3oZi4L02GynjjqlaIeOt3uzlzS+XFC370/HO9BrSFkTqn
McgPhm2js0XX77Td4TRBB6Ucug5RTcS/RvL8ySQJ5BTeCvwh4ZBKPtRtWOvfRLyK
SZx0yOxULhzbjjVeCUepmWLO9O+VKxqSMqNfwUahFE6NjwZbJTj/b4f1A+V7BxcO
yNRrNCKQfeJhb1s18AWZEUyFpp3dsSHF6HOBxjvro0lmt81mMtn9FWfNaOTlHChd
F0ra7MaKYM1+CAzaMBPnemkawCH0i0aqnELlEBwPbhpk44Csvmq82ht+LSU8pRRo
wCHF5I0hN3a7ffWvAIIAfyJkBQXLvtKhx0WaCOpvg4Vv4P+QxV8nxIUpG6JVM3AI
MEwvQCziX/4/0N2zBu3yGqDtb+p+RIRvvmYD6bIm2EULau6nZCHHamu/Sv3yFNBU
GENiq+ZDGbpjR2FRza9tzauArvADqWFRx2S8zydgC6TrBQ28Vg4cnkIuh1nuckSq
dLqsqAwu4iGdxSrssG5AcEpgMnNvFWh70VaHguYwHkB+X2NP+AYs7ZCl0NDe8xz+
uaqAi562V7jAOqf2E7M+YQMYFYpb+6EdR2UoG4iFOllkZl6vl8meJLUEYxBzthDP
zFA4hU6l7h3MIoL/lHFpwK2M8dnCr00tBiZCAhBAifFeCwgUx7LT1/AqYFt6eOW6
q3nte/6/JSFJW8KihWyP3RbMlbeUZmsqBkz6usG15dYiR4wnXaggLI225g5HdLwb
6Umh0dFAsQfeWctHa5mMJaYzJvC/3x823CibgXITqx9s4hgp21QVFM9avzwW8wTm
ggGS8S9TJIIf7pfCXT0W0SuJgiXOXEan1RN9xF8hzO5r1F0KMvwylPZXBUKOv3kE
+k8sNvQvktjGK7UdAdvuLC36Y8KkXjWpJrzTKQpNnukmjxaPbvpEo+lAz2zrxOu7
q3rOWVByJPNWvlBWQlFbeFMiiKBMxehLZU3bnVId8SOabtcouz7KhpLHVDbCuqmI
YhFitIo9HibvKSuf4kCLy37P6H2rc1nLIUUFtGPJf3tpGG8aBSbTaddqltWbJ+Ng
+XFTyXpvn3Ttboxwd0zsb1mSsoI3Fpm26SrSCrFYYfp+Bv+qaAjr2hM1+M4T62dS
JIcK0gIHp0mQcNuR/cBzxTzgOh8yHcUvRaBFc5Jhz8AvYrz79zZrPJYnrrEJ7wgl
+MnLm50l2vSlMIYYFee6K7X7DZONyFywobv2t0QtI5gaTc/daleP+K03nPEsev2Y
KvAnEYlSc9YsCU4uLE/inDMw0rJ0d7wDXkUpeo4cr1rrut8MEEpbMzf0R09svm+A
gK8Jw1ktC2h1trJLQa+fBaLaOkG7JpLn2OK++yC6nE/7guIY11rN8uEzAO6CDBPb
OUnsDr/EaU+QcF6YdVKk622lWFgucaryECvDbvrwsw/JmvnVn6+CvqKpcKyZrJI9
Ihw10nG18ika7yk1NUjltezzKDph1AXTQcw8UdrIAj4g6WtP+6NKovqcd5Vv9wJ3
zAdhOh6zrtmpKLBNe/tx4QzDWhYv718041itUOmDm7BsPeFuVy0kr5qDKZKrIZUw
5PMFE+dXukbx58Zb+8SCnSkG7ngay4fD5IueSEdgDSQVAxLM8S9MsN99PICnv+gV
InyIbMv4QfSoRUCqMzS89oBh/82ez9KhmkZJ4ivzX8deltq8i1GcNSP06eZbVaIe
jsdirNJrMVB70bj+UYfsLzzIjJbN9QGP1wh/+LwN9ayXMgs7+HYwu0wUHufMX5Uc
hkXBVXCnPZm6ntPIXH/x40wA8nH6w3GTlsr32HAKVT8vbHtkWduoBiaUVhlXBRyc
KTkzuYHu8vvITXfQ3t9DggTbOJwk5pBmztbCeLFA+oQ4eawAyWV3OlRkoIlZCRzY
aUcfq9FcMfjAsAi48xiM6LcR6tIvLt9K+XrtvsIUJ/YjEk/AkNNmkyTNvs1v1LmR
ZSUZpM4xaS4+a4T6hkrNBJNyiS9hrJTxCJQeuniwhSd7WhRVo0KRUkdC9J72kJg9
23INAxnIxq1eeISxgFzMOToFjHuszGiOVV3tgsplJ3NWxYcNE7agd0f+4tMKiYt+
NG1wagmlPHvJ9Kek6jG8eUr9Wd2T0Yyu2QnCWWW1tTIDRAm8ofSAUYdmuAUuw1jG
EWE1vGUCh24SJ5lUIArxhrbkDsOz6QiwhZUkHU67jviki/ubI4U1skE95AFuazYy
U6cA0hkBYT0dpoS5p4KzM9X9mXewPGeLkgrKZvkpomxHpbs8YpqpAUiLGj/PlNEu
RwVHm0Ya1MnQnEWEGcO/ZTkdPtZz2Nd6Q5Yf37EzoAArBPk3YuW1RMq8ZcH4KZDo
ZsagB5SOJXrOZSrg2HapLibMRvoXnSPaZfDbvZX9Zp71tvCRhyAWUcLcJl6RpYdN
qPSWrvSaYkNuposCcuvQw7MwOf9INK3GXgeHA/yxBZa3bAHIfYGv7xUNX4u8AnmR
+8rhuYQSUR1Bh/OKgEezW3l3ouodi1cw6ayQpaOseqbZKNcJc9nd5yfq3+owBTqN
P01xUEP29clMBUGdrQXIB8njTOOkueMTCk7MwKAhhKOzwMETTdCu+NcH/TP4im8W
PQma05AMQs3HTpkAChgoySYmXFblR5FuMBY+8mfmTjV/jjSFZ9qRDusX2L7yRrWv
RAXIkUDRAwBy8gUkeYdzR0dyxs7k7vutoec+9DXKUL7jypcPWLByWgTKe7x8SUxR
LQ64rblH7H3brW8P4Sdyp1tArRYWUDOnzVX58HBcnOSjqF144EtkudkN9AoFOuqO
cmzN0MWYaJb4ZYPw1UcSJSbJ9Za+YiuPVDCkGbrrqU7vyTq8zceLbRAnRX3xIYyU
nwufRlVjkE7yq1niL0I7UeEsAIYo6ARzzkpsmXSURKuwiUzjZODoPDnQiBI81er3
OfPpqWcpTxYLuPoqAoP0yEiz5BOYmfvYaQcN+f8eCADf1wSf2/YlCKJILfJ7mQSf
vaJ9A+rVXnbr2d0EUkbI995Ys5WOW92SY47l/y+Z5vjbgVWwzUJMgBwOEMMs+YAT
m6HCKsCz3psbIPPlq+P52dcYwC91MrONPOqypaozhIIieUmArk1yGgXGFluzmqxb
7Ulz4mTcqI80I3W2xTPCbXF760wmiw7XFUm56X7Ajw+POeuK9kKJ4qmxvlIEAFXf
PlmujSOf+/PzhTGkaewaVRA1zu8a5Y2g7cKjN+2TRNvLKsWvn9iQr6aegQJT074+
wQoz5PjM78Zv5jF4/9t57IGIQfgDlDxsdkl0dsCQOsK5XYK2ZKXNkMfRXYwrXiRd
eMAXQXEdIBESpq4Je3o+6ni6bQ+63jggmH/7z3NkPZiFNd1v8+hcLu8KlW/tezER
04a1Gc9YU+cgJuGiqotaL7x53l3+ahtBta9UZ5ttMmuf5PXX6o5LANXQ9moca1V7
hKZbceZ46kJlVaQryIzRNmG3lVEcb3HXiAPTwRz+nD2XRXEc0D1ekXCoxT8QK7Ro
k8177FJNGXUybWDiP9gIsdhsUhRNjqCbQY+kI41zH3BNfpJXpZzmV9yem5FZ4imW
PeQkGwc5H7cM46WYYPQLKbwLtDOZPXZJ4sCLn+E5n+kW261ZLhKHrrm5LedJQn75
1rZnegBnmSV11Glq9Ba0m16YovGt4r4FcwolW3zGXuumaEkdSHcZ4cBA2/VODNYv
VlEmCKPBSqyG2ZJUrQkCM83yEQLFS0xHyPA6amcDFtprIYvuD0iJm+2Y68iE0+9+
bNtL8OxHZKj6lOjqpk0mCtiwGOidToCWZr+RM02WwPbKY2OSLngD55wHHbWvL6om
OLUAmGRrituLxla1QSPzNC2xgVBpWgzoaEt4BmSVF74h6+YnnmViO9KaKMat/6xH
WxA6D0+YBMQuOqCJYDulmSbRzpBBT+lk27iKezUEWw+yFDrBmTbR2Q0gkKeqoWDA
ppp+ZllWMZmyMpWcDArxwyeAoXOrmqazVZIKAsVxl7zt0udL9Jn05W6JsE1nQk5w
sloImqtuHwF9MhpMDOFtbU/yWokO6xfHR0ILyLDxMfvBirygx/g8nqac8fkglg9b
d5RBYDB2OWYY+pJfo0h0h0Efn6rJDKLYE2o071uanO761EJWtKfjUgE7fbu9MFTF
VAwuE8wZTDXuRB522POvVjllXyiuyDUTr7w+8HhH31sPRgJc7ld3Od2BTcj3139J
O8yHSOBFSD555yz1gnfTgo+BseYO8g9mkdD0Ve1e+6JMai9MLV4WnRkMedNLDm7b
EjXF0FlLiYqrMvLUn1SERvww1mZ3/d64NYgdBAw9Zwy/hBuOhD1TrZ6/om0yhiOh
1tVnRjARI5PWuTIEw5AJOlgyyzdD/kzBf+Lp18/ySeZIbLHr3Z/wsO1mwQsuHaz0
xbHWnQAZCbgMrxkysLfrY0Mf0yOn5KG/SFJ2NwS7EUb+uTmOZIfnvKqRQXJH+d1N
ZAjq+fGqztzFNI8Aadlsq7s4VjnI9D2McxrG0AzqY1jW0Rat17bOVTiQ0ag26dfs
cZ3Kjhq41ALwJ7cMl+RhswS6zjNr+SZ+aXh6OzlZXEF7rjrabN/yuoHCHJ7X55Tf
tQlvEthAgSRqjsTloyUbyolirBbAsJodj9TPp6jNi/v+NROh/XdjgP0Nu/LcGOLJ
h2RJ0Uttk3hx0NelQfgrqodwdLx+SHg5QDsu9+CZnl5n/95uAcV3oDQO1b5Zs+uX
iH8tFK1EmgJ5XtgNuFX7Dxv1+u6XCcEgleK0s3V0Yqd7cQFk8FzhflJCgeQgaG2n
C87T/Ot2O6EbVSeZ9K8OyucO/YVUJ695TtGeycepEnqrn5SUAGmmUoGzwgflcfCN
PW68/rNLm60EtQsFjff/mHozgUK8gpC2oLQOGWr97ZOwlLnH9QuhzJOt6odLt2C9
JFGzmdZCphaBNzA4Jvplhd8zmMnjpLcxzr2HOZoKWtTQdf+ntzyyteEXrS6Z9xAz
t/8W/OZEw4zKpyyTdzNOOmBAC3FTvMe4J9YP4a1PEa/DcGvQaQL0TqOjt4VWzdSX
99OKWaGhlwY6LRMEcNm2HvHy9KNSdbTd0iNZw0GWfYDZJzQ00lyWQVrY0zvLHUyt
1I45Sb9kYmCM3oSg21rj9C4+wppFu9bhzSMpAdAdH9iEvTJvaniFH7QcV/VrhSGT
bvQlvz/JGLZ6Nms8EqSdl0Tbswv17Piq/Ahgbv/sfZiwEzTH4rqxC2G5a1WMp54+
Y2/HT/pHfoNWiRhNPVRgVuORW809CZXaR4JNiC0c3GxC93Fk2386HDE3mmSafrL7
IL1Kz8fc6r2/KaqXVAzYxdztu+AF1lrzEfUalGY1VXcpHd0iGYVvXOe6RJPWLiqP
aaT5XX/ILJlQXsJC7bR4Kphf6VOxH9SXqn27jQMWTmKfjVhK/suxKtWLGKJmMEuJ
Syr8JKjlfs/1jQ7pVKLftyKyWHGNBc20TcwYJhQhsv7T3gT8PvujnlCeBZy4HMQL
84c9rFbMMrtKyDAtjhGlF/DeqP7oGYkvD1P8Bndr2xi9505RZo6lPhb+9Y9JBR5N
x660sTINlWgYG9FG1WoM/UO9bv4bizzmgVWElkgT/RfCTQMubpPOEKEqKJJ8D5ia
bKtZ0LqBakQtQXzLvU9SerutcA00PTTpc/RMo1wVg4qBLkj7bkL14Dp2eHDiPGLh
svVZM2g1VBnJ1/KIEW4vTH6DPHxbiEH+aOYgSxygtkzvXM4q28uBBLxVQjKYZD5Q
Fby3nxA5vUnXR9TbpYNesSOj2IFtVYDCpt/C5EglWO4WbMRf6KTdR+8hwqqOKHZ2
mipowpy3PSGRE/rlW4qdGYBX7JddVH4mLIsIEnXiiTGNSs/dr4SXPU0CJvZVb/Gs
TP1DmKRX57zYrLkavhj6pKkvjNLKVwPNZ7GEuzGF/F/FWsXNXAjvMI49Rj2sQBl8
97Yqb/FQ2dyaYc1vgc2/DaFQkmosGVzXgWOFdijS3DfwuQvk+UWQC00ebfTHsuT5
kwHTbWfAy8gmzQLO3q4SmAHQGxjHb8Q7ChiapNWR7fS4Dk4rqdPwD0NOVPsgTfgx
pDC+I9drSX+JfFnKcj5TqQJuzJwsYQF1r2KONLh7zrhMtD62mBlHPIriGZN+fmX+
B00slhQ0ryjcd8yYjQsozMokreCxxu57Pgu/cLyxYB7w3B9y84g3V4GYPy5VppPs
SVusy57HYklfQeF3iO5Co8obBtphjU6v36hWmhojrFqjDweChzg2N6Yd1YVwSIqJ
t9V0VamARGB51efErS6uGaKKN55NNBW9DGr//ohvzCT3W6tL7nIVQZMokzUJa3tv
kPuxtgV2v4mTs94ZEod+6D/EHntXf/TKBo4kRVxkHnwxQ1F7cEt/n/QIKX1Ndi9x
tPYaP+jVNl00pCrYdwegRUJi8GNInF+/xvemGOpNNZT3WfTRMGJIhJvHJPX6h2Je
1Dm197ICjpM8DV1pITg5JbyU62YnnEKDi2GSFU0bFkGDQ6+Mx98TJekgvTQzFn47
bcPqNkPHrQdXNML25XgtoeOTYBTMMxQeB6hod+4gE8BehWW0c1taY1lS/hjnRHXs
py9OR/85L+IyLH2QiNkkik50gtORNUy3lJN89T8aTPVRDuQakbZHDBWtFm/fDl9O
EEOEjVqr3M8I/0Q38m3rhdI1knFxm8Edc0qeLHncG2p5TbsMgiEX5xpaevMC1y5c
3sGqz5/0HYP1XOXnQxmjNI54LPtjo5gUIlo998nkuL38R+lVigvcWYGRZ/LG7wNV
71DXYH3TnwBduzJFApH4dGkDGGFxRVc3QnA0AXZmNQLS7MHHBN0TJgjq+5jQrKzj
YJeSwzacs7UYhsizmAN9I7lkudT0Be65dW5o1qNXJXXzq25lOf/GTXMWP7APpa+V
bVhKYWzaXQ7R4Bmis3CJOwe+mDw1pzyKRHHG3z5qgjo1Q6Tf7FlhUMX/RXb046Td
DSyl/dgvxNkHpd5pcWXg2+KyfmwiZleI4RnYqOr2DRJfz6sEKwIVMV8cZnNZn8LI
THMh8GPlwfDwEVTq/fXPsD5BMMErIxTMrW2VIy+evTw1SaOuykXegKqw0AVShIAj
aNa5Ix0DY7YyCjqqJZbZXtc0CebU1C7J6HLPLxibvfGziho3WXnRVdDoUYHw+G77
f7sBbbqGE0J8qG9e3U1XWk9DxiukuCxUfOtm0jDmqNrwEPHxdxu5EQQu/ZuOF5Cl
BvTJHW1dZFwoQj84RJvxdGR0kf4QpG6/Ma+CRdh+fZhQDGRepsyQ5FCRkSGZxb+3
ExNrPKnuLZZST4qqkD9TPFEQLXz8HOhx7Fdvhl8hY7bAXo4ruWPNO7Bnhb7L7O9z
Br96g0ib5k3a7Rki3Iy9WMGB66Ao49du02aXLAjGPP/xMcQVBxhBc6nORViESCV7
/3PIWnfhw6bOR24UxrjdICP8qj1xe8emHXThy8fa3uT9A7ZWe1MRxPvB3sisxoDw
VeTquzUJStcBzTmyBKV7SnW8Sd1gfc2Ba0+az2mOln+8rbsaLwaaCwSDFyfmbWvP
0e/NxequERgNTMUewWGJCX1T03GTTSXbdTfnI5VAC/o1Sf/YVA6k0HoljCm3lq0a
ZW2ZPeGZzhPbylmnzQ+bb7OC3HS+gvqx2QNnCCAu9Sh52miuSsLx8wqQ6hQgre9X
ESgq8TVgAHfC1G0xBmXZkUQhRAlb+TZ2TFJGzEFn7hr+pBgQ8tF7L6/+YpyYk3Yg
yQvgLyjjA5RhV2Y+Pf3M37ECxltb25vRwIlU8skYmQRWbNFyQcAy3qkCWvrN6Qqu
yoGfGv9zqjYTqfPWcMmtvJQMSILcJr3RjUtsgp8GtHHL2mGF4bMpNI16Lo/XNffm
v92CLZb7edG3RxK+e7HikOgnkZYGGe6n8dpO5/xgMDsgXhtHDoGlxhUhZRMV/mUK
MLPoiGPT6ruznbypGSNZXPfnKR7OWB9xRedI2BAYWdqPX0G10tz11Ql0wbg3dTZs
wqEpQo+QVS7xYXI1RHInAO/XGgji/P6imufaLsQnNROXJcK+qc/DSepsPO4geEGj
RAQLgMwc67CrZAy68D8YxX/ZYdhxVD3+hHVnfm/OPopDc4uYwXVKNYfmbxGCYxYP
uNBcaH5efH3/zLsGX/NrAfjRYAZwS/CMpTQbo8a1xrgVISzF5Z+hthkpFk4mmYk3
OJyOKZ6JUrA9xK3uQ362N2cMWAKpnweftuyh4ygK1daek6QuOx1o/U5aZDybIIed
ddlgQtQ3Kqb9O3G5TxPxk0lDTSf9BD9LTxEVCd5GonmqECscClL2+eG8amr5sQWr
fZ01TE+W+aI16KchnuoAVkPdL539z2H+GEAO5xcad1GyrpQFqEDo2moAZ1KG5ieK
Xsuw3kb/OJxjng1GGntEyJ6a8a4z5V1Shq/mxai4F/jCt8Bsvm1udOV6lKUWb1fE
SYRLOABBxQdbjFfCWgCnhhFME13XW5ki6eT51Bfo2j2vZ5DbjMu8V4VcbDGiwyIP
6sE6C8RSiC3u6XtX8D4L/g1MrD9UYA9LN1XKB9m2fSGrEsDuY83a03aifeQ7XFjc
0tMvflCTwJ3nmna9lKKD196AFzaeGQiuW2J4awybVkZsmauIFf8FWbJh9H9H/IKP
30Xedb1/HXbu6AKAR3llP0fekYgV4rWeXL9cthnUvCBzZL98KV6MtzLO7M6nE9rv
eqb00KqF6eM4reN9VniRyGZTc6skUD2cF0Hewa9RaIbI+y2rS7suQheo9WzMDVr8
iIVW3pA8bB+ZYQeWKR04C9vNhrI5s8Co9rN+B2ZiDFsD86Kt/Cyxo4zX95T4a5Ds
uTAJErRI5QCDpzFHMbf/yjJ0WEyztUsxOF7/oXFbJJFQ/xOSuG9xa8emEw8mQGrf
XuUDLIiy2MS8lqq22nS1G1XjlcNxxN2WcaoXjmnkIu+X6SJfjwB0ODkZGDc8peKR
jKvEqu86+dzxrcYpKbUlg9XmzOsBlsaQPRFkK9idLZfG9h5SZ8/tRRN2XJvCuJ2H
GK3wiHGusoxBhHFgxiuGuo2sL4Gw1ImnBQzQieWZlYu9eAGm6w9w1XuRFKYORpUh
hNay0oSrwmAvA926Bz2odFEWG8SfffATaebbDO1oNns+tI1ahxyp/o+38KjwlIfF
mfGMimRgamhf8Q6wqrrvcdTK7xKw8oyhXzV0hh1GJR9zGdfD/M5dhAZqY/DBNt4K
1ZcfoX3fd+WbLCYCqFcEhKAAUU5ZmhhG4EBzJiRx/9tRuzobjoQ2O1Mhz9Mz8ImS
XUXJdxAoUlVurT6AYdrgr8oi9IijoZdv9x2YtG4vOyeO2AOfCY1/rTCmDj9EO85U
b8xb5e0g8R1EULER2vgK+ExvPp8Ox7BrehDqV02NKd+vcv72sDSedJIQoMjyXyHs
NGbXO7vb7lg9797gx5qHsQz/FQePQ+gcZc9KWtOa6ifmDPwA5fVRqEfL9etB/nIo
7cUC8hT36y/0OqncpYRjWgBy5uHmlqiY8M8xJ6ORhBTGMu/fQQCHX85exb+dE5Po
e1PtM/T7hjsTyigZkREe2QHXVOdt5urEwhZD/T5QIAP00yiRQa2D+WklXXPiQZvD
5QOWURANJimJgu/lUxalOo3a9VrVwgDVZK4/Zvu+8ysjwYr6DfpE/LtQRJD0CYOw
/kvc9PgGsajMw3cTR6f2oFpXlyh6lNuTMS1i2AvaW0cAPWn5yelj3l/iX+z3ZJw0
bnV7/c3knBjyKfTZtCqpLA1rRvSth4ESK93qGt8TA8wH1psxoQerrKfK4pWbi+54
vHg5f9UGaYjxmKcr1GKzWH1sHooHv4WE/m6CMiMYmnE0J74PXrl88yGSjuji5deE
xwwqXlnwbiC7LhdhRTtnq6JtnSb1dMsPbWscQZ22pTDZkjymbUZ/Qat/CI7dTQDm
I3sPeUmi+fm6rDM8YYMznoyNBK2S8rhkHxdI9/SUEpxpqP7F1jlE9bnvDXo1wRRx
N01ISa2f3VSiBUJ0+3Gbkigx8f7lMxSJbUEUlIB8Mp5uVsgWbeBxHq1crOFCNneq
pmB+JnffAd+jHdRF6TowgJPjOQCi7q+5o/WY7G7F5ojUhViYzIRqV4bebMhY9S07
3jr1iqWbehw+fYVi+P/mE0IaRUr3YJ0TBYFqXjn1XOA9TqAwSgPTdE+HiX3eTYW3
GmI+n8Cp0sj741D1a2KjSP8PZvdFTbsxo1GgFdLMyOF4chvShKXuzF6nrprbni6z
dmPMm2ani5Y7+0ZI9aZONTVsCNLdmg5o+7bnv/DaYKNaaRjstdmi2oCMJDUDgcPK
Jc4NPuClGOtcWdnIMzMhefA7K0U9Bn0bNSJvVE4bs714Q2aNmS7X1fGOgwoAQ4tc
xK8zj9QK/hT8NaCLu99cdDHytLSpnCD/N3Oxs5diLJsI17u0FMRtaHdCiKGSQ0tw
0kvkzQjZBrGCzuokYsdbec5NwErm2lwZ73knwKK5FOUFYMr4AJgA224lEYX6aQlC
K+jcMlZfeVehq1Wa62Qa5ARmm14y4DwET28zbMuHRo6ghugnuBbCT2pNx4NXvfu7
i4hayGWoqkufHLIDBW1AZeQFVBm5Zc/wJdREJyjRC9AolI0kRs/Y5xRvUIm5bS32
w93oFhxVzCb2pyi4mSPwPby5mM+OdkfdMtHHeTAdvf/L4VVpmCCxh3pnBBCwlHjd
dKYlaUZPA3FMqjRrQM9MSd4MfZYRpm93cFc5nzWDKkZCL/B3AazeueXCl+LiI0nA
4MO6mQwsEIJLtWIop5kWWnqX7hFTFQGwhPCkX2UB8uWfvHWKYPJ8fOvSbhiDalat
G42xzHbfbiCORIRcDtVWWVUz26KcKOtWA+BrrK8ljFQ5U+JXn6TPNR70/OwcKvH3
B06QlbU7WIizaCV7N/IWhIGNZs8YHQfMIVpFTxMcxDfeLH1eZJTsEkUc5zsFWwgb
37YZHACw1SqfDT+LRz0JG24Be0lc8J0szAELFMmAh/WVh8YOHRuhLivBSuYzOinr
xg7LvN5U1qSbs7LM7+OlCex+jACnl9ZE60Uk+R4pHBr4SUlgyNwSwahiy9NY9tM9
H7CIEV4EMJPlLMWb9ROuhuftlwLaeNGpXe0Ll/9/R1AKa+94HrtQiqIsyvysY79E
3zY0E5mX8x7mfvpeU29NXfXdFprcFlDCIzzPAmWv+kB9nvh79h+PKymBadTDWZO3
fz9ajfYRXzPHItNDcSGi6pqpM7AVJ+hGOKxHHug+Kf2yJABglx06/Z7aMAoWdIda
2qd7EVIxzPyo2LhgERbQea9iCcTbJ4ElHwLoMTGxLd5L6AEV/DQ61e4sDbtJiEja
337slud5++t44ef0jnPcytX5ljfPnNH87vDfwNmA1pxRt6OwygS2O4LvuYvHAgmM
D85TPFDeaIkKShZsUvWTixZ6UMBzhk56y/GHQYU4vZi2Xm9GRGVzOrrwIa5WkXmU
VlWLB5jMdb4uttvsWpl2voBd3Q6wCmDPbstH4cX3kAaSNctmHCZGCRQS649jkZ7N
HEYUvOAxA3frWvJzcugPdW6MNc6vKJiHF+99nCv56HcOgmClUgzkRPEQlIPfwpgM
UmcupCXL853Wnza+Gitw/QX4TyUQQ0L3baIWu4ujMBHAPKY3f7vce8XkmwLZuXKC
ZnRKoeAJMrMVbrHTidDH7l+pl9ovJW3Fq9uKuw/GnvFEOjGZaVTndjCEDUiapyIb
qrCpmcmRaagNZV2BCsIJ+LqgzBodLTha7/iKOWFjueCX25Blv86LiKf0FLJfvCDo
Ka3MT3DAU4ALuaXehD+Zd6Vq0DA7iTjCE9ui9rrtJHEjebYKH6QiD1/xwjZ7JIeW
En294vxnwSAYcl/vLwiePg0vCv1a/8aHP0ioAGRtF4wYlqXN3ACgJnbozKe69+61
1DpLo5RK1auqgwSuvsMXUJnxabiK3oLRlkDCeUmkOvGjPMH90YOzm449MY3UXfkJ
fZqRKEsZNkyGJMoYiEKcUAxcCF8l04qzv0AX/pJO4h9I3FzzHslZQpGf47rvP/J0
NZRPKIP+MRHqQrS7aLNfqzL5cGNqMMuEIPg/Cs+pj2j9VmncPy/k8BuV1hgcABq7
7ukTrH1Z4rfABaDP9H9NjDg4iLBnOtQgR+58iTDjE303HOvWk4RiYgLgiHenDJcK
sZJX3ceTrDV3XTKkx+Z1s0FPiI9BFKunAgEzt7nXXraY/1Oe5jk5vLy827ux/E/w
ZdFhTPjDI39RQuyMKgMg4XRKfX+Nl5ueTa/rnU45R+/4PB2vo6U+M8fAnTbA1RF6
Sd/GM3Z00g2YCbSb5DAnw8o0SYkREKWkP9L2/yzBXSEnwLJ1QQfJbpE03LFY316u
3sqQfg4PqvcXLLphZHkf4JsHAk9eBVMopEmfcQdi7OhkbkYO8u9oj7AZ/cQ4dgE2
ULRwVtuZyHibNVvCenIBb6mMRPBrfAHJWZjYcp7tqZiCaruabnzW3ENNiU4/2vXt
5dS/fC3Fk4ysAtRQThKoPecu/HbF9bTU+xv2hkyH7CEKixoMHEKJimMzDqpweLw/
PCtOEDQTpg1qxQk9kPntptl4CeS6ZO9h3fFjWYoZjgQ4JyFtIFHn0BuPfSfXQByY
IUmyNkCaHuTzeGoGEIusKUHushf56C8hHIf9iQWUo8VqEV3Pf/Bkd7P5g0HTgLq2
mvONN6sNzFPVPHVJiI99WFt0bT+hQzJDj9Y+A3VTPBjHdAxvCe+gv8HT3yK8IYrw
lqAS7a5mLR4H3g6Oyr4tn+IBnnFYZNGRukHVujO9vS43XbzHTg5Bp1PuGEd+6uCh
flkxh3KKV9AtLeMUJB03boZch5j6wVtbhjixUTV+TTpJT9TCW8yOnEwPYvyTbUVI
w87P2sxvvsAFVP2jg8DmAdJ0WGwtPlETSe+lxT+UkzLXuHQ252mY8HPUX3/da9fd
mJsg9GvkYup/0Go4sV55ZhGWv+T52hSKx9TorQvijUf3pWH0f0VWALJIZRAv38u4
43/kmKh6k4QCdgiRndXndclFSNgr/9rZs3iuGLgtO2rkekDKvtkHxOzf0mwz+6ty
ViTouEyrafaKGB9c8m1I4F0gytRJ9BdfexpNeDObOzomZxXlChWz3aQsClxx1Uof
SlGUE9Nth26bfVoOp5Lm5eySFb6MbS/R4s9YCyck2JNZuGQfwuLw70tOvJ1V2zdr
2DNlCFUS1gTvzLMBYt6oGi0lQE/m0FxsrsqCU3L86AmfgT/lfckCy8f/7t1f3cSS
7jmbpmBpIEetYytsNth6+Cl672hPrHjI1DVUbSjRvvDWYcYvtuweWjw4e36LTqk5
9CiluFzxVyHEIVvtJL0zlkUu6lTdL3A5xLPJqRKRFbfjg40L02XBaVp9P28qeQ7k
wFS4NSG9rNzBC4ndPuqQb5ds0pLlrRg6Z2pT5GHXUcors6KyQlsfUIMZ9dALZifF
E+uggNdL/Y1iQEBltG1iI1FF7QJsn0Kyf5EURq+wYqkwdk6PCU/5fstCjnvRTxWq
wi9zrVJWiYqqXEXKXBfub8Pj6rBgPP9Y5Ksj1dxFAZgwFpnFWK1MNDjkSFy1oLYC
O2Rjq6Qwb7rB9sAL3RR5BzUixUoC0cNGy78/edPPm8kmdnHfHYNBsHtMZh5JGNiN
1Y7uwZgKZybkbtN44YVX9/sSeTdR2oHt0aJqwuYPJiZb4dcvIMkxBYw2Rg4PJuff
sVvcilHGAEDj8hYchYYE+BlqLaOBSvaMcSu8fv6q9/RX2Ntl03/AeHSkp2RlLbd9
33WdUeGcwBiU+QVTX0bef0jVX5VcOWL+123ZntwhdYFNpoob6rgfGUK+pVKq7EGo
h1reGTRj4HPjlBr7vZ3QiOdDYR5tVrTWN9glgGjJijSkGiOTv3La8+Ok+FBdiKNF
Of2Z7kHn3HI6mJikneQ9eVInNLj/uBCIQ//A7erVRENP6phJSQD5jha6hM9hFi4e
lB+jWJONuedVWlMulftYujMu4i7yhtgu7rTHhmH6aMuDFpYMOxu3GHMfpPHLudQk
iR77MGN14YRlGJ+j38HFm0+rE57hFU15+fX66MNoaBwmTwnRrmRJt11c7RI8jlM3
p4wKmSA4A2yQO1Pd5sBRPs8hzS7VeSOgBp4yltbgx6X38Nxm9tl0m65ZL+3h+DIV
H8Eoc3TXIQeC6CxocoTAyPapsTPe8Irhg/DI3lxfQkWGYSAo4YFlBoj5WnxdY9ZE
IUvgsh08j4p2u0J/FTHJVeajfWcjMw4td1PpRmKuGu+UZb8zUlME7w5H+AHkkRHO
QZEbNwaCQYKq2uHY2RfQvGD4MzoRJu7/gnWdJvxoQ6w7PSuAOYs6fTn36ZQmwf0f
IZnUOWyDC54tt8vgGTMrDZDHhJNaBP4iIGuhW6/Y8+fL95eKeAs4+0K2dM2Hfa6G
t8zrzf0lqQHB4qNf+Zhs5HH8kLx+vbv31G5HFRwcQqbTz1PUwOHARMYafUTPBOxm
SkaZn0d9O03bit9zuk1RXSTP328gHaSt6ois3eanZg/4DerNkrj3pitZZnnMCKfm
q+67AYL9OaIs3V18Ka1gs9vymfIfg8TDeUYMWxu5kCY2cG9eYsfSYXcSsgLf7YOu
jC08dTrIdYZOKzip/uIDoFyGRI69Ye11mmrob4r+EftX5SpmU/25lPmR/ytvP/av
alZEY/z2hOqdEzgwxBYuJ1IiIvdphpVxUkR3B3WcFpMLg6WB0vVDIRLKnMhxRXEr
DZZhrvDCimKjCJBAoPw2X4E1AA32WpokeNidq4bXbz73Bv+3VxZJajNC1qYzubgO
rjWifo6TjoBEG+12QZsHE39zEYFbDYiVpkKJxp3Fc2xuD6pp5g7tmwaXkWxibCE7
3mYKJA/6Q7DxnS7NLdnuBWv2FO/q4HLb1+gPMlgDwgN0lDG+PvgoVnEhJfHaVQPS
zu5L2jyBnTn9ATABVXn+2tKYliPz6B1l4wvXkuR6+y76VfWpwF7/JNhLxs5IZPvl
y0rPO+t0pWbB+DBClG1ZHLVIEY5TPJdKtW6wIp32DrrMlQgnYf+XU+SP0KMQHDXk
Ya4W4kjFq3jHhQOhjkMkOAwvZiL8op25owg6btl7R4phxPQYx4hjyZv3tyXP1jCb
XZb6VZjWBZsgYVJwbQf2C667CsJqtFpePZurxsvFod5HloNXi2z5DwNgpAqjPlgh
VyyFU/3+xRgDpZfjrJ9SJlh5gqCgT1g7lwepWr5hBlTgmernZS265NlZeF0uAP3y
rkl1MIxE0v+bU7rhkRO8Lpt7MT7WJbGcgupx9eH4MgG9/zYIu3YDJlpIHqvrvBrF
6T+SK8zySrOCB7sk7D6OGBbx8lxuLlAu7sYCdnT7MBt9u9SPMmzuUufifeE/KrMj
JKwYQHI7A69gvz4r6skSN7NcOPniPcUnWWajQFObaYfNn0GQ4s8+kfTOT5uLjLC7
hW1Zi+U+GbUJMlQmk5gfFLo48ogKLhDfkEVxSj/gARPwPsPqVHlB3LVHfjiPODGn
1AkGcyqYQMK3bSTHt4I+RaQLp9imht9TMFfStgkaeNZdlD+bimnAiU2pdTQwfzj8
MJjOwY3HXkVaNfEuJ1IATG91QC8J4jupTDvqyvqpCGPMwZ8FPs6CblfAHOjSoTKE
2gvxi1HX3r08qEnG3/zWjKDuj5JLxcW0AaYO3EfUCgRitYc/lZtYUTdeLrS6FBEg
8iNT/hXbDdOBLfhF2ow4qZDU9whbzeh/Wk8FMI82wGtVxo4L7oEUxavFF5wNczWr
GrAj/SG/Pwn3DnnJd1moF27Yf+7+BA3iko9iyTwULZL3HsXsdDnb9NUXiayNJV3r
rcnhBJzgkTmR2Vp5Ds5yvKTbgostZ4hSsqLq6GvgUBp5KcFWcLu6k0uArJ4M/A2f
RgD7rZhG5dfXQu7jburO28tD2thAiXhs4U/wAPBzCB3fId3pOyCBX3Kb8t5BnHBS
/RwT3nPqbuTmfZX1lexJbN3vgKpurr6DL51klCoyoF98A55dSa2IeFYiQaZZGhxt
UERadzEv99P/Zp+vF8ctgWWt7GRl/rNQV5b0AKeB01YdsEjfoUhOrFMXVSorw/ak
ly73vDGDaNqB8+1lMEtx4laTR+l1dRKXGnH+oSA4y2yM4yOBuNt0H4Df/wHDoVjJ
C+NnBc3X9Z2ZBpJON8F93S9/8YQb/gEFcRJHjHnMG5aXX1mqbBt5gbZgMDfJZIVs
/5a3wTkQcqovUsGCaiOh8YslaPolApzNjf59k37sb4jldPsMG4HLT8pSnVD2bMR6
gsj87yzlIqJc3FdsPNYnMkBEgoOz7krQC2XWOp5EU9xCMZ7s3hOZlLzi+0U57ZC1
iEM6SGO7Y2++/JDugX/D9za2G7VLZo1xvd2HschZ1rqDltQniwo+BVmuNNfF755E
tJu0ZpQxM5VxDBr1ZtvbbRZVpl2Qf8hvr2qeq/nLr36SR8bgNdEfIcuK6ET5TWGC
kE852usoiZlWwSONlwLnypFcvfPcW+UVZ2J7M3OErTC3D3/y+o93Mxhxs964QqnS
c4BQUgTonJ416k2uwtf9+zCG6nGOHgtmjY+A9pDh1zMh2NDLSlBwWjNyykFgyg7g
oknVo3XdchJ9XD721jsHH9cs4+N7SdQ9rhWTg8IjFlpfnPM2Zf0qmhdT8l5jzAm8
d4nMekK0erxvso5QQYrGftj11+AMWoeIvtC0M4ga0d9lM0r9ijmi4HypTwuFCMbr
SS19KIRfVU+McDtIB1JyegJpMop4vgTSPGs7xTniNB+a6OhnL+fYDKrT0sA27MQj
0tJW8T7jRz44Dh23wdd8J1rYItdQFA19otaQ4YLMuj1oFuXo/cr0AZbqE9uyhGIt
LQykXoOWmc/v6KhdjNkCu6r58PBiL3pwSq4flwQpQvR20+hjkw3l3fwpMED4xxln
zh7OxKj2vdiZIbFF3AacOR//AT818WSETl8okrO7gjtGm0OzSH12wIHAQy6hMZnt
51cYoS2En9XmPQxJYX1jDWFYYwhZOu9sHHDZtsQhWtFDAw0TOMhUI5OYXmAc4/b/
Ro6NDiY/3vcLfj545bNDhDNZQkaOj6qpTNVbMI+FZhIn3qL5JmIROfyIK+wuOxJk
qO2MX7fphCM3HzoynHzOvzt0867HQdZzE4EXC/GXn5mo5JIt9YG9VTGWZ/3MoXyR
BBrU5dsWTRXSB8TPJcd6tA1Ijzq1NTa6oZsq7HIKSt9j37y1WGzPqyKy+z7eN55B
bKiS7dKFrlNUJcZ9ocvUxZ/bY37iQK1DkvXsYsX6qCw1Ag5/Im/c0XvgOACncVGx
R37qR62iXpkAhZSUa1np0B1+CLPm8NIUs5YYlSdrFUO/NpfW2lP3M5RdQhH8voyh
OWig10WMvK9IkDcoLFhTXqQos1B2FhzWCGiKHOUuCvLaWiMWQQWJqcT2KqzUwXxR
0kA9uR2ZyzybAZACU8XhTb1khDj4vQU1SRIY0Y9UhT6mZ2/NX+nnmMlqhA6L6mCT
3Zzc4t2K/jlNLOgRGEq+SMI3Juiu69GDfP3wXQWu5MCODm/jO/x5nhBgm2ZpbRx2
IIafbfZhyx128cwn2PvbkIQt8wH5hT9MSEr3r7nYpEXdbvmSClKXa+ip2s3NyGyT
eFnG8x4VqjmtigXI2+/WAfH0sy4g94qn/4/h/MuMjB5cVvn+YAvEfmNIzHkRZpcZ
nzt8iapovdt49x1NSE+EHW0ePzbOXk51n/as8sSuuG27pXw/YSrpPgNDWMZS/aPF
pQHY/8KMRUwjkNl77vpgwSxRDdHnXl8lNZG3wZsZoyWl9w9xoaqWVPOD1Z2rpWuE
n+1jmDTi1bYvn+KJ5B7lQIDdP4wToSYaU7ayLU6mp+XKS/xq++QOL+Vjo49b1Cqm
fkUKNiT7iSAVmQCByBrDkeOqONzr+ZQXf2esw62ZU97IMK0ZLHQKQojseEkz/rKM
Y3djOBE5pBVN5eyDUpvYkA0KQM2YrHaVxVkQKyH74p5hEv0BGt6HPiy6kj8o1j2V
+FsU5VOif5yUB9OyPP21oFush+MmtTAze3u5mSmDI10T1A678PtaaTLO5nmOb6MF
Hhi5jkSLwRYx6BtcpyVFIreq5cNY6KstKZNv5V7FhEQ80sNxsh0lR/mWXvDU0mJU
mO9PYG/3J4tl0l/qnuHoRXBxDX4miD2z0vsdTuzWeNIBhvyL5bVUJ1npeppehREG
HzNNLAf3DmJPRD3c+Zk5FxdYcE8h5CEtMKdt/Qtm7auNKUDrUzTiXPkYty76DX5w
Ia+ps0uf2kPdTC+q463FMoEX0F68yaiaOcEL7dxm6/41UQ2DxBC+V4YfBenEJkz4
/c09riaBlHIf9lljgIoBHA9oNNDeR+gxDg2Mh1YgKjt8gYeit5JyjUjTrjudVEki
m6NSpepYeNjblr9qSq1rKJ5eihNu2kidjtMJmFUuCcSH12Qzqi7s1HiQsjTeIOEs
mZU9fUCZB418NQb98MsHO9ywGEv+P2zjY9yYf+9cI+PTbZgLe6I2uR6NAHVIyM/n
4T4LWX+z03ShPeMIghFWc9gqcaqykcn3/bHTGMFExt805agnp5GXpv1RX37xKFFX
MsYinnRrRSeyuP0yEUVJejj6F0ubGnru33tmhQ+GbaS+C74OxZeaJyMBxdEHVWvB
CytAfGwwT3jGmogbjIl1ZGUJ4DLCddpBvoDZteti1wikDbIMpR9pgaC1D6t1FAu3
ayCeowotfuY3dYMyN6FZcHTZDubxVkBn5BYL4p1l/m2AU9QqAjQyxatWxPq6oEr5
LKaLsQfxWs9pWsvpWVH4iibIfDzdf2hpGYAkpe5pwIo3kT63yQf8DK5ifnVP1Yl8
CwNjBkz/4zJ7jKPrc7jIWr9PMLipZ20y15ReJpf/HW1w/uAzxCrG5TeKlaQjU+jq
mtncUdJNNHjitX6nOsnsi1uVgkc1MgRZX9WGBkSHhql9u5OnS6AYZw4WPvH5AP2O
9AFMafrqmS2NH1k3eD+/jgARiGWpM7ALNfQOmn4AhyzV0hmyn8n6ZIsT41Phdcbj
eq0Kjy7nC0YxeJXNtsPZQZz+4tvW/MVCnQlly2N92pxd3anHCNg0BpyZHMtaEvdC
G6nrtiEgFVf8KEvyTgElek62T6h2MXlZCtCSG2ZYB1vK160hkjaHq/mV+qPwHfoy
TxOh59y2DCyQB2oJQD4cTM26b8dolQSxlPDI+6iin5tFh9W9u7yHKk7XxL6Dl7yp
Uk/nUy1CvjymqLz3KYd/JYRl9PmnrDyrUUWGvvFG7uMw11wqmWY3nh9lUbiBVTVX
wFwZcPNmL3sqA+KaGjOCnYW+O8ZZNRiSmGoaGGtr8tWzbs0MW/JMnIk7GTHN1VLJ
C1J8GoaCqi2Ln0dLGd0H3Sr7Ky2G3c8s3YexrDypFZGJ2WI6QJduOSGPU7RYi4cv
eTmG0QZ7o7uBxYqSiFxCISASEJMiVzUmjbfYTHzdaM7HTW66PXgCIrXihtxHcqBg
soKC61cZRO91kyZ/exAHyqLdQboVQjPxil8lgnJ/jWZ98z+Bg5TkJtMyYwnUcNXm
yvaP1IJ8QichxqLo/UOY1M6CEKd9IX0/Ri7CB1cAr0AYmFlWzwiHdPC/qXl3TyCM
kBe5EmAzfkZDEnzWKYfrxeAyGJSzWZf21IqnVE2DXUEq3xYV4rdC5JR69NP9EmMY
M8tuRSx2P/HelmpPA7Wv35iW66bff5yMjfCL44sul38DLuWgynIi0dC/BAHwuKjC
bfuYJ04zC7MkuQlnpySbnAha6Bb9LpkRNIkVsS0+b4ws1e66S5aJVMnMXP1+ufwj
MKOlkW3igzSdfYw3YI+YrY6pGB6DNZO5GCPHnsGJViuT5qkB0VxpO+k5Z5sdffwM
dwGDWbrGVRO+da64FWYa6BmVPl1gkYuI/QpFro6dKJVU+qym6+CMZQwxvxAWmAOE
r+TsKA+ZnwDDPGMUCF6zSx3lb3SNglgR5SyydQEFNdBOzLxooulZ9I7OeIPmsWLE
AVSe14eJDjmGmlJd6vo3EAF2pNRVI4TCtmJfn8zDWeoDnhn6zTSLTemYh00CSUIj
UqcvwpvSMsQ3BKjwqjS5K2imkN9ygmhylV47dFRpwDKWGFSDnLpMAxMaiYchVuJ7
6saUwyjMJ/Bly6+QScG+kP9BgbAiHEDG02aAVvyK2bqJPKpKYdzwjknDBbtQ1d4i
Lf9sLf3n7/OjNwxE20ilRs4vtksEPnXLjIE0Xvpxi3wn8AkxwIfgESZ/mIciUQuC
eJji74rKaZQWVBbr40v3rGr4RlIH7i7zxsp7lijCMhXZWDvo8+aG+ZkDb+0MfUEE
6F1dL26UFZOVy7uPPe2cW/W2aQMmL34GHg+7jxvPA5ETS6FlNE0u6PYktonPIs9Z
3gKRUonJg9Qtvd6OwydoWqyWGDVkvYbgW/7v6zndo6mPXZ4vY1z0TP4Hl8uHHjyk
Rlx7y9PnPXQ2FyXZyJWKPklJCujH8GqBcAljroPvcnitlw20z874egdj5nnyesDx
W5G3f7kIlz8x36PTgV9P+8wA0M6n5rbCy3QL6RoLTzSq1WT2DfvLWMvtB0fu+wTD
4HtXLQmB7S1bz13i0vTD27zjP2jN6uQIX+BDhk1Of9Dd3BhgVUsQKqnEtXfvMgOI
whVRIzJr5rTJOfBOUb2EDoq70epaajLzYwF/Q/GvgxaSksWK3rZdqJg9nNjKpLU+
D+nk7aRU/msgL450lsQO1MFqLu8ZXla7QNMqI7Atlkr6merNooOh7OFxxn33O6xp
BKO2suggEVj5JKqv8lTMuAllnwQZYNoZdINq6IMhmKOr4rsJTxjj1DwH+3vn0sWO
8hEIveyLdReQF08IBXLnB9ttF4TcApAC1UfF+T5IsEtJqejY7Nsx7bKuTuNwnYkA
8/jdwpVFc7p4dHBjYGODc2cTeLIJ7LmeoXk/LTm06DqEJYWMS3H4kS6g3zmn8xkV
syHq3rdu2+OQZUVgrk0omRpn22X2C3MPIKhlVuMeBTJy7twSbBiBdfAjyiXc1Vsz
CzOBCRYR/AP1oV/gJcyHxOtX03uPBAp8YYoBr/aM+NR3rDX+thVMqJu8EUg9BKVf
UIDp2CPEMieacLjSpgjrq5XhWfOcvJqZa/rR83+5UzZpXnZN5I0yhPiaVU7pPQT3
+9k4vMqRXHI6OYrtISSKs9mIYvn6ew4PbEesQazCS+z8//w6lfseqdx3eusv/5zS
+aK2kiy42OrpYT2M2NS1Iz/gRIw6H8tz1h9s1EGZG7jSJUJaq3EqNTqLfQoqa10/
ytCyUW7vwIa8x/J/SPdUg3+jUHTmKX1EpUjCre8jomYtho9dwKqf8kf6xM0fGaCC
R90bJCQDRli8Wl18OeUviq3Xi3IER15/Tci6P3GPWDtrsPe/uPC3hRH7rIpjK6er
Y76d2V+sFmaA+A5SIfYNpwGIYagALxWSFiZ7AAoYeS7kxzuECQ6X1EGly3sx7PvX
g8gD3gBQ0BBtaQ1RuNxq1FKZyDmHIdZCUDlsrBsZV6fWqWDXjqLCcDDegwwQC3Fq
uxCsGdbg/UCJq47czF1XuUIi3nieCk29bnN/PjprJAzUdY/Qg5qWWr9l5H7aH5CR
v31/uA70MXZ/wCQFoEjyHDqh7ddIdATuqZ5PWx5ha8/8Gmi0GWCpEK9j+TBzr+QK
cAy6E5PzNs4jLFwcCLIW1/MxO8qv3uSMcDV7qOEg/kpidgqEluS4XSu2ARopUcGS
jjE36WB2Ymc9x+p/3RKJ/8TR20lcSt4Sv0DAXKEoBk00sCpj1PrzjMh2ms3equea
KNgdYj2KfYABWjX58EXO9Y1fqSavMzCHJ29VM+8AOJIofTuMVJynd4LTxmX9QYc6
E/oU+EBn93pC8JIwJXf7r+KOhJ+4S5ULB3O3lvnSt7SHNRnClXBA+65awXXPo2Rv
0EqVvhF6GYRON9Zb7lYg+g7Ws7fdbdCdIoPkaFyRnKS/Fpjo7DQkVY9b7GjB5h2v
rxR3KzDokl8bOKe1t1RX2Al/ATXIIDlc8i+JYJurdrrAVH6R+d2yslOhPr6BaQHj
0C+JMbswMrJR1Ka40+H7tgxW1Kq5cPHEOIP7JukWhodlGJa7FzyWw787dsTwOhw5
FQaOD1LXX5cUGkoLdE93sj/jt/m3r3yjU++KT9RnRkuRAsFD4ph5QkoiCzT+5ME8
WlHXDxKCGoRKfZqHuJJrAqCyynQbLcz53lHKxhmWeNrGjVVFi4yQl1u2cJ+xilzB
03R7WV5dbyPeVmw+y3d37vjIqzCh1GyEFUwHWxd2GP8U7Vl/I7PPEEZVf2wKgflt
ihRxVTpGX0afqJvV8lUEMYBNwH8IfXa7oeQVmMJp92tFpPM4CU5B505PqKRTIO1F
ifJQPiSWzYwur4IdtYeJ6198dlVZfoYcVilvigvKrC1V8qZxd9e71sL/I03N5S8+
XwHJFucpySd37euufjGYIgyRj7RFsrXsvmg52rFVYGNflyKYkqGPlwqoelhMEZGR
DJeIQ1cYmmFc2gte9E+RtZfJ9mta916sW1iBYZgwIg26ImYNP+6m8hjbV2H14G+V
P1FzHSLybx2X5tlPn44s9XFZM5aeW7vn4gbl5dIjdwivhutIYJG1A248ZRJ831re
Vfk3cYtIRgsU52zLBAE7wJlgU5GC5FgdNP8evcmifuOtLchHJTDyX+Cio/fJqZMz
pllI72SWPnBGtfG5z/zasJcDCRt4SfAawf3qQzTLlMlVD4Yt0JQiMAg/wrdnbOyx
SB+758RryngEJZOU32X3afPQVh952VAIaQfG2TG7WuP9T3hgYGdDACq3aHGiAfiv
8y1VZYiT3vysYbPt2Q4cKt7Y3V6qP72W8rxTeHwrMRcy2uBD3vXpFU9VQ0DuYmBp
rUgN0jythZoFz97uPLV/hEtAG2ABqnUTTBuhiPzWcrZpZwcWcY+Y+WQRzC9MB7GT
VE5G7ASgtpmeLoFNz0n5pK/Qrzbu8nZPBzcqAQnzFJZ3bGIeHPYujhm5yLXAM59P
VE8hLWcfRSr5RkaxIj6pjKSXmmm9erCNmdNnJu4UtBAYuT0VVXGb8dlF3Pfnf9bx
/W3DHy9z+/Kq4jrse35qPML3kcbzG8EZhbGuCJZaS2JtfJ9SXdqbM4DN2QJ0VRj9
jgV74CY8MuSKM3OiQgsfsOuZMbVHEg9nol+A5NTdMk9yYr/I1fYBer7pSP5iDKvR
QMFcEN6kVe1fHppOhjI6JxRZTq6Nvytog9bdrtVpXVNJUbL577wf3qosBK/SaX1h
TlRrUZHkdGwAiWdJJUgZCS2F6xNe07uWKSrzvQxQgXIRsi34L2bnv2L/R/8Np9D4
nciVcy9yd1edAMAx+bPuZaBgKOJWMU5O5RsteUQkYN9wc9CrEI8IFlsvtWlgRT0b
kv7HTSu0rjMUKFfKkUs9zr9DvHaI3lpMKXx+DQ3gvnlxw33OFazRChMMRj/fCfLP
JpxJpnrc/SNMjN+ebGGkBZkrzMtQwSvYKe40f2WPPV3RPi8myuDmzD9CGXCnkyxt
JOAT7DEaK/92eUtnO7ZieOpZUyS0t8nDqbCcpCaKcpmEOs7KXmcqbZt5Q0l9qRNN
rZrBAXcIvFaMV2s0IGdFQEvfHU3R1taRR23sgQQG6TGcK/gTT74khmDwglTgYzRu
VUH60MeAlXvs+nl6PgSLyxKFn58ggqjd8oY/xvQr0aOA273l+r8NBrrbbRzvXg5T
gNBljVuC4MWWGToJeyhvAchSbwfYGe/As6x4fZSvhDwcZKy7JQVA9cpUcAWy8HiC
FqvaCboBMmXt9KjyH+I8ZDAm82zC8qn2AK3AVspUaOtVTTPexeXMXFiYMAneWcaH
8CyTvTVvU7vFHjwxerPiFfEMKHM4wJ7GDOl25DfWmDNgncUTKY+ndqmtZZA9Ah6a
c0SCilVHz15X+EvuKxcyCyemw5NdvyhXvIh8lnteTKu/R0Q41fLhdxDQ8muBMooc
jXJKpW2nvKSNQ6yWq8s6sPn8tkF/gYVloT3khVq66lpDul/h3IPQK2sOak+kjC8o
BaibiyqcQePyhLsqWDYFGa0uiCv/s6KYZ9SMXgSMib6OwaTdf2d2oLRNLXbp7+3K
aZh6M5Go4ubgM2Q3oAwGIo2EBDjeLyKTZJv9nQBopM9BB2IXEAWnYENYVBG7lhsc
bqU8+Lpt+rqVHt/PUs2tL58/90nbjx5neOQ+idyRUydTlml8QJsDJyK9AUUPMVOy
FBcqz9l5xPxT7XeCk9G2zxSdQDy5hsLSU/h5dyGM+2N8Db7jD014KPyjwMxDHr2Z
6r2AY0gIPoVN77gdGry9kM0q6HPqzMYNymnItj8LtUqQ/JFn0QM1nspVdU8kca7C
ZFo6Jn/864hF18g6UmmLifj4oJ2QXzIOKcEG0+luttzA6bUTaJuLrVKt19WMwl1K
7uSpBG3saTyPslY4qhrsHtOSzUoSx2bF2IxqKDyjzGtjJDIpY1FNGOAEr7Vccgid
p8GR0IeTY11DTqPuHAHKPP5g+EeIymxQXXS1SIu6YF8NfNhb6E9TM+jpcObKgj44
/lU1TauP9jivLyl+EjpgaU4h6WDujIlRdunczrRFbnT31H5qJVVYWQ+JkGdhyesG
Ud/0pyg9GIOH7RXUU6Mj4RdSUMAOYPthOS0Wpf3+QyQhaSJvYkbrZcpi/jiVcblK
9RptxJIBSsCbItHmRYzgyG6LuWwszNianVDjDsd2l6HYOwh79A3BkMoKrMLfgIK0
9BsneaTlpUJ9Yqh1ccIZ4dxeDa4S1G2kYVepwwL8wL8/LuMjbxXODQ4378AH+YzZ
HDVkdtku9WfTLRljyplrB0+DWuO2ws4x3wkHHLpcIuNt5vxVCKR2Oj4z6/ZxvjvV
/2bwGvBGo5Frdt31q30o0FjyJ4rWunlBcM3t4xzYNF3rkjBqqkOhv2xW5DLBB64D
5J3jmHCjHDqW1bvMx9DZe2HzF2rst+b4Pkje2QwSqay6n3l3Ju7NIS7vCWpwKR/z
jEbX9IoZNmGuzXkI6v8VSIUmervYkrLenl2ilWf1Gq8MTWefImNb1bisDSgXfCwN
DT8aFFvvFajPXKd0OizHRuy84noGoJqT32yUHb/anjwhAiK/QWBskygN+6ZPonRo
/sMzukq8+Db/vyARYXTRlG3qy5n1nhj1I7H27dUiJBLPtZsY8IP5lZ4XH3Phzk2y
HjwcMVOu+5voEbrS/1R2cp+bVE2gXQ60qIZthoGTjJQq5ODPBqC0EBgT8EHfqgip
hNorLjf2KrL4S/UMoQBl5bPsM+u2XpWtP4kWr6HYVI6iXx0T92KppDQPloW0wY6O
yO7wOWL3x4q5TDoB5GSw5tHx+WQnRT8BZB3m5nR2DyXIXV0Ny2H8hQMC0AZgBYmy
/w9kiEtmLKGz4o+/2iR/pxfzZ0351n1wxBSs0Bqun4/gvnD307Tndg0m4vuAhRp9
170pQ5wdgAOkTJ31khGSHM0xbcTq4W8ZPBb+90EhL+56z60FSM5Z2Cf6nb858XcT
wERZKOmi6HBoNMgmeZA925JR1+Ds5RILx9lf/KjeCEOEE/ejRsDeAPiljUnv9+gE
P4HRGrCcPqsy9Uy60TWgtQ3VUhFSyykWksA1R4iFO9QQl2PUkldr5vurG+6EcMOg
zKzcbsYQBoF/dOIwS/oM/H543x52P0wZCCPw5oyO8vOHDS6hJiFfdmN4fqkh43C3
gMMa3cpFWGozh7QMQdiGj91KaMNmom9Ol3paqs1H9bnY6ELPhQ/UJ4yd9v1RYDMB
qndEnGmrmzXtSoLz3Cvd9fB2AmDSLDfzGrW7OzdigCRDhAXVKLBA/Yj+vEQyGOxw
OWOPWHaH5GkIqFluSpgRcYYHys02ehrhXwFSxDIPJKyS6rJGchjjuO6WNWsmNnfT
XOTjJqBTFGrTSgEjvPu+//2sfm7F4sST7d/eikObUDsi7vWedXpP1MmjOjWFyDeH
2F4LneHkT4ZmFbVCa8U872P8l6aeAu9GCcDsSeSDP8FiR49RIMQVCtUWTvzbpYHt
qB53FlmNiWd2t+g1/Mgx1IYbLdhNsCe1oaRQ12PL3jrLBfB5SzUajYLPElPJ7mB0
fdvmtQzepaDJXy2BUfxBPeXNxcG7mAO+ituv69d6o7ABKekvXGkhfZcB7tH2GulK
Jh+4K9p35k39uN3phIR9RFqsAoOEbbNEqvwEz47Be5AuyQ5eKcxsRXPj2OzamudM
a2aO1s9LywXSLMThZxtWcTbtPEXqw0Mlibv3i/5Ny20NITYWonwiPDvgAftbh2WZ
PFXYADJ7qAK03y4bChNpsWp4/OPeTSvpR+5Xm2QJILtf3durobhjWPrkxcBaJKUZ
lynpE4pwB8Pv9APNCkRlM+9NHTuOlOpWa4wvYTEVzH9NedEsC6vsmYPGFdTJVpcB
RUesoAKHupnCMXkr4L+KY+v2H/F9cBwfAuiO5ZQykQpwZBK3NpS29/nKgD8vF6kZ
PFaDVZ0v85inHbZyl0ElHlcAp7OqgBKqaFN0jnJapf/S3f8Mai/qTM1V7ZSLtCcP
PFyJKBYShAHx3IER2WBGatccFs1WgXgQKmLWN6xFeYj7AsbgFvW0UUuMOgxu4MPd
fJ1It97eUvj0uvY5sCYQD1JxrdzSk/hXWcDKo8omO0aO564dBGyxXYa6WkA8ntKI
mOXK2NKk7eHTDQ6KFmMnN731BOjxrWmfJiV0tt8W//MuR9xMCQY4jGyH0GbA8l+Q
VO2ZAzF1+IuiyYq13r02imQq7+NgwdEoSjXNr/hB0h7+ti/Kso3vYQJrmRJ0OQUW
8U1dRQJjnvn3ShJbnv5PD+CEEl1xoSZ9rXKpG5eVNNZwuPRAifn58EdaxBmvPC5t
Kfr4sx1zbz7O9jq8HXqjtm2E9LZ9TRp/Kt0jDOYAy0t1NB8L98fHdKl1r4hrKNlD
0Wi2EShNpip1oe31yNSvUuvID9uhF2vjx3S7a4b4N22/B0d0ZOhi+FjzlVh53I5D
KQw7pnTCjcQh41HflNxKnY5AaGiLFiRRl63VLnXS53tOwdr//bi81ptr1/VAZkVJ
d9YelPOXZt1OSWNLF4ikl0Bx6/tSJ0Eyvc5wM1ri4nbnRUYKHGubM1B/U6IDehAt
n1hs2HCSCL4pGDTHvD7LM03I3o2aGs/IC+dXWu6lFnD30MlaICe1gST5L5Tpr+Yd
hiSDF9qtRLblhxWxBtRCtQ9d2D36KTvS7rI8ZujckRlyJksTnc69Q6lUX+fCJ7UM
qOW646dkMv7tlVwg2ASBv46kjaSkHNEo+ok+Fqe4jslDvAFiXMTJij/23bNRQozt
BZOui/nNW7OFWf/0vzFQm8oCOpuYu61pzwavS1q8r8RdLl+F+Qf9veVgZL3Vm0Qg
5FwzJBMu1co/xtJT/UvMSYBZji3027vyqmfN5B80hu+/j+8sG4N5fc6H0Z4JRfRm
KbsR1kYi5UbFgihVym9WzcfJuS9/ZqY+gAJdqfaqJKesQtkKwfhVu8sPIO9E/Wxl
TFCc9i1k8KHzKh/aiIPz+Gt5yAKcK+RzrASkyZTpk3mpGmlAbTffbrzpe2rnP/WJ
Sh4k895Jx3O8uUBFrhjQfKJfLVwW3EDQY+JwDdJkJhsvBu26gk9xUUDGzzYV9mw2
N6BjRVBPhOTT4QUkO8DJPjfSOSJd3JNeEeqad01dsXNxVSFc0WE1/HzOnJy3EeNF
okDjaFZzku4G/l5cYT6W1nnrECrJbRmfpfUQxjYMKztILlCTxs7CTHQJS/VT1nng
dhlx2/4/nRg3ZSEf+oFRgP1n//q8wJTCMYoJEz9I8wPNtfQQ3t+ZdaDW3JLu8oCr
t0qZTpX7HJnA0Sk4HfZ9wVXCRgkiNqEPWIpOsbA4gNjXC1sw00wtyATK2z0c2oki
y21wPBUNGiH7JPvh3M05RDnJBy3XrBnDaS+Z8Krwld/7/aoSc2rdoNP/2CWbf4cx
geXy2rb4f+k7P+jts4NwBFZ+MkIXCHCi6lX22+1gzX1Xrxedlo6wvVpkh245X+XA
eX0g/aRc2l8XlmGNYqwL6gw9hzvIcNH9RZtN48oKYhTt/sqc2mYaT1MnqYA4Djzr
0en8t5E5HZVIxooAx6ZrOwmsYND+opxaE3JDbYdd4CCMv0q2xltv5mjvPH00Js9k
qRYRf4HPQWr1oYCd8mhN3CzrqmMm6ld85lGShEybqBr/HgQwy2eLeQFw0ZlohdeO
FOlVw+ORD9GuqRR1A69nSCx+DaM+lvDQOKCubfOG/bsaydaCoXBU6YQAqD2f7iZO
LPeAWW8wBZjbO1jLGR2K2OXhcBYQI44cCqU1Zul+RpjCqpgU2MJ7hvZ0mG0eysi7
FeNP9gJs5QcLPNkI5YUI+8bahP/7LSWZ0gYMMjAUAaRB/3yX9cUFmO5ZOw/r2lO8
GA0j5glyBjJANx1EE0j/bW0DmnRj0ZQ2fYYWoZwm2ScswdsuBO8aWw88LbB2D8De
hQ6w2eiuheqJd5Be0rJAoYg/a0/XH+SF5eET7CBrOJPAsAwp3+Ki3ztERs0mTGqd
g1irssPoJpoCH02W3cSGbqyBgo9c7eTjw/3AMrbUsQL5kRuBOJRsUpgimV1ZqpeD
8E1QzJS5KSxe+D+7oQILr5QQBm01W+qSF7uROf6SaUgbO3MlxKRm83BeUY7kGoUt
A6jCkxpCW6DB2FAdCPqnJtNTNpRjzGLB3LHTAQG47NTdKeKQ9GN2/tu8pEXgUEuV
DINNtOsRPOYofgcZLTTjQ0IpzFp5i+2CzH1ddAExTfPFvPqaDPop8dKfrccv/ebs
A5zpvv1NFViAE741VhAUFUq3xKaL+l+8XkEcl0/pw9ddbCX69xe1ahR6GxNVwkJg
etmSbrNAnpp42u7AZ6U+jD2EHXQvM1hXGGMvo5aQ9IgMIGpYnJW/HI7SdBtticVE
A7Xmm9l46AQvvivRT67LychhdSetegFhlOdMPI9GifPf3/FtayF6QpUPEYaQB4GO
BMs3qaot4W7DvCVamuPKTg3bTJYPaY/N+VG8gLUDdkEWnyWvaovfenaGurumdKAY
65QiR5kMNpcaCquN3hmB9AHuUhKd9HlTzHlBo2HU6hAXwvWYUmsXWIYJ6Y7Jyh/B
I3WrXSuv56S1y/DsQ0ESlMghZYGR3MIlt/Rqn2AyOF/BIFf7HQeFCpj5cSdEJJtj
2/lKWhpSLd7ss/AN4WH2zUyFGZ4/B5PI/R7XGD1sgCDXiizrCAzo78pZCHAwdzN+
714hiKR0IB52ig6UIa7NC1jclsn3FHgwF+svN6CGadl8x2gkPdlKtO7GJGCc4Rdx
mvA260MyPTHSCqsx86T2NExYqqX1X3uZE1f8O7ETOE3dU+xwxrJ2I9anGe/5xPW6
QM5/5VGRAc7mhEmXyGctfNuhjffwFG9UBKd7lOSqs3JCkdJiKZ3l8nsKNFrWQMJS
3bVGkHGYs8vkfjSpM9XBeLsq2A9rFWHmuZPyMGerWnGa6Wi+ss0DV5MikXDlWbFg
GygHmjPZ3a6J9Hhz5ErPz+sg82VGxL5Ibpyb60OwShsTcxEWSEHcZbert3Xqe/5x
Me7fBzQA1ylBGw4Dg8IaEvHQZ6vtoh+EmOE4ioUxVHls5jkouMxXl5tI1HUfimp8
4RhhCpbkUMLBnayR8yKSTUDQ1vs0y3SCvHSie1m5puCFyCO9OSpJ8lofSGF2/ya4
sJv2vg6rVV+iySa+b2akcKf8iWILePF52mEoJ4KZx09aTsjFwUTwMrh6/Kb0VzLo
WKEftXQrdiOeG3ANdmI49wFG2baosJfs7DzrzY0E28/Mk7wq58/bzMv9xMDOoGwS
Pzm+F1oOBd2ffUIzFnjXZ/0rtwrSPnUR+l0wBaNKhY6OVh0ttEdzQkqv3zJQuGLd
YZ51hBBQ08ZbUNAexeZws2o3Uv9XYkdV8qfdJKF2PuHp8hAf3q32E/Gx29olPARF
yc6bcVIr73TygbUqOKzWmWvxQErD8nAWkBeEhJ7MGCswDS0vluEX+oU2xdC1Yjt1
qJiAsQh8qwhzxLgQDPnAI80aNzEZoksfkAHpkl9oobjZF/32sySew8tuTAcPcMOE
Le5tM6Ef5JZVO9PLz+FJtLObzDhVe+LQQgikVSNLRCfizrXAI4nur5viOuwaLojD
QyU2Yw+jZuFbnVS3VBY+NiB7bvRv9qzqClLol7Uv2DUVQ9UT7YHT+lWXkBPdT7sy
iSb7SW3MWyeCo2xFtn6FbLwZrC1Z7GMKQmjK38R8YBLjhpiD5pZhsLnU/AelhMw9
QUGed0FU1cDV8T7jt1oRfprUpqGXFG23hlRsC/JkZfOKOdWkx/9OwR0h+rF8obj5
/4fWa13jOXcPbTuN/+2wIGmkMOZF7oH1nrsXYOVkKT4PFlPo2xfwgMKgdYThhMPE
J/xJ3JSbzK3oZGlorAGV6fGISiJTM9veT1d/KdEUPXSuSnOQVp7OFJM2FfTYV+he
ntJn+p+DvXgcOZu4anqP0ix7UvEmQ9eGk35Vjtc+27AcpRWdpS8N8oVjdEhYRUvJ
/HIkWMSpGvAaHekg1UuqqmSXdRQaN/TM4je5hQKORxWdVeMvmT6q32xUB86Qkl+K
ysAgIF4SU5SDqAbOCUr9PJX7+vjRltG84DJ17wGVtrtxtFXosgZ29pPYOhLdD9zZ
URchQtP5L+Nq9ZbptLGfGHodsOQAFm3fghwi4mI1WHomjrbN0b0jz3rX9DdzRI5Q
p6Fse6WNIKMT4eHM+27G5WMq2dSPNNXX6+4YSql5wxiLBJG3XvOt1s2AsqlvVPbE
TtHeMKVJiIpnjen11yjiB99N4DKmkYsKhcfSKoRo/RvvnJgLArCuTPlUZht1YdDv
uGZfpkGglapQBfFNZCbBguUYgX1igN5G/ROlL3V6ce7fk/i33Jq01j+BELTjcfRD
AzhQGymUdjDVes/6yl3w40fPkvx4nIr1zN5QVA14VuiSbCQTw8EZnnpzkWnufmsD
w8Q0wu6K6RuKAXDFhmWC9tfC9QIL3RdJOyA4LojDBaMwe+fBZ2uBfOomhKPKUcyM
x1vutqOA3fiH6MwnAQGNwyjigU/4qeCvY9ibjimisJJEq9jrbYTI/ICvKL8mn92Q
Roz4zAXTve85JmJpYQd+z2tXR21RSejAY3rFO1OxJDwbExGc42d/oeM2cO8YMH/x
MhOkaPjKDzXODEepwlYW1Idac2tYgRT1puXsD8kHtNJViUVEAzBDXmqGRYSEkX3Y
pwVTI1u+TJ1SuSvBj5/EF2sO1gz7dMbXUgh/8MFvz3RCt1wiOzGC+Hv+PUTYFD3V
kyvaiV93W7pLL00MtKe8f9UDnoMsPDoOme5auvvrNQ8j2DtyAx6PV1+VabJgmrnL
AhWSSi/x7YrrXr32GQrmVihJFx6V15h2NxxgiViAoiieeR/+EdH6WO78lcyDSoKS
EdRcU0/EU8RWs5T9lCwDVCHXqua5lWjW8cuU1k2QZn0eeImB0vkYRxWHeTAWOXWy
kUO4BuIJOy2S9v2EhpyNN2rbCGpcrWTAW7mDDKWxR/g7JxLaqEQsD0M7N0HnQv3p
5uVSAB/A+8zsoHlRSpd/GZKuk5nTaTjs9viu+rWSaesMtBnf8exeTlnaBMp4QyHt
smTVr2j0sz+z/O+1Akg2MQ0/9YwKyzTQeFuI2uy0l+BE44PFwggY0hTajCmybgfu
zOZpx7Q+fLsU6dNf2rDEJKPaKsxFx6XFL3qDJrRotjjWkFALYh7d/nI2f80RqGv6
CW1ipY2xZQB9W7gXObVVTXFh5UqMxqh/Bec0gY/ctrjv315Stk5dpmpiLw08MxF8
z6lIfsVSwkb/NVuyqPhUttOR6lw/95GYErPhBcQ+jZYUS4zLPerwxr9D0pJzF/ZM
DLkOgXFKlpSGkenaQcd07EB+7AIdOdUmKoElHecJpDri+nubDvb3Y5QLYnt4BRpt
41Nz9ULQ/QC/Nq5dO66QZnkZDzTLuJxy0vDJ3py2+nZbDK+enuz7FAbvPPzlUkiB
n3c0YJsJ2HdehoLMlfcl60waGJsev/rCceGjy7aRAsEmBwS/fdRuoTQytbNRCVEn
APB5CdkBf0Ov2Oy1G4LogR9CsxONmZP0YnR6aU9nXx/oO1FXphJIXpYUZrjM5vE4
QTMBeBafyDZnwUKZ2aIHG+Ia4egULy6zxGA8rKEdnckrhtUySCdDW5wcgMSjHhBc
2LV37x/Njb/zwJewqvl+Lw5IINSpbPMNBJNMayZCPIjsRLg0i76NrJquUZn8iEFJ
afCla4MvAKa+TujN1gSbhNDnvan72D8f2qKobB+wKkr8ZQudI+yvCVjnmg2SVrQc
UDQ6BMzY+nQCzOgDq4795s26TfC0i+LNzwfnBXLxNq/VaRcw52BfeQQxVmuuQt9F
C2G8J5GM9dQWnYY0SOId0dQd2j5uKHthE7jTewUbQsjmVB9HBanI6BHXT/Rwk/qs
Dc2n1FxAZcxy+NaPFDDRU6c1zhCxGuzn0x1v5jK59VJnvXqP/14eJguz6pNuX7hx
Q8iOiPiHl9qZSjEssUofNv1cHnvAkBvOM1Q47KIramqg8MrsiBIldAHdAYnlTcjV
cCb7XcJ6SVtV0XWTTFb5qyu6+rMC0cXQKc/smCZJ0z0jbFINK7LPhTfNAU6o25TB
bMld7vYlI7GLIReAbIOJvYsHrkQa2tE+vvB59E0D5knNAVTaDQAT3MWPpoo7BCR7
PpSMsN+ov5gqQTnzO1UrjibRh1gBYSPv3tZWgndhtUl6dSTYgWs6Ng1treS23B1T
Yb+2mPyR44iru8bmEGh/JOo6odAgK44tkHO4NJL23Fs3veFJ0UJlL1nUey41vPNu
XYjaCQq8B2jxOmdR1VPy7Tl0gsgShQnIAW1pCnIm7deYDZg2kykt1JMTbMruzE/+
S6Jq0ee9UkNvBrtflCgKTOxqBZdDZRK2H9Hv48YPWWjId/IAkg4HPOOyXZr0UsV8
ZvDjpjZaxIEzS4VxWcbgOpBv2/mzTXRflRrw5A285jC9D/l8MqxgRwhZDdu/vkD0
Tpik4kuYBFPuU8StcvugLsZH1zwItLD3eAur+Do2iROuBUAxeiNS90JNzMY8+oWU
Gb3iYoskPXQoc6W+ABlo98AVQWNsOGK3w1hBaARWP0K3jTjud0qXc+q+tfaj5q+x
UtrLB+qANplVKLyEel/hsshZjfN9UVt8ecYx7sEYNjg1VeZpgHrTl6IjRUBgpjzQ
Dptq/FWwdEClKO5p1sK3KdCr1bASxp9YFZ5RStRCP+8/V22MW6OfMjP4P6BjN+Vg
A1nS/N+JBQeNudikUrQjmMBn9YlDzKFs4AgNttphDYsv5hN39qyqp7CBHhhGmzq5
ZD6xcXUpvLEKq1IUFSHrhsS5aMGYFsWE47ct/r1a9l4zcjSDp+Y3F8nv60DhXoyF
aV8d2+Ao2znMgMjb6AgCM5EGJPzyctXs9jbqWChg5IA3yOfSMLdV7+PmCHAmzUdM
vQNjhnKLFIPOWC7OWO+Mnmpa/7SYOjn/zD9rVpoDiaSwYq1jLWmyqsxyHRDCyXG8
E4ynSbwFcnn1yB2wQCdihCYyCqfbFfraxQBeVRXtpClb3my5LPZTk/BhBMA1neGm
gjMyWIYZeqSDAdziElPVFDl8kMvwqlgQEhHUPTrErA1Xi0I+HU1oWSxDJuqtkNef
bRL9yhSzf0SrkbpBtGY4NMjZ48cdJN9Fjg9tWbhJgTt8yp831UlXOV+L5AqwQjz4
06uSvBzJ0pYyRskVFRhnjtm8/UO5x2Dw5g5JtOmzEGzS/j8jva3Hi1PvYAFLe1jz
tAFWr4c+qva/6T4MonSHzrWok3OBGetV9D4P/2DK6dRoALNuQPOlud9EXsh39L2C
XKvYAJZTi9/neJzM+cDBChzB20aT+S8nxUVruxf2ZKIa6voLRJR1jY7lO6wBkFzs
SR5RODvRQo+8iq2rYcnN3F1yFw/2Ye/1S5Kpullz7ElGC5n78nnjH4NFxzP0XS2w
v3jFyqdGITchlkrE60BLd7Ww2kEeJ9bjwTJ6qH1q1oMX84Hx/zdMwPflSNn6o5ae
xIwTshTl98XPgfIqhoJq+GfEZeops0tN/RBqP8oC8bc6Xw8mWRqRipwZVT6vl/Ma
rWs0uNhcP0GGJSmVwiIJTSs/XtnY7dTBmHhjAgnaKqT6C5LonqOIevrF/W/tE6Hf
XMhrYlqTRxG5egluQFNZHBQ1vtpidpFrXhU74W32MM3LH/F6uwngDNXRilyHvkrW
9ts6N/kkGGLOptqj1iWEuks0JyX7st++v1kC1zqYz/g5CheX+9eBU30URVt2WUim
9LETtTYRcIZdAaG6F1ry4aKcu+aD+3kDK4/52BZPJtKqiBc2TMrQ+ljIeIokqBDq
hGJF2++5taDv9FKq21EXiu56KOPMO4ijkPYcGLnU+yBAG+/VMB+r6BKLVhhCqtk0
t9OAyFB7u36+8qb/c9IPltdpJKMeIPUqEb4/lH2qizsmHhUrPMjRKUfz3AUALfcL
P+LI+1nC+NsDH7CzzB9H6cSvbHWjfKDKHpgMA06hTEBJ6kwCvjS0/U4ifgP+n4KZ
IJRr7YCVd8AaXAxvCqJDJdITPREdSBuo/xTo+fjRaaaQV917NTae1Fou60KDZwuM
p4eJ5REb7jP89rY9KO4tjH0aybvad9uhyTQAEgcSZ3mM2ivksX6YlQAMqtCg29Ym
lV/OYlXgWeJ2gc5GZT9SCtvFohkizHd9uTXe3PFlfZle66izoDgqhbDEkrVAfkjB
jRSkdSu/JgnyjXzc0oFLhJDV7WQcofvmhs1SlNGL/G2ViJTMD0Ppgp2/+PcAAx5A
dI6N5DeMN9TDoZuNvTQzkH8QmZ1SZ94Bm/MgrIrGyjhDMDgCIdYxrhdZJ115oPpW
WmmCpYzhIKA2WbEVeS336RNAGDTdKlJ9/jJjBw4kn9OlhP9KVNP6aoPbsX0eXcQ8
N3CK7yIqZAdtyLW2txM/3m3fph0JVL8+9R41paM3w4EXCblUHlV3f4RMVIY2nLOI
tsZfL0HJWqRdW9JWfsK82XowcsaH5GxuJy9DGq9a4beuskdv7TKxYGecUCILDPeh
1Mo8aPb9X1dGFCj3PFpgYsG6NN6nIAzPIIY9pMCGWVYxMtW1VVK3AMTUmgamga2u
XvgwjH4e+U8FMlGSRxRH4RjE7zA2UVs956077X1+DPBizzKqxaeYpMMmET5FbEo7
qH2+ThUcybJyy2M56B59OS/cf7ynne36vGPud46mPioEC+gE+mGzbp7igVep3WqQ
OFzrbkaFVlIJdYWrVZqyhjrOhwEQs14omPPECBcm6FYCAQ8jEkTyfvozN+kpva3A
QHn+dGBEf3z7lotS2NgWYTRZ89ozg9BzVNPzb2iU/6Dvdy11c2S9mfXtcFYjYXnT
NpuwmGe9OV/BjfvnuTvLBtGXWjFWktRYdpCuIe8HAB4H6aadfILViN9E20Euvk/1
HG5IvGAyD8AWWJNS99NxdZVKtevkAS7MaJprsYFzjZLm3VIRFyGAWOSo8jWr0jku
vVEaCYv+Myx7Tpunu563xwSd4KlT8QvnJxbgK21Kw/Z+2npZFGJrthvX9SU2LE+S
p2lpkJPz6UvtAs+B1oDWOGCsk0tHQRBjNyTZ/vNZety/K5VUNwKd1AEkHb76QdBT
2JTeDTcFErVA1XC6AoEFLqzgwBQsC9uM95ARjhpIp/ZWbLYzwr4QEnGL4xcA2iX+
CKYvea98UYO5Ud+iCIi4BEP4WYMEMZSOTuoxb7Ldci8L4mVaY+3jQ3qP/gKjrx3e
5BcJequpUJ5ltfTxDBQbEZB8GVEQkrHk8kRGXf9V3tB25L1yTR8AhWLscmHnMLcJ
7I4715x0LCw58/KjugaRuFYRFnmicfFX/G3Yom9mKpeyjAWAL50IROtr5amxHGcm
Aosnzfwn7MCHZy+45uhgMVp94UHo31ys1xXarz2XDGnbRvNAR/0od1OH2huHzIdl
zlpJL/qtyhyUn0+X5jNaZOztfKUo/hlCwq/5CQBO1CFa0bXBOOaNRM8mmiZdpdaa
EeLOWxzPo7rOvVn0KfxTQxmcaGKslqL1VaOtluahqj86Csv68Fo0nb6UNnMRJhJf
jix6/warHB2IA94YOeJKviOJIOSIsErIzAYhrsgQM6mWK91gW7ZFzjt4sXgplyRe
XN6P5jOqLKDr2mhDBZeM9RY4vN7XK3Ejrb3/Lpn4AAjt4lKNESmjO/HTwuP8/Lkx
r88YLp9k36UEO9HoHDF6Ne53GalnEYpmw0ZP4AME9KkzzxhcWpBknOM3lm58EUML
fS4Z9OQk7QKvsqLxN9hv04Gj5acfQd5UAUtd0HjeJEBNCMjVNimIMJfKFpcoVaGk
0WeLDX4V9HV3Gmxqvirx4CnDUGGYkRK+jPih6WBfYp0awG2eiMQxYUyrp8i4RkuO
A0OWOc5iFc2iMCdcEUI355WQjtd4zVC+J8yW2BtUq/YNLnPHIYzIhlH4MyIFbcgd
3bhY4MerhzMazIQFWQOKt7wwpbboF7asWZCJ0HDREYqQjQ6063NmjkCxdAzQLHgX
UfaHSpFmQNTTHDrUAzhxB+YQmdua4NL9K6TMfrehTIDeJLw54zaKgJzHFln4wqVR
oMD06s8rX7FGDeU5nfM9HUuFaiRXAMTOpEYSTP4gAEmENDsPt8ueX9zqsqCipx8T
IUPm7euHLJ5UO60+cbXTwdrJHc3cLBSehuNvI8vTyZ66TmGVPCDCa+XtNqL9NrPu
bf045GZv65yHTjkOd+J2EnwgdOpxEY6TU6NS+H3ACRVgdHYsjwty2qLMnJlR0VZH
nXWB2iW4C3loRwjqZ0ufT1A7i6/yf2rQeYLdrtNW1HSXtFayYqxK2Vt4JqYppApS
vds7iDmaNmsKdYvLWy3RCBnCGTvcG2dj6DyJwpuD4lEEzja7sMWNcdmQykdM2RN6
/M8lmIuibvXNqqPZHQeYxFx7b5kIAVXOxmJG4TLrrTRkO9M5hdayvEKbp9IIfZcY
e0CvYb0ADssuUBqRk2hTBKrpGfnPiHKG3OeTQfBqIu7safipnq2pMYRHTJ4WWJcw
UT13xz+VIWrAKCEJt1LxAAjhFagQHTijo5DwEYtMaGmYV8SAOXXsBmKlRmotqp01
Z90EpV+/xKj8GcQLbTY6eLDmN3s3wzii6+ErS8ICKb97yDpF9dF55sMtj49O+OJ2
6ts0zO0+SBnqjgPhO9ekrZ39WXNFO4Lnsa0GgQGw5UH9xvGK3Jf/V9nSzAizOtLK
acTXi+u27NMHSb4n4pv7y7QgLo83IK1+sCC+7ie/jQbVuVjJ6rezPkOXE7Xwdvu6
DNWMceJFjnrSZRPNe+bJ5C1UV0sXHdTHcUK8RQRlBeGYq+W7FXicVW4OoD1oqohg
FvC7dF+m80MWGowRpevszn2GgiP/Wy522dKFyZTSgtFPCmn0gOsMOuUoNmD+W8TR
XiUHfIT3QoVN7VcAyRNaMJ5J7ras1yuo8CnjlZd64kRj3edITQJ/mOIWdHHBgEhd
J3rgn+Yz377eJiuhbe+BxNh9nKEsB+MGQxNMegM4fLX7dGriFexrSVmarlE8Tkrl
c6SsnTqRHSSCYHPWeVGaGcB90xbYNK4gOOyJ9aQ/kMWmjau4Om1e/x9D2WZhG3bv
oY7Z60DTxAJO4wFjn54whWbsu60MtuodtzuQni3hBWeUT6QBq5nVUGVOzCn8ObD7
HU4SWSMxGNcmFy5XZuXfOuoO+J7mJ6x3uBWX5sbM58HR2Aio6QXo3T4hlbevgjs7
lPsu8M7kNgszPsDJKI/+YdUcP9vPOCozccdj2hAyUFglTrGiW6dy1drrGo/PQLdo
UgMt/VsTqKDpAZPUzBh07KN9fFY3TkM5udSX4hWSy4pDDTi0tzauRtgxMiWqE43f
MG3SdSGcjaagL3pfymBzwWgjafaqzzMLIpmhYSH19UUNk0KmrSFKf7GMCtMQzJ2k
7+MSMG5fHY4eXr3QapqJCQXNdZpeIQJ574QQkM4VXtIv+9WbB1GAshtE2/OaFjjR
4Yx26ZM/Yw8krbX8bRizcuOWcrNCKHWbyye/BiY6AmNEtWR1Kn/E0fORkIjUW203
KCGQ+RSU0YwYmqQGF2PDRysgGiAXo+M0TEmhkUhkZjuz6JEb2oTeICFl4dx2SUWh
jGb6JAJS+TFfygRGYIZ1lgjkAIElsUHlbQ7SSvOW5XIObJL2kiH8qYlCNcNvmy7F
rkEt+0vnM7G5uznCbFXj3qNBNcNaossKXbUll/aJ/aHo1wGpnhgpZBFdvyn+eTI0
RzARamolxNBSqF0a5LVsn4qQaLRDIgKJCfjZVSONTpSPiSYamlKLecXl7Bgeq3Qs
JahhE4RHzUQf+OUiWeFsjQmrD7j7P8TxwdpbxJOerqKbQid0XwZRx8H2bHx593oP
QHExBesCioFgHf0/wr0+08EQa3ALFcqg+/USLY4diqOChJSqaoGxpO4LsP5u9RDh
2+dAn1K1n71BPw6feBgC7DJZ6jtrYK5vqF8bNTdioJw6ufcKKg1RqAOaZMniv4xp
kGYbuVlbyJDkzvOd64uYh2WoWzl7v9AVLxAVwSxLjFnQzYbqPor0Nmi4KpXmbz8q
gUrheQf/xlOparnMZZY2eAMeX/+OSyS7jIcV4ArH8TURV9YUJlu1m8cjIhYdoiMO
YxF0xN3xrWxRA/2qf3YTDpwj5EwJzGYFzFJ3auER8vojAQZxFeFEAWTopoWM4rBG
47fVd3mih3ZSqf9c3TAMHhg2wpHcEUqzvlQdXVnDXYERx/91DfTAR/Cag7cE6TEb
/i0J1MZPCnaUFxSqbgA/xTudHo3WRu+kopEGG/83o9NQpBlBd5CDQjVUqznKwY7j
T9Bl/K2UphSo7I47Iy+q039DsOB8CxUgxU9pZwKX8ZbSPB8U/7xMovCK396qGyXd
93EEIC2UuepkmV48kX5Mndx66390S3w761uNGsA47xeSFbe/w5gpFY6FTV2FuO6/
lzB2DfQYpdYc1U8LkR4hYhPXzTk8v1CkbqwJw8BqRWfk+zQn2BMlD5K0Im2HlYyH
0W25d+bPnrcWPnTIrifHyiNnJsxtOD/CikRgUzty80P4XgfSUifnP0xlVp7OYqz0
peBedMoKBLW+6JrWQxcd7N9ypCwsb2PJ++dj4QCow4U41jJyTynaTmiertixCueC
eCUhnh92brPWQOjDdqGnaRdU3EMxZWcL1kpVD4RHlUR/36eH870E7EjGbc8c5yTG
wUhHlA8Piz/cW2riBdd63J4iMQgk0O/wtLROm8Ep7cKXY1Y/b6+ILAkqRfi5xkji
bUYb9tZRTgym9O5m9X/gUlx61fHEZt3BrAHL4/bCd71on+akwMET+gAFOPurMC90
tYWEo/Rw8uPDQUaPVeI321my1BYJV0IVKa8YnoyjgA3kq+f+ulQLq/FE3/gVki9k
L/5VVjkGojVQPh4MIGElFhOYgcRiGIfh1LSKMNYzBayetlQ0EfuSLEIIv2FGt5AH
Ld+YFCxYXSQmFcXGjX6bN6qaoY6XfBU6wPG2U6cs/A8RdGcL5D7hYLiVozewFdXY
mUhOTpLOtjmpJLhNpmfdcLSdlqmiVMp1zQjyctR2ps27IvQ7TG83UAmR7l7x21q8
hpm9c5XVucGsXo97TZfa1JBETvEWzCKg5e4VTg5aS66ShXFNbZ4fMNTlfcvozd5l
SxNqN345GPeVBTSOP4NuxqAcO2MXXWxsdUhwvoBt+IC7DJbST6cQOorpevTdzzH+
zLiXdP46J70Y5BlD/ejEPUoKRYpJjeBYWvQBZ/7bxrOjRKBOEOYaV3hu9fsOO3Yy
atxxb1NZQo2WXAgYkwI2fc+7LcfmBnZ8mk6YyeE5ibKmqyuD3My4Gjg8KTwiP7q1
5SSDrMKLdVWScpOXg8bLy6sB+kbnyLAIPxN1EqvfF+0XRtyhDpHuum5DGpRe2dcf
rKHvbR1Bj1VtxhlztPXMIbgNIDkovfJTcCnD65a3j+DP6VM0C/whiAMSFZP45HgR
33JJm2X01PT4JuJaXUYL83ymDQaYo2WpkwZw/dLmqISx4DGdLPKIdGuS4FxjllS+
zwFQ/xK0LH+lQf2et6ff4i8ifVIGv8RKT/z0CP1ATAiNPnz1p3kWObsbeNdd2kJV
EAebW6WEedpR0rc1T67Xoyo16JNk28v7vsTWPttEFyS2eXoSD54LkrbgVgrHyxW1
qcOwkMDsXDE6ZCw59me7QwdNphz4HZIuUNkqNXBReTgYyfqgXHfX4FlQxWoDvRrj
/VsVsYvtgfexseuWyWbkaVytPT+qgr86MTkk2Fd3LpUqBko9Jl8vdtL3wHPtrghe
X6rqTjPJ1KsfHggH3UV132rJvBE1DtEGw4JJNn2H/nRrCkp6Dvm24do+kVVQjtx/
2Bx4+P4HbbFP9Y88zoQY79fc4u8uPtTHRC9bEiVhWn3B73pUH7Ndg9kIXqlGWCaz
FvNTHBAA80ZkeAhTddeIKwOBBg7kpniiJW5gRkokOMQjsh0VizlNWk6SdhLocOQY
VmFgexI1FxnEPDp5wjNpXgfeQ/hy0kt64v5RxfhF8qsHzAdbbVvehos/EbtPcAbM
7WjMryzuEVsCO0pGbtaq7D5ILse185CyAiZCmtYMq5aeEVhDUAMkfoXvE7gwk0mN
k45iSkZTLMP7fLUndkHdhtHP2YMBD5z7tHBFD7Btr40+RK5ne0ex4KQ9h1Boqu1j
a6ECjUAvTM6L1T/gusD5AmZ+7J61Y9OoC5bfXcjN/QV8L5A4XI8bu8y+R2kwz0tc
F0IppAK+sAhN+MBZ9/OgbowFYpLYJGEIk3h9buidFTl0Db7jLSrzwpj8sSyEI2Vm
oF2Z8C9RY7SxrC1avqqOBT5fWcwnVjCnVWIgfILyhGLyGUBKgqieYRauOWLOAknq
jiX0jcGt5IJ/TjzeJsChgicVpkbhsLFvTuqzWVjdM9Icb8Nmn0v6kXFm7U2QCXNd
GTye1P0zsvOwL9OnhigJLKt/NKZf9OBjHqXuFW8GZz7ZQsgcu9RWX1UTU4MyQIuZ
TQzusmUp4JgvXOXpYHCKtuGoxXzJid77U9wPbjhnWDnJwhJGOYUxK7oiIVgp8tvS
lyz9PaN5H8Copw62NQME67pxb7yiR7rRjEPZEjAxMV4sScfQfxJpoEDV+hQWw3Nj
1BnZspJtBphhuvotPeIB3BXI6adYooijhaXB0rSmXYmPchEdrwMpgjXviuHUGsNH
gLyxmOL9TaNAk7RTQrrsjdFiFho56Ymv5ZnY6H8VBfyP83OFBbEkypUmYPqgY0bs
BGp6svk64CtV9dQzwxKryH8ATMb0Am3IVPs+X4kgbfL4VsE8mDCWVD0S4EQ+vqst
nJvbHFwNkxMv1UMsRT1B5YvbTAt5W+s4znBsJz4CBS+JFz3Axbncx4ly9VVZxrRU
ofplK8CwZ9h/S7dP/fyrEmb4EZR5WRHL9vvxB9DjZ3rAR3TMtW+f1HFJwvg3mbvA
pMPgBHh92RGP4Ftynqq1AgKcXfmzHN65JArc/zCdZ17aJ2SNRdewy9YXbhCCf0Yz
uXDzRVLyw7Tdf9wpngghlhLPX+uitCpDRkWKEU0d3Zxx2hu4sxooTzvfjR8cnOEE
OwZgP8GOJ3FqDf/bt5294VD6p68zoQnEiqgjfDeD2uT9Lo8rdHRTU+D3rZ+uGBnn
ErJMfylmQEFayrDh+tR83V79cDRHYOQW3MMJ0wIV5VY74XRDoX0n4wuwpvThh0PS
jTEwV+a4IPCoxBwEyA6mkTQP4dbFPbl0Mi08AsWZuhzLxVAtM1pU5eD+sEUcOgtT
T/53rO5LtoAmk0zr1EcRTMdUj3NzDBm4ZYxDMTocUWglP6mAnJmkjFzUEHCpqqDs
CoJr2op5Jt+RehsPNya2aSmVUSfvdYxwuS6cVVhQS5E9eUYWHapYOmoPbeUN2zGN
uUbmS1/aSxTCF/vIZLd3nFp9I+MH26PKWwECrgYTIleYlufoaSrOXaBGRGuTwwad
l4Zrk2twU5lPlmq5B53sNZiPRGJLcaSvlwbPxreVZWYKTtDaey7GLhIH+5s5qbXV
4KTzfutDXaE525JkkW3CYfRdbeD2AR3EAmS5MQY9VYVjZMMsQECzKGxdhCcnEEBi
3oBRgPnKJr30TOSsHzC/eb9HF5V8dTyndpj+FI1D5wyUEmrr4UgtDzPJQj0bv161
FN4QzAE5uTM+zTrUdelN1kjLSVvxSwoe4SyMwQEcHRwN1dxkasA8U/0S/6YFmAV6
8d88SeDag3h32EohLdRTfiLLbOxZOh0DsniLcIjnCzD/vxTbQvxap7gEpvidslW9
B8/9oC/H5K86yx9Bn2COZVz1F22Cwabf7r8V6M2/hPvIx2JqZrBIEWTqwUwtsTjM
fFe8Fgjq9uFlWOF5Rx8d981nx7jkwoD4yRLBxhwZpI9qOP3Be/6hMXdHX54BTc79
+TGAmcUh7trJUSwUmMGCe5X4ImaVZazkJwGkt3/OYdyAMLQ22L3AFG5DiJPEz/Mx
6Sl+qUeS6ZdauoElo9CQOM4C9DGk0zbxPZlkX/98cn3RKAMlYpSSH5rUlKL8rqGE
20Pnu05/PvrcLNZ+sJ579iU8AfY8ckTvefOUv/LJbIxwAY1BZwWmOUKLWClFjPJe
MrEk6FdcbPYYIZISEsUu/Y8kJn7WcRBzQ0tA1ZRiU63ypPjUUKmPxwuhLhQTymEo
dgA3euZSoOwXQI23+2z/JHV+kw+g1zXfItnZizCCjnMrvgM1PPGaCMb+H3XkQDaL
QK0pLS1xW8R87Af9xw3VJImBwq94SfI2ZN+45IujpJQ+a8/2vSvIKf/OwQQai7XY
AYJtpbDoVk6QB1ulh5Rh4e3HNEUGQSd+t8qQyhLoUYtgKc7X5CTBq4WM9/T6EDij
08SGMFpHQelo4dbo5GqmaJLSkki9K6VeLtxWKj308KlU2rAS+Mo1JqM5a8O52lre
/ZUZedOa1N6+Um0tDB1fwZI9SRdd5Ss7Ok7Pn9QYSA4TdsXb/sc5QAqma7tJZrmH
WNqNOeI/nwbV1rhanbBiRexyjwkQSL6Bwu7R41TeG+/BbdzqSmyL1pTZ85mFdVhY
Y7btdy2iLZrnqcpR8i3GgcvrJJW9jo2tNU4SgxXs+XReRGQF/hlEmvZhPtP0erJK
7lsxz1lZfKXKnem18x24ZpFBcIcuMUNJ3x3h0F4ljr5hlMcTZnDkgPaXG/wEEGdy
8+E3nwQJw5B/ln9O723qxzp7JEd79fFOPX6M4nhOV/xHLUFeYUMKCK2Vjxb4YHLC
WBRtm2nqB0daVl1ISO+5YNw35HoUYYTA7j6JUMUTlwY1IKUBjGMLdraLLRvWqDBi
y3DHNVQICL1jCwtbS6LxTSQlSTOiIN4DpDGBCRcWt8NDVsJ43ac8yIiCNY9AoOFU
9ZA13h+rQAL3iR3QeYZN49phTy5rhbQlWyx4LchXMZFTHEz8GOBGcezpn/XAS46J
E6FQki1DKCXZypk7ICvwMpSZB+3isX6sVTUriLYI9FIXMt/rF15J/Wc9UUWp0rtO
GxlG2GKCHOfLKLQBpRTvyp4ePlx87jO2QKT3mMSKmtftjr7aeJ+CT6FFzyfBb3CQ
aZbyg2ySbnSXrTWFHrbKLchCr73k7qej0qvvtuR0lK5CXrELYMeD6mBFSEFkUwEV
yC7tzElif36ckoP0dvTnPgRfSktniltpy30wKbYmm8SxqXfP3WSmN8GcI8mgdbEe
SZh8jbFrxbyrrR0cN20GKP3z7D75qvlgKbSuaQG4EZA/5JNTYSWA0N8HUuEPVqb2
BwzWuL5UVgdGcbXaGFwDReJK5bbIph1J4EiCmGK0xBikfstiKcF+HNL619HYiKOA
h83aYmX3+jI5cu4h5p4ao/bU+DOOBxpwyL+oqNXJtD83pDCFJnIhtemaLZOEcI9S
o07RQAN60xvpvlDcqAn/KBxIcN2wLCazgse30SKpa7dxDK3/IU+nFRBuy4GpvMep
jzDv+/fnq8mwD3nex4po68AOecTu2RywGEulx3V5xx+D710HCnnR076rfB615bHy
B0KYbhZSkSPLI3yvGx44YrOfM5oRToj3bQXgVHaBqZBLF2A2gMsG7yAs54btqUnl
ntJB612FmrKVSDtwzgSYkKGmOYudyq7W+0M5dCcPZ2kfVCa+N+48yKsQqPqaYAK8
FGVyRCBjooUnUU08CiJS+pzKl6n2QE36eSE8cG/hMEVOZ2wrM9i+Ur7wMEUWAkNV
IhDB+otoef7jwCdAPDgD6slqHzp5NpWRrGz/Sc4uHE7eIx4qdIeNxYd5btFsQ0EG
4DhkxXvWrjHsIIOm40M76qmimt1Mr5Femv1dJJgFO+Jynf3Vuu9ZkAvsvW5t+MhT
O+xec0odIMrORmWjT8VBIgYHOnQOPCOHDw8DSsTYuJGLsKOs2WgUJkfcjlGlaxHo
6J6cexcYn+EekM7xhi4zo5es33ME2E7IeiGlKo9IONIwVW0XTAZhvqxdJmNArlLK
1WNa9LtJd4IwIl4Fvnje/kkkyswU5BoeEZV8ncymNUzSVIGQEsriQWnrDYK9BxxR
4/vs2Z7cSstknOc4hAUf3R4NXV+OYKqXWHgrFONlnPpNi5VrO9sg0/gIzjYdUkf7
zBYQvZdx0LOyAyZwTDfYioUtc2PLgl/opcz4fXMB+Btngo+PNBAoMwnJosDS/2Vq
EGgOD+treCvP+G8R66Wp8hYoDMnS93Aht8s1wJ9O5AVmuRGbMqOVTiQH4pwxeHJ5
2ZROX4ieIkschRaHnp33HhJxyq4r9Bc47gjUgFFnRpNDNmuk2ql5VRlFl1yIgWFi
EzK2BmqCGaSJJ22WLBxrnmnML61N9yNPsGiqhnv222DSJPI7vvyN0KkaKtvKOyN2
vuYoiAgnq42vWdLJSlteDqWx9TQK3qrvQ9q18ZmiWgZtroreKmKWGZftpSAYc31F
OSu44PGBqHhLNWAQU3aGUPwN2yllVrxRDyhvFubJ84mvThfJoWzyA5xROnxqDOVZ
REAAuWyGylh8SeSbM9BMZWDobzvoywBELjZL4XSpCUw4b7sTBkhKoy9RCFJGJbnW
xLiovJ3Q/fKt/ohr1NXy5oRGLwHJR1BcyPSCaNGZt2eW63qjHB902mB5/ap2kIJg
b4XyQFrpgT7BvOHpA8b+2qrsqo/ODc3ZuWR0VynuGrbsZwDiTpv5LjOdZqwfAMlE
35JuOQmU5fqleXN9XZ8QpZyUhEXxdY4BRTWXjYPc6+i/FnFCPFYiuDv4+Qijrkru
KKmlv4O85s/IH5AtWmANakyZWMYoeB7vFvH5zWmh5SKVrkEIAJ47RQO5SuxXvpcq
Z8rqWmdxRBFyX5z6tl3v4KCh/DzbyDJnEtjQwu+ir0SzsEKyYWX8ROKroU/FThvz
gee+ieQcwi2jRdMluZJjPEFyK+pzYrTQjEI8QIImElpyn1JsfDzXbHhzHZQNT7oi
FV/Uw8nBjlEUGgty7ir6lTC2wyBO86Fjpds/afjF3WOXb0yfesktqDJyka2EWMKn
ZUrnUOwsRzER2MFJiG69nCRlm+y+xt4CbKDq1ep1Oem/XOhHL6Ft8VeK9koJFi0c
Bv9Pxs2lM05sT49EttRn5MMUvJ4yPUqy4cWw7ufIh0jcUauJicIvtSDPRL1mYtXv
9I2QNP4o+JKAQEQwZmixpOmY7xYiUrx8A4Hw1lSUzSKW4mDkiCEm5Qo0RCX4wzFI
BTe05NrFoX+7eo6vBSGoTfFGKJHHA1XTiTilbpEhUpVtLWjqhomb2WQ6+3JESjzh
NvBnOtABpenmTzDFK2GG1/GOqI/t1PNjL+HQcBvUePBBHcXI1uthGvCDmxkU8mpg
0IWuQO8xjYAfbu6w1PmFnTrqxv78h+8FrCCnSiWQzwi5tc1C61dKUM3/SknkzaRX
ptF/p7XMzRx2/GgGC2a8gm7AhlBgN7MSaaTonqdTjHJ7V0dYNNf2alsnai0nf9Op
sihMsGN2v1qlWcH47WsRfDW44mqBrnOONYKOuSE3EMfzRf8oS9pS28/xmi0DWi5X
ph9oqvPl8yjk3HqozJdg4T1POpfgVM4oQNeE7jdbPZJN/3j4La9u56rj7EdNI5K2
VpIbCSoU1hfuoHsPib7h1IBiCSXQ6R9yw757CEWPvzlHVl6rnXp6+AJwr5Kd5If2
+YsaGMH85N6mXmNjnOe4QaWUGW7cx1MyFyKW02XfUNUw8B3i6mv465p0/OSejCrO
6mZ4EKC6FrZc5WeNTuZbVEEt4+F8jLvNihHTTD/xIViGFos//xWIXFSAkoG1yA5s
uOqdV7IastmBMbwEEfR03NYxDcQdh/dmL80KXvWwiLYH7iP6urwDbUsloYLgJrUX
RDfpS49i0zdJjRQSZXe7uWFyJKBfjSH3rMj5RmBrOKEeAwIVpTGar515j5tLqkCb
fBxY2yftRdb/Xfa5WY6Yprn2fbGRicNIVttYYV8WFZlGB+vAnkvZ3hAuKBsUmy1i
qaoAR0zVkLcmqBD2L2GhthVIKi58nUmLrJCzKxOrIDYHkRX8SX+je539OMggeC4u
R38RgB+vZtNIBKPNAaWZPGy3DcGFM+nYhbmlRmQSLp+M9DnGTnN6HIqelD8Runo3
0qVdqv4mDKZyTGCf51GIOJmiXNa9TFXIGfhAJk64HK3uEglQsEalW3oq2h+jCfGN
3QlvczaT1kWK80zCkSShFL/BspyEOLWb3d6l9Mpp6+ANZ6nxleNM63LYzBnWmfVY
jJCQ+LqlJg3TRTG6d1oBUQ8K/sCA9M2KbxkDDcxrQNMIRxxwjJQ5akP24nrAvdIP
bqHOOm1uPwnAQ6qcWaJGsOUANLXNxzhrtD5EA0mFxCu2QQSoGj7FaJ7fOEEZoPcM
N0hdgV1JGRAGlx2IwFrLDyukl8IMvQ+WY7LGn3sPPS5pWbZ096VkCUBWPan8uMnt
oOwe5JFxyH/ckdXuj5UQ1RTdmjdlw7EMJl3homqt6C4Rlk/wLR9Fz6RXpU6h0sTB
dVfbEmJ2snfhsE1gdRYi505LghznwSxiH22DQs0toSwaiOSziDEEHh2Q3J+FyF4k
dfW8BWa4zg3sClc7Dill2HqNQVpnCNdkQHGeGqwyt6VEAMQW/IfUI1BkECvlQvBg
O4B5CuRUug2wJLXhEtpBF4micmXwJEa5Fze9MU6wWSvEkNhvQ8piRWRPB99fGLzv
D5HydQlggHt5JPsia8ctPLBHzhcOvNF7po3z/LHrlaIW1j+ZriKkCpBtdWakpxr2
3lI5r7LjVdigiwPIIDAStITr5xcMfpNJe7I7R73IRHzJeS1NBpXGO9DI1vzrfJH0
PQ7dm5sGtmiQqbKj0l8uDhWv04Zwz8l0RZqQFv2hqcHLGpWNQ29RNGOnlVSIMhs1
INmmm2ogziiBQrdkKVrzNm8tGxAqMUAsZ7ou7asDg9s2k3OGFrGF3it7hVEuSr7a
+nHbhV3m36Gx+zSo8Up/lgiYXLuPUxZYofmNKUD3zg6bwdRDV4OHE6tJgtbP+57k
D36iwTnLrpp7zvcDyMwqiJkacX2FcVb0ifobVeEo30nNRZBi0ipHy1cShxVwenqP
G1oqE0jaSeNo5arCOAsLAjEnacCZwLaujaQqDs0ZrYRua2FS4mU5QoJNbXUA2qJN
nDww493zFuNKgr4A+kBi2xIUACJBnjoKvKotirMtj4/XxPeoFrBQRyKXTtVZB5YB
t+fUdKVDWaZV+62OBtPca68qu/Zg8wpop9pZBbsSnfNRLOTCJ3d7Ub7oEnNSmjJx
oUX+bkG7Uk1SQ+kCj0WSp8BIzV1LzMgjuL51aQNXUALHtElBA5J9Ev9tnrHJYw4+
8yMdwvRxVsq+a2buSuSRZz+ptnBzkEiHGBUDUSApAEd2AkX2fn4EuoUefa6j1PIM
f82RickrniRsPU6NZzMkJ2pQVS3LtAroZvAoU+OtH8y9twsqPoN5ulkKarb/iV9C
ZTPtsqNid7E1kWt9jxf2BoAjyP9J64Sp6OLHq387B2znxrVarpt2NCNPIwnNz5Lq
yEAluwejQpu3wcCnxoLsXOlRrNZ2WnHH2bwnn23QnyWOtKashnCjy7s0xdDLzgTx
gfXemvQ26i785PA64oqYkwYKzGCiJWHIMxeUFiFuVwqFubxHc18Q12QLeE2NLN59
apuVtkA3OfBMcSFrkVm3iB9Z0FgDc3TSiHvK/n9C1SzuV/x4B8rYJxBrTjQR/zNG
dVhoPf5jQUTWoBQ4ESfbhvvUpOBHOVxH65i4tz9qFZVDtSRv5p3pHdh0ETEKLbyt
3BJ+TzG7oXUIy19pp5sev9gouwKn8xGi9WkFxzXY0h6HMK7eE9sS9idw7mZWMZtv
iCx3To5m6Zwv0JyWa7fdhtcQHckVhG3e7vGiphk75OJP/93vBXpgLvuQAeSgUFJE
y+1CO/gnC3ur0awmI00b7lhBepKdWe+yX9/Z2baNNDow2EyJKc7rMutlJscrKCyr
wB/+8pbyfda0NTg7D0t+xLWxJn6u7Qt+bXIAnWiinuucp0XGVq6BkCd3eioYBxXh
ej5Zf5eEmweQ3ivoGMtwMSelYqdu/Q8mijocjp8v79EN5cMnjaUGw5EU1BwrfE/6
YixBXT5cRM3om5lQg+LwTW440LFPV644PRoFLo3Pu3lxp3xjnMM0WDW5hmPyMcKE
cPk9OMfvz8clfVuo2NuvmETiOggJmxTByJTkKuRDoh8z8k+jpp00eYQExDIwxjwI
JnxyGzZa+SpPIQU7qmafqHzeDuc2Yz0eAf7qvkMYpYPQemZLZHqr46GAbVovoERk
4Jr6UPqAhhdBmk72Hpudz1r3Ebxc0hI6OwHSEgON+EKjxgCzWoyJDx2CMD7xbJoc
/ugzAsVUQ53XNtXjWnkIi0VG3HtayrGb7cLefUizWtOzrX2iRAoatIvXB1U9Z4mo
GUl1fFYAHri9Ua8zsGPqn9K1cqGaSYhwUTqYSPE6FezXG8oHFhJDqGaLAF5VRK5X
85UaPvwVvA35ZSFElEeylCEo8o2ruVP2w1s6z+HrkXUnrpOnjnj63vnuthbUugdn
ipP1aQ/fZrQQLnZwAnUgXBzXx9S3v5LaMe7sJGNEpEWvM7Lw96gG+pbgfCQOWFNb
sO7GizavEoLAgwYTPQoCV7kzCdot2da2BdbxWdxq9NEYDRoubYviq+rooOQdqpLY
FkYhc5KY+5qV9nduUfVOu765ZoWMHEC7QqVjpeqwwTiOB2aWJEio6PsWKLjfERzU
N4U5BSUP3/E+0j1lhu4mLpAaoL7vZ/G0tkB2TE7SSpzb+7ax/cNFKAx7PymdOGKo
q8hUHZMW+TS/hl7DMxXOHr8AqXfm2XjFrZbfqacw5SN3lANGFQX/aOGXOmMVqyAJ
n7mtmkHIo28lCa65lWxFcnGhP+r7YP6Zi/9uzNq7wb4QWfzpPxc1MMnCj+b06wSw
mZj7P+uh9uoc+mbxPSHnhQWMj2HCgXlYbtYdbU6rjHo0jZvx/Os6j4CwNEWdhCF/
cxHReKi8AvNA3CNMFmD8vO4XnRbTc4R8JqSLwUSMR8cSz7m05Erj5TZ2iMUe+lVA
x3GTy4bprfSsAylLmgMy3HH9SShCdqBoLnO7srqgoWGfxV11IRCgwCh3xuQaXRxv
js/eNsMBU/DeXOukKITEHx7dxnVspLdIIcUQvAaUtLMMTGE40ig+4IBftsmE9dJB
vJ1r1Z7WPwA2BZ77fmkZiEjZ9eiq52cMkSHOjQOXELf+8oqdhWt76QhGjUgTBMCT
oexX5uqT90B3f8nPpbQNywajktQxtEWhf8ZrwgSN4eIIYSpk/8CP4vcUnqFE/Yxt
r3grzpHxFefYEoc2SYdQsHhBqYWKmlxU2ZXKmbvvRrpmSAoDT17V6RwK2aH/ygCW
tx/hcF2bgfAkLRm9n1nJMWeXfeh2OJ65+j1wxYBlI9EDRWl5frXVUSzcTPcDUSsg
qB4qBCyLQ8RBiDCNKoqjRNd1B2xyikCTa3QnA3q+RAVzVTaq0H5WmKvjYOFHiE+S
Z+pQzymnd1C5CcW45VLpFfW0lBC/SJowbiZd8rdDDVC2FxCWVrbkn/638sXl1q7M
dzwyipAhCAXR8YHUfMf0YLXgqd7tlzYRH2wr/5aM8iGNdhpQj2gOSJzC37I2CZPa
OuM45wcM5thm2kyIhorcySd9DYyO+L+TqmKk7FIeRjRJ1z1VIAbJTKS+mjAPU948
4BvAA6xcOL8s3y438PZ33vU+W3S4ewE8eddXffq2AGrTw1ec1UIswtJdK/eKdLwg
ucm1Fqx0um+W8CvVvVgbjhCB9B8G6L3paw+YeOQVNuNvOp6DpVGDyOdEAKRMpAbO
gjYRco/P7kNG+uUT1s7rtSSZpo2yZSe1LZF0KnM88rwDgmLQSjyp+F73ntapayD0
UibSHi9jcDE658FDtQDn0oAEYy80f+BARTmUhz1wesVaxKPbgDyHvQ7R64PtFahH
WOZ5PFRedkT107QWkLHxdqd/a6wbFYlyEzaYJf1Gj0Zx6F+dSw5XsgPC8gg/d9Wi
ggm0Ofe0G6m4WOVyD9zzDZsqRaat22czgo2CbtZPnFnvsav4dAbJBsq0LHp1etjo
ORakusWiIkX4KlPT7dAPjofJTxs/OQSqDveKYR4Ug0ikFkoE8pFQY7Mzna80ghq3
kXcc+YQ8qIasa976+S8Bla8NGD4uugpEmFyl0Ng3zjhJRGjP3dqpPC89XvOOnJUT
p3Mksxjr1doxne5WTf1Rj1LtRu4NZETmMTxPpDCowKUxECqEZ2HBaAXlJ/13Nz0p
rhAibhFcovkz0tNCBmXuzfsWnb1y3pq5aWFaN4xT/YwxOQ8yo+TKCwPoLBzMeX/3
AjcPWPX7dinpARQKlMasmnm1C2YKT7SVDnbbP5wiAPPGs26Lhy3mPG0az3G5U0lQ
QLSc6R4sBzPMUYRNXLaG2zndf93omb/hRF9IBIj42iXZcs57Kg9gnwT0zmsIJW0v
3D0h/7VAkpAG7e9Jmb4N//x87X1Xmi56RuEC/6rrOTG9q8jyCjLdrtVR5T2GsZ30
NOtu4LN944FHIHTnOq0au1sepvkYUkK8dPXjxDCw8d+k3ZiyhiO/Vss7AdJQsgKz
nJhr505dErBxMpA+rCrhSE1sVGkk/f8Z2B4WiagZynleRRhRr9MnqRV7AbmcY3/8
pc+BeuMKpyWFvyl1/mV2PJgxnZ69FVROBzwHN+BKBMkmE5E8gp5MxLz4WTL5HljH
JTtpU3HtlHLsfXYx6CNfIH4Du3W7VSI5R8i0hYRZ7PImt0iaXKTpf5zM2scZlLP2
dk/zoyeU+XdxRLP8glWkQuru0I5wxaT5ksl0RAHCqmbOud+QEBzqe+b2yWT6rO7a
Y0qvrQqlgoMU0oPpAVeHpC7ovoBPjp/YVvJzt9f2iNbjAlPPWrtkRXlxE2E7RKs/
nAFSx9hJ2KNrFavmTFLTEQ67MhwCzCUAII5R+myQwsIaJwvPfc6vqY7HGovXX5ox
GMg4sa9K9SdoGP1D763A+BwEUj29ZmDvyP1x0IKCtgpmt5pqeATDsInXdQ3iEGXj
hE6DsjoqwIciZdCKxe/JSC09uRcu7FUkpNMJ4wpaLbwndcmC1QWPXSTbD/INNiiZ
o1q7x+x0ZH+K3n2bUEPqOTVJfKdFIA75HXJjsPPiozrp/ruE/EhBcy6B4nVJkJ45
qd1DNG8Fd3CIhlmUFZBSDY8UF4CrsntguyhcKJWIAEjmPHH60Y/jsA2f7sIMLt6Y
ENa6OXdUGF3f/AtL6JMLkA76xmvPCWdgb0WSDw0OhYcbKsiqTltD4Ude7UA0p7WO
SH3D1rY57Pa4NKXsYnHkpQGcb4Gl4hApgjuWWVwuz7Nu372bEhln4XQdRnTWF3K5
Jyu8Mmwn8EKeCqFfk1mFSgxoz5JpjtyW4+Z2XsHCMaBfJi31Znp66DFvKAW+MAYh
qVveswKFI2Bifi+MHEUxqkPBcgNE5X520V7oLQDbLDQ12cZ/75kZiZXEY7CQUArt
a9QRqKlxhiMqiHTvIwwdpHNNHpaDCgeF0WpZMSd3k4zHD6V7W9aYSBXQeAN1rb86
noiKd+s76Uy3pF9PJEtmKwbbcqURq3+H52u4ylyX8RncNid9IZfA+n2fYOeI+a7X
HmuffQEq8aPKjzLTLPQuzGmsZBJxn9tmN5Mk9q0cfJ816F9kTsGBpKB5VhHEcpxO
v+BjisiarDI29G198WgL5jB/pk+EIB5Bf1Nu7pP0W2njzATVQOuOrqkrkjrqLXTi
GbGFdOUT7ZcYQn8ZA8xNLG4wA2PUURu4Ac28OCE36m2j9qQFY3Uzmh7yRA+VkJ1y
306yyPIsoaZSVrM7HyLbSLGpHPViop97QLJMoIyUocvdb1AMmhLQf/hdEBKQXIat
yrc4t6W1h9uoE79FiC2OVYYETYrHsPuCqS2tiRNY73reuAWT8/V0pE3m0g50O/i6
xLYNSwjv7DpZXcK1wADRUD1VvkI6gjXoDg+IXcyyX2Nra1HzLjNh/OdP3qFp4fPM
lsmhkndUrTc8nxMqzJz+LXXdEIy1P2xFIkbx+lgjzVevAwkBaynW2DqYRryttnzw
OnIBqudjEgwFTJoqo0YBK30KJc4PCgZbWg0kDtYJ1WNH9wBnYleDdKn9XuVOLNCv
iwVq0Z4J0tb05lz2xXS35jcubjEMAgz4VfwGZLrzF8jmvVGBoOO1zfJsNrfLEaxH
M4URFyg3vtB9Ap8gDd+gRfZV6scWvdWjt02QsKiY5TYBrxuxydsdJisjv2XcjrIF
tBpJZZjbx7A9qRh7GzF3xkjKPi8zbDW1xmZtgobgzUDx6XnamjErYNupY/NOXYpm
hrJuWf54OJec+2ZaOBdsbVVWbpW4076+p6GROM54kBeCKHLzh1ewzKByz1i7Erqn
keQ9eneiKQ46RpQeynN2Eg1JY5u7BE7sCyR49/KRmrnL4du32hVYAJlaW5AReb3s
DGnuKTob6PowxWwRhcBW6beCSQjqHfeqLhNB1Rws0C2dH5a5+oO0hFKYaD444MLH
Q1M7w5OhDlL/EE0fZmuJ5QWzEChY4fwt+HREUbeoiAGD5ThstbzgnZL/UH/2oDCG
IZToAP2wDuyAHYTs2+1dI9DfdGlWZKv5zoT5L4m1zf7u5RxskffkRjHCizQ+KQig
5JfkVazg8SLrea1H9pCQ2C7MvZKZ+qSF9RrmZFtkLGdJ2i6YQwg1lyaoEsWXv7jS
TjQxR9zlbmES2TdYZeNmo9frBW8JluCr19wgmioNlz2a63XQhqwq/brZgKOHwSQl
lgl7tnPRiSRyE+f/6typUz1Ts+UfhtK9ZK+aqrCt92h+21F9o013g0drMnVVdMyy
Zp2aleTdHYnGQyWp/SyvbZ84cP06BUPaPx69T6MZkMbl76aWft2U/6lHSxsvg/6J
oAaSpU7ZH1a6DdIAtjMfMhmkhuHfFrVd/iNa107wTxV6DFmbP4h9hY5lWjG7SzoQ
0iZ27wmDMqLnMHQXfx+SNgr6Ewa/vnWlDAUxvbLobAKccTsEUfvwB8QiiD4nbY+S
f/KK0Q/WbKgZD6Xzi0pb7XgEpojufeXkZif7Gdrx8ECTvYmQsO/7zxc9MMXpGQgh
HqXXCMHrDzTfvAbclVuMiX0u+ud119cSmaFFv5GXY0zaeoYHbMgDSxJ4LEJhMWH6
346vuvj1oosQI9GQZcVVqdowlodyX5yctvU9+T4RmeLEqAwplTUr5En62VcesY7Y
vhiCa0T0I0B7TfM9jGpXRTiVLSqK809Rvj2jJdcDm6EDn4MJvW06inO73FIrxDqH
BpIvkpkC5Blb9jPOIF8bGC2BUwwCH3maLXC+CSMGUrPv6/ft3DsSMojcL6I7dbsb
Cigz2tPDibld/sv3idmEZj/JFYx2DcEvT6PFeF4NGaSjbb6vpHXwgNVobZNAH/gu
igPaAxlnvl7vEih6vruGFqGvakaUDA7bNl99tmHmMYKadjKlZ+zp1KL5hbkLzbui
3uMECXmZ9n/FH3TXNfNu+XH7g5v2B+YVG2Q90yTpO7GVg7p/JrhG2fbTsEyRvAsJ
yzibSAJIfRgl22QohSswYw1IVKqcR+Y8iL0T3zp1Ze5RBX2JO39q2l/KxLEjJ5TH
VJbltzQDgFqrykg7+V+P1cLwYNeAG/2KmLQyhl99r5eqG7YYWwYO2cJsg4E+mMhX
PxfNnri5lOU4ozG5GJu7djpPoy2TLOgOYJoXrxbOFrTi3VfPyfHk+DEn2FzSY6A1
sbbzXcCj51M2uP2l62f7LjRayta6480NkYdeLAoU8OwjcOKlJoZgK/wVpMteek++
urn7TdXBEu8ViL6dVMWdaeQcsSxaM3lk1B+dj+mRQHYoqcCcXmNVVJWVd1Or7VMU
KAVW/Q1O+UBirwwaLgG4CsnKHJOcJnLQu7H4oklk4q6gIktkPh/xbqBlhnHKzpSZ
WSXRajTjFMjXlAZRXBwa+EJFYA+uO8/FjwfNjugcJioRE+IWEBfYDZXNn4ll9WPL
IZL2uSomzJstI2Yuw2qaY8DLlEGnO6/3YFVRaJBIoOpAtZ5LJtYwXxNWBB5dHDYq
p9KZpy3U+QITO4xv6LiCJ09YxoUpz1WPhIWTWeAEKhF05A23gDWtRFAb1fd7QL6i
7eEHFF5W48cquXdX6u+5lQGGzL9hkyqqZsWDFVvLGon98LRTUQ6DNtg9IxCWrTYV
IgooyvZiuIrEVaVFPk8rwye8tjZQD1wC/8gwR8rnu5FlrZ3Z5wGgSJeX1Av5J5Ub
FI3qD3+qzfSGl08K8FMGNPTVEhe5U4PtatmzpHEF05sIMr7GaP9TAE2vpYD6erCy
Zs6FdXHMC0Lih9wPw2hdWQgP4Ri2OFxfzyyAPVOrb5eU0xmtrjzO5FEMKK4UqJcY
A/hKfetoDVPgGUZvcmUUiYoRtTPmOpvzSdXTpPa5CRpL5sL9dtZxCZh0fde0QkWL
o2i4UFk8dRJHVwlqaJr+BNiBp0pcYnVvuu6gJMIJiBwSpD0LQhcR5hpU+50OO90p
GVUJKbqbnmeyuVtljSeAV2yJcH3B8Jx4cDkPTUgiRpyYfOyihK6yQBpjvzSzOv2H
xq7kymlslFwHGzZRCCt2c+VL8FKyP2MKULJ3ee+MPMZCW+1OeJBVKq0FN7tR8t3z
FL/G44ShMgDdIjuMc/Op78Nf98dxVU3UVuN9aRx2wqnS1CrwdcOU4EyFXS3bMoh4
usX8uJPyf34mjF4ssnEpIYjjCRsHa1mFCl2DC9y3qbhhSz86Pyzl20r50v4bnIi4
Pq7gfrN0br69+mhK6GPArVTW2AR7Wj4r7KupMWWAhrAe6XJjsHFOtfv4fhdntR8c
5AZj4/on6/lPQZKmiFXHvlWmQMNuOwXpYhdBsXN5Q55vXoLTXBoDGwedrBQAGRw1
IutAfNWWuqY7TLDEIE9Epm/IEjDkUjqPeg4DRsi22wARzd0cbmPRdtJ2y7gCfpCI
vUZ3hxFGrVB+1O/c1Bt+4jB74bwPvT6qlo2CA8ZVhRNDyHxhjjWvz8IHRAnna+6y
j52IC3En7aAZPgZDryoWeH4YgyrGcHIlPh6XhRtH0rDwiedQ1Kw7cS9TV4p4rSbp
Fg/u+WMA4SWcUVKMs8miItGUr2rpZNwHDv2yu83SYB4kAOyuVNsZG/auA8ICG75m
KuluL9cPqprTMK+aTxmKMMy7g4hxCIr3ZDeTncy1dblW8s/eAm1FtxApGCx2Vbpp
iLJD9OXX346d3ToCNdpWKaEPshSWJYz2y9UsPMbZrgwMww7UPNQXTO2UmiHi8ud/
sdzgF7PjEZAYDAziNMNN+utrRjga+rqN8Hs+j+AxxJ2MIvs6pT6z7jxI6kZkf1Ku
oEn+11FgMSB4Fy9OJw40zPQ/LUDfcp0polJPUwqd7N64a3a6p7ZRHyw52EX4+Zff
hZ1EFkQgY7eilF7LJAKDSduKaal1sKQi+202jAq+6Fpbw2Fu8lpCOS4+FHdlHBDZ
tmGYTy0Y9VoU46muihVt7RcnSsNsxHvaP0ZDuffRTxZ5MdWLgHOh7+bhvvFEJvKg
LOFT37dygKtdp7Hvkegj84ogXaR6aY5BPw5RWV3AaxzNgy90TmTMRNSO7ROF5niB
sIyAXZMpoplEYy8qLQkuWI/SjkORlnUJbai8QE+E1Ys0U07CoPsJWQQN2dAjnnzX
HzekNC7Tzth4FXPKrWZxvvCGxZ7xJeRsfCeKnyQSRuZVPFj2STGT+xjtKLfgRkTS
4Azb7ga8tQpH6Bby2PlrmR1XJpTnGAScUs0hYN7lEq9jSPS+FtkjZ2mh3YBXFLEN
0AB98K9rY8mbXOqPNDARzyYyJNiEWT6ldZxKs0Z798aqaKxSIC/1E9eV5kGCJgAp
TjDR/iv9YqbMC93NgsR48WMnc33kPqjnY/WZkCs3Lbgup6eAYmBzD8V3LQGMXDTZ
g26hM2pL2a//spqHX9pxr/ZnPu12fzYIvkLIez1HNKbs/HMjpeqGEIXavoM5NViP
vg7Mg3+U8t+6brs3AUD9oujLrucmg6m8wye/I6QEK7o4XRRQK39CVi5MYu/GAJg0
2dRslPyUsuV6bK7ddWrXcIPtcmyBIRHXImylKWp5kbTXnk+w59Um1jm5eOcPACEB
OtuqtG4kFt2RzTCNITcQVuHokLH6g/DUN0vH6S2iLHsdrZfWYEnybuHWp88qLIVH
CvqS4T0HHGH7X4RNxy+UBhG/xWr5dwDQPYCw89X///m+OiIWOyLlcaq5AoGTLsdN
8nJqdpaoBFCBRVw2W9x7ez+yT4iriui2ee//JlzYWUsVeOOX1ZKboilMpV5Uh4WU
EEUVknz89RfdLDJ3Df8hnIByByVOWnm6ze6BlLsNyHdtsS7YzVtQ4H4pxyEgQB3B
QGufWfZ6Ge+rxaoK0NJFSS4lz11hI7MG5uVOTfbBKPe/t9B+eRKriiu2XX45o5XP
uXuVp16OYGSSVI14RBbvtavOg+p8do0vMMCTkKSRKbtVJ3TLCJwIIS0QxeoYjYPz
ATgLh2UnvggHE9lY4Erjy8a8/aDwtwrP3RUC21gGaCzij+YlX23LhimjAo+WTY/6
a9RYChQUKUFZEuGv/Giz1N22TvzyP59hDoHGrHlLqRdl1xQsPglLuCVEkLcNQyIS
64842198WGlVuUcR4Zh3sYRxBlXIcy5r6CvFnRsiEHSr9VUhmhbzCjM1JdK/G/0p
YBLle0uulqQ87oUp9W/djiXq3hOF+NHEp4ua2sJr0d2qJTF23ny3p81hlZVfBQZt
Y8KVlZtLvl+pt9BZu7bJmmJTWuXoChrhbKqzvtA/0yMrPghl6+vr43JlbdKh5nkq
hXDgiMl2V/5Q/BM2yv6kU9gFFWDdPOsVEg6kM1C05ANtLEJemttcfZ44ksCBWrG/
XkxCb/Mkt8hoY0TscVEWg1xWBJ7LwOGvMsr3auAAqeWpPND5GRWEsg8zAX+cR7UH
UaIPIg0W/ZE7rMFIePiQ4L+qbGvzUQq/5hZHp+lP8iVT7tQ1+Pny3OpubFqGl7zZ
YTx3Toz8cnAYkcHzC+OQ9Q02YTod+bmwedKyt6P+zPxLN+JU4dIFCK4G1n/wcRei
2NNM1nr8fjNj/x/YpXl/SciOtFEBrttJO79eYoDekP+N2KSdnbmHmywlcyQ/+shR
1Rs0XlAGOfphYTFrLEzEECc10wQHp/0EsYR39RjyAVdpuaA5bM1iPClh/wds5kH2
awEkAQPQ8QiwQXKW8DxJCusU57lcmWuInlEJ7UUPwPdrqIExAdxMjGDiCLKzRMW+
G3qj8en+fhjCaeyhH4oL6BkTJkoxIpTlU/WTcTWq6B8tx7lgtIS2uATrZgAtUBa/
bbm0Xqye+86f20y2Nslxlhtn9Y4gybJ012gvcwDCHBWfWogbA9KrJGHw+v6r0uAd
QLdVeEJpAb6vhheesJCh4hUOblkA7PXTcEVWEdkzi5LzjD9TlVJc7fURboLc735D
ghs3ICKxSNqB9GMMnoAlixyqDOX5ucBa5ToZY7Sqc3O/1c+XHD0NUnbf1BhoxgNO
9EaaJdwp+SESCMb3DbBXmTKjakc6IgFqWWf9n+PioIwkQb75IKySMG8EJd0FxllZ
B4ojU041aXPTiyhG3B/uTMwrKrBEcoU0mVI8jTe53HwkXlhJ9LreiUvNilSruyNU
Triyc+ugkbv6uGD3kVR/Ic+r39xUZ3FIczIcs/db/ePuhsqL89t8qxcah6+6DdUz
DLqfvq6D30cN2nhm7XhEVWuYfsVLiZ7wpJWGOTP+w8GcUFX3cyGsVkaTt3EiUwH6
As7uGXdrwLPLVxnYPc1AyVtBgbhR566fy/0WjfU3lp7R/PWRRS8lT0eMvmXEBN3c
gROiire+Y1rjoqgo5qU1dkLQFfb98JjeSuuPZ+kF+KsKCumLYCKLiR+nk2XT4NJj
Rz0nVHbpAp33Acqx4jJNPw44VgfKHA/wSeWhgaBlFlkuS41ygzs46KgtdrO9gyFb
pxIorsCkXBB7dt/jK94X1/2y+eMlBc/JqQQ4xzBk0mWZ3WJl/coS2+Fi0tkA5WH3
mK4Kn9fNVdv5sJtJJ7NPDUAEgAtwS85zCY+hJSXq8Z8xWbKDs5XfLnwg8/B11wOM
JHmcJEaKv6jv4nkBdJO7QV4V+PKBXKoOPnGxT8GLrDvB3Tm40njTaJonfO8KBsVY
gToEuHBSEHm5BxBdkGsYtinG5qadj6QsmAH2Bh3Xsq9IOKW4GatgLykZ8jqYNBPn
n39bgrWju0FVMEjW3R0gqPwhpaUrcCem0b+bkz4SbrcsTukC2dMdTTMbGxHySwqB
4jQs9ceegU1crBezdGjwislru+95prGlDhTGB+0ydWOPOZeW2w1A8RbU0t+ZCpJo
EfHQiaAKAdkXCWiuLrEn3juPfhyvvpOr6xi37My09BFNOS0npf03BgHqmcFv53b/
eSiq0RfM7KkyiMuGnPaOUoH+RTmcUQRGNDd3DFM3f9tMSZBlEU6HO1BNGzJsKFce
teFrqUi8kCiQnZPq+nUOy7uLL77Rd3OLvLvOPDvyIM0ANgeXklWeBxEfV4EUIlxE
UUj4uT2+L58b5GhAP0zqlNHSsgJD5coJ9Gn3yuHRi3lkSDGBusnIjwUk62S5JQcj
MSA48fa4Ghh2NSxPa/wclGhbZSbTWC3d0PJgi5tJsHhg0XRDxJhdCcXITcgycKuT
TdX7KdmGX99Ne4ryKSVn/XUA2ixfe4l+CS8+Nz6VO3qy3lwF5EQj6tRsccBlMZqW
J422u+7+v5Vb0gRoaKn95x0A9+yR2iI+3i3h/gxyNJCNpWB5c9UgEYwCwfkltkkZ
DAPew+nV8zG6IYPchSPElgGEukxV8Ba7iVDrEsCBC8h1dYI02k92NVgbZ17r3rm6
XsW073YxYk7IZHrJTGYQnLv8A7nLs5bx7gDdIMyXS8N/5/zvNhuuLC6W9kEmLqas
0HFmu4bcuZDm0bc3Cjf2ymxXGKak1OjfOqUkGBaTRl978oHZjsgx+ElT2E9dXrCD
hMVG4WQ/40mDhKuSPg31NDNO5nhn8x4DVkbdovVmMuERBVhGRqme9XVUMksGussL
1ER3hbq8nRen4RBQnGEkwoWWG89QDIXcAdgjBsITGHe8SbyicS2x8OUkHxKQJeC+
HtsaIfusYRUqRpSBQLqKxGVk9YLUyrExEmdvD6ioO3SyDY4whkabgovMHHgit+uz
ZRdE8RMSMBuczIK7kj55JG/HEgfHHnq3zvL+toGcndjFM+pq4eyXuz/9uN7b6FWI
cGE/z4HlwY0lBOmBUf8086LFVfFcSbxQ5+27m1AkHVSFsm4++CQjp8IXl/uYADhU
AcNl9MHgbMBrf+jCy2IuKuc3A/iUE+OfyOWoZC4RAMzTeot1Duqjj4F4pRir98Zs
F6wxXrF/A8hsbuOczX7wAjrQ+bMA84ci7qMVCftN17kG2Gr4YnPp1nKdsKG1wr+r
3ULOIgdRxlKWWbuG2lK2aaNkPL/IVEiR6D8S23LSJu42RWE5MyacLdV+RmiBRW1B
8MyiDkgWLllS/tEm56k/pOswfgIRgbdofxqaHwEMkCVRHl4OwWqeQbpYoiPCPBRp
ZcOcyt0SpRUK5KzJFldPQViOEMO2Tzi9kAsT7v17jfpNTSlsJYmpizmSsUU0sKyH
8EALo0ID1NuJ7GndM2hMvhk8yJIGX0mNfoa+MLh7DQVG2+BKnxRi0R0zl3+qhk9a
pF5QrmvOfijIxCbqT5b3cKWUJ1g05kOpuBRyZcprKGTcM6QSnAdgQMMnBVzIaRpu
ByfxNjHlwBQn0ef/SYx+bkKKX9G+Ctu5E8P5Il9Sl55QdiMhoBlMr2aqvtJEtfqv
VcHcsRqIRVCBMKfFsX5szpV8YT/UMfQbW3Gr48vKz2zlIrSVdOXj3opIh8iFJiRr
yJdApwcYep0hmrdwmjWpGYAp+YwPKgPgS7gLDLDVICdVDTz6/vHwyL1zB8HmZeZA
gVdbUDFiEKtsP2/TmvnYWFvA9mLDz1VobFZ4lgX5Aj1k30/VcPv14CnOZrcsXAsP
TmMrCaWGCpo5wQazjzNjKtC9Xa9/E5Iv/DKZe+DXNU9iWdLdchTCMCP3MSh5G8m0
SiSQ76b5c1yhRFZA4tK6HH1bmzWyFBm3MPNShXI1jsV6lz0n8v2aA1d96PvnaK5o
vKk/mgVjqZndjkU7Ut9HwEtgfG7IrXuIEqJidO2m9hVR9cDcXSMKVuX/9mzRslFX
OypBtuLQokQkJT6gsSJtnUIvB+g6uLht3BJKAgPyT1wyFZixZYMvOjxCsDYDCCNF
o4tpe92ckidkbEGuVpgGWtqjCKim7/dBEGIzWS+mUaYZDrYNg0h0KIfak73ynD7U
HtialiuyYzgNVapvX8DiIv+HK6Kf2JOwtQxk9zNIGiIveYhm2t9AbR+RB8Rgj+PV
Nk62oDqltgZP186XRgA5arG4DJTMZpIzESsmLp8g1WHhwTfDXXAnDXoQdd725p1r
DQ3dsmXFpHRf5Df1h97oLwyniuhjRMfkfgZiPufkroRj1uLLZGQDYysJRmknMmz4
ggXF8ocmw4/qgZWh6fXWSWXrZTK1uOb7bAQEWdz5NHpv/Tu1PgRvAHWuJMNd4Z+N
0VgZg48Fj7xJPqfLzKo402CLyikj+YsiLRdst9nFMw8TrN/6wZgS3xXAHxKopekS
rj8u/uPmz1GKQgX6Hbgqk19p/VHX/bVTyqKRvNC3r2UQ9CgO4T53xQ+vIqdx5wng
ZW6BqavY/GfYDhUm8dfN9LVEHspvDW6xwgjI3kYi5BB6Wu6Wt3JfvbzANgvZxHl4
RaQ1sGumiiUBZZxWgJ+/ycvI8HQAE6309PQmsOMptSxiVWvOwbpuMzebooMBy1E6
9zhoUI14vqgLAVoz7v9hmw9nyQoIqSCFWCOyQq2pVPkWpmia35cvmmWXic26WRkA
rYUtJdAid7JuKsVrNhO13ITekRAYoHQWKd/D6vJrr12vuQSWYQaGfJOufTUhMAeZ
gxc7H9gnrmaubiBXSaae4rtZqo8EtAZXoWM1+OJQ0gBKUf9tcr5X7GeGaegEuwOw
n9Kgw3HvnK/dujnYsYTCy6r7ILvJK4pjaQJldymKDdO6WPOr6X3Xahjgcoyt93Pc
miGtuF28qQ9br0hMygE2iTkg8hvsdP6SJGDC4COsiFGxJqDGcSW32nupIc27i62B
05yYL8irAVLCpki8ThBTkJMd9FWFKsmM9Gw17HxRs15SHNOV+E7CsaAO6DAGag2v
p424eHI7dmV5GsWVcZr2g2WsapcfKqs78QijhmkBj7WewoV9Hk6GP0LkXRsfpawz
K/jDDjg9IKmi/8hfK2x+nrg2WegpovdieQNHORKIrwRNBNP5K/kfVkk3IoM/IpqC
vEFuI5nrPoP388DLGJAeVk3AS5LdblF8dFcL/cSIJIdfeYv8DghOdgKN2QpRkfg8
zYIiWOc0AdnKTnnBS7dc6ZAgiYRMgNSHXHHi1vj9Clwc2+QhbMtIYymq9c38VJe6
VQZS8URzUX0E5tgHRycJs5Y8Tea0HUIXr0hpRUdVLS9gIW7pliix+/2OeKmgM8Tf
7izgXbZJB7lFyvrbxOCruNXNJs1rU8zFguHj0qB0T85fguwLvXE2UFFTpoe9HH1t
eykx0kdL3Xm32mCr9LgO+TN4zhOw2XEZDrwulgVHTEUSaLcWGU7CsI+8WqY2w1Nc
Ju6d3lrNO67RHOroWEZKLYLAJG6MGvxnk3mJdonjYLkwRefB1RfE6/a+48KgixNl
YfOtwjSXCK7PFdHV/HisjMUqQpBp9p5aj+xFgUYL4hoAasthOSkm8eENn6bw19Bx
PVcYYk5q58RDU5Oy9H1tIBKlTwnQh5Tshxm0Fb3Nvk1t7YR5daxi41hh1MzKWWqZ
Bdlec0yq9d8pJwhjHXMCm8z6943y4nrnNE8n+d/BU47tB6DpIfwlMSFq1M5j9j/v
LNbf49A46hn/jTpbaboyiIE4cFI3a3BI3yGjiQCDCn0FbwQa+ihIAhnw5m4easFj
Lat/Mq8AD3SCkkLc91vWKWK2wZIiFl+gLO5JwCmadD2dJIviR0uOyUWkw/lCYC4Q
dF1g8HvqnDlYg2/Qe+LF/vWmsSe7hzULyEO/UdXwqC4y4bP4Kd1DI/opzAfVs0dr
NWqiqyRAWdhuzuZ0FBBDJBnKbhA/jQIHPRT+WVtIP+dSU3ZeRbrZNfzQyS5fMdXx
PJUfItuwbVd43VsfqgBbTF/Ydm93J8p+tx3m+xsmm82UrmgT9Q+B5LGBe9pWfh4Z
iPNNOuA7VC5crSmGRkwO8lzQC+NwAW2He5yMiOV9rkgHFtJhNUl8SzWozR7we/oV
+rm6QUd7TAdAmiNsqkEyWTQcSdFghrhaqB3ZrflPow+pX5xvJYMxFbSqdBNxYxhE
c+NrvUbp/kklAJskJ+3T+A2fhhDi712QISMmixbRZrHeQhdf+RA4EZMDuFuY8Gm/
rcOz50xwg9bUIvGzO2GtbBsEUsO+u/LrBOxRkQMGV79B9pmR1wrM2Ic/1F2bjlbz
GVi/qgAfgjjpizeLjhyag1YIEtc2jzhNkzavYd0fJnpgcFPxkPZDIfEAQkF05Gmh
9nbHouctsko56ajwMXEC+Z749qZ86qeSANq73SVhJ3RAT8+pPALMmISfqkp4p4NT
fWe9OUy2psZ9Bm2wzbLvnjbKot1xCAp8PyFbgKsTgc7EirdfZfKsyELZKnY9cr9V
HAmHCr06UmA9HsA6wPuetkyIIRpWnwoTFCmIJQfR6BC8Fa+YV/bnUPKR/lCZlzy4
OAA48a/+l07TexMYbFbWz/kPFjKrE4dQCNYhw2AipOTlprN5Wk2rCNdxZB87FfRn
RRmMKCZN2pD3IbwtUczqiWGH4C1bYaPiJQbGW9neS4EHw7NIqofyAgpQ/3lkHX4O
kE4lpvA+jKLchNFqkHSbVykeqcOWQHRPhTKYeEqK8kfIOL6vEMrJhEg5fipohQZB
j1vE1a/u67IWlkKydQ86FOF5lJfoJ1tj0w+owDpb4PJbiAWgFbeUq5r9ouY9XpAr
AyQw/ltzRAEjCqYN6U4g4VCzhKeXcAnH1Hjn514px63j9ZjdPeUdrdp1iwXXnpUz
6ta/l5X8X9yaOrYBN+TC1+1P57+aVpXfV2L/Js0DkpJ3Tzjp+WiThamiaGxZFPKH
GSqYAnz4ZKHiT4MSbHN7KoOWlTz0zlfrx0raVvACXSUS3s9Pb6nBWRtcqF66ePKs
VDmJZ5VRWHW/nmwRBks2MpKkn11LiXRTWg0cmMz9K4in3Djm7YOf154AEWa4QSYJ
o3AiJanHWyjPoWo0yWPOCM8v0/pRRPtYHF5bZ4L6Qd2uG7WT0EN371Om1eNXDnSs
zsPpK7pLuPXj7S71bEuGW1am8vbwSmlG9SzY4KtWRtdQuncXJ+QUwi1XEL+YDe6P
5x19zTwKysMJgitw6JG5XgpLxOWK4qEVNTCyJ4hNgVKdkOltx1NY8AWsW4hdXRYa
GBBkWstPhwuNUUxM8r3zRJuMlQVi8xrhxrhVP65XIBFmfXNjOir7pBCDPFKbA0Rp
gUi9gPLYDzYWatLxlMAj+joGYcQdsyASPhry75g8gtcxuhIVgBzYukaMWn+M9Dao
1X67kqoWDGeXuoGkJDlWotd4chRYLDnUTS0HA1qE+Nc9Wx19OVGC3tBaR0oGDAXL
bE6wPxQs4FNmFaqhcOcAP3Rc1oZRPhbAzfN/07x0fUfrpSkRfeUyh4ete9DLeehp
NHSEOJe3sV/ohG1cozXJVWO7d4CAaGwKK4DWPvg9jYxbeCycYSGOXSJMVSAakqH5
gjMP+eUOfVC5RVAQd5ufXjM2ZEPX5B122MNLMCSkEZHg3R2VruCPpjiBPrqhMa5V
NgICQa6fFJh0NdGVdaO8OGDsPBWiiyAOpdMbAzLPmVNoIk6dq1JkC39pNLr5sXaH
yk94GVi0/HcHMl5b8mSH8t1jiNkIdRjkfn3bczZVjWe9enzpwRdcMhGR+RPRjY/Y
m2uO28BZjURHguOEp3wZwkSZMe7spaLoavRr9HYAuJvT/bYUFO6ykjrJjkovUWTH
83tBCTt4RmF0PDPCktqwFlZNUmsp0f7+g23K14fFeJN62iqMvFzi8tQOvyzYzLhu
QgH87ARJaFukmyAfXhosvddLoMGT0Tt4aOYIig3X1fbz8mDLHbLVPLZJ3nBSPt3G
leukZOYGxP+ywXsHOvTFoJAPsWr67+mHqAt/dzSmUaD+sTIccg8/rcBK7S5B9LXO
7fpyiRYsqjAIyipbr+pLjv242dX7iUc2NnZfzRPOys3wCD+leW4B2E5DUvi/7Pl1
547cCOqBoGOGbSiVQEIcY1OE4XeqF0p2pGnWhhkH6z7gg752XywYJQrMGxMT3jtO
eZ2qKmxHbg5idOCrgS4YKtwPdRFcHyhPCXiB4CyIWN248AWA/0IN0PZIH2WIJ0JL
C5kJ6ig4COMyDHcI1C6GAdJikMDX/abxLpMcI3ZnOfvHv5jKzXPUv31aKVL9C573
v9awfYvk9guMZYmd2NgdlyiknV2i065LCv42W9mZeeTvAQyMnbnlWsrrN71onugU
pPc5/jarHD5rB0tyoZSWIdVi9Dxmwb/h0gEkGnedPDW1xxGTT79mxhne05J4ciZC
03kartWUERWRnj9FoWPlISq64GUUODg/ZYyES0epmhxuscGRuX4pZwHD9gZyxr++
KNntGx2Gu+0mulpsiB5kUK5M32MeN0NX6v1/HNGixv0mhP3clSGUqa+Cy5PZMa+M
nbraMnY6kLdWWUePO/KUNRnpD1HtKHV5oMUesDFyS6XT5OsgDkLgHwe22LBuN82y
a1L8CMKFQ1PoGCggoAhesM1qbVkU+WfPFfbKz1amhQFYjXzO5wdO3M19PNG1vJIz
q7b4IQEMEZgTMl2VRm9xsvOjJUY2wsPx1MrNkngLaQDDTBpipKolJn6fMKHWxfsn
JxFWbASUg+3uru1/vsKwhK9b/NhpytympQn6Y761iyutRufJ4LZC6wjlyK+Rrhbg
cDZX8xbTb/p1inzNLI59zSiwGBRYG0r8nAVHDqcBaL12hEPAaODMAyplmQhIEnPa
/WEVm8uZZkUMP6kxiDHRH3NCVgji83j+eMDbAKLk2BkNHYySoLthtM8OCFDnV9pD
e1XFywdMFkf+E6p7Z/NZ94diRHZgTGCdBdf1MfbRGwxDw3Xcm1Ya7UGYLbaAdMNn
huXDJBvQlu2b9JoExSKeU3IodGluF24RR3ywQGgG4hlHS+okY3UyygsbmhH+/bu/
R+Sdddd05q6cbcwAaTF/ya9bdiaGDCPTh0kDn+zhHzx/lanXx2PIzMkkVAA6Yyeb
U3CwxOcewOkJrgN8xCetqFX1mPH4Zod29IakDUelgw+/h0rWoBeF+O8tgh8p6U4K
YGBswdPJ+tlAcPcn7QzuTS8A0WnOpN3Wf/IgJrureTDiIRTgPbjfQPHkxAMuXrAq
n6koASDfiVpJnk0pwvoiH8O2hbsF+gNjOKErCS9e1Fg+qRhJRHPuMGKY+p2S6/Zs
CbdNL/TvcCaMFdV4ihLjTtoi+0bQXz70YMMtUoEqTFBfSmlVUE8tuxD/Qo+WC2KD
/M/L0PrymLp0907J+wREr7zQkvfxXnKrWZR9irluquaQA8cFxVCVXEIumY9TwSGV
MkRabVuhvgCmFUTYt+8n8L9ml9XUpzZETT2HgFgWldQz4Qjsvmxfs+D4AnkLdBR5
oFDv7g70Ro2yejkA/gzMq/sDs1vVpqf+7HLp2ASfAkJss7RKW2YUHv5q6PqHB/+h
tedpaZIVHv5H9kw/zPQmfVTHxBLHLXtnfc4IIFQMfe1CzhOhqsAmwyHr2gQ019ac
WNCBk0aZV2eLFxgzeikwIMT7d2oz02eEEI+jn14pSU4Se7gvdBz7W+cb4OzmESpr
KQUnm9uEwmQJuugZAdNJ1GUfOxDTpr+ibhc1NEbe/qkiPY58+H9FlJtdpA8Doymw
BUWK+OM4Jglsrr+R2dujxRwqAikPryGcFZzu5VMMuNTK9nbzGrrPlsjWuHBwmlbS
ZAbw354EhqFgXiPPMY28xAUV5WD9aJE7WEvOGunSsV88kjYzIMA5xntJXmQIXRxw
aEbwB7kU3wEvS7l+Ut3ynpCPke8FMryIskow6gkMPRS7kMR8QVMh+2iIDQF6iTz/
c4uZ5FiD48fX2S0R+nzyEuJno93W1J9QD76MNjpi9oTK2lUwKLBKQ9hQg6/LjWHr
RMdft0pQrcRJJB1XV5RKrTUCnU+bHkhov3IHZrGD7r4D7ypfFkDCHy01BqpcoTAc
Ng/kCWHmMGaOKfgqWjT8ZR6jYDYM2jamuJO4NtviGATitiv70v8vX+3gzUUDY2hE
V4V2YfCfKTYWuqZ4Vjf7748Q/P1UZFxXLcAznJNpffmrTWnvfhR7F1+E6U9xn1xd
NdWB6y9Elg1UkCSmp8ADpHquL3muY4lHEIpLntKqtYkdHjXGBAs4zTpHkCbD1lqk
6XFL6sKscqv3hvvBCNKAVCp2aar/L2foH7DFGw9MZ4Sl/FdfeonbcFK/fZ50pI8T
QyGua1tu3zPAGZ6G5ZoF4Nxo3veZZNoIVaS5wVbChTQgBYdnl8ELc2qtKb/amNh5
a4t+STvSSVAahwA1o0DpxS9jCQpvKgD42RIOeRU/S41cyWkZU69iYJf7/Bmeu5i5
A+kODp9baAhRXzey5EbV0TvLSdXDnOmIJE3roo2O2RDv8KEMZ9cq7MweLxSPeOs7
zYJzhS0GEp9Y0YQ+Fi1D+i/VkEdVUOJjh6Caphn9EJAnR5BppQRWBN/onW7QEfAM
3z+1gcG0aPW3Wh2sBhFBa0v9i8EIZVDATYr76+vsylXWr/umjQ+HowFgEizaqcIb
OFk6lMV0DyIDWNoh7dKVdbtz4ir6jcSylv/tY9YA5E8KaNcOGxl6D4pWZ0I4/0lN
yiqDdfIn4ldmP/2fGoNpW9WUGz6gvXJRrbN2hCOkqngcPeePVAn8LEXDnpQ9ow3Z
1GWAOCYXz26yk4d7YtdqiZTF3vwK419tl4kvrf65AscydgKAO3ZDF7Mm5FDIrDkG
+ierefPJIKQlPCVdSwv0J/oGDvlkSDUnMKQyPRABEC27TBgLIQ59XcjPb60BW0Hh
aGF1kMWom8Yt4BgdQMnnJv8x9BUQosw4JeiokRGjP1DVsJKyODdRUVRcCZfmJjjr
lXfb/0a3DGd/Ff6Apq2nad1f4z45NlNjeFHMCN7JBi6ydOe1f3HTA20GfGcZEjb4
Z29VAi0BsrN3KTA8U7bnb759fvi2tEcXiaWbQbOinZJW4gdJ1HCJNuUlxgHeS9cv
II+ThJ28TDf3t64UUo3Vx4i+SCHoT9wwQzvj74K55+J4X1JWNSoJDP/AmaMMB9GV
G2++Dp3Uua8LhhZ0k/UKKk97UaLaXFyUc7VMCfcRNIC1Hblbq9Dh9rntDT7i01+/
5HjOkiS9kgo3BvhLEA/BTMLFPKEcHV1OX/bYtIlkTOQ8lyuEJYpmlVLsQWQZPB6v
OAfhG58nW+O+tlI9/FxbkhfM+pnx6xYtJGz7n08eKCpGFNpp6YFCtW44O0g99/Y4
B9CkzJ1vV+rIo5ueQHxJ/trLkGFJvEg/o3gydnqKJjZht56au0V7LJjTE56XU6yp
Kzsbb9I71VGQmc7Rj6XOzpvAvW3zsoabCeKT9fXbFdUfQJAFoANf5jVZeSPNGqdp
n7fEuiltyhwAGARvYDyEVeD86AV0WyHfyL3YD0SldJA8Qde6o2S+frvoU3QEpnWo
SvZgEebB+fXT5f5/q6HYACANGpT0L8zxqsFhvFVJjelLvkm8XvZgmC2TB8/3m6Qm
OLg0s59eRam1R3DWaziC/n9x10PIFhIBir8uWV+yc9VzpL/yj9tY8AiM4eGAgdga
GB64mxRTxySIVnEXR17Fr3Av4f3wrvBEtW6ehJuiFXfaYTtAlzxxebmbH48eu1zC
FSmmVWB08Wc8RWSQPBRMstvdeRySgBXOijIb0X6aP32dYVXzYsgJ2A1JbHc8yBdN
h+8OkaKVY49Qz0S/BOI7qVQpFc2Et/JNZmA/6PmH0NSM5991kjY75VqBJN6wQJnT
ayqtAoRrzKvSHlCv/KqP0bTrgfVSoWbL0i6lki5sFioeYhOg9BNc2oo6kJ1TWt+H
Dp9a9JgWn0XUcD5ovhUU8TX3uQ2lKNcepBDoL/utsjQ3CUrx5PbQGg/zryKhK6iD
jAEMEDqFbWyKkulnQFE38B9VdKDXBCQBsDnIsXolTYMdDyQ8wmGbgqY5tkFLQntm
93FNXX4GzZhhw1HCOim76hfcEU1vHgnd4cyFAp/ZmQb473X7OIwNtYtnfS4wjc6h
qizZqixn8QQLuWGB2JHJb/r2QESyw5XtXeIFIlosqbukofvAF0njDSm1THau+Fcs
laA2St8PLOyU2xQ31oPov0U0ft2ZmNkD76zXDE/GxR77a771pK2LSxspr1MdL0gN
XEu/e+1F2cs9/SVZ+9GhflYzVACq7NgLWWdw1anmJzKs/5sIc5MqiNTlEl/r1UW4
N1WkQR4EFi3bWuBrXD2YUug3B3DpTAxxbDuQ4uraN+f2cEtB/IkcXuCPrr9N7TvU
RR0fVwWJHZNoBYOQR3LuLC+7n0CD8I7yuPbuRgFUYD24eOEeBy6ogOBCjpD3OFHR
1B4JAJSA6rAt4BafnbwqVfdWjslCrA0stcPJz/V15HXMFbbhePW1xSA0cmqVc9Ya
+SQkv6BpXFECJIm72vaHx7dgRrjsriwdkF5++WDKZKiLYmwaiQAEvEPiDq5Qw6Ue
uTycFqSZ8yc4at2qF8j/VZAsiqAISLXIGYHO7aB/XrF6qII+I4vj8H8FetaezuwI
MR05qYTsuviCvQ06a6oXP41IYuX8CYo1BEPqNEtHrCGJq72ldmSYPGFrMAoHdxeu
JRNS39sjm2nUVhv+YlxJEXWP70lcyjSF8ApkcPJdt/nq6uf2E93p/rjIKEgDvtgW
KZIQ2mZY7sWMXaHfWiJhF0eul8UUPOpR1vGTZfOcSDsxoEx+novrS/IVglrhaqvs
w0IBJjix/2yc/xCtLu+kMSRPS1lGM4kjHeMasfrCZSCW86RXLVtnUbMlbZHwQvJK
NyxgTmXjATa/DP/9n+wv9uxUCE6xlsKXjjKbOGk/AJwA7SXWlL9d10ECz+D2g6A8
lbZ3g8Egv2T4ikIPhE/h3V9QKgv7sz5oEhGiEeo/SR8uw+bOroMDazPQ9gD/0nla
GoDLzlsCcD9B96go2VBIwjXl/kQz177DDm+KIldiiDI3VYegY1bZ/ePSIPtavcZd
t+0sJsj84YV3SJzXaL6tCjsL1T6nwOgxYrRvs/vCDLAgKMZYRUcY0cwJq9DLLIHj
zmEc6KrSP2PPV/yCDdnXCkULeLndClmgZCeiPpvfuWhJDbfASB12Ubns9kJV95L4
qI13y27A2luu1nzVrrtAJE++gpqZEdpbswguSYemH1wf8Ndh1xkbRvsHRjrbD8wl
dexzzhvJjcvBDprQSIcQkbzb6Wd35+5Dfbgj0NSYOYfWHIyB+iNkDZ4/Q3ggPg4B
s27oKfuUD6aPZcqlNu9KSLJqTHjKYDfIuP+IM4pKDziC337n2NCs0pZIY7noimLM
6pJWKkPCtqxA6d9BPC5FBHuuHULG03b2IIh49AbgR2EBxgbIMmljRLWdY6D+ieBv
RCk0Bmgi367zPBGdt3AF8+4V2GPHgCt+4P9QLFeLt1AsceELvkBrSCK8MGidZ1Hp
ujsayU/52HIR6+jvprs7HLXYfxSBw4ZgQkpQ0pHdBNdiC8dcVPrR0Cqo0KmlDzY1
bUzWxN+B3Sqi58+BxucJ8E9OILTi8PajiAoon9uzLGFo4Q+BVo8G/Iis4zi02aqc
sKKjzob49zLCoX8wP72b8BDm0safY/oX5eiZaGT0lY16Dbb6kyPdH7qOB9rSkZrI
Z+SV1hzPcLhTDhaYK6A1DmNSJ3fqRqxEGpcEQg4dAPwsRCIOi9x71yrdJnlK0Dx2
yMTTkWueHGcXJ1l5EC8J4hahcr5xcukkfX4cBeoPoXeGGGCftmQV2BFhYN7cXcLD
TuuF+fzqo5DLo9G6/QpZMpB+1bXtqOVkqXU1SABhpOBgOpHHVTG+t3fOID+Slk3B
zwNvwSwybyoJZphtggJK0TWMNHztkSlTKGmhGPE/xuqs6ZL7kGpcKISEp1+GTnGV
1969ARj//2+AE/e7ObIqvZKIq+SemwCh/J9rizcYlpqKmDvvWcC7UcgOMsofsB1K
Gitp3NNXhdQxm1BvhzquXZoa8hedrFgzBofQYQAWF8mPyVIzjksWBlEPoXyzRynB
5V0V1RMeXeTpK4mgif/jI2x1OeqdCJmATqVgmZ2SK0V8gV0a+jikdT66HGgxgh0H
XeDVk8P8Lsbwv8KZmzz+aY8PB+VUtiEsvsx/ADxo0y7iHlNzeAlwg3ai779Km9jn
ZdjYxS+KhdtCwtX3UXHVFM155cnpbp4zz9YJsT4HxsDt00XWH98oNyjwTFVL+HdW
VluR4hHp7wo6LhhP3tzQto5/NohFkODxYh0Gkss8kW8kV8QzTB9IsmIG+/GL4TBz
je7ev/nH+G3LRooutxKULwA4/NwY/Mvs5Z5UjoZUPpwWrXxoXtXURioYnjylFK8I
aEAl/Gwnz7qGSt7Ok4FxkrL1mc22oF1RlkvHfLKH0eE4mI72Op0HMcKnmLz1bvv2
3re9JssZDdmoNqWjsDzsm/qHpUtzeRIado7XOaO7RSLmDaigBAkHDI8xeDNMo14V
fzofaoDwaFH9Deo8zya6GdecrFXBzAiwRaZpx40EgVyiNk/wuchkQjVrY4bESPdN
FJ+md9wEMK0i5zakq/r3YfQZ4zW928cAPj7aJ4WJGRNR17BYFyTa2U7yFwqu87jA
fdwx0zKNNrjYEAqQgzu6exy+0BKAOGHzlPP5dp78FWEKXucjlCUaLPejNFYzwUra
8Ekg+/ssGHFARTYIcLTguN3K2jLdrcyWBloJRLAvnR0HsBaM/gvTxuHYyi3XLlk+
WGNhPTPJg7AR/Vw0JfmLRd78KAbbIry7XbGfNoGUP7gGxYzf9s/Kw5thPa/0VbUW
3qGCWumNK0/kWYj9AKnl4zV9ScvQdlRTX+ukukguwc5FAgQchmbSIP/ZhzAyFXNA
gqYPDxfpBDAB/Pip5jzM8CYthpCHuSd5DPZcXmNXtrEgjXZuTmCs68bO/3d/4Qq5
QAziGupDWihS/ue6T0ilasi6sMSv+qyW+VZQ9bVGeNwUmugVmDO0bITgxFDfpeqn
ZE1LFz2DK8U8V+d/RENJDr0uiA86RB6OzoqlJ8pYcNATb8gusECaJ6gsYCrQOP7c
KGZsLr1+QylkCcPW/CP059eJKlgamooD5KUmFEuHYnMScq2YTFILZIpcRmEu5xo8
eFSWhFH2z7DcJE/1FahwLkB1boZhJZZSkHWfnYjmB08VXVMb0O3vZE5eqYnDp/4w
vh1qlPBmTOufsQOCO5CpcG6pZf0CeK8UbqIfWacwiLMA8RC+nM7s5wJN/b24amXo
piisOF6zujVBxi4IRTXbvvYNmmLihIdUcgK2NOCMDquGYXtQ6YcZ0vkiACtnkpZL
45alEMjOjRvlNZTUWwl2yTtrBwgRXrcqTm91yY+YOt0hlJNWYprh/MQQGuOq04qL
DNLXvVByHnHlxZeI8cQfarW6u+EY5nz0yM974Rzt+wwK9nWjV+jdAEkzfwneeJLR
kHyAlWBuV9pvQieGbVX3eKUVKa/LeeL5xJwhcui82pdN6HF7RD0zeBIy2SKerV0I
iF77njioy8oju3V4IeWj4Mv/cHgh2VtQvoynY4CceJNci/bzpsMKqzi3+NKE6RJr
lUsr+aEUfqassVKsY/GQmhbaF972c7oiGImTeLnBzlaI1rqELhWWnv1CBhZXWPCH
V0qsn1aacBueLoOuDXa6gW7v8TkynUAqzgsGGNGyfDNcE300i508Qxtv1drdwARX
2GM+KH1hs4ALMPrpEY8Giijy6Pgxm6MIhdFrz1Sm+7xDw2XbXpjbBPbwEB4kdpRQ
POPzed7sx4QMkf6X65FntWm3HVhzTUQVjWCyarg0CXjH1No3ye94Tvx4zRFNp1ai
nNNMknYJhzyzmO4ZprFc0mrNtTwCivI9+KdUekaMSMmBRAYGZkApCjtJGjabq6Tq
CHNNuZ+BW8f4djLjMugHUciZ/FEJJRKZ1nSitD+p41AbEa/D4ij/68Rt8PPDPX9x
Q2Zq3HQZ/ja60PobHDa8T4LEMIVI3+Yk9oB/X4BbvKol43A3i+5u3RRFOgfNHZjP
IgVMp056RL5jDr784eEUqIX9x231AGH7hpDDlHo4IT0kQH0q5jhBUZ51ieHIxL+q
GJr/tvQh5SXsyziFPN0mjYiBtRAsZhS4hdGQg3Z8u68H5A9VNq9N87TG9tDsN0XG
Dix9LZ9sg4nvWWTYkuMz7RTAzDWnXCMY/mB2F67erwLr0zXpX93SYfkL5qqnlqa/
ybYLt/bWZMnWQyEfykY4MZSMuTne09on7I2gL85Cq73SAr/TvNG6LO6ZGrIq+mwX
tn7mKTfREWMkAugnkhseQXu7pHZhhuzY5GLG2npbrh7hCHkItLyirflB8i8O5zTU
Z13aqlDKMjkjtlVY+3iQaZy3kSE59wqymPNZzthHbQpbPW9SYZ4H3dxD2MffKrrS
dSl/uADXZSDYiv9jkwXBCBCzNd30eLZpX3m20XLhDgt/9c0Nym8zuj7cqJTPno3g
ADifpH+xsFY49jl6AaH0w0Z275frFNJPGEL0TX6izbmewmB98ELZYRDriNxguEVq
uUz60p92oUFQ0M5mQ74G6pHLsfRUl5toU7mjbfCZNrTFvom2hoJq+9exMAtpiPUa
jWCH8gf/YXSOpD7se2V/A7Wme/GoJjbgn1atocXfu9NaUNawdgTZaaKSKwP0pYq4
3OpM41IiDmNXus5Z9T/RGRJvEkbgpwm5UODRIit+ax0rNAKsHCLYpYny/HlwSPKK
QgiV202qOsvXeOq/HoCIdcruFUEwSKw4fsA++0DFyaxV90sKyi7ny7txlvNyPN7M
iMynns2QfkEHslcK4EkJyBYg0HqJtK6xtAzF2ccC+7YEqDP4yeI2h/pE7kY+vpZt
zxyZtXY5JLeeH63ns0rSNl5FbvwSisH4JnclNB7vXMdycw5Lu+7EIEt854iZuRVa
ifEYbhtJHiFwzoXKBLzaCFci1WjzmS6kIxANuz3u93IYvUfBFLSZCwoPaJCH2tM8
FtD6m26EIBwLhx+p7+QMJafKklvac66bY1wsIKI2lQqyLpFx+XXU3c9Ltu/bZ+YT
o+RD/HVn0w9Z/9Korf8RuOmvXg0MGSRlZbj3KA9py+KGrIerY19c8lQvwqG1y/N+
jk4YyFioC62CgXtreNQ9e1MdvUYIb9VvRdkMT0G4MpP7jWKFfb/WjztEVBs7vLJa
VUN3UjuieNK+y8yOqn2qGDQanEkarb1341oNFsx9wfH9hNxiJ6koRXUUL6g4vIEV
pqvPqXgViRTbdNY+6jfJU++hzKG95XnTQ7vcvejqPzF1YuAQZjOGGTGEqLlXiYcf
yjnG2xRN6fvZeLTs19mA40XAu4O12XlhuNOdEyJ97LTjNTKU8vs6q4UdtlPnfyb/
4MPvUU2h11yoUWDBTyMCbm55uZSiD7hkhmQpFdZuVj321fBFyPKJOCuSI6YtgR98
b6c8xdxGvxRpMSFgALcBXBSYa8+tqnUimYB13c90J9RUBAAedneV1ggy2I+acERu
O7m4HS0nCJPnsXiafIEaYNlkgPB/5pSrVSipIY4Z6x6LuedwkEl/2LbO/tfIJmWF
NqU0ctl0/bo8z9B/BV5HUaWBNg9Vkyf2txC2a9ZLi7z1xZIDKOcS4NRm+QXK6Udl
/z8GPZ7MbFz7PtoEZ+XK9rYDETyKiy2Cff25a4JGnl/U5abh4AGoB0sOn3omRocj
60ToUmBbFoiM/1wAHefF35hWHDCXEkh+npeRw8ofzCn1P7B1pFuMyZkXPu0roKYw
ya93OF4hxS/E99ZnT7VVW3qp53eTc1IJuKgSwJVvEZjGNycFnmlq4Mr25QBYvzma
Xc44Dut8TIQdqaxS4sVEB4gSqFL86GjBHrthqL37HaBycvDRmxWZc6jNXRUe0Pil
mMe054rMSqQj9UhMRymYcqR5VBL0cYceyjEUJi0pwa1yyCPApx34wWRcdhLeu8g3
Wd1a1wKo/5hig5dssJPpuZ6reS0a4NvFK+RLMM7eMNDeHVIdT62MyC40/M8Rh9cL
LARhbm1evCOl1qLc8kgF1yua7ru9oSxTYII8TfQzf2gfpXSzufaONPALpMkdWKlx
av4jjPseICIXnyfKAO4ovpTGN3RPTSiXHme0oFAMUjnGQDrUwC7L3oVr4LtYPlUd
2XS4z4htCtMXiDtP3EKsmDwiXmazaCe8rplaebfIIKMeS4xH7IQMYrYAUImMSVLv
QcrmXaanvENKTSqcDqraW/3akJmazOu/JjxjhQGme2MaqNyBk/FEVPgetI2YkhEG
/JFW2DPNioiHiu/hJTEp45J+aHvd99lShJ8oIoM1bqCLxWgyt5T41MVs/teYXyNq
a8lrDcwjP0x9Gsil53qJJ65YaCoj+ylOHZuPQFjcSNyenFSb1kB76OZ+VDek586b
s9lBKLHCM1sGchFb9F2K8fw+btoujzCgH5nmTx/DLGR+GEsQkylesZEpWaqLrQSK
5w29LgNvzzRf9DKQw9G/iZLtYvsT8blCak+6EDYoshuoorSfKJELRBCNC2h5jxwS
RTysrgp8VUDYuC6X/kMfE66bD2iEA1p9BC9yiuiXQhyvZz0NNex9WJ/BzcZmRy9C
xOjadAccn9AUpmZUp/vS7xxuL+Wa2aMTuA2MsgadRgrdMycVVKwNGcTXyD0YTOWo
kL+QjjyC8VODuV7RJLbzuwKIHzqFvxJaoow0Hz+FPB+QJ+6oiI+zkCZcekdFpGuO
oRlIf5cZjgI+2QMy5ARUaUG7vo0JiAIn0mRpNPqpx5M16VkiL3R0p/RfKxsscIGH
gZvLUYFSpP4eH2M0uSprXJ39jn8flIVaKjH7EMAlmsl/9asy0ULhAPvRjOxfn8H5
sZFlU8mo8Qt+YpbKMww9XUaE0BcCF/c9QaS/Trzdbw8QiDKZ9BLWRe4paPPyUoXN
BSMDsSXkqqi1mfFh/ZxKOgFQK/UDvCrecKqdiYmfyT+d3iHHIp3o2BkYpqYSK3tI
AevgGDcWzL+R/d2zlKyLyv4uJ+g+ZoYnHHqCgfhNn/q9/Y8A3PHhw72lFEVnjX0Q
DD8jlrKiUQTli+pfwem46hqD4ZQvyjOQIeOIhAb7YL3+mxsFa6IpLv91VtgUo0y4
nX+eUYjw5U9AN/FsTrHtpR2BlNQzs2bKt9vzU5bbwNlmr+awiScwnsTcmiQ4Oyzq
ev7U7LCn4GvG3gOPlyoiBcQEHKCb3orczrnk5tjZJF8e3qgzTw21ivgr3LQxMS9J
po2FeEsPR62CASoMHsC5VFsWdBYro8YtqI5nia3QzP+dFDNUMAftwyFFaYr91u2r
9FZ0zad6AIgqI/d6An9zuKJfrMFYiUnhuEQl4zn+WYJfyn/9e0S2ignBTSW15Se3
KG5u3RyVYFxjeNHYVHIYi8aeNCRVL8mn/XaS9aLzqhwuviTNAQmJMIo/K3zmbr43
PexSxwfpbL2VfUmkOr48GxF8DopyTN1F9svp74oGMofvBd5LESMSAKA1RjUxtF/V
xOA6FJMhj1bYeTlIRixvCEW+I17XkqUNy8YF/Ee14T9as5Z2KNxf6O3CbHOMfccP
TsZj88XYgiuyL45gqTcl1IPSBUNY50FJzB9VinnoCzw8BgY6EJXjusb0zgWzPgw8
mAfrd9R6se8K6zvkj8lSDnozYVzhZ3jLPXOl8+4wX9XndhmFUH8pO9lua/9jfalA
0trinEPy3UKXAu9ynyCrcGqxjv0DsQqpJsk+AqlCH+4t1oiCpzih8eb7uIo0tCuO
e4sojfkCcJB9dwAm+5oOYT467KLdlVII8iQDwcGxa/JWG5+HaIEObOcLP/8QaXn+
ldema+MdHbHfBHteTwZqGkHnU4s5y2z7bgD2m/4d55Vf6DYMwZN4cgWZYSF3COYX
dx6rCXwoGByeMiY/L+KQ7ugJXa2NFiGa/29MkahWgtOZqVkYfYW6xtn07FhylP0y
V6upiO4HnStK0JU+d4Cno97PBh7CSbC4vBq9LfRscBd+QM9a6tJldaE7kNoiIcPF
nSBr8XysqrRO0faIZFo8X2SGspLPCLPq4CbIUdzCWka0YqErtzVv6dULoi2vZLbW
rQgM41BxphkNUycNcHnPAJ22VhsPD9froLtMaStQCzl6miJZ6e1UfW5J1FE/Du8W
ZUs3HlJXgjO/jeZu/42uYLxV/jTc8K5b9Mi4N2yvgAM7LZ5Uc7UlTiBc4IKPtrnc
8flwbp+3nfLJYGCZ9cPKAhkuemhgk7TyBEcfUzoFwY2G5IyadtGnEnXtbTMaqnce
vEalgy3lAu1Icn6dGbkWl+DaI6SFDlb7LfG5H7pX+4B5I1HcolQA6NT7eRuQ+M5h
+nqMA7H1vuF7f7M/LVhJwHZ3mMsjoHy0wY2/pxvKMGeB4Lo35yEmbElq/o4uv8qd
0wOUjL31iyVNDb2qe8jqL4rCjlzDDv+xQaKlnEd9rDF2NClNKN1jxASEWq78mLR/
8leg+moOd4aopVY8O6B4qdYU5V5qup3Gh08FJmePjZ8yldyBE63WsBvfdgFnpiLw
F5HRYwwah/KaMc+GNX/dZjsAd/aFx+ReOboTpfwt5qichiU3aoxPPdDyxmIPSdQQ
mf6ntzg/jmWLZRKTd3enN94tUJkquuMkZe9yZfNRk6Xym2ZacrA2hWjfI/cZGjwv
wPL/qdqT2n8EA2no5DV2lSQX43Bzg+1MQgZcP7c6CGUYm9j2mm8ReMn5SAXJzv/b
8teht9BeCdK2oR4S6dd6bTB1tqvicSuZm08P53KcNx5cHfclEweHFeBEcFETo0Wl
aXR5un1MEHNRO5L9t6PErZ6YGy2vxXxEgRfAugvWRkJ153GE/2ibLLOtjDLwXyNj
XfzNFn8N1JzVxU+6wKy64LXGX9JXxFjhswNEVwP81VUPh1fw9Gg5CfLz6QvOfRAJ
p4LEWawDmajfJViwNVv5sK1dC/A5tyxiM1m7i6U/UOxkmm0OEkzugakr4kn8l9pd
yAV1pZU6/L27nbRE7HDjHvMnFNI9H1lP6naWZZrU7HivvhHdOFjTodqw9x6kg2Y1
s4HjFzLkNpuCWBEsaXYwBH/jpTP3oqzVMSh5UW2ZQM35vHGEJ94fBi8OBMQsfaY3
KHk+VvKi382cRdcKVwEZPLkZuz6CpYpT6Y8o3HtPH5wYj/8B5xvIRlVBTo6sffiw
9Y5MhVYBIG2CjuLANYuw6aXPBbasAFI4BRWg4WwUHIquMNQTwRh5kzhJBcNcu4Np
uhtUGaybAaSlZyIR1c3nH9KMAX+iHRhHk9Ip9GrGplHQdp5oXpdZExt+Pog2AH6u
itigtQTSr8ZjbMc6gSPGBG+Zs27SlXHON38yCAX0EZxeZPkOXOJFj/DbgGgb4NOK
ox6qg+/aR5ERWdWG8pbegKiTwKmxDa3nAIByZ4hZbIr0kRaU4fAop/FlpkSHu61Y
9xc9k95JsJxWzhRbdq0bL97xRPNxYwedwPGP4dmk7VHx5R688HoUIRZ7YVQgcx92
zRdIuYvnEghZ8MztofGZXgxHVFfpWTqNvUMb/p8dJvsXU+hTJE5qlDwghyVs/uQW
hWA+KQ8LGcRqnlm5FEifVG1jox9QQcTOAmAjGug5ReK/S4LqVreWv/jn0JhLPe4/
cXFw7k7D0rg/wk9HPchI5LVvvl+n9DPw7mXP00WzitvsOXU4LNLKK1ZejcTsluOk
Cu+AW/eQ6SWNaOLBB/d/aO49pXyUIpeHtDiS01OisHdfLt7vxQtLNzUEXtuoOJSz
mbuurVxApNRMkILRLJ7i59pKJ1iHlJUr8jYeNVVDHd4UNajdnrlUKvB0QzJB5Nzg
JCNBIeIG5aV4Z7YUlmoT5Dnc37UjiHTqZp1YKOABZKIWj41igLNFEYfJyt9wnwUM
pbVcdmUckUVYzwaJ/vtdCFA0TzWhklo11UNIEKiJBbofRIvw+hK9b/qWGbK/XMSF
rfj0Iv85BA07ZbdERpL7+W4CQI6uYvzDghTbhfpGjFNQIbUtZStBxin77zoPemI7
IACW0LQJy6C4XXMM0ehCbK5hCHsTDWUbQWEHaz8RhMet3YWZZmZ4Aqc+Fxi/l7rX
2GIgw1G3cOedAKDzlkt4Py9iHxFaFE5ML43Cx2N+iRPHe4tV2wbjfiZ0CW8/59S+
PrPftKTzhaL4Kat72ipgpd3rWvYpARPtRzrMWYgfqmChZRa33+rORWdmOO2ZtQkl
vdQD5N8mpQj23x76/XlCfN9rqpbwWYugzohIH0h+SiJyeK15K1mUJfstXpoIOGS/
ddYhrMQWeTX0A9MLJc/fz2wa+BOsfsW6QuD61W+U9QFuw5A1iE+u0Jc2hnbhiExD
A0dy3VhnrzBFu7xy0KpN+YU9JDEy4aPyHuuu4EJdaBjvddPXqSIA9E33gPVhUIKI
EXK/jYlxE8dCZ67z0RFmvYWhMyDNaaizZBXpnAS+btSB9iEHwl9nnQd5F/C/jUC5
Q2LRQRrZYayl7WzfC+yMe262Qo/usY0AzIbE78rqsEyTHrZx95qdNmi4WUKTVyQw
muk/l6yXpbU1yYqtl4yZwi8R4tAVzp26i6tyWsCcHT8h5ieqBDKsje5Uu4/gTPpT
E3KsTL5YLgq5X8WgN5RI3+gufCeFXcyDRnc0h5fn8bS2weHxrZQBhyrB9rG3CtZL
V+i4LHHa3O3QgKU16KQoPzzOH6eb23iZWxbYD22YcN31T7Ef8v10AhAHZzH2M3rs
X7CQ4OJdgtLcOCDb1TD7JgYqN0BbHx8l5myqWzXzjBGH11AaMrpUYAR0B8WJZObx
V7yXD7gaPV2bN72CMk4JNZacTCsoxa9IHLXzMpVJrFv22wBLgUEMrYLogoCOj375
bmW57H1fRk5l2IEdj5AbdjVOsT05tIYDCw5Dgkd8WEDBXJhbhWDdv+s0ljSctPWw
glL4EYwywHYtwcGcXLZBuovyeDN+CHS5TAuoqbYQrJQsMftnCN63yVfAZLm6FBF9
8P/dhVN7uXpkgtAHn1lBHzB1ltYzdPRSulED1EThGZPxW37x2bPZNaoS7o4+ZI7S
CIQe3uoM6HiwiomCrgUqwdiqS0vf66zPDYwsyZioQ8s+zImq7yMet3mLAhfvDH3G
G3lesAvElHeQqdw/VqeJrqnc0CCNdzDW0x1/ESQ2WC7HL3A9ddCv2daeOcXC0euw
XlqHsKDlpruYosBMZgFyHakK+fZiTeNSpffKB4GYfyg9QA21JIoDCaRAG+dD7uDK
AVzhw67stc5RZ7mQelp1iPfipSjg7iTEBfY4z1UgNoYgm3FUzp3eTJ8IRwiPhgSL
o1AnOaCZ+633RZrhP/9NxHw0r/vS/yI8kw9XFqiVJ7Iw6CjDBADHJZvYzjW8avV7
duTvOQ/g6hUxkta/NZOJefsMr+FWhzA+DwRIqeCM44P33Gx14f4QGiFNZWdwscH1
AO0WJfkBX6sIA3kIn1zT3W2vVEVTj6UYADOCv13e/49jhaqiRwBZOYuTJge3kQRX
ohovDvilYNYbky/Vk3cdeteEMp4V61TcKv00c7YyO30LJDuSeXtjm1IoH7sj1/0u
3BQH+Hv5sy0tZmloCeayF0FlU0pgRMj2f4z1TZKdUy8sSWqIf1DbKNWQ+x3J19MC
+K0qInEtGvAhQPLouYMGkAQH6Ck2ejeMmSyWW+0Lk5SCx2yDZ3eMOXiBkXE3lYEZ
rcV5qKSvHHov4iZdQLM2d2PFwrA+JuB+nTWxAjzKOkdoEtFHM3XK4BMdNhfEqaoi
BTB6poIylNCIUEvdOO80Fft9DYqFtACDFkR8PRaQxJuHu00MUevaqhnKxXEOzciw
dFxxOBAzltkg8kSQPi9KPQBsyzwBIBw3Z/CviHgG2D0kXb9ZNUkVch1LFI25nwhi
uFlWft9F4p98q52/oAYA1D3HelXUTeZUyxzh/fjD43yrActZEMa2HqDOvVLTGPjH
SmuFOUOOv3mziOhndW4qYX/ohu5eNC5+0OLq1irxIawxLWS5LsieQPZTC/OWVRqg
+pgnsCcVa9kzC44F/j9OjMbsgKRCAZE+Vxrb4j0HE9XUDFMhIbDTHtir6E0mBqVB
DYvGSKj4c+4l5pi840KOBre5HNV/4tNGOGdaqXtuXvKKhUy3wftiaayws/wr27wG
GDiiS7fahmHqNpweCsMu/lFFFWRjcg7FPBY13kEiS0MczCsiR644Vl6avWTYdcNU
ANjar/G2i6JmDb6oUFff9T/WnoDqqpLI2hxJoZACBFSRvnClAg03oz2P99EV7aS1
zfaE40OBx5BeC2pef0akhmONJZGlTkSvv7tDQtUwqR83nWA7Uv+uXqLw7k3HmPgr
il5YSJXyfk0EQW2VCVxTvqTO/lT1ZJzfXrK1icAk3kyuevDJ5dz/42cUaFP/K7T8
wc+pCC6im8LYpbeTqsjeV8ss39YnBKMnx0SOyN6VzQsbuuNa/wohW5xYsY7XeJvr
bLReLio1VLwNUEiEVASIGAlTQxqSmhzpxvDz9e4T9ZqVT6XSz/OpPGbTLjEQGwHo
aoK5F/mEDTxl1RGKrzZeJBA2EAF/Do+1eNDf2fSDOw4wnk+yAfGCi6uW1hCVxUxQ
HNl02NDFPIdDMzvuAW+A55yK30ixau15Q+UWnYRe+bOIO04rTv96e6ZVDJax5zaz
rfT+A4xZhbP/3DHj4RqwwvJwDJN6w8h1kWskO8Q/Jj14wyu/Wwi6c3aCAHDemQz0
B3FeR+l0Gjp+V7zLIN1xgVnNjavyMO3iGxplcanpqa3Yst1ZFsUUvFSEhcYeqxI6
xLIPxa+5L8LSMLdDZVpAkUIKRZVlKDGtM4Pq2PxaMh9gx4jNayZYl1GyvvjR2RL6
FvJ1+c6KUNO7m0GE4ah6U2Pyb62DzLWdsP2UTLbwAynNRQkKzzgLm2tDbM7o63ra
SCF6RmVuHy2CCWnpfLNj4qxxSQOaIylq/LaWdwNE+XL3eYmCuJYNfkiLWAXcVk5t
dfvjxG03kuAsJTwHGWS58xIp6tADJDP3Ac0SF4IPg4Y+qzS3rCEfqYgx8Nf96M+u
4xnlU8W0UwI6AGJzf06CXirxLE5EiuJvNOwHhUuMuvJslvNtDOeWPsC4nx0bCoH7
yHcMatBTbCGIKcNFILTTb/upQHxtFefkJaqzogcx7i9lsIjhiyBqRLOHQy52RNWF
V9aRPt/JLTcfsYyN5rYn408/94bwghQG2zKziAtB9fRl2KReMWrRuPfOesr8ZDPi
8QUFyOOhJOf3/0ZjUxN2Qn+7dJrF5XtbbE7kDwKOAeEfs8ZhKeHmSejPPQ0qB+Dy
RnHmIQKS3iaJpdWTRTb/dEd7bs83zXHAeXIr3U/FFwsNvx88RhCR2tLHTjDurcEK
QkAvCJAa3tITNP1pLHdJ0GOgZE65cbBzBsHrVKV73SxQxFNzViE6Uf4uIdosdGO5
jceN6r6w4Z+MERnLxjzdGU10zTlW00AR9krhk06u3URfRiSWqw0f0BoIL+G5XV68
9qdZ3Ls6qnltwaWEziJzVn+5QOBwU7b0KwNRpNDT5tbnLdg9g7+26A7bXZzmXbfi
ISBHBr6tdi7wcfU3BX7CiDt+ndB6zKo81IdGk74IA6bCFUtoI6bDNgGpeOH6Fe2Q
VX8AdyRIqOx71ZB143y7/W2w2kkY/wU2R2SnJXgTiMCZ2obwBNkCdsrqokumGgb0
VGaMo28L2GJ/4aYSDQBYgaA7adIcrVr0ZsBBR9j4e6d6hBHc0Y15gyLqvlO3y69Y
Uy3EpaOLfhsrBhn+/Bk0MYiq0MKhK+FsFYDJJmzfpwARt0bVgEWhec9UPz5Q5eid
RwMGiVj1R9Z0sKUc2yyzvGXewwI7mAr8DPxuDXGwjmuIZ2WfiJuUB3DEULmHnDRP
ruQ0qSwfduH0NoEEiHd0izFct1bDrEs6XceYva4X5vCwGhkqte2LwordSpKcGHAo
Dk1lgysfw+r4cxit/c0ClAdFm2lFVcI/uawE8swTpffhbKDIwpl28t/G2RQhnH4Y
+0OHDSbdCLg5AUl1itKKjjGUH3WFW4T4pdKjGh1GoTKFwKNxtm4vI8r7xHXX4zo8
5e0TJ0mNitP1qriXY5zQVzOiftQSwUC7YdDlINakarC1aLZfjrZDKsuHajbiQB/N
DGuVRc4WFEu+ZM/s03+bHGo/2igZ3uJb8FWHjFubVee3d/MX32UWP3Yeq7LXvHKX
yB7GG9RoUJpU+vPDaSOvlnrAQfyb7R4lYPL5ZV7RfJ9yauizofoIyv3VQF2TqwD8
gdv5mOhjB7j63whQCxdlp+aEtdj1Cs+qRxCHryEcXjQeNTDuakzvefAlwuLY5GxB
PDYLRqHRkKycyu06jrZG231pUMKIb2Zm8b0bNNXhZ6Q9pyYAfeIpDCb57iPpm3JV
KpGsWJHf9llnRwgwAlg7ISIlkPSrz6wrBV5UXsQH9E8wmRE0FsjrEToUw1lCMp4y
gj/m+TrqMNr5YkxXK5ympOazQ1Lc3414CAiY+kD+NgPcPigITSq0ZrJZ9WT22++z
qOK1LpQNV219KqiQOHLnnOegUab9edKJ61QGIXv36E4zKqhqb4YhlzDvXzkuEBJO
bYjGzasJDatEhHUlom+dMqw1TfqGY8vwNzuOXJEXNWzonWiUJHlC7O5cbVVGd4JY
Po1ZzQ9BCl9z7zBK/Y+VZMBfFwopHmyLrus0biPVyQFE08OYHRnbo+pibKZMIdzp
pgdvbVLF+m8hZo2NOWnor+PZ5tiDVsghuOFFV38paLZmvBMnVYM3Dc5oQKR4EKK3
U4szQzsfQxmzEwxc+ZrcXt/GM/kq3TJEoeZgvzGemeP2Zo3cX3ddGYsOVSmHIXeV
d8ou/JUoyfbLe/CbcntTSSN0yM+O+nUJ2LT39E47BZ5uZLSbEVQGmOMOeIYqeP48
BxQT8f11nRjQs2PopNo1A0Y1IjQY6EWzw0QKrNSPVn4ywOeLBzW/jbgqcTqwevnh
BCHFoJcAbhKGHYP+qtcPfcJ6FwdTBaH3QNCBuKYlwStxEODTk2c560sXvFMYKiiZ
RwMi7orLiPWXr56II/qzvbvyfeS2jdTFPkINNrYGPrWq3mNIXUvUE3QxVS3tPilL
q1Y1HTgw9d1l3hPltCLrcMtf0tFxI/c9K7kE7dVOeheUGDgs5Q1kqdq4mjnegBWZ
cKkn9ed2CAYIbJZl9nsPpR2bt3KpXOdM8AugpCVmy+K4iUBeCOacIxX9xJVFB3fQ
jBwR0bBM3ulDaCa7W2VY+f17yqiwoL+JmJsIePrgshxFiLxwPQq8OLzhw8gQT3xC
qqGO519w2a9Q4pHMavogN0MnM14j4oeymUSKu7bJTqWEbZU8SXoI1tdXGB9mrZkA
kAJkFRHOrOOPnDmPDqAPsS7Y1cz5CAQZR8CGSlVw0Zd49zJlbXjTzx20izgC5E6W
tNeyiSz2Fdc5ObefK6VkNRHt/KRz0+2AtPthGmi0Vm99y8cX5fIm1ibKrIc3a2F3
R55jHeb/y18fHY/VEaUwBoB8JGbm2/E9ySqit18HnbMn585cu4JOtBK6i1pO4CUD
SoeprL6lo7xPZPG1D/lQnlFqbpY77YJdEJUNsfQqXwvJ/hz16nwdCipxyl1zmeUo
QyAT4dgwU4wMzkwTdYnNcgH6WuFZH3dj09vSIbky1q4TDtwax3SeqxR3y1FKLOEP
xSxhC/XcN/lv9QpmA8ZHZmirDrn1v4e/CZCGtc5a3QMrnjYGO14dWYHbNu2mn17p
4qqzkbcpc4LTzDFSyglAy/RPfDU9hqBQR0a2V4XvSi0AjXYbWC8zplx0u/QbsQb0
6VDRdt9GOJuBG3CQASZ5ZbDQfMXT1uNLfEhAQ+khdKNLkO8hnYkQfsf+upyC/Keu
vv7ZqnOO3KStcjOo4uJnAfX+PMrThoiQom/Xc0mxhd7sIMiATeMRvI8jdZ8+BnOS
Qj21tGzgv3QX2QZ7tuwymndu9EsXbdfg+vzGM3QEGJHI9cY+SYU2TwuEJtSfD9gP
nQkSv+06/h95uW4q7SEU+Fv2iQLiOebNBIh2i/DaO64aQ3x9Ol9aVI9chPIKU3z3
WHzWkSx3A20FzT0crdEkc88C3GN8fAPLfG3I7CIEnVh8kCwpuGsmMG9i7B+33PqI
LSuP0cVXL0cOfhhSOrg2j4uXyFmtfdSratUy1aRt3Ljh0cECvoWnt28QDjkkTNy+
DaLtIG5ZUt8/9457oonqxRiHCDOVV6pnl25HLSYFtxLrQ9hd/wuC3asx4nacxrCs
A5kA5IlOeSqFzj3Eagy0aTGLkxMyXzZBKfu/Gl43V+flcDATonql7q4yUxsMs66L
aMHRkFVnk4iYIRrWoPTmopr+xphuiKhNFr2DH/AHRRL1oBP7J1Tt92kkptsZ9bWO
PT+Sx06a8BAwBo8T7wsycHEGJa6z2CMzDqLkgSIzOAiiTyXbVZoVCGB584uK/4Is
ySVaGCJBMDx4JrZa2SO79pfsWoiKH56lOossuWxDm20xeoMSnmA60dxiext04ZhY
OjFEWm1dIumkjonA7YnoBjoAxrRS21tRr56KuJ9yUwohMjebKHux8tYACeiBaSyc
/mxXQKrIucavp2/fCKi6PiyqZTyFHQpEEtlwaC1rP5hwxmAGiUqV6ZqeqHBVac1Q
TegfXnq2KWa2zaOAoclXxXCbEk3JC6WC2dupPo+TZqb4bIsV3Xug6LF4GnARVnXo
HUBzwb1IE8iad7wBaYDw6+e2mx4TPdZ9cEZk4SMXXpKY8LJMwuAIXivzjmbkAfdK
mcUfziRH1rNh2X4SKf0SWPjdoSW8olcreEE0W+aQr3elariCc1MKUuhVmOyXEQl0
XwO0tzcUsr2kWdjAr3ha44b8GrxZj4RSPq6ExFBA5D2Q629gVOEo7UXzdPCUo7J8
YcOGbDysxtBlBZqGuknW21lj4s5nhYQD6q99uIY657pnje9YNryyM2CzmwNSggmu
Hgn551tdsSi4od4vDCnSuG/+uJ4bN3fjMkfwN0xgXk8wHhibxniQ0Imh0wTdNSTt
P/WalDBQgkoS29blanxlsMaEgWEKHfXiq+mYpPvUHqSzpMMAgjUQ6jceM3+3dqfO
fGFfHvxxdqfXXXow9HtSZVy0VmCprbaPADfNlkeDyWZXHfJtlOfKgxh4tr+66jw8
y4toy0xbx5ojs1PIaA6tUvFPJ0gQAvCkATPcYYn8/TJn0AfPsBCP2X7eBUUA6VWT
4sU46yyUESoJ/6yuU1aPCYX1qWqSbuC4cxN6s8D3jVrF1nuKBA8jHYvTQBb3NwKM
fBAGA9ovoxAliWA3ByvSIOKPxrGXmRaY5/GuIyI3By30I2de+rY6KpOWeflNkhOX
nL0cZMliEIJwKCGHLW1JXMPHjwOUevb/u9XXZLslwRUemXUk+60D1idWmDtcnfPi
uNFi3sSdKSkhD3IitNp0OTIjclApB1lTzaga1j1DvfzS1nXKH0YcwR/BvzQN247C
LaMNKVxQOFMxxge7gixN5+30e5Ki83Z1OdD4ddATBYOtPBvJkWjCpYncwnNRdBtD
XNo5fM2s9wH1r+eCnrltkjU+/MgTDLXOMXBZK2MF3LmF62g6PJy4aw5izrbL+gn3
/PEpobm2FzFJcmt4BLdgUjRYDNxqLsHY8k3bxONL6hUKpJZmCT0qFp2PbMLakvYs
4Nfp6eibtuJmmbkX35iUArT/wA9M4XWi8/hvWrfrpn9fZWe+p7jjpjduzJqlPpkq
IGzcZuNO6zObqISgk1d/PGnOfJOFWMDfB4Zx8tiu4++wnVQLtVma8Tm0l+BXwi7s
B8C91+nlBQCbjGL/g8pscudH4dK8mSiKgtj9172bgydhsNF83bPOvbVwKbom+mi3
7r1hkX7x0DDVSmaqseBFzZQjnnDrkJyRDkuGig/Oix3UFl3rKz0y5lXVkGGv5RR6
CgItjoAKRyO22EFj7OOF4VmkTSKlEb9x4UJHHoDXUdqzszp24ImXNYSsQrX081Af
pcwLD5aDFM+x2k5lu+5ULV4lVaqe275Y3PA+y2SDQxQt13jzzcm1lq6h9YLH8R/h
J2al2jdTIaCwaO1IQuXfHE7UJdaTNyCz+xZ5zYm7XiDoN5pZmrL8e+4Tj/OpkBBH
XlM7lEQqAotMV7IwtVvvask9p0PJb5im4w5u2y2M9w3sMx2XLsayvjtiaCtOdIjl
hKixyzO66qEU+oZtQkHIyBtieuNV3XRNWEFJcuTm7+mtqVPpVzMedwbNzcYxiIGC
MZO4p5F58K4OBeA+qKEpgXN/7Hj+s2tNH2x5/VSabcwym7CT01zpRkBT5DlmMdwt
7BpxQNUUxa4io+LkT6MbJQBqruJZq9nCtUIK6SUu++6+MKOKDwNTKlIIe+O90Qfl
rwhtpBqSL6CtKfqGjbYW2msUCnqACiAa1aRI6R910OcSZXY2SvoAl/Tvi1XWaDyJ
COPGr64WT+X35lflQ997R/OQSsxW3hDJ/QSNQIQ8BSAbOGlQTILgM70OBJlArgCZ
O5eMVEFALH621Iz3uvAq2kfyLeoDuLDqeVYP9ST+eRz1lQhWaz+t2iIjP9Kez5r1
C2MN+SaBQS8q/JPLX8WE9oYgyePOPO/B5zmhsE88nffWwFrrF+TIjt5ktKWgsD8W
BQWeqSO/D2kl9tJzdQqvNXJ2QqCIPic5mVq9p3rzo+bkjrx6dc1VNoiQd3WNM49p
n1IW3MR48n6EYGmj7tsl2FtIicEZaTxxzxxPfslWQyvEUeo8bqZLxVf8rpafrO7C
gaaotLZwj1S+Ab8AlxxuLx8hpmFGTTmXFkDh8wm41GNOzmF2ukMMzyWzVQbiQnTn
P5hQJuaKnttJRcTWEHf8s8/A0ho4RRs94ugO39eQg4RO9Gj4seITDTQ4b/Usm2n8
Z3e+hTFCuie2jZx1Vr8ziBN+s5G7/ld5U47WK0kXQ0x8ndO+g5KdqhiCyVZky3el
6OB1D+iW2yOlQzN9xy/Kd04+hy22cmdWy++70XwCnSFUlOzGTjmKIkLi16pxmG+8
LukikmgCDRnmyPyby3AfcWQBt3nGr3yJg1jMGKHEfQBne2GSI8kpoHKd9Cd4mU05
CyMJ66kofj5dJE0dnItKnVPUCeZUyzyrqFjlIzVa21bpVZXInaKq52Hds+fgtXAx
nV/q6n5w7EyIZwj6jSbT+vg9lP+7s9HDlvFdXcOc5HWAz8H1H744Te9/E7T5yXGo
JT9Mv7+dLPgi5ST0gfMMMCa8PsFzNZvSVWw+O09FkV2ghk2NjoPYmtXK4cHhuqrp
ekKG7zQjkydUN4VLW3Dqfoy5cABUSSKuoADRi+jaI6IlSZ3LPkfwk9YLXT9mDhRU
qcRhnuEgR5tQGB9Yt6JsqyBIqmONXTklHtD3OsJRE4fCPDNjR2pCjrZwfqOuSxn9
B/LOtQucPvy3gEGLDjnhSoiz4ZkBMWOjpCibAep5BC+QUTmu2fG9ofR9DUdD4M7V
SSpxdmM+9aymSL4v8Nm/B+udmA4hM87aXbBI5WgwjqrwV/RQB8DqRcTcHmrCWHZw
GK7ToemgbODt6MP66NJpDo8IpxWpWno/NrgeEK40qhegcloAX9g4PsaQ2egKFDCP
a9NWFXKkv1NjHWlyu5eRDxwHqj1JfxiuOz1nSekkyh+vmtAuHsuAFTBAIemfKyhn
RKuId+RKV2RGx3cmS+3j7wr6IBlo5fqWOvnZFUsBE91OhGuvJQHB3y6Jp0xzzfTp
nfAZzAYb2UmMEEPifdRJOxAVpMEwhjBJzG6rYSl+17l6bFVhvvhBaAYoWFpqLFRK
Yh39Ec4EVj5MK86ofXh5jdNMoqkNedIcMp3Av6KF3W89UcGsRJsABT6omv8PByVq
KkImYIBbRRHIAW/UONWaAdBzf8FfwOvixmmnnQIS+U3g2qjJ4YZx6h1XF5bwqyYf
uCOh42VBC1vMXRLsxbRWRH4uoQx4ObgWsvFjlxy6t5LjRIpBHfhZH92ccSlRTHtH
D8pEI1AU+4HlNddzIDXQvYyKkpipERTXY0baJk8uNHAwr3beQct8iHWQpKMmYAEN
WQkYmlcbXaYjq7RLYOwEzc0ydqDav0JeKl0C/c7VgAMdLuwqV6FfzE7zDm+OrWZf
96aMRnRAh1mW4fHIYoxpvce1TfkgZeifzf10nVgcNvzFObHozRBZvSfAM+Gj/xQA
07b5HMk6ntxes6x/9S1FAbNZLiUKBnS5wf6CTol3S/H/vTs8jnb9uW831GXEmap3
cowAbqu89htoWX5W81MmGqh0qZnyHYOo8THgGfxfw3YOhVPO/h/M4CtkrHszfYnd
q/2aW+u8Jft0U1IVhWyaluq94sEJYfss6pIjF2dhMOwHZKHgc0g+TSkyOFYoqEQB
WumQaPnTB3jMZ+LesDfYdWnPr3NHoEBAt6ksqDwDmijDBZEnimCt4nKAX6M/3M6D
5fZXnUjbOHgiWraPsnRd8cZGXMk80ieuXncy1JlIhCaxAhcBP+nyJy3MpJj2dy/f
iekycSaa5bAuRvpRQ7kJ9PwrvZ7Fc4ySStMM0DTqM4ZGWyLERlpGhw6xechj6Jra
4NDbzfkNLQza0G7kYIfoCFC4MC+plvca345OCWP74m2fB+ht8WnxyU9DJ3qt99qW
gQNh+xbIo3ekmYw54U45N+Yk1lv5CBZjpmsbSg9X4SvMKTAKU9SDGUJjL++0nIrC
SAT6p3ZoSDbUfaIYmA3Fk2/TesNgFt78XkUA63OCCAjyCV8/KeguWftlc2L0vRFo
Ta3Vz/9qzxTJzw6GuFe3AdR7d9BTaBFcwImE3ac8QprD3TWibMsdfrIaYqfb4O1o
qHXIsrAU+5iFy92b6SlWvXmxZcRI5WQX6ieQ8oWsV0/5dPsmNPP5tViBWTqrZp8b
W8Y549kJrAY+1+GFD2NMKfvMq0Nh/v9s232NSdQQ/A6m/leNT9Of+CH+8iH13G5f
U0oLjYsk07TVol4l/2B0KZ3mXFeQ+MBCdKnIQdQb/PBaXZhNlh6RzRD2DY5yMZPM
nt9GKIEWPez1bJbWbb0ygiAPlXl9uRNycz7TMsjGU+o2dZjm1Jl5t6vcktUhw+vY
acFEronPUEGq0Zjbi2TwDzjWXmqUKoOLpcdWA+ikJnN1OLNmR+W0AoplSSYp2Piw
7uPOlIokCOqsgK/9IyeGW7GB28zsJ8eyZpB2gatC/xSYBGJ2lhqFnOTclm4mOvmu
RXTWARiKGRUbvg8atrLiDrvK59gmPBsfGY3/74wArv1Ny2H7KLkJmhS/TZY4qTIR
pplQvy9Fr/xp2PMXqt8BzqXQroW0/d+w+2ljIvsdX9gshMqwzbaYSpKDo7rp5G8t
RmAwosJJfkKqCuddxIy3242o7NtHZbnu/YKk9jqNKIZ4xy0heuxrg+HS+2ydK67j
9FRGySIohJVke/hC2TlQxwTIH1s2oentTWDy0SFgrx0oFCGL7+TUVyHxZzp0rP5q
/PmZYHnQQXr7zCdYBjrjqqf62sPloB9GhplPNl4m0fihjh4YvuXaWbosr21MIZGb
x13aWWbUdtcSUYgyo1aUktaqVCc6vrcs1lCE2WnRJT85Peh0eyyCSZ27jO2sJ+Rq
H4VDYCWpPIDn30P8WnaguqNU7UtwbyTKH673wJwR6zXMGwo2gDgV5DR21Z9GzdY5
uEZdNYuJzwOlRUSQ0znAjFF9G/hXMQLt4FS66HnKj5eaAgqjcdOk/Wm/z/enGG/c
PNbDD85FFRHdEgqd8WGfunIf5wyMpjYJcXoVRNT2vjb2WXG81RSJ25sYNLf/tmCn
jLbU2niJl5keM4PQt7cFWtvdOYqUWyEUXaYYbf2wPT+NgqbO0dxOoVeKnjUBo2Dt
Olijkb/BpKBwXrQoZShQSqfE7DAP6LBoUUy8ygTKD3on2FRRSuNQh/SIYGU1ZqEW
+Rp8Iba0euA6i8uH4K9ZHLeSM+uZbjExBI/EIc1GH5zw5KzeqjarD46aYnxUjAXz
3e0Q1itpvEZj/escHAuAQquAwvJiU7r+LjI/o4LlGN4EwppieMhkrc4vI7+QdRWE
xhiYZ6MzfpJ+7in6kRo+lwHcbAAYthXD2mfBPQ/2yHX2tls4yEaQ4oglTFaFpt7P
GghJLOKZWS0hUkzBm8uSHw0aiqCkopHhSqfo7G3QiSnbJJcEuj2k7CW1kyFaoT9I
xFvM5582ZB6VgjJnUwTontK5Q36mlPrRpIDX5GPk/Q6RfaUqxbT/5jzOst6T/qa2
kpCgf6wzWvp7uDBEXaLCgpVibZH9hFVauhNsLAIbM1uJozXMkwzA9WCptg101qtZ
UYmB/6yW+iVh6hzihhMTQavhfoW4/8NYjxzLdniHvF2dEKu8vqbJyDjFQPRlyPts
woRA/sX5/BTtbOcDCkJcJgVTGqrKSdlFgPVyVmDM1la/6Gu6BOA9TEjl+SSA41mM
e0QrN+cCupAQGORvVgsKX0dyndsYwG05k/aXEQ8D7SWEER5blaM56/dD7vw5C0K4
Qqvmq/WzfiBSmgkEITbqYfP8ZZQha3J2/GY1T0nTnTRvuUE1RWIaHd8B2+Op7YNx
2yCbuh8Duw+PDL3a3jsmbilL/y+SRU8HVY3xwMSaSyGofNhcr0g+JBxGkvhOB0WC
lF2nhiLqMKPFSB6xgqumtDUbCs/+DH2Q+7lRwdwHaS8g/qMw7zdgTemvjt7d5GEF
WcXZEjRtU1UGohDqxdDDxtO881W6cakOovJ0YJkPlsDt8uGxAc2dRkBoFkVmF2Ki
GcfpiyQm00l06b+19PIy7LR4MQ8Jt9aZIeFh0eDUXCgf5QeJozCZuymVZ7I3xdOy
YnMHrhHZZk9IobUyQyfpi9Z0Hw7gbQVXLRoAQWjg4/pulskJEoD4QkJqqkGjGfy2
LNNsUmSc25nOAFKwMlvfPSh8eADTlmN/2JyPEPemZ4Fj2S2lJI7Da4n3/EzGc8Bo
cBfRLFwMW6apJiA4rvKuxFGwmgq+RFrUxRnsOz50+3KNOtWllvxJXco9f8ska/T2
Djrb5wFbxffc79iO9WTkl5QMSVTKIFJ41wiOuI71eWu9jfg8A5THU7zR80LAeH9c
zV7WbJkMWXCZQ3n+B46bdr5D37kkDmEWX3j8uz7f872JRN2B2/4ZH/z/gA4R12ug
FouWDg/TgYXSOUcR70DxjnK8Vq/m4BEe5GNhl8jXDlXfHDhWpMAfFu6oQA+QVlYu
2zJydHv6b/zOI7l2Z+uaOIdtDOf2hMdHxPk1Tdx6rITM7SHl+Bbc+6JUnzo+uFxM
3NXAtm51oA/fSqNslZMF2cVTHVVgL77LjAHABnSHPwKvZe1YDMke7bGv4T6cvRd7
HWjrQFOtvCuudIv4JIFrQGOqv+NF3w9eWYqpJp/3JUkX1a2FkCrVodMQDh6V+3S9
Cy+DrUJGnV7ELn6UxuuUViQSLQxyiWvhoMVC4VCUPSY+ECx4OP+IgrW+Aif1dj5t
/yJM1xlj9Ye7ZtOv17bWp0M8pM2JPyINakZGrnBF50YOgz1mikmheDRoQ43PEvUC
beCWiEv2Qsa5Nr8VnCYHyv23vJrAK0fptZ3Uhf+QA+HTSpABojFCJJWHLKlFQPUF
EncdbCwgU8kH3s7DQgi/FT5tLxMYgusvsWrs9kyPFmqGfCNqkRtI/BnIUnYRes5E
uVbIezxTX4lk/61TTfznGRGOhBW1YZ59KaUXvnIsMq2V6BfjzX9CXnjsFXc1+VKE
tR36nQ5RF0W0MtfsH9py9BGtzHINpNtSj3kL1T4xbItvK0fJ8k1HdM5InGL9OCLZ
FkI0zQ5mh0WMFwnDhqug8A9sJN+WbpzpirVJDmPIbGM1NA+GlprT281W1bruYv7g
a2os3hcIbDpfkph5JD7nEBdhjMWB2UQvNNfdX7iT4I5IAcVXlgfby0vTTfT3GPUN
5Seq2vSpkFABGGK+pBEsal5LrpCg7rL5CP2SknqN3xAuYTcQR0YDHvCn8heC9S2W
u9UwriCEi41ObcHHwXP2ndnit42MPUTUiBE5KKaTBQawmbjOL14IGQtLDl5BIl17
aSyon/quyTnymKoXyaKTtLR6mGQ3ZMowjjaxHD96lOrZU/Nkiwa0rDMStSK1SSJ/
37UWVEA5ujjiepNsD8tRgjsYQZj8FRcbe9OkS0J0ngGIwhrwakudNk0a82lupiAn
mncKofCkPO7wBEb4uvc/WJ24ME2Cp9VejiRF8I1B0TG5WoJcacTCHz/rHrpeedTE
mL7nm/z0jo8lW/h8txdh47FhyOQoZqJGwlKP6uWuVBOGEfyEtdZz/j/tkbKG1UF/
ty6E/w+eZnzIZkUhaZoOHgwd5nhzDTxfmYuLmPsIc4zOaXfyyhr1mk6Rdj7MC1gw
/5mCBo8x++36x86pty3MzmZfssAKPv6VxhZEVjPYu1YKyxQMxr69XcOKp8yslXDI
rGXxX5rDnLqRiQZ940pHEv827AwLPzbrKaDhe1DbVjf73WIZyJQBjxGRSBAORBRq
FSM7WnIwXtIzDgEeQhgVDOaVDVUva38dDujeBabxhrMo2nncyoHzaEer3PhAGaN2
CSIr0OXQvbVsX0DBTmpCjBJ+SAdSJk9SODMsU7nc7IK6R6FTTiU9W8/pxG1k5ydn
JNvploMVAVG8ONdv/XMT34C34Ux1d+vuPB9psVLH/wsh+CcBI5Mmh1VYQnzjO/sb
v9efB11JaEHBqplF86lRvgXBWmPZR6nUNS3DtdnMC+XaiUYJjOXSApI4DqPwI/J3
kQ5Vb/F7RN+FJly1s+97prGndj1lZTn6bpaFBLn6kix2kKiWGKTL0rZixP13W3Vd
aptl2oBu2YzrXMtfTQTP9k8Eab3FcpaUFj1ZkweBjUw+zaOaYFAkVqYJL6Tl28oC
G913DGJJvRwChdKbqLcYLAJjSLoNc4JpdhXiBhYRt0YZ/dCVNnR/O6iPiG4gZVFd
Pk8e1XMkjYCyLDQxW81x/AGJ8Xj800N9pcvSvL4PcPgGbeVCCQo5/mXgT/+AtxaY
K/uiF1i4N9Fd7dY8YFqfThEQwY4rC6Ar7sXm9RnlK7BGQBp4pXQyaxU2y75sI34E
aDemAsEE9jdP72/L5sts3NLUQWH6n6xajxBQn9mg+Pd/jYAMjWV1uED8C1/8K4lS
E2RznIzYpIAr6ySHL16gVTZcf2HRUYfkQ3k/dykDNvRwTCdP0pEJi19mIWRcha4I
1uj7ZxZdMTilyHtCj164Mt2tOJwMTEVijywiUOkT2ezfX+nMUFofhksCwghORYqt
QNhtGD1efVpG/2GkAZ3z4vygkepeA8E2jFK2+ftSDgO/O5uAhApa8LrWyXaL8le/
ZyOWR34QLNh7wYbhPL7oXoANpLawfXEBSe1eejJ71crD1xj4pSqWgurXzdHHCozG
dRZIr/nDcE40AL8UUjUVPEqq3LlQE0bI8RVBLCpFSw5fDnEYtvlOsdgzRfdN6NCC
nuRod0P89RPK0gUOIdHZ2w9g84ZArjotDqatNyKjDCaREizyplOpy8+BzlkXla/2
6uDNNzBffp7gS0PfkEJB0k1dixvG20WRxA7mbmfHX+nwwpiz4VhVIE53T8srhbsM
3laRyz/kfm7G2uLS2v+gVvLrAuk91skUk9GbX2JlwhoXqD5dPyE+N0xLBZK3va9Z
n9KR2wcXFdn6SlxC9znmvCMj/kXZp5tLMfXMsrH5/cJoxCP1TqTzIgxQiKawtVNm
TlWA6IAQDcE8Gt2xlfr92n1AkMny0UfIhsAkurtHLqOKrLt0rOqCCj6YCqM8iRjr
5an8yKz6FXS7rz1sCyycN89aA+QEKYUBPg3mmD/BUDmGcFld3jRB72vjAUaHG4Is
hgwnBPI+zOS882sN1I2TaNYaKpOWcEHAMDlS+GBXnYwA0qTMqBluRVtPJDw8EMY1
Bo+bXbesxtyLOrtrB/jJrZj7u92jCtFAjw3lTF1zdCMnghtOTnguFePBq5WNj+OC
tEc9BP4eQIppE/0ukmbMWMLImq+GnzT4A7rG7nzv7Q7Mn84ZydWiMderrQMEGZAq
GDaoSvm+AjLkeSEUJvB6GLpWdmWs7Z8Ghr6LU9u/ObRsocFxKNxWz0tZq1q5mswG
YiguUmzpe20amosMKRwb5A8/6rs42c3hVgr/jtxTX7MAkdl42ATrolw/OHCqyMLK
6YNPWysxiEdQsMvW2f3nfMtEf8ZUply5WgSEGkTl/cx3WP1GfeFXMge+IO5+52T5
r8P6yuqioPfqlRa0+iZZrJYHzkAewaedyxR8ZLNhvcLN61L1EtyctYMOneuDie/n
kB7GvTI9UDTWritg6e0LLLhfjnl8h5uXPYIAX3XrUA/s3bVAGTxPtwDmLgHUlC4A
4RLoQ0XLge9/SCExNCF1mWlIJa5byW8eyDJb4qNAokCb7mpJJxihTbuTe/yNQ8Jr
wacs43huWnahcSdqWtlXu3lRBXmEsZngruZbDCyNng7H9UjsSiF50HmEEGJYajCF
IUxdkBVXVm/V79NOdfuteRJXp1vxzSND5+M2iTpjGVOdi8nH9sCeaaum6gOVJ14p
76n/zi6tUXgHIF3X9xlSX7e7syLv6HNXJ9jtVkU3wLPtrA3O86UKbEw4LAIYScsZ
dkLf7p5ofiItTk8oJFG5tc3M4mUts69EuywMlss+TONFiiYmF0J+hNzKZ3dFY82z
qBUpgxLiAflNBuG77FRlcyEEXpw5c9xqLivcmpHfy+Bupc2F5/7iI/KgKf9ohaRZ
3rclkIRBE85FF8ShCD2p+3oQzbuGmhYkJXDkVQpPQYew6RlZXWH40OCeG4I6zMyB
k6l1tvpnj+rovbB+YPeQvntPoskAK1DJgQh3UGoiQW1e2uP5pUHrkFBcBS6DyVIo
HbUUAoNNV8xa3eDVM2zcIXx4NBRhrTL+v6B+6dskOwNLBUio/90MORg2CtGLRPkp
YGTVcDmY0VBbt8qAby+bgYMLh2sqgRNY6AnWiOuO7KKBJxhtUp0RoJzJAWe802lz
1IlHMfXiVNHWpBi78cCPzebU14ATC9e+kb1mIoeUMi8Gj4nkqlD3dK1mviHuO6Zo
Lze3cScVegNtGlHZazZSKICkaXcHOkFJ3G4PhKaLn0n9l0RO9kguHPGwJNQVMwml
JPpP2AabsvdctZlwZcGW/9QzDGoTqGlE71oXNB/KFnuQAZSMeFehBXO2uA0/looS
xgqGRC5ts3VlvxtfMMSJB7hfVcke1Fbs6cWB+HYOirWPhDscNkOeP+6WfwaI9QRV
1Z/pO3gBtrRNMwv5UCvmaj39/XIfKHSDxoqtHM251Nrrr2ucocvg7awN93aHV5tf
ci1QoYA5aUysp3ub9220BJPs/P3myh3L6aINCih9CP9wQ7pOyY/wxPuPEy4+ddDI
Gy4L7D7rBw6dDJS7gRsX9zLlNBDwGGY7kcT6wM4tyLYnVoxfWoRjd38lARh9YZD0
FOr+F2/b75fJaMlgG1pVd3UYI5+CUTwTu5/tcbPCMzY49SEUn7o2sVxsTDCYK9FD
50wyr8Wwr6OAcaOA8EaPw9RjcrZsMR2dSbtFJBdHGusEniNY6Bg4mS3yqDuTQ36U
0A+PlaCGeitVq36k7xJpJCGNSl9r3LDKYFtZzYZ5icjyuBSrOBWNM8NQgrizxCMQ
BpQ9QGXREpQVS43HaWhyCVoh6tLcE35ax61H20k5WGMCcnWiVn3bcfousDrr2Cqg
Rnp/bKCmhRPPqyjAf74O1K4Pksn2uZvW9yhG9U2OMUKOXBb4pO1m61s2k35wszbI
AY04DzVMfBHH7YybAT+qgdFFXE2TMHrAuV+kyPr7HiZDKcq1ALaUpp8qxfgrFav+
XBxG+Y3MT9f7kID6Mn0oZ4y2w7DrPHJhTMM3goha2JylwG885R3/duYo+67bxQzV
0pHV0MC/4zPM6kRMnH5PR0mZYgfoRj5il/L9UW6eL/JQyjpJs1cTOUuwz8ST/H5O
KEEhJCxcc3ODHYqYEW6L6nd5CGtKxkXTNI68zgSreRkJ99DKuu+E4RMu+GESLRxd
qT7/wg6iOgGkz7D7wk3x2Kuk5A2q8YNu0FIYWpSM8GwMBW+RTvrmaaEXqDRZtS67
oGMuxk4E6N3x1JHGFZUBBFsgAaGFHOuPh91aJ2rLAeLC3qBj7oL6EFqNqWw2flJc
mIp1P8RoXX0ed4tzM61cG2GWxqP+PFpoEPlVdPwcOjz0xMqczv9rumv90NQtf82Z
NlSxQf5fGgc4kBgLxUtSJ+dEK56XF44gIgVyYL+ZpHORU6617e46bW9Ph9N7WNMJ
2zC548FzYKB/REjKVorCnIV5HyRRk6jgPtbCz1Uu7QJIEQ5+Om2cKT6Mr6nE0HXq
O+82IInGt/Npop202FNz2hLt8ke/YTXIi0VIMaUP87DiLW871OeyvYAp0fBHM22s
Kq9car733VeucWNoQnIvhmwOm6u3+GT++wAB8NEMIyGfNfU/PmeJMP0mOPgS6Ik2
hS5x8c1cTLMg6Nm6sZXvsifrkVn5nOaX9fY+XUfjbmkQDmrlgqoRZKexJJ7mqKXN
d3/WFiFBhdD0EBLRcZAxS4oVGo2+pvu9+rRDq1U7JERX9CblW8/ggcaumMh/7JJf
phbrDY0q5Ovq2qVn96rLbMPT5kcIF7SfSWzE/J1hK5QxsMtZgKAYzeclhyAP5acS
cLH//EHOuO7Io6VIYO7JAWaZglIu0WTETpQBf2HvmLrzO3c3oI28z90gF3XhxAMd
hQlo7KhftV2O+VBj1YQ9WkJPsJ33tI9pKUlPAffyPV4gv1XO0ni464wZR7faTDsi
cD9u0KL8Mr7QkdIX73gZwTt+0zlx0niSLD9I8jj5gboZAduTxDznb+KbLUqhxjX4
eS2qfvOqrcpIIp7uVUd8BPCcyA0PtHyxJl2rAju8FeQqRHH0EN8AM7btG3ikHADX
Hx03H7RyFq7lhFjCc7OVTzQhMtsJH2MocNTVWJYbA8FC38UdWS0tWbXaUOCsHleO
iLGODBQ7kuZDIRPsZPbrB2VAzwYyA2XjGgx3U6iggfhwWo53jwFS8lIUEtBwD73y
kR624QN3lxWSLjjoCk5uVay853yWfxVkGll+r7s27UvftMrlGcf2xLjIDzgZIdFN
L7jaSkWXWfdwyX0YpR9KzJmzMpYBslzv3xKGQHlVwtoVapRc6qZcqRsjhBTEUSXP
CunvV2cmrBJ9vTRI0PC75ExoFjpozSq24aHgvQd4rp5bIb6ORC8sN9f8GIrFoGjV
ub5qxYyMGeMf1bGZATfGqtg0CuuL2wT4AIR27Zg5Mlua2uDjhOPlVhBKG8jEp8rL
pOWrmZU6b06VI4nuqdGXWQqbcf5ef2md8t0yT4YFQEqyb1AaGDYwYGNJruec0u6/
CwHrqwo7/eWY4cvFK+Q/VhaBmze0H2/WPvXxNpPCFfruKi3L8rTiPegoabQee6aP
iodywrmztcb/OCUfCy/GFR9FP9dTx/2iLVkh2KKBwiKGgH+d9TEqU44O23i1L8JL
HtDo7V2Huo7hauXYS906vUBojBDNxzthja+QE6ojwTlGu0HYWt54jNK8hyMapzxR
u9j5GEj4nAt0MgRQfOpMemu2DPQBj2ojco//Evp7BnCf8d7lPXNy8rXuohjs6U87
wQTYTvxBCaYJ5lA5ZXw4Guu6HbaIEe3HicDkktjtyYEiZqhhOn7mDQgtCT4JNg1M
RpEpwGG59CWmxma6hkvm9GDMbVsBwAStC3Qm92OE6sRs6UfO4ParKxcsSyljgI5E
z77V/eHbTFu03NQnNIIj7ZyprFHfXE4W1ac2BSY/+f85phacNyjp9zCrCJhLsZ84
+kwgrGeOD5pXL9XnVtchA/BB4Rwuo2Vo4VsZ5xbak/gCBUCYA0qWj1gQ8fZB2w/X
N9zA239N/bO50IqVjgOtMuQFWGHkXmI20NpaQ4SgDQl+AMZrWmnavXOEGafwC6ug
ofnLLe0Ygl0ML2TRUiU9ec8IVowf/phWT1LcnyDAN8c7lFHe4U+XFwncMFvobtA5
52cUs39/ZbVjjOZ8Mf2vfpb2RNnZViJ25nRpWHt1nTsk+TvCWp4yfSEGmyF9CXG0
xHh2HrHKMRU7LEcSUgSkSjjCoaMgt2jWupO61ckVUqfen6wpX+Z20t8ouLF1EFBv
Mqlf75dHbt0o8VU4mqPEIfbL5xjqUZDvb2BB7PmGFnf0bLeQFbVml1Rno1uingv+
EcqhZWx2pinADOH6h9PdS8RE5shDdmN9hstO0oJr5U1hHygVQpgttqv9HExpsjQK
/1v2PfoploLw7H/G/dFqgsezz1Pqwang3Sbs2fkcd5brYuv5u34cC/SSaxoBOCb4
ptOpgmIlh+BjO1KePplxJQqC4a0TEMHgnG3nPHTBMS8oAuJbo04QVyVph7S9loHH
An5XcrnAw3cww4pst54W386hEIztgp/PW/ZfcDdxuCE0e1PFgGdM2qaSG6NKYrj1
9vTj6cEJUwfunSx/c9IjVccLejdwc4Q/ZnkMV7t20xnc/8ASq9HARI+uywqF3gqe
zIGQdoUuy6xqYM8YwF3NC4cM9W/5sYDJxr8V40oST2fDA/wMl5orfl/VKFRRekdq
oY17N+FLUwrEZtjC5B3s/polVM6Sk4lnpkKZ3NpfgwvctujG5ygRhYfh22bd+RPH
DL5B+MnmJIRRX6DJDA4OL802BJWce5vvKVkSrVi9or2BE+OTmcoFjPu5FKKpnpIB
4x90dlDG3lR/t6G27X8nDudYKR8wRX1ceGTBz3Ib2GhTX5Z0xGafwceiswov93kU
tatN0oTTMpl0LpRyL3+z5IgKnuoCTmIdrM89HblJQullng3ISI6BOiemIlh4f8Ve
btqmjH5DlLWYrMYOPx02DzVsfHOOf4uYGwWZc91/NpZiODPsEI3IxFq9rVAvJhCm
FgSx1Jl+DOWUVDnPGunYyVsrCImLWiG7XGvwjnOTPJ4I59/I0jgpjvRcsIorncpF
X2ZROJNs0nzBGdHRY7T8I3z97vavzkEfNiWPC9+DnyqqPXe2UwCZtoeP0cS+ZYk/
1phzybbEI/zlyX/D1gEnl7PfCWDCrQPEgm0mTR0PFyJBASxtDDFL2Ohm46jepzLy
D/sNbnglP1Q4QqcGglmqjAL6wd43AXMeOnqZyk9EP3XdTC326/Lfb+o3dLS/T/Py
53ejbby/fsJVZDAh4ZBBcFNQUO9U84OMj4U6i5csgVxiRxiiZ0JRFqBc9XuekTXZ
GXohko3NIijMoc/4DARWNMQ3J6c4QJFuAxpTLEhkFc9xGko6yFSm9b5Yfm/oLIx1
JFxU3v4wZXlm5zFmO0HyRwg4Mi95ySRrdHwTdw70jFmTnwTrk4CVSt1JD+ygCaSf
pVaDJIX+KC3MkA+xhvgXyMhPz3KrceX+hw9TGHlNuI7SXZUALfl5PkeCGape7pub
nDKbRLHe/zQfsQkqtKF1MzF1QPpSm4PbDKfLZuFdZ5fEilaTsef4r83x/Ma8mb/g
6SmQsd+refY9mQI61VGxmuKAYNneSSocVYrn0rL3ArRMN+o82Eh89HJFSeWs0rDR
q3zd2MvH3EQ1/3SLaTh9UAYEzMAipNHRIlQnNSsb4klulCYVaL2xYo8mhRiKpU+C
i0Bl6f958cYRr0nUGw582e6GtPrk4qsPJKojpdsG2ZmplFzqs81EVkBP9h8s7qL3
M3SR2mraXWiUaufTlrfn67JUNOhuHZfjX/KlXefYs9kA+i5f9cH4lrv8/JCH1t8W
PjyoTt3VzoxzMWY2PYr9+h5QRRSDJoZ7sMhAF67OF7r3r8htp76cAdqBLqzfCjVN
Swlp4JW4mb5iuSuomfxetRVkdfX0cLO4OvW5j6OAToZho+iCTQjj6Bi0G7ztCd+a
Lr2jgmF2QdS9D5txZjQC2M/+89Dfn9mCPNVSV+/SqJL2M8SASU74lyGclAFMgCtv
sdKgIc1hL+RaJ6R1NGrR80zm+zB8Z/Hl/srKU9LqxFePeHJs6PhKZim4VNbhpNRu
XWzyA2d8TGCnCIWMoK4HGuxO/CHgR9DeP2qbWRvO298/qK49aXio2jGJveUaNLpZ
DmP1HBEK7Fai5sVCc74XXQqOivNLHwS/x2vniA9AzwXeGTrk9YAQE2gRyssydhaX
WTFzadhhkdLpIp3gYoiVSA2Xr7pBcF9QAE+Av99y0v/LJOmGSZyqyDiLlgk16mAk
JZLDzSyjVHqm6wp16MccNKpecqFkCUPTOjRltMg+68bLqocH/KR8ovSekExbfxD3
7srPFkz3/mLJKtA2GxYp/6xuR33uZkB/6dj3OpBadtkaMYcGO3VWdql0QZ1gLs1D
ieQoVXEQssXlheQHg7l3Mf5gXuMkeaCNwtqPmkrC2TlwC0mysQ9I2kmxnKRlcxtO
wqjLhlRHvuYf4hJ7uJPFz+oYzR5Dz3e1xlGRPk40kQTZ5JMGhqGodPp2Iz/xb8MB
CgpjjBiYSrv4CO4tUBo79lZnPiJVS9dnXleqVc4mVb2rD2CFBCIkgfcEwCiM6YIq
x0OpyulHyzxz+ezb9E/OcyiiqV15pmnE12rabp5+BOfnB8FUdWsEj4Q+YaGz3PRi
NTbuhc4olQ6cusKltg8EVFxWifUIO4yjkF1oz/z4Uj/Cwzl97NAhPVhmqeBhkUN3
1o97/pQ2cBMU4UbyE+GQW8SMzscmn6xUH0Xk86ROsBODBrruW7EMF+PVCIbspXiE
Xm1SwL7V3zMkmdvjy/3+iZ7xpLqMkzZLkQaAO2O+WtHV40o8USzbrfZ3LLc3eXHu
O2JsVHsKk0bszMnceONo3wCXQcK4SJt5gbhxNPN6EZ61ZN//dEWPQKKLhY2jRzvA
mGRNj/EUCJL/hZ9rtJsPeIrw2K1/z1x6y097yFp0793eY0nV8t6Rlamv717av/tp
q4032fDq2D+Qw5DLWNweZKof3I+fC6KqlkWOjBZdih6vP8eXRFBrpt0gxDd75i9g
Q4T3y+I0KPJ+okb80zTwXPDJ71zkWWY5skFKUsQz48KmrmxR952zkb/NNtI8525s
TFHs49Y2HI/X1N4iMKk2DcmkCAgqTA/3guyX5fwSqnuq4HDH5NWCHM4RjLJ/2OHk
ghw+YmYatXZvQaxjP1WLBi+Yw1Oj0NXp81ODDl4TC8zmeTtnpQEGT3NWwp+QcHXW
U2ZxQijcf04swcuYgPMTAVeRX3OD/JuVP1CinqSuy77FxCbJXg4SyI9gIVfjhrbJ
O7T7JkcqHK13xTZCYMXKyeekNkG8JwdQYttol3LBIPz5Fg9w/QbBEGK0dAI0rhrx
MT5ocw06p8Ljevz2FFNn/fO4qwuawgcZ9bdRcVdYxLpjtYEEGhjlFT/TpgN6VkzU
zcgzK0MT+6fDpVkteSOjmq965PNVI9dOpiqwID9A4t/s3l4GTBrBEM28eNPhEZs/
da1BDTZZlAG1mtiPXbs+Nm650A9IGbocWLvpEqniVBjidi/zPtjL5kzwzikDGZh0
fqFu+8GInWbMucD/vELdEkqOvjr4HRK2ZvF1+JtZU1XaA06fTiaypfvrNxW5zSNz
DwLsrHi0TxHnm9SUNlTjRPD2EgflKfwvMhWElhQbPDDK4HMMEMeFk1wqMbQl6XiL
fC5iZaNWzfdIJzx2VLeM8StikLUY9WLw73mnL2G3qWsTosQAARPxdsvvHCOjLiBU
JFGp01wiF/TPA/BK7dBBNaP2R7njgqIqRooh/KCODYxcueMCjqg93ZQ3cZLA6w5V
M1KwW2W161OwKjh3p8PbVblCns73GmBtSLFXbvJnALX9K3928WvCCXkp8WIz8gf4
g2uQVTPoUcW+xGVZZDT8F4dd0Zf3Pwakvl/kZR+bbXfg6gHnqV0dMk3n2pSLVih/
Lz6mWBE559+cu5JykxnL2DhjhuAK4zmJQhHScIUHzDc5exHnkAgb04aECXippER2
+ybKz6iAf2eFe/cv35EchXaIzLogyCa6lMPEH/XeUaYtHHyeNSD+6AfSVcpot51f
V3zP7VaonIyF+jtDFmyrPC704AfInbGkqa0o+QHBgLi0OUQBdCpBNOPQjGoQErZ3
xm77+QsZ0f7oZ34lDYYKKvaGbcFgUXXPHIquqQFZrDKz9hSZZiSLapHJD11dGqb1
WjAWHR2hL7J2C4GBvBOM6WbJQgBZsVJv3KL2p1ja++6uHBWlElA3lo42rj58IWrL
5RAFcJKDA+sWJo2GRnuK4n7sh4JteI/S+0A6/U073kjRGo45IGaG1MzydTsNZ1TV
CWJyY/+rcdVxgHvqpq5qLiyowJD6T5dyXV1BmsJ5+S+Achs9cBprKjMgtmlxHtE5
QXlLicMMyutx+kAQmnYY3/ZZI2NELeOOpsUiomrURXpqa2yEHu/mBaPqyk8I2FhQ
fov9756Xy3qQNSFaXxsDhyLUtJLc2LUvcR7WliuzVEK4v8/bovIxRUVFZvF/W1m5
BWPNCicFpr+N+q5VOtg2dSWnhkb5kebA+V7ReVehZ8s/CP/KOyLk6wP0BRH60Ezi
D9HB2JFQg0k42tczdux+vFiBxlHJdKsSDcQoln6g5FoMYHkDPTQftKU8FVGQYMNl
8E1kA138f48J8VZcXbu4Lgg+D0JLsKyDPjB0abCSRBr/WoXokyDGdEb7bRymA7Eb
yI7udKBLOwu90qv64csTBvOVAtlerVBUxJHXcax/h1kmkbRl88eFtMYtxdbAA1Es
FWhri8Nsj85C6Ir9hN+hpIu94n2tehOPv4cxFoNFaIMBYmkE6c28+pFRwCj0GWP9
bHkhgvzKrB5nCv8rvLMmGtskWiD9VSQkjR5fUJf1ImRZH22t1TA0cnV00kkPqH7E
G37Z+zuCO1D2/G7e9hQY4F6QiCr1g2nrpUwXiADrSFts6lpbyNf2CJyeydNgEeub
nK/cOsAapdft84duaELLzbjqEI6RfJ5SIRZAtsLiTkmdtEaOvzAD8YGL58ukpGWV
7UZSrTMadrUWk4Bmnltw903GTQ6TxJHAw8fpu0DMYqb+jqhKj1H4M0cYe7/OoCBv
PLAOZI/kWVe4NSXEPJKHSjG52tCsRB0K54BNRhqOzWAn+JKhQXQ5H95yVB9kvv9t
8DAnfYOgqsFiLn4WGJPfTo42th0Q/UlucYiJN5EoM1V9W611nz2bwsHjTXSIiLAp
xdK84uSr4UK6anpPuwY80UnqNt36IOyzMD0cI2JOZAN4oo/NdsQ5/97SOYMGfL8n
fNCahKllueOqCofyC2ZKWT35h4jTbqwaoQDA/JsLEZMvXNnwCuAwteZsOI8gitJm
z8acEoSV9J13kUin52jgKZkcE7TIPB9rOHYwAiM9NijvX9ezGHzt4j+vn/KzqRde
LjHlUyrjk5rY9CDzWh/Jv3yXU+/e4RTx1RKzNaizzZb8EWNpWrlnpQ8GPXQMMGD9
giWh/pmTkQY6U+lhYCREMybRSEvHIqnYRvmNDf+RzdttNnoXVzAhxbBkJUzny2NE
eZvPGCKJyez1SFYCJne/x+6xh8xBqthT1ECo+JXo+vefMgxeAnr8vpk/qroo8Qjf
aMlYWcrkNLawH+QCpuSZVwTTiI2oSk8YrqyOt/MW7+t+gQ5DN84pj25lkMKG8fEN
OvxEMNR8K3B0z0AcJ0LRRbvG2hh4UQQVYnzGdl6u+tdG9e3LthX5HrOATN389Dqg
GqMzQbHsx1dRFxF2nbxjBHSX4h/b4kp4agn+xkkU+ZAu6prMOWFqLZ2xnKI8xwkV
C4HAI8s6gBMDDdW3Z8ZQyUKcZ8dcbHFV1OJR1J0y3pvsBchg9IVScA4w2j63TQ4X
Gyc3MJYgtPDk2va+tzlKo6KkEUjhK97BAFUeHLHVxITtxBze/MW/qH4D5ilBWDRY
x7X8Q5izRPCEKZzN4L7y73Q7a0wAz/gbCTKTpl7wzyNmQCRi4E+hnJVLTnMJubgf
AF28ja3E9tHHB0x9y8oGUIoAC+t/2qXqtfEivKcCDK7uW2vbSgNf+YQOwY3+nKjW
TTxHIlLKl53dtkzocEof+VlaOVqoBVNmzbLHNn7drKr6rwe2VSdcjZOQireRBUV/
cY9XzAu2YFKrI9JsZjTuYcXjvqJVYfxXhQPaBiwmga1Xxcp3aD9Fo7IFqW0Uox1h
hM400u/dU9nlALo4okU731YH2zHzbZ1+AwnFifj5so0b6lCZ6DOMiRyTZBrXmw+L
6t646wvX0/HdysqzNmRPTewCuwMA3/vzov0qH2NpzVOpfxzIk7pEFq97DBIcPEL+
4ViKBCjZwKJlh//+GJqRok6SoT90Xr998fNwA34A5uf6so6L6fhthmFQKNSQmq31
1TGddhtOyYty60D82hzCQYR5kwwGIczdn6MoEpLwN9u55TzINaaYMQ35LULt6VQL
cQaqDsAbgAtIT9iyputFk7jXgBqx7dImDo5xpi69tHaEc+PKMApLpj+8ne4HHsRm
j3upPApBQiusPzeO41+Chf3Rcx2/otcZNwapKydwV3Ns4XjR3mpON5JXDtQ+09Ac
P1kNXOhFwFansS+4t8Ewo26sH1jaoosJQL+lOR4vggLfGmy9ueAZGoZKOIWFcy3V
5nEwX+brnI47TpvRWXfe+bRR1Tr8Nroz1T+WTneyJ4XyqGXD+XeB5RCk/4RcmW+H
k6YRfks0fabvTBGnH1SnTcvPCBOdiVjXNxEKlekhjegRr9gbzKV0Di8etx2d/JPN
GUycpVDQsIBBZb7Y4pwqTCeZAiHv6f7rF01gm4ocrlpWoH8/2APAdWen+YoKhFpq
iqmISkTPBHseOLyztJkNd0gGDlGis16WxhTt07cUFn+3kUs21VvcBiPQ7QK1YJmS
6aGHKeHJ/iV/W1U4ju+WxvvjQmncoRrpL/GmlU+dv5/N6R2xYOkal2/+1Y9Xa1XH
AzbaNx4pr9PX0F38Fg7x0RAz/qTgczx8LKphp01EwOMTl3kLWdpAXtmX9oainNkF
44vrBgMxvyA0jiGpUGIln117ZVM8sZ1NytOFTwu34IL1s2OfjUSRLSoaTgc2fPNL
ECQ1k7g0LFBAQwtV7m3+b5b1dkkla7eIvW1vMWEQdLEV7dCW7AbMZ+n+O6cqL8bT
0uOo+Qtkec8xMVIr4oEilzm90JhepGV/QBwK77TXpoxpY8Aru2/e8ZG+4+4LxCmg
ygyccLGxqPOLSlXPJBDsiOixRNZsjB3/FA6QagxEdRJO41vJHvS3Tpfcof8gnkr9
aVekTO4TfR9Cj+s8k4WtKJpOAZ0cUuLK92DomK5yYg6WSELNpytWpndFhJjcpieY
oFVylLBQ69+B2Zbc1mF7CnRZOUkN/IyL1NJEuD2V6tcAQzVy8L6+re2BK6dDymLt
JzsusKhI/csb4Hh3sx65/+ROOcQ4V0kVxw8gMR0/etVzgsjcG6OjNk8pBOZC/ICo
TDj+xqMw5P5Jo0jIfOPYkZyLcwDPE6aF69KwsL0JLZyTbw4RJtFIXA1k6D3Y6mne
rdcdyQErkMEgUSuUh3gqcShWMO9ZEwk/uDM68TtKYVn7c+lI/o1HiJPuNncMnWlP
58D3fGTVNFxanLRkpjHTE9HB8BdTFNuPdpv9MDVIAiB8bigamCjjF6JkwYzMdHbs
3LKILaU/Y5Zcxwg/OaRjHnQoKb7Pm+Yru5CHCEzlipfgWXCW1dXPQJnL+FYZxHkz
ZGkYCr3OVVu9iD7kT1KzPIIgm2oQ+AnrMvYx5ZpBPb2sFsJSkVnI73X+gCrYKD/I
UP1fXnmbl+M7t1fYZ3N/Jbgk6YcgX4TMG1x2BWWQc5k5kVYf0kumrSH/lF5B72GA
jsMUWtUKjawFkZ5OA6ljGtGqqbisP4UtdP7npy8kjvX0uMR+V/MBRPE2B7Tw9ipL
Ys22vlNY0sGnI+uv2btof25GIs9Ml3KvyuLB4XMmBZj2dJWmlliO5feLV5LZkVP6
UliAB5yTCdJOwDdxet3w/aGzm5zdWKkwTmFqWscagxTY4aIoan9NJOt9Uca+v7iI
bm88yT6NRRWJ+vqxMERB/qeO7tk4QO72HeaL+wK2tGbXcfZmKo9/mfml0+3sSC1j
jCyMv+BRWHkjO4fuqbCJJOtwcoJgzqO3Zfy0jXbM/Al51WTttXxS9iRBNnyTuRg7
7oQ5HgtqlJ1kEdvYrK9/7FQ6+lIkLiXFRRm5dLzq4U9dFZNg+HSc/nthJUBoVCfJ
83t18edPzkIAyUIBSfLeybLJRryljKBHHwKp4NL5CY0o6yB4wxzsPjXez+++Mq6W
dpaggRcItHVaMRDlh/CFPwsCllyXt5cTNVS+67CYZAzOqP+2sm9d5aYTPDOe3HjF
TETg7x+oK+xPU5qH1Asegh79zgpShm5jmuCHNQS30NvztcYoLYiT4CdOblSgDgpp
izn2K6yt66zg+6xKAE5xZdUSMOrPZibnMyzXz331grXxJ8yEQLZuQRBz0Z2seMMf
ryiXmjIcWidc58jqWqmpuOw4XLJdjVbPPtqQgDuH7+Bvsc87FTdVSehR/DCuXvlD
CBaktrAp7TvEAPgx8CtIpL1ELQew3D5y0sOrhZEabNv7ToFSeTx3GYMs1RAcjDIg
yOLXK1tSXBUBQjqN+xp/DSGQzqJOXklKmCCjHNCfhALLxN7UDQZFlmy3v+x84AO5
Xx6qPL7YJWZVUBJLgR1pWrzISviKL60f+DBBVI8nO0MGDGazFQQ5KUR/GSxpz+Al
1q5gXliOuYJbR9snta4WFTrWsMpht9F+m3ghsrig3nzoHsCaQN+ivPEGrlhV0htm
MUfxL7aLqSM8ANq2neS/1eII07KGi362DV5GCwzoWaaSXyXEX9MHkI8ATkGSyhqn
CTAgGIGkjgPchTPPMYTWD7zyKl2cu/Fe8n06lNZKraPQArJkqBlCN2MzWoCZKcVC
yAAoLUbTPi0Ssy1nFIlfkVcXBT6560lgZp/JTIB+Lg69gpDfrQvBUwlQttBFplxz
6aHhECeJYBA1v7xXHJ1F3brgs01/zn4SG6eeqRzCIl8IgUKY+qJzgK5QJgnGQ9gt
yxpKzTsiemWB9SSfOyEFJjUN98XA6O0CJMttsC3BxODpR9Cdbe0mRx4PXGC6aWDB
28xpMdAMEmAUgjt1uo0+DZceptH2iTXaiZFvY5h9OwZ6KfEbefOC9pxcEJcSj6Qk
coj/Ot2dBSL/c7fq+YffJfrjtSImWJQyPZhjtqPSZngdQzwunENDI8Lh39Vc2nI0
2rEWI1oJZiqczpUVHeMJ1Arx3aSl8CJrodWkK//vUf7ZCdXlYPPlDe9ZPyNioe6s
eRka1rnxWbbA9O1t/oNusD1mkc75ViQMT2JwiZo85bEtv9MdXY5MRPJZyntMPNaN
tO9rICNcuwpYZ0SYIlJ/X/A6rGSQdI8d3k0qHzcAp9soRHq7kFB149NvyHzZD+i8
s2+Qrr9OZtr87LKpGAjc1QdJ44jY6pcpnIHpxkpxpZ1Ls6j9+EZ5vW9NaMWzqzQk
jXVcd3nBrGdGZzm9llgJvBLyhpXvNZ9wEFYO84bxy0IL7iz+EEXVo5taakxlSxr6
8eOtycnga+6R/BrkpKiHU8BhdSLvUc4pSZTgQQYK9bxUK9hzmFsx25I25OB3oFlQ
GeCykancmJxYuWF4SYdS1KkDPpg+sC3KkeIfapmc/hHbpaBAvkUgICjHgJvWqT/Q
ftkUEgE+L71xnaEB6iJ9Vw1P/Hwfmr3whXZoB/9UygMCiKpxTZV8zxS/+nzgcXap
TmIrVePRNL46s/+KPtq4NcTeZbrWqdDXtzLKhLYyHtbDNNugzWpM4Uuv0aG3E60Y
6E2Ys0e8SVKu1WGqx5iR/D+7GhK74dSu+137OtEYthT0KCk5p77IBhXQmrmFAZ2g
9XQoIirO1zDjWeM7PaOvzCwCQWLNiSF23qdpn3WSRfmlCrm/EdEfE/SzvjXAVxNU
H3S5oX+o/OuT4CX3jpBrN3ePC8e/43BDlUqdvIhHfLVtNh4ypZtLlzgVVAt3Vqpi
nPDVFuJ9TDIriqwsafv2dGcy2r7Kb7tNne6TTemnoL05w5jrHU4kYcuJQ/FvEBsS
Xl3YnTBKNBv58hjwgp4ANh36SG5N3wSFIY64QCxe7cXUNKsoz4Gg9G/GxS7M1Phl
3MpvkoHzYGGdrW5y+/PgH/d44+gX7QQa6m9umH+LQGKu82bFq7JFI1PprvKGLcd4
phT7josohAE/XTs33breHFD0NZSkWUvrhfwnNw5NWijyA1Wc8nZqhoGgKiEzOIwY
edgJzRu5PZYG0y8NqBNyQ4oK7stxXHLnd8pLFHUVqrgmbhRsuc7d71HowxcBqCBI
D7otF0y6IyxjJXCwz19bfGctntvYWAccQ+ICrmsz1O9bzBeqj0UzFqs2bEKg3vRr
MBG8elFExtB5WU/U2EnRMWApHe8xtrYM+rgvoIHDVL92pnF3QhYlMOjz4b8I/5lD
WKCFhiaRRr/A9tarWV8B7BYO8SwsBXi+h5D7Iu78zw9nQykJlrgvyiQDxwE7H7PV
nfyhRkjSiLa9SWRhztbLtpoi0zK7DLNIrcs5ja1KJHgIn/8PsjGsNEAr+OJmGf11
403AUEXkRLYd+IJD0+XH5+eUsgaj46hi06IeBPLgBmbUcsUf4x41ygceixRHjpEE
1zUPYgvqQxJ9jM4b7yldlwrUkcMiSaMdq16uDIiGlxt4uLyM5ietxEJPn9eGDK4a
7Qw8PC60GEwPHgzx3gxSFdS4ihufctr1UgFW3693vXLOYfEBBYzctTg3jWXOkjxh
ixI5wqVtT81IJBs0CgSt9JFP+A55HYsG34se3UQtIcXQeUMuptOYtCPCcCBldiN9
4f/5QxwbxonySJVZ0u/3iLl2rjYzbttEhxuXmbD3H5PQFAJZRwwDFpmV2JCTV8IY
QH0kJVfNkpE1gh58e0r7eBP5CdS/xDg3/52jeJOqgid2xNroM/ZDFYc7m0KrbjHX
69E+6iwvuBcXoOJtlub6H6aF2jm/s/k+l9lgrsBgNdLlzPQQ0a3oajkhAe7+1uz4
HPVoD6dKoFfLYPp1hAnFPKUkV4jRt2tcsnxXi5Y5eVdn24Guk2PxXMBW0YNHXXdO
QXBf8WppCRXrnqH3/FKG2meCqm3kmMteSvB2u9TcvnR79G98K6ZC+oa+yRUqJqoh
9z2WFGS5hkMGmqhwy9yHRnyYDRUIk25X5GhF9UvHlqpyXP7oB8AX9nDjvsSf3N7X
GNMzrsvZBA47Nj6Ej24t+oneKL21shkk0/AnaCCH7o1CWc4qdm9WMhgqVivPryI0
4cRD+7uPykykNCfgk8HboOHHBbtKbNQPlZIWF1QEeUyROAr4d6JXY43RAiHIt/Y3
str9rMVpqnWwss05iWmGuK0yNIYVuDfd+XXEZz4YYiBPllCbwVAGFsWEQQOnqW5f
Z0HvoYJcPBCp43mnAewcsWxx2ZcAzwlVPcbg1s3r2HqmsKTv0CakHrsaooPzeewo
Cli41OJ0cdjHzTphesuXhU29IcVwk1RoRcroouLnOzsN4FAKEaCis7+rg0eU+mOH
cr5zMrTka1HQ6eCHOzO3MHw6P+0865hMzEKJrWiL51jJliKWp1nFuUd34oL/Z0+K
wWR/6Z3px9SfOsS48gBBZf378c5NEN+UWGI6u0MCBrSgQOQ99bJfazUuJn95MzrI
eg1t/gc8ny+fEI19LadRzkPvU1Rf1Pdx1OY1edxvv8aBKpDyvtGrd2HIaRdJDxCz
+2BGAST1BVGud5QxhVd/RkKDQfZC4FSGwQ5Jv0EmW34jwUrDC5VTQTN2hfRGypSF
90kzltfTBaOF6xm4a1er7MoneM69BMi/Qge4puGg9L92CbGorfsBuPrTOtpRQYSS
WRbQ4FCHBvC/Ii5ODx0I/atrxF05Sf0I4cLhLz2sN+MCB2yFehBnZdbrdMjz3fX+
/tx7QPhGZG2VlNsmGqQ/LjT15P5M9VGCA70WaMS8CRzV59WPKJGfxr+Mam+EhRP3
JHWAU5LkGSWh6R3mW3yzEqz6nNpRujBUhDUVYIfwnmf5hNI48FfsM2zjCBCLFzXw
G2v1AHL+EQ9Y69C0I2wyFxryg3FFe22l3uD8Xl2pS0g/V9dNS55X/1I8e9UREFDW
tywU96Y+Ued3aF9hDxovpXqg4DbnGJB1HvgdVsgHZdgIK3Z4fly6F9VJ1kWAnRWz
VW0NX6s7EhOy30nNge+TE2NLqjar9W1lx1GJ1GN/mOh/+Yhyj5WTTbNnrZlncLv1
wM6A25yhry+j0AD4NXEBJD/gnkpRvmN6SKN8HYxENCPg6226iyaWhqKTpz1kWN6l
rXnaDb/4AcWGcznHgLcihcxQssTq3e0HNQHrTsuSpovHW+ODC+bnteY4Uwj8qKPK
wcNwwPJrDLU2QjZW9usbo9U5bnRGMPnFpDRHOlKm3Pk1Tt13aMmllyCCuIoI0am4
H52vjj4eXnbNIMGxP9r2FwS88k7VJKf6QbIUiMYXd/aMfD7m1AQYhIjRopapW458
4iVFREr588zjB7nWILAkSR/8ZaFCdOwEyrn91roCN5OofnVdhffM0I6XL7TFMMA6
hN4KmTNevum301/Lt1monqAIU6+ZzKWn7eNcJVzdIp72aKvCk00ocVeD3GF9ouuI
+xFjhaJs2UI08eOimsA2ZrMlMeglYwsyN1AVBz0vxj0FpA9Gz4r20AZoiW3x2ueg
9sIbdtvT4uIRnhkZOGHK3idJxj68VOCbjjZoZZy+jglFRiQmeLT8TSw0iSXGRdEa
7DisXgOL7p+rZFmfyaUGwsMgZ2teDtEN8bajBufUZUjt/lIqjnEucDgfM0JDZwd2
UDhIpO+iEr/wHPvc416P+39H9BW7gmbC48Ykavv0jQSBQ2B4iaOZNEwB6nAAgbKV
mD+SoxUNvIEHc5A3Bg7pKZ7C3UxJtqPGPKX9spQhNKjFktnT5tiwPDNrl9uv9mTd
XOxU8itaUrQ5Mah2CxT/zgRP+4DK24LLVfo++QFzv6r8A+A8Z+K9Krda8ZzJYB3T
X5/j/iYLxKBrszBWiJbt5B1It3mzGK9XOdSVicaza4646khBqzvcLQ0OiiAT62V+
V5cX2jdUlp0sBy4JzQSTRAuafvc62lDZIOYgc+hnc2a85tHBXNOt0QicTcKioNYE
Bow0njD+ggAhBt6d+J9jWCuesaxFviXyhE2TtJRxYOc65H06pXTXhYQhh2Hz2Csr
dpnxKFH8e2geveMcCnGJyfQSIFlWm/E22akh/8QkwCgRNIC+frPJ77C8XjkqDO+P
MHYMKO6uEub/oN3LxYbO6BSuAy34ghT206zrKL/ke2Jl5MnlumT+9SiYSooeI+e9
JEQ2GAZHEP1JSzou58eq538LTN9k+1DAzHptCYS39e7KHoHxMXgCpk4c5qXeDVpo
R/KvxWzU7yE65nor+yu1MvWZ+Gw0wiLRme+KxFX4ultTe1TLQwT99tWjSxuZxZh4
JbTSH78lFQtr1biVP/pbXOOMgniRIm1IlfyJCt+FFox2HqNYQk6Yd9HqmcEy7lZX
SEDwnCabUM34/JBxWeXdqaSwoXeoElrBvPpUsbWNy+96XEEQ8C5g5phl4o43Fcvf
aEwAYzZXOZ2mn2Rbzly181iFjGXl/Q4ahhhnBXelDR7zeBHJnMmtU9b6+jv49IWm
lqK62LKPBaZKpDvdjcaWLkUzY7anSudyuO/iHA1KDB/MpyHf+PyFj2xUBIkFzrIC
wU4euQZ1xoXYl89V13ZvbbRQd2gcAOp/C93PIGotPNvpNF9CAruExPrqntBK2mVb
TT1JTsJ5WFLw5rYOL163aNLQZuFITeYwjO1RO9M0bnHGBet1W2H69b+fLguyuPI3
7AbxvChMXQG4ZG6u+XhsHfLNIHE0tjUO698sdrzQrkItTpSScs0IHmO9QYEsclQ9
cT4w+k8NVWIiEaSuZEfq7TfXQye6MJwqrOcD9xGl04y0lMJYOhV6hGtz05Ma8INE
ozKQiSR3a9eb8O/zDe3YB+l09xUOavlVbJwiVGtq63o3dzwT2N56lTRcD+xXz3MD
S6eyPj1lcaFCo9bVHyHjhmerj5c+VBGC3XduP8knlNwrhMbmGBvMqWIGUiZ94ATW
0OVK/9GxdWpJShmQbB6AmlYqDl/g/XKvISlNhOGn09+WTczpAj77p9qSdzhF308A
V2zwoq1fF3W753PzFQVJOQmENsSDa8ZHFTCrpHvWwrfF3pkrbiAsi+xSdWHke7cj
StPulfurNXD4/TPctCko6TRnsuGcUYeE9zoxHfm23wmVvTzQvj7kZf7AAT5sMRy5
ITa3QVhtTuR1NrYmjUqWqNOuKjzwSkSD28UqQVIjzihu5BNMyYD9NspbBHhX+Rl9
KFfj3PiVsjqZ8lZHhk+V4reIE45g6xFUOthW2Xrpk63QA1s1SV1wGppxfOBdeuyT
XC8JiZmYHS+Falt0EYusuAVw9jvMyQDDf0CC5SscS813ZBFgqQvNbo1lCUMtPA8j
06oWhsYcr8+5rZ24TRajRMLzeIQDnwtSgSgDC8LMDiN88oINGNe/w10uufuCztZ0
9bgYk1Sf5HL75o9Tu5hxWgwaoY2uS6LJWEmOWMyVVo/sKpRDlpqSIqcaBliEo2fW
pcKBZyXYoaBDB5yLrOkJL0BLRpX+t8VKMfisjQPT51UCrYrccEkcnv5K9KlB9pal
OZvi3a/gpGJd5Ug6IZrcbIU06pA7PlpE/O7q0nNoyXmxW4Y3fomnGK6fm9zw65ht
ulRK6vNFQdjqUA3SLNlyp2L9P92en0A2QMFjrN0TX3vj1RV4e9dOjUDL+WIF2o57
XGJ28NDddF1C1703mSvC2t6gd7UzbAJxm9XIJold/kHXOD7l2NhYsjvmlW0nebns
52l2UT3FDY6DPchlealKgT/y4D73qbeIBAiuTykh+YNLub3qwrjVf2pyWSF4XsiG
/kjBjSyS1mmgnTY9FvI/W6plS/+ZPUw8lq2O3oe6v0VKNX5IrE+ZB0nksYoluu68
SkI/EQTjDp5Xjt1AZOWJ1N/Q2F+OEe6MjDArTLbdhrZOYkJe4g927HQ0plzMqdWI
rNAWHkrlvB1tXCi7GGfD1dTRMi+v7GYtnyvxcDPAs0u6Q+EiS9sh8c7lem6mgQ79
mOpukgheRRgzT7IIp6tnEJ+Vs03nmXOYBi8dQqnkOBjVzaCqkKwe2aLzUQ7LFg5a
zjUG0fAeX+9XkldRcjx+iiEXHvpYi5Ez67jfqJiy28kMpVEcHm2sxKu9B8wohOrh
DmP3xa8k7B+yh7UzKyR2KqBenJH9ZN5Z17c9bR2CLVgC1RERryihDOOfiQdXDc4C
A6eqBhMmk092KfYMCoEJb9RLtVE7ZDjFWCoYgq/CPFNppxE0+3Gt7Kt9xYQFfKpE
aPBH7sojQUWS8vBzSQcQ+CDqsDPkUyfD7atjS0MdsbKNz6LpfywZtE1orZSexoB/
CUtXrlmPvTq25AvhcHOFB5FMyLL5XwEaFke+OohdTtNIjeAkr8VUTTwyWo69jh1T
k4kMioS/8vYU2C3rIpyRIrZsjuox/TAnbmxgjkGXDE/6dPlBHaQ4+BV2iw+52eo7
QTLHj+Z9GHEvZ6nUrdxU7D57iSIdo3q+dM/41ZwVCxUo60i5m2avl1vqUwd49PXd
7VfPw7FdBv7AaIyD/MVl2wuqa3H9RDLuS3VhUJ/rWCp0WMyQnJYwO4EhaBbKa+bF
RLM+YHaxZUxDJd3m4W96ldl0VJaa6C7Aqgi9aK2zq6mbEGuVDzvn0dC2Ir6biTqy
qErz2V57TY9fN6L/BOJEsKitqnrAyQ82VrW455pXp3VRZvdBp0ssIjavWHghET07
uoFP48LYWLtRtNPcIpGvfZxokfSnvPVXR92dd6ryPDScWvRROod3Xoxy7JiZrqEm
Tv7vEFWz88dMjv9wk+ryMEJaM2GaLYrotMNdBSvgpYrPk+h4nsm+WAloD0NqWGY0
/FC9wambfDSA4pimDPR/mO/NLY0/KWCBBXriWDe66xXEjhMsr17Ym5lti8WbycCo
TsM/VRDjRPyUPxSIcg0B7K9a3wYzGQwvpzO1+AC/EI9iQ8o/WEfXXerYtnXIET3U
ooSSc7jlk7UAUq6GXpi08e96WHa30n66EVvlndUgB9RO1L6VPRxRHeOfEbr02ygd
1XFwe+dM8Wdu2Sg+pYoDTR8QRbcqYSZovBuh6/KhfeuBOCUvYcyhy+weKqT9IPGD
uAqDy9UtqMK6T9TfQBb677egCbMrArn1aHqR0geIiirnWo+EAkvxVoQevIqFNr4C
GhvXTjRzyepUR9GaVEWLQ99w5GCDR4Z8dR2PUBmYDIIQD/cGhqGolknXj/876Mxu
g6B2ELt9ApJiAvsAiIbvS1MgHlD7KRteIDrOrlIA4u6YttGbXFq1io0R1LIvI3Jv
wffvsFyLisCtg34Tmap/087SmTf64p8u06oAvyqck9Gyx/H4PJyey1ioggnc6ZZv
FWvH+x7NLBc42LgLYjGD5355x3WEeIJX8tJUvaYA+3ItFQIql6D0bPCCdHu0xdJB
LyCk22ttiOw7A4mF0eJ+b/hq1tlgZwm8CunsPpeR9Xs+Z5EKdaqvB04JyucIj4I+
d0PS77hTvUCcMaLfm3PO+/kwr4xuOxFI1aJvVFOPGCaZviyaddAaCKln1yYeLVoZ
FzSELv85qQwTRIxdPB95fPSDPTyE2v8orNE4HMVhLspTQofXwvfnxaU4V7fvl6sh
hmnzSbMkKooO6Wqo6mi/ls3c7tECt1mKq203I4HNYE2a4i5vS8LaF8zDZfad8l22
0HUvbKAbe/8uFGsrPceIpZf+UDMfCUpeJ0079B08DDnU5Lglb69FvFMKDp0AuKl1
/Amv5yEDN6ZG2hP++6mCWcKO2Kf35irJYTFDCarOQNQ6/VOUAu0nLOnpD8V0oVSZ
y7D6wIjVzNJs7gQAY4ipN6gSYVI/E+EKdgWWHVT9HYEfYoxNovRKPYg/U1nqjrc1
RKAS+msIRjgW6Zm6+39X68uN0Pnn52vz1C2n3l7C7JJ+0nSz277t9jeOyGdjky1K
fb84NcUQaKO7iZiD76DLiU6xiEGcrYw2gVWdiKZTnwLhBnvS0ZmXsyILbyX/xUwB
5KlNBbWbUcUZS2lluwiKkFA7dTPILR7b50C5Fgmq0ol/TL2WGy+hI9d7Q+Xbe+s2
xDdBIQzyGprUikRzXolgSdG9ZcGruE5XwWM7PNjZedhxCEQjIxh3i2fYuJ+ODwG7
M2nAnxXaOS+f3pi3b2/LRHwc/CHdm5Pa3tsJr4LDCunxGg9Xk8YoBB2gxo9thC0c
/EZwJeIN8ew8F4vEr8qOmNkMAqZ+TdpwKSK819BAPmQpLWA53wJai458cP8eJG2Y
UaXxNbW3c4PynIy8AwCbPinGmo6YXmcTZlkhJKsibqc8CQYlxUmd7N+5h0jvzxKx
fycLfrUC+W9nDl0Kmum8DBUux5clgRGQxz+BDkHHMjhWoP7WctnANY/FV/GkoLRp
/Ue7l639esTbS+hqCfF2TfACuGRTAyTFrzG1ItyylLQUB8polm9kuJP9Jq8qDU2K
bmDS1I0ihhxVE9Vm/wgq/Em/0U00NQ1I1oi+rH/CnoHXQQAg0BxXYgJxZZSTagD0
0V/p9iZosrsYCrkzdPgtFNph/vxOQ/t4189WGUlRZuufPWkxIhg2PpgKaePO9nP8
xhQotnOAvzW6U1hcGQ/aefebt+jp1JSJttNq82YhVVs/7pKQ0iUbCKrwN/aI1ruQ
gt+L9HSuXrh2WJoIWExpDNzdUp1mFMwJpflLx1rpwURguIDYVSVVycWkxfIZHmPQ
VCs6dNy8UcQxGNgM0pTKwq/kgIaHlvUBcyr2g7mrDPaLww8C/GL2fuFGBq7kSr8n
o9GMKQlAfKW3wflviMPk43qnTSJWDaXm+iPcgv2cyN9ilUd+81n+kTH4LtAsQ4qV
K0CKALvMqJhgB0M2n5wYGwNHG8ckuJc06+bOl8I7eHcM1rYkKml7NX+Il4SY8T1K
MCkQZ+MoioQ03YykQ6rwsjbC0bQWr+GUaFdCO04SJPnCDYsZgRnsy/JLEl7Pu6Vz
xvpDLHsAPOwv8N+u94O3AhsGa2uWBTDdE95P/aevA4nweoFpOB36mCoV1X8fyMZd
Nv3++qHDsXnCKK1XYW6LCs1KXt1ZaFp21SqCTuMaS1yrXiURtnDiyM+y/0+s34dP
PLJX3aT8Ygis0SRNF2eqckbHOFvE46TbRPelCc5gL+U8e8/loWJCCdIYjjaWjEuD
GUaquFgzTxiKaaqyMNzirOSKlx9GE/9npnmLZjF0Tux4MqPEuVssD/jxACaSFIN0
XVTWR6mZvPCYAPI1Zb4UrWxUcPcGebyhTRNENX+0XtJykNS45Vld/Hl8fTqpWKwF
aQMXtmYRtv/RoLXjxwWs+x3814e4ZpdJfVw7z7EujLQGO+g+MwbIEBAEcyfB1c/6
v0Vp/aECplqvBD19+fDKh6NwuMkxDum1fn3FbI9j0x5usl9nIR0iZhbd1/vq1O8C
H9TkmxQVPv/Fov3opliBJmjJQlM0P5FtI14tIDwskexbTVEyLcoa3npgBVpRrJNQ
Zi3G3CEL2obMLOGA5Jo4Rp2b8NmLr4OHMLcUoejZ2aQoVPIXmytDAqk8YBN+BCBi
nnMBtiKsM1HpXt0H1b1SiOH3giZSGfZi+MHt8VquIc9B2YojxYx+h9ekK7VkjT3F
APg+fkrwOwxmIKshLLCt53NCXtO61m3LIcm58TpxzABCx4Xt7MSjb3lgndZROcHJ
2KXx3lsHvTmCEaid5lAiOFV+KzMWpyjNibvK1goUOSBQWLerIKS2Ox/MWdql2LE3
bfUTDSh3IlOWAWPwugQJxTg80nSfXRce4hv+Bcuv+bumbvMOqo88mVG8m6LPmFSJ
WjphOr4zBFe/gYv1qI1eWNHVJiW5UY7W+f5x7kgTL0E+O6mB4Oe+QCKNMthXQTwh
3/cmSthXVbMnhgbG0jPgkXThSE5YEFE7XrvxSwzVzfUu5UjMTM51m9Ih67B9Jyay
iBQSewmdrYANjnmHtjEofPXU4Wr5b21xaApT5hyDw/b6yFMMYLq8tPurFI33bYne
/FfThRMDZ3wolQL0P9GsFHwrjfToYflCbtEPiBLOQC+dCPc6QNpfX2tAAgCDA1Vu
pzkR1BPwIY5gWEzR7BmFPG1ELZ91LFsX9kgLQBUJ+A8n1QF3GVF5P65Rik3Qvp0T
mLMOavu0K9rguVrITKUimqYdM0rswoRCVPjgp3hL25VrIVbDlLKJ8JuXN+SKWOUt
RdnWlTRNNrM3noMl/4Nx9K+vt6lpWn4S2drhoEU6facHYgBHQhgRXN66ZV00vjxk
zXyW99yCIZeI5Emy8Ps3lRdfukmtb5sDIL3nWaSkh0dwZGDkqy+DqC9RY6dIlQvS
rbOVjGLPNqce2Tm9IHwXPF6Q40b9zGX40F56+GRd5rRe9c4HnGrFhdXs/ip8xPeN
Pb77ZsJ1o7bf3wPt9C5aXc9fyo4YYsFYvhKDayEqy2ga/X2mT3hDiTzKWO84fwiG
KVwuDc1hkiDNMlyH6AcdMOTz6ahIGLSBX1+fcrFwiW79sHvlBmESbfJHrdV62RPz
Ck7tPQimro5hVcZmVdY3pYgh2ix2FWGwQ2h3UvcXQjM51l8DnW0JYZzwMYHOyx+S
Uml0oaBcR4SqgZ1Y742MLfAeZuIkRKcEIafgvT0Rkt+PQIr1xDwZvHM+uv33nrky
t1ut0vnPOdWKOTlwR5ZXdQfrQ+S2mQ+Vd8GEUVUvnnYke8IJoWQqXwkWTS3zj4Xg
yxr0Ald/ObgYc8hQLOPNLn7Clni12aeZz9sOAgJWuouEcl2t88RfJ6nyJKVtUrjv
NPSHuvX9J1k+QJeRARdNcOdPOqbMuoZ5dN/dzNE0tPz0oT/2ur8tEY4/DhjLQLlb
M5H0o7UmUEuR1bPs/XVJJfoy/K0GjBm2NYUZk+MPHX6W43gEnvAEB/Nn/F7Oay95
PzyQU+TLnteA6KFgswa95v80NM6mI61nH6TEo+X6cjAbqDLN9gFtWcr/zh7qou3k
3Sa/39FOuuP8ei4IrhL6j88s0yviXR4iBKDZp67lnAUGKHNMRgmkGa482a1p91x8
aREJjS+t3YOrk7e+X1v2tQBoDo4GzQkdNvArkuW05jLDnLRBx+1tfzeD5k2MGwIz
ZD+dclQq+GuYlVQfzmq64GLfy9MLGeK0iumQpoCtBNe1KaMMe8vexfU09RX/hN3B
Navw2xyJALs3RfroWlph+eZTxcRLE4K1vMiHvVWjA71P3FoNnC/SOkkDCWbwNRHy
Ct3ljV11MIXLkbN6uzap4UmWOTYCXyEuaJJ11vDj378OXQW48mPQ1LINXMuYwDpT
cCLBq3WINVrhH7ar94eyiRkoeZP4LFzCwEgM1K5UP6XV8vTyKxOb+y0Uz7JxcnPZ
/rbrbvUdL3sDgQxDVGf86AXenCkhBlizcWVCNlop5K+9vMAxU3evEAAC+EU9gJ3p
j0+S5xqK8xRpH1fH31C7t60gpb0N+6n1CeReeZnT5bLC8gxSJdA+kPcxIeKgH/kt
ovmTck+jP6UDJ+9eM0q/S/RqBPnJYNW26/7SQHj9aNh01cTviXOyH68ANPOJA3ez
ABsNZo++8VLBQ8CFimE0uc3QCXlXW6HRJ8+EN32fyF6uxNH69ii03cy29/C+Eomj
t1eUEU/SBLGYX6jfwhxtL2Aa6+PBNmlq16MHdVzdaMgd/Y1CWw6MmZm52VeJnltY
l5lwdWpShQ8M/PXEQftWX2QUktWdMQaxUFzscaV3TPzkc12WRS/jAu1nhHqVTVWk
wA5eEJ7e/JERWq/uyhiXJGr7SJrL2g/5WFZ5bJHaSXtWVo9b2gn5WMmYPH2T+IfV
7Fl/le23L/kvZ+CQ2x4vRm8eHIR+B4LgUc7erqc4RL9BsOXtNAn6jQ5BAMyLp66O
hkxOqvQIR5I4s8ZbfFOgv7/uAbjCoK8QFMs+JdqZxRzF8A//f9MQ5NDw4MjfSVhc
W4F5slCHqzd5l8+k8nY0NuuwujM55IM4rgFFWG0GXzZJprdK+iOtQ1jPm22oGsGx
npy8LdxMaGyvF+6b2FpDYjTIfECdJ2nJf0yCbtrwjoljt1eiC758Td5j5MWqX2S5
IIAefCeBkBHVzpBy9Hn1q3Phpjq1iXG9PsnP9MCjfAAYbxe1vHGeDRPRs3auEHI5
MmJazu1fz0MdSQF6gndMBRmBjHm8BCuBJYGo0T1ugwAo0xQ5/Xqn7OQHFN0OOTOq
CMSnXO1z8ZGgWszxyOt1AFxJM6CY6bXB3rEtWydW4yrSjqDOVwHl62aI+jFRngbY
ouxoVPnkbPnIPh4k40FViPUYQ4cEK5exfVv8c/qUhbJWW7elcVTx6PVcspCTKPAF
KuwwwqOJ5xUdujiGNkefL7K4KktZC+s+AsqdHPGeZM50uIGzte5JlUnbDltve7qz
gsZDCKUAPB1Zng5UrA6lIo4noRl2ZWHlSBSEcDOkUcciaIo19uZ+x03e6nHJpUGZ
Nznh2fJaVe7LlDZO7xa/dGa3U3aOitLpypscdv47g0d3haS5m9JmArOcCabTep9s
vC60VfeOxI3PbuEQFTZNxSpYeNcf7jf/v/pr5zOnM5OoPwxmgTuFQVQV0pmhM9TW
XuIV/XLO2akwOXXy9bO+QAdyuCZ7mIUMBM0zEf5HTNLjKtevaIFEpB6p6vpBYPtx
hjRZj63FRHk8aZMwCCVXqZienmvuycYu089xGOXawVcmY9CbJ3Bup4+Ck5sM4rzP
1bOS6+N3VdzEpXvr7qLTJNRwGAtoeBArKPw/Ql9GNQ1eI1AxAbvNEU9P3DqROYEP
ItnwAStJshDXlKH4V1xroR2N4vVuU9DH45FxUMOqWXGQXaDlXYdB+IcrbCGYrp8p
v4FWGsEUjgM8XIZ7wi0lvVpDIYyqi04jGf7yQGsqYMq3bM1x1M9g9GYI4NRwF8OB
G9V6pqi0NUPS9ZGe4l0bgHh+gobX38o8oxDWAywHu+V3ceFMcwiEFTJS6yXNeWwx
rkptp+cZAsfp/p27W1+DgyYg8haH8OSj0XM2l/YF7C9W8KymxX3Dzm/RnlHsx0OG
xBAQjC8+8HuUM8SmCbufhYvDVztDZYR8knyzY4usNyfHQIFonCVEOGvfNn5RCoHQ
lghvMTFTMzasqIBdVkXtdESPqj06WW1/kymUwGZo1JP4bHAsksLjVNS6VKRQeNob
jNYoE1F12Qdq6mZ4+1Gtth0vRYhGt1hMvL4Je9UraK6mozkEqMfQKDYRymB2Z48Z
/mj93jjYTQmIIKW8W7E8y/8dd0rCDJ3Ne8rYFE/XhLSrsm1dsdFMpQ0Mh2Z/Jovs
D++dh5eWU3ABzfXFFnnBcRk9ySsbZ2pE+bFR/HKWyU8VEslpMYleebS4Vpsa/Yqx
RPGBRTmdkb/+FoI3O/QNcnP+2M1KHnKCcQWmV9sfwOiO5Sno5S+T9QrfxnalRFsj
cITjahJG0up+W7DJdKgNeNi7SxMHU5AbhCMeNOkO2KRGXFrioHi3oUl2YeXNNnqf
oJzYKKSotGGLwROQdjRlmVHX8ZU0HhFe5UzGXuLmAapBhMxWzPhQjWnOs/5ChfbB
EYmD/w+k6BNTMOswnApegTlGI71Uk2Z7GmypjXhyAWrqVIYUV28UG4KEQqv0wVEH
Sz8kqHtwqRo+n7T4Rgcs0EjC7QWo91yXQdcoU6ws8NxZHB4Pm7aX08B4aEc91c8g
8TncwOUdt1CDFfJe8sH+nghnAxsphnMOl+SpJOLZdghGr4DxGlXI4uICocxzK/TA
X1mOoKGxDYZ39ttZo1T8O4P9OoJIrtbjFQF+r38rwZvMrul05l/mxS7Hi66A34PA
5qqO8uXN+MZsCfnMfpy3wI2gdsTUL3vZgMcvsFLb+sht4xVDPj7Fp5q3OjqwT/ay
UBxFwq7lmz5F1AXEpMLknsHZYfUb/mkV2lmmNYWFdbL+6qY9cYNHzS8mz7b932LB
jPSjWp98tDIPQteVOFR1+h4vKN8bkQn+uwVzHOnG7ALd+OrS2zuQ00DhCz4YQbf8
lxqH3YnVIOe1PvoHPVuDsz5KlJx3n68mGbJlqkkKCvnusQE2xeKvkrSjP9TaFRLR
2K45e6kWJmaSfMH0dwlh1C6HA5keM1mfay0osl8K9TppwLIdVKVIs3P7+I+IlSwe
ac49gxupcLjnvvdGMOMB3xcttkw2rrVtK0NH5lSKjbJdOdoK9QjlivRnloBCAWg5
vS4lzpGQ0uvRzA5GpYeor4xlVMxdcr1Bg4ucOEMJSLpjWt6bpI+OPtFZHbhb8Isj
oi80RVPObOQOduTdwRs7X1xHOcwk1cev2h6rrKKMtKS1nEQRKucrJ1SSka8o93bq
BrWsbAuHPm8/zsjyWpNDpMiayKFck5v/eYrdjTSKO9De6h9dVi6vE1cmagZcWWVN
rwVVhCD1BFNdtoa+aCNe9psGW76g9KLtItEcoXBGnlHrWx7QEoT4jKZkN9aPADgy
tEZ9dMUvsfdC+TMQ2g3Dnrxnxi+6D/WnqDn+euwlbZvpSHydyV6Hbt48jrwOb2Oi
jxrbIhbY/lhHhTim71gUXRye77BEpfGMQ2wAOtaXI2b1A1i45afCxnQIyiYxVw8L
7imJ/RGdEBcVncmZsxqUeWxWI0n1OOKHh6qIVEVVfMQhewrIm2NkSFsPQeOHWuWq
XTA8m61ETFk5++RcHmteOUOcqih9lnZDuk5J9H2R6RaHXRsgR0c0KRW7rpRZA5Ox
CNEHlylEzvUxN3hKYVWBQW6guK1fB9q4x7a1D0MDuCw7D3w2SH2zHa0lSOQw+CCA
wbGswRR5QUsDXFPj7GjO7+8+Ta7z539oWcGwa/TduGxENao+rye2JL55zu3Xqt1u
FTY3gwnDGEVi1AYF+VjCXmJobrGN2qV7lr31v7zbyCEegdBxz/CsQEKWG317EwMb
Q/5l3l9+rjSHxXyFT6qlZUYIuL7OfUgO54yp1JtNI6Cc1Ivs1C3kHuuMgeGousMs
eL+gPFaAxEJ2tB7CMxmuzwBil/q3fTlltGVx471uFZahqMRGN99DAbpZ/W1PS6fM
YGftkSQ+UT34KzBqyF0I9pw0ypO9p7K4hUQgP0MwBqtnMe+gZw0J5pmGDWnaV2yZ
XZX/nYQOHj+L9eEiweVSzgIEqeBxlxyyHJPLGg9FcNvORxXX7xA2GECo9Rp7veQ7
w9dKn3u11QhoJ/bFSGDf4uqH/3F5HzlTpNWnVO3H8H5BKJksCdogN71XfgjVl3tp
sEr+ElE542Jyxl6wzEivW3cordDyNe9yCRebrj9ueFIBuym93qvGAOXBzSmmvCvD
UpeezknNAq+p9vcng1uPvlS5nrMwU0JRnvfJF3Yl1JPepQN7i56O+GNe91iQzkAV
Q1NSZk2PewwEFnjqZxVZNO2vGogrsUrZpuy4EGiBl4SBVjFC8iAcsNsbZQgF1ekR
RYkjyl7LWx3z9eZsqQ8NTBgXlBWTuQvbYe2nSNsS+HhOiUABCWbIQL/77p51HRF2
2cl4csHpF17ji7ol+R3EFafFxo5WQIpk7XZV+oWQ6LEIHufjL6sE9O+YzqkEOYTs
eJRU8MYBiM6Oh/xHvf76qrAMq0rk0dqlTDa+e9buX0bC0VKDYJrXH0Rrgg8XixDr
gtisTO/gP8LG8aGVnGKfKzyvJfwsYombKjH4QZLBJW7h3l9rXzjuEwxUR+g7KpeR
CIwKDbJdGulW5MgijznS6GXIjBPLdOoDQLtkQdp4NOpEmFGoW2JQUXJ64QlBneB3
NQFm5gtZrmnFgCHjcjaNo25Lgwh6S30RYXq6Mp9IS+nW1CqJj/zUYWTOQaqTNfyi
4in4XQDwwzlJcYSVwOX6YgjKEyvGiEq7WsTCq0OB7Y2tFPZNTY88YXoM7kqKQxHp
M/WPIp4vwS85vz7tFKSLabF9L5/UdYLhhCW98eswM3Z6LgLH1eYnq5F9gjIvB4ny
+vFmGBEtQQ4M4n9x8Z9ex7FEEGdAMdX8TstCNWgYPzGQ813aReTmg4L/MB5WewwZ
LjPSRALKTcbrtM93vOsIOg2h2noJ9ALX3IZad29ybNBFc7NN0P7D10XPRTAdxyZv
Oj5gopKdxuNYJVmVB99bU/hgE4hYWODvYyw9f+n7haIofPrHl9QY/jorv4UzacDB
yQOEeHTH/h9ZQCbhM4kkQnqjlYbbwh+YhqZh0XyzrCx7A9St88yA20hW+Egr9+s7
lBwh84BunWMu1NBJyLFpZdHupE/OLTDMo1VMwUUndhdeRjvCSJlcNM/++6OMlavb
139+GBJ3IsGyeT/ev5X+rYLw2TvcEymMrl4F7Tll1h+cpmv06HwQMiEMjuyIlA0g
B21wrXD7Dc0rFdw0VCUHIZACAQGdpnC6+AuW+afFUjiQVVvkOWb5x2WvrSXSd8h3
D2ex/Zcxh2AV0v9iF287MXCFpYxSm3ceK5hohHwJKruAtZrlEumtWKHLT6FirAo4
4KMY9qk5KR5Rq5WYEEyLGUJYcv7WI6cvi35P/apIsM1zZDK442fPBADD6DH295fg
RJvuIOkJKfd9BaSZq2NDkVSKqBWfP41lDBi6lTDxhi1q/zHZk8SHyRfWOVkTX/vK
zk1X7luaEwb+40AZL2MNatAJAGu0aEG64ayQjqOqf6ORjGhfcp9N/J9Pnga4IRHE
52XeT7bCNjif/2p7ltL/xotdhPWX76B7DTft3RBmPDMNDxg2OFrzKaBSdbxvt6Ov
TjUj2vc+QoVk4LV6gKHGFkdwm0zadCmI/T9SQ4E8hl+5bC/Mdbv3PLbsjjQ20gOT
vPJrHMnrZq5Dcjg90bRwTIaFanpahCVkDhnYYj08+lJrkptK0V205nGS+TAdaZtL
2YQ6buydt+XUhi2d6xv42UooPbmmsC0WLKtOhrv58Qo7G+VigmdHL20WCgBnah4q
VeGBHrJyplrYGAUQBEXDD4x+C1gCAZZP/y7i2afCzDRJFUO0nlb00fVF4Esb548F
lr9YCXat0WhE6HqyVCBFPP+DG7qZribr3LYfosQ8h3Vct4TvCgneTXqmpmZbmLeL
+jWKK1LxHIv3edLJ+Pp9ESB1TKb0FZgKxccWNwZlgDr65dsJ4SVvDg+ya3osQVxr
YVbf05oSaMaAHoWkjKj39BsMn9NSU8qVCsvHyzCSlvH44n2rU8CYHwIeeKNnp9+3
kVn4UrnpcbzvJXN7nUPiBs8Lmxye2uRq8Z24mMP13pwzEGVDBu/YoolqIO/YO/7K
geA9p/agTtF+zo1KTcaopRGemFtyeed90Yo8BwIdf/dzTsInci2LmPYZKtvmo6PD
mPiIfC7pcK4zwYyJfkwPsmA20K6nWKub7gqC4LY3PUIUs4LoMX7667SBhE8z+mC0
Td3UWNDF6qHV9b+2DtFm5KOdeV9rL9QYhAQ/hjC/e8/S5homQKKyFLDkPkGi1SPb
AQ8ra1+o8BjHfV8GylwAcMJvb5MmA5+JbORQH/LckTvY2YqvvMCe28pbKMruWMwt
Iv5hPuTP31AJpuM0JnIhR+ZbmbICTTzllUy24u4prar3ME98eyeNrLdrI7En9GP6
3j5Uu+37WvFvDNu5WX4ha4IbRjwgOAvVBeXaHQPVFFKNWB3LlTjMSSptP9DUvTlZ
bgL54O4hWAxGZNQEeBGw7iqPP1J+8Cn6r0hTi4x7e8+egLgRFxOiVVW5rp9l828i
CKuXiXW2iICdPxihhK/Q63z6oaT6/XJlg99H2RICFpRTnSWB7HvSGuwRlDolqwjs
mWa9q9Jj0lo1CstamZkG9FFyUMgjJEA0Mu1+vll4dJZR5VicwBXxIOB2Cz60yCml
cMuxwjuZYuXVkrm/KeSz7XLb+Ew3ZCoC3IZdwpRkPGg22POgGSZbQ2Hi/k5MUURg
voBJgwfaTrYLdl5ye/woUGEgHIN+mdo49DpP/q5Og6fP89dyQjYzagC3/UUDRZGQ
Wr8KN5JBdfmiWCS7cHcUnH/W4tkogzVEhypO4QHyYBzFmF9GrwYwPfxoz49/4c43
fuivGhg109mv6AOwOHCwTIfINIvJfJe/xmLJzIcaOI+2gHY5XBYugvvL2Y7IuMTJ
Nrfzi4iioMbBrtfmdSeLOnfJA3/aezRiS9nfOHL6CLno6lv4Nn0oIv5t1go/6YII
RYphw/Lx/T0KBxSB5gbbCKgXcnLnVudbo5Foy96rmBWiq1TZwXmkaaYqr/HCrsh+
sr1pgs14KSlap7KhhgZnNKP+fBVbpDgzW3vw4Mhiz9oBaqgC/CHEbGP1DJeNHfF2
b6RonUtJKTbwsSOi7K6GTjE7Mq0idmEzv18uyRND4KwkqOJGyoEI0KnPT5iuH5El
3ZF0nwv/Wjrhj+jeFR15ntlx3agKvLk5b+DRQOirFai/z6lPQljoXgmSX/HgdYt0
Dnsr2wS0hwZgW/2xlrapr0cgkvav06zJp1h+fDxB53JUlJeHCQ7/PPnsOHVvqPWM
khdTdUrniU2O+ALWTelJYZ+H64B9UfOm0op3F7H9K49RJXiSE2fPWU59W6OTDWkG
NE0RuNfUHjgLnuhQ3aHKU3w/m+rFisc55gjz1oX1MRBXz3wijjkd648eF5n5EP1z
Ze0lT+Apu1wRmZH+tDNyE6dkkuBHG4HMiIJi8LymZQVt6nCCmG46wfX3AHC7Svb9
yQwnzEYYOu4IyP99QxI4TtwNLUevMlvRpy138/VngmaU8p+grMOkF2B5Fzy2W8So
NJvJHYQfzra+7WiOSJQbeuuxWa22/nuGIMcrOLIITlgUWRsjou4Dm5qr7yr7aFDT
CrEfo0y2CSd9geDO4DCAXE/2X/IwJSYQdDKEdJb+LFXlVMvJ0WuESNNPuTOTqyos
pDIH616oxynTsrPUDkPSW1BIQ4kcv40J46IcBdaUz6tYXyh/fR6vcZarqSkLljiX
+mmXG16ABaiF5agvdZ+Py6PXDhMz22b26EzU6MylZ6h5T7TpGU0SUAWwOreTbX6K
PRDq9yguHSeyZqL7w8vuV4PixDTHS04jBUfL+yr5eD2t+vKAhSNls4K6fD5m/x0D
nZ0txfgHHqfrZGTSoocofnO329ecwUT7QojHIEWr/jpDAA+oohkuCUinaRPm+6KQ
Hs+XgMKo20f3BfPlOIZe0d2J0z7o+/S50y7iLjSckx0Sh0XbHYR3oX8+SYEXxJuP
7xA5IAysSOSXnpzl+CtWg1FOy6QSXSUQl1gVeX+WbXVk8cVHcC+Cb/SrdS6QUuuq
RIFkBVAuLd5wElbXYmXZDtX4I6L/WIyWRpdQaZJIcnEAMPXb1veH2MmQLk0fCv6q
muyTkRzna1MZAZHPEJAvAg36HFu6LgQYGZJWn/vH7SmgLCIWtbOGoEWi6+8adww/
/vEq62KgXGhtDkC92xADx24kUS/Ur8RzzmOz2Vle7htx256rynxjyv1cfPF+mC2O
QTvYNH+0BLMNfWCnd1E4mzMJd9JS/R7VRFKw5cCaY6d4xwhDOe9sYn0lp/23Cea6
tu9wU4Esb+diBBASHavCKiwAzDwsKbeoUpgVDAGrUrwml4AKGg6cZ4MQgGe0IOW+
oAfz3Z4WvqLYu63NbpO4vGbYUN73LmRrmDP+LobI8EGH8/Ee/8wukVaslWvVrVmE
SMC8WtL8CUbYbn0wlDmMAFeZCAa7N1n7QaZ95+iEr+a4pDY2zfIzx1cGLypK2BXP
y0Vf02VdYI/kZvwYkllmN6BAWWT0VECELRTIv8etK3kXvWS2QW5Hwyk9QwozWyBm
zNL+VbdNw5TTUHsV18AoFCkZEVHPaHHJsyqa+UlDDPv/dNTGDUtSkXcIy90ubDyH
w9vRlJLVIl1KvJlQogHSoCUZIfrEsZ30Q+4sTCXXNaKqspmjHSvhxCaXuXMsPrDi
ESVWm99sJo+mGB+2M7xFO2VwzGoBIE/KeOwQdYkNdanQ5ITZrzq6KDKUo4NjK5F1
zRYvF+I8Uhkk3tcIfqA5O5teQoT23LYvXRsIVH1yhVMCWK4B0OJchRUGsG4YCxI8
4vhuDlsdE9OGOhcBLCDjn+8AI8veYcHe/1xzlS+2maczNX049bDDNFS6pjUtE2a+
u6VVxMTqUHXAGhbxfKWgMehlzhAGEBbcFE4kfmVe6qrcmZ30X7ks9rV48KQEsC+k
HT5+p/5hZ+U50aG+LijDOSGkdLrCzJtIgRVNXOB9yovdaP+0CVZD8pYamyW4dCK1
mPaz79+NCMxpxkay5HS4jUscTyEokzlXSrCcGut2V5ielgMvXAdI1u7oh2m5GCdc
yEfvUzaYAY3hxkLgFyK3ZAb1qZDyIQYXUNT0LckDD3N85t/jPbslQSDmledtWqCm
zML2ME2iBz3qDhVWH/Q7kvoPJgZD79t0bOOuupKIkNDIGcZv1GSOz0hB7u+mSHPF
5hN0sG977J4n9K7MupBAYXdGDL9XW5JDkWsc6lBfdEDtuDmQ3+cHZu0v891nSUTa
d2Q6VeTB+NNL1aoxQJMzq9JiKuF8dixsTBmYK5TeNCDIeyjHzrxU0q1VEOXE0qnX
eEYQYqzWSWu5jNkC4m1njIiGN+37Uz2bVNtdhtpCtYD5tU0kvlbfsfaFhV2A5xWk
aYiLYADX5XywWUJ+miBCAZh9Xx9MsvohB6ZOrij1sE9WzG3IojO2WAAyuAU+27j8
H1JlnDAWTprNwEtbLiLa5hpNcVfYeYcCfEdlodJ6IRm8oQcMUjLfBKvsUzT5g+Tz
4WlhWvdw3RmnFnKzWnYhmBYaVd88IVP0a0KPnkOa24hoZjqplUgkW4YNW93clIzI
zLrnTT5g9tF/qQJz2Nz8PNP1TO/3uYSQTIzwF8p6jub0ivVYh2ic2YOsm8XWuBmO
NGN/GwDxdkOecrQU8h1EawZaPuZKHOu4lCcQ10SHvWFH15ZychPfsYeHCjg8oWtO
36S8XoSBjhWwCu/c3VpS8IWRTHaAK12s2drMeXa500cfiP+HZD3aceoAIIy6R66r
b2O0jEdcx3mNhTIoPd+mrewBMIyinvAOeUDrjNMtMsK2gXOBr1/E5UqN1cV74upA
Ickf9T0e1ZHO4/sm3ryFkU7cok/kPuCuaSZi9Gz06hTq476vDBBhcMTuw/x5ZYIf
TX36Zc4bdrzJZaAp2VUAVCTCaCcxv5bfnEJ7WeTavY9IWpjDhS/2DQQFZahUI+a1
SkXrSObtAGaHBBh1cEbMIUCSRJZo2eCMksGBP3VtLzitM2k/JbDV3zIFAHpFbsKd
mIlixkvt6IN/PCZmUJiOxZatmmoS6vKpUprG6hWm0rBickTt0zwHjeuRx6l+7yDN
X+EAgXu4zXV9uFGtllCkocNJNbIyvJj9+Gz78iQuUL4YsKKxcujN6AopV2JNxzBw
F0CHqplJVfO4XtCy3lNxo3Lg62q7v0kk5BZCSkQc64kk2Do6ihps61pMwR6WWh1a
rdbqUso558/yt33RYCKNTHeExWT3wLvNsWGtCqqphbh0CPgjKS1JxMumrpi2WfjI
sn5jZOrQnAjRfe8LF1vlhPJQTo1woqb7K/XQWjGof/5uzDw2xFUBn1s1rXWs8MHb
B3kpHqoZU++YXynHNp5FiKBpat3pN0SG0EQSF060Am+RoEwlVMq8jW4VTSUnobEw
Rae2nqYkcdXo5UDV0bdxUKjMIcp4WcOCFKMKOm/Ouq7EeL+zcvh24K9MvmyVwp0s
2OAtyAOH40LyH3CZCJJDzcP3CNTVnFW7DlfSR73vgBPdkbymC06DGDV2icSaO3ws
F9YMHOZSLuEZBhbsjk9mOAwuRiaBeLJWpzsgCZJaGGzn3GWagUrUUSpnGcqEvcNZ
ljIH3YPcRQk6FOP830a0++IR3cbA0q5BIFn5i6wI7n0TUAPzxo3596cF2bYj6NuA
sWGk4uuxUHzw2eWMiwvwOcJFNl5iJwAeY15DhwreYtLPA/fmuEB3s/0t+veJ0LLI
rsT7QORbmfmBYHszujucnDv/oEmeCA6nMlHuZpNRw3H2MJvNTrCnxGkL3JdI8nfK
aOZPWff4oklGSe4M668P689h0ZGUYEAqJH6zzF2uxHVvuxcKFB8RfLkv2yWjLKzx
NMAm3DLBrYNmsQun1DWGOzgyX1Mr93mJb3idCYYod2fxXLyE8gNIBxpSsxSkRbP/
HZMyEzT9I/IXVI0wsVoBhTs06odjeex6AVf5srfXNBTgdzdOZXTG42Y/K1Yx7ntD
9k3Glb9sNEdfv4ItOFykDQkR//uYbxRDkcqsQtMg0iDZkgTaak6JMuUiGkraMh86
H9kSHumdaxMSI7kekrBMXI9JStEdCzoDAdRy2xV/eyoo0/vfGRSPiL2YF4E4YKYv
fCO3NjC2StgD/VB687Jr7ICefXQWDd80p8IK5DIBCT16aIGPekWDJFEUbbKAVVLS
tc6wYeuWMUwtmnmh07NOaU/Ny7GCuf7s0VpPoKQlBLilIYIuz/ddV8H9iiN/p6Ly
H9OHT0GL/G1GEteMOmsckMgWuanlVougawdcOfCz6rd2rjob8AljdLEBcJ4AebOJ
06FBv29mwpem2ol1GSTmAZB+eexZXTeeYR70/pX+Wbg6jXmNdg1DOnqR+eaMU866
Cv4VzfPfrN80msi0vh+DQDzhUS5eqJnGLt4Llqct5RL6JQ+fax67cgWWH5tqaoDS
imwYxA29aclF7DMZwJklaSxVk8apgL/w1/8GaTJmh9Y9SKRwHOc1vOau1UzI76vh
GLDnP74ECIGBjMekh3w0rUXHj/sL4Z7w5vhq4aYpUK3ozTA3nmGz+z8X6vBmG6f2
eJbuT6OM/bP5NEjEaE3hRDMmja4Te8ehsKzVe8wIcEqXAxPLGSJrOQavgqpMoBlP
0syGFs4wtzdrJJLz9xOI+EHxCKLpBDUbg2O90nEVRZ16lIzgpMBJLJBgCbDihIdq
2xONxVajxuuXjav7PEHhdBDE3hA0m34meo3ixLUwyjTBcq5LFcJHMMYzkqd1CyY/
CRnCGLovFBqbm714MhkDS9NFtXmnFJO4Yg6GFRwH0hcx7qB5sohoZx0NhGuRDRqE
jA6q25kwvlzO2F8s7HgbOAS5KJaWEg+0qVJVXNmkKWLsrxyc6QJYGOoZb60yb/Xz
Xqul1QGQpW5TQVchM24s6Xui+Q1YK2F75WX8eXrkDJdfahEICB3tHj8AXgFkKgGT
UX+UAPco+HY+OzO5/RZI/mOIIRd8MyNAfNtZZSU4k6IlML+hqsXGCiyCtUYUAekV
jWsm+bsQHxDM4hetcH4POqjETgpmhtB5wvRIL+q2PZHK329THK04qSxj6YXHEm4E
C0WfX4tFDvuUCOC+qxWFormPtUcYVWXzaEj4xDmO9EDWhbWECz8X15aDXiEbZBuU
2sKNKS5ynWt0yYhDhDEaEN3xT0bhsnsKOb+11Z4WzExXgfTRXiCavwWVUpZH28AU
O1Duk57f6i6CSauYLGUL+E3ZKwhQcWrTPkOVNGSFav7gDa39o4RuIGWyji3nUTWL
kXp4Oeo+brBXzLapTMrwR0IKmy4u0+MVq7oM5dXytqYzZyGdc1bIcP/dUod0PlRS
DDsm5oEdi4awfyFFWy26gLIo9vUjb14HB9hclv6JySm3IHVfwZlHlYHnRi/qmDbG
03PYW0s+sBYnIhlemjhTwYhGKh6cnnEmw0LEOGyR8qVbi2QQ3u8ADYBkROAsta3R
awdJszPhb1vizI9WY3HNRdru9VVTqTOHagrznL6FaKZqxQqO0F8VI+CrAIcNUUHN
udUaEKiPEsQhx4IHAJi+XMnajMpNlZgQ8Wof+0H/2MYgjd7q8UZSH2zC4v5yNeju
JspUabGRODfeg8viqv/pTTE+4OPRB/Y+2LuxLBBsY5+5/SsJS6Spw0M9ekkwK/++
/Ds98r9mhmMLVWIi7Aj3z4IygLmlUgt5iLRQ4VtlnnohJAMYZRhKVIyRUx3dxJFZ
1O1BaYzMe/1VYvWpyDWQ46wAa36xQk3Y9YjIgdC8jhCyEFcX/B/zR57SihT3RYq/
FPvrD4W8uP9OInA+08QDwJnQGA4v8uEvchKO0JejH801hEWlW4aNZMfgZaL7SmXG
OIo5RWcAvqZdhG8bq9MEuVogCjCktCM1Ps+kEzkkz2O3ocxW+BG+MGjvMMJxlG2o
9pI6qEJdxcJA7iM7yEV4PqppNiipLQ2NO0DDO2ZUcUGRXD+CWBQxRUDXAAwc7vIu
NNEwO6sgoG53a6I9VofXW8qDXIawPRTCBjhyLsKnH0JN/YnbYfIDCacy+soSIkiI
xD1HK6SF6Or24y172sshv0ltZJzYsYIHLBKeqp5PhzT97r6+lbLdnR+VWQqQ0uNl
b8AK6LC97krUwuaFhy6cBKvgdzJeH8JrdwtOTJUnoj/V8hpD9q6IhBUOH/PmjmPG
EZMve5eh0KMH2S9vUQVGPCLewyaa0JO05SRU/aU4X+nMS4AGj7E9Y5UrVPERZJeG
I17pRTK2fAySd9XpEDSkENLTI8fKujEvXnRjE5VlLUQRit1JAuLKVzFl1Njn0jMC
IwxDhiw8zNkeIZ7YeqM4Pdami6qoh2x+3GcDMfGfqRTWwVEUB0zi0Zm3/CcXLpWj
ByJw9tw/NOdA0l5/AKsTjzHuphJ95ibJjjQbXuKwTG0n5ls7Rsk42iTCu87rTO97
qJkFofmfQQbZ5QDtowjYHK4D/F7mpwkoBdkg59c7qB8cvj8sA5xMeYH3enaTGry+
a/rdFKEufytkxWolVE46KNS9YqAl/7uJel5e/4e2n3ZRJ7rF4n00iJ8I4YJf5JFi
KN12vW1XA2BSxHDRJB8pG6RcqdC4Vojhb5kaBKP6tSP9ZccaeofLkThnFN+UXYOR
tKUQCVxCTUelXEZXwLzeINStpo7KPIrCuiDIH6Tuvf8rsF5jy22KR8oMtfaymNGy
qoRpoAHS7ib76AE1lVYxOlizIGbpEFY6Cb7cjtBomspGknPVP+emQxELr88TK6A8
omx/f/ew4T7US6w8ehrsrzLKFT3GGnesngKqeWwzTfyx+viVbELfUOHWpcuC0HiO
0uPUT+d7FxDRH2bFDNfGfgpcJ9gX7yqhsjYUeCMAsnymaFwoGZMJ+5ctvgIoevx/
uEkYCYGm8naUhUMSZ26h2eV0/HowlObjXOFBkoYRICdZ6WcVYpf2XWvsaO7045ri
xJfhzVu01zNZbdijMIw5ur2gw4pZnfI1Bt0WDl/8OGX2kJh82keBDCJtYVkMedzE
7jXzGP5aMP6uO7nJTyzv8TPrcWqLRHuAI71DxK41tcgR+6nRRm6IZdg8a/+4l3JS
2J9vku9NumCJO6bEf/zRBGNnTugbCA9QC+A3dE0zfSRanJ+VILrm8rmaB3X5VrCB
JU1/Bs6KpE7Qj9Je22ekeviVNZ+Wa0jZTRCtTQ+bhS5WxUD0Aie0MLe9ff6rxouK
GegTbM+Bi5YI+RfiSFWMnrpWvRHIwsFZdRDAy4rgP1vNOjnDbX65D+aj7q2OwfP3
zq+UVIRHfK6Wvmuh6Nlkjw8HOPm4GMTTwiumcoOYCVyRxPMswm42yPIxJn6RDs4/
KFFlZAMN9EKnMXkAdL2nsjE5eorodp4PoWLIsyC6+ChRNrCg03rSGD0blTpghJG8
+niEmGCPah4K73jLm7OzKZ74D/BY3iFDY/6+ddOsS8NGWyA18bQqCyhVEZv3yn1b
pR00FSXeGboB7ehmrwNYyfqjbO+vM/f41YfuT1H47Mmf+9TIV4WUM0a75q0+nBLB
ITxSTi6NYxdT5irXaaVSBPR+PQI/DzXjbvx8djUMMjjIgwiGxQzl8YwSo49IMy+R
5hP00X0l8uDuex2oPmnMtjvPpcIzf2Xo8ccgBK7mnAY58MAlFr+GMMR0l91RBwNr
iEIwGQvpJjaabUoXHPSfaDw9txbo3zETcw4bISrWO4Sr/meW87Gja/iN/D6qq4aY
w2Xx6lVMAq4TuCvastMWASe76azjN+Evpd1axJm9u9qh1L/TOz1mGTaPOZbO7rnb
qWKIO5aCLeIlj0lKjgw8ueHLhMnk3r+s/c5+/wvndBHEx+95jKR5iVYBTTpVXuMV
gwr3HxuL58I86oPHpmnvU7bquqfG+GP9X7znXGWvd1KYuDmIvFg9a+20zOJFKjeM
vYMarjeWM/81WNnTsd3U338cyrVeKRxl2Jf58BmGH8+QrhGnG5nQ2lHgzfEO+ej1
LNWMTOdIwJxkaotmwrLj9vcGXbS3L5YYcxRqHFI9EsU8U+3aQU3wWKn3YXPoa4Hc
FlQLLQZahnMrT2JFXoLGLRe9JSmjM6NIYHOTJMpWrQn/DCp47xDnAGLxqHETI65f
jWQ6Ij/VRCDCue9Z1ohLEP136qbSWQ47Ma3g087VLH4eIhVFpgwf81qNQNgFaVdZ
Q1OMaMtWQMD6FDqCTWCnU1fCVo+yys1z8hDTcJdPnub3vW6exkrpi5EZWEsFhK0k
7zkCUVdPGD4sXtQuhbpZCbJMmKJEg+uIV9uP/J7paWOrtgRBal6cG0ZBNqol26N0
x6LQ5RpeOF36STDKMCZsbbrkH4S6u2XibKZNyCJOmCQSivXC9nT2rRG2K5CZDfLY
c5VMNQSyPHLkHmgb/PFIrMcZpPZZBMn3Gi+gtRIMBEG5u9lyk2D3esOL7L/Tgx8Q
fKiOuX58ykH6nK2YoVCTzEbJc0wKGXkhvV8/117YhKHya6A0fVbE5BUxNaCX6PO5
G5rVd4H+xjecOTXw2mMqkvgCgLse4Lek3y8jZLEiH8DcyKaq+5BL6Qbxq38mnM4F
SP2buYLrytg+sORvhNCx/ezegSib9TcR6AHLQ4mGX/QpuBnCkrqwqziZPGr8Md0O
m5neKVLuZLHQy2wT7+MjXNpYwkzilC5RQwpF5Fk0b2KPVeFXjdLiwXbU4urUM4Cd
wq9FllzW2JRmGfgI+KEY8JdjRjdLmrMK6yxOnq6A1hxnrlmkW4X+k1uHZcDlR9j5
yI0YKNjczedDM5eOPfjcN+BuIpLyI9td+rTv5YPCdcbeADCRm87GxtZSES9iYcTk
zE7QTKIYTbamiVAMfojL8A2q+Tu1kpIrIDwthU3l9pMQj8qwH+c9ddU7xIe+brsf
g5adEL6mGDDUvMifYLfmaqvZTMqCNdCl3qQJVEqezbMkRF/rTo1LoZvBTK06sVWi
Uhn5UanxiQFHwL3C5f9yn2/2dA367f4aroQ12vePF6VgBeZcegujT2n2ow9aqltc
PWO5aLlsVydhUx/wzAy0K42holwHUHy09oqKHgEnzW3+4T0ffuNu7DdW8g4ynSGj
QN7ln6uK6Zlgm7TooBhpx+abkg8XlCOY0ioWXAA3WubPzHQcpBtpL+GtUDSFQh4x
72aGW2PMdEnK/wpAwcgWxYfQ9KGLvaoB7rwkzlUX8ULfK0u25Z+mUZ8uu/om88YI
X1YE7o2zHrGp4poCcJOmkCoYghwgY5clzjWp/+z/hezMIQJRxOVpy7M9HjAY3ytT
mYzwdasnKjTaTJftMG4T00GuI58FYNjoXvxFxuS2eODrcqPyD5brNPWfwz/weRwB
Qf7XVIg01IQPSxjfuFsMYEkG9WmkVCbkd3TozctQV6q+aJED3RKohejuy+bGUrnd
/4rxOuCfUaiS+hDXafjNZRKwxGSpG3Qhd0jnnw5iSTf+mDzxYYGsDm6g38OLxToB
h1cVED0ltAr9/nFH/Q/MsZO8sp05Ff01z4W8Us25j1EWYytn2eFjYN0QmO/46u2E
Gfldc+PmSNT57PvsWuVKMFpiqtLQE2yCHfN1DCUSvk42PxC8m4gEBGpdy2Ia0J2a
W7lRKkTEBHH6ADPSSqodFJsC9fdFTdOXMmFrbuZfzgLXjXdt/WBxRlqmR3/tJzfg
FKMbebefQQgg8s9oedJVeT+45cGisQGkPEk0BUY6HMoLNa7yCHsUrJImlvmCAfDy
XryfGBb8fpe8OCUwjpQ6p/o/grenWO1EpLKX59ESOyLE+zgAFD4xNd72dQrO6pe1
vXnETSfwfmqaBZ1KpUY9MSWSkes44O+tEGQrs2GbOW/QBUpk7djv8Er9qpEHpapB
KpeBJGn+aqwYnpiMjfcJvR1NXwhC+Psxi+JUoxIoHK4od51KmPTlYQsK+0YxmbWJ
+YcP+9pF931/JNHXeUiftsvSM6OynlBeNjqCwFn3TEQn3G/6FA5VW2sAOtBbzaeR
e/s/NPpggmmbi2cdwuzsYOHp58YXAnlsIbbpqKyljknM7kHxSCMhu2BCGv31XRUC
+UD5hyeoDjYdkhkQRUiUtiuN7eb3IKd30AaSfp99S6ohZDaTNsXgQ1YADkBZOghP
ZRVnG054AnuiYSo1GmBzZvxZZVxwgzUwuflxZW0yj9pXhHagfeQUgcn/IN/i58B1
Botbc6m9SBxXFRkyxmyeUkcQ7O2paRZloJ3/yxIDq7pLYSmxs8c99gYqwb+cFH7N
cMJS/+Z4nRvx3bALxXTxyi+jzRGl0H2xXBxUSLE7cvjkhqmtwHANqd+JJrULZ9+9
GULVjp/dywjhz38EhMV/ix/+aVlJjgLlFab/IYb1M0pVeusLv1NpzEoO/spnjG/K
o/1p7O/bNOAc+7enHM6VLfjKKhoCj6ovR9IA1CjKgWqSr9iW+ULZK8Md5pBOqZ1a
Z0M8zV0du6FnsiIm3bUQ/guI6FwcrnCtrPn7EDtn3Kw6qEDBAMWGE8O9EtWTDDcT
b2G82paZDbEqk5F3bBCxEb57R94uKGB/5b7cmRA3TXSIriPC8B2Rm/YyqgfSsWus
OYsZ1FYW/y6U12gHh3EA90BOlSplMz+12Qwm0bHGzohAgI/6xoVVgJX908zlYylp
lOex+ANJYFFZ0KUjTmep3bUZd3qCK+W8cPYdeIVaCZHn0emrZjNERbs9T8+1yocz
IsvSfKbO24c+2Red2fc6VnFtVZqTf1rCTuRotOXh8qtZedDP1RWAGDkxWs+tCIgl
/CKHwwq5o52z7dmz6UMP8/QpJt6DzYa8MON2VCzi8xOkPHu1SHzzoCxYUqNTRPau
3D0cZv2AzUZSfzEEYn20udk3Y9pWTPrDmPRndDNEDXw7yZtwem6cklR2svOOGVje
IEIq61gmRR7w2ZPqu/r2GUgd4wzB5XpgiYR+n8GupaGZwIb++GWKZnlw1XMPDelv
z0ULVfEBRM9vNRxwvJahY3EplA4pDlmWQBM8mb1+rdYeFNkeiXHvXsN+8nxgP9jE
xytm36QDkiyeaI2FmJRpkG7HEZMZRoblsboP547A7T62cdFr20GHJqwSnPjefcJB
wcL9IzKFoBPsrDHdWKeyQCDsKNVSa3zLYHofG+bxItseMwgk5qInzOkxOQdZGPND
ujdQd1iPkKTK5vc8kLDzK46MmIuUDKgcb/Hdyy64Ar3fWgaSHl6cLFK/TWYshoD7
VUNW7euWyoT9nA8y4k6Lz1CU6Tbqv+vT07zwMEwjsUqN2OyfA5P3iYick8k6pSva
yo8l+0Q7tKqErrxjHiHpaQu0JKjIIPU7Bmghs/DIwQXXqBw8lQ6zoQlSEP5soGpV
7Y/F4CIT9Qh1fByJHMLdBlCtFfrdFB43v8m7IMi7yJhUxtXhiiUYDjwcnYt6QFw2
1DJWWEbVkxhLGBmyuv35jjBikv9CY5oyxqGOnqHjqlvMPfF8XQ8fFzW+LsOY9IOj
i3rOb6J2CMSAq/15st0M7DGCVwzGCDPyqjbozJu5HN5O81zSxdxNNuB3crH8yFXl
I9kJIxJbv8wQJKT7NoBhvrvuTiGD/fSE+4Gb9fFIdMmwZv2nta0ND28yjyLQ/wmc
TAWbxc2AZcjbagkrMa4xQNjHstBc4eqoPvGx6x0KGTm4XxPCn7KxR0MKMraTiQVT
m/ZGeh/MMEc2iBQPnHIV8Yd6naIYvtZVsY2q2kIOT8nPT19ElrVLr8TD+qcsilNg
XsFCf2sBmpr20Hn7myJ7zrRdq+138uOMEQ97+GtMrCStPT27sUuLXilVRRBZj9S0
8C3FGHX7kln6RdDTEda1GuFio+wMlliywvf+VAgujcsYbLOGjAc0TEyLhdUHOrhN
F9rZOM4wA0lSmPUs+QDCGovPheQPcNTbKZQGpMj1iRNzdePHLll+qCJ8jXQmz+ha
6Pcg/ChnAyBdwKX6xdKpqVUEbHzPi4gyBsNq8Dk7UUTuXH1d57OLYKHddAlrQ/Ap
hwxPzPhLOgb1y8gkB1MkfmpGfEbaHh+XIPQCfpmfva8SIn38cW8QBCsFqRuWn6Rn
1nTK6HoyjNQ6lFjOH8QZ7nY0fnN/e5jjFOSHCLGJYaPAtxOxDvoDmogT6kfEfmRH
6eMtGuQHhklJ31RH53ZMLtsMEaNNxRiVDvfHJEdfHe/iLd7RggANvT0SAtHwST+x
2z/ZFdDQ/coSViIgSqUrRAAjrWPqPQ8yRxJ1NIKG/GeHFabizBo7PTH/P8isDwDo
yai8p0Si5eg9ysgVufPIqSWIr10ktpyFJ1ZG9hbjHy2ZOk7aS298vRfoLCZkuxT2
eGySPJj2XYmSPgmdy5JKL5vHlFqIKrNxJikiyHfhyree7ZcFss2WLXvmRMK4G5KB
V5Kjur+sxFwGaj+FPN5xY7WezlMQFamBTsx5oKE6FGQfnw8rokhXfIMWOEGOoSF2
rKKTuYZIyCs8Ceudpcc/Iwn7MwsmEJXBj7o6she02YwhXKkftWNszzZAcjWMfOSD
zyCJDBisnbrlLRb6gw9T60hTGgyJp9xLigeAKp8RKird3eF0RxnlBktZJohKGGCK
NkTZf93Iids83yuA8XTxizggo4t7/X1HAL+MOiLpEwzhb8gKKETdpkjkpaXpgLcb
l2x9cQNqPDj5d7hrV/KXJRelsFsXQM34l8hyxvOUSw20QCf+GGUH+BtO0gNwyuo5
WflO6SbKd6/e58xoZt1jAlczOXDjWHsNxt6dyPedq3qyGZZa+y9JqD1jd/d/PhZR
j3S0UQymtx6FVsZ/31YJXsvM7/yXvA+uR58wzJtQW8YMs0if6vDQtqep4rqyIlQT
KrsHK45VJTcHr1aGv7Q3l5+8mXogq5sWPsEA+q/3WN4Pn9rQG0MX7nqyTIRokqdC
N90NFfps1l1yLguxJYqaFdUmpjdsUTsKTqVS1mCDfemqlUSUmUX97tBZ76iltxIJ
JhKrklqzstx5Qpqx/B0kIU00mCpEngeeiwYxCy5ExX7FuYGSORaBORJsiPPj2aGb
XgYmW/MEuFsItdnBHKb6OkqwlGfQy7L3lK7eFNXr2Yggp+2SRumWufq4D69urk5k
kMju+QR8NIFxmzWlwmggP1mDLXo1+djaBPG1U90CjqSMaB+nL6geqUAW8E94OCeq
0dea85kG3w9F/7lPdtAjhQOXB4DFZFmAatboMJgu8/P1PU8tSsJORW9TXRtcpqEh
NlkesSl3T/+wwkfMJMSREsR5Hl0v1ShddGSRFgdRo/ufa3Isb2Gmp+8ghRHXMmli
s7AFet61uWtPB6C9bRS/YMwwDyYXYfJUsIr7lm+agUq4lNzF9yRZ3OWBog3g/ph8
7LW+1B2+GSwIJDCg1YU4cRdEAffcNejtDYgF5UY/ExsqtUcP926kNphicmKTWPjm
Frc0tktLJy4wnYbOPEft4m+xvGo/JDov6Cwb1aGiuUrZwjl2SU5JwAYaqP9nCcBf
bBeWVkciNbfzC+NfMkZixXuDmYHLvJfDfSuUQsIWMn51DlyoOTcJMHttfm4GOXPR
tsL1JEb1BXKcp70hS2gH0s47ui5zSGE98u7TW/HFH/qTvuw4XFvcFvfYkIKIfeOx
IGW7J9/46Mir9YltL1BOqe+NiA/RrgiFI+kHOnzFhs/FWz+SF3XRNmZo2RTDMdvd
yP9lEmO/QGdgk4Px3L0k6QZcKe5UoTMKuIPDFmlXlSSaIavqp/jf95Mur3bgQsWt
5HK7+QnYY+Aq3a3WQvigmoXwA1XoWBAXpPGmRmfQ92S1gEUcHKkJDy5DL5XpvF9T
s0UNorWfsdhm8hr7nkC4MI44Qjug8aktroAYjRkcPUGneP8/gt+0t4rFQ4hxytyK
SowLXRdcUvuBWXzFlzLMSiqMJMfMHD4LPUhDSy2ArOpx5xnNTjWdiQEPKpqnY6WE
gGGbSmxxFJWI6TFs9xsUTo4kwtt3BPHC3cP84Zvlki77MXukRkT0SL0yAa4WJ18P
mWmShmgq6xXw67C6O2mzMHADLwH5dJGmqE6J8eHTLUhXs4b0dkqmW49cA0nnbVZe
662GhRfjlL9ccGjR1p2C8tIr0DLqMSiQPGF4AtT+XGgISoP4hlmeYXMUjyP+AFWO
hb4qp/uUUW6ze0D+0DUqkfJQG3hOew4FPRGWhwDXb1u41jqMOCiT1eyIprOPEUhC
DYk4ZzQwZjKh//9c0qhGgzdqVoS6fm5UoynsViQUVeAFLyR9P2Xx73I311G25d6R
pOHyrQGw0CbDdPlmtKQNsDXxoR7t1yWA/FybFyHKowV7OT44e4aqfZm/3fQaqfSQ
0Fslggmz7ZIVAZ48oJxZW/cXxtwbuuaAUvjLK0dhOZPSfV9wKJ8NfoCGgn0ZGjXn
/2hUon0G3HOS4jEXcs7Y8JMm+7EDAjSan7LgoOWtfT0+ly4ylcKGbA9aoC0/CE2j
MwZzU7SQbC68Jgrj6lljOlxDBfdRp+LgGNSS6fWV2BYoWytzfSqw33tqiBLUsnHn
tvv0zoYZ7b8GOPEoS7Qly1KckoyUYzqmdHpxqWe5Y2Z9UAZdV90The6+FQG2NgBN
4o/GeByi5zGic3BhqwQdy68Y5SlRi9m0jQAGMwmIuECS6RWhQayKFfHZO/bntdcy
Yq0hcaOn9JiAzxTSvMwj92mHrnlz8hlW63PEdS90GvPSUriiuHhJ8aRb71Fc2KlN
GXfIXLbpqx+q/mNfkMQQEgC5nw2rjfBtivFrlA8RNkLdI+HAZTA3NhxaxnmRWzvv
TSsbs89o+6IHRegaK5TEDpfyhd+vcA6hO3rpZt7Cf1UTtY2kq3w4WhpZeSRmh3HL
YPOtEZ6yobiBTbMgkJdfMsYQ84LMKiDh0uxiAZpXNHg+l/hOF8Pa8Dbey3Xojfsf
IteYLQla/EqXZqTbgBlBy/OCwvm0RHvEKq9dpa0soTsNhAOGAvJ2yicrEtOIsL0B
GDYf8UI3xq/RjTNws5m0J7zO/eHg8g+ciihGVPxQvSAg2sM1XnJLsBjwaqhwBR0w
G7qgQfzVkGeWZGWOnyCyT63iERXqj270yPFNLsGRHZk3orxPh1wqh/f2K3Bm+rUY
IfQtywyKP/bTavM8tkxP9eV/aYPNZAuBIofYDrt4HM16OzflkxLAP7yDQbjWgy+W
eOzkqgB0Jvok+0MDCJqOYydWSirPDx6rGl4dVfixeEMrnTHjx8DVE0w02kCc6tWs
sIFFE0mrSToVvv0EqGhpa1QeT+UDqGu6QuDmZkOPnIy5xBBR8amXhjIDjU2Hvcys
LwpelUHB8Re6ZLUFZ7EbZM1ifU1f/z6c1i67rr4b+yv0vUCerbTD0LzxbYBaywJ9
ilThOJGWsGw2wz8TO0zfO/PsfsVKY3+8sasECRLrfuenLeaMNDg2XnleOQMLVyap
cofjo1m5fO3lCDMm4QKGIhLlHw8Wilbj7FQpZtDv9HzQ9bkd37uHCBYegNJfacgc
doY3u1tqFtnk/HUL9U6si1zmjx2dS14kAJF3GEzqwXxZFd6ht1aPThdOzy9tqJfO
7YmV8NPuUueOHjECGiyHA9bAHbD6EY+Hi9j/LKfCp/OEyTz6t8fN2Dzpn71/DtUT
QzXYl6Xsu6+iLc2BbxZXXQ4NxMN4FWstIKwdam4qZAJ5rcJy9Er6qg0tbhQdptNZ
+NVig2yCeNiD41femlE1UJLy97Q5uWTFecpGLo4HfIKRrUecY971gBMj4/JhQbj8
cFoXbZL+0l11kGse4QdvUySnGnsJVBM8jbbhsPgBTiTqpMPtw0bFNLtmhy29Wpy6
5KW3A0sIubJcNHBV7ZJ5Kdo08Gud0iw5ESll0mlts6n2qa0TPeCHswBiGbVpowjI
OQkJEAgKgX0wYP+mpFJcw+uvwFHHWqL8b897mjdkDbZ1/3AmBrZmxP/Y+pHa/RT2
AklbW1OfXdkDSf0f2LY4XWd++Rttu2PZy3Z8Z198EcQu0QGNFupTPC/2pK8kw5Xk
FeklsZ7LkN2YIzncBsd059edGcahsC75XTNEBKOb1McEy8v2voQEIG7DU6hTEiUD
HS4HN3jVNhuroMToLMOS0pNJznEgwQPrVbZ+2czazyNB8suUKPmNgfpM5qMZvLHs
8/h2JlyCtih91pNoT2Do/cba1uXm3TI5PjnTVt4psEyf6/z5AmsttdV9X8M9GQH0
geBCNZllA3EoUj/wCmSxa/3fTgpiQR1Wtq/BEdgw+FKNnmQ9hXgUz+8PiovAYWSU
/dyYUhnd79C9PTkPYwoyYHP2vwRkGK0USStcusYrEnlmtghK8GZQLOdOkKg/CcRg
+nRrn5zELKd8+r1TQ5+FjGwsUAS/ka54a10vW+OWqN8DN6NpBOQn955GToj05ZLC
ccgWEzAevmX379cvE77oEEfru0fliBxM6wuIQTuYfn3pKxJewvvauPHAlGhyKr/C
VjbLK8yX1bCMI3WvUgkXcBbC9QdFSAZkcge1fDTjhIcJWB82GvYKh0pRAF8VYgmq
lRYWcy5N1llwK5Hd4eCvmW2wBIk2U4hkyitfIGV9q1QXJvL6eBjj+riB7YUWPOcK
hLl2hGxUbmUo8XxYT//z9k5LFNaU2snricZtMMo+f6sE3V1QxlO+ZWEMda2RaQVT
I8wiSSlvD8yRAqoLrdDAhc7zm/busE20SRGikzGCcik948Ijiva3O6nPJxNVMxew
MqbSj/NfGx8W2uxSDZsr0I3/IdwKqvUYbraiHqeYklDPT/h+Hy55H7HoLr7gUbNm
NzJSYS4FO7q4fxo0YNc8IFYT5pGUydIVwImNcjTQGWG2Too1a0Zvd892k6mU3ryH
Mz7SF8oHZBeG6GFYIQwi7BdGB0EtQjQcsJqQ0hWb2YuIzqf/6dzafSJLUU/tDpX/
4fovcBvIzsxIJCiJ6387ZEuUjp0IMczT34Kq1hQRscdEKYHqJAosT74ScfnnvU/X
AiwCokugilqvYuvdTbSe4onD8K3Iumv4XCdIYLcGM2YDaUzvz/utEZOv3Yu7H+lW
NVA6BzytrRzZLmM82sS31HbUzV++e/SikndxPDYUO99tdbKcUj8/IeymXncCsp0g
6YxSRaxGILSOkL5GxrJHvHG4KhMcKrSQzOiDCajFAm8PhVChPBSRVP5/Ed+M2I7L
SN6otkuAsvazEhGDtRZSStT6pIVMHuWKdUEDAPc9NuWxRU08Wsy0zS3VQ5gD/YZK
zFx2nYpTI6fQ+XTSL6UZYnnW385q85lKDJtboROdwt/i7Nw8oZoyZc7pefgfOrRM
JIhMPlq34OeUMpnri+itFwINPrJ44RLKvSRpjm9MoPvkOglFoNW4XK/VY6z8wMPr
g5qindM3OkhVpZRPSn/pTljp4oTWwwGx+E70yjx2sv9XxdMIONOOVT+NHL721S39
a9ltpJLg+9bvwq1JUsOSb1p/+fhfFew3CaEKDJM2w5qLWBEbR0QKqkEqzBFb1phD
pP45BTvewSat8Cr8a2nHdrn0JRZwW6bzIpJIlDiwn16YNXAJJQkGD07SYHCnk8vx
nOyXPnFf7cSAf1i3BLCuNzqXryW8zz0WMxyJgKg5JZZd8lz82hqxBjARtuETcfik
pHx9P4bk3VTFfRCqCCp+zSkQZYJeZnbSkIPhmeWNT5KOFJPLgQ5gwk595E9/ASu1
7IXIqOHzyxLbdTMXiLIdQa0T0RGL5whogI7TCCbdmbiASVOSjjHk0NuOLfVhnEXU
0Om0EfhJlM3YeLNEKR2heQ/XUygl3jQIcd5PW8RNT8+EinBwCHk/+itXnD84fkHg
jEE52l4yGOVcxO8B7rwyh5yOA+OYm8fYQvic8BpkvfWdLtWhePdLhbdv97j/f/O3
WsdmeNOyw/uv6JVVrbPFR4UolE4rKGSMyeYp0n1Ui44hdBM6fGCwYEfg06GhGwgp
ZWFnLMBmlLYH5QqzfJFT5DqYNXiTL44UxxEEWl5A0yTjOp/nEiZ/mvQIWqYC3GkP
3iuaBrAWcvQPjzPqR3nIz9QNBUWNWLuCyP8iWhflEf4ZGPlMMz6zBOPBAJ47JN/b
wBe6I4WUWYEeWoYnVEVgBpYlQywH5HkMyC3wgkEmlrqQKqxN3DrDU5vijJblW2xq
Sm4idQ/kPKOnFRSszFXhPsuNb67XaKvIutWFVU8RdGZdYHiI9+ClzJmEnXSEaW0O
QODNRcwCzkiWals+P2/Hx9nBXWimI4BYtOJmEmd85dJ+lcJN5Slo9zO2gg2fzcXj
dNVwWixeznduBtyTkvIjmVvzfbfOhK9X6CQjVNNooENnXNG9UeL5JgeqJGNcmcP6
sZ8wjX7hm80r1uDi02X4W6ZoBK3i41rDf+oTpawNiTMHQIvNiLMnxb0VvGD6p0Lu
DDDauOhinrRT9UHsYBooCWSDfukZXQrKm4s8qD485COH3+e46iKw8IiysU98qnpu
aUoyPNY7yoBLsss8o30jeuwxVMXVwvNCsWAk+799ZSlUmGNnRA+3Ll60O2+Dq5Jq
B6A5zsfJ7LoGaucioXg3i/2PZUzPORH7TmK6lhCOJvlm0VmoiiretUnTWqOjkGCC
eLq7a8VLxO4LyLGMfZnqoOx57z/H2pWFYdFSAOKgWy85bxI6rRSncC1hr/lL8UT2
TFKDUICW90n2OOHAGDhjNXxmqZr6+zZ3rC54QdhPV61wt0D3oF5gQsd80vp4jOr0
wNoQ6s/HM5zJW7HThPlLI5HP51pPdKZ8gJq4RBg4gKSGdNYMGtkp2NBrz07u7PcF
f5J/8F+YBm9uQAZmiMYMs0Ykbb+r5TjJJfLiyx+vP+oS6fWI4fRlcWR9l7iREGBy
IYs09efe32hzKl9yS8HqtZxLGtSMUxvjMGfUaYv36OU8FHgnWPD6M0hK7HL4PHeD
zUKdAXDAM/+aBfRknOIi4oIDYBvqRjOdCrH0Z8hyqC76tNrQ+99elU0HdCKhCTqq
PrZ1OCF7mpLyXjDHH8xxEEwVm6wS1qSSPbvBziblf7eGtS3Tj8eb4QJ9AhKmXIdD
JWg89FTwnI26WYM2Um2HpNg/oa3mcmsIvAHC05+yqnqEc1KUeRKHE9/SYittGwRl
8jaa/TUD7GqArHDQaP7hLzUuKjdfR4BT06JSXbHBlYkIEXn17njkR/CfbMTopykX
N8dANEmqkWEIs3jbndoraZLucmB0h9s3lDtpNStlBqYI5Ev9DjrfMyTzTNZ/1x/s
8b25ZN8pTmh/VfoTlDqoUOSA5zyLW6E5XpPyHUsDz6Q+DfZFwcxNPct57f4lR9bA
ly8hiErO6dMOptdCwwiCMTa8rarTr4rMJWTPfGNxO8sLsM1E4/4Nd1oeZTwuaK1y
T0defYh2yyRvAzcdtPAJbJPIb2RPGmQiguNT7dy/bZmrja7KKBuCZXIAuNmem0XI
zfB9QzAqVAGFoBUUYqshlHCURVJpkGSbiWe5bhbItpR1OOj/jbdKRRQ7Qio9tCP0
BvoC1V/pywuS8qbVqMaYePGOkA888Xrn5bdcQn5kf58Tf57XHyQZ61V15LmtvfP1
cC9HKZc9ro9Que8xZyGnhBOG9iBY0r1seCVX7j5ytqIWQdFQ+v1oNOLeK+wOcWGs
fQlze93ixQzzzeUg7t5tXoP2Q07TFmIXANXwR0dYTF94/7Lk5qr8oFaVNfVg5jHi
4b83EnN8qfE3S4mUYbGuW+LFGqvqzgeO7IsBzSZozqYXi4RiSkVZFO7XPNnoKvPp
SO+UytsPmjcnAKKD4VzZAnE968vq4wrO5kwAoQquGwPeUWFfxDD2twYp6tYcdKQ3
Vj48P+G18h6Du726MN0F0G7G9uFsi5oNFB/ATAslRUwMcPMV3J5yQC+S3jd/QE0E
6ziuGxFnbYaOvjOhBZkrSFnp0WYK8V96namkTNueNSEsLdVzDmYPyft123/lw8nH
kohEG+RBAELOZ4wJwz16lzc6Dxa7S4NaH4RKCOiKqMAP7Y5/nsNHXOzA8pA0aQS8
UksmEv8ri5T0Uh+4g3Q2OqcFl/4193Jj+2G+GF4LSzqAnO+rSS3yoK3dIAn32bwd
Zx2yTwrHUf+MN8XSr+wLsbmv4WLP7VmIHXkhkzHAxokQyUlX/LkGnwD/s0KBFFRe
dt3JnKshcy1/AWfGKoTdNDNLYYjkB9fpdMrQwzVyNQijFuM+lLhEkVpV3FllHyoB
kkZxvpy2VECS+QQMp6qvmJePeyFYU5B/cmx8Ed+4rRJ2GZ7xK1Mr5rxajAlGw79x
1m0KqZELZ/Mrc6V5mwxce7tJLHjJ1etF8Jsz7BIqjReCSwebRKt/YAbqFav0uejI
sYERkItBP1zoZAwIumwY2QSeb2ynd82EQcWngO5OhgHb7JX0xTDteFMqiPEgkeUU
VNZCkmWwPEseBO7xRIvxVu8/EcabMoVyrpG+huaCU3fSoaRtR4f5inuV6GygWZZc
y9GeYTU7teZ2u5zL50Tk0CEY5iuDE/+dQDcxa6VKuMdvWqB12rI1esPMZZ04GRnb
D/QYfHKAy0JTVtFIO56Dm4eLpg27o/xHS3T4mSr1vNVB3U6W7FmPylqNecdRiRNm
MCxIPqyqZeut/9U+Tb+JkQIxV4TbZTAu9rz8Uz4WLFcRWkcQp6j07Li+m1h9BHag
oHWgoLvt6seAQXBzM+Owpk+N70kNBOFVZWwCtwJ90V8KuH++vknkrsnSQSMemGMO
vdvX3ZjPKwDtDdQfugkKl/887i1L87X0GT86/rfV0OAEyZO9ALvl3cNdFE0F+igm
xFYy1gos2l92g1xibf2B5lC4YCq3OS1u3R8zBRAm9K494jALsTsQlJCkUbTLJX8r
S0noV+zKQTWTk+7j/lRWdS76bhfvWxYnUTAju0AmrnqIBxOw21BSmcqNutPR1NPH
kuiYC21gavelpFSvLRu9Zh+elPAXKMSmp1a/ICLEWfCsNd9vFd3i/Jiu7EF/qbCC
TRqiBl3n8cz4wIKp40fY9/S7TvnY+fhZs1XWLA1ySF0HbXpa5ckBn32xuLDIso4t
3YmqbWFZ4OdQE7zYzML/w+ATmOiVeBM2/olDFUht821lvjAlJ5Q6xg4F3npLouXD
QQ3qTFmriXZXFhZ1o6I9Uq8/Znj+WwPxiqnIAOsfD2nIdKcTk20qYPPK9DqshPjJ
YQaT8O5eu0K9RV+pS3EO9cB/85L6O5KGrGk+ECHirUS6G35DMS655Y8zrCNoJEVB
yTkVFuS9kcZB7LpaOMg2eWDIqe13HXxD0BfxF3HEE0PxNPPcc3Y6U1hFpdNKm6mp
hmAnIhSnxfOGlZnbxqgK5KW4+A17JuzKWN/6PwIIjiijLM4JhmWZvAOKo3Bsd/g8
5UmhQbLiszxzxyiK62f7Xc18b5CPLIzpdQxj4lEsj8EIkyQ9HvATdJilWIXRwJIM
FepKvh+SpBVXD2z8opk9aGWy1k9UQ2F5uR4gIgOt2CBA84CLZBkvhTDuw5L+K9yo
Vk+UadWHLDZoQ9rhlmd+qLc7AntYw+Pyg9RwpoIBRf/ttkWgWiyn+P+xTnoFcXve
5ih8GLfnSUc5vcn6BzrIZeOqUNgpB2VLa52eYT+3Mse8j1byHzwckBdEfIgchuJG
uVMSMoqL9iIOtZew5axQ8eusElJ6CvU7v66eC7lMizSOfe9UIceJjjA+1Nu8XJe+
QlsfuuM2kRUUDYCKnuSqh6YU/cTn6KdXmJds9Fs0ODwFfX7bKT0XcJ0JiY/CRxwt
taNgK31uYlqFoBgtFk5deI6FRZTdZ3luL3OQTvmYeK0GNvlJFyOL1+tcILCT8kpZ
cZi8W7SbwOQbtjB3T+QYPrH5w8LM8sD77bOPgCpHP2sb2Uh5fN28wZx5dhWHbryV
0+xs2GT9aDjagfXzbUDj0LCbFdDIxR6ii8zNs0GHilkCe6p8bJZDYyy+/PqjUxHu
EEQ9YUqEYCA5+A3CgCdoa1uHNhDtR1EvlEZUc9ti6KXAPtYPHju7CtmBQJJwOX0L
FWR2oiqVsEeddXjAowuvUEvyvRzTagjL1CJxv8kQzhF00YU+VgESHdQ26ABWK7/K
eoOCaW2AAzfBdkDFolPQCRleaDkCCLX8Ye+iUzvMlD/oZhaUu4c+AlgWPi2D4q2T
8oNMUoIeoFwA6YbT2MgXPd/xj1cVi6IMcELAtYWAuAXf2kPBOOIpCZ3ROF+xqPE1
LwZGYZ2cPv1piqMFxMFcFFip+y2mC+QiKzEimj4GCVYI3AIQ/4gHnoqBei7xQ4pO
XcwgmL7lCzKXydxs7imGhGMUoC8jTC+NE1pmXEp9b5PB6bq7B7KhybB/d1khvrKG
L19zmm+gRw7JaBdymw/kUimu7uRs10Wwa8ciMUxnnm/l4z0MO9KunBqaXRZmRpyE
1X4Ltag10Mx9ppIHmvE1uoLJqxvvz8hwPLdfeySsamRZr3vRTKByr498kEBITbs6
qArjSfGmCjE4HL9OkZd16CJpfF1yP27P4aP/uFIDXdR3fuf/h8u89OIAOn3FjMYd
z7hD+oI6pZlEfBP1BHNYDh/jx0bdZrXAapgCuvHPW+NRcXDbzET9PPZdxtEV+aBF
sl+31FQ8DXx4x7WtKHrgb+UtRhU1cmUtmSC8Bun9vhtMrXhJgd7NesWDHS4kHrH7
6TWBLC2Ckrh1mQ5nBCb26GCTEIcbpqR+H9M/rRiXrmTRPKiNg50fcm7iEQDHyjF8
nfuoX0JMTs4drwS+57gnHmC9L4/oVwjpUkTC+qegKukTrHIqRm3yRmZgipjH7LyF
R7EfIXLmmonDzGfAv4ylEQ+XKYVT8+9mxCDn3u9ot4gsF2boSuFjF79wew+Sb9UQ
TzqiD0/poFICNsCzpjpFzBSfXS2SmkKCAj1XA/pp7/qp38dCgkhU8K7tOprxQwYW
5IApHP49Hd1i98RuAjOcA6KBNyNR3cgQh/yTBi9FSI5ihsjSnVmQszYvNGFERZG2
twbZF4DkdrMmy5/W08mTm2zCLYSYu/KADeN4JIWaFZcqP/mB9mn7ihqCLyc9mn/l
ljx0dB85W/UMEjM+mg0brsNTIFMy5TaR11DCCER0j9+05MDT872NqWppJhWu2pCy
TOTKVSPw1lOP0nFBeCfeYTJE/1djcxZHjVxAKVOEYoQvEAu0h4kWah6bL/3VGStE
Q+E7xYRk5YHbNttuURwoeZ8jo1mqnAQVv6zgVmUmfaEC83l3Dxo6813segfm/nye
n4MmAyjtaE0g9Yh5FCxQNKxxwgqSbNk83S3HEUV14lKEbFAz/HnyfX550PWNaNd5
QfQLNEEkVXMZEAK2IYkyWku+X2HB2ofcAdzpA5kP3/t7dkhhPBGNLL+BIOCxullG
2anVca4EAnPKtsmOuYasZ6g9PsuziH+eEVlbI0neZOPnMsdWlE6Keyn+efDpE/8s
M/Z1nE5JdPq8f6mW1vbwdnAyFDOdSsTOPC+/ziARM0HnsO94hP6tlTQOXKzZBJ/R
PUBXI5iAqEdqa3LYE3qG8T2owBF7Tsgne3zhj74NjFMy44QEXWJnooz/QS1Ja86c
wBiOXkgcqz1DYZxN0IIjENo7luK8J8DvZPlGoDjA1A2DO2pgnUGckBOpjKumwqfP
FaPeOTzYfikHCpyWG0n/F8Es84/pkHO/ODCzYqMan9m0/aL4AvXL/ianZ8/fLzi2
g6416jb+80NBqX4ViWr0lDn8sx6gyv5eeTcLGzFLtfGaG/rPyxt5jVSJTBxfYPRw
yl/FLqw32499ge+nxshx+bcsmbJ9QtNGEkdbMR7I138M03UQotlSbL7oGl2BJFYS
2Mf/3nQt73fSmpLehH99y0+WPX5ZwcXBAQ1Gp5oVLUvs7GsTokYnc8JHp4400zLY
L+sRrYUEpsF3QvbFd6eRkq4WSHXVlYqHiGTPj0mmL3BrLYo5XXaRlZr+vQUZdZms
uk0TmZbhCaDZsnuXX048zR9SlygwZsoVV+bhC289gEkG5SFhggBDH1j3wYmdNISw
V9bH291N0rOiolWd5pD90ImMo9ZcF0fh22/4+LM/X24qZeM+/0HBYi6mRnXkU3TE
TI9uj3AMncVBC1QVDg7m6qaju2PUYB/Q0wt8iHzFccWEpQzMkunTlcenElSRCRB7
by80epFjwI4ZL1qMMxxcu6TUaLVSXChjzcd0Ymar0TTbiQWNtUEeLczD64jGPBYC
JS4Fk1s/cl0s+vDFWQUwJHm06vY+YmJdCZoq3LkDnvd2tmG+InytymeOxIu9h8Gc
CwT2OZMrbcOn/ajuO68YP4ijcYf7HIlA1sUo7s7hOq879vPME/OdYxpLidOENYqB
bWSrRCwBcwbz1daHV12tO6nGctG6zNW+j1T6VQ5aAiljQNRGTBRViVX8OVGrbPo8
YBbmxFzADSM0mH6bSn+SZDEXXTCOi3EsriH9TVy+jotoU9GrxTNplIHbUz1ArO1+
GZ4EcBqAkLDonMX13NmYMOaDm55TslCrBPkGZUQF28sOQTD3O7Th7iQexoQmszjt
F4CgVHNZhsYdUohRiNTyfMTpq4htj5ChGNVIiNNh7CF6JjRy5SjpaZvvKKxh24h+
OJX0WD3P6kh+p2IJdLkxl/+CuxUX7iSGKOe/nWrIOLWjuDlockw9JGtImhzbr9Y4
mslcm58BPFr2JIDFmw0IOgnI/YsmdXnppuypUMOumIaLRoLDVq7ZDlZpnVqq0GXD
sBx1nq2AkbWzQTaNcX+6O0ZDsoKlwh/Roi73Wkyaq4YUtnA0fGVPcbgU9thmd6Qa
FVtgLqf3xjjodCDcfbMngrHPDBVhNiFz2/LDuDDFsbkXyuskVsutWzsioY15xpix
dEN7jc5AvlFDQe3yKaoxpKupq8o/Zb0SKMyERoOIy+b8AmL/7KWc196L8/kUQkD8
nZM3fcHs3vX0Xbe9Akidqu8hcGX6MvHNiPp9XZRx+Cn8602hXnHKW/OMt5QLkEST
sweICYDcwsM1u/jf8VRfpyIz3Gz1hU26SiunBKe0RlHIY2AWef+o3JrAO9VixyWW
o+tVhFrnCNNkYydZSo1R8FIrsPOmj87aEizRgaigDXuhCKyKkDrqbtd+/LzJCW7B
aHBmgmA+ViFANn27Xm49iQE8q4JEGUxUhIuSaRYJnfyjESKfNq6wml8GjzayOOoS
h2Y2BWSoc8q/n6yMvex9gI4SNi/3sz9Jbe0u1FUXTboNuiLdvgqqbVCReifV62EV
dPhCs7KbQYvsN4zmqM9RQV48C/UHtNOGZyA+U5OAcPGcgywdZ6jDka+Wx2MgjIN1
CsaTKtxl9xZuCZ0DbwU9Reu82o6VZfpzM+PoVOT6KoEQBJRVA246CHE+kUMSqarb
1UqRjMB2P8qtiFPf7Tmksp8riYl3dSdI+G+Vwze965OwC1WkSNNnYa8WARkJTzbW
g5fqDTY+YPiillRwQXltJsJ1jodsHcz6xDTOPlJkT7ij1CkuOQw87V8mvwiuw8+z
mNK38E0KWRaF3PvQgn8TXEEaKTkUpEY6DudK2R4d21CynuSbO7OkC4aUuJIBHjSu
TDtH8YqtwX9HmjlYFo4kp/mfrwlCSg2/BfwJZG4NCG9db65W38QZkWWuuTMO72+w
B6sCR+GvUfWFrovH/MNkooSi6EEbkFz5ikimpmGdfLWHnZ+D8ytRlivQ/VgPp03G
khpU/1eYIMSSPCbbe4KWnuMJwnHAC4YCW9Pt2Av2/dwAh2nnsX5TqSvulWThJ4JG
5C/TefoxRNytgDo/PxnVg9R5p0vt4hgtSOWXc9vrN44pxyK0dYR1a3hDBaXOVgkv
r0DWJOKcV/Z4UcVpEB8tlfdNTgPTfapIqBXiyKa5zRMJneYh9ZihfTJbax+Chvyn
WVeP1k03lkGx+LChHP9jno6Ip0WY7w5Vsbniha9tQ42MLjqEdf2L8wusAhVgKAmK
ctU8xDexL7AiW+LFWHpyJZV/bVerpw7SYNbQHqKUGy8Ze7JKXw8BdMmoSUEgHwe0
a8EHATrusF/swaAMwJix1giq3bFU6v2dbNkIUr56FXXoIVAPkwoyK5CkSp05cbls
H4V+8LWmKVWJf61PPgk9fxST3mmAa+TRuD0RUWx/SR2xTJSLj9JfjnV2zW/t3JmN
SSMKyKpQGU1l8yWTFG7grsslI41Krl04acyh6hId5/48mDtizGjn53LxgSiZPZYQ
b+9+ZwAVHepSIcxTzgFjS+1FgyrAzE+9h++QwdyxFO3SgDFYjvNFsImepf3rtEdT
HaoxI0+zVf4rHRXJEs3i4cL+9XMxSvyHxD5zu/8/Xeq41r/OgpiO5xflUtraxtXU
6wTIP7EwcHUahmcUAOUh87dLBtICN6yFPhEcLHZuDXWVNFcgHACnCOFkO6+NcvcD
AE2TnVc8yy7k8pyC6ANkDH+dEM6LX+nU022UivsTTCn4boDp+dpcDrmjbUDG/fnq
XpeDEwpAY4RODf635vTfY00RKJ+zjG7YzOgW4BnMfEuyvZhQVLz7MzZs5ubXopEQ
Tb3CRlpBsqmM8XqhgeUFnjEB19Hvs533bBtRxQhYJpMw0TQv1S4XEFU6afm558EO
4bzrNbM8AQvu8/8JCO3OuuuzCjdY+9KlFaHZgK9/M9pKZ8za+fucvp4/N0qetsK9
zytpoyQ5GFahkQiWKxvcskSqdwIrw5EhkeGezjU8qQxuT9BRy3jceJwQIxfI/EWs
Qd5GaJNAzLDcTJZyVYQA1S3l1jyxNWB0W7j6rVOpXKewtVJZLdoSEozzkZLF3G/q
l7PnfbzKbEIaAOv2NgU4p0jsU5vu7q0JfMDODjl8GgzZTd0HxC8pScPsrI7sPAV4
zx7CSWSIoU+Loj9yW5nNVF3D0OEQBUhUDUclGk9vFG8LcVogZVDME3V63Kf5Stgm
Wqdrpyald42pNXPsJSZ5mtfNQjQmHcRmhENcPDpUiJcrlhL5YRgbXq3v5zsgcC0H
oPeFpTAPkYKdY9taxqjEIFSXEeCHC+TSDOTLjjrgVJIK7awZcNl2Gt/vTE1ethqI
RzDe9tvbO0UjzBV5sDxD8JYOpl2xtNTOGj802GgeHncCkP7EQJTT2NERiAsDNEsm
Frb/XGRu0W9kU826xqLw41SWTFfhqdlstiUCdOdwlTsL5RCzkP+NKNTHEehFAmKo
/n55YI1srxUcKhfaXtzW9KLXS8/oHLtrZy8lUMH4DjYGmqzNDAfA6DZhY+UWIT6V
oFRURuKgg2WKmh0MBVXszDdnYqefcHYZgzUg9lwg6jMcntsb5hVT41xb0VCpjxEX
LZASPJRn/yIlHbXKZyMnKMDAgYjSyrIOrElGzPiMDbqShtkzIwyulO++NV0u65XK
0bYJPgTAZlcLGwju/geE819C3E5ey0//ZQBooQjaSvF7pZlAerEiUEqKJBGUQIRR
W5zPtP7cj5B74CVUhczFgqR2o3K4Lr2cG8uz8ip9+0z0KOxOaxb05E0uQ19jvo9G
LXG3oiWZY1lIZ8QQWQ0Ru0JZD/+bECPd6rw7SdIKyLnkhYcmVGX4P2sg3ezDjy2k
FvzUbRspc5SquxDZcNz3RVo3oF2jKOdPgsh7NvayiBM3YD14QSiSa02jrqzTGP2I
vpejdc1eOt17FyHyxqwtqZPmR/POZTXiOvLvagtCjEgaYoEuvekJ+HqrxFDJXXMm
yVsac+qaoahoNcg5qlnBsZsn1ksV4pvBtNKwZmdkLlHy9VwJzL39FM5j2549LgsK
upkc3UvrOfL2I55y9eEVQPo0CBSdBvRebWRsLplIWxMicPQav/yNswj3heqsp/A0
z3thtCelo4KPa/reqapUNvDhBo1qvsRd2ajyxvkScx0XP7sOrJDFOGCvR6fvN3SJ
CgwvzS6DxZrMmDXxTOd7ADDwb9JNgg3leOYta74uJqCjPmtqIG2gfbVVTCadZmT0
z8AbA1R4E3pLG1WATJ4tqVkEFsqRTvNGiQ7fdTztkQaQHC118BU7RozJGXRM493K
iu0fNmq+Hue8uXeUeBjXdwzWR5mk6NWIvh1NOLGLPduK+wD3a/AcoJa4LqEXiqeu
OXZ9SNRjeIuVFYALoIIWiuUR189JwY2nu76Od5X46aiXbfuxiObe6RAFh7i5EJUk
Lj3e8bgjjadolKo8mweSAS1QvVQKitJTP24VAFmKT7iSWxCljP68STGgvO7QpVUl
/YUT2M1VRkvCnYWO6Sg8ih7/D/XDbU+ooEVdQzNpCo3TRyvkM49f9s6DYN0iK1P9
/hPUv8C2kWjLQ/w9LFFcP8nL2ZKiyloLxCj48LGgId5DQ74te3y521yenQJ86JUH
Hf2Je9RhNz4D6uwEvl+puktMfAcnQID7z41LNkvmdPglZOT7V8nixQc470ZvTvol
u2VUa1a3Nddn6SqI9ciy+11hPiBkFy29LLqukBGeuXVSU3cg9ri8twBru5cUslnE
K4GiXJjE32tgwvGsQstwW+AjUibkhJ9o9fQSRGLYb/Hg+DzSQSpIS38YXw0k63Tn
5uxVyn11YuIHkXcacG7mCkXOpOHTGOHjIAgZzK42EvrqGnODsJxAZcqPmjuDxEbo
Vo+2O64+tL9gg30pziXwaRPEBAr9YQVTXr+L41IDeNunVrzHMaSiOolcWTbHEd4a
KAoG8R/UbEXTDYZ2foVlAWC+kCcLDxPYe/d2Z2U4PnATsZXpQxg17CGyp01vjW7Y
SnNEhXjxSSQByWN0E7cijuVS5CpG3EOdJkCqK9aiLdT+8TeLhLhWW0LO5VmlrQ8k
vImNFybSqw8vS2eWs2pno0Q0p/2EOsgsoQTl3j9kNB8Zo81jLkECzBqSye74kR8z
EkZsOC680wtFuv7Hj5xTIaBgsJH8jhfOzbWkDyu77fquHjSmNG9MGQ2x1/Od7xbm
WYq0fbb1QSktBPBJw2f8UoiXBquApcGh7YcZcShURatejpEcopx1t8iVSlAotR6z
/FpvvcqMQXWoE6jl3Q7MHXCrit7Piyd/te8ITQDOUSsO90aEBKdBpUu82NRbIooM
mBYH6KJudPgMK+YPHmgNJ5g2OEdmdJS6X5YJL40yG0VsULRvCEW9+4hQH2kREaaa
F+img0WWXd9duPBWiOdPtF0KocJyfv37u9tbdIEAbTo1mofv1W9mbCx8ewUmDni4
F47Sl8zlAynqdb6wvMp1JYqgc4STa08zg2OxKfzkdrzpDXs+kx91Erk8LXr7Dvcy
Dhy5TuRNJx2Fz0N4Lr9CY20fC9lBQsD4ztK1PvWnsR7WotqtO3Liq+EIZs4aboir
zO00NSKfooLIRO//ZzGMuYreFPd6EvraZapWtJkVGudFF/rMnd65PW7k7ZdNdCIB
NyQnbHwyr+Xy9c1jzCRJVwsN/snfZt1wiYcE7jgDcMZSyz+dN2UzTYgpEgJxW2GC
LQ22cLnTReYOS0T4idy6eMrSGa5/Hl/8AmScFZw0RhG7H99PV+S/+dVdpV8v8pl6
sTDzv9/ZplhAzHPZnEPuezc5ESoaFv8ZPcJt54Zm7OVP6LtJSMxqpeqmNC2h+hOg
lRHhGUmYImbRo2uasE1oNWkx0VEvbbpLUqdeM4sGFeIAFzP6OEGeT4UY5qdW9NSg
w8JRXPByZDTnV0OnWgNF8129RNz9kee+0YiJFTwVB8klZMqBNBqFMxjvJm33fwlk
3Qj1POdCIgCRNrKF/UEpx5WipKUi2EEZYdqxt0ZbS80raBvLMyG+sONxQggIBRLX
GJZ1xTxsFFPZyKN2Vb/q9hw6xp7gzfXRt3abtuT6PrbIQBPYJGR0RGZQVijNCfVY
x31t2FgJaGq1vlQi1tBoQjoE9ODZDkioZ9EnBIt0oBIyIGVaPC+q0nWRU009GMjD
viphtdhY0KDYA/u1SiFKhO71PW+uQYGZHHbu0FuYRZ4HSuf8gAmDSQmnz2tJ8mq3
3IIBOE9BmOQ89JvKIqqxKZmon+5DhIT0QegAOSUygzb/M9/JS2P0GnnhJ3F2953m
bx1ahnLGV94mp/xcw4J94UHtRZVsXWsLd9M6x4M5dTk3PNsx9HcditVxFLyRGOrA
8j8/i0S4rl7S5Jmweud7GotQYGybFDM4aKFWiw4Z87W4fMOIgt5VGRSWkiHehFyF
iLUOiBLyTbSIyXqwkmoLo9j8g0Oqef2kjYwLeEo1vXVfXj972e0pjC5sQBCZEh6I
Al4h15oU+DIdaKReIUUh4fQ/3QUiXVnh+5tQFsrO+3xBQ+IORjadAe7i9i+t+wZc
UcnWyUdGSeXIlUpUOU3jjXG69wrx78co5XtFRcw30Sx+x+YqmH9RwpgHg9w/fGkm
v/36thaadEw+SzFwO0j2F28eg9GVE/JCp6yrq/OLCZsQs/eO5oxL7CO+5YsSpmzz
ZkMbCbMxtubo9cqCjteaCnPr/dJmYal09NPzyNDmBUkS6qkUd0h+Iy0VFsC8CWXY
tTKbK0W7bFr3DiE/eOxB6anH+27Z+tTWRPCxtGeJhRSA15vowIHeAmfyj8j6GooR
YwoE3pjUGXI4bFqqkXrl0fX/4p4qb+TEgyITsbsbExyEUMBVXvgwZvSNjnQ0ih/+
1yXxKyN4oWb6HCWDCCL2QjxZCn18DVqAi2yRPzWk4l5uCQBaDr1SlZHmDI3TAUBK
HOJgHL9tJtxySrdRIrtycrgkufuNqgVluhWGhjn/nfqNq0Z+AqGwdXIwVm0QVzR9
5FKwYS9dWL9GyOH2Z03Cpzsl9VGMCHWyiMjKL9psoYT1XtSdSoJHt/Lt4Jik4Bh5
LbB5gmxdNjB+hP/F3xqx2IoJ6jjC3LU44qOE4g09koWhd2qbBHPr+dnImuEec9Vb
4Dl64J2QkFmqgtePkjJfazOm/huho9fZ/vwUfycx3ZA+YdowOLjLE8xbF9GbEWV3
gajQzju67vT2ZtKsNm0G0aDkBAFSrzRItkwBz2IXO1ZVvwSJVeEnNP1EWqNIzPqm
4YCkLg2/Ua9bcZ/jl75/SQkPVonpGrDiyGA9wOWo1AIwBsdBDs6Q/a+soeBwkzn+
5fECQBWcZfrOIY/noqdm4nup4YJ0bYnTilXva3yhZ2ArohM4YJ+kNjMYMa5AgTlL
TUmaqJq8lf/tTeJMpeXGmisS7d9dy5jGPcLMOaWGoWC9rhWB9i3+t0dcikhiyf51
0Cp2hyMYl7QScAeYJQ4k3eI3XSJiZUerN1/eti8BYgAGBnaACr92y5vjK5s/HBxT
7HRWJBW93R4rut7ENSk/8PH3Vado9j+oobAMCNxvXPbxsCVy+ffOdiwiOrWmRZuu
UE4M9LUcNt8cLZ3tp16OhZr+7iARjqr+lZL9GNTnc2gxc9A04eM3kgyKuR7Dst/3
bmsydkPSsaUMoFzBMijgCUEnBobMrD9SoqAg62n2uKbNsQLJOf3gQeRdX8AlqfIk
NiQlj4tSCt6eVIBSS3SpD6r1Yvl0SSEPQBKodecynaWw0eE4nlTxJzbuLSAEEKoC
BBojO58efUbWZIXXssxMFVYD+6I0mKTDcWO3AuuUCAjkHSiu6rQBvFjpJxdpLF0T
i4KyxWUCg6if/CbGDDyE49PUZDYhdZkq0Bi66q2qh7kaiJ5IkjX+qio+hT7c7ZHA
agLw4mfmTyAS+MjJ5fksG1zwwVLEdXqDzKfouY8hZO2TsagrvQf1p/hxNnFjTwRq
/6GLH/IgSp/PnHGaVufArhzsvNm5dBSe+yA2xvbRXVeduK7xv5a6pdDH4EykhBVj
UkXGWvFRHo4oHBSVfPQJt7l8CziftNWum3b01IK8xAsQ4rsVRKxnY5sDltXUUJeD
ULg1snHVNmE+5arLzZjFlMSK3cck3+CiZ9cQV3IdW9vISIvEtqZRcyRONsKHpgRb
EPj03wBtQxzBPNWScHB55+peYZeRClNUDyJ5X70gDO7sLKXRp0vFFPRFrpKpJmxg
x0m3DK+C9jgbl0iE4/3d8qmgRCVdl48tO3lPOZccnXxqgEGd3XVV6aStZwT1rtet
tK+TK3YyWTxqXiYh2bcbHj+8AKZmDxLxj2FgcmQjDKDtTjWLU/g6v0SXpVQFqqZm
5owIS5gEH2llAVKvgj0neMrlk3ptirch19Kb3EKBidlm0RdZ2jcVbqI5SioM6LYH
ZxFlo3owpdlup9sR0RGYTHfo0zVNUrAiHWmBZ2ANDEDgM91HHI5FW3zql6bfP1Gq
MkQkkFySkZuJOTGlkIPBb63K4xRzBVwsY5Y+hBTv1B2MrtChyjCk4DLnAnsNN1IQ
ptuWiHhQKbhXGHv1V44pc8nLB/GOoBoNtmU4bdYzvwB33aK7BPYsAe6thp4qZ4C9
yOHmrJTiMRU14sYwXL7L20p0L3DM55zVcAqSZz7j3YfINhQrkiD1QqovI3gVicPt
YDiIgOL1PgfGbcjCwH7PILVyPvtsk8KdoGIs3wfTafqtGW1IhAryB/tlPXpmQ6PX
F6zEdleTJtuwTVXQaBLLZ/iPsVp9dtSGlUBpblpR4Jcu3ZZanvvG8DsPgKHhzbav
I4y2QIQfMqW1UBvNJ24NX6QPgD7iQd+7tCcMogC+61aIh5HW7g94OLXed2GKrqEM
ZzvIzEN8dZPNHkRBzU5hkMYcLU7Q6py/NA4TrOXV03Aedgw5cX4d6/Y5udEGn3Du
SlG+H3St/dg+GTqRxTp5F7UjWVWCWOc3v3q2oEx5rM6JDIo0vrbGoWv2ekZfql6K
f1BcBp0a61xTa/sW+WNzQEnyBFRf8UbSt+EOMg16rU+fxeDLTtiyXooxxlsRUzrt
q6ROua0mvDBY6oe9G02u5id+xMuN6zXDXN6QebqvXaw88QmD9mh6JN3btSDyzQEO
Jb9yAjE/25Qc7cwqIG5/K6IaLQfLEohJVeh+GLJ3JVEb9BWTe9hz0Z0EC5PkAX4n
sYMoeJ2lIM/4TaNMlHE+OLuNIGAiHGY0x2ITJVWP5kZxUwCRRdHTGaov2Ex9SVZc
wV0ZHId91Qd5U9JhO5PHcCEglbXVGdzfreGD41g3fKoUFW6KT4PGqlN3Y2jFI7St
Rtx4+c6E6Dy8vgKuHcLzkx9aP29D5vwmQvYhQ9xNw7TT5K+RnKr3JjyU7PxFbmei
UAonMy6gYveGeSwsRQG5/r7svtkPgbwO1UfJqIA2uw+SQk7Qh5M1xVk3Mhy4CT+s
F283h5pusFMWDHcCvuIGNbumSDGVlJKgzmFxH5ccgqKEWMhqPlCjK0O/6gPHkK0j
QX7YdwU5IGdinFRiVgWHlR9my7a6raB1IY/LeziSUdFk7kD4+XqYlzSyBOk+Blqa
/lsIYQcFCmQ9BWDei29nz45H983mi2fMhUzXr8fORvTHl5JDOfslb9kzH4CYvGt5
AJcJuIlk0rgpqATv52pB/gwSV2gPWEX45dRg0K0OFuO7b2gi4pEjK8+MKTBLSb85
WoeACqBTcFdNDp0AZO6JEA2RedD6gOI4jeC2ENL69M8Rpn3zZm+QaaGG9/n9bZc7
7cOhSIU57MoB+fVocksqglIkOcZgyKBl3tNzL7wNDirl7V4+8vNvk7owxy9gWE9L
GLapmJE/T5h5U008xlRexu8iXn/2QqfFN7oTVgo2Mn5vW8enMbxOzZQhEpF4rUUl
t1P+j0BcCoeLnSB/zx3uia1mjPpu3pkDqRsi+mIXCmTSOlVOeAmh2+hStZ/52xUt
2uC0LJNxBYYw4xNexAbO5auSkoryi+iqxckzJBRY9tNorE/EQaYCn9xmFyOGsDvc
U/iSyqlG1Oj0d/g8982PxawOWldHQh5jkvrMuG4FCG8TknxWA3YOHj73IKKcuj/f
05c5ZGvVQQbxXDXdhymuEihY/oD4U6vIurrGho7Z9qoJZ3zu1DeB1YoYKWWSOf/B
ab0RTgVe0R0Dh07lELiqz/nRZsc0klMZpB6jgH2P/WnymQzppFfIJdap675iPto4
Jugb6Uxv7jlS19hpFqA8xDD51U2ZSVK9kOURR+k2MQqzZWu6A1U5Wn5GLR+44AmS
5uxo2HjBMB+cEyUt2dTnZ7t8REjtCtkKGsVqpE+RCenX2kTLPfm3OWuGFXYaTfbV
qd9zbcRKLwus0ET6nxSw1try1XawfbD8ea3qyvB5USZ4YVPq7zUj84Sr985PkMaD
a/cDnUle4OwCisEBg7vuIOMyOk5yaGzLOMNgyS3G3qcbpoa87wkKp6eHYryZxokt
8Y5iK4ZTW+uMBDqaZ6k7IPdtDtBZiLw4y22C5YKfUOi89hUsHTXY1aKuCjMYeo6P
DiQ5HIg6tHs0SsLvHZB3mH9i1Y3+7KK9/r4j87wABObnDTjBjHIdT/pO1K9Jba8o
p1oUuba+hmSWXnoOv1AtlxIi6Pc+ngtaSf1ckufNKsy9yGoOnlpQSU85YdhQy7pP
VeK9uwCZ/Z8OjHLKShcjAc4/DiKwo+oiRvvmJjM943D/Khh3W4rDgHVhpqbDrb0E
TUxKy4KlX12MNoqT04mlq/ckTnf3CdnSd5nbyXdKOyLrp8ESGboScAjZfToVunSR
AKn7qvgc/SZY7A8YyYgmodiLzSDAZuVxYHUH+5RaBUKahcN22NvMMUnRZCjO82pf
kAEerlr7JEJkC8y8wsLV+hmEqh+vq842RL3XvQTNBdwd0iIHxvkd8waoVP37vZ/b
6lvsgZJyGXhSwV4oMyMWIq1tUUS6tOgGt+L5K0Kpczf7YF5gJsADVVQbh380NHkr
qBu3SJMRC9bDlUt9oBVis2EOHAxYwfWWgMd2GVKOgPg1/0UnpZfQnn/wXf7obSQi
yJ2WXADdMw5qJQQ0HOHGl9PKJFqS3pWVcnv/O6z3oolZiJILE817OYHiWnqcbCxB
Vpn0KMSvhTPusUneihAx8S79kw5VQwP4yQxOEDPa/Y0YEtilKoK/KnVD1baUQpv1
V/gIj14T1pGBFQj4YO2DuNBHqS7YrbT3+VYXvQblw9Fzbvk4oCdwENsOlsa9Da0x
jmh2o7FlOFSG/cPO+cfCnICHsyT0JVlhADLyWYx93BXmXV9AFvGZf0bRab/OhAQR
coxFq/b/18WRyLj47qWy5C7I0tYLYw83+LBk+kvGh/B73uxbDp7vvbTfa7dSfVEu
bMjHA6Nz1I+zKSusEKxBHXeU3gAigHuaWcfejz5Zqcreg2vl6Uue2x1pgLhB0EOi
nSv1+jIoWzFnnhFJbNYz/2nUtRNsOFIP2RnG0GiNpn16eiwxuFJynpf2RahcG+zv
0KKOcqMTsym9irQ0gPDzGlQxIeOkFrhkzFLCz6bEZuNOGTRnj/BALGVeutbMYCV6
XPQ6vf88AVRFNUwzf38b7XVyVJh2QvYm5s++bnXspqpsNjui4uK7wK8W7l9fFIi5
UdSgZN95vlJId8FmeTYiaS+6Zvsyfp1soGchlEuWlFGdI+oFlPoiRHyCDnCYYFIG
C12ETfZugN7oSNHhf9nAYRgYnkJY8Y+lPEf3WwwnvhVmPMxc1JR1RayBJiyFQTZE
jWkFZ44NNxQHoH6ujlov243/WDFv4cn0UCwb7t6HoiQjTu7xLqXRpM0dZ+MO1UsS
Fv3yrPidioJ35FUKeGe+t/L+i0rLgnWRSPzznGF6b6tOK4jYXu0CRsUUQoWHsV5l
U/7PSOaux+X8m/w+G04VeyNvkQUEMD3njlJcjbZ1UIlBl5uBDBx+4Pk2l53NsIVy
mmcgMXAxZQveLS9/AXcdhEUh1bnvevUEOGcmpbZYxM4FChot97AtQ1qlc/c+4sjz
J8kwjuQORH672vvMcFz5DHXPuqhGRdKP6DE79VDjonuSI/mJq7JAjnteeEBdQx+s
e8iZXbmlmvDV8RCFc88cn8m2mgQMtoYvIH1EP2trOGvTpfC78P3BcxJSgmpHKJrk
HPp7auIS7wQIfmJwRJ1vn5M9h+h+ut+AcDEcdrGRpZFG68wnMulEElGKxQyeU2q9
gmt+4l/z/O8ZYkslmKOyqJi7l9hXxignCDl+zoPTa68sgENuzZL2+sjRCJ0eu8Bk
RkfYGO8B2rJkwc83POtCbY7JHPIc11RxGxt1rHC1rQ7l/Qv7rpx7/A81fUl5Khfy
QqRvbKHIToZjAvQx+kU2B/MtGwqV/CxQPFnGyzq7surnuV4iM3bPkGCw0Y7Va9+U
9VtxzRExXaBwiJnC2Zp5QI8FTu3odn6dQhzFRGfRoB8PXaeaC/WpXhwrrjvgp0Yp
c8i3HKGpgDp/lZXTUfT9Eg1sflCMwRJRxQo7RfUidhhYZRly+iIVBdtztGnUq48H
Ezo9V0RWijq6NeObMTvYYMsVN62p1zQDZ3FimEgkoLwTbGKxq9ukYZ0hgO8Vz5Ma
/t8PVOoxXpBad+Zht5LLAedFGJUul3gntFwmhFd2ZQHfrOmKY33GJQSOdw/1suKB
Da5wj86dXYeGbyooXdfAJqpjZFybACpgSYUreYJBUjxXlDaqh8D5htOF+sztXSg5
Q+lOoqVkgl7m8ayC1IeVznaJunAoXsIO60jLlV0Anvo15pkvpWlEFb1xnjP1rT44
KGavHe/sNQWoRqlVrrFrdXqBE9XO0jaeMViH8XfULwR+hHuxZqXDkbfUrDbqwklZ
DIWFrn6lh3EFdksvt0XDAsvCiERkfPKFXAHcyJfespqXWQvG8V7LZJaikk/PQCYk
T/1f/a52BowIa9neYI06GLudyG/DTfUUpHptiEdfBfI53OvuGAMs9I4VvqoA/xUK
SQU0ZJsjTg/zV+opO/z9kdWeuBojvTtGrHokveownCqq3Xm7N/TpCFWEXxEUshiC
res4KDRwiigGtUMYFN8lptFD12XM2nzhbj/V+cnM6ZMmsaJjTPeQkn2uVq2lBABW
aa6h9YUuD418HhqUrDYNIfg9jhyElwkUM4Uy3aa2JpRYoGVOmdyFM3tFIrhPdxxf
L+hUB77uKK3OqFzm36XzQWDMjw56tJ4QIC1eSaUil7N8C637X3k/Bnb0MzsG5T+y
O/pV2b2BS4yglygR/t9qQVYa5BRNRKdO+pPcWZSsQ/4eguWz7apHEQMHa0sG/HSs
xmTugHkvALXj0ggDqy8s89ndIzxNWHljBGECWVvJt5fizJOR50qfd/BWT1ha7V23
GfK0aE7wr6YneUtdkTMAXIL7cmrsmhhUScDRAQm4QQsPzX3kjaJv4cQcrnp+5Jzu
STpZ+ZDiB5CF7fjuhKKdRyekaBke09KtIxDzyslaITNC70z4/xgzx2hxCuXpGwsy
qTrvowuUpXALRrW2AdfRIEzh6NYFe02XcQvX/3S8aP2NM9+trlBGDDqmQe+TlO/B
uFxYfEk0QT8P3ThaIKcjLHbarNt1j97ngutQpxvPDHJen0YgCStyeXLijOtMI7W1
Dw1k3lPpbOmeTDHiJsfK8XmMA2mL47tDJiVGTh1cq7uJO9lv0+ovpgB5nZvogoGr
VYCp9neU/JWpy/fJOm+ZYtcKL3Zr3LEaMCSCHr4jryzUNVsrrApmXdDAlXDl0EhW
MMtTfIE7pK4uUQ8Crq0HerT1nVMdtYyk2fzwZNnn/+13FaojM50nVp2vEx3JLw3n
8bHBN9GdjXU8j0WHv6WudDut42lK6y98HP0viULiLMSH4Dlas45KEfpvqe268H58
dslkEuLojrq3I98G0l5ha+3mGBfiHYPSXtksTaDhmakI5jW6DEPHkEZrqsZOld2A
uYOoNNUU4OcaEuLvhOUR/mIAZNvXcv8vpIu0PrLQ2dNZjUEoLfq0ngZSk9UFsS6P
Fwz8mMAYvppyVlvruzErf4kEkKn/hs0XqOFVOw6VTTVv2gO4jMKv/fuowvGVqs7Z
GYCjZWtKgnxZE0eQBFaH1g2RQFYqaWE5FQbInwTXBjy6yY0XX7RMwUb1+yaMpkNf
VIPx4aKIGUGPPALckHT8yw8tEvMMKMZVU71oBOYDClGKQFg15zWHPR15dEY52ZT0
4gtGXp7D5fxqiTOLTqnP2QRC8Zii39crY2L7b8HBPiWkeTvqjg/FklrlfLExNv0l
KR2v5+hn5QpPSnNJFCvzuigzMrExbSpA7xlHzBAVES/1ijvOivJXrYgKnbehSia6
ip5txio9aIwDvrevYjNgBtd5KdU9NChtq4vUIk6VrNutmgj/mP9DFB8P3q8IEy/J
T9LMCzBp1RnVUrZAD6RJ7emsaboYL5x73usn00H8g6Qi1mOA4CN7oO4/lpSeQzTo
hBFoO5DSGjzL0/cCY/DPIDw8c2+phaNW1dISHQ9QlAZ2CHcH8LqI1DxDNRYlWRKV
tUVfSnJkB6wXNWfBZ4eC1KkZNtz5Vcoy8fEx9dNroMoXQZqnUIPjzjtmoGwtExEf
RldPWWf9ObGeHiuUEjkk1JDXk3HAaDL08Tr1NwBcN+YyA98GcTzfzFAoFFMPkeXh
u4VxO5Xklb+vhK0G/WCYJ64Rnqnzr0hsFS5DahKWSYXP30zciZ2qDyjAoi5ZJWEP
s/r2YZW3svlkCNIA8bXEFkwWIKbABNsBbgmL32Ifz5TxtCgMh2y5RKm/qvGkWNV6
DmCFuCwcKAdLwzLp6wuJWLR3606c4SEpObUAthcl0moM1Q429J/ukCkwd95s0JfE
JLTViHMG5rvOVybzuxA7U5fO9LfL5I3OT7uSsF8J1d1JdX6ETSfxG1nQ+9H3EaNx
UrCKCJN5BiPSFIDE9dNUfjYNDouuZEIyJB/I7O8K+YfXK3ZDvmgtw3pQKkAct/kC
GQfYCyN6ZoZAKhyiRj029/RSnMLrgnVAD5VpksQOLKXk2Cm/eq7zIGRu4va6jH+r
mDnUbJ2hD2yC4PRYu3unGpw0+Abefs+te6+Meo48s9lZ1xo4cD1GPBOb3qPeTCxe
COGxvCPk1QrryrP9SpXh62I2oAotHVsBPm9ThaI35fRwL9JKmPqlxpUxsZc/8925
8KcS4PYHPkDTjsk99Fwx9/oq+HXy5W8wIt/ERJdBC1KVDg2NkRkfo12A7/oH1SGJ
cIn1Kfju8LyRqMReeAUsEx6rvuOmQPVIOhZwT0cXFtVFBKK3pHnmzHw9XQ65PpKG
As2uoRtzNCUQbpnkuJbeZERqjJWcyXCnhPe/YuOhZwqXe+uU6cNH+gL3DsOI1TLz
LlAC8DquOH5jV8acg+6oD/DIml5P4Jsc8v7aAbHgjWbcCGFDBkP10aHvjiUaXAwi
e2uX2Hxg3kajk8JYp3gxvxF+ReERkc2DCaGE+KBLkRDf/iBqDtbdjgAOF7wfMKHx
OLAZlHNLA+so3IeS/r9cQBoPjFmhEtcCZpdLZwg9hF26/9CA/zjksiBL9/6Lk9bz
VlulCvY3r+3KTgzDQL8MGOwAEjYhMudehTrWQpvdyeTw2mpZO8TQ7C1tGN4B4hqh
M5OxRaPIyBtkgyXD8Tc6FDX3tdxK1XUVYzlR1t/fcMBAEuDM6ffxHtIyl3KHiML3
xxF98pNUUxEV8HG0tTLT2+IX+XA6Z/E0fZ9+0i2552nDDd7VnxqYkpoNbZNa4rG+
p6RQUD7sdCnxGXA29CXV9lbPpgp3mU+XeEA4zDVxjqaqVK2r4pS2Bo00oW5jv1av
N+JBvV8DuWrCGlXqvHJi22wZ+SuVBbdkBR+sC1PlPryH8Zq0LnNa1OukiTCmsFZH
XbCri0m/RGIfYL9ZfRASIbDdUIk12Oy+7WYtqx+lwb4L9Xeh7Y/pCC93X2doGLgq
rW3+iFeWyyHjXysP+VoqMkUyQFzWkYe94hPxWheP7LTu0QceA5aNmwt7fYCECwgf
TUj0UgVwfu6WFHZxT/4losVaJqYiL52v3HijfwKKWhafeuMlLMbNnvtJ8wdq2ccy
auO2J8meyXM1QKueAsgxbS46cq8GPoYXxZC+RSsFijBIPV5XpbuPm7XueHloJ/5z
eoyHeKEhPLSi6xke05FPc+fVcts8TOEBXMQkjtPsxXHxmLOu1CnMun1c6DBYAZ0E
tfxltDvJqsd/x8NA/XV4nn+dTAClRACZg3eeP2ZFxvhgoqYdBjCYscfvvz3a+rZc
UnruHzZe5Q8WNNMQiejFtw0npEVi8Imuj8uHDnA5/JjswoXbj6Ba/A0w34weaBVv
XKcrXWIstqB+QpjcNdXE1zPVmYubB5S3zc/KG5ppVRlaMpwl5L+jkJe1o4PIdm+5
e0djADMRd9tz73jcIraF485XQjhGYQJb+VRkfgETUzDMRkgQKa/I7WJ+QFqdB9zL
tVCYbV8a/UL4UtGUmRbsktq0pzNkMU1U0okdfHytkdc+JRHea+JbvcgieDrhntTL
tFfKsPl5MAIwobjLkq1mYUvlsAlPNXTLr9ecmkONtvykPU+Ha0MGOeoOrCs0jwnV
M1kUJCMYZyxBWYh30yBeHxyEHbE0aLso35x/TrDmRdVtJEBGKEJ23jbY0PjHpchW
DQ3ol1nB//9LbkxcNBS2coh6hSVLEn5FZTwHUqU7SjbUG1FKzjpw3cDz1SoZ/xmF
ayolmNUcOFqVZmPzvCTCK4bUzMQW5PODSvddoP/mYGeW4zMLPSMuq3mvi4lO/3g2
XDFbIIeSju3zI2+t44n6vWSL739kDXaVxe7VURvhDbSL0bkuEPZCZW5ijwRVuyHu
gRUtcyYIK9JYajIfM+nlxNGw1L1CK3z6397kVlJTACWXtxhmI925NsD0VXqoCiSi
5XevrfHVnB0SPh9wH/afep0RZ9+cDV08C137spaEcOdgh86P5g4UKgv1E7T8ajAf
ZWdkNlfzRe6QEYESxHSblW+GL5UWbMVDcYV7V431wm/YZYlLQ+313IaW1J2EOpB7
YgXu2XTedN/k4X2pJMmmWsTTBK1E0QHMMeWBMP4uYwdExBKI83EtItURWYarfy2P
pthHF3Rnr0iauy4Nifs5fvQMESVqO4DNKPLNap0bh0PuyJQo2qYmnb9i8jTq5HqU
lA6r4ZymsgbbKmtVR4kZkv4kpAo5eWesgh5v8GD8EINfW2lDoYrpQrdyASSpOXA5
S++mPTVmeCRAgfrLjueC2REI60vErti/K+DkePuzIT3vfS9WVo6diA1+P9D3j4IT
uD4R83xbNR/EhSmnj4rhIpEO3M3TVnVGZ+hAaJjBLRnY5hgk/eDwr3SgAswgyHQs
Q//QJRBMggDn5lF9T970lYmT4bDhGjviFIzuUcWEu9GnRweryi7WZ8MUe0bblNXl
MzLsPB9l/zMBAH3xVo81SNa9hZ8TOS9/iy8qPU/fF6n/31YKqItrX4tv3gTMS43O
CJ3ALD9n3OsRSbjIlcmf9Jdvb4/P9NeN+kPr629RnpsNpH9qeEO5QwD3JcvG49oW
bdjqix98QNPUPW2JCRDpznKvvmucHJKUu1jQjINMw7MWDc7oyIfokbHAGTI+IpnW
qsm6j+sPBCfo4UE/ZwWst2ABrwxi5PPOnglRFk3VZrkPNhzlbyVZzpudyu+P//Mf
G1zaEUTX0wKccBLATv5xtwUGkcDsB+OM76WVitNApdqfyzWAmC958TSZICn0uk2m
+1/D8HqczhKrbXpMIpQfrAs7ahTzscXNiHaZ2xZ0mWKjXRPkAKlCiQttiNXQx+w3
YrgRfeLlbGX3SEe3vdsLdAqa+QfMXIE+UfXbZOuzn+0EzT6Wv+GX3FjD+An088ng
LBIB9pqZ5/M0n9EIeuhYFG2mn31+gqNnVmQ30bPzDAY2nHeRrnx0bM/lck/oTBoK
Uiax+aqjZCs1F+8M1y8ZwhwLQgUiR+LZ9/YFGJibBdvbgm80nUaO6F4ZEvLkcWf9
H0ZU0XMNh/7sqvYOnL0t0UDBaTPGYlVKqNRlVQaV7n7jfmAHftBRuxesNgiKUBed
OupONxBzLdfQBuugt148+GiDyCEFqdjH/ush+Ln7yTdwoX6fvzUp5uCRvIgyxWAc
hx9dOol6Z6pSDrp+Q26XyHmdE73BdvRD/t6llSshcpkh3unMVwSSgmbY9RSepq78
a+DIb1E/TN0CDNJI0rGSVDz4+uFEiHkbRt2HzSjZFaAq3BDgiQQlAmEZlD3jpYOO
plVoVgRz19UeZUXrT2AB0wcloSSGFEuRdCLjd52hL9pnOX+TTv/J/fk8/0XGzvxi
JS3ChDi3y2MNtHkiSEbG02qLsQZBdMQ2lGe1IlnNbynhCxRFwxpCsOk9IBbBH50V
anmtd39EZatckJbUifdgWJrWQEMs9b3Ib9jXqYTL3BUWc4SnPn7JGbcZ+1g1smFS
7JQ+UZirRqw5gGsuIhOXVf5M0kparlOFhGuYJcu60RYIsufKZUU+Ht5mLTtPLMum
wf1r8luVgGTFaUa3P+123aJtxivd3Kl6dWBtZ5wxzVs1G66WKNxXEvmwJPXDEv2U
tYbICIvF3AMZxlJI84llJPzs4Oi8vSwMJMZg3MV/duhE9z7TMgd/+DH7Oyjf0gj+
sM8Rh52Lx3hwVjr1KZiHrjD9E6d7BQe9tbgshStdV0w1xwvP8vPBSHSW5ls6fheR
p1y6zm9gMl9ib6SCzWtv+iHhQL3UI0bOkw03i52gcFhvivNSx081tZ+36ow0z8xk
N1+mmCFC1BUCneAvpKr1fKEqJgFsd3IZBbN9RxtHvwLZc1LIqF3UpHTFhyJBcfI3
KwbXAUyt+OaR2XnixPFyvUNm0B2dckCzqNXA0QIESkhi/LMFDNbcFU1bRH8FIHc2
hFltFCzlxfFmHhbyqmIe5yJoau4SFSmSJREobrMBaYV8MVl7MLubm2ITBKE887I4
WXT+UNjGXoYOVWdLXDkubyMOxmQq8Zr5quhRBJgFiJU/J6ai1uctON8JEqYts3DO
zvkKSF/wbM6D5fBB7leG7IOLGTdC5qW83Uv3KSMi/QvsXxi3JCS2T/Sr4Ld8sqQw
jl6wlu1J2ZDP9TwuNmUB3vMQUFfJ0b02QhFyE1CSAkm8hR/CqU375VMzUzZnrANG
zG/RFFXPqCGrLFmkfyRWLqRWw09H6jnXnC8/kQhtkM0TR3zHwIJ0P4NrXl75Ba9f
FQgCcDNJkuslF9wGgirAatlqTw6C9SuGvt5IhsQOvC1weR5J1q2EykPaE/+JqtNe
uJmsWtgGwcuXhZmS32witD1cayO9tEN3wjH1tn/tzOomLtE6PLaqaUx3s77qfkBy
2PcRjPalIA/oODG899G2Wiogkj9jo9ixa/ApJo8PzYrXkWUg+wzCt83rM5aXTRTp
MFpctR3FyTmhW63qACQKBT/74Gc1W8kuQ347neUJTEc6KLJQvqVLit2r4HXiGZ9/
4JoO/Nem57E1q9mwLi8kSvv3vSHwzABHg/Kp7+Gk8vLPJ1K62QK0DwvqhQlV2OH2
nCaj+qR7+iHnSV1xBXhoq1sgcp+9RYmVTgS7b1At5geCyEgMhhyg8NRDJhriH1Kx
lCwF0nO0xeitRhz2IKgnD+3tnjJGNN3FWzwr/XLmE+rVgwQtjq5i/gCJ5BdQrRrc
T9z7jUkE2LhmiIXbiH5Oo0lSNEHDe12OGKyG2lVL+RyqsbBNYENAjE15j3HOS8+K
Dh/8xKYiM1PammgjZOUIbKeijIqBz69xERy3uIff5osQWEEpk5ju5RVuVGXGhGVJ
PzgFXXy6C7pEgi2DKtviyH2+10U7VRfGxNZFYHcDsCZ/RpJ57do5mJ2wOxVRxwsg
Yjy6/0d6CEI8BGSH0WwpGZdyr7ig704QezmWykFOTXYw8VUTC/vKcJWwfEvWZHJT
8QlKPPQa32Gq20TYwc2aS+GkFlrHL/3NzgWSenNkP7REsQENpZ+4rCN1n1IZNIy9
nPi8aag5BhQsvswEXPacboST0zcDIHhQjdrzD3Y6DS+1A7MhTftczu2lRn3FGoyS
VEa2DIi5s0W7aIz1Iapyoqh3PVNlwDGH4VZ48I7Qe8CxCXeD1RUSO8pBUmWCPIxv
QA+NW6y6S7epYmmuGtLJ9zbTpk1Btk4bYcDLJ7o06XthVewzJXhU9ufcp2oJNR4q
rF6o/HWBfrLIkJxBrjTEQcNmxkv+hNdrZX4L8NzFnmyYl3ygO/vOSerRjaUhftCu
75g+3AsKj+LPlxrnPLJUZEFFu1FxO7pU3VbZ8Z886/MgTXLxhx3C2i6xcVRAdiWU
6Zqn1D/uGcZAB35F3CxZPvOzpXYVndTHq+jDROSIjmQqcKsgcahfCC5OegJWR/Sy
Dm173kGM4tZSObtnLQxrPX1/cBIdF9/q7l1BX6CgB4sMPzCCD9LTEo47EV1zK3Pd
4JEwgzHnUPsDeEnlgvWmezruKbJFCuuVWxLjdyZIZJj9dUDVBJ5fonkys5vUMywG
V+5bdhUbEMdCvYiQ6bckddjtUyTd0K1jvYJP+uWDtUsCtIW+9vcb1XC2QsH4nY4v
ksJ3nhwe3SCmH8z+euIY+FQjJwqSc/DJwg7y5Gr7ym/fKDRNOl/tFHAM/subIjAr
VAYVFaU8V6zWTEbUY4wETSX6ANkofmRAstVwesZV8Sd4narI5syrKnnwBENVlPe4
JGrMvYab4rZ/2fVNNZi0bHSm9RVKoIIscOsCnz2hfSu0g9815/F8mEwgJrvqAmb5
mjDsQF3ErX4FstcffD3scCBF6wR8Iqp0mQ+owbQlEKEmZ2Az4zlsWkoFxzPUf9vA
n/5efmQKvddNh3YBFB+s7DeeiMgIf6zVOrGXZk9FCa4ioKCTJplPjIWeffyPzabk
yl4ZIs59qriSlU6D3dOjAd6yFxexWQWIbyjkxle9fPyE54D7g5cRYgEryxx0xt63
dRJLEbtTsCVZ1LHM1M7cYZoTJafFHm7hC/8OFi8TBZ2e3/V5aw+nSWR+jjhfEBI4
ujqzND2lrdBuccZdXM9eNaQVXlaaTC7nKilg+veTUfxe2x529ROUyvSLhvdAcOSr
wpH2CHpacSEgl2gJJMtM2pa3XBf6Mb6z862HE4pwtJlm2GLJHs4A/TMrsjFiesgo
2+cWIgCgK+bSpWDHR9/QFyZSGoEs/CuEPLDOIjH1yCIFl/bs7GEgsi9T1X68lOQn
MJ5X7GbgXc/bE6exmTcqRP6knq1UuTmYFXyKq8MljsaSR8BGy8aZ0AmdMILt/3F4
aIxuDeDTb1kWdWNfAVUkbUP0ZoNTYuKxc62zGVySkt13JiKf6RTQmhAev+0RoJp9
j9cfJlq0WOnWYEovBDwLNXYiqFO/DXjtv/KxLye5KSP0Fq2wpNJ8nffLbH+2lRKQ
A5DgzagsEbj/dVmisd27HGlPMn+PSHrTM0VaCScYbTsm+8RQG6fQHtZxag4WR9rF
reyvmj+vgK/znMn11VgvAYZQKnuOel4uHifsmXFG9rBBhEbduR5Nf/gGfp6msRgO
gghPFZ82s2O7Xx/h5QMxS8DPG88m+aFjWUEk9xBGRG5lDG4lXdVt+iS/brxBVx+/
wh+BE3kQolXvk/3G9itSL/QQf+9U/JCdf+BOWU2P+3ISlqC0AFRprZvBlozg+S3i
IdlRim/GlnKfE6tI6AxFHWxYZO3qPrp16O0soBO5gpbFCTLuCl8F008oqvarzwsj
WqevkQjNb9C7vARWUn3oQdHBv7DNm35xj0Tdn1GYKmkpah0R4iWVFaPdGvJjiCOG
Hf/b8k7lAK5rRCmLEj5syf/7FiSYcJ/m6BlI8zLaMTlIJt6x3fp7thrmBQyhgJqb
gsGYsR3eUi3vVFkXR8fly1VlESxf4ujLGveW+ilF9D5YYr00/F2SCeNdjxrc4mKR
DK0FxcFhDdHyPf4kVYqrvUpeSWpL9YcE58yyi6tvyNXzFMXsLxnZFvNk6jFvRr2J
jtvrjxEXlHDRZL9/YZfly/fPHCzADOFo5SfYP1h9AzAYVz+tkKzcJetYQ3CxVcGq
tbrGrK3J1NTB2+WnD1GlDaj8TBAcYILZJfaj/MIj+JYfBxd3xfJd4ikwzRQTIKGI
OhWQxnebh7HHc4+yty1JZmYkYkh66l2FP0laDxdAgomGt+7tDvXSCGxb3VmcnR38
DVU7PHVXBldxO0Ic1GVte3C/fJ/4T8vtgz2lUVDIJGCheVnmzKa6COJJr5o3HYge
FJ1qvi9fnI1L2gD56A8PRPu0uXD3X1TAp5OhMo6j1jyGV3ShiryAkJXcpzG/ZgjC
m6zRkVI9rFf3ysPT0TcxA9+4KGt7TcZL/rpE83nX3XXhqB929w4skDoRPLGA1zKD
9kr4oWci6CBDMMJLa7u1oaAfrrBGwTRii5on88Z0lJNuUIF87TaULBTaB02kGMcI
a5b0Cwf7PjbC16hJ0wFzslJV/Mce40Refl9oCtS0gbtcCAQlYcg41TEoQQKKeaqJ
02/egy90tFXgC1dhN6McBmTsmrqhga7kUwMoEk9es5BOa/TNjL/1dPm4sKMtWjZw
iBoV+Y/RZz/0g7o1nItHj3KOIFxXhWb8ok27/94XZDpEqEUCvQP8MV/VeEHifRE7
pQL4f5TVNmeu/CE7zHEMiEo2TlKRsH9P/+U9I5GQmjTLUpzKBM6HjUN1GbXsUlgi
9ibsyq6kwowWdYPj4sT5Q91a0uRkLO2L0P+O3zHzFlTKaDH5onkIbpw8by+pXAyX
nPlnm+Fd4zPHP3JKVuDCYxgo6pBSe61b6IDhQrUSJ+kvEPQraK4QEICnafe5h19D
sDsiWTBPjnyvaqJinINzgls7BUdapf/1NEgIZaScR2Nt2g1YIA5Iun833T435ZMJ
g+bwCI+j1aVZIggtWwxhcU4aBRQ45woVJlUQH9Oox5EOYWWjLOHUs0U33WagNxOx
fKSQqkT0/Df4vkYSS7ULuBQcZISFmvKKiIpXqALJIkZfzm9wdFdbY9TkcNdvR/vq
aQ7j/G+4qCYsNEv4OJlipDGKsZmboH/it+w+yXL+VBwyRm/lK/URDXdHueIVcM7G
RfVm/aytyA5o7Q6GXhSS7nT6MjEyBGRBGEHSpzUmtU0trNsaUn6geAd3p0fsSEUN
OJrHCU2flvumqwiUDd01QfSwNQYmBjo0wk0YMqfJlnRo4utWPTSVj6RnJnLjrmnz
P3bQGaqZNWwNmYwwa5qIyX3AoxJ2SmenGzoo6QGfXm4o75+v0QY9U/SEi4z14ec6
s8jydEe/l8N5yx2sNRc7GcB/RHc+z03iQbzfMUd/tGfUjgIe8vyaZzQLTh8TT+ev
VLJFVuoXUPb52fqqzGfMrq5rNHgnyPe19vmkx1feZvxbLnK11I9UTwsso5cWZb1+
JVCUJGphpSwUoMJ1ocMqNEzkHmISZ/ibJf1B32RjLzA18otTEXKHmpWvJ8ncH/db
rXfFywG/FaIVAVDETZtY1BY2TMoVZJOwOSykXm33g3yFoyNjZdwGLBSdJXz3bZsw
tJ6x3Q8LzEl5tPBpAqEh6p+icI80Mk8VImi07WnHPeOKxpHgcWvXZ2eoJuHA6qXZ
5Gk0NgBuKIJaR3OTyiUR0td75U3TYqsXNtMcgZodBBWG7hRYJLl2/OdLkLbwJNpq
pzsKnciTJMtZ60J/iCTfddOV2rDrwqswW9Hnf2k5xXVEPMPSO4zuWV3Dlxw9q2GJ
t2IfHMmCrbVWkQdq5xuMA5SmxQOWms4ZVJIKQPDgICN/CBh2kXs9+NqYtez4b2br
Wn5maARbMpyLoZrejh/KVCvwDAGn0jdSvIeWus5DRLBnlkoPeWdOTyTscuBGN4Th
yGRsRAmfMy5AHVsfMMs92j8JKxUmtzjY7nClniGyjqXcx0ji9MlwaWJ2SZA5gR61
YTdr6lyK6Y+AKaEDSJN28+WO0GBUQSyblcPC59XVjDjFwo+z8PXYDqThuP2YFIbC
DzlAcDbHJSLb5VWnHhGiYHjv5B9xeRe1+LzDFZMSivt4QPONtnSptEltgBf9tG4b
uwgaaifGYHwNJqFIMz5oSHp6LmpP9wDELkVPX8IOaOnluuZTjrAwTygu6tXtqUa2
CoY0EYzHrg4qb+bEMB1NfJqoZYlXtGptcS4zR8iyRTsYz/NqZ8X5kb9T9xiIj/ds
hQhdee+I/dRY1n4nAuBEGdAUxAcI4p0ofzRFj76g8lTdKb+w3QnjIH7t/6M+mq+z
UHvLyWx5Nci0cVHuWp2AmOFFaQaPA1JGXAE7FTsh9vrx9P7aPoBWpHgc2iCTKWXQ
kkdYgWRo93rXgisC3pMFKI/dBkPYjpazvYojWhFlB75X1aCU8OlA08RZaSINkNJO
pZShTbbAbEdxLtlEzlM6CdFvBVOwHwalucD6Yi7AZbdISXRVAKyCGLxQh1h32/QR
mxnBVLyiDxRrzvSmkOXF+3w82e5SjByGp6OFmxfguR1J4DEf6lBo2ju+Gn1L7Ch6
dsv6mzzeUSlTMMb6+MBvpemrVSUpBcxyJPXIHrU9nRoUyfuebXm1uRU484oB6s7d
g6pdon2fRaUXXQYs/SgvKoKXw9N4KMPH7iw676sA9RleuZSlhAbdvdXRWsECn+W0
OCr/rWQ+qalAv70CfZuLu+GLuPxXA8zMdzUtkLPBEhPVT4YEPDTMIzkUzwRinjbL
4kxI3aBqsxOtMF1MBghzEmO+Oqusd5Q77LaFcfjGT7SLyJH6UvpROl2HK+3XI9vn
jAvjQvRsaBlN5/h0RgedpdV/Ab+MNg7w9bIDMydEGtVWg2CFsWDsxY/5mkVBckBZ
NEOF8VFMOSJDBjVFj5S/x/mGlfGg8yIqJQRouDZrNrPzQr/js4PLKW340onNmKLV
PD+p633ztlryEsDpV6m2ihSLE/Dk+eLz4FSE8fhJCRyHgJWn/a3wg7VWrwcDXGPr
vcrZ9BMHLQw5z9rXK5SbBXdK4Q0p/Ug0BtsKrrX3TWLVZEVXI6rbDG3sv0MnkZg4
osxzzpUDkuwy7YHxQCrK1kq3KP+TWFeKwBCnmW8u68KXlNxm+j57Cu+WUGyFFQ2y
ZCog9xkSTY8W4KBta2v7+HToyLrcX4kSHmkOrWI+iQY8T653Zz0MzDZqdk6zcv2b
6PRqGMedvLi/owF7uBayhI3njaoRpzbeXmTLL63r3oHorf1GJ8/wFln01M91z8gB
OIFycnvIKzOEvskmM97hdR1BKeipwIYdyFamWow47D2ji/H9lRj1YPPTickgC+lp
93SfpQUBUnP3eZrL4OcxhBBnnC+nwllYqvdmMTHaIjWuVdQeh7D3YdrqZvLPAU5/
JnAGHp/WTiiST53fESru9DSwlHZUay/L3adT4B0b9Whk5vYAux/xENSQ7FdkEuDM
mWZSdzi6yH/SFXjacS42iGCFTfzVg8xtGrvJKeRD5xN0Ht+7KswmA8BOYxuV9x3N
9aqeps0TGHiW+XlAd2P8bKDuPyKz+B0yDlkXty1LXTJ2KcNEN6H4cKHhoTsRgYt6
iLBvbDxKrzVl8FZZG0O+JzhH6DAJ5I+pc6s/ZogO4ZP6cUQoDSSEju1P0xvcIxZb
oLRyXOdG3tkSZz+hH5dLTW+lXvipigAba1sjkijfTqT3VbikDCzuUXIkyrQG6g3Z
82138fKfWCFU8GKyYbihDXL5aWKMeU4gl8z+9I8yW8SQO1FIHMRYD7Svk0ImRAaL
hpLK4tvPwIk2MCWZL+57W6QMXbuDw5mHoVe+mvBrUA7GVWBG5lZnYWIT2GLFgWcd
bD7pWsM9eNwLEUTYSOVcb9K+bL/A2MDEHBmw8BPu9KkWckN+uAfrORzhmMO/TPT2
mFeiPru4pHJsCIuscFK3IRlIR+RZNLe0z93AVr5OdwOfEqZztTYy1z26ntoguM74
BAfAOr9MYFy1v29G1AaRiKbmKQiU0QQ3ENv3KrRuZyMmIfpa5KDO4Kptx3oaJOTG
6xQr5jAg27dOZ0ccP6P2/9VeVZUgtULxemqZcClI8gjb6pmcBFoiTbXScNCC75oE
lshtc03abM8clMA5y5LzAVEu0aIj8Fs6xl+Vy4IyoRjCbPh7V7fFyRci8vve7DB1
ydBSBYrIPqKD+kw517YWBuzE3eRUwkuscrsCIqtPYR/g+ALoGUwFT2F2Ao/lT4En
N+RN/Mn99dC63+HHW22X5lMeG5zG2SoKIJsrCEF5tLlw7yYVNmvpFrjHjmq1QXmI
6I5jJRXjPK1SjzJkVJ5vgd/R+gZcU3tlHImGq667oN8TklWRTvf48i/l76sU+wyN
Fq9d/rFg4f/eKDBtUTNaTRoKbg02nkqQJQXlL6G6X7DjZkNvOWI7Kkw2hG2dgXaX
6oCCFVUpWGPJAMK0V04aI8ThFcjMHZEn1NlSVtGIX28Ci6G0Z3a0HqlrD+/03M++
+rOC+x1HGvPbojSywLtE4IW1ShwD7qSnRVFKJ6luPKi4ZI0o5AzHvUabNFq7RYLP
CCEAozdZNhUc+IixFWQ1k2LaL0JAPOxiOG1BgzPYGXUa2CSLZ6u9ANX7jjE48it2
fZme7pfo6/5w4gUP7qjBOW+P/huG6XSu1Q+ZjWZFxuY5n8hjzreqXAoETQbmkwkY
QgjY+bdok4h6wE6G4e1BbgJ891lICH7K4Xsyjj7U/gyzOlKGV+zCP13Dx75c8Jwj
Wv27W/1Y01FOe/dk5ocJ+CNhXVPxESzT6RfrJQ8brQuN9BeRKdFG0cvnDssfEKCO
9ObGXpfZn5MEnlAxpt4McT4zUT79UJqGGRRE10wEiOq4JSSpDOLjGte8c0TJgXtO
2TnjIx5xUcQ4yLEFcvSW+uglWZRj65RYP4T6kR4uKYEqNwlgQBFglPwixAgUFkE3
36M+6SC8X9z3BIavMhkUl4mkiZ5PCemHf9cPq9jcOMhTdy6KjDfGZh3IYD7+qcNW
n4jwuZksESJWxgu2Pp4f3lrUyppqXG2xU9ZvV7yWfKNRe+5mWJyMSUcimmo4sKUp
lLw7ub961iC3ruHDDkS4Qnl3L5YH1Uq7MJaOV49+cPt8hYXYkcaHoXY385YoPc99
l1ib2ZjFbAleMpoYnvr0qOG5eQ//WsPtiphO+h+flkyVi3iNNKP0BstTs9lPtW/2
pLgcwDLpLnLMkQK2qtIKPZvFvS1Han84rf87nL9nQhf6eDur4EgnWyeIB0NFKaIv
6IWANCzA20ToFKD/23DnGV/pXdAtEw0LGomB4k80ojB0ZopobVwE4CD3R2juOEGG
11eEzVQC/zNXe1/vKnfF5Fn1ybUqMeyAGEEzqssZiVn/HaAJ8+r6SZdE/VR0/EeH
KjGkMKhCf4iMtyfeo2sKd5R8xe6ium6y0IY/RPW+CndLHLzXx0Ckeuq2grRElg7V
z0NHigWt2wmI6Rm8F9+g0TSqgqjEQ22mVgnsy63K70XiwDfo1pnOZb7frdSMUk87
tTmqY6LzfY35jw+neDBvyLznAVByBxMpKOc9dG/J0qlxRRBRMioKmy2WgKjam9nt
R4SQupmjrAaLAPUUYR+5SfTG+zEOZS8qlLbooz7PfDEoGHVdFnvZPLKF7gRRsTe0
MpSQnKssJ1LlHv6LhSVSpG/38HfuUkY3rRgd/63Bg96JasHRJptItCgryP+ocMbG
+GwjTCt0J3aoBSIMIH4kMftPdz7pBy63JEAG+i/GfM+Krtlzz2nD16P9vmM3lKyA
u8O+vI7oCYcRgKBY77Su3tq7KwgeTF7xm39/ftrHWphcBe2V9PPNeFkL8UkxScdw
YpP2lYmvreZbAO9/jasNo8lSmfUEMQwH9qp+e2UZoRjQsvR00aoXkLGEerzUBeBr
4qSOMintaR2G5A/3gmkqxI40gy+QtoBbPZqcgPEKtC9WoZ/Izt4ofNf+Gvs/UJks
AKkysFsJT8DuVJV+b8dm9BWJNz5veGYZCLXu54c2Ng2o+5t5OSGlz8cCpubnvST3
wYIn1WxVI91UoeN0VuyEwQOtWtFTXZd589pmudx7Rf+UNLX3IpKtWFUWvuyxlAWO
Hk4w7fzW1shISLOq5snFczHh0IHxN2Rmj3S5nO0sH12kxmY1EbEIodDINXniRviz
MwJycnFpeyAzqh8ARt0YSLa/sOo2IsZRMCaCyKwfXM1C9CGh5+W7uVKp3nXGBQcN
VmJrpLfYKdXx5O1dSA9Mennd0Sc3RiyLnAlEQo5ciSajKneveutDP174Oc5rdxOD
qt+qJU9Tkx36rHm/NKlFSqUtaNvuzmKmbuIXVhlIJMtuyDcZZCp17VEyCtysgVwJ
U6HMEjLdeXvIS3tEO7AWVa9DnhTAWcMzt0thJR8fxRbRlbLFg+aokZ6wLto+udcM
QOQwg/80/lg3Do+JLXh52y5LszPL42IwE3YNKQNOVP3epoWAilfyvu7G15/f55xn
spvQ7EANJobBq7cPaKaNIMklOA+sVj10J15BRQFoLgX+8fUZmmBoObDIYmBhEJ9y
tLyAhYIijmimrifWiYhO8CByKafiJODbDBgQlEPLHOlF3I/chZSTyjrSdSQerUJz
7mB0St+tJOiqVMNP+qWhDVxtovD7IMQcm+qWze96ZiGaMW8vuoVF2Cxcz/JWAixe
SqRk1gelybNHSmFBOpw08ZGyyKgPKnRzVaOyd8BWEApGPDc3pOlkMnmosoSl3vUE
V99E/lb6TpFUDKFVcK9OkLo2ZBqK56sIFIwGH3ldi3OJGu5J8KPXOWoGW1R0Msvv
BmbZbLC/+DRQRmDndSPli/NmVrigOs76Se5cWG98g0FUpvnow+k2XJI1IPYWHkbw
wK3LBNO2LUvq0XqEwjxiqOLPHp6WhUf2LnN57VKv64eAZgdxruqXHMK9xx0Rx+yg
c9JtKb8HOg4t3NVXxJGSuoKPYvPPncXLxXawwmLF9mrgSVCAhZek/SxbkSq8dZhB
yCHIhofUKb1/6w6SAIyPYeVjxIybgM3Hbv1AmPpyzbrOYfLKnHrldIzpBTtucM59
KknKwmm1vQr38DTZgj1w+fSc+4xxyfSNNIQaYfqDRVBaQFIZnBci0WcCvCFvKWf+
K9pPg8y7DVRf/nnshDrDGvUtCT4BIVWcodtqsLE5LxPWiZv3ajQMtHgxkUjiuB01
JaizQOTWupuNJVvSzjDP/jiECRUvsrRLDltib6bXInpfK44C80aRDQBQ9aMBucFK
pjOSYEBqXHrxUYakeWZZajfHImZTRcCFrvi+35eA/1Ucxt2r3KyRvNbjqXA4KJZC
75IYHAHToeFl7zBN8TrMGLSwpXnLJ9+Ru+DTgzhNkOsrw+8skVBuZvs/UrA2uIK0
kf4rMjTF5prYVLkIaYvR3k38zq9ugWp6LJYUxTmFivw5YY23nzbfF/iFMeAyMhhx
QQccipJRyxRzm/6+/IJvoxhJILfa2hZ5CsEIZvHua9T+2QWKPW9YPFxn0cPfcsLb
l+mliYvAEJ0lFtlQSaMt6/yrSU9VBriQiPbO/Js+SzjowvrdE5SNRiF1lY9/GCUX
vTF0/2ABN+KsLEQjUq0zyJKIRUEumONZ3FFrrruclbdellt1dAPp8dljJw36O32s
q8b19JMqz+8AKurfYCnP7CUpGL51zyDFyUsm9mn3wkDgE0Ci2jL05Vz4rxookzzT
9ycsS2xGODguM92aRDdn2yr3Z/IMCHNMs1yazZjmU85lkjMmVIhqseonafIV9HlU
+hMZrhh772V9tFo87Bx3RgcQoCoY6Bs8u4kuGRrb077MLgZ3cu4bRrmVGbSpGg5g
n3n4MQ3U7QL2acn1gtoo0wTAJhqTcABsIakCJy7CGAOoqCHLo6FBUapXNr4jTG/W
Rv4Zu1COrVN8DRYtspX41E+rkKQ2mopX1aoMbVlCx5S773BY4OVR5lqeMC4DgDQw
bQZpqLqBdrcYbggtHmeNewg006ELcr3du9GivdsTSShPW9S03GLkyxT1KlC8cFMI
iXma8JmpVBuWBBPUYPQHmf0sY1O393BUZCe4p9w49FD37idD7O3AMpMpruA79o+H
jfKMZfXd50PlKOTgidp4xE3EEWfYdDbgj1/wMiK+H9egWtpS5RaHPifkt89KNen8
mNkej192iDSznVvlv7wWjVOhTSJaxW/kEZBLpg/SVhm8hTVQRjdzpdzzvDnd+OKd
ZN0w/+ZIafUa+fbaESYMWBSUfgw8mx7Kt+ZfmEjdFf5U4XTeKnnjrTbu1upZAa8m
1qn4L177GNz1dLMW4kTafgrjZulsm/Z/RJpiGkC7PCdA4CAthwFlgrAK46SH9ogh
H3MGLg6jU67QSBNv6EgNvv3r94UkxanKl30/dPZNflvgtnmE4ze9dbGEsjH1Phqz
rCsXh+ePReds07DqzctenaJtjXQMxL2JzkxP1JPb+Wro2hMHFi0SwUNjckjYaHyM
iyHvxW0WMvZHFWutkoRsmN6j19KdOk2rU14qsVDSrYiM/oIvquN/vDE2BrOp2abH
bcBszwcJ74AeGQKGmpdeZvSewe/5MYOifyocWyf4NzhzDVBmqpdqNWeG0mfsuNCT
9JYZnl4dIBxP8J61quYJ95ob0vhXSWr5apdaFwcZKn6v2gR3pjvBv7GsA3FzyfV0
425qv1FQiLwmuQmXjU+oh9C4h7C4nT1RT5RCxICKUYtSj+mTjg/vM/0PEKA2/ft/
Ty8UNEJb9FeJPittg9KM1sXVVJB/dXyfJIzdOa1JTIY5NUjNsloiPu03vPPSQKzR
xQfwJL/qrKCbakeY6SGCt9Us5xIBpMZ9eEDGbfMpdtW/RKqayNYF0STJzRx7E2F6
/1/OjkX3F6IvVOd2l6y/mIJPQqvExy2kv2gNNg9OTVQDa6AxgFM6yVVl8kR2T9Ll
9jF/eAc4se7n3h8FSh62OecMCSBr8h+71yV/Pt+K8S+Jvr3LwCWe0D5oNsH45CRK
3wRU/2inpcUMKup1UX8OxdY2HLCx2JftEzYh4MCLM0UtY/5B0PoRTkaoH37UmT/1
8Clpf5aQadBPBguuIZJxyjAeI+SeHWklKR4Swc+pzDIKuszJyOfj2DqA51rgstO6
TkiG1kQth7FMpj+Yl/uNVE7cAlpcLIkh+j5l9gId9yWJw7P59dhRXOQEBZ0ZqG+g
b0Ik1d6v0KLFJ/Njbf8V3thj6mfleVVVP1eitFT+x6pqXxpE1Q3CAZWO2kQqZVXH
do6/UnR73Uy5OlDAoFJEO/wS6W06fWjATu9v4F/hLWU1GA9/BToosiyWlhrmi2Ci
PWLPU+ggOuXtxifWASeNsMRDe+SS2/M8xT9OC5ix03k+vNrzjUntR2aKjkkxRuGo
2ZPoMcH6p8euWi0Kc163/6yvT4/4lyIvbAWwODDau8K7Se4KBn4c8Z30ilDrYc9Y
FWRnGH4EMzlFxZdtcmLvb8xJM0Qht44YNnWqGZIkBIGgdrC0RDog3n3gyrCYjp/8
fITdNLrL+xvq+SmcADswu4WZas6aDASvysxeKudrO9uvF5IUNFHRaX6MCDE7FeKD
1DKVFxk/bnDSxucrP1uS3MBhtDxfKz9BqG4FgQ3+svj+nGic7SjFIomiDLafCUTu
c65NnoXas/5EsJbGRwVGMVnD4pxXyhXSsayPL0A1NrAQd89xlo4QDjtobRaLvfNM
BShN848X9gQJyz6Vn2sdPQgLabQiAyonZ/qxTp1A1pF2CxnuLSI8FudRpxgdisRG
r0eIxf4b3JznLSPm7mrLzQp2Ly5H4Iyu3hkIzsPiR10VtQ6vLmR4/uZgVH4QRzQe
MOt/wRa2/bw06XC2J2VCpfqmUCaWydGmywFSdhggNJGLqo+FidXTz41lfvWqkls0
MgEKgDgoeI64u/Ml7QGvevUONUY4Rx/CMbj+/QNaWRz7qavr4ft5mGGYQZIhy17n
MRIhe/t28g0u09suPdudB5lrMXes/X4pzfPDMAczvIce18OMh3tpoXGrNeU81Y+4
DuKR4exQzkWSg3vWFdGsuS6xMMrOYaS/pt/doHCCzwBcx/Qvk5JNLsrY3h5DOQVj
NeNRftsrbL37j20FEVUSdwC3lZdoRYwJcvqDTMRfRqaKeCt6wHaDYS37yIId/FJ6
qaTGeADBDelR6RJ6itVLJKrf0qB6u+AkFkx04CTw67eirgk2FcpJBitWQLwkfgmV
sRxVJisqb1OoByTzw6XAbWqu4rKb6Oe/Fz2jFDkucbsfHmCjGh0Pqq1nXz/5AXKd
k/HCJ8sZXP1l/8XU0D8958O4ZbpF4OdffautRs/VsCsIqEjcdnOoRWxkCaSv7rj4
4a1cFLsJIo1sm6ByX2mOPdm8tFNl+ur/i1ZjI0Em+n9l3wsdKAV2bm4pm0BZJjM1
wpeDokaTuUqcFTbUkYspFRTOahiGSdeAZpVhoXgAZAEgEmEeoiKKxAuNFYRlq0YC
Cx79FtiZdMsJCp3HUOgYacfdxqvonMc0FpRgc6EJflKFH+hg8MO8kgJ3+7sCtXlu
4AhW2Lbvcd9sj+0b25lPXwjHz6ANHGnvqUfDe5pUlvqwNn3bG9z6nr2FDDqT5Mwq
AVwaOF6qkV7O++crNahCY1RPIN8Q6R4YzEtmxGOZZMbqtAR5+vX/MQcb5erZ8fzj
bWNmVCgmpP62oCKuNYpv/MDw57Mq5a7ZGzaBDfBgAOwVrPUONV8ttJuRadkK7Sf9
BS2XWW00faP2GhrDHJm+RL9RxLO1OLK9mDMqPejouTO06Z8uoEzFzIBxDUrqDkNK
qjXQwLOVINaDIHdy7Au4f51SkgPbeVKlmnHXiJORQsN4zRPDJAU8jaluUGhxJZvt
HgPUhJ4J14DGah+yx7kEYfTEOPbSVZ7ENEP4AQEECiXm8FpfHA1XUAPv8QjUHHsa
u6Vlo5rZB8JBmCo+HYOafQ5C1JgaYpbcn6+cgayEv4B+C3Eoyj2tYXCL5JtSkhlw
klPH0wt6qeJ4zS/cS1vMlWGh/L34lwup4YlEogNygCdCCCFYjXZ7flq6bt20/84O
v6K+7tjdxL2W8RVDAVZ1Jit2i+M6EkfAlKt7VGdritxJHoksO7pFJSfST8bB4D1M
jAP6Vul85iE4GOSbA7qeHkl/WayVFhFpb3v9A7KlsdLpFdj34kfEx0XLM+VBVryA
Sqg0dOhPqbYq9x7xNRMycZ9/diFtR0/gfIUP5ahuWaN7d5I8pqCtUst/mqSCiDMD
+aNrikDquRbEZLao2Lwb3az0bqD0R3sj9/863lsgXJDpX8l/m7hHhOWn+lT5QjGb
jh/7BsRnuPFGDXz+KTvlhySkUwUmFNjH/8vnkgb5NPmN/sTroFWpzEYzXKYthQ4o
IdWOTRNh6u1ZRUZuuFPKtrKzvDzzrlfDgQOEHaXeHXc9b4EGfFOoHqtWADh4axwD
75sthOQXynYyZsGX9GGU3YLuFbOzIuR/7+n02Y1Ko+PWHKD5TXjbclUPUGzD6p1c
XzrV/C1rU/vNbpeRYrO9sy0f+S3/C4w0GxE9nED6tRjPwbd65Xh/IXCsW06DLS/0
zBQ2sP+QotYWuAPlRhTtkeU9nbkJ314VuYKscyeEIdN5+u+E1+DErwO2G/tbB4YS
qjy8jsoK3KsFXE2xNyRPC7zRGYZu4yaqo9aG7EaqVKwkcu4P1mQ03QPBJc5pbh7Z
aFsRUvqABmIZKkS0eUX8PzyVtAWMffmu5ti9tZdEBxtELBdQWnCR5QzqCVnFDUw7
rVKEucRBZixLkbKJWZSbLwHvOYBqqZhMMnoANAnet+iPxKenDyadoTGi5iTh12/C
o0GR9sza7gT5EH4g+ADzPWYVyVJO0MFJHQC5sYiOpJ4GaIOhd0GscV738+1bzgiX
wurw7v12cG2kMa+WTb5ZZdheKJB5WhpXjKudQd7edJ1ur4dBEzV/JQzh5DayuqJK
r3NwAjdg3FQsqDDfX8gl5XvHpgNn9+TqZODvmHGB0XU0Dgcqd8iXNluBDruR5z+0
RyFopmAzXo3Tm8EmKxt6coAVlk069/ib2AFdlc+HoUHWs9tVDFkf60K9nEyWmKHJ
Vn4eZd78XIk0KAmKY7gEYGbdkBfv32zaIHZjdC1YiaMmfIrCm+6CwWU2t4uPGpQu
xDZ54tH7R77t5RDhYhUNTx6Qghfikjh3m7HLoh9DCY2Ha1RzoFcjx34+0P6pW9Z+
zbbRLhKTs2Fl7GWjTIfDYxdSJslynWcC2WDOxnZlO9Iu44/3zCppeVYYe7rGlaAk
nN6L6BF13j6L0MXlc2lerRaZSz0e8cbbcG7teKUGED6y8saK9LwuOzJ8WhAMGXky
LptUtl9hzW56WZts+OxcybxuWZpBFJRIRwt7HyBEipUt9UbUexMtOR+HxBDJSVtF
PR7OxXgd3lILDq6PtdRBYHyT1JU8Y6qb9K1aUnZmtHn7hpEoqNbOxWgKiHP7edzq
4geol76k+XBwhMcUS/Q8Frl7+Vx3W4Qgr71cOmPkxnhdXIu7upWhB0HCcS3KeW4D
sI97FXtPPdyw9rpyJlCo1HBMpNIXM3Be3NPtjh17MalOVuJsGTYQICqTbAtVERQn
ADI2bVPTDI8ZsMyLo/3iRGOCLB9EhK4VQyAlYE0D2gQhx0LPG0EZl7FSIoA0TKLF
0si1Tf0pQNYTjDVRNFJhS17OPeCNJDLt3TL1S5Zq5uv6T907U+lD+auw5OUCfzcG
3mt91K5sEjM0gCg5WmmRFqdIjVkECDrytN4qXxa/WBGSW1D5dzyzuWvHqFBtvj0A
LfX1jLRo5udjqrwR6Si4f73yeHl96nHEwtK2JImOVC2yywUPIeZO3VVKIum1Pl7o
JGFsLy3ppPF+kMar7N6Ox71CZQgCTistPXl2y7rItFNl4RX59Z9zxtskXkZHiGbr
dMQaWLKY9xscse4u9SSXMZir3jp+BQoM+jfC+ec/Jf5NVPdMg/9xzEkIgs6kXxLu
IyoPzq3FsMyW7sJrgp8t7ICM+aHIwBtfnboc9oDYxqnU+x9Lr4sVKcRTBKD4/JpX
gMx8ftpILSWax6abYTVSxWuDPirBkhSdXjEPzIhXCuS2yMDPqgV/+6fqt0uTu2HY
DCXhIjOhu11zRCwZOW+2nyeybp1ncAN2DvwOZoxZe9FVaPI8ZOQ2Js+G/CMtqwUD
DD+FaD9s9DBS2nf3IvXJq2MSQ9zWtQ01EyowF58kFKt72fiGYMymHz+km+jv7fla
n6NeUwNpNv89KHfC9YkNbvdQ+lAnq9W3sWLhPbjNN8hGMaJ71KrMCQZxeKRZMp+R
rzxm4ee5FuSgHA80PhPs1z8J841MkDjzTNkcUamtrbITA6hEr2THQyWadd/sUNgX
2ZbtUVlhtKvN9HsUZzUHvHGpZnDE+0hwX7YgDwHyY4It+UGcmo5byGA3d0ELD0pj
fHxeUg1XRZav9Kob57d7ifrz+pkFxMUw3Djh8ZdBdblO3LRsdtB7pvOu6f/dPrKd
upFLy9RNrfQKzBDlVv1uoGYNKSxnXdqXuj/cBZyt7Gbae4TZpDgoACE+geJiC8tv
liT//ilT7RvWz/S5UXekFDPnDG8uF2mM3d6Q5lC3mXDDe1x6MeWNM+RZotNV9LnP
iw4Tc7SNSdv3SPPpQWTdOKjlpJX+/B/X9lxapZoZhhhuRfQWNfi/f/4ZIZHOJKnC
cC+QSqbp76ls1iHfm033vdd68z6DaC8a7S/5sLfiDOvLd6x2WFxCvhC0ktUmFArB
1e/CMNnfaaLPAky9EGnwCkoSLMUOtN5It9YMiC97w0JVGA9Aldwj+YxaGvPwb7yZ
RA/PnJprjh/OWZZohsSS4IwyvlvTEO8djcueLMEIx+eZUPQMn/RVJ5MfNoKkhzRq
3/4eoH2FIMHmDaeI7S74JO7/UZw8sfvBf6kh6g2I0s2jeiocdKNKPsz4qAA50SMy
2mKY/hp8KRUohTftcijfYq6QiFU8pTvoEh+QGheshF3/DKLd1fg9E8rrP1cczUAx
mX4bLLUgY8iXSmgBmSXSyfx0BZaTPzd9jWYgZ1luShpMLOPT/5IBuSQ4qRd6wU5p
W49hiDNr3li7t6z5bmhVVHT5YTl0MS2H2jeDHZ398BfABHMAbNhH5k9DzN1zSbKT
j7F12Oa/D/eMR5tKNlZxCyFXCSkQCW4JBXe28NifGFxUqtuTCLAKndBwgA5MnnkN
s8MTN1/FesQK4dJ6nMEsHcHJ5Bp/ItYBC5Q2aLWXpph4VrsnEXNINqVBHCWcLxOu
6AP4OIkQhWbJha+E88YZpfKJoMfjFcObZX9HfJ3XuZMzyKOQ0GKyZmww05tzyntv
zOFFOn//hr+FTw7Y4wY9tJPEiAUDhT8l7DDJczBZOvtypBUxQXlboQ5qkGPCKW2A
C9J6RO3KU6lPe5u+Fzb77mCpebyPh5RWTlQOIFo/AQLUd2s2yM70XqIuW8Uo4tuV
Kr/ezHm+r2i0JuqKfRGEjRSGeW7T4deUb048/LDeDl8BKmjTXUY4w7pMazDuG8vQ
6dqsfyQ4tYFRLhuSrIEH/KQdnFB9aeLmTbRARj2CtB+J7vL2lIMMvEuFm9L0OyE8
QnfkXfT3q6J3y9NXZ7EJCyB0rMFS49ClathTqxAwub80KwOrXPYJt3/nCa1ozajg
jYwnf3eU/cBBoTy6auQmuHGA8fxTSrVKDCJQRuOTfu3OvHajgtNclrZr4KFf283v
/M9uR1dtI8xKI5U3MpZTHCnXCSzlWWyor144NHmZaW5ef1ihtKlbyP8AtGVYRjnh
ZOto413LqDVkbvn4MTfBVAZlxWzEOTBb1al7lc7ixiIdXR/2rJy/wh1eo27c6y2C
YBx6lTIqaSqmfTFndwYdwqc5Wgf+Nqs7KCPCFOofMx0XFA/MRcZsKmd4Ny+VjIxD
t4wSo7n/MU9AzWVDDFvTcV8eSrZnfR6nUvoAHI/3JDO14CTT0ZwQYkdgczGUtm3R
Ng3UD2fyM9ww3ObzTnKAbF08F1p+Ue9imTzU/J4Inc3WdU8bLZ1zWJ8QHlvhpkIi
JVHoxXzbSOb1dzwLVvU8RiPlz5g17Sj8L5BCwKoYJuBMVW4Ef42HzXdr1/U2rkai
CIRo1EODR18bcgm7r5wsGlKjkuMdmtQbJruPsLwAmr2gZTym/pjEdOpmAlxisFcu
ulwT7eqgghLJdCx8K4QDQzDHc8hfw3iSD+c6SDBNX4bzd3f5yc2kPDbZD9Mlmi2Y
2+OvO6qokBAWAhE2LMKcMfNaCm/SIMoAkbu+nMg4T4VXME53PlVsCG27tTkXSTgL
sPiW6qXEhNuhwR7xLqYXFQhRVBeiUR7tQRaiCL9i5a1p3ir0t08cGtsvpOxy6yne
3s2E887xARtcEYU+lszLnfnQbFfZleqG0rJh9/RYpNT1X3bMJ9pq1JQcEbQI5jOZ
Dive8iTpoxuFDaTdiYc+7VWV6HJl60SCAt8VszsxiCYBFRU53WSD5rI33CAmJzVC
iej9BEj/4S597UNbJlJwsyfFieENDjXavSFn3K/vFe0Mu8nst+j7BD4rIiVvUKpR
GUc6RotluU6OOZjt/d87CWnCc3Wdi/ECQvuL5+LQCZlA0iQ7r2PjzfRftb8EDYBJ
slMrjsEkBBAWiFc6ooljSPkmbriIqyEsekhnkI43eyrjKmkk7Tm+oK3I2CpDd1Rn
q8TMiuwjT9H9RKhuK9SfsZOayDclCQv9RN7Dei0ic1AZifNNu3891WEf7Qyy7dqr
w5M6e8VmIxhgybHMjci1keKWvt78upDcNsVmcxKAnRCD9kKciFqw637wbc7KrS+/
naH8AcU9EESYsqGoOUD3l1AIEbqNfHbf9f3SSSjZ/v+srd8t3GglOg5uX4r0biEb
hJYsBivuqmox46tt6OlGvceB+uuO+//C46A8Sg/J8ehU+bKmRPUDSsC4u+ym3LJu
miW0bBZp1kaEy5P8rbgG/djDjuvE0vLsvFdciFlqYHVQhwwyG9HdQNUfQUM+xsUe
ZcxA+uhqaUdD8GxU5pxq36SWPDLIsy+RzIr1PZzcz8hAxfJRCLzf3zAWSld8GCow
7H3/yg2Fur5SntSeafY3gmRYbe8sEqFBcjel5zwGW7tIA7ryHYL8/ixQn9fTaIIo
IklctYNdanSuHKWGVbMBNaWYK8krikiZGJMCe+1uSxdfGK7IvRmZXefKYzFdNoWO
Ay7t3suwWphTta8o+NISJh6TSL3agW7QLdFQ8vXVCmAXtTfrIOrXNjBe2L9pcIRw
H63T5LeHxOi4QSk71R7DG7dkOTer1TZ2e2N+mnkGFEZvR3J9TZWV1p2zkIgYEJ/S
5j0zNEXnAYI3UFMjg2RptgK/rCnKFBwABYZAqks02fHNr01X5fEq37eQKoiy3ON8
dfLxIziXrBOsSbvC5OeeZjExlHc8QorJq6bGNPqt93q51Rc38o/B00c996+DcIlf
nt7n68LQfgYyCt2aZe/gYxIrdWWaF0YPUzxgBLkw3m7hnq+cl8hZSJfdwLz8Rdyr
9Z7/CoTXsIkOGLU1Ift26aUm9xQOhTVJ0olng5Qa/pnQQ2Fvn/rq0fUGgNjOVlH7
39E/HJBybt8/KGm/7UE1xAZVwsYl6ePRrWwQ97NUDbC0rx3Nqb/H81ZOZ4YfRrx9
p1vY3+r/ceDhOpKR1luu02erxzcD22EanXpnB9Lox1hdD7O2rLCK+8kPvgYY9wvm
MSaaNxcq8NQg2YhDrFre3SBhrdK0Gtq1YQZYRkYSG11DcXDjBT+e3I9B3hHy/aYQ
SngWAsuM2Z50VkPoa7MIfquCb9VX0YbPGKDYYS5viKclJu0W3rKphFkPbyHcPrOo
k6STTh5jzbYsJBWf2pMaRx78lrGIBGy389sip0P856wupzNU0zcbPQYWiLGwjKq+
49v+emF9LqsInIItn9IwD3bJ/ZF2xhtmTPxhk+wK+UePw1NQScf9c8ja55AOo+0C
O2wJGLmwZKeCZQNQGaMkBWTyU3xg/C42F+DnVh0CuEsltkszy8ClaJbAzAiqAsTD
fG+ZuXaX61j3/3eTAJmvuAEB6Peguex1lAHqSck0AL75d0JwQs3+X5w6VTofUcwD
YoMcGLEhrjOOcx9BCZGzyZYzrbOMy4JBLSHziJDmIcPdKuiBHsmc9FXuAgV4VPGv
YAaeLhqQGnr7DOmLSCyVI9gs9GSuLQAWfZaLyrRve1/h3nLdVAgXrs/oR605uF+a
3V+L8C/uGoemYAjLoGYV2YZ5eZHw5hzPb62rb8NWnIDX/USfJLH5u1BroGqyuAA/
nPoQ110IRnwtp4rGvQj0KqMmLfxgaPNBXnEqIl2sp7NBsVf9XgvJNmDRiMsRYMhi
87pH+hFFMC4WhjI6G7L8t3mpaOXrMMlDrJUExQU+RLpQIuKsiDpXk0hj3qiw5fLb
Ftpx7o33baqHVXPiXkpY6mVCNWIP/UdoC1THhdZ3Qj2k521J2jZvRlgiHFuJxCCQ
qd+mHKoZ8fuHqJRyUGsKRRZUFwj33Og5XuQvcEYZ0c36G+SSWTXtJYkQLmC52CJV
JEqEmdFwFlAhaJmGT+TrCpEXGjhRlxcMEO1AcZgGCKDwCe+R4bzXrWgN0nykPVNd
oGGSk1EvvYrx/x2g76G6+YX6sh0NxZrgc6CwfBtBdJv0NursmQtUJE3h7wKP3QBK
XUyW64a49+1YEHGqh+ZlV3ddxT97DcMZ+PImo4VuN8/IbWb3+iTLjrl4cJrR1VMh
VexDiWey+6+YYKdbYikq8/F83Ku1L6eYkllQReWVqoeA97sVJHtOz8yLH4SlKDyH
sQSmVqUHGbHYxkpJRsd9MOhV8pBZTjpZYFAsRskoTWkNJe4UnMl1gS1HVMiG8I9h
gb0ORvrAJ6gHaFT8UeWqxNCinlfiGCE+89FFBrgkR5F9wSi7htBlQ41c2drCFAIW
XYWi98Ronxy1cURME4/3jdDMW34htbaX+wOaqI1XOgSChcN5/ZQWCnmKI+pHjD63
OW7k/2x/sIZ35fMxTibH1S+X6/f7HLgRwxmn6+McpR6UbvRmTTy5Lrb2SlHk8e6Q
CjAmz19MSviyqQROkFTOVXm9Rq6PtFHgwK3T19Cm5RrhpSds453g4YJodbHj2Lwt
uZ18J0d4DqDfpFws3cB8ZWs56GqWzmmhmcPoRhBCDqFMId5R14GyPc6VSWlasCJh
nW88vn2kJKz4C40xhiiCk7JW9rQP8nXFIYFUsARGXvmRT9vgziwR2R9itjweipyK
dtw4nkZNdkUvezFSxD++Tp3rd0ZJ3zwykuTboq9EmoU95TNX2oor5roZb7lhFQtJ
+HegjGA8T266y8cL1Vn6B8LvDg2ZuDAASW4uNM1dn5npByryWdbpDyj7wx4iSoGg
OGuk/etvPdxYmBb+ZyWnnL6LZTq/UpNBxAd4aMMvZV78mEX4LKoWz1EWyGciFFu3
ZkHEWBbIaSfCg26hdvejsVC6v9TiVrwedZyTL5bkYwCFAc1665VRzDWlCyf0f9K8
4hr/geYhsy/ReWMJvxBBICdj1IUR4zEWomwxo9tQBxZejfo6lGgO9PCRsK78rS34
wFYb/TWALmI2LNb1GaKWHTGM9MCJ1IQvcomq4etlewpBLquOk1kkgTgpEk3ldY6f
/khZTX3vtFlxf7XFbYvx4gUHyeAQLeJ0o1qPLuNSnBAeCz5pYzAtt3r6zIb3YFFg
F+97ffgqf/25VH5N+iJUGTnmeBmPN9cdqx6HYbbZofJCZc+OuIalvSYBAeR7iHvn
OCrWZVrwPsKqbITTxdJ8Wcoc9kTB+KWEHqA23h4HERCP25DbgQHH3V5+/wat1fjX
MRLP+nDbPXO+Em2wirM5395/IQ081998QaVONTPlQVrH0JVFBvuy0uVCC0+b09am
gXecKv5Hrl16o/Aafyz5ViOVs+YljRkZBaJN3UjrZ75uj26ovsJ4NeMNN+m4KRVt
y5GgrRLteQ83lzwjAEvV2xzr4Vq8Ds/aO0qUHbq/INUQzm2YJFxd2BZAepnTpEzp
oZHv105dzeDgtZwJxDL+8ahJzaxhfEc1Raf1xovmEj1SwBNGwmy/wuxfLIOCmHt7
m91GUhvathEtEGFkOjaK5D7V69tKaLdLybXFwvyhoMjiTeUWOixweREctVdxfav4
aszwmTpWCYoq4JuC3G9+NovYM3t1flgZ8lrEEVL2fHkTNgJK03WUJmmlzYD5QHe7
1j4Gmt/tX8Zt7cQ3Z5TrVD0XdLcoDNBgG5f6Xv2aXiDx/YjRb6rVqXdNwnyP28tC
6U9tGjGlj7ya/yYyZ7yT89Es1tGtbJzQX7NAhWwA8RtZYZI77aM+TB4NjcsnNGRi
IgXjOLEycb71dtzwO9K3rZ2CjT5P6yTFCTVD1sEw+Spouch7vO88d/XzVmKtEAOw
f9HuRWFX9t96dhK9LVZNNwU/i8URPXRsco1+1/6ACxm3xawhCzGDjjD+27b2rNX0
tGTl7YZ9TRnMbX2OZ70ogcPVCAh4b9orNDEvXkZNOyWN1CN9m5Nh+sRyBjFFA4lJ
NuvGFvH/vLHPX6vBRSr/UMNcsiyHGy5ypeknUQeGHyxHvva/IMdRnAoA4HE7R26b
2gaIC6anLf0MF3c6gaos8OzRlqJDDHahT/oHQkXTY/Nb6ybURihRiZ5b2ZtoC+Uo
D+TJuVxKoh/td5CUwYiaR6NmJlJUCuzxCF7eShsPZeKkp/3B2hy1bBbeL38nhAbQ
5Mm9dxauCAP/zGOpz3tqwUnaBMNkv+BvIAxBZ7yYl1GUmZLk/NOueq+HjNlzPc2c
BtH5KUXkltuqe1HxjIozCk2eWM5QHa4Yqb58d04CGsVvT3cOXcuagvP9seX9eQwW
aab1KVlSY6H6E727m1cFk03TJzegsZJynWxl2eSyLPJ5esubWV0zCTEyz/Vemott
F60Bhu9gknBmH653pui6+h0mkwRyQ+gyjVDyTA/2Iox0+0nEdYo/yxD6r1+dhQs9
phK1lp2pvS+u3rr8hmPOXkaWK5pckQ7+sCLqm6MEHANOOrFCeF3+L3sob4IVigRq
0rDueacaPIYHB2dCnzgKy/Tkt+El7esWtZxGIaq3inlejLQQCzkllbsA2WbxGmCl
FyeMhh6gaFxwCW/RSvUKeaJIHNVyL0A8PE+IXqHpeN4I/GJbkF+aiw6ulB1tgUSh
3AJZpU2grWJRUHmuWkTa/Di5xngI/QYA6sSHqxoBg4XBCXquZ6ES4QgOiJtU4MHj
xweMfcAIHmacbWALbUXtkXszWKLisOpY+Yk2eFm/00noEf4NXNzesZjN9iTavklH
QtdQTGuY7puvThuP7Dc0+QvWZHke/1Gp1kPj709FkPZNEkCslCjSh2uYouTwgcqy
I3KQhv5RP6vyjo9IbYyy66aFEgZp+NhWFhDAnB5QEi7jKLv8sKYJofNh6lUu69lD
9tOrMDV9rovuE0Jlr2X08HP4oXuVn6NrZilsDJDauNQN6t9tLC4jPHpWKvEA94zC
Z1ZnRyS0xY/MGjIwvFa3NBJKnHF2TDVxDcV/GWSShPEaLAvUTk2hAnBvFHLnHFSZ
wjYZbkpo4tfqMKPbt82BSK84YgLTb4V/vNOvdIS3rQeF462y2mkUePcTbXQL+E2m
rk148+ffCn124NQ0gcbtOTLF/b0xLmJpIzSkGRyLPQKCBA2iqUBlk+17fp2evUOX
VJeC6MDfZIG6xR7W+0mfK4KLTEH+SAb/HM5ERtwj2wJWAvXhTNOpit3O1vgD5jJy
NabbEJqOgMqKmTz7F+BoCKcAukb4zskTHH+4d6tngHePU5uPnW4D2S2evFDyXrd3
AQBLpsHnWoAI3Whu66a5/ovqchertjd3yRr9oWtdsWW3xW+NwM8EzhbRhnaAGiGc
yzSTj8430eNldS0iQSBSEs1MKSbOQT2A+DGzp8wihe5jgaQwGZgTJkrkwXuf6JCs
reFHdyqtvLuNzE1vRbbGrok8+V/gGHKLoF4UblUWs5U9Xl52YFGoOIvZq44RiTUW
1lcSklc9Xzm1MFmddJgUsXlYvejvuYJbmj2d9RIQqkKsLA4/n5WWg/mFWOC2CunY
dFiygX034wYNtmI8sxQim7j+exSSaYTku+Mhslnzz/3wYqllvcqLm5u7TXYs3asm
/62+o6dREkhSrgYBx/cW8GsNdQ7VSQHXMOtAGc/7HaKSNqtj1wCa3n73st1GyVsc
JbSVlf8+uPTSobWmzt18FcjAuePXKVo3g8C/Sgh+/gh1ttFRm/Vg9JkLVe/e3v+u
2amPeR+O0Tj0pGuYE8uERNzZoz0g6I48HCPnNYhYw68xHVzCds1TWvIaPpko5jJM
EK/pz3t8rwFUtJfzJ8j3lvXvDC+Ohu0gSiz8VrBuku5UObt4xq4TuL0pnYlcYGvO
AvCdU4m4fhn3rU84SfbChPHer+p9qJaZNUKmN/822Fd2IFBpJtdr5qaW5FEqdRdQ
3IeyW0PCrjlF2Aa+0IVKg2WHJpKJNWSDQwTNozWnKixsNNpv8QvgOX0r20BKIOM0
icbKzlhERpZ+EvjH9M950TjHPrNeCaIweGSAY2IiX1YhBEFdeoRZyozO8Y2VGETB
hDdeGH0RYYRrVP0jsrTZLquzp08ZFrBqTzv7mZGwBOz0bZ1cXY8mRIe4PvRC/2aO
krIoVG/l9+sxBFYvFjt2o+9y4ATbBJh/pGVCp/3gUs16iC5Bxq+23jNBQFOL5pL8
jKXrMrD9vUlmdH4C5Wphe5JI7f7HJljq9MV0qPA1RncTFB68Y8wpBzUpTxgkSiGn
w04w/lhoK1Aq6yDvkg+nt1QQ5iKgAH3YlaGLsLxZqlNF+4qVnfKBI7jQZi0KZahZ
pbLxTMwaF8kfE8yZh+bEG/x1bB5vk1GSeM+xLv/AopAFWuZb2zzMeOaXrTIC8zeu
GjpldXmN2bJ678IHtKyA7Ms81sXv6JGCekXN4etGVAcQqyunEOtKbUWhcy7BwR17
7osP6IT1Hf7Clof9EXXFB7VHY0ghmLAoUOnfQOV0T4Uof2GeyAUI1MJMvqfKndeN
IUKMAbRoJB3jxq/KvclVq+S3+UwEiP/ITFTZpCcjICN5daFHxbILmlNTKE8novaQ
x3Civv3+F04RpLZ3loMgDcK/uOsSwH8DiUVsPqJJJ9mNJ6gnxMGCxpMSkdoqOMZI
N9MrSN0YkPeZs70nMWr5r2jluylLch6h6ySGySf3FnIzGqrTVD1KhbuHswlimDi5
wB0/A9r00flOzh5hBUSI25maYJxXJSUG+YJy1hKslKaWzl7GilQKHgXcLdApM+9C
RcmwOP7m1n157PY5d6RTROTg6C2Y7ghnV47ltw4lBw1Oo9erUEoqofIGeq/xaC5e
FitZTtjug/T2bISSwCQVBzybjD8lO64dbYCPM+RI6Tvm/KLr1LZ/H9R3M98xICQd
8mRY56DL73ks0+z09PVpL/qkbJLkB5Rm/FsQK4xFR8VcVTt9i12d80GNkHYet0FU
ZAGgDsgYUc0QunAM860u1zA7weUbdiSWpxsarNXnYRnmqFhDPbPr4wO9xb4HVrHC
dvp+J1ewc3izCgTKypm3Un+UB29E6HaqwFehKtqr7JXTAHvhdL1HE3VYPp6yjh1U
YdQqyOTyiHQXZv3Y6PF+Y1MNYqnVxP2rpD8jDOynW30TKrNwN8TPnx3g8K24dyCz
wsGwH0xHT0e5CM0+Pl6L64jjLT9FrMfUJS1osotA4dbXvf8sJRnR/2EeS470fofE
hlnHaxpY0DzRW/6jVen0z32sZtU4WR1gS4xQGIiQ+6hj0mCk9eIw/9dCAk8CyQxZ
Y8ZQ8mewWyX4G+p5FjYhSy4+SDPh2iz34/My0u6WzPrYHRBj8FqgQNcy5Fqf2YuL
SuO3Gpw4jT11lh8aMqMvMfyOXLHSVSIoAbOfcDeziUB++mGNpA4wW+5bKMaFPV58
CBKTfDYJCVP/i/jJ1hcXul1J0L0MOIjAwIiSqgcVAVUHYnUaFzdZPhEMDaP4M0dW
5Y2XdnP5NNGeBVjKkT7cPaO4W0mw/h6uJOTpzsEcT5cE7y7298bNAeE7eEp8Qllf
Af6mYpI7ztLy4t3Du3pjzJr78LdZLRidxNSwl3nBh8QDhNC6FYMf6v1fSsZvo6Ng
oYaXD3OmawkiHC3x0ccLDlUaopYR2nqJ8HqkgJ88Ym0yDCPl34foCK5zR4JDAWo2
jaD6NAzn3/mYnsac2nfixJFGcNJ6baVyd5GlULyJqxVOk+7Pf6OesGiKtKedizSm
J2UIs1VefET3+WQ1CdS2UPM1KFr5y2Yr4uMtxc9rZHHElD1y9Tmnr7BuIgCqh7YE
T6/TZvsqpREERm3XlFmt+crNNzRKCsImkiEjxDqxjiCwK9ogIvanOGj5KthF2WTt
mf2oHoM71cp8r9q/yzbvfch7TidTHzvsGwmSSF0RTPl7JtdJ8FuGMByU1jmHrMp0
e7AIJ/kQbPN+s6TasxDaDtplhh73YANpA3U5ODj9PB/cJcZ/yz8h54UakMWXZ2o5
bb3k4HoLVWwfG6Vg8pa2vLyoU9XLzGk85d+Kg4TSuRJ78yFc10q/xxZqeX/UFOPB
QA+4aARyKGYnqRGTmlNPS0Fs+VVT2la79oAwFUmtdMcJLbruryTCzrl09rWwGYcX
PKcESU7UhIJUoH22X1KVw23mXL0ukyN1ZKUqfSqIIGwtEXlS09cRhfvIDZjv58Jt
x3y5ww8k3LxMYDiS7En1v3m5JJXFxwiQ/hECWJ0DT585LpAgsytLHGTVby4dKy7D
RAULjq/NN5mbubV7+Os+j/DKouZxL2b1Mij03FgytAKGFSYqPRnPdxfiDLsoStyb
hvnGoZKba69Yqybx2zXUxCK2KqwIfOphV2oCO6E+tfC5rXEuBKP8zEMtm3NWVX6t
6VRK2Jy8MJ3q1fGxKdszQ0/bD5jne+YkvxDKBQymeeNRlMVICIW+V4SKbQLlVrrt
kbkebx350LsE+l0gF/gBFC5eBOOr7IO6r08tR6Ys0jFB8ZQwM9eMoqYqN67eBg+b
RktFLil11ixZ5Azpq1vaSE63w85mRwoqu90vI+cuGMVVrTmX7f9fLqfCsEYI9DbS
jVA8pMYQRoLQUeId29W2KQ6Y8VaZua4u3dJYksXM00kJPGnztajLSGyT64G8EC50
KjGWYqC5yd3NIZv2Kg6x9/+9gt6FedCbWk66Mp0uEJ/+aQ7MQbc6E3UX+b7cU1Q0
4uLRRy/9cCrhwp+BLMhgIF0R8XGBe2alzVcv27ccXCxwEq1gzy3Ndhi5c2bhzIn8
g96ccSoQUw1ghD6i1YTsHi2Jnmh+cEG5q4Ytol1ex7Wz7Axdglq8sysu0NgnAxoF
L/k/RYO01Zq/mU+WFDZ/Gy66D9CykiC1Q5EzsXQPaxDd6W6JJyRy8bBaqHijfNVa
aiW3OclET9QSb+qrizJYENYNBHsJYEKKvQXenKg/fVyh1OMNBeiaqK/7yH0bgE87
4L1EuA/A6KrM5ceU34w4ORcgARWGZ9tWbpmX+YQyK0MeEBjAY9vkw3p3V3z1Muqg
vJ4fK2V5nGNkt1ODNHy6Ps6Bs9Z9aF7ewVMG8/V9s1zH6AC4Cw1qgfbzmEcJfPlg
gfKyshoGezLicefp7AWHW8Mkj1oDbkjVexy3JNZs8/yDiP7OHTb1kV++uL7WBm4r
ERQWDLWnfL35i64AsU/FXiUL5cHnqo897SAKR4Ri3BHCkwG16R0FpajAEhMTJ8C2
HNlOyRQJzRxlkJtV3BOB45iIcsFuoLFZrAWnIYhdibeN5aB5sCbm2pXU1PLjnDPP
e7RNWTon+okZPZmmHuOTnnC0BOPtjtpJBmCcNSq9wmCdIREAXdcjQcak795nF9f3
0hifgYylS5l4AYG0nFleTIEEPlFNmHUUGQ1ykAAY05WqaAVP9lUgDNUAlqrs5o9b
Yj9qE64FuHznH87VGTgnAfm++1M+pgd/4owdizN+mglVLrLqisQ3t57UDp72KTJR
OCOBsLU4+0iEB/y9nHnzb+8PMDhSYDRep8MRJFoZdPe+WrzTnPCdsvDkINfCs/MH
iPDtOXTbqZ2kmjYw2P1YvfcZjDjEI7Jt07DicDTQN/PbHC3bCm63QUIdZqFodcI0
SgI1a7F2SOQ0qFI1WhMoIhEz8Aixi3lrnF6WSEoOmqDCND/pPy3+8rPbQ8/CUHeO
kkHBN5dAkhmxryZmHT8CcUww8/k7+gyF5B6f5ce8VwWcJJkTVkL8EkzbZr7h8NDc
phpGGVw2t/QQLbG73HW84HaAywyIWUSlZ8kIXP9IllHCGTUHd+29intWTvTt8bKL
r5/+wjCoQpL1l+miKBwqazrxjPuxQ7eR1MJCeDrI9mwklmaA2AnL5CCLithQMbUR
Y+p7W1CM/X0G1CA4NW0pO73/4U+1CWJLzVbj3UqL79f6XXL9vuAup9oaIVI39UjZ
UF78ieYYJRkXAoU/ARaKkmLA871DWhHJPtm9TetMiP1EmEjckvi9bK3bdzseek5Y
F+oOCPKhjYWuyGlGeVQUw1LQ38sTr2aCXePT5/j+RcCKXvwcB2/hCC1t3ipDP/Hb
kURSjUy0H2TnVRtPhSknpUUx/WJTgjCFW5VzEgI8G1ZzuwdxA1AWX8TBtcg/dazc
NA7ToYdPoCZUASAtAhoUuH6QfVkW8I9vB5+cw2q3irV1AVNIBdi/m/0Pi81eo0Vc
1rytuyYZGeq+uKrUjnhtj4a1HS93CSOd5N/eT4yvEjDn4hoHWKKJgmwV82yiXEQJ
lyZ2u/1434yIrj7QJ4ROlqRX8legL+QoSfG27FJxAHOByC1rHzyB3RQPJtuukOx1
TPVKFJhgpOxn5STVAzNT2zZ/ytxbkN+d5uvlxbmB3hdZYWSxxTgqHC+eNAR+Fxyc
UcMxYQw/L7yNIwtDdSJWMCNvwV4TJBQsQf6MfAoOhCFSDmTgP814qItefyqgvmlC
o4XkcqTYp1bVwiycTtNKqKGVDXKlrhzi6LzMdEZkcQJGTC98TdUlSXyo4b6n8r7N
c7Sh9rfvuEs05S+r0lgmks8+FN+l/voGT9ml0DNyufWCWexwrrERJDUZjsL4xIai
zWznbvjXe/7Vyqm6ezwsTooD8bIy0yUYPs5+x1cSrXxMlQY8aQeJ5GtmQOFS9ff1
dxTmDUXAIduP9V7CAzJZijCgPixDRTxP9wKrRsrEduQyRh79g2lNDMMVUgk6b9ry
qIv+ybI/4eP3h5jcgFzj3ElX2lEoDidlE4S92UAfZSRp4bX4ykMJ3uWIwxYsT8Ru
lz5IZ9VDkzbM6RGPudUCfcQJnt9TPVRhAaHo7ir7OXcdYkBqSEX9wDbBE0Atl+N5
p215TgQR4Kmue++63MUyyZPZEHk0L456wOWx0hOHjrsA9KTxBq/mGDu8ck5JFfuF
1cml1spMFVk1OtmFEI56ug8VrYfuF6g8YwfjFfuNAC6NGIAmSIEernun/3ndTrvr
av1PYO6qlsemervfc2nHDkGOmfbAFmde1BFmf8TDJUpY/tz0uAur0VvD6zWjM6lZ
8pcy3n4njTgGPx9AGZGIaQhL3CReR7Eonp1D/omXvEb/ijAOHpXmGzxcCZaS1TYK
EPFzh8TJxlpI/Bj1V2OoO1KG8edRn41dV+GTeZQL7sl3rVz0xCaCLf4LLObrKEX/
i2waJdrch1AurXKctcORU8L1JYSecauxSUrXU2nfmbNnbY+e5/d4V5GxXiOX45zs
K3N0hp0L3vUNLjEtwHHFEyNmzFG2DqqLeGNrCSUlNGUq2gec+1B4Y9OgOJwCoWKq
m/RI8Htdjul0/kPIWmE6IdiZsPUYbFS5oW7x5t657lkHmkT3I0ELX1TGr/JLec+F
x3kxHedc0pt97e/mB0MSE8ccxNk7BXGgy733sq4+F/RTL68Ik9AoDnODBgfLd5Tp
uN5q+9K//GTH3zrwmaY+0IPrzrIBiXGXdl+rHPA5Atyc652gxS8c2yyhV1LJX8Ts
oJaiy2WEt9HpnITPG1YJkEaAYoViPhkbFS0JuEA603LN09A+HYhTP3KBJCwh605F
iuzAP13dBvwmhrsCJnUjge2ErI8eLQVuti+nulqNAcEvgZAg/XtCqL8O7Z3ymu8p
kDyEssBwG29eRYV28ZTodM9XdY7D8U3wc1mesWj2X0bGGpBdDLuo65+/+oWSuiwC
0z5KiLN8PUUkce3JmKGFQl2penUkn6G3bjW8aa+A/HsimMhIaazWKpBdcaXdmKj7
oJGnY4kjD//5QYdiZfy35FH18kZ/A9iTvipuJO6l/JZTU2Sg5jDFoypQLEBRf0RL
df3mA+9hg3RGpGCuLFGcTotxIxOzefT40pZ1q7z6Arxkd97/5YrGHCGt8ye38QUF
FfFv1zFNMLkaMxwavScNbbNiBdZi0oR48gkIDEJ0o8dRhwNZXfxR7W70DOVUWeI3
w4fJieijRKFN37D7VVDWrEQ99wNSyOjt9f1y1I2dmEE9uEH/cVxiqyUWdW66gmbI
x1gq/woLjVLgTTVWBMFqBn2mcRpDydgKov/fbiu1FpoO1eT+SY+yksPY0F0bmpw8
H6uRhCW/l4f7JpyEyD8M7m5pslRs7R0SYttk5mvT0q+KS0MKg4bd7lCk+tDAdkFF
EVuf62Vu7/Pz56uEMG8cDZ5HllZtgo66b7ll2q/lvbGxEH/ZAqobwqqkkObcl2Hg
AhYtwCJxHntGoPsx+ucIbBabj6rpG+guBtJBBoAfhVAYdAM9qq2KNXhBwPeEY1EY
Q68npXNNG21xe4NtKty1IjDjW5Rj5CKmzwB7SkhPTO2GA3Yu5fQd5Jmz2U4cGkSA
ivficms6rmt8p2itxN4OWjPWvCPTXOI2di0c+j+jZf99aJQ/HwOWg9MFO2l3/VFb
RguApGwlGu2GOtwlPkEYmzm5yiSbmPLKVs4O2qh5iOXTl1tEgWwEp4GGLCHvC/BQ
IDQHvBsg1/xUMk1DYpqIKhPCR7NjqCBQzm8utY7aQTKaCvzpsd28bcmOYBhfI3YH
rIvp9H1o7id5jQ6YEo67M9Is5wrh8JEHgYIVdj/DqI5cHUfC307x7hkI2pW7FV/j
XZCOOYilXLAc/7qJv5effywB/KQiq7II6VEZ1Mtxxz4yD8IPXv6dJki6JcpbWUd6
otVd10O4scXK3rGfI56pp7wuazpFYs9KSNBy7RhYcTLlDja320eYAibhdxFh3pSF
3gH/WqgmdyYyu1t+nhtXGHposHz5FzRd838Gd6OQOfWf6HA1iCbeY+hdeUTSKgqu
fZDauT8IwQaUk5Gt3m5J6PwVSVC2+zLjxVqfjZeZkMZhrLXjsK2hDpmlPbMMxNFQ
gF+J4MP3+PmVos58zGoOtEyA6+FhKxo6hmMPyJcugAl0hdRDMcoBEQGM8lvza1qL
ZvNiQFHbU16t2IMKegeq/4ZvFDhC2jqWFoNVcgySQ/ty4goG0j9gSplv8auA6UcY
lY8ijyrX7O7fiujpF/HBgXK6KX6NytO1sw8TlxTqXHDJvm1St450xswhx8/JZKbG
jihavirijCfmt8Y3L0Vzt98NPrFWIE6mHvM95vXecw3hLBnoRI0d/vZPWmYD3+r0
wSgbK6YOF7Aznij90OwFxkLRW3GOxOmserLnZxnt4HeGUIAiDNOjdHWhhs4ykrbh
61FLC5xVVNnoPBF8ibUNK5PXwpBejos1dIMP3EyNtHwTTcPyrbD01eID8ERY+T/2
pPXNyGOYZhbEW7UynXIJMYLP38M/Z7o9QBfPbK35FwWZVgEdvhrtHxoSye30mXxH
KPO8JIeFBgRKp6sD4c7Br6eavKSYJwr2bYQM3JaGSKVUOeDE+GcI6PB9Q9WyCtTy
ILrMRUnNLW5JXkYl6xIVtougI11gvlivyZ498ZPPm2ga5Gd7+Jkyza5ggIlSir/s
vce+MqcMTHbwbi9DgDiaWfcQqdo+3+ZRmSXqNfhQrnmILyhIIdli7oEqvKO8zknd
LmvJpTRv0XAkcUSC5vj/QTN62D2cJSFeNoOiuMJZbr7TXg+wu3AQT6K/Y+Q6CenS
IE4bc3J9b9aslceJnN/g7xvTQQFSaojWqOkFeYqbMKGxj+7F+5FaH70vWSrSjwuX
WV/DSS8WuZI7ySRhb/KOInKZCr/oaMWEUncOkrwhQ2En86mYAVdprsGjdBX6EklI
8fyHqPozVhNGo523Kp4QrWpcR/P1pcAEUlkulDThRE9YY9yrguy9GRR/vcdr7gdQ
0a4xVohdkcAbpMjw8evIDnvZTmZ+kY3dTj4GB50jQFVVIS9fCGGOuV0SB3jXqgf9
abr+0dQ5bIVmIlhfVyRVFrltCySjD61LrmqcVxC9JjX6RPkLSGKk66JBMC1kf/X8
wS0O6YZ5iB20OQr1CzgaJrIfc/6nyujER1xLhc6TE8OLgfKExmzC7oo2opln9wCq
M4/w09tNVhcVyf7Ltcz6fdEflwNRi+S4QkQp2lIa9X7Y9cXULvMJqJ0WL7SsrDEK
IhA1Cc2RaB4zZwtQzIqqX+Au8LKvNKrULNSkU/7X+ckXePt/jGxi6LB5RMsRb39W
aRtIfwDMQB/K6vYEzZ4PAzZQ8AkHoHYGo7jzg1FhSyyyNE7dO9qxt67iGgjGv+oj
DUe6e72Y9ivSsj2VZaN1GmZQiRzk8VsSV63SUZWh4YrWLAdz8DFWdHZVWuFo6tsa
1r/2wr8l6KUG2teKAfmIuFNqGyBDn5Xj+LhiSPrLElQyGNClXLl1+YIAwrcD6i4v
f4GX3XhvvOIzwATDu0hDS/FMvEcGz460H99emdj0VITdw55vyckB3OEDxLEjzFap
fuiZhAx7fJHY1X28ElkqOG7fZeiHdZdyMqdvget7sK8B7dbJBdAD2UrCHDXdT92/
IlfVmqe3h/zktI3adIz813CGz8w4lJLTqz5RCMfI3rCNfSLUVBRBpqOhUFAv4lV9
4bdFek9izpDSvtCSYUVZ93Z+FhLuunNqP7y5/vdI/iCqc8OXyZ3ic6a3NO+EzjjG
x5+e8uXFGWvns3hNG0tgm65RHJJoNsUuBjg6J9KHL2SNpjqeQoH8OUOZ3UzhQxwC
oYqFCQ6wWj2hVedTSm1L2kAVH0T/hhOy4E+bsOP+9FJcn5RD+kc/c4Vbm5LzhSNL
jyfN1FWWXxk/g7svv77JK7gJA7Z50lL4iPkv3TiT6VCwuxKyFG8Waleg/99OJPT3
K9pW3aclQfCZkarj92ixPocrYLz7jQiC3g3olyJ6FzAcscEEehN7LlOGWn7EiGHt
uS1d7sL6wOJk9c3JL61320Umekuz93a/cbcz5dkKsi8ce8DjuKff5gDiL7pL8v5y
ZaL/39lqQwC6JOughMwVXTofPhp+XTv2n8lCY7pPu5YUV2qMRoLbuI6bJhXDQSCc
t10xaGrEiCB9cXpfzMSbopzLPAuOtmqkip21XwoJYn1UnuGzO1Ijyepn1MwIO5ZO
yeE453An9NIjD3UJ6JXGD/MDTUx6bPLJX/zwCJ5jm5P4ZlWdy5OS9xZApNTPOuD4
dapb+dobnTBytfaG8KHobE4IQgZ3rvVLWh3kYhJVL4AmmZIDSuplJRMdiHCDXF+m
LFDZG7i4ens6tWprTuN49C5ZpPcLOgRALX1uHP5gmUzN09ub4iy4o1yEixITVARZ
zmRR1Kqk1D96eIFmZVhlzwOd5beOR0gW5nykTifvsnG4IupUwd6aZxf/keJ9sxLC
dw0LCCCmiWSbNX5X/d2cJPV71L8ZVorvwSKHB4D7CEh++Ut5IgmqRonTuBq27NFA
u0Lg+bvAqWMI2hfzxdPk6Izpz0PXDI+pkl56GZ6BQPIKSgXy8u37yilriZJIyWmd
Ur+DZzIA/bDQuZkSBoYe3y/646fCXp2pgha7orKssf7Tuh4ipjCwUMBM6V/X99pt
qFqfh4ztcta2Neufvjo84xVaUUINualMul+T0gAo/lu61sOSnsLPJVfa1c7+6fgs
AJqE/W6XM9DeET5wjvri4RcIqMuJoAihEDvK8dvByJSFcP8H7JD+sK1mhYRmbrtX
vLm2IKssW1aBQHO97dmE9eWuHfQDtN9s8SoQ9j7ueuTMlD+2pD3nnysi+GAT6yB6
GdnBL81fXHb5n+N7LKNuItLCSWHO9o3xdy6yP2hbtFRQzIpQDbQ2RQ6yTmqh7RO6
yJ/N+T021rHJuYhdv3eGWCGLkuKHvQu0fccKhdeT7z7V7Edse/yi1LZDaZquoG+U
qKQpOvu+CwF6so4O7xPDmQWDINfT+o0wbgRrCcqLU4DfMDeZamAKezQfw+3ISfTF
AnaD9NU/czhyW0m/1zTn1X6CheORlDST9dVmPFETNdbIBDVH3B/PQ8Vql17qlSpQ
WDL7VBfxAhr4P6lA2OSq2lbBqpMt7uHxHvFpMKW8o00XrB1ypYi3UERQq0t7ax3+
oVsPVT0MyHqWT1ZkBqQXVrgWOzFf1LswVSoBDbWz7IaKMLh6tcWguuANlsRICcdj
1Mduwxu5mZQUXxH44AXwsjHBmNXqU3a77EyKBHmCq7IyYaJw97uMgOaCXz63SeLs
PM5BiHvfO9iPHQ0GVg3pkfUrAY9MxxgAbhmkpZhO84L6ptK3Mz4eBVNr9MOgutwr
Qr1e0lyxn4rL+Wn37+TpBaRZk4AraXtpGtSZKxRbj0Y0XCf21VakOyRlFpQsBZRy
FTVLM9NN/96tVkG+k9OX8C2ienyT6ildaVZJc9iN7Fbt/YlJNAWFP78eXGS5PviJ
Mi01r/X5B4U5qK/GIeZCCjA1WvuxtSjyYomGYXnH/ema+Yyu+NwAVOpuyjLyqtNq
KsG3B356RogK1/Gduqt+IlqBGUj+1OUGFez8wef64iotcn5bql6XiSwU2fdPFS+4
lRca+u4lY+crHlVaX1/cGLLswjKTa0lo3RdxtPVOpjVFZKoNWuuhYBJyJPKmezgA
IPf0uth8+1vFJh0CuCSOM128o9WuqXaWWbKMOpEaC2JHcPSmQnoVqUxFEPYj+p5q
DiWjsEW9JFKE2++5BakdMI7UqvrqJelZ/NG6e78rcJoVMR3SmZZno8aAbFn4cjUV
DwCI0X8pVEc74sjcA5lhnR0hJ0zEqPPuJ2ZC8IcVlW9bnKIMKWhqNgNlnUzJR2+O
dg17TlVLWFfpySPGI8HRyMqnozJL2XAqc4NdV/6mrYf0tjGpHlkiBfapRn34XnLA
KAFdM4TD+cqVrMjEQZ9w5j+Mi39Esvk9cyAPOqXC38ddKP8C51G8pebZn4M6wW9t
aPlqaHdUpw8GQY8YygryGJ2YtAKL56pv/KoDOdS8Dy+8pPpYNGlb6ns6v7umMX2p
fxGOcvTHtTkZfougPZMBm6DfcENaQWmAhIcKIE4XZonG9+bPRiVSneE/skSv5zR+
gD2gVm10r4VWRWfVHFohiVQa8HoGETe5BugyDkxo/0unaFI+wuOFP2QWekCQqz9v
TnT7T3PR3QbHt4v9yVLrQKXCyJfTAYu0BwDxkW3KLfuL8cLwv+spOTwls/L2Zd45
UmsV4oPpLrhRgCIu9uq7TAsXcK5YLyFHe2Gy/22bsmht5DW5WSfSX8eHFtGaRBH0
3kNjWUzGhFjHnJkXX7m4We469jlGpVR8ykPC9uF5C3FIVtStf7ELwdryiYOu+tDT
9I0I0CUUsyMqlvcOVMbCUqDvuYljaKrtddCSaF/KTFAoNxwet7ZgJMgeNFx7iOKQ
D6Hmm5DCwtiF0o9xuzfq3H93y7zKlYgtgq83fDk2WLnCXnuCmPpU7BBNL/1d14rg
Prfp4tpg/o2ZfFJrADFfXFnz+Ti33+TOlW7O0XZ/ObFPLgSI8FHoAETDJ9wbLO0m
LzvybgHqngIhWEWD/oOk5SaPSdw25oj54zg+zND0bdHLRzz3gF2s6lgYvczoP3jP
FQOg+kJWFe/S1oJFUUNPNJwiO9D3x2V55AqE+xZqGTc6FRR+yg3eahm0zVfuTyOl
3Q1GjHBRkRdtwfXTUEPsVhmqQ1mV3g8SONBgyB+5ma8ZfNkCyCotTJnTdP4HwRIn
okXaxg128WkeF5hgtcGAI+rhhEVcaqr++4/ZCs5uQ4gcj3y0ITWaK/V4hysT/7G2
AEEhPWaCCa42LKamLd7HPHVbbBLf38en9LN0bg5QRcQR+aLfqpzNj7a3YsmtuPkW
scrgdWGVxm18pFimEtWdrYDo7g8L+MhZM3UPR8L1LiTgpUFdpSCukd4ktCccJ5Jl
nPAiXAw5nSVwYCrnGfCK9pgeOvMT8pOLW982LZ1dmiu1Rw+9jUtxj86pY0CBxq5S
em+l50YySYgf3l1DO4iNd66IWL9hXsyxwncPVF/G4EL66bHcK5TeN71o23EvRBvY
nuv8Eb7I7Tv/zDnCIdZaz17MOZTXUmsP4/Qia0hufy6iDFl51+F/BJe4ft7Zzcuu
W19Go9OPI62KZCrddDmi2qZkK0K/MIu2YSben9Z7CHdIqpGmaPM2jVpdQQyjJgB4
HP/X+GEMtXP65xLAVjT50H5IH7edGaQjuw9uGMJ7F0zFqU6B1W58jQ2o/vjb7eOH
PbLUnzj4AA+cqfwVqSIr23GlKsDZUJZKvOkVvjuFOCIM1ozUF4Es9ERNcKUC/S9j
1tqnbEuiHi7VXnCT57foFIIUTEtiy5KG861/Nge9onilaEMLus4opTehTiLc/UeY
3KvqfwaJoFaselGYQFEH+k6Kpq5hYd0Q+vP7hox4v5uV5WHfjsJ6f9Aj4ZQGvLSR
QfwRdofwjxt74STPXguVFh332e2MHg4caJ//abNecPB684PVqs7PEy5JrNqGsRxR
A38GoK3bvWc0A6fU56XD7bD2Pw4zikvT6ljJypRzb3Hfi46bMG/dO8Sj4FcdR8xQ
TmC08/4GCHC6nRLva5r071T5wW6BHlfSgDsQ7MoPDUUTxgkAH1DBmneCr06HmpEU
epPnk6QyVhcEVwpwJbhyej3T2Y84w1xDi5ML+GQInCvC56vG2yN4Gue2dc0xGtF7
9xrM0mir32QFM/ut/Ur35dc7HUbkey1oNbIgJXnixBoDEwAoHugR+jm66pHtLy7l
gv62LQBS86MrHpxxRbJsK5FDz0vfmC3jTV7UybnlUHj4YeWfpgWXoQYWs0gMIh65
0OWyOeVamG5sTwGnM3yvrYHieJn8qIKEqfX/22MS8+a8NLGHZJqRQwykPrKQoDWG
kpIO+bmU9W1bGILy17CYGuGPeVgnnQchx+ERRbkSZBhw3kfsesd78iAgvOMBY54b
Nj8JwQR+oZs51qmecUwNOXqK8wpsN+BA3eqBkSUW3zq9JCgj4fFiMcoOivQ1s/eZ
mpd0xJl1r/wLI3Nm37baGMiiPeKOz2Bp7GJ2lhic4TxnZJvo47PF+DCFQaMixXpu
ty+MwLumufBDW09B4wqlsBR+MEi6ZQjUSBLOCKb0wc45Dy5QdlKAkaLVHXeqbyDK
0Q5obGvhaRWKs8bdE44VvoNATXk5uI2dbT8NDJwHNuizGkIGBC7i3j1LsoO8aO4q
VigTSl8Eo2u7NVHsZP/RVEPpAtAnh3x1GR3k+GR4Yx1wTSxChh7rtFKRqoIQAD2z
34U22e9OEiRcZmQE2bm7HXmbCZ/ZyBJhSekfOpO1hUbGHTuOUhQ9mi2LAB4VOPzq
DtylSRYVJMmBk7jhqfw0OqSquLEp+8YABpXDWl8fijRCGA34eqq6tj2ivsENflQJ
Hbz/ouc54g+LMCd8Vct9lfCjt0te78yOiGRUoFO+kytW2Oc7P1kdK66mKTr62pOS
oXYXxnmg0tHt7NBHAQs5Tw+XJnsEDMjuuPw0BQ8Tmb6j5muHshd7PgkgAtQZmmhQ
Gs9eKzu9cO9ERik3Svw+82TZkgZBtd+GPZTNDioG0ixtqg4nE/JNNO7OO5uxDVbu
Sa0VwBdihK8lfiHSVEpDtGPjVMr3Va9yueIql7qnMZAYurLHWh1XBq1oHHmho/We
M1r0Sx8cFZuX2siBd4jm1UOF0oyPFCKF+R1alvqLWSImdodplO0v/qLnCdszR23M
ADvjtoaj1loRzHIEI97XiCvrLCrpiDThQtv+3GBieDbUav9mPY5zwikA4GMPOe5v
FR3WLDgspMlxaGxmwXSfv6FHRbP3WS03mmj8Ru0vmQDnFogbTHt6gumlP4Z2lIcy
bEkgGiio3p9YtAgnKTYxenvDMEUBpJ3tMq5BtELyKGEJReLhLFOcC306Ppim6GQG
jcfpAdf15IvhjQZfdXwYCbrbvuF617KublQucEafT1WnLxr9P5Xpf4qB+NEKmQLE
SYABOBkw7Ty81zEuX8vsFbA/djbOJqCHkEcpvcn+YwYO8Va1OYKEYkN39Xs1C+qu
a6zduHeJzjnQ0GJ3+deZ03Gprqoon1R152b7HTk8deV7Iyg1KYk2LHqQplIfK6KT
kDNmxFP7aso/R7LBKObWMZVsJI9myh+Z3lF9GkgCMQMRm0lILh/2wxhYRFwT4/vE
MzE93wMj5KHuOmbfXhk2XrYFlGOqz7GTfpF6si32UnAC71SvfaIsymHnSUQPxwUJ
bL1sgNMGSldNZWM9kiAhxO+Hx9nAvXEd+WzteS46m51cJOU1PtErxij0l9ND6xf+
w9zLTFxHk3FiyFnVWCEBI8DlijZU1zF1R9Zj5n+KNidsvsVmCoXUVZ+h5uzJk8xR
hlKBteN2B+MOAlunysTovEiqqn1pV+RrAPBBDaF2vunAFojRuDAYh9sx7K52EkRo
4yb56UhqPOf0fWdN6p3Ucf+KTnbgLTgfUKDz/aqAYPkETPiuPEDOoSmUuw/WcEOy
ez4OBBiexHuKVyxhxT7lG94+JrMXendbeRT3q+Jr1SdHIqIlyOZLdWnID+IKD+2Y
8QdVQysoRXDLFfAg0jkqvsavDkgIAp2J8f40YAGo3uvtFMG6BhvUIwb7Gsop6Fka
6kd8cRPCVS6Aw2h0mVbr1TUBL0pDbMMLXbo3CFRl+wZ1dw3W2wGQcSSKkb8+b+Qm
CfueKJreqvAQaJiJ+oyWOaxrd/1gOXijJ/zkt5xfK5FAB67K5rasxmmAlS97/pbJ
CxYnzTy7n32l4Bh2iTSxkVmSqC87ZamKfjJuynwi4L6VDBOggd+EhzuXl/tuPR10
Pal6OjMwJWAdipnvuyusBAJYLqWFaY/z0NAmz/+CEkr3Ls9Vzvbkq9TLQ/GG3gHl
IcVS/1Wc/3zDxBt6TAxjFqh5mwuCoeCVPH0YDDSyU/n3Ua5AElstkDQwr7Ba2GWH
hBpmm1lzohv6MtkNIAJJ6k34uxSPd8blam+M8U2ikKFVoZhoEtncqvj6BIubD3+8
HjVjoCnVEV0aUMIWZ9kuSpef37F4JdHY/G2Ns/Zp4C7D4M44bUXwOiB8B10XfQ9N
aMHiZerH+WUM80Bp1sYMChvlH04f63cUV8ju7gxmHNT597Z50eGUDNL6KOFVQ07R
+7+t0k4ZSJ/BvgFeTtDXyxAFxTRWo/MBcMrrdm/tzjrq3K+F5CzC0LEFYK1HiLGU
G8ENlRguXSQ5atWNWaurGWCd60/qdsYQyIM7DTsxWauxLIS3VBkrxWXANSiUHaNR
1qiR+o0mTWeIsgR/bJre4Q38Hr3Los1Tpd8/0hqr+NJlQQdm8+mpulQ26QcNK18o
4pbhtboRD+39kzAcrOjCWMLMD6AWNNbvdmjMQeKPfJCN6mNGEnh8G/U1rGzp7NI0
DnymtYij9v4pGf3XuBck9Zpq9nKg2xWj4X63Z8mBpqMQJS9VFiZpoy1WNtgAvnvU
HKw3ywaVOQi6RuqFQCXfxfcbQM6iSgufIHYebvBag48cVLaGOqVrZRgUpRLoehLL
/gzFAPx6QNVe4bNWsQPvLrtlZygKKGt50daAWK1vQO9ivMW1DB8tGc2zLITY7zzn
yWaJ6XEHmf3u+8hGDTTL9u1nvQzMD1pkGG060EmBfxxwhnYesFkaswwpvrMwRm9t
jSdePt5RZSBHzTvvYVG43eLgx5JSnYRb9j/to/rYocesRGSbI623k3JG8xgwtr+h
EX0aFL9Q0CCDZ1Zz1kcSDHtlWo4zMJFuiNNQf5AI0Z8ne1kt8BzUikw3cXoR9ybr
FZYTeZ0bxLTtrEPcpzKyT9shlDUfDeOwgGqZCmpGTWEAHansE6yOGOvyJwHZjMcG
OBVdL3wSYfqMLVeLk9QtCsiA2+amkkR7GUQaRir2mmjQ8UYI7QeGmJ4t18PGj0Mq
PWrCLcSy7bX2NzH3dosUuJJNy7m0nSV3HOlQHQidU45hcnop/9za8xzFn2tXd//d
OaV1ddsPzqsE2I9a7XfR1iZM32qaQWrZW/l3f4gYCQBoPqKBx7HLLDM7F84VI4SI
CIGV1ivyPHzjj8gfcI78pDV9qw4xGA3H3a2d+VhLCuZZHwq2/4jfys+be/Kf567/
zZ+L0zcfmG1lAFUHmk7d4Nfe4Wbb/wIrrO+wHfsBfoA7aF/QWLpYif/4/Kv8cAJA
dOLv3zJ/6PTYxJGR9sy4QKI/tOjs5wUTZKlzrz7iGMX3FWZe06yzMWHcs0lJYEO9
zJxOpb6hTZiWnr9wOPMVEpXYtmAZrCIEUaZi5aZBhNkZkQ459eGIue7aktbPMDZ0
BxpxOEE4aD3lYbhDbFJWh0Vyv+Xxv8EB6Yyp969HQGPD8ZgPoM6PhALUTE9uUHSg
26OqqKDQefz5Nee+mxy9OwKNtYiU3NS8iyP1ktEloYz/bHTWViebXuWHi/PH3hcN
VT3dJZQaEWw/MAGGTenQ7Mp1IBfl7LJ4ulC0ur5CDbJv6mPWuPssA43QYZmLqluE
wws8CLRifwKy1Ie2SpByBDoDioBSBg1AVz940f3S1fWajiHt09C+yOUpACgRDmBV
a6CBpUthh0TVGGfd4jBcmlHZADANJ3ICohSNnm0HykyEYLbHgXRoy9iTCWts9Kfi
6c9T5CbGd1v00h8OxxKawgRe+LTmbvVHLV93mDFNfrU5UE1ErW4XMfJz8Bok5Cfj
xUviAJlDvXakAaKlRFTfn7pDqNKeGqZfCrYxH7/jLdDQLhI1EZ6j808RiBGFG6V4
SMxCdhu/lms3Z9yacTn1eWt3IAgsZ3X6aD7W+uQ/SHU9RJeAgO2bLOAhIeAoBknp
rzBY3YCbdRmeDaQs34JbHo+4iRAx4Ro/PvX8STkwbi9g1docve7PAl0t0v4rgZXf
fqBrfRaIWTAqDouMyWCxNAcJKNU/CraRMbc55s9FdQU3kwBurOHbaDkO3XoFaxwc
4IL6wM10SL9jmzx1MPgZCq8NC5yifzTiDf/ybbxu++etIdLIzZTzOTifD224vtXC
2hoOB2Kqiu/VTMS+EEpUuvs+gjQ+fG6hH2W8qg1U00Yo6gdJJ6jB36nEjtd0u3Vl
ClN1WUgtvK45YVYO2C0WxfU4JKtp+hhovHM+KZOAb+RrEih74QaxUvL7yKhXMcBI
cpPNrn+sc+tZf52iQrQeUXyhgz5UcrkI0DAmtoDLerw2/Hw8i/TtXAvv4XbvA5vt
H4spGPYF+e6adBBdtegCXHgZy8O74/9C9fZgaEbRLoDT32eeF6PP2SFqJ5v8ZYF6
CYQTrD2aTBlw2qTh0apCYbAh9s3lCDeo8pZe0YMAramJk+n8XS6fWm0hF0GYl2Lj
+dctBwpsSkZf1BUbAL0g5fqQlx1/Xpy11siJhd59w9lbFEcUPpJev1cJLvoXZQCq
+7eBWbFn7uYMN9mioOBdilHWc2zje91YvAQ/YZdyTmDEfqP8l5AEk1NanGtXH4oG
hHGRDAKPY0Nvp/tabOfraWfHIXNXD9tmitnR7iZTxlRb5qZcHZ2AH9nIafJqT4p8
vcIkDChS3oPgOQfs+KFlIwo860/rxE5fQMEUWJqLQg3wMqo9UJskGR/5sfkeSj3y
X0yQawK6qQVGQwkHoOYs0VgMaw/ucPfmmQOpKc0R37xA6eWaYKYYDLLkEI2K8Y3X
f8xIUCC3YmkHnzsi2G4nJL8Y6gGNWammQ0lpEQ42OF/Xi4wiB2eq1vC/zr14j+3i
E4qXNFuJb68RgxXuCw4oQD1SP0S/A8JmlmSdJluX/Og/FFEX1hngeykkYU5iKv5G
6Hy4FPWzVUf2Kvm45nBgpUyWydGy/ACEmkeR8ZLqLx2KG2R6j5+1GsTb4yej7cP3
rfswttDhg0qE0t+1KCnRSAphN21KwCxtv2ntozb1pIcS4Ttcz4s8TlkXlONFGkMT
WlgCzQT0+nJ4tMt3Z9ErYYlfQqy+MF1pKQlBC7+wZpWzvW1TcWRkYj1Z/n5aIB6A
yJpsK/Z0Tmhy5fOr6G1n5/zxSGXXqmu912hLmy0BLx/Ny2+dnAVAsXfAor6wD42o
ONZtrnVRnO1VvW3icDqFbr0dGzy6y1ec4tJz2FVJSfaIIN4+uGXu12oUHCdLhmh3
mwtD121c6LcyEDq6D1KaWOhz+VP+YCrJIyMChhWeKRmTdH3xO3Wy0rwc6CJrPGG6
9785mcjGI+8DeUlmbxZoPZflpJLCfKRPu0WTYG3RmZoyVAZ7vl+BHmaSaTc7VyDb
QAegN4Tqraom69/gTCgqRyzy54NqmWwnnR+hVwn0gSnsiBORXEE0PHJiH0ZzeZmh
xE+rKY1rCUiQTFhyfWd488ovKDCFP9YanpckrxV1wmI3TyBJwvTCfz6i1Yu8jMg4
NGuYFZFx3hzcvn/+MvOVWUX47LbOfdz0Y12yUe0pjjIJ2Kz0G8lhm/4SC6/2R2dL
35k1KD9yZJ1lLyFnukIxvEN5IYF7oL5j4Y6PV6kisoGqpYRrfeUB+mYzpQXZvC6F
dIow1evO0SEtTf2yOcPuzSoBvgRq216zuGiboZe9TBShkJM6OqISAOsEp6LEKF5g
rCFxKsF44Y7emFN9O9wi+71CehuJY1l2uJNDguijRbaVTeRS8He4a1VnVlKE59/S
T2gC7N/ZhIS/yCg7Jklqk8HoHjRqe09aM3lwUH8sc1oddZxZ3J5+R2mYkdsu6WBG
LFEKZBbxHKOR6jSD2L0qJEmq9umRMna/Z+u+mvEU5S6EZiRTgN+PDNrh3dJTirTO
tb1bOsleHGblnWfyqtNZp/gcBPAoIAev+pErvFowt/CkdiEB/sG5SQK2qSs2cP6/
DU5zN+CV5m73Fpzz4WHgXa5DDz1oF3KVzOD2xYV9G6kv9y8go4ntodLCCiUsqWOS
y4wMshOnIjpetJ93OvuiIRos012/sd+H3E5gTzX6XZwheUU7Cjt05cFYE5Lq+aV3
hMLTdcidFhp2Vp7eZZGk1r/zu3y3bL06QE5hZuZSU/SKRnraR8rAVDHIC7LtWqeX
O2/wSm7kL0xUwykKaJHI6dKY3rWXa/EHyRoaGLObDHXrEfzCHZ7FUJP2Evsr+ePy
AhNshXbIiqFymLx0pWesCTuFxCmH+dy6vXW1Tr79K6HGNzI1yScGx3bC+SNop38Q
1kmbBmC4J/2EGCUDsEmmvHhn/VmnjAHCowhhzQUVDq6ptyQIigEEPnLx2HxHnaXM
Qo36dcaiVYoHLimQR4uyN6Qh0/RY4koc0zQGaVSj02veKPq41OfsQhmhedId6SdC
Rgk3Pn3WYBWYQEZaITP7Uqior2/cYT0J1g+bS0ZRm1ZnKc4pgpfho+GSyJAY6XT6
d8QoeTrYd5DqAM5VcJ24VvLj4iCrSR3NQvXBqaHw4LmfV/uftJ1dChMlm0c2I5lK
vxrZgLpqMMPqdJiNmU/G2LkDo98+TAVmVPCbUCG60TQ0IsIEYVrrStELeMIClql2
03IvrUNUYcvr8Jz3Vn3HUrne3f/GhzcsOdL3O/tJ1rl0O6cd0KssOr03m1n0Ca92
EWgdn0R+L52/MFZmisfVeWLWFRiLs/P4xij7UhbzgFTw1PwJbeV9qmoXZVCntHk0
xOYOFaQd8zh+buMdQaQmb8ewEDO0veWNWFKPggIHQL6utbD4tNkFc1wka0sVeABE
XCvdR1NBkjojdtbMmaO1kzVe/efasLVY+dEiHIguIRICbYdp4wyggluzKRh6dITY
yne5gCMigtJk1H5ELyuIu1U/ryJYnqd0z/v6NJ+AdgTEeMHdcgoutEBwJdfLT38u
v1RU2nG8KA/ZaS5ZBLNz2tgJxCSguOS5CNuONrNGCXjT1dyrG6k6AXWSBE5SArky
FjeU9j2QkVEIz+RG78TOiTcwwp8RP5J+Um/9SoS3AwBGRW1hP2cN4gIHIsZOPS+A
2elCnYn5dDqC1c5JvEfW0CnFtkx+UWelEHw7q8qa5oRIGdzJKIVXQ9EMPeW74Wfe
60C8NG7nGlZXlQ4joIPk1SvlJz54JwVro5eGZ/dhO2gRtJtBjZSlSsVoowaRQ1Mc
dCf9WhHbrgwrK7ufojandH9o8xijeCVzrvKQNvkyND21RBa3E9xwsEZ24iohxobc
i4R39sPsZ8GXFTuKkWgkSjlzv5+dNIoeemcsSgEyTXc+BC7X7Ka1Ievwc023emdi
tzsbEELRmpXTGYJ1ytammjnlkJO6T51TuxFOeBkHup/k+ZmsR8t5F//bFnihp01E
kasXyE7R4ASlPwKeLOHO/fqZJ/oM608eV1YnGlU0rJzVimi0hO7sCZW5qarrPVBx
n/zKmRYsJrAvIskM89nKFqNwO4+eSh20T/WqD0nqZCzjpT0gv8esyJvRMVScm13A
P3h9DmoltbZ+THFHWj7z3TnXMgQPaql+jT+JynyUBdpRCMB29G/SsH+dgMTZoFji
nzfu9P7a8mi523oIriwVHYoGmQfA3fKYP1Fmtg5COYYTr9A60nuOD5OVeqjtW3qX
ZKhd1kdb/FIXEzaMDzsJOnqcwZ0ul8L5M5jiPWYOgfTJ7aZ4YpiFkjQUKXZnoHIO
FZ/QsZEY39NYK16ofRyzM15jxKIgydRsFaCPds9uCGYH8SiUhPQW6TpGyIqGj1Vj
ujwrdwJ9xy9lO7ndfJUIcEoAKSj/Gjn1rw2fc2frxCozsI47+CE3N7HQsXVTvDFF
PQiMiVhW1FTU1f673z7CaLe6tI087aSZysvvOLPb1Ooo/fkYlObt/sjbKgB1sA94
rCOm1JWeEFRnSk1F1/bCo4CP439VpFznHdbmlwSzjUoWVMwZO919K1da7Y7yzVCW
3IHL8KiBPaO1XSBFLaZkLaP2aIA5XkGyBVWb+ReVnvZIwHfc6FPTFmosNa+GSn8b
r/ELkT5KS/EHiee24/5G+UQbkYPS+RUvtN897WDDbP1CNFd1gFLm6XigNW9I7dby
rJRFawRpb4lb+0mQvD5hIGoPjTmygo0sxCBlnRAF5YI294z+Rg+mw2i878ryftC7
6B9FNnZxq1eNta2whZvaMibRT9n2VZ0tsLt9wHEanvTDM/0DaZFAnLMbqmqMf6Vh
b66zK50uK8r2o0qJMZB/FjAQZp2qFi5jZBP6ds2YH9Ku1a+LhAGNWGGnZoI1JmkY
5uebBAg1ZFP0BENoOKkhXoPf6WPjFk4uU98+MhzMPVip4tOYoOTsVzZwHQ1OzC3F
cq2A0ct65SoFQSkN8sDGwG3PE+VVTPOTZclVC7RrSey04oghsiFZjLQBHJ5eLSwJ
xWC6iZqnjZg7Czdj77LZNVZukRM6of1gQCAJIlQZDNrVhcj1FQDc4FlQ2QxT/SKd
fGRRy+8zMRsDvi+s2SktBuCeE3ekNbecUA8lRm2QUoN9gl0GQT89VysQobzXHPNp
R4F5BOiwsELbqI6/xEBezU5DOT5qc3HoYurLcuGjIomajZwxNBjOCQHoanpKup4e
YD2UqNtdTQwLNySZGLTXqdd3WG809FwLrIByIF+ffW4LYCBophXGqCQg8/K1agDN
W7MAS0IJewzI5vkkMXjUGF8+HymWAORO6KhKe9MVJ6gZac5StNyiw3IQwuugVmUQ
d7MG7Nc8wJc0op1oJciZ6rrDmGKAymIxPGTE/3KyWqlm/uhhThjdoE16kryUiYcO
0q1MD2x6IWjXd9qxokXMceIY+PqFOqdk5M9SgTENc3W/Q9QiTf9hAn636ojblNKz
NjHWIs0tojf8hb91CWre57XRpUQm5/UqRYKtUBBlLwA17fW6fIFnBOZVDabNCRIg
bYhcnnmAO7Wg7Nc86pKIrdhPuE0PcOmUJFrHlNMhNRnr9Dc1eQ1nXdaEotg6yDRu
xUCkQrOYExAhzbKamTVxSfMbE0FcFOVQZDI8kkmvhQua/BjTCQx1173jtqMR29Xv
mO6l1QGnCPNRsF/GyNgxn6au5JtPbkfLGu2Ul2BtUgXHKRcbNqoghSaMPWCEJV7r
V2TKafQ4+XgRo/tM80nASRbD0dUEtJFxH2d637VMy4UeiWzDYlFAHo74avGPbm5f
LZKLnHPSWHnSKcwqq4EvUQp1B9kPTL//OqNkVNIaHe/lRdzJPD7Ekyv3KbvCL2ma
UNTeIW1mzLlHJ6a0SWM60lq6f3Md0rwjBh+5fO3OhdBUbFYBa40KUTbMrSUPePTF
rnUQ4PRbS7ZTmwV4op+voNZx9JWw8gwvl/zHlCRimdhLpilV2CxGNix8STe+2P21
MeA5uw6IzFWlNkr7uOBWJIUEqifu/DoPd5MvSteCi04xSt7osUZ5llf567yddXl8
or6Hb5hCEz0rMI6uG4uEl0SH9LZ+XQf9n7gz/kb9qYEjEUm15YZDruERI2LX695G
TNfkst1pLPR2N/j3X6lQSrvyRZK+wgQaOa+QMyRpLGQbd1QhOFquwfzb5GAcdSSF
FNNQeqdgf8RY39EcX7/SRaOubYlzU5qiLJlwI0SRewzBU4sNa3jn9Ezc5HuYQNnz
9ULBDjwBksW4nsFZyeCE30AlZ9LAkxlAn/YM523+o07Gdfh6nCiWv7+2zLew/Boc
GeAUrNuwZJpmPGdm9wr7s6aD48S0Qt+eVyFKY7gaLOpql52Kf37ef1KOUaHHyP8p
mmbjagV/vM/bRx42npWAdHhJggVVnDYFp/r5l1okAxKdrlBMPWu8fyHH/90cD+4H
QLRuI9UOrsHjYvFUyB9XIcYEbvEera6Eu9yxASdFizoWMmA3ybiXPZUgK66Z165P
wCe6i+sVqkJzshrQYlJvunHo3oCRCb1UDY6WLgLStHG+zmEL0tCeW9mdIyJRxwoF
3qEqwzYRGBwde760YD+GFaAgirdXV9n0IJEL2GpNxtRAiE8C3b7r7BJTz3ymXJhW
UFReJl9EvMqqW0Irxx9bHd0kLGcJCEveXig9lMFm9cqofss4+B29JQ9RxEQohcao
zZD0hJnCNQsemocnXVeN1RMoBJHzndFjDVjNdHFaJYbxfJGGQp6xzBscsXP1hrBc
E2zpObbV5pHwnpasCBMxhFT7D6T/zhBkVWWqEUB/gjYQKJEpChAv3WfbeU/kJmkr
NoTzbr3wnRwJ0dx2Dn7IR3oWDPDZ7h68ouQGoYlWY12Ut6Ppj9C0KTUvTUZt7n+c
8wEtp8yvNnEw4dI2eliZ4WmOunrUyYfODUoZCPsIwJ8FQzrnk+zrlWCJ7nTNHdkH
MEuDHvxjpEwkmbXrKemVernGGMCArz72FpWJw32myvSJpT0SZbSnDe30qq+TCEwZ
XKG2K8XkCxI/xoPHk/lHt5X8LHMu21OQNFTD3rsqyBxBRutaYzJ7OSfjRCeBUHYg
xkCQvNTAVfbJpyqesk4L75Hli5hP9W8HxAYPIfHuMmIOOO4bMMStIaW/pAHCDl/K
TSZznqbQykGANqmjb0EtNaPMHU1LPANL8smjFX2bNA44DMxzG2pkoLmra2orIiA7
f4455MTjgZPJv4Mh78pJBAFWwuv5kHbZVoVPuv+T1JkA8GJV9XaufAh48QWqLUyp
ynGJv8m6gJzqXoHQElCX4niH3T2U9aLTj43yCqwvugxD0/ltvBWC1byP2dpVcm8j
N9dv48rVGz6x58hP6zXPHHM6kjt8hLO27o1+h8tHTgwtZz831EFsJwZ9mWddogsb
256DO3zuzBgsYTxhnnfvA0zBblCMwX7o+Ut316ahzPinqjCAYTmiWOs8CYy17VPf
i95eVgWpsNlC8gCGJtMS5PibJHWm5fo+Q4ztdo3jHp6ASIxMKyTG9+ekWZnZI0t0
Vc0Zihsc7qi9L1QutElh2er8pznoYBCnzmdSNsYw+5Zb+cC2jtZtUjlL4dBhpXQd
PJbhsEILbPkKULDNKWE0ruCzWRzv8s/pywGKnlkyeZ1XtpE1UnhQ/svW8b2xPq4J
pNkHpWvDcpkimEvv2ivnCw+OqT8TMvpLpdgBc5eIA1cBfHyjgm4wf1RFVtKpfXOs
D+M2u4Eihv8Xgou3nVQd2NB/6X7Pv3JI10JcSeiqm4jKeLzX9QImniQd7dmMLhlu
1IToc61VqW7dOz87BWqRLmEFcqHBEud9zMX2CwwTk3I/NSSDedto6OV1gtoOADq3
ITmu+UAa2sxNmD+gzIbvNSwIH4h3cGaXIyItXWKc8JnOtFeH7+IOgFpcK+Oz8vct
nqZs26S0OVrkoocDj0bMn1hFE5VlOOoCgpaGaypkC6DulwDWvwxfqXYeutLGq7DM
+DhnnUeTblxyN/MBaEbWsX5DGXQc04Cu4r7bL7JC3ggMcxMWnQzO6ZzUZfWFkd1I
9w1bmaMpMlQZlldKIZKZAKccehXCsjfd7KkVvZUwr1fsckjDPo8k1YOFuPEVGlVl
qtT/GU8PGPyIP6q5QcOqCySA4RLbJX0fCcgP3YfOdIp7mNW+5ob64SKuKymwF8f3
nV8P+pf3Uehgeyv07bEtbYxs6MYVaY+D2g3vg++aay2+wc9HrkneIrmNJLG5tkkH
527WkTuNs1UYpxvfcb+0oK8Cd8Jd6mDFuU/Obs8q83cOpGwUhx+pVAdZmPHRnDsz
4alr5+SzJGI7QHJ7c+bnjdHbyThlukf4nq+5jg5XNpBW6x/R81HS39Cil2Hf4z3S
Ys21uPbxURPfdJsidMy6EBALxd3in3HLvo/nUc5WeWeE5zbLVaK177Fa41OZwMn5
LsCQzySpt4DCqdQrOOKLLbv5z6AYS9t6a3LzjuqsK0+301PY00JH18ehvyWcAXT/
kVE2lDN+24m0pAsKnbO6vemdpX/9RKTV6bolWmXf4ZB0JkOtQvu/fA87ycjXENE8
s8uJ8GuiY85Dd6UVBqoeZWVP+RqM1bi974Df75Xat8XuyjZT1HsA0UAX4OBW/g3O
MGjzzD0wGHFQSSzd0zDfF8NblFvLMwz6cRRlHMGvnZY5fykXlDr10iz7Sea20Kwn
WVX9yMCgu2lXbhgO+oeJkVw39hC/llezvVfSenVadJ/okq4iOObBqpHSWM33pIGt
N9r0cxULQlg55SFypNbyHNtKgwI+zRA0n5QCWbnfd2kN+ck9BSWviFD8DnZffqqq
vEJvUyy/v7G5jIJjZYsTDHOLD628qS7IbvE9DzupUjldiyGMx7V32MkzD9BYy2xh
16G6sTKYMlMNTwUY3sTziizQBgmoM1QioMALhMk7x5m1fIhfOSZhQrqalrPpD2Ai
OiXvvKByMB+bnaakwUEV6zARoOd7x8KsAut/Yq8Pdj8gWwu47jiQyEK0JYH58OJ0
VaCY16wEmbZVBgxSO5WAjf97ujWgkYTZxXz2I+mMWCC7k+17JMtnW29hphb00fEg
sGNCHK1j4o5uIlpnTnTX5z00oamrNfncSPg+N/JLps6saUdfF6tSJ0c6pglL/o19
4QAIimD+dSrG7B44kRAbFSi9rbHj3Z6b9SPNz/Lrg+aWC+r7JxcgmryQNdARukQu
1RMM4OhF0R3kgzpKv8Z+4uKR/WBkDJNx2q0LamkviUt1rznuSzyk1TjCo9wq4j7Y
gIJTahDBiXqOgIT6xd9Cu5yxlrCdRdY6MTWngjHJVzXYLiZ/3MAVy+lE0/W9pro5
2yyI9ujf0XMYJbTFO6sLEDlp8y6Ig9YC7dpU4/B6JiPOSpBgNNf4fSfdzPpRl/dC
bEW2ZqlaBZOw4wKSVjdl/aRIg5C185mDmy02MGvFZRLLK/BCDyIkvPm7dZlHjrfc
aEJm8QQrOQaZ0FdcJfwy1a2mzPJgKNso/t3dsoQH/HzG2YY5YjCYQQZORJW+LSqR
KOXQ84o2KjRfDILxR6jO2xafAFY0XnPcJSoBP5l8o45+IpEm0uP9dgXHDULAWIOq
uLZsEBKn2ObRp2zHZEer6RzFjKoulY9m8duQ08o5nnQGm4gEP6sD/DeAUKd9+/7f
Kkp1zKCXF0Yoa/rSLbhpdWn9PLI9IyK8PHauZ18vUSTRYqxqopPUAr/wSL7y4qKJ
s9yXsUXPxcGnQDOYUOHuL6Ao5vZYNzrbDiaefqRrDRIucpGsLENYNTFzi0ZedW9H
erWZdruuURj2EZ/FfZ0anvm4kOoldGOMaqnuYCydY/HF1OxDtAgSHPM0mbTXe9Ba
itXWzbb6FBFx0bkP1FNX1cjSEde2KlhKyl2Ju+iLSInxMIns0NgR69OB4P8VqvZw
Z73Q+BMnf5Yulg9KSrzcfRDYPrkHYVjOTNlsu88d8N/MMvAFBm+/wPSXa3oorujW
quwM1kO8N8Fsb/aJykIwaMNnApgC3nijm9zbvXr8JtK3f1bU593SM5HnLhogmNCA
YWYAy0olddhf7sRC/6fcPazLDljJItfT18+sUSUvkDjiq5oDwEAzMTt8gi5rAfma
CGn9MsDgImenBioOTxzbXJT0xW0LTNpLf5CQ9q2iVQ2zfbitpEpfpW4gwylun9G3
h3lMRVyB9XaaF7BocJE3OTnJnz8j34EU6EqmeDuxzViwdLw0AYJLKTkdW5Z0/vXJ
tqhvCxSN4D4QwSs8NOiu5K0spVUnJaXTpGZsvMrhtOkiLkFTx8NiBDFHQmH1DZMF
3oCElK6lsHzuAcdP1dNFpy4fxQ7av6wSUgNPH5whHsht+bSl3Sqo+S9thp/+2iBS
0cLciBemJq4eADb3+qQubAl0cW6YA2x5GLK0FGjhltpN402L/WmOb1IN2aMQfgq6
zankUa+oRqL+ck9Xjq0FdkjKI1OtgRjMdHiTJvcR867b1qWYuRmQfFEzGS2nmZl1
jLwF4XSbkV1LOY7sDij6aX0X6jIFdKEgRmIl9oPflpRo63llPHgsmGKhwe6BqM2y
juOD1ASBEVz4g3zhHraRoVRdskUNFl/zkIrQ35pwUZ52Ax9kx+7oJj5sQt6T1VUC
ULPF20AJNXVov3tuLwa5VBEfZVVoaa/mibHp5gLSulqTMJhd0m6SNyq0ma/GTyKq
haK2OJUyMU66TXGH5HE+r2nCe7weZErfrzMYAo4dVmIUuZunhQQSd1l2bbqAoFNJ
xt6dB8eCWHdhdkFURnv+YT5/UY4ciHRY4vuc3iHEcAAfG1S5uAJgTR4xCQCaQKzu
OpPAg8wldfhmY8YWsBEuUcs9/4izyndTm9Nh1XP231+ENrMaVeJbi1eAI2QS6gF3
TF6f2Poi0SM5vvIQENpNW7jhVeSA7aFJxteWy6RsePlhufu3u+oq+z6lIpu8aFRL
KtEivEsYUZAxeIJytC6v/jzk18o3rkGPC2XFEukU0TUbJFVMMUYQdTbblrsyhgP6
zK2rB9ilRKKj9w4Dzf6kgtCN761nXDorG19SPdQ/+qFbRqlyh4gKdjvLEhaju0kf
KCH7kG7NWj4mlVRgE3TrmR/7yNFuFj32R31npcnaSX4aXQaFXgwcimvHdFbzgj+r
N5RI5wvsf/kWKOjmyZKmXXRFdhbNXWYYAmC6mzVPitSp0fX1lDh+NlGLEM6vd21W
nxFDwKC3wCLkKbzRmk7Iohl5VY1GdiwdrwgBHZDGABcocIDYpZZzxbkH+YMAdxFi
aId9t31CpW/Rz0CW0ec8WMCTlNluMEPQ9e1qP/652Vcmghy7NNkq0Nhr54iXqIA5
umvq3ViAWD2yD5NNC3zKLT30HJF/misO3pVp+gubHF3lMGW7BQ38WTWJeVVpllYG
8w3RbrGDCJ8wLMBpkj0PC8umzJOKMEVKmrd96oTWT4nkjWI5d3kG07jtAKb8oOhu
rk9FVZvrhdgqBftvxl4EgsDzB85Zm5DlaQP4Wst4/+Wqwl9rEK6veHQKjlffFI0r
a8WGwZZymyYspUWB3Sim4CdXYIjhI6AhHeKywSNaEoPmqURsJcH70MrALGEPRbYb
79AmYsYQFYsREUxFDIHH03zg7nbTuF+S/fKwDwntNkwZue2rdKwFlIQKWZf56TlA
3KjTkuozH769tkpWXx4BnECHaiZWx0d6LbCCJ6Wqzffp3SuN49NWGGuXn5Yj4FOM
Cey4dCJkWGarMjfsr25GMWPyh0q9+fu3RqqXnZQmFZfQdrarSqJrHw0/xLWMyuRl
qcjDv34BRWwsd2yYcP9hdNXtix4Bu4P+ikgoNm32bzqnUrz6fdlgVIzzeUXFNOiP
ieejINyayLO+Z/U+wfaPyHpI44x6QlLHOQQxG3t/Mf6tewSWJKG6VV0xtqP3cJ/k
fP0y/ABkZ37tiSR1ApD1J+wr6JTe23z/ReyyPq60l00Pu5VLrqa2EpNWWOUEj9FY
gy34ZqeXtOe/zPJF9jhqHSWL7gBT75RD9NyGsXF0FVPzlwpihnXnY46o3Sgiz8Ti
ouDloTPBHYRsz9n/paWP6iBA26D2lIVBaQxaUQmlsDSGClmljxj8KBDSsSgpV/zv
Cb4W0hwqwpekrDgzuqjvkCOVezYSoABD1hSLb+Vc0UZrdW0rhRYCzOkSPRsScLNv
YB0Hp4IPeZBtMPzHXp/hHdv+12g3R4r0AxFGgyLQIKhzMwvvCxOa/88pwx75znvk
YM9PWnmmR21GlAuI/YSG5FpsnfX+ScbdYv4bMSpWSTKAborNpf3TvhvQ5+TYSsIy
oqLhkToVNcm+d8vQ9vy/t9sPKYZikk39MLC083TXagvY5mZK4Uwb5j5yrePItVL9
kBIeMMUFc60BYm4XkhaMSOUS7ufOmAaU0LZxwtY9eEs4FGI29G6URBI19lbOLFG9
Zf+YVuCtmjsBAnsBZ+sYAaVQFySClyYOjkSjcNlEFcHkWGH79iQ853/ctkKOeUmE
W7zQyNX/auxXArnzoM4LkST/HmriGOXF8q+mQ3yyU6Q+1lcerk1exkz9LMKEmXyL
IReaO4nnQO6dO8FxzDjEd1dvBpwxXI2IT3B0Z6vxtux6hyLZEFlDpBdt5h8Ls37T
bOyTcCI6UJWC9miDhyojDUwA5vimalNW8K8ZsfRRCJLYVHvkT645xTVAp7BWueNH
eJIddoHoE9LCYZk95Y57rrVSBJvPHpM0j6u7kiyvpf5j+TS4kGHwwI2eCaVMOTN0
nJXwE2z1tGKq88ZtlHlPUdIhKXyAsA2uotlGLd7QIJ4egLISU73wIf5a+rE7ISlI
WQ9c5mNVpZILXUA52LwuHj1+M5fA3OSRtNX+jzoBNENKEY2PkoAOrY8i4LlmWXNj
mU7QGyBg0yKasH9BeQ/vJ0kjoYGVj71MwUMGJaIFIM5SCBYjJfmvX4sWW52ugMAi
LEv9DqhQXyPzra8YNZKzAFj4hyOrFHApRE3PAV/RFn7t+f47MF+ItI+EZBFpn5UR
y6UOpNVPWSnwmzH8yP8NYJIXne4NvrUAayGo8BvQuC2uXsriYYmNm8tW9piKnp6j
AYdL1tDs9UR2lJI6EyLJVKyHzvaVvgoc2Q4faNoiIhJcHUywgTNg2GwinGu3LG0n
1bHDpbQcbDi5Nqn+NWQu5PRhWonarjsOL9DL56C5cS1PM75PltVcYNB/sqM8GZmz
xTd6Rq9Ph4i6RGJnvjR1XUbVInxTR+5XUJwZsBElwo8neYZ1ntl4loRXijzXqYG0
L3U6/KFMbGsXD0CEVMMbPDOgDWJk3LhO8GSE7RjgxA5hCyxvlNtzegfUGMYSvStV
sY1K+SUNkzUUAjnQ50SlHh6o0BmbCPIuPM7u4y67k4pHPN/F831gszeOqeLKNOB3
l57V/pG3HShM13kreGXfDwO334AutJpyLhuN9eH14D6/7UdsxRsfX9PJ9TobUlrL
FbB5wzuV+wmhDSbljhaj1puVnJUiExSfVcp6ssKPawQlGaBskU0hMdRPb03YaBE8
bakHM5GeXizV3YAiUxGAYvRF3BJSTf3rseAgJBOMHhEr2YOvX4tsrYKwzAOcVX4C
CfglnEKhtYjGIXGIS7BxD/UTQj5tLknHejANVBAozxi3oCJfVQajUNK9KqlxD626
Bla0WBAP6ffko3BDx5kKe84LFiiFNAH0J+lRjEP59RdVhNuvm+D9igVGoO5TmGGP
iAR3jNHx3e90jCi53PvFe4BXvoEmKCbgG/NTL9hkVeR88qWYGpqPT6AEAlqgihsw
Ygl0Cxhn4h/QGmpwSX64/TJ2RDH6Mfbx2WBDc1FdGoUT9mUGS8VGVlrWV3XX4Oob
Tbxl0kYIQH5SstoB75I2NMY8JbGOnfR5hf489yIVvVLbU0s4+NoHGY62z73eV137
momKogbmJh2eVzdu0IJMCbB6T1aVarfYaSwcIncFzbMI3PVHMHo/gp6obqW1pAwy
nFZWbRtalzmb2/WKAy4HMprBhQh2xcnZaQBEfELJuHgOVixzq9zCK/6s4XmDU5eZ
aevcGlQWw5bAPCtazyVl8UChPGZ3gLos5pOBLturZzox4THFv6xap/U1V9rGZ9Gl
jfnJT8rQasfIzYp2xpQI1XlI919vX6vhsoDbMyqycKTF33fApNm2qt6LngYDov0d
rH0wnoEqJlFE1Rxa1IJ+2Avr0HQdG1jLBn9tBuFcydVmhIk0uc9VXCHj8F5b+jA+
DP5MGjPXcDlBQPTUMPB6gwaeO+13NKRgZpMN8oQC4LKS7aP7L0IzBeIY0XDaYopj
NC9ftBqsbaXQ8CKFBOpVf1uVmp0mYsrAjjvYx9I82p12IXDNTGuNg9hl0oCC8FS3
5MtQNrtI0/BENSdkbf6JhIfcM+KDrrzs7WYXDt+C9moFKfbBvebp0QnBwkJaIlpR
Y55uGKDs0PMe1qdPQl3faTwuD/IZuwya7Zs3aPExoTlveUf3qi+bgUFGpsJH7iHM
tyTo0SKI30HMFYgojtdO6J3y6+5AFzy/hvmwyOsYd0B/MSN/HjfoseH+KE0yTti8
/F0h9gYISfuadhSF1LiDp+8XCu+eIG6zmUOi0wYLppMuOvTGEbdBrxc9iA8meoWS
AEiA7KEHwJWVJaPu+G6o55QfTKQUR76o2D5rxr3dWRfZWER8ZULPiweQKz9J+BjJ
GIxVHbVOl0qhN4hTEjX2UN2zvELdWU/ObmpZ6vb4lwDv8ss5HcjtYAV5xWCtf3dl
3K2o2Mqb913WJVDvZLh77UuG/RaCklSzTlONcpPDBTlOdm1C+hOcv5BDLAWjrT45
IbDJGZjcLv0HqTna3HY9bd/BxHZuEwUavxdkQUEPHy7hfKnr7hpAhvc+zQUeuLMq
D8z4LnOBm4HO2p0/vKOZyEeQxM304CKjAEvEAuFiwey9foPhuLONzwY6w03/W4uG
5cZWYvcC13NKq1M343h+S81dwxyI4fSRCUQlnxTpcCtCgY0UAmKGgTec7tIsOpm/
bgbAauzus0ArAaG+ZeynyNjFJaQnK4Ov3EL96rjYiu4RubPypgA5PS3BwlgODH2x
7PL7aIwdxaMAaro9XXggYgs5l4EG/bdYZrHjK2GiNXuiTbxpBWj8t7k4fCyVJdMD
gG456H/69WKLKXiQ2N9Lmr2CEq/iY5DrgshK0E3R1f/A/dihrZCC7JxvysKhczqD
eGQqwowYmA3Yte6/5nulTjV1B7k3jDWoJv3czecTidSYG8esZ8GOr9w03LIdyKi4
evrlbvPGmV7mxRmfguLrLTOlyrxxxO7ZSgBMf0fSmB5U3qYf9tsAu0S8D3vG7NEm
x3f4ed7VppW/2OFGC/xCYqu5l1REKfpCJm3lqYNx5ySRzm2bbBKGkSSeCMQeVJ/9
HrHneRam+/GwY6BTJ+xcaKqZOXew6VBE0puGO9y/29USvYSLsDQ8aUBm8sbkIfDW
7bTVsPdkLYcLHzuDIRpxpEqXbLz5M4tBt3V5OSPFMrRTmnEhSK51/ejEA73R0+/c
aO8Pi7NFRDYCS6YQCkxHCdKlVuDZZ/jqTDngU/V4nclbt0M5oa+uazBpqJJoBsCs
xrai5vYhuXjp0sedQ4a25rdzN7A+26878grTn6j51Yp7XFOl0C/TODpRzU6W6XKq
av+N/6/FY7m20habVoYiDeJis66bJQqZ0aPDFG9FQQ27qP8VMzCZM8W/vJ25Ss01
/Aw33MaHVc2kwgWZJPfWPfUwJJHqxVAYlz7Lbc1ynJ7t364WpMR25okgHqystq8b
h7Ci7cvJWPT1YVRcTDWPuWDEY/kv9yIxh4FDJC7QAXfi2d96jQKl7M1srkI+U2BH
XTcXhR3WjbidUbemGmM1Abi0ySGE2dcxRCh0u3mziU5HeGdk4s+pdkcFVD9BvWup
W9FExI+L2mAWFAHZhufVBZKJBwq6OwbxKZQ955B4cQBG2Ap9N3CbWk9KSQp321kj
7SVYIz6iu38B8mARb4wACoU19yIjYp9qwVPaZmfZ7DEj3flKbmOMmddlxDsp9cvD
/j3b1TZtTh0t8uIWu5egJMWdq1Ny7Aov4qtT+QfKfbCpknmj/s82OJ6TYzJPMBh2
SGJ2Qw4QoIwkuDeHvxlt0hsdQQja3H2Jlocv8ViFHd8TSFkuYmk0Re8nrnvQJgQt
blmGNiCT45p2PrInBeRfdkYEGFx/dlNFi81khS/9kNgRed9xH8XFEr2SYxDMZLcW
NiMxaBPw/hE54NM3E7EFIWoXnRCpgx4N+NQoXLVUkDxw5ng/jAP/d4yXY8VXBUL7
GRe07u/qEWLnCvLi2xLkEC5bWKQerA4GPp77EJInLUsCKsd6L/v4b7ieOy7IJE1+
BMLVX/juQROs7lKDUTpzWw7Ze3eq5voS7EhY/r9ybCOXQkz1EOA00bVqhM04GZlV
Pj/Z6V2DcSxBBIJ3NXg+ZNjYft8QdDF43yq8jEHJ8Am0lZRh+jdDsIHOGoWQYpmJ
UVgusAtCJwQC0Yqgvxm65pd28KWcDD5Sor+OinVGW779aMEX/2VNOhc8TexJ4qOU
XL+4g+ye9w3xg+YMtlKzTOBsaJYiJnahBsW68FSEOXwIZf3LlblA3KrCIdolcQAV
IeCLLNCfB4ZrF99uBj74+pnOJLfxh5sSenQjZtSKeaisqPjEDGeAhTdo1YoVSAJp
ZzlQMM3JZFOE0NT7SAt+KO6/hivxchhE73rk43smRHtyyxzKDsHnHs70Hpv25EFu
eDj52fKwdFyBwshLifwiARjagQOsOj779VWtIQSIp+QofiQy80fZt7iIM9dC+k+X
LnojYT68asAoY5wM6M7MzcQoi/F0aKekw+xd4Udm7KIkka6f1vfRXOb4oAp1qSJf
7f/4gluCtEQ/9r6t+MZoMNE5xY+tRCWWhrQnbPWQKsATgXfj/q9Qnhu1krAHoiRI
sN0MO1q3daYY90O/q+n9LhDhVfBdjLHCfMKwjizwCwtykJIKG8lmvoJjH7I5yXua
mUUq52C2gcLWkO7ZtDl1voehMqEKH9NiBoXjDiL+u8T8SnefMuWhgq3QLxQawT29
nppuDy6n3F0eyjfZiTrCkhRh5LAp/ugDcMMPxaVQijGjhagVzVTMBrTs3T9TQ6Z5
B7qC8fZAn0Mb5DT0XJ2XrGrfNM5a0hOejLDVrwpExppBBoOF+QAvgJGhd6k+Kh3v
ky/XzWyMiVjrKu2MRVL4bKgPRTX4OuHATjMqa6f2eeQqG8EMSbG2W72/tDGcnxg0
85do9hwjMcKoVf3P2sQZqCPoCIARMdEvBivFF1GF9Ne4b273GGCRtWcdvKmR0HUu
yN+0MQYV2WxV9QBKJN3AfVvcOGDPyJogJbVBmJaFrl4j4BTEm9Ess8sFRR9cpqTJ
QCpxA0i6hnw2ZP0gfuDDHIl1xHu+aW8IVYNqxuvQ87RVYx9ZZRcSuID8kSPduXGm
KWCdHnMfCQNznWw8uaEnn4rKiDmEXw6xIT1F91maAudnwsGaFvrSFL2jxmyBesYw
ZlYZEpOv9EUj/x0uW9bXRkD/9LcO65VRiBWjIQV4vMj41hL3jv7MptxQwuKdZTNV
P6sHm5SImwNq6dSJjnWLiBKPKbPQqAZhpS/O40LkHwuoA5JxzkpDpBILc27/MFv1
kPPGcc3ULI+vIUe6ZQxjSQZX0FMIpBN1yHgbO5dx3zoSCOkIO5xo83IvIUhdcQfs
dH0xnIUpcY5PRcuBbCSziTAy7QDjVg1efplSGqRO5dlxd+bqoCCxBkYri9+dGz0L
jWOVpZOgslnCDMmdy/O7WprWrR5MALKHiRJy+JLHICrzzN01ufsSjMulzJDljNEz
mZhatCNAqDem9ltuwGE6u5KZdiMk9rkfivH0IjTZAJrlv0hfArnYukZRsZ0+ooJk
pMwOEuOc+pn+VwzeHSozQCpXNtLBlQIKgVs4ePEzBeHaKtLJbXZpwigQlHaVRmYt
N4Byjdzb1ZLqnzIY9XqtLoE+oNPK3BA0gMhypjtalV0p238I0oKO7xqgzMrzrP8D
CkqlvUxVf4b6rPZRKUlieT/2I3AXJsrzQqF28k8hDNpQLYT3j7KWKy7SHGuZiOwo
2Ens5yR2BLSCPjOAnz13hJTNacHVdk0U8/WIN2IvHMDaquwbvXtYWsJhNP+ygQ2H
YeFFeH9DLuUzMcknSggfG8sl73+Z38FeOT6MOsq7ozDK8NqQ2rkv+CL867mnIkca
Sz+P9Zn+bzWIw485ur3sMvCjmlfVKvcKR6ZlgQvx/IM54UbdXmANBMeCwdaSiiEI
rPNnjJxpYEIRSQGfV6ANZBLSV8s29ApspyLHdLmTXjbiGmM6+L9DLPR/4dDCu0dl
OTOa96m1/woCp2jvXoviVRfB4kVTbO/jQJkmjNj3v7JV0tGhzCCB4mgQsLhuEW4s
wkZgH6/ZU/qV4aCSJc1ShxHuFHJE2GFICmtQltndL2zwIdtiLcUwiT2B35NsqnMZ
N6Lgq8RmyiatUN6RUw3OpMWGnTZ6a3wb5C0z1nmqNaMPGCmRi3hFAKB+aYRL0KLz
GOO3N4r4hO45YrKB7dCZ+CRapm7/wlKvofJu3mDtlTbckVnB6hjBNeMwW2t3+MhV
Cb4kUuCQ4OePX3tuhN7J2ZgMkpmDCriSAf4ZQQTmLzvwtEchLDMrBNy5lFr707gj
OXfA7JwfMzrfYk7nL/AUBtNmT5vN7K0h9hQmMEmQu/RpuVroNsAdn/sahQevA+d+
+UeNGD51a2VcoF9dDT2hO2pS3MB6bn/JqbgwM3pvVxFQ5+M4gMmP2K/BGkYsCvF/
uMoZN3AeIR+NPa+9tdk1tsZmCG5VtqPf6I5fHT5I7gvxXSruCk7dwgp45lIlhzk8
yTJ0eLWVltr8jLzkfKnWTZEGiNWixZ40JmA1UGvYQwPGKeuYIJi6r0umBUncAvcv
epW8NeO8uSNTmtjWkrllaMkIfq0yiXHQ4eGM7kos8Id7Vbdi4/UM6wKJ4RgqBW46
gp1P97/msQMACwMk6nX9f0hO3KsfMhZwrWy1T2cNgVbyenAMmN6cES7XJYI5yxw8
kIZNuAk+og7X+Upw0fmUUdp7iE2+P8NzzT1Tr3uqucB4N4Z2UJAC0zNmVgOnxIPN
n4QiYHc32+PgHn5AMqNF832pMszQ0Qt38h8rFZKwzLas5CLEuk+Rdjb6LVaZCIOx
+xOfFubFDoyAgVljmYOBt37WCdgVP0TIcEHV0HlBBHawWTFqRXXuTingWeWYPAlk
CyOQyU0ojbLK+IldliHn0fKDYBdFUWeTOqrXHFv5mbeLaUl1sN/ZC7TIs/UhmsEG
x/kcclCME9yq9dzpRgoN/LlJLsJtu9FtcqI8oLGEJLyzz/zKGSvzFFoihQyIbAYe
Gud/LrJBgeWV6P/9tbe7+VBM1zNHlYumvMsD3cnwjAcV8XnHtPPBiMZu5RuaDgae
CeUb29c9pWsywTdHFGtWmeR4kMR3+2M/j/CFf3kvyfH7grtKSkvS/stprZizZsBu
SKpgynQKYURQmwRXffjapBkJTUt9JHoWSSEWYvAmz1xuJ4Z9nj6gdB0FfVMpQ9Ku
24GkgeXRntXgMu4CNwX3mKnbpuIoGXk1IaoBAU9uFY5BEisEMdeE+ZBYCWKvxWa0
hcRoCNUOi7p1Jw2Wu6UjKu+A5Zrr4UrZAWilEOHkpdvCFT52xiLvtISiQvMy9z/m
yB073Ya5fAQJhn9lhyZs3uah+bz99Ug6yiOyD9lNIgANmzszNoUA7RwD6XJ31snA
W8yEqr1xME+RDnyMArtVB4MFntxCiFHDIPeQN6wIPbNfv4a5VVD+r+FrmYDVixvT
CT8K9X1bq5dntEk1TZ/95/W4NhpdeankxW8lYyitIJTcgREUYWMIDUuEug4Cdzkq
dYNodOJpPE1nGZu8z+CepAb3XbTJohd6zYiPCQ6y9jnLeGrwxkPvPD8FmCeociHv
Zv5BijZMzt/HtJ2TKDgLBG6L8Xai+rplP4kqCx1M5FttaXekNl5t1HrMcVZehn//
AyKFD80SKSumwlLQUr4U75YyQp/aiMpGA5kFJ8Nb3V/RfhIrDsJjRE2hjl0g5X3h
SmB2LhhxKxoc0zRbREwuzLNrzaHlsqSbTW9MBo5Kq1WxZYL7eww+tvMNxyT1n9eY
RLSyzZKXFq02TR06oVRZJz6LXkaZzPUBF/HYsekaLRyYux4qLUXTeBNyJxx3dIXL
dJ1EoYQXdlt7exYGjnWr2kn4taxT3kpfViWwUewSXvNGpjxWFFm4VQO0PpTeLWQE
nTf5RowbLvn+f0LYKNF1B0U90bZyirpH0zDlAo2zSmqLMVj+s7w6iJKdgBucJmYK
yMQV/BI0g+DkGBEgybdR32csEg11Oml42wB6YIw30l2yoHryIrWeDpQYK7xNpa1X
tgBSFglzrVxcg8zpzE2Nkw0q6Hx/cCciH5fK6dadPd5LHXE7VLcYqRM03vZqgYGl
KKP/aT1r6+0YQgaiUZQbBviPUjzcIHNhh253+t+voCZahlstrZoXC8NfYJs/1Pnr
7JOC1IDYbtoJFrr87CJNpoViJzH8ziPQrZDm32tkE/lRSgWt+X8H/S+ryq9PB3n4
9ZiaOJv+dXSVUx6ulGSQ7x5I519jrrWqt51RNy96IHyHSyKfeEppBr1BCqbMG57i
+HNxZmj9sa5QLMmYWkPhOD4Q9fhAVyibIQ3OkaRidIFrQ9hsUkIyw6vBmnXpgWOm
NQNhTKnOWEXP4ZWAitv8kuVLxvkz045yvE62QfFPK+dGVo/ooBta9Yz4rQVbvcdc
jKBTj8K7lodUJ7QhPJhf01RYbNGZkXb+1nMqjGqlcxhglm/GxPgRbLip4T/9Y7y/
D9bQQrI+WMHvCB7Z4dvM9nxsE+Jridz49Bih/8S89ExX4YnDh2zownZXS/TtIZlB
GDqs9p7Cbc0tpb4HJ5BMz1ofwBvQ/XKzqPt85i7EIS3e7GaVXTSi8IgMyAiqTEdT
JhsPLd1heiIXO3e8XNL5J6n7zOY7bH+/HfiQXecHuHQAEEty9n2djBe9X1jOQqMd
yczhPrUF7zFubO3YhkSSmASjDG92RWkqa0QwGjoP0Qtt+bxHo4fHw1yI5auh4Yti
v1EVFI0g4cT24YFbcnqmeJhYiF+hjZJM+8hyBEeRrNe5YfzTSMh2Y68wfjz2PQXk
mfpyqh32SXreA0dsydgAiBwes3lLjsHboz3e0h6nBQ5QU70ciEoO2osREMqqWPUO
L1t8s1/zuKEvArsNS9za7FnGqtBx0+teAtujfcTrQZGjkXOmM6fIDieGtPxKOq5U
UrSDCtl3C9nef+CTlc+YIcUiBPVjv73Ek/igDK1UDG4zIBBtQATmUsqmahvbOED2
nwkvIZXv5dLw56domagpSR1YuqtVJQmShGyL5xauKNgA83oXbdOUmtxoSAhi9VT6
C1jtCdolGz5wfPmyBrG8ezv1SO8q6HkQG6ONeezmxeHcPxwv43Z5MHqpdNCOhL0w
ox49rotLj8XAG4dbqbLY1G/9rWe6DftYEgEjSurL8nKfBDbq1f0tgfhy2HQ4D/4V
FPatN9IZxuLaH3qX+cBexGbMPTSN6saWsxxMZgTtXvr0fzvJhw8+QpqjgbkJrKRT
SxdOFlPmZ9y7atxbLDDQ/NIike7EhiOhbBTYPwZO/2Duevs3gm2iq22EitauXxAf
KqO+CtcqaBIpzvKtKcrp0RILLyLMxzynSoSaTSrSzJ8BCJsu5R37kSCMdfsDehdE
5ZDTI8jrriuJobZJ2tYK/3b3S0webg/n6NqPSektXtLcPTkYbrkFEfXluIu+CfhS
P2tH69JbF93d1utD6pyqr5kdUf5xcoo3tanualEOPsnaCAbFrbmqTrkl8oeyGwFu
Qiy+WcLeXAntzjI7YZvUWzAnU8zH+qW6glQPRbu2ci2SpnVa/e5VJBhUY+JiHFrW
4BU5aMkvSuFEs1/0F+HINgWfB4NESo0LS+1xQoWFPgJ32ZxKNrAavTPX2ADgvFNx
VeU37o13QZsXDK5fj8eb5UIKxyGMkXujVs6jCWnz2SdgAoOuU48NFv1sjZrdQXVI
L59+uyApFjcwITpgVrR8LIE1IP2tnEESf7fFrI80Ldj0NZSD2W7U0BB8LtKjvHYi
siSI2DW85fGLgjc4C8PkoixkdyZhjuUwsBu8nfbAsBQURkRFlkjw/RcJyhwU8hdg
H/Ga8z6CgNU/06Y/aZscUtAo4DQ/+u0+kL0HOxOq3nWkb0GQ6uiswN2QbEZ31AE1
cx7bw+ej1y6KvzbS5TVnJ2F5YoImy0egsfIg+HiCCEp0JD7ouzR0YOx86fBc2pKY
N++GneKBvS1b6TtqEyilMoiGeIsEM4mH93Ji4o0/O957Ln2LN9Cl9SQE665CT+k+
b/U4bhbpwcsV+vek2JeZ21VN7Qbdibz2O94G+tDcYkxzI7OScJ2mNOZxejmCx4Ug
O5xUkOkhU/BB4nKXIPMJwPOXiJFD5qEFlrFVH7XsjUP511uGcaKI8AfQge+xMMuK
ntvrEzg0lnpKGM2QApAkCRg2gHLNiTSBOsg1nC+p2nCmyLyUhjucZY+au0Ykxnr7
1OVNMR2jJgqloOSpOQ4sD5a1lfaKiO+WYx4Xniygov9UW116yfGW41eHmuOzC8ME
rI0JrokQbLL5EsBNUC3FNHLn9bxFQQRdMyQKf71tccAO38fQJGexVtyI8/kNPyxh
29TVjABTpsu6YAQHaejUakyBmSNLfPJ6n+7udf9X55mCLcMHKJemjUSfnUgCrAgH
i4LWa9alKCIpScE8ohItpDZahYCol4m1Nm4vCUbgJXqYM5q0SRVEDkRZr89BP1nS
X0PVnW06H4SeG6LamseEn4+As5Yn+4afJbtGbm3i7REblsbreyae8bdsrsk7qCht
akccdJj5EYtWNsBdEcSyOoR2W3V8a7Xwplc0afspoPIcK+MPN4eFIkuzqRegm5b0
qaiFZ8a5/edipS2J0JnIjBjqJPKfa6SHyAFKJptLTABtER855eO22Mkq37hywxS/
ZduXwQbP/aZAm5ooeneBS0S5BMGpSH8rig9wCbjEFT1Vbh4iasasY9Yb0zAe1W7B
yqeAEFsgSN9DgOXMAavWx9g8jhi4QZwztr91ONXc2hpKqwAQCWE58vs5Iq8yIB4n
briA+Y0aip1Nw7DX6I9bK+YYYPDnEPphBxc8lMuPr0Cy9HfYLd4iD0BkjqLGtgVu
jij64eUxDApkq8gsA2WS0r2TDSgxloBZeKHkZErf7i8846xm/4rup7Dp66B06pdr
ynWSQYPaLYUnLp0tRruSHjtmillPpTTM8juetzAXhtzk1Q+FcA/x9MF8x1a4d5fC
Yrdgl4apHGgIpXMUB/7SLYPqcnvcwn86iXKqmSUk+SX89GQ25Wq7yUvXVWwRM67m
J2TAqO1rjsp2UnspCkCjga5J7k1akKmjlTDMsGQ3M4IjI55jyMmwoN/xpbhfCLaj
/3nXbfOIijXs/BsXmL1DxxhJNANB/awFYJ93QJsnAJKIH3WphUusP+gV975N085O
lfZDfN3BOSatDxjRhCP8GbuWLR0JcIT+1AxjriZhMRk5XQmHMFXRVndqA6/jFn0+
mNbncSlrYRJzxKIN+cUUFPq24nsB4XJXhrtG5DLkDqVfpjPxeVM4LlVWe7Hs9Qxg
B5YYuv00x6tqQ4Dd+EAgkBtfDxdGDnG4fJC43hvmGxOSjzazassqgUWZLBqH9sS0
21uREShuLxMV/MJcpKXrPUDJ4jlB0+2qUgwZaLZgJAdO3vLBZhE0KDO1GaxgcLBr
ix19ABGeHPwe3rtqRvljjkGfr1lDwx9UJQqGYR9yirMB6I17I2pd1MdpUNYWBaDc
Ca6zIlCH+4q2M+/1jAJ9Uzy96aM3SWwwibPGymHJqirxR4Wb6bWyjTtBe93h4r5J
R8DhAEc/NC8ikTVf44k7OuAx5FptgliSWTfLU0uSH4dFOJWbX+fPxrCU3CB8TvGM
eluDwAW7gTYY4tZrkINF68peTZcR7VR9FbBexDpIRqUHlpbqtWnfocsp9ZmMGdyP
DVki4aMzFeTApJrWA3tfYk5IgdwLprmr+T/NutGZnbmr3gy43tmeT3uZfSOutrqD
JBuapGvm7Y3PX7xDwWP8dKZWvwSglRJ8HXE3O+NUhCmbfL45HFQ752yS1XfYlOAM
UEuZh/tpRMsj4IJnRKf/hGiH9nx0TCZms6vcO0Bk4KJpxc7WRTdoj50T/qHfj876
Pj/1xbGI6M02mV/hC1AJeOF5ryUn/6oPUeVulXhSdzVCTmOtLKIWc6hbL5jZ28W+
jzsk6qDjuy+U5RGwf1Ow51n4c4maxD55mepziZXdMUmCSmi0USaZ/LJDOXi42ht7
Moyy7eSBcDx6kqdkbOuZgDGTozfxBtszER4WFKbQ5RkaUdmAXG+LY1OmoC1yWCbq
v97PstGykLxxmtZlVMuEhr3sx5UIGPrcpTR3wn7VsHpm87eaLAur+uFeXSLZE2Mq
qbRbB4tD+K77WPXt4wRFeEmZSzNQp6dXtHEFaRuhufNKyVCfgAqifozYrjDxywyc
Dh/dY6cOfTb9LEgNiiZyncSkpzAgpjp/Gy4Lq8bfi57tvxuM0bq9x1KaVEzamlFz
iMqV6OU9KKOhNc5tHvOrlhRSCYITXgtBB3Z4IfAvzhOrMo9+wGuWKOERk/hlvhIt
oUDibUK6F/ek7lol84rWSOiMAQ55idfUop9K4Q7bz22OfY6QoqYE+KimYFGoVf8h
J50Q3QJom1hBGlimCzss6TZ64xBANu0CYkGxXaEMkyHr2bVh9pYuOlc1uYjTJNGP
eInVrRqohQj7onSoRWhmfuxtTrCerf+6uuPnpNrwHL+kjuW+/oXf+e4CZkDKFCN3
oSeNydYBS+qQBJOLsb7wavX27tgc5HK8d22h+XCokKDxhiI2MnKe3cD6aL6zPmtc
iVhjGIjERm/a5T5z94W/5OTjL2bcuFgvSwz1yyjbapBlIYML+uVGwZX2yoFI5UZY
5uZWdaPwcM+oLq6IR66K/HrtFakmA9ls5lmw4vSmlLODkbgyN+Tvc6SikgJuuxqc
jwwvHOlRxotgKQ1JLojHKR+tckIcGqGvnpzWZmQOOj7gSxpRlperNU4rge96Bjid
uw5EtsSZF5eJGVimYJ8KYgz81y1KqF3YDwgZWfvtRNcbAMcIWYSNi+iVZ1MWVkBd
EhR39jK+xRXiwkEbosksp1cLIM63R21gGAvSvLDHNYu+Qyuutc+Wazb3Qx19euOS
e1MuGQy1YdrtHXAKQB2yxF1as7emHPqEEpQJ+01GIo/ICFqd1UZ8GDIKJdytO01u
4NgUIK44f3DP8v28vJAycrd8VzP4Z9gPDKBdMVwT7aU1s9SqqK6jeDL3Td0IYj+M
krObF1cHd2EERA/IiPZUxRu/UtN/GNUph6fALKoJBoUTcxU7Eabg5PfHFQueQO6D
sbrcZUp1EnsfsNjBWABjcy7j0ayX9duLpqdcWWrO+CTR3jtsufpHqLs9j7EV1FZg
/qCUrHuFkIpOpE/55V2hrAR49DeUJaJjDBRE3r5D0r/TERyI79tlGWyvxuJh1nMJ
AaqnONUdQz/80XWjPobv2UyO2HziFN5z6w1z5mSt3CXgAOk12v/uJMhCJLy0o4YT
zS8GSfeomp+XC6YkccIkUk6YTKF2RlHU5FspUfuFEO9wRT5u6Lvhtx4my0T5rHtY
Y/pdGn8h9P2EnoSBuV1SmDFo/Fzbylgq/9HkDHCqqwWuFX+fG36/lkKDXIh/Ut98
/SBXn21yl/KLDoEWmEZlot4r5NXNDC21H6WHQ3ci2HPhv7EdlPBdYlE7tp6hQIA4
+k3tWISMMdPjWLIMqHYvAhsyd0cfy+02YdaXIoloTLaHMgBADCjnFx2nagcAroVz
jBM33B9R3aIwTlTdLl+O2ZkLQcDQD1lCK+wwJ8AUT4hCZx2BrkPHvppf7s7ZCtzU
8zkgObnsKPxG5k5qzxkh1Frvnxn1Vnk5p2Gf+A42uhea4d1gWbNiFpaOW54RYlUB
Zd61Me4Ppi1BVYomA2MWAEWEngnAeCrT2y+1x4apGgq1ZxMKsEEh1vrTL8jL7hTT
ZJYoW62HfxCjl2+Qi7JFKeqL5w3aa+KVi7UhkjCrhfQqQNgv6LglD20fv9VEmA66
WFuZJyCEHgSnoE9Yu121/gUFSGAfTVnEIOtKSYPNurLEfEuUV4UCXOwe2BsmnXnn
+mHUuH2UMR0Xt1fvnuBW02ik/OoHp9H4UBAXgVY728FmTTkuWbjZINi/sQNKhvOX
0J0UT38MKNKs8Zd1c8ikLCMKoVm/e7GOWKLzuvdtY0ycnWZ0V/C4navTUieCKCmK
ueBkbNd7l+hjIRWBby194gFEfxdZPoJ5+lwh/TpQu3wRQoUj/+VHck5IjWl/ISW1
E0f5kFnajjU8bemoRL7R35/WuofOwr1Yp6Y9OZSHxrHrKJmeYyC2dZbHl+J4RV5P
6G9rsvbnilV/gBcOfO2a3HjxoqZ9OVjE0mWaE7Gr2UICvSFGB1ABnA8aFySM/LvA
XZ+97lgg01DCzQMYDm9jIS/LVLTzdXMhVL/bzMNJU79ZvNiQ+MPTNUVZ7qWaXrxC
cEKuCFtxovhTQQU2tSVRMNPcHMIMvzObgJ9zfBz8Fp4lEi8sjO9+A9Xshw2s1sBC
szakjQkvxWx3Jgy4MD6TueRzbHeCqP9OUGoLWo+wmWIor4P69lBZ+Xuk6Vx6JgO7
O8pEnQFmt1rTL1GMujwV4NJfgFTRTYqaGOICj//7pJcdwtn0PSd87eyy598Ldsz3
R4GF4MQ/FynioMKZ4lJ8m68Q3PB8/ii+VGE2NOypIEn8OAAVfWXH6Ly+DXti6GDG
qo2u9KtbWM8KsfLiDFzqHmbJ9ednXqvSi5QxonRQlSAQtFYFfS8xMjvnRDdoCa4k
oRJKaMkooWZy4Uhy6dspRo7t22S5qCMW3B4dSJBjtzbYcS01p68pD5pznY6dktT7
c+EYY9a/GKKLa0kOffWoxbVPxCstji19UJvorDLKTQAqORnOD3Mkd9Fmd+lW1GVp
luOJEsZrR4+00pCdfkiUURG67wKVjH8TZYsIBJbEnQh/FVPTNTSXnQGRsKM7NGkG
qlopNnjO69f2koTUwL1Bjt6PmbZhVEq+FW9iFpHrkRPKTMMo5vRYoOQpTx122F9o
qvxoiCx4Bj9aWmZAO6nvUOfUs1X22Zwj/YkWs2IyoJ7CgXjsVfFLEHimnZ7vyv1o
x+QcwcmVaP9TILkuHC1hXy76rKtWSSyQdb8NSCJIwAJ3pyWa5fwcQbXSH3zO1b7u
E/VOZg+lq21Y93ZeSkgZz6Q1I8XI9nmsQdIYL0XVyROZOf496waaXqz7f0JGAaj9
dQBEt5tBfbEVO8HXspyQy7DtEyUCEuUqFEk864KczkJUSgV4KPakYFG22kXGxEmF
/sdFHSN9meE0OpAGy5C6QBKxWnnXdyvbnGklaMs3WZHB7m977f8KuEwb54OCC9xn
Teqfvl+VpB+cpHgyHy44r2tVgtNhjwWEGlDQNPFVs15Q3F6aPP8MKaiSXfXH/yCP
8gYDdh+sv9uDKIP4WOwPewBAJAWWnSLI16pwv3wwSFHmjZxo0IxCwXhK37FAOnUH
51CeX1Ylp6hUK6I87neN7OyN9IcGVzLU/3l2z70bQN4B/kUg5gqXbEIOPxfoQvdd
Y8ZMt8Rf63jTA4FMq9Pvm7ysCKBEMYrqxue8jyMO4OftuFXutR0sDr994mmHBgf5
oCyxEVV3Q0zPmKJNYsfKM/UQVeDXojwBqwc5awDBK+ZfVLH1dXqgfmn1GPmiaju4
vziRT7DF3j7YFccJ7hEbyqocEnHGI3klqytyHYaxtN/UnFribiDXe2cfw0Jhhc4R
IN67XTyWsLk9djEOaeLUZ02a5vJeC37GqMHlkRNBAslsIU2bc+/GiI8/djkrBwgc
nNpjaLXqYFvuoqfrJ4R/Txg+kkj9ZmcewRzEuZywpEcmHv3aBh6Or/H9mzoNkq3c
qXJW0yRPYFNgOyWoXiKMC9R/KUouvuXbvdSuNZyOVX1WoK1u4JnbFTW3fly1xGuM
w2ftC3etZ7+loyP41KumdviFWA4LJjn8QV3yufxFeJENEAdw5XeRSP3ZCImmJcBm
ueIwytoB0+cTMJvE2zQ/t8kI0KMAO+Ky6SlNudgZoRcN78bv0ZV8FWnRMG9YFEcv
2I6UagvJek0+jINljHJRJVH8g0ilFPRrG0akj5rYEFiHYIqrtvGnZS/thNLYaH7v
4EFcJy7wyClh4oZXRD/fmmAg+mF6lnTtFgqGUrF7R6ghxnwxtSY7wYcvYw5h5aLO
0ukRzO8pKzQJca6sRUGjZ2PSre8HSaa3MoLG5y/Bj05cDjVCPDoBEFcwFy8PnN+j
l1l7o8Ta1p6rIcOBuM6L2NapFbmcL+2ODt8eSoNIKjviCTBsOdmbe8f3AOSXbecX
aEs4LNMWDux7enAzpjW5cf6sPVSwrne3mLWt0bDw60T+UaLiosNJNsZ9knY2Oy5n
ioXyuB51YxSMeqYnXm8H4tEUpi4HNxSgN4THfO4cBqfTH5aK6AT7z8ymHpywahnT
9R+7mnWgIFnpfaDH1zbjd/huVWWe+J5S2z6alk6JL2ha8V6x9E7+wtwE6/o85a46
NBqL8s0MxCVTEQUUih43d44HTZ9fFZQJYe/5lfOu7qgoROZnptUcm/Q83tIJsGE6
ocYHHTesfN2YWTEz0VpVp7zevdPPNrVvcnc1om7ZW944iyL4Ly1ZACoAyFKpUIKQ
89Nd+V4wUBZ5OsJDHApkZluZD3hPxQP5w5HplJRWd0g+uL5+qpeF/Qy/HBS615Y0
dwF7vuCu1LDwFtNzS5vxsP3TRHSNSjAgXVFLnJUH/45tTdjAokv4If5F66LhvJX4
3nxnqzKNmWmGk1WEzeWtAlJhe99OaXDkxu4FjFKDjqCluvVFBGlsUi6ZQixH1c/2
VxfEJ9iE9MzZMMG5g53rdvR5vsO8VfDykFkrCJTreJ8QVkQH8y1KuQD0QIFP7jmp
rBmbkQUfIHjj3fgex9TGOwD6ttboR4zfPfjAak3JiHVNhG8kZkdfgxx8+4y2xUbN
fluBClHDCK9KF6f7r9m5Lb/zGAhTM3BHM7ju2f99yOpiG8wYlBCn3HLbN6YdLF9i
iiaTmtzw7uLVbUgr7rjDWLCdXpqplmBSpkkNCV7cEQP9pHEpsSmjl/KXgR2B8ynN
q0OgpCw32KamjcCf4ScWCABOCX04Q8w8ZEP0xVKEfwuRyS4XZA531eZgryCjvYj8
XSvBGE1EBodHSUI+keul89JsMVYQBryl8oZR14+p5KDEvNuDHxgm7yP6Kgoyp3rT
WdPVyw/GY168lsnt8gRi82VOeuEYxQUMhibril9f/pfsBDXfbdNokUiKIrXWVR9+
PwkRGRief36o7JCckaZiFBTRY6rRnmpxDtqUZl8Ak/WJ5f4V2yeyBJkHFUE/lmr2
tj5HDIwyweSktAuoLwXX4Lk308MmSWC22wVwfVVrwdOnn5X4HcnvsNiP52MAAfFG
i0LBbpWScMsajqmg8fDDpijTChpN5qz5Uu5qdF9ujlYqtVB8uCgIUron3TL6B4u2
NbslsquUQRPrD8l4p4jE/Kq5qyhv+x92PRsB34RyPzTenoVBAM+a44WjzxkF9VIu
MJqd75KzPTIt8fj4nZrwmsRWH3WG5jdmp9NPSxUMgGf01gwHZfkrPcowJLBPQFSu
86eVAaFELAT+5tSSULT6O/PLZgkqFlynD1c2NBbnwA2NioUTzwkclvKIWGAjZFF9
7FdKiuWt+x/I7clV9ejyStWagp+N16Nb5k5jPtwklm9JAnRRa3LLwOZFmx+Vxy8l
ryJVMCAmnYxm0emk1B6Prmk38VHD8/umlynwChFVdS9j8EGMd3uduueZnqYN051Q
/2sFIPkNBIpoFWw+PWHWlpR1twGOuva/1lr0uHlrMiFgsO9ikpOYMAC+UEIS/PZK
QL6NYfIuF3wr6ORfyg5zyL4hX1h5kUAOB31VDVgXz5xXWLzq5eI8FL6DazW9zSeZ
Bc8nrQ/AsD2XMTRC8sbaPb4mpPgaN/jO2lODAi7ZTjcxKr5Mv5TxCALl9eth234+
XCLW04I6wjbGFmBOFPUnUtEkW4xn6PWOHjw+8saiJ3T53meBFbILXK0WHfbeTd0l
Q+4CsnN8DyoMWAsIpihrsgVOlTHIm9jqWJWaRzHMSvh7YSKJjM5Pxma8XoIiM+v8
BKTS4GqOyFI+hjZJsCxrUCvBHGr9cjmrD1WVFcGlu/7UCW1SuLg4O+V4GhIMuft8
adD90vwBRa+ANqlDu8iYA45HKzijjzFRuJwB9wabVImjZZ34C8zmFoJMuEq2tOQs
QGI2yhv8XrYQtEdS3HzNhpkeVge6nh9y54BUtLZAIziHuvrIHiuLfR7rxJHyyI7x
hKYea09tZJ5v8fWnn3Q4njopy9KxvXN+KmZGHJqmlngVm5z3lZmDn93T9EpumPyK
NxQI4cXooSOu4/ENbjeyo+rh5FjnVgnGxboC0P8832/dhwjRrrzVvVBxLXhwBIG2
zWhViR+NL5a0/Xt5YoTj6cmojGD++ToyJ7N2MdnA3KsJ0OH254xCpCinKNFap6/E
YINZzfdwgsnHufZgDL/FbC7FDWf47sle+YzdzRmCBabZ6r9LXulth08jt5201FiA
vF9ejx6sExHrv2gQjaGswgO7p5zwddK6lERb/g5a6CAClpHblCJROh5vFpea88vO
YgJv9f9XKx9S1K0kS0yqevAt92HoLh9lnW8SeR43tBeRBYY1Tiww/E0TBw17YWJy
hiMh3wo2R6ESJ4bQX9w2RS/5YQtNFIP+5dJ9XoPQy7ny8qW3RjsAHQkc4TPOvZga
Np76sGE4d/YClnRmr8up5UEc2DAnMJa2lt7OMPOj/wuphwOJPxveCEEzKeHv37zf
rLKyfRmDJj8lKarnWwlXar7F9FWuWhpshBcX9d6Vy8b4XeeX3Ac666IZMHS4Da1H
j88nTUA0paYQk897829KakIbMvrE3cEtnzrAITZpD9bZpoi4mkMEmFD9UjviZ5SY
w5WcP77mpBIo5EZv7XEpJLYVjWOvYarbrzMu7lx2Xv46GQh2tgkL4dQitaO0dKqr
NoxuK1/LLIyeGwHRuCkTRIJlLwF5VMI1WkRuqX2Gkxvnmq3mig0p6QQdrvjVDgT1
3YaQeFQ1YkaiozYlH8QYVllWRAx1ycIiX1rdnjXgKMdOwxeEUACJDaKPrOo4nIKZ
83a19xxFFrds6G01vbxL73FLOgqL7C576495cFpqq1pJvj30tDpqq4iRyYJ1zzaL
i0iaEZ8d2kGHnH+61i3onRzUoxo/AnfJgrpSkI9Xb8OwlRMWv0lqNp2Yms6E0B+E
Z7S/ux38sdQja5RJvxmUXzB4WsQq401MD1TkIhPxiyb44wyUk+hTin9vU+OYUooE
JEm7At25kSYZXHuHrP8bMiV/ghQ+Xlsio+WlK9ajsdWP8KoTK3PCP4J/LhL8m4S1
znf3BBjS1ScQFoPBzYf7/vIV5Q1RMbE65Wxxid1p0kXqax7pDpmAJdAe6ib/mWJs
sJYAxQ7ZHadFRe0fAkbIvrEMSJi7hkaOk+0LqAZSR+c7+RRpStC0vjFlzTb927cv
oIIYdUWkM+AkOn4jSlN6JyiI68hetnUofz5N9RAP6YyqRo1MgwRJwtDEvc0J7Y3B
ulTtTJJ6uSBuSDm3i5LgzG9XyYtIj5tnsiHjJZS8PjCN++NRbpoNT8lJ+NQLx5/H
UBYHz1N3p0ppRfjsv41G7Jl/hNfxbNfNHYRBVgNpmHsXHpeBL2V5aSIPcaUP1KCq
lI9F5uDOmTyqVMn6OQLNCOhx4PAJ+g3ZOOfDrEzbAIfpi2jA7N3jSbZyxH49NHeH
G5h1fiV3zPjPBQEr+ftDT/E5aBh+HGJUQqdlObb1nOvAHeuZwUAa4DXwfrlh1JQP
bBJLUzhTPFNaJA2u6VTrNY+2YxmUDgW3yyJ3gqQmjdyfC/QGE+b2o36wJGU+yliV
LCFAfSmP117SLeFr7wxyvTAnAhEs890qsLsW65jtoUMvs0pJhc/UMG4nFMQAty0z
LDRua6PTtxDgp37OMCsv3OAaWmE7xWppBmWC+bxFB5G+yXFYEe3Cr2YWoLTks1WF
AToqDS6fSgLL2xgSP4ltlTJegqW9cbJhgG+01Zz17KSrPhzKs+u6oXmhJOnwtj0S
PDRz91SJ/aJwG5ObebZkirkdPbnopJRsLypllaMw2lYaaXamDhq9rFs9z/wBINLD
jMg/SePuIZN3NPVZUu0UV8rBmnP+9MhJ+oOF88Y/F2SF2sjjP2lgrQzEfntss/JX
jVBO8FYw1IAi/UlEKvaxTOCX2THjhq0Z5aMx7O+/4TFbYaFUdW9oSX9xtuEzKJyy
Q/zH19t6Wb00lBUagm0UuPLFIUk8GAHH/63ReSt8pIHJ9oNtdOUHTiAyT0RkMwZ9
uEs2ByypMPkJKikQak8J8rWyl8LOFoQM/D9fL61STG89nT6viyes2yD6AoZrkmMg
TuUCRSfvWixcdQBbin8/xCChJ5B03OWjtF0qsEhZAuGwsGdzyf0CyuQIp9InFB+6
Vc7QP1rYYGWC0OrcmNlazRwhSIsiJLd2HFXukG9XoAgkM+Of6q/KyCF/YQwGw+fx
eiDZAIuSVONVYkJzhNrVpEY0dIMnV6BoBPhRnysN61x2mEdTKHGRWwHniVa2vbDL
TslMY4j8zrQfx3alhaO/aZeLwG2l6xaN+ZLc0yKG832Ondrn5c+9S6ttFH02HYlp
Cgk+UiD18iJRexig/EXl/TI5H/GdKb5Trjg2x4do9xssqZvLoiEIe7r5Gt9o9yr6
SFa19t0bblI/H1pyZNKd5+V2toj3Nm5chFUgcf7wr3NWKfH9PFrHuKOze2SDqfRf
oo/NBFsUd81TOu6hXWRfNbFoEucUkJ2RblBs9DbtQTc0FZkBVbm72zee4pgWpXzJ
CogAR99I2enEzNJtJFOZ1ikB6TFJADr+3qQ1KMB9Vcwg0umRn5/KmlDO6KqdANP6
L2PAS3/7Gf7fgpKdEtjGye8oYwG3N6GBOf9nzijqqq1UU0FNKHOUdDAbMoGj/738
IHqf9qZkPXruXbzkdSVS/pt6zZe5JsTDOBFaU0hm6wX5ugVny0iYt9l8NKctAPCf
Njac4y3AFX0RONk8mZr/lxjlVjqpziZmwJtAaaeXkX9SFAUXzPSGD3pm3ieX0yAB
hFZupNSi51K5BobzB2aD1UgkO56JbwjfvqbmIE/CizIY6YcIxlD/idQYsKJXc8V8
OzFgCx3sz14doKqCHt/ndWw5He5Qoej5Cfi/8x+m78Vbc+UprscBtNm+1Wox4DUn
eggAn78mIhIQMj0gs+btBu6NLnOSfrv/FgOcuwiNceGUdeiimkq31EFOXDRDcIDQ
9S/49oY7uElTbWegmFgqWpm89co7fLw2M2fWo6WguYiZ5XbG6bkOiPZZGpmaZmUT
jzjrkoYNg6i4giQjHUsIhh9Rv3cB+HYXV+W+/8/xSAuQmCQhNuGBYQwCCPJt+ycy
eJXWJg24PeoBB7RFrKPt5jt+WuFt5yy7L5PqGbblQGmlUrDvHdh/8xvy5hPro3Db
Rj9RdJfwaLcbNx+gqWiPlIJZ8UxABzuBc7POi2axDuCnKUbt2H3InzcX59YF0fip
Ezmg32lPRhwoPl89kVAcXrA3d2kKxlpv37/1fKMH7WgBTVHEgOFun1yX7cRHJv9f
6f38QlgCNL/3rsr1pNYqO1ZrVmNEs7qYnW+PcOVhhOV6RJmRO7hoLoHmCV5wZJ11
2jOWJfgxMyrk2OGDhdtb6DTfjQ7H3dBi7CRTTEW6O+MdCha4dMjyp2SnfWsi6Wle
wpXK1m3q4R6lT+drAX64txK+L1GIZXABEjwaC5BF0SMA8ErrJUaDCiKyiKVYucn0
A7r8ZDPb6Zi3ptcIBVlBquhX++rkK3yiwlQtJDPOH1xgu24pqDFIxk4gkqsrON0B
wbz082SMQQE5eUAvd20bk0iEh8NUKCCb9OYOZS7hNL0DvwU2JrSFNMFk7zfSCPzK
l0iY2FSZ2W+Rg6Vc1tiZIC/gEjMoOVA4IptD/cvUPmyj++MvO8yZCEGjK7wbmYbG
h38doa0yES5RoZT2xlzu8WRdCvWjNeXUcWdwfc8gFGM+lOzSGUSfstf9LYsLqhwj
+kO4b0q5QDgJa/9xog6PmJnXokSJm33QsnOi/AtnSzOJnPec0VlqclOQ32CW2QbZ
XOVcggAXZV1UFq+vLftamr6gt29xLeah5waj6v/lUAJc6UBTECD3LaR30TktO25s
KrWQIaIrvsNWXQuHhE06/2kJC+erYMF6KIlGz8Je0HPTv3VuX3seUgCiUhQdrX28
Poy6LWieNwXdLl/Dl0BchUiFcBAibs72EQ7XhdrUsgL0G3CpxjT6iUDsNRvmxZfv
lbioH10xPGOo34Q3EWuJg4t5vZ1KzCK7DJ+UB6i9lEODGwXKN+yAd58KHifDCu0B
8j1fpuZ3klgYkN9kWh82x3n/YDnl4ZiEhJJHHP6XkR/Nd+zteplXQiJcYCCm+9rG
PHAhU82y+LFDAFe18Zi6nJuU+1FUPgthVC4Ry2MbL/dyCAhMpiccmxf3ySQyGHsG
PjzjyQtx7P4uyBJIBKvU7w0x/r1/dawvKyZ0rlvah0CF/sMSmPxuoCM8qGxqFJy0
zew5Z82qADN1xxtp/yxdsASAts3wLTwtOwLs0VnwnLR43KsgqNOhjXJRqvRxq+xa
jNsNF0uqoQPz5uA2tOJCVMBaDe0DZc8e9LB3dY/voWfl/3/9YSjz8JkmhJIeNg1F
onkOW4SY/5Tc6GM03Qn/Xcwmf3FjM0pFdRC7IS60zq44NZY2TtAYvs+rOXIGmT4J
Ok2SczE4jSc0A7CYLX9aItWhj+YMA/e42bXEw9ydS+cygLQxt8Pg/oMyJgoQE0mc
0aEVpYHWjHnmkos1E4ZP/fhyYbkOVFoEPrdTVQUfYn1adTHD1c9jGutQtg8MbHdl
84j3snBL6649D9FGrUpO9+JPdvkOuAJdjXyGfoxRxdglAhq7GI/6iJ3ynmqrTSMq
9sAMtL1SJL3mC7xugplKBhW8BjLP03LFLgzTK4n2JTw9eVE/0RxPCyDxaeJzuWkY
3tJ70hhe+USRsZYCKN0VhoM9eKvbFWwwicQN1QfaAnp7T+LoYOM/PV9wDEe5tr1/
8GMYmnt2CArDUB/+9nK6lgjv1Bzv6HFxrN2CDqXyEDMnNWGwLpLLj2hHqUy4Mek9
IO8j0IQXt/0P/VXyY4EDCy+mW3fHNVCCuw0i6c3C6jiO9vNzSz3ztS8aZgdW9fIW
C6GBZFx0e56/YUzJuUsxxUyNZLwaWQU2cXaNXTmM4XhfhQB3aDMoManF8xH5JWhU
MBksL/1y+W8iI2jsWKHtvS5VUqidYlT0kzPrWeOE3sah/7QAYvnMq5DqqobrPdzT
yocTr/1rWMvmiVM2CjA6LnkzzwgwD5sve5olfTD6cLq42cM5LaCfarkFkUNhpOBI
Rtv+BBtnfQFd5N1plTIOVhAzWVO7VEy3VvzW/DF8FfcGMHXUojHie9qaUJsjTuFN
TUR9/I+X86oVpJCUSr7gwVgSeaCcOvdJYLDqcbeUCbFgW6pLPD1of4x9crfjwxMD
/1xsSMPwRwsmHobmoUPnmr9sMEYlgq/00cWGpDKLjTdlytu9FxCrAIWI/fVUM2o2
ndKul7Y3qYEPolepfP+R+ZBhN18jIGyOyshCknD1YkmTkCHZ11wWDXIVjWurBkaN
A0P9zBZyLjyLhcNtUJNVVyFBuMJV98kOLdCMJzZs3hr1Dybegjz9G8Q9pYkFsdnN
07s7lVAzxbyW3WvrDp+WuvZ9UrhEt6ftvTZfqxS7MAvPt0uWLrebN3VVaJg1B2lH
g3YJ4w3kZf5Uoubl3iFvu6PNZQwzEOdoS6WvfO64qmEIkG64O9zVAyJZljcQ9m3y
uHo7l6Z3Wy4IH1RSTNAqHgR74yO5fWujTkQLG8t++ppXotDRZb2TmyT4nzdf5cPt
nJ2Nky1FFA1ktzoDN4Dfp32IyxiJnceHC8ulp0vBVk0r2q1IBZckd+I56yQjGBzk
tXQiiX6Ho7ctuebE3UZGbIfZUR2XP6JBHuwfAsKZy+PRuB2w0RGwXIag/HIWL7Ie
SsaMOYuKlsrzZgRWHDAPMSdElLWfKzSdxJs2P/Y9yz48QdJFoCTJcQlKPvKUkdM3
2W/wFF3P7qRcAnseJmD1T9g7ess/K4/LLMxlKxblUORJ2OR8QUlDJZFEDeAW3v5g
1+ilYGh5ppHyCgAPgP3N/sW107i/bBn78GN6Q3ELHPqHehGnuF0HaPve8U0IZJS3
emZdbc317UcU9r6r/JLYIib4BIXC8EwssBJpkGSl954Chw95Z9rMC0GY3nAyVYLR
E7rNtK/OGPPkXo1oSeUgLDbEJh7n0hlI7N449HKFhzCEJ9yZw+yPhqcyfDHk9V/2
8d26oIqjVhNM/PDkWsj/FB0fa1jsar7Kg5s5C7u1vk0/5z6EuD6kwON8KDYFf6pl
n7QdLuVNgXw+F3OV6FHrkdka+o8nHtQv3YUB1ArdlotEXUkBY+vAy5o/JCiRFZc6
afvxKBSGCIFeseCiBAtJ9D4GGByDqBW+m3su29vONlHWLs4pEhIWdjZPF+QoKSU2
NiRnlwHeDG3xKr1CyoZUcaIYhCT4pnnHh5Yn/5uqLadxrSxdUNjZn1kemXYrZRaV
Gh992C2LlhCIMON8BzZSJ6Zhsl94PEM/AlvrYKmUtW31/jRYqJWySyJOYVQ370dg
iiulK+X8b48+yXjJQQC1WRrBrPkMW5JmcErP/T8GO/KUWsEtli/aZbTE8nPv+RF2
d2p/GaQRhhzuoucW5eDRdVYDTWIVjlGK7jCvahtV1wQKELr22QPn7GD4I8uTAD/v
c6CCCpFE2R1kgppOtuvtFeZutR+pdJEyV41sSqz/lFeRdYKccokoEWrichvLvSyb
8Pjpq2S/mc6Ial4uD7AV6klgQ0Q6oG2WerdPF7PuVlbHU1VOlAfLfHarZOsVj1JQ
yFML9mvB6MWuD2AGhA31nmGvBwsLt3Tcj4lb5UAbDIiXv+Mj1B9SY3KcIf8citdz
ZKRzgzsm1JhXe7fvmhOPdGT25v1SOwbITTQLX6N/cxqBI90WwGQRdUbWtqH3zE8K
pZ4cbd3jd7VkOyUI1AZLhdFGTabzx/Aei85f9GPxjNLLcSSHnsSBnmX/D9LUpONX
ubIDXcI8o5x4nnQ3vRVidCMqGXkUn/gvNJqxtzCpfJdennoVaD5raQFH97iZijNI
7Pf2EvpIHsJgzLTMPKUAYHAThooZJs5J185JdMDDaaBHYR0uwyDv77o8ZxTQSjM+
6t2+2MhPY1cKSw6TKkklCqHNaYxD1NXzYxBdJi29I8JBQv8u4R//4BmsOKKhHIbA
HIb9LUve9piCmooM/VgrumtojRS+TMJP22N1AcniYIK8lJoto1NQINPlltUwf7Vv
206HZwcpdxbFJc5oFFQndAAsvsDyvic7DQS4JatJ0Rsw3yGkLLkfkIlVqm6ysB/2
ZnXjTVH9Sx8hDzxoIsVxeiQUzAYdVQcOjz+DfzJg1HizKHUKANf/2aXqzat+S1AP
dtiptNMzeCsfyDPe3aJQbhhgEMAUDklO0wi+R7EQN6YE9Yl2zzCoAmdeGYyCHMv2
qh9iWbBJSONYL6UGINC3PgRx5hf89778gfZsnU/NqJBnuanA+yY7MQXF+ViQ/8M7
Va+n/OjUpHnKe9Xi2r029/vSTLAFfJZ2YQIaNasmA+JzFKyrQk07tflMno+t9sDm
TfSP0Bk5viS46+qh8VS9dYW9b7pOlPPfuIaj3QHb6K9jPXwDiswmPEAoaEWrP7/+
5qsFPelz3TEPaTLolImJcUfU/HAb5lR6af/vD5O97xy8N2lsroLdxPbStEweFDWK
EKLp7y31A/1J6BzeZrS8Jf7pPFeJZdddkJWwID1ELDpNosP9Ft9UlaK9IUNf8MGe
VSJjvifrGhu4X6OOpLcC4R/uIObu2ImWp4xe9KKzLXP1YrCWlOU8HRhhqVf4bawn
e8vngOp93bu3Rpy3NaZb8gYoFDYwmqE2OdTdzBUZUc5WGvnlEFOZw9wJxh0uKnAU
v0Fe5DG76UAuF1Evzv/KR3gr8Gp4OIORBA9sxrvnU9l6Us+3iK5o6LINHSHQl/fv
NZFFjgrmFjzQqOy46OBtrOcryP6pmimEgGvMEaUHa+pzPFyyarJ/hoZvpqwrvoGm
/WLV1ndSRm4c4+GO9dxvqYDeJw619kUr6cpJzuswoOApIoiDpzRc1Gl+sbBY/CFL
kAY8uFo6trZo9XouFGo6k9Xg3KOQ6vs0U8LHz/yAb/qpYwQRx/oOs8KnFUoL8FNs
/IYx7ZVcMiRLngt104Jcvaj51rxcVL5wtH6ICJIWpI/fA0fCaT+etc7NQFi6TTtM
kdPD8QPuCGMkdTjjH9Yx02EvyxeEKwhGLSq4MDjVvbzz0c8BzORT3CeEp32tOL/w
ok7xNK84yT2zTwEkmfXxiDj/Js3Pwd6eSX18CLqHimYz11yWBVb2k8NjVfBgayG1
N85hMWV0IrcPJ5J2QGYjIgENdjnduQzjPVcqSMH9giI5sdiTsrrz1ilOS3pT71FB
8EPYj4fcZ4Q1GHloEhMyx/M11CUUFEyyrOMw0BVXaJ5QQlzrJvsapycr63wV6rIU
K7h+7kCu6X7g4x16CdEy10nBKKSYiv0mQE3YHnyHcW7b1gG2Mfl8hwPECwO1VNGA
9Vd7H3+zpy+3Ps7k9/ePkqSt235e8iy7SuzPjY4r/pjKnd4+vh8T2QeyzpF9Dnio
dFDasbxZC6M6EpeiMLjI60GQeNArBKRbztcpu4+c6fZnNaotnxD7Bj9lo//QJZFw
+W5wLkn3aWVFNzXhbC3ZkWQCv4sXsHTu26zl8FCf8lug6qU4WCUbk4s4qIxpWdpN
1wvHG2QtCGjN5pQ2Z3Bs3XJVi80Hxs7G2pUdpOz0AMwEewlE5LK/iEUzq65MxEb9
eGT/tfHHY1YOA0NXrW4Qb2mMBufKfFxLKftDPsFHJrUvIGmfvtzDk7GYb0pJa3OV
35zoEKbMQ88bTKgaJioZwIPdkVbO6vSSIMPtxmoZBMOyRyoYuhPLvQWoXd/i64Lz
yCfTA253kgHiBCf5VXCsICiIx44D2ATX7R3aRyCicDQftd0h0D2B2YVIEj3vijuU
UXXsxqvry4Zk0CATk1po1TdZSJkz2rSC4PbMZM8BG1dXy+8yC4zYf7B5usDdDoXZ
Yz5czdSk/CdDnhWyW+TDfAotcrHXmd4ysL1ZrViLzH92Pk1BA+qFglDK4+eHU55V
qbJkUFGvFvfKwo2BpTAktUDjr8Js5zV0OsXGh39oQwFQduCv4zo0vxLK9pLEWv8z
VGLRRdrB2KWVjZQCMwGJHo/i8DtAiTU8P6ovbq8PXaFvFkmcKO9tBCKcnUXCnZfV
hc+xd750d7egf7peXmcYEVuwULERvEPD6t6qYfnjKZdnXcrvBa7jxgzDk0NKexEq
Oc2ViDIR9YQhKPv5QRqz1C4DvafIun6Ni4jnUoFaiw40llfbUQcb8v+djAKFxUlE
S2moB7pMr8MYZpyp4LmpGTQanigIcQ9QwEuDu3FrZ8i0Mg0WpvYAGKle3lbrDdo2
qnLLftevaF9xaZ3wR+paXgS1bDBeQRAhTCVC1fyj4/r9OK2voeHo4jbkIg8mq5bB
pR02ar8Fuo6d31d/lp09jD5tGg2PsGMwXyXqjLrqoC6JwOUvJde/3c7cW/f4fBGk
iEtah/BAk6vKPxrDIlvpQwSyI9eJ5ZGGZdDFbaLqKpouAnllgZEQcPX9BR2VfbNt
X6HwoHQoAflKi0HZHuoSg75WsDgq9iZE9Fs8S/Iw5tvMsTuy51nDtlRnM5FqzSus
8UFa94m68VwUk2Md5frMWswssh0K6JhSNqCKQ1oWP6uqrqAOv86c9ldOL2UUVTA8
cqlx06EX/qngwyEqSqbYpdPMmV8SHj6GK8zbbxuLMz9S1ewSnfMcRlBHYJ4hZQYa
f7bFxoHf9IDu8EPm9u5sAO14VL+xtn0HGO9XVbKoiIwlDi8oMPBVTqFLbETcbCiX
PvlSpqwc9wBlflA3gCJWxQs8J3Cq8NFE4bpnRs3OaF4iqameGt5aK5ZmqcAObUG5
lZUJ0ZwM1cmdyNqufCYCOBE04kwbq5ypplIq/cd9LZfAAJoVTVEvP8JLn3Cfes94
Kl5aOWMn5MnLZQjhGm9fgvqrAaQM476r3fWJSh3PX1YUJeXRHX+3fZCMLyr9anRL
cu8Nr8KIgz1xScb5HNtPIj3k5UPUHsBQ4U9PendbMd5AexgYvZ4foYkyOPsDB7++
56PO2kmKY13svBAwMe8hcAvg8uNUHArll0ukS9liKn7kxsFcjmAFCN79PlbtjVnY
PWT1IDB1qgbZJTukH+oob/vAT7uoBH2S0O/FanOXQvDPHZaYS+ZwpRLL43qBqnjt
SqCpYpSaL2QA7YXASDfj+O8+N07gQTxp80SvfwAOoNU8fScbIrKn/PUOpAdCOKYy
qWHxk5oS6hCRbj8QElpeXVN4JkBY1D7AcBBG+KTJKqdpMjF79Pfbhg+mOf4NP4vC
Y6WBZdFGxA47zkEhaMQ0aHOoPWgkXfeIV1R0kIZt2/eq+LhNcZWbAPHuoRIiAuyE
6PkgwNfFEdi6g01zkNTExg11ou8O8wE7Dao1T2L6jvDSgLjZt3Qj1cAQOJZZGHPu
sfgxEdMMOJtEMK0NQH3Sb0hIFcV1HEOAxnExWn6uhYRmZWj5tAuxVFOdGs+EN7T4
AUYc715jopIXM3f8EKTUsCbiD+C8DwKi8rRygOMxg/Mr8RGxOSJeQcHIGXy0pNYy
li9RiSqZBweZ1bJoaJXD82SBxJ10HzGw1IOnTr1oXHzRZZkqQm0FyarHYBxqEvNd
D5SlWQPLimK83LU3uFFQu2bJY8KOB1SoaFwgTMa3H3cWGJsWwuMOPA3xDsm9LqpT
l/03EzFx0ndFHX2w01x4AH6kD3NOy4KlXyVMrFEiZe3nZ/UFX6hC6JH4fE/eMeZb
i6vcr96ehJU5Yn0F65dxg6/SY80svI1EpEyuZyqyd6rNkvHwAUkqYWLMZO7jIVSR
1WJQUFKoQeeP07E6txzwuwW5iu0E9xz0tKHjpxwpPs0b+gSk1Q830bnM6rm+blg4
/CaUMSUgl99tOSIl/WdL5QDMq/5b/pVgvDGJtIO6i0khNod9031AW0XdKOXWtA7Q
rNskJCO0JL4bPRr0oEAtvj7tjN2Qjx0TVFAxW0NkyDY1hpoClwUd0sAmpBt7y6mj
MSMrKHNg2gjVV3N7y0NHpQIU5KFyU5Z0AXFjbKqKCVNe+TH3fIJIvhD/WWsajqLA
/iyIZmYjfeZCyySpa6+Gx8l6TtsAgB2r5ckQaQYHIFc1PXTvwA6mf4DJZVZXQgXh
ypATDdmJxZLKYlsOBle3QK9Ne2hQ3VGsxkGf6kSVkqoZAWNy8/eyt3fwGIuUSIef
nPsCa+5xBw1MTLPupi6sZZIBFbD5Fh6WSHEiujrDTdNhZOb+AgyWU0d8hdwwBA5I
iFtf/HrqlUJ454467JBvgvTuAnglgZvfc4uqMf/UVsGWJ+UlTEzwPywUCHOL0qwB
1ifiZXuLkx448RhoW1EPs/wNzGKHjyhrCTMsb2FoxAzYkwSJkOqAT0Zni5CiufLl
4FY/AklWoWcdQPVOOqW+r0UrabrNO48t9GSzZqHlFDX655FzIy5p9dZwJn3Notcc
1LbRsduWWRzhtX90+DDsiXImrA/K/1WHH71iNq5uwdyJfpcrDOPooedvgB5bm8WA
mWGztLXo4VnwLskFpBWY7476Q9/kM54gxpyRxj2VQxilkI/BQZ8DQLuuTEmbiwb5
E43xetdY9Rv9UsRlsApukI9L5mBgTPtCxQbA7Q5rQyuMDKhOWh0turi6TXFZWw+V
L9iJ0Ix4A9Ut/3lkgXHVBxp439igkx9+3nVy9SgdcbM/eMmkzI+xqsG4ICoYGq3b
3qtNh5aUkdeWIw4X7oBJREvCqlK0malFO5GhQNGN3QtguwNc26E6C8oV+WPnc/Vd
HunYXEdCk+O0TZZL/tRSf81jmgWqW2W3oAsenEwPg+DnUsTQm2htNNhwq4ns7Nc/
1MC324d9WfuuqRekIOrv++p6g68rYGKMrNUwVBWYC8haWpaUT312xEkgjscVPBxn
/D7dFKoLTZlkGVa3j+wuFxEPt8ai7zwGeC6bMPLLVqbw8VbQ1HGQIwimUXG5lSLm
ckwxx2cDLCldENbKB7bH+QE0K6a2OVRNSeTHLDI8QEgGSOrTmV2BmY5LFMgwtnPE
+bf42k75rzznMPeHuRtDuuTo5rAR7Ct2CzyOqT+M7p3llwd99JfGsMJf3AayWnuq
BZa5Kb+/FE05WxVfp7GD0Y5jUct2EJwEWDrO95RZP+2DsKRyr6iTms9CfB7hab0n
bhjUnO2d3Ew3d1Yb6UrZIspoi4ab4yzUFVKogTbskMlbDEu8RjoS2MBi4NbdwAM5
hSFCGkWUl1rVIjjolr4JCbMMdD4Jw7KE7tnNMZ+Kr7q6gtSlid9hojkAcby7Ws5w
l5zGu+bbVWy9pd1rzaoL5lbOkRcZqhTGaWGFBhFa8x7rHkmDKC9DtBuj3ZEF69Pb
U3v3GpI8fElS2hraLdslqHLsHBIBrT+r5+PyP3BPAs6H1W2YJfEGOlhCPuskZ21S
3srTnZ0HKMv+tP6X7FlT57TCznn+iREKflfcsaRt2TzhF9nEWh50jl42FW3gzyOI
ADuvP5snN4jYGl15Iux4oA7gYX7/vSyFqdlrdea9q5mQncCXa4BFYL/7f1YBk39J
hIAlvq7keHY3ECEY86gyIxgE3CnHBCjuqIkbF0i2AcsyRUyCsO7SIK8B5kprJk+T
WDh1GKccq3S/i5LQ9MpV49Ic9GUmZAqG/Eso0EFUTOYdipcNoE9dKOYZ2dM4RF7v
0ZqYBOaSoa9iI+KWg2VNdt5cpP7GyRLU1u+3OAT0FB7keugOEFncZzB6809Xq0sr
L249F1d9X1huMj6ge4lQIRhj+PxZoggQZltTaJnxIiKjSz2kKVbJSXYj54dS8qBs
xMa1sHJ5niystjp2M0rycmxv9r7beqis3axIIrB/OVyyiLbEqIGoLwgQNxNy6+aW
Y3MYRuCdGhzG2eXdyPLIKWEvIu9ig/Fd4kNSyGy6wLUP2s7VXilD1pdbDhr6Bt/4
V4EFyXxLuZFBaKtADRoQdfRCA4figyLKjRqAFbBflrSSIElv+OQC3BsNs6/pJ3dO
69vf44/eTDAtdaloJN/qGjqV96n9C7BXRxRMxgzLNj9yfboH3uPbJe9hzGr/IY3o
NLHwa3fWHokG3VIrRwD6Z+1Qbjakx+Qg6nM3c8BtqWRjiPAXeIuOsunFSb5MZxmz
5o0nPhTaLXsJU9GLHU9ehZOYZgCa62bSrHNVr5GMyKRj8eUJrD8Wu+x2LSgbG9yA
eJuxyzSPbZfywd7IGX07/N+OdOcIzYFamlLuCSOb5bv1nnLEJ3ilwPTm/3HkfP+p
UOFg9cQYWQ/NByHiC5ur9W1iHAoWU8XhIwdfrnetiCMVjXLIj7QCkzlTbMT/M06P
NAChfcytr/M4F9pO0NqMBcquA6G2AW4rFXaLTMatd2bJjSfPglpT2OVznujn1q0J
v6yn6UbpVJ2epn4fHMlBWad6HjOZJmXAGMgZdg19palu2tU563JaPGxON75CCa8T
acFt2clU2wGmosvmfKgkeQPzMNghyPh2ijyso/aUaa9CCPztP3o9K+HAQeSV2I8L
rV93frE2dI/cPomgw1XJSOxHMrk8AlVKMoiUpuXwGnTLJ/Cr+qksWY4WS28O+LII
qzHiqcjXumjalimVyU80gouHcRABzv3K/cnP4KISL4ElRYEX7vrLgBl9R57AGj1M
CV3MJzWL2H5J30DpDRczb/tCNd6q019m8seWOKCysowXake2ssNN8Roil/5MSOZM
AC/ioXsBwGf7ZuULoM9/yZqBhJQNMlNU3Gp1xOsrFhpVTx1MHw3HT4rn01IKNPCj
4ZWEPRaUChWVMbvDeEEM86B1wquMe++/MQXvXjZ3BYWHfZucYJJN9/2IKurdhn9v
CqcwKSs3puDMC9zvGVZjiy8MB8yXlED3X9b4+kVlT8l0nCPISPTdKEohh7cW/X1v
QmnCLaTULo+3nEoChkbiDIdqiVq5nb/YljKuX8cBGe5cNgqSd/QaMQuLgPRvGeyF
mNE36bocZQ4DBAWF4RYplAJTCK+72aTF3L9I7u8pyZ9pXAbKtSKH0ST3c552WNoB
hyuza4t9BWY8UTOvI2ubaEhcOzEVpyErsWzRe5zHbEy1vwAfQSCua/nmn28azWpP
T4Vyhq+BVvBRPwM5fLlT8l7iY5sKXfhE7OacOVdjOxYwinNJoblvdZlKXvj6tdYG
dNbnaxM4hJvfe0FsBf5O0bwx7I4veqEIDY67a/6pZ4MeRvRI8QuBIS1T8Hv3zJed
Asefammv0O2kASU40nSKrmdyzVzIr/VSzZDWVHNkhjPeeR/L0tasPuFEDY2TLRwQ
9PEJHhDf0U6P06Q2Bs637Z9k2jWa6MVRe7WCqJFBbQFVGrSRpRNdiWa9xM3prBxv
9BeFHUkwYbJ5Vfq8VXxThJa1EM2FZBMAvwAP210o+0OSUve1L9pSyFcdWX7FVXxJ
iTTvZSkUMjr29vI/Ft7AcrBxlPl2JYjyFCXpNdrvdLWkkeTt2Tbh1u0kujfDxT8k
bgC70fws+FptrjNcN66YHyTD7xGUVDPeK72T5fE2T2td0DUBVPARJWA4QFP/MXjm
+TGWSSD7i0md5ZAyiJGYG9snnCbGYT2OLJMh4IKyuSMM0GOxg5RCdZAXG4BeZpxx
V/u5RPGv/vN39NQRyN+ac1jXlF7gxc6d8ZHRbGZVQb2EnO9e4nbc6IaQ5GoynAd9
+y1D5pU8Q9hccZ3swExd14bLLTeC8qlgXi8bKqgmC/JrQ7Bm7QK5YHDnDDfMmZuW
bvJU7QipUqAo1uxtU81FMkw2BlRqVE5ji6J6yccC8DvVpxZjBmIrkQnaj1UnuH16
LjLYZNTlW21JQcAJEzKMq4OtC6joBCCwPosT825+wOQWaj0eGiG+uk5oqNvYZDNF
WQJtuI0q0sHSp9r2hpK51R+vRk2M4apDmc5pM8imaPQoGCanDMOub7zzEYnpWSg5
tFCcOt0O983sjqMofkHKkfk8TKwvYuj6NypP9QCJa7M1OjQrH9SiNc8DADqC7scs
8/KrPIBwSdKyc8Qiv4QDotXadF9tbtlcy8Di4DqZEju6qn2KT/YxdFK9JepKw4fY
k8sSnTMe443DW6qLYltXe+EhqQljaR8MbkYx+uZtboTnrV6KbIGjjcN2Kri7NR+H
8m4i5R18O3tGYYv0cGK0k50WDnT27Tq4eimvEhgqJMCBFOYvlk6BFirUy4AXt13h
AWSX9B7I7LL3whIZMz4PHAJKye1dUdBGnvTt3Cg7lXsvDyjDmiKdMBuzNhn+3VTj
DwTq8RPJtwBOehml4dxEaKYQ66Gqoa6zyLJZyS2orlXsh4osch14b+O/zdjRpC0b
UaDnjtvKoScqnLOXnVeIfw5bZ6zMFWsmOJHCBIwSCqUJuk9CRrWgUSIQbwYjvude
I/U/rxxb/ZVLaMdwus0WU+PgHK59p/T3hmgr6lmcZdN2WF4xUHZmlHKDnwJ4O5Wu
CFbcxQReAl+OxYb/rA32hxcVN/Af09zTX+NUlpb4zj5nrPFSFGuC9eqEKb3INJ0s
8cHzxPzpJFEKAg322W+guahEFI73rTnQ0JNKM1fVjunilo5d2cexsGNJAaXvzMB8
PyT2KeFi3aLdxwrCJzElNaYmoHydbRegju1/LE0u/PonRioOSdUtqnTMqnpuy6EQ
5eZh7DsYPjrfRyYpTRMhAMagWi9OVY5E1+3WciWRmwtIrMKE/3V+7gaTqcPDw0BZ
RNBl7BtwqIMTmqi6nb/u0L7ZZt5LGQFP5iHSVSQfiGNsmPtc8O8iJCvL3bDEuEoE
WtDfbrGp3jZVb4rSNai0/sDY1Sjbgc23xXRdShW+IJL0tmRDiXli0PbLJro5oiRX
xctfWY660dzsYdO9LP8FdNZ8sLNJckHNzHoAOWVtWCbMc8Kqe9AUUxVzmz9d9uST
yWUxQoiA+a1xfuKEWgz9glf3IXNfjv9w9HCL0PDglkzAWP33c3tWscNA6Y+7di2Z
HAoJBlE4iJDVlrLdKT1rcu3zeuk+q3syvMEKSI/+NnuHBefJqKlvWyl87ntmIp7c
lsrrBOouNLq14KCq1CgV6G7w8KKqzBMQU3YNc189F192ooV2hgxypHlxpYxHRwlU
lzl906SBIS3LJ47GjCMT3VBtArOi6OcAFZP6XBMumv1VrPe/MDhKHAYJPX/5OSut
dUvXnOLTjV9FSIundNOY8Bayfq1s3fnmnJapB7eKAi1GLXs0oY/YLXARcxxr9WDZ
yd1n9im2bXJXKPuhYgXYXsq1WiTB3+Bf92+Yg3EJHQ+aeBKlcgVOH2KMbR5htCUs
uZ2XoahyCxKTn/wjuTbiEOVo6fqkbzsCjeDdyeM+FJDK3Xf547yRtGRs8jARZJCq
KiZe45m41eruz+XVBpx2gP7FePQMbQHGJgVVF3p+R8E65m4VsSM8XZXVrVqf2kk6
zrz94CRI0mQJGTXnnpOAFnqsxXUV63laTZgnEyv1of37x05HHxYIt6MJnaJOhg/n
C/gDJ+a8mdgUWgMIhI/sma1LjZtrBUdwhAmD4IWC1xI/+uUfKMEN27JSBu2XR8P3
JSjEw7ij0wsA3xY7jIZXpNxGGgRZU4qRNLI5Clbs4PfvB1TZ7aeaimuyg31z21eD
SNkEyKXLS5kGwljae2L+0lmZkXPcQtGKhds6Tc8+EGXmjDh5eYzJas2El2XLkhBP
zeueMuOfeIwlF4/jVtH/UJSmFFL+UabqciZ4xwefpAWbQQ1zYM0qzEPtNpaiovcT
ftsAO+rUp4Jl4kWM2FSDBIYdRkYP7ve9X/nrS94ZiX+cpAcdnAdCD771pZGb73e6
Lv67EeVZQhdkhZU62xVn+3b8uPtTCH24af6iwg1DWj9wW5ZYocYD7+3BM2TXwlHs
+IyUIWQJRDwuiCMMtPcOSJdqfpHRnCbDjlRr4HPlkY/k1r2+xP4zM22t35V0nmlW
HXSEx6EQL/uakQ95BhBQQC8f4S5/fj6UWjEtV91csAdmbLScVUngZC+PnWP4rtoX
atdBTbrIHWDnW5XXnKsiDYz/KG4uvXo5/dtg+L/qURFDZ3hkKqz88NXgOzEOSMUK
7QqMaCtZ7fmbaRdylcP1nAKyK3PTpnz9QgMOez3Kdil7t2+pc3ieiqANaaDDGWww
Nq2WGahtMrKeAV/bdEOBaX+bIKAFIWjygE799PhKukluXvjPqy+1+Rco3Y08DM7e
kA7kK1C2Vm0Av8mEEoBo8WACbdpNVwCbsm3W1JtEA4FbaedTxgAjrSap9czLF/4V
ohczFx6OPfHUyazNzFP4CVblUZh95uzAZsi6jsSZaKVJs3ge+RNnMXF3uRT/UyES
9OJDEBm2HqMXQ/qwWZ3BoxFosJF20nIYpyVN9tB/MwRgEotMI2fkcrRn/Tch5Qlj
HMkrwijB81zOWBZXLIEV7jTENqWHN58m0Bxe5cBZhgQDvuofekYsVNpqJaZAD27F
VBDy2qI291ZNC75Y8cXQlfpGGjKPuuGaFBFYSEBtCsd1OfAujvPk5j7sA6bAFOYs
rqLPaYJ5LKaWFet5brTqAgDddORJMLJdQ8yhruJTmB5S6GGTcyM749JoYCqDWB08
qG+bw11YlN8S3uYi4RBICyRqvwFGUKe88HIPSoCa1cZ+2rlhsewS9+zhFNT9srmh
U+yxuGYVUd5qAWa+TJzr8v5V/fSzlGQkNemCKJtvJ2dKgbxVUUYvbvDnv6+vzduV
z9JYkPDPN4IxUyuhMHM374Hqq8QiwAgDeJaLi+AEICsKTWazhLg2dM8k7+fygm4I
6XkfZYwBxSN5eBkYaLPtRgH1k7cD5z8uDgScfbAYHeWjWzwaz6rDN8AXkmKTbDpD
dOFrYcmXv/8P0oZtkJntN5mtxQ5QbJqyyPUkQjDciksTDsfDBpe2EI4L8c0sTa84
k7nIN9DW0hYVanQvKEu7u5trC5WkDpVeG3A1jF2ABEEnG3Ili9ESdP30mZ9sgA49
gM+FXcGM2kK9vMJpf1IGFlXBbbgwrTLOL6F+0VWUokmslUeJ0LJgjjWbg0XS8gNV
AzAzsKQH66KOj2GIMmat9GlAdmXat8OWcYfXwtgItrF7ZjmavIIdTWJri8RYAPz1
9VTkMGmjeo83fGttmErGY1xh/wJOzEz6xNdn8k1x5NTMv0egvpa+E2dwQSbLqns6
SYrnQKb7La2uEwYyU6selH4fJUjcHY/H8nurVeEsVQQx4RGPjwYRPNJ46H58lJiD
SuTsXd7UD18hZsKLk4VkTn62zuw3gxX3BCvu0HmlrK7/hJCg4klFe7iGJiyPgBEU
fYQ9EE5exgSbMiTB2Z0JyC0oLOuvInB0szRNt5xIXfgndU8bf5h3AKB1q8arOLYV
3WfmUAWwnOisAeinGxj5H4va5CusXVV+NeRZ0rWqP+etYVTyF9iZnUCLnFO9KYb6
5rM1YaoJZRTziQhx7hHUgRU4UYyQlBfuF3Eha7JHip3R60jsxw2PyNfEToexV1B4
IEzwje5cLAtjMpQK8Fl8fJpceXquLTc5Xg/qQ0FZPiKGGzbz8ARv1Ht78P9BBMCd
Fa5gPEBEyPgcVim0nln7PPaCWrVT1S27GLtdN0XooEFdTcLv6bXOJ9V9bAdAAruH
qg9sifgZLqhJNaBdmLWQFL35qhsXBJlndBOw3AuPsdA0ungmngm/20dHE6S4W7it
I55ddb12UBeInkLiUF8nQ0msGWrn6f8vtTngzERF7HZqY8hmh6AqXmj/pABZsLV7
Lin8HC2RHrAqnphYGIRpDM7ccTC5/y0JGrMMto1de8VB+N7rVybsjyP1P+tWCeUW
VpWtP/vH4zi87Ly0oySClGdhpJtOKVtmQc5GztJohKzYdkajOLr/aZS7SXjVpQKG
sHGh0edfDNAMxp2F6bQCJ2XKvEjSry1tukyDnMv7/US22BOGFhazQWkxFoJGkJ1A
cOlDoaf4F4gxoi8XThldhzeFDI5tfoYDPMMdIBA2PR8q/76FlyyhC/wGVrHkR35n
XriQcm5eKLhuM5n+DcuImbBehLZlXW4fh7mcaaqw7TcNppzJCokDA4EYr3efPdYQ
FkTsW2p9r2wpILwf9d1LLwglwsix/V7h54A6lzutdDABlP+7VIZ4+kxDLZ6OGM4V
2rLcH/s1lM68Br5OaFS0CYJz23KdKyE8UFwItOebOPbCiAH5iEI9BdaUG2sAw7wk
hAq/ud4WoDihkIVhFm6XAVy5YN2qNh7yo1P1d9bc0A0cYKsdxM6OEu1Tb3YKAfbc
YO2xhd4Vn10tGGUTDFgU9fBfPet79P2w4aTrpv822jtTGI+bhjN7tQ0UGlRXTj/2
XRdS2tnmpZugDrcmhoB4I5a2c8CN/ot68z/Sm7681GxKx65HusVJzD7bAWXxaQ0q
Re1maeftd3gywqo3Hqcng1i9D9KpGDCucE/hjd/DNmNLFBo6PNS5phb6DaTHh0d0
M/VtISanmBBnG8wTbnbhBaO3etzAx/hoK7hMlEtMlZN+758PI7vTOBDct5NNl95k
ggADOBLo4PeLadsojXXs7tpM5amB053xRRmbTvkgj0Mi49uixQU0YbCTLWddBD99
3tbiX+83klo4PINfwKnxUHoL7i1R4zqWEjApVMBFDErw3kgKcPbU6WyRxLhJIAuk
7o8sn/T5frOvoPv8ZeuBcGd3XYch/hRKu88bsUQdnQMSoZ0kpqC3F6JRSa07ecbo
JHjEASlaQrz1p7OHDkPomV40V+GJi2oGOXcoNZF1I+/8TrIiOUfisL6vshRhiOEL
a2n78xz7ekP8BxO/F2tLSV+4XNMfsTdxsvjtfw5NvdmMRj29/56TTuMl2Zeh4Hk8
ppP5+kk/W4W/C3S9DZ+ZrjIZgjoxzEfvxsD296frFrAkZvldloMovYj+tPsnW/xI
POePmS2a+LevxuDwaNjdNaedHFQbWd9HNcZMw4vnlZyyewAeWcSAn2DF4in6J18Z
hGZLl+cMC3kV6qbLbFFvSRTF9e6/5a7HNFBtlW2QbtmvQA48CSvmN6aNZq89OMsj
wqalKE6ECZq3aNMzyEZ+xdfxF/6ft3tBK68+b0mgWOtmIfNM5sOAK8n31O/tCxpL
DNI9StDrac1q5fvTEi1oxSZ6ZlTJjnlORJSKEDeYyGNOrVI16hmvWdxWU33JZkbw
VXil5a1WuO65zkzKkYCk3FWvkrVDPrekYgYtsa3VMu3VD1LdIA0gJ1Hv7nFxrQEQ
MaDQ/uWaMTBCFK2X71AyliIkR9DwxADH7MoRE3upZdgMqXyc4WLqG4ibqbXrlIaB
KwKctqrsek03KQvKDW9tI+g9Rtv0C659XpCzCaH+ovv3+Jp6WpwVkChwuIR2lLK0
FeK2FVszO6EXFhIv6uMEtX1v0yGbIN+/Y/ZPSBvVTvumGHBIXnz0rn7zetyt3YcW
Rhcl9J9QMT393YgK10jsUVebAItsEbI9DtvPRH9woNhIJg7V3b0b8WLsMFkD6fHp
G0YdMyQ8xWV55nKeBtZTABLVMPd7Ow03/rTSzKO/8nhpVnmRHFysoRoU5GBYiEjM
zpOV4NLR2MI1IUOM7vcbBd75roL4jqgQ/szh9+4LfvqEG6002DRbUvm75MJj/YDT
66Y+vT4LTTKpanSNF5jlwbB/ZYt7RlGJx/AHY1h3CEP6kwbWQPDEkRKg0S1LCkP6
lDtga8DxjcjFII/KaFwVSTOnnj+Z8W/YlZIa2bhGRcpNylUxPej9RHtmbA6Mt+f4
p/gAVMcajvoJ38Icjm2fCDiRObad1ZAW4QDsCha0l2OxMzHVtOVSAOK0wKapaqws
MQkPQtL5SpMx+4tiy5DcSs6Umxn/v5+aav6D83agt0vx0LgnpUAaAOVw/QXA3/m6
HrtXUnHadjIS9OEjcDRRWD3d8g+BGLpnSwUXlyrjTq1lhdP6SOhb4Nf5ucDcIB2y
7n0D5NVahC11KpZa4JwTGYD27wNpYZyecS7ApN+T0P6W/8rC8dl5n7yHm+U9cPTV
bzl+ewtAU0BcxBRlkM8gZYUt607SWYHg5l//po2uekCOA8APZUHqzn7sj5c0TSq+
49lDAHwU1A6SCrm23l/CjPHPaqvl+CJIIiRD+6HEc9XnaQg9rOdG5Zq5pcIUAb2j
8h5NicoYw+5+iPj1CyueJ464z9vcu2a1rX5Dnka0m92lauRo6KlM7xEm9iSAC7su
BNcdHbfnJUdg+fXkKSaNBf0pNpzpA9vAL8r9CaE68MvWP80AKWVz1wF/jGR3I5TL
x1sCYnFK7LhsGwnVQnUxtN3w4zkXhRt74RwtIzHGtpZAqe1jQJiQJPXBzhoiWDyA
SZJbZOf4eJMKLh/ZeXDfYf6/9HZv8nJXG7R9VjF1FBebD1f8rdjWAJ/0gEDGYbMe
SIn7nvriI7dA5trI+Rz8Cm01qnUorUJ8eWTRqtWApVPjrGjbAYg6lM3zCYbc41zN
FPmUp4pWuwiUYsEgIRZY1/TQVI041jDshv5HUHnKGYmUAmzPHQYYHWnwoOFAVYzo
SoGnZI8LVRyAyfk2A4GIX51jDGsjRUsjirtUzJUPgQxkW3U0kX8KgEb2L1QnXhOf
RsVYSbKDQyRIJUz2ja/3ZFAIWr1fToZdTD2zMQOZsG1yaEorknslUziAb5zj4G6a
paF78/3M0SBCbgY/XUMyeh7JzzTleyJ2h+qKU+GvEQEEXliRerDRlBs38JRr68t6
h66jEhvK4MplPD2VoGlwz0mPu2VtQG0T6KWuSEZRwn2iJ+7bHEcMJwz7fvFuV+RI
JbNTtrwIsQhOsN6KG+Yat3o1r//lCXObhG7Olfi0bg/nk0beYQTzRXX2O570iXmP
VJvlxI0OH8zStbhdoMJ30E7tJU7s7DwT5nrVQdg8jD/HyyvakPCM1rfP9ejGeFF/
NwHThCpwhBFJg6DAZtOSiTbg4MslSk//8QMavQrAfYjdcXBTXP6lWBX5UK8Nok9G
CfEMXyYVoFsRcUBp5toHajX7b4EZgUXtX0t3ESR8cQZA2wA3RH0mTYwoJDXITwsN
ebWzAbTTbc7CusvVDd2l7KB4H0xjsugKFGxtJsvsdo0ItiuzPZMmkwN9tnjU/eug
yZL7SmS6yXWbwPsXi5Nq+aUDpAPGhpPaCva4ML0OS7I6cUFD1yT91Bj3dj+JwA+4
bgGfRxNYcuqCtWpPE/2thk3yXD5vWqMG1P/Luxm6kr8iwykTzl8SnGBUFOULNusm
GuIBvZtGVQZr66ppRnKXVYqPZ2x/k1+OaDKQ7cJhU+Uc5+Y/NBHKP2nXhXpdbrcj
X8QAe+OFRzDXieh6tqY1ddXvrtZOxASBFRvH+Ccu7ji+8DFWsDAvwxdD2vj9agl3
eCJ6rQONSQYZkP2SYGmMq8sUn4Rr4fZDsx+ignoIEYfp+ozUuT4SHobcAsiuH7gH
g535gc466HJeMvLeui/32PcO5Nfn7IYMN3LSebldY9xohs4R03oa3oi+V+888f5Q
QpF/ulCfLiMFyCQvz34bgQSuiRlTOiOt2yZYs53nf0Kz9oFVhyZn0eElSvV5xPLA
X39c4Z5PMfDGja64X360bL+jkBTp4lAM8ikmk5trzLVsPdFENWoazL1EZdLdZBRT
uLze7UiPKEybJ9E/AHiF8yDt8Jia6soG7LvIiSigibnNyBnwwLNjBSrK1dqK3r3S
bJ9xtMJiyRFTCSaKLQLsye91+nH+tjxUGUVzUWrsG6hb3eis4MooxWM5QM+BzQnT
/idVcUBOtDkNoHk5qAzBQvA+eH7hd7LTYjRVi3f7aH5ERAdLU5869tuTbP1UgHyG
J5/a12qvCih7OAZx/DRfnS3gu4+zNd7IWtTWH6y6aD3MRpMH0QauO0n/mOXrm7LE
ZBN20rjQMnMsfyHmMKWQQ6Ho/OMUK013JwTnmRfP+NDMuULH+05SK0w4akarZ2yk
lGCfF5Ef5kkxOmsEfefweTLjSY96U0SwsxGpAKYucHOVrWG3Rgf2KvdrFX7AUDEt
bF7HNzmvRFIu9Ij0Do23giYVcEbX/8IsXPzQTolze6bcu+JxdI5lY8GTwkmsqi5S
Dli661nl33m516AJImAXnAGvYg4pdYDQSNDi2wDm6SSgQ3D9bksV8Jn3E/3fpOld
el2Ca5i0Ykd09wxKaTn2VR1hTzz/85hoRQ4oCKN57edaHhjUc3xBdXsErSdxFABn
B0Ie4LARMVTFkjhj84TbN1TQmUQYvwPHiEB04lT21LCy48sY0bPc9WozoXCs08FE
UMIDVqrNQSg/v9ScLugP/8KjybroD6c+0Dbq91PTBHPG7hdauFiNm8cEa5AdzpJ2
CryW5EZ3B49KUG5fquOUDtAgQ08XqpR+JlKBfcO3SdGsb8nnay+Gm8cbpi+W9zHl
hL+Ei0AiAlw5Vjit3ARzU31JX9B0T3zqIpd4Ig1cFbCzFdwWlmgWVy2kqi2pMp1I
lNubxKk/OJ85WbOV6yLTbB5gyz9FH5k0P86m7kFiLzRba96aIbvTfUrkJynPLahH
ybsHhE1neLnNjybpDDAhn5HP2P7dcVMOTzUeCfZO93r/JTbh4q91ro84dlr2r2cz
6fGKIYHzVpMKR+IvAKbc2/cepqsliKMF6a/NfntZAPQSZmT9IAG/5umxtKlek+EG
XW/wcYMJzpkkU2M6Q2yTi7TjW5k5Jjoy9y9ENlvoM/kuKtRFpbrBwHzAtHi8q/hY
hyvY5I7UOnkQ6sN5GwBnNH1HHkdv06BePZGkwg6GDfUzMIsmkcUIT9R38hovaX5n
1OXjaPl2hIdCy+cgnZSM+pQJHtcl12C76OYZJEwXQ64NV+LBdd2m5Ye2gQpdgZIe
UM5xkl1/sabYXK4LIUzD2qjQ+H+Df6cH07zxOaN7eiPmJ0/rnLBuvwOpX0aLiIxQ
jFfNwDHUgj6siBkuf8U9JA6H+1ah/0NgyJ7mzIUpTeKUFqkE5dG1TpYwXBz8fJhb
aqxGKIzLq77YPUWCDbOFvHMi8sWwScK+gyPrdZDgqzc5THPMb73UOr3vVZq1htGv
UKpog8A/O5nnbX0EJ2Y6rEa1WQHoWreFJjyuA3L85x1u1WCSNDdjEbTsotI1mv0G
lDtEab+T1xGGt8lxJzd9OdoH27p2n3KstdWQlr4P4oa4Ir8OvUMAp9+RYBI6+QH9
lWZQSQYzBjPE7sMr9KwcDm/+sZaG/l+Jty6ZAjvDrrbd+hsKkTgMvwVRRYyR33gM
EV7QlszZKr3Y7kQdsY5gfn4vYBhAvxFI00RYLqUXS51+rA0JRXJqWvAO04RHM+eL
3IVoV6ge9fRsqEnz8IvdKUPDwIH4I8G2+oiqIgX0x0ggKQjKgL6g6dYCm2iltxpP
VpEaCIhnZZ5t6EtO7TQHyFG1a7QkuLBUcIZhPqkG5FPJAf4pKwSyDonfJoAQr99x
TDWazrQ8ilLE2Q86WFvqP9DRf1s97Lhx9VSwPgQtVc1uWBeM9hQtm92jaJaUv6hE
AROcYsV3t5ASlGuxBVaOi9ZTjM+bHOTY795j+gYhFSoct5m/Cp0Ss+1c/rIaNmbi
jCKekI3+Ikm0F2B85y+FpALD7XIl5BLTV4Slgj6tNm9kwChs34AgXjwamSYiX20p
+BnKNuVc9/HLDWmFYR2rZxb0PMG2nT16g/CsGgGBNwz0Th9nop/uh3JGu24FbMeA
4NAh1XQgdBPsSBwCiz3nDWCxGIEg6KPhTEqGd5v4AZnhiwgmURyKZhheNShm3sNs
x5SDpUrRCGbMhOhuHXoF9LIyeM1pD10eVz5YR2pra26aoeS3hzNpGXFHV3ZtCIOP
CyfpgmETX5u1M+ZYQYcREKK1TLlApv+e4iOApJOV46dWm9NUtuRHkq4Id7E3tnNk
+skYxJSMOZLlpFIWWYMu5iKPWiG3doG02kYlN4ZoDXWR/Eanin93q0geRguDb5Ax
T8hciTe0LaOXWLHGwFVY2ITSx8lGtwrY0hPqRyoVoXJr2fnEfDmEe7t2FDgUFrhz
DpI6YBvwPM8ii/1IKzSTGoGLrMqIvNvuoe0ZYT34y6X7d6Ds2pU+gtLFO9TZtpSR
EEQuLKm8TfFbSJw4jDSut6D96Y1ZAygUbbzcVfcmMQ5NnKkY9yHzbuITKlp04YyI
vNNUbiZn8swjBf/A4Z3pHH397topHffii1LAs8UFxdafHZ58pEDb1hxlKNO8dk9R
3oHuWAcUibAIcqs5fwCp6QZyJrA1F4iOjQeaFV8aSOgvT88ZomilzzurRGRqlAep
afJ2897hj1jzr632DqL0z9A4M5ASFjN3MkMC8m3gT1G0wJbPYNlkPBl40rl5u82p
2wI0uo5mSDMSV8uPLKtmAg/VP4Z3YcMKmvp0iGWxZUkJhfKX3e+ZIUOXlz1NM1uV
awgsIK3oZxcixLhhA4PJ9H7FRRv+s1R4+lfHqZ7W15JnxdT5OrhGR9N+dV0VyRFD
2bUXgWKawAsHUOjaXhavZYs+/df1R/ckngUxWCdxCLkVRGRDTtVKm2emKClDeEH7
mgho/wn18cXLtvT8ottCNZFNnddm/15SvIfE1KAAeEu3U48GgKT3K4TSIZisgY7L
Zg/7zJ6lmvPplxDfXwwnrtibf/0RqvrdTFcP7732kt5bzMCMfTS2BVWKCvpy/+Lu
Iv68Zuk6p4HR+99dSbb8MMvB7liviPzjWKMUBgQW6jKJEmAKgpm9wb66FLh+1Egv
7sp60XbKI7lVud2XF6OtEIlR2ASg1lLx+Maf3CYep3qiNvCjVVKEyZYO1GkR1RsU
Gxj6Je8ceGP271uffQq0nD5X2rXM9h2C6mL5UITbSg279rBwzdNH1esUnDRojuRM
16wXdPFuyWQoFLLKvXQtagXSCTIbzo//rUMXpTLItEBhL0u6ByPQA4dJ79EpuSkP
LQrW+Vvm4cUqmCj0JTchAG/gy7GjgOZ61OTS4FykK4ZUdM1qnud5IgpngBk8m+bC
pixlOm4QHQ2Sq0qbAE5msA0nlbOBUH28YUISBO97yqozi2TfaDyvMFoJCSRbNBfJ
to91CNEjJoPAYoxbtBlbxMs9sNuC4Wb0B7Ost5G8ihkR2jVVO7+wOrs10hZdh7fY
NvegPh80z/AhN/PZ4K/Anl/6o8rkQH2Dy7iI5ji4KfPSEA4DA1HADxarETmHzY6j
Nf55TamjqFw6vcy7vtlve6k1uD/j06tlaQwuU5Q33h24hQ7LKvDugy6vs1pB2AHx
ik6m/Wt4W3WrXH+cz8mDpVET5r9Rgsb8sech2e+c+jk1gF6HmxWFlX9G2xmGv4/m
ARYnVWNtBqk9eMT1UsCDGRRkQbCOMCpfWdt4MNmp69yUFfmMCDkQQIoVxAuNuwRt
BNGtYN6MYdt0OCAafokdgfD64yjhm9jBV00gVjJV85M1iAfiDXxQu64aOy/Ujt/s
wwK3iP/IuGBtX0/fYSTYThtPfsSA5h3bSHTijvaZEzhWjJee+2Lm7qWS82LIG16V
czzYT8sZ82beqVAtMRrneudRiUZvCDLi8r7MkUAeXFoVAAxyO++jkAIrjgHvEdA+
hKUsvXVSZKGByspsyvsYVpsQTEgKA7R9hwiyxgQRXxBqsqJ8Pv7qAplwHjGLbttu
/Jxgx2QrwWlT6h51gvoNTWM/kKORAI9dzTifZKkNTmRF4J5GmBsr5YhSA+xLcCZ1
0h90rifItr807pnMc2oPWTDtGhXbeYXPgk5qQ1uUTDyaF7snW7E9+5ivwqg/22aS
j02E3KIYJcbPXpQ34/kiDcD8zE6/lMomkNKsi1j/h1gzC/Hflz7/l4EhXiaqtUz6
1+Kpms1vk2QP1P5tRRNXbZuO5zmr76wUVvkElgsnvfNpOXMKOD0BGuc0orWdWZLk
sW5oqEJAkLgycITTMXtBHRpSUSmhgMHCVFVptwuEog4K194P/ax7R6IS2kAFTLWz
Xg37Zo0k9RuFXlL9m4Jm1gfWzEkRWqLtfhsfb/Re4Qwb/SAs8Pef+VVNLOCZARZW
kaKsHdrgSZzHC4EqpUteoE796WCfJeIROGWNeFoZu/d16JtnL5PhOw2h5jWm0T7w
ISjaD1llQP4IVPCd1ks5xxI4Oa0Cske5B2/psutYahreHUNdFY/2AodGHa7lZyQ3
T77WjzDj3a51zRRM3SvTJqYv0VZ+dcFjyUL7mBA5tA5jMjMUqPyeVKL0Kvqgsuab
fAw3i6gStn5HpbsfapN6vLzrR9QapImMfRAwf/g6NDNFSKOjHnKlVSs+TG/2Rj8v
AZNCxZcOYnibswixwwdtvNWj6JzduhLGe8SdBvgZeOS7k5XzxPnPRfC6OHdtzxve
y9+xE9gHpv2dW6SUQooTxbjBhpLoQyTsfmMLdQLLNUGOWNBilxwHTDtC7f6DD+0h
r4JtFCCOiG4gtfUDebH+39c6+RdfzbAyUy5K/P/GTpoDdmsdza260+Zjanx0GuyE
ymnp1FLf6AWMi2GztuVtKwk6I4KnGfkEdkHktaIclzONaJMQI6Mdwrgdj0a3HEd+
65ePXv4TElsTXZZfG3LpxFI0ubGiip4OeM1uIfix1KEKwcBXm3ffn82yj9qx4exj
u0WPKchHVnIY3xLMAKJgfs2grW+O+DWetop2h6VaB8L0lmw6R9cEpZDc/nzZctnK
W3DYA6j9tlP9hI9vYOjJxtdW+505bip7S82kmr9wj6QKOg96nSDjTB00w+gT4lUV
sTpIet0g1CJcNbVO2MUf8oTEfDrZ9T9rXublMPgh7112sLjmlPCV51FiRyzzrepr
13HShJ6Viile3UBCmRAA2YrwZje1JGxVOTDklFPugb3q7X8eYzdCtiwPDTIY74Zg
tDuv/C9fUff3e7Q+WAC2jFEQlVxJEXC7U6ieN1KpbfnEzDIMtgHIrKUwGPcn5jgM
EJHFCoJCY/vKAHSECUoiBO1mP9JesHq9WuAnuGV3eUxjLd4CpIyy8KR+DSLnHb9m
33F5r/PziM8i5G7fPNVhTi+12jPL2BbMAultrINd/+nqn4plzpCOstqVI/eKeTUm
2XX2+msaFVs+4XHXfAvj4dLN30vslQrscPsYYDNEHl6yQHRhOXPkzYtioCpf3car
+AMIZ2NYQa8SyuC85kimKSct8eCLkeRutuaTFxBtD7sqqYif94RJDSkPHetAfEQ9
PS13kZY4fUYvYQWK7qizph02YZOihKCeXGGjEOT0tW1fIyk1DsDHdL5crV4E+X+F
jr5EZJZAghHKRn3sGG0NIYDDj7dPxGPayutPNJabZldlGyaNfzclbQQtuwLuZMX7
10HtwAyqC0M6I52gd017rRUrkOmcKIMhpEj0v8L6xMD5GSffcbFV1x8HghR0aSc3
nocZThTjd+up3W/vwbguzcc4gGAqYW7JXUKefkmRXJYt+GSXVVuUa2UjIl4itbaX
lDwZ/AGMxt4f1XeVj7Sbb7wZsI8ebWXr66g/x1fPxhu9abAVr/rBFOk5owOBKPZf
AFjFC/UQwZ6pfLusVmrBetD0xyA7S4vuvaaA4En6t3NMXXgqwguDGJBmKSUvnNmK
MDRIyYZ0iXveGiqGOC1Cot3qFTSbeS6xbWLsjGkn+aL1SLGZ0HGT/LJD8uLV3uvy
fFtaULny6s8nsWz5wWLZ5jCrTQf+swcJ4Mxlo+CKAGZz2urW/K/DP2Ez1TwIPxrX
TGUckskSRcXItbYlm68a1Gt3ybXWhEl4TPbnHCoZkOSLilWEaY8fNfalajARwQTD
GNBdHurJuROCnDOcdpjU1Pk1GqZUUMfnMlMybJVJUZZk1T2X72WuURU1jpd6nW28
0jlnNdqonrcm7kbxfZFIPP3BpzbPvr5PJ7Ox8tx84icRtNXytRbJ+o00guE3uYuw
qG42LQidc4xzj97nq5ntyOnvB0QUsGMr27Q9lpWRRl3rYl8zsHVQ5zmeWbbVp2KK
08/ExoxRYQieBkaZS6Vg+tCoyTRmm/604pYjjqDSCCWxQJUF43wRb4Mhm0rkXosz
RgJ7yXKdOOmCsnuUn8/dyvMI1Q0JSP0X0PIIi/vhJo229pNi01ksMRyuL/anClkl
8lVohO/h6fH+miCdw1pt0x7qyMoLBDCtUDoBsx0+hESRSIZJ+8OXGfnEHMPVnCHw
JN/pLoDDksg4AzprDC3GejrUznvfxjQQgt8UrbwgvTvBVNWbosjfBMkGEB9Kpo+R
Nk5dXcOFQa09TryYayLaCQNW8obWP+dPyxDhm/nJklWW95hOmkrO1s/YPhkDW+NZ
37Zd2x9VDssE2WqtWNabrMJAXLYuY2Qmqo41rAJHfiwHC0B5uxx1WxgOKeLvmpyY
XNXg6sEcqnjU6OPFJZMHyfHx/7TVKOvDWYW3fVUlF3MZsH17p60noXY7EQ0ybff4
Ycc6nPxueMG2ieG3BcL/vT1arBrdNUfNbwqJfrW9jYIjunCUzAO0TvUeAlxHGBQ7
RQBLQbEoo32xC2AS61H4JFoMgsOpmluGzDok7zMCeEZIQ/5JLbGEOqtQPx3cHw3H
m/z9Ggl+R4HFZNk2zIsIp+0JytwwIiJBSvXQE5LM3yThNmW8SflNhdqFbk8XcfUV
soxWqUXEzGJsymyXxi5BO5FEbhmyz2ZaCKCTK7WYsUlkOMqBPwFQK6KxD4MZ2vwx
9gSQpehwyGq0kK52mu1ZZ9PGiW6O/Vet6lwRqrv4ecGDteYSUfG6cyMvMt1IDVSP
SJspyt1NVvZhERi/FmHrqNVUgklAxiOwT9va0xzzckxBsxHcWvTzelKHa433EwTn
ilDWplNRGHSiW1o81fLQRsVaYo0SR2O9uNLZNuZt6LPxuwjQjl2A+YSqUcnFVhv8
oZYS815TD6T5H/NnGmY7A8EhIyvIVvyIz6glh5ydeC6G36lDnmLuKqx+RwGBF5ah
8pdRjwQc86fEQtsolRjYhv3p5smwTh8HMcPHdcIjpotnoEBU8+iBVCd2p550aQcL
XxKoRcUujsXXCpnqrVTZAXk1HRl5O6Q7rU6b2qv0xYFSnxU25Q4y3n21qt/jEuHi
nD2ydWOkIGTp56VLwvGY79myGj3ldXabTnYmZM0b/5Cfl5hYJ7Ub55Tew97Xyeu3
UGBE5Kk9TB1g7CPYnZo/fvRqo8ubyq5z8K1O3v6hJ8vHEHWdzId2JIUs2OY0hKWS
2qp86jmbbydUGBHWf7jgn4VmD+GJj5nTB/kz0UL5ExepRmJGvLXuCppRoSsinMMp
H5l0RdbnD7SCx4mLxWaaWmt6hV2njPHanqy1dXcK6363sEahTARhhKJvT5VvGEoX
bnvp28w6liwmOEXWfAk3t41K29EZe05WEpmzHv/odByTWNmRhfTJpfQ7gWJvchQv
wmqLPO0wKeqKYnL1BkZ50Zcr51dubkulyqPZyhKQRLr4D7OSaq0p3q6Ek9OY6Lv/
+WL1RdLnUEmyQsxlh5F+Ff3L6jurRIiYLphVwwQnZdttsVW/ukYZXg+by0G1/l9y
GukjyFg7mLCb0Hh3dFR6duXVoKy8xR8V02d0Jm5epwal9fUe1SIIIfHE2Y8nmyui
afYjJ2KnrWcUdJPy0BsHj57RaN2MGMlW4Gvle1cFtJ4EDo0zCXwgkGGC/l6oV1Np
qcuf8/le+X1CdLKNs0ubSt6v8FjFOvTmgqLLriwjrRO3X8gJhMs3k9kK5Cm0GmO5
M/qXXwHvOg94uBXqrhgLNQM7RCIsqpJjPg8T59UVmVBAYOp5xIVEv0KYMpHAGEq5
jkuH0CJToSOVXnjJx9lRlqqH4tyrXQ6Dn0nTunzqXFtcR099qtdux3fEuLfnZG/I
XJyu1Z9LzXu7EJ1MAukoTY7NrLkiRIL5dDNzKyrDnYjmtPUOyiNtrvLi39M+LqYE
ARNjtW3sJbAKjRgtchS1SE7S1NqNd/SRCgDdpy09jSUZxqjEAYfc/zrKz8hGz9ok
m6LXpxgMlyc9YoCdOnlTfMZp1cR2U7wLz5eRdJJy3xdsfMqkGLeeo8fCGRi+tJPG
1aXpODcxY4/+AA+UE2DYov5Uj+Ev7GMlfCuexG+4Ypu5Ff2Ov6YOedLVfAiSHvMN
e/OZst9cKfh+rghTa5l3CVCrJU8YVfyTqcs7VTKeiLjVyqyZqoEQrwpbdIvosbdM
tdr6McBy+Z8ZD13ltGMKFowOkwonU3QtWqyW9ghDXR283m/BCYRYS2/lNT5dleDN
lhqVoGJ37NhhysdvYGYdDseygicNtE86RVSvQ1gd44y5fhuJbT9eIUFk1cMhoh4i
s7DZngGYswYE3RUKumaqP861+mGf013aviCZvkryrrzj+UFMibwZKVTWPQhs2icp
2PeEiKt3931KBEzoD/wO/CJt+Vv/Il05oWiaANlZbDwHwbFqwtoNoxSQ7yyfRVNy
b8vvz9F0AnWzIBpj+ERdplS5arChwAqc9XKw3T8s+pPB57AR0onoUGJZy4J6SIIW
/hcB0G6qHXKqGUBf2BLwNealuw7aVllixiWklBfn6KiCX9HMWmuLrJyWxH6TgObd
xBwDz37ytVEJjYiPIBTx9LPq6CQ/VA9hRwG3oo/wQeQASuqrlTL4fzpbq4yZO8Cc
kSNdZKL7WOClxK57RZ2PtAAyW6OmUfe4jDEn3x6H/j5XzX1C93nVRSsBB6dKFv6q
mAbgujQRsGcI2ibUcAmZHKf68RkmvmwcViCXnsUYoIRMyG8ythVcRo+QVvt1rPYb
YFe5mBDatkZHQ/rhzXMY+PKT0FA5Ca4aXitPEj7Q8W4k85WB9SZwuB918PSKwVx1
cYKDNjj6DjJTZbWtR8y9nzzzzoiMtxdZ1CLiVkKw27eo+Pz5H7gf+doyuGabj1TP
GcNFs1S5HKo2rO0FOhhg4B9fyIyv7+W217xnF0u9rS/kTNe9nGPzU3+CnLGI4br5
J4baB56FchEyO8v+F2/4w9U0AU+CVfLDMMh3ryNJ6Mi4ouJrYfPL8YXvFdOWaean
2afZHOJJxSkmRU8uLRwLtx8v3bIBRJDBnUV3GtCavXFcPL9Z1DHdSifbPtLWESHN
py8+6jscxnauaFWC9BzJaRc6NmvemswUDKCrff2/DFddYvm5UMdxzwuCPV0IqFNj
/scgeHBE3ByutxabwHKSIgzayUSx8A+IP/33aCrnKmGk5UfpvrmfwSsO3Lp7EZ9x
shGMJU+3lCsb1Vt8P4tjRZam1E57sab+IR9AFI4W40oGxJHssRn00KuGaN9npSyq
om6IRg5kll811R5eJP1sXCAfOs0aeIFZEZnHXknnrUCu1XxIPMDpk62/sH9UBJFp
EzZ0NJTvdt2b9kIVc0bm+E35nXeyQ/p3Aqc1JYf65E3TbRfPzaaP5EWi0f+pmkeK
RRfSJ4ZpWlZeZVOkhwABxZko6C5jpx2LGM7b1BG3h9tU6t+TIvCrmUqo1kJ1zquz
GpOAg4TEiop0IvOj4jEZqgnD9/Wjn/2xb6QDrZIiFekjz1dyQRs4VfGQBYeXUL4r
Xf0eRYkYSqULMoZA3c5vh/DLc4rcDahNhxua91suljNxMvxRv/c5GPcZp8zxM3Ix
FPkoJukK+e6CTl62qsh/c2qdhcDhu6bL6WKPVpGLBMNrc/9tidvM4p4uCuWug6ZM
LGk+CRvkJABe6+Z3i3Z6CkRJeelVJEXltHZDxRDWohzd4BxwXz0kLW4Fs6DAGcwG
TNA8mLo37ps6/Vpzfg0Idoj+e39eRbBT19/5hBNnVjA8Etx+sguSAIr0t87/telt
F7MTTYXFiJR6aE5xfF9exn1D35cApCbyifx29RAWfdB/seEAlhByE4N2RqrTzIXG
DO6PFPoqyjYnkEDIjidy1ajyRs+IBjLJNVXc8xzjUO4GicJvxF5d7VfOlqSRYYvK
tgug46UHs+v+wB/wUfKp4DtpP7JzERH9XQjm5A7serM+5xvyrFQDtIsnKEaqgdxN
/e5ENfAKV6Y6ko/wKmdCy7v7Uqr2qFkyqjZ14DIsnfYGed0pB1RBYgeGDE56OU8l
XPWXJlPgxdG8i+cHouOy+N2sejsA9YDZBWVeUhJb2JlTLfc1hXlVmc++SN8lWa9R
OtKNuXhNFOrs33+S+cLLqucAj65/R4Z1SCzyEHOa4qy3wQp5bpcm4Jtfy1Z6elZV
qiTs2gYFfasExau+iOSyZ4eO0BjzmsxpJfBNLRahk/MkxLtkxxwIFABx9+pzK4Pz
AE6DarphxmG+5zFAoWCUnhOCtlkBmQdY7UWLamlyKO4N+gpbtHNXZycKDpv80j8Q
CjPRrABvVfLYRtuLvI77praX+y+HlvgJ1jrTaVZwXxIzJxIoxzuB+nLB0xbUHeq3
LI7k0IPgz19tp8gCLYwA5jQEwPOqn/9JkhsXEWlNlZR1A8L84TNR8dz6Iq+zwIAz
hdztij1u084CR41VidI2zQjYue/EmRvkXAX/iPOfYe9RrWSCHu7cqR8des3DkrBT
b/KHMbL6voZVsnmB5Z8Gze1P8B8pmunHbSybVPYL33ouqairOOHfKKei8G+CmjX/
IoL8P6lr+3SDUO04tAngo/oNEFh8lClb3I3N6OPDKmAgo5uovxFqW/OPgf60gy5z
K/s5bgV2jR3sbyUQad3MUvMAFEzf63j1EBn9yYC3MyAMqEC9/WyFgSXMDnQko5QR
xms46TraOQrGTnO0p9uOdDzCSHks1xNH2iWJeuaIXZ5noK12K1kk/v0ehQ3PfMhc
3ppd1Aw1S8cZ/vltEUp1zTO2LRemaBwKMy+T1zlzbvPxNyKejwQqtuK87p8GFMlf
2TNwpVfm/NPSYVHXUyYng3u4v6xM2bjYBbm1VVEkCMYDFU+5YVIAGxUFmGr0focU
+9kSmCeJnkuep+lewR69fbptA2zzEpOBrtsPVHqjowW9BvYwYBSK3ysoKyZKYYls
j9fuxVRZW3E7+6BsAIM92mM4FupjDu6hNWzNXNiSWIOsnHbpWC1ZvDlYjy8rBemy
50bSj6i8GFEzTGPfsXSbuIBxK0C/j3Sp7opJQDg76DVBsMiOEGBWHMl12UWBg4WA
6Inut8I9XyRejQ4d4dUHIjmFakio6M1Ax5rP1URaLb1Rz3MKKOQJqs3EHzUH8r8f
VerKEYr3j6uDYBVRdoLaEMGVJ0fZwDyaNt151q1WR54qpdaFFBmMuaZoVmQ//dOd
VNqQZMeLE2whtfKBfzEgzzakcdkzI7TzbN//o6UYm3QZ+O9uYR3v2TKOcvmBZXEf
VHuLTf9u5XgXNvpDXYohxeBD4UpyZSsi4WaV27MBigV5jaFj3KYvN130jvElQFMK
cQ/nIuJoqqfTu12zH6+3h5Hi6p/p/1FfFnu45oNLaSrdw0hxi9YR6n7I9y9WSJwB
q2bLEgeTD5/nGKuuQYVhp/IOxvzgyp501Nk++KxvGOUl4QQK+v6fbmYCZOTSbTQO
QQYZxgalhMBolc9Pl59bJ9+ejAF4AEuFS24HSsNtziqFQmf8Ez0dxUf1zlclAZK3
1udVd2SaVPO+8RkTKaUQyKjmqNyf0L71X+znL7ZYzyLDR7JRjRlfeO5i3FpyKNw+
DF9HbQRrMfLBoNh4Bmtrl4RD9eQRvJmDfuk0xCSinrHlku+tQQHNYlyy9z0/kubb
WWxElGUdi7a84PHXLiVxQYqlO5O9iEuIfwZb/S+QbGbqHn3ZEtevyO9U6f3Pqb95
/IXolJu6TSMcGFQE6+J1FH9wAw8UvT90C7iNVlOvXGqKwXWtDq6BhlygIGPtcgPi
lTtNjmJ9F9GzsIOkrBkJkteiItY2Br2nreE4WJHYia/VXCJEEh0tAG4h5FVbH+1q
IPCs/mWqlIad9OngYFV31TRw2P+rJo0Lnu6Gtro4HLY4YWCVniYbCiw0Nd6u6MTf
EBPyqNAWuLh8i6Ho5V1nCI1CxCuenckXreRL8sH+UdgVaSnl7eIHiS6CyIs0+wi0
bKxpXzzxAsE+wJ1gLT9zRQm2tKIsyyQHEcfim2WV7cOpTIRIuU5zTAdE2Bm8g1fM
3heiwp2pBUPzrPyNpI1psHQTHalUEFZIjkCvd6dLB4tI4bZc4K3xaTkeFuLeTHlC
SC5YV4G2aF0Q4bZIVnn86b1xUfoZIMYYWXgdwG8xT4rhAypiu3XnXLWJ1zMzRQOY
KJuZDqsb1apeq1WrjuCuswc9JExFTFRRwi7UocymBAZ6YNN5AUMrC6wTBz1l784G
k4VDM+xN3tkZnvSW2wy6Q9HqW0vv1XXQYAPtFXJN8A9wjv+V2eo2KIEWRmKGpxZP
eLm9JkUHqfsvAznvz3b0Ntaqxlxb/ukeyJ2Ssrk4m5hJg/d5QiY1WKve4LmZW7Hn
I/Pru3G+AG9Q+NZABR7THltd0A7AgQ/Jg84l2v5AFJC8nawoGp9cN30MoCOLKIKd
cRjKzQlV/k3/vdz6UqUIMKXf3pxBJKMsjYR+bakqf70VujQhvs3OvUqRJVczveT2
RklipinN8bA62Abn9270vJexCmFO1ZAtp9PrgdBW6AVSDu1Pgex4scDczx3o9R0B
XMLFJJohKJLU/dvsjaUC3WNZKqA6QH9mH3FulfV/wA7v7n1xMTgvEQrzjpwVMQBi
aN0YfaeWwAxrfP/85vCQIm5uxnx0ZuNLUwsaOEUNbFdFlULNv56/BDHVIkPPQ3bn
m7RKpl9rTEskK7kd/vQUKmC648QT/+lExEu67OuOq7CMBgBmY54pY5YvyVTGDV0l
2EXHN+rut2kLdvJ8IsDKF2iAbdJG8iSzfJgTLhrj+pD9i6RbB6rk0Rez/6INhsvP
WNJgYVnxzupIZUEImVfWMMbGyi3ERBR4MsBerfnGSGzUiwcIQtGNrfC6jGs17tt+
xmWB4fdQJF5i9rSsy+hwCbhNDEyPqh+U2QhkinhGldnajJJfpBCO30mkuWm1F/RX
2kT8nxl94KVPOJCmrvw/t8KufA7E4izTZANgUg7FXWSAJA/ZQ0CPwZpGb7w+v6Ty
XiCGMO4DnHtgI76G2o1fS6TSIecp4UiIHKGF36oZkXZGMD77UZHDxXOpsVjhpEHj
uZuZReflYsSjDZsUy45cc3+ZeIQ5ObAOlZslD1JV3mzYnJQg/kW/vTi+1uKQlJJT
ganLbYUSEu/N/krenlGS5Kq+I7lp+CjXyR/ALD7PMizG5RKTU/726FGsawiDKukO
xL+3GnVOBO+LFzzCMz5QATrL1onWG3tRYzsTTjowZTRN7J6Yjpnv/uKfTG9Q3pFP
Ol4GcaqXE0WmSsJG92tliZNOrr/MmPbaouZ+/MJv03cq6SsWVHKJ/wlCBlePuwMS
Ks8SU1dlR70DMl0bt7DHzD3catv1HpXJplOI90NAOSyKUnmCj/vx1g8kSBCzz4Jm
yLZYD5USi9Ds1165LXa81gjzzctWC5IV+QPnLz2BzB89jKI1i/Hg1w8elItONVCX
++WBy3kKWNfr1TIQq4CzyVZQFGMUOmxWx1RXnYUbepEKC55QpgL8/cpNcwBTO1hh
ody4/bsUsaDu23SBVI/LcQgtU4UKOFXJwr2qkmS06DzA5SYWAvwtX+o6xjEBmKly
X77kOFtmU/jptPzIPK0otZQTm6GSlA5CmaGZuHkuMs8SStZKUEfQaK3J9NEE2/YO
15zHoQhU+1N2HX4BbbZ5wGRdqi4Fzu/3xNkkPF2c3Rpa7lXNyFE9zHNHlZwahoxO
nD8xZAGYdLRnzkJaEDYZgOAJ0v76DI+hNrOOOql1ro+ZkEQ/A89jJr/W2WIA4Ott
Ii1QGYhi9khTylC+7Rha/uKmzopL+3mAv6Nrvp3SslE48LRxONPqEw1yFRtHN5GW
xr3yNjfg5N+Paex1c+mgPYcU2A2ifEYmrj9e9E81PhS+HLZub9N7lp5DGPtx4fey
H6T3Ki1dItSGuoR0iQJNGnDbwme4VUqN8bAZXQHs9/1/SHd63QhYbdmj3WmA0Ugb
JplNzqjfgUD5meT+bjvaaehGZaVI8Vi5/yLhyu+zl/ULQl5L2xSbX9s60N7w36tn
Y+MXuuutKPfZJptZm4MNAH4a9Pf6v5+bGSXPMRyNX4WFcruEH4tee+glsBTubjUN
20C4ZdUoA7zHSRIaEieMxPg60qZZI1sEPo7tkzX43xxX3NYRoTBOOK3toK8EYuHh
bBtqA/8er+XAiazE8nhV0hbAzVtssg2gHj0maZRn1tFJZQoVKo5pdWjBkKg4G9fr
LmfXYetiMYy/v7CRF3GUZHP8IiKJdaL4xD+IYSbfGUHTUzdDjEEc0/UvROwx8WW/
lKaMb1Jv3ST117CfIm64J+Wpv+vOLYhxQ88hJkkkvwL9RQZOfGcuSSIvcpJq+YDa
RYEgXeseE3HEdvqWYsMC1ftyw/NcmT4ETxmwHMvuHZLhX8T96RFQCDXVoqIvPvTS
UpMkKzTuSJ+t18EZ7vncTnrMpovw11Yb6Dn37FPLhWZRKq4IPtJMDgJI+oSsR1ta
9rjny9qcSc1euaz6oOSw2H1s12aZ7wPRkaIimXpu5CeW52iHL2/wkVGeqEAaXH1j
v0ORgdUtBYQJIaeZor4R7+TEODUj7T/U3dichDbX0KQs4lLRyH7T0vJ33BWp6+4d
JYk444oBTKtUnGK1Hf1hu5EVwGCSqsBU/gxANJN40f+2/I0gbHsxoFayZ8QSC2AB
hYodQzgoEHgJ/Fgc3YjNJzVpfu2OxsvX+XKqngoGdL7EZbUdDU4nXHyHnjAHFQXW
9GkgnX2KYc7nuz/vKY3e4rLg3rngSbS3YptILCMNa8+iyIT4OIR+ak8zUXEfbWd/
6ytiqGeFLShEWw0gBSXDt9A3qgxCt0x8XSXI5hKFErnsuFhnR50HuJIDUK2luj0G
isGrz1XwJk4JeGX0T2rtq+2TriT4HAvV3fPvWgShNcvYBf/UN1ddrF5tcyct+3Yb
ux/gJw6shLl20N7dFFR0Qxp/DhdYFk3mTSrlU6cPP2XZmVhm6TOu4Fyw4Mesv5b6
Je5H996is/L/wexpUtq75jXGSc9EoaMITT/aAbx1H8sV+z1JG2mpVRdM7r8jvFPU
URq+z16sDsk6hX0yzuOsQg/WwhM4OV9/nu2x5lIN8Twtu7XSMH2vENjmFhTqak3B
lruHuaUsaCOKSAWWsXpxZPEcg0UFVhIDzwKBYUI+2IJ2VAq1CZ/hBJI27i1uPgZQ
zVah42BNZv9x3pOoWpWFL/OJgqJ3BUAh8CbaX+M4w+HE0L0O1qVFDDEWRQSiRAIE
VarWKEiHf+JSPA7ObBrKTtLSKvws+EdFIV9YDZuzMExFJ0/BcfqrK1Az4dwSuF6u
The/JbEaz5Ycsd+HXCQKxlgrYZl/dTdlxlFlyHCOrPAbwBWd6/JddMivbA+6PdGc
3ZBPBCoc+HtiV8pT7n7aJZX6r3XKdfmaz6t5elby/xtLxo/dXgZD1ei9HZX1AORa
+ae3wqdyvr0d97uQd01MS0Srghx6xUt8CiMO8bcu4/DKXH+SuB+O/aP9tlXjVBEW
At2JiY0+AlPpgGqCRJ/Btpe+jbTCB+dRKY5rK9ScSVEMxvhVN1OtUV9jlcxQdo7s
gpslH5kmNjnerTKgvCzankFpb9D5OYMA7oM3IDbX05ZJrZbM451iB5mKy3ENfmyk
2vOkq8p8rrssxRXLeIqOOtq5liF+4HaC3rh7dXO9NftoRhL2Hltwwoj6JkKm/5M+
ng33j9bdsKo1O+6Utl+6n3Y2RP9hSbRimQaNB1/TOQ5aJ/nI+ktrMJRqXUI5l6oa
CfVRJs//KfqY9Fwq8sLw4C3jwsPlSrFqk+sHNxm/bVbG9WzJG7cP3xeDweqpDpu4
TixV5vWWvC33FyHgX/2l1D59l63Y8jPQM2rmLRegFHi9vQC3LzEfW3qh+Wk7v+JI
UndI/OST8AluoMmnzZx/R4mH3fHKk38sipaNmFIulo03W76HEiPbbsiDbij8EoLd
G7bkJ8ynm9Dqp/uAMCqSLd8VmDM9BUtaGQJDtJijbFbkT1IxwM9nc+pLM89QVz8k
vJ785zFGOwzBUa6rtEgKzMUK9Y8qb9zAs6Lc2DpIm+74lzhQAsc4TlQidxhK2oH9
HMFG6Ri2QrUqQpHsWx6bDNGamdiZksTxinD6GsMmQoZ25udGIDQN2TRyIRHxRrRx
woFw6XhwtNz+heGMXkMDlkAlS2dnbc2UiVX2ZFQTBRtOkfmgTXiuJ/TN3D+OdumY
O8tpQFxNR9kpKBwYQjJge9ISR2Tcayc1/XiSJSf3uhs/UaiG2tuOL3heIF/v9Eaq
KIlRm86QzK1ah3oBXlfVXbzOmvzmETkHyblC14d0J6NQbN9vNrvhGxxE8CObK59C
bVHn5LpL6TNVtwYVjX/1KyGBnwXXJ6BEZJDoQj4Lb2m7W5TBmmL3ShU9HnkL3qhz
uXpb6ZOJO5DPWaCpAXFBzPInp7dURo5elQ1qwlPobOFIRYrwm/fwvR+8ccjRAI0n
hgTvjWce5ksX/kD9O8BLbdRO4kczJBx4i7J8/cUxCvCLPIzkD54SPo/PuxXlxDXZ
6u7dQOctS9TIl8D1vPjNE0YUK1bNrWFpR+yJMalN+C6p/b8sDfIwrCm45lGCLVzW
mgOZMGigQKYp0rW+b5rnThDFUi98veKVdvqZeGAgm23LwjdIxNK3ys2AlH1rI7At
DGIAwQI5gahnU/TS8d6gfwBJznJiNTOx79jnegnA0rhaDOm/fgM9eqc+yidXvbQA
Kj+TXUyczGZgTv/aKe0Rx2Kc3TvmYieg6AqfCmTHE0nbzhgnU461+GN2H8XKTU9N
THkoqtRdJk9tbPsCXZ4yvCNI7NbkdB0GhyMQpqZ/QfOJSiWbM+thUbmRxy47stdy
ATIaYt+KrgTxROfy63L1W+Pdp25+Uk9zs0vyWvXgT3vqX9aieSzpM87QcmVkWVOa
l7apPNAEGdpLk8yj8VudLcNx4kwrnX8H1HWgRIMzFtfQYx9zuYajQPbvH3GMUF4g
Gx0Wi3Ylucopa7CasFv0kT3tZszNyUAl7YRFlq/m4nCoVc5/ZKRPT2W7zsZyg6/e
AECe+A19r/hFyAV/BsnYKOakGtAxzjwLfWAUpmZYn1kkFUeB9KgFhKl3zWT2jpp3
xFf3yspzd/GMBsirgQFCnislJ21+NzktpmqV5gCe45BflBkc/jaCsuCXx5IaH8Ib
IIwiTCiz+0v0pTGGtEfm34t12wHWywtjMNhj5hgBfx7fcjxIXGTbhecmEdMmybYD
lUWqj62elPK0HKyZFjlQAAiSAZbsf9YBaudPT3K+QR4HbHFYpXfNh75fcQpIrr64
h6Iv2Too6j9zaD68mybFmQ+ZrY/HIAK8tO6s8ySXrPfWkGOXvO5EdXzzSaH0a1uB
34kpMAdFopGi9ot1isdEYC/hNCz8D8VAklyDXVpOGq9KaKkyDbEgl7lleddSfGVE
VYXKhoJq8R3pC12LgKtcqIVkcPfXCEbujGaJQqkDxyn4d0u1ZHEmf5oopfm15Ct1
4VLWO5n8gWVv4Zd9DYtFlcMhSQhtkP9++nbGscqY0cy2SBBlIcPYkKPX3FPkXaRU
MErbLy4RSfb32DQudqPV+0MADCt9I7ANFhi7Khht/WicXcd233BtpcJ/UcDwOxb3
Zxuf42cLBLMRtecLew1sLLL0h4wpzb+k9GZoZfU5p9PHPvvY6K95etowPSLVYZrS
zQ3jVNPdZG7HCEDJneqAQXDi9pfQ1xkoeUZp5ACS/aL1c6vp/C/OIe8FB68/rrIq
DHCCS3as+a9dDPv+NffCMxhbP2LUPMVk2eTfKFrXZ2YWMeQxmiMfq20kuZpc4+49
vIfTthVck81ViDHmhwwsXutwUYBbdnXQWiP+1nQOZ650Bv7s0qKT4owz6/i/xQh1
CaXcO/H90ks/zxBWrp7u+MGGac3fOV+j9srdVyu+gjqsGj8Lsp3NBO+r+zc9FshO
FXZQfGIdAL4r3GkjPmIjvEIqY4Pu4EV/wdmxxK19pISBog3LbHqyD+3gmNXwF7/P
GdTUJkdtW1zEkv2YbUZMByrIxpYzDzU9tKdJY/nPw0AIZoK7eBxq/3E7V9wl3lkf
ps3lq8m2qTLUkv5ZpNBXjOnOSmiZnJ9UQ1aT4EGvaxOJ/PvjaWMJl22Qdl9vMcny
idGnM141g/m4SwTC5tVGB3dlJjOVwsQ8DLoh3vtWEQM0toceIBZK+dLonsCxKdWm
zWPspATLsZkGyTSJXRLPdIi3/Wo3N0JLoA80J/VRbhdGit2+9ECA3hi4bdk45iEF
0zb/l12PISjJenHHvdw1DhLU3oQL0uOKStgP+cIHqtaLSvDtrOsy7k6G9Bif2x4/
FnJMQrUGLKvIRafzrnIwlZF07+B2AGZ3Ymd9U6nO6k9RAT97q5/zuovCESm6135T
2v0kH+Da9aolabqPHS0ff6Xj7FVrn7emvUVQtGBKfwKTAK44sllbIf97/0+rKStw
zJAFtleA6xrBVgxUoLHqX/M80+I3CA/HA1i3ef6NAYdGH64x6xwm4KUN+kyzK1BE
UPAAu9Xipg+56c6+vd3bp/cHI1N/rlGAIVoTyRbSe+eoNhXtWwFi3bRokjg77B1h
U6a2X1lTXZezBFUTHqHbNab/mMMfH24NWQg4FVxZdsl9kywJ+WwHqT5gIGn4UAzZ
qCfn/nfJKMILNMzWGq3vJtwEzvtLTfl2NCSxnhfetGdfc8VH/PSYvsm8HexnwMMS
jMvVoKNlxJzBgkgM6tWYZaYD6pBEzTHKWKghB82zB5ghmSn6asCD3Hvc9M2rWtYF
r1HNf4mrkQrwrCoDcvYxx65eSjySKgTQbuSouNC7ckAe1jIxQbMKAj6TIywcLDdg
m327MUU2U6Be4WNFxLaSfYo7wfp1WApyWfRWjlFHitM867GXqf4sxvdezLhRAcBi
P0/Km7F29YMkLus6Suj2MTOyKjw+hamABIHJNYOTUMyuIsclv3fqnXC/GE/MrZ1v
AqPwcEcMOCSLJal4XUR+hybG0PdofU9kn440k6L2Og0Oo23uzSzbTueGoUeYEgT1
332TmZ8TDljeDVNzn3ZyCOc1XszxeEmDTrtdmFLaLId3juhYulsXtQOhvCnGJlJ9
cOY1te1bur7YrcI0xb4FeIrteYAGKCPpCcA74QtTrgX0tBcSp72Vzl5+mr+Pl/Jp
h7jqbOtPqbLSgyabiLxgkAG44coLTkeZyJQSyf+zu1P4mVQ/KdpgePZtcgebytr3
4nwn/hUyhc1uR6+s1KVeaUc6VszxzpvJneqAQLZfoMMtnEWlSXdk21hW+aNJI86M
5rHMdkXhY2AOGG0RYIHbzO+OYvY2Lsok5pOb6QKvhlspmxztlpvk9PdtMm6VsRxg
O4oU1bmK5aFZgF9g3rp01OkIwPmHlooeyM2UJiT7MpRy8HVwQtnBlRfvxo4Akqmu
soRoo4pqhLVEU0EVKV2UYntnj8L4eI4FwS1d3NV0sLNo5SHnphaE8P2GiCqahnuI
SHjgTZcIE8u7NoL6YwANOkXY3iM5MPJrOO5AEVDDH44McWm+SAZ9+YUss41fLpZC
+JMYqDzPm032zpuPSr9mGTp9ArKP0ASWrbO9szoND2VPY6rCoNYZ5C2LfXAwCJf/
92hoaKAjvSqC+Z4yIozCrQ/wIG+i4kW+6atZX6tFrnGHzCSl4o4oqLGJAJuYQrFG
yTRcdaNvmjtTvyF3cCW4ROs1EmYIAAPUi/LZPUaR7tkNWGMWDJJmYdIK/wsGReiL
Yl0mU2Sokkr+8tXK+3ii2nNwx/nmsP02qQr32ylzsDAsmmsGYyN0EpkufCsQ5c0N
sNl+hmQyG44d38GgNg4+u4BHGMweQgXMaO8wmZIcdPKCuT5IhC3zIXDvSRltkKZR
1ApwMgGRl5VDGZmLzMzXMBvpupzwsxklEGtQ2NtvVcOIP/dI2op1+l0W+ROm+IJp
Y98WPmZn9KOY4jvSWwxs6XYbs+jePblNQa/RoqfJsKUbmaXLI039XUXGJRwF0IYN
xn1N57/+Hp/r8X7+4T8FovMghfeStDblgd68cxI5bRCZj6auxkl3HFHgQJHU5U76
fHYK7r6wqRNHQhh9WM62x7xGzan1ULLgyyWWIIORYJ9K4e6wm4hBLElcB7+A2Le3
pWqoh2fszsVbPgFobUBLAVrkZ8Hs9YnsjwVwsSq7QfDWWxyKvSG1MtGSbVLGtqUI
/xLWoUW7qT8y5w1QsYLx5xjzjm1P/x46VLkfXhdlNvfP2a8d1+J6TFNAzQ3q58Rh
cugPRG1LxDCCbkpWm6CpdYgyv7LDc8cLwncJsYuLCMJqGzSMrMxtnKnm4ntxQ7X/
PdXdisbbL5/FCSD5NS4HVTIjOd5ChDZzMbXV1da9EsK1VXw6f9UJvPun9hxxelBq
f8+SEtvoxlJDYhl/CFwSPKFuOnhGE+jwj0hsU/3BD/e/wMr3ghAA0Lk7pPN+gd5d
2pKJGYC2iOoSTrYt2PZGUT9jVeDJoLb5RBKcLIRxB+Hvp4/gMCElr/dltr/EVvl/
9IHyLskmH2kY/1XRs8JwV6GOkW07RegxrzaXYvvZUtN85sqtpu0wW8+E71s+8FcF
Ifwhwj749HgCw+Thk6U+wp2fYDSf3fCnvHMgI7lXW4a6JzQ/MFAcBv8DWCYmi9KV
ElqEjC0RYbhomgFP3PR/SdhLCGzWvdzO8UBweDCD1BthwAGmbnIiDls6zg2wsEJB
ebtkz5dtCo7QAoMIbPkmUk5my5gBYls/dZy79QImFxVsRMgKAjP02/+ZNZ3KgcmL
rfkyhgYdDB2vo6ELQav3vqXUAhhw/2wtd8aWre0/yAKYJhc2zOCyVpiJ9b6+RgPD
4kNmnhC4hTIguar3O3AEGgsRcimD/k5FyElpLI5c6t9yWzusSrgjoqcvhJG0s9EK
7K4cJzEXMjjI0gVL41Rg/pULrltXXCOtEe7HNAxie8vHVvcXKKmYkxC2THvKk+3H
93OM1PCRAjSWeGML1pS+/iVfU+1g4Fp43cWNlMJ0Kr5cJOr1kv+FvS4mxI1c/4ZZ
ZYgWT0qZstHm4vizZJ06P5Nuqyxjnt+GT+1jCGL8dYwM6/Nph7xGcd9Ol8TX3EJI
s4wuRjs1Q8CgeYzp51RRloYYMGeFYz4+lEyhoTjpwX8oCXPEoqhzitfYA/M7Gd0+
U0IUxGU7gqy6tANtyMY8Nfs8bHR+sMWrSXU5N5vo0VQ7+RMllHeNElnJQLD5I7o0
gHPy+aqY+g8SRDzm8zjygm2fengAyPkUReKZmlMW/pPbR6st4eX9a8fS+CzZDqZZ
vrm+VUqPb4Js2LEy0q4kDdXaI3aTyoeXybpkTgRRAAVTK/hTXhKwY+oslqmz+Ddb
Ns1fIAz/odES7RTCq9FxCpE5LLTSRrARW9P6ueormxGReHwrqjMR6vRPVzavjvRl
zQfcD4COGlYDJ/ZlO68DOHO52EbT6hIptSqqzJ/d12v447gkqIKv4NKEZLbekOVM
rMHh1dTb3nSv6Lfe8KEFVn7mOewDgZMN0QL0FqvoJxW5+9JATxZ395v/PDs0yRMl
6M8dUz5i2eKuXfnrFJRrSAI6XYkLCKcY9tMYwaeNZD1j/y9BxzGQZSs80nTXfzlE
0JkdtZLTPompNKRFIAQ7/L8wv1Rua4f5WiupyCB3N5//UJRca7o07intjRTef4xN
JDGixj5tUb6/jBXOs45sCkqIl+Nu8d6tu6bl6A59PE8iAv8hk1CfWksGKc5HfTbq
I9Ipz0J8amDUcDjkCmQ2iImIuIb2M3lU9Y9foBsXv/R0QwKj+QpN0eNzDOIM2yTp
CK6nuR32zuHSMbz0PL3H/ptzCWDH3eF3eZV07avpozJoadrfqO9ApYlPD0ttEqZ7
XxS60CzWe59BaBcU9O1b4JpClNIbHwHeJSPQisbZiIz+iw9Vjeq8v8iaCiViUMc7
vFSPiiq/6v92mp9chuHDzS0wDneHqGVwmngiqjp9XrJDp9CpLywvkmqIQW7cJjLp
9bKwSCW36S9h6+9FbmznvTRXhe4eeAvorz72FrJKKkSWYMhRekjPLw8B7lWgVqxz
FcLz7y2fd6AgiYifSQSC37KS3HmNMJOMROpmvKg4mLoAP9xxaOfkNj2UsO1vNvNF
eZ2guGhoJlwbQUnuDjxs6Zfi/BFbq3p6XjjcTFx5xzPCIgpk6qCzd8RUJaKrH2IP
A+eOIA2tYhmZFk3vtsM8t8yFZLt+tVMqdktSaOoHTQuOa5efkfi6vSwOnP7S5c3N
ZHMrapNFbVPAiP8EFBVOgNijx6BYplHoUpJuXqiyXLzHlxfreP1EOft377BkjdlR
G7hOcarfp3A7+qV7irjXvDwFb+BCd32qEz7hpisYmCF12S4L5a/f8eL5UVOZgjuj
dLyj0ia5qs4bBdCtJTbJCFPbeUNcTIKtggr8kEgxeItvpU0wDq/RXxU4R23Y9iWu
2ilgq5D2Oyccepp/8DSTOlQs9vo9Aq/xtsiEeKEzpHlFJGSYbT8WjqmIjK84J/M/
DU/6p/wiaci1sppLWF5SUY1WrNwwhJEf8xYB1FIAJQmwIIn9jX8oV28PFpOLfSWS
LMCdpBDuS8Er9g8ePXzIKypry3+CPGCjEnvGjiT7ss2vQw69u6V5lJ4HnX5n71sk
oOtVFoerCWsU4JaRlswPdXUFqqGezRnbyNEH+dlEBkn0R3YB4DgmUVK0zEqzo5kq
3NN+YznClSqzQvOZcZd15UNL5ZTEmLdOeQrRaOmUSetUrRYeOtisz+Uco24eX8sY
AzlGnBAP3967A4R2/AI++kUjCwKbHxm2pmNutSiO00bMqi5k9tD8GV59eygWTRDv
PzB42FGFJqTeE4PaqiOM8+jBWlhnR5SySr8zDdr19V7m0EZK16lHdJma0pbaHx6K
cKwoSqmbdx8Zzvqxz+FGnnqtYqvvD4VpHGGTx8Y+nYT43q2xZzi8lDJzv/B701KK
og4o/3vHAPv5oBCxD2irdec/EOPaxJZim293rexU2VY2xOF0prfS+Z0EmBwD3h3V
gUZfSp7ojrC4MRd08SWuaTtnZV0zycl0A3ZUfxAMz5Ch5jmb6/i6GSs7BPCzgtJk
9aVyumnaGOUKvZlumGrZd9W4aZRtybwPHLrpXGqZN6yH0QGZG48XB+JRMRq6/CVE
hgbZcb1k7VMk6GfN16ds1JGP5DKn3manbHwMLhZEWffF9eHPnMHK3Nd/A1BBflgp
tKoTSDc24sATL6CH8tykbmc0fS2ynfr4MZBlIz4C9jdMVezT24W7nkXeYgkIJ6hc
716/BJtERZccJCvNvWG88d28rVCDwZxJamGEMFD1Z/XRB23KMFvEZF7mThvWJev5
9u6odj10phI6JFO6GuV/XVsCk379bXJ4aP00Hx+7w377ea7KR4vdxkX6+XkOA+Y1
94RXBY/305FImodcy0elaYS2rHgRkKBUYW8bMgsyuzSolC3d6yParMcWtZm8b7kv
O4VXpUsuT28FwlFVf2FHIvadkvjhykC2+lCj12bY9ys1josQreyIZMzke6sBfUC4
jleDPyhLJG6fFf8pFpfI9GdX251mXXmdjFxPu7+MNQ3/2CTsyAyypWCym3J3zPTy
OZrStTF5c1l2S9A3o/Z5tdst3mLLflTxpB9J+mQa9lNbx+tjDBhk4x1562AIAtCu
FMnojr/pQZPiNRfxwczzMwHLjviPW5Nt2SbzEWursQly1VvVPfStpZyEPmIti4dU
hSZpfc22XEwf6vB3muuD7ek/mDe9pEAxW/A020wSA91xfKMO7y5pCvhHKaR+Btft
94vP5+1mz4G4Q3C3erZ4Y+TvCBzEmZ31Wn6slgW5bbdnknQ8NkoyhWJPD7KDSRSx
pW8jD9JWaLmHzlj6dTXvMpZjy7du4VuZamJ4zUBeTPh4JKRJCrwcCSYAeHeJGXvn
5c/FdtnBIYh+BDVbBQ5UmNqNgYU54lMRnNT5luRg5AP5P54IEc5IXxOQrsxhFB4q
G2EVXu4TiUGsMhU3T1IXy2pGzEmuhE6GHqTq/ufEN39vKtRldr8zbRee0zcrQgKv
nTyJ2XfRbwRBhsEvZTiOZ/0eBfHKrnPUkQRFmK/rOn94hzSLqpdfyOgHv37inIJa
cl48WxJ08JVSF7g6NTS7UMbjR1XGGlb6l9N7S34F2Qs4D0FqmnAn2zgz7RsY2Y+h
5tUNceyhluZbEDKiFcWiOnTbMkbLdjYCowA9aCjhN6JWZVggIJs5n48x0kcPgos3
OCN6Rg9Hy+HRIMiLsXzT/RiHvkqqs05oAgT3r8rLxBNiwAWcUozZMHf2iJvkZ2EH
CEyyWx5PhnOeMCfwCkoLtboraIOmubg+yT0xhknhuAIbj+8fPNdEBhJrOHjHvdmq
U3LQ0MW/v6G8fvcstTHIPIh1B8Bn2Z6egfK1Qmkz06GWkmoGipRP3qmvbgfwNFrK
y3z+y8GzkbATxByRUSrRN/MHT6TkW/Tpk7aOU+cCyeyuhnHpRzYC1/lZYPkbFbQ4
zRDVPujEkOYUpgKD6VL/Gv6Ld/oW+8CdVCDTGOxQk5D3+whVj5md6ZRhWdnOL4sz
dOG+J5zjIqxQLHzK9R4bA67t4f/51NDnjzUhfsljljaNNr5vIeq2XOrfpEIyDhVI
A4LVktEjaAOWuaK1DNNYbPFot/SeWtXpMNnnxtszMohRUYCcLmvyYxynAf9vV4TY
hIsk6MBbRJMcLHkQ8CGfdRaK8kt1zbeYHU6MjdLOgJiSHMDzpQ6pTyxk+tgnEmhZ
Y9DaFrd/i7wd25aUlWrvckluXFk47xl/PqUroGSB9p9XjTtDf+fwZyqgwCiLntm2
QMNp/0445AH8YH2bG97tL2DFxEqmbxqwez9nk4oZuSs3G+F7mLgbooF7r9/nhcPR
YyopLi4yitdUwmmWM2P5sMFFt2sBgFFKT3+piX893xjaGBm/1teZZZbspdtNwVS5
AVEsmR6ImCtn8qeto7Am1+Au85MzmO1iZqYkkq2478pcowSKEZVvrZKVTgvj9PEM
SmJKluzlnUWg9k+N79V7bV8vhUJqL1gh82OpJ7fV7AEfLIhGVkHbWVDQyAFnAOAI
go2ziY2Rx074JYO+bjXXJdRs9Xp/WVnFgRIgSbpfE1yCqqfJhkiMFoopYPjCs2qt
ireNgmiOm7vF2qjqtw2A6fZJ0yiCOo7fZQS7HU3HencWZLv4ulCUw6qP86+wUTfF
Wgk9vR+HwrBgeSFwwoMdF7dABUfknLNvuAc1g9WyS22WbFoCAbrm+RlUIcwqGYTm
BzbXIGBlkcl5e68oYMlGdGOwt+eYnruZcg38PWmYfasOOmC6O5Zi4jji6n/VkPqP
3JgeWLw5hj83Fbz7hw3gN6yylNFb0XlFeAm4nmal34C7KxqfyCS3HkY2N7qgj77l
4wv0N2uB+c1X5kwW6a0QiCSznmHBnwKX3YZlgp+uCFEE/iot/8nzucbfAIAp7o4P
A+Gr3TqumhsZeVHWbiB+NPaOAmmuSPGAVQj1c6g9VjuO+NPYg0vN/Izv0lqyuRtS
VVOCMsUyqZ7tPc8nzQtCSM1jv5m8XN7fm2ejElnAxdlLbOXAS16fsHRmHEbr2ZFa
g7jQY0unslK/+Awa6MpXi+El0oszjrLMbfhwaCtNYjpZes2Mf+0IspvFKmcBtXAf
PKlCB5CJ5z+DMtGlun5+7gvbYN3cBDPlJ9++O3jHMkUlhPpdjTc1AyLYZ7a4nj3P
iHD902w2ngM00P8tajo7AVdZvL2vtqj5WRQRyVm2uadiW9YQAKXf3dH3nqhyCiLK
HX5RvimZIrje9ALXIeX9pfN6c6UntgHmcy5Ruf++sGT527YTdcjkeUbp9PRNRYM9
xJVmEzOm2+wRhrCDrpXKm3rhfIgPgcXbczxSzbBvL50ucVFHXGV8DMNzte46gVwe
Nt5fmhbmwVpF6h2J3H1h5+117yzkbEWpQ/vnriW2m9k92hrcji8T7lNQ44sCJqkn
LdTYkrjKvaRXJ+wj7Zmb5rptCUCpXLc0y7IjvXk1c/N4zLGy+kWogboZ060cmLt2
j2NfFACTjIcTmOE1CA3HWUz08j49D0KNqym7xJ0E2Q30OmY+API/M3XInd43ZSDl
6TzMNaUBcgyxCw3LM3vic5xAbM7lChNypkadvbEEE63314P3WHbvFNlw2VniETdV
ohrwAKs1rAWVk9N1NhLBgbqRxZYD4Ej/Cduqeh3a5g4vf5p/p1oD1KA+zrcZzxhI
UBoiLXTVBoCi32vXuLNQXu4PKsEH1DhNhKer+oGwI0nyFpdUucQOzi3tby7+Bhjq
Duac74SxfLalO+G5phxMc1qIvVj/FRaywxdTJBuVZ396lYE53tYKzYWWnpQCESWI
MFL5JRMZIm5a8O9EXCC02umpEh6ffI52Nr2274v8DhQ2UsuniQOKtMaPg/c56VLw
acwDsG2ldTslADZPU1HvhccE09BsOsi4VBjn66U2WUx5O4sJEjVtEJhWWOyYSTDj
8PdA432+4y7fntPfYOskjhINLIOxKD4pTBN28lHTHHKEFdDPy4yIVWjbjb1hiA4a
lk10GC2Wp+8RvyZe+P0RTywQUfe33czbdAXekvdjWmdgHRiWbBwQpMwLSTq+abJm
/N0yM6W0RAL10qEUwpqDJ5+hBcY+dGeMo0LCieZJOvk4gQzb88P5fdB8//3SWDQ8
Wc+1A2/xfrIZ4gCYZVuxRAANd5ZX6NrWZvnqSRiUu0WDWMCKM2l/Xw0PROtz//Kg
xzIrZKj4rVNTx6+okrxZPfBl3srP8hC37RBdQ3St+KvdVeq9IEy8QwffZfuic+Mz
/uREAGB02b2KNdipY24Xt3eKgfKMHDds9bzcv+YkrksX9Tte0vgLDQvn6AsnMY5B
WQl5cS9BLuH1OScM6NdsjlODSpuEIERVURgF//Azzvf+pzxLQsoqMxmfDluxKNax
hwIe92tUQUuECLzpGMArQhkJp0fAbMB6COxu3jAUdOKUl7ir/mLiLmbjKLA21WDq
rRNEpGHZRCvm1JTRj0r7hH7zN9p+AzLKqj9Uv/dWYKtvFqejsSV1ajwk+4WSBVFM
iGfWmxN1s4IBQfEsgMzOJ7pFsg4L/wjuA7L42qSnM6fWttaXtV9GqheV/cuHI7Ss
vE9B3mvsK2qvdvHNNsVqcpeGxd+R9HZwGPpCYM3vVC06CIp5p4ttKEbsrPgSQ9e5
bJLVmqQs/fzhtg7ORMkFWzr+8BktRxW9WR09q9n6/ChI39DkjwYbpjiR8DzBl2CZ
jix9GGbVXSF4poWm+HpM6d8o8aJZVtDQFUqSQCO0SXNUsKbontN1EopROO1YbNGr
mAHp0EpCmIWws0HdpjWdVf8215YrATcLKnUtUywNKUG7DrLiFLGkO0iRFTZIm3pR
6eeLaUT6y29ZUPcEUcJYzMSxpOkVP+knqk/d5bXXxpYjU0iRSBJoSnIXVSXbYy0D
bVdxrSJ98p9hIXLTb8QxxPxagETmlqF8ogQTHDm4dtXW5UI9i0fWdLCeVMYpa+v1
quWP9DOIie38KGPKPk4rAivbb25t6FDMyIRoj5pFvXbJ8LowqykUcVYcv6g27trr
TmYmTNyKxLVfLRmdCmQ3s0Ut/gjQvgThx2OTs6+YBidUuhiKpqCMEiVb5c2SlW5B
Geib60bVF1GWm9mUo6Hsm14RI74AKG7ingsR87NgWIVZkT7Zt/rvmNlGaXzPW6Wv
xVvMQYupIdPAPYBkWiI8Ly6PLa+Sui71YIA4k7zktoUipptjI6zlrUTi6lYrZ6Oy
+xaCRj8txxBIoom/qoCKFU86kVVeEdao3OCRhueeJRRl26F6MXLcI81kmLF77eYZ
ZbjQ+IMfihbp4a7kVfdwYwWnKrAP7/DWJvRDPnilr5VtMwG5YgQAEJl0niYt9Oyp
UTka7ZwjIDJpk6dhA2EFxapg5VVBac0K4pCxE1+uUDNF7Maguq5gRNcnjhhkQI/a
MUU5Ob6xQ2roKrtG1pnMwmtLUy6d2PBF/amIGMZB+Kv26nvJ/i/OOJQAsvgJkQ1g
gkVRNLhN09aiGxNIDjiXLFuKdkebKdos32j5Ht08cZLaQpoub9qRfqrJOROJvbTO
ZKg0NKTzJd1aF7GvlrrQPqT5sbtaN/V+vpjpVJ4AUCzQV1rZCprQ36VOjo5LKV5d
QQBh75ZFeA39pw5Zf9pfaV29rMf56VQO2EESCCkgLEa8rrO66sNh/aOuTKocTylH
HPNLOG6newsFBM7dTb9q/yvdXHDXsar3ayIqeNyFzFioGLGxmK7/87uQh0Y/2iQ/
fMU9p/4imUQOIhhJvy8pWvezbzoYnh9eXD+ZN2Baoe7tm7hn69G6hypm3Yj+cXpA
aFHx+dusN3/vecW/fabgMs7dBSUuBj9+PwaW/YFws0zAPJPp5cNkUT/EZ914JFKY
MpEtd7J2stFJSSxkqlfqcb2g6CkyAYHovg28Va91Q4+D4EIujWUiT+c4zWvPjeFV
gHIDY1576AxGc80wcCyQ1q56ed3gLXzgS59iFRHJhLiszcLESRDBZtKK2LK7+4uH
hCSQcGEfi1dwh2Hsv3/Py+r+yCgefwCL9Ka27izw4FqbfC+7M3KGyZMGTGATU/0+
jsQPeF1cZEjSLZ6ImX/LsMmP+edQibLIJ2NH//nTZEf9ftG753HE3+5sCjZaIOr6
Z6144Lp1hELA0eo+dFYAOGaQkMXV1BQLExGhKuPOnRcvfslSZyXcwjYcWoXU8ehW
+xnfXCOp4YE+sZOysGXdJl6jFo/5DTQ2QtVjclNBO86uTDfHiB/MwI7vqlgijKeX
UE0+LOLLTLpYiTKirpIODTSZzAXAg6f2EZarsRsyBAzwu/nhdQ5tZ+GPU0yUy2Sb
J1UVhLoBNeHLkGCKXKFRkcQ+lFw4bBUatvOaWIlLMhbGxQ69Kl916U7RarRlgjC6
i5iAzo2/ejt/0UQdpGvYhEb9w2fsbeSRh6UxxHVGbjf4E+aE9lNBtaG5HMqGe8i4
TmTt9W4ay4ad/tTWh0ze48WJ8uuE/7+3p9ypdYqbYJ3cicSz+HPCIZewwQemqDsw
odn4KeytEAClwVTvOVktAR80aGvWjtlo5kFeUDAVfhfO6Xkv21UchE2iP1C6I1bU
2JbZIUdwcwrxniX2dn2FN+4j8sG8MjauWy/BwWNkJ3IbUZ3Y2+OK7gHnxaRncXKr
KwgYFYxnpQkXE9esU7osyWC8k0ksHEXAaE3Zgyes+sbdewBpUKtOPYzRYL6+w34D
hBUeLEQx14LnxYbJRgw1JdIIgeJmrdN2qs9r/RMQjntZkE5aciNj1mCIlQ9q29Nr
rVTSHvZANLFOlGOwnqrMOHlCm/O9JOWOymnKw450v7uVU5KxB5nJixT0NHu4PV+a
sl++/XX+vHkWFBHzQo0lR1KFJmCexrTf/Cuy4S4pyV5O1WynLLGfZGrGr7wYIkNm
gCsciYM2pDjVHjtbZpzNbFJh6HqG4hKyCEkeVnud8lzJSgPq36Ta0YeYN4A86lbx
/GycNs9j/jGBl3GwrWtZh+egdju66mUfgskB3BdQD/kPGV+TXHyVoYZ4AnBeoyAS
iIs+GH+jQb6VkYJkyADFQ46o/+0uLDS/ACZgseZwC45ObzlAQgsyCa/Q6ZRnbtIA
1Idfs+azh964P9rW2M7TmZxIQKkh/u36iRugwW3ZfH9s/clD0Cc/7v6aV/te86I0
SIcBZ7a8TfJ+0LiDmmAoS92ajYaiVbsvYmbh0ouCDzs3+AC4stZwo4/wznttBJgb
/6kaB6c2MJft2RPq73L3DaPpCYzyDqHnlVL6SFniUUHQkCQKHFjZRDgCA4Mf2tlm
cBlJVXSFINV8rn99SWlqLkzioVx9IyBwiQpC9PBPAXAieJUzqcz5v3pbD4hn5LHz
USjIW0qg54RdhGzEDARa3edmHQnHneHsPXEm1ZHBJqukoJ1eGtgcnz/QBnPyAtza
hkqk38rZ4C5WNzHl5YK92fNCuqFkD+FK/8P7jSuBWPNrwVg4hXMA6CvU3i/OgRsq
fMO4OKKCBYDoz8kug5MA2ZQWs7fmi4+xOjKhmquzmmimVnmCVEop9L/MhDr/Kbyh
d9v0nRrTCKLGBICCoaYxsUQpk83MW92r1f9H8Izsg1/cniDxPh5P2Hrd+W9ikrrZ
MtHjROBWUL7cpev3LChlp9wl/ph/zoWfpyl1qF/jJTCsyHWZsk95hZI0Kb8VNBKY
TyNXVyCJatithX2XO5Tdk9IERL7J78MXUPqoievQKLhKYDZJz0Xdt47I+DTOBYH9
VAE/SIi3XhxRUqaq+PaJLLNxDkO7FVlBw1OA2DjeBEkvUnG0G5PlgUiPHF3YDMmj
Z5Cr6Ll7CGQDc99LZ0MW+rq3+DOg6ox/g7Ox85ezyWtI+GWVSXBK3UdgRNXbC3Gq
jXGmqxpY62Xo86tpOHmC/6mv3AJxhvgGuBnLdYK/1vZSXLwnGHmcViRk7SYLcp3D
+jG7JzT+hLOyQrdJ5ZexsNSqzThxQpvuR4pPmhgtn3C/wZlDDHlt+8sZK0Tp6xqj
3e2BoIsZGAReXTL5hj5p1D96FkIFP9Y2WyklMafPGG4P16MgJvWa5e9cqjB2g/Fi
vsIFJ13l/+D1qMVzJFaoK2Q75dK2lG5AsYdEpXknOF1cyeFeVWMJPTwRC3j+i3Um
beKlna/Kft0Ea5qY5cW3RI8zobZoogLLR2zB4UQPsJBFdnB8Cmdig8hhnWXNop53
HQw+QuNQwW5UW2eVDzm6B88FVyCe5F+5RvyVD5SSxHgB9QbjOxVDr/cGwpmsjQ1L
A/TaYrJeBTtxSQFs3Kivgxotds5vC1LsUIVvgLoZ37EV3m6MXlyModp+/TecluoU
8/8z8Fsx5j7d1bOcUZ3xFQxuzcvVj/qS5NfmGDIY5N9iMK94oNHZCOQizB4jZ5I9
lMrGGY0iGTlmDsWdsNfuq0IRRI6UhpSs7hARt6aSIfOg78tmY34vh94oOXuwhq7K
+NpnFS4vHt5iEFUD5Ep1rLx7JBjWJ8hza0tOFwWB2h+Xl04quGsJwJNZH9WKp2Zr
VyRk1qDuTH4/irjqdrU6ZAZkmcWZiF2X5+Wye3Q7FSxZdZF2kZO4RzcmMcHhFBhR
R+LiXraoKiX93AEtMv8xnfOrPmue2/wiRhsPlKntH3bxE77tFrzKJhn8E8m76Pp0
WTU7PS0lEnxhDPqkxEpeme2fepKbgkMDVe2I3+8+28StYtOOYFdFDZZYEhKSFCJj
TjBAQcUXn+1DkH95ssUVdB3hNuX/R3WV1iCUnC0oAWBP8Jh8GRFX0WrQFxnE4AZW
M8mk+MMnzMsttAe28XhtQ6MB0YH0mk3HFJrM7U9yU12sQt1hySYtQ/zC3qq3UWH3
mwMHQfeRpABwpZ9gYKPWjWBjGI8RnQMJ0R2whyqR0yEu+Nbu09EbHIpZ0TdSgi7x
Tsh5VDlR6p7/6DcHND3RWXiasstAH2zfB796TbVZwOGcUhWf0PKWkPr7P0e3MlBP
daOQCOocNB61x3M2725V5cZG/xU/K3HCu+qaPLSEtTwforn6PPJ6gBcNdcqrGjlM
9YKAlXeiewaVwSORkl5pRLKYz3G+z3eV9jMNhRHfUDzj9oHIWBOvNr2JHITxWGCl
/oPG7LlfKyOHNomBdytfKHkk+u1qxbYKTBj9zffD/+SVJX2gA+HNnHlckOaPeAwc
eDCywh0yAYSBuoF5djB5j+0AaY7SyGcrwwCIlG0Ims64bZGes0s+WnOLTFrHXO/K
6/qH3p4Id/K98JBLY0OAGvuU3UlQG0dvLvc+onCy7haNVQZ8pTPEwDGzpXcL91qp
9o4DDzaaODGEoW0JVliN+1zabGqPMN21Mh/RLcZsbsIBzyKGvL2mrnmqxuNImpI+
ZsfgHzyOWJVX6/dj2N3s7xTkUWauRLUYRdv8Z2AJXsluRqsMFribGq2aFvJkG64k
mbsn21K9b2hUKIPLabdEHM0j/ihbggcI4Fr0X+vzp7V/rPSsbHmqSobaNNQOaxdN
c9av///Hy1zJ6gJtwCbI7vvTZ43Dxqt0kT3mPN+jwk4ZkB30kwHZxF0Wutq+/MEc
w2LM2rD7TnbHHp0ZQ6w0w4I5YmR9A4Yt+5tL7xeMRwrs6GOKXSnVOhumXh8B55p1
XrcITwXC72syC6W046yZT8L84pVrnx5Fe52B6SKsFaytviVSMbFTJf0csvogm0g8
78ALhGRjBDpVzVwfA4o3fqhFuHD3JXWrcWPr9mMZdTBn1TCHNgAG/93v9JCJhSMz
Z7wUXty6A8H3wxSPKpai7HNqwPlwEedMO5DXMTRwrgtnSiUvPLOJBIDlLCz2D/3l
gllt2GQ+dKUWxakXiLhzr7o7KmV4rIib8xqNR9ASAM33H8o23EYb7+tO/XUaLFwf
AZ930rPP6Hx2bNclANE9McYmmhmU5HY/8mJyU82yNJqutq0TKCLNTSJ35hfh1EMH
BmIUIdx9+9VmxSwsTn2rZGsESDaczpXKXW3vqwDtEiXAHhM7ENla8C+VkmACHVTa
3i/lo2XYORIu0pwM2Vj1aYk3n38yDw42gebRprJTLe/GO/pTB4ULoukx4KW9fEbW
4920bThxtnwjac0IuJ5xVg4x/4mXIGUFOgIdz+WmXXmcKmrImTIzRZTzSCGxwEUr
IEtVDWlAvQr4i2xvNS7TsqRiZ9QhHMt+HrGR8Rcy/dMs3NoqeWKC3z1lPOD/pg/R
I22xDbabiJn6u96WqTGdyqlO3KnL9hhdpZATvI596bAjqAvbPdrO4X8sSdeUWTog
+B3aLPg8fGtn193F1zPUMak/AXal0EB0UFQzYfYdUSoqmkEDdwdmBQEll/oTIvZf
cJlK4YU5AZHcynp6OQtxtaedVIAit6x2GRbl8JKlV2wI6yUUGcPlMuCnoQ0UCSfh
i5O4Ub2VtSapR8AVNlxxXlCU55hA8aTyyhvbqVPSGDLTYeA1AqV3L33QJaNon6+5
hagLRlmtzcGub97s6y4MHbPL/YWX0ng0a+UHw9GyUYodz20zGm8PIuA+oN1w4R15
rNWq44Y8GJPSUQXAl165yd+rbbehOX0UOE9+Nr6r2g76sjcvrKy52/Z7ZeIAZad5
qZTi/8h8Zk2M9BbOUrO0q0Jwwe2LJpKAb+54YCDHKyC5siv1QUzfiwVXdPcxphUe
QUbs5mOl1Fei2X+gJLhugBd8PrQteSqN/7cuRl8vNUDyJuMuFX0F7lgxOf5KojrY
uMYbVadDE4rbO23wGF+2CYoZ1p/8aPld2F0W7d/mla762D8vHn2OfNhWnngSUrZ2
SfQfaFHup0QcXqVyIfgVB3C6nSN/HlCNU3OiXJtrcLzIYgDUl2un2DpSUo/rK5BH
f4LBB1wy6nNnV5xSbk6BSZfYAxWA6eUFruBFr9RRFfM4cHPjoc/hjk2kn2KQu9UV
esbJM453YDIjzv5usVn74JN6kLgs82m8zHu2PmydASLuBjY1cGLkcgpKYDP0GCcI
46uau0H59aUawALFihqBlyD5Rk/XN+2ynwBVjmz53v+9jcb9PaOU6NvlDA0nQdoE
hXWK6lfH9qlkDd4CpVR7gpEG7eGujzmfXGrGu/rq0H0RzzGziTyzIR4XudMBcuwb
XS+lVSWsJ1DIq40G0zCnzYJO2nUGw2wFJFTRyD78nziJ/oAE11eh5TWrYPgLtvyI
XE3mHRFRVRbbcCLMAcopktaP5jUMkgBgSHA6xuuDdWr/obXuS+Z1beDxZ21qzcHM
CaoeSl1KhTf1GchENT47ThQp22QSyTjK3zy63m1oiOQOSiDLvz+E9/h8dBbFkk/Q
WVp7a7p7NqsPu21P23HUPh77hQKPwFLBOhq8qTCyYFA7NRkJD7e/1Mo1Z62aMGck
9MJaqulS4PZkdkNM4OQc8t6QGuq+tWx4KkC/nBfc7NdJ+7GAJ/9xigsc7YR2Jb3y
E9czjfRJIb1JnmnsU+CW2tbLJxxzdWqTJRaycf9MqLpPi7IZAhO9SHjJ4CpHDllK
2gKzjajMAa2ZVe2WPLOtIAJs2n+6aktlpqpwaH3fQ0e8EtcFbSLH6N/cF57VeMJS
+hMrIoYfzhJrodCrPbYIonSbY5YUD7MGou5rMwXRGdoTWHFDM6Hk4RHTDASdnYdV
U6smbOLsBfElPO7jTWOy5ZTMOGEBGTgpBFMCGdh9T4mzFS4iE7xjTgvksrjos+Bm
yjD26brYNBeaskDTxVS0qUPATehSmACwgCqZVxZp9Rtrf8Jza8tRz1FcWUJ3IUFb
E05sfyIMbtyj1pxTp3FbRjLGCgqgBCEs4SxtDi/P2cs/FPweu4/Fi68kG5xOT6Vo
6xSPN6m08D2mQ8FBzhPcV5Zpov4Q5xC+sSoTBd+JVKWuLnlmnVk3HwshCin7y8U1
ke8rg3Hn2bCBrfOZXxp+rGlTkifL1zPIEp0aRvnIZ8qWVMEPZe2PA2jIuW8ogOqo
ozinmKvohoEFPJrXrCA2i9aQgdJTkW/ISqJwNESdyBkBztTf0MLGVW+ffbQ6e4UB
pxq7VdMjNavILb3HLWLmdyvXZ/0jXgJS3NmkgTR0kphAS4ivefdWB6Kg59eRLg0h
POz1VC+CGZ3QG6SIrqr6KpCNA+EXYlxQXtfOSjCjdzix0CDG3hu4ofsXeueR4G95
LTvOFcGyHB0TscHiWsDYelttdn6HLAjyG++FbCEgxUCaDCSw+2kdQEhAEW0QeU4U
etC17+GeiGl1Cr80jZdJONvb3HCuzJkD9d0QYMj5E86PK/KXdOjQ4QnlJyHIX2wV
/UxMciAOpoQZKgonnZPAUBukVCGsuCEEuU72E81/FmxP6Vfxiq8E8qqR4HkzJyF4
4Jxh+I0B6zdBV15yS7mqxcpMzRGLxUT0aL5UdooyOC7cyJMz9tnD//ZjZMLvPXku
3BowBI7T/BbTQGKVTLpzlyFl4e/eh2a8qZBiCeUwODakSKDq24MWbcAgvwX575lH
BxW/kLjGCHiZxT+okYiABoSftuRzDCsVDhN4AFTFkD6r+F13uR1IpJFgNT+c8Tq0
DiJ5Krp15CkLukTpzOvExkZNp8F4nfAkzWsaex59l5onT0BOawLACNDF76D93yEV
87lrFqGQeAcDPYtiybLAR91I9DTD6dfsSlXcT62etmMXdcn3oUtYgorAN1JnmzMl
LzSnFUguMF+r9WqlzmN+jxombVEXLT0iClxNhfoR5VqguQzNmh39H8gJOHNBCgCz
YDE26Wg07c1JAw0m699P8nIOPMWlNR16UVNJzrp01QZra5LyZW+eW11V0ZK0QJ8x
wSahLJH9nxl1oprqygXNXMNbb+aXzBgzPKCmbLZPhBx31bT3I+CfT2xUsAklRlfy
w6RwMIn57iLsWS5TEWLqdEnJ+XU2UycniGuWwxs7CbYkjqPL5JkT75+n2e/XeqEB
PwdC7cgtmgB8mzK39ElTkZudaulfKYQgFwbBoq274eFcQ1Hft1p8ATMsValB+Qr5
YFL391XQIPmVCTIq4BpC0zPlRoDtKw4ebOMUH4wmPoi8eKzKo/dpUKWXJO4iSEmw
h2INQJ39fsr6K09r91vQ/8EOksrESk/pgms+j4W1i+2o62jYNB4u48bazn9PRsi4
H3vnfoNWO2GngZG6A8cnPkQOvfi06E84pRE06naBBCtUX5JaT12YzmAKIPMUbU5A
/uLUPf4FfEqxYU8BhLJ/zALbQjUfLcnwDEuuJIeO38a6bvl4H4fnxez4trGG8tDo
3fMVopvO7msHdkpLDLOayrXv2iUZL76p7oYgm4yFuxzhVSGnLDzssTqlyL6KOSYR
vqhJCQpW65cC6HQW42WEeU1jLXIFPyxbSbN9T9QV9cz7NY1pBg9uTvBGwGU9if6C
PV8DLyjIk/V+zjaWXvzwK7BKuy/PQwnpm4JRzKV+BsZNLmtCcdooFeKMsAmzD1wu
yWDkTK27opO8zXAhmx8IvR1o+ipJykkiultyowUbGdibLuehTGG7lVy3B9wSVFd0
4vvPJZnPlHZlImbkfHNwWu7UvdlH4NjPSB/D15azc4K+1ML7JCNjUY+7dXpY/OsE
o/iP4JwuRy0cRN3tYMAAdbs6V1v4gLvIWnyZsGJfOA6qMZj+TXlSWJ4xwiqfVmq4
ROnjAXVb4t6xeCb6y/WeDGcqF16tTea6UlACweFWCF3APpvCzCPN3t+AmxbdWvLf
8kb93jwWADwAY9hup+o/wuYtuycFscub69HDOg+yd5p+z4lIQWoeNQpXuQ0mPkP1
LMftFXADkiZec6wnfsXVya6n2+YjzwvVP4PuYdIB7RYRH/6mjBWiRNgI3/dznTT1
kUjWVC7yOjm+LElDr/w5ocf97Cl0P8wg2XnhncyC4ws0PZuXVwWqTFM/ptaQGNWp
wDtzk2Q18Tpd07PhD7NZwPPw9n19zrOSlzZ2vbBvReMTPZpOH9fnJfyULzUJ6/eN
VPT227eWt78Qz/WQadcUSdW2ipGJYntPEI2As4N1nl6eG6GN2Vn81d80Ul8RYQfe
EKlqyBL60Ud17FMVFw/Va+CGLnB128VxiQMnho8Cwm85XoHl1V9BHwZJXiK8ANvD
SI/vKRHtNfTyWbhbVoSkcd3sACS3i+N+5Mc53veOO4Qj4xvY5eKTepC2hhEFU8CQ
mp5ZWGuvwZ5pMbmNzLNVHFzaoRtZRfvTzxRp0/WdgW0WQ+mfoDy+BRi6n9VAJMmL
DnPsaM1pS49n8VVSNqlSfAejA159fCCZHVvNeMf2k5AadM/WA0xM5l84K2zCEgwR
TjNTeDIqxTiKBH1yZa9KJjd4Vx/SxzT1EW7wyCMXysHF+a6ecwTXo9HIB+KvwSo9
5CTYMfhjHFpQnkgfNKaLhABXw85dUGks2WybNOzR9bm6UiZdRLdnroLlceHadLX1
kfXVQr5rvFcz7RLE5Tta/vQt9Rmna+FPfgsUPrv/USGup53O3VxG3CYuLXGHC5nP
PLA8I/MkQ7akIzsYTj8NZchVzKc2n8kCQSyCbBKEA6h+O8BdJxgJxu2h+90ss4o7
R1bggbN7NrILNuDGDNQi1l9ZddEkK7Nxa/fKAquJvGfuicM7rj8jakbuyswWIkIJ
D7/8edLzntOSoTBN3Y9U63hypZiwFMe66lcxQXIsQVpDjwvCFwGU2XaDVPdWnYQ/
4ZzR6iB00MHf8jYlstg9YeITxf+0fUMnmluBss7p6KHQ+zSq+GDI/QaeFwKAOtgH
zuaL0nrRbp98CaXCvRTM2hHZc3v46yn1ZQrNSvUKTkLjtcxJvGRqMHur+6809HfT
XuVc+Kg6yLw+iczGDr2GV7NDX397jUYvzGqAOz/ol4M4kpOf0DSdr8KSSA0OQb7S
ppEHxlb9V1XaWOU5P8idDZhFxUSHt+4+12vUrt3SjzrhC8yybyY0JeyI9Z9EGYG8
GmThpR8a6hUkkQ+XlBk7ria0/kCywqu7pfSVDfK3bQSxphE89hTXDM+XiWWxV1w7
oq+vpkxm57z0xx3DM91CcAFtnjihqY0BPTpmQI7bzVb46xf2qb99n/tS62EUaMQL
My+Rco0fRak6J2P/gRw5dRSLA26j83mgyIMDb4DjDop8hcGUY6U+S1sm4JJDes81
oUi/3l+/X7TvH698VKxnXmMFVRV8Tgw3lhCv52MOVtgu24zamzaC23cxbKwDFiix
wZ6IGoWsxm3OzIgFPtTWi1B66mwnBeZP7V0vREXX8oN/a2iuCZQfsM+n7EyvbmH7
9VQ9oqDjI25wflCuAoQLDN8jr1xtRAlhIeIjHLKT7w9pNnWnGu419yl9huC4qjre
DOupACbTDpZdUNidK4A9tlJbURdyWygUM0ltYw7vKIk6UoTfUnbLFiT3EhrV9EZk
yMgAdl9VFTOT9QWf4kdMMNt7IsGSVXfSSkZ8wp5agYnYLtfXMCcBU47ofEtuDheC
FYtGUJbLofKd2iqUYvT4VOXgHsyT2tlfjWQ3/9M3Km3RhotnhLZlR5rToqmAzGcJ
tkZ2dPt7HPG7kCiL3qigPCIxVrEf/Q00AU4KiaeCGR/mwsOHpeuqlUHm115RhMjj
67e9s+/pQEJFi/R1W0IrJckjU9qX0w+NvZljoFParOe5IZGwPnAlwTnp/fhBc+bv
+gXyRmMsa64H6bOooUFXez8bxCgndzv/XVfqvLYvPFwoNs7OcGW4+++xF2TaRTrL
2ee3UFhKHLQL6FZUB296LpiNI3Y95Qj9C64D7MFZP6fo7T7bUHdCdqTV9gipUZ8x
HqeAbZXgHLW2rvv/ogGDOJeYIx5hogPlAbmFN9vNrwM8dNRhnM43WxsOPDVOk5BN
AUG7g/DOwGlda3dQkSCXLOL37ZiAO4NIJdo79kMxDaJfM/IYM+/Rz1l2YvGdWBKa
Eubk/xoqQSzCDVwyJ+ioMlH89A/1ARaoAA1GP2uxHlGxAIvynUvgFmxhYQEzI7y1
mCAwPXg4TNvlAOQJGnyF4c/3KH2Oiyu6AvJzdOeIrpDZ5P0TYCLNcWg+MZ+TV0o+
QMcFdceIcIDo1PAAT6qiHMotlZ3uM/1V/ZLHvVSgb86u+fYZb+mZNXODpiGQHOtB
tWiJctQWpf1Sxs2rZsVmtaLpHXU0byi5w9VEEfnHS2LjA5YICA8t1Ryi2rWUst5n
Wdtp7MRTp2lH869JlfH7nKyRYl978/atL6LMjIH1z2mgJTvGJH0USawEZdYvR+pw
OCbmNb0jeu6PLyCwbS4+BqyQAdZO0KL649toxSBfZuwgaReW5UOYBFmEl4B4HqO/
Eo8M0QWP6hwK4xDCidnI8Eieaew6BYWgiX7z4XDS2bE7VfckmiumjFMndTsxPk/X
fL6hmhibWaPLSiDA9UKbhVE3rRHyozJGouAuq7YlAhbB6sP4JLEWJodDIzfMYm7K
nXGP7K+sO+kfil7TarrbAQI1+Tidpp0J7INKup8Suh+SYuxCBw6NYE1i/J2HCY+C
UP8KeYuZdC8BZyU0IWFL04TwgrJorf43aMzsv7gSpxIysOj+zvTKyN0SLuDba1Xz
j9H/BboSOuW/u/Cn4WwVaEs4xjSNA6tpcdVYDTphd+X5bRIWj/5BT1beRwrQ5aP3
uMHtEGuTnjrqfg8WF/lzT+neRxH2kF+x+n2D35xijZbq34Iwqt8IOkhLLutfkbVL
mx5gr/51IGyo77tnwU927Ft80eF8bxtGdKD0TafeEbNy0sc+Gp3wbB8PDjeoLM0i
Hx6KnplK4uJaknMOpYkVr4emX4wz1mPIvVo+GOIli356CcqiSSfXDbcf4rSt10Uz
nzuuIn9SiC7MFOLjdT/xcJM0QS4Hk0GvzRkfJK2eWshxOL7UNeMWSKz6uFkJ8uVW
rIdZpqLSJLAFfV57NHhgRMf61k3FWtQElNsmHotO758zkdaDtRxHLwJKC4Tl8prW
6xgFafB36QCVxvneuKE7HbBTLNUj8YO4I3AClz2uPJoPaCgr/4iMFsnyKr2HLELL
/343sryviaJ6Iy1oxzw6Zh29nI60YJsyr2J4tD68ge9A9qqJhVeDVK6142+DRyRm
AJ0NQ4T79+dTtDpIKHzjyR9jZGYr6vOl3cdx+gD4gpLxIKc/lt/yZH4urVHqmqGx
/xRXn55lG428kCqMVwIrMQeQ0bBFY1/5IoEmYv+zQYUJDvm7/aiITyMbnaWjMWel
9cShcOBkANo4nBOtCu183n1alOV/dP8wN/w6dzyz4BMweVjhOZZF+YyTeOOrSHFb
aDeHkmPXFAsiKRBEeRTh4H9NloZlOJ9Sg5He9fX1GymUQ/vUJde59+r6ljQCU8+D
p83GWrCnukEQ56WIryQPzYGVcc/LZMltzuwqVYCzPKbKDnXVcDxDoylDY7ODa2U7
KAlE8AY6gfuwbGeNXXJC1H4EqNLgvcFKLRbVkiBsLCHZFfxGt7LGLLEAld4eAt+A
28XzqU2D/9l83Kk6VuqdoAC5DLkAh1Xs2P1rjbjlJwPkm2kWjIPoffnNwJ0erOtU
zEdBjLRxTf+Ix6lA5Kl9uW3PbNYCkS6ldcZ8lPJEjvwN2dnawTZj2U5xi5y0Ay3K
Hz/imsDnvOGSamGPdmdl3yk8eoVTuO8QVyc7FDRku4E/Nu3LgnrSEpT11Xq8UDrz
cX6SIJuli2MJY64BqvgJQpm8IAYcZPaVL7pbLquavEx7vqBurrQKzt0yh+DKYjhm
kku03H7qZnFkiQgmSDnsiXQG5xHACflOpk//racDrvTm6EiFqnWdzSnmsG0u8kJT
w78w9uxJcxED4aVGR+TQpmoEk/XE2Uj7HaPIPNA/vBq41nNvBB88IAju50g+auVo
SbulT0xUDlKE63kKWJlEVYDHpl0QT6gHSYtsx/p8Ik2DFZoO0n/PVoT7KSDMAppQ
c62RE4HHGr7kDGKRvAa/hnwsUB91HvBnE01lU839EnWWivJX7v5BwSaME/GNChY+
FPm4njMcilmB4lsBEMw387E6e0QHJrVmoy1WhhE9JfPrFYfgTMFBtq7xKBDV5jCE
L1TzpY44+/xvcXuP+ViP6eLiFWJbdbDVJo7FQmjgy1KqmTpf2HOXhg3KqR8LrbqQ
8rCN4+Iv9HszcQxyOUZbc/N1qLq2irBezIUXlLXPrALLyO+UJCSQc1DW7q7xvMeQ
THWvrfcDGGeKNMog0OR8vVUOtv9CcnodxiPnY4KUjnraLZreQ7nzi1YRxiiHw3+A
HvVmazVQ2iJbo9V8jdBmnWH+jxIECA3YYYtwW7ErStrrAARbjxHjBrxa2n7sRkaF
ZawyLCjznprdWLx310M6Fj0DyYZSublHZ4lVjuaUKzSd74jU6jdMLl/K3cCOPcmx
dGyiMvrG5+kzRFkT4C/OnbuqHNMICIoiJRi7D53CeojFJInqBwD8aSws/uy3cAPx
ceDqof8jwSmMcw7OSgRzEjW4Szk4f/4Wpay1i7UmtLblukCetNLpp/d+QztABjms
JN+hgRL45YM84OcZXaurNRzftSys5khSNcu2MZDAMZW+kGgcW+zWd7r/9dphWsra
C6MYa844e450kcK/d63v8BFRy2vtb3BXEceQv6grXIM5S2J9/4ls/wFhm9FmhImv
pNqqG0IV4j6ksEs4N8Qzu+EOAO7LIVBaRqXHO/umQf24qOOW3eABICWintDXnNhK
+n38pHSPNhQ7FFrWW0IfEKggwaoy6v9wqkUvps/tWvmahQp6THAos6XbC1A35Qe6
AhVWDx+6lJWx7IFbfd4V+GAhrO5ZhrhA71q1sdsY4P5ucQzSnEMeqQMQEz0+ZRVM
y/tDlrUNQgEG/WiJGG01WCCj5dOaXmLYTDTW3Mqkpzh/wFbvkF+5kYEO18cIeOTB
CYvEmA0mKExgTSEc5g0pootJRCQwBnQb6S5PfK7pwYGhVM5OsfdcjZk3nc9ds8MH
8TO65eIqYlwnz9Jhl+RSDepdR6Fz1VYDG8/KWbj7gyObJnfgF6YTo9s3//AHkl+R
9BtJCwJlqwALURly2J2jvrXxCRU3D4uB3QJALcoga6WrG7gy69824bwmkZepWmWH
sWVFH10RNCB+hbWujIAJJ8BkdsKfbwc3v8hZDcptAUfK7oP6eVsCQIB809TcjBCn
AaKt3mi8j1SMiTZunGkcn3gDgsxl1tR/ObwwjqZLlhJaRpj2RV4NE9/PNcabcJCM
YOsSv10vVb7G9KyD+2QTN9JCSWgsypH7m1MQaSN+qVqMgs3jCPqmzB870KIO+63I
adEK1d75otVkTovzocSrDBI2d3alifCahjexm8wLHj7AnTxVpzAz0Wl901OEpa43
TSyE2Qcvk3JxD+lfFgh7TFVqUQNlztvkErk29Lq/akOLQTWODIScgz7JkpAssVx8
NDdBsLoAaTcC5MhYyxRnCdQsRu7L2t8Sv9XMGEEqta8ucu//ksE1Wnu8VSY40z1D
MG+1ORrqM19Ftaikyb1mHHBbANcBB/iXgNUslsxlZPe65DG57WkTb0an2/hPOWw6
GwJuwSiaOQdFkjzXse/mGePFYbr7AKqR9pmzpXXAOkBOfKBTjpiSRt5T0pIiD6n9
PfFpVp5DW8pKfZ0K0htBIrc+YNW1tOQ2tw1ae7dKLHLldq0S62XbgnDm0Ik0btJE
ez75jzR7dB98YubySwsw5DH0eOTpT50SsEP6nB4eUYYhMKezEhMgBO4/Bw+OIzUl
8+ovAKg/E4rRf9ZJnpMa1l2Z1m5qW9e6pbj6tOJ+aEeECmWIMa89oV2iij3G3561
Z7BdvpG7lue9rIqLQRQyMZelSQ44aoptjz8LcRFVkYXK5McqdHal9IXA3tMggJoc
AShREABLHjs+GQHOLaZ9UMWTZ/9f/fv8uemhRT111Bz9sFhNroVrJ4hBUSwWdMlf
DOKf1JGLOcU7Te7MF/4ORIfKOIo0vHEryqa7AkP5Ub1FYQiU1LZkuhB21qP0erWE
wxMVaBlQc8DzCBJ4kvysDevm0FyKFjUKEj3h/nAcB1ye3mZKkgrtbvtN3t/AUzch
pQ7jke1QTPXYVQi5DkwNDqsf1OHtMTRb9mm4GdiwK6mLnEAgNLpkox1/01ooaBvL
E9h4EwuseeXyMP2KphP4uvelRTNuO1gaGyzIx5FmN6z7Vlr6TAJfHxwmnOZCpKzY
xrtb+cnkLIgymFbbUm5L7pQYbGSnZLkMMm5HLeWPbFpLKMf4sHmoTjhNtGcrmGjL
0CfF5TTrOl4zNEPxJZ0puL67mJIMAak6owKnmSlTYevDbmvRB6yVtoi2an+PchTS
NZQHVm186v1vuOBlu2MduTs5DPjn/kMHcJGLjdRboZwseQPoovtIk3b0jJ6YVARZ
mdOjs2YNX3BKVb9Fwmuon3OUdCIrYcdZ63u1SQfejWr9VGB02Y5ax36z+MUbOfsR
UnoDRsrmgreC+YqJ3FItGGVew5JI8SFqV0oJlxqZWr256vFFC/y+9YGv2CE/053K
IFV246IwoW8DSR3cjRhhQ2YwMMbhz9CtcPkLAseaFEFGgWh6dRVJvr7hjAtMBEuj
Fhhpx6W8p+VmjGeHKxpmVlbjW8ADr+jhIDBsQiLL6gLtkI8/Sd5v1oDoK3O8WQuH
C9lSSsdn7TJnua7UIY0j4u47FGxzOCXe6P8HoCc8UFYG+ns9DOwkrK5KPUiEZrzp
cMOBg5DBS5Nk5BPcmXJlazOFG4bcdhtob0uIpN3/vcrYt1b4GSrPue5CIOoOCp4P
vZrpNoFPPYTC9snqEaDuNiNdT+Jx+XyhyrYDdjy22v9gUVCKzzTGAjGs4aE5RzcN
UKkvwTSNopojUcRbNooBsSFq7EW3VLc1BgG+QJQmTltXoCWDV76UEYTK2DM1LsmC
r1JHPnTPUbcoZpTTDoRoAnNTzOsMEZf1rjrFJ8AaKZ10hgoTOElBPZUhU9aiUNTm
5AGNKYco3L9L8nW9I+SaOoCq8TIKwxnqf6Z95lMCamHoj1a73f8PGBrw+pYrBKcn
T11WHS5mi6JlYUAsSpTobaiOpF2DwCpQXYzkyp/+OMPktGvFdu/bm8gz0PjQNs5n
/u0kIWYPEQPxw+jrQ0sJTN0XcawBcWgf4pZddLNLkT1cID9qdTabJMJYU6dX878y
lSPffs0jOxGgRKKps5lBP69Kbdxy8VjKS6wm8VZ0IPvHuzsefhVr3k2gE2btz5S5
b7B043i4oce4eJp67b++lYHivkt9wFHMks+u8O3YLb7an8pf3QNbpsqc0hf0CD5j
3J3YGONsMetlu3b5bjYYARGWPJQb6FIUbDO95QBk0LLk0Pt5NFIvq4CC6vvfehFn
ecwrG4+lRuAQ5Jlhe8AkXufdue6mLNy7hBbsnRIPip/ABcrycrRtnwbNpEj6J2bb
75jzaeHGyhs3zseC985t4yk56SWgFEQI2aw+Fg0kajpkYesPqO5SxoDFbaT54TNH
buL0LwqYNupkyFXUQtvdy+jMy9XOGhx+rxSqO95GrSrUgJNvkkrI/+jlmr/QBUGo
6VIv/B+mp/PcMBZRarxMYMbcPEg6LxWkLsTVnFt6ApkTRTzZfphZF/1F2Wbkwd9a
8qkwnhgnfUYoF27IXhwVKGARK2TGpFqVSut3l6Z7V/c++Y5Kv5Ww+LLuweEKtfWn
swNbuPDCMugPX3T7Lwhe6rAZ8RB0vhEeW1IyGv2dU31UJWSWJkXE7+ZlGdectr4p
4/KWyuDwvbWqLDsrZ+mlRl6CjWKKq1VBtzfF/wOpROm1hLuf6kcrwxtkaZ6A/h66
WOSxPfSWHpv9fkFqVeCcGdyoJrWJcIUEYmifMKXm4d/z1HuYrFuE/nw9+iin2c7f
voJNAyVgIezLoxvDPuV+XlZzuk92Z4GZixpNhPJnnWtTrNjVtKFy6//QkUfKd8WV
T6NWaH1WmlNZ5R2zKoh1WSgRxEHRIGcDiHkMumAGiTzCS0jkUSeQroSj5L8EYZAU
YYCkGJhXgM1XEw6lKbNea82owXmthGPUctkMrJgaFbOAuz+yqtBREdCMFAq3WJwS
kl2kz8XNZ1tEW59haiT1fqG5E0b2nq/9fTNGIW0BE1MGKCTlKwI5g2vX4NHbxJas
+5sS8XqKRqLGfdza8FnSCl70/WKlbGns2x6SdAMTFHiKqZLXQl+nIQBPnV4OlF2f
HQByKGKrr2ALNvsHf/ob7V7odrqWW4oWF2nbgR0UekkgxXsIUWU7JC+kK9p0OdLV
IeD3O+hJCe/zMhIrUUNF9PzUauXl1MzFmf1QD0YPJr20OW7/zsUdpGiKArRQFdeq
xxXkWsDCNLyx0xln3WGCfcuWITT1b55sa+fixA6ul48+4S9DsQdO95ArRRRS/1oT
SzsUbCd5r1MJhU3KBsxS+4+B9u5Iu0/ZdU1TO8EEDlBVGWylFgOINz6zhojUvJQG
O9AuEDYA/OEncZvBRE3t+dP3i14+TtJKS0MZxY1yPf0yogD56FJde8ArJLce4BsS
iS+mTCX/T3ks/ct28V5XWH9znjha6jihp3w3RRsvk2nlRkdXfN0WkQpni0LnqtjN
9Q+o6FnrkSF1OJpdHfz+pECp7hbVccqMrp8n0+sRpgS5UghZyukjvbttRe7jNzmO
l4ea7lDIe/FN8bD9QlU4WiWlhvMCizPwZ6tQZVgmftMQ+I8r6cXndH9XcJPji3ft
Q+BjI8+gYvhtDikdmf7A0ApV7j3KuKcs1sJOFIAjqF9onmnx1XSBx67ydPakkNhe
TkoIFqEI66XyNtxjKLZyhsfK8iIdOVhZMzFDBKWNVeCoSwoduHV7pqUBdfjFPlX+
CKZkU21/eYMRN2VCKhgICioV6u8btCf9TTh6xLLXWp+HB+ne4cN19qIMdnTCr/bc
HfWDphy4+JEb0X3EjVkVY2DZUNWr/31twVgMVhFV2MHamvEcyo6+PoUg1XVQc9eg
GHPHW832gKOiNpu3M6EUsBbatmcrJDE1ZN5DBsO6o/CxKy/sLlbEH2AfmVp2MvXY
M30C4JVT1Bnh019e2rCDRC3TpfsrjG9SexvcyGvCJ3AxdhQxFRcFZnF45HWamJ6/
zk3WduDMaiPyNv+w9PFkq+99ZHVjvLlErGC/cA/yy8c0X0C1H/J5+cIIC+4KE27X
N+GJ8z3x/iosC28pMFeRgAfHXlk8UvILnOoY1pjA4kHo4mN7QIeysZ1YWx5jgS0K
i9yiXN1WVJz1LNWF5W4VQ5R8sBVSEt5KUHbkvxe+8tEYc7F9v0mGMEHhSEC0sE9O
aLRtLmu5jjd5aAomEGH5+EI5yyVE35yJFM9B04wtqvCRQkqUlzKXWxPqURXCJIHr
xGMCR3EJoP3KZJ6K6HSmD0jacuNFBrw/MgtoCHWtjT+vvx7vWWJK7xlb/HfDPwXI
uB6yCVW/Y8ocxsBzICRswy4AjXFdhx2X86yGV27BE3LPNuQNMqA/1kBOjebBcNo8
yc/Lcjml12+/EqZUDUrsgCkXmmUpUfh08dvf/p+VIu3FRnPsiF2srczivdJsezLz
tv6anRJUmsgHh6+mHXhDsFxkNgKrAKci4d9qy7CND10Hq1q/1lGo2gbd9SrFdsQU
Cj9JcdNlzurDTK61wQDpJL42rTR+3+xFhq8DmXA1phX4W1GzuEHsYLEcHmApFPVu
Os4Hq3dkbrPs6za2UepuV5JKjENRGAmRAG/aCriCbY+pOBK3ysFtKCzzSlZbJiEU
IEF7Tg9FWvGc2PWQyElwj85TPwCAWThPe5QfxpLCnKU8QNvLMkAj/U4qc0rouMbo
5Nt52QhCY/zSOW3/D3wFD+TAWFT3Z5HDvm5/U1dachT4kj9HUjTT8I/FXJxuG92Q
RW1x4hNlJFr1Cq77HleEV39KlkBUx2m8ePDT9m0GUX+W3+awUWPuL64wd1jzK94T
SLckv0RyvnTJuM0ObF533LAH5QJwGlFWmlVdc8M6dji9YBiwvdtjIevaKol4alaO
D2GKuJz0Zp+P1qRgvuYz5e8fxbGcvIHaSEaGrD7lyKFn4f2tCMTxbjZC7sfYvQ2n
wZpY370AvZHPF+wuOoXas1KxOejfrHkoou8EZw062pTQnnjIra7b15IVqhtlnHGl
OMne9yp9MfTxT6rQ4OkUKi62f5Jbhbpghqu1QkZ2uqieB+Qo/+lpdfMNIiBiiW66
QrFDar7wt9h/RQwGNQMErwwb8amEhV6FHPNYT9dGvhkE2z70HxwUSg3R+JwSo+2W
KeM7ubXz3qNe82ONoJfPXeJ6HQCDHEJt+egHjj3q8rJ/WPkAVdkwsmMkqql/yhgO
oxDj2jWDPTaUX5maozL0xmIZ1VNXn+nHnQmIRr5+odq8zvO/mkP8Llq0GMMcVEEP
dCebzMFpVIepT9qAb4FmxPrdVUufHq8pTYp96yevFbX24tpkAjmL4Qw3nOstfUf7
O8/54covt+fWRN/U95PS7+BE1sehBu9F4BUKfjzQA7pHUI4ZZQ1NsJPAwuaGiKlu
mkrAmham05CmOzWOFubHJ8J9Up84bRsUf23yXtPBoUPQg6QeIHYHV4NeTilu5AqD
roOUhaE+CjYx88AfenjZQOlv0crRUo90YCbt1yQFtdk/XSgKR5/rbdlS+Al2DxiU
1Ex5aFBkuXehEeOyW0er+xLUGUrZ9z3aKvOjHSm881/znP7aA73wuW7pqBUxCK/7
u7J3Hq3ZhMqj8LJOMrG1c3vNqV8KZGt8ug2KK/UuRhFiZs118ptcqcaEXZZla9JQ
SlAQF6K4M34B9/AdAAXMTN0EPr0QP53nWrYKsz2D1kJn8W2Cyapk6LxO0o0ouUDR
uyiTYAlDYiup3Y8jwX/H33bUAX9V0U0NAUpVeZvljP6kMGfJ+gzCEWwWmrQaoFYU
yFLJg8GzIARgmjqv03GbgDT9LCEilUzzLE+p65WCIDwAnvaw0Y/OEHs/gVk33tzQ
eURT5PKb/6BdklTNrAZgm3zUnSFQ7npUnpl2QyQkG8j10BYVBFNekLBGDvDuaAXy
U0jblIAXJBl5pM+wTBVRrPzub4IE7T8QdEsa/U04Z+2LpHhe8OiuKfmMFcBSE/4+
U45x+u+1+t2VbvFo0Etmvik81E26CUTDl0OoFQP3PRYmoeuC/vRHORbar3XWfF+B
iykhBHXWhZu7/I2JPYK750/y4jXlVjem7RL6hs4ZLK/AvlBGJBUvKaTA7Uzb9xb/
JQxbtwl/lS1vRuOqhixRQ4guWr5o3pf50V9776EAE/gVCZLd0oIbLRrRap2QGo29
2869d3nVrKA2o9hFvhlQLkSq7wNmxrvu4yVEtFTtLPb08NFb0XBfGeFARMKJFi07
0B68E0aYDn3vfahjHbp7t0co5XKnhl4Jk7Wnfx2rZOIEx1rnq7/usDTD0Zizl1TH
M/hSiJehor7rBSPBssy6Oq1uam3DwCNQV5Y3+5FBttN3YOU1JRS68NxuVKjSFeo0
u/dKIkZ7hAXySeeuNL0tGT44sOfeZt2uItZFbRqDRFRM4cRHW2AGX/EvYwShG07V
q0xFj09XPQ+OzU0gpX0UNLnPjpgUJppzi13G8qFB+O/8cZytEqMagtesvQdhD2tJ
uwmHI/DkKucs7R+Ie8f562BgERbS9a2YXgluMzlERfm9efxE90HTP6dF4I2UxWCQ
Z/6RaY+PTyWVLfhHvlUp053QFlpeiMtX3MFCDkLNBqs6HAnfaOcDH7G78/N/9NrJ
BMs3QjafFGD9Te5CBdHlXwdoXUV6BFetRE+M6ZlBJnXHScNKTWUy/e/mcCGsN7Ym
l6mymnv+6g/zbFz/XRkN1wUn1Ssn1Z5SWiOjJ7hO+7ASceSdmTbt6g/1JaA9Ooxy
jVH207qtZ6tdUYWtQi7P4Ojd3/VkLsD2xPh3iMJ2jH7AulZ7yhjdRZxBtcDUqQBX
WEeoMSoKiuiulSywRzdlew1Ba5j8OfA9Lji0yZ/uhYAloQCKo8PBWI8LZbqNhvc0
v+s54Kktkj8nJa0GyDZ0ijgd2xZ48CvKIV+Dbkb4r0wwOf6asR/EDqFog2oA/BVX
h/xxYCzfWtQTLLITJc/eZ7RaqboEiJi2fcN9tFvvoHcE0GrwK/NP4duvQr5p2KwR
S+h8L/HvwqMzSfrFQJNOue8RzTkSe9DmnAXT4bji4BTyuKIz6eoZznU2L0aV1GsE
7WeTH7UQ2XW8fVUQnXulp4s1vFttshzH68mXWvgRYUx4kGiXWxhOKhZ8Mu1VbdR0
0P4vVoLeFyMJ8dRpb/+UeRsu5IQFIDvwzWHwnnc+dSGoNJJXlYyj9nAQxSTZHi8D
fON7AvsipEQgQ1OvtfLN7h+9My7+plMNLGUa8Guw5XDHtAETndcd7pFEZDyCqzSt
O92+0gneMHLysu9hjOJteIJxlZ14rbtObtgEksIztXV/MdwuNJ10crndLQn50ehH
r2HyVSonfFnjWD9EjMmKM280awP0ot7v6HnheN8HGTeHDJddMFahFmOblMwme6/v
bCljW6jfQ9eAHEMgzlEgdo7IKWRLuJ6jw+puatLarZWFDtvO4A3y7sOT0ni/IQG2
1g5iM3BGrCFYK81kZ380q82eNOUSC2dster0dmquEYGo8PsnL9+vJ83bL5LhSFsx
JJH1o1Rqcl9tx6Fgr/Iff7BMuBHKQIkJ0g3nK1oo4kqf7QbG/rI957ubEaqFmzd+
yQe8HIZverpDkBv0KR1/hFAZwj1lJinDoTKEaGAc88TyRU8kk7jDogokoOMOdK6l
7d+Es0H2cltlQTxUXh7EMzySPnVARyyeEV/eyIAxROXmHvIJHBi0HbOmsOE5tnUp
XEZEiDh5EFm8GauEgDOwBbmWVABpU4sb6VHXuhjNaZiD84TCP/XHkAU/PqgQS2eK
vGGgwF/32ZNm14dkt7J85KxVx2P+Lhfcs8qegGxQWDxqMyEcsbJdmUmiWud+yr9M
blg+9vhAJzqrKDP357FmuEHGh9T5zsZuSEfD9A1KHHO49ClLLarhIicc1fLn0fWx
BorNRGSPkrdMCL0GgZXyq3H6DPxaSQqnc0GFKdR38ZFiq7uiVMvTknBqPJkEieXq
2ecGz9mvM4BDTe380lDyHREGsuQUBNEo5RliUW9t+ZWaS45duDD2neF4IgYzYguE
ikSXb6AWAJYGCPofrp1GT4aPMYgVPpTErPZYsOOFw2I2m3G5FFqd3jyxnhBlYTuT
5XnD48N8vl5Ap/8dpPWGcZHcKmOW9uto2M7awumqfp6qH7UhHhnXMZZVEMeMfmzP
Ow8hTiKkwBOVm0q6sCZb8MVRz1aAFfqlwD7sFLXy69ceIaJxQ8LPrdq9WoJvZhln
ow3KPeQCKBb1+VcNFamCr6giNr9Bv+gHSPm5uq7zC6nJCes+GQBDvJsv5GH00kve
XeHFrajVXEcg54s3tCxpIzy0wBi8EggEo5znz5TdH65MHrjMz6A7WtN5wtzF5vDx
uwf+PPPbWIeucdYD86JG2NXxIK83Z9HH7eWA+ilvFbpLOxoUUotNLrVK//UOYGCL
lzA8O8VoMky9iO7clrgoHtHeDUZYsNO9b/moir9zLf1/yuphp4/y/UpGF0aqkaGR
d6l8tDrrGYqGymjIrRYKv5gFqIF3VGnBUU2CzixK8S4PYZpjCGSW5nH0TP/KwghE
jrkjggsde/k72KrMohn99XUH+xwBao1z5qIntXu4THlHy+PxMMPlQB+QLy7CNlTe
ntqyfjGG4wOK5AksYD0tHhNUoXlWNLtiW3FjI+c05S9XPuPtz4K0lYuL2Yz75Y+j
93VXg3u0ECMhC8NqU1+LUev9oAlA10J2Bl+jvcI7sBBJeTWKsXvc8jYGC8bnn81i
qitxgPJQo/NWf1ceCB2XdtkSd28ha3ZJYAkGqJIIxfl6pBK73ag72kUbrUIY9mHM
0f/E3E08ZNA/7DeVXKYY/VRGAUlWO9yy7HtDSwn1xNai9d2zlp2zvcG8sLLmVb/H
emZB0B04f+JwNuw+mJdc/r0yrOIQP2OREE8V0QKSkz5WwVdWZx+kgcHfJHE0WIHc
hnm9fF93RmgRVPoLow2T9wiYLuXlg7sKzJLl9HGqFcbufFYVEbWN/wOEyjtED/Fd
rav/ZhzktZ7AVmE0IgNQHI89S3RBTWZ0qUnjee/2HVvEqErQRsNLxTODlUlgfDoX
WHHremIM4Q2+//WdRFWHx3Jw33ffwtb6X0S0twQoV0ZxNr3HVrKuNu48HRG/wvvA
RxcGQsEeFHavU10+DAx1qDIv2a9NHZaoF6D+y4lMObUTTql29Jzwd7SqMw64zwe9
p+9stSvfGEwssX7Wcsv1TKhPaIGNZmII/Kk8uO8vtCeKP4VCf0uriFi0qZdSFFE6
V1xUN6AUAFPXJEiLUMbZmSLs1qawf+sUaavOstomz7dsKJzvaoQTvgITXmnL+3vE
Mu8zsw3Xq+HoJT8cEYWDReM0n37I+HrAnwubASPYlV0060wQ5/+V4U7G/a1DCdlW
CEO31ntJVI5EnHYDJ9E1oLaEDNCYpKSqO0M/MCo67DeISlZkoKiui2w6jTo63vuv
5bMHl3eLLgoVyoADXenGtsNFWibJNGCRwtOCUctT8Rf6TxWNDP7FxXv8kXjeH94R
4mcZCOxOnE9emMX08JZuiLfIgDnqnHvd0ifOO5bnJ/NuOnKT3flFNwtbyRlka2gY
UnAFSvZUhWr95RF0/27P24ekW7N0UjOE1KkpbarqzG4lMwncrG7yYNJ5FnFE0cCD
OgGrSddt2I0cWv41g3uqQZsKl7U24D/bA7HiLD6KdE+Kqzdo0AS5I2vu+kvEzz0+
RF+iFQA7pzEYmDi+PQuGE1acIesNjH3qwu3W0J1Q0qUAK5yD0C3DKGDIRznO64cm
GrfQqInvnxO/n4YIBG/iUd33EvvcvF11TMA0N4X9jrQaPto+/FNprKqfmYB13Hsl
tLLAvGzPwVhmCjdXZtmw883hGGttz862zeEV+ZljIfqgtQMqz8lriedEpSrm5YNd
SlZ43JCVtipnHkGGJE6bviOnLvD25nPcVFI5VC3gWwXH33RWGm4h89JPjJfo/0/h
W94fkE96RT09ZY6Gtv8aabJM3H0N0DuLrE4bwXaeJZir92xGJf+pGAdJWuiuW2Ep
R10EDwyWKW0jw1B0H7/R6XHDp7cZDbLCoQfo0ksRmn6q32DY3yfwEQVEjqZD8bqd
H3gaNK/s1cc6mzJHTmBQbhAq8TQAOHZ8FaCuYCD5bXlB+ukOqeuFRFYt18xQvSqd
wQUWbxW3DxdW9hkX0FlP4xgPEymvs19X+43JCCmwwkBA/Qih3DH0qcrvmKuoOQod
/0vTFbtO9sXpOAK93peaCIVrOTFwV8JAqzUedYEqD1X0xsrrltSVHk1viML+O2bw
khIgCldEVL+HC1xl3qDtsR7JJ3oQKnfJNdtqoF5q4bbmWWpoEhmNlbCLZCnMaD6v
3E1fschLFt0SDJfb6F+BZO7ooNIRuptAyVb6BzNQxdoz64DYYyFtWPRVWdKAE23j
TmkxPUK2wFYKJ6sZw6hdClijQ9hMuimxN+zGNhDk0sjNjjICnIqqeAAIr0mmXogs
uTOqNiz3UbwNb3Mh1nZuz8nO0QJT3F5DJeYNN3JMjNhU5DBHo3Bk2CbmKKPhgGEY
iVDxw/GPYTo9QcoJyawufbJA7k62oclxUC/paTrvN5mwV3hdgMrTKKs6eZY274vA
/SNDmkkhgOBPwO0qUHYNOSHdp2/YsvCcOKlbtIoNDNGimQRGjj3P5A/f+i3wkd05
vndoI/kYYAPSHV3331/jVJ51B1np2XlOB1chZprdBvfSo5jLzIUcIZdzSec5rTpg
tEkPXyVz82jYiPJE7oHhh0oyPQfsDkE1U9HKJEQNNaKBgufzqHB+30Ln8yyDhSXn
I3YAH28RFer01iMcTtlQVry1lfBnQrDqvQMMibWvkPHFWqc1p3JI9ODZgWkhrER4
0mHcvw+tskBCSm6NIoh2Zi3u3kdhvoOKqI6z2q11ZbO3o5rPX9wYiCrczlNDBiGI
Gfv1QsS7A9RGarkuJEiQJWIWtF1UTgrBiOQVZzHfMlHs9Jc5LWPxgknuYp8C9rKe
RWoWeHYRjBsOhWu2rzlqqwWKQjnQJpn3JCFzDyUWdWzAWraHw7ffzKOMZf6yiZeK
PxUGz6+/NB7iNP1HoyHuXHITh7fAEw5ANLXuExl9iF3icrM+afmIsuyKf0BgKNoI
7YEDsmNF3MM3VK/A198yWYVM0v7PNK+nqqwv8vGJ8uN5axS7H8zDoEbjDPs8+/HP
Fk7h64sX+RFd2MLwcEzYnrATJ7n2SsVExP7h3BJzv/lMsILlmNBsK/mxPCyq3MNN
04OVTSQPggMkW4sfjcf1SM1EkD5qxTVjYF7BEtTpMkNnGhB+OkBlhW8txtrWoPHl
XUgYvhCeDUODECAaG3NXaXWoUFtZuQAfeg6XFzsTdFowY91YVNL130m5WX0uhWlb
fLskxHjssJYQW0DPtE9boB84rikqQFLt8CeNjABPXy0F2J8QT9m5XnxxzexPM08t
TLJz92o/xbysaMHmZBIAcmluT9FYG4qBiO77VhDQ6x8XME6CiYFL23tunQqwWVAs
MBY/BWagRtYmGJo0Khl+p8sLjkdhMzdNKeexCpSRxL7nJuWrZ9WGnUCetv5CJYfr
BddDzbSWJNFWUKQv+X7aY5pVrjrWOF44nWDWAQPpvhkueMfVQqIahlcK67GgyQQ4
hDIRpgRJqidhGVgWOoTNh3FVhqSLZkYWUG6Qp8NNki5Q1gpp2vWhWjDmEuqsDo1c
x8K2Qb9Eo02+Wy4HNiC+/+8rrHrooqUaLC2UwipBHqJWdxY5GpKy1bPAaSXPygYl
HV0RzED3dTuQZ9/l5afAYOi8W+ME/9dsewV2GpIhBMOeUMBTb0XzX0VAcA+rJwyZ
42CyafmWp7qHwMfqXrF3k2suvf389dbk+BuISKC0Wwoe4ULwnBa08As4tRSaGk/I
ioBaP5a6PpsdH5Aoprt3Pw/ZZia/oGPuwbKTXh4NvTH5uQ50VCVt6bczv4MtlxTY
FxWbHg5RuMIahimrrdWaHPwGwFSAyHNk1BSSIQTlQB3tPQraLcA05hsJ9wVBa3W4
LFnaPl6CHXdCLHH9L0iLGdtjKWhCCvw1FIxQxdW+PxanZZdLAJhZN0c75Fy2amhy
oYPbKBezxnCIvc/JQQLqrZmVGtAZBifqHT8vgeWhBoVc2O6wy1mhVowNaNwttClt
3AYdaX+51yza+HHwe1md030dyFKqn9OKBDu8bW1FEmtpuXGDQ2xAEAbhBV0bzGbe
gxIjGFV2Y32uPbfPGQp6n75Ia14VZ1/ojGWIjhKIeUBVCegh36H/IyFBZ0wt4Tou
cKKMV2+a2jMhvHCoUrhvGuCS3Cew0J5wQrJtJKh9Z1+XOddpj6kbbL6h/PF1szCM
AYajeM/5MDAbrTvdx1rfhCWB8jMrWBKAQJigoH8PLr6Fq2vF1DSTFOg0MUWqV2ty
HZ4meVxuZL9ghbv0b3dkOtWdiNym4o2lIRlpCzWmos62v8GVpBwS09dxFBSlEew7
qxDS21+PNbKP6hCwYaq2z2w+OHdYUMBl43cm/mSLLXu5KMknCEkaBhCjBS9Oxf/I
ibcReyWKSVa06Rtd70QZgSE0TqdTFowj7omBdzbNMxeQYq1g/PmYdAAorq0Zd7qp
IixBwYul9As/9+p+DJqgUByHc+NkHexjF+Yr/YXMM1LxUk7Icz9b9K5PUK/i48GW
Gi/2H9cfhCW7Ba3cniTsmv+BinHulmPRb0BbXoKpfh/nOEzvzHBA+y9/9j4JBCQ5
YoHjpNU1EGcrjswIwBvRDlbPD0e9Smtlx/y1rTgJ+hjGOE0gC1jPwZN4hdqSJ2BA
vE1lBEWJ5sHlWXg+QbvUg5zL4z34VDU+Q79kw2GIhV2ANRzwAvUk8rnQ8vKZHMou
1aVXtgbYYMRCqSPnNE912p9fxTLX1Fgp56YtjiFURCXSF3LUp24lR62At5/4/6B8
gvZ63kwhIxUZFfc4P/SGxUE14QYnAFhAk6jE95ANIOAnytExz4xgmvZSakJRzosx
c1drEI4QHjT0KP4DBNFJ3pNgD7kVQBqaF0PJC5OyhoJrL/0ZF27HuEcNtwf38VOY
bkpfO6e6aOZfqCacdt+5MU6nIc8EazVCwZT/UqBAQX87g0Btww0Sw7uiJprXCI+3
Ic4kMnh9afZ87hUkTc2Y+Rnarg51JdZngnC0lthgm9n6S/8fV4CBw2Z+1mqeFJYu
rTQBSUVI0hGC4F/ru37+k6LCH1hQyH18l7Uj8+RHuYET/N7m5ww2Aao1yY8My159
JqYSowAuRjX8944DP2hHk4fkpyAYivybWbCIJQWp3ZD/oaAtNxdAj4Le2QMvpTKC
2hFuN238iOjctfh36XtsvQAEl32Zkc1UxZ4GPEM8hWyTOixi1o7onLkrpRUTMldt
k306/ZCLZ3aiwWQOTtAppx8fCugRBjIuN+QReHMY4MygwEFgqon/fhvgDpJDF+kB
+4az78L6UocYs78PjcWeh+J+2BuFpPMLMfM68UStzyNEMXg/V0mxWVTlFNw12fd/
wh0xyOY8hPAZe/sNqnF8YTnmBEexJA4ozFcpAe1XwJIt3tLejjARIHn3rSiaeJXV
LG/iON/gdYDbp6bBBB9v5K38E5nHvn9fso5CCzkPbWjnyre6Z2uSBOuq8so+Zt/E
zXKnBpgifYi17K3mY9wZMB9Hsx6QBEnJt7Xp/zgGkX5FlG1VdONlF8v9Lq7TM8hc
65mciaMLcxJkXcGQadgJxrbF4pbTy8iesgBRNKmsLEavhDAHQ0GmIVOl88yJP+Rs
7wLN3rYY4Lzho/uoWaNIeNLWyRCrPBg5D59O9pjse7LYQUJZKaxxpYviH2Wyf9Gs
97GPaO6Vy/lqnEYvudKZVJL8s8pl2uEVg/t3Gu5mjvfhmvgE3ie/DCjvy4du/Jk+
RGROS/h9pDdQTut26vmyDKI/TghztpYbm2h2/TMFdM0+vTO1fSZCQ03Ff+28HBGu
EvwVNgHLIykDGaTt3bvg+FcUX2ccmIzvPGxd3BPskJta0FS+EXPaegEI1c7+y9Vp
A300Hl/jP63LOeT6hbT2x5OY14Dl4E+aZ6agSwXmXUfExAju3VxJrlkw0rnf8gj+
CPGZsVeSvDZbHoB4GBVCEIVUQoDzYn1q9jA8/7DgkYJIl9nEc3693LT3NBoGxbZW
iTaEMqZdfONdWY5U/7L4y+irfih0F51PnmzMc5YfJSl3sfmaGQVmFPfumCrUG46i
RzY01TQ7tnDhijMVYgyFLGs9URk2tQF11EGTJEMiOoSjIFPKXXlVbIWvTX6iMXQ0
Txea+SNxt8RkAqkhGGPCzQ6dhF6dIR6iatwRsF2ieVR6/923zv5VEkv+7BzPOMlY
//566pOAEGqY5Wx0uW3qM8IGrq91DFGdvuZwwCGD9jpqjCAMIK/JyXmxdTCCGLlX
9S1lQ9KXfJB6/tiT3LpL3GQg8Ni5yjKqqJIMGZpKKy1rbAM0aWX8lpqoEIvr1iLY
1I/ZnVdSa8j+65PfLi89FcXKkH3qWCt9C6I1szXJARZrzavY3btKCv3+nlAHDfpQ
7RfJ0ol5GnoeLCcqzCM7dWPC0CclcKQS8P7K3V/TRbVvT7eyxuWBhg9q1ezdgkgC
pd3JaD4Xoeb3wG3rYeFAL3af5coU8sNakFyVXUpx26c4y5x/GXGSw6HXqyFZLxNG
KKBNEEeSYJCHg5ZM0WEMz6TigeIK5biznMAx6Mh5TN5Jed5D9puxL7n5DTwxbIoV
lcy2nIDDCdBWIo+SzAckocgN06IYOmX87bDvyapbHuCeBF716VM4Yrp+cE348tvZ
DFyO5jOyS56vL7ela5HYUB05XprAprCwJ2igMNNRfBigOOf8FDnXwuxbJGPrUVEc
J+WR8C8ja8lN7iy6EWNmTyZyd67hzTIktxeECvBq5EBKTs5EKbN0ZoMLQV0J6Gjp
J55DvqIE8FOK80PWoCk5loiY+uSMUagD3JMcRnRqKz1Sa+yx4+T9xesG9Ck0lZVq
vQyNfb7irt70X7QzgMRVixGoPR+ZIW8PiA5ptCQWQHTU0TkSVDucFK/MwoDEDSrQ
6k8kNlMgzxpOhiJOmwDSwsJJX4M/cHcGdWnZ8J0e4pPcQ6C/MABfx4464o8IvvCI
4mscwfOeRIVp95zzd7+oYfNpAAIpergoFhgzlKfLkvrpviDEP5+zf/nc7UHdatXf
IQO+26VsROHs7rmlc0cmt3FhMbcTzqZK9CU25vkyr3Zt/v2TF/oTa6nJsiSkD1AE
bXOopRs//j8EihDHcFja9RtNmXmXRFCBiS5StpsrOZQ2hTmFL2A8nUJZKv5arpJl
bV0LN3vFcJN+bF2KbY6LGZd6gQ5sEzIAWfNPUGeQCoYOnyxC5xU0P5I7i+cOMMfz
sILKF8NhmwMfci+GTlZijud4v7izLfZZ9bnFPbcueWBLezm00ohR4MdfoEZ/yQri
UUP9QFMGMCW+lT+SG0ut6LdblnZIknBoUtR4KEWQcowYthHT4sQ50esn6mnVXc6g
RuD+7bw/EL4BQrOF6XgB0r1Frwhe0IPtt9r1qPqJvwUhOmerD3rchOwJZXoPElBn
viI6H7Pj/WQx3O2Bg1rwWZveABrsicOsgp4yYHp1kDMzQA2a/Xob47s1SPsxz380
QUO/NB09GhPUqtlJR386oR4dtd3hWi75Wnkj22/LRkV2comNoEiYhW0ZmHiakFEE
hBrvdjC9qLhPWe4/xxTEn0KtivwCMOCjdPSCeJIjm1ty4POvt0roaaAaeOz4qIDB
Owu1LFokGlMXGsQIWKeIJiSNB2ZRPjrZSnqEjy67tkd/k8/iZq+jmozxbVFojZnj
Pppntst+aoJhLTYTA+YuFBD5YNRWp6u2Gy4oa3bEG7tvJt2XgIDyGM0n3crkm/WT
A4uMoZ2fnXAT7qqLQwThpn1QUxtW535XSHy5+3GR0sqE/6qSNKyCGJEFMxjyHc51
CH8wsRpQ7fOjP8H3W+5oPJ54y25/eJ03xWEmsDJTvyRNYgX25miKA0akc8sU5Dla
CwcbnwqaB+99MmxJ+Br1YRIsqb/5f4Ihcyj4J0eq/8VK30+YxLm86A9kOiYniMVe
DEOFxqAXipya6iQKUS86KvrFz+1NRBCnT/fgsyYCZIGBCLqyI9k63WwbDYV6ZFTX
tm+fWjyEbz+HFTluLna9fzfjlzzXfSixw/dyjxh1UM8Khemhrn16g2Gbhq04+QUC
TyOKjG9KhJD6/iLYkQQ/Cvd58qsxxeHZJLLj0bpSbj+DYFtE28kVSEwKQQfIi3bU
zHT5EK3at0s3dGnGscUD3QtJ3hppMZ393md3PR9rWS5d3YQ1LFW9VslDKLLUqUbM
mRgXsQPtBoy7UO1nJXkV/22HRhO2+4uE7uMfpaA8gEqGshhpkMS6AGF8ACJfTgmX
ekgsLyRtzEVYHltPhqCefOOZph+8rKEzKjKDru+FMB6XYlzMmByAMSlF33aah7lC
jirsU3L5mtiWdC30Iog2Noch16a19jd1ae3gnMNGAzjihKtYG2OBrWeckMASBntV
VhQBLPPNoJHnM4NF1WV9tawKAqFqznAEW/6DakygFP5wUxrymCUzdRfc3xC0Kbq8
FPkOyeiVnFCBBVL1x5oWDTjfCrfOjT+D+qf3TiepwW7z2dg+FNxkMxY7g7M03I/T
kh6UWQKRJjzryqebYOBfye+/da8+b2ReR3zINWnbwkTMupB9IvRx5sbdRnw+38Re
gqouWQG3nhiFL+7OzksU0NoHtFiAm0OAktZJDrl5x2n2V+5X00Tfef7qJqxz+liu
reld6devC3/I4lOTngsYpN6wSomc5KURNDzzMROA6+UzRgY8TkUHu06SCkrM0YFM
6XQIiQCfnfzstEeHhetSs/dOeAEA09qlheaqJ9bXsHa8tFORYcVoM2kIw81yX+x/
h7MBX5ZBANckNoZNNtM5w//1W2h/v9KbjqhuoC2u3RWhAGD7DEOcQC5toBQ4Sfih
igt2ouDITCC+c10x1sNfpVHTJ3Xf16/iuJ1y0jHtrWCoXObHQLIO/owzzvBT7P4F
DfK3b9EE9pxT1IcFqxgWvmsMRr2v1OG+FLSGZTIYGX6WGvs5sEwodY/55h59yBAg
8bcUt3zuHp5HiGnhyPzqYYsiGMMhqkzUbAQoqjM1pWflft/Ke+TlEtSodwg5P5zt
4X/I2o/G90nRvtHzU/XNHRsbt0tX7gBcRg0u5E2+D8aEqP8IkPNhRUxnHnxHvlu3
1mQPF3e20Ka9JxjCa1/kRwmtgAMQ4oErj5ZaoXHn+37S1FtO1oiYvxe3PfUiWt7D
D8WVly0SRzjJkGPfoZzG6l8pXJsElCdBjxgkZfrhdBaiZgWt53n0CSWLoKDBKK2O
1Y6eNYuN0dmgXEqZONlskThx/4aD6/XqU0BlsmIRBNPuUcfGMUiM6BS4ykn9gl+0
4fP3q3CN34SCJeXxT6kcQCFV78+Pb58PtG4BTDra6pCbuhvKj6dv0NsVLtOVx9h0
r9bagfxLVnrm02N0HouE444MWc1MC3d8x1+3U7BIAerbyI8fr1H8GmSpXIAUwieh
Q3reLCOy3Nmol/Nwg3UBhV1h79uPw5sfNgThv6XunRMPNdjZxpVqVGi+qxRh52CA
5fPB+LuRRTgRO6ir9imRxrLOW5Ovo5XeOVSGtCHIB8jqYIWJoQp6NvtdspAkTBLj
M+TlXpxzW3lqWXbQKmGqPMnhYyR15U1M+6jjwNQvApn8FxdqYLgjQGMfsvaOeDgW
kwZjLVvZRns2AtCFxGHGoOBKtwP2A/D2q4RGV4T/SIW3JLxslXx44SRmLbiSd9Q+
RsNsPcOGIaqCLgjxbI5LKfbHtqg9u8/Df+YOW0Zu3gqIrqUxLCw1xw8SsuoJy6cg
kOliaKKT7iV53GIG0dBJzNIw5SiChnkCKEd6+F0/jsfoTdnGqR4CS9vJFYRYoEFF
oc7lHVH2Q/76wrz9uPUy9Ls1Yd3o3zbwi0+YGMef8f6P8gHMHK7iwGDcyFK5GNbU
YFpq7Gn7wlyu9eXOtfCkjHtc/wAfPNbMDn3X5jR5Ui+B4fmVWGR/56weyJM6S1lF
7NNCg3M+XXkGtCUItvZkmRAF3UkaPQnhRT1G/1DPHhgCTYQpdl6pgPcIUnnjTkvj
cNx98L3UrYqmcu0b22Jylke9sApzJhI6oaK3fgwwm/Z6sOmZUz6rJOhVfx5ZaEkc
whhCIPMBZ9SnzvbxCPV5Qv0iNjeeVvxEnWuvUaL8a8xvsbtvOKLyCyDV7ANu0Wce
GoSX5voY5hY18+I1XHKCgDAPqMupK8jL82LtlWZPd/L3TYa1viwCnaeCv4hHLVkI
BHtbGX7v7IAPv/E8eapIrVsxgChZWAkBz5GTdImkK26ZXaGRGRWbohnHMcexC+Gh
/XWYYAo1hNAPjy9I7wCkurTRl4J0kySXoGl5zBreoO6kYkOQwBN1WrZNK/cFnPTl
bWH2mj/sP/T40zfHvtD+nfj2PRLIsLbDVle8j+bkmAme1Xe+llX95DVlpKj3o15C
BbkDtoMhbwyH1M9znGD4egarMIqUAwu3iiST1wIuNmPqE7whKQvLPnSQDJ6xwNrG
1r7s61Wz4dYwcMBz843bfH++7UfWlJxob1Jxb5om0KMqR78p/pBKf2jddo8VtxNG
ppooUJfDaccnETofKOFhyAVX2zF/W/DXSGVKoywMs4IWdQRuTBYkfDVV4Wq9hRZa
cp0gtegnLIeEiRPXvtkkXc3yapjtycNEyk9Ryw6g3w12Wlgl8kmpo02ssN9df+wa
JUYH3FQGNcxcn50UrU4TzBe9TBocLYBO7qEKhcpIgmra2QBtYM+q3Jq1SPSnvZN7
A4LQGVK3WuxS4Bnk24Plhwp/kcbhawQ98wOOcvnzJqmstpLCskwIBFggItoQDmDP
eE0uhBvd32UZA4FnA8WDiRoikNe5tZLv76FbvBGxrlt98t1LIEHdV3hrw9EHL1T2
wa2p4m9PX1o+2VC4fWUT9YXZbCTS/vOkHBMY0Alr6iwl1To6U2HBiYvxbhIqEeEe
V2iP3kB3N5Loe+sQQnyCItDBx2ijDp0akYV8U7nrbE2JOJIdVW0qDXAwXevQ8ld9
3BwqDrgLwDbey4466FZA8lOTIyreEsHqvY2+Grhxj0+VDGa91Z2Bn+O50mrBNXhh
qQHujvItNQko+AyKXmmXPmFhgvZrV1tFKO7T7FD01Oke8kGfxdR3y0wXon3wUWOD
n7vJXoakHUyK2V7KQFHFDu9NYED1TSit8/RSJjJE5NSi3lE/rSHTZcIAB7Oam0D7
5d6Lp1MHRhWsl8RUYk6fyJrWflmMCUT5jAYVyZog5Uy0XJunf+7UI2SGUf5l4VZ5
2QKMvjiNz9H2dSQ/ZUGj637gwKwSmZclhj/ny9YvjN//Xk6ouN+GdxsoGKDPgmY7
711bxHykYeRpf8R1EJ7h1IqKoxoRLIwxnQYeYbux05PlMCHMVjiQI6jvbpgioTSr
4Z/Pxp16gyd9713UsLftv3fTBNyZ29XcBc4Zn5ACA4iMwiZPWJM4lPgFVzuGuDMS
LyKHxTZ7AOggfdB/utXpAC+JqjNo4QJQqv89wZ2Osjopw6atyitIZD+jAgPrtfup
IBCXgpc7ISWT0WQmEOeE3gJX2OFrWo1T+Iud50tDmlr0WwYyMN8SIsD6s81t1Amw
f5e7a2Sa214lWMwvygkYSVpr2qvTwJk9FWbwxd6myfztmaibqeGjsg+eYfROHt+2
NBmkqU37hLWKJPhH2rhsgxaYhAUuLMbj9RY51WHvj07CjA+UoFjMyk1jq4AjZSft
TkktQo5nGOFhfoYlg3TsChSx4ob57N5ZT2sFBFQQPjPnk5YiH3+5LPqAGRehvL4y
pc2VaHpfhLX7OePt1VEQkZVQjt4GBeS5oBIdopeYbwO3otj9NFtGkOj4+wm6YSqZ
RPjN7AXHFnT5DKK8+eRvy3yYTHwD581TMLk9NrLNJIZtSvhCtLUqcKL5FP4u68YC
HtjMW/AaHslIZ2Z5QeiCRzm2xMxNp7dyjQbDCC2FU0/ay0FJCWkFH729cwbQUdi5
BsSFR97gkgPQn6lO0SyyNQcH0ldwiIuo3BX0oDAXjdThm1v3GvSugOlIo60cCBLL
4efo37Om31ykOB+yjenbQ8dGHIII6BeiwLsFWSlRu4uU4dFj4rnJ7hqEeF6lzC6Z
4fvdGdG8MeKI4MRxAniYNDcyM3CHe79BZomwpGp7HBhe050ALfPZx/dNodljq+bK
lNITAafErVLsXcIF2Eyy6Di+Pz7R8grZz4YI6y1Rj8/iJD+UKKbp/x4sH6bhSYnZ
WM/7eY31jkJ18LdvpPmcHwyp8E2pM3c9921EiydzBEV8WDTwooKsIvTR13OLnJj9
1GWBiAxB6vxT6Wya8XHNjO9qKCb/09jNzOP847tScC/3MN3VGCcgKAc5Tk9hqHFg
+SKOAZwBPKGjT0iLRza3C8GHfBgOTdGnvJoqX9n4GXeuB8+CZ2dSTPIn6f3I1+kr
ixFKyEmQcdPamMnQX8b9YWUVU0+kuQPGrHWxhwhK6lSFxkDU6RuivIBv68WL28fS
gywGlvC6VIQTsmqZ84e3r/aCwNIZRPwMCA1ZIQs/Xb39853KifImKskfVqb+6Ltg
TShj4BvQkM/gZ/NW75Bd1sw33ili4VX97NSHrW6sOznjsBh0Qm6loPuQ5IHyNKRt
sYeNnn5iU610DIenr+NJBVkFW6yuNVuqq5OnxR/HvdHn3wzxYJv9fkapuSuRyNh3
Bhi1DLwnwsaZLjBJUl3/yWMykaoqhR7zNCfqQozmzmpRulGqwlD5dpHKV7JfZ4to
KDYUNiEO2kixtWxALGzjJzuuRGTySKR4T5pRYOyREo/EqqiEcYRbg/nKuNYgeLnb
KYVDuF6/2t9NDKJol+tLoPNeXiFRChRsa4PI7ly+RQbs6VnJAZb4tY+0OV9B979j
EZfbDwv4SiETQOcMp1GDQIzwfk8V9XDPxy0Gikv5X795+KCYdil9AZmj66KKs4t4
WawnLny/UVwSN+TpHXJCeXmK8tkm2L/kBVKza//dVWQlNwr9dyEO4KDr/t2vRXgM
R8dA7/6PIivaNui2nBLX8t+nSthoO303LOH8+yyuFfFo5W1abPX7IzQI9SRaTanC
UlRlG8EDy0xj14D8Mpy6iibcHMYxUsTf+aNfOAf6oFpMhHDfFllNrw5Wj8Gozxmx
EF7TTtkTOOMGe/SRiIMgJMspLZFDFGIKzuueEgnSs6ARlv+oqjUjZxEf/zKVYDFf
1dyy2hlXbzAgRxJ0bXX1oSh+Qr8Y3AgviTrPTxs9wX3mLjI49epIJHGJg/VfoFCI
9l0v7QzmCl2SmWRR2yEdzXy2xx/x5EpiHy7MYOm4P5KYjbAXuis0OR0ayd9CpMMw
NMe2LUE/u2AwzCb8WDPk6GkHQAFetmwfiRlkgW4+6tW5bRJSJNvoTT7t1Yhm1jKb
Utqg0RDih450bC2GKb/jUdetNa5YeIiwHua12mu6hqCta+OM0EIu6vdW9nna6TXk
U9mcKlwmYSwD3q1wN9QueAXQNMN06zQcObKjFKTqcRYJynRDi+PUgaQHUc6xSdBe
3FtdOFa+r6wdMA8Bwc+hBmOFHGOCNKp684lt+kbqLw65lVI7wrDHXn/gfwEXqCip
u2KfLLoIQNu5OddBHLx0491U2NWzHKcCIcD+SwNzk1XUch4RFpLqq8MRHRJzNHvA
e32AJO8x/7zipdNCMCjSwG/0wp2cdWKB6uSLepRUQRmGbCGx6/AqqaKBblrJMeP3
WcWJnp65ZmWcThsu8NSJJWXkUV+xBhkYq7o+1fu0BF0e2AjqPk1Ha6E60Z+R0FSG
X0H5i6W0r5CUwjuAWuvheStri1QLHOHrpRLuQCBOdBTXacNj+M+rMbehaK+gA2If
gWDGF6eo9Bs/IbhOjhbHZkQw6XTjQVOAjN2t1Jui5XHJaZf9CJcI2oRTsry1FDC/
Lej45tLY1fMfuvLZJwZEMMBvYliENxCUiPpwlj7a1WkhhX2WYbSTHj+59MeiSsmN
+rFyweloAanW+oZuLTpxgbaZqsZX3mmrGzWK3JKgjAqvHM9cGbIKQohMSu2FUTQ4
m3m+D1JoG4UCatZjj4VZtyB3WbexBql+ZBnpPTgNSg+XfQOUkEKa2woL52E1eQZq
hEe7jJu57gsVpeooa+k8idZ6n3S6KINfV9qEhow85J/fL5J0gWIgwuPzFmOU4S5r
nQYYWRe7TLU9DG4PgdhUK4flUP+87BqioZVmLGosTlM35jStsulH+QMB6dPF9PpX
2zypLRt3HajL4I0TDxAf0Alfb2qO94bzfYPrn2LaWBQM6kwgpFea2QbhlMR4D1nz
sc01k84ySzKqmo3vKUdOcHCrSvZngI+uIqm8FDzPyz0r5HRFh+ElGnUKwnRQaTD9
YM8jOe8CXD1EUMZpse3PW9I4T/K4boaPrGJ4TqwcQMgJfX6GdPNTpjMKRiqFuM/e
4HLdlMvna238xFAMdCULNlvu4e9gyg0YFBT24ejwTV/20Zfgz36FTWr01BivNbZ/
tRzdFEXQTGQMy6BI+ML0rmkL4F7kMXMI5e8OPM/HWsZSV6AvhzvZaNFi2HkBxAt7
T7H/NTaPyLny3VgYe7OGFTFL5ny7ZsweDRr+AtWDF+PnaQjMof2vn+Kfd3InZ2mz
8SaHpdAoz+Szhae5FeNoEwgbSpUNpzHJFkdA3fL/VxGakWI92Ap1rp2wQOIe3F1B
izq59aN4JZMwJ9C1qmFHa/IjMJeWLYBwvPFwogTmijjDRYFl4pArx/HEbtQDEC4z
6kYuiEQ/+s93ejZqNEDy/WMhHIaQG7Zz7iU1j3LgNSr9iG6mvu0SlfZN9lTY7rDy
z6qEq4mjjbi1QfAG929HJL+KYlQrDZ5TnY2EBK/jt+S7p0SWlN7BmXsm93rT7MMN
PS0vOlIm4ITXsgd6LRA77EJklvAd6X9tz2OnT529WXsQcFGJrz5lzy0wxS8cu0oX
mnfFvtIhuzmxD4oa6evmy3skh+Ov7rl6BkQt02S6Dn2lLUaUfDGtGiEpo+W2jlu3
OnmCIQCJismvcMXGpC21Hbv1UDvW2OK1g8lYvcwnEnAMrMnlHHlguwP9odOR/83t
/07segAiY+NCWdRzrE5KJGm81qDisCd4Jljy1XkrueQwS4t+V+JYwxCWxxffrJzs
K+YXnYMwzcvHuU6WMMg3rXhWOru8eQsnvG9uKj3cb18OompfGmyfY1MC1ldLU+Qc
qp0KWotSfql6xr3Xs2Nfu6tz3iNRxV5cGzepREwxRw2n65jnO72TeTtz8ba7xRh6
gSuNZ/OP34sEtvKl+MFLtM+PDXAOWHxhIMN29Ag/2M5UKIN5zhb8MJy4pjaiYktT
+SjYH5upgmBIOTbqTP32NRyXjYEFCvToU0dF26EdeNqr4CpFAn6qiDS8P0B+T7f4
6/SofRMa+mbhv4fetanh0DQLNwknXq9fcM1Ww7gCUZH4lI+zNvgbkOBFocMZeEi/
6OVF9AA4vCamYlNiSAZIicJ/P3ifw5zcEraFLSx7kAVPOkBgbCP0ji4vonnO6UYv
hEjXUDmDII0KgIze3986tp4hrkTf06xH1HSrY4REei2kyk9UpH79d7YziCvbaIqC
V73n93ANTmwWksozU4kDPz1qt1sgqqkwQ+wEhVu+RhKcYh4xS+EUeO5OEz3hAFeQ
JSva7Gl8aVaGgnhXXE9hIUUzNqew6F7eM/9jLi/kgyxJkaZtEBWEMNpDQWUYRxvw
QRntjEQhonHaxSCSBPPUc9MX0ge/+d1BhrZnJcMfYVgWkLXlwY0/6+Qahk4rsQXF
TB7dyz0MXKepRcOuEIweFCPnErI315HHKVXji77CsGWQqmECCeJj+1RmoSqcHxQp
PVjZsDAvQReEKT482bdjxM7LZ3L5Q7F7kSWKV2okdRHBLQ+eSgztQtDtB6CccZ9g
j7+94c+ryw7E7+CDjmdHDUZchn5ZwA8IkE/8DrHxVE+gSZFNxD9LQyCYwQlpIb2s
vRiDe2oXiByMT8iWHyqaKN8Ll0zZxFTm3ix13As/xxnTD89ZgvG/950P6Apk64UQ
TT6SmHect7Y9THU78p2dwUhtwB5Mj/ShpQkuIvEm+prAFDFIOR+/j1VMY3EpZ13y
Hdj0jWeNSxxXPzALXQAfU8G7+TASZih9CCXd08OJdDiMKur/i00c9oL+Hhpr0oMV
bTfeBg333z2A3isuLgrktiSlaO8KsVCjl9xVYthtkMe/7YQWO23VHL9vIEy/mlUp
C/L5LCJ2TrMVoP8IfnHy5EMxNBqtv9EuZpxo8F5QVDJwFgMio6ohTOuhV8WSfohr
gIgjyzn/31gL4Z8+mVCRuEIYiOWnHjf/8e8x9JgrwR/kznmX35ZPduBb1RKQEq9l
agLEp4VsqaS4hhiDUby/8lzuSQnnFdg7/LlwPReyRsf6VwnG6WsSK/tIuzXnopLt
+teySRx7uP5nHQJxDz/xcaNQspTxF6JB9JoJvExOm3JSFAXPQ6JXGCAfGbB6mzZo
gFNBaw/P1FCqFm9sW+0XK1m5J2+y1p0qS9tJFS1wDsjobP+m1a3ardPMVXnhV+Xr
fLbadrWvNHqOwlG6xOKS+eq4+SEpgH8/5ta+PO5GIozqgJ0ju0tOhf9rRtALSRxb
wxtSqi15wP4HfQhOrlsAq+AtT8WWklGZ6xTNGZlw6jcpui8mgQb6Z5acbRTVKSe6
7yraPOC/IOoG0os9JWedxIOHWO4kHPbm+fVn9QBvmjRMZ8J8QFkkVI/3aDHecMLE
NcQUkJtADJQes/lgELrLtlLilTcv3bS7yDqPqcdoVqHpPBtEcYOJHhVIPsCOZcsJ
/ZXh7nAqYHYe6/Y6Tr6WoIM4T076pXZ4sqsa6Ymkdjb77nsVNEyQ02E7fv2eSk7N
pmxSlBMYqsY5sQobXo/Xj+nSTuxzVC+dCdGww1IOdtQ7V+C/DMNEweSS53DBv83P
IOPsuUlzUTdrto4DMrkbi+JwVkpcDfo/lmi/mbgYwcL24IFgaRzlteLhxbUbAYGf
yb4pGCERwrfDhNB0wv/mwTBSGgnlNZq97D9mnrS+RfhvtHn2xYZIc0OoJ8p2Va5c
copHSLGoJIMX5dpXyYd+hMarTNYKRXpRMhIL3RVDArkkbF9sC++Wi4JgWCduawku
TioZ/bouHtjrru6tCZat/Lpx70PdQw/WQM82/jKbliAb9E9g0QkgHl6YhLYZwnrM
xdg5IGSTQSSqsADy8tE+inMJEi/40+xOsmGo2jAbO57/Phra4oTltXspC/3GM7Fa
U4cVJckzQ0CxllyGECGoLZFFJqASs0FTqkmhCvVKkRR8p8FwO7m+OlYGX2uBVQgR
HFk+/1entRgqjsT0aP/dQZydfp4+VqjwDTDNIET5/GpGnV0jW9vhDtO91MEA7tnz
vLjNk8fxbecWNU7LM+Wcy73vwtmJtkYWjULpbyixTbgaS3kpS7C5PbsuW55IAv5E
8MKnK+UYx4SRwzin8oVItbqPA6KCQuHNBrQDaM0zVNcYaIozFp2t5vr/6YtOFgQG
lxIohyl5r6IFOh4r5VChTq/toQuu1dnBTfo5DWY7EedUTu33HqfhwHeeMtkRS8Hq
Zi0gH9GzFKPVjo6+kDMpcaVM6R7jo4vPhOCl6Ue+43wXITMAlZvnU/T2Aeo6T/JQ
LQ3BHi2sXYnE7DIgP0CyHz6/DA921cm7bNlQ0XgPcwZ0g58Uw2CYcpGvzCsrtY3O
BMSp7AZuVNY1CuiazjF5AbdCldfV98QrGd9IvRBi2rats0mf2cSTcc5TBDhtzt51
YnfbrF35BpiljAKGrl17yWB4Qw8PQY3IUv+bL5IWVjUl95SBikh+5DSD7Wetcm1Q
NezqaaPGj5I9KwnWiwog3nyDrr1uWbeJH9ONuYrow9VsaUvFfQUB4DOFLH5Kn+Es
02AgcKPmcEMvK/wYqr86HNpUzZeAlOmn22wYB8SWuBdaU4YiO1SQkNlnM/kVFd2s
sypv6CH1Evg7TPjp38KPiG/7tleW9H/ll4jE1JIhllllKPYcyLhlwFjhInC8WqPq
7CC/4QVoQponCyYtfSbclsV0X5+lTf4An8ThvrAIJgwSNfXbAVABx0Q6AlQqcAIE
NbrH2VcHzN+cAcPDdfMSZ4UjroVx06Gteq4kYeRsPIom+CpnHVUTs+vVhp9GoOgN
zArpM6FV9eid5mXmLG3HderEexy+DXfYCDE9gRxBQGSKB+LRissEE8HwSJ/q2EKa
HZzEQQrOQNv9D815nRh+Xlr+J+NjrvTVvuCzyQQIX7UGlhUjg849marCKztuY611
cP1p0we1rsk9+7+k3Y0OlvmuLJ99kWgX8crb9rt0UIPTiwPP9KGTs0OboQptN7rs
d1pcP0zUC3PIZCET3P2IhIpPFoexgIeuG27Lxlkau27754u78nqPgvq38wqkA8c9
hpXZPiMOcgmyT1f0GYQ3kPLxzeWiX2WNHl9MF7PblElw4rdBsJMW0Yl7XhdbUzEt
eUy6kpYEjf8cdL9YQt/equr5AfNN4IeopZ1zP92HG5rynF+QgOQZRkvrazjteXIH
V4EI8bHDySnpJLu8i9zL3R4Yu0o3DNj3fCll5NGvojpyva9jMzLQlIQlQCuD6ZA9
Csf5FcDH2QjRa3OckqMG7bfGENiIeZZdBDApHLS9l0khqFsJtyepOhsgBxcPa2iO
KWqdW6IJ6crOPwmexkq0G/e4sESOdSiP6YliT/hut3svZkTuFin8R9BjyUOR+qiF
pKZO40LKRaLijEOEqOj91CHGI/ZSu+uGgKWJM5wQsEUi/jb51vrf3sRmWUSYt3GG
5oUiUK7YwRlrcr8IoE6vpX/JfMd0E8WKwHrC/MqZlcVCI6tGTIVB0mN8rVjQQWfd
VzwVFRwGinIBhyQNeItqbmmbfbmfGwx7Jg22EMXYUGViCtyv67zSk82/QB5Ec9ci
YFa/jFB6hPWIG9r0HCYQ8vRRj4TA4PBIhUoTBGFpfN1YpMvP1JedfWppuKcCOP02
dhI/QEWqHDJdjeW/euFrhcijBIrfyN8MpkuSLr93SoBgl5sW0Yju6kluPjxDqC25
snMUgyp6ZmM0pVl8WkmeFD1oWarxvK/ugwbBaNEyA2J6PGfEGmlLlbEdarVVyiEt
k7sdfo2hQbEjiN3U4ZCPLLL+4kcryPpNjxmu45d+89l3RE5XDRYIxl7ioMAs95Sl
CyRfgsDg3lw6kcLFDD6B4kOQGiewASyk/bIioTx10+AuWLAFM+AHpWsfyjWT03HL
HxwFiOorD6Av6UYdbSlGLN6Opq7M7E2Rbfry2k/TOD4/ZzltgtEXld21xK1jJhvf
2uR9OnPfHWsDxm/zjsSWe2UTge7mxfzH+NjcxvU2fhc8fFjnUI4PEUpmF50ag+bC
QhZI9ri4v36wgCMdxPo0ZjV097fcBzinkCcVZ18DwwH2AAtkGdWcgDbZKkiQHzkE
qqack731AiAWdyLTfPRqztPLS6RUvyyihxnjTPgKl31GQYKqi0524kiVbjGaGpg2
80BPyqTwCx7dELkYjTjkcgleORozRyPctL3XVsdqNMzRmYQ20+JLKJ0AQzeOIF11
G3aD9AwVkNYJYYK8Hrelwvb4EUQLBaSX7hF+a0gRd+i0aWdsBu48oGV+lcZOuha0
d5yq7QvcndSX48uWYGvF8vBwgknUaD8cF8dpBZ69xEy+EaC9zGnxZ0rpjWolcXIR
5oedx7jL/8EmPpm6PjdYp4X3uYbsSiFWDYlTZ9MkJ6/DTpRq1A1dvUUkhRvEb5gt
/IgojP9t2dCANTIJ1QCzUxL6FBqpa9/628vxdSDXN2kHWkCSIpwSGsRPm0cLqUjD
+c4n1ltgmt/XZrgqJl5mE9GRz2YSsprf9CkEjmoucs/EuR7csp0PyEGf3uTW2vJO
cJtmVqakTAy5JTpuqNB4a3qUR0l4FYGNe7SwZHlGMaled15Ab85KBByYOco+YljF
8X9kPwpxo/H1sJSfOAlpdh5MN0pf71Gw/vj+OY0xx+45GbSwQx8xwneWAmNXL5Mm
YgQ9f3e9/WohoqJe2qaoGjq5Jo2OSbGkNJfUwHsnRvmiyBqG5KsMqLky0ty5EGnK
9py7NTHroMNq+BDXKmH9bdUuS0jlCXOpzc4Y8JQyh373nw+5I8opdp5vDyXxloI/
XUMTuxjzvoQP2DZKUdWNiyj+tsqJvxVGNwLRljSvevpee74HPNz/n1WQY52Uih1k
NVxmU2fwMUo0sKUziRN/x+UR05NcthJtNf3AyjZXWIjTAUsH87iVfjjdaDIhVD6N
te0WDUcIPc+Mf1Clgof5hn+zIxhVPxqqqbepJ4Z0rX+uH9MeR/FbkT6BNLWda875
CtJ3F4GstgCzjo8QpVzgE2B9sM1w82F6e5yyvaAFO3rkItFpbmw/p44YTfs+Jo3Z
tXRuTmfrZwsu1a6uDgBFOiqyQVZ6Y7Th3rOTa00xcOHifVUfeUubyXV/03FMTDws
yWb1V9BbdVckRCKHDb+ryFQdlPkI/hO1tMRtV28wtWx+/1L6kK1tJ+FXWpyj4Lcf
HlixDFInoVS0eMrnuj2dxJrcZ5vyCMueA0FXDWpP5fHvzNfq58cJlrwA3wbRvDmt
jjgm5lZoKAEtHqsjRriWF+hZa+L7FDBP/OG6+ATPph57xdTtTyXZ3501amT0KXKS
iL1MEZujF4/mVunMwEgCJkeWNzLU7UZYgBEhJeZCrPD1r5Riv8/x0C94z8dfd/4k
3E1/eAKbJUymtIOkgX0GAYd/NsMZhQs9Vp2MU8k8znK7pLYfdziJeArRos2rLLaF
3YwA/PdAREaT2nVfxmn0+KiaOX5/LSSX9RlvaKihY4BHpivNXIZXTrrstMIzE6mJ
WAk/zliwhdReIJEg51OGE8BjFxDvepeCp+Brc3PzG10Pk7vyLUnw7sKtC9Xdz76n
CVJiNLXlDljo+ASH1GF4SsrQFHrOJVJQwgjtDqRm3EILT466ITYT52Yjr2PV2QyD
pH48vg2GATf6WeEqUqslXN6ygEcHB8bRJk8va/fbLOWgA6usieSYvmzTSKjit1C5
pU2r2BD26vB2Nbi6Yf2Azj7VATTx3UbJ7vBkD5Mby+KCZkEtgLehFgj9Uytic/gM
fjkNkhIFnzPMDfvjOv1GU753qXAQ+x+13eg/xDmI4V+1XE5MiFXvkvqQuZshaoOS
7FfQrXktGb+Crko+D5zo30woejL7W+wCI+eJpsK4EgJb/5HNwJosPJz1hM9Wk8m5
G+rGIsGt0+tTq7Pos1V4CABbMdcZL7amguzjKeg4u5e0by85uaEaKHiKrKfpmglj
DbY4Chr2G+HbBkpI7U+IL10hZ88TaLoigjHkhrt2GBWfPS0YHbktDAmu1tN/l3P3
+1eNQ+ib99Se7mfSVscYCfqRu/bpvIDYf8L9PXE+z8epmM0RREe8/UOyDryjd5sy
Fq6QQfw4q+iG56KD1e6YZhnEr7u7gkqiEO0vN3eKsGPu+5A6uvMf1eY4TYz/aBi1
lIfON95pqdjacnS9F2DQxcqsavy5XTZvOGB+JKKVMdfQpuQc2C7d64Cw0qvxDPKY
hTSxU6+prOOrBn+c5xwsO+1Im7LjbY9n4ZpFZ5XnQtt8JJR8sIrvR9UJ1JJHED+K
81XYZ9vqZjZR6vlpSOnb/Gh0sV5tEFFauRptvFTkslgEL1asTMbNdTO0GtfNAwk3
G4WMsNSVmhHJ1NSKJ62YFQzl9rJzP3XW7Ee0jxK2HsIBhM5dLDbaM4qVUqbe9ddi
lW+8okOo/wnsKjAvkcoPVy2N6hilGlh47Z/AgOpzF8bGOkQa1dCBoNrzAnVkclzL
2CnObsb7q31l32PngNhoayCd6e7e+2k4I7fHLOeDrQVgEB3FvgtN80FKnjwf26L0
YDt23+jn3OhZj/NYfTalQD+aNrz0tzS8UND3E/5R+UbdSp0Oy0+Y3oWASZH/KjTX
tW6AmhxhodF2NHzr4E+5sTT1MFNuD1redlAyuOIhFlX/91TBWbwolR7IPxSzBBcE
88iptN5D1LDcLEtDmRwUXPgnpjdowJdXaUdcT/g9IIL3fNAXJRowIrqiaRVj6BNB
31+zreUCrnKMGQsZOwe+XlLwasIKlUNDqCeGH9WZHl5B9ivwGK+0Ty8FDktBA8t6
vm017WYBrAHR/+48/z3PQXzoKxN71iazysf/Z6Dv6K4R8fwFEsbOcaMg/pxt5ic0
fxysWBcbP5O+FFcKs4W/SFrf4tAKoeVOf16oaOmCiAf9ODQt37pmjf1E+6J9xN75
w3vnqmuNQeKGRIR+2yPLS4+iXR5LxwVgki7GyTw0PGx7WBWny+UWXABLaZ6i+rhV
7q8S6K93flSRC3avOF48RFS6TyrZYvRCI7uHS8xJRnb8EwDKc/atkGazvp7AR/cE
AAO2sV+Y2nPqRy2fBkZRmDOAksAfxWEHczAXSPvLta+ItqoYNRgOwrfadnDQ1LrB
LK2eWR7UTGMKxm1Cfx+n6kbra8DbBkmEjqyd40ucHN1KbMHjXMgbwV0ENJpjI7GQ
z1Kz7yz7Ibl0YR/6gFZVtxtK5x6gYuOOUlTn5PsIFYMZ2WPSXi7kwSlCuNMPgcae
ypaLWDiaFyIT/NaMgLz6IZDucWx/vDs8bo9EfvB7yZDgQoWwzgUlfUBbB2AndzCz
rZhMxVCNMdCVC9H9PA021MHli00xbK6RnBRoZP8dWBnHN+xmIAR+1uHHbX/KRjnp
0md3ot7O+IFmxVtKFjBMgF91J+GD7bReHN8Cp12VFNvXjtK9uhcl+8jMVJ3875x7
vKbkbfXdsrp6r2UyKEEErh5S+WutfshJfC5NowIdQPakQRoXNoZqJ9wwBbmz7XWF
IP5e9fjqmRrt4fi9qmsZ4iRpZZq8AUIdJmB1pMZdTsxsySau0pBhRX5dV++XTMf1
UFmK/22WWnanIHvFDO4v3bhM6W4+rrzLMsBHUizsdlx85BmtIdQLVd5N5EU3c5W+
f39Wa9+4rMUKsOSiE7waYzui9EemNzpq4O7mCP40uf36HK9WIRVQ4qrzVbitHL8H
UkfEFTPa8L3nRhjLqZ0LvJoAsq/9cIwfBs8TVLE/CAKrrbfSFZ0njDCAT+ONLvYI
Fps0sqKKLqZpERV0C2BNjBwbDOP8Aps6qmfEzwkGRskoCBilKNEB5rfG7Lb9Jn43
F98/gkDLDKqLB7xT2x855uQjKBszM45WaxASsBkgQZw6B2Qzdor+m6dUxAzqX3xC
M8kLndaGxmQV51BFX241zd/PrKOTmblEqsyOosekgE+nLfOwYLn9aMJeMP6vjv89
p2YpO22ghCUL40TqQm/9KzQDGfIT0UAKK6uZ4xSeQleHmEL12nkDd4YDkHZqCoGP
/OMu1+X1TA3tsESaKxyP6EmraQfWcJ8iPXSFhQKnvluk8W0GhR/9G95WkwpFgE4T
PJBv0HMK7W6PZE3AlEOT8Yv8/tlUvs0bHZTvRE/jo0l4etLLZBEssjzvV2mA9Do8
i3vkte4xzEYF4PhaZLpSt5+wiyRwaGS8zERfqFuFubGqYLj4AaKKgBP3fTXHiJtp
vqyN3mwrvOa5Eu2ISerKWNXRAWUASPpqcyTc4VQdh1kRGU8/YJGkhmtkamBI2d2l
uEh8/tBr1TM75zLyPU0pU+yr1xI2J52sAH0jZE88nF7qAbKkpips82dgCPX0QIwL
9m9N53rWYs0+iJD7BzpaUODeFRMeDdek8Yk9MxHnpCQgb6MGvVccLmNLG8YUJxA8
RHUuYBUGCee00bK++uF2sqmgnd+6jdK1niqHlfLSe3rYkQO9wyRfN2TKlryxyxqH
0omqweS0w65mVfEWaXLdlNdKx5pOJaoRgT2cxeVISiryxLHBUqMe9j85yPjLiGam
TIqToth9R+c1bLnwLqsA9UrCp0xG+VVRKqd3UCx6TDQgUykKNd6hCXLe+3Y8i1v7
iGs/f3qf/k2D38tXXdaPmnaIYVg2loQeLOqOZNLoCeOKayzLXLfGBz7la5WT+fzW
e0eHNZRMzOUdXoc8peDD/A5in2ZyF6dh3/hJ7jvA5uKVZPeE1kG1LQLmw3kNZss+
CzoI3BxDZP0OOh2MRnOQQi5F20oH4FT+UPuta1Ss7ESv2Ty+kN6HKntdGYWBO2iu
zc9hBGWJQi0ZUXOxponDArqk22igRqTIL3i8hIRWNsjEliDi5hxB6ku61Wp3m6YA
RrcpuTrAUOttzrLtK/gecgT0xu62eaEYripkFCy9nmVQHTAuoXEQFZ4MrUEwWPYP
zOrrU4f1N9NuaaCxwmB6KpzZ4ynHuxFY97ZgOWVfTqBPB5ON8Fl7qyD8OMGMgEWv
TdoZ2Wxx1L10uzxlS2z12sRnuFZ7PG3hRqJA5UAc0KDs7807FVdL5fPZPaskiaTM
cvv8JYw1GfObv/YNJ5r768isnLTKvGPw4iBjDHIc2pmmrJZ79DttMFIxBTsu09rM
hOiQN0whlqq/9vtKdP2QrfPLcP/dcZmpsilJRoR+nEtrvppnPjbcx3wEs/+oKaRx
UwfZa2AKMQx1hrBNKnmi4IZptXISA3umEHfAirY8CESM/NO1gB3PyVilVNxuLLFC
xd+aSxGfneFf3kttp0Cmb7G80DQbh5OG0ZEknIgaEp9SIeUtnmMAP0G+WD5Yfs5Q
K+gHfskRfpW802vA+U+Tto14357iuk2cWsep7gYdqp2d41b9g9Pa0P6+Nro7yr4X
0IkbzSxhe63TzTs4qj0XT4xvJQfWsBEfbyp5B8l6PcE3Dde8f0VP6QtOi9ssEhT7
KBHXtpLgKM6YXwL+MuE/jlusAjblcaJiy7sQcp9aA1w3ZBuUyUTcsUwMcoL3DEk+
pQT4qWx6BMgnv9m7kxMv/Nj/NzE+D4p+XKaU/56ePoKbALgPMruTuuY+VWm2UWFE
Kr5McRrb9T5EBWDRGCq6CcE6A/C2mGGxPZiTXL+7C/Iop0+XeZp9Lh30LsV0in+6
ubv6KYb4d62iwl5WDpKKw2eTG7PNPA3xsjF+oe+ZcX72y1sHcYizIO49MAEV9JVW
WDrIv4E7HZq9RnABqHrUPijIs1dcqf68+HYjm2tpzzgu6Au6i1L2Rqwnp7V/2/3K
vosOewyXFtfPNqQ3zk81p3tWwn7EVMXljV/sMYu86jQXVqNrv1RE6ZA+4EsPQS0O
bvFSJBQgW162fKAuseUztZnfqN/uMi+6c6amh/yvMSlMaZmNAPu78d7ld3gTr3YC
p4ZkYxCD6hrzgMkjN5/B+dWNb9v5JDNArKLS34kQFM+1D90o1RJHw9cWtaLIavRM
3bhZSTegoxCIx+pbr5nZkHxP7vKoSyeTHMPnR4DOwTyKSTzTVtAaMUdadR3mPIId
irzIiPnmZbuG/neFiZsCS9TzN7vXFQF0X+VD1E8DLSN2rMUm3Y1mTNYetsO8GbXn
+5OGYgGgyLr7yBBjTpl6Jp5cV1sQ4eH00ZCVkbnrQpvo6z5KzkFHyAVzz4HhkujL
XGotbpeNdLgsrzy/adrZr434zG6xeEEzJauhUkVUA6tO+qrx9eoNO8UHXuaPmxh+
JdSqs41yBUzo4aSpPBuiFPrPCbws2Lhrqp14UWCxCiaFv1I6oTnt/UFAVUxQSfv5
Kf9EyhXjwYo6H16je6TEfTNcKjfOvyaHykWd8zFUndWyqY1hSwr3JH7+qFTYOscM
fuovmzUDZEcVtD5LAVEU5lgg+x0Ky6aDRKrr8vE7jkrVZC7oY3OcCgykWqN9nJp6
gZ+eonFOM+ik2Su3fm35/hCVnjuZTrZ0P2OnTw25uPhOEH6B+lP2HTeWf6jLV2z8
Tkqs9I4a0IqcIECBp+ypD78xoQFGHE3cWIK98xABl+TOJ6KgnFv59lcJIGw1IVXd
HUZMtOHdnA1h/p2FKUKl5x1wv+TOqk6V0l/ZpQljyuHxo8P61S8VC+LFhy/aj3aK
9SpatQjQK9cooDwM+Bevmf0m8iwC2yny471j1fBg5hLFlbce9x70Y/hQvW4OAD7v
YSVY4dbmDpdxm8Mnjsfga3A18gwEZWmq+IrXhDhw9RGC+KQ9SGn3ycckWaCO7yns
uUZvbbL7hx2v3iYSrg8shz9XNRT/6k/hYo1Id3EJWvt9ZVncsz+y1Nv5S2DLWEmg
TKBtqVWJ4dkbaT+RMaCwieTMn9F/jO051THxfkKQathBfZZLu93kL0fVkKo0udZv
ww5aYHGtWs+2W10by7hDCN3Vk+ALXsqaDvjrD0mfNgnB6MP3Ek6EdgVjeMu4MXJ9
CWD+djF+eaPR17WZWMnEvJBS+uUcPP8WpY0X80By4OvZWrmGC7/SKFiY7IAU+2O8
PHl6S4bFT9HQApZPK3zSxIMk8XLXpcLMXSXb7c74Bz0EctOg2ztS33WAQrgq7M+Q
PB2SWWUqjoVpLEBw6a6FEVsOrczbXtxgGiPOurWWPC/izPmO2bzTTGlEn6H0rYpe
rgrE5YZlQDXhCvBlf7iPOvvzkIe3xDCK0AjPa6wRbfSjJlX/ub4VwNKaQ2q2RvSA
lH2WZ93MwVeQwvmFW2NRLrO95NX1kYj77UEbx/Mbp4FuC4rguMYbzdaiktsnZEmP
auEG+OheFbEzuSraR99sxAPbczuGn5Xa2vBWfPZq+jNih1YkiD1zSMnDa0ZujrG2
HEGZVzzULV1xzERhmJFRciDvl9+ZBzKHRMNZJ7iLdab/giMXA/yyLMvcSNx1elih
+tqVXNh0tO7SSmPEDqA5rza0bMLOjqvul4NEVv/0ZjfsM3Zm/wwu3jXRekJmp0R6
2vPRl7/Ymq4uwlUn4VAgBx+r8ogVqgppx758S2YVVnKRgRpJBi4xp45VWseVHgPh
29fbzEB+4+CPTf4kXoJU+UeiVEwfPwJmYl/tOkW8QzewCMMQ+6xzZeHANWJJNA/4
JajimJSzPAF6lj48WiePASjGQWwee+ijT3VB0Rg3YvZehVuGCpPvHolBVCZ5+Kty
TyeLVA5aPw0cMNOHXvK2BEkwnsjdztoNGQW+JQkxChoTC4Ee18lU0yUhp4uNdmgS
HCOo9UjHgG6zAp5MSHbr0IdB51xEXqYBKuJ4v/OdieW5aw3EJoHoJDCp4vR9rt+9
2VJV5LiDFZfV5Zc1vpWi675WbU30dBatFHeLA++qqw2MeBk9G71hfoCs8jyX4yCV
OP8aBLvLVO4+3VxJH9cQ231JegX2Bl9StXQXxiJrrFgslE9Mx/GkcR5XGNv/tMT9
IF88K8GFl9NNCLLz6samxwoEqC9EKzeRFuEW0ok5BtNBgfakpoCjbLdT+/jh+H0w
8CID3BimdfxkaBEqZWX56A+CXTGjraT300e+ju5VeGTMFMV513ofAKwK/Bt3Nw1s
f+SoqV6FwRtTixZilbS6yK78fyqoT6mkFwGPXQS+EGetZFGmCgCE4qPrl2ka0ve5
/Mnc5BckD9b3UqLyPkW91tAN4ctVBKYzayO6ZLENsDNGKlQEZSR5D8AjOs2n4jSC
LS+mr93oAwglR4tjATYYDESOka9kw6YbNwApx34k3bplxt5CGcXiy13RzxC4Tdoj
5jTLg5FiKNnW28rnH4Eq0ltlUPMrdNwWOpIqNAgI3w8afWw4x2IC8bZtmL6pLUfB
sFku2Ptl9McR3Cb9w+hJMkmk7SpoZ2s7Ss0L+VyCg7xkpWsNmhNk+QY2AHATBglP
WDb+uaXsaoObmuTW1ojIg2mX9xZEj/6OG1JZVy4Q7h175lku2XVcGlR+qaFgc+cJ
K2C+ryVTHLPWnpIixoG0H6k6nQNoIq2b+cwAMDX+vSkomGwLFeMivpNyeeuUIQn/
CvPZPnbxoarixrC40FjChEGxjBoGMCXA2lpcAZi5kyNLLOt195KlRe6ZMQNFAF3Y
NK5cGMsbwcuVj0zZtG2jnd0etbE8KYEzFzLWBJlzHZSMrlKTQzq+axfBchg/6DV+
n+404Kd4nYiDVABwnjhHN7EVplhcPwoH2ZMcpmdeAwOxqVTKnhacHRd4cznnMOG/
Xt+nQRV0x47FPh5GXz6QGM2VArmChGn8mcWDvvn7xcnaFmiWbB6KSh1pr2jyI1s8
wtjRSS8bd0wGxvZrSmdJ0hHxBScJZaQGmYSBXvj185wmbTRGy6OV1Vm7PAWBA94O
Idx1YF9nh6BoU5h9dWSp9IiwjYMfka6Pwc9tJjTJiUw1I79FbQp/ppreB8hyCB/D
3id/piOeedwSOZd0zRUu66y4eY8nt2IlaEp32i/C1alTeMRg+SU7lrb2X5Bg8QzZ
B4qi9GfmbUrWTFL9Ke5wU7vhv0GYCE79kNSGJEjlTb+5bOdcUp2JASfMu441a3qk
gStzSC8X478I2YKGZAJZQiTlEMeXUAbUZjkrKL4TgwSJxo3do499tKSgpzmeKllF
tiFeEsrAXGm5ydzT6fu/K7svz0YR8Jh1oRX8tEYkF32IvXoHOHNSrAP/7n12l4tY
cXx/ptSHbt3zEEUbMCmlrKeRecOcRUd2/Pqxey8wRS8Vd5liTlbn3c1SNucTvX/B
IFLXsCtSy9Y6gAKb23ywrFq8Z0eJLWHBX/0LhiyXhXCBpILaExK5EdHq1xFI/w+N
ob3XmWg+Pea+A8YOKc27lR44VVIsC+fnPqxnx3LxK3ewT6tHxB5Gjt7TkT+nHNF3
vLtCntVHyKMIvauPO4mO8VRfHTi1pH57ugecWy92Js/BsZKAzSdl519YUTvSZ64P
jrLDAqA2IKBNRY4S6Ri8bbey8KDww3bwzr94lx3h4wofSPfCytne6/wBdVPHMjgO
UbYC5oXUFaIKHajY5xsslUSthMn8X7Aa08m9guZprGkfEynvoI0iu5jbhUh9giQ3
M9hLy/9wKYgGAMsLuDXOcyB2gZfZWmacWRZ/2KkBM/l0qLzGT+8tiW+EYYeRQxS1
1imoG2RNT2QGRJEuT/25K2X3BHLHYchEW5+wlKQc6ybqDkm0cPWSZMgOrLb/gnYH
pBDqFTGYRb5QF2esW9mIwgpbafQG4gRHn6XrTEgUwR+j5c/wUrn0tbu4xq5/EN1i
cZv8UyMa+Ra8DTd2hMR9AWvBKDvEv8KYrihqij5EJcSLCkjsG0PSPc0seAeYK/iw
gdHLm5mBiExuuj4wy9kRo16kUkdc5Smsa53hwhAe2Sof/PKwGbDYdKgvP0jO9a+z
6fRTfM+KrYuJ0tlj2tarIolQeQL5JlCiU+eAgihg3IiTg3aBACPfXMnsYxUMkw1q
PsL4WiSFF6xkZn+itkbmt+3lQPv4q3Pb5wgrhO5bDrCRCf0fASm03c4k9Jpq92lS
RxTqB+IHL3+NwmCAZ8+M+UQeBR3btkAKb1+E953ygTUZ+L/GPfD+5Bg9MouCIONI
Iipl9gxesip1f+gf8jy4CwjfXZyMeBTJc+xBU5fQyhqbSwOChQii65gAT7SRcp6P
mMQeAcM2NAepvsB7w9HKqYzuu2Hu7DTvZmePwxeAH8CG3iHub7iM4IYQp5FJg+UM
JNN68EG2Ov7P13N96c0LCG0yfy0Qqola5xDtmBjcF93dUvfG63WBkUmSzQTClpfv
mnNSimfNdt0HKHQWfX/shDobsruHT1n028Cnq5tZhyVIuvqkSMdtwATkNGJGVzg9
lnavK5cCgUigj8kVAdY4hWcnVwwzQafdJNTw0MwvyTrlu8i/qm7IjZ7NnXzSzLOK
G+v25SykUNATSVbfkD3HV29Sp+4Qzu9CAV2oIG58V3ZnBauY3lvOvkLLg7g4WQZB
mXxTGhkRVLUhyFK+JzJNHf9BKj5gWzM4+VudJ7dZ0yOktzQNGXBsjgoNoZjhb2ht
kd/fjGjpY43dHf4NI4vSr1boQsc5XZprWdaaLHKpn7Tjn9wUFT9lI6naTSO1fEfo
iPJBYqDVL++o1qGOCq15mHFA6AZqH4MlL7rXXLg5IX91LlNU0fIPrK3xJyGnMdcw
3HKOqbU4rn6dDcIdPHdM2gyKrhnu81ILk0fCn0jgrbj5+AknZ/BNYc3OWWi3uohQ
pcA6aQsFLFuw3r1s1kyA3VjVkRSO/Lj5rm8kUGTEgERhtYy7NRdAbgWYvymL1zRR
XmXLi4Cjg1+PAM/OhWskI5fVz8ifHh5cZnKy1mRKK4VossbZ+NoLjNoT0/+cqKUr
psFt/5U0yqTSvhtUn/oNdHaZR+s0kOW5HNiQgho6QYHDxS1X3l35daW+UI4F8Xz4
IuAxzjX9wJ10s9dYHDgycFqyzbXsHTM2d2nFLH/uAZxSOU/8kP7tTzfJuYUZkS2/
uiTwBy5SdSFyVrym6CVFHUuS8uDofTs/Sovya/MvdvLscYv7CHkjhUNZp0obfRuz
T7LkdXI3riybuH4rRkmtxJ/bs510BedHXhpeh7kPwuLXxr1/yNoc4TxP9KlsWE5P
/jyDJSPGGEX7F//JVsMA1z/+cxHBcZ4iqMcHbLqyUqeJ05xSKpn72PHNaPQwd6nj
4J19RrL1evywY+GJZQhR53NUsSz9gxQvINI0gRmDH5v9DjzVzUj773U021Ovfgyd
hvkPJH4tDBTXPUN6mdEaGw9uKME5lJDUZRMwwCifdcV12t2p7HATGA6eNQrRwMxf
Ql38XlzNwGOKDiQaxNGERx+fd7J5mzqn3PBO+MOSg57wItoQdajZ7y8jeoCQ+9XK
k25yqVmNjK9owwG4d43+p2A/eeFyr9RpX9nYgequI5YzT7td6dhoElA0hn5WrFFp
iJ1ZKBaXCfR7NlKhbZvXvAPA/fZL4/ZOHgfBgaiAoQlAEtf9XifFQlCM3emMEARF
nuAeiqNEoLmUd8rL41PHx8E3bIGb+7lrdWBZkYd3Q39TUvxOEGWvwG4F6/rJf7ft
rUJqEeM2l3KzBGO9wIAPnUMQhw9t5GXv5gybEmkq8zPqBS8WOHpqlI1F8pxDUnaX
R/YGzjgd2UvhyakloiD0jn0aFU4SPu/mvOeydZ4F6ARYmfSJFxrW226ekpjdsJ6E
ZB0FrmI8Nf/RnWEhbNkD84Z3x5X1N1jaZv7qj/oUP9O1JEqCWSLNl6uJ1J12ISYE
EIdPIjxnhtay0LdvHnuzJ3fvTjKRb9BCYXz4kpNUSfGrqBjL+2Jx3/WpldIk21hY
Kip2HrH7Iu+cIDJva89LUjB1zQG09CXOGvODjK0kriH2PcQm/kGA3w5i+C/6w4rr
mlPGbh1nSTlGIsJR4Bm+zl+/YmM6Piwx+1CpgKeCSU3elqXbWFPoUhyuPLj/eHgw
Q1Y0QqA/V9QuC0v4nhuYjhtLEcmJwH8rIdBTYyFcgfN/MiJtzT4w6hyuLh/Ff4vG
BchkWEahkqfQt5Aw8wWD1q13gn7VCmOdQ3e95309J7BWJFIJFlhk/muhk+mAOJjO
RC+NSW8RzFA5r8W+tAc1BP/xC+7YLOcs3J//MhdZ1P/xlaT10Iyh8LFH+cru4NWc
f3y5YbPsT7dtrKaRvL8xkm2dfffpw0VuNAddi6zPWUptumeQmL+D69WSk2x1ruvd
BN585QLW7oG4QMGJgRNfMfDhNMPCqN7i/JEGas4FptCCo1lNl4H8eSTXgddF4AT1
kvVYXEdE4UJCs9/O4bwoqox/RsDtvQV7U83WeX9YEUI6cjlVOT7RNXxpKCxo/3gd
6B6JVYkM/BvspH7ZQ/TO+LZkqLPKVqbjjr1VuvapBtk0xTwcZ0Q4vQr3vES82yP4
EOOMYlKwL5Y+V9I7lPO/ZOjXY5ci5NVDDmXX/LMJeNuW+LzWAckfOCvCkpZRd5k+
ssWdqCmPdb4DxdNWUhTVEv7i2fHI3wVfcNdczZS2dXFtdduU615Xn+OB1tDVk1n0
J//yjpMN0fQ+wvpU7gkhbD+G3I5aY26ggf5NbGyD7ME9wh/IoTL7s84NrLVE1ODJ
ZAH0nVriq8IZwAKM/aMdufC+mkHQQmGgl/TWAzNMkTcwTUMHn/E9VtIBgmQEVCGg
szrFyRrFmYmAHJ43fRntth8/zmunMUOKJuddaG/ehYK/NJhKrBg/vRu2Y6sY5p4f
BOqq0hQe/eXszcdl9PqaKRfKcF1MvkNHv5iwr3YABh/OdBwDugfTMeL4lpXEYMow
/zMTfavg+EzmCSv9p1TzTWeq1QptMFVvw8udwJAJpEQpBA3ehjAn6XrCfRL048WA
msQAZIQxA4n1W9G99jJlKMXA2V7TlhJkzdOpVkqs61XiPUqHXX+vo1+0VV3pJ+zI
zVHyrvcb4g2jzOH44t9sN8yUPnQyjNuA3gqXpQaLv+KN2WJF665GvjkL9QOFH4bX
MkPsSuGhR5J92TeNaPzPEXqG2/kovs4Jap1rObE6yhPqC6z1tpXr2Nj8eVJqaR/Z
44Yu3Jb9jDsY6qAqrl67oSV1DWlyJPASb17BscJXPbKYvSrulPTEIcYiPBQWXCqS
1h9m6azJnhyuTMTCV3STiRHiZnp7PtTafRi2Ux7/q1vAXm2fF0VPGEwL4tiXmLQv
VsiqzurHGibW7IfB7KVU0CuZrNtVvtyIYh1iQgcPlM45AFxRV6U0KllOsPzVVea9
nTQfIsU4qV2Gp//MIvzqAeXlyQdVx0GUsDec0KJQ3BY8zBXjZJMEuh5IcipgE/94
zqr/D1SYpixBKQBZmN/ljP6nNA9gWdslEie8ZzftIQ3LdccW+MWRevPNtMr/jPqX
2Q0+6xyElsySsH90UXzkZxjur3/7vbudoTppKp0TE1yUBISmc/7mh8ayp2b/jgXX
tna29J46qKKweX3SRSlEUjRIA05ChHOmB+bW47UYMMpJtBVpGTQ/3CxSLDjCLNfS
NSvm97q30E1SQr0MFNJ6F9FKlVxDFRBCns/QNNeRtVWpEKocYfEAt73a289/tYY6
lkB1ONhD7pnaczYZDBEZQOXjWT3k04JyKHiFunJKeXt0ouy6NYWx+JklDozzQf3w
oYq0B+jujs/wm5A9TkUcd+/zbhAcPgePKTFjaDOCigkpz1Jw0HXWFAQ+49DiISB6
rt7fz0/Hc/2y+rWDl2Mma/93NHwFyBFx0RPE2tw9B7YnnnNRoeZpR1Zj612Rg9e2
rTqhSYucNhocqP/aQhZdC9s3AdBJVWZu7IWX45qRVp4ME2wgULkOizXjlWRyft92
vOnrXXTVE3UYek/+oZWQZLxtqQeDggOKAeoJKXSGsOEvLeYznAWWIMEKh2XJgALi
R+N6JhEZDCNpHKI+tuyaVWjHxmL8/GcH9Aa8GEU1lUgrAADWWTwSZrOsVZQ3rA8a
twLgEvC45BNTQD+Dw/mQ9GTdp3pdMlJ0wmtkqB+PonNiJXYY+/RMlTIP60yC0Vek
G4tT0N2atBN+jnAt376/V2vfwuCHPGsd89JDJ4v+CJNb976+kwEs2z+iPLmtXO16
5BjeaKtE2WLUr+uqwKLiN8J5OjH0bgMVTh7m3XkVp67S3O5hTuAx68jTap57NagO
ZFDx4Z6hbyc/83dyFh2dzoFYeo2b28AuVt85hdsBPsd9EcXusNI1g50sNwq+HNQq
7fsCNhpztMb/Wyj5ioAYDxvqeqeYDhXI+yZUa9QyTYA4UP55Zn9Ob9kQVMB1bqbO
QJOg9qj7gs9NDd0Kj+wHd8oOjy7tuD74kRc5cd8e35Gvytau1L8onUa8ruO8cduD
O0Psu+Xio4nW1oA7A31wV1uvUz9irXWd+6oLD2AQTBDbMmVbNEtwho3pLYJzMb5K
jYok2cdt32X7x8Ip9ArispjURpOgeH8htzEWzQQU+fRjZOCmhIW3pfUYBfYKKe5M
k/ENz8azM9iDTeaqQtpd1RCjFbeqOlPTBN+2OxRTr7S7fJjkd8mm1mxYvUL2wzos
Ym3JoyVbe9xmj8mPfGjkzTi3wgqsxoLTeqRzlDK+lvoIB9EDkaCqxdJKKN30TCmi
54QD926vIEazvRNAIG9tAnChz0xSRfxEYX4CDFquiu6ZIcPfOkz6KtiVtmlQbbj7
16s+Ogb6q2UxzTcdUcRtLWma0Qia9ZxLKKoeg5Q4arXzSxV5vjXaL2OmHIqjkAkq
dfhP2HmWxHSPjj8eFyrfHoNudyfpOYozE9fHwkErp7oxOvrQHTYByI383HXP7j6F
fhFWFyVnKPm/sVSqsVS1OxzFUiQmSSHztEJktDbMngkXTwD9fwV7Dgyket20r7MO
lA/lWqJHnx3ljC6ByjCo7mHlHbPXVbN+XIr8scEJBtyVf884WTpQ800deVisGCbj
0mxxibIglEWSU7hiqnPgUMXQno86YpUMlHOFhGFqYXkiSls/z89SYMBb+klrM7YM
8dhzFLzaG7FDyeJWvezduBWp8L0TZ1muAT5EP2baQkZM1vGa4WhqQT5TclWWkZ8A
Ksrpn4/FRKJTCUbqsHBieYipMRQ2/KecXLtTyrHlt2JQqtgqjKFaykAugA3DpmDE
Yv/383WodgOZO1R6tjlYZrPV5Li/rWWTXQCLeUJ7W2e3fQa/hMCu8T+OmGgABwXW
tZnZBdqr0PK5qjDDueGdRqlTeqIjwx9cn9ATbv+FP1vAE/arq0IzDMFXJyAaLZ4R
MQ+twaUUFq1BKidxPcJLvIBtO+zmMTOj1fc5wADrDU8DxodoxlSCqJljGxCufK+I
021wnS6CqIggqL7ctEF9c/NHh/QODNang4lGM0cRCqLV0soA0loJkUveHkF+1Q7b
EJaVi+fQ1/Q+2yD8kPCH1uOAcgBDcJmJtBERZgajR8yf4T5OA+haUUUyKHZUCCMp
nDg3pcsGp5mbldqEfICeZDIPckCXSs0xMsrvSy+Sij315AUgxDW+xLlw5wQOLE7A
nprFSbc4YRBLWZEuk29Obu7WvH2lyUaAzVm/S5Fu8m7Zumf1Fpk4ueIFDw2JwmiP
IKwb2vJIBV5GLS0nQ5CXuDGhs2hG1DxC8qItJJglEAJToMySY5gKreYE0Mb/zeI4
L7qewXNlKvK/uPFOrPKhedACsNymsMv3levuNR06K9XEM2wLMq7Df+ye20P+b+QL
8pjBK/LUd+u+MZpRPM0AQdiIsIiEKCMgTCyZa8gnVrWpb1G8feRAY0qjYTCxZwkj
1XdrjxH/4ozzvsAucXinRWTbPlNbK3strFel71qi2Ugi2CqajzwlJDhy+yITGbPo
EruWVNaOM901924xSOM+VGV5Dxy9xgdbe/M++l22G1+oEfRBX6lKnNek9ylHNKPW
sissaBz5CzgL99axFQ1BMOI8ABgkD6Q4usObFJQcFEmcPgnkl9hb8TrIs4fHXQSQ
0XhoMWyUwhJw28rymWtUWGvNz4jiHknwKRRgdNoQG4ngIYsT9tayUO/o/foGowXS
K7CaG0nkRORu6YC08tTNx2ASmao2DDv8TD0kzJGaSu0Enp4DwMrpHOp0zu7719S7
iprajETvhFSiNFhlCUn2r9h9D9SV87lgLG8dEHINQriQOIASl6cl+pojWTh780gf
oRB2+lYzjEmpZGf5oomIOvGIsqRrW22gjzcO2EXZBCpShZ1T483yQcYmO1iLHqtU
eMW0VHFmISHVWL8B006DCWY2Cdx4IA+QqC2a6oo7cQ3tXyEa6Xn/A4vauvUqaY76
jEreZlM8UiY0OdcuE8OOOskBSzA05Yg6Qhx0QKf2yFmPhhoF87NtGwaO6UjQOHdJ
tCEeOXgRwyLKynnnEhG/J+MvOvvvbNajxb7m3oGL05twM8ySoB120sBVLVnlDHIP
YZbZZeO2iN3K9Ug3dhnXInWyC6jj4b2pChZQqpMoNgIkcBfXnWqsLY+jvS4Uc/mi
Eqv/QHPcCaRXgBqhaCq3vthM5/2apKVNSawmL35WIErVvq5BapvbDs9utlRMwEx7
0Kf+DLkVNG4NwK7ry+9CiXblcfrS4hrZZoCfomw7CJ8g8wfkT1CbZJ8rN80Ac0Hg
ntSlpuyvDxm5E7VlmmfvMU6biwcx4DO9uvwxcTwrup1e9Rn+vef0LVHiqXkJxCwL
baYz/+SekJudnVqoM4is6v0aFXmzq+dRejWRcDR6q3ZQ79RaCQc8p2CPG4OKVabd
lUK0Lx5jwGByyqKc+x1skqaepj1DgZiN8+l4WOBBESefCrv+bogDGLJHEVGVUWmG
fEX8bhPVEQG2q+OQLkPcgSXeypTJkm4jxK5/xOJsgSad9/xJDNUYfNiH5A6ipSh/
Bljia+JhFof+z774bAatydxhfjvmXUq6Eyl34w7Odq4Gbv9/Mg1SdQQmA/fteSH1
6AyzGCRzVcBhcxnf7haMDIZgwQVUEpzrqeUk+l2zukFfsIdzH8dTloqNZfq+AU8t
NLZo8qZaTq0jeWEZxXJUrVKcaK5ldznPmektdXFB0abfYu7I4kxqTrSsqUI8WQL1
05z8jVCovXMdN0aktit6bE2COi/O/SY9hHWt/ks5Pmyt5fS4m9+r7KsWv05cwQR1
8QtXZg4aJLH9HVE1eEnBwp2xEi3GPYQ5tZSJb5jqLIVIDUM/0Ymtdqhtp+QxOJSI
5Y4x+gOfm9DHElG7ODBtXCcbNV7nA5werZ4zjZ7TXGXvpvleJ0321AOrWQ8j+sNE
Uuj/9N+To/7tftnpDRyy2QLoROJkrR9Oh67fXm1V0I0NMP1SuFTmKkperjr8VB40
2XJbbh/sHmsrtPUTeb+cyD6Espk97bTvyaTNDB+AGHX6LWh5iB3QJS0mcvE4nqxP
QNf5sBUTCBKi2qCZPrnHGPXHnU34UTVUYzp6dTO6Uzk2MDvo3V66NnvJpAyOYRYx
Mqhsh7VsgRWiRRl4SCXJD1NLknoe79b+ml1nI0LIO75Mlfnr/OfEGYsWbk+wHD92
FO8RjAsEifQ+ZjENA2xe9Vnvp8bkOzAkDhorfUXZka9TpjP2JwgkII9Il5mEyA85
BJab6OXPidu2VNFTwQShx0KwTAsKax4vYMEq7sXIeNrGvRCFAiEgmiIjdmrFXBKo
xMGw6WdTIvT7uLyUjsB3rvInfZzzkNzTs/4UtW9JgOMNy14h8MOlfHP0lD0ztHHY
k/vdm7ttLlqtbRvyjd9oXW1VgLliVMhG+oBoyFVPcdFw2gMVF6keU37TSrItnuV7
XiseNogeGYYSFrlYMaAwuvLHVACxiGcfLzTtqWVZaGkT2Q1FmZQ2aA0IlyLA6PZQ
674omrcyBKGLLK7Aiz7PaiqzJnA+a5/nczDb91aHNJVIZ3TWp3d8aXHJ1ucrqE/c
JtzlCF6e5/onDoCUbCW4vp5gr96JSRdtiRfZDQqZahNMhpdHDZ2RbCE/RLOT8q5B
3MOr112/V5/VNrB2oH3PFlXlF7fT5MiU/BB5KcF+SiedEsgQEULHDIfTeQy2advX
R0NRjfYBlLfeJBkuNnvuoVQUnXHJ0I7bZDtnHRRwAI2aYefE3FH3Mjrka8OjEiEx
KO0gRM+iid6HPYLX7VT5nq8DN/O/0pbDrDvFXdTUk4mlGlgY6c0h3rl/er1XcX2e
DtA+PuiFJCy1VEIVtAE2A48H56inmuDJTy0XVwdZBuJeE4ga9Qjbd4laiYbv13m1
nZhOzEVT5Lp0dwsm8UsHdjJeDVbbAkuWd48R9B2Xj9tl1BBPp5iRLUuVZ2ZBs9cH
GtteFwpgrYNYOhGCTSFD1njyt6Ra2d6oFh6FPl7JeXErNE8T3GHghIRieUTSzsld
TRL7OUkoQ/XQaoiJ2AhLh0UmJgA9fnPj8M2VfnhwecVMaRW2xMs/wST9kG1Vg3nH
JocdpRI1DQ0qPf5tG9UHGsZ3XtFfRFQNa7aDimmLpU/32vZFgRdfrjq7mq6x4tOl
TPjYIZpgUhd/55GHlDLcB1AICYNbqHKniGR1LA1kgz9YWlesrvLnneavqznI/Na5
e1ONMxSnVCCHoLpN+vaGdEZF8Cjpe8prv9rBmV3angCQeafw6XuFIFPgBThSKwd2
G2gf4555xYD3AE9bxz2lZvGOOKpSSHFBmC8ahWfg3gPXEP58had0Ocb8XiMY3jVJ
SOu7qL4HG2uUaQ7FazdVakxnRpGvJC1UgxUWR9/q2A6nX4x0zrY3kNO/edY9SWHp
f1fRj6koi/5bM5JqFy8jj/FxPGXZOLABFyg1uS5PWTf8vVun3mofMmBQBG6cjCna
2plBrvSTPLE0ZNraSidy8SALka7BwRgUP5cQoctt+DJ5yZg9KSo2PD8gxk7MZm6E
s3wfNsv4Xa0wv658mb9aWyTJP1SY6be6ylLoImQWPVmuL0+aSygBOEBT6g4+pzYG
997zI61crFrDEqd6+UKK76IrsO0wWsKEyAOrWTU8cGVe3GSh3UhhALrYyg9OmH7I
TI/xDjjJSSXUcUfV+oWzMMFhVv02X1OhakcKekerYU+l/fPgf7lekexU6n9UBVW5
9qetsiAeF/jDsFtJTZ469N/JsqPVF3ofB2tNp95FVjOxwXeviekDKW1tL/lEoVFM
8AXxhGF4rQOC3dRKfFY5h8bZC2Zl78PT1qOEmddcQ+Lgi/ooW9y6pFWMDmre/SzQ
q1Aw3f6xIKlDAW6N0EkrUw3EIlPagbzzDwTLhFgrvpRPaZ0mRz6889qSJsZUbM14
2oGWxxKfU4qxzVNZOxjJ4us9VAmn7+Hlq0sLkBulVZTkorBmEqXXWOJId4S5VGW1
AGePclyfPtGxZDQ0drndIzQmLKc1fWhjVWoJ+4CGnUtwIPo32MW3PEhSFaJd3UvX
mU/9K2PNyU0Y6iM58+W0wFFujqkK5NDASo2BkCTheZFvXOTfpxaM1hjkiAWuUpyt
Ln5UP5NexkImMmGZo/fyFsM0cQocovRF0geuY+LQuztg2ujgtV1YlDV9PQmhC3sq
rwRd+4rHmfKwIZewut6MaWYQ+FEYKDI7C2zZYSdcHHuCUbMWBcbXITib2EUgU1l9
op/XhjsxXz2Shqm8cObwqk+fBjUZfZ5eXBGPP+dY3K+YDhmX31lzbCWnGAKEJGa7
FLeHKvzkG9tBycEBhXojIcqImdxXdAoVOUsgbIpmpg9EXkaYsq6tgNJbpcLczp73
G2aUK9HIBXXTa9Uacgfariio8ZQdeBMGnNFlKOIH7RpUsIiKs0v/xtXtASH7y+QB
YwMx+Mw34E3fPFHE7r/lOWGDAxcpgNeSm6LiN5ekFq6Vi4QSrlw9oxJx7LQAClVB
XIEeLYhOn0ho00HGFEhgisrpPVr41DKcugNUg7mymdE9yGM+PCHYm6HjwG7hbL+o
5x+SDfk/pYCju8a270Nl1b9kgWGesxld57ZA99XA0kGB9eu31HItV9eewBqYPusf
6++45IKesOWcNMNeecizAmfwiaoJ08yjESv3nrxgjh6PF85jQcWjTabbffGO+7Cp
V9iQIhu1OgcUzn2LkpNmNlI6kKU2o3h8lqUcrDkmhnr2IZ6lJ0Oy4+9ZPDpDi5bv
/aOliTvN4+z3sniwD/VJW2KYPfGo3WaBC7aecfk3LreFu3SZ7MFXqf7EfyFgG9AU
7q8R1wIkfy+M99PebZlebLna6sJsK7DkgbqzEkX1e9h7nGfqdhUdpQlbgXrmrO7B
JtDhuCXIFl+f3bKcTsnrwznAXek8j2JzmfH92RZ/mTcgdc/QwJ8gMNC1QBPrI9np
8srKLRAuSVl0YN8SYZKN24XXCadi1eBAtUn/EXKF3CF/VPL19p/06bht/Ebdp3L1
xTrQlaQqzI9O6VzgVRdOIFDbAOifTlLPXvxeE3OeZolb2B0nGQ7MSif6M2ekvxmN
ahl9ggjSpUgG+dI7q1Miy16PCPHeeEyPqBfVE74YptAe1YIBiCD6FuKlFyNzH51e
yilqKlYpupHOEYX7kRa8pkl4Vc+FsyRXubkNwt+keBw1F2NHz1rvHYoJCMBBjMya
zKnYV3UKr15J9YF9xGREXeuROong7tvA4V9wylD2TrZNPBr7wvd/PqI/jGF6rZ71
gz6jN7dwy/jvouq2QuhQt9ORfQGK9/iSpM3EOJ8lnk2sfJwI4wFmPnwCqRRYd9o5
W7NGtDhM19eIIWvf+NFVXZemUvPHHmF+a8mgcDJibjq5hQS6QNeZCNSS8s1gTsMm
CWvHRH8/faxG7mRmhQx0H74kE0bD22pIbXmWpr4Adi0hUYQuqoG46rG0VclPi4Z8
SWzuFt2FrYc5JfABXQzoklBI9zARYudzjJmFrwJdHQGcEaRHwnqwtpQHwtdFJKFH
viMmp0sY4WnBG8EWT2fnMOfJJETLt6eIbMlWrGhVa6VpN7JmzE3G94CiJ0S67lnU
7q97L0vkVxfgPmsI8a6fV+D8Ssnln+lypxXLT/4v+eGfgyhlXAbzzUwdgwaOL3g7
wYcuV3672eRTI6KuMr2t0gQSmokUB/M93O3/BRPnCWdR1EqyBsnuhi9ktxNzB2an
0U7V3sbmtugB8JfGGc2CMzqZQskaIYgVBQ8h282xKOADa6b/1eZzSMKyl1kzN/Tl
zDwKZ8DJRZ3I+zCovWJ0sBpENejGYASRo8vvM2Hcx78uvYJNRo8d5R4IwsWKeWG2
+/xzfw2TUrqwLCP6Vz2U5JYEGsRoLr0bbuUiiBvb/23ssswtMmvI/zQD3PzxSm6P
JrG/ODH0tlDAtTGoG5OKk5JQ6Ob/giXgj1XZ6/LjobWzAjTk/zmAb3ZATAxK5Zhl
9Wej6St0xBB8+9y1Nz2iUwGL4PXaXEbhvPFHY0kojFu5YZaIub2zTb72aOqMQQ9g
7uX574QCqTzdKNguH43R55i3BQwr7XlrgxdlXAWnM51SxzEyP93AW/EoixSJP7kr
3LVtSRrLY7Yj9LsdBuc2bJHZ5hn71MoML6fmm+d7ZvDNyc5apqQ0f97mxUDVPorB
97mtVn2O2V5qGn3IvehCysy9ZIH4vpdALB0rjr9V9vyXM8XXtuA1hV+VvbX+gV6C
wMkE6mqgwRoacuvhw7lmhS1n7Z7UivqWy+exrbGXnQUhBXiqdcQhDVe5KLdL/SG9
q47SZpy1SubvCqqRjQvrmiUp5Pbx+QL3bAGCRnUJQULNAOsR84pCONrSlckILI19
TwJMgczmEI3gn86nUZtDQ/i0uNLoTTPYKMkp76DhKdWR6WvCd2gkK09ZUEG9DZeX
9OR+XqloTjylpdkSxdcJ45xg/kPSXKVWUch5D+S58lK05n/2wa1d7uV/sl4vj9qN
NRWCaXwvxOv/FDoG9a8W+8R0QEjfuatoDKd21Gb7Wy7GCHYYPxatJpJnF5fpCrqn
q9vH+gdqQf3p9lFqnnebyJ9y5I9D8puB5zu+XZ5KXdvl9zP5ivxovlnQymj2uaHq
5h9EWyJfh5O0GGKyqz7ZS6m0RTt8/TvAG78t4TM/pMoWYHges5Rpk28ebY4Kz2T5
mAzGf8ZtozW9cRrxinTRwQTGq+mGBIG1n7G8VQuOXIJizUGwnA7HzWFZ1l35iCmc
cL1yXjSd4VepyfJ1Po2Ire/1EU8Rnb0kOW5a8n2ERYtzc/spxzhUD+dNN8v5opox
jNfU1qseiAjeCyEeqCutowi750gDdMg0sXUDw010E/MUdrY2cZdHxC5fAcKeMB/4
o9SaNZJ/oL8XqXRImlYZA/GEaOcwo0Nr9gGwoDxew5efoGEvPEkcJOiqOQ9DDYlE
Zofhg4Xp05qtmgveou/XEEVckLuV4DlErULY2dHPRPRY7Yw9TP2Iuq4wZ3yjMW9q
Mj5/b4x+28ycbWpNnVTyLmK+6WrXQIHsPMYnzM+c9y1TPB6IvELN6yhQK04GXkst
39BXigwZyFBU1xMD4L5faNc5+5G3bOjqmr1oIy0KavmSdMmwUnaT85RvScwgV2ND
/QggX3bF0sUtzUPuTRs8jgknda8wkXjl0ZeCAyZfzyERhpMQRrtdT4txLr4AlE1G
bYmG/9Vnl/mXwQ3BMVwsicDg0cogKAuYYAKG20fjvzdp6tjmRiaJlAkUb49QzxiA
0HJqzzBKCa3q1pa8Y10h2Pd9yE/LJgA7phE9gQ057aL8RWNFiTdIFoTvqMgTOSGU
KBqM5hqBpv3XpaBK50mitoK1Pg6CV2oy8kdaBqOO1/HR80iQSG1a0SR/34F3Mxv+
290+fFBP+f6oJ/jn1wDYvpIuvUHPzOVclSMczYPrvU3tCclAUN6BN5hFnwCLi2aQ
FkJTTRBegtZqOBzqbBAiOlWwBRKewHRRAj5pjAG7q5kIzpaGW0JEco7F2ttszUr4
p52mHKnXs7Y64O2AHId9DDrYvdkMsJqqN9jAQ3CSGpEiuJWUsqqmVaxLmBvHYHwn
DfcWpy/gy/UKhol/WySZumOX/KpvAwpmJVX2VwzOuOCwtRgG6bEmE9a9YHeJeyPS
ldVHqgFqKI6bQOnnPXle4bHPaHBjgAkZ20VzBhsHCofXD+05TUjTya2muXTpr4rK
frGMUxWc3CV7E4s4hJE/lLyk0YLajUjwV2/bcb1+9lZbLwooCJgRhlW5wYA3/fuE
osGZ0CO1NiS6IPa2WlKWZhuLeActaJolm7tbJzRMoIVEOUbVnUCe/vfA+HrxfcgA
j+hz9fcPPYTwdrDuU3uxb9/tujR1z6MkDXCdkYUHhKTR1sLA8SrlwbuxRYjNZqIl
EYYya379q4lpD2WfmzjhZrnzRrmXsckc6QzTiWzdCepfkTb4d1/HEFHYiqLJQYlI
sEJcY0UFmdOFeZnvCCglVIUwYqTiAt+L2GcpAflSE3SLUBX4LhXbz0sN2ozT9kNr
Ccfke5XIsG+VP+pWRUH8lTa2AsfV5V+97q6ddqAUMczXLzluIKuM1olb5aVuMspI
wIgtQd3bfAc8PoHjlk1HgJC4gfcEUOL/kmAa5mNiEYV+w0W3ZeVWfpjszM2g+gEF
plAuh+J8+K3sWODC1CcfqzTHWGCbOOW17UYEQQh1RmQuqKRubDlt9UQOv8RRx1YW
CEuU23ceDsQX4bC9O2qgemZLao1fYsmUmJYbScqqxpST1BiL/iBTg3PU5b+mtykq
AnRAqsfLUgqwP1FzCOG5Hrli/Mv0OGsKf0EzNQSFYC07GYQJT8usLFAe6aUPWMoC
xQQvKOlyg26NV7PLvuAJWv3rDo3Ybl3Zcsg2aY7ibSaX7phYyJjPweOD2RnVn7cT
BWI102BKHu7T7ZsDEVXa+/K/MJw/hHo77MEkKxshGZPlCLe+j4723QtfQ1KXt3hp
txx11DmOslJ1qn5h+o3NyN+u5wZpP9RlpyGVfCp8TPLMFqgPYvbWWU9RvRY7lPNa
xLyu0HNH/zJuCs7WNy+xrqEyCqZO954IsVJhdyelviCbw1XMlsvUXWhwIXBeDDcH
Yqq1fWBAJEaIrI7eFkUiS1Mmiw/I11EBw/IKszKcdr2VEriSTrQV72fvJqh3hn2b
PxSStPBQNq9T1FUN2RvJoxSEOnWQrPdPA9EX0qczfLtqNh594aRaM1rJ98UPd3+s
Wseb/6SzYuZnsPuOBr/Q/3YXUQYQEvugnkjOkqW1jMRQUBUBEoF7oot9GaPOv2Fy
F+0wCSYYES1VxurCHkzheC7/ZPOcKxJiPiCr3B9tFVVxNjpXi1mY0KOe2RbxMYl+
qqyjCD1d0jNaZtRyRzmREoCs2z4R4icDIjhN7+ttWUvd/+KUqj3vuW6nojM71zWY
pDOxxxilWjogA0XNaJYbQcOA/bbVQ6oEixbgNmMRWgNQgwr+VFcngvuhOZ3SRdoS
DnIbIdTuDJbJA0US1JG71Bl6J093TxdQZ2aS6EkaFMn8UJthxET8NoiBjVyhJmCq
2VH3a7i8KM1VUlmKsTyDWV7MwqAglinTF1q4x6AnWf4qzKQav7ADAXAhmJgDGHyF
3tMOlNRm1pGGcHFy//z73kfXYMR7Y/hjmpJyudiaJVyaGXgRbCLkqgeCZUN2QH9F
J+iuJELjcGNfBpaMiWI/PPJOKZGdpdZQrQ8G1AkVFU19q/CUSoGIvM1iEDyHvIZl
vFNnBWuOKrVjV8Z4jmUOlemEsdAuVCSxHTqRdJQqptYo9cJwKqPKA1ikwF540cnC
26FN6Yq0CdtH4M5XALCsql6BXiyJFlENozYfRaMHxya/DT6y7NV6p8p9eaYB6/z5
w5uwj60Q5G3c4rqnX/UVwcrA9Uqiq1BrFELurMIxLbcYZ1xZ/FaB5TlM5SmHrZY6
JXrpZqTNLq+jc9vOGBu145yXanGhoNkf1+RKahINkEXpIhqF2pbVRVS37XdNkgxC
kFAzJNDn5bkjIdKQzlrhRrKZu7pSR2rYZE8jdO1t1EbYm9UtneO3tbpmiE3izuFE
tZNKofv5QW0SnRPNW03HiTHeOyfYg0Qb79lVpw9jyiNcb8yESPnGnl+ZqJyOp88z
ZZfj2En9hh+aS6bqXW4SmlSqQCSrK/tRDdP9/hCRMUfzhrT/l35HHk5o8y85sjlP
iuDGEGrd99yH9Zeya8skwZU6Db0FKWmuqK0CKTnfpJSU5yFIWNwjSMzKYaCkjQEm
p5lsT0MP0/CyR60RJTw0UKg9iJLtBxMVcH7marSdyCvClVXmqcsYTbbFmumbJkaB
B9o2/QR3w98gjzJ00Vx9gpyxiqney5UiPnWGBQnq8tmkaTM/5qoShTWXu1g0/1xb
X8gWnY8EWwHzHrCwq6z8AvAjxqZNX2nxZNguLbKudQHp0rA13xTC4TdJPSQO58Ml
pclCCXLqdRXNXVC5u+T5FJA1ZQK3j1jGjYYjZ2bMQaglamWwP/z+lTfcQnEJMmzv
PGTdxZDgB/phgLqYdclLmSxA54JVG9rtbO3mNjRB06a8N7GcYYorRjaMS+R50snj
nOuGToeypLUWGXLeo6bvvG2JAEjrWwyH6z1KUINTSeucr4F6NNebKBTdoQwYXFFc
WyX9LuK2lvaEPjsNXcwmrxH3eG7ZN46n2Hd3LZZJWn/ZjIX204HzW6pvaSHDOvqk
lEk75wKW8QX721K8e7eRKnT9qnKTiuBLBRWw1NJmUi0MkRkvcnv2cgSa3jUtZDWI
YxQG50aXN8ZUghrS6rK3IoPYhjniwhwK4EyyLl/vZb80h68dp94QZQBtvnlWXh4g
tDfxyBcc9GOjWTQusC6Dni20dtnY0qQ+AfU+V8TYrNRG8Ovawk+CGGp5fZF8nKA8
SMGWV21CWL+PpAoH2NjpPu4hf8wL6hpzS+m6rQh89pRJLCX41RdIz77xV07AAzk8
1sG2EJ1TAmprBf5LlhfVKEPI6xo9BEoAT7GR2lx7/InY/bWQqymelFvo8ak5QVCo
ZoLgd4Wii6Sb0OjQ4/lLWbFK+rEErmexY3FSaNwPU+5nKZTLTLd6rawI7/EGvl8M
62XCJmrN6rWf13ZStSoMur7a9l6dce+H+EknH7SOwJTync8Ie5piBCWUY07EQIn3
jB53XNiPGuqI6yp2KZq2sG2si4PgZG6yxGWm9B3KSsyWdhl3nQFK8JrA0MeHn3Ri
XSl/3IPQayF6UTSNCGo6utTn81gsZPQN38C8fzXDvrqCjFPKo1+iTYNyYHiJ52kh
dETqCvU706oLFUkB5caw6GNsjcRP4SghMzBQkMGN1Pu9zCjseVXoIRmEu41/B4yw
2PdgdG41CPBOgkd7qUOxtLwd6OTdF3qayLmeXJvicixQkvOK6W/2OzIPbXhL0OgQ
f774hmde4gZMkf9SAY9q/HLGN2OMQOmnjbERXuy4K7kxLAtUpV3DZc01gL2l3x5C
LFz2RHNxgU/FX7f3ZNWTcb8LENGUu+lopT0SPUn+Dp8SqSYDUmzxJPGaLiLPhHoc
T/Z6OOkGyRDS48Q2WfTgiwjR5sECq1QMDhe5eT5Pfc6ytndyTOntDZLwcu5eDT0/
kwS1cPy2TDqyp46XBpq72gDV+Fc4ehUrRsi7Y8jq8Z2Wx8I5euiNE7Vlljtn9tXm
4pfYWkGV62rFyOIEKIWqcAbFyxjJJMfRwWSvggUGjhj29sIevVv7n2QzO2kYobv9
uzZ5zQsK/5fZyARjucVJ9ERYt36SxdrVAeQc10SKwiggZ5pLUMb59DbpB++NS2xT
19rYD3G+OTCrZSJhjIUy/DF2+BFnqyonaIvrbqLzwES/1eX3xwaCO6CKYY824t7m
hlFb5+H6BbQiOttF4RP8omO5CwGGd5XDEg34UqMPJpHw5fvTlngGP80lsknp256X
Dj0lal/0ERy9weA97Kak2CPxZUlMgd3qH+mV8BpVABPaf6U2jfSebrbkPZDqc8uE
2wRaKxp1BnCn2Y089Q2vO6nWfXWBGVYEASQhIlZjYqIad2Ff1R7yAuqgXxFOc7yq
XiUG4pfOt8B3dAoP8bRrcYj9tFNO08De0qEh2P6asa+NcK8ErVF2je5fAt7Ooa4b
4Ckj9QJOnoshO9zyOxIcaZHM160n/eDpI6WF5GPX4ig5KDDdnJmi7kSJy+Xu4VnF
WZLxenk9AGxTQDjo4XCJ+TDpEk4P6NeAWyJIiOEJDtcpd8Pn1nBlxSZZib3+dLev
crw2cJmavAsDZLRPV2wS05mniI4cgJsKJn4bCNdc4JCGIGWx1SNdSAv1EM5fYdsu
+v0jdTxnfQVFeNBsW1DvDWUsU+tiROS+swlNCEqPfvd5y3QBbGjsFBvn28To3KDN
+Z98Te0pUBU0+7ShHzc1TNKLpPOc7Lf+SQOVSnDPxV64XP73cO8SETZUL4lyifwv
Vz7ahBSc1WJ3odljy3TZfyT4szkwkUFNvzwTA1aGvFePdYc2n49Bqr1KIl4+Wu7b
QcnHMSDMROV8do0pILgT6gUDm7wrm8PiWh+4in0nWQZgoRGNWz86ZhebP6xzGtkI
CpL6sEt15LfPc91c79YQfejttanLbCWimOXFHbgXHsHsqDoittiS8D1umGS6WCOz
gXMWJhXIX9LB5GuLBBYVfv++47xOPscEjcR0YP3LGlO5WaPTSO8KrWMor7UTYHvc
4uGx02AgjR5fM3uce8eJd6orlOr4Ze23A3uxeKK4LE9SgVFEfUC/INx15KgcsynA
bnyBD596aJPf2W0JmZ4QNwznMS2tW0HZzLQ1Xwcr1m6jsKWPHDU4HovrwtLvjgGk
QAOKpHuPvuL0SEm1BHVg3eXd9EqvT19n5Z9a4GvG3i6GMoHL+j8CJvsdrmDhtcH7
D4sc0dEbpic8we2azPK66D6BBLfhcThlSzTboduwgxDIsGGL2zUbzTHroD6VjvbC
s3wSe/u/Y07uL9G4cvhljc9BTnD2H/7sVfv2b74QBf6kOxbRFarliXAoLjSppUpP
xjdJWDuH7TJ5pjNzyKjfdGzBuOVAYwAlDTRiVrN/rNhqhbnA+DTwwjAoipHVgtFG
eCz5KLLZBC5l4izIvWHiCZSoytynmApPKdr6KCGXPFXIs6dda3yNKb6bW4Kjx0uj
r2qz62qpYj5JiUPWpJZLLtDjByJqQbXRgmMbLYF28EBO8Nu58Gxf2Lddtn6dtZd6
leq1go3c13DTmUoBMemFG1fqNIWSVLuLMUpIPM2dCb+ZM0aIlb/VRYneigo46sR/
9tIKM4/B7BEL109I+mAllbS4F/MnjAXpnhHi/AfZUIMnSA8t4S3qIBtQhwZLMZLX
bWvPEodeCLzm1kRNSottGN4ZUOdxsgrYcKJb8e472dBftZzt4dybiQCvaE2eZbBg
1d3TipWo7ctZldWRtIfrk96qTUHw1jAdAuS+i48eq2hRf1gCbXaa1TfOlfa8KPyM
a6cNeLXcuh6yvQZ3LAwAmjId3eJw6b46onU3p2lHMEJbogayZrKlpKEZy7QHC05u
SIlTs/YBxEe0yXzA/HlXSrE2kiT+MM3e38SGafx592il9FkMK6gyHf/0phUVvOSv
QbIPzvhxJJ2vIIFDs8kllh7IqBs/HYPNJ8ovNN8DvoPJwcmOoH0AsGgJW40Ms8fV
s+wqW8flsD9tbVZUQoxbm5c6O5jdwgCzFnzEY/jWK1tMbbjboMo0l8ULqP+PuOBS
DGlpWweSQib1A7W8fQ70Nh4zqWOn4/1WXpur+pAojE4szTJnUPZG4UMj9RLLldXj
MUBWjyAYLDHfHFEYUAG+vgGgqOkxJXRnwh+prei4N1ChO5UizCLlesDbhoYfxjA5
1vb8PFvJmFWldtQX64FurD8TUlfE1mB4/A7HQ6HLxfvB56BHEdxJDpVoqd/xCHtc
vvk5jrhONtwdPo6QP9GlwYP+7dbO9XeMOJT7439OBh/5yNpt4lxoAlTwo8QA/2y/
4Ers0rWt2Q8rZDaRxxdG7c1+2d9P4GGNLEHAavomrNuXMNQ8AMk56eYxBWXZ1L0K
VSOgDZ/2x23EOG1qnbJk7wTJHtrWrzBEdcPqWrdq7pxXl2dV5GY+46gwW3f7OVQo
9ULnNoMprPq4f0QXdb92t8gHs4KH6x424z97A529OPRTlQ0goHf/qeKEDHqDT4r5
lhcM8/N0IRZNJoiGQv9Chaiah0cgEQgT4m8SfH4RvJKhRd5i0cC+pxuiodatea0v
dXcA+N+bKlT/1RiWk7ySoBFnxP6WlWG/zJlboOQ9QgG31U4CratcuJ4lbAHXG0jw
k3gnhkqYlXWTt61qGXOMvwIrql+ilx0sswjOa51fzATKgo5p56OvaloYp5oR2aDJ
GX9QFFyNr/bSVtOlZ+e1pNBWHB9hzHXhlEZNPIEEQH2rHPFt0zIpVADC3IXdjRUw
2RS/m8hWo2DWWygthECqU76v35ERU5ziCkWd43NSuPAJRhgUwyGiu1hTZNx9Y3Jk
okr/eHZfEExyhmwsM8jjCPt99dnmbuc3xHbH6474prqEQOUZbXZ/lBVz09J104I/
+L6Jq2PClppqeVqenrb+kfVryCI0N9SNXp+YO28OlZB2sRFHxrLnr082GtI7vXkm
5O+83p9pLgFHjH2ZsIXEUo721GHTFyMztaxAg87tZ12KXD+wkZWDU+mbUj6iSsVF
3T0moPcbe9nOJvb9wAJuFruqp2p4Zqchc1b79B6CU3XnrVCIuQEEsiOFqroAcBIw
440YV4c8x5Tfx/U6h9E+3qVWu2whks5JLvi5YbVGYxWVxMSiLF1Rkljp1W2v+y6M
Kx+gU2psSxffvJKDB1KiMXruxOpcUdLHO9ru4+Ac+0BJdTmBtqNj0Mgw2cB9Huc4
ahxsHFWQJl4In3ghQjqiciUHvDpVo0O6Yly1qxFifB2o0pzr5TCRkUvRYOJF+9I+
Jq+5EFGUaXwjjYwZyASL7Y2B+JB6nS+FvOOdEPtiAr+0cIUTYSnK97oX35e+Ondq
lhuAoUFs8Bu88FymyQu5CX6WM1IfDfawB/fOvU2EGY/aEDAt9BuZAZ3bwj1icVPN
2Xr8AEIIk5cS/mtaqZlA8oxQ5o/3tVPZhb2zzUFBCdA1qTbBPageqEMVCJfTiGlt
5pVRZf7uYhwbcl6zeuxArfcZUTnDlPQ+SPGBApGarcc7EKscoJBYOpXfIuNEAZ7M
HBczN99Io6Ia5EpqWM85t5T23JHkM1rQnEkzUgV+YkynIbQFuc408rA/Np7EOZCO
pUxJ0vgOR5CYB9uRvdQpY/Jzde8dJ4SkDkSmM+dTQ41BRuIeVezZHFBO528deqiP
huQt6OPMNnAUxrV6uu5sV3sK/WxA1TPIA/yZgK7jKCYJOeuFD4GJmHUbFBSoOKhM
/E591mrJdNBbcGxqqsKVkNXyGQZ4jpaMD7JDMozzC7J0HO7m730NmgjsDzN4KtbW
Jqv81CnXJRDbI+nLkFpEUID/W5fgjxErUycBTPwSkFcehwLZ2ACM1dHKXFJqyZ87
byVkOWgbOQSuu42RRzyYAt1K2TYZaIrTQ7njIOtK5akjmUPt7AHs0SE9dk16x0M8
YMFsXIj71dSj18Bs6FOZz69nKVlq7azq2s9j0B8DmQIUq0fUHeIbOm/b/T02Q5rs
FN+yiUpP65Vxs9r+m24afXVVpEJTQ2Aaur1M6JMwDwqw2nmRhANkwlP/iWiuP5Yh
bclDl5LBYF/nFc+K5H7uyV4vYtVj3m2c3kbblM3o2xP3zH7BTHPGj5J/HLm2tdM3
lUyr977JkCgwEvCUXizNRnuC5R+2ChhXY269947kG66SriVgxOPj/x1Mv3XtCwxc
7p1s2AA5zhu3xi5VnggtMmgAq1JhbZbl5ZwT3nQIkRUUfJ8Cdq6RDLHS09OqVjkq
7pMD1OAkxhvT5iEXBDVonlyIvkC0rTg6haTUdivPhs52nrU67zOQScf6a8cgnERy
mGqnLpGkacZI0SfB6w/18Pe1TFMCMPlKW8gyWlms9iXs/whmYpSd2fxvdBaf6C1r
jTTr940Sp9oudc273Am7VDANARQurImCAJcGTUdkwWfgR8mxI49geHXwdqQqjCUr
sbHrnR5a2s2w/HmTIhOFQ92DU5TLBUd/dfDMofcVoWJjoqwlBNk+OSWIY3ZF/0o5
Q5BGbpp/t9Sw7EP7kOqSf/KYmNud5P6Ytl83SykT2jI221pvN9b3S/C0FwSnXgkV
xpKydt2lPUC69oIaxnQleP4eXP8rgWpyAT8++v7U7ro+qhHbVG+mbJtrA8oBz9VW
6HmvuCipHkuWaRJxRJnj/5ODoqUCydxskv7uQ2eNGHUFvQcu0iOLF1uVFV+kP9Mv
l7SoZI/a497ij8ugl7UoyLWVRVx2zHx97xBwTHS59ZSu7wHlrktHGyYXCKuIYioR
NxiBb75/wfIWgMeJCL7qrtLXKK3QfdH/hYMSOKaJqbxGMb2AH8PjK0yeeu6RvxUz
WOP9KdGgtaNg74YgTDeV0P40G55aVh5Kbwl2p3ivPgbY8VWDBLfS+CY0xiwL7eGT
EtJH5XZQofU3FQWKrgu0hipSRqo2uqd8vKuhz9cAug+BYUXWlaUoGEjOfMc9/THV
l2KFAQatwDdtLTt1xEmQUiay0HRGVuqvlpZ3gAlZ+JBbIG6g/+SgGQlwFmPcEDCM
m5fyIgaWc56t0LK7W0s2cxVXMQGVBhqrcDZmjYFs/gDSiFQU3PcGPVxDJSa0x7NM
/OVQ5cevyDe9/0iqWfgquilCCGAMh2lKJiCsUEIXGO/D84MojSWmol2IMnhfvCml
/dCPy5nugTILdveZ9GdQQGZaVIP/BvJMQPgxSIL456CZJo03P/kJ3m50r0rrjk3q
MVGUjSjU1oyzaaYXmhtVeTWqZ9gWS/jirPcSjIIDjdTv4L/JduKMez9WNvoMmV7G
tCpmfu/hDHwwg9d0wTPlKyzk0jZ4p3ARVuHGtCEUjoY4BFywEJ0kSA7OXi4ND8E7
cUcT+9CsFj8PxacxsU5zJX9z3T7v0XWGnegEIPJWUVAePlWdGxkxuQQVXERHxru2
Zox/O395UR8S8Q2gE94HuJWrCBjwqvKKHBh6OVo7kYdCisWJLXdbH54ATF2icZsi
rrsMzqGnNuo1uX5Z5Y3mWdO9RivzLK7/kODLEzxdCyOiCWHI1WYiP/mlQU35R/Tf
JKYrKq+8UqGEA1fnPDnvBQ0QyOjaO9euf/RNoBjGj4OqnB+pYp56cB0WpraJztKR
AInaeoJAx8+B+Dq7GX7aBO+4e0QxhrPPqFs61lsCMx7ue0WPJAE0vkik1hGqVMuR
2w91BsnUWU6+fAUFEp4NFs1BuzSk1ovLHkxwihW9t6XH2m4rmEvvm3b1+Fg9+0oo
aaWRHSuCcdHMTdP0tvl4FOPdkxAQeumTUBo/zEdvtBF1/4NSdeP+1HY++TViNLFq
5AwlLlgJWrQdt7/Au9nK2YDSXW+NxVYJZuvFGl7p6SpdKpOx05QAHpaMrmWazxn7
HAg9IF9fe62oqzZPpwDCy3Vakz4y61LIj46NuG7ypz9XaX+OwcHbhCGQ6wh5bQd6
kGS9N5W48R7w1mgtj46Q3n11MmtPE7broN4OfLwKQIZHVbeZubu49NKDUmMDVO6z
FZifwdOWAELLIOdkxxv8X3w6X3UbfnozjRBJMzuyc1WbPgKdwAYgrn2b8dDGhHO3
sW9cz57jJBYQqAxwDJkbdFF4lFgvKoyjxLte5umII/U+nKE2UrHDlqUoEiPrDTD5
5GX2EZx3kTyGhoFGijA79aRp+2nEx5bfwPfZJ+LIXDlOHcWJSgSLQeWcB1snLG/q
cAGWgwtZLQ3PqJDqKc9jcMMTj62Z7p/vtI3asVfsh85YIc1+223/gRPKeTR2u9TD
NLVs3RpnnCQh7A6+hE7gjG2+hL2Hl54xBUhmthgtXrEpl72PXmr7Xa3KKoCKu+sR
3EuHLWqrsD+pPT94xocEiGRtBC1IaJseOm+wUWhwyO888NbQbijDClW1D9uj/QoL
2Yw2NXFehZ32Ksm59H8EQw54EvgPjwZZ5Zg+0I1z4m9hdgLrsm4EkNiA15XkGirb
uGlMx5F4r+uOtCwGQK62zXR9zHpU9df/c8WdxMQfskwwrNNoWX/+iltawrFYzd7o
BFbcLWfqdkW874U5SDtGgNwLz3tvKobRv8jMe7W1Ce0vroM7s+3IgiVpcjEtPn37
seSGH5ufLRNaaP8uKzDeKx4LhLWNisLwhKbI/RipRs9IXGEkKZNgMouTfE7yY2WI
abEBzGRSCBzfdi5Wtrmw5NOzrGe0dl8ze43ujhf7JUN3vjbjMikCWaFTCpXgIYoT
oVW28wVUa91KvOUjW5S8Ye1pEt6BxN9mFw/cEbJcXFMQaAQrBBBJVM6U/pnfiLTO
JEjmePD/E/WZl7J56Jy4bm7gDv/3/V37BtNDp/kwPr8KMCFx74NMj8WpFuPrHnEg
L93zdyVvlcS++HN4NhBCt8CuKdFXc2sLFzQWjtdfErt0GaLhESGGuvGqPu9/eeKt
mI6ux5l6GZ+h0zB+zv/yZXVP67nwjd7N/EdLvwRfBEWV0NTrjlCr4nvmCYVqSrtu
kBuGywrQID7eYqjcJqEyye2iucvf643C9qkcuz2pPUO0naNee34anaqi3Rwzydd/
Tu3esW1usDMJRJX32x8Jw/iR+97/eRFlyxCCwsVu6M4yI/ktvnncs9I3qB4YjDZb
px7u2lq3fKJBGG5ZmLMG98H6c9eg10gNM/35tLu9LudlfuQdgjI9kJByZ4HAo11e
AtST7r7LLAwH/HG3CTp/Ok2Fw+k3LAtwl1fFCWrNR6pWH+HAZeiQ/EfWWRMqKwby
w0guyHHyLAqHHh6vUzTjnonPQEDnrvX3xN0amEKT8JgocXvxXoTR8N8fxpKX7+cA
TXp+/EL/GR7SqPBkZQNkMFIXgbkkH/Rzii1ndWtKcg73sychftryYb/xIZPKkjif
5WFdIHQplCKcBfzz1RDGdlQRouNMb3PB05SoB4L9rghBs97OvRekXxwsdg9OYJNE
jFkoW0PspuhJt75Tho33HsxJwl3Kt/ylIpPqvYWaHZXssuesYjWZI3lLGgjqlQoC
R/kunZTAmDOqoOJZVjYOb5Bw0H6iKqi2IhJ0oUhKabaHz7hSgia4oMzLqz5QT0jL
zPW5RtM/+xFlcHM4dtTjoTWVRq71aWojjiJSrM4/Wh0u1N/rx4Wa549fVvEMlp6/
9dkUm1NPph6WGaKa8qMnFOEpDNmfrGNg+RneHzGyuLjAC1qMMOZbxzw83EclGg0S
behE8udrHeltNnxWm0PRxqEZd1Kx2Z6UwtOnnInd2/mn1f+BUAuqVyA9FH83DH08
3Nc0ca63ZnID7HoCIza3TWHLTyJAKGdmGwV8Mb9tT5o+1RCWdztKHDGnXtVDB8WZ
GEMT1Salon21yu+C9iD+UVAAkf/GsXS8GZQ8HQ9/b0ved+0pmZoZrMGviirsBe7X
6T+VGKbvfzrUuIMNxVicAKCQYRJahgcxHnb2I/Q1m1VFn+J57xiHl4hNtXmknbyQ
v1zN+VSeSKsZJai5FMyWlbAcFn6/Lf4QTeG9QetuNNf1xN5Bc89haAWkIgVuBQHv
QGnutwnXvt5gYmpKFVgqldqSonax1mWBdOCHW8fmX39dXfeKg7Wyc2I97HiLx8Vw
usBiTrTebLMX/bHrIZujjDVv/QspWScInZ9C5lD6epzcaGiOQlKl9GsyFllPRD5/
Mvq5wNlK+tLFlnWVAqxLlw4ISOt3apnGLj45M41ckHqaK07ZxAA761QrfCqNbWz5
FVZyXFyXitOn0hdZpmcgxOL1WaB8i6qydC70YcejhZ1jXVJNGaMa1w+xQlo26LUy
384hGNB1/Dac7TDCSitcQlk+Ia3oYZIobwG5rMTPJjQ7jUGRiZ8ZeKlRh8NBv9xi
28dMC2UEQM72wrTqzS7HJYFTC9qLQqZXEh76Sg/JF/YrfvIefHVTztE5dX/ft5eI
vXBoyFWz3NVSyABur/Px2irYqeUGN50hx3HBd0wfF0eewaBeJaX/vOFcyEIpzh3v
WmEySD4dIk5VdkvCNyx9LNRBNYsD5Q+yR5/hrnbjpRTfVvrmzf4gGtN5nuQCLlPC
p7WuVMB1fU2B6AdHPbPpvb83mWq9k2jZhzyMecQWHsFfV5RYjtmfzKCUWNVPme2y
iN0k7jyYXsWo+PV6MQKx/q4IDjQZxMHS8TZIZhz5XSIkmsqsXPLiPZwb+giuQHwA
WCfBVeQvRyvKxMQ3WZ7dRJFAQExwW4qq1Q8seyv5YyX4rkaJMpB9iVL/8IfA2Vz5
yAjP3/X7Zjl7w89Y8bWxCYfia94gHEoil9yRwlEeyyWA4lwf7nqDPtCtCNOR7U44
rFWwjMZrJmX7R6WUApwxE9FVUN2OK+jnUVAs77xV+0uokjGLwaaETXqzm3F7XjBF
PG61LzgNk4+FVrSPyXoTAtn4wKFKydMLB/gbliC2GeDAmr2l9V2m/fGm2+MfOQkW
S/BDJssFMwoR+nTW6hJAk60cZuXyE7/FhSmAwiTd8tCqfpZJ0lTxZL6jkNyupLNN
IBe26rNB0Ol/UjT/K/12ZfmfpNagE3taW6enpG7A7qPpJ6/PZvBvxChh7Bu+oksb
lJcMjUqMSkk817pQEfEPl/o1XdWOXk7LWqCkN8Q0xgDIRnONLTKJYMPp5V8XNAO0
4ga1drhDAvw0jB8gwQMuyyV3jka+Hzu/vOhjtRwSrmQIDSwLo3O01Lb4z6uDkWbd
VFQdwM7pUQgDsYZPiUKE54ZeKsrgR4mXlmrpM1mPTcPWXDk33D3nLZqfbGQOvjup
ICpuWJth8OjPYgz5nc8Ky83itQewnT9oZ1FND/DnWdA0lpDmgN8WY8HyY3ANq5h5
4ejz99lcEfO23FL8Qn9ECEaod0WIgBuD2jJ20wLZcbCILfFHmifcud92hb5EGZRW
BY5j5bL95gKB3HctPNzNJGkCdgvktwZNuRQBuca7NXY/mlujG/xQq+7QYrzCvu4f
+xKOaNea5+3TH12kN2IsIChBDreicLTBkin1wKgDYkQVBdZD09LZWOfrfoSYJIy7
iGfQ3/VeZm+2jsVD5zBPekUuW40vBKasRqm0bzyg504w2DH/xABHyDciSu3OSfpS
nPdozhgUODy1xufHugTjR73BeDpdovchnm6/lqCgQhPt4ahnrCwaksqKXSJwQLN0
YVV4Aqg/qvDzjrtrjpD3vFZz2k3H1ys+Cm29w+JzZFLxwkD6B02zMZMI5oAYx1dv
Slss/OLOkT8EYl0fNi6Y4SKxf0GknnNycbKS9PbUJYj+KLdEiONAh7ahrGr1LBo9
SQDo+Xs7l7ZuWazZdNPxcEgAssMZNEQ9zsOfEy0Tn1RaoCAmR1FTn7E0K5XAcMqn
wkmNMxn2LvLgLla52DUglyMvEe+fvHGDA5swC86k6oFqJM9YjMGlZEC1Tkekw0b3
qcZ80Copmz6fiN1zGECIYa+AOlLRuH8cgUUqNMJtSuLYE+Dc6aMgyxIokM+YI6bv
DxHk6LIm1A34pSzsFoPhCZGib/JnNbDyAHCJtdIowdEI89mw67qiHrQpU31XeXuF
XGC7nP4rPGP117LblJKDpKjzSeB6jG0+krf4lqW03+bNjLJUOoZz6ILG5J2N5OCz
dhf1NNaj+6/0UkknRohR4cby/nm5RNDF5AWzMxUV+BMd0lcTGJ3Gky3qhIKSAiMD
mUd/DzCKXpAVuh2Aq5H9/OuoZ16OKijiIfv90n2XXKouC/GqVbtxh/VdVH3Nn3Bk
kjzZEc5sxr+jP/70jzGycUpxM2TE7CKl7nR3yhm8cGCrwka9QpDUyNt01Nfh4hhF
38I1HwQMtQKMcFPpxSrlqDIzqsmO3WUs3ltvSr958MTzF7fj1rfYiv+re0e/pQ4x
h/Ep1A+FlbGeuF7FGoMy9TX3Xz3PpL0eIvQnaAmIZ0jCo45lzuTg9GmNGg9vG9kI
4V8ERF7/IMJUL5rp2cQ4upX0Afd326p3m2x+u6hhpmlsGpMo3PBy61Gs8A73jmMb
eWX9brXHIc0V/IM2OEjGoqZ/vHHL440I3Eyj655MiBCOTfGVab6KSnbWlLYVq7D6
LALVhNVcp/h0MtuYrHgrrQH2smqdXSqvT7XAE6YDazErCJlzxT5GLEgoukiFNXpP
P5rmy24BYCCTKkqtazdDHjA2GBELDDcVLtrquNS+uAbVxNU1XX8N/gYrhCppPFAH
wxQJmPzy0HLYMkK8YTUGbSvRCYPNJ8nmsYV+Sn9jKbJNSa2zf1vnmZ1mvXafMzYe
2oBhz90Ni3GrzhTj8sBLbxMSuPjWnMEnFzE1TCmcpG42jq68xVMEg64KRp4lfmRb
azTwPGeJ+YqBp/0XfyqW+urtW0W6Jee+/J4zPZZcbOMLPMdBbLXeLJaoZbJokF2N
jWmxHX6Ab5RWuTPXPuLAtbZ4p7CramHEuTPk8fyLjAWUaZrO2hmWA8n6n+GU0QUo
08osicY8ZS97ZG9kUQmmyK4KrLQQErwYNO1tQTcjukCW63POLGT3ycT9AOBZLnFl
xuwDeP/dCjbOxyC+rzaayPVx4BGO0k+rbr9xe3pbVbjrolriYGYjZ0SrOWXPMMwZ
XCfC9woM+r4CMOkCkt0VkYyPGWVsfVymZ4s7/LoDBeKk+0/lix8zBzleuSrVXSHk
SfzKuEnKF7wDZhvfU53H5Qn2ec58IrgVf3erOtqp3YjkhPr4jjZqq9CUhCEfHWQx
A17de1W7RZEvR7IZzk0P2XLnVx1Y34wsoAsPxw3FgDPx5kJC/hjPA8CzZX/RtYgC
RqZTVLiJBHoYADQFJF7mY/BmuOS1A1oTpyMo/lqP4EpdwC+bq9DroJspMQbLmrB5
XRdVgcgWpvR52UVasxgpwpMmWrDSDTRugJKAL7SiYKfWYKS+f17f0A7v4aIwIMg4
/OGeer+ZkbkocpqheCSmh0momagwiseHcKSkyOhjP1XBlD2nqO7esrrKjynRFD1S
v2JqS6tt2yP2e0r2YGcqMZcwQH8+rcqqKUmsp29EB677ec3dWVVFjxyqiksoHGQx
rJS4WE47YST+zBnhlrt7l5LL2z78APPVByRGE9uzVyCayZDNnENJEsq+E9Yo3goD
6dno46htaCs4Fgq5QzASazVLlc2usdhoDSl+HvFtgizZpnHm6H6fJkhUW7bQyKJW
cG3qljVHUPK7TxG/o93SylQYuyRciSCFNK3g1y+t4uqRabUqYXJLig0nrcrOQD5Z
TEYHmq5oD8EPeBFWBwmIEnHj+iunYmWaRYS/ueHtuSeNHWYm6s1jEZaz7++y3NQs
yQct0DYJp7pFvua5HqdxNNWlQS+lMpERRQcjiUswVsIHhskd197wvNtGDgVz+Tww
w298imXlqvgmEPSGvBZO84hefvRHxwo/uNOcHRJKkFYl/5JCrN/0C1Hb82N60Z8j
zVCFklT5/ptJ8ZJ2H4K4mv2AKE+xpY9XxflcMtEO8l9I5vnaYmjytI22Vge9mMjU
0RjqwsqrTuDSLR1BPuCcPoSCMqUHUmP4kc+VxYqmsvFxPb19Xf4FKAT4R8v+lJKz
KFZc/g5XmwLcJ6pxyzcCFlYxo7UWWwWpZ+DqeBEXH20J6mX89hpKbJ31GQfLWbr5
U6Eq2R86i9A/8c0QJXycrj6W9JXFGfT8jDbMWs45ZR/20x2Y2VxRSqc5X1NSGQ3f
Q4mKYr4/goVzyiKBSqY4RpduwIDyh/X+/mKm8qR1r2Vcoa+xuBXa4/PlQjnf2XU/
3xePk5sCXE7QyQz7QUtlblsvbXGpMLmbqNBYOy851MpkdQDmNxQGnowyDQCLzgCS
WRX6Et1UYQNKXH1W1bopXmBw2bq72b5mAp9Ga8X/BYu/WQMKB1wFM/SegpTwk6Gs
GW3FXM8Bzk9jKX7dWehC+g/LVx0sZT5pawbUD9h0IeKKChNfJUxo+gbE/5VaE9V7
uAV9raOMlEBNSkSbW9zYp36v2onFzYML9q3/ZXb61RJGz0vv+Rk5LcvuAXGlviGO
LBRwloAbESh7S6S/AYKW7BS17v9WhE2cmxDJkQqdqid6Ya7uxLLgqDuVeOkEEI3v
LH9zw+ORbs/SUZBN7QLyT+siuowY5/cgwvga/fI6rrMK4hGyD+nF+/O7+8aDRhMA
5Yx6VJ52sXpXSNJ8SRY+STlaL7f+HUX9dZ99b0OYgKaNiYLsMibVMcy37Rqf0NRv
rvIqoF2FH/VeZwohAO2Cn3JnVffaPLN15lVcK4P2RpvDJfi/Yyo0UY7+5M7o+Y2U
/pinaTWXGUe7zE9UXn95ew5Ra33Cqcn1FWius32AUA29+/3/tLE+hE/MgfyH5Dji
UMSUNMrGPgcYbjqETAkXvLh7VQQLUvcSucTyHH2eqyKTkR6VdAlv2ffiPQOFzbZ5
JboDrrjpJaaoPIgn4SOhJXT+FJuYp+srXNmtB2FH8j6aOlRetWrPNug12d+zFoF+
7a4CowdtLVgTqkqmTbK9Jhza+YP1HDSi67nbYX9BgcLcEduPWyAJwkPCCiBFe9lB
S3d9uelWxUwoh3nMHO4h0gGmPEJPkn3CGhnbH2Jtexy0ADTq3KnWz/bs3GF1zb8c
WXfVyVgG0TonHxWZ+Lxfo1u+D9XWNCsfYVIPYR15uLI1wBgBe6fiq7Q8fD1GsJLb
1v8sbzP08aBDZOIe144Db0m2idQoy4DEaCDG2b0gp7k5Wo5FAsufuN7ZpTNTU3N0
oLSEIrQNMe0joS4U7Nhxwr5I5wBMQHov87hZAjJE6XW5s4/33fFjhKLyyNPUlW20
/CkwMsJEUUbSqb6S48GwXi8svkRZBzigFe3g6jb/Yc4J9z+AJNK0NGG8hbtJljo0
bqEZB4jhl/zlICHq56h8KhYlUn4fnYCXgPcOtkx4u9V60x5xaE8yQQ+GQrEWcK+S
eQHEikQdnIOaYy01RcDqBBnsljkmBn1w1+oe1AHPxfZmv8ne5vMG7szyE6EfHczm
jbFDu25vGJ9vHCqkJ90jN3bp2QQ6fq5L5CLShzpJridlSbDa4jWg4/+9Nem22puw
SBDEOP8ai6CLHjBtSD9zzTodBYphJtyws9AWW3b6kct0X940P1z7CnkPA5GPoMfk
4Xy+WVKSUPmh30umWzY2qcXTYrLMontnxVfCnnqX21N8kqngzt6ZGdtvrrHnEaJ4
mge9Eui9bgFKKvLg4I0tTXmGYNF9JZDWvDEJ2LQVb6J3fxNTOTCMiTrVDG1jRah+
pMq+RbtcvbYoMYFUgwjBl5lNYU9ICzXdzmo8Kjo9fT30lWUZGKpromvU1vaiccui
ozm/Cse4fsjpPanhDY9thnLfnVEaUoveME6/xGlqGFKxclJ3cW4PmoHEMlAjMuZK
xFmD762+sq0dd/AVgq69Y0JAP4I4pMjkPmq+mLLg8hjPLgkY01jYh4TsQG4KooW1
C4SKxK5U8nC0QqchNJIBM1+sBD1EItciI55qEl74kASwMi5FBa8ijR2x9qui3tFS
L6onh6w1PlvomkCxjmZaqloKDE5Q3EmLy/wR8CQF2AYJt7UNhrE77Slos89d3DOn
/Dq4osWvYGDL8Bjc+w6UQraPBq8KwEmCXfkHazeFrBkoK4mTnczBkE4HafxPkiQe
kngt9LEsuhLDuibPn1HB55Pk75xqfqmLeWWacyjaN8FFj0yBxEIiBPBjFGCXhRDB
8NHCchntd0g98OLpDxlREK5G4zUrQDanaeyTRrlvAwXdpdkruXpgWdNj2T767e48
13ysWXhZPCJxheGjnH/FNpH9magCsIhN7A7l0vbSWehLAqmiLY2jCJLg/WAanEx8
W8Jy25niD0tSG1LIhWFlnhyT05LHy1aTgdMma2vyxgXVzpnZVHpfWh4+VAZloqI7
2N9U/1MWfNxGKCDvTJ7nvmpXFe4VVkv7XF208d7MC75FABt78uIYpLM+AVXcKbOj
wsvQDUdF46xFgBcSwBhqRSn6yDNDnM/fUX0TGPyczSqXHXmEQFDpirR8qdZDGpNo
JgYDrPXaZyLh4ueYHnZQ8UElcEtaewSik2MaNCgOQFpr+CwDzklogxkkFaPKRlIT
hPCyqODdTgv6L3VVlEuSePDuL3xtoYI5VhEOH42qNRiaX1Id6QAo//QhOKi1dS8R
dBlxtBoC0B43lj3YR7Pkuvvfdpu64lOM/d9d5/5jmb1tQUldKqtmZNbxz9dfuyjp
ZEzwgIoqG5yfiACDArwtWaNYGaSmW3cvM2H8SE6MyLkGCu13LzIO9E+8BmvBesYN
xGXzT5QpJDHZ4ezQetz+LovUNAWZNwZmA8/Rd8RU55csYSzSWAB+ISHsICMV93yi
3dvkyqpkxgIP2qb6GOndZtXngx8VfiHz9Uc3eWNH3p5AtehxJC2JdL5TM+Nex9gw
lHoKNvKMeyA+c8GZO/h2UMwB1pRJ82bhRCB7p/MM1K5/M124lmyxENeo+H4OqrDS
v5LtKgckkWWScPd/aaayRcnyFldxb0O4bPnDzhOXrDzw0ji/nDqF4os38O46QSWn
1Gmrjrhn6TgRtl3ChLXOGg7n1jw8b4iCchcjacKs6d6/7KSyU6p8NUmupo7JKP28
PJvfgQYIlhd1SXPX/dZwh7nrZvwqDBjNXNZjmzNtvi0bbQUrS+IsHzCqRsmzwYdQ
mdUieHCKz2egHD5n1qHhtSp2JNx2p18yArvXr6tx9MbA1O+TJzmYetKmTFki7oNO
Rw1QivupEMmK+mPyPSc72GsosDq7ns+P6ZauFSL6QTfLgWXyXhjIUJA1zLrUrnt6
SKXQpLwKrNAXFBOAhrwgGXJ2e1g0DYsU5+GgIinTf6fJ+i78RXqJqMaZi3Leojz8
mS8FvL9WPHKYETgSUAInBZYK7DZZ/4DPzJEFS3dPYWcRore1pYjIprQ/K95tF5bH
5nKouf1RiKnmcFBUYMj8RZn7ksxeLnNdCmktxoiOFUWCMi2oygyjcrGn0TeYczAI
14iD4byJSKFcYYvvLIosHvPzAXA1pq+Z124RCEMOtdcdo3f2kcHOUhvu1IBczQAS
gBXYSOfoN5dpJUMZrkSmAxzvnfJo8fFeRVsXLL+1au2QKNQk4h3toF7qCkhaGt7R
woJk3GhRFs0yeqCiODXLeLPq0gRRk+eOE5wGI5/QJjRXcOP1dCscaz0pEe0Nb6Zh
WqNAxvT2ILe0yo7ZsdQhX6z46590cMIpTBw7FeCcqMcy7TuRgKSorbYNl5S/2cl3
G3hdeCdj1fxGlRYp0ucxTdM7T4sKT8PMdPBjl5b6ojS0YQklrHo0VqsShkov/IM3
f2UsAOJWmVbxB/ThN+sytR7sk27z82+oM4atBnqRzWhamUMYKves5hZ78Vpq7/O/
o9QQcGffXEH4HuePfAmyevGy9500Z+SsqSnmN/5elJEP8J2XtaefUi3h3LcYoT0i
1u0nzdBcPTGLRmnBt/wOT2JbQ6sjmoK/XBHHZu+2pmeMjrCZOLeHAg0rGxVrcspa
d0eHR/5p9DXl8g6Ol8DKcyKpzRabwMwfoqTcps7C8ugDo//AEGXmgWYUClAcicDg
xR4oLB2eRzrv2eMKIPxUSVJaZZxMsr+Y96sbjVaRi16nYk4F9ziCN+LTCkPte2DS
yrfBTNItqdbiBTlmVlhQLzM0OSiBtFXBR86okBocMRUzXwr1cbmpQeL3UjEWEaSe
lX+DoVaSkT03CDLzgR9iFauCiBW9v7qHzt6zxV3dQlWNgEQmNKkmgyPOSNEVtVjF
JMOxrrf/28na9RPWnycb2BUiOeKB4OwnRVnsRE5v/enNWjlnnYZvZ5MG71ctfWJ+
tFFpDnSNAMwaG5C1J534QplTu6Gvirkzb4eYNF2ETPoBxdQ6U8i2gU9Kec20tLH1
UieoD2MsqsgOBbkKvw8tJSEuA++wZAFjldp9M0ldvyi2UeHVn1+3c+6Cpmtqb38N
LRNySDAN184fu1lvqw/QBJp6VS2MW46EGPN4NM872n6TfRtd3QG42eASJGlMCkoq
fAP+9y4YpwknoF9vwRrNuu/KSUouLwaWTNivdYXY4tX4GwMfX+rLwkVkp+bfCDuO
kBN5CFvqkrYtzaMqQHdrujHcnQEpi0HJmSUu2L5JHWwoq3+u8YQCM5PxsH5lBca5
H7tDU3tANv16s786cuVZNuojxGA+x6fw0SlsLlpKqyomNcecF+uAbKPG/H4UgX2O
s4DXYIjXvjYHKkVrPRUza8sstbpg260XeQL8ytQ64RCg6WRRddFej06Ssnr+NtqG
te59KqtcDdx1+beHkyfc9y2IK0FakqAqwlkp3GK79HJha6A3zK1yRFgqxt0n0GnT
LUlwCDyoQ9WFVFkOy+LfvdU0+u6rxyTvi6YG8CcpTerkNTRohDbIv3bkVLWDfJya
LmLQSRnREG5IhoZeKjgJRu6NfaBxvEiMrh4lehjpgxobgrk1yHsqo6r6VrLwpfs3
Zl0TCDJUDeJRFKsE/RNEawPi4y4k3o+YI7bmkWt+xLFBJKtlCOd63sjOxQ8MNg92
8zVHVQoKGAyYbkQhdukzHsFrFlzZ9QtclWDTqe+CqgRsJQNli5GMMZGcANtJEWIt
+x4u1fonzGsYXcuHl+sSP2ByV5njJPv2QyYS1+bvQY307oNuDcnh+0e/7gmy6TOw
IRLnqmNxLP97i6O8+W56vxZZdREaaIN9PJedKxXkA2fbLVADcmjbKP+Fs7LZ8LlG
QwbnIrdvLz7jLSxB59LnxNR4mkQircQzKxs2MOgg32z9+K6jFcuqOlYCS/lFjk4u
Ie3EYJmfGNi962fkp9LAXvEcQ6Hq9hGB5TARfwMZYTVQb41NuNpCXqRkEee67wtP
ss5sZCsmw+DyQlLeFGG4bQqcPSZReBM8UhNDsQ0xkLlhuPltYRWMJv6QMfHkrp1X
90KSRl1IdAI6qFG/3vQcIrq1RcWDHmF/Go5mRnCEyetU1g4tVd4q0XnoqnfAzX0N
qVh8tyG18DIY8UvM+jz6cKegXQAv7b/K7XLS3qN48YBUTEhQHOOo6GQh2YjQNa4E
F/lThM4Go+oXZdwbp7+Cv/INE/cGOQOcF30skTHYXOk3larAGLjYESPygrXkd9Nj
6/jSNj/ox/KTmu0Qlee3P9DJVu94125xjQlQDFRkKPpQJJcAuh1d5nilJXz787ti
EMz60F3FzulGtAyZp3TXBsXhjFj/shjTSHBBPP+LRR0ZELOwjyaolxvo2rZWTGMW
r3vRoZ8xlKe5qRev8zeWffZT66R4Qb5Rir3+Nadd3q6T50uq/QGvlBFiXpoP5Tto
QBaz8rYj5W/q5XSJhXSp0bW4dqgwqp3RPN18vFA5nqbi2zO+RvXgY/Nozj7OBDvQ
dVKdE7iF58eHmGeeX2LfjL+bHowtjsmFM54bVCT5hQPiOhuj3+/7/Etb33vY2dWv
5VnuXeR0U8e3WmerzS1juPk/sPlFbljM1GIuinP1KFtZ+Cd6VIqrgo/wgTl6CEtF
QqiUz8ED7vYYNEuYZITU8YXJw6tAl18Ne/2PG64t/Ti0KCTDIArUCh+qnSnHqhtl
td/OcQXtn4ZTXMbBXBvJZTQWVgZ3DnLVBjR+HJCq/3UGhWy5yhQawUSBKUYGFZDw
gPOg2ODoBaHmMPYofXdq4WZ4vLxspPA5ctnYyaM+BniHO0vYosw5AxKv24CST2bC
xwD+GydJlb8yrGErhpwJob1Tr63e8nNXQW4WX84Ha2qiZS7CCmdQ1E71xMV4UXKo
Jp3ZuNt8VDdZAnDHMJk6tCYLmUQog5FzNgKh498wWpu+ha1AHBwMP+2abbi1h9GS
zrX335Uoh9CdqDODPbA6nVaasTsgtYDKn1KHbrpfgfRQ8uMkXe2b3HATu7N/kih0
C/rw9xA3gQODGeDEeXWdOmKgLSQeQfYFlgzY/0mH53JXNTY+PA7Qzzvx+W9o2+iG
XwjazUCMjeQPqls6b+C2C3wQMfACZ5LSCvxpAGo8DyxBU2d2iFKxEB/Cs4VFR7wT
F+Iyc28CHXT74uQL/BzhNrIyQ4LGR1Yukd/JQFO13Bv8X6Zh8+OypuPYp+oazSEM
+routt7+28lI6yF+PXQLnqgDH4OXygcmNAf1vQZjxLh73fGTyhPhI8BPLuWKoB7E
lkkv1wWLYgLEUW7IO6tb7OfMwammNq5UGbAFRiB87jIU5qRfDiLpRIAHKRlSU2+f
KUuadv7QakwReJjK1Km3xk62LURcnbjdWsxNH/eXE5Bk5wpzSY4p0rY8Ms0u9AeM
CbHOyMUKIp2wB3cFNQRGwYycmzd62jxTs5eKWUxTdb7XRLVLdic3SMq++jB/w9CV
t7vbKpZiRvTzeDopaYAy0VLVfbXMRJ2Bp1dMSijGNNHVZ4kPH7l9kjqBJ+FEi8Ve
rfF5V7KHdtiK++sTX2FCb1veb8YAJWwy0WG4o8u+Mc2sf6XnaSY735nc/6s5F4S6
/nq4nzydxkS00BjoVRMV+Bflbthi7jcMKo8gGLr2HipdQ2w15mP09AhPAB9CCK5G
u9EcGlo6rEsb5cnkY+df51IMTfY19bQNeRf7WsboPpMii2DAfiTXGvS2icVlH1T2
ZTjGiz5xwVXY9hQk9qfsBFjDiOIdMBV79xrHOKiFsIgz4lT9Q1+0aQ53InZ87HIm
W0UNRUg2LeApX+N2iJ/jMjSy6UG04GWs1huFif+3cjmDGqzBob3PYSxOQP4gL0Qg
wTM3jSdzYPVUmwWEWCBLiM9gevKrgG5J+w7tDopGmK3lV8DEXCOfoThr/5eXO/+D
D4iIQ/f+0LzvX1wh1egmtp0nRF7sBbfYCl9tnM1pNXomJFj87JW5x+ezBYdlCnMk
Ys0Qw0g8pMaGILKxPn5tCGnta7wQVa4t6RXuVjZvUGz1qpfpHqt/aYx8f9FXYmHH
vc4kFGTJRWacBr19Pancg8Ri1tF3GvKYmsTXh1oaljGqMAbvV8nyyXm5p6un8x3m
J4u9vDm7pwX9fiJGk80mlu0yQMfUkPriMBwpYEnxhpgxMb0sqlBmVIWLT2TbCpAI
tilWgtIfu+XSZtRc88/H2FVaw8BReH2a3tSomV0qfeFeFzutKBtylRUjZ3krYeXE
xTWg5K0XSs0oyyALSr4cwKXqmObO7ufBP9F+6N1eidowZ+W/OPE3qsWmqG4Qe8NT
alQuxCnLlYRtvFtY68xyDrSUyEs5+3l/tENHGKo3unpYW/RmIugIq6c4jSu++HVr
HX4r+BkOaQq1VTZCGoxyu4XP9NIu2dYzQVo22JM4TGBKAmsMzx6zpoYNp3TWnr7q
MK/8aisbVR9M+szwiwLJ2ziowmZMfGcc/1Yk9Chika8HxHA3oTXskO9njnDnaYhL
YC+KJYUwmiRoVWPqaYr1S5dqkIkfwO35gxO4xIpcusCQxDV5zeSfhNion78xkOVf
9izzYMd8ATjxJTf76e6HEo9ukjNhemT47b6PKdVKaPNlOVCTZN+dsEcdOU1ruTvX
dx9zVT41qtxLwt3oLE3I0prum62At9ECYk4Jy659u1huOkDEaP8z8I8AtrkdDbjw
WOCQehE8A/bzh/ehzNy9fveas+NigKMLLAgNEdhElo5IUFWt4ptuD/pD3YKFh8Aa
ylEne3FSVuPYO/TtDeMgsaF1171BzKTq+vfcA9zHgvQL7DDSUI0fLaqqYS0oJQPh
Hhk9W2d8gyGy4PIByduA2RxeRsg9P8gUUcjq6b3JQyumJYMPa1tplaP14bHhwd86
jIVUfBQ+XE5S+ulzj8fYqoVeUKGxE58rb78EgOTY3P6gfnCwxEjHerzBJZ4zEFTj
ZIQDpAS6JcAEIqRk6oRWVmlamVlsct3A0CklTQ8jAGDvt/FRw3Gc6F6jjmwqYmZk
PdDTH3zqBraD8LsXiEh3yuxA6IYMkV0Yg6pHrbrHShqSj4uQw0v0E1NO3qVHEYHV
LOdJh57GscGNxLNBuwgcsU7n/2loiECSIhyLGbvYvN9VRgBNeQsL8foTGmW6XV8Q
KxFsSFFeMDlcSIm+bka1OKr5ryk6M5R1VKpPNRbOd504tl/5xeu2h1E8tZxPm84I
v4vMSnNjx86KFP1oDw8dAs2zQBzuZvGSnMDWhjKLYZPlmZ3OWb4BnQ5S51JNWXNs
9oFuvVK/eNMObSYLPLwRFc0n4eHvzankTGg2cy75XpTS62JVp5i2Ua6Ajyy87v0s
nzoNFPUvy+it/tgW9ll+djcVBl/o0Y/Fj769Amswg0Pl9R2n7bktpnPpB6u0W4nk
f+1vBb5L8vRoXZzy0Ok1qmYG+putl04ZiZpYpepRfi2Btidg5ZlafiGgWgaLxHPW
Jpk8MjgDgw+pw/3v3ypiGi6iILPiE7j41AYofZ36RmMb2DOHglD3UwpZG1lL60+j
LJ3ofGxSr2m03+3cR2xm0LknMSNSnA4PfzJp/AGdELtSAYd8uGxPt3R5mSJxt3Ks
4qL8qAE4wO+7a/jxBf12ibKETpAbKa4C1yS3yrDmyybLx1Mr5YnymgmnDEPmECeo
L3SqM/Fqevjdbd7xzStiT8UDs2xoX4oS9pJ+2wpAcgCf+++RXU3qKGMaI9UPj3tx
EAtxBIouAEnk3y9JnNh606TUSHwThf6rh+AHmc0UM6mC/nG6sh+D1kVSGONd1z3q
nIUDCmSYcyPyPI+lJwwlsKFNGgIVHYiJaiHAm89LDZep9oJpCstEV+9KLwKTUPt7
2IbriGUkqfasxP2yfNlsBk8xTvDvFlmS3OadvLnja9+HKxK30IGPsTmk9k7gLbOr
MvbV+rshzUrjSLMiH3RHGP/BsPtpVRQepAyDlbQfu3QVgbtwcOZDhk6vY30lMRuU
wazSn63HaTpzvCtN3lMHcEJgfGhm0onPYDyEO/EmJwT6n4iYgtWc3jBJ8qLS0IKP
ORHWIzNvMVtVT9FDONvwJVfToYqljjENBlkQ7J8FvUuB1f1t5iYBJw6lZ5ZINP0x
y4jISbjlethBJGlNoWcLI3goweO4KW/5H9wEufyxBOkE/mArYVX74zmWdsBFiH4L
1qpvQdCL/u+Ch7BmdLMiee05CA0/5Kesl55IwqBPQEHYEuV7BR2Oi/4+sZFPNyoq
4ygYTOw2CJ3azThMHD0MD0FGKPWsKH4pNu79o4P/XsCyFGPos4jXNWGnO+EaH1bo
S1bPPQ+IZNZzO6GfWI/wqtrp8bZqDSYiLO/HdCBQBU/oSP1O2ikJy/IE5ZMP3Wv9
cxP55dp0BpYMwGObmkXjw1aFScM+RTFYGOcSempxMvx7rYlCMfJeVcVW5UjPh5uA
UJMAfCFonGuy+8sAREzWGGWgFjmlP70frM5PMNeKkjcrF6S+JP/+9kc4ElVzGgAG
B8AUWK1LdOUHKjQAqzY5L6IRY8k1tROaMHSqHXGc71VX3mBoat/oCl4KJUFMFUNt
sKM7ihV3qmKS2t6LZOTlyJMCNj+Qwahm862E8ci72W6oVD55ET1Oi9jxMj3cFg9o
G4S1UTTCLIx/WlYs/DfwZ2ByLmIlq1f4dusZGHAemsoDl5LuV/FejaU7Ga04M44+
XChBTXyRflAMF12h3N8ghnxmNizGg1LPrkCCSY4h0YOpA3NbwemU6iN/bB+xCZON
jXiuN+KJ6knNjGAGg2yY/ZLTHF9Lrr4NYzK0IXVLIOUc2G+RVB1x+nUbkgByYXi6
886jKuqfhZNMniQcnDr34OF21YNsBTAbiAj6/3Qr1MQZtdrCW09pJX+UF+Xun5aZ
4onC6NJ9+o7QCDLC71ylPirVW2kHjM1bdYOb9v2kfcUAvGaLp3TVcnSIjiTcm07a
+m4QeSkqbOb3Cr9MYeH7bUqjkpGxzbxQfy1q3heVFbpJ5r9gS1xbWaE6+FOz9DGX
7gezW3sghXTtGJinEhS1t6o8qO74oQzlLdFaJUKvKquWcXW8ZOBXCa92rUyVaGVC
X6dRKLvMsicYA4g6wv/cfIuyUIo0dXtu1ITjw+HsHdO+xmBH78u+mcJMQV3yWYpu
rVu8foCwHDc1Ts/2DhcwuB4k/jsobZsF4kIZ9Blha08yFas4SsapO7XQGBd93h9v
IxyR4Som6yR+GpBvjKs1VgcBerW6F7CPw6+lS1AWzWg/vmZ3wI66pyos/ySQrqRB
gX5TbupVHkY+xM2xxkxYSCadvE9fLZS4PhBxPYwJ3G4TUV4gB9BnhT72f1hiwdcI
NjQkRV/WUxhlrz1Wga/zQmq2LF8NDEYaeVYFe6f3pPIhTJrpNsfiAFpGiCN7AQU3
Qlgn4tDL1yVWB+JbHLupClJAkX13x57nZgcOMhK0ITk/4Yy+mDduVVJXk+CN1Kii
X4B6GAofHQa2VeDqHd1ZBHAfj6Qe54TdW9isIERX2sYTwBEMG/cb+XRQwd5dXOQN
+ZqigY7df2I0r/1xOJ61GeZrEvvvu8YU2rJSxgtKLQyiPRW0UK9m4D+qhR9vi2ip
6CDSsqosylK2BU7ESyN3DqpHSegxLgUDztGLkxw1pR3xQGizugGB6QaNA6EYyQuM
SJLrVrtUGh7h+6sXKbZLqoSMtW+IsmUHg4y2T7T/JpgOOfcS6TFusjHosNrlLUqH
14yB5ZMeIJXeg73sbGXBub3OCdFWggF9Jp2CYLWFKoroFLWZGypCHYtaSti6/CIl
QKhkYvxfFXwCNT8N7Z4avLYXgg74e5JB1X4VoS3QSHHZ3fJFOcIZVZXiEyNUEHif
2/pcoKKNC2yQkUFFyzZydF9hSmJeMLdP58swq9BnJe0krbR6mVLq3t0g5xmwPwMo
ldQ/uGHt9bhBWdqwAMHQSqt0CduTeSUbrHWPDap0PlM/GE0BOyy9ZY+/tRImR/PT
2WQ8xzluHdsUNG4RxipITPn1MzmjpA/5YeHk1f5ra+rv72EbEKd4EK3Zu57Rzz7Q
eNPLX/AtRRYhy8czhvI1Av1oSIHTeZPr6i5hkpFdZGTz6Qp41h0iTi+mQQuyMpZY
uJ/TNJMziVZd/PS5UXfX9GdXuvbcToxcdbU+jIhHj31cWib+BLz3V1+MpIsQ+7TA
xMoe7kYrFaHZxBH+2Ofw+Kx/nQA+qAqOlHP5855Q5/X6MwkWT14mnj2XaeXaESEQ
qGfH5czqy6jvHedFWntWS295WlgOSfYliRZZO95bKvVbZLuuI8QecjEJDCtkeiGh
OfT1iwa0bk4CsanQVUZb/A3TWFyEzfmpLD0hdfbE+Tiz809GgL5dxr80MQ7aIXSi
VXjuLRAMNpdSUw6ZPzFr+9+yTs0eip2LfLFCqCSP1cf85r71asMpJ+XzJvUfz/N5
fjU3eaRP3c+1mfEK5cUfwto9E+0f7iqOavBtIwqI+F4iZFQIczwH8S/6DlTKD4gK
WQguE4xVJLQld/lW7gER9ciWbqESf3S6KF7OZanm+Q6sjE76AchQgk3G76zc+846
9ddS95VVowrqFejh6Q40fuOi1bCyPV3GsL5AwzHsICTiFq1ICk+GBpvjiP9uf08m
+9g7Tbn6oB6oOvbbEgasKyiVzX+LwDjczygSPLvuhcuhuoPSR5WtA53qUguzRqnd
Of2dESEYsS99dxOX0sn+LPuNIqytVwlqZcir8ynLs/6R/5QCgM/66x2cibwKRFWO
Z67iOFEfJpKmTbzTjpSXsaHbBkuhibL3EKrEZ6Aa4vn00XMPiRDvqNL2H0PDvRuS
BmAKz99PoNvFwXFbp9vjUHJVuIyAJMsUYyvmaRmfsfbO0xFwwG5PZ1iWlZ7DaOeV
1AD9A3Xrmwn2dz+GkWw74/P2NHtMUdPRN53z8ItWNOoA+fCs2irXEqJlSdIN7GHF
wb8suQ4HRRDO6yYBUgDjWcDyIr7KDsCRXf4hA0NyojyFhxjG6Zr7bf8VY7nC05kg
e9Otunx28XMImcb5o5bH1w7jzB6PgXiPT4g0tAyLl98KWlwAkroTEqM+5yTH+ndk
VHwqvGkcHWRtcwh6clXclByUT/RATMcg5xtXLHD0VbSBm9jRPTYwfCBV+V1YxmLs
9SGY24J712p4K5nuHtUHIdnP37T0QJnRBhLz7sgvgx+/3QEy8mWNvI8tfq4iG3Rm
TlpHh6DnfLGiBxbGwySOYXsep8OrsIS+GFul+KgBxkk4J1xiA8aNnmxCGk05oDDj
QfISXhgK9MOfsGzNI9M6Awd9cD5eG8IQySDVE9H2g7HXvctJxxc8nmAIP4mDMeeY
WGiZ7ZH/srAOgIEKqlfN4c/W/AvAQ7TVjqGMfJq6CNdVh6Yj5VvlcR3+R1JXYIXt
hLKlv+gTYKzNn/KBYXMwnS/LaN1PgRSjeduiCFQn1hP6sU0SPpUt4Z7uoLoNKgth
kkFoi7IgPKscUyl9vi58boNWZzy7tWaIw7JxlIj+UGqt4gK6SDqNgeOi3AkC5r8i
GRAlsgbyb74xTZBPh8G6xbXaLckzuIqhVqiqKXN0yORsdvkNcA8UHWMisC5xEWGj
++QHT15oj9po3XlMsos7/Tl0a4wMZNuyb3e2uVKsUPnAPTTrFV9+DgzDhJg4fUIL
6DgkdzWvZjOafCn+eYPktn7V6elYLwXdqbeShQEsJMorYcDMCDIC8/pAAEnYhVuq
+JjMF8VM3SnlH2fqjzLoelZmPe22Hk5jRW6bZSOAEt+/RDZBKR3DBpbUa6t+XwPs
sA1oNhPpMJqbSgutVMd0nq8+LjotyVmUaFEnOrhtj4DfxUZ4AaBY/T84fNGBCkYy
yh05IuObnm+8hpLDPPaHtiybiqee5MB+a+uEoF/NRccZO3nQB/45Xjb5jedQnwEc
3PwuYGcLuQNqbkUTT3CVGR7xS7KGCHtUj1Zfuh7mteLEjOtuRP+l8Y/fAYTnViZr
2DVeG6edF4a94BdprPP/HBCcJ12aQD4gGp/wKR87mVXYrRPH4ILYNs4VYpyN5WMY
rdXmu3S2EE27ktcToXrgzTDXYI/HPdQH+35kgAUmC+nhVoecLMuj8QUWkDh+qxFJ
0Q0zNUSE/5ahbnO4zlyjEdE7k6583AhGY9PNPvAE3EuZ/3FnNcMT6y5sdK1jvmMS
yniaqjpK164ppkP3jaYJbgdGEv6E59VtDI1sIVLZYGnbgeZ77l652LiVx9areNjK
ZtyEFKatk+o4OD5PfKpBiFmDaaLDrh8KPMM5jR5TtWXtAFBT+dlXSIbqoAk6JXm/
NaOHOgsfTdf9P/KgEePSEuSMk71pJMSvSpa69li3i6IgKCoF47+s3tA4LbPYPvzf
Ai6knLVuApFNAWkHBRA59ExhdHJl+oQ5qgcokaQh3GiJk21CpxRUu8SG9LY0I+5n
5gAd3J9rRHMifPFcyw8ncXZjqDAW26Y/qDB2kT6WL4qOXc3RQFZHgJl7sGrYBNVq
rcXUFFaVUPMaOMwfQqg3ryyFowgN1J3FnXUC+uFRNqCYq7KECAa38wid73dw/js9
QtRiQ6VRGaoaJ5n0hQfvml1OM045qzKpjS5ZrEnEcV15o8gr+a4Fd8+dnH11HfqZ
5zbRCcNMCTsK7JdTjP01ZfVOGEMVylaBCUq/PSk25OUA6rHhdtS8dfj0NR3GBTGi
rcEB25mf7t35ANf90mGt5xZ08WwNxmMSXkjiTeJibR4lHT1SUcs7hdsCEYNo+BkV
YCaJMRAqPYgEFRyckIY8tUQkPGrukSSoB7dxymmxi9zwInwga+Hsyckw544QXUlB
6ID2lQvH7woGOlc5UO57S1BFu66+GneOkZcTaMYzY1CACvewK+IRJAnkCCHlTM6H
DGm2nTmJDo7+EYwlvCURaLv7WPQvnkegrPuozvH/seQ75a3Jwo++UgF0Q4O1BfAF
H9NmG9kGyefd/zWIUBF+e7E/3Amwe2G0XBPVzCbMsLEHp4Tdsi+eQGB/ISejjB37
Xf/dGd9/0TTVGqyoWzJ4kMIZMsGEhe7xHwCx7iyGCVtmNx3XR9mY/S5KZ1OHvesc
RbhvlFwYxUzKjI6SYV1uTLCZOV9OsCCjzD4lAEXVuwjZRGdd9J5aVGciC3+iCCqm
QWEcrXjtDzZC2CSifOISpAY+Z3Jh62lTdEvDjh7c3PyLl3QAyD4OPiT9O08GpxNL
Mv0YRQRn1CRKm3s5H3IOQTklu7+5igPL6VKUHSkCXKWqR01PS5UNN8+SrglGt+Ho
hDR1IHwKDEEWL+eo28ou4T1rI+luRI+XpmonjbXBmOVfml3BGhM2eOOf8P8U8AmA
ozB63YW3cE+mvDj5X3qVUTcJwGAkEEexxZougUWuzam6oIo9zfVUX0vuvi41A0Ve
VK8ydoLFPRm4zGSZtOPIGY4MYJEHbHav/WS7fPGXS8507QzpdgIvngkA/oZNxTKb
57CGzlKqYz4+vIjCFofA15HThvTv1FccDSlXhNqhxxJ8QbWv6qBZyiK0aSTaGK7I
+IehH+iS6YdkueU9pBa7FML9pfJUEFvDQsWMUC4FRiQ7g8h/XO7whWiu2r1vjli/
BsjAgYLYrrRTyHoETsVyCF83Ckrzuk00icAdmOwDu0iqW17i7Gp/0bzLDVxR3Adw
IIN80QwI0v4OSzAJ5bj66ZyYJXH5vRSWVkw0pQhhzud76xIgh6SKIEzm2Wx+aUFe
95dJPYPz6Os/yJjtgNpFna5oNT61QDdRO8qdJJz8V2ycWJbY2lFjPh5ikPWIrc+G
QiwNnjiiEHmvALbgN53gXQ95Kl62UvuHIiQujEW8jZNd+PZ6SQoYBNGNPAcNmHP6
56YiKVoVAM2V+0xlIARV/AmxSZUtwvAv31X5f0b1TPeln0ZGEc5kRPaxF4uu2Kg8
iGZf3AdlNSpdJ3XEHRbeKAgSCPBkkO8EU7k5oEtnPfUQGiRLhczfJq48ARBcn4l1
n6t13jRS+COMr3XeHEGI0wuESOgF0JuHtxcWwQZ1p3N2mSWvuupESbpYFDOjvggu
pyb3j2elphZh/zsICzcNndiwfX3CJD+LBQ8QD3H6+68Q9HSNxxJQUlqlOFRqq+mO
M5TfweQgGBZhy0JXHkLIfj5pt6pktOhaTc+6o8fCz4hgX0pVb2tJnlmKrI5sNH53
oerwYmxt1kG5O412VJ+/uh/IKr2+4JIHwf1dQHZJvqdBaUekdbBS7Y5VraA4tuyn
vC73wmpAbgHwJu63yNq3Fxc66Oyl9ZKzcNkAKMEp/bHTEAA2MpvBfVqMIu/6FwrI
88/0KtsmZysu7RvC+pVGu3hl+qdw0q4KraH4ud3Rdx38LWS+8SEakCLYBYLhDO+q
V4pgEfW4iGfmV41HLxTNofgFqObxB1N4zBQP0jmXIgWqZCMguKzQx9YPtYuKjfRs
9xYAKdGHbpJosBrTmZqwaWcxLR5GVOIPJJFgoy2sUXF6rKlb6OUts2p1trF8CZOS
MOc+J4c0VDKzSrRmqAO0f9rRQGfGjCPF/7nphrv6WfKiuSziJGbeEVJADWBqy1fN
cl66QmhhyFYRmRosHKzdLEJLTfK0O48GkzPfyYr7VgF9MdwrTtPBafRBOCUmInjm
+rQ0hWeBM9vSXsoQGJaB2mvrhxkQ52L5ucIZgDDM7rOtrQMTr4sumyT8GExSIGk6
mLNfVIR557sQgnv3rTxnScQL/TdCkuqPV03uxD4NyuHEyDHuVj211sImT16ft2fI
KJE2aDlyt+2rGmegitHHHIvIXmYr4H0VpEQGIlJyusPK7Yzo3kgKD7mz26A0kp1P
oEylaKm1x8EyGEx1X9PEobhX1E21jF2YBLU+M3AK27HjhtJ9p8KaXxH9J+qryJ8y
vSa0fnDOpGc6UkWR3xTlxQmBhsnDFM9RZCiKu4AOGeAjfDv7bz3wAE9n0Higtav0
Spi7xXNqI522i16om579AyBVK5LJvyGh7pAtb2OLhXUqBbAM7S/TcohPBHolnkm4
uwzA6L6D1+42BKMtbj+VuKPQAFfSpgLWonpGVev3cvrTmAoymoLesiFiRBDWFEm5
PpayVzopL/iaXNTe0Z3XwriI8egWF6Z9a126FkQNhnXLl35m7g8gyK60uudclWbl
neltcx9V5Kch9sAdx2ht/Gi+XsijgItOUsOIgMAPX9nPnIx/cYid9IBwZSe/vmnl
lU2t32V9mF+dfDHNr1O669+4RgvC6TneMbb58BZXsR90v3g+iy6Frw3CACT+Bd2I
ZGwiJgLmQCH9t3kS7ycvmLd4Smy1ZHQ1fFJwvT+I27x3Pd1P56n1ALLi4K0auw/m
rId4ACm++PX5MRVZEUwjO7gRGEZ0jF/S7c14t6A2VafD8MXIGX5wrk9M3SI4F/Xt
DssvE8G8sJWBdFaPmqdx3EIbN4pw/j0RQ4ZaqLsxO/ZBUFveUApfN2vG8G3LvYY7
BiYXrEH1bPTL4pEScqFu6pKTUwaUHgpg2os0YximZimxLJKuHVne6w5d1Qi89YEK
dWm5K3rUI7ZnmfZU6YQ3rrujtpESyGIgb6PVCeJwkGtKpyMng9koODqbdSn8YCR+
+nyWU1bpPidlZeW/VzalwxBoSpNXeijJlpUZ6npyFGY3oUMoO7GwtiYhcn7U/JLW
WacJ2H1sKXqEjLbeiogaJJD8IxKfhh3wgHRY7akHVBGnNQTkxjgNs+LBHAiGOgxd
ZZ54tdo4ebd5xjdOnePN4Ti3RA6kDvRXFt3KlhxV7p1oFiYyuKJCUOjEyHayaEeI
F22XHJvhGPcmb3VGLPek0rdVB6bAjl49jy0rKhEs9KfSSen9LfUzBhl09VUM2ka7
OpC1qKe3oCwhyWh0z2wXupkUMOfCd2+DRyxeF29kRhzUj1TbpF2VkvMqkdsnMTwY
hMmc94xI1SjwZ7skB6ktmnkP8av7ikGLZ6Aau0LEYT5Jl4o08V11iOofD+fS3e5Z
Ffnu4mgaSJXhzVbkQRxiq0Ri21dlyYzR9pDgSINsWwg+JqywKp90K6LsM88AFs3N
B2SuI3nPMlbHN7+BSCN6tsVoT5vEEqOPBZhCTdk4eG94LDlglA53W4tGS2LcPX63
LMIOr7mwKV+6a5F5K2TtnSgvHD8VhIu2laPepTYKe6xtdD8DgS5umrwPd9xBgdc6
Kl75j5WVCcQKwW0qPvAR0C2tIE8IIGrpb8g37O81ih3VU8nv7OKFIOvwGBfeaBba
0eTfIm1kwpv/ShlX8kw1G3YqgjQrATV12II6JDK99NhJgTrvrJvZXPa37bYZXSfc
ivn3EO/Yqghamu6/2JVL1x7r9QXpnV6YuBKzIFO8aFrI+s6KnC+mafqqTs+q+pqy
uSyWJFFu/OF5tTrAOT61GgOqc7uuwcZtc2KrgK9oKSN0KAoJmtE8Mq+CkBpileK5
AYKjX3q4o8+lU3Qpdya1+pyQx8hEHq6sanMRhkLs1NDT9PI3WFw2qqIhinEhFNeu
6i0fLpN8nA8DatRmdgKKWyAmM2MGrWEtfLAdSjP7AJzZsaX/hlCLaHUj5zN8aiYK
3dY0R8zijXkqf2xUmL8aBrm8bV3TNWfrshlmAXIgx1fSiIpZxFJLUeqkFNSS58WR
40Oz0NIswPFX/NzzD9y8/q2r18/3c4r09mQvsKTmxB4FCYGEKKoA2eAzz+r5748H
wH6AI+HKRzhCRNIgGt0SYM5aUEdJ5UpVdr5TA1WsuSDzw+/sDo5luon2isN7Gmve
uGOwj5ZxZKOFEcn4tunxPeCd7GBHZLjgetiSTvl3ARq8c70lttVJRHVmlj+5Gtva
ENqPEotLlA93dzNQkBCymwNjpwcvlbdO5iwV4VE+XetV+pBzPOxmTJi36seoMgHp
WCOIy5xMa8zMJAQPdtUy7Wr1BEKTLCoiv65gCUjD2uOJKb10bZWfHYWyzzn3R6r+
tvrVHBT/2qukLFYu3sL73ihA2RfjLwcPkvNPCt2xemu0FtC1md3XA0Eh37EvLTjL
J0gEcb8e0pQCiGRJWITRbWhQq3AvBrrF40+bRBWnh07ehW1JP8STSyKcN3wiB5ve
ZRqv/tayUK3wUWm+tXNOguN86PAkVJIuvI5bsYPhshATr41X79l61lv8lBN/Fx8A
LOyzTmIfmcE5Or9CCnbiIkAOTwJn/vRG/oIomcPPg+q7/7pXJlPIUyg7OMiaImKp
5H7mA+ifI3GxFIPELp2yvEX+zBYp1ShGrIki/mJ8u2hQP3NiwrNJngzu6apHJUuM
8Bi5/SFwA5kMygdsprz6832053PNw6lkv3+jpPzCOKIGuWbm4xTOzlb4FE/hCAQO
b6Ibl5j8WcrourLsvh8BP76nvOEMOX2q9xDJe07+54U/w/tD9LEqOsh4Ty4HPI7W
J6CJc4XU0si5S55BsMA3eQEn2a0ikK3QvQCfc26Z5BCs7YuiipKXC1NBbT4Un8WF
P3t/b75m2av3eXxDEkBayFrCU9fiTo24OtRLmBFgyCycgFM4Wu8ubZ373zTtUUY5
CBYfzfNPl3sbmV/TAfBLxLB/bIfC1fl6P+abDxvQe5rNjpsARICmsKafm6XCw97F
vJDSpAlDpVCTfiIaplHRbEK6QqGD47l8boTNyfJVtjwe2adK69bej3WBwzuihOPO
v26H38G3Pu2zo4JoawefhJVcDvULHaMvSQlBX3hFK9cWYvSg2cC/zUzYoOjpVQVm
/hPoyiNb7GNBXSkcfTQRpbWwYutHLUTBaF445OBesV/MXJHTL1TEg60sn7Jw9z/4
GWayX5Bw7m4TYKfwVvL+A1GZhqicNBOmJxLp+CQcBP2JC0AVXm7FROS/TX/mld7+
Xs/doMMBfkcSDp9am/e39oa5NZ5Q+BoDxKxkJKYUxMehFvZF7aIukpX21qXhPcN2
abHcrqx+QdJ3jxxmloP487v4KECrK64ZfvRycqFicv4qOtUMkvmrfNa2ntc7lQt8
JCkoL86lUgu2uXbCdytA5EJoDV2vltwLt4qt2d1OWfKVCtjKUXnLJ+lk5KMCLh4y
izSPmafl+8HGbpNucEiXYFLG9BuN5vZ15/Fpp4d/lLj/yOUQmOuai7zTf0QUD6hq
sOpJnXfN3XzLku77mQHJGLeIfJ1ac+7fX+yKFWaI7tgS6qv8X0Nd29NE1ONvxFBu
sd18tjJSpvZ69COoWEXnvaghUakvqoWN8A7jwJ16Whm1KdRaSQJVbA8a34l0gyzn
WM1rnHbgZsrjWcUZCMWeroMEplEEFREAosAxDBldc+F4Uu8+/Q740VBj8F2Nvo77
IpM1nZwoz6SpX40q1O5qyoHWYk+c/+XLPqIscGSIpRG8Iu9Z+gw3JJLY+B4HRNx1
Cr2N2nBDUm++ghBmf22guZGdmbVBB0kSAzafDF7keF5IUVpKr1iK3sv2SWnvmBuC
2UM0n4gZeCSq1OO637CNQD6m3EHftJIC66m52txGSQ5fx37mghoSnT2QAZiAh4QD
18bLH7FhC2l+pyMoMNUj8k2vymQUjKhr6FjPEhohK8dhUcUmDEKErRD/5WY+dX+g
niqXtzK36CiUItQZLVjwCvOori6RchIerHvmLYZKA122BmLRgcogX1Cmg30D1bfV
2/812mnhDXlL/SbM+LUW/vP6vPJJaCzqzmhoofQRjI/qgY/g00/EeAOscD2mbQ1B
I4yh+EmoWx3yyuXzWI/5dRxQLkRYKitQjpYRI1KXtvIH6jbp1lCAts8tZYqGCag4
eXT/u8Z7oY4IrYw0HNXUoMQioeanO5N7OuAsp8tsn9+pVyeY76CNxoF/ixfTnYsu
qCVBmSXb4Ml8XLz/Y2rCrpYBwTUTyDibsL/xKcmbpGScnbn/hdJDUIaEuyowkwhn
0xYiUR79j2PLL6ZbnBRbF70z+YazueQQCrJJusnURhI4+wA68xpHqnb7aqCy8O+K
uwx0dabcnEGeqrw0BN3d8mkpPAthfmsvG6h4f/WcJG6QZQxC7elkiuNbyVz7Jhaa
EYUBt4QK1d13kIMEcsJOmXcdDpiW1o6OnH47okgbHL9173C4E0eNQuo7tQrfIxeC
+B5w2lMS5iWwXtyuSv54OVgAIUv2naeTwBLYUSc9l+FefXWG7PPkDWL1PIIGtD3q
wevnIdPO1lTbzh7awze77iLeRFgvwBiZB+1bVo51QMyOec5+KxmKHVAZUc+C71tl
MU2fqL7AqTnxXWNdHorhvt1I3cgRwgEWk28T+cNOL3i8dlVhcawQO7WXG3GJn1ZM
y82ja3eH33O4BQjTS4tcfEp3SyQdMWJyKoh8t/8ryNHQrnUDaPMeNXFIe9QhoTVB
mVwPHGHgkS1kbbt91UInGgEUSiy2uzCh8b3evQHPSRowaBY0MZrpaZVxoOWYAHO/
efhQfL1xUvKhPsOLMzZFMMDsNSuZ2erYvygfc2jTBIMnUbaxTjcv9oY2tTlDNmEr
sUiDrW9woqvsMeJH/TzjUKK7ilM8vbrXZtCE3wAPPzW2yNTZ72SdhT+Xd8jbCzWc
vxWKhM2GymfRAwFqpgH8d9U4/paPLBuRV5+ZymLgLKN0envD7gi7hLz+bREmURmk
bEEO7cWLVaeFNxQEqiZ2mcphkA+GglBhe0hnsmLVhcr506bon6rB5qBNqTJmgo3j
lGDxfaxDHk9btH9TAbkwFjFwSeZBIL3qDbxhxgaK2jIYbnyDq4qS/aIJ0TU36Rvy
Gr3sAtCqYGo68xhoHqik1sKkCsYsjAEzk1zNcE1vNRb3WhQy12ECNc17GTL+vF2s
Ml78jQxMGsodVsnWo1GUZCtQ2cCwIQ808Nt9ESkkt1jGP7ravoL+pWLvSxP2WDhw
U098OhljY5h+ZcpXjB5ouoXcC4ccYi4Re1R/QAtlcNpUSDF8gN9DtRQG3K4oSiOc
JNYKkRecvUAYmIv82+jwu27Q4mIUvW/5olSpEsfd0MJJrLJnnFKM+7DnUcsG3OEc
jYf8JRUBtQ4bjwds3ky7WV7B0vQyX1KrQZR5JB8rBT8pp1dk8HcGKDZlqfZxE03+
t7h7Ao5E1q8m5rljyVj42nXMmdx/AY+0zgYC9xzIHkZk0wshER6r6rEJZuBlapJ4
vJc2Ad5xPCUBO6B+EfssZ2x4g3+Y2f3atPrCeXXRjeF0CO44oaBrhXVwIxg/Am4e
BR651DdRMcJuf/NvQqj4asL09kd7xg9SR+ssFk1XUVqOX1cJ+UdBcxETkYw0EGn1
vIg3SeUDk3mCQPydu2g+KYtCSuzFJ2oXXTZTvHzCz33/E63ABG61iTgQbzz7TICA
kZEAMRhmxjfMSaczAY1UIvXSfpVOHEJUx8ffVg0UcaF3ZGVcz8Dp9vzozqQzmKnQ
FwaNHytNIUfeW4YTdUM4aAaPwaxbHkPaXELgNg8cdeyQmPi6QijSAT+NKLw/q9ir
8QBkUIdUFv2a4J9qsAssURGHHOMIPjIiLsLDvpHBXM3D7AWzVsQ3PPwcYB8zVywg
Mqtw0Mk67GMTuanDudqmlVeDS1Z8MTUA/ZcDdmTvavfC+L/PNFhINkLc5Jm2U9cf
J1RTbmkpc00O9HrhLmwKueeJYw6lPDE8mqHgYFQbr8pTdopqIMa5kHEEXWIN17OD
rzEDVJFbC561Oc3GWQ5KOkxRYZZkE58QS8M5sVWP7P8lJcOdH5kZoiFzhDw5Xpc/
eGFOvrvX/f97YCh0AkLvq+6uFwyPcdXM4WuLTiWo5fD9ES2HN2tTe6mYjDlf/wCS
nZ1oOHlFercfJ1S4pFZ3AJ8jTRz4oiQP5QEVrPggHb5IycJjQwdJmE/tq5mxLx7Z
omIflHibzgf7Asysu4pAVqIiRJLERorYLTlngTAOilN9s3pP6rWq6tOymFpfWShI
YW2n+xRfvxSTL2wi7qUGFZS5zXkZyDF9l0KbQSOvt6zvguUHEM6NYP6eZV6q48a9
6xpOOIcFANZ+qGLbLZXWgNvwlxuOQmwbPbvE9lKRNfMChRTgGkRS+5Uq0yyJC0aT
i6oAUltVMbrImcJc2hmKgSiYWqGUnFPTSpb1bJEDghrPacShvJ9GhcUNLiS/6Fb9
ByJWUPNZg/GLl0w/iOCLwM27asQAYULGgUDyYcnrORl/qBmGcQRS8hEJNh5r84AO
TTO8/cq3t24K7CHIpjM/QWWjK96jc7KcoXu7+JLe5KByKrU4i17wCv1otzMuTja9
8I1NRv6MzlRtDPCGheaupyqTI5CvNBwdBsiJXUwp3GyVspP0BjzrKx/NZmsW+9Gk
oHk3jdiq/3fJZ6/cYt2hhB6SOJTL9SLBhV4HvQOUvoh6S+IXMPm3/9a7cicXzEm0
FnzUu7K81sl9nAUaRd1FcMzp7IZCEl1MneuUX0IpLDGlLOTO4Yg0N7keToS7N3JW
4lQr72TgV7cNtVPKFme0IOVJlS9fgQ3USsmKtIVlZmh2WDuCuBe9Rsvv1hHex2Lf
C78YzdzlzGJdcd8zdfBZMBbm4UQ/1/5iXZEOtiCxOiyaElfOdEneUy3PioxoVX0C
Um37Ly1sY/KDYywaV2IEYe7V13DiLhqBno+BbR7xpmBZr83EMHFjv6IXs9JCRVu8
bDsLzdRgRRAt0D9AV5SxxS5GCnJ+Ary3q18jfyWrHCDQjhcHNIod1W7nwHie6Hhl
6jb7SysyO1EHAUj78WHEomJVPZE+I/f6l9h+JOe1fDKJu7eq9Lu4MUGtc4CjX9gT
YXm5CUxPQ1kQJDMyx0z4XGzr+4tPQS/CQMjovrOBEKZI2SXx68Kfncv+MaIMkVfc
PjRbAM2v1b5eXdGN/5sxu5xQ5fimbBA6qkqRfj65r8uVrp71dIlBiou+IF73u+xE
77k9cFVy5/K3gD3+y9f46xI5sx0D5fSC5NFNIMsODGPTozooVhr7rMcYik4hxBGv
7+So+EPfkWU2SmEj+sDc3XzUzLKkvhEb1Fh8a/udnD85QQ0tyZci1Fi9Zqc+2r96
USsR2W6J2qKep6CTXX671DY78TBMlLlp5stjKvmHpYRIy8yxITF8xDGTHp/oClzJ
+eOyCM/uhwsOMVFyKygqt8DvxoDKUTo3BqOH9vZ4FuPBMHD4ydpOogPT63Lbn2Nf
g2anvVmKaotHJDYrTpEACfDZOAp3TDq/umIwtSOXYxnxYjaXxjHtiztU0744PECy
g3o0CCNOhAsIaSsK8IZ+LyBZFpWgUQ5O1LaZYiZgxL/Z6SKz3otO/6t/hnhU+PDr
xW7Cs4NPjxRNeT9DLZ1MmoqVfk2zDGkRGSFedfam43YG4fmBF2jJz0J8swlaeLGn
LEcdHsh6IoPGsA+IuJaJARKWYUQRkgEh9ZwYfobBPENY3i7DWHvr097uujDnZWFW
ejYiYW8lriv2xwMmY+AbRlfRf9CA21jS4RUZD2p5umTTiA2m1JMSoesYhkZdIdh3
VX4E6kYHsDY9qqqWK2A1qsnSRkNE/8714cgEmhng5RB5mNCqC2WXanKEjco8kFAA
BXYQr6xJLaCcFu0EinjG0kiSVz2cWvXbYQp6WNlhkK8JwkyJBKzI68d3WS0D6qS3
50jludgO4n30Gc4kaxH2XcSNPiX9zsDKP1hmuDzIdWQkhG/1HuIWYKLmFsRDMSch
zdMr2HfnYtp+ep23+M0eDpnnWnqii8142/Cu2U1PNypwA/pFi90Q8fiN8uhpWy+5
I2wmNoEDE3f4PCkuA1LL8ggW5UMYqpPDgUSqNHJB4fBfOsyLtrHKdg6GagEjp55T
H8g/fERpXKtpsVCTW/SOSnFAM52SUWAXam4N6MTM9q/sSmKDeimfJLAPsFLNyREw
JsnDuQQfFC9lMoqBQ3ZgMnv0zU+8UqLqDu3FIbaFwjA+RPILcI68qt+xyI++GFwm
bH0ljHgjtZEsVlHBdYSvL7sHZ4xObSCL9Jvt6lghB8UvEOQX01r+fCQxcJPuo3d8
pW7SUz+s7lDsW87EVH+Xlf3xzgpoFttJGqEvVPlWS5CBRldMXev2AFqEk+p8oZfS
oe2FeXsmRKISRBa5HEuI2EpAZb12Va55noLQ2tbXjt21p5t4kueDxqgW/LVKQPSx
1J2kOpySzkccHx+jIb13jnEIAi2qGQpWxRjoUyeccY17PDvIK6qnDBv798XbDaIA
2WA6PU/qwhffvnZXkrwlhJ1CIAhK7pDaFco/s7StPXwoWfpUQ6m00+iQmrSrMbpn
vLGIbm89sW9kjrUbejCqDCp8b1bquML1ezrhSMI+bog40BQ58y111KEKaDy17yuh
VvmLEucnx9G/WW5z8EdorG1WOoZilZMlfZDOCMPIPq35ImYF+xIxMk8XSXAvbjeA
+qKz0YwcHcuoLUJm8bNeAEGBB8GLmcHOr/Iw76SbETLpRcRVH8vrSSDsFgehuTKF
6VlkaZX9EfZpDzA2L1r+ntiIgGt8KDHRstePodkkOkxQ0Jnqn98kzvQM2xDPuJwL
oEKvJztre1+BK+NH+dSEYFGGWwl5NOkwQu6TpBmNtzgGaZri7GBPx4dA6554vQOk
fwW4C2PEZLj/sfys0FMOtUr8mPhOSC5l0/iOdtPHuTPeKA5poiogGk6wCTdia2mc
IVjrM7qwIpoPQDjPL+LvArLxBID9X+UTg+NvBeY9X9mizwv9vjlJ4GhLlHc6QL0c
SO8bvPCzKI9JyMZ/ARKcifjA8AcGcJMGZWo/qsnXoGiMXJLr5hVtGZA/s3KlNjyV
5jBs2yiGvsroa/aWqz+qKe8ka0S2d92zfp/GFotsb+pPqt2sNfPOPzddHSwpD/tR
j/Ji+Cn8ettt0CY1gbyALByp8gvoKyoKeDd+0pcVkU2EMzncrHiw6brishcz+obw
ZX5odNg0lhZqN/qFIFgxufrSabniPpX78YNUHi8bBJt1M9yYjxsL4622RkwPc91h
1BMET8Vs5nse5Eok0eefG6fyBPa0Uzn67CkDJg1PDFcWnIdypRbW+yVnn/Q7OL9v
QCAX4HG7F0vZUOvyxlVX5qwcooNg4yVGnxO8PpwDWi7CBR6mBbKALJVV/ytTtCjl
8YKn0fAcw2KUW26Yw9p89B3GIBunEwLIs4CzD+22rHi59Ib6WizHxsbvOWPXmI9E
JKVEW1k2br0KoqD9p91SSADFb1PjhBvc1fwRLWaHG8O9uImx2bw2jgtkU2ABnB2s
CNPHJSA8FpOILW/auLu4UMmfeekFmz4/VWiRJAh1LtVBNQDoT4L3Z3xJhN3ABdRA
2GiHsr2daIzBO5sA28XHJI2oSLWWqwLSYRxEr2ABa9zK4QBNHD3ozoyppHX8qS4V
Soz8Bxn2fHD/FhzO+2FjJoB579hqoHZSco3yH4ncx7ZldleUdI6lzBLPcT2kcjNs
liJb8ACpW2QTMXfNygFSyOXRFI/8pcNvEEzI4CfsClUtanZqxxFg9NItPx86jzW6
JSXu1YdoiVvdB40XpPgqEbo2TKrcPx0WQE1ELVOvNRy183qw/4BtDU0vu3DfpMbx
EXoeJirDYXRJEgPx1Dlgy+BMIyDl6OEOTrCjlFERXYY48b1ZAIsFq7ySYzMWZFYt
o9bdtpVdWUAbXElGyEV/O5DPCzEurMQK+zisPsdgOGzIgEtoG7XPuwZM1S8rNZSQ
Ae9ZGibqex0j/Mb1SzRsBxxM6l6ISRD8Tzakg7utMaIte3rEVayeSTtzXnAemJ7S
bkeBOQ6e8z8NXMbt1uWK6ieSbXJmn8TQYLLkYhCvoOdUciCmwJqpEv/kih8leYtn
eej2dvc861cqbQYONvWxse28aBhWRAviQtty3qvdUX5URJs5PFXsrOIyC6b6EiIZ
1RwaWZx5OP7yEMcwX/BUZSYK2f2OnXsaAt75T1u+/QKrMZnyIizfCyPuqaNz+GX+
LUYYkjHv96lVWGpcBpOk+bUPqEaDZyYVMqwnl/FraQ6pqZZ8AKLU4bwYcbJhTkfT
rG43Y4Wiccs0p7h1QrvpoIJVewNIowek4/0diRMd11J8TFlWp9+NOez4zatsPnKE
8bWNzbIJympFfvXFahvbx4hU4gGga3Py0yifRmTuct30aYtjmsu5ZbMfU5NpxRAP
SCj2klz7GwBGSY2Fkgzq4+iR8fqAenRHWQe91kLeFtE+BUDOT8OrIzm1lKCHnZyR
bo2aoYQ3pLR4LuhK5S8Wk7FrFAv+a8bhGYxE5OutX9KzCqyS3ANMI39nIl/w/wnG
LAaxubdECAjf1J7/6sY6aF+XXxU6ct9TNJ5hn+oygckXUobwteYBMARTfmOiza/F
/WVesd51rSn94R7JC2fFuFcWeSp0umXTtVF/MqmFx3PmJJjHcKO/cL7bi2dxOkBQ
+i9vnV9DDvQ4rwSoQlrfupHFacca+Zda5tpDTrG0JspSeEaZkCGavb/6ucAKDXUh
kaSLmIyCFkANk4YEYKryJP1vkCHgSFGLQOostYSlSnHw0DiGi0ml7+s2VN9nTJV1
WfviUhhkQ5lVWF1dp+4pYPu1S37tesPPpal1Dj2xyDkdXl54OKJNS2cf+2pm5q+X
jSwRFvNlMfqw3l4OiYFiddy7x0wXqyZSUsSZ/rZABkFk7ltUINDOxHPcB3CZQgpw
UMkpGEgOOy8alfDp7f79VOdSG/ZagIKRA4xygcu9r5v6S43oOhXH1UgjCGyNcXbj
+kY9iO49jdnBiUsZ8m4QmrLJ0+VNU2gWfUScBpte5Sdunb5SyiVq8K0Q+5m1Jqh9
VuwDhisgh3SHWzCmwvcjHpYbT0dK1zAeeLnV4usVjOM1KYUYyrepy7RZepYMqUvW
7kakGwjLpbJm1B6PMBQW1jFttximkWXY3x8SYf1JOM/44wYWThuxwyQnR6vv38s7
ZzjTRoTzjuzT9BfqGB5fd/+bSHOS96WT+Uvp+AnhnMEdKIOCc23Hk1vrosNCPNQF
9hhebPBrSrv6rVGTfKBAsClkT/HzQJTzKi5dcIjkHUm8EM2FYUg66YUN2sCO7Tng
lyVrReJOLQ9D0DlYe1WG94YU6OW7cV8XeEbFjVlb+WbyRnN/TZ3spzTMBkACrAi3
gRW2pR50SOF6b/XRxqnvEnpGUTNLCJ8s15cuwdP5hlybLbV73/2dbTvkp4xcI/4w
H9Q7ZRwqlSMwt4uHWBlC6ftFZpCDq0HzeiEAtutfHetU7tyI4FRZb6/9aPiw1pKY
C5s2fmstWwOTkJOQn89e59oIXhqI7v95XCRYNmyxDAq55PDQBs+xtZYQe0gqTakV
SEqTtTYXTXyOFV51EXrSgYQTk4TSJq1+uh5E5KvZks9WtGnidLxRnT51F/dIsMK7
8GufQTAS24qIwG+l27JdEob9x+R1BnlRPfMsc3vMsT7/yaKHF1AZ8XvKCsMNdX54
ym1MbZCF3gIqYNLqKoJEn9ty5Bu2igoRGfIneLG+CkiVTo9YOkkgJ/cwpJq+HuZU
FJQFT2AKka7//Fn79vRaDM7hvg6tqE+FWfsC8OpDuk7Nyr+zvrY6aaTGEQ5kL3WR
DC/KkPDy2krE3RcM4ftH3Uy2U+LFG+gJoEsY+ha9kEAGlB/yQYlyRIbAXS4RPAwg
CzH5ELtFtBOIbRx2SNkd108JWaTDya8FwjMYcZKW4EQtXtTqFzTUJGmT+hEzQlr7
H1psNxczpVRlfcw8O4oF8KcBY0a7DRiU21rATWr+QtnPDxKpq7tlbY+9auHkS+Ir
c/4bWXkM7vryJ11il7sf09KFgJKVXuxI9i7x9TbimewGlU9M233aSSkcUz2WigMk
OzxFUmcsZhrob3nmho1ay9Gnb5z/v19Iz+tl/aMT3xCxzX9f1THHV1qGslYxic36
bxfktvvB0ct9PZJvFWqS8NvvoH2MvbLNZAaOpg+w56jehtDpH1wpp3Sfw0SKa333
ANV2bJvplujivUFqnWCLIjDjbKMz1iZGtFxhkG8Dfyht95VqF9DTFsDknEQReQlw
EVHdsrdPcboiuReGbSUy64bHis/PH4DSEJR8K7kQzfKnEfFK7GhGnnpjmBgP7NXW
9+XsIwXiHTEd6Lfl0KuXy9mfbtGoYNTmD0RXuH6bqiYUxl6JwHA9BRgsghsJGjYB
y2vQFTPgUanNHpoH/qXj7ifvjYW3FhtG4ezmIThX0dEHED5NaTe+6P0RadkXkKro
9Xb1/Mdg0om85W12KqR9YyHcfM2AzLjkInWr8Aq+KsGwDgE4wtRfw8v5Md+BqlQL
8nLSSyAzceMkO/H70e03NFLAk4iVl8AS4049BH5sj7vARRGc0VMVLnulO/p+Obuu
q2noSTBJPg8BlX9zIV2Sp5w9VfoEGAWFjxpncWIvK6T0usKdJ7NYzGOKRVzJfNDi
iVkrDQhgL8f/mMD31gI3QXsouoemQPK6vlqGICi7TD4NSyBqYUmj9IB649ZyAG0M
c32gM7Uyv+NNo7WjdO7A+5VaFgJEJVljZsKJtefWo4TAk1ciNYvo0bBfCigHVfAi
XzG1BXi5KBr7u98xMMChHoyHGINr6i+2HuVgd0cOGP5URPxmOSqZ534eTcWeNNXe
Xc2lgOVOTik8bMMPUC9WvUyTqoJjcyr700Sz8o7lyqv20ypfah/2SOggg7cp/vR+
aGx/mAUtyyvg8KCbguPFwMutUzAYpJqbO+wiAJuVE+Hf8+IigWgJ4/PUgQ6K5QfP
Zf7op8OZGjHgkiG5APdI7NsqgH0gyq/oZ0lRKfULg5As+qWcbAE4BKUhKtny1QBn
G5Ggc2jhqzXC94w1iYdQ4hQYZyGme1aWFKU2JjEV9sRNekdgzNPun1BmEsIFkOKv
U3MOaqQtyApYMKRDuWHFbWuieFEB690szuRY1buJ17St7J/yN+fEKLdjyoX8Re/9
XdybIWzWz7R2h02x+XKaLpsl090DyaJ300SORcCgoDpfXbC9FA9l2jaKhBv9bWYG
Xciysjl6ltwxBBTlUd9T0B7+zv3tjO8dCVUW9JZoIiiZsjAS2rK7or3400Q8w07J
ikOmWBxYqsndsZuOrAkl+OQYrDhsBkgHfbEyujaQY9vqM0TAHJ1ls8yc3+Psnf22
6NoCEZdSbRnBJP1gukt502y20SsuQN8srQ3UEGxrRzd60ygveT0FqUIkfcvi6i7o
WtPiX+2VhFnUawmN/iunXPJQ1yIzhhyw+pcWd5/gVSRMDBck6ctryZY5KwTcMSJ+
zU+bk2fE908CQFezM0rYbREUQ/1KRSVsUGvE67S/PIGUU/PFCjdFVERlk2CeCgMW
Pf+ZFVQIsKaQbpFxjDtfDYMq9108IsmuaoWWf7kngDSD7tgHJVJ4zgz74GxjODNv
q8RNN3UAVsj9/ISxQhpW1tRfA8pZxgT+eU0rsO3LDmxKRlTksSG1zt4CLo54MnPj
HMe3cuiL4UfMiWUug9+6xunhj6MdE4UWMGICb9HCtvKyiaRhAcZxEvB2myARxzsi
3C4te8kovbEc5ztM9bflSukWS2qfruC/k997wSarK1/zbOn0BUESudIf8LZ6A1yX
XWhOI+8uHXFdKKTzaHSZ+dz7SwmcsSoIInMraev+oyGE9AIQvzY+HVqCOY31di5F
UC8Au0qHQ2mIbMG7KrvnYlP7JxtZbfyx4zBg8pb9JYBzCGwtYFwnkw1VZ44cwShN
P+QIghNKiGK+ROjIAxy4uHYk2lkCg8sEMpZgeV+q+vQXYjgUVCQ/2TWr2g+io0Bj
MTcR8TAMhwFv/T4g/4SHV0H/Pra1Wq58rlSanom+l7d7RT2CAr61/8DjtXsZu2qy
lOhhMgui8Jy74EkrLOEO5CreUQClFXdoSHcxkxGBzUYgVe9h7lcRCwIr8uuViH5h
myP5AfyOemRNiVnXpCium1YDmS9CSpQQ2udLiGqUdptr+QSF83M15GgeNFxZYEKx
bLfedM9NAgR8u6UurIpaRbsOY5IaRKAwU2FMQeylfqAGBj9Ufy1GIV63Zot7OS9C
fYM572S00fdB8+nI4QqGrUtNyYBh7U4ruaEwO6wJplaEUxWIC07sIryiysBJPAna
xPBkZa0Ge7AD/6tees7kM14IE5LGhNSOXnqi89Q+E+dIabS+O1W+Adq9M0XnDjeG
//mUpDXvfwwwge2sjO1C3MfTs58q1h9vcfKkTHUxFiuy6ucllv5V1zF+X4Vga8kf
XmEttpIBNOlD8AKKz6XRAM38BpBF33Qp6jqG4wOwO/9lfXHr9ORZ0pyT2JxvgZug
/akv4vOgnpd4QgmgA+COW7RmjaJ1a3CUIJzcj4JC9U8VFXLhHULdkzXOC9uZ9OXt
qCsH3psOeavL5248brqDSvm458YEioDsUlI3y2vHxJuITNHILlYce5lrRZeyLXWK
pHgkMZ8BREEDF2gfEg5rSlTgnF8NQqjFgwYHHNBOF+ZeQpcuV1v9XHK9eyxjnfu2
xZtkx339yc+LLiXVOAw3p15gdrmoaS7o4t3HmJ9YnFtJfE03cERo1yvNgqTrc69H
4FXpMmY0dPVRDD68PyXyh7/4XlQKH388ZJOYguBNr0GveJJMQce8cBDAO1AUUQr7
GJUG49QVE58TE8xVmcjj0KYDRpYBMtk9li2cj7sex3TkoLLG6Mgy42B3RKe3rWhI
aycjFjd7Mw46pyOTlk8Ksz6OeLHWnfIMXKly3gqiN8nHGVkfSbsQAayjlBISjNzT
yGFYoXcJBRLtGxRxOh7Ms9ijx9cIqpqkeexJsDk6BsS59N8+1giX0VuKcn4ztn7a
ViD1985RtNQ3ctil/nuT3qsot8NZLTFa/6Nra0Cd2Se84fIWLPgFQ3PSkBcjEto/
3maygpPYriD0ZXE8bEgqn/nVSdawtJv3wOYYkvjyE0fyyY+Ts/0QjNwQVMMX2ESZ
0Hh8UX/9WyU4cAb9a1GPUecV5FoART7bFisOBDIyF6EFKNXWXem1pmbb+Y8Y5wO+
PqZtgbgDScj/mk+etlnyuH2C+YHbtnXHXWLDNQXPysPHXX98MfrjQdYKIAcEgBw/
zA0tDgNuU05vUCiYmZkyFREGqGHgg2ViNwLrnh7dNDCaq2mJpln+CQwULoUkZNGF
mcOCsF+8KKqWAmQk+BLSqJf7nBMXLwby0Nd+UL88Vf2EN/Ei8MGbqFk3fpH6AwnU
jJ9dR+SJ1fcvFGRJvrExMfFfD9lCe9WVhFt1RIP/Gll0A6u3gbhLGl3k0Q92qo5h
LdbIOr04g7e8N8Pf5KFjv7aZ8cox9jpRS4M+VF2rxDi5rrcn0hG+wW2Zg/x/r7o+
MdEjpvDes7ayHhY6HSKmVBgY6O7O5XY6HaT3c6Bpy9qGQP8x76G/Q61EENes6+YI
GLWMq7TXn9lAAgcbjLGl0jsdF0G/SS0+C6cDqLKOR7/oU3Ab38Uwtd1DAhYAUjOg
m8L/7fmfLhyjdkOH32Dzcnc7SQliRQxamhxeNlrDFfERjPAiVRkX889XoNiEHDSh
vMxgNFhokBGXq4TxLzSgSfsI8g5vxZirK7Pgwmd4zAqbmV45PIhxUQDy4vOfru7S
P1LT4OsqSSlIMGFJIwhUbM2ggGqeTBMCXfswEcgIPgKDyQzL65WdPp1F3UV0MH/w
F3QX+dNRkSR0etr+ARck1wknfMm8FYv8S0mEv0oaoCrhmXQyEwEOyldFZJ9m4hW3
IaxgnG6JyjZR5+5sjXzYYeKhZRU7YD2R7Ht+YiXWHTRt7Rsue94vkJb9ilXuXCR0
bo4cqB3Q75mjmdjNcGAoBtPAN5yz7DGUh2qhRqv0LA7IvHS+Dheu1ko6id5kJRck
D+vGchwTyVG/ZEbooh6S5TIKXs0HzkVsUhTEupTPl/D3quBLro93CCHFx4IqybQL
F5pFIfHIlvws912wdh2RzYkvUrVwEf55r2llzzPv/MtlmYok+/NOTnXZEbKAh9xt
6nlP7eZLpTKsx9+KcICADd5fuLWt1V7QsmOQTTOCKUT3hwWY+TJGhONndlLDzMYA
49lwKjkys0Ihl7xl2Y8ETvGNnYIXcG3O22cU2nUIQeozwYAbZ3nn9Q2sZjJ1Js59
o6wjj+Aixa/OjjzM2Nq7p9CEqgzxL93b1gzYVq5Jst7iGqjIeIEh+W0WqnoYfusO
otNZEEygvl6ICFZq2z1VNfO2cN7qIlhJQExlCf/GfZL4fP1b3J5NE7HxNdhHVmYt
Ikq8fBmecm/OTpU+JNsoSmyITbCbFgEbWQNNXbLCLXg7i+LczEDWW2KbqOm2nhaq
f6L5FLl4fUnm2aA1vJhjxwK7bXIhnDcpqw9xv1dsf6c2Kc4Pgs8/bQt0sV8arVvI
6g0ePwceRSAZ2S/1D4C1O9BwIzJHIhAxapAAzAXSjMOGI4KMwuf3C8Ehk0n4xW3m
uVMKdy8FyQzkrA5oBZhvb6bkYTW5hHl6XiT3XjQd1khID3ApI30fMyGzTBpcKIdx
W2MWL6t8G/Q4LSEpVFZg6P7nwuO5JabGTasA8lQTFnZr8j9/0u/Wd1LshDiRPNFX
9FZNZGJhkKjAbv6UkfgZ6W5lnXg+AncB9MTU1Zjlt1DweRr+hClplIZnBI3rbYxm
ZCSSrbcjAUAr8wbsV5vv1PyHM3CcVpDPzDia1P8tI99luIVjvLqXq/mTq14oB96k
IREYfFeCLtQKTk9Fmpp4GYwmk/rJ+nbkCMOkx9sbFTlhtjwjngQKtdotFd/3uAYA
3yLanWuEmJi/eIscDoBfNdxiHcSS3sBrT4Zhe9+BaKf5v9zqOzcyyBQpO/MUvPHP
vi7d4NY8yFIYjYtypmvQaTxRwlIDT+i15YTMG+l41wCtBuP/kXYeBFQ8qkSS5/RK
jFbIRMG1RVRODrtZ+Q5tFshbByv0VxktTPd05MpMzSYfFU7iH0JwB7JDUfyDsTZu
Fy5vr+Wf9ECGStWnl+WWsG4AhjDCkNqtFM3IsyBn++9lu1KpPcHbgnN+N8YI8Wb+
gM31YXEGj5cOm1bo3VfYuJvyK3OkqxukXhO0G8pRN6NglJG1oFoBtGsPHM1t+qko
5mLuH1vl87ytEcxXUsKyv8UR5tgIRsSKjzNvp7osTmSDyx352hD/loQTDc3notP7
/qz3In4QlfognGeOao0fNQtAX/DS1E355U7qkFATKninutZKRk9VzEUkshmlBKQ7
SbSN7TGleeAXYsiTOlme5Ag3tw/cpO1Q1xPCeIBbvr9FTyU/tecWDkM+tnpazfVK
6wut7xtTqJaWkrUXLO2tsvY28yXetzHZZFFiaNGYJhqGZehGvYWoDm0zuWTmUaXU
nDfVPRqh2UDnNbqbeRYHHipBFPTkVI1zQOIUxXELoSaXHo/tZOB/qiPjVCYElnhd
G1JYrqmSkhrM/ToY8g8HK7z26SwfJdaK9QQx/2erb7vIRyB+vKNHpIWqHMQP2FXF
fKeoVriBre+7iAOz4xWbFLzGOQ6r5+qcvy7HYXVwJPBQSW7QrLFx1nFkZBP2+drQ
312Gc0nARrVmTtReGZgjnnsMmAjbKZsD4eVyjGNhBFvl7IfbJ6CNcbCOKf5MB4C8
iijIr09dk/sPNsWQTtR7bMaTh8cPaYO3+9ZHmwuayu6J60pGp0CKCKGn1spxhaPX
Tao3BGJy9DU1qeyUk/9yhXDTXnnMKmFyjsJ30gQtZykkWflpo4EHY1jY7AgSAszX
XcvoKHj7iFBcojJzH+cD5idHYij+SJnEABzqMXMdAxaA6b36A402IPW8SfCZymIk
wYq9St9BtF0V1rJTTX/ciT27HMUdx7OCndyJL90BSu98AWzNV0eZvFpCRjC0J7vj
3ULCrzBHzwCcddtGx1yOoWDaV/Zd0IiQaG5ZR19Tx7+WC01Spqrj3C4YACTc4VUV
mAVNbo51/HPdOr4RyD2GyfqNTBgfod9rOvbBACdRswzgG2pm6DTf71NeSntB/jqu
/fjpUPwSblSAMeOQeWAclENKG1NNLpHludg5ZqyPDa1mVhrGhzqNUDV9hKWqt1wM
G1qbxCSMOSnDLQcKJt5cftyPiplLC49eUhzDAGfA8ymxB/+7HiEGrp4u3x2tsPj8
FypQ/RpaU3DH+gcqYSLNkTkuw9Cl82dodUkV2kjE21WCGSAq0BTscYyq+9sxM84m
fPVTO+99OCf7UtVlzTMGtN/Wh8V3qRQ9xtv1ZBDgG/NYgaSsZK0L8bePgTvCqANX
O6ctCPID/KqfLRZCZSm2Q1neQKVAJbya7/S5XJi1v1j4NQGDHzP6Ou8ySU30LSnh
kgplezSmY12Ukzt6N30ryDMLktj3BGeME9CUDPmFn9xgvUHFBC2qOTHHh7/KlAwa
eqlTs2DxeLh0Xtac9vqCy557v7qVNyKmBsYesWmzh1+muXA+koTc3AQaVdc4J3qM
YtiPYWDZkcrS061A5K5lhq9gIDoPrKiv7FRjlh67SCNJJ0cfZ9tJ4X0n9p0U1UhY
Clrv0u8jjeP0jP5XUpb5CtVphcqAMyCO3d0jH9QgFwZYxR3SQ3tCXreWc6RLDTqK
35/gJgLfblmVb3ZzguGIkb+xooWwvwKhp53ANd8LGnEfwwr0YSOIYi9qOp90zkiA
qxsZhSfYvZcRVtG2zfIeAQfFL4P1L62MQGe4pH/mhEjbDo1Ru7ljxgpKRZUu5dif
onPxTBMAan+d/ioeWEU7IJeQOXr3ZSF7Qb8zo6iJaxOPflwxQYpReW5hWi36lfLV
ObvLtuuj0vHRZEUxJ6tQTLM8ZgUOIoZWYNjWb+91ttZfSQTAPyArlorIAqGCaeuL
KHklDNi9eZfNt0LkHP/CUYhxtqp+UGo9AER03+YfioQIafraiSGAzAxB6BM8OarM
cYv+oprbJEVrqEY7tlpbvMC3mf1fpDb7YCYwe09lKs2K16+dYLhZHnnO4LlW85uP
RudahDIeFNmXMUssJa6xHiYMe78wSa0GDqTbb2sapEXu4gyk9nwnkUgvUCc1mDDF
+xR4Ydy2iZ5f1CtWh2LxHhTyhpdbQ+553vx4trHMK4CwcVFXS/FkNNOZGZhQ3i1m
GEETxvB3rd4kS8up4BrFR/ixHob92zdPNHM+tjcQPValYnxQ8iKZHzyYl/rn1rs5
B8+K85m7ns3aJicx+aLDhUpu1t0Wsasm38HLyi1KvQMHhqxw+YILIr0Sxz4tI2tn
AQ1FbIXhL/cva9AVsd9A+plmpZWPbs6IU9zmyo99U7oka4g5ysMyAxQZREAZGGYb
4ZXzbuqpO30QOyb3MRHz7UfQUkFQEhKNslufhahNtLezGkAzG3rEt7N93q+zmT9Y
vrFWFcZWgxdfROhNpFATAgYFVYoExLh1AqxYxprgg7W7vX8zDWrtMqMstzpD7H/i
soyiEIXNnANHpiTAdTflSPI0+CkbjY0bsknzPLetQWBGaCkVxSDdQSSYBvJERx70
O9Ehe/KtZwxA9SUsdwtZJ0DNKND3DtqHAiyHalV4pOd0qAoDEayC78IDR6XnK/Os
H0S+cG+VwirZuhmqgF52UN9qHpzkZMpFByvTJ+M7+qvs59BD9zH9shuRPANOjXz+
c+fHIjkVIn6Vocp2ziliy7SIg+DLtnA/0bAGzAYpy3jADvf6t/n910ya2wBDYZKC
hmnGKqAY9opAgUemdciN8bLuTsb2pRjfRQ0kMem933o7Q7z4fNgTK3lUo6OhGkbC
xk1fgRMseI0plGAM/MkwdhVEyRSnWD8rqonUR9CqOq5vV5jVWLA4X9u3+3kYFpIf
BpIS7Fh88wVh8HDBMoqFW5iKP1p5YSvTgwTrKz9yLv2q0AD2QCz2lAbnGxyjF+rw
w954XU6rn4GaM0dog0RtsmANu15cY4lfebgbSnyfaH/XbNwz8/NDH0LyrujtdOTq
VNVzOgSuQtGUgkdKKesq7ieh9ar7EAbVMYDfJOgJizo5WSHfZwt6RiClgGoVcDOO
W6kxj7/C0DWTatE0h+iRuJg66qFI2nuZtX0S9raP4BN814BoiRiFSx7tjtXbrqL1
fnWKy6E68U0gRq7ROPFBd9cpaF1K2n2MgPmJWAKtk3fMFyAKHyAIw7Av1pEM3amp
p5zIRlodnPRs4JlawzQi1TGKXF5aiMWSGXGeZB3fcBKyY03XApwwmszhzItpHT6x
sP8XGVZaWqejNxBYBfD3QPMFrYnyHIH2Gf9sgHAMUwUCXECqm7rpDA8YxZCiYynm
J7mMUdQv0vceuRBkVO4n3nfBaaTj+jLNpHsYrpSNTdXiQZJAUYyih5wRdPv4HCc8
hbNxVCK1WCYi2iizps3EcmIxoLAExUhSs33UbYK1NrINko4wosR9GhswiV15a46a
XlHoGMct2GTaKehFpwUNU1X0cWl+9JAMli35/E5B5E8eLVzUant+DM5FWWHsKBk7
oKSTxg68koxQa219ojQank6rnUNAPJqoEPEnx+Ww15ilg48rJQqRiKIKFiggWFO1
8x0ljVO5MMCiaksmhglYkFZ/0HfrfCpKB3rClCjNmO5pFnPuMQvJtlOcbu3OVwMy
pCPved01CttJoMAPWc0gtPB5EeGCmGPxo2UA2JGzCBN197lvkDyrMl1m94Mf4MQ4
BepeUeHso91PBI1Kom+gsmJliSgi2X2UDHf5klrEPxpUyKfRdbjgNDViLSqGsynx
v2hGSUHGjPTQx/hHycGXGvGXUMBfdodNwy3jIOJO3vb86WpcvQ54uL+U7atjx+ZK
cLWhRbibNGm0pLO43cyCpX+s7PgY2GTd5VL4v/LbwHb56IVAXIPlJd/P5Xg1O6xS
f752m2qefX+/wYTQJUReOUN3Ky6m2g7Wu2oh87D51m+aEIeKyo+JDWxkGIJhvq70
MiJYkNRKmWVLZcA2ar//pdANGfaBY8Nzt8986/AHbFzYeIBHQ/CaTV6+Y1LvBBrJ
iiTYUA78wb/2zYZ/VDhZhz7owalVfKPnoHhIc7fhIEqh8Z7ns867VH80QDIH9Jnh
H1mW/9eN0zvioFhK5sMmaUOZX92K35+3GUNN30JA4GIdC9dFjhc5AVdV4lNrLudC
JFiXar7RNpJ8LGyV2CNGxttJBiYLWoUFa1umKRZKt/t11rwqBXV8L0l0QvpudgqF
1f5pzJznqoWG8tFu9iCvCYE8P6AbC4ft4WOLm0XPCD5zbRmlupJGYcziXi3qpVRC
4Y9mtKkehLR3k4Q/IuPOSzIqkCyiKdIFI6duLCFHkQ5J12KyFjGiVXhannqCFh5W
B+/P84zgI+aAe6r5yNt+t23hE5h6nOQlyXXH/c1kfUHEckY1ZrlSTu4OI5rGB5eR
+BnQ+B/rqqkVc+y128WHIOAKWxyvPWh0IiZ478XIP1F32p0O2X3svLQrHdFAULHH
YaLTb7OWPfof3iy2OuXAL0wfBCmKqV9m5HJD9la0Q0XPkcNSKEtC11BoLd1Wey1U
nCM51qA29jxyalvtws88Qa0WpJiDoXh19PvFoG9jZiAM6M8Cx+ibt02qRP+WZMvE
RPqZo8ZaWPguI5OcHxFBJyw1j+3UM90Vp3zeho0Ixk9OBZyNDp4g14GIZ+IcN2zh
2+EYOu5g5WBEc5EstCuxqsAkhFMrl9hhp9F/vQYSVzKc/9PeydwDaS6GEEFGgQZf
2n8SEV5E09MitHi8Ak3SJzYgEOmOQnQqeVN2pgS+F7wrWXDIsjlAyoY6khFtoPwZ
SWwBvCmiV0zHdMqFh5HgWJBxEziblCU0fn70254G95JFYIJnK1ogppweHa11qD92
WGaGYHQsykpiv3n5/byfGLemxILea+anedi5H7ZnIR7fonKbl/ooqA0FaanfeJva
8VNS1wDf6J9bCd5RWtqqDniEf0WbfIhRJXPawFEmRcZnPfNrvifHXHArfFhHSG+n
z0pIiseZruWuYOlEFG0K7X0EPSw34OWwIYBdsO33Vovj5hP+zReTaVbdwtRUlCs/
AKJabNfrEswSHRcLn6Pjgdyrl1LoWdiIAjqW+i7f08DP+wwXkLUgWKNQNAASb/QA
ajusMN1/nbMXkNl8pczRTN5h+AFU2ISkg6G0X5CrVNkCq9spbNWvuK0unwzNe8Kb
g9hVY1iGQgltK/mu0EdKoYziI4UVjC5ubdUBoMKQhhygSs5DvfUo/d+PsQFjbxP5
YZTekOmaWGTLOgQkkczI/DLZxvLrI8AI3lDM4jQx7r8feCAWp2nTHdrIOOO3Ybbh
986FoQnviD3gcC7wBj/AhvDcM+HfKGmNoyl5l1ZQNO2Y891yfl2ltRVo3SIgit3R
QbkGKaA15WO8ZVg9NP6pC17wlSI6cOrBuS8cFbYh3hRajp8dCcCruun1a7rQ8bdQ
05I+dxXgAvakd3JdSMs54bn2guhVj7iEArb3ygfaMgXaVuWZhPwr9p911Pb0xc3A
BCF/0nzW1RjhcXOy1723mwtGcVyigy7+vGUgZOq/iXF6WuFvqQ9xe4g3Q1l5QsW8
W7MgXjspwo00gL5MBqcBItRioZarHXhn83SXjfHDA1jRfMbiz5xBP17FOoawszj3
0jLLw/3gu1QUq3o67G8BawziWpscy5LeHil0RuPFScQPmdQBdn9JqK68BnRhd/IN
oo7L81y1WoXViMipcVhJVMn78ifFcIaCpSjWVkP+HhBr1xQCnDuZfMpF3TUsl7Pl
y3YDFet1aMtGy5YtsU4exrgto39FZtW3r4zK8VHMfNznfl7qvvH8jY8Z43mSePSb
Ox8VLtYJzkvsnaMkAiOaWR2OwFMIz2ZBHLW9J1qjgsXbhAVYgOaN13x6nNQH8VsT
4YNvC9WTBX/zYWVHftW3X503Z5XHMnopX0A3icr+SagE/N+kXGNQy5PhweQNiOUM
lutw9l4Nu37cJuxzFgUB/kDAcaWC4ZQz219ilmduIix4cbRtKbgN+Jw7J3RO+96M
dJh2ApWtBnh10ewjMA9oNFtAqhKacAt+E52JsLypXKQjRmwYM+hF794EI4eh6yu9
vGJE8kcU7+g46Kd87eWdPMO6R9q0D78lOkR7w+hnVNA04YJqat+LBVdbG0DIAOBu
zezo1rKCne2tzKPO3G35SukdbNlbxAK+OEO+00PWvDyOT/xhyPRn88rrV4KdeEr3
4RRaMmpZWdML207BfZ2o3spRZLKx6q8zLC5Gd2qxTzrrshekehjxU/1hvjNHCVF8
AJemAGMbAjT7goNBkUSNM7KWIDBF7+5vws8DswUtM5fNdPWvHqiWZXt4TMD11d+L
fXbuAJKqxU5x1gTidZ/+6RaKDK9QexQv/Va2LsWbfFQps6klEZLRepWkOnGV0rxL
OFX8VZLmwlUElQ39AxqQVcvLI0xp1RS8swI/yIFZdWkD8+k+nS1qimxODws3hbRE
/00WbSpjikZ+6jSJ/n/KSiHxGb7eqnYNup+foYlPdRi5UlDbJ2Sq8WfKu8qe4K+Z
D3vljcePUykJ8DaQ3MyntE6rvVLWHflCMagMuTtt0KBnnn8UJUyxDqdzV0ns+sGX
cAe0T/CFlLuFHvCWXGH533clLfrNJQ3VWHJu+rOw906jNKb36pa3xyAHnujrXu7P
ZWQVkW3SbWkgomaMROs1ZfpIXHCVkBJOlfGiv0C+mVnfcuJTFPJ6u7TDGTKu29/X
SjN2J35+dtjT1o8YMglKAOTj9/JRb5eEkvwFR+89LNao5kpy3IwbcbDFO1n1ymfJ
k4NpdbHb6hJg2w34PWr6tlfiR90bz1ttKcDcZtr0Lt41W1rSOqAv3D+pisRQv0BH
jgysXx08oJfT799q7y9V3JbJYH4HzEx/jShtxhtAPZW3AnF0yUo+jYiSeefze7Av
GEtOvs2QfuUS6k6vdc1v/Pr6XtIz+4h6A1RKgDqa6V7kuRkSr79bhWmxpCnfQXQt
UnX098ozvWXXjPUVqIi/rIJODQAETzvJ2MCcjrPP3DkiSHK6VEsaoTfWdTf7PcvA
9KnwLgE6+vFDimWDXFzS1SP3OlzpE3xhXVWUg0O8POLlpPsFctJUlP04+7QCxWQk
oYPK3X+JzINnlV3Aox24RzKqik5uFkNXXhOlFODdhNHbzhFc29gu95d69QKroUBv
SRcvozog+RGSDOkRFvvG9lz80fyXZCvyOCpKuVUqPTZhb2DoCYwML5FHcpBHmfzh
2u6dpd4H0yauryChRUgho9gpDIcC/c/R0GWKeSXHIiu6Qb8iixTmMTmjrOVMaw6O
fN3vTCwD+vqFODc89if9eyxfZP+zp5upJSQBm+ZkiUxfHfawxd8ETNtOM9n7zsbK
96Ui47bY5dmmCck6iijbXtYux452f/e908euxpnBK1n9AJCVKzsbGk/SiyJWdi5D
US31fdDlonNBQqy+Wmg/tzhMHXs0kjXVKXpH0eVw2c08NbY87jpes0Bi4pULkXUu
lNcaQWVkEHobxHftr8PK5WOknQiWvaQUc/c6a/Uv4psLT5k6wyWivWgs8Em1IB/9
Rg9M/cCpgLeMlt9ya/yzNCyDMut0oBScZhX7EHiuu0GQMdnUYP8+RtFW5Zgj5yN1
J0kQadc3wgt31GTtM+67M1jr2bOfRyml7CQgrcRNk91vandSIBCzoGK+hDiPNHdH
g4cJ24nU4y+HdCY4GAK1SUr5HRWyqobYckvGxMegB4VBuTq5NDHRntJ/GAnMvZc2
RirqmMUQ5XMeJStZSPvhiEMWFkZpKx6+UeO3ORc9kzBjE12QqW1d5buGnzKwWBQA
uNabyxWeDVjES6XHd681Xkdk98Dd6Ybr3u9HAM2O5iwTin8Xpm4Yl73kQE4G1Yad
b9owdI2wecG2EvNmIIwUZ1h46bLL1zkvYma0ZNZlcSqlb6alRlS2NLRQKJQD1LV2
ZkjEA8FFQ3pJadlE5GSnLoZdvjFYCHSZEJIhcw0+gPfBzjMaRS2/7WDkQWpfbPQS
9j5F6t50GEVAIHfiJlF6aou1YJtYfgqG8uVoLS+syK42e65msTijM/KmMT9TqSgC
o5spOytAoNzKUJ2D/Z5auqoF/JQbbYZK9VnidwH6Aw2IUevlDAC8GArsHsazD/vR
Gh4TwIVCPJgmPYUjEJmmV4adfXcg9bnBK5bd3Xobr1Pxx4xDN/UEZxktt+6BsDAV
BA1VWWmX9Exa6LGVrvdwEfP2m9q9qyIJkv+6fCP/bZfc1w0oC3Z5m/hhxMaTLRY9
vTdjy8rmIyD3kQJNDsjObd4DINTfrNe+Il4BOM9H1HxBm3J8wFWXLT+BYuDh8w6E
ZMoT4ewxD7N9KVOp3wvRz/tUkf6vUg8oWbrzPi2TcWkvfTrxWlkLbXVLXfKsEwLu
NB9tsEu/MuLQ+p18INGgx4W3gLvTCvmK0LoIGBXH8STtABTcd2GnhpFjToZCQG7X
wmKO4Gf+iVuc+vztAmfffC57B0PQjr2TWHwB13E//JgjCwcKm6cLAXtCmmPs4YB+
9EIZGqiwM6fNCSA7BqhQ7RznnfX4ebhkm8cCHLG8xR1ntv3MVg8xMGacHhxAM7hA
RBU3CqXwiZbWesI056QFp/fRB16KP4Tmlj3fNISI/uAK+y267ZdQPTxomexSfm2O
FZa/MM87S+YeuxL0WkgxXefPMPVao7ifEOiOX/Rn9BVtPHAXXYz997AANlKITis4
J+jH8Ct/BljtHHB7Jk1BFr+/9NwrzBtQjJLuqIi0R3GHbPhOXmSs2gk64KH8I6nh
aye7xxZLdGgome5uzx+JKQ3O286ULInrLaTNhpAHr70hTIiQgVTV9cPz+4dchwaW
lbv22RI0Cvhyyo/Q3jvlH8314gySpu4Dp7tQreEA1J0N8PiNZIIDncasDTSlRfYh
njiDClA+TB/2ZXmfk6bplmPRbQZ2+wZqarxZa07utr+EaFFhjw06LoSAkGyJxJ4F
MIwGedhMPipE8l61awrDlMpWQNcuaCNnYhHLBRlpOxu8KQCTddjmRz650NZUutxl
mI2QRR/WnuDgaLR0k62t6snrNWWVnFSQHG1cs82La/lROojthdqUVOlczVJ5etc+
LpwgqIwAyszpxN0p3cOiZf9+gcjlLwLbvMDtXJwPWkBO/LmYiqdO8hi9buuo0H++
MMe1bcw3MvJWJeppih6Wvh4rtmcgeqpz6hsFYqmu7h3GrlOcqH8/DzNzN3SRdypl
vTWc2iFqdNWlu45Mzq07azOBUAS30cQGVoKLV3zgpRH4HyGyU+Bao08CVXPJm+Ep
gODmi3pBQVXSF0zKSuvkm5YW2tWEiVC5DlUjD1Ksk3XB6NZ9APEi7Ig+swJzojtk
I/l1Yp6mJt16dpm33YOtgvN97PhPLUb0UIyO4Tx4U+S1eaNb1dy2s7mu9TOLx+A2
Qezm2QBvSsQFIuh0rlyf/s61YQWUTL/1jVTJcGeAOFr7ga1cIFUQqyAsOt4+37WH
P0O+BRhyAULjBt57maskiPIlBj973tsFPf3vnXvE7NE9u0eMGbUKjlWOlxnD+5bl
9duWXjL6K7g+OLpxU0pAOG/TXGmxOjhlFfGF6xH1JBsJu3oU1JYW/v/8zXq+a3Mk
z+Lx4np7Gi8Mwb/iYU2pMjgAUPxMZVQ+cjJyYLZurJFIQ/lBIbGZapJAq5opkZNU
tijEy/qEPUyp8Erw+cT9pzgBv7btB+DmNolhJR5MoCiQZrnJoJhsOjAC0QRzvH3o
zPfjnKt+uc9blqtDSljr9av7Hi8DJ8WZ0r94HC0djF4/Qbu1FZwQ6dlqo6155lXU
ePzdKYgAbWktGXkUdXkLSrRhTVxmJ2rwtVqxF7YSxT+pjKgtrqxaxWgosbsDh2/h
RO6lWGpD2uVIJuY6h5fj36SFA4PQycXi+YhCiGOS3Qk7kheYrUHa11flmIDFLZK9
N3p40FW6K++Hek21SYXPXAid7xtmGGyWPf1Y1cRTMdlEboDueKHZLWHnBwr0o7I+
KDZTpavhjvXjXlG0sJW9NZce+ySyvQVAAbufV24ELy2tLci9PrisxDaaa8UyA/pP
2j17EZzrlb+s1ktF/ZHtbsJdut0GQ9o1GRIf6x1yF1PgeJSxCymn+wofrIwAjIoe
1NXbe1gU/trI0fSEyLdvoGNlXAf/cw1YvP345CH6ND2ySdUCOFx56hZ6MCw2ICQP
RtsR8LV2eJtbqE+VP+MjLo2KZphVmsvBNqeg+9KkXvxcRzXb+GLIVrDReLkQ6oGI
ZMjWTiU8+hXc4gFBJcPGrE3veXdZs/6vj2ja9+ht5A4YtilSrFPtm/0GKfYOnsIA
KVMWvty4++kGQGyUsBKK9DxkgOze4yoj17fCozjze2N5P77fjKgEabQgGgBp2ldZ
gqW8PcIcX6uAEkIpKJXJHV1Yll4CyvCZRl/YY0hmhBiPKqzKphZfLxkACSdYZxOv
nwE5BclrCwBJ8bTToimLG4PWsYFBDlj3EDvgzKc3nKIlb+AW520iPHYvL3o7KaqC
7lqRTCSJeQANHm8H4MBTn2LASNEQOWAAJ+yGY9efP29Cq6kOK/+4cU9PcaUmcG/j
nmEUbVJcm1ZyJJn3yfkXw0nmRo86aWHba0oHpdY+9EXdlXs1Lx2BI3rgkn6pdx+A
lEqMMwxZk1YR6Mnld/Je81J+L0AHDBRGxvzSsaYqSAvWO+ACThWL06QJlFKAdzlB
pRZMJoesK3BLKq2vrEAzj3HiGPSYb+whaW2ZbWtRTnrwnBOH1Ale1lBhPvVdoTQ5
fckzixXbir2GGlJZrhLD41EVGSYWupRjTbNWDmbhnAHMAjW7IUm/ubyqF4BGKUmo
8nwMkNT45WS8YckygBsnL5J+2WPgUhtmw1OGW7p2ThJ8QqeLzmBE99s2SCrQePPr
u538iEIoZ3KftWeqTp3O3TpuX33qtRvPPiKmuOeA5vJGbeUvh/mZrKUYboQP5r++
mCc6gC9DtM89ZSR4eEQRxc0/xgppc9K2/+2qRMRbqDkDNuTQXAG0s1bCwoDNlFI9
2qUHjpH4NIoDBrSggsF4zx+CNso0uZD0dW6LZoF7kghFMedxEGYqFQb2QyIw9NKN
mrFK0vu3WxkkLRm1Xs/1tzlW02sx+lKyE0/GoRY0OV1NjJ0waBcVn/WQTBbp3QZ0
jjO+rC03ntwtuZsq2pjr2hLY+6E9h+aIXnpvbNmLZoOsp7SveJlwtKwLVkHeSChc
o2PatzKkTxkjDYiarYyeEI103mSPSuxXnvVLlPUFEWuw8+odVas0eundNRjc9AeL
BrlHK19hTPWgkj34OePzmAE0rsbWarRy6vM6zmk/mb8mQ8AnpLk/mDzLUDvgQzH7
7FIIcrPV5Y81VRBBzwcaEFQOxghUimwY9eL1P2vLuFF19uszQJUKRvHFWmtk9+AN
iQmEo7Tqe2O0MmZBEvnu14DrAkLo+CALjuY9kCp3PQqDkXuHYDZLA2hmWBRmCAa5
+O60fNot+xP6GmKOIl0BStoqUToJuekqSqSFMP/87RaeBVTnw97jM8hEDBkIoLV8
slGx9SaWmMLU1jsJCrTWerx2kw9ToidWEnhkxi9ifQj3u/hMAUemp6hoJNHGkPaI
hJDatM8N7mCHP/1PmGqoDQHFChwrDm03LGR5GvMST/fCwLaNy6GSwNkSjkdVt+9A
dKmGHgcYTZPKaIepab9jr7aRKWZ1Z3mRS9fnW2pbKCjIncGyWO/02K+NYa4ahtnS
nlwxpD31xJrL4rhHVEyLRlhZLF+zShX74t7WUTceUUzZbKEKEToY6RHz01v265AY
xRmDJbASovRtWMr3pj09R+0nSzJkbkRGU6TMeV5Dh2WRNsyIQciRZteF4Jt2NGDI
mcRcFCH1QZ1b5lwjg/m5jXl+fV43C97F7HrmiVgIMQM+ObvOS+gV88TD3SUQzOkm
0W3IX6cEgBBFcTQxremaYcOPwHiQ/WMsqvsdlOISn1Y7r39D5X6OdvNQu+U/JzdS
hasbfbM/Co5fiZ9Xp9tDy0dcG2sAgSFsDV9cnXHjOamZsYsP2Rz1Xp/KLHgbyPRl
WEjWypRKhMA87XDs0qOrZrL6MKIkYZz83eglqxMbFJHe9359n3cZGb+JJ0+OPJno
RAUybbgp0WNMW+xrzNlPp43KUbk4ryStz2f7x1albMNWhH/e6ImaiHdO+WQMRayw
vAVGtdnLAx9Ovc+va869q6i2nXeA3hWHgpwbzC2myK2OVK1JtwyITKEeM4YFCYzE
cXp2owJUdtycCxqPcJBEG0tC6mqpEfk/gFc9HBa9q9iEHU3s026XMRU0jbJ/q8M/
bcYektFtkXUSNgrnpgGRHERqGdjmCHN/U2aCAeuNZYjgODrRBqfBWWgteITpdWqF
rUFAQ0XRtnarVLLOWY6JpynIuksRCOdBKZZVCeDWrbeNGnJxbPFrvZDAGJx2A/3b
uGUhqi2NnvUYYmdL5FC+c9j4HVprJC2CPVpYPbi2RwWUQC/i39raXFJY1Zhh9yGz
xblBvqkEsWmhjsO1sG/E6GQRSh6XA5Fg4gXZM/Bzhwyg4gr2e6A6p8iLxAaF4NJQ
mpcNMPEaItecWlJhT+cw6MBpbnlVjin30SFl46QBf4ba/22z3jUWm/070OJ587hY
GzzL9zDRBoOrUw2loCUEot3XAilnhYgUU8quYy0PB+T1yC4Ot95ZDVGzaa6ovs9C
d9RUj4iyvH7MxmyiVz5CxvNRGi/odHMY9/V8KBNHLjI9Z9Sc1Cj9uOZCp4ElFQCY
W/7UWD4pZPtw9j6LoD/neI/ZCg694UXFrdLvLA+Jcb3VXTqdi/zbdwKRPxP23mxC
bGSSfj6PGGDHOtcPKlOEQcqc9eX87sg9efLl7CAjBG2YwKbnUO84mHSnoUrE45gI
nmMWniFmbNh+nn4Ygu6XekJaJhd3GsDcHJpQ4446Yk11p6ggI2OB5XRjTe3qdvx+
WN9m0Qacnuwg4LVTsTWnslaNnYH1UdrFBljXeU4XKKcLsH4yM/k6trfAZRkXniLw
9Sygr0GX9Ch4/OHvUvivSWtgbcGDWfhcI8WmQ1ZQwezYX9yaAo/gPGTMlNOHAwEI
WesGzoCXi6ZmFr5idgeks7Pa9WiA3ANv+/obqYLcjkYrCZSLTOBTjf6Ps/a6cZdS
PdydwMxEpEKn3sX848oiVFOy0z2QRktqWUpxNJerzeah8JLlJkulE3TiKQrkMisW
tF5BRqbLd69yhexa13ic0N2qL5XDF3RqIr3zTgFC8H+i/ecjglvGlGQNZitJlOCE
JTwUJwgQGgRh3LQMZtibM88H1kCLp9ucGg5WEWA6KUh1jxQpnW89v4teX7AiOiKs
hloxaEpzPzLnuDVcsWmMmgm7Zl/lsKya7j+gavOegrFE7FwikMSXABwtf7qV/6gx
7BiK3WBgVGIa8W+F7b4fx7ApOoH26ueddjJBwvxvfSKtDwvaig8XJEN+dRI4TFKD
byw/8ujigfQUAq+PfzA0/Xeobkw6GsbFVsoGHW6Aktp+TW6AXnG1rQ4cqGnYxwX9
BmkQK9hBy/LLS5pyx/990OCmroCWsQBr4U2e2hwWLAHvqUS4Qo3Dw+GmbyFjsf0N
Jxa06KV/wt3YEb3zmU5G222ztbUJhaJ61EvG2r1vJZrOMMfI9YqudWKuBsgJQVri
PtM4IqtugMoim6oBWzvXCusnpXvv3Kg02hOxXXrrmQaAH2/ZyAKrGLXlXDScjED3
A0ixCWpGPe5aTEWoVn+EJ4y5pFVIHuKXjXWnMEe0HDxntVnsXY7YE6a86KDhy60C
viO8DBdTPUfP/Pw8BIYyIPhjMy7QwkPbVYGnUMFG3bOo6R/lvLiSC+wIlZgvvHG2
M1647X/+UitNfCsmh2sQYsG3nVngpqACPPpgrlz4/F198TOafrs3GQA6hGbR75GE
NzPcQQZze2DSEFxnDriHE60vRaUhYOjfiD3721DV0hmH8seY/J2EV0GHjvsTkIH5
yGxn2HLLURkBcxE+oIETxMNletDH1XS4Grb2erUuIMZoHd090SHUDEAcnZEicB5k
u4Da/pTNraSAuKGI6rxFWgJdKBzx9fBCAPMweVL7BzRKnZnj2jmJ29m/gjcry+Lf
DdPX7DVZu1aPIrNgPDHiGw7xS40Qd4ydweYfDqYa7//D+rKWu6/zT3skD2UJ51g8
Kw+AHwDH2Eqi3+SwN53XBPzVv4IgdVvqjnQ7ExSoTQDgwNw0EVrKj4XJWIPmeHj1
0jlVy3F7Jjb3K0rAFztsA3XY5/1q8Jrp8HXCcm6oXDvBSpDZcJSmeghkKFn+oe7Q
xuKm8jULHr9apnLjfsZAvch3ckARSPEXrr8DP06lt9o8u1fGyFoKc2JK43HqEhD4
+XwXNVtyEvnO+phIlbOf7OE01Ft+Dn+NnKChD0w3Am2oGvLAtPGx1CxZni+kdL3X
zLHw8rhC9c9h8qq4ZmuZnvMLAzkTGKgCuZH49GgVgXyEbf5V+qC/VmgulDsjt1AN
OmkrSQIT6zNchk4/Ssm9hP4Sq93KuaV5Z2HOwWIG2UwRfBJtK4OHGiMo5HIxkGvm
0ukQzAMmxkcodIFkQJJkdWGF6Ekt0LEpuoPejaYiOGE1tUPygToDbDoyUWgNWcN3
8NE77w1zuKirj3u6SO3Kapo9gSaei39mRY2CwwNJ92ndV3v8MAXaiYYAdWlF8nLb
WgPQ1UPPJMKSOcqYykeE4UKQCpbS58LoyCXXjQq6Bs/L6PTwa3oCKvWVrYIopAhb
lx2Od0HrhZZzBpKtg9idBhIeyrb5Q6ZV+4X1OY4Mi9B/mPirwIaN0+lAYYsl8+K2
fyhZS+HsgLERt5e1IdNOmRd83+bueNdYm/xJSGcuXPh/cQRe4C9DemsQ5Z0CSE1/
4UP7f8K0GCdTl2JUda9H8pTVItynQ66oPsHs1D8y18Ja5X/3xxTpxAmAtDRqgpmg
hUJZw0CekDpE6H29ih+9hz9qVl60K4ctrzZ+sGegaZUeo+8gte7u9ZjFFw1wS5PE
+4mAFmlseMRp1ZuopgDEfTUNz+QnbUx7QcAEi7BVNAJC+5X2KTl2TBZ/61gR/XBk
8r5IA8CSJi4lm60s+0moVitjI3aYUNELV1TdBQ2Gt4JeL0WJSfrDH8irdiHL6vjz
P6qSivRisTgxJjr+G5GlsZ/FgBxcoWdd/hKyxlsDTMovvvxqynnWgNpCAnPxdOLe
eDgbzLY78viseUNgjqq0rZHSMXtbVQv71zS82bglAQxXOQylK2j9O3b9aDo7adfP
ULeka9A3kfOE2LfxyfT7VO6FjmBGbpAleULrrgHu1ympWwx5LOyAJL2rPwLoLxU6
umjfCPAzlM/vd34QvtK/FL6YUwJywsr0DbOn3ssmDmz0qxBKX6KGhqu0Yz0QD+L+
zhC+NVej+RW5rAgWSTevmQsoWrL3wpre2ENixZTTnROW86ftOkHix0Qi8teAPmIN
PiA+mLxyb8xP83NmnY0OnGSyay1UEOb9kjlyqfPWxg0XpZHvgwYWjg5BqZM8oDZH
7NcuVGkGE+8KLBuQezAWGEOxGSKiUbp+zhg8D6SEkh3C6ZAWfOkw7CexGwRjElkn
tg4idS0LOqObNAsXJt3NUHicwBs8x+YlCzr+VeWkZ+NNzmoqH4ExxWItvEwYEsPB
B46Pcev43Y07Q277jbYgnXRpnN2m9IcsMb+2qxC0JXue7IXUOI/G6lbOQwVISPug
PNESULJH+s2oLFc+5bS47nW10unuySdeE/+TJFWgAo3FcCSEmV3fwsnv30bT1z44
6DclgvfAt01agQQ17jx0To+5a4sxQORTbfIqrEL/wwrGcU41EPDNPgWHfauoS3kK
gc7AwHe48LqQbH1VfCDYbTv71+CbUk0LtXgIten2oaBbPbXWEeSLUHRj3trtvZvR
rHskey4RFqsAPBC2EYAPOsuYey2Yu0W+7Gu8gr6P6IL4ke4PUvv756yvQPlNMaLH
5MxzWEnddpi71UgfjVaJ1KR18nleIhmZ2BOS6e8/YoVon75YZG/tAMRxCTU5ecQt
DJlXJF+QLLjKNc0NB317aoj8dSoxr02DyHUsEs276CC+j1DxR9BXQ7529MiS3s//
9GOVWh/+qT4FaaxVtbibrTjcON7XU4AgNfafJttsmYryHjbWjUJN6PYqQryGZnfA
R23KqAqvhF8q03KikEBtRxEPcravmPOtQbWD7KmAbgn9ygzs11ar6/F3At0OQ7hu
XnYWxz53gvGwvQSywF8+qn+Tr2bhwMRSGxIXi30KQocl9RrdPEaG1gMLA4YxoRzm
grTsDEMNcrb1L/zZsVRO4GGPaVvQGoJGM9Eh84V1VytuyJ7flFZpLOIKQEHHPlsj
svLyChnxSd8y6blvj+DGhdABjy04POoDocrDHBsAOD5UEcTTyy/Vnouwx+mtPf7u
0sIDv4ARG1mKH6lbkshONpz+vr7M49coUbW11HlRZWOvIrIg8Rek30e64vN7cTMM
+X9XhoMnzjpirfIai0vD3fRpEeBWprfk+8lYsKc4L7emXinoJ7P0kj/PoulApHwV
kk5aD2I6RkbDqC8juqJ+UMlfLVkT1Oy6xAwuSSGLXKUaFzmvrRYDddN1/uOeFMd9
gTLxbfV0cz232Cemoy5kJXsT6QERiDJogxXduA/4+CdBEqCM5/03CqJrqHwPCqPc
uNoTtRt7AmdpET7Fbhl5ifNsBb+X5mUg7XHzOiqKUa7qZPLIkIDNHp9e24PACtLT
Iv4Lmy86AVCIoeKb2xF7vmlFjV0c4V1mMtz1R9AECiTCL2PzCmTx2YRFsQbPPrtH
+SDYdfl9poyc8Y7976IL5juWr4I8NGmi4eCNYbcOC+mWT7dORl3YaELEsCTYAQmS
n4anrsvzESn++1+4FJzom1tr89T33wxsSau2Jnrnjv62VaqBnXZ2RSF5dyiOKYAL
5PdqUGC6J11gWGnunim5KPNHRq0RcclZMmtofb0EtnrTuOl+k8gLjtOawafRUJm4
ZUIDlTYvd2as02LHVpF7R36joeqqcOwCgrkKUvpn/+RDzroBG24SofOFV64b5vfd
vb3KM1oEyxrmm5qcYrqzpGiTFveq4LjNx6pFnxcreZ+C+FcKfyNLoJVwbyJfYKkY
/s3ojfuf1/TKqjqWoZNLAmulUIp1UwZwgPtM23IvMfIkIEEKpbvLiSK5Ds324vvY
mrxJW/4xnb4mcTJOl0Olgw3119UfbitC5euwU9ba+5E/pdlu3PU+4ZdTwVIvxwTG
A/CsKuzgkzimCGSU2RiuR/+k5pqo3cM719BgtodZRvgf8yd7pP76Savpg3VBHfKd
AB/AKH+fKveTd+6zLmLzCH9Arn32VjpWXUDWvQ1H6IWs4N0jR5t3l7Xc/fE91XFq
LXjEAMCs7kkJ3miRRHCn1RgXbSekIU06rqzW1rIrk3Tq6cHenIk6DHu/udl9p2On
TjaSyHAOLZcF0BAwVRXozVDj/nbbDBeLsJ+N24yIgPo9IudgnpYqsnLTDH/rJlsn
tFdEyeHThZqLaCNL/l2sLRoKSwGQzCxsg1EXlyYatGON0MwwVkDrKKR9xkN7XMhe
Gwut6R9mYUdm1e69EX2vO71FhEmr4/sVNN8rrxXuDun7vrjRMGREaEWgs5X2E2lh
iQ2XnMv8GKhNiieoGtuf07f4sMMszC8kBV/n7YIdc3pq0Br+GtYu92esex1jSrcM
asuTUKym2E9TE5Y0ayW6vJqj2pvH7hJ4q1kUmAzk+nxkPtG5gQhxFGbm7Lo+c1YL
PK65JfTn9rM9e4CJrkkFsvYMSN2mwOHGaxdmTNuc9rUBWXEgGbrBUrWiDIVykTrz
2w6dkvFcrZk5fphM2cpTTtkDHble1HcjX2k0wVTOWG3/XSzxFqiezAMS+zDgG1VL
UiYDtk5lAh2Tgi6JZ6Y6o2co906Tz1ZnWcUlDwyZ/txt0N1g0uhv84i8iFeN+A6p
9+s1UJ4i3WFbsAd2A8uaPmchRxTpUmWARyKB/ocZPhYbaW7vc0Ea9TwVYTYXtor/
gsjq8L3aJ1LMU0yJN1V05jA5Xdz7Ls7SWNXr8RC4EcOB6xD7Mct29EzA46wjVKi3
luGFnrttKCj/f4JXdt5FKFjbcJw5mMD8pYlceJnhUt/y7FlsNykFLpi/bqTs4sDK
12bUnBet+vN3HtCe1eM2nzCcWQpJ7zvFffyCciNUZ1/MxZ+Zej69B3jkwcbb67aO
3oO5hOfQaeTtB2c4zKNYGr+QoHeSelr+jMLF02NqeFGtaBDMdJwAxFxWc4G77NyV
+1FlHML76gUiveWMHRIlwY9emSGd9tfYkDW4YCdm3dN/WQHamUWRj3OZm7V7WjRb
4sv612ljBjVcnBO8TvkGb1IECc7uwYz0ddfBbm2mHW8mRgPnIP6xppZTZY/gNdGR
r1ZzGFkruIIMKR7je0sMpv0yPFH2VEbxtRxqzqKqMuM0OCpbvxV5U/S1qr9nLm+y
0wBy7NuSPmonSd42QyyWjqSD0OAUtIrZluukKKUXw4dbYgpJDqOnMh3jIsJfmc4E
3yZUz585fy5pSV0e/OTG49z9pulw0XAhjXiZ1qmXQhHz0QU6xmVpXmnz6FgXsvFQ
ryFvlpSmOGjnHkChlArpPqUhc8MXu7y+/UiFeWX5jGpXNgnIKjH+fnx9Vfr4Q7XX
5j5rHoNRmiRKaO5HwBMtKdbHLVMjN2CebNH5ay3d8PUGcMDMxJ53S4eqDFex/BQN
kzU8pBYu7zoMqv6k/zfVCNyuKOFvkiHjwyaiEJDXKDBKUJjQRpaM7bAi4IgeVjlu
0A59MdhrZfb19L+YQlmz+pUT5NwlM5DaWHrxcQfNJ5VAXIVtvgnE/FIUXaEsvulX
Lfc3BDxDrBppWz0ZQ/q89ifBfi1xWHGIOhQgEGBEM8YXM/TijU7hU1nTEnU38WvK
LyjKbVzNf7f0QIQHr4fP+rFfZINn/7kpkP94t+wgFCGbXKfXcu3NSerF5VDZtiVi
UDkpKFAJzkvoJbhkXRzZYyw594bzJZVutnMulyluh66EkAoeYYT/bO5lYKxJjD93
IFMOBOQ4gWpt7FDqm6Li5ZR5wz8utoZ4h6Q3R1xu27F622Ta4JqcyCXBImRRPwSl
qh1CDQLZD37eUE4KLO+a+KtbWSoT6wJ6mpR5/GP4v2YgLTJQOAdqfMAgyG+02D/v
r//5sJCNScjDIe1eKd0fjfErEjpg5ONKflU9FoIMlTBjEzt0GAtGFvqrDSRasJ9L
jpcXBj5P5rKBIQSrX8mNGnM/lg4Im0qFlX1LY3O/vJS61U5htyHxO89PVQUpXmzT
c1B6usyksfx3Gb4+G2zHsDpU/a3F1i/GI25SCdU7JQ0p3+SUntSXyXWkKjsjfncA
UWBF1RbGbn2aO44lmp7KtxZDXOXw/1APRAf5f4VbOe1P1Z/f/A1seg5bHnlpNOwz
CeU/ukl0fuzNrGoUwOWhBxXWxNlP9wqHYyyphH6uUTBuQFm1gQW8RuZLc+yIycOR
vacvw13o0jgjkIjr9DFbzigAEFFXG7doBH7oeGGHyfXdGaBBv5Imv23OgV0YHcsG
BThGoIT16OlKNVRwJFUJL74g9wUU478vb598YBNaPqJV9WME6+Hhb70cmeuxKY26
6TnK6O4rOgutzDU8UmQGKWVEHB4E5U+il6EuaeVIutbris2VhRVvdNk3KieanH+J
Iqvnj/rzrpe5o8u8Jr7QzayHyn0ivNMLzEOQnHLzqRHUvkcACzCekTUwZrrwDonZ
afvVyr1CsAdRdjuHxFsvnN29FLRwRecsLdlMpbAwxccW1EFakHmkaq8Rd93kaT2Z
dsYmeofrg6gZ/yxEfpHGqDPZ06c6sPM8+4f9NpdTEKZCrPXRTGxnKTLC2J7jwLv5
mnzKsKhn5bu0HTVO8NnE2CPc+NpUIPU6Ruck1EEDPeEat1o1YLJ8lsUshEPOg6hK
91zG7WzJUH3OhSVyof/WDECL/Zje9ZrXCI2HOjP1a6KFSJnUzdISSV1hkVEaz9SY
+Se9DGWPN4EwNUHyEGKLeEeVCE7Iwa+fjfbBcUlXBuFpUeODUyWNXIT4uBdp6O+U
cPiw1tu1xk7ejJpRnOT8+iD3nUp1EIdK3VLNr3a6Cse+dw55/zlVRu78XjCosGEu
qZRnO7YFI40OQ+w/ILLCqrJXPy1xG0l0+OkH9PPSTzGm29tQnvxVikGppEJAv7Kp
ceR8N7he2edJUqd5jp8/dv2RjMMLeANjZLnKCrNS41srLeh8xqITw3sJMj5mUU0B
LNQG+Kz83g2Kd0ukegjlGZB5f11hWbKZlTaMN1D1J4+6CTBV62R84DBK7FBRECdc
3Gajmye4J5bFJdRX1Fbqcgk7Hr0NQ2n4knyA1uvyGHze69zp9+HF64PtoSHsgaFE
k4fqHT7K6m3aE8KBKnlrSKO8ncmg46u4UlNmJjDT8CECIDBKiQdKWA57mprYKT2u
O38j4hVvQ0po51kBOqJXnWnx8zlQfCNUrRTxANalIxw9JkGC99HxhFm9jfAGgk8o
+N3K+/c3fVcnDES9cet5KoQUgVOsyVZ/1WpKwNVIwcfPEfwN+rQHF0Gctq2Vjj4W
L5+PaMRz1ymu3OYDde5CcSst47krF+ISmRn+Efyo+kdhpNI1XmXonwFGrXDSVFya
FjlHveperZcfpsPMv6qtKzDf3orpSaTcLqPmAQSBdQ7orWsPUAS01f3FLcIaGwvE
/an5EWT53t4rIhK/uOrX1oj7uvnHfFN8hC/pDQpFQHydFsVK/92axJGEvAI9BdKt
EPYiVgybi//dNQTiRvoRhM3a9P9Yct2bzEKk55evAqZH9a7S+z5IKTk0n6tlnNFJ
qHHzx9c//BKuJEkvDK8N5UyWm1hPdPwAT54fNFz9V74oCGeziGvs95e1lgyy4GjV
PlR9M1mZ1DdlGDKWYIqN28yNKnGn/HM5YKBZdemgP4gOqUoYxuhjH4zEgkh0W4n9
4smtHF74w4Rf4XO6ceFzec66GsNtighYs9gGQeWZVn+Fl5zEErmrmd59fHUY9Tzi
hfkd8DqtC46FDf0URCLnqFzb1JIHEQYS0RT35jaMbZGqjesyE2JheUa/JC2UnXJv
OWZSd7EF6jPLhVcmOvR4yfd9n+Djfcon9ayJ5vcjNPjkhddptoQWIbVQNYM9OhWC
j+dlQ/GC6+A/THgiDC0YcpfsV/je40HVQAQw5BlmAgFcnGSy6tLHh/6DStfto5rp
gfdQxOvAlSXKgQnIEpzR9zSihOnf4lF8d28xzsEK42E0z4HWlrbqyk5/aaFXagPe
2/5aUjX6wUGUsrS+dL3wT9Ta/RxpeOpBLJYZZfx0Bm3hHU8cQIj9Oq3hhUS6rAPB
GUBdyA85oxyp8IZ9XsxT/zJMAqfokvf38vOZ9j0ykzkjFVywYfqKwQW2AUIzC5l5
UhyAEx+AzS0m6lercVEwqiOcvHhYqUZA+N64zXeaP6nd5o74A82d9Yq+lFbAaOgJ
FcmYjWAz55LM+BsaZZ67yPHSaxKOLRSWHbGM5bcNULYKxZ4crJwazeDDyoMqgs/H
Xt93P8w1tbNYYvXpP/eT7ndwEYsmLqbrGLSbm+Tcsm1h58X59fyTc5nJ1ydgmuKm
jMwj399cJHq1Nuae3uncBXirptHF4Z3quRRafVqX32ZiyWCnyYKTUmt7wJSyC4Lw
DyV+21ETWDo99ly+/ddjL0kJ/ESYb/5PTMXIHGxEKELpNs3mXbTUrc0Hr2kJRpce
C9rCAGj3G4DCb/4uRhQZ7VjrJozl5VJC9N7scCRU12gz9qAVUaT0bGFQobDcHQ4s
oWEYVz1PDYYmvleIbaMC+hBBJuxX1PKygSSxNlMNYmxm9ZTYNeyNyIjQ53BwygQ+
80CVGXzayDoYIKv8lmhE2c06u8dUdkH2Dks8SM9iKMYaFq42vQE62d3cqYusEAvu
Fk42UaMmqcr55Oq5Aa7EO6qe/QwCI16w9z271+JJnvpUhBlK116iLoGXYGZHl+yH
+SfWrMrx9kvym/CwLxUlAvyEl85bpLW4NOD2C+yxZYzMb6/2CuZ5KyAtCBwjLQf7
mxK5/T9097yOtbkhzr5u96K8VHgACf1qzkpQFz5/tqDB91ezgHEU7AKU1DUDqgbd
Lo6BcNTVxops7prFDq/TW0ojXHJ0scqJaCV+1w5s73viGdxyIAoWG+d0ZoV+mq1W
wCXhMdC+DbiTka2H4Hzv/RgiYr7pNEzuCg5iuT49cdzV0ugUVKmtT/SnrobDEzac
l+WBXEHhbaturbIPq+YqPLdTyeS/MskiSfo9LTo0bXfyzPTAnxVIszfFd7m4PKPU
fbxpODwTC1WraaRqm2WrSSL3VDZe+p/8CivmxCB4qo4GxX/s8m2yNwIGxjX90jYl
UB2S3+UnvahvPdM5q0Yd8yqli5PEwMFoRX5k98iFlhxHUCBqQ6O4ywam2vYce8w0
vYQVDuQQTGpeuGl0A+5LIPM0a7C2ZTzdLayCqYe/RNLvNgD+i2GYBvh74hzgL7pX
S25b89K6EQWvUKeH8Yt9ExVEJ5a0PMTmD1N86OjNvjrLZfmaTmCCGFkBOu2qdGet
JAw8fOGuHvPZZ6QQkTMpBfjo0+GYECeud8Ldoec2yHLuad8U79FFCnt+KHiTAbXh
SAEE5l61pDegNGXHbgWWHii8Fz5clDLreBscQk6577lk6HN3vdtnwOXDxI9n+6wW
6zwR+GokkNKCb5Nd3YYGoCAw7kVQmuRnWQ4S2uVmQbFILXleYrVBaUHSN4nsOlH6
BFqOOCHZ/nsR52+IzAn7QAmAFqsQDe3RmNjw1WgKv57JJ7wqv5eKoaGf3WuAKm7N
CvVNRsg6QBxp0twXbYDk10EOPG2tcybQXSsjpn1jyLDp1eY/iBMuG+Pr0PoV8l0w
15+V0ljf1/pBAgjV1qmtuB/b5vCeYPc4tZqlQZ7k/Fz0AcNaZDw6puYXfrb28kWo
XhvJbPD56mUF8ZQYO7bwVIm9dIRE/k1+edCVev82ewrndWh3uWaJLoAqWBLGlBYn
ZMVtbRw1+jeBKRJM4wL04G//lGXfvvi5uzuyPoeMhg0W+tzo6xDmPn0N1vVWdALB
SFyx2oSYkXNeO++yo75unE5UtouUYKBLydQWypxNd195DJjwh/CDyhjQe5QZ8zk+
Ej8BD1m7+7dfx2JTetZSFjeiO0VBB94SLoejAwBxcQNhJRp6U0tB7e/Yz6wvIm7S
kHd9IOCXmRfOt3+AUxqAXlW0xexDABmu06FckdvgsDqVQ3l6BJSYsPIP41ePZdOO
0G7MA72kM3ds9niQamNgQ3RuJrwQVdMzDyZPak/FWVW/ftr3T5RvbZR8RQYkMdU8
5vnZvdMzuFecgGajm4C9Ol93YnZIOx1NTDFkNpLv72N1BHfDTIyEPKE4caUwZlW4
ZRKppaLCbALMEKaM0qgf0mQKgENDfFhLTbWH3Db1LpMzN2p0dt2Yf5L7DUYT4bXc
yhc96r15TWHOzLDy1SDnLiam9pfBmH84Er4vBJR/9LVP/uMjmNpf/2+DvqOkPsKK
4uDdLNcD70RMbNH0WmdDEBgvcNy3dxr10ZprfHZ2V35LoB9SKfo6pjod5yIfY5KH
hZ4GqUYUxYxHCnPDP1fPQeEzvC6VluAp8q1kjBs38iEOnqBk+n9ZpXAt9FbRR4d4
TMRWHAYhdbm4qAtNdQHX3M2pXreNjA329/6MxWkquIqbm3o/vjA5Be6WN+il1Q+o
95sL2PY5t7pxjwhDA/1a3zqFwReLbYGUWbRvPQK2rmaHNO6G2KYHbPY/xsAYXBe5
YQ5lduRKwwTpCT/2U8GYWCY2/wG0f298znNn9+wUaFTOcd4yYXCcrdvprjXf35OV
10Bc5+WJo9fSmJfFte/kFq2bW/PgLfhQ3yDX2GU5ETD8RQqpdAmIubpFdYFC7v5d
0cAidcHBMVcGpZcZdk/ZitvjIyOlR7AXsdtuDMts710MrQFRE+aDRLgXEUxonPNZ
XMmpCDb9LS4nM83TjDOGEqFK5FHJsIpTopohprl6GaUyA546rDFoimuCs3Ld1Q23
sYQfDyEk1bU+DqQar4ZNPzifmGbIplqx0EAskpERsqSwQMQWbTm8yRybMChJ70H0
xLiathshIXPmRWwUamAajTWA4NRv65WxbO1TSyfi+CZVHVjPIhBjqRlCBCOiLG2G
Nh/xV0cEoJtG5EWgs912WEBzqLrwFEaVRDTk3n4OwUHTl78K2jMuUywwjrcuQppQ
XZLC7bCv0liEO0KsBrSAv5OYVR5EzPC2JDpXXXnFQAZ6OLdTv2rRiKqQHADZxJsJ
JDpMwoUbVufnCHTs15z0tgbXQgEyYYDYCGJ6svAP2ra+iZ/O2B/zuS/cjwFK73H6
A+mUJ23Ri44Ye+iaWW4jx3a0YRrgVgL0POBjs2NRMrLMo/ClwYTYUcyyJECQCogp
Pg8CWead/elZJByn1qmWs78+qYkGmMxUFhHvXcANpc6P9wMak0Qsj3NI5TEcGGCH
0Qa7JcXpxAjdh4CvseyiQEeoNVJZEP01P4NuHcnsWGmrAlZIAlvyJS0AYDwHzv8M
I66sEFRp0X4XyI+h1G/hRbwUYy7nz31mt3tj0AFu/EbmxVjJUtqCF5jCOtG4Vl3b
x2+nA382B64F75KT/gSTjMfIWDhjuqOqsxZSSm5XmyjYzhlx5QrWy7NvWKe063NK
unnSl3wemV+xzpYQoFNH2A6oSJRsYY3q01D3k/PIdtIaXvtsG02+A8paierV1I+H
3/Py6lnA7jkNZcsquupAXQIquGLqI8Ldbl4hsH3jTc7oxxzXQXwTjSkjxvD4NSJk
Ndl+BPkwun/W2foQSEr/yFJAJ6YC5iF3Fgtr6BV4ykDrLwi5uspEh0VoYZeuDx8g
t8BJBK8K7D749SKprUsqavusr5LmX3r13tiVw0fC01HeJKZ30HB0IK0Ve2NSL2mb
z9AVyJY/kg23mg+kBzMkEmJ/Fow26AsJ892GN1QGpCdknusxrtQpNL/dRL7wYX7f
wRSkp95t+wsU0PR4cAycI3oFIriB53kPay/RZaITb9UW3jbQo9eFVNJIRYOZi3+f
BYNIZPFp6dt4ywixNXt38TsoSVJ+831rBbSW7Nsc8v6q3D9ssaNWnH+qJp7a0fBj
qdtsfjFvRofqPHWXCxu4HPWZ789qRYejUMiUlwTV5n+u7+Kj9sq5rh6CJH4Xsbkn
0AsOhCwgoGGQyrR+eKMziQKyOOXHh4tc3kxc32ybm4zdPxnNJQ5k6qEhm8g53AxD
eG+f5VpB/E+SmtYwuDr1lN/1S5gMduu9bCYg7MaU/xjVE4ws+uN1oA4X3F1aYSfz
xxpCvs1xwKV5kU93VVJKffAmhaK+dbZP1HhRIWTAtZ4HXUkauRcmyKdIKAjyeYur
RbTncBvbY7DJDRGLgxW2JUtrfKzI6htCwtau96XngQCYl6e+TUzJnXgBT07VwWEF
R6GYEAnYg2qHLPdu8smdfsqk5KSDwb4hLhrW3dlu24fxB+msKtQqFYl6hanFwo1K
K40aFsBTU0xxI4+CpwN2mgyH6qzH78b3hgjNCJw9bLCpSV8HC4hmQq17I/Adl+EY
zQ5LacgoP37jJiqyvNRbDmpEkAvyqgpjrC44VqKpahhqyQYEvJDFwvDbXVHpe88C
UY96UEUV4FE2qoYz3iF9TOJzE1iWOw5/6Iy6foJPkUWAShPxqG6viHuH9P2ZpG24
kQTE4Qt6+QJkbIiGcYYIoTGgW7y1xm09igdXFvCA82k6EcrlWbHWF2JKrBbCBMtU
tOJA92EAvEPNvBVO4XfP3mNaWD3Fus5S9IKZ5/AL0GIbyO2CP0QeFzQq016WV4pR
rQbE5Gj6NkPJV67sFdZHTKFCTQkdIzZWJYbG2no0/++yJaykwoRXFFjD7pVWOeiv
5f+sWSEWqUEgxDXdfFmKISJ9Se4q34oi1nl/Yij9U5ZogYMhjP+YN691ZinL0Y7G
OVC5UCfgUVwt2Y2lEmDXbJFenGb2D0ltlzJ4jkGau5YTRUrHRVROOh7r0KQdasKC
nM443jgGX/KwaUsO3u+iqYRfT/e8TzjpAyXi7+Yz62NaT9FBHVaoayNP136VU6QW
qXK323UcLleV6AMC+n5mi6GUhplVp5l7kKPhCU0GJk5TUFEeUhJcqSNEEvO8q+SI
h+JWG6WJgk6lDc9O3pagVaxsHvBuvjft1KjfVQS22PqUa01qS/W4lLP0pjtMbg5X
RTRJabYarv/vTeFRPeCroIE4Oh+OpzHSvWtDIPTzFAhziCrVxv7Is0V85CBDbTEk
KSZ1W371hlDn0SnF4PBe+5mBMc8Tq9Vn+Li5QUlqg/VzJ9kWyGZrhdCxQPFXYV1D
xPJY8y3rXtSvy6aEH/Gr8tcT+Dq+9ShRtN5olDI+Zm6QKyV4F/u61w6nq6uUEsGa
kyf+aHowAzuZsOxAfgLMoDswn096Q4G3ctObgD9miE+ZiqRSB1nLWxqIWcwUsEJV
vpQOLTunUnxsTLCf/OH1xIB23dxV8XYK9jMV/etZd328VbaDXWU7HcNlXIojd5K1
F4LKEk1wRw3O04QKVJ6cyb+MkD2QBDbPyc3UhhiF4v4P4B9bhjDusBM0+avUAImY
HMw4BmKWgTMHUgV1WP5TzyB2UnGxc00DX9nx6/zo20FQacVIl4xbT9YDEvMZABkD
vyXoqNX8zMbmm4iIkvAySCdH9NTaWKGwWUIEv7mzW7HYPjUq+mtJfYoM5ZhFFX9x
DziQAgXknde7p3zdkaCUa4pOdOHlmacLMsZ+myXK3skX22Wf1F50skG7eiGfu4G9
6XQd7mKC7UgQGkfNawY7K9Nr5P+QyRtElbJ0l78MOG3xn0c1oU4w4jZkF6Dz0uar
PSXwJAZ/qW/+0yfa55redTTwqZztp7XskS/e1ULebYYA9+5sKsg1WDN5XNw9ia+f
g+cE5uYZNOboHIl02LjOD4P+9A9rn5V7RUrV7wAAHJP9Xsb3OoxMSzoSP5InIJ8b
Jp3OWR/jE4dR60evNtlg73LNvDotjAPtGBBj1yXLivg56iJHYPIf5dUyrj1S6OtD
5WqRT22TIrawzbgeRsRHI3GI6uzD7SUiDiaYNTz5lAazzFNyOyfSYKVBiAx4XeWl
vY8ag5af5BuPSL//EVjgqn8t04dm/RbIYsFNLQMBcCVuskUxZfD1MROq+AaRvDyB
R9nMWlllqq891i9fXWb6Hg+zL7qRgBSmIGDnStRbGvVtoQy+ZVLE/fJor+/oxnWa
8AfF5AOOl02SDs1Nfmeob3Sb9Qvw+6y9IqvsnOYO86wlmaGmoQAic28gwwwbqy7c
W/O/s7VLP9fg443MnwBpM4Zkp8D3TvqQfWaP7QRnLEY3HQ8ovDeWYkM0GUc45tY4
QUr37mBOxCN1+c3Kn8eZtQYGb2Atx4Jsl9CT0EWFnz32n7Yajypplkl+WYFeFyQl
WdeFTnBF1RrSVGyrz6STkMnZXees12aMFMIMY1OAHSZ+5RL8DMWirTNYhUlOikGB
lSvnKWltNnf6XRUnKKugjVq6f2trrbHZQnP/kcatl1lnPCb6WMvaEZzSwlcmK+s8
/rZPwZLQQO+WYtrf+ixL8MvR7/iF4T6/VCFZ+tni2GO7/OAw2pIeHISN4k5Sr5IO
j70JDf7/I9SJMN7u2ekLes6XZICPSl+Kxj1362F+nKASJwm+Fl3CPoN5Y5f2SSmJ
GAMYH65pvRdydRanoXpFqnMIvQdwWU7k/oop2PXSYKlLzChiHGlLUN94jsUGUmfs
kGCvQ5RglsAX/o1LY1pylSZOXpaxNFqwgwwXHRvOK66Gal75U3JbV3cSCXehb5Hy
xnajJRuOALBLlC5Vfn48mkHLmxN+1TdUCxvtivQBLFkS2fAS4m/qG5htMhOSu0AG
hkIvQpXi0iUMPvuUqbERhHOQDRdO8pBCsRG6x3JdtN2CYoNxMo53lFuaIOIifkvB
uqxpaUj9WSuXmSXHBd2rVSlaRa/SJAS/omaJ/7dIp+ZEFADJoi1te2wrrT9HirPY
QSE3DijFyjftOi1j/W4tBOhJPREQgevXbhahcnA+kQRywo/LwVjHpUrHzOnXhjCD
yWeki48cuCsH9gppuriqJS1ss8Iy6WfXRZ2nRCReL1ZcU3tYOb+75AqNLvNtgcn8
QYRVfw+tHRsTlpRvKXkR2tsAUoDj2kYeV4gXtX1LewUdayNRRbAQ5u8bdH7dcJcS
HiHeyN+Cstj7qZ9ow5LjNymVMe67FVqomNvJn9kNy2Gyc5FJhVGJPghrdrv3qVN4
6C56ikKy/kydec5aSqmS86GEQ2EjQ8CCVU5noB0UUhrXvNJ1bPAGtyXWmgIfdujz
wGq1U08FxK+7e4Z5YR3PlY++3cqbVcqjxUfOIWZKDwCHFGztqWV64RmDRUDY/Wkg
usYQ+0UfMqvrDK9yvBVLCgYBp0AdyxGTp0NdnCDPSdhReu0vDqgvFBqVnDgjBkdw
HKasDtm04wcc0ZZlC3hVKLs3GlvftFuv4hcxXBU6UbGiiGxX6j/YuFzexXqRaFZ8
ILAFYfDCzUaMaqeDA379cMFOMmMv2RNJN9dpZmWO1t6V42aOpW0Y0ZxR0M/51+MI
acFLX1pJJBiL0IktipDue7b9Ce3D6Jk6+UTZqBWvsqAt2zYs6PejsP40Qzr6UxCb
WLecYvxPYAMpDAE9iXfuvhZbn9BcAm1vFDRvMEOPGhEL1Vl3qB3cGLxA01Ke17lK
fym8VdtVDyB5o056q88SDxDZbVAKDb4QXhZiYUb+bkH8uz/AnOJdKNcyy2JaoObf
8fm0CNY1xpnlo3lNdqyROQg+vqz0IMIbMNRlrKYub4NXECFi5b/qkV5C5TaugAi7
zpcI/XzJb4Jr01SpNo4micyuIGLlboRcLAKqMYBFZCNVnnYLC9yAGExPs49te+oy
+YkRxv7Y2llf8zpdYFnyVGiDu+lnkfyek0h+eFokRoLGpJttPP78a2SHcJScpwBh
PJQ/+ztVyLVvZAmqf1s97j2ARQg4aMHtw7FnQ0AmZWXUzewC+mizY7aCqospVLm9
RX30t+cZ9PSbv/cVWEY1Q4AMuJU3SDG/awXcAmVbUmX6SAHrtdkgvs9urqSS76BD
CHysk+gw63U6sOT6VnkF86CNV9g2dQy6UvgRokCTq/09lBU9tH/dNC4JX40MAMNk
GS9FQcj83N/qdVbDXEwi9N4FBEy/hlcZJN9ZFwW9hZF/ZjAqOZSuCgOIBC/Bi5qX
WD1/MpREloSLTdaQ+cTOMlQ3aptfVviu1rjstf8YiP3Kz0n366QSkQCDh7uliH2Q
Xp9qioPo8wmgIVaIgmsU60M8q2vlvfHke3vqrOmgPkG8etKwtnAjthcgZNGVpwll
xWLMgMAncJG9/7TMTxmLXnBxDTH/1V6uJ5cB6pwSSJt15yYMjO/R7gEWlduB4Do6
gKyCJlTLfhnz5NoEd4ePwYomjzWEwSPEUoTGXqdvij85cWwPlbhreokqv2Of3q5v
/GzjQAkMw+1IPY/cJTBDKu2gGKDJpElggub8DccwIEKEOMbsmWlirIzB3M8Wf9Gp
HZ4t8bRjqwmFqqh7CUaAdf6yC7leTS0CJBu99OSVFQC48z4RoIiofboIHBjokBlY
nVXdtJOqaIcnVJDSaE92FwhNPuSFwbXrRyGTn1VMphWyaj9J/qiF4svA0MK3Q7ba
cKBSLEiIRGrFv9w6wSXeAJz3uyTOwu4q2Xd/cvFbopwiZF6TydyORdBC4u6Ol2IC
/gz0FjtbNWJYpe7hcNhomYoxXMSKyNDM2zdntSBMTHRLuHG1S3jZJvV+x0LAWxkt
Ql1KmqydqQv6PEfFOKC7Zv2+okqegrsxaVbLFA+iDF9BkgOkSoXEVAlM+4FmHAuQ
WIhdH9ew/vv2YiGYz12TziG8mP2QpB8yZqj3EgmLmescOrGWpI797Yxjl6/z9SYv
dhcx0Zxgh8aoRh7I5Ku9XXtWTwreRzrlrR4VIN2lmtr5PnAlpkx1eThoOxlgEugc
ZAG7poip6pNUneRtHRfU9UhR8er6hrDppqeyFcsBrF2BNZTUVNurgL+DMqDYHjjl
ZjRemxU82zKF/2rtHp0YL/6a/XLy/50k/qSwg1YjoXppMI8d258S+HHB6b6Zo/b2
SDV4pRVIJAtk2zDgvbThnAcFdMAiudetPJABkvgfBjY9qVj9w40vjlRi8AVMmO8p
pmXnhp3jUmo8cO0SKL95nGn0YOs/NME1UIKkSlTaa5PNQEFKoF6STiJMDB/UXapo
Tg04QMbYX3O3qa5Gj9rfQmRGINwFqa/Nm4z2TV0oObcH8VPEOfX+J2GsDcDTQylS
VnN6M18UgW8EplswHBP1zsjsWvXKhhp7liH3GpiE+hUbSMyYjd1H5USt31KMPCUM
z/J7t87Q1HaN4o5j8sRjIBTfP0P203+SHaIMiIw48pG3+RfxTaiKro9s2vc26pU3
hiANv69vgGFnom3nDln23D+h7nb2QEMvMKv4WNbDZDiMXCv/9g43+AGU75/bS738
sLGF5MQnnAMK+8sc3dHlHQY4ZnG+qB/eDXXxid5JrHe8Hqo8aW0iMQUX8eflT61O
uzb2X9tQMKPzGgGRx8kixGqC4rWGHz2n3RUbriOCF9GiUN2D6+Y3GfoqsJ2KImnD
Dr1is9fyGLXJrprQl0APdRz8uEfB7DYdjNDEFw9s9wT3YIi2W9lwfcTvDVm+UOo5
rxcqDMCR1wZpn4oRF7KbnYd+1m6ZeR/oqqFkagYmkUq0yF7kIBbFLfrG8X2QKPRE
6WxW9LcFQ9ZYkIevoTx3A2WvTVif94K9gFLXTQzrapeAn7Qy/kM/fAwxwyb5vtDh
hqlEELeBAxEi/9Kb5M97m+IHVjgoRGBi3t6l5PEzHyIQpdnd1P5ldpHBpAEuDODG
0AZiP0jX7rjWZbZot0WWxzMlnmYv0V67OS5icbHea6uPU6SmSXWA0WPn4xeSG6rc
6B3cNXsRtluXkCNkEJLu3axb8+Ymlsbl/lMld+MQoqmKR0rm2iB4qzSVPPKLbYrA
KdeJBcd3xhtJ3E5ePnzX7YIp0lJTFkHHKCCkdXcpU4CNFSM/qmJ3g97CzM/wBNiw
T6viIrdZUsbfRUBMqRiOBTlDW4RpkwMnXU+jPYpvT42Tr1inF8iU+OAkRKiSwOoj
AOf8JjRKEaqN+U7RgJnNwJ6B0UbnDycBtR8Irff2zfBEnb29QiETU9bzC0e6rfTA
q5JttCk6sKc4oWtAAwV6hXog5GKYUgtAGx0gWb2SjBAg430AUU3D6+p0MeqBoyRu
9uoPOph3pjP7iaGoNR7XXYT+hQ28IDHrX7FVNH3tKbq/P9hJitDL6nSwWnp395x9
kmwbP76XdxcCAl7ruV5SyyOCtOWyiu8yNOzciy15mBtFXA685mdy7VQvptz0eXjI
Ozvan9FNJI6r23cGXvc6mznPCNzjcoG5MF4WiHnLFPxwd9OowBoJSmhLm2hzb2rb
nJFfsDCBWoC7mgKryF/DManlIxVRRrGfyXR2AXiBOFetsEudrsQUGy7zab0+2c6X
uUJO6Bi/IVj5XbYq/LKj3/HiHmedcKtF1iG41diU2YanzCfXFRCXkC7EybARpzSD
rZ929j/V/zvCQzMMm5i7LjwAHVqNbFxI1gNfFFZs25ytpjc45QcncmupAWkr+0ry
6hSlBwEG6q2n7LpCuGLIWRn3FE/YJlOMXT2LPTSV/KFHZX5vTWgunkSSTU/hrz1P
2KgOsnh5n0M/RssdDJ9xCQHZMQog9JBS6Jlu4cr5oQtCpTMU/XzRgDNw+TJNFB77
8VJBNt2aMgl1rUDBSeML+Hn0nT25xux0gn57G5XWkVKzCy+xu1cZX8qAqZEDwSLz
7MyHzZhBISOxo5oaeH83BrijtaVqSJuoc/7L2WcyfRNlTWI6147fhckM+BwIdE5j
/wWjf54r1DCFLRcmYDM9V6nOecgZjAwElSGx+mCPBuk0fzp5bI/eJyxZ51o7gt+d
8q/HfUqkq1/miuR1FVkzu1AyAIajNQIgCUzOFkDtwfIiGRxIjis6Pg9hLYfl9cV+
ZWJKwVx5HgoZkKDJ8yiovTgNrdlJwPGowbNa+/RwovXLKuc3EBjrhJYurAkGSOt0
uVka2G6k4L1VXuXGtJ1VLGMExE39v2jFxZpseYOU9AbcCuFfm2m+EGlub7xhyszs
wIS9el2Im36litz/5wUt3n4wtYWLvuldg0S308QvwO22xClJjd1cAOPoAaXS28+I
X4jSr78a3sCRN3FZfvEVYE9+t28mL5UOgDB5HXtC1Kb7OVohQUi/CLDvMC/V96aw
kGrvWd/KTZW0uSoWn3LG7wcbZFiPQKe/MCXq78QjaD5cMf62tsP/nPiC+xxsh98Q
bdMoOQhJXQnD0iaZvTrgud25vh5A954iqCLYB1GkTBRzRTEY9FT6a6gydaWDe8yt
q3b8Wt74lKaxkwJyHkEqI/HupTs+BXkAl2k/vvoo8RabHp84WC1ePEnxbyYEc/EU
cZ+ByTsAzmLopajHjKoEMqKBV3zVNoJE/mJXsp28U++vx/fPsDmTV66kFISXwdGL
9KLOcDq4OluirhtfUh+ZVI1diWIeZ4gOHhzD5TCd4s2B89pnANxs+emjrVsg3XQB
AzOhJGLy2nBhEJiZx/xYXUbfGG+vW88Y81GUBApE8SpkISELIPf9x7HOMox1JuEx
RFJVOygNLXTH8whi0Xps0kLJE8jb/TPWvHMX+F9lSZcKPEfvmU7oJw0Cg0tXchLI
zs3+LMIl9W+CQOZO4RMQC0lECg70KQk0RuAcJ5xgJjfpSzOePhv7crjAZSQXcleE
nIaTg0ZYog0YsTxw+aykWvbV35dS0OJSNDyeivZE1hvkCCbBHBeeKbj3WPEuqFc9
zfqkZG3OuLteK0qHV0Mm/ESK+icKTLCJGQC5o3+DmKasVPLal4oFvY7tK/BtijZ3
Mmqmn8JN/7Lh+ooly6tAJjx01sf/gzWkbbvFTB/T30JwURC0GgZhIh9GRnY/0j+r
7U0e9918BVTgetpx3duT0ScM7fvsxeGlyLzHzUEvn1X9thn4K7UeMgj5sRkV9go9
9f5QiDf4ZQOJ9vRfAERtZ1WXF6dV/LzezW+zWEKA405VRVYSpZm1XQX1zFrtRBGW
gLWXXV+VdR6w4/Ee4F1tA1qNHIJU0Vfo4nMRCc5DdnDRPXBPxsBogBbKRrKwmeC7
AvZ77ce/pQ39n2vF/Hoei+D5hDUYR7+gYhItgIukz79uxxLx1BQMLYaMs5YvM65/
FPofuGSQUciddidUscJn+sjc+x5CvhfKJjmMBtmasUTFS6kwYQH/6RtzVxyj5T2F
0kSFSCTBrtAfN28H1ZJNPpEGsi3syIxJTcQ/H3EzOu5gG+93nDpou/bDi+m+5uGr
YDdNxdmjes9fm3hXWhIlqtyn/omrxbhzVYhsifT66fm+jZTvITv5RDk4DhDNBMRO
oDl0EkcJ20b8qvt0KLXQrMt3u2ksZyCjEBGhWBdVjtqjsHoh1yPnexn9CgaD6sr4
mIdUfkWDLeBc/7gkZE4zqpc7ybpvGRK9x5rZhsAl2r2lix7QF72E4LxKhQY0nQjN
XEQ5uhi79ayW+Wts+TgzOXI85ziFY/f6V/VbJaKl8SfUgVTenssFOCe7BZOrzJyS
A866teJIIR1trBEeSOgbCmsIRM27iXo1WlWMc2TZ40bobzOnSgh0P27/A2tJfWU+
yz9JhMaI7wKw7mTv85ddUYwIc14iM9MqCU1wXYjQQkBvVr4WoIGa+217l1ofdCLc
+lvCg4tMpxWlQwyUnr7H4/l/hsA7RacVQzCcmlXzSH6UTCXK+xuaKfQnxL3TmO8h
jgswmeMenYUQNf67V6DD39jjiUvaoekIGUFwIcGZK2Ig7FWi/lRiQpNF3sgsBpay
kaltbrDd120N5GfEjk8gcqY0gyTCs3WHbl0hfDMlPLSMuJSlcfmKgXvccTui3dqp
KbHmd4b4hv8c/r3IxHDgYtbAVF7bd3wp4w1+maNik8HW69B/gImQW0yoIYyKs5o9
twxnZ1/h1flpP/KyHOpwxNwZqoM0jasgWyCmGjjc+kIi+6Oxp4p88pOutoTYJuf2
KRPgu2/Rn3el/nCKXrIR4pY3FCGMNuHayOQQV7sMzngbg+0O9chnOQhGDEkTXNLW
HVoNSf80OL3zsN+KDspV8NlJ75HjqF2C84O95xwinn4R4+Tco1nSm3/kTWirah7X
q2XAWxFVGzJ/EgwyfzcU4TaiLeQ0PKkdFayhypBjXqT4kXnWgWwLxityzq8mS1rM
GB/qxSRtDdQKLpxUrPbT387UNkv9fQe3z/ph9o/UUqtV/ZogOc+gn/UPmL3tdDUw
CBfaUZyDLz7HIojtKclo1GEOPHBVPqws8GZZGpJPsEHxhn/4rGQjMkGmqs/Vbq/7
zzdAKDGCr7NqQJbQq44UNhs/j5+XvlaWZPPe7LMyE3q/88RO+wmQZeIoEjMO1Ozx
xN/rV8TlAgtE8RLz1ginDfPNVU4TRqzLkix4pXllIrSNySFUHGn10G9arxhsAdBr
32eAagBHEKUAxH3X9K4fyRKxYEazofWjVFj3I++fkOCIEm8ROMHCu/3c/2z1FYV2
NHWOeoX8sCbam+7YhnXbwMJJh5SXI6wMQ0IcLUHIpbSV4iUac01mxwH30A7gPi/K
I7chi+N1GPrHJvw1THV38gzQ812UCvju/EtRASng7OVjkOVFKT02cYAQLVgx7mnH
2zOLXqxjhcRlxdp1OkJ2bxnQHCVeRalLS3IfYC11gHSWEFx3b/5WakQzwyKF4Coh
CZz/FVlnBjHqZBGXFimVI5Vo6Fb5OWezjtbN0LqypsWaD6u9RqfbpodYoyCnkQ3X
hLx2hd0VHFhwuxEZ7dW3iLrlfmcL20putYdyTWLh/L9h80j0+U4NITqtYJdVtOic
3XxVzkvkjalcstxI5U0ODXvoGZH1n5TCXwUe6cf/I/bZWp0FgNbBL6mXrXY+cwFZ
U2IjT2Chkg1aTs8XfmoTnC33S1K6sQMEZ+1evfE0QjpUXXt1zYkdsE/Gl03w4+o+
eAlNbegosMvA1vJoPHKRZeCYKpQ3m3oOlLfR79hUIIKdwdfr8hDtE7FVfB64Q6uK
2kP90orc4IX0ttQ/6WbYzcpfM7FC6iLyrBHl09z/cot7AzjSk/myWk/2onhJBVdQ
Uo+aWPQ/7zGmAWJ/CIFoGOAWtUe8BGtErWmUIO8wAzp9i7o7RHRX1V3QcgNEVbdZ
cp+injX1KaM2nWPnRDu2HQL2ABANXttNh8aWKpwy1+fzX2724yzglouflMwjz23o
gasJepUsPwysJZpTNUpcafGXTBvtxJD5KOK3vyUWHmT8mrKYugtYCdRieX/ihePL
Ln6z4JEFFcIFYO7utn3auWHyNzIOO0PDFXiAUG7i/DEArWcGQNivnDk18Qlv0rwc
LWZ2/URlojsvx3CpSYbYadJJooV0ecBfUcctYZAE1ZHuTIejYNBhM4UYHHtONGv7
MNoKXzI76CSr1w9vEM2FVFHF3WHeVldSOFL2opT7PKfpV6Zr9c6Q3v/Ngt/tJ1uE
tq8M5rlkVIL0O4+v6/RgQucF3iR4G+/OJrLFkSdq+6WfB4HKvRSB1P87D1wOsUMD
NsPDS2QM+Nl95Um4Vl0l9s+jtgiFz+WJAwGNVTO0Bt4cGym3MOy95a+thMq8QVYa
/DIUvdO20GUfavquI+knM6OcmQfJOMY7TJQmuOmJxTC3/rVi9rroTbgoBUnVCtbW
W+todjp7z3QbSHSjOzCcB5ZBKPHgHEgoTleKInqGY1XqLIKwqYtDTYZCpF5t7jiz
gzhV+09xk0/CaWvccwd7GffBAbjJxuMHH1yTSaazbsCdE6Tcla5xooUxOG6VxKwy
Z8m3J2HpCNhe5Er9wETyhIn1togIO/nTHQTNAvpTr49P/b8wFkxtusQodfcLAXu5
1/UB0xlRcUTrM5uSNAWP9KRJuQalT8qIHtlsdfhMXs5N8vTewDXKR+h+BnnkM2M2
aupbwB4akZ7DuzGyFH6bD2FKyPKyz162s4bmI7wKfJ6woTkPgY7jpSU4++4MChwq
+bqW84NW68ozs2APvtLO+ozCF+FHi45uM02E7EO90Nix4cIWzn8/f2a+/TdPYI77
C71sGoOEfNoXkWgy6NHMeaaLYdYw90/lOLzNP0gnn8TAE8mtWVl+bFjokwNXq4cq
2BzjWGWxPhPS3gwc6u96CIp0nlMPZhWe0uBs+pqKuybSNlp8Z8Im5s7xOlZ+aKQ9
5Z0CAuFx62hSfzWWJhrGj3iktLVyFnkeyLzSDM354cCNWzqR/NycNfev1jks49DY
GRR82d02/Mg2iB3eyll29DJXfsRhTZWxp7p2Faf+wiGqzR80UOY9agl4pEtWD/K9
cpJY0seZRxVHVRK5TxDy5yDxmLWrzhwc2wvZ0Eb+dOOYZw8aTQMFbZ5Qb7kQ+/JZ
RC8T4o3nN9eHNStQiBS+/tjPKoftkC+3QRwLVKNSFHgsCdM+gE30N2lUzVN8h0Xd
HRlmRpEqcOKyDfOIwu+scf3Sk5DzHZHhhgTrNU6le8n6Y+kgmEzBFtl0uOJStcY0
PbbAlz4+tkgBD6QRumf8MZAUlbPnAwIskGNqodWs/zSAUJwNKZjm6V2y3GEd2TD8
YRkBBz5eTBUw0bJ/+h0bijjgmB0HY1dOlHXbQV4oC44/PKqd7yOG7647gIKPlp2V
LNISLZV6J+WqYH9yLAvNE5OgJNVbhwh4f1/SVjwamFRvdTBP4BW7OzBXiIIDG5xl
huOJ5cuzVEqLkh/0MqqgOeUCgXK6XDbqqof2SfNCnsm+x1ai4P6LgUL57AEuiV2k
wZJShHv3bFVBRxUV1r8+ayZQo9cu9EmU/oiBi9xad6NYp89u8lH4dJ8Mmd61IcuI
OGJq4xL7a/VdEeunZMvsExbMoWG1EEEvC63Ana0gR3PChgi1vVpVw48LVCW9FoRG
ylIoSisxWBa8P7X1SkFjEbv6rFspu9jjduWKNCDSW3sh9byR7eLhCm4IrsHo+7cQ
snuD9cGqSs8mA/sBuuRm58MyinyxjDXBy6aC6JsAUi1dWbbpmD7BuIWxhiO04rj4
uw2pKJ5Jr24cDW7mvbjQJok3FLmw1yo4y2TDQAtB+SHcydG3mSQdIf7s6qOLyRke
tDxnkwKyNyLGRfIVV2A1yr8P69kkF1CDiP0vlSJMeUiKdjADXMiTmkFzYGcVmZYH
8iHBQQ6NqG6ej9jd8y2ry8VZ7ssF+qob5jw5MNNh0roBKU6YlUEb2ePAMc0R7OID
JwYPvMOIadQEFWo6RpEcufufjtI3xkVhn7/OPj+BNoBlJmEZXDDU6a+lYaWbu7Li
B7A8qqbL2Gk7msZ/WHrBdSJczkjZR8DAuM79xS25JlE5AUOcRajXQC2p75MaV1f4
UO6/8F5KXOCooaiT4aMJ3cfeDTyF7jRUhLEYNjBpTqpHwsJfFRQDv6Ckke7INH+s
/uhKaFvQq582Jwfh8pQeNndDEuxatwumxeElaDcAKH9jWLP+xqEw4A3NAfBPsgAa
EYW5aexuRAZHR1RSnsM8fKxuA5QtBad+25b7tgg3NFV66GrjocaL9ow5r+ZBSQmM
WyNzSBwAPMOhfzojmaAq+gXUAUPZsfa3HBP3D4QeCquxduditSvaCXVfgtef+Vq3
vHiiOfhvMExTnvwdaxHf2BDtZyhvbKX9Tcoazgyl4K/0s0yWzPyG8BEbYuUB22Z/
jyvgE7EO9NIavYKaef0mi0N2hS+UQph+84Ryq7D0KtU1e409gRmqkxoywAby+/AH
lgvFQhgT0ob9wsNglN9iWpOeyL3Bh7crKrAf0ztwKepblJCdVb0zvPgawdXj55FY
tJIFQ7OJ+tYf9H6BCjvh9G/YzisRy8w4wr8iyaLGPCx8+RtWY5YrmQ+lZD3h/86r
eHJBNBtOUrDXccPkVdZHaAnYOti1ON/iDTHP+RS4W5ujxdV8v1bScwYtqqMNB47v
lus7h6OnJfYHKHYC0xqAJ3+r32qQqnfEuhKVqVGsUimDogy1NVJaas5r9rzBErJ0
4dN3WdQxHp6SxUnKm0u3beP6IHYkbcVy8KSOmnKI9LaSGnzLaujGdJLnvl8uzaOz
cPz2CfbwUzhvU+Nz8aaO/nM6kqJxmtSN5rZDlwlX+uL52FAXY0A/raG24wd1Fo0i
i9mayeAn3RHkkN25CPwdqoQNN9eG2SrLVKPdqTZGPNEveKeevFRbQXIBdKJK4Y/i
hDvKwf38HC3VJyNPL9/mCPEPRYyRXf6g4PcDINaxzR5JCaXF12jDIvAKnZkZo49D
wKeuSEJEr02f8A89UP1kGtig2dIDwQPonVzy0Q1xFuFeUDBr9/IJdjZDaQNlBZsT
yB1f9l07TMWh/JTpkufgF0GpCHFvIZPm5DSgwImHScL32EYU+aaPcJLIxq7yBLKb
Bo6rReHtTzB8bW7xci4hXZOG1FR4CRpgyjhiHvZeyO4KXWvQBsLYBnzHdxoyjepZ
CTc6r8BQZ37KpR7Z/FkT8wMiXq5eRo8wMFaiDsk/cGG+wuN4soGOGke2TDZZvpgC
fPech+3VGJ9hogOitQDR+fPKTjE0GqtEEh+CdEwiwvLdKDCtzV7SkpLAQIcBVO0F
Rc0fAW4t2bf0EewKOtqpjALBr/tvBdZTWPC9oQ3ZzY4o/4n1QkEXPlIrnyeJFYI4
T2Lu695egPSntXDhw6ly4/BIg08neiAXmHDN9gGxbMqms/fbgsCkFecZjwZ8tA+Y
m0SvLIUthgZdBlgJlj14EcIE15D5+suZzlj+m2BRPqHKsyxfvI/E0LxOiR6mbX5s
bfLE0zF682QeIaSiEgTCdZ+zVcSoX5gCVP9gyogpJX5qGy1tEIEThvr+9/5pZ5Bg
zN5JkFdEi/zz0++lapdF5zPYhqkeBMMt3mwYGKmVLbeeuT+/5h0tPNKwPS7bW2X6
s89HbPObs6jbQvEyE7P3Oqz2AJlhSVhwqHNMi5yy6hJzuFN24Y/hJP2DtlS3sDZY
zUcjpMgHsxTHhsvPN0FsP+BO1MP2dkmEHziwoFJmSnzN7dsHxWzagZJ8dHJvfXTb
H3HnM0AENhSsf/Th+aEEe4Ddmma2xvDYOApZXp5uBhTWc8axq6scRl/c0yynPM5i
IKudjzQDpF6wNPznMZmWSA3LS4DAmUt7B4FdwQttVBQIrO4MmiFEfbzxI9ymGdxR
yDOicCzSmnUsc/K8PGyZcSY7Q8sQftzUoQClU31uYnQ8rOKf22UMYpgdj5JxhFw5
oVUw8P1nltkRjw6Z5az34CcOOmb/GHIY1jVsdJHPRFX8fKt5P9Q6Eau2zRvm5guT
EJ2WZ/II385SKCVL5UuQTLSPEwcLBy9xxpb8jUkubvfy3D/ODpNHAv26JtxVJGc5
7YOi0JQ0Fr8HMTKkuUFkI9kPRTkSXdEU570h1cxQTPKAZogcQcAufBDM9rlwOq6B
Q8L2TOtSAuXwGwuebDMSORJfxQCmlFwHAz6h4N98rLkDycd8EpkE9glyKzl7EvHx
mktZZSVbVm8M+DoY1OlTDYSy62rtyaGPG24xShF0goLnDcrKf9xmocyfo222nQVI
cIW8bnQyCgo3jy+hIRjFAIY1D6SgpuKPbDm9K7VS7bKt7uAUYLL046s+SLAQ4t66
lP6WZw8XBDVGevu5yryErUI/lI4rGqy48wojd4X9yRIVBiOAredIY3YvZMIBDUkw
NCYgI8tmIT5OYWG2egW3ON1QiU0+wE+UF5hREKUPflXLHr3LUKAAQSxkg5R3yOC0
yQqKsrVZkaCw+DePbJ2p0JerXGERWI3Uf6gXj+O7V5T6H1yAq8Eqm7K/waa5F84g
QJBxMRSSWStF+HvAHjdbs5xt0FzYTRF9YcTPN1kQ9CRrMMX3fxMBgldP9rv83+2x
s7Jcv3nbYk0FGIFAVLlVcU3Ay0BgOUeksv7nZeMhF7/B9WU0pFTSMZamNwQmfegv
HvujjrqhJ8s+QXUMZWFxkDk7Zn0OFdRddPRc7Oj139aji8MxQi8uwCNQP6dI30OJ
mciugnVSDwUXZRkca3wMgoQ7eDUKcXmVGq1peG1JYcQr70t6x64g4p3d5Yu2T2/u
63gu4BCxb2c3/EUHKm+SPATrAOELjscqC2xKcLrgX53jVdlMsRnj8o2iNFuAbAk6
/D0yJNeclwMZ6/edbNl8Rn8lFSe5zsFe2sykw8QKGikZ8EzxB71mv1LhS4LmjPEb
RLQr8FdBTZDRwlwC2jlE5TkF8Qv/xUHmWMBEPsYQKnf1WZ2DdjZDKV6FKdhAxzVk
kMmEKd7Y9/3dXQUd0gKpTgljSd9gwB6jsBWfd78hFCKbIMw97VAvNoq6p01Gmp8s
zZuyDDaKiipZEt2y8b3yHxrtw8lEKuue8uGRLM9l1vJMxhc2uT6vTwdrH5czwZr0
hdRtrJIkNsU9Usz3JH4pCR+KIeNGCPK/SMwuHad5hqM1WEWD27zVfWXEwqrFhwfW
uplQsziRPaESjwOY1+AnGXdb4L7OfZe6dmgQMFh6gjoFLUXYNwyJ2qFKdCzZliWc
f6wLIJbOd7DR3smEHBwCir29qSayyf114w7e36QmE2vxWEzGG8y/d5ZfTWO0m/xa
wkfyO3Rg3vjW3bz9wYc4ixcDa/sjoT50ZI1/Rb/GXkH6OLkh2Qv2pqZACrF1Ol3a
KNWufX48Vrr9EwpNVAgqBrsIZ8rQ1lmTRLa3o/jjtdmVySqxntxKPEbPkufNhMIg
SIvl1rPz5Ss2WctCfrNp2RViZVxs+luempjwObk+AGnrq/+4ilZbsVdnzql1aPYn
fvWWXSKjbnxTOTX47V9z+f1ptVoovceb1KdKqUFnd5hQ6cbqtS0+oiuosK85I34q
C/tzt2+CMPwedQVoKqLqS4CQ8JQU06JLQhPf2dclMhTQlFcoJY3XNzk4czlrzNM3
cnoxaj3GafRCmly/eTg4uUniblC++CvS8JVZLUMSMlEbFBYH0CIKYO5+/3kq9AhH
BLtZfivTqRa3yzrmtJiNLeiG42qnvZ2F4cZW80nwReMd2hZsF5qIE+XNdEcRjbTX
nY6Arx3hqoV448bHyXgnI3dZXUU+Rgt1xs6pvtEQ8unqKHzPahNNBoNDDU6SD4yi
gbbQ4lUeUDPd3wJ/o2Yptl2KDT7zICWlMmGZwVjq0uciWnWebei4N3PGjONpruYl
QhgzbCzRD5afs0zXKm6pc9CgkZSvtuZoLQnIFx5gFAngycfqhW4mYEBn2MyooDcF
ArC8I6HnXAVr7w1lS50SNjQpwMd2BIP8fSV6aLDuIVw08sx16jwzzWpEvjT8BcvA
ojzJp+i1Qmw9x1jLkx6GCGnZow3E73euKzJNNNWJvXOjJuE8HHQlpk2cdiZKSG9a
EnOnvTyeEaZVD0qJZsm+mnYzw/ygGkSxE5yYtlY5u6Gk6zB9zMidyyQXmv4WPxzG
vvgYcY7b2MAKDJMAhL2QpUTJbQjRGPIVfAyD7r8BRjwUlxhhPiUGlT5VpEL9HvuL
3Gf+ihfPX/JKlno6+0NZiFP0jrQwQsdbQhNjmgadRA1kdiFvZYOYVl4Kz7IAonqW
O0+x/fP7fpJtcxDN/mDdC9VG7jrHYMvIkhdSRqK5BaKOCLQfbpQjozGy0h//iUnu
OppCJ+jSV7csZQX8wP3ZkXOZzR8ItZA23pssrrWBV3zjmWyYpFc0n+LnZ7WbHESf
s2SyzlHFGkyACdJGbKq54e+tk17yYOrlKXz7cY1jZoSQTOAQT4sqaN+dm9MiZ4rx
6rMe3yeAVNfRw4PL1s1ZnVX0ZK786xyGq/oUDiIFr3hLJwD6+qDoVHd3PlfzEcFG
FJ+3EswFOyuYOUL+6ByLo89HI6U/tF9w9cflY9ip1BJ0ppTTHTf6V9Fo9qAQcu86
/qSRZatheTXi/kRj9xAnHseYrddnYr2J6eLsrULKL7Haq9AA/HSaS94YjKb/+EER
UXuoMMvT93pO5UOv14bBAdObL09OhJhg2D292VN0xK3BOkjUIlOwhDLMehuCbzkP
0zyMHDmOs2VJciFrMCCKyXkYo704pBsDmegUhXKffhOlstsiPanpvoyt088EOnNt
b59ZYFr/tkH77oQanasdv4ZeVQvuATLCHRUxHoJpeP0FIRzLDWOHhIt2h6GAH88X
P+JKSn5mVLjuqtKs20ObS8NlS8H5esTHim9wkHvUk3uEOM4vKeH4AJd211ih3xW6
kmTjyMG0Hty9nrK5R0r1BffscrxnrcIGNtWjF3+1KNmJYir6sUfXWfc/6tDvTFPh
kMBGFkx+u4aiCI+NcFtHmhD5u+z+Xo9A8qJigPyF5PUdzZJIGczD4jqV7dWMf4LS
R/Z9/QoDAp7LQs1vvkupnvqmV6TxjbVMcL/+AJblkU+Gxdt+a7+mhPxFAhHjaJWz
b1UaLPUx6LeskoUznxab/FeINEZCNheYmDt8ZaQkNq0PPlrmtaYtuszF7OtbviJe
C6H9Tpy5cHCdG0xMWzvLsznEWrHu4WRQIzbggEERmrDdYBIF+d8XNRVYZwtweEF4
ZZ4N/PqBUBU1GrT/ZLN61ZBnq0q1TPDaycMHCVUQsRVGUuLN5ypT2YwIuuCsxp6O
sDuxR+czxekcJeP5Kn6hDScgjklu2slDR5HXZ5Nye+WQNcJbWp1yLVr9MGfCk8Sw
f1ickxr8kDbjsUC2/74GoJrDgnVY2oU3eM0fWEj/5YeSLu8XetJNaVa1hvAf7iJq
+lVgaZbah4/nHxbtshgcf/el8GnIRQJO+pCp4QjIDxnxEib2GpWWdx3fzTJD5Man
BCcYmE7R0fLkSrs4vYVBLAnrAgDQzi1eGrf55PHyq4TKmhKFHxeean1VvgdnMvJ9
xLwCdN2A2OVVOwY9NUyRR/GjGwNkZzTmYpOIVx4MTzDXq6HvXo4teQH71w3o0fKg
gn8wLeZygSXQ6HYiK82JN284fHRvP/Q5TJMA30/a95sQlQnmPUVF+IiUkSnzznBG
uhZytmBmZOUBxDWpHTQN+hJQci2ugzM6Ma40hW9uEVFiQYKPEN2gpbHKpsNU349L
66rInLFnIdD/426UvvGw7SXGjn5tbyQdIEc8XiNVneCOxg5gxbbmsH64ystNjyLu
67xgll/Kn07DLsyHPhrI2QYn7EAhNsmUEwmXyN788b3ynmIkN6Zuwf8qoRk5JLMy
rMWubr4856MdwJuwlcBQIFbGjKqnzyjcXq2w2aCYLcK+In72x6ASH/E1Pu9A9Uoz
9cnsKGCnYeOmVY0C8xj37+j0vGw1krrEX5q9BfFSiH3xbPUf4eWmOO4B4Mwd7EOa
iiwHs5Mxe6kIIrnGA/8NZ4P5vonS8+b3PeBvSh0SoTX5BPMfI1dD5a6+qaf2EGIS
Om++cZjaGJvxyiMsJWUS2282+JBTDC4kQfANK6gb69Zyn+mUcXzr1ciHGuMvwW+Y
r9w6ESaR+eDz8S46lNF9Lq+FErXHgL2Yx5t1q9kVYJwen4c87Ld0h8o6ywZi8MBr
4WmU2rB/8X2H3K9am4oEOwnrAJiPaHixoezMGch2fVzxAvbYhR7ziqZ+Da9ZAKjz
YVqtmOnYMzM0JI4BhxR0A5CO6ChzbtRLboeOaf3l03RYfqn57M2ee0omKKT4ggVO
k8Y+sgV9w8nXeDbBfLUhOsnrKjIL0VCyNhbTytCySJAY40fP6XIcixJoSE+bhZh5
nyvCdrKrRWdbiYCoRC5OCe+RdHL7q5QI4cm+a0jcFkXq2b/g5UQESrCSHvbpFJ2G
PmwcUE1Bw/V3n5KFTFoQnj6wIw9UOFdKD/PuiRDDVXZdTkPdoRxfBws8k3wzyhP9
jgTdd78Rv7XrHQvn4lgH79UyNVuKmIACkUIEwlNn/jF3jnGsJ+7dfw2bx5r0WKYX
8gZCl9zh8IUH6rz2AhGZwsCcWhfREITyHf4FM/PX1mZsIbXDcGnOKs+AMAoL/lxM
hmKbV9iiGQ1jv3cnTqLy1OQn0lNqQpbBH1g/zhcGL/rgpQSHbIl6NwNsXq/JV9+9
D4RU+NE5MHmu3W7zVgtcGsvh4Y7qBam1fKRYsYwFGFlOYNs+Km6n33uNAPW2PZG9
+Q9mF9X4GlUo5phmb0QVt8JJfVfRxr6h3IoOmaeu7iW7+0TGCj1/mYGy+wV6IauO
5KYh7DKdTfsBNftkCJfswah0KgEiJZlVqGS0B6k2wHYQiwYehYj83wU94rpZFL9K
k1mSWkmGHHUOKJ+eNPsVEU0pirj5xFj4PhsHq8/c0VmUfub4h2MXe5gwZbozEytD
PWN59MLEZdv2hSXOL40QWofafFTUZi3jGxvF3W30AsrdzVr/zbCNaVaTfQtQ8Cf0
CKpd4EyQwxQOKfQZJ2UipgeQvSOLTa+z+EI8+PnMcTw9Y5sjCjzttGRm8cLl6lhk
eaoeTAnWrIrgkwWlhmfTTeeJC2TTqmYRT3qoha+dGeyEUqxxQHuxOWjl9y1ZSy5Y
IYC7vs5TaVF9BMSZgaC+bMQ0luWGZrs5HyADGIlPmNoyH4fBENCdiQVz9IIyKHqa
rCAI4sFvbf/sKiTojBHeE54OHHOIQeeE7szWB4r7kfb9i6wjBDcxVTBJKWPNx033
7xDigMNRakkwU87NDt1XfPsfHgzecLpgWpTsQQx9kOjF7XpF1iY7Az4GgERmfc1w
msEWQHSfis8Bqs5CGWUxwAy8n5/NFI24WsYw50rrjtmoivV8cUiWUAhbH7872LkQ
74brAwTphqsfl1zHMtIRJwjoljS7BFFT4AyQufcjnBR667L3uoxs7x8CN72lukL+
t0aMEqJC6wkg6FlsGmDVvScHpnU5GeNtEGhRGIwcldx6XmMW/YLl9/vd25rv9q9v
IL6NqGobQtmDDADVSp5auYS7v7+yK5DwYJ3rgxEnSqlwL6yDL0MxbH+Tdnkx8tro
cehWzPQZM7nZg5J9dp3PU3aWKGTDBxRI26KN7xi9Zutuhy+HE9DFJr3GDhu/myeV
UPwP701Bg4L4VJ1Doqqu0O+UnjRFu3ezwASmlliHbxZ3fBV1K+h7aUF8LNvrB8YD
OI6cF1sM5DdJFWUv1pvIQKE5NH9xZySx9rF2knXLibJDimenJ4AraE6m4GPVu2cq
YtD+rsbxoLvq7JNLauTCRuiGLSxPBabevIp9PYtVpXMd8o36yQ+KrceBohqB3zME
Pnl4zMCUfj7/QxeOw1okF3JeyM6p+qXCYx+zjwVVwuze5Phyu8+9TUjVdPJz3nOg
oJyLc5Twtxx/ziUFNdQNKwNakVvIs0gnlyyrk7NfQLt409q+LuBzIEsMA+ftZRAv
8u5z4TfPa6uHhEW2F0lnYtSgw6EBX1UKFJdxIGCy4pdbiudvUULoQAQSs39/ulz2
BpMa8OP41HAB3KEgI31T7z4CdV7gH4h0Sy6xidJVFGM+4Ji7w3qBatu5SpmB4rNt
pYUHy6xALqJy8xcN/sdpkZCgm26fBSBC+QqHtB8J5wBbuAvo3lxv98+mk8ssBsbN
olTGGR8nU+l1zWJjrXi+sZLmEELGNDmslbgB4Kk4fwu2ir1aEcVCSxshw3TG1C7K
AiVMXgXP9Cb5yWvlUWqKd10ZM0Ids15srocp+eoi2cKtJP4SQ8SoQeCxgZkiGwJv
el+FPqGumOYT9O2OtMa9k8r4PiGvujAZ6pfoYixiPrcbVDUUJps4s5WipLOFe4pO
bl5ziIZpdmuAAPBLHkCtUf0GEZqwysTmhYh2uAga89uxK0o8XLLz3SkUSe1eKskU
IC4dPB+xs2PyQKLFExEBNNSyqvC8v1aEW1qUckcdJoWBV9kXnpikKI5xmIvuFGZH
xxOJDxox/68D0HI4tbrdGjfPmKzkL8bK8i8JPlG9EFUavnmqNaR6E31G72MaSlyE
EPa70n8DvYWUtHgGIZVGLfaODncrdY9NgB2byGNp6OF1I5TVweAXaG3/FufBlVzV
gaLz9iajzrZPTceVD08o4AZuxBNtVIapjVl4QKdfbqyd9908/rQOy48AeOSP2uc9
hhtNKIf5baFdJ4QIMuK21PYH4qX/vlv1jXAMB7Lo2NkBssHDZF6NxroPEivg6BeS
vVKk8edga+HtojmDkqiIQ6J3vDPN6W+TDVL9vh307X8X5M5W2jEiTrbho3ZF11/o
FA9sZPbX0TyhSMlfp2BRvlHgrA9GQbUeZvYCH1ItkjDJpH0RikQ9sg9mu6LNOvaC
Qu+6HfXAk2BX/OF2G0kRj9VPRFGQnyTBtooCooEWW7zn6EGTs/nqnw7H1cc6hdsk
tnDoc0KHUBpKCAOdvklh9uqPWVrsMq/+qPqP2Xko4rsnUTjQpYFqssSr8P6LIpG1
zKIty6MbB/mjXIuaTULARkggiMa0xwUyAU63VDAnuDhxzfoyKYx6T7lirVOGd36F
YqV63Ym07Z54S9zlJnJTLZcV2k0uticr6qNe8W839aVvFbh5NonBmFbEf777omOg
Y6Q/9nZ4bbDot56KM9AAI3XcIpvjgKC3x8Wz1M5u3idvlH89M3lXOAnP6RxIjqpr
jBV/WdD7bOcgL3UCI7Z2vc8rFli85CHe1HeFTMb4Q20LN4RvJfUZ/Rna9Qb8A27L
ZayXaXcPeUSGzirMhDbNpI2ek9UKbgFtiScDX3QBudQ9eOLNBPDbObjaEpPCBFmE
zjFhEQ+aSwO6q341LRXStaPDBl14C/ivd1NPrMMsMWf1tXQV+d3AuWiUUdU8AUKL
jUcWCe9EC3XRx67W63dC7bEHPhaCLoc9DSy4zkmJWlevs7dhhd+mjXl5o5GrJrTo
wku24RkHxd0ynBkBsNBjMJ/rTvth43jcsGTfzRx+T6K6PcTzzZVfGpqVBjJW6Z4A
HYCo7hx38/YbgUL4SEc8rJcPf+kK7LIImo2dWNnUhSJsKwcBZNVrjAYPfr0NxCaa
enzrNK3a6txVLlUs750ygXm/nuaTGdRrH4aGztXuyyJAtq6uo8UzpHkzptKAhU5B
DBvDaX1cSzDAdTC2C24PvUctkNEH5G3hoGt9dOxPWfb+nBK/XastaXMnpP3c55+n
6ZKSYqPAqvurXxSGH7iZ6cHJo1h1uk9XHfP+juYxMn7+aPEXFkoHkxDaDrNnc7Ke
AsFPwrcACIeW1t/lMldgcKyzQhgh8xsrCYgt3gDRwu8/seCjj8/QfpfqWNsrYs2z
uXWtpclgst0+eIks4qFos7TeK+Uhl+6xy/wZL0nM8By6yzNd+Wxn15k5QZqCFJhU
GGet0VMxvNtYpQN5mCYtrRlwLJgpc+0F18n/NbzRc2hJjRT+R8TYJnkQJc/HBUoB
8B2Z7lHNZpyXXH+Yqi5dO0SEIPvQVznnYNKVeAhvrJHp62glNFHeXrTHoggKXbUI
DJ9Sxir5Dee+u9V/KZafJrhoC1vJVpuRpEAPYrurkqGfxp3v5/0mffV2+hZF1qOg
bGiM1uvTsqGqHcPaysYwgD6bRjVNQZbvVa/ES5vTS9VEnE5gGuw7aO970zqvq3VB
sCYYLoesVVFKOym4JYfW7FTyBdvfmtRzXiwx5GxlzqXcR2Fm4Q7K4aOWDOoHumhs
yr6/5dWI4/qVH7XcmRKkxFLlG1ZOZ+7W20QpOHOmMKpv8NmpcOA5yZqG2n3V4j/P
Fr/pub4I0kAcSAEf2Tru/+mbwbyKEpyuqVhlAuZ75EvQId2jQvL37U6C+O0y5/zW
qMKuXJ6ojj/AVcWym4jzjwYaqrxkSMrKsWnmJS5Fm7ne5qlJYswzDEHFNS94V0LK
2vY51Kju/hcuX6j/8mf6Z9f2Cgyu9lhLGwsbnBV6ZwdEsyuuB62UI8+bGDZZ2i4D
EpBCcOx5D37qbH0nUUaknW+/BCsO2iEU3VL69RWDCMZXP3vjRLiwZ/6PdsEFNDpH
z+pjR1O5sAcES+B+/hAHnBDpAYBrhtTXi8q5BpIG4P5tIsrPYFbULDnun6FCjjJ5
4y+vSRD/q0Ov3CFYZsw05+B9jTpFr39T+exYd15r3wjYMWxY9tBfpSX6sp3oELS/
J52hYpTwADNSMsEsCSMOholVNKy1N7+IqF62QjdyVSKbxD8rwqpQNrPR7kpMysJG
iviurGOywSZ3mMclp+VqRFSNumj83TtvdYdW/jHYHA0ivlqLpcI2hhZROAWJQBmS
DDP/FE7zP8gcj7aI7AzVa0M3x0XgKS3AY2AIbXFYMOpJYk2NjZ35elNHaj+YQwYu
gNzS2hJjTsH+2eTAX/VldJk22Xlz4vDTV2KcoYJr57Wf7SdXkdC8jiu9MSeoioDE
wOCDPHmTGLFaAFFkMpoS7fKRawBZofHDGcNHDSV2BvAVd+g54eTn/PLUyUJPcGvN
dySXTl5XoUWRCYbJu92mD2W/CIKGKivWTOSFizn6wO3wqV1X7TdJc8AtVTVt5tAg
OmbQhuf7kmGKVlPIg/9de2U7bbSguRNJGIa8KO9pn26/CJURIV1RdSNCc8Y8IBDz
dmNeHT/pskKJhHxEw8bonV1kvoAPP/NR//clpXFyWoDaSVVsNhJM3YyYMxXBveVq
XBF3vP/mwG/YceLJZy2UlkjJVn3GYPj5ti8p3/O9/mRYlXmxxZib8lnCvfsyP7c1
TWnAPRxAIJoer4+XtK7j08K8blDEblndAv1Atz/3QphAWW70oa0Hdukz+fkPCuIx
wWuCeSgRxNq09Mi7kWr1hi53TNbqn9aLsqHfKil06ee/vKEe837uw+K8elpjDNHk
VJaPO4l7416yDucCtJY/xdXD/0k1m8F6+TKGhoslti7LvxUJRB0HcvdRCssn1l78
iCVZZzn3hM/z3FGSBh5voXGFpTOj/6mV202Haz/Ek0Mfg7X4nHAj+u6qJuSFI2ZR
TdVyJz1gx2yGw0eZCMqTqrGlsMRdvLTQi4Ad6NlHWyvzikWg/zSfaM2qm+4hSfOv
HSw6JXnnEuwTUSpeHpKPeC8HWSUsi/PuKjpUEM8pMM/dFU2O9JL4KmwstpZBiyRs
sI7gosN/RkS410cQFG5Pr+al2PiU0SveXF0EXTmOWhtRClGqB5EYYkCU3VAa6BxK
Y5DVrNXzxF4Y1UeGMZDcdjeCcFZ3IW+8KvUpPzJGfZ/NlRSE0zW639crZMt9GRG8
AHoKXyzwWhHwoVoi+nnNF8+uAEHELB6JutrCAAQJ5c4cL2owbFlSnigdVkM3bOBI
2+0Q03VxdpWryPdOmxrdLsTbSWgqYchjUnM1VIbfzOsUiODrDTvcmeRry+niKUiA
5CpO8ByBYHGk3fGniZiB++aE4zD3IrTHJKMHyMMT1HzzwseDcdI07W5BrZP7kY8n
WnuXFCSjCpvcHZRsV2cPVfZOLtEEOH0JzsGjSY/SZ9UE7AgjzUg5TEZoyEL0wFmB
RcHoWLX9aebsEcF2tQP3iT2+l10X3VThGYvZK1KRI2Jo9JEqr10TxKf3VYX5fBlB
DtfIw3aqRcfSqEJk8HcW0xPdy11MCbRuC8zF3uY3pFVvuSoJ+L6yQTuCanuuZmPm
sIQwwCqs1Fic9BGfAcNyR7CcO+/Z4sYSPE+IsxZlZK6c1+DCIas3cO9BKSXikg+O
uK1awWfOLAZ3Fjd3XCfVRlv6YjG5CIvMey9K/DIBjXFF/nMFfRVG4OOKmLw0cAud
Wz2HgV5MwsGUU8lStKCFROylKI2/IBxqu2LlBBJmfYWJP5+AK0B1VxSGzCejxQET
7s+MkjmS8LzsgQtbThxD1RVVGyqrL4aOVRX6Upl1j56kkjtRfFwPYGWMdCdX5YQC
yLG8DAlUJBQYg28HKAd1rVVI7vN+daCTNifm3sV1iGGcCXshq84LP9caZd3ZeCq3
J/qLYehDH2+h0ltS7LO9nREYruw3u5CLWUgJAEkxr46R4rshGDelClyn+z9YdJHh
xLn2U0fCN0+nUPuY6ExWPrDk08wml+v1e9myCMOEfi2NhEGchJ9K19n/REBxhBQI
pu90Jdv+FUQ4Pg8DbJodq53uwNW2nlBPRLI7s9BkfXatkBvWuzzngjQp1Zpiz8WR
Htkv8mKvZx9RolSoDK6pi24I7akZ/TYVC9sDpJP4QtIPijdOq72MjgH0EVHdpOHK
u5zSQ6Smhsq3Zbioh9BoDyMeVm5V0/SZMoEVA7EZHeWqjA26Nrt8W30NTbzgWM0E
0aZ1k5qX700omU9oTZsvdn0/mLsWwOGBwA8oo1fm8P8WO/Gex5xo5Q/cz96q5+j6
YpV9Ojzmvyex4/XLBfjLRSTfdrQhL9Az5EjsJMfa2PkyoXD3znjz5AMxa4cakFIF
/+Dbc5oJuJ49tNuf3rS0HYcq61RkEX0DGJpi8uqyxBQs2iE9D/7dXLKtlEjQ8d8D
4iZiylj27EyxQAbIH1N3DnQE6GXZSmeI8TqgMbH10Vfp/tqoLYvv+rLktZKT9pOg
llBp2aScZmeou17FmSNk+R2EU4a9viqWSWxWJ2fHhLtJmMIBfXd3BIpB4t8WI4oT
GZswB2/5eHcWOi1gVNcVtX4cUv52jrcL97bskV2oVZkjEuiRey7STQHiPHKHBdfq
AFkwG93WoSrmjwMu/WHcv3cZpCIJSBbrybpNdZaCKzspJGvVvr5YvU/lJnDTJ5LH
laYNDu0G0lAMqDG6iL2JkCaUnXHyZ8qBaEYcWZUzEL+/kh0ZYXbDKpg/rH8D18lw
ZtTNxAir2Hjtblsv24FIIDGbpVSD02sWf7NYYNJlEAGelEK1LGQLWDJs6j+zy2tE
wngmTyIgSRpZoxaTz9sO+h/zT1ImK4UlAP//DtAmk3XTvwvAwk95IdtCfpFdzR68
K3uGsnIECMJtfWZdTt7upct2m8pB6hLQ9CbZVndiWjIYqlzdsJ4NfZHzF5XCPDoO
NTlxZ78ovQdFBQ9xX2QO9/GqJuNf3i6uEODPlitzS8PXIbootyZaYu2p/iayJzQr
9fdiix/oXdPv7CYWYJ0sp0Y3lGrtMXgPZIaiMjJ4oMMC31OEXbhyYOuqmuvRhiy+
z6aY3MFt41N5CUDifx52PzhzJATzLGnMxbXlBa3DLnVE6L/AYquFD7cl1YazRZR5
OL4Q5RzK0K7WhqigpIaS2HZyFjEew82oJ9RSyQvjmaasFuqBYL8mXaWWMptb21yZ
HJsgOsZyD3FsEtt9RhkiugfVrKDG1ZONiMVTqCHwVLlUpvH5VZwruptbdCNC/qGm
NdOWepm+40VUSBG2B6qPgD0x3oV6cWAbNvESq/df4sdWwu6m/NEbcxzt+dv86xnC
QRz+zD+qxEeclysGhHWtTFm2Au1WlU22F5q7OTkCR6mF4YJq7iTdNp091RQYUigE
nV7nMgyt6WkRnF8q2r7WI+sc2q3+DRqDeyCv//2Flf2mQqD+tGStHgJIJbkgreml
ADQUmi/lqMpZba5+cf+rxuW2BH4gKbgX8TMfkj4ma4CXIN+Sv5KB8EAhXFEvjLXK
Eg/biaesZeV7pDSGTZmUSLeriTBjLHYGSEkfRCo7KDUH4muTfmmq/c/TKeUcUzR3
oa/GxKYl4c5fMlPNdCXwZTf3/5uUZVUDNc4On3edBFH92QRVhENptMY4rMgNRZSI
s7rNd84Ew6xAw038vOXv1XsbjHDHU74S+82+L9Dyx2rearmLNweYITKag6oPVL6w
2u1WbETJGrY7JHtPoN0o2EGysk0g+Jrx2b2FVU8P9/4cDv8AIQ7+ypOsc0zXb0wM
K+ZQDuoYK0M0wHSCZmtqggf45OgaaDDJ67eO1fVtenB+srwo8gvHKQoXxV5jxXOM
GSGm+2t82sGgK/U43yBMdcmkv0iWJ9+ymdYiYg1kYbFcPBfcxpkqo6JoKPNnTK/q
8MRIykCDxqu1+uCiIYeaxbq693tgUEThgPRoB7Y0an/lwI569Q+/Ftc53+61Fn2G
eeYnsPuuh9FP2GRxZZc9G50iAWaMNl8RlUqPtnBZgpj7PgL1k3hTwuW4WGTedWKo
7VZIr/6zrnmBzZ2aXCE+puo4UA83/GCIBFjx9b/jmVXzJEWmP6sQ2IQ8FDbHK8RV
NZRVb65LtgjtY/aKKArye8KxwAu0s093KTPZcNOv3jnNttnMeqkd1YAUs/+H8Qx1
3rxc0MlzKb1tmY3rptPYiFIxlh/z4XaRVcEApCnSYlj774FFXt/SUDTczWnhrb5P
HWZT5lNpBoccH5obnrtvsQs/wMDondCm5rbfoEuN/ERoelOPriiL1SVgb2MLe7+V
jHvzbfOq2xAZwoulQEw8ZXNLmAmt3MoYA1mLsbWjyDkgDCcuOUnvxd9mC0PwTV0H
bIEzZSYpY0biq9izt7PIcK1lmYUHCjX5yosvGli6SYvcXiGQqvpT3Z6pKsxXWIDW
5RMHv59hn9u/Pl1wzWDpi9xW28BAzkZkMVqgoZMeKMfiNg+CLdUWV2Q+E0LzwlmW
DCRetO+CggP2y2f+XZlceCHcgN5V+ebKob5FW9oIX3GsQ2hGghH13RiqgUjyz/VY
WfNXWJ0si9f6ldNid9VvxdfgvCzljXUDK/KMC3KYZTLWQpBuQuTN7YciRpcT3iTC
yTXT0ZC4D/MAnIuC2IN6Vpk9N0jRcIsHow4/TXbTAQ6NwklbyI95Ku6aiPlMCCTD
tP5wL/yDujq+kGimRQFd+EGmmFBT8X9sEshVioF2ExrIszWtwiCUNT0Y6sCjGIcF
jhQik0Td3YWLpF/WHYgM08vnkj5E6ACvrgMWFsHmfZK7sBa1/TghVYTmrPhsxdUP
wY+RnSjJ/nTBWrKbQNnIU1qxGRezQNAYJpvDoUdaHvHhIsRwYEmqrmZfH4662rZ2
0yqIjFCIBtyxls1fb+xSrC4OP46AM/zVL6UigAOacEXg2Kty8pRxYL3pHD5Kuakq
Z0pqlGmFwEjH8jQR+iy3dh/1cwwEca4u2gPqnAxHbNLHZGPiHNgXn/iy09G2A+Cc
FIfVrwLzIslnXFKDz+qo2+Q6Z5hjOJ4R0gjNOwf+2UWJWJTWDf23G6+xU5hXMTdn
1KKIIhk4GJTTlYgoxv96quEftILBHDJW7KGMHjM70drUGRmpuXBEnxW/MFtSdsm6
f0VGlzqgL+QNrMkOptEplAwL5Cu9p7AgQFQMT4ez5cvthUOADLXj7GRAJolMHNOQ
b1CqJNt8CKFxkGvOwzvVCb+GqLp7kCyxywMe1b95EJItprsyur02g1RM6UByRHbb
kavIh+QiZix3dWEY9Rxhp1dDMm4jeM8cToFqPgW8Xlr6swJ1jJ9dF99hMqjuw2xz
FdrrmezcZ47PeUCGP5o8wyepv8MZu6xZKaeiDFmuFw1TWeiIlte+FXZk+MEeR67D
ymTLSTtojf0YneQQ90aJY0sF5TeoK3q5o8PJYAjlIRa7DvOHb7Ktx83NyVYDAJuq
duhMwBBnSPz7Rivw62xlcWA2d2qa62cKJF1XgFgKyXM79mYr1YcdlGxYLPdpKK66
rAR95IVO7u9pedZz5eIF2EzyfT03K10pKKvPCVQ6OUwBIi946HIr5o/CIEnhFYC4
zbLYIC5Jgmomitfkk7PyADO7w/Z0N6Ypp01Nca5+yfA3GztoYEjG3PdLgxfKUUAe
8dAat8sixdEf2fA906p+jkBEA2xVVDsajvtPZaloS5DZiVmCpn/HV8qymuZsJdqW
jj28EgNlbnDJS2pZ+N7hLO4bRdcAcuCqWp3PPo2WOmpWGuOk8TglVsSwBj73stop
HxX3B5WHCXHCp0UkVcDnYKVxDAPfLS3xJMwfHNlsR5iZA9yylSxKwcjgvPuzxmCv
CC9VXQVNVfW56Qu007qQcNzewgJCSzf3Qs74x6cMjNzyRsOWjjXeYp5YyObtbnH6
FDTEKkhp3L7/foqGMsz26rvU1bpFaei6jNVIBOrjkcFa/Z7N9T6jEPF62yZwcBAw
JKqGULKpgGTWfrJyoLjk/bktp2tor8KaMjCAAiUBoIrM8+JdmOXbKGHJow6pMk00
hsahPWGjH3nf2pbMywWsdrgp8LPDwyr7ZWnDPLXkgKvFubCO5XBCHmGP8m1biydO
FZNpDb6GDYeefmxIrrnZ+tuWpcAIpu37y8xw1s2GhuGmhXSC1bAQSgvvcV7k5MRh
w4TQGNxa/uIXDFpSZit74czinmc9eXFNEf4hROO3GxGZKsY/bBMsM6kP8HpCWf1g
BIOEX+C1iB+naJDgn9mEwhei3VpCgfqiyx8JTXh0v/Zkk3wmARbnj7VGc5z8DRRG
710gkyWglXXFJiIXPmFmmrUHp1jL5MGqTDCffs5+tTLPO98+ozgoHr5BFhuBZYwm
rv1L2P2N4teioqJ16lZRVzVzticxbKwl2C7ldl7Uw8UGnpHK9gXrms2wKcrnj9oz
lFScIaiE6A2SrgBy2oVC1qJ0zpaMN4uUz7O/LfiVHlWHiikYJXARwzaMY0wANCEp
DzisugGwTyzXMWy/1QeoK62tGP8tQMEMytXHZaMKJYCGb4y5g92qVe2dIpQlNHQs
3M8jaRitRRetfb6FOwikxWJvmujowbIWMj0qPtr4dia1GXTsTBY66FUmoi5TLRg1
zHnMviSFEek/BOzmJZOzMJv6vZBf1Mu5pxfMm1bH2atiA0pyp/LThGjto6snQwN/
Q7Xl0pX+Kk7wdx/RSN1Zm2TUmUzoy/j6rxrO17krh+8aEstPGvz69WIvB+orDMcE
7Qjc7qBLXexRqhzg2doIt7cGN8cDusautD3mAZpMR4QYUP5GX8iOw2Mc2Jbo918p
W6349ULL6ZGzeETOEk/JWx00JRCc7V0PwUhSl6TkNOthD9RDFzX2IqoV00cqY2gD
eZClZJTvazyvheATZeT12BQzor5dWCuHuhMUcZrknNoELT3klj4didMhO2SY/9cx
Ffi1yAllbWQncr0cDYwAOYXeJC57UlRku9JLdT4dmHSeyamNUQ7GZaDXJZCO4BIo
7efkIULkug85JFFO4X1Dh6ZucA9WyCvSj3MTyP14HFLapL+pbKZSrxfmL/z/e2U6
X+iUz0F2WWXjB2FCWY3Ymh4l1kXDVe//GE5H2GfP142dJGfPyqSVDJYFQ6wjgMz4
kCaVKAEWOrk44BfGHkfJCCsGA+5pprgZWUWpQPJ/do5fqlGF3Hyc3KdwdaKZ1hZD
RMjZUy6YvDcjaSqG+9yuTgLE3s61UJqTE/IZaJvdcN72RNtv88ENlgbcKtBOcgDY
d7QdmRZ6fL4QmfSaUPVtUZP42lwzEdJ/5xryjgiEy69zJdkBawuZoMdR85zh0JOt
ibajnsvK7hTKGdJKV9D+bbZcZgyzWYkLUudUlisJ8HY5Cvkz4rLJlEWuLSoEkeZK
PbsupT7zL/j2DoVG4k9qHfTOAFosxDOfcBCZ4Q+a8lMwHsuwNZ76r4COTV9pbmr1
b+OGyxK9pWFVVVIjCcelKMQ8MmhoIj4WmvGVy/1PTMYrpqo+zmnDMBEpc6uuONZT
+uSFWPXQiwxjod5s+cEB33tApdewQHrGjtYhld7ps/3137Y76snGegIWv2HF1fKD
2HDA8D3H8fyj4DsLdlgL5FMls0tYlrXbdDhS9cScwEUWtGxfBL3ywGxebVLQIqgr
fr5EQ83NlTGQsQA3T5geAsyK7mx+rfpfQDRNqv3u2i155uIrSC64Vv2Abib4HI/F
lt88i+58ATGKTtnkD8bVN5ClV47yKLKw5HsRWq0u2yxeBJtCY5GT9cVYAJxazVg2
dEEzXT37oz1PeLimSyfmmeHLHsvoKvP9+MDw43bJg/Ob78q+LtD2R2dNrHkppAU/
Hboha59L4t6D21y9l2vkx/TE8tSbce/diUIa9cANATe8mmFLM7kzShWwlIvBuG3s
JLHt0KY7DvAmNNSU+l5u1UPMyawrv6bwEsrKJBp9bJc0NtMzvk+0TBSRUczEd/17
pYK+QeSz+qHJmziEiicSEyTEiSPAyvkDKD+rxrkygNsfgW3G7vQAqO4JABcV3yzV
dCAFudajulhOl2HwBL+KM0DlWEa3nwrG8Y2ONbRf2YHSP9GWxTrgXwFSzUFDX9kl
vBg9k6RASiqDQYbcH4VozP1e+y9dji/f9os2wawNsPKwDgUuW08EveWdEPxtqDQ8
1q64FpMVaa87hBtph/P/ZxEZC/59eAoH5FJgIS/b00E6zwIgkY9sarG0yqF3oG31
B/3qWVJZxnWfiXjibp2uJe3oOGUW1aL8dikevcB4LY6TUZ48NYL9tVvQ4dE4YLmE
McTZp5JW+pz36yFUUSfHf31p0rIxNwRZKujABRX07TbfYxn/sl/OpLUTddXBGa4Y
DsI2R+fcVxFLDwGGiYWM6O4Z5qAJYYXaHjcHwaSL3BtvxKTJ48h/lO8bZsBQ7OhY
+AjNAKABJUecC16bn7qIx5QygALthrqtfwJSlJO4rvclVtkc9jDM3C1QT+WzUH4n
0KzBKVJaekngaxiixaQ+Ge5EWi1Myigz9NFns0mgbJ+iqKGoMPyeMSdU/18NAIyA
qWVjx0qnkHFlqCUnfqdoPsU8a3JV56WhNeSqLBb/0vX2dhxTvaJu6tjLJYocW/Tm
m6+g/oiWLx5Pi2PxPTwvusTJTo6O5Tyhei1yq25S0WTSo5x7NNjTjwvbXdYDO2iW
UDPhw7rhdNXpmzUxlH0qo+i7mrpTq648NlKby7J3ztSKvW7XxP3E2o63hjU1zuH4
ki4Rt5x44t4b3XZj1CCxKGOeaKVKxrWsl7G5QhIlcAjcZwV+GKloW+aFpb6WZ81r
i6TVQSsNovNl9YIGdeNZFP7LTuu5M64xbuP5lkvKCo2Syvn4J4M4/4qQQOjGJMM+
TC5QY6WFOn7PHX0cRJyVLgs0jCZPGwvXxwfIf3B6tpAnEwXxpNCHkObfNzY1d10R
wm+udsUIVKmukbkwUVRe1ip2+JFMXeyIJkOjQnHHpqLXc1UriyNMIZ4U+7S6gXyP
g6aygHZ12wF/r1b8S4Tvns9YtB+NDLZJjuFglX+eZCI/CQZdWLiqFlo5vVMrtE7N
XrLAGXxXmyi3yg6ZHKl8XVIIlLYYYZnr3JeyqduFK97+D0357iUVCHCt2+TEU+Nx
ajaaLI9Iupz8pmsyP/3cfRIYZRdg21mF0+KK8e8Ad3IjEkaB+H6o1/GmMuv0sa8N
Zk7oAuyfPCSbwFANAw81JDP4VcW7z2vRU9TuRua15iMLRcz+izjtd9kln/HdudZA
64zhOrup4pAVUar4ktvB+28bSFTUkzqkHv6+QbYOGRPrn4u19dP4sHtGs7srF80l
kFoKPnZ+rUqD9jle+PuHR/1W1/BSymUr/QUO6TKy6Caw/rvMl04vSCusXyDcemOb
WBU/vJIb24c484kbqObMFAu065x5Gr75bb2jsX6SoFeYvjM+9PWTuGlOgJ3Jr577
dyoMrqq76m2uKdNJGUuZuwk00nllSUbWXgO3sg1fZNXLK+e0wtHt2QzmReEGjQDJ
8BO4xVfc3K18Pp4Dq4xDm7G9bQ6YrMxSq1A4Jztr9uLm1VWJSJetyvsZRLp2pzbW
Ndi5XV6z7ANryuMHHzv5XLZMAmIgU+J8Oel1yoJosWwDXbWtPASMsGa9cpXGwO8g
QdM4hnEKEZszatlZXpMHkWUkKAHcvyTC8mdiOHV88vqjcSqURG9LZSzCiHSCJev6
reuE3v85UPq/GfHe/1Cw8IxhJe4449IlM1FpO1UP/AD1vklj6icu/TXNWAEgmjSA
3keH4blA6kJEjVYAKE/f3io9Gp3Ds4EiSvPE6R8k4yEOQilW4xBdf3pUQz/YpSzq
H7RGb//q+hubuopMJWPGLMJurR7YVb7ykhH6ncgJuKEey0fdrP/yBIDKeOHEM+9R
sWYlJRKvB/ZEoe5AakwDZAhQT6MZmWYTXRZuQMOW3OqKB63xXQUFA/VfA7H1wdmM
QRzQS1tDy+gFU6QUiAqriqMbXGv4R1p9C4m2+NhJSmBVcntinEkECVl2dFYJAgxI
ppx8X+Mbt23dAAY2aNUQJWGQpTO6JSvmBHF6dU1KxeOtOxteJk1Nn+0w8wvtfjEQ
M1yu5E9ztoIIayN0mo97OvGlxNK2/kLi2RZK+zvBAV95xe/mfIC0s9bNl8N3FOYH
YuQLOvDZrNPQNZ2abtrwbrUpYJp9FvfgA21ua/bt2mIrUldBbcDu2iZHL4vPj2Gg
AfApgTEm0tenotMaTY6fCL0yIU2nnJmJJiYbR3Yh9zr9Eq08NLXJHUnk+Be0tYAo
9XObIsKYfWTKnNeha8tJ6R9AwH9KwO7soOxXGroEla8pPZ8BUUgj6s0bvANjcmjD
CprwwrOfNEYXnf0JJQkGMfF448AFd/zN+z1BU5fbmPaa1/9x9HqELjTzg5dp0kLz
GSGcB4nmyR/ZzUr3nMs+4ErXq+5U2ALFpsGPRWpwnXFxKfhhdL2+vi2WJup/+sDB
/tkLYnCHv1TXRIf/wQ8YvjNvj5W9i/9PsvvQOX2vyzCdltLY+72S+CFWIifZZYzc
cAOETlqhY+bOXMw4Zor8UJhbhNpF+92MpHDxGEZ7vk6T9GS3iqXYeeDkcdhqHHVH
eMKNsMRP6zQVv0rtI5tZxtG9WiQFDoosmv/2JebkZy4947lsnBENvtn5uNwuv1eu
Btd0OgrD3SXJW90AmcCKq13b6Uhf5osWgAzpF6wbYxNYVv/X3J/QCoaCbj3v4gTb
OlMopy+3SIiDHrNlOzQfoaY9ggLPDq3UUMxscyi+sg0nhKzZMCTpTha/Kr+fp5sw
QY1utgrpdaXDdDUNAggIJl3w5Ir+WJQ7X9HYpPSw6JQG9xuaOK0zvFlhr8yI7RaK
aBsGWrTulQpB4BK4V9JiFrexIR8vmd1Sg5YubbH1xpReIVeDOrwB+2Ei+P+IPC6r
wyDaEztjzQdMnqM3Wfd6LnkK5h7F4RTmpnYeak7oIdpH93gx9m5AuA3hhBe4y/x5
uaaxM7MHzIPtT1jPJGG50wfhyi7gatJ8fpUUdnzZ+sXRwucz785U3JLvaugJMPet
dipzlYKOBsiXxLMhjkV92+awSVUIBRFCDqRzQneeawj1qliPSiePUdMgIg/NHD/K
3fYRnCf+8DJQff3a8TXU6goVAQqmyPRZZjdKVFYJLpZvDP5OF0PAV0+L1tXrME72
77iS/KqYeI2aiO0ZimSpS/rKi7FDLJZvSSi0zKyGKiBjrDaY0kcccImbVoMlpAOu
LXJp/13AvI26yUIemKC6xfn87QznZR/jsp5cdg6YRtlosHQUUuefMSE5c5Z8iN0t
yDet9qebPJNoT1qaRQs+U+OvTJGMJR8JwfsCPwGXvAPL43YIKkiX+ZB1BT7bh5Kz
m1h6siIRbwS/wTUGW5SIGMxB9wgb1T4H+YbHTNdmewHZ9jgb5InQm8DOnA8y5RFi
MHGMN2HQGtAmr+9ESXmzVah6OS001Sqon8oWmkz4tvV4uwUpEloItGrkauwfRGU7
hADL0Hou/j8bndrErefiiWt7swJLMp+mVe//xiGb5JrVAPlZe5iLUT+fBXK4qFeX
5mmVqTZtYYZs2S/DfzaGP1b/tLLlJNjVWe15YwzH2p02r8wfxAepI10gG1xZGiic
gbAOQRUD3weCa2qrksWvsA7/mQ5r2abmKZWw6VCSx8ra0JGxHeq5Zlx7g3ZiylUR
yzAVr5VsN4FNdhN8jyMlDh13IbUZ8WdNQd7L59UG4aGMUaZr0TB4VYiR7i+4WB/f
QP4uZWCbFn6QRvYCfDx7aGurltSdYE1Blb7GVHXzsNGf0e6zxTSZ/6fu0SJCYgRh
3D0KAgpdAtpqwyxvBgX3RsiT5t004U48SEfKJfKn6oZivvzqNcy+2xCoY2qY+APl
H5Saln/+hluhhrBttNfy2RCtXGmCL/WbHm5RV/Fmp2zaI7Bk5nZVn28FObAlQ782
NoOIgnojNbg0qvKvcTIM/jSrOpRCbNNX6YVUWIrX4RsDTx8BaxCfSU+357DgQaV2
yuUe/+VA+Nij0ALAyiKZx4CEKHq7liqg6wgnm1PaLKfYY0m1b7Ebdny00j39mIEN
96Bqp7zj+Y50ywn4GtQ602jbF4yXR28kYvRPZ5iCzlAA1/vstYoOYccfgWbyZAll
c1uRzHcx+DyqV31u5EWLVhDBsSuypJsDVeCAzPg8ck7y7bno5uKO/0EDuufcqCa0
CjDpdPf4cICBQe4Irn37MA5caJtewHuGY2WZNDXWCWUQO2vCNV2cHnCAulu2GI08
OYmuDKAMMkEpnstntPKvmMf+kBy+08CjnNjb/IOsBHaz584lIHI4T64V38qTZ1P+
cnWnD4SSikkQ5d1UCxe14diwtYAgPJU1YqEo123CI8jPDTB2LMkRZacRNs6lmYbm
rIxKhR8TVoT6DS5RgQttWmxlk4ZWQr3+RcJrzOAQJ8iiSCqAt4VHkZM3eb/pI42Z
cLDPYrENgRgVFunntYG3SPWfW/nr9OXzjnnhqPyMlu4wl1ion/I7vvP3shxsUn78
DxpqYLMsp9vk6GJVSMRKkq1NcJlMUC5zxAsyd+QR0/XUUm4Gi1VQn17RDi7vaJQU
rZEJr0x5GziooffFmsLDmN3+8pkKDTI4AEiOxT0E/da/rd+E66YqPtkUEsaKxGsJ
ig/74PlQPcHK8OJWDRNHpHZxJLlPj6Ky4mYO9H4X5ozzLAT97R3x18ZzcpTZmtzb
GQYKK5Cdh66sZvnoK3MEtzQXQqILb2TAKL4CHGz9UgzNV1pTrXVuo5CGS7mXBwJ2
oWTFZ+fuaFHoQFwgsKMSyQP0CIKRkrqT94jtNpwFkZNHm4JK2AGjWRBCiHZHwxOn
6s8SXk14X5aVdVi8fV8xAYomtXZAVZgz/B7uriDAmkZ/Uf2WYKB625EqviTAKi55
fu4EZlf4lHtIu7iCxLWMztDN3JB77rSDKgRX5IdOzVD15/qkdTZd8GDzMIr03jCl
npdTEE5yMQLsQTs9XZ1ySi6qtemZJZKlxU+NkgSvp9cfvvbJWmVuFTF3dVUkIPq8
d+WckB6yI6XYQDuF4mJWjbZJKewoDor6OWJpvzxZm6Vmc0xAZHTRRarodi4nQknE
aVVqRrPdUbD8q3IggnJAszdOLpo7D7a1wz0XvEolgFSlMnY17ongBFsM8osNsXgl
J95GCbzaqO3CJ6mft97UEfAZDdXCo3v428+hU/xyQuGWKlqzkFLU+AGuu46Nk2xv
21m+JpxwSabc2NvjOLge94xKd9Ef3844D6A+1Q7qBJMX6k8bjn4ngE6L2IsxgAwt
c0e5Rsjr4H2lr5zm+qiucCN8ZAljzW8/7rVRl+BQ0etcuVFN9cJKGtZVnwKEBtU9
3VgPPg7cV1H1/ci/IMWaXslKJ0wqw4VEQhETtkp+bOSijSiA7EzT1mj3XfB70Tub
Wa1WRNp2e5Ycf4XzfFzJDUGEDRTEGCqz0VgPVLgqUmfHF3ALcCqTmRzRs0nc8BgZ
Y5iTUcANsxLNr0CI7joZ0uyi0I14Yw6sdATaq1X1oeMkHO18foL5pTQ3wjf/QxKW
Mhp17y8lIx3r+nSnDHNEqHfykBLIJ9ndGXbJWsNyLYERDNl4gH6/LKAO/v78J568
mjcqcocYIOGi6dM3o4Dx1Y9xICqk6zFWBmsKaCn5ylEoVKqL/0K239MB6Q6RXRRy
8+35l0ng3NA8lw/u7dLtsYKYd0caNjoMMxuil3XA2sllrYwISWo3EAmg9Lv/xoQ7
xYjSZHNymbuKWSwiGZ9xLFQ6XoIGtYFhGLyKhy6lYCZ3ueIPmiL7N/HhtkEynjnR
14HLvAzmMJ6uiHKpY7zMDO7OcoAJ0KNfhx3Lrql77TTkPNWsOC3P360QR4mEU4M5
bnJdfXYm/Lkqg1l9KZnvDykq8GXqJ+JWmG3wjOClE7p1AaIOtnacjbCEnQsw1e94
+AbGX7gHbq0x88dSE96wXTx/mHx4A/qYI2FH45Hy1ReBDKOpdwMXV1aLfP4H+5z+
4ceyxWgRJ+c/DWE625nMDxLnTnkWtpc2aJeZhd/0/T2wY3BxE4KLvsVKkz2g++ed
uvamRkDwqeGIKOwMC59LXmSoIZ7+Yq8OddxpNn9SvNVO+jv0G8vTOLEC3GcpjYrp
nclHr5DZfx5bim9uJ/sm3FXZfFzurJE9a69S3jELBgvwCwczy/D5OR16fxd6/G7A
A4wAAbEv7/CRmfeOm9CK46OGy0hDYWaC7DLj2xDaW79TCKBWIgEyGx8fvWsJYSCS
KPPiYr1KlrjnFgSBlsl82V7OFvhVUZpC4aaWZTScYNXykGiOfPX4hA31C+5tIkCY
RPARus/BgcCsWQ03kcFQmugNoYMqtmYmXXyLtBkblLV3XiPsbW3MhTkBjwlKsRRz
jKrwSrHYYhCrCHwvle72lCA+rvF5oZ2W68PxFWxylmNt4B2Oy+Aq1mJ6gMOnQ2pv
O7mryQbirfAp7xwE3lWaWPylGAfFKg1rt+i+eX63lWLKhfdxPgg3kDe9GN2EDGWM
eXPWuHP3/jHUFiZHYRYo1Dtn2lj5/koQ+KX2FULVJk44BB5+3knhVtm1tge1hML0
yPkBJ6kQZtIE8L1sHph5U71+FcXzUkBAa8vts+zfFwZLbXButo5TAUHmFxL/6k0L
9Vt0Os0cCuz25T6nA+urZpKcQe1dR9KxgJPJC7cKR577rK/MvviyioP5u0OJKdbU
OFDj3e5+kjQ027dSKvRb8AN25CQRPOHvrElLzuDXvUxR7LRVYAOm6DoTaLx8rU9g
dGmGBxqwTAJOpQwZChKiTp+7DQJ3QnovZc2oii8BtwrmmpiJRRUxK9ir06AhkVuB
k8RtZIVLZb2Qt5r5t9znXuQwPjmjIbxVWnVFLQxO6VO5EGrP1wjCyOg7B51GPqyy
BnL/9gVHivt5/tPDz+h7YvuHbAUQryjSvLA2aQYcVLWU4oFQJOYABgqHRooK8U1D
xjMwr53tXv2wKpWrGifFOYk5DohuHW7Mj7NksBihIC3QhSU6E5YxTuo++iOD3ZVu
lBq6b8GiWhkuC8QqbLQvHXeqOeXJV/6zdgrSYMDsWFmBoNJF6vp04ssNoxgKH8P3
Y7yYFsMq1115t3W/ElRVPeWWJhxFKOT6JY0MGThCUKUed0M5h5iY1WdVf/jeN6zH
kMlt8O/SEkxdBZ9y/lLXnVdgBNjopdUb8Mk7WApFK7jbVR7+/cywy2e71qyNEcyG
47tIv+0cD44sv7p4+qvAA5PmDKoacfjsw6FXh+uX7BCuVbwAl85OL0X2B0dIid/g
QZz8ITN3dINMsQSzTYyCikTnJRJhhL+LGi754gqmk8WAqGoqOOvejV/+Jc59e1pu
Q9KRLZ23Zj1nggQVfgO9ZMxQqDz5B5LwmFdI9GLWWT4wph3wk+zVxGni4NIAIFrD
GvU6EzyWpXZBYuQ4elFKNOV3cgBBzRsTURVzGV8t9R/tuA3LPPSZaxiwpunPwWPE
JvBV7CBvxIyYvehA015X0vIhmvrPTRX1I2BQUSAsfLm/d7ssYP239cE10RC8LzDa
qdrZTLMjTNh3/K6PJMRiP2aQO/PYyhX+K+FRn6x98duQfakG0B+yr+4IFFMh2xF0
X81tCPa/R8pDTvvlMjSHB0pVvOWPGmQ1BGpfBktEV70Gz10VuWpv4+WrZW0pOu8B
3atAaudv72tjUkYExKJxXbSQSE1anqxSTZR3/tpoG8ekz30cVZYKzupXJxq74a1Q
RyTlI/Z+I0scl5Zo/AZjkPVpY/iG9FowE4tZ4nVompUDpMZpRxLvRbPdB6FMVxBE
eVlhDKzYBGV+0ZTQZ4xvgEP9CeA15la7tr8H4fczqyyU1zFpp4yUUlV07tua3P65
mB9moJItoNIC9uuOjitXGoZpZTtQom3FaquGSo19m0+fZycfOd12D4sDKhfZLIBM
HUYXaJi6CoHZaRt1OBzUzJrzgZMBqQ+dAoXCRIxj5mZhG/OnEKzFNUMeof0LfWEb
Iot6FjssFqenTuOccBNz5BTOmj0Z/pM6AnHOHgWnhwPbekvflLRCzy51p8wXf51Q
/3uCsyqtEfUvpnujgxByCznRldPnWqZIwu0LoQMvUCsJVFge8HAgHKI8Q372jnbN
/2MPMjzoGv60U6xYlhhkwGGKl0a6eZVcru+qTdl3aqULXw5VsiSELnzbpUkJAZzD
AHXL4OiiOFeJHAoj9qHrcXmb5ws9cdd3uqgq9IhlAeJ3JRUdcnqD8IzFOapNRhbl
fWaHR5l9zPPMqW/hJYDbl5/DHCy+cOIHggGOSY15K2qV9HmD7WLj3yjRwTs+Bhti
vnGb5XbZ+qBSOV+F5Pw/ggVR4MPoumQvs9C/gnkK6i9ECcj/Alxs1H54gKmiBEup
B6mtfjzMzTP9YaXEwx9kflvqiUWZANz4g+NbtRuFp46NTPEJqtZdy4gAkdNcVy25
w2cqhiKsUnHe1JIUGG6JNuWNUuoZ+tU7rsJpYdoJZ3A1xaHwdg6x/dcmPgHzionn
LzRZErbNocG9BFeXNvNIOeTA1Mx136gJsPvBJz5QlJVsIPLnjbVoi8jWhYE5GgS7
z9sopcHIU3fJncyyJivkzbpB/nPBpll1rcgXR8tI3sMXrOlRoEj4ACpuJZ8MFU3I
KjL26jLflkwIMQaFtQXIVlqSriqCGophhaNkH7KaASwhGZQ/M1B2p3dy6mRMEp+8
K2uUEbphcRn9AtMv0TqfOz9hmPcLejUMPsfs3+rgwdWYzd5v5JdZEHpfHRJa4uxh
5EDEfks3852RvrVLQQQyac6k2Vs9K7Jd7Vc4eUtendcCEbpOrmcXLVVCw65mN3qf
aId0CxRfiiC1em+ifQda972XsMTQjyyaNxYt79Qf6teKkRz0oBIRaaU2JQXWgHuy
r1o+21hMq4XuAacnTWXIxtFeBU4/lpT5F3dq2tYuM2ZB/HW0iLakWGm4WmQsmmX4
oiUFGPLDGavIOrToFWtw4m5UOmIspuyug0hCPP3E10FSD8kbXziLW/2UbUXeClWR
7TAvyB6QGs2H9eDPcsDaUhSCTkokdPDFKrfluCNau8qTxN7eDiN2Gh1NcAv7bH42
eijhRMbvHihiDIPvk8+F2rV4tCfN2laDeQ3LO04hQOPLcNIMnLqlx88mfbX2Cj5a
V27uIxJuWgHO7YZuK423yx8S/hIvM9WHoQ0zMxo547rVZ0Ga8Uwqp4WSNGj3ca+i
Oz4tFfKz21etYfsHN3qqf+BPZvTK1BC0JhpVAIiHmxefguMchxV2YUjhHPC2Z11V
gPIE7jqTzUiv4PiapBEE9zBFqal+3H2nTPqZIM2iFJ4v4IKUPA2FfNRd8t1hE4Zc
LkSfZ295Z8XtdwqDK53twEKaJn/RC6whDznn1htamPwwoECReLLPl8JPuLzb4NTz
qQ7QoVawHPdXLUSoGv6bL7zsJ1f6EzSi+Xl61b+kNTyQxvuBtVh1m01E3QkoOWjX
VPf4n5mxq+RqotVnObFyTJcKpo266uLUXg6e3oWUCQNAxAwhIl8Mh7hXxyjHNF9M
wcfyd09IkqY7OJuKsO0PrJ+WkZpchN6ZcCrZGhDDaip6a0eg6fHZBofraffok6Ho
6+BvLPpqRIuvQOSY97I/KqqWcAWAeQUMK897TCPCZT5WKt7V6BlHCqRCjCo7dbqY
bE7Sr1TlaeiJ3Wm1N2jKcELkdWaRz84J+51mEDNNG+SUFbgBolohJmQy6y1vIH6B
kWutNckd+fVajl1rjol0zHxJCrzIkkn+L9gadiVl3KL7KQANyGmkX8UjoTcodzCx
4bMspEhzsZIfhX1051yezTQdzlL0l1q4nnhG1ZKogA0T2jI3PUFIhXIpRz9ELoJk
pijs9ooAwA1ioH3Ti2hdaBWEZE9XalXWnhk4zv2yR4Zb2YY4X8GBsxVAHe5HYgWH
xPmmRCKvUdARrKNeV1/wpnf2NW+ijcZ219v+ZdtO6vsnlxpw/aHLVywyNpppyqrp
rIyKkbjkvEut8iCyRBX1a9hTjpLnsw+Bfo9p5AlvEKuAKy4nqivxz1l4do1eWsjo
NFPvyOdIWkT8yK/MYdZqlmOA1HtBQD19sYnM0Q9HlrGwhwS+bMeSjleQx+RLZFmP
QbJ7yhZW/z3dYa3wqOrrVWb+l5POSj6z+ocL5KmrNquq6VPZZtL9TjRiIclNQLLA
q5iCDdQeFb0RBXvnsgX0NQMJ3pjOFcGnEPtz6fU7PnMgKVZ3/aZU/9O1MU2bQmPa
FdKaeKaXxOPhAm6oguYCD/tgESU6xXwAsBHfaZwlMPrIpf4y5iiE5HI8czGerFOb
SpfSG0CDs/290+2eBJUL3UMwQdWhwU/QUP6Nk1zEDamuzmSLe6KYruFEfjuL5C88
l6yoJggdkGI0g8S9H7e9Gp9BjByd2dnjVZJzYTXvRmCD6OsbZL9Hi05cvupOy5Rx
MiSrQROeYpBq599j1V9doNxea/YYZ7WE9H1TidAcOsyFD3/N8RqnihlxfQGDm9gs
LTRhdpKowW52HC8SoNzvNit6b7qUSgALLMyKXBTrSuSwdQdsBoHs6bS62Qojm//E
UdTt7pmOOQc8f+A5j7VL+qBlYalI2mDCQKRL286XfbmwGdDhY6paL0+DibZ7LEf7
Og1sJe2cjP3Rhc/UC/5L5NqPb4tuyJPvbOcUapQJoP5WtMgjZ/6GFXVlEyl16Ijp
D8+amP4Plb4C+GxvdlkCyWlyaij+WNvsSy4SiwOR+3d3UZ0dHk7o2S9t3937xSCu
9nIaRtJ2ehgHiC8AHjSjt4VgbIpWCfWBjo7WQM7Mqgguuj7sCamqh5x34+d9zjwb
JIWcMgrHxJitf8nuZAOPoGDCGt/FN/DyT4LteKUxD7BhbUl9XFvUsN9b78iXNyCK
yqUeBqDPqP1k2M9SrRlk26SAVJ+8m85psFx1j4skP8BlamlNV9wKShhvi1HncOCU
X2q41xVzBz84MTGKdWf3B/c5rHhDsqwpZyNOyMz0yWDR4BMxLHcgHKoA+/RbW4yi
ebzhUU8Nni69SeFno36M0ByQ5SVv5lY1A7UrhAzN4LcNmUobjh9ZypJOnAA667MD
HPWFY6+y4/lPMs0FMzjeyBJZ6yRj0uGfBlXxzJ82tJFSXqb/VTxqwCxDPotxMlcL
sE/ssBYugrv8YcjbgNOf9ZIM+nXDlgLn3wUScx0JU3u0KVOUaZBywANMaDlqmfcK
PA1AixIPIkkudCh+Ka5KTf6ppQoFiMz+buNdrDaOFe5KUF4MRbiJrOo6s+xu5mil
4bq4zVdp0SiCb4z9M/Iar6sd5BXPJd9jkzktph02/EUI1tYmDP42nnDbk7l7xIMc
+76heQCdHv8zFEJ2XmfnaWivLXgENryPcocoJktuxvaMaj3yGTJ3q0dgo0LQr0kp
ng5WkqmRtAIKe2lUx2gq7UlQ+DQhsc+RIY6JK1aDa3xihBobffXmG7orqjPOqw0x
f9UxCHjAUwxp2lvLlgquYqk2q2iOFrAUmphh5/neaM4HzTAtTVFwEyr7y13n+RIb
wkFsXLNNitjqktocbf4w78R1m+X7SEWpxl44zIrvNaCQjOvPjS9FRuNPx8Utvb0w
f6oQNjpZ3BcWooKpFXIn0gXW4x6Y3MHtWXrke/lDEXYOeFyLelUCDzOKQQNCJlKY
RAevqNCFCsX264EDyDWZYC9MD5qAMrb5fwxrPymusn2v5q5S6yhVvH45fuIsZsZu
yznuIqJK9XCmLeT5aECSaNRJDAY9hD2d8XBFMbwaX97wgslbTjjHWDCCY1+yT0aa
T5jzfJYR3Ygswvjpz/q+YKfnsLxRubDZ5qLuwuZCHGqksOyuiXoyISIfM6/6DvLo
DRiEeTNc8szXq/0RzNmYgEhTqWSh7N1FRC3koH+y7xOBFnyOj4VApFoaNJRuLCfe
IrY2vxn3aDCm6aBFrIxd3YGFIGvbhOdsUoHG913UdrOTK2RFayd0edt7mX0Hh9Kb
NyLb3WvSgD6hLAk46P+0e6DOap17YmauR52wCJqglSTEo5XOY/ah0y0QWmhPeuGM
NT3kHrdf+ZLlH27x/ZtAmOpwf1vw26nLPYf+kD6fvHRSrXcijR0oesWeXNTvdrVr
f33bbIEqeiMpZ0TwLJUzEC+NM/w3LiwKWMlNEkD5dwhOiuZGj28io+Obi3m6WOlP
ale9ieIxp2Q1J6QwWDlfTik4PeTgUeOnY+M9Upn08+EmEZlzr394Q0BDSzT1QmaX
CIwRHZTfH99whejjSLUBObdu1V+xJ65Z82cSBsybwFIdC6ol2eBbQ00ShuezpnSx
yIuZWD2WLPY88qK5E7XemmM4z7Lvpx1w+9rrQuuDTlLoT48f+xJMw2CFsK2D1OxH
eBjzI0LfAwsl4l/uBmY7YHnBUzyDH2uAH+ATARRBVWn7rliNOQnV5AeB9koAQDnA
beZ0nUkGM5McX7BuUY03fY2eDaTt0+cJlxBcnJqZ2Ih4daEuTAtl3tram3w2rufH
uudiInRS3G5smrBrl39TL618EXWCNZp9e4r24iqRiKAIi92/4hFIHsJJcNnRvEiz
8EFFo29qs5i57PfVwgqBAy6/Jr8LGjSsRncprm8s7p3pzr1rdhbh/HN9GhuKiKzr
efMjRKMvF7OzKc6hT7Svoi9HkNWQgl97Ny5X0qNW68NW5lE5wADT1s78dEPUqCpw
gpfvKxHwVQOIAhvoG3j77G8Oymmr3NhxG9H6skb7ICsvtndBkADPGuROXwmkbQzL
TI2UCbnYo5uv0x1AuvjK88a7rYGY3sApmsNasr58WCVzw1aev/7wR1qiRAfHdKgx
7Ok+fQ7cOFlxV7V7nIIeHJXZKkab6CYCFWSxEfyTbi7lLSgs0uoV1rzxNUcMKE4+
jJ2RQ3hdrd0uz7EAXkwEH1nNDunkwPEEeSePinmyvX2gfzMFwsp092TBxUhCLM8x
jaRXBXYEoP97A6AnEs8/jxAhML9nT7TK4UTsDZwz7G2DzoXTBQl5rmTBjt/lDuVo
JcOzQt+ErQ3xk1Qtb0povym0lQQam4P7998xuwDmOOKr/bCGqoPaCp1Ik6fmLabT
uFWmaQZx976ruV8AQpjgUd1f3aWWWgMrhKl3iUdwCTgplfbCUOJynGij8g8Lm++S
gR0po91covdrD06mIt+Vml5rnWJpGJxYgdZAQFkiInQOhcLeLy6R69n+ixDfR0ai
TcjVVUl7/TMrY8aRb+J5mQOgqtdBBY9J0cXyMQOVxks3rCWSDRJGRvLHOY4c5rtY
HYL9oh4m3oWmOXIN2aIaHvFPKdO6kQGywlgz3eInQ7vbkR/36mkDtlPstkXn+Pgk
qUdUWaX+FfsZAbmxbcMFPmAYYYB7T4aMpQp63DUSHguQbXcX4ixsqyG4da5WNnU4
wV8VJy20ULrpw7j67BhP9b71fpPknd04/nvD4lRtTooa6K9pq7/5xHWGws5dxVll
1I2c8qrTDNwyUQ9p8DXcEGiK4pHzuE4I/Tc5UbkDcMN3OZo6k80l6544iEZuTitp
TvxvG7EKZH4Eb0YjCXFch67Tdad+0ZoT25n6nVrRjWbR0CwCRBovWembBqfz3xll
XoBSHKCOWGhU7w9VsN0dP1nNaImkfDgBsoU69jQ/BZVysp+ktuaAKMUGlbQSY/kA
XEx/d9iNvPOjyAuGR2RF6zuoksF71l86IMvY/duynRWlTstCy0zeOfndzbqNLRHf
4LgfxCK3TlLiSDtZrhEQp1HyKEAPIdxfUCzHY+tN/HBAjV3r1+WCJIvhBiMKiPAK
3+Ki7SX4QFqc/r+fB5Zlsm5ORcZQh9ckhF+WuhkmLmUhGF7BbkquchLWwaZfunO9
xB34Lpml05vMWtZt+08vu9R2QxjCmmzvBOM41j5p9acPn8nqABuguR72mVH5L8SN
tLM9OZJpAExlA/m10foQ3rocYB1g1/LqPchjXyqyIqHf0aR2TgO+QIrr8xTtmB1B
3Qio3CcVkNQczehocbrwuD+LsES4gDGESVeWdu2hK1jjy0SyZbPxRvxqTp8VdaiN
Wl/czBTYwh3jsUuXG5tPu1cMC1dd1sm1jCHGP3Shi1j1YGaqEs63A1sjiFLmYX72
vL/MjJBjAUoSG5VSt4ePUUbAcGNlAbjhJcn9iReSfRCtIWrnFlmy/6tPzeO4kcKT
YtatpqO+VTbCNCoQE6ZbM/qYfij0vaih/Hgysyh6W6sosZATDRVVtMZQCJBrv2ub
8j9z8qRyJTqrcYQPcgO6f5ZHHkeYRUSn1wpK+Vt610NLJfFEislbyTM22ZCKnGNw
XAOw6T/G2MSsjtbWYJYNP0RhTKznSg11zjqMQMPJQxbxh3E+JrtBNYZiFrBqtyP8
0THBf+Y8Nnv+d6f0fMMtwu72wu2Hw1wUJn/RQT6JxfIVkxOTccffMf//1VFuIRfQ
o6Mx0N64sdkvcNQ9DV3uRntpIkYa6SvjhOYYi/eTmk/qSIFzd15gEBP5nmEsQ8s6
JE/YgHeKzLCQqvBtwZHhL1BLbFgNRJPJDvXAJw82OrfWsbu5ZW1DOGKCFjq40yI7
wi6nK0fiDKJSirgvinswusz6LaGObUOd6s7epOPMcx8ZkSH957ptTPj2jYFovXrw
HWJc0xx69Ki4/Vf3J5Z7x/1pnnVM3npmnvVV+kiN5BpTuo5mkU/aJHqdX3fGRI+n
4LKQ9U9xfVoEfLPn1np7mseDxUsnKOwyhAgowe0scHDg7lrJZMWJGDzaT0ceAqVO
JGSsvPxeyo5L2i0feHpywMkXy4hiD6ikVPPHhUlrFcx4bleCDLWbZglbE0d/2oAF
o0tqcTAzukXyLXTUWLeHY0q06u+gvHZu60BuztWsSmn65w/EAF+VykMPeWHvAHcM
exFnUPL6V5cV0nhe5H62jI2wEN2YKnyYQgVfB/xgzVZNwG5MISpxGvTe1uriC++c
18JdZSIrFrJQmGcpw/TZK58CYUuxSQuGJuO7GzOsOMlGu5wTNMNgaOil/PzfHfJE
ERPq1E5yY+Uj6eyg6BAbCdSKXJa5KXoVcxYmvYF+BZMKggnmsYw+ibW+rRrpULw5
Cv7NRFY37up8xt56BP2TxhKZmUOc9j7c7hHyKXA/mJKammYZmfi/gKhxkIcBaytM
Vp8wKfs6iXglTkSkOw+pzYh5qwAZ7BGShEXV3TmxjbXI41hxcEGas/S0djckpCCs
HOeb4MRX+KsFsiQ2lmI1DUq2CUCmzaefczEoa78zPfRI6G8dRPhpjYk3upEHW6IQ
3ppR3BGKfJudE11UbtEF0RcJtWGPDPSiy3zfd8WU+QrpkNvU7D4zoATm8B88tUvK
bAswzKLrmTw07vZt/H5ffNwRgbAiBvgAYHPj6VbmqbxD52bN/E4IDWkmwnGAOHhb
dc0m4mx2GnZOrZAVcXhWJGoV29ix/QYgboik99eAY+QM4qFQILKBuKsrWa1c5HmI
LBparh9TGdVfKpHW3g7LYFxwVnDZS/pOWsfN+HBT7NKH7GLKOb0mCbPDqjX9vsh+
inivFYzU8BAM8xx8qhcbiCcbvuYIT4l6It9peZYuozQwNskpFm8mYfZVey9FGb+3
zvs4lNpfDoSdU33zWI2N487KJfFt8HK5VMmuSm7CPcDfBQdZ7QLlTflco3BAajMj
eOACgaCyvJBfr5G2uvxy7SPKmsZs9AzI0FWFW+WZ9PULlV771hHQNftsrmO0VLY9
zT7TC/+6EvrfGEgtloXn+vd9ti5J38X/DX1jr8j2kkCFa7vdclMEA0u9e4VKz58m
NvWBgOS0hLtn7hb3m8unNsqS+pF9Xj9frT87dSYhWlB4+Nszj16BYUN98jNsesJq
JpAlSkma6MiJX8v47MwY1xqj2hU2F1DrKCu5VwLusXp3cpZEADfrvKFa2IQ37NDS
uE4LKmUUoIfSYTtu/MFYfzKkkc9DDlKDaRTv/X+7+gMGNx1V5zddeDzeWwiuounI
sTiNZEqRU5/i6LTLmJoeU78lVCmKe8RyDcBjuBwZt8ZPNGoSRuPDfeVe/njzTYuF
TmNvG7XTB7qNBEG04UbTEsOeULK4q/26vVLsPsRzfTxdxBW4zJmKA3LRMu5jopps
U6ZmQhWsMrJ1bA/6Q4ngZ/DVrumIw7Rw4Ndi9CTDGgD49F/NvRWwXcMK5r7unWYV
9P6PSq9HkVQ61+zbrf388oAyJRc7DzD8RE9PbSHLV4u/5v+MmJJYVuPB2mSLC8jk
0qZdMXyTqkakp/g+gJs5PQsvgbRgHA0eMgnvmbtYzUgqwTi+waGwarbkgYl69NWt
/Ydfq4uer+JdImbCawZG6oY2EXM20IvD0eaVr2OIdEXAr6Fho/rl3F0PogFs1e4R
fUoBy70EG9yoBSaNXG0fTiaKiYCAyku8vv+3jyznIAoRJ+i5uTvXi2YYMpXzMAS0
VY0jgxngnGlHKjLzpwLXRrfCZjDA5mwn4g6uB/ScOJas7tgi3cdlGDx6s7PQITnc
cfG7/caNkCIEptxGdVqf3B1uSygBZwSE6omGd7/nH5zkmoxQwIlIN7U0ImEjYAZL
KYjtQJ++ghgIFymh5nxBC9+6Fuh8g8RVu+Gdcl0/qsFFfd7/DRz7PKtdyaMq5HmJ
iB5jLFg56OuF/Qj8FO1q6XJidzx715zLhaCEAz9qAyO/EwJgKTOien9UJFPQjGlu
09DLhJKXMxKtMfk5GL3BF3LMHKx4y6RmOzIh1tl+FZDkULHuKsXJyZK+EUrUH3nm
17+d5zJhFobjEC/JMSsY1y2KlPXM5vzmEqsyC3HjugINllHQ7glyYqsv9RvOVYzl
u5PbDhnec0ny27X695blQPJtcqiUtsaIQK9qFFXMemC/rGND/GBC1Gy2SSaHBFlS
pX65iw36+pIXjpn0mebiouGcND4IA55NVHAJzQ7nHlb5dJ/cTlFfWLTxChziGl8N
n0xVKbff4RfYQeeUQqnwUWYCIdo4k5dDUGd3Ruqh8J7d2XeV+zWdgnXVd3+TGLbk
xRqMfAnfbRLPQfMb+68NTCV2ozmeuL8kFQkJojXlIqQY/jedGtSrGRFmnVrscZM3
A4vjR8rFpXqlniKmpuGkBKaxQOo4s96SsSAMzNRl+JObvSJMIfDar+MUSSyuoM05
729p902qV+oboO8KtTn6SVTYZXyzI9hplgQK1LQ2cVCNOE1zLf0YYy94JuhsI7oA
hP2S38xkEu1FkBfGN+SBXq++xN8iDnOnFBIa9IEBkx+xhBPOlYvltviQ060V+jzB
Vj3EVj7lwYVT93nuzKKYRjezLrYW5ohfmGKIBLlBNmH9u/CFS5UY9FGyDSl1vnb+
Tg48/SCSYlAGl31TIBywp9mNDgHDUR9qbySr3GQdq9Q/CMsoIFw17rkR+oAVOurH
5ewynr/a8SrMfxef6bWpnLlppP8VSEBZUJ8EgLqm3uOvl4P3mU8b/ftu+CrwQFWE
joxxbPAl8zEBLlT9hdFJwr8vZHambp+aDdz7E0t61UsYaR+ymwGJGYQeSt9Ejqtl
QmQO8H8+zvkJFew5CXj8h0C3uGU4lbnH2i/AtOZSXQBueedVDRSdvWA/R1TZk2+6
5+hFjAmNFXYijLUIpTQYHMVP45MMwCv+6SMXTDrPljL0Jsb1xyyax0psFpPOoaq8
9t5cNUEoC5MzHqvSCLbq0CGlqaFHnV4NYuSjoRx1LghrakiWnNOlt9papiCZawD4
R9wEFfwRO+GMgw423MIQANDPwMjCYWNh6pBhWZxiXeperV3bBl1cJg+dYcBKsHfY
sycO/Tn7qmbv/tchRtNVGHogyUppLo+3GhjxO3hYNX2K80hAVk16bdF9qQN8t3/y
sNgcaNTd+hd9djhLRpnwrLesB63RhyK6U57yu3TiJPRwfynRQDld0Y8tIcpqJalm
JYoiE94v6dZ2ccPJ8U3gkQNqCFVOXWp1sr/63cO1jO4+NT8XRYGGt6YyU9Qv0Vfh
AblnCmTj8YjI9oUUktcxa7o1m3wlTsAYeVxmW4wJy4z4F2ay/NCaBlgpzM3ta9PE
+VUfNSjuAtN07AWlUePw9CcgTAVxDCTHvKw2boPkL1iZIITFe3js2/++zWJXbwwj
/zwkfZzG7pFg5lGKHhtbZTKcg1mKOyyOCvEVyQW+eb6Cwk8wQ6apDdxbU1p3a9T1
KmCPTNxB9dM9qRGu+emd1vZILXKH8R3mHr1UlpMP829QlbZCPLA6eOsDui3sZQUm
lwGw1wi7bE/UkX1wRUHaDM1uMSX1Et2d2pm6kHAa7rI9u4LeyDNbG9d1Shl6LePR
wEtkMtUUnNAnFkCytpwZmY+WKd3M5hBMwyLIzkCF8fMyl1rSHCtbxJQu72NPzU8B
kvG92zNkGrPSbTlYAIf1/1+NVkhBX7YTApAVAVGwH7SV5EoeCWUPNMIr5LXLkdj3
gYAEYtEtHWiU5VE2z+Ut6bdaDOiXbxx8zqJK8RvAqP6I/dUa0lw2pW8msp3QOfan
dF/8rBgYOvmdF1acOUxU4X21/zc+OS5baT4Dal+tp42rKdfBzcRWJMrNjWhYdBEV
KTM64t65HAhcMqbdgNsWMwB3m8zziWnWFxXrnlcoQ4sFC3+ddyP00mnua0pV98aN
eM/sRYrTS9VQz76tXE7ojVo1mRRi7yuBd/Qd20/cWxtAL+6fhFNsh5yVOy39ZWCs
BdmaXvvfOAYlcu+U8XLSRkt91HmQWU5MB9wat1RDp4XacwtDPaBwbhtK/mLVibqc
JcucTXZrUx+lHkOKFb3d9OR1HyM3PmdVxm/Z28hf0g3pHMF16DOyrmbUcdbtVEFb
1EW15Z+kFRmNMgGtDaf+K2dI1TbXhq76x00HPcMrzxNUTMi+pZqJL9y3F/lBCPLr
NfU+0BAMutYxiNDSWlL2AojeMcVS5TlrAkFRr5Bmtu4NXPYEeSjBW2D/OJJds5zI
CIRoBoUq0cqVKVqNGBqN8jQT9lSWn2W5S57v0hy2dejWriwZy2wFJTfWpdz4QXWD
d501f0EGivNVqBpz6NIQL4+dGdgazrw06w0v4AP0gL2iDyK7ygBEGykaCeRcqslb
63FsaNXzdBLrYKo6FKzCwSKwUm1PXKyHlFP9tpQNbg/FIA3/+nkMihUteIoNIl9u
p+R6aR4m8mnn0CwDrrKjFWdjE2tVVIau+CU25K+6HQVmr26Pyh4ZkbwcWZP6EhNW
UTiTXVA75Is4zOunfa+ZkbzzGuMRIemqUN64Ibho4YcmGiBYU46LESt21YeAruEK
UE0xlQIBwujOrq7CdAYcbSws6ZV9ND0Fb2/wmddrdIKQAtjgtvJfML5q5JpNgsjQ
XfPMwIRQ7Yadb+GN/+H5MSm5mmaTysxQmO2IEoqfz5xCbXENX2D1jrdy6/5zsSCR
Pr3o8gDnFbAebdWfexh23VqcEEiyQqWiaQ6RIayK8CCDsl80pH/b8BdpcDErxW/i
dz7qLWzZLdi1q2C34/C016jImrUH8pEUr7x7TblPN+PgqTGdnMeJYtbZZGOAnJBw
7z16+/S9ABz9OfZfmC1+awutIhDVJtMHDPWeHFo1dgYCejF+SoP3dZ1D7SnxiM9q
zfNm47V57jUUJkIXlif0PMFr1CNo9XpD526k58Lyny80YSWkBb7yLJigOEyTjg21
A3xkN6eKJ3VSthH3GjWK8EDVKbpVZ9Kr3Bj46876cmmkJHY8gmrzoP41B1Q9aTuo
Fl4jY5aeBUKuJWJ++MIRYM2AYtFMPFa2P6+ui6diPhGMaZoDLYYTA2A7mJ9LJVnF
9t/bWM2JzVvi2/wrOXhBvVA2HdKsscxX+Er7K64xHI3HfOKy2G7NYutri7YGl8l9
f/tibMtHZVuhdM5NVyz3W0A7rAXDbk1ZnFtOWBpXja5PZaISbkF/GiFRlgJIkCw/
+lowVkR+X2ex+i++Cva9/sdVukjQ2q2OJsg8cH4yt70hZCK6FezPjDTgoBX5UuK/
+UPQxawRVmTX/T44sHDxaIIG9fknI1vwcQjSqEaf0Fu3UxC0ncRDpj5GSXzgzfPK
gZtqvRvxewM+uYO3I97gS0bE+ODMOm3PZneDpCxFfo7QeHhwcnWfqrqd20jCTVuI
JeKfUQ6OjOBbiMA24EbK1c7eoy1yfSllGAVRV48sgNaiYXkWXox65vPalJZuI5e7
itfkeH8WSfXOxepxLPNAuGzwm9OEcl2q3oMKzorH6dQWKaMv8LO9a9okDHwx5/Gm
ltoweNVUuqffHg6woiR7Qb1BlLiVPd/NaqxC7I59UVc+Xyti1n7cRt1kHVS2TXab
dWVwX7hETpBzCY+F/Xz/x8r94sba8qVfB2HTxq+78N3LtkUubkXPY4/la51Ux6F0
VRrTEsDv8RYfw/JUKZi+JJeO6HMHSXfifXkgOxt+4ESm1gv2EtKBTfC2YN4yg4ys
kZhZAoEuW2BYb6Cy7c8oAY0PAlVTGZ2/Pwb8fzLsIZO3hsBDR7O3WzhnAUKHFyd0
5mJghD7qqguMCh02Af95hlopsQVIZNn099l3KNbxoe3M8eoiXdeX4kvAXDj6CPPl
ZvqP02fGfPMxehXBRVYtPqTcXS69n7MKqKX3B9Q02YU/teVyK8dalbfs78stR8Y9
7tU1oMe+F8li2syHA+7p4Nuhp+lVJWYxjRwfQqHha/UVlPSdnYeqRg1v+szqNWdI
PMX2awyAF1YdGnK+PCp8WSd9WJBUz6MrB+4yVmMA0I1E4r4mL4mhCeXrSScaqxAs
VU2xv3h8ZGgiqL27v5UkKtoGMfoKugi5fAZTS+dQ2jwIdbGkgSco34cFQGeOPRHz
NzzPa4B/pk2Ral7lrR24O1DUQJVkXDLZVgPuDCNZDGFZGZ53ggHU1+q5RwZaLXNc
VvsS0nJ+Zrxq6k9JdCBu1zA7sIvRAuwRT+PFatQUXAabYxDQIMlFW81xIpJRWujO
DrcS+F3yjxlXFpLQcel3ClBrvraPDjirWNrTzfbMIx+nYrtl1/92j5NyNPioEnag
+yN7S8z9D7E66H8Lznb/IU9JMX/BST2cdaSVURi/7kC0seoWBV1IWKe2MeGEDQSj
Bp/7SOM1z5nLkg3pAXvm1XH2kGPM7qcUWMXpoqL3gZGJqEuddotEKzbZrkSH8oU+
Q2oc93jt0LMJAmeo7aV62IzQHJaPWvtRr0RbiJlM1MkVHCtHuNCS7jATgKQZc7bz
Ygq+yLnhZ3bdo+sGM8N8O8M8v8fx8Mf6eRw/Fa6DEXb9kuUUMwNil3IELGuEMcQd
J8UQvEGlwzsXuPW4I2j6L4sS4E4QueFJFtovMY82ANneprDyYb52nTobusvGQ62X
ie07/gvDt3JktchgKEzQF6jalksYrCI84AsxrIloG+6p7xD91SEfvXEde6ibfDk8
g428h2YVugVHsFa0lExwxMYRMmIOtIhRY4bTXZKKGLN8TPzLPX3TjIRMXRuwHxV6
4/PS+xAkJz9+vLh0nw1YrDij6xVFOBBJOL8/lls+RzAQLKxCw+wYb7l9oXCaYWSW
6gP7H+5FivXv+wcZrYsg7pEU8Xg00d04139L8ZPfqpql7puTbCVfphhQc6kLYKLP
hLrSlSEiAOoUNDupc3M7+RwAImijqPwX+TGu71ALdIUTjHfAR3lfX0GIgZ/hXaxk
WIFy0p/gdk/Gi/FXIWWO/I2+eM8OySG0HXSX0wNxXbuBEaDvSvJTNJJcyPHBULOF
Jo0Q3RrFYWKdq3Tg2Tnb6W10nKG89OEF/wTDW8tEjcUvUfxtV+sFwWm+JSfQUSAJ
QTD1YsMvHHkzC74gpoLxOZyM2hjSVPAV6Byf2ZrX+F+si3KjjRnhpE0F57t1c1mT
JChglU3Pgf8LAAL9ZegRqF24VVvoKGnAiSFqayO7k12kBnmpyjvw9If5f3qWZByU
Frfb6xRNI8F5Hx8gor2t0Em3K8CIw5Za/CasIWrGcp3NUTnGv4/reB48L+EaTjG+
pYUF/PnrxjLOpRsgm00OR5EDd4P2LiEoqtrJVWeCWaAIZm5PsHNhMCLls7po0Lqk
mRv2RkrslhvJ2vCzi/N5pS4dnQyAkRcAMjxIEcIug4DRkD00xDaK+d7bA/73Dwn+
1JF57rfovxgQ08GrYI7pmXcc8qiWNEn19kVXgY3NKlauJRry88/W4oIfLH18FEwO
yydHrhgfDuqPdT3izGd5EnLoJOZ3Fsz9gRYR4pTyOBfJPn3cXmVoCEBdbcSg8szg
/5PgibRrr7n4vuyythQ+cicgQHVr0pYOVyGcvEJQz8W9iTjlWYiYQ+C0nGRsoM+L
TFZ+lMKg+vLzYHbQ5J51kzGj4raSf9zeqMvUNFVNywi5qrFlQsTuPoLv6QMoygSb
xxDm8bltg2/Q7H0NXGZmi4TSm70/qusJptDz2SjUtGDdR67VySCZe3JIi+CpET9E
Ch4BLGSjAzTkvj4sRbZhM9+1GMb57e1BXMRv+qCzDMp+9SLPreDOuTyejU1JhqBo
H6RvYL/bDO6Z3I6cGWQZMgOxmP4D8is0YuRM/pNnOgn4N5/fVISN95g3Rku60/YO
gOm9J7QWIN6fT3KeuwHntwSpaPWNFxq1FeXcR1bt+j10zgaQx4PSPNcUOiHkktNW
nJA9gJoFwg3fOURNPbAtNWUkSyiu/4Z5eKyXH/HjrGVP1nE3V7m26vTCR/nP02mJ
Br9L8NyWzrqyTrqUtfdGyo4PsMzHAx9MW++8Q2kIIvcziran4AZ+dYPVmzs34lbE
+rCa7mZMoSvDU3AidukeGU7DfHYIN/8hxMD1gmCiFXI2qM3JYXXWd3vZDsqTDDnk
hyF3WjjzxIDLCc75feBo3yw5nazG0FgT+ICFZ4ZHnvrT3w53gLXjd6VkW0dMXwEc
WfUzptnhtfDxhilC8rqLkEdCNX1sznxL5ilmuC6J2NZXvwpdkK/fkRyZUOomKVZW
RAh2WnT9vqIUCP5ehH8tsCij9dxfFkyvF+rcyFLPF0k3QVjbNbRuEDk3noGol2Or
K5VB3kr3DBWwLfKDmZMftUgUwquX2Bgp2dc5eBFGlBUnBlrxvLDUtWBB7HUeRqyX
PYwhcpIsqStNHM2F5tWmiaTdL801eKTR6Rh9UXZ4edYeYb4/0+77fAGtyfHrdf7w
bpP/sWO2kz7RX5KU2jRskPQpCTR4VaqyEvAZITcNU7qi3EiX5qGXHq0RJ6CQvErz
S6AQTekkWRKIN1enLmE8iHIWoMOU669fAXGPcfZKyHoFkEyERgxJQur8AzJ5ycqJ
mB3MjKIMcx2C8qAGHPAvHhnUdwaZETzh0sazRRpzEd7GwVmZc4Hx928se9ecRk3j
QJkxfJUsewEJVZ+F+glVlzKgrNDARY1IBXuVeIcv3rzqI366ojODDLQug85Xm7he
dqE2tXbOLbShOrXROkIN4JL39bHqdfz7OiduVb89KmdSZ0oSnRPcsdTCRVjCYOOt
PzfcZIecK3gxHlfnK0j5W8q1zx5CsGts9oTHgpZkHQO4XlaWvj6mGd4kejhZimeW
ScjvLy+5HHKt5NXXcUonbC2r2AxUcCuCHfCk/jLtC8b2x52pZVu65WW4YUkLD8g6
5D6bOEkR42UD9kj1uV1mEeaD7IDzDncReffW2NPG7MEWCMZTTplbNKD9fzyBF7nC
ee1nNHRpPtHnJV1Al2HShMN5ck7S7Yw8HKIOVa3JELOr5WyFHeVUvxXaKGvsWQwm
eYROPyb3hDdWo3LsZ6pLIccLHCz++pTFAHMshBkDDGEcA1hWtfpncdtUyhO+CnT1
+XhoDiOAh16bnjZ8xV2KKaKjOP9kZFpcaJhY9L+42HyDl2N2qdm0RgysRYMXx+7V
VhImLnpqD6+Fi13Qe8zVQKJjn12MrHtaftfl4VBugeeUpxfbfL6GTfzXDSL1SMFJ
IrZVhqU4HpdFq6cbJwnErArtG4F8riqHqJzSwkmVgjan+ENcXz4lWjgGMfKlbdT+
WmXmd2mPTQEA4ZDmReP36BvVKOq03Love0W+9Bsd6HC1M4kyjnDugBcpdb2eYntP
ST4Rco1S0mIcpuTrgpqfQoodMP0Iml3JfQW4wGubBTkP59IIujIgfe9dwOYEiHVo
OUJZ2fQVdpGoPcnV4Mmi5d0Xp8MAis0UDCfA7K7vvWhml8MsMpyvnfyElllIlPTb
wAtgBDlNXDSHBT1pjUwlZtJh0Xk0U9LjKLc7Vg/lHH9sRgJ4UNfpkwtZvqUxxnNW
6uqQq2c2Ng4IdFKEomwjyCbt1W2FXsyp65t6pbdO+x/YjjowrjCSLchT/tytSozR
Fk3kHtHjY6jjOMmCT++/A7/aM3MjzFY/jLte20NrayRUb8lzmnr4mBpw/01kNpZh
qyDt6eVYIKxa1tbWmOEB5iewEV+/nTyoytgylWld4ODilg6oeWps9XaWFFbAJM2d
cdeRhYiu1Dj5ZH9JNHDL6z1Sngxdzw7ojUtSK+yXEFdXUcDvrxv1rnPbykSS0M4Q
U9YBjNXyxfCnFbDXLgKNyzOztEUrKVhqHybQ9762aXW76J8GQvpujzrrukgvV88+
0hCH2L91C7L3EBjXDgEOaeFJ005uH07glwvpQQxVNFJn93Onc25X7MXJcCrQ1e4C
HZjca9/oCGI/jqF3VSAC7ex1vWPfSBVJB1rA50ktHrdy65l3pCFlBji9BHzEh16a
sj0bsIG76LZGNjJ+dNy9y1/jHgpbffOduatu7kJ4z2DCoFS2eQjZKkmq/Gsdk99V
eO/mQiJk86+PwLunM+X2iB6OTjSgdLGB6+b2K//3F221frnvtddMvx6h/6LSJaeG
f8+2akxpC47cxBa5NiJdLxWs3VJHJTsVYMr+ZYERCDuS0a+OJlaRfDn3lZyxBqiC
gJXHWSSUnFsIN8O1V9acwxvoSz3MUR1qRNePIFqxVDkoL/iVE6a+wONLDVNxNBwC
CpkWapOHv33TUaZkqfXlzsJgMyYDFLkRrCnw891loOpRSXKcJLVWoBiFfP2M/Iad
H3Xo44yoou9o9+Vfsw2mxsPJ5/ZLyQP/ZR5Zz8y/rru6XmEQhBWjXAfo3rwwSzHY
56h+dh1qF0VGViPy27IU/n8M7H1iXjKk6r5vYbHe3CbVOJdL1WeA8ci86gh+78Ab
rDiS3DtLH8sQ2gsNIJ1YYaX/PFREN3CqGYJwYZDPc06PGKHcsjiefskeTSF4VTdX
gL0ICjUd6VMw7qv4EQUPWS8jIMlMwPMoxE8i7t+THKjQF410MutI2nEEV4jSFBvb
mC+fG4yPXuTYaboW0qkjOPwegWo7aSyGsGRWHdAOIfn9CYwAqezN5L6kKZKOoBu8
I1pOaS5z3y92o7xoEjyWmwBeMZT+Aci7KXQ8rl09bfE4JbExMT9wYKats3GTyuiG
VcKClUWMW0iL59S0mxQdSxzqdojdt7sfmGqLuPo1iaU3k8p11EWu+wcSn6jkzIYK
peAau1/loTl3zrTQpy8/fZB4IiwlF3fsVfEvLaMTNs0wTCYWGAUy2oby2PdJVrv8
puwo7Dw76H5Nc/HVtzr21AY7atjZYZJI11NrkX18N754iLKckaitFyye2nONc8qz
nxDiJINhCqF2IBM5o3nvaA/iefQuRJVJMeLHzabBk2LsrgMSs2acPHD8O0WYGkEJ
ToTf6QliUCtEydBiU1/5dmpBAh4hZR5UKFppdLqJ2H3AZIllGtCxB+hj1qHs/amL
Co2jC9bSU0NFP9uhp1pSQfvsr8nUdKEqsK2X83FzVtnxaAyQV+RGLW20ks9tx/p/
zwbj7jxhAh2jQVac9r3rcPOTysInkXQm766gQaHWYHcvnjUAK5b76q7VZuer6dXg
JloJJQ+uN5IqxuVvYg/QHEYtYXBPGIx6aGqWu3Bg6V1MjHvNaYU/hZErmNAWqvLU
mfx86HtMa7CsynVwfIjZ1s81HHxIfhvOjNBirB/EunB52/4ysHwsgqyoha57YWFc
s5uylVlNdLNrT1JpNUmA6l+Cg1OXGMh/zZhXEWVWAwKVLnQd6asC359xnbrCavAP
Mxiy7Y7gohfrbphq9JA2qeiP+6wJTU9HON3p5lYuWxr4vd59bizpbCWLIrQYZ/g3
nOBizeDv/wb9B7MG8s2UsoJp6D0xoOMVP2XeaDEPxCVX+1NHXrsfxxKmV9nfu9le
mfsyKQXvJaMapIYSre++2m5/ytM3Im/ArM538RARNgtt7xvPy/WSvVtIv72/6X+g
98iz4R+NpXoCIkHuOrNabMSWBA1MePPI034b18HKc4v9gAtDhJ69y2PpdyPxU6tp
97oYSj4dwjyZCV2DH0frnhCIwJzPukb8Q/5mGQ5ZTa1Q9iO20Erd+1nDfQ5+XNPA
XxXtdLrQN3qLQ3ujmBkGPs0LxBRuiadY3rIFiYRLeVY+b7WIKFIb7RbtI/k6mF8+
6mcHUmJ0Nw2hCwgFY+5Ly2LI3l5RklY0hBXm6sdSe3EnP/BaYDqOWRqGjrz6AJSN
PLGL1S/GUGGSF8waNhjl0buGEenNzxU+cO5kzto61dpkzjYotEwOS9p/ppsVWUrv
3sxF22rZ6DSD81Ph6MzYXz14kxsBLgjav2Dn+X2AfnPjo2WbTTo+ShLxdSa8e+iU
eSF7Br4duoFwuuS3h4/8QzvkpcO5vpbFGIyatMyJ8nVbwtZtKYpC/3XjeV55f/fD
MDZxWlv8xogEGj1tjuFnMbw1fFUBTXEMNqJUxJX5XqIvxrusSs6vWrq/SSPCa67t
vp51DfqFSdqMrfuUJyOm7E80WO5SrtM3u2ZvYANrOaFPkyRiwktga9yGOMaFSGgB
1CToGUqExodDJWWPhDisfsYXP8nYb1c1wpxPoGC0pFKxNQHmMwKP6elngMGSv4Dd
sP/hESCvN8SMKAs+z7w+p9FXa97eDL25aq50A0ilkgeMFWxHd2Yk7AkTL3WtwyAD
XxYA/kiYanP1GNszrxO3akdaoupmZaPYS3Cz7ZRWXj0EgXyLFHPfAae1vURPWU1Q
59H0EVHt+p5DHPzf+x6p6MjCfUOqv+vdwWFiMvijZdhsvJ3RHd6nqLpXjkAh3+WI
QMcSSnE4C77aesxIFgpfp3H4ZXrpyNRFHZ+UKsAtFeIxRbgf3x8J2SoYDTKzZDAV
DV/mUWJmgd2sQnODllnSheg/pGT0aU2Lvd9ka5E6iaKrKV2yioVgjcohR9oDKVvo
HFI45bMxEdwgAyFpCjVtaYHwjgScJuxqc0bg7cC/OKn/noiTrBEE1oIa2f+lOQks
4OMPvX0ilHqhtUR0kGXrbBaAs3CHaUZrJRg4+XgbNOW9euH2MttaHXVUTm+rhJzv
l8qqiaarZDlKcuqNcdq5KEPl9QAq0c5vKR85K3V7J4VYtsM8dOZe46cPd9k1dNnT
cThvH6JC1PeTZN0Tg2rzJ3I9tr02j6VSCsudLo0MBLnoyLlSjplHjKFOEcCmT7UE
p0jOrrMGRz6+F4gNnlQ1gvT/N+8derQOm0Z0FxOvLWFvejAipX5B2Ik6hgXuq9d4
Hr81++c6HcpJqOe0sBb9RAkIH3IFDzQrpo+TQf6iifzGUnIRHpyUoabWhJJh4hAH
2pJcJ1K/ydW0WPx/xKFDa6sgBV4XmDMYjUz9+NV5MldN1AxfvYRdiJohzRp4x94h
bRs762nLpbbWpbm6a4dWVfwRYKflQtlkGEUJDbD1GXiz3TfNsIV1o9z1l481WaJE
GOo5iDI0Gpo8Ool8BNyp+YEEOwL6L+zCrgR2hZQeo5XoiT1QOAwaXHk4BcL3WTeb
3UZBXkyafKmz5ODz5fcGFnKiYwgP+8j+v2y+KeMc4ZbnvbCVv0jhpL0dw3Z/ssHj
SX0bVWDW6U89hxCtJFr4YArl2NnzRVyH8RrFvdw+sbSCbywfgdUm/pvp1Tj5wkNo
Bg6GlXINrRyuqdO0hEiZuWW/oORASSyVtlC4wcqsu4WNebJ70Ez/gRyuJXTwS/9x
m3sgnfz3ApEv867FlZLR0uBhTQeNv0ZspJC6dQpsVCA/DjbImyXbVJAJIRSMAXeo
8FpzBrrkT+Ln0QV2/UZbzccslZt4fluXPTVksilZ9NxnJjgVA3jVeZUIDXtym4Kg
6FaB6h7E0m9p1ePKQ6IJ55i9Wb7a0O03BXgNF516fOrzzyZZYRxVzjMwKZUdOZ/H
KAgLBa/zBqKfaR3FliN6YB3gKr3nKJtz5oTppTPhGIo0T6ZUQe2vxtRhMqnemNQQ
/tKzqudC49Rqk+rfGv1d4l0gz0QGYxtmAjxMnPbmA/111BRLfDDvmR+IzSbYYEz6
1p2y8Xukou/TgxkQWaDH1DjJSvNiDTvHwsKS7RBdKHf9Tl1ik0Yp33BQloUoT7lb
wetwR/hcezCf8nr5p+Gx52NYdW6BP/K95I+xr/NUUg19csqeK12zYwfo5CcRw+bH
r2TdKXrEAGJYbVCOGdQaSxhCLSLrsWK9hX0I2xqXfi8SovAaMYxsvnCu30TM7aAF
omREymNHK2B8pD4k528J2TSG5OnIKE1+dD75BEEgQ3SLk+P3BENmK6Hr89l6R2Vb
e/0g1CDT+tlWA9UpCCTDzYilEPolXZhWp/Z8iI3YnQKRwSyukdMUtkOV0TM32vD8
uA/XxInXXy8uIDR9nT+70EfaCmq5hLr301Ydyp1sCW6rP742Xk87g0bMOC+hvfHO
kiNuyac866+espB0GS6PWwLRWvvt2VBwfdzPFjMPHOU4FiMSeEyXsm1LUagDhaQ5
oj1UC4V3GvA4sFq1kSPJN84x9iKTDiJOLsSKCPGgRqOvMsItVOKJyPI31MHVtzJY
a3O1011D4Pz2qIx+aTa0MZhwYAH0qxAdge7ShDjHq/LphKyVqosxSf6mAezYfIpt
OWTSfdBbWgKik4m+rNB9XFsQKuMwZy6QXHtf0eSydj7MtxOC2a/JXP7yhtzQqd7r
0sfDkaOFb2i9AddjI72mgS/+ViiqMtJ94LaKGFdpTA4jdZsmyV0RUc+9wo908IzQ
F29B/+MumOyh8Q4mSK57PnlSz4TwmkWAbJ9COHoS2mqh1nlyTaTdW5u2Si8Cz8uc
MVN0J1cELUCae6MGlFNna0wT10IBWmiqu3EYoQpUCLx9yXytgj8w7omlcKaxLrQT
85aQ3tSSa/S1BOPnZ8sEkK3r9SXP8f+TURZsaIn0M4KtpJrgn6nDJ8MZioNH6hNq
tRPEHMBuVOoZjAxJBJ6hY6GcYivzfg0BHvRI8SU/Yn3uDsNUy6eFEbAad/+A60mR
ONZTktsoAtXZQrS6u7+eR+Oe1FNfuBAz8wL/szs/T5U939yWhqMKo6t8uaNfq20o
kAPqKfI+PB+bUHoI8CK0NTYTyBTrVZ6RfIMOGGu1+aigJRIavKgeE/6wVNlkCrMc
QdfwyhYWyHJBJPMSoTsxnNNf3rHomEFvfqLJ6GGYCovJsimKa8y5qDsUA5L9UviD
kO8zSbwLVGxNgFf+HUkNemDUqJwlkJT3MNpz7inSAkokS08HhO30nv6bAmyyMivf
LnKvMtxQY+6yG+NKa1g04sPbDATioFDQ/Sb60jyTrnEuITNcF5I3KOpFR+azbQ6l
ETpn3nXX067iNYeX5ZHBdYAjCkZ1myOkVC4FFRuBQ04J+S5Ph9Ymv91+di2iveiZ
FO5iLIIeQegNOOD//deoWMo8kaQBpdHIWUb8MwUUc7ZbkbFT97jYvTpHe+1UuRIO
0lCGgIpYXN+yVspXo3lkpxqXIchsYqUds+gInXSKrqKGZ3NayZVU28AcBZapNCv4
JXNr/ka3XAHWoHxInVJSICdPBwINp4NAwpmgotAvPz/22ma4rx9rRH7XnD4TtLBs
It5U+OZ0cCZrLizFpvSbrBQ/wEACYr1q8uK+uPWbZs4HWFQJmhrlltRY/S97YII/
3Ra2mzy3gVaHpVZmBKOyA1KKAj9J0QXIQCGTTI/auNp9KsGPcKI7/jlqglrI+r9i
rzcLV2jbkGNg59y33zJmBfVs5oaGzy3WqrYgR0ZxzhPA/b60qLa1wWJPlDwaTZrx
nREPhE3+w8DJDl8G1whAS1Ih+6iAG7uJoremkM8lcFASsjTsGXW9lIbpybQNn6fh
DJ4IIVOLn6HgChevtDa5/BpUbUIDjvD3eitVjWUB0/kMEmiBsybr4SPy6asPAsFX
+mPQXQoCyQrzatZ8Ab3hayN8qBDUmne8GIpxdrIrTezaximFonuHPbYos1xgJ0V+
97qWCdJTDwy9piBKYr/N/mNKtK4MYQG6fUnHpH2m0z2jpAn8aQJZ7z1YNnq7Rs5S
HN+EDXF1mldPRXN5ClqrWFBdHxVAE+uWAJFlrkNfmbqFgRam6IxlBZInV1ZoIrVj
uy66OQJXbPJVG2LjRCx/FDzjDjT5EfGUIU91bLgI0mFhyKPBHovW5jrrEKlB5iH9
2eBzKSHijSWRJaPfWQlaaMfaCLvU8IvHkJPAUc6VSOGGBwdMJSIjmCpVKpJnqoPt
8WKk/g8toKuVYA3BIZUCe7Z4HhFv4ill1mrHOmF9lvPWXl0eFFnba7aaytm+QG9f
d0+Cx70mJcGkQ70FBy/ZtiEi5HuHtkJZinjqzwdIW/lvJ7updjHRL7kQKj1j1iNe
Ss+BwSO6WBQ/BJQmgMh4aRlz6DyhaWrvYyqNw/yMSLi3KnRkGMBw9bCndj5RznSM
aGJ2+aQeZ6K70K7yt240z5I3CqlS2Z0vRwZGxR1pA/TiQNU0fgxMuCnz1VZhR7F4
pO6tJKj7zyV/dcjpOVNuCULR0iwP76WT7MpT6+WGX3FEADNOSL6XYVsGxmC26fKQ
TVF1WEvocio9VugpAYAIkGGSZ511RNjibnXwmJj+cHzzdZNvFiWwx3hW9TBquok5
RqJPaW2paDcI9E39O2iYtWW1ms5yXf+lpiiKf84TnDEoYe0+jGk2HlPCv9thmVm0
XLljKjZ9BlfCxyHTA4pD58NAA5/YCe2RKjMUQhh0GGNr28XXjJkLrvTOiAUG07ga
u5O08Wwjh1lXh2ml/auN4PHovAhmLa//NK2yBXcEjlBslshVSQZ8OqxRsS8sgXnm
O7DMtwSUg5YUfYq6LogGdZl8A00n6drQCLFFNuAc0miCadDu7YvKNL1IbMulWGTr
3LVDWL00UVrHO0rdyUXOrDCUfZsN0Va9Ax+SBkNDnQpX9WdDIiqRro90ekAqM7F+
UJnoDqFAqRTAkOQBQ/h4TF2Z1fPNC9w4wr6pjUsqyLvwtSeoLgvzjnaTgc9xz8qW
PNEk6YkT/QZUiZjEN63B+G5rvYhvuc5KCs7Dbp0n9RjrGKd7nHAG2w5HCecMbXjV
OzZ1ZoaSkDkb1cADrlQhLRscyXW7uA2GymHIsRryVseVzy4VxbM+obAqdNpG83YX
14vi6bE0P7XFd/2G2LPR1ymInwKD4og6HEd+1iy+mmyec0Y/X5ED9yJV3yvfrNPr
J0Usr32A3151irQ7VBNwBhaKEomCpbDLNKF0nheThtDD/SC2rMcD6LVFPr2hWOFG
OQNfSRTX75RRpb9Lum6sx+AmsSPeUiVTZsryuA5DTj8m8dlkeXFKEwcvIOCYGXxV
HSEuJHnjles/GZgKB6ykgQaLfN7UyzyBLuOiUvw8luhGM+NzTpdTnY/VTEqrc9nk
rvrQ57eSYS4u4opaLZ5V1VDo/6bLPGj2RzvAXHZi9cN2Wr4IiZukOgLAKh5zwYp+
qFUIWuMq6YAa8iQKcJfxUFCvc6PrzT3KNTtm0g8+WIWik9JhyQf0jci96+Gz2sps
ZSrLSroQaXJX8C/EWybMGnqbq0UBeBY8xbJt4DCkoH6skzuXGDKLGUvO/CFk4I5P
8HIKOg1iIhVp+pbdythdSnK0eFLYrMKT2ao2Eut0xKGMWDGfqUkE2H8TBD8rCbTh
YxM+DCI7MSDXP5cgnniSilF5GXx2wVpq/yu5CTu0J9GbMfZosb3OgIHVvKI8Pze/
6utgcDapTg+u7IrFB1FTnUvD92haPHbPOBnaw7T3s7wtcHH6u9qYkkVeFT6OovM4
42XP+d9DJGiT/JUnBUQmQ4vD94Iruw18DLxngJutpjL2XZ45yW1waxnr+/agB99r
OV73I0ypeWG5sL9W6JGFyhBrhf1luUteCNyBNhWt0zawpNUkQDXfGLaAMQihFFC2
XxRLDOaIJu5E/IzxSEOGOGlijs1zdiRSBMzRMcA6vsUw/fnx0W5ipafZdlAIcYkt
06lS/S6gxHS2LcHG6dI+wzPbVk9pIcuG1Wu10xhsKe7zk0axZS+zJVe65AAMN31k
B7BcyiMCiY1vD6wom3mqinChGLr6sUKEydweb81v3w5jFaXPHoB6+cCrdtaUulVR
NY7hbxZHtkxN+yes3NgTNOVJr+4UoLpN5WQI2eI0OelEA0wZ02OG5NAGcx8gFhuO
gmwod42DNHdX9+79w+ZzHaABg9P2hNIOYkrlGQwL04t464TnTOj+j8pzsrPSrBs4
7jUad2bWPsu3xE+zjmh2v6KarNIj9xp6we8qTTYM5Y0nj/4ZqIlb0Go6OwvyFj/9
pht/fatgiWrkJfBVhNG1hpLGoJ5p5PHlVe8KIOCMP344xTl20XlEQYaJF6E4wUPY
LFaFvfgk9LmhlXqIC8S0S7nmejT4sg6h0TQPRBejG0gaUlwCEGg7r2AG4bU0G2O1
B69Id9288IrVsGCukIReFOb/L5epv9nJvUg8ZkINfmUGmSD4ir9kz9NcakewrCtS
lnbTQnYbKdafLW8BMBTXpONbtA3ZuQ5vk017xzKCJhQQioMTfHahgAuoPi7Pq2rs
BVJj9dcKFCbOkVG24EhT6hhWBpOt8q2Bs+UdY31/M0Qb/4kGHGzhYd0hF49Ccxyp
ESCS78kH7BJXrBoBEFm74Z2IIDwgzo7fjdAXVYXxoQTA5SnVZ9bwLmYz6//YZQBX
05wbRx0gbgFs2zC7jZydkOhX2jJ8lmP/XDeIJqjh5hfeC7z2rUuzk6v0WePBTnOn
kyEKkiLEkqFkJjAqhSzA5VFbyflbIxIvE22LMUDJfAYteGExvz844cTUXvCe212V
yI5eZNHHVnSLQkKohlk+0Bc0NvR+Z1v6gaMKMfuyQyP7rHr9E9N5pgu8uqHykQfK
CMh0T6x9XbdVxvUMATID4S55Mkvvjh+W2e7y1+tx6+KhX5ixexdRAD0jFEYqFfhV
FHI7VuVkR7mGNIL+DAtInqyoZO+14oZLKIMw8VskaTnxdlOE36yMpjjQ8JesHkdj
jQ2lcfOL3L+19V3yfqXOJsrYyTxrLASVJF8NZEIkBZ6Ha+9u7ZZbP78befPSlskg
2JJq3jCd09uiKd0kjoS9aZXqIFeNKpO0T7E0gFlHl0SHrEShjY9SSGKEpTq9q40P
ZuZhh9KM0fSlJzzZFNjBr9FaTFiXMMhd86ti9cYH40lNbM0Kvhk1TRKAdAHZnJll
fOb3AxCaXe4o8Gi+6vQbmtmHYsgTNtT+y/t5M6bcSppsHi6YcbLf5wlWa3TLHwFj
pMJINhs/BqRVaAZow433n23NMTC2LZUaWqfcim4bncHyaSDg8kdwos/lxcX4HaKv
P/kTEBkhXauHvHfp6bdxh+7eycighdapNWrIxVzy4eugyt2cNohia1T8h/yQYaiT
AqVMY0Dt720v6rEe1ylsQoq1RwaOQn1utEiuCdy/mYapoq6AJ7yCRm4y0/I/a8FC
k2/Rr4shwTe22fXiAEqlufOWP+ZXZ4w76BRr8ePD9/pjEVtwsydwKVWvv9tCU1wc
SiolDZP/oVvGrYBWVpyCcpsq+q4q+ZH318ZHR2nukb3Z+wnXVmWgOU2HxJiWjBhu
ycBbxhbE0/7mEc2o7gy25fm51cQ0WWmUIF/UhZqt34jyyLZeNNPWMiSiB2QKZvfO
lsTTFnv4KxP1aQBPOI7yYWk0jFjjUFtM6XBTSuTDZY4ZNG/aDLfK4nw8fhu4cyAx
cygoL0jceE4579c6F2I4rM1+bytWUd1XSHZ62thEOAD/ajHU0C6VquboEH+rU3PE
ymzO2xnefVcZU9UKRvN2x32vK2usFajWyaZa0hPC8T8E2qsD2nWh3kW5SRyMyQ1B
TLoF2AN+NQO/9dqHnkeY0ASFnpgQwtJdcoweBVxk3ZGRV+qycyPLUTVfzhaiIZKo
izyHyKoWC2IaH9H9lF13ltFM5FKWVYDHduyyDqonF4IQ1jw9x/1hbDi3FYfsfsGa
Xu/QvjZm32uSie6R6jbJ1qTydsWHKK2xx/YSMeROLxJOX5hFmnk0qaT3Fv9UbswB
wP8xU1h6aJkHegOx9IC5YWNG2uf712e7vKRgY10WCOZE7W6SyKWICpjsCPH7asht
v+yq82AAizrtDeOALSp032BYPSc79HOPwAi2VhgFBUVBuMXx6+2Lncr4w2mtE1MQ
6dMF/zs4L3HWg2GwmySerkWAzglD6YMzREfSF+bem3A6aKJk6epmNDClNAp48dJN
ONmt9SmptYJgdFNPFNIScuDqhFRKHhrMiTYsPpJmz5Uel34pGtD9mZiKdO6vB5S6
Bgk04PFWCTkO6t9zEgnxFFwAO1q6zgA681vTCHth/+a6JJlxkIialn4kaU7ozNSu
RhmDzNPcih20yAkz9tuPmO+XATas3f92TFItNjo09eA6GUAswYdJeJpPTUo2ihmV
lksX9XjAhNSDdA+DRVyvSqMlUnyNPCUtR6fVF1sMk9Wh6CbwNV2H5uMwSvmVNlcS
u0kqU3ZDnAj3BMNgRXH47wIhuBG64q/1MCM38VWIaWaPKkrWjDgAwc19LR2bYryW
7pBDaxv7VW1puA0s/eY8jxGmKLFYZX2cL23anG2N9Vpgu7zFoFcYZqhiqfvUSyox
rs0VKRnfWcogg/cAbP2TXnnNNOpEejSRykhCCqZ56OH+H40Fm0iyRODh4G3IkoIi
mOJrWfx4a99tKLf7lXLMm/GAxa7/bqvS08omBiZFmJmXY3Mdpgpt+vDTnWANtb91
OJwuAQ4IAHNJ+V95a6IVv9I42ISatztPFrNMNIZJXEQCQ4BYmjZUJ6Ra2JZ03CLy
irOd4Z1Fbwy2n8WGqNNvl0rFszc01lJrEHoSBzN8+GstPohI4uypkixfZRDmW4LG
ZYWgO6BgvRp8C54V1MgFM4eiN8Fklq/wguMbKcOtIQIGp66+Zl7MW1bGQkXK2DP/
cRKugFPRQiq8IiJpNQ/5XhuX++R7i0NSUrnK+z78hEKfKqZ/oi/ahYphUcJ4Mqvs
7So3aKSQkPBrTuGgq4WLgPi6QggfrIY7jqTh38q9Bi8z2t5oI0VC7EszfVHRDYkU
MuBrlbF3dmoTeuGQurO0MOuGNuIioP2ZhWIMsRz+nkas/6HvBFaqd/SPFPh73zGd
liObwuE6uxy/mHMgjb897zP8chXhFoe4vTwk2HkYTasHX7QpP9CVV+mOgmFVXNnj
GI0jnG8uC1oAHxdUmKd7qRTiNu42iLk67WMO0XPaXUudz7YpTNvbeawNY/fzl2vo
Yxd12JlUC9VMMd6vjjJ63aAr7wQXFy0IbttDIRa/dDjRtWrcWa4PsP10gBcT+42J
uwlRs/19XlCuuXfgmxe7NTp4TYv6MaKkLznILkQLL+sN53XV//kwck3yYSF+vpe8
M87dBjQ5asEsgVebtqifFqN2nYHVU0yDSroKizaOHrHHV35uvJx6zumOYT7mGSKL
fPHfjj9yj9SlqUNUb58OYvBFWSzDKZ0JruPljzJGZYtsxrGaS1roScFdx3s9lgsF
cG7G2/hwi5GNnkm9nUacfJkkU1zH1SSCLIDv0emjhdKE4TNpZR+O/DNhfZ1hGb5c
ebqJVft3IPk+nVLOEDXgrdzgBHHwDUX9biem0bYA04LImxtl+99Fxx1n5Tcwq52i
xhl4zYrx9bNYmBtUeV0TdJW8gfohI1l9piVsGpZTt5RpWYYpGR9LCeTEL1zhlY6N
xSToh1tgGjk6CX7ruNGF6G0OkzYH41tarZqMqN9d1DIEcB8vh3C8V5jvXlQX1Wgc
9XOtnaNI56rvMtpbz56N0hvZQ7yUXtmW5Z6pBdw7hYz/DbYfBVaJdBvnI9lQk7ry
n92LxJEtixZ6G8iD0iw7g8bVQwgAPGNHau1e/vxWOxicR9S27uigbzcJx1mcCxvN
/vWDGwT5C7Uom03p7uQGFNNpDQWC6Y6r3rSJB/oVEiNE+zU7TWQ4zullZ5akClgh
yxgeWQR8RK0uQ+nla9x/CyODFSlnFyhTQQ45HmjNWZ3MjwfGES+54P2WjTJfLRZo
fdXsCi4XYluw7mBI9S6PUVMt/KAdeomHI5jdqe2I/zqy2TP/S8XtTcoEfck8r/tl
3kXJ6jWkQ5TEIu1kN3WsiAoZIjJxSK004mUc32G7b4bEkQ5Uqk9DMlMZWkdtHUqa
d96FIhUL2TiZ3IS41ZH7eB3dHWtXRexQXAPXcb9AH4pR9MfQjK6hEyoJdAwDatiH
PZ/JgX/LWJHqRjWsTO6tNZsSOF4GHCMCHFJJIlopEg3uxx7oV5Gfs1RZU3g+PLVr
/oIzh38B//cdhyrcazhWxqZ4syX6uqHcGH65rbjjNP/Hb6xcLC+M69VoSpktdmit
vQCrf8fqJU+Mv/+1eVS+OAaIGaagQWxbY5VAOfqFLuKKFg3NakSdRsKxDY/jS1Ea
k0QB5gPdHMrY4JIolHC/k0J4hdyxCMhS8w7DiUF/QXy2ZYSLHhRK4YyeS400VENb
64Trnm8y9ugVwIRNiNb2ySlDjFISPV+5O0S6vOGe/Oor4GBv/w+NZhNF9WQGlRLc
iccTLVWm18ANYd0TnzxsJ0A0rAWw/4mPKUbePLaHyi2xJd4clL9l4JXf9R6koj+M
N7cADDxcp4+m1QKkUgWhlY/n1rsLeAMcc6ywMnXs3G7S8PcsGZ9L5efJ0Gj5dl01
jbBFJCgrrqJv9K3stvnES47U5FrqtbfTgJYuRZpS/x6bvzVKYEfIlfAAtdv/EdJy
GjNLdLK3pBvL6YG7MUEyTr1PAQcVLoycpMK58U0uPfewc/62Bxf1QD9BI+a+QzPS
L+wlArvvec/X2rZfT0IuhvZgXWOe/wrHcjZlHda88U3/NTMgRVGekBkajpSCwZ8y
pyCtO8Kb34nPsZePY29ptjKa5/23G6tSg8f0vPL84ycgqgVpIReckdz8CBww2LV+
l3qGr2SxvueDUMhcrkAoZ8sTF4ezrC2tQe6OGKqnkHDQV8HfkZqTLdzi7QsSfHae
ESX9+bkCF/oG/9TJxyd4Z2vCpeJsCFbxe/brvIrjB8cdLR4TPcZTrVVKDG7Yl7Tv
ZTno7MND1KdokL+fRKYeo+ze9K4eo9G4jhvUffRTYEIsJ1fOFC++3nU8mBhCpZRb
X9rAHVNFjzUDbw4eetQUsDwHfbLNvX6UKjaF6mcKeMtqu9D3qQAksN8q/lm/1+17
oMNf+tmA6Lo9g/bZ1+L9gAkI86Oswm+nYTu0OpJMv8VoHlpEcqD5LRpHxnoDYMpi
tSwdVTh0t0iau+BvMxzUvjgRrJgtOA5XgYCWjXQ4ROISVr/kDY9jADS2/sBDRtk3
aWB/IELilZsz4/g9clITfdKzxtFOdDj2xVemjX/xWguhxcPGHwLe3QqNqGMoG+rB
O/kC+JYhhVApt6uHYg6RcjREf9GZISNaaOgevFMxw3Dglfv6i7n8KSoSYWmsKP2k
kcbX160s4C7mJndHGqFZrw7BPCOwJPDNhRKzOGemHGAcZGNzSb3FBHQ1lBl+hxOY
2LowSZeoJHhpGLW36xodjdZm0cHTvxCC3dlV03OlxS47G3D1dxYW9ct/FI18oHqh
Mk+wYTFdUU5aTrWUn38dg9KZqY7HO5MqdVbVMoCVbadJ5TVssPXuxi8HsH5OKNB6
xQkj4T/xHY4AJRHAK+scw/QKAm+pdEX/ZcIG4d5p+6MbtOe/kf7vae21uZw7cU0t
qpjMc9lcYF2LpYLYnRT5V0f3AtI4HhvD4sDTRGcRnWhqLoW6MxuFRkocqp0p6D7u
lgV9L319EuagWQsumYwqdfjbtPMNIvktfre65oUtUgFYY/nvE5Z89/r4aDgU8Hn3
imjDPGhsHyamoBiqqSF/pCy69RPyBUqJNaUTc/7Xo06HxHHPJNUL/IB1ZsrENS5m
id3kxXjvLcJo+IVW47fxJTp7WaGGllnuvzcYABAxIYNQfjQSa4C/cyUKJ6mN1quQ
Dkf/wR6cRdGMjsBsPRd3bR4CKd14kjKl7bje2LHpUGJ2AHseBkjj2oUC14yBzFVv
JcV7nnRtqDxICn5YOytdZNbHuMXrz6DRXKl+V/Wlb/YXzNxJkRC6CVcGKG0aqo9K
bQ3ygzTyeUaJCksF15Io640728zyZpu+NSCEipUoXDaD2g/pcc7padLwNT1kv577
GbDIRa1On2dHlfouxbgLr18tP6q+7PQFdXZPSr7mIoWzaPfhsnb4Z5Pr/ZOGBE/9
ZAysX0GxOdT0WPIneOuCDTckF8HRh7D92qppwXwrZ3KC110KAJWSHRjRkTdC6D03
PtVm8wSJS8StzjDr+JG57jICGdQmq9c7coMuA6qmYTbUchNz/bM1x9jfwzeMm7s8
n0r468kaC7jXzXkKF0JuyrGso8NNaLsQzF9cRrn7oGwJ7CAVWNZ4GYOrOhJ/WGDi
/BEIYMX9MXGptlakfab5abpfZRmkZZNhcwG5Vn4YeJOjJVH4+ya73f0xeJ8uvyNV
3IlWSUVqcEwEEYLqaNSbEcd9svXTlD/X+b6EQNmGzZk6odPQZQq5l5XweLz1f8MC
xqVaRD3xUyFKiiItMLBbGxNNP9vyT+qNF1vb1ZOJbEVhGr75FSN0D7vUHn9Gg5h1
1A5pJZS/iwkuWP9kQ1bhjIUwA2hKKID4pS2KP7LtUIPtXd0JrT+qlszAkDtCgMoB
LnB0SBZqlFsqkgV0P1Bpl0aH29ywB0BthBbS+CxgUG61ax1vsqA/88DUJc95xab3
C/P7ybM/roPPTvOjXRRp3PukZHJI6m6pJMSx1OIa2UtwkVAfcFi987/7v9OsfkUi
N8yW9m2gqPUZNU3Rz9mXgNMFih5s69hGUrH9aslJAD9P9d8NalVKJsikyy4pn11l
wy9h0v1IIlv06mcwEy+TEsnRLS/FnM4YNR1xn0Q1vRoV/MdJXMSBEBE624F9jgvZ
ZytD1EmOoJchDsWGkmPQBGt85YEbIKgMKnqviioL830Wh55PWTDu6FWhsiqi9xfX
+mPOgbPMmsvDUTJRZVCCZ0W1oCDgcMeR7GpZ43RgvuxUCNG5mPkXTT31UappvmnA
a5DLytSf9PiMJvtt0ZsgPvlr3oXmXmIXVddQEPiindkVurAjVfCgmRckJHu9rZR+
EODT+K5dBFBwEoG9LStKY4dxFKcxpq55OKUReaLsDAP+4lwbJSpx7jGah5GOi7od
lhiRs7y92gp9x5gsOwSVQ4tMKNSLae0KlpnGsyLkgm6D2OaDCXiDtci7YcOdkppN
49r3rNFynaZkIRQuWNnT2+Ap1x2JudVr+oSHmIdFk5vytvR///7QAfkgjXvv93Jo
46smVKZAvJjLZS7o6NXw7VxVbTOhUZhpiwHIJsXPG2fLzBXtFujqmXnG9HouK6+x
WMQ3tfv4VR3LqBkycKOemzRzx9QGoroyMIUyG05Pw6nxi6PzXD36sdLn4AZVm9PN
fX6k1p4q510DQao364zr3CytlAAf5IXwQ2VHxHmSKH7/07ewOJuKdZUDPLCB8uAs
lLW8x+ggQSk2QdKep1NSWEq9SC+WyMqOuN7GsCHdp6uto3uUF7o0jb/pqLi7xDZd
Y57ieraEP8I1PQc85HtMpicJILkna9LWX1gBYXh60XG6o897/wUQvKwx7wkzocG4
1ejpF+mXVNZ9PCLwtNkVLl27AmQSHxEyc3E9nHcUJ1V/uKQhyUxQhi8a4qwBpbCD
go8tWNgSvbtmQJn9ftbxasnIwoLgIhmWEn4C2hUBelfdb6iP1uowMgHfP6cZG0IZ
zSVggmW2MegtprF9tE0xdX0Lxp0amDgmfZejDGg9L3fli/hXeQjEE7ulXP86Spdj
luZbt8E0sqMaoD4F4cF1L/etoXexn7KkELSy4DcrNIa6n8OuNm5AJ2fd/8zEsSza
R9K2kQ3uWJDTB0TY1NgitRsFZSbhEuZGvzZsLOtuSHnd06NPdM5aq2WkE4SB0bWj
7k5XkhWbBFEbKbrkHdf6QqUqP3hDDuqR+P1fhtmQZPlqktIkrlPQnBxoKJgR9RGJ
mMEevPFM+kw5wv0JhiQrDEALiWVYyuBvCYDNHg/MgIbtdF7PX7bs6WzfO6GkhKxZ
pvQ4LQk3c4Zr2AsCxPh3PJiLfqvTOnIgYxov8aI5/SkW6VSTXm/Dh2qwfZ81jeVn
CoYyABF0XttePV+JsLT8TLxOZ0awwPEMGwy3toJXNd6VIv9FJv1JUmXMna5mRj+S
z2HAgf261zKq3VBIJwBbV+iaxFtWxZvgRBM9QnV+1C0hScBDuJi2Y3Vh7iQkP5SC
lm2ysWWkGFpxADzSXSAB6h+5oSD95e6pOf3wyGgxNhqIRy4ZRf/kpaX/ZjBEd0gV
elFjWo/WTc+AF+MZqhUunFbBK6Crr20Cg7AcVCAomRnSNub2gNSkSEkiBv3nqBCa
LdBvmi2Kg6lOlglABqXw8bADflAzACQRraaOLGhQUz2DqxWl95PXWYyOH1e4lVEM
1xS22oU3KE/oh394ROu+itZPfRynELTE0D1LZy+NJT0ajdQhnbX6jU2PZhUREu63
yo6YXdyHQBlZrxWebZQZLgyq3x1v2DLxgNErebaxZF0p83FqzuLUVqKoXXe7Cv0K
A9ReTXGinwLwNnhItp/pnpBVs6LWoWZAVLSOwuNzoMpZ/kRgJpkEHbq8XtDgbh8h
8wOXiONdVfDfXDd1cxoE0eh5fTjk9K6duoMR6P5z/3zYU7x6kj9mmpBKbQOF2EdX
xsrzjFuHTfxtciKGWAU74LBSlI0Em037jiWroCaSnao0Vbg4YfWsiUvPeUYOt7Q+
PL6+nxTJjdIYR6XepqZ1NHbkDB2BwH8SLdj5XzT3VMjfTHSuE5hy1zCbRi3zqzTR
tlq0ZlZOtxGcqnQnxhC5E/6ev5fvw2WIwXF4G6or8MuZKAujeiMfJ7uuce91ry09
kXQwlnDQ/FCD1yKcEf3LeJGYkqREue7MxFWHA2KtrD8wrWylwKQatKbN4UpHLI16
Z+gs6Q/OZAQ/LiUibV1OXpYNs7uOfjJ5fRydwZRQDLTts+44d2uOTsHlTm095PUF
nHvqra4ACknVpkziFYGhkdueFTNYG4sS3V9tlkkuIqPvLAI7ssnXf331Xe4VMrEV
r3lXURQjAy5n0nM0Mzorv21qKvBWNweK/jDnQtnY4HDIhxqpjJcBB7NoQ5tp5BEn
UHKbrC2xqSgHY5lHEy+nKwXNJ8TGti6679bYKz8UCxXwjjX+zEad3sUeilYXxBjb
RHJZ7M1p7Bpjhm84OnZYHovpiAqInKA2h9lRePO070pnjs/GvewQE2/26BQIuFnl
4Dy8jcWMiX3i2TtN/WOvJ43PFzd9KuOnzk6kfHtQLSr2dwUTJWKDZ2SXl+cgXd8H
MNSxiSW9M/mPprt1zZW8V3p2yNxHce4EbkPPnkjr3b2XdStB7zua0MPXj9ucP/ES
rQkobwV3UVG3usMcC0LvCVQhnZiX06Wj8Q0BQ/+ztXmILerJDJMe7ycHtaM/l02F
T0ubOez9KN2AKKj28p4xLzvuOH1HjpO7qDoMZtDg7hRk0713c7PS8ezN4TX0c5g2
F5pwolfxM9AAu8cwYUI1Tu+eQ9F4eg5y4VgmvKCbnpxJa0zSqRUO/Xq9A9ivCrhu
BzJyydXdK69ZND1bLVmLQv4UWwnYeZnKWGavmr9Nipj1tCU7XFZON5D17rDwy123
kH4RVKwSJGidFqrs7vaEcXRVXulcpxRJjMxY02kDLB7NB08wdsvhGy1TyT9uEq5/
4HO3kiTLAPq2cbcth3AArTF3NFN2QoMbFdBgV+k+Y4ZlPviXgsokA4yCc8Hvcf/k
Qp0HvRl1vlXDnEe2FZcpRZBAZFs/Hthl7UIxQLE5Nwht2YwoVAVlxJQPevszL8uj
HY8IrEVBixB+2a6DvKngaKZIDJFvUIbzkb/1VyoxR6icd6XOyxrRuK/SUtCriXe7
vVfhueZOW3aw7OcoFI9FXcexxRPw7iSRWu/wv3QBZiu94uzqDDHWmIKhqP+inm9K
CP/mrIsErE5lo6EL6PIpCGgoUaYbKVpok/vY9Q/0YjJt+ZkqaS3RoRmUbSOt0Mln
mqhBmGRRU8k8nTkYXymplX4zXThZXUFv0KkxR7PTuZ0z3nBX8gsYHxZrM1ZcZQf/
8F4M19QJa3NPgdwSBrWt5ap/aN2sJqmCX2aUB3BiJP0JNEecPDYEq6zrCUheyMrz
8W6wRMGQPRJFUp0iRLysg2PA7w0K2D10O9sHglLnCM8D86XApwHINDowHFMw6aBa
f1m1N9qYGECwShf2bB3ZTT0xiCdiZoNBzVrbmGLrTRyV5rHB64cyrFrVSdSOtsh4
skhwzju2kT+wF1RdGgy5FsmyNfT/NB2XQkTbqkjvdsU97TaXZwnnCB3Ejt4mruq7
xN8rBPJe4XVwCs4dNAvmMuc5iEKCO1j0LiwReulCLsf3UX8miowiqbcNR/N95N5/
hSz6CpQCLt8Vlt/p7RRJryTerWyGnioJ1R2swZr5T+EgSCD959GI6nRP2gM0yT2A
epMgCq8oR3JsD7Fax11moNESGEEpNL6wgZQIAjOHrW2r7XC4RAdMttMmHPACKNq8
M337aVJpXSk127gIK/s7/4+ln/8ltChBOBhV1TBi7z1SCk6XDtIlu6Fnzwu9670y
lhlrOIjd3FUx91QWaEAF9RJ/3jUkSFOtCZGM/CBaJUpMeD+D0OyY9GJT05EWN+zs
gWxLPE5AsMc15Asfjq5RjD6wCdHeVkwzq5pK7H1hDcgUGNsVXN+thl5L08xDqQlW
/T710Knioe8jJed8B4SL2nI0yDU/XoRDJP6UYaAesY2VIlYwFi4o/d0e5wyBWwg0
qXcg4yQbtdk52T2sIDXpcXPMCF23ik1MTFm+n1fv/avkuI81rQ5dEv+V41OpIMMn
I/IOykzP2EY0TlJZTDS164S9EcmOoDRBsmul2bHLqMHZpashekDMathe/EMVqNBX
iLuy/xifJVzsCkSJAXAN39SYZXDR11GcZe/EbS0qNDX0TQiYHHfTgF6PMH4uoCGa
143ZEKTup2zbexQ8Z5P7IcM39sSOWBYk1GZuIDTTleGX1DPxMZbL6SGew2SUzPZK
U9nRRkK42LaG/wsbc6jKr3RnoC+CXaiuBCAPnBsnL0yqpLLRaVSvu6mq23ASpAd/
CROViSgF2VN4g3F1BdM/0FaR7GvZ+JUxq5eTBcWcHCkPlsAqMHWj6Y/1Q/HFggrS
PXEumji0FA5lUXTftYNzoE2v4bYOOecPM69ri+bT5huq+xQlUsB3EQAvIT9ZmBR5
GbgxBTA2/h9heaq2RsM1xdAB605kym50Q6reyyk1tr8ZmDiY5HPh7hP78ErxyoLo
GH7Fv10fQn27399IS2p7uuuAQcPYasPKd7lv0XEBs5QdPHr1KbQkxUrkxFWVxyci
qXYfjI1nbNmdjcmXlVAYgusas/8llIKTrECIVEMnYdu/T3GGmJYYJJm7yUdmarQT
zOKp8fyv1ZfsJ/zQxStD7iGEran1akEaEW5azeXuAezTxvJZHSBvZhnHQEwjTjMR
aVhdFp1Ykr7Mi1Ukpj0w5yPkxxDcvYaIVabnMarRVpMTRvsbOvrln0+PwM0OIGTI
5gLZ/2gQGAs5F6LZFaCYnWo3OeRDmSYxioMAQZqP2Sc1YKlzieG9RoqkQ7UHMqPE
xt2xPt0UKzHo531OXKwNfIwjWFFS3fymKc96WoK634pnsBxtPdS3qr3pwI1X8Q5O
WFUGByOXU66ocPbxhOSYAfqUesfYf1O/lg8lzS5br15Y+HFA8CVCUGBi9iLc0Zif
Rri9w9WMEfJsE+XIhxnj10w67zEhd2keHp+tE6ROi1WdB80l0eniWbeCcNCFi9y7
W/lzyjGj9l9rxA27MqPltG9Rxxo5Z/BWBojbH5h2Zt5g6Xyn6T8G03tntfoIi+lY
dRlyvfq4oH2u5+C+gdQxWZskkabfPhKAaOhiwKG8WWVZD75/7beXGGQOtmf1TB+L
/r/wwaZysnUJNiLpt+NaRvDo/8rldUMaPV6dMAT8K1hELuNb88ZE9ENGvhOEQsnn
uYLG7cFAqsLC5EibiU2aGL0Fp5fXjwIrN2NpyIXgJ8RIwsZHoT+GHPBrvCU/BEoJ
WRCRPEqTwcHb0SZnqEMZO+wvyNcYt8S0NlCDapbHKFppFyX1BDylCkpr0/BvKExs
CYyEU5KPLXuoF0393pYS+MvjP/XfMPLpDe2YMDCIHPnb1BihBl0MqFYUrOzoaIeh
kQxniiSiopGVIy5HBiduEGdm4boXtnWh52+4w/EELAoXwRaKQpPK1Ock0C9xf2Qr
yYbpScuLwTVlprJW1Icn2plQDx9THpCkIlYGhcXLZ+rI1+HOjzq8jPxGEa8IYK8T
NOxKClUKy4EhPS1eWO30iZndqGX5ZapzL8GnRKH/9x+LHp3K3TEBUSauJMy6rmBd
6vWDCbi2C+2bUDM8YUqEb8iR72AE04Gxg1+meRP7gyBG91usG2oIaVbJ/3TWuQBf
vHT3IBzV5m0uGBIh6YAzpyG2HYV++vSJj7RhfULs7NI23mFkiZNvR0SHgTj1gVMT
fnqhbP+DVr+4S7Pj/xPl5lJYv8TnJXydJqVu6MlBBDWB18lbZqbJKNS4bYNzD8zy
BkqDF++pQKDpA6Qxurl3ZDL3O7ysIkR4OmdOkcBO+kP6z0cf4kDQo80Svr/ScTvk
AIjmMpWR9ZfokTNUqNoOy29VnPhs2CCmbZkG7FlDJnrLjyBSJMpfgfnRTLmMNZG1
7Z+5+qxvQrdbq6CsgmQ7YYd2IqY9jbWh8tkNqHPt6gx0eVymvtgylHJNwea4az4K
6KnJWWIUVZA+WPZaRxharAKzgpXAVRDqJ0oD2f38spWOWja23yNg4j/4ZCng/QyK
rogloXXt3+1MZ0A1kALh0nYu6AFVc2YeFtk71xflGV9TK8gbdzQroeTIKbGLpcT8
xeE9HU5lU2s0fSUNTRL5XqeaCvgvdwifr42FSSxn5cM0aauBnCrvChOsP2ofyxwX
oUKqMhb7CIim+iuna362F82lLhbKOiXBYDn1DxGYy7csZoUR8B5NmXO7hCC99DI5
j5upV4Giydgm819ElIeja+PeJoEOd7dj/10xEi7s5LIlRu8dxhKKt2kwEqAnxYak
Qa90xy2UzJuqF9wcgjHYeuR25NAxAlhdMsI/6d0N7x2vruiXsEg8PEGGPTeQP8nK
ui4eybC8JWbPs7iYet3V8SC/hYccCayQ9XAh1tnmJQ7ckVvCXjuifups0gEGo4Ec
nem0xpjv2XXq05uqBpHNz6vFRuDbinvbHvDFzpNWeBd0XJJSAG0vjndRCodNCG0k
n0x5uVIZbf2JdXxGz95vt0MRZAph2jOUeEpLpWtNB3a0pf43suXZzrwPT5WevEeT
A7/Xrbvoq3di6Sz3tPaXFBzbEjFblETpCur6ev/kfoidoW6hEmQ4tnSnBAC/bSdJ
u8wGEXS4YFTgR743CGFKZkNv6RzM6LMsJI48Pu/nKrUNV+dHOgw7slWt++4AY81i
NefQjsn/RWR0V6lsPFt4ICPsyaZfCCWHRiJbiVeYugIqepY8cU/nPd0VeAuQAfBa
yMOXr5NlO8C/QjEN/OxIU3P8cBy1TnFR2a9m9gMMrkuza1XFn/frLPalzJvY71Wr
SJYG3H08cqep3aD4W0Nv4LhVRsG0vQSuB5Ws4+AvwC4MRo+qVt+EMHtfynuHxDT3
B2N706sVCyJJJ0cqh5vGNPNnkD74prceLYlKAUCE7x1s2+OQhJeVfG0jU0V4A/KQ
diC0nliRpB5Ad971ggOkI/2nt3Q7CbtvPfc7pZTkdijJCQ6cANqwXBIPjoOM76Ta
jed+q91qLV0hwqpQaG12z8jjJs5+hN1lBHJ/x7H54CHVcsfHVLjut42PXKsfWbZj
HcsB7RCMdNHEOG3wG8Za0mXP0Z/ZBbJiCNQZmREShdlo1WCQ2jEyCOQJ5ybFhm5F
c+MR2PA0Al+O7NTPhPRZ5AhoJhaS6cnJeCDeloVhhTXxXhz8F/GKG2GGNReSchVx
gakgW43plOz0+W+hXk2m/FB/BquZayP5WrtHjIbovi1etc6tIgm9+LVGjiHCv/YR
Uyy5werjY6eNW7XMx1xBwFC7icLNdXItuQmEYLR6IPX6frO160wea1Gx+MwcQBBi
eV0bQa9/p1OCfw+zhXQ62Ji6hoEpvO8hhDAALdw8L6Kg7CUfccEj/kUKP/KDb/cL
E+1hPsbRUhbFdovzVatdYr3bAL1znWRWJ59OmWFy5Iq9sYo23858jpdYu3tlKpe+
c3gMN1duep0Tq7pH3BlY5Rsh4qg3ALOJ0o+LlD8hQDvljTav/tarZY59/PcPwuCr
2BuMEf3mEhNfAg5MZRxsD+NgIaLeKpAykeMKFwS8woa9dw7KQMmNhKMvcDz9cDq0
tzVjVnfF4n9ttUv0BVw9N/XfLSN3q3pxqg2KEp7RYvtGAo3EVOU52Ivgc4CPKpJw
GNejtGjUtb//QcbzupQucuJp3/gsyMzdEsHEJmQTj1/X1UxMRgX4gBUME2d/mpuF
pNjXFzXXeegn900uJM11VYXA6oM3MGLQwLU5R5/0X6kwwRoLNcg5ZM54VEaJTb98
yqCwv03R8HLd0aD04dF2pFa0lLsvuvk60cimfBJUIXM9pfw2nr2Mr5i3kHscDigx
tEmNxHEwux6ThLH4XyUJ/cH4cqHS3cedIlhhj8RtCqTYwAQwTDQtiOvD0x8oru1B
o52VjjNrvrWlRk2ZN3+0jN1HnTBk+N6FWNkFpgPDhRohg8XrSlz/Fm9BvScFA06O
IttFsa/vY0Kx6mWxO5G+FyalJeynAewQEihBTdLZnlKfLDu63zRYA4d2qkAapZMW
TwtUfpLJ6MARZQeaTlErU66DzB8dMalVzovRsAFYuK3DRXC3N4ob/fo5ybU21ATE
S6pbzSFSyXAITnBdzRPsSJ8yDETcBvptGrgy9tLa54oys1/lKCbX7kXtMhNtRjUi
5FyFx8KkFfYkIglXLXngma1pPhXc/KIUybqXOPpV+iKyec8LRetXLX2l+h8YFxpb
gWci+LbcnPDGphwpOnODJnSKu69kszgPbsk0r/Rc6PamGSvf93zoUBDgPFTF5efs
KLsjaGavKeVhcy1482dAh4KtyXIs3upG0fJ7JfyArnTMPwBpTu1Lkvi7WqgY3vGD
dofad4SLJOsroQuLqr1wNbEYXjYzFY3VgrUCHXtXEGXEGzur2IfHLO68zh6m7KJJ
WUIG+fmJ2nGD4rebLCHjxcwxFfgbaTqcjrAofPQz4Gr1LjRneAWYWCJQVXQjxloP
zYAwP3CtATN5oLlL+kBIymX8UTzuRS6UIWO51RRJDy2pXCnYo3iU6USHaeuCcPJ4
rxmq8MN3wyEw/A6wzQB6LGkY1gEFIMoLW5oQNpT79og2xVoFPhfjpCLgRy7lb2nB
MoMTOZuENIoKwKo9opLDl1EzgiML1n4PEiMIvh8YyX7wpeJbuwavWREoksfDqrBZ
4U/wD4XhkOTc92Ovn3JK8FAdVEPV+kLdngPmkEJIElPzeWbbnTFSttUKCcRripIm
9UEJ5fWx4Vs/kK3pznNzDxb7ydkdKpidcMebd+2+Ak8qqoyb4RnDOBCGxYN+mlZl
9LnOAJk4FHKHx4vXNQfGgzZ63ND+mRmgBlwF/Md2LaA0UwbNOHbpY91AuVaOx/Ci
axj2eAc0gjnw3zlq7/RKrZ3iNt9nxKQY2k0ie4/gymE2uFZS/F6bX58Gajka9gGO
GVYK+uXchUZTXeIpKDR99+MzyHlzYDvyEEU1Uw0qW2+FQgnEr1Rr4fjuHtrOzlC/
dFAJY2EK0yM1O13ATOeZbnTGaucbkKEoq5PeRntbTJ4XRJizbgAru1Ss+a/6y9Z5
dHjLIVfD/BSjBrq4QvLDQ/IsHVoNhr+Jt65ddg3To80REjnfxxz5RoeL1PJ8xQnw
Gd27eeKRwVFh18q9WEFwPOImBZPZ0AKa/STVT9DamVlPem/Yb6Hw/HTtlwEMKawa
LGTNMPhp1M4HM1ouXFATlcveEbOuskA2XKaCQsOvwdOCDgooVjlpqP2P2z4nyaoj
dBu73/etlMbncG6zJPR0V8K1dGPoKoFHBJzMa64nB8HHOcngQtTVqOeieQ5YhkCY
SEqCWGtMnJJWLKgP9o+rA8Ng08peQxPWpNMW03QKVVNgwfHP6fkg7aOrPlU/VHkx
kMPSIIMDaADFVmT6NPTPlxAJG9AIIRyw9JTr5a/8j7W1loXyvC2w7ERRnfsAqoIS
/5UY7mrtjZP3efpCMf6BrR1hksOWOEkrgJfDrS1gS79OsH8vohtJlQO6xHE+8JoZ
PD+xm2C8ZJP1CbDcSA0rkYxHPDaUP8YTbPY0OqByv5Dd5ikUhAxBceONfC/2Q2M+
Yg+6TuejYXZ4WtZWFKeg/KvvyPviA7Zj4u7kwMVgmQGjiMMKfEC0SY6xaYINkKz8
o1SS8m2lGXmnG6Bsn2x8KuszubWzIe53Qj+f46blUi42BWpyRsVtcsmUPZKLmT3E
sJ1FJbQdbB59m93Pjhj/nWk0R4CJpWzHg1XGNvzVjEagmydsS+P9679pkHMys606
sFWVABZpXHs4rUamnjPSobFkzZ+llDBiWabztY54Ydtxs+TGQSjJepPcWCTpYIhv
h4t6zIYsmsvY5Xnx4md34zHK34EOGNozb1cQg+ZGhsj0fUWK8xmuS5UvXILORewM
5aJf6ckVRAihUlzpRbzygPya8uX3dXES1Nc1/YYDNk/xf5nMQ0Y8/WYL2q1v6EVF
pwx78cZKIXiiXy1UUTXBd8FcbjmJWyFiyDmYyyaDr6bsd/OwVRdG99W/X54ivasG
gCiMUqwK6q4YgxIz+huFZP/uuFKj3NYeaPMYbmeka/VCiuobMk1EVLQvT+MHmTqa
I4R4QPBS7LRSzrM1BBpA07SXiTGXgugc7x/5uUkSb4ObR7qiDNL1fKfewmJK1EqW
m7y5COi7MqDPzZoH1eMW7DsZhQ+NfHc9FDQEL/t0WcMWMMIYD5/Ti1rtFqdsh2sx
qIt+Bk8ALMghdXJeMWA8+A6Ighau11wD77tLwtU3eD4lOcpW5fmq7++uqnihcp0L
0lkAMOcfe2FwY7L1dhdCeoz5SpjDzsujqDZocBXbonbkCzbb6JoK78p/2hVLiknZ
jRch4xn8H2eJJnA0FGOjZznTQv+FyN/DXT7tAtZuhy6LSl+LZBCHqN3Vw4KRiSbt
eYDXvv1yY+4L8+2k+TExKfPE9LW9+uv1DEbmRFMVmFAOq9/SgGku3gkbcQHlpZ1n
F6EkVJ1JAvifBY+18ZUBr/Dk/Fvh8olnQzOS++o6W8eajv1hi3t65eRsEs6O0W2+
OSBD034eBCQ+OMHWCuNUmzsHWwvE4wgON3opMzA1IQn0x5vBU/sU2pQZ+DCs74yf
JuNF+bAsWwmBDeT+Cb2/auCcmqNhe+xtA7/ZngN6zLS/YzMWFhxkh4MNOB5xR9ba
Y1ETmURH06xKCp+rOvbnq28c/7vwKWGJKl4B8jT/XDrOVazDSJI6ALCTtNAgs8HQ
Fs+hcv7R/uzG2ltQg9yfu18rl7H5E9VpiUB5LaMoJtiZo3sm12L6b2pDaQed0SeB
V8CqjAhbY+gcdT9WoHPHVfMEK+4iP9qk/IbIdWR+iylo0eLVLxFBCaK5wOOfdbZk
4NpNnSUqud6lLoNawM0MOJT2TgYa8IAJq4RviQwIhDb7yknv7XPxIr+nmuhd0PMB
Pbrc0jtTqkM3BRcqakiuAjrkMEtGeiA79EcTUxmhkmA1hR2SJ5/8RCPbh+FzHK8u
YHBrtYRUIMDtM3SpqomzPh2TD1OVOVZ4Lnp8JRBNCG84+yvtfocRDajEJ3jtrR9P
jWFqSbl2Vo0jnkmHYk3+nwVSfUbJ2n1wlxZaaIL4IOAzmASegdKU7gEjnowQWvrn
9jYjSPhVeMpfKwM/tiwbqXFCPWqdjDtnSF4xYmqD7K2rdRpV7ueGTTh7Yq+808PN
r8vc3oWfh/5j17ArZYQ4O5qhJBA4Rf0KVDRZL5juZSIBroS8xbkxg9rdr1Ke0wo/
2Y3XjU2ePUBN/Vyf/8nvw4+sHcuv50EWSCMXREk6b5cH0QrIZVTHaLyfRP5boakN
huyJLLaDLmkGSR0y1zlcEufugmv6ZNctFdtKllY3eqMID0lOdzh0e5xeCWRL6zIL
kETaf2rYIsnoEcadJXoCpWFwFu0Ogl1NVKPdGekd5xo+IQTxWUKtfWZpoqxEAo/E
v1IAzqgPdg+b92wz23xrshzmMd8Gxd7nI1crotc5y5V8VDxhW4XL4ruLSlqZTMVm
QBthcDrSyV7aQyqk9Lt6uo6W5QqEXUSKtCPArRQV1b3j2t5oZi4Qg96/cdLn6TF2
oyGl0+EgbZkqIo9YVI4DpYd6c5ABbF5hwaNlHHEbNh/py7GX1xybbMWS/eBTjjVq
DLwDRec+i6RYUX0Zj0pHqH0Qu30Kq+B37xdu/8zXL6DSa904XOSQPTS9eGtpvmue
KSBwGteN6yQQgaktQ9o9c+3QLAv6ECPYPI2ZahSvjFL+mcaRL6bI2gEuDWmpeTby
nMWVsWZpZ1PQabPFqmf9Mrrfe4FSN5G3qzcnaPcsuVq3YuA/xNmbrP3mEtchN0Nq
Lce7lhiuVgas7QkCChukuyO0wcQkXZuXpWWNQRgGFTjyfsbEw2dPTv78PPvz2Gac
GFlajDuYmf8cf/HBuRIfsxzXs4UNqi6yZdZksUWiWHa4fWffEu0JyZvKxovaT1Ce
3VpuMsax6Cj2gLtiaz7ulKOmu7ugRlmLu/3kXKWE6xdVzKygWvnlopEaYfLU6YeF
qOS1LPYuM+MZtvEkwxriqX4/YMEFJ2KRA5Hedc3WG15Q+u6Uyfl6q6/vNA8NFyed
cK9Eu9WCHIf3Y0u3r6GqLFBSIdFoJbTDD84gaI3onKwY8LJ0Jw7lGkeytS6r6lZP
N0X2zo35AEmN5wm8GnD9miluz5aiOWITLzLiVb5SQ7Pn57aXm3qqqcYK6BRFu4pP
9WIuiW8+APeuyghkiRborNu6+rD6Qbj5xTRQn35gt2U4EkVNiDWYcE9W4sX48VOM
3Fmrag5vWV02gBP4vE7hWn5QVw2fRq8NmhElMZjPqpjCh3ZOtAWOApPFAYWyw7+P
N2iO+Y3FdKHcgRmuOtvwx+vX/Mja6qipvt7EyhpFow8UjyAOeO/AOYORg6lr+Fvx
lQMrgnnVopAfzgqfijsVFRMbpi5TuzpqHUgEunLVbrQqwc/C96K/lTmIMHayxo69
qCATnP4TVm+aR02RtDD4VyNCtprWTgXWGlcMm5FLc4RDW+72BmgTMXG2G+EDmZiD
qHHU2+9pz5ST6f5mOwb4+igIoUwBBYd3+LXj+8Sz/mR40LU73v4qwvBUKnGAbfs1
8J1ABbU7dCWgNpcE373mUoIiRJVnIn+TnNbid9eI+76cOnWCQiL7sFK/DFd+MoEt
OVHfh9A4TcGk1OytrwYiB+AqTDxX+unKSz6F+Jc1bTcBMr8yThtK/aju4mp30BHM
56dM/0hEieur7PXYMEnd41PNAwcUpXgIovtquLkvsBHFy3GH6tkei/lO1Q9X/7vD
CVroqgl+2uuclELUNL+TOPK5lvl+j/9yLznZIzoolMSjBrUe067UhP4tIXRTy1p6
OnV2+ZHRJ0o4NC2Vh2Dz9VKoQWCoSfX2Ab4OlbwOHkDG89TI6CsT7vI6MSqgKH39
u0nOR1u8ca+/Q9Mi+4hw+TX3PjN0anp+eeyzeaUk8IT3f5hdzrmBvNIBLLqaSHPZ
rsJHpliCTNdfmAlq1kDntli9d0ZP+xVLgBlPiciFePOid7Ge6G/v+c0akJmxXIIq
u5i7o6ksxsxGf8B5fq8OrHVMVNOXdnWr2iOQrXzs+xv24FmgwOqqJsEKL7phygdp
NsESjcjXW5PtAlb/vY4lC8/q02ZuoD+H21EWwhBfdIcGiFBYJideFp7l0MDT+1kM
LWWEbTBLmkblMcDu5c5il2r4aXs4uIYMppfWXverGCr8MHsLZgJva3CY3seVd8oG
Sk/qb8yUveow5vGEFLRRevG5wk6ETiC3eYT3ygm5Bqa3NEqAL5/d2kpZpP+/F6ow
dprE/S7V9Fw2IjXfDVm4yR3OLdvngcyt4MTSy/5IFH6JlRCZHoWrU7H5Ti1cLwvf
BieuglO11WD25VMRPmcE7KB9i6Shnq47Bt+sQ4mYEyp32TqOVpKBiCZIFo9fte5A
xtwkHm50OCH/Q1Lec/BqYDIjKgLVJUB2tCtN6tSLOiU0EZGUimxcy1zeaA48d7hH
doKFfA2Ji9QapMA3OiV+KACa1b7WqwsLianCRsQ1kG23LODz/9qriKRInenokyeH
8FZPPh/cvVQU2Z4HsQRIEzrmoLVW4rGDbvjjID+659PhYJtvdRW8P9EfMtC8dM2Y
zljbN6XpShlPG9jupFMaBFzrJyRD+SK2gyVqNjlvd7rfoug81NJ2XCtt7zxEFN6D
3tQtpSruI4OIgpF9w0tSavkG1WrIuIrJboo9qxUyEa8pebPlSh2+x4VBPVUz4Q8T
vqAbEMEc8i/Lu/NnPsKqie7syzj7soHo3MFkqU07ZpuN/not35ErhPYlTLOCUm/u
5QxYAbU5sOjNhvVQ9oRHLqtkLP0kRrMWMSZaKUBPazwmF/+9zEOlZy1QRhEAfkO1
PuO7aQ65xwzbW13zeuFLeiJiX/WDlRHxduVK2Bf6IAzJ85SAPQR54cXGTj7MPSlC
iXlVCjJnw5VfAYhX4UO8KvlEvzx6fM10qehaffOwRFuK7298caki6Slh7rFdt5Dh
TWWtP9xz1TjXDCdS9HQ5qU9Kg7Zxy/atLtZbkp9vAxbPhcQgYWyf80hQhfRBMC6S
oF5cboa85KlMPZxjBQ/r58g5Vza1Z0hsmNHQ7vLkUkthg18lX4CCQ+XjjJbpIF1G
pOgeaewotLN+c1ZnDkvqAq20Ahv66Z67YSZvyuRS2LDW4DM8zVBfoDmmtyszOTYc
Q6T9VVOoBOhiztdXX/m/ldleWcMruSOhui5mPMDetyXSMJ1K75AWtrg3NVqb2Xpa
UoqDYfh+Zn1gt/C1SEZZg4yJ0xwmyQxJT2CH6rZ6KUtdakHYGvxaVMZ5RS2vnXRv
wnEwXiMtiswo+JNK0kHRgON3yC0boNRbbFQTVpPptCJl5KSsn8T+0F+dI0MfVmZi
p0rWFhJw5K/ILK1LD5L/fqgwdo3EUIVl3Vdwo7aQHKW/nGUc+WpHYawZb94nvc5s
DlykFqm8MFqNUMSqIFe5mWoZmhJL6pYK1R9B/w67wmS/dfcxGiJTUkTGXy5MKHID
uH5wy5O6ay6pbBbZbuZTElFYAdM4FSXrGcWUer/zrtWiS/IoIjkTq6t5zXb87iH2
0QiEqTppzcNobhNgKQfaJD82gShCzG2IPYb5VWVIEdTRi9K1VxOTmI5kf77p4YCf
Lo0Qruy0/G0OwOdg565ceJrlqT41l7N2KsNZ4SlSe/yHFxdSeHqWzzonVoEegyo/
nU/FQetRHV0c6eFI87ucMPN5OencIpokGC1F0q7vhxDkEZi+2HrRAxFpx5q80byW
6aBasVppU+D6aoELvbUkjtnZRycu76jA0hQNnDq7uR6MPNx9ePcY4cm/SyeyQcoN
Nx7QeMHJXB4xHBIk+iGubblMT3sseIkNESFo9ww/+jXdcRsWTmt/Si2lSgM+wVZB
YkJJd6HkKzN2+VYa7NA5iKHQrzvEBmwOtC8Lhylk/urCegfQDOQigCwgqWQzc8Nv
ssxDe+pZqMvXtlAV9Y3G6jltryITyTikQ1RxAYLZyEy3CFAtoiojlhFOttXWhFPM
PXPEL67wxok1pa4QdQSqHKU4VfCKqxDc5S62+1PItD8M6+91yIxf/mCCsERRPv9O
RaO6DVcHetqQ5ccY+jHG9CmMtUF2erc/InCXsIzAh8kpxCcuqICoUQ4bxgDFd83W
F15zy56pGWC10l9qTb7O628J2QKUndZuXNlRIH57wK4P5l8Voi9xUGmYPH5WWNDd
VmOx+pQbN5rO24ihHHpDd+TJiOWjHZ+vehO/Y26G4bCFP0k1s03yYwBOf414EPpg
LWutlnTzBYnTPNPetXsb5ZlEVQxhJQbcoIbvzSDDb7r7rCH4izhIEw1eP2peLSLp
gA/SH0tVXsw12u+l7OYUYtKDQh7IUwotkejCLzD5DHQgbzmsyhSIHk5FWDNuE7yW
IIAF+AniZ8g1hxjlwf3d+Qa3ChQ4vzKyrpSQmzMTZcVnDPxx39+4UmYc3kG9NiCM
ykdgaWc187+dZdFl8x0H/ME+fumgOTeKtSkzoSqjePxAL5rQ7TceCvUod7Zny+la
dpHEgxFV5cofMZgoaVsMJWCnTfOA+cUuZdCq5rWsWlHoMx3ZQQ9T0cA6AWIvMoDU
RsUGZ7XC7VY36s7kaN+FmMzV5HUvTDluZduaWPyDQA8a0BgZIpXCETbJEUwDzkcP
SY8dsSLC8Wv8UMspZhWr4PnQRCq7E3icYKGacoax/9YnSBeVwfh6u+x/nX+DqKdR
6u7jaCDtN06QDTD+ovvchtxNr+1bfvzVzOhpve5KQzdj2nks4J3s+ahEJYRGCzg8
jSaCND2QXQ2DsZSHrzbNcVCduMkW4/lG0U02V5Kpnxipc9YAo+m/ixDAKavuydkE
lumdLz6NhDyq8WMdy0ajmC7lBtttsj8wOzbpDzTTeupxs0Q0GWKqP50g+5yFvChl
IbvjhG+vjMsK75g2vxCNsncY2idJYmUEV0XIW0QCsg04v4VlvkJLpQuC7vb2g7I+
VpHi0k2xa3/wjEeRqUomoTBBaFRU8dhXsfDIIC+IKiH2OeQC0EtDrAoDaiit4QDu
rMwoZChadxtKpxhq5yZExwcxjvcKFJt9ms7A9JQgEDBXD/1mChpZ0iLQ9Fs/xoua
QlvHuKpVpkbP9MaQ9ncX4WC5bttKyd9wCFz0Z/AOqNm4fwVbbm3KL/BvgQjsseQ9
VUyjVqwN65YrsBkEim2oNjV4sOl6JjfOhW30GepTxO2IWHkzWh2W6ePEBZyILrH3
su/E1XG0GdQ4+ig1RK5QICmpmWA5vj4ASO7xt3pGIRSoDyC8ZkQwWuMOJIOAKwha
N8tZaToQrcZiLfO6AR7FDTVdxlpG8dC02UnHWFTrOdakUlp2OlMd/8LX1i1YRRE/
KEyNsI0qZ587q/6zLITyOlJt0nWp9tjfMOE3fB1EREx5C5ZIscuWWKXOSBx1lhGa
z+uadHKAdRYh6efUDCU4YH0VLbiNK1QNtB4c8+Q7oIqxozusxiQtAP+jr5c2S/Lt
x0D0C4Q3k/C/TZ+BydLV+gOuWu5Z6Cd7Gjnwpx+7/3NftZVBf4+TMoVivDU3Er5s
Cbr2RbQIrqhMIWN7mSs8arsqpEjP3zsRMTeO+n1L7i6lu+EK2hNVSWx2VGPBN+D0
iGbmnHgU2fHoPuXD97LEZ7wPOyT2D/o1l70MeXWFDxnL3Rlsdu8VcIoKp0rKRZbf
BE8w2hps4/qAJJaGXreLV8+AyId/VzSfl0td3YW4J20eXRwSD7Zp404zeNmSQPA7
NjpheFsHKuHvOCwf3xocIdxG+El1s3Q/z7L7Vu8/qrkME7YuIyF4Gts1U/JM719W
pjsKZ2waoVvyMAaZHLhVoxbY3GMP2x0EV1nL5g6p4zAOURL9F+Yh2IfRUxWj3EGV
qFF2TaGLIUPFvTFxrV53ZgF88EbYdybi48tj6fCGU2/pRmYnTsHIRR45qzzegBYh
6nfFNK6FPzg8BwANlEaZP9YRyuSnlvG9duuT59kRTI/dklYHSoTkBXrThq2HWGkf
8Ta5oV8j4q95kOTH+FJmO4fs5lbPl/Y1D3sVb7ykSDk3cIV5xtDAqo7B3+0Gdm3X
PpmhX/tiuN/DsTJKPfK5mdueCMEtmBULB8/mvzA5g8pfNXOx9yrQ5BWZP69Cb+ih
wIRSypynWn/WzMowCWHAshcZI63tc2eBcFdgJDii0uScLQh94jjCfNUbfRziA561
SOpnBn/FhfWWjD6z8hiZvxtpucvGyOeocR5rVKZMTvR99T/WXkRS9kt2pk7B0Lc5
8dGFyom2H7Yiv7/qTq1ZhE6ENOhbX6MVSMtMdBFoD/ZBHNIPsC0Hw6yDwCwXXjga
YADfTTjNLkP67H0XmlQ0Use3fzPZ7iUK2IEUsIsGFBwvt/WkcvdFt5YMXKFe3IEV
Ulbewh6kMVcVknVd1IE7J3+sPTsbprMb4w8DbDBWp9Iz9nC5ym8KtHXbuv60nJoE
rRe+zv5OzAHhT2CNhVhiIgHKyTE+xnwmkQvRVMEXGqDuWFL7rWSPGp7mM1gbkO4E
Zp2AxPZdl79JvJQOksX4pep1x2cSm4ry3SxrekFcIhgToSJMZ/A/cwMRdtbEgqhH
6tYbjE8nu9xglbvs8QVb4GrfhlSbSA6F5HzSyvPuzzHvutKD8UXpg6EynZIqLzrD
qLNtZ0xFF0IaDkWr1vrmjrbgo2pYAIfL8sy8KGqIIGXDeDDwK9lUzCo72EWjEXyE
S3evMNuMdTMfao1IIgDmuSyAvikmfb9Uo4LoaGoSL0/p0alwQUVga2QqCH2dTlm/
9EPAIfK3fvHlEIspVuy1sFz0ua26OwP92aNCdvZrH6IIl/sk563UDYPztczBPJ2F
zh/lxcFFuGRHJ/4yeVP0rw3HObqY3d3Qq91y1/4Aj6TPTfngvxxWbOwWa+2vAe0/
Msqt2zVoBeXuawxhx2PHDmIU9phA+n+bRpBEBnBb7cJQYVgLSXebNTbiItenGbEt
xU/MB4Z17ByPe7ZcAIaAdIs7gUdnPhzPQfsAMayYv8706/mi4meplARtX2DYdoCu
ewR7L0HdYKD66jrZTkm2yiKR5bWl5wutid3b3cJEmLxK8W5xHQFhhTEnaXQ2KoS2
1KOuYxFR/1nJ6LKDXHFGemmaf35V8HVXBnTMhtOF7LVwN/iqKOv1jfAxdYIprYj0
2SBb54MVCnX2vhXpMCVNCh04NFjPypRh9HclQxI9qGwXpTbMnYNjVVwFhe1GTuHf
ya41LehKcNbEvC0TagB/yydeuAT/WACssiJfqylnzfiOO25+33Dh7MTbrBJBIA1c
zYQLQ0QtX/AwwMbRaz2Iz2ung1ZxIkXdE2TsLDonKI13wfxQ6oKYkPzhfyIJeXyu
3/JYDCDd4fj742jNbrRni2OrQjy6rnK+KXtqQhGDE5Kopb/3/Lp906zOzJf0bFXT
U3sFT3KdEbAYwtn5mpX34uvJz2r+u1+R9/9DZggSH7CTQoL5roL9MEGI6NOQTwf3
n9kp8vLSIPmcE7aWx85vQA/giTxN9I/HO6KY7f4N0/LYB01sr0d4OSc310UuFBiF
zllmBmjBB4BgTIgAfJ5Huopzolb/T7MNeyPWYV4lHFmDZz9rBkD3VAfwmPV2iIT5
J2hRz1iqcbuUbpZ60F/0xb/LWrEMQIwBQrcFcm5AZcfwrbsHml6wrJwuzA5QZcJb
hBAyz+oKfgPqOo9qEKnGB/R7qT5Haq/iRAQX5Lg9hcN4DvwukQsdFrOeXarO/TwR
i3ObpJhvSG4rXq2BUiQW1IcwoNicvAUyfu5EN9jNhEh9bem3sSvjuefxzqBxpR94
S9uXd6nGcX3ce63tbHXwcs/s9R6sZlkDaYufCV+t0/6Aw54mtuiCvgG4oFEGkfX0
urGHjDSnJNKKbuFenbWPWQVWe+vIAKGiG1EzJSR5kfHwovIWQd2AyCBIvokUXBa6
0rJlXg6SzDQi5M09nWgVSN2FONRZOmVZKKtD5cOksgJj3wIlOCetgqq4y2dInVnV
6YhsHNDyuGmOrQNFumKvCP+cMfTL0QmXi9X89W8bwr2nV++5eqG2aRbYFgvvUfSG
f66dS1LOjzQ1ts0GLIPj1ahtcThD4ZmEK7sUhdD2CvKWkmxnBXHECGYJK1ZJuhIK
S6aMiW6sz7fPACGoXNUd6goqIt+k+4tp5tsxkAU+MGkkgLU1l0DxQFa/HN0acy8B
iedQ9hNs8hlSE//NxN+qAI9aWTsSr8Jk1ufLtQOiHozkVVnhHJMvLF3waSZwXhnM
6g7c/RLhvYImdGPWc8naOfi2u637cimcxnL18jh1hmO6aIjVAh+7bkXhpV/AiFw3
ildAjqbuy9p0ExfttG8sT994pD8M6/7HShoMjGf7MFimLaqVJRiCqRf9L7gQXjKj
ezIdvBVB1p1RLeaU+8DZUovpY2BJZI1OQt0KPLxIclo7uU0iBIUsq8HItJQQ9ajR
OgPqolfZKBk5pclXLWV4+8mW4EToKzJ4llw9TBrbl7OW/zYvkWn8Mioh5GoWVuIK
rJkwnGFVvVE5YJN03yG8X/bpLepYI4+cdweJH8L/N2ReBZQv3Bi+zHGxU5+xTviN
O660aN737J4mSxjDYMaQnNCmg1ErgTs+mfamBtTOLJSKO435UgU0Tyr5P3llsgri
O2rAn/MGfVanuUEzPSxCmVYlX/LKOabvCFzIdpjX1O9SEsS+0MygpKGTLfXMfo0K
ePX0Or8FWpkrOP9QGvRv9Az9ezf7SwUSbtIQ34XIvJ+LvEMW4K3kvAlIHeplGs7N
cMyXI1E7jIlBrPu6Ta6TElUrwenYj5Dm7To6rVr6dvlcnKVsv8Ip8wvuraTKh6CZ
ovZ7+KJZ3q4J0McYxwr/D+Nbat+Mz+Tqnns49i/xkS+Z0gUOntBCXNbJTa9Kg1/a
8sH1gCEUY2NcUc51BQRYGJ1MNnYqvEmM+LxdQUbDZGFQ43CGjP+PrwZnXSj9QGWQ
27Dh5XhSdD7RVanU9cicv/lBj70PIWUGOmC6ykXLSj02fJljQwgWuOJZsP8KVcVu
oxoyP5wv9mRpc5ba8V86FT8L++4BK+k03OpGvH4nC46xABxDYlsBZIOjWbGWYg71
47HqBv/NwDgwtbLrYbJhnu5BQndVBksKuheJF9s8OJMplmf7kNQD6HTMb7CZlIWr
UEYBflUZLbqXOOxehKvbwGM8HB1nOF8QuoPmafUzxvku5v7OoDQF5qkwF1Z43TWK
A/VvL09geLobCMJ/zsIWB65t+lGBJ1lJkMpdshmGmc4PmVWpgFi5Ilexo/GXkjgu
ZsocMaB4lugOUZJ+NqhSD9SgMfRJXiGwc1Hd0KNwHZHDZWaUMABFCom1i3qUII8e
ZBlngqipZPB6Byt6Y4bbxuWUyO7D5CYNJA2WV/lyhBi7vC/xufKZQes7REUsudiS
Waj7mK+Uy7ftoxA+mqt9JjVCSywnhcEoS4vMRxRm2LmOeAd+odkqCJxSfifermHp
u0CzYBQrAxy5jd0MlyvK9CxNvV+tKUoyI7TXIQVcVqqUeLB+J9WdPDgCzsTdmGj/
zasipM0IahfpwPhZ/RgleL0RUdrUYRn0k/IIOGTdzU+AEYlT1fKZLZ6pCQh9+UkV
pNE9kDidpEQDmD5EpCiBS5UNtJ1FxDQw3IdBFWvWYruOZFVv5XSbPwKoxn7cMUKF
K91W+0c6KD591QWFXZ59MfRT0tEPBg3xLfXUF2MaREFQEkDXDzvWAO8iUFqYdjd8
5i+nxRaEGgg9ZvJZap/ToqIdVvm+FvdcojkZELd3JNS0sP74SJJvsgiGL8uFB1qu
RjUg2UqHZZ5vIyDwFN9NT3BsUwuMsN3ZfY28+1d0St0wNzgB0Os+QbsIUalfiXmX
j+3KRYux4Y4nGDm7OosiXgbyjwC3XdLGgfvEDfUpaenUZDdWR8pQp8FLvF9y/6TD
Q5JsbFfY4Ek90O6lH4BUB6xb7rZpnuY6Diceh6GRMEBh4HlVC57otCK854v6sGOa
1x9g369f1RxP7ox4IlF96kqj2bcrgk5/0iO/0kQpKyBokOJEmoks7/T/0xszn49G
rVF7c3F4sLPuJerW5n9jrW6q8SI43JRCh9f3Ppvk2n8jzTYpowqtiJaluBLlAzQo
8OLXdXK3e5gl6NiK9HGFOz2N8jyNuLIkC9iMH07WC6yte4o/N2Whl2MH5hy91ZVH
e6soaX4/z01DWmZmhT/1v3jN93uFEWe56/Fcz+ToqlUPGUAPLXAaHRANhH/iSFRx
PvGOTgNTl1KymgXdQDiac4LAXzgL8qyt4BfzwRdvtGK3BdH40ekHaym5kCd0xAyJ
BX0TnwVHa4PHrZXoGqP1W0U8uCQlG/vqci/8xYvkHi8YVnfOTP/4FsiA2yBubRfN
+jjE9Yg68wQBxMHKiyIVStMCSFa1jmS5M9lcUSYuLShLglzo2tDoAaxtKHOgxsnC
1zk957NQSXuDtLOYsaWMg0MtVJi6NX60RjvcgkJFM38liNjAKq2scEbT5LDd7L2t
ih/DCaKJ423YNpvwEpw5stgGP7lfbadwCTCY9wl2h0iMtDnEioqD3BXPe6rNhlNc
W6EsSYfDZw1U/Iq6PzM+IBiJXoxLciNgehLhs/DeSqj1tBhlAiBHjysLDw5lMzhS
lTrCoBBe9VivfYghmYs3cGNHBnfkCtL66+dq8NnXSZSraQ/QGR5R6R4HLb9q3hZu
+VbNf1Xs0J6TG3AoocDIRrMw+jBjYSggLb9exH0viKj6I601igwc6G2ibgR+OuUt
PcnDR/x/NaVtB4E7GiMJXAyyanNCAAejSlclkAMVmr4naAl4ypr+Dy4VunY+rj2G
aMrE20QbSwAZ7X8ovS1ck1k4M+WIcbGPjhF5hYkt772UPARbyeRS7ubArYCXimZ7
0Wm/7q8JGE47dqX6vBJ5EK/bLXQtl+dNudU9haDbWGhs+p92MPmixN7SuG7h3rnL
U6loylb886F/0XQjre1fhFrPYV4Af9zWyjTBh80jCvcMhbubyTyyE5n7nz7UnGm2
hWxqnr47zClJSo9heY4JDBX68PPAxpYXVQmPVM6PCCXuxHdLx3uIsZ0BkFxTO80N
o5r88Iq06V4cUYygeA0mWFVYiIitynvnYuCnSUdakRe3+uElvRjyqp6lTVi59sb+
7DcPrX3MCpPP6kjpVC8tnBaQQaWzFHZlgLPb6R7gw8PQFg4Id48xGyi7XCplLo1o
C2F1NQoKp+5z90W4qqGfm+BNjsbsVLXpKPnFXBxkJv3wMYtC+HKgYRW3T9/KftfQ
/fBqdGwLdxZuFeI6s3XSnSCIZv6Igkfon2dxSuZjz3yr3z9I2jdHhEWf0++15+i/
eQ6CjzSnRnUFNoiiEWJsYPPyCQNBCPus91Ak+C4Fy8wLwJWoiNNYQE+XbK85bZGi
YQEhadmieTev44JmRRAMl22FYIc5h9vpztrsX9YG8l2g9Ktb8YpQMH1zKgpiJ/+a
NybMDymMdDceKGI8HogwUgyMmd/xyAbGahYxhPzA+8mQgWeHfvj0dosQmabQlP1Q
jx8smm7BQODngufeHGTwrPJg346hPOa/+6qExNNtSa3j5huVujUshdkFzWuCNvGH
2MIr249x8R08lhIq72d+klUFXmJdKkj/K8euj6pi2iT2LgfodtqfC/qPkUuB2x3V
IY7JF1iMcyh8XGewdcRSxxc487sZafCA3R/J5IS51DJRU1RnZvZ9/LVE7DBlZGCh
Y9V3ISR4OrmPfTfUYCKr2xT8x5cSgnP07bBjEHRZQD/fObaGb2iI14remVHKaQFR
918/EK9e/libu7BDuEjvBoVza3ouvfgWnSArH03b4r5abU0mDF21pGn9ns/U8nkt
wBBL2+Jj5E2MmHgSZHoQYs7h+Vg5xL4X5Qbk8wpRmmDn+JUqMqGE9gnN4S2/Fsu1
9n4sIkBKHEG3BWYADlIwYF5PP0s9tJjgTX4LjJU4LdQGUPwRyJrwEiqC67BlJLlH
fu3mupgt66DkQvjINgR1tFiwAUpq5fxBRHf6TLnNA9Fu960Zz8P4X49RJhSjMrj0
ZDFqPAJP0qoYjt9TKmDJHQjAaT7cwznwOCPnkFk5CqWcEXqE0+lE3Dfs8+R/m2EE
ED4cWZkU9si8CALJxyEPq0dI/DZ3jAxcDzTT7k3sQAy17KMRd0zcblMhDzKgN5OW
e4iNR9affznIMIb93p+8UUdz0FE8We5oXDiKjt6OHMZPQmJPlLG/j5h/Nk7R/ekt
RWtA7GiUbg5WH+EXZ8K5ZXhWS8cFvhWuWIyVaPvD9ykF2WZdczcui5vV5Vh+XqHM
AEpytt6w+6Air33tcMkErVQA3gnjNuvQ/XLy+2x/wjzntVbcjCrm2Z+AoiUZ2PXE
zeaNHy/8qpL3m0mG0rqBvtG5TAfC2bcrdxxCd2CD60saDwuOARkmSedKsngEAsy/
qqPRJ0FMgNpf0vActQCtRvGxqShiEtrU9XSx5QI/UdekGdBXg6NwIUKRkrGzF9ZC
riRs0066UXcjfW1BeuacRu4+lSKldQPMHe6Q7zoZOpq6CRh5z116mfA9nCzifjGz
vt4eIlGnTCjWbevq3NvpB3+aw/9HW4gOwkO3wjWjhVEpstx6d6SuVpVDHyI7JQqG
pjPbYCRRkYkP3mNC2+Y9Kb9Bm218OtgG/eSOlFAQZJdLbOSd3olHIBdEzV/uyoD0
kbozjq3XXg7LKHcr3JvE8RfA18ScrKCxNf2U074YcqSW5CZQCQ1qNy6IOLdgh2sZ
dHAuVTD6dIslJ3IKan3GEBx3bLIKBIGFsWiTCPWTAe1wwNOzVnh+p/CsdGHP51mb
BSWM/vhbgwmpi3+WoTO48plb4y/9hGiHHzzzFXXVBSf/o3vOK0otKjvxHRqjhFYM
jXhXA54BNpNY0ihDLrmebNDhZC+5+AS9osWgaR1weLIxV+YDdHdYEX14LJQ2CEbW
SVRsSviJYyu4YIqUHbG6jL4C4p1t4+cqJRTnscySisrUqOa8o+qTlU5y/Cs9Xaot
WV8QTCgIvhhSBBT+Oi5r/usp8gL1QyGHO3wJZP4IxvAhsCqjfD2HgYVP4BWG4N5S
zIWA9RhBf76K8EceZ8MGRu4SyJl6V8OcGtyaZkJ65bPfxVVXsfnUCFeKUeSgfnSM
lHjsOqmje5UKUBpbx88sVu8AOcGBY+9WugbFg2osNYEyTVg56N6Lw/yDrXvBuhqV
3hdkHOdk4i32zTHK66KS0Y3qthIFMOKrJssMnI5RNEQgNicB8/Qv9DSOjWYzkTkq
Fja43p0T+gqxE230WFBrgJD45D/J1JdyPue1X5LimfArPaS94JEyF8FRkaPr6Sy/
x9t6cBocF+q2GWBRE5kFxk26aYPniFNONCHPxqikvGal3QD0u50e3hATxRE3L/RP
35Vgp8hCRMVP2mZSnk3gbxE6ls4UyQ1h0hIn+fAVTv6yTB+zZvhSuWwzBa0TH76y
RAqhROS8yfaLi4zkl4acTm89lw3TCnrnt3VhU60toOOfH63+UQSke40yYTcpzesp
9MjVEwOeQ0SdbL1P9ZDcmObEJcGYv8+hpKx2V5ptDGM9pIM3nSkUMYY+OMSyefLT
tCVTrg0K+JorbSR26UrqVLIipRpJhoK0FttMp5Ytmz9/V/7hqhd4FcnbPuQVOI2Z
YxfjFbF3P7K2I7cBEG4ySkUvSyCYgTL6ULzct8KDWaz/pRbfavD3gjNu2j+l3SYI
UEqqwv9nEu1s/ghPw1+D/6nz/f6/UwSU8g5v3/21zj90u1G/1MNyvmjI/wbYP0Zb
HJg4GJ/rnL4b/56Ug72CdjDsnnmk4rtAjwyu9d2imRCwFm4r+VDrgWzkQKi1vt+m
tApi1TbDXBR/Yh62EOpLwjUeTZytENbv0nmS7dPbd/wQKjegioS27ytZhTubicWu
tHXBj5vISvvDQwgVW3OxusQj+9ap7A/K+kFzkLI2skJr0MRgeG/d0rFMokZ/ZgQ+
HWhFAcDKZK790D6/AFHvAJOLpICkvJCmk8QwBBRwdwLpXsTNhBAyM6iHe3/FHpNt
V/MMLwtmOxXVHMoTBSJegaU8MP27Pcmcaqh2JWBdliX4jurIEeexCsmGMsaS0SZm
Lw7WDe5o0Kx2p6ZKZ5JY5It2GFTTcIZBFF2rPWNvjry5hHbLidFy2O+lRqjWl/NL
J1C0DurG2+AXd6Ak136eqyxNwpNgTFD8RnOoNHKWfxfE69lLfMaxSVOHPPSBuWas
bD0JBlekBuS572QXH6yS50tqIIw/ys+nLB6lWFmNmWgmpfxHtnXz8Xu+qVd+b4xH
1BndEcGNe6hkM82qkOGUpnektubVnWS5WTD+Ueg74C6V93ePhEI3kXua2saV43qh
LhWq41DvWFpTOisDzXiIgheYpEFnDyO98VJe0MH2u4NpLLbca4khe+KOF5+h+onS
TNUHdLW/++Ypm2CPQZW2N6Dptvu+/9vy4g/6UnI/rxe37MyN7oh0CYmCxa1XvF/B
raMDnunBJz4nSv4tIU0UFOE2/sVQVGtaoLBflyRsCj1NQRUl5egsu9LiF7cAYv0c
OadiHHHt7XI2SApGhnJ53XFPiRKaKpQb7ZM3BDOacwiJ5FuXwFyfF+QJEzAW4k0L
BDwrwNZd4Tq4+zEE/wJM7qkyQbbpo/Am94bmXSDMeRaC1bGnpcHlmadWuvFIjbu4
0HEpyuf5jndXIyq3LuZhIS5FT65cjXEU+UMcH0nyhAAF5fNQnWp0irj5yNEdb9S/
e0rphqls37SxN6ed8MM6xH6cbwG4Y9Vqq1FkECtV5w+ItiNsAIb93IA6PnS640P+
i3KJktuMYEK8j2d/P7/TpO19uW2uLpPQzUaxL05ldrgiY63RJ7WT/OGPVlgB6XUd
3aDB0bptbYTebbZtQpLGxawtDUMvPdJNFB9UqVw0AMZizU/McMlffOfvg8fVyQPP
KK67aUOsLq7SfHr4C5aQ/OepSE3r0W4NXGzHjmzY0zbqbY5402a6Kyz8xTbViRzX
IjuRNkYX84xYv4Or61oJxMyYhzhw2VtXAlONSRR1YRboU6XYAY2/mzs2AaO0lQCh
5Hkry4pqzAlC+pzaHhU0A1X+3WdI6diTZUbdXfq6J34xsu/2PP9JDzaYLzdbyPQs
vcbTZ8UrgWfohwRgeKluhyGhzHR/JDYN6gUyE2/a6PeErLd2yG92mp1lB9eUeKyN
ddjSG413CBE+Ea92JDwH2TavgA6RhCsx2TnKC1buhP5U5mtedr7RWs7IBLsNzRXJ
IDBArms5zPTvVf1+9L8a8Fm9muQ9M5YpaA1H7LxHACX2S2UVC4CrKWG7VEBxVuCf
WWiU4rpjC/deFMbdaYs87MVse63qfgZBvfELfk3DMUvb/lFAF4IG38zw4/eH5XX8
9uEesUx9pEeQF3g/bVBIe6crqKVpfi60xT4K7jJkNpaLP/I5hWZqTJNIIkmOf5dB
0YF1i6ibYaYVQpIjA9WpgvZ9trau2S0cRXn8kpVKMLKva2rUH4vS3AjxlbqTVHiK
+c3RhOxA71R7gtPkPf2JYScHRKvkCpOKcy6c5A/y0UmxnIEkmYu15ly4Q1MTbH2t
oYlbMGbPg3IyBS+Ud15JqwzWsRmyskAzazkYg9JHcABpTH2TlWuNotaWdNHuXPwU
c9dUBciJZucyQuT++p2zckSk0Dsjv4bjDxXtS9XmgOSeND4Hzif1+WvVN/lJVr7r
8BF9dnMSPEeBDlH6Kent1Xl19IMOTJIKDXnc9zoDxiFKbw6VYDrk182PG+Qeu9Jx
E8TJmfeBdEZC7aQAxSANx/s1q1d3vhmvSCVfmY5XIhqLCGGECFdkmf513uX2oGFW
/xOmPzitgOnzTSS28OTsP34dOsMx0ail1RZ33hGdiaOj8GIqPJt7yb/pEPeRAGQC
boak5M3LkUoN5E00RrhhUxaAPC1Y2OpMWezcbcHEhpcL0A163FxxV9DNEDQTVaf+
WvJqROla4N5t1UKgqfUJgOEIDkUsyvkRDEw4vH7t3ULJoBJl0QNOZfbNe/IeiNmU
3EsBVvwv0IXZrXVAD6bH2lS0isSTowfhCMFbX6OsVIzPJDQbCKptkO/D5bJ5G7vw
/+dyPasaImVtGyRQBo0babXY7hDIVGBmGwLR3wNV+VEvci9MRm8+G9wkdGTwl15I
pQ2B2+4BgskPdbVKr3AbnPuK2jxqvYsRpnfLabNf70IHxI2Qx8EVrmBDyKjziQ8j
YBshJFpcNMqBeJt0t5hilj65tg8TL0FWMCrC1BtotCw8E4OQRzy9rcFp7gnFJbW9
08HZ5FbC71rHVi8CTUHbomZFtr9ri5DYJ0tKnhD45uOTNbrPRcRa/iCFvYZ7kRTQ
utCj3L7lbuan5QNZvblsEpUCDRLobXC2afv8TDclg9L8bljqlLYJPflybHvcePas
yrkPrTbbON0T04xwpPT0x4QHue7PtxOWONgQxecfitBJcV6paX8RMmfl3oql/8GB
r3p4tYzZVPKWUsh+Z3brSBu8LFwb4GClhMqk15AFre7Lw8Zwqpl2YNqMhNXAxhMq
J3+FrLQ1FFk0jLaRDfEPUMviuWG8UVodLcuViojVYP/avQK/PFARBSyqN1/oBNBu
Kwe9tNGzdZHqqthREt82sXqsw2Zex8eN0J4sLJfV5+52262jf1zrh+ocw5NANIqQ
SNVP1ZuvWt+ZOIRxX4Z+waxqoNpworGLvw/BlQOGj3e2UzxIF6NDtXl1lFDfVopH
DQ0JPWfbjsmdGEbt+Jiypx9OLzrUSfs9JvoVQvkVd15tbZ45LeawiR6UH5nCHLgA
6TuKAa53giX/XtX6oHfS/Ek3Nl2coV7me7YHdwsRwd/EabESQqSzirY+ap3srLEU
1nvtvVtClZ/cd2nHeM/wCBlvkaHeNv7kkYufkRFSSc85s/iVfanLkvNIzIRh04C9
oyJi1Ep+C9nwfITi/sx/DGhwUkuVCCPXwvXDSf0fgCTJuPC4YXRq19SSjwr1mu9a
8xLbjIS8iTai+0VvRhGKUqz9iTCa71e3QbNF9azixFhF11zTMbHZdduZlQQZhFbD
viBaauhVzNHl7XjRQkKTJXBg4gecVlUEg8MWElhQtcDR6dwMGdu471uiQ0lubOCq
CCP3FD+6mHOp7XeXCj/AJi2iHc6yb049LnO8kE9dtwEYfgwOoaCQehp5lI54K41m
IQKov86ikrwaGmdnx1lNZODN73uUewQHlV5iUl5tuRri4DS6zMF0NnaWi+49GGZ2
KZsWBileHJCbHnNJoh9MmzQ8VlmgUXfL3v0bfUjFfqvHzF29lp+szmboUSVNm+UV
3bc3t5/6JY4NijuaGrNIWKFMnqXwLNvVrIVPwl0gR3iqT9cDoKgZ81PsYStihwj/
Br6hKYgBIgKWOuzVWduv85cf3dzi3lrtGkgs1vG8NgLGj66wkKkrDlmaOCPlPz3V
lGRVBSsj6yuuIZdToAFDe+3k/iekYYeinKjsnDCxCYloRnqccG1npMuBVKLshaxw
UrJe3LJdSca5IpBIQYHyG3maSpX3R4n5M1+G70jJuwCDcs49mqxrTlsGziFSIpTV
Q0x3+0CZ0e72ZmHwEnahV45KqmlcRAVy/ZsyqZSfo07oo2tAQ+pOr+O0kgPTfWfJ
0PC/CyD7I0yaVW0OshnAfTImmI0gxUd1c0wfXLP49m5F2J1mQhHT5MvnqRwLJ/9v
mzFpL5G/OJA8sbnnHKQmP4wmzkluRa78I3Ly+zSc0RylAxzYFaR+2LhrpAOpNwJS
lr4RMXJt2jzQO1Zsr46LAxKMjOsjJZh3zYbt2663Ftz8I6ITH8WfDLwnAASM1PGb
0S2E/seMMYiiZAr+RjMJT+wp5TjDJemA4VlUujkfNNJj1Ucf+2G59w4ZlXGaxEiS
SBrLSs7hvraoi6gVw1t/AHL/9ljAY/YLpey8T1pm+hNWjPTRaCypPcSsn7sNwuqc
MC15Kcyntx8XmdpRrBchY1e0bl8YV8g++v0X5AvEdCEf6xDWfiE6SCz4JlXLWDkS
azU0Aym+rfFHJXNg1Eil50/haYiRBwZ0UculQEuygrc5r/kQMe6Y+LSHNJFSbusD
Z4bCfXvfayTR3vyYDbG7OyIgEiAHcU6MOliBJCu7VfRi5W3udShfTe6Vx7ETr2r6
FsqKOR7bpE1naYohY1FpXJjolvOSRNZQCgfGLZgLWyIeureLZoKTJ1zX/ncsB8af
BFSPrYtN/r+1crLkQq0tD6vpVAe5J0lXtdCRL2a5eJkx7wszQoO4cAxUFiAk5V8P
/gLU3Z+PmsI3a0IhJUv3pq4g7F74ROlJvhx1lN3sMAfarHwXaMtQLEnYjfbYUXMU
UPo0aS3BLA//G2wFkKKbHVAeqrPum8PCS8JrmTadBeyPOW+FdJKtl7kPJAZdWWXx
HARdOMGUGkfsQDYr8vM5oz3Gk1pwn+PEaOAr5xCpdNSKPaxzSmUpDsHa0/SxjO0V
yoB8bq/K5qNkb7xYEAUca3ID5oWzDLefxmnZ29gOTpLhAyLOreW+dv/GuLZizFFy
n2KxmEgGRL2khXrv4fcvzqq/35P/NbBHoGOKytdKybtoY0xSKqWBOm4Lfm30u8md
fzxRyCSh8VDWrVEGOZlXFY05tsmTv5Sg7SdEXg5IC21dqV606P+5kJtNTsGa3tE0
PPoxy7J1g5JjgBf1ureubc5AIJROalm3BIeT1lD2gdKuruKKxM4+ujliWCq/JqOh
eO6K2+Fek0lUGenyP6pLcS9a6kdcTo6HJG+Gs1pp27xFZDdmAfIreVaDKoxP2YCP
nvVH7TYLcStQ+/jmNfbEQUCeoS4cij3+rOt6/tioJXkhrIDEbbh/di3Xnji5d4X+
DfNpZru3bOqF705YWrMaOhdSHLiNrtDQ560XbqqqmL4OsJ//G7ZzsfGVTIJst5o+
zKpczMeZLbFoGATi/zBR0tAtMHskv+kuMBW9AkQZeO2syonf1/FUHC0doeaYfj2w
zOp4XCDyQMYFOwOUG79pXF9Yc3A7V1hkuW1IYsuTg7OD0laXuK7FWFnWUbjICns2
tk3CjYg8wRjyJl1Qx//FIZUnRA2s3LxiCX8WWGit/OzsHFrLPlxkVDUNpnmV31P8
qfZ+/YtqYcagIRgnTIQY2SMeDwA2i0aOCqw8UQbyYEsNFJ5kaNWQFfIVKIGp8jwB
3nsXHHiXq7/Tpg+OvUl1vONLXTeCtxfMg7bZtg3DKWl4j1vRUkLjp9APpmMH5xT3
S1fEmXpvTJhhqQbqRffh77uYB3qte66m22e+X64HzSNyMfs1ISNTbGCgBsG9ktyB
oUv99qdbCgSFZtKWQ9f/MEdYNL+S6ekSmcx3xrbQwsaReN40D4KFJsiqm++kT9H6
hBLGBg7IFhG8nQslJkdlAAKTcyyFXdhEHwrjjNvskM5zLSy8LtpJBhn891VMe3kt
JL5+zOLp7K24Va5Bfms/8vcFlwqrCHEkk5JW4hxrTYlTTAQWhxgjvh4Q4/341okz
KaMHFS2+BnBCMLnnQQb1SPWNFS0anIRCne/bbbKy3a8sleK15pCj8pT+vpiLT/4M
1c+HX3MWDULQXBvys4Q5dUUAjYK0dp0vnNxAW4QS+H3inaH9HXxkPdUpHttyACqF
dAQJx3O9ze6t8bwSMb6v/n1vuTd8EeEPg3ZRQEYGIhdPyqN8jz5b43mS89Xef5+Y
sOoDbdCKKqaI6e6RQ5HlIGfgRMTmOdeXOUjJG3J6o4pUlfeHZ7qKAvELmg42+kWF
iPdStH1BRwb/IIHfbLVdwXk7Iwo99IDVd8Zy1nMASf5pFeJxMBm+MnPU3VL/6PPP
Yw8idEBcdLGQq0jwJt9EW9KqkpStCgl5pbrLf6L3fGb2s945oohXJJOxgBZYRz2e
tJq+F/m0cbY0/QwpJbAPXqixAHUsKRQC6HuEM41jedpkj7MmRfQ3kOssr9E2vRh4
hVkS2laDOZVvizlvzOsgW2kUtMFduCDJMsP2UaEOvjdwixB5xxbNjJJqUoYtg+Ca
qkWPZJ50HufKInuJlrJfTw7RH5M502rvPQlWe5X/z+7KW4BMO1Ho+0PmS9o81ANR
lgkfp3pONgvjDjF4DKQJgh+w5tNpt1ewuhRJdsZZLwGH6SxKGxRPoCaYrLbwYPWV
IuzJ5NdCNpSmacLSeffvUX9My2SCwSX9fep6sOwmyc+jMzuOWvcYZBuQn6Yu4MPI
9+XcjJxZe4oWEKs0gHqrdWO9uFNSH3lmvExJCn3eckxL3UvURA4YJjBnviThWnXb
WgI15UJVnYdQsKE9ehQcYHVnq88637d0ceQkFgFwHaJlVkB8NVCvzlzUfQ391Ji+
SgzUvS6UJH7FXVtNOd1CVSwD3JjnxH8B8cVII571dh0m/S3fED1ryK44MjnsQiFt
x3WapJUKJdngf78DWSkG6bi8Ztq6o9kWUK7/VG1xkiLZmqPqT3x8boWMgW0LptVl
NeSmlcQLeLZji9ro+Ga0vZ6f8I1fMYFZC3kn9F7MXjJlYRRPLdBoFYn8m/U7mvlC
abVIY4P0v3HAtQ/oGHo4od9R6FdmlAufsw37xKWOHtWKC4NX7VeF70opKZ3r0VcZ
1wZmvICWoQxSl21DbalVde/O4aoAPKllXK+QiAZF45D99c8XqcLGI+dqTq67VFoA
byMXUUUurKswmI4iMIH5MBrJthRSDifE3ndjJo+Oke+FrA9mquazZ/2AN50KE4ZL
GmcYj8FUyDlQ8/HuTzu5ggkePf4hCz8HC9LZLcF6Nf5IXtyIdccTzALJgBRnyeNw
i5tuCu5+J43c9BetizQvcZg8j1/Mold3NLqQKS1vnNjZ6JgBCkLQLoM4znvYJpG8
/8c+W6/KQva+6gs9Zat2zi497xOqN6vJPmLckWdwFo8CoMjLALS9gfjDWojHHuRZ
HxrTMlBpH1ZmFQtC447KDJDAY4i2FzwPp0vcl7EI3FrP2gK6lYU+yMz2/U0uGBYI
aGWKmGn+Eg1sAIEXz9gduZKisDZYm6yxJOlrp+jCWsRlGJ98AOrUBgh0XHxUo2Y8
nHPHvg1NTMlG2R/l6X9EkcSl/nE4JigjJNk75+V8xC9XsmitXpe4selAa6ZhyNOv
QVEQlDIWLuItxptGtih/qr1jnfxJBwXMLaFLCSm3tKIH2eNu7ghV0+8n64yIsDDa
xTvliza5W+WUdqtqlq7syJatIsiDuT/yJ3YDNgIIkG92rT+K+c3zlnRSeUvXj5tW
fQZvzXdmHKokrPS+F3H4kET7Kk6HhJLK0UZJcCfb9PUn3ZqfPDgnOUNHlhaBXT8c
7DkXhd5nxfI6/+sKNiYjSQ1yaWySLG+NluzWXrZXmT/V69dD9CGzpOTPiZE7adba
fzn/e5f9LoIvioQKrBSHRP9V3dG6wBkV+2wqoszCApNCYd+YUZqutefg/c2pzeNN
uRQIjtzjYdGh7lVwCsWpb4Pqlm290Jixkjf2PZQj5AN2DvK3x79ra1rMA5jX2tC1
mzLYprgbrIX9w92sunF4zG0a0tJy5v1XsQ3Ds0AN3NAjZBVqUQ253bGO4AIzKe0i
6zq51YIwOLEJ9XhJ9t2uJjNoHwQH8t5oaUU9bVQW2ws3S+x5fdPq9HC7EQ1f30lK
+gcLbuIfTyKSTM0G9/q9VV+NwcmVBh7IJiSYDez8Z2LP4QS7r+rDB/VinlAgPRpe
7NacK3YhuVvLYMd7AU3sHTj94UdbFIvjqRjSxgwjcNO4S38hi0dT+3MtvX35WNmq
cWKJDZAfAXda5ReoN91Sz9g1ygBhvCi2ynBBfIn90XabJQDbtACaWEcsgcs9LrTK
YmlI4YlCHUWpe2qBsgKgjK/cePo6Gjln+Ftdk4mLfgZNMVPOOq7d6XOlMj6tTswO
PiYvh3uhlXZ3pzrs2+n+5pBVbfYQOgO0epccoROFUw39OsuMwYN+dllnYMgzNX4X
mqdG38qijChrAkkVaE4WrtW9Fs69gG/pMkolwdatV07urf+F7OhgA9NSuDxu4lht
QUhUlHf0iP55VH1vj83aW1d8AYEItbmKGTTZmWaKev7s8tNm+JkfwXuTLHS/OI9X
sfMRi7dq1y6VHm+p8J+Q0g+mWQHZWTo6sJPJZC57asnS/bfcaO0b0DsWBhXHabXa
/Mx5vr7otzBiXD9PRhf288+vwJVKNh461Wgcq4jGYNBZevdNh7Q8xgjjsmRXWGkQ
dPqACJdcW+c/QZa3ln9KoOe+BhZQ2chNxQPusqW2AL4AyUVM/g72j7HJP5Y9H0fZ
PlU4nIP/m4dadw4QMBSRuxxaDIAqUe/T9+FWAsOikZPPFcmB4mkwVHvJhljaXIgf
h7KF1kyIHna7RitoPQmPfDKWqyKhdsOKbP1yx33Z2rThgntJM5qtc4fMKlsWoFuR
H2JjDxNA60cXEQp8m0hxNMVgBLdVkXpBVmgHf52xo7FBOTjcXAYH4ZDBCfbdhylH
/b8FPK8DHlti6Xh0GpwDc/4Hyo5vcKf7mwcuYiK6hrzTwXwvb5mArh2osRXmPf8N
BANC9WmYk17mh42HVax1uX9iLkvQzNQNpDb5yYpdANPHve2ClyiOAtxABwX3GiD2
nROnEoQZcdnadWBa63zCFrC53v5rOBy+LxBKEFhYzXQOeIVxh2BN9CR9JBmm6NL7
Nd2TpoNJXc+UJsACwchbZH8rDyFlEe6ld4qsUnHSVSNpZdpDp87engEUvxHL4F8j
7cdmxJmYMqSzebx8h9WCNuwzv0GzmWwoD8Xc/GchnLc5g3cMxQoMZMeSDYj89PWk
TgpuBoclPgOUm4oxIadPOKT5j5mYnDwaOHkU1Cc9VTU09L35Ym628lG3gghVbaFY
2aHz5cQh5q+dGOU2kBM9oNHdl8gIWsEccTYtkMjya45/z5JIw1Rflcp+bpVy/kwc
hp/HRM7cLwex+1AVK7lgvhn9AZeHJCR+TsRamMVuCcsLGRJWtUk6v7Im0jJhzZPW
xiBUGmfBdBtWhPFHE/Bcq+NektqefcFB3fbknDGcdz/NLnFyFlHU22EDXRWJA6cI
EB87URjONsXOGvqwaIhq0VT6CwrLU4Ukq7YDU/8x8Bfld6DaitiColpeVS0eYxzN
hTynqGLpjRDsk836H09cUN7klVGuYgyWvqtKMPtFSgjy022AYHeJYxcNXDBXaCy1
fSO2YjUwUzeRYhxUhS+KBsuMMWpTQBGRkk4EN0GNhf6+9Rq27LlxnZG4ishxPfds
LU2xx8ZDAGWuXF6aixrxlRW09ySKgY5WmeHTj0lNmpbk0SI1K+l5ZlYKhIboc9sY
gsT3QK91WmWU1w0gAbLRSK4YYLgUQhtM8lSk+s1wRO/YKviEvTVUaNyK8ND7gT/7
brckXR6qslHC0xPD7NFxwyi+oe76t/Yl+EI7/mVmZeOCWbq2mE6EwwO1G3VcO0Yl
jsnojNDfIDMKSCotzJhNFra8qI8KrtPW40/jEZGvGLBVR8OGMF+tcmu0i6XOmgBU
wPqlRdOnG7Ih6NVhuyY2xdNJN8FWVBpNmpNHyF9GOYQoEWU7pEHinp5xkMdbb2MA
bZOD03nOz0CYmBvyM+ylsepaSKs7brTD0u3NKhm0MZGGg+os9HQ0l3RHzGRP5ljM
55zrkE9jiJ7Jq46T8qnwYSVLrhwu9R8v1uxE6K5+2HNmihiutm3SRrIYvJ8bsqRQ
iMlJP/msF1NCnKlCq6jwmXO0D0zZTXL6uqkL5fsl152xlSTCpzxPN+og1IBhkbNK
51t3tCoH2+loAILQalIzJ8y7ps8Vod0PEDX+PVaFf+AFpSi9zN27hHGjnMLgnl08
6rPQqYN3IKENGbRdxF+mC80n4DkH6d5IEMICNUgN1+2eXs0kXFqcvY1O7ojQ9cc7
tURCtwWJD1hvANM8wZfyckY+FR6TSFIGUDhx5QtB5V+UEhcDNXJz5v/xR8TYYx9d
/Ny+fS2q/RDVaYvEQTn0uIOIu8kudFAA20bBZCz1qNtBmNfraQ0zIYwnN7R4YB6r
8qS6NZCn8VpDPf+hJ4BdoC9ewMI5wlbrlBN516LqbBU9mon/wnejFfUDael5cZaJ
CTOdrFcmoQfcx3ka9iHtFk2H/fZOKqYVScwFv8MmQPjINGQAuOmLAltPKqujBiPw
uNTEjV5yXJpQmMmv/qf5pDVz1AjxoYLvSsxnW95GUeIod59qomtiukBrSDMCr36g
iQe35NQANCS8Vc5sGU0A9ANqDbAoWKEYQoPlkdnKtZXQq4DiYQHItNCpAxPOtbIC
gMgCbrvPHPNbmtPvxs9+1mNLui0hfd+tk37ra7U9ggCvypf7LsSutEQqODiMf60W
IP8XfR/MZYmUnXiVDW1ITKnYDwGZKgskCxutXpq+y+9G53YuSan5yTiQNKZ7koXG
dFa8y0rYzyeWqKKmLOl3voyCCm1bjAqMCCWxbTWsSKbibewFWXspyPhOXfB9Z1Vr
O9ajNrZG1xluCwoArfa7FuUfZP4gCEm6b3MZTZbs2dhbgZUIDmoElhw/E+SQAy4O
pGN9oe519Jq4CvYc2tHM1w9FjunCqBEJw8X6DbPUIK81mqLRo3dCbSTdngDcso78
RRgJOGL0o2gH5rhX5+iNOeGy+1tlluqfv9+HzJbpW3UJu1fksewYB3E5LX8W4OUE
5PdVEmSl1ne/YhY02e73rLb0w+nFHDW97lvIlyOBCT68xep1PUaZAD751UqqAEDb
pfibQaEogOI7sMzVen8aPhz2TGbnl/oWMuAe2FUx+Mm5wP8BmP8Em+2Dbazuzuil
ZYPxPg++1vs3h2DWrlR1axqknIMwJiIeeZNkKB8uhYG7WuS6q8xpXX8EqxYB7jS0
dr/oXKvRtUAFUcCd00SkajN+e97rFotXqZPxQcvI6ap0lQuzNFdeT7x3v/TXasWX
iqAscgf7rDWec6S3aUcvXj8UdACKP0lBhRqe+FkZuMiUGi8v/lmVTskUTAvzhw23
I3EQgyybyQ7yaD2BEKSX64fXw5m/oOyidaoMPPdMZHkKpLI2WdyoM0StYfjKOo0P
bqnA345w27T5Zm6KBLeKxR6vhAq9GUQDFbZ3TUClr1kv+3jleDiwZ+DCRI2BkkuL
rdxDUdL4seiST7YiA8NGpYkfo+SgLyVQ4GWv/FVBazxh2kWLJy1D7eXeaMGBnIDo
nj4y8p6I3jDWQsR2O2gnhg39YEPLLj5/urUSIdxVNp/RXuAbhZ3YTnGklVex+jaV
H+/5kkNdq7MxP+Tcn54Vyoq14aHppGqNFV2mUA/yquFOC8g3xQiCkywRRcCx18zn
IcuzmKchY5sl3ETmiWFGnHQUS2EWFgYHdTlfv1p7Lf0vKrmgsylERMQYl5saJ5k2
4hPjkur9I5LdGMh+kJk3NbF0hJ0tgjBZAxhZxEhX9r2f7FhX6zv4DsWwby7IVBOR
DKP3lX1liyUXPr9IfSMl/pf4Bpmlzh/1aEuCYFt49a8Yp4pJXBqypMZ+6E5VphVx
i20uKCeyXxmD5xb80xDKydMgXHxEHo0E0YojiXnZ6j+YHu7B39fS44ih6ZlW5hAU
deESBdn8mR+/k68z+RvHhLP7pvBGHvJRLuR6SNxYiKGfXgYfa+01TzVezsIjEAMH
53CJ1OYC8w0OeK9limqEvP/7wN/jK+1eoMngfbN/+eJWcW0HN8ciovFd3JuOZQ1q
5fpEW2Ls9cW0RSv7sVylRxRWGXL36TguTzou4jbysQmFAMARrQYJkvNTFNzaF6TG
vhamE3+vqnoZce+vaOYJxBrv/XwmamELT5w8fEJgZyXbjfqUVoGPIplvcQSksOH9
h98pEwbpjvLRw5gM3Fae79DP5stzI3ljXUMkhsInLijYcV0o+Lj7ifSeICrktVa9
Q0/uCowTLa95VUJ3Dh5+tYxIYHI6aXiasLsmhQz2L3BZrUUETc9iWSNIJEuREsUx
cr/XDV6kM/O1rFALwMPlOctYbcBj8gZkuAdnt350Iby86W6ZyAnfU0Ds4m0kfW4M
5QD9iJhn7p86jTRttVnuns5+gX471LHeswL6HXgGy0QytjJ8RXVmZF8DVT83c1kC
S1nPdsOZVljyLkPNCbkQooaHdtG2zALr4/OShNgscKpwd/5iydOdWzMZd8KGJmHB
FgPLUry1yNbwsZQF2MvBlX0EauQrKqdbH8zJZ0kNijCd17BGSxcOxdYgddxEsBcH
xJiBI+UJOXCVhTgpa3IG/spp0Ao1y0xLSlFu6VE5iQcevSfn1H5slj2jit5ajzcU
UJIRnc4pCrnMjtsyDQLxXXnFaVcBqNYkraRXHjDirLrY5A/iyeiHEzbzxM2BqMhn
JI2/iMlLs0SdT1gBFN3tEzBcpvlX4GGjWnvXkRWgepdLf1cq7AH545b0DITsf8AK
K5xlCo4h8yj3NRFczVw9SdcOKjQWDPmSahICM9bJvm0QfYRGKK8z5eDX2URV92qA
jfyl2Dz6BsBYiPF30J7mywdl06PTt8pigPeiZdLKrwn6MC3poV6dj5/i4s5qJ4g2
y1dNKTfIRgTjq0xABP5j7OVbQiiKfmmpESN0KCyybFcyt0g8hcaL7fIy753T0M3K
3JMk2WJdxqUCboen6/BOQdT2xiTgYUVg38W3dl5eyHpsJfH93bcy8aqX31B9J+tZ
tIRaXGTSPPWaPqt3CxhocuGDzxtWOv3eqghljMAIS7m86WLkAD1+AeRm+La9sqie
zJ1M40siHw65nvGIR1FzfpmxlbIvaETKdTZZU1kSTRnso5Z9CL0J55k0nF4DYuOC
gE7YeIvjPPUazjoFSedME6xbnZKKJgSWh1DpM2PYqwOMjdeHGLME2ZVMsH+otQlY
HNvzO9x9slNCH3GWk36A2w+z7JKnecNjPYdwSEk840nGbi+aZo1HU4sD57o4gl0n
roeD5Q9c2Aeu0ZwhTzxPqcoNRW/m6RUEJ/J4PhpTeiOqDTPazDWnSTuX89v8HOa8
h8Az3ckgwJvApeUSFQhDiLEUe+p799fC6hi7Ys82oWZHZJH+puR4wtlTHgiGnHaP
+5Pc4PM8aoIme2EDAGMqJJSgCmFqTPPJqvk3sdNtzBIq8A4wzDj4sFZgGauwiwX2
UPPq/FzDp1dZ9tJn2zW4CIh++sn07/broEmFOPcxodefilChqayIFEfMnOgvUnJm
d7T+7yOFME5IG5k59lrnRcRt4VsdxNeQd8I6W4vn5t3eDYLh2Knmh92ISZ1bKxmv
EEBdxScBV1Xwb15hLDI2gBYVjDKQLpr4r3WT00xkR97uJsfCTCNcocxZTC4/WOM6
GL2rqjkkBWOEle2Ajq59p+a3SeqNxQ8zQWjkl//a51xmi83Zcb2O2GcJh5xCQU43
ZKB8wCqb3gpnSe4mGXc3LPPvkJV7cvN4JI4ozUq/fDt55UQ5HE96ulR/MWzUMKcw
cCR3OwkrRAH/evqnjIijwxcVLDA5TzVuZeWpYyoV66Aq1Xr/AsXErbuBohC6Z6G6
r3Nspp/CFdRfbFBL7J9ggRGOOakAijICzv+Kk4Rg49MTW5J7Dr9s13HsgSfHCV1h
ZdNnz2DyK2V4BSpDNT4wk4nBVr/VIcWVMpGYEJls90AlrgdsgQQ1ZxtUjo3Dfr5S
9zfdO7OB5j1GhvUMOhWjIj1MFwbtGJh/ApNugOBnmQNZUJiOMfa6er8a693E0s0S
p3SLqKtStQDn6IMVafP/FjxVMVqLi5ankWfptLDM2HsnX3oqhuebys1U2GzfDyuq
t9poaUBae09VfEBTRB4ra3PJyXVWnJl8zPzH2iOChzrOBKd6ECjZrhovkFZ4anOx
XUdy40GvfNWvK/lx03NaMVme6sH2MY0nByArIGuf4DalnM+i8YD2EV3KxiWNfOMl
rTX/fbnaOwOQZO/4yJGMGzOG1l3oTLAyyazD+1MgZqckgEhPmqA4QAf6GdF6CdTs
Nl4SR2m3mgGUnCLM0twBmgh1VEoykEHAGgxKjJ/Hq220ZANfxSsoX+SUB9Iix+Lz
C/i3qij41SFbDzvVKZ8Or11tL88amTGn+JZt1UnxcFLRo6ky7Pg8Lla0w2CNvYq0
fN/DSwwwhEB/ZUQ2UnoeXqdEOhB4CPOK7Iwu59eQjCvM4+iEraf0vrA6+RFhjjkb
Rg3i1nUqTaifWLbh8UJ2aPwRX42uwyuJq09LulIi5V/Q+FTXX0hEjrjW0PhvPeor
Jl3aWrvafS9nYRXFZ0v14jWpodGjpin9nrH654J9Zt6VyCl1O5l8Lx7tkIcF18hr
9C8HePLIgExT8OFTYg+UH8ZURAeRlhrLAMckFmxIsXmwEJV8usr5yYD2J12/yRV/
VVjdR8cwmNZSVzzVJyo2+nn8hbBtmFdgvWub1hpuMWUVdGKN4A2gYQ+PhXZ9csZd
2iF/Lzow+wpbciiFac4Ke1pb7I3qnM3FBSrlBtNA+bHTXCnyck7gHZOEQ9Tq5mMm
ONBIudzKXjJ17T3dwHIyWMOD24LG4LK5PNFBfPJHr9a8cbyYRPe68vB2xjjUHSFs
PbXtGuMXOyhbpZTTSpu/bpzgM2n1iLJ8KrMUr/YUvkthVwB3TzsPrU4PRXXcs8bc
/nyn1CYV9T6YS4TOl5RSrWgmqzQxY1V+CPvhElLclMd27NAWoZN6iMao0E+jgyIq
nRcoupiyajxIBrmnwnCqBmD5SLHmtxIDiwOI66AnHI5ATRfDd1BLkdxFlw7Ah0ig
EHZa0oNZQ0NmZMt6bOayLEtZKECgUrqsbQgClW7WnwmG3ASCoT8szlg0dBJ66KhO
CMmA/v9wknv3Fr2TMP4ILQ6xUuYCtaQ7yUEAYpl6iVBY8Tg3jLxsNA7sOIC9zxKR
JhtmI3XtsR63Pslh93tHlDXx8QcWpJbfrtpY0T2JOQ41pT9aYEuLBWZ2ESD2pM7Q
dsN30GcDksMyn8+S56cbX070Q1RQvlos38kaOxY3MQ1Q8VanFTzNbuywHZCziBo5
LWEI0+WS2g/TOq9V8G17hXgqm9xVR8A5CtQtRSfUnhnxqz57scydo/5+jbx4QlzE
oPOmwgRjjMsaVzI6RMdeHNo6u6IKkOXNUVRuKr6tPZUfIpfcLCDpwxg6QofLLJwb
eHPkz4Hp/xdHqMSvnBZqGKz9HTfGRNKuM9xzYjSym9V+67GabcGsVw4e4RMYJo94
MvpHEoC58N+Ov2kHwl06cH1CYVI/Q9CgWRqv+rm181ZgNybdD9IayYiOf8a/5ALJ
9f4hAx0xn6/IXl5/BZ72TpA5gDW2ErXn0xH1lHSLWyJv6xS5SFYTaB47g+0fKkqp
mhssHzY+SLGwK0mqeeKP0rHsVDp1g/PQCobZADxIV6uJlC6DR8DhuPP/OlSVZI96
QkzmhNwKnm9qdayxJp1MMDkoT4WKjBhpmcLplTctIqRTnMgI7SukmqeLj5d/GVtv
1cLgR66lbnarPHb1vt8Of4hQYtC1ghUF+mEK4+Rzj8+Eb00FOCZkXjmo/IWKHsfF
75abWV/jK7ILh8OVvkcCO3W02A9drGmY8DwCSJm+F53aJpObCHgsdkLtdUfjH39b
MutFOkTJhd6KKtADzZhXt4/DrL+vN9lDkvDEb3q1U/FdQwCow+Sj/DFOkT3Ib3A9
jivFknhvpNoa0SxtFfAhU8E7xh7ISFYtaYBHSY3D6L2aIfrTn0AHJR5pg5kpLSaq
etXeUbAr1/qxw/06F07XsY5wG+ks2i5KK/HjuoBIZ2RwKaRxyoiJ1gcq97LUsHDT
YWDLd+c4hhEPuDuNh1YNrDijxc4f95F+yWXWTkFzpFOkjFm9h5in72aNoru5yMBf
6/uApAHekGC+h3LcGQLC8kZOUVgzFUBE0KTiAmFL5wFxsBVpHXQnxLZOiryTTO0/
oO0fokpCDIdDVNaRVm8iS9YuJqX1tvKK6ygJExG5V+DyW9BRIfleC1BlLkq7ld4d
F5rA5X6JIXBp+hXF1b7Rd6w38IUC7x3BXvMDk2FSerQ3lo9/wtplXTRepztEOxpj
lnwA0lljlnuOC+mjsd8m7g+WzThGlZqiwoj8blsO2ZytO/NiXHxDBfK6YwGAoJNT
6qKRlRx+CbIaAZpQldESdLpWBSttcrjEEx8MXz+6eJ5R4YiluLUSaGFzYnAw9ZYD
7VdZsvsY15OoBOItMQfjlRPri/6PacVChYJrQGtR5Xp36unhnNPG37jCw7b804km
VMK75Dg90tSqOo5ebWdVBOaYKtcD5KsoO8Xqy3JnaCdsrQDBG4G+T8X/qYGC7jk5
f9AlbnhmkIdITs+dKLe31mYQSd55HoHMLt3mMhdPvepCLav/tv/ijL2xdxxYUP+H
puEVayoIeqHk+FZdNuHb0qj3+Ed8LZ6ev2/DVjRL9gcpvkRw1ErgsgB5JE5X3OiH
TaRMWHrYehTAHmh7qtUN+Ng+v7SmtRzO2xrTdoqfxh5WMcC5zWiOftctXbglg6KL
G82mQfTr8xsJlxAsxA9sLakl4KegX6HwCgCyD9AKXj0lRrkqFezfKftW88uHcR3Z
4w+RAQCmWE/2tP+7xRQ997XfQsjbW2NnLmnwHva/xq5mOsaMDIKjjGL62e2OPFTp
6RzQ1Ss9CQD6p3yVnHX6RMS2mv2/fDfzAevSl7crELolRV1tXzGY1dO438HPnSZz
utp1ybbZyHnhGMw+aOtEjOwZ4D6/kfRfOgWdyhXATpeifPYcd6wk0MjjxKtHZOB1
QR7t0SRziapbnLGCBIsU4GB+oaBhOCXaAtiX/HmTRJ8jE2v+q2M3Ife7TcuMKXpJ
H8coRXkJ3u+5knQlJA7kgYwxPRc+aEPqkyfycaKuSE5as2G8W5lzNR8iCALJmwL3
Pu0iYe/XqspOPyc3tT12xGrjwUrtY3ge5RCVlBsHcSg+/zybbuIFkew+Yequ1Qib
QnAWRpgZaVdAHKXWbFVSZeqPOIYDc9OFbTXsIn9vnyqGpWkbc6KVydYA3gVlbeS1
qSf7TTo+OroUQ8txLcxe9vL4qeBpgrp80S/W/22DnWy4hlE6QEFk0h9173cm0VQ4
xPHJFskjYmcRexZwua6Au1vCD2fm05Wt+cGSMtgZ4erELT5cqiymZZSxSSKNwOPa
pg8+wWBmbqQBIz1zB6YJKx9HhJM/hKUU0BQlN4QpkG04nT9n0RX0rkZthRtkN4bA
GdkEoWBNU8VCBepF2zvCAfulalwknGicIfLd4wbEXolYkk4opxZcc7j4Lc9bkM7c
hzVHjQq0R05q3RC0Yh4Ng9N2fMVp4RY+ELtrtlwq0nHNmrIEOwAOTqAvSvRv06HI
5X4Y1qAayn3tH7AvOeWylewTdaftNZBKFrPb2LPVassULs2RxoOs1IUYTpwNvoVH
2faSZixDClyavIEXlUn2HPv7pSdnDiMAc6eGTPVfca1ZdUhXOTlaU8E1IINXhRKc
l15RDVbAruzSCGgHLoDpV70PGdgTUWmP9+ezwF4Jf831KGnGUahJzaXZTzWLFTus
DreRR31KJoEjfFkrPtsjR9hyaz8j+RJDw+HEgSUjNzoZQyiZjTIGln4apVMn3+uo
YN5NaJ1syQ8cI5Giuy2C9YS6QdPg7jBCLVFKjgYiUD8bSHlNdEOaE4/xwalEal8y
mzK4S9of/FZn069x4PxjhOVugyi8PrEXOg5QuBEqfbe0YiCf4ayUXGk2no9qqOVB
yh3OUBeKVht5wGYFrqsLbfkRCvDbEMOzd/ji0189qmXHEvbQ0ss1ubrIgX69QcT6
Zz4guOHPNWWRxTLuBVesFKJuOxXVmsE8sjb9Gc2vNK2e8upINIS38XZOARGGFhpW
efMGW2uwG43ERi80Yd5mUQd0Z+MmWoATtQLNQIQ5wpND0rkn0Olpbr3ro2aSCKyT
GcSd9Jjd2kYh54HLWBwFHXDRro+b6k0JE2Va4oh8UZTXaRFWw/dtgdpZ/ntY+HTr
Xe/TyJfYqi7/i9NejEyhbjAK2LkMDMpObPQGsmECJp7zQm6zZi/EZQmtW8bO/R4T
83BFizx8k5NiWfQCaB18yV4XOWBMaBl74Ifb2CV1E5Yb9A1VsE7+J26sYhK8OH/K
rUpH8vHg5gVuIxnP+rwDey4vR/lp6qEHXpJGq70hSXHbMoM55D46RD/Y+qUDYejE
uM0I8TI4hjI+/NIodT3cO5pnlNCb1YbHEcPXQC8NGbVvwJlzQfYHCjZsh5OWz3Rm
ImvuTswg52mwC91BRwKWhaDdLfQcBmj7Qu0SUVg1+gvGcO807jNF9V9vCPipdl6+
q+1lx1S7agWVHkuYhELCM0IX3aNcwawQ7LAys8aGFh0qisaJWv3qD7TklJrckIyG
Ig7QzDnGrKaHBZ8XgUBgXqbw70TK7IVbkII2FnH4d/vcGCM6/odqaJMYWr+G3Szx
LJgYgECj1eA43nPzX5FrVhnD+MxvzlZJlZ/NoAlXztSt+m3/o1P5uIk3duivA0I1
AkQrOOSqYjW66WYBn4FE9FIQHL5uKDg7pZ9l8hxEuLX1DYeCI+EgkP12AQeivUCr
FFvfB8QJrDrbZh6hsll7sRve281/Va7tYxwy0qRGL8FLbQDqMhT3SVT/LT/AryrO
lAGoYqDDXMxxp/CZ9qDH119UldSXpea2uG8AEUmF6JB6k7sh9ELs2MV1wYOwYBWg
3UmqpdH7V19LwpO+l1+UUiBSlpcVc2NVdCm1gAwFMuXQD/l+DrJKOmcwVcpndTjL
D8OWB3zlmqM2WWBn68TviYE91Vy/tDwWBcYXPDbQwmxjVG5sqyMAixjhWo9R1tqJ
LMJhEB2bz8xrTEH0kpZzKo54FtWNBANS/pq4nUR6McNwGrq+dYfnYGVcJEi9GESo
5bQiCyx8YJPdffsagDuRHTwYpdtkgjl5H/n8AjaTDXYOP3Uu4CoxTVlENSEUxE+l
WzxNEhOlzzjlxLfx4P2HaDzMqhIHS94pPAEqtbA4iad7W5ssnjYcD+pEU5ZCrf9w
zCwZnplKOXL6yBvS4M4iaVCvH4wOGN4I/H+BQ4nd7TT1/y3NkOSzTs0TMr2nxGAJ
iOy0JtCaHbfCSTymhtroszEuQ/qCd9Tz8Ag7QfYLs1VVv5etFtdusd91ivl/m444
ypapWUe79FGq6xD5jNODsChtujdJdQF2bxFsNQQbqF5XqKxlPmIrvsD5crJoIHyq
OwfEbnvOaIwhEeYhMid1eI0qxZWltK6Fj0PD8dLn9hZzvoaSFf9t8RSIbNpXmgqJ
cIoRmnzJB4ISmakfroN60JVOdqZl6FutDkVq3TB7NfnJiiVlQLnkrBTPtqBKE6Pj
pDfLeSXDNIG0r6ootjhD++WfzsgM+XDmFZkZl7E/7islDf4D6N0ADDVdD8KbDaQt
OUj423biXDZG9BI/Sle0XPuL05BBdThH9tFNb25lseqUTIW9q5wef8aDyTXh/3ot
Y4ClbbnEtzENheZQ8/jt6tpcG6Ovv87lV6dvj+sAtD7uCjAJBEqzQeEs6HpZR3rd
HG0T88vs+6mHup0nrNUN1/RuGbOBJucLz1gd4/51zmevYQJaFJ/uxwK4urB+FWAw
VCGFgLfznCs4EkAuDrwE20GlsL04QsfT7mnxG/lw9eTdkUjkOBR8sDfu68mtCVgK
GQ1DOD+tZ8Bjfx2SeQFccULRdh+gaobX++VpcAMtNMUzr5whyGI1fHtoocnGq9Vi
0L8jyO6AyTrxLNU7nF0kNRzV3OdoODy07eYMNRp3F7FFWfnqK3M8mW169YbIfA5r
eWR69Ps/AiHAd8nG3HwgGWOzD8MWPhmz2Zdb4RHhLzOSJPmNueSBm1k8vXaGqCX4
c2Je5UtaZ8HsAdyE9943bwui99Jk9RQBh305N/qrz3XFitqbRCRnnzsNes8dUbdY
8+HLf7URNIjuR1pdhmNzJ8yp6iYgRd+DJK2+hNq7PKq1abjft8axE1D7Ql/UmuS5
C8D65uwT0NwwNKacgwAGjIrxhJg2A25DAEtTxKkfoIeqLkbtE8H1JC/oEh8Kf28+
e0UcE4qQ/mhxSJAw9hgb+tnOaB5ERa+f0h88F9Ebo43LnYyLC9gWSKJacznifR5N
0TuzfPcgCAtxNRsfrFjlYqAM8srB06FxoWftKPa18+4aw8paZGWwdSEHCMB7Defq
/0lgyCzNZa28ZXbGnxCzmrafHRLR1czxvoju2RJIeg8IylGadGrK032h7zFrjJtp
eT8dn2V88JeJrCiP5157UK+XO1AGIoOBcT1R9fG5vZKWw8oJjVG7krhFG0Sz11N1
aew2WfD8rWYXBHi7nyagnUmBu5QGISq+ty26OQOLt9v7Q27LvXWNbNjgcR2l78Mr
qKimMSWOMSUL4RfudGyO8lxCRUkQpWJ1Fzu0qxRT9hpQndU4dx+Dpy3KAvZtVthX
LCiG5K2S4ToHsTwllpKJxZG/N3as98VGU/0s+Bl7ovm95IDilnr7pqgNadcFpzDE
3VoWVzbhHPe+VDcIiGqdOjSJcJFUlaZqillBDh6uAjIj+5yfP2dgrJ9O7bIqYicP
ZSe+aVSHlX5vv1WFf3q+n3uVgmTRaFtGK99jE3YEejTmClbm8SEIXsiSa6NnFpKu
/Cfe6zH1dW9oW/eI/BtvNUyzq6ERDmjveYPUCFBUEU0wFADpBMiuCCCqEr8TBowb
hbV+dBFxIPZCqG/H5JfaC+ZrVg9KUoGcbKchvIIp2S0fA/++afkFNO2d0jC5nQQS
CIGvuDYwmvt3uGjhX8yWIOPFtNgX4BHwx2oUsASmEgHx9rYutAekJVYxk3Sb0Ckp
5orp3NyFKId9rlwY7ZDsqRBFZe93htbWB/Ys5zeze5AQkURunb9OVSaGgj800uyL
hiqO36JeiAgcpWLrZIozlnWSXmsI/y09sVXaqbj0GCZpm8VV1QIsk/XXtpbkR3iZ
HyJ++c4//hq5WDJ0ZN9uG+JmOvdfJH/n359Js6A9FU2C1qeLoiuXKZNlPlUS+kY0
vwScE4coFRFGGsIo7ZqDHYTk4DSwwt7s4HHLb8plxuQa5l61tIQ3u8amLCJFICro
nmnwlQEaufHA+cQQFYfCWX2l5pLhVJhYXoSrW+Iv35kuMObHUYSoIwn7cy6H+Inu
uAewpTFOP4jT4kocmnuQFmzCeBgip/4j4k3yTROP4LOmkZzHcWIXKeEnU22KAEN6
5LdO7kloq2B6SARGMF7u+eXfRaVUeS6qke78Is0aBFBu70WecQe/GA4DAz52Idez
O3Xni/Q+HI10g2m3l/y76kZOUatDZs7Cubz2pTcaOoSomY0BNfDLFJ1IKgTySuTh
RpyMvrie5PODzHxs23/CgMwt31K0LNuuEvLLmzaDOQce2DdTRyHV1ynaWyeOG+vS
geCeyPHjRm5fXSpnpD9YjGl2gl1QzpftzfsqTpgQXPnuIf7e6y2WzzKmRQ9cyqcJ
WpfR3gMzcBY0pIQRj+ABOrxpWAT4CIn38o7p1g2CQfJjd6vs5cNk04VPjkLajja0
wVmjL2MFbeXYXHB4DzYLnFmVJHp4EmEedAi6TM9QeT1iYtTRJb4tXBNvjtI95y4s
npXgHAARVBbY/Tj4e5qjA3JzslLoRl7IA1zHvno1vvbthEmRD0pnk86fxqJ4AuMC
qMer/sFiyN8m9kBr2tzP40LaMJOFPKGDXNPLsSdBiSEv+udtuE9lyxpcUo5wef5e
DDGbZuZRGUIrZA3yBfkrF+K7ZWO6fjF6t9ouLGMrGP76MTpdqQVN8Us0pGMqCiuf
R9LWlgYoQhSlL2MhiBW7L3kGIiNQci3wxaAuZj2oe+L7p1qTlLQlpO6LXL+A4WG4
goa/VKWrS4Jar7KzRU73theUS6E5mUdA6ZfQSruCedJ5rxS5JTPCKrGhivgxklyR
v2gyhw5JFgdJIks5PE0zD5/FQWziwl/bCLSgaf1cn5pgY1eX3ng1IO2zI7j+Ze8M
iyEc8WvGP/rfRoy2E13oIBsf/W8H3Z1vsI7SmXEjjSWC37JEp8nke1kRwTb7Q4W9
Q9a33VzbCwNYw7LPgmeA4QFGkTA1gffVKZtZZYuJPufFXfHIWoUebjs6HvsoEqr8
SAF+0UdR/gt2pcC7EaNKaUeQJTAS1QftDVee/KEKkNhep4PFCXFKFYdIqOI0Jraf
if83+Lx+3D0vazLXLZ1BYKFwIBKFTEryDebRckWGHhNxFKsH29azNjal4t7RiAHE
vYpM92VbSmmEpUypU8YYAHCJC2j6Na48cXQcq4P2iusH+2uB2TA1RIhcRvVPF/ge
hGueW/bJgir9RbPaqHe21cSgKnV4F/sDtKABTTzon8rT/pIwKMq5ThS0kMxV7RSB
IiWhCEdRMtha29We/ZYDsdgbc9HuA3HrPnWuWZhZGHLKKzhizFi4sMyriuyRQlHf
+eBwsRpaNTXxgauqGRSjzF09687MMYJOLocPshJW743oS5iIHfo9V51DmvpREMs2
y2vePZ8HMA0n+2xvNU0e4g0E/SczuhsZ6EyJJJ5/ZK/VKBTu1EfILeiVwH1AczGA
59hqJD6bMBcQ6Zt6jS5F/yLNrWY0Eu4cfQebnn7vxklmneOR6RoJ+SfV2tu9FIT7
hG1bKgFQ4kS3ih2KF5v8fVXS8fXIXZ31Htx061XNU6vc5lKaD+gvRW1PrJKJC4Pv
WOjqpr83FroYqBmFTFQSBESEAHaqrYGufwwQb4dvadzbOkyCMb90X96qgL34dtfX
v9jnXc+9xwKB7tnTAscDZUXAbGCj3caCwFNTkBismV9L9e7U1n60hWbcoyPBNsLV
nFo0QjwbZgQdBci9glrjd/BHvHwcMwzfG+PVhW/NS4lmEQkNDlxZEeAOFuslOq6D
u0pmDi87+da+fpcT1nYFFxzK8VbDvvgnatGUGvKXCmnpjD90hLX5wjRZKSL0dgZy
MHy3WD8NV5BYu/KhdOFE+W6pojra9iV6uSLBv+HXbGmnyd6Rly0RReY5Csm1Y3vw
XJlHPleqKeAuSWObTO87SCDAu/+eUjORmJcHJM6ylU5KF8Mjzrrsf3WpbkDupDjS
ddRFoyI2rKKOPJFDrhm1BnmRS8mBMsuLF1HSDaBKjupe8a9SrT95sci8Fz1mUZPq
OyD1kJ+3lsJJ1Rfkeorx04wmLoNZdn6Oy+Fu1CFlut7bIpq8mQ5+1BIIIQ821K/e
9qsZtmsgaxgqFkKlF8CZ2L+kbyJ3uGzDO1ZQgIUqaIBmZh7dAaugXTEMVfGNF16+
VTcvqg2rz0szKrFvd8yYXz13dL0RgLpNr1ypWdQmIeaAG0KCp7aGp3FKdq8qgpMl
HNEruMDzkNr1wEOhQy6JNcg9Xq8daCDctHRWo9xNcZ7N5CXBOrZ70t9iZt3b93z3
afVoIomOPSyru0gsvUuXEDpWwwYHPBPJK8dA2SDHxy3nST/+/yqFEsa0l2CppUmR
S3ERwtO92Foie+iresrLpOR/qVMXCTyU8WgreKkReE1iCPoKFWrvjSC21gu3OM8L
I6JvhMB+TKzNHA6pCGQbm2ZjDGHvTB+4148LnXmhM8XJkRo+8uNTeVx6/Sec4cv8
c914cBAwW3bjcPmtSLhve3sVkTQF31RKiVU6YZBHXcdlYDJGnfbMGlAPbiBLfPSx
4wIaOmSP/3/Ty4ghsrUTVUYnfKEGZ6qxbi6lIabq33ZJVg+0cuRuosy18IAoo6EF
lW1Q5Mrfu4zBQP39I1/5VlQxbZlg49R6GvWSrSiMFyfWa4nznZdQVHez6J5c2duK
Q0A4QghKZgaV+xeTDcga2UgB1DwDc+GWuiKkrdHoAa8EGQx6YFx7VUVKOGW3Mzjc
I7J8gueejjuHXFTPB+97uSC3YFSFuiz1BqHibtZa5Y3wmXJluI1NHpjbRM9TZKL3
ghjQXjr0wwA/YRSzs7UMQBJaErA2B/TYRTobSWFGUoZtEPWQwilTXSbj7hlwShN+
2NCLtY3ZKjOHZv6X9EiYomy/OBDJJTakpkKKCCNB4lUUHB59N3BtHFg1oYC+LS5r
Txp530tTml1BcXJvmt9c6kaIa4SZsylZJLbrf7s4jVLXHZp4oM0HNsFkumCNsjf8
iyzcaAcwu6MgCX5gPUn0bm3LjQ/XBkF3tlXRYhuhq2q5nEWGpYPuJAl9liseQh0c
17tYiyDNCsFo5B+zL97avzLel+S7ScF8I2YGEFnRCz5S2dfOyFws/2kKFkQYUCg9
k3JiDuRHZQ4J8sOKkZfOCWcj0dcZaeT5tF5T3krm4C9lcdls6TczFtx+kJa9rpcX
UjFwMbq2Byod2xZd7+bQBpIBOTy4IeXkr5tOUZLP+PxnSjJFy/ec1g14b5R5pmXk
vZhivom6h9zmf46gYmWyV8G2oECRRDilis+cB321AlwYv7qRFFoXrC2vI6TRy9Kz
iqBNrTkaoiRyrXkHBmbV5ymUN1Ny/penlnrREuBRvGDPja9CciBvVu2nzIwPVwxi
2nlH0CQyM0ScAuauDdoS7QUFdezWKYO4GrpfFcKr+0D6PFBOHwto5JIGQfvaz6TB
UvgV5sIfWpB09Z0+GnjsN1EfAgiymnmM1cOj/qLxJhALwANCM9vi5wR2vXPSQ+dg
f+fMYkKMevY+N03fhzVI/aHCA5FRrP8l5Vr2d/Jr/MCJux5WeJj4PEJ50CGu08r1
K0pcHoXLpnlnY4EmVWnhJZPtiYlnGfBuqoZ621G5ozCKozQRM6DZ/wdUFkyfb1Wx
ZvS52QmfLRFPD0WWeXGFXd80uFn+CGgtFiZo85iYnuQpAVuMeIe0A2yGsySxAv7D
c/fqtJvUjOaN3tO+iGb66Vnl/Ghb/8aENauPiiIQKqZilcDMaTFMF+M36vEao1o2
OnXDnBb1hObmzIuctP214VIdsDUubngbckIYmqck6EL88JJ8g5AZ3OMLBDJBzo1g
OgwTUR3YVqzyzVP8Ny5Rq8iSigGHUGswT6dfMkVhY+Hr1FV/RQxJHurtVuAM2AYz
wuYH2faiZXhZ5elbnMoKB1Wl7iw+M9XvEyoVr0tfDZzC4QBAAB6CxTGlNUBwTQzf
jyUa6D1Tp4k+ifgxhwpc9KOdP+TT+3kVVEUGXSTCJgqDajLFauNzSsFWucRCXhTI
7DdJg/In/4jrMfLsKzeoyyEp+Wy/XfQEHJc3gcu5DeKGrKKjWpzZNB3WCtaN7Jyk
p15zgGPhJ09SVsL0FbuzZNaR5tMgluQSSX85qBDYFz34ncMSAj+DoKZY4ZmW3o6n
wBgbpIZrU6eVHxsUfHpysV2aVjjgBFfX4/xfSDnFuX/RIdcEZRricFIxU/vSZX3H
jw1A0lopQa5MaoA1hgxhGQ2tbO6yruaBc2KkJl1qKo4rWcI3Lx9lreSsZWjMkhPo
F0F3pic8ysDtpXdrDbYCqScJZ4b1k2ZILKDgf3QZf1yEwXh4mQNUBqzapr17ulj3
JHDQge0Rfq5HphQWkjMj1k25FGtaly5v20Ke+0iv7MHrgKoP3cLbN1bhSl7QuTZH
nSohdG0uVnHQEf5EtpKqYautRBw2mJvwk0867nK6ZZlOXEAmHWHg5mxIl+CdO6ZS
jZXkEC0K+jQEMEbAOSrNnrHzW+z38HxZ4AloATH6myIYF6SYk3Ntr7lXRzp8udIS
6YOiOeAZv/5WeZzK9SDmjd3m/CcMuywYR3qefIie/Q2/ByqvFopFTF3KPf7XK4bN
PMfaEAfEOLMjRKe1dKeb8mMOjmMa2aUU7wdZwsIPNbb7yQxemMRNcmLk1tuEAKSE
V8bPcAiS+YGCfQ++MG2UYZeTTHjWWLTMIA9utAlkKYRRr1/CmzjfSd7aYlju0nzj
CTgtDPgLWjUvvVqRqSqUTX1VMuzMZZQrw2i9ksNl+MvzpL3JjKa7KeBIAZSSC2u0
iwNjUvMqAnM/3g0gCOSSn7/+waxBsGnZpcPaLRHL1YWQFC2uEHOjV7xSZ0BY1Pki
6/WuzjB8i5QbUxxvYRiHV9wrX/fu5BcoEZEC45wqZznnRtNwhTdsR6KZ1wv4fv4+
pmxPccw68t2v1bZ6nEqjhyvtDOUJo4q/gXOqXhkSE02iZT/Bzn7c8HkVgI1kVJZx
BjhDslF72YBGDCe637IsXQaB3/bz6kzbGpjjjdFPAC25QR7AgILcjWkGN8k2EDEh
Iv3XzSrBTZe6m6FymRmiNPrqoKAPBsjpjTnv72+Nyd8I/TyYKm5x4Bzc4VWVBJKM
HMbn27aEgOE0s+FEV/COY9/0wGf4ZM1zubzM+R9PIAEYTBxDHyP8qOvfAHup7tQq
80jU67doy3hg+76vw3eVaVsBmF4+9ojokvWU8ieZlGT3r7P8RVsoJOK9s51hCDKz
YdRdaiqHIvVTnY5UZBYP0lMCuV2ayU1tKBTa3MCeoT+qRtJvWFhZybXGGn+NzLya
qz/sb3qz0PPtDNX7mNZZYgXq2kNbGh5snLKnPr7yVfhGJJg2j3wWlWdzgMrhEPVk
s5cmbwHEP/D9DJAv5m8rTE28RycfaIV5i59aX06Ujy5JTzCQU9mELP8R7g2PuP0+
hM7YsgGDVdsFhHC+qrBbyaTVV6zdRdOFvi4FKow/UX1NJCs4p6DuCvSBlrXquD/f
QThqfagmJ2I453ZBFJyI3ee/HCuaZX715xD3dUatefMM+11N5Ampyb13E3kO3ahA
h7WNUmD8UTqcjoedqkp4J6fD5PtWuqv7LB1w/0GcyEKDj2uUGEMtSCY1azcMdPsG
bpwjWkeE0fAS2ijwPy38QdehG5VATEwjjLEdl4f7KeXO3RpacdcKRqhCZreJjVtS
ybQdG6b2m1H+VjZCn79v5GLHkIT3251Kuk7hFolE6F0Bk6Xk8zYc9BVO4UPMMSt4
6V1AIvTJRLxKo+dKr6t2qUi27AwI3c2xUl3gNMqGCp9Dv2jaX3VIg5Mi7Ar+FXKo
84+CJ0zWH5KOs8KefnFYb8K/OWTLvhmtrKL4tm27mYP8mTPHTg17IYGHlJ+0k8vs
2fbpc6zKAROFO6eKG+tbszY95sk1rPASLuf8MTrcKTJQa6I4fsRDJ80U7NdBMGyr
8hj+Z5f4qR/pBU3hHtS2ML3KafJHnLkE/EgCUGmyHaAQMFX/zZifegxNkGn215bI
wwWVM8RLVxGbFQamkpbK9yarbUd1Mf7mJEtv3/p5w5P/rXJbxq6R14wiQNW0s1Uc
2QXqdtyCV/njGzmcD+KBR7EIfDWmRe4T/4ckOi+ZHsIH1mk2iUChOdQSHOIHLU7N
v8dLWbrTl7Z9LRTcMRcmQSDyBSDHjbyT5XAzBEYV/bcVK8uJaF5VCB7N/wZkE/nd
zV8Eoq1sTYiZIUG056n/ONDPoiUfGL5LQdiVhv4doMFJ4eiyCZ93I7IAeb6cPccJ
3d+111WuCmKnM9ZY/RO6AeuT3KEglSLvDIb3+pG2hFcKXQc2OIbbh8e5F8NRkJHF
TtgkpKl355KTPUxquQzAjfHma8EFq1dkmSYff8smiViVGnIGxtn3xozhPApcJ6vi
qxc7CvOXr2VeIGIYRoR1cMeOwJZqhYhKxuv1gHyzWGnllzvWJ8zRmLnSvZO3HHO1
D+sFV8c5QyXW5JQdY4oWvU/a9g6NTagWMK0pT7MB0qKN/23jS97g6CkhN7x6zsLv
QFfoKZ4LD+wQfpcIDPInmiK4xnp5f7/nlVH31e9he4NwIFk6dkQSoUj834fpFQ2h
sKNGAul18FmLtD4uXPzCrMXs1oTYogk2lKq+P+NQT2n1DYjKsEswEByVeQAh+51e
yVMitnNbbHvTELR0cB4JCCBWxonhomfj4sg5Gke0GY7V7nI9qf7WfHsK6V42JJWw
1T7vDerH1diccdkIAdoAFB/KvA01aCy/iC5XPIKUUN+8bzhQTdXrSSWZzGFKG1/F
RF13W/yZWGkupd+Stcf4vN9pgHPNgRnGl27mJcUwGtl9ANSKbTjgE6Y4ssVoS5s3
NQdOMGN3DJdzwGr+ps6tWpCpox96vr2ECTa2VDTzB2S+kXqWhu7qjDppMLyM8M54
OeYbFC1oEIB9F7mo49lT2quONvw+xaB3B/r0TvOAgmXBvjn/0phWnrkz/rgy6aGX
8oElFlFABQUYp8HSWMLfa+PSmd2EMz/2TsXdu6ytmH1x3R7PrAsRo7N2e7wi+bCf
JZHka41Cx69VXGLcbnxKv65ephXd6uRb+e8wRgXmsqJcrxMCR7NBL3OAgX8Ime42
GyttSAygxEC45zL1pUjbDrFW7UpELdTuzUE3L/f8P8QGs+TAOBADvp3E2xWpdBUu
OvGAACZA+IhM0mUk5CIhz+pe2sH4/h4eBWy3oMCjDi1a3WuoIm7XNe6E2+Fql8X/
piCR7r6deJa07FtrFCwu2uaoi64A14jdA8YAjLLcU6OCVtL0rFXHutRRQreckj/e
ZeexpX4qw3mAXHZS6j4bls7fx9ouNZLCxrXrcjSoVvzuR8GQZC4Ag/eXJjMvRsfl
Y/E8uzbnA1VWG/XgKd6quxWo7/Z7ULRFt9xHvUdQ9rvWjPeXeBI09VHLYLiYe8U3
XQWRAOKhMSgMazTHIrMdZQQCOXGgSL0ufi/o7O43xq1XjjKsKNy8w7jwaBXTyCcb
XYb8a3ACdW4F8j9c4/sOw9O8511k4MsH7QFeZEyNPJHfasX85FHMCdUT0zmupvlo
+yy9PwNo6YsRjgaBqRrTV1M5zrGPasb1GjlrROcH9inx9eUdFjLMB3ukJyvrkTMC
nqvtG2cfRYil/qF8+rXQ6MyTyDXSPu/aQ0rgGC2t3U3fH+YEYnjKHv6KntClfdcw
HNl2WeXMctJCaBtyG+Y72+CDhnmN6C1tgryoknjkAqYHC3EuXE/5J8HGswKCuL68
jRtjCodTZ6Qer+ZbTk4kAB7Lud0AAvu3GUJOlNl8EKUVSXeYnoJj2p3OMtPnhLDX
VwfhX6hhBFDUVZbVsmOxgzGC3oUhi7t0d00j4ReQX/ysyfx/NDkcL/jRhAYobQev
aa73Ti293OVJ76xQtvhAHFtQdBc1LqVdJ8uciJUMkMGtZ5F14x5a2lqaL9TXDEXl
bGUy8JpWLyeWD+Gqcee8CsATzwaCr57Aou8qaWErE63/Ul3eQ6wRyiu+hceAz0yD
AszQPWDhF0pAgdHAKEJPneLK2yO9y4agQw/xQLJoQUAS7aKunho3pFmv5X5WlP6D
TEMm7F/ba6dHq4IxZdRmqZ4paMaRbZL/O6sXYoKdkHAfYC44q8bhn1nFoF4Jumvd
iuV8yM3qJ6x2x//syNMUjpIfp2G1KG528Xe4XhDfhhkv+zbK9SJnPpk6Q9U77kD4
Ua80cSc6nB7+CwP6pcmqehlG4J5LBS5+u65FN1YvzG5coUPQidBqZL9hwRh0rM2K
hcarWb5aWDNQxvn1BJCKYOScFKzRAz1Vvtqqw+PYkcXSkmr5uSK2eoUme5920KSZ
vwSBs0viK8R+McLtCOrNIiNAEtfaNDJ7H2rPRKIaWD/PZi4IACDkrtL5X9+gE5Ll
GlGsOek1THr5SHPbXafq7IOwEsroc+SILmmAz0tX941IisCnrmL4fFL42XLzhm2+
8HEZ/AI2wtTP6pS3JFjF7Q/B+uxK+GzmNEI3ddJIL93bqGD0zNE5WietRwakOPFJ
v1WFQPl8V0HZLz58RV3IGuP0x8DyLwYDTiHYWiVI+YzB52cU79qqoNLNG6kXDQAk
K7Ho/+MBmuCXHNclBOImRthvTY8A6tLD4KvKKCMbzJ35YNg/7wkYBoFrFjTDIRN+
ZyzLwJi3iRHqQ2Weel6MC3SXZdc4ABrl06hle74WTqDndlNNp26NIpuAcEBJYXDp
o9CDrcVjyXFyUbiFrJUaZqWvCSoShqPVB751Fck4qSkAhxaaatIRHS94ijEfmN3z
vdO0brhIRVZyFrtgIY+pXQf74KXQbSJMEJnLma58tcBp7tKI1Igcpc5/Vt+0JAmQ
4604onCW1bVNiJDBt+oJ1tFCpQHwpsc/gI2aXFvIx56vytJCkRjsauLM1MLSzeNV
lpQCjUvViH4Rh/kvMHoXquWMLMUMx8ebwKn/ARE/YdVICH1kIojB3QRKXmGSHLAg
HdfwFwuOv/rNe6KOK4NYQdOTcmb0EBoGu8m2NJA9RYBfs/BaAFTWCJ6qCD4aHqgL
ncKlLb+c9Xfr2i7G8H239S3La4W3sRO8DR+xWLLihVbZ5O98n+aFHirAPrpdlGRT
e11qmQl561Gpb6Hg29DhXEJt5NCrJE5v6mgnHZjIJoyWGmI6Uf+oZepXZilKdeZW
C94gmDz3jz5DndSe60AtYAsi2+aqg90dBLw6Fi//xkRXTonW54Ue2ISPgW9kjmfW
jSD921nW8q4IR2pe0zUGKC31alVGONz88LxRaR4sCYvG8/qV1it2M+2fcEE/my/G
4hDnKkrUL5M9vwOAh9/ZYwv23FgaE2ko5FUmEz9vDeEC8HCQtQd4y4Sxkn3VdgvG
m75hTrdVP2qO7IlvBEShg8TaZZxiGoZWvvnNqpWnOleyDMza5ulUYhfxLZWbM+xc
JUCIiPQYK6B8dOprGfqpoQqnrsvB2ov1d8YZlPgB18Y6Ne39Usqsst8nWi/KsyEv
sTfJp9oX1iceDSTgvzQ1NqEDZVRKSVRGhGRUMi36GuVSFiwgv+JTGVbOB02FDm6Q
wDk1uwofYoWKwP8io4tY5LH+ZEiU1E3ehxiKjN0MJpzzgWtHL6bYSjwigxdK5D1K
SKRjD9vSXNIzc87HTXeINuV6pEw5timLG7tE2SniBOXcyLCy9DcZPSWG6/g1p2V3
8Bm/b327LNpmrhLd48pX2eypn0IdGozhfLnEZckKwvlOV7dYr3WhAPqLfquA/Tzf
aSj4OvMUF8CjA5zu4Wx4VcBbBUK3roa5oQ1QfoJNotX4pD+1oyb4m49NR15sqGAT
J8ybz8VrBc3c90mUy66Sh/CujZYTB1blDA0csn/QxER+25UVWWlJo3mJQBkM4Xkb
0ytIgY0AFjpz3rKitQ+/TwzhWdI6IAeQ34FCJVOFmxRq3b564e0i0tYgcRb5hz+L
sl2Qhh1GwfhdvpPfIu4Ivh3aVQxegZe3f90lvf56grTs3cpPWjPFJjAFO4CvT/uF
Go2r6PgLryHbKDhdAXZzq4yH2z6tr0xm5Q2+skd6fvYDzp6EKjBPLDqVag8ezMUC
vpv3v+5qUX11ebWiAWwsC/zOhYpKFnP3SMSXglz9LY8Vvy5Ls+FO4TxcnW1wS89Y
ZVLFya1ZgVVnxSq6zB2Paf9eU/reLcaU0MckvR+xZZWRKrNYyFBMnzvnXlMr2QqA
1IuqNZ34BymlavG+1IST7r1x1+CD6qF8hlM/TcLDwqLhULuRJ5GMeiyCqvhfYzyS
IHpxTUcy5CjJ0HwwmWL0xuNhvgIvgSuZpjEkA0Fray0e014OR5/zqVfl0A8cGQyo
O0Tzh63nHps7f2/mxq0EpeCIC1GbFxDmmaoDdSg/EKGEl2jvb+7R36RnvGY03pgN
ZFVf41qLoSJeyIaEXhjBb/AHK1Drsd3o/hkOtVurEDIwkJLE2YL3ZQryhT5xZl2C
iiqfhYuBKwy9yB8ZijfiB5dvvJ6wS6+bRlmGgzFbi27A0edUXJDlZAvlBgdj+Gbi
kEnENhqQvTDiJHKWHlwOAPnIFI0fozE/56SmmGtyGNdGLBJMAgr2kVPKaPYlfcRM
ReAt642QsKbXOIWzR127OYSi06LPUQ1MiFKLvFh1VSkBg5aNoE6e/xUJfEGYWh9I
AXSs5mg/ad1Hf0QgFE5tWV0WuPKbIZpuxLf4mF3XFtoTteKRZ06LU9ydeSFvj5zM
JoRcaGp4EGSXYubARP0pPbYqFr61bRwEY4YQl6kbIeRuBDKZr62inEaaW8mjDmT0
aX8BXMCAa4RNruKr+3gqfdKe0S1AZnBJcqecu1iw3nC7Dzvi3qurl2CTKYn7PfJA
sHsxUXXU+bl7RvmH+oK5bJOUxJF7rJSbUqWUgirgDPl7lHKJYFHWIxU1ugqNlmWt
WGPQ20sg3MS6ZDsxEsE3i367rcWSn6u3AJ9JCQsBvDIcECGHkmyHwuHTYuf+00xl
gQ6OVVjdPL8MOFb1jpdUcD/Z30rYHxQqXnNIarLrdjvYJkEecSerR7Lt5vcXB3iq
lfRYIqaxS6RnfOYSDUX3L94kXvXxnYwhP9mElFGIDvkSZwfKBr9JB/hrgQDnC9EO
bxwzvntDu9GDDJefwvLgmkSakPenLsk2T/Ef6ai9QvHzzcTxxZ+SHmgjwmaNTCxc
RNMiAfejR8cpHV8GHOAqH50urfHbSSzWm0zAn+1aVu5KbY2gTvFPsxlYXxzeyP40
LxaG9XdBt7OmMpTeM/wTgRh/fsapo2dPI4/OaUiPyekORjAUjIy8+dAVJJk0ZlVb
FshKeCXrXWGk4uw/K9AdUM5XIGls+508z6GAx3j8LPcX78AigP3fW92V3DD12gI5
wRYyULs725XHIIb/yopWHhZFHqn2H7+TjTclU2G5iPWNJ7vHVyB9GAIDLC8CEjlQ
T5ejuTRrJeAZW/HW1KCymEunHvxTYMeuTyKcr4ntnffLz6EKBdOpCMyNbMJr+Wy8
Ytzx02HSR0QTfgzEGicuVpFbyu5KJdGCyMsvcM1pVBENL8EvbOlmpha+SOLQmMeI
tKIxvlS/fbpwQ0j+0lbTQeWorb0HK7d18L4eTnrF+3UZrhyRP7D7I3A3vA8MVRmu
m3/eN3OUcYQOj0bgUB4E5oH9PX/Ex7vptc7ys4ktKQDQdIwkjLZRQf8hMQsjNG3L
esmeh7Fz/rPDBzM5AsVLefDvp13WBizTd5POCPwhEFy5Irtk9L5kXzjQc6oB/4Eb
dv0/pVvV4+E2+EXbb5OWxJ7loUGfhqhnD1nECyfA2u5AP7cFA5DrLRS95MbpLucc
lodR4DHmekg2Pg4wTgTBcSABiFLGO4A1GmZHH4bEWoRPL1nAun1nxG7352vQQnHF
ctWXGPlAhUNAIk/is0Cq1d/OqYBikRZkGGOqM/olTbD8sH42ZYtH7YXOb+xgG7QD
8ymnVG2/VGBNAfMOSO31eqMBoU9DIptUpHcVnP1gsNC4eaRHhq+tsBgalLH3KbTp
Tp7s7Q5NP4IjsBnbiYjQdF5Ijx40jstjvYR2r6zn/y0NovhaCkiiuEulTO/yTEYc
WHxFBrygPwnxrPzYR5Qpd+GPq5ExXd4QGx+V4ejjk7RZD9rJ/M4aL/jmUryV8gTg
axhViSoVko0SFZ/J7Gjzm+H1RQ74g9u5XMwB7csvp5qzZbDoVkhYqxNPuQDnI2Zx
t9gl3QXLt3D5ZUp9qv42N/chQj+W2vvd6USzZSZHgUmJ7oTJBDGECh1yP0qq8DnS
+QcKgHejrqZpk0BV4C7uc7n0FKs+1TJQCHAaXC2E1aWMI3Zq1Mz0ixWu+6WkXRSq
jvb6jQlhQtT2VjGMaA4CrmE/Y+OWAh8JLbonWNktpAoN5Tjsi3VRfru90j5l7xPJ
JS3bKl7RSPeOR7+hCAp62uYzwkTqkSbLVLOJ9Vn+PbK9HQ+efpSbBzae7Rz0E5Z3
pWZ/8JMhBIf7aMs7Iqp8pMvv5KbktCuE5WOJKYe/sRYLSOtccZ5zpC3RrPR8P5b/
BN/9DyoTZ0uwulCkTEbWMUy1DvKrttluTYn8Y8vj85p596SgfZVsHXOubEXr6TYo
kTlMztrNYpOY+V1TlrnMeN+DfZVfs4eq7LFlDPCJ7oOkoIUZRM/90JEJCizKY4qd
0ztjhcFNLLTcy3+0+mbn++lDqs7BZUkBtZoPqho0XgsBaQxfCdaQRPQHjgeAwmMu
0qK7qAmtYO1eB3vpYo/OWau3iGVq4dhlsYDTZbPS7sxZiW/B+33h+xp007TtcBpv
M9udWgB/ysamhpvUTyCcEI+qGe+yIvItGakDhaEIE/bwz1q2rBOurb8KC9Qt7cqV
N6bOAnQOiJCrT4qmgsFZ9HhJzqP/lc7kG1r8T8Rzs/Bc08Zx1qAbCKluE/Lm162j
a2+rnwnnkKLg2csfYrXXDUYBdgjfb3vzhHwwmb1yzup7L6lEe1TFIdQDLfnu17p7
VDB4BMs3L4AnF9j6p1PlUclwwMOPH2SCn9XyACoD+5ZAEDPhNPXQYRuoIVON5Znl
wU34MCBELP6rYb6nVkivzn8C67o3epbuGkjZYhFeLWKrGaq4aUi+PAbvehwRpV8q
9wkWNncnZXWpi7mw1efzUff3LxvX4k8M+B2CuQ2AI22LuAn4Lk/2NSt0gybRYAkk
FfVUScsU8sDBPVL8qNO3zERHQyF5vIB5wdnWQzCM1LWSJmTM7Qpn1UxIaHsrdrCK
RWpGjqL/pkeGuMovC7gEK8Ait0qDC9F4CBP8eqk6iNM50qI9gS9fCI9JmwLQ61jv
mis46mNlf0igV/avk/9qGJgegBSMpGGPmHsN3ldvDSK+C/gTki3IKLcymZ2eFY0l
ZMWSYpqELepP5TSKqhVYWcq4+ZirpA4YqXxPSSxNuf4sXha6F0/Ab5dkpDNum/D3
CmTB3LWARfTcNb0iGSlVFRBRAQlu0wBgsYlcUpzR6j6WBUUQGD3t6Ir0eut6Cn39
nNXfyW4alDM7mAGb7iQrWhlwXraPu2P15Oi0AeMFdAhjyfES0RcNq769u+gKBeG4
+6uE0eHfWYCvvkIkZHtSAQFL9Qgzci38JFg6u2AM0PR6VALEIO9j4p/6f1kCSOkH
xnlUA6Pj9JJ1oB9pskkyElabn0/f6evKNJqdY/vY9vUpLujhgWnKcFqehPy8Ht6H
Ew8zTiT+MeugWbFP35YdHOOXDDf6M5N7XnYy6i6f7Jg76wqhjwhRGXvQUIpfol3z
t+iOnY6g13F2OdzQitWJxBIKYNx4fMEtE8SeDCved9BHBVjy3nu5efKbTZJADqEk
Ot1sIlH074niU/pyGRlgKBGJ1PsXy0qrDo4TfEynUF8CIk2ySQVwfba8M5dG0Fwg
25G64N+3x1oBq9TC6f5lSSkQTKfBLrbP1ioLf2jj2Ms5KzmOfwUjpta3C9rKXKtw
/rD+9Mg9DJHouQODwoFaV1d2//x7Ub7CNyoQ8cDw9/vavcQPsgx9fBkdwSgCN868
KbQQmN/iGyv5GvYz/v29o542X3CSR9a34oET6MGMrNC/3RBm+m2S/1DPdZJk5Yt2
AT7g36Kkv7nz4ezoKHHFMcajJGzSKwox/AMqwYaJB+MUro62pqChjFJybdk/eK/g
SReqmxgBPlYPttT4KdHszxtoSGt8xFpeUg9bcvvAEYgKJlOUgArNWc2H1yZprQsi
fxib6MxWZ4W+MP8cSPnFW94S272KFuX8tOUnDHvsZV3lJNYeb0d34UDyUMRD1arp
N7fEyhZiFygLBtUOgqPOMBTLAKlAOUzV8TxIhX2bojQUQ7ID0wjj5TALjn7gVOKh
7+2YZBFBx/fai1hSdCXg587B9hNi7mLKWDsmUPSsh6RS9Kvz9Kn4j2/YquaDnAaO
NSEG/unqfCakFQ+A50/9Bomd7rZvbJXxeY6y3QH3uvc1mEikRDVB8wEuvZdPED7Y
gueRS4ujT93y1PJd6fGLOUJdy5Zm2Z+4Vi/KmhtpZySqwNdGsO2xjROkGtEXLk2D
AOcGqz2BRGWohRRA+WjuI5h54N7iQXOV8wNQYaNCd4gg7lJQzpiGrnQrKM9rPIiq
Vt1D8TR458gAaR38q4IVaajScZPCPmAsihKF8roXpOqRfbf1oiXHW+OXxQG+Aji8
nqSqswv6/Lao5IuXnPBylm2Nwz0tjf8LPR5umNHxStmEiJQe2LQ5T3YsNn5Hhda5
yz+Kg7Misu4kWTROcR/a5waFfigIZI8pIhDyC1dH1sGjAKE6BiSowWzpPids+BFD
i37iSWCNBGADiHjf7R3fLnwONEU/NnvATnyFi1WSEUguxQSUoPjt/nIecCGA+4yE
49V0qWjiN2oSEtI3l+rLSEMqBvi7dAaiTTUyiLRA1/sNHvBoIIk6tlg/hlcDoct3
31gosDe5UA0JjUgGgr8fON8fCx7pCTV9Je9IdTifSSmAq0prcAb8KT7JqcEISG92
f3CxUCoxCO3gcF5Mg48fCvqu+GuNMFgDsKZbKl1VnT5mspi/UbAXjXB3GH6C9U7H
IqFKSW9AYpz/6U8LUVnVGrPXYfDH2Wu0Gr0dYOubR8huXqhWXjSjvTNKrgB5Y8v7
EGkqzPQjUjUC4vRBXPgfmWG72hi7S6AQCHAfhLfd1sl7+Dupxkf1MsmeXW08yD5w
QmxiAWotfiIk8bfIQM3i4DrZlC9aRa3ciTb8477l6qafoFZlrDz04zQGkk7wl5Zp
p+0HOpWxPijS6D+uJY7ZTY/8FZyDMHuH9Jeeje2ynrfhUM4r8INUk2eBLrBL7I+z
RyOu8WIZxpRGAxaJ7V1MKCbb0A/1OdJKDSN+sXtL66WgYAQpmlAcSM1FjfTDe+gl
6KX89ZuobTmpg7iwxBvQmpRoA6GMq0KfZ+KJjkggwpLGyYLOVIdarRqXaxWQHNA8
xID8bnmNBT4SeQmaMg3NwFGx/8jGZseWJIXsm3KVQOubbsVJ3umWXVP+zelBGAM8
WIFoZRcdcbw0l/gal60+FXnHJOaO+HmHe+ypsHMqkBBBFI6OqlW+wOE8KKna5zoZ
3//ckEdpoMOwmdEaU9iiV+F0SvNzKG/JWFZ6FNQFPlrRwsHqNtWI40RRitKnHBUU
vOYbKLTysC8e/uxfO8S9mkzuyQjqpELnidlbYDHfGPvY8ngvI1evteyvFxdCnlSJ
bANa6etbIell21LP64tsBaJx9AxTH5VTm//X+6udtEYCMuLqItIWexy/sIfpKp9q
WcPsi3jvc+mKXxVCHZ/kgBSvikb8qWvLfsRAvJGyh8Buh+9Lci51/6+Ka7dGXMHZ
8B4xwD4aAqg8RaY3QHwSTwLT0//t2MEmVNgEdnIqJF4jUq5hJVfH7Q91vvNPn/3f
4wnoIIysuIgj69r5nUhh48DqEoHIBe2IILEqca3QXqrd/C1EMlfKIo5ZOWSyKY0b
oeyR2X1mKuy3nhdYLnywdqrGsiaAxxM1FE7D/LGfd5VbOYJcbb/nN0o4YcaH4Rs4
xKjKxjO4kbUyHUB0Ly12xLl0Q0YbVmPtqWCRUByN3xYONMkhuuELJaSoezjZuj0U
Vtm/PncUUMFlRrr2cyjGiU+NWh3ozpyPf6gYcpmQ9LWOYmgeK1OQof1j+xM9h6Ln
OztopM9Z1f+aYksRuQytXu+RJqowxV9VGAoMRH0Rv8QT6xQ3FKp9xBmIU53VitSz
e99SGoeiuq6MGA4Ntlvx2HXSy09Wyn8cg/+5WpPWXq6HJn4bGxFL/XrfBM8XJuyn
RRCrEpSjKb8mQFBhA0fdeV7d01Pip8tfm0ivkvqMDA1RMPdA2qtgTwhRz3OLQWaC
xK6NTJB63Zj77XfAy1sZXQI6Eemj1aHwIp8IMUjy55biY6m0sHfTN7yOZrLdNGb3
a0ZrFwdtyPyw7KZpmBOQrUu6jH8rEQKujLQbnEQHof60P+Oc9IHGzBuJjSI7UxWP
e+WflCCySHPVb2piRmdYPCmxG5k2qQ7Wnibul1l8I+HBX/yHIJ+QSvGFbJWBix9A
W+Nl/hLUFv7kcc0ZsU9kIzLlKy/WActKUTtdNc757xF6bbtQJWUb/VD/09CqHeH7
scUePbQRrZW4ij8QIXFN0xHddzEHvRe1ELFhGuvVdHZIXQbkISzgM1I60abz7C7y
k+0Bv/PDMamQH84dUPT6oLWD/xnX+zcKilWxpPbqu99xE0/W6OyqEZfF8qO1Mogt
qv7JYmFRj/WJ//zLCc3tW+HSyWPzz7aaQUKjLfiUy4m5jhh8+699OU80p8S2sujG
yizsipZQ7lv31Os3yqv23qv+5GAhjQioZ4VRwjhlDq0xAG+wGNYnSqur+N43wcpc
biXCGNYP5XWiLJCMd2NUvewQ2zAb13mhqcRMh3OCe14cgeqYk3624JtPu0/R9uFn
xti0VeUHAPZJN6YZUDocO+vHKZ0VRzgkhw3enQIy/pZc5PPk4pXstpRbIJI/HBef
j/PkAeOz9HzeEUlhIPazqoXYZfLFGxf6LoVWAV4FmO281WtenJA/1HkehjghzWdv
306d61QG7PRfFQUB5MENmTY7/b2QLFJy+oC1B/tRPqDiNqnVxNuoTbZPFMyQdXpV
kY9A8mPK8OBQ+zOlTycB/jD2s1RiURV3xnHelMerVGvPIhouTKbcD9EGX1gMMuzf
j30REBistEf5Q4tnZUWH0jgmcZKogtvq42EHMk0C52BSfODrdVL+7A1zrZoSw5Tc
djks8ljMZ5iYStSZcvH7DsrNOEVV0zhWXCGRjBJcdgBRV5Mn4Xvx11iCq0A9VWzw
OXoAhu/QO0H1GcLfrr+JzlP/+A6pq6lNtz2D8YZaImv7zy5Q7Ff8MlnuI7pBDOns
j2pBqiqFn1vBpZZk7Wqtc0XT7I7pXp5BHdn8tV0ZrqUlpPCpBV4shF4joqp5jyDl
rCQq1d7hTcAbKok6GkUpszkfeaf8rAfHA/HEWFy3YmaPLV7R7dJPMQYQ+tqDK4bi
PQYLIyyVMK1JCLOCEbwCNg9IelDqqlfEWf31j+t10PBk+h2NuIh7RtNEjFnE1JnH
bEuIUk7c/rv0VvAiL7dzcR78oUO0V+Ajz6yZeob0OxF8pvz0Dc0dCvD2F+EzAQrX
g3vA2ULzR22brO/uPn71JcekKbvIrhlCrgD2045kZ9KvW4GI0rGa/xzru43Nm6f5
wWkZ1t/wz/O+/NzRTrVgzbYWTbA2WyoOFzs4nrbtO+lCMdteU8Y72D3d9Obf6TaE
n8UzWobHKt1WaqCpgYSVCxRyJ+VXJv99QRYJ78FcgXJ3pSomuSJFTb7lDgq140Ge
bDzJ6/S5HgCPLC47ow/qm+PnMFI70u7YIUEkwT/1Q4fsE7aOyJU5Mr/u0TSPGD19
xvMIrAx649a1SPMhARyyVgaCORKSDYcWUKFWY22Qd7oT0NStAGFv0bD9TzZblzg4
9sYIwM//tEPNTFb8/FUVS9LCQKURn+v4SdIhz7x4kRtl1ICvbRsfGNyxwySTjlD1
KAA6GHXlj+luW2fVOUFxdiDdBFQh1DIT47AbsOL3NKG2MPiCUApYVFqO8/xedihR
Ya4osAXq1p/Gi6vHxWGbfXza6MbepEl5C0gcX0HCFN0vC2SiqyBUv+VYQs+VDWP8
n99xrvOXbQx66rnwWcLda+gW8+IBTRV5CqV4vAS30pklWTveHEadNTmu+6Pgtv96
KbqcBIra5yhQ+XBIsKRiMmuHIBVX0kV/3bKFcBCIc9teH9IhFVYha2UX2RtEDFVc
mCOWswLm+9CI4vUkatVXPKZRImDfPovyPmxq3hBoJihML2wrIG7EG/OmitPhPNwQ
CMNmIQQn1ptndSODNqmgANHKVWoW5ez+25gGmGl1aFoI+cTme72+rREL4rthQz4h
MqOq+K8beYN9KuOdZ6fowZsThwVSXMZmXEHOVsI0gpBcbyEhV2GW1XGOhntt99eY
4IdrC9EByvzEnIScwUuvxZjWJiGVND8SD0FvrvAgC6c1dgigQeaN93nvxVYX9aew
6Jme2d3Asp2/tZmx4fHr0ql1Om7g5twA5duQCEdDEhpi2wByw7EjNXv+aElWXXvn
Vv8yvgfDS8k6I1cCMF7dAEe3SCtMDG5M7iG5zZvq7L+L11C//VhO5FYc8U2eFlpc
6qCWJCO9YVSMTB9S/E71hhk9QCnI0eYJ6djeGFFbgf30Gl2eWiGptQvLvgIjJuXh
u21KtUdKDW/7YnhOM7vRkgDdp1RnpzKzP36h/643r45TZ2BMEdONVptxSRie9Hlq
o6sRxEgG0eM7Wb9nYy/iEeBb9Sk2HsD6p/uaMXHvF+Mm6PlBsgaGuJmXt2z33eIG
UZsgXCJXFdbO47tYdMsRV6DCEYkfKcJYDwkSjmoAq2No0+SN0vgvYtY2XGeyksRr
0gHNwE6IYpBBxpRB60EiSYdkfqbCQLipmK9TNMWIlhFVe62ZbwRMg1fy8TpXchdv
L4sq3Fth8gMKCbz/HgT3NOMvst5opwvxhTFbK6k1057sXIB0EKxKCDpv6YEyzJ9a
60W7jS8gVAp9q70uVjRvqUTQeTbativhMi65XGZbKBXsv3ULL2t8+68ZFroDntJt
kuZ+lBAuQMV9h9PwVVtKa9SEtDuyIrycC7KQc62qc3t+/JC67YW5ZdsOMfQXOGES
WXNzEfgZfDNLIaIvBN6RxoGkNcsmmPjU0ewA6tWZvdyWP4LtMXrgYsP90K8vEBJW
57YU5fpNOy4qzR3BZGJl+qAuOOlCwV+9WXYrzIpBheXE70MoFk1dCAebAS5RWrOu
s65OImB+WklX+646TY22BOWEmOpRgYBe3stYd858lLhertN03eV4S8C2vWsWDVv+
JpYQ5mMJKTurfra51LCzXtW8yI5XkMgNZS3JtcLR/X+5ha59AuC2WOy5GCBT6LAZ
ynpZGBw2kqKWP8aC36IMZItTjXQsuBo9pBf2128tzHdAaAf4iPfUBH6YcDgfl0nI
lyscdLY6ucEah22/4pErHf4r0KtIvHrFEh7KFgC8Ppk8QWdtkOelwCAF31f1h7P1
9fI2/ymjPWEYcKs/icm+I71TrylyX7oQpMKqg4ttunhkGanShfyP9RIatjNcw5s1
zMtDRihtYDbie9mXjXzO1V+9A89QMLsv8IL/2k5UW8l6HZTOBz+7t0HQQ4shJ7yC
3zK2rBWNNlcN9TGkNm8Wx8JX7gNaNUx7UWAg38+Ptpdae0BHohqFI1oiGkpm2a+u
nf4mQuVjKzEB18zFYbSbkW00pwbMDloR6cw4SJM4/SzMwOV2gjC4WdsA/8wuhDlw
i4sklk8CbbOAUJEvLf17eZIV91KRgU54kTuzmJfExeVSEQRwumw3n+MqVXwCmX28
1SOpkNafKpDOyAT930r+9jrhtKiKCbE4ZjKJsLMC7DHPDnO51HqedeHGni130xYp
cFV0Reost83WG4/GoF5qvvfd/xR3qzSwXqR4P8GAjczb695nhVWAjDgKBjOdYkpR
O4W7rpjiIEp4Ld7dD3sYKifUaFnG1xtAcYHMbBIuzeHRcJ/ByW80ZMFj23/NJBXx
FEwDs5qT9juPEUrkZOq+atysCxvVu56vFR8jGMb0mMJmQQH7MBPQZDcItTWcjh8b
XTrg0+WkE3L+orzrYA3E+oY6jULBSDZV8axSMjkX5y6dMUPDc8P570UWoRf4cIvE
Q6hspCawhW2TMJ84tc41S/u+K8Hiig4NZLvVfByEyd89TnyGMsyPJ39pGK/oseRe
NIY6qSvcaz8mbabeUPEoG88UHsHgXZ6JoAgJD/N1OEyc0qr+slIwPq71KZpWGa1w
wgLlVNBGiqsAxp74osF9JSn41h/ouEsP9A57pCmpwW6nr9SAgwEWaBRLDhTjSUm4
2+ptH4XlRqfxKmiLLdhDN7Qe+l2c1yQRad0qMaeezVAEMd7TKYxmy+3fwtVuQzDa
jc0F92jYIPn0CiHX/2WCfI8KM1ihYwRo2dpAj0CeHQoGpipol0omRGNH/Tlu9GGa
/iyBtTyYKLhLZT9b2sk69IB3UMWrRP8cj8gUuZ/VjI0K4VZPCLKm0Luq+VNPAXRE
Go8AGt7MnmyL+vMwn6DUb16TSzYNGatq3hb12JzAHCWpnQPYBxJiT/Bz/s+AexVR
X7WQPqKlsavFY9BVHDUeERhleP5O6Z5huTi8xD4BUQGpA6E0JAOgJRhzGs93sByv
3c7D8ycs9D9nMueW4+KhhDW6Ddd9zt6kGK9q9FYQg0OOiskurqKMncQpJ22bTklK
cki9fTovvXRINrNB/oLOYnfjTchPR7W69ouLjrQkv/4ks4alokjdEl7ZVfPPpbET
pFsqmZfjeKkJFRPwa7U6YuoJ3dvnkphuaSqZQLyzGIojg1jPw8LkoalISHx9mbhX
Jg/hSvyB1E+m9B82JYj7Ahmc49XYV2bCf3rhEYTF8b8g+r/2FD1o3sD84Exk+Xw1
asrgXpzQ0Buh50fkWKGcE7ElnFafPotqbBOFcdd9FgLIPh8oEAfvnKBP+l9xIohH
h+IJtc+mK/iK5p4WzLOYNJXDxTHJLGVclj+jxAi30CBvqJc6arJe4oubdOZ7OEdG
a8RYhDpO+AE1vgY7f54OT9XyN7nbQcd6kOvWzxJJQ25WBn7bO0uch5u76GFxZunh
4QHgIkuxQybe+6X2kLlA5qWIJlSjwHd0LwCu4W+SjLElVv/OdnxZEYl3hoeBZBv9
jqXG4GcYIl0uQZ5gIROg8MgmDLprhoqi/HgPm2JAftzKd702KEM9hG4v4xusbElB
/w87bnrLTkLbyCJ5a05az2uPAop/Abzf0JP5tzMiR6Ry9jLl6KmAQ9yRLO90IK1y
LD1OHxyAZIcuydQxWKLzvZpzofEpFw1sDIj3WZlooElqabWXezZoYXqFHL+lE0W8
CqlpEaFmYE3e8m4X8Mlg/ULH5aWaLC7a4XCLTxJ2Am6eWA3dIFDFakEDzC1RJS0a
WTNp/n+DAZL/56kYHkDnkEQcME5GNgs3yURQbjxcgK5V11lBGva76ypAQHPj8Nvg
jTBxDczXqrig8D4bykKHHwWlMfiZaNT3A+oaL7NZ6fHrbXmphQS6f0vqq+/Fnnhv
M0K9G8s8E7BqsVNcqwx1NzoG50O893fl1cIFLYhZH2/JMOZ0nNkrkwcXkBuTeFo7
6ia/jReWpULjqdVgdEK5DCVky4LaSpedvTcqmJGL5S+87Hkly5XxO5ZFTNLlOdKY
7CpcuPmTobo8sooBTTjpo8plAOkyxWKsZc4ay8H13sTlragG/yxZ+ek891HyFwSL
MiUZufCV5pULHyJ8UatuRh8azCO8JzCDb8hoQheLiqRWuocvXcdSiVYVBe7m8ssC
32dsz+JG0pEK9LUGTqz9f39Z3zVyf/pZlFVTSw9v+PT3l1ODFj5U2cDM4vOH/lZW
Hb3uztlQyoAAGy9X2huanpf3A/e0U6P8AdlbOQuz31IJK/dR7atcGftvvEBRjHkc
itsc68po74MKNh46FSD2hIY552CzDWeLmumGxx/HzOpk7xz6TlOyGMFTvvyR1Env
uy07Of+FNm3QZvz+JkrLI2maE9bPrDMV7kS7OfMdgrz/U/qzjRwoSTll2LheTk6m
fSItdp1ZrvEpxRDChklKMItfgWCzg3Qm5r3zgF/efaQiA86QnZn/K8g2RhwiU9Wr
D4otKch3DmFDxr3eeTlrcwBvIkLPaQH0EwobA+6tjGoiz0vaXFoSfz8OJW1t+VwW
OAZzJaEZuR2j9H9lwc4iFVH6fgRizIK+O2vQJAVTyCPskE76T9I5DKve6o+O9Rtj
dNIZsLiamkX1kXo4nHCufqv+h0JzKGKeDC7tfmv7rIJJmk52FvPkO2lBUYjThZTg
qqbBN/dhNdP7tDvKjX+imzpXAwRBnBhc8JvifI9DYIgaStt0vfz1CyB24CkuB8LM
hO/P0g72tXUC3LNySyLuoIzRoqLxZks3gAwq1NzmEWFa8XG0zTD75iwvPLpRCaY2
KgqOA9SLBGqOhdZyCCUkEw++2MQcCgTPIXZDVVKutt4Z8oH6o9Xhp2IH9NHKybzm
+2jf3bErW08tbSfFN4mJ+Kq2Xo99fdcdm8heNDrIKSYxR68hsT/rKYYpMYrr8owK
H0fekEpxSobEX3Fz5fyVcFNigkqYIS9EhIxQJDqatrFmpBOxPlEK1eb56+jKkEv1
re+I2lcYjOgIuI0eDMY3+8AqwrQ9Lhlku5bZhlbx3s5HXbCdw43VLFUAt6/LSJ9G
NWvhCDJf1bih+/oK/qWg32+9Z7Xi45bomeNtunO1oHdvYKbSQKCgjAaitKM4EO4o
Gadx/boVTU4q7swGg/De9eRylKA12hP3spxR2W9C5v9DzqvLk2o5Sf9x2KTdlnCr
eh943gEcHBpL4EfR/d4ZRZrPB+m3KxHFBVa8jawQQbtB6C57PVVncGnjt1XRugXb
gSJkdKqkG6fP/B66n0ZNRcoZGjALeHcPqYBWi8XrZrBdMdsx+pIf5MVYU5BGGVHk
VaBcXmkGLePuI+RKGlittg/9bE9gqipE03wnreTjCs248hrUZqpOJC+U2h8vQ2q9
Z7nuoTUfXjnkESaNxb9lmG6XFLLX41SSjJXsfpnMByTJ72KG8DZ0+2LzGpJ8ViS3
/oJ3hGFO+4ViG2Tx3BqJ822BwnxIQIHorYWBMnmCIjByP4RRLjreaDe5HfJEmd6e
xJB3qCHouS0wWdTo2SxbFcNoPNHziOQqTePAteA35j2sj3GA8ouI84UTYM1dXXLs
3FxBRPEtgAP/SaQwyZZsE6wuQ4/f83cK/qqD6BTrYrkceLoy9JbjkSqOJiQ7EJB5
eDP38rmkOJWjqcMRgiG1zI9Xk0PAq9NRMw6oP42ftI+gxl9AtDZ5VlG9V0WLrQ9b
PmL0u2HRnlYgMepzq3MmMuF+AyapAx+DNGH0gwg9sjPuGDngdYkgs7STlQSj2vjT
L1opaF4b4q09QthKy8UGcM9sWnFkrwX0Q5EyAs4i7vDcL+126xO8naU6MwLeSaUb
oPx67jMk6Df35nU3rXJUIbVT4W70M0PwAhdC/RsHok8vsizT0kYfRNRY9IVGobwx
XwoiVqMNFeYcVzWPNwVgw5Gz4caT5MguTOt6nvylyS6oDDnSSFEof6vB2OJ5W9ql
z5wNFl2BKhwy/16MUpBWR6/foSvA9ewF00HBprbVC3z7DRTR30vEGqyfY7PA6r0F
MTicheKDmlq1ZYfZv+jp/g7VpjBjql3R3oX1ZHKGGIT6SxRF3HcC3kmB23QcrDaZ
Zfc/Wb89vZWt0ISxPQnYSsuvQ4Jk5CT1Us1ht10xg/snsL439Wnu9BMFn5aTOvWh
Y1qC6Xcb25r2Je3mD1OqzfssoovtMQIsVUjZZwWs0A2kPCQoo2t04776X8o1lYlv
F4LXLo2nlkS3KhgVDh85876uo8JeaFS8VHNFbQ71C8Zcec/5UJxuDnFmclWZnd1V
yhLeauvhCHF1zRczkvqJVlcQLg7f65afXvdjSQ1iTrCqIARm0Icy9/BjAv+0XGhe
csBhtWTUOX2PrwcJnWBNhR9JDGvRuDghysDds6l3/ECN0m4ugKYV3aFJ9N6/5Ihr
5immsRKwBPC1Rejxxz9ju/Dv6mBzULgjFWf42mUwaOhxqnSCAiIN3JLukaHQm61P
hHO41du8xBYJm30nAww2mq9pARKaFndO3oIGBBO2ZveWb/rFP0mN0bfUoOgALj8Y
ojpauUPcxwb/7PdvyUkvQslvbsC5KPZziFpPvhHRSMi5bCDvySVZtcZhuxidqjIE
DMD1t2dqs3w5gdZdJR1R/celZuI4XftH4zl74WAdSv6FqUbkxCoo1B4Cvc4vwH9j
n5XP285vQCf4TUYwjTUomVQP9GiycUFNXycD/9rZ9cRUYg/Z2RZPLaNnA6UmWDMq
WzJ9QkNOqkXwUB9PILxMU/T8ryZvR+ZoFwNCEnEsqiSEzdoGvBWXDrTjsnvyI0Rf
HUbp1GWxFaMrNTOdqGZOkWNXONA6dpzJ9V8T+xXlU3O+pbGCy38Sgz1cBx0FhOBF
C9FwYgC71uZAKP8VFjOg0UomFeXs8LWJrwr4gEtN315xE3gArB+1JMBo4Hh3ej/6
hJU3eelIpG+YZ7d4y2BRrcDHfH3Fk2UTFKT7oBqnDq+Zg8Uc4S1d+VmQf+MtTYUb
EBLad1BYkPXr01yFD75PvWNIQ32Q+aQl92iAlXBPcP/OlkGev4KHWVovyjCKT18G
T4gpeFyK8KFDgJnoQRwRCDjahtRHepTUFkShJ6a/yBVVCIaUhjikwJXn8+U/CuKs
xUP4d0sKJ4Q8TSvinUanhFGZIlZMeEdejlUdvPwbgtA11vs5vva+/qcB1iyQAh8I
3D4T+3j0NxiWE9x9enokVGp+uFY5Z/NwobqJyiherz2GU+qIR2z/ZkdOisVc5WS6
TTXmdmm0aglONl49k7QHS3YXbcQp3LbyrN57NOPhiPuIng8HU4b2KSBEY63jeicK
yMwPQjLTn/fjBXsSBm+kGCVlfamqgtmqQhTzzdmwauRf8EgBwAYEtf0n8yAwrltv
9swNFRs6/yavZzQHwAPbOkoyelKorgSclergfzM36UJJleQ9iczoF1KEn6VH8toT
ChaqZFKo4ghWleK/UY0EiUZx6Rtg/s3R0w7QSefPulZUWXaYmd2UVyCEMJ7sqbdB
VYHC6I7Ix3bw8qWn1/lATmoJt55GgfDgTHKT7Urn/JNqV7HFleF9NSQFHtF9SoUG
+rEqgre7cDP+1GP/bZ3mFB6mmL8AK43GJQDK+0WKOGyznA3PLM3RVmfIo9LLYAk5
gae4uBxDPy8X7ELzGQtR/gUIA96kiAXC9KM8VmcneZe8s0Djuw1cVkORyjTXsMl5
Opf7lakr7O1qQd2VxkLRsnvq5Yee+6fqEKQUq/95v9u4MMhvLkeQ9pfIYnpjZhRF
WD8OotJqXxbe5dAkFc7ahD69CRjLFLLhaXwSljQlqbGf6L3S+GMlLha+Aw7aBHHf
HAyhpy+V9EeuzA2ehhBeMlUKoKryZec6S9vlH0HK1kFLvsVMpbKu2hn0o2ZHa1z1
KZqIqNN5JcI7ROspKTSG9/6jmdlJTDWCY8MsNQkMnBGhC0rLV9aOre0KHC0Id+7C
sz0KQAW+jwLwRjB7u6y8DwSIhr0eeNSjHlsMuAbMQjKoKIaPWwkor3Fi9ftYXWPf
X6mFK2mmGP4Qef9h6p8MXDTyffT+u0EN2REmomyOJ07g6xAbA1dsaj9G/yiWIYLq
i3EfIQP62jdVzTwTluc4jqhpBC5VLY/Iqpo/hz6gu3dHQE9s1xynv/XK1r1wPiKx
vE/p2btQ3W6Fuz52wYq9WoErvVk0Milv9gk1rVSaQ7GfQD4aPwSYUEAZEdBC/zDD
T1jogFNHU9un3ZIBDRXukPBSSrWyEDVMEUK34OaHqOppz30QKnsFQX12Parx4i+L
vS3gZeU4I1A0ztk2xo68nRZsYnh3nGmDDjrxaqtG7kS9EFI6PSdiOvzKNVGqn6hf
rMqhNNEqFuIU3MEgSeg0NZjPkUi4x4lmTxpxkX/PQvtvRPiy2X+69rN9PA62qxMd
MHAm8Y7ppZMF+a427mYl5D152VSOsEc2iYtc367lmeeJnMa4XufV5XK2Zw0n8CJB
ypHKtfKXMh8hBRbVmCS9baf1tGxUFaDUYitk99ybSAiAeEBtCdMntOVPmjsmD66G
HpmnaCvM02iC9gZ2wlcpc79sMo4Cr2eDZkuhZfic+GanUPM3VfgSlHrCy0YoT2Cz
BeiZhNhYaCg2S5kpvIjdySOJKEilPXEY0DfXLwB4NHqXzFWA1dWDQzhP9tcaZSHs
KrOb2/n48ZADlct6efwT2feGHq9AWspeBzWgLxo3ZMMmuFyJ9ahdKMPZAZF0QCib
GJyYL9AlkkdZaaRkoMA1EA1Zt/m3TcKveLJGqa1cGtJCaNHmjwgEZWzhuKDyURUt
3ILi+xKOpR4EJXbfwdq9gg6z961pOF5LatqO38PX2GDpH65lNK3jEw4kekpHB1ZC
XxmW8a5LM9hU4cdSnf42qZNL1lKeieUDsZyAiifQo3WL2c7bym+JmV2sY2al2mYc
yXqH2zCirkRg5LX1xMnUn6WezOAcAVeGk9iGDcStI9qpXnhej8XUjZrhbZRV9z+n
MD2fYIOKye/RQWpAQuSFg/Pskd0WfBA2tuY4jcLZRp+uj5cRA6j/vUiwu9ntnczU
r82eHpbrBmI583JsUEuCVjKUv5EX4X9FSlpCmY2YQ/u22fd4qHmuUk0OMbl9Q+iU
rAlapPOiYDkhhrmk754PjAAc9RLThfHjzatgD50Fx/6a6jWevqW1kSy85AIxCGyQ
rk6jiaFOQu/MN8QaEdLxpUA0i0JiYa+sgg3PipXf/FltE0/pm/KDPqb0TChxe16Z
xPECEIlc505XF93FARPZJWvszEqw/oqlMmmCWB7IOh0xCJmul4Ri1TEbx4trLJF6
Q/PPm29ys0vyqduQHp6dXNKJjRAEEuPQPkXqxglr5KDX7SnLsNc5F049leuEjM8J
R65IKQyzlxy3NUo9OD+6KoIPE3mnt/nKy3W5B5o4ultvRoWpU+XFR81uc0iaOlV2
L4IVhKsJyiN4Z3o+nUlZg1LF0OvEkdMyvLjsAjX/LNrOXRRObr3hKCsU3lQ61l69
VbPh+Qbmx5fe9vndDKvGN1+vRKypRZ697kzkYpZz7d6nualwVt2TXiVm4MPkBMde
cSaRrYjDqWrpYzn/7quyKeK+QcsHkiS1vLqgOYO/70frPaDWsG7DBP5rCfzMjX4M
9HTyQlAy6sd1VaFU5Sn1CHXnpvsw6iKb7PzztPub4JB1NJXP7OneaQJBiLUV4KoB
oLSna5MJO1yIFVs4lsJx1v6fWpuKkaAI5e0ESoGabCrSggpyuQoyQgvxEf0LPxvM
5lwNju96PwwTrc/9OQOjEnkonayjKwe04LWYOBmeI9P4KtZ7SJzr3uJCRB9lQKFI
/QW+j2N5ixdjTx1fp8xyHKLk6k1+S8YnlZlAZOO+HeM9OHi9XmcTaEnyqWQz5yq/
xrKAYUWFGMz/k85WoS7fNexEDochYi8oH72gigXol7oaCqml1Bjc7oGdEvml2TGk
Y1BvAI2fLb+oCP1CVkFgtdRebrugygsCnMX0s+BgOwxePW+qQT+7zfYeDzKNQRw5
k8l+R7VBp8gkP7Lz8IllaSz8ky/Z5YzYhloLBZmqbo5irQCa1IOhs/++9dmkWAkv
wFr4EmjdMR5oPQb9FOVxHL7zXE4kP5cNYgt3wQRFEtZw7+5jEW0Ur4M0WyTwYO89
dNK8ZrVFnPBdY8oDpG1hox5Q088fIfy6cpZvm0CDRt3HL/c09AnoZpXy2eIVt3Cd
dDQWGcf7KkV0FE2HVv/WBIvHDVzHws+uCfrgW+EoXXMvabKcxJ0PKrqpj548FlOS
D+EALvscokWTTxlj2GysvdOG+BMz0BnLOVdZeMzk2mztY0uw0Nd4R9cWIWddNf7Y
n5rZoZPGwSvfvaSpOavpk5WhjXUwKJMlt9Su4m2fMkHLMm2rpN8JeU37ld6IcyQ8
kpts6a4DMBipY9nbya4+CpZ0zfK0MlqPYcEKomn1d3NFsvJ3txhQewAqJk9ugQDj
SthqZLaAF6tQBB4yrQE88JDnxh+7dwKshGy+pPkWmwXI6QPsqsC4ndYMxECMI442
LQXKRX6aKrcBoAw4MXP45d2yzHhuLfP9+ZVGBnrcpNNeigK0zgudocgDtukIKb9L
582UlFp5bquD8qvcJTCag5Q7SyFICdK/12CEYtnLRxDGdTHgZ0xeMjIOxg3B+3xR
8so0a1HCJNCLH5k9LHfW+jYtYe9IjhyRTKZczA08INtv5ccQVkq6LLeJwK51V5Vf
4CAzoWCfuMD1zb69k8XIRWdv1A/uFmYWVrAs/hIs6FoMTRUehV2jJAuBh0A49uFv
znqm7Np2RIDVV11pSLGuIEsAt/l6U3bs7wvSU2QFdz1/9lgN6z/2B7/GQU/ZauEh
FXDK1d+sUBQP3OibZGxuXttd8w02uIwTpMXUeEP1JhZwRD99tKLJ9Io/h5wwq14F
+SRIF6uPKO3hy+BWFMo2ZmU7k7l7fly0ECCuFc7vtqqZ9xu2ZJaNRRElbXioyrDr
dEMG8/OO05mT+68L8JICrHDjlw6d9wNs9srNd9skz9QYGYvdevHEiDf48ywMXWym
FVL7J7Y36zwK9iFivt9DnVmqrFmvGNbRl/wsy1Y3OH91lxWgbSXh1Ng7r0tNk/MX
8HGaAshaFzAcbKIKlT466rxR++htOMVTQYVk8dg3ondzMgCOJfJ5t9ThVIrVORFy
CquIyolBnoIiBGxfNGO1Ch2F7Qc00ZL+BOhtcPoYTfo2rYd3jp6grp0aSXQ3I7a3
0T83VdThL3hRrcgK8o+1V5HbjluR7/JPo8hUYowrZgXvmXx6ZvvrPmocVTdHaNkO
NPDEJro7rF0MalnkVev6v9K2CKGpfS59AaJUEBPDdCx/rCwzuQxDOlheBhxD0WTk
Eg4f6qlsiBbL7y3bVA2fnpP9anyeCwD29JOGhCD5pTa6Er00eDHMoCU2uNthwK+X
b8OfHGjZgxqEykDqyGK9zXXFxkgHZg0gVnBK9rMM7VluahT6xE+qOkwgZ78sMlQF
ZrjOKpy5d7cQ8BoHKmVn+PzB9tAMqLiGoBTi63RxxZZh5KKf4oOGMflEhRoi6yV+
zR2lu9GZUdGGXRUa9Labq8cz3SaC+pz3ZGXgJkr8venh8rxTl1PxlDF6SgBMAa26
0Jiv56wC5hruFvw1gDwPKphIGWCvZewm2KcF5U8qegNjy6dR1044+wX88x5oeQh7
1hBRKigUaUboEPfgC2Ulj+6wREXZ01tDpudrPz3Wpb5O0ZgMhjSM70X5oKcAIk40
fAD24HnxDAHAF17qL7AdHIEEF0/g6LxqBla6uNCf1HTeSa7pN58/deQGoE7zY9xz
lgWd1KiAvSf7vDWS8elTlrR6MuspWvD30wq1ULfffwydFXxmaIaoqPLjxhGwtw/7
HH0MNL7W15eEkBCTTy6aPK1Dw6FK7HK8ZxoZnoFP8cFDSeTwrVB2vc6njzhCX1St
vvM7XdXXje2rF6u35b5dwyu20gc+ANIQ2mIomHmLcble13oLOCAcLaOMQSLLt6hR
wE+OVQmzIZ8M3QNZb8DAYGnH9m1oz541IkgGOdXmVvfr+MIZmLFSVz7njfXXSCqA
qPjFAzsknhlFHEB5wzGB2A4t0yYml8SXI0Vfbld9eji/1o6KV/BXfqLp9a0svERc
lGPbvhNjmgkut1BK03VHewzCZ3tNf16gXtyg8d8mkCnsobDcFL/9LefekE44bSes
T7K7G1Mn5656gr4WpXmcJz0hEua9pxMmYbU52gq9CCTuofSRpIV9ux71O+8eSq51
9P3/JqFQ+uCmkWj4qfCf6ZUcQ/Pyf0aaFy2EALh2VlzyYib0rQYGaiERqePz02b5
7zyEHM8Qxn6KqjZNAUqN02bzDfKBtUErAlYenB6KvIYwLnnnDCDY6Fmj9ZAZJuv7
Ghs0PCZYaLWuk/h4zsZwe/Wx4jBcb5Ocxfqi73QZN99FRPEUFAMYZKbZ7xHW99LQ
EacP+8nHsiB804NURliCTftZBFHTNBSAqe1SmfD7K+ioi1gq18DMTkW70rPJVieB
ASzFkBO8+zWjWaLoW7OYTWMd54MD1qqCINzIVKeBRxVDAaT5SgGcAav4hkX/xekf
d9FZ1WWuUCTPRqmptq17D8767ay4MIBmLotHOkeZrCnEhJgp/etUuzHy3B3JgFib
vZdaZ3MXAFQfp/Bbjqmq/eHP28yi5pX/TQaVZHSlfesrmDHLGh61Zxq8Ok+PQFEK
ZsUPAQRfSQetgQnjYvxAmUo+pp/UT9qEiNVJwdTFncC71aFCR535n7v7oKf03ag5
aTo4DlaAg6nHhpycwA0wDJgQvwmY47B49f9kqhfkOGS0spWZy68dZd4PjMxP+dAC
GLJ5bftt5yRd/vz50DbQ7d+8e7yJ2/2/TFXWdmDJ6lAc0K1pE9GGQBtbsiEwEDZw
HssYYU58rurtE4ceVgbp/7M8jLSkzBckLZjE43siZimT0/b5XZQyVOAr1C67pG9Q
ATWR3yl8uquzqJpRd0b60ofUyWcmttVqjgOfI6zyD5J2fqss9F1ud+JgSPCV0qNT
AEd8Jex0hyPSmBSfPMyPDWot676TZD9fQYmegvXwSopyLUdHVWnEG5y/Pd6HlGZE
/5I5bhCo/zCqAV0dEt8d5owtxfDz8vOLeUCVo7qNTROAYOJnXliJ6PDPxRsiEMUc
/tfo9+NryzafSPkFbIwOCiKqXrlZ2kvORAZP5u5pPagCkgLRFnhLcGKuEl1xITCa
ax93RPmN6o+m88lX8cFtPJFP0mamYVltbwAMFEP0ll73Oxx1Uhs6vqSjwQG0hLAD
SXzrjQmZFOIsz5hY3J44LJU9a6JtTHAj5Y/StoEE6TcmvFh93KMWMVPUsS/SYF4h
bXPSOP1yIiki6Fp4qGmlvpIrF5s223Gt/FbUQlPte750s+IddP0urBIMu/521TRn
PplUWo8dC4S7qYITFYsQxC/QqiLuC4DTrieX142sJmhTycGuRSeAjRVbw4e8TGYW
5V9GrRVlxGKvKtn+FZ1YeoyzLY7eWlGbCZS99vuWjV6RkleVYAy1f6dfra5YgNjb
cAX9xbICIeimHc3VY1mj/CrcBYUWf30brlORTST33QIGjayEELp3a9mI10ar8auV
yWLTEdXsgPsFttRV9aVadV3Fj3owAK/YKXOPWBsRiCMRp8pYvF4qzMJ6awJa4jfe
1YGTVvkoCrmQPZgC5wrGBeFRx0DgBD14qiCFrTscW/hQ36B+Yw/Ef1Og0VzreDaW
3vObOlv9zdeXnqTxZZ7dPiO2dVCXd/1BApw4Ky7CPakbWkNuVyBGkEF3qjvmcQPS
bG85Np8+xfgnEiHEFrX/kXraaRqgpF3B7tLh420tlznjIYki04dtALCoj65+iOnR
j47vcuFbGTkPfFkkuqj76ZhK1TkXRfDHisjlrxmQmsbfF7lFQ++y2wVUuvCRosrJ
0H/bV9AmyjgSI8++Tcr/12huFoMheZAq61cgkEdiOERBSIxrBB0nw2AF/RhbKw95
2xhb6nqiazcwQwBdHsjOPKc3R38tj8QQnXOGuSMYe1239QkSiEn7jFIQwrxF28uK
lp7VyhxUE83qGydfR9nmNA8k6Ya6bgx31QozlH7hzz9v/ahOIcXCf00yB95HcjDm
eEDcLVQmnespMq4igbjKcvnqtvWFcfdIYWS2ZnFjIh/f+V4ceCMGffydx0TsLiBj
f7alZ54jYuwtwAJC/B9I1P7Vw4YnGx5TdQtMQGVBOJZ9wrnqhTGvx/z4/UAt3F+z
IjxfFdmqcG2wk8kmbXB56qQhTyt5z0HrjW78qFDJAgNZMF6BhVoBKmzMWfYro06u
ksToteQKgSEzJmsWmyPwyinz0u+snMGj4ZqjCrm1t8iDfI9+KcuGgWjkZMYC1wQo
ZuwvQnDOQbL1Yr9UqCWON7P/YnqlJRsfdBQOCV5cPy+ZHLXKub5wZI8otCQNXi1B
Lb8tuI43rAD2TEJ1MpDJrN2cz0u1p6Mlv87eBVvdnvMar9GGZ/5IV3VcGIbVvO47
nOx4kjh57d0ycZlBrdC5g8b+WGrQuQJTd36ZN7mdfUOASvYqJHncI37z4geZw0ed
BKVq4qyAiaiZHnxIYAuKRw3DLf4uhqXmoKal//3pDn3ZZF3Fr0jA6hq91alpyKEA
D16dOETWC5CmIV52jKbRSlyTyPP3oH85eo+sKmX9wq26150CB2d+vEUijxC4KVLH
sgbpBU+v+tWYD4N5y//V+ze2kMg+vVBVoU8/DXhN2euAuCZw1FdzcVQJZrljbAb5
CkBNvGdFjCnuFVT3ATXLUJzsfkXz9/GSgkJfxrFleGBKg4JWNRCIuIICnhpEpNzD
mpJzPcuHciZkS7o3dCo6XmmT8iekZOdAgEzoja2nXjlvpW9bfs9oq7kSKstZSBih
VFA4ws1jZ0F2UPWjT2rVJRqJlvDAH30DEDyaJJ2MosO4nJyDYCavW18Z5RLUPLBE
yoFo/ZSFvwvZ5jyMdsXxDZkL5E4QkHBHDamN6fI3YcPmy0d0ioAzA0mmg3ZcMGkh
elqsfQai0AJypxTptFBHpZAVNaT14A/8QEynuwPlY8cNAzwodbZRDi71g/g2DVGV
LawociMq0Iitu/BStP/8IuKq2FWx43WesJxM28tIZBXvh7gvU/IU4q9KfOlbTflw
XLa6U3pgbUCpCoPXGpNnbtyzorC3rJXlTIJ1RKGz4VHyc7prqGhFJDEhHRbKApvu
9Q3Fvf8v+xdQF0wYQtzYjB6w3CUquk+dlFDjO8+MXzNt4hXpBDaLpqfI7l6+YygP
Qm8DRvsmhC1LN4paOtrLbmCG4ARCMrwQQfVDkAn/xC6mdZmcmIBuYEpXp1TDRSrt
uUQ4TN3YYvHcRkGNIXsPBY8drlXzx477acgT+zeDKh0wmnsDnLEZ4l3XXo1Lwo2d
hFdkBS+nYjA3L4XZJEiGaiqYirDNn4sK9oxqu7j5zxhIacG+qmkuBqk5QusWbpB/
ASdNrbvuQbETojf7rJ2FfhAQnIhN8h/IO6Ii99ayZKiF35C/REJyoBc4VP9IpdaV
LmyDFmZkstlIsxUhT3JxiJBq4dfUjB8drAfPwF1Ngk1Ge+038JJ81xkM/sBXBnJZ
pTjWkFGQRgsoWdXxq5iNnm8sqG0t3wcsbL6bYaaw87U/BwE30UkQaiKRihbi5LRI
OrkczPCMhNLFXzN4492YSYmD3ZLHhmCShlbKmByaOQbNT0dJrVIIfEpcXjpqjvXw
JioD4rOj3G5O73yl7ghewx1CGzB8cowtBYtHS33lLj9pEtiwzdoMMSwMA5LfRIhG
QqETWBK0tU1BlgkcOy1YuQXpxX+do9749Mk2u9rNw13zlXqR8lBXijq4fuMT6+oK
2lTROWf3KQnFDTTl5Y18kufN9L+FB5umzzX/kqENdJN4Cb2jRFQ2wWQcsm5aJoYi
uYQpO9wJLm9dL2xldvdnUYSNO2GIGfnOYe35qHaJRhQlTrl6oZxFO/Vc6ksBaMAA
bUkOSqUwz0I8mq1SRdXxtfLG6+9D65auSZ4oN0nKXnHZmN8Dd69TqH0b+Ga2b8wK
4iLgZQQg6qVntUEQ8Kc1OdAAMmffjyRF4JRoDSf6jnS2Y+yF2b9Gf63pp/+fbFn7
VW72XGaF2TfGZlN3hqSoqNdj/utoD8LGK5DRC0hJxG17tseLVYHHwC53n6r4s+vM
0RiMqqYDajQwPC57jwEYMcCRX/e98FdB1qmIoZDFIBkL+ptDfWGnHTlNIvlD1jJW
tCyzYJYZFwpH4dKOM7sXXWNnqyGT4ZGy4f01DMdRC4P5b+7FkccLXGTo9DfWQvwP
TJp/EIOnT0L17a983JZvBSU0B/BCJrBTcT4sUpYwIo9a39IcP2AZGj7fnmq19/Dm
63P21Ih/o4jWzHGL+rphRDuCmblVALS/ZH4QiH8KzWInAMkma1W8kkfztstvi9zT
5LY7bKx8eJJ1h0QPtj1WnirDUS52J3jfru3/4sN/QrtMnThL2RaEsulhG2CRResa
wXkx7+6S4HnZIHhnq1RmFVTnUxJuiqpYvTXrQZci67lo9L3BWkH+/QVRdwIzfbQ0
+eYne0kOi8n/PdYfIQ3yw+nezMtMt8FEkO8WlRz+YwWm82vkekj7d3TGYabfN9g0
2NPtUR2yljVW1F9QOz9odgysmN8ooUbALCYn5AVaNZo+4Bj+B/X1TEvxHDPpsxnO
qF+MeCXpu8F/aQeK/LoAORmdWwGuglHK3OpBxUL2s/N3O2mCjRK4EqnZ9Jwu/XiY
F8xv3rd4P3z4ddqOLS16IW6XnHIZMfZXu4Ge7D+lFAm6I8gyMAxKcv9NZP7feh6o
aT6Kv4RMJTIs8gqWSn7O602g79AJoyZjh2EqmQYPxh+np7TUQIjoJDpb4cnJPchG
cIqyU12/3E1V+WN15cbvA8ci884d2YtSGJ/j3ZCCu98JLPQCLleK56JxRMJpezBZ
sY57Z4RLb+0A1zQ8i2b/7JcjBEWvXUcmgOtfsVmv0auE+WeaDFwGZBugz2OWfnhB
ilWOtvtXcW6VN7qv7YHbfosVjZxFiMAjGmSvqOOgG6SD1ICRXwlw8PETVhOrDhG7
5VwQEBhwFN5mz1z1MvLAhEpcikpjnM+V4hMn8Nv3OPTDoCK9i6/dNSItyb0gVW1a
PdDPLn4v4VxSIBT/8zGAvlqawZjtrkYp8hZFoC0izGsjAXR3BzSvoSLbryevoiy6
oC3Y4oXkL1wvYBExHFKyRa+2re843aO2evyqynDxeQXobtrqJtebcDclspcrfaBv
Z7amw4pujbPbcTFL4p5uXatvHkt9hNlGNa6LM1tHKj7OaGYplTRWeRzIZQgEw1ZK
/hEzpEdSDmJbYHtHsPMfnFfOqQPipQselCZH8A+aBGId61GIX5eIDw9SZ16ZhCxb
XsNw6zsagXw02bKJnGv+SQyQNUhypA3ktBGaA8ARZubCS/g+zRlGcxCdMm/dGzf+
/Y12kaaKImu3GSD5EibEAKHhGSyOkEkKu5nyXjO74nL8bVZ699+c0NFbPovEONQG
X9e7u4hluI3knjCOye7XALwIn2HCthS+jlYdAD+uNTdsrtkLdTPyUmZDxEqs9krK
VyJkRN6ySx8WNa3fYOFrNHIGaBP671Q5g7duHulxZGt9b2FrjfgLe8QiuwaYMOTv
qc15QzLh68GnYcOnDob/ab+o7WBgEHdMNOuGO7MJFTjHYA80aGWS6Fdbn7TZSopC
MjnW88vU+d7zfb9ETZerDfMBlNdC0E3MkwXLb7of4W1PRyaz3mcFrVd3ZsG+q5AU
T+lFQRBvw6sx21o5fxkGWyf9HtM8EC8FKKkhcrJ8hGGP+xMCb57kqCxMyrdx7Fed
LK4FPpQNCfQE1fHgtMct4Zdisb+tRIY8euX/RJPsQxsA4/UVbADdHxa9m5kfXnBd
T1/uEevUjJre6ECbZXoR9lHFbY0R9Z0/IwTwNHnvgHzTpt58Eeca/5B8TyTXwkSU
lgduyF0OC2+VjAA9mCyedk9SvydrAZbxOOxUQTNaJKUDqZkqzdMhz9/tGeb+laIm
wcZj3UvwZ3lyyHiZ9DKWahTzuEngo8sfv7aLJ2otJxd6h4AbBUtziWwc5dzfU4PJ
ZIuD/acSl3cc/QNH/gTizDKh9NPMBUExmVSPxJh36RAmGFrl45YQba/fPIY50pa2
4+H1H4S+IorJtzZLMDuPB1DSEDT2WHAEiSu+A7zywlDeSG+OOLsyyuh1UfgEYWGz
M+9Ae8BcS3wFzKV5DBchEBoH7Pi3RFRr7ocfqyZp+NXLfRFTW+2kXnuybI26yKUG
HPXMgjG6Qfacoqt4ktkJ+lD9s8gWBD23C5Rtxg+51AkfUKL3Bv9kDWGgKjgXjFpu
UXwPoYqo9zndoW0QCRcY9+oNXMSFrmzURFSAH/5PR7CNR93a9jHhneoE9silnKYA
EM1zNvkflsKIWsZPks4BBnW311fMUh2Lw2j2EtU5iriWVVyKb77E2Uv3RuPFhCcu
OqRE5b4IRhO3tuKcBbz5r1V7MjJVC5ncTIgMtJGGE86KN+knOn7Xxn71eDJ964Vg
lBoJxbJs0Hvs7cWpTq39x2Z1smQ7QXPPeNErsEblymBRU5EbofrQEox/pU+YjAtj
t/0eioV0VK8mvLAuw2Q8ZqvOUEbGduEeTDF33EljORTNdF5Ii6rB8bc0IILV/YQU
A++yfcyTlJ4G1M7krm3HAgGBir6VjbW/VAdalSPhBjf7g/LWWLNF/ZpkO03OBVIM
t7yl7jbZ8PFTrmhfZm4XQVF6UaPNd3fh1oNvqNZN888crbwmJdu0hbgoODvzhrbw
JvmDDMdE3Teke6LisfU+TSrFY0VNqlFDsnJGYHzXmm8y9P6c4aaj5+69uwpT/as+
2eoUP3Oi3fIXIh+zXdW0h3py0daTkUbt1Vykexdkw82H3ZCNIV7dRsXg9D2JXxz5
XCNj9r0Q2zER7vgndpJ3ZUzqydYxq5hbxTzeo2W0KYHc7uy1kX7kSLH9aZCymb+0
AjjwR0mYf3FZ8/5wZB6Pk75Dbz6pzuGls+OmGVpA+gLkHZPw+f0C8X8kgeca9cJJ
zXtvH5Plz8NJQcxD6j/lBgIIObcGP87I74ek+++N80YpK2X1N6bcOINY3m5ixF2V
RuSMCbAfOSewBTyEofJvO3I7ZFjfsFYkY0mdoTGwPzM3N+C5YhxncY1ZsHz0lzv7
pm4csJPAOzPcproVrQi0Wyt5eCSWuILbifOdsz+HlR/PQW2d+iA/l/R7cMJWlQMY
+1SF5cW/mD3ML57QGdzqLWNly+0dkuyCN2by0iZo8qQsBsRBivZywJBdyEN0T2HA
ERM8HEC+PunepfNEeYP/n/4vRZYlGudje2+drBG7PkK0nHyrl0WdQxFhyf/ncvBn
U6msTBsbjOEdOvXMUqrhHDhGjmhwLvQg0xd4FBGtNyFJs9dop1NrOS9J1OFMEDZF
eJZtaWP2Y3RV+feYuWBGvJGx6LBSy825q2Smj4pr+0WPx0TcPFpCtXC1YzKApkDJ
85k31XlQ2Mz/BDrgsECqMxdwl136+5QE4EWturOvyz5h65AKvuISWO/aj9Bf7l2o
HXIRWhggwZtGDddtiIFgB5FGEQQhF7s8prtLB/yZl3qFZIOQhNqzJqpiKtJs1JpX
weAbBw0CC3Xr7nBh2lvbIPbSPL0QPcW5dz/Ex44hkr7EJmW+1ZLKVSsxiYrIkeZ4
REJvHLjQfSdEkUdLqXib3HFcgPA/5uUuiIo6ZcVY0SZO5WOjo0pKatxN4iJDyvj0
sHlTaxjEtn707nYcwfmRI54WLNYXu8Bu2WSATh/jdsXKj5pJFOSkdtp5dxB4B+IO
JeFkfKfEO+7fVA31NSaP/E+YBvntBN3jP4ZFW2ryauquCHMKzHlZ/tXljE52IeuW
uIgmw5c2t9aYIAaaRkBcWZpP7QdCnj2kxnOYFGlsVhYcFlUuGRfijA8QEGk1+C5E
caLnlivR8R3uxZLegKmb06TFzbRcWsQP09epyY8KzAOREHX+GrGo17RCNdMf9RQy
zImzqP69J5/9mGvduiQwCIbQMtjcWKEwv3xKlp5erWv4iE8pM6zq0s+mbW768R7t
gGGXE+nNyTIZZxWUarD7/yVbaFKkz0iEzcTBIFIp2R+KVsh7l8JWCwbRtfmOzCsu
UAcNcSUCMGkxxR/mzrAIdn5XN2s7RI4gJM3LHyVqLzHJ/xohV+f4CUSy3Oc9qFXY
eU7ovIQqlxW0ILvQ+XZCQPWBcQrHIzTWSG59gSFtL0Kd+A22rXeF0Lm04bmZSk2V
DWssz8luycM/vqnD2GcPEFwuCAtEtQUiKkqdk4v7mM6K4n2211mUJbsVMyFdYojk
VHllVvwPU+gNckY0eTVVbfbmbkm0Hm3i4N1yhTWr3Q3MLu+7nZGSkcNI1gfUR5AI
VPAw2Z4JBugejrCVDgtJeR7VkjpSF3e7zKC9h5NGkA1c9WVKuqQetrkDaZ0iCICY
a5E9RvKvj1kxNJJl/OmRVjbZo7ipoj9I4oIQ+yn4yQsB+mcLhW1cQt9vLhuFDAzz
ZlcXqL+aqnZdYKHHCHk6HvKjiGMMZvPfTLmNNzwr2nAE1MIwkyPhjnrT6lBgm7WN
acd5No6aaNNYaNrM0ixkz6kpwQSb9RcgerKiR1nmEojB/DO5wI/CsKfT5jfb3723
WhujlBKC/MDdcvdh3KAOddKxYd6vEihktR11dUsmm1wBzrE1SaAUNHTwqvpP2UYW
0zOicV+cKmfRov1N+o35QAMHCR7baDdf2Xe9s48Pj6wTSuEFPwaP1/A5pbxriXzf
C1pv61cEkXXLKo+M5z3PqhpIZ9PHeRNiu/BH/RJUCO2QDlvgUC6CR5qk45VVIUFv
in23DiDWlGa47cu84cGCBQ43ptylV66uKD2Rg0lpfclCxBUU62HZfEghGk8EEU7i
ncoh4WKW7sf66oy3ZSj+LtR9MQX6MUs/D3qq0KDhrq6H7Ey+cZ2ZZXj0kSeK3lGa
X/EAPzIelI6zlKIWr5qrEhzmi8S8G5AhrRFucf7gOp668eCv1b2Vb5QVkyDbDFhe
ZH13JoUlOR3s3DpVXAwJ6FbOdIkrE82cKYQRudkgqvPfhdIcFKHUOXUfb9LJoM9L
8EgwewXVi3rB3pk04KWSQ/4X/myv7EBMVdrOkU5i7647+EjfthnlHzfuhXxKzN+w
sLwgQdxIF3TDL/3850EZhHtFiGqOvh4xNu144r5mFGVaXVpiX8tDSqVEflSTraib
MTnNEqeYvsXTxeuOGHa2QVJNWO7LQhi9hjzNGpAh/o3296TEvNabgD477O0x8cz2
7Yc7fc+x0JRpBAkY7fWs7GmVSxuPjPpv8iVP7X1CI3e+g0Sa9vtnyiklIY9ovClL
e3UgETs+FwjBwwoio+uwdpwk3itETxEQwo2N2MD9GxT8FIYJJEeXzt5JncK2r2Ta
eXiLZfZeAZKMG78bdiXbKwmoDg9f0CjOZ7W7L87bvkVSALEIH9RNGhzBBzsrkaz6
1ZpIJ6cPT4te4uVO9Y/fh8sDHuJcWOqb/HbVokOFtXANPzlR8wA0e5ejsqMSdXxy
nfWKMtI5FwNN+EzXM+LzADyQVSzAS5PAnvmovCRI8zTstbPoFWg4XN5mrjpeR2JM
aOy6vlVUR90C3633jZbgIfTCgL7ql1VW4q5ckg+wO9RyOgUDuZoGPONMt9urbj4z
cSXs5uORFf9m75GKm88qCWrWbSpFYRJ7droWaFnWMeqa21uCd9fGboS9mnLSuSeA
/S4hJwSPAAplFLqhbXlZQ5hW85yqLbGGNlgxpMGZN+bbBZc+fVgE0IL6jMkwP7WX
0xkaUs9qyxD/qtlMFmp50+73ZgS2B/iuGDcAnZBoLU0U+1+kU52tvyhqgMkdy2W3
oAfM0RA5zlB/uLt7pqQ2giBnuXMEq3s5cjeFkGbHuZ7a1o3DnQgxGuVqgUyZ8dXE
Wxja6WFaw0deJJryG1giJmYY0EPS3bIGqc6E2USfzBoNG1e/yHt0PANVTNkjPtS1
Y/6p9pk87eAuC6n33u9FJ/C/4A4wqL5iCRWridp5qs9RxMcn06noB4qb9YT2nkqm
zn73WjIzt4Ubyhr3ektgOpxcdCYBo7/C1jG92KTVTfajB3TNQRqW8XnQdEqy3IlH
4OWM0A2dCUPtPXXcyQlNwhly+0/ZYTNo5l3RTxQu6ruzsCCA7Ir/XOeM9vU4cZAo
SKkPYaBOOp8VjR6SEyIRMiYxr5L/AmenP8CTBxKj1QnklVvh4C/eCL0QujryCfO8
ZGHEPOYK8aJyKmF8/bQz85cRk8MfQul3IG9oyoAHZ7AZM5QjQAml31Kc94InhG3H
YMVTLy2sCgttOYtZicjZX4P/wzeCLccmZF1CGTQ1WUOjQCg7sszgCiPlwJs7prqz
pJyBYgz+CzQM4dNHTTW2PlMyR6/YPcdBDf2FZx/J+0DLN3/8IPZtK+TCp64qgvzd
2Z3n1EPs6WQpUxruvRbPdYUC2BFfffey/HjEjp/2eYbYxlKDOfpKLpaYLh5N4ZxO
uzomXI35EEXBhQAOtEyasoxMM0JeYgmiWpYMNw6pz6nB3CAaethEKMzjVBy5k5Le
/ct5YL9RwulP0mG/PmIdHuNLyEvqFhX5N9o2LNaj0dyGcmbs4SiFPhFzS9s9tF2t
IkH1CQzwB8NhboPFkbZ30vo3+s+VDUPbKHJQJZj/d3asGOfo9bmopS6lCqN4sVkD
Gighf2cGqapRiMW0XLI61wl5oj5CQtFqlPhBERGWM9KgD3+uaG+yzLassVUnGR6T
SztQ0px4519wJ9Bud/ycQSdJ/bvHh5786k0jhyBLr4cv4lAshTpbS/JLR6/oCiZQ
ceBUrjlJ065ChJfJslmeZEKhvuzMsHb25wsjBW+kfFPAgRKjU9hLiv/j/cfpyNnn
yOOyNC3iQAmVSsN15QhfDDpjbVl/7FEwVJV3Uh+yeAJQP/53U/4E0nLcbge605r4
FWA/TdvaZohyM6NOkIZCs7DdNaON1ergS+1cVjuhMxYfuplhtMLGbzDljeQxBq/P
OoHJ9DV/mx+YkiIyWEI/WRK5m03Mn382QymsIl24MMY7Wa7L0m+QUxxmNCQCq/LL
oqUMayRLpYWwQrKx5sZbmCgVbhwIcyWs9rJeJdBUT5aBNTN/vGpVU8ml28ntRsdi
xleRleYWh6wqji5v5MiOuEjBPl10P9Yo1bd89v2rp9rh9P9Y0nw7hybnm0Dy4vMx
lohTfIiJtzIofe9o1N4UoZLLZzifPhYk+ipQhnknj/k083kgS7q83HZueA6lo0ID
lSlgVC2ipxJSQNKAaKMk0nNyEsb45VHtjnBSVzQO1kVkiYZZn3PW5UrH0h1k50oL
sOGPaWTNkvD0/9Bgppqiz+nQZ6TzqGHsq1573E6GRtXXBbm6aBe/975tDXrxbrkX
etfc7bGt7lLRcaF+Xv/sbhprEyhaERGNE0FCCRtVMkvibckQ5Jwa2pwdnK9A7nzp
V85P9vY4FYS9MGKdZ88H3hiBn4ZaS1JWybz5aAVcmOt7U57c+iuT7a9fwP9IsTd+
OsRWoeAWz1B0UG7Crw+luBuFOlZM03uZf11r2qoj0F8xgjoiB5hSAFsuuYUBE3n8
K1Sg558ApuNpk9SzpGzPxT9vGBIfuZR0rO9shDv7qzPooH1xGd0ibQnpiXT+saeJ
1mamM3hP6dn84TF0ctaPM69n+LBRStTnKkXUaG5vzYlZ8qcd95V0RLIpGmn5CBFr
bDNOAPIqHwPErI3H03NzVl71Xhb0pYH5wYDGvpPFohAKkNBTJP2ylP4Qhw/ixHba
XF6aXdwjxKWIH/gGnH7KBKygjUCTppWD14yvkAoejboCsud7R8GxGDJdZeIPqnMp
nBBh2TYQqoQJLFZvZFclBmSSVdJsC4awWJOIickmRP/UMRQA+USi60AyCSht951+
v1sqsptzSvXCoHt5b+3GzVCu/02HgjX+/Kl7NNJlcB5gpEcCnM49UPb4apb+86PP
sZ5fRERb5H4fpsg92hI0+KtWL++0xYL0qyge5pVCEd4uYHVlqb1PnjZ4xY/iMKgU
Q3MxZ9ZMtmxw9RZYD8MiuO15osm7qt/fTFVPuzLiD21AioMmXMapMBe8jQbinxcr
5no+MHVjCbs6UVuPUQ4LBlC1wvVrZEfk3xojGDiX4EFdsAGjUQtKfLBwhwz7Ad29
whXky6VrqpsQH8AdUAeWd/RJx0/xCxdZ1Ery7Y0QqYgcvtALa874Ht47Vlkt74JI
M/QUMFkzUDm1Hal3esDn2NXTvYLbVvyeSmM960SziWVsOArYE+Ce+Al5mIW4eSzD
csUZQMbp/JiGTDAvwV2wV8VHr6i1pMWywOQNL9zw3ce7cQMGaorBFCnTVBz5yAx9
eXdEXpDgtrF72Era4Vyq4knYal1aNt569oy7tAax3+ughxg7pjvC9W3jbgIbiDCW
H8GmNwyf7xVD7BTcWT1P1AaTohcvSFox3eVInxSCSL5ZJ/8TYetgmQ2lIt+GQujo
WnaIZurXpHukoujNEkJV31vs4gCEDOZ8VyhsTaaWW5Cpu0Rt3U4V1onCv5EQJQm0
CeM22pfci1j/Y80RypuXZuQX4snQZ5UL1F8sC3m2T81j593XmoEYWXzF3PM/ft1p
/rkBrXpUa3nIF+1yCZwDnNlAY8iAZpD/MkWpkBPgbJy+AZP2HB7fPW0DTKXqUc7U
E51IDw5ZBUPz7VqzYFECdnKtuHrNXksRnO1s8NBjbmhX5T60lRH3P4H0CVWe6w2o
IxfZ8vzz8lx9XOJ111ExpFas8v6YA7Jsabbvw80LQhqmZIaGPjDZLNvzMaSRMOQm
vLN3nlBtRwLdz+4pJOTnGDzwl0JkGdkZdmp+4RKXRtB9UZPQvtP3PvqFr9KaCMjA
Ylg0tjoOrRJQLxibc9fyTZKNnX9AVw9RoPjykTx2acVQCVnze/hxjixuAubuir4h
yDyi7q9V8Sawiw1263kr+8qJRwleim89CP2QD8RGFRcEfZjD27v09IBtgFU2ufeR
22i22jBtb5KnQ5huj6PWz36XSIhGc/TSl8AShGe/kyUyPRzZJ9PTYH2+8RPGYeXC
Hr1L2FMWivj1HGRiMYxTZDeBE3EQUFsycMeCsyFY3liByoDH8qLNuu0XE9gXZFBZ
S4bTzGZ5Wiyjykn7+DvBN8rILSf+IniRrUgTMIneiZjN8GkBfYLN8xpV+QpuF2eD
kjOgb/Kr3YUnULmcRCcYj3+as6iLLkhXWVwADWn9Q/9CuT0EYAhO8JsVyN35URA8
c+Wub0++qlCltEjXpnpPITZzrTZOyT3DhnreWWG2DSUJfpOZIqNFzvAQhRn1dr8j
8CwmJxvJnPm0ZXusArOuM3jO5xYiQtHKBh8yRsw+3dmKktfTrRYl+WGteO/tiog3
PimtISLoohJLiXnzDtx6EF8/iWTlxOFxd3dBnPxPrLN2k2WeSO7Saz5nrGc5cxHO
x30X78D61WCazJZtEGelq75O25hShog4Ae/cixuJugF+cUdb6j9777CJMVOoJXjL
EWDaHyOW4wsSSy0L1WyDu3rxjb0ybBW23+tcSHwn1rOU3WfMjGow4VbBk9KAfW0/
2559+jXL/CQy/mr/EV9aBSFus7+FnzVovaDAzBABiNYOwB6QYaFfZfoh4Ljlk4Cm
Il2+5Vuhw26+xrdDw12Ecl6cAvqkxOD/WzGD5kub24qcbpBZmFCmjH/25UOjZOOU
dg/9zIDdhtjfYiRz6q5r5MKCVqehi6NW6TMCxjVPtLCX0c4GimwqhqWxpFbuKDre
G/ha7tk4cVH+UoS/CyJkY4ZAydWopBLAlJlzr2/GjUkJdVZe1iDBTm0GMni1Rv6C
/itb3VytuQGIbhSFLjUq8OvJl6bqOLmo/6+kK/ii/XgXnQTXZMK0hsp86hoxShpI
+Gqf/MWis64g+uy486OAcF5KDZjzNvgrDOGjZXibJSev0u/p7+YlG7rigEV9coCp
eL9mHChHsnH5wogUn8GUiQyRVIjUaXdtHzxD2rkmwSK1/nib91YUzhtIsrZ1BkDw
2/4eSengGZnuVyDOInUSn3J7Av9Sh1a1TA9grsVnkA4iWQQn3iL0PeFoVLkmon4s
OTPOPFUyIHupYKemuNCT/Vcqgxw5uyzqUFLo3bTVq4nBHq5fTTeg6lT5eUsPoSEP
nOA0cR7T4G8rdQVZ0E9mXfCq1w6KbUxN1jc6yqsD42Wlrd8e3WdgpXMU9Axeq0tC
jJyoTuX52T/ik6F+9QJJ1LKm6unRz02Lqg2v/hFtyKjhvzVMMVENoyjr8Z/AIUPq
TGKUxMBn0UapZ+nP537kZ9JnnZ9Y2jhJW/nUTBEjKqk+6WF0KwwhShjz1a8Ittw8
JdufQOswpmUzgfOEhgfkH/Ni1ErZLv6sRDzfBMXP/dm8HZXwJokS8tK4vRLb/m1e
9YN2tTujXIzZIiU/u2KqkeyOVDftYVYoTOlMotLp/qvuAm8NB8cTErGNKKg1rFa3
50Me3rd4im/9uo6ji5RKFAqHCw8TV6Qc+HbYGwTtTPs/RtF1wWULrFaBA+JNbIwh
f/zrI6BA4WHd2u3LuAxCHWcoQ3sJHZJx9mqry+6J2vc0raV+fgJh/XCKL7IvqSMs
In6b5yVObN1a/m6pU9/yX+4EB1NDx2cjchtDn6MUtfDMH22D+UKTykEEeD3NgAo+
NmqqhhdUBvQfI5Lm5sSbTlMGJWsN7Y5Q9zG9AOT/C8LvfqE0GoYKXUwmxmIbPQnp
G7tivj7GW24oN2MsttqQ80XVNHmn1Hoj5ThXa14wrF7yFHF14KToGpnRMEUDDsDi
6BpSxE4Ce/l4vTFvcjw6Fz72r06QiOtLDhf5zybn7WocAP1z7oC6y+EiGAQXGtck
u57SWQe5wEtibktAffVG4CFhQ1ZArzCGS2TGhJ0VOz3ki4U++/xEKJ6XpUQsRwB7
CAu7FcmA0qUWP62ouRgI4qoN5fblNfmN9V7c42wAagD38ZMtXRT8oKfNwdKUukeZ
G0NlyuQSiVMehB6QSz5IEjfRRq65V6Ps82lxcZCMr9k5yBKvEq3gg+4/gNsdfxRG
Bl4g+/LXTu0BkUgo9mJC5aIWMNELtQsEWGoG+NBXbHSNQCh4+lkqwLxLkl7oRHAX
pbSTDr2kubwdzDH4prQhVIRGxjRiHY8FbKgvXqMHxR16ASsPTuSzTZ11+G31WXom
0+wvProcBPsdbhhonQmTiOIMQkRCkmCOKDvziY4VocCuOuhGlGfSu7WaMMAI8158
Gx8ELaa9R8ZZHNMm1oevBJGqcMZpgRSLf8Pwiy5UejoYlEek39cVJ5hp7FUVRWyh
9z3O1SHJYeu9FjIhxU4lk4GMF4JFoIzVqlL98Ckgp82QT6xcYe7YGOKOzfN0ACmQ
PH4i/rlkQseiesfeIyM9C/NvP0agNtRg0rMdHx+NX43EJwUo1TKCuyx8XJBOMYvu
lo4wyU+92Xddt3PyvkMw3Xv+/gkyAn5e5XATWJd9mioTMmaULq+Ci64QwfGygprQ
bz3AikneAvQOMxirQFOvHfDCFeV3jnY5u5kLlIIHL2FKamuNj9G691smCuvV7kD3
qtDPE26/+eZcHhOLeiyn7lM/pGcmGTUfbEGjQPmhd79FTqxFe86to2gQJAnJfLXC
P4okVMXdr6gAhbmkuQLVHkHUOvIHUMlBBrYHjCCH5TnMd3X0Stpi8xqJeoWD4cCV
mPcIRqbdA2c+An00IkpHSXAL2l3SGl/BzavvAdUoAq8XM85a48IouSXLOYZoHH8H
OQKIqiAXF27gbzOhWFXcCMb8pYQoKCqNSZprW9r4PMtnqYnm7sPH23453VVetQEt
FDnCkRu8zmmGzqtzfAD7eWm+EVl2G79ycEveQT+D58sAlYZr3WK2xihkQScMZdBd
dXZla3bgkyh6VbdVR8qA5YFhgycgJKN7/F7pvhxhYejstJQh2PrAtT2LYAFbPTLD
RbGpf8XiXHgLnwzc4GP78/nLQAMb2rcNIpC4FOX9YfmbSvS1cjzD36iQgvXvqFOx
vBqXnoJN6bTpiJoR+Tf36aqZLifVteXTpNso5pRJNpT7Jo262Q5dXDAkx5uvNkeF
sCvYrEzGTZZzdOzpsqAOIPYy6u7uhaZw4pjkweu16+ICms369XZ41KBno1NJxe3h
u1EUAf3OVyUwGFm3pqZPja+rRd9jWHQ4yw88IEFw7fD+CylRdNqZv3j1WedLdmNV
osHOvxdk74BOGqN9n8kmLuQ9hbIo8UtyjU/HemguA11yuhX1j+261465Z8DLmkXl
YjrkihoNA4+Ayu+nGNyZOYkrM1y31VyzM0cBWB1DfHFyZqbLzgwhf7OJbfjHECja
mxkBGOHCmsddFUeRBUAHNri+ZHSbl3KQcuXcM+ulHTaL4ynrEOwJNNao3mj5sUUh
npiXa+K0G/OjPV2RkaLa9HguS9HY1d3S9e8Z5QUcl4qAZnSExB+p8sTXRFJrVg45
WihoH2Za8B1iHUgCx5+ao1DLa3taIRz1tUineipooczl3q46Ct81rXD9AAcHvV7/
HFoQ+OeU58KD1Soc8YZl3cspOmd1ul2tMx443CEz7YZcOM+vxPTRdCDa5F0eykx5
mxVdxfdD0FjV5JMJqu/0CXriJgwBZOK7O7/nb1iHHbKNlILhuIR8HmH9IEtHAB7D
KzXlR7nXCxILeydoHG27PYsICIBbRcty28gpKKsJt+jy9pg1moOIXk+Nj3v+TBob
rjcmGP98o0EBYD+sa0YMzI9BZ7T9tL0l3LF9FiJV2gWhI9F0oVbHamq2fwTUnNqU
LkMd8iLnOiMS726kafTrh0spUBxS6QhMOkQ2vV7Pc3jh39tp4zw+WeJ+DcPPKNEF
9N2CLXsX1SrngadiMX/vfUaQEVNncOI26svJVDGlNGFS/bDoEjoY03lfa8OA9Usy
hKpGthfLL3Mhnk2H+PgaT9brZzCHlX8A1eN74ovxhpQvl9qZ58kZYDMfFAV0+j8D
/dfTDHQISH9/ctPFNH3KbzmsVnIifXQqQkCh/lyLKM8k8sgcp+8RV/PbPGSjSVM6
Pf7LFJ5oRekpZLfM8j2gOxJsO7LyoA6d+DrNdaI0sFysfkXix+Pz89Tc8Qve55Jr
LFLP2bH/5LqRABnYgDGcMEZZGmDM5OLfvqb+75FYh9oXbuA8DucC3KXGaRaO8EOg
XcJlNgzzzilLJRv00mbKXzpDK/MyMk7arQwpKi2lfzZMgkrARLP+cvReOUMLpR7W
7OV9ugmY+EqliDx69oZUx6e/13tzwgn6oqfvGUSyuvlfBrMGxm0SJvHgSikUJ6m9
bI3P3UaTuCFVWf5z8NKBiP7IhpwKPbLhgM9XzX4YSSobx5YHiUavP/Zlm7q4E05E
Y5rLnhs/TdXztuZXyD4Khmd33yyQbqMdskGrdZS5q74Qup4+f4HZ9lmkeq3W2Yhr
PNPc+01ZEdZk32s7ZNQgeOOHNbvgP4wZse+4UhvIBEL5fz4DnJj/UsYHmpzBYtf0
t02jo04RrysvytOdSO5/9hwUqYihpNkg1yQVIjJJoKZxTw8xJu3LfofBYj3IM6h4
6ZeiMqMeB7z9UJiJfXR/353nQ4hCBYNU4ky62cuE/6SBJVtUMWa0rHule9WX+/97
RnmqiEvnWueXt+iAAeUzxf1ncMkqqI600/t1RRYfYuWGWqMy1qzGbEzmL+YjsKbd
FMZdGU2UcDD0e43PqyNer7ZiBGDk0hoDqlxvb2FHOLi6PgWQDpV2Mt7kTiblFvSh
UKSBYHa2VzhWfzedx0Wxem+D8EggzWlE4xA9DvfFYeNwzdhvgxtvIAturP5lCCqm
QvRvohy53lBXyf588JShN9z3JQmHha3nYDI4eh1oClElhcmZozmD4lKPUMzmTS2s
QgHHc5RhktN12c5cXoq/mr5W3cmHsNtZ1WXFXw1iY1+PFV+izTCg0h6AhcUR5TMP
OSyA1QheXsq1ttUs/h+HECMwjA8kGqH92tiX8dUUuCyInOSjLPtbF/7Q/1qVQehr
jd4DVJqDQY5mrAhE5YL9KT6iyBuly31EnDtYrrkYXVP0VPjdjm1Mo493ZfK3cw6g
7DztuurN4ErULfzYgACwoFNfFJnCamopPQp4nRgpK2El7erM54mm9a/29nZbXybz
hb+Cc/KvlilhEQPurf8XPASY1YBvRhylPRmfUk1jyackOAZL8uYOIoFXLQJCyASy
q9n4zjOqF+b7UEhzxjFQDTyRcg/WA+0JRBxzT8IMjQEi0WcCkILP6B1/YIyrCM7d
pUbkq8klsKKoIqV9TUTMhD5ZmcxPr2I8KIwOeFGCNQu2hrI9LsCh3/MFDcZ5RaZ8
Pz0zdTjJiNp7/B5bu/UXfNmQTdHqKkUOo4v4poylXYqR8A637Q+Jwnlo1wWGpE1S
lqLqHLfHj0NUhuLMLjCDxI2URRKHwRyueIQR2f1AuaDqkE5twoR/MPxFvK7D2/NE
agCodcE3Fc0ydTMJSwu+tp2QVVZgwCLH05zDK4BxzyECnl7I1MQRnft0DKWLgF4y
Kl4Mdht3c7YXr1g8juWcFgmtXFEG+hgj94QFcocnkZSRryq7OefD2Q4QNzxt04im
+sntuZpyUWAo/2s0Mjh7BqAYSXyr88SlOtxFVmJ4ZYGijmhPIY0SN2h9YGONUG0K
ZZ3GsMsbgCis7l77JQkzL7ldd/AaazcY1OAutyUxTi2sxZjJavTyzC+HFWNcL7Ls
utpB0FaeDb0Zp5OCN1OuCF6g/bZ7RLjLxOwcPRNVJSpdQ9b4NvDi3sWi83WDpYAV
opJoE9IKzeKBTIiShK5fDg/hMm4PdrJu8xJ1zXUzp1VwqVo2s94piY0+x15P1bmM
vJvbKXmgV2tlwCnf89wLstcWgTOlr6zx3Y/p8ON2g77YXbZSVcuuIkz8NER7O5L0
npaO2ly84pjXzkzwRoAWasU39Zu8PDLUdgjHw4gGcd2cFPY6uHn9nwNuFl8Ba6dv
O90C8Dc9XGnux4ijAP31AXgrnLZmunx3JgP7jOTs3l31im4yBm2at4n5HduCZi24
UZ++bwXIxTSpjvfN1ude35UAohi3XodAYegGQXnFiw6pCToaKkA4++lRjPxoLTta
d4jIKiRTsYSW7pmZCvpJzFgfmV2tl5pUjqiqQG32T5+rcNBhPRskVbtC181NZxgA
+8SQ1vjfFrEUM73s+iI4qCSnkx+a9rpbxJMkHK4x9+957Y048/ydhAS5BbICEorU
YWA24/OkCmWOY8EZ7E7tBwmqZM627vvp/LSzEhamh4nioDf4jO85xEyzc6lNT+M5
9TnMkr8jrl3IFMwlNqWRladeINSfeWocUefCDnnnjSFEvvasHRcGmbrNE9wAgiLP
aH7ZHNCaGmfbq3QBNKCrU9pu8I2eM+NuxMNiMHX0RLnUULri/RJf7f6+p4KQQr3o
0KjfZwqsxz/GZbRyzIa2DkN2Ji5h2qhwzSIeVvE7+Y7Xvbz/p/oo8weLyVS0TOx0
r+gR8wuKLjUpu94qO4++2054FS0uxbugpe9fJckFQscfCfsMkt+Frtr+mNWhnw3H
5F1kPaSLeQuZAIIUQ+xBhwYL8Hm7qO1N6yxbete8v8lH1gzmdCTmW7EwPDQlxHmM
PLDvH9l0wz1HlL0xP6Wlipc2rbpz1V4Gc4jsCRDRRmutTcir/5WtQ8VNGK/Y5YNe
vvfSVczqtddZ4PxE6mPFdaNKtiLm2SWzH+7a7shlXwq+twyUsLO9EqsO5wN90xDO
sy6prKx9YrZxmdEDcxHEKMA+FJyf9FigOn85qVzPAYJVt6OshsgyApYGQGRBbSlv
wz/9WSE3gCym8wiE7xrsq7OXQhuoH83Wri9sY5ViBH4XMqgTcn5Z0HPeQr/fqkwT
pBqEEd2dq1iIScUsQititcdkxy6t1hnpu/Cc8nh+wFOeZYH54mZpKNKXY/NsAroa
GZJj3AmW/nryruq8a4P64DaKb/tKFSH2KIManhkdFLvnVhiPDGCCTD0Awh/EYWcy
pHAJHXAhqw2ilJjXls5QwVESBXHoAupTsyZUCsfC9wL8yM1FJwcxTLMO1D4MVuNH
0ey/CEpZ8dsnZ6ymVrtODv4DTffQ7j8Sg5QPSTafPBMeb+T6pDxefYNaNTUSz734
jY40WEr/ODQeFLWdKk8eG+Z4W7mPHvtaKdGYJD+WJQKr+3H7uu4Ml0TIrRTaT1we
W25GOmdVFu7U5ms8HpME0GDN2dQanK7tsAUE9EC9zEAwIDtXW4ggpf8tbfMzdqNx
lPC7qdNqIJY3jzEpa9iA2q05vkXTy8AJoVZ8f5TFIbSO625rX0dqlCl0rpOXGdwu
T6g9OLkk71O5Y/Spj5Yg6MWQ8T29aEdDnm8JRMNzIuw7ZkchT5N888O1zpXs2ohV
ySZwYGmuL1CvmMTUjwSYl5xssT9wzre1I2xe6OIHIGNXtG35vWBikznFQme0yLV3
8S9E8xQA9AYhHHxuGsPTCV3uq3EKhk718Lhs1MqUmc+3YN7W86c76cYYW+z7lP7A
G0ibtwcVdLZOz05ej5J37CEFVa0RrKyvbGOh8dDW2c9juhLHL9PNafMg/AAyAgIn
eITF11FBO0mnyaozf2GzZodXUCXklAPK8wmbKyImpX3HG3jbHGNqdSe43msh3Fq3
+Omw3/wBFZ+AH7YGZKNix76OrSgDkvL4Fc+WIwYMfmfiuD9uRSsoimZOmij1df+M
YQ9SR3G/VQTHh7rMovgFjNzba02dIYvMouHSFGmn96F25nH7oNPmrmEa7hM5IZnm
Ya4F5YLrb9PHafgR2dSOHqhRRHLjImCsV0/fJ+4LlxAZwK9E3XBudtmiwqLaPv7R
xAOyESwo//ovFfy0qzIW85PbJwnwoJNpHC2xUHp0RvwL6WaGXRjBSycQAwocmyi0
x8b44wkBL7Gq9ScZGEuPTPd7PJ3wB/OvcdweMIw5hVQtIcjFeWf7Ygi9AK5YGDls
xy0I05jbLjePjd8wccQu9a3C5yOLmEYxCMxdySA4Bc+YH0O5t5Ss3flpX5ilxL4u
J0l72R9+3Pxc45t1UMIdKFea0eIAoTOME8Kaqoy/vTT1NSq2RS3JWI7oPSFbn4ph
bGdHA0JUhJshLUE5IN0fvOjoANk8dyPQgcj0QGrapXPC2U5fcE1FDrXWA6GYOgfb
fsv36ZbJ8co9C6oQJpAl7ZkvXN/lrE+kP7kQqs4jNL8hSu1MC0OfJviQSFCSIEVR
azzQAjla+wyWzmjBkx9RB5QUcWMY1VjEGPj1UunkuoH3FbYSovPaQ6043g8YqRsW
TIHfXMZV9P1Ky3J+aKOap6Uj9RH1i/tJSF36xg2QPANHhzYC4ZWFd70vs+qcstpg
YaC7gqVeWD7mtUuJIUxwYfJsjkxlALVtvgxmzIxSN5mq0ErIwZw2zw5fmeKwGTEp
gcalsEl4fXZ2JG5KuCrwJ5VKUegbVGb9DG3/XfrmN+VPfSJBh+3lROA2CWsUyHnv
ak7EsithK1lkMUGTvLm8Fj9OzXzMND0yD79zLqTSfDnShKjZqXa4G+Rujd7pFCsU
LxcdXs346rJsjmM3AzLY48tl3xALwRR+NYDMCe1UHqcl3RAEEIAVXtvvhB3ylV5x
xYVgu2ycqRubH8zdccJyexmcvMTqmNAW/JUEqzd4HLaY2csZql6HG2NU3cPST0aJ
khTQ+qnCCbzVY0kclv4X1fe21E1CutN7C92qo8GV2ICSEKckVsLv77u9zYAkdQue
dPlqAdzBV9QW/ZgIDBza1YSgWrsDXSduonjWgzYpINupZwpYR6FivDJYkVWl5D4t
FhiYIYIwBFFFFH1n+JGOUJirDGZumdBhWLFo6RvWHIHTqTi0aJjbipHNy62PuIXG
Ilcgw7WDrcXPLjmm5rMJYhYQlAr2V9o1d1RvdKUPyjmf4OaQ+bhMtuuK/fCEsBjz
rGFKADPDEdM7EygYjU/PqH6P7Ly2ziIWScAXmWB2KRhhV5J4AtvX7ga/nhljAM+l
kHawgJ+Q/0YzKqsBjV8SFYN7fO6EaIDwhTBlt7r3hOXCHhjAA1bGotIE6hLqvi3r
EVkI6b4ziH0bzv/Iz6Xj1Y2lK/CcEUMwGlJ46+99A3SOGaM1bGU+L9SmqPA8owmu
MzbxQ0+yIKRtQPkjXtY7qOOtDZCnJnAEJRVnt728HMlWFmwo1kBC/IZEuCVB40O8
pcbiMMSJJyfXje2ZS6owVcKqJHMEYxMU8f1SHtIcO1bzL9qXoBmhqXAOzrGn2JIV
AXp777GOZLWlYFNDO4VRqyhrsrfu+OjMaICRKpMxS41QuWNNEt1zM9NnEwI85ybc
n32WN4c29AEB8S96D0iWE519UtNw7MQ3zSjPOqrqV/FU1OhCXgvzObGhuE2mG4tD
LFTbJEzwaHUS4HACD3Bvtgbj2LMHUOIpQM3csavx9KvErThq/O/WZsepz06d9Edm
Uy9o690iUfrZ0nqH0euNE0ibt99gw4dtz32E+Ec9GdwgU3HtpKZ64yu7jxIPzFF/
2k5z2Ze91ZCjrnY46C5BTTew6rNqrLHVQiATzZWHX2QgjdLaJL62SM53ntTtmsbu
OJE0n8D3+u+AZFW/ixHxaGKV5vE2XgZxqAxaZP5aerqP55vKFzU261vznsoqwlKx
U5Gf6Vd+RkX3yC+60p4khNJL2AbWSraZSDMpeT+SGxFKnh9l5CLKzHqsZBeTM9ee
u/QrwD+vfuwupfnIOdX0jUz4IWCIRGbaf6/6jGHUgMAJ8YHDrQQJCAHKFl6nInOY
nFjQMiBPxwiRsajiCiS+3uaPlZMxgZd8VZAEgH9tN/6I6NrMmGMZbG7NDOgjXP5Z
TzdEudiNjoDDq7JqRNjPysjeG3DVzlodi6dij/p5iw2hqeawIULODC3rm6Hy6c8P
wDlMFQDeVduof2kGbDvDWuP1dIrEeQAmKOlJpudHIqL6UKkb1RBWtnm6Ap53FRzq
4Rq65FqIoNMcc5vxfHplfxC+4TPnug+rDZPctPwNW26cSqRa/rGZ3FE8gFt51l2T
m96Y4qkWDG33nSswJ98tajjsoUFiKhWK4/R13LW44Y4kf/zAbwm3Wt1DFQREm0pX
9N2XbJgGveOUWd3VeTa2M+bXqpZmlU/naeyLIj5uJrc4/0i160T8qi0Tnqj3QKjK
NdDOT2VoF4Nzye/XBXpuL8+F2F/TtlP1G0Jyifxd8tF4OfdNNWdlCEEa4G0Q/Rem
iY7O+kMAlACdO8tk85UWLlQEeyAG5EkhiMAVFiBFTi4+rfRrT7dq2pspS0FCJc9J
zNuG7Wy+zw544GhNitxQLOUiQu2dMcuX7N8A/gwJnwXD99R7LCJ08GiaTfLd2Zky
DralZP5AxYXh5Uivb3pdPnVmxJfqWJIrsnw1vC4z7KxRTH381gxXfqrLgeI0eP73
CGXQnsGfYAVf3oYdxBhZz70UZtZd7ZEXDauJEnEVFc74nymvSYY1SCRcLBqrfdDj
GntehBSf3gp8ABYOY8Hjaz1Le99Kmnbx/sy5E9WzOyxOI7BeOhykUDy0ebuy5Qqx
84Y6nNAHClrKXos0XUm0Vay0WjI9bhovO06wf0fzHnP7XVluTihekUksl1lJOsK6
Lrc/D2u3PZl4OWHVa//nYhAyK+FnwgKxC/Z3dGHKyslPjC4AXkANinK7vv/a4A6N
oKBc5FC3OwtVmxEajtOq3JL1uxjDWkJiGKOjr2C6bm2bMEUVY3Ef8VhHfb07oosj
XWs0P1+zJxY0IrQ2+MMnq/puTf5HPKx91nTFB/qOuV/0hVIGdMFAV97kSEUIWeOe
V8TgWOyYLcJXgVr8lHtAo3N0qYI6B5HZ8F3YJcorm3NTx+lTloRW3EqZZ8FMVUcs
OtF7n+z8wFfGNu++49DYGaFf1y04/2wzy9mGV/XhxpwXdCK51HBCiZljfjRN0396
5VCp6/Aezukw/VZocM0rud0BENB/J41bRFUWjaaTCtXy2iQIAbitjUE2xDmeTVmN
a41pE+hd0VZBmxRoFYy9b/KO/1wQUET1xUeYJ2uJAWSvTs9UeMJLJEElGaOAqRUW
8jSYNsTXgnLZmF8QZbd+LDSwZfwhF7PoVSs1L78zmQ9pQArd1NrchHeSdyKTW8KC
+p123gvfQ4XcdSSqOTgobnz024B2op9PzwFD9q01GaAhqFBUKvvW7FYj5aJQI9kI
X6qicux8rItDPxsteN8tX2hK3zAu9s5csWSOrphSbVFLTA63Q5vKFeHhHKGHiTqc
gME3jya2pxpVHwhJahHdcNoultilQmXFK0FL6JHiRQAYJvRBPTuosIx17RmVtcwF
0hqf7N5ZLRHLqL+/hvmoBJfin+XJAJMYr8lTBUXtcy1U5TElEi5nnyGcqx5s9DOl
HUi/JPliyvjPaF/pgiB+48Z+aP5LyehUOf9/0FpITpfgCV4vUdzcuBkOlpyhwhdf
+5WY3JO1DD7hVpUmF/8esQ4FkTfDeU8VPhYL3J0b/5G9rd5r4E1CryaXQZcTwgcj
9vCosE/w5AoO+nXS2APDwE3jp0KW40tqDj+Fh1bvud6KhsaYy3TfAPZCxTTBnGma
BAhrFOPLWqLn+hhWrS7jOwxZMfE+tIWvCzKhvfb8VETpgtoO5n7w6aJ7ClBr0c/k
Y1YxR60dxhyKAQPUMykLJzTQy7N9tXVqwHKtkpvgp21f8NR4otxKZQ+L7qHyBJhW
xySD9XuEDXS8S6oCJGuUlhYYS7Xw36qszqzPzK3e64qZhatDI1wGVeWj289I9yjH
BqtX+BanhxkZXsBJQ3SIzoXW1oUMDGBqmChfFmlxDBjR8HAErs9+Ylwi+xUMvs6W
d5IMzmWU9vINZN+C64KL+mqMprTy7Kf1762cwpQEfd7I0iJp59giDv6yxotQWVI4
jcGNYPcKi7namo3jHefh+K1RsC69Uj3nN+76x3elwMIgzxEvMODCcohyeLNDq6up
VgWDmvYz53omq2I1Spgzp4Ar+9Olp+XE+jdubxobiseWiB/j5M63lgE79ZW8YsPt
Y/Js/cjbp/fOW00/TZyze6opHDBuxs3NjFv2nO8aaujfXJGMI5xo2/5l0dV8j1nS
5apbp90SVIWouCZ2TT+vefQARxRT99dDWP5M5b3NtfcaCTG/EFPuL/XlUgMbGc5i
ChTlTDSKRhOO8Y9o3z1fzeQgmu+mXTu6L4b2apqdLQQ9ROwFCdnzKYwpGEzMS7TA
pICiO3Fw3tPksOlP74TNSwdi3JCuiGXaJH2EpihidImuXlTyec8sAdmsUTAMBHI4
zvseRnOzVHiP9pvDrJ3Jexup20jvoWPTS84vXPPsPP9dqEp0wJR29pO59wbWcMXI
tPSL8fTBYkofeMSk76F1LcbwhrJ7huE+FBYKdFZ/uUB0cS/5vNmgA9UgnifmvKxJ
JTOsk9iYVkzQrE4UwGQxsdqAgrdn/bTY46Uh8cHhzdo+nU6LWKqm/0J60Q74f9Uo
SYqyMrSwZ1AZ73w59+sFpzvkPQLK3JoZr0gGmP6hm1vACm3jULayIN0QxXQ5W4M3
7noOxg4qJmfOj8TWEy16G5wWuadhZ8OMBz19tR5neYyM/ysdbIAOOW9ahSi4xRQz
nExnlfBN6cq7Jc97IKTcvt3x0x2zE8Yr8djUTkZy6hjlSFBwhTXPy3QhCG7afuAq
ctkHjf2IaU8alkf0VI/RyHvNvvDyBzBqNziRpCfe9gHztPg5r4yxMgug3SapPkOp
OBNCr/Piw1RgvTTsyFTUDoQcFBDaSpHD5r6pebClvFcrSjAAp3oNQ7Q8B4AZKnXu
2aBndqeN6TgiLcDh8Dv7jgcgNIAZpSR+V6C01YrImGekNvpew3eervbwuOeVpm9h
lykFjUwSeAChsgAiz0jEtJDKxDDtTBpvmzSZKGwsLX6MQ4AZz4pd2wkU3l4Pn1Qr
+D2JAb/7u8UclioneMCmts6SN0VxARMTywnbvK5lgSYTPv4mSN2wzrnxQoALLkPA
V/DUg8r2utu+AVQFd0WXRrNb1RCdCHSx92n3J5FRXfaxzMIyp9p9JUfFQWirl5tX
2irQXl2QQsK3w60TD1e4NGECI/+HXfVJh+V64+oHdpzJSDjPmGsQg/4Ghy6Ct5bv
F1Jn/c8g6QspUa3t1SQjvE4MZEl4Uc4GcGAB8IONc6TE1JuofITrBxHNBF9QXBNA
Ye0nwiO5L9qaCrH01IkAqG4KXmVcxvmhT3qpcXIys8jXfgHWpBG5rhCi+bF/6SoK
9JfPaiHlfOXB/lYrTuPk7qqoGMyq9RIp7V4fbigpWJJd06FyQdnXCJCGgs+IO/i/
4XQiikzACTKmgoUX5luxpfyESAjvDb3apv00svjhjw12vL0P7vCbzHWFOruLmHnP
hIrDrntfyrDHQGTWlKD/WbdPswXupRxpOUk/a6IzYf5mMzrVUqU6Nxzv9nC8YS6x
b9n992wFWViFlAn/fxGsMIzbAxWk71/sJkORtvqB2OWIb/OkmWjOkqg55C7zGe+K
Px3IFyS+Nvboc+8LzcBF9f1qWefIIykYjEjWGQdB6tKFg7AxxTptm4UMo60wdFDQ
dCpvXGsffzgA4z5kIl1r4DpxfCj+HVTa3IMNlQtGfB1CqRthnMpp+HiNFI/wQI85
pfpvIZuVk6wMt5q0BS/NXaiwPrlKrFplyw0/HDryHSEZvj6jebI0Yu15BUoxHXZN
4kJmpC+HGOnUPOExndwyNdwZdHBjTVC1iPUVU6B7e074QGCNnkvdIBoKkJiYNvOJ
OpEDcw3/rpntW+AsMb/FXsKYl3MAMKGx8Ty90K4dDpxASfamfeKrULH09WweAd3/
goQMLPWkft+fuHCA4CUu7EzBwIPEPZ4T5tyh+CyEXTBV4/7wiLptL1AXdbUTe0GQ
DVhj4WkdNWOBumGfzZV1Vn+/r/Ve0SbsH2hBfdjHSDf1ONjImsI50ruc3fx3XLBw
0YUTc62yUYB/kTo6YroSvOmeegpBA2O8TlWR2OuItB4eWCuAaja+aYomlZGFo/t2
gvYk2GD7C1wFov9+C0Os8CBeXpIJW1oeyqRoF3oO+yyhhQhP0CtRnNs7lfkMYxVz
L5fL3ndNFvAvNk78wvktHbPUVRZHqvmnOmGDlhwTWggwU9B9XkyzHqWYnObzFc2P
rxPPYD1uR9g0AGh7g2f8S+KsHreUI4AFh+vjJt3vVKCStkFPhdTJjcRARvOZ7+Fj
riWYF1myFH10P8yLXEBOg3/2pRDFQMbwqF61x7dlvg17LtTVB8oN9KxCPDnmIkJA
C9ba8qnEZD4VTJQk6yBxZ9dndgsjL9IGdDCWsN5Uo8iQlnlORT0bJZWOvj0SfA0H
26l4Yu/FLd9r/MqCcBpN/6WizXHeUNNXzc4/YHFyiZDx+sdMypXt94MY8KWkBFT5
Tf7aktMORXfefuSjKfKErn7du7QiG5uyoi3cIMqf8ADlpH+r7rP8RZc78DHKxEe3
JsyMcP2JPqpNJNnrPoqqwtULyghyNFIsYR4o39V3TZLpr8pDSiEy9eamQGBUAuEX
TJI80k9UVgZSIeGXRXPnGcsWmmjQiqp3gJYoQcbWt+uu1ysa7U4dDeprT+V7RaMl
k8YoIy+RbtYUxVIVM4+PLVxP6zCo1ngHVO+PqVCHeG/wuaQzyO61s6LVMuTmEU0R
XmoCINVxCNJauHBugR9u4t99PdNca6jwZtBOv9NU7KFxuUYD5uuit/6wCZuIckc7
N6a1ZJiiS3mY0U3ettD1bNT6T1VHBEc/fG1Wf1od7zoR+BO0hVzA8NIZ1NVy8tmb
+hlDjLdZDrj5/hAus3v5p3BIFrVl/T59PH9GeVsCZRAd2ksXQFuKwMCbXjEW6I1c
gNlKOiVeW9CZJITW7cD9lhZY42i10DaE1U1ThnCax8T66rnr6vBGuvF1ogHn/+zP
EQmo5QhIVxjTrbqU7H3CnecRnurYmSHn8N/TVQ/mYjQrR4Fgd+gzf7g2qcvwdT6U
yOYL43uQ0U047tz4LmXv+sPQ3LF1rsEh4NFVxFs/hjd0abFKJ117DBi/0RE0XhME
1aGH31N0xQX0A7O3Z6dkv4AaeA3N5iwUqEnlRRxqH1E9CWpo9LrkM7F5OGrOqr/v
gvSPvMGEfJAnr9m9rlz6jAEZ2fSNOTP8qkGeICdPhI7qYjEfrniz0Mk99mc9Bo60
dwj6uQvs+BRxQEM+jqHQROzru4/K4ng6GgLXOQ9fkD5zlO8nO4MvCFk1feajBl2f
I56kMiGZSPmbDUAH6gJlSJM3WrexytXst31wsMXnZE5pLleUNszOjH1q/CHBCvoq
54dyHo+/B4nSCm8ft29It4Wptg9M3AGx5Yns3tSqbXCwpmGDfOP4vpLavUYgbY0q
jdmAgBbW/kDwG53CNyG0TyCu+8mYHC0M2+taqKBeiSW2c3qpkhb71H+A+7SbFfw+
rXaQASgUAB8YPaTJI71D+WXb69yCRRk2YJAjgGEohSnT8mLTxUCs4XRt7TPgWhjP
F2paecJU0fafRWNHzjcVxfFJXFNMwf4hGVQcD7hCkxYmBlVdihMii7FaVVGcYAmF
KKG5Rc9OjbZZGBc5QGNSZP/kM79y5Z+DAkYdAiXk/WqbnfVsTH1nrwtUXl8jLFVY
gMbjJVdoP/b77R2fxqZdV4jfus1GG3Aoj2qephrWnP8pdZwoJp5tOrH1ucms+TiH
AFNI0GtWZiOBC3Rb58SDJx+N4q3MpZ5dTxGhPZY+Li9qgVAGpbYiUgxBnrJKsBHF
PL1EM5B1TDc2hiNmV55tCtaNKNd+QLbxpZuNmypM7eMcZ0TQPIjUxO1eNy5BE5mL
3JaJo/Qh+qLlJisucgjULkDmBhFXo/KjoWWht58Y/PRUXDAfI6/WeJ+HGbc3erb4
O5fNS4Ffz1y7C0oqw9ljXD2yRSv4E6eMcmariEBi1ufqsSJI9maeRnZDyiTuYqvw
Cngsqd2MxEmvbMm6Ph6HBZ2cCiDE5YP9RH5fCjSliUeIjZuT1vs0USQ1dryqKwkP
/yVM4ImIqXT9gUPdoAtFDPWykXlNkyo9RXqY5bhSUqh13ny/pH3u2e8zCVHDf3rq
qjC5rirea4nJiM4dcsIGozVNJLF7Vci2F8F83wXZuESC5wBTozS4VgKEdDZe0KAW
SufyP2WJD2LEyhVGVOHcU/zyd+G9PwnTiO4CpV78ZOj/pBlAe4lRBYaRgog6732w
3shyJLES8QCpTRYi+eu9ZftHNWi2tWKR/3BNSIuDD/PBv7aD9kzz1LOpmcC5UASr
SddVJFQvtxahVqFmXEN3Y39Q+q0Ld/I9X49mLk5+g/L6qnV37aOdLST2lGa7uXiC
vMZbS93xGt7yKXzGjxq0W9A97d8HLbOzCU5Fg0ZZ1nfYDAUDNaMyIo9GHaCG6YS4
tou0OJFeJJtt955eHRGGI+THrrijkE61jlbXPlQWkJoy7dRigjE09Tle3eeWWSnj
lRSolaV4C5rSk8FzTrMqgXgSkNXT6DBVgTxi2S8DP65Ay+94GOp4/TAh9BDnll3e
4WipOyDEUhsueWOefiTcKf/Py+xaIbXwHgiCOA2AyBlLhTbHGoR5o/4c91ERQhRo
bk0fjx4zvmBh6H2ocdOF0yXURefmrsuY42L0MrZczQjUp+wypJLP+32r50NcLPAw
mgdj95pF6tt146WkXoZnWgRnuD3OVRqcUFKzTgK3cwQKRze2VP/abwSEEq61F+YE
LKtgHXnQgHwNdcErtBzI24UvxygElHoNJJ8Kunht7H9+Dsouw8uAOD8VyVYlqS+q
Wlzpkc3RrrhnxMWGtlL4iZ96R7hVbg6U6wrou8Ti/B6ig2NsYxUgkkal5D7+m3gg
6wOHmtiZosBsrVizxhJ799oW1G4Ao1sVHzSHvsC6mB//Py2UzJ9TZ+6gflQLGTHQ
bA8E3pKUljDREsw/ooXK6qnOD1HBh5uVIBxyLRB4hOcAOuSnOkVkxX7Bv1XonWBr
mrwvr8buvskhMKQ3YPyb8a22i23eawDONdxREJ5izbND3flXShqPxpHmDVPdgl4s
51zpiyecj5Mw5yTXONjLlICZ8AStsE6zwmEGAoBp5TBnOjxrAL7OyIuAmve7CPxm
MCM1SSygtJdJGqwbfxmKP8rOIAYhym6o90AZcUMxyAhnzhHEr3QbSVja2VKwT1lh
Yo2shsn42hfDef9MwCC4C5db3pTdnBO/MMtojd+PvAYtPDfiJ8AFbNAfJEQVTc3b
4OouEiaF8i5Q4B/+U2EyP5AbVXq1kzbbxjo7Vou9Zq1jYcwpsw5GVWAvZzRQtwdc
K2ygAidJooue3lk9HHYLqY3g4ok7zul7sXBrbwKn0IXRIkKUrNbL9XAf5szf9yYZ
6JZaG+TZNVsFC8jb/PjNeXj8xLIdz2COhSlZpqgTUqkWL/outt7jy9+x0YT4x9MO
DqJT3AErTiEeLZTVFfIS8K5yijJ0RjtZQk49ocaKNE1VokCKB0+mp+w8DDYX675o
mt7dJl44SFLJ9Tn5Rv9pp+A/hn+2v9VsJPGTqpOakG9hyfedGaaZIrWr8AOKkyrh
DJ/f+SIgRNw1IESQijC1gu6Cb9FNj6yqWAixi/xUuEPD2rl2yVuIbfjWgcj8tDC5
t9KXoR/WKZU4UAUgZwrv+QneymlK7G4mDhq/TzgMVbTOXDqyul5NYQvvwi28w6eO
QekZ3b7TS+F1+nyihZzTcao/fWnuxri+PNQsQFB7xRBj/0lSft8aloJl3f7zXoUQ
UWI2oaqDXm3AkOlkFev1I7pc3yT0oUmRnggftcXGcUCdRSSKkeKoU/HboL6+Qc0G
mmKVW9ZVNjr1c6cmCgeXOB5pK3+ZPOuCK79zsGpMuhbJpDhRDq/OiSGxrLeNnADk
qYgwiK3hr73xkpQTwl/xA27yNZvcmL6uZvysv4gz3pjVFwKQ7qRh5n9KmNVvi8tu
2J7iSwgRhqs4GvjQDh2+BtrekL/oISfizSLKNnALwX9Vebu8cweqcO39rHv576gh
7uHsp4l3BQPLK3WR7zSSEODbkgB1dVcXQ2KK3JIAjQX1OLGf2+TKsfUe1W/DJdLl
J1zAh0G/wF1iM2qytMZNcdOaNxUf6xSL8+zJqyh0/2u4qsfMa/4mvQgbD9BEXdI/
lDJTw6BFLRuGkj9VUt+s0RhjqZT0DGm3WD6iSjw5j7XJAhAdRrJ/i3C45W0E4f6V
kxfqMhuchX7f9e6M4qcce7IU6k2Z/t+SXdP9DDlStZW0Z1cyAOHOfrQPzAWFYbdn
v3bB4WhtY1nHC2K1LotwsXuZK6EJYH/W/0vH8AxWd7TqkcmpBPFNI3/MUnbcrasf
MP1+oPGckIlghDawPNEMgSiWSA0/pUWg91thq8tVK9wuZ4o3a20M5CGrI7Hc4vzN
sXAnCIBQ1B/xs8VPqdZgusk13bIC+BNAF2vBc/ZaQ9Km9hQo9gc7M34z9EUtbuyb
MlO6p8QLxFtQgmUlEmCZFMhIaGRiQAx1N8Hgk3iZt3S6GB6PicCcH5F+55HubY9/
ydpVdArtA5DCah53OP2U8ArGhaKEQsBsXfn9fUe9dxX+WI37I3FZqTkmfFfWyZoD
uStdhZKuchCJXOvNw2Jc3I7RbbEgBfBV2j2OZfwe3q4Yzv7RUTnNHSwlpOlUOVix
ThLnHSlu1iMI4o+YB31uONuIUHP6+Hu9Usu/q3eu74XX2jacbc0nq/J2pUPX3R8+
MoA5gRfjNnVlQICEhJ1fP8HplAyUkLY1qGItGMphBRQHOaRD/HsInimMuLdAdIAr
JeYpLLFz9Xl/H6UDhAFPKB+wZzuLPwgxgWRv2BiGDgZttBCRoai2tUN4IBBRLHWz
B9Q7UynnGHUtEUcg7OhepQhVVZFLgjkG7oTdwlViJ1N7Q8pDudiDythHWywe0pFb
CNVDzTOwJblWUbY8xwOkNe3EZc04sgUTDnDciGJ7+jkUilCUUHhvnWDrSjljtS2m
0RGqmy4GfLSsrqyzm9CvqiPvSlQoPqjGkxDZJDn2YtNA1YAIfCp2G23hmK1Xb/2o
skjFcLVdBPidBhKTt1MOLvdvDA64aki85nO0Fc62XDpuedG6kU4bmM1wcSh9fDkH
VXafh8oozxgdby3WF3lsWTZSYDuf5AxMrhbMpRQy2XcVF6vXiVxu+Fp3S/Y2Wdgt
DqUZc1+5yI+0sHZkvKwLAgdUA1b9FBFP1T2JFjwJeP/596f0A0HYABxOhQ7AA+8e
w/84V7pBK+eQItb7Kiu6MS+A9Bnf4a7imzSnnBS+hfkLEyb/D5jtTvpexkPmYPR9
Z9apbS1rbgXPImZgAJCgBnimGAfAEsyuiyQ6ffHnbCzIWssGJjdMzuawBEGskb47
Mnci4onMFXWRjZ9q5YgPhQXa4lCJx8P4xBCPNeO8IrZCmpQk9WrnKG2ti8mG28ZL
JUcPU8c18qgnEYzDWDdw6LiP/CDaEvDDNTN1R3jdzNy3KEl8pHr/zyGpvOnp2xUr
sM3Tbbej+50OGnjCdW8md1rZniV0CRa3p98Gt40bq0+DrwUTd6+o7ryBZSmlYDV0
giswtLLoEdBl4rw2swrk3fE2X3g6nUwyeXj4yW1kg+rwi/OqNXy0JNvEoWqfPdmJ
8bBcyu70RyP8EwR1P2JSPDLgsgIvXTxmW4jxPdtmEP1l//BlSWAFfnX54jOWb2X9
oy4emiAvJskgoiZrDcNWrYtxQNF4iYHIXwwrjSsLI3BhSzGbDdd7UZswyGhqcgO4
hDzIVRbjSjTEkMDTj4EpwNhD6qDS18ReIJlh5RDPnzwvCnGU8Cw0QhUnUtY/BhFt
mJWQNgdMRm5+xiYHUidd55m7+BEjRQ2ARMoGExJJV0Z6IXVPUk9mh0sGeeSZoJ3E
9YPN7Yfoge+1Gjvh5OdCHPGlEvwHXaD3TeM1K72Rr9aXZNSzmTCYkTUFDNRR9QtZ
yj8zvFFRP3yU6WPyL/uk8SSyo9JuPwphfuD6bEodN+9fcPbleg36uyPRcct04CDM
sEJvhdIGDlxyHoJuP7QNzBZaym99mbeGwNccofaNRAem2UoyMO2wfs/e8JaN08mk
N+LzEoLcdtoNCLLQ9YtRh9ZGTJ54lJK9L2mkUzNohvujhFhh84kPOTEuxgem/DKf
GuQNAaN17P14OfLrM9cEd4PgUUkvKjR2N4S7LObegxgWa5smQov6QR/lTepi4zrD
xdU90i5yPs5jDu2N6yM8kjdcFS9lpLMX1X1Oyc8kcw491Mw6+ofekxL5h+Gwaklu
N3ghgtWUcUl5vRS++mIeiWwN43sgQ5M3mBTc3oyDHcZ0e/4TFn3h4ncjZTRQkWIK
xAsc29bO7SVRxNp8qoCA24iRB7DrLd+n5X5wAXK7UYHQVpa8AJdj6Gf706YSa0UJ
m6TAovZHVJ+3hHDXjI2cZksdlBWpoYLSuDCz/BbDHxtUBtHfreZnnQKKLqMA5ROi
BhaPvv5P/w+C1LENo6p7ZAx95BzMxwKBgrbV/+R0ehOSQHvZ+eOchvH3nFJYnM8A
Pljgb2MPL6cGJ3zTjE3uH8NXzav5sBcAobSkaxH1g0sXU3QZFgyIOs3cnzI8HnYc
xuXwrNaMUbgakVuph3W3M3wNyt2lTYxvewXHtEZg4Casrg4lXbaoSVWMZTDEZEWr
t6ANio+7UncxCCkKVnBek+DIe6H0zPMfBs247vGOdM4jv7RKR9DpKvbI5npsqKtn
dkxOYY77uKnn5N5SCJk1G+gaArJaQ+Tsfp8nZuWgZ1Bj1n0dLSe59Dd1pw/lT5eX
uCS54QOyTzOgcWvQe8dmivhWZ/PsdXNkfB1bfiI4P8PWIjYSc38O4CLHANesu+tc
x0TAKnSjdrZcFcR17H+Vvi8me93KlxPR4f8p3OU2opr53Lp+g6lXLmdoz5JDBhO/
ikZNpkdfLQLhCWlvlOJy/6LyTX4xrdLI0NJFGvM06CqFukL+7kg4FS1QqgY/GnLx
CAfhAJOa/8PLAOmAMBW3AjoALhzMLmIy6w6J5Kw/rEHcB5CJSR7PIA8/Ve7+S1el
SW57oWtFIo0991ZoDZvJNVW1Bq8pKareeDU1whHTMFi3gYfI0Q0G5G2rpmAmGKrQ
XZ7eMuF1QEfJKGJKTcZ4CmVhPeQvVk95nij+x+XhbRDMy0YJjwomByNijqkv77/m
SJRNCmH8xzKGnXloQIIWAWwbtEPboVyiy+zi9jQPf/975jAtjbCOigtx+4JKGWby
Ydc8EMsEhdFnIf9UC4JwQBcG/RGwz44tWW9e0zyaRdrfbgNMVTEJc6LcOp/wyOEs
Wf05kqReeasIUyVVtP3p9SlMdMAmgoRL1DGIeM1JM3eJBqT1/2DDaDqeKHdbjYQG
nJWBOe9oU6oRU62gwNZto1OrHP+7HZYxQdaWNMR81nLTPNiAR2VfqcTuGWDA3Kn3
qHJGuUuzQuh9bEE17wjkNEmF1KwoeNFtrz6ilzvsOwwt0Cx10MTYi1U0TWxNKQXb
gxT3ftIIU5dFojf+ymnley8htYsUyUGFRfzqMkvId++my2AQtdzsszb+MFWiOX1B
iM3gzerjjsqBrprz7qM9UzM5Br8OUKnsffGzqn+6P+HCjyRIdaczkg0ulXGOdgXp
bQ+fXYZg5t+uwtvGXq+Gu8B3hjNIh9wlMOLI9+ZiR+th5TOCPQ0iVFFNHkxDuF43
mOSrvi9/4gCq9oyZo2THHroIOpitLkPaiAFoHca2KLIQcijzpDUrYLHH446tt0Cc
obcqut6ZOc2XfOInrWcrLXLc4btafbYDWSWVZiclJXnFWtdjtn5UcGzwR4i3kupP
RyI+y35u5qQcqjg380JOvh2P+Vy705HxGRI9JTHZEJhcVwR7+FpSZjb44ReQyZSw
7sehlkWn04nlt5t5LWf4eKXjAxVRwgJYIHQtTmtsVbVid5ut+76P2I2q178wvCYc
A+9HRgIh+zwiAt+gye9vGv1r7bmmpHSSijpT1bpfOd2lMG8eRlkbeqHYj2JmAZnZ
dg7M3Q4UMY0iyDmg27+GaQHau4Lj6ifI9g+TtW7NvY326DGfAbh1JTLd9wRZ9z+G
n15qyFmGO2w7gymy4G/Cic6CIxpQNAy/Regbh0d7eWbn+zbWGTcyZ3oUR/Da9SD4
rc/TdIF9HKGf5IdpAxh+tkb+GRMC3Tuv73yMLfx1mpIB7wHc36wNqwjDmKyf7gzJ
3IaL7X6qhi+ZgOVELUw20UutbJH5xeM9nixQviw9y58DSfE1LI+xS41GLVvNsMyP
22ZqSgVNgRbDJhk9bFJFBuqF9XYgKa7uF3/yGcySJbwKycJZgMxEY7RAkLj+aUhl
kzJCTRYyEOJA54E3S9akTBJ1PBOpC5mVnagoeFfRq3SdLQjkZwkkhEvXoGKuGXXl
gN2OVdt1+ya2X/ah13TOHQ9/qGsDZP76LaH8cyEiiNK2gShf02xiT4EI/LNK+hke
73VIeu1aNdvn2WANEI24wqNB7xIJc0Rx+Nev5nmwjeth0oYb1M5tMLjrPm2vAmof
H6EIDCfy9oDcvK8A6KNADz32pdz071n6G7H26HBGsevQByjc47qYsp+TaQNWCfv6
5RzLOXYgSxsSk/stKitdFQUM+w17Lo2RpknrOGK0L0AR+WzeyPK9cWZWu2QL8sag
ajet5sZgTWg3bRDuBWzRToJbrGUw3SNIOffMV6aEJNkmYpsnKbc65BS5tT4UP4hr
uTMcEnhwPLPwvSTwv6PIouf2cYmpkUrHwRUJgbQYSy5dXO2zQx7HJiwiriJ7+sSU
IVuY6C4yKM3mq9DNE+smspLPAvQhF2mMmn9vuEKai+eQZaHBAwlJiLSJOODX/tX/
QCQhCFBIWOr7pZwvltd5cXUBMNHpl2ye3yJtFHO9EwyNgNSClv5eMxLWURmWgPRt
G+MUAK6ca7efSq0fLxGEmwt34hc56Y4DYoX8bZmWXhicGXi/kE5ilXaZWhPlzBJE
Jw357qbbqcXO2HJP8/HUXBUB9VRjTGYuvykrF4byRfL+3PLVQe3SuTnqFAauNSzz
xDn6uYaIAt7BuZllJEXgxtXU2wM+3hRgAqRiRmi2AhkLliDyOYLMWUqJBtvVrQF8
G1z2bLTV0/McTo//4CUSVZ7UdGrVPIY5m6yztd1R9TwigtxrzLIEWNPjoigdqOUy
BsXDQT5ZfZr7TnUwlA5YZmHyCFsK30/1NxUj1ayaQTC7LkYBrf5dXpK+pjDal1hc
V2ddSXG1BqGP9RELHX8PLjUtEUqW448vaPIgDsrdWMFRUVDMaJDSD47kZwGHW1ZU
XSVsrSbwxoIONCcz+CHuc1Bsm/N4SmsV1sADypX0CYk5OVjfOughCf00VVFUIl4v
7TIRM5lUP/PvYIwbhSlLDq4d9I4f5MMPF/jCLPd48a9FG5qI50vGBTrlKMrHa0vw
uca0RN2kzh6qnxHIZqCN1nwpB09aCWc22pDrrp5hJEgt/8NXZ+eIZHs9x45O9EWf
HvTo54D3koDYV06GR3YZ6wrSg3/sg+3Fr9RCDT1K2NzlIgkPLmjBPTgM8D2eUvtq
GGr0xkh3U2M5AR2ICHilqaydLg1RvXjCfcwRCeu6zDSpa39LLZcRBNEQZzVGCEOQ
/ChOmEEOck7rX5SpPTlma4Uokd07ycLYW7UprnKoXGCH1lIcHeZEvEQY+4IkJogx
l4GkYWum16imDUlTsVam7R6EZdWhd5Fc41kxWUF5CQ0/6Mfu71zsRNLZ9+PTy4BP
gr6tDdM3hDhyhcblnU98GRg6RaJmaFlsHCUhvfCnD2PlGW5x9s3HCLyQuRbD6Q5S
Fsor+URXJzqSjfvCxdLocox0AvtmBIHjs09YA5PnKC5YbWggeXp47k4+6K8UIGoB
DD7By8M7gPEgln8+LofpAvgVAvBWTm+BnEOOHNMJtS93F96P5mxqXshME4UUhT8e
qalSS/oxm0W8XuHBvNYKwayC21yBb7GNgQfXWH70iXyNWgLXDGY94GHCwz2EnMG7
LFtjoaar+XEYHEEaZdcUGeTAYx7hSf1lxWKhyiF5n6n3qugyju7MM8PT+1rnTNRq
LXgkcYbd0mrgQLtQOMS34mcsTWtVSHgS1KbvvQQ+7BOWBvLYlUcAL+wPpytcMHoz
HIB7sES17dCC1IaWi8XcJgjj0UpPt5FRMkPALReULjuP8Jx1eJde4PrONn/GHWtu
vI6QeMqF4uh+2F/k1O0rVFJg4KVoJvyFPt2eX3QK/3IfG6PoqQmmbVBrCozUTPWS
z8g1HnDxDg3OcmljGlCYbGAMXjkbZ0juFhQvuyymUveAULbGcP128kV3PlyV4wqQ
MH9qTwqK2JldcsNuGuJ0LtZv0jGAkcXhsqImeMesmhWDZvNk0uydszI+mFZs7gBi
Kc8ewQ/vvbFl0/e9CTlR/ikiidpSBi7zX51ojRTuC3iydXJlHUrASppkfy1MkL+k
1rYG0f29FoeI0Kff5laNDzFDF8swqBx6CwqzO+1ivjtAxBUgY+BKr02jBf42HpIj
ht+/NHwtOFr4DpB3yeq2QSuWhXFHpyLKB1LdiwbYFXfn197EQ73GxAL2sYPWIhNr
zq+fiI2d3rVwh3DC75M2CoF8rxmBWNgFYM2rsdsF7hUzXP/nAHKl3FqdvqYjYXGI
TgmQrl+WMl41YgT41oIThsTrQE4RC0IKefFm/1IE2LGbKTZ6gBgfZFjzWDmZraXY
Ep1bwsYvo6kPfypZKWuvbVyHt991C0Oy3xWUm4YoR3b5elAPCOULowRoOGpGftot
SIWBHKeAa0YGOhnr7gAc3cWkIm1Tl2NIVcLZGV5l1d2Cx/ujFZ+ZOJM29V9o3rIL
xG25W6yritIbTeCOnj5lSzWZisARwiCwgNGI5XhqawrZlONCs5A3rI1PEPok84K5
QgA79RyyDyhNCs19b2RlaFvlxorZYzLiYWIzvdAftE11oykH7HoTcbac1QyFGowh
Xz0RiqyYbMxYxzES6Yy9y5DgtdsaFbihCJT9KuzF6nOi/6AEo/Z2w3OOPKVcMZfo
oqD1MtWZkhNkr5jVs0ttEtQJe3eHveAH2a1EYM6pBKReS8ikXmL7qIIjnz7ZSEDL
IO0V9AwlYqLmYy/rnALemfANXZQWQ9lEEcAub3nwIJsjpPgZW6g9EbxpQS8JTUdp
Ef3J9XPaL21bt/nUoa+uKWRdqFBUJn0FSNvwzJQwdI1jsbQ0aJD9UUqlr3CRuEn/
2cdRU6ZszA+tZh7ItoHeIk/VPE3p1wC12UMDayAxJ6n1U9XfQIm6bQcc8Z7dr1Wh
EuxwMexZqIc7GbGDuRscinj7exnoR0If9n1/69ivjtO10tSuxr+Tu9KoXHcsTqyU
Tx4IYpBXRlT2ty7AipVKscqDbzwq2PcsanXBqeopbc/L1gg1/ALWYFXGNECcNF4M
cw+mNPTzVnWHRD7cmSPtkGKHx93qXM56/8RgUAPFaZ/Ix4O5j+JgVHZ+kq86VuZi
QU8zqrvxIU17DF5RisNehvYPij6lAJcZFBzHLOja3yfgG+VUNdxnh8Xd6MvaLEu7
6U+Q1mIsynWzKfsXvLOoAFtq4gko4F71VY2iJFqwk6WftwiuHcI4Pw8+TZyYkQ1m
y1n1upfOCBjwGvsRVwA13HjXPZYIDloW7Pw0JgQImzfuqy1nAjFoxG9ko5gvh4MR
WbQRFRuFYAjhNy/2lwB4T5URoLrS0Nw4q3LsCP02pKWbVhjHvzUPMN/FNXxyBDB2
xfaLf+PIAY3L/QsgAUGmyeABojqhjB/BET8l7sEITHnCxHAXf1lALzAlpzAkvPoD
mCrm34/2xNOhwD7L9mzoE9l889I8Yh7wyeB4nfLzoUWBruZyMF/jsW4kfXHf2VjQ
j6Td1CeyW8FMiBy69tLI1gofYZg5xrqYTQ5JHREq7S3UrzZTrwIGYh7/mls6SWQs
dxJLRV2gl972GaJZkaYBBvbUo6Oq4xqV4CvXqNVyn1FD/a6IYJAIBvflis7Tz9qO
nGc+uR02trYV8BmWT24uHEJlSmnaBXPm39zqi1nA4RSLFlFHZ/4RkMLloEQy0Em9
XgQVUL3aKINug10Dtfpu4x0J23u59bvW5GDljt3B+TswnD1mzVzK3FNTJC9vIBqE
qi/pMEIzHRFACdibTWLs2i611/a/HGfuDbzHoO9V7ZWi+MSoBsXeDN8CNA6JwPr/
SDud7rUITJrL+mSFbx8UVWGrE/Pnv0t+LhT+48IvBHUnhG/2iO1QyxXZWI6A2KZb
QOJaie66gXXcAtn5JuABoZUPLXe1yUY2TZbDmMfMDMeQFiDkyWIUIckDJ2+MsGL1
VMUs2eHjj+R4zVV3Fwril65gSL4FULhEXVWgKGaWcHiwOXg/tYGQsu79molC+4pQ
ShqLEyJx3fIkabPHcgBqIpLvoAVe4XHcIpTVoVJFxKjiyZn1ZNUod2DYVwgBOzZu
gkaeqAG4leK2hCheJNEZRWFiwvnpmDZxZWLqCu3EO7h/E7Am3v8Wvu1dxc1XrpRf
R1WYLl9p0TEPaL0sTWiAB6tVF3G10zSp2Zg6jRZZQwuf9NZkEAcKG0b45QQKc9Mn
ERq3S1QBjQLcYf3Zo1H5EFeWiDWTGNBmaKmLG9QJZUlFKoST46E5mBcAiyNT8x7n
3aB9XDzEteA27d/5K/gdezTEUIfimH2D478sdukREbHzjapQuaxYn8j3DrdrSHJt
qSJ6d0r5A5MgsP/WnOjoczX02fvvBY1Cg16dbg0hmoLXJ7mhXfGeH0ZPhtjXhVkE
sDfnpBxdYdPdlfaI4pZima3ANXyI1AAx/HO+XI+/g+IkQK3GJpAR1HGqIVqGbCqi
OaKnW5TN3d/psxixFEqJ72mIvjy2UilkCtZ0kJNlnLQ/rDVlne6pS4mqC+6i45NA
IsHNsOxOaY5CCqABy/I9kCgjZASHnBuYN0YXW0PEbCOlUvkzaGHvk2xu475hoRR6
J/nOa/nzioIZRifTrh5Qu4YB75wAZmyaq+18UpYqJjGPslC9bufvAbmKxMCtgEP4
xU67NIGpR2ZBvz0ZaxaVJGkDRQQ7mDEA2GJniurkw+QEbzlb/RRqqDvTf3dD9ulA
dHp3ESGqUbC5SH4GHdydXvY1KCeBNUSNLjsS7keFfEwaGZzVWC1M6hGpNQt9qPoq
qGFwbLaIO2i6bQoOPyiU6F6V4/enD+633cbE4wDQmIDC4T6RohTK8g9gB/rfv9VC
eaB8HI0doZNXVU/iR0zworZiP9nbxqACHmN0HgOJBlJoCGCN9ECap2syZbFcsa2d
bS11+HIlyzsAcEn6+E5/mdzJmqF6LhZBoS46XLHIGFEorqGhAhIR09zpDYkhFmog
j2r4ruEpcsqP/1Amx0rqPz+6494Ra03N1USOeVWaJyc4+8noBsxXVg9JaiHbaan6
wnKtVYl3i52DFAnIzuDy9Tprq7ETa9XzlFxRAssFUiXBUThbaJQljgTQumv9ZdEG
LZV/MgCNdOFb8tRabEOtjMwLSJowkOILHeth5dy0m+AqKM5GXK0ab3sijlN7WCBx
qZZCJ9RGQ9F+l9pQLmnO8x2ibDua+PFdQqxANRBeg6aet1IKnd6qS5JjrjWXywRt
T+4bP8wPQuqMx5j0tC37nJeduZoXYkqEtNVZBrP4JdJ9neXQO5Wfp1A1xqMiKyoH
QAUYH6/1r5/l+RPrMwNDTi8RFgyxr1w/FOsAN/WGZ7Tdm3e1cVjaBQnwXCunPCI9
E7ZE/5SoIwDBknTy1jS8wfqSB+yTLSJg6tvsBAso8Q2TRHxQ5E1mlJUeVYv7GzOx
Xa4tEQoCiU2UVNcZITXuTc1Y+XdTwaInS7eef3X7lHKbNUCkNkWnQcpc7GSU3cdC
Uh9im+zjmCSEr8vn0tU36eCd1MmXZAJpSXpXRB3EVWwhKPzpQMHig4K2d2vxEjrY
iII6a4pAT0IA5ocsi1ZQcm+LUNR9mh1/PsDqzrN5oCGHcnfN1FZKP2dXkrOF6Pbb
eBk2G0wiPhmbbWWTXZU6JJealChlSMbxP+fTEKPzU3lrrm/n5CevobKMZ+ld0PQ4
HenP+U0Pouqw5AbaGBhq83QRIEU36GCesomNXv3nbK6Dq79v77ge5xvxlm6l6/il
eP1IE0OOG4npLRLeLQsrjrZEAijrn8TRdSepfGjOVXv1x4qtkYc4JzMEBHEae3od
iSIXQRdEbWF6n6WhRuQvP58XJmThqMgVP81S45apv4luKwl6//sr4SPaeGkCcJQl
vItkZejHGusKySBsImWKw7Pk/MP/6tUsZ+rbWG4mMKq5CxeRfAjVkAbK9JOK+Uvr
Bf9D6bjThMB1STvI6uk9Rc5JDgJW6u0Vn9eCT5QpPYnM7YSgRQzLoF9TqJ8EiZ8G
urYitpmtnPOxhHvaaMaT86kO5FefjX/IX2x+3dL3J8fUa1OkQ/pLudef4jL6jV1F
LznZtw/9NAe4//kCARwlbNnBT83mtefptsK6JmSYHZ6kcVxRuugmJKW6xgZuDjXH
SnTvDXfgWLvNp70d7O7CCSjVR+v19CrvkA5tKkJdVGAlSbWQOfaZlxYPn3uu6wQs
Cdpu3zjA1lQxgP2aCZUchbfbjcxoepHV9SqqZpk0Fal+f7jZRcHvdu9FvLaAOdVh
yJhdOmv32lWbfJXH1YDn3/6Yv7B349JIyuErVDmn6p8f6uKOA1XJztoCTlnIxjhm
KfNGwX8hIc7aG5ykDeSolH5D5sCisH5n3+VbzBm0nQKVhFeOm6kYEfSStWlpXEyP
rDdCMzdg3oIe+WxtsQ9plLpBg62FjEIsQnWEhUdldCGOPh0P5E9hsqCE/dIJ3f1G
w+4qEg8IcRb36OVcZvkK7+FM3S5Rn1BLOI0sSPZP620wrbLcC1/DpVD0CSUIEEEa
uADqvlz8XzlxccfkNFNIMWp187/+YDXim3wXAjCNxKQQ56VWxIqqoDa9xX5hjYhF
wxvOnZJunj0/0CQuxGHYQ0byf0u42akyuLWAUXzZdviASlkFeRo7wo3VVZxteo+o
XcCymVk6EWf/w+tCl+6Wa1PqdDhG4E7Dy/M6+ViaPD6VQVZSjaXW3KIz8dGfDo4O
SQf7KTnh0KJCxHfEHON1GRXcs4mv8hEsP4bTcMEbtVpCUM6ED/jUxj170NS2qOnP
j+nFfzRpd/38KLEnZP1KFVqAtEun5pWlW4Dpga6Ch9erwmuRk1W9AazmldiTnmIs
d9zlOb5EYHhEOjI5VBKkuYY1GiauJPjWK2jCOfsFtsLiAA6BGSiy2qIIpXk46m8G
Hcw9btx3gxfOtHANjqW/mAnwyngxb55V0kqXPux1Q04LAl6QcFDkteO0kF0nY4XY
uaSF4wrHd7YbfwVGPA7iX2U51CAT7+pDZGHtGgZgixjq4H4Gmo50Uw4Hxb12hPq/
27kVCulPP2q2r77J/8ewxlPwhwQTB46WYqnhTpGS4hYQPtE+ZAu5uHIloCldZshb
iTBuT2IQmlWqDWrjoXECqPyDin8w/0HfXLgB+G266K8sH3CdcI2DelloyjL+1CBE
umgGt6gpJV7dguixL1u9KAo1/+8MNmTtCGxvST4x2PNW7CtE8VbiWFrN8TwwcteN
iNL8abJd5jKKTx1qa6lYUH9lwit8MpPs2iBn0MF8l0Bm7N0Wf9ok5xUjJBNqUzcT
rJJyHCmjbFgc/5xQw14Oj4VdXv7S2RWBWO+d4vfm9HQ5H3l42iqp2+1SAhaC0uZ3
X4v3clNzcIAwz6Bg2w5vpY5QLLXdLqnjo/Drz2Cfzfik7G9BQBxMISJThep9cQRp
6B+ZiJ4NB46kUy2apdF1Juaz9w3rbyoPLBAV0tD8YVqP84Z4gpLaBKvU7YDv8Biy
ftemSDYMbsMzrxTFjW0piC3lA9rX/m0QjGdDL8vDb8Kh0YNqh6DQpXs5ezfUrdPe
WjEEjhO5upcvW8sCkSup6oNmPK387vuZ2ZEbm5HxmOp52OkCcWIT+4Dk61c4yNfH
td1t+PL+ezAo2NilJ1oDGb0MRhqUyhLg7rL0XRAKArK5ufiR5x9EUecbrbPWq1s6
SQXsvT4ZeJmHFVPisFb54mU9upADW9gzjHLuHWLpP/jYZQMVkBhbApV1qp/6FH39
aWFVEK1JR51HHHTvDJ7Q22xiv13iq1q3EGt4QHMvCwKtv3HB7cM+9ksB07eqQxWO
So6mp8ZX76HjgqTJfVdk91C12OjTE732kzFyGzq3RFm1sWbCXFWLyNHpMzGSzpn/
W+stVxKzIT/ZcE8zsqFpOYZBAHjz6mDKwL0iuw98fAN6Z+w6kTKH7mWiLxVyvRC/
2lVyk6Ry1SbXglVs4VKAkncXALiJ4Ow7PzIAuQYyKJfij9Ap/DDpqQ/m3HsHzGVl
/xUm0apHD0S5vzeAivv8YJat+SFx5eS+1nfbIP5y1czUCRNa3214cIhexOcA7gMF
Q3iG7j5R9/J0K0tuOvnlS2x5pKjpR6mTshPVAtcpnx+BdkZbaMlck5X8uMY3hkfh
BSRt4eFsl0XGkOG+JzepNUnC7iVsV6w4P5foi9DsmVr92H1wmqhN4GU8BvXpX8xq
fn3bw5yjg4kMHbuow4+azZbxJ3lgzcn/d9rErTM5UZur/SWVEHtMOd1LPt6RsaXQ
Llw38X6WRDOF0Xc32BxIoB2wU2SKUOTgobfAXPcTy/FyR6ZvQU/inOCD5iHZJOsL
tOI+1AlpBhi4z/7I8Wl/PuTdn9n4dwtvfBDymrV+X2G67dqOI4sPeL//eMOeHo1E
Be863iFbSOanNGTO7B8jCUGhsu6Tepho1VCedjFKmr6V3U1yU9AUJSHIU6+k8wOC
NyRg5HxDWSwXcMdA5vvGNJUlNDyRZn1igynAbidk8xGG3cws6sZniOIr0z5+08la
i+tRisLdFzA4vawNkcCkCgOXA15z9NlkfbqNV/rBcXw2NMX14L2360s1e0WBTZeb
ggNXqepRgcqLQalzmXHlWCE08RbHvZe2jhQK8/K65RPi8mOBo/2g1G3rw8jYqovS
c3NfeeXE5ICX4VYyizc0B41apU2fDUDjZfmRnI4GRRYQc95p+yB2uHDb6BTlLBJ7
Aud4XbzsUNsbylgXR0D4yQ7mpqhTapilxIoVECLpeKezr3DPkec9W/+vFuzD7i2Q
G9urXxskcK8d/D3zRqPeALDzDdSNu9v3HtuXM/2kbHeW02hD+7U2enYtV73aQ8/j
m+yYIp7cdWBsX/OfvaQsrpJpnACyyaIMHsPP06WBo2g1TqkKtqfM2FI1z2vezi3C
mmZsYGgoh+Acad5VYFYI92Saff8DwG/lQ83n46g/hp3tBI5I/TvrQPt2F38VIDIK
VocwWZaAI83M+T55Xn0dB2EfwGoS0HY6CiAgWWAmHH8mHIcSaDThnRJrOF2SVtEM
ptSoVlq2vx0cJ7o8/nuAnJ6dcRt8H/nwmJxO3F8scjzY7B+3fZRX8R0HsoS6oBc8
Mga7LxAM0qmnM3kFtVksV9hiziyduvXdQSHOuW7HNOIPyyvRNP2cnWDWVSriBl17
2PpFyAUkAkCyjA/bweOV5/WgvmO+Rgc02mNUYTrTiSQJ9PF1WefKHbVrTG4z+Vt9
oejzwO6RlcAaTCJNlrOwakyE2m/zrRxt6jAAT4y/jCZNMgg9hk1KMyfg88i/qRw/
I3WedNDyMiFW9SDsWGdf7JdQyGuwJ1sPSgpiIsPaGGIhIDjHI17Dhphy6FcznzdZ
hCLjcljRjIhdpaBfM7XQJAngpvYg0nD1E4jrJ0MVgbLzV/sK94s7fJflPsdGoI2q
ggqnlQAkP8BdsSRiv2sRwQqyNYn+/sPHYJw1SIKuN7hIPnpeHqhuuK150J+YPHdX
PhTQUVeX+ac0U0M++jaV3shlDJyXseo4QGaM+mDPUxoE/b+dhv+/svzfd6NfUhr5
2TySiy1kVoVQ/kCxen1kl/DRlbtp5labMa+5KHxXf4rDnAbs9X4SaVVwwEn+FRQD
wvO30/v/X2/ms08wBn1nsMLx0S+lqYOZrsO2uSjTkKUql/Z1kvVZllc/1eXvZiNj
t7BvLzf++DZkuCzzV5bROzgJVEfjK9Nv1iOnOWRQ5NU3iDMpMyEjeFUnrCv5cM43
OR+I+GL/gts5hBGeDPT7rGyGQwIIUacVKspLfrRKAZNyWDxSzV/QrlI6SNJ57eaD
BrPInrwl1MxoW47LzxbJuYhSrFcnC3v5t6OYWKvZzJt6kEcJUrLSfmGHCtS5cmrZ
Bg0FIE9OOJYl7dMNla9okuxJWvaIc4AvmBHVPpzxyLjCLBaj6Gx/bdBRm/7XZrD8
eZFNNPozrPrYulXSW80Lcbq4V3lJoGWbSARk3z5utSEqQemY71RINZb/8L0o/LfW
TFIOJ5yhK8T3Xg8JZt6bE2nhvUQlj+vNEDqNBsVOzxx387puh4zHuN7N1X9oHE95
qskYMbOTyEuwmzQk+lRUcKU+CQzAUDgGIURhiFyPpGPogEs8cEsxZEAXJfG6MdAZ
ggS3tNFh6OZACfUKw3Fvj9etuW+rieIIzyQx6QNaBARUNhGUNy8uzc1y8IdcMd1k
iZSPmh7PbRCoDrrJmsqlYLsHmidYKbONrrActQDvc+lk756EodyNHZiIwRUaa6Zh
yVhrFZw+r1Tcr+/i5WNTOWituN0TLz4vTRcS4yM7qsr96Jmhqt7Vaqn9qFLa+X/Z
cjGLrvTQLbXP0IT5VokMDMkg4t3zqw9pLq0QrMokS+nE25lAd3+DKoPJ8Ca5FPEm
BFgCmUgSOb6lZSLX6Gsw7MKQCT0aIJZFD6Ja9RSV0ybWAdTbWf5c0eUf/i8TZeDK
+AFbJQJJzw1gvr9hedVFM2ZjXPIhYiuAqKb27UI5XFYStlSq2O8IHh6X55BrzMH3
tnGpBoiH7vXtbqd3EdtdWf4ucxurRQkkT9ku4XjcxdDTOIDWtzeuZplPBaIJrnQK
EnIJc8RfDEEo+tsjhwZsKWSKhYVD/nxnPIZGkd7Gu74ZlnwxrwsN3ijDra7slDwh
f33Dvg2L6jPgOUhsfK931+vFsnAu9/gREQ7vbFB1AmlNeyssThzC4TDugoj9SzjR
1FQyt47GzQ4p+t+leGPEaWCMJmCGlnPPOJPcpPkKB4zcVWaJ0eXCRnnhDN7TuPsw
/bCOsYnW9pr3s+cxCFEUxu/8zxQJXu6UbDu8ab4136tpTwDK0d5IYJTAIlidhEy6
Z3DNom85+7JidV5qjfzh0nMXpstMtsiGLFIU9cQIFokxuD1maYGQloUqOOYS5ZNW
nAxzWA5TpDBSyCiNCUUkdAGio4wgCBO7npNN93+zYeafoSfXnZp5UcrVNbjIEkQt
szD69QgOT/JvQ/PTI7DarXYiMrF9b5BaX6vA5E+HqK+eLViR1qfxZ44kTRZqcTts
8CFuB62YxVORe4r2t7vKSsslyHQf6iVlGv9U1TBJ9UYOMI/0EGU9D9SXTMO6TVod
XO/3Bv2f7Ok+Iux4TMEJNP+4NTPxk9McMlmIoi7YwOlKY6cDvlYE3g+WhCF45pRN
090ijPBAdbEJmYe7m0KsdE2KAIboGOJtlrPZtfcqhtD4tDpHO8u70QThYyfH9Lo2
hG+l/BiRGDTBQd7cVWsBlTAEAoHkoeZI/BZHMrDQNXeVk932/MoltqCoWsSVa5s7
IDe1wJuwDUWk2u4EfXwu7MvmqJbJ1p5jW7j29GDd+OyPc7oFZIapcTWFvuhJLvUU
0DO0xO4neabyxJ4l0Gmham+nLjs4PxVqMT6bZiqnEZ6oYpfK8oCrPG7CxFIJxtVr
N9e912xag6s0Di4C13de6Y8n7xkd2FGxKHdHTGFiUC+rmEFR0dCVP8iiThVtY7aX
pp4mY4osJC1vdGUp3tzlI7/0TZ8qVKgdkpgNdEfd+Pe+s6p3RQmx2vCcCZxFJ//p
MkTDHrhBF81ufcwwp0t1inchUrgLfnjucKFgSTGfcgE6GLshEGpDnQUPvAjf7tAO
tr8JzQHd1T+UZ33j15N56e/WXHXbEZ/fYrEJne3cthVByKQayqnZD3NaMtIc53zU
22xNB+O4oFXwYAG6vCLeOq7hyCQhfnkqYNNDpq4EKe5OXBC40kovgZW+n8f4seJv
y3WTCgS7Lr8Ncpm0i+QqjQs4lfzS0RAp1kcjFDKqXx17a/LTRwwgf4Oh3kPcRrQd
pSmlSmJS5BIPg05J/0HRV2AbuDMHaYmEveZm++zPDc99+5SJa9jBljAfnilehZ47
aeA/uidWuq8cXGwhIPZPxzgnudeB/itAxCJpsIR0pJQV4Odiq+AuIN+xwTHk50we
xUR1EVyW0zf81849sjbns135NmySBrg0S9bXcn8/wC5r1x/7R7vma4JV9GtpeEjS
6Ymsv+YdlGjQosO/TVWcHqmIvJ8hXTpDCUBIJpe6zC+poAeO6Dy0m29DhYU1Wtd9
C5GaGKBYaDMdHsT2THViP+qh9d+f0Yb7iltqj2k0lXKw7ORtGm8p4KLHfdM5elti
F//wXZkyO3tIJrGnykjOjwylTfyo1nCarF3Y5f9pCiXKJ4APxTEyvUGCOKpS/hqy
pdmFrp2UyKSk2KjwewFGa74MkJv2N6TkQrzIFrAWIjtQsbkHpxxkqYFPeV83VEJa
zHlobZzGDVUFQ3kOWF5IPxqp1paiS8BxfLjR3IUCuYnUuiyvqyvdPQfUBS+ghHic
jP/jbsKAnIFebsaEUrilt08IJ8hm8iITjg0c1kUlgtjIJ3wK98yqwynBHGtuhPUY
a6oxxn/QlNkL1xw2TOBTxNtq4aUNktkkoy1LlYU3IfIPIvpekM7nN/KLZSM4/Pn9
LQ+oKgVUZKkRN8CHjSOcJQG+AKYHAUZ174sJnUYLNU4Y/lIbDoV2/2Slo1E93zyo
RtuiUWBhFIXQiX/alffIL0pdhft1kBravORuYNEF8zEr7hDS4iiwiI+TJEmjYcfQ
kZeJ7bJRlaSKnbKTcB0RfX4Z8GyHnPMyhhN+BUbbORGNHApKFaWrjHyLyBxn9pT6
K+I03UpOl1llTKCeolh3pyvt0EaK64QcHEdMjLmR0OLNZgt1oyNYkvIMljlLf0H3
yKEaFZZwgjUclrUfZHsbWtPjAq1DlcWS8hWcr6z+zQkUekdR39kGAwcHNTJXV2Q4
9xVmbS7zXLNJzO2qceCE9QJMDsNOeb17FqwUvML9s6bK6QeN7cRhS4eoqHkEoPHu
zGAjjOgRXEjAFz4EUVt2mAuodTlL8MirU6TrRLFupS032zm8DLOE/CBF7X6AKoUa
6pB+ut+26Y49TSkv8bQHaFZKshLBcUgSny5FRvL4+X34MEaNnrtqexd8mywCJtNJ
xHgsGvLBdhBr6MsXYm2cL7BuDoFT52DvTYvat+blhcym2t/7vIC3egy+18ZSmMH3
KBvHBBX9PCgawiq/47TmlxFRvl3v5lCTLLRTWtXHQu8PQmogFt4JTyx2SUBHIMW8
baGMEj0JuxvoevNXU2P4LqyCLhUdNWV3OqkfVFyFZD7IdsR1zSB64rWl+jBgGGRD
6tjrEgJaSTJtedJosENZedkX71uohu6rjWwpPRlTyKwiMulHI2+8t4rLzh0qNhQM
G9/emAR6jefeWR6jUxoo+zcH+MyD71mYsZskTkaF+DSjys5kHfAlYSQREmgRGvC0
z134+AxOPEmHcVwcBno/sfgFxWEM446S+WsankGAHfKC7tQx+pJAH5Y9ha1SU8lC
LNQgFlc7L/tHlU/XgXRASbLkIFTTIG1DSZyJBScJSJTkMBOaOMSonqiYwyKYtT4m
cg2e600iMU8cXpeUPlLuPBZoZOixF1IsksPSZLf6MtH2y62+9ICTZeRtPjqEaygc
NYYL1+PyE0OAYqoV8omYLXAhAiUDTRRZY9wYOhLceLlX0DWEgoWJbcMd2clVHedH
KdT8iWSdmHP4hVIPOmK0q4tKfSyq+9DhK0PNpszrjfIzypiMDOPxm6D2TPlki+h3
E6gDWOxKZ1iBMK0TrXWPnXPdfBcR8nTtpYc2drnIcl4s3gaBbTaJilCA5d/e7Fks
KWmula/HwvAwj0iubjnz5Jgo4t0fgbgd9/BZ3nLTZAP6oDzQJ7+WBxbuWZ+VVsJS
X/9wPjxncSHXGAjiYP4f2Y4sVyP6BSkWmnmeQAhxypH1NMPv6RYpUMiF36MU29SY
Nlv6fVbQ/CZB7bcKBP49U2B7x8B8FcJd6MY743KaXKkCyH+jBqvvfnosVjpzPPGF
PhNGaxzx9XFe2m0NXCPRXDl1dkUlL1PajirRyMl+ue+tfqbKgTORb35/Oo/ygesJ
s5SDEcECkHmhPz7Hsw2Hy70Nrbt8DRcXRtO1AMcl9vk0++Li92yyU1O7MXHFyB7x
7LJxMoJpKs6Yp4SuDX/5AuY0heIOmaw3WjE0etIggKyBQ5u5SMKa4ha0EhLHzrIR
Ajc2OIg/kkVZH+3N6Hb8FS8I80iYmkcqwsjLeaBfCEzoq+ivpu56An80X70Nxoge
NGTklGCpzjrc+RrWInYCDhVJPnqsScHH+BaK3PbzrcvIug+YX1YkgLp8A6ZapCH/
jfdbuCEOPhDNlsdV9rBaJVw0x8Fq/mubDeoknwu8goRtymNRuwE07t8ljZIQFLmb
xGea1BddYmJAXCpXMkHceBd5l4LWMF6iRBBtIByQytz7Myl3y+TzV+TxgRkCtJp/
qtL+zUb7/BLX0DYU/Ux6Jc/dcycVUC/4vHBqR2UIZVMcjBlowZJLVsy2l2Mzzj3e
LmHWSgaiSvFXrEVVl8IKGk7XoA7mziRue/4u4fMd+rrDfDImFNsTA1iS3LONz+Ef
8J6hO5VyL+KRE2YZrUEmdh5S9pHcG84YLMWkHrMXukQmvRDv5FPYJ3xibsaz2kDE
32LNaE09mmBmY5z33jsQ/ceXd4vxDaoc/QcRPoEAQWz0wm/wYrHJb1mfCA+upOyg
yHLkep1M6Haz2oay/67XMc6cx2vUp/pT19ayBVwgmLx9lp9r7sQQYVC9x8sQm++f
M/yARRHZSs/OdJrOieTVCsI2EjDWSalwIbNFC8ChFZdSqpylAn3oLH2Iufo8pqS5
AB3ozHCQmvAfZNt4B9L0SinoD0bQ8eYihfx2MCZqzuhGrQviNeQRkL0swVfcXtvH
0KCEOWOLRn4YcmV+BHrriGdiHQRQl+vQ3NGcmwVa5rNBHylaTkgV71tuCGbYaZLC
Q5b79VvZDRwi0Sswmvp06b9yCzApBBAjtR2ZXfEclNSgLqw/93CqKJ7e58VFI8Gd
R/BLQ4AWwJ7csvyl0b0Ey9DdcVci84adbUyddPcRH45DluUfu4wOhvUWzi8En89N
t8p8rVapw5fJtobmeR5cLLgkoo4zturaGwPtF24XS2T4B1AHKukdGE3IPGZ7sGhy
qwWWpz83ETA+vMEgifpuRCphtGlN/UF0plq1A10WQ8vN2bUFVimKPlruX5nZVW/O
Tq/W8p2FfBPn1ee9i011VqbDrZND7BNc1vIHdy9qh844qZsV6ZkbMm08GL5XjP2k
1D7oYASVEuQ3TMpkW9Jt+T9CMst9bBOGuKFPG6AqmUkIydBrW7CCAXI8CRgv2g7K
yTRG+Ipr1Hn+sRYOIKG6oZzyvlSkPgM0ZwQhuZM8WMdPy3VpNpQn8kAKhCDMQzUV
h+CzT+T8XkkLvZ7rFCt7FZWBJQvfoWR5B16Le6LC/h1+v7p9TrQUhQmGJHUffgjZ
fkUar+owuVSi93VSYeURCrm6m+YuF8aCPIFP1N5qFjuBgMbVera5aNxHR/CdnY5z
B0g6ipIOagwlCdYZ5ksNKCGTc2hA2rcILRqT5Pvx4ri+buhTxjP3+oyCyvkFHffu
fpvuadX6YQKzl9gUVMrPj06SfZHN3ONf2EM2uyf83/Eu/GrguASoHNgf3Ty0fXsd
9ipxFhjb1un0QKBhyTBUhwLFxGqjJg0+C4t/gm62F8vbXHgvh8LDp7cAKmZcufnU
/8FnyN10NwYyJ0ROVqTM+M9AGg3xZnrQscIUQyOC5yFkTDTrp1Fc+6eak2eT7MkA
KgPAPNFiJJ1aEaC+LMLZSBoZHqqRDuvo/6eCLNXXiUASYKJ9X82yppKYSlUJ7G+5
REpLfXmPq9GJ5B2rnpCw8yMbIr8508oAYskMVwkjJTUZuahD/NhwloxADd56mpd2
RdHHr/GRTKpZhj+Ij+arxvPPYJg8gbpfEgxmCA+MxTUJdcvCmifEzzjjuYxv/wpq
NTkJK2JVBP1EkFdQSUqUXTWseB/zOrTkcvpn3tTTyX84TCa7rxeIim+8WyjdpLWw
dc2MEe9BbuCxor2wtBJHbFhVZfFE12GwBx7xJld3QQVraS4K0oPzYPGUvdjTT7HA
HuV3JkFei06T0FpasnXw7MzVh6m82INPKarB6LnITP0+h4g1gmT1+TEKeIfxR7nT
yRfqeH5KGnuJqb0qDQ467nIiuRyqmGEugg/NmKvlK3nDI1IU8AUMkxzRVxUWUw3I
VWbD6ea29AFROuNYScM68RHZydE5ZLVec8XY4FnleORYWC39PWG1OzE4sEvl5lGR
a8ApWkftvegCY+2VTRrYStI3VRuD3/pyvwWDGz2KAJ8FHhOwCkOyYMx7J0vNY1zU
cmWkZ7jAWrEQG38bD4GMzRVNxnYK53uMtIQoXV14UYxRLJjDZObPp2ezg8BeSmQH
sCheMWDwZ+D+dM37n7/wQu1IeRTxaECBjfoAFcIc5kB9rjsixgP4TyZJ8KtJw9JG
lec9xSI/yxkqk6As2exqzb/WGHevix3YsHvmiHMyV5EX6m3XYpyzvXePo8z3UkAc
7eQD+mYOH2Mz3Zd8GIMa0C7XQb5vy5xld71MzRfizulDhf87A1HRcSwxx5aZMBz5
j1tfdLwT9OhVd4nxG0UZVcpQRhouwEQiMP0ysS9PTDJpjC99SHddEMraNDL0DjxC
S3ZVE7G1P+W92z6JhHb5kZcnBkNNEItJUHhpZZA+Mv/UbuJkYtaHigibS4Q4VzCV
+CrP6QbZPNnfwCww413NwjyUuEL+E7CK4Zw/uGMtiO9FZWsMUkDrtox8SzCwLFAV
7afYEHqzee1V1/aw5xRY2kIejuqxZ5un3LkVisIS0PhLiP3g1emrNaiqA72qDTh8
QQcFV3cS0+rzABxPIvBqVYN+e3AstDu0DVPhW2q3ue85xlMIXO+K8wu9OACGs+T9
qQtJc+4KMi9Z/WrDUGlyrRneyISqddtFVieqhVulhZ1Uw0KU9B3akeysEumAQFUA
MK14HtdSNrTndEXQajVM9pWZKoK16XYIib7UBeXGQJsYF6rj658QmOGR4qnpp8i6
VgP0vUJrup0Axt7Lmt7aKlW5lhMUmZdTdpWwoVHSaqNXsg+9wOMU7sIo07O7ctRs
/pw5y3ccpMsxNEc9vlZ35TWnAzfSLTP6itKr3SWzuVf7HLTHSj4uQyYPRNIXalsk
phMb3xsPlCi52K0jEHpf0xsXHUeuraZAdVnsS7iE99tcr44ATTdOW2PeuDu/TXjN
xjwHADfm66qfXeUcrEl4HlLxD7vbGcW9nuT42xSmtSZ/nCAnRT3HasHIJTYWLidg
l/fj++1eXh9c2ulmZC/jiqdqKGyRtckgAOA6R6O9eu7kPRTmwL8U3vuQL+Kdm8UI
WnRBYO8Q4tEkDh6QHelKfzttYgh9H3XlyHAzQCSj8vh71Xir/VDQjqKEv62yr5tM
Zbn0ZfVx19B9aSjOgdiQqIjHDrVZnDCGwh/0lUDAbCW27B3qXCP+ntEZJ0O26XFF
m46pViwQcjIUAwncuFaYqIpqb1cwBhWJ29SMTcvkqXV2PNfIGi/bIiKhP0s11ZJl
nmfYyiq/cQYSZDIMkAnSOqMJ+HWZO6NOehUlRHa7avDyrscrQQmnI0NXdG9vK6/U
/jC9AbNifecXGTeqmENcYLmwH4C/NZsv4BZ8qgUjWj2qC5r39PpKWeIUyOTTRvKo
F0WRjB4MAWq7xZpG/ZHphE7v9LpG2NMfEcSyRPHKMvlBNwIcQ048lo390xhG14EP
2XyGglaBlpuScUbDt7JekkQPpB7zCYXyhls8/M9htL4kpT6BgWLzlnOHrqnTAKcN
ODeQJvTOs+oz5IfNmPTY8Y3SWDe7MMYWp0KcTGPUFJ/iN8XQjuhGRAh7SuZVB1i2
CrbzWnP11BtwhMQ43RteUaAE0o3HaMbXkSpQ/NeHTDJ7zj51JIQ8LoUeujZR3LFS
0R59qqi6IBy4cbDm8nnw+4v9FhhLqIqql12Ho+Im9mhNoGLvT3mXchTrM217u0x+
ztCd+OooAU62Uq6aaOf8793+TPmJt334d/I4wspOOWN8uuA9YzrOo0CBtOZkjdkH
Fmvqc0I2BA+gml81GXs+2WSph9Ry/2X2O/3RuzYAZ/nevkWZwXeG9dnz4mio2Rfk
rJoYPm7ML791cwoF7xSAo08MUCgp6VvIrA5Xp/rnpjlurMKG2KzeQ2/IbjbCEwsM
aQgh+12JE0d+uSKrMDh1iByrLmhLSbbRJyMeG4nm1hkBht0rX4J5Bz4i/w4rPsNm
QgWvGbirDcmOTOGfJFYbkBUik8BMF60YggZh5pj0RhmHwFNXxIGDCxBnccFPF0nP
eU5iPePM957ZUN/DR0RiLcNwRkA0u0N8/0tNAkKF6jpxZK4fS1Ccp1Mtm+oEcFI3
fWZ/ILIJ61T0FfwcHVkrM2glAKWrLnsFzA09iRXWqXES41s1ee1KDwI+TOtSEjLs
jfw2BDbswxDwp8n9fuLcwlAScC+knr3Udw5vgYkbdLCqNCsI2YFSFtN5RKHNw9Fy
QjNDrCCNPoNZwLwPV/858R9SOoonAdFV4jb9uQigjxg69ci7V7SuW0eGAOQeEY6+
aslbDXs/RZCWj62yOSKyjVaynE01qciw8RUl2sIHvnIIzm5msjxSPA4GH3TBHeH8
b93gThjeVmJn9rxLxDunw2SkWLYJZv99KnmB4GmPLNC2Ry06PqVNhYu/xeoW1GeU
ug3mKJR6POA6yqIVnKhBl8teyJgSg335iGQVcQmrLlEoZplJuoF2Q82yIwDye4vE
XvBQcvqswLZHM8un7h40OLmLGvbT36DhH73W1rXRziYFkCpgaj+W5BCGoIm9wfLH
A0cHp6CbIkZIPEmfGkfGUL7y0d+5QYkcUoZ6ELVCCD8fFeS433OzyhAeIYJn11VE
Gscwi2BqvvD1Zo3l14oW6LyL6FrgEW6yBkz9fNYOVjVpscrCqj8Ec3yM+Nqii7tZ
j0U1y0TypC1x5OuQb4WOzNewvv7wM5stVQjghLCIAgt2CFTkrTs9PVeKHEVXSfVx
4RSfGjACppykbwUZPAiE8RhKHY8TBvvBFyNH2+ReYJgq3V/wiKO230Is2qi8Zt7M
mnaOf4IlH4I7vgN+pY055E3ziZaztHQUaIMXrTyI0vgPLNSYj9mZpvwsZyp53ngI
qNsUmc6b57CiRg6s3x9RsJgLTwaOeirXHCPHMrgX0WYBH6CG0FRICcTgy+nCsGeQ
YhZmgowT4xtIbomMR/VpwL5DKVXEy4KDBjP0UV2epcIv+CsxMCXKn2qsfUcOTakJ
pNeUbMGI8UAQrrQdY/GVKdo3RASUSULwpJwNAv0QICxQJZqJxnQE5UIqMQ+VSSUe
zCIXW7vlzJ5jODEoPcZ2w742uxHUmzjDXCi5IWJFjBka3kv1yq8DyR9odPeJY0nz
tZH5uXK5T2GjO/mhE3eckzvjioAgVk1vUp360uM0eFFaC2FqykSQ/o+DYIvJlOHc
YvsrpCLB/EQZnD//1a8mIk1l4bcJ/WDV4Mhl7lRKelMZgmETIdcTnRHca5InBE57
2Ri6cKlrJjH1IA1p2hG9mR3zRFZQp7jZJ/KOpZvYsDIvnI/vU4lAHcq0xQc+4LmS
y/GtfM2IQ62SjQVv9gwYaO77mUFSTrfEFNZt7FznmyQJctcL2VLpjevrVdLP/b7h
YS+MWVxvrwTmmOfHcf58pFC9QLqboWL/Bt/v66xnH7EjEDB7ql7SIG5OYmbsgnk1
2kePw9d6WwB08rLpEB6y7I2FRkXCKcXDLt1am9nmAh7CTk8Nn8JoDyRQm6pK3TNF
Fg0zMYLrRcnQokN7DJIiBY44GD/KXXH5OfCbOrmys6/0B6EAwM8KBJ3gkx3l4Bp3
i8rafNzag8yOQHM1EL+5hwEFcLopnuVZsU2fw/QkND1LoZbkMPamqfCSCuOG0xo9
oSpHJZIhvDCWE3J1K3wQhR73NrYWt26TnNR1if26rEuXlLxXlqHl2svVUi8qz7Wb
cCVCNhKQtZDKyT+3sCCRx0NdU4ASlV3rkb6B4hlkNuurHp9bl56Kdgy216JKHZ69
IjXZbik4IVfVDJPTdn2aqCRQPj9PPBI+EJgW4qjlnFXIcUpmsPrXr+OVhmDnDmbp
K4ClBFUWvtDVhlfdxl+6LBMY/Iquzth9VWZFVNdKDXPwiuoeApRn8DKzyLUjRP9Y
NKKRy8/Qdcg+isAHHal9JluTIv30VegbNKXX7cSj36Xha4gbx4wHGZAG8fZ+Wb/E
2JOLvHSiP1zM95I7Xce6x077DS+DhhYIOBSUvpXoh9/vRk33OgnyQ5x7h2vU+YD0
Pa+OMdEN/gtjpGJQoWP7nCS0tjYOclvWOrWYlgk7tR4Rt2BEHoVMcv7fqI6ByX4v
6KzVcNvch8+TyzWsh8BWHDTWcmVQC0W6xRJSo1SAWdEZJ+v06xrDUUB2u3clxrKQ
rBXWXlysPPri3Jx3mj6816ycVh8KaT1s0J2DmkCm3hAZUR+M6oqUq44LiP/gpIPS
aWaFRIWrZ/zd+CqmPBCAOFwr8hzHvsgD1UThBBZZSI4LYnATRjTA228htYdYXR1+
HM+WDmXkhoH9hb8WggGN8uBSZvrikE3SpQNb1jWTikjsiZXrCsNV6KEd31RAVCnm
xF5wYuG4ejiU4DTYYkr3tfugFmFjETPj0J6JyZfWWKDG7Axo+7egNT4bITmxbNd5
GftN6M+rHdkpJViCEsdfvTf5JjE/yaag2wvTHL2qx1XZaMtI1VRuTtYQh3I62VAW
vbLDtElcmsanoykLXJ3YD7OZ0uKE6AJTTK6w2ZUnINX6tg+Hd827qpADiTb0nf5B
qPEtix1/J5Ex53mhfxIDvfECqsCq17B72eUsOCcdWu/BaZ7yJi3pYg5OwHCtZEk/
JhgwNgA8PB/SnP1AaPeXt6VvwSbaoKhTDynX65JlWtNV2Q4voNJMbN0G5B2G3eHb
QSbHZrdJEa9xnEuOfWtvGPITjMxqt/82yAFjP2EJlR9JJqbuWGmP8KjmaiuIJj9d
dRJ0qpoAMNEK2SbOdKEGjY404/VcJAZQ0NJEUdeXdBj/AVEGHu9Eotp4xPVYcT0q
iezEprkRqxxMBKIXJlGbtwnY8OSIjHv7uzWsQuJ8CIEYbVwD+Vh9vkX7Ge0zsfEC
8WUeyXDYPnLUcVEGn1uvgi+UYxojvh/g0Jqw18NiZ6Jp378w684af24BR1vxdI28
EY6qv4rsZDkhZXSBwMKw0B6uebOuE4X9YmvNCqiTvoSi5HgsvOEiqvK7zFrX/iOx
q1oqEQCaoKMV4AqdV5vPG6bXfMljga1ckr7t9jBoh+AJX5pyXFsTZ5AglpjOrR2m
wvmhRXLhj0VWGR47b38RONzqiaZX+NSW2/QS3qc/OQyPYTDk7oma0d5qd6Dasadw
T7lfojq7c+NSOxoqciWxiWO/6XK+nFxh2cdfj7KErC8WJLoj3TkNAVK0bKRVBaiz
6psJOrQvcSH0XNIE5Mq+SMgrfG0lxGiohfr3PBJkB4awCxvBqz3kPyRTSBGwfXF/
Wli06vldeRBiMieCfpomcdKlLA6+9gpJ1YikxOebg/TRi1CcaE0Hb4xJMWIkVhsx
fPrQRaCAEE/UKb8Shgx89gdNLdhrZkGY7eZEWwsHo5Cfq1S3p5MvCx6KE8DTBZMm
59ey74bsu1Iq9nSkb7W1msLW07UnjWzXivUC5FU8n26aofoBSKlpTTW+emUpDvqS
m1VMXrPKXkIm+Zs3QUqw58CCnhY6wOMrkv69XFQ10H2A2XzVcPfewcF8tt19J34C
nWSAwGSoq1eDeDO08y57ZBf1uAHzQM/x1zAk0turMU+DB75t0H8F10UhO/LL2U+M
3PPf58w2eNdC02TBvPSB4HZ72DwAqpaesIQKTPiFwH5DrO8w9OwnUh0zeHRpGrON
UB3NnOcU+IpHEAoEgp8JR2S4kEYot1B713hVUqs8AYPWrxxRwhzAV0DI7ctjvXny
j55FQL/dOigwECT/ISAkp32dmfJPac7f/+iG2Baa58VaT/q1/j1AVDBloczreWt6
+kABDUqKv8G8QXh9BhRgKgw60OO1Tt/unoAFEhOpQK3wGoRBQuyzCAUnEba0MtBh
YIR2Nwl1gdHWHC5But/FgBKOuxdgEMgcZPn6DgDsVCmHP6N65k7Nc3TUzA0Kqb7M
Wh3ObBwHzoS52limC8Mwfn3mCwF1lJ5qVFozEyqfpiI1/bpGsC7CtPa5B6GOFcJw
hutpPtNW6t/Dm6bLgd7vAseid8B/JMeu04TbSvGhj+hB09//6i8vXlZQotnCKe7u
PfoAoI8+2DwevZG3ISUJ039/09pU8Rwq7pb9Wa3dNk08u9M/uqp0sEILgyxYIaal
+9TYDRjFjX4P3PLV3fXfRE9KISFTnStKgyGDglNg4MBizRmcRBqztjRFYfMxXLzy
N0hy27B+DEDWNnSlrgjwcsxrxBwguQPukZh2dKsdfb2pOIJ+esh4re342u0LmZwS
xfRS09F6YFsGjkYsyKa/b/8QtUt/l84fehCP+sj/RQuX5j8y+EhKMKYldFuGFKOR
TEyUU1GKqebFAZHPJ9iNVG6LPce//FrH0TPEGZVju0yCyr9mF2iCardhi2nVe6GM
7HFsKMxTj5DJ7ZjxnQj32MaVMNBZFeLBprc6sD5Eg+Z3v83izJNWad3OlSgvaSAl
TN/R0cWBD/KaxcTjgX7gInlHqkZZbRPxyaQc+w9N051+WqkiyLWNcElsnMHZ5Yry
Sh9p3MpAilgxqncO7sWVQKbF0j4Fq9Ex/o/8fGmYQu8xsRyTgA8mzq/mO4Y84CgT
nfO+7TfMgcw2cibkN+MvjWgUHOMDzlAzQcstJsKEt3LNo/RinV3s4/MchwZFJem3
GGNO03EyKfY7y5uNO9+2cHUqX6X2o4JCUKzThCyIkhy5hfOqhWne8DrhAb+OTjdS
C7ixAU1y8tm89+vxCAa4BrGMlbB/QOUxlbvQY7uxmG+63MOK1Afti/8WvLMQnIPX
HqOpQ8g1uROhsW0XyYIFdjk7og70HSBgFZRKxuFo5S7pUeymT16p42wxbEMFzxlb
hEnEoXw+RoIEmVnF9dT5DikVcqWDFXZv2wzthGcOf9T2kO6hXUlRjtSzi1m1VKzI
IeMEuIbjtNkY4//3y7ZQ95TjpcKy0tsenlMjUNfbiMhcovSFljEbQ+k0+eRrIak5
AAueH2Z9onzYV3xBfw7GwIB8uFBTseDY9nBubSBm+kqDNRxdw0RGpjCVOrx8yY2A
jn6RCGX104TcWKcTMxlDI3wA8ecmp5Txfb2LWdRUqQQ23fPUlypsk/OQ/DBwyccP
gEJIJjB9hE9S5XRtTsymMs8GPfcqdkKfZQVYqK4MTFnaTB7Db7QwqEam6nYozopH
6AdmQHnbSmS/FF2gYFmi+2ZjmqBme15u5+7/aZZBvDLKRIUjf0Fx/dri7tuAHG8b
tVX7eqCBmdEP/yKS4S4G6XzqZ0Qj3UUEuZYh3qFwu1VVAPhQZ2YkqhcbtxljlZy/
J5T7uZx/51RfNcMx4fHypA+0k07NXrmoZYbG9EeC6gkgslceMOu6CG1wbxRQ7DDm
EH6109HVEpoFik9Ozrh+2BNNfq5KX9+8WmMP3pV05xqdlajunS+DmOMHW8nV52IV
9Pw/0LzY7IxyfFWsHdqZK1TnhD+ZSFe+8WKn0ZrHvLUaChhr0yJRqMG7RANa4Cyh
VhBr+wLI+bxEGIxj76rR3j8JydajrV/omLD4cHRgJ6S6Gy4WphHwtBOEwx8qD3s6
9MX9eW2NV2U8VxXm3eHfR3sC6cXDiQeviBlzbHWJHHxGhCsLSQzRJ2PhQeh+L3D+
oWsZEU188m4APHoH93JNS/MIUX1SAUq/DMfDXgwO37iUMYWHoIKP2emHNhR2IKwz
HxqWZNIV+OmZiK7UEGQktquVmhQkfe+bYHEMUyvH6Bag+c+w17h78UaOYS6rJ/xI
OmFli+7tpUdtUaNuuKxRoFzNwsKEZLP3GmvyWWWTpUtG5p9eWw1dWNBFruKXCK1A
uMBTuuu7nuY4UI/zJ0H1JGZxjxuJNE0lXaFcd6aCSweXptWuM7y0ZvA0OgJ188S2
1XrMtXGbFOpxIZUx3hGjkYX8IsruswVAK6dSbPB47XR8ze2xx/VvBNxyl8te6gRl
ji3q+Xpz7paLd4meVEkxn3rw0fspwacyJiX4lhvlLDX3mcJEbD9UtuGeRkdH4sel
GXjT5x02i+9X9NrsBKMqmp7os62ebXdsOC+ZfsbusdhXXBCRXPihN0JwwPh+m2l0
a6llLyPMGuwcHJ5Jp59u0mzokcb7lVnrL8ltiua4KSF1EBe2K8mK8oRbR2nzAkkE
3pHt1SP94PyiiDtmSYq/mqLyrSy8lRZE3WKQtXtB/21WwmfPAYSq+EZTMqeh0oV0
bB32PKoJLrZQ3SK9x1bQhsn7v9v/3V1swBwoE+tDO9WbgZP2Cb1Vdsaun8fndSTb
CJiBkQOmY9umMywsoBlo7Io5zrtejJj/bVbd5RTXyQt7tFBo4ffL0Wf2riP7VpvK
509AWsxt/F5WNC59iXEWQQNXlZ3yj5EnpsieI4OCAKxF3tcmAveFw6/X7rVsk03u
vK59Ag+FpGUMHiYb/rgCFD3eVNFi29Acca9c2TndKpGzDg6EGrcWbEGfFcfD3n6q
nMzx2YCct/iZhB2+k7ncTuCrYDzBXwuwbybH4gXmFRCLOVIu7SlIreO5BFG6UpQs
waofIntn3QGcwC49LK/l0IENSqC56SCvsHZUy7sJe7BHSbkJTTwaGcXyoLAOQBtU
6IkWfZXgEdql+P93YOeOFSJBVFriKrSbr6HlTUyX9Cbonb6oXICoxjQtOLRU08d2
VT/Q85BMGY88HXnAIvEidLg2+ucnqbHXqyLzEmABlv6vgWjDrCLYcNR6P3vBl9iC
fCvlxlULlO1RSizzmswKl1smD6ORacGuWZXYYBkAIxQSJv860tWboDrhSoS3O2KM
S6AfA3MQ/pYREuldyZgEj3SuWyzEeLyRjqQeDDCwK140wB+fR7CK/ZA1j6MvXuPa
HN/e1kB26h8LOtYJ832evo+jFbi8NmKN1ArDQ3pN5m2ib4htY3Bmr24d6hr/lyNK
aqYhHlaZ6oa0Q8caU2xosoED2G7lGAXlUmsq5jqTJ8BxpOzM2vrHMIqq4TiDVHOm
IgYkxQtviEWLfkZuNOvg+zhmNBSSy4fuzMKCfKRqdquZ0GWMxgIyghMxNlDTQbSE
lqt+NNDtwLs/JXzdkPDa5Vmwt2uhTSm3CFVxKfoK1mJGoj+XmUzU071Fc3sUJtAK
BtOczHRhpEiYRFs0RtufnHkWKqfyx2PyfAvBTmNBH8njT8TUW2VC4MvGn6a8fCFV
upE9WYqf8X2HNVS2LnTQw23vReuRHKpO62uFmw9CwhE1pb5Kp8ngNKA8ITOWxfOP
qFGd17wxErwihdHLqBTy7xpDOrYeM7YHQZ1FXlsmZr9CHzyptxnggc9pUfOttjel
EHTbrTC2ILnDfYb0udSWTsrvWFIbsfUCO1pPvYK3WGezo60KC8Dpp+iInFcuZ1JO
NO3gKouWgIVz9vhOU8Z+yk+urtBRUU8gTQRwnuOMLOrIIu7w5rIv09KbrER0Plqn
QcaLk2gBbud7aZ33D6Y1FUFri6sETplwWN9g7I1gq2P/hijBfXTk4AbsvUx1jfD7
vNOFFqzIAAtI6NOXlJ4ZWB43PtHTEQru6N9loFX7nukVXX1lurdApyvfluIHOFiB
IEu1Y74sFw2RBWsbiIZ7YFzn7c13E0zaHfj53yTYTuzRtqmJbSuw/1y6Q9jZCbWJ
NcTVGE3Oungzc5rw8AE9mM6Ua7/cRtMQ0naWyefFcaHAtAGulgYpxxFrCkh/RUVI
66vjNzcs1gCzamZ8vYPFTOHQQXEhQwDa0GhimNg3Bayky63ekXoxjeGg4+S87iPh
Qp5aRTqTCBjC/LKxc+fok5rhDXZix7PimCnXqsxrdZL7VjygBCWYUvGE0uaWVsH/
tCTBFC0NvNIciqmj4Ydw1V1WtfHJOvcV5Gb8c3M+Y4CYZw/ETgV6+Y7mAd21gY3v
3IKWZ2/Z06Ki0Fq79VyNxVvvt6Aay4XFoBXDWACzI9j2qi8cBX6JTWGfBRf+HXc0
cbQYl9IxU99Qe2IktMu5X2j+2hA/vxe1/8d7JESiNXswtH6hBv95ayHeYAaArjwI
DIXoblYq3xjc4Cw+NLfsPtJTEN9SQjwYMCy0i/cQFAPFz8ydJZLzuN6y8ftRzYwO
rvaMe7IA+WpHbaB5NcDBKhrcWy+1k7BF1agsoMFsZdukYMohlKqBtlonHaGmYqKm
bVvlrNDZk4HkOigTpx4r3ZgRB17EDt4kuGyHJwZhdWx45Lr8DiGYmDw0nSAozz9+
qmXGsrKOvP2f4ovEtfIURb/MBb0X7RSavM+CD52FZvYUT2R+7wQiXOnorWUsgDuH
qpvqHelzSNdpzeHJ/n/429lG0hN4NuuEKNAhAlKzAiq4q7bUKz2QEQJ2RD3U/GFP
dhtlVZdWyjEiWiF5CH0ke5hD6RvjSigHReUCxm5waqI9M//8pZzwkUh9iK9Y40Wv
iEoP1CgGSnKErayYZxhnzapZdI16j7AlPzSMZEixghqNGz5gxCOBKKUMsWKtC8Ow
9oHwJ8MywZcPzNBt1o4XtsPPwPgGPitBAJn6Ob43dGa2LEv7aZPydI5MhCsigAUi
ChuUb7K/AbhtSO/4MJF5mV+HQzl3A//zjK5vzkbPl4bnje9DBbR5BVGb50ivUqQ8
WHavxmwYBDyzm8PhH17PoB6OQ1pBD+Nb66WA7jlDNLha634Y17T+PuhNKUN/p62D
spl4G3KKB5qQpUZDJavl0SoSBwZEI/ND/1bXnzIwm9ai6ZGfDBbYTtkAGZIwnB+S
Ppg42uDfN0M9LNG7Wf+Gxpea4Y+Y+3U5UH640u0140sRJeUM8pZ4q4ObSAv4t3ry
bAr/DNsy6IgVzQOnkCGZjkbin5iy84jEqGH5QlK+/UC/pwSC5zinfhRyXWAyROQw
5mwhorIAngMSuo6pHP/XSvB3M1G03lXf4aWY5DB+k92bCQt0J8AuBi+BNYNhtt+w
Q/JivLp3QrTn7nl2lwAyURSuI/x25yjE/IFAWcqmg0wZ87k2WfRSs58Y0dfhOrEq
E6XkOJoY35vAl9JNNNUW2vANw09AaQBX3uKs+KXhepIbE1flejnKhzOrMDQVthWb
Eb4zT8zgk8JKzFcVC34iMl/Mc2UuN+v6C/qoz0mRDN66IhlcAxDm7ACAakHFsCIk
RsCnPpsjUYV9grHwttLkSvdJ/W4U18QhM/oMfjd58nm0s1udU8phuVeWY/WfLoGF
7Vt4cGQbHhsUSxNDo/7iX2wXZmIhjYm0J4YS0UZqdAqXWwUehIpW2IiOPvVjsYQF
aEkbcUybDXlXc7YQMTC5gHnUO1u/1zikgupQyN9DZKeazKNPuBuyLT1mTVhvq4cq
2Y4avnSNhKtNVLJZpE8ZcAZoMBsrrkJcOkBsqL6x7htq/EHrSK/8TicpOm2CXB0X
zNlk4f6YFgAcLYAKQ6qgOl4rK10DsUvs5R5UuCvjYdiYBKin6AL7jCOr4IqAzofq
l1XHIi88/oTHhC7JZILPdu4OF7v0a32mlyFFc9csyC4XiFPirU7Ezmghh1CG10rt
pHiuzoxP9ZQDW6BIv2Xe860S0pXvuMGEt2wAeRIfafFt3JkgqB8zkzePFxpEXLxZ
KuBnd7E8csz91BRMfHMOJGTIySXT1xbYCFwa9x1E9F79IkWdmaDvVTy+FS96shmA
2gnyc+l9QPl6TrdGjZk9/QZt1FWb88hTAAw8E05cN3paEwOqC4YsJl1dxnv/oUBy
USiTYM9GEB7LEdxQEazgzMmziJ1fC13a5yrDNxrF77Z9VFjYFnrpcxRvXq3tiEEu
NEt95usgTXLZMrzHL0ggMOL/2ZeXT1qoO0ZpkFwDLupBxy3FgC/jtn71yEtTL4/1
eQeWvGekshO4e4GDH6puRBPPea+SYVTU1g2jmz6FX3dLjggpXmckrLXCxKT8O7Mt
Y+UTEt7AEd/HLAA7A/nMnEOmjb1IxExZMQEyEVNcFaNTMNjAsTAtkt/yQd0hDy1y
Cl98a/mQnKBvJ97vd22SUxqGhNyx38aRWq+eD6iuwVLD0pQ+Yn2l/ME1Ys+pQe0B
qoNTL/0v3iwcGGs4JkQyoqnSVqitsVFx3PEL89PqVqcenkPAu0UZv1p1ymg4ek5S
XInPwZqrYMJkD1tYAb5TdruK8mp1EKzHrgrzgEkHB9LfZXWl2DmgGrZ7BJAy15Bk
8uegq/6guJ+BEsxXqfEH+ymjxketZoDN9fUb/WgetBkrYYO83Ts3mIUPW9g6iYGW
q7dAnHaxabujuvNAuVoPWdIRiY2yCDJ0C2mqKAqBId76GannZRYnrtvOn3wrw1i9
lfpe7xq3CMU3VblfyYElhWEjhtA58MXhQrarJDZ5b4kpxG2LtQthFTgy2khhzvdl
S2fkmkDOXjnac28sxPAmQlNMRSTLYQWYae0uVLQTqjnQThUjX4StAReWAolXbgbJ
S7EmALz5JQ+ARhiDwr4ZRxe4TeOjlOHQuQ4kKEPQCTCXDZ2/fwU+CbOu6ICvhXwc
msAvFKue0eR8KEww6oGUDGbTzd253/Saw4HIJbUdWCAuRGYfu4ECv8RrPp3Rlf4F
vSXPaA6OE2Hrt1qTit9wQulTVy0cftpeae/h+hH9GZ9beU0kIPhV33FMuPm6Iskx
H3+ulK2bQH61DqSdcRJSXqKz8nTYRSbu64qwYMs4yCDQ2bkio9KWECMCFYp8ngKr
elK6u0TBhJ/+y2N0rk2dhYN0mEsSBmGOq/Ylbg5mb7XaGtJ+65ktuG0og4/TCIfq
GhxvvPEPK9j23YciQQtluiZZy801tr2di4nys8FEW8Nep0IqODW9hd/9h/5ScXbZ
jm+7V45CNfZw/IAYa4ZiEM6F48HChBoMukhPYhNOGbEiQaBHbWFsWA5FKXpfSVcG
PDMdbuCZWWfMc3b2jVCrye6KJw2AiIHQ8fMdfn5wPRSngo3ZDzu03W1d/O9JcXEz
1b0uF0275Kr0ugh8Qpwgzq3Es7T9fXCxNS0fNOq2fTxLU0F7/+7Tvs52LffdFLIq
Q0SGKteRo1b7fpIAMYJ4/7uBxR2nCOaza3kRnu8ksfqVixYVjoUf5FGaUpxprWrN
hkoisgcq4uvX5+3yF3VtG0tCtcs/98Wk6LokGkm2gN6xaa2Lv2/FwZDAwxl3KInx
x5kN0e5QsgEHaXme2/OlEptJIbdUsJVqMCgxf8EnaALFZna//5BSfFLTapS5hmSw
GmqlDz2pmx4vJf2AWsFWGqWOaKTDM1t9TmZpLpJ5R7D7A5mq3eDm5Y8FF3/S/37K
naYEdd0MIFmAH5REg7Yulf6i5V/fD/IunX6e6Eq7zrjU2je4Lhy6yfkTl/H1JS+Q
W/7MPOrR889sE3Sd6AHw/kdjlBmHsxDvqYcPqZVKGgwwW9+LGeVgXv+P3UpAe1kN
4+dVF9CE/QEt6UmcjjN83WVKEbLp5pNutajB/5Gpk0f2qOFc+6hB398ZryC3G1XI
1vaYAm4eL+rRLMJs1WXTryRsYRiMOuhg4FT2EBZoT+XHsvxp4Rdw00JBlZQD1LSS
ujDiXhB/PVCdatHN6wICGcYN9bryduqFLAhzyqP8n6ix0Kq4xoHTMZJEq7IROZje
XEOd3SMQc0tEi3AyPMMe95681uqkZeB32EHg5pQOOfaJK2q5GiH0SnYfziIpZzr3
G224KwUNtudSVBWuhjBM4+8CqH1MGvG0joIKrrMjJ/YgewqzuBlRtEIfFKhmwNPG
Yh8bXfjpVxnYgY2s2+QmVVzEM4jiHHRFMowWG7HCa9Ygr6+njQ3AXV0EbeN4XSno
Ym0k1Bm3bq+9ON50RqnhxCNbr4djzmW9HiuLc1hFXSEWZ9le2iEPVvPDNSAfo/dJ
aUgQhNDYPfefgu9Yqy770mecvNV3Rh+CgJChh62diBTZCKsKBohfggM9i9ulagam
2TKK8+IYZgbv/KCFLHKotRmDeb8Ddqw+N7WxFDaF2CQXABLIIkNlHA80ndy//kEj
nhB9Ik7i6/Pjazm/MBFnCmp21XI4EarfnJr2UUxR2o1I3hw0c2BWu+6J/mDxL1xm
GSpHRl8tAas7+LASuJAyF35OoyyZz21nOT5lgohnhgmjSlgoFvZFRbpdblUExaT1
9I5jbmxUfjzxr+OWpv6GBF1PTSeDXZkfrFAnZspEogh5ySShDV9jCqtoZBhqMVFO
XFRsbdAJbPi2OyYd0QeX0Jh4II9TY+Yn/c4F78m9tJCHa4JuVs3c9zYE1tKYLrxU
+R+DX9dt0Ue4t76VS6K8Pl+tiYxJPrCHQMbF55ixqW7/23d5+Scr/BOtN+ZR6tVW
10IdrPJ9MUPU/K8xUtezRRoimSqPo6ZasMnvv8aRCxQF9/eAJLULGSAoXvQ+xHA0
kTyUd5ChzFeHCGKCRn4iSBgLCt1uL/JNWSDJngRKiFHEe3ysz1VgSg8B9ftThJSs
hw+FnVtSaNToeLDZYK6fWDqef7Jh8V5VIWCKtmNllDW+NWgZ3A7m5UhaL1PCSxbC
ChYyC0iGa4Hr1lTOop+31oeY74Hy1a155MuBOKzAeKr3DdttmUxJ41iH3tHvmNGw
yJWvDBN7CG6v27b12ccVcfL9vF/bpF63cSu3pVE8WLxFjk99d0fWlODki/aygCQ3
3h4aT5DZopsUwxDAdmp0cMB5Sxgibc6eJsIkfpc2ggVScCWCTXHaBts1KEAsH+qQ
xXavhhQnNS/B+aWMduvFElH+mkM82A6HkaEVVd4kaeRWmHq/dh17IBeHzXR7pNLr
Pkqjzife0cDNrEiIi2hlvo6AnxivJPiIiOxlB5mpx8J/hNspjV7W8z+RYr2oU6gk
qO+WINje/C9MS9WBkKLAh+nKnqRCAMwSJ2JBg/n5rD47xmX2qQwfYE4tyhXh9jVe
72kVCI6gMqwXUnSdTKQQtZOK9LlCVBxPb4a++jCcK1kaZIzT8bOv3Qp23Wxfubq7
qQkfw9WyS3apqFhDNfvT1Ao+PBEQsIYynUWPWyXm7/pvsaLZm/sMPubo9Z7b7b7j
vLww/id0jebtAk+4v2xc64sk7YWtcNLs+lcdk8mk5Q13Yqt8SErbOzFaSBzzGWRz
g2gPDNal828IJ7uzlbfHEpDItWAH9FnL4h7rbRNltbcHezsNd5up23tyiYNeync6
Nulbq/zUl+XSenh83Wzj/nTpD9mACxhLn540elm0ddqOi2V7Lu2bq7QWW2jVv9Yi
XxLgQbAtcq67wi/BavXpS8XVWay80okLxicsVQ9syQvo+ANJZJGDyaOmrKHYONPV
zL1okTM6Kf2qEGCmbwmbmxjnOb0jRvy5Y/8jEPcaJtNwKDei37DSQypOD6ZcYdee
qQMsO2Q31nQEwl2EScqf01BhHk6veeSB7dZVUD2DA9FhM6yYSqWcdUTxysefVKDI
QJAxytVyXfGCsbxXkE0lPJAaKK9j1269I6o3KPlygT3cF1K143ZWRyqdmZOI3JZg
kIHHgvFEj3VQzqlNzuWdTHBXR18y9TOmuyW17hogrEYJZ5iL7ogp03Syy4YLlhlj
QatsFkZWCdwXctTkvV4EkGzaxA9zJr5gr71XkI/NbflbqTMpN+mr1L5xdtv8Zq68
Y7HAQAs8FYBdwERe6twbFmyWx0iWEOQl4nHS9Mh9NuZMmieREvOm2ncQykkRXpu/
na0pZrlS6Ra18VBQy2t9ihD4tIi7e8+0XE9fo4AgZM12uLTKgBcqm/i0ZTZgdffr
VC5HUpxIiEoD4jFC9P9W/5fee0d3aBrqz/QRKNiG8hpgciqbsw/2QRk7IyLvg39a
VRthRLeMB9Bii5Eh9S/juYRORjqfoBkgNSx4mDmKnh4TfZWrkqzfntt/1YT1gOi2
h6rUo11I9WFPgIzienMeSswoWunXkwkbIGytnVVGnj5bNmXaxZv5Uqwma6kXO+sq
N0wxERI2h+L5ZrG7n2a1mNmEtfXikUm3+jt9WUK/Y4xgZQcOc33rfvKH29NiUq2N
4zZaNX2PRVU64WgaY1RiJFTi7L6alPycAdkSyWF53Mmss/lvSOAvFgwWgKOl2IlJ
NLQm4yKOrZJy7VHwN6R/EIzV96vh3H2h3PktfAySXZbgS6tRFu/rrnA4OST3T33q
QvIsSMEQe7YnmAU9qlshrTwcQRkDAkGjpjMHXEeXaQM+hqqshePluBG1c8iCvvWv
NkgknmIIPIvMmpNnPtRkpGTFZtcogaWe6CjOOKbb5cD+uKOKGbxN/9FmssveEJsK
oyb1F/NoO+ATF3rcb1U4Z406HH6OnrG1/eJfmnAuF1bpzjd++K6yd0ViLCOJaXsi
YmDGy+ORNd3RYexTfmxfsE4BKWAoLic+QpFPnwTV4h4AcoSoLrlIR+g7xrcQ+dEj
agn5Ie7ZyxNIiTWdEjRHQYmU/20kCGlTMrzRSxAaZny53kaLFlSLS1jDhPSO1FCC
ZcFEH7cyZssA01lZBe/veb2Jd+OuUc/MXtdbPCfQWcDikQpOs7JNX7mU1rW4sZhG
ObfofkJ4iUMEz9RVK4BYPFLNBY+8Qx1clLFf8Y+GJtE+9+rF9VRx/GQNMl2J65Pm
bcsX9DV3l2edyDI8amqO46JUsE7XRhX70O+JYt4dSzsdRC7lOm4nUTzxjNnMVsEs
1N9ZC13xFEVnYXyNUP0fkpLWu1gqbF4EBWXyhfUGeid+YOR8tE/4vLVb8YIOR37u
X0ld18CUBg3llMYixoYbOddn95DBiopARy5CqNUNAm1aDpzmw5Ys/PZP0zVafeli
6Ijf2bNR8OjVFjLiwtOjzVan9DcSbiaf+XkCS+ksQc08D5m5rnqGxXdROkBNph0r
D2RhphnfoZEPqkv+ADO557mcOdDdQbqAGw47u0FWduuf6bco9hRwQwrmXMcSVHpG
GLnxGdeEalrXBk6BaWRgjyOl+ySVcAFX77yiIdbih+Wphg6VAadUYVXJtNPclxXA
Wv0SorjRFyJZC+qpi6KeRJVf6a0AX5VPY2fb3u0qnDnOJyiAcy4Pwktp417dooLn
RTLFWgwEi1T5BTAIXaeWfbQVOFgJ+BEYx/zO6rMWm8T5YXCJS8e3O+bb6VifMu1t
R6h+Ksn9TSeqiFlRs+P4DehKMZFQOHl5hrhe9y3tdRGbmduUn1a+MG41ftPAdpaL
JqYN03HlYlRXmeQi4f2wQ8isFqUB1UM3KU7Q4xMbh6NOT2upeZQaZLis31Y3QXxj
C2uoXpVz0fw7CnWrcGbfb9gF3dgIVDWojHmbwyjlDH4iooRA0d4rcQ+uUMgbbZY3
i8DgqlEvbH8o344uXqTe+IvHSJj93LgDOF5ZFfEOm7bce2jqMeMY3NLv0uG0iYRf
eN2XZ/yGYEOUg5YiTb+DmmX7eQgcYWlPm23nYzThyGSiV7HwrRp/ifwmAul8xzA6
PZ5k8ryTU+Uqu4EMjbQebTITrvEM0jo7QhboqCt9u60FhfGGSmsn8JgyKN7Y6vEP
5pT9GuWasEg/1Q88famRDks5Al+ihB+Zy9FOm1GXwT5Jk9EKrNZIzqmZySSqWRzX
9cZzDdh3tL/dKQE/yM0csIf2Z1CPgqPjLyvUzvU905VrpFmkcHdeb6wtSuoqePzC
cngtKnbSOBAI9NUK/U3jwkX2CaBT9I5ByD+IVNV6rPe+epD2rmaUcMq4ishboYqI
d5JQx5FYe1buM4w8JlbI7gw63VilJdC4wcPNXMFLTMR6QVhMn7jfr04z4ZQtVGQ/
AOzNQ7wDmGJHoX8ZueadfNB3dK8zK8Yi9gqPTUdu6bWyaSIcWOdS1IP4q6fLhn4Y
W4D3SA+4WOefU6gZmJ67zJKpewtmSYDzPRCHEczfsX+1EqKJAAKbe6nKAg7MeU+r
nr2qt2Jt8Rj5PqjGfes8P2LP74A8iZeyaPKXUIBV+P/G35XCflNtGbRGSWnQEOnw
66Tz0YyCCB8fbHpiRl6GkEfSsMU0ZKR5HNyOr4x3UnnJqCdkamG97qM9kVTxxNcb
8Tp+zsNn4nMQk8FAZIW95AVPc2r0kkn2NcPT5LXnB7V7eIb+E5RSXbKf7CFV5piw
QZI4kgETl7LfBjimugSrE4yh3HOXtEjx5JfyDCUEdiGUjulM6UOCzghUU0+KM70A
Czi6sWdPpyqtQm2CPNREiYHYzY5y3k4BLbdlIryO3yG75DCSdZnJoDJ+n5s0BeT2
Ejyn409W7lqpUiL6UDWUEyUf0j1EFVDNO3G4Gb3eynlZrPHJ1XqumuAxlSdFybnw
9wEufCHBXaKO63V4xiUPZehY5nkAW/8QOqzF3FL/6l20KRPTsmm1sR9C+NWgwagh
3utpUWXcyQIV3P1G9eHNxSAMHU3Eax1QsvjS2HUNgvRge7QBLxAEEM+uQ9J08cRz
aiuJinoBg+aWxMfa04CcFay9wQGwbciP3c+trS93VZBH2Dyxn3y4AUWolkJXPRUC
ScAVo+PrkgL+++Tr60yVjjAactF6CAqA5UNm0m1qnUKEoXVX0+bTW11ZjOt1fi1t
dTU2lygr6NWfHSLp0yrtEOVL9Xm9j0GDYP9SGYUP97ucjL3H73033vxNe/HU5UI1
GOVug4jO3q9ShGSKlKt4DU5nxBvoAmT9OlGSOrJ3RnMpLEXFPFtIsAuw3H/iEkpK
nH8PivCL+BJ+F5L+ZEHnGzM2SgONTO6cZT5tc37s0Oun0aUqN9LZXaPBlwHIM1c9
RJ79NIAJrbOffWr3mFyuWd01240i+FJcSzdO6+kgzod8SQ2rEpox1FX8JuLh4sjw
tgEKmFRZrWKwfs4JSvi3INuLfFfGfr/h8gXpH5JZo6veVs4K+oOI/1YtH6jx4c6F
u7IO4M8GBX+BBBEuXturCjDHG8ODrC9UeaN03bZfH/h6I1DOtsw1AlQedtaTlTT8
T7LfmplqzCp7VX9Z4dwgZcw1Qiebdlmb6ZcselIX21xNFzIAGUSnwt1QRF8OlMnC
TfKvCiCks+6MB6NSzR1vg66BS1zugoF1PhuM6As8gRd4hdiZ91fdqxaWRPK1iWcr
U0DGrFZ+S54RFl0RfeMjavImcJpI1Ww0LJXN/KMqf5+tdslbaEYgrvg0rnJh7yho
OmdLP1nMGOPHjo5m+sKenyoRpfgtUv7KzIydoBMEoRz72vQwZOGfuAnyGfopAYwb
oREcZ9mIWZzxdJgPbBDDsO2I0XhqPPP4pO7vUXwjk5rz8LHKvekurPIiLt4zUSE6
t7oPTEkmggMlprwYP2fHBxt+wd7qtRyklzlyIdzNifEjT9d3D6GndoTe/HLCgflR
zIU2qfkN5NdBAyXSCkliCUwzs8YyO8EwvM3dBxOBw6TSI7P/OZGJMm5bxSlTQGRq
8aJv0Kk3gnZjTIG+l/feJX8OA3APs24+c0OY0aodQMzCsOVVR1XNzfZgFr3aVEQw
Fz7oJceyQnRCIolrFTrNyO9KDd0q1wq1ErfKITVcaQkZ/SyJszLQ+icOg95Exo7T
6dbOtpz93UZez5PZHXwT8n55vj7zBB0pwCBoV03NGdT+2HJzNqW4vfs5r3NDx4ln
evlkh7AnZr/hfjqDJHV1Fkm6uzR7mtHYrcXN9I8Jh8qUDggZnzbs8/cGQQxuDP3u
G4SAshpkDShwwb8JcJPRJ0jBGGgFYTlO8uoKzKlMlLLf619VUS7+rpr6sG2ZOuoB
7FIN+dnTIiNDTFt2r56favPImP6cxPJ9KNoyjhv4d9B213XAY+b/GHhx5flhUnm5
KK8wMKEcMWy26OZoK15otbmHyWx7X9Jf6d/UMP/YV6PJLYd+M1zGS99mbOfTKPC7
UwOAHtX3GahZRPk/jUVOIcSv/GGlXGC8dvlmbKCAJE4u9AKof9+y98dSSk2kD3g7
/ruqHt+/9wHxc2F46HL0KMwV5x6DLrz4c7iz2wbEKv0jqC5w7Q/OGFSOCSEn1Ohx
wlBiWGYZYrRY0CH7gM53i/UVJoh9B1+DHfbf37+cFPIy7TF52pG12ny44WhJsjRt
5diHmg4RJnR0e7EHSsQlqYHcxjFZsDzbBbmrORZh1rpwtUy/9Njo38CUunonkj9I
PHLhYEnmB14K4+aZPQFaAEzAYksTBlsy5ckMZHqHGOJTT2P1hOX9QvCIggUs6kHC
BjJFBVyXNV2c5sszF/aX7+z86i+3XX5X8wlTYy7QPiXb8d0v+VmNpAb6hRJzNn8q
RKcw0SF+KS15u/es/I2+ffEiuhCFSPONHmOz1+P07DHj7wQU/748iQsnTyiv/U+f
345Kn03ZL5q7TdwmxjEBxqHROLxaPg6IcIzVtv4q2nlLpcb/B+mpPVGafqMqQvvo
tGuBUICo9yCJHwCiYZr5DqSs5yqApc3Rj7RGUnAPAApaIDYAHZdqukSUk7Mi1Ic5
7alcE2piHrX+nxzDLFMNZ57hTW00Ub4h+/RKRt2ZXtCNtfR4M0tTL1cJhUU5r8Rk
S6vZC+I+aBd1u6DKfNme3BijNZcbc7AZJLJEQg4CWq3kwO4Jbq+JidCkmtttuL8p
VfSuBsBnk+/uti24TSeZ3WJe5nxIO7hdMP38tDKN+XZ8PsdKBoqcQJpsV58BuijC
V1Ev21GIt2QN/Aa5pMsd2DgvxANpjyT2/E4Qwb5LBpQToVZWdVhNjzJ0+s/xh23q
P8HYdBJBUDJaKLXQtvW5BXqD1dxca7v2lP+FQLgeSMaDucQZ4RZk4kawICUCb00P
W36WBgO+w4EUb0kFZ0s9MNS7pEuDug4tD1e394LNNHwQcGvMYeCC4UVMXP2mFLms
PFndHcMS3yIHgBboUXP6LivxQaDUdQRNxceNxEzb8U6zVeYlF+cY4CsCpvKJ6eIb
aA7v+gq/n5QO1cu1MoNuKt8fgqxTXIaBFIETOUGDJQ7CCP65KM3uANeZKn9lcPDW
0/I3jetl1pyWZ9hZUC0TVkb2g15/g2mkEBAoqB5YdREyj9ZXuwNL3f7Ks13LXnUS
jQxH3Jnzw8gINsmBWkWT1LmxFWqzACS05zrkNxbi0PvArHL1yS+hFLAlAj6lAbpz
etTAdiIbvGI9lwYYiaydgmGyMNFgXee508Ev8isCEGacpPSF2+0ccJ0To7yIdxzp
fSporwANhVCZ90Cujk1d3MpjFHy7fKkNKbaC6dPLh/aQl+o2e5u3zB/2z3zjBN4a
hx3gqomGw74fUEi9qUlxHmG4zICZYVmCBuLr479lZAS8TyQrK7Nr8MZZrxE1YPak
Rhyk3vkRWFewYOsbrw3WzhQZcS1yOgWKUK7PVC2sZHfgqXXu9e5hFBweGxt65vZr
M7LJpJ3mT6gHpd690oQ8WsaVYZLi90s/atXByWP6gACGHQrC+vGzjy1yKGU9QKTo
lhmNCYPLIY5kJnkyq8maF3kaA1Kus/dwOuBKAev3FC1YrwKa5/dNXPPOV+gYkIBW
66Q8AC7SPSjByPCxTCaKsYsWNAmQkfJjUGzqUakQjGgzoYG/I6PtF2oND29o8R+e
7yPShtOtmZDin2TC4acLE6P5cSZzd0p8B5o3Zu/pV5VeLYdRCDgGZUwXrJ8CQpOL
03MfXX2Ft7nVYIYmGG9V669CKCx24vCbgqKILXCUc684Yd1GRTq1K8bqOl2TyPP7
q+PHBYo+6NBOT+73j2LpDNifWFAs3v5OGlWn/PSSCHlQKtoqk/i9UiumnNJmxDjd
R8SbTGPWqxqgWjHs7/Ag7j6dZav5U1Apg93CezfcK0dZ4uNurGhhi1ciPvgY3rf8
udEfnvpzEHC/RmWHnJuOjF1rNwFcSSyIydoZXuIdsXfZ6qM/L3s0YjGQHeZfaP5I
tWI2TL2LAcv13f+JbUA7tNLnoqSaMmRiUTSJm/ezw2BspLiX7EnsGynP5XygoqoB
HCjO1A8wTuqlAmllsBUUhLV5t3/Vkt+/w38jOwRkibv4ZKt83JTVyL8/hvZfOArf
eCZ+q6ilVBiBmVgGAgOMbJ/++MQPYJlFu+RJnyTIqSMd0ydZLf8Ig7GiCJF6PsoO
6QTHsCWu8fMCmJoI38LD19CJaKqhLaFkqkZct9FGeyy5iMGFo7eMMUqPRVvBR6VQ
fWsv2aicf0imzuNYSEQ+GvmRvcqKkJLU35qrUiSUFlVzM6yPE8d90+0SGq+8xhgH
+qb0MX4r0dKR63MPq2w2LhFd3gZ+cPjDTZR4X3ZiIMgwrsintUvBPhWRPZZxcxjJ
aQ+0oO9EZ7v0nHJArcb+iNeEeWJgKZ7IhkUCdkH8p24rR7pbpeP3KNkNoigoLbob
sFQ/AKfHvPJAX9vAhoWVs/Iq2a9+dSWV6MJ3WBAHUej4bhWsvBGgHg7H47ti00zT
1sf4WnvCsl5XrJ4U4vdThNao8rw71ygW9/7fyLnfi8D5XdzRD+ZSrSUG7iFVCp0T
9yebjL6/QVCZMj+IYfoy0d+3JiQlfo3bFOZira4EuCyTL5rAQbY1s52y3yj05qKt
u1qrs8+lw6YMRM+AmF1oI1TlhDgU54cOCTjFguVyiH2isgYb7zTkJU4IZwX+Qo3o
EkYSlCF+TnQstoygvuW8ABYBXIo9JN/s6DFW66QHTNEpgYAKaSJfHohEdHddtVJR
OgF9REPLqi2zab3CrLABG1wLXdkMum74w9oILzmjBF3QL5WwgrQoFviPWqu5xJ3d
KpDgrVn3cCAgpAmVz3dKh0HnW/nPunKi0a3or5YcHSr7yw6gT6OZ2Shxk05lXL22
9mrO9whKrBg1WlJ2JxSkA58ltAkArkCXYtkzkDvEfS3VB4MydVdMM0V4x9SLbAlI
k/R49BPLoE/sO411dnwYMC4rKfBulnO0yUkNrJpgDF09ZgzbdqfxBS9Nj26cYj+C
vOf2+ljgfaQNFcaplbeVkaUEbb71DPn+4QXvOnt61YuNcHnpbGT8Br0Jmi07PaX8
0UQ5Cq2tnzTXvPhfKhf3R3XepYV1rEhFOXkKmuKr+s1ielSP4q5068FqLRyDAs8f
NfYNNh8TTOGYnB8QoJnVzyb/9/4kT6ep+Y6B49+n/CJgTXE6+k8ZoQmf4m5+0b8h
e4qejoxdhBQ2Hny+xyxYJMeGaXa+21ikKsElI5SP8Axys2ucUAJc2juZuDbNO5Iz
Os04ojAieKX1DtazI3B53yyC+rWyjavgVy7vH+arTY50cXVRx3Wx+LaC+Vx+MlwQ
pKuhKvFuIIlK+NdZEpDPd+3g6j4z6ZW2SmnR16MCFX4IiKTr90+kX8zaxgfe21qg
p80L9DXqIo0t37jcM2hKqLmhk9SJgAmcqFMR5XuZoaO2udioDZMwoWZJeSwSfgw+
DOO0GbGZm6hrZ9y0KSC/U9DuD4f6DWlRiskBqYex1yhPBpPiN6Yz2UOv2tpyVw65
zbE32Kz+i3jktimreC4MJZnIcKVlkimy4Omwk8vOpaUuRAx3GUlHLPyjQMABmgyu
JR46k++4u9eb8HX24re2Ly0Sp7lp6tQgsradT02CkAXeETx8/TDxkF1tmuMTv5ty
XXZvo1ZQReRI6si72meavJSP91Svb13H2fmsks3Uie2ADjSV1lYz4aLSdYAKhSvF
NaG6kUtrBAukwbhTn4uXt6JPJEIFyFX+YOJkMchrrmhuieAsiIU/uzsWOkpIN+hm
4pr5O9MN5OUyQyREgXeVmFsukiasUqep3u/IivK4IUyTcEpG8WWTns8aIps9wSGU
MlYevseNni5na4wJC5Lcfs35GYHdeNPvy4aj3aM572iwGrKNzKt0wW8gm7o7k3nx
AoePM0HITDpEhbU2zNQXjNpoXw/c6R/saDQcyBAZ6m/J+6pFblk6vPxPKkpt1Iy5
58egGp1VCLzazYKwZvAHwxm0icWWijE5uGtlQ/Y2MfUCrWJcXmYL57CpuN5NjGmn
zr6XyWDSmQUNfkwPFO7W4spaYVoN2eXbLrpqYBYHfOMCCIUcI71FvNEZKJL/Xf99
W/Yjpo6qN6GOeRmXMTP+Yh2qWVdr2beyztqprHSZkxN3hGDypK7kfzHGNyrpB0NF
UWHSGobIYPC0t0ByS1du2cM6ZCo1mJ932Zn9RJVJQGgGXDpM9SBwkydObe9r9PH6
UtSbMdVmm6+SyOnTcdGTeRgh7SAjeoROcHilbTbODbAJ6Krb+Z7VtdL3NFdGTdbb
6Vq/KuLWEiSWrvg+bBiHHtnPnbbPQ3KEGMumROfwlwqlSI6EkdrYkLy5/E1yjR4J
OjFVZF4wMWFEzGz35Yrjhgq/vQsXRLFK6u+YTdCGWRlwUv5+O6mLPo0QCJA9SWmu
avw6FJ+BvHZvTAKp8x+1Q8pr+fyV1gFNioaxrtgt/aIExnSe9ukwXpUq+mBiq2fj
48sEvLDOO/kDnlQ+Y5fjrrz0wU7iyRmU19j4kuo/zUQWrVKe2kPWkkvY+0D3H2m/
UjfU2Hq3vf836ly50XzGq75MHoFdN1ey/hYRkOGgMHlnTlBu5OTyKJPjt5dgQxJr
UmTRe3lFZgth3Mkj0rYowgTRcu+u1dmZqJV/dKH6Y9g6wJGSX8G1wrIiqSMEIcVO
NzBAyH4LzzCL03EKyx1DM5gtLI+uZQyafnNUfCAVXWeZJRrW43eIKF0CdxAuDOqC
rrQQXVuJgQCO/wZ1WJ7cPL8cpvdwYCmuuJ5OJKKcvbo4EzJ+ctegUqo4fqbCNi5/
IjLsEC+u5Eab+ihnWdCV3/1Q/F9ltR6oVoj9N85GGlkKNUVp+fXqOliLzwHHpVmv
ihYR+N+Ji9lDVjrqGdhxqLVxuYU5HO5oDojniFZwxN0aYACb1t0fbpp/MHa+Z8i+
Tn+IA1AbFdDo51mDOv4HF4m4h7/KWk/KHpRmXzP19oNh4k3d9xsfvxB773cQVCDf
iIMIWkR94BK8bJERafLCFyrIXRdJTSik+zf88YHEPdjPgEsnOpDk/Ff4NIJ0yU1M
Bk77lV72v6JfVrs42IdyPdGM+YV0h+BFS1tQ/1BEqMKqBTnJ3ffJo1epVRAz+KIj
plHumqbqIZR2ZnV5+SY0VzA4dJjyXYxG4H9giImAi2wxNlxlnf4G9r/Sr6OYNp4T
LG9g7M5teVfBCy5Mql+2WbHNFlDGQJThOCp/u0zw70ivEoVhWljsZ12Ru58Yb+a5
8QoY0ckYEOnMvXs2Gs0JubJMXD4kZc8LVv53NR2AFP3bCGVS0+NW2CdXVjEcCwrR
OceXd0ITcB+e+ZquxHyviGiB8TM7amFqqr0tk8dWruYMerSTV07N0t0iMwiAX34h
fDiVlUFAp6DUmAg23r/6b3sQ7sB+EFVDVd/SBcWwiosSrutBpNbrYS1+o+vWrN20
jUCPAdb1SlNvnp8son8jb3+e6tM1mNvWBA5oTWU3aMggQ2obL5jvv27zlw7iYLsG
APuCOPudvD1/J+6gvrr9bA5G+txIUDvUyVZ46nn4+J3djP7qoWHX8P/WvrHS3wRS
ZuI0N3SLI9O45lGQ4rmi3HHvQy5xw+KmksX0ak4TxpkdYvaZGW5OEItkay6ttwml
5tejPOe1W+N5FvoFJVuYdUJ5ZAL1JDSqLE9iCbsAm0K82WE3Shm1Ym4PLAAzaPfy
IR0hiaG6kD83KQ5b4IBMhujx+WNp92ttidS2a4ZBr4g3gy5fvo/3tE3fjd5j0oG4
FaxHAOxJtYN5nDMac6v7ZpiRGtnwrWWpNNa070cqIiWcgVSD3pTPPRQs/aMklYIE
j5RjhCjseOytxOHsxlJutDBXSA6jCVtRJfl8/b87lW4jTKIsChTwLJ6isesZNYQt
isSg7ySARq34rtm5AD1nGicj8rMxb//Fcy3UOVIEdaBIgIgo7IJVTLH6sEISsQEV
g7F/HCKhTr+sXR1V42XRBFww4PMS1VRuydN5lMizTUbvKirib7HTJYgFIAUUObTa
sz8QMZSdi68OcDmUtDnweqkrZfDX/5XEeT6IMLG1gvtrB3p2MX6BFb1DFoZ1RKJD
oZqZTbjzDyv8ZBVpSkXfdnrnm8CXKRQtPC3/gfX/lQX+NlpJcUGvuBBqYlFH4RSQ
gv+1aYpSQQDzZiQ9CiAvvNlxmksKA1QG2sk2eHFy7gmTo06EgygcizxMJma7Efpm
k+BfrtN+0XTtetvlTTOvVdPwQ0VRS0gWOm3RJavogkDTDvZ+Kb950MkGfOTbN9tk
FdzvUPvNfEtwplZMQupX8C72O+KDc4YCVMcS6JIGuaO5oKxjIT5J13TAEQIWR9H9
3X4q/nK/n64AG1KGaMb185Mvx6JIUNMuCtnPySz6sIabaP82IxUamcVVYRfFFUDq
XhDdWf8tGt6p7KPJ1bS0yb/Vfb9/243qLUSKAd7kVQ4N9/wi5PQDAH8796xhiZXA
RHRe0esu65QWArO6/wgiqvmQU7yk0FGKFRBwfVra2CEOliYWNHBejKTHRwbV6kEt
elreWXn0Qa3w2jF92SPhSjXs2T3TW8/PL3POidSbnpAuug41oicXpxGb+EEL382B
kOvGSoumU0mpd+C/rTOCdGercnJtb4mm5TydLR+Ey7CUswNd+5z2kmwfwC7s17aa
399MpJFiPg61mIEOsBFyXehzTO3cYZBE9nRU+HheHrFNqwexa5h/GDBFXva4clTV
hm3awdWMCgTEbDoNw5gdQdjJ6ADfSIYNldfKYIqBmluFmrKjcRx+LSCTX9m0vr36
UqWz9F4TnatTsnyBe+RrG/GyMilYwb0GWm8C98lePEPDCRGQI1wU5x129QqjklGs
dhGOHRB4lhNpjnhyb0sDqmg4bep03ePDCH1pfaTkS6gRH9PIUc8hU19yCc1dX8iq
WRNEKZ0ub3gxOrv+VsNx1vfzgI0+rqym0EvL8WoejJ9morlsfKVTvYmdI3nQpcip
RCfvujZNtCt0lZk8OS8CgHRSuTQcrCFNVvPD2LHDdF+e90C89GXzp9ZIWE+X84fH
YFQ1n8BqMu9uOlmVGvXdbWMA1Cn2wgv1OyKZ9UDmLSifEK8j4rkif6VfQht7vzIX
yUcr5r4Y3JBgh6DamgjwtEzE0U2QBxeBL4FEvUcEiH2fyzJJ69VofUmEEu1sI6+q
i3maPgUK4m00qubi/ztS7TR6a4g7PsEWr6nZF5ptRplUbE21NSHV9nBOdzdbaw0K
h72RReeRSx0sJEQhGVBYKl54f0SmahSf60x9/pUZjzqMT+BvSO//q9YP/vwQ5E2I
I8EfQLi0oL9jQt1mlRDNuUTOcsYV4dn/F1q/4tEcNRMgHnGj4XeaxohYE7u/yIHX
SLupFAhYgZN640vLdGh6YJCQ4HBnJnAPqOvF5XrUJv+wROcth7JsunU8PlicgGGq
ZDsVEnY03DXLAkRJXJIH/YXyxvyZcq0LG5jPI3B6v0OPeBfMk28kJNjne5cY6K5I
sDy+WklCtgtyj7uGu8jglTTMTT2/Khp6oq4YL0BXTbhOBfIpniFPmNbxsQszgMjU
XQS+stimiJOrtifytzntWAIfxI2OkdXfiKf8bQZ8J7XxsQwoJUXPdhJM4Ecqt5gI
JZtv14Ww8xls7iZKtB7mxBcfPQ8O0rRdAZ++riv2dAKbuKGJTIywaIe26SucG8OH
f5G+iI1JF2A8e6fzFy8p2j9PrRJIfNQ3vQaMmEPsDoDfrUX8wpY43ZlUHcEtFTP0
0GhOf9bo1E9wj1sVsQTaxSQi87sEnK5enWoDcS7wHgLa78M9ZairWwIsquP1Xr8G
50MdRNdlrfan7ww8cpuL0kba67GMYyyyEda4wiO9G0yGSnlrAlPitL6hq4RbQPAr
q1JByJ7Xam+dDGYG2FuUWi3xj69IigfiYLfOl8l1GsJYBAQTfKOWyMrGuJuj5xPP
W66xW/CL+V56xo/T/Z65emMMGxJOtUn6BF+tWCYDN1WSKCgiDiyO7l2BNwoeViMM
mYju19WZrCZxdNi5/+AqVXDSegnpLvGOewH3hFrjZRc6HbGNXmVAubyxo5Nzjhd+
171MHj7qx/B+nqaVU4lju+KnWSE586uzZiYxKEmJBBu8yiJ4tXDhMfYe02KOe5Tu
JlmFPl938f7Azx+tkFWqzqL4ZNvUu/hAkjoKN7jH+2FE6Qv00kEWuHVh92PJ9t7Z
1IW40YDbqqjgkJXoCtrWZ2VLoMue/tI+kByy/bs9stW83K0Plo5ijtYIgWJ/U898
QAM09Yw79rc8IWfneTGNclmMyuBWnJGrpuGelmiJMkW2oRLPiO34A78SpM/mQOfK
FWO/EZsOqRzduj6JlkGvRAr2c9D9qcnH7eF7fojOWRpuLGa/nOyJZDWc3Cpv5tC5
BVEH0mGeJZnj+X4afNywCB1t3G7lHv8+135dazeXM0uMoiCqwFvMdeVSbujdRX8s
I0RwEqZM6OvWOVzduUL3IhLp6Y+Pq4PpJyrctqCdRXr1BNx7SjaXFTFhRBOkK+A/
bpjBVGuRyewnMxd14rAo48y4LcMCOGS+eGejlV++A9Ysme4m7SZ/IrvawesVHe4K
fMfZuwhe9tSeZMLWXTbsloDXzgIRs/WxnWxVqaTVDbaXiJS8MzVpwjTtVXN8/+z4
ErlAcstOJosq3AU1C//z4TcqluwIz1n/ftiuGS5F5qDo196oGkRStUvnW+X5D2OK
dJdKd+gw1RmE5HyOO11RiDIvAzh2jgXrh/5/FvsXz4W57gTu72hSNCgZOB8oLTHN
fTUewAJ7mwP02YTNjzU87ULm6oJ/sT+A9GXG5u0Cc6Hu6DQn0YmVTZsEf9vk1Ty1
Upj4jLXmhVeQNTRShDhIVZksjoWYkbZKKXblpK27/6FiJfAMTVbTULllPA3/+Uqc
iihs04aQ9LT0yzaK0SDfFbTJZS8YAlvmD7njfnnroUgSxqKJOYGyhGS6DS8m9Oyl
4unm6eN2UBoj+X5dBQZAnQrPdqsa0PjXNRjbEYfjFwjx4My/y2LsaYrlwU7Q+Bok
gOVunNeR2YfZC8qiQQR+nR+jrqW/UnUWac6frUbRUazpkAwD/I5kDEaDWTn1TRzX
rAg3unakySm+Ip/AIAaM35cW9LFBCTCaUwpNQXeTd7bWna81YK0CQ5vrhaSUnmq5
KRCS8pzBT/YkV8rJCOXMFNrpdcsu70Jc/I9LAttqRfEDdZEAaX8kTPvXu3rbsUIl
dSxEmj7cblgoXSjJ8KpIepfeVARSJuY0ihR/VHvqFj3daUgNi4wTTjhc9q+OpU+i
sZqR3vcgYI3mpsr7UFqwWfMjvUkuSK4AArTgAS46BQ/QStwKzBCl2XeSb0itAWdp
aDDacHyC4vj3oqHpQD8pgWJxnxra4X4deRXwyeOexuqcWjQCpXQQlA40vpHfNZww
mqvWhzfGOcVy45rtpYBCYrkMiupD2fZfODeBRZ2ryspceYwgZPzmNbfA/u1hEJ89
40zxCAhCaKY2Nqvz//mTmOLUGiiEiff+4db0iNX70nASo3q2nxop+dBSgE9NO6zz
0K7tmA/XFRfYQosufwNo74uR5ha6aP6ie5OSdMt6YyDgncJ1eQZqMxVsR/ToMRNs
cpfsWWikUX+5bAphVmcB1QPtonpIMn9f6S1VxTNhVqq4r1i1f++tnP/ULi3/dOMC
xyKiVhnsEQ6Um0MllMh92SI3sni3cIea6+Or4eN8mhIdh9hGxsjr/mW2sJSQmA3P
JVFeNC3Vr3l+mJjUz0HJJxD/atXkI8ZUyTtEgIHxJLcN0tCa4EHy0ogDIGQpuW+B
kk2tCPvYyKqQHcfE8jeE61IBxhH0Ip/hr4QS6/aUOTSPFrgmWRK8lrXjsjusJPP6
3Aa305iDzacQwg0kApNovPIP0KfLoMu8raJDmVlaeComDtix8hcKM+JuywasOdhv
sxax4Vt65tHo5BE670vJqJlfpbnThIPWwxopdK4dj1RuARWy/bWPYMMO8IR0aXSj
EaD7GDxnPPCxJOdHQ3k4SxSxxl30HaG5bKU9oNk7nNaz+oaQ5uFdW+Np5Is3tDrK
sh38vn3WVF3teMrnqRmlzJ5/5wzunnbVBTRCyuPkoMWAg/Njg9U4M4bPB/UXXYwc
gUPIuxLI8RE4w7ljNQq6a5NA0td5fX7HyNkNNisFXwDuGldbMPvxUgBMCPK+niRq
1tZv31yEqcmliyjhh/KTvrYJmPNw1l9P1VWlNK8l8g/RCaSEr9gVvq8UfV4xoID/
X5jN/TSkvmOlmIrPW27xhUkUFED6Pgc7xS6pa5ys2MvXBhseIW8wgOghEaA6ZfJF
Rrt/gAgRF48TzRT0lQDYJRW1VsUqvfbWh04G0cz4C8olSk9Wx+ZtLsnSC8fk17X6
hgHK4DwLcKwKbAn1QMPyiAlv2T/GHkdVX0ntECrc6pdkFbmIB5jyCSpuC2U1HD03
vmHQ8ZF9f2FAlXM8DaP8VsSSMN3v7IpK+vMBFc0Nj0bTHRVjoAnqOgtTGQ7LFNMY
9owSAMVzMyu/RF8RuSOjA6gdXbO7yn1uemsUMqQdnBWTAZP6KuzinHHOQ8uwZ8cH
B1aXOncKQCdWPp7kvd1c7EzCLSt9G08fgVEeYIE7G+iXPMXEirUyKTU+zojP+s4V
PnqXiIjoEP3+8/V3iYgPDGKddyhMskZvZSRbcvKmVukF+d12O0QORAJGsXJVcV+l
+nkZIHwgw8Aj8y26cyiXGT5Jh1vyzV6SbwI9oUiUkK/JJS9ErIaTeSuQj5UiwYVC
8EZeINEhLIsWIhKDp0NPd6ohTwCwFo1/RnJiBZzQVA0Qwe+PGc0hyF5bGf+OPwG9
vJr9jPnnWdJNtVGCLbZrfwseQaBUnGN6lmuJdKFCAIpg0MgNbcYwvfyG4tRA/qN/
U99BpFbhgWAWS/iWwHy7eVXIud2zX1y9GY2AZO+OxfPCHyuj/x74uZbgF5GUHkrd
lsZUUrQzZOerQkJAZ6pxW4PyI89Auc2j7F0Z668a/YPfx+D2C1pjHF9tewy8sNS7
bp5uRUL+FbdIKBEqm0qz0AYStCz2uykjm7v5vHDnbWbfJCPv7CeDJtHD/qq0woYr
XFlJWy/R6al/8bCVF+/qi42xRuKEriMU+7B8qvtjMYuQmqarZMPJ8TozxMs4YecL
g7TQtyTx12QDVjH/kZsTOb673YDUX+v1LWHIKoHhnH38AZm3ZFY0wGt23ubbrkat
NWU2Ma8jzwxAsWQEYMf8gKWAFXYSfya0VCI2VNHeYA0xHxlsy4TmAbK4fXrdehpc
CyZ2r5B1P8CUOOhk3WpVc+p+ldmPqP4r3CD8SebLbVRawXO9p8ufhzShkz92cJco
cZeFJISdvxIXo/eb3SOpEUxkNEMo10kSR1rivb/kpdl9CrUlhePo9IxwdzEhVILZ
InowF06lKATngm5fgmInv4EfTJBrNy534DhUlFy1r023MTvBb4U0NBp7s/hS9fWm
e7uzJ9Wve3pWW+M7FBxQ1baYCAeQE4MgT0EHN5DenDB7JoLG2O13mTIZZR97opi2
baM2j3633raTPb14ZScrARlCgSsJLCGsHN4Ng2vccmAVQJq+IAEr1xEGDODcISae
cXhOFLNDJ3oAO4QcnkIZFPzmv1uCKOANFVeZ0qnCDxfyaafQSYHSRxu9aOX3pdCF
dOMkBKBQjmDdJ2wLQBN3uQJjwVHT2cJ61TxwLeHCAyfuKk4D6myml/mKieK8ZA5S
49V9cuP6XRj9QWgw4fDHBb3Yz/2rndwo0wWgDqI/dlJuLiRr8MZPOxfx1I9rrEsY
9Ftmt0E/30s+iuwzcfj5yb0KuMsXZbQrxI7hc09++xoSyizqFhNtNNdMZnBG2yc5
3E1jWorCzDTYO9EXsuLnlsce8goF9OuDoqmiRzGNy0Enm9PsurStuPnyRIfbDeBd
VJ361Wwjf/qxhbSieQ/z/JRJvJxR5C+Undhk571iw+s8tJSRnpeF6g/I5sF4ej6I
oIinQLorul9gbbg8J62EdgMZ6QTdZi/+BzmiquH/Cn6S6K9MfrFlMJWfgVnSRX4t
Cx5b4Z6pRYd6WlC7RqBc/7q3fPkxm1sSxDA5PzMxU2Trt2+LcDPvXp7ql9QNGgdM
BStHLbSRg5Tn5GVp9Z+x8JhWA59KM5vhlqGBZ/avQXTMMqBmxqgyjkspPGU9Tm/2
VADYGHzlPcqKdxKBrQc19Sd+AVpMJD/B1DhWQ8Z8Tbc9hHqk64Qroc0Ip6jwwkXi
opNBLrsbJf8oNioaGvEZ9jQNv6pY6uNqZatcvuskk/8EUqeE5uPrAhYkOS6iOCF6
/pExLZNIuS93vdYQOENYlltSweDfowoW/MLNwwdxhmllVAa7rvflNFzTc92fUUdK
ogu2XwTi5PvpkyAjMwNnLBKkfbZqVAsThXOhkRTEFW6mgyjqQQPkMtHQfamOUAaB
Fkz4EI7ciIynYXMCAD6a8CrY7/2vGdLX4uAI8kjNESF4QkmZWQZZWjqHs5NFU5o7
eRmkecB1SR/h/sDbQeqsA+3jyOkybh5VGX+d01KqCUpZCmiLU3ciELmHG4Qfceah
1t1SXzf6fVIhgyx1J5PKMUtwnwdkDfTMuHLIIRRpo40b4dQE2g7of4mg3ENf0jaB
VjLYIW38Hq75zGVQr5rZXtqa/Bx7+9vWmR4wyID+rxjrNuYLO/7tF/PC49mV3xld
D9zOK9k8FJ3IVZKO077r4dbPeI6sill2Up+oVeCYGHOUSludaAYuWieFkhNdMlgw
NOn9hDEgnUH8DPqq+9c2hgcffThBiE3PzLPBSrAcYreiEamL1ua7aJ8sklSEVql2
CNCyrCD1ycNQUaCc2TkqwGlBOII7m5bM+CjF7dJrospWPP1uwqFqIl8Fwpz8SgFi
VkyDxc9KuioVOxn6fefZ6qbNh0mYq9pVJpsmStH9kGEx1O0yOEwcnValBUC8xNyY
mos1Pfpe1X3XRnzwlEZlFqJWmC5AMe12QHI5ByLLi3EzgkYhdjYc2EyQUxn4re8A
70Ye87JZgUCjQzqSj157o/slp2L9kyYjl6lgq64s5F28Pad3jnKg2Ml1foRT+iJk
bVhbWeqflrg+qbel+e9tzK/kGLBa4p94C4cQCZAAh/Kd0bexYnNBXD/X4lB0mcAi
g9Oa20374hf18mpmbDY4TmsfwaejbD+16AHebYzmc3wT3hbZkMtf6RszEVj0lh3Q
UAwktxd/L32nrjiG+Gljzo2//UNaSfDWYDa3Q54G8VO80DgAe0T4kMf6E/fS/iiO
oAL0voortljJiEzwebjfzy/raReXIBxwKVdtevE3sb+jMCNZXKzFcSjkJZGVToOG
8+MS8OmCx4pRPrbfw9TfJGMdFB1th6b8/JVDky+oqjqOiDNH2/aREFPBSgmHdpbM
cwN6Pp+wmqmBOFiojwOeSZA9cXsvOvfrH5Y7OqaS4ihcXxkJbuA378RmOuik8OlP
AHKXPz1wSWRnH+MArMqOseb276xTISYk3fnYYgeEvWE6Dz8kgh1Oqc9aYE7W3Zb2
vngK8BZ8M8E7as21mFOYPgUaejEWCJ/WKQ1OXf3wiXSdok3MOvebYwytuoOI+/FQ
p7BqIgDIzxxYxabqtsR3KPQobMbMClCqbtjeiPhCdxPnls1izJW44EgRf4tyj26Q
IWjMPyRV3yX+YrJ/yvkbb7fSEvT+VjF7/oXNwlTAx7y+BmjYd/l0ISRzIDxPFxlm
u93M/oNkuA0ENzzCWjeVR/Bgosgoji/EkgiQZHctt76hOBqAd8LpsY3hvjSjrCAa
sRlJwODaMP6z15cBtlGShRmfC3c6c8WNKg3PEHqYH8Um0zugX7aW9SB3bVasCAm3
tgmyTx5SkBpwUULZ8sX/X7LLnn5KPRUmcoHBPFPmcnL1jOJ4y4TsWqC42qdVQl+L
HfO484rxk4DSUiLtC2j2sDCOhks52VoPFEicIUOw0cfxGNJuYDmcEsJoR6hpSVIV
EHlArfJPEahYakB6hWWOcc/EysXjyOvmmZsW5I1SPLNldhfvSDYcuHoCEn7WDGlo
hGwxptE4yNtBozQ+DH7VLnBz6lvEuwrDLRCJw3npZNpxzz3w8+obcsAcy+aEvoLI
MkX3TWnjnNN7n40FbvcAmfAV9iCH3BIovWWJgU9j1kOhXflzlY0dW3Mw31ogsQpY
rcRWr1PDJBl4p0k3UmIm67p0KquYWBCHn57wyPbfIUxcWco0OSb3TNHWmZq8jb9/
xNdCCZ/cHKJc7YQnbkjMZTG0PV1R0WkaM056GjvJzsC3gn3SPLCB+7TOKB5pLA8E
6dE53Z15Ul8+K3dAXlB9B1wqF5oolTwrkipnCAayv4huoWdt5g8lHyeiOCjir6WB
o11DjbqJvUrZvzjkzRGf0hmsaWP8wDRm000coLLSBjtoRPMjp/CR3vwg9aP/xoht
cB7QlMkz+ZzjE8FFYvR5uKOzHFcTpudM4I+Kagdq0EX91GLp5CMNxkdLyun1MJ3k
zdI0RMrVsKcvaVUpl9pw5Z9sxhVMdgF1fJovSzDOimBlY6LXZu7Ad0mTtLpG+l8J
qbHFROJzaT/GcdZq4OPpiueaDru5fdHVRYJtEhj4k+FAM0YSbJTVcU2f/ZZnFzdv
6YQMzoL+0SUnV8Cr0QneXWtnRrsss12iQ2adZtIW7plAWeHxn70vZR/AVlijzEoM
wAjxdLAgt5+jbEnBjEuhrmTUqv3x1Qoscs0OV9xZsqsAlfffZwUEXqBeVbcksUlb
pz2wpL+6n7uhK1oxBtpw4yjSVd33AxJonSBAjMzxGcc2LElBmMlWHHx+fRDPWBcv
ApIaVGW5ZR0KITpoEbrRcVJAdXkwNnrGMGWCzMorEy2nMjExRxnIPNODp+QDcA0G
wLBD/fXjCNkU4MExSQT1TTIfRZV3RlTap0bHjSTY2HybqDbv9HyntIfSlkneaOHl
cdF2z2+P5I6dSDtIIVf4Ztf/FG2ugzzHVVZIqYj6x3ii/IBQRnHRPhFkgtSQIDMN
rKnOaAd9W2xO7CRhryw8GXThfmWNNHCPIIoGZQvt81JwUS0zI/C/S5vx0LPJxhiV
wxFv25gPPpbMpp+BFgOy2yGzhTszWwcwcWUWOBNl1oWTUKenlcSYz41Lty2b9YDh
rIjuoBPb4D2iZAHqqBcgZy6wodKuNKGF7H+muSMPxNZNxuLBiCMqw3mmMbMnAhSR
KfbPsM/UyleXsvyhpcvcNRvVJoq40JVmgNViwoMeN8PwRYLf8XTr1MpPlKoZ3tcA
iO4pdc49ybHBZUzCDrxZazfIk/fsHGymsU0nhGaa8UPzyDXYDnUcg8cIllnGbRd9
275l4JZgfLpNNFZZ2bT76rxbpCt/EJnEVSHgyd2v6mPzZ1y7hInvv7tMB7oQZFkn
F1hsXGrfPOggiqi/e7iQ+XUlwGmpRGD9Hg/krXvaKmUuhChqqA8DNr5pzolh5a5K
RUpeL9TQmbUucJYS6dYBKZJLnXj3dKUcydzosoJhzKzd+tlJaIOfotf14QuK1ZaW
TksRGhVM56u1BLuclkT48dix0IK7zjA4osVrP863zoO9V7fyt7ZHBn4cZdFteHhE
7k04jMl2boLw3p5pXcucj21kHcG0FBzOEFTrenc7XpUauSJ64vTrrEFbBCC/TWf6
xlgx2ong6gyg+hUJzNiQbk5/61vgJdIApVE5r+ZaFSq6uAnfAgc/DUdJYGw8bSL2
Pev1nlEadENmWHghOIDOGfBSucdSzveRG1u8AdbA6w+j6+W/lMR4nZJG/57jC5Wj
yhU+pPTK+ehGU8/IWejU3pBLZeaLrVK3W/AsjgxhJ92wUWKSkPl+sWkr8ss1lZmy
qhmmZMX7iLLkG3Utbi7pYz5LOXgOb4oOKZtqh1M9ptb0IqxVA07+IselrCA56cKs
YzdbmodiSpsxs1euBqTpsZX0XH4/7BKflonasM1NTwnpHupw0dSt3IEuQd7Vac9d
mItwPBSBL7XOjlSnGZsQZXe4GBQshCQEK723Ke09oVb2VwluHut2rGcEEskpPlFJ
ACcgiMUy+3HsYmimWicz72VoPmRSQjMs8qTn//Glhc6bviT/CmrscVEIbDyvEDbk
w8TK0pSiPSrZki+JMwYX8n28pY4i7zBpPP6Gna8jBncWHlNR4OipWgyD5LVQRV4G
VK3xy4+F7mwYW+g1ZVSJBsllm+jj/qTb9jyj0Xw8pWUsj2fbkNmXjJBtJDbNncVR
46+gKHA9Akom0bzGro0vIdMaEUJDuo2FvowNeohEJgPc6S1/a8GWX4u6JBmWqa7I
RX0YkAkp5kpLmnF/8p6KHKsdU5nOU8xLBQf0T0ImIoDv1r/GWJJPqv8blJG+rf+g
9P3PlfmuwPt/ioCnyCI1iXcrjTeiM07QSG/rVbD7TynVVNARW6PO9ddZweJqKr/z
6JekqnvUSEMfrcHxU/l/fOCVn7V0NKb2YqqWcUyQZVt5f5/qSMzbif9J5stTnpLG
d8dWygZx6ghyUTEofb+amPVUgtEpIrcuzEnmWwQukE+2dH5L+EzSf9vXKxrKMUee
24EzJ/e/N0IUhC3Z/UqzdhS5UdKo5xhCZpKQvBNl1MPCKvujzfQTab/LENwjXDIg
3A9TRqSUjKiig0XrEwsb2jfQQCdOi2rdKqKutZkqVFGxokAK46m85qUBayfxLAvg
yO6/qqxbIl64N+Qofc8/KNSqYfyxYoLMhEolZMwRxN3iiZzpmgm1Bfh0INANATqg
jAYZZ3GSp9kkQwcVPrZQjZfz0FaDjMa/AsXFo6PYBs/w7g/UxnW8ZOZ6tzIl7xt1
9XBMkKCHWjUtb8VfzzZ+xNpnYfi2zzG7CJJPdsaKiXvOdiqOutV8L0Sfgaaz7qWn
N+JnbLhN3iA8xec/tgbfuyfRLKUbMQ1pw42kjv0Dm8l6r6VNhAT4UzsYLEMJ7x/K
LvEJWDgAKCC3Aa0zlIzi0uAjE8Am2A96Cpp/VHBEheQaTtV1pqbEJt3p7u0tKt3M
vRryA04wg3pG01PSMQFrF34QFrLDForVpzkpVsAThnrGqAkEFivVAAxugVf3c2T1
tPHCzICtDaboUX69T/sfUvaSEErsmWunab6ZTBudLHliqs5GP2W8mFgJuVf88zoT
/Rk6gWeal29I4ne3mGGcktkbr9YFx01HFrVGJ+/ghutwA+P0q2goziw6e4WE/70e
uSBFjwx7ggdKt+jTqUD4Bpgbyuhyw5Lw51Ty9qvE9rSz1pYa1HbSd6d/RQeX8/yQ
1bLQl9bsBYen9dVdS0LbZI29bZx7IdlA1P9QJqLEwhVMzPlxgdqoF9n6IbeAEP01
7Q797BQjiGQQvRgp6u+qj3mQDYh2Rzr2bZEHyRhnSD6jizpXTDdyqD1DDj94+S/T
WmEgO5SlXqceIMTYjx39H98OsF2hlqUmlJo5fqwZcWvv1vtFC3/oM1lj6DE6o2Hq
c11OizWPj7qqlmBPKli4kzhJasyam4aJYv1MAraHSnPEo6jHRi9ZZmYW70MNb8K1
r2zl2WpyeqEzXt/VVgUvTuZcTHSa4hDuUsa3ie9EBX/cR48thxuazb0sssWed1+M
/g74agSSIrA7hs8P5CjRtfPUQEwhrrWRHBj6HELE/rVoXs54dD2Z9BMNZZlbRTst
BGWdYXGSiicJrcH+2b76I5Jke29obn4EAlv1Sdk87UX98Rr6wSgkqfp5s7Bcg07k
fGTjKMoQDnhAPNyNI4QCERVGKz62BKnadjUXd3lC2jEgcWm5hy9p5K7FKCrISfCa
DpFZV2MUjwzR/S+LdAbNpb6Gj5bLhW4X7mZKdSLLkhU7Oecc7WpeqBf79wMPu6q6
Y8yppL2DT1DfdYtyF5abdlnTQ8Czz/XpRp3TYL3EQ/ENOGu6thBT/ELTtbzQBhBC
Hljr4kFlVML+Dg2+uBWvAtdT8P+bJWQr73Oc24YnJKaKQbp2Zrx9d7F+kFEWewzU
d0QK9m6Gzfw7c8mUED3D1tLtBYZb02vAE0G1BdR/HgBeATfnYnG2uc/Mf5IDiSud
IuH8pwVR1KfTcgjFzds5fmy63pFsipoXrAzq4lrtD/U8bTA/BolohKxfekH62NtP
XrFAOTlM8r6tS6u/0cj2/qcj/9U+f+ug3v0LrglFZw+DLm6hJWaNLStA0C6yHAds
5Me4uAYZVtarCZhVTroUt/t5EBxTBk8iJBblE+EzPEELBFZ2/wbB80fF+HxOjit3
WyqmO4rzjTCVHCxKJ0HbQnA7muAsa2LF6DiVtKc3yg7m/F9pbkY8tFfKHk7FpvRP
/jWyw+gO3kZCeU++iwid0Cz1UhJQevyuGTPDH0BqxwHAojSQeYj8R6DvgeyqvMzp
Rpm3fSlRp68iTGn58mOtd4Zb3gjUeYjRVSYY0+OFoWjXL/+Lk09R7SyPc9xpE5GP
Bffv30qzAC9GdwkQVbr+kZ2o9fSbWQwj/ngR6WSKOrGxUlIUTHafFUcVEFtRsFdi
j96NIbdOTDUc+UEEEw8ymejmU0c0ws+s10okTQOOlPvEzuKvutp5oa+BjLL27Gu7
+lto1/YEI/HFcE1aP0jKyZv+iZWRSDrsQdqNp+s78/TPrYSw/uFSK/1DRl3K27/D
tdv118CtvbgvhKkdrT4NWWadW+4ROVckKhTsnwY+b+PfmrhYJQPigKUiHCUf+nzs
EXff0JVnzEn6Knr8qRHjUEskvZHYzhiuXeOag1TftLk60ktmOWkYAGXc274bwQad
z5noBNLpbz7n9L1DoTU0rl4jrnaaUYD6eXVQuE3Sm9xBsfX3qb2FHP3/f6AKdrYF
BrfldIXn6BmlSPHvn20LOhDQRvbtmzYO/mc6j8ZUifK2xrriec/REq7ocrO9ppD0
AlKlZH89Y5lrAscGs7Z45U0UUyusKRNghhpNf6ECNuMC42rAdLmb7LZEa8MXZMaF
06FXpIxvIwZZQ7tHpuy3pUQk07KJkFJ1G6P6GuOeFqTBWKdqQp3OLA8Fly5eGQ5H
FbEuFgKfXhjgkHYixofBsmc7z0CuZg72Vw+KolUk786nt+442HhQpEwLre9OuKcF
xzfBKZJMNyvXAAoFtOaNwntoTj39WgLrU7Gcz6SgGWfNLTpW+gwBGO4IcXXGF38Z
PGKg9oumdD4RjHijDjeiFQXjb4jNM7I9SsoMmSK/g4wH5Ii+c4qmXPpNJYsHxXvB
xDkxnilGBVEe2sRyFgYvO3+uI3lN8eIU6zLsR0KBTGVeZvaWGPN6M3+mK/VS2LS9
m42AM9cm3HbMAcAJ4xhjQ+DjLzRDGopTLXSGS+3/zHNx45jBDMxkmoBS7AzUSzN+
ReltPv4tzkg24ZVq2ilJiqKNib3NSZlPQd1ZX9OXzdp++p+hiakmQe3Q70OV3Dzb
nldDNe6Hd6h+GQiGwfAevzywkBZOv5oklVDE3IX+ho6u9D6mqx2R8+zWhKlSWSED
LWOSRy7378wkCZ5+zvXfhHqw1hIz9NEhJ+PsTfJ9oPvJZ3XMserwvJaQ90cSYpTQ
BfiSa08DPAPRDAvU7PGeBJ2SSKO8HvcNIa5kXkx2FtydJHNc+ZB8xjRnWjP2ju6y
0PnUqcTfmqF0Ad4tQ7q3LfXy0YLEezwdwFaSYeHT6gHC4TF1IPKzwNhgrK8GnnqC
FAuaAvETqhMe6hv7p3rwd8WyizeIusQe77euqUeVBP9r3u83yS1yr7IiiUmMvzL2
ho0VMOxvwY4Vpb8pGgS64uq30hE1fjfJHl0AwTRJQ73UclyD2rk6+jjjKpEElZBS
43JHAPs91hr3bvsJpU9kp3LJeP9rqAOGRX4RM5koXpaLWA27VGt8eKRxjxOZxKyJ
lunrzsu0Xmber6iJZd+TfCq7NIru0sZqBmdp5Wj39igkF299cE1Vn3KK0QloRTKk
RCdFEE30wwNt/zHPgEeZ3S+fhrEXF3+eL+TIbE47o3NmZ016S+wOy9GXIfwUmFYe
9avTkl1KXAUAFId34nT56t7L6rPAoXD383gMciy5Yx36hzgGDMHyjzWEDSwqaQNj
QdR86dBxL46Uby5dQ2s2P9co19mI3yekvRb+EAIVBr7B7Fqk7tIAyIq6dwoETiSZ
nbiMwObcc3Tz1rokdJ1fSRkD6xlThguQP/GPnUkiJz7DhSUsWHM8+DT1DGR5rbab
NyMrESIYCkTLgyg4wd/y3zF1qb6f5CPheN3Em1s/BCY0X0iBvD09m6Ul5DvT8s6N
4lB8MLEh4tzdDxZxHyoFN84zREcao8C0TPXSI1jEg1a2NLRe6PwQgBQOzy1ITpn0
dIrO+qg/tBBrx/kJ571ooZ8ofpk/YeYrLrMvDLTg2o3XqUZXBH3ze+Sog3pyfmV4
tXR4aalfWxsdsxK1J/BbZFvCR+r9F2W/P815Deas7/ApxPrAC8Gg6baK3EpBdeqo
tZ+cf+IS0P7MVoNL5PQJs5lrRhUhL8FC7JE60XJh8emimh0OG/XMK0pg6chaW9kv
xToMcsCzHCslqcbCy0ceGriyU1FuCLzGlM5YwiO2BOW7usOzdHzyCi42m0ov1c6g
bW5j1SxDOeTC72NoUY9rE6cSlHUgdfKtxhzDiVP4Z9k/uRPoBi7T1RsWBIIkM401
kT4i3BXLWB+7N7BUirRqr1nXQW8Fr1ccar46XdhAFxQ4q6lyJZQDxx9bQu0/yExb
pMKMIO2S9SvkjZLT93lVhpmUol6231OgGaB5Y1oXKAQSV42XLR8cpTGSDRiHKA/E
z7iTTMtOvkFWfvac4IxWxm/Fvm9GWuVEKz24+5G2OdvAiAcCcORJ1ejlPkHxmXG1
HUf8+R9sz2Z45B8H7F/VXjsztqYlcqbq4hSMsgSbjgeT55tOjSTq37KZM/2X1HvU
pKuH6ySiOgxWhkDwJ49I3+UpxP9j7PaXfwPA06V+iM9l5Rka3NUSWQe9xqz/G6hy
6ES7tSx03UiGCaFYu4kwiyZBscEe55hLmNkL/SwKUOVN1bNCeXBMj2Ex6DB/oZe0
sC6CODJF63J0tRcZHFejBoR7F8vl9qRSJZXCU+E1JX+vMaVYbi88WC3WN+IHEFWy
OwQ9Z9bJk+abzMYGjnkMplHEXnRDuogNd37Cuc4JH6GtX4UrXZ9DX4y4bqX2vf1l
44U4qUML3VH7OznmTxDbjOT6SEaHp8OvIJ9HEYqZqoQ6thpphQBpCYAuLuOjXTjA
wbxUihpNyYw18W+szC3hETqccvB6Qe0VZ0ED8r0kVpWGUkgV3ITTh/Phb5gZOWj6
ojCL79LOzwtzjYqVEDyMtuRTtaz63y1FQcNW2ivONztAfln0chedu9UG0KmJD7S2
EGkSJTYHQby/s/fHVvD5kEUlQjfp7l+w+/IIN1o1JMXT/uPav1txG0flIhp00S3r
8cvRk8TZtOw7qGff57EhQziuFS8SRqpWRm9QNh1phLRexpz9JjpHAjzL+uMPOhlw
1H9eiyqZa8tOYAI9jY1zUhXIQpb6j454uTEJ+seOg2HPBDh1iO26yuW4r1JVxnJZ
mmElj5R0xMeNbh7uV9eoGkSUgBL42GzRD2QNEjd2a0lZIiT6Ze8zg0DP7Hy88oNJ
0PSIfs4mxeTzriKk0syNzkS9eBlEsi1XtU5NAjI6T6IX0mpVOfWa0iiLzpxokaz1
8msi6UJzm8fYbSD9g6K+UesgWKEvGn64ADEoO6/eCrQjDslhqbCAxvzs5cmMFRTo
82OgC1C6kQo0jzCSe4j+tr1No5yk4QtMHDda7rsqRfaEqOIfxYeHSb70cy4s+HSt
hoj4XsM/hn3B+cwrkWeUwQZd2SulKdQHkGTMCcnZpJf9cbNFV0pgyI5spHwRKqD1
dB2o4Jux4K59w6zXvlnKfRdeMpi52gXZC/JbMlF7BB22c3nPLnGiBlw1Y+cqkore
9t1xTo5LCVR5BoqAKYZyePF/XqXZp7iXdIRSTSzAo4r6HYMZqCN4WdhNQJ/X7xdD
k9qvxO0sOwf5qPrzbUBt8L+ugKPzGSliDxN57mH48WsBvbKiGAVeIVu8HgSdu3jO
trHRIMaaTt6FSc0artqp0HVPc4eK+FIlSsIdUvuUr2d8WDxzo+WFxaqEIeAoAnNF
CAgevzZDM3MvUP/45kc9SvnUEuSKMIOxl0wn+myzJb9lJRPfjcn3Y9wn4YNdgXNo
Lhdd1tUcijecHiTLWCrrMHM2qgBsi8oooDzsfmqD5BTi/f2tauYXK6sWdoq1fCot
QXV1ufxedTqAeDvbaHnvLFofH0ZKHOgqkOUOXSWVhP16Nhz3VfORrPRXbtxdXvOW
nbyaYxr+L1YpjuBz8ax1Viid/4ptNlIInU//8nbuEd24cUmbdvvQYFmLSaRUuMKa
yRAS0eO5r3H7C018CVUvLeAQXB4n0tXjZnpTDdRAM0qBtL4Pu3vG4E9B8pfomFjt
/2micbqtPmQ1QQcFzs8z1PeepAFrR88DNMmf2T+5PxwBVB+yRZIUAiKUOEm19qfa
4UpjTHXI7u6lBsPepkW2SWzYUX+ZYDey/1w39VTYbtxlme8YrskTfJMPSfF5uJZH
bPrJeqEJeDGs2wmf2U4l+ARNGKUnIpk8I2g5FI8hQ3ZePWMGkrW0HVaDO7AxHcAN
XzMcJZbpnNYqmzFikseHuLz2NIeXNXHdHbzWnJaP4msFngC0sRp231ulhOd+0RgP
nG5hD1Di2ovyIsMbwJkcwrxaDICk0e9+kFUG4r8ws0I50e4ZF3SFbXC1I7TgXr7P
jP0m0+vf0RXOIIpTOVm8zs70nmwHBbpxeggwK2EqvlJVi/gUXD2KCkwTVyOkrpeZ
QgpkVNm9m4SIMCp/bs5bTobl1AlnAVIHobmum3+6eDEWnmOWaXMrXIf+tVRyLIEl
ezrjS1NhzEsKHIWcQmuG4+/erSN24wSm/qatEh1AaAK1zfMem81e0j/dsS5Hlq9c
RiSHkSqMwocZc6PTGS+C8bWdqkp+jMlQVdOksfQ8WUT2zqh8iSRFt6vIYFeX3y0t
3FIFO1kI9JzDbPkOKX1VuqBxSa5Fowv9bYVUuVUAlo/TtAKHwVwXIDagwkAzJgB+
qnbNUoKpO8BxZl2fsyv+ykyfSV7EHoRtS5ZfhktnAp9sbdgkrd/foRGuTfjhU/Jv
cZmw1zjfPK+KXbN7urc2VoVKCqqbEenNPX/a8B9JqAS8igB9rw9Xdk8rD+7/+kMu
AElubmdAR8ULnX8P/eVssuiw5SEjO/RzU8HkNXKeO7LUjFUkYCzHvqJ4rtzMfF/g
2GsyKvWP5jTRVCRZEzWedI6g1L+FweJY8iap9idjmWynpqOOW1caUdC/vEifD3fN
6WnhTcaCXaVxL2wWXWR7M/m2YSVjz6SE0VSQFzVO0dA0Zo0S4NfkRuWrBX8JYq07
24hUwHXwVmUoGxjFoiS/pDQv4y/H8ryAXv7sGntkzHiD1eVXLz1L0phTHWCYPL+X
zimXi/pLQyhAtZ9CFPC6pKoEID21xkSghrHYxGQy+5sdp8RAGLg9qjFO0dD872+S
a8AilopAGHQVHMccu7ckg9Aa+FdtRDanbJltlglmvB4LtFESythGRJI53RlvQvs3
dEgUwbAoBIh5f6QvFTL8M9GEU6uGeekJYIT1qQ0cHVkWd6GniGUApSqX/xl9Mdt9
PWHcMhSLNtKcY7Ppn9BbW6T3w5r6qDsis/tQX1P31ojOq+vxUkf7NkR9xM7xlrAS
Bj34H2JZQ0aA/3qZWnRZBrV3YMqC5p6z/bI7PqWl3R45nmgGb8GQw60Bw0+TlGrC
UqP72zojVoIkfvcR/rOIn2GNjW9nXA8ZqjIgLwh/gi/MFYSYy0jNkoNY1q4ldq17
JPyZ19/1wDr93rbgav3xVkKtyBp1Ghqf+W2q1GDJ6tuoozMzEMc8wqg8JPDMP5Wb
1Ne1kSQseFnZSlLfoMU6r6ijfL+HZn9Z8sH4iW7K3eRJJMxFTIg/650LyYPEChFV
udwkKaRet2ql6s0voScHPXjVhUaPSoJmXGQT5m5wpLMI1vTgmv1v+Fmc66TmNU7A
rJlZpBmkWJGLpbzN0+eEfwSzP5YW7Wkz5pIIepb/jJqgUGZpMMMBiu1RmDwbL9Sd
QV6lNvl72+DIIfoUEoFQ2rP96I4JlXf2MlOOX8rXt/zuIFnm7WKDQiCTrOxrKl9F
p7NJpayIzCXbRu+d6/WsioyotTpGsOCQszWFC8Tn7hXpjaWsCqePlWMH+pWSNp+F
rfs4KrWgv27EzyGMY/LI+KKwmlH2gSKR5DV487wEb3weKSLrgIe9g/3K4ATvKCkY
iRa8M0MPGPXZHYJFMWjAfK5g4ydOprcDsTnVqudwj+2SesoIQ1b3i6uClh4IZ2ki
XKutF8gT/EAGT/f0b4pC4XcfXU0C4DOZ6hZ3D5ssgO9J+aPZMoZBQZQyTInfkDuw
AAFfRFmUuiHuPGzRigUq6de1SIMkYKs4r+lgtNHzwuKx8aYgDoLdATg0HHsd+7v0
AkGw/irNbS/HGLlsHaFHhctGqCUDZ29cRji1915IhZyEBu6qoWI/HZ7imXccmSvP
r9+vB8SIQ+3avHLHWw8+7+9XVkIQobLuPIgMRDfz5te+8tFRWCg+Bam1LZaMVzN6
GfjzHe0aI52dPic9vC/Cy6ZkFh0OYEr1qgBGkiw2WaD1qJgi2JLnmW87W+CrC/vg
r4L7SjcLikb2zNEDrtP39L6yFI0PtA3WUEcXwcaIg1vE6bofTGXwinn8VxKB+ggm
VvDWK/+AAoQMGGki72jlV0DtOnawkjJPMRuf20h90Jqw7QMnr2METjjUnUmh6HJt
R+oAe44+VsgHo4iTCBPTWUdyOH3vUBSM7BwCPvn2THvdi2URGTo3fqKcp48LbtyY
Ug9W6Oj4O5onac3ySnMtsDcsm4YUQtmvqNsjmkKMaFmK0sJHdYDqvs4FXJOV2j0v
6519j5m/CUyY4vW3iEnlzQvWnmLjt5JFBjS4DkVtHowv9GlzYS75hfEiMHyxeusj
n31cIjreRNAZZ+Z+9/KgNKtjP69znpsDsvkjkogGj3P/Xe3XdVZsYgAHcUMOOMQ4
yr7vrnOGKYjwJTaShWltZHr712LiU5vDm6sr0Ono68hKJJUzbR0MQvsEYiLnhQrE
MN7sXtBm4nWDJn8XsMK93aV/QwjbJf51KyEPXjMQSrd1eGiv5JR4Rd7Nxy7MDbxX
9ZFM+FheUvl7veA//C2e0wOX2rzcfwiGwKF0SX243gaQ025T4j49B+M4lKVQ57O2
0PMc+xVCHcXo+Y5xu0amBUplGz/yeZB4W5DiGm3T2BbvqA4qPP1qvN0qvzMyUkfJ
f+upqE15CMqx23mul4mvd4F3grxW0QB8vFnTP/2Cas0GmOrDr0dmTbc1/Ovv4WzB
u4uBX8NjJ//XgqLigVHq0LE0/G3DgLBEIIdf5e08z2ym4PHh/mIrWghflrI4Wezz
osLiP+rJ7opWpbevUNxXgkAuS58rYIAiGWt923IZcfM4rafoM3ZGrWAMqEWnLX8R
goi/0Pec7Ahzmw0WzCoFS6uSp0FLZ7hS+5Zle/p7QyUaOVekJ7fhR9z+kpfdZnQR
rCBSXkF0WdE5q35ZnCGQSxueCns7prny8i/bPoUU3Yeoj92ETuIpadG2aw5tj6Qq
ZViv/QWvftDrk1PIvEwq6qM9tZh1pTXzdFGEXYfn3IHChR/CFyp864YcvV8hNlKp
vseyGT29qFcM6a8muFWgLQjL0w3KDWaE5lWFd4q9ee/pcpXhQz+Tdjkk3oY+RCcz
G0Lx8yqkuTgIgWEFOJiMkDkXi0LbFh6sXHegCmydVikoI252LIksMskd50+XSzEN
jnxRUNuqPEYSjEeZwFPRQmtyg3vxL2yX9F2wvLtgH6of9hWTGEvufHrpWfhYM7yH
9Satvr4o2UGV9wgGRzV5E3n2nlv9PLEKVxA+U9lPfCIUCs4+ryvq4lx9Ihm20qJC
wx1G4COtkCC5qDh3rcV+Ezl/E6AkjZ3peXUoAT2PEYXeTz3VDFLF8bLJZNHcOZ25
6Cc7g8bvXfXIcVEYR6LC6t1zRfdDocqujpb+QvuwaVjIKd+1/WvkETF37XaT1hVd
CWpkAsL/aE925U81mjrxJpa5mjPlVFHvEcZHslSemDK6Lwbdce6S/wAsAOcMaVQn
3CGjlds8EoddCiKrJ4oxQYLnmLd3ZxJE+7Hrh1kSQkKVoeLaYh9nwmzrdFrTapnc
+++niwEciujEzTq/O3YrF7C+v+2mLia/h7ci6K3MMYEYAuDrPPkup9wcUAxGqjfD
UG7njbNoNb6CQfY42evcXlYooApHj+0biADgjPtgLLomkhoJaQuUAUqobyWzzHm2
XA6MNcjaY9ScHsvfeSadsU1AWFtEbCXNfoHlHe7lGmBuxF54oK1nMHZILAClwbNa
FYu+ek9YAjXB/yM2hD6hkltK1kmKT4ENxgAms5G0QpVSozkI0PtOp/3tqt6LdpTO
SG6BDxHFOTTv37IHrnMLSRgqC9zPsfAHYTDAtA361FOvwsdbxYfcukhlawe/PQWN
Dm07r44TdQWMkD4BkX1NOYwMgNjj2n59rCmplV1IJQbgvHotAGFkKSD3hzmCyLRP
Fjb9FEirIb9Je1lwBUvDoh0tsKZ7z3FAMvkTREWYiChgQJiDLYpWWIQLcst1Ho9C
c41S30wzXr49tx1N/eKpGHhqQ+yuDcuMGd2QMSm8tL67HESwRJafYJPqIHbRsYcV
wRkHYui4brVllbbxoZ0RlRM1YKhB6AoFVcBE+DWzsvEjm1Q8SvbIi2NGiBULjqXP
382SneQNT39QLgsQ68Kj/mOv68D+Ce2ONf/2wNukC207veSgX3FjjKX0bjEvyQFd
ZTv/r6a/GE7LrVdMVlCzDj5yWxqrqBVhsZECILU2boNo2su3mT+SSuBIugg3EEPJ
N0piGdTV1T5ofTiou2xkBDY1qyn43WVuSczp4SIvxmOAEl9G73WpqtLaq41wE1If
u9N5c5Lhk77mGb0psBmE2k+3CmH2hA5XmUHG/DcaUN9eCtxsRoWBiHWyCsmITxiJ
uUDY9g0Yl4mGOsfwP86+Q5rg/4dul8e3E8ZlG03RTpbxOwmFVdRjihBgijSRvWXM
cJwJSEzGA3njmRjrVQzg4oEBvuDnl3GBO6Jqs1bULh/lsqEq9IXL6VtHs2ytWHZt
lzzdTjSFXE2mMs9zmNy5AmJd+/CmxcOb0XCE9fFg59mLS6Zwr0KOZ+m+pECINPVB
mFLJ0FaBfa3icmqXvcyvNkLpO+ooCGHZ/zDr+dZ9+HeHIEtOT3gW2g8/8KJV4pyu
tFLGdHfL63BmlUkS/hZq802gf/8uja/iFqHDCkIsQvrU1lot2VZJbZFK5y0xf0rZ
xmM+ej9VHjTJXgEDOa1yMsYKMDDhPZSXEmUcuXNajE69qn9lZaq9ioPJrb2nrtuK
IoGbLAuX4XT+cG3eGVo4ZYVzQVSJIthHcoCJrFE0+nLSmHANXfPiTb5T6NpMlWEf
HqxTqKrsrOUQeTqkKoiBEpwKtIMXpPHybO/pLH7e66K7Y4t8lvz5+fjehHqpHebe
uqa2O7m9PdFVKqhss++TnXttSDNDa03gYXBrTU8SvIh+O2yGh1+Pg4aSEpFyN58X
Tdtq7KY8+ACgXgSKnXZcvSmkQ4MllqcilxqfUNmkQPummtXtDq6PvlUawFHNeRvS
+cAHEFrZD0Ssd7spobxF4XSwatkN2d6T2Ez/6wWCz1SpNN6PPw0+FdEbQWIWUTqy
iZ8ryRIOFIt9LARNULr+mb/sb1k2xNTr+DlqNl8TH7aOtzMRQyWwwnz8RO6IlpFl
wV4TbnsGXU+JRzDNtpzHd2xIczGALKiVfFbuEPINj/f1cRDtna5dgqocbzMbs/mf
T4H2cOOdYxpYSWfteRPdz/xnjt49mHbUzO2qlvrMrV9DAR+FsoCxI2fUdAn61EBt
2QMT2sqJG9XUIRLYreYwjzn09kmkCL4QXYTeGJ0GDbQ/2OM6G9xH/AF7VDrDD2ef
dIp1BWuQizDmb8fA6ee4eK/KqmSmhDaM9cfIIIoTaGjsWzqSDv5Ye31ct79pOwNl
L7tlZUZKDJr7ago0V0cpi9eFu9F1N6MH/Hi7Kl0dljpJNjJgX2CAQgDL+i/C1IyP
JozREe5cGf0Q6vecovp1MXXPSgvJgz9RnyjQTZG8Ayw/nt41u6c0AHGIyHjwKuYg
YxWIs48yJY96YeMY3OFQF3vGkFbr0E6gtNCW/Wc5pRS2pPtFl7rahLkOTMx3VL/0
MR+KLJh2Ym5SjZntai8mIQyEgMuYdL0vwV2tnhMWBSIT0RwDcw9jIQMOu9omLoV3
8XPxB5ZZbBoUNQS/0QNvAYvHUWBM3lUtXgFc3x/XeykzL+fujEpUqBIHuYQxFvNS
zqM7gY19FPQdEHa21z3V5CRpZsLYh+OTTRb5OTXklB7aRfGFVvqyjSTV9Xr6hEGo
GqIeKNgdcs2fvVkgoVa463aG5tvcbwxwdMQggtEN2/LactTf/GZNeXSbuWU9ra4v
bKdCOFVOT9imCUgdmU5frwjm3Stp9TEZqcpHY+ACGFQzmTPkmfgLipG8SDNNkrGz
DiX8vfjqtaLr8MrqoD+EcL4v9gttWWviI6vZBv2unl2L8+doxXZO9964hURLfMr6
wtN8BQDI1LP/TBLhEj4ILepj7bhe/MpWsS9mtkwguY2aVVhdHTP2OBqmqdt2o2JP
FmTziXn4/GWpQoibdyseCUiND1i5zLA20Wfgc47HPjhP97epxe9PFmzBOlHXLl1e
6zmf9BFUMTfXyktbn8JdF24NKaWvBAp1TVAnhecGDbuXhd7ZiCD9mCjeG9caSjgP
H8ro8h0J9G/YfbrfccmXofdNTqF32OigHdCdqOZnJ47IeXOe7NEh2Ww8tOdZwOFa
VpaAf5WSFL3ooX4i+79bTLiNQBadmfBOE+5o1OrrrOwGrcQE7VCYeFVVQyZXg6aA
aJvTLPwLw7TnIjU2nTr2sw46xIVmTGCV6qBLipTq1IoRKqrtgEuBXc7jWttuBVWm
N3rzc6lubh/rLbbei6NiEmDt5MA8bmwiH+vrNt0od4nY8HweClpwUiWtT4aSpEmI
bw74F1+gh6u29/4DQzSwKOx1AOmjEqd1UyKzQG43gLl9fVvGnsnljv8eyF/1B1ar
kfIUjWthQvulaEBQs6GFMH/3DDv3RkCnCcZ2KNFBM489nuYxeG+voWuzqaGhCATW
MthZNXHqMUsTX+PrfIvMw3+CXq07YxhaW0LX8ILoDsKN+ICMfDOmQJYaCt3IDQRf
JK8n3HGc2fNJWXi3Q+nFGWBdvy7dmQEp8P38hDacvfgTzfO2DInBQCwFdVt3Mu5O
QlPokepTVHFIa57XFISCU1u0GBQQU0xq5zNNZG6fE3VncgQWQSz4bJ1zhjbS2Kjl
cvA2qUCkWDh/uwkslSQWgkptFfoQRbXYXuky4nd1nY/NSfd0cNkYEkiyyD/RPa31
8GYRfHqwuhDnKC057KwW0B/7aEwWdO6cyT+TVc/wOgkzEOJPgzBbW0xsIwKP+muY
fBX5jDprEYGVdd4YjmxWaqxvtWbi7Sqn3p+nRDoswLKJQxc25mjvak5uCZPdesUo
C24ytRclKTsEQSwvozXQxoiR9SL19UCY5BlZydqWBH4jR6QUbc5lgkd10OJDq1uJ
S9r0sZf7XTCFzWu5sAjabPn7SUYe5SOTV93i/z+zXOT8VQKnYIwYQvr3eVxK1yoZ
0haI+/FoaXmIGnv4oBh9EebQO6gtIiBWcVy8qOSNTWDrSC2Pz6Vhwr6/Jq3M/zpG
dkDEZcdfD4P3qfrQDw5wDVsdh1B1dMhwOhSOFC5fVCkZ1VlCPl6kQoCjorStZXPR
iCOgZ/dDCVYrnXp59qlCXOLP2sD1iUUmSBSdY5w4/v5SCRcqDRd+wyUpY7ZLx4cA
/GDPuH8u1bOccdB/z2Q4FWd2Z/FK0sjmyxyHE/o7PfxQZXNFCgPPiI9Pq/DtI3QS
a1IP7/V1hCEIr4M6UDCyW8WOEo8lIvTcD0xOQF7XDG4slcESDdb+c9aYqxOWRzaZ
jBxIftIskvHlBK9YKCkhynyvPf0BLmSiuyP9Z4J06U3EtNzHKoEmFTm13ateUs1e
5mHokProN1EeOiZlZPQ+RarhX4GS7poGNs8xRw79WbqnfByo89IegD91UhXU7/q0
e4Mo9Mmgh8uOM/OJuhvCl8cIdyVMxX/OswIOrmtFWbTl3tbyS+h3fvZhorxnS7bi
doHoc17mf+fMpyJ1KNFzDhfmpTWsz4+lu/2M0xO5po+jUpD/iz4RRg9mb6LzNWQb
sQNaq7wf3C4NtFTjbuHeCYxbOd9B/S/VsDrSh/VMPf3t18TSsnSx3CdXGqwON6LV
q0m1fjbJHm4Ai7VN+o0267wjrjWZPubw6hbtYFa+aT3GkNlgilld+Um3sYqdycxR
FDeE30WA+/4SSJzvAsVt6ZXwRfClbQU4Stnz9T11zOvME8Ya9IVYwdX75atjv/6t
XCzJjRzBnQq8h2dc7M5jZMMT6Yi0XpzZWPUlRQvQruIrN011bDGk6ycdO2tmpw6X
7PRRd8DwSZACfuTeYDX4XadTkA969EnBUEu4EeX/4HsALvRkGjyN9fTtqxa1Y84d
6hdgZjrYXCLXZwENZx9y5igvJSYsM6nKTZ7gluOiPVkcs9L477ydnIvMuvJPEr1k
q1FJDe2rSkfjGInGBRdMu2wDuOmP3YPEBgdVx/4Jt2qKyWvxPhZjE1jnJXRR418x
eBUYS8RUofwZh1XumI86GX44iFzH5D9Vub4DAcoqDFm79CHefcHFG4DyfJI8JEre
QAbr2yrR/GZveVgSgt2m0xVWmjHk/n5+K5h7o32/j1+l1K9958vTZyaoEDrqCjOG
m7+pc9aVFoZNDhXTRAR0sxnIoOaR6GKieR1XuuvWmv5AVFvHd25jnETC1hpkwp1v
LSatU0W0OTFKSzGlh1FMkfRTDxCnGY7aEinrV35LEkT1O0XH+PKoiv07Zz7NfhcI
Vzt3XWth+J1MitXXOCiIrVfd4KaSVC57bI+vaHuxbo/IxqwyMwVtrCp/fMSyYN5/
/w9eAQVYhjRn4k1JYzNqy7vJwiLRq3KzrnBvx6vY/GcO4XIEVNa1bd+mLURhZLnf
gbVofEXkj/D7e7KTGEmrHjVo79wbNyjEkdSxixlLxtSiBI385/8gs0oEduYlp4Rt
iw4yPrtwJKLu+EaHZDOgB4blMyw7cWn014eHoBOIdnxCQVLkdy/zAm7aaw7hVz4P
sanq4jQ8R97kOJyBx1dz/DWcNg2gXaHxhGeLWPFf+8kuxKu50PpGCI3nM2ucfFz4
+7+jZeanyquTACjbLOqikyPc1D1/pxs+uDV00ON32ZOqIPp4seix3pyLDou8gywj
Ecs7W6+nYQxyNzOQNq9nbvoE69tEmFzlv5YbM/C5zgFZKAW/gwZ6ofwK9PCH8774
7JB0r+YoZUggsb3vzdhfwC5pEMPVIsI7YH9yvhbCHc0F2/eMlyFPMnb8EDJUQJxw
BHiaQAtqMXD6sixV39sd7rZuAho+ag19RpEP5yQdVXCtG9ecY2i8a3/F2GGR/bvn
CJtwZ4ojVABDefsRKVVstuAdgPcH9zAsXxWSaKLCYMKgPaNTByzuRFCIMyjJLLrX
Lg9Y/WIkS73Fa0/HB9/lLZk7nn2ghZO/7TywiDafgwDaIB708c5kH3MjdpTinLHn
koq9gUDzU8K3I4rlcnERFhpP2UIrzE905AgKl7QnC9E7smNtKFj+cx9tIX6osD8Q
kap9HP4zQKB9wr3V91+9LDqtZNJip5Pxbfr9/clnjTrgLxXiyK2vMe4351RXjo78
HcvhlfRx52E0hI/DemK9nQFhbPDJIKutZcbCAAVW2OeZmfRT/V3CjPZSNTPpEVX2
+x34+Q0tAnP7hIcrNoEbE6982+Fkds3jxlwfXi+q2GKMrTR2V06BnOGB+otkQcT4
pVoVLoaGAMLM36dTGWU5vdbtooEKLmSFnkPUp2WegVIIeB2EPqZZmIW5xHzORKhA
BZ8fG9EmsoVb4mWlgMkKVQzD4wIQe6wg+Arwa8v+8KXVQS3XIXolsJi/vdOM2OVS
rwoRU767xcRrYkaP50vnCciWjpVhmkdkiXGDgzbOky6zPoQe1ZmcAbdelKsCQKQ7
9NutOUphamnhsIfzNEuoTlLJ8U7C0r0wqE6dKlAqw+zOZ6jTpEn6t4260tXtx+OH
kdKPSOFMMhQpK1l77UUa+6RJ2p0g6WIa8y7IF3P3skLWdTJeUg3eDUFeYUAFlHMd
gDUdmB+LLDGFjn9OcLPHxWHIeqM4IswabeGUEexTb60HeQK8Z5P7Y9wFfeIQA+y5
7iCxCNGiKqDK8bOw7mLJVME+mWrJedoPMlonoHI6cyzrNQaOLdfsSW3081vXMF5R
45S4YAHvYK9zkN/oeZBPP51gQLMqhDn1T5C4vAdEXsROQdpCdMzOjLOkN4pF0xRM
76SuMFZqGtlQVxR1N3pVTNvFwbueiZFkwe7pgfaDpzrCd93Xj1nT8N/prWzV12Y0
USxKndFOzuLaoJPDIQZBgKtY6dbCJc7hv9SDzIZHYbqLttbExm/N2KzeDvMlAUmE
ITEFedrQgdaJuXM5WCJ/XW2Fm83LjG/rcM1lxm+bmUUVNi3SBfNI3x5o32MwoRnG
1R+cG5O0nyTnWn0xv8mZKSETK+D6fiDmtc9ONFJFEzT8qbZEAbUWaPpfy5du+7BM
/LX6TacKxwR8lP8mHFK+XeNK2ci7/A1pEJGqVWhVz2mpmx6lF1RCHxV6SKkRDwpg
nioNXHKdxiX7Vt6jqsMWo3ptQge9N/J2O75HAVDBw35vZ9f913OUg1SDHagd7w0/
23TSd8mImjfxP3LbH/GJ+62c4S09TrcHVr8lFI41tTYIs0rL3z/Z2ywEZunR4MMo
bdXfmlpExHhxO3b+df6D6Y4xzL5NHi6kzgkc8Vd7Qxfds7dLBrl+Rr4whKtDHFfV
IsJyeg4O6ySTVNW6cyXy8i5XU7gbLwTf7EH2LPHthBVeW/9TjSdgZSEPTZk0mCm/
k5getAo+dMKCGxyIfGsohkCJ77YhMjcqqICcfsTD7d3W4MCOz2EajFxgY0iXJhGT
NzkNuZpmRBBHPpvRsHb2QMj/N/h94PKbazNJV+gQygOP23xffX0NapYpWmM8Rb8U
svRatXXCsDlc/ETAtVb1LE0MKjjt4oDOYKk74sldJKZIIqwOERjpBSn8A4iHG33q
C0w4WeOcl2MpQ4MQQv5t0QE0WQT9QD3HRV6TjGOyitghQuCHxxRoiPBENxzWmyKE
eMP6NlPv2oc11DN5Hv5ETyRTn30tckTYMJuicxr6pjBkwNFxX/u4szKq2cIl4RIz
DjKWNh/DBYHdzf5fgpt20WS0YEEOnr27bC+kzTfR+I7f9shHCkM//mLKNY1LCH8/
IteZfwwzAB+Bn3Kn0OCWaBugHSe1r6EDbmmxKRtQBIAFMZSSfvf345S7xTCG0Qjp
THzJmjyv+sQ9AXEpg+18OII9T9zJhiHrBHPrHmN/JyOT0u6hMDRjnYggjBbjZcxv
HIW/scco6tdi1TbygcdcyIql9rs8RWOrTKEGiVFzgX1DvJ+rq3EUkeAP2f3EVL02
7lTcSd2L8aL9Hs0Pug/Aj60cunbODmaCqRZuNu4nV2Shtje8PWes54xKYynNt6ge
JYHiOhORs3YCD1ME6n9UBk1DWT9P9rM1OFJZpqfrfdqZvVXQUuXLzQlCP3EHXgSw
VfvCkj8ma25HcREuNveriyT6TirLbVDB0U2J0rlQ2shJlEkR1iAbUii4IePfJzkN
9QxcLentsYWth0EXlfcKGQkHrh9HmBcTPdku24pi7fV4Ihd60guOYnaE81piA7Em
MJW23MUvgtzAj9da6GDxegXf4n72YZQNS0JdSxfAJXBBVk3DWTTBxuCNYZ1vPaea
zd4XZrZ9Fg12SOhGOQD6D6CngOdzVmiq6R73NB+b99tVQL0q5ah7Lql3FHgQv5k3
tRIjyphxINI5G72KUFiQTpB/sO8lqalSVkwdlvt4j3c4Nv5XxNUQIxt+2PQHuVtp
cKy137kGGCzwtsPsbILE3u6rKDhEh/biuRsmyAhYMAISfDegnfeqk8FzQ+/umRgD
JSCemrh8WzbmK9bXhkYJie86GFUiGAzIJ1e1CM1rIhBvd6IAJu45BGEqk2rtdpI4
ye818j/GREfCAjS7SyJMI1oy/xCXg05ZKJWszF23xDzkqurJKdEY2mdsYQPDEZVh
tdCna9hUyFxeRkm7Zk3GgxclPrxmzBeXBuNFOQi+hDBUsFNxjzQE+IDO9hzo/URf
h5KrAlrBgdmZ9k7eVZVEsFhj0Rv7yPb928qJM77pUrA9vqTZtUY/r2IVhjAD0FNU
CwalR4OLwZJUsfWsoUY7ZM9OlM/Cr8XOvzfWaJxDo0fg+k8PWlxBfuORBe/zzPIa
Is67MlK6QWHjJdkZnZHlJiNpNRQMR2Y/nC2/Q+it/cdaTroR4z6/uujn/zWqgjte
Ke/0YQVrb17uRTFFlXjhhhnCjjw79RsZB5SQ8nvyY2Eqv3ilMl3vbD51oVWuaeUB
1e5I+OPx/RJdjweZNQOC+18Jog9QLLmPC9WfitWbZ+UdeA9NNS/sMSirMEvG+NQ6
uMzFaLq4eVZJwHlvBvXRuP5sEoBa1v86683jw4uWUGaQXq4GLdUUY6U4wh5gxWcT
M9AB7bWCBiunWEHmkk2N3UkUI1HYozazKd8JxjnqmMVdhEOQesyqFZIt5GnHRMxd
G7EuPV0RhbOwUtZPFZ2xR14OO6I5QZsYLy1uGtdEFCASsgpb5RusxuxN3z0Vm1gu
RBrsFZTeLus+UUtyMNevSY0HpXEwUXakuAfqwly3j87qFTmUi2K/o95RxwhYhYNc
8DiavKeiKSlu7hVSY03RtCHSARDq4HYChuV/H35fh68kQ7Mr0MXyIxwO94+VV58Z
WOk2mIQAL4L7ID30IOzJ+1U6V40pXgLkYUEDvTccKRHIClWedJGRw7GPAVTWiMNI
yQV/UT/CGTubJQAVwlmtfOiRdyteIkWQx0BmvOVJhD7QiYycAZa/3qhNZuMGu9AZ
R7bPUsn+pigs4JW+APZHb92k4Qafgfi1Ig81FL2EkjxqwIZZbmSyq3bzzG32NrcY
9hMztYAsLKRNmKfzDn67yadHB5kU+kGJVJk3bqjPxbluEPNVkuHP1GjmCMziICPw
2UrzSxF6UpWHqajgndkfA41u0e/XMKgls+KKyH3FjZF6SIEHVlwv1pAO6J8hP0n7
cs1rLBSx2rEJd4kcwLn+WL9LKe/7utMvHL9jOAv6P6hTTyzA3n2dA0o+WTn9EcGg
+LynlV4MG64mMOO9KLB7cbO2USbAez9LZlfXUc+hVwT1wgqzxe1tP3q2fiiQIwtT
z3Fo4qfPfFJ6O8q/JXZY0dXj90KIzTCAlEG+OwNE5UXPaQ9IZQ/vomzcVi15BJT7
TTDVyQMmdPGTl2Upah/WtA6a1Sn+OyoDY3W/hYgl6X/k+02JUr98ZYpRzIVuGS0U
yiCvZWQsFGj3btixa4P23CEL0OMNB0wpKCSJWuuPz+6OEZJUFtPA0pNe4xS70ret
4kbM9kL9DxPpGO7Pqo+6bcY8AJi2GvoYgStP6Q/yh5AUjH9C805alaBqIlQwzoop
4O2MUFPaSb8KM1EzLnrn5s18mHB6V4mqIduDJg9sFf7zgXs6YOtZIgHYzyWquygd
eAUdcZGk2N4mC0bnbaV8YJ6bxRV6zjy8rH/sVoGpLxla6c8qX7kGGauOuYbbYTvv
o0xi9e9ZflddmdXWqkngt5FKId3nRyo4oV3URkjeZGS8i4khJF1kLULy5vTeKl5K
caLzTgseuyRaebldAbg77JiwEDAqHaj5QLceagnT9eccp+wSpYajvGVsIYTXonX6
mZV8rphhC5C4iHe+rrfbGIHsN0cMSCcFtpUOSYeg7rPJo4dikCd7SC0Rd6sDbLhl
RMwdtRMZ+8GWKhedu+8w7UvoGHa+7a8VT3hSqNry8BgKZ/umIufSPCinuICa9e9l
UiC1OQBTlFiQeVyhc5UZKeK69PkAbs7z9Zrgg9kRd/sqsa2iTb1IB5OL3lm6Ae6u
+plFMonZKAfYZU2UaXEapsdxN+nbDAsnfhcXlhaar5oiW/xNVGVRa5Z8RnDRH8ct
VQ06k9SaleNZEOuTuxfs54kUTtmwiAyfWE4mOB13YZtuXiRt6YCpIj7yP6yd27qG
xSTrmOzoNxmhkKF01xcY9DWEEHrAcgN5IXgw33qDQtzNNjFAM9lFfpnlMel+dptT
lxTNtNQAVlEpXeA5eRPgIzEqjLV/sGo7qi/JuUcGVqoqY8bTvFse9osiACjpLiXz
xlfgzsAtLl06dZs1vjL2yhmTYl4eKhpcYkEgcpG+y45PutSwqmx2MWLy+4PHy7S6
IdCVJVePSZK6WBQvrgoS5mSYObdlwKohYhiCpv1b2HKdG/atXQQeGbtnnpYuPK3k
wyo7JXOsyhDPH4341C8Ga2xufUO2+pQxNKevuZ3irQsSJm6jVEDySNTwo9O5OKYK
xSDWFzUuD84OYW1cPXbFhuqJRIlBoYbKGHu7VVV+Hwj8u5xqxuzGfFmnrvVRfV8h
IdH/Br42ar/D0qCLqlEdgBGa2T7pGubn9QO71OjLGKAIU6IrsnjNC49JXIJlDmkE
l4xl/mrFag8qMEicOxuS4In5mRg2dVilYgPzBym8kfQLrCt+FNgXmEI5OOFYGR7s
K5Lt8qr9mYC1iqzxcmUMZM780kIhClZ7fYCqUeTKz+2JyldexuXY8/2zCU1UxTLa
hOxs1WClaHrClFijEaQ4aJ6rCvOLeUhauzGKDfC7MRSatlwGD3Ku38con4jsRTjC
p3UFvVAhdYY0pKO5gtlGaRYy0aiYzMTwZZPP/YK+5oC3dmUp4HARS8b3ulx308eh
15Q6Hixb1N/Iwybj9e1bfETN7EzZ5sPwp9mZjKpzHRH8TnwPBD3IyKcqRGxoJIRc
1Mkk61bbe51JbnVstivZut/AFQQk7DmFI66v+DSxTYZ7CeX5495c47ILhzsNPtxd
2fhopK3m9CsJ/06yZVWVe+GjID25cd+usAvsHAXIMfmAm4ZPty3iPJ+upcOhUc4W
pvSmv/02hglQYkcWC/BQbxN2e7K8q4V0Wav55JJJ5+7ctyqhXqGkAu1Qvj0XuxDs
GVOB++SA8Y62ZZVs/L2kns0w/yNaNYbu27oCtNYhUCPnTtlKpCMSHjp4mCpj6lOK
foRbStLUJKPIdfMvUrvds0sLHxnPkhBK3RfRmASidVqM8UMqRtBI93omMSaQlZjz
AXi3mJthsDwewFr2FuSZo/TrQdQH+VEVUKLrVbmoXTLVGTspBRPBpD5C5KkQSC2H
/qakPY8nOsyk8EjadCLfIxmk5zwAzjm1jSV9u+7oE2QO25NB4D7vJR9W2P2UTHNI
EZxr9qWckFfx0c4BKxl7JUszU03AxR5b9NWq4Mk3KYrsBFdtxYweRuAuyPfiyAhc
Gj+aTnHNRgTjOCysryWIIg8kV0RYaTyvgxfut7J94QDCArFfL90mR6hnZBhttvfO
CU8AWocvkd/Iv0EO4KY8kBqdsacX0bvjTR4qaSXZxRxQaTiPk8qa37zeUtwgzGlk
SmvurS71RIXe5Q9pzkjYiQIB+X3KGXpPWuu0O80/HaqZ2oifV0O6U9NN+iOni6PK
lMp7bOgceCA4OEdYx919ok3IxQVypRLzWxKjnNlJFpdOb9o/zqZ8fMsXXZMNpg75
ZOr+yjelfafPgqfdLywyETTDRA5i3B9h5gNQTB6D/DvDCIysBWZCYxcjLXJWvwik
EdaEja9X+c+HXSoq4gtqQKXdcY3y5EyX5p4mE72IMdtEnEx1VQmS6dYIpGSVKG6a
W7XBA9967N7kVdnUMOrSJgsyB3VST/zZQjXSI8/9TORcwuOBwZIsD/3ObyZmVipX
tz8OllC9Hsl16z1NAUCQgm9aM20q+M4yiSv8eQp075OT7wCi3tOE7VWa6QYmA6Ci
pmipWJ6yxRhg5WdNu1DwQtsXHvACpjLwzOhK9JsciaE82rzjH9JSKgAjqbauN/LV
tMP2GC9tNnfn3Tg/50DqyADLufyXGnd6q5eqWM9IrAoxTFPcX7c5jFsEqzLPH26p
SdgI3DgksLxyuPR4p2VuVBEHdj3kjxfIIy+IGQTnLXns0So5IeiZsWbWIF+5yv86
XbGgDdH1yMu0Hx4nlwTzSPeaqeG4HC4zfBnH+wguE4iO89YF3d92lPa5NAwQwLqm
8tVd4IwInPBFhtYY7JOoG7HSJF4FHrBb5Xan2kPjE0LOtlmF02/P13cEwHp/AOup
vU6LIQNFPm70mXWxhfowFXr6J7BrRNWLWgUj212YZE9KnTw1umbuR/Hb4bARUA43
g46aKGU+rJ8MuyNCnUv/KC5kLqyXUZkZn2Few0wQop5jlnejJrrEmG1ZULYKQNm9
c4C3hSolv04Jruv11LX+14AlXKVBScJ0+3sfH00etrh+Ogeh+feRH3kIrRfVdZns
bzsSEK4orjTNvCplfilhQLeiRyYvrsGbiB4HLR5KjYzmDJ8ct2L4AP5rNGG7yNeT
sL7tfKwk4EcPxRSU20EjJ3bfo0u7r1kOdUbauvXK3HTBStupGIP6I7/xFw0nbLyo
9/AgDRih+nC4NetgVAJUgtMoSVT9+pAKba4U+rpJjBLnyEgJcAhUvntmCGV8J/sU
cFgWB3BMkZPS9PiHQCctMTQy1td22ZAdYwp9L2Ffz8ADRF0qnhRdLtXv+u5/mioa
8wfihMLLOLhjp/sETlk3zi5jIPWl0Jtb6cOtJH+BsOsiFBNB0RNC7iFotnn7ATDN
L4DF6fO/BD/4BbYXw/Ac6Pw4zJVwbWbXNfxzwLFPXGNFV0aVjkSEs6tLLRiYNfMF
I0Z0+LJwu5iZKhWYo5PPKiT9vvieCxgT+wd3lAYZg5tHHjB88ev2iJfoMMVnon2G
YjjeadsrJV1P7+XdshGNEbu9TcA9XljiaRGsNimexvYOevzYQOsLaC0usSgVYDuX
bY/UtpfQzB3ChLsO4hMnqecD/ivBbnfs/G5A+/wuPdbbccAy7klDCrRLbiWdg2P0
dPZ7YYIPn3K3pdBvRQfjyKjtTxuciyfvKQKlga06sHYTLHlf7K1bQVtGKr8pD44C
5eG4Zp+aQ38R2Bp9Mr3s03E0nXttmEyinxmbYtq/PguQv0e2ycLD3oK8+nhTkI4B
9jY9S2x7Y4NhJqzeT36OiqehOIjhfyn4/IEMD5vt9gEnA88cKZSxz26mfCsp7QZz
FMeaGjJH4iInn1EPrWXjOz52qXpjpkRB+w0pB6vxNq30f1keVQKAlOhTi9ORXbCs
x1FvVDS0iQM+xPQOFDBFGsD3xmJd46fppwNfwWKohWVeoQuXYNSjHQ5b1MNYY2LS
zWdEU6JaMzy8pyjd/aJlDTNDZjIUiW3aQP9WbukRsFTN2YqlKbSQJGHlwkwBQVai
KRkRDrsgYpO7Z2J6JkQe9t4TDloo6Mm2cwbbx3bWlTx9fvZwVGr7CBy3dLMp0L/k
oDDbkzCAH5no0MIn4tvlXtUC8nyX/wxRT/0Bf5NgmQR9kDwmLT+uAr0JIr69z1tS
+Ekec3qRmvuTZ9Iy6Ne3q8SPMOViWsZlzE/QcFB6Ik5F23aY5W6qGSkuHJ+xaXQ+
532iB/7ytBsHte4Tdwd9RWY8k8T3qH1X0fkiYf+OhSXKoPHy7VXCxrXq1cCM2rKJ
D4LrMMsCJka/s4mwxp9CGMMMEtW22ouGHh4Aw1xciD0BYXDV57hwvs7LEBHvNmEa
UNzGr/TZ+sFw4QLCtseg00hry3SarHme6V3wrfgymL+9+LSMXLUIsPh7Oz9/zbTT
lbSrmEAQ4p8OJNg1X09Smq4KwIq6qUbvKSDZleM3tITrH+aE0hQq1TKnA/s7EcTF
iP8XMEEP0J9/AqqGXV4e+VpR8OwQZ7kvQp345eikBL0Dreji1j3E7Z0m/8LaqpaA
n8vMFFnsBcO/T6rszKlJfAHmUcOr/ucjeNJPOTFVcN5L9IO3KfEtBAGrBtug5rvd
QkV+njKHSfP/Lo8WWJQYclaSkcjdbQtrYjsiFRILkKhNe+u/VTEoN7EEVHfMW1If
h4PXDlfIuN0rP+/GQNOOx8TVmSOcJzPDhEj0bngTK92pmw4tcbi6pUNGH1btWxlz
iqL8o04t10rNrJGXWgo18F6F2RN74luqbXNHQjrBpvdgMGANEL12tktR1Ye792yY
HMK9jQe2dKRigbu1LYaveDp9fgH41caz/wi3Tb/Q23ejRcpkHgRayh7WegqF46+X
1jquUHabMb59BdMWz4EBxGWeCUKav3kLLZPRJDnCMrgKOVl+3o2ssRYXqeDf8eGd
mUxD0GbqLa91sKfE2jsHfQYemtyBSgLB86YCDniHdxi6TjrWVWU6IEgMFoVNY2Q7
09ccRNfRl/WaOxD14A9CjuhEI7vgtldFnE5Rfv/GfBBxyXB8dLa1U7tKxcXjntmT
bkIKi0PxY4AKFGGk+64LFnsStS9e9CC2kmnsewZCO+DcyMglhjCGTW1Sa6uDr1+x
CfYwLtA2A5226wkU5T2fF8OERmaOUgijrQZDH5yePNNYTPccgjl+xNG8lvsTbiIm
ojMuCDc/gprJ1gWbZ9S8JbCG3buCueBV2mmvexsY1E7P4zhEHB6n1bD4HOoGy/jD
53YEmo2GR1r470SOr+AgIMkeSSCjAXXZc9DlUVJiVnZeNcIYahUGbGq7/Mwwx1E/
LN44A1PosL3rwkS+HoIF/c4THnWdPeQmHgrWBnMc/XTERQHsJsBrWl9opKhMbhWa
NBcd975tmaIVEAFBxkFNHQfQBppFkpO2eQP6aLPc8bNHidGteQOCaYkUi/fEppTc
ESGFsLPx+hgVEzoC0uFatz/RdmBHgKCH6bYBCJGTECbOL6raiVMyVYqkodLnNEQo
93Su30FXBmlzB1/58p7DBF/cb0CEdWrc1Ee8xSXNNwT8oQ/QQcn+aOPLO8RwFoRP
oIK3GF88tw3Bwe5KthJgHsGjc8+UVs0inwaSmNMg1A/n7del5sWeow50kOFczJhU
6txMDqit1fqs1HhiOOZvlMyA4UpwieYbzcQ3LhSjkuzZTJKYLmh/5LeScdP9iXLM
IoyYaA1eENtAEWfCKzNyItt1hyoKhMQxUW4cJxav4HUMhTAVG3vgxoaQAO8iqi2E
9lOcPVdXc9Y61TpHC0sDgodMbANpHe/vzA0HIddGPqXadE7+bwcSAI6NiEHAjOQK
5noJmcc4P2kYrz3ila+upTgseUP4FljuIo4QOF6x5B572/lb2zAEjp6/r/Jw5Ja2
sXtt/16Lh8IhEwhq8EPE2IhjcV05Yrq6Bmg2YN0OdZW4iaCBdhM1TLuJKb35vqQa
vUnGNOgLtb/fBAAxEko7lWSlCzdU6Ih1TxGLxqyph+IKkBlvBq4JsQgF/WwZk+Bb
GxMYQNZ8yxrspiw8jbeaFONdpk6hBfej1LXSc8mvPStDOyTWvuNWVA39anTiyL4S
9a8JX4UR71LqIXux0GRkR4v4Zcs8F9KgZjVZqRPGR0BOKB054RT+7k72hhX5Dqg7
GLLNCz9CrbukUkOv8h2KWaRcTLIh7DNAME4okkdAyLImyjIazD+nSBMqICXs40P2
DQvabehMNujI6gWdU4/M9UzWcTrvTi2IaN409r66+D0S7T3b/pGfF3Oe/7w3LGL9
Ejh6VamCWm+cgGzYY75lyb+fICjPl8AebKjgUk2ju8RAYxsIgK0zmIWzS6bK9j4V
chkLC9fdLitXruE4+qucmXQECyBfI40hEgsF15d35BA57aZYgsbZKOqV3b3/scO6
5vup6hxJ2KpwKuGfnY01jM5twqI4+QiYLSu7F78Hp0qBhjXXV9bT935xWwtCcKpv
i5fLC3bLOg2MqtWIn+AS6gGtU7Hi4bdroRVSPc0u21GbcOVa/0LK5RYouGCkKmtX
fAhZ0iIO+PzZUac9a1+6OzvNcc35Fm2it9T/YXA8hbB3k0qCBwSVhZdySzAo/U/E
20HbS1Im5OlaIRRN4y0dhJEwbVuMnih1IRVwlD1fzjMpfJV7RqFk2ZEoTTMcr/qR
6d1s+mvz3YndWPPiK6vD6EpbTOa9gFxXFXAmVr/zFxsIFMQW+Tq2VqBGe4OyeaiU
vIRn3c7nCUUVryjWLeZXD+NNXidYoN5ktP5Xf84oVD+NVwriVulqxS1sHr1e97d1
Tm6Ix730DEgEhHNiUpOxgbGaXaGTUBJUfGhtgQiuQq1lhGsYrDIdNcP3wBvMfkJw
bY1NjWsy1M7zKtR9SA29pgrTJUggM3zOQSBOI5zqXUy0XWrataV4kra1vs1iEm9g
y/tGQJtjErcSRP3n5hSd42VN4OD2ULw0nnzNHFQTwopFVemhGoO2BCaViTcDd1tQ
fwkYVdDfisLhbcWAIfLY8LFo1o2EC4DypjqWEB4+Yh69ISaDFpn+xV58T1YWktUF
nXU5ilt7dp7ifhi+fABQTVEHfXEdCVTz5/j2mMUCKxvB/MC0yR/7ZwR8IVwAKVI0
9DqduhcDKZL2gJErCk1x/BtJ1NXyIMp0IfloOilNJbTgryAos11AABl1CYlv2hG5
Gv69rznBiUaD+wIapzScUO65N9bs2qThFo+hA7oDZ144jsUQPKEGtph4Q5TqptXY
C9WBswVzPaLz2bLM9q4/EE3km8Kc3ndtIISK9C4bFPJh9U7dwn+4D49rndnmXkVq
lOI4sDMEdBZ9XQn/n9eTFabW4jryNRyBxlIC6GRe3ngGEY2UatEYy/sVzEwXXEn5
twmS0fo1mviGrC32LlUhzvYKIOHarJu9ncNpMudCgcrwf7encsXzadoUK8ZDOUSE
7oDSeGTFJynlFG7fBnarWZ7QStc0fQKtctuXQmcIk0GFTgA+7Z3BUM/vDIewl/io
uYre9kjKxK1Gb9U/ivxslfDymsg3vUPR2jY38ynh4mgg5q1hssFT9vTXgnpYQLAi
LO813ZQhsBVkuDtW4RXg06nuX5gZqBdaBiW3x5hQ3pRQ1+heZrPG5xlmVo5AqFMo
DSa/m7Ydj61PSVu5rgFIASCD/6xA1pDElmuSho5dE0B6Qag0/l9mnZoy4NDatWHa
uDYWQygGXqMqFHN1Buvy6l16DnZemz4GiCvN6PQXK+FxLkM+PGmJ49xBfT2Rn6Sw
EdqMSOVCfvN3zT/Ju4GA2IKptrf1c3cZpGag/BjcuS8s08EZSA5qjDGhW7y25CGA
YZa/YjZKnXg7OO0Lqv8G0ymzRil/lanpgunYhJVuQw7ql9TroIbyy0QqnfholTYg
3NGar9ESWF/Uq9y9y6+aoJ8dZ0gvSL3PQimIywf5t4kVW87IcAdzXZ+ScKhwywut
1+cE6VTcoJhP1Bn+bQWpwr+yE7clHZQrUPZvRmhA6qgFbieBkJkbIMypJDkOT39J
DUQFWEXVgJaDIcGZ2mZAk9VQKmSjIDMYs7x4q49BDK9DlI9LK/eSbKxb0Vutl+fv
h7iiiCurVtqLTwRNbWHwSGqxRagSTBu+hKFLzdR93KaPNBZ95mpccE/p8Hn6Syqr
EXvDPZmCxcFrVR/BquB4UXf6cO6aAwVNBPx2MKXsEexNDuqGIyBaph0NWL+HUo72
zsLMyjmtDVMNbLJ3qozIxnXKZb7qWystOA/Zvh4ThE/vpHIAfVDMRvbBJjsfAQOI
2WyOqk4g0hrLnpFptzpj9d4A8Q1VhlXgLwru+KQNtGmJAP86ThlVAQah5vanoBkH
KFgJqku1mkBQ97pcc/Iq4+R3sZhRcWweqglkxb92dBllCa5vKT6bvi6J8sQkuNnA
pDeeLZBU9jUWiRjxPwbskThRjPfDIaED4h8TgPl9l+mkDfP+e6UgpkFwau7fzEeQ
QF2uXQgiradQFa2YHAoUju0oYeEsRm75icyr2aQ11X1pOljNDs6wnBk7k8VQKUQc
UHfTfx9gdrsJ9FSxO77EdKMnTc4QBhzYFanr7SzrwT8NbmZc8rd974A9+epg+W+l
tHLmo4wURHshlp0h63TbA+CytUli9lZ1PD6aSMiqgduNe3xTCd4RbR+jbpTgy5XF
ArkObWN+vlMekKE8+4lkyhyE9mU2n9FmcU8KQ+u85koeGJWpTlK77Hs/JdqYKXy3
aVTAlrwQeHJEnxnnA2NF1+xl+smbsCdazxJUnCU7qs1Wgf77ab7FROXHo0i6NMCo
Ge7nuNV3lNXlwpPRdFbEvyIrtoHwQwY1AaZTMJGbUnnzqhgSA8zc0fF4I+YgEIqq
mdcogSgPC9reOYTXzak7sHgix+X+yhnjRCfi0blN6SpBs+J+YMZ9YosHnoVjfobq
nssADceIoffkHJubp6rTJykAzw7OAhsW/wddUTn/v3CoWIYNeZvFc7k01Iq4H26y
GgoM5TvGdEumm5prS/gLKew1kCIUzmvg+w2KSY75dA0CrKFLva18iimKT2FjmXih
+y6qiCc/AuYyb2QfDda10szVRtNPynd8Dr/DWbGIPod9xA1hv7EI/qGGHM3oGbOy
uHyJK9702eRW0XCrd9oavvt7iSZlvHBERmfU+n8cm6q7LEGYTveN8QsxbkWU/B6i
Oh86IO0VFhKmmU1sDe2HjdldO+Jam3mg7LEy0tvmwwb1j0MIps7KQ93Iab13If2n
UATJc0+qBVLAYYlenEAIRSUe4ykr36p/+9h3hqSvWJLpg5qX7B2AvUJ+6IJhxGCn
2UR/hWAhZcG8FY8wU/TcpeoT0V4G2jbhsj7W7K3TmrOi7GyqeifrirMMrfvXA7JW
0DCnDZeVSFvAPx/4O72bDGgvw27J/CZEWZDezimbCFQtSo3lfk8T3+2Sje+WyVEC
uDK55pq3eidYi5l/1Rmi2AEZCrKY/fudBPJFRJQozRELIAV7UN2ZlbqYsEzFV69j
ExSluFml1scQ+GptSFp8Kfnt6EUpeWW6XFfVqVgAhifOfmXg+1O/5zecmKnl3lhi
FVhfbr1ibeq/Abhc6vimDPozZSrLuGjKCf/6i5E1XDUyLcSEDSPS1xush9b4SzPH
L8kvz2nsNnQelKWYejcnRBWqmDbPWjOTbSfaLp3W0tudwPfxSBqvHoHIw1pCcLC+
pCAqfkfbLYXtwqiBbo5WJpBMkPlAQaYsbeCRKdwYZgfuwplOE8SM35+nm2wUtwYS
PtSJ0vddrpFK6Z+tGR/1LLrgHGf6DHUGWxnegLhlVG2Bv0MtVEjk7+G1gTTI6Pq3
JJ3M2ZclQS2P3L4RH8M6tPqLx7HC0uQTKh4f+XtmWMDsJ9Ho6mY0mixnbk+o3a7A
H9gTB04OXebS1TUCwb2lWws2jXs9tiIraTChGd7wv19ho+C+YivRyRML/ZZOEMpL
sYX0u8etlIk34jqdRlQPLda7n5Sb6k6XnX6wcHhzlxzdNM7W/l65DqCqsKDlshC7
SLplJMWJ+wqG3QmK4FBf2XtDSmgI70SDi/NDM1ivwZ+zUxSX1YwZg6q1xpnucIhV
IPBUox39qtWMAcOynVX88WX53dWehmgDOqQEq2RLmlk7ZMp+jK1WAgvBZMVRqmJ7
vZZTyr2L6LKaFfLo8G2ahXi4iZvI2NLRHqTlJiFZmJk5FtyITaeoPUmQybxBOtf5
7cg6twGTVz9/BCQNf+THUpEidBh6YUxHSAX3ZjtnCYVx6y/7PT7McLNw1SbFYynx
wD75CbvtNd7WFj9wx6kYAPu3yPPtIVhAftHz+3jssSOo2HCN4nGGdjaCSQO03GXQ
IBDckN5viTyIdHZHUzv7a0WOnGIFxMOj4UZdZjzi9jWWLD7q9mU4oqtegCJq0mpO
ncffzMQp1cCGjOQvLBAkkKLl9eywYLzOM/4JYfl53SyAalpE6ptwW57WOtz6PJqx
Nf6NfJILGOZcmXQiGe1rLfF/6we/zWesvvKVrmtFKTlPcpAfmgp7vOi8FhjRAAml
vUclctMn3w5sEgKT0xJPjC2IzOvWXb+LG5KdBclUwVxEB81aYpbxErkRXS8sWStt
E6ELDZ3GW3HrOb2d4xAhGd1hYIFIUDPczYlKrb9RLLNTEDGadVjTB764im4IaX60
MX3Wn3QXsHv3To+GsQBNpWC423QeVeBrbGPI5C6qgflSmCvXfZU54CKUIds+cmwq
iy+/7K9BC3lrIRWqcNZuO6YvjzSsEhdgD3yLPRLHUtWqhytRL6Oo+HSEnMoQirwz
UACus1x0hW1EZWHwdL0+Wy58bwpSFFzZIb/oVvgNtfiPMog3gTJGCb9cOJsKVA2T
lgNZtoGm/Io/tmrdhKMbEudVFk07th7HFxH/lc84Ic6swBvUqR9lMOwBMdlSJLat
sCJWyJNdnqVr17VLhksb/2apFJZIoP3i18qhY0EIblWD5Rq+AYvle5F7kVw++lcX
RguA8w8N96gWPPViWutStzPtQadZAOitlvPLpVEeYGOODPy1mSlReDPNOUItkIjt
+/Yta+vq5Jum+hdsnvt8JpGSSXq2+SDUEsza+lho6wzpM1omv2fgihSu264q61ml
SX7NY4pR86tLEIZa8VsjOp4iFfy38NWlgs3pnbJ2avlhSZNSpZRCJ2iwI4VnrD1e
s3mKIS/kQ5tgxS0Gxha8Q6gw/ndboIcRIyV3yGYOERTn9sHhAYlXMW0SlOlt7qmV
utx1vTioq4QCLMz9dF/xaGV5qZUA6ypcjvk0B8G1YH+ld9/hacAnc5KEUFuY/B3t
Tr4TK1IWf7GE/lEngX9J/MG26vxIN4XltvNH4IgAbEf6bAggX51xC67Q7f2jeCrI
2raRL5qLn43n7Oj30zIRtDwNT73xjzenSWy3JxT+WMRiiWYSbGN/+Z1X3owNhydb
kFbS4Jfrp/CeCksX9gdYJf9QRQi54AIwOQlFXgW94GSV4oLdil/QskeS/XTVTUfp
x8X+0qCo7OsLURUCTc1NZcxfAif4BPUCsxrHc0fdBUk3oc5+obel3agKqJ1ObLBU
cqkJOz3aIyE/CxFtVz4pv48NjPXV7MEhJYE8ycrszP7YhAGf5EwX0XmvXfTXpyj7
qNBzqNsa0RfEHT68BW0Nhiim00gfEt2qbZWBVbhV1kCiA60FmYXhttb4bR2eeBja
pK7NXCgLPfEOMuZ0S/gY3rOclgUPSzpb/fF+FbjiwIZOmaIyrlejarLNkbxW2nMJ
jmehm4DxR2Ul9Sa5QE8h4nJ6AtQgnz7WAFsrCiyXiaryItKaM3qI9fvK/lpezY4J
o0anfSfOZ3s0rFpyyuaBFLMMDQd8AeI+taYslu06qdpcIPvb/uPgUEsivhqI8gof
Q/axRQnSK5oeK2dfh3mMipUzOJl/+UO7c1FSE3uN/UdRE0EtIxjEy3PvOJ6JXW9X
VYL33bSSFIQEuzsOkCHQ4noDFH4H+6NLucpvpIsOkDof+rYfXgdZvfnCctO5Ai34
V+cSVGqJvzJ0fmgto63jwRZRWm/z9E0tf2DUn97D5aoiaGR+msvx0x4SzCt4XsLg
WZQvLwA74BEYKlFtyygd15HAm2yns7RhPkuedUg8hAcSKjFEYgK0F8s9DlufJXE+
gRFNvEWP7yUJsZMDk+aHnW9/FWQbwNMpuzk8XZG3NggI6s/O/uKZ813+mUBtKQkv
HjL15w/DAoYmwZdb0KxGjcL6Ewqhmyv3y8caUm5XWDpopsjnP2fOqKLePx+KhKST
TPA7psu64D6a+pJqopP5GJ+cnd3mHjdLlHV3dCt61QmHVXuka37HVobCGTGBynhX
5h/fP2p1QeTw9935n1AFr0Wa8ubfu28u4tkZeONMS/F1w9OWl9JcvL/Skzaa56O+
xoxy+p+6aFr5wGQiW9qSvMEJB5d5TB1OpUKyyV3z84iKCHJeeQr6kR8gSNNvCWNF
lL7PIxGc7GdnXoLZewuYG907xhSbgilchHLmNBxRbJPNGJ8mMSDatfiogwlX2ZX7
sesLGNvlIbCtKV5xiRgWsiyLWRXkGgYgLDNUGMsdmVYHvXe9m9Xgtwd+1iLlbFr1
/RfF/ZA1CCbFGyGf5hQdxtroLMkTVE//WsS1sVhet65uKrL67PMkmaahuTme+dcJ
D92qSuSmo3iKYGjY6HoboDOMZwki4CB0x1Yk1kCvYxbiqpRdOzwizAKdUbztaxi3
RbWagLf1LLzIy3tzY0CNfOdYPpahJXhuDcEcJSV8mhUsAzuOlcvcXpD4E01YM7xH
gOtirjaP5wlxq4KhfrCGcmj6a1NIJ3+PJP75ERBGBVSh6ackIvx9ri2ogDNAGkHA
NHLo3ooYESzNTSwCnnUUULlAZquRvoBCd8XgjBR9kjOUVfOCAsfrXwCu8GM2FvSy
hPaB/VSlHeEskkDt5T7zP5GAJJO9KhBakDXmtJHNqNf3ZJ5gVWSLau0HbbEmrFEN
KRA+VKOCdhbMxXBkLfCK5MLXoK2eRsp5FeZbfYh9K7uirbqsVgvzJGCgy5v7DPwQ
AjZOq79gCfThtvpqs16WBamQvGNZAMSd9mwEyqOdC9CjxHeCASZjZyzn9/xKShwU
JdNgy9KryiBjxwYhzfRYKHuQRdNOJDS2hMQzYUJ0SVnEq9vyXs78q4shmkJdP6Oo
2CKnS0L4EozyiYIaEUKbRDYrQy4JAM1+HCnjq0K96hG80cxqUT7U8cU9ojwcMGO0
wn72kcwS45d4o+wx+ELg7pQy81jBipo9r421yV1G1MW+o0dCSJu6CgFGyZveadtz
Px9PuQK78wO912crTkYudiOzo/b2jWtjuPfz222tD6aIv5m/LnBXdkYiqUrewBaG
wl7kbxn/rn7qFZxCHcuC4kjy/fy2LUbrWQm+2QMxHVda/ufgAaMEf1SS8FfI6ZLT
pat2zLXHRGtjzB+D855hExi1yHpI3XiULQjwtFdnyDl/vCYLJmAaJRbA7WxbKL8w
GctKNkvyDIpwOPHG2NOjovwhXLxFErxrdfBSQvxttaHNvUJQHinbruYLu613YiCS
G482R8dBeO6qJWjlU3Ry88+fsAYpx0N4gwVQuvLR+/sRM1RSf5rwa82xZTw3tL3b
eWRB5neUiwEpnMa8qWh+cMrt6PEvVxw23avFPdsoYVsYQUCzwaXD2gTxID35D0z8
Qw7I86cJZG1VDDnbYq5ZpsB5M+x3Yicq3mbuD8RhgjW01QBR5lZFiSKaU/R3KWSo
bBfzgjL27SkPhHtDJl2PwhJAlDTpTouRH4QwkaIgXsBOAd0fcjINWMjUmpWJgAfG
pgHEF6WknRfqoNkU3oEvvjhgMKJZCXHvQQeXjXq9xKMWFFspYk4SJwrsNJDj3qRj
H5NUabv0zymfoHFl3DRgOBliKcvvpiLNz4d82yNq8RLURu0H3fDMAviiyjHDZxLf
HX0c/MeupzYU+376YZHYqxoioFoY2dMpJAjZ1K0beDngMcvshHwdsBZzs5H93OHq
quhs5YlDbE75cYPdXhzPlhoJFYmjZT478lUlCKUtqTv2sxOnb0KZdHt72s6Heu3i
mCynKX52yhqAQZs8lQ2cLu07I+vzQciPEXFWMdI/3bvOC36bF2qELPJBXRc9p9qy
uc63MaagIqkGQTYmdoCA3mTQnSwIFMalSpybeBxQZVjOwDMMcNNlphCJBs7tqyjn
Qh0NNXmOK88tMFA9B7KivcPMRzDH5IGPZMES43Fzae7Aw002FqTADUbPDThF6IPc
K6GTWhUFtyEAsHAeBMu0xZbbVP9WyyFADkzhEvrWY4gYlyafsBY6ivBsscG4vDz/
tG8CpAkQawK9I/L5f2nVyEiw+PL1tugDm2WsmbhWqDtTfTraYcvx4WSmWBaKwJLw
DFUOBoDjw6Dm3j+mJJ5ZEcXjrmlNU6nkU+DQVVbN2lDIKDW59QYPh8nhchZt1h6C
v0szMlrAcRZx3EM5c8xAmdctPvVo9cEE4KWvAr7119w75d0RZMp1diUumETuf5jW
IssaD2YjE7u8tspJT0HvDzOnPTnKHlh5Ch8JXwfdOLRfUPaQgKEHFtlkKkFo6Z/k
cCJu0FlogLTYlb21uHoCpEkf0naE91FjEiSoD8dnjQQo3+Om29TsKkAoXaR9tBYN
Rb2gF+aelsI4n71fkzIAWcaF0U8lCePtKmzzQxJ7b/DNQoa6tFNKhnjsqbVT5ti5
VJl3yfhLyo3z9EveRt0VhCBwCwMGTWDYaImSWVU28ZgohyRHVwvV1Ie/zG+bb1mO
9F/rWDtiZvt/umBJzp9V6DKLuJ1pdptvedaFoD0lh8Aq7vP33TDF4AAvEy6wSuTJ
bV+8b4kIf+HcIVYf7+UY5mCOUJDM4rXhbzFKkuc4ScSC3q2jBj4U9chlPgUhXWNc
wegxMUy3FPQGLlL+sIKXuitRumr4SEw2/kpmmIQbLD4UTQagpFS/vJMxTc6eDVO5
/yqj0p42tANo7FJwpgyovm8VHh9uus+9PYrd7FjkyNPmH0Fd1Cp3LBvCC5T8zb95
VRBcvlW2M3ONx0Nl/DtsT/5oXmNae5GIBx41kFAPPv+QrgEkUOraIXuQljl25JIN
aO33YhvekWaTp3+REj08SfgSRS9RLaCoAFPmC5aVv10l3pGJTXAgEG+VU7a7zuXL
QmLMkNnVCDQ8+AbhjSuQcK9oR5sK2MQSqNZVyWyjBCjq86U1eqf+VjWIw/2SdqF7
xb89nlP2acHtYcoAuXxMWWnv1VKPvUqqTLgwxDojJGG08pV+KgagP4ECFscnwkAj
KZasLt2x92zn6ZYEskYHoF1ISTveUHb3wJO55fDnyLi03+MYMrslHHrcQ/w3f9+a
EqAnhO3l7a6WST+kDj8zQ3iY7tKiFm9Xr9OeokA4+XzSlfGOFEIq/FqukrpcXDQo
erQYYfHPkvprEwrZcRJD8onrg5cCgcEklKYdj5QUmh7Q2hkl85+q4Cw4Sd9jsA6c
2ar/f9QQWLRdFAts4Bggl3WSvHXftj3QECxLNdMlMtDjKOHKY6WJ7riW7magMay1
fNDfpcllqmwfGAYWqdsjICCs3OWsUrsClQfLWd5Pf+CHlFSHg8hlS/tgoW4p+RMU
cGM3Tq7CKbfDHhc2D0/7+WaKncBkWQLK2xMvZB4boOywEu3fyaRKsiqMuXWrUlaH
d+p5CgQCle60p0DwRBnDNrWXZpHTMIkU57iP8hm3UwEuaLqMIpd/szG/7gQ4czXF
KBKNfW/jrv19vdkJvMTbH9ATIBMgKDFLXy0dm3TMWrE+Gns7PC0okCuz7xqAUUf4
kr3aiWzoeG6S0aJdM/aakaMoROTEup4WnLZfVLwHN6pU/edvcOzVcxrUVZUFz2f3
b2gDJwx9NSilqZCOWMnqAjQX+ier4TCEdpC9oJjt21w5TcuWMGOSVh/FL0TjmEJd
eaKN3doco/IG9C/cNB7ZH2LhQ9tY8GJhhjOVN2dmIPmJdB2L1jDGA5/B/VwWdQYP
FsUYYHGnlQelkWmTmF1JNhtJLs+TejxwThmEGLBHMpNxeRvxEeHrpj9VrCJvhhwf
m2Lrlu+Bhy/49pBArj79xwwwyIDLrzPiRkfboe+jDoC8n+7jhwShF0ECQMsSiPOM
Gs30i/0WTcYc12Bcf3VhoWHB9BRsg2NNhLV49kl9IjPMZh0CJ2i57TjyfmvhWU/K
TOhAmPtoRTGDdJtwYCOWcMInnpmAD2KFDyiWrXsdZ91D/Ofd7I0YM8w3loeA6DEN
hAVPPhdcBUY3w7GfAFuN004LGQO24aF8WkvNj6PrKhoW3nUWi4mETt35L3aSiDdJ
UrWk7qGj/T5p2A/eVCKUCgzG+2Bwb/2R0pHAg+JDqDx4zHIF+4SxYoG1VCuK5i3X
UNDs83CJlKToZifEu8q+LNNlQy2RYPSrreIUAiYGWF21ONHltjU6tdVKJ9U4TLrH
uXHRONcc3kfywRRiSgghWYDL4R0zPkalqsmpAHFxHs4yv5DnxgrrpH2++ZcGGvfs
r5rUeTIGI5JVzZjXMOWWGfFxXdD4fr9IsIgigTX38SF/ik2PJXcLXs87jlMRsLod
iWmGZ4H6cZT3RzxOMTMruNBOTsT6IaCypotU9M/6RNBVSkfRvr1/f1pHd8JZMpSo
Xe9McKYLyZGRJ2wXxojRXL4bP6z4Nwa9ytO5vxsZBQv7budm9+FvMEGEUiK9PZjX
teTMewCxB/Wj/N06pIEIg0SEZI+WFuEb1NJzeMcbPqRw5SfThvEjLRl96V49e1ep
Ae1EOCMvR9PgSxhg8a0z1J+G6Rifcnt4bPOv3dL43BtXW5nnOnqQ6daN1JSiErZN
/iMc7Od6+Sxx1TzVLIQ7Ln+6sG6uv4goeMoM/UsCx0V9l55i4XhYrBXiUFuaZgUM
wQ2rXqjR2yCFQLBMURFDfZ0W07/xXvX6rvexmDksDHSqCUMMFuVtYRrpPpPdsf9M
aYJNYyu/z62Qi6MU+iOZ1+Cb4JnTsg1AZ4C0R4jb2X+m1r5FZm5iK19S9yfALqJ4
vBt02MeSU/I/ztudFDnXx8aESUojlBHYybDwRRCgS4tA+0C569fNJTfvQMHYdhtW
uNwAc0y+FrjhOu+EYx5TtlUxhdiKXw/WW4XEAACj66YM72tHwhbCS+MwbizZdD5i
/6jmO2M5JeuA4L5HM0N62p3tmHLz3uPz1yT6XVa/VW2hSmeAes6trq03dsvNdZ+t
amn5E2NZvzGHO+uZWhVCLz3scZ5zPL8pHvtXbTw/6UhlWFFsYn7yrsoidbgNk5fE
+Uu0wpQbazEEWWT8hU/YnMOUdpymBWrpzXVCV6GYcCIKfPhVRnrx68snrWMRoeG3
nR3OZADhdoPrTNedE4ZQ06WBg2SenDGF2N8gpNQeadTy9W2dbdp8VTZQGz5zbJ19
4VP+ZzDV9DbotZ7uhYf/hl3voaXeyBkr3XyJ4bANH+7kCPsRjFAgWJmZ6XwAXid2
xXyk+NH6RbZIVG6sDwOS5vizx65EMh5uMeJNN95V1HUSdi4VvgUpje3w8ET+kEgk
1/2TURMuVxA0WtRAqYO9zTOXCIXXXC/BUOqe776fdejzEhz01qYRkWTn1ZvZsMjB
FVDzkxztEf4HkKApPQvEx0MTAUbmrsyPoXAvqwi4uks2kiG5XM4T63Z5w3Rz4YXI
+fdbB5uj0iQ9P20Isr6MszVcgdFFHebinZk3B8TvgjXKhEm3Jb9AvUDgMMDNe15g
4QfCHUCatCsalsp20qNjNLuBg5pAMv0o3jbUGGKacbqrlA4sF5yOUwYh/feXo1rg
l9ImsXrGr9+FXKY7cOSlLESzlqqRZYR2VIHlh4JObzIrVM1r8+QHWhlL7WxsXKet
b1aOGMl4VqRcoiwNRTdDLVue+mLbRSflByCTJKIAUVn3ZWs/TXbRSjVPUNgCMUNj
v4Z/uZCFmxA1NfMmoegAZJfb9kHSfuy/P/TpHn9CBqqqnbhB2HgKOdvvVhakCi02
9oaFy8DP+jnH9nOmXuz+tm/BSEbnawSg0W7Dbw8G+uUxL6ygmjdhhXkg/7cnvGbg
sztg33vBKFRP2ZeWBE/B9j5nHzgNDHCNwBswFtaQysmIYU5hUHWih+uSS1ZrMpok
D3gnRQkE3kf5zmk/anoe25PSCfjvBX+1bJqssGp/481UwQ+xTd9ETNs0GvZvMi2m
z72HIuKY2+Cyhp3xTQzKpErakHhDcDFnbydtuYzxvSGYr5ExMP/MF3uTqIwCTNWp
QN3h13TS9vs3eKzX7Bnn2NTtvHJWbfDyU4hY/tOlbYlrsTsObzYXXklEZq1YCI87
F8OAQc/kTeZ/EVTbpVFrLL2O9GfsDSimm+6cxYfLNNyNSKuxy6cqSg+JeRNXr4y3
ChxZY4IuVSx9+rvC7EsRmYNi4g7WTjGdyuOFlaLcw3J38lCVjy0uoEczgUtPOAlZ
DNul9h4lHaUV/eRCP1iH3/X49LKWLKMTmx1I9JyNru/ga76/ikdACd5Bw0sXhXKr
me/GYQs4ELyMMUHnc/UfryNvkUw90qbBTN88PKUxpXy/RHmEb6jt7GgE2IEby9Qa
FzBJH/2mbqZqHV2P3L03AC33AQiMXAx65OcrKUbu2FmYp2t6raGnbCLmOOIYYxfB
/ECSICr0Bxal/UFDEfdgvQS97eUt4kSpcGUl/fQwSLquqK7taQZ8z0kIel6UGeJk
cTTuSRPvm4mEwdB/pIaDE5vKHaVYNdvrcL3LW7ESMDtWlDx3gHejAGZqW0IAkItr
zLWl5csb8fEdmLQDEH/ROZOypmKJZLJSLxgV7DGuDpTnkEjOKXJX5pAtk1b/Y7pV
oaE4uC62v4ywPhJp+AlNmraA+EYh+0aPyhxI2EOGY+7/c5J3PvGjRfgiygi8lwcb
PGIQOv/W9jVkkZJ5pjRvjyovSpioiCLCOJYvx4wrj0/nGJ7tq8hmzW0UfQY3PInS
on/kPKGu3zq3wFzKHnANYyD9GhjKgWzy541yXcKe2/LZx3ofDBBNSBfmkoghR41Z
oOM7xrm0IvhIp5w4YQHn4cQt4HApdQT9Hvu9z0/I2tpYfFQBMa7avsx/e6DsM/Z4
rdjja47Y+UkKcK+R4tjNV+zUF+KCRc1Sw7CjXDc0jZjoUlkgkqVW9pCNt0ejUbqh
2zAAxWLNKJ2vsX98qSF55ZvPTMri1LN8kIt1yXDxotYiWjASP957Hr5qdoeV4apW
wmiMmdV16HkuNtL+mSNrAox5JYr4G8upeva6pmFbXv9c+KDyg9KgPGy8KEkcSerM
YzETGvBA5g9KPSYdgEsz6gDXdpKVqbGn/7zU7hqFiKel7He7F9UpYxrDCRzxNR3B
3kyNdwqub3JVJ8gObqUrnoTLs5X3aRv12t67VUVvx9Fp6iD+Q+8TMsnhMD6+Zfvz
dp3xFwmrJ+rD6bCpi546Owv4CfQGYL3AiMRTujDSrSffbOs4a/SHqu/F3BILx0Bf
BszbqNNJremYjypyEDIb9n5/H0na3xt3Q1dYhR85IC/NycKItnajUfHlmft3QVwT
p0MDMqeJCbqT906180aifHriuUQjxX48pkeUvtjTte4ZIcS3XkGPBRiguTDKPtW+
gmdBpEJYKD1snTIkfqx6MgouAInrfjtub+bMW5dAdNsY15Q76/l85960ugrLrmQ4
fipmYm6R/XiNHwhkkgh5oUSR5FHgPs0UVXRvjnOgxFnmxRgHQkVbJsNQDMrA+kqi
pvWrf+sfkPDjGativ0DBFPiLESBkTmF20EAe/tJExlKoQg/Cre+T2GhGVi1/HOC1
3qgVxitweO8kZDp5HqfwM4TmzDxCCQfgetEhPiJKos8FItArp6NY49Eh97S1Zwqz
UzXE5aXdngQiMdhKOFOKkFDY6j/OUL6JH6AtKvV/sukEjvmarqnofE2y71gFRooq
wTth0Xom5hSObVnOJpFPxPVoZ8ZSi1zj0TMs8tkIQtJQvLU8fdNUrYRP8L0GDy6H
2j47UB2EUWPDtUBzCIS6DHzZsCMP5o8YI2F11LbwDZgMvp9nXWD5wLrR6XgQv0Mn
ifnkS3QLSuu9RD4QV1rFCmrlRbDEcJOS1p2oRj0xspxMNLUr1wzSKgKL6cRgi+hm
/fg6+q/lBAlLKfy3jvKfP6c2ZAi5X0r9xGHagP/tos71C7RgIVnnQo7AP07YLQPi
if6nuSoYIOGL5KrDZZAxRnGGzkpMalIf1SrdcWhwqxcSKaGE28bWOUllxNK2oqkJ
uUJ6tz8j+LuDGdLt/z7pVIQiozVdbpaU09iv1/hHFVn/73nRv65SZ2rBKZ8MmDqL
0l+uWUId/Y+RiEKD5elHP7Ov+MvPqgZwty80CCfmP6jHXehtdfFuKWrgGfUmBOup
7ma/EIz3GBPe+jv/sKkBOZVXLOgTFuYTEBzIjVOPsq2vpuuuesR4+ba6JCoholvp
kU6z+M4H+MFSaVzBbX9UG86pbKTaOoF+WtDTDyCqEFd64LqNnYYu01CSDULZEHQV
LHUh9keGXHjeS6Sl6Yu62zdTAX6iuUemmh0548bpGRG131kjnMP5hUFMM+yg/+v5
ykZbaoqx3rSLXJ7U44dbXH/sxDRMsSQqxvOc0DCM80LvpV4ogvHRdZsL5kQgEY2U
wsZBcRYbBCVANs/4XlXOW6BRtK7zm9CD8ZKrP1o19q/JuSkN2Xqv91P3aC6rsnVN
alfwV+n2H8R3sB9bq/gVr7phmsA1s84uhiJ4jVRjWLU+79pl2711K8xAOdHzjdMC
yQxbnHuRJDtKniG+eHiPux7bsGim4hU9Z2xqrYkOnfXZcau9IKYNZnwO7K+BkIMu
JY9+q+kJHu1uovslAJhdiozUI6XuuWRy9bnKniBZHSPcPRXnvatp6FyOlR3v8hbE
yPmSWzpcFIgUai8PhWXgYI9nUKhr2FbObZzhZpK1ttlbh5YwP7Vpek3o39vkd1Tz
yBc545I/4DOhqoYJZe+4q2oXTLAs7I/XSSAv1v9rYdLB80wthR3PbReouNUSOWgk
35B7F4eXp244qUZIMTtnYC6jj4ZA9J1n3ZWn1SMm7+RlMFt50QVQD763ShiFqwLF
zU+qBW9tV/qN1pu2KES/lbhnFVP8lLR8xMhp9gV0gVtydwLUWULEptHjnRVi5lLn
RbGUZrgpnDm1LAs0M9Nzxb25vvKtIdo2k5Us5cEm7XYhyLqblMsMnfgc4zURimgc
mpm+lGV77PyOgA6Vb8hVfvHGbJaMTSjHOJncU/bV8GW+Yxj3GteT6LQfIuQsJ1gf
LUnEeAkTzTb/59h8/TtU/ZPtVD1S2XsaETzaMLezibhcJJOCMc0PXc5+8uH+ASm/
PHbKzfXkpILcee2uA1mNNv5y+8cZBiEM1HB+7ictcRZARMNOsgbqbgFyfrTD2+c3
R6ZMJJF1me0Fwk5bFRbKIAmGrrlkIMqeFUJ2b/KDX8GWk17cuu7b9KOZfZ8hQGkx
2hbiOJPVcE5U8OimpVmpUou7fUtpc2FVCqX9rBpB0QkK+B2ADulRwLU4SFtxjX2K
1uRsDQqz1tRmoeHIPfNd3G//PpLD+C5Yq+4ecSvnT1WkWcTzN/zV8KnfCHTX7GZp
33/qGJbpiuFGQR45poRTzJmTHLZNbnIl2C12frTXpbo588Cqxx4rpEERZBY9jF4M
p05DUZXrEAT6DoTqtVRK0tWjW/BDFiJy0BBMddkHKkqcnzBCcPvYfbXVxlDp3puh
pvP+a5yDI5Dy5XlF1fsXa2EGpk8FwZgjp6Z6z/rSXHAWCEQPyNoX4AcyV3wQRj4Y
Bwp5sKbkemMQF0NRqSqb9PJIGEcXmKCEbrd3w9y9y4hoiwjmbH0/WSnNrPv4vrVP
MmXYNCibGE+aEwMWt4yfQ9EpdW3oMGp7UpGyMbAhF8Lxhl4LRGgZrw7QNxl0X5cr
nItac2SorK7z9hWyQruDYwS9LtnVUr+1cqMHbzliPzzBFiFS2ZlxfkYuc4pUXlna
ZzIbEM3Nd9GrD5zHeErrHB+6hzm0uWxK47aUpcyszvacVnkuHR/HJ8In/pKJEJA0
7Gz21R33hkc6jqedto5rnrzJp1QGaFpx7IX5m8NECkiriorwn1cCVfjsdAJ3JCNW
sxdDgNJAPjn8iwKIqsmyQIdNdKQRTtYYw7XSkPs0ZnoHs/yCDsNI1qj4N1Q4moWg
BGozG0s9BxDCWsYye2cadZqxI6/6VaK2inKiJxNS8Rc2OyyVwrusvTJaG6NZFyi0
8wSq27KwotWTadwwNRUHiuS4WYfKgrH7Hc9b4L40vNJurqBZ/Wb6aV0Gr/EytBX7
a8ht+M4QbkpZlUQS3kYjW9HlRd2uFkiOJBkzAwcCsFDpohdutUd9bIL2M1v1ywMn
XJfc3rMErsWx+hipdrqCyhnnVvGE44zAs8h5FFO+TteoACdbnjSgT10MI/U1gfW9
TJluB7oOlORfzfykwtvipN8uxIHTB7r6CeAkW9YPekFmP2P3kBGebIvpgSjPXSjj
PypH4E/XfZ4DSler2vfGoeTrbw2nqM8M+bctJgL1S7dKqEDs0DhpPZxUmdL1uEWq
5sam9btfoAvfZtfIbAddDUMHKZNEejdWu4gqQ/IRo59pHYEkL/gJw4QRKLjQLZU2
eUorB7O/bcL03n4v1Z1gYxsNElxOUE3laon/okMFYrnt8+0Mu96cj3BAPo9aIcbb
q+oI67U5KXKNZqjWuRLudQp4pI+b68TpWAA3ESzyGN2F51GrAbo4YajyumVklm/q
4bqt7P2HgMH+k5lC17/wsxetRIcNJOlsUDDu02zBuXPDx+wfn95DixRJAnHAkCt9
xT5/GzbgYG+O9+XY1M89rkt2dv2ZdXI6jOfjk9c28AXv8LYuZ0sj8J2+ipWQzc9t
D1nPyKZm4ZVCB53hMNZGxJFAFoKaTFVe4MM52ixe98jVXwtc6XThYA2NblK8Cmka
CtY9PtfTzs9aafxKsXx6JAaePm86cD2MzGr09b1arvqcUqj33/BCG/kG1jnygf4M
cCYCl7UnLa7EvJbAU5wQHCaFED7t4gVCJq17t+FBVb4XwhtsZlsSuxWfo7mjz5Vp
znl73RNxIGXip4CpDy/wPvpCYPjOWN8An9LSkVv7/eEx8xv1CoOg2dyvryzk+c51
i6n26GQXj1KAniOp/GrCUJdibjAiHyKbnLQWcIKYABaG8w1+/0KjIKmRSZtjDejI
nNBPZsy+n01zSqEPy8vEQEwitHZiwwCvQaEROHlzesLdAPqxfAY+UInMkAi+yA+6
bW3XGrhhw/nfCzg0LRCi930V+bXDg4xCo5VO5iqZlcK/xEMiuohAQZqHXg8zLrnl
v6rAdfPZXO0BFgD/MnQfRA9lNulPnsES7LvTVQFNToSALIDcdS84zNqA6yc1tQqh
qn4oxLbaGkxxDDMK90IWpKk92kzfQXR/ZHuouhDdyrSERGBTxIPC+Pmj4OPp6dHq
7GrX+o8qT3LNm5GED5m086Ah/804JDhHL1gBByAjbtUXhm4rPhfTPOnGzewMebri
Rg5drTmfbJTUrN9+PkWm+BdTBGTCh8esS64x16MDuICweVjloznBi30GV89V3Ft6
FycDuabXYbqySyRrhcSY1NduJ9NRd80pFcJnkuq5ZI7nAgOIM8OZ6wMw+Jg8JN9u
HozQSCEgy5Q3qob1nQfSrrNUGHb338Eq/lAuTiDZ/ZVBNvEbqgwZ49CoHildiTkj
Qh931fUFCNIL3MwVdv3cK4y8Z/pPGeHOdd3Ar6r0BPWMC7WayrYgCVGxPSjjKo+X
oCRn62+QjoBeswiNQ0TjSFJ+ar9W6HE6NWL5BKcOfI4YbD1BxeoZ6WuEkxZxtTht
mq1PM4LBvY3MwoT8uLo9o+GhBqhMsf3ZbgrdS/8FEDMdgghp97PCPAnvUr2t0+Nw
a3zkCCW4ngt1QGBumka0Ln/NSWYpjARLE8D6Q31WVaAyudBn9Z/N1jGdNYOU33yN
oSK0L0wOecMiQ7ql7lwWRtWmbz/1q6fzDAuVe078FAokLlddvoUsDkPck+D8mYs3
oWoqtp8Qhb8RAkdI5DGluDxP0jFRSllWgsQgWo331aXEoNw+uJ6hr7A0H1GCJR3Z
EdgPF1h3DgdCRhr88jWIi3UGQhrWtbyft9+7xN5jzRXfvGjRD24DY/mSouhoTOfM
VYk1kuqeseKF+UaaIpEg3qHA70UpSinVKbbOCHyGeyqztjpnqNmqqbLINTimIW2G
TxGkgj6hBews7LCBPYx83dmIQvbF1ZzVYwug3gCJcTynJ5o3+uKmGNtjgB6brNFg
bUb9DCfHD74gM2qgt3Jlmi+d4y4h0gF/eeq/zhekL/Z07ByityV/S8QxbZgA98Yv
VAw21cE4ShoIQCGoHeRm6nKG8PZIh0bc/gxI04idZewiOkopTeeutHZ+9VKBhzji
He+Fv2DWVvsRgAIS0s1L9oQxguREZN4YGy1pdDRpWN7vode/j6UU0F4yTO0Cvf5S
I2DcRDfLGHFtOs9iAyq073+6rK0bni7373MTjh4i11BN6SgZBG5qUl9BirwDEWSG
mcHetv05sC+jbK85RImDN+x2cWR2N2XAjF3U6svzrFJoHkQ1a6NVnS+oHHFf+UHp
P56IXzY5miwe+8XBHeR0bCPlz3R10xSBbBcflL6Fs0ZCXjCgm53EY1E7A9yORYYx
tIMy+XSf+1MlQ4SBZHVOzHoknDwpP9S0+fSCoQ7XKLseoRKNrWiGNU+N+6nqqldz
6Nf/HUzjfgIhIMWwcinoK49fwcaw5V10wsnloLISsUDbIwwVTf32P12yIyJ02CMu
Vgz73UEkH9pc4lGtB/JwRLsfeJ9RttKUAQTf4qJs1fBhhnKyB6anu3vD9IMBKoyD
xNJqp1zoQFii9mXfCvT1vN47iZW7gwsD4sTukOHRH6NDxR3U34QlOQZzt4cz5AyB
SsrGvTWgdbWaUm1pVbKiegtDPddCd1ww3bBztZQhjHE/5i7heUt+Kn36mwP1paUH
w4NHN9KLhmwHv6GDeUOmAoJ3jhNOtlYJoevXWcj0wBFxeeWyClX6KGrT6OZXVNdq
fLnloA5t2UQdteUy9YxAEFqh7nFuqXd8QbLB+RHFO3+1FWrx2sB/zsEUMVuAgqcb
zzydnmLXTgXGA+PLUET/nVx0BPd1zzBSyG+SgX8PJyY3wGuVK4PD2jdL644rlKnZ
n69hrAajjKkt3vg3HTZCGSZVu8C6dzbFbZw+yTWzIo2k5DJGI/b7KYlbZpN39TGE
FAKAo+1Fw6SCQujD8zVySLlvSI32MNE+wKzK/mnmatXexmVukE2lkaic506jeCzD
ZGUj/4UxrZ+rJJurG57l+zKD2Auq8isjNs4pfH7K8dGmI0HzQPuXHzmbKzeYAO1N
MoWpxdH3UshgUWZHBX7HSbh2hnnKaZi5b/p4u7d06p4htsIdKKJ3tRAHKJgVUmoH
KmYOnuXqU4Hog6/U1bIciGH22Ptt2Zhwx18OT2Kf5UAIcJkiYcD4tHx3OjVoL09s
dZrbcYw0l2JZQBwsDi9qe5eSnLhrctAtVL88bFkeGHub+kKz3MR+buc5iqGv9pal
0amv7Baf6OlNlLaoe9XZIlAM4d7bxvRkCjv85qKv8l8RvNXgWCgZD+jUGuS2G1sx
7uGGCotCnSTQj4ACYaz66YgcZP0+8dqvxl3h2Lr6EbQXtMovB8yjppHJBSj3PSbw
DlpaQEvLb/gVb6GMFjuqrbfi1TwZ6ozxCAjgixEGQEumLS8lcuu1K4wgv9Bd2qXi
tjKwHa4SoEL5LSFirv21TyykXOLUYEz0337/GToA6weBag1PPcc5rHRUPW1OGa/6
CiivZLS/+JynaAijbBKdUNqMxu+qTp6PWxB4RgONye2LzacA5nbY0St6tEJ4h3r9
2IeGZmxh9Wd1gRthg5c9RO9L/IG7+Vt+LeM+lFCaEcCrZgHMIcjDHp0BBn6iQuJE
TuhD47joMmn7kzFDfqoYciSpyThsulEW8+FeD9kC8R0qYzw8kR94DhMdlQqn1W2i
c4P2/5T1HXEPQ2BGx/9NlI7625SGROdOQQ4Xy1AV5zjjjPy4nmvKO6oncDEuc8VB
Qjk/a7AeYzj38xVdgK80aw3Lmb9dD97++EHIedMxX7z/tVfQ80wIWyaP4NJ2bhxG
OFXZPL8YbvtIvrv5FBOyldY5Jqcbt/S5CDpkKeYkfETjrfZZfCvHd3debQkOnRpL
CawP3a4SILAoZ9JrSVnHuqHYSKQtfqJxBqcg0WyPrcRgTgEaZBm/Ysa4QhcQO3KP
2hWiH0bLJqEvJZZO3C9VnN5frOdr2AEavVKIB1Xf5j4hx5+EEqd5xL6MImNWZGrc
jH0bcyOaT2qbxJHrqlDPE7pk85OgVrKsNrSGgCBAKkgGRXEhL6IKAIgXqnu96sGv
E539LsPeEPsh1E87AnMeqHqzfX5BquEvTROoBStT9S4gge7mIY/FC1luPTUaUcFz
QslCz5yUjJBYKKTi3dZHidXeb/HP6rcP0azXOyj4iyPrDPfVIfFwPHdOfx6kamZZ
UnQh7NzK6TJwKzzIzI7KwbaGKNislonWkZFkenGqfOp+w3kHH0djDpd1pT1CVWlg
7LQxBAiVK5blQO69uzavDq9uSj4gl6qHoTnkVFIHDLefTwF7SRvk98lXzy/dTTNI
f7ZF2nc7moi7ztZeMbQnC8q5i63rS/3NgF2a3itKdfk+msJsdxaJc/1WMIsDb9S0
4ipGRdZmNcCbbGQK6E7LNdii8PdBBaBlecqn3cBCVB6XQH0Z5L6V6aJxCYLSzLhP
SWtnhU4vor1b3XccTPvDNMxBhsUbzpRym6x18NzjL3390VzJanAb/W/fKGmD6Bd7
+tJBmCQp/Lo2LaREn5C5NwANK7CYyq0iyCCw0qMmMiCiBLP4LDa3YIhM53HnIL88
IgVr5N7YsuchO5q0x1tdBY4Dydu3DD4H6SpBvL7YxEXnZOeuA5aq3bW5Tt+kCsM5
Z2cdEcc2aJCrFJCIRXoNwvKL8aZL/Oxl7DonTmd60uemmjLMNtcwJtrmNsRHGVnv
42htO/Lh+Sg/fXUvEgLrMqRSLDLsteXLLuFXBNE85TL4NQbib1zU928S0cP6ZAl1
nDH43Tt1YFKwWX5RXdaMX9Ugphkph/0h5U963qhG3xPdK5k94CeZ7dGgzLBxtjG4
nMqVY4yg6kUanUUoqRWcqIL1gU16Fk+3iYimbGngQv05FL5JC3GKuF6+O7aTJ7Hm
mKJVopCe8UnmZvbpi8mjoyr4EXhbm7EG52/m/5/APuAQQ61NPvADS1+ej7cbBx+h
coYrXDWL60sSCidprAXfJj2Qp7JbDLsjY8FJeYtOKdVMDAPLLNokFdLzJeSOmoul
0dOgSC8bKorwPxVf9LUuIUccgMXh5z3wEg6NdUQpXtfvCPYyiOKSyuCf3GZKPQSO
fC8OFAC1JXL+b82b6SZ/bvavoNnpN9UKDMuytAEMty1SBJ1qi4N8IZcUO7IhzSfD
WC1d+ksKDw8WLN7SN2Usquc17FZ19+qbdVsg9ZMNlusTqgcj80mnGgvHIPNBLnKN
7lmALFwkbh9BvF6mvWNlfROP8qJwX8R17vLzhpFi0AS+qHERc1yZKYPgupsdJtah
1yXNkETllXxWYsRQpzaaKNR2trY6xlVoXv5Jw3oHQihKcK53u0y+uBbkcfYrxV+E
E2zASCHnczuT02ilHnxfk+L4VUj2oVeWz69laCu62uGZ4PveFTu1FmDSU7ZYZ6d8
RVpoNaf1ukxkBlHZ8T1hkM45eLl1nUj3vvWq8M5Z4lEPX8wxLazpZUL8W2svQhEf
POM+6aiOoTHDknWezfv6VjNBremxbSnpzFjRo/9WVP84b3/t9hwwCWGTCE2GZxIC
GDAP9bJxan0lhZmGkl5CVo5kvOI616Ayz2tXXFfyI7cPXJq023f3SMaxT7o5UKIQ
R47nyuouvIRnFD7AaV9DhpeQCjuw4RpRt2OXFBMrYZDqolOx43xpQJcZp/TV5F2P
e55JmL3RaZ1YxJxOIiopJAsMc5BVM5E45cLSNi0E5nb/OX+pEVu+eEr6gM5CetNc
wTRz00y/A7AiNPGkKzjzZUITYkG+tq4R/RxRp5Dqfpuwko2nuR30+I8dGYTxoLhq
KDinfAukvysphKRlF4zj5+PBoNL5ptgsqAtVaYaX3lV/EgIiwkCLVJ0CgOp9S+x8
QS0krQKfeElsxTs4EdBIbhnNyCUWWMoiLvwRHTz45EvH6JGJ1vrvBqy5fr6praUW
Y0dFQavy9M2ouQiMzJUOEQsAPa6WEA31NvTGTonz4+yzOOZKu2Z61lNWwOfPHky2
mVAlq8iXTL0phQp49sSF4Pd7qaPxTjk61vZpFNDLYBPv8JfjjbmgI4Apf6OvlvYz
vdh8k0KIIwasaSJEqBHzb5rGJvRozIN18BwzDHUFmtJefTasxhw6+sLxOqxvW+A+
w59r7QB8d7BeoBKNrCKisI55YpcPWEbp9xwfMwHOC02krkAp1y4J8Oy8JQ6xrxyQ
j/eoJTmNhyP/CkylVMtCRp/91DyrMLwhh4kAFA7ISHuXSTylunFqBnn/4x9hVZcK
7I4dMqtSniDHhmuTiBnraV42sXiYVlRo/OzG4iKJaUr2vJhtwUQ7sn8SCGhTM+34
X00b/iUukuwkwC3mty9Tig9475EvqNtTQeEs30mhyR60XZnoeaaaNBdDqRdlWYEf
/hgsjvmHKRtvQqGLzyN/Ao9vrycQVJvnmmz3iwl00cSv+paIBDaCWfTukbEOHANC
amAEeE3J6mhrmuKt/MH1rQqUuKG9gJ7nBh7bkIUTJVElvnODjShBM6xfvFB+msJA
lZmOc3EITrznrvk8n1yqcFZ/uCufIwcbMZeYZCGURuz9RSwhU+Wuofn2Z9EGG480
NEzT0JBb2XU1r4uQG6PuebyKZFpRp1ZXpKkjO/epM51ZsxUmIVoiIxqYVff0kzZY
5Fri6VhLx1/2kZ429v36ke8S+H1Y4Yyw5GluXsFHEB3l11+BAu4RAnZpbeh1bg1p
2fCho+YdDxlCMXUZ2Asccih0GkFI9dpPF1A2hTPXBRD9iR5h7h+wkDvpmKlgIwQS
R9h1iZEwK/Kj6JcTx7owW2/G/6bbDvs5F9HTJnlZqOGUkCVkhqt8Is8sWWPNAK8X
TMsRgR0MyhSUBTUVaCms/olYlxDAVj7Bv/RMs9QL0bve4VtmeiJrU3ECRnXotQXQ
9//ULYiMaaVPgmHn8BGYKtwakGsU+wEullDnZi9CqVuVMGxM2TIVvV2b/zU2T3q6
yKCWMMGzfKdTG6qE0vEJkQ6hYWIuF/V2m6bYLs2vhi5gTLQLBstO1VcROv+oVuMY
Cz3UuV0KFRob21eJi9p7n8oOdBw849gpYRKfz7Fsw15P9d6g6AQKBP3Fib2Q/kOt
rc72jzinoHJ62KArAPC7m/0xqQJvdO9von4O6xgaYMj4GlSqBnUccRJp642PhiwL
hRy7qy0h4VDtgwU6ZQbk/YRVe7UWd1juIlG4GEofmf6RJmcpkjIxni4g/Kjv9PB2
JAQgiikbREfEvtH7J1/GylrYMGSrL/Q3GUXKBHac3M6hkhsOxFB1iK2RbsJ0FM+D
+JGfZhFMr+rbmT1HoYmv5jb4O0XruDbckTqyddRqcQsFrqEWg5z30TfJUaNtC0oq
uwdigQOTWd/VRf46G3MurpSknao6dfBWRtcji7cMvBZj1UfZaz3QxCDtUqmXWsSy
hqXdY3bgmaowLZK86gN/mHWvxspz/HGj5dnBCIIOH07fo//76fsZtI6d/STwPJWx
5NRIT8Aafor86kFkL5zewrHJVJRuZxou22uAg3nZhHr/7ZmsOIEVsrGVJXtyekIP
uP879fvNfMjL0c2S/lniEh+cCo9AH61PDp0gyScKnbUYynq9xZ36waMPWfcya+kr
3DGOTcF3/EGdV/UAsSUgRpa4mYiqxc8fDdZdlaXQhk/7W+PgMyd0+K5OYQE1/wcR
LijEqBnME6W+HRsb1cQ2W20Z/Lio+VJUh2nUVEThoWthL3G1ZdWdCPKgzH7fw6td
bKz6/kcq9mAptMuHVTVmHRzLK4pNp2HAfKraygalwdyCU6E/aJosJkL+1XiE4LEt
YZLj119hcQbomDKfHN0TQSzoru4Gqtq7aMgmTKgTxP9QyANRMoU+C6VF8IYWixho
bUF3rgjcIQDG+M3tkXCg31dWEbY5i5TQy7hi6Ic81VKX+0AJoxctIYyfyi740HRA
hZouuVnbUpMgAFwsCnN7Q8vZajvHTj/RB2BXVRoqaWMmxwJK2j7gm38g9SCoQmuf
DXf7TPktWQZTDESw4t1li2lODlraOSqqPtp+C6g2vk2cILD+1fTyM6XAccUB298T
i23+lCX+QH5MgQDy9Bk/Wn19c5vLfIPV3ZaT1F/TFDfspAqXtx6OqAoD+xaCQg2o
SGpdD9yLa6/BRPj1vxCY/AcQHCY941PnceFxd0u8iiE1pQnnubQAgezgzOs9Mxqj
/PA91H2o9eSGm+fy42yehgGebF/qvV5R22rRzBTX9TW2lE6rwnk0gj7hANpZ0hsO
nT+mRsObk4qiNofweR1qu/BW80Bk+bqJKodud9UJr23587Q4GTXloAOb+dl+zsBr
Wuyu+Wa1wqRhwV6hvFWjYf4Zmfcm1lxnZ5VnvOy3XJ/c3Abm25v1Mw9l5djz2G1l
a9IcHJV3IoshyQj9qR9Pmiz1fOL0DCahSAVg0LC3aj/obhNBmHJcHnPRdSCVAwLH
VPEuogyb3gGcpwv5z4qIdGGEpIcW0vXHlOfxR8IPDjT4aOaMuv/iWpYxpGSSRsgl
vpHsFQZhzKCUDI6hewYMlbdEq68Krx7Z1o7kSCud6dEUfdfpoXvl9GDlDwIfHwcK
3lLYscB5HfEFkuNoU7V14OC1gbQ4C7ENR9eayQc2ezVKcsAmdYcNwcs7siQ6gOw5
E19MFyqDTXwzJGup8s60lfGOF0P9Yu1UwWnOTjVmOoyYlZWigpZjKQ83KYX17n72
9BBvZ/TNQeAtqmN+IeElW5NgATJC3NCbzNqHvqM5hq3mMo+/la9IMxLCC/lcClSV
zi2pqlOTmnDGZ9dlQboad6Zhy92uLv9HMPhI8yHHTmHj8Uuie2QVAJRWKNqgOfvn
AHjlvc8s3JxzNnp9OLFQJQ6ddlLGW7fEhnVkGdiLal1Tqf6OYWBEcmtlbYaHOmxF
8rpqooRJImBpNFdeEFIB84T0FfoP782A3HXXrRxAszh4MVXARxiKhGfZQjx+P+7J
UWegozjDlr4fyVHNEesuNxcSWTwozzZsVTmS5qmsS04dvI2RgzvNwh2WEOlpFPsf
t6pqTwJ4lGHMMbJq1Q6/DCbMHQWh+IPK+PBFYU3CcjXPlUTF1doLRZFe3CDmmj4s
Pbhcl1YuWyi7Aqtj7OPYSCtxzS29ZP4wqncipkjoyH4+v+qhmvsiiFfUg3m9dSuI
asAxj4fsITedIkBozmY+POSG4Gyc9JJaWn1ql0uz4c5+koOJ/aeymQ0rXMFnWc1H
m3OdVNNq4wX7YvHC7P7HMzRCdKn2K/dkyhdKFA1qPBcY0IAzzALyMTYzmRtaEZjY
pF5lt0LmdjCvQ9pe5IHxC1DcqFYcFsOyxg/wFgnUAR8dCChnnEUGPVVe85jqvPcQ
X0GTkAROxxps0klcG0aZARg7DnnMrIKVs43M/cbiqkj0/8rh+96fnEF9TUrxqf0I
Rm/tZ11MEnIMlJmz32tbKVAXNhMfEaK8u8sKjMurigZtYSTxYHw617FnAjDE1YK/
l3VtahoOG0D3dPm9do7uvC9Y/mmhr0F1jgspJDuBEM416zZM8HunvavDkhS1r9Dv
VY9jUMVOr/fqwqwK+DECkDnuIM/2XN5UZkobkOct8C0SppqvvLwwX2NOaAz7UJ37
kqlxcBpBdH+KkUcc9ZSn2rTDTMOo2+JOMYCA/wQ9HVlG2col8WhPofDWLQMxExsn
sckBNblEQaor2LS7UIBAXMD+Jlh3mK1U/h5/p/tHSpBFTzXdIuXhJ0xctD54m0vL
W0qlyU7hPMZsQo1ZOz1SKNtsUzx13KWYdjAaEck5ASw6xAt7xhHS6QlqaMJfkfjJ
ut6J3PGWRBogqdIWHmvev+8NXgPoxbgtJMyr/0GxJqDWKsZB51pX/TOh8XMNzNQH
qRywz5B2zVuYYNFOMrFsZrvaYDmRBgAG34k3dYg5AjUpCG3XO6sbf5VBbwHeC5oT
aFCPGRtw82alLXIRLz+xdTDCJeQXZ6wXV7Ks05m+fWQXKAZD+27lOwYv6kfbQMML
oACjlVd246aiq5hUtlsCK/oUu3FLMHlGhOs64zHdUKlSct2U0zS4pbZ6pvFr3TqX
7qDjArT/Snl7q/MZ2Ko52v8MeRF6jCuF+iHSjVc+LR+sMOxns2UE+iPC05H349S/
YuOvfWmKR8LI+4EoCSBERWcnA4vuw+1cZUXNgvhP0O1GTcAwukKjnKBtl/qRUSnr
34rf6YypCzmHJyvXK6EO7gzyvuqulpevRSkhOCea4USttuIxF6wihdEunfjtM8wD
dU3YDsZoUe1HXkqVvJ4je3xUeaWRzNpuFK4Z2WM7N4jtGT+v/3T7zOaPpxMhzxJD
vt7X2SS+zHHficd8btIbFnbGbBNO2T0gYr+U7PiK6RwJg9g+t5jNEi6xNmeGbue9
SPqK4lwXPxh6e5BpYgKZrz+1wmWdF2e2mGQ8CMdAbHoNphaPKfkFp1OhJ9TiEt+r
dMqNy/F5/sgoHSegmqPxTaODZZ2/DzLJGz+zlr77H+ibIs32sJLMixakY9F71nmm
qUTO2vEe60SDdaRQl82W3TAwKNosYtjsfskKGtKpV2Mb+YHga8NuDTdVn3NVfKrH
olr9H4op6u1E35xgOkbnCre60+d1wByxwvgIWD5lk1U/5feZ/dkKe7IiQjv4LqPb
xcmk3j+Z9Igl5GzAJEWI9dFLvIXnKohPX/griq3ni4s3lAXvk3SyfuA2MKZTA61h
SgEkSzx5o3p81Bf3rbUl2V7PN+6+6Drs/tZ8Q47HN/l/OEZ19yb3hN2w3yTQ8MHt
5glMBpPCJSg0+pyEi6moLfe9UuQsy/OfAlJDU0syWMdC9h1LbkI7i//v2Bb4QDK+
s4cs85lg3MyFQ+fYR0dngaa/c9/dJbSmzJAb1I78YYx2pjlwwShN3jkltWGul+uR
MIz6tROXgSWRuB+xRjPEdtZwt0DP42AJMlxqZQjiBd+RWz9AGE83bd7FrIqz416b
nGCodUo56T+Xo2EEyqYxuxxWw9lU6rUS6QvUhYZ/3oCITB0IPSW2hymAr349VUT8
oKfWbxNHjx8cIYVF8EnBVrd9trZmKaElA3R5VXuL8/Owa8ajKGjfUS8dnQTl1b7m
ad3B2cqBLpUVfN+SkL5TtUIZLHT7HkpMsdz0xhpWn9H4PydwWFYI8grghX1H7Xiq
KYSiz50Yl79I02w9MJx8/UXI5103Nd0ahK9W2xvTnX+pVp0ZxcD37bTAkqTFnQ5y
cymBhpq3Mq6LKl46jYYnGWg9ArDBE4V1/Q35j17D1wZt7U7wTUgxxWR/Kio1e+eO
OC6MMyyX3D3gSqsaCOHIH9q7zkkcTi9unp4WLGPRtnRlLzB7ithyfSlppdnDUMD9
7+Yc//C9qDQNJen/4EQphJwj6CgtC03Sj6n9HkEMcUsCWwRfT9Z8xojs5eY/NFUX
NEEhIPHvhDPDZOe76IQNf+3ikfx/w4J6kOpXJOiUWZKy75xVGj0hbaD5+WBu2ziy
xKR79dqlXt42wFnpZmyaioulLCkHN6c7gzE0dItrkwWQ/82VylbvaaUkg/6fhYs/
25GqY47x61EMpu+pS0+NbBxJWQ/7Qd7gNVu4E5fSG6QsxFctUuco7d98UR+nsykF
YJgr9ClAhCdwPEi/tE4sEpMUpnuGh0DXaRj2UfzzImuuXd93mafzXRANr+9uhcLB
8GxrhcSAPFJhA7nGVEoCpt4n+BHeEbShK9Xtu98A75mVooriEAhfDpEZQpjr21me
k3RkyU1aZlQnKJTRZZ+Ff2R+kS0dWxf+Zo2ZRXOuS4K8TQhEfBBV0E0J+rPhT2vp
XfcNuLvB4f8sa1ZOxUh8nw8e1j5HzWaOnaJs3TW9qYCvV7W9VhfZQqMVD20ZG+/k
HgDSJw/XzGnIzolNvencSbHEIY656L+DJv2UYRLfNAnMzvLQ0+Krn9R14fEDQB+a
s2mDlT5VmY4HkD6f7k1D67Z5dz/do7HZgh19kLFUj2Vdp2rkSTv0y0pYYCwE0mug
3Uo67w8/60vjzYyx1xWHECTf38DUyshqrwi2Iett0mlySRICUnNFK91tyjICg2yX
Jf1b4JV9/eQ9l/Erzsxs74YYLB0V148bqg3m2PuF20JyV4WZPNzjS63qRx5l0raS
NaVTB2bAbdzv+HNM14PdPjXsXledeCEDP2kmvkToeh2br3IsXqc+hpxhBWQhYTpo
eQeupd7z16fZi+JENuBQto00sFClxIjRfZZLcirZTvMqbQrnmpmujF/DJft4/BeV
56UObY8ZJjqkMbS6VvebBS3iNUFl9RRN5wOqO3XXraGKZcndiguOrw80lbJQTQgR
XqdSjJGNH7VwrvDx+h+mlEWrhq6JABzDxhUBSeW6FU03Lh/TNzH9O4t4okopjk9f
4Wpybi8jmH7+Vr5LJrYoeudLH46RnHGY7VPkPNddZi2Ap+ti809pScECTJuFmE5j
5HmzubXE9YKV7czX2Bi5bPaC7M/kRlzsgRJfQW5jsiLAOEh5ba06HEPrFmSg9bjH
uEvM1cjeciA5W6M5X7j3nnWKRcImXT2EOI63VSnDa+zSBbwpmychAsQtpxWTdKs0
A5MW2nlt0IIsjNb361f1Sp5bj6FplB6UDobGa4JxtJFz9Zzd0RQuDk5aBZ81EJ3Q
4tX8wQQL7SMv/KEr8BQYqK6N4k6JwEdNuOCBHHVy2LjdsFLZOyU8Zs97DYzdMljR
desYVCbGJ6Ni1EGNJlCwX3YTbamchwrqNCZxBFUTKKogp9p1Y/i96Ps9y0p74268
TZdoM5SdCtmtlADXssYHX0POexbgBvHWbqMlknI+beRGLgzNrNpFdbVBzRzTSWCo
uVcnUFWUSJtyX5wTwQA4wqNntaaP04Dmei4AXBascXHbW1fo093YenqHlqeUL2Mt
V+AAVSwUtaRsxGOVm0wYKevfZinBvPnKwhGkHgauKvsOXOYuNF/Xmq0dKonyy5yc
42MmSORYRB+0tz+6Aq9cKWzKNbxofo57l5R91tNg2s7R7bNKU5CY+XGHKSangPeo
V/OfJqmydjCBvA8jqzWigV8cZi61cYM8Z89L+fxy6JG9aNXpRHoLHH5k2FXmWRQ4
LWIwfU09yhDTkwhvao5GLTPxlSt4r7DCMZkSHRGPLLdRIWYzyBI4tbaPyNhprnmu
QETFl8/xIppxksRB8F1bbJ01idiobx3FxneIvieG1wBKkOGZCapOw9CmwAqsVdyA
d+Otxrqq7SdE/y9U2FKt6L/K9PmiiifDlHWnI9dYci0BDnTxrMPFzYzcrE6osYu2
+mJHAm8f9PKK+v/jSYCtvn6yyPHOupaaF5XoQUrzM+Wy9iEQLFYLFS7Q2IB6j/5D
ENmJjsof5TLKJkdVZAInDZvNjrS+2hVJNap1WH9vfa5JjUCyE560x2X67D+Xe0Q0
lPRzUGaFRW0ZADU+xJ1vdeVpz+ydRFNDwiEVUrHClOxzf4P/bP2SSbtEP4Fq6jUU
hMnzINwkLhyE5AhQiofMHbKwL0iQE6sHd3potiKHwAOHB992YDAPKs2H1B0Kheql
lOQql5TemGpRp1VKTMlZvclk1RQIUV8qjEO6sH7/j4RFlsGgQ1GuMPfNaYnGhVSj
+lRUJCFCbq2fVY39tXhtJWEVMX6QiWrzZ9M7vyJwPctC3LJhLcDGOizuUCtOLCPw
R5J0tyRsBJzt34K3noRj7td1CIK1qVJypGnbIEydGCwfSMi4KlatApPro6QSWz6T
AKP3hgg2T+Nr1+HbDYEVNTqlMAkrbdfgfk5mVok7l3vPI/2fRSBw8/wbuCXesyWd
HJeiMZzwR/AkKpzRXpluKpLvbr1aQs38ojbmffzD9L/7uWF0JC3FCjmXv3XWh8Ko
Y6ZsBWSN8MYOFwuvGtV3gXFLGlABEt9fKD37o3VwNLyDlMD53DVlyyk8GNH6idSJ
VWaS3RG2/tbJ3ka7YTe+7MqyGbdF0LDSTZ1hzUeg6LIqC8osqSDwX7fvK5NY8bQS
+49dEu2ocPTf59KJKdt8X9COoxIqqfgOSAtLxVEWBjdfjgkbJYtKWs2BG846JS0g
rOk8nyVU5CqRes/qKk2ABkSOwKklDBGgKp36OezWsNO0hBFi567u+W1ZZL8Z4g1e
BzoltmjZ1Ho76uSGvlRcAvNV420YOj4YQWB60kbr5TOnbAakK9iOAXGDMSZ6/kvX
lI6FeyUIQxjJct2nwxV4YSgRSlLpI0BiIsi1nb0LwHgjdMi6+EuqdevVwpI+uJEz
xNNRNS2dnB1vS5Llc4W8dmJHgallV+pY+VLgTp7ouDJ5XIPBi02BVRFvj+YuDxUR
fe6ee1l6D3Fu4hCTQvb0vXLZOGgH3z70i3GCkVLnSoC4A1rjQr2CeEu9GM/zod2X
OyO4IZTNdRhUyEkxua1MFb0etKACZrxRq50DnIQWJZjIUmK3RUyLLQrnEyiYfmSZ
gq4BGyliVqHz//owjhfrRUoSgNnexJiOY/a+VgtskTgmnk8B4q7fuRuLTCuMkJRy
8pO7fIm8+skUke7Ei3jxZBtYJoJ4X2tl/erf94tomatggnL02VJZ6+Yd/Cyg81Bb
TJI8xSFNuhQ1IBqGnQlxmSKeeRR4ZbdqwJ+OnA2XbaT1QATndoRvrOcLgoM28CA9
uqfku//Yfdvif+OpEwgb5EDnOlBPOa+MP8NVTR9Yf7yM1xFFnuVZCJUI2tNY9QWb
6yrmaVuqoE5zGPyIRxKIANOJrVSrteqeFV06Mvt91aphwNZz7I0K8t4w+xOPEPHY
wO9B0bZMAuEB0V2YDrAZgXq7ZLnYWT572GHIPQINeXMDeYAujJkaQ8RuyQjT9AnJ
dMmFa9YrPbyF5KA6FHQZbIaO7TaJtLFLIvkBXPmmit8AATreOm6qqF/inRNtmeI2
AjXJbm2JG82Gl6jTTphw0eAP+u2PSODWn8fNd/rvIGdCvaa9quO8hu+6dgOUcpUo
97ROHtLqS+hw6qfFwb7rakoMLIw4sR9NdQUaBwLNgzD3goN4L0jqpMye0QaMMrnI
F2WftKmybH2tOQdVgAdjwiiJ5MZzqlUW7VDu2yN7P7Qz/3xoEyiL62vhaQsjMmyX
bIWIgsaxFLZviDJY4CjIHfMNXHp+KLNk6i0Z13wcHokRH7gQsZkeVlqV/EkpB7YK
UCWwIhSE4QlajvS0O5eyOVy8lPvGjpCE/A/l7iGu30HMKA+bL4ksJkYt0MtAwTBd
2RfzxZpV/ZRwIdxJuCrEWf5NE2h65rqtljsydY/83wbUvAddMMc43NgeSnbMhSU9
koE65CF/p9fVrUIN3cxdIpTgiDP0JPkgusa1TC/QZJxCHJIu6AoLlut4eHhiFZFW
Vr+7vR2ygofXfg7Y6jAHS+dry5svvqPM3NZPvBCc7vbs3SkjorStMPStgAg5pTcB
y2C5wzfs1e4drYpACu8vQksv7jls/2hAvtr6Jcr4kZWMOrrQxX6OvoYNCsPYl3ch
TUINXVT4M59l6kZSys3h11pgmmrPnJ2jTRjptk88L504tyRHM2cD+KYJ+xiBXIQv
1XvVjduOx33FGNYZCJ9bBvURMJ7cyh6vRsyWDElDzWl/usBedGr2NbiOVGdmzDiV
ZbtP6wFg54z9jkVeh8vDyoEXAUIEPC12QHdO/vyYAupwvNmdpvUtW5kcrWyCb3gv
IGq6RhcUhX9Si4PGgNBWx5iaF/D5m8LepTUM+5ELJNyOmkaEjawENNVQyRflqtuQ
lCxOmVJWDWAwj9k5pSI/qsRQbELYBQl4pFQpgUVhzLDgDcUyGt7h4RBwdXr+WThj
kWant56WCHDw1HOHc2+UMTxaWSy6BcOmc+D78lLcdwuJZulQz5ILe+ghmURUTmO5
2RIph6e8+2dqD+x8owVk9lga8bs7EVhDs0JUpxi5x6ErGCfoO5vkG8z+Lhu4nnle
82HEmUeYH5/zAbN6HsdbZc5qgl/kCwHVjNT4WIM+68qdw6Olp38xioImbSDb/cTq
cjaKpgvxf+DARILlJo4+4Y9MMzEYEyZexf3O26E3aqbFch8BUW3+tHsW+Vg3Lh+F
5ch9XP40Z9onFRgwzzdh+fAZHPz/Bm+tcP/phZd8fu2kEs/qzwe1SiqgxE1PYLL3
Vf8ABSqG0OvJ6rNHVkGEECfu6rxwZFRaRdloi9Bf9i/rkU6WKsjB8X4ydOUJURm2
0iBfXT+BSH9yIOp+3koiArjNuVBzoW8pfDRDH6O7uwDaBJlt7NLUic3tgWBIQy37
ow8bOzLjje0L/pTmv8PTtuvhVgeqs2dwd2ea19KfrQLmbsPbFu0enwAbjK6Gac4a
0Bt2BsmiHal7JNhOfCXzshoOcBTbgaioB1Fh+RhyqEtX/J3VWAHwBiskLEPy7upJ
Mwm9rXz26u5O6/iwkV9JAC6c1qv03aCEOqiCij6BFwPznGPcY2Zkm7OVAl0Izv6x
y35Y0oDWFYgzTe/isee/Joiv+PGgifrRHxk3wmFRkZFSuYXPGcHXmAZrnx2s76JY
Ipk/e1pQDBRC+ExnIJ3YmTXjed4aFjtRYc39vFSm9PoD3/Tjy7a0SXOmwg989kKr
pnaoAKYcJuA9Mo+np5ipjFloPTKYGOJdB9QjCEGAFHptse/uKvcb7Y7xKzAI65ly
Bm9bKHs+xnZqOVhPZiCsqrCDl9kPzhhFzLL9pwsg4kgKE7g8cx307V24LgL5QGo4
WcC/b0sP47wpAAsSbKhtVUqCV70XpDDFBvsUGA+am7CP1r6t5K5BjSScaXw1N64G
7IN/YjkIqX0iiy1F67Yq+roXKMmQ3TfefqyCdrKyj6nbND4JcgXea2ddH8v0uEvq
g0pJMpQUHUuRPSlXbVqJmvEV1etIyd0Tsc4btfbUPUFl+wbssCi2y95NvcZGSVg/
3QMbI/PQQ+yODTQfw3GZkINlVtyWuBlkyvUNCS2WBE8bRtWPvWZcLLQ/gpWeierF
L+73PcIZ+ns4FQ2zjE82vSg5gpGFrzRH8l+n2H8Arbw1Zmc6v771AmpFH4l+BF5x
DTeSNdruWIdNJRcg3Xxw62KL9eWWjjYFON3KqY4qf3uy0Ir6WmfHbac9WIzDNnHL
tio+Vee/UnLx9Z4l5sf/gsZ18wwKWlL/KbnZm0BylKlIf7+PJhx2+46zIaym82bB
oL89nYCIohWgLk8714JHwludIRFp/hJAhmh+VDu2Tjpjiu1hy8MQxsmcUF3FjH3R
wJ5XO8boud+LlkeuTj4FdZEa1y8yBWPLaukj2Uit2b3NFl+mluVCSo1ZHSW/ud1f
3fdsIxuf4EQyEUB8cWtau59W5ELum2EWkGVfvzcuF7Y4nEc6EN6+SPVb/BoruQS5
v25QaykNWXHjpUuNZjk9GXp5i+i6igMY8ETbHXwiGVRidkcWwLYTz46KDjBDLMGC
PaOSuDTCj2+LZXI1Hx0uJbPFmf6H2WyqQGydTUUvyvxnYab3JcxgV02NCmP/lPuY
5P0aAeGQAbDXkgnmYdLHfhkElJ3Lyi7DOcS17MBvAtUIrY7IxbbWJyqUpCX73z9k
7kmqmEeGFYEH3lVyMTfnHasM72IhmNbM8ZjRsc26YBqz3i52qVZqqU9x/HfGwHMY
7ixBV0X0GYYFGzonMp/eHG5r4RX/6Lrc2X1tNtLOzuirXq+LhQOOpACwXRa9hyS1
icplw/0kL5swDYxs3syzt8/VoygC5wWrw9G2U0jqfL/cl9Pr7XJthsBIEmJpuf9A
Nujcdnqzg7QeYhyMZJfPxeEf54q2QTLD6f1+ajwgPFK+Uk4/C9JWqAldGN5F1ear
oJGvm4NrJf8TUiFgBQovd4/PCzGT6abdp72zKul4y2Ns0kwOrc7B5ks1EElOhBB6
jQBvpp40vdZZc/ByRe5LpdcMzd/fnG2DgxjGr2XvQCTpSyLaciKPW9keKHP9Ih6U
EBDNydRYCrAqQTd/HrOPXoGrgAuT5tcJie7o4nsjquWPaUOcxF37g7nLZN1n/rCG
hXP/mwFNBcvOdjyR7L4Zh5YApwztypnre1xw3e/P8A/Hy2ypSYSOUhxHsX9u5jzw
BJWMYTnfI/txXgaVCjRgcf+l9g18DniizM989H8g8aT32NzIueKK6eXpsC3Yldrd
Q0O1Zb75OoKGrEx+1qDPI4xXSSGERNwhOF1Y4mlHfzLg7j5ec/7Mk6cQPCVMOcQx
HDcrQm0tvFDrTyxrwdyB7GRUWhnFCYPHquxLyxeqihPB8KBPMazrMwbqjdP5Upn9
rmQ+adQBb/QQ+n6+cEbyTNvd8j+IPj5lYqaH+levcd6xkElz94923hpxURNM1Q/g
sdQ+93Vio0CniDZFe9UwGCOBbyDyjgJAw7QxUdWzQGUhspvWNLhvxEm+JIZDpMSn
HDjtQc6yusfuLgbpVAb7FHOJL3o+xbdO6ryOYLGRszymKuxHi+uMJJJUGWZGe25b
y0kYq1Mqn9V8+2RpLFvCXO0W7s8BHlBNrd4+YHMYEPnqy9Ou8cnNbVFBbW9x27+g
yQ6TdaDWMBN+uWvYKuFaprtoroMUFRfFJLsDZrcWIGlIeY8bUT5W0ky57ksG/SNj
qdqsS4SdmmSCiqZVIuAbhEixRtif7cH2ZaR9g23ZgatzyYDH8/fZij60mkAWc26M
iQfMd2SO4OTzlCj1QTyfyVsI/9TR7fu99oKEU+HhrCWMFen19r7ircqavTtRN6oV
64nKt21+iixMWoVnUDcugaWylz6kiee1psEPlYXP78gOKk4rb07dOBpiKCKfc1t3
sumZb7xXpdUpflzcXc8CWjEwWCSAiTzRZmOaQaDkUjdt+ARk9N/uLlK7Ijb4dVnw
f373AjMHzKQp/UszoyA9gjoyCuPaBKWt4gOOqvvjef4Iz8JRHoAaSoBZXrjka2Ah
FW2QTyirjZcdlmCA441b2hsW6dJq9xssOuiThrr3FzSdDdiq9y5e4NO4gSKlmftQ
ZQlUdoeFqXf5Tq9GDYwls49GOEUSJQfjWiLwuX+TwHnKbPax+ZqvDCEZIs0btZ3a
6IS6bX3lsJ9KfEu66f4IWYJ1Xsz3/c1s9SbFs6/9xv/9DvCFPB+PpgAuMFbYz7b/
UVFtthZCtF1Dm3Mw3892pol2fIDB23/HJE63xzNXP3eD1PyXYrDMW+g6kYbErc4F
rJOs5nlgPnRSqBe4HJDbyWC/BqmEZ55q6ob0+YkntMbflVdIm0rlaxih3RNh/Fqr
o09XOQs2c9TNdpVEE48ucGzbxcZEYps5TNx5hnP9qLBJlUTe7NPM0N1FkrpKvOSS
ijmSvVsq+K7zKfrYRhjBIGIbm87wVSe6W0VZWwKiWntq8vzHXjX7ApRjM2ibsytH
xsPleAsexTrajr1JplVwth+ln2EvBAIEppImA47cQ3zWCBmYSvsrI6AFX9JAAaOu
NJqgpXm6B2rffsLez3237czLw5pDDLvl6bRVVVj/KH6HtJ/EDyTQTucK6H+tKGGR
h+oKm58m8PsubN/Dx+3u5mbBb0/AEbhWux5KbvheqAr68Tb3I7UC1FyNoQyfZPHY
T6cvSVdI//aSfY0Q4wJJgROOQIEhCXb9Q0e3vOMqwamContAf5U2B81cViw93xDK
B0V2VR/QEu4A0Pvh9jDsOCQ1NUJelOthaRHd9aefPvZXWTqcU9XzuyZwbWt0zhxv
l5aPmueTBO1g0qs5hJTeSyS6YrpW1ltSI2Zf5hpHt98ErzU0O0VZi1HsMJXcYf82
x7AteRZs/TooGldlxJbhJOXkHpOXennk30y1egrwR6jyPGJW6k5pG2rQlb3tgr3/
c3u3tBJ7DzdY2KrnnVW9VqrxmqMp0eWmSc8W3hD0cjoKQf6O9pJDIfGbIgXuqz1x
HFb3fwEJKgMNA0vmBDAAqVE287DM5X8C4SB3JDNessWh8EtUxKQttlOI3T/ocydk
GjKiH1v98JwjgvHxvCzwfbu8iU1e503jcW8xM68mAdRPl434P1Y4x84Ym0Tnq5ne
7E1o9F1qoFMHLcp+S+DaQKOC1H4qIsocHPYYdbO/eH40CBArAAZFmM2/4is7QQRM
hfN33SdyO1FXVucaT9RRnhVooVc/iR03VnwRaE16sEpEQcYmhrn8S75a8TQJoTcj
aWuCR9Q7m3dkPucM5J+SeXUxKiz9R/JOi3ylgednUaiIiL2zQlzHHVDLvA5KUFIc
2a7oAVTyj0txevIjh8kn4rOhqJMoy4wSGyOSv4L6ZMUtc6CIucQnFUBO7PDQKbBv
en/A+rsIdlj8zzd42wfsMtWfqujniiYJVJYb7kaRqY5Qvb5r1Pb3zUt99zMGpJv/
y0zeVOiFJYYUAVHt8DNIUZLG1ICgzdK8WD3LyI9pVsB4tjmk35iNdRh7f/HT51SP
UwICsk8YbpAU0MSouHKCzvIcSgWedzVgozwprnGMbtuBbCaVxmbLxJFs319X1fBg
mCZrko1DQg07Q8cBDJ4R6Vg6srOHdWS9oC/EQv63rEr8sP2MF1J5vjaS7Opb8j7a
PlL6lh3dbykegl96nKMbVZruiEDiInHZe+G+mYA24Kr/c46YtTGu/dKx2t4SQACD
1nBGP7VNrmaEfHK34PGnBYerqvaxsdefxI1hsvRCWxrzegQN9J9vVjH7I0YxQgAY
52bEKawFcimiAjkZLchroyYfH6ASlDYnZHSUkWmyJv13z3PNS6wI46FrjNBrt9bB
iX8BvRXgFeVdk9KVCmRc25S3l5GBC4xJNznm1bc8NQzO/oyB/OGWQeFx43040xIx
EQ7CFiHonPWNuZdO8Wb8FBJa52cXyTpQbfAbBfpwev1TX2uqLileALbzLsqmZvhM
1KoiLShGIjGdr5KWcpWw4rIaSJFOmfiputMz7/Q2S2MTywr2mDkXlSDUaZPREGpW
w94tHv2Dli8/5ckwnk3EhY1TpMtze+8XnCXTeHzZki9U0U/0o+U47fj25oj1KYMG
OWdo50F3S2u2h2iG46j1aROGA4Lx2h4lIfuLVMv4IxN904aXy7i4n9MgD6moWLGU
DSFc6RT4RapoIL8foAnZgO+/cJnEUXDIvrev7GbRvjzBBLcFgxtRpXbW07Kn/4QA
o2hBfTrbnNrMc2kuoQm1P3xsAPXBSQbokpe1L6WnM2gbm9BY1yvMCdFuInZ7qCJB
oewqGFQY23ywe/nf8qgHOlUEGZ+Nb9N3dnRjlazSPskI0WIGwaONFixz+WGJc078
FAf7Gcg04F/kekpbi0xEXbpN3FjlR1jY3/QZcGCQhA530OOSDOe4D/LgOFNFckpm
CJATofgBJr7cGI/DO1TxrtPWCaR8Fbv18KDqlZ4hZlO854TwMVRLEY/aoO1g7tD4
BJvYFtD1JCA6HNmY3B0drPTEN5DbQb92uFZlY06X5BfOjjXnZDJJ3V2WpcqKkjT2
0kj6liROezNMU1dCu+dKxbAD2g4+59hd9asbK5Qvx698TVJsA6wykaOzvEZTGDu2
z9tZU8/N/OIubql73SE8AEL4i5yYLvbRWoDvxJSnsYRwgnaYeaFJ1zLkegDfZeI0
M46ynf3PwLah/Z+v2DmCDq9310BjZTeosU8isIsSclXwZvwTmekrtCQ5iwMFKVWY
Vk9Y6BIgatURkRT3og+cvHsTvdNQ6wyP+A/qnoiDVJXn6bM3PZfolGOZB03xmS3j
0OTiFIiKwxm+49Kgg+IkQGBv84OFj9r8CtYDNZzzwBimQOKqPQ+lAPd4ls/BTYqu
RGMq6YPL1uGqB0hct/OxmdJiYrPaZ6AyxoZe+ZPMNNyvkRo0elEW1XNyECUrL+9U
YGafOoeN0sIg2qf5mYt0Bz6kL26hb0xtcOQtcy0+iFe7O3t87Bl2riRjAuMe/FCp
IX14jPqH75ZOO7at14Y4w9W48hmwbQ0KBy2MN1uqK1VgLmun4u64Xf1kbJ5X0HzC
5hP4mbceo805dWpuvaaC4tuSIp/iikvSCN5jbYoILunQ1vRFv6X2bjvS9g0oSj+g
idGflMejFtkzHWOSocSo8Qb1kolfT5NoSOFOCmCh1i/2i4LYxFkgwpxcs7QDgjBW
yIQ38PD5WI53ajaGWNXj6MfKIMzV6E1EKHFOz7IjWn9HJyKChmvGOJ/sE7IYIN4r
I9XaPIyRGjNNg5oJFocePBTOhPXA4j74Nw1emQPlXwQ736lAm0kvnfXgnpmNGI80
1414mz3P8JFf9O+YizZaIMMYFevI6kQHLJQrOhmRTpMBemelU19JpXBwDdt62Bmf
rwX1LuoCoWEA3nBasgZjpTNcv5XkrSpIDBc0LdJCEE4itGJTUaGO8CNeh9qE8tIM
Lem9ltrAGu32q1ov0WOZXxyIGsW9Vl0FxcTNQ3RL8zwWcXvLaMRB7GLu3fFUSi73
CqktWQnGH7vfwbrAbraA3QHwpMVSeDn7h4LY9Rp0HpLmEowd1dZI2byB8z2BoO44
Ra1SBAAPlqrmFKJ/rRQYl1JA4u2/3NpadcIEfgwcvqg2PusppunF/JCUnfJUlUM7
oruWMAzLS49/YpGLOLsmSs1ogr3OIE4ZGcYiXdBAUcMJ1LQpSgnRdnCGm7Pc/DJe
8OPbeW4EoY5UCBvmceVaoysRSYT1DjyfGDEuYwlPHPJ4QMeEe/jg6Pn/wy7x/uov
/VmdEeaoD+FAtD3PUb1AqnsE7RRLny87wi/FdxSTSvctJ+1z6a0X2nlLWnSVz1IO
OFv4H0VmsM2CSmuchdGakJ6KVRozJN2upgChYuPoJORHSRfiAbHb7p1QQh/CZhgU
enEuodxtqOTtcGzSmG/XfeVqRHNOratM5vgqLPox8NFjFf0vviueKavJshlAPAR3
R6o2HG5HF7DXr1VgVRPGx7c/gA1nKHg2qFyXFU2ty6IJiX8ywq/KRRhbZ3Y9rrQ7
1PELkP3N6CLGBoSM6GhA3nuDF5+veZDv2ciRQlYHO9yAWDvCqp15nJsuVsBgSoyB
ZS1IWQ2rhn0AuVRz+V082FH6ik14wqWu12QcDkD/kSbpVYxWS0AydfTfXZoHIr7L
nYSinqnwLPIFtdleuX6tqyFh9s1UlU5Tfycy1NE0V0HS2HJujDggF4NYUr68lMg0
1lWptGkjNi0asP4W7RVTLZJtxSTRJc+8O+xkRoni/pdPtGjF2lnhNqC72HY5Kji6
H6a2tFf8tzTabFe098q41/1fHR/wJm6kCRIEA819JU/Ztj/nB+G3GBAfE3bD4R+s
F5fqcvrpyBQxA5pxLfdo5STZG2uMo6kkbAOpAywP49mGIeAk/Nbfn2glgu1NxS7u
VyaUZjcV8cmn8BGTQIDl7mvGPysOVY1csYckAqTGSPNlrBp/3hDJjfGNGEHzXLuc
3t7XjXFLcMf03I04uyNczQEZMp104vEc0EZEemzU93N3DRKQsTvh+mMyUSwUlPlm
pxnGJCCQS/OhmKMQS9Te17GXRkasHE/1O6s6X/cd2WtqY6isRLjFa190o/Oj/oVb
euvqLeTrdAgSl7We04qnmJF3GSeeRv6ecDGDmJR3AtUXCGYQS/XKuTmy6JkHVQuW
LOAmn0lq5L1Nu8AXYYQqrcTwAQPZ1i04g9lXOfH40YL9Hi6FYopuSMHZ2Znm9OFk
dedRYow6bZ8x1OPHcPXb2fqV6qeMaifwr6FV/Idni8jrbD7hlcP9NMa2FebkBJQ/
AOHZh1LRSSk+UL5tbofPs+SMR/WpHNGNFsZn8DjEHFen68/VYw437sTT8FGXBcaM
9xRPwgAWw+6LvKR05HrtJWCv9lHG6fgB1xsg+6YHzGjNcn++28nkcBlcGOMuu1rM
JhZ0QFFIA0uUnVASrXy7JVjqe3DPDMyoongSilwhdIUa7jBTDjwlFhd38cqoAwy1
aEZzbqCZwBvYp3BSZaWwpvaURXVTiugrFlcuSR/6+itZtaPbBikhoz04UbRfZn/l
NxUt7LME5wgQtY3o6E933dqZiq3uo2kdh7UrzwJUKajlQBjNI2ME0CmI12q1c/JT
XHzPUHCkWUviVAVacZFeVYUz5E27OKgh5VMo8xMLvhtJuDLSbvuX7FIS06CxHmqW
FrsO1J229BNFPyDfoekJfs9k2WzM7dNajtN5GuYQQPURQOk5soi06o9LconBLY74
e5xZbB90Ev66QOVSM0YGMnpTFW4BIB5rsbm5+t5GVDnxXu15xqSMJwi8MrihaRAy
sS35BbUq7cdZn1fHTY89gk8GTj3uF6fhyBlA+jcp1mGD6zfgeU2qkIlwxN8WmR/r
zYwulRGhYD9RAyNG0WWzChv1Bpi+kMZQ5NzoSVlQZObA3mRdG059JD4UOfcP/1i7
9nI1KydPv1uvbZHBcmL7QPhKHOWu/QpLK7URTgXpBCVhnXrUWU0kFvCHpfDb2fWu
IA8Ghy8LVYSEANYHF/5Pp23aD+dY5OFhgEcqE98UCym5Rv9ykih/0ubEtPkNGrBC
7Ha26T6BdHKFV8sW03YpaA4aQUuDsiRhM1HcqjgUEIisI+1pr5wE7y53jg7lj58n
9j/3LLagblcABE/YcDUQggUyZIlvfDoatwQLxiNSGiZyBI0ammLvbe8V28VNSxoz
IWoqDVJWUMXvA9+EH8jKrLsiAmrwAUfEbuo0zeKhI5JVUkyLHcjgVKJoo3C4dNgY
LBB8RPH6sJfNyGJNYMCxp7km4MllLT81VFI4Fe3ZMDQ7SPWe9RBgBZodVTgNH/H+
rDHLVorqSXAqldaEUO6ULDUZi0SBzN84oQK7P6ZQczJRZ9qLYK7Q0fEZV+EcdF6e
3oupvNtxCxZS/GMfDUS8DYtvfNnQ+S6N6fm27cj48Vy+Vwh7EbvKF4bC7vX+654l
zmJB9NEj/Db57n0q2lL1LPx26FmGmRmifLkbjK0G43ElVFD1giNVsjyb+Bb588dA
IkFLRPP3cw3plIC4e8Im/r+Hv+1wK/koKghO0gXIk5eIKEJL7iYsUH+R82sfDg3M
CMuw9bqzGRqCpxVjRaK9+z4PqiasKA5o85/IuR0a3aN95qcplOrtgptgBe7YuH++
yPAnRpNJ+ANmhIv0bhe6hukv697P+bfAXrIxQkxl3I2zPV1T4SsOz1r2f0koVM7q
NmMJb0o8jsJA1E5FUVqJ4CxGvebEPmcytEUDTfgl23VL94O8ZiswkmXk9RGx3qTC
pWR3VSwgYjC2acFc36q/RUlstl5ZWoJlIE7c7VGRsdNgw5O80xe5d+8cKbDOhRO1
Of/VB63ho4MGHEobieGtchczbA4Khs11Bzbt6vXI3OcTdOqeFG80QNkYDmlfUfyi
XExMgMBLNwtz2xe3ZF+FMrtCH/3d00663tesM+qbubUiNlXQ4zxB9e6F71c5XblS
UWviQae7qPIfcQs+PR90ZgE5aTM2nDoRkP3cXBqFAjcUtENFGB9TO2y+yrDfWddl
wyaKYOuWGkmlmkO8XOTtkZFNo8p78JarkLECItN+gZRoS6xZdbRm4D2214yOu8Tu
/t35Ykq6dVh8D1vVKm6mPlqW2iR2ecVL1U9Gsvqn2PAekhDH43BilHQaWEqTv237
uS1/4/TJ88GfQ6Sef+ayiFwHuwhVQuRvnG6b5MYLYB4G2WVIetaB6Zi40o1Z58gT
7dvg18mKHXdehXafLancxmy72YDctAzws4FTeRoYdufUV0OlhPilAPZJ6gf38ggp
e0zSE9b0q1BpwLAb99xZZlD30hsUXSypg7vJ6NYqCBLTLEUrN3QWEGNtDEp/8tWO
p1pmL1qTVbU2aXACH1RenukXW9DDu7XTYttEAAs6XAhcVDOzHPp0r45VW8Ot4yZo
LM4qsOV8yZi0vh8HcUhqfj3G2QE6+2jLYHrBpg5SwPLBMxYJMHl+0B0jlUWq8nb6
u504KUik50ja7AdCwdfc45GlsbP4k63YLSJWwqBfpTZGK4OKAYIEdsDRxE4jlA+P
q4RxfhJUL4B4dAeXMtmT5ecoftSEkwUC8+/zwmsU4ItmumYMZfoV7GTX5lHYuBfX
lXHAbcOBiXoiN5SQ8WWpSgOVj4X6+hAZst01gU84MHOJRR5ZYpEbaPB9vk7CBv+Z
8luNaYrkOnLKfvyQCH+D7HvAdX3vJzM68J96KdFqazf1TFMa8p4wbtZQBJI2lYXF
Df9Ca/Y9Fw5YihcJ1kj4NUlbaIAOox46gwS1OxCpXcO3WCbGEmsVmHlmZ2a06Mz3
kIGkfk9s1ZXtYjTOpkcZCTbE6mxt17oE2Pd8lttnwMBNrai0gfvqlyRjsvlAuRTV
AzKCRtUQjD7paxRazymVXG5Vw9WsM+7WNPk9Pwfdu6yhIP2nSu4R8sJe5D6ICcvE
RjkS4w9k5uDWiDKVXUloW/8fEh9J8AlxINJ4SaYPCQlX/A6xmc7t9K22UaQ5eOMM
+kO+8nceKw0xo1ZM+f+XGR/yIGkFLHdZ3QLJ6LxhOnrbF5M02tTEwXyqTI7gdXFB
BHH1eO4zIeYkWZLQZQhzVrClDF+DkL/QwghdCArgAHbRZVHyTDvg6rKg955Qrq2G
aAxBi31yEHw48g9sOznB3/lwIx7ShVWdvJmA7yzfGdLH4+Py8sZQ87IgLw7ewA4J
+V0cFQBHpwCPOJ+qfndetx3VUDbKgfWVgAI9Oq/SVG9KOqIv2dGCO3w7tvotIvn5
tJGohjB8vRWPyD810R/bjVYIN0bLwrc0u9ICaqVmmNhX+hvj2JoVYgkar+7GHmsd
mBpITONPUjibo2tDKMn6leMvXt0uFd0meYyEVuFHZwTgGFxf2iriO3Yyh1NZEsVL
fsu3/m8vPYpOcyVEz2N/khDwSVo/WwzzKFqrhRlJj6kh79Y7RrfKtGk/Tm6TApPN
KiRcxdP7SozbA2azaPuE/S9MXd/Yq0MfdvczDzYXiTZ7QZpjCF5N7wQ4DP5OcnHn
4TuT9afG09ufdVSWZZu3lGzXEuBGcJWntVIgF5o72Xghsg4E+SGRmRbDcnyDs/9h
U/4t3J8Y1fbNiip5sgIYc6cNGou8fkWo5mhR24O18oUvn4Ld215PB2KCeK4+A2+Y
NyjrHET6nJkSAker9wR8dYo1ZoyRfCVz1eoZBxwHNm9U29juVkaM7sJRqhi9STkM
BgSUFkxAtC5mXLDQBqChqH2eMSgXx39gGALSh5WV4EmGFTx0fK/rvSLRdGzqGsXA
iD/1rweX0+1UkzdzXYFhmOf5lhaqJ7Ic5Cj/r0/zQg9fXxoHqXHW8sOJEjGD5QQX
GBPHbYMHl7d3fQOrLpSHKYLy+LtKzMKPb15qWbWmdpWx5ClN2UNtV0YmUuC3eHjL
mBsVaikIpyYygTciWPsCeomfIxUTtZvlDRx+BVOpKA19ftoZs+WyFNEeaecDVEy/
ug6GQmdWhgn2k7PNRCBH0OhrCdYfgBY0KzhD/96GeHBFdKMkFlaSwrHvD0hoyb4p
+dwB3waH3ZMyrYZoEuHy7lL9WMBdO72sNyEfboC3PFsmWojKWNamzodk0hpOt8lb
AgZqfUZAfjEYElTLE1mnr8Q9l719ZZMcXyxCzV1WK3W4PbrpLhbE68Y1eNffju0Q
8YwtxfcSEV1HZwIVRP+/HEuVActg4E2zpg942tuhcONtdDbjxIpf8/GsMEHZpi9F
x2Pj7E1oQNaCIljXCBExm8hVt6/e3Y8nnjxxzOJ9poO+uoquhtHOSq/VBlPfAOk3
x1RN7HvxJU4NjoKvCQ7uZ8U+XvFlmYZnJDCuOc0Y9gAgizLG5/Wxd0cuOm72PyuW
Mu9H4mCPrq5hojn4lQTbohWz2pmaFspVnDSRQZfT99gHJV/E3E8mmFqzZXOEdQvz
LTdbF84h4NOT3KTg6LiQ9A9/1pV99NSzIUx98PcYV//xwPo5qaop2a7D5iPtk9bC
GG0R3gSCSg2MhRgc/0posGIkDotSdiBD0blQEYR1D71SJ/NhEk05gs40tZjc1u+i
tFIZwTiNU2MANf7QBpnPlR8YJV5Hhi208jKWSk5XVYqsVBaBmTkGu7lTclrjDXnm
kWlfgHclHAIkklUmcL0ARsq1H62B52n9sgyxZFyt3HqLMxpgt8IY4FPnljoKlfq+
449qpcFllLixeFn/OC/UVOj50c0QEqnCuEokfiMOQfD50qkuDOUejJk3jP7FMLoy
I6XwWfdg02Y2LtEGN0EMzSIrTBjcwJHXV2lk8zQWiHGn1gSTeZNgTTB+deu8UJHj
MvQtipajEEnIuJwbAq+gtA1qvWe7o/MInW9A6N3PB1I7CK7ikwnF/H1NtbMGuR4w
OVSNDRphL2sjZ8KCwouLMxoIkAtjkrkJ2sHID2iXiA4mOO51j89YeNAG9BYNvuGs
LlkFWnpWSPn9UrsgbP00+HtBg4giOboJyQ2ZW55PUTsB6UFl3rSO/YTSmRXhkNJy
ppja9GF63c6Nq9+V5Ng7MomSTD+CQLRpLM3Y2JlY5fDsblucLOvABbrvZiMGIvZ8
g5yiDbo0klrZLsnRJcQQLH+WKhkPTy7R/lsmH9EfYzXkRWD5TWmn7mx/r3aSi4uA
0AhLsu54k3MJsBBhPDY1oaztPqG49h2251D7/HeLoXVdScBCWw3Dt0jobND1I1cQ
HYpnjBe7LTIRps1R1KPZpxoMRLxRIDGCULd70y04Op5HX/cexRxht2th9I2NfZFz
lsJl0MVo8nV1Lkic94HbyWCmvYfs5mKojuRWUu7lMqZcbwRknuInP1wWOSMa/9HH
vgFGnYxxu59I7B228gvDgN4aIAzoRNj7+xXz0PfngvyQRIqpn+oJbb7JWeglakKP
G4gqiecdywHPS8LF2Ao/cB+SMAZmozjVZdiNGajyVOKPYRQWS3kQmLUd788cFoOm
9Of3tlniQJQUZXAaDMM0NyyIqsUVD1W/ubhKu4ZL+oHoqg8WTj/QhlS2ooVUPESF
yYAhb5VfmjAJ/Dh+bmd5sxJeCNcPfLziDiTHkCWXN7JCJWnAqB43iR3OUhQ+X703
zGtDc3YRUvUhGlWLHM1khPZBNSMKKkhxyTdHm78rhznRXYINggOPcAjbw3GZ2+Pb
zGUmKCTx4P2xcmPoz8WyZ/rpAQ+eHNbYpwJSHhXq7jAZFa1bcISZbNbBOlrnd/4m
uWPBhjSSz9aHMWnbYxTdlH/6vVUolttdPF0ZPmOF8y8iqti65Ar4Hbtavb1GE5Ht
Kposg3ngMyWTg2KN391WjXijiFV/KDsUtdgjkxKleIBbKYB5ICYDY2nb4x6q4K57
SK0W0sCOQs6M5OvPAPXvDYjluAunmyhOr0Ihx8/9X3+8vALXXieb9aef1hFUkkJj
/MqLqNTZhJ0Gs6F8a8Z8buSbyatKm2eCcnmZcxIu/FcX7LkOZjLj8zi2DANLPs1L
E2av2ilSv8AS+6cm5svwQEGg37MIXfcXqkVCd54XHTm/noVxzUaUk37QFWEzDFpa
OLGBF7NSN4tmZPVTpX3qkhsy3oRiMWspaZaSG99O5/fFIQCZFOLYJB2/pYq3QLdo
zyuEmNYnEqjvKcLPabDv0sIRXPwz0Ss4rP8FxI+DsMQolC2rGaoENT+ae4swSEy4
YOPyyWfG7ZRPd61+RO5Y00zEwmfCINmJvFGEiB8T+HBVhTahKnKMlaBMwY5lJQm0
FCxM/OIb/N5GmtMN6FX5jaH5rlulVw85aCStiud0PG1q6aXqZIacJKzj9SYCu0xJ
kmlqEZth5V5mvrsyAlAF0dulqFC0jWE+v0stcVMZLB9zKEuWEGOY6IEW10WD4Y5H
HWq81hoNDCNPVlybrBr617+b/HSP5GJwj8bitw7ErksRLUipnqa6mQ4Bua6YRHWl
+I38Czt9zos1cZewLqjaBfTzpySls9vXl549F/h5v5ponp63xBGQyJ+0zTmSrd5F
/NR1ow5gheJq4ncLwrXJvBnr8mSu8ywOXRg8O+XzPrlU1a6w7kvugn/V/yIFiq74
kahyICIIDjW64FYxIYZGlZhKeDBlDRhoOEQtjjJNIIZ5Og5gqZGX8MvOHkHOPEzm
KWQmwHZMgj2cXlF9rAhnJy4PCeqqtqH/W91KUSDYoCkL3t7DPT5xaskD6HfYeLJv
ThnmrF2g0iL9kblcPY1yRAzujxvTuCVNiJ0acm5M2HkA8E8VGKeW7IWtwv6HwVIo
47G5lRYE/xDTY9I5tZo85jl1QZbs1haOQyM7xSTEQ0B1jaZ5uOb5PzmcgU0owvHj
0VYUAuQl0rT8ewUQSpMPYwuCqNUvp2np9V2RUJuRiHBbDMiwcE4tNvu1ykxt6a7c
9ds4E2H2bbPoFahPQ4zjgvUQdTD7eaMN3cGl1QVfrXA84OktIzfege2Y/IFijDwm
kZfhAD7fzx7WA1AT4mU1NHgeOdlIW4CT0xe478AYAJ1CHQwScrFhB7y11yM+n+vH
Lf7mMyOgKde1+A97Pu9935YuFgpc1s+2rzV/g4KcwKi55I/p7koiCIMwLQWNfTNw
SaREmJgNT/AbTSLAICszfuGUhfNlZZkfOiTD4S/dqB03h19eLiyIGpBDDhKXyUr3
gjSCcJx/dU3d6sCB708jnAk45ieNbAUDaOGBpcRsU8FEU6XZLKeU/3TANIPBqMd+
Y0HZ+ng6MfEexb+SnHo/TchrjR0oI6IlUPLik3eRyzmkklRVrfZpZMpVleyKS17t
uSqaLyXq0G8O6zAwLkkss4Rc3uSp3b2ozJklKT0sYIsfcBCCW7mexKJfs3euPaO/
ehmcMPSbOHe8GeJBWsHwFYQvgicQHueXb+3Ho9lfmaKJ4uzW7qXhfqXKH6lTLtjM
5bCAMC9WO2U2LE+7EP7Mb7YiSBXXRDVcU3k8FZhtVk7AW2mrfMTqVKjlR63TFBDH
JGhJ+t8T6nitTzZzr63iJ256Ohe66U+RJf11Fb94CiTtlxbeevy9imOjkBVj8Bwf
w6MaxWiArISuYrqOHqBBwtOHDUWneoEezQnCRAChzrb0MnnJm/rREVPJFyDE+PK0
fM9EISXBu57oMIZvkQvmwo/oXXkLRqLjTYG4uPV4IB0w4F483APxGR/R1AEl6lKx
9FDcKo76KTI1ZRUlMIno5Rb/V5vX3Xb4Y7YgeicxZod43sV2eHcCGq76iUUPgLsg
NI1W2CAnCzuK52jQSOR3KNkjC6UUAnbflQij9Tqgr2yteeI15YK0+ZzS55SfdjyA
JyWQVgDTV+6CL2LxlN9s+Y+EoPJAgLH6q4ks2ncGSD6S+pGZayykUoV5wkkragFm
98wOOwqIkA61D/IYcjoa+Raif3Xbc89Szl5LadISgAo+PjcKUeLy3ORBi4Fzhgpw
zRZDB44h1nq2mvMEvEplrAg37nZX0nMJNM4LLgbTfHV2MpvWeUQ5q+6RxpsSqSur
oRkjm27NnS0ERQbhu0X5dw7MoExsSWgdIVIr57CVVUVrG/5Z1yCjHPkmnCgbe6Pn
asFXkqewY/eU3fFwathAXwJgrRjYuoUG9NWy6UrOKfzNakappOUgEfiLZk88ytjj
qHYC5BCl/ZtY9jZyZkHXE7fot1vld3Q49iQnXQJfyaVRhRToN7//j13lUVBT/fFu
HH+QhbwcaFiUmN5Ar0m9zYnT326cwgudxo2XiBVj3qwPPSBwfBaNjoC8QwXhDSlj
CGJbJgmS59mNH1j6rQ7VSR0rFUblG42FAQ0DL6uaRQbLe8GtzNQHpcfqzxtl1Vlt
dWAJOiGgRBR2uCcXu0sRXeRdY7B9+G/eBSa2p/gaHHKe8HpwZOsEoB91v5rFvbuG
9Qtl1Fa54ZlGeIJH/CmycuIOf9XjBTjn4C+p66roK4kc6vFkQJJbS2oI3KeTjNf7
jUFCqfm890/s1HqPbvM6viJjCapX/5618ukG7wbJhMkUN5NcrX1bIBABmCy1SEb0
f3GoEer7ahry7iJ3Nv+XOzHNeUxtYWE/StEwRaWytYZTE6zjzcNHpKHL/9UCBGiE
Bn2cZIJFpS7yvpFDV8n/3DqGjL+kL6sDlP5lmnWt5U5C8Oqji2jVl+0gW4zTrLNl
OaIA3PIuppul2sZnlKvGCnD9SVzMJKF0SXOEdTTArIOBPqMioR4VH4wdzZRfJRY2
Hsjpj0516RiduCVUpgJA+au+1jNkU1lImh+411NTGqYg7KDqBDZMyr1e997xkLvI
y5He2ZsPxSGJYMaGFn1x9fgoMfZatgW33mWYbqfBlKRoFv25ZttJ0PEnMXwK6QRv
ejWpzAdBQJMkzX7IWFSBOi2Bzc78yyi7M9NAzANzSrFrIEh9vj1OCo07ct1xSDRJ
bjwgzeaHsYt8xc+UCHV6mpfSgOoFl1EzGJ97gxrRkUE0nH96e9CtQ5+aDq+qSMpO
rY8R/ThqO+cbkNj8/9TxFwQxJxgyUF56uT6o1ojbiA/9+lVYltPN8ySHREwgFksw
xqKNlaaiGbdsmIrQbnQDoa0yF4u8y4HmCAMap/JBte0zFp6c1nogVTIsx2o+dHfF
EaUbXIhGJwQ/sN+nCk9vv+tneyyvK1n6ZJuRZ/dmsLmT6IPFoqcczSsbwO9y6SV4
WekEOFue/1EiOvQgVFcF4IBcgt8qbzrQxnzlLZCmuKervMml0N9F74oMMJY/C8Ei
Psk8xFOn/ubipfhhHM5lv57mwrfGcs+42b1cJjIhG2ttSTiqLcXlIRZZ6R/Upa1D
vJJH/wJOWFtcPqGutRJWpwaas0UY4byP22Ra69BbDqoX7bZ8JvQHNoOHSTYdfak4
/TwIT5wpGoQtRRLqU33NxHS18X1Ld+wKEWPmMIQagKTU7cqGjLoKkg9d9Kl5ZnlE
gvDKikzxdkOdptVgA4i6clJR8bN7j2KzGMDdfChYu5vGV8Cwv2vDMy5SQVhhlsXd
pxxrEFLMs70SEGFE3nk8jOXHOtsskpBj2fG3FlRlXpYmJQYZkRP8hoeoXN+MXK88
5+WC92KvNhCNMSf94nRBtb3+oYd3gp8jeVt9Oj6Cvyse4Pa6HnetqtpbdCNMNEie
SHyApX46IL3miOiMdQWrdIDy6aSCQOgSb/CUWVPs69atYZfjzAQJfbzCpKoAUWod
ZYzdpg0za6oXXYZGtoYuxMnc4YP4NinMk+su3lwaS7EhS1KRDcRfTUKr/884sVqT
PA4jZfMyZMjO+F37iwhby+B7Wgue4gokFdycng65pjblztXHRWqfIOmRXjBIRENq
R2Mw+jnkOTowyxSzGxhghpdoxhecd8KSJbcSLlNHxRYh/ICWK4w/RWbVAXbl8WX3
A6KJqAAH3Ffemuqd0hNWiSaENA6zdQ9790ZGg/pM7qOcyEa+lQeKH/Vq6EOjtRxC
7oyj8oPOvpllVl9XrmyAtmvabE7K47JKrCKlENnRZcSW4lUIRRuvCrI1CgpMuyMF
oZxSXP4mA7goCAoi2Dq8aQZ+Lg9QDmG11JLpsmsCkjjGEvCo1CM3IxGvTa6+tevc
jiei50X/+enkh+vJI3feTIykE/Ql7xWMIPloFgN942bJJZGT1gjzxS8ZJGm8KLha
LL7ZP7i3KXWZF/v/WsUQ4YIFS95ENjT92mEJ25mrJ9zSiPF1LGMDJ+okm5mtQsio
deC6NvxU12/2JYNmp1+ZiVkI6IUPe0bz4HveoHuj8MsPOR/bXeQsCwGW9rQdjplF
YXTt1f8oZ5WPrkd8dE7Xdl5zhG5VId04Sk5gMrlUC0Iaa0Hwht6Zqy5aDNtNz/76
Kk7ImRvJAaCJYrzq+wJm67Csy/KPFLAj+dETrX9OV+nWi20CPfb6ppBc7ZgBX+yz
sQv+0PvhtvMe1o8eNXErEHQbpyZDU+Qb5Yvl4VC+ihjZ8WjysTz06WHny+t4mAwE
nW96souYAuOIQ2geXJKFA7Fllm49hha8AQXj1xOsy4WeWgbVS3mLOXoB7Gn09iZj
KAgmc+ffeg+5RlolTtJG8f0/BKEeBYKbi0bt2gGpxj1fA9A3Oa4ooITLl4sI6vxY
A5np6eOp0NEc86oEik8lIajMb6uU4aAEfUrPW67e/N/BByBvlu/uEk5Pv38CavrD
etoyGArdE/CZDoaJz8HrG8foEF1reSbsqdebn8uzJDW7YhqdHK8HjZcMqLbQDA+V
6tXXwmqkR5Mx0BfRULeyapqdHS/398f9ozs1Fi20aPBvGNh19j3VEu99/Qont5+y
8ZydSbBb9aVGUMQY238kPNdc+bCeLOxfqg0X7PGz2EG4tYzXvNN9H4N77uUvlCm0
JfOSK06iXgmOaodphMAq1Fjwai27bjQXA9f2AUGLM0LMxCy3f+Ah3/srzjF+mLr8
s0m0OXQTydoEX8clo+RV5Son8d63YLPZmPmTc/wvBivSH+zbyY/SpojqcFIWFt/N
mLeE5IbSryOBlFzPrZrKnhzsguDnpDosHyB381YOIUfxp4Sxtt+RSdPnkXRoae59
HOhrSLCZ9lRb5EJgm2V/nUmkz8ieNjVgp+J6STtQcW4KYNorI5WQL7oDvGkLuo4R
BFJS/OBUFaEetnVkZPYj/DdLGoQ+z7CpT9vND7xetuOhEAdKczDTqjuYL2kANYn4
fvz/EqbwfRVar7GhqXCUoiK70g8+4EGWhQ5jntCKb1OuT6yZEGzgsUT4XvQwb69j
QxnVY36pMaqIyA8cTD9/5XwI4cCWJxLOpcK7QIdvAoBJOParUcGgbCmunWXBbR7d
tJALRXL285TE/rMcZQKfRSbtaxTAKTgSeX2vUeLv3YJC1g4I7OQqCiJ/3mQrGGQf
WkAfrdAFHaqME6prZTWKFts5H97xxPii/oQlwRlNka8Pn9uhhLe0XkCWY0YLxFgr
aXpPVOtpqICM72V1NGGOHq7N92WkJITqOqB0vfKAqP8xwPcGgtszjDOkG4ch7zFR
49tG4YLHB8M3brht0i2aPxSs3VNse7N2a/bmXYGEUCStQ311ZpLwE1JX8WA5q41x
d6HZNdZJQ4wPqwvqvBuPVx579pO+w8OqAgWbDHk7q01vKo6M6XU6vzK1txDJmu2w
HbAZppB0UY8Zs9Fu5NAFntwkZl2rRe9D3QzAXKvW9BddZKtR4NfDQiXgNGCrmEdO
A+KRaUFfpVCw9/BQPg0Tq94pqtRrZRvUCu3//royBNYdk0+hGJKuYDlvub4eMuun
gT3OLvfaiVpbR+HCfIMGmdV88YKzkJcKm1GZwIl3Z8C2ZXm0KpFwaOLxUqq3b92q
lTxQ1yPfa1/j+TEyOBLCXZYgOE49sSHj1W9GMIXTLHyaX2m3NoZlK8wFGj59Jt4D
TXiO3qIjlThwYM2gy2719GZIbbghw/e2sPWzNLmbGlYqyIHMdrwdfA1+Oi/Mqa4d
GxL0pPY44+kexzMug+KAlI2yACL4IjuFIRNTkdD5VGsfN4J8brbKs6hjQIwkpgAp
Ds4pcPoMtaoaeCcrsey4MpiC2US87wYn8SmXzAhEjXltow+KwsYSeffKme9FicVH
S7SR6OZQOdaMDcmOfNsJi7lSUZmGgkwsdTEaIVdhPPq/tZo0P2F05ZaisVUBGJzm
lSiiYIK5049cNPTCQyWdMWBLxF151DbUpe2tPrngDg1HnupkZ5bt6P4+XfCwxfi2
tNcI0d8c9V20kuCWEKinHM2V5kessPfXDljuSLfgtIgmkarrCSiYp/GtW1DTCWrW
N4fE+wdhqqTB5ZG4apmKATgLm6V9d/2KPy9VU/fuJ/jIoeaN9pJXuCs44c5ap55c
oPVks7Nyc+Hzu46E+wITTJYGdGFejNPibsaJR5hjTL6vGfWHMsKj8x6GsavTQNw7
1v+AYs6Yp6KO2U52NJGU8A2NJN9spOD6xuDhIMBMjXeDBx/o2vEFztYqcdzrkvcp
K7kYfVszQxBAFtf5IMgj2bQv7vncbGVn253VqImfoTEk7gTPYMhUQvm6LdqOfBhq
9xpfdVdyXYDhBso58eXe16Y4X3EwKVpGs+spk1kK1UGYcDUuU/DbotqkNxYQ2vL2
U8FCqxW4psVeJsCdoPZFgIdNalVI4dfn/WDWo6CbwPtyQNeG7j/TJTTOz7tSp95b
NVGV+LNijPbRY9cF+e6m2o2oNAHP9wywtb6uGNsueJDoVmstn79Ec8hWYiwyy0Bo
hkXBhJYpWKMet44eSx8yYxC0m0Hy8HU8+d0YDCyF3KjQfNA1A7G7tmjNZIycl9to
aquDT7x2mDswT7BqhPIRKGGWZCYmQRL0qnLVeD7UzkVxy92XSPHgiKRwGPl8Zd+U
NuodCRl+r0gkNMn0DvKfpJnU3+++cDoW+PorB7Z5I7tq4f1M3kZcLIYmZDkvd+DC
Dx6rxTqY0d31gcpO0Ad3R4j5Os8y0WyV1FKST9T8uWJkz2utxkebB2e38upcjtn4
CuddvRZVVI81rQDo0eodYB51Hfrh5rhBxd2tlvctaQ4JMoKzU5fjjXxCf8V3RR+o
F536byvsSqiPxjyuiixuS4SelOF7i5ihZcCX8Knn7ObLX+5z7c73cSD1JUlsbCL6
YgOe74rVOT3vSwR0tMuv2IKWBNTOWVGB4EOS48dc1TkexQ8u0+bBkdn3IIsYKOgo
rAG30qyZcKkeF4QKhj4AYjZStoTr5kW/UuH8Ma+OqQgEr7ch6yKgpKmQZXNCW+Tr
wMvIQhB37Lxk2Dzio+CYOP27MKRe7HAz99uXaO699TT8TUociVDxxpy6M8/zVY2C
Qjp3g/7ABuZxGXenqo0RKtHJEIi6qgoSXP0MZcsZ8wU77Lo7v8HpJ1qmex1i6oK9
Nj+3XnErolzwUXXOzE2RN5l/D9mscGiMjsxmdgnGdx3ErMj/bi/agtzTDVQ/pshz
te6L98y4STPd/voiu+XmLlkgZjrHFOVECnztmiAW1JU4wXRJFyLWfKsD1G5u9t1b
P/S+kUslPx/xvjFFp+8K/pdFAlzq3XTNPuyzMYeVnASZU/WoTjqhbmWncCKqu7dE
FqOFaD4VGd9cAEQ0BkUtduTlxxZxkE/RMxcosZHICdzCpDxioYcguuYOaRUrHwJV
BlfNizGGseKzH88tsUhLuT2ctMFn91MO6vSE+DK+wR08qc6A+wCDXOyAOu4hDqST
mmY6Q3H5W50aS8nF4rp3kHGRcC4DQD8p9KXXC+4WzUsIKYU/WD1yJ39p37f12LiE
ikatNW1uvbO59713n9udF7ltNCeDVUxaH9qXcOTzwMzgfEjozdiGxljfqlqSG3qs
6QCRvGM4msLj/CfNQKUsrHrdf7Px4kkgcUM18H+9S6luIFQWNSEHW2ovX/pcuDYm
J62BJharv/ISn7G6soadwoRV0czNvfI++7UjL6b9PUhvB6wzU9UdQlMFSQJuMOcS
RIcnkzUbM7SjyPK+c0hvPkXlriJxw2lw7IB1GbmQYefSkIu/g9AXIqGzR0sjQ7ie
65232vpKcu+hswYEHqAgpNIc4RqQsLGk1ZYoj7SFl5x8uWhW/aO/oM2mCIiUmmok
sDK46hkFy0948Cr3qNMJjxoz+oqCanmgG/MhX6KsrFOzH/iBJmkabm7NKt/K1huf
LWLyKsJjD5eUzrG7x5A/0kTAUz1LTXho7edTp/8e9ga+3r9tJIhsSOzMc+PDDj6F
bIqg+8jvf1R/aOILoHV1EIbKIaxxoe64RUEtfZnI1dDztNg1+K5d/1IBS5oKVn3q
o+RfQSG1rBMLzlvaKdNEHkFRKy+uS6LMOnckaRhTUxaXM5NnRuiut8kUSZ9pz1pn
6VVVlSEjQcM0d0ej3au1Q/GFV8xzyXSadSSIeWpcEpksU4p1DQN1/RYnN0F/DM/r
JJlskYxAHYjV9fa803uDLEMIL65ZfKegUtolqxZrgxXBYgmgxdksOnMXYYO3yHTk
M5nAkCFVfRMX0B5QyGWomqiuWMmn+5xggEQzLKUqyWLKNPbatPCENyIw8szRD+c+
Dm2nroYoP0NaF0T/ypC1lw03LQ/a228Htvb72p1aHixYsh3F3H8IiZw8Y+bugnUs
grBcCZaqmbHDYuqXks40VF3byCcAcYSSNJlAqBGgnGiwqNDZ4ypF+U7/lIEb8ZDt
HK/tbZIt85JXvb9vK68RiO5NuOZTB8knr0I6vqt5RjhpMhw3VSSOs8QOOBE6QTe+
+ICPF/JYgrzcmntLOy3EJ+49zoVzckcg5f2t+7EOGwFK3IYT4RDQXuzAaLzvidpc
11cvtPG/R31bu7GMcLZHDmmPEeW3x2GPdmhKkQ5rWfr/Nn7uIa++r5ov3o1XEiaJ
oMc6WX1mkSK2GVVfxhljskDltaWtq7tu59kOnPdvft+cbF7ffJXpw5knlpX2k8nd
oAf3TMMpdjQ4++IbOP+5syeujsDuTnV45s0jowpLz2LmXT9B9ej4zL7w/mqyTkzT
sDn3v9bxBDlo2g6770yDu25IBtITiCPgwRemV0qw2wINMvof2/5MgEDITBQzTMWw
tEzQr9MxOdxfDlYcaEpBfbCC1mg3HtvQidcSfIxfilbgqrNYRS+cl6EwJWbUI8Z0
sAu2ib3GXm8mZPRLU1945J+KPy7sIZLCg8pYZbMbEQpH6aVllU66V/41dikAapC9
47uxsyLyNGa66o04lp1uahgvPQm+5VeGObspAbqXrCek4a2r0UUeokK/UaOYEylM
MJPo7kfATj4ru32/NLQvpPSGRL9a1G5Ne9fP/ru9lovrmc7jpqw5e3Ob7hr/C/+f
6IKSmhzKWXT2FncPemjGI/aBMlUrHX5XUZY7ifq0EuIhyVzFoKCEoybZna5VGc5/
FLceFXydMJLlUT3b3b6cJp8VEx2+VW88kId777TQovm1Fm2l6qCKiPMccRnoZu94
gVdXEsIUZMHSnWCXWkBPJRLlxU9q1yuBy5lrGH6yEQ+LXBC97sjNQ5JU/Yz8Myg0
6/2cyGXvXMUJlXhc/xmwanX2QuNHfpKRF/QvEepB9NDRqTHNih3r/yszBcUI5U/r
RIQtznDuLyz9dE4b5p4hPawlJ0C8lodOCaO5kjL1ZeEAzyP/NpfPNlT1Ew4w2w2L
YPaeYIh0B4OfREMLWv3OJmzqxhiNYD3EbTdM+R/7sKkj0EKtGp41YGG55PjeQaAI
tUlQ54X7QKAH2lS7PSt7Q2/N5oKDKgJAidGZEScaB1rdF0FPT/+WjKoS9sNVtMNo
lIBvn2X7He0Aqkveqr0iBqJA+Q+/Zar1/l+N3IDXmqMFhQjHbPcsc/CbydUcLRkJ
vECH7ReFvQh6sO6NpFARWvb549qmYNGpIH4S4zS97hJQpo+vMYxk8i8JCPc180JQ
QpSmaQnyoYFsctX205YsTDMVJAeLdW9ErN1/bWp2poD6yh16dwCU2ajXfiisU8X1
3QZeWIvzQfoLAMPQLuxy6n9I+e7ejBDoCmk1tKjzcTlvyyENqNejfdcWt/Qy2DWg
uFSJ3NJs///igno/ySempcai86dYoX81DXXj+PCLIFGw8qf4k9QMJEV8zLkphG54
SJIxDLBY9d4Ef1P4b6Bc/MK708ORezmNi8Nw8XrDEr6X8wo3Emm1gEykBdzdqbhg
gtvOdu+4nqZUUjbm/+OBqLzB0Trq0hT43dxVA2d4axQ2XznwRu8IkiggmfgVJRuO
csEmriWMX2vU/BMeb2RRMn0GrbWlar4fZuY14gh3DvCaJFh2HdYh0G0osb24/x+W
ls4/es4PI/GHH8kgPr2fLRePkdMYEuKDXWH97+SEEeItbkGSZdoO4qS/2J59LwKE
Fqw8fgKZH/OBeLFZqBDmom8NtrD/DtaZ/hpFz7zin2i3cz/acYWwx7KtA04lY4AW
jEfpKfOYOIoPnHCm8EjA6F4EJAho/CUUPxTOYsZMDrn7cjgqMovfacDdAT8d6jXI
Bkt/rYi1sq+H65HUHVL12SJCX/54AV8a/bFwIBxxlla0D9+G6+cS1jbkHotVFafm
EegGKzNejyS2V9J/QvxQ5hTKIv9xZkM9HfdUUlmCGnr/KNCEtPsoW37ZncViywac
gIN94KwFyKI48Ff8Z4qMBvJv9kRtvLWQDKVXsBYfdFnle7m6tJzhTcC+dc0UJ/Wa
1xcB1V1QTZfCCkzhULonpvvdlWOTs5llj/ccWo9ZoCNyfL/c68yuKJgx/6KKZ+7X
3cyOYR5P1s+viayMv5XDWvOvbocJZbAoNft94O+trpvBldNaruouA7DUTbLztcu9
CeitunZOrr2+Go7Pri+6O57voz/ETbwdAyjIrKK2uoMnYDIu/7qNsIRhgmRGw/Ax
7F1hJs3h9wyUyB/QKnXhQESHMcOFPsXzwj7rRz9hYXOIQuOwzZCYDiaQSM3qzE8B
pIsmXp1giatf8oeWaBwI/sO5t2S4uMJJTFauWV1MgSwOtjJ0j6d3N2dvlFX1rNBL
vRDuR/YmyPnCU33O6aOXFnB9pcr4Xjz5GmOSgThnV4dHpk+ETuDMFUXROhj/I/kW
AZRdTMxCYKzVEZQhwVwSyh7XTG2UCLtHum3C/IGY0Cs0zyx19CPH/nLFA72vDefk
X1lknR0OyTSV8DiNyUw1F1gvTe/zj9sPy99Jkw6slZG1U/3eSf4CXUMmpc1gNadm
tYRbYieHiE5Pl5NCvxvZWOJ8TuRLCXioGhLvHpi4grdzYaaoevM4TUVp9SiZ3lFk
5GktCJ8rCewVptXRPj36Bg5EJ9SgHMwBkbYxMR7cYuIgFFFIwmCGvhvio2l6GszE
J7rRXBC5tDZTw8kjrVRHP/FegUVhg2CQPCK3ED2eosqQa0UgDKqlRlDCjZmeH8Mg
W+ReeC4LBkieBrxQT7nJP360sfL3sDKmstp3XIC9MqOc8jnJfLXtkNWqubAXlwon
XA9VuBOJAkVmM5tlNVURbT+P7to8k6WlwuX1riYh46NzYC7SPUGGMD6OL8Vu161r
Mrio4dy1cez/41OjJGOOgmZNGHv1lOPxVJQPb7OkebNmELL1lD4NHXA3KrF2q0Kj
y2kMlJAvcmGl2OyegPY8W4DGOIFeH/Loi1HKZR3cXe9e8rnCXSPXpvYNFNWwRK7c
gdS5AsxN9NGrC4eovV4ZGcyjrvg++ae4h98tN37ZCqBj14sv3gbGl0MHKbvFxLDm
qeEb39sqyXWDFTaxgmKri5jPisp/Wqx3uzy5V+m8FMMwvY5y5EUmC5ikrpP+QhXu
xTbbH6Mf9pRb+Yk8rJgqHohFZnQho1h6PeO64FtqenXfeiIc6u2oIiqGxEqbyzPC
5Y4QH99ZgRU+kMuNC3lEPw2XMDevKW+NAtGdqaXtQbyQwBAnpRu2M/HhQytP29dv
Mhn+fY6L7abBE0cGBNiSVGg0lNivwxsiAZ0J6ErrsQTwH6hmWLu636La3y8IZ3E1
LQozdeg0woFGYk1dTrxbTAHmNxVsxdBFjzBD63kRhX4DYutv5bJZb5KXC08a+6Ib
x3BvcFT36ZeKnwF5IeTLtQiVBIBGFfrVA2WUgPemw4U1qVN8rAiPTHGkQo/wspLx
hgTwARNMCv5CF/ffVdulC3wLDKxig4Z06VRGuNyBl1lUkTn/Eb3FV1A3FKtDL1Bs
ODscWkE145nWMbkwknL20YuPBpU6OEo5VbptDXDMEnSNbWCxqCvuXkS3si4tsGg0
WMYg/G0/GdeC2SpxrRb6XjFqsqa22hxAYn7b0S4gbfqeMyVbwwlh6FNUNTXFZElm
trg7vdJ1qTuiGvxgbQqCXiE7KdRT1FDf3FhAalMFKq/oyjPEuGUyMoEDLJmFTw3C
fb2ZhKo5d+GOx34n917R5uf4rQOY49DYdRIhoLCPIm2WoGMFC8d13rhT1I+p/2Gn
1CMa3CS0r/WQ5FA+GhcPATOt9IghwECfpX3pYxn0rYVzSq3Su2YcQJM4zW3B/hPy
oB1EFZSbnI6K2Pd+uD06/3mTrCVSkxM5ZKjUKcPj1VGwin9p5LUoulzvzP8W8bvz
X29Lj+xKgXQStwKgzC27LJR0WTtvqOPwG/1wAA+ivi5B7sz0seOfONJQoxtqqm/F
4irDTAc1oer5bMYxNZMEu/DAF1sXNkQ9tOJgkNAYqzllh9uW7fjxovJ7yV0y9DDz
ZxPRdP7g8WbMVaegJatIgVBh/akyEIXhU6XEIgUYgj1xVxR3/e5Uvy9QbTqS3039
jTgE41506uCaErVXuhfBGX+csVGfrWoGin/VgVhb6xuKGPRDFkwPYxIqVZ6YZNhI
ji6pyt+QBefZJaQtw9V3Z0br5av/wberTuCFpB5iPUt6egnhoqxj+sMIIluY/Rbt
n92uLHHSm4nenQiiA4+swobDiwEi27Gcc5vK+mqkv1CJx3XUxN+oqHNK2UuDQ+et
E1K5orl5Qo91ieNYDc1oCMDwVhAzJuYQPscB9z/BzCHc1NCJgb2GY/VmJbMQDWV0
u/MzMV36JsaznygnKyOfyfj+LB6YZ7XHp3NtEQOWUpc8O9DFF+9HcjVOXFglK9GL
8bHw3J9kaU+PanzWHhkr85z8CrY/qFkB+f3W64tCSQTGHRrDbX7A9Tlsojr2J5c7
iPGUPPc1y+cO8uDmLL5V3yLm/8BRvL4OBW2Yk3tiTKnRXPfmffDG93MGxLgwdCbq
B6+jseP1M//Og58RXIGJfzC/dRMXV1f4eWyVAIU3U2/Ev93ggMl2JKJPA1mMjAfN
RojZ0zUagci4PLT3Loal58xgXhjSgZux6Y95hRaQ1+qPyILAyRhlBPwtmbRm30Kk
SSkNiGI6FnXi1JVnI4z5VUdPYv4te0oyP8axVaV8LwUDxsiUVrW7CBBrGDfTpUA8
H+9bcX/c7cfQdHOXfNjArm6iPpcfyKMvzg1spBfmEd8beZYQquUIf1ALWN9JqeOs
DQvvyAK0JFF9vwnZFCwzjFfN6zRUanI/+6JT7uGgbTn4OBXTe+5r/EBC+ru/En8j
RKxjhVEfSR/BpHYqTpw7fC2ibdgChMfG8WCDA1InMHzZmY+LWYn1j8/KF+O7/juk
qFr65+iktLWMDQQAPGLmKTkVDwom1q0qUwFrCQZPmemVi+q9MUDbMMZZJ+L9iAio
mcIdtjY5kZjvJlj28t+6ooyfb2LKjgdLccNeYEHTum43gm4wqzvfgYltBUDFKTB7
eYAEjREZimstO6P+xUSrOhr+kKZQJ/+q7nAAIlFQgKWzfeD1bLdPupGMEsKeA3UW
/PeYchTw//S2XNuDUOAYLGQHGKkLn0Yd9bDzXiPioVwPq42KkkEwom4yLKx9vZXt
/2YTAvVz9oLEcBwJuFcy4+BGER9wsPdGvkySxc7ZMmKGaeHLHrH45ObTjR3jIKfb
oHkcWbv28WeEd4NiZA2lIjsd312xTgeFVk/Xa5j1uSkPUK5UXHs7luup5dd7rpD4
+8avXwhJsJe8R3okeUfJmLilHAokPQOs2fOv5OYrsWWfWHAas/G91BxS35/ojN9d
QdQu1kujZkQBxf+KNIjxpLFT7UrBln+mcdA8Lzb52QuXA/jAvslA2BKfGTCdd0JA
Dv+bKMouRvQ+gTns3oTLpWXPWlVWl3Pgd7hJ6Q+/pCk+c/gudGGvgAacfNIFPDPB
QyE878h3plCpTERuVIbRQrbU3FVFsTnmWhiZu1Te9A0y2j/eiwmA9QAr6QuXi9vv
Cb8YzEDJ2Dg60GtiJhPkZchLYnM6UHCVn1lT/KjubxWWuAkrlKTI4oA62qw94/Az
eAMF5zKjZpoS0F1asjCdOLdKjxjkinXK1NzReHKnGYaxk3GvoNrnlnyQ1fFrYAP5
qL1sPFRPQuGbwX7FNtvxAMfcCbeiFtYyb3ZYhozpe2LGMtIV4ksqTGc1jMH5WmkP
k86BAIqsDgdF8mCslnJpmX2jjhWH1eguPVfEuhhznZUpfTjU/pOvlrwMYAvj8lar
Tt4crl/dgM+V/1KxG5RFK2zqQ54P21A9J2qhwVTHPzAFO5uAU/TWvPd0leKCz2xk
3frMXAzDtYCG+CNfVQQwvHwYcy3cAJvnffzOcL1Y4HXrSWcNa/7k/ZFnNbEV+jXQ
GK3an1rjOHtwO4BtlGajlMIl3GDVebUUweZoDN+sKU7UALExMJYOvrU0FsOIYMaq
PYwQg3tKytrGBAlHhDnVDmLwWDbAkuICcmGF1UYnD8AhE2EysJQiCtLzoGTa4lHV
j4Dqko15eIjOJ8xxjGam6sCtksJrVRuBZpQG5WCVIbiZazExTYGP0xg+0MEdOJJy
QnCBC9+8SkMNO3YJBtEZWV3bM1VFUfYOhDhCMP0Q8p3BlUD1zhzzOSlifQDxLS2o
9vroixC6qGJ0FEqXWJcx4Yh739G7hVmiA92I5DVBkF3FnPTWPBSDI0WQpTdztTL3
rAxjl//0bHw0KtOlxftIc2Xgo8J+bN+1084lft/nQII95l4Z4QJnpP6Eqc+XmdtK
VdQRao2mBoOjyjmEJYAPwHUEbFqr4HR7cMfntLIOcdr38gxfO654C651pSKjyPfq
PAVXC09GRn7vFjd1wyFMXgrr7OZdKqyc61sYjSRcORgUDfovImJ7HnZ52uyB4c7S
FeqzM1RxwAZF6aTAMpc5j1xWlu9ehWpiBh5eRPHDnexq9u6u+13u4ZDClfOa9zfO
RGSlSeyozSQamKtrRrjamXGtSleJG34DoF3UdGZ+XZQWz92QwzDgpwdnEiFilBA9
RIyhx2B9QfTtXQ3+tCypEbvX9Qh/YjQBMtrvplMtGfvL8xTPiHHyPeaDk4Uun0gS
P3pRu6n+a5CIshscA3ghpfgcpsEp6mlJHwCcRXLv2LxDe5SKseKYKzjiiNjiFs9Q
Pv0htUeNw/RlcclCUGoXN4xyjbYP2InbspsGZJRa8bQpkkDhZkXVCE4clS6XFnaq
sr5CuP0bAzZ0shvKNdn4O60vRTdXAkyez5t3xVSaGSUsSybl8gDRi/2S9kZxOnoD
kKP4zK6AFnLgHH4omzNR0uNGkuFdTNE5Bjn23TQLvbRIzVDyewDM5OW+JBWMzfYd
eXuPmSs8MeE1DfOWhYHtWtJHt2htUDncfJZIaLS9ncCi+FGF0StaAmD/ISiNzqS0
xlQBl+3GimNKya940qy2ap7MB+2M6j7jY0tdKkTI66nqx/lrW7I7ZWf7eboEvLvC
wocnOOf+Cwz7BbENF/XxhPb20YETK/DM9lCGjnWvgCbmZI+ipoLu6ELw8kHyVnz9
lzxL5l2ptj1EOFoEqU7AejWpnhNP7Zi2uLl7USszECowQGZHyDqbM9pS0L+cgqyC
m6UPW5NNQByQGwnlcvjp8Vz8RKmU4nYe6n8ShxfQtpfkJ8YCW40cpC4iBLJFe9w+
zlxk2yp6hV/AhsvzYW+HLFUXKkDmwljVdoBIxD11aRl7TKZa50kbZD/AGXU1awDr
GzPOxiX5prfCEJHBlkAUSS7jiTumj0+LLL/i9kYzOkJa+sz6RKxjHgYIFcud6SgT
JDMfE91P9WkkT71leSGrVRvCO/sXHEaBGuLRGMSfUQsB2AMqgVyuw0R5ti3QcVWa
XShZfuTe3ShcVGF/RBGSP3j2dxD5d9aPd00lnC9A5Qenfdd706iawsbfAWXMGrdv
Jfy6sUy1TYb5EqdtwmuaRBR7mqmJyHSkrUE/U2Me0MQK5AcM81GU+NQz9jD+YZwl
glbTQ+wjgiGtlQNz+uM2ryzIP5/CIAW63fFiMBZzTDmZLabOR7I0ZfvDi3xk24PW
N3GX9kHS2sR8OLVlIUNsa061xnc40ZnBxns5xcoaeeyDLN/Z1UzxfLFRY5cbN00t
/oQmeRl4xFgDUy0NDNv2LjLRGSYp7KAWxnwG+q2kcYp06eGJV+CHXGjARkOhNyBf
XwbhwuhBSAl3TOXywZ6U4fYmCQegVakXUR51spdpdxVTn6em/ijwbWR7MGsQ8qpv
AQ/Kx3CG//JFoPMnDOOlwGo8EcwGFbB1x1Pxix7My+K3545SpnXtj+PFQojKCzZx
yzh5+GtuZIUgm9DLDrjk4V7XbDr5HlJc21gLnukkc7DEvCKoOgCTyUvoLNBaWQ7Q
iTdDGHCVafRM3PdZvbSJf6gmr2sZmz96x2AC0Xlmsy0WAVDDkSl1NDLV/d4AhIz0
FnJgRuqFS2IAFDjNFRT2lBVJHycJLVUTT+BQ2Iwt+/p8TWGLt0ze7wyYjt6jiExl
COZ5aIuGLWy//SNJEZwPG5NCEVLq2KYNUvF/6ttkPwqEU8mvi6zbggnQl5AMC9GP
sK4vUKONyQ7O0DfAAt2V/U7wBRUMoAdF6Q0nS8lhP1JtUm0Q6tfnAEbD1//cs2LE
r++kuRHXySFcSvaBx8OedHFwihNFsM7rli7J8K76hYgxYLnWC+fIhnNgofeEnKWL
K5KQaZ581nu8BLK7MNj72eVFe1dgjXZFQrltje+cmHsszsdRJv/wv0zseT2txbcM
Jsua3Skm1e5vYZqG93kmKWxBneyJtUkotAOeVuHcXSFyv3uA7BWONSxZTci30Oai
FyRlAMR55wJPATpdLT5JTwI3xxM0q2VVAGW+FNkVyMWlEfIy3clZtujjuH6IgFho
4PB2UrHqI7LzF4B1R980sxu37am5NznAuaqtFUZqxTEilrVCSyRRKft1Z1v4/jXx
Hz6D1Ht5xoDAa46yiow9HQV54mK2DK7S4+LTKp1nWQk57j9/BS92UGDp9RruNxmm
Wcxq2K7NxHiA7zWcn6lzAy0dvJCf5CagCshM9PItQkCzFTO4WoBezs/flpLfZYQp
+P+Y8WpYgefWGjE13/GGrTK4daPtepM4THD3Rul1+C9v4GnAszj6gbHznt8WsrwP
O3krEziPioCH8EihXJMwGS1SziPSbSIKe14WOxx0XNGWa7CRfEZEAwG76szT7mfl
4vrH/HisU/nkrvPQDB2Hw1w6IhDnsVztFtMQJUgfQ7/5gE2tO7qKEvuaRWDWGD0H
oy734jd/Q6NCK+lb2DfkvBO+nVLi3jfejrl/hG+hNbpu3waS4aIcO8MQ51atPn5v
xfxcGxo1uv9oBUvdrjtSSR8N3kxRiWJbRO+CG7HgaBWgnTu+/+zrXXkSI1/WsWCk
eS6JgqpvenUyxj/g0nvQ525n7K52V9PuMPUxnokCxX7mOJ8RoBZ+0eECByf2bfqo
QRET4dfOy6ygeAs7VyjQ8k9I38OKfKPX8FlbR5yD2z08wF429II+/HBbQ4s/HlDj
gbSSeWZnwl4Moy/nLgxd6N7Ryfx6+95swwpBU9Q9G5wYiW04b0VCvglQ0p+HU0KJ
wQAr6rzLCwbcuERAfZDFNzRUzTHqi9lZ/pXQBNSptbveG2so6eWDCeAwAcHuPigx
Lnu+VFoxJvQfbFrGdfWaRZM7VmCGrxaSUFkKgjYSqVQACOW3P4OTPfiqVNcAuztc
fr8/zKPooGbNlv4JAdou3RPglyQtK4+kqzxJ3kWbJ2/R64yHXzzbhjQBmDndUIQ1
0Y43Gr/V/LnxL6VPB3RYqddvdeRvCzN2LE/k55an/41L4M5H65zssxLFnUQf/Cul
EQh8R6LkQWNR3hse12ICOUcwzwLqrjsHCC3soB9G5awFmXeiJV+hQxx/oR4FfJoW
wEC4lg9lc7nnXaJlrKl++UBD15rOo5cYupVrLJHeoxNFk9UpLynX6Gx8rF3D9p2h
6xsavOiS4a/vPFyl9/X5jPaj/XyeDe+5PjPwFbIi9pVVi0jb4hro6+Y2LnKgdfLW
86+OEEjhsPdmWus84et+gej9TpavfaCuRHEql2r8G4CSZQhHD4RPOXnI5QHf5OxE
fvbMxcVAV4bDJtYaWhSar6TlW8KnRLdQjd86MJw8rJjDoTnTI9+KAQ+sHX/Xn/8c
ZSPtjvpwVa/U8zKSWho+oIL+V3axfuKumo+AMtD8zk/Gy6J6ox09suDCmGfN2gGJ
t5Br/OwmR9LcA92qOcSklY8lJvbkMGlt1Ol5Oj3Vwr6rQZ9i0VTmHQuOlI9VazGP
RigBQmQtLKtFYTRU74RulZYEGyzV+q9v6updm0gfd11tvnZCvnObHjcRV4yCYkdm
CktH1x+CGI4GI8ZxY30OctXuUtelmWllaQGCPD3uxOGq2qYdVVTdrmpqdocryrir
uA5o39CbAauZ5bb0tN0C3bItt3caI/RF1Wo5TH2dvk0CwORfIMDgJcFEfsQvCKS3
SLqMq6HGgDYBNap7zh5Lm3ZvHqGmQiTttMV1LbFieZ7IoXSpGl5wOwEw21sCE4J3
amKZL6dx59auJ8JhRVMzz5/lWwXaoRIFe8t006tdFvubbSFVPL41i3ZuU6Hjum7d
9koMVr4EzrIS21FsvCV7txjkqqyODF31vm1Ad3xDa7Kcz8PoZE+RHsPifiLzA0Wh
ShuyiOJYk18BV1sxL5PH4JgF8hWvVRXZGo/JkRnXIi9KUCmvDWRj9Kh8YeVqagXw
55RZ8y2X8exWerOmAwr5SDJIz4it5VOWojjIq7uQKamVcQ0lAt575xV6NukBDPQx
IDRlPQ6AuPAIrfKCeV3ZHigxn+nFKWZmHQ/CjKeJM8xm5orOz5h+j0QVCNZH3rR0
DMQ9dbNRaPtbzCuxab/apvyQl5113IvvIimijolzqI3nz79sPvLoz+b6zIwqXGHB
KyaReia/XJJY3rQpWEutDT8C/TKw0f8gnqKBqSqGcMJzSJ4BadI14DEx86Kdf/J+
K8j7NAQ6lihyFsYRjyIGbpbazhvTJ8g/KOSMEkxb6qJ6NRsIIyJdh3SXMEIsmorn
sg/2YFAogyT0ZSuN1UIJmABIXlxLmgYlFUsxsJ37GCzorGEh5XK+1EZi5gjp4PVL
Mt6nTqohisTTDbpZFHJvIKE0Kp3JHRWX/lIpncLK4rU6N7gZuSwbdzdIE45zUdG3
pI/go6wgNd+0H+EJouoZ9KlkG/zmKgwCHCZiqvNbaw8HbiNojpNHhUb5nX1ZJmXI
/j3eV8lBXu2eP1S3IZnMc3T/H/mSVbA3s9msbcdRTjz1X1jXk0tCWM4fBnFZiFRF
x1N/73KFIhRIl51HQhWatrQwt0fzn0ii9utRe/1tw0YScQUKYw11zqyyEI/WXxD7
pI8km+KjHC/jvStr5k1Mto26S+pA7V2QTTD1bXznSDvCGJ794VcnjJYkJ0NHEl54
sAfriivDPKcoifYtbo4DIZLMJ9HawivfpAHqBWna/Iqy1f72S9gWM76Ai1SrwlwF
jMi6K/jYowjQn16ECkBaOJ7UkVwsvIF3jz4YSt4kUGxHTS3H+cclFqg1JDd375nf
x1gjt1WsoSpelxZCY4JfrdpYJlzhQkSup3wcRo/cB4gJ97qozf+Wpb7aXV9FH/+r
tLQeklVAwTWPCEDAiZDr+Nw7A5cX45br6oU1lmrBDI+9bdm4GBrQti15KPTn8CpS
117sdUuKKhkaPscSeSb4qMbcSWTP72gcwXFb4OlGgiq7htPeIqYtdoNnoSt4pZbP
RK7Qz9p9uSdeVMdsQUWBgMe/CY5m/Ghv75Rn2FK2JMSeawjK7kYmlJf7spU0l/xx
CN1Iv3BIABCW4TijMggIdypu7p7Y2/LcOOaPzXXfvXL/F19oDB5tyzxEOvyaReY/
z6v56TQw58DU7ca2rJ4EZ2uIHLrf3djUbHRzamyxHYRSRu2v6rJ/gd1plv55tByK
QbnFaslVm4pN5mGIbJ6oXw5U+fjkqmO4686m3nzy/Uf/4tqzhexS7/Y5QfoxATbe
d7WIIT4d7gicFEkgzuWQRzoEqRl1eRQcIa8y7jEWJG+ej+Wzwwc3bzn+jXwlE8MS
lSbFL1qCzNt1LXmyaAEDoazQPHV58d3ilaZcGHZm1PRwGW6MRzDTcSOqt6vQuazU
72b6ku7KttF0JsL7cSltb1yeVbgJIZcCoMfn3rG82/E8c18bNO8kKTUF2AF9n1Sx
cc/EOGBM9aduKQ52BamTSi/dp/y6v44o/L8t3v37p9GZnt/ukOrDtmvhrEtjeY46
rsUG4stwv3hJZl+79b6MZ0C60GPMrNtFP0gnOXBVAX5X2t4uDMDO2DbbMdqR3JxL
x153wSURbiu9MjtB7KlgdHOozO8WtzPfuMEJQWC1TMMqckaSuHK80b+/Hf9EiHLp
uXjhNAdn+bMEjhgkBC/SGvc1jvlTYt/UbHOefug8nBicGzYbCRAZofzJyLLfS/pd
yLbih5TJHIyfTKE5woGqixKD6l8Vkpypk/v0x5HZlM34aak0pSv3iL3Osbvc30cw
jStc0BGbXw6yCjzCNpD7RwMHlAWdg/bUvFXwfX5Vo5f1PeFp3Gs2437g9eqadOhD
8W/oTV0t0qsm0DyL7oOIB2CVJd9OeGJOtGT0qMaL3GV2uSBQthAzclhMqFyanvOZ
4ucmvIp7ZVGaadqoCydYmFIdkhn9MM3DSi/PKq8KDyXAt3COk1puC8zRY34ohF07
I6gSJCMLWHdwxKM4raQOBbNuRzBYdaNOlrvSH80hB0h8bz9HzjU3N4hwi78FiWOS
ilcAtxtEPCfX9ffLD7jCSq3Kk3IPoxftysA82p4CcmHinsH1OgtPEgW/eR1LiqwP
9SBHQ+ZSV1HbhCI5N8gSdfa/C4Q3Agun3ZhpIEhPkiyU4XgmtVmaOXyTPsWO6ykA
IMA/oDGajg7yLTBhjk96Tk0XSF4SpMIC2680zE5euPXZMIXMhfDGIx0THyQo0vqi
EWY3kOAdr0s49jdP50736QtAeH1TJLAHF+e8PBia117wcGYjWpFZTQ8TKaiEeZue
8Jqa6dENiLxaNFajVasUJ83fv2/xwjj5vOkgmiF3x7wHwT19FPd2i5DAXkUo19QJ
2plWln0cDdblspij4BROVLVmXrtUAEW8+OPH3PEDI6mJ8C+URpvU2G1IzdX7+Xo/
aaiK3PNInN0137/TnaSb5oQFvfN7+Y+QZteIVv4X43W8oijHPnTnCpBsA8tRxoSi
yn9Igmg2UEG1f5JDolZX44/QGZn1f70HGmMbQNcLUJyQLX11yLQkqq8trUaMcMqR
X1Xt7YnPQkkrTZErPQYaaFXIk7iEvLmLyiAr1hN3Q/NCM9ZZfTwGFCC7NFBPv40S
aWjMX5egVW7+xMDnMUNg52BOIxBg2oJ7fCQERYpGsgI5Ya93KM0ruyWakIU48Sot
yXoi13Sa4R+gUN2CVRNfCHq7f3K9BfpqqQDH49a87NvGebRi2MbH8YeWbxxhJNj/
Jcxnq6mCUAo+RQnf3X8/mhWGkjeqMG5r+2XVSorllr5DD4sALTAmB2JgTHvHN1So
EuZjOIrL9yJGWKOwUsnh7w4EUm83uyDqmpyVWn1tS0R8n2mxW8ftBoNwq2UbZWbz
4KVKcAi63MiJlk0Z0/cjB6lUzyyRQFtFKMOc9t87YdEL1ouocd/tk9bEw7THI/iy
d2ym5wbFrA2V9HLBAxKvZ9JJ0qgel7sCggGOnbZlMnuRui6Dyp731TMFIk+IkNKh
YRBdQjh0ylJGGuE0LRcuxgIw0ZZ17967wCte/299H06aV7+hyjlCrg1HalpbrRnw
iXWQEeEfsJORcoPVHVLs9LJx2/V7a7bzyEgioIEJdZ8597bauleYiY+FxdNF7H1M
TnxSZa2D+Pq5Vn/Co3bQOxGCOXQ+/CnShwRjm3tBw/oCOwgM1ciEZgcn4rydE5uI
p/SBiX3KYs+4w7NeFx6QgNHZn+FdQHQtRJLc7Xzxa+Q9Qay1VVhIheYp6ZrMyxqO
kWX/NtISMgD+0PoliGMEBPoTmWkkFMqN3R5W2MKjjFLHq3CL0+zW5wQ6rVF7pBpe
pPI2xCxrFocypXIqs/YPu/L5cC2/QRfuU1Uf3P5/7JmYzOOXGaHaOGPdHn26yHrC
+dWcK+lrljqBF9PNKxNJpgGBkzLCLF9oRJb1Ek/ZfhVdbQsLpGbZf1pniZQ6esXK
ub8krHnBWWOYLYUL6u3uQo3U4Fr+AFQLG3Z9ORs2Gb0gMFg3QOLDyzGcRuN+WcBX
WayqNcMvq/ayADcokZmOIjN9J/9Q+SM1QjhD7x62xL6vc1YfSRfmtAtgVW+0RRWP
QTtHQ1pmg2BvnvKcD8WEH94wITsvBIGa7/ulnwYU8CwhqwZ8N+G8puAoQ50EFiqj
eaOajgfxjBalWwQmZ28Avd1AMQlCMoX2ZU7qWde1od3a1VXKkjL23s/ql4Fp7GcR
8aqSI1H5G//5g/ct/QN3D4b2R4g3Gk6MTmhYYn+LVBJwCXRipz/bFbujcDegC695
ej6a7WgjDOQMwRY1WKWS8zfK8qqqdYpLfhy7ROSKo3/nYQiQ3CmvGXti5J0bLYaP
NQcCq6at2nKHBIdurOpV2YyxILp61eqMzerppgicHxr+VuStXvJ/9PnzCaBZ+COw
7HOgENHyNtKh/s4Ik9Y8+HMx6b5UBWA6sXvo5cNBm2JCVV/aH1d1sdRAqQLgStWG
7mQxk5GATrTTKuOHPcrBXsynQufBkrz5IGjc9rRhOn5F0AqDyWEIBDrvAjJLIPns
ZRmTnI5TWquhItXGBzxUXNsRangOfLhI4YEe4ZvMF6PdvzJlLK5GPPcMVcK6LG5R
8OUCR8pJiHjcxVDARWOYYD6n7e7aSEMM+3HtstFQjWIoRGiOVMGEhKkXl6Rn6Cbr
0AJiZqZioegUBWU+NzClM61s5+Ish49BW0Qi0OHWOPkia3o1NYv6C9INQjG8OtPC
xWAK9rpzO3lsFonlEMA37yUQ7mXiKDlooZLthvJRuy/OE79M5hSQJgJsM6UESy8g
Cdk8G90gE52IMCiKZTKtzoLu0DDh4mFRSuW612NaweouOntnUVaeOpwvkE9L+ngU
iIDrI6NR6MlqSPpL+Wi/oixX9gkETIIK960zXwZ/2q4prtRU83NSs337Svnl50i3
O3ra1MctGui8WYK6RPSz8X0sOg4ZfvF0CuFi2m6gIuhLJnXk9a6DypxXH59QFnVt
hbj8zQ6LwRL1gOdnxAlgIhrswyFvwW8nnFxy/IIQLMAV5ER3CSvvRVc4wwxjKPv8
uvs3D4lsOlU2OKa1y9dLNn9QoE5nZ2eV9jzUdVd/HInEeMDw1gk+mQHy/eBNAGCH
5zXLqtcqlRJajAXhiwyyEzWzM6dQGZ21wSyu0oZeE9bv/fMpsPrAfM15oaLNL0e3
iDwF931xGJ2dTZVE6OPgte+KEE6YJXaudzlqRcPdEBa/AkZ4sITYGnyfNhRumeiv
u7EpxVx7U5YmmW9m5WYhTZJ5weEaqtzBpzL7Bm3L/Ahc6lw5nRSYttLHC1PgtzcX
Mwc+WU65wyXnu1bE2AsbBcDRayZUoqkRSnv/PZwYYcT0at+SjV1mqWDaFwVnAqOD
7JZZrhNb0HLVC7z2h2umjtJfKVmD8LWkXYXG5FRIOQ9Q89AuLWklVGYaLTrfeJT8
RfYnUDZqZ3teFyRiPDofLQ4errdE6PCcmWaChrYwuT+6g0vWKX5IMzv7TTn3PYCr
nP8ZADd3nDAkd0K/aJ1NbEBR5bR/iopzvrpv8B0Gzigr25+Wnf4EtsVjmbiL2erd
wr0GfYYrYsJum9UY5/Kfr825I8jIYs+s+rdvB216paeZ0kpF53zJpL2vWHDi1QgL
XMwydhyIsmabDtF/q5z9ifvWwjcw9z+2eHaP/zkPhBMMNf9iqegyaMgJOr3yIk5D
kzVCBGEsZEO/b+AM1eKTDghcOZs2DOPzWv1V+XBDz5fwZXY+qhTqBWz7zCmYfOZO
R1QXKgm2XGHwwOQnr845eyrQuZqA0V1TiRDCQmbfLDDIMykEYGdzoHmhBQQ5dgkQ
RqbQ/x3LC8/yxZmXALjijrV55GnNzHLRlSG7KaPxm6xMBf3YYczC9VLdswfRv/5h
hd0pRGiyuj55pPyY2kdhTjhO896wHc8SX4Zlzk2FtNbdcdm0yQAwws/B08utGVzH
I90jlOkffH9pyOdiiAyPF3dmpmXF3MSCCSPFc8BKFT9z6Q9PNTQOc3828AGM3DCN
SaDNFZAd+xUGBVsJuLkACiflVlw43JacNY4EVVYlV3CQ5voTdM0Dn4zLWKfLP7AQ
VAdxM6r5/7y+Ao12hrw1ZpS6CcU6f47K4s4QIGkEIvY85UQm+THzKceZrEr0jfb8
byGKN5UErRU51czn3Qz9myS0LqHtbzvGJMIqUuWm7h8XpG5OOxXfK4iNnjF3L9rk
QRGhmTEx05Kw9cDLRr5kww2lSVCvKEYgDXsObQzsD8x6wgdICzF1RiWQs8vdhvCV
0RHaF/CvM8cTc10CiyH8BejjvpE/5TcYOJ77uGgyQ2t+48c41xxHlLfnfAqS8qSV
pJWQlzxhpUXOgfXD8qq9Rq8ojYuHU3BBZrkDFl9pV+3TVBjS8OeI1OEBqnhPWvBF
izHDoovtdWbeNiG/gaMt3XQisYJ2j+NmOg6HbUrWBLLl5DK5jalA+4L7L+6+bCCj
LQ8RV22vGQmahXOrLqCv5HmwahjzilqrACefytuMi9E71xAJbU3/lMnqEMy66JGi
CbTgQIXpWBvxA5+wb2HznN9nNK3fDQKTuFnzEn9rrFh6AozL9hevSxpclctfOa9p
LuhGO28izYR9R6wfzQMQgHHRgjV4g1e4UVg8QjfveTKZnhF8pNV9YquhK40WzJEM
EiC2yJ3HxYYZ47zvipjG1E2klkGeB0jahcfrnwTk38SwmrPH7ug2f7EbDv1xEY8/
GTfrlmRqNSSKkUZFnhuywT+FJJUwvq5p5o+b+UI5p0x+eu5rRGRGqw2h5qx9f4Dy
quK6kQv37tL9oF9a0g+8D6xY74s5sy4PL2nEmu2fOxgVc+4fLpUxrfilCjqApHDD
ow5w+odHZ/5S5h3n0vs2tWe+XdtBlK4FJi8zGBHB+xO9j423NS5y9Smg4VJsE80P
SYJawl2Knw/vVGMr5PylE1ER7JpYIIFIPPPWKM34cCKJsWoseskBI5NddeaxAALp
gkmYSQvZ/uO8hE12PqKC+PNMj69ObmN4aJJVywBnt7fFKb07Nm1yOFfL3SC0Wx8z
PUYhtI6HVwHyiDT/UBCcjj3go5++ptVkTtgTSQG/5I5mqJnpfmqyKvAqryTlZDbu
y1dTB0nhTOaeoLGW9mCzNUJcPq5vIrFT5oTiVicqqyvBy0fRPxcvMDhWAWDce0e7
vabOFY1AJ2XEuxoJyEqBRxbea9BzBiturso868fwQjZcAjxzsttDYsIIAOJmuz4K
083lxjHw/bSAFM/gFFI2csY/AEe5TsqPPWBTTIgbN0DPyM8p/wuEEvYYF5uJQOGx
+EZtwJzPYu2xyGFVzOIPC4DMfM9q46Br4qcVN4FT4Fd1lTSEcXktFgxWScwCCtIP
109HL4IJUhX/iDwdWDv9v8q4IuSwm6Mk72GUhetu1XeWPjSb/4mTzDhQEZvFR2yW
QBe79KrhKWtX7krG+sV/TDLDdKLEIB1/Fn1H4MUuWxxSvUIPoIsNghjYvG74azUz
+OqZwuTqoCH5XJrjyHv0rOVraxRtx0H5BVrvRdJwNGekARak0k6jm+vdXSlGoAM+
9+aFfjQbHDBn0Inb8teW/a7sLd8gikU77vLytVAaEhuqyGVentm16+JDL/XTAJYU
jzHWk6rHOnWp/fxl3z/5VE4C/byLXkdP+lqw2JnpyG/z2mZXH+Gh/lS0GTusQ6VN
OPQJbOXuyDq/UL4gO+Tkz6WL+41QHpk0GRLFH3vKMmoHy9ac1O9xAownzLC77gF7
tmyDwwYPDPhhxCmHuhk7swgbulIUCtqTpT52Y6f+NhmGYqJoNEy6Q1ejFlGR5s/7
QbIQ7HdESXkjzw7/A7LhsJ77MuANQ1ZpEyCJ5WgO9gY4214eHfzogXQAKniZpC60
Zm7eKj2YqejdiWBBzQlN6O+DqHamnbnLizOSiNeReAtaKvfLkNSHSotRLqhwYpCO
jRsO7roD9TGUglst3o2Yi1S7eQb9eYSZ2FOkdVRNarDVU0AQFwE5BtVLKLl1Vdwk
qaZvH+PtFaQTBWYRFbLNCUzB/HAfJL8EcUzXMXupYnlpRMZzbCpj3RzpHZ0rEAEa
LKgMh/cIhAcipV3mLqZ/IAljqZpovIvKofWVl7bxY3NOsDgBMPOchNFLcsE7Qbcp
wU3IYQpy3ulcrME3w0eAfMc8ML5b/RNDcshtJgkqZY4qOxmon3rwMeb0C1BPp7zZ
SHzNRZXCeZBPxw+xOFq5/sDhfK18O12c/M7xqKczXP9Ai3KLsW4T9BJ/VOHiNinB
6eWwU13Vj1uFuAzw/mZwGSP+QTlRZarOUhNoQd7geX29XcE62SG4s50foxJ/Yiy+
YVzpNWz5dAp7AFV/TErgUPCfTAPXXx6CBFqzRf7OAMhzWU2n52kZbYZzycZ11rT0
5XYDefoJdo0kNvTw5zujOBFqrHVWXI43qlsXcOkgHYK/Pw/m2+NGYQBVxUWFkoue
DaT5dZh4KBVcK4UFNFQkFAAh+IUTOaOiQanmNunBhuwhnxU7JXC/DzvCy2JU8lj8
lkY/qMVuTRil5Ny2pqEN5NIa637uYSjkLD2svWD9waMFJh/ocsOn9BZiS26YjGyA
iS4tTai7mt9AJV4QqLTpnhu+G2kQXJaC13Y06Dgpm8yWN5vjPU+kji9Nkg4mc5GV
iusFLk8L7RH0Ct/PzZ60cuAyyN7gHoNhdhrpSeC4dtqY27f2FQ8T0HQyY1Ivx6wL
+BV9sJn21NtqYypbN2PajLRFgk5nPY5Fu/qsIzWkqECnrhWxXImZu4i3JgrGB96x
FV/f4DodE6bamh/kzLHERZFKCP+Ih1JBzz+IP6IdYm+AWMNWbSks7jEfvsxxQkk0
BI4Ducwp44DyYJtWg7eX7bsZJZ9m9CSsVLpJUkm9ct5giE1155oDwF+ih0ZH+vlM
lrgMQmOWa7dk0kMidrgEnJp+xxMvJRetN4rX20Vmqx7q/IJzNqOKoty+LvyCmu/h
vUTvzVPQznCb9C6R9Fe8ZiEOaXEOIDk+pQGqHWwujpVUJa0JN02QXMMKNu7VcWvC
YRBogMmD0jM0rwT8RBCkCSzhbDM190GnDahOd6tVrxP+JB2KoC8QGc4AIjsyh6w9
fbRFO3WKsk6m/87zdLaCGRuFGIra0+UGDkRECyt/5mxRfZoNpHHkdIzCNWnH9XqQ
CU0pJY9kerWPLJUO+hvYOcPngoo2W3G/Y68GmwZ1o1oxc+grrfhnZ5lzgX8fu/2I
OPazDUzZO8GSd0gj1JTr4G6b7TUwdIWfRQxnbPgrpP6N87asjSP1Lq4mEOZYFR4R
6LbcnLb6YuVVC+o5ZkI5ngk3VBhoili7CsVQEw9y+JZHlENe6X47zXDerFWOJqmi
SN8TmhLk6ozjUNm7cOmiYd9WuogAf5cfnmPf/csuU2gm00f8h6YrzJwj3Hs/yH4f
n28jqow7Jddn2SKo+L+YFuVH2L7e9Dxkvv0ZY5Iu5zDWQpaoJenG+xST3VDk+0ap
P+5UW8+H/jBWutWOa6aI6I5vzuUO7jF2YMcQ85fKAwMYwxjYx+UcK8YxF3V8YRCC
LMRn4CVyBRO8tMTIFTOQd0QQmU+04RysRqF9tSIh0CAOEjsd3y6z7K2v/3jTiflQ
UiZr05+XdjRR5oqxaRSfBUu8v2FMr6sB33lqTkKE7+ojssVh49sW1vPFAUt+9z5e
tS/PttLouWuTE3lm9D8jYW3UeIHkkaJf3slOFUmLiQ8ahb42Y1IC0KuPK/uPGOL9
dZVGxLpXBnh/SPMCsiWxfB2rVwGkCvqm2DjxvLB0wxTroRgIwe5rRMkALg7BKAlz
09QVQY3eoIafTjAYHIjHJb52mGhI8S9uw6XfTB1gaa9foBNtijoy0gSy6tXc888X
yYFmumdYAfuSmy4gnCIg2fB9+Tt/LOm/xc0kbQta6I49pJtmkmlydJUOw6Ug2Cem
JCdh5XvxZEjL6dmt2uv4Ix60qwuGi+MI6VYv804AwvBUOzW6zSrFVcQq1IldAENk
IRfyOeRmoBy2j7lgNv98dghWxpiOwdZSLyv7hmzX7v5H5mcfUQlZwgC/Qx1LTUB0
mUU4NO7ne8kkA+5VLu7KerxdkZR5gSQ0V08UqmfBxss1Lxp5p6BzbS7dP8RO9zq0
nJnbZArSBHwO9KcV/LmQLhaGSs1oz/JWQDvwHzs9GTEqJobEMROL/LxBgzHngyVX
yORGN55Ze+OUuEbIGzeuQ6Jbf/oWjWTZajwtLzK0pRqIah57nlR3w3Uy+nQW7JpY
tToRDU3UAM+r93doUkkF0d8wrGMyI0pLTkZmSJq/6CBo3a7rx9/7Z2qh+Y79QFoW
+/sRzhU2FxcxWc2X3cP3sRIrDg3fK6/XmEjKOvuhD+xP4rmVFYtjmFtGAZFzu/ot
syGe7ziRIEd1NKwQfhfuL+gd9ITabzZqcNORJrA1t3+CB0NBhtkIsMRI4As1KQks
TqgI+SaSg3+DO0V6YWX5HMatriSNX5ywBghmkwGy9gFZTnryk5bjJaa53UudR21+
1tulH4EV/jTxxzmXFPf5LZ0FID48DgmsqwZMRSGt7eYIqLW90Pwt2/+lKJua8+si
gZA/bA22KA6NQlCbBVHJqrbBbHcd8/r2TXApkAPOTNIRM99wTgM6kPY2Z/CPrekR
SGyK91GTN+7kSuLaKMPsKkD0USGsbouvzLnbM2axakQfJU3rD6nacRiohhclUUZX
bDQUk69qdtjz4IuDrL1ifSRDe/8Bjhf1Qyd5O7jb8cRiQIRQ5bemMfy8A1HmYU60
aWtmR0Qb41QPjZHy8ILwxVlyJdnhz2yeLWAQvjQFdo3Q3kuQBYU5tzEPaEjezLwY
faSNBZwEgL1Z2ZkxTB6eHR2lmkPRuAMayk16/wgcYEw+2vfgqqlti4m4LX7q6Thx
V+yCPtSTRF7q4b0xeOuZcDuN+sHTZ5nTd5E2sfrsgn9v+9hfYM5ytMvSJsZsxyK3
Xui9aL3VzRz1rrAsOTf1N3YsEMwjq8/25a+pvB7fyzHs5ajBtpZOm1AMyPWnNqQN
bcMe7hl+uH+jDy3NBGXA2LcTBdZV9pW8BW9uZL8RRN5Oau2N9BCMuPbRWyTd/kPr
+rLavIvQXz2DB5vTIoa+C+7UmX8av0aco9g8jjq9dU3koQI8CVysDDT49bdHUhP4
FTstsRzGdgnoCUhaMaiGM3Ht0fZT7JVR5n+g6AMO7giyZwheSF3zdQdYvZpRNv2z
HH67P0bWX92WxyvZBGRN1rwGs5TegKw8AvjYS74TzrSUgdpBjy1JhfDwqxHFVEKM
aroqksjmuNas76GNK4et2z5mrqFA9EuzTGZH3a2z4yrcHI6xskJGnF3w2PlrzglT
5ODfiLHJ5QahDLOYddosqzwkZbHhJTgXUtSuDjx5SxUchtcBrmStaGujzgLJ3ELW
Q+PFqFdhIlSa9xEIRZ5Wj1iEpyWC797WQG/82ec2XsWZi2GNOdHC8OUzD4iLbXRZ
emuonyNm7oZ+MZUpQzfIhZNvYpx7lSs3/Rbl6UKhN+tG/AfO7Huebo4FaOslo1DL
On4Si12cC6r9UYzCceywQr9Sj0nS0VzECVppQpC43AmaZFP+kxpStb5BRnwF0D2i
xsGIJ7AoB6D2y8AnsEuAn05skSXZiGzyz62iYlWV71jr/d3eKnPhBxL3MaC1vi0L
aqJKlHGjRfFnttw5xp1lp0s66hsXxOq3R4T5G69NywcK22Bt3gkiLqumWQp+Pe/z
wiTNEVIsZISryXWehMsv6N070bkbGTZC2iRk1GAQHBdIq7RccbqTnKxSu5xH+59g
6LX+86bviUpK09dKL5TpotE2nXBayKFc17gYqP8ApRV/OUcwSNxIb3r+6gnROLIs
MsVFTMSXEQUgAJrRr7eS6cvh3StCWTM6L9JsfpPkvAqrxT8E3IkhxaLl1lap0j21
P8EVe2mhCkQ3z1Ql3QSfUMzZp9hXkGusp7Qqp3YbMmGImIOmk8cniRNKvNuiRQOZ
0NLmPLM+RA7oGeWw06328+rI4eplRg8pSNkduWlVOV8epfDQJLLuEZlk8cyl08Kp
qUwK3VwUqubHsPcSz5JDfuvTVO5ShX+DkWaahTML8+CZp+e4vIPkCuNeNVzCcL9g
5mAUAjeP4nvUIfAh/c3FeMHCkN46GZf9nxrtS1Nf6Im3djM4r09CKQfFW7WUJKHo
iNPbLp0iSjuOjDwLuLq6Vo1PpXAZ/FItORkvF3gmlxe5jYxgK5Fbs+JI1f/mvdlq
E6rNSilQRkp3E6EKR0aHcWCVL5ozxQ/gWe5bkCpw9XD7MwrhA/7gY5mwx2rmebaX
ppFxM4tTIdwIYZ2970aqW2i8UsOOmr+rn9KyuQGZnIlduznpGGMLHVu1t8jFZalT
cM/TI9aJUg2b9MVDaW/Mj5KWFttmRtdknXNFv0HdOOI6uOXdPhBV0wCcazCnWc/r
qpmd4xzLYxxCdX9TedYRdv90pBtB7hMbKN4/MO1qqVa2hEiHCmEaG9TjL5k40VPh
kjjHGjDdoi/iwAjEmkjx46IarMam0KrdPg9UnumcPV6GyNbQs9UVbTB0rtQ0cqkw
yiRSY3ez3GekBjFm3uC1H+t7hMl5cw3nftki5WVERIpdADkoi7GOGtkAx9Op4AdQ
wNmIrCd0LX0j9EL/+CDynTcDqsS0o4VPGrKQqlIo7lRkZM1wV4wrnQuZh1zaDNLD
i2yKQz2CuulPM+ljIaRxzCt8OAdJjqUhH5dotqBD05pLNH6qWfpObB53sDbUvy+Q
RU+3wsSxg5Heiqjz/K4pI1HVCz/M604CFBX81HemdGl/+cfwMMMIi/BHyVal5vs6
0tVFy/aeJ14mtUse91qNNztofAo+Tus9aqXvQ9yJRiHJmc2xD5KwT0xrBDbEMgM+
QfoJrF7XrNuL8dnV3QLh0Zv06O6xOR16cB3TRHyuhnWaNTUxkYJ5cNGm5jeeNfHd
e7KTLjkfWXe81jSNwQ3Xog72d95TTeb2zapMC6Pq6DktIlN6Vuo6YsVkSRQGfQcj
EGbhp9xmhCnXRW3olvOmimgCT250e4g6yVbFHTg7VFhqvg155eKr2WhBdTR+Sx39
Ig9lhK9fBZp4Vqo1OwAWK4PquJ/CF94cv9izEgQ9X6u65FIJ5vsGrXK08LFDFDYp
LdowvqGfJ4Wh+CPt9D40wHTaQhHKeqp80sok/ZtG9o69r4JCG1RiTT5WhNMNoAgm
Lk+MkYqTKIdBQdRokH/KwdcnJJOkFriJSJcz/F+NtzP8MOFFPJz+8vwm+fn+QWeJ
TXIfc7MNrUSllK6ybZ06weaI/gz2JYtgV0mD0GkxU989xR3hpGdOCA8LpfEFFu4k
hmOKDKkRblE0tT3CQ612whniaNoox+p9Ww4ysCuxjoCkv+N5eqVCIjGWzIkBULcN
7ffm92O+tfwHsgT63L+uHyPfVeZD0fHJvyHOighTiOl4bvJOYOmaSLDO5df/mE+5
/Ew9vNUx4boc/GsY0IDRN1AhWFq6NNhzfLkFOyViLpKAn6pbxuKxQGKMBq3qg2iw
kVRCKAQS2GSXV0zQoVmu+pgBl/KUia+8XKnpbtzFK8dr78AucgYbMZ/rK9+v65bK
RO17iD1dKaw+T1ZiI2+OJ369SduBT/rTC53Bjr7GPR15J2A64U5P8O6Jezx0znvp
eO89wawxi7KZW6VmnqconZgW1YutIQWL0vDxULz0s5eqjF0T7YUV9Z6BKnMtUa4u
6k86A36S9Ub/nthbuAz5gRrvQicdKym92gYtuIcPg43Adn1Yau+RsCcxkvKK7Z7R
Gkq7nSas9cM0hlnUa9+H8mZTB4JDL6D5Ui4PRnYo2MnbUDHDpw/7ygwYBApszJ7I
Rrw+u9xXwM+7iYzRaWbsjaN60dk1HMyVVh7pKYHO2tTwK17luCOYUjhdgyGgWbsj
Y3F91KD7q4D0sKG7jixOWDdZDhtKuUzdNK3gw99hIDXrbc1SqKLmjgnaPxmsKFUY
KmCEmUOQBKMXHw2uw2G9fkUfwDfYbdfu8OBRNweV94lE6yriK2dausY5KY0zV8MG
jIScYF00CQnIm4CvAtQonWMgmx/fH3F9f4q3VNvwgtMdZ30PJvbNMz1DrKcZrnHR
lqzczsqPssWx3A5CCax5N+s0wxFXByuRmH7fZP69kOn12xw1YJzCdlIbvqWyYi3Z
Zw4Wc6+X3XOv7NT6WPJC8gAYJTU+KwleitbwEcRgTH6iHQN7wDX17AyH1I+7GTWY
mMS6XQNJPMWG6OsaXsQ51Ivs3WjqirZN3mhwqwmgAP4XP7d8k5Qa6b1MVXalBRYy
dr42CXLk/IWt4fZxRAcN+91ey4wNdcx4vCJYv1N/OzueM9kdmrTU61NHyzQ4/fmz
Zfld26brgfeUJiOX/q6qGCt3pSB9U5kRvJPMt2570VXRqCfAPU1TqHxwBCwCbWIQ
mcc8lo4n9UbzVYoOsQGh9CjHnqYhGxKMbtycAm6Wht2Y8hPeL7feXUNLYjCxtLRN
pj27S5OB2mk0lTlp8V52oU6thnfsqbFxpuEpZC4odMewXZV/jZbSXHc8k1sgLn2P
f0u2si1UU989GWVMODTUjiW1oJVY3eGehof5veDkK+gGlLGClm/45jMJfbElaZkk
f4Lv78OolI7KBAAxHB44gvFhdIVQDYKEiFm2LGahvhcpg4xw+55o6NCAcAf5UDGX
TEt6sBRju4382NPZLkguiY/li+aRcJcS+Abnlg+LeP/lArRUPFjPtFHBdXlXec7p
DoMfqy73vMKOxcZrOWxF/ocnOH8M2ESDp2zjcDwEq6fywy9ggD2OpG/FBnr50TSe
tWs7dmNYGtbjAyfnO9ODvfkiIjJVOKr3/UW5NK/ZCUeS2KruErgh0kDz/sYQ4HQ3
hHTCLpwADb+msxljbGTgphf/rOwVoVyJoG1XeJZrVwNI2oAqpqz3DlVut5BZ9vMD
zVZ1aUzJCSLcQpAQ2uDiFw7QLRbDW92iWVPKnZsgRpoiExQryX+dZuFNhDmlsrNW
dbTWawQg4rlb0yKGT49Eq5yGVOVVVSUG33zVdTmh8e5OAfw/7JAdWEvWIjA8fU0X
EL1vlN2RcHkkCmYAJWS80pdnw7GFmlz+9oPX+TcGCwlWwe9BmartYHZZJT7/Fh8K
UpF2OD9IOm9QbKElgwb+5Ns48C++0jAcTb6k/EhK1wvqrJMBwMbbpkWfKg1o6l9k
j9iteZVYTPw0CpnUsymrcWOHfV+WnQ+lB2WYcLdsOwhfzPpfOYXk58wPutgkiV7a
tjmP3qVw4ZFwW84rLFoOTkpgezoVFdwuVDhGpDiBqo2mG7WxxUUun1olDV0d3Uqt
+iGFaIxneAao57miE6bABVCCoSZ4SiExAEd3yPpV10zvgMoQcVTt0WXwmRFU62xZ
wCTk5mkXD142GcYdJRQ/DnJJ3Zw6ez1tJ+hgYj8hG2kdt2WqQreWtyxqY9iOkPfc
s8nGOXeyFA7LFCo222fCBWNeosLzt42cJ3cCWm4ejAE6yfVoduWrfvwegFny6v57
w3DRv9P7PGrlfRIMAlThbUjhhSu/phd5THb5AiPeZZT66pkNkMY9/6Ee1p156N4C
dudCXUUYo8rruE36kusP87VEmMi1XSyJqJOlM171uHpxirAGXDyZTixIm9a6Bypz
HQhmTzLM/uLbB2UMwEneK8gGCxUaqOQmH0CUbvqLuBBj0oNuGrjAhqr7WdBTQlye
plIxkQvu1R5F9c77WMd8FNucjVvHFqAydvpVEJkdNxmuyIBqn+Nnww54uL4LkX78
Kvwgo7VIHnadVYT2AnglsA/okRqsbJ2VGE4qzkWETKZyfXVYPDFLI52CvB9kXCeI
jwCmkP0nWcEf8V2J8SWKRpiZOR1X3Zld3s8E9WskVIozv9t/X7hpeJVubTSmBoQL
aQ5wbG8+sRMMiS1QicFeU+Y9wYsyqhivEdse92JBkNbfqm9yzyXG+0SH+6NGrGc3
9/pBz7yp6df6sDiRwjAhhgkHbCN/xOPCuK7d0S2zgtuErxrqWwHUBk6syj0xlaun
25OU6tzXyuabry3p/YpWkphwDmz/AYdtPcZJfppJ9nvddml4Mzr1h/h4Ej2S2n/o
+3uf1dcLKVNY4ASnxhqLrrX3TkVAhK3qyHhkw7Q0NvHj9/Sthb6sJpEUNHkGhgb3
jm1WK6A2RHqk1Kz79C3UkYvg/k7SyXdCDfOg1H6SjRBCsZKMuIod9GyUWOIO+DmI
hlQsjRHDKzfJpCzWQ43f+/yaJS9QYBGuGL5KK6QAibU4KpkjAPJqaVGEnLlAYp+5
XjdOktz3bKHtynJOihxOUQ2w/C8aR9YEZWP9+cf15E4u8ppnVEeywgD8A7a+lMzF
8uWZsXD1sngalVXRZfm2j8++1Y67eirrFAZyUe+0tov/XGRdez2lW54nLUY4KfDr
Un0ahQBl6fZ8jTGA3zaHKOBIp9tGximHY236Jsm+eMbwsxlLAUcyWwT5KF8jSNt6
VE8bOCWY+iQBENDkfFJgQWIrQWpL2oySzvz8hoNZLnH44VX06cBvtSI/VyDIMxCb
ueIr/lKuPBJPheIoF4Lbhw/XV3AK7kmgHjeSceol0I77kQUXz4YStAWw9JCVfpk5
3UPl6EJPrGtSCrySe78iwoGsImLDm2FoOmR0Rn5yG2dLXjUGmunM7OhjWHPJ7HsB
fkBysAbN5AUc18dzw0pwp6OLwHGiDaWP+0mZtl5GCQsD2plxjECmcBPIC9h+Zw5N
xBf4qAzjhD6jRBsBb1tEb2i9AW6Z8o1jzaMeDUb8oiSZE/alz3wmQ7wOxmirYora
N+eZ8UJ33glpNZqTAmPgxVS+MApFN4ZkXaefhadv8aiafy2uuGNY55BDf0hQdW7W
EB3hijhpuzcD/58/kAWKwIix/kTrEpOAUFH81sLUexeM6DbeAuRvYgHa1uY3QoBZ
cyWHe4zOCJKtkChoaK2+O+Kd34EH9Ib2LbuvO8Ghsb0BW2bW/kbXo6mU0cXoh9Tt
Zd+MOsR5C/Ixw9UZPY1SG0lyYUcxTg+yBVReSFZtHrX6TLeO1il7xEgrg34MdM9j
+7OyWTBj5dE+BGpF07ivkRaRnV4U3CHK1Z0deu6mqYbxwLr5VtOw3iUrFRyxrxU+
3cBZKhnEnX/6/+xGdQncmId62ZM1IBC2PO1Aadsqd4N7zAvVMw09DTQFGmpORNNt
1qwHv0EV2SD6XeTiu0Lsr8UwFC6YSRYghpZwrkgCapMDKBCmIJrM7l4F959txaji
efabeJvUd+pAoNJtkp7NJdhLH0TSqnj8+zDWzcTDxVsRLSdVfFPx/D4202OHa0qk
mbzKYc8fTtmLdT1pTTUAArc3uJmWYtMRKPHmALf0ciXCatpLjdXLRA+K6Mxu9Efh
RvmCkBe6712uYKECbnV09xwtQeAbTgrGrW3DHCJIJmqhFNDRVezk7jLcfE0rM8kV
QUVBhMn79nZ8s9n5dxPJYuJkEQNPjE8W9z0pDOF3LlCNtXT00szPfsaXNgwyO+Gn
jbyz1ff6aPVPE9JNgHkVu4PfQoSqbqgbB/kQHrZdlQVPG6p2Laqcw+DDI8HxXx73
/SrWwoofopca2dIisnpbhUwNdewy6T4xTJ9jh/405Ohqz1ZCIlzAf2KjxRaSDcbJ
YRX9S8bED2Zos6K3lMuN4PN4x6PoyyPC5EVdc1Mo7WZG0jALzLoyWAhB9gwv82uU
lybsp4cCLHgzdvWvrq7Cd957c9g5fSqaBjNUEv42iEt9Fy9i2a+EMw4M6jNNGcZ9
FUQ9RzvL9ClWIawbhcGjjhjJDt59++CLmwsvArjn0TqhR0yeA3nF8sM2MJTD8kjn
bSUg0NKPvtTTSY/w49mJjTIAFaaAIcvGi4M4w/SDB0DflcWzqKyt84cyFyTUvTuL
YAL//pVjdXNeVa0Nr5KaeCN+zHFyr25w+/FiPL5GCd/lWjx8j21AV3FMAhIfWBJl
Spi2uPj/l/2wQqksiagCB8/Oav9mKAdZspI5MlpOEHnKH+mGfjxULk9Vk0dEQtbG
AuhhXihEn8ELhwy16BiOQgghijGleDhX9BYC4wGiXuMRMeS3P8DC8UpZYgbNhVzE
KWscPXk31WIVXQ1h0ipQ4ruhvHaX0J3TheWmirjaXMbhQjVNzH3pIZ5FG3qvJI2O
DeUTgQ9hmbDcFajPNIziX2PTlf0VlYOa1f0u08aQxmif/rODQnYR6uzc9ptyS348
KhpJP5pMprTPS7g0WwQhpYfFvrs4SG6+3AHW5LCBZgXHjfonkXQprO3lrpyDXjLr
MuWqDy/tUfacCO+EJ/eOW4qjQvcwYfxPgF5paGRp+Rg1gGQLH6m/5NLlmq5j1ptP
TkWABJH6575Vh7cKp/QOEiUR3O0ST7bBnXlQ1xx8V0Xf+bDglBydjbcdk6mgH/rP
eydX8QhnJ+h/0RbYO//23Ss0wCNgOExJvMd//wnpIRYt4NjsonHDKJW8SXi9mNVz
HWwihGvO/41ld6P//LHiuHjST4DFtA2y44lIvjRAtKH4RkALRtM+0HNDJKqexwJt
LpqTe1DYUB3yLHyRFJkt679NepWlXtAVJsX639vwxcKX/z5cUXo3RC8P/gKHOjwc
ka+ycmK04Iu3vygT6wkAOKvVdmyiqW++tLrKvl8rieobwit2MKGZ93Lq4yKLHg1w
qwZqkqVEgY+pj2Nej/F5PHhfMghfyaj/E/YMWPuJZVYRPsIXcd4oxE4mcBnCnpyn
FXwT9/qiGmMadXShcZhLTUHBhauj9vwhjD6tRV/w7k1IpXBrn8NfiQnkXqY4T0y+
eFdoMcyIu9il2flxGHi1Pz32eiJWiqJyiPVn50nBB4jk4iVCXLQy8Uzm7EaX6HV9
eOOSabbUb0AXxJfF2p9n+l1xu47acvJrxpuqU+3U4TwAi9P41lxe73XdhgPYR8th
WqBgtLQg93dxWxuRRzZI8H9GVbTd7A3hndkaJZ+XImFU3y+hLcm1zD4Lnaw9Ia4V
ZdK09f6EDYhqak2TsP5j3uusWkNheg/4OKZChe2d/vrNVGSyc8XUE93RfaRqt4aA
IFnDp/pIjWyNTc9KViHA5KgaTPMETWyphr4gIKGyU234lt/pASybncOzY/78QnG0
FIVGGEh8M9gCKbekCH2xFNGvtQ+sLEtEI/AKhNSZV1ioGLlHgAl9sS3wPtU7sI3D
D37Sbd1wetJx5OZ6oDBDAVTuhXK87At5o8XmpqvjBp2RZCSgdNyvp0WQ6JeSi/Xd
MbJcT2YVipUxJS/NppJ7F0qFL6/eOL95ZjEV70BwKA9VqihVS1VeO7PdOv0rwQlU
9W7PdpAPfzNizZh9hQ1vtjf2uXqnz0UpowmOHaF7top0vkydK9BzE6PKtrZM9jhJ
KRBOxFFclGh9qjmAMp6sRvAD4kpYol9wEwb+DlwxXOmLRFNa7pJSz/k8aOF3cmZU
NU/NkNaw4HeS0kTmNXUBLXhAe7/xAM518l3oFcwFdi/bRyEUolT8tEq2Nf3x+5mS
mibOvyoWf8RMPk6yRZRkra+YNDEIMTsLNtNzLGeH8E6NIqNXd6UnpC4bLHP4XSXM
7i0pPo1qyliHUf5fQn0zKvEVZfCBLb8K4f0M7b/MwTVSwFg2uE0QojsY/Efaiyud
cv8YNlhVOTallaAt/SEF3aSZzZ6Wgt+xha/wKytuXvvD3P/nFH568JSOsbUcilKY
gHPuLIrxTw/0chlNkIzwS+1StOTaoI8xJ40LW1Iy9vt6Tc9DiZTONrCHR9s8ycTP
Xt31mjqW6cot8KH7DPgywC9t44zmESN4wQGBwif1fFBFFxbkbdkLT4kSKBQoQP28
OcOZudtqAkCSVPpKSW6eAwUnlc/f//hmk0Bi8aUSpsadA/Tlf5Pxqex8iU3Wbjfl
OhtnKIfrknD7b9B0TxnO/KVfgBGgPLfYO7fevk6hQZz7qDM1l5umM56fKuvgetBR
Ix92aR5wf93TaqVjBT03y3bAqjM+mCtEwoUMImj2e2ZqOFWrgNzZzdU/AIiljKp+
h+5yX5KU4wvmvgx7tM3cR6xijfSkjRSD0cTuGeUuqkUY06sQwSoxLcqRUpFPwgx+
j/iOZ5QBpDPTq+UeZWu6BtI+qx1DCm2z8Y8Y7HNm9S36uh4TXwHVRSskShmfaCf4
x+T2vpLBvzmakaESp3bhJqHAmsDJD3IofiQ8D5DQ7zY4JRMW2JGJ16KzRmkRngCr
7bvNn/YUy+8uj2MqgF5Ne1RtRkbU3j+B3UgfxXGxuNShUswkS0ZTvc9WiphSSkrZ
HnAO1J5Nuwi0PnubsajfLqdTp1cG5ErFSiqRcvxmG4wkf9JtSXpAv99GfeOoUOI3
i5irJP+sVDCiK+O35Jmyj04oxgOtrPiO4fzZsS4PEy+xbQoWwlLeQIJq5RKU7wg8
pIiwLPr0oPHzYw0JkD4aJd0NA6IRaDAeauwkBWVuvB8uMytVS3OINPgwE0Vaz6fK
WGfy3+1Z8RGfgRUMl2INg/Yh7wvI82eeUEWxKnCcCe9MCM9XP5JC65s8kP4l/rv3
OB7ET+EbxMv2tQP9fEyQzlrypO8jpCO4/03MsnwC+znrcJA23sV8AFe/ZfpShx9Z
DxPgKi+qKmK4+xAbPKfPLFMoHaeFxb/hk++ySnM1Ok5jWRHFpLgyvdhUjChRQNln
ZcXVv04fsPUKZx8tJEyeB7Cxg/aPk3l8tMZYfXDIKWJ/DAPy1YBMe4aqC0gRZB9G
DKT6yZFgKkwV9Emsz8TkFAp9wRwOllbwN18zai/x7OdwXR+UV7hc8pAG9XNkWJ8C
5IF4J6VzKbb40xq6h6n4D6+sC7K5HRspGrEDR5gf98gcl867SdQwJMdW2ok3C2FB
lZNJvE21jNxtsNM7B83z7vm9iavcW8o8MyDm6ZF7+dy3YMC39dBnXJFgZ/EmmCVC
LHNx2fScJT39EZ0TPVjNbsaTG5P+C9Z0bZG3rGFoUq3cDi9gWyc3+aN6gpIrrxPG
1Kd1eDEmTZBn+dnFxifhbXhLQFREtG3ogL82xfLogLDn7ktqgjKiDNZR0osgNxzl
Y8OJbFk5d9wbg/Adg0Ooh7b2Ky+m9DJkFGRVXrACSnllxz2OU131zOnyXpHjkvOa
/YHZVpoASQfbm2nVtor1CHS/FAw8rWtIhaCLXdk45541fNFyVcZaxEfoML6CCbcE
2gPE/wDrAg62IllUvDdOv5PuW0kUoXSL5xeVxS2szO4R8r78lZPlA5KxPhsKy3YU
3S+RfoC2aMwlJBu5D6vRvhr9S/Vnpnk/GA6vLkvDVYKWKX/2DLmIpID2mewXzWNA
+Z4d99+YJ43hRV1X4E6pflc4ALuwJFLM+HZFB78N6zaPNjf+ESMmgmD8bFTgn1DA
nJTci6LRrgQEQmBiwTD6pmloK3wnhoACcjyxr8Q7pZSu20ocj2gPjS4Es7jmrWH4
hjN4/m/Zvyy1NpgNVY4C9wmZF42xzfeKwb6vG/Y/uak4S+jhv0IPle7j9g0T9QcM
Hvh3kmSLZOrYXSjYgPAtKaIEHuN/U0WeEiOrlZCKFiW8ZvFjszwA7met/SwOsBsY
tSAHXnVKMBUmpqVx6amDfBWLOZzM7K7oPOMoPdqx6S8STYH5cXgbDjQc3Cg7HBeF
XU8RNcS599g9YJKqnOwDgtrPNrEFOXs0Ziyypk7hxpZyDFy1pxedIjY9oKZ26JH+
zph0K9BTDOxTrjB9my/PUlKwLlrqkbY8fG9QcZ3BkkbswKj9KulOIG0x6KEHe90s
+WPnDYl1ysyiNJ3GvKcPD5jmar+GMO9ghgNnDjyRDBuZnsKAVKvu2caxnYC2Ubgp
Mjgnb0s4bESveGVTC4fb/D4vxH/G8ypHc/qAkHBbpe4+IIPj9+Zr0VyFFzXTLNa+
0kM8vNvoVlW0dB3qwRxpDSTUW3JJCDIrngnyAtW8UrOLAYZbU3h/8mAbsnTsOkeb
qWXpS+uPBSmpSycacJVP+hVN51FDdYfV/mDzspqnHmJAQj/bFkIUrXMJg4+P00ZO
IrMT5DBWNdm1dBwG0VVK3qHUh8+W5twGs7/gnF+c6e1KBJMp7k+31fXZGbMW/+2l
qb/iZSZSkQ7UvfM0UM/RuenPRblrQJNBpkzs7JDFVLkbzYubs6d3f8jS3dtS51Qx
JVi9injyPiWepyu7zSrpdN4rbSVOSZ0fspyZ8Th5YGXvHRnZyl8nu/mEDPucDSd/
RfXR3kMpRnpGg8pVk0BLLZvZDlxV47bLAGGeNgMTy/oz80hS5l2zksbJ/tOlKNAK
SE18ttcnSDkBxs2q5VYq596r/DGIWit8RJ3pLdkEr7BaAhTN9MseZZRLAEKB2NEE
rFMLVrcuPKNr7JRmRUWZpnKzKh3klfdpiEoUfVEE/l49uw1hWWJDV1pi6NnXCjsM
3vFfOMYTbwk//gsYp9PVn6EMkUlwAaayPfRvkeY6ojnbp4tJvwsAjF7N63WAWz6h
ZRTL5KcmDH90Wimd5IoxTmH6weBjX9Y1943uTSByrNytzBmHGhnZV3DjCNob5gpx
N20kdephE8ij2gHYaKH9RpdYzlEwHWuYDVcLhAQfWW+d9q4M/tNaWPJ/Q8uTAocK
dT824V1Pu9J0dqt+moIheEF4b8778ozZhoetvzaWqUdNMQOvnzYlbDZXqsreDiDt
j1eHZjdWp4pY8ZJCqysFJ/QuGZNruCTlDhOeBnB+iuVAYu+GDsdXl9899IOuFR6Z
64v6tm0UBoH9vxXFCDsq3RuAhAEK6wF5DiszEQHRw7rrudnALiTil9oRdE3++hUL
xcJa20qI8ymy+vT5lUSleUtJ8VsoAB1hyFk4OwPalpDCXdjRSCM1LDaj/MbtMeC9
732yPhfbn/RWb8Xl/PP2uwkNt/QWswtMBYUDSApaC/qEw5X5ICPgh4yqTM2mlpLW
TDHTK88TdknPRQHE9438NzX/7ThpGZKADOfBk4+u+1CkY0Jn1MXozzoZsNAAWqbi
Ty4CHhhIk/Ljnm3546vaqcK93Khrcf7gNICqpEG5cu1H607vE65/qVtS132iqfxv
awm9AVRZ1aNV/dAvAh+wWVKmlWJZnKMYjo03rtAPByRZwi5yqXb2AmzMYItauf9j
x3pTOcpMcVXgt4/hPmA7WOjVFvx6+ur/W2ytEplwHejRVdYuvc8+vgE9t9Mqg3dT
7HqS1tRYK2hPAdeF5COynbi379UgQdqyujNX910q+u/FlqF1LjWji2zFVrT8EYDx
ZGw0UYdqdf5lfH1JLvQltu/AuFFxq2omB9D8YdAtO6KsdFXKYh10+Tj3N7X9xH9i
TkJRJmG/1EpKJG+AGv0fH6F5uUo1+nnPVsxD02gkxm86sEbqcGPa+Pk2u0Kg0gYK
yWhf/dB8zKm5pG1s7EU7yAf5rLqIye5OSy9N1j3SLSHkZ1wWVTCaVyHgJ+NB3GuL
ESj4Dh4lHFgiABaD5k3KvWsHmF8TtS+5fev5U6wTGQKSkviMRg3RhBVfwUmBg9iY
Ler5kn4OA93t9t8BhQCtWUJOSXrpAyXoJ5mY6yJAnWwpK9ntG8VrkHEv62sJ3Mvr
JknjfPOV8I//tk14sj6RkDZDrgGbRPBj8UXT3FV0c5U7KqGKqraP9V53infg3Opf
Dcg07Q0CjG181u/Ft8VPgEgOROFHrP8KXzEF+/ttxcC0LCm3TfNZ6FypgWHH66Wz
BritkyT9ejHTyH2AUUgpxqqnW2WronzqfEs5t/aoffKcSDp6lx7qJJZ9r9OiSCFM
I3PDV9HjzO5b0SeC5ZOAa5dmcKBR7sQXa21Yk0cy5qShjph0LosXnMSu4r9F1K6T
luHIpFTKc2ybdlTpAHMVOb5IlyzBhs2dk8OX5HeeWtIN9ZVpv4diSkUTVf8Bhtyy
7gOpE2Ti4K1/eiABOer1LiUyEL4wWqZzn2BkkdasS6oPGD70C1zdbUZECEEbA99u
On0+4/otc0MdXHEiJjN6sTBktepMokG2tvgVO9rmPmuCEAnzS/+eQwrqMRaTm1yV
iDICdLPCzSHavd8slNJyh6EAxsQmXzC6DsE5QM0Bq/A/IjPaEO6haYgbd5wuw38p
7lAZpeMwjx2fZJYVu+2Ug1ZsV+GcwjxZmkbYlM7ucfOVObPSg2m0dMed++Rtli86
p8IkOpl9yIuVXdDKebyub5t3kOHFB3QhEnzubwc03H7UcYQXcP14CMcD1TZ92Gj0
VCRNvdixlCjQcN2LwpOYL6h1WI+0mTZRK961v8hAZpJSMWH/PIr1upXwv5Qsib6r
4YRTkk82MiTzDkCIy2e4abK8ZpCZXQnBD7Fb3cQ27xQilZBAXVqxFFgFJ57FXlOz
gLX2R6ACZUbWTU6IOpnpdgy6wjXch5yktnOqRFlODL/UICelz6cZCh5VDwc2qExE
Ek5Nd1a6Osac027hXeZOupIU1wc9Bg+zlgOHMoupAH3uAEZUyjv1Wq0uVpxXAXVu
paJJA2ACGvoZCzADi79yDdROiueKy8ziY8PnL+Mfm1bLBfR9enffxSNvmlezL73x
6fAU1ewwgrecywfxanGry8IU99KMx3LtXZ7d727JIEVa2RPSEA6409+eU1JwzI8u
MRYCpgCC74v3Jft4fmMeh2iwC46b0ahOWKaptp/5QFj37uJAqVH042P36eiDkrhU
aA+50sYYOflI9qGJ3AvgOmx0acW2zUpXnmd5VVZV82h8aDw2lNMqz/4h3rCjGRiC
iIUpywSeXksP+v5PQno+erVrOkh/jRXZR2GUMqxXpwARJqBXF7zavSVx7LkhkvsN
4c7BW5AbOmuK7PGj7O2G7ddxUdfrN5NHvti8rYQkwKs4KOFskvmGT3ikbEMma2RM
jJdKMIjFbuZKMVvKfs9DVadEyPD5L2o1C3CiPEnRYzYf74jIVv0VPSWuRgdW2YhQ
0gGSgY5K40e8NdCtAUwrk6AGzJEC87haM9HI80DLpgvRO5JiaBaMZUKLYFzaXthV
Iuy1aiwvfx/ZD9ANwvhqZ7C8cU5YGWCmxXRqs4M+yrTsUQLX+Abt9U+xwdEem2QG
goyY0ZiCv0LKxSTtgEvC0BcwcfWzOhQLzHz3CRuvGzsKYctTv2GNbfJCmdAAUaNa
LBnd2VY8NXUNpAL4gniuSXIwipOpFSStVFL1Uol/oaq57broHaHOcFqiKiJRJPp7
xQO7GdP/6VQjUXYZtJ0O5LLTt2rUrNB1N+PJnE7N5xKhPV86QT9eSkHW8P0BSzGa
d2YSZvzYKMm7M8Rb5fSJl0GCafOVzxAG+cLWBINC2aHOMUFfWrxZQaqRzA0RpbJ2
OyGvq5zk9hcokHl7P2zuUCbizMS1moIrywGRq+OwCVEFQXfDffOLI1/wyFsXULhX
9SeBP5YC+TMcsIedVV7I9nX8strlItWCsSZZ5ubgM4klLLEZNdQhAY5d8jXiUqA6
lZSwrs8Gm+TfqwHdv35AMiz+xNctSdJBMv4YjuCuJxf+rKCi9SfjfHE2z6gZ3X1x
DlPEDleUfv43890X8tClgvm1JDNnD8jXzSukB+g6Yalj9SegRv3w6Bus5hd5pCiw
mxbB2QCRsu/AY4y6WNPsa2bgFYpurUejD2zHm8uW3kNsijn/GzZ1x4b7tQ6Gp0x4
z+/il8Auea3Lgxz9uI5P2oUU1oRoYweTH7Q9GYH1yoB4k1MCKh+kymZmVhFABraZ
DwOoWN+dNsJPudbf8pWEQwNJiJ8z3pU5T1JLoWNOYwAQQXyZq8Q0lJQ7Z3h08MJx
o8QlV3KNCCxMYFUoQqQJikUbCG8csmPI6qCv1LqzrA+YoNkecYDLsXBqLmOXE90J
xau3KvJBpbo2RmBj6NX8pHlxk36sN6bk1+GqiFyI0wq+9baEzRfD/MmV1GdN2G4Q
a1oQjPfNCsVnpRehaicdlTWa/OJU0oXPm6FbIAhacBMi9TsBKicOnIS0SjIRlRak
hSkPMPkfkt0LW3gDU030DHgVg4HdbMDcCUu+6RGEw1DnggH4cLR9eb2jIRZyWdwo
705GZKHQ4kBxsOjpb8XYqXeBndx9OwQ51jUess6T3+7ws0jSoT6KFqu4LsO5Jmc2
7hKE6Pk5jX3yON4sP6rez+ZAXKuocsT9e6LeKnomRHp/cJFdw2lakxd//qZupLX+
OiKXzeaVlfWNjq2hLtOSuddgcVNARy02Yncdo3eER+fyoFOmr7lEN7EU2VdP7wYc
91Zfm2AlmDEUlooDurlToxdvhgRWuizSOcHQsg222L0bRL/yPXGBZAeo41Vnk+XF
WQvvrhmT1t5eASFyl/aU0CH5AnBgTar7NwJn3FY90y2bZa3BwSynnd2+UuVcwt06
+XijE9pk4eM74Y/jT1B8F7drbLpl6hKm1bk84qN+S83iS5uHkiMGQdZTeckkaRPX
DXIESuXxas7Is3wNv0KVmv3widq+XOyuY+A0Ve5QhJtz2zi0smX/xFSBqS3M+k6P
vGlNtwCEvgxvdxgIAxBLH5YKBn0odIXqCi+DE6WH0EQPKL2cT2UoxYG5PJfCMpPz
OGISNB4dG3hljOaq40YFHIZuA2PDhHtp+dCI09aZ6P/ErY2cYLJgyfTXSY26Iecz
M9gcmgUm60qexWcz4jNAzu+qHPnFQ4JCrhaOfeVw59FK9Ff4Z9Ozo8FKUtiBtlJV
yKs5T4sXqSrpAhEaSefWzDeiFSQneGVpiHBaTPe6M8L7B9ddKRYZjoG4l7pF2Pyx
IF96pCisRW+3+B03yQqPd5xcDgVRrWfKn2JgHMsWpqVVo501Jp+5npnAYvPBe7Q2
U9JSuH6Q0RItBOZge7C57GpLqXjkJTHWmsNxAdC0UHC7cC2xjBFRJihDi8o+SsP7
jf74Gld8rInW18BaoWXd9zR7z1t5HerWNLuf8j9+fSHeGywC0XuVL3/qJlDMjWs6
qlUaVLbsIHJEXaD+rcCXupZgiHE7VWXU/5N7R3I+jIAKqv60+JcQt1fr5UlCgqGh
cnOUfi5jeImnb9xvVY3Iw7uEyQySM7ggVOf0bVaPj0A/1vaJtRp4i9OM4Pn3fP4o
RIVgjIaGFbu6xVOcAMoyup4OQwKw7z4Fc7Rk1JyDg2Nej2KAMpU81uwowsRi5AiQ
/vR6KF4Y3+6JGBVn3ZQp2OT29chFJn0fnKGAc5MPkPBbknhpVTPYH7tkueZJQOPR
YDDS3AVHPNoM/cHJApS46Kn3bSxML+D1XbCvitzBbjatNSvZyggc0A+Fuvc1nTxS
ODWh9R98wyZZgFtCiS9Ow9yEEDuyOQdJ9aYZKwVje2jFGSnqxXLMqgxROYUPvmfZ
QItJTngTtMILcbVr4PLK3QcWZjQvSgL8xFTQaUU3KDf7vpkUWqHp00XeBtOd+8mm
t+OBDZP9oR2dOhe3H8oIwdgX52o8NgTmGclH5/8lKxMlBc5liH8MJuvsA52cVKVD
djEUHQgTkBMaxdPf2tkERf/5SV3ZZgw9A7oy1QgkeL/ih3wT3oAnPqc6BGfM7+i+
3YJ+kPnriLLgW8XX2UggRqREOSbwVwkJ/7CJl/wNbgJp9QdFBSfnMrGuK1mDpbZv
SSzNRCQEf/7Rz4ypl87a4kkHLw5P7Mn3B/0o74D4XfWx9SgksSn0S9ce5b+ReRHn
qUN+oBt6MQE8R+/F7A28DfTzK09TVmdShSDAGRbjXz7RSYmLhDeADAiB+EMUa+BR
nB5u57PELL+MpOyh57/3u34oQURK8O1XbdYAca7BJnrqMM7zg1sMd+i7jDRqe9Cw
tgcxlfIkeEkSkl7pYdbCO/HkQiCwp8av1Qk43XqFzDCSK0CIIyUVD/6S7r0FS2u1
C9w7yC5V/q7JTFpwRVuJej5pbC/QQmeI9GsIlURplMnfcjyHDnBM1dxigthRH3o/
oyISTo5nSMnArUAzLekAXL4D0o3v5nFYJStDtpY5XAX1xKaiMg8CUvXLss1HlzQW
fkDRksiKL7s9ycBF8pHDV0wzManJ3ognHJ4HHo6VK7bHFFwG2NYL88waDO5vFF+z
inTRU/78w5Epm48TkzEu2/Qb19po8SPeksS3TOPnZMD2/e/HSoW6mUQmhcDbBlfJ
8JVjIZgJEDBXBKwqKuA2bG0v66p01aWwayozhuiBBrMUUEaf1zHOhpNsQV4GxAr2
yG+2lakDhCi2y6EiYecIp1M3OE+BUBf+J8F4+RRdk+umFgMy5zk6qvPYvNz22zz2
fNGLEoutdd2RyCwWJBHv+B8LYBAtCTAq9laSk4uRM1w3tXzvd/nNmfyI4ksRp3QC
WN7trsGGvgeLkcGZx4aufIlSbq1oczCRgRcrjJX8TilrO46rfevUwzXu800ADPT3
zlIBisquCTRTtvYT2FVDp6cIwn+M/tqFSVTlWPnikdiwG2xFuuwHwIvu5xvLXAqd
uSmonOj+AXZoaZ6dgV0hdsb8T6ZDK8zaVQee7/rFgl08PYds8u3177wESuplloc1
8Yf5aC0pYFfCmRRw0FKzfqaFxbYoL+vEf8ily7LGF1653gpfkSNnPKUGLvntMYb1
4wmOYNnpyFbBiLdZyZ2pK2rKQD6iJlJrCcCuhwq4hNJEIIDOSCIBfDS0C6vGt2C6
ES96pehxsaCwjXgotXqXq8sAnS80OGEAj1HGrCWIPpIZhuKICP2hyDz8d67dssCH
08CoY8iLLrFZNJw4Isa54f1KMnPk8EoiFwgr6npgJITTEpHkI0cIKDELCQJMVB5X
/KECQ5atIDVIWSYNuNqC50EeVVvcyX4V0/HuJkDAoDJonBEWnavqhTKS2T/5m9Iq
U8aiF1hvcWk6B6/j1/k4Uc3jXGBJPerrbfol4PwmRz/CiPCJS9rvnv8ntdxkILIH
GPTDawLYt7B+teVAl1+DFrTc8q8cY9U574DTjDPRjqI+ukKI1oF9qkj4T4PJI8fq
Ny4q4cbDI3Hz+M/oP9vOTMEYO9q/20XO5z8K4qrfjh4WFbqlUmhXKSzcYMJVoTGT
DLHqLYey/MNQpA3onev9WRdNEr/3rh5Agz4gE7F8X3gm7t0n9AI1NiSluN0VRbyi
VwqSH0FUNVkEmbI6aaCrKwNUv+r0iTLMTadwNjywW6bHeur3rxUARJwdajUCBwxx
VUM894e+MdC0loTu6SG13mkGK1ji2V2wCv++K3jm5WrX9nskQMNvW7PfR80SlBGI
IZUc+tCu2NEUx7MNq/v65tWqGddBUxmNwvbfrbMJHnxAmx+9r9Pbmg29X1zZcxT4
EHWZzUPR0kvVqIoiqdbwlA79/8g8Pz/iixa8Q7JN2hubEepUpsmghAyP+NIpS7ZR
dp+ltdjFLc50FLJNtk06jukYTsdV4BiLRXT1VBNMw9tHk3c8I5PGqAclZKvHINtb
kyfOLN0ZO4PREbM6jVmly0B+nJSEL6Z0ou7gE8RvoLV+ilzTB5QJttRXse5y3eH1
bZ7Yu++xCXWRH5GRrOwjbPvqYri0eDqeS8WbxyvL9ReaU8J21Xt5SDZ/BydM8cFv
9nb50ZNifcCjQh6HHj9pYQALdHzadr3mSmGOqYv7o35sqibWTBX8BDWH+0OTGKuV
2V+FhoJhdWctCKN8ca3e29xTvR22C+xLeJqlbGIYChgvCKJimJ7hyQdfSqA7dYTY
IZ3HVFrMVu+Lw5ZfKlSepKIbO3Fkvgcr1tORu8HY3WhrcPC1tnYgxorNCuWtci+b
eiw7erbq10LoWWqjDZMFJXX7SST/UFzcBLBuCc3rtITa1/pmRWhTmIsWK+GOACp9
t9krZH44xD8Pk3/SdVem495opK3D/rGzvMLVl3X1KYaY0fB65lj7IZNRj9ynT+n9
3BXOvbFNpcTho8U6wMCUCWhArRDPwNNhFU63Yy5XDlpMT9K2Ne8tIjul17lr35O/
KqifWzpBSwWX3FfA63wqxcjZo1yJcuQNpJ3UxHoYqmdCaI+Lt/YT8zWS/TVlmRPD
eoE43EgljcntKuC+R6wQmcYBrGJKNqzRpaIb84zdT218xOaVMkH7Eg6HPBtlHzHt
RXx7eYbp2Ieqig14c7Ayuc2ds4zXZ8DHt5e60lEdXpk5xK5UAe7E0fYf67i5Pk4d
aFilmo46xOBmtERXK97fc6/QCLgIM9EKD6xjHXDdyxp5j4nlL+ZMIeS7feYH+8/e
We/IlsJKwxIMcf/arDiFmyDE5V7NWEhJMiF/BdyKtQ53Td4chJzx0153jF0wDQB/
rK6dO0jwgwB08rdlcWaO5BYhwcRvJIxWXTgHA9fj2sX5/GLwbtdc9x539xpMD3D3
5mpW3EgkQP3Hc3XiWM+7QPyPeMvawX8GNm2pNKHXqGtsq/nm69SiGG20Sld6vXog
UyUHaet1PrkzjpsQMhPj3Cd+ilafOB1xBSvVlbfBJDOsM5UTt/R0qc6kJ41mJZCw
vazQnZ+HYJyhQOjDtAZoM8dcMtX0Pkrwn1tduGHhndQsOzuTcg9eSZ5+DDgmpIib
v6Qe3C5EbJAwaFLVAzkk/5jmS3yhWaRdQboBkB7UerAHG6I1Zl4xq2VRBAyzCIio
1Yda00kP+PSJjhq2N42QFTjROcYy8BMJs7ONdH7l/Yzn1s06zOD42B/hj+rnQm2C
JmkOeiIhJicDkD+hZHX1lTkvdYRitBjZ+eV6ER2uBqJuH1GW8FL2/SmST85p5ryP
B/b+NSmXXeMf/GV805fKjf1hwJhmNpCnnFRRrDJR0ZL+nyESRholcM8tmKc0vC5R
1s3Vf93Fz9JJ7fY9b+FMNiLnuGf0LHj/WIuCSW0UZzv0RL3wWcSNDL7pShW/M4Lg
k+hhZJClpvq51Upvsaz+fZHOpbCgStDrthSjU+gSKS0dj+E+/X1Z/WG+WPhJJYAw
A7An+hdfz4JzeK0BCHkd9F3UyR5gkwMlaPjXphjEbJ3MkfJ9ZqvwTwoiVwK/9VG5
uW3N2QKvauqm+cgzIE2EOmOkchAzCLeB1U1bhvtjaP0ccWlwwkD04pgi6I1ElTB7
0AfzGRPx39opI1OAnQcca1o078CxmUsULj0KNns7hzbOj9fPHxirJEMYNnAhpFHk
46f8hichTejUPNM7xaPdn1Ff8hZNUJvSTYgSgFDtabufrSDtF8d2nO2yvTrzNbpM
J2aFGT4m4cXk3TR9EbGolyKbWkGnuqFnv2NfIVjFWxWXGzhsgfPfCJMmN752vpr3
Hc+Te4S/MsLyI+YSDPA9vX4HRelq8jRGIvMW2nRrXVmXGWnzaATpM7oPghkbX/TX
/G6+vObapHSybRhevFESS/wQnXe5q4aUy+jKOhWU9I9aOsoyb99vYnmLxQ43bb9p
yWjixpR3COXVP2PUfXZT2wubF/GxtUCBQUJKnhVBqHvmZl60xQ+gxpmdrEmqiENN
RYkax3aS49w+71IzmyC4cthF9R2WqUek2btgX8AeKvykFxwbReP4XqRtAsciJi6B
y4fjJcFK2l9apFXAZKaHyLJ96WzNtvA0n/8XMuVpky0pgvtmTWWO8gIeoCjdF+Bs
sSnkSp5cxEmkIfQjvDZRtwb9ZSwYJNxJih9GrXxpfKPvhU4jyWMjc74OQXVDn6pQ
K+a268juavQVGxUEXlY3JJIyfgl4H/hahCOTjVV2LO/YcKWgH1G52igyFZiZYJk6
gxRrglXtg4oZHt4h2kZbabmqssii4+j4H4NoS/bq2OvZs2AUF5ehxjm5KH2o34Fh
OceFtQyn7NQwUtYehrnB0jxZaq0JmwT7FN8zdG61uD3ESEvKnPdqAdsCLVYyLP4W
Qh0RCjmztTf5anEh9zgqPuZi40YUEgshz0jw2xBKzxF7j3Ilep/LAoTeHtN5gJNV
mWfnhF3xTLc7y8l3VhQG+tDou6eSdRqwHtJx460CMki3mzE3Eq+zteO7a2lDua5X
IDvSIYGV+PtrpoxRxC8CATEqFN8dD04GSnwTB7BWmAmMJ9zbxeUzLBOI1kqQOIJC
NSfzaW8r52c6fDWaH3JiNXG4GoHslTEeILajYRrM+1he04r5gpWuPnzdKyb0WKQL
ssuX9BynYEY2rgzHuoCPwDEoE8r3k+tZqAwIuOSw+3W4nRJ8v8QoeIsZIxuvxiMV
HnxHc6cZQg0LhasWds6GB6PVkC7UrfHTpnpU+o7vyqwDdpu0YxDPjT6QmhD0RW3a
HeTc45n47Q1oBQ9y4g04/W6peI+B8hvUZL9Cp7I/86yLDvByz7oTSC4FJZWGuU3J
I5kr45QyOYIEFuYB9IwEgo3Z01/HCSoz/THickci/lzwxjpi9prMcQLhX6cNKAmS
ifu14PdtWPOroGkV4kP6qbgHtROFuifRlfCgA2MOJEvDFS9xutWjWpsSbTXj+vGT
9zeipp/TU3OYGaTCSj5qZpaJoMQhtoH+f/ooexpnF8PZKj0RoV1POYUwqNY8hzpe
3z/iBsb4mXkSz6IhMAybuq1LbapfZcmPsSw7nbe9i/3Tzm44mbW2AwYjb0bcBOsH
cZPWcaT1epVybYxxR+T405z2PSOd5PsWMwPBn3iPVwO5fpOh21bHC3vO+B/6PEwj
YThNXhHqQczv6NfF2c9lbvCfzyypfZYsCMGtuqnUOMr27+Eh/Prh5qJKrM9YpMzp
NSi9OqIGoEMOsOanGgL+RPXGPwarHSYFBhh6N1b1vuTWABEvZQpO/bZJzfeVCWZJ
P2Vm42dAC1xzjO7WHu5PVX2lUAxEFDkA+bGKgN9b6gBnNeqbcRRuZtT+si/fOrI7
TRII2dph4XwtPesSknqnBeFirwn3J/8nFGB4pgC8fbC/t2TqvgJUWZTNTMppAIUR
vow9nm5/Ims2YiI2AIJvA2OifraMpxH/BDPvdd7TCpW9pUgRpWBzj0ohbWrTtw+l
KS+1+P4Fp4C6rN6RpAqQDHxboAmBulf3F2sxeor8WQrry87NaJ3pSS0ox3Qeti0q
92YyAsx2uPBJZNBvR8hhbNRyeWp4bcU1IZ6uZodM/NjO3+e9dCXOybMjeQNG+8UD
8ok3kZbx9xIuaG58pFbfUwYI8dMPhMA386pSz9RaxA+K75jLDxkTDD2giwp8BlJv
Gp/aSfNyFMf1dg5S4llySuo4k98BSI4qyMUgNTa7KtYDb9ZftzIg4BOF1KrzDoKt
vxNPPWuYKSxSx/ENV8kVqNxAFv9J4lFPoXG05eX84/cwaNHJoEBH2ZzuKtIZs4fr
J0341WXV2ql35WYaj8DKpqhbG/f5FvTZecGOZQF6JRJtdod2VCKgeDnCrCPJFTlq
Uh8bN3is4Y7w+vsw7oF6eVdtEixkHmHSxS7GeD9U9Zy49SsKJZ+Qi1ASFkdzVzXU
ud4umWHIMfQpaX7Zj2Up0wZZVX8asg06XwVZ6/spRLWbZlFv+sZvfHiiMtTo6syY
DfG48e3GxjC5Zq7SkhsO8s7zFgiq4g1tiOfitWWYi8gr6vLvRjEQj+MtoEY+6s1e
7RMUeUzwZ0Td2vGL7ECo20gkPHWsBmor9qx/gwjcZNRWyM6dDU1HX4LujMi7hCNj
dpfXoFmJc6u0TYoo/erSF+d4+2PXo5Vr7DxKCO6lYAeunub3XyiG0gWBdVoa6UI3
bFjwlaQ6mnaq8oNhkXftl4gerRowmvoAEZG8j8gpPB9rbnr8i78f/ErnOEIKVOdt
EhdPf4ksoKRKXoqWz8ugCEAUFZCatvarqAV/YlqloXAhFoiqYGUl0lPX9lF+4j+m
nZxNju64mWeF3pF8TRN23flAulNZSRH19gSZCKQDWHhJTfm+Pgg9gVc6Ac51mRlV
elqqygQ50bxqk6e7ciixG2TRkfQ+jYW103M3rv9450I7YvgUCE1HPBnj+5/HsLt+
18eIE2JFcGdrAzXlz/SqGhbC87BYSbMD90lq4yiLAZpwlvwqmmY31WGIKc2//zdK
w7DfScFpMMcB8KnhzImlULXj25OgpKEYM2Bv8ykPMHTpqryxl1PSFzDuRxG+68L1
wit+qSY52iWcalGfKBF1rE2hcyegmrpQ/sPSKccsjeo55VVj8hcnbahTJilNzoI2
eYgaLcea0223zcxFjKNuSYiympAV6YzTOEZxbqAng685maab4tGk70KsCvchDQUj
q+ATavY5fFeKciIvkhiK6fahdgsrdlCEM/kcOMU2TJjJGqNUcYNbCkyxJ5b4K7BS
dBJMNS4yQlk5qCVndCh8K/4MWlYfyhCofkAq7Adq8n17MRQ08RjBWWW9l3G/cvNn
gJl1m6PuCOz+iYnoiEjmEj16DvoEK2WU3BvsMRP/aUxyGS5ugtJMiKyPNAZOvuo8
xg4M6NwaQyhsl2as4GIHTvo/F4wHITNKyXYcytuURlNJoNuss31IT4gRpRKnz2n7
6+bxsREfCNUSu/MAqRXj54qXm/b4SOKl4WklhMqSJOsfyBgFfuerapDDbVcjadVd
uvSb3J0LWzbz42FO2/PeQ+qFNrP0xFXFZffj0R5KTPK4biHWoV8l7tl8w8rxrta8
mG3dwB7GbSa81s7jcI8CC0JbaayUqzT/IpFEW9UXasCx5fXJI3nQp6QTSAPn2Pbi
5xCsgiJVpZpIJhG5Yryb+gxuxmSNfkX8HjYaXZ1w5PAAJ2G3EpnbfShr4BVYnZ+8
WsU5nGpuG/gE7z2Ywg5D7J8rT0zLVUUz94zQF5mRWg+0ugGAQ+T8zm9VhgVGFL0I
WI3Gjs/5v+Gws3RC4euFCBWbTFY2PhV0ubpa7tvdfsk9aus9Xv/UeoQr4N0rrAlq
cSEwfh3e9xaPTbdNdP5FdgKCjNNkfsadmeMyUEpJcFEiYeZcx4VwxTKtVxEuVEaT
oT5hljfbP+fuKOGMN0riQ6vSXmgQuZh/uQozzZ0DO3KuT2A2usBwBT1Plq2Mdkn7
py9TffhCs+jNBGbMu4XGxFaP2cQkX0nVt0b0UFDi+tbyfSuMMzemwoLkDgcYQXP2
wOPPFQDSAWqmh2ytXYLLbh3NxcrtoeA5AwIT5v3rM/02NdOUlcAzduA8XrkxYK+o
KEJsTzMU2JcToD4w+yLFugOwUmDZKZqJLj5Jb4e0jDuWcv5h2FRHnroTF2VJD4i4
A8g/SE3HHyzwb7DlQeM+RR+uRBca9KCDyL7HMaaf/JR/u/e+YEbGb7vWm+XgGdpW
7qXLdskAXLr1schHfb7F8nQsEx0ZS30VjdMHRRqAErxGMI+EpEW9tVptKjdDgGp7
GwI1187CpdE3xm1jLxquUjwhu9NopUz4t6tFOKZspCDjDJGkf8ua2RTZVHlIHM4X
Ffauq3fuY+V4qdSsoGyvbIbdk7g2OpRM29AR53wgfEHpyFdukeU4UHpi1HDXwl1j
+D11XYwjJa2WPWiK4ho0NpBsaZhhItSwQ7Hr4Ot5qzXVggQovA55aE7yfeU+qvza
TJcPLVnWSn7C9SVADD1ddbeXQ74gHqFZDravzaPrfHHWtXwbJe63Mn9vcsdHW9zz
v6ilVh/bQDT5F0tP5YktYUeuKkKtLZ9uoiGtbY+hkGx+9hMqypBDx6vclv14VY05
cyfTmmwBks4VC1PZz2u11HuAW2uTM3rcfaE9UAXnKHl7bqSPLPFq7S6dL9rJxOp1
ypjgI8d02K6mjPCvNIAFhzPH2qL2TMTWl+KuRoG9gp6svYNSsvBSmjp2yLh7TNzJ
QF0JYDZE8PniUjR5ir4mJomK3AmfKp1tM2EXF93jdRMfw9KrBBkMb6d5wQ3ArejU
nkJQTjQ6J5GiQ+gIYgVGzZfs+fpfOLujjrlRkqQYh+yk9zpdN+9B3xchWHWQGT7F
jAxQWhS3W/cGMoeiIhfsPDtKBHmirl9tr2Uc0DwG4K1M6p6LnGdCsCXo1pCmNXkX
AL0zfRkfxxWkKLIDlNI1+IZBrQAIhGNc28UYzWIY3eA5EazzmNcD/w8q4VIXtuhu
GmRJlmdeEF3xh2qwRoROyCDO9QLFCLBJo/MgtUD6dSRuWXZMYWK+pnSEAvRpOVBP
Yn0rHYHxnveCLPo1bPh04x9zQVJbasw2M1r8DeEskuexbxfDzVAeL12fEadUDlOw
Mj9h7W9qkaBBS+rnoq2w7OeGY6KMS6q6Vcye8SRjsLR+ppYpnR77StJg1wRV3xWD
BvF3LQVK13UWuDibXu5UzOvilwEtwGuFdkiurRbml9jmXCg9qcw4M3iiJb/m27Jn
AtruQDaI9WULtGuJ1tyJXCxT3i2VSkYcmEq1i6G4A6cYUkHr/eOR8Kt/qWozxOBV
tqgdNE7wV5o21Q1fnmLLbW6Taulslcvr/VLwU/gChegLqBkqt7DxipGyv8EdaK6e
YfzSXIIgiXb7Unv2+yOu4AYLLbwQLHg2Dwdq95ErZE5IGV/JPAlYNjltJDXbD/ZO
DfI7vujdZrrGdhsNpOVR2ik3sYrw5Lc/Rs939vl9vJ/x4POehVdtT6rRQP76F92K
Al3tUgsLmEmlRJ12I67JP1rN0F2IRdwj/MN3fU/lgUrcH9C8ohC82URNw2UAIIya
2LbIxUGY/01eLeIme+cBsS83vQmQEK8N0Ij/c+vvJtYIYH+WCstZZFHylJ2pd2UT
8mZeyuW4N7uPYjNPVtIlgprSLWXeWpT4Uic78MjbRqQlJbTkcPIljC4Dw6xWD683
F8FScCzlGwkkzA13IJu1GnMhqbyjCotkKiLwhTgznXmxF3wQFSlSNnbsYsAVzSBT
/kvfw1Rc0LcYJFcZbHwBoc9hWk1M0qjEHouSjzeA+Muc8SMvSexxb1QAOssoaImR
zZrwwFwc/wZNKDznZY+1TjYQ3DAnK4+Q2UqYryQLminyyD9FuH6fKn/EescJLhXN
mMKV0DMRvnzgIFEenq1Z5iuz0+Kgim28+J5SdKW67tzT6iMQF0wFLtY9Afq3Lbo1
cJjuYBhRKg/yGk/xpmDiWOf71xtzF3b4CCscNk8j6HgH3/cME1FnpMr0GOScjbgw
YuNI2qb+OPdeutFSvKSkYJyUvvodF0ZxKCGl8/6NcyzEoRqdm92ftUr/QCH7+jS8
0lvc2VeoynUXHnlulP44KeGdtQNBjnQmQbJhNUEkS3SaAa9tHYM++lYboEQhAJDs
/cVgGErCDFIl2Aovw1oCnpbsvZCRpaGZ3b31C11Rrlty0sHN6mhA3Eea+V7h+7+X
ygZZTGBuFM/3k4Jfu0+fpSqmXazpFFrcN8Mmcgm2l47R45PiCtMgqlrBK7FPV/C5
W9ly5XVnk6wooUXLNzaiWc3I8g0dCiASrF62gYnsvpR8LeJc+1c+4uH5PmuOvYpD
H+LSxUinCoNVBiFquqSZvphbGrqooOqh4bgE/NkR+IdFjBUQi/Ju6OX3kKs5IwGy
vfZjskDNY0/+7U0T3gS06pdn53fd9Bc4cfuPNo1FhGbd5z9t1vnmBQ6rYayVZDdK
JZXcoNm1EL7mOaVvv+Tz4ZSGLLZeCVVuoaJG0Hb/vxmVAA+FsMNhkXmuq6ZKV4W6
CJVexQveNhwtXsAbSHvfSlTwtA2/CRXTTtQFM8FjSW4ffGON7zpiv4YWaCNQuNjt
cotCCLu3EJySofEk+opbpgY7lH/gUbh/Oz4nb1BP3iThIcY7vKyrRa/4iPuwZky7
O2fJZ3+eYHpJfhI8Pq62s3E5ezK8vPbcukOwNal2/jQJpKM45/fNnk+iwCn0h338
eFOZfYF3spwmegE9A78mumyRtYGaTtLgJVxZ21LLCtfhr36jh1wUXXqVsUqPds+o
430j6ny4ETlxR4OciobK4eygQapbOLazg2QhyjcioEQTXI/mfcmLgnEto+UwjB/r
wiwh//EMt0a/BdXXM2NFbIY4XoL/VJy/7kDvVN9mMPlSDRyZNXPm5AmQLPHOuVdB
Jj4gua49ZKGo8RJW8FTIRNDdCorV8ieYm/j2CAAtoGwsH17GhQMGO15FtMNeBz+G
R9LI6ZolTber8JpTjqJAYh0zR5fszZLOT0nR54U8oEEbE96jeAGASCSgrNkDNmWt
5C0/ZDtYEy6MLj5f5ZkOmwA1OMSC1lWluAwYImJzf8AJYRyO6fAAkjLWIRkvmXFL
L+DZQEeyf/pcQ3Ay323a3JSCpdBxNsnVieJRuwgOWFFy8MLnBK4kh4XW5vgzfHjV
vn4oIObpQIsLIgdTB7QnKnJjEnJWX43gKmQEt9bUGhPyDHEuURKxu2sOm0p2ezvk
FR+Hd0Vo7PB9YBtH4Om2ZHXsh5lrfJTuD5wLjhDEMuL4Sb648OVmk4MWxGjiUpHM
p0+/eBwm2lXlDayi4+T7YWk6XnVegqX9bsa9Veij0od/geyAAH9dqGfgEsXPzrWK
pQDFeiFKUlW1H1foeIi9Khkxe27cu2xNL2FeZuZmfJM65ja8qDY+02RSKGQ/85GK
6wCdWlZau+C8JNJRZCIb5cgOK59IIRcYj4+xfKU/Zip9KdDRXuFNwgxUrW+a/S0c
MoTKBkuLvmjM8hvBFiw5bRg/qwPYvtzhFgwGtxAdbdXEkGHVm2rnRGqSL4z/E0nm
pxeQQOt1yLsMZtYLtqEbTQieIVO7MTEToAxS0Nwf9p7pUkSOm858mEJPfkg+Asql
tjLt49VpAQV0GW1f0S3UQKtzVittRslqUUxWbjD/wMUbIRieLerlbv0kNUB3xIw1
YA99iwGZHIEUdrnWHQbZnNTU7Pc24DDUYn2CF4IDAj/BrJitC0jAtcuLNPfikDLR
3ccMtn5n0UClYbHGrskVSw3yZVIgoETQZrD9qC3Sc/D5dqR+PVYtjjTJaBB97IeO
w8bPZY5ZUMVDMq6t3OpP71B02fGpKTR34NfJFHXbe3JgYK1Q76Gflf7b+YMwYtRj
EHZ/bzqSb0gz6o63aokWNOS6K6a8ya66tgIiU1TONTsW2oGHR1pb2tDCQJqI8pCZ
UeSer10ALpJkZ3rl4ZWd3nZaFCxYk6udsuWX6x4/+DhY9ZvrZS8/TqVftfM9gdJo
yWhwn4hmwfxx/frdGO9BuiqQqO+YXczY//WBuP5rpm28YQIMQ6Z0dXcxQsFhh+/j
XY5l55tp6Gpk86ywZdg4iTPfVx5VC0iSAWXIa4J7dXfAgPGsXPHczYOsxcs4FJne
Cw9u0jp04wXMtwEg2z+KL7lSXoOL+A5LmZ0TCeH4A2o0H84Ji0lPA//x2WVCTYAp
Uwe8eD2KKGskCGFArlBhCPn7dqmsfUWCRqLisAWr2p99ftez5McVOYvSSNG0pQFT
EHE5mBg8V0boLvOW6dmpKLToSWTsmr7FwZkdSh8NY9diHj91XdSNfUPdj6i9qyPq
32j3880VV/g0diEckHIJz2KkI9DkBYw6sVXg/qQ5xYcgQPBNf8rI4POMUJXGnTIN
Vyt614GgES72eVx5klSHBUg0Z4G+xgckNjare2vyMDvyDPx6qyz3eAAZmmPY1FNr
Tzr67fMfGv29t41MV3n6WtlmOnnfi3wlTbpHFg2VmYEOCUx+NEWIpafTXtTcYlwd
+Xxzo2jz7T+6L8WbnrUnbUhVGDKQbszcl6zqxvmY+Z8iVhFn9CgKWYomS7vxvGMJ
hZj1ISI2UEivE+VhVPp1ov73ySg1xs7Wdgvb6WkWredkI9NvgoWUG+Cibk8r9oyo
bPAb3zTuY/BSBVTueICxnxnF1bxxCWSZJqM0p31pdv9B62t2q+A1hK39Sc/2WEVM
SdNM8ONpCtvYVLpvYDpWTvuZfQePYTVkARFn+gsaANzvBdnf41XPMWeGDCXzRBYT
NS+zc4KLeYB25Z49du0PDxPZ/vqXBZ00uA1rG4e0N/HTF0gNgNxw4J9+ERNZvdmu
aCbpfjAreZYiWe1nit3lIdMMQDuTW2Z0lrgMtA5A9OBrH5OF/7xXksG+tKRTNacl
k7hibbXcDxt2c/6PMMpYxsRSYqY5W40q4Y9Zis7kyi9hiRa5CzHPKCyxkVACNEE9
74+ubohb3xzGruVMI9YHvI5riVHqzWvvXR5REdYAH5GVgagdyHoL09wcn5jR8OUg
P4lF82rH5A9alEFMnsGKvojoPgq9P2kl7sBy2jLPj/GB3OtuBzS7fuoaNjyTMmC0
HeHLuHuOAoGNGLaTsVNfPmL4LGgwpw9TOblmmKAtxFAkrxFiCMIPhmUrRTcRQMtq
GBolUVB8FXgoLgR1LI0TEAQD3DGkK9HLoiRXYbEgwRaV326AHBBR5Fii2sPDQcOW
T8Vq7gn/iQh5wv1i4jwvozqk2JxOQOKuLjLyFLgy47Hu3JaM5VTlpelCCm2MZDhI
98QUmNNVs3MHC4hlYFfX8aLdhSqbpsY+2I1MDgX3GTHp9ri5b3yeSzcUFYeMkTUJ
gQZIzVQHfFSSXt1dJGqrhXF0DqXDcd/9N2arK0/JNz2gaCTHXteMpN04OCSRjrxY
HBEbUVattUTW0unCFct6t5nvrpQkag1kIRhggJ5BAY2iC9XmtG9ynsDj0+Vm75Ex
qTc6N1sg74pkjOMAnbXFJjRVy20aeW+/00uXmwko7propqX8+70M7q97eNfRBpix
AtzcjY2taUkJz+3c51xD/EUEgqgD/yJoQa2aSApENr8E6ttybnLpJHODFwvuCXT5
Mlx7KjKCtvtVxMOp5kThiEhWRVvuWYrmIz0KsHQjwfrUIH1l15QcqeSoGbahvzXg
YOSkMsUz/xQGX8z9jfdt1Za8V1eh9PxnwQDXMGvoNTw+cNxv1T5wR632xcoW3L/9
6YHPO9FuXskBK/Y0iLEGC0rv58KqnsoLJ87yg26roa7DqLQhdCb6SN3lwev7bw35
NCIN69QxsYn8rYyNjkxr8vmxM4kKVD3R0aNeVy2Jea0591EvZbS/krB2vDbykInT
KNSuTVdfWkWTT/CGTuVmZYJIi9alY4DHuO13dnPH3JVlT6ngToqjRLxglFzuOteE
NZSicMk5mLpWJTAhBn10n4wSIHvieQh9RyV9NWFvpuPXhMemk/RGHMwFkCPO0coX
Pl+0k96rKvScMqS2dxi/VvT53YnLMvsGe6U4abRCFsFDqoqYKdnlxluYip28I0YF
0vxreSzrMz6YT6J1pu0j+u3/x06BpwDJ0ymAS5ZRA/l9Im2XOU2X6ficMlKNcs3e
W813YOQ0sCY0yYDKwGtfEDmylMduffONkzr4rVBlA0hzv9cnErm1kAMcKmurktW7
8nx7gi0Rq2GEZo3e39LxS4MGkKL39831FxnEwiabtdWmAf1GFR0d6P2hMis4vsvN
p7VcyH707oqXuWvjpuGccK+Ks3akvidINRftf7FuPuHE4ih0tpSPdhkrxrqocJ2z
OFO405Mz1nNRBVkAUkBJA/B+E5X+yDExBFwJG6fadgykNEkJmCGquXr1h1W9hwsc
Ssgoge83zb3o9ESsDDAeYsykcVFcrVYU0NZlscL8XT56l6b2qdOROE6MBwleSa6K
OGm5kR5m4jFGn7vFC2qiBXV/WqYch/oefmM84ZLtMhB3Jub4tXKXhDbWAOBtCvWJ
hwyTUHj3WytYLVCpIN6ly31BiUiZcu20cjVEfyv8BL4WbIrA8zvaNyvynXFoodH4
lAVFJ4l9XATw8ttxNmfqe4djygRNfNIFDIgvVarRzCqA5s/twx2NiTpwIyun3sij
GKlrqLkD3KkO4A85k6mNVqzof68f8bTQQSXaby1hj7B5Xsq/+SdP2KkgojoOxeKZ
0K8WFj7bpCpGA9BZL6PTC6HMk0olO4SSPzu6xSP1kdiOZdL1swnI4p8lksIGZK05
9+YUeQWxMt5r+QC2Kq3zkxs3CHGewg0isIBGXzNJzWlvBEQtqTPMvfp3XzGqHLi3
YENRMjLra5J1HqbpV2sv2ri8x5J7mupxg1nEvLffY72BVZVOhs0b9Lb3sN4SbKx3
7aC5SnqZdPCNOZ2mSCDApJMHgzOvzhVFL4VRC3+4u/aZJG5oX6lZZptKO+re3VVL
YdVd7EPD08nEyIyD7dVetfty2w12Xox83klIZIB5Feec3eCvkaiMy65qx6SfyojB
2tpuakw0kfXVb62UGtQEzMCvctHJlyJOxT44akkEoTWEDth7/Wo+MtC2XQU6bLKu
H+VEyLw3kLVer/2p1z4OVV5gtChVtZKOSG2FsqgDp5B9QnMb8d3d/MOEYE+0rYmV
Ip6fU9mx4pFL+vVWJ1LJpGz7Npt4OWhfYNAdAkYlHSSC6xYuZl9TGsXMJTH7rh9E
vZuaXapmde1F7gRsAPK/0DfD2VdjFPcQCw5cJRfP1hN3pJg0knhlALFBBGMJWgHH
RC9fNPPAGBDtoTJoEOD2FVpfavKekKme7b3+EpCdqDTmK+X9SdMEs1xqGW9D1who
Bu/Ks9EnPaLV5lP1SfaF3P9h5nOfRgEmY1hixQQDdpJ+aBqmckP4h7FM25D4Wdcd
/j47PcsqZ+klOCLb86lwb6qpoalULZsmY1hbSYhbdcwaY0I/POBb0tTeFyB6gjQP
J/uPxN4qZSK1gcMNiKcMztRCeKre8LRX/9YWIc9l4975bISAdMw+7kh9lZm3sL4v
6Y4H5fevt27klmfU0C/jIRYL8uU2BaQ3XXoe5npxcxLJ+8YD9P2P8pO3c23pf+3y
tm/qIEGP69ZiWHmKBxroUW2uZMcP3vHz31mlzHhGPEZpjCiCmtZ0nWO1Qy+GPlxG
F9Uve1PItqJeHz2EXfPdHZja4K+fxvR+f8QaNDmHpMrzxvImvJ3/lVVrVRHMGsvw
kdMFsQtWlrX6oFAMo0IZr8GSPA6TKQ8luusHsUU6x7JiZDIN4+EdH+sqftfxCufD
Fw6eijiyM8Nhd3lJUmBSDzipLcIXL6mMXoJinHagjfUdhnVme7+BmN67y8xPWjbv
P1wdhzHwMXBKGmPT3/J2SijsMgoWygbvlfnEUc+EtPC4LtQHt/B9WImPzm2wAjgB
wAAThSIcEdbVLGe2K9EZm2uavhsGKlWRn0Jv02Jr3+je4RHdNxF618GOivnpvCBU
VZ3Zic0M9+WAMB4inmdvH0O+uzt5fJt+AKfLE7L3EDeYAN1G/TO4k1PmRBO9qZiH
3Sdo5Lcx5ikj4LgyS6A9aLpZNJOTYyuApNgx1F/FsQCvOs6LYSPlUAKND6TUFi5O
uDwTSFE601S6TtyorHfu6demm3FAQxONLfUico76h7luIWlpVM0AxJ5galRNPaBw
H4WOwBnr0pTOJR1m+05qfjXbF14hNH2Oiwsgu8Rt4KqsEFNNipa4aZIxylLgFkYs
NEdQuSAwSAOu1T6901NF1SwjGH9/O1fmItRVhtgKyhU3bC7VRJdsrPOejHwQu4lp
7WAQGn5dFxxyc0Xdu0KfiN7xzdIi+D2d3TTbnAC5x1sZsemOs4M7xT7sgsyVs+Ec
tITwSzBiWvwebNZZ4WGbgHYr1MsyM6KHADAdYih0+Ikrcgvf3259ShJ+PQzpaJ54
KwTD5V98CFlf9l1a3V4z8u5CviqT670OC4T+OvsL+370Rl1p84wE2klm/SCwO2Hu
EKUHhfW4XOs/dxC5vfHXE2wzafwO/xvzrl1AmqzvH5AahvrisT/BhdJ6Q9beQdys
F1Vf5A48VwaAdyYc1qoWDAtzYUNwDfkFKIGz8DURs5kw58lroQ3omD9PYiuKeabH
IP7C4HLmAltPItz85qkVA1DNlja0Fvigfyxg9Rn2h11+jMVMjbKNYQHxM9uuvUiS
PThZ8nxyRZ0w1Xpjlf9ZeSRDbD7iJOvfCAAex5OZiVqRpMtciNMtZBNLmvrr+kcM
V8wqCKd71Y/2TgdY4BfeNPSzx22OHGiWE5P7qZBAFl5BwT0/VgUmik5iBl1BPdhK
banC8mIy5mMACgJ8wrdiBB5M5LwjJR10TwkU7KC9h65YQIOd7/PtsDtt95HR6MQG
b6NatJULjgAfDYPQo3UjhfZeysGUSD/pNX/WHadFTSGym3jxLPP+GZ+IdI5sTxau
8+I+UKik47lY2JPpFY0mNj6WS+tVu6Y8uLRV47e/IXczG2FEqjqYRlw3U096kQ9W
VNwg2sR9jT3/ktLDbAg5SGPJM0R6tb7JMbWidDKOLK1tR2Lra1zxYfHSO/s2jeUa
72S6B1xRS4Y5svKIblWCfnnZJ5sV6iE+oiaRIQ5E/aU+P4am5BbjVuUMqQjIDug3
0JLKQcXBbEkDB0kOFfPBPervF+CWqo7cvM5Wtia9PTIbDl1m2hQKplr70dTu5Wbz
w2ueF4ldzOz6zol1qWw8LNSxAz2ivdhAQwGlrrv7eN0WDZkhg44/pj1Bx7nF39Ae
I1I0USHa5YgdJRZNQu2bvNeEe1kwor9CwPskRwM2cJBipsqKGM7316PO90BUY9NC
Zvib9KY4HuNoqHwYNIsGpViiwnrZQGqPhv0BMQta3JiWICoZmZ9sLkEa63vNx/2m
HO2VFXjeWRlg0y2GZn+ir7OCxNzJU8xBPeIv0QYAVEDESjyzB1N3LU1wSY7Cuhsa
HHDI4uSBb1CNd3JPLQyfda0u8uR8NcdSWjL8kQz49mG1jnx5g/0tq5Qib4sqMx89
DT9r1naJRragBhQlRk7//R8VeEI+9acOim5JvZ3kS1qsr3EBaj4Mi7BzOUWaWJtx
5wkpk4YfCTzzrqHAP8dLqNulV1hNxPLBR63n1AJW4+VR8B1n3BchJTOX/4tVdCj/
trUSeCHi1a+M09s/hP2OnNEDyTCyQTM9tOFBXvqCnnyPE8XWn99ZN8CaqBV2Mgwl
LmF77sJ6v1CY10C+0vKkYs+Lpiqxu6vboraJUEpOyf+ZJtHG6qBbUgcAX+IcSFkR
zYfl584IU406pbXh5IpQwc7WrHlOVrztLsA7/QelhLo089KKsR/jveo70smb2MG1
tDTwGtsvu3lDnJLMMglJODegwATzPiGKiClH4pJxUJpPsi7PYLBfNAxqJ7fr9qTN
5njkeIdhgP9Pkc0R0QoGMnv5TDO1SAld+CMP+r61F+IU22nDJcap7A25YjqxIC4H
TjQTeN/DL59gMHm8JsIovVQiw5SNBZqynBBWiV177J34Chitd0RJmCjCBfrI1yU+
4IJfkz225yz1tqwMnNtZxk6p8wqDqypjTeJb2ZBNWKhG4q3zgDY69vMjEnxdw4Xx
WCuWMtJy12NS2aSK86PVcgwdPPePWXOl4mFJ50naJgEzF74j+HuXbiLBF7pWkbf7
h+Hw1lSUucLRR6GRDkXmNoe/t5wCbCLPjytmP32ewPHiTzuj1/CdmPt+9e/8lpM/
Di1xoRKO11hM1PGhYvwmV+n1D8OBUpjt6YI7BiPsJZ9ngwPY4TkBZK3DCluvP0Ed
+JqRpfmN0Rkoj3YY1VFUGp9Kg+4ERrAZCxuvsTS/FUj+GEQMm7BivpM3EwGK28ph
iDRCfAz1z4gSaO8HEJuMxhIc8FjR/a6yT/+bk9BopKyYmd/BN940feD36EoHEYef
cTts2lxEZtLDYfCXOt/5Eqk4vyoig4Bl0ODZIhINAS/tUdYqCNlRyi9m7cvFgVeW
a+PMc5GsfZ1XubHwvALhCkXP5SJk9cbZU2emQoNnLTPJ7OvDicdnlX28j0W33mFA
DGmciQ8YT+vWGDv7NNd7vWYixyWKyZGxxZCqiC2zri9WASEwB+R/pqw8wnq6NIcM
s12Z7gRjjv9ASgmDIDdNN8//2T6LqqEinklXgUV3dRrVbvKWjdFDq2uJwKReCp8B
qtdt4+zRxPLwa/mXo6wl6x5Cbdv3J6Bh/zol+ReaUzaYsjakMf7Ao3lMUGPWNmp6
WqLjdApn92P56g4YVi7oDCW0CCrxXbmUrMBZuYK9HGWctQUtmVjMhiGD8SwxOhWm
SPunlLOgdFX2F/S0Ljv8sddzOe7nZt8+f38NlCSQ9B4DszMkSW6Ts821oNZV0e8E
dkP+hc+RrS2NbrUonU9xpZI5uUlplc/HrdQOORGB5OqFzjmgcF4of13K6srE3l1Y
c9TGF1XmePWciMtQVJIlEXrLoAIKlLwgRMhH8kiSGw7zzMYWaHeT9TzWBQ/s4YqF
u4ttxs107kg/zzH1KCy0ntbZABntHiuRcpgY+PDwiSkYLB9QxO+sxtu+xZkAJpcq
C2thzP/6hy0d/MQY8Lo+7vm76loWmxPTFk7JST/5JO0BtPiPFeDDfKRow5/BqkK3
0zHH20Jqm9h2CF40bHD6AuRlXFTSVaT6gg4kskBXurGFp5L4JVkTlcSTKh8+auTq
WSrtQIWEGA3QHbsF4YziQLzNKWMsz+xXlkZGU5RwJXTgT8K+Wc/FWN20OndZt2av
Skvf9Sf5GqzsmEYNQCC5D/8oBnppjRNAU5wLeHJcMSVHkbePrRyrrlrAoyvZNpsc
C6brLENxGeH9Pv9wXnEYOvk/BLf+1R6Ntg2TiljhyjL7TSe0avlFh0h4NlNLN6dC
82sXCe46t4yCDsE4Rychiw0VzAV+OnjHIOLF/wAr3jo/KfVKzlLo34Oqf7ZZHSUC
2tcylup0ICyMBmGMub0KofB/MuKtndPkZtONuUkR49tTlPk3PavkJCvku57YLz4O
4efdj7q+NQctKkyUI9HM7cD2fgyvDoyCbj7raCgzFTZZn6ZM5w/+whm8R7Em9nwK
CL4JSHS/zGWh4h3nvpaydn85mGOPgP8oa8U75LKq7GDhW+LtEjRCKTec/N/yKI/8
YTREzdX9zqFAYiqL5BQ/E1PGOwkZXd36V2b5tE+cdSGbl/4rcwLosZ5YK3ezbXCg
e1t3nRA6k2eGmUYcwgefKH18x2HY/sTubHNmyzTG4AMo+sMkEFlGVvOBBcpjTIY3
0rb8uC8p9VqKiLIfM9A4EaC2tfJB7JG2xVXcOK2SgATalpjE28NordFPwCGIW1gC
2X5Ls1jGHN+CqGza2LXu4R3D0avUuiOacqWNYRMNOlFO/ers1QtaOJliD6UvxP9X
9FH5/cas3zHHFVCV5+IKyGJExC58/4i3NH1yDKyacCIGkfU0M35OddjKo3W6vEYW
bt6wYf9SFQl+bRBcqbfN7480mG+UlZyjqPajCzpZGj3S1Qpezbh5WRIzgJzFjONl
1CMHbWmkJ05AzVEWR/gS9oXoXkOCBqQnKSUC0LQzYf9GMpTRMqgMF498yMEjAC2l
D2/OKsKq5QtvMHDuC87vuGp0HoTHsoCKalA4TsStnieyB6J7F5QgfheWEINH3UO+
njGxGjkNGImeTZmxAyZseyL/RDorxj2srTSJzlLXhoxO1fB5oEt1O0aYLuckDOqH
rumNgcYL4GLX2bpx66aqHlKTk966ApLXpTYb/84E/Z0WxH0TGf3YT866rMEm16Qy
625DIOPjJ1HM0x1LIeQLMp3abLBPQqidmi0dRUlhkojT01R6vUIedTxtigDT3vPn
2ehXC52Nt0klbNEGzT7nM4c1U1wR0RNtOvjyqtQWkUO/NvZxNKIDA9867ev14Gw1
aqNcViJA9SIQwQ9IP+fb7f9EzJ6NpoTWshgUdcnq1bc7G+LiJd279FUNgX780AKI
SqRxlM+0bOlY6b/wmLfq82oUEaamIopcTJPWLJb6qixRBUWGeeWbxBE/HgXY8rFE
m0OguXbB0fKUo4GOyAlNqy+K/uIGfclgU5l+7MUM3l8B+iG51qJ6uhHipcftlyep
7tRMqQY7F8+4vykcv5VfCTcaGSFP1VZPM2wQBpJxeNAbNUYHKDk6YUIt6VlpM9gP
087ZwFwwNIc2Gx034QIFpPEj0q8DmVdFDIGbdN2MWU7BQ3gvuMDe4A3cVhE1lWLe
cVemwHZmbD0XIz9TC0+xlmD9q4xAzvEjjI/7gCVD7rwuub/TUtPORJ5LOcw+8IdH
X6XMneiW4lEw6NoDiA0HcP40COSNdYBJBsnE6PbDojg2DM/Zed2e9lHkRNgT7MRV
vqGljVMpVJjgT2gN5NPThxwRkO4lZb1K6uw0hG4YL3kR7I2P1h6Xvi9BtRxCxJp3
ZkUiLas2Ij5WY7vuNV4sinAWvn8zzbiPZv5jRDZfFWf71DAkPZ/96G2LwDh+U6kC
e9+N8fVpZ9QjZr7bkViEDR+XdRv7szrrMU8r7qy40vMfZrYqRqfzmhb9w2YMlkmM
PdDeEvCJBpcLscb5uOFbeQ8FxLKNuE+bv6jxdzQifiDb3Ns2r1upZfE4T+u4LIGZ
QXYCIyp378oGXSA93A6ZuFt4FIhjrYVp69YYiWCvDkshylxp+nGaXIYjjBz4T3oQ
DqovszIKgsVLGAYnDz4qPKw9GSw6V6/JM81NdaXJQkeXv0UAhpp7jEdUpCqGkbZ8
t6HcKRyqdXLAmy8uUIFqvERzFlp9U/fA5xZyZzvMZOPgx4y+0OqauzfMGhMO+AKg
GGwuGRIQyjWhL75KPk0ykZ01pD2Sh+B0EZpg4jvEdaZg6Zkej072Px9IEKUtLaYi
TBavM9FwNYw8RbOJR136JljpuCmWEj/HXSWdQdfN7TNcKsAEiLhKuh9nmUyuFkYF
r1ugFA/i5NMyNovDcgVsv0GTCphTuleOAqf4LQaFirHH7RtaVO9jGhjV4g774ZeU
Pz99yH/mB+TgBuVMkfIfAafloDbp+26UW/N7UVnre60m0xtbmRITamIP1+KVY3PE
j7rDLYJ1icfAUJYhQFUuMzDH3Cei8IOGAtpJ7424shur4RzInp9aNL+hM+9ldUJf
FSUZAXOoZxOsQutIlB2sWdrwbaAmBDHvm76cqRxGDlj/LORtZMHVCq8LJkTCRwsJ
ZadmIVKg7pB5dZTG3gyobV8icwuN4EMFMtxyNI8RBUxlOLn3U7hJXD/VjnT1nF64
gL4DaS19sLWwCv/A7qaguiOnvsZZww0aWMN9R0shMuTxWWzF8Dwxq2goeno8ykRb
Cuz18zzrgT7YF0LFxjsd3VEdOxlPIUFMGf8gpQQwRA4n5TAJX0IW3KRJBmdsXYR2
q9AyITW1LzYM5brL/D6YNKNF5UYadQD5rTJ3II6s09G6IWoAmUz5LRyX1Cxk1z9U
2fWaBkfI1ASfbcbiAlkpJIlLL+em1BBNiZCwJyjxekYFKWgqWd0noRaH1FMg9kJj
t0d+5Yq9fVy9/I+9FGeqTZgcFLsrmwnsVaAHkH7BG1XyR3MOVnL3KYS9TYq6MOKp
AWpnJFGHBtOmysqVsgx+1CQs1t9C8GolR4V/PGQHFBAkJ22IFFkdUFnG0tvgsZZr
tX9nVkBoII93ThfKHL4bR0LGd9T0lCY7STz3ERIEECMv1d7pZsrkq/8pmVah/rgS
DjLUEtglVHaUSJ91oAs8iMpP54dYoDoKs+YMM8CSrjczainD91PGKniVcaKDcEyj
jWuPu0FnZoO75P+3bNDuuYyfohQXDJXL8AjFQ0LYNDvnsQZ67PDas3WXWFPgf4YM
dvHVcRVxWkvwX4pbQI0AeY7w/WY2dUkhQ1BmarlEuPPK81fd4Kj41m9+/1CqxJIr
Z7mcoo1groXVDF5RN37cxX4EUlpY3x0Rmlmfs/q+GW1Y/kL2B1ac2+zmMoAQVFxi
ca4NCDBdHhzcoYUTF8bxFyl8JDQoPNPjHrl9++Hbv4JINiet5nCzZ5fUq8GKPmkD
iktNo5Ot4+Kx/HZEU6o6vxDhKmO+M7EPmnLu4bhYLnjm4bwyKexpOM9joDNrpilv
d7kA1ccHjs5tA3N+TxKFdDhTsxPeMc28lTu2B5zaNG/R/1HmYKrKg5lYuAbChjVJ
GIOVBxSx4ltxGPdgwNEVizCKGBw0+xQkFCH8t84mHi9XiPDfNLicyxmtmbsHDayh
MlGs/bxmQNIJAJKaNrt1W1qnJZDH+ZYfU77D7igm09+2z3h/pdyHCn/aRHntk/fN
L1socQ91PiCITKUPK/C6RdrwUlQeKlQGxxCnwN7kCCu/OzXi4/64w1ZXsm/zirH/
t1S3euESYY1vJQSEh/guGyjDb2pfeVTGKhKkge4o3Xp56rNOhPSZC2Hq1e4c0mcp
Ixcl7F3Seq+Vu6z5q4bzplxjWlsoxYs37fem9a15bkp7eQQlywDtO3A3EgNBzCZR
6AnPKkRlaBkaNqDiSh7DBe5cdmfPSlnaeAUsB5gicOsRhYgG98w2H8Eu2RuVnC2A
rbdtMRLdGuenW/5Zne3K93zRJ5jFSvXWgbI2WX1PSiQa95ivfdcZsWmw9OXfQ3Hz
+brPeJrtVIHsuxZ5Mu8dyKwoiXlU2E2djlmwdLInNSFxT+JiJKFbgQeamkmAnoKx
Db1zdW2TjvsC/WDgvnmNTNr8/bSPNonU0ZpCSa5hAu98Sgk3Q0hgaanqIRYyFcKF
sWm8Zq8eJ7f1nCijIZucVEF6R2+nnwOBdPMxhvalW1KWKFD1Jw0+KE+QOaXLj3L2
YCeg1FwLPHNhiXp6m4rZc8NoPrq6p3rmR2d+NpsgcuCelK4vBXrCM4pqZXTJfk5w
RA6jq49/gpKWwYl/SXvB9lc3CjlKSYXtGp60j4oppoq1I0uQJl631yh57dL3So68
/RGupA2QdglEfN81J0+deoRiY+wfkwROwTpt26VmA88HPBWDRMWTJ5sGmIjwIC0B
S/AMx7d/NgSYkw4orRZa+GDnzTfW+r/RGyQFU/A7i1BqQJr11b3kakiY+ITT5X48
QBaWH7z+WPcuSSsCNsKgvzBariptvUFEc4maMF/zdhkQFHxReg+YLJoPIkQO1Zce
0iuNGzuEj52IHgp6zZ1DrhymooKQS62UTNeJTcUD84Pmmu+clLFhxy20rJfjEkEG
BMNQb8SgIDyuxA1PmjCBEoUvA7YivfetKOTuDfXSnzI/1WgaIF8ltl0a276nUXsD
s0etNOhUCc1inT7hkCHWM36SwD0htFaEr7yWKkPH4H6NU+6wc1SubB8AbkciiaLO
K4RiTOH9Byjn+jwW9ChwAgf4Yj3PPtztn/BDZoQTjZ5YH6KavfhbpI03PasL+2U4
vc1wphKrnb0/CxmzRMvgqUcKVNTa5W3ZjAQagm+qQ38Oekk8M4gwEhb4g5fVDYea
LNeBmmbJP7mceMMuvPY6HWJU3eznzRu/BeydlndYnagIZ7XaualKL+NvuH9q7Z6f
LvXyTFtx4YoqL8kNHXLR6XQEW97X7Qh+VE0u54iJuXKtx6dPvQOOivGPyaso4fqn
stmm0wnHTyYVbhMKqj4suHuqMrlyxggglyKzU08QLK9HSdTzCToIjnRVY5SgpDRe
m+tZR14Sums7HhMVH1b056aOtwPiS1xWYLzSLEnu8eehxOteOrw/O6v6NuQNFrqC
eSqNv0h0JamkuG+fIUZPJFORv/lpoDR+h1XE52lPIwCYfx4E83zL2wSelPK8+1Sw
e6hj7/d3vRQU5y+V2443njNifjZN6tfcq4rKkmfrxrUrmTN4bqoT+yDdSHkFhhb1
l3Yq2lA38rfbdBrOgMQBF/JbIRcwpQ1WIvfye9tg247E7Z0sq+rRV2iXNFvDN29L
adCdbMCpWo66tOJgM5jPLlUscMt2xeqjahWFfd4mXJ3Om1oMPoRmnqzva2oxbfUN
LBR02BrjDiVDZOEWBEuP1kORFC6+BdFzDRv/MwzWswLqK+4B7A+nySrPhdCYxU4Y
jUtMjV8QehFIukhGjLPl7ml0wprlNWiRV8WkvE7PvHl7O4ieTZH6n9fefJ+2k01y
4QI3LddPQYJ670Kded5p0JaGMTPvBev6TyY17rTSEieeFyASuu6zuLGtx2AqJ0y7
+q6JJZoSxvJiq1/semVTta5dLyFL81IqKFeuoWhbSRxlMbmcml0uuuFul5S202QB
PG5fEvFTNvVwOn/ftxbnY7v6DxCt2l2HXr30pN/IurHasLPz6xayXJoTec3Rsv58
eGieTkJkEeDVsOTCttcyV1e+5z6CtyuXY50kaiGEasNZtzRIQ5pYe2Vu6rhKqj1x
6yfDd9KXOnzZVuGwtV9sFv8lJEH7w4EeSJotn33jUbCLJlVk69A9//LJJ2hpDag2
wyKC/6SAIYUKGA8S4VEVJ8uQ4Ovn6KRRn0n9UPi0P5LN4uYSSYkbdgwAtLrcGngC
pRwEDQC4PtqxlY5VJm9Mgh8tpVGqYNqVhoBIpbv11PH3kTAJZ1T7AMNgCVVEOqpP
qxAoz71GBnp5lJQAUtMZs1rseqep462uRrjqk/UqO0zx0HVoKUFF9HN6oQQmbORM
90E3QugzSCuGW//qsrnbr+PgIjamuGKmELAuPBjM6LZR3jabwmkYecQoQ97TLnZc
S4WG4H2qFnbiR1DOw96RdkB7fsnU8zY15tMay61yZD8dZNwtoEm19suQu7uEpAID
MUm3OGj+Lh21ToMlkLAo9/isqbV+eMTDVxTLdhHnUfOoq4M+qdJR5+tOoMsil+qJ
vfBl32tdhPWYN9D0qRxJhSasGnNeCqIYggYNNBFT/2H4s8gEg0gN9Cg9KT2Kdwow
uKHDXX4N9pOjq+wV4hcQ/vEuoWkq7W/mUyIRI0lV5FBJnb2fo8a+UtfU/RasPMX0
epUcSQlXRBvctxyug6hlvDFAB2CdAGDxetigGqymuHrFQQ0LFRhjNJ/1Wg0hYR3R
E+lx7oj9qnOlmU4joDCqSwDqGrg8bRaYx/5eQRzFe3/sN4Ie69wi+++mDbaLsJT8
4qQbhVVS/9Kwx4AM1vQtgJbgGXErPV97vGtb1UFP42hTZo58nY0crN6+B8K/JSqO
Ts4SlwuzOhl1Sm6GHYxIracI8BIwdPzF/teXaeHAG+xqt4tk5GgQTgmU6jxGDPxh
AJL0AtHlyxlnQsKlHQra96YyRIvw6kVmAgp2y+aYiX4iImzH9h+CBxROXPsCvrQk
CzyOL9jG8ivUaw43GGmeblhen9OU973HOnA7OEKx53C+bP+xj6gfT4mbSE0A7jBy
ddZtanm+H64ivZ9bZWaEsDFHwzM3CQXcnGgx2rnJ/jMFqO5rSiJLSIs7xcRuh7nd
7XqtU5QB3nl84C809tU+S+Ax/pMczYRK7c0CIxxkGv/DDkSIA80+BYxk3MQaugay
vzaKe/KzcefYiwRV8gmyKnHzza0SxmhQlQmwPxxu7zz/QaSkW1NOvSh9EekIRveQ
GEiMJ1BlZ2tgvtrn6L/YMM7yXZV9N65GCp4JdIXbrION3Csa9f0d5cY+LFAHUo4h
D/rhbxp3MxCAHZK5GR58tg/fedVIShPKUWfSsYbqHqs0uinSI9N3OOdxhebBfEJb
kPI0ZOY9bXGHg2JLwe0m3VYCOeHfT/2KamZGEZlVviapRrQFdvZ3bGVibhV9MO/p
nha5u1FBUSN1xeCVH5yj+CS+OAvrmT3pZWEulCggOrjstlaFduojRMPnsbOs9Vsz
ZVrWqBvgPWuRSPN7hXDyecKpaH5b5JTQDNmopSZiY3l2uAz0QTWkckESDj6Bplso
fr4OiK7iDgHGV+hqVIyKOA3YPgQDZMEEEWAIJYY3tnHLBuMyqj48oHt+wf3pfQ9M
Ab86wmxD8CVtfTUy8Tu85Ja8/ImaTJFTxJzgv0qPfIOJ5gU3KFWnDDt+LpmxX7NH
UiPuCbjHndbWUaHcQxrp7vVTigRBy8ManJIoIE7Wtb+EFMWTB72W4Bg+JmHaNHYy
arJjPDUe9eE3yJP0iIrP45lOGdg0PGyPnY0zA+GuQ8oURNzFs2KyC9BKlP2J+FaM
ZmLeXMpkqHsWZptrA2rlb07ugpuGDB7DrbBYOSWb6pfSowtX+3k84uzGammvMK9f
SssYIeRlWz7nzUv4UptaoD/4jJbJ58TmeaKlIYVTHNqoP7Z4PbDT3ZUlEDJ/WJ3p
iacb2DII087Wqx0QXNc92xzkj/dJvUnZBqYZ197Igfsk2BzR+C5IbvXXwlnDMM+S
nkX6ZzvFeuffSAjMXmizdaU+PqAPFID04xikL+CA1EeC63W8z/QAqHZIWv0xGAZF
dLpzCOwb9QKY1nWNJ08EQWuQNBrv28HVRXa4C2a7wdj2yYoIVQKcI/QuFBOULgv4
NtBA9i7Yvu5qNDNT3ldRgi0GAaD5+UuRbLMMYUmpDdYz3IKPNxfANrmrOEL6BxkP
4l+HPo/tv5QijeCAOgWjyYnkvMzA9dUd1KrmSWMqUyFKgwf1xNTpcUsjxSyJyx2Y
Ie5Aed65nRwhHTAh4SFrx193qi5Nkp2oZidTqhbJZ9l7BbyA4xf3jhoPnkLRpieC
gijQTauxtSY6UmasXtQirANF2TDIknVkEjLJKbBg/4oFbGSeRdUFU154zE/lcrqp
myAafz2BphB0NybuG3zZPyyXvzROwsvAGw59klCntzICR2Aj4S4BlJyKAsaTmAQC
z9OS64FcYROB/GjyVyw9x0uwjjEeiEiMRRGE3V27e4ZzPpm6ebWF6u8qI+XIBw5x
yG1Ax+EZxVSafXNjd6jZJvDAtmjwEkU6mgwL4/37o0PoYgtpSn9bSzx8OfVM+lzb
OFDQHraQFzUsS0u6a9x5KPuPcQidVfbYlX4AJ6R1WRBbCZOHJqrSmJSkZLjpbAPE
vbVyMkgSau9tMXKkzlTz2E/Fv55nYFWsYYi2jpQUu2FCYNeWHJhh9e8aA8cznFuY
tItTrezKbYPVMpgHA6UO2jla7+cpzd0a5geuEivAowAguwmC/aCeoVLWkRS1NQaL
DyQDNtxpW1IYcyxnHFxXHohfYuHNXMR792xVPuFjSbw9lBr3muscm2UUyDnMbKlf
vx4+2ScfepYtzklvPX45avi4JNk63tJZAGZ/AennwRho3zCndAWQdjE28TvIPFqz
TmsuQvJE91QOt7YohfkCI+AHP59qQMWgpx35/QDoOxViHcBxDbtD1Jx81Uw3YLv/
M80q6YfjJucRv2yvFvqDg6r2WYOSL8Kd4XJFrzAaAQPXMJz06o1uFnV6FBNbh3IR
HYCDboSeNClkCdpswABJiITQvYYi0Cvx6ls4Plkr+45Ogu1arzQTSEkV7btFwNfW
4dc/CznyzQ0B7+z/BqR7W//qFZCjtGoK2Z0Swoopirr1FzWzBj76jh293wR7gVGW
rYHA0WA7WX2KpI2r6l8KYh72r9+ZoYNfRv2eYoGfroqisYJL97rb0zYLODOZG0Kr
2afOa5rXPJ/yfrwHbUABixtIwJ8OnYN5L/wkoDtOo9AZBV+LY1ZkbeODTXTbwr3X
H+VLIrl90MIAHMN/bwEcdiPZnD2BZCanouzwuf2sEQpQSP3tCluxgu6BgJi6KgLe
oa80IjTtAzzM/tWS7acaSAm+RACMnN2uDEcUW5Y3Q8hW8eq6YvI9XyFIkQTcwdDa
dFbuH4iyO0GKCgCYATAcmg85if1k0qsWJ9fYbnPFnfIYtiIkH6N4CkDM5enGSKMM
pJ+3uf3UAnLfbPUnKciJEVq4hheDnob4D3NmAxFFGV08g8OzIDL40lIlPYudZVtZ
nznv5UJMnocaPQlT2ycFZhfLmErPH3LrmrhjtgKsDgR6j2s6tDy7v66rFLO1+tcA
hbrmxe4Oa1o9fNyDQ+u3lc1B5ttrrIP/1xWo+Ldd3Mf06r8gbfpJA0pdRuACWkJw
xEqUadxWogKCsZoscRVevhc7CCm3gk4lK4f/NdCnd8PpObfuCMJxB8f6y3PFE89V
xNPbxWOvuY5eHNJTPjpMra1iGKsY9WuphVuWJBJPhTAYhDmqlaZ/LgEAbnU+qi9y
Id8KNNXzD749jkT8C5ifnWdg1dz3EhXAX47kLk31RJYvm0SdikHYQWyglLksFVs/
oBMkPHxww97CfZGMgNBj5SLTRHY/BH8WQK178WR8LT58bQyIwEtg5v+n2A6v9RBz
hy5topD7GPTpijwn62qfC43HmvnjqJikGZgi0n1kUnu3dn+D1nIAvODCa4kJnzqt
ckp5hCQYbsjPQzKmhX1IJ4b5HuKove91HiBuLxUWorHaDgWpcU/cvFNxrqlQQI27
Duh3jQliBNVpJjupWnj+t3qqJWklEsSSYVjdv0MymIRFmWgHyFUM7jjcXgOQh6U1
44eSRFadeTFVM8dfVZqsTqS8iVdcwxjXRwucAWsUfU0ZU6Ze9nF4Tc0xHhCEQx+i
puf6XTT5zf09zQpqdLuoiv59X/ouBqdaaddaiGl7iW4/ktZfuQv9GJzI+7xorWOO
q+uC+NaFLn4UzwPgZA/f9Wv0c+fhX7Y9MRO3XVFDwqXXqGvY63WnjCYjgQDIpvYz
wWJBqmFA6hpTjKA0hHWGJ1iTFSSn+jTbQrdf1fhoE4oRB4RAQA134z3gqnyqArFf
WMNcTzihXmFscfj7y4N14RPynqhkYXxHjpztbxnOMGaPiXpJARrGrXaIRiL9SKJz
ILiCNOpcdeCXpUsWrJd0A45IAx1n++f7Zk2+SxedGXAvTTppvpY5vWBFDe9oJUhI
Jn7bxKjrj3my9oMO1s5jx0IdiJIrcha3mwh5x9kaAEB2Qgc4Wbny7wDtGaBiGPVC
Q+FkTwKOW6kDfAvFnI+4VcY87OSY+0sJjdxnvhschYFmTKuhyv4oOanMcNkytXAn
LYfaW+J36olQgfaizTWSt02nFBjXn0b5EjNt8lepkbrhn5Qo1c6+edd/OKbE0P/V
9aNtiQoRSFA8r9znZaShYTf+c47OFmfz93Odft1Eo6keu5Irb1ZBNV4u6P0mVbVt
ssWr2JqchugH7yObeZ4vfoPMvkUjVfFlyXLy6GzRSuShpVtuzg7gBZxe8TLigoeU
6AFVgGoRK7zzP4K//vI6NWaa0pKzmP7DL/9rtA9OiKySJxfQ+0Kqyk1Gwj/o9ZhA
U3svqc8WohVDZfThwf5AA2Krm7o2hfP9WPCflekNFuxZwZvtYaa+JnknXV0uax1m
Vb3IrjnsnesGyQ0U8MoVGovHTahe9FN5RYHp2dLo29NYT1AIXIAgyusWxDnyL2x0
p6THfGG/LvlHmoOgcRqSYq5vyYFsvyfOV0anCiVLk0SO826phS8Ny4Y1KBlHaoQS
ZjHIkMfuEm1qlXH0nKihzmhEq7CTLpHrQ5+5yo/+HccNlrm6ON2Lm0dvR7XdIauG
POcgmfdTqyKU47LCEHrHx7mHzgdASLPgoukxNnJgpTVtTdmTUmPlNm0IC+xxBcJ5
NKM6AGP9odhYqFa3EMz1lc3JDZaZdbIt5ZvyKJnIf7VIDClRxsgwCfVqoiIWMU9o
4HDgmqd7d6oF111JE+X00utHZnnkdvBLkZPuZIXwaFFuGCwlLrk1KnMLjI/gH5CC
7MeSW+loQ0wZ/9UauL/3EYixUHbwMuUrJklnXuZz9I/n5dknM0sU77fEXJ1t/6s1
4aS2373VP5QtWKQ2YkaYobFJkqwiZPLzXVd5IC9N7AiJ8i0gyHGBXWpzqgiqs1jF
2wUotfNqsy0S2GZYfhIih9Y/aiMPZSmZ9a6V0AuT79x/7pt6APVVXOH1biNCcdvB
VJjyI2QnYoDA1rd3qPt6crv/ZDk7jjKzvZ9G4LtmFTy7HY99HikVBjZSQVxFxfIa
G3xjbR5ZVYs3cmJJTntGpzNlfaX4BgAFZK2dRNq9+DJ/jADvRkw1vjOuzfRG13C6
hPOzVwDXXEz7r3HEdUsNByfrGOdB6gdfFT5PXOsuWX4bZmgvMYSdic4Uy8qlVJjN
SRoXaH6D0TDHwMH6J6wKlnoRxr1M4Wys+VVyuh7zV2cJgqawFvWXG/R3SfXKQ9tK
qw7rU80/Wcgk9czEETp/rGsK3Ku18jFLvnjzInJV89PARZ5UL9WinD+/5LGY1aA3
AVruW+2oQWX7qAbq4LYnz3/RmVo8marJTmBh+YwTiR10pwSfI72xj6eu1tRamldK
Kmu/rKjn/VH8Y1iVMe6QWkWp51QSGfYo7AGtD+O/pRmOy1F8e/+B3vtuhvHoGG52
xz9g8n6qmVnes8boVptRvxoZ/E/L/u2jz5xJsL1UXdn9J/UJ+7Pwze/vdN1Ho6ES
o/djVYr+/GTkSas3pmLXYR6SXuHHwli6cSczIkOZbX+ehjVEltQkU/GxUlw8Dho9
h9fWcxCnW5x3lUp1hwPyuiHvUE+E2zW45e5l3z09qf8JsOvyZaoRbXBTxoKT1W5L
pzpfO+7ccozgDuGaKWYRHoo+QkExc3Sbe3U7G7aot/l/PA+EipVIw1l83Sy3a0oh
UrRg8ckaNGq27Lq36cEAnMbsm4QpM5S3dOgJX6x+vSuF//o1Ga7+nkwdSvCqNn0o
lU3BB/qCAK5GhSeoh+mx+JryvkTKvj/L5v+yEZ+HzbB4ZjeC7HrAZzIJxjEwQOEu
X5Wd8T2eU0hVePWq6y5nwyFBJy3MkAz9NKp7HBG0I/8341dt3npqY+zHMjNuByI2
Nk7fanTHsvKx5GXRiLrxVOV79bxRCHYwFCPh9iFBsCMwnNWldKSZNLYyZPaHW9/G
2znBgL2MWjMpw3PBtSwve4dlGezguy2X0twNVl8ix0zxXKaLqLjjuIVCdYrZwYE2
jU9/aQ6+RrJsFV6DE+LtX10ducKsGLST7d8Iya8n7zjbdhetqvRdd19KD6j9UhGp
zX3MOwABSaeO8FFXLRwcukNf2Ca1ptU8f2sE+LPnvul+ljb/VqL75gghi76guXxH
uViStNhprwTBJJ4A7vPOt0Elaio7m/aubk86MJmvoHpX15yWvbQAhZ2cyZXL9Y+5
cVcs06PfInDj6Un7X1NkozJ3dHf16uaGYzto8Sh8g0PkYpb48zgYv21AcVphiihl
MS4TfM0KDTSqP3ksycLJJ5o2CPVh4Gm7GGNC5s80zkcunSWBpZeNpJ6QAIq/Clwi
GznuLiDeWUn+2kxSSDpsVDYk2t3wvojO2645enpab20fbFU7urM3IaIZuUQjtMiY
y6DIlt6Sd3vt2GGNpjqoi+Vky5ka5u28Oqh5zyOZN+xtjZTjQu0EncmVNggwAKQ4
Oh1wbSe4WV3BfUwqy5J8LuzTJcLD3v2FHq01k/0ErxF8VYOaWGv4i9MgCofcgK1b
cO9Mx4U+fn07NWBUe+ddVm+flxXS+2SEz0PikSKa33DxKQyYyp4H5cSSWaWU0y9Z
lMDZVATpxGM6GAkpAUmfK9Qy9v0EbmJCU6Hx/MlTs+6lk7BUsfqX5AHpWPvwHOpv
WN+LZHe7JrU++65QFF+PKIeqgwBTjMUZm3kbBrByhUV9UESuRmyDlGHzdmoCZnlR
VbE7dOAN9Qn2XKO6zfk8guCFvq2MAEiTw9nhOMDmviNVup9maJCZfieLimdMD5P0
FtfEO2s9jJEqazvxfY4jdArB9hPx54Me79HCqFJmwZhqn/PzldPHW6ep1kMYWAFn
RdomAQNJ/ybsna8/R8CmlVbK1oIZ07VysFlHfO95kpSmMv4QPDh2a75xrrOoxDaK
Y9vwww1rhPFecm4xt73n8bq7qrsiPBUSG1E1CY+Sc8EUdox5H4w8nGFP2kQPALpd
ECKb8b8PhPqztxLXLodCQ6mul/hxAuQE2VrH+lfMt/HM7XflqR1aLgw2KMcGHYnT
GydD5QmqfPxAVK2h32nxsoSw/adNM5Yqg2bnWIqt+ka3Flzar6nRvBVarEOa1pfE
0JOnu1db95vlacOE+ASY1AAFq52jQKAc4HWrg7YKcrOGLuUSG97uXme1cx4xekZh
nBH5llIhj09bN48Ed53sDr2hEET4FQAk0E5L4ixeUMhYAhnNjIgj2rF1xr4bLect
eU2v3GXLSkYxwgzaIvvX9Fvrd9pJSOGEHUGjhV8hKw0lFk/jOSCvGfhh5BIoEmhc
UUWtnN9PjREDfOoce+wwENOLbG4EmXeR8/H9i16ZzOqoWDe4KRJBqNGQdhhHkC70
ahU9hrqgLespDQgPmceosN0FT5XQ67eqR/w4oC1JlyQOHYfrO5xEAQtkrGPFuytX
Kv9pVcKmVL57yj2LbBS/fn/WuZcpZbwjTDyavUrcF58NtYlWuN4s4F2EK11K8azz
zWxgwf5wDLdYSMx8OWmdDpFFMeRypPvV1MO4e9OJjDaDpcAkxCsHPZSsYZS0B7yF
5O4akHwvJW4FhH7MXOImfYE69S0bSH3pOCHALV1yEpwetQ01yEbHLYwQeshEq5Q/
0P6U/SxBhOSKJ8C2OYX+wdPOiW3//RGsUqJ9T+ldp/mav3Jb+B8kt/cos5KUeb5b
56kefZ3sIPqYAfLl/5/nHPwfRTLe5Vw7Eha+JcEWcdDCXWqMJE1qD22JGD2Oo3TP
gnCqAPXk73+IjVYUdte/Qd01zGy12PlwiEZ5HgE42BucrFgQjCruLh501hXuTyt0
8IB8Nev+l2nr7U2loFNT28vkDc/pWcEHVLptoR7alJWxB1MQo8KSNzS0oRgwMsOF
uKErMzHVq0wU60KldneyTPqWjTmtie6iA6o03w7mRf2vbO92YpBgtPVJ7cZkfW+k
KOtIRgSSbGDljtvAB7BFftKbQYD+NA6eilpL/1utwOE0/cG8Oa5Wk1FraA0o8JNS
naB14PjSssu2drGO/aSy8HZCJjrEIW9Ral4H0F8YwTPJqzSFDd+TB8J9w21XBUYi
SJu9w1h1f95yMceimMcodUrdzrySHf/tGSk2YG6uTWAFG6f6K/SPYb4P3jWNtkU9
X0EJKu3zX9XvSUDVf+NiZkPMiIQz9dKhATRfZrNl5MgYpVSgbYgxRYCJr5S9iPtn
rWoRsWMcgRzm9trtMrZpiF5TAflgLuY6x35A7SCZGKkvkO+cH5cPetETmc5zj8eT
G0Kqs/WsR5s3ESOGXmpFReoiyu06y2JeM39Q5y9zOxtsxk4T8MyX8r7LVHExODOt
G5cRLWIMlzgg8Fl28asuFcn8F9uz8p4KC3mwKV8+a12TSTcETvcJQ2yqLf5aEeqQ
28SO52FJfTaw1iCsL5UYI3YGhiOEHiYqr4VLWPwClBqoLH+nBPpFemrxMPNg7iCN
LwF401+U2lrAZSG0ttuxiAL0fjSsoBZLcZ/jiFaGGf6nd9udrFmXUsX1U5FQ4qco
sOtol1mfk9lHqehm9Y2ofmf9ToWOoGYrwGldkQEBIbN4Bngs8DtVTG+BJm/iVtNK
SykepV6XZ6PESrRnpsV6rR/dkRhdgSNL5WGVXAKdXuc7lojeoo0HnS7yQR1kqMia
RA+jUkxwTqFZRIjExo9CrI81kK5A5XgeG+Ho1AeClf1/3c3MothpjP0jxHHnNlHZ
AgF1mCwDsqJRJ+G08lS4LvOPEku83vQb7a+zWwHgi1meOcBTRNk3ifHPEUK8v8Bq
6Fk+DJ0sKdEAsL2UVm7TQoLNkGkqYOxtZkOcz1uXVpzZsYCcdzPzN5eYy1nj9ypK
l3xTr2Fk8nPMb6olUT4dyOBvJ4ylqh0mAA7ieKps/ZYQWMEWq+6LqiA8IksHjyis
nGKtJia7cl7dfZYaWl3FvtQIkCCmiXwhnCtSOANoeNuKrLRdUv9JHcgcPXPFiG9g
6PUz/UVJI5ynf4AXECO0z2kRVSy1LZH1k6AomL2GV59IrDeJqfCXadpKbGmHPAnk
V3RMayHluaMIAYWkq6Fgid/Q6pGlFyyDx/eyQjE8wNLxpippsmubnl9ZpVebBgmv
USHzgxSmQDEsbKEN2rS69RtTgiL2xzNhUjF/rYqw2uZsg7onziJfL3RfNDaBdFmP
Hrp2B9zMLp2gZJdzJVz9fa/4OHbL9s3hMJu6fLAWeongWA9GY+AQRjLJFv1PLCiK
9UojHoUf08KV2mOEfpdXV0R35rYqMfL2sjCG01nIv1IhxO1fOUyKe7o3ZcdW3URH
gVRF+XKnQIkd10BhQLCzpjM0NNW3TK8tU3qjXUe860/YFA5LNlYWPfeyjf3EViT0
jLUhuxAuKz8VnM63gTA53NOrvFL/uQMLhTqdL58jA0sCqx1DQqiF+ytAmE5Fr0zM
K/G9jB7uIIoVJc65OXGEf0E//wHWJHSbMJWMQUjTSirre/ViBpdbUCBqyJ4WXfBg
s2k+Km25H/SKMI2jZtxJ4qxuSl4/iObu7YgHEtu4uHhp4PlrLRlG8BfTr8C84W/J
skoaDfHbgHVWIYqwEIcOMq3S97rgkYyH7qah5vRSt/nEt/9CA51knJ0Q44/N4Sc5
1ttGOGoEA4y+2ikYS/BAtoi+78slERyRTGOuvDZz9l1SqfvwuxRv0YijsvI1kn03
evJ+B0TmnWnns1ttHgdfEO5BRopusILWqzDbQV+Vo2sedspoQePYt0Ktt8q+5LIz
c+Bkupj8dOtYazQCam5+653ou7W/8LaGtbZLH5TQIJ0B2aIX9X8bFN9r3Havmhz/
apEIPqXgk2AnCySmuh8lrHqKlcv4hGLhOaTL9Uw64TAhgApPGerX3qXkyLGkDw2t
BFTpQ+FY7bFUqsTAdios/Hi6+G6AAcNORdEOfyQ764DyG4vR5oGobHM/z5nIxveE
op19q03SICgFDJm/7KrkvjEgj5+t2t08akNVoC1FcMTJTVeMRFG9sXqZpCgJo/oo
Syb6Ciro1tKyixac6maVInYQOoq3GbZmXiyMF/PD7KrXSKwe8zIfvNMpg2vJOJwP
ZtX6U09iwzp4t1QlBB1AIo6r0z4CZWAIMHo/MFNIblBnJJuO+FtM8BwdwuZFYhxW
8OQpRLfnPrRXPabj76TsFYa2YedtJUMwqSx3pzqpGIAgmGj72+i9lrnLY31/O9rx
qXH1Z4f/vl3tTU4ZWG3pf9azmBhynVq/JRMnXgmCKXEpX7LjGvSJTG4oBpB4mMA+
XvBAvTp2HFz04x735I4lrnXqv8ye4qJB8/v4O64ktBq1IWodQ/PahO8PTHQbHZ5k
RlnCkIiSwy3EUol3wzr6HR61D/u6ObNw2TPpD4yLsJm73ExZzX2h+LdYxscwWu+z
ahZwm9cLBdUexNBCcKjiBIQAzqNKPSy9rP9oIqHSbR6Fm0fvmhg7Zfr5xmw2FHZT
+eVGg4S+Zt5czfWinCXVuN2dUANVmbB1hSd/oVLGng9hjB6sVbHA8asgM8+aMFFY
Lm5plxdft4gC9cC4VCnfGqAjAfMRHbQR4kdCfoNX4KcxqwdwDyStmMbq6glv5ER7
u9wSULrDyD5hdLUb8VC325l5ek/un/Om/kPkgkwcO6iruFUn0L3aHHPM5EyPzeF0
e0Zdo+TVhZEKBbv4dEu85KfRC6lr9rFi+M3QaBMOJIHPf/9n0+fMYPjy9K/ZELnD
P3r5VnGXn9WRkC2SEaWo0lZf62J8QomITkwdIDLpHH76yYtqrUNB2mUtE5IH8eWs
A7JEFtRBixSDSbTF90zUR5KJ9G/NbeQqKygZJwGjbUmepcVixz6eCL6F4Z30nc0E
ULmPO0Rp3mo4gjJobNw4Bfvi/SL+/L6CrjfyXCS5lZWznUIZDQe0KCUHckFVD1Md
GfPI8QXNfQIJSDsChUu606TkLkzDbT++lSAl0xWKhLgmOkFfRjNhBoKY4PvyRMHU
cI2xfJzVivJzSV3GW1odghHTX2PBoXJsaIMBNjx1joKaa4ztsL8mqmjmA3E3jnQx
dTg6Ri2SnQPPk6PXHGkHyvnZg4UJgYLvGrtIhBt2tnURouQm5r/12gSje8NyADNc
dFrP9sXFpQWP2r7vjGyUOGCrUPj27MPvk74GCg/uu0EOVh4cpbS2G6Rg0FTDJcRw
2cTBg8A9m8+vosN2pjomFIPsBEgngH5EWyqs9suNoNvkAlh43GZiHrBKvi4lQovT
824wGrr9OnRrVbACqclK7obDmsoqg/HeDadjRI0xxnnSOaJEWryoj/kMOLAEF6Oh
qsdmZYUEigZVTRPdv/4nooJbhnNXVN1orq6/u2UrKYVwGVT0gNiVUSHOfGLYAXUF
uOjD8+3+kD5UtBoKla45YhK59EmPX2cD2IbgI7pDym4S6WzFgRspH8KAcj6WJx35
nJ2SR4iXTEw5eWzkrOXgJQbQFIMvIYm/McBFPvhLWphhGjeLfBLQm8cugScXxyKH
bbzJjAseVqnrR2/mrIaQBGrbPrP3NO6nJ/L7d9Gn0KPLRLaexAnkHTqT/qVzA2E2
69G+S1Zdo07c3YVt32bX6LcGsRd3oTKx7b/3ee+valZdfuAgeUZgnkzbmbF5CsXv
omVhPPsdVbDZrBlugIJUSKEodVMPp3BEuyo/OHXPIj+48eVv5UcYdC2Uwceonsr4
DiRFOLzVfYI2/lcPLT3T2Uy7pr/n4AU6dfIDaRRf90LbGpnrKWyu9KGlI+NPfkLR
DMV6HycK4PfFS6SkKMQ+0B6+QV4mjRmtKSP6aPqilsr8oDDS8RhNmGK40drknf1u
5drytG0FxiuyHvdXeNJif+q3rU3wTNQxkL/NEXS3XIInWAlrp0hja0QibEw3T3kP
el52WFswhfGa3RkmALM6IIH3Uh8kCOfVJXop0jkFViGk+62VXZqH7iqZs9YmuyG8
GNFlXHiVUMXQVpiAZn4iUaUKdmVRujUtUdArQmptGXhAfv/rsSi+6xw1YiGMPQC6
BkblwafF1WYtsGO5Y1yCu/6CRuDZooq7UgWRicJCJdacTgZqKWV2Xh7LlmlrIYSo
eWFUMQjzEVVOjc6HZGhYcivGWZRGu5LS2VCHZH+k14EZ63VWleECNWOTG8GlpN/N
JMckNJRTw4VuMfxDqzQa8m3AxwX+Oay8u9B7gsk927RKI0Qnnhp20UT+ZZDgvedx
Pf4tjKkO2ojiZ0cGEBgddGv9fjMwzaxSRyKbd6hNVevKA1W1t7UxIqsx4nyu2I89
mbRd7JE2pLXue5XRag7ue2uUqWnURTcvIkaTaKfWCqaQZTUxqcAiJR+FBQ+l4jQb
nh/pz6mTGRdexoO4DhGA+GZqhMZlQGCHV+uemPPJo8dq/yOs6XVe6ende4P4CTR4
5j1E2IfZA0GcWloTlT3amlS+FN3s+v9AXuPJw0HKFf8NT46dO0M+YJ9RqfMSSHFE
ZBKR1+JiKq5StoKkLsJvRstHPPGFtezOa9/dtJU3vM9Pb100/YGFrmAqil72ecoG
jfmGCS4Gsp0HEKj6hZc+14IL+EUJD0/D7qVTZupu6v45IOgOSHl9ztkoxVZyL9YY
fCSb3Vsvmep/XwPZ+34oK3dc2JdGlz/LbaLGH2TRrgDiJDMausP6owkpRUZeRbnj
ToBNcmoTnTxrrggD2BpwuqEnn6gFPy7IItvdlFXH2N6S7sNo1IiloTT5QN4zLdIx
qAsnroVc+0XFF6+l0t7oXYqz01Iii1eguxzDQjq6FqEwJIZRkDlmK/v0uIIMRjh0
v1EzW0OupzAs+sVQXITOUni/libclNUpT5nJXRmuzDZP20loROSJM3PyGuKs3fyY
k6h4mxthURHmCyuLUQp1hpashJJ4ricSSyrZHXmA+pWIYZlCfSziKAlGsPh6sCj1
5LUR62W6FnWf65oSQ900z7q4SvhBmORQdAqD339Aq3h2WYB0QIDe8GlFffEoKGPu
JEwB0swNaw5RlGpTLG1HFwQqVI21oBu2vpfDbj/X+iNWzvjBPvFVDIqNqvZ0P6LY
N9nTN34zvDl8F0ue19vUnFY4ZoXRLcbZfHnXW5sx9MgSyqyuvZVWkl4qcFkP8LJl
zYBwDvSN3KbBn04eFfks5vg5MT6FUhuKHFVjz0hBxeZHw01z5ac9BG+xp2Zn+ENL
UR4OnwQuDU0Zoo+Hh+NR1EHwBKNX803VDNaBV6RxeKxu1fuJUzyz4gmoMx6gzskH
h4PV1sMjnRaDQxCOfyY7z9p+70192/Fw7yjFNa9EO3FEp8tyzZfIF77CvO+ehQgA
99/N1QV2wjBnIE8nY5mdmUkoUZkaAtUKqcIWERNW8Vc7p1hp0buNXIWeto30ORL/
VXXIHqmvicqSsQHnmL9a6pVfmsMt1W/7bJ25oLl4g4lDOnKe/jhbo67TnbqmKUoT
YOhBLRSN3P0PbDrdUhg/uzmxCfI9hVvIDAJp3sJkGm3+y2l7tkwSFDid2YpKCkMU
gB0ymlT2nQl0g0jvG6pGu1bVLkgO6WEPxk8PyUmp4RUtAvGnMPSv/IpWuiaTuVQ+
4mRHBS99BFpo33A8hBMS+2VmzOi74BCzEHPfiMXzD5Thjju0Rb0yTxOP/QXRVTrn
oGzTT3d2JS1LbELJIRkF8WX7cb19xvNglQJ0G28ns9lIRqVJYlHgeS3EX9sdOuNm
ih+A1Wp3ZGZwhkPI3H59hmKlFmxZGwKtOhFKLGNw9Ndqa4OoRBEJzKVTRPGspv2o
X4En8XXNU3sthCEvwyEwj7/C3liYglLxuWdku1SNIFpSQNJite+QVkLgdqaTmaYN
7GdXO7NzJfpIFUWT31feNeB42j42Ac5/yPrubwVAmn/7cR/56sgi4vaO3A8mmgKY
QGpBGn1jFZG8IL2ykU+5HFSOHSIRz0/RS0QDwbUaiNY42JNH04qPXA3aidjrXS96
yJISnCpuEbrmU7GZtGSYtj2FCKvCRBw+y2JwYK2KkffEECFqX8IJ+ZlspY16Q48d
nuB8aKcHj/UXulPQO0VmK0PLsW5GR/juqyIwSJEi3DjXEi69bdhTfIxvbymCZuCm
sMSI4ybxA4AygXH4bcKEHCeQCt22SY2CJY99onVnaqoVhLlC1vLRbI7nKr+JwdBv
Wz2Ss3LAmpheai4Fw7KgM6sGyJ6kC5WsB7WKEqkq8fmpHaqPjwwD7oM7SCjQcG16
MsaHe1r7KDjhyXjucWIKeNBN3VXveVUdVuby5YTjMyGeR3t6cSnfChQMj2ijSrpV
b6mIUEf+EzWPWFuObSjC0JN6feXeUcvzgsYxbBRkEGtA/j6VssMUelScahiaA181
7uYNT51mIgCvmUgw4ocvbUJVbBy5qeURVS+t1Wcg5hRPZ5JSEUeGbEtc7GZhnFxo
TZXl+s9nSFtFw+A2aVa9F2RpTx/ZKpitIHOZa1Us/l4d9x6iSUZm7SESNUoCFW2i
ymI204vCWKmu4pl2Tk+SBRcf3rWqcbo70oQ5ETmULrGvzpyiw2KWvYWtPNUCPSCu
fynQjMUtQTG3sCnszjHwnXouCPCYygdj6I+KYQotOUDWO8pE2FnlrsBEO0aXKC0c
ICoDu1JJDdE6tUN9aVFtqszmFBz1e4OBcNDQyXQX9UEMKG35gNJZDA6sqtxdygBh
NqiEEBwpRi9yp/55iM9QyganszBXUK6lcgRkZtyBNqrZzqAzosi+JEiS9Wd80ZqX
zgAElo8wEsK8Y7tSUAhHBKjgBuakfu2o58U8NGUbqP8qU/YzomXFAEUMPsUHQlvN
pxgqUq+GN5GrGnB/3tSLbJx8YJhvv/2bpHD7gP+kHCDnth6W91XXtKT0CzB3OP1K
m9QFc5xsKTy6ys5pUGD2DdAyUP1M8GD9TlGWFt0CWNx6M6BzbSHVW6CDHjUpo+88
3G0QwrJz6GGLV6Mgq5juGM+C39Pbpm2jUJRt8RpR+kaY3vLekXmIbQt2++LBKLXA
ac9FBppeeb/REnKpoZcOZ2nHIvacxddPnw1n0AMtUeUoaZEJaycQgJhO84HOeKz/
lTod6BfkZTmU//RKlVS7LXsaoaTdkXU0FWksbNMkTMnI78J48pPla67gVeCwadoH
H+dnqJsOk5kcubH79valFvFLKfMdQE+83YISEmsxAg6m/3ep3V9gQH/JRsB5Z7jl
DhIc5KZr0e/I8ountlwkRAKj0p0YeJnXpfHsKlX5ereaJT0cu8UWmbqA+22BbQ5Z
HGWhCRWHobsG0CBrJRmX9B0KRS7OZ8KvSwykqzHHGMzPrn/kZq+F+KtAkcr8Jufh
S870LDSE7bqRV0SihQAB7Og8lMiduKSzwDVsff86r6AHn12r5RDkDSEukEkaVcWG
F5h1y8d8MX4KwZ9iTb0u344+98eXkoNOOHAV80xxYjTJ2J7F+TPjdmiqBRvMoBtn
W3FfKRUKtAeWGwRMYxQsKMRf6SmjEpr5TSFZ71nzkyQbFTRb1twNjl2eVR0rIyHA
Cv9bjJbJKTsMDNsmQDjS+lgVDAOePhaoHPv05qn+nYpt0GO76R/NNQMX6nnMy2WH
qucBPUY1560WW3q/NXUyvgRNeKKwouwMPzxGy0RjnnzqY4UCnwnRZPmIqnx+I1Uh
wo2nPSjV4n/EKL6XgX1TVXcHmiXQT69tmFLTzsRGaY5gOQm0xmjyUyOhpOBCpP2S
6PDuxLQbqnt1DwW7aq5+duvuAoyUd9vySkxo9WUPp/V5jie/EobKlF2RyCMYGrt0
8A7r78Vycg/nKW3mfPTVhkYDDh/fyBSxgmUXxN+8hZJsV7QZkbYcYfpuITW4U1Tr
Pi/1/53GGzj5346jIy/cmcjL0fWqwV20bNzaaz65tCM5umKEh8jvwmUBl5gZdAZW
hyiuSRjTq6JzJWnsemkRZFo6/bpl11Zfai4ItcohvY2bMAuoB7rXi0621KBLUeZH
fFczc6F6VJH1b5WYe9RST7CBs+eDg73dEUwuVs5jhdWgrrU0Ez0ijNSXUaqn7WRx
hjacZHLYC6dUgU+OJ95RI4aexrcbGi+1o/hBCEWqdVcNZmiQewAIwzz8Qcv7O+UO
RZWlKngew1HgCGWPbXJgvRwk70mnoOunySAjxybbTnYoW5SThxqlJvQCUan0Nzlw
ojBM7sbp7itFwQ49c9wFDlqBIAz2DwPOA5JAkPeUYVnK+a+vn2qLplm4aQGmicwF
AlmXsDat80vxOtPJT1kPyo7gmFQ7FBplzXCgB9xCq+rU8I+TXCct9EcslcjblsTw
etDfGswpX2X224jTlWSpuzZVBg+68zI56i9jFImTqKeer+ODnDBom7P7m2W/Tx8k
01sRDCGaBnjPGz4ammVBkxIXNOmzfW/QNhcphnEBkwXp2RpUYJAEd/amyuVs2QBd
EYMbY8sioamNBhmSxY/3OR+ip+5l5xn7ttDCSTidPO+aOjwPGY9I7zGLyaHBPbsZ
U0n1NN9U+rjU3RvZvd1h+qYm2r+rqGbZRAzY33D+Pexd2Tey+sWxS1qQr0qSZejU
d49hRPIsy8P51GN1XOf/aBHIuwPt0XQiofgC2T4sqr4RCNEVdAwMEjKlPERrwx62
+zW1P8X9Jg8/p8M1U+XH0n1EStdRG7aWmICEoZ8gruZJz67um3p1V9tXCZ2qYQoR
NchrKHs0NCZVXz7evtuk3bcTd4cN7b2GRsKkwGZUjdy6PkwjtcEZZthtQmt8mJ4F
wiRLcHKrpM6fcxX1dZwnLSombtq96VeJfX2kVUMs5ZBrI55O91orH6TXPAJoJ5pX
t3NMscWou5iTqJD4VeiBvcOwRk0jG8Oz6lJ7M3VvpTkngkLdmZe0jkFdw956c+o5
Z/iv40R4iJscHk0aaDA25KqH3g60CxiQ99JZG//TLMSOiedtGrTIXlNfeegGHM/J
4nRQK6ni+/rJpq8zErUwpCSeU64ugt9AGqRicYYLx0MJblFGC9l/SGqSwFonDx3M
Mg0E+n4kme/ZbZ1t+P/2caNaP3Odl8qpBXOUdceSOIH7SG8VZQV11XzTr6LsBsgz
HueEXKITFsJ6snBjgq60zwpv8AGgGf9Hnft+/ucwu3+yJSx9Wd5+D3cZ/Q7tnaT7
lITTbztvsrndXVZOxAbEHeUcaKUVp5kYKFvAJt3CpHpa5+YlZBu1da9qQGQI75JI
21QsAq4b8c3P1VoODLjduxdTyi61m2jSNhakTYIEX0nKm7kx9ukafVHOjyAe2EZw
6qJScK34h+bUD6C8ZDVza5rsjlMNjThT99NqE7a0HzjoLtEuF3nMnmBBlLbGeFfg
jO25HHwgRqUKsmpjjLlSo9fsP6oy9uYztqCqQTUASLpQvPsRgdmsBlxTq5C2+x2Q
SDYrtP1jiWXH+eSPeVGZgddAQtpJ2lnxlAhJqbAUqpI/9GK8BvWRUYr53BjSDgfD
6ztzBWRMVOT1xAlsdXO98byVKbsAjysPbD5B12R3IHwyrpbkXWv8IZlACUzQDaFy
SsPvbbWuk4RRpGPUTmmDAHO/AGmL/7KlpPquBXmjGFTjbKKf6wDBdtUWo70pvLye
Bh+g2gKfnUnWFODPZ2f0JOtfeuAWdVEC3yOPIVu2sRPCq7wh1RC/n+vxO1Mb3R95
BQQJpaakPsLHKXPwQUUqvXWR3voIXF5X54tjZX+dW0mZogC2Ff6gpq8HW+xTvyBS
Y9oLBCVJ8XGN2JIcEoyS4py/BNZL8rYHm0FqW8Suh97T1o6SWHZiedFsoTCZUkeA
OCPnkVWgMVIogQf6h1rN9XDO277fy8v3fgyA7tGB6GaHKi1UrOrJlr4Oqb9S/zfV
6B32kLe54ycYvRoLk1GvgNFdzNr7UvGA1CCwDpE2FPJ6/24X8P2i32qU2bq8OESe
liAwAABu2ZKcm5PhKCmLbLC7DScGcv3iuADx+EXwBn9GG0l/0KcD0BFNbHN0SGfo
8WsRAz6KwNLHUXq3yAsEJNYfSXh+lxFebIjghrmYVPJS7ZmHsmU+VowHRnBrJ0uY
UyOdPT+W8WvAAFlEE4ksjklHRPsSLKynAwxwHxxDv6d1WZzXuRIqSk3UkiJx+pP1
M5reMWSp8ojaGjqGrzQb/Rw7Py4NGltfTD7YxTpg2AnTF+MyU78APdYG7iHuwLjM
/8bB3N7gHb4YUX5FBtn51QA4rWPS3mRyLG+wOABonRgvlj4HW7nOThWuy53hS88a
uDUJAzgErK69zJ91fa4eFTWVv4XF2K2uH5I3uQaX6TGYu+mJwrsz4EMkjrf/gTJB
TA7nEFKz6W81uuWjeqfDTLdExw4F9iIghDlsQdvrRPFszsQnBtp1HAjqBd89N7sA
LX1wIw444e2RwX9KF1Gb++qTlIdQZREm63lSRB8rpQRuDAmpkshTfFMBRcj7EsV4
14MQsYn1xBQa2Yyv2A8GDmlwmm252dHA9kFPfxl68cvPhadDxGhrRpzIU6t4H70e
pLYawl1T/gye7pNsXEK4j1CCRTWzNi6dNNGUDlB2tbEsPrkgYcnSYLtHPou5TlnW
4aVyHQiKPePaIAncbt4hJmXzLtFv47tuWIcsR5n7Vkast+cTYIHA4mg8ARLwegbR
Ag+fhs+TXlEwt8OgJ1+kY9PGTrz69j496se2DRjt0RzmGzFS7hWpD8v1AHGpIViS
o1Wmrz1suomqVVjUkQOMXcZ40IGRtrOAWIrdjVmRUxR3fGvXd8qh3QwCbn3zGssM
ToorCYAomKuj7C1j95RRAXpJprkQkj0BBJP6dDOCE2kDC7Ubqf9CnF0G29wtxChw
+rAMGSXzmvHo8MCh5AQJ9QW6Xxw0rlHgjB5eYqwpZD0pojzflLYhE6ImW68OrDH7
M9RueYWOCugPyp3kV+P7cuIbGgXAlBVtEiuKq2gCdn35GGxRL6N+b6B/936Mk7GQ
uRg+WfVIgcEgBNUCwDp7Fus956xOSBR5eBb0REweaD3mSUmTfMoIffb37i3J0NbI
iUGbww7zaKUdjXA8P7Sgdhi4jDkrN7nF00MAOxRlzeShgRV3s0ycGEkg/oMq5q3b
COs2pVGsU8b8xrWRBDLAd0rF4tzcknSy/0nuxyO2Vr/KK+qw+pi1SJW55v8isH1u
qKGOFfoZNifcvZyYFVQSYrSMYWQFs1DFtvB1RmtD3eBtQ+i90DU9qJ8zzzoUSKyq
8A6s8+R69L5rEa9IqkZFxhfpuM4qGAePZkZt7CGoofmLCC33IrRGhAcOqlnKH7Ys
IHGBHRWn/zC3lmcRxbYeO/G6ZUlhQzFUWDrnU1ehk2OLGLkZRcmmyS62YiecPGu8
Lt65KzL4a417QAVtOQ1XGr9ZsU4sGj4QvXfXBmlhcGGn1DsqPI/Pd9bbqNg3u6tm
NxDhkRHqMQqlNSU8G0MP1dIr6WQE3EJUhU4tBoHRhvUkuBSfHwvyrL/C1qg6/pm+
4CcceXm020rt+bXKXdtYSfmDutqlf8hrYJ51+PnjkA6IyOlHrdx/fKSv+JKrwq3t
6AWCFCd19fqu+/QLLPkzj2Ag1jkKvZYrwDUhdEsJHBxJeHdsboObS5TEZmIkzMQt
UqFTN/T3n7vhFhJ6Ry20T2Y0W4OVwNRNETfDYpbYKeZc687jZ7LuxXhHntCEfNTQ
itBXj3WyV8fJvVl8SP47EMLUCP/86TfIq+CUcySfnZY0FzSnPc7htw6F4yq+Ytyy
EJdWlyY8wjcPrJheGQ4Qf61sHtxNm2giUBaf0v/FM+jB8BRSy9EltGw0QXi6HpE+
imEmxRJZVEFcoh2cKY1aFaRpgdLwVX7RtmS2Wx+qmw3wJviQV0s/asEuERlT2fF4
Dej3rrPuwyLgM2OnlCTco7ZcMIXdISZY7m08om9orIBm7UN/OaqkdFol1yS+dKxU
Omqt/TKW/D1/kxg/t57833dR9sjq8ak3fBcZKsTZ4/GLGCQfp3ku0rjZR+v6X5S8
oSnu4nba+ZOIv7BRab4rmzd8Jm16ZBuVhXy5u0/MIq0zQ69a64xdF9o8roICSPse
R/DUZ9XmUpPdWoHP7NvfaoABAQPShxPReDsQeqCWYVUzE2wPTiBh/lTH1XsfhTIs
Cd+zWxfsK44QaHZ5Cz1S/3/OCGZx+PubzsoMZ1O51gMR9XCTfl5jz+TTB3AP2T2Z
n1Z4bbwJdRrIsIZTIP8A2dIxYcDnN+FgG/Sug08AnNnXxYP9nRJOJm/ZyXNq0lMX
jEr+1f0cB9/2B6htunIVh2rHvrEPI9bVbQd3TQltjQllCvFPJ9xL0GiOuNtz6bpm
GGKs73Mdh88SxUKFEdA3DRxBh2h2iuB2Q5jBCUdpmXw08rSOlTFE9poe61UwyiDo
J4n3AgH38OISoo3esx2am8zV6gFYgoHv6l8RiDc+8ASoJuBM8L4jU4McH3PRpC+I
t5WUhGEVnWwA7HtQEBi6FdH4+HO6EswSqMhRhzyrCqrMOmO4QjPvFGWSMQBi1e89
0s/2P/+iYc366q+qwpy84eta5uTv62NdW+Qma72F3XQqMamkcnlPYoOCZQwkPb5U
JEIA+6+OKfwxiUBFRocp3zgQcSO8z3i4tkuBM7gonH4CJLmZZHSIlcxoDYOJICFy
AhNqt5+f4ITwtCA0X1/PDSkP9PhFabZwQQk5WA+il3IRyFNJmEeXdNlBbN9Qb7ev
PQPHC09jVIBhdJokpO7tlFCnC7auvFRsWILrK8F/ZtHIHV+D+y2Md/4qjGnq4I5C
Bk3lobEpj/AWVYuiKl3w++vu7lxQ6EtkYJPY/eBDlxIMY28eYJsUlTuU0EaWT4s4
XLrVOlgyhOEPsnPDTBTmzRmzOaRpzIyk6rDCwibkRorMlCYtktKW9cZktFvJe8CJ
TsteCw+0hycZpefMJ90zQptgTT46o1gG9uOJGVivqgYttSwE6pvIa4EKVvIHx1xr
ThFhZ2t+LhEG2RIMlj7A1+LkuvLCexl5wDs1jndyWU7OnLPemLXMBUIH8YEtwshW
gCGc648qiej6mQX5zu3JerG+8afsuOTGmcmPv+FatirrMYieT00PvmgE4gcuGPAx
SVzkS0UD0BWGkbT2j9K6ybUrAqxO7qDA6U0JiMNZHWiwD33Iq+ZHNvX2mz/5zwE0
6cyCfh0A671E71qKy5R1gNzbPEUykaYNheCrWxBXIizKs0nhOKQw0hZCjl2c25Ki
fBu173YnHeysdOu3/DsQ0U2pWNriCxFDwQBOQ1rxKLFGwap/RexmXXdPPxbYFpYQ
iac/r/imERBeIuNmdSLpb2gArNYJZn37zbLy38LPoynBb+o570VksWgfiXGD+i0r
QR9X6sPO0poO96Ix5nTbVao0MSpi2FWF6OkPKE5OpW883tgDcOqRTHa2WdllUKnx
ifRiwM0wPFLuIv3COGgsSh47qUn131ia0gviEbWmZpsd28LWONY2QsoxPOz4OAwv
AZLZsaJreztuDK5naNNy7rLFk9YjMYO4BBilV6czXNGSAZuFC5ZXqkzRdkzL2NFI
Q0Covvsysvjxjj9Gd/zsygx5rcpFFcCxBR2mBWo6tJdgMUyuMAE+M1AVwlmeukYl
u2jcYAYBSMvoT7/+kns9zZPcbQJpFzoDNEw2PzRHWVGEg7R1z/OhjyT55YXewLmq
yhv3vMkrMM4QwIyeiENsWYB2VfcU8MmhpsOhDs6hYqqAhNlSfxy7L3MsaZe+Yq81
HGqr4mZiEeeOmD3+bC8DsLipCa26aMAQMKijrjgrp5LOppGKuMFV8/KRGTstKtQt
OmXUVkIwYi7dLjQzL9/2HjEq9i8S/VD7Zp4BpaC2eHkobZp01GPM2NEqji9uxwFu
SruCCJT7tLTUWyN+0kwE4klFcE/LXsztQbUM3PGhLWY9dmuJ/2VvncArBBkwLFLB
WCV1Duvf0lmmQm8sghskuAZnQ/1eb+x+C/tmmPWEoTHv85oCCcWGAIFq7eHTsSY6
IzxJWGlEJF0L1yo4w2+qinw/uH4IxT1ErWlpzOYTwnG3wBpRYNj6sMh61UPsNv73
2ouLaKPOIpT5IUuJL4HOKQXcnf4EJDKqAmzJK+BoRthZHdKrMn6g3FCRfBQd33pH
jQbkVTVjpTfXGpc4utbXJI6RyS8RBWPT7G4Hq0sIvOH9sRph6jAx25Eqr+wFd0o9
fF/U0CvGLgJwKUURuxPL1BbXsMDAat+hKRVhWauJOyxZI7lNOecuI7nKEZvZad5v
lClpw9aZgQv2Xn0PkdXgzRzBwurTlUJu/ZxqiHYAEbKPE2Te8Q8z33fBkpFeM16/
BlPUll3KrNOBdzBr0FdT4/eXTEu5I56KvClc3yC6eD9pyxkqroZqj5Ft1ua+Qvuh
7/7zY9w3nYZfEni3jHAn3UitDpWYtmz8XTIt7KSqFkPh2jv/GBw4GSfjAc2AwNiT
FgQySbCP9q3lzXVTW6h4+MzPCL0yGtm8w+ta9rZjvOsd6EDRYgmeWtDKGhuA1Jcn
eGcIa6Z6bOqkqw38+MlW5VLace7YSfNFfx0HDWqzT46GObAu2XnzLZJiCgwUE0gB
Xh1FGK14A+jbqLOttG2KKOnNxk64biulP9Vl05tFfyYgAP+7lHrHIwsTpZmw+Aik
w6CGXA3V2LFnxqW6gKP4rvFsL6UNdOG7gHf3BcDHboJ9phGxQErJKFAOO+P2mIfA
+LhLkg4G8Q2ST9zzfxqviR6Zhi97krps4xFH+RDmnrq5q71XX8xb770qtB34PZ0Z
Ko1olIWdKOBy/1W4jXsryFOpONEpvtLxjHnYmYYS6bCutpBQbpYAvAddnW+h6Mxp
EDtJ1MtsIVTUwb3cZyaTKhAu3I4PFjlh87UO8lxEACDGr0nsfBEKXR5ZI+06K8vK
Q9GbBCqHKrnmtbwCQAuQLLDMh30LcwxFoO+cHxSiyh/BjIIv77t2LMHovHPSlS/N
4KeqraE+CdFPDH11edz6OmFpS2jkTv+1+gyY/rKUhWswW2ouaoYRliwNau3Msb+f
tHXDacJpp53YcnE4kw0I/ss8mn0zZCQVoudMX4+KUtDR4frRp+5H4XkMfRagl5VS
88lwonfcKLISr86HjmZGY2hMvJx3aKT3KEqHzxlQPkxVFVqW3wxjoJmdZEVgiOhO
60I+y5yPYspV6nL0SPKPY5tHCvw1aQVnZN6MfoxmZCDCU/eYTRb838Ng7dAeLc+P
cDKouq/TnI+sgTrjTa1ZQYqVA1VwocciHrNS7UgqEh+HQOQoQV5DwYoIZcUhK0Ui
xIF2QGjcnv4RrnbmWtT5ULvK3Rc5Ud7rEhgocsgcuIvA5HUaOQp8KowE0+tXoUcg
gyT3zzmqGL78IxIw+jGlAzMJylm5APzTSolvXDHHtLn+2lwbtiKgw/PPe9h9BMcK
jFOZcQtzApOaJ9ljH5hjdfO+VuV0sraDlfl8k88Neu5tO587EmHnsbYfq29pFx+r
0FgKLL2D6LKJ5LknEnhOdNVvMPamQ5jUGS4dWHPmd31+R/79RnhgViSXgrIdjaa1
2I5Gg6QS2MZPhwKDW8Z34xHjMS/KkGIqUdZHcudSkmyFi77UKIT7N6C2KdIS4NzU
5o+Vt0f35wHw3+e+FYMQMsLigK7R9hWVx0ShqKqABGeCNpCrF5MpLSen0E0xNOyK
lnFXKlBDIN/BT/Q8tVZtWIM98YoqEYt78Hycd6KzHFAyX4PpygvfvqMOIcukqlaa
9g6IrQZTZk6i9q30qZ/MiEEigVbobexP8Q45Q0MR2fxG/5ZOEZOkVli4aPqCAglz
MgFJeqkwrVN6XxAk/HxSeGY3PGFdanMR+NjrmAEn69O7O+e+8RIboXOHseZ7lrWi
KR44DMPkBaOikQl/yn3x/wvNdj5Oylgx7Pz4sbLitM2/A69jEJjt7Qk/hrTtWvxR
KiukkxyUBQUdDJ6dv02MLXGW3ervs2oORBmQrWk5+NhAabIbMY2N9VSQqXFztCO3
BCkVrVW8gU1S8YzRq0UDlWIajF4QBW26nX0yjLTwaCg7OvQegEYKy99PZMj/pEP0
FlmagyBDtGh1cJvpRpI43KL24AXmZz2i+BAX+JMJnYFxVivf+r9jGkVeh39aZrRC
fneNumpIZHd8Kfk8H8n8EklR8poc6eKVbECj2M7F5pT7WQNc2Q5Qrvj2NBRH3MVj
byPi9XZ16JGd8EwiEDfELqwhnujrp6hnoMOg+lfrVp8wgM1tyKhMKau9uxT7LgmW
UBtwzXxCDgWSGvlb2iPmMCkALt7XVeINNY2artgXN1Fd05P51ou/zayYxo7aPjif
wjukkbc64kYgc28sGN29lGNyNW7CYhM6sYJIAirP+LRQ2wPBGK1xhOXE52s+khyK
cspnz69PFzCEm4cJ1l6swPjSCub2P9UVIr7ycq8j0wDUEVoHv5G+Fk0YoP+3yeKz
YUqA9a8QK3KYbSby9Q64PlkYkrXvvVfx6mC3t4Hn+rH0lsSfkNlYkMDDFU2I9gGU
Cg+sghjmjGwlvpJBXVwkRVye38oKxyzy+SkwrZfQzkBC4ZKbTZp/kPI5T80oqYPD
D3DCtlvsyPIi+1l8jixX5Olc6GUUxSnykEBlAlS6fB/V+OcJGagNEACI0NVDVujr
4aWTESRUIQ6468dY5opVqccwf8EiR9MLwNwBXWQyk5owAbXLGaWP5UvIZoYdAYmb
/uxunAUixvs4iYFKSR/trFzymOmSRbEwOxTJGyAl524EmJx46wxOn+bGQmT+yonN
2roYgkpcfWXOM/bQRGAerHVu0k7yUAE3M/CrwvGRTpffzFss6rg5DUbGx471xoyW
TfPw8Ktn18I3IpeVAERwSV6Z/b2139Rw1i1LuEzUCb31/Z0J4A0blG8Ak07bG1Y8
SDA+Cu0bnYZO2VO3RIyIm/F5ZG/RimEetT9BY3ydb0T6lbnkqEsNEp6s7HP6Z4e0
30TEInkjrOpNYwjPui0U1d/JNw6lNKe91FUR1a9lb4Y3Ff1wbY021mknyan0/GpC
XapNGgYxJizgfbTo9eTZjZbxBFOQG/P5kwIZmTKJoIvHYjdDE6xekxx4M2uX4Kgp
F+Pj16CPmeeGJ4xChbtjYrsE2LBcNpbPNVZ7CAvFSyze3s1kf3W5OGMa3VNUadJv
UPIRS2jSbTEo0DiF+ICuwk0/dSmxVGVbI3TYlkwAPRBcQSVeTDPmpZuaNdF+T7c3
UVq81Ku9eNw4FiGjAPVv21UnLrtGok0lpdMZPhSdb/V/iNXRyXS5InVv9AhjiA+z
WTgDxcJXtLZIk5I2DGCyM73MpPeTdZET4GAQVLgOHwpar9e25/Dsv+zgBy85pK/L
0W/CGalyKCG0SVIIu9A8hGbz99D4O3cuBptG+KLXPl6fVO02ZgiIdLf5lcz+7ala
wEfV0NPNpJeiqaVmGdnYY/ZKp61XdzvJ7klUStPjygB9G7KRKNbdmwHuNtFcFeDI
uZAqJj62FxI8VILhUxPMF2N2uo8D3IBJTgPfxwFU38rZPcHGKz1664CdSUliopKk
eeSLtYasdY22AI0FbLPX//3jzzeXHajIx3A0fmJRjarq9BGJksQrZFO5TKldyOzi
fvg85fcuHUkKMzIFnfzVV+oM8lV7XQmJxNZWgfdvoo5s6z6TRrec1mK4i+sInOo4
HBpDsMGRTqFf+qD1STJcJFWrUu6o+upxi9vu/qkygAtpIzBow9PP1crlzVnSrg/U
P/ImkLSiJxzXPZcksDXxYoddNoGMoiWMLeKjntCr5nQxmCcykNQzi5tDMTC3gXeK
AJkoWoW/TobdmZjW8LXcNfKJFX5+cAgKjUlXjIDtX4CCduP3cFjiHyE+DPHYpLec
p4wkYdkCLJ2Svhcw1GfHD9q6qUtdZ22FlGk0OSEj0L008g8ASzyfL54fc2dqv449
mczAaV4VKntJRIxg7NOi7CPG4ej+VcgL/POuSk5WsLGtx2Y0NDdTrcL3WeLbizq0
rgrtDgt5Fp3W6wS3rQhisKFk4ucbyX3jlzCh8BFFbuv0iLfxqehm71GPQl+fZDFp
TcBXCfJHXECYM8WpSQNVmd5Gt51k8WbGBczWcsvKS1Xhd5eUtBCnm7s7IrggsktR
0QkaDfjeuKKix+zvP//scLBwKugeL5pbbVY+GWaWsLNmTSmsBj78cyzh91nwkB1X
P3FOlpWTNKFmmKU0+Yo7Qyo5e/f7wqm74DJqfd6UlMHj9iAsOKPITqD5kRqXPc8W
zt2OE5v0UI7+Yk7Coe1iydcj79bVGFGw6BKGcqr8hOkS0RyGyCRzdxBITsNm3yV4
ljCqgRSJXalKwKU+cBkGMNW4qxPb1jIreFjZ1nHlQ4/+suvqhLDXbqBPGGkRT4vt
9JEKHWjr4YJ9s6ACjit9LjEY609Y6sb+JXM3d5cY/IYGeqczYq+Ox9QTyk9c0s1/
vLkcv3ae03VKaxYrxkoHaJjlOcHnbNO3IPGaZs2YN2/9M5WE5Z3MdluT3EgmLK3X
Y/FHDGnEIp0j/Q//+tIuLB5e40dMCOG8L7oWBQc2q040GKbFUu4lv8L37zf1ptRG
I880ti2DzqW+tKezHb4xWpWa7sXYIFZt5zXFLtB3SFwDnjRtU9M8Vp4TeJimOehT
QSU4652jBGrPSGApbT228SbF8syp+wX0Vwes3p97/f4YLT11BsB5XQrb/jk0EjwK
L0Lj4zw7zGRUIBtvjBG0HrXwLis7IHonlmDocdz/3oGeLJ4FGE+4nrVdpBTyGN6b
3AOg90GKV1cvots+VCvgqCXm2svGW+TzRmXiVpX9FuQzSgkT1Uo4qeaBT8CEP/x6
o7I7nZaT4ySEmaIJkoFBXGGVD0yEopVeiLNV+Y1hDA3yyy614TGq2//TLUhY0fwk
X8uQKrQp9x8y78fFjWaUjxYqZjSLwrML0UzKiM1TlXXuqiRVvHNPC4VhgC6alw0X
gi/UnF9FmPYxXqOmGtghYfog0jesFQiMOsuENr7BrTz0xUjcZKqifadM+hBYx4ie
9ZBJ2/wmeYAN1/ReHBKNKZPFX7C8wGMHrJyVcDtgRXp/HXrewDoHOBzfMQChr2QK
7f563ipsQPhe5aBf/lWvRKn/anur3p1aAWogGmr61HWYTMSR/I2OGDAO8VmMmF5t
LBwcK0JbrMJX8MCBoWF/kp6SBv2k227ywmfeDnzIWGf7kp5KfObV781MKTnqIifG
NC7GOlyqqQAtYzZINnb3vPRo95h1JUYS0gBiXmlkDIhD6NuVzRWL6oBktwC8OVP0
4tpxq+hjtCKEBgPZnJUWd6aGKZBOnyaXlK9vRgZ9aoI5e6M3IVtuscVSidFeK+FP
pmg9i8kYJPhVbXXjyqwdr0Vs89CChgPYSmAFO9Rk+fnioqTK/7ItvAuL9BEw1GGq
FnNISqgXpPj/YIs9exPbGDksmX5PeBQsGdlOAtEE6WJ8PxWkkv8YCXDcO1kd0QSg
YubLuBJWG9vy/Qx/LPyzFmUOYNWmqh8RXWaznZnrVArUM8XGp9jPuJJs/a7lx5iY
jhN9O++75bS1z4R0MBjl/nEeprvNDxDt+y+PNYHIM/ZKlUFBiB75uY7yE2FIMig1
neKibEHUyMhA8TTRirdPRf8uUTbbMPj467IpMoMEjp+98ITU/OGVltsAda6Vkc6u
3Ku91fQpA+G3vlQzm28eKyU7efRaPbsvK0zKqqlk7vx0AGoMYlamYpAe3powJVKt
5XR6cE1kFtQxaejp9OWj4yVd+YIcJkYtshQmI56VrrleKl1+iPJOTGwAoxq31pvQ
I431q1llbX40XSRIFU76G6oUY7UQhYUtAMEd6Wzo0lrXwJZhEuRmH7Kg0rErHeLU
yuq26xQ5xSRIjsKJU8Ttv3ktveHrQiS7ntTyVevj9eoJs6eV6yX/ITLtho1tCFsL
UuID5c989EbsSTyjsohEk3VKE0H4b2fyjDitGBOioQZ3cjG6zUAuQIpdQjd+eCtV
6S6+anXNVZwm/eX7F0fwGBVBRoXlEEaBnnTXMY3IguBERIlnH1L0zLttroeS5Vyz
UqwswjFLMeiGFm00gpN7RpiZtBZFmRQ4y7qCthzr+5XJ2Wbi6wAtCpnS5zCt88/p
nZDRFmHo6oeomCdsv23+jVgiYkSz2kiMPuThaQXDbvuho1eNE+YsRRaN4JfZol6n
y/WLwKHAqwLcQvXBkySV44rLNVc1Ltx1dR+khtuPI6veksVhChUgw9JmLYOczMkp
xr/wbXVtEKRdXsWtmVX01X0SGovmOP2EphbozEkEykeVg1WgymE5o5obO9bLZ43o
9puIh0ESZaJUuRCl8gdVgl7K0LlH+Moc013zXwXOWTe6aYPOtevcokdvrNvXFRi4
BMnoaZSjcB8EHF3vedfml+d92wxtLhZA/uLTiC+yym0QO0hn7eEN2x0B5yTRFZ8e
ALLnwMoQxifyV/y3fTmEeEZuPStHV+4zTnY8VuYkPTyOdq98xlqR9IadJHlEyX1m
hJrxTOucPHcKh5LZ1WOF3u7VLKs4b4xS55pZFk+ccLZzdE9MhFh55Zyo5BpDJM4U
nM7V/f1aLkRSOjR38rOrIuM8o9q+sNZ/1GYfJpwRWsvv48RqSjjdWQIQaLt9r3fL
a88beKfyN7YepCcypJWeTJvXhAJAxOePfVEcqGrpKMNWUtVhmuK+gsZ2IN2OAEM6
dixDl+3qnvDWt41iMXr4GXnLOL+aLtcNxQe7OiAegbL7MPq41hBmQKK0gVjLwSe1
mp6CpBHnrUOuOxgsKFpBkkvpzZQttd8jxu1A7xrWEd+yj7aiTAzMPnrY7T2fOepo
UeQ61oetHJ9D+OuaHRW1OCsTc5G2MwnAB2I80i/BCefx1vST+2M3WIbiyFlBAfnf
+ru3N3jh79x+jczrAkFy9knGpU7XEcCG2slzoPXXH+wSWd8UWE48HdcpT2zQwqOI
pQfVgVZD2EBKJ5UTW6F+4dwWLCBwA40Et4y8TiFStBND5S9yYZhrNRLnzHWSwzcp
06ST2+T4fqT2T1qk05Ex6XBB9YaPQ/X4MwZ/sITAX22Xddcx3G8J10xil/QmZmhS
LPh45hDkdMdG/xuWFUvS58OgIy/OfD3r4KznEWp631alKlk7SX4pJunGXYmdRVal
P1CzoLSMt3bwvbWZxBabMpQHe4GYhPbQs0pOaLcNLEHMnxXpoBBmiRQ15spCEiL1
spKdw79aexM5lPDiB6drTTtoPiO9LPR6Ao4DzbAkT2kVXa7OThcA5EfAxPGzT2wp
F0+QjtFcBDZC9V1NDZArKw3G1H1ZHMVm76WxCt/u+cYzie1E3q5x+hbYdCPekb2b
jeQyuDc7jhnxRGSPd7kCyMAWnvfBm30HM9LJMKy8+NqhuW7FuhfuNeTibonGyzCv
wvUI4tI0b7Bm68mVhNY/eQfyoVBW6BIPFy2pMMvY089uoafWZXlfj6ZjP1avzIFi
iSDJ1nczVLTZOt9dRN3GAXPDR7O5lcr08fNmw8FiyI1lJlsRWL6pgWNNAiHawBPH
iEJfZAVw0OeIW4WZihOIOwlSqt005TVm6vwn4TnYmezap48WBfZ/WYN4/fubUHZv
Rgq6evZG+EdkKDrEVUx+7Y3Shg6TAmgIv+ecxBlJktbF89jwNMEmVlFIupc6mJib
DkTXaTtJn4okut6w3rlzCX+3guF/o+X7eXR/dI6h8xMkmeoeMj1e5F4Cga1yMW78
RGYQLOJfTyu0f+lU2BqPaXSQ4mZ93r/qM3Tt+EccEWFDWqvRw3SCoNaYc64b/cEa
CqicSFf9CFqYH39xYfzElrle2PiYVCgPLI31nB4ahkiR168L6OT6hXYxE/tpdFR/
5jOLSlC4C2aJtjdFBLqqQYpLjXpdbtOKjnKu7IzBLM58xmTrmoeEzBEXo6Ym0gpb
VgHdvctCOBv8V4bmZn7SPA3E1Sj0iNYoeLqvs+dc0yymTUgt2Gtt4LiDte3UN2bP
3+20QUa7SfkIDlzLP+Y5XGKsT3F7xnmZPuQ728mX9LlMfNRjIHqZSpiXoV1AhtGB
ehl92WHxIoE4kWt4SO3CEwPcelOuL9uHIR4JlAm+G7lrmX677osQcm8hrGLNeI+O
Dovp+3lxRMJq9GoQHkXYBvc3h1SIIR1VVQi3m1geuQvcZ/oxosCAqwixbMvO9ymD
aSyJsiH6/wZ9wRfd/Y5rWt3Qejo5Q8A3Uiuodl6wc9rZtPzxxLPJDaabQBIYpi9V
WTPSDg2GdpHfvpprT1OV9ju/HkgJ8aB56QB/yjIZ5pXctA4FvqgS/HLciUYekTSE
yQAasziYj29bSPeRnT9xKS21AO9R7AiYfH9IHm2uZ7TkcgY9hfdWQdpHiLxXiGVH
qlFaD32V0hfxyDOrrOarMP8VF31F2Vu5HhRJw0JO+Cl9dz7adA1EKU1GsNd8+0zk
SVgcHHv75tvLpLfA5w/8PsL8l2BHTMieSHzzZgGsoZTkPxSsBcvKR9CM54R5QI9p
69tkFebV/kK0OY55uqIsC8J4cshDbfSRZQInyUbnclXDtGHjygburBsniRDyPFIY
7yCvLG4d6fCgm0HoZTrBeBmF2MmyJB9MgSsC2x9g9alUnztq0K+LpDI0Vp3lD1iM
vKXzmybbeoitlmoKzGD3stTfF3N70ZJc0sIOv6OYs4BzgqcIxLTvjXx7ktD5WJzv
DM7Z8ttlFWaBWrqdhtyZ9KLS5jeKwBBc0W2zpOxpBZUQ4qjgtNAacc2Gfy0fjxlj
XQHQBNQGjEd8VF9UbPFGkxTawjRG8vCsWJW4xMbNlWusLCTfuuOXbDUkz9slqItx
eHa4e8qFEFN6naFVT/DEji+DystoZCzOwFFJuJMqg10pDlAw4wLmcdyCx5Jb46pf
9OwzHv2R5M51q5o9fYVWPEloHMykJyu1zYVdx6sDLGPcExg1TT6DctvllsDuD1Dg
6gMWL+eXVE6xEu/XjJfpbLKWwwziSmWnAmbbtk/FJfZWzhWtDP6Gsnu9QrL94l4r
G6ySGbyO+9gZuHvxJlTB0eEpldFHtmB8j2P1TAY/DlRoRqEp3Wt8GfeGP64X3Qns
aM4pbzfftCrtI6DkIVAa+zzc+l2OPiKsv0bCu6zQjMqY/YX8oyce2xOCtan7qjB5
qJLbmt626lQD561gcq2DGabOY8LnmIG1aNbwe6KO+/bBR1/GLkGeCkTSNHruMnLH
76jTiDaw5ZkfPLl4LHO/2bzSPlk6ECBpPrJGViTY/Net9ooFZLYcWdJlAD6Fd907
hoP5whGKcgD1rQnaAts2CayRqcGIH2ZerF9VQvrcjW2UIeFZiRu1Q7MOwX4n9Mmu
bX25dDB1QpLlrkui5C6tnAYEcKrB04WtOH4uyG05jcE/lRgThIyaVFHIku2JeaxP
Eu91f/uXfzxuNGrNZrX/qmu+1/yXb3cbnO6QOGUb1Xi9qOxvNURbZrYdtIql7OKm
ZcTupm62qIpG5mbbDyTYDhhxW9YL8k9UloDyk9vXyQf90zBFr8WVle1Ja+utFELs
tJT8aiPXXcvh+ihvQOK6pgrsH3s3yLKYKyVjEnfATlRNdNGsYRqWm1ngoEXGRWfF
wJi7BiCmgDssHhXhJTlqIMEZsBDy1x5fb/21Ltt8Urrie+5XBNsk6eZWrJXJbcuW
2w8y1lJ0XEoJJCMO9wdeXJpOo376b5Ylk7qxuVgYoOo2/iRa9HsNOZh/VCgSImtu
9W9NOxCKO4i5TiHNwlpkhhtECBsqul4yDUyUQOB7GAdvMxQw/70zFyAoY99ILkvy
tU7C31WCwOGw4ANWYusnv8ade+uFyT7axYCt3cJq4A5/GB2h0Zp8uivFo2Eu0Bts
d6uI6MV0c9w+gD46/hckfLwBjX1m596gYh66DlKsp0JsvDUYmf5ZF/W/okKWRWXM
Sg7OnkHhtVqsTLcnTQNN3+2XiKLznMwe9u4qO3Em51RssASwa8r8PTwdhZmq8/FR
PNmGveZIWZtMw+nMo73uLvtqxQNPQ9gyPK+Jg5nPFNflkoIbj6+j4JSZcaQXryms
6HLwSJpPRvD9jfTFvPaEG6Ii3HV1O5gae59Q5gKtPt++QmatNZZM/Pdu1EbsKYI1
VW7jiUWOVqodXkhQoTMCtycMFIoeQC9k5idzJ+QrAbT2UqyQ1KpHA8NNPB0wQ/C+
MFPzdO8oMAzRKwOgZYGJIbkoPOumD1MbofIrTqUysd/G7f/x53wpRgINA9gWmuVz
uiNImrkV7Z/OOcHVF5pbhU4thrWrULR9931aUq2uc8Zxj9oG7oOnroMzy5UXq0xq
q9S30dHOW7fVmNdr2dl1pGtwotQqqAqFDqkk4cofp0HTnfX5hKcMROxkuygIIQeQ
49egbb+L7uyU2kTN9ZHjbfkcw2emPS05rN5+3xiVWaPOOjmYZTJeZB4TzoplSPa4
xMvWRkmlUb6aCwiB3OpJV5pYJWS91JVwMVx/7VlEA9gHQehBR1S9UQsCIEoMYyx9
HiVE8+RVXwEUX5g/ufTWgx9rbOipeFktlx4Xi9/7z7sljDX+j9qd0Mj9Hr9hnY2g
g5q4yknxVv4U/eVyaaKnQjuvgY/T/6Pe0lyj8VPcrGCF3QJIu472Fm6WuaCyeD8j
H3Wjtj5svRPnyTgwP8zEQSwHveSfCpnLV9cbMCN0X0Rk9IQp/wlJHImIXfk4TmdR
/hr//qzLBMkr3nxnaCJcv9rVZO/G6Eyn6eYBubfYUR5tbgVEzDj+xvAxcaTdhHn6
CENjHltU2FcK0Gc7WdGIM5r7YL8drBW7m4SPI1Wf8bScMr4TzZt7i+8kraQMHuiI
tLvq8zpVZch0MolZYbSdoDMrbSMPP3By7U9o1mNw4J0xoXd+l3UeJ/TbT9zjYlQL
+JZnlnIlkBfXf48JCErXmhgZVoGsndu0NECgMDFSFXHPT2cpmXlp9QoaM8vJzLkk
6VCfzEpxcfBMDc0hJKG5CC0OwyluIYkOwRCzQ3T3NXmTbirl9JJtnG9dgMt4CRRA
NOGtqLQ1QcwrH84Zep9yN6TwMjwK0h9jHnRgpL8CEI7E9s++uUn4eSD7Zq4JlLUr
XW/5YqoFDwlkDGMFHPWXzunaJCe4tJ08utgvHGwgMhhPSViHd8Txp8uPxtB7qIsM
0E9PQyY50ZUSDahxFdWXyp+8ab+zhiABtctZs972oPdvpRXE42h87UEdZSs+wFRm
+H5/T0PP8rX/DyZ7VSwdSeuhUcJuQuRmj/wr7qG9hzO9dk/2s62HBqhcv6hZAAgk
trO20Byhpt0wxZEWJWbsI8uT8Bvmx0YGqWW08YL3LJA8YnonxyWoJEcRcnQuZr6I
xs4cfVrljV09LaC3SsKfd5w76Qi9aP5RAq+2ROhD49i40I96c4jK2e1Bz0/i2y4F
03mbfkK9RCuu6Mx1nfJzp3U1a1aUhOqwymuQYHzKLYNOxzHFZD6qV4V3v73l3qIi
lEUbnKTksFSzObr1flDU/WEaNwGDPYhRZg5PyvXDp2E16bzzDRPH7ZIcW0U9dX72
J/fnV3fMAZEdaHNuQFVN0u9diL/j6uCipRE3+/xpOtbQuoJUjwbiFNVYmJGwYe6m
CQybllQGutKt6/gLwasQKBezvOHdRAFhNQJXk2FLMTXiZuA5MR3q4vqEYmEnx8Px
qQVBhxa4FQspFtCQrnLqAju5/7QIK0ZwetqBdbaSSkWQAH4ClF3ondNte8Cw9TsV
rSVl4BuC2P4nIOxxL0XHlP2zb/cYlrCf1fUFmaHiRzBGZkYAepeOil3A+erjV8GU
KeJToklWgJ5Hc8y8Zl75Go7Rarf01ioHrjf7wje6mjnS71raMyN+yh4+QAeO8yh0
MGceA5TW8/lIPh5FHe2PzPuDAWNzsHU2ab9xJgDsb3RP0iR8q5Sen29/pWBesVk4
yWclv3sDxhhqQe9V2uLyKyBq7KGXbWF4zO2RZT9BYo2Gv2EmathaBEX3Urh8g168
dtUbH5xJB9NDPVgZjECGbPlGdUBpzqUgLMLQGm55XeYs95IjknzD6d+TJgGH+q9a
4s1AS9Ga/sNP9YebCaI0LG6kkkdjSVcmvir7xzC4dizmZvQMuWH2DOPNlttYWo8o
loZCqig+guIXY+6kw8rSnvbBZTlNy+UULcfOKiXT7MEbAGTV0HCDiANzlGlNXHF9
FZwWLXPr2cfw54++8Te82sQ3MQE5sb0DDmaNnFUaH2UypJEXVu4UtKUmQd4bQENV
nrrkX6DdJO5IM1j7BAa9fZ5LIKOZ2Qp7fEeE1WQa5ufhtLQA3BbHOVEjz0tmvYzj
fDHMpgbaM+xm1suy2FoHgIGnjrCYJaY8eEIue9pKDTvs6vXEZF3yyhJ1dr0gMpFd
wnhUZkaeS3JTf50+wicvgiCQtPlsq3fBRwFGP9Hrk/BTEnblrrGwoHAxTWftO7uM
HTqU6ClfeGN8wR+YEjCKmvE1AUKK+t+X8ce4hNBG9tSNhFzLSyjZm4EsRw2h4/GY
HaofbL5y4Zb7uRqrM5JbzgPn2XyES29LW0Jix22t7BaRP/lUBLh5v24SVjUXnElC
Y+ySLKKmAnxVC5zNKazedt4HAu1eaR9JhQC7IT+jm7kjWjWiQsgooSk78oRUNsgR
rKjUW3MdLhurGGqtADhBvjDxD3j+1TrTHjP9ZYnVpQUxOdplNFmDSAMCx/kz+DdP
65unCbnGbgBv+/rJn9kEE22HSMpZQMlRYfZDrvug8pC9bE9KM1Wbc3LpWvT5OsTh
rd55t43Z10mT274M36mY4MfXFH7TiLNmP/77dJIPKBfG1/nl1lXhXIRGKRcVoA6x
n+7slAnigU+vUrxx9/mN/VYTOvtRNVZnVagdffblYpf4lm0B8YLUo7Om6zCsl3FO
B9gKhdpfmei3QQ3B3XwKAajtK9E1jTcKYGai3+Es6jeXfEVNdnrYpUcxtinu2IAS
Cqzmtd5cAmHVFQOGShHSeF6NGYjpyIKcYauekz2ugomdS+UWpYm6N9FCpVVV2vTY
HIFLMYpFyb7J9tH5GK1/VjF82zDb3II+OjOqN/wlKMhL75VkZCvIfsoiG5RWCnQQ
alTpqsOvCU3iwFtcuPQVa2MZc4cI8BKm5MP6kaAX9TK4RB9rtjduzxuvmNvtTf64
t0IpLMHaPM9T3+25KSuySN+GtlWN12jP+rcrqc5OnEyl8IncnpeuZhAjW6+U+w55
Xb2qdKkpOwQMjDZ9Eeqf8bgd1G3+ZI5QD3Vcz7HUzRev0TIG4iLEUqeTnFXYndwo
zxrK+eswVbbnX5g53mbTZ//+ZCfhVM7zzpDqwtecTxvmNMWuSCZLHDuyLlxK7+FO
OKx+c7ehP3/JZr++gyRTzzSka4FMkC2FYTRJoYV/VBOaFQjWrmh1zl/VLgl55gvU
ywkvuHtiXDKivl5hu9wXo3JhpFIKD9x3mTAKRtAQAI1iUi7fLFaMnWlw897tGL3s
MK/WbDOYWFmmhrIBGvZ/9kjNqYzWuC1tTU3/l8ZKyWjTE/1Y4//ZsQUDzYJCXl5X
mWL70PGGiMIfK3orK75Z+4j2dOZeA5t/l6tf0gE23i5bYLvAKwF6JTPFqiHSh0Ww
XvMLMRP+pOdD3PzQbGfitXIQ6+Gqgm9xVtoSZc2qejZ8EE8Y7IEP3wqbTKgbaNY8
5OUNEWuU38o3WmW8YndZbPnRteR98F9VQTRDyhRGJP0USnxGMQ3vlcv41g82glJb
s2E57SA0OIgbapIzpGN1eerUyEokAMqvmmPSkjqyjxDcZrb58g8TrwzjGlualFab
NfznuHDpwqnb6Nmf0KfzP9S/pKYx3pBqS+rrpqdELJcj2lkDPkYoXpS1u0MAH96N
BA3C9fLmvu0fppEqfR6C70jn0rvCJCdOTPVejl42OBahYQnuYRij4WcrxJ0mCV/m
UJon4be0ryepwGGTA9OncT/UNVJpz7opb75eAH7d/EfOSbZ5S3+QDNK35YIS2zYh
9pHOa+OmCBCjE/YzAuv8PCcFA5AuSjkXZhWfrSORPcdp1A7fbzZJyKagLx2qQHqg
wlcwQJpCka5ext5KiYFHZTWtD++mE2gfZRWcctZpx+a/Bjig0Vr/bhO4GOmMdO20
6HaklGZ35TNFtk1pSkkaYsj+RXN1cgQF8Vd0SKBjbYbEnTuzwSQom+onrVpKguVv
HLs/YC02kPRoZudJ3OqE7//9ySZc3mQx7mALqFNWzHPQj411ndACK+lp4Nbb+vfm
fTSom7I5Opo/KBEelO8VEwHnx0XmxhV8NO3bTwxD7Id9nd/Zof2bsXr+TsPz4K9X
xoX6Lh6docBtifISRPX7ZlgqF1RFSWLebyMMuMBdaxQOhKI3g3kR+QMdX0e6oz+l
+c7OdZXArL4iwk/P4rSxzizpZvUkBb+NYlR+PdnQsdH/l1rK8qb/83VWR/gAuxs1
daMrLcbrZAM/smVjUi36MXjQfpWfW/V9MYF4XCLE7MpHVQNbHcRFB2BFxPvJ2DJD
GFvK8ZCl+qmRMiSzWzdwkjgPDLPm0++4/sIT/wtqnDY0gnJQb5Uw5LHuvX2KOtlG
u041RciQ66uhTObgjHqP7WgSoc20nGh5FMYq5AImjI6jnDgtTWaiZ16TQ92jyHJc
n+RmGlxcWrxyAxp1ktXLOoim0Eovmkay0BHEdEMrSAlq7tcJp/qYUgZMIA2Opkbt
SPACFHHByFEJjwypy49fidSob6Z5JFZaNA526AFxLIVi97ajDibX6Ip1GaNL4bLV
QKiJoPRCr4GlH+GjVukI9vZDHlFFwkdtQtAFY1G3aBAifonNwJcxPfkMMsAM2+Qn
i0LcWrdV6tbH+Npb7DXeqVOQr9G/WLkE3ZCh98r7n4A1BhdCVxNQcnmUJPa4qkiz
gKMYCbgsxsK/pxPAWUsjCCMc0s0T0LAIFsDC4yq3lej+wtOZH2kYowUDD2OfY7hU
aiOaOq3mO3+ifvT5ygSJaqF+uITi1aH+vEm18AHjRBr+H0dvnymTFUjfFYZAofxK
mFRjkqX1tCFJJDabun58r1hnseOSddhXdpSGEpZ1C4jPcVf82fDzzHLFJPdviGCI
1U11Nuw/Bx6ag5RMaiFEa446rDv2pW8G/EEpgA7pONP2WUUjIE/UX4Q1QZus19a2
cjfDmfQfviqiXdNy8v0HXnpt9wYmlG8aZlr09ZjfRG/hCCynSpC9BTUCXA+8D8AZ
W5yl7HwEMXKP5QEvTAWNxgWT8DEUIfGooMj5zdRSBnKljwYLnGDeroJbVDoRc+U9
x8zjKLPGAdcUPSciWnNbvNF28TpVFcKi1o9ukuf+Grxl9l0ZEcAv8oC7YXOjdBTq
2V7v9PQTQS1nRzZDQl0biBFLe+5xNYBNSbOUHU3x1blVWQnW9eqoLSOH+9pkLQPl
J2OIElaacB371frEZU3Xl7A7T1SbG3uGEWgsHs4griK6feySPIYevQEoZm4Sxj98
8YiuEFLsBqx2RfcLNTfEdC330LWPPLvv6Mx+aDITsOmGR6WzN5cstvaSlSTC1fHw
iB329BScVKiOLnk5FZ2nHLN1zEmCX9z0eOJcceLdycrm4fnWx6QBjbNZoMp3zZgY
5QAmPNm3aOMKKFJxe1EYiA3YP1B1kcIicaUuccgfN9bDO+oPEawlavF2+HTtKCvY
uN+VNxDxLLRn7i9EzwjrMz/S4ZHbGj+C19JzhDDkhuqZ/5E9Ix9aMkkqKnH+xvz0
qXZhvFdBC9Tfs1ngv6Zd7srAdrwk3KPvyOHYtDqVgJxOilSHrXBBQio2m2fwhIsG
+PQEcT+ztz09PZ/YsLDtkUSaES9DW8F0T0HIBRHy3gCuPAELBJLRRT1FG6eYnGDB
s/IqwgCtIYgWtV0vnagesbCYBVb3j1iPDUYpo+AmTLGsV0qIcAsLyeKZWsTSv/Pk
Dr1+F43F1seN61zQWNY5jrYHgzZwGtuDxQdzYbgOdtR2ODi6aCyungffJoNSG06t
MSpYzuxxs41hc+hZ1VvzJfKQ52mDjD2jMrAiZpPnwfA7nen8MgmjLb5Jq+aR0kjt
Oh/oq8injr5oWwnHFfdmPfeLeFbw9yBNcMXLhSP23je+VK8j5KDT1Mk/EhDwYtEj
HRg28/9QAkbqzb3N9WP2/nTH2whoZOuT/8qASA5MLU08/Z7FFyoSAjOzEHZLoCjC
aYKD0YWQdx1b7QEJlqloPg9XJUCRgJYkm3FbiR2sYW5Tg9xri8c+Bd7hXAgEdb/a
2WwsbIDaWb9kaC0EyA9hwSKvfgQKKtzebeAI+CeOgdbzHzUdBj2ab4sdP3aLJseX
qdSFppMUjMl1QxZZSwOxCaAaDZ24BqvNWapo28z9s2yw70HutUvl7NpTJ8F2AK1i
ikMQ7AITNuDbE1rj8lIIPX2W2tli4tiKr/tG07jYTgAXDb/rm0GpdIMj8RQPaQ9e
ifsk4uk312D7bMOjSblp96JdZw4ZUsqe5Xk+ls1LKp54yW0X39JlbWeasRWC9GEG
WTUsIneM0QviuLQEmq5kyBEN6eZdPEFioYgvf7ZXdMINdm5mLQ/Mg+WWg+Yd2Q2i
nT1u56yPkotGrthmP4yAvWFnipv5XuiqD7bFiAziN2Nyl+Cdct8U8rR0UntCGMss
uxAs+jPaHpGLWTQQFipNDI91vnLwbvK/flYAMAOwoE4RDDHACNWbmyv+jY/mVALN
Vz2UdCvxZFtlXyEWeUK/jTchRH8opPDEA9dtn/FxDKjARuNnBeLP1BVUCcGmHX9V
r4hEE5soY6aE/FHngAy96aIhHpog9sW9Snteu7AYo53IznEtzn2RKUGJsEMm4UbI
NCNrMfMhVD4jTPAWQilYImm0sPshP4LgacQTxuMGD4huk5Aghcx2cVw9Cn0b6UfP
QQgyPn/X7IyzPbxewGE9tz/gbGSpoIwcig6j6D2R3HQ04PkFJe4GqSEG+h+6pY8Y
Gr3cffS5rHVIH9+hLzYTKWUwYBJJC+3OHhNE35BRQ8hBmMezUEkTU1C3EFKbPPZA
xu1wpUlvS0BnoXDCTWks3LeBw8wEak53cFatix8jOvSv5mq9k3nwAEbEZ6F9g8sA
cv1i//JovggxjEIyWA2qoG5mRRthUuFskl+SW8ttmy0nClDw3jdQdq+WMAANjnhI
ANbO/CkwHvWnMwMpwY0pY5WqGw1KSpdYo7FFTHqwq1YN8XxwqmkAKsFtnfGbC4V8
Lxkxg12d8MaHiaRMiUfT6uERMiJLg6kBE1qz663UUsznX1G5lkBBWJai6exJXpvL
YZCmVk/MNJDUaZuYpWpH35+K8Eb09qmQoHkF5b+u1jNqJOwOy5gm8MulCClepD5V
eJ6M08YGvMmsOB6tDs22TgHZ6AvT2RCILtkACrZheIouEZ94Wp3PygmJ/4r/G4Sz
VGQarRuPTcmvTNrjkf9EUvzw0q3/lInEha5FQmSmnfIWRTLiMT1B1SpPeCq8nUbD
JNqUz4X8SK04VhBzV7do2yZ7CMPASdzFlhxOE01XiepAzFr/hzAdJ/WTMkLy+0aq
eRJEg+SiARUqd3Z7Oz+c2/M2pNmCDe/Uvj9uKXTqvAD0bKgJOVM1wEE4yKZtSTmT
xpzuul0KMD+RjoX8YBO/uLrqloFxUehSkWxfkvMWRBRiqTNyhLPw+u4A93PnfiF1
2pEHn80a0qEhI3411xGE/YNGjM8YL/Cp6IPNXV1ZptqsNoJHtzf2BxrF+2OtbeFI
IOxqwM9AAfHNFrTTsx6h9uOttNTCHpNQ5o1v7RYq5Kt6nFfWcBrcofYxn5UMxn9c
Q5pOEkN5bCIkWq0zVPwINTqGCE/1n8Z6z/WBBXij+Y9dLu4IK+vvPdInO1dKbp74
vpY6F5GhEFPLlzE9rQkDXKOfenCUzyG18bwRZruMVBBs0uL4DojYOFrl3bX2pbtt
0a31dy4qaFHM2BkND9oElSt6PFDLgVvZVd28uaZU2KlvZwXZfGula6rMuOS7+qqq
LYDmNe8F/N3JuqLAET1HdTh/TG7mgCTsJ/gwgNF8OQDyLGJX/C3gmTRTzUSI9DPw
bKSZjee/lt+W4rinhhcqMd9adwGwiXefaimEMSQdANVm1PMfiSl1oc5hzKRRC/6O
4pw/xKtqlP0afzeCoFD8HKpqop8zsMziGMoDqcuIRDIXRa7wrKbwqXZcH2L9r8gv
ZnHzYoe21kFFeV929oP/7A365Lkkr34eV2od0qXiYFbrg8G7+EZG0xG61W2j0ITQ
OcS4vXZLR+PMjZKTYegHDaDtZAqr+ACn/uZWcET9rfbIVB/rpnVijeQD2HoEz7ig
xcmPIqxPt6HML5dcoQQbEkJbchviJq3rd77B4f/ewcchX0LOFnlDLwL7CXIzTdXh
kyFoQ2wgC0dEWjghh12Z4gWEjFEaZhcXCRfYZ0/cyGK4r9ioGSfkELYEjrQVvC66
coxnOUEDAywZAtuh3FSoB82OIqcuyZDSDmHUM3FZr1zz8TIfCG8pxpUJI6zDk5Ad
+/GWc+nzIJX4uxZ8nCmYh0SCSr8XND5eLc7vm9ztnu0v5VCMve5LkPqKnuQQjEis
80AKIM+MBM0oi59lu+OYELavFp5amDgAPVEcGZ8/3DmIX0wQyxuBC9gtwUI2q8kP
fb9lpUvO79Z6hmGDWfExkXZghCMEh1YXW9s3Jx4+ffw10KFuglww5uD/LReBQsYV
Ms7Htrabq3IW7H0Iavqw+oxskMq9+NlaOrDDt4gzVJHgoOV2gP8sqIrs8Jpvxonn
eRrGjig9QAK+4+Fe/L0aeA8qMsPqT0n0zIMimIPBPN63JnCSMVpYSgPyAxpM63Gc
4B8v8B6ZowVz2DNqDzOr0w7rb7GV8serr1pOlSoYyjQSN/Of9/5svrVMogCSOEsX
9F/vpFEYbDeCZj6h8rJKt7HAbN/IZkpSVrSuXNDg5IefQXz+6vPpeY929oq2jaQ3
v9cbtH6TDmxBWx/01EG3cAUk2SMlCJwxs0SD+kMvCa+0qb0vnQdYBQjx+VUAaa01
AuCPIw+rVUmR3Y+Wyx6h46Z1mhQvDPT/ayec0xhvDDeiYG8v8tBZuMVmn/eno6po
66nsuIIMFYZ06Ipy5npWAFuhfFlF+5/8ibV+9nCW4qj7BqUSrR/NSYcL7WPC8Pwy
y0BG837/OWPlw1a2VjO5zjsPLhDt7qBdFC/o2XAWvI6ootRjSLKXaYtex2Ct1JdG
2WIG6jyz/AbCe+6BTO55kSFwWb1ALVf5KG1mnM+8TgdXQoC98vLkGLowoWZG+t9S
CcV9gttYe6kNa2RhtTyN2scYNCf1GN7vtuEG4sBPa1RF6sBdikSYptjsubkxALyj
TQC5nMydLpYXDUuj174+OU2XumcUFdvRjFqiDr9F/QsrOp7CbuZdNcOc/entKr5m
x4KM3j++rPKEtPQdk+DlWNO2tA79T0+E7Z3REr519hkkn3QZt+kbipbHg/MOMTwQ
y1cOu2L628Rc2QlpsVnSDQ5lQh4wvriMF7RD0ONNy3QgkxwGK45cy+CWnDjbl9Go
cDczX6lPNgv4hBrXKFJxXvfEBlLZugslJoDla9ryUy1RR9yT2FYM5+58X51MCrlq
Em3XkM2cwup5O1VJV/E2uekKGEXg7Xt/M4hiK7BHRbRw+FdgH73ovSQicjEslIEP
CGQ7orOIdNfmpICLed0YZdSyFtLCdr0qiLhuwi3VVdOlGcXblYPZGHizxLt1WsUo
TcISkDNm3uxQQl+Ns5bKiUI5YIucnAk0QQYvWD7w5mfNpLf4vH5Q25rPCZlGQgqP
BPUz2zv4SeJ+8yTi+Dwu7SjZ7gADiWcjb5//XjN3GVEg7WH7N7Pk2iq1ZcE0QH/H
Nk3t9KVAowUzjaCIwu6EK2xdLtsjCJNzXfx/EsMkJ2KQQP1hZeJDkkNbEvXN3PIA
91Gcr2UCfz6wpMDoYsd4yobd7LLt4rNDpOCbzBNcnRkGtLM3mvypYAb55/jaPpcy
6JvBD4GDP25uU7xPxY+07UQaKQmLy0RjiRL5Ubyexu5cRTaPXDqMS/dn/t37uP9i
Fe/2gVQcpLi5onI/CSwqJanyGNZsetebvTa9ghUlM4CD2NS7uQgXGqBK+8oHP1zw
WJYg5jbDCCbLV/YWs+VjGjfSaxPvHgb+S/AVlw34hLjgUnYnPLUh1v4Y7PL3ACQ1
gwc0XTmI+ESOhByM1wJKTC5CUAIIYdvWdFkKvwL3DYRZWgMJlcEsBveZGvG5vNaW
SaFkgzrgkIgPui5y2lOcD23YbgeUCS9wQv7C9bbLZmGptdWEyGurrqzj3sAthc7h
NL4XDpFZKsVDfx2/fiPnbUYqbNQDHlEV6GDVFWstPmpw9SfDBj15O4fM0DHR03ta
xXEgbekmq+xgwuJaMY56WWOX7wfI3whHheIshe1D4UoMDPfejvFtHXrzhcmNNurb
6XPoVMrlNmffjgEKsehSgbAmLCOSsOeQ/SAH1pAXypd9Nwyf+3s7d+EA0KfJdbcQ
lZq0cLScuUvtUN51fK+SiIZK9VKiI+QP51P83V+UldK4vivHJbosOlUu5JDH8x+t
MkSM//nHGtFiQFgvjfuxCeMXTSGYfdyFQLym6BFPk7N2JKcwt0eEl2J0BcV8MWkG
kfIdlq1kJUu9wz9lq0PTK1Gdu+nmMkLJ3B+QtxB/mZLCGJAgVcUuKn3at9eFDjPh
JCWk3HfYlRmF2kwgao6dGS1b5b8dQ63alibNmBbiV/uLk96Hu63U2FAlb9bV1VXj
XM+aJlDtpdQmA+iQwVB7GcxAMMFSdxgGMpgCHfpStJxlGHaVqa9ja08QYT7cJ6+f
NQu9IV95KIgCOapNvZ5vWDZdo/Lf4um/iad52QnvoK0NEYeRMQVsDbVcAYNra5M7
vRpEaFiRVu04tdMCHT7ytNldt8Qvl5As8QfdXELLIeWSsXqNmNYYCpbJ+jkf+XG9
ZCtUYDKYu93m0lWvA9U4HRS/V9ZNr5lioevJu6QmEVU210sMJLNe1qdUkbqwX4Hh
6NYLj14TqHuCcIYM/ktg32ozEPntMzSPd0YqFYveFfJ3iIrGb2GGyq2SdoJ5hOED
5+PXB3qBag71IrWYSJTHZKhrkKHZV2VXCxc8O3i/aesXUuMB4PsrAtsPnJPkD5j4
cYAk+xqieUN7V7wHh/aPRZspbswdy6qP6F4GZRxxLbiqfOkerhVUXyVFf2LiLVhR
eLNA0hNUNHnmIVJ77g434PhkHVEB0IjhGJick1GvmN3DiFt70IJglgHDCXlFaIna
/GpXtHayFLs7rpHBYqstSCOtyXus5Bwk7na/+BUzXrt5LeBBtfZoe7c42oDUmebi
r79AJNgRpAzbXZYCOGLkH0Kqbj4/OvE9JDDj+Y6Xu2IKjAv1FzWpNFXYeSLd9LXj
PVxzAaWgr8aTcZRg/LDU9O0uZEFwOdBGF9MuIunByBY1fdeXj79yjG67wOCk8hyp
Z7GKbuPl9EoQei9CtlcY67gWbeqzWETrF+BfdBFozJqzuNo75jJ6tbov+7QFqtDA
B7AVfoSwEyG1Z2dkHwJUVUOyRz0SAclXw1NCe4Jae9RT0HguUzl7Ex+lnLjRhJsj
0X3ZIp7axRTNQT4dIYrNBmeZrD44MlKjwshLtm7DPI1QIHeB3iKOeOL/8VMO6LKN
bav/yOLMiWZAbC8PYb3APdwLEBBWcgNA8xyXNoDtpTwPs38JfVuVKQiTZsGwJud1
37qB6t6dcdEfhOp1X/qSi75jzs7b4inISaFqYM6+L66HYEtU6Lz8/5gmqxPleUb2
2vd26FXsUJrKE7+wOpNkuV7xQSTHXI8WFiMoIHzeMtdG+YPvMlpiTF4s9QVt7xLu
6rROYrPKy6yAPYRMmNp4svdm1hCDyPgpbr+pVfhFlWndVlfhwFVEq7Sc96csG440
WhPlKHN4ljNkWFGhMHvYifw6v1yPAZDuUKegwmJ7WXqIZDdVqTy8WzkblTuDZ13Z
7aTblQy+bc7UuByBNfHzuV47zeD2SewT68LVCYUTuniQbRKAIyiNU3JJCsbNAT4n
zAqfnfndj6gOF+4ZYZNsIkx5lfW1NogGW1F4JXoby00BYUQPJu14xsApmyHmoAKn
mtv4uIxgW9T5meo+SwQeWcLFlmoA34SbWR1mKRtl418SOzGk09hwJzmJlDV/Jrea
+YpiOOrDbIyg8jPkDrat+kiwx6TEFJxd70QxL8C4o0Ty3q2/n1Z/3TcXWX78QHtk
e4Q47EGLZk4kO/l81Nc66FlKU8Tok3qnQFk8d0n7e7d6iLCzoULPMhHpMMIkqOro
Q5ShPdQXWXMxHjDrN70Pa38Mkok/xjI3KvBwzAYuw2NwnRQL01+GOnj5JxfCMVxf
8o50EFx0KWjTVy5eTfBTO1HxLH2+zSa0+8sxGevdmX4B6da34fgJPEr8msavRAQQ
F1BmS2p/NHDi4kQFjL3+tFQKco2fQ+Dv/Ou7CVkppeQ1yB+h2UDXYYM0jNsuYBsn
TEhCiq1lqE+RcKVTjn/BQAo1zxV31T/CnReBKkbjAPIW5/0kcheQmV/3zXFHvgLl
7PIcfTC+TppAzZSQoIgByPwD5VAOZAwh9/8b9PSU2ZELMyrNkSbDCUJ8BcafTR0o
lYeRpV7CIXxQRUG3AnmEBnwevQgClN/X9xg+n1Z1tvMQUfCva4UsSHfKcjDxQLBK
QIe0iYiAWyFEFepv9YMvrT2yg7nHHFZ8tS4+qP9kO5AyGo2nWPy0aiCtKeQPFvcM
1XjEiV2v2n9JVF7f3CRZie/v1NHT/epKQ8V6/pPJn8yn0g/7gO4GomsAIe2MYGVh
uqhU3dFNNrHq85j6ezD/SJivwk5pw0I16vl8/ISkcu16KeXVdyeLotSavBED/d3v
GpwXT/VKISfba3gF9zKYifsHCDrVh9iGfJUUnpnPw5cFOCyqae3cDyZIEetBAtTU
SCjpsFs6xX3WUk2Z2PiM1hnJXgp63YuvfJ9r3YbTCWqXGCYgR3jzgNbENyj7gUN5
qufLgLw012R4GG3CXPtK+OF+phoIJpHL10QfFBRzsjpxwndoxkRy2nUqN7AZ+0CE
fmRKDgKVabu0gMZ/4awKkD+bLpWsulKQi2zyUbOfFEjKS/NlcY2W+mr9+wasDkdP
OcEnYqJVpQ4wy726xBXLTAk3mKVMz2vmk4qU0sCSR5apL757WnDOrMsHdi5As84L
/nc6tZX4/8yPne4PWRNK/bUQQVI7/cFdsiDUd6wrLvlAO19RQ6NnubbpG9aEPzgz
xvLxZL0HifwmW0PqKDMqsf2fK9r4xWBwE6FAqKFSU5AD9rwi5tC7pf8/UCiCYbxW
wx45UOEuElTBqy81hypBQoXjRQ7zi4bLNe6cjqL9Vd8nqPxZV/xrV/vzakKfh5V/
sAGDIWrSvnnOpttxZo9HG3pnhcluU4b2Kt5okEoTMuUl1XIo/C/igHN5sl8qAEpy
HaQqCUR8mVOrWs+Ab8TdGVEr+934SV129MxuqhwSqTUKOAPfp9zhSa58mCU5vkYc
fJL/Ydpij6mP+8bVG59RhQYs63muwTW1T/WH2B+02xuLpXIR5Nm9/wrJg/TLAiag
xkIV6v6UZBl9Ye4GnC36N7JDq5sMIx6GeTerkX2MaYof97DOBLGjA2Bo0taAkH8Z
Qz1M10DUV7+ltD5Sh9nWkGBhtvoXuH7LrXMlCurpWyZj1HBVL4iXnQk5F01i5YGn
IyG18CFEbcqMW0kxf/KooTAkYSVVZWqDRlLvYa+I3KqvCE2w5t7HkKmlsRR1VRYY
R6eLyum+AJk3HEQXl5WB9H6yfvBFxRivHUPnSuOenqvyBpuV0yOt2TDAO5l+F/76
4qAZVXszKTv9R570XShy2Yt/d+d2vE0czVjsAvS+RAu0ilMMUVM7Cyx4Tls7yoNk
CqAp27nXhXT4Ccqm75IdQyRxH7OCdkYlFXmcXmzMJV4w+f00aunykXc/BWCyFkTk
X9SV/nMiTW5oPk/iWB6+KSFoWE8KjW4BDzo/G4iqDt07qo0zC0xdBRNBx4HyJvm+
u46BGr+uF8zkLVjqLGJrOETOtFM9qLv5VY5mDKoiXA7dCB2tNuIYlNE3XWz1Q0Gy
DMDo4q+40ti82khmgLK6LzLy8kbmbgCrY910PYCE3/O1eyRIKxCEz3mlnmZNh20/
ctBMw2sNiAutcs+EBIcc5d34BEva3gXVoStaYyL7PD0Pc+4PZTikwHAkv25G+cbf
ArQS+RzX7KaZXfih37eIeBWOP3CbyZNTCCst4Pn5tSn6B3rqtaJBxQSuqcOluuQA
glJjcGWMtnWykOKGImIL4LHAI0SCczIn6b3RfRFCe6XR4NIc3sM3I2qEwEVFXTJO
sa2w8GQDCi5ft/8T+5xuswE4mMdMdNDtZ6+3c7QpvmdZ0wDgSe5XT4FATNcJVM77
Me9Pp1tx6bxk3l1xDjvTaI6gnNzjT5BAx21wU2vmG3M7NiRHX1/D4lbzAS5grzoG
vm7eFHPBUYAe8Ofky3KGSMN/oCkl34AStX1oC8USZJVZn8rHZdWMJBeNflX23knI
faobQTt5jO5qwtEx1zn1Kf7IcMhBRJGyCKhll8PtugU6P4bfHw1DAxHc7n8Gd6zz
55/qyeY8Y1/jsIWq9YfOGBa0Uptn9n4VjtmRNnRA8sw3Ms+j6QJWiCTdt1XgwNmA
84URgRDad2NwmI0MjR0DIR84v3sif4w0ukvOiuSX937FYqwQ9gebFTAgmA6w3bXp
h80TFJJN0UKxAZiw5EKOP1Rv/4rOlm3qmsYz5jigSbttiHrfc/L+lcVV/SWWLT3P
gssX13x0drS/Nf+8X+qh0ukum+JTNlJ8eP+IkUj1SiB0dorS+w8oSE4UtPHSHH/0
EgXdxsF9labYSsKGx0D2GGWqmZTsD/L4upsQrE0OcdYKk6sb2922UOfda7aO6YTD
Qo6XgUvZbgUpNdCkiXodQ6dG9IXzIC7/HQOd0PDg3OVo5FrXidzDzjb3fVrojWLY
eRDu98kzlwb1btBXwJUrfnUDly6nh7/czUKtV/sLV5rdFxDwgaTWkiKwsrD6Rz40
EeJaSd0gldCBf6DYqkiNVEArVuegsfjUuW5ER4Q87ADQmhGgfbt2VN53Z5cKiXwB
PGggo0yw/ehhoxFhawvLHGyzcHnEMw3UVmneJw/nr6laqCjTxT6SRLPqfksyzeOp
kFac8WhbfmSSX5JJeDxxnt2sZg+TCPf073WFqYQLgzwVrabobELMjdH7ezsSx63h
qBAY/qFTfUnfShAyMMwitdF7Faotflxnk7wn0W4n9UbucpjShPHADp40pe7RhqBL
20FxnUrXaLN79vkiX8YPF9YCQ4FEpslkEDHAHaZT9Yu80uAGdtsJ51XHVPEpiv4A
7gXkBtsd4ZGLRbVcvZIcwuieWhiB5exvDPX1P84VfUlwgmYkpyiflj/jnkSfb0iV
7FWC1sJwFOZkoKDo4piYu3Vx71llgHKvkqX/pO3dQ7Lt9/14yPMLILF9wJ8Juptm
RwO2IGYw21FossbEFbOpYXrDk+GQgBvsAE+JfOjjFFQA73OKkwkpipx+vNvQdUub
HZK4JI74w4Z/IUTvfSGWCcdbZrHmJioNs/plLXg1+c89mQ21CT3Su3Is6MCKx4Wd
cNnM8C064kL9ocyUAFPA72O/UG5a2fFTOQ16mWjQznb8ltxtm/lineLuquJODUFZ
VNuK0xUnixpLogde68L6Sb/pdGRLIwFxhYJ26sSMhWtdkjgee44RsknjT29wD6pi
8BAuOFxyCmi9Twp6+QoAJjuiqDLf3ZWWDwEj5GdQ2nJXIDbFtAa0NkilcsLSLdti
o6Wc4ztWAVGsSLxUKq0gUZ6eLMKPP8kmKXIHij84mihcVaPe3S2JB3yL1g4uxUzX
KXIbUTLCsZ5TfSKBT4xfW1XN6QQmoAXfBvUmFkfMpwEkrNa0z19nnMBwja5HdRvL
g63QmnjHuaJWrqcIocDdteNdRF467J4ejVBXoLCG7wqPsDpB+wEhaGEalBk13EpP
2O9UTHX/Hgn29pBGVWicmXCRQynn/di8y0V4YOcRiP6LCZGYwGuU/0Sq5JZz0o0f
7rYEP8gxHfS1Gl1nWcg6KidImb0VB3FMy/bKln3WBLgF3niFWNfqNUZ2FUkA23JK
f60OgownlwOMtCf769lLMdFBRPGHook/gwLbQjd0XirVXyDmZzQyUYxe/Dif1Clv
OXFvXWPNC+uhzlGiWte2wcoc1ZbgbVidUr3eE7IjpZhpPninwRsiaXJqEG/VDpnv
9zuemlif+duhMe01b4FTS+j0DzPDPZ87LKT1q0Of2gefxIeL1a0y4JhqTFOggyLd
Eps/se3Hz612hIgNUm0SMXy5FakIrs4Kwr1i9L42B+Aiz0RzGOaV/almM06s2+MT
SaKtKqcPyQXq2WkmOvxVPlnGrFMbDuSLHfHDlcbwSC25HEZVaLCXJEXqAzO/SqAb
a+DjNqf3fzefuxkapBj8KlE3wO+/i34sOa/+2xyZnolA9utKn6qZY0lyUcoSfk4Z
471uWjTn76vpf9VWmnsawG3YyoHCrfw/Tc4WV55bI6aoyebEBb4w5RZeMfxItGZ7
is64BS7ku1NM7lubp6G3UMJ2OmxNDM71hUIDSpOpsgUDDnSSs3k8S8hymxeWKzmn
gBNsNPk56AIzifvkDYF4MZOP0rovL9tCFaaUvMrDtl3gjoQbKbgBJNG0zKe4nZ/B
wsolglVnZ8xRRW6rBQcSsj3s0JVfQCG3169MNjUSpYdat9KswmbPH2BET7Oq1noO
h6gGesfBFHoApMZi3X8bo+pw9fAIR9pT0UUP5gNB7Kf/MkvUM38SKBqkXaysnJWq
Kgcy2lrj+vAcgcLEVv8dxe/DtDvCOC/O7L8Uwu33HZ5Vb452hfV6AAJ1m0Gb1gTI
eao04s8G6QR3wl1k1lzQ3nYVFYHyuaenCiWR5mO8kUC7XPyvDRiWz+3NAUZYo7y1
kWTfANOFtvpZpqk+NOofBHXtMk/t3CYf+wqgBh+gezFmK+DeXq49QEEERSzki3wP
xapSzBJkxfrz3oWqbBROI40Xs13FUz9UROib6EY8syjmJZco0Dw389AXId3PYH4q
VBeS6ZQmWmNQA6/f48AZxlUTt0IKVBYrD/nUdYUUugb2cUwMm5DFr0x3a9mgTiBa
OtWqWWDw27ZErh6bCNCd9+0rNsm0IiVBhjBYlJ4snaxxYhFthL8Pid0Bh4mp98JH
vge9DAuy3SFsg2BkVaM+3eCjUxiqRLvCoJuoz32jRpyFUQVCXNZx+rPd7fjJ24mE
isrwcV9TN+ZMlO9suX3/F/U+73WGIp0rWpO9z0k8vJcf0RzHlAXetmvS031CSp2c
Ita7qR3I1fDq9esXLp2C56QAnnkC0eYGgAA3iNFh0zfJFRhNajjSh3e67bv+jdFB
+5YfaNwbDxdi7ca+baqth4AMrzkBPZ3NN5YuQAdYt0Hia2rxkSPZt2Pb+VmCVLDA
trhVQ2ucW+Q4HHcsLzRvvhmuDtzNpX96jLQaPnF8Zy3vKNJ+gsYRBlN9iY0eFPwQ
OSfXR0X9hXRIfR2zdJ/ahdbOLNohFKD838yohRtRAzz9JOitMhdsMRSjOqUS1L1n
CXBH66A5GFxumOoF8ZdsfRK8D69X/NzqeUbBL2efT+/SVXrqXUBrzEr5SPgoczqN
2zxOwB4dLb52eB4VJjciOBx8DHzRXuSrrz8EscGp8s5FKRUkEGilx5oiy7THUrGb
dP5uN/itLT/M7AhS+yD6NyAiiiQ+jIb41gAPnEMaZP1J7ACPcx44KxGCzN+sQrke
TIHmw++3vGL6UK9LpZaadpB2Gb8ULvabogCskon0TCWTqi038gw52EN3P1ZJ2Xt6
lKCI70qF2tymBqBr5CwYSVJCo5MzjI06H7oC/5Yv8xraZ3cJjY+g43ZYuKndZb+d
2FKIEBIajRUO7+9xCDhNrQFyW/9acygXfNA3hcVW/cx2OBxHnauw1ZP5BpeGvnNR
0aNZm5dzgG2FLsjguXsG6KV/dgVdj9bKlrrGJMSkPyCpcBn/L7tlx1QV+bJoOt9e
QblGOTuPdWbTjY3zX9uhAAa4ngflDJ7j4mVtGmwh0WYO+wcV/Gz12Zh1jcTKTvy7
sMbpEpbB19aKOYiv5Nzyjgi7XlTYuDRf3TZczZosTKRzo+nq+LL3O22Tzv2V2i6A
GZaQdMmJ+pVRxffSklUn1q9PAfWZgLpadN4dNIQjeeqgdA/Des4Bf7FrZXn9ayE0
rgxf2fsoIwAfhIUdkhPKYiJYXFd3ce9unUDP+WExzwXRlcvxx3iV3lLTTz1VK+ma
AuiVnGVnq3szmvevJplVxk8+kxpZarKIrws0jUmmp+v4PjQK4zpOiUvciEY19zWN
vPdQUjcukxiFJ+GL4wAtzkLtYm4DGN91pp0X2cV/OVMTlso5K4FLtFWDzZeLiRav
MNdza6TTq/p44w57/Qz9KJdEq00jaT7LawQdHB4B07uvJDutSEKlK+3fgylgCTuu
zKVNkfAvcyXmuWZyTV2zDfxInnfOE6SG+cFBDJn4wK09bNgScawqpuyVY16JWddX
nQrLmT2DAqrGEOBJiZfhG0bM2um/5OZTNAy0wt6/pvCmTzvMf9OsQf5N0LytKQZ4
q+Yqut+dDLg3t+S/CYiuOtGNrel/7kDeFrr6l19HT+0uVlL/yeGxD0NYIEGopa5T
dhxr3oiuD2PLInHwe/eMNyiuTJjGCN0gM9Yru+/lno03ST4UccgIH8yxEkLIO0Gh
k5t3YOlT4RL8x4xtQD8ANy85vOC+Cnu7Tcbxpva7ewmBnUfuXWxUvIpAV+7dHa6I
w9vrSlO06q4KYbT8A9ua/xEwaBtAX/bP5pitkQzZ9/hvnFXeLRODN8BgyMyeuw/S
TqKB1i43pmT21W2ntrFpheNVs6mbih9BVHc6b7FNtvk5Z+EAVBZMwJDYS8XWdxFy
R8arl454+3kEIL1fexidEtM23wdRi5KBvnlSUN5T44E6YJ404kvfpqWJ5tN1ck4F
xsJKvtnRNUY3JD4EGodsnpQ9ts8mjOAad0P3YIhTyhTLYSpL6D/abLKjaTW6o0by
fjFILAvPntd1gNWCMtropQKdr92Z74cno0TLqRhSnOmchwvWoRAAswuwRg4iE1JT
LtD2/xssT+7p16Ipq3jqqLYNRfjpdIlT605zC0uLEwea+z6iwX9L0Mk6168zRr2v
x4HMB+uVlh6HCIGE9f5mihQjQplyna7xFtmB7/b3+aC/m5MWSAAUZTPoFZKFubIZ
IVi+9YmkWGfSTPGPB9XfkrV3yhepzo3bVVn6OH7SbWQUEMOG39FXfFX0YoiaR8JF
LnVwhbibe8SYK8CyQt/Vu5rz1sX7Hf5YVGZOQGjXsOfS7+NIG3aJ1mVX29KsIP+X
Z1GS4IIIC5tLuU4N17Dw8/Ohre/HHNs7BWHsLeaHTkbrZ6hjCEZceL87rGjKT8IV
Xui1ZV9dUJH+IvGEh5EMTwU1u80Ijxswj/Oea0sNoygrwGvuAgMdpv3bFZnzYNAR
YqHt+OeCW5s9K4GF0YrJj9uIWnqNLOOvIrbunqqT4eYFDO029+Ry4N6Nbeh9WlkW
BJNF0vCa8AfeOHAaa3WTOXNYTQrbXR81N8hRppnyq238AambQRQMjoVZxOypS3O8
Su8kDbcbc5mFsfgDtlJ0Jj+9EaA3t+DkS5Lz8nzIU4fIMv6NU6+5DsDXOyXQxj9p
sV9SMKfEbtKt/cZDQegDfl6EouW7KO3d0pvSWr9cj2KPMYl05VrJid8NEw+z6vR/
gZV5PgJuJ/dpwqWEyhpkxw5eggtUfTfrvOOmTKqJk+1/yH3+Ih+zUIDKonmSmYpA
JoKGUhElTk52JCuKHMOW4MZesmeMcRE2AGmm9QRygxhsGsG0v0WBiLr8Ce5SrUWn
MgoRj0KO4nP2uVDsCI/haWfGZbnRQizAWcyCRHFFVcIXN1rhCSCgjoKWLnD1Gyh3
CDaYX4H8qNFIqqga+gOnsz9WkvmMyhWgQbdq4Smtq7efcynnwi4XzPaSXMowZbVC
ge8OX9L49QLseqf9N2ZISnjnYWP7FKKFN9VsuBv/M52xAqK5WSjIA9z+JtKp7fZg
aBfUJIMVB+Uu9sYYtHZjkr/WnBZHIRN61lItHkSb2A1ldMJOwFrSHFlNOMqWpnwY
A/LusfyRZwDLFDJaz8/Z5WdiuM6+45zgl303fPGXmRYVVP/xm0ZhYjbmRhQpdX3k
dQ2060j8boLVQVh+lvZFD+fUlFzSn/nv7LVp+WWwcq5PMMyZWUlPWSmdKHBtV2RB
Dankile706ehuLvbsNqyLBm8kq1yrxPZbenhiiSKQ5nq2iXv2S2Rm8gAu2gJUSWM
nPidOE2Qk6TNgfRmJdBJkmOxVga81C1dp+JtghyMRiU0Kevty9n9Ls3+CkrQDhd7
7nGK284Po0Yc2CXonvqbKq2wneMA2E+LFxmG/7ok5UC7iR+cgAt0bbI04Fytgzra
XQiPiKvze5FJE8tNMcAGgNHCnrYQWsBLtcWEiAxJdxFIn/SbchPSOx2CHSMgl0Jo
qP2ro0pynZuT9lQAM92D8OwemUIEyk3eU9ZE+vxjuVCzQz1vHhzNK449FhqfAbBu
LLgPa57r5XjKZp+xv/QyT+SDA+MmRimPmyNfk8G1UyIbj133dtmZ7GbwMBO/l5ac
lG9ltWpHIDwzU6mWOc4WN+0/wUiF9GJ7MOJqDgnUTvWVrahIzneDplVLBxrhUUhS
q3REEnhQ3H9vtZPV0uFMt9wo/dZYry4tFDNpVuZ0CUMOjjRTbIKuoZSgeJwSu9fo
nFUukyQSGG61vgy7WmmoUwqIPBOSTDSteYvA34lun50KcLrbCLoWkGSxjRo+0G2x
OG4vwzs++uT04ww27MbP0bN1dioe7qupCATRlGVQayEh162dEnycXiXhhXtokjT3
BPufKYok2uW1HX/HoDm9N5LFxZ4VDgMFfck4pBd2B546jzsPTSTs0o56mJ+k/0py
iXoHjAmKJvY+r+V+nTH0Zfa9uVlDKnZeVk5assS8aFVygBSyPYGC5HWP9xYod/L4
cWf2YoZQEX6AfABH+blNSM3EszMw14ivBHJHh3X/rtjfmEIxgLBcA9+hQH0GEfgR
j2Sl853WMLIVMZiznzr236VvpioLNR9QuWMd/so9yJj5lEpmXymNNlQvx8XIkfyr
OYZV1NZNeeMV+O2i1+gP3qQPG/ozdJM8iA3dev5Tb8ehmcBRN+v7eJ1eWpSrpZXC
GTFnWwTNhiGk1iRZGqZfgmEachOIq4PIpz9VPaJrgX2oJGbDPCMj5KKhAZcs4Xs+
XHUvLAoeDmPeU0mIyGKpG/BVPmymTGB1N42mcB898LbcK72aqatX+Z3dL+FY0k0h
TqJHvbYYmhW4FMBp/ZLcgIbZ42z9fLru7oLXIT8V2a2EnZlulxZATs6CIKbpIkpg
nl9KCxG28yyRPVAMDj7m7TWt7l+byIaUe2S5Yip05eXZVo1PL5M726QeuegMXdtw
U5MBZJvyCe3GfW5cJCgCz8qByzr1H9QemBN0bNiiLs8/8JfYoPfvX5Ola+l9yizz
ga/uEAOUkZg1x39I4OunaThJQ8WGGyLrms+Ggd5LHtYTzYXo8l2rY+1V0E1dicvd
AWshKwahI9TNIv+9R8c2hgGeUY3ZpV+pmdYw/1A1rHM+yVz3g6SVKEUPhpACn0l/
XIUPbjRpD6aKRIi7o4rJRaTQBve7qLub7wgiqXMqeecqGzWiz1g0ZIidh3vO3blI
gaABMlHC2VUDrDkQi4hJm6RwXl5zQ3yxD92s5+Y7Z6eXKSOJWYiPkS21AnK9+WCa
QJVYjJaaduMX0TIKrTZ9ltDukbQQGIx7IE5Rrt3kzufGXWh5zMnN0SBePrI5rjEq
9VfrBgabcVvWEcQtE+P4wSTlkuYZR20pXj8QI05QSmXDmrVtweeuDukEUQWr/F1K
VuBfUw/Yel361Q2f0k5OFFRLmOueQ4A6Rs987O4+3tXupjlWqkb8D5C21X7na0at
lZUni04FDHVFMXkcRDJVG1dQrBi7vWe5o1oDeU/BvKOR1qGeA5Z1IeNESPPbe7Qd
FlocrDe/tTNCYPRxS488v83UOEELo0UA8vxi/hOE32n6ojJphD4R+e+sz97aQ5DW
b/EDvlvkVa3dTjNY6kMYzO2XA0cM0DSJDsZmqbn0PaDPBAoFRStWeeX+9x0YUVZY
c7UatLQ0Sn7UatpCNB+wj3GWusIv48Ev4CMsroPn5/ZeZEABYr/CiKTSFZL01K/W
zpSRZmOUI/qZTtzcK7NCl5Pb6L+LlFwQ+fBalCEEDhhORXYDE5tI33K1oPuU1L4f
v1uVZ0UH2+2A77KHi28dw9gA2ROOH4cI9IqIhu5e1bKtwPAOYzTMJaKXeSNQ82qU
O3/sTZtUdrT1FCv4R1PESTMvJjcS8T8XGtMUAngT3rSRZXBBuJa0vJwRp5qLh2Tq
ecYv8ObfQARHEQYbdFJn5hD7GQG+MsnU5ateRP64nCgaswEZWRX1Xwc+U9tER4Bx
CYBtYDdoSQeQdyM1+kZSufjWVI1Aqz3BD9z9p/gh9PmQzrSGkuXV/SvLhfBWJhs9
yA1gTYyoDSjP17sd4Fkb9KQzyMssaUsu6zwFvLxd4LhY2HMUqmufqq4/9hopIQpy
nSKMcPsXr6ANvOKqMU1flfYia1aiey4RBk1xmSfYeOLaLRfnJPcuJNffGw1LJzzW
pzPg+e2yQSw0VDvYTtebkveBFoKy1pkrOi9V/LDLkuyR+/+AtzYKIfAel0uvXOEf
nuDvV7jAm4HG90JdllQ2Z/IwszBSctYi3AbEHTPmPcJjYzJDO1uRNilw8jzd7XuL
cwLHG93WLx+F5FlK/iXxjWZHKRUyFnsqyAEHSbKWK9LCN/iI1/XUaEIN9PqcchH0
uL54MM5oc6d7d8kN9eYELbgcqJ8xMIsFAg210vCzd8wG+lhVbjw0f0EteARv/SV+
wJy0xDzCtEb+XXjghVMNdd/msbwsXgH/kYtVemKxwyAxEUEfTf9r++UmfDhWOI8L
f3FKRgvK8YNygydvrS+Pdy+d2AYVrk/n+6FOEp4Bq/aH25vNyQ27x8YGI6/Fq985
FIWdiVQZ3IN6MFbPOfBz2ODxZ18aJL+ZpPlWqptDMklVXvHaqnN3Tr2uB9KHZMeo
kPt3YSW5pEaGp1ywpivofmAYxzkJURjM44RMoKWQMii26pd+uFbOQXvw5oaLvnuY
XnnFJ5yyX1Gv3q+FnU+bDQZpwzV/pmI84/cL9MTIwHvChQtfoRACmJoZaqtiLEDZ
LcisZwdI72Z61fJ0PJ7IWQucvTckXu46tAtqWgbSe2dcM/DM9IKQeq0AJDbGFux3
ZLMDJgScMgr+G04rf/CrOwY+ow/Mo4E4UglZF6ztV95td5dAOPaGfxZPGEmtKBQp
8QtxftxZOuCF/3UELeyS8HdK5WgGt2iV8R/crDXIev7q3xV2gWE45RN3KQDeeC2m
YtiVpcwa3mlHtmqKdw2bef6eS+pwGrSUSjgt2K5UfI+E+Qv/MwZvacZaoQs+4/bD
wwrvxlV3eTn1O06zpPcbTV3QS1oEQq9mpQVtMiMNxNOkWJn5rH2skjIeTBcHvd1w
hIsAClfRRcBaqYuri+KpXOWPcbeqH8xcTlGIoro0+MtDOgh6ePWPAWN59kfFleAC
dJvFJ2tqFNG/aoe6XKY2Fy2yCFsSYZbp0Rq/Zs1h4advwx1k1oYuxCLHgoo/9M+f
uxhSadKr77gjX94xlLlmO5SJLbiTOXU/Px17q5IEp7RshQ9IAlJfQO3P4yuXfv29
6sn9nW7+ehVrSeisyg/GQ/+TeTfAP/j9qRgqlJbrnJ8ZwSlVXKwcmMiAZcEsAucU
X11i5STUKdN9GGhgjt5mxevDAZDXoeSWI1FtH//9loxUVV7etVFyv3092cBkIjI4
SqEX2NdZk87YD6VhUVUKxg+8CxhwbT/jTF3o6p2CxGWcTkK/G2KKUX4aPtSS/q72
vFH6PXRxSZ1VoSAN88qw1OKQy+i4aJj9YP46hDsGnsFYrUcLGs9kSHqS3m+kdLN2
XWkpgBDcuGutwcFyrlMActBK8muwhtsyv/r6mzx+R6u4Mr3zfBYbckohcxHJ30ci
P0ntJHvNI/zVxsx9xPAsrdb/pqIhro1MVI+Swr9Oe0nCk7I/trBCDsDFhZdMqh+j
uKU2oXCgrjqluDkW4s+nnpPtLUQazdbEYN+rj64CbjTWk3x6NxT3NX2JWs6nB5oA
Nw5em7vgZkLAMP+mgVUP49gHXj2RkPnrV2lkPdF7gagNtlhFrBiCBPLarE58gl5O
bthAlliEMyf58qBFpT/BoawWt1iWHYAhq9LadJo9234dLbCWOgLfnZUxyfQYa3vn
Fz7Uwqv9XHSSBPOpnrEk8guhfq6LAbPMOL4EaZjbY0bM3rJEVYEU1Jki8dOnWn7N
rZI3edvxoeVOjWZTZjkjGJ9NircQhWdnsao8oYXDGBpEEVj/srLr3lglvvo+JTR0
GbnhB2YEYuW4XKxgZO4PTBFsCRLqAglFqqat+4r8qA+deujmVBODm2Sybnk4+Af4
VxmnGgYE0A+v7JmtkWRv/muQ52UFf0uAOXqkA7aDjC0eUsfrSeq8j26sxvsvAduP
B6LEPtXy+PyKQwAmbb2UTn4QF/8heaQmNLLv3ulI8uTON+ChiaOq+FEYI6r6h9TD
19HwMXx2X12DoYsnoN2B8ZF8xiZY+Uw0vsp8ySXlOfWjydac0DTkW1aK3unyqwb8
5sp2CKf7Qn1ct4rQkchcwTux9NdCUfRfDypzAP9QWuNd3ONc8UybDefIR/qxyKfH
xCkZ63lu3AU7PV4QiLOlqk062CWI/JeoJuJMZ0UU72BMth4k+ZzCQm7yxH65ShTX
ctKfsd0u9ZpJe9kFUImlfPxkosg9DeYJ+s8JGEIJ+HP99Gi9MEMD4V7rzXNbX2ai
KmqzEoMIolDs/ji2+DvxbofiDGnpzt2P40dp5aFjfkPzu09KpBdix/Vi1/SJPObD
a78tyxw49Qf0Sfn5GN96CbEbC0VTqn7QSGqjPONuIa5/vvV6panPbS2hT7KgZ/8u
VQdSsaPlKoDq0flXNChxPkH1E8HuSj5SQh5+MAa2fED0ZF7foernIUQv3x6lUIuT
AYAJ/6ZqUdfZGaoOIh+S6xlcP+dkGykOXKpxkJYPHnsG0gNKwd7ZSDfUaHPxAxn6
3bQUh0MYzdvrr1I1ENQLh36A52gaBjJ/dPcm5bUwWzbmAXR4CDBlLq9VF3hmjJGj
DwIVWRSbJrXcYUCXK053BXuggQoDG6rFFULc2CYbvhi1Ilro5nmW4HuC6nU0G4+i
qxDxqemgUu0jwMsDs9rX4Mw+LMHlkQ2Zwjy3wFoXeRnoS+jhsevgnxly1dAt5c6X
YBznlNUKILiRvM07+rItd26f9Q7SaJcK6c1iRdQpTzvKBE+HDUruuMUANpa/K8nz
CrwpRdbRXuAIfyYRllM+LUYFTzV4VumNzfZZRO7G3L4KrRO9p1l9eQvCi8t1cuBD
ljDetRBOsEq+obmnxRmLyZloJF9VCIVS9XcbMUsNIuAeBsTNpQOrQQByOsni0y9O
T+3QO3xG8o8xYFyUN2j+6JUpPkezDso5xIAFBFgNasjKsrJ2dYoTtoD5JLTAEs14
1b87VxwRyeexwzJZbz2aYBtLUo8T6wl1w3erNcmdjxQ1noqMw6aj81gHqwp7hONB
XTv7VMb9+zrFDA/RP2OVV9Ja+c25rOet+xq5NiW/Z5cClpEpgChD9TvoCMB0QoJH
K/pZfe8uXwEG/Olb4E+rBjwTsVnELsdnAx++tQGPQ0dhNBTgqDasUhwfwxlZ+oXS
KO+kPZA/gYKHBAkGLgjGNyXbnxgDi+QgXRhsln/QPkcCIwC9vbWeom26axuub4Ut
rttoCX6yeY32vTIkM98MO9zgEYQbscVvHebbhh1h7gsiUf8jLdedqi2fRKba2pnD
gziKdPKxHPKAyjWggxzYCfc5FUKfGsNlwIBhToPqwy5+LMSg5Aupe+XnVcZlyIFr
6AdoFILj0yClapF99Kv6S1bSu9G4c9pOKN674LfVaaqhvoN4yLQ0w7uWh1WNbFUS
Zzfo74Qli2o1eVFgTVxV50YG4TlH/8OSwKMRHktgoWGgE0+pf1XcvLe4gkpAKTfw
B+C9gqVVJ/TkTh0ygVXNUBJZDo+YkKVfvrv2/u2uRZuz68xJtL0KrOTX15aNp6CR
iC/ZS7uYobLLZBh7aAce+F7hjpbiNLqF/KI1ABi9J2/qzPqizmVsT1aTXq+kaYzq
BKsnAbC4Kd5t8fn0ci3SaiOPfPSkDzNwFscT7Bk4+fBmuABIyrEwFbI6WrkjQuNz
38Xq54oiyZqQUbHKK5GvSvK4yxfyCQd/c+WLcwdyTrxZ6cS0jPGPnldOlIFUZX9R
RxvRhdGvJ8Tl6LAP7cuilfYreMkYbEs1Y5OE3LHXKCZBEPBndD2npkKgyS7ihlkg
CeTUDmMjHNwArNy62IL8fjR6b2gFdsyjWOfMSIHHMDlIAdaIwRaa5bj2dJTKrNGL
MPKuIr6dZC1cK3hIel6SliogHyiR1WTfN446xzTGHJ2uftAYCkZPLqOP7+6nBjyM
FT7YAqeqWS0K/j3N8XOOksZP2nl3vL4gwBEM5/9bsNUo2da1pBHjH417h4YJYaQD
tA5xxmDxSz5/7soMKdaflSFvCfBe+FUPjO1arjDXDW3bcQd6mqc9GjcnK6uv7dYn
g19mhmMOk61jL3U0I8XS6tY5vAGiIljKCji+Ruic46WpuxLqvsY5EZgTaKSpl3JP
ewxV2sukJYjHBcA2/R/g4A/Vz/CLjnCAo7bblgsyLkYnw23miXDZWk65OuMURm8z
Z0XUpDJ13pKw5CyHVLwf1iUEovmQAx/aB8Hv/BkeO+lVV/FqhIWIjWveKEM1/511
MfPDkRUKi+kAGO/ff8s/tWiG6JLJA7OzR+u1C9t9I+Zwm/91iqOeOTXsw5DJ8IHP
cL1SmYmpUHVPs+uFFx0hAcYODXfMpkwJWPcFWhMNrzK7d7FFX3KrZdQqR9yCwpYR
QZm57A9Gj1CdhBJ7LgNvbZV9Z6kfBF18nBvStpH8Odjz1JLnep1dqJU1n1MauM9F
by4u0eH0tLerjuRVcKfG+j4yJu8A4wEjI4PK4TAIr6IZiFjHMV4/mMMSjlhLJR6k
rcAvSuC83bsCh0qz98iZD+12BN4nvM4Mdsg0ykX9bZfjeAG7IQhmccC0AeaFomJ2
hlMf9+hKWXz0npWUzgy/84tl0RVJQJCmKR03wc9p3Lg0IJBcqIhIdoILFhRzXj/T
FamI4EqLfYyQAVHLpqkFjTGajIzQo+O496XnA2J+VP25f3BUVmMOJkXz8nYU4CJ5
93KglL0zGXsGwIfl9ksMGG9oB49Wm0vdPtp9B6RscOoCUdnhJZOwHMVAB18PTcPm
2Hj/8MvpW5Xmdu19/0CER96t5YH83DqHs37Iw/BVY2Iufo4O4jnkOvJpngKC9AMy
znMX2YCBVOPJPa/1JzFJCYk597IzG6J7WiQydAp1lEG1lZCUeJ0MwmaKbxBBBHZO
6cMDc3k5KogUPTDpYKzokJNbuIdAKjQFSzYtZYYsLcIwYAGYI07QmZ49jsVDKW9j
L4sMYT/PfPs+QQGKVQIJX/kgUYDQ81O+Yfarki4ApuOyWYJTMkesUdENtApGa89l
UXgWb40odi2TUOIkZYltsrgesD+0GeruToLM/Tlzti8QjpRQDOMxkQboung+xN/Z
i7XoQ6mUVK6b8P8ygO04Tn4qljhtImQsEucjWkj+PrIPMenpbiQDgcc4dcg0PlQk
vtU0kDBd/DdItfqj50GlRb/Yc2uKyKws3q7u6EYZa/84i4lKP928DzqsAMW3RlOB
fNMnlefDO1H80oDeImrKRaowUlXmdSOj3x7kNbIHuFAl1B6Upx5DVycJrUKyb/du
oCpL3YFcqTKNUOAKPUC04KLgOBxCBSmmS2kkqgfrk92HhAdWyQVvVBTUTwNwY6Dw
bfZ/NNQjdCvsKu8/WpqtIPvB4agsFKhO1cTjdcMMDVlVdJkq7etSXc31JUliZGYq
V9lRj4tWzlvB0gspyBNR9YNCEZo2c+xGoUx61UUzsI3fSEHxRp4x/J5DJfvFh9Nz
KE4bciTTN8IUpjcbP4cQBHOig+h4cqCqKZPmuPiMzTja16AFfqpm2ljcpu54NJEt
Ny15t0w8PNDWkExOg6RSgoNSiU4MKBbrIpLvCyDp2G+sCfj1AjKcEq2zQE9/cL2E
6XOZODGX2Shq1vcMbmItwX9SHskP93lnHwJGRIE4oMAjkP0YJSCav9e4xoWM2p9b
1F6unm1g6LTRNErI8DUWoOpuAQs36XjpasKJBLXs2Iu98BnCkoQ/v+uqS/eW8owr
PtIpYAqm6KB03ohA6365uoWylo7TyDqF9BEuKZrkDl4SKeetSkbwiWCORTye76k8
82FsFsQ6QcNH9b2kz+jYlx/Lomy41Wjn6cF9VfocQCT6va3NuFxQoqwFFGTL01sN
r4mksB34wZWCuveXSRJiHGcxUXyuwpPXsaFkuCFc2lwkeRFezXluwCNhHN8kMdYx
p0RsIlUF2j/iBCZUM+DXtb045M/T85PLycLJh6cNiafiEE8I/Nspp7x8PFpsuHpI
whGmRnGeo8ZXTrlAqaY2QJ132/1PKUJrbPq3K0dBFe7ZkkyUFADqOLBQ7E/xMDBF
Db4AtL0u5udNlRblIuYt0Ki1hTRxFUw0RrQi0+r2A1OauFucupGXs/g7iOPnw/cP
SuRixUl44WD0qyPcIb4CYxYjmguos/AUXJ5i8cExhEENmCv7xsd56HrfNtP5TUvK
v0yOCc97BYqzhlyAi3Xq5sJaUACIgtidXs+RzAXKVWAck2yvcrBe+VhN8Adgi3Rr
LjqCaXB0DD4ZFX0eccm4pyiBr2B8UFQwMemK8r/GHGFGMLK7FVmRFEXF60UYp2kh
qakQAPz5VU/e03LU0NKJWRDdL08F435yaOopOcLi5VTE/5Vd+T0VkM/4TwuihWKU
XxCAvYEJh0/o3AhFLx5ZYLjGpAbNqB+YPsvk/OTFXc/b61XwfewNoujrF2sWboqy
wcdIpO7USrGnI4SmF5jtWq52/P6M/4tueYKafG0MRNZj5FnXllWJfbWaOybKQRxO
VtDxYcU97VczSKfSzG55HMfnMihAZuKxr/F9ojxQnRV9uoxvlf+9kdKIQ4TQNrj7
URTz8RJ6qvDgf8x/v4jUjXdUJnp6uW2xmrb4x4vt3ljgmOFWjJSwk0l39yqnP7gs
wuRhzR58dXTi75G7+QCTZC8KZxjvodM6sT2uQEz0u1ILJlDKdalozH5N/ZqELlg1
+x9E0Hf13tiNx0D36PFBSPCj0RN8UyDerI7RcIRvUjXgRr98ZzA4qNv69Kos96SM
qR4X4MhG+jkPvXtCXkZQvVNFPK5MMAgQY0A9FA1El/ETc2rlr951aW9LkUTJD4rE
q7M7A3Djzs3ddDFiHjhd1Bi/QziU1/Pg5kx4Xuit20I9t6a0Z/4CQD0tiVCX2bcw
BbSefLSs9YOBpKA2qS21UXjtQdH9i2LS6asjYzcWN5pIz2rLfnlvuT9AHZCZ6XVY
FElhQD0DxoEK2NhLCKAK35vfLoZG1unGBwJDcgTM91PxEexmeFqOZVr/PPPumb3y
wXWAXh6hbDlt5k+uNyWbD1tb2J5SIFonUevFprXc3mwlo637qP9umQtJUHZdDBB8
o7SreYRHdVnzqprEMosFuDtgaTQicNI5hvuKSA2gRRaKqGjU/fFDVytIDMLlcry5
rqhH45NVa9shqoKTzt6TuDulsfyplPsr1f6XrAD++6EaaUno72TRIDig4qX/zE+0
B59/6FK+zQ8uGDDSXZEce9aLAJn9rIBp/O9pSiZpULwgp12oE+BAXh7Gva5LRYLG
4SdLXEcVZ2oGe6cW/uwU5fH+OCK7pCb3GcUa+f0cB72vr1u/VkcXySBr5xJV+UDs
gifySNQgHbcd2QwCn0u7M8hwxxpNIbKn05hC0RXG/DHxU9B1APv5H3IpPccwgVlS
kFHrdY/JYgRGE7/9qk/L8Fy3DYg8KO07cTy2m82YXpNHznfbsN/0v01lKRueqZL+
fa8YOUGjiVNUe8oO8lRoNEGsKmQduueQjTGMABJ20mkl7+YlYOuUOagYSz4zSv5f
54GaaP6cewWbMkM/I4efkhjjbmXmEsPCY/RBdqJ6L8S9zg6dRRuA37UnHPuWizsO
uvLLqK74U1gDVAsnVdTgL/EH7bnmIscGbmFXk7MnGBsAFKBpNTyAcdZQWmmuaRD4
iEb0gWB8mS5SVCkBy/5HGH3/J5wTKvh4AMTK6EFg6DSvy+an4qk0tdKOdgC3sZ7x
Kq9pkwoRBB7cSvbGUNr4OCFipST6Dx+jIJO3xRQpaKtwZ09a4E6jJMGnAdv9h1IK
vI+uMgtaRtMwQugVG738fKkqr2eyb6r++k0dFKlneaVEqqb+fdvjzsk7eb1WFZEF
TZsOW1pbK2cRuMM8Wv+iD2UAwTN7c9q8tf9aNWRy+br185Q1SopNIkFYIe+5rJiK
XY9AW/Maw5PGRu+CdJZGIjo6tyX7VJi35D2iCvUQhVN4AJU6XIf2gHBwHXER45sm
1cyoKZAzz3UITSd5Fi0FXRQ3tchPkY8RSFC35csNSSMOY7GBr6w4lJ2ujZWA71qg
pws7HxOH67hZsKIDJtJPeCbXS0RZPc4AT85my430DT56JAf5DKMdFnRtOE2/jrts
dfkqGw5Fu822CaLQGk52CcytjQRojpSHUUNc1I0nfJGAVT2JwYY7Hzm8moYyDAo3
Q5xPVh1udZV8PzrMdOOHchw1UrjEeShloBDKD2udrkgHsznRy2T9VTDO1F4/WGpo
E+xEp04Pu3yrbF+KQWaZMaKMmyZmCE8cEpEbdcYMAFhTlsTNi9rTBI2jyqLt3JNA
16wWaotx0MR8YCVi7LNbTpNS98w2844vyZNTCGdnU6xJDcGpLuuKWrk0goNy3+gF
6pZO/LQ95d6Kmok2P9iRunhFL2TIS9fvL/U9s0/H2aA4bBfuRY9aTydIhwgMLrFU
BvKe3KGMjdfRIym/hUp/fvw/W9svbGT5J9aVPiAbaj3BBLkvzh/3Ggt8seWGi+KD
Klesgh1rjcGaLhYN1pFZUMzRbre3BpRp0IRbP8sKX/WHRrA5j/2ekfZ1rUO+dK27
XD1qCK9jiPbDGDVyD6LCDcp5gP3eBbiap/jZN3BDAMsbsdXkV9M3xMTZ9q6U9/tN
+Q0gY+2eqqf9lhzAmND2CjYsj07amsQk+mmFq6Fd0xz+a4fyk8JOjPI8i5DABSLc
qm51K8FQaRQSRay5ZxpwExzen7C7LHI74aEeFq+Ouh8j7U5PRTe0kyJQ5B0Q4uMx
uq2aHo8dUvb1oBRxJnKXLnBxW6JSBZ7qwQ+Gy5kT1i78/ZqlIiVHE4rsspPCMe8k
d4O5IE8GW2+TWsqg+IBbdNV3DhcNgMC2dCd8TbUavPwrFmep2oAPoIhnvmwFD9Gh
2p27vI8YWb6ULCnEk3haAHF5IjKboPlFgvzVpqnAirZJ8UClaSMqXGSwBqUP/rXn
6aIzr5j0HC7pplewOxRkGIRMqzbJAJz0axNRX+wncpSmYKftnMX39AjNbzh7YmKd
1OBxAuOXsgXg6YxzROpylM6OkUSV0WjAyRXRypYnJI1pki+/3Cy4RgmccEtiKMmv
d8olfDyQoaRNa4O0EMFtuRgNfcsHbmEcqdXZfpG0AxT+MtQu1yOWAvWmL7CaSRh6
oiE9Prwf6uMxas8CplChMTShmGhzA74TmcRd/mi3juYpG9aoZaidODzw9iAJ57BZ
uzys9+M12VbmlBPuwoIDRUwbihOPtGbkRIdIdJz4+p46b6oxgbD+pgqMwGrkHscO
ctkWp5oEHot+TQGmScVIKtp/6AhN0i5SwbSqIFs+/pwyNJmUAq+6uCLadxTJe0Lp
3dddEHSy0RDl0+fLUxsd+/aXQ1OiG5cxDm0Bohlp6ar8a1ZVE44F4z1uvnWGXnQ8
JcVudvib/zS/9AD13N94Wqufq2npMOCNK5aH/jEiChDogDd/pUEnrry+S8OZQYtb
3Ycs2kgKSWoZPmNVuwqqdk6YxtYGzCArIcUzTLIWXZUTnllbSXWc2o4nXE0RDKio
CefAZB/yxOEXERLEOeRQKbj95XiyIiZN/2xT1ll+JaGvut+y91xXVeqjJQbBoVVu
AuPhDH+hEfdE56d3rdRSQ4fIlZKJ6qa8nCEEg1Qk8SB3mo//5LBVphtqKEjikxYJ
KdBnT5tQFpYeFtUFAymwUpdXgTDAPVN8wf9nLoEOKlYRz0eiWLHV6n8rimGT7V2B
27pZO5eSJ6DE6Fte5/3vqZR99klehkhibNGFhAI0aTCFurE32zzOBQOyUmDjd/yZ
Ry+a7Q8CA9YmArnNBGYFfS2/XQeJIYG7024Fpw+3L0tMqw/VmkvZdYl0uLkdbwF1
AwsGXHiAhFDoyR0naOac2bBNZa2hXGNVa4tYd9z3RfaNUISebiVJ4XL2wKKIkGRm
5iIUZM9JQ8TRItXKmQHXXwP7upozd/8QQlR2zdmf6iikS0AhDKR4RhqRzAWDersC
TdsuJehqrwO18wkAdAWTT1HC1oGaNhc3cFobegpkZHMgT0vhIGoYDnucyl6yqVo9
kO60t2van44UIPrY7fKCxNmSPKjCsU5hVQJTX4C5aTDb1A6krwD0NLWtaKaHPzlA
O6zZO5kXLrNKLDbabJkmmOZFFO/IQppwJ+J7hohoNu486UyJE6/89sK3wsBjxM3Z
EbOl2SX5CwLZM8iYLSNoHB/tTzyHbP83I3TRMjUQBtu7SNECJkGMGa3fb+UWRvca
j12X5tnj/EJysi8vITVJ08CkWkr/AJx1ggUsCqT7dHtmodIV1FvEXhZReeNOeXU9
b+ezB26duHTYY0/HGlA6IKGIP1U+b+E5fQhMNp+5NPCdBIqXIbzJ6wVCQUyf1UJy
7rDOcSHRpECIaJpY2IVPoQsrWSCbkZSY+67s558nHecbMZ/vGOzs8veGH40uNoEz
OOprdAskyIcE41xAQ09d2a8YL3odj4gUqk5q4cGRSuxy5z4e57W6lKb7KWKZPFSi
H6jLhaZt25FhMDNviPsKMTIlDnGTfD9NcYRvGaUCS1ScBFAuhh23LFchByu0fiz/
QoKzSq6BR6qhW/zIHrRyiTq++hNQwkimInB18ZLXNpVrqu7ZyMuaflxYIFI/yof9
W/zkclzXyYgxtTXnxwip0KvJytZMAoGtvAaNH2pGFyAZXYLEZ8YN4MrnQAzEq55Z
SeisJe7dNLWdNjN61PLj+JI3YyCe+JiSdP5B+B+Q2sLdQhkpFUXydTDRGVHR9jkX
78Fc0V3OxaLBXO7cWLdtX7kee9vFlEMnTF7UA5bpqkH8CqOjGaxEuSrdhOY1FYo6
hv+XbcwQMBKq4YaKg6SSnYEIv6MzAz4tgS5GG45dFut8SKdRjQKKJOE7EwXEnusf
P708GnzOrrqJGU6eKzz/QBSVe+CaaRd8dUhhdadcTpvdVV4LJE6KBjLiWkyFN+Rw
e3SnNTJnP97u3GlmV9WGrI80Kir/yof56NBWvvs5kElJQbmmx+GnXh1HCfAKxVje
ZQLyllkDCfGcuPbihx910Y5Sffu/5kouCG9Hg/k+koDXTBSz9BOMav4scQHiJxH2
zkgD/LJ05+PWA0S1Z0xt/OmyrVcY8CJ8jvpiqJ7BQd6J3deDwnojuqs9z+y3CbEQ
Ajd/7gPWQhx3Uwe4iRZH4dsRJEMtRWscZn6H93l01+j1kJNtylj5d4Ih1oumfqXw
xNDvrpuznVdwnKQ4EKIUliFZ6osLmy2FemfLWb3CtoThb4rqIzzjilgbu97SLyGg
9AB68hT+hYEjMQ3dC0Rmm1uPEECu33pJn050HEdN1B8DhmRljhy0rEiiVvB1T4TT
YuXG4vPKC7pQxcHS285+2sVmahp9m5peg2lCfj+w60nNRVs9zGvHHNXYYkmObRtH
xyPrsVqqPPByCpEJAcX4M0aw4IXLhqcBrE1hCPpIpmdcdwEpcwPRnW3uYcpbnvJL
YAqW1nMH+G20wO2NwRWE3BokyHiFIWA4zZCqe8wO/3eaBXYZEPBhU44cWME2prDQ
MFaKuRK0ZWBTdTjmksBIuQSWlCZw4ZSEAPgTb1TcrsveIY5fUMVDu290mrgPzGKF
XLkmbLi9Im6DECbxqeAFMDZiECF+4YEjQX6l37OY3n7+e1hQkWD8mPdFGWU3vSpG
2OK34FC7Ky8GRr51jspLr9gSDo4QBfsZKzWBdaRtfOlAo53VCRfr7Xv0WIjkvON0
sutspTEm2Gg2Asr8PMnG9rwynkOSp3sq1pNM8uZYFYTstPOVDyfnWDHmmY+tymVf
5M9vPL9byFAsfzfFXfBp5OSWkag6tkGh8AjjTdYpI8uoevTXBhtbaNAJ5Oga0uap
NMnWTjogGlKzU8zo+AbwLHsA6gYtmrxDgtcEwYTV997hTfXMrMIMoDHvaMGxaTNs
ZJlhAuZRcgG8uYb/DmPQGu9c1dip3cC22Tb8KawMQ1TRJuOmWf+eCqeZSPxpE3qs
Al5HmGOLr2No0KrJjEzPzyragIag3qduKHKwpnaLLeKgus/qY7CeTbGlXoxZJEFW
ehv/mAtQKeIzE73DE2vsdZGG/fd0yZIkVLWwv+9AYb/HjWJ84g33i0UFWLtrBTKV
Ve0bemAR3wGhLiLGXTsmEMwDb0I3XFZvRRH3sknUA5SXLOhQ80/Tc1cNQIAJ7OBY
5HDxaF+SMvtRDpmfgrl1slUVCF6/kWFmxu58mT4utLM/D3Zjmo7o7JutVwiAEF/w
IcK8uCISGEau99x44paqqd5l2Otka/Qvt+rhcZebkRYcCzaKdVmJEMKCqUd6X9YP
hHuaxipJl0cawS77DNOIRvaSxLVYSRT6BsTbdqb1IYh2D/0QleR7Ga2RST2G2LQe
ZJSw/70DzTIVPSt3SpeS2+DkqbHcZm5LjND55cUTYCGIp5fPFrJP+tk0pg8pA6Nv
lIO9XO9bGKAl3/macC5tvA7ypHDraf7WmlIOjlAnuyqUR1tmz4+Gp9SGiLlbToFL
jkNHCuayu+NKfBLBojaxNXVcJiRmdQgS7Lo80vwtjy5MOJGzsjz69xXJb2WxGfCM
R3NZzXZrwvkW3Kl+BYatGNexDuiXSZpfTIjOplExcRgT7GJP2b/+zlWrpLcndrAn
1/8WAt0ZPLA69CXS+z3XF5pmDrwmM4pcX/YKjv26cgTl3AJfOq71xY0nwexCiGyW
+TChl9eRzEWY1EGb0AwTHZLxt/0v4dtfq2+JWytq1vtS6aIvNV/rgkZsT6ya/9ro
xHLRYquBD0ezHk1FyfyNL8WvDsBwkAvhX1NxzF/QjvOBbLv52ojtf9DC/hAZWvM4
I9095P+1GlslknEHwdWlZMOGRvCzcdALYRIICWl7NIRiu+fs3E7jllmfI7JZCc7a
PSRWrXD4O+kqtRPHTCmP7hNfrSFR70qI5ewlgYX9W9XOXUJUM1ixvUGyRLyPmN9x
H5WlxPsWsrb06bIPsFKdsktgItOUUj0JhVHZbpfXha6/y9giHcwybmthqbJEu5cQ
ukqQbvxzxkJ9QbVZEmTqja38J73CRd9IkPs01BfUjjNRE3OWalZ6OExYidI/+2Sk
BO/PTWkHpWu77fy9vYzcETzieMnHjuS6NCMPLgrIbMl3AwIE4FNAlwsTyKqCW0mH
IVdLN7gDOCTARVPHiavCU+W66Ph0Ni/foWAW+b+zb+B6qAMlqJEJ9iklbBd6pROI
V+7hS5/Hc2fw5F37tJFAevocov6omE8ax5pYEbJkcD4RX1I1t6LETte9fVUy6RM4
YbIG8ltcZOwr7i37XwpAvjPbXZUD+TZg01gpBSGKfMK6PPJG99bzaRxQD4ZGutg7
r5Y7tSNx9nz8XWiCl7qe6na68YAsmAxH9CcoTIbbfrclMI5l1am738s8GLVNq9ii
MKAswDXTtTgd7pqwZgJa8W+BgPZXW+VHS2jWo5exEM/2uvMJIPwDK0YU2Mdc2LuW
8tSNNU26S2R//331I0iqljAXq5VcGPLFNkbEuXov2+6Qbb8F2X8JDtNEQuqc8b1X
bFZhsnWWfJv1Xy+dMXzHVhjHrpx0bVtNV+zPrJ1Wu/lifRFoiFPdD06TlJFFO2wr
DbDTzrvXc0M5OIPosWb8I2dn3QgD1vRDO+7NZLQJTu8YPdF1RBrUyUCI//n/bM1b
fZdVoFhQsgDzPXIBwGuuoJhU9LlnqYvyTfxlfp+PXY0JXYrad4fICY8u9xEBlsjn
DJoHH3WE2ePRDpv4gzNbgfAiP2XhTn1w4lml6GHvuUz2aEf39eFiM9cB0EBc41dK
p8HfurtVcFJsDJRlwVi9iimDZQGbv2mCyM06NOUqVIB9uboEU+kuvNo3JVVRSky2
nBr0Zfu8iOIWBYie1u6V9isoOSwsTs8P6vLmZM0FLmpIRnB8UItJjr6ncokYpKR3
TzxhdWVZnqdD5i92oHV7NBgmhFLvlFygpr6GigqFwxDRB0YZMSbrGLKLWNTIVfpI
ILF5BPrZBEXtlRmlQPfHXrLXy/UQMoP9MPfh1+5WIw1kPeGMoO7FnfeJHKVXrcld
kp+jL5/PL5kbpa9uk/Jy/S5Md8G41seRItEEMyr43Hj0EobMKjg3ovSIjNSRDwZA
EmEkbpfyOB7wVyI4AXh0QMz9FlbZLTWWqlP5miOx3UfWyUCoadv3k8EGiT+LyRFT
RSRII+hGkbmKGAQFxd9grUss8Yi2zGuT/+43U6XCnYNA57U4lbgNCTDzvYjkwLoM
THyA3J9M3JjdwpUmQS5mrg498hJ7z1NJvQQtn4n6LiKnINl00r3ChkmHEET0HESM
5YRpKDEcZ0CnC9ZZJQdcgN3+vE0dqghj4tpIG6bh7TP22rJ1TPOESYnuE1Co3etW
8SfosRgt36NomPmVGNb0jAC7TCdLW/AR/13eAEt7koV53r/VvvZ/NA4n6Sb4DgnR
5Q0xXZlCg99kYAGuA0hTUmKctvi12p/CJn4O/XTMBCqD8aJWfrCXnydoOKQ8qM3x
F/TZvrQTojmy4i4Xxedotnuw03c3Qursdi9JMf+Kv30vzHmisVBIdwJt3Q+g4P85
P8FytaV08JjdL6PI6BPuh8ggVXhO1aLtXv9jDBfqSKx0a9PC6d4G8POLp5QYWhdy
LIqWrUgWuObZh3S3MgIyTlqLEcV4uWzQ59+HQQzdLZ7UTRdWM5BW0If8vOTuf+hj
rL00BEXZVX4vynAgB4pseowGjHDa4O2yPyFRfGh3IM6kmsZhbGZ/Wf+3Q974/3aF
aTLQFUn4Zuux0a29Ocy4Sajsky0uvpQ8Xs7PFBtd1fms3mwmQXRcR3QklEVJYDfK
UcFPb5eeBliKVfUrRA4Ll8/B0VSM/l8IlxStye4CEdZNbXfPQdjggba27Rw8zL8M
pcR+dsCePfUkCZyJUYO3h41ghnpqNhlyCuhEcKLkQrnrF82fYDiDmo2ll1c5Ibbc
o3SNReMJOHOqvkyQ3hceFx91NBawJ1gN1c6NYKN/hZKPU7uxIbYahdAjv9YmyXff
aJw2cJnD+uiwWeC0AScnDfvQ4E213zhWUDktyCgs2Ko+Kbrj+mYEIaqhgF4AN8si
3KGVTEIZuzLadQEUsrhAnmksRGvvRGmmLHotdz8dRSS3302nGX9FkYYqd1Y8duBE
aqarhcoFk2lcJ1omzHnzvkdGeye+bt5aEs0y3jE2cZYXoDV1aqMoZlL/i8xRjTFS
gYAb9Vl0Ah99QlGFoCOfraGnA4tJUdrnDpTpTPFVCz6rmqXpjSV4ZvHaMFlnEL/r
FD1UHPOGxB2phgaP9O6064CVTZ2mjkfGjz7vI5F4bjQ6xwLL8VCkmnw+5YEpIZIE
rM34/Endyq5Yox5ecDT2YtBMonDOHjUjyl/3DQPNlUfEHx5WXTQs7G3rIukOfLiF
GVxqsLqkRTuG3hzyBbTrQBXbDx0ozGFWnSp1FNVcwkekejq3KbNQGGJDFjh6gNo5
+H3Z7W04tSJKoP+96DX92jc4hUzpoq/v7mMPhaazKP0GRR2pE1DcCYPXUcEpHdXW
7kI0EOF3gI6ZlYNm5JDYV4BWGu02nhANLyVvr1HnZwZo2pXMV1+jFbRGaQK5NlIS
W2o87g2DCMz5DehwKHejSTYyY/MdAe/3jscR+bH9Esgi9gVeCkb0rQFGxbGmI5lm
c9NMPM+f5dgsqJv60WZ6xxIsjMQdE+OKhmCwsZlNI80/tsLE4CdG/blFU6EjNdod
26FfPoxXzbbTe/H1DZ47fZNBFlOKGgC3U6XH+mQAp4MovVkIn9Nk4QfPKztawkP/
GvLGVzNA5ZUUNPuTTVBk9Zg7U0PWY7Uv0U6bKWjOeV+Mt9mDeVx+PbafBBuCLfuB
JpaMJB4FWEVj17Q/vmT+dWKrInNR1yHvXdu8dUth2XELCfgolweTaUgL38SQ8NNa
Q+1m6r2arXa9cdF8p0XPho6uUqxTIrAk7/SE8h0NYFioUPZm0Tf/T/RbnQmVf93W
SazPIaQkjrkOGDc3vYnqANar69P7wmxdzv4w3HkFdvucT/fC9IFw0QeuzqSwvqe1
34Zdl1QvBzNRY4YyPGXvVQyinLTKvpMaGAdrj1ERtzgouaMbWyvPL2MHOsVj6QhS
d2eDAQOfl76etBf8OWlZuBnf0BkP2EMk4dgayvTW42eQnOfGFqfN7ap8OJTwM3Nm
Jrg3Z0AOezGUMB70cudOCaVTTp8PbKUJWtP60SNCC8qjOoOYECdg1kGRk+hsqK5u
CRXSf4CPUH8OMz758jKiLE5Aro4ZmwCcR/j+4mc28AlcKzNuXjG19KspftU8sADK
hKUd0Q/Jd2ufgp9wyZcIh9u7U0wXEds/YrjI278E65AXoptQ1PnkxuefX2hbgQlw
wgFn6v+o7cgTqFjzNrIrYFIFrggci+j/88t8Pie5MfFPqlPvLMPGtUAUWMyITF9q
ucnFzSu2iU57t8iRhpf7qwGVvA34iuP8bzB+eWH85pf1wR/c7Axdms+YLb9Ya3E0
BGZ0DGlLvaOebDDRyt36TAb84i2KSKU+I5fRmSscvMUchegKKk5P5Qxf0gU0FbD6
8vMVlzIgvgK2sjQabAQVWT/dblO+zMR4rGHVlGn2BLv3iVQSNV18DYuHk4C05Xzz
uVBk7IRqK39DaksWUGF4DFkOTepa+9gFX8Uy/3qiQibo4rXot5+iLmZ+p7/D3YG/
CqfEABdVxYhhXEQAiALW9gJCUp7u6u97ovdPkJCNhbgpx4RLC62mZWn299d/U6m6
m++QcLMKqUuE0L4aZk6igUKx38X8YIFMI0EjE3+DNDQVQxkzyuWfMpWrTABV3DKz
PUqgL7nzqCnBDpw7QVahvMqhXr7OT7NgJbMuH8YAhArQlQKG7dhnTty8OwmOoNWb
DR7gNJyyAJkk8JGrVNYK5TindSWF1HjxNoBbPyCZ+52xuO8OcqGdx9OKsKMwF9tu
3N/Ql8vSIAGu6qUpTNKjcDG88HgCYWo8AJOD9jRB5nA4FYEFPb3AWPgtrvOyFPva
Musd6h8MG5i8oHknZ8c6WELMtmrRkD1V7YoHf4DugaMELBtQ6wSaNpAlCCkXnn2Q
1naaQLmRaQPrFGx0MKeRgk1pSyzfZc7+TGCYqQbl7MwkwOs1roa5mMHDyxGI+Fgr
p0DKRM3pg6ERAcPXpNdZYx81H2s717UfCoqb5Uoz8lCjJzB8Esw5QeMxyywP6l2f
1Juizy4UC/ujeCQHo3OPX9gvuk94IXZ2jsoWWw2jA/X83AhgY22zE7C7aGt+c3Kz
Fj+UQw28cRTPv1z0vipfBfmc8i3ZxhWBL0ixxN73nadT14pzwQqxP60yZTjmj1eN
crunPVBUkEENTiwYMZR0IA1s/I6Le1/tOEC6Iau9NXvNUpOdjxxgD1WMxN68+FNo
qmw0vVJv1+XKybPjIL4KzRNU/mPM3CD3On/+qS77Xf87c9udkTZ4OxGs0Gla+Ofn
b/RCbrVbNA/AcEe9rMasSiv1fYo9YY0W7XsZrkF0uLRb91aw0CgSd5plnoLcxgTB
NFy45ZaEDMDXeFcGOPdR246cxzdlt0LLge26AhJ03nszYm5lkz7KKgRCv7A+963z
Boa0CUBx4MBKGRlFLhLqIbYNLd0kFjtzjmMH+VoEXb8IEMoJjzWLZ97uj939RKI5
LA36CPYN/qEO6PbUluHEMWVzgu9bhnkmT46SQQXACvfdy2VR7dtlvBGfDOdujLdo
8BxzSvS8GZJeDR5ggQzBSrXHIbOQ9oEMDLf7ZJhdNwvEErLpQrmcngbP0SCMgUtN
d28dwAxOFNosERrLU3OHjIIgMMhQO09tQgR6mqZxa515Rs3mO9at8UrmFv/lFix9
MrtKKCb8OFI/hheWYYt6GlVtHUoU7MmxggWsnjvV/fxSmeJkBCMBahskSjqGYOVU
6JQ3uKMb0rQLwds2J3EYYCu8m9VpQU56gTE6B5zGP/aCVf5dCDouMqxCKlG792qg
GKSlWFHHNN431RL1Cj/2JJlWFigj7MNtf8Gha0ETSCEZxRzl6svsZWAMBsMyVOmD
qPSjSYx79FOwEQ36SG5p7UpLAXwDk5Fi/8n12mbJevD3oyosiyqDumIVnpsXXbFe
/0xkHTIifsdYQp/K1+9M6DQ90/6bDrzOecTvGqJO2S7KeMgtJImEZK/uSoXtRIub
bPYsP8ph6BAk251LhmS0D/ds8eBixvk/OOvRdgUTK5q43scd1yQhWMxlmc7PoUoT
f8PU2Er2I+j/Uxs51nHKq/IQYry12UX+AN4eNqUhp/Hoq72+etT1pEXuVwSnr9dm
Lk3R8F2xNcKtUVKaPV2pqAB7nbMsIP09TWP3rMTgre4HpAx0ZK5/6+LLgaLXCFyC
DulWEgUwzjNS/SsOx9tzajMgXoXks0GfWX5pZ8jj/5+6YNAes/YyfLMuCcne/b9X
c3sBsiBaElgYbM3S+UVNiJWQMF9NViybyd7AllSLeN45gHA4Jra4Oo+prdtUhlKh
aO7YClKQ9Bl1W3yrhLaZkzbUAz+MGz+o3V58ZzhC0eibKMLOKu5xV0X2zcnMEsZL
QR5zuTp8yokMjAkD9sgwUT3kNhI4oYRloiKvCBzWxcOMbCPY6mHmB4Flm1HAa88H
eXLoOHyekxIMaTaXF9GMWZzoID3yGxPa06Tckx1ouqVjWh5cyJaJcV4H6FphgG2b
rt5AF3Nzwpj0tUYFLl3NwPF3Y1lNigDz1taNrXPnxag18AectlaUJqRVmbX8rO/C
bA1HsqeQyFOE+L7TTi/dDIZHGGjGZKWOH+3fFbmwRmgeIbnIZrXNftYNx5JSQ0B2
ePmkMFggLNw0Ui+wnNL0WbeTe5IdM2q+jEFp6P4kE57Eyhd6wxpAVMWw0xvwiFVQ
CSuOne9UxCTRiVuNIKPE1Cqry4wQUPRs8gjVtWe1ckUaPeJN9qA/qLQ56KZPctiu
8TPHdOrjW31FSb1M415j4PpoEA0KVZ9/+uGxqJJVZCBio8G1C4zxEngrpQdUkIQ0
fT85hREW6AknMp9o4nQDlganRF+tjXo6sHvW/pkb13yv4cYNMFM/l7cABPiZUXeg
GNHEhf05h5pRkVkeTJ0Fjw67BHEb13gPXDh//eU4YW+/GmUbZ6JCing2pQoNW8lu
ZE8khBIxa/cjMKQ7+Wy87uh3H/jsh4Yu3c4mVwlO5sAxUW3nYuR3h4ID3FcN6qLa
Fx8rZAwRV+8K6Ci3XxN7RiQ0NLdkiAGIKUXs6d5RdNgUwbd+0fxFGhtWhRkzheve
mRezxoCWOCZrBYxJee+wXpxUcAiI0bBx6Hz+WsizFQ85u/vzoKdiDYjDqFYbZQTE
BuQ/5Xr0y3frblxG+AIMMl+9q37w3DSGuhdnUy4++AuDXJ1YlnbenVe58wzz6E9k
dmJWFiWZqhttBny/dbqLaWdypdI9VWiARjXb4sYykLqlARRI3FWq7JTdJxC6Vup2
CwKz1xSsDjYBjwpKmNALoWbQCvUgmgw+QyqjEPIvP/y6sjWeObXuthKd0GT7wzQG
6m0vc3TEowKzEJRsfafJKjE2ZKM3Pd/gFHd6e7hAzagFck2lTjy2+j6a4vIYbmRl
9rnAv7m5cEflchXsEHH48ZXpyBFVkg5PUwsunAZ4rWy56eEyxArbXjsdNCJFbvGC
k8YMMWS30m9mRVji4Fr3gM8k0onElb9h2zp8NpRnQE1nLnuaxZfwNxQXhkfRU5zc
7nHb8fkzJ2FC+EshNX86Gk9vMYw2Yce72KSley5PwrDhRQ2sY9MWb6O2HjMeTHnv
MwPnFwa0+8YfbVD4Gx/4e8GJPfoeYYI9yhR1EOJDnFFbNmpvyM8LZeUEhOr94YnN
CJf4lVKc9p/iSokbeZhHaNyWCH18LrmfIMjr/C5COj1Ml0q+iuYYdDp6x2U0ES5x
jfTDf/jUAxN+4YoVKBUGqUkhfSWy7mOI7zWSIzkJJH1wQe4KcdhkJf/emLyTEHuA
WfLUbRZOnHfRDBbCYc0PNXTtt6cYh88ADkgeBOyKkOhwW/tGCajEogvfiJmgqRiG
QIZckm5WffPZJzMKhQvcmYsuI9t1V2WhywWU0WDEKaXe/Rk0YaFof4/P823NhWpo
7cR1e1QkZxgKJ/bUmbHWWRAUmsNrcwNfYEauMgQUmx69fS1+kFYOcNE//43s9Scl
oc5gltJR/J8TCz/NPf5RUSwe2kNWG7vijKow3pgElqvgiauFiwr55qQHiBvCfiHZ
KO3eW9B5bU5751jWzdgJKf/Gb8vqXCdLitw6LrnOfSsPOSXnoPlEsDh1aUBScDJR
u7uwFeYDFmphbKhwkt4dPrISMDDIBDh7bXTqciWgdbDDh/TdTwFi+8bYtHyIEOnF
Uv7qxJjZ6JR7CJEOlQRsarS6IqKbfl/yPiFtp+h6YNLAaGFJzvq8WaKkWLGG0+zn
vLH+KfzoB2tsaC4JXorDb+LkRk1F63DQS/X95mzxhiU2L0SOgD5F7OmJuVxWzs6f
l8qjEXtiAWTkh+0rmSQ5GYXWzO5648JSuVIlm3nRvvXBfIpjwebjrhr977Q7il0f
1gRdROn38Zt4uXt+T9gkhXGVJSYk5QCDgrAWkjDohnD8xhtkApG/2Ovff4H8hxQB
mWVLFuMFb/s0Yuu/rm2Dl+aQ4mmHdLjE0+tQ3skkdyLJBL3X9/V4PT5VZmtlTwUy
Dojjp99kKuY9oq1aEAADdVmlXFnGqTzG7pznlMzF7QUBJkmxWKohjPrAeX4iKNa2
rTQDuQs8kqG4cFq8L1NwhPF3yX/m87eQ2ytLNvCUq6RKkNIdVYTWqmum0hLUCTYu
rCCb46tdG51vE4NC97iuwa83qPAaEkL322DNEgEtI3zkWty9E0u/r7lUaKB9O4wo
k8XM/n+D2c3UshLBMNKpwsHzfuXgQlqWhbiPUe5EHZJyXWui+HL4ZNvUJWLtYeqg
j3KYO2bOOGGUf/MfHtsh1CTjoxhyI7iJmut9E44HnY1d/xmnm0ptCNc4HIqxYDtl
+HgMWM50m6GwhRcKdRFDl/Di7ZIkWZTgW9vydaTIYjOp7baWm1YlWkUA+xvDVkEu
0InS4lnPqpF9Ityt2/GCWYpu/e+Wj81dFyHel8pHkhe1PTq1/klwMJ1CZLdK0uND
PRXO42vOL7DbCnz2Y6Sl2EtqKn8I4YnRMSscuH8C9EWz0zExH0Wo62FMV9FiOFWO
Z6tHZ7uKaiXiirZgJQBhOuBJnPaSmQbF4TgoR9tGBtPoQcwfsKD1G6PioBPhM7GC
ywa3hmYj6kQ7HE5zhRh6AlPANdnR7IoBbqongF6T8nOf9Z/5GugLrYkcM2IpbxVP
f6Cpq8xMIYV5n0FwzwXv5kx2gdin249z6ryv32b7NDadkbY/USwVUCTLJZbhEgZA
gVClyhA9Nqx4+mjMEMAXjSoeA5GELUITq/F5NWLrTg6by5Fl2hRYFXoCTw8AiTZR
1TkvlOOLHhufPR0FYR7U0uJNyBSturtzbhJt/O5d/ahjrwB8b8M5cUqPlBBSs9ju
NFK2vT0YYjcQAjAy1raDkwfKC2EAkzC+qELZiArfci8YToAP+4iKtjg0iayW0E+7
gm5uqxmhTdCcOmwuCW4BKzS7NlYXN0+Xj5k5ZcWttuxEBrnZNmB+TgOTmp1lO7Fj
LOk/UyGXRFifqs5seV2sALd249FNtBPT8XX1ZIE62EdNuoNHWRuew+S5pjwqqIDy
+sGTo2bQyLrhBQpQEO0OmUB7m/OFEmk1UJpmB7Vfr7BbmUCMKlg/g4DrSOV3NUS/
O2SPoQN0LzhNAzEjw4PbzHCFHoDIZpBHsO8zp8u/NpBh8BWECEiZgQ2etbotoHcx
E1eY7R7IXMIGKQVnuyWjJ+QQzfuZCzo/P9j3WaaTVj2HiF/3hJjD3RM93Ics4tbs
ptt13gnrDfsqv319Iv0tlYoC4rPLcKgELwJsqRtFC5CWNUz+os/sA0Hnah/ASO6D
pPJdJBVGvC5ilIGkvKbPq4V7izATYRIkpO+bsJ4slcBEzQQjiUQIZK0+pigYU9Ul
4JGjElIfX728Yy3J1zSGQilX4JLUW5EvEaPgFg/VAINMWAeVLS6KBWcPv3sL66KL
y7y/I3PXaX7iC8p15bmVrTaxPYXQIEH4S248DkTaWYdrZB6F2ZL6uHZE5mXznPAc
rZKapN+knH/O+P/FRH2W2dr+Bqy1KPBI0Ed8nUv0qGm8TuvhAu36P0e49u4ddqYk
JCh03D8VVJLr9DNdETmJfvtOU0ZTgGfkl/JvmMLZMrxcmtrJ129WzSNPgH4HhW2W
4LtmeVTXD0B9J8qYaQe8XUjFtDE+smWguzsnIxlcx5UCUfA/39SY0m7j7DQTAT56
Cp2S3KrsODdGO8bL7dOCiOOWYITjGZzF19hiKbwGwDdMQTw/2YRzyxwrxNcMwdix
gqGsqTQgTRDQPX8yBUyE93CI3wiYDDGhTi6o3Xuq6P4XVByjI1XkYVQZJvnMJ9FK
F7d4lBAm9QWi+Ss+z1h2BvWOW89MN3I1hIQa9qjdtbokwyxqj1YSXyuuPltZzbRU
thipClPErwsiZpTYI0oGxbhaQsEFfuKutmxWk2dBGSk0lfWTNlsdOshX9uVDDcol
n7+ioDwEsCxT5ypRPIB2q9+D1pIXhDZZlT+xbHuyqyGHW57oj/bQOtMDlVUwnc9a
klyWDeol+H4bNBKmWUE8XU8ds0/IlSMuAStPkYyJCq79qR+YPlxjKZRQyUNCuksL
tEwzJ7pPEnP8Ktbm0FhaSvTsgXwQfoPcPZNtyYUe3UZloNNAOcn9llKvY/1pMtOq
r3meVNHRbFVP5yRG8gSwfBzZG+0+7yvVC6jPx9oLt5J2MVCKMuD+KYJn+5mXP0hD
9FOejrImmwrv2SKa5THz6LSOx4g3w/QhGp/MSOJY0PRjaRxZFbXdMnjrXZWISqsZ
RauAzqF8sDHpxS+B5ksLrQSuHZHC00bd6VH0mvgxJHlhqo4rPco+JRtSpF1D26A6
9KAMatehLrTis366YUYC58tMXLbKV4XMSlRMghU+BZ+zOqatiNThQ5lPk8bQbcoi
95Do9ybxgE/kFp5lpWx6W3YVLkA4juiNX7RZ7zp0xDgSCbHADb206AT+8IS1npKB
AmoDL9HSJn28Y1W+ucDUOicejVOhDCgqGNMgjiyq7wENg155lsxWYYP15zUGrs1v
0BrkuoIOo0fJovbpY6ugHQKfj8JH6BdWtQTxF42muQ7UpKzVX/QncrhBQWg3Zl6/
qNo1qVhaE2nczF4kI4F3NqjNpag/kSmA8+rjXwJZLaIOj7RyTcyEPLYXDgJ/OJ73
FSWWy3lE/KSgRQSMgMve5NAWNxtxiX1ApgJuCvyyTo+e30BEOohuJZ+mI330o+Zd
H+FSsn4pnOui/9s9WYGyRjdYSqvtePOO2Cl3lYcgmvSgMODlHtF89H0JRB/SyWrg
cwENGJGMJQBwxDyglcnvjsRBcT4uoQqHRxtvz3hwlMxxMILZ0Cbf17MYql3DyjLC
WsV0HHpR/Iavw4vVswZLAq6S6uGlKMjNr0R9oaJcw+JNVEp7BWZt6800oEj/hP8k
Tl849ZCC85DGmhtNOz0FyKFOSed1kF3a8nlyeyVQr/0FnNIkzh+Ym5GV14g4LLf8
P5T8IwM559z37zBGBQ5Ea7a5o8XpS0p2aJgV8CR+HBG4iRTWt6WZG3b9Fwp5SM82
IeCDtyE494YFkKjuzmo824eJPLU0BZHJMu1o5gUAv7LwahFpGr6Y7pq5WZmMd2DA
JUn32KPZ5mhJ9JU1b7wv9eh6hETQp0AjAVFiGp3gOsOVbZZY8IGwSoZtfje6puxB
IWmE7/gCercMTrzHTpWiXerpoOjvveIIQY0ObS6VsMOSFxaLSXaxVFV9aJEvuKGx
mdJztKysRcsUKtPnIwy4lXTyEB1geeUhqlqXr4dN+Z+Q/LwHORFZmJoGXnHogEQU
JBiRxuz6r2D4ev0niCXiTqQC53J1i3hTRo/7nfrE9ErIxuV6r1RmA+6coGVaa9tl
IkX2wItzj6+5LZqrBuWruLNeB6UL6w+EhbLF3pugmaPgAFzDzD7laiLBJWhNe4kw
fACM1Oh3kHXIDAiZqeb+Z5p+I65J30Xal73I8ElrKV7rdPgT7D+G85cuK76G5vN6
vaxJGChhnA+caR0NnqeAxeIysu3kz2VOiRhFKcLcbpMEue6+fpe7OxNn4coUiYJp
Dp5QzDioLqisoV4Svc6sfIs7bKbK0awVKMHKgQ7Nyh6OkffDWrO4S+ulck8eNHFn
5D71oHqqPQRMMbLci/WLu1iA8PaQZaT9zIQCiyMPXv5ECgZH3XrXA/71kEq2DFzJ
a1DFydL2JmzMKoh4JbEh3UeLnheS5/g/TDsVfWairRAsylYwe9j64pMDS3E9Uzn+
8ISmcKBufMFksx3t8UP3M0RQN1rPsSeLj+5iUbbijLx4Vn23CebB+JYrbgYkRGoG
3LMawvuehRSMYPQmdxt70gYupEcpbfWMAHM0IZNqk6r6693hucEnMgYm8bVP+7+K
SGYorER4sxRCLWzqvBFuXQzdgQrwjNkPNdCc+C3N3LG4j3meZyqsXLakaDBBU1FO
RXKBKrD0wvT36gC2WOp0dA1QuJmrAz6ktIlXiWDvteVY0m0nyYWHYddWOOoGbwrP
NfbrhPT1fTCfALYQf1gXIVqgAevhrw8sA14QSVWtdZp9IZv6sWrcFwy9zO8uiwn2
l9YdU/xMVnjRO7NNoJazIaC7tT/oR0zD0XPRUQd3CTMnYtbUpDfvDhM9bG6zFwt+
fLEEVAUyocIYh5I4KqnREOllv87N/vopG37PSUXDxYTx5P2bPEaiTe2c0+8ar5cv
Lwf9CuLM586zeiEMolQj9eGDL2zQ3D8bd77dT3FnZ+LEC5EXLt02tvdWAuQ8Vl/6
wtSnjxmA2KVicWsdeyiP2JdAu6irimtsmxWSVwtZIlhxIQMsDwLo8OyHf0CHMzgO
RGCP6xjRvk8PWlBGsNu92hi/YtHjBX5KilFW1YJjDuW2EVlfri9AgRlVoPLQDQqA
c/+rf1FSCB28XMtzqUvuFPL0t4V8gs8rCAJhhkD6bHs5z725f/rJiQc3QUDTNC17
vx4M883RbS6WoFhj2NX4k/q+qkI5FkDUHDzAuzwF8DDbHvMZzT32/jj+35nNvesH
DVKJlng+PR9o1SVo4T8nmJWziWQnW3nuowna4l/kdd7U75a3G7BMxISy/GdMQirg
bRanx8n9d+93ou7XpN0F72dAwz4uUGqYN8aEEsOOpmfkPgdKLQWsllAgMmgyBJw0
MXgoF4mHgcIJHNh8csKIUU6Va4AgQXQB0iYG/URPEkcjR3QebhH2V0z/M4rfLeTX
4yr3mG6UMm7A7sJ3zdjvcVIM2U2LemncgYUNTPISr5gKA8Kg2LeUG6KW78lJ5mE9
pQXVfYf83FgaXlToPcY8yRLjbPT1inYbEN2o+9H6ta/CrToPp4nFlOREbMCCH+30
wP/5wLS+AGlY6cg2w+jT6YuOEIxiKLGL+iwZ4dIIAxs+38tnNgwd6LpJ6L37RdRB
NMG80B19jxL8/Uf4P4c+YP4SWL30RheaV2sXGAAsDdHMBb/ptAIjXGOL/g6FMhyW
qwTnQ71kZ59f/Gzd/pfK/ejO20KqBb0/tbnHIZ6aezmm6jhhqtojuS7nQROPVPN4
i7NJaYtMCKcG/7QhpP3HQ9zE0TMo3k4S/rYsY0lrJNDmd0pWTYSvSSB4+0itOw/w
DI573lcZB7APa0N1vHkfmfUlPCtVMh/yOJZO5en7XWv0hRU2npa93fMlJWqvtdWf
j46mBAu351KfHrDFFM3rtRNPLiKDEL6Ia+Qw2/8dTR25nO0hXizm2hLmVVE+UuJg
7Bni4eeHVQxWfkgHqkoXPMHYwG9vxVOC/uxVir7XQU6TC2OgtEdwp7lx6XrqZ+aP
zYYCUd9UuMb0lypREmnR3OEVnsXgpD1btYgEvE1ug7iHV3H+UBPynW7VyaL85d6d
eD604vPMTsY6SDARMJgmdpecfghtQy3lUvdXeugIt3RDl8LOD/qIb+L2R03sRk1c
PdP4Qima/qFL6a0zhCCdIS3QQFD0m8dm93zhhwKMV5Ygx0Dqr1D/h9kNNdZJHJW+
56oM6hPQQqWLP4jq/21Dl5sc80FWjbPKvh6CwmuVAMfddE5RClA+ESSeU/jreSGA
6YVMacfWYngsBUk+cFA112Fgc5cQhMljB4aZ96C+f2psIQwvefPU4X9C+GOeMF17
M/AlJ2WDyDNUsluI1gbIxIOptDiaLsIKUpU9mEBvOxF+iYWFUc51LRBsL+LZYfyG
ubJKVPo2XUhWL4B8EePhoxdSL6G02ZDjisQm0+t6TpBzpFKh5gaGYYF7/NarGmR3
xcHPAVvF++8fCVZWoVmJzMgEmyGE3MdC4JNC4ITGbCzl78jNPi0EeStZfgLCfskD
XrbpKvjmHn3npjeHg4h8VnwFqLpf2HSHIGatRDn++ppRsuQDFGXaEMGLMf9O+0au
Ed0zmlH9RcbuWqZeW9B//9K/cIsbyC4yF+V0GhdPUp/FZ2c22CrPCKmJQouVcZ6A
tJAUJJos6YGC7xVQBvH42piWX31zKQMxaaz0OTWwIjRnhUMpxFBSWZ6MUgLFm/Le
hfzf1Pv7maUY9YpJdHIVmENokp+tblqZOGnU93GxDFzI9OWmKPESPDL2aC1i4Uv1
gtgxQ0c9OmvBDNK6GlemAQrIYdCBRno/W+uOAkYQxUePriDctD9AA3a6b89VOksO
8r+o2t3U+cPw53lcDkKt9bLZNlej9SZWAAMHnMlEdKenWUhPJOFidZt9XSeGfE9q
r5pf1rgiIfVnDIZ/NdokCRZBJAmuo/iw7AMPJ8ZhY6206pzrted4W4zv1zhgHBRW
h/CwevRlIytbPPfxhcFfwssFQPdxui8/mHArlNZNVrgwU1AuVsEztH5/tzy+1a3O
4RdoBTBKlaGI8YkHnW/V8PuOtYpGIP2E+LtBEB693dXdQdVV4D33x4GFWr+yzOge
DLMCDhbUMM98kMvUJUjrcpubVdZY5XwN3DSDVsWkV+AR7zIH+565oRwPs8wI4gcW
eMcfa0Xq7hdXHfnV9rJLwlE8jsNcBxvnViKJSpp07ijWeN8qJ++G35vKide+vKDv
b02Nr5DqPFMI8mfHFoIYig4gennllYCoMddEhauCZPweg77MbpKdSyzswrSmmJ+9
bw5qW9EOk9NUtinEK6xlHC5ztKb9PA/xdtE3RfnieFqte+n9lDPm2gwoA3BvFOln
AFOy2Pa/oEpo6PxwExTYBHR6bcSEc9yMx5U6gBL6QSnHyVDQxO5x9dd6hKrVLoJC
zhhCh12fzwm7h591j1D/3VSFC0TWF8qDEtEdb2r+xFRysd/iKX3YGmvF5JfG3YDc
UvoR4tghNAFZGbKVFUCeDOhds9s7WQQZWLY+DS1fJUkfLDjTCbFFFn8BzHYnObc8
oAI9ZOh6Mgaxa5us6NxSLhnoA9ems5Ad5kcTjbRizTMaMq5yIlK28QReFp9JyQpR
yEJ+ThrSfkHsgBFFJ2pevqVeE81ZRCJ2LSsQsE3ehID9UhOA6H34XtHPThECRhGr
1n6NZk4/kGA4pNz80Ak4OD8yZ3LGWNzG9R0cXMw/b2ywoH4Evbt65bBmIE8w4pJu
z9D6+6I1flfoVg8CtRdYYVSrMPepdQtcSt6yXLBdwbwZ/MVZUD2jSBesKFZGwB8O
KTCxLN7wN+9M29tq4LHVbGyJQmUQvdEZ8bQC7+YZNP/uej8hdO1olYiXiNXJNboH
4Jn66c4ZsE79d5jj9aWXCCA/W3czqSt2FNJ66i+Rk/wYS215sYC3njGTkOVzwlQZ
+xZoaYT5LR5bd3WlDYdRNUba0hUYJejr6yG3z9cVyL6Ge+opsDsS2IHsO02m5+6o
1jgKNNyo0XVaTd7KAXSN8WFTx+x/Tc9+hqZSNOSr7iBYtZFsCVqqcX7SuV7pcwi2
4xcSqo8ShXkQYwWQyJoThsC9F1ih2h69f3qOLQ1SGa5DF8fgAJc04zREQYgke5EX
QwyESW6KCEvJUGJopdOAmFix6l4qAMhD6xNMB9eFzQR/W6uKvFSFXT1NmoVb+R44
7c/x6J2vmh6/EeJzaN/AYoJq07+I/Z0D9T98+a2tEIk84qIVybZnrGVJsCl2vdF1
XCnZZaiPfo9+ZgupwBOe5v68e88igNPbuZGy1xvai7l1UlqVp8uUVKnHUc9hsow1
q65vbuoYDcKl61Yl3mfB1nVWcV800CrNmcJUWNOg9LewnVLiCv38XjlZq33u9Myn
2HmzxnRY+vSLd2uy99/jIGlLeXUoqoHEmLL1UHZ5ve0Xbre0PQI+EKrfz6tzH96y
k8avKQTLrG4k9yGjcJDayGKL1l9qpMqV4vC7Ud7DRSVmtjcpjxDembwAnqJvDHKK
/R9NuM219lSZ9TqMvbMim/QfSpMXHm9QywPvQe5SMSVTK9DCvmflBUoCQzNSHN9T
apU+evz1exjRea/nKQJ+D9hRl+UA1TcwXYVnbIeM1Oj8Ivd7nN8r2pfFwubySIss
yZ6r+sZIOsPro457URusUDTHUlebmFwle/7xC0tuM48eFapg7eB/xhBKTzW2KuNb
62tNq/fgeHCg0Tq+1+6j+or5LSmJUn82E+wO+L1RvCdbrDTUxy4NiBV/8Y3PcS7k
HWYmuN1NvBVGhuMPJTlSmm94c03cWEj6cRQGgpT2zuMbER3y13upILNAr2YutpjO
a+j6WZAxHaoBznK1V6LeNojspJDIkCnnB3mUV/knTFLY9VFeFay6VwJm/UONpcmp
YMIZh0vBnOMey18EQqqSOebJkUtD7D31IFDr7A6QGyt4a/Ow4pKcQe8eyTbsOgoK
ietZXdrJN//GfKPy0nO9/6h06dT8wPKXit+UbhYjdOMg9p1LSF4QaO9OAVgAYeNd
sXygd1Tu9O5yCDWMaj+weJ7kYs8As8pTUsvtVcw+WcKPjdXJlD3IMCFWhAcuz5qB
6lCCOMcqPZbcT+NTL+5vMX8es0AfBUeC4bU3FFs2L8Dv6o3DS/1PknLoB8FJMLqG
qTV8SJHW3zfzgahSP44L6t1n14yaysE1P6Ksw2aC3epH/YkwsSv8pAVq6yVDeoZI
8h8Mq3SFibQS7DNUCg8WhMLDzKjAvDE8wNo6IjFDaPrA2y7Dum8zSfi6bt3sFksG
NE0v9ysSe/gJq8RGQAaGXdtaLfNQlnQpTg2Q1WPhgURIE7kBZ+lJ2qHA7AB9nMDI
hbgkNEpIlXwgYgsdK71bFkWSwZ+g+oGQZdYnQ8VVEYgdo7Q7GvRrX41PTk1bi8Rf
9L1+RsXoG5pvUhB9sULtl6UlkTVaGjFm7NIoOHAU6LE3KN9EUkRU/FGhN7Y23BsG
D+WUC5XgzL0BkzRyTMGHdXa8Udra/pZ1BQF9eQ7Uva5jpda2tDQGck4kep6ipdrM
NsG3WqWww715pkGGwqrxtiri/JSSRWBlOB/qoSR+987MizqBitUu2D1NwHbIy07S
STFhhNhs7X47QmQFck78Y3atevYVDsOe+h2+NaY5bDXsItKXuU6U4zwvP683Thn6
hxsEaZ0XK32YBEquokmNqXwKkRrvrIXbm8e+Kf1PjLBdP7x7p0V9LKNFQ/wqogqq
54spU0oVNSLxW7Tmr2S0UJORjsQIJOweKjOUJ+YtcdI6YDc4c7xiT4OEMS2qNcoi
34PvqksKjdYzhmOzaWvzBFBu/GRhgNXDcE7HY4hE4R/1cE+HhNI8Hj1rr7lkx30/
k04Slun9t0MPzT16MF0SvxR0w2Xw73Skd+v9Q/2UYtPAiibBk2bdtXA5GGwYRkPO
r5w+lQTidfVurfjmsOkOmS2qcFHNvET6r4+i8hAWIdRqVjn4XRR/6E4bMaCHw66I
uG0MjVJQId8nWn4HWVck9VQvCBTsZSBg51wrP6o7CAnDtCurxwGaq65vN8cCXTHf
hrgH5Yl/2SWITds6WqHEdse82SqOjvC+tsNFaj3fczLMK6B5LyeZhaY7GV4WqXRF
iRPW2HbF+dJ4XWi2651a0890a+lnWc3/cxbQYsMSqWFZ+iens3TgqOTtId5vG3EK
PaDQRJYo2SJ9FQcNWEk6hAB9jNmn8bb09VjbhM9Dfg1nUM5MdCh5deG55r1E9BF9
n63RquC5S9qEvKgUjKm4859u4DIxbGqS9FG7R3XrF/JFA5XACN9Y8fg3V2HFa/K+
GcaFo0fJz+xv3Wz4oaHD7/Jn29H76Czf1GKRGFvoS40V74AqB0hkXmy+KkNOzbnZ
SuX+of8ynjAAG+awXzjiJYGkyDJapXl/bBakRi1n0TtnUh5yojs+Cf4UjdRZ6QLS
IpUxi7GEnDT6eTi1KTNngAwnwldwIg2v59H1DlfYNoOkh2AdrAh54pmPwwJfytQK
bvUKPPGUwJ7C4i8iz7+YEBNYrEYrJIRAKAcjNTuaOYhQFmCmuL7Kvo9i74i+hV5T
vaezLZP8cfKRiUhBkQ4wE6GGbi7LJ9wxU6KaG8puveRHgTkpdDq7BShCAbJUq4k8
7gJqHCB5ed8alWOxmsFy2Zr8oLuVZBfwAtmlqBDcOFT8tIbfsD/wIuklt0GYq6sj
2S6ylin7Mn1F7oIEBImdqVg7mz7C1n2vx/zEdROiI5qpA1LSWnQzpi09cXCebwTH
YhDGOC7gEmN/7nq2nXxFI9uc+dNDM4aBMSDllcw8lhglsP7PMRQ0lsDtfJKQpseg
fQG3ARCs+F8RI+m8IBpwFf+8lgm/G1+uObGc3CSDO6rGxZrO5OfplS5ESXEmuEER
x5wv5mFYtdBwEgkPDiw5e7Ad285GbcuXOFjxqxu+YDDktBRscYeo4ye1gkWFWqgk
Iq9FFUI686qI6zIXtywj8SFearj0N8iOALccRIeSAg61ck6dTKFQCGL58wFibbqG
nT4tAOMKR4YSY9h86Dk2+vZGe365Zb0Ikt9H0NBoQWvD5Il/VDZFPeMBB6Pk+mh9
jYnV3plneCp4Mh5slzghtafvOKSsNYj5FenRghqQgHj3dXszt5qsfgzhqPtb2zno
SPUUUkTHtDRJzvXplw8aP3qgsHue/OuKatf9H5moO03hpRD4/LZE1e/fUu7TsohK
JUdTcTqFwL993tgbgFH3bC3xZDmpjscMCt8J04D0bvPy+KTYJyN4QkM7SLPkHv10
7MW3vRbvbl2RyeijfZ61jzbfenID9EBrzIikEY3rznO4LNDhoihR3q8Yky+wdOKM
APaEWgOfjZy7p22cZoigPApt+8d7n2gbdurFUnsJ1I5eqOohmjcFLcL0ZohC0eJ6
uzjht+WzEzghJzWkWsZSmDnRw8K0LYQGBmEg8gV4kDk5zBVelOelCKk23K4gDSle
JqWnn6zrAU3Dp/11MNbp6nFTojpFpLzLxlFljJ0EDuJPqnqN3WpORt4/OhVL4g3H
ZnbTyagMzjTJx5U2MMw4f90H1+JD7Sqns/ehNiGYz4WvLMa1SATF+5SNNzBlLcDj
DrRxYaPN8avQEkw4h0tjMPst09jmcc0v7xMFRLAxcrgdPdznsEwUoQrPxtlSaqG1
LRcUcPoUlZM+djsu0GYgyMWBJhFGB1ZEf4fuugMVkj5pR3JJd18CKr5MQULNmpdG
32NHGVjsbjbqi0rnjz9n++qk7LF8lKlRXdME2m5jnH/UnxUOBu5UruYp57FbK4mg
z35wmG5fF+jr0vWvWoKJA2PI20x18/nt/ii0VYGiSvihAtLL7Zkfb8GCLIOWETYa
xqmohOLsIjnK8nAEDbyJQRdX19xxuWXhLcDW44KCC4c+bVTzclmO0/Kyc1/woUCC
k4L2DD8IiPfYtB+C0dr3TbuonKRRppWe4XgtWN7uND5iMdjOvmR6mBHPe+D5IizR
OX5xEPZHPgfti4fulolisgJZvbXhFK56PxSBnPsXZeCKnX0Q+xsSwFYESb1j38iI
DWT6zStLT27IUPOdQCoy+uP2qp5CKy55q14SHYEeGhIxTbacyWOlj5k42Fpk/oVZ
PMP3uGgxVFWxAzomz7KzJKNr8vBEpZ+mtg/OLqAHCW+NrLQe/zxo53hlXIYUj7aJ
nQd19fbS+zZPswuDy0E8XzDSPqJjUZDnX5lcMKoyGu21odE+MA/W7bLCPzZLe3Qk
k3SURI80aQnN8Jz2mUV81zJqSi8QQmyrSkw64nu9K6EHUuE+1XFsh96bv62qS3lH
IBI9oi3mEi8+n6O9mddWm2T3ZwMmcJceUJLH/qEifm0esVv0aN8J5482Z7bC/soa
CTs0E3JF7abH2XaQn/F8+e06/19v2ycay6MCCGK4C3kAUdOCF35/uzsmmuh4Lvks
CJaDz3j5xf5psneWya5UoWJs97qloWgyxS50cORywDPq3UReaySMZ1xb+wUwGMJE
2OvVWEK6YR0THmCYFt6Le5CCkkQ/bWa52AdgDlitUYQeCab2zMTjZV4x1yn0PH9J
4k9J5fkDO3SLwW57ImAAh/x3S4Nkx9gWWSghzY+QYqivBzr9Fc+2/HCZrZHW6asw
Eqg0x3axMVVfeYu6QTfSnm0J6/aq1AQ4MIDN96U0whEce2UH2JiDCrbtetY/UNWX
qL0nxC+R99oE3RR0M4vQV/ISSZfjFDe7axgk12TufI5A4KaxAK9igHO0bz23RwIh
WsFIYqwa1ehoMcnuUewT7NFMyOmyNdMMc2D48+4qaIO9+7k+6c3QqCwWqFgps2MU
C4VKnIe8VQdTV4ndRZ3rYT8nloIA+rTO8BeB+UWYQgiXh3j2LH5uLWxeQh3UkEsq
V5scR2WkKHvULK8n6jPzs7InZG5wCJy/g2TxCOI+FVWLjxTcHsLpV7FW67tdg75s
SbrImZ1s/uR814oEA8Q5EgC58S0uo6krBRv5Zh8sIw0BPYLonM8tQWEQWbhyuKdH
Prmj2vRATvnQELt0IoepI08QYBvNm3jxmomAXrnGvF8Mb8ajWVxRfABdnONznTny
FBDnI2jYRfS5xmAkDa18cDHGa53auWV+iYA8gAPMyGp5BJY/2ptqWpj4meRcExkn
n8L0jWXfBwl8a6/5jnusRbIvw93RBMo0yuVhAzhMOOVrf/luoEUE+IEPxHxFT8UA
27gLhELcVMFRTi9yX3CHN6Gh9p0Mqyr0KiiUFj7MNOJL1zuPPAG/bRd2/bfpdu6F
5jwOZE/XNeRGGMgfr6Z166TjlrxJFpDFuTApnSmQ54H2j/7CycVkS54Dc/BRFuq6
yM6KnWq7vaCB5pLY3DIzyYFFNvDAltW9alkcp8lDrxxGl5xlZ2xbJ3bgF2QAfI6R
1hJxT/BTf7YmxSdHqfL5FcuCVzzxvdkeUol8EEDlZDZm0y6zjG5x4QI1MiiFdE+i
r5h8i3Q7SXCah9G2VMvAG9gMyqQjmhRviH/ROnNNKuuRYWd5nIK1xjGyMlZsZNBu
ZQwaJ2fPVPyw9jESDlqzMmYwOB5VfKcT6BeuYPyzXFfkablePK4nYSc28b0KIDYS
qvGDWck7ot7wYY+7UQST0wTNtEYnxTvIKzvPkrBa8zcbgERDvUyw3jFhHMVGXo13
ulInmxr0CjtgVSnEs/6dm8oxe6sTuswONe86FKg6qA5/ltaev+h9BY+oiQXc62M7
oMSk3v9WGHX131en3d0wNcCbXn013Nu6SmUDU5Jlro6yS/tMi16vKtPdwCeWOv3u
0zePQcehdu04zCrFxtuvhlrTXe4L5uXXzkZfexJlUjlFxtWpO6gjpuzjLGKvw86J
tIRTnkCxDW/DJ5nd14ioAN5+eO/b6XkgL/Bu7rJNULvkiJKDlmNKC84nuRT56MAl
D1qO/zr3bm6IbcJHPSQmU8dxacJdwdJKP5MumiiHBgE7tQiLBgmJ0dCoPZpWLKiU
2rGrf6UEr9UZHc/1yrfFa+HKW0we0DkwVsO1yUtfDhP61AUziOQSuKh2qQJaf6HK
QYDAcAWUynMezHTEjbfYiiww9fvaFcxoNh9sjN1M6TuZNowFJEOuXGdFYK3OYo2q
pG7Rp+OfwAjU6GIFwELHo8HCHdo1m/k/d/jycK9ZmvADcP81l4OlrrQwC9DMCygC
ebMOkFX2JqF1uRiN4o888+708kxOhjveAquK0ddXR2le5G/p5gFIV/nuWS7oDB2Y
g7HtkGRtszWgjo1mCA4zMIJyBv+B5ZZmR5LPfWX3Vixtg81rzKTV92/NUE+mHyQG
5ofLweXM4+4q6s6nqDkvZ7+km4t5q7PsAVpFkRQ3T5EpK03Qb9kU6/oxTFwe3AWM
jS1IFRrUz8MntZ3ECGVY/VvYpQeOS7OTMF8J+ZutT6E/4OPe7f99MmA0VpVXmGbn
UDGlMCLcc7MqZlx6n+nDG6b9wJBEXENLdyM7ChLLi15ibTB1wFrSnH1vRMw9W47V
ixHDTXWd4GBJ7RzpqWQyx4JqnAcB0hNlyo+Cach46qe6Q09X8OWL93eCZ/dTtB3g
RerHSKRhDJt6cnxLMJHJV44NKfjlSjaH2z4BlFVROyFFkOKUvCqbFQzDa/HOyIfd
zjFsAUnmyp40ghTXwZDW8qPn038XDPVXayVJN561gwwxb/QyNSoPYtZ/69Ny1zmQ
+03tsRIvOsKTtEA1CA3hBKfgILBLdLTyIjSaUMqF9oBGtVBLEUcvEn/3nLiw3fnZ
2beft+W6aGHn4qxVxeD5/Qjiq4QYUGbEVf/XrhL3iYOeMsqptmEvjDwOfzoaE8gp
nVOfYjCQiXY4SWyq6jpXnVUrov3aQ6kDXMyA06ehuH6dKaNhm9oD8zCFbZObTq6X
fEr4MqSGkdbvu8DmAgw23Hq7yH32FMRk+5uU60+fmiK5rsZ0DFIG0hHBMu/ky1kX
iTSnnOxET7QPpU9LKF5eMiAFbmveXcoIn8cN6nuBuH7Va1NRRwuYxDqq36DErXRU
URCuK2Hm8V8gd+3WfGYV28w8P2Hh8AwwLK57OqIsvLi4ypC/sf0MQGvPTxfFoTnS
MpfBQLiOYfERp1nr+niqij3sNIpLT3AX0SRE/R2HV2j5nd2SMks1ajVCSAIwKq21
UuIfCasu15igqiNqdFFtjMdkpjWnUdwieD7iGKw7oO8XU73U597baHkY/zYuL0PB
xjR0TkIaSxGaju036REkzOpYuNgx8ivdDg3VPkC98Hhz01/hvrR2qCZ0zlvISl58
sqzUCpDsw4/cZrZKCIdUOb9RiAwyERHED6CzJouTvTqRr1aT6ynNyGyWZm/xZ++2
Mt7bctDAecyp6P9cSg6c8ZfXbqgDxUd++idqmtf6S560/mrm123pgYa7qAKW8JV6
rd/pyLuD2Raxx9SbBdAwqXKmhvhBs7uG60+5gVmou2DmTXiuPBjgJcI8sKZfHB/E
AwsW6fBQAA/dD1MG6wGGD5dBRcilmOl5Ve/R6ITjNl1UwzVrfsAUW7oGf9FIFdAE
fQg71CtlHTl+yD/+XPXBZN658gl19a6RswTjqiM8E0NBoBTyS29YknlgIXcFsI6q
O4aCIej6HxwHyABbWBio1qvAw6FXePYKVRLf5+p5+ofMVSSf0gmmAMJDiHvBkCLg
KwzfLioy4ZBNakeGNEeu78fnR55nKLVlzOzJoFCBPO+lq8bKD2mOiJHGRswRGdsW
gmTXi1Q73M2O/tZRMxnyMi+/pd5SHARdzMImw7aMIRzLK0IX5oT4H0Cfrt+KvwoZ
m16POH9lfwQ+zS4LFxKmkHOykAkqOAcF7ByhCX9FrrjY19NsL1YHQUfdk1k7I+pQ
aIg1gr1ViImhIHntePIDr7hYgMUjQHUXqYzQRZIRrEYitZNsJDBPlUIDcwFEERKM
1VDPq5x1ELZQluLwCHXikUCaeELUQjk5Nwn4j7oXppZooAWQYwv7ikAMjbs3eLe8
vgV9iUt214hBEaJ0sWtwouLm7OgBopD7NKgR1s9Tyx8Fbf/omT89vPGKGt+TzASA
X/R9R16luiYkjpQOvFC5thYxS3/LFBRufhES1eOEGCjf5Zf2u6cajIaHkJYdLJap
0OIQN3+QqipyjwhDw1+8Nkn9ENYXNjnppYTZkjfE/tud+LtLsxw9XB7251b6d9Q3
NUPfkL8aZmTfuE0dk5RUgPoP0C0Co9rWUdQb4hdqpx/7piZvXo2wivWOAfHSPI6+
N/FHUEGFg5UxEWeF/8SSSm/H858oKXMntP1c4lCLd5g8FZBRCcwJUtDgvru31cM7
w0KQaEhokz8di9gFe40ZB2ET3V1FnL4Hhn/17g2NVGxaEXPl4Qz+H3gZQn+BDoxb
DsZtBmYJOlnKYqYU23IFsXBZ+8iSDQeq1j7HCbkMeyANG2FXJt6PBHsr2KZHpCu4
WvuBwAJ+ymNUhKRuGYWGldgJk2AB8sJiD0PcgepSZTpvu/3C1OL5mtM1o6v59zq6
mTSF+fVg3fTKRAgfBUtI5qPKtQz5456WipNNS55HmGiepHqX8Ob6vH7vN0SB/y+8
8Bg8GDfVXkK/O/yrCFaIL8l47so4XY7RMUCgV1DMSS5gwbOMRWWIAvd+HVhfIjIw
taVn+QEx269T9ohuxxPj6PImwngJe8qI6MvIB6KrWoqIXn2RwkZlztoLYxejhBX5
lrDp4eIHELYHWfLyAPdXCST6A3t1laskBBacJqHUfoNcpn3+NR2wTWre3zeIFICL
RzU81O312vL5p5Ev35AvS5Zp2AJpFV4xWzL+TNF4GJbNKAciuVXCb4How2MVPbHo
AX6NwTBLwIUPN8w9KVYvpKcBWR2H0cm+JnZ0KQkyaL+d/DGH76REvpsfuDkZd2eK
YRkIMq9f3unNMuiJfo1Yhg7wMZVoAZUTTlHjyQfYaONLnZtVc7Xc48BxOfYcxbPO
rEublDsHPqmvZ/TPOqCBBXUQjZ4JfZZJrCbv6XjmXHktsRNjc8b8lD60k1Lkz1En
DhmNmcmij2gZHpqBhUUEPVDOTCb9GTk/jFmx6iVSRVlhOmf07eRiTUFbo2QiD+6H
4HZMg776vky+spCZOUpnwG0N+L5BdUbp+9kL1i22lpTNtLk0n7Bn73AEAnTuwLWF
/RvwpO/2xoc9yGskOIfOb6JqORKfQTil2bUN+8M1ZeCFZglaKI26PqVUQ3Wd7AiD
921SqgwrHSj2pw7WvaGVHP3kUd42alHVQTEsIMhqngDHbc0ZL7ZYejlNzas8VpuP
2z1d/ncSZSohOHxtrILmw6w+PqqDSpVlIQCsntbK6501aHaPrPose7USY/P46724
+bN7yk6ZMOS8eAB3OkmWIdjYcYpfyQ0ye7XMZm0Ow6Wtw4ttYpY6LBe0h/19IZBQ
xpU/gl3qJg8+t7+ATB5nzvGT8uxGhJB6lxZ570N+Z8A2HqLbQHpnziykXk5PbLhO
9Pv0MJ75cpyLZhfP77l5MeDK/kP68GILftHUKxB+lfvJpMX23A7v0SA7TACCNzap
d0ze4JkjtXdpqS2R9VCd8YY0lZnXWapl2tzHy6RRAiWDJRWsJ5YoQ/hkLf5K99jA
HMN09oTTne5cGGDEbe9xu92IHaKfE3uksbgTwK0rzIQdJrPrGpuCcxzxhR0S+sNT
NKMHDJFztcRgb7Lyrh8YEkkTD8I68bx75bzXpZ85pLcEY0ZWMdnOq8g/2sp+mMmw
kRVEuPB21Zve6j9F6g890KtJKFzuZAMF/r6j6mrlhN0E08y/krm4vLHJKJidO5n7
HeRK1xaRkQNSZKuZdDmx0OD8oMcSQcw/I528yH1mFBj6MfOoeBIklGZJgrHFxi2w
LnmgzmCE4g0bd91035SCVMHKoIZQNZRre1Tk7aUbGQqbDbe3ALJnQN/HegtdfYVg
Vai81UWqaR/NEzBdhI6Q0nao075vmPszpicGWh7kb/qpUOtesuhZXTmaqb5y47hy
Ma7drIs62w+3BLzC2LjavdR1/CANf7COfs9cJNrHBxhDxHVdxVbWw5A5oMhpZMKD
zI92S4ODjjOtuq0bYS1sRN9LwnGFDYN+TebUvRgsiuaI+owuv7dmdGjCsNMGOAbY
T3LkwRmQMB62z/dyMgtcu9vYN5TVAHGwyf9EUDnXWmhjZjL4kWbY1Mpwlwm33rIw
Luk3jj8j7Vc8Xg2kOtM+qy+NQmtFw7c7VPeictRKziKq0nglolQCL+NOP9gYtsgV
h/3QUQqB2VNNYUNUT6CRlAJUnKXXNWIFmQDWCtFsqsPk852H9gUgbmDjrIqdoUft
QYWbH0AteJ7xGu8JA8X0u3RIyjdw2DYK2fLYj9b/n10ZkT6i6LBZnwa+9jhkmCcZ
oGGyHLCFXuEqNJu9np5k/8kbsw8PywHHEMAAQS9/tcmAEyWohl5XWUb05zmdglF2
lbogN4ZQ0yMp7rTtvJIhYWUafjDiuWUaNzym1Hv1+UUxxS61+hTxrGjhmM93wPzj
WLKQwjwpjZrV3Ed02La2175xVSU46Usrx5E6KcGZ12+YS89gmWHzlDzRIloe1Z6m
SnaU5ODYDf4U1EhK7D7Ukx3bXlgHOFzMYWoM8lrDK5d40lnh1zv77+FHxXbWKu9P
xHXR0dQDlbzyuXHu7XgKz9t88Z4BA948Z4Hb4vpPf3hv5DtLPWHOOXdGS+98zKN+
w5mZcU9ZNUnrcd0SWrf/KuV7SaL8aFxUSdZA6iE5GS7+7YQt14ojt2ZwZYTpSu1u
L3K1+6vFuxCCZw0opXSfoSYuhnWtwq/bJcA7wBP6hxyNU4HSN2FTOsq/3TxAAXkF
p2gep3Ugbv0ItR9pNUkxe38szXMLpIM6woNidSPP8zOuzxULkNMpHA9gTYSDBZ4n
sHxPmygKX9NOzvThG8rS4RCLTxlIVx5cjKR7E8f33QUGVAhLM/0GgwjgXqyf0BNR
hdG4XWSXT61nGYvIVq+Jo8DVTHhfOMuPx6uIVbUjUYWObtlOtGWjzHI8hNFIyCCH
avYe7fwz45CkdEZLVGqIO/CohGqMK+8zJuLZYTVqRKdFqTzDPVTJH9lQf+ujb3xc
Z12j+cFXHmRmcNz9O/jrO3VeNYfEH5mM+Fi97H/7/yqyVztvcldplJimTKJkCYZh
EGr7fcquwrnd5Ta8mkZcdLy958l3jteyGWrXC4pV/RCOIjwSqFcMCpZDcxefgnax
P9lpaijX+FqrbaKGDDswEMfdqET3c+VaX76lX1ma0a2SXm9YDWZoypg3YAp1o+Fq
EbADgnqU3fleqHGI4JPC1X1J9BM8eb2Qn8pqrARKUt+UC3Ox1Rwg8g1ZERwgxtVc
WTvH8mD/V6suNYEsvOMi6pGRiULiPiznbhJ+XTi7A+fTsa0+Ux5JdMb3THhohNsQ
fnZEeRRkEbeMGDtjEq38B3TdeYqC5DeBeNQTdKRhHrFEgfxFiRY4O3kaftZFyz03
gMSqSfvFqBFg8xhIssbPVlOZqUxBLkCV4Ak6Vje9BLaEUReGweMbnVZfp+MggaNY
SD98MBcouPC8zrsT00xFWAIfuccaScjMzGYzwtfHJOudvnlWQYMSpV358oKROSo9
Aw1VYW+eXHDzNeDAoZnq7H/Rae7ideewY+zWSTucqXyZJw87XtopiR7Uwi2tM2kc
E4w7ySDWR1b+6VJpZ9bNKmtw8PC5L5xgxfFbKUN1ugRdA4I6BstCiDxokczxVtCQ
kS9qy/NlBHZVtTucYWd3ufw8WpXA8kJr+Fw5n/siOd8UJQd4PJPfc6C6cALqiZZ3
G8emB+rXzK4Xo8h+3ZZ2TJzCsHajiwQSX+lzSU//PObp3PMFvtvrjeAapwJfvQ2L
mnMs0xoOLDJMI+jz+2reagUEOOhMuny2SjLhWDow+fip9xK19KCH9jf1/W7kktE2
OEKzUbS+U7UeLeBqvVFcbYIPILpCcoiGJbfU+QhKyVFuKMd0HZKngrsm86fiKTiF
RvcRgQ10SVwK2K54B0M8GsSPs7M/XAsvoaq81e+7TBcHRg6DNjQZkJYQZkOpun7W
GTHcpYchdFpN1SXXVHAWFNlU0uQDs5L25XTaOsDff/zBhYQzwSOaQfuYt9dmoKR4
1jNmpQ1owSUDmSwPpstk2nAzlLwf+JjIaaCCZ4B3lyZxEVKGDSGi1cnxRD0ddxsk
N4xH2FwgOicSp+TwZW++5FQYPwpmY9vMD3eux9kEV+ytD5kmkoQoJXBVAp0qh6iy
XvI4cL2sHmDfR4m3ASt9FAhgtTwpMwwc0Gpl8QJUtX6OQNp0943qAMBdEp/dgsfz
wYZ/xZBGyXlieV7N2v5GQxDdGN2hUvibXZHVaEHILNukUsbjXUBJUlOcZ8GJJjW3
xOFX76HU7ZwAJf9kz7IGL0WACFqDXy5vpEFD/HIuJMbMEcxp2w25G4FS19aM+pQe
epqAUBpn844+NmU3Im5NVUnfsmExDpH3qHSlu26lAOW4qIKaGXEMqG6p3qR/0EM6
wKD8qBRGS395n4PzynhehQ9hYLn9NwF8M27/n4ypJSZoJ//RUe0EFwWXtolT+1qG
Jt523yU0B2muSLRgUQf3QxP5FtU5ZPTP9Ax6ZgCU7hu0PMlf5fOK3xMEpV9aM2YE
UfOBa/5wGF1fZgkfTW/95iRhjsfOBAsYdJ9ohzgyC6aRxrTM+zluTIxB12+LXgTD
dyU+XDGDhm68Llno9DMVhaDg+sqZE9GJg4SMkdagcBionoKYc6FtCbNLwY46NMPw
KHWIUO66TGVwz8Q6pYa/mdErrH4KSJZ2Q8fkd2VnAU92FYU+xYki3ACB29NTchLe
3mjh9WJV7OrDciAlGvZPADeXA5wEDdlIbRkBgQKlzZUYSnVlAUz9JMva3QFSa2Va
bCmqwjQB6iHdyQ7lt6xWFe6mYXOqgz/i33YxYpTyUbkiw1iGfqrYT/YDu7sl2JK2
7ccn7d0EiHLU/jfNTf8gaR9jhUnISS/xHIZgOp1Nt4cwu+lmX95TvkGPRgJA+I2M
N+Tx1Xh2d8u0NTmgcNlzlec4462na8guKwjwjMHBzMNe8E3OetBb0GcCBF4h6Cso
oyaPuyQCMwa0Kwj/j7t8zg0/U6kmSmYW0I58kcnbtbG0N8oVE5IFkhcOOJs0oi/t
ziUz4XZLiB3ue10yg8KuFSJUQEbqmphlN4KFmfa8SOQaesrSRqmWAYdsC4wan5nP
qjog0vprZbHN2HDpv1Io2wJ3+dbyzndBtBTZTJNk3ovWTDsW1PT+zuDKESPnu71Z
gjjON5R+QDOLJ8MBNQlG64+jLmi/LBoY6NokzkVLQFq/Ewg1YqiTWHr0lNjvaKyH
W6rDDeXVSy5Ktl6gP2MzSqmT7xSf+i7JahABKXMyirJ0+09Ihs5tdufUmbNAPIY+
bvPpHh83vhprlWuM8X70NyHT4E+1Mpn9u5zpwRIqg6gskeKNb+079xOmVJXrJwXN
wRJ3abjWeop1jb0ade74cNOPJQR6u9TO40Vo4LF9BVWpP4wYmKiUn6CzZkXrsra5
o/AV034l0l5CvzPwT7HjZssT+CNAAziox91Zjo/oeJoJsi2qjyG0h+QLxVrTKXgE
DmA4k1f/JhIOBvWPdR2FC6n96yzAljNPNjhFETYKOMotdESYcSTl+EBhV2IXBw7W
9nO4P1pJjvQV/sqCxhXTmi0qwiybjA7/2ScEw5tjPeqHwvtO2yBt9uOLC8RC4OJx
1/5Q2dBESFyiJZoHvKZ0ZLOmqKT6ah+/amvDcr5HH1qLd3ZGNhMMS3p6hlDC43Sg
WlZVofA1UZ2R5X8XJdfs2y3HglpqL3Fw/9Z3SdXVqB/HCnkzA+EgEWqPWd3E7tx5
APprmTeAGGLmKgnM4ElCwhIBUf2gjjUqGrjep1o0TLWGvwfP3UR2Zjf7M7H0nR9o
3mbZ7+o3hul6GT8PosORni22lZMk/JiMCgoQfMEo/EtNf3fFdj5HwDIeHvrvsSJu
nLtbQkIG2Uf0R4ZDl+bTDjdz+AWK5+Aj7mt66u0TgQANT999fmAA++m4kMNx/EDc
7ETRIg0f4mQLNSvh7a7mR6ZbsJJl5hE3C+VF4HR8/zchV+y7mkhoI5GgMDQaaGwD
B/LYu0p8zK3/m9BKLU8WUXakd6DgFSzc2QgMHdA4Ui2qtTz3EI+p7C8VfspwxAFu
gPgKJmGZC2DIMl17JZ8yBNwcftltEeFakCcZHKgZ05tEm/cHkM69ST1rabws5drt
ZASq9zEBqn/orgf3oEyenG5WstwkALvU+1yhj1ktCaSZaVAc8deI2zAOXn60ugD8
lkBv3vm5g+NPxF8btu5zWR2/BBRXrIvvOoCM8eOfiNZJ8sNwFG7KyHrFbZ5jg1n6
ZKaEz5Se2/B4WBAa8xwfDdrbx3O9lul3Oy/m2Xv4fUFaFHA0MIvwMnXpiBD4YK/m
ikxV88H2aSAipXM42KB7CwxziLY0mtsnLHKueydsPBC38ZiZnN29ToIxRNa3c6KV
HPyuqVYB60Tpnpmm9IPoIOAJCpL7CEzT65/vBLs/+jPnd2Ix5rBdU8JlCfSW8Fu2
mBLQ2B2hrZuskNagdAODi46qRzzUuZK32GFI7AhFQ5ZwR4hAqCGC9Z+b9eYiYk7u
RPM6IF+lZwqoUxakzTB8HVJjVxgGUy2ODj/e9IaMRpSGLegqZyHLNVx93V97osOC
/+gUSdpc1BwouKh/bXZHyn/YYwF5DW3AoWmdWcIObnKIIcHWlH3iv0ncemKg1JY8
aXI+V+cP11gSJMQf7xBwWvYU9YI15NAgcvB9ijpoDE88BZtj0bmw/BHwVIBK3xcc
XZ/zOqM+LcqLnR3FW7TuPtK0YNJELycDf/7cBOM3RWyndFZhxuCsLLo8X9UYhNyX
5HS1WYVFZgJXqyk8eGxfTBTmdJwNUEI5hJ/6IGRcgkbgBTcGFtbEoE5y1fYJ2A5w
Vbqc9UVSCZNIonkB/OcCNJ3hfXVqv6qqxFE7UP84LQqvx4SQvx1YMEwVoee4tdCm
cnHcEiyPTOuZktUuxMGqkCkp4TTbEUuMK2AW9Ryc8ZPdP5BCYTH/yHpvkBB8yJqH
5eM3AjuBTOGF5/HJqnv0fb6oMUpBp+tB8aRY4y6+XPCROGTrs44LRcI4neZ7O9g9
eJyWZDUGxLW7wwTTu6XUnVyeZH7HV+jtc2dW957jUHY4dctFnaI5GBBzNXvDk807
oHjQSUENyBXj7l4fNWxSul/jPvwdnSMs6MinW8OrWSuOpiXEQNZ2DGyyB0QbzZB1
g/DaCOQpJn6oKme+iuA/x/aeRkZ8Gifg8TIFn48bnJ1OqPEQQfAd5et563DH9DpS
sYcZ8MKY8GjAqYYdVRIrP12C8xNkUd5Ky/aLmAGBwVHEXkhpL1utyAvvAVDYkiDc
mYr+BC0P7ix6kZv9uBPnhC1pV5SqbZGG7OUBKfnSkZFY8oCis0e0cXO1LLIY21JR
gNZA0NRCyYRkRKyRJjnscRJcw8S235s8Nk/hu1CzYIatwcCASsI0D2VFEgVpn18H
OCx/wzcp6y8AOQZS5ZMuysQtCAYyEYiVDYQeKtr4x8A2IOZWLKx3W5eia1U141dS
u2xJgxGUnPoX6f0kXmV3EFDtFjXrAySMr8Ce8Vr/Kv2uO3Cf654YNQowYKTnZ5YH
4HQm2/CJxkKfeYI/1hk3jl1an26WSB8cBKUfrCFN6y1kKdDo418h/CKcnwZ3NztO
KNu6Y43smSr5wh3J2B9ljnm0POR53CB7yaH+T2IN4PcFXqgCguGE8n/pnhoPy4/W
x36Dp/vR+PzA6zAvfTPdlVZjjLAA/ktWOiCTZGKEHv3qyWcGXwNx63QH/zakzX4G
145co48qLPhh0C3jpnd/J8aMXCZWr+ReXaOPYZUfzVstqy2dys96fZoiu0B6VoOU
dy9dllq5srZHjRzcjuzWjq+lbuGlCpEraJnjUjrRObdjgR+UM9Ari+HLCnjSaH1j
cr40u/6BTGoVN4nw1WlTqvBiAZgvhoSq7HQXmgUgFOS315k9PFbr43VBVxUbM5Ak
i8KHSEAg+6g+dBfFzcRqkjYxhk0J59PXhRgWQfmEYKpLw/NiXD0WklhAw48vTwNc
36Y1nLW8q08wukTdCErLPBqQiUCFA0+Im8JNP86BvMQ5j+gwjJVGOPzAUuxK9SnG
5DTdaN3ovVucih3J7kIAA/R7cMHbl4oXKm38etiofGVoFiq//p0vzrmHTSp9apjU
WgSZE+elvK31SxF5dw5xWFD0VaUpgqwTO+SdCOKdPtMZyZLk06nkQ9gXbC+FqiiA
MgUtkFJtq/zhaNYijD7izBSX8dnDKGD7G8LvAZxsSwkpDODM8XWtCuY5rNoDtsDT
4m3WM4A24xKw7Du8rWo3HtGZMIZY4Xl2nlJfiNSclNocBxvx/pCPGw+U0gsuEfRz
V9RIm6BeN0XMdFXst43o6hbbTA8z0b43i1979v5NAZ1XDpsoVR9zuGlGW/XBiXvu
yJTTytHsfF5xmuU/fXNsWeOBL0q5AqqaecsM7W1K+qldUDPsgqadvP+f9940taZP
5dFlnvPej/2taXBb9G87eAWvlNtPRYz4erUalmyOe/DcmelSYUb4vc4ZyZlCr6Ty
4K+w5g6NiGselRj3i/eZvsbmNHLED8/EbjQj5mq/E1y/djdOEQ3CXi32sWqRrryV
1iVnFCTmQKzrPvTF2U8B8Q3KH69unHSq1dXoeREOw8A+Iifsqd8Yn0ONcYxLSWnV
c1ORA7/a8kl/jp2ATRE7RHOgcyhV55/5bO+cz6IT8MBjF0r7kkUmKnNx7o7ffBn3
qKRiv2LHj281ADdt+GfmA/eSrCTTYHvJigyQAO3EDBYYnJ7p/DagYyLBfTFczRA0
oYeQG2bor51L3WYBWit7nLSXjlT0HS/a+vMyX0R9+ZIT4R7tUkYTk5L6+10qnsop
k9K1dKnj6Fwf8Y+TtCQ0n0fcGmZ3wTbH7cauDIQIru6tapyR4dhgkQp8X7OEiF0g
YAq/cqf150MRnN/UGa7hMcO4T/48snm8M8YF5ichpy2lWKI1qefgq+3t25oRDjYv
A4JfB4tZuK7jUnJVzhtZsgLidx7q8ou9xo58tBwzQpBWmwnVz/FInbTW/kw8K7zX
2P9MY5DWmKLI8POdNnc0LXUtnmBP1X0E9wBWnjNdwUA/969sD89NXrf/Qph99zyt
CR+4yXj/e0R07Uo8pucxuWtAGMP5nCcAroFQX3LWiVLyekc79B3kSb9Xo0kKYlKp
QdQkoqgA0YAVGyz3cDy3VZXRg4HjJdRVWocXMaPOC+YxcjCDCpDhfYGqrU0LixG2
ekRGrA4iGXKmVkB/aPEz8c/FTyHMy4M2xIHuisDaqB/vHDMnrgJfRbxJa19UzrBP
IrBhAmCOpDO2dKAI+RadV0Y36asWyOkp/iYXrzUkys5501etpYemnrvhaYjJtQ/Q
GbLiJlAKVgO5fGZpgOCTT/u2npom7YP4C4MVwK20A6LjJ28TGAt2XnlNN2E9ahoG
5YN2hCLKX90j97sPehis8diyvMD2/We+FjBHJmMM558UrqaiG/CM1F7PqF+ch5yM
qCM8cNbR1kFQ2PaLab6kLZ4W/M89mK9aslAclIr+Mum9iAO1aCaJAC21mJ1Ccwvz
xJGyCw5NlGBJ+Nrr9x/X7LhSVbjfwCZ92cGWeqMv3jBSTLmq0S5T8RHLHNhvsSfB
pLY1lyxlxPM0i9Cog1iW+eAFoWNQBIjplyP5jztZy7QzbUKkZeeniPu1/ZP11rFm
aL0Wgqz/P8sVREs1mxVpaQr8ioASMLe591bi4Ja2NI5C4FzwYRNOAPdqGe2EDr9a
FXOiRR5lA9zVa1NmdYOmXxL//JtWMerBPNWX3OoKN3mrNtDLblwF/UAhdV7fUzHr
BZ+HLLCFsyhyfRN5glovq7DXCBBX5vo4NYSmBlZarMYQKYbuRz414upk+q60UrYU
0xe9JAbteXhJ2c21PAuvLrNnvvKFJHv0YyeVpu5KkSrDRqrIb9jShIjgMjji+qJZ
+OcJ+nZZoA/Et7N1s1KmF5rSgrneX2gQBtgz4ZyZetB2tvKWSoOHb10hJqxhtNX/
W543UlylKc37hAonQhePbgbV0de0hqHO/U/n180RgjEdCWRYNntycKv08vf/BbMx
LAiYsMavME3JxU6QOyVr4gjYgI7yPevdVFsEPVr4lzH1FdHRvlw+10mhCGQ2JS04
dkpSIKFeNc7FEaj/OXZNOUSq++U9Pslnf9O5bnE8F6adGcBVg981oc9xTterRK0n
I79nM83ce9n3etnuRoXJ9KH49MUuGa2kW4bcykQIYAUmxfSwc61YT04aokwQ+c30
UK43tGoVxbK02GuffpKfCLOhGt0QwxS6SGpqRXKWhUP/m2M9Jmc1wmLrhObnLdNB
Wre/3vjqe10L6BJrcBMQDKHJAp/9beDp2BPaILccI64slZg2z1yqRqwNmhtub0We
303zn9HF+d0O4wg5yoDQ+UqevO/vexl057itbit3sltw8OKfnGGq2tGzcgHgKbDs
F6MLjHB2tug1M8JplGugLkOQs0oKErRKEacfMnlptbdk+poqCcsqmlCPd1TnXz8N
jtwP0oMQtWNFK0geyeIWeBexOA6/4aZ6gL+Z5Wyyc/LMOowjOiy+1VIdGhJ4nB4W
RugYhQ83P2w4VuYGUugZBJKYGyJgv6QEpEbOzE36q+jux2aVXgkYec9mPogjaU62
u1dTtUHIKPhzbbANIXEvb0A/Hj1wsLnFfjoZNfYFk3N5wjyioYHnqsbmp93aWkcx
ikpHJCrFLnYN2AISIZQOmUUapq7YhPT4QYdJJNg3FVSXE0oxFyd5UBulUL1jBl+h
mf0YtPJuq7uMLoFUa4gkRlWT3A+PrQanpvLYz06n6UeuPPjqu/53LuK7D0717/Iw
cQtkWpU/nLzoZFghYH5FZTrbgDJ9mGhKnduxncdCxtDucq34udXj4oceIKRd8Ths
DDhh+CnUR2JzSdamiM19IloM2sOs6/ReIujVCxvw9srf0w0c9xHIVcxnQHmKE3NN
tQEuMrfR1kJKC7fSYDCIkuPIESc1y2Mu9Gu0L6dblHmKG82ZhlJFEZYZofP/bkRe
jgwfUVfFdiEFoWs4JV7mHxNPJ13vsc9Em1y7uXKrrRPH7q+H3zsqP7O/ejSQ4frm
OYQesDOKjqUyuPeFVYMSp373s1vGIlrnzPOP2ysJrLotdbGF8ACIPXlkwnBrB8zr
GTyF6fjpqD9yeSzvYk3EGbz24qXW3FK8ecuqabuNPe3R52JYnSUId17QoG0fSIbR
gWVjvVbLIOVnBU/u9x/M1Q8J8Xi3VVYzNvVtZSgg3JBtbFkM64Y2n1Hkv/G/COiJ
amCp60J/K0tXBFwEK3ThN+r0Q5M/s397yNkyeu0Mjm1b9aSLov0yG2cVMqoyNnyj
RvIvcobNgfvTbF8VuFn6K9EKicZHWBt9l2IAR2j11lPjg8HFpuIS693ZoMqhhH0d
GfRD/5Oc7RFdUxpREFKUcDxiNi+fu2hrjELCK8uVrp8guGXDGF3FMKybGMyTENEK
AAGAUSW/V+gyVTECgoBlqpvmPYxakqc+Vot19GJU5A0RmN5qmDbaHrHkrBWbNa1n
aTEcm7G/hQ3hu2zgAIDVcVlGzF9d1UOQiMkiEHBnlgYZ3wJKvmLk1mFGIQfgqgr+
GZz6L/Ac+vmu8mOZaocSxnWb6oBWK7wSfW2NxqrthKpWS4KgFMhoIKv7asiACzCE
69vnTKvtAxUENHihq60VDsaui5MZQlyI3swfSFv+YdSEnk7h9epcF5hyDqkmB+Cg
OmFPSvDwFQoIORSVoX+59TFwQ94WiMI2zuyVMyg8Pvil/XSWZE6TXiDHHmcKO6Yg
doMqcpAo2tXDbLDc5t4kgQWJsUsnbABrnzjSTa7JGGbGOzwBneafP+ShRavhQco8
7hjGzK+W12VwWX+kOT65EVAGSt73ch2NzV+PAoZ8CBV6F9BvVVUMV5HwhV4jUbp4
hdK1YFwbwa05w41YQrK5cjMtLKX2MUz2xZFsKgGr8keuO+Tx2g40xrPQ4rpfU4Wr
lmtYuK3go2+21vObI7IQ05aZLyWMC6ryhnniVFCexIRgq58JpP+z7Z9DCfcqs/xZ
1Aw1ISAsHKeiWof0xbXf5z3j+gLTlu/OkFLFxED+mjOSJsDYpls2ZJqLbk1itz+5
6JQ7DIljmanDQS9A/0k2jnod12Uya0bGvwRzK6utknpuTP5z8N/H3P9/WY9pPQ7u
LCcXLJzlnhpFB+qPFeyo5HJzV7jqdAqzvYZwGAZ/DGbTAXC5l4zoB+wpKsvu6wuo
ozokavDwtHCa0Qe80wioLmHZvFziE1mWw8m9pRCaY7UrNEAGkS75HZkjAglbVJ5O
Y+l/1QgdN4jmlwcj+puNmnpH/qu8Z2KXis3Jgs9BqSXBr1e8Avl6ndJGvW0spA6w
z1rr/TmOcWj0n/F5TY1aEeqwy4ugXLLOO3bVBb6eQUH7kK0twcHtz0KgAe7wAXtg
nCqZtBGYp5AG/gfIFmAMxZMBwA7GWg0UZJgp7mU9zETsXG92lrOV3ZDj1lK5CMp4
s/d3RkujRQlt8KIg3LsIme38YycGKUIJ+6cTw8bB89PrHKM3G4skbhSSsnDYqhMO
zjXwYjT8WfOg2+A7nOo/Y3VZm6pVp3Qz83jH6zGH3uyYMxgDsBZdjcH+oIjnp5vi
wKwbX2qoO0efxjx+jgAXEGxOwYxHJCJPsPSmU3YPaYh4oGY0hRKt2GkFhDp/k/is
YVopU3KFGz1NcB01J6MGU33+UHFm9vfhlQh5LGUCjGfjhfNlOsbQ1ne8iGxYRFoK
Tkv5bA9lgRqJBgqfJbyaoyL1mVEdTP/gaCB3beFo3SJ+yCX8qGOn9hW6MWRb1x5T
sD+OkC+ehCeqvA8SrXjNHdNfy/+C1++ulg9m+XBTKmG6fW/9cow2cDeflbBEu1ip
OPbhOno23bY5dSF7M8lCO8s4Qm6kw1UDTHO4tps6hsg8wgsaod7Vbnu4+0b5AT1k
wDi/m/pgpltrAZI/K1jLnxIoQteHz6F5/X2nZrpgcfI/btErrS2A99Gu1bIckQBq
ujO6qZNZ9+DIAfgyXbB2CggVi5SdRGPul49uRDRPq2kunfRoTA0Fe6gvQb9hyM8J
KDYsCemj/GffzamjXEWkBX05lHfoHvTJau2Bbl69WN6zAF//Erq/ahc9UWbLxkGI
8CvSYhdv3mfM7lPfl5XJ2htH8pjSy/vr1rPn6llBZEL8ZemFDOUIMPpYe8yoV25V
rGpkoENfVFk7SX2EjunPa6a00YXd7SbO96pVB6jPCxn3npvYJqMKPQf9D1rJHET0
4e2laiIG3YxJNmWPm37u0RlqtlHCkrn9MuZ+oVJr7VmJ3kpP7J9e0FG/D97cnV16
ZhSsbb2n1zklHgzTHggk4QrtGhq8UY6dg8vhbNFmH18JGy4ovA2QG8OAt6I5QiXG
sUEsIRt8dFttXxnhlw+fRifo0tQi08BgIR+xx5ZziHC+SvmADx4x0BUyXfoac09k
5ZAuVgY/wqnGYDOhVOLMliAd82y3/A4yolx1BUrIODL2zSSK8Womxves+hD9vi9t
mGUU6/ZZjxekl+cs0hBc4DoTQgzHj7n80vUrFs8XOWGmRcnrzFQCu9aNCHepSrkF
6oGyXBRd52hkG3RqTiBOE4RY3H+UdiX8AQ3yGxDX/d++KrMTNMjLYJee8xWyUk+t
W58z6qOOrRu10y0WLtYE+lhm36WoIHxpa6vef7/5Uv4AJpPGxXlgz1tbR+Z/ViDw
+KM0DTDVPs9OpbQLixV6FV8fjzpRcHOL79/BgiY/ycyRM9ljki4GX5iszZeFfPUO
vjZdL8WHntbWGX3heOEEPzQQd+WZSjJkjb3TZ7KgmKWORVQDwOe7jEu3BbrdJpg6
tqCvfE1ZcMYMaStbdg3qVnbSPt1DtRRPs1Akgb0ZfVteFK46+M/6V/0q3+SofWOW
Si/u3JBhNtrnIcNaPQFtgrYYXLmNj/Fk9MNrw3DhwcBp5U+TFWf9/JvB3nAh30Yy
EKuf8alPbx8IB9l3pqdROW3Z2Zz8ko+jWjp8XBsRgYhA7yk3eeW1AUfYxxp4tb2g
O71Hm00Lszd93+TyP2K7G710iqlfPVrsdNdP7f2Fiud6MAGsnCns4D4bI9t4xs3I
Ntik5Ythbs2OyQRCBevuf1nQGo46ZSiR/sRGfbDAQLWRUbfxb2kFtpq6q6WZF2Nd
U7wy+AauhvSlNc9zNKakTBxpwfD9h+JAOfZCMqKr9WQjSHsdTMKNa6JnPOdZk0VC
ihvxY+P2PznJgNde2rUffDeU7rzAbJkNUtOnDR4ZmECo3dVFnQgxYhxRzms9oYpk
R+n918FekdsoN/jlaCnqhKCMKO7yjAY+ORnJCaf18WxQMYHHivfzIsthmJaYjYT6
tq6mRjRz71h2viONdlKQ1ld/lBe2DCwIBs7CaTrbuZ3tIAy2W/SGpbxjizTrn6To
mbQFhZfNm6yDcS6PNQhmAYTNmz/INQZ+ZFasKn9fk+lFYTEu7I1FN4Yf5P/5haYB
5VmjXCihQJ4t1UjNLkhxsySSMiwSggdO+25imZcwSZsN8QB9VDle4gSxcwl47agE
vMc/BYZfIsQsV0Wdra6tPX6k4N5TkQNQ0SxLr+fXCxDs0NAqEjludmN1MEFUMlXz
p3z/V8+APmvDgJLfhnQdxJnFmIse/dVWCoe0L6DVKb+AZVCIFs3eCyHuNg8+OFRh
cfe6gTQ2z2U+Go0WdZat3AVvJdIYeGiY/i/eXNHycbkLlP5zgSFqbqMoIsVAVNEK
qz7PZ91iCAnAcqzC44lX6yGzgvmgL8nlsWOvEDErCuKen4ylQn5uoJtL6PdKvkM7
cnVQdHo9yTqG9eK4PQBYabbCuu67mLE9gw3kZEwgbnlds8DgSubEx5IlMxk212gJ
/ZOMJ+7Epf7lRgBxfU3nmcBV3a997eldH3ZL4Xd3s+u3JQtY+EOvJ+apmWNqGDZc
9rw32M+p4SlBpuH2eyP3lj8UbZl7iwEbU1mZs/Og6Ppdo+9LKSq9sCumThL02l1/
yiywIzxWBlmr+hszs11sq8TvoZdFXnWQuMmYH9lSkyRLgjYbbse1uG20XJ4na9F3
QBKGMoh2dkYXqIO/XoBZ4oAjweGUlmjr348Q1I0wUX1yxfrgXvS572vCJGTHwTU2
7oVfUsJYbCr8ZydR84JciUf0ueHNyXrAA7dytGija16GpeFrNmzrvbK/N+5FdPCC
uRNU2MOPP50uAMYYhaUfukAmQIKt9j6JpB/XJroWLEPgo/ytpGU3h0TSIG+9GwZi
q+Yzd6436LFgFah5J7bWmXdLzQi3cqEaO2L90oq7I1CvvwD9Gmk96maHOcbvyUe6
EV+2dYMYKrQaFAhl/5kduRhIZNpnYIQtpw0u3/oEYmJUc/XB6b/xiZ8HRIRWbgCX
SIrHdK0JXh4VZBYrbRii51TAMk2D8AcFtZwEdOCnOBDCADsDgvMq+GoADP42nw2G
s/P6h2bGC6Er0EFAiNwfHe/ZaqQLzmg8+X20g76Nluts2c4aeq5MLm+zaN3W7aRx
yPSHLfo/1r1y5pTwl6EjFooUhV4odh4qTgNb5uCobt+wviUxb9BjZyr1QATlJZ7I
5F2G271p598rQJSbFNPVCVoRufJwU52BOvwj1Vp+n0rY7MFZh718MtCLgNbBWQ8g
LI7bdOZDMG37VbJns3oYXKKSoo2dRD4PlM6syDA1jDW2+6Y1xK8eHqMvK//CY34i
DxyrmmqKGXXU7NMGWf8xdS2VHsBPeVLWXRn1GpTKkBwj24CNwVZf5/hKMj64xKqG
MDhMXXyoKK+8CVpyjFIjUmJO/Z/gErbXAOou8j4dAzA//QUOo+EUXJY+MCO1RdFX
9RjX+DwT0vH/QZZlP+AGizzdWAqIPHFH/B2UyD+n7rKwabSLewLLGwzI/zvn1WrE
/uyslj1VU5lS2EuhnUa2F7+QmC/nK007xYc2Dq2uLUhACCLbT0kvQDHukwhY8hEt
MKoicH6ygMJ4Tg+VBdQxt04cVW+jr712cW3ex2L4rVBZS/8JZpS66qFvmPzjbf5m
eb8GWE81/nuSZErRnzaMTxzt65OI8HGOXlJPKesDXqSK+zIhSml+84UZEupGUFKh
SWuuiEZ0ooeJHMZ1A7pAulF0YELEBY4fo0NVmJqVXxS1FiOD0GUJBUJLssJQNPHQ
+l2sYcPa7rm1SMfzvm3wLHtoNFSS2YciGiB6FBNc2u1K2qy9+1Jx/PawwTMSDrU5
p7EuXs1ruVKQ7UmFspJiP6/5v6W05eTpZapGyOUbFl7G+8/RFiTmHss8+0ILmYvE
bSA6r/2YkIfoAPj/DJzuptfBlAoErGeLjc6Gpv55RzPqZF90zd/W4LUAeKpApHDo
thD+bFT5XiPLQalsP66D1B8gs5EKKkx4iw8rhGiuitmR07amvducJ66UKBuD2sar
Mncd3vCj1U2bmKDL7qr14xbH/uL3Up8APs0+toYrqVSdAciJ+UVqxvVR4QZucMTD
0K7tsxrty6sj4sjoGNKYrFc/n0l3mzMjrqNUlJnu1jyeLKg39B0tXfUHLLqPqQ49
clVMr55UI8gLj1rFpF+j5xC/cUT1zFUsjQa9XttyBjpHFRtYj4wCi8YBeYO+7FMh
CAxndKeuZWmT+TV03nUVuVkxXoV9eXajTJ3LFyRRRsO1HGlILY30IPX/WqzQVBzA
U9YebUn1hdL/kXWiZoMTEXd+JbP/rw6Vsv6yh57E2MCYV8V5uWCDSXsFRIuVvg0x
fqjOQbfd37LgLSWahxKfbNYWSeEAFZh6FSc+olN9qgZLAdMtIFgW7YScL//nqF3o
pH1lRV7bHNc//uNqaJjxXgA9PCYY11I59INyMCgxAl5ylK8maOipxO2v41J+ww9/
2Tg/lc+4aTixxGhdICqt6Zi1GdSwW4ZygSGI76GBQhxU2McNNCZuGCi0seT6pYAt
cCa1hXFpu1/dhdXySd8n+Eg0tnZB25PV1Truw+PIMFPD7x4haYBEo6xjViWNqP0e
NF2ZlojtvMfMA+AmO+FrZt8toE0Z18HiUkLQxLIRmMzQts7h6fAQNvRI1PMSjvxI
cxfR8M8C8nuQYwAIwpMl3d0hm/3Md7w79arGTX9BYGSccfIauKff6dQwun+bcfVx
rDKxRw3Vd38Mceho8L0u3HxnfPemcDkQAE6jeow13TBDWDfeKvAO44ptaUUoPOpJ
ig+zJQU6BtSamhDVOiTD9R2m+yY0Qt0ODo7fdwxZ0/c6GRBIszl5sdxugbE7sE71
3Ua+P9WiQNxK8j8tyfliMKrgzhDBY8RUhsueRNav34MNVk6MhBcFtwZ8pmK2JMAo
l5A2DAcb/l0wVSvClTyBndpejOxVPAJJztNmxyI/SbHQaEgmf1Bd2kmAgIebSdub
PvWliYiZ7oiRF1lZ0j2yU8chQT9uBeBslKwveuJd4BsZu79b3pHLxp/n2MpqvW8l
BsXoBJhLrkk88KDUW0znNi+VIL93sG9pa/MEQt4qq1nmobYkM9i8D4LBw6OWnstw
3TQMD9xwOdHsllSIXP7wlh2U1TZJCnu+Asp06wJWr7vANWHz5z/Esp9x8+uwVPiR
464yubvgPy2PmU56sMVd4tXZiPw91LqVIDXyLBPvkXoUsi3MZ8euwgGmvXpsRCuG
Qkxl5ZJ2tdTFCq385CxySjdvsJ4A7IaJBBN4BCmZLiH9tcoXd2jYJinIbShMXTDG
HR59zuVvtO1kjZ338TWsZ53CHChkTiHt4iebhPSPBHGzORR/lckwqX0p9XUemEAR
bMdwkUc/3v5gM8KVIuZrU9oU22Pngn36DjmYFdNk2wr3Yeoh4gWFkL/gfHFXDtvN
kHdL+A+R/7O7KtbRp18P16nmqDJF1HMPbIVt3tLoHF+N5aLpQxIOrciuqaUgvt1c
+7mx8zHIt4fQEgJEzE4+eWh8bj8T4HMv0YvR3dckVpG0+FQrehY8SnNwEipNo4fq
ctgWNY52Gw5rgSYFCuTp/qEbAMDdSS5qR8yKaGVqpbeEqCSqwvB+U66NIDW+THIU
Gxhuv3iuiE0x9/kfX43Dds0GW+OvKsJ9mb+nODkZmvnlKRhzwlXKCkK2A807ol+x
UeA6vz6XMPpbhl5MBQUTXWYi37/tUmNfZEc6gdukzld0lO0TmM2PTkq5n4sCZzSI
Ce54ZcUPccLHiIWsV+W4a7SLsccv1qf0IQpps6RpLVhdKIzjt7hCDJxlxQWkZRkf
epf5XepRCHbmk9BjqY0lUOBLsBpWhO3WA5dovNTyWgN77SwANw08xFihhdbfbXJU
6wVnl7VcPKX0zXdVuQ+zLiDFAFpqpU5oRI/bhBeft//KL7uiTzEpGK5sVN6UF8Sh
uJqTRlk3TLHlZNQWxBXJW9C1rDXqtajsBApKCQeWqRXjBvIhEjkPnPID4NK2tyum
bHRUwmVTrs5d9vxABtssrsaulaX2KrV8wMBt0FFqSdYhZQk3vN+WM78ocJZXUNXV
+d6tj7wiWjXUpnbhKYRA4QkhUsjAVU+ZdmlC2Ajsm5QhFd8zPEszt22kTw2xrlAx
6f4HqLDZsR7ZHx29KiX/oIskXDcjN6Ffgayqg9pUQKsWBhqBiflVTAelUjZU4c41
di+H5oKptKHQjbohYP6YzON416g4JRfcpQdpnvSmPrY9j+tkld7pcx2zWGslnaGQ
ooi+SGxC6chSKG3WAK5y8b0m0GwuewZ/TVEm89rr19DHkjD1vNshaldaaX7jN5zg
GKgl9yhru2GUVnzwJc6KPJObpSqc2t2VQmGkuTRB8UhVJ1PrEVmzmrhhE+Y5vRRe
OLt9LNoZKbhTaA/0pYlpW6+W6FpRi3BPDCR9ubSKM87z3i25vBqCpyJuWLGksM4V
8pYIhxc++9uAxHSq8PNjzeVjcEhH0uRcDCN31ygjEhbQFLe7rdBVsBqk1gaD4OKg
iQTPDkApEySG4qCCESAYsJH1SJKUWyJcxbKSui2sicqVyFcd+6f1+nIYVtEbrR15
mqm6Hh5swiMoyYygbktmBZWwHhaaHloH5CXWlfGmORCBSEFB6Cqpv4rQnDCp2VUd
ansxsSzDD9zUSTjDQC4SgWCBir4ssjk708gHVRBHB2sYlOunCYSp8OVEBnefIWdS
sR3FOTW0kKmoG6bZXG+6uTzDf0RuTtBijOPZ6gSGnVHtvQ9gGPB24jxP7jWaV515
gw+ZVzcxNxPHl823jCOIERDvfmpJdTMlfrg7Dgoudv9SQkGNvs5QFrxhduTLNPh7
oX+i4+/tv9Tu3/Xu2hx+mlYzqg+aXmiFVjytPX3k0+FaVeFB9bGVDLAj2OxJ79wE
yPr0/jlqK+3NnAbggx1BN9j3QnMtdfkMSbj+K2Ef97Q++5MQY8PmYe2CHNBi5dx+
Mjw9I/mS7GvY3ByHQqbG92yRui1V+A0RA0C60AlKOJ08+nN1Fz3Esj8dcFT6VbZU
7Df8Cq6k5EA3ugPAyE/yR+/OqWSaXtL99LJyc5T2Bu5YHRy53ZAQe18TAugsk7NM
KUM4PDZQquc4RP9Eqjl5SH+1GRtMvR2oJdXJ2XTNgkaUUQQTDODUzrVW+bkFlBxq
imnhZbtraiWpIn7Ak3ILIJPyQxncGkr49HYE1JBpcp2EQtT4o4HJWu9b202u2xPh
MCKZ8BY8UJBaxW5R6uPV+5GTLSqSrfPQSGo29HRUIrallbXy/DRh1lLaf3WJbYLk
/if8csha1m0NEX0tqSzRY82bQ3NDSZUDowCcSkiWvW7RgihYnVONzzsbkvJ0q++n
jwv+jmHFhTjdX0FZoWGHZTav3KsuNCk9I9rYFiCaX0hRXf49DNFtej0x2dQ8iCvv
HoOAl8sX8E8vTUmBmLJpbbyMytyRytD291tahA6hfvBDNkaqBfTAxdsIWMChU4P8
MYBNjoXxmHfajRl2IKCFnddoteve81rfRJ3ktOYGtuDoyRzsN5CGa4d3VwaNNMjQ
deQoaQwQ1rllfOpZ6uW+GvGDdU+3ffPPCumzUJlSx+Q55yL0DA7/7zZIoVrwEvp8
+mQw+QM4nSD4RvHQ3ASzLD63igyGYRu+U9iMRb8clUOJGx2NXFA5jGTaf4kKwVgF
FmCqp2V+fFmI/bHYNjFZN4QEoujTg5/HwRoJhh49STr8rQDmR6wm9o7RfqK53BPR
9Z22cl/xchapVhMvjG/EvDqJRVnIzH8y6SrBFyda2H+BFLIyYwPdeyc63ie8h5qb
Scj5Jht1whhH3VMBx80SZBRFzvaIm1Znwy+tqSErRHk250i9T39A+pW0TFYekhkA
k9IEcSD1nU5SJgrcH6sdITj7xsskaEkP3bM0VuVi5Hbtx3iUtmHxJ/MkTZdS7ay0
k/EONPcjY19PotRDV/IKSNkKqwAsF1xl+JxCHLGc1MWAHs4e8gI5nbjaEABiwAc4
7s3/PxXsjwF8VqknUJPfdKDfVRGc+u+l5bIlFAATP6H77ihp3262vUUBq9qP87sQ
i3BPc6Kx3+curFjYTAlTk82cBm1wzWXrXcDcdg4hx3X69HW8kpQPY8Kj9/lIed1o
4yKHmQXbMZ61JHWfOQpYo7gPkyF8wDf7pIIMqFKjrGUXOO6heepiRPFy0S3L36q+
fqWyhCM6CupID2kjAd7SmxPxo5sWbS4RX3EOkk4TaN3UPkHtVAjsRKyJ68GNk1iv
PAeY77RMh56YnKTqlz5Psh+/ZXnq48V3b6WfZhviScl7xgTNKq6N39XzURr6W+jq
0rqTgT+oVORVeMxLjq+2f9hz3EGvWCsmmBG5XntJD7Zx2XkZ56kTiUcDIbdKzYvW
NLiC5QSD25AudCBicpHmnXtxIpj1Mexlju/GesfaD9M+3a0Gdp2Zsn1DrlC2jMug
EZz6gLWxhCMNGrun+6ZMy/FmY+tIA60TxDwjNOehaHHAQfIf2HEIR5cFnhNmjHUx
BTdgiHTJQR23ivCpRssANMVQymT+FvBXcO+GmNYAybTZAcUJutCPU5027aNmOcFZ
TnWtr/MBbwzi48o/TOGjbK9/Xd7RKKnsyrhAe6JTLyL07re4e1rOTRi0vTV0sItU
ojENR/sEa9Yy2ueZhgKEsqzTY9UJV5i7gZOjK0jeZ746XVDTyv743TxglHY0Lj7Q
9mPlAAhMgBJrpzFbbBk1ZxoB865xx9pDzO22yXcmoFhwm06xaj38C9AuM7VxLUCJ
9HwKUbW0hCxuUJJFp1PPdGixl5OnzuhrZpzMWgcs6I8ySwgTjLhzRYjS1gYydMjF
8WN/HjcPd6aICkkmC0WnNyRMpKz1IAwMJMKZMmSvqFMWWTNVJJiXaLPEPM3lqIsA
NpXs5b8UY5ltDvU1mV8k8QaozJQGdYl1oIt5rppBr2wFJEukwvuxLIg/bQEnH5rZ
VsHtsO0swu3m7eWcu29gdbssEjn26YNT0Y/E3jgIyqRWH8OJTjzC//YiGxhSZvkG
vf7QzsJFXO/tVbsWBjK4f+i4T4125+mhdE4qRcjip7ot+4mh0HTg6egbg/Ucf8Es
D3SNV5F2ZcrQX/xHmdAxvPLhVO4JCDIshAOeci2v/w4v24bhjPg2JxAVgTG4p3FA
MwzfVgGMCbw5pvJ6dmlRBGtjYP6XAqNLlMa9wRwU6uFG3D1QNAkJMqRighRw/DUJ
vq8fOfEZ4G7wLwxedNnqeRpatTguyoE7s/Ja/SyEfzl2LqOaMsn+I3i5p+6sk+5W
sU4sg4XnfmzMCZzinrZrRl33cj6XZsxYVfoKpU4/hwcUj73M3pEnnGSi6SGXhP4/
QfGV/rWR/3ZUIH21huViWvbqj/LuKP5x0y234OuAOsQ98yy20baA0oc/XqyGqFVd
baEywwNKVIQuh98ZG1vuibMGIy0SkEV62gMGpZuMe7LZLLwFODGyCaoDj7PH4KiI
lLCVAvcSTC4H7sVM/jaNjku1dZOnUZRQyVAH4v9j7IZQncBUSZC4PbbluTM+Zxod
daFLZmO4gh2ynzN4FBG0hT05K7dsQi2gMYc+5jRo4ACGrTGKD5q3h/VGhHDhD4wy
8Fwnu482xQpJ38RRyE6zYVSK46iJ1WOcQN4kz13fiSWDrejnKsr2GaN9QycCTSw2
r+n8OsKRVEX0CyLTk7hgq8NhCJ0sHKBfrmOJy+rqYygJPILq0zrjZCkNgtESAyvq
2KQwZNpeYdDH85RrXBzFwVnPYYH4OBBYiP82ES23OY0XiQES4p7Rq3mAkAutn02q
ZeXycvaUJKQamh+Yxx/78bbxmN2JszEXa1UvUZ0I1XmKGiJW1M7XV1Gp2xzE6g6Y
eXJ7luto26H/zXvaah67xXNDZO2PWqy9CvotchiCuiinn4t3BiOUrcGPMmiie4Yw
k4hS9qXg3YI1wZ9D9DLkNaSNiUHrltTd/n31ZZmfT8v3rkq5DRw/Zz058KVGB+Br
8lzqtC0PrbMom/vsOpYP3n92+jM6ugjm96tgPZWfN8CYLHGH1Vibf1pTgcV+0g+d
w3HMh3UOvPww9ILmtaRBEq1Txx8pA9fhsttJlTCtKnxgQIkByzgGM7TBAKojCGtV
Qanrh7/rOr3wrSSil2D6tnhpSISy9c4coOp+dCC5Th8NzaLjYx/TkgEMZTftyKot
tYQOEfNwpq0C64uj4aP2WjDkTlyj5oePzNk3CDY7jYDDf29Ye7OFzy+NVMVd5Okb
jwTXv2kOHwqTxGvyA+vC63sCsLzQXZhWLgNO/auIMCHY78busdcT8BjmgpZQxv+O
Yu149vPbwpN1CQZzleoWqEietYROT8LKcrtQB27FaSHx1bJHoIK/5tGhcpMILYgM
v0+rONV+tE5GHaB7fGx3FGpC6ECC7Y+3BJ3Wee/3xauNl1M16MeKV0Vt9ZIaKe1f
fMOl8xVavPoMLvr909dR8sP8gr6sGB+5k33C9wz1T8264KEzB+cGLLFsuc9dyMjo
nWShxnfyK5IOCVSXJLmPC0yN4+cpxB6wk9Ezh4Fj66Xp14ieWHDBGALeOk8BAiiL
RNo2dNO6iR8NHP9NqdkD4GSStUua+y480eaAYM7XPVAh0iLEPTo3hVUQgnb/QBPE
+S5tUEk0BCZwqdNXQOKRUdCDGtZ6ne8bWQvKQ0EvmWd5o1KLc4rxHIQ/8JCxSwWj
4/fhnHXmx84VPXF4lIfWwotlnWLzUUwfC+Qjz9CbLwxyfraxDbnbQs88+3Vp3Jt3
2CFyl2p6drAvbn7WKjqVdPiJAvYk1CSPu1SZ19aTTpVIuLgmcmg8Als9bZYnkvrf
g0L8K+quk7SgYdNld+LN/gxUcchIaGNc28INB+xGL+kBns5c8zX6JvvPWZi1zyto
W3Vgcs/vHqeaiNlE1J3ExOrxm3ESNdew05DMdgH+0pTJtyNsNpdArQjhCimxZiVa
mbVhb8jA6KuwypniUwzxWO4tTcSbbuUE65z4TG7MlNtHdiXS5UOiGKCxTzT0QPeK
dXUR3D3RyuDGZp24yGZHoR3GQGMS1zHKNnXriLsP35LEXaxOlSz8V1m2FOSfuxNU
nqmjgDK+p970mSihh+1VzmMn12Xvk5EE0VvRqhZ6Gcz2Thocrx9FbDHLVLiSqoG9
tGTtZdCr49Q00m7j5/wW6s1meCGYBdd1etYKMpkjzyplWSycWUMasL22qsjclDc2
kgXMiolBFEUnHN/VWgC9/7CTplU8GS8tRTUpZ8chwYX0eB0ukt+CLYOrnT4L2FWg
NgsYDliSpwa+EUcdhZUC+2m3jELnk/BmTZmnmLFDVeSmuTHO1hNycxekZ0SkAw5P
zjYCKlb3E3jLZZUlr6OdyyWKCXrwEqA3t0ELcqkVF3jGKpfDL83qQTk0TKXtmktl
HXTq4hCEO0EisKiwBKeafOZlw9u+v4X/dkFz0RxyFf8G8fG6qSZ51pSRiNXjM3mw
uTnc22QNkM21/Sw/21SXVBAM2juEvKIGmkZoKxMWFg3vnFE8aydcqVLW3j1LZ660
03IBtE6895jkLGqT+T2CkAOEcREBBoM97dMTRBo9enx1HhpPFUJrlM27UAR83atp
KRuPtGgywKE1gd7EwlseRR3OVt+VO/jnhakIPQ+Zh9JfKfo5jB4qse0THA2TC27E
Cb0H+PiWhlw7XOqYN0t5uDCTF4esxjIxcEiP+FTwE5BI4RHZ6mhTcxJwmqytsbCv
TgI2VYQ9zrQtr2yxM9cbmANtJ2VaMCJ4yLZ4imIrvinLY6C4IF72cST6wsfXcvy6
659xorCtWt9kIFXhQRX34prQO6nCu1AIavhB2VFMPgeQW6Nevjv11WHKJyBEN1kA
qroaeY5/Em+/M8atIav+FCairvvYYihxieIxNcrxOjTAeYI/LiU8npuRbJ5/mAsm
UhM3nhGgkslv5PrldPpBK2dxbFw2or2NuZnnr0kmjmCzg4cg0ifMesFj0a/567Il
mDhB50oOC1G15IO35kTYb+yWkO8r4ATxPz7QZ324NJ+QJWatEp1TgthC/uvifL2s
KLy4yaZlrVn5VhHZ6kSY1P2i7hTojb2jyU0ywkxArhhdRtXfnjRV2k4BjrNA0LK2
Td+wnGc24YhK+qz9Ee1l9WQ44OB5obisNvGZC57wCkIRv8/gZ2Du1ktMqj2RQnRe
pm834eZ3uQDA9kNgrLLxSxNcOoqlw350TFc+67qmW5Yc2IEg4zPZLRABYkmvReux
qZq+H+dcg2lQi1dJ/lKkcOR5HTgH67h1THoRXQR3JQ9SBoNDBIR5GpOwM3Ayyj3g
TUca9UcwyxSil0zoTSCkIqQY2xIJ4ggcAOhz84PYvQUYzEqo/2/1qnUSIdVlvbaJ
H/P+R319oz5/P8ntEW223MFcGMh46Q//qYY4PRg1bboRxbQj8o6b+Q+iaGm8EfWH
Lcv+vhf7NqUIR2hhedzN4WovkBsZZ/51H0bTKRFn/gxel30jULzJ5en/kfZ8Nncm
myEcELINUBbBKmU+r7qb92wA+GSqgD6zXs6UUeGrw4un2/XFqqEdJkGlYAoXbAEe
inENYkX6DdieAda/jQvV9vtZE6X+Sax2jcGkUH7fTVNFC/yQSLbM3FW9O0Bj+mod
g4I94EQklvKc9e8cwbE4ByGWa/diT25mUs+ejAONQNfLfEX7X7/t6dY9mLa0pzxw
8pWhOV+AyOLmeVY+M4zfBIhsaCQW2lFqI+/Hj9iDKu1KmU5wDkBzn1wWVBmSytNq
PUl8Jw5k2lr50DQef1HMRtSDma8n6i8FF+TZt5/Ni5MX/cpc665G9+9IGnkvKqpo
dZ+TNHL/gAC0TO+L5M1ooFzXZDp4rivErqkHfYNZ2aA9gkPZDGuR2MjgRweZ72rH
SQz4ZdxW3SS9iHupVuvfg5foyFQOLYtOSjwhCjWyJZnUC5SwthUXR2lQjFjYcvo/
Nh90wBGpdC30PO5QoyntaqybT6QKbHMWqE+pPIAUFVAmmmsJWe8v50raVGrN97AM
dHGO1J8AihsTHCxFLxVLQG0n/5+sPCQYnWQYNrXQdVdzmYyke81MKEAm5SLcQjUE
wKQM1PXhMfWoYTccJu/JGbjzEE7ngB2j7PdkqXw3e3YCdRIxzOOzRhqf4StEHoX9
2PfCVbbrWUd0cMTmzWwWF6hlYwAokyjuV3/rTnDVmOcwAG+dex8g2jQSnUWOzMJy
955tETiLmD39dkox7GnySoH7M7GlaMb8K3Uy9v4iCEOcaPdywP053oVHrYcC190r
2GyTdms2VamXqzYPO/6eq3OUzRph2Qz6cSnG1/chSC7rhSzZwO0qFjHd9CcO+M5N
Vl4H4Czcl6YBOw6ywGbh1xs4sMLsuw56PrPBzFfagQ7Yr9oInGC6gWwQ2Tpevias
f+gJSzLkdVtpdeZ6JeCn1d/NqEeDRsgooWmDpZiC8BGAgCohcxYiOE635skYzgCK
5zbO+/RJguvKOLM08q5oiQdeF+OPShxGY+m3lLJE5lKI6urdrwv7GiRxhoCJrIeF
frWIto4nVwjFZ+Vm2spXydZ0ibjHdytg7w6U9Xjm0fIdydFdnc6Wl/20tpT7vhhR
n2xOJ+OCQkYsrlxktnmh2NEZ60GIrxzJp1/Dk3ctam2ncJTGNj1ppekJEH+o3B1+
N/TdUmudaBfJqEP3gvEUek26wTrEbWPgBXL/J3i8aMd4GMoPCUY2pSnjl7MCHBzb
s4eEZ49UPSEOzvqTlrJ+/IN8n+TGwS/fapDpBnLh/fbvWxXD5MhaynEVn8ZBHHy5
+RLjrjB95Q+KGjBhOeDw4RruTkqxfA0uV/rgZVVBdX7ydE6UQNqWHO+Uji7wDNcg
ODSLq2CWH5V+FX3qK6DA9mFmGWI3C+KMmjrL/xXjSyO/exl3+YjyG9HMESpJJ8Mk
bfYhhhGEPPcJHqRuHznvsh6fQIyZUpGaxkbCFWORU36tjcoc8RX95/ZpmPuh89Pd
CJvYo//OK8+B421XaJYkkm5TTG1i0iWgvYDeOF/6XMVZxjXuEgl1dH6XXWt6ksnt
r4YJgBYNh1juF0Opy9uaOrkh1h/oW4TAuae/XiZDyll0usjxjbD1gWcwdo1rKz6C
YvAYLkQ02Lyiy0j+ZPUxMa4BVFcOZdU1m/+XPlf5sGpo/lI9U0PIAeESMCB7muP2
99qnUkjhTk9G68sBfQE+UP4ukDZFfvoeTTMIHovFvy9Cz3LKAtWzP9my7EKGluBd
y8qSV6iiqZ+25tX684AvIxoXPxTDWlsvt59H3VNVqxNyFNPNz+nM2BTmn/uBN2iv
CS1OQzTsGtAPptCG6hKA+gXL9DD5Gc0oELQCkjopyAvbfXP7kPbZLcWoYR5EV6YJ
D/RPAVaBqCxVDOvCKJzLHDB9MsOw05ozRhWXk6cwqaiE5QB5L/dC2Gqqyqwxx+ka
15vi2gfzohxCmUu+Ys/CfQeBRc4sq6VY6hE02JC0pSDcPAmgDyI4PzWz+kvrltaS
LblmSVk1BgVrSlzJjF8D0rRowBxe7gXHwZwTRQCBYHR/57Cu6q9JmlC8jhIwXhAv
obapr+j0HVe40QI/SPzSSQ2Lzor14LAGKwj9G3+/5Edxj9txW+NtLqLOVFf+/Q4i
81HGf/N+9KZXQo+sNgeJ74ztwirf4km5pPq0LA8XrfcGP3NxUEmTlDGIqfKDZI+S
iEFKSz7hFzATuU8fdLOYErLzLX7rbQCyBSB/GqXQQHtmhkYdI+Df10pH7kfpe1gc
dQrF2VBiSeukxC1kaYw5GSdpWS7IN0ic9I1pNUk7+FUeaIFqIuDwMkWjYsPQnPv3
o87gxdsXYVIpzYj3Xoil3Nd7ejlOg1Bu/V88fZnmAeApC0Nhp0Btd+jlJ9+Ic/eK
eUEKgt+KTSRvNrzsAGEufpBJG2CiFDpknWC3rOIdmTQqMZG+8PIPAoEzbhAl4N4c
8CCHacGDsTtI+lfCCwD1srEFDAEumwI64BTa2G0JTjTS7qq1EL+PfMbAVPR8tYaJ
nreN8rEJLrTk2pYKPun3QVLbJxrI9ctm7vmV3CQRVD+vxazF/+cRtKYMQ5OhA3MH
sgRiwI5dCZm3wJmRjqOXCm7Mgx772oFjlpKXXjIEw2WZ1X2qsweNrtJQ2wrAe9Kv
ONLPeuh5Gg+UgSp07xp4olc8APdEQUL2JZL/vv3MVv8ASCTeH5yoe5PySKKckNCU
vrmFNW3tl7YjCxj5d/oKSMRhiqA+4ycwAnTu80XtMqB0AR+6OlD6Xzta0+wZHDiU
vX/prjzHSJQJ9u4CCzWqPVxyhY9w36R7pBgGy5zZPNad+s5W3qhtUnnArKGRRUbg
kMJmffoXJ07HkyXK2Y4b8LnmGXa72drCTE+WlmNdz3AaKlLJD6co91vtaDnpCZ9r
ZBaEm+wc1r5kTcX7Sbta8RAI534iZyqPKX+zvwZuaY/uXncnnnjHME9CN+Y1Gq8l
EYi9j4Rg9eTC2bTR+zY1ojz6SLOZAPdlmDEC/G6RokDPBvzS+sVEKI2Fv0KszfkR
HAVcvRKts5I+SyK+QUYyAd8anpCvRYFlpsdBaECGHCPAiI4OMmecJbGdcXX6Rn6F
T8Xdi9nsGl7QiRLKlnkQfUUW2g6lmlF6ZlNVoFPGsy3L8KptnIczvrYWYd+m3YsC
nPxnIi7jdQdYHC2dQN9imMcu5d9KIDd3lgOa/GO7EiH6OxJAMfIHuGIMY49hObXB
N14fN5PW6qV+ClneYcWqJLI698T7+FU7F1CqmOy9dHcGhZxtmEVoz84IsE7yPFWq
2zAM/XMK5dBXxPDlkzD3W77Ye6FtoJMoEM03ZN5VI+2FzCu9APWz8ElwL3tssP+T
TJlzcFU7739juVmxXsLXRGyVZ1SkNtBgDrSIdNYon12T2mg4DW0abHX23ry4epIO
KffVKcUxvyvk9KVqaFuh+8GHoeBHZYxuBAl7EMbE7WUWLF5yVlXicnf37ImDsV68
kWicyvt938bq3I7PJfmXmKnRtJmaJw8pWQ+QEGjy68vKWXfHrJd5D/EGSmEIKu93
OKi91NfKXz9nBbGiXGXhdY+tE41pXIFhFT4wnPDD3YsNeh018cb1v+H1fOI1NM+Q
9bgfIesgDGOUOfbE7M38UNMOQgHPzgiKbyIl5mw2BnAcjFSNMPxwdOcp2dQS1Rs1
JZyTq223P9BkTpNwrWv5/2Nixl3ytrVKPpmOykFECD/oZcjIiQCM/B07KajrnuCU
ehwWryO7mihh2BS1YfmQfXzk2cy/MQh1tsfCsiu2BjQhU0XSwBM2HWD6Cvv3GhrQ
3+hFgYGQIVXmVywXpodaqcYrOIVEE2LQUw9PuA/IuWjcsZV6o/4v+wGtDo6F3jvz
IwGFZLZsEXocfCn1UJ5OPeA/mKV2gvoaMzQgRiYcE21vjzbdDk55pWHqh9+928k8
xbrvLTVyiBXGK0oE0UMNIxKUvmJcPpFjDTHj+Qlv77saZNkxQxUsednI+spFy2rM
wJUxue+eGgSDSPib+OSqcfLrnZqANAXceNKfgUAV6QydecetrcYLtFECbVfSbgLZ
8WliMRC0NaWc5j1M0u4LranHAKSQqB2XxkUCkoRqg7mFL1BQ32GB2kPJrVbZqV0d
Y9+LIyWuBf9q5jV6FZqBXbG4lhckWSIrRMxDLqqcAQZSxDnWCLzo9kdBt44dssR5
RFndgVdBy3YfybR8QPOSUb0hvkWR09hYDt01VByEzIYFPqxRnn7Bm7ZyZMk4eqp7
9sRFKkw4G5edPgqtTlvlflwTyQh97zZsAp2bXS2aFb70/d3AoTipSAJ2OQM+POah
vYMR2ljVh9ty6aoXJkIbyloP+F1ozxqGlOPN2FravdGvQy7K8wPoAQlsQ43EMTgg
1bt1mmsOQZiWGVQBkquvifeOQg0s3BuTfC3uUiGgRWlBDTDCyWCWpXOpMiKPHk0F
yc2/l4H3vZFh9Iq9a5uOWmacs/NbumSQIAkon+S+tQvUzAdG7t2FXX/5GNoPuKu8
rZEQX2gwA0tgWCY70mfoVE4clgMCPZ9HOSoFnwnEGBN76ticzAlyH8g59jWu7AsC
DspCeYaftZ3KPKRak+3afb3s6o3IMhu+KWyfIgIVb0qDFYW4LHM3MJwOGDeFyG8/
d+17GC2YLrUE3UVJ5eboHQsS0IUhJLlmRyrhvGg7Rqrf/Kvxy6S/XF9x12xALfOd
Rpn1IzCT2acVVt32zM8kC/1OYTu/4835dIiHsZ6WczdICUjsViyT2+sW4PmnLIix
BhWBRtwDRlVWgOucfbq1/7IILO1cqYxJG438pANieWqpQ0SzKqS0XKylOXBJfH4W
8iLe1bFZ2pCkLNAWTt/OQKlz159OSvawdlPjSVoe/UvNVr82kQWtlPVX9TKNctiw
xD1iT6hyfVfV8tEWMh8Jk+84SylbtFxzEFSyJ1Ilod4pFU57jl9dhwxh/VV0ZFYP
q+q3+yNeqs54nucjePS0fC9WoV6Sy91OmTR3V3cMsFoU4CoR+lfApsSIexMsJ7Kf
kFm6MacmcktD/AJcUyW3E1CWQmk0o7SP/FYHE24tQNobSHTxFPTiUZakwW4i8FuC
pnEmkyXlAg+iCgjvDbIl5X20Xf84Hqxp8kvYwrnkcaSCUB273PmuzdovWaZMdybr
D8XR8aXe7mzziqNZqTQzD71m7Zu05kV3cv9LoBdyp6hGShuSw9r0ImcFw/jfwCGh
oHfN5oLvvRGr4QhEB5v3qpdDm1D0N0L3NhArdv9jOO6r3OH8kCopPa09+lKKclXl
fNP3pOAkdpXnLTVbhA3eYy+yaCml3cB3faskF+6FVm2i4WrA1xSt9OPAjJHUTEia
ih08fs9b3cZaHxKpJxWRL5PLNHRMeqvdqGMupJymgW8h1KYs4wYAzU0q4adpy5hw
bi47IVTsFqjy3hmLaQrEBnydnUHZsllSaFwrIxpmmtZL++p9UNp1eUjjRVQJv7Re
KnHyEzXCo+B64GtIQdk+BLFN/vmIjw2GXbpyiE7CM9kaqWBmt33hCfI0EwZOlyfy
7K2F2TUZqh/QKTW0Usx//H5Vc3sQtCfcfgJeSBoKTZxFPI9Kv7djbAllHdlftgcb
xb1E1Cif8SSxDdPdKe/bMLOS/34zC+C4ImQ54ifUqV5ZMgq+NWEGBDbst3OG7DI2
wJY3BTprMJeGM9vMoBC4Nf5B/JZzxmnvMdrNKGMSUikcsq3+StIe1JAVWfrU34ZZ
VecoLvHxCXflfkWsxvb9AeBDngnYIpoyAmXFhJjbJQkQ0M/XCtum2Od0Wz6lADlA
iJ7lPseIMRZuEp36B3sDgAyiaxr8TGV7JTn/dqJWUIbW7vA1Oii2JDFxmBs901jD
HKgafstsLzD9jXy7Vqw5JjPV0Ko01BaLLbXqdw7Z1vnlc0VqJEc0T8pkEnfJ9PQw
iLsj8yaIGx6IdSJSy+bYFLvx9e0had4QY7rjmFaINdQFU2poI7woAGNbmT2N8ITF
sjmRBbWsTjXmul7LDwV7o7f9hBFfBRjbv/K8+rEmUyw0gRwuUnlqqPvyAOSm7lIk
+/uEEenB4mwvviUtckXm6fn1rzx6YuM3nxcA1cnrG0NZNXuPYQJ++Oh4IVHVBWUC
4L2wBauBWzs4vmnmRrCV+g55Lg4d1MuqTBgC26y6eYFPdlIqxdKoSyiruu0zVyeY
er24XYVFgmSVdvMMdyWfeidyMs5jA9+nueajuIr4kPolmuteDidt952FygKBsKSu
qZO3qPAO5pfoKRyrknO2A7Kdu2gO2rf0lDXiZmS6qHyui8C0fENcKnRuCdTQrgKM
wEAKednIQoSggOyTmAuYevgDmp5As+/fvhV/IP6jmylzIcSn6C+ZtBdEg5Bo3QrD
kN68R35/1qcMGb4ejkL+8+f6NkQVownwMSWuGq4SNOTSS6BKu+cCoqPWv0wfppcA
iRuQJ3sLATB7vkJzME0xnMCmupQtptDS0dhgBY4qsJsyi+7FKJzuZHUCkLR9ilgk
luD8XBJBOjR6BuxJ33pSmPEe11o0rXxY787AVDuMkKUTCPdUB4lPmFukzMRxQieP
40dh20UveYyI/RrSXCwqnEpbijUX1hzeHG34bl5E7lPOT/6SkcNwGLarYL901WEe
eFFB8veNHI2fE+BELYOCE/c0UJ/Qnsgnt7NIgHcTIN964i3BgysAdtCax87rRi+D
BDb6/YEAblNl7QAJVqOSUgGws/6FWzGCy3kCq+L8Zryf7UUyyRWCfPxf0UFAoSg6
tFJ/kvgnic7+c/S1U2Ar8ehh3R4NadwMYBp4Hq4Qc/FZLWuAjUVX3Q5Y71ehtttk
uhyPz5jutIwyqLn+386jeh+3NzFKeDH5AM7/c08CrIR5IyjhaFSKpoJ8Rkroifas
+RGsmJCXroghp3WsdTDRSUx9WF0IBmBnXQ757HPhbS8MNs5rDJZZM7e3PFYlf/IW
d0jGcuctYZqbhMyGUEqmYwWtsMg4Y6bOAK9mf9jp4jkFspuenHK96ubWHSroHc0C
fx2DSPalaaYgyny1qb8H1bSJUnThuCPimcoCtS2nRHbfixC4WZGu7LOfEOJwH+kP
YeAnfMxfSklu2nuO7nJ4fZVLC/5cWTLgm0038HUZnSSfJHg2S/8sEVjISQCoVAAX
sUxT/RIjWxBul+WX4z4OXiJLWm9jIdQHI3CfLlunVagElzXW7HdU0yU4lhQdt6/v
3xsx/4P4ujHosJ4NvtAfYHQdWVGM4MBhCbAin1AJcnf8zRyqQFnvwpyM6nPQ1LdP
TePken6S11cBlhgHJo9ulJJOs/OCx1kMTTKng0y2TK1s9ykUTesG5uC+vIUgvHp9
VJcynZY9u0vSjiBOA67QNNZ91IDkropStzdHdirX986jLR/64D4ogQN5P4DcLiVv
rh5cLf+9V9rPYbUwRE8gOjzl+gblPZljMMI2Eg7YPx7wF+joRUNCRFDW17i2tynU
gNuTBpEqTzzTQ4E+N7DuGnR9tXiNdduak3b6847Y8fA03ahVeMgZb+8ReZXozvAn
2Q5PR1v+i4eztuQGe0XfgJkIXKDPRNDXwu5sdj+iTXhZtxM/w7UOv0wMNfg59aWG
1xOh76Nw7G21c/bq06nszeNe2FLyt0LOw0gX+EtbrcoWQUIONPS/cf9Mtt9jylX8
MCNbLcj/TeZnydUllclD54myUr9nC99JLfRj2t67vhWxCV8g8fYOFbvhdr12LMW5
fQcotdQOOY3ohzlfqBL9TJXpd6TfD1yXrPKtOYB5r9D4akJRfLI8s3UntZlzRybS
hay03qci1m/bf9UlVCc09RfUjLXtj9eXkiLCmVlTCD3yiAUWnhgJsjyUaaJHOyu5
nb1IOrA2yiLy+TuLciCKkNvNdr+ZzsNQS/ANyE8M14ZE0rILsn/lNw8lzT0SomQG
zMBsd/auzFyaMeD63qtg5PaKsVAVYhGNHbE3NL/JVUPhq4G2Ug7azN/8lPcSapf1
wjsmC6suXHutIUPZK6m6JMfQfDTtmvGZPjqB2i6PcIvOhJwzEhzpM++p3RIOp1Du
+HWO6jDBqijak/HG+G6zXKdLHb0HsyoA0oRF1KqcapkMoCrPcm5MGbguxk+OAVfS
j+K8xfKaue+2xNjlECX4FV9BjQxHkwXikCDstMbrNX/wZgH+sJ4kevt8PPjswJ7X
7T+YW4LWXKXEz9s1ciRqC4/8itfXPFkAakfrfGJmBOoD54K2IypDubuwK+mxGw14
Q5qWDz9UqVs0hFrrVyxTMVeX4mNYGiHf10DOAOhls5Q2M/Tm23oljr0uMOKLf3HV
aHJeW3m6+WwyG9uPFzEoYNHKEUBzGwl9bEucu/mxBnyWGA29pPvwHv8w/e1s47Vv
R8xLRP4Fe4ai4nfFbRgeMowQ46x0q8WlyD0JkyWWonx1a+PjxEGnay4fdx6kp/Ny
I44y45GnlZnp5N/mFbsuYuUDio3sKfgI5DilU5i5X6n7Lpr6ZNUg71eDwQV6LBsM
+cl348GiobGxEvrbVwgPsAOUcdGbsuM0NOKyFBDERT/1ysCKIlTQ2tAIcePQp4cS
rXLXHGEz3d13F2/j5W49fuJCMfB66qh5zDxcSXD4iIcEQ4uXsGNPBtJHJqA1VzA+
s/ZOojtESwmPS7wmpB4TLUj8cjkCLMT3+F58UU3W40Nveky6hUDVCih+dD4QR8ZV
+0RKNyiMYNkK+pqQ1TE5fSAUD1AzRA42iP5qVB61vmzeiZGDIbzX08FMnu429JX3
0Y+pYvgf1ig8bMEfiJ8+LH5CaOP4gSctMazSi70VvTiPFAn8GLVmBPiJ+HSEb+/i
IT1wRObcw+8TYY4l+FqzXSEwTyMWh4kDhrmkMtxLb9XCX0Pq3MsTO3SGgLzi61E7
jtOU9ewNLNhWSaWqzIOYJMB2gsKisJ92m3N26J8JVU6bySu9Awv4BHbRW90HXXs6
JQ1PnqfzJhLfF68IjFcX07Fe1c5J2AU466OSG86gDxXbNaFAIeKDlF148vzuytv9
PTprcykaK2JFOHlZxoxfJcWbtVqtkTVYwm30Ik8Ybg4pB5gLTD3XF7RHquSrWURX
h48kuC65gficsAKt2keyRwIfpfQKkIhxbyQjIOCw1hYp3/6HGQb3nxQ+iv2XOeZI
mly03ET9PS8O+fpUBQhQ3IxnczwdgjNfTETL7cOU1dGH8MK7WVW/nb63nT1Xb88/
WPWJfXIrBcazCdkQsHAFgl6CLt8Yz5sjDLHG+orYAjXxeIvtyUznczqOw3PUJt3T
uR69Rt+2mdfbj4nWB1SdFk7doE4mWMtg9to1UY2gFAteKWrM+VPn8IMl9XhiOgew
8rVZ4t5hYoYVvbe4OjSUuKP48pA7S1ropFuk54lOliVxZ0zRnzC94LAaeqCS4Hk9
z7eOpnBoRf6nGpMnQFpemFswYIyYLBL8QDctRAqkbEAh1Cmp5ODe3b3mUgJo/4xX
WaIDex9+bBq/X0UopACLqOrUMt3syGMeSpfJtUQpNDJfaNczU31Jm2yQ4eV47lpk
WufdbK6o9RgO9dAA/UFt0S0w3Bmem1uItnNm/dwrekt9t56hh1F6wPu31kAyBjKj
8r4SZK6JCWU97iXuCBcS0eJ+x1wCn/OgrvoA9dc90bFkM+GmIYk60207OiEWE5d1
ohqw4MSkzXTVcfB4TaP1IC8g901VqRYuXu7BMmiOUxa5n3dxIrhU1dLHPPvY5rhk
XRsL59DVKPJIjfdqlxZi4TZuat3hsMW/7U3a2rb11vD5gOFSMx5COMjKWEb+57OJ
akWLM7CJo6elemU9zDffZDFZzsd/TY/Sxti9QvY9SAXMPjWjoQeTE69CT1o1OE5w
QySUEt9NNSmy3BsLJnyhOjCPzt6MYP3W06Nr8L1kxCVy/9L4ompMq7qXML5x8YZF
fEWHpSGCVYnqDTiLB8gfsAuI2YkTbTEljYoOnaTJDRtavRnz2Dmv/ZzYXzgyRZYK
ByKi+0Uoz1qZKig0RJBnVBZnOPdCu9EAZG75jAwOuXEwG0FLu3sLVIw6cJYozt8L
Z6yGInDOAPmxqHvNX/hLdC9fhqDGhDVi5D/7aZR4zdOOGlvQU0WOFVIpaDknnPmo
mhaLuZTHFRChpzA87IHUwDj1e1HFwkeiwbm0PoSEt2c2NfVyReZTnnM7/k79qVc6
jCCqBtjgNKOf2r3yi8oZhUhWWxSu9xb5bKz7wKQLCvWrmBPmQTbGY1Ai+8MfWhd3
Pgf6IRAP/Cvh/bvrrkraXOSOJ0WdEmbUPfED28qb9QouFrDs8GEF1b3l/e/kDpCy
GKhv2GNyEzVnpGJmiFOdYjZ7bpHZ2Rmezlgcmp+fM3ruNoRz2rGt2I5tGqo6kCrJ
oOY2jjtcCAoSluZFIdJl+aKkRRYjEwdQat3FGD2Hv2bcau5Bj+lKWrHk5oW+UqvT
ZC/sgtCIcJlg8V8kApgWVndpePSOWO6e1PQhrr5mWDMHrZOPqHJbF4QbS8OMl/4B
1RCvwRAZYx68nWfCAKRsA/sTbmJsQhgUN3rGc9gk7OViRjWHNz+Xd6cKXT24oXzg
L03wAxmpf6SLt1qWezU5ys4Xhjo6e0x6MuD9D2UblcaEPoesBzIQXNUYvmmumXk+
QsDCaGfnsfvFb8SL2+WS0j/+fzAQLkBgc6mY33gesoZymVETTwuvJamBoPpv6mDT
X0jG3eg4/HXI8fivWkCctbIy5ViT22VC51Itsy0zcnptkOfu6oAdfR2JO2Yw1Etw
EpzfHl9V9HxQTMFGq4Kc0bE7cupNH9NrbqcBSLzYeVjXSzW8cQSwiD0UqVxx/KwI
I6LDGwYDmF/KxhDTK4Up1Fp3ZaDXwt+2lQI06THO/Mhnsi2y3bS1DcXtOTt8/AuT
G/DknFJy1MY+5IMjXxLwlkpKz6SdKfKRcy3OPjLWFHkDQ0JSWDSw54W/Na/IMmev
PQvjmp9wNJRB/dVAOwOU0i1YD3S7CA6zpy+AN9fF+oCWA27CTOIdefP26beSB+Mv
KfZ5M9FE3hYDK5HNitw4kXz2HsUEyoPoGhNlmd1fYM7Gs93n6FU1zap+9QAJYbra
hTWRI7Y/wM2cq5/JEhXzoFhIIVXeAiDIuxt7mtM7NTsm1YO2Xp3IUjsUOEvusYIj
hA4gp+XmZ4zA+nSui4ktVNbTIhT83Pgog1YWpZCcc82WSufvRM+oPSeS84zIBQcz
TslOECExbUIQH1yNKDSOxCuhwXpErt8FrZOXvb4VlXm6HWo2ER/FmeGQhndTlqux
WNZWmv6DXbbfxq1rgmz/H8Okkwmfq8OT8XmJhhbs/Mn9IDRK8U0gJf/RoVo5XCiP
rbaWqBSNaRDEl1XxWkIPpPzOLtV/6hjNxiYzB9tjxloq4dWOBQzBPBvghZIOJ1d4
ei/jligkO6HrdITxbUAQ2A5G4qiRbYDv4R/Uw+A6cxpEEGTRn3Uh1w+dN0b5Skm4
2gp3rS8PILdqXJ05Qk2dG42gxemTvlxRVROS3bfTVqNKEtneBX3zftvm/ezfBzM9
XVq/vKWwGnfRcaz4rH5J3AJji7W9Jiqj/s4oUQp2Y6jnV7Sq5W7QXHQYhhTfkQ3V
TSbG3Mp6TVhAOZjC+lymRGUO+EYsV9A5GW+wjS8Dsm/Z56t3NF/y0zJABG5upGUK
ifaYePZ+5xBg4Bwrug2lD4Ts3UzkIDxkZtd9HAEsvs5oZewPsA1SG+5+SYHxH2W5
sLRnzB9gu/UujFvEt2HI8G+igerGqWDS8ajrmnPfcGqVJrIJlKiuUIqjyfiUpnkP
dFANiyVk5FZ3gFEaJowC/AaVjn7lDTtSusiJmTu5CzT5/nRPBHDXzx43w4THfDxu
SjdKxxkgHJPm82xcAE2gqJWGeg+87g9MQP93QNi/306DeJjGq8rK101gSr9f6cSd
xgNoNcx6GGjLb3tU7RZz9LB0gWRQXrYVddQ7OG5XSwF3d3KmXatC/DpHeKlqF2n1
jjeqf1RtNpUueMj789xlCp+KMEcnShz/y/embApl4gowJqMhMtZAKpWz4BYb3Oq4
j/1Lez04SkN2Ykpd+7KpndXKVL6VujaddL4xc+K2FDiYA/4RweALjcbq4NhaqPYT
ooHeSexFHjWSio8TmUpEtPMfv5hFpmnyccWBH1oMm4ZdzfdksSHA8bbUZU9KqKfF
/vIuEjCXawH8dNTpI2CqkX3UOnaWZKumunTYgympclST8KiEiHJl88eucVj3pVZv
ek/p5iD5rdJtsLMAGG6EB5IuV1qFi6CI3HGtoICiJcBhn4oabCUACv5nYIn7lanh
a51uS1CKg/On4lZE0OVZHc64r78f1SDfBoUvUm+o1Sd8mukwgk/fd4f6hNrBGNYN
0ggdpIrDwGxSNwkRVa5tHwQWn+Ac5D2qq5Lj2dsDP7L55dwFthrhVLeL3OjAbCxz
9/k+uhpCnzm6Tddj1VTLi+z2GwXwBOd2U7icg6TuiGcXsMkjcaUXZuSPueXqyPnC
v6atjL7PGeGs+1ushvqyGH2USNZBwUW8wl6s214qoZevpA2AOEE5dtdBhN9tfcEY
0fzg/9qGU2Sy16ucjY6og+KKeiYMuFSt+gRuRt8IaYgIZ5/trxzXbluIZNKSGHUQ
sq+hNUKBBvg/Ja1y1I/Et3cDbTGJBnuindKkd56yUQG3jb8nd60vX6/SlPy2oNHn
C9ArPr3WimNlg1RJFj+oMO8HMMZKq/7Zs3UmtRbyKPjK1VFIHNL3osuTKvHmOTqn
d1Xrc+JqDZMgDi26PmzL04P+yer6v+jIjbGrqj3uRlHtKAZcYOnXoMaVkEvn6Uoc
R3H62nJE4Ruhdnos7kISAycO6kbNPH2sf/9DesTnxhwrTeZvpg3+XriPNZ3ZRGpd
UBZwuqpPfKTK1PevXZJ4HbNT/ueSRGy+g6kYTAx0GPHmf+c8pwp72PoHm7jH3q9i
lgqRb3M2MBhVrhJKL/nhvFO38W8XGDsn4J7qr36FJSdLlHk34AbzZx1CXwwqz0m2
sxckJn05cernn8hjoS5uHeRlQXBe/gE5hr+H8ihxvWC5G/Jpmay2Jzr4xp+hvMNV
UOifR0wjEoqWPxNT1P/1YlTwBfVbhtW+SsI++B1bss8YcRH3SbqKJ3GYWSyFuSmq
9epFfApmNO/T4mEEA7vycbjDFPmi3r4BA6ZhsIbx4MYR8pV6HMNQkpGR3bT1zhlh
Cv9JCun85X0USe13I3h5/KXfqe2ZYwZTqyHFiuE1DlxJlavNV9vuNhCT9L06xaEy
GJs0pmmRS/Tw3P/yGk+T9K2jWIWI3rlC4yZqBfBBn64SrncDzqRRoLG5dWjADMJ3
5X6nXa/TE2F9IQCWASev6pAir3iZi1d7FFYLl205rE+wnw4pWWbOlRE7L47bdqc8
mjz0BPpcCJOiy/+O0IymmL6b5hGk54RNCtR57rYhfHXom82jgXIGCbKYI4C2eDGi
NG6OADuWhpPwef/GNxMUTkvi0liuNnxzK7I7B/yl1Fpza2rZrR5cSsMNyAs4noyM
5LSzlrOf3EqudjnF4pmHcgPns/JS3BnkGjgRw5Xjj4IZ6F1RTSfpj8pIRZK3i+fN
E2mNHrjIiz2o6E770/2gNcGyZuJpQNVa6f68u7dAp315rL5InLNrK4tAwiK4ScNv
LY7+YyvCyBBd34x586Xm3jrIeB1iFUjfr2iGLbzgw6X4oWByFFg1huQjhuvcXJQ2
lkiKtN5P2VZoAOKmjNhmj8Z/PqJ1Oqgo1SutS+hP+SdBb01++9Z9eVdvqAa4RqUN
/zRA/sFpvFRvPVyE/NsH7zuRLtaUsS3Um7HQFHGsy4t2x09EXAhmy/EzO1OO+FRW
bUo0cYkWmFcPhL7gAUbc3OuK+rdgxHdZCfHHA36nncSCbdSOoC3t+jjWtXXvZQpz
+VP8vz5Id59eXjc+XwqEz3MJnv8MPMtUfw2rrqhLQhmHm2G4wtHN8pIquUwhUroM
T6ggZE3yDrBmuldb8OhZsOFC0EE8iL1BT3760E0xMxiEUkcwHmUQ86Q65O+Bec/a
jpwwmnRuORSjbgC6sR8akI7oADGA6AcmfdJUfTlfXi829QCHB/dVLWdFXMAQe52U
F9pgjLruXVrEBCVuQSftkcUxe100asGNfgQb6IjjlP2KjWm6L1BKqHwsmz6aisyB
Or1ume+svJiqPuNXubL6Ea3yvDrGtPQ4xMOot5L6iAgmfy19DO9jLwKHiVJpohqw
F3fY475B1F/wcBvemqwn4qI3COgjt3mVJikDDPEF83c5lG4Mrx2C6c0SxQ80MIql
MgTivMy+NCAd4T6spqkhvoCQpI7wkzoE+HoIRLnul4PZ80Si5mx5QgXTVVEkggt6
s3MR7xuhP8OvArI161pp5nd6rDU2zGv9xQr4Cxl0a1PhIzoERaSqgYDw386ivtbn
2odVjMnrQ9OLie2oNXal+AX0JI9aozp/4yoQ4dKl3GPnvpvwxtcPE+OzWyH/K4nb
RyFl4/Nzc5Us351Pa3W5emdlI+fVxXR//RjKlr3Pzan9qGsny4m5nG04Tmnd1dIq
z7KxKZ1Tv4U9CLjv8BCVtYqHlDpe8jyOH1yBSiiGJFt5v/C6W3CH97VgWOPcVif3
fXuPr3os5y2hLSohETCPotvwgsKGnkEwiazZdyD1GWTKCCk/vQD8vJJ7/4/9QNC9
dyGzaQcmycGldOZN3eOTmK2MAMSaEf1su1QvP9WJf31oO6yPAsi/uYivchnrkWI8
/6dVtgcPo51qP2825mq0GLuENgjzBDvxHe7kvO+az5Qxmx3eTDtwLs1dljtbzX2v
pAbC03qLhG/vDjf44yAO9zJlP8WaX0NcFxXkFDtkOUhoqy2l7SNaQ2cPT7HyF9L9
qQxqnQxEUUS89F7lWyFSoG9fJhlZ9jefU/4gGr0B7MFmXtB1HbFX9+jQcXpCeR8r
uzyzAag2nZBr+gZLL5+7soPZTYoV4ij2x62NQXTXuCuBw9yJCq7EHiOkSL5LWbe2
QBZvhawj0m2ayuSlId+SHyyqDzSFeuG2QjD1Pcvh+QIxdlH63TPdh5yD4wLfnKIY
Bt6ZfeB+KIKcCO3XNbCIbqnoEtGexIAma7GJ2cOVOj2wfz69P5NRn/cgt4Ol0MnT
dhRoRV2gnEIAzi5VVXkriUaVbwcLQ8dcOGBdrMuRIejHmVnQYrdUBtdRkxiEemaF
Vly/uyHUAJqV6o/eG+o/ysG/vWBA63EGFn8CY9VQuYakMsnPBYjk9Gdmzi00rmT8
e5sdkcVRYzO9sK56Rl2MKRPwNL17o3cWyUgdQYUjiTa38IY4mmzOt+aHSh4vx2kE
/jeNrAIWdSHOKq9oG1hL513dXJ+sKaTo6IJu+C6csLytvHJ5MKdobLHWV4x3ktub
r+EXCBGwjulAVVpC0ROtgMjhC6OuL6LArwXZ7zy85Wc45Eje4Kb+2n9FqbmUYd+Z
jG+3CdvNfBC8C6d1IJhqEAJ4lJjdzHTF8Yht4DnOjSJoMQ8EPLAMUWbjNFBRBgg4
5NRQ+WKHm46mtjxDRFXy2T0hq7N7h0NlR7RWKlGTYGEygwaXvdpg2k5LfQ7eEZhi
GDPTf0VbZSJLPtVNXJMg5jxuMAoqApbTUPpreWrSBESTGbVmvxzRsMedEV7896aT
lQc5j/e7l/6QieG37P+Xt3Y8d9MRNkzi1LXDuNfgAEeK2/IykddI2Eyp+JDnbMij
Dyvb67TpfBmcyn8Pz1HURPXiWWuvSFvgtd7X5Jo+1RSv+n97QdvhdbVpW/OxaK+p
y9GfuuGaQxX6mhY8L1vGF1CbZlOWmslI5VEPTXZfFQK8ibWzwCB1NrmRRQr1p9jt
ICkgzIz/gAztgfCLLdX1QHWarQqTd+p9OgkWYi+iw/RJrcQSo3RppD3iMKK91pnh
o+qD/RLwy27iRtATp9ANBziqXLugbzUW+3+oe3fyd0c3Ioe0eK2+yfr0R5ySyxo8
Ds0g5bvDeYTHFEZQsUk9JxyRp8Z/2EZv7/t22gAWtGe/+n44Jxt5hCfIQ8Ab7Ahx
bTeHBYmUdy+odtZ3BX1m8HZIDd/N1FVbnfSH71nphGA1ZGHVyfLyTRKFiyjli0I+
QPdq8JLPswKkhNKYpuUotZWkhWJWKViL14Cv7zy+70WSVJ30OSjSR/F8JzlMsV5f
+jpCRVb8Y+FM1wlavfKoBNxvGsRJG1yjYcGyezaAtKHwq7GuIpND5jUWb7UZu3zM
kEBuLah6SrrtXNPlppHGK9/J00leE6xT+PHBquo667INvaiZU4EiEsPkkXWuExZj
6662JqLQoAywtyfTr7PIa97lxDEMZ6PWiTCk3w3Yf4x8jmWq4qAM8rOLxKno82Qg
t4OHLq6LT/n5B1z1Hsg6scO15y1IT8UVHiIJpn5Zi4kW1fugzyGqaiWRSLjpehFH
uZN3kpUW76MARSwdM5a+uibGLjMSe7DVFvcLXIz19AVeFB907QjMfdNtdkHljctZ
oKv2FJItWuH+rod4FkOBg3jcpxR+tR/IJnsu7tk7aFkYFGPjhwbFaOwOX27cN86X
nrOuLW+D10X+SUC5lLqmm5smOYV/97fdI7JN/X+ey3bDieG4Fjedyt//NSD2QJ2W
1KA2vnuVcnZ+RO1zdMwmQ69Ga/P8aVsXdUIyZPgrNkaw2JDbMSUFmcDwEKxxXyey
3D0Lq5ZDO3/8SkQQ0sXkbY3lQNgrjwetq0oqopW6v8LT0F8uo5qmBIbiRbrwBEa+
x2DDgzUTEd5pWTY2k0hjLb8QYTDg3rKMaF7y6STbU72xcC5GMUB718t4rn8+8jEL
aa+NuHyqb8Y1npysrly1WnYnteBZuDpzKMMzw2w3IqKjcwlobP52Wqucm4wcJThY
Xvr37FWt5uZN9aSMLkYoRLnb0N0W/1yA/aoBKRPOb0GaZvVYNWQdSfea099truyo
GOSLhGchdSidKt4jACcM5UMsxy4iQpQi4eRmnWsFXG6t8JbBOBMiqAkVmoNGJ9G1
spLPTPyOdh8/j4GIncLi/+qJRu7sSnBAOk2NaQNZ44wanv0alR6xzPQbUBfqGeeT
IWOmGfuqNC3ExqZ3Ds+Rzg02qQCK8X00Z2uGwKN4VRqV4yASnXquUgFTVaJTT9N4
1vt1O6czjcO2NlrFyjImhfUXNsqZI9N3GlBkJ9rwUql6FW5F5ppMe0UsXBxqh0CR
pC6oMDIewApk4Fs25kGMMS2E32GIklKA98Z9uesAqb8hDZ1E7OD9vT3QrRGspvgB
zpXVvrIFTb/ySeGLPqJygYoZGe7BwSNy6Hx0t0BuVqpM426dkC7b0Ao2hrrflR0p
jECdXDNoOlVBh/ar6ADpvpjL7JzTHe3ZmtHgYAguHDx9DRwdUSFEYuWN5U9WQB/1
Mg8WPJUrURNwSS0XYpGc4AfVV4aksNI3ug040eMyAWMAzBrO5/K4PTXm/cqJd8mN
yzrXCqfJ4B8Mz74LW5XvUhyVPuzNYet5Ki/TvuY4oP3kKqH7LVliFWjOE0pkKLJm
jQRpaQ1DjFb2U0dj0XjpRCM+fyW9zU3bEOuh6ArxxQxeMARaMMn0zNp2hVRZeAtz
Abq+pm58j76HjfQKfkMS23FrUegsfQhrzOHLgeLcMkXc1rYoza2FvVlCyoxB7mEX
vmGYPg8C3jC+8OFj1N1CVa+uspmKhdTBPEkv1Yf9BZyRUFAXJc6v8xMSgo/O78MB
ax6NjmLlJ4hAJ7dTuTwsbLdccTj9ABS4XEyQXbuL0AycDyd+Gw0Jr5P4r0Na+8FV
rbPq7ceD7FB6AJe4h+9SClcc9ZYp6Ppx99hXhZVKPiHzZvQ9uWWfKZ2QrDvFNiLW
2EyTtB5GdziO6874Q6zTYNI9tCJ7l352BFNCk3n6XFiC6sa0NpBE1uL0wkOhRhWq
MPC42hPE4VA63oLvyz5A9diy4KrboyJ+kUQiYRktBP9n6oZCm8qe9LdsTCpLn/G9
YORT3N6+D4+K6xsB2bqVpnaxKQ0BppJ/a4L64qv0NkPzEemMnoplY9rvDXinw3TE
u9WCqXJLkT96fJm89EJF//ki5UnRJTz5tIV6PKYZ4DdcBD4gvIuwwrkeV74av3k0
yvFZqWlcmSvnatrdfgsaHwvXVZf91gtj1CmpilyxJd/hIAJ+ojntKc3Fqb9Y7oCW
F7tqcMvUVzX9+iTDRX2Yz7ihtc+MEAzScH6WGz7CEdnMBZlr6hB5+mKiyp2Cvdv6
2qdKYAz86jGVWt0WZ9xDFyOCshsZad3oJDDipEMvymLfat7N0uHXWLIZduqtF0ZA
8LGUWVq+shlNo6drwPDXZlvSsQarMfQ0FYRcUN4VpSVwhaFRUbhLZ/uw7JBFwbe1
KcN0w1FmJX2F/TeR/pEiQsZabGUZaSPxJIprPxG2ybRvnamMrakNvzTf1lJb9jGf
6rr4mk9kjxSW5URA3KzMOAzfCEurgUr0KrG2pDEJ8n3MPl48uI723YyPW2BuzLjN
80R/IreNz0qW+Qily2G0k//sk7KCmag1+7ynMaaRFBGgqlqaaDw5QLrS8GZJEq2Z
sf6NnBSif/SgqfT5UT+5D1iQXDXlMMVK+8iGObtWpryl/2AWqwM4e8dQEtertcXa
yZRK5fB+BdHQV+bO6eCxpCS9Sh3XhK1FCrysTKqWgNTn/GWpWYuaAmLf3JgWCxyV
YUpeI4wL2yUcBF9r64FFJAUmGNd3lP3QlwCuRakGCkFs6cNUqlJ8+QNLrlIb+LwT
h7y6ZNNjw4v2MT57to7YzqXBs/Ty4iCTxEZAX3peJ8rpPylYVCimePtuzw4WGK2m
61Z+1w3PZYwYHFnkt2jurixRD0nB7miPoHZ5xyvoDQQQsOJ74FAcogTSrHAKgNlh
5hDHFBYBJ4zuBfLlmEuzqmcAf2i+cPfn6gO6oVNrQVMmLiqjkhKE8+i199RyA1Wa
padH5fcsZt3OI+vwsGzZxo7s3TVall2Gzj+Z4A4aNt/lfBbP4sw7biJYJT35gXLt
fSy6qrWyZpCe7m1UTSZOkKjMcp3GVSbrqpen00Vviio+rcuX5pw7uJFkvlLk5D6m
tHoZ+fb+lg0iWF6hcM2N9pE87kXr7ys8+xVzw+UmNHxeJN3ziOujxjA0z8tbFhWF
53E6/yMRHN3efOOyQQfeKzR3KHzc48SeQz7f9k9zt1hVzQtbrkL+bkzL4Ug9Pav1
4g3wI/+Yj9n33A9dD9ju2ikOPlcSBdxFMSkyqYf2Ic07k3/zomXjeXfRQrLDrXEk
38nJ7+pbJJWS38afyV+IBhBmrETj7Nwkrg04xKH9Xw1SS0AatIccwYgLkqLHOL2H
cW4jWSbZyllRrUTiCi2J38hwyQjWFgPu9D/S9hzCVvBsD8XQCD2br90s3opPJwBX
EGALLIhvgNozm7LhQkS9mSE81EOMpjb03MAkUzd8h/luc/JW3wmwmRKtc+iEUn6l
vw7jflFpRXnrUklztMjiCC3CnLdFI1ZWMFxWwZRdByUwTr2YH+yANMXKS7ekT5Ov
2Yy6Sda29Q+rkXRQLzpdLsnVYZUae2utpkIGxCQy0512SmkhdDFhfsUjZzwyJNNe
0B2LIS16eD8R7rUgxMwxA48Ud9O0/0ViWDkCIAztp7tTMHKnAdUElJpT2+OXRf72
8jsLkOR1yQSS6mprKi6DqJb4w2QA+NHTl+V+zap/oWeULTUHOCsLo88CbenPKRAR
uSzihgyDqP3TPWOjyfszSlLfuLlWBA0F93ksYtQS52Fim4DcS9QtlX7IPAK/+OwQ
W1fwQ4ykeGuRD717h9fYPPK+mPa+T+bv73RItCaabAuUSYiJDP6uwJqT1vfg6b2O
DjSf/SplUeRnAh3REgVZxspaVHtSHASshOZ7xvOarHqopFEsok5dnQm4kDxR6L7p
3nBn+GlFs53ViB8LxwUUH0BhgyV/P8E2oYTeOyVyuYaW5+6A0HkcMj5F37CEDMdE
qTLCUx9da0U5BHWuX+fVivUJejcU5XFqHUmeqezvVn1n4bynbB8eA4YUCFI5n/K+
J0RzYu++6IXqiRy2VQUTsLgQgL7lEBKJ20AWw0vUrR9zXy92HpIl5ai+BFMO7Ins
rk0+enBHtikNLZzySG5kKc6D7841J1HOmEcqo2rnJloa3gYrHJiPugobG/lyJ64x
YxsvgHWREc3kcsxIxx4Y6FYBc8hge1m8PQUo2OBe6G83GbYY72cjIqbxCtUm+lM8
h/8Domq8pvjYZEW9PKFxvVcMMB845apULdlvxwTflN1ivQKiULK4Ma2oaZwTFzd8
Zuai84gPEO+SjYzMr4PXyK1P5ITNhVn1LI+j7fujzStc2J9XZhX9wpkq4/5Bs6AO
YIJM+VsslbRZhUrB3+LfjvwHZq6qtZMGjFQ58B1KPUi6zj7sNL0/T+nIJRpA9dWr
d/BaXsmAuTKJe3486j9K4DSbegXrItFuhQ0AQQ+PfXFoNqaPFDzO2gjV3MdzQ9Kd
z7QoqowDo5qAwJ0G0q5o2XbO+ANgzCfoAVXddi76/j++jDJD6h71kZJ862JdnB1y
OOWhANFb/Mhvw6d6vc2p7sgcsISuF61Q4+yCiA3sk+pWUK1YW/Np2f3H/6gjIeKE
yzU2U9ANeqn5Zb4L0GziUyiw/x8mfmTnnBp8QPeQFTwVTVsmHNu38+oC4vJkvsBc
mQ+wr9djmH37kspZhG92d3NGneLFpjBqk28y0w9msjIv52Pk2XpbXyb8ENM9YQ6p
ykcT7N7FSuzYxUaHkCkf+F+wt/JSIf8YVXoCjYuY++JUcWCJMpmgsxaramwv+SfI
FvZbwcRBiWoRrI28w+hM9tEQ/e/XH+mmEnf37PsnmokMM86XiP4KQpB4Mt9mU68H
gjfUxu1BJw05yWnSAWGkmg9ekSCtOwR7xb2uZsW3xvsRO40rlO07V02JF6gzO4xf
qeLZvTKVDy903IODL+HGcVfA0tGflcUig5Sr/SWrp+sZsYHVP7b3L8xmWEiDn1Qq
izQfx9rxXg5sf9SL4E89KjqD4FwwyWQu4mcQo44BkYg1J+XmQl3eIt8Wa4ZFa5Ay
H84eqKjxuNfys+w463d+n4TWvtOqZS8WUuvq7LWnOE2p7qOh9Jpqgo1cRySthnSu
t3PEuNvscmqB+kccAfLt6nUYcE1/IVGdQ9cRAIGCC5wFuqKCDLQ6P2lSZQqxNWLa
9dwkNkAE0eOgSD83iMyE1f4S6t2VwBlZ57arlaHD9i+HzxNfdGTBhYzAxU3nG+LY
JN2ggaXQJoQtrjuSVXV9usaYocm06khAgqKzEsHqH9C6Z62kEi7WWjufF0B0YdTq
a+sGYAlYnmiPis1YuJn5ZYbecPxnW/IkqUckQQC74lIGQAWl/wcfIhuB9xiDChr1
MFVKMtYqWCQ4ahghGyT02M5HirUyfWr6lz5YpDoiCWnH1gWL5nPNm0Kv32GwFNDr
cZFZUsAMm+B54t3GU96RCcw5k9zo+Lc130rFQiip69D2YZCFbQLC6+gL3NgSK0Ce
dtIw0d57MeaqiaHn7igIc271T4NMPthj7RT3pX+RL846h2ganJm/JgqTYuCxKitM
Z7xBDXOnz4nX9cwLkthk4HztdlOR0BZNB8q8y0oigdQ/nvMlivtwdE6tmMtgqruH
1d2cywGVxwlfZvEeXd2bAmRq/LCygZ4OaIQGvJLmenIuD5qWOAJ/FwQe59SH+PSX
r/I89i4YAg03SpWAU4m9bDFY2tLjsZoOziC94BLY28xeEY3+xZZaA2FvM2BVONww
FNl/dKxHifyVUruiIt9l75VG8M7Oju1w9YbLdt8Ydug6IAJ7hIAogFZNl8zz2Sn9
01iUE55/z+wiKjISPgk9PQ8iacAqT3b6QKN0dVSiO72aAepUBLaO+NZx4SfK99d7
QfJIxZebfE3bOtSCLStRuss9W+tzf08l9o+RN8lnUZR9FFuvO4Tlww79SW0Iztt6
UQ7Gat6FAGCTdElZsjWdbjWL1Z0pQKRCEumaMItKAQI734taefMLn8vGZaquudwp
J4K2+wzFWrbURMrIuII/Z2J1lZo2Zk6Ln9wMuqZHQrpD4QJcYhtX1BHOMdyJK/1/
IcVzk18Y9BDUWb5O5mPzZpvADeKcTcIMDr4jHRNP8CFLwr1912mTW+CO9uWqOGwi
t1gvo5Qlx9oGO2HY5AZmRALcvF4K+RgmsTNQcZqcYm0fZSSbqc45z7btHop2WqtE
BoRhVCZhFdbgAurcF/aC2VVx6rwtSDIqffGHjLWcKoJFSCFnmK/Gfgtj7brF3adH
1+kYP5xGKSWiX7BxhKdVAnKuaXg+fdELRv8IQHxZBeWmDE+dTDkubTWJ5q48CWrv
mPuYimVdT1f+wl5iDTeFFtiqAJcQPSq7IGD0K4S7IIc+E98ZEu5/eEu7hwdTKf3i
Q4nGC3VLvNrJmj1n2+0ET8EWlPKXhrHukOUwQgFm7v8b+jcMOFpfHOF9CyaRtLJx
2r2uzOH5IC+uVnOhZk+BVugpW8GKQkfSnNW6cwfjOCR2D5moDIYhYKV6MD1CqOS0
8cMkBFHBA3uUUjWlw3X7Lmu0X9nrFmwbrZt4mzs7g8TNS/ROZG63P4s+E91alhAQ
kVSZo0KRHELjvW3LRBlSYlilpJQ5mUwFKWnE92RvT3VSFrxKL+4PgVBO4R1EyQFm
7m1WXp2qWjTDHRNkMwHZhlVSkb5iYAPFT2412OOldUTLi/0DnumjEjr/T3ACVPGn
3VvR7tnQDUF2/FGWJrWttNY27gxDSmGL+nSc6ESW7JyBxUy9u0kYcsmEvCYK2fB9
nwS/LfkEavp6s0VND6GESvMeTM0//E18SZyv6qw9QtUK9cMeUIwY8DKvZvGE29xY
3mQIA+IszPkFmBBHTYHG1Gf87HzmS3ZNE5MYYQUA9LHSd/wJIB1k2jJoJ1UGmKvo
Vv4hv/lLkA2Ry7T/BtXyYXkIAMLrm+3sb2nAwHoqFPA1XhtYYzMgKn8kH8oY4+Dw
wIC8Gh/XH3xk1fLh7NSzEkI7rqOFjPDoGTbriknMVxGGghiluRIXyoV01VWmyQn8
dvQu56w7qGvlNT7BEolxq663YfB5j6gldIubmaMxGOUt5QbLLtzRADR3go6wjKaI
x5Q5jFRARRWAM7+ZkIN+cdF6/xuyHyozh/xbycHT9zUN1OYUY9UHQNU46pGdwLfi
UBDxzusETbCSbY/KcKp6sjOwHX92zEVVMiCw0aNdYu+gxnb87a9ctzfFUgyhHl7s
WrpgBtn8H1zeAbe3iqJjAHzcrDAqQ3v8FCGJrl5t4TakV7AhAKz1r2Nfo3kKeyAp
Z7p3Xt0Efp3EoE/ux0iYkYKWZR4v8aOy/HEaoLP63pbTIjCulWxl7UpxyZ+qsOif
65jzjxYRuntD82OrlEaUQhX/E6ma3bz3Sx23fkpPJWKgriQKu46tPsSW3kkyI/VU
GHBmMx7Q8ZJ+f6EUwAb43r/y+aWhKXmfC8iAKmbxRVQMQ3DO1Bjw9kubrUQC4DHO
YNsXTL7fM2lxAtg3mNz+dL5aaCpSeAshFmq4c/lODROm/MrUwCv36d7+6QwmYRiD
YKpbb8YEe8qQwDib54ssUeQXoT1SHvuj3ushY0dqE68P2nkdvIqSrY5+dMW/AizC
wEIg31EOkj/h8s1upSaOBWF8ExEhWNdSX9HuzJ7A6xBQh6UXiZXpR4jl04oYuLTe
PIA2RxdTPA5SRJ8ktnzt9vOM8rAH/z4xhhall4qNUc8FyEfGlmmXpfKYBF+yoLn6
gvTiVKryY1hj2s327plohrJVva8ttVsFC2cF5h9JozsoR8/qJ/lKHdrMDaHlXMfe
n0MFQsnrr/Zo+O4KMltBmC8s6v78Ro8rzzJGZ2QCNpzMzUk4p3Kpwo+K2vtnGE/e
FFGyOZHkCkaOpo0mbHGOUWlfc0sqUfItVkDM7vRgjJqlw9oQni1InGgY5WqZujyO
/PEe/xCXWZlWNbu6ARJ1YergMf5x2l+dPndcc5dgujgiYpyJdQfe0XIR8kLZVeik
GhlWhX6KOAH0QR2r/1caHw+hmCuB55CpqFqtwF/xToqBMipUTl4aeFVO8eT81OLD
NmVUzcl8oKJnq4SwVFV1b37kQdSkSQY+KbYYAImtyevvhAbOBiIlSej/XHWy0lbo
fXvp3sUBwpIJHZCOi1W8i0zju64NbvH6QD+MxmkvvMbaozZg9SJIrm0hN89cuivQ
PHBXXDu2zSA99J87MrYwI+kgMnUApQnGWe/aW5Mq83qcWzb70cANxBhEKTKyQlqU
oX0kO8f8YYW+t5hWsIG3tAk3R/oiNRFtecKzLMoYlD3POw0ctjTxuyozIc5WxUSE
gOqUUqI2xzL8E7tXtsc7t/0ymdoGO+FY/lhZMVfGFf/+kkpIeOX0e+iK7kPtBUM4
JcStsUFQHYga/Cj818S+vyeOIkcuukCxQrYbxFQcDoVIu6Y6IsOTzZxv/Y9qKnex
FQ43oL7fwCEvBtk6ud3eTfl6p/NjlseU6SP0TyiMexx5kLufbSBZTbALu0Lp2efv
jVQ/SQkBwm0zz/BP8Mm/e7BN/4gKJj7lyAHj6xkQ/Qn/2BDSs9NMv2ip6v26/Xi4
4JOXUu7Nvfuk2E9ipDepn0yB//8fkym3OP/YckQ3jTsZHHC3crilopVA3gN0BzTJ
fu0ZZTrqI1iRdmvm4Le4FhIBxawS1xT7xtw7QdShAqHcvbZxVOo+l7C9iPLU7QVA
q+C/T32dSJYuNve0rYqWda3I7O/WAlQml1cEGuCFUzok6IN2qnTdhKrjsrlaahFN
N7hKe4pAqbo54x1iZk4k8GZUPMptbGa4hC0T+SPa8m9zUItKs0fusaIwirrYHPfd
1A8kxIOGx5zXoCvLjxngY9Bmf7xnWjZ6PdvCrMXEB1N+AoCtEyGw7V57mCw1i8cP
IsMIERsDFVZXle0BKWUfa/1S9INikRAVBSTFD6A3gMH7r5BDspoQWfntnqkMptHj
AN20l+hbeyrRadrvkaLtODJZcIHi0WLpGuol7CMIy7/uUfJLq/FB31sl+QKdJHMq
RTwIW/L8W0pwmEtvf3L+t3fABkHUP5rCOpiWG/Ynuoq579ggSiLxlBu5D/XujQjI
WO4xPTFj+VoDZ8nCjuCgAx8m+G7rejlX0BjZDxkdK0M4TcVqE8dF9ooshBhLZI00
qYoxt4r84HdBNd15s+kz78vv5mmS8vgXQFHqZ+Vjm3ClZlH5gcqF070cvnox7/FZ
W+PzyN+w9pMhNrU34OHi/t+thIFYskI7EIJfbcYRaYrLIZOsXSnSSmFBLh8bh7I7
DVj2ZOlQ5KpDDAQukXE0znq4TjM9gDsy2lv5HxHK3EQTsiTn/ebMkxHriybufStK
3grQvhpQhl5C4mSNCwhay69LvDzdC13jPW4SmjYUL+TsKx/iDjgtsA/zs7Kmu1ZK
ov+agiSUUtyqkt+y9IGRGxUKlTNhaAvQUOCPytQtCBjb9FXaU6jfi5mwDGNoKP4f
BxG8KMjDmn0OTxl/hXeGIGR5iMFaBlv+CCjwEonYcgfG1TrNaC2xW3GAvcZyHNJR
+7RMuxSpvcbwiY5H2y5EfOiStlczEr4KRF1Yr6Zk4/1/qvr55XUU2w+ekQUYtc/4
A8s/G/rwCJSPauOYxJSE+Js+a0w1e/GXvmLWUKklAnI6nrcOaDeUw9NPm2EST8FJ
rzC5dLiwE5zT1Xxo+5Ml1qPE43SRZf5BFELH1AAT3m8Vf+NZye2l9e79fyaxMF4p
VXN8YQS9ygL4SfYBbvfjooYLCl3R5gJgTFwDM3FCXrqMIPwmPpLmOc9K6QCN1LpU
sZz7q3EhNCvOkVQMAjUEClvvp53xZL/acDUemfTr1K/5SumQdhrrI4Lo9SFRsgPm
n+4CySvrvavGquHSKLsgPzd89FzEoejXNYA0kJ9Tf5+pxF6EOn8CViw/iZC6mgto
AYgveHoudJMT5G65Mwdyr5Isg/APvV9jmu8Vvz6pIfoYiGgNtgngCDej4TyzVsn2
L7n/b4Xs5mTlUeXbQvqpVxLGNGG4ghabBbygRNWXOb/TP0u/OWBXHiyoQvY6Rs7A
ZO+PYfqsYC0Vp+c+6q5vDUTxmKPB2lYpQQS7iF9omvJSdcDQCKXfD5mFVyZ1BWp3
EZMVviTTbSTXq+RFxfDhEilKFJo+JB6GmvmMh4ERVmMrJ5OFnj3CrTmwmNr1rBpc
X7OXvaqtKvgjy4oHbe9gz2lAIaCPvAbNoaSPqN0/ytdyBLZ8bJpqSuhPFWsZQD8d
t8rlYLHwqKqrwPgCE3iTekyGZ2JHg5uvCXBG2+S235GU/G4iFetZiO3ZgFWIQ1ZX
F6nVs/NDmCV70+3jCLXD4NHgUx+LUZFnzCEz6gB4fZ0ZE5/yi/ONAS0H+9CoLqa5
hdcnuNhJZ0NT1Wj5m55qwia4kfQnPbghX5E4d+wEWSbxa8CggzWqu/Z7sc3T5BMp
IrgaZ0vh1komSOqqCGA26CMHIPa/8o+QMdrDVNtl0I1e05d2oJiTbcO5h8fFb0OJ
1CozMLyvdmgnjt5Ma3FlnDA6CoXCHZdDbwMMa5fAStfYbYBQVlbDS0oo6ak2uKws
aT5YAqY9vQ6Ob7O2MdhZKufjx7ClZlHNmkE6t4n0rSu/tCQ0bYY18rZF34qrS7Wg
HZsjASQDe+BNhMw3g7I4BuWHD4L3ii/wKgM192Fe/Wu8M3QUjGjmb6Gn2UemdVQO
/YBVf/yDoARhquUdfUztiA8sBBzAAcpd6j04PSw3bDy/zctwFd43z9ii+DjeQMx+
lv49kWkpbVVRRX7GjrvDYj2T2OJyTWs0qrlA0JPme+C5Z4vb0Uk4X2p4bW7y6qoS
VoQhVV7n6SVUtjhlR3zgzS+4dz7hHDadChYL0euYyejxQGB/a7zvlIK2Vf4erIml
TlDY8RbiV/9ZC521W68YnVUZKRUIh1Z6OIWHeyuEzrlrST5iWxrZKo8BToysQPYi
vvV2f7VZhwDl08Yumk0U+/XrvN5WZD3rRxltFTW1PjvvRAyDlGU5m/HGWT35t6sC
0tknApn3PEi5pIYqqZR0157WLx00Rn0Tq/vNQrn39e0XufjQwK9C2Z1fdX040PM0
yGHIwBwvVyPPtaJ1QUDGp1PasfZ9CJoNaOq+OBs9xYuaAqLJvzdfts/y9riVfgC2
o6qBhAMqp3Lod4NIKClNqy3c3NqNOD5V6G7pAF/AmW4fE9NHkMwnnBS/X6XchvuO
SFW+EkraHjTNsvpVi3dqs1L8GKARa8Rt7cGmVNyy6LLqgXEOi+RBLYqfk07txQmg
kA/JzTOYBfVcMMIyTT4R1OCC2IDRPPMSnVO2sfInciNHMDQoMCiPV9Gl/fOIZViM
F3HDVc0nc5loS0gjv9HFXCmhSMwlLmAVL6iNRb9Lk2ll24cAY0TKmQbsFTH4/oiD
XB7Stie52scovjx4eF2J7yq7E94SEsqroM/udaiOBVClPuySyMkPQaGmlmvIOgDn
Aa0/zmnOGColLrIPb7wiAiYkyPqmVD9tFWHCu7jLXmXoAVbuyLWlQn0Pa2rW8/ol
vtyuglKfeB7+xNx//qIRlGw+zHxqeMxhfaDQcwulbxE58eTAMDQ6ZmKtAb6u2m0B
9UccLv2PNt8khp8abxkujcy8wWx8hMQPwkwTLFQGS74DRSGrb/YRF1K7qxj+/NaA
etOd7AK/xUtSoKQdNOHOwXCKPtN5m3r2gBSXuJZ7hlktmbur+glpgsxGmxCZiPfa
4eSppwWmDoFt5hdS5DB848TKBFzeFTj1MNvRzJalLNSRbQXdZRu6JRmE6Q+EWTr1
ZZ4kWbdM1hkv/rKKFPZKqhdvuCyDRnvK8t+AcjN3RjENcVT0o5WGpgBriCBijQp2
kHlHdfFpBJttwQmbR1QyAPMtEUB9XjbfJQIHldIjgm0YuabWRfNXaQwOz8oziEr3
1Net8dOPZgYJVy8usxNv4BlLjO0WhpLkaE1JrtfpNDiXgThKkZ6q9A2g1wF6fqLT
+C8SwsS2tkcHhYfGt5eS2xvMDNHzuxnIZG1lIekDxmNMefEG63LjdBdFiRB/yQLE
xwnzl5LzbrxvHBdoJm+Y5BEtiOOQkj0lElCMGJGblCYnHhYHKBgikyzCUPMc8hCH
feGUjbz2OMEVOOZ325E5APrPCmdlBqjnF+QwoWJ+l7Fg+dPScpqN3/hGr1tPzpPz
oMm9U19yAq5orc5UWPtnKjv5+dnJtsmpFh29371WoKlug4HbZQ+1/eHDllJbfPlZ
zs7OJC0jHAkulEG3P6QmoqiXbXyPF7U6AQ4lVbSBiIdSQs7vPU8ROasdquknBnB4
UnaMWjvRo6k3u8n+vWAjr6tqO16MB5e6qMtJCF7k7QRtI4oW58ttcPhce1TNY1Lb
as19mTIofMB1FI9DOn4iOf6ogDwMQK3Mi4LHVpQTtuGXKZI1F+FGXxhdOrrAUSEi
LqrVXe97YQdXBiWF9tAwMzokHPrlSUymL8RMfDeSqqjfk7pHG5EPrtsxHF2peaEp
MuYLc1p0IfB+IDrE+FiIoBlrzkwYwQubofb8SHVmNX2oEfNOTvzcPdBKWWdiZ1gn
BquwzF1TWqn1ojot46nsbufurrglxvWyeZjyDufCp1glf5ccTZ+9mGtkpdg5fct0
A7tNC8HN3RPpZxsBAGeVgvQrrfsRgO1//Qzpxj3eSAx9TZZOISN52pMYEJqR8zJ+
p1HX85AqmMq414ukNbwK6yoJtbltaa/O4B8RHuSzH2XcIKSCqgog3joO1n5w5eu+
9ocIJqspyILdhB2nmSC8/n6xT2HcQ6cJqAbJ1iyqnic7byPJQEzEUjqTR46nsS24
QkSlO3F28Sn/C28adN2B4eeDuMqTQdteZMqXzRVjuK0ieEv48l+z7yc0/rJmdxEk
NfYFQ1zJpT5A97uGOHjxj5GPDbljouhEPHmItJDeyPt0EFJVEdS08wZ4URqOqcy+
Jt4LiHDXxPKA6qdtIzcwc/5A57KbXQfnjqNeOFPXz9J7LEGhJAIkQwQTpNkNZLf7
k4yAQiJmbe6ThVFEIB5DpUU8bTzt/m4vdfTbBVM7OyTHFs9+HxF6PE4AoOc5Aoos
aFRd4ujGgMfCoxoUg9iUXRTli6PsxZtgPy9WcKTgs9m+ziUBrZRmdccFhcR8mr+3
jmcfX07r/FvPvlUvjQ/J6pWFFSwewkta391gn7EaD1p55bXKfuR18mtAg1JDTXVA
FRlWEZ6w4bXMBRufX/Da22Qa4yqdo/bDmTTOakU+KpA0hceRPoCLlh9hkijIQzbn
raita4W91ZldLB696Os1EV5Y9bEI6C+4mZ6UFpBtIXAf9oF/LtZL+wZ6Ff9RDPnl
7ctyiFdNcVsCHq+k2w/YHs2Evj/mn8b85pyo2D7gQSq5G7iKZIWhnqdUTrYtq+4V
37UHGL1vJgiifEBwyjQikc7YrAYFahSh6+T984cgOGlr+c3LT+THvoxFt6CLOXK/
vDl6oAASIu0LZ9NtlkPAPgOfuqtEA+8ALEL8ptxu+n2L6gEtdEu/sPD4ExTiRbal
CD9bbTuTTrkZzWCijMQom4Dy+90mLMHrPDrbEGM13kFPBqMx8zUf2KO2n1njr94Z
q4BacEHanIQRYkkIYNxqGV4dHE3ImN68FhqBAYP01N61o0lS1zSzUGx3J1LHFCfl
jWxJBjM6fUuERdjmtkneCzHKmKNxxQnjIhdmX5YDd9kwnYxw3g26QBXN7vaCHmOj
vZfKUHdW/IuQRdQyDN6qZSIw9MgB7z0delX4H0yXOMk/FEmDG40evOpJ08PTiPbU
yoUZfnV0dVkvF6ezJBNQ/8W+nEQn2b/Zd68nI1iJT/DWZQ7fxRWg6XUo3365IqvU
04pC2CeDr5dA+y2moYpiDi5mMf2HQrkcljq1PO5G8r4lQ1tx8hUE9LRx6wsLttJz
rST/sRqllVpZ0LhCV0wQYPj8w47/DIkWs9nPTh0BWv8EqbwSkPknivxEV9ixWcdz
uN58RBVYrtziFy+JCYxRJXvS5fkkrIrFcrjPrU0UUq/PiBiYh9KCPCRSsI/gQO72
fDWmJCWebDHPgUVaDp2oSyyMnkG7RjQ793WCxoFQe6PyfZhkBGI221ja3OPPEjkV
5oHsaWqNzPqQ4s04zyDIGwpDGS8viRxJ+1CBdD2hQfrGrflaj+JHjpwqJrdeO9Vb
9tp20NdfYsmGxitEsQIjnZKFfuZASp0v8h6Y7ZrFnqCJISiqvcd8yajLF5x9Ja+V
Lgz6wrJkOPohPLcrfv1KtyFtI/e0QoKtvOCKbTiB7aR3pxkNorHmE3rOGpXlLiFg
0cBOq8gHho4H7OJMuYxZawsYjT3Js+a1hOO/bL+SjuQEV3CtmQYTWCkAVl+obC1Y
fegyT7yXJ1jbGk92bgQdA59Lg9N6eXGn/NVROcxg+j+s0DeVO38/TFUW1of1jDGu
JJWEmyFdcgtFVomiXLwBEc+oZY1MQGmypxoodZPKRCjZGAtGu92Nl6qB2vkwAbm7
3Zq115uNiZ5G75+0KigIs+Sg2fvO1PvPeOApSkDcmJAifCdVFkEQ65fZM12SP2Aa
MInnTV+bXqmS0V2nXvtSoKWf1024h54ZtfQAO8RA1OuZPZN3q4Zg8BQw0DYkKDGy
bA+SNwv99KitgWr224xbLstxkHZZM5pdBKrBerQowyrrPiKZwYHPFg//F4eKfS8V
aDM/v7g+gFUITHvUrnrvLBxmH3dTOSIPxV5KyFQtijiL6p2gFG6xKOqSM5zt9M+N
Rp1gAnaTbr6ZSZwY1KAgQnPsJkR77/Yzx8yaRgQHJuQqwInPY+GVQHxh9HVyLdHs
flCUFKORxmGZHCB1UM25xnFjZKRTnaxuNzizDkmVv7YJSJXCYmoDIZSRRU5w9NeU
0bE8HUq2fUKjrTPw2c6RBTs5JN0xqjfswlzvydz4EG0WB1T49TdGc/LRuw9+PVYA
ErLF8NY/isWT3rMYQaACkQwOtuRJTREVZxj074p+kd3GlLf9gm7BrY3FLd1G9KCV
YLgFoCWvr8905kZEfn09C77AwSFhkxAWX3cwl6XN4DOe13AYB4u+DvzZzHVxDg9l
lI4EOIHAAi48Pzo+BOqMKvzR+B8Yrb7n/ksa+HO3dLmedFMueGDQ0GLgvUJ8BCKa
ryB5sq8EFdx7X5xAacAKOZaQcav0Nv6TeHZGtkabf3yspC1xYVZv7CeMiyA7VfMj
38ybCXPCoOo/oklgUUJk5aXQr/TaxCYT171Dfw2deo+GUNWXwdlb45jWpfHO3ZB2
+ZrA2DedWprfHLmnivNuRHc7zHdSiO5u32vchM8cTHTND1cCFi+80lDD4YwK9pWF
dGfnbZKBocBujf1W3CurRAbx+WkuK4L09poeb73kyqOn3VzWq1LBbGfN/EbVefSz
qCrKoF+nkfGHuZaCQs1QDQLkJx2L9Lig2nJ3d57sL3/CV3TuG+RHcTSAT7jkTWuM
gnXLCwMKstXzkrQlLv8Hsx6UOnPilop85+D4JQSABjVB9IgumDhNYnBvNtbN+6Wf
oPaC8w2JeTd4l8o6/XAmm6+Wp4m525sCN8uJj0DWLVvw2ABXZQjgEWuSQ+t+VU8y
8KSTq3coVbySckQ9MoOf7tMNSEZ58mUfVV0GlI4nIImSINt6BuVN+IiTY8zwW2Zk
sxMLbdh2hsPYR5cND3g6ZrRmHy5Fh58FYo78vmmoJ4+qcRbjRl6IqXCM3jEDLCG3
uxQZJg5Gsn6BEfwd5Jp/lg5y6SK63zyMLTQoIvaHBihgmM8Dnqnnsya31/TRWshg
NZlAC69boSjmTSLiyNpySkNRMB57HW0aZp1mz6n/hpYgvj4aWwZiSBl1BjZSK4IW
tYPsPBMqTmHfv470TE1L5JtkyXuWcRpolq3pmJi+2HqsZFkohZMz4uw+JIefKvuj
mJGBiuErbXOIEU9yi5/Zbawk9hmr1EyWMjyeMVIPgJ1fgI90CjnK2fFeHbT36O/z
4++uwWJbXdEPfL+cqtlgxd+rrBx8wf07fi1JMyIAs0/b2PlA+qWpM3SpIq6PhoXb
qi3FkWior2u8M8XHUVtvlIellD98B5TpGFy4888ZV/ChXJDchhjsK2aZZBbRGNl4
OoxxCAIBogyjm2xZxo7Wsjl3OSUw2ohBnZsZn9OqYOCkA9JEvllD7xf6seeznyV1
bknYBnAMCemrVlXqvwpJQWTxxMJ/Kb/LBohrJQ3kBOVmWRaOWdxh42mWG26kCi19
VtsnF/60xfNsPkBcUw8tKBf6oO7cLLjyWKp9Ed0PSyBSAv8rcO1vPQuNwSvUNLrm
U3msadhTEKbRPIuLqwRwWa9PeVxoWPqmDFbHBZRHAH3/q/zYoSMpAVmms/inw5qP
ORaFjlZiM+UaGeBpn6+7+zxPa6J6ca7aXB9ajSimoAwn2bf6Py3nGejAz/S27M2j
XAB8yUQIOAqvGIqBr7t8lR0amP1MA8ymmDxMIy/u21x1mkD4s9HOa7Ui9AlFFtpq
G9N5BcYyUVdta3kX5RBR7svrc6clBE4z/WpZp5wlGBK1X3NkBm/QFspoz11PCsQ6
uK+Hm4yER8yDi7jaKDt2H0otWoTUNFz/ZcRWMSj/aXcrMLLe0NE94FuQIibpM+/v
WhjVgjw/kY6yNniktusHHybpLm1WuC8AZ0Ac2XeghuZGrDZQIhHZjEOmXQB/ov1q
YkSOupid6DlBSvJui5hoODmd9+vbBqbSGezcofh0h0HT4XZfYQ27aRxvSiXjAZcK
85yRhZIC2O7eVNhKphBM9cytN2tgy5Am1v4sCs6xUHfmRsPGYWVF8I9QXy481Ulz
ojJUwcVLgsmCjFbJt7Jy9gMEWFnP9Vh4NtVpUW8l60Or8GcJR2j6zY/V15/yuu31
5tPt00swlhq1kMgHPCE9qZtWEqRHE7E6Jj0fVZGuwgJftxAAN+iRhUSvO3RTqrzt
Twk57VbzFpUMMVhDEt0EuSGwHTBSxJIu0OU4zAR51drAcaKEQL8dif+kVIPCvZyV
Zus4H5U6RwG3RO0o75I9aiw6AeVfrQdfZtnuLQKacqwKNrdQ+wgwKDnDN2LiNU5u
d9CFuhcNX+XAfG6HTfQZPPswBA/DEmBWKRqrQCtc9lc4dTUuQgOiR+1nYg+JxDny
4xBE7mfLuF7xbxATI4tXPTOx5XbV0C8MQ/0RUHX3njRA/KhW3mUhgs0cmneIgqba
235UwejWGIevZQFdcIoG8laam9CvhuG79o+ReB7tiwsLKQ/2k7AmwYtetKK2VzdU
64Y8QZ5Kd7yFpB9P7x+4dnosuKA1r8U5m0J+7CZXDg/3FFekVjPkqJdcQNzjgs8k
jDBYYPm0rhTlJLjqUNAMqczmLYJvSfGkNNPCjfro2wLqgKnHdzUC50Ed/m538kyo
svxeNn19g8+VUD4Rsknq6lqtvussKgcPB350A9SXBlhhv3Z5wojeRA20Dcynf6Tu
csOzYKk8CuXvpagGWMGEDM7e6X5fmqLbdTNjdsV+ZuCwNxwHfe10N/G2ML2uuTAq
E+N/wxseLWHUAvcAJGns4Do6/PPw9cao0HLWFXdLUKrdCMJWDqq6FX2I7mbZdd5i
5HNNUW6+OOXfA4GafBlmlqvzkaC8qa9engIT+xrabYWPCr2pUk6IYCBqclIn66gr
ENxGdqgPL3vAgRYiheJx1S9zsCykK+LvqUfvMj3Bruk5cu05DEt8eRgktc9UzvaR
ATfflBSYBcLJ6VPEO5tqkaku09E0f8Y5cj2JovwboQhd52Y+Of0jx9SLpYp7p+e+
xKBN8mFp+cHIiFUsYrZhVGwOyuAjiRYxDMrdbto8FSRjyIpqmmV3kExwjGJ8Kq0W
TqrbeZrTRTPvxnl9VWM+Ibwg1845zgOCD4HGwiAapai798LK91oAkteryde24eh3
FbSa1W5M3WbTSZ70FIt4bLI/ydTuktXm0P1g5eGGI7Fb5OZlzDdiLtEBWDfEUvD2
7cdNYoR/q+QkNUz6wi5vweXszV0l4KMS2ZRRVAM9x3QdUBiyBLYMkQqIrL2eIof5
MH3YBTgqGuTlIohpSZNHRTNydaXfKLv8On6YCiVEWqVdSEhyKck0Z3N46FWvzx35
4W5RkuDO/zWaIh4rijxCGh1TJqTiEzHM/HNjTcrmax7vaC9hX8Q81kQKHm16Ufnb
KCg0/nhgYlJBjxSfaofUtRjPUoJW6c7alPWPvDDdQLRU7HMEGHbbhTQ3d4fvvS92
o+fNRnyqYpF1WxNYf49z9w3YMaqbfstI+a5+s4odsL7Lj41iCEctgppW784qncEX
UdIIsjmwf4P4UDLCbP6/hUIWt6XhR/J5C9bi6w78eEJbTvkfXZiENjDO9bz3mtsy
3xVl7UD71ibdaSa4owi2mAZquPE8WGfQilu/y4ayMg2R48o3UYO2+6gmT7ID9/08
aXsdQxzIrZ7elJKiISccEl8lQlSS/841zPb++NTmfXz/RejGjaqCQnfGjyGaGi59
nY6BPVRXWNdwe0TRNq2e/L4FuiFe/LNMRWTSDn7jIh9OjDG+xwP9u58tLI1rrPmN
RkZ+rAaOKgq9AuxtXdcctZ9o+DHpMe7tep9En80ko4wBbDpI57pZyMNpBHeO0RGw
TAccaAgAO5w9PCVftCat1nIwqXtXchOos7ED6GyG5wWqf2oBv+gksTbYlj9R8mln
gVQ19zNLLjMn63e7SfEyhUSEdiKvt/CoNonX8VwqWB+X6AIybqdqIkCcGcXjHDu3
/gLdwnL7z2bUge5qBIYZRlmVbQrx1bfndkAViHpx/o3v3zROjMq9t6qm/VyA2nDM
qcDo3ti3rwTk7mheIykFDAeI3snZBO8Fi+Gf8IgpWiKGyhiNZkvKjtwZkF7v1MEY
feXXR9kjh5l0sRPNhFJmYNjximVWcv4k+SeloB90+77KmaM5UYLAKwpNqZs80/BK
RUKNmA/GeTyUVvmWxIkCrNHRQhnRfTp0tYzS/CcD3wodtIFtLd6Ut40mIIrkQr42
8/a4v4+shyiv/avNNw/yAZ/akrqZIxfhp2pVKY2fsj78KXbGyQHn4fyyw1mmfYNJ
LLLdrJGS8J7YAlcTGOIg4PCtSGwr2BhdglShn/zVTUTbfmFWP6HSzKTg0AeSDV/a
Qt133ZqcrdasyJesV0BV/piCtTkKGh5WBG0kpiuuBAY2eP1P7hy5M3f2JfsWeXbn
mDJV9YPHpbuOPvo/fx0iVoF28EXSd3JkdNycArEFv0tAiGUI27Q3vgnnAn+W57/x
+KiylZqC1tgp1310fJMftIgBhvwCSlTMvjALIYgHzpSAeWOyB9eJeHr3dzmfZ7qe
8pXcTbS+bpzGDJPrm8Eqb3KelyyIK00qzCzSRrquSrUiXzNV3pBZflbO//9ENpnB
eMqGZR+RTaejvpN2929xyqgLBwQBDtQh/T/ywixoZ1GpNGcDtbIyJv+XD+VbHgPc
PlU5hYvA18+nooY998NSh6L2yFGE5GvCeim8yIShEofqxKTRF5qv5IJeXfBE0A4M
oEiIoloBQNNR1W2e6osN8LaPw1TJnGb6al2hclclvVRZguA3gWb28Urc9O+j7zNn
74pcxN9g6qUt9D44KpmNPt+tARd3JAH0NZq2rz9YShtuyOD+0KZQrBPbVHir7AiQ
IkJzPdFo/qGBZUwfpIwgvTIH6X1bD1SfvrcSSAiJzxp/CkxIj4rLxKM1TdZ8O5fu
EZ9+Qf/vwu/fV2gkeqjeehScDPglkuh+6R08YMxO6cpckc/fF9SQVGEdNizdoUSw
O7XwUHUUfDKtf3tS8hJNa2hEIjou7t/KSe3rAhVz8EP/IP1gRwvqi3vm0dWYJeoX
xzgXYoDG0J8LNCNA42UoaQskjzRNo+MeU20g62wiDdC5fOn5hGk4TGNxVL7qkMuQ
MXERW9qyMjra6HgwInzeR053Rx6VaAPuJAIZfHRL5gFsHRAGYj6U6pNv3eGiInsp
5oIkR22t/E9Wa/vHExi3Tw8x9H4KU3+NxufpKG+tq/luQR6ZcfUhhnT7EfLrTcJR
wxD76XeMug3Dfrt5gkQK/okLhXzpe3ShDbsuINxcz83C3NpwR/V+M6nLq3UoAhAz
qNjLDggZqtFOmk2aZcbiNIZLhAER5fg+UNSEZRsNoArJMWYyQzOyITuOT85miwVe
lxG3G9CqSS3ZQhd+laJEf6rlabMWB4PdFwyYcIx75wQnpDG7v0tpFGvO7XprBZ6Y
mmoWy9Sn9tUYEXfEdZsxsGVKgB7VGbFXMCWBz1IaI7qPNXOoy8rHgZ+60H7UkdTP
hdqTAVATj4aH7B9zYqHODGgsbsC0lFVF+Y9w0Q9Y7M3gJSB0xL3TtU7XK9Aus0Ek
feHcIRLjMn3NI+4dMC3I1fbdsp1UMgPSBhA052npoATh91vljX0OpE4m8IyiIwIW
A2ZF6pepagsz4BpBWi2Uh4y5VKqNGM+G6uaqMZOF2apPMirJb6YzU9sw0B5fLBl9
8kuP+MUa44A1rvqbdmceXNnCb3ke4Mw1ZHJm+P8LsODVJaZPK+eI+zn/N9H8no9Y
in+g4jO9so3Y2qAxVAHYfA2fKv6vmBYAELvNfjKzUBdxGpbqnQwFDStLLr+2cceh
bY6LmUac3hOKZYbayPvCl2lJ4FdPG2WNdTfCsxymN2ddAMLsdmPQFJa646xQ5JHR
TZIYaubKLcARANX0Vn8fHgmRtylGAlEKo3Y7AKldZeRS8KCw03wdACcjBU9FKQyi
DrqN4QpRIa5Ga3ixCcXucjqxL7z3vOj3QVxOmnr8JxyG+pBl6XG0CjIrtpgQ3ne1
fAextNIfwNbGtfXIjZTGEpAE0r/ed2WBRZ61tjJTSOoV3cWZnJ5+s5Y2hc34A3Jk
HainTSBXUjyvj6aBj9bH3buJBxcKPZ+y+SlY/VAy7sZQH0/4y/Jw+UcsjKQjVYAo
YHuEwrakYvM/bKtv3kX3Uh++Q8gQwTi9sFzC095mJ64BvC1cYrXq5qCfbqkcDG4G
wwk/iIleDk5SptyuCVk2dAiKMEftR7s5/7eSZ3xnrTqAP6sm1WPVda/yzlhiskZE
ZxPqs0RuBkx6bvsnMyJ+Ev/Tp+eGSakicIBT2pwQDkECnIoNKjuVfzzy50AOlJiO
sC4uELcUrOYz3uSDKLheGY8XVshZxUq5AVcBM4YAJgMRhbBPg0c9xdiZuchZ31mk
J8QCZhdlG0Db7KEzFebNjS6Lj6FC5xFKTgQDRpbXHA8kt/E/fgM4ZbMNVeqY6WYJ
uSi13C3NPfVv7wohNVTAlhpSEx98I7SyDtXz/Zs2LQZKEdEJZ5ZwEeQshQrevVwb
LKOQw5tNI4mEb9WNTNh5oJrZ+f4MTaItqCB6t2jGIOHaFHSkd53KAxncc60yK7QD
uCB6Zd6b9u46D90sD5P4T3BuADUvBWXsC+JtfgRzstVBLn53buT2HamiC95CPUB7
dtSN3gm0TmmWEdr2NE4R+8F/ta0dvYh0oJFIt8HwrYIF4yH08DNLb6YWfui84+Z8
NZQq59PpN9A/0rQJQuSo/g9qFFepA7QIXV6S9rW2iQixZwLT8hQreZxV5udWzZ6O
vrAM77Rq4TaMuge3ELNNdO02t2+prRbdehihRxb7oGmKdn2JlUCy8Hu0KuARDna8
FNgGHnaMJpDbZ63ylsclUKoWXCSMa8qZqVZjvOxsYwyVgJaqgHBTRN46+MVMeycB
Wl5vY0L1sTLQ8Q2tVad4HvQJqWb1So++hQsWWcRA5AfvTWP/lwchFE0gxNUcIlkE
KSamJkbGlY9sR0XE07IKyx9VBqKQNtnjaJqVmPPJWxPaDLBpet0Mk7m2WEoRDEh2
Zgj2ijHMUnaQDV6U55M5xeRtnIJuCgIAID3L3snseFIdgultj8Undj+TuejknRde
XLGidV56J8bcI2UaLy0lRxSR70Al8KyvRl6J/MoE2726CdXggp5eNKzwDXZecZnA
f6eht5RvtqaY77IjOHv1oB4Ly5na5WpLRriH3d5SrDmz9B0VwKPNtVy9+Z18Ciwa
bGBbe4iTNQElm4NocYSBOs8NKFKpv9/2IphFZRN5t4ejHeO/y5wCPS8X5Yw13yRf
uWu2mxjR9U2WpegKmDZFss8bNA78yEWpy5ChPh14T9axULHoqrtm3jrh2RTTTxaW
qm0qFlmEObNH3rAzfZIPFUtEacxWzpSl3KMNwLtpz2APVjzKwpNdiRSI+gMQWsl7
XOs3AY3y8Br6NnuSQW5+APaViRBuD0O1xndzcGpO85pR38NA6ajuezDhj25mDDXs
aNSGW/fvoSrsIu1fT1aP0oh5HtkCm6gb56PX7eRREJmrHiQJMb0C5QtwDTQz30fc
aY7PEIBhj1AvtO6XEv/SnvHsWIobRWn4xzUweEfRwgFmRPs4AIslYLbf+769mkxL
09zStuYcbgG5HFEKDY8y5F4tiP2vqeB0vDrwpxydVMxsAdblNsUNwAdmhmCZZ+Is
mUnRJi2HoPuoXZdX1gcGvswUDxRLwmUvtErs8kZEozJdB6kHfETxIDx6Dnch0U46
Jz5H9WrrAo4xfQAR5mYs8VZVOcox/ZN6+q/Crybgr0y7jKypxNiYEwW83cctaDq9
lb7T8PImR5VS7FKRXFvuXmpyvvQ0ndIBH0B5wQi5/kh4n60SkWtlCLmyM8n843FY
I3WLmErcOHB5NYZS02wQ8K64VetOXjVF1Oz5wM56BzLfUekb3hREwDDqAd6Jd7kj
o1UT2cLubNJ3KpOyKhhOHe2GzTFvti3M0M3yUp1iUGDlhJLpy2rK+iaESHgXgI0C
wn3mOUSkLBoM4CuUxZ4jm1JocFXWBcT3D9VewydTxT4Kep7Tdr1SYwb8HYTIGNej
BrGXgMBuUMkiPxPIWYVKe+lPDGjG6tAwpjvVyNjqFqPK99m7w8US2mnsFI26/VtK
zwmqiA61XOWQpe+pqO62i6+BI0+F8FLWDixQqeeUHaRB4JKALSSa2PAfbso0Zh0M
VzBHheMoaXFCdgKmSlBrtL8YmE9ybTv0ttsNo9xkPq1VSUaf+EOLTi9ZyNaQxi2X
jLHHHEWIVXxU9v4GDPSHOHT2T8HkhbhRdQ9We6eE8up/iOHncolq3r2Hlr0kSo3E
Xc354O7x8yAca8+TNsMSZdT9Mt0xzTCDmhoi7924JxHxcVz34fJ2yiE/Y9FXtwWI
dsC5sBdZHfOGrL3X0xFh5Unos1qKNg7Aiawyzcz1QbRVtzx+DSOwzraw4KIr7Jef
OxCIrw63xHY3FDmdcSJt5r5sicqKwICpaR6XglIlLIuns5hsUQc+5+3I6d872vrF
zZgVkhzHiuRIzdAUFK2h4g+WRMcTo3LNdUoq5plJTf5pNHei4YdKd7C/1JWmERaL
vQfGfl8vfk3lOcR1SreklzGauQeSmE/Joy5a58Mm+M1uw8zq8MFmFU8nWsnMPND5
yH6mEsjRSLG4Xsnplom/DTO1skKQ6PJnNzWSnKumw88TDaUDmTQo0/TVfXUwSDvF
NradOABt/5+l43jQYF2VioURfLo/JxN1CGDVn1yp9YILBsfinuHHGTjRdD4iZqx7
VW0ePK3pL9F2D37KR4+jyIQKhDeJY+DtqqlevQ3n749UCozL2Fcim9Tad8LG2BvM
t56GWShrGnO04rykGXGo2I2nqyEen0DKLZGmjtdQ6Mt223sIgtAvVD7ycbHEqSFX
FwTv8q3PyBoodRBLOFQaXbanF4gCJiT4+yCPNBpiHoTkgClY9vvcEXnVyksjQFUj
0vQiqFDxDayTF9zBVyAvpyOn+Rno7WGl33wCNZnrh74APtGcC8YjBSPazdwSzo9+
7kn2I8HKABI2VCGHM6w+TBtX1wlEnqjCJcnuIBk/IDew2Cp4zHeZVW5TiucvD7E/
T/zWF0YHF3b1RRn6HOmv6PJYK0V0yL6V2VFf05jC0ZZEzjRDgV1gi6opRrXIEH1s
Kfeld6zBetMVqESduBX0s3HD4Cy5SiHMhTfUvy3yHlOi9Cy1C52rSEhbKkEqEiAe
3lkOfS+yTR+YcMnHwhTjVcZKg2gq09t16l3BQ4yT+WeQUzF/WLZHKkdKxu0g1Fkg
Ctsc13tHgA2OypxHq5Nvz4oFLz2H1YHtTaCgThMiKWyZEdSsSsFJOaj6Sai9Io/R
MSNQi9eGbo6ZRxeo46t0HZhEBRUnVZnP79uay9kM/r3ss31derVl5rT3D9yDe7Zk
pGJvMWjqSMXjZncYV+MLf7XpF6ZuRU9wzrfP7BRVuJPjlPevO0dkfUkcY9FzojKC
CzgBjzz9T38BNJxc3cvZo+5FPY5EvYpcD+oC9YM6hgJz4YhwT4tuljPI6Xm0TnPH
QS5m9zi6TX6cCw333mICbPZFaOkA33oAXAOdC1JkGSfQuEqzUebmOgnCXcuFQ2la
pYATRq7O5MAmofI4pf+eYzdbz9Y32AU8hmCV8O1P6DKnk/gNgeLVNDfnuxTHhKoH
RVI+5o8aJplrVKDabT1Yigd5N/OVG92qYoA8Y2EWjIG7SkDzFb5Hm2eer0uSsaIA
10AZBGdPfh3HaA8MLBKbNXEUTn84cUfndwqOsqVpN2H3hF5A7+JJ6trrFzY0nVbn
kKXUxwsHBrMr5hb/lXFHU4GG4pykpMMi8Lv/znzDKIIX0UcoCGV5ubHIRoh8aLzJ
4qDxEuLd+7tgJcxZntXgG+GfMIamOFzky9h8bye0Ei/Oxyd0O4D7PEkWLwtFhBBg
5cnK2NrCOG9Ux2K3WeJBjhf9oRVouxcZ3nCLbEES6jFebpC+/J29X7eQDT4rFv1x
mtb2Z4i9uH62GkLIxEcVFKjA0ZR5ugmSXI5bVZP4TBNNk1IqgsiSHf2CyB26V0mN
J58L1EtxFFi6HzOC+wsfZqxq2U+kGw652W4CsOrTBwNWvkGn+oNL5lNbn1hGmDgg
b1nRNh5eTRIa6S8FdE2D8dgXwHLtOaLOQ/Sk0MjngcYVbM8uw547e2CSOJwxkv1A
up9+3G4phrWY+5T/0WhUWQsU7NAeSKq7Uk6Auk5Eh0wKdBEPu9FrHo/UDhY68aen
wd7aaRvJXYYOd30FOkyCYH+H8DNutRR9Fxb5EUeW8aCDW3a73Bh4pwrCaJouZXqu
EbBGpbI5z72McZUjN6bJT4XIYrOpOFO0K6dmv9HRhnHQBfXcfKWbglg2I9dNNn7F
B4gdOSyjBQbcbiEH2fmcwWPbHWWs4O6jWZTjkePPvB8O4hfdHGLaypyTwVdnFFLs
oD/esbtg1ORrHv2akbhFldwVGNwljaDc49V2Hza0wxr0qITmNi27zMoNQVq03klA
rVeDmhm0iNXrtmI3gJGIDd7Ys/LNUgLBa/U8+AEc/lxxPhHYZQJ1Jv7CyPWizSgH
gzNpGmyVEOODLrgL6mypuzg2kDFZT6vVGopB968CtbPG2MPv5x5EwO9rVRlauLPT
wMeYowLO/NDX7YY4rZ9xqWI5QyMbphY/VJScN1RAncCMsbTmG19pWy6t10vjdCPm
QzSoJ01s17MB9Ux7vqR0qHaiJ5PjN7z7kdvGyjWXaFwunn0UY/BiYu8guXCU+WYf
+UsGCft5XmOEh53BMLQ+weRsbGD5SYfjaz1MdvWLfXyZBjgOemAk3ZudGN5dc3Zr
Ts3bb+yKsC2MaeqGZ9sNOPsIqtXwfjNHm9PuS30YnmACrwc7mARg+u0K5P81MAqd
TO1daUEWyw7wclOUnze3ef0DAL9mmm2qTk12NavNlm2itcHFcMH9uedKEp3ZPk0F
ed7jB4QZOeTHMlt7VsVvwlsyYVONTi/R3/f5FwVddIDIxrDXR6VBrtkN4/a2x8Oh
CTs0G6h4bLeGkQXaIaEtw5V3vuk925jj6MD3+gav18ctF0bvxDZF5aaGm0HC928r
QZLZr7mPzqlD4Na83TfYAU9tsTdVa//OHyxiG9LL8bHNldWo9WzRyEqbkuHzh4z1
R/bAjiN0IgkJej+mEBDDQchityuAaHRhwWSy3veTo87mVL4qwYaWYfVI4cD4WNTL
6sebKTetECBrLPTVRtInEGxyRR5Zh5iY8gQm0FH6h/57ghrkUts6Tnl2emXBkp0S
Xol+Du/rYpYEwf7oLojf2IO5C0Q7OUFBiJf9pik1HFlSQfK9Ojc9pg2KkiwOXDik
BGk5Ouscugbfj4lQmbqXRqoKT3cdU3iOi3n8BXW4Qd1tKvSDHykCh+0xEIOAnS2o
nolaF5JsEwOK4YK/g7CqL8SrOWzwzhbOaRgfan3Ep+PxyRUrT2ICwhdCEdWn9OI6
eUtLnfzJSGzCoRWAc4fTilKZRUqQTb4d8VNOMg97UIXBKJzhR1vRTrQ/WOx6I0bB
epIkAz3DK0CsmwD1PU93vbGTc4EcUpZ6TwjkDmOE4doUe/wpRiesVOo+8SWjsowC
/0EXum2W4Ddp4m7nrQKZhoNCyk4GJ+1fdSJJaGP0Hl4JX2pjil2jYzzj3SO2Oq0s
Ub80Nq4Q1U+2kixvn/245weAlTPOko6txBf3NFg3Yf7KpU91iHhHf92iEv9/gMBx
GiboSaxJ5p7WinytIT6DQuwWU4wz5tR26tvmVl0/aZ+kGMUBqfGaulRsqB1r9Iq1
OMGVxZHbDy5TWxeiMfQfIZWt1wqkMGpcXMhD0HClpYUd5zSNXXUZ0SNcs6VLEKr1
oZxkCGssTq2mHBQxIAlJxMIh1SPYc+KsoC/jabmFEX71UcRWiv43CeICJsSvZLE+
9PYa+xq/TjCVOsfvTuBUA85gXMDT/K+LYV1fl9d+C+hAUQ41mXIUxwkqeGeiL2VR
Z6pQVJv8pUcjyx5BqbXehGCd6jzC3E7ActbeeHRPYn0aGkq7R4QKupsTOS4vqF+3
Azi3UUzOBzJwzbRP3LXZC3wlLT1sVjNnVd0JBkyJbE+mj7bJhY+ABJe9+tBqcaHc
PqreL/UTghajZ1trrRlnX8Evd3fcgwaXVuCsJSKxpTtpj8XOninsl1v38LQxpFHh
LsvdwNC3C55+sg9EHf4ouHtZoFASgxKDpW42TiGyrm88Z1kQKGqim/tk3XNQRR3y
sP5QoYqRLUPbZPkHEI/J00QHVkghGH6QhnzZsuFmYDzpJFOuBRyZFRTOGiaHGwk0
iw9Xj8GRl057HQqZlRocOZ9Sy2r6xIsqYzmp0BX2Iru6FSDgRrFQ6Kms+iBBAwTt
3p+pKLDye64qv89QMcsckBk5ZLri4NjkmHKQnnFHSFAzO2LZowmGY5qITvHghA3b
rsHFtA8XzvMiUGpkSYGbipjvwLHnyZTHpsMglogUqZ1UuuB41RhyRrWu2wUnTvhK
AhkDuCz8Dleuo9G0jP4GIunPJ/sjK9MIVSkCWjLMPy4FNZugXvJAVKO5ql+R+d0R
v7ETSTb1/k3qkeORA4YBys8vlfXKR42TH2yJB5ElaPzgEpyVSOAFXkjYLEPqmwpD
YRU4XR45yz8y2aGRRU/hGGDniwt+oCa7TBkDz9QzQkX+kieVPXps9ggO8ED03Jom
nLFOc2or03ALTBOTn6rX4qrq393G5a/YW2iFqtplfF3qkCsCcYIELCnm2JlmbeCI
/6sd9iGl6iLdAJVA4XzNaDFEsv0zEsRsdm4tWEPx7NDlg6B+fSR3N0pL0VUtaX9t
JndYGUpbLlc01s7XNTVsIhiqBPrk8uXsjtGCFxZiyCshGxbqzcgscyiyZxhGZu4j
fo6DcaM0fIckxLM9yfyEHhWHlzr7VsQ8hjZWOATqRhKpzJfRAZhVJ/tKD3qvT6ks
BtRv7NqEKfRBE8gOKZGVduv+Sh7iVxDxqpZyjXpHTwmGLuCZsa/eCpdkj+gLsXKC
6LyfCSffxX6sRHnxjr4AZLBosteSjgEwBI1W+bcLnzT2o0TCuEdlqOqelTvCrxmG
+zXbgs915sVFLIxo1d5auW7yGSbOs5yT1A5mcKkD6bpCLfgxyzXjf6CBXoE+Lf8P
TORiX/AMhiboVCVj4vCn5Jte3YZrucoOfeY0BQz01HqYXRn3jL5GiFQOrwc4uyTw
OfMnqL6cTSWkNkE6XeEZgoHvOmI1mgfrTrF9OYrhMXeOHM+48elZF/Rt7n5+AItH
AY75h8e/e78UI5lmXMo5IBkzBkkNxZcp39Z3iErIIuKN+hcXlKT055J5oxQhUgYC
hm3zxP8wZYd0eIwlcqhLZMToAh9uP89poxI2UoR1KTH2QxgNXldQTDpaCHf9v5Ox
xFKdLdCZXBTvEMjbcppbvgLvVmJW7zlaUrd3bdzlRzw9meGRJVguJ5744IBC2oXz
uBDrvcbmHmlSI76er9L2JkursYyrWG2Vyz5MGiElDoHviDHNVHrXxnMbkj6Jww+O
QLJ+VZxnLjGXoGL+aM4oFjxEryJmqh7aCwfVAcRJza6ng2h8/M1sBeQkgYYmEqMA
7VYKx69tnwfHkh/LOlUV005MDsctqu4zR9eC2moqnCWPxjWISFTPH1zKmmJ8BIHc
Hcmo208LUSPWmWuKrbPAzyxEqUlGcdrm16GqCHQ6cU7Uaivg9zI/nhaNAp0iSXR8
G7eg1w4U1J2a0PLAfKzv7bgsZ9qpdi8aBgMuJdCWEZsW1WKZm9qX73+PJzjBUhDk
WQsIlgsIralcnQwo6dfiOAOj756kXoaoHpGeAYYs44Pktuc3KXaW0TwpX/A1zbTV
+owXKJ8ae1dVP4VW3OMCDsDU2DstK8ZUzptNW3cfv7BWeAoQ3QTpyn2x9KtoD16K
CUkW03NLLv7dmE7CXAstwmudE9DJIGfE/Waom8U/3EIodQ5HlhQPLrE3CLtw0Jbj
esIbAdZAbtaPpRBreFXaHr8krOT7RnXMa8PX0ZuDQc9RIibXmi3F57WLMg2zbe4X
FstVADvaAP8G6qm+TLvFKdAp6JlFEMUmrWpcP2vXdnByLvbEijWc/7tnVNW+S19n
tTCRapW+m8GVLgR9Us4nYVfibtFumvzuLSt5427VPxCc8zvxvOuigYV544RNFX6t
rElPVXDNgIoJ6lgRHtgmu0epq8NtXg7RDszPM5A9X7vbJfJI67ZxpAoSel4JaoC4
OgtYnajtRFHOu180qM5yB9oZ+zrf28bHFHoDg2L9Xol8YXgbUvrAOzf5SpsdtPBK
/rFsOgktG/olZM8HZ5lwIQUY0iecK/Ey4CFv03fe99AzUtlfklZbq3H+XavVgraV
JgbvRfQBzmrJc2yzOOJ3sLNZewB0e23L13h5jVT9Sl0Cvr2CNdnVEvn7cNtYzKrd
C0zIP3lz/Xh+CwTf+/bmD/UZSZ3ivq+nLUVhtfceLjAkbLfKqoq6993gt3xymgWX
7hlPs9kl0nqWQmhDD3LmB1ghUlDrQLLR5Xe6xi9iCS0aa3aeRFwBQJlbjeC/ezf1
JrWU6/1f2p+HeA267rUHLFgn0OMt9V9Jct61TEsEjwHzb0LyBxRLJBO6KHEDPRgY
Wu9xaQXtOFCcvobhGSxUidoLmNZty1jPZCrQTMrhVVmx/6ZsQFufuLZcQTBgkFI+
z+fZq3Y/W648a73r36U4cF8nD2q19Dq6I8vjmH4KHDKVbP1q0UJyubnVAMEYs6sv
4EnyrC5HnRjSxVPQEfE+JTSKZ92nbx8T81ukknj24Dev7ttlTGTVB2615WgFNjNg
AWXaeq8Jb29IKdd7DKpNNnod8CBwX92/bS5eUncjmkswjIg5Op4KNwwD+wvSe3sU
pOhDAEZnjBkkH6PDBzA2+EU0Fd0+gmHvacKSToQApXElBeA8V+DFAiREQg4Lr62C
A0wLiwr+E8cnnNiPPhgSoEqrOlX2IdDc9g03sCXFymEfMZ0cbEmihB9seOcioW6T
ZWPUx/CqfdfSp+doddxcuaQ0o3XQ2kU+rxZ0PYejU90XZGyYFHQObW9J9/4naV7D
flCYnXvW06jkGou6yfEz2bEjeUpWnJjmVgtLV+2chFbdlu034UdeyoLma8Kn2VyZ
2HGB2jfveZvqnuCqSGz0jjtRX4/Cc8BAzuKLOg6FEDzIIpbJBedc2A/IyRP4hvk0
OGM+JkmlZcgwNO0lhldeojjEHvedNuxLJbCrn9wYu3ii576SaNEsEN7oZuLxaXt2
scxPfqjkRvOcRRRO4Q9l7hdxhTZK2k+rX7fdjBm6cLAMoIh9r/+1mDExoWgFol+d
rlRoHhgfroRkqezq2MSDJFNO1605Fe3Jg8/65Pc20SaP9BD8hFfJuZ5p/QGQidjw
V7b99PT9sfq7w2Q4XHXIS6zzbNgpjWK24RVczYZ5dgUzXFAgOYvQyYMRAUXiXhSX
iqMqo0FKqDqHUGWo93fE0QL/bgjmiQ07IXzlnjN12e9A25csJpMlFP2dXcMIfC3D
4biu2YLQEbihan9xQW9xSDlDrHHgYi7b2DZrnVyG9t7uOGtJC+djDbtCUOXyW+pk
cxUi9LPP9TL/26OGwGWVWNFWBir372qTUr1byzZtivhI9f6+mQcmO9MgckgQSSQH
YAkSE8eAqDUthWNqDsSfNoKMgt230zmg0SIJDQq+IobCm9fu2nvi3X2noaRpvk8l
Yuo1k4WpInIXdJV251Uw8CYMJNKhMptyDRe16Q04zHnRBg/4Rcdj+aJFK07DpGq6
WRO99pIBD90t3Qv0qVwIRbtZLTA4cHHIrTL7UYCMozliwgSw9E42QIu8egfEgWYx
3qqpYeYMlBNcw2WZ9ZTDJ9oD0M4vSJeUovREfyHWCECbyMXlOQwnqcZtAYf06CR/
oSRGEHYgX+nVJPPbjkVUceltvAztEOT+xL8QpHN/Ytct/xqCnHp5a8AirnJaSzqd
hpDZkJ5+aHbkJT1CEO158Q0OVgxSvywF/5SRNEnPWpQtv3qAQxd1FhQ33XavcAl/
CMzqz14cJRnvLF7tQnbWn51ImsAkcvypkpJxDybT9D1BuYqNVCmGYO2MJS6glAeI
vWgKGvVB/Ku/Yzyso/J1cr/2BC6c7Ktlf7NfN99NZqRXq4Xzt5aGcfSHNaDoqLo6
3WCo+g3JFYbPG2KRcZT0MNRFCXI7eiB2CiumHkhNxJLqjhL8IpsN55XDL2XJ3okT
L32xqwhnsb3Z94UFwHA4Cz3kVZ6R6Z/lOtEhiLwRCZCewUaYjWyJW8McA+Ub0vme
IFS206gRu5VaaFmk0ykutXaDuFf3hkQqGQEIEYtlq7FFIahS2YmSeXTFVE4ktXpb
tqhTz4f//OCG3E2yiFLdr6lp3GHAQ2BkOqg9StktiTZNh1JmWAwoghjCAdDOqgLD
Goi85tK6lj6asHCwQdks+rZPAimOFxdbG+jgQaPVtJAQg6trJJELZLR+oPPAcVgj
fwAofBJvadhssPWdjqDulexB19PNB4D8kaP5bZc0PG4v8qGVaQS5teaZ4uzqDT8B
SW7ubtW5yP/Yn55qwoZDJs4OCAnFv4vJK6KBk0mosIZcFlAoIriSg8oHEM2wtCeC
wnVz4h/TrXC7AEnusbuMFQNaWeZ0n9Ulyrl6/75WlerTNPdl68z59UZ5j2cRNhHp
UUzMk8XoX0i1GCQuM837YuFv7TyUluJFnvC4qmXXw68ztliAmUkzt8cug2imkow/
4I3uo28O8CUejqQ8qkumtRimZYmbwiGSJ5JoolUTh9HlG/X51NO+0x1zgGshwz3q
tB/O2h2NmStLnJfH88XhngNlhTAlVzViQdgF23sUiQN+BIFLgDMFlQHuRUv6S39u
YjmhlTNUDpma9N3fTtq/VU1gDqNUKeKi8AkIcyutPa7gLlo7W4RWUENDD71aXvcm
QrjxdM+drWWmqcuV2RWLB9FiKr0CQX6dSt8bnxqFhSkPYGbFOqMOqWbRP23R3HkR
q+deI8fglHR8Eb02nHs9khCUWUr0DHWGRrGirNROlx+FVx0K9e6THpvViv6A6Ckf
ghtDoiy13US1tQM2xVXZXmj3pkwu1frNpP2QEfcyC/cnrkcqnevm+dDYdNS3xtfG
CeZQErcQsNQfGfvpcDEWDAC7R4CoYeUx2AsYDs7nHoSL9aNTw1SZzRwExyEo/udP
67URFLnaVa8GsMUgKUNl6e4Zg1ea+VhWw8CdACoFi3p7cnOeQ33APFW5arFFYKhB
tnTBKLc/GSA+xYxwbkGEqVmqzorFKrHkGwW7ELNT/HxlS9Q6szA58eEyig9INIuW
Ny84WE1kFSvSMXnwSUdO4c1h9EVxiLuxzJIo/zxitJ1lt6Tg7x49YbNrf0KfiduQ
xSL8gQYDEH8K+NLNTXe9EUHiT8NF+EF2JebBHdavWVup1S+6OfztBCvesDS9s6l7
wBtAYsNPBx4k/HTbBzeRH9r8oARp3zQaK2f3T7WvmJUPZ0MN7VSPxEnhF+VLUHYD
uy0W6P/5BncSDX2xGMHctFc5oEcqOgSsG9lbpZN0kCME5qJbeesluZ4clY/RrC64
XIkVuX1PcI1M5WDDdfNplRLysjcHgXLgKQxp64ZCnKme4X1Vff18Z6cRub6IgwB8
QDEz5zDQQvRZMwf7e2xZUZI8N8sXErGq1OGxRX1WB+aK8c1Ra+xu9kS7+Fxhk23k
mtS+32SfeeO3Dytd3mX+EO4mr2Yv3i4QZhfLWaQId7voD+ZaOoIrmrIzjeRBnv7O
6dNrMB1N/D/dQt1aT6oS1hl4e3sP63VfStfNSPU1xv3qcHOg6+npp7IDg8rL/ZJi
uoUiTUx/NXbmyL6hYXK3NTnN/HpFwwaSK0hNm30eMVisg5lmviP61cnr6bEV4jlT
sUkGHb9i28N/0vNgNbrvsoHNapQO2kQg1QH8OGRUD1llaNCwX+76p6oAWHBdNmWa
9k+PxiQNmvrjL59kfMiBYMAEasHBXvyxg7z6njY83GXxsAq+kYnzv77NtE+YmcC2
m/UyAXDZ3MwgJtb/u/63wCzze0U/w3BJuFyDWRquDB/1TgkgKZFPAycUH3vQnCAd
tIXoKmZkFZFVc2bBGvbKbZyHMCCltSpxb+r3VclSUFjrriEcw21wW6QT1G6n2W46
7hzNUHgnXqUD5dfnKo31CRoPsYz+K7m5EhqbMX6WFU7l48YOLUdjL83AX87kf36S
jYRYjSs77wbi5GPaX4Qt5F+uWuZ45vRWejYhU0oEubRruBl8HeCZ1syhMkjtQsW6
Z8mFNRGVllUhFfs5EifE5bKFfmKFyMQRCr+CT3/D5WPzDH79gaVSmMcZsEbDfmWH
RNxPLfBNM7TComgdaU+WcsjicFo6L9eoh1C7lzQLjrfXjAYPYVmC7hLUw1LHG41H
yQ0WAbVyKKu1THCaQuCY95LXSVF9eElfK6dQQvba4PsQvDbObekhsOrF96+XBEDM
kM6AsLHc8mvPTgc32/FtjQTDT6Kjsr6l6X03HjElpINiqMrlJCCRmfhebTBj6oGf
eUsaz2UvDgjZ9Bq+7weTRJGrPCpygTu0cPH7cLrGlfapaBiZ//yQdnzfKU8Nlbgk
ZBQ3m0qSoY0ODdtS6/cVs55F8v1JDgFYUFeUTa2TfUCyKzBsniUM2pbZXIufCzMJ
jMWeIs3e7I2GV2ELxjeDIzGDeho39C4PlAq2lNwWpnIoOHFC8nBKs1mMIcnpx5Sp
Yjqb7lZZa9wAx/IxqwJX7XKkPva7JM0XOj8Qwehkfl14Upv08opv3y3Ixwrx7/iv
1V8hBOJB4km1cgfQFNTg/VISCc7L2ubcMUdj2p8XyRKHWwmHGSj7obpTS9PGOj8F
gVsdnDXpMXteD2AFj6YsmOoiAYKD/gCI2vZitxR38EutX8uJo4vy8vad1hnZ14yS
Kui7NS/TQunFUK4E5pDElcthytqqWAR5JInXYAusESf+Lh9NZ2OCFUmnCeonkkLC
x+d1SHtqM0zMgQiwgxA2UpdAsDHYXdonmS71RlRRRpqDdAk8lDza47mzTbHdKv+Y
4XcZdmEbztq1MLgVThxV81aEJR65A9q8LWNKjICE/geHgkF3p2Pw8JQxpc3NmWis
P7M79y/58f2IYESp/g1f1isX/GJbb+EFbLGN6TxWutbvjOs2Iv+pztBtY7zjQm9y
qgYbZsA1v8hgqXc8ZMkbn5nKHWQuBas6nMuSAxE8HoT4Pnz+zO27bzNOqWY//TGO
t6YPmpIqKSrttsCavUSEtlppO7SsdJE1poQD0tYwKNz/X1rXMeqgWV5BpMUpaWjN
a4SzyTKpU+/V2RvOAhS23JSiu/I7gzKh1yi8Vd7Zg/P4cB6MWnyH4b6skf+0p62D
i59CK1Egz9oQBzWw0+d6GPnFizZ60iBrQwu6Dzj7Svdi+efNvCDrrMh6XzhpFfab
xDBrjukCtrbjOrElsyqqxJol2W+inYS3/6/tzIRsxvZzxqdVcGiRAFB5p5Bv19eJ
2ltiz7uncInSxujoNjJcu/oreE1pVbSuC7gtTufWOYnikzjboFvrKe3ZEPOI9WZa
3NfL7Pdr8l4zLvFhnQsr5PtA9r3kvm3nmM+W7P9XKo2Si3gKF+Oosz2/rIagSJkf
WjRbKfu90d8+GnJ2hzTTWUEK0McNBPoDz2Qr8Ynw/99yKViGT/pp8pVnZBaT/jcn
7lXLCHW8e1b48wYeU5HDzQYnzafaLFcDrExC1i0q1iH9gvtqjOMMVbpxSO2GrU2H
0DNMBG6bR1ai3Ckgw2yf3IQ0p6gHE9FaswmJBTApk8mQUeOM0m5uM/513YLup8Fr
mhxF1Ivjc8cKpNBsuuJIFzicabC+gUovD51U1gO8HAPGSssU3lL2oH1lnrnuHPw5
wnFL+mwrl13Cz57YGI8xFbGRmOGA7/Ezs7gCBKdBBY8fQUHKgJdZQ8aNXxW5NaZN
rIsN0+yu32Nzo/0Pu+YFtxMIRUimwApqSU8Le3ocXiGM09aYgevwNyM8L9LpcMbA
uMEWL4vo2HcKCYBRVsvpyZQggTV9p4UbFp0eNJ5BfT3oaxlNIr7zTbbISMK4JL6K
1qXXRxv2GkJ3bn3KM5sDfxMdSOvgndyPDCEcKrMCLfNNyJwMcGJ5Enw+tq7A/Lch
wvxzfT8BHOaomCgzZP/WjwfoyT8gPVDjg2n/q66pf+d6RaHleacXa3DyY7e/GwY3
xqRz77OS1epQ0dqxxAzAggMwG5cPUVEr6HuTVL06kEoJt0lu+lSNikhOB+DQmROS
Qh/9JB+wKOmwYd+dK+2hVUd3gEuInqbNU5aUt6LHkBhNW9g3RlJg3soVTnZ7m5l0
OOOHcFVwl5s2oVUATldFZ2YB0XEgJCKdTroTPe+brVMvGjo8Bq1LLYS3VSl3Q/v4
sg47DeIBTlUm+l/36wccAAMxcULkvZSgneQve+p4A+YJaRW9lyc8TJFZo6mVZF32
BCyKsnMKXj7H7kyQ0dSRFOfmlDAWubxZcSCXPXwNZiQSm5/2yKsP2r0J/CkYVk2B
7YOtmWq8VGxjTKXnO38iYHQTy+I1FtGku+6yKq+ulRd00dxs//DYA/NZL3+w4ST7
TEvzceD+Obu3hTJmfUs6GUEX7a8dJK7qQjfibC5IISqKCUv4gMS04AWFHPUUSahh
ukQtT2VGn2122SLVYcpIRO8N6w9z9Yc15A1zPDqky/NxPyvFGhWDyv2HaqjkPaHv
YEzqwfbrN+ZsVQPNsVxcwEy/KcsE/+/ZMgHmououb1pbWjaifNGABlNsTBKLJNIR
/4Lv6mlBtyYYq4SZ1eQbCAS4azXPVrhnRT53HThscVOHu9A78PJWsRA+ubtXdE1c
6qc959VAG9Z+DqyoiD2tD75tyvm7YQk33yd52t5uXw+/J1rT7s4ZbFkWfuoFDvK9
GFR3MlP+vO+QK7jwzSDPPXZA2N/xbYA2gLChNj/vlaFrMHbQq+iCK3mnxcT3lCsG
JnhmTUC4cVvVIBRXOe0uMl3fE4oVUw+P8dpl1QE36EpmIJ/HTpY9tZmXHjbxILm0
D5d6Qc5NE1T43hvcswgxBvKlW/Q8PFBgXuUoPm8dp9YPUFaUNMlpE8XXSuk0g9To
PeZF6Mwnjinel1cUQZc7MU3/Mrn6XRt43VOvS1w/WBjreWhBpQ4Zu8mYxmRqoBjh
0x/03+Ch/LoEHXbvcPPTkFpCgH1iw3zzOP20fd0tsoV3B90wgPDhb4HoI0VVDy4m
Q1+0hmCsrsi0TYzrwGB9rHoyhetVsYfVHVCAMv7TZ8hQ5GMGkUeCX8jd7BCG2Y9R
gaXTf84JuXg5Z7TPJBzeQ6ApGCUeNLAaUAUtJ12jj4yP2oRvdrsQgU74MeYL52HJ
5NZSbH/M3JrCanBAKGS20ok16WLHpaebhHFbMlH5haWC0fe7AVETF3ut8tXGGSdj
5EN4eWd2Swhywyz+3UXNJnKYm/zqV8Llp4XRtrt3jeyRe+hsKOwl7gTSPg4342TR
vv4k/qhSBQQlDTUnmDkE/5ba5WBhFSIR75AXeA/BZnTaFKQJPfD8jEcM//VHpxf4
tTxsLoQ6wwzJkD0TiL8P8iLih77OvuEPyT01PHS4XRW0lSHbrx2lPdtZOBNvNKM0
lFnQS2pSJWW69Ci3nwa+xSB7yu2gEJtURwmgEf7NmF3abqXEPyd9JbRnFEkRolgG
SSVLrHe2ttfLHJM55SijXAwNn82bY0bAsuMy+AENspkWgZ1J7/uqZBe16rmAAyRp
wqL6AE2TSnwLnylfVFTXGDqkFZp/zbO65ium4C2M4gPIZzCPE4vLYpRDCByU2CcW
IWWwr8Gk4KT5Ms5pzxL967Q6VbbngIgcjgD0NyvL7zYSep+X0G0CPNmayGyesEhN
Z/uUYyB7Kg9tM1uDlryRc1pSI24pPKZenCYeBuRnA3VgWVgYfKAMgEaLVt1z4F6v
uHhYIpMi5V3PbnpWKh3YidTZdrkjDHGFjOYaAHTLF/yIudB4INxa4R4xp/RWXEIq
a2WxtczbKTwiQfmDO1w/DztpUiUVYVBcZGZVMevVi8nbHb6Xv6nNbscrw0GMdazb
tMIEwZ1oGWGuzZN1i4EXiIQZEefPwqoJjxSYjFNJKc9XGHjRciLUxJO3cDC9YzZk
6H/xevt48kou+Wmo3+jPU24AQVaX71r9T7p2mJT65R1VLqnTheOsfDphIMWNNZjX
gP+stgnTP9CRdzDOxe111J5iFmUTvSNbJJjJY/TjDi2LU4/koc3QQvlH1vrhFGmB
3S/q+dSch8VJLnBtGV+yUD2Vqvqk975voQYvlbxiBfXZXjpi74tz8dYGfIZowO8r
AHpqRpO5oFEYiFUK1I9KuA+So7CsC+xPF06ewU5ovziyflTnde1kjHzQvlb3MM5s
q02nJQTchSPliDzMZe1ia4CPAcYCKnGAD1EwEGVE3v9S96m3pnnLG+BcTWQK6+HV
sbhnjFZcXvu8kco9X1OiKMgNGNuCHaWliwZLK618MWDW9N2QCvEnziLia26FwLKd
gGuZGOrmsEQ3rZbudW3JS9Jkajvx0d/pzTX4j9A16xe7HwdWWUMCen3rRVZzTMA8
UL/6S++3dvIV17Unfke2tES7nFH5TKB0+3QPzB6Ho4qPhww2a05wSwMEYLzTL3gz
3DTz16aeU66U5fX4pzxwRBBvOdmUcvj9IBFxp1wkMcsNkY915H6GTNCGg8X3k26p
63g4UbY1CKaBjKVikaPN273zXSxcKIv7ZwJlWOB53qMV0VlNBa7SZOoKmrsPYuth
OzbQdmKVq/6HsCZwxwvN2zNYdkfOIBnuio2+2qtX05ytg519O31OTTjSo8ZChWTm
D4iWmXT6MTQwHT7Zhr1G2KNLfo5in3Tc7dz+T7YQ7BNDMtkCAakJEHIUQYRg9/rd
RNSYlv4wA43Jd6WXux/C0E42u9L7tUoLhg4kw5WDOq0MjhWWwtiNPh2eP//c6IMR
UD1wWZTSUjP0TsoD5G+ObFQo/qKJRmlV2MKIK0UiVx/5qHzD45BBdDJQSp1NYw1E
LBKl2sq3rPa9cqdleSvurd4v7IFOOJdIPP1dmlabzF1WI2JwQbWKPS0a/6vpyXtZ
HpRptbyrY1UHG9oFTuK/3H8e4jAF1VCnKLYJniryrhmcMjbY9HEG8gnq8qyGmnAY
4jyzp1doqS0U7+C/e9dGc3NhWQrRzHNspG7i24x5m9i4pvbxCM6Ru1f5CjJwQHTA
ktyLcHwu6LAic4mrUgNmfnyRpCJ26xufi6v/vB9L7i0MmJ25wRpTKq8+fKoU9MMq
hGIYQ/VTQ3nNbyJTpbG6ZbxQ+24fXDiX39sB77JDypm+d8VO6st4QJ9Y7nv+BY75
pneOd7h6zD/vm0Y2ificW5Ve5UIB0WenFOqO1bLZc+1f7dfCwKf3Gr0uZPq/pZGT
3R27afn36Gjy1BhFj7VUWnGrrE2/HoXYVJqRClKn8gOifWWVyuiuhhlwReeOQ11A
Taci5LyGuHzwNynFvlbeGgtPnlhxSqcbBGGUg01Hh8Kl3K9bzQT32LCmbmeb3O9B
uNGq5MTNLAmqAwn2tId70aJPLKn+QAsQ4kDMcaguZezsgDAEWEqnPAkfBbDucuqr
/u8iNYBe8c26GN0P+jfQxI1cO+iAledRtTsemjBP2F5Ls025JEyO+vAUN9niT8fo
/QPJ8877Rl2i4oFrnKqw5GOBACx/CfqcuiyIsRmp3q6pMq54jLoFcILoUJQCCIsT
HayETM2bXGkz6o2Pm4rjyxc2IeJYByKWlww4503H5Hz7Ro4HhEANtKwH4K76Z1ks
1KztVske4RdMku3WPA/3EskfG6Ik3PTwFlLQMc4pTOofGqo/fKQCGvZEGtfMV+/S
GkiErvb4fFl5IYsgLZ+/VZdFUoHTnw/nnXQjVv1BBAf3MWk9XxwQi0aYDaizXzKp
zbp5pxwEB0PEGYZnZBzmayKrB4eSsoyLqd0tbzE03a7DeXmHqE8p9cmiCKQqxXrn
kW0TBqo1yGWG7+0aWIIEF4jExv6wCXVjNdUEqR+RLFzwf4i286y/HJTR3WuZZKZ+
kvfwpPk9PZsb9x+eFfCJ9zF4lVy1V8PN+e5GeV4boD9SGkKuVntaF10CZEh0V4M8
ESqyFsZdlHkPuAusTijrI1MhPrQ1xhDZvqI2+fUf/lkKeQBdsOQ0+78JTMIQfzJl
npa9ka3RJ/oQJ6CXFJmAw7x4V6VjrDQAMTokFD8cNqJr/jDlU0WYfl5TNWZJxEXU
1gYRXPcf6Sz07PqwGcWrZiX6schi5JaxlLQRVkuYzksNC0gCbvGoioAdutgczXi/
EfPEN1VzzRhbNmHStvQABw+4OALJYccCzjbBiOI7HYxN2CGzi/lmc7ms5Kdwb0hl
YNYyoukhgRpHRmF+QpAgVE3ABZ1gG/M+D6uYS2xTQ2kKn998rRm+t/Q/1khKVSkb
FarZFjNCUhj4Oiszamzl7RxlQAyqKSABCuFuz1Vv3qS5Fp+4drftdvBkv5P9FQ70
dFfSpMwiEwvSXOORs0jY7Q+quG8tZK5BTXw0foSiOQgHDrDHAZ3WwcI4B3KaGACz
y6yMyW4QdbzMolXfFwBnsPCEXMIKv0LT9VzBQyA6jz03rPVPqlHa0CCwLl6vZIPf
S7K3Vn8i0JOnWW8LrSo/4Q3yZeQ8Lw7M0z4r62ako5MLYQvfYcGrkkkS6fAxGY41
zaMjQNUJYeyi0sfOXfLQJZ/37eARge+zxhYFNE1LK/WyMy6l38ZeskIRsDPwsPcx
1QOv8UE6dhodyEOp1HH0/roPzld0Ix/JkrvGAqM0wyf/ip9zExS2E3p9X0jalv4g
m3cn6AKyyrYQbLuwGzpc5zepaP4rbIw/F70ZzIk3IfBNpaSaQYmWd65J+hACEjBg
gTQ+mF64wAnDySQWCHbMyy+E8QJwgOJL1brTPmjhlir4PXafTKaWezfo8dJ5MkL6
6AA8J6UZ/aKXGnlIAfNJ0akXd48f6wFCk7cnfXWQTP/VKF2crOccsWE4vYlrlYG9
HW+YJp05fV6sCBP5GDYBw6vwoEUShT44RsXclHR0HnXVtPCuOr7l+fX2otpa+gaa
QVUrYzrndUIOfDQmxGW8Z5KPNSvWUptaTsoZc0u94oZDOQOFVlconY0JKR6xt6ni
VDsCv8OdgJC6N+ZMvGIJIizYvxpWp4AYsIyst23Yj9/u0Oqp3y29UTxvCm6vvxse
Liv8dfQxzSaNBCCVEseabHsFxoy5/esJohjJBlDvi6Cyu6De1VdeBXu87Vfwa0Co
tvLeIt4a5iXGUxzzStaQn1i+I6f7GBAkeP5lTK+zNYKO3MuUDutYm1ulxUoxc60v
z6oAxGWzLYVMhlsubMcDnrMe1qLWb5nHWpgaUAzBbh/iVs0qyF0Q6IVW5klurdNj
mSiOWGSTdL8razTbopOkGXTVowrzL26XDuYlhsMJ4yjw57tvah/FhV1I05vs+8Xu
Qh9XkZzFccXOceedH5dnEn61Od3tqN/lgZClP2ex76XqCL7moVBfIe2AGS4KaOxv
sRPYRQ3Q/tB42cwR+PLpnKY9k+EzuYtUutQI92GFhZEC1DhWAQKCTbVUrrfIxci8
X62TR8T5uaYs2P05a+I4ayiYqaAavfS3DH/+jMhRs6la03HFENyoZQUFuLZr+MRE
EQbIkogZhtQvRwAkR9lH7KxAFTtDc/UXtF3Ie+7AkFAo2uaQKh/rrfAdOjHzNgQt
hnXdCge0vjXPhfLlgQOL64Bm5o9QcOAOddy6TFFdf+kW3hsDszxD64mfYU4Anf/v
NOB3S9eUOFeTt3Ftbe6qEUw/G1pjH/3DR3W4T/chjnWrsNT8l0qH2+T4VnzcPzkN
6/fXk8rODfnuuK/dRsZtyTJ4X7eaTi/GEhb89M2xHnT+5Ym+oTfyKHMdaTyPh/m3
I52qg1Us213FWEJIgfpKA5/TSZcOX/oimKdqSbExyeMZayyVjd5gf4j1WZoSgOr/
HknBv8kGlfAmRRB15whDDCPxEnh/WbVPWqncDAd+XxSgvI5+2l+OymLQ/0YFSbzL
KlT6M9jMmIF7XYse4+yn5rltuFnaaSeS4wCxnTR4flEZ4EY6fa/vZforCoNcYYJQ
2hr+btzq3du2nj+4j9hGGoXgOqcsrP1WKTp6dv03ej6cmt0Omyk9Xnxym6slc2So
Cszt0rZdx6S8JvdkY5E8X1OEqd2FHUbxtvUXNYeS87cn79JkB2nLJkeghtYwYZ26
GtSgSZsJGjAo8dzBZJPyBW0ijg0niRe7LUjsfpAg4vnrqyVN3ApRKcDxxGVNV1Rm
kczAv6y4FNDaUxWl6c1aA+9wSt3Vtc4WRTT8Ob8jpL9azH1lCj0neOsEPX4gF4cy
Ij5xKuziSHlS9q5MYb9F2HnVDvvhxKuuWiikVUQUvBVh0mBBuIGyaoY2BdTUDzB+
Vy2m0/634QTM2+ZTALFvxETdTqGjuPwxMrMH3ua8mg2EbliparDXPxBnMtVVs4/P
caZW6UkaUEpWbHW7UTGpXz3xfKmAoHsWg1gmbDHM7gqgJ9wJbvzg810WpNbxK8dz
pd57xOSvP0FkQlYojddWVIy5zuGoI5DV1iq3DXkK17+bm0qEaZCVHFX2I8nHI0rf
B938Ny9UURIvtG74sESvKxZ80vv8qCcuJRQoEXyOykg/UQQC1/A23Dlrvyy44O4k
46huq3PjsUO04/z7Ie+b+jFQxJjFohsRxmMecCW2nsjiJ2ke7qZsRPI5/Ew6ZYAF
g/eq8sQIBQsJpdynJXK5zYsHeGuOKqt8lUSupz4wTKON/V4YVjD/2EvlKfMQmTEo
cBcqMXFAdXPlpHyn2Q109mIabRoluvuKEcgyZK6BpdwXh66BmnYZjKrepMC8BYn4
5L4LJYVY+4++7VWG8+Ig5jnt2c3Vmvjn4cfUWpbTorZF+/E0jZ1P9h6/cdD2kWPU
wQsrXoSAN5vJYgLY5xrwZY5PEkOVvyrVHNTM2Kwo1XHPEiqqACQa3DOAcrFEO82f
Rqr62SaSiApaDgySFy3fYBsr5Cq/ZyQH2WbIRLD3hfiAcz+V2AkUKFgL96bv1poB
soNGNTkbNaHHrNzeg8tG1Co5yAF8zE0eglqQgg/mBVhz48ccJ6nCxuA4Pe8W8/jU
sMPcsbk1jJlEVrAh9r9bZ6PCP2LWf6Xpg1wyTXeFth4t3j/51SwtU5HSG6/N7zhV
0jQtE3y/rTgEShLgcwVs9apVItChJWYQFphZcjlyyJBkfD2NG2BFi+MWPjHwhU0Y
Q0p6Lv/jgxAT6/d9Lw6rD8dHkJM/UQ6GLP8s/lyVOuH08MuEw4u60EShO/lmI/YH
59zGN9XuYeOyLjwP/sJF8fPKA7mc/Qg6UbImUagDgx6NgdvwBvGt9ydQ7Im2r4QR
OzdERvvqdEDjbT3S59g3KH7BpEi9O5ITrvx2DU7kZfXK8Yq1Mmgdis3l4Jho2pGV
qgKTCaS3pwyXZk49GgiJBz5ek77biDJUrvXp52Ziw2LklKyNh7L/FbeiB9+xoM0r
1Pp5+5nOp9zYBCwhuoaAclS30Wsvsc90WxCThIvlpi7kmKeOLwOKZ3/dcxaIKlCO
DPNEXuo7MQkWRDl/0YpNBZ2P5HS5uxwYMzV78lHJDTw9sX/He2tptwXCoQIJr3+Q
vDNFXklLQfPAb3/HplKxF6CpPTEIdcgjfdHEgLkwoesOvMcei9NsVD5rUj6QUYN/
JoIHhQT6cArA+PQQoBjex13rtcxXPBOtUakjwjCuW22E/2P2t5TsAecj7jyH7FcY
MlQhnRIEYG0oW2hHBLCsFRclf6+Dcqd4zSweupN99hqzUidSRat1huH60wo4eWZk
uP8iecOSRPAoNlwoRfIp3QBJbh+5mAyVPCs8zuvr1DPTu4iECRfsO7K69ExKRQKD
YXqzTsJ4+Fl5bSMGOuEHy/K6Ck8US7RD19ho2TocEKNleA+M2mjuy1Z2C5eRuC8g
NbJy1Pf2JKTRHnwntTJdLM/lsisJqa9uRdfk92YpsjQE+SoV+OhoZGt32YydCJ7+
YhS/QIy8wfHGzGjs0Zs9O7Hd7VTrc3yTE7xhQUw/o+l1tXjAIuVpku+y8AoiTN3X
wKeVOwnWaQcSgm5A7UlP5P2QS+LWudSSxMHNsM72dE2uLipfs72juJs3XXG08AD3
0rIuI3Pm/ffHloxJrHLdcttOY0uqThDKyoldSnCHedt4/AYOzfDfw/KuPqzOLicn
NmjAXq2cvjKOXg8nJ4jafVXETVPHFSo7L6eZDoHAd/dqWkHfe3SB7ldn+7zyUZnz
ugY1LKz7sLsUWmt7eNRinkpdNY6r71ndVdDDK6VzEvknKt1H60uXvv0LbiioUKn4
J/+SqgZeF6bP0l6AYsFWQLMIQPFKS2LoldjrlJx4SfNKAyXcx6lE0o+eS0kQsoQW
J3jBZFLUYsNM/O5ZL3TvcCPLzDKvyzc/tb1xVYLeNDw9wIoT6ByiEC3ZBnGdevth
d4AM1tZPSeNjoIWidrS4xhuJKV8Yvb8DF0CHUOC1UJSzLl2DGWldCrGKr7dr84bO
HenXhAsM6FkTjZZmB1cd4ss/oRSd6KOJrRbW1iGyOe1GsLAzbUWRsULQrCd+Df4D
qzodiwDSoTqOy53gJ1AeYR3JrgTWWC+IGQE+ee41cv0nUCFHZY1QJpf5Q5KjcAHB
BtXaKtWGUHPuM5xoaP/tNQSX5Bl+B4N0qVhjgd1dTGH3oPCnwcCg5w+pl1QbGs1u
9MPI+wzcT405sRKm5Nba3ae9Tk0cKcyOwS0sdcsS6YiENfSqLvBbq2DrfEqPa2hZ
EoZdgoq3p0ivTlrWZtHfmEwengLTvAJ/Sljh50pfYyBFoflhYwyBnCIyEkpdi/TS
k1W+W+3eLBR85DD7XG3KK1qolOrv2PWNedAjlSRq7Vn5ROEgL+h2dQ8QVioZ5bk9
mE4SPfl3LmBifyTgZvlrjPIx1e2okoRKFygzgmLYydZ/8kgPHaVLAB6spSBVg9G6
45Ud0S02Fql/RZVE5Z94c5koWm3p+a9yyJNr65KpLTjxDdT8r4W5JzvHx8huAizu
BZjU7ImFvC5RlJZ2PX9YB6ZnG8pHe6JBgDBp1yL7XW09rv6kDECZ43wey3//1/rG
DJVxmKwxtVQw6of34BKb7yRb31ZPXgessnhokeBIwdm2XpOxoLKIyMnyYpkdw2/R
1A8D/zw88nQC8MJlHk/WWxQ+Mf1biHIwauc9n1vIiPQTMVkvcOu5/4a/YcBTetUH
KY+muOLowthB3GeBYtCd4JDeSxrIEeQTfbKpT/x9bwtmUvNW8T9vZU2bDw+AvNAG
Ta/H1+h/7IE36xKglngBo2+nhY73US3ebprOsCvTsVU2c+jH4lAMgdz29y2M3tkk
kLQEtLxn9Yuq4TRV8PiGD75KSGK0Gv9U7mI2bLjxzxh+3eTt17E2i9AY/wS0bv7m
1qKqENGmVthlN54B1Vbd9Q0bFs1V2LAaAFK43MvV9KBwOH2rs6B9YfbJzcp8MF3K
4Ki0pkzCRLfsJr9vZARPzykZOPH2gKXYxiSduleOxkE418pVqoSGK+y0lVdlGfWl
X1EwkyrzLv0SDROn3IImCu3yVWSPKZ9+GxE5mwz3CtHsLXkHsfVCni3fysH41Ka+
YMG+Y9UdF7vqDK59bF1rOfC+e0IwDXH8+pS4tbE1uMM8XAyFU/Vt7J8fM791SrrY
K0js+Bn+4bGhGT99SiMMHrlDsjE4pDJK4YTSsNy+aL5sn4P7HJ5MTfJsDS8f3ds2
3nV+1a8YXiS1y9OsbUNPwrdOLCm6Z9M6fUFZJsnHww7AfCyFKy9QxGyn1R7jpJsj
pTr6i4W+mJSQtWPaAC/LIBZ4iwpj6OooVeQH4aFNB6g3w8/CAaiOs1zFcaJmcRul
QspTdbPCil/cWlxspIzUbt2KYAwjh6Zz8vrfSsLVPQUjax2zwlbvC4HWKBXv9Add
N7OAp2MdwiyD9kT1lhu8wdI9Q8/fQC533rkcRSJHS00JiKqjS6uxmGOstHNWglqZ
3uYG2uq2Ibrsdb3eQXH3Mu/Np4kl0qWtgm2X7dy2uXqV555UJDQIvsNdBX19S+JN
MgB9HMfdtg7nH3txHPbScjgymBSpjQMPM3vvgKIWw/dfbDNJs7UKreJ0wxZstGvr
czsKLTgPSzvOQ7PTFhG9FlU8p0iHlr8BNGeaffHQrxuYT0Sq20Jb9nOauszl56tH
NTx7vauhwmQmuptDiJGpbQ8VlJjn3+Y1ViK9ittHvNLYiIOZtSdrNoKZLODDz324
OFzTo+ENmmU1eNlQagdWe5CtQzJEpVkOZzXVCBqzRGGeheZKAUG4eiqEcanBo0Xg
6c/sAAaEkMgQcCo0Em/LuEHuQ7uXKycW7AwuSyaDz6FIaSgMDSutLdNpLJHatzCl
Zm4UlsRMWA3QmatT7vGyFBu5/jnWjYpJ8gpa4oHEu6aJuPMz/2tTZtNYBaHjdr3N
RCq7fCZfD1N4TBeqD/OkfyOBxpcam7Zd+wJ66eXIcc89EzOhowN/gPlT3unBbqN/
cm1A9YrGQj4zBPsIZVYNAJY22LV1jjOzOehBmK5ArRep8aiiOlI5NVsdu7sE1z1h
4oz7UKDdSK7Qufk0ef0jFsgvwzoe2EB55Vh9brwVii6cZCmZYij5WF+VE5iSAKWl
pke/mcL3SLZE0njUMWXQDApfWRCArVzK4N2wXBSaSC0kiiAE1/AxVz7LQtdViD8A
lJhho5LMYjo04L6zLGEv+KznryHcUkzHcDIyhzHKQl6OzuZCF1utw0mI74aJnSZn
2e6j95cupDKap/dHxi+6XxTbZfsOyIEoVBfJNtZfA6XGBH9bUnSeKhgndAT/o3nm
h0snFyTY7QS1ymeHIolS8uy2SPDZphu6t0OPNK3GzOIwF+8hXwrZFoFTrgElBU1M
lkM+OogMgrv4M1f6s86Gt+IC/TgQ5vFJu/5Y1kCDx7PTg7AuP2yldQUBFSzDkmcb
4+swErF2mfXxaaesg95qeQMB40cN0JVg6YUnQtp5PpelqHhju5DUujpaVW5hzmfW
r+tTgwqLUz104fzvtU2eHZPSRY/RkGQNevE9m0CZzTIUMpS91CK3TfhhYlgWAaQ7
1eHEApyUICHE4/DjzWC50bJ1iVs0gZ+Hh/x1tGiL9QpphWo8QBEGt8r3F+9zYHsF
MB1oy6RaqfRrgl7QK0hlmm+EVviepD4pgnxhVmseNHBHjHLaz/oeGjGWrDTUkR/a
9kzeGE8TTAQh2aNAjGXKohWQ+NYYJYqR31AoH8Bc7ZmQ7eN4vecQrnlbOY4LDZP3
bbVejM/kiu90JqGQcZx6IKly5OQZVUkg91AJjcbzyw63izBLxazyzYnJTv/IReBm
/DurINZb89SdYbPsPgvg3liYOLc+daBp9VtxTJjE1zKtr9ZBuJohqy7gLJDaDpGg
p4G0nKfYfoWIZMBOipvSAEp0pldlXxCeGu3QV6t1zcqb4zmkM9pb+l8oW13+NKhN
L7bnGdxsf7J4a16DTM/mjYO85F6YhxeyN8HuQit6twfDog5olOjxJorgHXtOi8uF
XYMPdgk7QFhJsNi8VWyEnCxqjls0AOZYaloeBv6WCz5o72rVKv1W4+KjKGb8qvzS
mdJdefG62ABy8MOqPwCL7U2DMWbesZ5PHbjM5Scrp/q82ytB/gATq9B7UwA1ZKRW
I7vt6P1kUJLZAwwI3uB1bLdqLtGagIwtfRee0ysAlpgzJK+sIGVW3F+1PiLQE3af
J35ykqNCt2rPRYpSPu+BVAoDsLemt3UeXwdEW+KYtGq0jdnMTiPIFFNw8K4GvK4k
n6a58wUruHj/NXuXf73fwTml5WXnl8ud/yJgPQ2AqzdghvIioz+LJowGs8LqlWfB
9OIz8jyspMq2GdU7MgT88Ewx6soqDDDWCRqHR3ApY0juWQpQwkxqlNU1w7YSvCXe
bR7M3xIA3KwiaDV/Hk2ufIkYqn2HEcAnLnT9gkh9dOr2aABd17OpzRCaYOEM4X56
GsGnLQWeOFCLCAmF2S2AWgRy3EsYF7ebtiDwTSS70jx9KaXgwmPUSFVgC6/xrI33
aJ6jan+wTQsGSl47bKZyO6HsSjfNb3WEa9P2ZUpe8yuPftO2mis8fiTW9j3FiLXR
8h3+0sVJCPjAVLLs93VzGVyAj5ErpipwotLPwSEULSiCXHTKTzY1tz9zKub9/C4S
3xC+8A+pFFA6SDi6Ip6/oj6U+tkUC04nfdfzTKfnnimnwXmRhjevBfNMikJrFchY
dycofKvAh5ARuScEiRylRkbABBGRURoLjO/LXRGHF7sEoYb6L5lW8I5SrrIpiRag
zQXIFGDpCi8a2KHnBpDvo5UtDvBt+NB2/eznHpsbcvAMCMjaVGjrpp5dUWsc/1GK
UrmSEwvBhAJnYcw4CvER0qg7nJX6uli9Bk8/zpHETgb/Vewb1aacfj0iG9qRCSbC
+EFNpywBKwD/Zo4Y7/UVqccVqt8aV9FfRTX6VsghGNkoB6HUQMKyPdm50gw0JVwu
egUfOjNcOMsRjZ6JPIlMUBeXvVAIOSofickUhUKKabQaYpLUxcXoFFL7faMkknbF
oX68kZEsDHJ3HjhrvG943rEtuSaTGlP9ykJfpABGJPzi2b+dAzjbRvimbNfgWVh0
frejYq7dTkKk5uy4Av7yaREeoNJYkzhA0ATYx36AE6O3hJ4pDOpvsryDy/9gFcmz
l87oXXYlpV+rxsZvet2W86RblRWG4LPfHbfTUWNGMsNyGjagUoiatUkH89rFAala
bYAxh60g5eD2D6NJ2kFcvI+bKDbJ+/8FeMjlo+duBddFCoWOFIYYnihNA8mxuYas
+LRDT1x0Qm1+aO/riw/ywq177lMVP2oU1GJ9exFzDdlgX4g8oWsILCzjHOr0tPLU
2/1VcJUTsZxvMsWhYtj/LtucXcpTd/e4mfw09ciXjOMdCGzGBoNANKgFuLxtzmx9
ER394oyDACxL+8Xg9JvIx1UKzH5Ttsy0ezoCu4JYLgWQtpPn1zjU1/4zRGM/QMaf
3e3SvZPV9INwt/Y6yeJ1LyPNnkVVdzPJVmaHK1TbizDr5wfLKVtD47SyGUBYuC+g
y6jrb9mPxHoFY17dhKwSQQGZfPDjfTIDImmDbqxmNX9TBodXoaYFW6AjJ7DwOncB
UlabN/jxiR4WIzFe7U9I+l6afwFo+ee/5+9HcHy3iwd//cJOwaoB4aAqaKP0JKtr
9rKTzRaDa98uDamMROl8vRURlwON38GVnkVZJjKYfc5EoWHqPsR1FjWlz/nvXE21
zb8sj2K0Fzbk/601i4xRLKY3qhBL8Dk1GeLcX+tLL2ra2sqOCqMBGDFTeKr1GW2d
SsRLndwqev0AzOqi7hgT5NMXYqCu232VpZ8Bq1/NZtFkpPd/+umuhw8T37Jk8W+D
MyHRAhKGnF5vU92Ia6/OTohkKI3FlrLybhbN5vg+ZPA9/Mr4Kb6Hn6Wh9Je4eMX9
e4OFL1nsAxUHuc2J9mPxFny/4xqnlFn62fU3EEdKjgpLJESc1E+QsUpZ8STp/DRq
+otZQNt5bdKJOOpEJO3vGxHrwQf2TB5y/Cf9ebeJtvk2z8hG9TtUnNobfDJdWKH4
uA1s/BeIhbloViOHBP31ZBI5cmvpNsEVj0vB3MFMtc8hQhsc5ze8tdKLaHY35nit
zlBlP7YXEv6A0bPMzDLEEHl+wVf9RykcjzCf5JdHLzA5GCUwqCVdKLIq8b+L5PYY
jSE+Xs9OOZAE/sfrwHeBPfYOfbUko3lQ3V1RhnJKvO9/oWFmnhu0Qm1UVxWKJH+y
aiY/pyMPRWb4HUfhcUYLMbcMvjgl4cAJMgbPF7fBXD8D7MONmOSaPCAkIz7kezRm
lc55VFR7wXtDily5d7mwqzG3hYCx8ya2i/43lSUOETGeJlntC6bPh83OJNWqVtko
9/60lDLVE0MU4xPetiGHNjh/wrAU/8sX2hFbdJskVWbvEXYOrRUACA+IhjPEcLc7
Tf8vHWnWWJaXSunI+mAKhYPbbpthe+rZA6JtZZ0sAabvPUkN6O70oXwLEUWaGMOa
dhgsBvV/BiognV/fJG/2+i589T4nZ0nsiLa8JQw6siHlm3zmBWtW53joNRGeZp8C
SFXDYiRIkkPsyV9CQ9JV8RqssqtX6uMeOv3CwgpYExAPG12JqYYJKeKw8awCSwZ5
olH1CfuoZuOdV8ZTcgwDByU/tQNY9SLU5ApbZQJqIkuVyLd0y1f7kasocjjGRSAo
VCs9YLWJPqMYOrqcVMpM2GtMLqLhnUml9SKr0OxMUWsaexDRyaBXaJ8tr9zLyIgo
u8FH4MDF8RljZalUcT3eZXcqTXPYJINZZfzCl/pD6velHq40vF71XcNDflbyK7i7
JD0s1OoLJGkUzjvwqbVks5ayHawXfPNQf80h1WZOTAkpMwD7Cv49leFvn/Eeq4K4
d55tHzWcSpLKG/CZ2fhveiZLAHBwb9DsfkUj2US5Q38b1SgS2GtbSq9PR8aKThdJ
CRFOS+syBpsSpVM2itHE4tecRl7+91lCLrXtvudEHaD8YhHGZ+htLe8tDRkqB+Xl
x1SPiyEJb4wzee3CL4JjjevNnse7/I6h7eK2iTb4zqE2edpn6SSI2DBcMNIxEOMy
yy5L5p6YqRybNZR4iu7nsSzblOkZIht7eRM6T6mcE+3zZR+4UqIOqXloz5Eq5mNa
XYjsZVICWfHT39yIHgMGBiIAfklmyFFL1nrb7hRpk1YcnvVoKevHeBo5DD3j8B6J
eqzhrKBDLb9OIyTcZbCY9xiW09Fk+ktrCJGR6MAC7XXo0qvP7yMSjyNRS87lDRb7
UbnxX5GUWDVFwvwzJOSvISQ8V3Ei3XHaqjC8djFHxJFep9/14Kil1nlzFOoQpn8J
in07+Qh1/FADIkBqKrXs5Fln5t1VR2GJjBXpWTuMwKvwp+CGtzNHbKsJtA0/1oKl
F10tDdzltIRwdyntBm0/d/Q8M6+s7AY8II6FKp5pLULO9SHsEGVi668i3v4e5e4E
UAnCzK2QuQM+x4It3U+/WkfqjKy1ivEDqRx+2k6FWhVsDW7zCzjyPGIlrwtca3DJ
qZMbWeCGrNC5hpX4zvgEVbfig0D5ThLXXfJPwFdTslsZRRMShUThRNT74J5QgCK5
D1qMMQzJ1iCF8XpUNY3BzWs/BIIzIKPf4OSF3+CIpumgjaoVRTzOz18GfN5x7HpE
JPQajXBN6qvJHVZY8yL1KVDR8fL7vxWyRx3H+oMGdVSPfn4JGQKMGjd7RwRziMCv
4MTEeuubvG1EgO/S27t0zUy6DKQdsL+gjCs948/Dd07OoqMnF8Z7l9nwngcZ0EI+
fecHS3ypKflQ4IUNbgdmjyuSSXs+LnboQ4Y4OJuO4zxmna42iEDv3OIX2d0wsr+m
Gb4nLCqv9fdTyZ5Fm7PVohKuL2mXvcXM1fIYDNV51sc068Ra1KV+aH/K0dl8A3r9
FdsSiSEjHdLTts4bbtrabDmPX/hyyuK4l4BE2TsFtMXzSF/PtVGf65+zGi8QXdHb
9y/G06tV0tmQAsv12WnJdaoNd5YHYIm+9pu868FLOMk/zrwnW1kIz887nfnPWhqq
2zMSuQ4YUmDKiY0flYvSNGaQfW4QBw1vSj8qxLhdW0ACINxTG5sPpcO5oimkqN0D
kC4yr0G1VDPCfkvQyGA5fWMmb5FwAK6Tc5BPuAow+nCOUE/xetqIuIgf9TwCf1Rt
KBPkgr+M966gS+yrkq0XlvG53LxwaRtgO7kJQBgkR8YgUXTkdBsU3WLkpZM4i60Z
IsnlC4P0fmOhANEVMa9pLfmbrjrsd9GBXoLCE9YX/N7CiXL95lHUmR1JmPQzkYFI
4TOED1snSUFzAnKg+NE9QSvdZfoXKKPCq8FAVv2sOsV6nE8dV6OfiPxH/vp22vXV
gC+9i0g5gCdW8wWMNVo/C//2m64KsszniqO2P7YNNaxBrSdbbvhbcpEW4x/xrRrj
SfNYGGsDtPX+/8jdJAF0t7J1bKdrWXEe8PSZo6eoZNNC8172EgcYYjV92ooGmu4j
/cVv0l11/URd84QMgmURL4mp2MruW2VkhZ3ZBCdAm4ivx0zV08sXfC2aWXpGNunV
MdLpGeIan/vuNu0hYc5E7HOUO4M230nnj+GoIFN5QDU/gc2CCYf1aR2jczV4wXwR
gma/PnDyx+c5wZEIm5AmkgMKWEMYDvO5ThVETQIdfSTIkmSkLfExCrPQIWuREzHN
eR0UfPtfRB4ssziQ+qm3Aenm+6P/5phzYo6uuisiX+k+XsYH8K0TW9lY2LIjIZRZ
A9mNNMr2UMEm2BCK/AikOw30se+w9RJZOjKuJduL6cFiWI1iQddSBkagn/7JyjWG
0Ppgr9eMbh3Kx1iGn/TlI3eqlt3ZCpV1XWz0ZrasdwjmAIdZlQ9DsusnEMcI0jrm
6eaoPFupgvvY2YObxTd3BenS9mV33bitUcq7jyGruA0qFgpEN74NNclr5N9yLCNg
gIkUzCfeeHeNqUPZmjOvS5AWoYlzE2LL/yqBdhWcfalRpiuK3PcPsmNtNtEKg/WM
tEgECfFvgq0Yjy118h6y1U1Ebr7z8VpVdXDOucTjGyqkL5Z3mYTbmk2T+gEPiUvl
k9TblXJqGiy+Wy/dmoCIVORuvszPgTUPlFoyBRLlEfSJkQRdBK28eJQOPgADSxmx
HxhiPwUyQi6UKIl2LAwS28Xx0rngEkUXRSUAtA+mTk8uZUydKKEZQ27DN9J4Ads/
IfBnaKjzpsMktGSVUS1x5ioBvnZbgBuvca+7gVcnThwhm85i/OiwoksOgmB4F3U0
W5HB2TNhI0irNm0edF1xss+VySliC2IwQTd8Z3cf7WOesHbj/yW5rufHMBXBvvat
OIrR7LeiLixPJEfRP9F4hQcMzLUqV2/ZmF1+uuvlHzBtXZICc5tbQ3mPOPBcKcJI
P786E72Qu6g7BsGyGZ+8EiFqhTjlxr1VdOyEoryAKU2KoBmCn0pyfw4DW1oQeWBH
XwYCo+Fq1TtuewBZMNtbLGNiiCM0W9Vo+Qr8WWc3cu3tejwrprE9J3RTPRFScf2o
EqQxNTZ5uewJIOTGZloOrfSMkEYiOLb92GWkJUJyQLlGbSbmx5ihfZQNgy79yUqN
qhcqUkUPntvsq7KBf9PvcctWa/xSsz17VP8iZBJTKpvj4N/kuFZX6QBbZcnwIkfO
n8gSZBbIr5q6954hXBrJBDXG9icvT6wZXS7LMZqBS9d41fwXTFYBuLBpA6LR8Shk
pIJf141kxtqoCMy1WRwQAEnJSo/TS244UvorrQc/B4GTgGDpgP3EPEfr6bhELPhy
BqZPy4L8UrN/WEowG2bkoeXlMTlxiZaeYe3Kla9IBWdMqIiwvurjDT9wxwQL2/I2
hqNQAavtMA7IEBuirM1onAtStlgrU/OMq1YFpH2JUf47E66qVPcTP+iDl5ek4Tpf
4j4234QaaGudv0lTq0si6G+3gNi9KNhPx6cbHbnOoxcc+JTQvA9IO5Eqrh9CMMyF
MSEAKFp9DEHvPyztazSz8lc7TRnYjRNtu+J4W2jLPgvGUHTqC3II2bRaVirPLMBd
Jb8iSTl3EgUZyegGudjTg2tb+MTGPAmnMw91WfFyo1OoGmiQmL4oS8NZbDN70xsY
Yx/CNFJWaWembp4c5rTkusgtIPpQYpFHRdTmFUbbKzrWTSHKvFcSOEe9R6mMgJkg
fcPia1baoiXPRtE5ZqzAh69Wj5E5rts3BBmWzQAVSp7MtKDTBJXQHxXGB1akRRvE
C5EpUI7qc0puByhggG+j6+e8LiS6N2Oe4I4X5MqAh598pbhcw1KGZloQMzxP/hYD
NpV25vbBfZ6jZiB7fvUxVWTdJ12oFsj76xyNOS68rPeBV84LCnTt/64P2yS+EGCE
krvlmnUgqHfq3pGh2k4+n3cn8VS32wAq+pq/L8yT+YXe9CZ3BBk+nwzB2dB6hjc5
JU2xR+lG/FsmRWiTy1OdKGugOWFim5xJtNPNbJ8w9KRVInw1dMuDs1Q1rh0xiA25
bi+U40jPqqQltg8pnBCCkfM+pheSpJ9Uhu1Ja9X6F5Y+gad1rYIaY0Q+k1c7Z+V0
53hLOQQQzWZj6yIjdI3W2Ye0LYxpNwMnCI7BzetQHht/p1PbwPslkPIKUZTXLqep
KliKfSEl1TuUVcRCEpWKCznRWFqgMAHrXZeSyghv7d+Nuuzg4wR2jvtByjOdZ1XV
EHczhQaCScjfo0+k3odMa9ABD+LvhNW5R8J5pqcMRMdursOR0Ku1x4lzJ63WJwmh
1nvn3nN8B51cWNCWD+lLX4r75KfYGlOkN67Ig2OPQZ4xhdORRgxA66PzyYw74LZm
tKLf6rMVOEwUW3CC5zBeGSrM5akreCM2cui9O3OszBBMjC+d+5bn4+H5NsegTOzl
5JtkU12WSIazenRavVThScT3Z9/Wjwi6i8J2ewu5mSGkuSzHLEj41SdoQ5zDMtq2
yhT0vjC0LGZMwDbOiz9vPXTTvvEZEKDMIUY65TPYCapK5FR4VpirWQteZ7vY9l0P
robOBfFNUcdtzgzJJsNNeX7a9w4ugtqf4lS92tHm151NjJUigjlaa6mTGINKU8dB
qLuPt/uU1FrLggN345tUbBsiRowNLxiWZrGI7m2Kdx08aeyBwPWbau4CSMM/JMME
PhL6VTDITMSJQ9m2xx8X4QySEhSsctl/jYed4ZHjMLPFPQTHZIOvJEk3Fo9Nnkub
muKikxTP49bOK4XWfTrocwIU8ff9vCUJscguBQ3UceCa3shIYYL1BT4qnF1qbOuw
6OzkeM/i0QPvW6XoGPDTC3KZ8ylfVK1X6dyqr6iazx7j3y4H0et0YC8dUr59QbtH
tLFEcIbMyUzDkB6IyKlLM7LOpb1Th/vD1VroQi7giO37UhCPvgm5MrylpSA4kPyV
W4xMs0eQozA59Vh50f6r1JpzBQLsCOqizm/nH7Ps8ZGpzSAxjsaDJBN1SIHzLbNu
KCPHuwh9of97GJHQ8GrqQ78t8E3cZLPkFXYSSphA0DuHOSRUPkFx5oGoWMg/AaNF
djc/hT9uQUUSIfx2X04Xt5eGQF9M5GUY1ROtUroRpvs8ZSX2IFZcg+pOgUb7zHt2
fteZoVC8tG0BKprCQCYim/fjtqYZ6CnyfqGsOrsbEP8gDjTyBd13YDXmvkOswSUQ
pf888qy0pWkCmpU8LwlsSNxF1yMvTeHDh0lw6IQd/d7ByZ99gZ6l+9Ysh3gbv+24
QgldGgIEhW/HPmI+MpO6Cir1eiIBofzXDQNls4IyXikiGJ5NvDgpLbrWp/Ps0Xzr
hPLCvspFiW7rsAyawf1fD3R4zIcsZiXN5qVdPbm+ia/y4Dt8ie51WNhk/IPgvKdL
t7p1O9eA+3I762bsgrLBZdDS4RCi1EuQE7T03FI3EhqHJC6QVSOWibgO3Md7otXf
1m0uvPdhp6QRKReSrvjqk0VWqNVFfktybP1TBEggPEsXfgw0hoQRLCSXSjr6/wVk
XttvPil/eBogOFgX4smTXVwoVvxPcCHijbdwmgbHts/qJDGZUy8oMpWs4oRqM5Em
QZ+WWJdyBVegJm3TfLSV9Q6HwDzUAwwpqCW9PaJkWwlhlllswKqksqOOEBUAsL2S
GCgeG4JOu5cnERdYJ1QJbRLy15XlGRLs+WvDxrcKo2lII3Ogp8l637g7mNSEke38
iNbWGSZftoNXM1GHiJrIyvd3989eDxMETg/NS++FiwwEfYCYyujZBTQHyGORA4YU
bGYQ46Z5xB8l2VAeGDyTsg/7LUUv8evNoXkg86mVO7S+NHMnuCcSfUD25PQ/Rnf+
UZS74MHCxXjubu5KUa7757Gz/MyQc+06ST8B7nfLGpCPKlOWCn32F50NzMX3RYIz
TQFWR4qcKkb/3mhYhyNQW5KdHJvKGdJ4FigQV4x/nq8hBha87x5Zi9MQWW3jPXr0
3HGNgA3bydNh+R1Sj6+RE8wdp3e2qBQU668//cYfuBgoeEprbwwkJWJ1y8pYYKVo
O8XbPmM+LuTNrrJCPs+bsAC7F5q5a/E2G/2RF19Eocsu34bxlcT/x44/m2WpgrXU
3cBB/Yu1REiaMXfFJqy4zluVx1b+UmS+wR5RS1o4c4/CSl93g9GBWwNBjsue7g4G
aTco5IFQIsOTQ/+K6xYso/2HE5awU54kaOkhrEO5DqVLtJX+HCBwesNtHVcYYxjI
Se6yn5CzmwMhfdhIThPf4skEr9IWMWax5nECajmFu2KjKPkSZDrWAmXfM8i61Kux
JLsUOduO2O2MtZCDDPCRIV/uIxruMveAnc4rmRMsQ1PpJ2F+Hj98sXWyNLpz7BS4
BSMOmMh5OGDux/EhAVo03Ld1xwcJXtDgfDSiBZWV/Tvx/dDJr77YaX/WcKNJ36Xf
psdvBTqfzQJ51GCV3ZCTyQ0Fxl9FBCkjRwyvRwH0LMGhSGk2Rnlgr7o6zgxKS/W/
CF7zO0Z9YrNY4jdqr7XT8k71LTgloV2d08XSCNEuae8zASMMhjjfKS56J468skvm
DAZtnGvRIVRUixCJLVFLUYNFV9Lvqhbqa0EyNy078v/CC9DXjgwUt8rlZVAVBJxa
qH19za9jXmydGE9Djq3Osp6J5jVX0Rx+gvDjOihg5HUWO3mIgoPuXIOlP1sUhEKh
KW5XIcSXB0+x6m8H+G5aEYMk25jRDocaWEx0OSlnGPOTXwaC1YUhUVihun5CiB76
cbwrDRBwXI8Bl32/1UkWieqqRB2m4FCD/jLoNQzm/INcdVg5YoyXd3UgsIBFRHi8
APXocA8i/8ApVoqS/u/S7ORLFz/qAlGLnfDhPTk/+eN6w8hs57JAiNzd+wFYYdgZ
A32DQnrnQZHNu38fqzqKBAZ2YUVlPGXyhQ377f/RYzAQDZ6KFTF6w4bFmantL8ic
Eu96vHEDqQcFEPYtTN29rB5+H4dEzwO8sl5N2nR+1xNc3TzWn+kh7weOjtIutNdo
SyfT1WGaglb/WUyvtxH8WPUepmLYTxbKiLlRm8vcSB/XRQRiCBdqF86u9HskvO8j
sWovaw7mu0eykMXtTKflcBk4jnd0ol8E12B8P3YHkbOqQgK7GJ0UBjv9ZQUNb3BS
RWarBkbfNEWBvZAInjn3ACejzl8tW4vn2CgTwhaAnxW+lv8MkOIwtBj+Yasy8jRF
5l4BhCLtg0PGvpuNPTOwexwsjr1nzIO9KFmsA2BXK7zOG1bt3psRGZMN4+5yQpYU
wa38U5t278ldvkATiDiL6eXS0f5g09TX8fG7UEG0dTCdFTqkG9ykT1VUM72+fvn5
Mn4bud1PfcW2rtrr1mSbTo1fxyHE4TAU7Asyy0ASr21wt4bzkAG7ETZBb4mkw3ZW
0klakizZvKoODnKDdqcuDGUsq5LdvYTBDf1eIUIIN+1XUUEnxUB5PUJ2UhOaDtj0
JmPiliafk3/3RIFPvlvEFG+WkyjXm4LwRHfPD6KTQX+mqmMPbp96Bx/t07u5lAjo
fA9VFZXZYYoIQCleGNcCHFDbVratkOVQxnE9mGYuyzweCIcVUj0P/1WDKsXbg50E
+24Fs2Z2ogVmEXtwROWZqBdmZjcoG69fJnXlTx5lBETRTdptPQOtqnp8J8M9iD4S
RNTO3pIEvd0WsG4nhG7awFl8lECK2i9IJIhs3uaAiT6cI4dob9asAbZ1qFpKe+o+
kJu/De1AFqRsLy4ibjxm4xspCizWPhBvjHSNOF83swFehBwkwLDPMTG4IDkcK5Zu
bIFYpCqI+6svPXj3/4vxCIsGWxBAOa4uEaZNOpe7QYb5ibgU9HLlkaAB7GLjvdff
iza0gT2Hj3UF3Ny5/zrYYYyGWTV17lVNbIj68UXPkKdtttQregYmGBBawk5DJgQt
tUSS9JIj6yzJSouMH0wE3PsL3gPA9YXb7GR4d1Nn0lyqZbp9qzO5TaMwnoYWmTaZ
DVyNA6hTD5dAmlDfraU+UZFRcDueeeW0DkqsmuNv40kJxM7waiQ3HP0ZVQvQE5wU
xolLmUwAOtRLxQ7EZ3KwpRlOpRRQhbc9cUmXN3BQjO+pczS30YbqIc353friLaM7
I4fsX6Xc03pN6ESqaOjN0vcOnKrkB0oSssmwtnC6E2aWxifGe5Pl6jM38NPgOiv7
vYhlHagAL56dpQJJtsmMOBVwP4fQrHmmwI7zxpdn3F2OTqlncHzaC13JUjfv8cfV
9HRE/rlPfiokljkA3hcejXanFN0Nm28V17THzlBzGLC6TNvno3DuUnPr+7yF9mjA
Zvuj4cXDWaR6yps7TgjAv9HHP2u3xziQla4m0cntwlq6fcxywLVrNtMnfoJO4s5/
yPFlTZpuOmozxo8eJsAjyZOPfza5leOyj31tKeCcG4Fs7kjGRKU4eJwC5q67/mCQ
RdxmkHVKHIjknb4EAw+0tBOK77rKN0xyj1gNRaYeTNWlxZ5k0aKgQoRlTqDnJCrk
GcfHx26cW47G5FnDUDp6vNb5IfHejX0AL2dfiZel1NnPBvmDAuGikbttN4IL3HQp
o63AasH3aEImJrdD7bLtAtIBOOGGVIQ34rYZJJsk+44dHecf7UinpV0Kgx5/gJhW
/u1wj7w+61lIroQEGuMMjpzbuXxNW75LTVGYQoyRou8kpPy24SSiNfBBGZDFIxO1
iJud7tUx0nyXPxLZL0PaWYCz1CEE6ftiZOZyu+Q3FsU+ZfclIv7nFcIy+gRzJzJA
Z6fImyNiHdqyqDLsaqe7W0E0jWjubFDTp1G64fOwOM1Rniq4EMLRLrSgCDjn1DLE
ceSY1vAAUUFVilUfSxY4YgNqBWbsIA3nu1c/IqJsbcYNhPYaTd23I5uvc/DbYPDe
+Gi/FcII0wK1gYYz05mv3wj/k3htcAQjgf61MnS52olAGyVxM8DkjeXPPun3t9f6
hAtUCjbZ51/eJo/SDUAjxBMgSjBCLkziTCPGfjxdzYtMtAZHx7DVgVm3KrG3N89X
UzNnTgO4zFzdzXRYMm20Lzoy3KqHDh5hmq8QmDsWN11SJ+WvNz7nXHQ7AT1GpsRM
PrwLP5aTK4aSTmnpKWtbQ+g0rTdmQSXxJE0bb9TnStGvajORTyxfhEBNKRMvOd/b
4a5TXTdakUrRoetOfLYjQkoAZjTe+AKLnGHleXQYESUqP4Vt8BGnZ7m7sPcKiKlH
B7rUYQPzNMktmwxsBkaSNx7ruEF5FjmzDxklGP/iRcVfrJJIlrmGUFt3HXUuzfVL
CNyHEnrzzVu96TtXe52fCG4wIDsygfY+UqwKSLAi2Pjz9o6H1LVd6DwlUfTH1/qW
yPUMYAMSAcY/WIeXW+AndYj0uZOGdhwO+v2dnH3JlvNsKXH8L8G8cvEsb4wVnaEa
Tosmf2/rk/Qb7yPy2zZMhj//0nmwbgrMVZxeyia3sb8xZg/n+h7EAF8UZLwEhhwj
B0Y20gF4M8QWVcg4GvxyYoTcUNHp/MrZjKXNqAYNAtSd3VBIfoeIFsep/aTuxQjJ
9vDaA6nlueZF+uQyTO75uIOCe9ppVBpYMMqDmBwyzgD8uxfj5ql+NpSxBlDRoeNt
h89aRE74vVzQJO2pfmanRTF2lZXLIIFpleGHERAkP5Fo5KRdAhgql+Q2uYCiGDYI
4koa+fznyzJq3Mz/5hi0nDhJ9LZ9dIBts2rcULmTUAUckE2TiIdMwAcnTAddPnVc
8T8yNXcxJr7u0AO2M6y/JCEDhGAk2UhCujmdUnpwp3ZHmA5CDhZVZ7n5iQ4APiAA
SoOiLT8dovvN6Q9rwopLc2E6kLsc8LMJoA9PHL0C/JGyBHR0rephyChAu7BogQLU
mPrz3hXexpzhPtjnwDmEmTBqmBxtkKt6jKN5kFAKWQdf9PnbUIvvPxZqXv9eh/g7
O6fYJ/LFQnnGIJoKeGwpnHSDFlXwRrPsixw9F3/KidOu2iTMgYXseitHrzFCsGfK
jxFJnJ/lNUGleGfus5KlLWjP9U1jyhQSLUC7qeoOZA9UiObob9FpKakonEwdpVlG
zjJchoa8a1mhESStr6uMzf2PFIzvOl9YR359o40Q/civznR9qwjSFYoGwTF8IHgv
3E0wn9QV+1873/1p8z7Fm8phsYw6VmSxZWGloglV/Sg6vp7Mmnlvf1P7yzLOhyct
7vnI0ecOOjAHkcQZG7KPniv3pBvWMq7DCVGm+8ser02MUoBWBW66tVK47RPM53s2
mz+t14HG+uhTwkxtivY2kWpt84mcNLrqIcVfCzn2YNRRx1f0c9NFaEw5vEL8a/rB
QFXqfDn4XZ4OUKWBahCa5taqm8Z+XOICOoOpVnwqHzmXen7UG56Z0//XIEdqhD0N
QWtjDMJtf79jpcEvd58emGZgkm79lcjSiikzMhb4piuM8Nx9HDgXDrFlB/Vv3Aev
0kElupcId3nIP2kFvfiGqk9Aby3nn3WN5VtGyJUSdbXJ17+ODYNWlig52LI5rTbi
CorYLTTkBUHj+qPJxJUJjMHKNdoYMAhfPrBcAtRAIp78SaUAi2ofeOAMIJoHnmho
Y6+OsLJYbqx+2sC8oW8ZuUaaPXkeuwaasM+hgcqcUuij2GDxOcW65X3996SEqT5W
ljf9bboH3oyiOGr52ARL/OcgapVd+F5NRSnowurw8h6VUHbKDlq6OBdiBUdjfuau
j4OqV4z+UF/MkO25XoBLfqikiKKEC1ffB1i0mVps/VEbNT9nKiD2eb7x8YTD54Eb
OOCyeMD1wJKDab5ICpDh4AyqGmz29Nl0rrHAlQv1PtYA4d/Hrhypj0lvYbvc4K+/
OUTazQUpeS0SWzHhOo2y1kQd2BCeQkIAAt5jlAu288O891Mmsc4dIidnDhh6yNMs
crN6xEnZ9A35bED2zBvoJgRS212qBmV+S3x1ewyUfULdTRSQ7XTQ7yudjlo2CRqy
Ni6V7Lzklb1ttdqZTBP+Li5rRzUp47ePZyKjZAqECRH+XAGtITmfy5h4f7HWfUzJ
h0Bvat8FULaoTJvdYAimoSWTLD+bJ9nomHB5G4PSf34uLwrMdI6YX4ms7KE2xb2S
pKVcdj19Dxyv+wCALD50yfvfwX4zKxsq04hu6Br6PlQmaibKUx2MIuyWz43IvXYl
zCfNwdK0vMpo7wfW1cjOyaIVkBuqBzbqP41mFWWQvaT5amTFgfgErDRdundOpBxq
SWp0M8gkL1KlsIhJVLPBhGUk/mbA2SRcf0q9ls/9/j364jL421D7pMYSYaIHk8ew
ryVoXqJSoX7iCiwZ/HOMniSYb0A1hBFpq4pPg+70aPjvJ9mP+xf5Wgz0DjsSa+Bt
R0HzbS7bKTdJ21nZB5AlKZolVwNhVYGrmkHr+JDFbX6KbMuFQw78CGF1ZHSPibSl
WajHrPWLnPRTb3+xyWyGhLMaCAziQzAf3eAg1jd3o2o37ld4EfBcYkG3J6+qAjMR
KDSa1fSs8kZid9XSWmic/feIrA4BdMbmWPwhtwGangS+TgFdAcWkD1ruvoJKKaaw
VBum1sU14TOAbvKnRaGjGAonJXHdiA/HAl3Z6i7YtwSRXsYWBzHtrkcMeHhhZZjz
Lpvr2oswC8v8wvN+RnvTZYvYeNid9MVEWgfg6tJOYHNtI2uIG4SWkVLzWuKQ6JEl
362o+VTE8IiG9TjG/tZ1NoFw42n1BI4bT9RmoodC/2JylLvYThqYfYFbFI2gn5mm
gqNlM8D5E0BQcvL7VkzItHnQCo197R9bZH5NbmRzbQzDSpbKCMRdwdM3H9T+Qrqu
LFUvBZO2lc0W3tITWzJ+KcfoKPRLjyXeB4odWhqyKqzfYdl1QXoBbY1pklR+Id8N
LUELSD97RjY7a+Eg0dHye2icapLAK4wHzIPNtuRhKfrGg1iR434OKCUOD6eiZFA+
eozfpvw7x1zqq+hMlJDWCqtL+94fhIOVmjaa/81ffvig8pUD6TkVOgajXegrObZt
bqDv7Inhi4bOS5rWJ5l/6c6XsolO74BFPrNFLPhZVZMALvt77lnWGn72WHvwi27i
4KcHrOvxm/BtvCqphS4oI/j6Wm9hlJZsta7yhJjeQ1GyKR5Qae/8pp3ZiQGcPyAz
Ljcoo2oVRMQFBcEplyh29sG2ui9ewU5vT30tTaqrQLXAz5F8BTcqCT8VfMEdO89C
qPCSw/K/bPVbad0bWrgh6fzEiLbF7YTkGQVq0x8Nn7czncLyAdIgwPBDhdrkFKv+
jhXjoY5EbqCF1DAnXjRLpURMLiyNkaHoRIEoWdv1hYBnhdHc3yWiNUb5IXh7smOj
tQjGUIOjROj7baIJErbw/I0LwHbFVkRJ1kaGUGefLDRR7UYT/ykIhsSHOuEfoU7m
3qQJxKm7Sw5WhHYMo+gj974buXi9StwR/eBTbfC//RxeSFPOYEWoxW8Gcjyk+XVO
IcWA9EwnTbfPC/1syA7BGZUWRiQzua6tGWn7JFhfbcOE/pyCjsxZXPcVIiL2f0f/
QJVq65Gc7ldqBo07w/Z6yYmfs/8CPytMeslSXbYaJOFYxOOLoDMYvUZFfHjnZapP
5vYSr6Ns3mS6yIUj37uJoidBqJYE0u8GJR72oAlbIrQsHCVoMxQ/Tw/XAkgGkfa8
BJKr9Zj0xVE0JoBkwiqeXzXCKtl36Xbc4q8TNNigDHiUvunlSiSFMqNNbeaDxKWx
Ig1B9ujuadfk4cB1SGG5JonK9iVWtLTne0wf+kkGZYVtEkNyt8CnHpKDyV9fsGaI
Rlqag3yTRqQbf9NpLRio1QHgfUIVE4H9ln+2Co+8Ngo7YM05WLYntI5A2MagqQJ0
HENGAsZtgEIW1B8TLatGS/V9M6jSWRy5B24DjYv2EZjXC/s2Or5UmUmp0mRt9zvc
s8iqhJbS6cc7/TpIgmSFFlhnmaouqmmhxKmEMun0SfsEccKePvIQXg1wuxaszkQ5
hDNOgOc/hD2VHKckDJpTIJ24Gz1vH7nlTH05H51NGNTl9ZVTyvLWbJ0IL8EqvwBr
pBiS6o0sFRJiVpKZ2D4kMM6/USRI0dPc2JWbZXmZ4WtMsrsD98gBaPnFSCjvx5jw
j5RRkd363d/T5h4jAkX9QbnZPZ3BFQKTqUkzv1kHxTGDfipBo611uDNmoaUhtyfU
hv10QrvKm5Nr3GN20Pvv711XXzLTJzTXsDe4tkYQPJW5lfhaknvWWgf/vh9Xq7yA
xXXVBf32mN/5oAkm43TasTVD0yzS8Nqz3QQdQ7IocJIUWibDsStQor/ZBzW6JJvT
S2y7JHYC9iOre3hm5iPv1nursEmxVVq2mBq379rhhHJ4MuUENLCYbaMYP8Ebg4Gw
hHrEoj0BCT60PWQI+nRsrGz45crGyCd9ZodTn4JjV+oFS7WMLZ8GtQpvOvmp4VIs
3FiuWaQVtBW0nyrGPMq9jiRo84FFLO75FTOLUOWUSo18t598DbkwLRH1gFIiTfdY
l0NloIAgLEbL52eEi+wwEKM8oDo5BpdJ025aTQixwpXJ2pMHXlu3Xgyq51nOF0tZ
gwWjuaDOhwz6zvnR+rnbsBtuOmPYfs5IdIBidFAvcTC+kygWCa4V1+r0PjxorEw2
qS0XSeVmK4QAjJA1xVZDC1B/JfEXgHFdR+bb7NVTENyakgGYoK/qCDdKdi6kMW0q
efyBE1hT9fnywVShkg2OK1DFKveuFmwSyOpEA0v21GsO23pOHSeNLJ6lFqN/42H2
O88p4AUUB5PaLpERYY6IoPtNjw1hRp2JInDe402BVxCduwhhrHSyUC09MWA9Muq2
yaZlsmWWWocQAVpNyMqxFML7AOv9fb5zYPCtQ0tjNqWeUczx+wvrAu5ZGQD32cwt
OyiUVJPZZydfCorMuTSePJx9z5q8gWE/wiDsZQGsDEr1z/1B1g1uLSYQHa4ZAipG
kiyFRtH7ZF9EzNEYWoKywvrN2XPsBCBmFUXV0/d0/9suh+aKivChIyHzVWAW83su
l+gIt0yvkMV5+JsIR/P5CsgEAfc+ODooO8VZMvey7ntCMNFNCN7vrAZBzz+Pgtei
y1uHgCmS0q19gRxrI8a0KHmz3SCZIx3w4rLW9fjma1WA9dDwysRXL/WCfa9mI83l
GxmvgtKztpbY0+mB1uxoxNDT6A1kBCByx5qpd3B5msrAAvJMgI269O9HceTQCoRq
HKp38iOmQVm8/m+l9oz+as5LMuIZI3R3E3kZxerFvit4rGghvNTJIkdmEDThB18G
SVZD1urGEkiOG/mQBXfLeXFGKoPhGrzbh8s+WeemnkY3RT1Hqml69Vr8ftlg5ALt
OS0NtDCf0T1YvKWnzvyXsQhsc6uQpHLTUj0SmsYav5HcY4ZlyrqhMvD2I4a6qLln
wKxGKEgLt3o7KVMO2twyO3AGSMP+c8kJ5zGczikimnU2CJzoKiiUSN3D1DVzAOqx
HlcYJB+0H67qXlB3a1RoLoK2pXmdHbkZdxIJrKEizcy+rTSMPpCat9UCV4AZZHdO
5BcCbw1e4HggKMvgjq29xkIlY3rp4EMEQncbQgYIi+58YJT42zv3nzYxpE6gs1Wn
UpPYXZIoDbfirVaCLPdbIgk0klvonj0mO4qISMkoQlYvM3/XQtuv6Vvm+D48Q1aF
6kemZqLPGlQ+yK7fXCmm7PaSWb3jvd9lXeETMy5b3VkG7t+cQAn9+ZR6gONptle8
UnTZRSYtKzZRdBAR34xLgDUVv8Os1+a81Q1iMI5gfcyg+6eXEe8bMXRwN2p0VxL3
bbwX+Hp2o9avoGzsPX1bl8NwKBQ1aD3Sv3x2VfS5w7LByqlgw6w8D9B3q2R2Rb4r
fKWyDRgRL9Sgnkitx1ZOcb6qhDR+fuPIOhkMHYpiUnLbSpwB/LbwOgFLxV2vQsP0
huR3S68QcSI7BvaOgWgB/nN9NJEmoqxY6guCduKEg93iUWaBE316ci6ORhvTzeZ5
xfjwhoKOhAeQPhHDtRjxe9dloPIB1VWttoqPQiV12My9J5inh7zqmTF0YLgo6Qud
JcPRuL/XP+NjIE4q05f6xoZL41AXHMy+sEsPEIrAv1BtRfhHHDxSzH1GscOBnorg
MnCAE21VGYh09NFcKXZeqhYHG3f6fhlAEKJItEhXtNeBZXu5ynuuTv821RXWZKZ/
CwjGYz/z+byV17rYGJzS+0nIe6Muu8VvytxQGS5ey1kVr2X/fJDglR0/20MlNSsG
DUWzd+vUdx0pUM4e8IIfoBMbciYpeE4I/ed6Mo1wY23GXANG7I35Bi41dMckeext
MEfneUKoxuyypVxdN5qzKkn44Au+awf79AT98AXPFxaZbEk9dIO6G+SYxETAnTKa
39kbvnsgWEl9rKO1FNI6XxKYioqgl0/mVC3j7jX5kxRa8FpLqHrebBcURH7wM0bl
FcA7Uf3744QK3l0GsXaFWz6MnU9RPPu2apHr1bg6Szhbd36buR28F2kKSLmSUbyJ
JI/woU0M7UBEs1J4IwEjbXQlL7dOaTZhRQRC4MRKcNCVqGLNwmyFEoCrYmyK5JXU
7pdqd4Y9SsvugcZMer0reuAsz4pvzQ6ClCmgfhq+LDYYL3X+SG5qtHHr9ddWoZUE
hWx58Wk0j597yxh7xR9CAmYOw3uRwxo4dhVejitHfwRAMALqWt6jc6Z4kACAa3Io
yQD9zaDaBhgw/JbvxXKGZyizawBqS0SdMGM7kINTLfMQiIasM3TGSx8nQU7ykRmO
zqJCFbK5qtg4SATRxEbwO2p7MyWHSVwwvQ3WPlFgxB4fuTM1T+XafaY4++1cAjF2
8KvYXaPAAczhcdn6S6qPZaztk9WulPOncCNgK1KWN8vlhRdl7527ETkdETdwc//8
ydHAy7984+N0C7qkP9vbRpj/TlYxc3q3ks/YmITLdFiiOYApNZfdtQN0XPWreeg/
95itB/g6hAJNJm7O0y/Rr9/vt8c8hc5if+LjaDQVI7wVnq/XXh6QtIqF+854BPPg
YqwPwSn+WJ0ENOTGDgeqf7uW32QPOXXttF7FTqfwd1SngvelylE0j1DbQpHaYpRA
kjOQlDgu2Yj0AWjooigrdFNp0ztKg1sEaO1eOi26Iz6I6+qN5QCuh85n1dkGB7cC
P6eEeqff/nlMRbhCXY74bbmX6L4ZaZ8pL4rpG/mqkgVT20WZ60htL3Wu8Ucz1l9u
h+ss1kDh2YsoZji/SnFIBbWHVz3JkUJEI0SBVyMxx6sBSpim7KeQzQfXjZkVW59v
Y/h+mZsyjkHoZfgaR6kt2Erd6+4XPQPhHQXfsAWeSankF7pCAxYv46KzK/P+EMOq
NUxUCRtCo1CK0tg9LxHUkrzZp/hxhMgXsN1fkpwjGTwNSofB9it+lvtCVvaaJoVa
vbHU91lcSKkDbIh69RkiCmsKkAtAEtAKTdQlS/mKM9CQ60wXgne+wAzQNF5fd+6v
xDgIaxXDRfycNfIr3LVkLxAGOzpvonhElKM4KFmNCasK0NPjtM0tui7e1tPwwFUK
qZN2NSaeEluzNHhB3vqnQ8uN+rSndp+p+g00nd73cXSudaDA0k5W+OFuCzNWDB83
hC3oxG4FawWsrE7Q8D4bf7JeBG1cwuAS5mnQGgm14FveeFmn8ET3vWdesWg5ZNg9
ThIL1Mk6Mshw3LjWtrx+2aayzdYMnodtN3ohUFkmBDY3TcxsMmElJaWmIk3BkjZD
IiZI4gqpEgVdmOdQCykdttqdjRBPGkcaXYjVdXe6hGO8opQI9V6KGQ6EtMmwEUzA
g5XLNpIJGiNV//kTp3NUcdwYz4I1KLx+wFNM/lAjn0G5euDamoG/PiH3RYecOeUO
Q9Z4TvsKx8o/ElSA3rCyjcVmro4TE2tgen5pA77PAql3vfUsSzdhiSB0fRhmh3mh
otNfcD8fVVa53sHEMn7M6rygXaXa60JJBsojmBr3Y9Y4+eWgwU4nCdxs8D8BtT1V
hJWEUI+/6chDA6NGXArGFk6HLvmq/aTQJFs7Q1aJ5onSTDdPs5IN62jaQTrwm28j
ftcqUpvLShluqYKGKCrkwC+FQqc0jPF82iRh+MXRwFRT4ISJbd3zm9+80gBTmehc
Qk46H3gg4Jd9XsfcniHRx93MV4jy++3hXTxgoFrhNceUWxkRCyQiPy2ZQ/QSJy1b
kBL9Potfxc7CAudUT5m+/ETAoMwMhY6LLqiC+/WfkoyHrkLEVNeSoepwkdJZtDHO
b/25BJL97zF/iTqL0M5JrSi/ICZZoPAHxxLozLWEtKbiJjxRwHlc2+IDbGlU3VeN
gANu7pjsIRE0c0S8aW7UV6+69fD/XlgJ5uk5MmoYkB+KaxSZ2EyOFjJ1ej0nupqH
nMb8aG8pzLWxyltfr0eHNEcMj1/YpD0V+5YDe+oqiT6MrKcTJLwpfj86GdQ26B8H
NeDMZZ6Qz79ubrExhVSy5S/XI3p+RuQjyGv6lxSstVANCL4ikUpDV1DFKlNW6Xul
oEg5Ur/pFE0VrvSE/rNQpNkW5puHse3iRATr0I1ntJXEF5fqY4DkzNiBV02YibQ7
qz7hIifThvcHusw6n1zL04cPrEyMR1GuBq/UXcBNPscLjUY6PTMdY9rvoDcZaeew
rfuA2pGiYfOYItONB9GP7p2hZJgzNElFEQv0jSCz/2LnhqiIy0cE7OYLB3ZufL5n
vtM99ko5mKLW91JuqPIkRYhHjlkcTBGI9EcEmYis5wRE+vODcGHsNkgzdddVWzfr
YdzmlIyzSx2kGaixL3LY8NVLjPrnvIzW+6agUkhhW2FV+btQGve/pkatNK6ykPEh
O21eW/zk2W4ESp504IefXjg9AbcQ9BN5uO36+TY7PBimxvum5vu81aEg81bcc8UV
5wAkKVdQsRcppQkmvZMmxASiIOWOqFOgkW1RXl095T2z936s4x9ztkyf6ODjr3in
n619G6iM5uZfFS/yeaApGQjUWMUf+MoJJ1T4e2+1xNzhj0NLGj+tl5QijFxuy5cr
O8b6lNGhxd3gLQMJ0qh3qRi202DaC4sG2798s7louFZ36ohB3k1MkqfqlDdbKxcJ
FtqQ02i7TOM4xyH+SRnUTJ7SfhQKbUx32ms9vRt+PcJ4AXQgw3LvxCj0wFsJR4B/
5Nt21WB1T+Fml+I8R25su7EMndL8EtIiAiMVK0vtcMxzKWyVqS24+qNJN0Bd2pAv
Qvk+BUwhmdvsm1V1jnRUR/lk2BhDBFKF1Zumn8Lc1a9Jmmy5nHpWSYb55t7k0LPw
WQvkDebgWkrURiYZPqig6uo/ytkmR4iZm1EEHaculKqFV06K4C4fS4/itSohAklY
TI8GvQGL1qSF9Y/vh8JFm6m/9jMtsi32M3s3RfUomsiHFJT5MmECJHhKoHrQMJvc
4sfQECq7lFstKOnH9Z1+kuCaOg2KLSFkybqQWtbmJMuvGJWxlT9GoMcvW2uXpreb
MKIxOoZhVj1oDf6Y2P07rB1i0Sl55+b+dwRB5yjFm2lGpHXbT4kMZ84fWPeafbK0
M1VZtpABseY1kabAa2H06KnS9Qz7otqA27Z0Mu3XSm/M8YCMZZU2NWnHb2HK/95d
usjSwK+z8HNssOUHxkiglQHUThQciKoBo5raVXtT89ulDYWRilGcXc35yTfcrjOU
Or3u4+qEGDrgwyFZ31QI42EGRzJTJtaul3NMzfJ73tgTRy6n1OQTO2muvan6Xsoe
HNZcmCDboooXx8vZMxKYn6+ZGTA1CcDW3rvSOqjRwQSxE9zWTsQ4IEPsidC8yYC/
5w9to6otK5lK9Sx5R+e2/V2It5boQqBTfRAYas+a14PnUMye1ckN2DXVpjA8IrxR
XhSUYnByMdPf4gz+ZDAgZJBpRQ2Gf78hIGEx9tUcuOGEDR6qghgWB5njOI1dJ8Gl
Tul/kPLrMLPI5hBFAU63KRs/Ph9/Sz4bcl9Ip2nBwqEL4DRTIDo0GlIdavd086DX
icL7VwCzFUoBXtI4Bz9EWkdFoMXKX/dFMKb+LQsGnDuPY5w5rQ5z+mjZDvJOhtXg
8a132tQjVv8wJqN07IySPcH+gcfKen9buKYXv1g5X+6CctQINhI+MzPQhBnNJ0Hw
EEE9BZ+VYObsn9lwcxae2RGR9BCVTvdtWlKclZ7AE68nzPz75kUffJ4msh5IaUC/
QYVx4/2Xe2zJvDMQL7caYFVX5OkFgZ2jikd8aafo0cNgx95djheAiUZYuF5gcK7u
CLtq27pHGEWnvl/1O/zN0BBw3rhzJoCdaUplS/TU4D5vXRGUbyQmLyxCQY8hu1jH
s2M0JAtlB2ZqUa+ComYMfV41lOxHIlQudov9rEj4jAt8PoNLuMCVx0uHLJE2B2aQ
mqGjhCHHNEtNKfGb5P+XDsDW1z7H7k+YK/JPB+ss+7OlfeMrmKHYOMmsY9dPGI/a
abobT6183ozedFOVZodwUu8h09rqYWo7Uh0FU0G1nluNlAIhl+17bUpbnR5kzA4D
rGbcFpB7pvw6H8uIhn7OPXcxm2z9go1Zx0Cei/p1rr7dTB922OW4NVrVQJp2GXKN
cjoTNcXxk+NnWCWpeyzLtLYPS5oBuqQrRpiSN6VNmlZrkc98nVyzgmarD3edB/Uv
LKjkCY8UHXrfb58RoqamAbaBEdAbGUYIOiEJYxJ7cjvdq24OZF1Yp1Pm0j1ZaDn+
64amQqHSuQX1hfUmJvUXKvFPEQ25qo6PzkWxoGIsP+JOQXGzCu5sbemSNjICT4s7
+xKuWfsi27HUgCySRQQVu48/Ro/7yUuY1E3yWEbiWap8FeNd79hXcP5xHfyTqxhq
0HS5otUxE4UwniLqwxPjhzSt1McuAwFmufvg1b7aaV/V/UJ5tqpD2RXaTbpcm6CH
V+Yg1pMw2BSbup6BQgAQqPs0xTFb2Ch1wnk52TzJ0uHDl2JoQAuRYnbx8I6l8NCk
0v7/Zo5GUjXfpVjgaTWMKMztLWCeASIJAz5D4ikieDic2IruoUsiN7WH5ym1FFLD
kwojV62VBaURrKPLJxTW06O7ixeAS+/BZ5POSYYD363tIyg4osOP5+/VP4qJbF6H
4TEZKs7A7KSghwCJ564HM2VWex4H8z8yNf3gKDxp54SVFexKN2NgJS4ne9n1S75T
6hu0lMVeHq/41rO8FMkZImojHEOtVzdqHxfJuzBglf9zo50EEH/9pCRXNFB5AACf
FyizFqBPyKa7JiXOLvVIQM3uGtRJtDPyCAOOCVE8ucWWrAskxfn1hdREb1Zsg2VJ
LN3gbcy5abcvpsIi3fiQ6ZxsluWBD6i+7eW4py8fd1oJ16IsozyhRFBCo49XFkjc
+gqIPChacoLu3Dwkq6MDC5fqbySv3+7T5GlbKQL1rJRQtVrwOE1iXCKqpmH3iXFv
fkd8ryibQR8WK/VntNtXfFyts+f5r2FbAaiHPK1xTPgtfooswlDJYgNQcqX8b2En
q3TRn20ofx1P/nyIlE2nf0jHLPxrvWfP6DFyf/9UOKY9jBNoZs/TcLSeE1I1nhu0
1xuXbz+zhTct3rw2CYVtw/JAyiKqwFWxPUCWaKEbIt82h9lEBmN41WQPp+b+VH16
qklBjY5gYTs8ZQak60xZkrNKW8u4ERO0ZgtuZFCvpAVmbc0BxcTbt3M/iq756zTY
rCZqFVvhXch/kftfRq6LUkIpo0gmHBT/D+C6M32iaur/iHgenXHAjiY7KMARwMZ6
TdWPm4M4pUhgprlU0cOXDBoqyaRfI/wCo8kwDrWaiRMJty9mmatSSCewjkkl3hlH
eVbH4u5tswiZ9abesRHXmjnnbvDk5NA46RV7N+rXyliPLU6r0e5+nUNtN1tw2rlH
hC24Oc6tR3fU3nIu554hE7OKEP/1/dPIOF8lck5nTqzbG5N6A9nIxBN3rE6YbVNP
D5kO9Zd2s695g+at/BTMt2EDrjh+w+Arerwxc+939K8xalH99y4Mb4mAZcbRlgIl
zewtdU6DVvFwpcAFfD++LJXybgWHbCdYMqcj4Tm+BTNdF20Mtmm1EM4ZUn1maGbV
PT0EvX1GkLXK3peTG6FJBTF4e4vpi+Jcyn/Plr5Ea8aAs67ct9AiMmlvScJyx3cj
KR4VXcIkdiI9wvwUx7JLYl/ERk9MmCEK60iUbt2XP4Pj7DVjwvCM/AGEOwkLrOqk
HR+rZEFLrpL3GmoGe88g1KjPA2jU7ljyzJMd99CxFtDSrOOB7oScCbL5EwbKS4H/
tiAU3S2gv+uFYf5lyYBYHrCQZrgDJgVur8bqOopL1hPeImTM5MFseic5bKFl8TWN
nitB6XkqhwgSyeqahFgEOUcp15QqdSgkjcHh5pbzhoUgKUbN6UXvNqf3IgSf5OeB
aeh5xJiEjHCvhiKzLVCz+li020RLVneBN5q0SrjUfG2kgfZLjsi0vko86T+hjHzN
nM1f9FUmj5zoXV1YtDQG/yJ1dO4RrS5PL8/8kMQubRQRaC2PmglabtP1Zyt2PSrk
hMKb3WmLHFDtcn0iarZKhBdDFsQULjMuDZLwa9gyC3/xaXr2FaMwmkqkSe7pWWZG
mQaD+AtHmeuO99CDset1qWYneP/0ELC4KZm/ekGIwDseJa8nyFiNysJVw6dI7jdx
PFwmh6xNGU9r3OoCd095P8IAjgBiBR4iSYCv09Jqe+wm5BaHSzN/Ua0SkKq7E1ml
S+3ZTo1vKVIaGrGLdVd9GwAS/mupcXFXyOA2szZqXmuZL/PonmSVEpChV5YEaFLb
+TOSLeXWZxwFJu8TrbMZT7jXyrSMkxL62awuevu+hb4iBdoH1xieWBxo3jJyRjA4
Zp5kGR3scobI+CoWNL7gpkKcsdklNCTG6tp2XiR+PPBnabcfFzGE7A5XL6hB6z6J
GC8PIoYy1SSaS3uSV7HllNyxp4fwUl6bC54yw4a/mgM8OcBPqn5Lupr1oMCSMZbo
f2AQvAdj7lPbQuKw7/djuS3t+WjenzmqwLxhRip6lHscSFJjsNv1TBEvnDlmqAL5
/sG2Tt3gOUymcUgI1PFZtjWZmR7tTltrYP4M8V0NrtEzGcaSDEI8tCFvUbnNvGtb
/JHkpovntvr6d4JE8D5oIIqfvjkuPXGTJUxzzgOLwtkQn465Tw+W0TW/gxctjqr5
wd1jnIz1pFsIhUJc9EHMOev/3bkIWMDe59oJld4CzRLsmeQOHn3EXPxa5/HBLVYg
kDEegwz04s0zfS/PP4MizF9Xy67sWuxHz1CDdgCG4EIITrEKezy2PVvQNk8bJfJN
hxClZd6xVJA5IvIt0+1Zu2AJwaEwWW/X1vDs5sMa4gNH+VrNVSumbG8oTU7L/QWJ
L1WroF7qAGS5g4sn73hTO5BNZ6iYCzchKqBFSAboGLhh3W+yBhsg17W6yZmejVry
rtn52ju5ksCwHpcmTb6v711ST3nguT8NqNKEfI8IE7p/8ZlqLb5qudMq0PLOdS3p
MCAcVpSceoO3ETrxPJedPh62eKDb2s+LYXJKss3CgOZ9X+s2iSHo4bLcymbZACX8
A3ZVK4AOKhKfEE13y7cC3TdLtR3BLryKNSVcb1OyEs/YoZGd+N2BjgqgTNyH8Wbj
VpiKm+HYIzgoEpsbFHWeTLTx/LkI58NFYj6basliiJX+GTC/iBL2BQ/5xqoqBrIv
EJQ8SuZmhiGThcdyP5jds/G1VHozEQMXjALNT8DGQbGmPTnlgH8A/ZGK+K6m1n8a
u/GtpfosyqdI8IWS2SalMYFg/8BQw0B9PSV9+YbdqgKfcMiRRMeF2yXZabFnwAaa
a+PCGfhQj5lXOUwn1TbPb+gb8HBp0/OIDGOU7Mu4rmt7+1hdVoxpbsnkdX9TWSsF
Cspsxt5FM3QGVtF9ijlxn9T+ZDnXVmgZ66dmUfU5y3rAeqkS5ny96AUV0SI30bcJ
eW1DDOa7+Z8sGkBbMMKDifFmKLTEri71U96HYfXqOtb8yt3Rl6Kmjn4Sf35yGAtQ
Mx6Lc5kxTeNSGmBrg2L+7gqklCYJnjt8Waob4ECXUve63x1V/ZynMO/1sM5IUbGt
bxuE/CknHZzRM0errYtnzcQZA3K1cIWnJK/G4Xxgj8ZeCzFYC2OeiYe4M5iXDa0O
WXTfjzmvCkCeXIftN3o8LKsOvvHLN8468uiEcwie5f9c8nV7CrkE+gvJblf1Mg25
kctAKoBB2l9NXVeHawrCvzFwKwbXlc2e6hdqvDhSz6iyg5Y/Kjp6wxohHQryHWRQ
Ot5qp3vCSXa1v4cvLISQc08cX/6N9yxlyjfrw7Hys1bVOLTFEMUMD4TbWUnw2sCI
Z2kk3BclaxTymA3Edli/jd5ZGBxJKI/h5Vq1tbBIktxM/0pRBT7Ro+jBPipn64Zu
DBbDzvy0p76F7fNd52m1Tu7+ohgH14vK7RgjkqsL3gx28DIV69+TnsdWPanqiGU9
JZQVuvGCGGxkuhLQUfDJHCeCJxFc1pMZx7lK/MlTQEyohSWpnrl28kpmwYaMG4SL
SSr4mKOLIHtpZMUkTh2D4P4r0HWTsBJxOXSCsgxSKrSO3lGjGho6UbJmEG7dmxMT
PQB1HaPYYJJVBvnpbEfNTFA6l/sNJskGOQZJ0YoE0TLMIy5chxnJTDCQcaRnchzo
hzEHgoIZjK4qwsDWXz5QEkarM0eUqK0Aj9kqOpwGVfUQ5mw3OG1mXyP20mWsOqVp
ERHR98ZeqkGUgPfwnab4MBWRxlJAwE0VtJNABlZpZpdWB5A3Tp9C8kSNitgbKFHO
axBu+FX5r1X2R0SXkGPMEanXOTZIHZVMLXY1btAExUEzy88dSV1Li6PnxwNO7ggZ
FPTEI6gzXaI07FVdHyCsAch/WYbZMUKVV9kU4a4ezz1HcVvAQZ2/uqeJ/jyvRwtl
1to7sounuqT1ielelqjXlMMrJuxYh+4psagevh8w4X07KysmOSf2C4EMu5TO1WFP
tGKTIp+F4LsCyR5OnbKmHmRXCYaMv29L+/kvsqa+w1i9cC0A5VGo4ZkeAIRUJJ+7
1Q6TLqWTlqAfRMZVtGV/IE8kOLkguJdjop3rcvD4iKRPNxexFu0ilkj9firbwFek
q6vFzDnu71PiXUsmPrJd2VV4HKjKYsrOQ/euLZylYXsB/a51UwedXX8SQ6X3tmEd
vgYkCQZzep1r2i4o7bwu/jQNR7pcC4E9DYHcK9QUeJR1lHCmc7WT7jdk0X7RiIuz
Xz/Vw7V9/p6DXAqMdfYs72Ub6a8+9I8UUR7qrGrWBU6TgpyOKIoE3cOYpQitgAfs
Ybki2SmAkR1per6DCXUiIw9zVzL6reZAVIopGkJP4B51oyJL+FnmLysi1uOMsMEK
82Atj+b65qpFzsWMw3WLJHpJ0u6ky3Evaen+yZu+pa6MOF1MEeLBFnpdj3cKMjz8
md4QnE5MYnWSJdNdKPbdAPxw/Ivg0sOuue5W2l1JiYekuxQFkuFf9QHb2cm03mHk
NMyODbabJjv/AHnp5Jz7hcOvG4Tu5LFOskJ18nGc4z7slJzqx/2DpsNGJAZP+Lfl
UsWHjORm9iH4C85tlRCL/lOeu2wWX9h9T0rUNlppXZ3UvDP0Us6sNnXMoW4Dh5kp
ag0mLfkbAHI3xf5ebDRKd6okUePlJTaAzSaXSXLbF2L3A/9xtasEL21qvAq4vm0Y
KAXQnQ3+rMtsehxfdGdvNHxBEAvEs2OvuCTp4eZEXSzyADFhstqTWs9m05p1nrCX
e/vV2knWhbSXcEGJkwC8DtW4UcspxOn4KNR2I+P7Otwo/7pkKTSI1fjPRGdhnzhJ
NAPQwPZjRS3rAJcJxYAOSc/kushYqmoSAxD3nQceTE6ScSbG4Ar0fBh8KS38EFfG
foYZkCNFZ6Y5/9ifqRezlKXx+G8cTrTpKkYGrVVJD3XyKtbETGO2Eko/xFX+KB6Y
GisFSSfUftSJwSj+UtX7sF3ahmUsCqj4iUKnRLZvx4RPCsV6afdOPm1Gsnh8TiOL
te05VgNVI3gdAiDupEjk7XSWnwHRtxcMesQoW4clijPHFPadnCkjUZx7r77HHgVF
r8N1zyQmgsfQPTEOSvs/hfm+DLRTGyLCLA6pxRBsAitfR2LecYWKHFJGty+pH6eN
7Ov2XVdfEo8m3ftRGURd89D+3kUNnznCHaSM3YIuClyQCJM4MHc5jLDrzTwPZHzb
Dfqfvyl4K8R2RyFbvE4NwK21DfXKz46Rohia1MPW8BhA+Lz2rqX35JwdOyYwUSgQ
mZJ1Ql0FV2wSWgkb5g60jsBKPEqLmvN7MpQy0ogYQYmWYCnNIhjY7oayGn6W2zxg
ayfjd7JxhL8IALnJbIC0Skbt3DvuO2NsHmcxt4E05tFkev5J04vCDJTanJRjzynY
L5MHninQlBvmN0trRRzSqoMAjty3CD3Z6HyFwjmhg5bl4kEx0YHkY7yP3gsed9Jy
RkRRTb9EGZpRqirJkEnjGByZ7I+D4LP6dHKyzJsfhP+r2A79830zZJYhW57BSbxt
LUruHwsRc0Xic1SkcYXBtW32s+XwGnVXQ1JKmD7QlE9gMQQCUXzcGO1HLkPXFeQ6
G1aOXudowa8L187kTRU0amkBgP1q9UT38aZB8jO6PNYynPDC0F2abWCf6iR2iQcp
Jp6uAPaDtY1p/QwZ4in26JUmF9UeO62I645mYEc47BZCude0nlf2kLS4E7/QNZn2
UJMZj8n8d0AjWYigmIj05iwuH3Rs5f3EYWINDZaM5W0353jRHRaGn6D+bQ6uHfaE
SDNSdW7PNIa+qq6WldFZTeDMu/9ASMYuVhBQ7aFZbUgU4CyiEg329Ox8wCmQ0N2z
lWBvqIPARa5Ugqrby9cCsVe2dwTLFkSTY2cJUcTDKqatpkz+nREjMwDl8dgFBu2X
n+weOwqXX5OqO1pC51ZQcunzmnOT9dU+Y3JbzouIHq9d9La4FxIYYt0VFkWy6iYF
d75EQeep8eYv9KcZlQLJNMP3F43VjeRX7Ppzg8wHweqGBTGTYl6AVLJ8bdf01p84
D5jnE9QBEtiHhAcBSO5azNTrnSmXE61dl5tGqkJkcIgFubE+D4TYHmWO8AVEyeZk
lBwiOD+4WmIAm7LESwnwssYy1uvMlRp6vobFFXSTkp4RGqom1eNJtVczgrFCQsLQ
yWiHmqSdWm/5ehmPPl2kWdJYXzg3g1v3GiJQKosySuex4ENp9KAt3VZIRIJrJOqL
02xpUANVEe/ldfL23y5/jPmbHBLuYqVcm06I1poeUkHwyGO7musgFc9/QD9tCy78
PSu+TeQHPTSmNfwdT7SDvZBiD5a2fJjL73Q+ons4k5liMpn3Zj1gb6X+ilS5TDgC
JQ+cK/PWlsXxLR3S1UnJD+Nuil1j4y0LldgU9KmcnyWzZ9Clq/FSLeitwqL1NJqE
JZVj4Yl4vbW5YHSBByt9cguCVeegqh9nebzbLqlSbOLZhpueVIC5FV1tnBZQbvft
/QFC2fLpFfzwb8e6FzB5VBuNTluTCXXUj8LQCLsiuKAraF4XVk3ELVUbhbqiupMR
OEh2/Cq0ltGvi5N0VbO8HYMCFttcsuZayAe7ObR5uwSScuB8651kVG3a48ZsvEdC
xyKqp1J74XCpco5pin1HPLlvtxANTlPphM9pisG7NCsdhR6D1rb02F2+V8AE+6Ek
xxaRra472M7kciQF4117qzYJEEtCXGk5WvQV1QWr5RFZypHDhZGUFUxj1MaYgisl
blRYT9sadSEvTHxAy0JWWeMoGY4r9/Bq6JR7ImSesFN7qivyf2TrvhyHmBx/UmQ2
+6p1p06jVgRK3bprpwoZ1a6VWHJ75hukkv++LyDzCMfYNDePNxSZtc1Ac/nvgWkE
Ic6IVRbrHrSl3BBaDW/9nme3+eU8a6zDaixZvG57ndTcoaTsXghKLueujawom6cC
nL8hF66zaMWZ7fVbAXMa5RXudn8Vrq/DtHx1O101I5M2dKu1IAtfqWypyJodaitt
FRkYSh1W66b0fGCediO+mAy4PdkN28zKAvAFHhjrj6tPLnDeoBbf1qdnG5mfqTZM
yxVEAa5ktfoebWpXT5yI3GDUDTsnN9eRU/cmhEajGdHYUXQ8nUP9jo45S7nyeQOk
6waa8md8NgKjOouvwB/yoy1zzpJM1Wr5xjgwxUCZMHsMBWycBFiHZ6KXeUwf4sH7
hl9R8gsWmHA5ZaYHLZiNA7nDcODx+KrYbR9I8+VX4fRZbdgVxFjS+toRn/gdS0pk
0OcOmpywCQq75VOuEviww2ue7g2/s7LjbXQyeAk4zoZ4UySmSGZt3XDaFo7MWsfa
gOcGAq5mWMa579Wi2TrMOJqUOrpm7ylVHIl4Fl81u2HwK7Gq4FqYE49CVs9DKLhj
LZiq+eUTtHF0CjF/qkxg2mFHk/7nYw5q3BI8FiqHSL9GHOAyXV/wSk/dCFPyLCjO
IkDKQQKuAeU2ucAh9D/G1UZaRiIpz8GrzvPBHD9j6zKmJRiKHVYxbtAY4MQXTfnd
M1XgsCN1fRGjbUS/3fKpaXFejCcCPJbIwb1i3FN2C71X4mh/vhG3nzMRSms92Ea0
CvKB3qLpcki9W7pSKo7Fyx/RVeSZ0qVGQ/hJptBc7DEFfhMylLAJhykRuXMpgBm2
z3Ge6luqs7OuRRd/oGU+NoLaEqT1UutfHmnvhkNDpO4nP7BjfdoxvaGDsHzT3Xp4
0ZY/ccbJczLq4RIEapjNrrRk2kVxUsc9GEd3FcvhDIOnXnUpDQ38xzIHnwFYF0+2
zkJZC7JJEVODdxbkKe7DPok/upBfDQ7kK3qhCLGpc7oHstvXCly+CNDI1xz7Zm50
/CQuNCW4PnqeqwKS6EcaXgOHGKeROjNX5jeueosf+R3M9IHcqVaPcylhp2kgQMfV
7yX7uFpUiD3DcAZJYTQtcJIRZW8+iR/MF7IRXJBAxJbHEFyZMfGnEgzGN1ET0HJS
WmRwWO2wkG3HkHCgbNajDBDbql9Ime4w6nBEOaf6KlM4yQ6oIpWRHq01rko9xmWQ
c2tnOATTSS8obe4g2wXiZ3morRzikzlw2WckiXdWSudG3tnKTSwmuD/WAiBGaKvF
6ahnXXESaiwJJSUGEqTFddykTEiTdnBNrXvW8BE79tmVyUP6f8GVADQjhfhg21x+
kEFL21/Sy3FUZ1H77b+keuS5uR0C8JpEnWgkxygmyWfpVWSd3Zj0Wo9TytjE09EV
mOOVk6H8tF2G3IIaLFDZG4B+mevUizFl48unrF03u7lIccqEvQ21ao1Sci+RwiLz
pFQg7+D6+0O+7YyTMSO1AtNVVa4jao7YEszDpXPTZN2d3vbR27reriAyCLnDtF6O
ONiTZZO2robZGzGs1j2BLnnHEM0ptLkRQJM+NzKsjwa51muWDPqaBfxzuHN6iKw9
ayQjZwj5ovJQmEnAZIhWnWOPXljbxLJ624VKxKphWFvaJiHx4B9yU5+/agt+jxuj
dXLT/WcMwCMFUB98MNwsE54FFdBKF4qTr/FtWIbMtXjPzryVRZb9SqGtGKtZE3+L
ywAfXNwoWNTz5R2I8msxLvb7GHH2T4lTvTUU9u4dmeUrY0nRoBiEQFrEthYukpi3
Yyny32W+P25ODJeeUWY+biveEHa6kxvBwxpU6r6b9mh5RXvO5Y6+jWcXc0AtuJdc
SNIMWEM6Ufvbgeo3zqRVU7nml/vYj5xb1tvl/60D5QoKzRxYqICB7WHxeJwcTPkG
iUsQSG4yhoUbVwOof2XaxqFQy6yWLLNydgrMp37LZ16VWMJfBBYVqu2a1HFWzsXk
fWoi4+mRBopULV8rOkwr8+TCs3y4N6xCDEqVCO3PhKAWqSkhMLS6Axovm8WMMPw7
Aq1s+IeyJEosVGWqY9K2HSB6Erg/TsGI3g/AlwEy+c691od+3X4kMl1m+0LvE9yx
DgsV7POHvZMZOGZo1ih6QEcD1QRATLOV2FRyK5DBAyJyfMVm1D8nyGEofwXn7d08
oURwNoIfgtrlpOClUYsQdfMkzKVJ8mBhd1CPeQyU75juN4lUAE06Lo+g+muFxZ0a
b2Sy/+XW6k3mC3xhhDqyXuOPaTXI/CNvkANuFAzj4T00UN/9wJE/MgdsIyv/wgP8
yYCGQpPR4u9ViKDAUQ4jgiZPgmZjwwsdEAZoI5Q5koZwmpKNT4Wvst2KFnpYDClm
PBDzMjWf8GLL4PuHUhYNBJYbzirtFN9t2lb2Dnhok9zJjDtrnVDf45m11kOd2mCc
RDmbz6Qs4LZ2e/wjstR6FtZruYyAG+AqbUO8DnkDOUmm3Xz1bWkHUd4CC0GERIz1
MY4ojyFW1FgWvVktVGjQYOBx7OFYI+zWIGyX5STR1p7erWF80Pw8EpAq7k0C9zh7
p9CbJm5oFVGKxCalJLaNXprudvY46La38/jtQV1patN/t30yQ+7p2HtNoCR+Z8zG
y5F7C4+t6dQ7UCNDCOzAk5IMb8U9za2Ut/saljUd/ZaaxbHcMQ5N1rGrfCICF32h
Bw6qn5KMZ4Di3qk7sPrq8E6D52m7pNKz58uJxd8CqBHlEHQ1T6Dkf3za58+l/6yY
ipUNxD4wnzHyd5LtC/7i7JeLRTHkXXJKu1DTyv68psSxT6yBpZItc9afVPaC+yHE
KE8oFL67xP6wlI8bojZZaKtTme3s8o+C7qVoWc20JbxQlspOJ7S6W7rmVH+Npuuk
ENIRQ00jkKHXnVWEaH1gB7q37vJaUB3CRvQvMN76uTGRrsqfvoSC6Z2t10EeByEj
stIXr8NMSqFsqMPtbZxa9ujsGIYJOig0HtmHtcMr5cmr3OPp+7keurtfJiNGWPtr
QuUGU2PuLf9dcEUpkMtT8qHwsYP/3zRkM16YLJEbJSJbjtTRTuzxAoHDOW/csCOZ
NFK0idC5bQYwwO3D8qdBjEexo5btLrrw0dSOk/Cp4NcTdwdFUYHzo5m1mkXMCh1E
tRX2Vdf+OXikFwZyILMWY0Al42+OUHwqKt57VUwc//qQLaTju0OkaCCZ1++2BZFX
0xJWeD1ZHlCL5noMjudtd0SzFQvRXhkD8vkzhorPeTnp51EnQrA3m9TNgCDpb2j8
uaeJGNGlQ1IK0dLdUYCFQPnuMQDcOBepc6fcTt6kbNJu+hm4X+7MxMqc04u6k77k
YdKOCO73Mj6mXgKN8rRjz6krs1P2FE8PKrcPcvlky9ZX5mxpA2P24vcS8CmStord
kyjuYFgel465qGA33j1NCfPE8IUEQ53nRidAbltAIN1ccdo2P1ENPOs4Wni+IhmO
stLl2rDHMOMBOgFMmZC9cT0p7zW9u4nMa+sWEYNlpVJcI3NfkWi2b9C3syd2J2uV
w2hbuM5AFtK2Ozt3OhsWdmpP6Bl3pVgdbPErzrkBBabqxrU82xyUvA3cmy1pEybs
GUC6uMWXlrfPGbkmJWAGSRkEcFyVmULMkkl0gRwYCC04cgWJms16RPWwtQ7drq4+
+CyRcwNf+hoEx3LlrmkkjvJZz/G7Mlv9Qxc+Bxxuo7IBZe4jeJ8B8IRre4k9lHi/
xmuzRLDmOS0MBLs+jthptK7EHkuzaBeMEZRHrgZ/VYSCJjzdCn7ZzalwKcIIkH0L
68w2RwoeOgxz27TDdkUSzB5utezY4OKz45RVYTY/uIJI7I8Fc5AJuJWzmQXtgBAn
oAPb0qcSB/d9U4vzDtufEMeR5zfUBPBiVNT3CVRHfHk64u3+gygjJvpZylnYsMK7
vFWk+LYqDkkZoAYyHXas2PSuFBlPAH9wUtkvZeZ4hoUiDVN39o+Q5l/aQRCboo4V
2Z3pXWj2KT98m9qom8jcZa43C04yDdN8VWjK2aXRinWoYbxtDljVp1FdDFWc0lZg
XjyoSrSNFInnuL48wR2v+4UTZPwFcPHf5VTzMPnY59tKJF79x1Cu6JCC6359zh4E
xK7JEkE/ikZBJJxhOyxW8i3wjpW2cDV/bf0l4G7feUCOLhhc9YVPBAxlh21DDHLl
fb/00SVemY1DJLNO8ioJ0VR+GxZybcxwhOmWayQr4j1L/TXvC46Utz0NIk3yHDSe
445mKA37db9gBmpYoxwwDS8iPvKRZX5q3mMj920vBoVvUUxadDZKNkILYPSfuUzu
yX8GwTQu9LWQb7HQnXd/zdMkTiwQBLNe8/rtDOkKVJksCVsUpF8oexT9pj1RmkmO
vyj5t/53t1TJelMmfUE5bFOPmvggpk9A85C7Eq0tZ4ex4C8NrVlc62h4JBOdQahF
wpWLqh4SON8OYgXyprJSfhTnlVexFlatpbKm6jAwB9ADjc76CK3vxDqsX3worvsf
qNlHx5NdNh7rZxPopwEG+JoDYegHwMLfrdPW9ELlUN4LUO5j6ajSHJ/3rac68JCA
thuwlljmlq875vSYof3tE7G5DASf/MVER3nnsl+nkbHsW4msFUgWixEJJeRRSZlu
Q60CLE+mbO8VN0oTGzSSbCEkr2m7c1SXLdM1anGKBS6QdfmIUjwx3nDKz2hL8gr0
7nFWw9yZOLFGAb92XaZ/inizsztk5G314xIdiaM2qd2D/jdw3JeGgMDMVE0OZXZF
CPvA3Jo5RTrppnwBj5QMhEgew2kW/fNUWpV0lBweM9S9pFANDPl3Pr6U8WJoD/Fn
wFQQPF/4EbyPPh4Yt4At2sYXYBvApm5BtCr5KZQSCEs731W4RaWgcWT9AKVfLcLF
bkkEA8tKYNXeku/wqDQxRftgmlQaccylAMC9VKUvWjFAl3mw1OUElYFN+6dYXbc4
GEX3rU5t5p/9IpobOkgaMPOvcWXxM/5eWYeT9qDPUNNeTclGOEshawmH7syG7nCh
xmTWLBWbj1Hbvt60HaFglXzGAD5Alw1K8xfpcStp9FCByxRC/7VeWO4zi2eJknsO
/ge4zl0LZSHiZzcz1KhbQMC6X9b82sJE73O+WY1uAKPs2pFF+suu+sV+nIUvanUU
CG2Ty5YQT4XdNjiZ1h2uAVqwl+AN7Y+9oGoZvToxgK5i/q9QEtqDnGsV3FXC7NO+
C/CnR0ySnDgAMdwCNcGhiwkpa3I36aQezociEiaHw9kc3GqikAR5gWxlbJ67jNDP
zkLJCim/ck1GKBBKqN5eXZMzF3qOhzxEYnwwD9O3sb3Xc0DS2ZNfMfGKAHztB3zC
QdVg5fDCzMqZDD3ftU5ggjmR2WrXzG+TI1P+/haHXSg/1aCYXhpk/leNSlmwCGW+
aCR+37j1bUgQuWZ6TBrkVEfWPE6W60a1bAwGaqenrh9nvvFn08UnCL5Cij4obe1H
ZwNIm2SFGlG0VBLdKYLrbFTRDrPdb1FmvxoH0Uca5/pYdl8S1bo/FcBcwzr4Zumj
p4vY65k+NDbIuukAL/NiVxPD4AwyUK1mjtUqSwfQE7XfxshY3uysfeofvPY9cXjC
YXjJOi9FKQM0RzvTwy8ICL/U9l5Vq7sWMj7WEIBnHvwoUQ/zyoFR/ZtFK2RCOZom
1avRgKiXuXOOf0AI2Svj8oFhwpX0Dk1HuSyMj1pZkQvjS8W9BqWxCdQkR72q8Ms5
uQMXUNg0ekzmzJgAVU3Go4SDaUSbbd2WmeJkLGDpLzksG0hPRYq8tHZvGqC2VApP
z5HhuvOep1soNtgXno4KCbh90/DABzZ66D5a7kBc/VEwymbwE8SOww4T9Dw7jO3s
zQVPIjVGrDD5z62uyqE/TCgze8Od0wyed5g1e+jQhmWeCPIxhxwPYELx4jWf5NDP
oTwqrP9fpLTSZoFG7FCRvpKXnrpb581iZ4pxRMAuPlxZK622G/tPdyILoP66Lb4u
gEbUwYnN44Kyt/aciCvymjqx/f55tC0WxPlSh8mruJE9UBXHCUu6majD3yloRHY+
opgf3CpUMLmUrwifGx/W9Cl/8PQWNGHasfs73DqIYPhJQG2SFozhvAUxOov/3YQT
CIW7eQFZMQo5y3erKErnUBtSGpGzObHKqchoT5/PAtWG8mSzP56plErotJV2MJgW
6sRrrmTRCnCZDlELLGeQTuDZyEl09WMVAmc/YC2wZ3f/412Qbz7Z/yb78EGNcNyC
bS2RkTUsbqsgM2DbgQcVoH/3h/VbNoeu8Vh0l3BoOG9/nktdzJerW3VQAzD4mHoq
CivucbORSIGOw8dGWX0qfmMntl++GVbZxUybuNoJtoVYnvbCpaGS2egdZPe8hcgN
eWOCGmY5YT9UW9o1rSTLMKQuCFn9n8lK/p/tuswcSJ+PYoXkB9vpKssJgoTwgkms
D6G/qTwGrIkdrDl4xGVIfTX62Rw0dvp29xeglO8nvm0q28PxXbC5v+hsoG1U4EQY
zSE5WV5COh8Ul+iEsh3tvD88hee3JJqPHzDmX/isF5nkK/lrHK81eRJa1KSJ8tcr
xqnjic/W8c5RdH6vQ9op2bb04YKiu+UVFBIWU/Ugx64Agwbgq+MEpBLSEXG5cn5o
SE3O8vO381wUjQ665YVVNxtgTttcEM+5d8KsYGGIyvWcg/sOtZpB8LGUjCD4JRYY
LQbb2fObgU0iXTonafpbbS6WjxqCFyG6hEGdL4Nz4lPXD3s/vrenmzNabm10IcNN
jf7D6K2um1mFvQ4HEqCzIh+Fbqh27qLowupQ1wvnmc6zt5CGObVxkYTkru1gT03S
NJ8Nt15byI52mGZASC8A5rznWypDtlP0MBHyk8DgJUQ72MIHvHGFkzjqAHbWjTLC
+H72NIXkPp1yBqLx0smPgrv06In4sn4+h22x3sG2HRs0xSxee1yWLIHHh7yl+kki
iVvTxFDOAh2D5Xfklw09YfjsvIyOYKLK6pLKvMsY3Nq94j5YcohplUSG9lWd7+ga
qoFNMT1ZHMyZqS48AX6ty97gUaIIba2cnTau8ob3xgZx5H5QqBkA2CtONnJV/Gfj
KnJfmaCpzMLQUtvvDzr7LfN5hW8/GTxQIVm9lmUAV8zmwfJbYLsNz9kU938Cj479
ENkEv3b4MzztdOs52ZthRpAYUhZSzej9qliH3J+88bA1vUlVBoU+17Ow3iVAcyH4
9cHFtZmAiKrqnVxV9bNHMUu/frSP5A8j9+QYPX7qvIb5V13xVFTooEIFWb0CTOMi
KEn90xSUeUtvE3iUIfFDkl8UPgSFHoc+vm49fHd/qmY4j72bNGPH/sE4qpL6Vraj
ybwuDxTfsyZBaRUPUuXomocMuk938rTwiyvODLaEEDN7mW4LTij4/gGRDu53LImd
WoixTfrilVF/msgzz2PM1zJ2+X2k9eDMmt+7OYoXwLuSi1ICKBYHbJ5+SE5Dum55
vF9zk5G+RCfp73h4iFYfUuVDWYz42+nZQbmJHYFFQOXakVSp8J5LxEGH913GFhTg
ArV0EpY3tX4pbFby+f45v1fMVwbncQtjfW6fwUoJT8eG51JnI4tIYQ9Iut0Dpohu
W81KvVilCTJ4CATnKjdYWJ1HI59yk5j6A5XyU6aQQFlVCsDPboemdASrurZRSBB3
joltOtlpMf4ekLG6flmmc/Wc0zo90GxzWjBI5gI/vVSFvYn7L4uS83RySLAY+Vd2
V9EfY/RzC7WtkkrrlNZGsDK+6yvS443KbMSdUOZgje2l4DFMXG7u0DEes1MbHqfb
r/uzkdXOB9ov9jakwNjlGE5hBcnNd1gs6pxZOjpnoMra48/jsDaY36UaS299qP+O
P/RirQylCMjucv1Lt3Ehz24PXDRZOtRTZ6L5QwbfhEvdLV9rk/e6Q0PXb1+bFBGd
3jmXFxo02SqHC7wcF93uPaFatsvlB++blRe7bux60FfEtBOA8+8en/5/I9qmbIWA
mysD5vEdlcyRT4sR6wh+t4/oGIF+7ZFMoJ8WmXAtpYwJd/+sg3F2DRISPYrTDmbn
IVVCu0nMU8HCjhZb/m/9ARc6GtOjM/KCzVyG7MwW1RG/+d5iRvZKDLhz7/q9Cxli
DSGqVf63JXZzEioOcyrJ07rqSw0KBYkcbzYNK7bj6n2a1+Ucq2RssaThw3+e6WHi
sIyv2CdRCg5jM57bNlhB9979z+Mq/XnUYMs6YimvJIuqPVhcriems6p4Z1hdcIaI
ePWsM4gwRC1pdorPQPPtZbPg6VwhL1AxPBbsL9oT4Tv3Qs9gwxUFLLjkwx4EiBtX
Vl4gwG/WzBm3aoBWVYKjT3yS2nw28BXJ53+W/NhUmjijLRTMwVEAQ7yAMZhnYwyL
MVBojILdM9HlI2qVeUHLR8o0QmdptenS95FetfMlQiCPubPRN2daCNrL3BQ5C3tE
ce1u+79zXMO4fl57rQOWhT8o4BqJdHI59xQZj2sW/uKH1ay4/q9HhFuvA0bh9GLL
fNv0CyqfQn8Rh0hAgyfMG3nkSsIF1yhE64AzOd2cu7l9dq6pU3pHBfjrKVzjU6yy
lHdFS1gE4vmmdSU31AsoSbaBVad+jrsbSaa+OaUYUqaG3GDE2b8nuhfaWMEvOT4y
dOCvDBqOvlBEiHJVld195ccfys3Ianm0eDIFA++0H02/bmBd5qlDvq/mXng/shio
u/MyBOv5UGMpGVprInqHynIuQ6KjPaQaatxBR46MgvtSty3oCxvutW2BcaqcH31t
P8Z8s6BjtvrFm+moN6BtvUF89UFjLwWc+Jc7G1YsfGr49TI6y+mxNcwnjVUzt9Q9
g7PlOJSXT6sOfbvES6BBhGskwCcfm7Ra7kj8NExF3y4qNAOwAIsTRsCy6c7JQ1WA
5g6/BjwkdeKnlgnKijhbYXgqWqsb7l7TvDU9XhVj21pBPTESGoAXvEYD85oeipgS
yJL5peAr/YYOwrrQMmH7IqqPMlAEUT5hGm1/L6nXzZVsc4bbVHJI2CMBlcbNOTt9
3G2SMpSta04QE3lb4T4wsMOUXD6bQRMVWnR9AL34AIvyiLERBMcfbCw2HQAnvIbe
ytzcFpMM7sfRSyAmcBxs6zpHHS4UeCT8gUf5shIy/9k8kFBwSA3qnJVqydaw5Vi2
4cBYQe7OI8snebpRxQufTAbmts+fr2fWkTEniMfW0URSqGylVBpkLvxaCZjtrshe
eDiI8Wzp6p/MClFw9BY7lRCBJh9vtGUevH8yEicMUOzWSRSKkrvbwiQVydydasM1
khLyMqpIvmdMwqhwftHKJjigxwzR75kyzNQYc/1IdRohZ+TtyPZJHMs5bSrCkIga
mBrFXSyx6Gw2xNw4iYdTVtfvXmPNLbd6uUcDp8scGzuDHNHt0HIyi4Dwr2xJ5W2X
8V42OFxSB6ngWCZCIk492t2VNa77Tlt4s6hK3C+zpOdU27d/CpvcT0nC744VZQoE
VzVl0x0jyZuJ/pbktGYGl4BVmRvQ9RvQ6hHnEZS18hgX0WHCWNmFY62LaUF+2Oze
slewfuTl/WS5T8ensa7RefY+BIT5Z86v+jFMo1TgrBN7tBHp4nKfCFAGjVcFlCtN
CQhSbqCif7SQuWa6OyUeCxBcEo7zkdXV6xyfhb9ZDJyQhBcidL9DGFedToZ4bmBZ
d+QjeBZbym1fFfczXn6GbKo8FFzCq4oP2qU3z5LbM7841yVSE4KXQcK31BBRhguI
SmgCkqailVbeHshupdEy4w5tjwu2wfmd1jPEg08weMIjfqgQ2U5ACnRgflbuWWsk
WcVrHQdoTEZZ8RFQ0pNZ9aoNKzg5C2dRLxR6CWC6xu6nvS1mXB1D+/ruR+X/7c/q
dqy+wLowsnU1L8pMpkHHHHQkXGcqrm/wAnCnuJWbRhsduZYCjDRDnFbRBCC7ykGJ
uPKtXy20UdHfbidYBZSUMj7C8yuK05Wkd3yC7Hn3rhJqKbumnUoks3RNPYY5yeEw
wJ970DjbWpD9J7tpZS8eH3ZMtrUjBAxtBwdPJNZn+5I1fk6HdlDs2nSfpj7qj4lO
U8P0jK5gZCakJsPTfVjZ+efph14oYJjgu/oHX/ZxRmDhHq9y3f+zSOeAiCGOsre1
ITJNVHeUpuqtAJ2U8gAmmuZS0ngToKPVme7pRqvzShvkLMmQcJSArwZxyfae5/zM
nywup29JgaoJi0uPJfd/8/ye80xzzAYDzrvTMaV16/zaHLyKIFf95vc4O/l7hbNp
xZ1GRn2lpf//4Kz2W8mktMxPiQyCEr2vMPaxp92FznXLNK+4AYm2XfM93OwEMbyy
GVFJ9sDuaJQW+JLCT+0Ny9TWkYi701/UzqvSXv7dRPKiMNRgrROna0u61G069cEE
H7vWQG4dPyJ7HyzsnxprL4jWsrzHdpm+Zk5EwDRi7XT5qwKcABtkzelUMBj1yWL9
PUCqxBGK30rgLUV1V1m4pFn5l4CYHF8RibfB5Bs8Ht3OLs9zFk25kMfRaJEBHBLi
oGhIKuxbGb5uest46nzHvXmEPjBTJNlGv368LjVvQv3EWadKBlJ5whBUbz8IMRwR
keIUpLVtpoX+DuXTKWbxYo1dChO41/zzGA/oqoLFgPql4UsnFprGnJJU/O5l44jY
uJQgG5bIizKiINQsImn3WklkxTjGo3Hli8NToG/ES+GNWzKk05A2wduo4BVw02WB
sY8wEUyJGUuezCh72IGeAgxAaiJ1ukiwccq6eQOyniSZj0cK3HUZw65JYL4QUV66
g5DQNr3F1cLeHBE0F/R/+8D0x/wkujjGFPIKwBl7+j8U6d27EG3mqi6bugd63gXZ
+P1/SzsjTpqZRDnvmZzFz8L5XeSwGenCHtegzIIfdgsjorLRoGf9cUxlT7GGVePK
w2RPCzLB6MEcgAKivrtGbML9zeywihVejZJXgopX8JgGw1289n0C8g4A2zHm6+pI
moeMG6v9sE46230AlJ0dOTi1ibk0xFeiZ/0eEGgsyM4Bh2OFmctegGwyIw9sel+c
nKuThudWJ0MfYgNmW177YkQKbqaDkjz5OZHpZa7MgpGVhWUSGY7Wqa/+YObYcHts
iozJg+E3IOJRR6UVed/cuHgz5eiwYswFP+D3ta9fP/AAb67C8Jh1o/BHxVRIr6lG
sJJV7pKQW226qeGwleAsd3A7fB/DFcKp0bRHNRnuZzW6bxTnwaT/nJdrxNSKHxN3
9W1IGEj6iFTYYstYwELcYrnh/TQpO40Ph6zfKCTUyrSnyeDZi4j4ddZ7tQyTTQHx
X1o64k7Zq08kieBGZ5h3R8DwAE5C4FXojBspNl0LGFuHBoO3Ed4tQnOgOWgKsv2c
rO0M2O2buN9KN2h8vDGbnHS005nZjqKqn6NdoYrrvglqbPQItAWjaST9IU2JKw24
5AmF3N3VTUltD5AnaI93uoXxMQEYdudK9mh6TQs2LkK6dZGvJQS2T05/sgwU9yCn
AZdwMSPlC+yg2s66/mBN/4B0q78IwEZvLHfbMct2UW0qPRNss6W1HuhKvFYC77XU
q/jSPab/KFK2LG+uMPZTv4Hj+MZIsTRMAd+OFmrpaOqvmDiIMNzhd2lXNa659l70
bxJ18CcwVrydzFue3PgO0OaQ7jATglQmxFxF9SVlq8zdomyFYI8elcTB1c3VEZRJ
OaQ5N3ujEbx1aMmJNX9nu7dbXMhbJYSBBTGK+hCdivbyqjOz0BNHO+swJuyAMZhu
3oFkyHOLoGEPDItBY3Y7wrSpW0KxrWGojh8Rp/Z758G6hBrwEusBS7FXpC0sPRer
Z+Ix6HE2lDb8n3k79WG8ZzFGOAZVclLTEKmqqqp+zFkU7VZEVDezKJ/xP93EwhG8
TJVv1gFLnoCOb4gkG6mW8L3OdrLHAfyyMZIGgypqA0D3JqqTG9Gf0bVQWpeWsBCj
brBkvhSNfxj/l99gtNMDunrv2ec+KW7RbR6jwvjZjwtt/R+6NpoBPBF9cwDC/IdD
v1IlL8jfJVDGXxymg2yFOCH/n6cD79CONVrDazivoq2xQaMNNXXR4HkOTgK3vHb5
PA5SZhJlkZx4pvA0pba/tjWaLoeUDo6oBfqQGQ+0VhwG6UG79aTWKBSKEmFuR7s5
0GTaTYeuN/DcrWeb+tWGNfwdhDrBCQx6iUUAviDxHS9gu0+9CES5r8uIIbZRWC4s
1cGyi3rRXt9wopL+xkh6rep4/cSbe72y4qNFJH7C50I4jxoGYy5g4PCMLakQ3lEa
CQnxArIzTxsUbsLjP2HYMgoj3jWh67P06d3oWCAevu2ZieBDZV4F/9vVSiB4QarC
CQMDirCg6aASotC+GgDTqRpBQBwt+6WeG+Ljbi8HNd/UrMyY4DEJ55HubzTavhkr
8NDcpYGDW08lmOEsV7i4R+lfgPGBj71EOpR7QJHo0LO6SSp3353dW03kOb7e0RpV
kNQehXlXhakABlYfZTf3a7AH0bkU4aBYANuejEwHsPUg3rEH9su9l2c2bNmTJjfi
5iUipYelyHa2h2Ji1m7GQC+zrwi1NHK+xGxKHaLAN6IQc5nkSBis0JrAkK1Z2foK
PRtMEugaB6DLUhaDS83Crtw9ao4aXGYqoDuzsI4w+BGT0IeDUT2Jh22b4uO87K0C
3nk9xTLQp2tsujf8kqZ2ubgJh1p6UwM4gpkhJsXm26VNU7vJTalMifTO/S0GE2AJ
h7gVJHYw6hfJDKsZXcIsdXGFPx3bu9AIKprBCBJr0aSOdBGUA8xnAGK1jQUUGypE
LMPTR+6aN988sdI6ubRjJjZ6TkhgD3NyHCwGYNR6mb5DdVKyUkrDxE+20GZnah0M
KtA6qMSWWwAyQztT9YftdRVXxeXpEtGX/LDGc4QD7rqZ0RLfCAArmMR1IHaEdMTl
hUCHjW9sKbiopKqEzroor7mleyo4PzJKyZ8v2BPSRlIF4aZq5saYqF+3n1UyBbA7
UpGLkm4k/z68qUpw9JbGknvTlAMsDCSPEnocSe772oqoVPNZ2yQOfCpC9Ymq/dLQ
TAeBIhZrtOwROqfJK8blS/tyBOrOlX2zvxhcuucXUkWsXrZQIWOnkLZkneOo27Iw
TBmzliQ3g+SBfy4W2AKMhtvpV/dBxgow4uNELE7lMj3+8S2CyeOidF7trilJfQt7
0ATiFxJ+5VVkDFNd1QUHEahZeobgPPtCgJ99e2/vqI/WLIZXwmODDdaq3J/vyQoJ
6YBQWYwsErms0mCy6W7hwJ+k3lpbew1ES6lBVttxWCgt8iqKRKU8dL6Sge3LGHoU
t1VTinYmjS07FmJQGGFptgrNhHb7gysGObk3LdgqacMYZL/1X3MmHL4eUn5Y0MQ1
UuXugmhkLfc6O2SigM7208uFQPwk4w68c4A+sqF8spf0s2WCqzfy+sZCpEMhHtNv
fdgwiI+j6wl2EyZ8nu0uIKvQrCNmCcHUVU+LHVGIORQsfWAPX25DpKs9omUTVXMd
HJGa9+fl5gfwx/hgPwI8eHTm/yqsS/s9kHJwIV698bHDyjZc9GmeDe+MUwmx3wRw
WKXM/1ldhOskfE63xGGYH2UWbjAKr1brTNUPasQW92G0FKTfpIXi5C9QATa/d9+a
atcckiFydSafuGHInmRGtTO/xJ+VrMVquArnwoZ2SebAOMniywB2f8ED/22VE7O0
jTczDt58pu2rhulcbzcdob18sXzvIHBTlQ64VY0rhg1QijdEiA+7XdWsXtu+KX8i
j+t9cbYJmSql2Ah8vNGmX67zTfgHYSO8lQ4YdFsH8KFg5Y+8jEaZH3Lv8/rOUhyJ
1BRuIkduLRCfvDbMZ8zQoLUtojTtKwBQ8fNXv2a5+5F01c/OsVFrudH4CIqLnVHU
W1hPgKT45egtWOB6Snf7QcxXg4BmE3RXlYy0M48dIdNOb01Xv05pr0/IxUA06YKb
9GCt+WwUanLxDJF4z//HDvbMTgKGZji2kNC/ARpw6Uml2x1BgQJK/Mwyx5t/mGhR
zzP3lD7XcsK6ReE9/7VSfygi6RT6qXpW7S+Mj4p0Y4PPZja++uhCubnruj4wQV6T
vqR8WEhyipDzVxAwhAIZIJ/BpVqBer5mCZqWm2kpn3F8MX5wIiiZmk7xf1hOjEkf
3295hEEpPaZdRV3yyYV1Hv5IjcB9+nmgJeY+mBaZuPtOP5ymi4if3YZMzNM7fEoP
fVYYHe84xxky17+XIz3f89GDIf0A1y1pNyL4UxSgaLlGjhmqiNHcFldwjP6TCpR6
n6LaaMu/d3ArKI16SMPxoN/67EYOlFXCr/aHSJXXgNA3MwVbN+F/y0MIIXvqtUJo
hIXxInLX3Lc/cKfud7+qgny5zxUSivyMMekcgDpgUqDiIOk9xIFMrfnLsAuzh9vs
9vCO00A2n6kyO8HnMQKFMKfEPhDiW9D+JwLoKxEA6bp3Dk38oW0EIlx9anCv+Hsy
/FOQCD8x31IeSkzCtxzelPFhYzH37/cjkhOWYL4DpZZnSPpxVND2rxRQ/2oU6sLO
gtMYMT/UhBNyHSaKnlT+GOwTKCgQg0GtYaOOCSfSJlci5V6bNA36yofseLgn08YB
pLUPXfbEa2ZzTmfp9LJCxyE/tgc3XU7pJ8GK5vIFF1+2g5RkQ/kAXJdcpknIZCju
3Yoqqj2hM1GltX73SoQIzCAFH2I8iXzFXSikXLikLCN1Xu7mlC72O3DFuLzCdZ7q
aXNhsuAALyGrW90qC5Z46qMHWHW42RSsoTYcdE0OSNvXWIZikAceh+v2uADJ1wNe
PLeV3hzCummQPeiPvXlh+XqxMNU/6UqajRpPIhdqrcDKXgyLvEWutk/5LfQQpdJN
9oqwm/BNVdLzcZjhHLTVJTdF+hz9wGmKM5/PF9ZU/OPpfFNBn7NwK8/YQbCoHW02
Zwa5NVyThsZgeQfCalH+pfvVvZ3i0AG3pNr4p5rIMrnVQRmMV6jedRqipYrKCBlf
XBLQafd2Mmew+RzP0qm94lyuW1ohKNWOcaQ1uBic1DRdXAeSUTOMMvV6WuHXNzfh
nOHW1Zt56cQsA6X0ZdhJl/Xvu0cnm2wpMnjwodBP6jajS5qf8ICHF6QgxixAEC3B
ftuP3xC8bJ3RT7gA4Yt86ODZFCKNZNY/AWGWkGrRz74CCSiNXU438QWIDpSInmS2
Q6CxTwGemksCh7lFEakBpCs8wonFg0KkTMfv2jXbCn+cE65dpGilmwkHj1YSwxzp
M6/Tb+3+Yy0FNAnVoj7UDjjHCJCt5K0CQKEXfYcYGyIAT/jWAFIOfOIpAhktluyA
LqyHzeO3f+NvuY628jQOVVx085EtDny8YavpCRZpwCOo8XtWKT67vDb0SnSfipsE
sU2mW1Uq+1Ah6bLWTBht4kXoDwSRpvFiKF3DNLTOJ7dtlwB0enO/UxFjTeCl8gZP
fMXXIck9TiMIUS8VZHKIzwH+6P0IuNGstonUbE6emxOazKrsd2u6KfEQshgWVLGx
L75y+FQfxNXveqgE1kbV0Jx2QvYi4RK5QzqK2CFjM+qo7LuKowPugghgl5NGbGyJ
hnCLMAPMAnDU6o1CUsK7+MZI2K1R6cJOi5OHzvh1WX93GUTkRPgreAv583ie+bGt
IuA3IiqF0T2DSNle6UYMHNklN/JAtXOpEvYbAn3IA5MHefyZGxQ/jXbDfvphWR6y
v3R0de84rYUKy8l20BSwQYJUFbyi+nNNi6TVLgYWzC2wFVpvUGumbw6UgwmJl2Vr
2wssKBhVAisBkEbpXsFH2MfiESJuUzpA4hnxUoz0aS6tM6vzS8FLxPK1Bgxxv0OF
IsalsfDIMbEFBgcQYx+QFDpIkPUcsZSHePduy8WgtAHg+8MK7PkVyB7ikm7qT0Cv
7LpyQJFSukEXa/9N7ClOE0JlFtPcmYWU/WASUODYUJEkzK0hVTPnNMJHZUapBfBq
PfghU5AoQ9MIhUXrSl2KsvVrLD1O9UzuwZCoDU5f4vd2r3BjxxRJiidGkz0QOBHc
E0PzCORf8CWSuEDZODE19fudJVe+0EmQ+qzXbZUDUsvzLxgQEYdN1Fzzskdoaxje
LXiRCBRnD8dYOtVdfmlRKCrwIJaRXiWnk7kV5mSLWL71UA8/dXztf5LiFRkMz6cr
BwCHyCx01fXkTAH3qq8mWeF7fOq28Wy/AOf59Q/Jj+ez6Fn8I2qID+hS4s42UCCa
Hj9G/1k+UfYCWQqsEpPrTnUOHsqapwnfmhdOPJc3Q8dYMzCCms2/TMSXCVjDx5Z5
acemjF9AzOn+H07O2lYxVKPuTZSO2O6WlESO1N484WioZCmr9Elnps9cLm7xH5vO
43qmeodw/8Z7bCma0ZjIjXG3qGoE9sMmI3NSX8Ghsfkksv+slfuif9M3F/N0rI+s
4HRh54cfAV6WHbYUAqT5fpT35qG2gxL/kQeWCHFFqzVZBQroLkZiwlhzvisgLORq
nMN7XXZtV0VkJwpi5OocWQXDb2u6OCMr9miM0h2Rfc+8WzTPpS49pF5HbYxsFhFo
ZxemCd9hLXBFam7T05Qpiozm7gT2o0Q9nx58tPY4aNmyfS8L1Tb+8/EffC2BsBmd
rUpzTYkgdXl3xIW/8b55GLVOxnKGHlIFua9VHC/LVhwV5zNXryUQNjl/UdlgTqBW
OKP5TGgt0EzdiJdx+w0AxpQ2z2XqzRtJbfhBOwqdk5g6wp5C0mvIfxbsmOZTS3QN
Ifm00DpKNCHO5MU27h23CezkoJKZLRGV9qbddQ3k8qOdN0LL8bB3LrYITac6M581
Qw5rR/TILcuCVJgDBfgMK37/bu9Wgf2CoVwG9Sx1Stbd5TyuiReSNfWWhPyGiE9o
4PJXiUHEDypL2E8J6sD0Am46DDmy7E5aPnOAUCm85xD9owhBQXooZWobbp5w4wBv
qJuydWEZb/f9RB9AaXEFogPUTQhdsV1O70aHstC3SoeQ7InEn1kMUoB5fmX9rRLS
vWn8ZrHpWWMuA4xYLbVYn0GIak1MYBuUY5YLToB63A33xRp6+yFZHuCLRBnO8tD4
LTnSMkCC3CjaNtr2j5PlqdV+UW4phwefqoU4B9skB2pdh7lxVPHpjTtpVAzE3S6i
ZlK3kv/AUHfc5EBR8z+lECnDbiUImfzS7ioCoLSnfSGw/FLOzwG9NtfQK4iwMK5r
ld7JWhu+dK61QsQgnLqOtL0zANHyJ6ILiOknJJFNWNR88dK4RVDLm8vO5YC7aXde
X8y6okcg/2guVGA5msPVjpvua704MagLgzFlMi/bOxfWfujHFH30yB6VynkKjK7L
hXLwvBdJ8otZLcS5ZWo6bmjkNoA+slv18cGTfSVNg0ARmCEahxdccefc5azOOw/O
N8ooj5FD1ECnNYqD9eToDla7INIyX6cD7mmi9T+cA5VUwC53xCG8YX5kdy1HFCgb
Nph4/wCpYjcawphqRMnChqGKxglHeops7n6AjPhe3zipVQETFUf38i0yaEPsUzpN
HdB1nVh0LvuZC8T2i5J26PToUUKEPIodlMuTxjKo+IW2wATKH2bRFinq7AJgAwAY
o40tEL5MhuV2oDEieyMPkkyUy9FGnJuRhvIR51FNDJRvbv49sVSjygQqZsJ16ZNQ
KiSf2K+UfHrs1mSRXlVSGDdeK4t/ibFxt1VqL8ETjYpP9sqF9G990HRPu0SGpyr0
ipf4WkcJtCqabt+umCyKWWvpeLlry5MtgkO+9b/W9IbpqhgsY834wtP3yVcOoyjl
Q9Iq+3xlJwSmqmFUSqloAYEBWmfR7ZEAHWGHnn6kW/UvRIqqql8a8zCVZJz6psaT
jrGRvwcQcJXSgpoG28wp21JwP7xqwFnlfhOQpoMaRyHt8leQdZGcD8L371HKoHrI
yIHr73l5beTlsoHIp3YBnFizv/LH7Ircc30P2AiQWdFVzGbCn20zHVzvvb7aUPyh
OZBmQT+7aiREI920uzukRU/ihEbM10BzfkpGBOfNjP/YgCy0rRSfJXkppxKWKSkR
UW4Me1xRtL24Ij5BV/KdKcWHIG2Sv8+uJhRcCJ5UVzatc16/Z70J4ngn2AS2wZVM
jDhkX8la3aSwV6hQiJnyA/T1voKTgIf+6XlcBossN/NVmN98JqrWJn+n2aEr/hzT
3e/WeSpPrb/GTBAjVBlvpeCaW9CBEaJrSkYZRYoDbWYnT2+gStyDDIrAvVpWWL8H
7zNCt3+hw2e0P4MLyMbj0BGIVyyRhdA6MnvVf54OFF71bItr6ae74h/u5xW3cukc
8MD5aUbNsBimlsJhbDf+22wzaoinxayQsreD+NY9djJhSkBpGOb83ckYJx1hRBjJ
Ok7gMS6gCNwhtnxmh/wdImuRuUDi0AOG822xGrrjqbFqEdp455ovvhsZh1fj7wNo
P3Ma6CtE4S7f2YPEd/MSlp3ecbDmOpN7Br0tGEQXok5BOah8d2NP528uWfqOIja/
+/wkYZszOV74ne0OicoIKYXAW34Qmt/W2CL2llCyQISABxLOeAICsxts1flt5Or6
cofQXAyfHt36m9gs4okuztE06ykk7sR2B5cYbNg5lPiVxmbLsJCe424N86HTKNF2
9WCtln8z8ldd2BON9rLguhtMInrH9dl+0uSUP5nCMDoewMlIJvAxltM7HCAk1wFj
7s6pnemb8rpH7bnbtdnnQ9RYMYEcIivLWpf5BHBMfnGbdJ5/NeXpQSxiRJGOcagn
YRcnCDXX3MjQ0XbTOiMor2IhL6acRfuvweLshBsg5HCrHCB7KWHPz18rGoNQS/mQ
N84YvtAsIEC901UfnHEtz4asvNj49HkuVHS5g++OKrMYrrPV8/uKE3vH4EhqhByo
FqDtg3RUjWuWECAKo/y0wj6rfvovC6Uo60UBJSH+7JeZmivxLmz8i06o8K2uEJVm
7fwEghtk65BaEnJGrNrzImDNLBt+3sA6ikQCsULyzUeW2xpn+GsiMxLGNhvxQwru
HpsiVPTAJFH/63xdLGWQ7VMCM+O9KvfVv4X/mtG/WkLo8pXtx9JmiIfRcM7Psv+a
z6Zty7Do2OW0MMwPCsTG4ReE+VXFF84hOlnLsLUmOMLeWVQSYaR1LTfoslGYsImG
tu9u+x374wNHL3lT4TwOqLxuOrc0Bo1O/udSu4BcqECxbt3Jjteg/TLrpAoUkaet
r63ZY44MSb/Q2qDQiwgBS4DljBK4Wi0E6tO1W4AvKttJkanjNhH4N4JqUH0L2QeO
h2A16pfhb+r46Hv3xHsStgk7fH3IWhPLEf+sqD5IvQyQEdf7aPrIaqK6wxjoX2+1
IxZW8gwfOAGanBiVulzU4yddfSepMWGx7grnSCNrmzL1YDE1gTWaCdhe4PFllf7u
ehv17AZv5/7JoXsRYDoZpQ/eUn6omH/enfaMgmBbuoQRjoDyj8WiLs2dBn7xBieV
0PcSQT79m0h6MU48hFWLy19ulS3REVsTciBoxKYbKGiuFPpvDd45W27MZ3SVY4WH
YbhC9jrOO7mRuWs7ik3zPLOmKSax5O3Tm22HosOrT4rxkJv/K+oKT5Cf/VKkhW8j
VEwkOAZwgEppxNLVXX5NszptLvGETupJ+/bKZj3dfSA7ihJdgmUljZpcBbJ3lKqt
5+UTwzL4yaXgI7HIJoa1DAtCs1NPhS//Hf1qZ16j4vHmtiKSneB1MMYqXTnEQlWE
2JXLm+o4QZapzTg94tc6jvDnymLNvfbeFf31+n16wQ/z9QIdYG7ZugixS83nDkqi
20YiQpVueL90Bja1TlAm94wd1SyUet1EfMFL39FAtaPhl03uh/zSpoY/lOnGlAau
u54aqHxzFZQWmStdo6IlApgF07tr1QMkZ9mBQR2eczMj1Jy3RkTj4QT2pfW8qpc8
07ZiGKLaFx2axLh1qOFR2ZTf/V/LQ4fDCgtH8ba+eY0+xVtN9Su2xBX0bZ+3Hg22
VyMAH7NwxiJbPRGEKRb15VKUT9e3u9QdYrAXGq/XYJnn03WmgPPJwgUnoR1g6MoO
lJxgMGbGLPvWWsZ2TM6PoTlJ4ZUhogvaPuiCQTYzHejyYWfshBVpgdQOa6AlZJzk
M9JPi941swkLXDDM0U2EcMiPDEVMZj13UM2jeItS2m1rD53yGn8BiQB9kKf3Ovyj
guNnYAXqZcd77B6rO/L4hAKKTg912OT39yXavjqM475U9G3sK9IL8QzJYXeQYqzI
VTCNQf5wL4oLS1EdUXt1R7qR3LLL3UazI1m4jWDwBsVtpeATvKv7zBi4xe8LGVAM
DKPXqT0GSpd3GToNDWYNlg0g6xyWHT5UHs52Ztk3B8AfBfnKyaZMUNqa/1/fJd1Y
+Q3gk8m9KwWNckyxJo+S/ZP+XPB/+bGmw+LTydHU9aH1E6Z9AT3lD75wOE8tIFrU
PldxNQHbg7drzYnUurL87uHj7ch5cBVfF3snOuFg4U5ZgYs5qAwBUMM/SZAaEMju
pzwsHAeMFauyxFi3XTB9g1EkrQgopAh2PLeqj4JAmR26VbZk2CJFGvCkY8FFqNcj
6QVfS5LtkrQ/eULVer9Y+YrtYpvLOrx+E5Yds0Kl+K1tADQ+FL62Ga5XrTpUQ3l4
ke34n4CclvSdteVKx5rqK+AWZj8Nn42NFrLo28m0Yxu33qHtuEk/lfPjH68xVTvI
Ff32QFacIjstaH4JW8hvy+j1TD+hEDklqbO5v+agRkMmSUGTlEyn6lF/lfe08V1r
78AzxSdgyaSJ/65lT0V2YbiSpbuPI+fpG5uspr2b9diTnf+MRpvJA8U6s6tgWxEf
69QtJO7H4JWOqQuYTNEpQKZFG/XQLsYwyg47+OZFe0PYtIxNeytak/FG2IyYlulF
UyADQMl+jPaN+ApVZ3pH+/PO0Vg1dLmI5zmOcBjzFl49iXXyyp8N4mPiEAYJIYOU
XKOzk6cNhyX5yYhhDw5Py8HVigA6LGw3JkPypQTPtKM89LZ4gex77dhAFVGVAXN5
XxNrwu3kgi6td6qyv+zCWk0N9EWfLKYs0hsqH/MAsGF/nmM8Tqu3Ytw8N7HJ36aJ
kTpS0s5NBOkXMjIC3M64hYBTv0Jc0O+9qCJmaETeeFokTqF0x/NuU6QsvDZu0r8M
6mZGczB+muLdLPGkM+TFVQn8wva5SMTyrz+QhDt/Wh6RhT4KU+2AIUcsUsCsTPEN
QX5vKtnxaR5itk/dkx2cCC2Hho2eHcWR/I24B8sWAk4o+2Qv4zpSDBBmWiyu/q1V
kmM7jhHm+cQ/CHXjOhRc5XG0uxstLZnVq/oSjFmn/32d4dLDbLFqX9AOJqSKtsZX
XzJyIX6UKsYufPk0z0UXvsjWXD2SdXI54IQo79LVvzCdKljvFSOqddcEBKt0gvm3
bngenMTBcvoAXlZ3JdJBVSkDH5b70Ec8LHMcU4ec89cyG50+w+Y1No+FVm4MMai/
wnnENOMaIIEnjTaGtIovb8BtJ/6JlG12jNYSwCsNaewiAH/7NwX7VT5NHMExpJy+
PIZw2omnnQFwWDEflBAneUmcWDjPGZZGZ//27Pz9bSN8W2la8+uTSnlSzu6d+YRK
rq1StCJG9/mCfPhiKxtOoUYQWkFF5tykOoBUsU5EeAdxR/RXc/RDvxObHPXcg635
Rtn7Tzi7bD6i2SsLZO1BqU8v8oegJCL4aA495z1VqJ5Je6spUZQp6dGuKQ1GXT0v
Xj97li5WlCBfbW909BtVc+kXC9poeI5ecQwkZwcw9Rl3aaitlo8JvIJpp07blErG
OMLpKpng0HHZ0RKpb9DzFLvveiWzZp9hLn1Rn83ITItDoE3rwgG43+aJxGDWZuBG
phf3WpmaYE3FrL2mWGYaX+WIAdkXjB5+KzVJD/8/isKXOuLV+AtvFey02dPbkyff
Xi/J1x7SeEjH14XScWMTjY552r7YeZqah5hnDGzJk1T2vOHGrRv9g+Z++y3F1HwZ
E9RpFs/v2WEodjlPK0p/+uTmbrMCcH5NAOfZzvT6U8S/8I+76TtUb6RS+58tnjg6
v2Vt20O3yizP69OoACo6/6/ncVf335WUBSmPmUfmh97M77BDbjEoZn9J0UYbXNYY
xKmye9Ts9VzmuSmgCgNfKxJ0TpmllZ6CzLOuJf3oz6R2BvBLKy1lB+/NFoCO04Kt
xeFIZ0nj1l5mFB71KltoEqvtJwemkJBu6yWmEC5NDXDz4CJL2VyWaCY0O9edUcUP
ozyhDsyA43bFM6XAqGdtVN3lT4KnDTewabjmkuJp107jgN3yWivJLb5ICP9Ss5qn
oFUbHbPuWM/GzvcIsvLvKnewSLUadv+UAnr7xaRsRFnHbfiLgFe6nPQBqI61kXqN
cRWciY1Q2jp8B7bGMT4QwJub8Cmqu3/XwYx7vLbhvNYOg7l02xvFV7vIYvPRD3LL
9x8o+eBonbNaP9zxg6CGFaOcN6Ys5hyhmzbWhNNDhEOt4gZtyKjS2JGmNYlNcMAq
oZt44Jv3GMGuBo2KeLdNxsh+FqO9XF+61xCx0hX00tJro7BRzLdCKgze2dqUAOxj
RhkDS5nzpsgI14Xm+YonkscLo813RwzvOY9ib7jgJSgOGBBNdBjVvArJu1tRPxsD
07bXbdK89GTbZuXcus4xuMM3CRXJUIxDOBJyLdO1hvE0c/UQGy72soMyeTbzo6Za
vOZkhZDqMDaE31B/tzkvooyorqHYz39CZXVDogtd7OtDMCbJOT5JIaV3njvIWifU
XYK4SLwU8gQIg3adrbphvMAqZReyNilWgImDJ2kSofYxeIg7pVIkabPHJoxyMTh5
j7P4GEjktnN1Td+ydDCh2jBcrTHNVA85jTrKWA16EI4td65W4bEjtdJG18L1AtNd
BaaNhy0n/YqTicr0iTtV1R9mERxjg9JI1QbqLG+whZPH+aRgI/jaLFZgHpDkunLc
agrI6ORqvmvWa8QrgFjgW1v2URgjczfxDT6JhzzSB99EVGvYTTG3BWYw57u/i0yg
MQuej7AnE9GGi0K+GM0ecxqknGTWE5d+cwua2yVZKCFq/Mk+xRFfchE0fGVu6m11
gwRCPzaJvRD5fpkFLdz/4NWJbWPygeva5/6O/SHoSh4SQG5h/DQSy5zeZuHWM6by
La/z2oEEirbzLDyMzl7uLWI+AKWFKyHfKCVc7aJTlTDF/hLBzN0L2TxgFMTo9rKz
b7wjFc5vDohCfMHsP8ZQBfIOH66lS+cFZWIt3EZZUyirLKzWOXcYlrD/5bZZA0BE
bc3dpBdDnmLkbRfMyzy85UjoR1OYdOyhX9FHTceLa5Sr/0q2tT1PWujWNonJWwUl
ieWdTmjZq2fr4VyqQLp/+ICkPEkHBsodGpyaffAol97uidEADEGs+Odv8V3ij55k
BhfipO9svNLo1j1fPfFt6b7oV7wc0eJYW2fUzgf4iexOut2FEzAN+jB0vKagdfuB
DBSxnAKPhes1y4fFUTJBA0j6wvyxpAbCV102+ROdk+b/o9KPGbejPqJjwNtJyNBo
YqmgsfXGxH3beJsI20UxXQc6yun1iEW+cxTFXZ2QK/L7W8ZrAzWTei7iBFirrOOl
oc5by6ujop471JkOaxKIRCf74NkNtrFphgOfFvn6kNRIuIy/TruEpX5mBLg//dkr
JCphJzhf/7PnBvRIJYrmhIczrcA7UytWV4y2got450AWek4mgdMFbDYCwEtbgOS0
0ECQxszpQAaOsnSrvpr0MYoGaOsZ2FZSNq78ZSlw8zxTnkzodKqOowdI599z8zxS
rjxtGAFjsg+sy7LfzdvSArywoQst2nGG6lpneWydUaYv13DLVs4k8nldAsxYfjpk
WceOHhK1hWLiumKBr4UF769aOO3Ggx46Fjl8CrDCifvrEwMQYxRGk91tZ9bNVQIV
YbAftpnC4eXrXB3CLczf3r7B/3jQKtyl+QzMTNLMtQMwAxDDar9UEA7uRSbLlcid
x5eTtSAu3sq9kryN+Nj5MuQKs5hFdKc50l0vSloJFtKyw7cscPf7iYS2kNP1aT6l
lgmeGbGgY5gypO4DFegX0sIHhHTueFSpPWMN3FMJ+YwXjgQsD2VtCJtMeJBn/qN/
md8oCumcyEOs6h1fBJIrQJjxQbRzUTCyeFiQ+WQzzmlSztuOo7aN7ybySSEZuWdq
+S0Qd1j2aem9M8g69nHHMtw8qq4k7nnDYDfNmztyoYm9fu0v5gPLutvl3++MFqiI
TViFaSMgG/2b9XlfRJdlm4JlDmdsmbSLNGIByBPlRMlJF7MFNSmJybAuGpBHG49y
NjmkxKCPlTckbydRPJXVhAPHtzmhtZ/056wBijXWl4Bu1wG6gxQyzIQhsMlUVnZ7
xzuHJAy0go8iD70fad2Sinh5pjFGkUU2xHxjTHRRS7gHeKle+Rf9TX6XqatK6Zbz
sLa/5F+vviRz4nYI9EJ4qAxOxcIPbwbomvlyoTDxzi8Utb7td+QpP/wYURP1/LA9
5GZAh0fyNvr7GZwOmIVkj0WIJEoglxgBmfFG6zz112d2ZR/MSRo+HSvULC3vZXpL
bGGmGl46iNhdYHxI0bZNoU+r6eAxay2AawLGrl/79EPtXSZXSOU0HXitgy54OVPv
6OgQw0gDDcE2uV/Iv9Y5Ij99743mUoT0ux0aZ/7WcGrwr7DANw5oICrLOXFvoUKx
Y3t3k5zh3znmJuKoBnF7B1gG6cethP2TImFqmSRFigzSnJsR8iQd236eRLQNXLDe
/b8qWRBG6eUA8LSrTUVKTue/39LgVhVQCyX+8WwNZkZzDKi226btXgfZUkKoJH+W
mGcbMaGWEIJbB6nP1iYqFJV/l5nBiLgpWzZ3WRlJ4sBKTHKmaj3CaJ2s5krMu63b
6xuzsM6wMT1nQjLAmD00DelydlfkGi6ogWb8bJP4C5qDMq8XYgGy5P2KZh7HGzMN
LRnQNRLg+HV63rIowsf3v+1HJ35LMnaErRCBnB520I5QKIdHmcUPy4Rm5HBROW+D
Qv/vxK82Vx1FvOq6NZsEdGQe7RA2CXWzentKYPzwbAbpnNHqj/13CiMkNVgDu0ev
Q2Jd41iAbU9vZ+IJWQ152ya+4NlnLQkg2z4G0+jRsFZDyUwt+WNdCq0DEnJKcwju
k8K0WFek1ofwX+D78V+KCKkp2NQgiEKB055b3NiMGoYVjiabQuVc3V4yiQyJVrkf
Nr3vQmJhzi+9ui/8Jp0iX1KX23me5dykGxJYxXuBPj5fV9wA+rQ/qjbo7HmNj0fG
DOrFRCV3mfSM3NETB/HDlSuiRAjWlur+/sGx6AEHBpoqU+tmQTPUzB053Llsu+IJ
B6i1GxBn2Jqa2VGaXDLJ87Gk5CuBzWcMlF8keNWOj62W7CqDtc0EbhgIsP+7lYF1
Ya2UpndAaP/8UavxH2ycRnFlxxLQJzXPPrYvpSdxBJsJeCR3q3RDtZPSS3keqG+v
lyDs/HUF8DzyExFGPJ0yYBvYedkwT6n7FXgUwDd+LDb0tw9PQD0LFEAeuaYamM7K
5XBSGxjbxB7rl+4XXwMFjiJpzYrPdNLAyvY9sOH10kPEAPAuuzYIeA6VQ/Z0togg
FF6QyrpJqt+9miM3kegCBSLPEGCt/WbNPKXWZD7wPLF+eJGoxWWnTeMIkKa4xaPP
wGDbHlTAiOqw8uoq4Yjyu/GsPRFPFKTDB46dcMqcunyDc280/rR/gE6YriyFyWFx
UQhAm+4aKH3CIHViZ3FC5xD+cTjuucjKnISYlEW68/WrRHSsOLUqw8CSpFV/mvLV
ccK26ipRdsGHDGKVUP3VAo50N5hZnPSMdOvDfIFC01L7n2XFHbz84m/FqUmMxz7V
1hpTo4g8JyTNfT4yMK7fhrxFSM2cmczPCamTreE4U8Au5grYmwqLWy4YN/CEpiOh
yg3wi1KCkdynD/MI+9rvOZgwNCt1h9S4aE0OT1dwbn/49xlhj7NbL2zSBg/c+kDn
EsQwCHL4YmClJ+PBnZr2jDn8FJlZ2NsMowuw0xFfGG0ZU3EoS+2WSnkY5rP6PtVO
afbOrxQXnkgxrCdmEVQQBgQM50GxzOKA0q5Dj7tgxV+8OXdgH9E3cmrs4o4+UA+g
nBDzdKNDkImsOH1OatgwrkiTiLMVX4sIeMgUBawExusZz3bbvuSQZNP+zzegho5X
OIfJT+d8UGOFMwVO7uKCMCaGos9n9a/h6vbW2l2KabiWDz152Mi67jNkCCc/h5ZN
kusguZiHQbo7AlS6R632SwvocpVixkm9zj34IP8tEua2wJcutAQt0p2dtjgUmcFr
Hw1zBIwVgx3AmFC12YNSNVrfjb2vMJiaRMj2qu4QIlLrJEsH/rkvcLpr/k6Xj3Jr
5Fa7/ZwdtiQvaWnUYDN4qpfoGfvOSqz4YCRNHfeeE/A2aLI0GpWAa/Zw22izw+iC
JBgqhgG28VDQLvpWPJ2dLPQ2bNu6tuA1Ygbjx22kOKjQWxafoiFZBebzktzfAKyM
am2RbzeLuZbUTy8Wywewxn/Dt5wtHm25jhnmlYlDmpbE9CDZL7G3gO4MmtXss1tb
MKiaSGxcsC+y+JTKZ+nvPVPztkwjz7uS4tH1+vnr2mErwvZ4gn3XiEmMCvFyw+vH
8BDFaV3MhvpJgaYgN0cknfavrwwQOpdGDD9jjGnfePi1kYwGC7Y8SlOh/8vxU+4x
4HsrlILxjzsp1KW7o3jjFWlutvNhpkvk84OPLTbWsweqoWZ+Dab4e3yMgOmyEZes
Pj+ynNFZZavWnIfW6guKAw/xiheZQYY8wU2dQqEOunpHCRXX0Z2gU9zv6lXUeHE+
DiaBtGQ70wThugbGJefSzGXU+z9V2DxYZt3aREM2ptelKV8cgoBRzQqgFZ+rslzw
TdfdOtzySlafcmuzy95fLjFqlFfoLigh+FGZKN3vlshpxKkBl/wXsEAuh8MmMLXk
j7ioAc+13XJCaBOYMOmwPiLJzqNNh+SAQhpcy97l5GwHbL9EEdw7Bhs+vsQgCcWC
EKuF8HuFQ7ZjfSuafRbBOhnOHOf1snIvuB9lPCXuIr4LOU44xZRQNwkD64sLJzIZ
1zWsaFxHWP5OB15PNBVG8cN2WNriWznI9vTDIGPRL08TfG1enUTND/SnjP1OWef7
xnSrZ+6j1bMJp6LH/EGdCWKhiMVOaIoqsTpiIfk+DXczS9dd/lRo9wY5VUlZ5Tw8
yMdu+PfOKMMD9ArWLqM33rRhgTCOFhPivZdp71xAwFrvqz8Lu1hm1IhC2hDQgwUE
g4jI2q7WpO5hsUCp3SFSUFHbMYVDFp/aTjseV/6Q6zX9Ei8qCk3sbOgkeAZr4W86
fJIV2TebhMEn/K2KDx0N6crXJe2TA8G5aPDIdgqK4o8JmFfc2ud8Om3bdoaA4H6V
Qvaf1nJyvjxfLfpQq5WIGBBakN99DROqnRtqgFhTtsCYRcGHZsxBFGgXMy5lMeVT
vnXyTewms0pVU/PyBka+kyAnNeFAuhc4m+TpEg9oznr7D1hhenJxiUOm8I7yOHH1
7WB79rwZgdyprYGXJAnaCGkPvDPk6XTqvSRyF3bS0hDtd/+g0Q0A5+ddzp9KqgWr
UogOXzGMFyfeHZGUzmQQAsNCFxYoH16ErDxFz7VE43wUsy+VZi8vi7rwCklqbuS9
rYQ8XB9bs97jpV3wpCmhLnAVVlEQ3TJezbIUVVtXq72CBfcW4zRqydmkLL78ZLl+
TB8Dv59evIhwyhwwXNglrbFWScQP9BqHtyztutwvLYF3W419M/7Vg6M5/XR040HN
ERNizB1kKrPzdY3K0kIt89/osEOsDgTJ29E9DlTWcY2DPQuTwSxw56X4GOOd3zJh
hSUn226PJWndICeiHoO3JcgGR0EuhYpREwV3XXzPxf3Cu+83Ub3u4LKHjA5TGkV3
hVE2cssDz5r+qjUVyfVKYhpx2f1YDJHz8LpjTVifYGGmqJvpqdGmR07BfxluXEjL
0itl4KnosNoEDo3JexlaQGKtZ2BQeb8fQ9+cBSTk72zqQFm0aYcR2ionyxJH/j94
9lbXg7u3vrkvJKbNBZr5+QzBJRY+H3+8IsKd1sjfLBd+XONV/BSWx9HOGxIxws+L
Bq/TBMFJ53DqBlmXGIyF9+J4KJbmPor3VCDZiW7V0ewYaQG2dSDlSE/Tq0BeXOiC
rM593zVLU7DUJojhmIIrgd/zWkxNHy27XUToLpr2i7hcQncZr6AES8Mf7e7n9CDm
S6jfL8nO8+4LamHjBNJZarNz7eCh8h8Qe8xuIQm3HWJ9SCIsRhImnbm13szoOa2T
jv4bmjcRcQQS/vq7xmBEec/HYvDcM1WQecarc8QJ0aham3nxSYvo0Lhuqw+KZ0nk
pSjoy1ZbuqAtC9sSCEfPViuUKautOujOhpFNrAxFkEeR0mw8rKza2qcbBtpVAqVJ
Nq6qsR147P+kFIbWp3PQLTMTA/tmiaIHQ7tRUEOChCLQ9M1j1iUTs72/Aa8pAUvj
s9mlxW/I9wOoQBE0+0ArDCoEyQ1mWQr2OfqB6o9eec7aDgVHWk062hZRojPxylAI
6Ke8qoFT+rwfJsdjCkoonhFzrFHCBQ0gEo08IdSAUFoZMuUgLUQmMuPDcZL6qqV2
EfsvA3DnOELXfaD5dCngtEChwLzLw/Ipu+qqLHy0LunslieafKGOrVR0YjV1DDvG
AhZ40+cG1KbeU8Tcd+1PXbbEXL9+eeP+JKjsaNqE8+D4XaCiNHbrrMdp82X+3zCg
mHMTqYznVZVFz3XCtAFJTUWdjkAhhaOr0kTKuHy7sSHeEfDKJ3nD49kTKNZ68p1h
//x7oQbijVCHzr+DqBqGmVu6jSGGUSbk7PPAGS+WQl5bMPbDUsKsyiR03PPU/wBO
aWaZc4o+w6sDoEpvsPrqPA30MMGPWj0j6PjBeooTFcoXuz5j0bXDn3kIzv/H1OLu
dUpNFF2o3yVu/MCpgG37OHNm0oU+gvbHqh7uIT3BPNviJO2aMgb1cNnf4dgNIGMv
1qyeuaULet8knhL7eZZZrrutY7g9ux5tNYkCjI5peG+x4xR2NR+ts25bxDCykps3
jPH8mlEUMoMUtGkDwGBaYxezGC1S7psnhpTCk/OhtKvxgYOsF88lLmk8S6juUAoc
DRLBJCR0e6PwmbChjxfQx13LrpvbLzGNAZjp6yCLy+aYbGJlcHcMbB0GCpLfI9Um
cR8FBstv7dgQ9Kr8yW4EIZQ+U/G80vb1FD9shA2xniKCq2PIgptuNBl52WDXaVoY
zzIqsXHAgNJM6k38UBe8g1hjW/7L1EE3CqAsnBd86wqSCCUzM4B1VmNq8t15ksEP
7pgTVmu7EaeVqWPmGZ2cMQ8Q4g1jc93lzXtNJs8o5e2xVbK1/eAhOP079Z4TRmKU
mEeeVF3dPqLMG9ABdF1743XNxgu+AiLkeH5Im1cKdo8TNxJymMsmmdt9IA6SZr75
2Ydli1p1OSluhbsILJ8JXq3aQateSLairIZiAqOkbL1G5SF2W4k3GJUW6GQtBny9
dB/oeGC3czXDwI7hOxvF0jhdKYmbNYlC0P4S9P/Qwsqe025p1VT2DH6bv5CxrTRj
SiLaUY8jyvfB8pPODzKZWVkJTfv0ik4k0OsFZkk1suogeDZdRdOe+tcg0nHeCmcf
4rpLCbnjmUxugxgqg9yMVU6J+bZVHRxIgaeBB1XhSn1lqrQsSjCaPe5JdJAx/Zvg
QgSd4Jvl9IrNWT86eBgM4QEgnMEWloensPmrEbqNoFsG6bgufXXXSWeTcAcLPAV2
3acyVMW/d0AqRgeruDkWYvYzgJQLwwMzYI2lkT3gK623y+FEcOvk7duWeaxZFD0H
MyU7Nu82P24S3J7MxRxPb/iA/E9Ism4zTHEejSY9kKWImRAZbIMBsamwAAVp7x0r
0YrIFGLcfRLl9zWu7SMVTNVAsuz0+ue65R/Jr5THEzsW4VAbHjo8jIdV5V9QgWSb
KVuL+81hRQlM3xyfElWZF2AZjd3Fha+po+lXGDV9i05QbcBGKV7+Wub3vkn44o2q
GH9TVOAyetohH1gGqAaauasRfJzmMvhPaqAkSPfn8U4BNKMcharyqAdEx8OgRr68
E5MWaw2VYFQro0PzZrADxqWOhsmFLBNuUhYaXdENB0zQvQpbqyKk1T8JDKVhxuzt
gNTNe2v/78dFjzQLFYfLahIAKwy/D310MgyNH+36f+uGL3LDHSyCVcamBs1YMEd6
m9klr7nmE41cIgSL88oBFW3RBNo1e5IpmLJdmrc2RoG1Nde0krVW6G4DVS2J1cQj
T6on3uvQFGkH+9lEkv0MknN8CPCxSvj4byMrApHB+mhawv5SbBLsQqoyejs8l1+v
bOVV3KoUSCVdzB16TZoN0xEgr3LH45xc8SH1viXP7aU1ZbIPAPZYKH/4qGLYgwyD
4OHxVk65z/9BlG99xJLaVndHrheCAdurh8qN4FEiTZ6+m415KwYI8Mc4jFjWZbi9
9UFit6xDyv1cbHX+XEQ+XYdks7DNtUHUokBdvKya2cyLXWuksvJX2aRhsu4EUVlA
KoCEDSelAm4RYlj1CqwtDQa3tezrB68fA6EB72dDao2te4gdqIbCqAF+Q34KKva2
UBr5hsyxbbvFYaOAt3w+hA7YRTEezb8bOIUBdhqfMkhvyklmswZWZY9RKfxw/8ei
PwDedpp5Rxddf4zMc1Cf5hJvaA6+ZUer7x3Y1EfnF+WqrXwflfp6/Bkj3NDUSeUz
ZnjJvxEvZMsJkX2z0K1ZIt4CQWQONG0MsQD0l3CxAYvf3A7zWz5zwNbElWH0N39U
OQjySG7c8q2h4I87M6j/Z0ch/48b1+P8yBT/J1/H3bYDfBttStQee8Lo7AE4E5Rz
cojZNC59xjdFG++l42vR9BsNW90ylA9AWGyMAZgqx5GvSmzN02ECymCmMXD+QeGf
mUfQAnLQzmMYPsKmx7SqBmSi//4q2Xf+gFdDtymSUqfKrMs+MaJWAM+wMKT1hO4q
pznvJ8gfEgZe22cjKNui1KJ4jJWnvIChr9FD7UqUI4TKmR3EPA2NMe2Y4/75dH/B
1W14Lhk198VwCsVKMz2HKP7Cr63mU0f9qegzLnxL5xfNIpwz/5rpqi0saJeVhN8X
P6RFEmrMC/z44ehhHVRTbZRHCI28uwtZXS7z5SSE2Xbm4eLGpHWA7XflQKiH1yoe
xHtaMsu4k2PDSRw1MdPNnRV1iCJrxkkR8OCCBt+ru4CCfzXtWcaUvJlpt7vZWOj4
Q9hHIDPlZiGfcHi6lMa78qBOCeUHWJtba9lbYqX3+xmP07mD718LwqPvnKqL90u8
1pcKKlBz/RqGuyhqaM/2W+Top0uAjpLwURoS+P3Djr7ik1/3WRwoG5ul2nfwjVye
lYdbScnp4PEUrjKHJqMZa+4SVcqvHxgEtLTDk3WSNef3gyR2FTfvoLkSGTAO2PXl
fzcbZy2uqcggP+BWNXdMa5M56I26eRy4zwsaJOZoSSNJQmp54/OR4mWcGlU6Nubc
9xZuW4dEjoOLG5H1k/YTO2+4PUi8OeO2efk7/czsE0Jv8kN9P0QFs0T8BWsAZCwo
bqgjcOSRD44DdfdeB696qavUhSa8vubmJ/ycaY6gL7wdIamKy1By+rafNmKVpgGY
OBvTkNPTUCgL+k95xKHoVGIRefjbNPakxeJMLV21PXkihZpK2srp0gavm4S7FPYp
025p7tevNu6YnRl3U6z9zOtIZyb8k6nbxa/22B4QFzp1jE/eEpm54mRxh9IL8CrG
wItuZxhmfV+JRQVo9edA/UynthG+19Otaw2hduncBzO66YevgjYLMd6OqTede3oy
67+/VPb46H5JQO2f8EsUbL7hfXXCKLXW7a/0MnE7IcbNXqaaCdqXUlhCLvjkb2Xf
6Cg3Xle5URwHv2TY1iLvdzMU4cylQ77m52/DTylLSMc9mI4fp7oqI5307fKjkc3V
R0tyid1/SV31xjzRIXMA2A9myXQp/wLoRnMqCCx7/+aWFicUj7kr79l4E9BoZMwO
c8Wt1BBXbVqKrA54mym3ddPFoaN4nPNRd0MTmYeXzKOFkpwk8D15KAhyp7sK3lhh
RmLwuzGSpZAuEwKjYHvi3RXSnA8FH+lx46w+fB3FWOq91ATb8XEtXkil3K8bQQvx
pSfVMSopJNmKFcqdGRRfxzqj/k1zakcFvjdwnbUqWTV1XUAmS42fK8cDfXgQpedu
hlb8GF8ki+D0awedtkA7ME5tR8wqXFiVkutCvnyguP4+tJyOwllLFRqu8p88IgaV
UIYOcUmDhY/o9Pqyre6NFjjzA6YXtvn6f7Es2MHOFPiDh1qPISy1FIyexf89HIH7
UjMED3G/LOIKZ86p+aNgKqtq2kQ8xApqUGm51T57PQQs9o9BxEVlG5TrzPJ7u+iV
gZzu0T6O4Ad0Kc2UE/EjkyYlfb3GCJIm+ptBRAXiGQF/KSZoAFOOxSjc2YSK4ahn
WrcQSjJImXwPibZzT6MtfRRAuh7xNp5DtlG5ccTFzBNvqQyC5H9fj87cP5t1PB6s
fu2YLv6hJJT2mgmN1wWhTn5AIZOsgRZwZ65WX5rOcPJyJBmb0zbKpMe2ztX4X3t3
ovmSitcftvhCKGBj5aYahVI0EYuYsymqyBxyEhPgAUxVstNpM8Uyb/SwthcmL+dY
HYJZx9zEJMMsTUtYSiCX2WRxlUqBK65pXt6GmZqZORwKaCL30lGioRNxZIQ8EWWs
WMipgrjG5jMeTk87qKStdVNZcLRXqXurIECmncqtjuxd+fNtsUHXnlKaL5FtfAKW
yHXC/FF8wz4Sb8RZjQ7NSJVHfWNJwPICa/75pG9+WVtrQRoLmZ4Bf4vIiB0LKxKy
b2NA1+rUa3B8ftrNzPx84VE8ftGZQxTi9mFUkTTV6iBbPbrgfzrVttnTavffyggM
Gb6mvqJqNwuEDtAm8qO8czok5JGpVY1SlxAuq/KApmy9gCUnsBsI63cgjyAWoc//
lH1rXRKOrPUl9FFCW8s6NJ24Z0OFz82rkopwaGZNgfVkutOWXUnzy9Ts6MfKajaY
9snW28C9sbTP6ilEO+pY+jOn63jaHZEFtB6e7FLN7A/DWZZMueGcuhkiIJ/MimQQ
D/a5/MYelGoAHt+o9sedRelp3FAqNBjjUu3QK7DjTZbpo6UqyMU/u5y59dGDMwmD
ZNn4vKaYFBTu5GBawV61hcI1tm0/GtERtY9LRF7IlEOp1rQdRjKYp+U6v8b765hp
55AXOa+gXakrKRL6yv3EqIxI73m0hQ4uKYR+/rhsvR5pdcOxWuumbYq+UbOoNVu4
J8PDpTtRV7LXSVjCkeoeIFP/asdPh8vM+ZZc5iQDOilyf+z6+58heSCU3VlWFWRw
uapQMbwoV2TiVDxmAX+lRXa7zCRiHBz5ttyLm7LEtL9SRbRB9MaalV6tG+92suqY
iyneV86OU18w+pL2IS9q4ZMh66+l4D89qXSka43teHNnIaiej1YyBaaczbdn1o5j
ADsizGhTgMtV6wWo1rCWU8qO8UjmV/VE60oDjAmKbSOyQOpEqRDJpEax8jwBges+
okHjgXZSLfxn3FcaT37eCDB6rLBnbqp1bvysuBLL8zPu/UYvXtdPCBmYYc8Jf02R
oWfck9mgPeevhoQZZ3mkrgyh5+7u2mdQSsFxCow/pOXA09Ax4Hb3DS+hLdHgU2/9
S9Yk0GBOi2KZjvkPKxwG2FGMSbXgR+ZpZzQgcSs17v6jUdu9FDrMIVTRUSUku1zc
PH/rjjyrHrp7SVKyd0mdwYrfd40N/K53XwzE+I8z1re3hQHc2LS3IXHlSrYL5b2s
lbliFxMyALYGUsag8ub2GWQ38ir+YKMoPas6QcL4CnUnRY84tAkwhJ5a3MmuovUJ
myu/MwdazGjEFtU/gzyl+tk+dHte9oaQROf1U83cplIwsUFVQM/TcRWUvkzziajS
p/U1M8ohnyHxWxNm+UQ4snObEZnoYS41U92HmJajFN7epiUDRhIyPCkGgysz3B1T
0u70aEd9BRHuoeoRoWaJXzto+Zx455eU8XUyxQgGGX1OEJpRSG3nOo13OcKlGeWf
IfLOi0mhgWF64jbZk/cqrv5VJtVwOHTf9EzZy4fdA59o6BTC835h0E/DQ9hhzkvQ
FTMfrLxu/N4+DJffWWP2PgSfmlP4Z0V3BCX1MYKj35McyXx4bMowvUmEXeN3cP8k
hT0RX7+6WykY45+1dkFdKSiWAgSK94iBAAwGA88P88EY28cuAwzQZHMc1Q+2xOMS
wAA6OatI8ykZeJOy94ghdwE+cEciHta1Msqkg8/KAURtf0cl/xvbr5ZGXYG+pre5
+f+sMOwEO+EbSGZ9ur1Cru9u4FIznHiUoLjX04KhNpAaxPhSvMaB6hP+iHjFs9qv
TsuDnylSBy9Cu/W1d+rbpPXWrUQ7BwbK7EY67aEkv0wrw0Auup8rpV9gTyvauwjd
wcvrHfA9HxClcsOX4NFDEUlO0JHKlIB087nFTxkwgwupV+lhjfsnAC3/EkC28asi
vmL2S6ef/aViz0yNdZAoa+4e3V46Bv3Yp4cXN5+huV2rhUaX3zZ7fSyxhgmTTSWg
XIfbZk4cdtftISgmKuGzzS4z0qSB/9Bdp5N/1qv4M3SBbxpdSjL+DKfLNM9V8Hc8
zD5qBa8jWMEsaGUvB8TFDeQ16WBuOQYEthH0GfFNBD5BWNDT63n1SjxeG1aj4/sJ
2b5PqYjZZWIDxPt3t2gcOLbb8JQQI+0i9nkkMKLOxBedDhBjwS4HoknjTluC37NU
rK+FArqOC9rbl6Qv+/CNlXAMX50RLkSara96Xa8R+vQ2G796j49PBMMqwCcPH9ET
Iq5IP1mh1BCmMvniF0rFn+m/E3gRYzY1WB5LUQBxJwudbzegT40Y8l0lH5EJoBqK
gAxh0CAe69ShijSDn9dm1TI1hDwl//GvuJab9nSbehse3dFak6qLk2dPRoHRfqQO
4y3aw5XitztCquEgQ40YnO42Nrun0cl5gepTTu0DZwSrwC5Yu3hfZmokWbkqY6Zh
B2S6avzS5kqptdISTGW4lqnJb1vuXhJm2nu8It4FhQ09Qvg7asHdOB1c348IVjhH
dnlsEaWVO9HKj6zOQe3bxntPnxJy/Z1yXu9IirOnWpI9ZdzB1CsvhHrGWJRdCMFE
vbg6yX+LEEWfR+JHOIlu5rl1+zx9OGJjAKiVFSPYpSCpRQQYGhTlZr6W9MZsrLpq
SeCDshOj7ySYDkUBjD0ofNfXqZosPxx7CKLdIYwotQEkdaAsx6NXhbPTjGd2RKfB
6geUROx26imYAs/fJ3jPk0NeuIEWRiEwVa0pr99k+rNxRGyanLGoHcRP/motgwKM
LA0J8mVfcDevFuIdmsqEx7PWRdPx+lTl4+nGjeVcEdJW5UpIUcyaUJFTK8adpa5D
q1UmwxNi5+AH3GLHssD3ZpRlMaTjiaA4P7Uio0cwhS2+IhW4nVT7w6j9Kpp+qITq
GTEgr+NeY1DJ4Y8h1NPBxHAyVSk1HX0iwc2h8SoOM9wLRQEbX5nPZPmWxfT2lYrE
c04/NcoPXNaxQYJXBwbYI6B0teaFlUC20ZfZC/KSKQB+2sA5RkYi7xAvBxmuNXRi
rKyrpVzDJba0+cprtcQl+p4IfVPeQaaS6ynI42oVeucUnA+58Onlup5DaWIJAWRV
korQNj/ww2tNBPHTJ08DGv0ztA3z086fsOnVXQXOyzKPcw7xXvA2j1fxOs5P0rFd
naK3qMtwCsH7Ehznsy2udQ0AjuE1r0lwziH4ljwWDcpokMyPZ9d8QmDnSRAcHyCX
IKbfSn6+7vNxKhpF0F0wXzNPzKd3yCPcmvyQ6kCdfq6jLJXmJwrQeNY2fxSB6n4h
uFTExRSaos/fjGJvGQSPv9dlqBIuhGyopaa8uY2HfDnI8w0eBx7zsqKUk5RUEIYj
BDNXDjqydL4ptcDkEMaKLofSFR9aQluzJoedwXPYZBPkZzbzOlh9zMrbDxQdBfiA
AvoJuO6biK1uY2nst9rh8f4xrhM+WPflc2YPzcwWihmKctvnfMtGzrWygpOPQGKZ
jYxPDhq0+Y37DRXjj5xqDWjSg35DMiRpisWnJD+ckA1I5Kj07fWpZMnWcMMAopeh
4D56v6RBNkGSfBEooX6w+ZHbvDrUuVEsFtUVqcqafCUrDGNSaYbDpiRbq1HAd2Zp
wxRDQL16gyruDmjAfPPGChn0l0QarDClK8irk944e6JJzGphpEA/mdMPi8xHzhDA
V/ZkAzHFZQZVGAzzDGM9akOPtoC4qT1/DaDw6yrlKJn7Z2Zbi/ihBKnKRnx5lQZm
J3GlQbHGYs74n9d2+PPyZBx9EgoRJOLJiL8oUBOI8IkwhnFcY8cVZgOvSLb2OqRu
2Le9eqU8rFFpiKrc393oWBZM2nl5TSzs3SPysXaPwyipBg06hs7QWi37uPMpClZd
NaL0vsa9vdrKr8+YkOy5MIoBbz3DxrW/Vu/l2g/oRB8EY3zSaFlo+2uO4FukJhoj
YRQh5H3tfFuO7tZW4gGcx6igeoLoYHw+BKKMY9aaPvcy/FM8mi26vJ3/bPqjAMrj
Ah9ukwu3vfLHUF98KcJ2nAt2OQnzmOxMMn2Po7hHyz0aiIPxV5cMMcsMYu0nIqlZ
YWm452AAlWZ+Kkplq2UqXxu8wT6FDOGMDWZt2D20HSxrM5LM5s1gmXIDqCvUFN8h
/vSoypeuk6C4vwC83rHSxW0O59Zs6Q2YL9JYJP3p5R3YyQXbcYTuttIkigD2Stbj
8UO9JorO2k+zwunIldOQ5h711sEZRGkELjLM940n72VfQiWyg2esyCSA1VH2PTpN
ufavYSZlf+O4s96IHS8bzCjsWiztzieRkQbCF8/l/7As+hLeu4BMhgC1atsrKNqj
XB8JlfiTCHw7Rc9fobKQLtD3dGvgMHObsgtOpzEkIgqfxSJ4TlBwFL8wEYQ+FPNf
bpPinv7r2HnBRKtqrMakdgm5eiLj2Vul4BSvsJX4B1tV93u6J7rM8oKNrB+SQDOK
MMd/g0l9qnNtjFqx3XicBSZLAtGd4PbcByfNH/vWoUaLRp7j9bfpq5Xgx0uHPJ7e
OLdAKF1YMd9RnRC0fHH6eJFi2RB5ER5/UWSp5tAFir0v2MShMxKMZIdvswDE1CGG
aMXrrryzrCSK1dAZHyX2nkCOJlQF5guqFr2A1M6LT2uhnRPtANSQhFrtd+mZnDRg
ssw31/jP6LV/U9bRtyLEI6GG7+tylMuAG+4jwZEFSpww0p7ytRkVtAxcybut5MrY
Nry8ymTePyykUtgjsFqEBHUsqQQQZPr4AjhpvU6hCe1vzY1+JqXjEOOCZ5aVXE3d
7PdwJQPjmLXsIyS1vd2FmOMqQy89W0BAnt0e47dpwB0K/tinovBdDraLc4Q72g6m
cV3V7KzIzL0D4v5QWGqPlCb3jsWGIAS8ab5kgRrBCpxv1iQF97Q53rMz0zGu9RwT
1CqwlcsWdTlfiRQ4Hy+IUIzkENOUcl7tVdblmT1YJFePeMQbZTzqLXt8gWt2Dx9i
5kC+1frntqPxU3l2NjmrSC9224217bTdrZGDGh87zSs8bEQrI2HQRGhMgOeF9A0E
cbtRRnT/e293GBy/Re1kW/m4OaC0F7lqv+VzCL3m8LX8yuDYCtsFTM/utq3+LQfV
+pXZpVuew8UFNsvwJSfXMRe2XMO5nIeKmW3Dcde3Gji2uXrmhaYl7qBpRu6PiNan
18vONy8D/04PzsmBLm9drAaRrW/s0s3p8lfULWItckolr6c6Lb2Ke6/gJI0hS9TZ
C2Q/b+zPe1suhiJtCvfe9HcJVOtHfq+dEa9lfpzSO9NGarHJJryv/o8In2TgUCKA
C7G2kZlZfq742Jiq+SyAxxrSCHd8pufi/dqGC5uHzC8u2FTKXjqlcvSDUkJODC0c
VQUADzVGhQyO7BPZ/HzUSIffX53CIXtv+rHzwhj+hg8oa0m/jSz48Ul/WWjSnkWc
G8nZHW4xpK8DywKOddQ29AW5k/zChggvk+AD5eYgnWVfjAyLdJCya/eT3rDB1kOH
EhViwkYLklZepAvVSdOj7nBKPAoZmj9fI09AKn9234NuBnUQcm+Rv/sT46VFcSwj
aPjtodvSQb1d3PLmcP63jLWYH85slzL6HmhrtkfEadSeDn7gCukN/Kf2oNJQoBbE
/axK20KqWdSTjqSTX4/eqd9QBRzPQW00pHI1KOtWfZioAHH3sw1jMvdh4u9HIZJU
k8gGFwA7JEiIoOG/tJbJFej6OYqjUJKdxnlARjtR/6zuRv0yogoDaQBfyVqmDOmr
KgPdgxNSCrUUC1J+NbbxfAH4BjpxIrroCvOHKXkEEGYXV4ZK+gBaIo19QydcZuTJ
31Z0EZ9VsXUfo3HrB0/2byIZ6T7CnxVBffcVEHVmuQzNbVrNwm0aU9QH1kRH+uuc
czGHEw5D46XnxeW/YF/Fbg12ncgs587RmewlYyc0lNAofC+saHefbl38U4a2D4S1
w/iA4f14IW06gsGWn9vu3728zMUNNTPgjSWeqoDbYGjMFasigzb4mPxFK2tak3VV
0nfFjjiJWRMJ0A+A68DWwmnyVijeRa1hclXxUwBJdkrAzhbBEs6Nn6hEOED1Qm0A
eStwD18VzW3Shnp65EdqNCyPJUfV9r7rLqiD1Vd1G2uMleLP39ZfhM7aVD4YO7AC
lLEFzZYkKzJaU0TrFO2iwVNULWVSHt8SshtUv8FqNIpm6pngMH4lyctfEkHUUi9R
Cqeb3xg18lU69BYVbE8pt20CayvGsAI+DyKJo4y8W+CfhEvzIUIwBMr9I82ZvoFp
8XAg5s3RD0VrvFR5l9ovec3H6tVZWuNJiqj0OWCgy3UQZQT3dh38liINvlCbEZMp
aS2bVyjQMuHeBnYA7Tr+laihTARnlMDHz0Ftlbve3RVGB7jjuEs8aN/OxNgvhYOs
JvPrvBu5x43HZFJ2KbpM1eWRAyEAno3tS3U/cL7PnuErtfeiyYO7Fm0DV3NCHtvD
tUNTc/eQX3K9FFQGTlH6yMAVdoRYAWd47BYazDlL2ktpJ1XO1eVw4Uk6zwQcyGUf
TgDg8gJzuqyNGnJrUSg/opZmXfoS0bW5PRzxtwTBp7zfg5fu28qX9DOpxd1Mu0YP
9gU7uPvzyzYaa9K0KXFHl86K6nQjYPzgZ42CkXrUiSDrNufqDuH2eNCdDqVAhCn6
fZdHi8khMRMV+0T9mjDTqp6dK/5wyAKNBfI45mdtrd3/QBtuqvpUq5dyxgPomQ56
981XlmrDvNVZS/ox12Va8DvBQ2G3Qzfdau1qOLq35uN1bc8o4EoVwHy/+2pc0qH4
nVTr/ZpEjIdC4WFcla/BUPuB3v7ol5G57tSZqnFGTQkoPka9Iiv3OQUnv23DEz6s
b5qBkxsLSIPjQHZOzcGbRDC6TN41eKaa/CQG2O8NIhol/ogmQjiTnUoPTeijWfPS
q6b+oUi4jo9RI3uVeEN4mhJW+oFfG3awFbsmoCpUaHmeyeTxwAB0H1ja97XVBDF3
7nMEjGIGCOiBGcVLiiN4fmzN5799d6LnHDp2nWk3JJmkdSkgnmMsmtmoue/i6Jxw
4UvZpi4pwJeidQ6yMkAjOJ0wP2LuFeAYADF1wtOGlU8FhkxD/8kdFjwP1X5EUIQw
V2luSTsts1eN5dAw9xNpbeuXNrY0eYo2rLMZPSDSdS/C2KCCCCUw/QBDwhavW8LX
x0x7qcAiXwl02EAmQZzRDBCVxgeoCTiCVybqMfog5vGtlFQQtcvlFabZybJriKxr
MbnLoNwjyQaSIw8AI1zUrZL9ZMpkaf7dK+D+yKtg5v7nRvQctp8XUHKNeMEqBdAE
zmpkhrzPEVSvrH4saeI55qO8WIacbgh1gchlRRL/sQ2YmWI0iGRPO6UEexpTqmt3
UZfq1S2DkDV2wNoL4QIM256BJHudsu8urie7FMk3JdF/ocrGRplcmS0WVUQdVAGf
tJ2P/awphMc6Ih3c2+1LSYNtf31QdUBRBM1bbIMjU7ZGS15dJy8pDAvdyg3A3htV
5fWThxu2YJH1+p0PX2izBjfZ1CZVA51VVNoc1ymVnCzi5Cj6pxbzaApfIoxRajwL
uSC4xAKzXbNyQ1W1n1K2tfxT/nyn/SjWHa82g9pwexySHIkU65cYLccjz7TjIHWP
xTy5ZFFMVSTyfefjPXmnjjDAJjLFN81y/rfDoM1pBycCLuOxWP/PB7cncjEZnImw
96YN36vwq72aWQr4dxRgknSldeUOuaLCex4G10dic4kOPAfCaUTaO2vLc+siXZvk
WS2kmkaSFI9zv0r536vSZKx5E3Pxxe1LyRlQUQgLxdq0TwicbGJo9hWIm5BChUL6
2qKWy51bTEC41BlAS086+UfRGsl0BO2MET/4Y1Q+WFEKIuCxtvBXcQ43PFL80dYw
6wdN9OjEYTNA3fpyiTtZU7uMwJcJdFL+0xHOs8b5c+MwvFOIVGnhyqJVOH503hfe
Hpd9MVWeZ6H819Fl6J4tDzP2HmKk/iXgpNw1zwiLAb6Ilv4CvCXI+IdnYclkjRm7
HrO4b3LooPgDr+EUTcHAoDFRA9iS/oUrhMg2pVoct4gqHLOdxXR95a4QFnFjR6uD
1Pv3bHy0R07CvgCVI73HZq1kpD3YgWG2iw3/YBYeiw4fT/9Xz7VqMKmjYhHxk3Ee
i/8Xn7DkG14k5+/1vqUbOUZPLpoyNm6TgHfH7ZDQ9n5phzN4fatjJhSWvMbZRFk5
VOAbJKsAPIsNxfG5IAQsram7fQuw0P1vVsEgREOQ6U/9p/wZLoHaP6UBbwjhK2m2
iIbRc9csI/5gy1xhAzNXoLPHmSnL23I54+rCIWlTC1V6bCSZ9V2UG/rws0s9MkLw
0DqodRIE0Vb/N83Mh5kNxBhJE0jd2e8aGycpZDCFuxZQspJ1Tv0/py0CfKxohZWC
tHbKJTlCTWj6tuqMFWbxu2h6Z8EbWtY9RlGbnBm87DBvO1jx7SMCcHE9BEYVvbF6
GGKwaYfvfQlthjA9ZBdhSiwhdtZFUKSPLpW85ABDqSFXWr8wW+59mORgViFwNamG
LZZX+CcGLowQH6PzpB+rZncIxWZUZTEdOOwqCtVMj+l+R5NOcCuobMewLWZAjv17
JgbQrib4BVGn/JIKk+rRDl3vq60nt63gAKl2DuinXbiD8Zper/H3kZixNTXEyl6x
g8LWh+cK6dG6EkidIcyJLPikClnXXL0vo+/b39sIJrXosvkJllroM0JzSWzaSGxC
bp2hoRF7ANTjNWpVZyNfOvn1f+gYjJkxrCVk5ZxFkHJlMw12u4T27+Cm2MaHPhUP
9dIaKZeR2JSYi7uQoycgDZerdV5r4ZefyqFqzeXUZgOvfcycjRV1YrCHrC6lCFKe
OJfQPFL8yGHHR6OS6FDAzUy4I5zoQ7JccqR7zFu6spCtbevcxjJM298Jwwijk0Gs
QhxYUqvNQF2XcDvPTz97V+2brfzNng732paDLv9l3MjoJJW+ec27IVEAoNl2AWBb
yXbbAWhDY1uSEs45hTKtZ4ojWZxcou5H2RXzPC2dyIjIIVRfY1yBTvyIlIFbXAY5
1IpCZ/Ank5/ZOqIg2jLCQVX+roDshxOaAnbHuDJI5qQsCGOkPqsX5xFDpkKHvRUS
6xBvAtWTLyB53mfY5fVIa/V3uDYuAkNodlCwVo21TuKGP9idlnrn784FgbB9zrOM
GQSGNEYBb1ZRPhhDsuWyeFhKcPXdsr5u0GzmKCnnxrBJWq47nm64ayOVQnekDiOT
qSrAusZGiSrcbXoQCK0WnePDpBCVm9cojBnv6iEyBZYch4JvCcQNdaiWzKWUz5u6
inALzN/jU1+C4V/L+by6rXmMbvZLDiLDiQ194cn3kmXa6hUt0ZsYxRdVnzWHkL9y
mEYHnzCObG9v5QllqAOd6zH+kC+O6V/2846JNc3UI4Rb87VhA9xO5jMg+kBkHq/Q
f9uXwWgYE2GyY4C9TCsykxrywkJKUN40VY7Op36DMekOVz5j9D+LnAJhPvHdrDSo
KxgRM0W1XfLBpd2Iu8PF7HK2x9MNYie+Ock46PDJXsWw3QkIogmnbNw2R/SURzpL
SiAMyP+EC3ydzWYIjZiFEHkDpubCbmPIdwGA1LKIkwUlVFicnVosqkWjbkXyI90+
Fo4vqdShNaSwVMgXyC8KdPHpT42E33c39fyxF2V7B7IdJWJUdMI2FvWYCgT8n75B
VAqLAcxUOBa4M22rJuA0fy7mqyFoD3J0wl/SqT390WSzEcgQrjX+o+XlZeuMZ0ey
r8sg2Ogi88Lkh4YLb4u+fmb99YHE0EOSppavoal1yAf/36x+DTvwG+9FRI3+Iany
m+qD+Co+WXcM2fP2nyHiXBlUrMo46h38HXiv8wUa9j73Gtc/2IB/kzRFPpjvl+EZ
DUs03H2FiI9IOXau2Y3tZMY1rmsb8fH5y6FbZDJXy4ouhDsJqDNGzrLcBT+WibMk
GRNR+ENUNZkFI8Dk9zx7x/oRzgmdDfnwWrmA0mHFDQCpkTOXZF91GLZua6cC6oh1
kWDY3xdTC9uvoxYvKxOXRUUTxQJ6FmVVdX57Q5I1HU1Ui4oBUyJhHcvsFX+u5O4m
bcnx+E34HHWxJnw+WRSrTQXyKkrRPJ/NzMCaWpd/Gaws3olkTYl1DWsd5p0OpTm4
dOWZa4nqtoV/wHra8k1vkeiEJCVk701MhCfXYzuSRlAKUE0SMFcnL9YGnvjJsCG0
TuTK2HaXCMPUVINTzm6ZzUn6zmqYSHYm3LyHGOcgJZBRr7k8TXIswtkd57dHP005
WRKAoAcDIchilFF6B/xZ3OVzSZ8gwc9BArXogV1UbyAFB48jQBSMM/UZ6cDl9MEU
7ktTajJtxCxcr+UwyjjmziL3fBJ3i8nAv4brbACjyCcgQ3TBygGk9K27i8cY6zRM
/4BWdgLWcBGNLEpnHyLdulZo+9nkJ60PLu/VII1NIlMNbi+xuUk8NmL46TT2PM1k
8ZDk9ieVPILolO6B45TQeXVAuesvnH3+SiPzMagT4pFszx897Y/+iOvL2GwyJh+q
hpsKTnShc2HSejhWAm4hbPHrwzR+bW8lvU8H616AC9PLcBosyzaUF1cRUOt4THNh
t8AeKhoZSuqq8Rc1X6QFECTPN/ZXuoZ/YCzTvexx7NqEJJ5Th16wYNDmhwksr6ju
vYLvbt9HoyqBK1awhOFNTdnUZ/YD50/NMBTAw75FLBg62MB+T3cX5EfbN7S71Q1/
iNSwPv95QHfR5mF4muaCqe4BNO4/+Fhy6s0MGUsckzJV+Jve37/kigTxT0Z6ONdt
y3x90dtOQV1S8xonqVEdDJxFt3UQUW23Ie7rezsAbEU9fU5YOpRYenkmtxSL84/g
GkL1JqyTIO0qdrVpStuyIQ2SnV4AB8G0qEEHxUL+gv2U9R5yhj5wE7bPWGN0i5uW
8WSI1I1Y2JB1ttMUQf3Jc/jWD4GEr64Ou2elWxhujBX9joLg6RGHzAw7AM/anjN4
zvJtY6lJlWt8FT24+UT9e9ZfQd2OFYJNfUk2ilb9F+JUMZ34tVdycgkH99lA3vaF
8Zwd67k4WLwMvSdnHZ+7FcsrzyKnSD+1BcFMy/OjUslhp1GvOQVrHvILM7l3kCU+
/JbQ85N9HgMMpjVzmpS6Q0VT9+qEmlfDAXRj4LmsQ/h+Q/t1Zcn+Tty5m/7cODH2
UvY0DDLlPEYrreb8YAFtjB5eEYiGmpd/hDQyLjjb6NGdjDQbSV9sLTKdJt3whZDL
UtPMWWNNoEukFZNIJMt4Nn9L40PZnbcFI3KwPxC99+LTPFEaw5lPR9you7EfbF1f
TBzW+qOGf4bPkaQeya/we6FZcE0C+EV4g63k3pMgYfgd4m7L0WY2OE3mnBS+vYwm
RoVzpwUwJLz7/3ZmS1Or8yEKnsRuUfO1CSKdhdZHfwPW0aCg7JSPdacgSUlKPOaK
6JM6jdP8aP3NJSZWCikA33EMQatjFL0Dmqfg6S/ykujYj6nb9V/uomD1iij37Wey
ztjxvxTM3LlZ2n8FZu57dlqCsAvyBk2uHFxnYooLZOyPgB7KtZIzltwSU4Vp8vqf
6ttiUXl/rgAGmAn/D1Uzps18jgsxOfFc2LIZx8wwJ3Q8arIZxo6FjBsfaduQf9Xl
ZmOesKKHsbeUoKvf12Qc5TvtzLuXiMWozoH839DNb69WpLUPLE1RoSJsCdXE+jjL
Jos3vY0oHiGA0HxAJ5azlMKXsjeraxMXLQV98A/W35r6zKhL+elnI2JCm8mPKkAb
iHfqz86tUk8GziBdo4szVplslq6X3JKEGiOeGosuaJ4nwDkroatW5DLzOU/7zKQh
vHYcw79ogLwIMtDaWG8qRhmknHQ0PdeA65adlQkXNKE20BeVSh9o+GEgNaVT5rnD
JI9EFkCnETTEQuF3Eo31xxdquru+QujCSzJZwXmC3V6JPv9mxNJgBFm8hKyvV41/
7B1RX3zF0o39bYgccbvSbzNnvFH5ut9vtVQne9pJu6hyF0CBO4Xgvte/F05bkLpn
lsdTwtw6MKg/VhVZfSj1FxOD2QbnOB7tLajW6GFoO7fLaUALQzNcGom27xJQnecT
N4WClPYCn6RS1HTCh1PCwQ3tGXbCYQMCTlfChoBnpioDVdTgIw7VHhiRW1rErB0s
uu/PctTHidEPqeQmWLKBdIJ0ikXTRWMAD4O5oamecmXyHIbAj5K/BGnC5uEIA9CZ
bV4c703u3jiQDIyybDLe795KXZAqaLtd23VrCn31JSMBXeJkffhFev+lbHn0Jqnj
fOSRfZZ3sA+Fm9SNeprrCoPOYI42Xs7OfNQnewmrN3CSZUNsc9EVR6UVPYiQwyHQ
MAI6/YfRyiFWcorfkzudbaTM3vQb0xcGWqZsd42IIgTILbH7iLRNonGEGZ3fNNoC
kKixqilxyjjWEUN6AlvFwgY5u40z8E9L6KIBLFzu2YcVp7ic3qoXf+K2cGoIcYK8
xRCPNA8DhBeKMfNWxhHvoXEajE8VdeKDzBUUzn4SD5QMDDdZNd00deo5EXQRlLCc
aZfdbPp931HMN2Vk7bva2LNbY3HG2DZ8y/qBU/m/dROtpSekImCPk9PAPFeRf21h
WIQyDJpNtsT5KkcCtWsf8DqLBlXNMD0Ih7+ztxRTg9usRpPsATqj1F3FEZ6i8sDD
bszUbt8mVOgjGZeafhxWIIgFTYFJChV+4JGeuuo6GKyfhs68XtCrO/EEvt8sFgDO
Psaf99ZPg9a2XnJmrNq9BHF8QJmDvqWLwaw7W1SJEo+6wbce3NTQEazQjgHVghAG
jeJ/RkTr9J+Xu3aNd41fg8HEv89vw+WhNkhwsKrt5NNSon6K/9YuY/Hb27Zd8YE0
SyNq6TIjA1LtVDYqravgtkgkNqT3jcvap42iGxpxLu3EAoUMKPB0EVoX3amrnF/S
SHA92gYRp9RHWtMst0fA+CbrNXcMJGPo0Wa14uhaYFLC5KwIJsY41/uxLyrsZBg6
50baofXue9NPSETlF90PAsjKHWeIDviWfQdSugs/XQquTd3zOjyTkeuR7Fv4NVZs
F0fPs6uDoohWu2Uf5XpDiMh3plDjkuQrhPQOEaO3VAxyNG6lMkJg6mZb+OTONzRC
A5k+/DF1I0FhYx21CnWYHZS9rctGjrSEeAbr8BePVDK25IEK5e6if7Q8/04U54mT
s8iuhENzrg0F63s76wlfZP5iONROsJ9iuJjoc8Plw2MosnLfy9GN1Tuk8asLrl8D
y+O2Hmv6tJGnw0+/QigGtBRJe3oiY3Gax34TqXww8rA8rFddeL3P4KwIFcPYy1q6
T+3TNKYiSJS9Peju0pBfS4iEWkvRx1/BzO1IdpUIF0U3Ax7PRMJ4BmRo8888LldL
oEHbg6JIep+/TMsNGkQNIllNWdvN6KiAutuVXIBjqo10kjNWP4DxZkG1mYgW2aLa
d2JYB/Ar0tiAfxswM7IiZcBULn9rTAyI1KA06bVl5wz1C+tIRKqbCi3ChSSKGwta
99RRi6ptOGQ5YBT0XP3uIEcZodsPoeuofGHPeErurFx86C7sAZgvgsPpZpqOi+Rn
9vCOQPlG+GS6jX9v76TX62J3HH6m5LB5OIK1qFwARc7qVYBQP8BBbgLi1p9qZ5fq
/N7DY1OK+Tl7OXhcUHZ51MAOPmI8hcTiEpgGzafqHACAxUnfuh/TkXICTgISVyym
vazkV+v7xeLo9K9MtPF+2yc9e5D2uaK183U9ZyQx9/tzC0kKb1liui70d6otsM4S
4/TWWN40fdZVh28U2AjJ1AN8SIdba3Q0OkGoXMDcGrVyeOW+vBkBN5qx1IRK4uQY
qan0WFt6KIekWdNG7d81KjEKX3TtmUCH2RWgZe36HMlJ5Ws4PlC8m6mcFgPK6opK
x2ZgpMmhnrnu7K+x9hTQgY7lQLw8470xUHRYUB4G2MFAmg0P8itJfvYIJLtdZ1A3
K3VRiWgJTVaySVtKGqcQynKoLouwUGFOPgE3ZN+KOLZpRNNBTENgRslUwHVThqd7
FC7/uEZoCRK484gQKtjQ5D7bfn7tiL/74QZdu4LbeOyrKtBAKPzrP9F+3lsZc6sJ
vcgM8D4dUhQQIeoX805gPE6lcz1KYrHq/S22OPNFkH9IRWy8OD+345l3TGJuvSco
8X+02+QWP8ay0EE7Yj6aq0Y4L3xGvFvx4v6AQLwzaFstz7kr/jwm3Zf9VfIQLTS3
t7gqHoUYXfh1KZ/Nmxss1Hjs+5zc/d3j+Gpe5+/O7pwXWA8+IaSXOERS7wZB6qhR
6NilHvrBncO013PIP+uD9OuhZ6L2UpCDfBBY2USOX7pRJSQ9a/bXTzHsRPGJ3a8A
BoHfw4kpz4KMlAXcbHPAXXyHk9YYPIPajGch4qvs6m0/SMNG3qY6gQErEJpIUmLa
/8kOo7wzm7sjKHMcIg47xS6LwDQXpJfR18ddKj8RlxORY3Fy7h3tsHOGz89A329J
LPDbfg4w0jgxk5V//+zBe/jHQVyuzo5CbJwex7oNy026Yq+IqQcuNSxCPa16VWhs
M86u/DRerpKl4hm0IzbO7mPw0i0Cm4e+oh19cs4CxYp+teEEyGUdkNH1bw865Eig
aNeOLGMVyuL3m4P1SAra9OhUfnYDcWZpqbOm5Xj9b+q93D9RLNETC2liGBDuQZ2/
v8bQSw3Sl9HQ9ud48nDTSmeo0XX5W6yA7cBXk3/LSm3KCX1V3GVyOHNposNCNYJB
089PMxW55zjEs2XMVlUk1Jm8GoL7uMaV3kCyqzzdZDIUk7ZEMCLaxwnUPjb1lLg0
CNRloklFQ62R5sKQ3LRt7MGDGEqhBUZXVaTCZryV/41O5mXBZg7MVKcldMXCIR1G
waxx7/yuSFYTLjHvxu7D/M7Mjvwq1EM0Ymyt9UG0lnZXv63UuG8gmfuoen2JO463
54iwcmk91EIk0N7EHtqsSzR2i+50//9w65HxUasvXUQd036JT88LzSljM9VW4jV2
tM571BeZBbs8SHqZUwPS7bOg6yZBaLDomjAxBawuNUIVr/7wHK15U+Yei2MA7QhB
HpuI6lJyQsEL21PxHXyVCJmoiMfOSaJj8B/qUdAPtnJ2JIdaSNHOJAgf3TqabUAd
+E0t9SKoO/UsqeDJieXg1Rv/1zRm+X3q0bdMsFxkoYy1lTYUwBCYnV78Nu0O3QtR
hoDmXKHZ/bsM6kGeFneGpy9ftqY/sh6YExPHXaO77t4YjIZtK3n7z0+vAHU40F/8
necOj6TX2phM8bSvqK4fVCoJalLt4K3m5ZOCkZ22q7GgqYm3by/sfvQkatStoTut
FK1voYhlhbqwBFP01T5cpqNqq2Zamysnse6U+vtX5snoMYEmMNDEXLtBWN3NMCb/
6aVoYQznD4MOlDKzqxtvFXikTNY3jz7NrEtHz0D/0IIBYuVezkcWAeFL5g2d0fAD
DgBsYbiRTTlw+Nn+sUG743KjJitGixRuFgO6TsHxZ95v783OSD+4rrmLwhpcb7t6
MbDK0DdSCwCyN5JADoXAD5nVH5hN4bL+EUcew0qhgDTc3tAl956T5vJRm5qjTy4E
dZ4QkirjNkeACsxJXJv+wQL8fCvsOqzc00Ql+NY1w3wY8Dz2KWGLjRhRRUSOvWC3
hz03tKSY/3w9vKZ3PHR4Vun4fk9kEeT2oZC7zcgtfJRHf7v5Kiu2QD9VwxFr80Ei
o+GeZxSpnhcv8G3QF/9BUqzYwaW4cnGf//5p0eJnzh5AbCzjiglUrrUUb5Tf/hWY
w9LR76Xr8VxZE2GXM7Wwuw0fJYSWwtFmXYEowzma0vv4kGnU8Sbo0j2t3M+byeMD
JCzJ43FPHx0qBZuPyhUV0IiSZkcP/x01DOickT+8YPD3HyDEqsnlt5x1/y4KMK86
vI7tcFnrvmmptG4JHgzNk8OaIc+dfStvgCix8elnNCVS5fCMt/2gEIKNWXZDEfDt
adOabfEc5S8Q+vrB2PEXJuVK3IQgD92sJPwUh4peMORZ9Ez6587zMytG1r5kVr43
k5Sn/1tjYH84fpr7ddpAuvQbeLF7tcmPx3s7Udg33ketKE3jGCaqjHppdGntLkog
21m5n+iwqX/Q7Vy34hM51XQFdldSV/mJSd6wFkkKxI9QGzdVB+9F2bOPHaXvsKfC
gHFIcCbpiOxlDIfe35sIEfejTVuhcTsK96xA0Pud9rliNFXfRFZTAQR9gFwjzv8h
Eih9Se1gRYwzFGBYTX+ipxRjYUNhC6CpepuFz+o6wCQkOkzNxUTJjuC+nqfZmnzt
ZFYpX77W2d0U8NanjY4UnKPsNT1V/2W6b6/0n/YREgmS4hKVPc7tQrwui/Vsi4R8
MNfna1hntwQ46WunQOLCx0lf76CdNUeApKR484s990HZB0SC15o6g6/5a6kXEpl5
URDU/c/UnS8S9oRkKdH0Nm4jLmQvz5GWc5kFnmv5XjqmdhbRPALqgUGP42WBRocJ
aYukG0wFPvFdoYgJzDKyHKtHX0mzof60dQxt2Lcshdcy2HYlnVAF7GJWoCukGX9Q
uMJsxLWZk9dAvh/KcL2N3T107s6XrxH22Q70zwVGmkgzwKjVP4pbCl+Es+c9+xNZ
eEPy88YOSHgIQPsc0EmvO4PW9ay82BGij2PcW7PbOA5DFr43RhyemwLqE5eEJ4IW
Bc9eouRs5OVs5QjyFVCkcvW8EV2KvKp4aUA9ADHZ/rLOcnIFjhk+Ae9vlSC7mhXL
1R151mZk7HmdXSXz/IQo3OnAFUvGxA7WEbEbQ3vJ6iE8I0TUUfz+ngeRTVNB1MMR
hAnJzHTqHmNOGR82T64RMW5pkhihPJIPqb+kUBIKnG3x4oJrg6llr1DlM1VowZcw
lSGORHSVMAONcGHHYHHJd+FRziziEzQQ8KhVX78RAxzeZ22ia0tySsYhMqOTUKQi
ip+WvjxNCR9iHNb52ORNdjaiCuYe4jbm7pBCihYjpj4EI8BREVq56Rl3iD2iRaRG
S5J6CfELm43zHvp+QjVfpTvOj9nOcGe7YDbomUVpm3M0f46dzuRCpGTgHL4qQOcC
gB21+65g0DV3n941wu/2Y1k+fIFYXHhexpvyQhK5PP80QAtHKdLtrg/BYKeKV1qz
NbhCSt3e26zt+XpwzaEAVuu+v7FQHgYnmEbhHN4roc2IiXKCp+UrCCZf7rjzdygx
Sy+oqDcndYn7CokvNLJZoW/Vh7oFEuaIv8iMOX9U4A6WdetxH1T6Ay8y1tI697Z/
Xe2SJfMlvlJQEJmHSKV13jWaFakL9l+1cuWFC2fC1kv/D9U/RSxWCfXo/FqwaEvu
KnWED8G/wO8hggVPBIynF15n5iDhXyRzBXY1+PgV6v5eLcjWMSwRD5rfEedsMv4b
su9RQYY28H2it7YoYn6buRRgfuPSc5ArGvBajU+a326OoIVVKj5n63fURos8lsNE
Hq0nm9tdz0KzbIWVMNeIn911qatQsevYbf1PK1tPRsTk/BDitoS5zBjdKZ2ewAHO
zFdLPoz6Q///S+W86qLPSi7m2PT7v9loVs0+P7rYjJ3A736e1J7s7/CWWLftCT79
E4q9Aj26uAi9H3t8gUNEQoXSNhXe7nzGWiQlMnewAE0ZS0UsgEjPbdH73J26MyUe
mUyFKt8uHoUufNdWb45B42ujj591H+Lv5Wlb7+NcstUbVraShpdY23NjIMLwvYDm
5JPdyWSFHIefF8UUuoZ4qFBsDyKOk/620lH6Y/O/E1CpjJ4Dk7UG1uVVcxNqVfaA
o/UrCSoGXDNOM6JRQpP3U4uEZFuioGuAJp24UxI+E782iMWHKxTQdGjnXz9MAhTr
u2ozb4peIxyXjmagrOEfw2GjwfOvNhZARmdtEWIg+kq1igwzKKX+cO9TVkTNvTcN
fBFxJvVGWlg5C1sgcZnWoZxmj/AvLuRI5MrtQkfKdhvmDdoH9zHJc5FW9uo634gf
a59pESwEViLudCUhfuierEZnjkqHjPHXKqcQf9VqD9dB3VfhYNG8VCBaUwTTN4bn
zrVj3IXmdzqu6AYpMye57sseFwRRz2LSlz6ACZQEIIUAvggQbiFInwI75zCxxuyA
i6QmG57LjG+G/PTTl3TtX40lxlx8zXoeTTht69lVWqDFGaoBSxgfPeLNGmZInSck
hzhUIrABtKAdiZYCOitHoLdSYf8vYg+0uf6/BXsmQ5T1f4drFfNVrpVRNpuyPvyt
0c4Ed5eIqImL/8eavIEvsRCehH/P22eh2FKu6XZgr7xNXilU0mLSZmUgkiHVfhpn
6L2ONwP/9ooFXeXNKAHTXYKigK0bouNARiDpxhVyQ6XWhRkqk5h4LkgSs2uKjoHM
+lnfaUU7OxvQs9ttMfSGDDdanhZa6/D9KnI84RVfGQ48DdM5HO8xppWsOc2JUIY+
0DIaqf7qTlsRpd9WHTkTH+7QNyF4Hxb3WAIh8+uTjNwpPZwpPVsDD40s9Y0EDS2P
d971Pz4NanzPAcHvoknEiPPoGmTB3sUNPJAT8cmR9q7pbRJDk9KhxbT6onm8ynto
QQYHwhiwxihmHaSa676WT5xepW29EXMCGJ5tixkL78x+J2j5dDK1jkofRDjzzFuM
JQp384fo6HmAEaHU0XnrT2nPyqFhBeIGWvTJGc2a4er+Fkn/Gi45GkihV3whlVGT
zzpzfBJP+sYSHlXQZx+NQPonYitT7LRk2TXSt3qvF+Eefg1Jj3JKCDPeiwNnJhn6
4Yjava7ezjgp7iGK51Espqh9jsUd/ppUI+DqfbtsiG5o0bvKAbjQKhU2pCcWSJEM
aVmpV9XrQlYczcdp8gq9UywGPQdYELJ8JYXIQB457P6qT13K72eNNNP2JolryaDE
pgsOpEF1/A9KGUlD7/02UjaB9cw8NhYtVKlEpwULNWduz1OgKA3LoASTYvDCMJ2y
FoJhM/OB0hJ8GN+rdd2huZBAKWY4TLGo8L70VDpPLkBrs5Jud6sWbqnMqQwVtdgt
+OPUxRv0+kx1Sd2uxI8XJdlcq6aMPC9PRVXMHoMZlKEHHbUB0nqiI1ri8wYomxpa
/L3wv2ZA1ViscKQVZCGuAp4hbhXW5RT/D+ogiVLuGZUgnPnOr3b5dLJEMCF8Mj0s
F/e8eHZKo9xaxM/m9agiw1rlLlqvtIuVIQw/gX+EQW/uADL6WbshuVPnTuVz9uht
P+ykuuIn5bMHj88vQR79Ncxwh1N1bJeQDyPE/+uwucX+TcmdlBVmZZUGXSXvqCU2
c46R7QL7bi2rVRhzpEFTu2oDaCKWJ9WsfO1cKo7h4KmRtqkOJ4WRDaW/6TMeJv8P
a8FimEK+fiqNfI56pgMCBYpmZ+XRbfUvSPPJwe6e2nD4/1gWridO4KEHRcXDtfFZ
Ew8wrag1A2o/8Wif0E7g9nNy6br6ZZC6qxA5io41++iCLrEp4UW4PRAAgWaQcFLI
Eu1iL5Sd53bP8oesH0JCxEtQmXskKIw/sDw/qBu7XyCp3MHY7NR2lJjcEuOQUYj1
KbF6O4Nso1wiSuVmJCh11nK3LlormpenEtWzE46WHukqGBvWjRRrAxU7yZjMxIHf
1pNyEY6zVWawclfM9z53g1vEpCVE+S7mEU3KEdNoZaF0Pj17oU5T4eTtgqzAINjo
axgaTF+3AbUkAxNWSFsmFfwNSguTNOIK5C2lAKgv5/UzsdWA7HqQGRjUS0u/TGrN
Po2FHY8XjgdxU4yIXU+oUsM8lF2zqEVLM2NiuAKN0+hR8IPm3Su8JEPenHS+QWle
xeX3UCO2/UbIgpvE804YPAX6mdFi0guYAyth3ZsKTOtFaSlpBLLZlRByqUxgU1w4
uwCAAtH7osp8QApalIDyTF7uw3d8hZLXjw8CBCZHYVHyGr0MTzo7npF0K1MeUlCL
x+cSI+IoFvEPb/dChu9nAmNrADDGvR4p+1hAWXHa4jwo5ZkLRwsj3e5GOrAWAp0n
ubYZUVm457UKVcJZfj7LCtt+JsOAAWsp58VtZ0lmfSkavAhQ/PlwbggKXs3Qwbai
ZZQUZalgwsA5cfQBJwNznAoWM/6fxsjsat8s/4G1ehcAj214VnmaLsShx+UwJ0NC
MM2hE0XMcBH+6QKj7PEUEfThTLMlQi1CgjPesjaas10++UWg8ZX6pe/dC5lzUQXY
yfdUZZ7TYrG+4KpZZbEKFI2yu/O/gYmbyHJTyJk1IM2ViGoA8S5L0jamW6iVyBQX
6vjGetKKaTpOLK9MvVJH8eAoXRjK8x6EEzmwcaq+TBM79Ec5NP/y+jqKLZVy5upU
pUxtRqskl3Sg27nlD1Xt+jDLukHeBDPMylqIShYyJeuOkVnLvve2yS9Ugh0V7OfV
onvHSbzi7MJ9ubFiFeNZqUP7xPIMtA/p9s5Ts6nxGH38eo2CUNcJT0rSu1Ykpvgc
icO9d9EikR1DOYvbvIFJpyKsKwENcrvzqP0JMox10SEotN+3B9klTjAYnv8FSVSQ
bNnBDqjFjUQKXTAvtP7c15weQqWibxn8XML8XmMb7JISoLN8MpdjR4p/GQ7HaI05
xN6SFVYy52fIkV9XJh+T/yjx4xVRzGh1dIledaeeex8uaFF4l3vT0OVbreEfjiyi
wdFyg664m9kcUiqQckd6iG/dg3wzsV0oH8gfayYH/UVB2R2RXvEClCK8OBZLTrMx
hpJbCRkv3Op+gHh4bNc/BAimaKP+uds0nIeelAzU+Yf8pfo4mOpEn0nF3szqkh5U
0slsuvM9fzIAeChGiBbDrCZ3sG10n4CDxRPDv/aEvTY/vIHw7qnbJIbjhMspPVj3
+lm8T72suNLonDW9yyvKAhza5o99bcjJ9y7MpyT55jM5uwU+Fjh0aaurGv4/iTjR
f0LqjmNUaEtz4sD+H/MGKkogfu3dD35xIbgBm9QG30RASz6eQHY1bI74P4SJ8XhN
xV6y42jRXTaSFNDUUukrzhGVZQ6ulPIIuRjeMbZCmI9nx66x9CsprNs7trtV8upg
3Lts8Nmxi8Rqb2a3GLf+/wORN95IgOIOUNyrVlmvY7AGrIZizI9VoZov6boN9cvo
wrAjiH+C6zwAcWzA9nR+vcw8yu3dwVp+Mgi0EPkA9mcGnvG+JMYFvFqeBkTcFQnG
7vhrkG4cuGpVu1NOK76wW0VCwN1XJaficbFlp/r3tjKpk8Df3Vb4/nDFtaY22gy+
1Oh1InifvoA9RszNFmDfmT9qrm+gL1TVNq2ndXUvRxHmm5SvnruevFnlg/dQmkJh
niSGWa1NbY+of0n2NY52IsuGGnV1lYbYBW4ve2XV5w/RqRzqlyHxU2hlJG8b5x0o
ytkt0iwFgarWBgl/5u2yVJ4UXwAYlGRRLHlvw/R/6TyQJYcZ9Q2devdB6gqGMxtO
tMlDwiy60uBC/18Jwr9Sq4XhNnTIEkOGN6KGK673BlQhauS9g/PzFcsIfylUoIZy
cSHNm9sggiCiL590oXDf2a3fpibyMsDFzPV6v+/KhQOMjcIdpqplAdhvjuI4ZWc+
KuEB0t5mpAAmPU8QMzziD9E91ojMieY+5abPomXjq4muy7D8OD0Sau6teoDHPhgv
BEvufBqcXX3sYjc1MEETcFdz61raCp46WP/YjxHSiRhT1OPWBNwWnuySplRbsBlQ
Q70+eV7MYZggzJZCHP1bO1l6eiz77TsYG2X2bC5bSMkKzO5Eihe67akVm3cVqimI
n5KGVnaDnaF0R4HKFlNhYvKcRc2/9OGzWsu4qfJvY5vGLtxqsjpblWdg53ALGkH8
tSEe6mK8RtmISzNrN2pBH+gUE1U3+8t7BnLtaiQKaTINF5mwHc4s7EmSTK0zZ4IL
RigHHe53lkGgP0t/DBH328pHGeUsTXpzeb5Pl3i8fgQKkx6N+BAfIhaLdV6kI/xa
Yh0XRuvrb09FbLgX55apLsbaBj/8cS8FMZCo/dNrXjNA4KvU855CVdU725RVNscI
Jy+HHn8mlbqmgsoQ26DooIKGSEMW9gY7FjmYntuiHxybuBrh0oL3x3Za24SLyGdb
Ve2r/2SMAf8CsHLsOlWTuOjHHkFL03dZPz7yilWgRWk0PHtt4Y5woqB09C867StP
OtZJY+Azrlf4MEbCEtgbbJlbcpfSa3HNSqhc4vXvlKSrwA3rEk/1AecvLxhzrSmE
ar4a6vrE5XIbrQv0zL14s9ol55m5BAMRXkT2YVDNx0HWXrPrph8S9wTx84qr05u9
Xz/XMJoU9qap6CRzQNfSCuGFQFyAk8yOixmcMeUMIwmeR6CjtqpDlw6e4hxknjEH
9EhK1YorXncQjowmvBJbgSILWgSvk6OQE7PxgpEqUfLZVQVjXLTWGEHXl52EpuNk
ZisbMAEg1cmrpoQoiw60wj8Pw5I5j1cFGDHaj9CXhtVFUAGfmPcaLQm6q4P7ncCE
84CzKjt8//IwneJ+KjD1CqPzscpy4mr38ZdYoZM8rd+z7jakxK5Dz7OznrtNGP4n
zLURPgPiBWb3bU6SAmeKThhK68KvjdTw/hgXllbvO1kVHL4zLs8SxIcT8+/h8EX4
FAgc7jvGaYNUnGVh0YuyYtIX6lEivsuh7DNMjP4i+KpqvpixqDfSK8EiQDduWqag
QykbCF6wz2kOIKZUBbzc+FTeDtzn+TR+DcUVu90EHpR1piYEg1ZPShC6Gs6xDimr
1zJNFGNJ4t/w4HlRxmrvZ7eMRXAspTrfgQk5aMs/mHvpkCKEBs9s7K55nl8GTBwZ
IERYhU2m+rpTv951hhZLwhugQ1WnRgEkjwAtGli41UFuFQ2qREi8qNvPaqKTA7V4
yNTGB+y3o/yk0QtcbDkk1zLGVbbyG1GmbtnPUHMmm5QSKryrrLHSeZ1sxcdMsYeD
INCeORgkLp7OtXFPjCd2ZWBOvQ/hTjVZOrqXaY6d0IDMeqyodEW0rN6CF31WsdWb
qHdCrUo8QsMuDuK226dWipVCImoTZJjzRFcu2DZIGyRWDTm71HgcpfWOyUev0xTy
IWplS2+X69aw9BIuJL2yArnIq9Q9atMXErTN45YxhoIG3ODDad4J/wRxhge31/JB
c711LcMt6Y2yai6sKZb49nSeCDuhaQYYTufoHbdkhlSWW6kD0ihBoXBtGlyyEF7D
w6hc0GsfDv2JTvnCzN71iWeRZGyjkFcQ+qd6Ovu5ZS0/OCqBTdTRgzAk9qSSsu/M
rB5m54CiQ6YhebFlqBgnbki6slSRdIpbywGhce3XD5eLxnOYZfBHBj3CuVHDBRVa
IZmG4ydvn1L8M9LiGBVomZl8oN3MsOm7rfszAOKdS0l/GzZ/AXotgzCynKVSlqKe
fwjMBqFUWPcHJrQEmViKYsEYh3uRARQolFgwdjlDkusNzkmIYJGu+W5EWW5HiugZ
QiWGv/b1mHak40msb/I+8pE8OO7U9EvTfmlQy0CXu7kOQi6gkVjCaiWJxGbtW5SM
gPrCXtsxyrX8Zpop/MwmMl+ejq5pELY4fpG/K5w0crs2lGhdz7nyoSgwVj9/Ja5C
q86t+QI5zIImzFwi7Vp6DVXjPzRJ7YOZVbqkyFXGYFD4ednes4+KThRIfqZiatCn
tChYkSIa9BGCvuZOFh6zypm7CmJJCD1mhWfQ64hQWuW1Q6qMy0a76GAXltQccwA0
BB1dVRI7UySAyNNfMLP99Fc/3FDSJK/lB6w71PMLRVWnxie3NtRCr9Sge8VDI6Y2
v9QO5gxR/g1jy6JXCRnEjpb1ht/D335DvBk7Lwx6oQ84I+/Kvlgwp61qxFfHhtIQ
G3n7XpBn0hCL/yCtJMHSJ84g8kdcYLCb/cngoMmRnrBnNF9hsH9P1P3g/K/Ry+B/
hg5Jl43x1QIP4IQCZBpsJW8iRcVk6HEQF1JuQgmSNCXn83ApoKdLWaRgX3PFBV43
heIBeNGFP2Qx6mRva4G4j0bQKaJUFqaDJkaNPwJz5CGPgJq8VzWXmA1IZWWO2xkK
pPk3OM58dux+eVzpdw1dO1vmItrHcdnTJ7/PbV/qRKkXoPg358D4S8iLx3RJzhiN
NpCE20t9wi6A/ExSO9EKqkhtmFsWqHBni8kcSFx6vb8xGVXu08JKzJhrJOIv8Y5M
X1OgBaD80ypPGfWQc0lqbEHbgDL7NpPo/00rgKB1+ktHVnoeHrbrNlAmLmzU70ks
Y2tS7ZaQuhk3zfkf4goMUhc5DkDiNgrxxf1wX+MW2T7l0PF1Lpmag7Yp8yP3KBE/
B449iq5yo7KnCQ2vYd4jJtH3y5Z4W5m0Z//hGtNB4qYSeaF+BXMyPsAxeSW9Ev2p
NL4QkRJ6GoItDj3SjignUj7fXn0PPfN4lyBd8I3CeZyxa57cwvJNlJljRQJcOoyC
6AnevZFE590WGIJNRK0CwvBPdXzSbDMW8vFkCEnW9Kkz+YKq2vsiPRDvNbxe5vIv
VFzv9qiwz3XZ3ZSkA6k5dKJoJG+xO2mzjoZCBaaTqAjOVmTitU9Zi5Z5WF2l81La
1Vr+ojIwgKX3ROkJ2u8ohmgFq9Uol1y3TIGM01FNj6kzrwzeqoCaO7ktzAgn++iH
7jhluy+lACfTKUXZod+sogTaun6vWVfEzI01NU3CSe5uZ7BUrzMs7nl0qPHoBEQp
uBb4Rx9Ews2+NZzTdTUYbcnQeeTGi3ax7HmUYXnYsRmxQFvseWo8o1BtCj8D7dp4
I2ALAnNVVNIfSUs3a36M4sFA6iriOgGHvDxvH5uPHV5S6jvWKYJMB34loadxOLgB
+/ssM0DG9frfugjGbjOnEGWF/pDarvMihC2AJpvhf0pQ1Rqf89HRW+vGdungMXBx
XaS93uiJTX0xWfLDsdCI5x/nUn55jwhPLRf1c8LLKYSaRzhqLebTicaG1xauo0ey
0DQ63ZWeAvjEGQQo9zZF3CcxnS/U8W5VteLNbgYRBoELThGj9W6/4AOXYUSiyKh9
i8qDdtNPea+ZOQ4L2duw6WwD14ikcXmIuJYFEjdvMAmcN1ul6UTngNn6ELnEPQlJ
g/GOYdS1vzaPljoEOCQsFjfAMHL1EemcytL0DzhISsZO5QPCc/yjDysugVidMNZ7
wHoSaVDgpbiQmyYpqypswTC32nt6snZBAs/9D2CiQ8vYlkQC8hCn4WKJeXaX3ywe
DB6aAY4PPhcefaqjUtJe5Y47UtJtaGIAYDW12UHU8PCnc80e4EPhKijQaWZJgKOr
I/wP5kUu0cvc4NFZjW38xJrtQPv0/tscwbouhS5VW2O//O+VtQczd7JDQeeHLLYg
e2GfSrx8uQr1EDQOOD0b+zkJqx+JqSy7KREVF/RGIiGo8l4f52djgPj/W0wFScQF
LyY9xGc6ElY3N89fyjMeHNWzYkOAcQEeSb2CwTPB0x78BRiSRSkxdID5giLBbbtX
5wQYUzDSx7aDvG0jxe/xTF4CjZygES3VQRAljDHfj8kzhwUuF/3uGZNsmo1dtKzN
YjoHWeCpijaSCbn5WZ+1GxG5ZpmAtDadzuA0/i9RbELh+o9qUsJFJqMyG8j1JSFJ
1iiafrN1wzMPP3M9KWmyHZbAN+koy3gd7wmlCJirI+zumt+FBZT2RfwdjKkDs2Cw
Rjz3B1pMdjQebNCW/1ojKMMeiJzzO4c/g2wpVdMxRey0/vTIP3ar+7awUV3HksFM
4ooeq/jNK4Ceqag9fGTYZIElqkYRiVh2vm98o8Ol/NMogoEKCkqpu2dnTK5Z/nZj
FRSNXphfB8uI2fMzUL71+L17G4/LoGH3Aaz0U2KCMjkbYFr2MXIC6Nk3VOTt3cmg
Y83M7Z/ZnqHjrzZ2Sh1089RqVJZvse2QyRoxVTK+D6g/lXmpjrMTwd0BI/koPqKH
KP0EV5hPkfTY5s+4I+YCvJPPdzUyn0y7ukFcm8MO30ynGYKYB4NsEyRHNIZxT9Uq
B2Ql+zm8AVYlc1WO6cH00s5Htn9wcTbgQ0k9cqOf3A9cqHYuthHDUGL3FiOQX6wT
lM64hFUDphapsCb83DUiE9SYu+E2R9dWQeCfBuW2DX9tczBBMWrJYYmLTWHd46HJ
G2yUr8wV9ghSv/MvBxNCiNG5sCCaDHBlJwkdTLE525iRaFJLlG8UD9DyTWRudmA3
QTwX7B0C2MNpPi2LMG3o8gqb9o6s5K7nHeoK8i/tpU55GgquH7mhI8Jr+iElPpte
iuEJ1DXfwanIUHWl/lX1blNc1f6d30+tqXHBSnXwVRTwISAlYMvLR/mmDdAG9DU/
1OcYErV9/yFWseEkoZR5E45jMhEOYZCen5ve88m3wM3qYdVNrZmgv+xAXDPj/a0+
l5SbwWqOEZu+DJ3AF6WQZ98yG55kTk1zCP/kmZ7DgM7vt5k1PytRDgxcVZo0biGa
HfIlRSipiYLxs4YSF9BfhQPfmcdYY/B4qJdDoA3DXNPoRbJrs8nHex2MQJ8Wyvnc
j/XHAjuYDWunAYrpIFqdYaq0Q7sGJ743JGyEjFRTjTdGlwB6vtX9pX23MKheHDgm
OcWazFZmlafKiQo6Ao/2Fq3UTnTHP0aXxHo10YCAgDV5BY1SYWuReGnOY+2D8REK
R+GZA0y66WxA+Y++95oAafP1rXm1RrvSz+7uLuKwf/glnRt9WG32IbX7V0zFqRhB
wGwah6xR7BOwloWsh39485PhGf4vUjRiDi85JE4L7QvHZRKix7Ih6io6B3V8rQje
UHxg5uUzmEwomdQEq3BeA01Xm4v3G+iDoHbXhWJmXqGWXbzI/1SNsau6FCzA8r1E
0Tqyv1606yU8/2uShBwF+7ufFM22lnTiTo2J+AhaABIro+y7awZ+M7rZ4OkNsYWp
eAfIBBJcl9AGcn70Z+xbadSorwdONZ3BwjGNuxjHmRFWslMMtPp9hAI59LSi+78v
SxyGj+Nin6a2Aqv6MOD3gL4p+wI7Lz3zk0uaclfqiO/lDAw/sDPmWgEBrKEctjSI
Q9VFKykUzO7H/AicL0C9Hz9MpzBMWWMnTZA/lzhNQNSB1r3Ny8gaDLx2WIPi7q23
ETgEAiXWK/Ik2RoczwUpyXT7yqoDXaPDrdRroxYpb3S1Duo96fne6d8AWNjG/ZwK
6matO+jAYRUO7CsJtrgCCsL47ZPn9SsoHeWwhxo9slneFJyzoDuJ5pVEB+j0URSv
CYVaUaeLiwEW3f6/oDsyLqH+nTY6cuqONk+OuFM4fPnVE21pl8q4yEe91an4fdpN
NM2woV6tyf83Ye/Bu3i4v95AFpynLZjyqqBCCbWC7pQqzYFRT8xiKDyuDBf2p47m
JdcYghbLTK1gcl+Zh59TTjqnI6pEyiaeRJatrjf5f0rW+idHmeVXSWQtIfdHAT9r
RkTvOFXoId4PJgL/shnMwUCLjcrHTexnl7HxBxzYPTBpBKRMdgkkGMEQni82XMF7
I8aINy6YDFpJ/r5w+v7BUKZ7uk/IHTTHfIE0XABixW/3A8K60wJK+AhvU5qt8Kmh
hOLs7ci72oxU3KzrnLBdUp1ruL9WsxSR8mdlm/nWDxFaog9oLMpfRZaeWRfPB5g7
11aOe8lrt3CFAjs8IpEkZQUwHc+34QBXzbgmQ5BGjhZ5njnbHa1CxHhTVPckrtVQ
LCdqmx+ldNYRHn7y+FkwY4Wdy0cVLe5zR61+7wFm6P5i2WDLJXyLxTckMl/+yVjh
nWJNFdk2AJn4yro5tMjfmK1mWDwFek9BoAgcGvG54tYnXvJWgCG+36cnxbtVmu/L
SquFamGzsdQ0/WcxVQZ1R+gCjF70HqXVsMAmNjjqKz+Y+hessSvJYUxEtdi6ckeU
/bM6sT4FKbsEJCnlcgd2ZsVq/gG/uWoohKy/+o1yMh/bKqxJuKiFt0SDhWlRey0k
jDij2QlUCr9GyTJDFZWkYbdQmRPzEd84X8EKEa6S/y0/OUwrnl+QvDZ6n28S0HyB
J3hebHGEb9osIkGwS0xTTxhNQG9IyswC9ijsMbcNKqpMAM/ZUOAKxFPAUh+4iyb4
ilBbnwxdtAYBN9njuxMl9dBkXt0ST0fOzbwVslKLKp3sHbq/UlZUBz3SJVhxsvu4
7hSgEivKDqKrzKfQYzuJXknzmx5jUi7PHvCTK1uWIV0wKtdAC/TaHqjeNms72shR
76cWSE5wxa3udv/SJoLin7aPl8fhI08wSivVjewMIxp0wXAartQb3ABwQQBeM1WS
CZsH0dBnuSteWJjIjAKCKNb15de9Fd7dHIWCIeC4lhcWGnrzEg5R5Qh5IUiQf2Sq
5+t48vCZzs9wpE2HLtDqFViwlUBLZOl3TQg9aIjK7AUL9cQ1bPUs6J4E8SXINSs2
qrBSXeqVHu5ojXIY/tTl5qqDoB5CStzt/kuObvEMYkr7KvaDHwv1ttwzNmBlM7s/
X5Gl0qeZk8QMhTSqNJQeyl/SWQLE9If5cD4oufzkNA9ripVnJH6DrR3x4qeP8p1R
jpqGRMuTJbeSH4cqlPFHmR99KqsteiKTGimuSmafjkgzPSdafcpcCqzPzDJLGwp+
KQMLeWzSnj3SE4v/n9BuLF4u5yPUqdJX0gDzPisZDq/kIa34w8fPiSqhUpQOFOTX
0ULpFiOyUrDGSOiRIbUdHbbpKgE379MUj+BzDV4F+9LcItfwXzruaZ1VDlNcmWnN
I3hBvKkT0boFdHEXI4KW97H/a1F6KQXy9kdvIVGgxSqE7w/LEEzP/5TqUqL0Kaj2
+UUmXSMd87vMhoNRl0V28GTEz0eqqI2PQbCtA9fZDpHJKR6NMtkbqrhBPAndXGps
Z7l31fqz9pj+4bJ2AROeRenwFF2wlLSL9X03gPPsHq3gQwedH4sA167nMWvs9D7T
LL9SZiabE+ni8XdaW0+Mq/wewXjdLOlJrz/6S6MQsFkWYU1So4CK6qYLhY+EfWCK
9iOK8TlBz+RkYBV+TMnsgvWpSQ0bX1ozc1/Sy96TKjbm4is69vh3H3H1BWfytPOW
WzSrv4eBusfGCJy+i50wM9tv0a9sJszMAFGVwbmR9OLuQAHhDm1IroUV+U2dyWnR
LonrSwwhwFy+vxrCK3VtJjal0kIKR5SL6oUs+p52cf0EZMYacsdYIDl5hUTM6b74
CQqz25hYEpbaRhIVk2yK2SkcCLSYSsvlohjtxRIw26oqbQd30UUbxRBFRXnfL+Bz
OB7Ftaq8lnxXJxF2uJaghouPsfYWu9AMAfi2ixEahzHGiAZMnbgqzETMlIqfzBpb
cQRxnwhsYVelBRjDE72qLgFoDs1yVMIKj0zGLGJb9cjBxY7lxAFRCenYrom1+Cf0
dYnsCDs074FNixc0mcdG9hbjdPi82RlE/wADVK8okf/+MwDXDONRwP2x3J0DU+n/
eYIJO0lIxx8XBKSQe9H7pe/r8tJAXwf1XoZTeDpvIsnGuIKw/Gh1cNIITOTwAHCc
X7RHwzvaY1mVNVcrcaro7ljbQRvJZZjpAxX6yRM0bt5WfTB3inSkTrIV9lbAwHb8
l9BYlnwUA7HEsTPuymOONcqdRMf/v55xA6K8mDSJfQ97I+9lmi2AB2/JxVXUV4Ek
0IXJQvD+ofTTL03CRmCLP480Vn0qRaLR6CokNDyK45MiUIuRd5i0G8s1bbdFz14w
hRYfLVi7IH65oZpdpULZjqsUjIe4+49wBommZ5lujMSSBYoXITE4nW7lHo3+4r4q
ImbSSFPmphoxs3nMnk282ex9kCa1mdLircg/dxyl9yHNexmQ1r0tc13+Vjbxj9Gg
EVata6njQhTnT6vNAL4au/Ce3ny+CwOIpp/okrexb7+skD05ywX3cGGwZjks4vYq
D/3fF5Bn1sK6WPGKv3NMCIF50GotR+HSYmQIN+TXygA50pecfCB7cBq6INZAZ1iF
mTfQZx4PhiXgiElOqEDnWsvMf9w3qDP4n6bncVIUWsPDh74S3e5P6zdlqSlZEYL/
ik3lRU2x/DcrZ9UVSdv/5BqxQAfn2GedZtlgtClt87D8Abm3Nfc7adz70Hl8kFX/
DZu+TPI5inGa5MhC1/7KsIgw1uV/RYa0fRTrO7OKJQdbhraPtrAI6MhCCEZ9RbFy
gZ4SpIDB8Wh6HbgDTaYP1bd5oIAOqSR3cKlEQ069jEDxvDsOUD9z8ac0SWa3NmW/
t9Vg+RwpNenYEQ+Sm0gJ+Gj+IxRR/iWeKdyrW/7EBDsSWZAr2x80gWTwhtRIFzRd
8WY4P9gUVpx84HBDE22x0L8JsSQgsB/EH/FCkFo7Lk/TU6GM1ldDj5UWtbMAUeHc
jMMdmeGGhiiY5WOi+yAD4tKI9GmaeQyApfInyRIdC5UZt8ArTYndy/2Wcgs68Q2M
qWrcvsefhicFwNOhuYzR0tI09w9DRRERRHcnuhkqT+h+amFh3ABjnEBGxM+LBSvb
BOsSeu5tJTZ0WeruiiiszFkYXK47nRCS0huPqZmrlFCCMpiDZmE/VmzywmZTZcXX
4dJykldG6IL9dVj+JSwK/TlcgLvywoy1vTi2bjU/JruvaRpC1I6akerbGTk8FHg+
bgJniaY4IT8g2Td9/uzb31TZIMi86X26lhQEZAfubYBFfgABW9flNAQaAMHzsFsz
rfqLEC3q8U75S1cYBK0logYMPuM334sJXJlNLKXp2dSmR8v2njEzHdq+wj0V0s5M
f7EzBOkKkipYJjG3L3mPH2/CZyuO/jvbmgh9q8o4AdxrQhbLr79JEYJXtB8VegMM
CL+UZgx1SyGWjIEIE0XIC+N+o/tc0GdWPXnks0CDGWssKlkEru0t85fPKcukIGgg
axzBz+Y56TwVCvI7BYsglnyCgstVEVZ9B4oFX6QdP3X19Aetyxw6QsAifr0gihdX
Pv7wUwBda9StYs6uA1znNBv/0D4DMI1V6Sv1QYrz2FzIqsdqeQ8o8IahmgMzoyOp
yfFBtJwGaD+gJV+F6Y9T4d5GWgj3XWx5kLbBwr0oiDmhAPVmW+nb3BmRbpDINB4z
cgVSzaFbM4l3phdfMa3ZeWyNDSCGBb0/SY9ADYICB8nGum4eTf8e30HYMCmDuICi
loa1U/1KU94005bYQzgYUjYH8gPzARHMT24KW78T8g9lRq0KbkJHVdL5G9amVVQ5
/OVFyyCLfg5psItxetHirQxRlWJqhMFFW1ZXPVTgjEKR6uK39gpwoW7VCRZDAl4C
fv0NmM3wPy50BUHglQuOyYxDzYl9KuCDPCqGRHi7wQUF8SFm5yZ6h0molMlbJ5c4
paPYdFhFtPLbF2LrKFyhdgTUhIX4/Wksk9H9PJCVbgDrXdjRzIFXAEhJQwPZ+RyW
Q0QkuX12mpuK5n+gQqKhNrTtulqMlWbA8K5W6c63Moj14Kqi98jTOoGJ4npfnMIo
eLQOIimX6PIpHsLHTU6hMFt/AdXSfcAK9SYgcNsVzDWFiAY5kXGrEzB/89xbohyT
wG/rVVENoGeJStrMSLZ1vIo/ElgYYVHOKgxjOswnpUONm6l2xnLiQn8h8veDx8Us
xqwSJ0zpAZxwiSDPOduXfUWkgkpZK+poffaMDy87VwlBZVL+9RLv6Jl8yuujfjB4
md2KbaxwZizXnKF5TKn95ed2+Q5h6p9xO0ryzVFAXdc1Weu3WhdlGIrnbhzQMCNY
DST4J42sfsgkBJQCQUFdw2lULczj0TsKK9pKF3zf/JK8Pmk0iQF5IU9S0egf3rQt
QGznV6L3vIqMUtC4VYaeaFYcA0hd9RIYtTzv3fv3QQRnlZ9ETCrE4NEGBpZ6Dn1/
QvMiupr1NOg2QtioeIZcTAbisDTcwcke6WxYVVoxgLCh71Gi/EO8opJoEbFFcxGb
Nts9vNNX5gd85CZK/RI+YjHnrGDYW/LBNrz02X58TgjQAutNyYF5A5Y4Mrr+FgOO
2JQYW1PHFkDY1SjV1neset/te47uKZ7MwR90FQ9tZNDAxOlKNw76eG+oBmppAs1o
icXb8W0YsE0rdkoPlWy2bJeQKEa8l+viv+8tAnnLj1G1C7sVMJlmSxENm2X88Qs9
HLXE1bv5l4OB2R4IJzr/hAC3O548SnhSOi4uPpR3TgHEoUn2WZIhLzb62TSHvOMH
yE9EvQfQiOylsQfZgTV3MJc4zDHpeXES1Z/mbOGlaacLmLAivPASb/E2zb+I5k4I
aslAqDYGWWFKcW2IooldjHqDx04T0o/SrbhsbPkNs/jBjDR9S7rN+0L03qempZ7o
/WsC80MRkzu/EQ9F8qKiPTzDnvhse7yT/lNveVBa9sdJirqDghzMB+ZX+jpBxpdq
Bcp5Er+FxfuY2gwDtTpBagtyZ4+2jHKE7T7Sj4+EdSpbCnqCV7iTZLhKOXl3shcz
Sj+SHlENPOFUCmgKn0HsgcO6kKR7uncbx3jtdvGgOKdlw9HvVWAKSksqcbzyFyg5
winaa8oWRDArBt6kuBEkI7fIpn22ro0zR1mKbTN6Nfmip/HLe5yEbV+213XAP7mF
f6m7uR07AYLog+EcTxqatzvyPO4KjBNiB2HjpnyC0NCNkTzJll5jgdvlk5SI8/5Z
4GOuIfU1tkwvkvMJo16xgTkzcMxrdPwJn9oBl51WK8EiunWN9js66n8NVNJ94L/a
6bvicV19tTDBvlj/IQaR5Hrd/eqG5jnu9sSiUN6ia/RKIOP0Q7M2WC7msN9OX2kB
Kb/02qC2zCSoYtirhM2PtCv8F9REESJOnatZvvwncmFk2iUQDsdQYPZ4te0qHQKI
d8eBFrNjOamJuwZErBmbkNwg+zd8P165OsA7q1x4tejPpSD5KBfy2jN5zSlGCxEW
XonrkEtaf6kilw+RF0y7QgSKYAjBI0RqwiWFIAwZ/+r1cxQjAFICWJnEXZv0F7VS
lw/S+lRJrN8HlJ8ToACdx5mJUoUj633eYWwiBThV9sykLWx7xDZgNLjP7IzJUAE5
2Ly+gqTkitE6fBSdJyycWBEbf4R6HO3lDrMe/8q0raTYSzdzgZbUkqmbIahkd4Gt
58oGiSeowB8AKCdIvPw2EP5s15GYhWnUTT8hCeT4Y+hjj1NaPaAlZaTO5uW35T3u
Hv0IIm47c9LMfM8LoflKRJsTG+6yby9MzHgaCjTJSjs7+YSAiA6HgvAYgl9rsu/k
ubpQYx8c9nCr2Ixun3qVd30pAQpjl/d+8PyG8ctU87lqglWU1Z/qVFSrttnT7cfY
ONWlCH9ZGAmcD5KniMP5l4cTsTvvh0QNEI64bNNjMg/7bFzoAWSThbGwpSxtbtPX
Oe9ylMRsL49zYhimIatihBZAQW0MCfMm3IAjIjw1iTV5AbRJKmdjrjD6pnNm/PLA
3OOBjkX8C7clWHgxxh8xpDe5P7IEv3pdc46FsIuSlxAPstmxcQmm5QjpKVR6UO7j
dndSt9iD0d+NHW3KnPMYut+pbTc5z8llY73JAL4/7rF4mX5dhDs+bi6vbwVWSuBF
WZ6m9N7jN+CjEKMxCv/yVGJX3OhYLpSZPxEaU+F4iQCOfssSQkJAtxB/ZIy8sRnE
OIGbC2RjYTgiSwvcAwr2Ei992L+uRtkPKmUaVms4d0O/bSTH5QGhBke1FWFZni5D
Uy3z8tg20HWcFHA0S1wWm151JfTnpvsi+7UjPB6z9CYCK8q5/EnCU5uliMbCQzhn
QUN1N1cwuuj/dggfwQJvwOQMUbRQyfnpPoMqUFm85E9O0UmT/ngPPacqmzVTNYVP
FbnrIEvtD6cs6bZDa/AYQ/RDZG0bjC5TmkLG9LJuIY8fC0wOnqVRecBUQjQmp6cD
qfwKAuk/teVJAOJ1vWeMx3ylnXNQ+xwFnH+64pQItJeTCWDlsm8awKhFAvF8hO6y
wCRfQnkNdddVGtw1n79V9l6r8WDC4ZXg87qfjC12fx1va4W9XmxqrbScizw9oHpJ
wrrcD04BMF+GObU3GBgLvUvO7R+Cl9MQ6N23L0r4sGXp3oXzMkv5n6UFHYindVYo
EYnIksueff/Gv8o4VjZokG80tmPF6LSaXitsI7n/OAc9EoVJZrcxeL2NJrG7fSAY
HFWhQSJJr80rF1jFpqocFL49rWbYnW4kK0IbHICb0ne1Du5ucVH6/qWy//Cr0/IZ
R3c/jssjwqOuAN7BBMeOjTijrEuBCgfTR54wnT4VOp9Of6gDD9EkFoukQqmfhWmZ
/5pH+vOTiyl8gQi3o6Pm7HB/0Q7YCnA67/IZRUtVfHQ049i5ix4tHkpmSFAJSKP5
SjGz2oiK5/nLZaec/CNFCkhQZG0SXQbWJ9P4FigNVSBR6rrEYpkD+txuFptWYQA5
BWxmJaODEzqcAuEBdf5oWDUO69TZE2mzKUWOW/aq6pdYLsT5PN+bDyhdaSMQfpDw
ABESZvCybZKTq8smh3XOLl6coF1q9AwAMPfYTFHta+x8LAT5JMQcO6TSoz6iy0Wv
PVTmFa08B3FHStDPyijcL/5/05wvHmXZw0r/POQX/Gi94PFnXRMBtQESxXVyYie3
/O87IX1DL5YwcNrykqed8J4Fiz2Wk1ANiIdUvfGUrvEeCBUvG5eq/sXz838uwbCs
vAqq4AVgaXZWGG3THV8Ux9zzIPAbd5fWQHJBKFKLSMRxHYun2vhu9V6gF5WROXiY
b/qdXgjnqRUSzJQnEoi2aCKMOKNam7eZDzpLuZZtszqt34p9pDeEVTL1McW/8dUU
PRoNT52LGPz17ZS8car9VIw6JWXbob/WNrE3K3PSOlSWuqDXZvd84ZSB+pxqZOF6
I0jMpifpvFcxT6Ko0rf5OmI8NqRa1xz75kOrzwcXpZBOVE43cixKPqloEI2/Dw8B
jVnLNgcoAG4YshfZ3s8P0JdoqkvtNv7Yatl+vyrKAtMHMdR+phXlCqIHPr1wTTU0
1u0hhrOpLhUyOtxnFsepI0swquYs8PyxqOJGCanhTwzMkGSJwGTlwyik7C0xU5gv
0MxiNXJ9eP1dZo+ak9Di3Y8ImGjMwjCcEx9K6L8vNu/IUX8aMM0MhjFwFd8wMi0b
nFrbtWcbsfPAHTADvowrodEtUxB6U1Ij5F5DOKEQRu2rsPZY3b3Xt9V6pupJspOD
g8o+rvN4qoJbXO9JPVs67gLNJGOPfK7jCIp8iHXX8InwkLZOhlaAGT5mkr061+Uj
V0FZKHpN2P5yaIjZ3cn+AqgBdf3UKaeRCzwB4s7HVgvHRs5hd7Av8OQHMc8luUbW
Gpf+++Wuvy6h9gRt+NCdK+WjT+CxUMVlSZuUk48i+5Qpjjp1AZYgezY9XzfZnZyo
dpZrO7md0qUKawjxDTWpbRzzgqPp2QEeTKKzgEFk57bgZi/r1uvz7oHvu4W/LwMY
XQq7QDnmstO+TLIt9OWiTq2Qvf5Rg2KWM00R0QMN2svpglzp5icNfQFdzFUMFc2P
lNXbVDEjzZ+kmw3xYr7Wug1FndpQ5CSdLfEUx/dUxqvTry4bMAxkwZgSmxl5lE7b
RdSOu6UO1RSfJNNfY4j5Mo93Tu3qi4mQw/Of/rE9n0c4A7Tfn216NBi8UlVDy8q8
tdNO8C9576S2SYpSjwwe3GHpDHl8PoZ2ZNuJoUeC33vLDAJrMDxyxAKOS8TQvGlW
y7Buh2OBbOKlpzPGqAmjKBwcQ7Fgqwr11imqd2wObi73mWwtWLGuNxXkJ/GeLQul
KnSmqAMg1QQb7juUBfW9d1IfuHEpKNTuCUIPaPu6ckjlP6nW3aQ0EKgy/6q7xAgB
tkiA8vFw3uJ2IefAvDKrCWrcmZknFHsraAu2KZpiDXS6Dunmtn4qzgre+rF7qM7P
gNefZJo+SH66Jy1+yG/AnrvaN8IDutpcIgsj6D9BAdxWPgtl9RO6PyeE46Ctl/jA
pj6jI967wbwl2XMn/MPVVwNVhOvLAFI9DpC3hvXD/hqTqakuU7A0Z+daH274p5bO
2JFZwFAJaFpvzotFzMEBEU0Br8FPajVXzxcposkiYZX4mYOZOyvv26iZdUlRrqrJ
xQ9Z7o/fAAs+oX1iL4NZkfzHHuJKbn0ETLD9l8iegBepHq03JIVKE3SftUH1dAGy
3m3p+vcWvvSA7PZhcroM3BsvjIS7CqMq0k3REBLXq8tiKmRKCmOV3Yl993Bja6q+
PgBLwdUZauHEeRtkuyp65I5uxzlw+yNmY8tJXxYTE1Wq7o+3mB7uM5HpyVSdwrqu
2X/rpubtLO8nTbarXCKezgISZKsC9gVU2db+heyP8yAMtHrROHkJanysFfMO3Z5X
OLq15Qk23Y8dcOOUmzlVM7cJCOZIIZzlx8fvrdlbvH4bNnB95j5G+t627/TV2/ws
BeMbMD58LCBiG3hOxdWqop97nxW70ZuMu0ngD8rfrt4dfVvaoKirs/QZyy+ihiyf
AGvqVf5YJD76iyb3mjux2OlWxt9Zs3MJhwJDde7HH/VWNzWQeCkGKV+dA6xum/kK
ie4B+WSn9hFEtRMr8ydBz4OKxpNyJI3njXQOencNC83GiNQi3kjnHi9NGDTeiivp
z6YL6e+MUAMv86O8bjoApCPezaBabH7QT/9zdKJ5mWCw0B+Tl6wXFUfhwMyNbFN0
s9LEXbcThQLF8SZ5bKf+rS8p6utkW/CPS6kpJ65BF3RZJIR203vTHx3MWRKNxLxh
Vp7fKxj/YqH7RbkEyUvf8PUhOUpGXfGPHOexhLU8qDGM5gSWPD7qHW6vYsdA7Asj
fivxaSP7LYrH7NUnnmML2nHCAR29/z8xwCtSVaIV+TW3JDLaGWTbvrQ9eGR1bk4j
Hj+gBjYAu/0ZSdLAABv/LazGBS3QPce4LFhfWJTcRrVioqc09jtuYbXK+QpcXwoo
MQz83604qT5nKfvhv8f0ag4TEKBKpRBz18cgWPC/evtS2S62teQ1J6KY5We6+fJd
omx6KwZVz6JYuY1s9SyoQS97zJbeAFMlV2TEDrBS3ERF3xbP0XiUJx4pYNnEnJoJ
GKA3HoHDet1Ls5h+PhbMCSbnjhnq6IFaLkIGlX4AgNkbEWRsLqXH3ui1TYf+koEz
P/akDKlZg1jFwc1vqybpa3oiUlBhESKfVT+4gAT3Bq+A0BGZbcO+DZL0bJGEueHF
R8pZL9W28ql2rqyMuQpwFAUtgX+Xr3h6Omn9Gsfd/cRo5rHpkGPwSroJIpspAO5V
4pIk9AcxzpkoCI+YF1VaYEFNWc8ZEP03KoeLRg3x7UHjjT5a1lHIGDeCWrtlSyLG
YAJBLoiq7dpGZpTSZ+uqQbfr+Z5wAGb+EhdL3qSJZ9CnOVFa/k9sSC1SErSjBM7g
qY0KCFmhLzVXn2zyJIc7ViE3wqNwM0ZmV7rqwZep9qrOJU5Rkrup1OJVSN+47+xH
UoOzHs+h0PwXauZJI83RWxh2v575PTHvSfAfvDedMNDdtW0cXl7rf3jys63N7vjp
4TwWS+lPOdUFoGXnJ22Bzh3OYVUQcZDCf223A9LNH8FQw1wWv56x4j1UtWM78hfS
jBARz42iM+jIn+QsYdN/qsaMJvvXXBCAIy4/T42bw1xou0n5/SYNwKyEa83tYpmv
YwXdTZvxVFgLFz+HUATvbg7r9grTvYG2ZWqe2sEkT5DWGPzkEVGpUb3DC383k+Lu
5W+kfR0i2O3zNH5l+mehJfUAdQEwe2pbSd8D9jKuncksXKRo1Z/vC1lGJ3E8TGzI
oTA/b3e/9fTRgwVtaF3a1J+Ldny3X+eyEvmTaEPyvTQBah9b97rFQbvC0b+eeOUY
o3CbYJi24qifBsCnPow5RgS+BMmSr9Pb2PVGAXDvOmh+h8GlsWnpydzf44+6GhwD
U3vVo3VQcI+WNvOE4ULZ3lrK1t7G4h49ZbQnAI/VuBQ6lsQ/QOib1u8zOmMY8fHG
9FfxmDwRnSAMDcL9obTsmw0ddFtddNP9Iu3McTdkz3u0yMSHTAi72w6AJJGC0rq7
LOFzaYc9vFwJXJ0VUCO2qAicv16uJbmE3GRDxl3OYMCQn7VA1Ivp6JPPGIq8/j92
Fl4cZ5HwEaP6+ZvliCp585woNt7poE91p8/DwxNOyd/44CizwtrJJf6dONajR4A1
8GTrrvJ+E6iWI9VwMRw9PZW/14JxrrphMmDbX27O4UG0yIkUt4+rPcf/GBIL5WWj
G3/zvch3OLHWmWj/SeQx25YXYxT7CodhDEjdRj/IPv48PovD2Clhj9mZlhoCPFyU
+u1haWOgwnyYWuLpIYZkqmYSW2o0LhRsk3VIto/oBbkX10nFLYw0AeXgk531KHSj
XlyjhCXRbWyWKvMMmXnAfMdfWY5/nHV3fVwGU7tT8NhmgoF+333tmVKUW1MILosp
2GLVLqS6bQMFk4LcHPPd42aEV1ZhG4OB6tZRSjIZIylCv8ktwp9UN0+qD6Hi+aQu
gmuVrgU8rURIXZLGLgjZLOtsc/II8a+8Rd0CHCrt7hKSS7trF713k7VWlTu4dF88
krHvDce/41plvsf0KaKx9UdmvdzrcZH1AdbF6G92U3GR6oYSFWzrLiNMNqzeCf+W
7M3ogwMR0Nylzyoa06BGEWErhTy+PomK5YlGLEka1Quh6YQbyckQdjeJsZkcIFre
8kIRTDNcKhCZh0SgHntoNp7jnZk51UmMw/WKlmlDQ9ND3lqHx/ONKGkFbCSfTXn7
FZy7BO7PHL86cM9SZWZ10NPdZSIxqqRAvrBTPkG/B/XKNSUSIzVjMo5Ubi1SRJ/F
ROKhZ/KHIs2oYhG8ez/gQv1fqRy+D7HKe88scb4UL2Wkhfgf3amaUb7MvC5gJRn3
uDXVduXoberjcz4uDfre24jNvx0iEQ5N3t2pBb8MOSEJmBZeixA5OmgTQQh+lnZX
6WgL3ukjcOBcOyCt515y6v8C4TgK+S0j+4c646iKSPBvoZC31OexrIhjO0MvuHkT
5C3o7scaRdgdp9j/583AVOdVWaeIYIhe3qMNOE0J8HuIqbrJ+Q8WmGWyratpz95M
6xFW139pi0a9GN8JaHP2KUXe+qzqJEZCObzh2IhXgk/xBrndLqdLTGBbHQ6TFzZt
wVX8U/Dk7tHMsfQ9sBxNwkldjIgTCUwdrvvVT50TX8lHvH/5nxrxTcQP1hy6ai5/
ZlvgdSgfJeITrPYPFe7A1ctgL1fpe8ajsiO+T/rtPDMSV2bvZGrZHVcV5Fdt4R2S
pIGeIF4gJc9KqCsusi6CD+6r13nG+EE2ToIFkNOVRIjda/NlOljhFnh2Qu82nOv8
k54fck7VbsOhLnyBprIUapVRLjpIaZxfCWKtmD/gsYuiBDMDz+prPvC8hF1DN5Hc
FEPtz3GtwwLyiupUWsOGi/hApT1OtBVYcJfvs7oLGnhtI382h05TNQI23TXEr9wd
tGMRdo0mFIOQGilHO7/dldIavr6MsKxaP0oLyhKCaxF9r2js+Pyr4mla4A1+O611
wVSjDDuSuX9rLCIh7izbtYYfzuYP7RTKB3B9Db+PX4tbEaLPRAQDbG25J5cM9rkh
ZegKKH8V2eKpU+9pQpN0EHiN4YRj4SuAsdjzOQlq0hi/xcck1hQtn34x8d2aIzR4
8hsFyY+xY1lij+Bg6AiTBgVXOLHSvtacAChZBGTePyKwSnOP3f5WHoopy83xri4Q
UKmPE1ymNtB8NS28fb1QRZ79t1Alf5SdQF7t3IpYln+d71NDrH3eOvajwKO9Le6l
tvhtacNs1dJx68Pov4OGYGo6U8LIQgEOkj/hr4htqvVJ+wkMNLM3hFmgY848fszC
rGoGs7GpKMADU+6JXTMTN9r8K45AP27ojAnyPcV24OGexVrytoKAY194z0xr1R02
zcaG5GPGjDDksZP20ETcNAbPjUMNQBo6JnbLZcIIjnZo/SfAWO7RSxp9QECNv6Bb
szZz0VnvHeZd9o0CajdGoY4aesNLyaH1GWgM1P/5pcw+B0kUU5/dFi42SJy21JwH
ZNOVtQEZ2wNFJ2tsiUNl3kLW2BHhHJMXXhP2dIXMoaMhEBY6z2B7lAVyY0bWWMth
djBjSq+0dlnEQafSjtwlNrFqktSav00YOFvewAdMISby4Lq/dTk7AuYKXcLbgxv0
icMUUYmChc7kNKMkRcfhyjXE+0VJCUdh1IOLh9N7hc5vrEERr8tJujKhM2nl/Lyt
Ksvu2+sPHkRTwL+uiscAVVKc0b7DwrMxnrx7rHjrYq8xnRDTwlnehZGV5QO2FpOD
0iZAMCGI4EVAawlQre3nM/zfogaXHFprHR/ljFDIyAmYZVI01Xq8W02EtS177CWR
xd6wvWhc96zXzeHaMJHObDUiJ+DDG2QoQZa3qn8rE7zEcdI+zzlqlSuRjOrAd4g3
BCIe1lvEFIvYf+D1h+nqdkTk2sMp2NSvwLb1dLF94eUEkrdV9PjUjepWC++rrtWF
tgLTbF1fcdWQ1QRl6TgC1EUZAUx9Wc+M6Jfcf0XeFXyr+L9XDGKwhXoXdvq6QGXw
ZW//oAVHkKpORoddvCxUB5vHsDg+3YhZUi50xJbRDXTH/6pU4gBuodX/JeVRawUH
BRQDGY90Hgd7q11S5tNzy/sYGzWfDSf/5GuEixivMijNBNmoP9TmNbdxxlSS71Wd
dk/AE6fybHlI4jootfjaQ0SdWqYmfzVJgtst5cmMU2tBByB8vUjvOoSREV08mYdO
FJ6yaGWBcK3ppXZut/DsNHEPyA55HIJHnvTVHN1XackrsSeKM059/uoSArDqft4l
XyynOlCfR9DeNBQpFEJOFYSS/spqy8H5NntkBNyzAJ4bo9Hw6qc1zqZiWNTqQ/Ux
OHfsa7RYmdA8+Sm5SJUZLnb+JqoXIZdHOA8vzOvlYYGrpKPkU/oep9e/SntFAp2s
WT4TYurfsi2txuasn2dhpUtLavr/h+kbjIMDSARslMx03l3RknEZ/Pytrc7+hVYI
f/+pNC9ZAkY3hZFOADuI8HS9nHrifU4sUqf1XU84Kba0XFuDR2YnNqFnp4I8egk1
QpLm5+umDxsF60rRBqiD43IRD3HTZ25iR2jrIzVY6kX4Wwyw5f9LQdA8iAANV8w3
74YQEp/YLPnrZZuwSOOEtSXA8wquKJyzK/6OG2bOTtvnV6IxgFZ4aw0dILJPhnLE
rCZR8NKnST7irieXzTItV8H4M6TwCiDF2kK2Ru3F3XGw2nkAO2IbMvVaaQkaDfOF
IXUhLj/l/tO8Yq2LeQs0jWBz7CuzHiE7LJX+/tE8l131jdjJXHRTno8Gy3XQOPWF
3lDEyhYlfSsymeIHB8CwDLaXrXTR/5E7xhG0W2/Nko3xKH1KqgwihFehKqhSg7XV
4X3A/Q+qhXXoOnponvECI8bNg0nP5mlK/dR+4Aw3RFo+q8PV/rwaGGoKC2rZxiE6
Qx8YwlDOBF4Q5+HZz6rxTwVNnz8oHbdwhspq5kPQofti5E0Veia/4u0P7wXVmRYv
BnN953FVVAUAu8VFDIopP4uN1EwKsvLYp547zHXZzT1E/EYJVyLHKmwqd6FjYZwM
oGcS/RrUdfIgQSo5moUGsugD2W+AKkZP7WzzJU7rBFglKXgLzv6Q3TsZAdk+s5C8
61v5a6DBRgfqMy0KkxYx1RWa1m6ex0FmDXdfsvzs9ZVV47cjjO43hfe9oA9DgYsD
pD0S5py7GWvkFf8tgdwbCDmypTzEOtjuytwKW08WNuzbx2YymbDK3zQxcQ4JoGnr
bF718/0kkU++nQeSLt1TqRZTOnhx5feH8GGEr4SUE78l68u8A14Pwr7r5/DqMyLA
s5kLjcduvquLxR1EEY+BYY5GJO7gEYxsycNs8MSFgFZf+9LARGzvxvuP7Swm6MrW
feHpkVTJOExuo7Vvga4cBA1MymlAWKM30e9uN4phVZvD4Ln/Xcp0mFsMl8H6a9Kl
J5n2VluCAWz0y1lOQf0U9pLxcWH+bq6559Nl7R0/qICPnSLyy42Q2AZhJ4/l2MC2
oHq1WwpGB+/mzZXKZjILdskzGJs+9ggRPsnKRx1k4WsS+OyzLGsfmtdBq6Twqm1/
a68NLGYw1OzyYOJ9RA6lN1O4PFPkHcJzAjRhY4VAUKGRtFgkivcPSI7brGOqxwu7
xwnEW8oU1lVBRxzqahhszrBgI/FAL0llMfusOrFBqDW9hc82nzamM9NXddIw48sp
Pg1E/4k2sh8vvogtQtp6oegOJ4ZWEAdkPVSAKZvCm2GsTk9GaG2FNSBLjValHnuZ
FlSdyik9W5/a3qDWmvlPMjvPMnWi40O1u8Bo6grsq21lmw15Ip/Syco+aI+aJCwT
xe8Uq5a71b1xwFSKE8Hu/3Rp6gGp2g2ykpM1n7ZXWkK0kYcSHP97lnXa9v3aK3F5
ocQsoNyzJzzEg1HUw6Ccg1sD91YG1w+ePruaxX33ZLmQQujPiix3r9ehX7ItG/cR
QKBiPot/v3oRq6hrRx+MaDuJWODmkSL1T1MmyIe3hiOrREgizH0b8NlrI3A+UUvw
KzodyQNYgEj9tJD3G/CqMZy2Cn/pzgKNS/RYpFiKFfKneruW3llezYCwiJZg8c/G
FV8ytkrsHndND8UKJxwFCjniIT6dVxUtxpCKMGxMSZtDppMd+vb5oMeKgLFohlCM
vv+v96fw1P+YPXZsFLbiZ5cqHuZF7bal+uI/5skUrPgOdAGO2XbRBJz2WQfVkHR/
op2QG+yZCzg58uMxW8cApm/lPQPtu4wbg5WtlN73KZZcrup5L0raf/eqwXp0FwcT
834KOySwkTfjjKEuz2wmyBgM6Wtyt0roZXlhkSdlnlBknIxGbDSm6KtepnJm/eaJ
W7ouzGHJPBYEVV1uCsshtkmEVOa6KfWhH71qt1SriyeKKPyA2IAgxu+Ge+stDsvV
Frx+Dcq3M+aTFZsbJATWgtJiUK3XJGlVUZOm8ptJbWzkBXXRJCGFTznEmmz9KFKn
JOXzVsbnM7bmDW1XoJsuYUUaf4XZn0XSSBUHXvC74yhoz6a+8HUVenqY41bQ4M7y
yDqJGvJV1hbbm7i0vcoFAWfyd9ndOYiQLG+Rrke+fxHb/9l9eLKeqeuDpZh34wqM
9U3RIYf9YFnAi/yW5ccHiWgv7JiQq/b3WhUx/2R+ci2lq1DeYroBo2/If3L/inDg
H5M+KD6OJ3w+mRYOdjt9MDdVjmKYyvGBSFYo/v9sX87HL2ijwzPXPyI7ct4TSQ25
a0b0l/zccAYfZg0Q2AgNxvDdBN+5WTFEdFL2t751eC1HpjDu2D4flinjRGvNZX3P
pGnXqcDXstRbcRcYJPQ6FKBg3PUUE+KzdGdWO6BPpfjSBsNfQiu0dtb+PDIxm1VQ
Dkjo+Pdn95pyQPtUTs4kyQuvg7xQaGcsW57CcRdNlS3nE3PruNephUjy4nzecwUU
w5iEnXz/5dre8T0uNYRS4Dv5SNB5prmN73I2FJQsUmcjVm7HrtUhPbIIo0c0Hd3D
Sgf3PuhZXlQoyZCHuIXXAOcjGBbxmkrpVpirirlaArd7uTXvheJzEffzen3xTVjf
Kd8pVWhZMDLeqid5DR/DQZXNEyDHUSFlPPpCQF1zwfKW48fT16IC9c6Wp/Vvti/C
Tj1clfC4C8Np0Deubz96bJ5g6mtxGaSzVXhfd0OH9jsA0X9ffis7ujdBIaVsj72W
MEPvugBOEselg35oLlXsadSxiJLiJoB/omBbQosMOu1CbNV7bEovtaJC0xlzDvcS
Z8eOI0KZkODquu8sahkBfgFI/58r3OAr1g6OMOjE2dLlhtnIuvtVddMcAna92vC/
lT7a2AF+fZsySzOy3y9QfLE11lKRIRjbGb9uDS6gNB0BcTPkSMkNOBOWEz1eYc/N
IFN4uJ7LaUc+eAXV4rdFhGwhRIgw2qOnqrd3Fqb9vZDgizKUZfTshh9rfcaneftT
ivxvK2JfJd7Wu8/Wh3v6KJhX5INp8ZB9UpaGyIS3GS62HYRO5R5u65Odk14dP7Ru
GwB8vzpMhwtaAaeYmcjmgpXvkmFR1JqNXIUliJY0ZAUDU0w+pqpmJNrolpYsw3H8
LlkvXA5N4KJphLLhDAXDwGIYt248pxIUSMCkHlZCoK8rBRyspxZbC8PjAa68qYiw
R0Hkh0pI6Kx8QBpdLGgFICma8snQXcqCGk5qACTZjzdzE0aRM49tVj9NuvNiI8HM
JkgKb6NP6FT+EhA+7QoVNtLO73WOEaxIxD2JzBm/jkP0pGU0WmYjH6h0yI+0WyvB
6r8+tNVsuvkKtGcH+4j6rFjDK7aLMjb3lwBwEp8wbbskGsn3SL/BAWEdVIZTnXri
tQO1KH9+Oq/ARCOaXU0ywBnbKB7uXOu1NPOEHw2Clhvq7bSbGhTxU5cXNK198nMk
MUwivNUAX01qWl5yr29Ndve8pre/jEJlzN7cGhpJaQtU4DYHYtsnLHYU4yTNlB7u
XMRCOH+TbncAWauiUzzq4bP4JsC48wwiM4HCYZ36aRmUQwTzK9U+qIi/zbd0ZvYp
bnsk6PneOV4Lh1aTuHK1d0BbQlInFj86r7nj6C/FF1ydVr2ekSEotTP3ZMIhpbqK
aBG6WzPYffQAR4WOVNoRv1DODWTbfDwbPdwklZOWUlxW5B8cVY0JMs9U86LtokgX
iwCh0k6sk7MMhLHAjvzhTwK5X10SOHlb/U8pf0k3WUCdZXKSt9hFRLpboZ61Ikwh
Z55p1HT2rnUjDW/J2wjMCYvJtSCwooxXtTOEXgPO/wDfcTDxhAXlhy1+fA86YlgP
AQh9oChZNBCZTvYJ+hC4jY05/g3kH49WWVLZuwQP+np+5Qk0PWCX3L/x06241iaS
QSqR8P3dPAf1HTd3wB3NsKFQaSDlIHTfSBMlZb13CTLiqyyldsPuf+KAoKYVxz3n
g+1YTqLKRFb/PTPpe6HO8zVtEYjKKC0xle/DEGgOPcC0KElAnAeE9SaK0nREkmT6
8XGsFmk4WacJkWZR4Oo6p0ida1tkPDfRxDH0bAbkTW2yqMueBgNTfngej3/rgYok
tPNrXlo7SrFuv5zrkLkgvdpI9CwqZG5U9hBUYMi8/7oJCCwNozQWnefOZBrFoyed
PMHiu44sLjuO9JOIP0rwvQ9Pn1T6ATNsfffwSikMoPDBOFeWDSnXFteSz85lQIqE
zV5BIMjRj1QAuPBklEFH0fsCocbtM3ASz0oiXHsJ35h/H5dCMTtifrypXgzzWA9k
szqHpdWTpn/GvQOHv/67DkU+sx0Z3Xi9XanXYzNXcA+GD5AzbudHS0X600SaK8K/
Dj++RNkzOS5w2cm0R+fe7LMxSOq9Lzm8eQy3GwndUOBa5ZNbQXY6z3gf1Gz1ONAV
TS4QX2xdqS9rTPHUpIGrEGvpgCqzcHlGfvt8b9ZljTSdTiBp3h5rsTjEcogsp+GX
uMnNSo4iHzpiRU/Q9PTa/Ab+jt3K1XvxRAEM3+XuoUjEQJgyVvHHvRAKiAgmUzVt
IfzrlHYEJ9bagezSLnnE992JZy928Cw5pxDE9s7F7dx4YX/5+HcNYgJwodtttkaz
EN+bUA3f+JS+/EYscesS1tgM9bMyaal6f1B1JGTK+wqd87hjMRj5ifvi0i0TCe0X
0UB9hvVY0SP8bMecB6UUQbz4JAUkCkQ4q2f4sBnCqs0VUR4TA/5DDKqUfhoattkE
a62KpY2RBFKVx6lYfZ9Jey2qpW34lid2RKDs/k8PG8kBpb4A2+N0wPj6ysnsZGPj
/xwd4PzV24nWhHf4wwRc+bdGtdIBQ4FQzalK+lUVLssJhIbwl30drzj6Q5tucO43
MlTip5bdXYXPvvegtlcGv2gKPvSgN+CnxBQ2LJV9NIdNG9Twa10rN3EOAL7E0w9j
o07dr50cVhX4WO0T2clWsXitdMfgY+aq6RSsynUQZZ/2O+SOH/gSqcuSG70oBInZ
6qKFku6z/prKAe5RhxL4gGLkeWiOXYzlflRxlqYoaB8uik4vI5HeT70fn/oS+yZx
tuU4qCU+d/DIQdqo5DY0O6K8ljslC4ITX/fjVP+MFEEpp0Zu3XgRRyjTgkfPDJDA
lS/lLZ7iucwuKp4wzLKrOrQOxs2ph2TAO8Rm5PhIY07tQoyYFKnKFNLgJvlJkz1N
qctFiTHisV2/ubKpzi0j0EompctdZaOQX+UelfWXxjuHy8g8Zx87IvEi2PUZozF2
Onv5+RNtl4BJkUc+o1T1KsgNe35HtJrLCg2vfok6V7/rbgoSHo1QJ7+8E5fNl9eB
Gk7p6MYVxxksXJrbRbCedvwWS3qhYqyLXFkJPWtWLcKVFwCEM++0ob6HzWQv1vgh
EEUtzvDcrtbYMi8HBNtjH7F60chxIH4hnxkc/0ankHuNe2o8DLNANJDJ/9BDz7Jg
Py19JDHqFeyVsppTCpcLnnQOAiXFWnsy7sk/F5rMW+1KXxiR+J9Tf7W6WGZVmeLo
wZILktwnui5AycFA6SEgIzAhPRZ7FLWS6KK+asNWciqs2nwtZ+Cj6WIlj/W5S+OY
lqr9Q5M4V56+8Mtgm+3JXrvYHIxjbfQNtz+XbHLKw+VP2SIUHHHdWzXgIbIQhxNF
RLgp+KU8AXfWgkbKpFQO/VCxnqITvhNqz2vCrps+c7f6o3+quOhTzS3v1SdJhmPn
wIZwUVgKfxGA6pXi62pbI2wLD1freoTw0r0uPupI57F2H2HIjzLj23JBPKboEPRx
5zYiKTou4g3dcIvT/aYo04+cU/NZaoSGLJKBQiFLy4qPjr9fBb5mB4lGlM0iCLOc
ybSu5i4IRzTkryHTKNtZB/R81yB33Ew1gDKSWN6hoBcXvwjRzaOIAKQpaUYAbfMK
YWJaQERqUdw7IRXmc37LVYoHC8UqczhWSxg5e3PjPh0W/++sUbFUksb0igtwBFDR
+4PPVP9e6t9+MxgnL4OK7UBLyX7afA39eAbEhlTFRlZCuqcq0ZIcMLmKdMz0AZ0I
9Qn8olBI6BJWGyaUfx8BsIVSI6hqMgL08klS/p7SrqNfGUv3fV8efjseECB0NNMe
L9RTIO7d9VXxRdUmp2p8FkMonYoIY4Z+kihjFMWqmkxOshPXFdsmkI6YpVjy889q
qAhuDGuPFUi9O4hWy3Dk/OPszffJQdeS4RiVM7w0SGwj4ntm7C5B1Jf+0xxOJSip
/fdjz5JX2nXkUDT4bldHYa+SEBLl+QdMzGIL6w8sdOn91SoY1it+bxUxvZoYlDR2
BlyeiWTajKzA5JrfkRcenWHp3UL/8fBmvmju7GokJUKZHaEdbvQ4nj3YsLSUFwsV
q3FRP4Kpiyv8R/0lg7sDsYMjlLJknl3YJ1X4mw3V+kQbyHxj0lMe/kVkeKpv4gIQ
pSJNlElUuxNtMClQNFo+e8d7JEPL6um6epoDSIsxp8FdXXw9lTylehy1QZBZNruh
qRGQMFzK5rZS6hH04xLYItcLVmA3Ea1/33+PRPBiAPA6zlVaZdfcj/c4MQFS4XZs
gsWmIBW3fj6HFy38I0eLLa1O+wnSxcPVcEdsp1MemXETN6B07tOOnpAMBdepqncs
1KxUhKJN4uUxryxZLbyiBwhxIFts6eLYj5SKnj27ZJozcs3/kRgJbscyn5ooH5fC
h95gN8VfGhDIrAV8okrMK8pE5PPRFRmsQJU0dUew8EEFi2KpZ+YgUlQxaYobejQO
QRnzoeKUFoGwrkS77t1BxFeHEyHTCRaMMtDLnXCT+nrZqtJNkNPaClKKh/psO1Rr
zJZNPCJak6BGx2uV+n0F76xpcTj3BHjGIxm9WXXjusqb8AJlr9TGCEOX2fgVTKbV
bQKgqFXewpQ4Bp4juHQjAcAn+G40Jb2eI5I4xRJ6cAuw+/YPbm1MPsL6alenTdvH
TiNVlRaT4Sy+oFh498T5UOe5EzZTPfa32M1kn8ybrUUcZa1mfVU+430hVqbWTU8A
HC1YPrkB+Fmd4H2fZIkcFU38i6FaPYSoyiT5LJ65vMF+K6k/DnHxJmm777JrwF+q
hW5ewx9lC++D7oAsZNeNm0nYoOxykK3nEdUswUrCzr7A14tkxbt7jG9lCvp3FnHE
EH0s2TY+vauw5jW80l/hFxJQGF/OeEiUODrjt0bQY4gKWR/stQ8dsUOWNjRzyRYG
3ifPlMFtE1EjbGV190ueqIRhJIa1mlTSdP0sT0gW3iy0UXomawSq4VhGdZJYUUcs
RuhkxDrHg9MFad6URzOFOc2rOhs1R07R0qQhN4Z1ggCCXu6IIMTfoxpJ1C+ZSxwd
r8Lwa11DVFVRRY1D959ArAAmQCTsKhES5oeAbheiWhHrC7fmbcOYVwXDUCyZiySc
V00081Na6pp2JwWT5kEaa7JJJfyW9NdbIU9SqIuqtk0RRcrlT0+seHzINfSzMQ/V
el+YyMbaoh6AIwK4ylNk2oisfJumgCYPRsI4IF1bd6TfkZNyOpJJMEc4+7mlRjDc
pA35m7KguBe33oxQefJwhCgriZqI6tgOMPFzOX+rtA9fPdCMsy6eKQbB61Pa4mIJ
AyEx5Qp0DE48BVDnJ+FRnHTsHt+v+pDVVzw3D7cUuMhvqbAzfrFur2UEmSz4CRhn
LhqDoDfKY7vXp1gYXr/sYFSndaS7xjeUhyjTQMmLNwT4GrkSS+dzOEFoKs91xKN3
tqJzx9Az5zlUHrclsdKidwC/tkM1D2d5DIDa39nP5wFknZAEBBl8Ks+H9g2DlcCh
qnEzyQw/xNrp0D4UGwF2Q8fn2DRa/qlUixvKYtMAojXvhvmYwRHeZi2iM0O1JFak
32GzYgw4OXIH5LN2zBsWcO7ZACN0gIqQANvDwp1mEhqJFTM5aUKjEPv0vzpxfzCs
r8VxH+6sY5ZTn6VQ7rI5XGR+R55UAU/JmeiUo98WGrVQM4be5yv4Mbxv1hfhjx9c
cVXiXno0pjLd9n6dddcG/9YBaLerSu4t6rF/r5VMTj7M2CjSR9Owr9CmaSwfLSb7
Zxu8nB2Be5LpO5TpflEHTLGmAJ9UHvE3chC+w5Bd2pWvnYgbb3jMbndhnN6mpFWC
+l6UbbhVJ7B5CUetKXRgopxkUMB6cg4gdsliA7wBo7uxSGqXxVTZ/ud24f9VBF0x
4eWz4dAQiS3AeNN8WE1rg/ZRVZPFVq7NhmkVh+FTqgxF6jK2yrPLTvr/lbgXzfS3
/6WatkI2pNJB2GecvtNd8uWUkxUouw1mw3/ph5Q8Wz4bIyDHKP8C6hJ8CxbYc2BZ
Qf3hrJfk/JJ/4uOAtUulHOfDMVXmwGm7n/BrmxtWfMS5CU39w5vkiIltH0BDL1hp
x9tR0GPNarEz4WsO/56Y5ueTzaGZZ+/s4PZjvuNlPb8JNNC+94fV1SVZf1EdeDIT
nD5LP3F1eLBnzfo6BGRIlEUCix6dcgKD+4fRdbP6VMCt3UzlxpTFp6iIUYBVY5fl
yOR3NfiBDrfsRqvVYtmEV3J0gIB0S0mM75etYiWbd594xehRU561cULUy/30V7D8
ktfgiqTr1GaBaOMyFBGVUZvXM35IGEhyP0rbz7xH+zMqAqUKLPMScNrVUSUj2DqR
nZ1f7m+7maypVYb8vjjrdOofc0qfcADIJ8tluzjmsUbpZaIyCcUeEcIXQ/IeJHBV
DIKHNj21e356DIlXDNz028yvmfOhG58MUZwyI6pnZoMmNJ2FgeTQnDmdncXBweoV
L5I59OyXR46TW+VYSSIeS7keslRkVCM3I1r4zVWNtOJujsPTST0p/OjX3EBVnEpJ
OIKgqkIYgX2t5sAOYUEqI764n6kni2nB0q12Hz7YWPGsO4m1+jlQZTo/vCmYsQIK
CVIIsuTMYUEOffE457qZynnkxu/evu+i8UisybwPTkN7RFMjpL3Bgjigffh0Pxem
4miL+rx6Avz5ZWZT8JeM1H+cUgXeJeHoPBHTRBXlUYusqKBTs2PNMc+6aAGnr2um
frz6sCexYudQfZGI7Dxq2Xn1pTdj4mycMwEbIyXL1zLnX5nfTM23x4qrwoiQYYZs
SWSMJCb4K7BPbwQjbZqKqYM+CkE/cx2RxGubtipnfTx3Eymn6K8ThnSz+lidAa8R
ePLKKUbo6oLHuLjeyQW34RxX903jO40QTDoU1gORplsLjUPPDzcO4shOB4ZD1T46
MebrROvnGo8YMhunlHBwCiUekOI0ql8pMCc5ixvFNZ25BaMYIexo4W5YMWd/RWlc
GwXGUqu8z38eHfof7f4TGVbKuoOSOexoy/SE0LHeaFB/lCT9BXF5i1oyz9jbtq3D
HPVUJrLfbgWWGcpdIYJ2b/OcBRZo6COWE37t2U4OSJ56nfturgkt5CFBKTYL+mL8
KWjEWa/Ll40pLT7yrEeHJ4Oarx/iCoGJbJv+VIET399Kt83qzAlu+gtI6q1AtJ3i
FfxhAokoQkpyqL1ky3ml43wmwF7tyF9WGaXkNGKOFfAtR42mPYqfmVQkSqXSp5qD
lUTdcVC3iqvBNXjYc/2uxAYZtxIfykbQWmQa0KLZXzhY3Zc/4esyvNOUNMGAh8YS
SnUgSBW6tQu4TJQncvj5x2eg4aG22IMv+d+Tj0SCJIV3ob7yGzBmwn5eFNkPru1g
orN9AR2LBxFZ5s7O6ZCCMCASaOyFqcjrqeuxxKJGIxIlgZURw2rX1pbdM48UUOB9
8Y9eOeME1qkr5KVleS/MCboCJdeEPPUuQX4H+a5lDDPmhiMWfuEZ3KXComGFtvVi
dpvefjhT1B8CYQE6vnq1cD71gNnTb3F0A6/eIrKgBYSXkKKJu9iCYhWWfY6yGEWI
UBweLzVIO7kSZ2DoTaWisYwSICMktRfNH4FsUn9nfuAPtrCc88gWIwM7PNSKt85v
eq07SlbjnjV44gwdScq+m5Qq4rV1jvqRspRoJsEYxbaGJb0/v0hCM3fmv6OynEhn
MYyExAKLa5WFPqcR2iatNXs/9EVww5l7tyri5vs2hel49jIEI/+r2DqfnRM6hqjx
N7ViAmdnfblNBQnZV/0Qu6IVljJjKKkZM9mE+zgBHFh+WqzqV9B1mJ04hd5/Ty97
3FxYySAPRoqAkxSJGa1RbLetGq6oNYxhCUpfHH9gkXUejnjXT5ffodgAlUSLUjll
LMdM1MrEDyRGZHxSVKnoD8/ez/fCfGjD96jLSTRzr0jqIDOAjFdvVUekIwIaiFQQ
EY7iay592VSRj2q/QH+6XnVkBTt6dYzLp9PEFCGJRpRtKCfhS90gcOurkZt6uL8f
75EMdWfH2g645y8yhE1SpI8hgEn1DexfYHXzBKwNjPiqPXMlmczn2GeZIo5LvJwX
ctYGw4YGzG2tbJMEVjff0h6BTYCNy/2pE9hEaen3rxu6r3fl45V3D+Z/xPd/1Jii
YdqDKyUyTN+pQCylZhEmeS0uS3i5/mJekdxyaapFNeXAQqmy1m44xhPHq5TMQT9Y
jIWxUreHaIsJgDKEwyP2ngLSpTbPWRiw7NEgOzZ1UNUiGynGBipc+/dvsXB5Rzgf
t9eczb0S0K/iKIYda1eJl3epwtZ3KS/i1uQjZ1A2sF2FJJuwtvKhpbpwPZt02l4T
AjO4mJ2+odEJ14NIitzt/TvUG3nH0xidyt0S+hNgyhnThZokPpbn9wwNx/3n9DSs
MGM4krwcg5vynCRdhpS4mMFWz81WVtLgm980v0XufWQ7JA3TV16KMnvCRK/gZ40X
1viAmYvNFez9sTb2uO/Y2iHqlyIt6CROl1/HUihPvu0f6Khp6apPzEH29qwRDlpd
Mm3lcWU8VSfRtZ48cFF+dAxaTk/znzLp2+H8UJn9aFqvp0kkuQA8ExwfRns3+n/c
PZ57uopx0RMZMT1J4lwgXXad4RcF77YgZfbphREphHIV4sQFJxBUupXGY+m4OHDu
ZYZQJOVtFM/T6FxbTW0OBB5456XKCa5Sbip3WbXsKFe6hpNe6GNBxVc5Z9U6lQBb
dDD+fSJkD1vq0S06YEVcLBvVbLQm0YyfHRwQqnuQ3N4fV4/2jAFzIp03/PSweUbb
ZAVF+KSOmkKK5mGts8bgSrTe+odaQbBTyWreDepFV/1n4VJauON7sBkI9LwNH943
hcU6TsqHfBvZF5cNo26L9r+Nc9dG2nUuYz5AWLKtua9BLfbYlUBqfGGEO+G5aBLQ
fEIweynrKYvOuDCuHva/p7UrJEAfoiV7nYMg+Qwi+FGtdiCIXmdxVm8+NxHQpT+S
4f6TLIZ9fHsWN1ziYE9/krFWI2F1qFhB772Zlis25CtnHYptVM4+5SQ8zzycl5GW
E/XmLuC5nvJzLGObjv1B1yh9zjBbswPQqT2HAv99DTvLdenI+dxn43BWQH+KSvJJ
Y+rufHWhI4M2tCGbhi4pSXh7NO75GLjNYEr92GJYMMsG/2mBEAykiSbt7Bd4T2U2
VdDx4gh3muFXdfchTVk2AY/TdObiKUOroSrHeJkxDe8OyYgxIiHITQSpOZd7t65e
oKysBya1RESOgQo9lq1QHpu2YZmst5sWr2vCA0WtpsjW+m/DicOg5CyKbKJCu/Iq
f38djCqGt2LX4En+CHi+jHIf/gk+wN9hct21oSacrnjLs7buGZ6NrXuLyKHKnFYT
zQp6e7kXNWI0UA9SjBCXHV37TnWjUpUSm1qDFEQiuGJFW6eunbi4K0BoAXQD0ACo
kZ308HB6/glVntSyX/mDW93QgRLksfRQDrHV70IeOI1hVuo5x20PNAvSMGi9X6XY
xvfEdA7z3Mqos2TwDPPVwHGuUei98/rNfh5tsjPKYpTrTkBhFrPRCZmpt0fLHS3J
g1eEkHRBvx00KzfcFcnFWZLY0Jr4w67QL+jKQzNmTT6W4O3wP+mOeZUNdZfAqXVL
B44ZBykirP2Kv+v0c4loxq5Cq8S/B6/8AGPc97T3HkWUKC57PPIL5v2vFCI2EQy6
Fo6QVPrbiXqPp+Zoj9vxivubVtVKRKkXLrMX/klA4D7HR180L1OjJpDGd4fv4w6C
n7kZvAN5dgClPVtLshe1MDRs0f795E399bAiP+l1Dts76w8QQqYq5scmKLf84ZNT
fYuVJ7WoApPsvHB5wZUmFqvYpIw17alezJxxCkzAKnib1yWLijJZFHGlvQjqR8Cg
4ZG4REP7mUtqo1K+wV3B2qnED69l3eDohH5NJNdnoEpEMVPIlt756zpd1seprVe9
5YrGyptA/+OTmUOXsYZrY01Rhu1bqzVKdor/4QMFKAR2B3VlbAsiNnbX2rb1Wo/C
X5EM9pLQqpM36tNCjVhGt3ltipjdAhBBxZOvQyr+yYhN0pHcwvh3SYQccvv1kzHf
EbzXWbG4LArt4v6+YiMw0vdqcBs9NrwXZ/RlR3mszrJMs4yQ0wxJ3GGKvKuxIZ5Z
2nefQloeLTLv3/T4kyW2p5O8e8pBm4s+rN+ARPoukC31Tr2EvPE+1V3byNKNzPNQ
OKG4VM6uLMVAKerkRFUYF3XyNr8jHFb1+amLsVFNZObiYti6QgV7igpMGgp46WA0
JS8T3ncrqArnw0V4Nr2IwHJa16TKfGmitfzxSOrLN0YFuX6WndqQPmZcfOAjt0fP
ISJTC62mfJhcjFpsmdHIsV5lQv4x7z4yjVrsX646UHgZ2umWB86GipcLG8y99t+I
6SuG/F0sQ2Xz1br8CKEFQbTcl9j7yqmItdI5zRAcKU9Bxc+jVNCdkUWzhwnCGyuU
Xn8vLfvov7vUr+WnE2083Uqw8y7/zTpidyAHXI11wy1/KkBGicJG4lRIF8LFEWnk
029BvhPn1dGBgU//SRnzoFJ+KMwOR2xFhHqNAYR0BHPBwuaJRC0O4oXC3g72FHS/
28QwxaA3xfQL4jYJGhubmpsd8y/NPC98lUNuQePy4XzKJ2xrJXcw17CeJFUXbuaS
efY+YDN8yer2SzWi0HBuzyiOIUpG/AuogBivRRWeJQSGeaiCqU9rB3WoONPjA4tn
kwlWG/tfsUfQAYwMdgrfwnV4SwGjfn/BeNbzxY3YOz6jXiVJbi9kBoGThVIbBidu
EKl4hFHFOpqGK0Rzbhm6IEO0utgRULyyHC/BdcZebSNzhdEoGookI969cY2CUeTL
IloJdx5Jd/+sWvWJJhkR3eX0+HR6dgApgyjJd2JTdN/dQTb12X54iYD+swIH5fA7
rUXqe1qTGln/ez1/ebWl6zKqNF0bTz51lYJsD1Coxj6dVABnDVmKWP6JWCtYXRZE
0x5dfWUYqfeAW4lfqC/hhH9AyA+eKfDpIkeeaKSmayWPXh6tS5UI+trCd0QlTPfb
snzqww01P3GJuTba5Dj6I3oqcj0yjT8J7bWQ+904G2Vrt4sEPTW+0eLsgHg0MDki
ZzAQmreLDzuHYOuSniPcH045JI6dZfG4RrUYz2DmoOf96iuNS9pivf0mqNFmrvSD
duHTuCl+2KzKWAIp1aPhdTb7DYjnrzLWVGY0SUl8a/AQ2na5nz+4gsdB7S/LiWJ+
7W3boLU1ft2mskmgWHOC59Dv77DkT5aHMg92oFDhKAxfbgSF1ka9v8FXg1onwk/Z
VLqlFo6V084TxC1LcL6qqIggNJvOJroq9Rm7qmOD7Cx9tWbDHB57bZxt88k4FwL7
K5Oc4c9bzkWoy6GOD5NWz1tjETrTQWut9rCTpjWEtwfNLzh7kjnn/40ZzQoVIHlU
kZuo8EH5x4DrYu7gO9PGer/2ZEtB3HLfv6butNnLcxlyl5PpOK3pPb3aqz1iMhcG
HgOyvXjWJqTcHjAjyM1zklqpw2Dz4Gwl16eONdiymsZjoRaS23rmPhbvKzu35D7I
fEHOx1ReJD0oTEMEVH9B/0iRWLZZwuizX3ItPYJll24e+SbmTwm/bmMZLI4fHRbR
fQ43Iut4nqzArbNqCGFnshWPay1F3qqRePUOoLjuk4LyT1DtcFYx+851RW3Le9eC
A2Gt6Jg9P7eAXaYzvqqYpTUmGbpURRqihuLCQ8pY4fn/wIanfhsaaYmKLEAI2Meh
4/AHSjff1ILalcBJrFlnBRgkjIrL5kOQgjLK4z9k/QM/i37IMQ2iJBBDUYSRQztw
DeYxxYRVHUGA4tiP6uz4TPzymHSCn37P92ymmgozUdBUbz8GWI47J4gg4xHFiH7K
SGN7N+JsPAMqfbU3Lm+MUbZnGPrXS/0tPoWfvsDqIfdkAxzhy5ZeFy8azk1mO4VC
hF8fIBDMXXy5PQmx8SEYJ9/H/VkFbnLoVq/wekWtecwEapcfyP6uC9FET14BE1ZN
asKR0L6YrMc9Lh6LBanlvp69laskUkI983FYCpRy+1GKXWSaGbl1iEHUQmQWepKW
XxzNRUYXaKMBAHSWeQp66mp7UdnyfcgLEVgvk424HH8fDmsdZtun4CesGcX0WzkI
deZx2mCECpgdVmuGqp28kge14LY40UkbdggADyQJMS1B83ffM9jRmoGsIHHyQk7V
qAQfW0X8JokqeOn54Tdg6mXCaeJiXwiUJXU1yYcEsbCqesHacYcKIwTi8auQj+zA
8ye+UJ8tgv2MOXJ/CDl1nlwRaLE3Hmkj8/Ey9NWMrcxgpfwP2x+DwEbF1NgDJ644
0NhTw4YXPT7v4p9y4lYCcr1L3s26x/RWMQmQzTgsIStY8zYvrToVIJglvtmCjys8
5OxLNSYFgqPaeQvEVglDzASwPm4fbRkecQEtnD1DntIbS0wo4X1koTtvU+LmPPMa
sOuUky9VcMkB+/S6j3nLGydae0Ye5HvnTRCAB0aMdYIxvUY6tPUAnu/0h2O9h12W
v1jRZWqX0yw11nmqELsg/2QbQ79V1u3fbtAVT2L4QOIicsSabY8ATyd96iSnRw37
g9R5HEa/FpHOj8V89oYTOoPUKtZ/ysvOONidzro5K3rUfeJL4e+ETcZNQY7vEDog
S1IpbQlW/c3oG3veaRD6zPKbgpDyZ5oofmmhu+r7xVleq4k3xJI5Qcz8XNQR5zIF
1kyHu6duvevKHXYJCuf9Bu5O47EmuNqm1sUbLXN4CyWwMPHHyefMZCGlkho+OWxY
mO/S6PuUjG38d5frW4eYWLIH52XJQcM24wPH2ZATiNiMOYAwSsobIdnsqOeVJMvH
Q2ntTp+8KiXEvIz4e+2IO66N+oePZhYUUTeBCe7X10F5/pArjiQt+7MskM9+aXyU
0ucy9tPgJlwPenVwoBx/q2OQDXzyX2RoRbvcPngVofFODCC+nLlLreAftICrXrBH
/gxywoTnBXSqcp73elYWtXV/VL/tjPU3QYgC6kb6MLdi2ynDxs0ssks1Uo3gqssb
ALKn7U3w3+LJWBQkHF0Wgwk2+JR2NKamCVal3ZGL/JnBbFonHPamDI/B8hrGzR+N
kHY3pbC8l/RxwIL1a8gPgJ75EB4XQPF5vEn/g2EPRk1kBHF93UAFnZaFs5ArJrX0
hnSHf9tDa6FfUszgg8FDBiLDOEI+ygST1B/KNS/pCGKOizRU/DBlvMiT407pvBDn
RVg86la7Wx589dUnXY96q7DZIlzttUZsAWRL3uPLbcEQtZpP78NTT7LbYG7V5t3b
3kzwzoNmyssaXKndd7g+ep11GKWCtuw2TPC0/OfE4WyCylsiG3ZZAceh5EdCcosB
h/6VJCy1xG0LcPl6FtSqXlv7GLN8Ubs9+srGLCwWVKDgae1l5o4nrP6uXVcT3aob
gbUTZ3MD3v8rIcLibnqZ8U7hpcZ75bcqJ+JxXdf1DhA1D1i/BB/gLE1HOHVT4T8e
Rjkj9Wb1WeER/03ZFHly6mGvviDCcH7a1uf4ndR/g6+gO86m+5p+kcCX7Ti5O23+
MVillnO5IScQOvNHtThNbpLhNR0+1VEf2wIW4NziYIk3/8cXlc4gS5oDIy58eeRP
WyCvtHRMl/0Qinrw0JsAXqWI/DfDdMEIlduSXcjZc//ug2C1tdeIyugcwLpvFjGX
bJknP9TURgg4Lg8urjA1/wWd4TU+ntT7IMKwWtv+N4dAQvSGwSYLzbLnyCwKSfB7
2HHY5modEwDY0Xo53wm5V6bQJl+X/3avQ/SbVVF8xczoSQy8SsXnatTwp1kP/82F
xiPUmZkOD8nLgxSgCK1jIt/584PLix0rNaXgnX0zCyOtK9GxLAGgUL7NXNr4nx+F
vS3H2WEOknAEIs7ki3Fe8oRcXIdpgICZE9NGCdMG4IdI9k40RQcjs4ADNe74cWm5
SUreBnGqVqbFLxAxycNLaorxvdbiE+ZFH8i545L7omfECd/uBKFHCoVqBc3x2ENL
HZtUSH+gEVD8u6ePwrazrDAWNERUI5SM5EOkUoZZkoX4CSWYYFqu/ZCqkn+bCLW9
vsYmU+sGraoVUxRFIPvU8K2a+6saf2lH1dAL1wCry0yidKIgS/qZCTkKh+BDH21y
3sls9kjXIP96IOT9MjAx8z14RK9RAAt0SIxEVOU0utbeNIMuhFeYkUhZGkooJmuT
GhHYGpJHoeqVzpHF0ks96xyKDN0fiJN8jHe0j0Eks1qxK8uIsrvj3bSGAJ2doKoI
LVhEKR7/A1428LbZtsEQOHCzWY/OYdi2y/XgbuWZs5fAusiGMvHLNyqzVAAsGRsw
kHglAZaTV3IrL87/SpcLglAo/gfrDdGvqKjT15kq6//bbPdqWUKh1SuVGnyRfZ/q
xxEYPqIvjxkKhHq7FSIMrCn0xhLjUNFKQOHSOzeWsiS0UkfsmXkV1H5jXtxDBjfg
bVj44/2OXyIT4aXDS1TI7piCljV1bW1Xnx6MlKDFpFDVBBUgy/+JclJdOnkHB7Gn
R0mhpHv1jyHieE1CmS8B++lqponyiPYelMOaN2fCLR7ZfuXJ8T4j8gFGo89iMpvG
UAZ4NSyJrmCwOBvknVDnHzghpLypBz1j5K1fERqlCAi1KKHd50aNMpqwwxIG8SFO
OV+krgc2P/Qspt6sye+G1T3f9tPe9e/vkr8VsaW12jmOVTtmzdGz4aV54OoNN49J
SgwugOh/JEuWihgXlLP/WaGacb8wP28bQAyhEnPXx2/MQuei056cXFtN5NAHw2O3
49VRZ5YmGVS8tEonmUvlLu/+OQeZhHToNsZDr6x54L/Nql8F0SSwI2KwaPsQ+k3r
+jUKOiEe3/NrSC9GxKdhMXbDO8wlVTL2KFP48oOA6rNAvs6HTa/lhfccqmEiKv7C
E+ziVKmgLbUbhOQcxmwNP9AKhONO2EVI6R4ZE7nDrZHHqx6XZ2XKgJW9MLanJYEL
DkxgEhLbNCkBr41eORuNCsBOoB55C79BVWxeM84zyaNIADyvKyB1ij4RE9yJulTr
ukaZBVV6CU3oLRVM+/1Z034HAL3Jzar0KWXr/NecOiFLy0dfVG1qE1HRy6B342Ui
tJ+wPW1tZL3LPgT/6fUKGVaLQYKyAIMtYQdvwK7LQZnElEnJfqFYNUyJ1ok5RuJ9
E/bGLHcutfaSXSnso+Ef+hCJfmGCDdXtZnG3wEKQi62D/3MJ5NixEOARXjyD+WpE
d8ReOHeS9B/BY2Rg37ck7gN7SudC6Ukb734YdXNrRoT9XBiRVlSdZaRT1qM6oKJz
wIUhSLVvHFIqupg+wFuXqapz2IfQoiGdb/o0RML7Q2I+ZT2wZHf+mB/CS6ycP6Oo
rroJ2IOK2Hu47EnZW7PfDJeSR/IGwHL6XZjpXjcvZVvakiH71gQAKr08kZlwnC0F
VqMbWI5PpgzK5O3lMj3MbOf7NpNVkxeaaBlZJrMvcFQY+K/OtvCEAZk+PVEKS/7h
P3UoVTGdUEG6UxEhEQcRNVCVhUAnZC21nZq09o98dlh0e6WsrBQQKhrvw7X+Rwhj
ohrApQo1DCf2yqX+hCSLMekft2nZWWf/QdssM4iz+FWUzXbqa5gvw2JK8IGsJChq
ioMLHGPZc+NmT96Tg1OqG9mPZrsmKexq9Hl4JTvVojkw/Eu6Z23+c+T147RsdEzS
T2JMvxV/z292OBBzxhvtAA5bnbl37BiUHoqrYisiLoNX9L5+UOgt5z/c0P3rQqVl
o6ikNynfDptK08Qynr2v/L3vumkpk6m00CgVPpfPhK3HqqrAoqkaMQ8AQJ6nf4Dd
TQUkmp6wm7KNqC//732B7Tb9/WxrgEfPGTI1B88Ryw1F+MmU715HOiF2fjgsToJ8
+lzzV0EuBCFjAzDMI9zvPSgGqJeqO35x8Nlpk1Txq3gH9NtOOLZ237bex1N6HPj4
gEBbUge6cXudnzaqOeszwfcrrzQp5cjUn2dDiYHuBlN6wwkC4V/bJM7aYRy44nUN
yyrNnkFYRbnH3ReqPRnIEHA5s3rAEBRRwb4Ablri6ptr/iX1tuSblSgzucBUHxLt
6J01CjgXt85Pt8nreb0rCxn/Txiyc5qxYXNpPgcAa1CAJLX6pascEjvLaRQiiebv
3GEZ8uTJwJMXYist5LsPeWMlsiBSKDSVNztOBP34at3A8H2EQKAusHNpGE/AmI2Y
550oDhdGrjiuulE7zR1lCgc8WLRSqgwL6DZBzpS31YZWg6g94zl2mmEFwdX3t9Ga
X5oI4oJ+CWSwPLpc92VEa+rZ4L+TL6BxU86lbAIx83jAZ/cYlIqCxzgCmenlHgCG
fNH4m+GUpKEQebqmBbBb4e7dnb+xkdDqBMPVC9F54iEwHqpctObbKiFbaiT4OG16
cdGQW5xmgIdCuzmh4ZX47fJvefu5+nFi3Vo7IIgQjxQLmkbnjXq5Ro7XHFoebMmT
xnGe1gUWpEHFqgeSykn76rFXWmnydsSFu1XofVK7XaeI9LHZCHQE5omZXJFcemJq
c+7XnwHMNwVhLMhCDw4o+ZfvUQ0/FRHY5obuFz7Gvc0E8U+7RSm2DAtr5AAa5V+g
TGxlke0+CSTx6urXHwYgKIzijG1sVAEQwGo4z7WoL5lnEHyxgfOKqbeu7RbXzOJ/
VecuPz+CuDJY6ZUk8+vQPasZ3f4gEy0PlT7gud1r1yuJQ9CU6/v5vVgxTjx3yjwt
SLj1Rxin6qFmhLav4745LVetzmID8ebhmIgqnJtMlX82t0MOzz+i1KeIFnPLAwaO
yRfVrGKQrCFxrrBQj6QjquLbOmbyxntcJcyto6xFPwCaeD0utVgcLDAPp6uAQFBF
o8Fh4YA/tZAhH55nryvonSpWklAm2ozjrflEHzztpT6yncm7dIejIIKj+tnKioqh
j5iHxBxRxb1gYytdi5/KM6nqD3uWHwqwi9WnaKiaGrDBuUy5TNgQdd4T4YaahUm6
L7BFK3/H27vW4k1hEwMN7FqdmqcYA2F7Xe44ZAS9G+nE7JWG2bsvCQA53TZr00XU
g9NLszpAEC3gBvHRtdKo+B0mWTGH/6IzIkznQUfZM6XolxrMopmFOmcDJDs3hnu7
lZJUpMqmFAJldFmxRS+Zzd1boH0raQ6M4++3ZIU4qQnGvoEtX2JImTa2r8PojrFD
pv3083dOD8LEs5F0G9JCTCAGOnsocyRsIT/DrglHzl9TcSrkjhaEdC1ogSeotHZn
0QimQbkzqvng6XUaoEHNZzmz/6+uwzhebHxn1TkKVi+LypxGHtfCouOpy3y4q+xR
gAivxM5Fcp7XKPBYIbuofTtMVryA8QoBrywoDc1QyA47FD275XGWuAULlkWoSR3P
0czTHA67i7nuQWtZB3b8z0EzWCV+rGXWnMJF+Fxs51/+nF3XV1nyHjfkgZfCe3az
Wgdz+B4RF55hO4tP93FQr74DwfZ8rCdTviK4gSn3UZhmwVrhmDjp/fDHZhPrTu6j
1pWRAgzCoBSJLTCV1UmDN39ziLqYM2PvmBJwLcIcxvCgsx2QGjNkD7RZXOLYr4ry
SCgltsARcSuYYQYXMNRCOW5g8eVJMbhD8PxFBYADDnHhYCIpkUbLbd2HFUq8u7YQ
72nMAGdrP1BuxXN8mDJb/bfXKTlpPFR9G9ItjXKBhFY8Yx2+JpWHjyMV1Px89+Tn
P4eZiECz38D0qVH8eZjLOkfPcdzLlncvs8QesHqnqyLCPoAkzjfd7Z/LBFva/vQq
sP3ysyGrGv1AbBng4OQpQsx5a62bCCt6L4s1Fbu9WoGeO6KEBOY2sHDhL1kgmmNF
g7IQus/i1J/DVqm/5AYNgcb7/GRF0u/Y867rs+P9pMoG1zIsfUWZdWHG0t1OcYnB
2ZU26TGiKWkn2QZE4KhRpynbw5cIiwbX+2H4UMWGhNWbBpt3bM5bwsjR7hDtuQUx
TSCTQ725UjLBSVM6fptkC+VHPwe47OHczy2KebQ1lhprSU6C074pfWxQE3UgTpEO
g2z3AupvbaPQgLUUt8MBf3e38WqlWM45AvL3oGOJu10vEl8PlELYH/LcVgNx0c7Q
LtL0W58je/N52TWZgKm/AjiOoHRFM4iIcfKcgFDSg9gaOWOuAZgy/H/FHvywByGS
sWbBs91wLCTEQq7zELiwVLqbOrIzLMy/zMJPkUBisvEGQ06J+uXfL7OqpIPhggAH
iCNe179bUuHI+FrUevpO5XI/fBKLbm1CXqYNPZYlei9KefH8Zyc4X04vueHcgs1a
d9P+2QHIkB5/3Cvsm2s5owRmOBGRcCncBJtEEj+0H0Zvq0nz7b4fWy56PXfymmhx
1M/P3M9eTgyOUPeSrufu2wcgs9hs5rR0EzRY9DUfCbx9Gd8fCPw5Rjcip4g4crKb
tTBVV0gBqMGRQEOZcVCgHDaW97ijzdsE0E6V2xMzoR9nZYalZ7zsgy7Q+1EQDMXm
GXCvVLfc/sVE4wSsMcAAT3qTPMj076jhHslBYn1jy65Wa5S47nAR3w+BGiya5S+9
2pzoeajYZ3pRqhlV46niEQp001C2K/ObsBUv0pnQyTvBnayaWuFvjkQJZUwr9/Dp
nOw9pIE1cIlDJqKuoHKVu0atOUGK2LuNnRpeL++GAwe4fhOZN2kzoJdNQlNKwIwO
iBbHtEK9QrGh0DoTsWxO3+aryEAkrCSh4phZ09B0RYHUrL6E9wiFKt8+o+DYpFa6
FW2djteILKExky27HA8IJTqc+tortk+DlmHQ802TY1t+RBMo9pimidyG/ObR8Ula
ZkPe1HJb3mNg2hgryP98P2eIhS8G5DwzUMX6IjHN/RBJXhVkIXHtBDRjdvDQuhqo
MlgZTUPgLixP++cTqovQihC+dl6E6og/bNqvmNrsPsEXsG1EcJkxCfrZ48iMbnCb
s5EEUtvAyM/vCO0KJ/ww62Jf1KJdaB20RziEB8YL6HwJVusSPFolx/WLCbVemByU
lC3GWaAefAPeRXEu0g4/WPlvGfukEkLTdLJKESaFc8nNd7++WKvMI773+5rZQWgY
cPRfC6mRhOUmIMw7l50eqc4HFOhCrGYvRS7sgxU48DuhY0I/TyqM7b/y3PsSwT+2
2NlkaDvk/TcfODmDxdzDuCTVHiAKVs8uQSDz3vBcdrNnEkS3qG1rXkFuVRDeysqJ
OdGttSdgkcnEeN0PJ4TelNbQrHpYi1Om33jHgFumXB7+yr/cynWUs5DkMZSXVSfj
bqMyLlm4Qeyg4iAbkQ23cT3RPCWqsEtilRimzXk4Bl29wl7cAES6heqVfaLWvdAS
VGlgD/tlt4SW8stnFUhFbw3WwH122JhQAj9uf5prIzVVmHVQ5cSWJmj2/E+ZMPyy
IrzAj/zdl9TkI9RHfAPh71wQFde/EkvuGfh7QtymT3cYd3PSPbC6J7KBz4ZAl+hi
B9+lL4HsfZ0PT5Pvn4HYIiO48xMVO3oNQgUo5/1jhukTUzz7pOJsQVpRMqvy4S31
+ab1Vue7ay1MojVJ6SkpWV5WKd9viJQIVcAJ+U3u5yoVx14084nr0Vk5BJIFscli
vyB6Vb0rL0HAahFs/pCTkHViZt1qAw00hYEx8Ru0lwmDwOwQjim9sxjtXkI+83iK
aPT1PTq3iN1pp+a6fA77EVdAOD+4gc3/TG5z3G8jsPjw1pF0OK46iOkeTN3TfWii
d7higt6y4ds16WOZ+tQWYt8kfr4EN+ZXcDixuMKZpI4ZF0LAQI3w3AxCSmLCcfuB
nRWou7pF9jN5kM150HeYebm5YRl8XkWsu2Qums8+Ie8K5qRlEthcJHlyO7KHOvd+
u8q7zChl2Aboac8kaFolY1vKVBGh0ZNLXoeKzguAzs+eg8OinvF3l55ytY6YcgSM
XpOKdF2uJho+WNEf9V/umhgvr5P2Kr6onAi8QAtgjnr+/IKrrBPG5PZaF4cBTP0o
EFyIXkasrbKdEc1ZqWaGWQfVdHHluCX+o3BM3rFRkeqh1JAhceFk9APknbqheLxp
cF1uP8nVuPstq3l4qFdp7CSPO+ahsuuwOSgzdhxHqZSSBrj6xala0T93M7I4vXm5
b0b+rr8nJHqNG2cDx7O374nJ8jeM5H90uU+6FagIAnhwP08Jp0iKIbt72+vXFM78
KQdCbfcV7jkATx5bg0SOFBexeAg/y5BxgunOwVgVrpTbS3L+uUG1Fh1Utwv7+2wI
IJDIqguvAiPcvix97E3RgjuKgz0Jo10qFNIplr7iUvwv8Hp5aAIV8j9bMYx3wJYP
NGcLrm46WOGNzOaWo65jf5/rtfy0q9283fTukC59CV9HUnFrDFVP//m9NO4zUVMX
g1UkNkxggFtdjk+1IsKDGPTaL3C2vuFFUCsWFs2e0e/J5+6N1fOmx6z2mPIi8aJX
NSBuGtXCCIzxXNZEJggDWFAOvYAPC+7V6az6G+EOJSAFtadm0IcyCme4xxytkrRD
zEmEFtOCbgCQYOhWHIn2CGIQDbpcOSibNq4KrLWlaw/GP1l5hJeBz5/225BasfFZ
EIKKrwAzHpuVoTPl9PFQ2AKUEn/W6ZKi/FpCj8jp4CRFa0mQAIvFAoLk5KYdd0DX
0JacgrjD+Z8//4FJXbAtBKSKWsInrLZ2vORe9AiSwYb2YQCfXTv7cgaHc0KKTGzc
NKs/4v45rhTUSVBBpY1kOniBUx+vtL0nuwwgykOMsSU1YAcB1DjW5VFrHDsZdg1P
wfl2V3rFST6g2Iys16N48bDipk4HpkLAeCRywkWMb1AHPuBz3Gy6GkjfDca7svvd
V6IpTmmYjbesTEVs4N0RDMIplNuPeloopJZxsa+13wQ2WVw4OedlVJkJv+MQhPPW
dg6YQi/EPoKvhUeep8AEyWhxoao+LopbuCi7+u2m9FxeEqeY1dYguizTZ96A36i1
rzpPFC3+0E4aOeHnvQmaC8ZIN1v1Wh4pHnZrN0zF8YI7yW2bCBLV8Z2EpZANZSeD
dZPF8g5gWxjXX4g1tBxXjVxZkYBR+7Ar7CKUF2S98KR1sICrkWkijrVN75ylzXcA
g0GaYOiliOdLK1xSPrcalgdK5bvrhKNEzuVXo8wA9mQOv3cGH+7wopSNVccsYxeD
yl2sK5lVjOX+tVMsP+Gz/0PKqWF7vMOMAOagmRiOGWwdaqnDYykoeoc/unk+05B4
XFDy9y5Plgs7x7vR7r35MNRnxUJMFobBQo5mDFoKFaOw7Pk7xFfWXEasUcHZ4ZG0
A4Si1dgm+zAaxcT1BWy0aa616tM2eDoG8hwEUheYYhrtPTMrOmA4JukIycWevD5K
WDy3gjrNIMbcslMHzfgQ05Soroe4O4sJC85zr06IBcT8MjLyeqKTXjs+6JPow9Xm
5Nsb0Y1QZK4CqIux0KihoqIqz7bw6/EI0EU5nS7UYeZytFGeZtPm9k/IS4sP4xOA
kMJTKl33kgXyVk6zAeyeuKu2OVXWpERu+AiugUSZXJUdcjdaX3a+xPsBQUmObWT2
QN9mRcsQKvJLoM4XUnpCyFA836/4C1LPXDisZ8Fm23qLtFwDMGjXy+/IYFaKj3AK
hFT/4iQdlF4n+O4cB7NfhzmpziDEgPGQ81WznNoW8vp2/gDnXKMuKHgvrQ+0/XUH
qD5pcp+Fc6nkUgWWHkE1hcO3iJPG4M2ZkESP79L7INtABmTnTBt8bZkwB4Xeo9Wc
VqH1A9rtlVNAi8iskMfL4N6VvghPnIltMdbavV0NbfyTxSPz12piiTWpDO9rbJLN
qcABjFObrx1O29WtNjlpmXqqAGk/PzugxP84Vop8oG8z2jZ2tPALP6X1lK5KKAaV
NG5tfVSpA7gHwnN8i3grBhsXEgKYncaopIhQsg5bJMD5y8fwIDR2DHAhRrf3eS/w
dVbIBmmumwGwAviCcRUWCELC79upTRIXTTRC20ua9XZnXemEcynXo6ikt6T6bNDa
tZH6Uf/3+T/BCJ/DXYmwzQKDmBpi7SoLkWE2EE3PqKoVQcm3r9FyIm7xJPEJY4uj
C0keWmTHmq10888HZSHq2SDMxgCkyvpr5nXPtk29uQnRC2/JYbbU77nNlTgTklnu
3AcVaF3s25r0QVD4utcIWcqr496AI8350vOec65P6G9o02NcowezyLlJMT1i9eXa
0rA7twJZ/dX6KWBiMYtvAwszkfVuMLM78McZTYqmUsu1eC5uWoa1GRcMsJNit4BE
yaXolNjguLc7CgOKB8di3It5ydfmvGj+PmU+NMaJL+sR3KzzpbhthdF1a07fxStm
nrEhJrJWEtfdmdYUcvDEXLuJTBXB1gP1HQHFNWy1YziNqGuYHLKZwdkN35V1WTw3
hy+2RPiM75nH54+9cv43l6+nAWp3EcsihaOQYzSYvznqevUg+kTHNuOyZPgAQCXr
CGfSf3ZLiLOYXG1zsSxFqEzcWZbxzIJlTO9Elkrq9TJ/6NR1DbXlfGTgykiby5X2
2z567iaJn/tTq7FfwHr6fzDhgaPEPiJzxS5mIO4C0XM8emBlJSn+fCkHREeLCABl
vEXgkdBZOSV7LTnyDOBoBAwo6YpzZcyu7AnvA4qDaY264N4mOpjygyix96+Ytpg5
ckDaJxs1YAgXdfov26K0y+J9/BZostrJc9vx3r2Yh8N9KQVQd5UEbdXxrktKgJfV
nx/sAHiRQB/Yn6gE2IIICvBj/5SUj77nju/TgvpQbqOnLoIXiszRQUoSyv3CaMX3
BNYq6NEetk4RXTMsrzu2Ck4i8HB4Rjk6p7JZMSIhHUi6S4vzV3C9ZdT5aNHXasSV
GZz6jarOxpsM6ETPvucMyJIopIZtBQYF/hzHQ4/6xw5x1gwyneiOVQNsmj6iNUov
dzoa9vpVLSjKPEMvcLrj6uiczb6XVut/kPMqcUKn0/8y9eKT6T0Eu0VFBD68ecGE
kV1mgEVv+1AoBszRSEOx0Dz7eElCeqDJGcoIYhrBBN/kmWYu0EXdXY4onC73NL5L
+IKmiNM4uv+sw6dm58NVXGlnitDsWdn0+rRArAimmhyYqqKNdKMWt/ZAPQVMNKCY
zdmRyj3Ad4D5dny4F1u2jKCeNQZmh3KxwfZLOaPog+8y+u20TmDnmYfNQ7Fgd/g5
AeS6ty3stE8/zzpQLdXZ1QKDH8e6kYSogVD2HCRqzil6qO1/D6Zkz8C+gWp+YWU+
KJIK85tLzzJ5JLx5xe4+cs7fS1F04IUjNhTYhXeGaT6KnLfRYYR0a4V13ZySuECa
skL0wqYr5nU8jKDm1Lzuv9dcgSfWE11NiaDA0G6PUjnuCk9mfKM3M0AEWUJ3j6tI
6F90OEquZ1x8veiFMhgMvWd+p6a54ST1n/CicoAt43eGeFRx/3tRvswNgC2Izxiy
mXQjGdBCUKGemtHMm+NC6K3/zZ87NDTjXGh0TAhSGjWB2vFucZpyYduKBcJF5APE
VFKOywLMspwanMfqvyhbgu6MOd4PbwC7qAgN+L1gyn61MOuMVvt6yoo6vc5Pkc0n
oUKP6FvlDzYNB4lXb+aP6eIvLMMSUc3TsFyTDDDbukpw69oW75UYCHwEQi3JU2eC
KXSnp1vCP8eNyV84Ryevr5xsAoF56haArd1C2BoEeT79wX0stppbcZNkDSXHnecG
T97gPlowaeF+gEMo8K8reFn68gdxdXBrwxVJWz7WyakrCxxd4yFCD1KFwCbZHQlT
NypThAW8wK/zx7oj6QdZWXLrHdA/24P/di/GgYNaT1OTQhgTlDNtCYTtUy9iY0Ly
MKz35cHOEQ/eakHP2lf5UFAOmIFmusgziMpmZYn4L2/FS4/AhiACh0Zp3/xJ3CTl
qSAuUHN323SUPAciFTM1kovl1cVIbAG28G5OC//esXcKBX5PXsWfq0LxOWURtXf7
28K/ojguDrl8jyNq3s9/MQTsmXOWNWfl7rhAQiUzLNUb3B57usoImYwdfUCQHizk
nuzoBPFubTkZvT+WzszZZwx7DrN/1JnstWAzdj7TQ0CLGjllFoYUTtbO171KTAXn
hiwL3GOcKO/ff7rOgUlODqkPxgK/Sw9S8YYA0sKGFK/mVkTTPV2RIVBZ3AcDfnDB
Si/lGEW7sttDRDU9oi77t4Q4q2Q9qyYWS6iW/Sfb93GEgES95XOBCSkUYclep1Cn
F0n9CO36/jjgHBUGBU3GKqMUbPiARoj1D9PpYaSnRUT5aqOrxU+ebX1WFO2LdO34
nfMQDjQ8lyXiyTvP+LUOdGHsDaSClKFLoAxa9AIXKAA61BtZH654bblVe4dO7xxV
4LsxahG4R1Y2a+UAojw6TbY6hhfTVbNZJK/1FWcfuPK2rtNKsjprxm1j4yk16UbI
LZ3bMsbssGWd7zbvof0JmVCxjlM/gkJshtHKf/8ymiwWKXhjvy85gsyt+lrjuJVs
/tAljgWD8KJ4oGOh2cl8VDCsTgTIlYtwMFKbsuFqaBvBdt2cfunYtdoYUFXEy1i8
EhYzbZKOBDLxZimhVnJ2LjszA9waRcjVpZpmefECgN5CHg/3pyO8oK0NjLb0NNbr
PVi5AwQMvopUWWsraNB2VX8ceUk4brdDlXeQJ4sqX+RBQ6EUAJ4YQTd2a8eLL6Of
GUge6QTOFXCrUzCbicoYi0OzGO/M+Bwq98M89PoDQ7OPUrNoeKAd5cTBPITRZJYP
430Ovm1J3Rv3o5dZLG30TqSXNRtvtQjeHY0KDCoRsFZ0jl6Z99Zret4oHq09tQm6
qwRZHGtB0BLGE1IMScV4u4j5RHs0nKl0noZ6hRd+2uKJc4QX+X961gAPkKWy9yGZ
9GDH+DnnoPeBtVMNSoYCiKsFCg1nSycwHA2AH5yrEdoepMRNGCKtS+AStMvfytDD
rtSpWhPtWGS/oTLDmRuRUnRMTFEU9FkAXuY4M1RP8IFwTtS0A1met813nne515Q8
N+y3847Jmmob5kiBsj2NxY4pW83SJv2oIrrPW9v3hm3S8+OqqfmoPfXfNyzkznkP
ZAC7FMlIfpUimVd1OPIps4gA9ulJUZroAxbqQg0FA8DhEh9rFAtNmuSCdNYL4urY
Q++7AN7NvV5wVG8o7aX21cfbktCDsEBgxrZGf3ktdCuA62YqmO5WgjzPFgDxxrk4
BMrNtixhHr0GdGkUI9MNjPFR19C33b3eSAKDybDy/BH2GH3K6QRv8B/rc7DbFMLd
EsVl2gYb852G4XLeWK4zxLkxaIvkBk9l4xOuFxScIYTE9oYd7SsWqSqBYN/dxM5V
VQgx1fu6Qw7HxNrncrGvCDe5u4kMu4hxdewy1LHoR1MQqsQRS9KNtdAALB9QxHXM
yHpeH68ZTAeDaoiORNpY9QYxU/mzBg6yt2LIx8SPgb7nce+TMhenvaEd/fEsunp6
/lTTFb07fl8ebI50rBk3OWI7g0hF6y/yyg7AT5GApDd7FTs1Uz3mZmRo+YAwFZP5
jV4ubZP+iKujrb7ypPS/Y5UDb3pya1OwO7Hqvp58WFixewHSTqkYLudK3g9+Ntb7
b6zaCx7KxEV7IBFKTrop8ADX+BwjTnGgL2btcwETeVW9SCPT7CWt49Y5+Q4PsaWL
2wAMev0sZvFL9tDWlW8c1C3ij/qG7SeUfibzg4Lqe71QeN5hksilaktDd8X0KQX9
7HG1dEbvbMH910i+AcziTQtgmHfxUR6gFZSjd9z2YH3Qx3E0IeixhWGbxWnSUS3t
Ib9f0rZ/xXCYMMnJWX52SYKYEyBXg88i+MILkImMIjB1gxQOuKxvh/4gLJXgGz5X
VC9X1URUL1VyyGr4kCSRBQ8+bLaqHzY7JRbo0QsxkDMvieLmU2tI1aWk1lFKCAZj
p9s6y7kang8AAWiQF8linfRLcOIGdbAiSlDYuBp4iBw1r2ooh8TZ+VwuZowmOpli
hf+vlZkL/YV8zeIKRgDYx3Hhj0eHcJLc26EQ6fN3SI+hsz32JK8QiGvDc7/MlL+i
SX15KtxRmDdfRNrBf7uKFVFAgNhYCosCpcaBzIZWqSfn37exjedWTsA4kHXU8f46
Q9NSYoLbKFtL4NMe00VOL4AI3mwlZNF1UlX9ULPAuzA6ea4rlYcz6Qfou1NMTzpY
2zhTGvEZFvXqNwSGZ4wu8oNOWXGXWxdiPDw0kSbUIsYMhI3H87ApexEJ8aCwWFFp
rIUHLMfRdceEiyhOWkpZ3pE4kJRC/08twde3hzfwVHTbDxT9qT2n62ts2y7hGDWc
3wx5eIL8iIuNPxbtVLN/8anSnZseTrYiFawMavpdrJzUPDuPrsdxtP8foOYL5Uh8
OdffSCXNpUa9YoWwnwrWOEdCKQDwfvaZWBDN3ux4dertsf0c5qdz31PQl8HgX2hj
JKSLbMw7Oi3w7GDFY1+0dQ2Yq0mVMYmsWuMIwu6UeFRTwxNxFJjLWNZudTILMrYv
MeZ1Y6gAu6vR4k92nNOTBw0cTrpaq4wOd+PpBd5GqSi6fdN+SUgmZFXhFlEKbKg4
0GvCQ0ShAVG3ZzaYH0VSCWEASNqLcP816ClqrXbsNE+XdcQR4ZsvVe7C6zYaTbdK
osA8YNeMSVFXXMFXiQbgB34xMFOmMLzdiPFUdOlxh2OYW+qkyee3pLp/MZy+W8dH
wMJJe3eOW/x0oW1rSBOitGDs1paKBgODPSjBr5/pJkpXrp7NWdifdGX9Mlv2esBE
zKXOYWwXEUSMtXcLIWJipohywPbLAkkqhjvnRZhosSdKgU0dMXCTlUI9XxtuBpbF
spodFzv7LpHjDlS42SvCi+ZJ8i10eN4+LKTW0WuwiO2AaXz/IhDgXt7uPdJ5zMHw
8xEk2/KSZMAYl/d+3LH8Zggg9AojtswKE7tw50SwM4QGpjyGP4i7UgFQFCR5VoGQ
MgzemRyBWrW4fLhQ6RKVogoIeaOBR0jTjPJYLyJkLocYTq21HtVGZu/s6zGKKAdt
Q2uTTBvzxU/OhzVii862XahlSEwAUlvh2cEPIobNepNFO7kYBHozjgGvwJEMjJTs
W4JynDGFRTnbTAFHtzB7aYfN0dlPCIw4OUrPrCJ0ilkR/1VOKYqdjcGVIY4smiTq
VYTTKOHty/siTvf6XHcLdltRAbv2oiEXdlhl/i9ZWXOJjQmypCNA5csLJ0liirFt
mjjv0/k8SoQrYRfgzNErw+evFj7wORtQN2kRYOaHFKkWRrQXjIQ9nq5ZsytKFl+6
N9P0YIKXTZ7g6hGaVIiPIk8cdOxcmNX6pp9uALM/z+RZ92q1xGs3WGN0Q98aY2vF
EzbRhxUAVwKhEZM22Db2DJ/g2j5Xz/sN2/vikvhBURvyVhOpVjF6Q3aumFPXZ4XI
r9OOiNWRF0evgVKqc9SZyvIZh18EH2oQcA7F27PWt32T1VZiBbDm92LZgRRFdrll
2Rfz7xybkBQEHNHCnKQWeB1b99besW3N6UYgrOn+n0wo37/4Zaxs9bK+TFw/NJ4X
50+IoFY3ZKobirQiAT6v4RZLZrZooTV2xMsrlXRXKxTsS4wELn0oLATSGfLyTifc
DWGiR5EHb/6x3wOpvqKxxO+a/DYi7PW0RRn0/vqNl6N6sfmFfnJ2A7OouwaT44EX
bSNaKpAeaKDI6siBJCAr/Q/SLllgxMDf4DDhNEcsIvi8NYqEIEklnPEFVXD7nRED
Xx6SESEvo0kyqIsZ5/Bjick/mMKegpEUBPodYwvRVf7Iqhb0Ge0OtL5wu1428Lih
Jp4xqTFjIubhaCVM0XhtWtwKk7MFkuD1B+/ViZUM3Vu1BUqPpyJ45RsOVL0bVdR9
825ZdP72m3LL1MExdzrONoKCBJEYnLBUJMKpuylMgfezFPl161zECq3h8yoCutR6
GrGOzSD6+G1RRnITxo/cawMnd8GObWSi0Bm/Tz2zVMTVeQctGz2ZaCvs0FG2Wmv8
wJphkk/I2mUyh2obIJPCGyEvuplJGFRAT9j8F/TjaHs+v4j7NHZ9Ye2mz/8gH8xL
sEAhysQLi14eClBYbe8JUdM2IrVNE0BtTXTMJMv1fiXFMIP9t8AQ9Iw6F4m+Vpgh
jE9At7DQxaF+aLsQf8n7ievzCn4PcJtQE0GdsAv1QkQ0bq7mo5BJObL2/LhZi+pO
4F/KnNfTynWVRRpM5URCHfD3w1QdEx8Ik4Xc7Kp6y3q7ybnIPJON9zG34z8sXJAv
fwg1z+SXMR42L1KNETFO7MsqF3hBu385s/DWaABoE04TzcJaAElKIk4yV9OyyTKX
ysBao1mQZ1AuOLeMkLAuY/XfmVV7cn9aJrlIVUFU/6SdOrycy7PCAJDlIKwFFW+e
SgVHdDEizP1WbARf9kqI0pGVsaqteKLbzFlIflxN2Mspj4rtV5nYIRZUPvnc4+Vx
Zp+zVEBfqC55bA+ogzewVm0LQd05fGBxuYbweuXITflf0KeJGlx3bFp6z4asufIT
MCeP9uCJmD9dpli+3ntixI4F0tsDTaS1Xt0/3+Vr7nQLcjy6BGpRBnL3CAdSXf2d
FSvsO3J/ucO2tl89A6kuKY7GbRYlzWTZ78iU3udOBnf5CCa3Sre4DsJRHSZqSGQV
QzJU4XIVA5XhYd1szn3tw0B/M0lafTh33TiMOJD/LO6B7CzmA/jRbJoASqkNNakT
i8Jbqu9qzNMiiXvYk1lSmwmViL5edcQ6XHoqSMLFL8oUz+M8xPaAIdifTQnfuyK5
HB5+amZfBfT3x6EesuocB8CMZiFJwU0CYv72REwvmdOcoJA0nAzqokYVwYLstX3M
mxVCwpHn7x1087728yGeGzWHNW3SvjITB+nEAyK+f+UJlt+OYpVG/+v/4bokcAlx
kbI9KUDIPk6J+8eYNDzQfpUcISGJ3tW9F/rYWDFbzBxOeSnYZXABwo28SeUEeyob
vr6KQMOCByrhrhUehbTSv2OzmxDI1h8qL1k9v4rlsnPMWcLpsklR4n3hYv8pa3Cr
3UlFq3lkWXED0iegmCYEqJAnVGH3p67b4FTxYHILFKm5A3GlC6ilGpp+Ei5yu8Od
l+IMJwD9w0KCQ9FA7hcysW6+bXQ42g4OhbbcflFXdi2T5EedeKW3k//U4KArLLaK
WH6x9QS2J9DaJeYCX3do+HkczAz7Wm1E6oSji5bjqxuNPmwPI4aRLOa4ceOpvsEp
0xuNlXtwbMbDArdTg0CvCYObcghIqX99pU2gvIO1sylNFQXZCivqr3zrJZ3X1H55
8+w7uurh6yTIXoFWbzlIk69ligtP98KFOb0kCELdmy5iDuXz0Hnrci2x7lU+w//N
rtLW23QZhJMWNRM/rcMf5LxTdofAA7G9CvVh8luB9oPHE628g4IK0BrA8GfOBuZE
PJtVKSqxkknLy1XYl0scDcUtBZa4mJTuM1rdJSr2CaUq8tYYlHKiASF+hEY77al5
jb2ew3p/3JeZi6m8pbb4Z9V6Hcud1rVhXYSuLnEy/exZKVWtVg7TJ5etRIUwRFzQ
pzwNzsHl5cOt/udPc9mUrYnASAZnWTSmIpDk1xMSiu4gRjoojGRAJr5QDhZ1RB84
rCxZOP43bRkCwdbpJL+gATSrEVNLCKzBBwZoxy+1xjd4BDHKmv/cetbTfauYdmvc
OKd0/cGTLlL/luE6/pjUta0y3pyLfHL8gOzFpJ/HGtJ9s6GO0F2ztt8GZrpctEKH
7znm4Utl4fGYDPaUGV1izsIK+3FdLlVq+71A7TvfZwimEOLvIw7ho+oCSTRDK4wS
cyvc8nhEGzE3JFv2hUWlR2WhYTH4npjDSN6kznvJ1c+IwZNIaoyUmxOTd4u6fLwZ
JZjWuI2QnzMUBRuxtra3n0NN3IChTlGX5St3l95UHKDXVY5SzpgMkQ32cYdhn1iY
w5/nIqTu3xTKNm33SoDydkpckgG0SgyqXNt7sYqIOGCiQ9DIlXJW4QHo3AAOMmuJ
z21qCA5nq57uh2p+fS6Ro1XhUfBGh+k2ipbFYx52fD65ThASaNBwS7cfRHcUtTcy
zzjZyzS4HTwYhSEmdT1n1HgjdgRVinOQre4kWjW2lakmRV0MP7n55i/UNOmJzBgV
vnmaLe2WqY4vKMg+bYTfLO++yrkJ+1EuGOcl4OL1hvizp19Emkrp3sRqTCVILDhr
DPNwoar7Y62ojfvZoXeD/wUpg+Lr23ia58c68+ND8+O40S9l3g9N25kJtJu0qXtC
BzS5YetQR6CgCF+rkNgNpU/cVy4/DYNdPHzW3+LPn6aEAtjyXbDyGAUPeyyZwdeR
ehwnnNmwNpv2MP3P4Ieo/5grertSw/S/3m4BYjJRSHsiWi49YYZN0KzvM/Pks7x+
0Fgxs4xMItrcQHhrOfO2H0wbDmh9YUJw/4/vyHh2iy/nPBTE1kbDVNzfOfjXbAsy
ebGwv9dN1zXwxs33eLyqY0VkJBLJ5D5EN0sqCWZ1t78yUYqlUMZZ3FjVISNFF2ss
xcwK2c02XXNv5lwLgnmMeWUgcboc2JP5WrA40L6jn7Yp2jPIXpf6v4BAfZWswNaG
JeKrXyYaPEwXdzeDtIE2VPmPtczXPvJKJagkTgihVt+vPPNCZ9a8jcVHyzZ16wsI
vhZwLiUj3MA36ZQXeDKy7DdwB7643FS6QYhuDVjgUqufeFP9ayJF2cFW9ORUg2z/
IQIsjKbQKxthxy5lXw/kzDrWyZmVFcVhkE3RaJqR8s+hFavPGweH3KZLJc+L6RS6
eFRMFVppKMRQT+JBC7xbbnIVhWQgy8GbAu2+/Jrm9zPDR5XKEwZpqQ8SvBkCoW6W
yFxfm5DbAi/7+NT8eIjajyuzo2adQf/pKqJ9AwcKojGAJWxWK9p8yCTIOSnpar0q
0p63/MLOZ+qVtBsgrZ6GTBQDpFV1ST/oFc2c2yq4tZEvcpKJVKI6OutTZ8rNCm0E
kiHU8Ic3NVfmtiSyYqo/q8FD23PeG2QfFPMCaX/ZYtqC6UdK6mB3hz/csDTU7H9/
EgNKqu4lMxeDODJcgZYnhkdIxVWIfyIgAnkTp8Jg30AQ7ZOqh6JFNCRQRnx51Lv7
lXsnPLWUQvb3KPrQW/zR9MybIIio081Vg+5NqIzzYyPoCecZkDCjerIa4xpEuQPr
3i4sH67/lgZRenZoq3tNuJ3Mp35WDcocU9k9cazjvLbMF/k9G9Mrn531wy2Mq3ox
U8KDRG36ddzJCtvYx4ijhpOV+7CrXtJAr+vHH0TKEIejyDhhbRDFAwD8lcmuZshI
rEBIZ7LEB3XuywObO4Weh9wPECl2QCTTiorR3GeRltUEW4Ip6bYR8qBVyvC9ZgPI
5rFQVzDS8oQM2Bf7aax/DePzmnBJ4GIn9zhLokClN8bu/2Yt+gKtd+kBtizHVkgN
OexGbXohfjQJ0Jh2NBKlMrf4DZTK92lqo7zZJ9mOTvJ/UV/RD6mVXBWrFYiDSHhr
Xo3Sp69i1F6zDji5WfEyZoXv3Mu0O5oYYTiqWXl74GAaOWK79MxWXBkgR5hczvMG
zQWNl3cndImTG8JyrK0fgD/meKK3a5n01MoB3Kud1zTIHhrCRlOQHKHIhVG2wu8J
Gny4tEqrqjF26538wwipcO8g6ob3epakA/BVkjKHvYS5gO8iZxF8wabNUnMRLAyy
9+veJw1BASuIbIAhwSlmHyR1j9W8ubRMbDe8VT8PXEtSWiI4REc2+a6lDhS+Ay8G
gElm31znTfB/AEqAnOs8Zg1w1yf+Q+FQnfp8g5RtEaZS6KFeDcJfFPo471rkWQk6
U5lLLtk/cLxDdu+44QSnmw0l1a8z0JMCO5DtoEzkj4ePZzd64/0UEWROcmYwOiCP
u5AMfbgHDanZE5+EOhidBwJaENgeNZIZ8icvMjB0kHr34YVdIAKT+shvyDfgJ5gl
JEXsicjTYJQX6fBcgd+QrYvMXocuDC0V7b0HxHmMeZNtYLcM+CTl7tCXFSxO+73c
vNs9qLr+3axnhQ6IW+UbJFkW9jaXJSUchtLMxuWE9K6hei9mHrx1/3A4sQMzmdsA
/086S606CdPJhS2yCAHQVjM9AtqG8dcu1jkd4+0kUOABefC7L20d6UmMMUlITGXp
6tJ+0t+xiA3MVSovK6+YlKHlAGRpQ8pRx5/8u4/9YfpUz1QjCWn4UNYYz1hCgRSX
sJASCZPXwK/hiZR15GWh+oR76/AYSR3wfDD6zO2ZaRX1rfPA80GQqkqw1PJPbXiH
sZUIrPcQLfxpvGUwe245EqJhlkLtmYHrHkkt+HcWYpRW8B8K8WV4/TJ5RqJ8TdtQ
iar2+2+I8Mr52gGVqTBpSsOCV/y2S0joXO6/SaWSoiIxM/AofnFxPTysFQojO9um
9191zgofPCuYhhJiYLf6qyAhQFGzV+LiX72AOpsEzR6cAFMZzTDI9I7VPAgK/pAT
N+gnWm8A1EcOXtYrsTlRBBM1Ubn2rlhIyer3/SfY41PBETmxk3gTRwBp1HCKKnCc
BZBLeAuoDL9lW+9tWfr2Q1xspMP/tTnqhDkTOldbpRz8tpKNhdK6VMcE7dEwGLej
WT2+fpt7iSvuI6uW3dZt7YENuQAlEcz5mx1zgjsF3DxfqUCveV8uOYdelOM9wKLQ
RL+GcahtN/DIwovFJP492YVZZISNfpEhrVE/Zi6MLCe5eMfSWP/nAc7Shdn709Rz
b3+WhmNgQShqCs07+Y/HGAetAtPN4Aia0Zh2gATqSUrzkhc+UOZZ2lqnNVgVSyQk
T4boNcz6wbO6E8gZ5EwINVidfFTKpKLfVEHtGfwbKiPlaJ17XD7bOr2IL+7ZeRQc
Sf1OMWdWORVElhbdO/ZldQOT6qBJAe/aSjI9HkocyffM8fLB7J5lTdOh10g/GOBo
X+46zWcRQoBjJ/mZJqfwDTx03UriwInf1x4mVeUcDJ6jpWI6Rjn5o/sbIEj/FhQj
K09Yl380umc19eAlUocaAXTv2Qn54JXcKfUjHtBHu2JBk3NuAPZFAuGp+63ZIIEl
a1sLZ+/G7AkrDYCtByZyon32J0/lg9rk8jcQ5gCFNwrFy7mbVrR6tKg0IerLieyU
l3NMy3JyCHTHuVq24wPx59DIk3Goyl4u2hDvTpehmi+1w4q8XoOt8qe6Ff7wNmNW
z45vDBwd+74fKf3HQ6ptdBlpZ1yqiqp7YJswv1oUmqw8JDQnf0lu7d8wUY2xbh4X
cUAzBBtIPU070RSYsMsj8ZaQqr7YTcnZz9GIycZuBGcREa/eJ/sXrSKnp2vBwKSm
AYHzZx4oLOjQ7kfXq++kL8LlOKrtgpbgn85V/kh+oXUKzlvV0Nwuugk4wFdzXihe
xh9seAkg9FXaVAKRPVvgcSMUkbBENr0/9luLxQm+tmNppSiIh64yNL4cbA4tL1ZW
NLraYtvIWJiNj3gMKOPHUdTDEYkLuEDWkegDFI/DZcmKK2XKwu4zZ/dgtaCQYQYm
plcjxaliYYToiPGYv9nN6WJDBEIFvCsIwg1u05bRAVBkeK5HX6KVancT9YIP8F6H
1/mae6FF4oQXihX4powFIvEFePV9t9Rc2EdEg3N0FM9z+bySp10/Pxfcr6hUYvJp
Y/Nw9k4dxbgLUPYxvJjDFiaBJTnk2TPgXZj41lPmvtILTyFsZsej/L22KCLDcsdQ
BviYD9APdoDjbwCcS7i+0X7LJNeHHBmCfrXGPRCj0UuWaPRuz4abUxHIhQVaAfq5
2HPdRNmdGUzcQ6hpR701p1vIuhBHNYouHk/nJpKJOROxaYA42y8XTkmh59IrCR7a
4g2V3b7QllO46sA7NBUPMgld5ocyrzbCUi1hngnu6KE4WmEZK2bajTnR4yL4UPtv
xKXTuL4ZVde0ye6i073iXWfJK9fmmm2NQ0tkL2LCRSmZBzf+UGYmppAzUXJeiN0n
mzwho/cPkpRAx1WWc2fEj/sPAA6ehXOhPnJZigXDOPST+D78nyRKVUvWH7G5ejBc
zUACPTSYQNi4GhTqGEOCJiInoOcqFV5vbthtcuFtr9oGO+FJ1uDK2T6DIhCfkD/N
eNM473mBC/do38TutGVYaqrYexKFLYDptPpPMtVxBwiartdKKlv2FOawXZpMDhsZ
RSoZcn5kgArp/SHA4hg0Bw1FD00zI7Ur1wpHpjVe5vDv1ehuvVvcBjAAToPnU8D7
kAACvL1nX6HwY/cKoEafeAv0Lf+5xNXa9aZVuIMrzSZ+5FhM3L9LtvzholyT4tIX
NjqHuqkfMx1z8mjwdUlH8f+7toVdY5mECwVgmXB2f18O+GboGU+AMEgGOwQMsyQ6
9+q7E5pS/MB9BuntCXXoj0QDoYBJChfTagC9kPsp1WxY0c6TvoTx8CzqqFDh7Nc+
6e3yrNfgrSKVf3KWQzS4wx+nsxfD0+hoEaRqvzTSXfj2SqnFEDVoriq772IBHOBy
CzJggsUYEgcRA0G7HIXDBrnY/8tAGmgpVYKOwIgJPqRTq9YbuANG1eMnwJvWhcf5
6Q8VSOU6T2WIM8lBd4kKlH9cHJPpMCswpGOesQloKi3f7dscdeDXpV4Q1AHrx1s9
1vf0bWR5yBxgw/SHINEpxClLUl14/RK7eB6yL459TUHcbvHnQ02vE8eoJsvmPFM7
HbzW5x5yYMuTy5ACFbNNL/Xf7X1sse4S6TtleX/bc7u2JVRoOiAMDxWybvAg93Ai
hi28jFzjY3zDKXw5hUOnKpBVAVqBcjcdH99OG/NLY2Yx2A/wCruZqA2GmISw+2KY
CzAsj3wwk6Xz3QzK06YzHSEYSUfXZIHn8X29nNYLQDJYG0k3IkxB0MVCJoXSuqqa
abm9cJ3cZfXimIczY9BJLWcJUHdsyVJSQTpBptohrcOGp4B0UMIw9BrPy1U9Ko+1
nxnfrneAddzy77+e32M1+OaOwxSXWrTWQhmRj+TzX1tr2JbAI1N/7jbz1H2iFfpV
3nrkpATGYc9V0aPWkozGwj3QRLDcMHZVtXWAC7TKMdocSZ0ZRZ5oSYEFONV+OGv6
gdtZWIhKq9Jowe+73Oa8IMZpLxCaeX3R+3QBcTaCUSB6MMgcy7V3GBbledCha0Yo
ZdlY76u3Jemxeq/v6Nq/zmyOIAeEWR7gnahxZBuN8BHv2fRwHsbq8Peo3Ll3UhZO
jykSDmP9BiTAHCGAaDl3FxANdlT3Wwj2aTpFE+325gdAyr0GbJ91Tjpiv9aqdFt+
Y1sUWBq4VchmsD+PR5RXzD5U+YcykesNhJofKligTC+lnq/pCSC6DDnnmK6ejXUk
XUk6mSoKh3qiqreLw/opdChgRznQ7RNpkPBG0Prj3LQz40i/qFfoTcuoIJvQvFSd
fDcmUr0lmgInY7zZ9l7iUzCLmnqor0vaVM9vphj2Ii9uN6Z6kOfur/xmcjFyRIZU
7kW1GUlsIRpyIf8PTtE5jQrDs6XLeHz901TSPoE1IqsVUbX8ZTSCJUfMKigAekTj
4x4gJgHfaYPJi10pilVqHCIo7XuWtPIIGhkNqvcLskLQf1fm0AaQ0nXLSXIfJvVP
i1mTGAxj+/TThpe3co5LCAPmihDZeY9IOg3h6giPx1o/SxZuPo6I7NYFbJ0/BVBQ
dFwLLxmVcP39giNLe22jB0VX/mkqUYgajhSQ0p25yG5hazPj6myOpl+f8mkMzuin
Z1pNor5otGGtn8gxJhi5OtuQiZcn02XxYrFOoeBOkBPy1mlNvuE2XXxzqIANjkBY
aUlclBAc6VOL2YM5Da9yBGELrv+1/szqZe5Xf6e9KcBW+owadFsuB90oFugbjpux
8hFfJ+y3xzXxuCD6Ex1YYV7Ua4akPvTrXJ0v4bMkmpIPFSFXqL6PYy/HNe2Yt1ru
fGK8AL3v4cXs0DC9xu66wFRcI89cEIjNLFTGOydIXquJTiKKqQOpSKybLNKYy3WH
subLs954GmM3Yv96oVtV4ujQAUzD54CnkFINP91qqq2+bIZ0JXchlEUTCOyB72ZD
nZhZDpN4qVpxQNH946yUsbC3chYfHQOZhmMl80AeG7fx4lqvIntnzGnB2LSN9rHZ
noQm1ix86M3Y79daAa44HcWLWUwHkXXqQOsHlK2AbXng+4ym75aVIXYmRBPRqr8J
VfuFou/zyUksB9cK/GWBs2RnFcHg+7ipiBVsfvk0CH8MyA3pLemQ8SY1fifsaT4x
gSgRwcil6iua8AYzzRUmRsD4BGpuQddS7vWnKr7421SjoouYgqz0bIW8dg3k/QQY
dQyCTkfW5h9DhGRC0eCIAIuYSprfueOxR1v2MA8hTNGqPysX24uzGotNkSETedR4
vXzKKF52Iw1Mo1RuKbbqy26PA9IHAQJJUDIH5rOD3P2V6Fzu0PO5hmZ3gVCXp+hz
h3hvO9ko/cHY4rvuu6kDezbl2u58wFWzeK7NyVH98k9YBmYIp94BSj5X+qtTcqV6
wfLYXc57cbUPtXjMLgYA89wt2tfzeeeg9RTwEtaWZFAmnHL01mXC+l4LJErOT33A
s1+s21cGZDxRcJvefFaTqShXaSSUyMq3BiKt28AN3ea4MrZ/YgOXbaiZSH2bpCm7
/Zl5B9LTlBbWnnFAIHW8Blcyx9lR8MmBYMU3hmi9Ea6+muigmSpWBwRQFCMCIkLK
f8ppVFIVoIDCIjH8QVOs8yNuJyfUBG2qlqyCTzkO0ZTyHjv2dkQB9HUDmwtD0ghn
DeGaOUudLi/g7Ag/YtGW3D8TnrZEY2OZYkj+cptwomcT5JhEf4b+oESwqZyc5k8C
wHl5mYWPJ7uyz9xMnxSVeyt0x8djUJntNGPPFTKaBxjQf3tWsGF319edqwRHvWtn
p+jB3ZiS/D3RouoGMvJhmzRaYyytkgxry3mqIdhHQh2gkb+sTR8+Ctrn6IQBvL21
hgmjYcoDkyghGcYBfCEOpGQR6NnLSWZZ/k2QWK7v0gbTGOq+qbG6Fj94MEc0tGG7
Zza0lHQSu7w/kWdxrZcZrkCcyhVtiW1/RIb1O/UxsFizyj58x06QMvKHDOUFdC0k
C1nV/wE32IHRjdtqm777JPdoLrJOhkA3KL+QoA7Go4O0ou4G0D+2EB4LduVlRLrC
IQUlbWhT6OuAL9kGopUgs/UHsEh6/6bThdOrTFmL8Fne6alhS32bQ13w3fNN/E95
WgvRU7SuuUIw/Cj8tlpSL0F1/HqceQDaUfhm6jwKsyyp7NQ0DtahxtGHiiagl/l+
8yDI0x5lQLBetk9y8v+bacNMjizpVrDSLvy/nL1eS5x9FdfBx8j6ugsbR5SBdEsL
wdMI3DJA7KT72pMsaTJuEbTqD0MIpQ1jX7YxOSzlJcivOpj+LsCpxRkDj2LYxm8I
tmYXpRi3qy+zOJnn1D4pBslzwtm04ZMarW9taNLlIXyK8WEWcMEMn+2kjrQGLXDU
nrGngaI9tP1d+JWzTVQWiloOgQkQBj6JJ6hfYGgR0OL0Sx+/Yua/Xk+xhtkuiKDg
Zt4G/dKRlpaLqOXPtcWyEMmBzswQ/qjAmpVkwwFevKZgA4C9hOX0ZFculWEZDYSi
Fkd/vdgFhyFlc2b6NFWWuDvjuO/wD4aYtdU6mON6c8XoX8aHe3EzfDCE1oju488S
/jP9jApbpgdrLk8e5idDObKtt4WTkaSvgBmmrJJCAxndmH47YEH8TVe0hEMVYFoN
BY/qnO6EKtXE+0WjnYkbqgQXl5HopyLDGnob+1JcGYmbMw4UpoVQD0QG6dobF3cB
OWCEu+Xb3rbRDED8tGj8VgEw5AiKQp+xgOoIuzlwQ3JC2dYeFBDYgFUvsN4zGt+F
wAWWwcRrQM2hAD3C0HEL37/5nKDJMXhA05eerDWnN/EuYr1EYIKEHdUDEUv76Rgr
vna7Gu4lJCF37Pi45ptIAYSrEnFecm2Nb75mgQU3Q6Vrsi2TDgT35/UoRAFE2fGj
hYaFQcGowmNLVjvyPpJ+48ar0aPyZJxJ6XBFkfeSDfArNILUQnvuwdlFw93DFs7d
TUnBxUWkZjZAWVYzQZIpdH0YZd5A+kRB1kBYcVvvUnoKvcndsLd9d2aC02t5HsQs
/NvdiwlmsmBJU/jr6+l6sAp6lWxlh1VunIEXVKWJ2IOsqEAXVBuseI3N1K8FlQ0Y
uPbgajhriUbSP/de4vTO7kK9mVMbt5gzRWFM+5W4eIqTBX7fmpcda2bwNVjol3J0
suvTX6PAG6VQk4q8TQlZHUws9MYAR3wYHZnYS0FSAjvbJJboTpI9MeXM2sDx6rxI
yohKECVvFuio586ZALLUYy2YBsw57bQ9hxQrq+SML7ByqVFIWVfEp3k3f03RXhgo
96+Iy8oiF/eViuaoOiIx0+sZQJ/Vfob92JtEe36xDEuwPrdSqHcbnppsa++uYgqz
Hh7KMhu6UeRAPfwtfj1sr/VBCWh7kp1+yr0r39vnldM1Kzj3poFPzGmUvIbJ7eMP
KDyCm3UY40ycjS6AWDSaGU4DXN0K9fbZeqSUfF03lC6LdNeaGdPq+S3r8xPJNqa8
vQYhmTynGvAPX7mVsdjcTJvFzds/iu6io3iUFDchb0LMdiym1XcOyRvHf+MicfIH
ulShGTt5+4exVsuXK3HTgzixN4iUJVUYWhcaA8YmYShcO0bpdaFtQhrnyPTIreZF
PVHkLGygiZ35Z4lXll5O4b7c9WFPGVqi2VmXKNigkCBxEBLDPmgXN5ZGHZBGxqLK
e73Ngbil7xX2I7/lrmA9HyrwgNykpOl+V2xU75H9RY8kJY2g3u5CreKU24BFcYxm
6MQ7Rcmj7PE8e/pA2VbLUggCEf8mvaWMVlRJbehDmy/OQ0/9FKJkNCAPjIsu3/qv
ynVPfC/wmYqEzw4g7lyhR12dzV4acOzdRUUs//MZ7eulMejKckRIhlEqETdkWVjJ
O4QRH1UDMNK7C1zn2jnlt5osGjpE4fJXlBaieLwLuv3cm3n0ebIn8emETgntvmxL
0dVBBwmN96ZSQFp/mKN5tVQTSqLgqSm7PYtWwF/rnYckMiQN0ZWGIgQl37GT0krg
sJ/nGWaXfZ7iiKwTg6oOUqVoMOPCTqvw5AfbF+7VkPeeUp/QE8NZeHRIkNg1YJ6z
3dtNk9P5SiRgscPz849JoKlBD0c5f8y2AjeKCc+xWu5ovugJInTrrTb42cBC5Dl9
wafVlfzJELTFVa8sXQn6NNhzqjwgAvKTjLgKqpdIa4vlVvB2Wjw2TaA0/Z8UqokT
UhKJGHr0igs5xA4hMRJ0O51G5n7yPMAJOKhoi0e0UfSTPCaN84ST3gVzhc/V7M4B
DlZ1wMTAmwsO/QHOL32M9dlE8C0hn2WaI5u5l2Ll7HsQa5uLX2HfKAKYsAchY2VR
3oNFv1HzxChFLAq1Ca6+1CRwHGJXxVcAqYcMvZcTndvaWdge3Pqbc7gBnBKIuWSz
LLBrqAkwjWCs4gk5vo4lDT30PTyWuAb7EDL37bWzmWzW1JspJY0y4x+6FZU/l0Io
7pXvpBECJkXVdRmZr/H0NVk4ulQ/c26dj3ofktvaQEI5EvZSZtnNUvPvsSDo1HpZ
SJLYxNmefW5v3fvX/R3+fc97K2Kr0HanDLCK9P8pJfOcZxK0p2kxtqomj9lniLWk
1q/sMPulPnpeuxZev/sQslzfo80SwGxApnZdLI5b/ZOrmDbYJYfSkryQTZd037tF
d/h7+Pk3+aN2k8VjYJRIMxtXcMJvjRlk3SfOAxB0NpFY+Xi5B81n8tCxisdKNG2J
I3n561PsIoXMmUrGlLiTQ3b7PgYbNHrrLMoGrz7t/52/ySYQkmyRnKpAQNF41zft
LxSx5H3q1YAsVdLqeV7scokEC0bm6z9JN+UmMKqbH58bFtnwXJ+QJDt21gqQtRKA
uyLqzvSFPLSGfBs8nAJLhUGZERhdvr1AqFI/nbN6bFmQl6KkrUktJ3f7590+0rbG
M5v5YnAA603IewGML5EaIjhNQvfFHwB2/38m+UtMszGBFYyoOIyiNLbWS8aMJy3V
OPNdaH8ckpqyeqASXQHAx6C2Vq71Fuw7zB8d2uhwqJKMk496OxOVpUvm7sPO44JR
mg1pNMAHlnTquQuGXEdLUjBUj+OWwZJcnth5q1yxZQPYrv6gyTrUrc/2vzGql4Fi
9X33mUueV61fBAR/tJTBXLMcu12ti9D8lJrpOBbHS52RHj8dQuVtNrAHG400+eCv
Ju7CKVI83otG39epS60xqP2aeruwNbH11aYIyfKNITp4JJsu48w/FqlUi0zBakDM
YlaigqbrwASKVZkSX2Tq+zRb0FSZbOIdMPqLF9x9iggdXWOVMEd3ECRLNuoVEMYt
C60BogF8E/rOBBkLBhzLW4Nmjs/JyBghDGVzd2cDzvahjVc85BLe6OG/PUgiyH8I
2oNZoOlqz1/fQbkuKGYoxAolhyBCGSgjkaWjMhjis/0z7pEsQGRkgunpWKKMCC+Q
EnUQk8F0gL4gLBGvIxC8biBiXG5VfC1tNFft99ay+7W1bxCph+xAlsOWjtU1oBhk
uU2i3PirtmAGJGTYMdqEZJRIbqTp6sNSJ59AI0xZQ75QDsK2qNBgY46gYWGAAi+j
hHHQF7CIFx2TJBks3rwXVX3Xeq1Su1O7EObtkIJiWPRIq0CswjdlhpEdUKOgyXb9
/k2nn1K6zgEuUqxpT7Tfx7oMbfGfiR7ptWTbR20apo0aOTNP5UtAa5WHDy8ZHqc8
eS0rJACalSDHUQv91+hM9eaMD9D1NS/XPfQreMMpJFRGmXM0mfG4uk5AFwmXZc7l
oy4kodub2b1+N64HJQ6UfQ5IF9vDFqyKGMxdVsTekcy4Ba+3pgowXHNq/RWG4LPm
gaQfLxOD9D4+xK1dHP8EUjKFVKyXVfbimS2D2cejrIGaND9NNFvQdlBIKaBhDPPE
8sRCwwjTttTCiD9DMnNuZHlJ5y9LPDTqmqxn2Xwx0t/GpBNr0GuBX4hLh/lsJ49k
bnNKNhBd4ixzb+p+ueUh4F6kvAS/Q5/N+/2BcYMT/9DwqDACF5UfccoSu4qu8B4h
SdU5QPhOwifOuO0NomEzvQXlamILEWWDRPw5sBk+Yidw3Ue72fsQND4wSvMeXiVx
nBhIwfbdDjGdXLl33f1E+rUxHwVUjj08gRP/lEjKH+zRyqfc2KfE4GeZZLHG7wZ6
RvBgan9d0nPQsQMztJZSteWa5zMYI16HdazmoHwefcVbkhCnlAKmlbBMNl0H70cM
ig1CWh0UoXcn1K9JGKjy62fg3IxkGi269gi4oiQYXZMsg5CiCqw2eNj+ryY2mLLL
BCB/1H9E174mRXAqUAaOfHBipmCgSrUz7hFphPexZZjNYDnAiiXoAGPXm3U5ku5K
VIQY0IjmA4z4mTvN2VfFRdHfewkdxH2dnshDpMtVksI69DeZA+aAiK5vt42371Ea
F1gHQ3GiMlU1s9t2KgkS0FRjKBjjRLpuyMYeMR4bXLJHICGh8Y6HjEhdQhIySwOw
hL/B4wiR8skHg4tRa+lpkewOMHcW9GeZ+IiE2wuaUsOzmiNZfl0wzh//LxI6bMaZ
lAZvrwgcKKf9IyJba1tk/dTr6S1Y9rndvneY+B9TtTE7inQTcACX3J7QUNhppvzn
ChmAgKaMpndxQpWvNL9sLCHanAn66ltVIZtgfJlZ0Rox1a/IBBuZTDJGJ679t4yX
LhEcszLtY8SluOCjjv1wGV6BocDTorWmYxrJVwsL7cVr5+ESdCGt1blSmZKttDgH
sryHXP6h1VGk6vPVRs4mW07PkhIg+vMVyKNFBVDCcMuGLeAeCO92zBSBMGNnZrc5
T8vTnelKAL9g9COG9nSAv5BSWes2Fjc1uQIc33ZspBr1nMoTAgyzGMIs6nNcaDv/
sWzLxWIinwvoOS3IkXT6lNhBYO0F/rqtOVI/B3TYk+f/dpcDcxcW2chm98hMFeCU
WQ4LLvgv/EZrvXPcUUOrGZuKXBtNrOXO9v/lL4UdQRtYoUkZMMlTfV9YPxgum+pW
CGgC9GgV/nsDWwljLTh9m52loF/A1UpEJBxCFjO3tQ+9wHw/76WBnLRaC3EEdArN
vPJTgM7n6RLXiALDQ2iveVodNHmkqBoIN9hKV1RG1FuZw1PXE3ThR3Jk4YObeP9A
Q36yR/JFmeMZweYPF9FktGw/ZKz/a3qSh3t5CbprWB2pD2HQZVd6oVtNeB1NSlYY
PMfwfcCNtuGKEAztUJ7f6z13OhtCjez6MiXtPUjJbbSsvvIqnQXz5eNIBWsdDOF3
ZJ/fftvKoN1pFgg/DQqmGfKFglP1ulYoxmW55gU7UQ6AVn/ta+1bmlIjjRusskBv
XqRO62CZrICOsSGYm+Z+OW9Qs+I4+d6EXFREJdvSo2dFD6QFuRZke/68aKiAEiSw
BnvLjSnxAov4xJFMe/7Otx7U9qiqVTG/AgaT5ZL6Z1ueQSvxLxNpqUNtBYa2z3Ro
x9usTz5ZQpcz7zBDe7z9vZIa9pjTSfrHluVEHBHWdLYrYgtqY9yr10JT1ZeHWG17
5/Er09OekdewCKLZl6Cgw/Mj/PGdMBNDIxzkhA6d11r9gtDZHyURcUk7rNKNkwMc
jtpGwNAlBIBoFLyrHpmhvuXEzZq/TLNaExINUtHaqL23YoequP/JKrdMXWb04yHe
4tToN5AmQ6Y4226ul50VFsQHBbICpiUrYdrD4nSMiE/BtEkIafgEQsMvpxcGsqD1
85zWNmnRczZGYvSoPBuWIwCQfNaJCtyxzyHBAfowf99e2uctKLeSqRvY+ZkJLDbp
TRQz1/ihrv8wsrxRSRbDER1ExXOVuzIj3UcnOxjDZlvS5Sm2WbQpf16x0SCHI+tV
rMeyiuYavlTPd+7W5JulMipfubBzbXtPglu4EDWTPMyHLqlyy9T3mJb7OvM00ya3
QCjyiib9deHVJ2LTMpYJF8dIr/kyg/hSDZsk5jxYMdjYUz6eHN3NBaooKflQBk3n
yAEu8wCahekmpnjbYurXPIQYGvoGEYQ3xkoWr4P9w4L9vliBGGudomOM1hQi7xMO
FN/1UVoH3oBA1Kalpsh+ySBWMSa02yH1wi6OJu70yuF/NkwQ5NPJYMe0HjHjUR4i
ShGxPrBJ5Q/Ga4RS0GR+auVLUM+1tw1uEUI34MWuxmLfU5EqO04kjMdmRNevUHE+
6QlXESHhj9EbYLsm7kl3rRY49jm/Jixdz0HoZ+ziMDtTWPO65NVch5/H+PCIhP3q
SN5jofGOqGItVrip4MZVnTL651a3R21MvvzdkdJwJ+6YlbU1YOGOZzrOVoxkOyhe
QekAqjQYiBndfrmtEyewyzRYN8zD/TOF/B6edsbw1LMx0mvs1IANkRrjGf/JDAmC
HLNRjZ0Cs+fbw+DyAZuttyj/0uVDJmKsKvEcVP856clXBdKsB0XXKBL/VYjlPr3M
JnLyR84mzgLDqt7AoPh9BTekAot5dmG3/wL0StSwOxnvOSe7k5+0LsObucGGP6Ar
cEhjtxNq9BlttqE4Z4YD06v0WM4Czw5NYOLAqkof4lPZMo4qM9pwixVZbIGwn0wD
FahvaVv2T78asz3Lo5h8NCmEbY1+kW5tqGPtZGTScShi+DkBrd22BIF7M7MVdBoD
HofElC1xjp/iB0vhWpl2ooV5znsSXou3pVT29IPIN0OpOWz5/HCBKaskoRpXyBdI
dhcihl7IRsICu/1bSFwua9JUONELfFNLRqkUtW1nCNwt/7s/11l7FVbyV6MmAN4c
dfWf5AMJC65plxrFLctagR0q+qRo67Y52+kp+RP9H6B8NHvK8K2fDsiC1Va/hZWw
WEU1hF6iWI4chOXZPLADs4kNt++0z1kXR/r+jR3vbfov0br00+3GaKb4uR033vYq
WsTV8bQ0UqvTFVwACu42bZQORE2bz6JVT6GOb4D6Zw8WtmxC4/69DHIuven5OKgj
r37mBBijClMMq+rgEKBcojE093/FuoSiYBGxpc7KV4u0lV8UMFO132biqZxFPbNM
Bvk3YhRDl2jGGDgd/vN2mE+TzcaE2b2hf60nY+e2op+6GSYDZCQiGVH6JzwefVmX
9KXfOwH4RcJ+7Ad0tKKTJnsbsyAkjJf220IiojXErJ5gGAhOH7SZ3bNeBd8h0S+T
wHP87mbngAOODXuIwA6vY5XzN5IcQF9KgfoIpx0s785fvvwvvuqg4OO+SHgneYBz
vVkpUF7A5ACJ6VJCld3OhxZNCt3ng1EHCmYVOQpsuhngXn99GpmCBPyT2wMtF3ML
N4XJ1LsGWGtHCymW0bSeumcEq0BXhWtur8USuDWwfRCs810eWeYqN1XInmlfJ9jP
eCzrP/qDkYADxvcQr1ZNdiu+Yk/1TsLirJD1EIPZq1bn5893EBJqO7wDk8+K4xXr
NXuSiazEfOphPk59AYJSg41nAICjgrJuBdxMPN8uVAD1zpB47/O3C4uTyp6Jkruq
lQN2rMBNwV8qDwp1HKpV/fnt93gRxIFkU1hVs2zOWGTIbDMt4o1l6MUzbDLK56sA
aFoRSwGFOVLs4N+1wTZs8atrIv6L6Lmq8qP6uBy+qqw0Sou5Iolhv5hnxHEa2N3v
64rtN8LOT+Qq+jnlfNcbN8vqLjcajRSqBHnOwt+38XS1gU20N9pVt7qqrOhg20vj
CUqa7rnULZfNgkIBx3SaVaAMPri6/trdS7jpluXwpwLy5Ljao9wbsbFE1YfN9065
wesseuAwemRnkKN3LySLPWZOU5PLg2N4+IJNmEq4etD3HECRFF5xpYmTPhKWdyKr
nORUa1WpTsPjW5gPPBQlh3Qo2aWztJOShR/usKVbJhCwO/AEQvEwJOUBNOZWtuL0
qM859vlPTgNt5xh6nU/QEtm1JQDMFjNabpO3+Tfu0TJh6iqXzMW9UzAH5fIq/qIJ
4ykylEVFm17LJS34juwTZLgeikZYPReb2TVsKjuPbPffG7UgLWAeaJwCwiJCUwEL
SDgzj/KwGijVSsbvvfRZgkIfgZS7OurUkdmHAoCByLk4yenpy53LFlCNoLiZ7wjB
sj4ekH0MUYHFaEHrN0FCoUc0yVqyNCrfqykiHY2c92sEaSV7djnk3HNODB6A9L+t
d/13wtk71yeeskdG6USUhY7do07bRS4YgUb3k/YEhDJ/wnkJj06C340AiXeDezou
AX4HcSYsuinb6hvJDcU0b+S49hjtl42p7C7jUJ1s3pA8MvX4HXiy8xvmJZ1MDGKj
Hwq5AxUh3tkzOJmbwvp49wim+CgLJjQj7YERpBDMbL9nQm/3VfQ1uZ2kSCzWOJUP
t2Mwyz0cUd7gxv2/YCS8rCII7Zibru0s/y3/q0ekVzgKF4Wsvq5p3XBqaXdlN5Y1
5OsF8tlYsIqqfc5ccWH8rUgCGPUXwdukFj713nHmtiAtDkHSfzgekRQVN4/MkuGk
cSq3q/8bzfWx15/20g8IqAYhvz+R29ylnkGknKzlynpr2SbxkoBFAezwO4hxJmA5
5m38kIajoQC+XL6PiYRBI7hZuI/lLMjB1ZlTz3Tj50wpd0M2zsMgKh5uLaxexrGy
oVwxMgmmeBrLr5/M7RT9LUuBwAlqhBI+ZajFW3sYq3f/9fuUrWBqsUzVAMxWlHhF
B+qRcc4Dpj2j4E77DSS4ZPWwlU7Xyzhf2Pv6a509EG+ysvvS1/1fMQ8PX+4RZlwH
AHbIfBeWt+fKq5w68UMwFdxaBVYR4v54Zfk9wAHaRPv6DLA6J4KscMpYfY1GRETE
dXjRbJK3fjheXkPdQdVwEHLL4mTlcmvcd5PduUpASJOrkYNrE0O0X1yT+CGYwA80
Lg9/YiSFACQW7i/1yLsVPbMy92qLeZM4Wyo0WzK7oNpCDl9LkgRZGyOlHv+gHjyu
FIq3K6QeS4wwdFnp79XswucL+hBwPYyYdWUQL9dZ+UDwY/PRRbyuy4xGA9+eSOjo
Jnz0UpONuJym5fY102DAWFEUId0OMNMUxnAzNsfW/S0Apyg2Cm3dpzpAB7EHrNj8
ENR35QQ5DNdvZsbKz8OKXQ5Pqcii5Yr8kTjfrabsS6HOfLpXSr+N3C7Hv56Pl4OV
NKwsKy2AS63IKvpVOOtFWpSXmfdPx3l+Uzao2l++rcM2nhdAVQeAFqdu6bQV2CVN
8vsqiwVCRev7YWa9mxF8wmxngx7nEsVnj1Iish+vUc4/3+DYCQAUOTXxSqfd5oyD
hYnKyfOARupDBPO1ivsUULD5P8yrzgRBnWq5UQDn5/XhHRZmIFIsa7VIxx4i07n1
wqRwnimFSxz1aKfuUwKxAVpafcLLXhY7M84efbtHAeHVBtiCLD0OHGnY+LxcpPez
MpHB42uWw14qJdX9QIzZBT2dcA7/RtO2PkPrAM+QznNn06aZSGckaqSZrUycqPxZ
glJpNuTWWmA+kOQOUh+uy3F1IBi3d4KmtMR48hIPu/kU7M/Uia2GAr46le/hMVP8
FQpclkSve03y4NENx5hN9cSY/PO0Bd1HHn0f/A8vvR/j2qQYvrL665AxPWG01xYX
CFJMwHPoDdvOWoCeUKE0fF0C5xAWJndLpkGgfZI+pMmfNDsW8yKCdqaBqMVQLcEJ
oWRjjQ++U8mfakBE3szxPifEPZkuMqopJWyr+lbi6bJ26bCloVuPEbRQADogY+qz
582zbG9SiRWOwQ02rMOyJJjYz4aWts/itdaLrhTlpnvt19XZZVjvMqrNzQ5qvsy0
IgDpFWzJG0lbmN96zLe2P7b6Iw4Kb1BE3bXUyzEOkO95BCPyad3Aiup0zKo++xim
iyt+meXPIDeKLNBLOLrRKV0Xv8i9ANAVA+YTSQCQzcVynb7kLxHWiNuIe50biP5Y
9bUHFM6tOm0iSBdGCp+ur1EXdWDxcr12njVvpy/s/vzNsHM5lpuUNMmFaCeKj5WS
COUK/xPdR9rxhRbaFa1+FOeJ3+wudeKM/hozn2n96Alp/q8CiUmxTTDxs1D0nJ3/
FltTUI3XDGxsn/fdI1b1kcg8FXqXxdJ4RC50LtqoKPCBNThGkPrShr5ndDJwNY6r
FeO/M7SFa9/TouQ+gXpEBczCv3zQoBeLOjTQihdO8ykfRxos778IEiDPwkU8Huv/
7pWW5dp3Xn69o8hha4gdjuSQonUY68Hd8hBdPnQwM5Mp1ZxDleLW0Vs9fjSF2nGU
KNLgncPZfUtV2Sf42TpPSS8OUb7Q6jObbhd7U/bDK3yZVnuCgoWLckKoLpP3jdxN
KEih1nWOiZ/WfHZ45cYaVscOxpL1rEq+3pt0Ef5vnWiqgClr1lkrDEm/EYXX1UQf
yNi8oY+ftr+hTzks4oskWrHOuZxz6q1JKVTCQhZ6CfE+Wr6foEXp7AM1TeGAYJ2P
OD7NzdjCXrreeuGp7EbQAzDYL1YyCK0KPOAaE8RP6ARkJCu8m5oO606Q6+DJFlO0
OuoL0PfXwho7M7yCo+PTCwu1O/ROcR8y1uzQfEzHcPjBA2rvadNApKzAmc/sO4Pl
ccaW9BdUxr+Y7jl0Yb1FnnFFEx4I2gRCD4qOWg5HClUDmtdki00X3T15X9/o7EmH
6a3xp0gDwT3dnPb1ZCnLBsUO11XnvZo1HQ7EBsp1EqOu9K714WTF4CsQqXNgqH32
o9FT0J3Osy3hbhLmQkjf0TLPlouE+E/D38d2hZqYF4jWdPdi0VjgGSfxz9xR8Q3y
wpX0cU54JTrL6RUXnMLr5E0Lvt5uXoZCRwo01gtUz3j3vRMBWXJ2Wope0ayRWfsS
abTOcc0e68i/n2WkkMfU0/eTc0BvGHLBVBu44BIHMjFX7LCa561YOvliNY9iaeiy
x+KWC2l6T30rv33lOraa7jPO1WuzsXE01YXPy1q9Qxlr/Vxu1Nfpr9vkvak2AGL1
QsfP9NrM+RUZthe3P6ecvkMJ1hqJleQH4Bvlr0wdfdMent3UIKGVSQPLNIEsUJXp
AreLrfiyw5IAibuelrTrDuN1POxCBW/KYdNn5OSsyHE9xnU7AJlCSnVdRNI8HqKn
joBkN/7rYeyEbLESpempZmDrY541oNzZcraguOOWozUyJmLGi6gi5zOsUyp3TEMb
0KdsSOh/VRqon4WN7yNMSalnRuZuozDhlt/x3Mb5G+T9VZohf7+6iol/fLnB1X9c
LVfzoe8WfjbVG054f8Ji5E9VXl5Q/NHYbxtOm97zEe+7A1Ss0OP05lcpI0xHGoZm
nuVokDV+KRYlG4WffAetMDAM4jnWSq2Fn5ajlXU68NvGnZ2aaEhXD6moU3LvzGis
BiWmbol2AOucLO4eKLuZTx8f8KU+s6rHC3U6N8PB+qFVG5L4y6wkThaN4SRqwvMS
WCBYHnvM79Ions6cI7Jffi8D3fvAasAev8xWdiJhPWs7V7CeI+fvaBT3DjeKnaS5
2/GgLQcaewAHt0GRRZow2DpSenc9ms2pzRYRhWMKjaT40hEYCH+C5poGl+vHkyMc
V5df0MEfAGkKTAQI4KnLJjmTcoKILdN7m1fuoO3JauDN1q80Kfvd2LU5Ykx0XZlQ
Al1EunCqi9gxi+HxT4gB3uEQ9w8LnI/JMSb2D4A5581Oz3UX9SmYqfeXO82A/gMz
4TWXg7m6euhbANtI8/9MHZB6R5DsnWrwOgg+qCVYoJ4IVVw96oR9oQE+0uq/9mQJ
KQL+pdalewtPeCz4PTEuZIm78u5r6FMPc+h/u4kV706L/2F4MZhelGIosJowL6h6
OrtPt78hzZX3vU5RcXc57mIA4r7SzKAeXt6RZFma25O3RhcRQ6y+xJqF90tDs68l
bDm1rUEjZrimqh1EK9Ibz7L/TAO+cPhgIl3rTJqWzqjqrggvEuh19hpPD9vEeGng
woWQEUm0lTBB+HrIW8ofYLyclZM+06sIpCmZABJzf4khZIQUoX0TERzuhkaxbkOW
PIjhbEeoihH3K111UmCtjejJDbhHgPy6kZmAakPwDUCZ7CKd5FIlgmntx3kwpoL0
FZ9MfCPPy0USGd76eOb8dMw6MI6D6nUdDZDlnYgWlXujRjqFIIzwK2J82ssfF37p
VlSymDlfco8PLFcJ+t+9cJfnM6Wn6IEZPV92PNsWecYySyCeZAYuzGw88CEYIHUY
8DHNK9EpUdrMOGIb5BB/Em0bH8eA0h0hZN1A3YqpoP6fUiMPh/UZbGdQzFld0g1L
+qFU4uRMniLRDYsW32ODQXH0vDFvK+l39t4F0iVwyt+6IBdkZ6OzWLBxXMUjOK+7
MKXy888GPpnW63SrN6cng00hL8WWc6qrbjzZW/TuZk2Hml7as3ihOcdTEMBVWaFm
wCdCUenPm/NRCz/tw9A+t/lm1G3ZG+fq2hpHioPtZBnb2CrwvW0nuTnGIXWcvKSO
3tj6WwfDKHiIZlO989LDjhqy3lDFSEfXwGg0c2fjv63KQgV/InWNV/DNkRALKwv7
5i4b4ACEgn2GptHh1tZcJz9dwHL9vO/Ycxbi22kWVZlwZaT3qdSu+uK/aU/crqrH
bdYap3oRxvZv27mb085unJuw/NYvf5tItU/ZVvDZhAzhfgEiehxPXph4vlFE5gdB
gLUZ/58My1hYXt/I3pEoD09n8XVoJlSQTnVYKKmu37kfrKRqdSc49j4bQXLiMjat
YfnEcmcV83PPFFJepwqFMOVUHWnpz5wYlteX9959ragjG5ecMBfdXpt9gKmDlEq8
I9K1wbihLoPIWAyihF7N+Prm5gEFAhXXUa8XqtfOcXuSvS0Yom0z6ct7cGo7WcIb
ONrjOjgOUS11A7w5d8Xl7ulPhLN+mJbo0jPSzUNFmaBSOUk1G4M8ZzZEelRKSrRb
0eS7b7gFoNxfKodUH4K6NVrY8ROsvOs6tN0knqXfvJjNYw1U4qqK8Lv81V6bgmno
T6lD5YgZRY2EefnL/+JIPT+X2jea/ggZnGhKtIa1i8EAfNj/82G2bZLwfwj/ezsg
K5DTuO1RzTCsrkH6ExBl5PqbfF9w21ntX2AV6iRxGRqlMlZXCjOZfsKKoy+O6H1L
uoVVig0IsX3SkpZlaymD7kaCT8YaOeqO4JQquun29jzFSHdHC+InxC2PrWEf987y
cm5zf2oHHbXEqYKfOxckiQjOLbjAVmW3b/QdmhDvk76ZOP+xLZYr71kCgaPstVi4
2mDyLj+TAzn9m9ES1SeLRJ3lpCDD63FejEwTZ5nQe+wN0i9zujE5nU6oMl+nZTKm
kXxn4YUo3nwviwn9oTmYQy8BdZFyvbRjfFP7f6IZf13buBZz1c+HFd4R1arHaeLW
5Xpy084QZ5c2E9Q32fxPqa1CP9Lsd0IjD0s4biFBY6/1ZnWqc2Lc60ZBj1zciJVo
9ThzRlipXvM+mJzm8ePSi24O5SSYoUw7KoFfP3qtZBPUIr/l6pRDwQflt3BtTNQd
dUUDAFc9aKXfduzWOQVoa9i6GN3cDyvR4Shl7tiy0/lGeBjoppd4S5AgVbqQwc8e
1UAHN31s8HnazJnuItaeUIDvRsWcUHc0CgghqnqJ0l6e8XW3cZzhBT3w5AyCp0sp
ZkF0SzqdxbwOtKBWGu1Oy5qwshNqjfs5KoaaAtE1qZ3WGVqC2BC11+9FdCoJKKF0
abgylEbXWK3dbe+C6mXdppM9jmfStj6qGs+X3hQI/gSeXRuHvm9yM+gldpbptmBc
B1ZBWl9db1QNuzNDqtXf67shC0bQLuPAI14tSYViUE/eCfSR1NJYa5LOZVZ/R1B1
UggQm2Ne5nD6yhHNQcS2VO5gzGWqFXJHR74GXpJOCWGzRtN8qvCqlcwAztmIJCNQ
JHmbhFJh9oDN7G3hLx/F6xqx9lkykPqnvM2r6DA/0aCFgbn9B0ujM9+0Uy6oOq/C
dXHx8mnXEcOyj7x9zeDx6nOZsKfL+50j7kQHufxNXyP3rCgjdXXJYiW/YA/fnW36
VJTATxnqkG40GL4SkFKYeCRPRkt9YBiWEl3g7sTA1grKDrnfRmzPNiyWcjS0t84H
jsky2r+ubyJewVVcJi/PzzYtHYetEEC+iP6Bc+chVsOfUjZ6I3sX/6tlialt5SKX
RHqixZwDh3Hsbc9zgfMR9qt+EKKHBc28vW1qJGfvVkGTQ4N+I8PFaB1OLZxXHiJ0
zuyFikL5DjyAnfRMud924dQ+6nf3HCsuuw1tszlJpCXtS82zp3/+w1EtIbdeBiCO
EAwqdhOUnMwnF5/tvIQ2PCJQtEJRuNEv3dHQPjcKC4Dn9D8xz3yNScCQeVpB+5JI
UwyVhOTd6CfD7WkUfVgskerDnKcOgoEB86t2Z1HCL4zGuaLMVb+83vqpNKecYZW4
CHFIqmcHy7DuBoGAuby3KqcP/PyLjWuhXmMPpusaGZVV8dTcXg2+LG5SlEPzNtRY
pBLcp3b1XvPJiTpDOEcLHs90ljJaUFRJDFx3RBy8xLc914mHbG0dzgudhTwxz3oO
2eTM8ZK8HdSOwKuk0ESCCdEZ358o+rkwy7UmpVtL5PRAd3U9CpEIkOaThRbf0Paa
Ww1//r9e0GuLtXvCg0pz/HnHXWCCHV9vd+JnRX2axNmHcfrelrehjR9Aroem5ObD
PkyZhAjkikiej7H3wlsY49atkuOWohmhlHqeM9lgHKIKLe9CuSNRlgotZnEwWsD+
PCJlNpRN4sMMDsrIt/4mQAZWs54VU5+qPGhvJ9JrUlH9i2PyeVqI4oWGgMWyl2o0
PTeyD10Pxx7cfJuP2ZXGHy4FLRbW5LVYNbsr49sIZVyHjmEPZy1cnPmHHEK1OlRG
1aGPflmC1kZXRzpVYz5vUvWYxWS1qMnQkWWYb5OBWP1W1PRe0++d/9gaMAfH9Yo2
1pXDXN/N0lXtAqZX1MQnmiq9g/oDtEpajfi5HNUdWNpa5nDh7E2NEHOxK9V/51Fb
Bkn1sdRhbd1sq1ku88lHSmW0vJcp2JeVY1O4aR3HdVMdYQkyT9XtclddXNhXALMx
J+iaJAHv4MxoF/2CWOCe5PTfaDPB2F4p9Xrqob4XVIWXgx2LYAzRq3+Dkqb+O5HS
8smfKbiDt9GynCYInwVyxMWlwKEm1vTt+ecrWoVJItdjjc/b/93Mlgxx179Zer10
0aU5afo2OAECccmpKoIVVHhs2ldIBr45FD6VrjGQKFv44is74M+3Hjjo3wrBFRoL
7F7T4/p2bGzbj6y/Vo7SxKUVgRDxvjeS4ggiT9ayOA0L2e7klqNWHpLlX4eTo3/1
SuGgAb6OSr6FL8Etr8oBgvuwUqbUjOFEe9R17J7+WdQd5PO5bD9Lz66k2srdAsxN
WQWirHpCnpjvhTD3cfqu7K2jnimMqFi53m2C5pAr1+J0XeNlb9rv2ojgWnqaUuEq
NT66B18vIuIOtcyMoj1eABYjYBc65gJuq+eUBuRVkbbmPClUcApQz3gkm7poVRsF
AFf+eOP+pGi06n1Z22lCChwMP9HKRGo3ynlmvDkKrb97AVf5NmyavlCFyT5hVnvQ
2sUrSStaO0LMs5Op1IpOqE4PAgI0iB3A1RvYIFmeS7/zQWZPp/wjPWqv2bxI7Wid
zzfqB/sl5m+6XlLG+azgi2EaWgQLwS7oHNegVJQiHE3elFzfQ9v6fd7o0ma3mUc7
YoGhhATIFng0yTtMjuq768/5zlDmFLLXUpaSouVKWbl15+DEeLK3z/ltijyAF80A
Au4iYR4HrkeXmpre/qaQXjJD569fd3O5duUVRN8D0pJWRvywgMv9yLsg1ausQCpQ
/ZVby3GZtQRUD7418TfysWRHO1ZuPg+lZgGhEeI1ODVN7nXE1YGR8YhKdFFY7xwM
GjkGQCkn0/gcBkANjg0xIQ+oqHfvf6hDOJOYMimfeOIABb0MmtgvplBLfZEO80tU
54CWk6f6HBD7EqLd9ec9H4U3rgd+cTnbzJaFkQ5ioNTgAWkZdtsQomV/PMaKtlAT
h7bUnYrcEZr3ADAyMvc2awl392VyuIfqn+ZaF1zkhHc3O62EIquq55HupzxzCERf
mwPVI2FzcOWeRe5kdmV+vW/RzCWDv0FBNVujvrzRHgQNg0e+uyk2G4ncfdu94XZV
JKqZg2eej9LGaJ85PO2XOEGfqLSgc3aIusYT9scsMf57SViBai5obKrOW+jmOgvn
2ucKKPyMeNn8AxvbHBLjECaZmMeythxoW6VqfkAPc5MSk2zM4nvKCHFfRzMQzufi
GNuZ66OFvd+lA+CsC9D/3Voyhr9dDRnMAN7lJ2dQH2ho6RyER0eN8VznVguGBI35
xHCImRZYBXSCx7goWXBRGjqU8ukpQVYZenJIUOGNhSLJCetKm2r7A07w/iYSQxTj
qz2TWRHVXPPM27A86c6G4i5g9nJMLG9aJUEooMboQPe7G8Ht96yisaQUjAhx0Ota
OQhoO3D/54Wx6Za7xA6eqXmcq2pTUxcxDMlOcuZn2GAORrgD/WduyTTm8kH5yiK+
L+vRY2cOZbR/CQfhre/5tFXl90G76pvq/VMI81u/D/bCruLPmjQYnPr5+UmO3w1s
4O4Wn0adI7yW6lE5WjlZr1C5YV7+V5qBSqM/sRNUpXeVHSqy1xqhGb5R/PU/qe1o
8YvdYpMX4BXcXnDzrho22o5raCMiqj0Y5uB9VfGRDBjJy+F3f9ayhzv6p2dXWaXS
GwtcgOxhDRiRyVydhke9oT65XBqfyL/lpPW8qslzWsuog8a5dMD4dSQVu4zlOK/F
19WwWRG3+l3SqRd0tvxIfzr88OfMmcwxAscYzqB8RALco/rmnGFdXziC5jlofIjk
bPVbvlv0xYJGbWbWMVVxCAT89MnMwhPw++J0MUHnN4I7JKYfzEvfUQVIR5nf2Bum
eQrf4yeIcFIwcZteRfxMBrWw91Ax5A94tLtanEPI+qzqWnoZWeVNudZGwUKfhPdp
W8U1rMp9/KyLpLVs+WKEnPSXnLY4B5e8d949jDHnaznPrk9uREpRNap+Ae2VvF1b
DxFnanMgMjeEcdc9pjotPrUGfW3Ow/kdlpQNX1uEFO59RB0e31CJYF/ulbYIRfM3
ZF7GRWvnoW0APjCTNnB3Bh9XMNNTU/xJvnR+hZaxa/3lH2JxcVWdf9u2NVyd3Myv
2H9N0DpHdjRhJE2VTeXM/lVciwQMcMZmCFsp5qPwVRcwQAF0t2hVCxRRAxTNRK5H
B6Lg3bGRQKX4F82APS91bMxXSLxcGCPmQeRSqMdT9GbuikPE7RUET8r/Chn2GUo9
0QahFq3X3hhg5ZwjKUWr+fLKiPtp2z8a9WKzYA1ljV89pw7cl+u5tsx9C4LbOslE
zPxPLZ8DzeE47ANZr9EK5J9uVWpDO6ply0DLOKWnmDGVckK4hxc90/UQ9JwvnmwG
mZifaq1/s2M2V7FkWniwkTDyk70RviPhHzxTMrT9PO4pctZTiif+JgEen8LTrwpQ
XOpWk7dQOX5j4XdbdbwumQQlNcMbEyfNS8jfAk4QzZ6Z39HCWjAlHBFGOFR41vWf
gr8vrDgLNrALfK+hwB3UHc1hyCc84FxpkaQA86+QgDycT3uTl8nkIvHgjQhMbyMm
nbd0hMNwUhEySLsHTyWL8LK4niHltq43Ka38bAlzNCmF6Tgo2d0/U7N/LU/SrXm+
Rm8qgwgPg0mhaNX5PdvubYESYR7Gu5QO/G25QoZz4HP1JF9HRp2n77SZGqV94uch
96/5yocnJp02y9KN9U7jtJyCIRJuUfQQkXmstHe4rVgLCoYH1h89EbF9ilap8zrm
W0445zyy3+n7xgAHlDNnPa702DYkKkiNxGqxFnkS76hl3hLaIjgGSt2HLwi0DmpX
IgkmGkkTRk8eMlmm9mQZ0OMuLoRUTTTq9Xwbs1zYTthT19DZN4wk5Y+RoRaA9Tbi
fkylU5b+E0AAs1hPyeq5m9xQJEtbi9oooKib5UHT5fhOkjIRSZn4YHF6nibP0Jxu
cqaNNdjJfYnvTvqlcBfzxhuaKg0nB0FqdZnQ+YA1eRQzWyUTnitV3VzIL5g8AlDJ
CMMZApTP+Ncoo/vFGGoJr5ndvsSH98cakrxv87sPhNuXy2qklDtLEQ6nAgfH+QmG
IVuLD143Qs2larsx5rVN4Jn1HVQdFw5GTPNMcaM7GQgzW2bJduOzqExa4EUIEK12
oOR9W8tmJPTWH4DejMCGira5fvmgxXMOU3AyoVD0lztBCM0TRFiR1sa4StaSdFfN
ZQm7rxb+572/uClH4xxzfbidjgmuL++8/lio0PKDW6PZ48oh716kLy2opbV7azy6
UhVTOB2dYAVUGXIHZMMUFP6UFrQWghNcZbO3cQLX/p4s8z7aZ7hbliqUj8doaK4E
BfXdk4b/AbrdnI8Cc/rMzkd0RwUgDnOPrm4FXrizE9P6xnAcUphOJ7J91PkrtMR0
wH4lHyAZzg9NExXW8HLSddsaG5sTnCnsT9mO/WlxS6B+FZYYylvL9BHV6E5v2eFi
yv7FzzgWlN4WsapHlf9WZG74ipnMhUcQdMn0ODWhoXXI2Ft2y1T4pf1nubSV7tah
0oUlqwtQKNTBOPV9kN7BSe9mm4ytNqpaoPtR7uytfyA/rxoRUn0XKq/T+yWeVLmv
iWXJ17bH7dgJzbDQ1za/SfFoAP5RbtTvZIZRPFAB1DPDvCnVjVPnqTPRSQu6y8cV
it7g7bIW9+8jkbDOiPX46qdtNdymeBez4DoMeKaeUV9oqeergN6uRoTGErd9ELql
IO0v1GVANcZkgekka7tLW70XtQG7pCVRR0V8fF8iw9zREPKSuuNrGOGsy2Q4oKng
QVHocagcuo1lBpI0OcqEffyNFSQxHMueLeztTm1eY9+4ayqlkJxQ85DNNx/NRBCm
JJHORHm7rhuUJC3xIuYvI++onYPFQbNfWfWbJB3GdyRQnSeaInOGH8SqZF8uZb0V
ymA1Cefzu9wAanQpVkSOGt2SP0CTO2QxbbpUsPVvkgsNWsmJdenOzGYSjsKuSc39
b2qX/MEsdXR6/SHwKS5Wp4KtXbbb0t/4W5rJ+/8VE9QBrrKxAJa1vJ0WdNtfncFw
mRyqpCUSwv/vnKxrfumo8K3hXRG9yuiOYkpBYb75IVssKd7Rhnkacl7OAF/fdE9H
guocozjhr30PrVntEbCu9ZKRJFMrtdnr0L8xs8MrwcVPy5/BfQ8FKJd6e/W+3nU3
Jejyx8L8TLmxgku3aqZgqIRBxS1/M/0sRdspg3vAaky9UjKmZ0qF6oHqTccWKIr6
aZNmta4NQESVs24xFp5KmZ2jiLAqWeMkL/zrHPkIQdT5WCTMDnpJF28TgtgFFKeg
pUHy7owQHXQOVWeP9sGpf0BmTXVFMCxPCYOXlt4drNWZrnzZdUbcWEyCIof93B5t
IK0aNfDR0TON5IobxcIvE2XXjHBnVEWJTSEBu3SXtWvXM19/IDygoSpW/BVNa3eo
yhQKM9lbeFfICHOhacCmmLELvCjLPn1nbfdf2lB+lZbUrjI1kchUpuDFwaUn9dUZ
ACXptN8F77vS2rMf5jGpJuR764YbGpt6v55qq7PCO+Djw7II/E+fckW5Wm3hxvnh
t8qJaavfBeIVbfiproX9bmnLO4p7w+XEcM4bPsY2TnNcevoHAOcWIZ4eGzgzhkLc
juXuzhG13FhsWZroUV3Dtz0Jz2CkiYZ1jGsMcfa21Rf521fbDnthmkMGq4k8/YqE
YbRo11MF7sy+6oQwJeYW3HRb5YYLXiMdZFiFCRxmHx7u3w5dsEKojeUzBCnFaEE+
mmJQkPtjUfn6VvgGu6caZliMK1KhZ7k2hT2Xq6lm7+Y/6EGxGDm76Kdg7UQEbDCt
sG91Wy+aoON5Qp4ZzCgbOYa99N/4nidwKDCahzCE2A1N3+T0DNybOI+QGveEzhWc
/q2jz5HGtJTTfK8znq7slYo0zFGIz/s5gZEdZAlUo81CnF5WOnJnQCJuU68RJBrC
Dt2kzJzgk8FWo+WPaoStW81MNZCayK4ifKQd+Wg8AWh+ESEml8lSkaHP5LmoWCfy
WU65IyJmPtrEhqYlmAvhdSeJbt+Ca60nMucr3VjfdXE6gGPYh6nz1s776AOsmSk3
AYXh+wkhMOigaZNP7nZDypDHjU2hn1EP+F7XvXlmgPrAHzD7zv2q6lRI836sOFs9
r7Yh1SJGRBfV/aHUg0vzQzCmtL3RXycuw2cCc7ypxlotcEsgJKk6DEbcRuqP6hmH
lQ4nq1biSaHjkDQHEwzZjKSm/+NDbRYWjWuko/BNKwGTrlWOporynPsBzCDeHzjI
KhM/Vxn1psvvCh++C3Xj1JJxQK8JXW8NozX/j/f0750UYVnMwjgE77X+DPQkwp+H
/vsW17Mqgv4OmyI0hDHU5BnquVd2g3Ew8Wkqy/VTGNrT8AV4KD2mS7mDeGHo6JLK
1jyoAdD2EvBX3SZ8NpqUnmH+cWKvagUJFMKgYi5usP48ySMSGVRu/TS+Xnsx4Z4+
z2oUAHRicagwnwMhTw3pk4wcsd1sT835rr+Bje39vGLNvL3PGxnly+UQYf1VPhkZ
5tUawKZFulW21YiOnf7aVahFNmn4V18NpIU4iL4s4G5yfyFpLY5x/AqMzOqu0PQB
boozhAWUkLUJTsVvdSOvEopr1EuaIAlhoFxJiNySvNB98qXpAM96Dc/jIbKV++w0
uO6ONTC6CTC4IO8i3w3ujdI825GffLip7KRizz+xsW+3dpP2yhqKDSqh9rYaD5JV
aHbA1vmKzNnW0NQNHpGnY5g82n8VbE/P1e8mQOwBohxN6Ai9V2ZtShyfOffC1O1j
fHRFwXPFSGIIE4hHAUS6qf8zHIngZ4sWyzfCox2Hb6xWfIqm/KR2BjUqGNgjTOZg
g2u+4SI+I7EGXkt1oyb/5qJKXYMuPqi41iVUtVQ57WZR/qQt5TJeOc2a88ERJDAA
bPgZbKZS8PKPUZufXbZI+Az0s71vhcfXjk4JC3+L9CKmRD0Z4wO6NIA5clYsHA84
UWJ78wMQkiEK+cJar20kgll/8JM4rjMqvzDzzMCff4VP9BLr4c26P1Y+L8gHlhm+
+ADBe0HJciixkSz85PIEnz1rrVl5JXZwbmCYJ4qSo+Z8I1HP377zGTr/jHoAlXo+
UxixGyykDwcV5Gk51gazCHMnABjv/ZsWn5kLQYONsCglOtaEfGTIYJwZLFLV84aT
U8s8Z1ms0XqHT2eUGNVt7W169mkySEoLiBwDzCYXxxUPVWaeYl7wln01a2drJycZ
VfTPi6CEbC8tkxP2gFLi9Ju07Qj8j8s+7D6iJf1YyfuutQEJoaxylddtOKpHE+xa
AjyPIMsA2W5dPcPaC/438jrrfiEsYVMPg+W7inOCP18octuPDBKcoVvUVgAhG+RI
1TJLZt/A+AD87n8xHoapeJoC9By5p6A5mq16CJ9QVlUrNsVAZ8nsOXWzLUoEs//g
xXqR0EJUOqiinWu2yHmBnhvCmxF19pqcw51vtDIe3bBLQYOwh+Hxo16Cunnygmuw
+I/mr+uY24h+F2zaWlo46a6WVHXx91qZCSZixzYjU44f6iVp1HqMRsPN2kNoY668
4GW7Ixfimd14/ojm9idOni1pmRSFPHoCx4UqWGnS9CGuwHPciuqFrICIpimGQbV6
5PHrB+zqDAz4BPIaphnLna3yikadIvhlIs723aJ+3C4ThnoQbqHsoWiMwHgJQRb2
i3ITzDT3ny4JvnVKO63+7x04uJrA6Gbe5EMhgcPf4KSwaMP++/2gVEi1Wkx9LnA/
9yvu6/S8BgrNEUDHxXCcm05ou1ff043Sp8NnZHZgjMbGuiL2TJZgONo1GbAd79fF
yFGXkk3F/9E9KNSqV7g2snMqUbaJBFcLLaUbQeaqjvydv2WRz8+k45f4o6KcJ1AS
hCiS8JGZ0Qg84IzvAKP2qPO76pq2sz2zbbIOfqlrcYDvGx0Fb8g4XmIBOncgc95L
ePf9+Ok+rqDzGSZFH8/qgEcjU2CxIde8L9fLoXznPT47VQA8u+rFlMpj43KU2lwh
FVRrrackSLmRlHP5xLijC0CvjtpxpX73umNTJiVs0rv9ek1ePAsd4txodWZryZmq
fGJlubmZXsNyR3kRCIPjRdpcafIzFrvixjGFwKf0fFVcYU+9MR2dSgM6S+V4Lj38
mJ23WUDkdC9VVx+GwRcz5n7JW7gXkyQYZzzNgrOnalp10xJVE8VsWhFfw1GYtyKL
AuFBn4jfj+LoM4WYXgbo4M3UsEUcWPHlAaGlTPtkJXX8ppbI9cPA4lv1ITSxECAb
4AceB35eiONWmK5RPCKzxqF3gpTj2v56RoWtwmED60K/jlYndXAV9kBso/vrHhZy
xgFX7tHm2YLAohBzcEgdOxmbwbuDtOckmPdD6wxm++Qe6Iw0mUsk/1HX1QpXfl+Q
5aViU9Ht6z9b/+taIYAbBVlz6IgheEk5iDBBR96rs1yYGxPQW0ngKrg8p3Twhspo
CQkBK+t7y+Ytx7LaHn+1Cxw0pAf4i/4q6ERYrKhej64Krt7Wb5woQK0H9QCu4lkD
/Qs7c7chOixHUz4/b13LKLsxSaP1kOR3H6hW61BGU37m5p1bZVvxyzLm2qIQx+Lf
4uIMxu4l14TeR/XFKrFesEMJge8TeMj/mdEt+mw1OwqvxoiXynSW2dCvBXsPO1ba
lL8DQ9w0V9SRbxgWBl7fLqVNykyvs2SF4anUDYKfRBP0nxzjPtqmUQhOut2gmnkl
Xb3E5ajqgByMbIptwYinl51ySWpyFpkIhGNK2wld2U2010mZcC9lYhPNhA8ktnuz
zq0b9fDB2n7bEtZSoIW3a99W1pSGWujtr62gM36BLWJG8EAkFk+cj1+sZr4tvrMr
H//w72OWCUX0JpjMKcu+V+NJKDzzJc5RshdrePFcQwGEK9eAIcd4+YHIeSGKjfHG
wTKw/WwPstAZbTPlPDEnxSL1z8eO2zO3OHBiaP8uwpZlnq9XpT2dJxJJy+8R2vdW
NaC4IwuDbtLXbBbget5ABbHY5RRw8OLFLQNRZvG3CcRZCY+VYz3e9J8ly4FFUByI
Z4I+h9TkbWHpNFwl2phNI7/Ap9dbSDa9rDs9G5HxEktwXJDWNoxljCth5LiJLPXw
20hfdjoGeLKaVyzCyfKFi/8g9dMh6ZwDnOqJsFGfFvY7YZfMFy76MRgKUuZK+6C+
fUzl6RVO9udoFSRoNy4sd1HmFrkaHxXtQRCwioz0mJGW9Xh/IUCIkUpkz2XcXNYD
pyliwwz5uYPfZ8ZoRJxrnN1NhzgVV5hxTqK7y1Gy+0DGIbaA3mM4ePVevVx3eqCO
zkr92s5Vufzu1SXO6IIS2VFl5Uo2Vo9Kcaa3AgicJsJEhHQ+QCYxqERnwi6gsgN7
P/c4Ik51FoINAMTYqkDiZxoWEwKZITEqbPrwYFAcA27dxg6vKtfDE7SpKOFyB4k9
m+wr3hpBtvLFqh6ixQ7y2qq/qjZ3la/mxBBK5H/RqkU4CkkVa6n5kdZfjUOkAjI9
wBL8wGLU2sVp6qBp8I3cahf/k454hLX9tNmGvf6i3i2DMImFceQBnTmnwoFYxPcq
sGk/2ufWR9YWCsxo7Mo2enN0c247/uq7k9TG+tadGOLpTPDyzlEtwJoUcTz0Om4b
W6c5Ec9vpgsX4mzP5Ya3Bcc2IPnl217ydi7n4+BI/P+WOuc7zr+PuJSzVNt89elh
A0/7mDLVGNWHukAAgpOCbpPOYauRiLmeAD24v9I9YGxmKZ1FeX7NC5bLQs1avPiR
hcRS4V0zwrPYPjN5GbfwXmzBIQxDuTwVtrOqWvfXUEO61NMqz9DbIqWZH56Dj5Ct
iUypxj2Qi4Rmm3m3g8Ze92BS2bfkCok3Dj2zD1yjvlFtQF4MvbeUt0mflHlMYMkp
kZ52IA+qHYhN4H4nwdo76JGuIlNrghH2i6KOo93AepPNNz2Ej52YLBQxL2BMDng2
5RRRh10VhDevtkD5SgNlH1wmrSB5WeOR8lI5biHJ1JIN9fNnfz0JGgDA0ekmpR2X
7xMjaJIRtunGtRSVm6Xo/pDu0vGQJnN8K7kfnSqIxaRhj+28BvumEgUHHFiO6SI1
DHAbtY06kztCrGgEJDVwACNvD3oRXFkGtMh7MytMEhyJgv2LALodzMyCe8ei1N07
/xscbpcwKq7X8e5PQ772EOh7nIZe0ni4aECeQoOSjeil9BA1tVnIjDR+lDeR7Hc2
4PWgzv/VGeGchzjZJdgzPsO1cSYo306co4B4KLKY/rxOgu5hk/vqmm7Dhn6UiwP6
ZN4Vp/8H7fLZwFuVoF6d6lf9G1waowDi0UnJhh7KIcvZVlsgHK5gnigUqxU3U5or
m8VrI+0dKRuIG4C1QvpGRUWyDm0EpDpSCHGl7eS8xA8TwbxDQCE5gXqnzDjAnEPw
6Tnkr13B2SC5VS/KRzfTq2I0/wB1biF1oEE+G9GS97DdjtKtCcMlk7V26GdxCmG5
XYeEe9XhWC6OQk5Ju0ReLo2CpHZko4RvSJBhOFDBwJpKICjZ4rjOQddLgrAvA2VT
OrvE9xtCk5/kP2tKE+RaYbeonqemnfBY2LnhLiQamFEN86uQPdldanX+VmKLPq+a
3n3xt9at5Pvk9HDhxUt3FZ24n9L01DZ3MS36v2unW73RlgOEohB/DtoNJIxt+KIM
rbWho0cIXzt8qEE+3WnUQZdWqruEmIm4H24Ttxhmz8ouQKk8bQ9vEszrXajiiHDl
Ur/OG5snD7h2K47k5GOPT4HsPIKSiI7Q1tcHgtPTBPsYdQ18ZaxnvbR74IQoD89M
igPnKsAkqfHOVK15lVzOXXWg17FTRKFqQRARdltFOln3hpC9PuHw8CiLL1WRRlFG
uf96bvyHYpF9eFdCFinVzxtSX+VKSUqfylGpvUQpsUtQuKSFM6/1UidoRaisKjV9
iS1RKtuKMpW1f+e/XaqAlj6Jrl4jbxbNpBurQ7tuJBDw/yhhKuINFfNBd/29cBI9
IqR4+5p38AzUd0gjcAXQ0v0nPbv23V7yacX1lCqbsh39yhfgvJFy6JpOdD7u7yjH
j5qJxrm3hQ3QnJzwy8kRnCMF1AlgmvU9+VDc/OtQBFQOYX9XpdqEZ5m2B5VFDKoQ
P8hz09A8JVUd3m2Zh8DW5owMCI9Ue0pzNDZ9hUbetvP0E/NSAyTjARq4A6HloA3B
HVeDDNa5PRLYMa4iufPZZsZmltYk1nQR7yCBhhuJbOTjZFCUj3LIBeBB+eqIRBh8
Ps2hcVHBhlF7xkNwlxZ++ONoxeFvMaE1nQBlun6pGm/0UxIOW1sk1LbmcVTXJwVa
vQidAvummsFTZ3eRlCboSxCvUBl1yDg4bk1YixQEpGSLlH+S4Wt5R7dGne2mQ6aP
mWKneRcZUqXaxg5sxfu5qgGlEYEnPKnW6JyxfC+R3+MrMwCWtwAponbP9VdNbJD0
fvvVfj808aO1wUml1jW4CADSULvUHDMf+2G7YgNLTzMT8fKOezsz49ou3YlPYeGu
b11t7bKYw7lVjdlX37Ec4tnKIyE6jNmVgnHBarl5VTvXEwR3wzX2qSlnPF1NfBHa
2JeyPvVE4nK++ck9Gt+oSr6jXS2fo+v3vWZ0rlzYGsnS2MNVbgCacDORaZk7GTZ1
lzHiCJctX80LUy7vRW5n459WIsoo+VJeuJ4miPlnIUqDkScU5kwrM64+kSNJzZsp
bH0hnO1hVDv6Od1NTP7PuW3TdGrB8vII8pKg3Z/NMXnmoJ/vVKWq4NSLK6GCBGlG
0RkPCqcXnxtSF8V0eHwpLkCc+QAQRzmOM8X2ofKgad5H2wn6GBcPoAFVgpqESq9c
4nsfeH9cTSA12ktJl8h2YQ/jTOr/gohIkFiZXoNTYz2/yBcKucYbmDhz1rcdzVi+
C6UoiavF8QBmznkmv95GvTlODSqbnNzSZugPYT3jdFKw4W4DUhopJFpV3wifjARf
AyyOuI/AJDBSXq03PekuGeQ/T7ZN88I7zx1NzSjNC6yXwBaX6AEsv0RlmeLy5238
ZXoIH4/eOw+TTAzc8pFXi73Cb1QtFSSc1bw2TYFMC7teKRdP38d/HNwhNYC4p2qu
ybf+yEn1MVKbzMw3u1HPqZtduS6TYMk3YvWTr8dtWcvxw/j3+ajKukm5DUQw1v1s
HwD53IO+lZFD/x35W4peDzWFwubr0M0TasP6szzEsg+KVg2xl43K+evrLNS/uA3k
xMj31bnKu19XVwO5juDdhq1zm8ibYO3pqI66ADUV6aANrXYMhOCGQMn55810FDrn
+Ky9BvO8Tq/WUjETdZBjwZMvJXDlxBOp1qEI6u3sJoPlG7jvPPT1309Fu9Kyjiau
rSbxr612SGBg49whkve7KV1b5xxacqr6emqBhzlt86Aj/vynAxrs94sa+nM6WCGd
jqk+QCuCpJMCXksORFWTV+SDb6LGInFa55kR3FL7XCzUbFUUz+G32Ox0KDlRFCH2
7gFhofoPkDC1tx58KB7d64nzRF88rbcZUnNaaNEXThflwCCXxYyaKJciLV3g13JU
y1ex2oLZVLMERmC0L7cr8PNv2k50+x8shBMfG+HFfCPSodd3/1f1PmvubdMRVIKc
HCscXR5K8zsjU9LCu4ZSYdqaR4JTK7bipDim0kuL5bk8UziZHTziKUWbcIY4MfcV
FBAZNgu6XUzAHXDdguBKdAr05VfddioHpw/ck6uU2t109i1HxMuviYbCbWl1OS7Z
7zg5XowwhyAVSpBcQsIy6Ak6ShFFUMKnRtuEYKqP1HxHCVLJctmVc/VCOtvZ31Zv
9iycIzQQZBpTA9J0f/vBA7T7NK1N8slKX6OkU0qT/uSuUejHg4NieEykdrTZISlP
zFAT7yz1gWgW89BVqHf30am3srO3eFGHumSUCtM57IKVnGprz+KgwQfvaMoOEDRT
Z/pslmuXkMgrtnM/gRVWGPwMzjb6R0dhSL9c8+T85egU9CQv+RR3CMsYHXQ8Fnng
pz5eHmurPzI86N2AeA54vBl2NxflUlqOcfD9dw1QY2a4n0MaWEsfUse9wt7GeXrI
R1neFIU+rBBaSZNUbQX0LI+foAodddvPGexhZYT+kCvYx5fIlar1IjuLhiFj4weS
V9uVY90mhhWaNemSaQpAr24TtzGqqEzYBMlHdf7z385wY3GGVW8IkY9z9llhRxjy
0Ny5DuMcwcm/IGdQjL4Mg5vDAbckV4+gJRKVAgbLRcNXwyb1JvsDJxPS8iESix9q
7SngDVdhnp09BdGljHIRLVZgBUbg9lawuOoqj8xOQiuNpWNqLht2HiMT5VfWacnK
5Nic0wjpYWbfJIoAqh14pM4Xvbf0HaUf0mFlCYZGzpfHTt+akJDes5T4ouH68IfG
59F936koCfhYzjyKGAAovZzmDGCRi0nTiFDEvHuAvOYcb5P8sX3p9DmCesvcK+Yg
jjOVqlBYJ6BGTT2sYLEM13VjL6UmfDSX6wcgXa8CrkbGCo20SDNrGfbY1buK2rJP
feWU04w9iG62tscAzRoFXu0B1pfsdBwWr643Q6fTHT8RWBtL7+uQIrvWX154lyFD
EWvb3RMqI2AU/6Z3F1k/c2EXV7cFMVmbuwJgHp+kQFisen2YzySCVEFQxByOIWyQ
Glxyn+38RGhPQcZm5KZw8D/3rm91I3/dV2jlsZNCqz12RkavoRkIkGeaH8eNL9Lz
55tm+2ATCPPKx9uD1B+2/rjTk2mkt1nPpUO5sUoGM49VMQuRFW/YdsLKGCsTFxUQ
cGJS4STeoBniVA2m5MRyrW9dhsQr1zw6LsphrToxw3UiThrGyGcRH571+0M9blk7
ey03Qn6QuqKN91y8qDzX8eblo4pxETsHW84HQ6zZNfSgVoa9xrL7Gf96oxmJxhrZ
W8PfqEBfWJgIlNcDsL2cIank3BUpRqfvNif2qXdK/oBC0QqXJKf5Q/kNDSdXvg79
JMBNwZidlMkGzJpx42klbRn9Dhp1UdKK2vWRf56QWVkrk2aB3uEg5wYVSnr5mmPw
59BjXTrKlr3+Qhvyx6qrwYWatThVrYwaunxuh8qkMXGXqL/8Xi6kPM3qflBUTJ+5
N2XMiWtlCldQZd/Nf5cBcflHqnYiPB7UwBZJ7uCKIdeEhfJNEQHMrk7uMaLBFBDc
LIwHOCGazaHpjn4gVq1OHLqmCvXJK0edqeWJHhRxkfYKFveFM7GJoQDhODFXXxue
Z7hMkTNsrW8f4bYpoW7gCFIDm5ZoDuiebbwc7vjrfzfBURL9BuZq52KHqm3fHXh9
7kjEOqYaj1ZnRhyHSgql+wNp9RDidWgc1XrH081mIcoUuggrV+7OW8BmNaR1FJtj
6BkmtN3seiUI0XyPo/FJFLZtw/VLoYCGjh3r7fWZiRNwKg21pKeMzgWH1dqLPrNZ
kKOXChIKyw2sFCDT6TMEmApU7teByv8EHcmlwddBUs15wkiO5XsQEeKXJZ8pwh2B
87bAEUohVqeIfwIBBapT+kkfgsV0xmmJ7wtzYdwGnZZdikb+WrYsyVGF1kE0xz5J
tZUAhWk4ApLm/hHGLwzupwp00jeXQylpYpueQRDq31VojNZHjPW9mNmtKeU5I+ur
cNuhn8mqCpF2AEo1S4uO1z1X1RkxQt3hjrSVuZDwkUeIXNfOkH+JgBZcE0M0LOZK
ammSTHg58UnmsCLi0WXZVkhHJ4Vb8OsICfdbaF7nSl4w/xGy5HM7nANtv9bZvZoD
MFW8CGElDlrJ3s9LjN/+fqMYXaSXMmuiQB+6KYyXmCxXLO1a3Mx2f64YbZSTXAU8
U0082nb8dhsFL9MYxK83FDpmbR6zdJZIW0NFcgGYqb5dClbOqxvytk1bHxGVMIbT
y30MI+vRfcpbksCYoi/qO2stPfKJzyyKP+9YYTSpfHfYayejuWwucdsoX2Apy3cl
PRHfT8k1xMcYNdW12RalsMAiEq4jPidhfjPrutARqIjF2+oRoQBw1WUUPvuAnBmB
a0CPttYnv2BG4rGCokEqFfvc8ewfA9xUBsJwioCLaCOaSNvxET6LeE9ROpzMc1YY
FoINLS49D3d+2y+h4DKy0VBvWC47IjcG53CQ9MOsrtHM7H8dXwNbNFeEE51rWpnZ
WbkTvaw35i64IHUJCOVomUVRreLIhlRM5YYOCY5oXM7B7A0bnq8W/AJojx1Bkwna
iXcOkgQGnzFANLV/LxwKqhaD0v3k/CML/ouqL083Zr+KG7MBdubqoLp4+w9Uan6w
zMUyRPZAq5yhJORHv4IH2KAl3geejs/yyitwFxuyMBZb5t7F6OeEMn3s8zrLa10O
OPd27ltybyVdho5375pMwcfJn+rpMMGYh2YcoRJQXafHzgkz6nLozsEmKJRy9K9D
KZx5AvUPBKO4UrVkgkjcAPwT4usoNz2YNvsMU81VaoTDszV2ZOFbZz/++65ogKnU
zf8jH7msVUg4tRQmDS2hW/3cs6CZ5TImuGY9wlawNjVaSWdWNLh7wpzpa/b6xJhB
hRLPbmXAj6NgElJstu9iXQO9bBsUMAlJc9Jl88ZJ7rMRwWjfbInXVtVohYIo14hJ
oCIpdV/6x53RqDVHrbVZRqzbP6BsHbsYUzRWSYmyusnIxfw6AoTLi84IjNYoiQP2
iIziGCBXwmEkK712sIbrvy41RGMtzy+L671K8AVH0AQRGS/etCLtenqnJrXCFd+p
yC+qRV3uU0tg0zZV1yaUWmlbqVo2tdpVUrVX6XDmMOFrvJ/W5haEgNPmiXyFEuf0
iXhOGmm7K5/XaYbJIZNpqiWM9Zz3x+Z8qzibgd/WGkB6eaij+/WyBJgeBXT1FWN7
/SkueEIQAHascz+229PbZ9T2ZygXKgTNV6/LooRVRnjauFs5SxoKYBsjEDakssJj
f3RHDgmm5++1D+zzn4Zca92xlmWRur2fjXntpPPN3NGXF2EgxEhk+pxnc33kuVAT
82WU3QDztostVfj+Y3wtT+veYQ05oDEpjAp2ewrn7Sb33l0h2CIyx7VfmibxFVID
KuHkll7UR6qq1b+97aebv9ZoW8GoofjbkJnXS7XLQ78Fn626oIE5CfX8Kt7krCvg
bI3uGiNADeX4lCJdwarJ3y0R83UxFCs4n59BV5KaFVwuUesRNPwCEedm5WaHQwya
O+SqovkOAMyA7wCSRbLzD367VoDf7JWkErHBVheSmG/72B6AVaDhjbBp6l/bFXQQ
T6nWd7sJcJJbpdknwQ0ghU5/oTvVRDVmHUIZjZk9VKMiQu/dJaNk8342+R7sXuUV
qmGzmhUF2MEJZi+sFZHaVsmGjg1rC4/EmjY5lQ5Ub6MeOv3PcG9+KL6GxMB8WybL
32I3PIIqOv3RaCsfPRo9LwzYHW8PDcfAi48ViRTd4tNl92MWCSiuZkk2ZuHaDY3B
4LCers5ejHQ5DtrJVeSgjahoP6PW//L3lDAPfd/J4TK5z7c60YvQyRviBwsmPnfH
DmmOy4GjzcXEnPz2AFaPtkIt+Ybhsp2HY/UD8AVp2tvvfrjK8D2YcInQH1T3cgEl
73aa8lvdwq63F8E42SZ+34VNeGHX78RLuo5s4uBSy/MbtoMbzX9Z1eDl/geNDMhb
sVHQwlwyIlQENJkqSlLfU69Tru2ZOamtxUoem6Gwy5C0OnIYJiGmHCC0ygHuO4d3
V72RdK3FGTCH6Hfmzoj95j1VMWS51s1WHVfBTiCAdq6YY98OJg9isZD8M+9GJw1/
virBf759zhUPis6a46tHTqLYsKkxx6jzZAPXqvG28fkxzr1kK5oyNerJmTMeficV
RpE3PiRYHErmAhxvJT6gAyvRyuSbkswYNJZexa4o6UWIYC4wzxakqhoN+7Fcqb7f
kSxXrJF/IlNvLGfFFwre55nYWzIx0KIfVywgFxYNaI8RioSaSilNVnGRv7+l3X4T
2+BoFFgGpYQDv68WVBZ/HQErl/4jvbSaGzvTYbRXypjLbp8civs3w1cBaOmFgM74
gIDdrEaw+1Bn6uoT1UwGvxl11LtMrJEDF6Z6wt/QEdUcx+YAPNYecBJGljWZdZWr
vs5FcPIyksWI9VFd9wx5w5QGqAAB2SCIAS4QXL0tg7Tp1t7mhmbvy6x9TwEiDFIS
cO87ugIDsowVlnlBpxuoCxWCKTDdjmIKrNbSmdgFej/g1J85EyfGxaU3bmdhc7gY
X6PO2ajlfcr9OaZMw6PGGRQ9drv4hJLwTfaqi7t9ntvchpthE4WvJQYXYnR7ew2s
F9ul/VBhmqEK+xXcrW4fsSa8mBbNQuglKCVkBBfo1U8GT0Jh0H1d1vbgAShQJhzM
+uiU3/5+dznSKXg8nUopJ76C1XaaWKzqtwoV+EXWjYzfarSic+ILf8oYL/EC2bpa
z/pV10ysN7Vmw/MIygwZnhkuaFlKfAxHCd7h51Irl5lDvIPYcnaoAfzGW6xWcACS
0aognSVZpImKbyuv1D63v3Q+Smkv1PcuxRYC3RGjxVcbM6oc5iNdQDgmo0c33M4d
VYeAeTYS20crKRNKLbGkdQGY2xwDwbJ5xWiubXvf3znp0IAq0DpqbEob9vmSe0v0
uQ8AK37HjMlHwA39znYyTx9euPzjw9p59fQSkKhWn7qmlnXjU0e5LhmVF40OzllX
sX6W/TEQK4Ct+ZXsgvF37E3yypcaGm0+kJAmHnSkJcH5dJU5mZrnh2iGr/NRCYZo
mYiemCdMFMu+1sotCCbIDsTON3s1FBh4B6Y1JUoBjjS71KHLVnfmVZr7oxGkmHVY
UsdRbd2jbcuveK6rv9BrSzi6D9iVr4AzRu6CNzPdtkfhcUbcUgGGZZd0le0oWZks
s5xyQAl75BEq6B1PDJpa2rsR7LPmmys+tQyVn0bXkWSkr+rbyymAAOFglX+LGwd0
db/NhlSB9KRD1hzWw6gmUyn1wH8o4N6AJao1ai6VsAugqRpTIvmf15sQQHofvJXt
+Ep0q+chkG3mh4SdC7JzOsCZMCj1ELf3ZOo7+KYRcy6Pb3rargZ9hXT4205IhKno
kdMkhUh8Eu4hkWuf5G662Ce2e+3lWYWSA7xJOJc5pt3VLX8MVUSe6+/7FGSKOAYf
s1zlpwZQXZV5gV9V2bWD1y049W5ZrsPRxgKK2L9FoOmidja6/oECtEXJ8/emJuxx
OkIlMZMQ5cdc6uoLmWoBtBiKam2pFSPJb/dBQmhzCCrCMMF5Z9fIkAKpsTNsYYW0
LkiSHLRLYNsffSFWiE4xx60jCObcLRX7lhVmlm5YlfIpsuzZ1nB83qZoPC8sqllK
+KOL1DjiUkoi3meGlPPGLtnV6uvukfVIci8UmKRGSUCZpmNF4azH1JZNCbcHZQQJ
4f2DT+ArbckLPkxwEZaFs6QEfuS0pXA7GbsLExh0PCzFubnKhJ6ZCjOe8LPm5Xoc
DXIHmwUzXuGDtMWf8VMRCf3qxMLTACtpORyrvhmiI99u9SSxdtWvKCDCsLkpwmhh
kcVts8RhdtJaxv/PGTYI4ZLE7ILnEv3rBKdiwZOEZBoYclZ/sXliwnQzPJUYiRJv
ps53RRcvVXmNxZuk9NJrzD/OoyPQez9OaqDHF4UNN/eTpTMuTiXoKFc+5W1ZLv87
O7g19MgXkt9m5Zo83IJgmEoabo0jM50EjjEw4/xLwsbrIQiVfa0SXF00RcMU1TyH
S2EWp8Eouc9kT5/A7Rf6DFXK2UfFjBnBlHxFi815YVqIGACDF1Fg1Yv67Mv+eD16
IfM+LLAMnOUUdzvJhGpGXFrsNScGrtEiuZG4/s+83biq66gczIbUlCkulBLLhc+8
j1svCF1rs0sQNGjzCBaMozNewFCO1tdroYz+ZFD9rzaGpofmMG2Pbwnk/kNUSglC
UwJ/CJzaa+28z/IgZIMu+YiDGTM8eZcu9DmFkaeY9f05TA7IV8BMYvorSC0n9S+j
chuTs7CY2A6+P6wS6NCrNFkb0QP29FNb0Xp1+yhENZiizIP9bRJmK4rBGfLM5AiH
xa99lZHCT03CWwCew7eoLcZVsK7XzXVxy8ExUUQ42fzvfX3kY8inDLRC5ecN9zyM
AFziJYogxp0kbSeRgjbzAwpiH46bbchYfejt8cNuDhyjV/V5/gAXI592tfN1f83/
cfpnoCIPP3ABdgn+6vw2b6iJc2p7lcje9EJVmVR3vMoMCV5+a1iTFFAom+PzRhF5
wfqUFZ4VlSXE+47vv6L4FVFZGTIoLcMeP0ZyFZbPbkOWHWEMkzIXH8TlYPXyp7O1
y9n1qTHfJhyuABUV2L9zI3z+QVvDvaRihgscOQacLtHqftIiq1soy569MHYS1Plq
6VfHmB3plE4IVVoYfD2/nsdGUUQQIEaApFlhk9IHbGD/10nLPB4fQCcHbgt4IVZH
KlCrEa/8yiszMrne+JgjDZOv/wvrwsyVnAUUCMmhbX44XD4xcYPHxTgQJs+57Cwi
xYEeiouRYKlslpsQqJ3cGTZhFGJzNd994q5/AJSohtlPBOeS/Q7C9voc4keECd45
LKuFYvFPKAXD4LrrQFqUkysjmTZz1ejdSeOv4K13y57Y39HWFNem6lGi7GoGVr0J
aD0WB9gGjUkE7/TbXumgmZ7g+0DKVP7W2GL6EW3xKZIVImWhdsbVfrKu4jWHnomH
iVClXjhdCSn8luHFTfoHgu2vuUard9TXU+GnSmiikJ9U4gDYU4tOXtKCK3wFgDuw
Z/syxo1toCuR+hsu74DAxXiZ+GNS7u0dRAH0uke0rvR0HvTiGFqYFDAAa1ng2til
v2Gyp/DnL/gK4R/qjq8iiT+C0+xxjZspTOaL6rgFMBMxBFf+ZNccDqPIPLWbgpyn
v8dYGODbkp+Dms7PaMIwZ+RoEHlP6GP8ayT/MafXr8NpmAU67xwbaKYfEfBAZSF2
VmdbDZIoUpnvkbaYCNMFYuIkw2+VJc4mV+MO/JGYWL/Ui4EeZqqAWgGN7YWLhv2A
VHKsFMGTR+L9kz2YUBJdQl9kW9pwzAiBFJiP4LYjYVuFT71OvSorH2dYy9avIfMV
wQmOYD4BHUY7oVK1Zh/2vaN5Z+pKf4chg3icyIkC2ebwEKLKds7AVbT+ebjQJ5M2
VgGZ015+X70C6I0Zch29nhkwEAZS0Si2pqHewce2zMR5lASljCu3TG4IR/I2ULML
pwQeyxcIt9zqNMrLSWa7kUW+GHpY7wdPSxI3yMeNfrVFOSyy/hP6ibj2Nr2wS0n+
7GM8z1XVsHYCBoA3FdMWQ9TmYzMsGss+DqWJNObOCyEL6NuHjQnh70IH+xIWZ7xz
E/9mHavHO+802l3apPdytcK0H4jfpPx+0SuSikOfwnweL7LxgONo3IoD43WBEbP2
v+Ghg1DdyMBsebTOL8ibdqPNracycGXOI2Pkt6JWFDtpIcURxTXTO7MCxbNAG5bb
wXMyj42TQJVgAOFqm6KtY1qFlY1SL48o8J3z7Mo33WieMHleX0YUJBy2YT0ga9i+
tdgkyU/aEzGmXb9+KGrmPi8Nm+VzzJ+OmsGHlTbMRh5li2y3xAs2Vy3gHq8a3n2Z
fNfE1oBzNY3JpEe1O9fRHUEbQWqniyO0aoJdfvRV6uZYJwW+WxjZcyfw4D08Gqpf
fSbpd5O6XyI2dRFyQK7k07mCTfVQH8j9pTsGr+GZlHuYkRt635A/stqwvbJcufpN
Gks4OeBhurYhMJ8AYUZuU6lbrTqusU6uzlY0La5cOVCTE63Wq/VpTByCGqQLn1uP
wAptnsOIy3ByDdTeTwgOu82rhFBJvlx4vHfq5Wbu7uXWWfkEUFwvekF3N7sp/Ppq
eDybxnPGG1rEJX96Nkub9x9RjGTJqx7ywqiZl37cdFesH0YEOWgcmyyH+hY5tQRL
nhR6HGKQueu7J5SJR+7FHHmHnz7Gi9cNm3tIA2FymW1t8A9zQWwpK2ffYtMd0o9p
jqB+4GUGibOH+3sCzpfFsZCHIKIig2bp0H3/7V0W4B2Tqlh+4RGXpxCefIzwsyex
Ye/KlTCRubDPiOUfWuGbkXsE6craizvNWpkbWC+u8DR8X8MBaVi3ai9Yfeg2Z0pE
afkxKgBwgr0zsBnWaCAIQY56TgoK6aMMYdtBg8+b8u3k7sdOCtRUKnhea8GbKZPq
d5K+HhHfwfF7jYkVThbBB0UHmE3unjbYa56zEso7KhfJMKs+XsIvDZ2wUAA/U4Uv
NqdRk4/nxlMLaSfkopNIgzUD+ZOCdJhQ98EF0l/sMmRjw7BW8Wbv09W9ciT9Lv+t
n9RhkeHGnaIy2uxztusJg38NLStFu9w43HC06Pe6hYM2T2HU/T8B/v8LtpSnsgoA
nTz+QoWNhtTJ0JyuOa7Eh1j1CujJIPxf4OM0pgRe2S6s9BR74n1iMJF3qzG7gokf
a+xW2OQTSyWh4VZDyRO3fD/IOxOc4UpYqS71S0SwQn7IeEZI1/MJyCOrAY+E4D4K
p+DBrbq64OfPoaTH9jlCDMDDmBX4QKQaW6W4UpStITQl8CYUUFOnryfZOEsXGhkV
4AXC9cJ5rZbM3KWB8F4vAJhkzL89ShWtv0+Fnr24SDUaGVggVYXzIevV8b7RFilh
XJfSIqSRXdZUjrSOrCrx1djYUti5dMrSfaxpJS5huD27eicpuAcKRPCjW/WZyOEN
Hh6ecGMpDuQA8pamTgJxfEkSTT0S09dCvQBghrnzOhf9Z1+kkxE8YaLjuu4ObnNe
tVhjjmQLh5Fsyd3uh3SykWYbEEqmah2Uud9CwqyC3P+5uNrjvXz/z6LMQnA3jFi+
JsEYZgM6gg3ch90sjDFcNSRzYbktjoLqVeIohqrhVtDIsRAeMR0uEbixgmhGajvk
l4Wp+gTVyye31uwjlrUdb+iYiUDuk7HCWr7lYi/xUZB+yH8yHEOKItA35nEj3eBa
B/O8K/HcUcpKe9wJWpeFcSQjMyf9Gm2OQg9Gb9chYTV8hpfq7g9wMcmNpLOk0TYh
+8XIcgFFApM/Mvl94tcdX6Af5qWA97KISYo46zJ+r4MZ+AmB24+z/rdcfaJK/u/i
iiIm9u0QakuGNz3f0KXJf5mSeP24OUO3Wh7t146CMx2B+XHXhjS1ZwQQIPEyc9xL
TL0JZueMvzzMIdLkWMSI+EfUEYHZ2Tf6T/YA/yX72HBJNmSK1KkOjVGLU2VxnELV
4TYonW4/2XH9Kp8kO4NP05jyi/ZcnP8TBNuubxZdx67ClRGL2BewZMFwVDUn0R7M
/R6GGmUyeFPDjS8FJmBunonC6U7AB1k6tyVAy4jVMhKJWFXC+tNfR6tZnpgsJ1LI
vsS/i11vsH8E7FIMeq8iELoYw2gBSDEnJjXecHmtDiOFLdPk4P/IrAly22GCPdL4
cLbaj+qTd/bK09a/zdjLvnISE5V+xwAlY+qS09T4BmTZTY+aI/rCtBlSb6nL3Z0e
lBcdnD8SFMYgTqg47Ms00SkwWcE1pnYcBH65KuLQ3HBxw+3IT/ZqeTNwGTebRxrN
ddPW1A/27C9NwiITQM82NARwbNooJfB+v0lJQ85d1Q8GWSQlIC/OwaRyvb/Z89qz
4vGtCXMki+kltKVs1i5SzuTSlLvfyWZFTLDR6hZxqx5e1GvMPVVF4nSjz36Ivz/W
0Tx92q+rttgZBr0qDvJu6C88tCzWMTZMYoVGdK3unO/tJ/KcEVK3Z9VXYAOlYR10
+rfpT8UwXEVZEje8sYoHBT+WNufxewvnQ6d1kX+vsbCBDDLCbxXYdOmG8ue49fLC
HSwegBMgPJZbLj7P91HOivTBWWXR5Lvzt4DKn4GvomskNurldJWNM/LmABJ/VEm4
01nIjvcCK87qKpY1U2SNKvY7C3Ccl7Hwx/gFlCYhBBStJ2DS5ByTekou04H45i2d
ESEj3vokO3bVHZNhzeqguq/CBcIrStpH303uHjXJNISLLw+ZQ4YK50i94M6uT9sN
ki8WXEdE6m1CWa8WPKRQ4YR+S6Ybom/uGqRKs4vyqAQJGKz0OLkQY4sNaSNAu3tr
YkdMLKVOF7VrS47Mr2loBnBl5H8czNAxkDMPA7ZDqbIqks9M/B1Gro01VhSopm9U
fXhX7bp3oy2VPy7GDxXmOtC6Ub7E2GyA5zn84jgyNligYhNngMfX3wpUv2WoEmSt
nEPQ9WPwTNIeaoGmYnpcpHTu+ydtOCZfegbjQR6qcQnG79YCl6avG4RzsLV3DGPt
7O2P6cSQE7p6Iw0fYciMhQkhL6KhuaKAQPWsKOWrQvrPZyo4Lidn+yPPjigTqw5O
hNEbNEQYLDldJme3e7juChX93daD4awQVIO0EClmVG1yTVCqhX2qZCy3YIqch8N0
mfYgDd5nDwB5SSr2a1AAa2uK+NR6Dlv3CVgDgMnf4f5QF02SRe2MfFDCnlqglLQe
b7HR+ObMglevUP0gFILMaTmSvwDu3c57RDwbHfa9ZMWFgXtQNqZ6moU9zs/JV3Il
yfvJUd8IDceL8KU3z9dgSnG17/gL1/gAy5Kzl1BLd8VC9mwm3KRcdKQGYICPZdCJ
YaWbStEAbd4wV3x2CHAg1QPtireBrWKp65XklsFFSpx1CKqPcfdekfdxnxxwNeiT
W6eGQRE35gH36YGS1ZkgZx9Wp0y/PEyR3vvN8yfVuWgHrI6m80XdtflnxSLoZaiJ
+zjZYBEeS1GS0MmaR6n4Abgoikdj7ybxomuE0afoHqUHJw3umsGtTpNbpFXo46Tk
gmmj+xhNbAOgpHgqolXnYCja7/XLrcA9OfvSEN69aJBReExOPXUneuowK3u6oaov
M+MhOZ90EiI4b5rERmUbBwgGXl/Y7trJ6elGsGonzx0tfXVagmM+I0urcyzNm44O
tccrUf9AtmuIkN0KfFo42Ogc7TEmcNTMt69umlgme5FgjjZW3qu95/zJqJoGF6fO
UKztZ16caGhdSp21pW6YeyetAffjbOYoC5uliz2C5H3zwoqacAvZAkW1+IgXUmZz
1mfPlBAxYGDLA1XSZ4G1jrtlahcLRPT2tmzrj3crVe+Pv07IozmmXBHno3LSafsS
s1w8n4nqF++c/x4s1G2lzyqlMF9I37w+O2hS44QMrMHY/Pqt39efiQ+/rUf8454z
L7hCx55DJ0GpSL7JWU+lUnGirAonIxUui82gh4cqNkABC5ykDRzamTidBGEDxcOE
2PJAsLH3Y0xrfiuF2oxHIU/WGV420sheS9A4lpt8uxrBNRw6o5efz6VNVAYsBcg0
yl7IoOTMca5jaao6ewKMQARZBEqo8NCxsyYKRi3Y/HGDlN9hFxguXNRWsBAB/Ex7
U+ASyjZa95MF8Og881foi8M2C9x5CPQXG8LACHQkWT9P/DlHHOroT7TeI4pIujLg
8hYsVtDM0EyIeGpYj2OB4XZrOuFerr29Lea6ICqklyAylGyxeL9f02w4jttMhta9
zDra7pZiLtyGiJTweV8pdsaNgxGXBVa1upTFiofw80wE0OC/w4A3Sk4/luHwxqyW
3axW1efpsN7jXLtKzbshE6QY1zYzoMMU/dLSeQ+zmLqNlm6hUIJ2ilQi1IIyIzDA
yhVXqbkarS6U6KSirFc4ZRCbcXdapLrnqIbTG+UcZBt72PV3W5mbvwZqIVIKdVM+
cvLC+aL3hTaCP+ZqoBrTUTMt8n2dgXg40p381UeVuSMzAn8wa6n8HPpnmI/APSBT
EjyXPw16VzvO4UYp5pynj2zcNKbyCcev39BKV6G0rHp1Zi6tT9+DSTkeiJMrXz4P
rwNqMM4TRBRnfrwN3Z46cPJgycy6mGZaa5WN178Km/Igo1ZR4nvrV3tpxwgNu/cx
8Zu41Wpq6xgq0V47zJB1jN9zlo+EEibouBXn7BqJHKxzKeU98Yyr4IMPkTkdDpk5
B8YDgqTKNhqNVYfPCOg6Enhyenma0V6XR6BKIFXg/EevPKooj3ENBFwyxFDbPaCI
4JtzzazCDrmdNxuYFXnJAL04FCJgH561uWIbaqPqQH3KJU6+iZHZKFqGwU7Aahrp
D27Beivt49Fg3p5WAnbmKCcWkYA+WRqQSQgQJxLN71ZiYXlJjrYA08pMIl7+e/Uq
p64sdD4lOGtMuzXI2oo6BqHkkY+Eps2CiEumo3iupawbiTf8YTZ7xMKVvuYq6ri3
qICY1YgMT2iR4N5Ui8spMeqn0CGOTCmCYyZMHeh8hai1WUuHeWtuyJffrdiNsc/H
zO03bY9CUF+WISUwtGqca7fmTGMu1uhcgqQJVvha63dQuXlG8zZrrRhZmqNczTZq
A20dA3sP1RNqeAmxntQGD0RzeVQrGSseDN90lRziGnxafo6hj1zO2Vq3AafJtMHX
RGuwcCChhYvwG4+JHBrY76sVe3+wfm2rt3ew5/Cm44I66f5fBHUIOTQV9boaeDvy
ieDOkm2V1aMMOyGP/hZhwmM3rrfHVWbkeg6qvgXvZhP6MjB8y++BwtRhipMZFb5k
JHYZ267xRrXkkuAdHkRD1xkGVCeC4gPU+rnfhf7uAkfRfmf73LtP87t0pYnGrCyr
0NhYJiqDGj1W7EG1VD7+8OTUULIeR/ZtTLdhuIdYDZFdfGCGilS2cWC1dysjUT+F
UtTy5MdTFX+L4efWzT4rIsVS8PtrhyCOVNLYmSDwQQphBO1P6XDr7NeZ1KtC7oun
6mTBHhEUgYREZXIuOn1vsYOkW2s8+F4EQ4bHlD2zIdWUpBLU0xZ0QW6WSR9i47cD
UfwPXLh7+vXYsa9NzVKyjjV6fIyy9zXZDHfzeu8fPiBBp7Qpd/r2ikNExDn9FViB
cpf6x/PJnZJ7ymDt+LJU4JszSFid0/fhaMfdz+kGt0hhZH9s5jLAWvWQvUWOUgPp
CaYRggzAuGwLr4dGUlzFNV8FwJWKzXHBes7VNlCxrwgWaVLTvzNcjDmye6l4dSBO
7jfjxmWlZ0Dj56kE5yFZJ4sxkyCtfwZW8kE4AEkAin1bPeSnNOPOrh5Bh++P3WHK
/OAYR3L7TGW8EQfUIdWKHdVPGeg3YFVM4227WetKCwrN5hFoEZN7nb2+yhbtEzYs
w/5VSp0LOtd4Tv99kG9eVMdWrXTeDgBB+1RzHLmqGixf5zWuZBQpsOX2pF3kPj9v
DYMlo6Vp7FcHkgYW7t6sXdnkBJmgvQM/WRNiFJiouxpxXqiZ3++MQMTsxtDIOsci
ZvvOIyluciT7P/faCiT8xmNII6iSkLCL3Mec2yTiE5nYgel1LCrHSErzMQW0fiNY
WCylKBzpGZI0iRmdeo0qny3QCCz5l11cUazrOEZPho+1birY2/pYrRS8yEr+rPXO
s2xtkMTlgMhVUe3DR2NEuH4zIrwR16IFXNc1n6DxyI1GnviMHrjDnkEO4QkmfJ6E
gjinZfMslfkvZcgz0Xs7b8evuvz9pvaytqB+tWw9Gb6B4Gl6lUK+SEkuVoM3Wyx/
4Ejqx3Ag1PZ0i5GqVrT4Mkk3HOZcQlwPQ143ZZucOkNvLeUe5QTV1aMOAmVWgyLj
y+YKEXx2YMThPJfp/95poKR/GWEVdR/f55ZsW8rYQKvR479MTft6jmoveO2qP0yi
8dJGn9HOgw6R31FwJ9fEzdPZSMPceq8I9QwkrLzRVDQRqZpcJwta+zq6501lZezj
47fl7TCm2vHO77Tg2PnPAGBj3cYlTpkY09kn6zujoBCL22yWxo3vKqF/AW20WU4X
xb60pqltd6bvGYaNSF3IzMayhtbLeS8xisvA9T10SCI67tvT2IY//HJy+scZnSqJ
vlpOwvMpydYgRsOP1RnS/KDEFb3td31xUUOY4eHurc7tXAg8QV+8wk097GptxSMF
ESW5KUOehmgkyhqUjgXfkczayPbPCyrf92zAUfG0bxVVtFQqAyO/DA/GqVEeLICv
yoEK9uP74Il47LbTf79nq0p5+c9WVlTHvO1lQ+tGLER13RfQnAFygRhmdYOxnTyU
HSk+PXt70yEhIQn2tyx2Rgr1M0nItiiCJmIK0lMqZA/vRNZqQ+jqs3hxAx7OczfM
Y8etU/l2NenpZpBJ3kTAIdSNHPOkufR8RxG2jy2glvw7JqHkwNjaNr0DLmXr3iVe
frCte76txVKGoz8X64sixKujPNIIXjAFy2b8pUmQSi9tUK0KCzWYKHEob1WD+rNJ
YV3Xe6BPd+Z+3FDz3lGLrw8alzkqPRj0l9MUOagsNO/0/Qzi29Rs9+I0AH/kYplk
rTaA0I7NX8hXDXzrX3XzvgbWmoJZe0Yi8YSVXucNWgA84q+WNKFqxNLhGJp/tDBO
y3tUG8wv8eL7x+XBGnmV5xdmb/+w8/T9+OHKr0qqOjyC58g9LQrGyggz1RTH/tuy
Ie+Xqvy9NIu6Vwgr5j/y+d9kQ1SQ6gafCyvKYANQmZUxkuL1nXoQk3x6SZAXZViL
wuRJWsMFBgrLjvYXvTqaFzS7SRS/6uWE8+EcpCFdv1XINi0qKrlqs+XL3rxMqSrq
JwKdAB4JeOKyYE8nxVJnTFbF/BYJadGQ7MIig02v1gtQQXS5TwoHBfUsrIoP+W9j
0CWsMRNMw+2BsyvzwPr4F2EshTW9IQZgNeu0l8tld3myrdWy+C/pMaVkgCbPxrSj
baizWzhd7RSd3uV+xjof0w7yT74P+hQVfEmdPl3LTc+MNjWRIUnDqA8iF2a1DHiq
uvrSPDyPSzif2P/QbwetIt5a/ZoVetLc51a7Nx/PNykY2fIZirknCGSoH9kIbax9
CGsF3ILX74KuGXRuGz1F0tZUZjkMpur8EJ/8QIfDfSYR+cE0o55MhA/BmL+3aZjO
iqN3DfzUvN8RmAql94FlMGWvQvz+8R6nBbu/g5AWqA6FQgOb0gbeIjSgVTBRofsQ
N6QqvCcsQNBfaV9SPrI+wKgxFimlXdFoPZEw1IcJbBPJNpcWMy5t+ENA/3voOH2R
U7L43PxjBPwDbhU9hkZxfzFqnsSFjDg5lUTJg2d6r8O9HVcn7oXWlVtEfZUbwgSd
DjS8SQsUElv9qI8gDlFTl1BOpRp4rUKCI3934/y7MS+SHMT6AUts5cHeklpViPhu
PqpKwLoJw4xw0MPNYacwdtezo2rXUz6xnFrJb4D0ThDkNld/HJk4ypeSZgtmiR6k
erv8BThWR3Ifk5w3DYilWTQPepkfcDW82e1s4qkxy6y8y3VIUFniz3j6+jC563uD
fqSTlQFo0pp0K711uA+s86oVlOdOo504cjQcWSLjT9brHS+JobuoYND6/OcXsh9b
FzFQFaRAromwdHXbbePSNkXuqMEywU49GnEyW4sRodxo0sSKEFXUr/t/0I8R/4Iq
zt5yBrz4MhFmSmw7Wz0/zjQcGKygzhDK9Q9l1ECMCU1L1Olsm0QUdftSQr1CHOPk
f1CAhTmdJ37HW4GRIXmGOrUXKAF0b8oTka/5ljfJs5zjI3FJy3ckVyk5ogV72BI1
WvLYh9FsmRZyS3Mk9t2vdFz4/hJ1XaC2y5+uMMCJYJP6q8ViWlPGfrLo0tQ/NxGM
xlKYF31ZZHyXpjowmZ7I1yQlgceLhVBazOIOupCLii2tGUgwkVv71B8vBCrIrKNC
Qsdce+qtLGAl7+Pt+R38CfMOAFqBeePLGneECtdxlud7HTzDRFv2w6dtTZa+34pW
bGDkFv08VY/xgoxY2kO4sliMXhevZcnV8jzlyU34uM/axkksp/hbN+NxitdaDnH9
K/OyyqrOx5hS7wN91tFEWmDppDLMmjOj3CsNVZMGlSreYhGNzYYbGnKVW+7ZdLEX
X/76X83YyZUbKFeQngNYTVXWfqtaPtsViIVNEiz/82DPtxpv88jVgHdhZ7YF5YUZ
mLj32SVpRTDHN02N4jrrToXDL9FdbWE7BqIT4Imi4BD5AnAjJQmObszo5DDSrkjG
6Man941gMrUkJmfHfbcJXBeUjtMGmmu8cIDSStfZjEBrEkW5J3a1Izeistch6xJK
585zdwPT+t2Y9hSAKtDuwoPYa+RaU/BJNago8YvvkdVJ4qluS5nEP7gig/TekGvg
QwsT82eX+NOxHw/kAc5AHLxX78P3XsKry0XAWWMbbOINiop06Thl6QYYsnHwFx0c
H24Kg/yabl+mTmgmlFoCY4Oa6pDc+JzQeJNLlZeRsVlolDn1e7RrGZHk+9XpH+gl
bL+Cr6D1GzQmXlSFaR70zx945CwkY7V1Z1bfeI3hGgD694dT1wM8adQjw9YTHPax
GtsSnPQ1ocb0WDuWB3gQn2jjfOIaQy/uIxd5E8PToWG4HYfUre6n1HWVrfW+4T3r
tJsIdoh0HNmZI6csuEHhGgn/utSxlk4S6Y19re+gkOSVP6AKwF+ZEKa7U9vMHGkz
q5pBU7Hg0+TkLmgfqijKJF4JrNArQrVve+yRaa+4yjxFPthk+/mClX7IbwUZk3fl
gm4K2R+JMFPaVEl38ixjUiUbp3jYjExXbbLR5tdtkcuN6X1daWM31NK1M9np6aa3
IY5q5RGv3OScSVmfGoQhsCX+g4Gx8HvSdQJql2tI3nW7pjstwl7sunb8LBrH3QFJ
G+udEtpOk6+zU+oDXV8jZ1+xPVNqHQ/e7LAgWNj+EXLcITLi1x4MUp1/bDQdhOPw
UTgrYmkf5nzNcAU8fxrnwH1O/A6qCoU00gGb+uxTNSMJiEwuDZZz08TyLSUMUMNI
6cDAqXzlTjeRvhUGBljccOiYuEZEU4HueDh2hu02glx9oygjVVBD+SZMvDJmzVoP
V1OEEzbTIPdLkPmsVbg9uVnVJzbWTJDGfT0tMQu49iVeXTGUNNLptfer4LLc/nru
bsxctKufYfSJyc8qUR0QVIbJckICAUADeZItKKxIeDg9RAiyLw2TUYn5aqoCV6yW
f6JGppf9PEtu0ds6NE7p2Gfi38CGw0aIB/zuu1SchLiP/Km+XaRtC6YQrub3L4lA
qgnK0mtG+exZ+BRmApo7saLhWWXbFh4dceTLkg2+n5UE9Sr6YeSVMcUc8DmIQF2p
ALv+JaV825K9m8juZn28uyBLD5R6b9ccDCjLie4+JPii6QQxqdIxwkK7W8nOERLr
TyaOALlGc0Ff9EFN+JZUNans4bHYviYBCX/jH53LBxgeDHIuaPGDEOIlWegfLOSL
ViALxEZNEeY6+DNq1XyFF0+a8b76gZHfTJCFwTwiurzQjcQkqkASDi+Wgxggj7zj
NyxRrddq8tty97fBU4SgI24TX6yVPSEzham0uAZEtVsk81Y+y+v+YiUpT7+voT8S
B8kbiwzuxOnLBgE2f7cx0qEmpHS3fek4wdoMDL2jRYUPjxiYHpIQp8zI1fpVQrNK
CLD74kbL7Bb/G78mRbrX8V73iw7S5NfDxj0t2IaoAzWhPoIuLe8KibxcHsDE7y1c
iN+ngJeV+SBoRQHxoFQWqHhbPol5MpSYlm54YBS5cNef8o9izEdYi14he8GWXAHO
/n2f9+PB3XP0pRjmOuXlDZjcgXFqBYkXjsOX3iHmACQXZgzrP+Ja0XHhQFQ9GuAn
sAFMoGIdDaqW4hy9J+jCSOoiNc0XdscLkUaHT9TV3OzZ61ku+UMTOoVhu1i6Kw4t
veJLyuNXp7yeix9X9tg26j80aRnElG0o48dJdJdQ/0PZvEnowmP7dgXaikB26Mhr
AMhfBwFH9rqbqK3imx0iUiCWKJT63BWA4IaGPSKCIm44G1IytyNUdt3VFe7zZwK5
U0hBCGdEXOyrUWBUS/hwneRvapNHcRiKP/u7D0pal7MVJVJo8YC/kKScmOa1pl9O
76GfgA28mt+w1QWFoV1pKDXYJVYg3CNts+jdItZ0bBRAz8Nrh3GfQkUjmjE4R+nT
q0010+FNt1qnxAtQ9wiGKy59mlSwxCAGvxCsG8KsxEACyx3W7L61kI5fdWxoC6IB
NWNOvWjxJZ63zaSaft8AN0yZEpSf3PCZhCgERpsrf2Ejntc10XFlg+gEaMvBhWVi
OS+8vrlALUluaZjo9nD5UJKDBARmIagWWxTsebCUUtRa8VQq5zK52Rv2Tvx2d/u6
ZVM2gLJEYhwAuuFgMvuNjpk5IjgOXmA+h1yx4EREofMUSpTdcs/vz9lU5XxinSOX
hA9KkeQ3UdbOYtvoZ8OGw/cugtNZL3057SPSrBg802Z7MzB+iznqhJpgM9N2k3Rd
yW9QDjCf9o5MGzXfoT3H6M9XVSsnJyFzVvK6zAVKHvoBhkVlUMSCCWgS6fDoABjI
MZVZ4aXZHZFEKRincE22HUKyhSM2taui0YPJJWL8yuxNzObeQGeW1xoBlrVg+jDS
PEZTgQxqO9i+dbdBNUcmOcdcJ4QdHV5btjKmrpwO8PkbnP/yKShj3k81ctNZFMla
ou292MUSm6FxLWB9b4f49fDrfzSAfZIS7KUqY/VpFAQUdvPFy61Jn1SREr9Not6b
SyrshYja46m8g5iS9qa3csBZ7JdAGVpNB3gmlD/TgW9AJrCA/jK200v7JAZAgJAd
DfHiA5ltmQMHwEk5I2CdepW98Zh0Y8+49NVkCJA9isAxHzy2bNwPnmU528qw3EC9
C1YPkmDBOrsyg4XhlMPZ072eHEMQp91S5YElRyP0DLjEDHm8/pAEICCkkfK6w8lB
+c7Ih8xeWSBuzQM4qBvMj+JPSnh4fFmlUt7f6/CjKkUNjBVWxVz2DcsEH35Hj189
3bkTrPzTxwF7OPFiqy+fR8AgkqzkrIk4Yahix8xT9AVaPaiebJWyT4tVFnUvJ2F6
ET1yJKFblXKI+h60fGoVPW3dNqok/Gt7plxceR2XOgPaKyiHQzGAzs/UazzvTvVe
6PfW3hGsw0KbqED/TlHt+uXUnCA4hZda1/PEhRv5s8B3xous4Dj8SmxKlE4DtStT
SU8OyQ8LosAvPzVnhCnO+LEHSTuUNpyoSgqmqKeAfNiTzQ0/3kambDVMUDA244kp
6ObwTZo8Vkh/l9a/+nB/R+n1yS2N/wmL+4kmNM5R5/xHYIQnCkvEIkDjkcqe6FjJ
yzEns77dNyaiV4aUu8/xJ1+n1IzgCk+m8rXbrq4sYRkoORmEOyUUEwergEvJ1Jhn
Z1uA+rhkjEjnEcWPvA/4cqfqi0hK9wV2XcJ1rEfHw2205OVA3Xkom4PQQkcqFcL7
/TKL+zE7/LObBQapck0OZDjjvssZwbMFrAzFoJtq+VHG8Dy8Ba2gK+1jpyHtPob1
xeYa/E6acnKzv1pyU2EL0LRbI/U+e8OZhUNn+jy61j01BGm9HYOfoliNJKyMW17c
pSPtYGvodU4Q4CFWuJ8EBfvuautbociq4a/rB3IakYE2HtjivbWupvzzorGZrfa1
t7g421wO9jj6Ifvp6e2dY2IVPDi+z2bPgrg8eRXkALkwNA4lTznQU7oD9sG3gRPz
6rWcE+3KUWzWGVOKhF+OJJYNDO9+fT0uCvEdjsQbFaTIBF44zaY9SPycUz5XTNgT
9bi3MBcDAOvgC1DXmwX5DH4GfQkp+kpOH7PKuqGizn8ObYL3kIqC8fX9Q4f6UqL9
k9UJav0OZr72Bz5otOA5ekSytn+kgbSaoiO1RJhBsl0OhuhAs6pRSu/zRn+Q1mV7
FJ+Lu63oHRuZREgzJBnBTSaLSmVGa7W/ToiRQHUslgqycQPyzfmSnqia7LDZCCUs
GQd1rzP3nBJLXjGSEitGDN/YlakPpqszUmtwFkk+kT0drx8J2SrNnyiwQnmhzd/z
nODk9nwZSY7QP+hx0hX+a4B8WhfdON26pZxQccpmFtkyxFCwg40qaYv1EVava0OS
pN1fjg/EGAXJjR08oy0fpM1JjVQkOsOWmD0yNr9hWa4vOV3rOryEzUUytwEROHw0
GwLmYtrlkcmaI/xW/hNNPiR+J0Ivd3QnrpiR0+wDFkZk87aVcizys43L/P4JeV/y
UoiR0Yd/zdaPNCcE+puB5r0CfAN2hI7/mUcJBopd6VfX48jZUNv9FHkpFE3rUCja
D9BvHXyJXSHpi0f1EgTY02FSe6cSeOjCbcsccW8YUR/IuQT2e5s4apV4Ib8agFOz
aez/EcHFL8N2Sdm3ifjl2PSe1jJxzYx0weyxRZagiNsBlzvw25EhS9axFTsiRLV/
fdz4thGSNbkKCKRmOhj5ay6IKv/UwwQE4DVqhNlUmAszzp8pm2XJ5G/x29IpC5VN
NM62VVLYQu4/XvFwM4d5/+PPYLfdsqFPelTG4CVmBFg7Z20fjPIzMPfN2upuaDYX
Om32eCZq1WFfI08P9vi/+RI53MnQsQzbz9WTrfSc02RH3JKEpfR7033cufjtHfXc
ZZIm3qj+a0T6/JCaRvO9WPu3jNmB+6BXrG+kfsqVgx0cAISrHrAXv83IO4Y1s4+s
1lUYNwLURp+aACeqBuC+swH7+xFyqPnbKbve9G94GLFBnGetq6FQpONDoqgrUuXk
Bg3QlCcQTE6VGuwU+26j7BVZQJLjiUqx137K5Va3rsauI+dlCWUjNz633G8X5lpL
6rPCHzUO7h4Z7UrxOonui46vXi6oxMZRB4KjGJdu5UWV0cKtcopKiAeg4oNHUoTX
cIahKmHysmi8OC6aERjOcW4Roxfy2k0IrKvM1mje86EqoDDPT/3O8lg0aO8YwSli
Xg4QQAZGI9YIU9iH2+T8XT6Kwep9yYdFlwtPs6TJyjyOWFkaLf32um8NFWDtVvtx
yWB5VuLIMLPtBSHUiH00pPLT7lAvb2J6znNDiP/cwnYn4xJEM8kq1Xj4gFEcmacM
cndcrh2fydY/AB045kfKvDPt0JJwIMg02Jl1YakIYEMzGGbhuWvJ4SXEqJ5KFeOl
EE5k9VF8UcN0IC08JaTocBrqXk8IDGcQ/3FdkvEqERyY9R2ErMfqT21WiXzUJgN/
gNg0G1gmgbJpRYhsKDSPvs62qqBdFyY+yKxXLa4NIV1YqlhunJlHko3K2jjFvgzk
B5Nj1QUxPaNc91meiVFy7WaT5kZhOuunbmiSprtgABtOoLXcGRgTaYgvzcoi/E32
tQfbv74FJP16gH9l5Aso7a0aun3WAW2VhMyODnsRCTCqR3Y4vkvg9jQRuLe5Tat5
ljr3D2NpsJZJQgbpo78nHbyI1lDgR5xGklNzf3XTsw8jDoujzj4Vk2yXk54Zsnbc
Yay1EV8uQf1JMHBuN1VONiHZmcmou85/s70Wl00LqvB2+kDzKrK5vFyM4DbVuhOh
puWbDCdVqx3FjqLmJC52rNn56QFS0ymKd60HmW+FK+A2pUeNGA/WOAgIA3wucfYq
aKDL1V/ZwkTsyyybDefr7xe4Hn6n0WOJw2ytz2AEqHDXpKJiY6+TfBPVuPg5LW0K
S5RoZOmrk1lIcHXkp00rvPo36HZtoef6B5Qam/oKNNCUZLHbI8JeubrfZAYlpoMY
kyJxQZNOlmZpXHxgymQEqmrBoCEsUyq52LB7IIjkdkSIxk4vrACG9oPZsZMvyybi
cAxUg+IP7LLr6SSqA5SBAROsIY4mbFbRi6MxA822FJKtQhFo72+XG1uBRMJcQue3
NFL0ErNWVa8agabugwNOUxZNAcdcyYuuVYds1B/ZHEvAFFIc0TQ+liUN1kW5johY
/N/QpArCxDVqvufv33DXHZys33pLl5casJO6fdJtz/T+OyYFbgFDs/3kEFsThY3q
vDB5YktYckWspiu4JAU8fV9Z/+CCHKmKLKV1QfUpguVFaTvXkDa6JpjAyIWwWJgg
4P+Eky+u571IJuwHUTChoAUtGuk/55qUAWoJuY6FrL5qTbiiDk9T0n5h/9PG54Jk
o6YUfoMzpln5Zrnu0dh2qk9ui4ZAX6sXzWdFjM58wD/71j0IftYJ6El+spA30xVu
mu7B51PfNaIs+dKfIuIkV3wgrtww8nHQY4gINUtjWjjS42lLHZ3zTK874SDpApbI
5rcW0DcsXybXRHYVRuRMaSGrOvhQVy456wz5byCNFboXLXAnK0cPFse3rIQzV42n
uJmEDuv/+tuNMrTSbJfKwj+aAJosUtGRqWA2/tI1WR+KeMNPSDymtiOtcvBUj72U
0QYhFi2yZlYgqi42A71m2oLSVgiti8PCChcTFKw2tBZ0X4XGA7jrqrJi0D7zypCA
RhmbvG3C0t4Tqe8iblw+BLmDO49rlx9k+NwwB/FPh62VUDtNCWlG1LOUg5mpucLF
rPJZv7YZ7zYuXHxiKGZLSunfVyINk+zuvxkBvlkdF8ZBO9nYq0ATtTMjg2O5UoR/
aisePZqFIOZSFFnLfiRobnQZMadecz5Smzr54soc6cCIkTCtA4ZfjbJpNxtiDHUZ
JrO1E40CBBWO7RGxdEGYXSA1ZQT42WljFEDFC73Qx06SfqIotyHqThYIsOa2gcN6
k2Cmtv+GkisZrQ9fEAzesaVy8ia8sctDwspnOYDRwKaQ45J0Qo0k2uElYB24ZSjM
LPlLmHzWdxdLJKl8ATRcdR8rkOEVsuqOpOAg5OTBib5JbGcxGIPXCsuRvLjWxxuy
N2rDJxgcrPuiPtcrxDAsl8kB24lrohetjh7wFqWAzKIeN3RTq7voTWxerlTui+et
c2mMmcuN3CL1AINPh04ttblRlBADjhVuFZkhUC8PFOtJAziOVlGJs7x/40i0Jspm
hF2TzHJsMK5DozMkqXWSo+A5XRjZtXKqPpekG3f6GQdweGiGk7powrxbxGGWibmo
uMGGuudNGh5eZZOx/q6yq9I8RcZaEd/xTP+CkS8SIsjw0rsv0sasTztdOsO9tXjc
P72e0a2cVKIa/RYe6db8gy+A9dxPIYQhKuQuUq/fxj80cOHnwjcnDlYmJJ0QauBr
UbG81AYON449kOpo+ShRqbiGktYfe4Pdu/IFiBd1bW3amiOAmByZmlbTdeV9LLOi
JAnFIVF2p28LvHMN4C2wHwmWpGpBSyT12mWhkaUHPU/E41mK/SBOLmW+wScxvW3E
omxnFvGh13SATdxS5lmwHnHl40sUuq52WGjXLAOdGBKtpUovOx361S2oFqZtGWWX
Wethh++0Ey3XnwF2rvje0F5/CchnjbCdQPAxFKOQejc2er1UcjiD+TmEBtIzJmG2
XS2TaQHVA6+OWqy5H9ASz6JzkZNVLeFVGIj4InxW660TnbXNByjBJt0Ho564bk7v
lWOdwuevh1nrEmsmzNUjnbp9nXDl8BKm2+yaiBfWpDCL127M99InpubJvJqsRy7R
kjxchjwqSx00o1Gnr1xSVFdq3zpVWJVhlbD75rW2U9P/SBWlILTGYJ0nugnVjlTZ
iq7df+rWyVP7cfjgJA7qwMnDs2xgfUCDxxZcPYvI/Eg9yv+DNpfVjmHH9UeB/Y9q
zizxZP8N6MF3pG9YXCtady+wo6DUHu9IkyneKJY5lkSxZJPcUskk3SRoEbcrDlhB
/qnorf3kwzzHn3c9GwPaQjYbf89D+fA4XSpFPVU8GlXYiawzlqiyFMaLDOUubG8p
NGOfGxiLOxlJmgXaCXTmrjkRd1U0LZdN2VK3uydun5nTL8Ies5Srzc736o/mC+tb
MRM6brScORQ/MwC+pVSJCgKfV+FhNhweWE9L57dFUnlgm6pvmtAXzsMNCivh5nmz
UNa3r/XYey5lzb5Tm8s64AFBWPmEo2+YJg+1PyNMymVrCd/kXYQkQnpZLR/MI3EP
AEbIOYNh3WVhAdcTPh/V+klFY4gWwOh2CfBOv/+XxMY3HNRGDllg6uSXdygiO1E4
Wlv8TdLhD9VMwdGOxPfCiYxinlIZWThBvm8dPbkhEZTYXiF44r3SN933FwhmrZ5W
PdIuhwixj9x5MI4AjBpjm8taZZ2M1FnVZRLHQg+c8GrABJWWPNLPQph6rmQn1kW/
Lksz6RO8VXX+nCK2//x76bfQVMUIhXPlzZBaEn9OKeUONB1Iqh3yb4qmgUTKRWdS
tg0AGo679zT0fLUhKJvoNwF3lbX8MD9hESfgPE+vBdz+Rnt8L0iQYVv0zwaCBil2
OUSKPNihEtfHmeb9YIBTw+BNp83Yf8pusR8VAMjqmIV/vPmurUqT9RyVYIkyczMZ
EBsjsy5ceNZE8V6verdnJuS2qpNKhPw5bqzLXAxbEh533EFKng3zC9OeqSABES+j
gs4BqpwTZQ68BsEXIIN3FX1TTwH6wr7mFWuLW+R4Du8UHSvk1hvc5SSJhQoLOsXA
VaUYuNIelvd7t694l0wMTEthI7i/xbTBieOZEDBK1jbWw1A90EvIRAoDBwZRQeFQ
9GQ0RnBMLX0XcAu7Vspt7uOtgLr+edNCbuAy9OYydOoRn6TMuQda4tjmJtEN2PY3
mltet0F5N1BW5DilpAssBs+eB1QA6+OdwcyVwF65YRJHxr9n49kvq/EddBjl5DrQ
dG2jqB3PFo1mUfMCQ5Irl5fC10JEl9qDi8EAQV//veMNhaOmryFdp3mJw3kL2E8B
pbztUABtfoJ4fB7YkMUuaD4v/SduIqJdR9i1Wf2KL8YIn0umqDNLfVhOmduYy8WG
f6qR/seXCbANNzPFN5m+y2H+ftBPEijI6AXDoEC8okbcwLR/QTh32cvQy1WHbBmA
JjiWXPvr+hScToHJ4ExkMYdrIRpMPKKww21g7kohq+KucWCsBhdm69xf3v++3rOl
x8lny2Z8ekKMEUL226OSS5vbBBztjMJG4eVN3N2ddcbUAe1UPyVtXFooW93bBsoy
JPdR3i//v3Egktfia3OL1M8CzM7SIA4xuEiGGFTyjvQv1qdPYsdgNFAXpeLsqUpu
pIIgOBX4VWfinBqj08WhSlwDUnG8HwJD1l4nK8e84OnND07HiyS8NxG3WIW/uaRU
3iHLCScjKl/3yce0bjrf9w6H4H+EJdUfNc4bW9ZQh/QhJHo5Ov9Ks6UeEBsRQDuj
xNoviWeZL7Acy1exLK4kAnATlCVUkkmLBzbev0Xttpk1pyB2YYW0HLv9qN3jTRZw
NtkfshhIfZKJnelFTTbLiET4crsWWKlmmNZ5ZZdi7al37u5EBK3koWD5auT4fuCC
XrYYpvTIN9M9A/QmlvRaAC4kq9ihad9XVuTWJH7PjXxE/FucEtrALlp+zENQapP9
P5OdGSATntmGJgHqEUU+c1zDCukfw748Yghy4SX2kRspyL6h32TN13//D5iolGTV
sco49an6MEXy5eSwsk/XVkH0i/kTd/at9Bt22TjRnFtY91xU2js/Zn7DUOCTqaJ3
BZuOF5vRd1x1BybmkoD9+sEuIiLVSO4mcaSyAoYItS+ah5jNGLy/ErAMY9O0Nll6
NasCUN0feSvmLrvnuK5BQWBd0vg9sObg9HU7GPuRotHm36X0ptG59fPC+T2s31MN
2nTpdoxB87ha0TOPC35UnaFeDP5Gqh7LPWvp+dUy9ZfaAyUhISmcRAlAae5CIbkK
00yUhrLMGFYzADLo3WjsFKdZhNaZZKBPZu7Hf2FUXN1gdUfpJN5aU+sdfws9gJR4
Xw7Uz3PNWmjgMr1DKV5FMwnPoZR5yF0zpP4KguAlv+f+mUOPF57BPEXHzk3pZanZ
hmToj2shugzZOGSNXWT1Uy82SxyEr2f7UCAQV/vO4bgawLWdywfrgIPYWhc8Htdd
TmTGqZcZYUjnuRbe+T0vPfqKSltHuJRmga5dCsicPxFeCSo4mz9H+nzQe7cS1Udb
SVPPAKcIevrYSWyfqqpsTF/24nvp9yHUyXofenFcAVRukxNGyXXSgWhBQ3hCB9KL
l/57TJk63PLTfoVI8a3hQ51gk7UKBXrqW5mppxTYBC62SDH0iXCb5vK8oiFA6azY
XxFfidLaMR1sCHb0mWRGhy8dHFzAHGbXUhoOQkJ4hnRhwJacDgJ0DtDgGqbkd1Ts
Ot9+ASUH9pqeskSBZ+UjWAglyZbfMmf9lGP72K2arP5n4YfYUQCZsZ3jOiL8DlM8
OQz43FBWS+KhRT4mEUxbdhsugUFF5dn+0z5YIQXKXcIhb0oqYPP4VuY9l0ctodzJ
ABeEAcbCdV+M9x4wYDSltTC4aLjsQ3QOPgEPHSzGsurwikBIHCmgpAd2KCSs5kum
bZysr7YdHpGwkLFM1YMUboZMZnVaHG+lY9pyyRDl0ULf2rRuUhZ5PNVw9kMIcOjj
KLImm+RlvexGDqNJ2CI2DrRtmQ2KADaujj0tpgbJ3IbStQ0r3wHkKIExcsE3eTb5
v6fl7Ublh4PsSbTqpec0KlOMfatB/ATK36PXIbUVWBjg+zi2D2Qz3danKEclgQRc
UjrVb++SdTQHkkrmzompc+InM+hYIrjN767hi5/j3SHxFeZ8YLf7UI/dHAlrN0wW
XH1+XQmCILQTwmYz+jutti1vgyCvZ/++5xSY6UCKtD3fAMdMAw5RnJzNs6vgMi5+
mpjt3Yk0u1Gw3galFp7TRHQJmhof/L+g9AH3/aGlakebje2tqPnkyLcabbxliOGd
jDem5AuIJ79IR0RaAq9QmZLns5OXelIyLy99NjKFdbY1BZAGoNFXZ8HX1EwTPUuv
nyuf9v4NKpfYomE5hUpyepLYZRnzpw/ry9OqWWpwHcQOB+bIIV+j2zX3zL5GDU5z
KFbK3d2wuuPny3GOgLowje3hRTEIrodxjlJ8OOCwLrMLy0N21BHhkwEEk5KrvcO4
O9uTTusnstrHKU+xSKL4BFLJI0Wyc1gpsDWzW0+HsppJWthsYrdGeHJmLet4O6f5
e1Pt7AgsZlLn8scrQLrEFvFag2w3o24FqSX7GZYXBlBUMFTGkO1ShITibVfMSN98
MJlJNr2BVcxPnItvVcYw0+AjNAavWxXT2CA33grzzomdNnh38WQT1U6TPvVmoz5F
Uctx+xhcdlrpQfKDo8niblJjHnYTJQCaWtrBC7pWxyeJTekkW73kWurBIxYQRled
4zMVDKAxz6SEr3kRiNLY+g9/7GFlrDhsvjI6qkFvBxZ2eNXrgNhAqfWN8/ZbLRUk
CQszlWa6pCcB/zgn7R1dlf3RHzT0MOfvQKaoQ2ndoBoVjnVtlr1D1ZKFlxTFc0YH
vOrUAr1D/BTMHf9xUCN77+ObhARRniwPr2VQYd/0q4nAjYBpQE7YeS8bkzwm5dYq
0SMzkufcLZREgRnAFqSzyqyfvtkWVzrYPTMKF/oNurOM9VTnfNePb3uX4VVuJ0XZ
a91fWaCh+WW69RfoQWsVAC1KnV8ZTAQqpw/A8PZfR73VgZU0siAUBucy7b4A6MiW
VQrNgUQzWqgYK1dgCaPc/gXax6UEvJNVqjZ/Tpkklipnmp3QuJVS2415PjV2a7Ny
hFc36LIQvTEOvi1dq15GAzFnx/kXwCytk9dMJDGMfwm+j6KvFzpkAT8TW7ryQReS
XAoaz3GHHc8YZIj+jxMTKazxyu9JzDnYv2WBFCZAl7TUMmfBob3Rg3QA7yLLJZpo
V8k2FpEDVIhwahChD7wutYbDBPh1o7Vhz0p0xJ3cGLauma4EB9JbEj+kZrGHr3GJ
RoXME2tsFovs5cHVx/cblgqHn2WE4/dekwlb4oV6OoUFQvQaL6SlHWk5qudhFuEZ
sCaGuyZRzApqxrFwsXoFrukobbm1floN2TyWDkqdZgHOETPo5oih4juhZrN5l3sN
x+zAeKJYevp2ERN7VefZ8gke9NI7ANXgGHz02brSfSEdRE8flLNB27c5PXsM4g05
xIoIFfO08zV6iyECSHYscFyaG1EjlXr4rEBsC17yJXcoPNFMmOJEqsU98Ei2ZEYa
fIptd4FO4hv3gUQ1cc1eul9pMLjn1Yzk6ZKuegjn7kIpn5jiV2ZyJFez8LyypX2S
vKImljcmry8FPgI62UuY63IXseTUhcru6YNl54iCO5CfO8uTBlZDqJHazvzYgWQs
yLuOdo8YXdgJNJbKyHevOKh1NGurlEYnKBafXB9+EzzBhTH+MFMh2f52p2oAPFkX
xanqOmrCmex12L2iNfU4cAUqNqpXGOTLAppYlLlZaC0+XOh6RswElwiYRXxe0JLw
eQptab9sCvs1XlxOgNva9IP1x/S9Enxcu4KMXBhC9UwPU7GvOURRWqMpTVW8FS2l
j0pVyLU7WVuqK1c1BFqJPOOL519MyII6sCDO11+trSmNofOxY2fcodTPPZogo+H/
4Fj4/EnVWBRwVPLfNTr1WApuIYdzGBsbJbK4/cfFjr9bW+JYByytyGtsMW96MSO4
OkefFp8aIPLjhzPHMeJgYR6wJP+2os9R7Lcd9+Kvd70vHnq3VObBULQBm0I01Art
nxJkKF5E5TmvYUUxoWsMLBVlu/b+iqsFQMC7KqxEWFb+0+42KRyUrgp3dp9sy4WS
mEhszM0tqgKv9h0nXG5ZxDd6RW+GKsRUTzC2KTUhNFkJ3IKb8L/K7n38tMdNY4tZ
w5g2JUwPtUjqNSVhby5z4i3h3rdh0TrckNZMlzE53t3laDOfroMztftjFpRm7dW5
+0HFvLg21DZF4CPpnk31/hyiQZgRyfPcOlhqoTQRFkk0+E1GJVyv+8P4T4zYJtXk
T4B+/F6yP37vFdtlNW2Ot49DwQJhwan+akyKTlex97wZ0nJHXURi2oJPdi9PBPtk
UxYnGAdbFOmYaITEQ+VLRBzWZ6e6N+R548MSR5etXT5iOpEfz1Zgq0CdKw6sjm65
p8BomMNnEH8AWLdbmGjR137Bf0qYzgBEagfaU044AG389rdvbziLe4Faj6DhUDri
BDK4JT+VgNPC2F1Qg8a7Voj8YBO78FukZWPUrz2dvzfomef8KJyrRIAhh0SQPVtB
KtzeYWCmnzj6le4q189w/2v0saeoE1j/fd5VsP7b5qK7/kB6V0kr8AC8NMrDwIRH
YbDEib+j0j46yO6Q7/dt94liM9YXf7BYSUmCXnBT3AcnJS7O9329qH4WbpuvrMQs
TiJhV5P8nqwImOYyYGLEN7HhDcuJgQJdoTjOLitQ4o3m73ghgvTcB+pPVJdjGgaE
RvNH8N/Z5M3WhZZ6yMarYuxSt3RmCtNZpTI0NfNI6Zf1YYLj2eoIOOnVomxzbQN3
44U/zvXHs/Gqnhczdy+oAvwz7OJ2XmrzmUHgm4rk7wEuYlJV257f2KHp29ddbuVI
nPMB/cmE+yHpwPutFnngA4FakK6UPRn8m3Y1BDk7vZAga6/l2GaRqYH4ofw5jCN6
9m3xvGPIe7gLYQfhN7hCMR874HPBVuMbtA4Q31R4YkCgdL4np30akSJoC6Rd9Txg
X5NCp7b1qxXMpRwgr0Lr/+EEcA069JLJg4zd2PmYPmuPL1UPCzhQfswS/nfRvPAT
VhgBo3ofkNnsJNbMDCuQjxtihSWR8+tP9ZNd2AC2BsYo6i7yvbDEeqUFWSKw5fWE
j59K1ko5V1Ek1W6POe2Q234OQKXnZc2mlz6mAEd+0VZyVoDhSn+iLdeLb4SWKQ+H
Ofz5o2cltZfK31JfEpbiJxpF99q628JK/IlccEhA3lPswQldQRD3rB1fNEvd0FDG
dszxRmkoirTp1vxhaUY0bJzRtHaX7zJeRnky8qHnTQdJ46imjOyGktZDkR362HW1
gyiOVroBknRxN1gwPDVgayv1gEt5Y0WzAUO43yT3OZKbGQqDkcii0lJtZwSRGR1a
1vnSYKBuWnel8oGxsD7yd29nr9uXhlL7zmxACMr0oeWBDj4pB2WMp5cqOQIEYMtM
8HhIduMe8BAZ4mZhzBT5IFAa+Yn1xQ/OBMxLvccA1zrYjCDplsqM4JLLxyz983EB
x6guTLuV7/YoF5WktwPgy0+yfz93INdVnowb8ztvN57n8E6eOdss6QmaDksC0y+5
iHnPZ6sTtgN7Y4w2kRZJR6u8gZNxkgI7qnRHNowBwUqNvBFA8VNN02Tg0Hr2TjAd
sgG2DlyObDIIU2l7Sf3CRYGvi/x4XLgg8tnhxnLKOvt9vFHOYHc0xXzNbqKgbG9m
63PQTG04FmIKntzwfuzDp++3pj1w62FWH5go44i890WdfM57cNIaBtCO8KqfNgyS
phgRuff6RQMUadAjFPMb9DY93ZnsUZWFSrtqXV9gvomLfhb+5WAB1Qpj9q1E1DcG
UMMVoV6zfUwr8W0N3Essdcww5BOC0jdRxdc3zRUclBiqwqo0T9JoN8DoM8FAIx46
um/+iXktbCgqb0bo37mtaQ0BYps6rcgVih5NRfd7vHup0xzyFwMKGyyj7i3q9Ht+
DIAVS8rPqySR22ZFkasD+mbbid3ITrRNAzoKb3uBD5BZbz1NpVf+pIEXZU4ZT8B3
G5x3aP96aM97J4hVDg2M07e6RrniUQY/BNnlycwU6TSv31NdlzZ8e3vf04igb7m+
1mOttdDKOOIWMgGDpukPEliBTFTf7uGQDeHWZfiKQz9ACoaJgbUw/0QL2b9I2lWX
rNezBdVsaS1EIhgo/s4FtMQsvbqYsSHzIGvaVLsI40UH7n1P7sBtHyH8iC3ChAq7
SPpN8ChNcd9i8KA3963Pjh3NOZfVY6M+0402RUZeDKK2qszmhjozwjDPBZYno+1o
OOWXPYAixv9jCQbgMZmDMpNebytSanFiRHc5wSIolVGHbqiTjoow2lESa2L791eR
Eo+uuZVh6sawU8tbi5SUOQyfHZAo6iNNVo/iq+6xCRfG75MgSWXyYTPcevzkhXND
8574CmDhnxSm6fPowziUzKPr2p9m6R2XGKNaowjCJsPzb4AAXmyRP8q32MDouO1R
f0POjNEKDjE5/TPa36pEcWVUXpBrB/mZrQoK5Z24vMKASHPjMMH/36pgcdbCd0MO
/3Guoxj9ztL1bl2Mz2Kj8bnFT6FV0iFIwICIB9HWLqL8/VBxGdAE/JV1D8ZFjZtB
QxcQPM9vKr6UokZU31bvrb1Zi1H7BmAS01g8XXsIcbY14TrciXPHn9uKuwHVWYw6
zgkM1P23DYlagNRAsEmma/xcnUoT0r/xSEy/yuE/V4J6WCoUxeNCTXjV1Xm6KZkv
1YUOFtc/QtwiIGd6V4AWy38Ph8TRmoQOQsdajeBm7FaDn3Lh/fNQUV/pbhEXnuHW
NROM9Q9rcpmuoOeEgMBCqNDf/LPOrsbtXaZfpICdETGw2MDSK+AYPAzK0KnxLDT5
MJg3ZQxZO/Jz/Pn3M3UTz+lkHvwyQluqLvp0ibUxQnM5IwrEJ86LYSkkB1YwPWJl
tOWlRqbc56mna4cDJFN0LX/Wfn6J24iYzAFN/8dD0wZsVv59ffrw2M5hClHtBMRl
Gq7epXBDJcRnaUm5IkGh+tbR0kToZJ8h3txoLndA+YlCwx2F0cP544KmdDU4KncV
+Fs6B70MzBXhXboXimREc/xbTOpXX02mxq65y8S4oEmQSfh3qKl3WXRscTB1pzGl
0bYGP2sMa95UrLLK6MGRt10SHeX/HSbzJk2mVdrwutxxbG4f7/Y+bxvSV4lierTE
fC+ppG1oI/5hFLu6K41sSEYZu8FmhyQksegCIToTY+HFuH6F9kCeLDsDdMKTXfar
W+D8qUvmjvDd29z9y1FE0OhDwc/mRIyAOpbYHx2dv0bIO57umYLTNGZFQ4kB51Qk
c4iKyrMC6nJqGtvN13+3Lsb+VprOCISgXxziVhr+ehmehQPm3rUIrikNUq2K+e7O
ntZHgmAcibDDaa2S/bYNU62EcWG2WPzFa9X3TQjs9lCMNjn5yPOYnKuBFpPGS3mp
YLR/7vaWOZitvm3K96Keji3W9hDzrcObldilEKmvGipK67lS/FhdgR0/8ZJZxOU0
DsxZWx2hGWRPail7DW8oHpeRMYL0iueZaR5M3+EWnse4sRoAwAcPvwkfCL8Y6DGY
D/6NkcJsM++3hu4uzuvXf8Jd5kDdtw5fu/jStxOEy2Wi5rwkL4Wu0qzGUvqBzGCs
dc2L57uZYML4yPlCXo4jl6Kp6Y6UTd8PGrn+qV2hW+Nb+MGQk8GX0h/X6k5ANwt7
tTUmP7++RAwe7K0hAvx/Qq2iUnBBOCz+WNdKOD2kKLY8sciAauqQJswsNFQoFOMi
X3VzwXy2x0UIY6wTymUsl73mpznRYCyAxyH+qRRDoRb1+5Zz0pRTPXX3C3azkboa
KJ4fPw4vqp7A8nFks3gwZCTUt/po2lrm8eCw6WlZgwlz/83seBDmcJCyW32CdQZu
rFAxKBZ2jI9ikKOoHWCLJ2662ojwIkRfEnDum352q+tfxZ+MiRGuAm3oCTEb66dQ
Ca46SpV/7uN0518TAwW/lMtLayiZBXnnDM9An+mYYbkT/030PL+c7V4heUiFWq2u
mMTeU5jUGNqq3SU0GmIWtwaYEb0EZVE2q1wT9NFck3uBJ4rpYQVVbvUeSF3/RFTv
O83CWBEMInj7Ukkz/iVmfqpF/jMw6bTSV0lEh+UNnU/jLk7X51ebc1zPbAYQZ0mv
bc7d5Eef6Lx6a3IpXlyvazp3SAy5qnvpzUjzdIjU86/4MPezfsQmNK9MqNPAq6vR
o1BkRqjxH7lIwkhzeZAc89D5X6TpSi7WD/q9UNiRZdOO9NgjQRytNnNuv9lB83JC
Xz8cNJ/VVpA1WRfj5mDQ70WdgEUGrTVAat0m1DBAg/WaADobf1VVutSBSU7AZt6f
y4sna7rBjtNGGUNg1usNhA3BuYEqpAR3tMsedF9vvPz6bAg6Cbk5xNwUGBNTda/8
LR2BzVrPtR5r0eNV0zcFfpVqKXwpvvtpPvxSy86+8AoipczXI6jwMyi355lXEqYS
SGX4LiMYGn4ZBMN388fVYTiScI36rJj8yracjtOc7dMIunJdqoaI6pOZaBXjter/
mqTBiSDm+ysl54BDZyQYrSQpCQhLxTwsneA9TIjw57KUsPr3Dd/gCck+SvW0QgL0
kDA0PR9bvNZ/wucLTKkTZ5JIrz/h885ePbfDN/r3cOFF3xQ0P3mf6ZV6r3DYDgCN
WutwVFELrat2GjFvzc2ZPXhND53RSKQK9z0uyuQjp54MlVb6o1m2/+HK7zDE324c
QFCOwES4gJUY2cpc1KLv4F50092nQL34SBK3Jxks3CubzSWUqMQFGD4EY+zhUvDM
YO1Th3Mtk4KPyneGXyFsamMMBvOGzMzoDs7w/FnoA4wZgBmh3qoRVllzqo2sMBGH
3rIlT3SugNV06S6X6ZLKtX8eRs4YxXj9ugjvfk1993OeNjoqzWwzMkjhLkTz6386
0vhlOCvnm7q22Ydu2Tjl+fpCZ5eJwbjm2xiCp0dLCV4Pqfii0CMPn24e6UFcn472
CaQD9ZuEGH76pyzl2chxtP92S3UqUZReo3oaI6++PL/06g4NPO7L3Wte3Y/TsPGU
Mlp7vGCmSH3Wo7C5hgOxIt0nU8Buo5kETg/E2FpUmR9VbHAIocjqls97p9rXOHV2
TOeOQBeOPf5tcXB/ek+6sCx6zqZ6snqIh9Tvw62cRi6foq2lhG7hs32zWkeUjg0u
1jI6g+uXjbTYdp9IqKOYfTdU5mWl19YZyQ9MWl7XF+J2BxGYQGt/DbCp+/UKJvqP
b63H0jCjdnJqj/yM9vutytGeDvUuv/WxJS8zX2cVBUfZfKL68H4grLWozSBZpINE
0VjY9ZDPjprpg7txEr4R9B70vwj0Ue9t4QNKcvYHYgApY+Eb0ZobYBkRu068V1ww
l9c1D2J3ZSZVMjxWccCVHnmXEy1NDYHOzbD4xh/A2rzQ+f8NiUi1DoiYbSIJaTFu
6+gU4TfEuXakv1KPE6pCg/MotjapUb/IhlVn3ARe8wJ5WLTyOiU6NmA9aWGfzq9/
t3pSLlFBueCa1T2GFciPpfTsdfiPVn9V4nefjqFfH14Po16Ny62DA7yskvpl9EL0
5NI2gfljUYRAtjSVChn9poWIjmqXbceZQZbmMFnOjdWyYEldTOgTpgA3MbwHh4lL
dkgPRPMa4hTmXyfJeIIb7x3fPEt78YgbCAgsBaVcjikrv0lqm4UK0ZJU0itkysSR
9/YhuXnq31hUO2Oi3Q2nQAM4iofcPyusp8NqPUY5XOT6Fn93BScs/yAEKXQhgsnI
R/GlgqdvtvQ4L7DSr7Z3T2vRT1EZLyeE5ErTwRPuV7LPuJDxDaGzoJEVGqNh04zC
XHJ+k+m6WcMl7Q0+rTrQid5QQjF0wbyP0A923pX9BaQp1CwGBNiL2n7D0OFJk2c9
E+IMEGOesZ7/iff2ZR+GmNuThOMzRapwab2wax3iFXFpcpAK4un1lLd3gBAivHcV
l3UsS+ybSoa7Yns0NP8uA5A6VKpcbKPr40cp8UnLCh7zyDVqpjbO31X8drCHgVPL
PsbRGWfZC0ztGqdRehcSO0PkNnhXKxVRc9IuvotRnjM6ZC4HBxvvEcwduqtjQrQQ
+8VnGO61VdL+kJvCi+fAX+YPxOQir38RO2kWryKaBLqaMnsbakbLjKfKce2AcNFU
gbUIJRq1+q/0nnWXgLoktZ1j6EnAfzlPb7PGR0Pk28jGZlN8OBkzNnH48E91TOgV
x/VpR0pADVC9eEZrRiitwQ9bhjphNMioiS4g//Chz5eL/4wg4r5ZlCzkMzMiZPI2
Z+VlppW+4iRuHAAzvuMX+Qo6iv04oZHj/rZl17unc9ZeGPRvbSizfc16X/Uj4CR9
Xr9GqI/Yrifieuluy8aPTVzv9zLHF6m0fHZxkQtNReOJAaS1h0iXAmEAHPPFMYgM
7XB7zGJBMzVpIIbCyW6vpca9IQPcsKlWvZFTGZd9ZjsQnrEhwsITdGzUZRIq1m/I
4/XG2S8MjliiiDiOVKomHAXT3JLFjZavs+fL64jNuuk85UNzU1UGuYEPk3tLa0lD
PBQUB7wwmPvID+laDqooQ5ew3Q6iA3colA0OWuA4CYW180qW85nM150llO9LAhnM
yuQ51MyLBh3ag0gBwDiG/qOluF0rZ7f7xmclefkHJ5pe32ZSyl44yuanWSDpVLjx
uqW25I42t+/z3ybW4dnViP0cQSc5n6ZqSeb64SBcJJxgj2luFvmjL/ylxLo3IcP+
KXSvVeukQJU+mOnHKAffnxw0KOSh8sKivfCxhx3/98y9XDswV6aO9N0VdII06aJ1
EUkMKiC70e9BCb6ZDEp8VgEQ8D21q97z7YvK8T0MOrwzeQkz0eCzOKD2rwt9+wjv
vm2wROhw0FwsTDWi5rwWO6eTvPNOzn6pUewTjKRCqbmknGcWWCZFaeDwNsgH4a+K
U+8pyXU68An1HbcCrI/BICRDlyVu2gCGwyQiLN5XvrTg4IhUHRnn8fhP9YyJYLPt
R9vTiMs+ApArOyKcfms/cs+px2Sq4JF+Dt5wXtPi8ICOMPZUoj4LpeZa4SSZCYLe
Ut6ilz9f9UwmX4VuT9mJ7Qpyy4fshEXg/gVoVTX1S8W1ZquulL4/g1JOiqf10PW9
MpVoszDYzLdzySdME5fcWSnDvXUaap2GGC4tUpSEj9Ja8cslkPM/pcBKJNa0+oYm
D2fTrcKX3q8QcC2YzZh5ljBgzB8Q7XRGu5K0Ae5LT3Sb/zGBoEJVAxFLa0tzp2Io
WXLvOw///h6aCPOIboEie2AU5nSx+7Vn7P5fPjtXyU/wTFCKBS9PzhKvyuoMoxHx
mnSUIAeATt6N6zHdGN4YTWu+YGWixtdU09Li/sfMkarjSjiATxNfiKV3ZFaQvcDz
Tys8eizT22Qa0GxlWulebreogJyiNK/fgiGy/uUa0XFPOFGq8qpXq+GUn6V8xdCH
SLs3fYsiK7Vt2k3V9AgjgbdjaaU7dGjMdECg8TCLKdZVEBqCwKttX1K/IHFy6wSl
BGkUuVbhhOYG5DWhnqmo5HRZsYFtYXTAhPavWI9UySph1w96iOTyyzqhW/li3qCA
Xu8lz6ZP03RMGxlRhpgUNBZcjslLuel22b9y7RvgI2gWyljsS6T0N01novG9r3HV
2uP85wI5N10KLWsStol2XltqEIqji2JYBmBypQvPWc5M35uf4s89OKiszFv1QlJA
5qzmIuWoYyT/JSj9q5e4IhQsDzGTJmBW7D88C1anKfV4f71m428oVEiAf3DoSFcB
6UB0W3RYXjqx+jNGF1t4/vDB0gMQADZxQSPuZ62NnYdgd3BXg1XLhKHmLp48ogSV
0BKGdve8yxf82CeN7Du5NjS9U4wnxwrvn5vbrp8c1RBU3/7Ylj+VSSvLM+0uqKGF
Q+AiZyFd1xtJf0NkRLxlJdIGEQxNvHncR2PwZadG7Ar7w8reNY2GfIDNH1Yqpm0r
E9MLc4CogqbMLyGurZbA//OmmcRfpaJWGM9EVGFZHFG1zwA3xkpjxB6Tp59Rr22q
qqTuHKBsdFDJVP7WfBAqFFKTkw0b6nXAGOIJwKmkdhpes5U5GeB1LrWv5mjJ7ydv
Cyo+bVks8dY8/Un4FjV5PUcZ6s/tOPbzeXcZqsBNAPsAmFKD5N9ZC2R7vHoFbBy8
cdBkP4OMVaNw7s16l27MBWie6Xe1EUQ8o+uXSMYtLmH+k1whRgT0D1S/5hfO4PS8
U0RXv5UDXa79onx211U7VmDwA7rV/Ph8R67+qHXWiJB7N/yavwuUBslytJjDPFvN
ReDges37ziu2wVbcFk1qcdHIMWKfuijh3OA/kZrih1PUuSIFynMvoysqyrX0HzZj
OoDYH47Lq2gVlRfupgSMVhckt7bR9cdF1uyX28aiDH8pFT12PzckjChgUzqVMhpL
wQs9cCCHz2MDY/vMwxfSWKgkkU3znUMkesp51aAqqkkmxQg/frmq/dmJYjNrdbir
dnAoZdsZaKrJW+TtN1IxSWjUZ5mWKrNP5Wa6FMtuSDHq0m5Z/53AogM/QYJPN8CJ
E/iNZ/W0suz0sxFYKl66U8kxS0Uhe+JoeIBxmR/G3yvxAtTYxw1Tv9cZhDAI4V05
NMXpmwKo8R0yEdux7Gnvjv8nAGtLalZTBFKdCRzI0ICbOBD986VAgr1ga7msu5+n
N5efjB7SLWQnBCrzwcpZRb5b/BFSj//Iadz3geScd7E1vMUY8TQi5SS5v7627FBP
Zbv0A+y8k5ntoiaJeXRJMJbqPAhl85esbT+Z1ru1V5H5+Or9N7lqHXsNyNbOTFBg
c6mEmDaN6uiYuOqtluY0vCxvO6xRx5jKIYh3S4KU0On9GsYswm1Eyztf5Yp/dB8A
YCyy1W/Gv+3YI2v0ZIKVQXovYPqKEDixn3YYuCMKB4X53YnPhA857FgY897OWJ/z
k1gxK6clfb+GNDfc5RGuLnjBDJ0+JF008xRfgZLAGYTPsPSF7nk0qhoMQpU12XHb
7TfVfazihku+2184jR3Rt6Fi1gn1HUSAjLcEYp/sGXCzpJCLr1YCGbv70k+CuZ4+
Vc6vUpbFcvZ6klC8+yW79uhL7TBwiS9z95q6D4Vzu+DcnVD6ohkpFTYF0BeX/ZHQ
HXfPvsnQDV8+VURHs893wfscM8VRwYgZPmKnBtKheL6AXB5+i9pYpE5jaO6m1oer
zUw2RddH31YNTo0OFlbfvvjsxKWrmEFPPp4Plwy3E8E6PsOkOyBWkEbUwyphkuk6
5tDy8UYG6lYBFEkdAfOkBORlkSf3RMFkpPHfi+ssc+FtgCg0x6H9DaYlNJSVYTAU
sYhQHbJpiVYf6s0q6Svy6V/2oNbdkvxfoK9tU9MUCU5nrevu4oU74dvUcOMSLjwy
3FGR0zwrANb1W4DYFiUOMd6E/hCIzXnAHDpdYbO+zmUdjQMvgR9juE2kqqBNiNN3
gNaXM6c8tvz9HyfrKAPa3/R668P3qmKlWTzYMe8FaLgfj3cE/bt8RuXc4CXXbqPT
KoOAmbtGqJ7G11eFxE+RpngZQsSg4zzi+eFutga8VnBz97jktyDAR1gk5X5DRZL0
QciObbzmTBrunQVVhtlXlKodDeUv2+hnLNt8nl2JznsdgXUMakNQrv/3aW6RaZuC
y8KUDEspx+6MDGVCTx4gCjCAE7+A9WW/nYjhjI4URELU/X032tSmoKuIIHn9V9gQ
hui8Aa/f50kovEvJmuhDkGEEZrsHQfB6n0aVNI00qFNHxB9m/yholYBTHUoVMt2m
24OhArJT7VpP+PAFOgb/yJNNd19NypEm6Uk3MLVlQ2APfTnrMDZtI5cXcWWhYjv7
AL5i3ZP6Idn0UfG2xGO1ZcM7FnYyUVkn8ub4Rz9HX9w9/jcHK7rjHsQO7HJw+02B
opMTpWwa3zvtnGLBJUobrEOSyIoxIDuNDbgi7D0nb5oK9OcEYylvT8MGBAwEIS9L
slhXkLtpUl+yTVjsDbC0VU2lpzzOsX3U8gfk7eIf3jIMNgG3US0Dzj+DOzCydX28
RK3H1lWH0e7l4ew9bAdWOsf5IWsuNPgUNuCEl7bGWjRNN6rleKBw7S2AIqaup2FB
EVgdd69Bn83JuCuPMQ5sNojYyUaXxwrfHalzoRLGqz0Ow9bJCWBrBkaVLBlO8vlc
kKWUm1U41hJ4DgML2Lcb4X0bw2s3gdVRgUcRrY8+V3aZQWew+617JjP9SsNuojCW
cWhQakQCNysf+TMSl1003IGAdye0hxgUIcC9n/8RolHQIDw+Jv1bvobcQY2qOUWP
73iOjYG9mv0Qj7BDrwN4fhwSaUnn1v6aLIg4lMTSxdu0V/3ahCHiJZeD5rHnBFcN
AMVmiYGG/TZUIR+T4t0IB8Aa5un5UzJ89kR66QYmP1YgUH0xOd97RtPQIPRf1DTO
iqMxizbxfFtzNqxgI6/aUz1yb4myxPhqGl8Wsii7B/ue+i2nh+xhulSrQXL4ELG0
+0orOhGcoTmR0q/WlB8/KZ1NBSSDGpTSth7uVQsfas4S28fQV6lmfGh5+0wBfPXq
y6APii8ho6yqFr4w4z2oRT4UPLgSnQwGENsYD42hNVaH/Kpkun/v1APXEWcV0GiZ
h0hMt5FViy7Upwr4XJK6yt9DQhp+xeE7EMt5gMcn8whNwkIYcNdGl+igzMfH7NT/
1n7afQ//8r9VdYuNYSHRzJyojRfxkD8qFrfFk42urLUUzrX8Bu0WMj0SGySAjFZg
kMBh+BFURBr/G/SoFj6BmS6GoCuyfhrxGpzFGPQcOSmV5I6i/GkpmglDfHuRBzc3
6WooN8mIedPV0O0LPOKUx9BPq9mmXKLnuUK9INmTlOjVhdILnSbFFamnJ9xSJSEY
aggWoECOf4/zYnJHAAt70SO4i/5bNUF3f4JwqSGdoUyxcJflTULok6rqon2+FDNJ
QJLGCKL+c0vr7IutAtVAfyx7ol3GD16fPee3kqMlRUTEyDKG9UlAp+anXWImVPbX
ZLtKiMnOW6lI5ldhLeo4aPsFfM1I5fOA9e2tkGzJYvPAisdiHE+bF7mQQO78TqvD
MRfqVj9OkN9JOSBnv3jhxvZ7GW7lvnieEl9s8NJMnDkGRm5is8dFqWrPUoG1Drkc
ojQ/ol6uRqHcZHLobIVCLbq52ttU83Tv/rllqX9rUNBrvHRgnzAz9/FJY7WOXiy9
CxkmlZ2grC1m6NE8KEzRF2gtGUMiwh0fpyp3Glo2+pIR8lNhDd6Tay2XVfxL6l8S
okmUnPczRCv4TRKqNURxYS7xbejOddrHrZVm7k6NGBaciUOSSfi6s3KyVuj/lyhy
IBcEf+ZJmZu75I0IanaCuJfmqBBwW8p3U4VmlcYrdQHjD4PlHd7o83rjeFy8Qn7p
KZoIAq+FTPug6bi7qawEarvTvPej7cCqmOLwIDueJ75APEBg87PkkLdUiBQbHRly
yhNeBUr7tEWxaDgSr9G+JYEZCJTiUivEQThiR745PfFCSYJJSvGIO3j5/t0BexWc
idDBq11FVG4qG25pa5Pl9acNKxFvdVN4XWmVgC8Tc2F3oJlQQvMbcp9CX/BsrwwJ
Hl8MvIc3LyVfbvCORfT4K9gUBAx9T+zJknuL5rKuLtHYDorkBYfK+EltvWWheRdN
VvVvCmsJu9xgNU8s4Qi7U8LV3VZBMK84KWmSYcC7cgRv8/+xk0uMiWRNWBjUHwMu
L/GJXop75j0PkhUS2tJpE50aeejkyO2tRhPZTN7lF9zFCTtWeT+U9onHuI/4Ejmf
kwY0nHHz2/3aIPOwVWhVOSZjS42LnOt31P4EH/T6uY1W0JhcN0AdPbLuGzYBoqOx
XsQJD+tW7e5eeQrzZQ4tRkpwOcpJcXz0YgaxigVXVq+7d0bWWxUqpq8nXyb+DWqi
YOD/hgLDAu9RLp2124hhf2QDJGZ5bS24fzfXsrdiBoyzPUC2+t6+rWrjyBYHZkz7
RpVi6s4b/Bx9y38Y8v7wA0KWIq/DISE74YuQMKG2wpxf7OFkOAKJ0waSBUCRXPln
hEQAoc9ZuPSrjE4p5L/yT1L95mEtRNX61x2PC0Yuf/h59dVtOw2o59hB9HZBATtl
hoi+gkc+1dozBGvrw+MrkgTyDk5hqbkJRDz0mh7xg5TWBHaNnCdpe2/2hPf8/nRi
OjOOo0o2LwjSR0LQ6GtW0lmmTzaV576CpNFX7IgNi8RDYCMYELcYd5B4ghSjR/sF
hkBm/HWdJyhSU6F6T6c4hoObMlKuOCSVI6kmdjEeNMrGLoKOSpMFBaarEZqZa/8E
MPsbfQRA0/wsKSlefse6ha7W5cdAitkVfn/jszIGicg7KNlJ12JqA1mP3HP/ey8r
AWfuvhgq0+A64UlqEmoXaCGx2vOQIIN8Im6B5lglU1wtYULP8Rl/xKDOleB3Tn6v
oHoDud8DRsw4acQaJC/quC53xQKak78vZ6aXevuWK6er1wsC8lQDNMdSfkOlDbBA
08xe/EigIsaHv8Ji5zRdQNKm3JULRA6B/1u5/wpe6WaLPFWyue79hx2E72oajWa9
h6VC1JLNjdK8xwWvXRhLLBwEapUqr6NVCA6OtBuUgKOzlGAwmrg+HPJKbIWtobC5
9RSTh1fHZakc4Hkuv4MakkjV36+RbBRClK2e3S5oCEeYkHOr7In8M5bGUjNxK3Si
ghKQN/ngbPOJ2bJTwm0aLfW1dwKaOQ6IfmZIoUoyC5dmf6DNIlXDgkTRckdgSiVt
rpNRC4ErQiItPTn2yYeJKIKFAChGmEX5ODUluRE1SlpiGnicRtJFJRHNV64/kgag
J/iRc1aFPdkOxorLzhc4Owh043YYIMjYVtfNUqi2BMlEzUO+NuzuEbikCCA/b1ru
oMN5FR/NM7KlMSmC0bkJ89pgxapM7HRcYjeoRLqQn8bDK95R0RBC1HY0QnBsrFUF
v28anHer6mBykcb/bjbn3evpy0hdh6xPNvXCopXHsuhYIAP/nHZLyGqw7UrO3J9W
Jadb3wnJfer0TCfA1E74cjz5Uco8cRy0ZAtD1/+QRjcSMukYyGDw9kYGbHqVWaG3
JgrMiU4pgZKkh1deuDJtEKaulzoyelGaFLYDyClgJiyJrYEBOcm0n1/EbtBcI7/v
ZMyS0RDIfZNgjAkhlOAhPQvfJa930hDFCQJWPTx1Z6jWgRGEr/0wu4BoLE0kj/WC
GcixHUbYjP75vTW/xMLPMrceb/jUE1DXO3C3ZZ+nyYCsiFMpo4baBXXwOSRspO8W
ZlkDeAZt9lr+mYfrScw5lVaTlrkOT/3dqCHdsz8QXvwohmofJWuxv/l0LkaE+cBa
ThIrQr/qqZfXKnU9ABCA6jygX2/2LFsR7i/GEMitjs7R/umY1hgtoGh54ipBiAXn
nDYjEQRPYY3O+o7mLnl17AAMNYhSfbb+WWtAnx4xOJqYdDwTBR670GgGWclZAwix
9JftxiYMlyBoNo7Sr1mWg8n1O1GQkC2wxLJGPOSfGkAAHTwNVj/EINFnoykmEW3J
SgtFP0ldtUkgFEMHfaeUTJpj8MiSRTfyYGzOm+kdiEZi+sIscrwTM9/gQF2xrl9+
sMpBSMs8wQeeWU034A5AttgGLAYekhRBu4PzaFBvQ+LVQ++3r1qELMUs85igZD0n
EYNwusOr2OOZvQouDmwA8BCFZ7c004I+qab5MJ1kmCdWTGGznH2+xUQ1qs0V1QnH
9sZE0wqENL/yarPZjttQ87CtkY/qYNpXw2EINYKJLmUn6JTESNK0vjBvGqY1euwt
HACE/qAcHnkYs1nrZcwV+4rPrHCuOLlJTHiGAfhayyzVCq8pMhfe5mhvEFzjrSma
uVxKHUF7pfzScy6QocXfLQJIqHdjS8I2zqI4VoyTxWLzcw8BK/958KYqE15pfvDe
Le9oZ5TEg/jzq+ar3zGExypmgNrgr5JMRrZgTJZ+3dqvnKq+lS+n22vhj1d5msDi
QieC9m82DTqfKmjn4uEZPRU+0GXzQ5LNC9yHhx4HkxHdO57y0I4GWfWgYU678ZzH
ucSeTnn0OJvUuRcpR7lzWXOlHM1kVNwVQLavW+Xa4Kap4IucQnu9G3YAupMjCG+L
RIQVKAOWqTaMq0Vj5/gJbRXJMHpUo+SekYgC49tJ2tKRGobQ6kKhI41ZkO58dwIu
fzoOMYoscE1F2/jc4GLfZLWY2dawyVVk7x7uTz+7b/G94L+ouW9/7d1k6QRjQQi9
85+pcTyX/wICiowOqTWRNNMqzuC6h4kWdTGxP1KsINnZ30Rz/PWXJunBQc0u90FC
1FuLVD33wnf85zvhUKR7+nb4czAw9p5xaJZ3L8H91owgUJrIh43GB8MVKFF0SYqL
cGPH2fwjTxCOCd+Ttm94SmwL/Nck3QLrXoC8kD5ILH2Ly7UN/9L7K9QE3BsRkwNS
bZNN6cVJnwYhqeIOytCnLMSOf9CidzcBGGBQcJjFfCRYeoYKdgvoZqzywcltVT31
A9GCbdSjZi+srwYlpOTUDvqoJUs9WfeK8o7941ztnJw6pPOx4/tly+3s45L9qISD
d0/0VGElMS8TTRje3n4rbgbhVZ7SaDgHJatCpzDAu3sSOmMvxcY8uZXTiOMd3Ege
MnieB5kU8cU8CIDEgKRMx+xeSp05YYOKvJJBhiityvJk+5ScRf5peb7RpQUNUfrX
L+KkXyovw1ZKFnR+S8gznL146+B+w+wG3ITVzD0d6bu9BgtaKR5gNmn0N2/uaPG5
dj3gIg/MNqcjovyXg7ucL507oz256+gDX/Oo4Iy2TVXwkbHtdHEdh+cmaaDxSwE3
u9oQSMTLfAkV15QYB4Sjyh6I7cqDA3Dv7PrEb/3vSeu3fLsLvUx+TkRmhdR4HoSR
tBNgRXMDTfIY+SgdvhRdEYv/rQWzYF1BgcIp3vRSLuqJ9GzVBgTyl4p9hDQOgLmx
tp5lzVy6/r3GhHsUGG4s3xCo6Eeae1DX3Mn+CKx5ISdAc4dV64SPuMDK0cD9vLDg
2wa0IMDN41hHF7sgNRrIrJcKri237a6yeExsvPBf0mnMzAhmuY0XMUl/RMr1sj7Q
zjppgc5WaKwUrEGEEzvPEH4TZ3AJxbDHWNrWNq5sj2jYC65G7ZaB3RdezGfgpuDL
fZbtn/0g7Ct/ZeYhV3lXmYPyhZ3bmE5iVzTUYuoAezZfx1c9d8201Gv3P62EYTCd
Cx1QrSwSrdQAepZNURmeoJPHnzfBGPAtSIM1T6oqm4mN4NTuBSuF8OZuSStVU+Ln
GbzOuW35l1vREOd7yRHkK2SFPknKBmAesYBrYAoT9q49fPD3c7WeUNgRoTzTX00d
mOJiHDA4JQepdoustzdRPRx6QO+FXzRhOfZQXkM5myF2QGZVzzXOZGaw4SAEbaJn
k9aP2vGOMX4ABILnmz6z0XUQDTRKmIKrrZxSmzn/wtJ+gZPA0DoVQ5PwdtuvJJfU
IWAQsMvfCxon7tGFVH2DW1X8Uvyro/mYMaDT2AHtCch/UKd6YW92JXCamGuLhcuQ
ECes684UMDcovuyzolY1W1PwrOxY85Em2A5btHobqtuGpFJCj+nIvgiALBsh58aC
YyRmX7zJ3KsFny1NFjpkA8bInzlg5gJYutEnYQ24eYeewDdjR3eltTHzSKmABZZX
7H621AB1wFadTeSIGP3doGBGaPEDE4cF0tHYCi/72IvxITEzj/mnCHVlsSldfq70
YEXEG7DwNC1VYf/BNT/YMG/WJpciswxHLg1FDH/BSZkS1espAljPd1iPhPkRgGib
bSZS3qLOtG7O+HJxYQoCbtXEBsKypYZl8udLQkpnD5NHsml4bdo/bhlF/tpr1S2X
Rp8JByWHsLZfTFsNclr5svAAm/dT1hXrTOBamq4FepaiDdo/RssX734n/wvVNi1D
KzYAdvPHpHnHCcrIblHpr/5OBsGWK1hRz6VVI4THVuCzp4S5SjZPPhlALnJozDHp
tTx6L9v4kVXmr9/g08CAT9jU6wIY9CV8po7YyKpGsB+knxe7hmNW/t/h7yK8iphR
deMH3WngHMEFUHUgoFRAkxlS25T2Jmii59P3GIWQVOZZoocLdaxI9P1+u/p9qNRg
/Y1Ofq8k+aI+9eXA7RbhhX/2Oheze9nzjdkg8e+mdLUahX7pH0+O4R63qtt3H1MD
IXwfij43Rq8B6xIw+lLdG8G4bLvCPyhj6n9vD6Kk+jHn0DOefv0gjw5pycJS5euS
f/bLX50OvzKBfCLbGTi9ThYbQAX/PFYlHsTXa7EJjT73VjiXiZjgXf5dt94IWl6r
qf9Uvku+9CHo0lSIe1JwwwlSo+w+rS4Hmq1Waz2a5KGphK7PnCzASf/lUQJeVInU
4Ygg8ldxVgcUMDc/1tlY4PzFe8A60bCywVm5gI2NW7yV2qZTttew0gXfOnPrO+Gm
tSgb/A1vXE+RZRe9Wwv26H44JUs5Lq6835s71qMfCOvFujadlT6CvCUSHP2qPYOn
QWYaQd3/jz/YWnv7mHx0IxTIyRQb+rTTWO2SpMPiuv9TjqYNNHMckXYjnPxQe1zx
KuK2LiHFgUxgmFz+NBMfZQlruRQFh6xZ16zNKMykFF+VvI4oycIZPKVuEZpiDbjg
15l6zCrLTFaHmRolTNy9NhDF/6uT/ivgMcfb6oNPynivDNufomYqOQGpV7wkiaol
d1M3UmvxLeyyQlt6RwoAErNA4ErwVZqHbh20TtyGoWu7rEoAMWe/0j/6VSZWvyEe
rA/qEczP2H4GzSfVliRhwiP4kyVmKwdiwi2LkZXOGyMFTl6Jq3GSBI9pCDZxRbXt
tK++l0RuStqAiN23y9TRxAWIRbi/husjCWHrXMz/q+D/iPK257TBXKsrEap8+mav
49j3nuL3eiTVROUS/iNEIO0NpOAk1BpbO6g59dvuNxPJQ6+bb8sJLAvBrwaCAb73
8jJpWz+jCoXAP4MyDvvROzboJkV0LyjCycLFPOFssSp11cetXD0id/+ewUdcXvWn
i6UxtSVlq+EDBTErrY58LzeRS8RHNS+69QFaRlWWnrfMBWS5qYOnlKUOs6n6cPno
IQ4bRhSEcEIgNlHr/wmokxGXD5vBJG355/ge2Wi4UxkMUONVRl/lARe09KQ4DR7u
BQCeXrJJF1B6i1nbpvp8nZsqX8xL4C1IkuxpyEArues+UFOvLDEfmnS4M8HzgXeF
PTHEh2A94uoLrg21UAGBeeeSpB7oLu8O9NrmYMMqWf/Y++l2yi1ANk+ebAY1RaW+
xbCUTFrNcaNpoEpUv4wYF0XJCbAXhcDOIx2s67kKrmoDD4xieYKTCy0jxatcRdEk
to+FTPc3WYhzr8kV0tFQu3LGMA+TlHmF9HW8JdCWXtoKdD7h4xjd+desn/ToLvVY
EUbxQp+LqwHczeaWSs83MyYvOlPo2jQwdU9Ikesm6WoMyWDbdTVC31T1fvNE8div
EL5Ue1WzeH5EBzlyIY7ds6wyIYXz8a18/rJMdQu8B8TNdw3JXBnG3HsK+UkrWTHL
szBoHeFatIPi0Sx+OJRvSBgISYhx/XYPtC0NFHMXYBDm8jpZfScnB75yBfRxcrMu
rCPyGYdsgRedeQC/Z/5RIkzuOqcG8bOdSiK2AwyQg+plYhB4RokuAniAy1vU/ATf
N6L80SEhWl4eaHpweY6TZ3cWuYvkMAkGH3icx07jZY1llsEu/7i/g0FxOoPHtWXq
HxOWU3x+Z7V0GM/A6IAX0MxhB0RvqH4grbyebgLJAX1Qk2Gk13bdodqV0tFj+lIn
rYHCicD5Ychj9W4Lp+oocoKY6XiXp1Fi4mcVQ9BNRgCRiirsEQRjmo3xLstorjGJ
PRwCawVvN2CCW1JB3vGUxuFOLnO65ZfQH+MJYdF+3ObWm3MkcYGYLPXinn7gXdAh
4MdJkU+dSoG2Q8yEJeTgnkrLemZh2adYaJUqaCZz4zw76nB3sNv+TlS6nVl/1jcS
YO5Ma/md/AR22SDz5Gjz8XkwSjE61IxhvWGu1MIZK72oJ1uvJo9q0c0DR6fB6d6m
n6RoguIENOqDMG3uM96bNuyPfkm+qiayDJDQkND+orPV79C8vH9atG01ChAJywQa
1zDYn5o+wn1NaGEXohtVywMU6CJxnvn3JsxEOOZoy2i6Iqdva5Q2k9TkWpDq/EJQ
N+apFbkOBFSwXh5dr3BV7K/FDQWpoVwnBf21Qr/i7gzp5+pB66GmaODdrlvyf77k
IR71Eg8INKzaKIjduSC3ZBLjrjnNepGAzXYSLgvJ6roeHjVXU+CeuSUVvX6Qirsx
Y+2ZXXIieYjEr2Mf/Z0g8MQZQ4JRFJU097hpNlY7gyUvt7PMpaM4R1n/SG+Du3bs
YtTc3V2Ww/2DxPKc5mjWEbq944lW9Cw04z/dZI9+B+f13A8+bACckB+ntSTlcPbv
fJ30FFbpGRkjM4FyExQIzkG9bkCL1d4uSyu5g1xlu7up7do1ujZFFVEJhqedpi1x
c5uT4eghRuCnJTGcr7x5MR6ZuqyVADYyq7tBzcwbicbcxKg5UMZDs6iHbxytqRTf
PrbfrphbvXZA2MQbM9RAKOOiceagFh7GXQyqqLUmP/KoAJB/8wk6dw5UsBniBKO+
DNPKE+pAWT4ztXjS2LofTH+652jY3N6F81MffZ57XHhfF956pSIS+JM+qJHQgFIg
Ca4TDuz0FGIJmMXeOYnQz45Z4U9HkKXv7Ku/fZrDf4pZNgcGeykV+zcUpKkcKTgA
mouvgd1Xhd00V2Bu2iuWroz+bgJEeNZJ8mWFSVjTdKwpsn/rRO51ILXjrKASzcgt
fi4Y06PpJzAM7ZZhRekxT3+rO/GI44AV4ApHdEbhbH1HFWKMascfvAlF7J4G37/A
EYrjs+sDXsDIiaTJ50miwOY431cn7c+pF3DYstTVm2RixbhHta8zH/VRz6EZmSvD
JVmYUROf7WHt9sRzCz++rgkT6xHyYv6WztwBn0l3e/rFY3c38qkLIwN9TSOhsJFP
4FxxcE1ToXK0bNr4F7C3BKs0ZzF0I/uaD46NF60GAWrWpYqCoF0ppmdWNSSDAnhO
bhEKMeg77fnJ4QTuiU/xv7CQrWFquiRQbBARP0pyIOybRK9huaFIpuNmn9C5Y3Us
CDTPpJof4AyZ1clfUth8OcEWN8EBX3HBzKDXiJY8doXWqJKrmGpcG2bbnN6f1XPm
7YplkHxq2XQv0v2Cap1FFu/iRCOTRAgA/PlIl5uTqRZrkpCpfKFEigySruV9+Mun
uLDhpcnW5mxUTcqoTtUSV9m5zOX4wrWr5tk3IlkGULWWz4HH9gfY0yyl8zHk/dAe
7WTMRSUCrL1MGbzj9Zz1uHs29z77GvhXPd4LgdOYPycBIKKLBowKc0NOJiICZ+Ep
yrbID241VC9OSDvFj9TQDG3G7qYSVF5GLBIXFL3SCCA7MkWO/cvaNQez8oOdBsw+
XDaVl1V881nOZ83jRzdhBu7y0PmYv7jjWnQclpKN5ZOPaQ0p+eytuXlyNBa3TE5J
i91FUMC4FbqSOCDw/nHduHx9bxQBJ65JzkrQv9E4ycWPCDDe+YdzBb9lePuZGLZk
AyKrbuTK5X1lx3vLntbirNwdExPnbkOBkEUje6yEbq+U2cUL7xFTsKnbqNOAxMuN
FMk/ByalEvJPIn7lfJ7w62TwnJXVgsRHaLAhaiN79thJXDNZYG1j+G047VFSyo+2
DrIYhGcxmNXoMDnboE0+rJyvL3hTJCwuJru1honhfVkjzqQDx5C7mMUMPLRowJpV
vF2G73V7PQ/osjRpTo8i1qfsX5JFnM7uYKRFn7NofbCHHfWgBgYbdyCUgmNLbWAv
2GlUnXLcTSI/Nt1UzdJ2zjrZfsLZOPdenQfrWJ9u5H4uq2hPWXC+6oR4Sjbtseud
5Afc6ZjhsVtfhiOhj6cPBpLcJVbQB4Wl8fO4EVUJZ0sdOw5hWN+cyFozFeSvbW3q
DnDZe1v+55wb0h7xCUVoKwFI0stDDibAlvfNQtv6Bd+/x9StNcGxOLvLijfk9TVc
0f5AsqkMOw5O3sQSvokiq39AfhQomV28WcxVXq2QMehg+Df5IHSNrNFY7cuV7gdf
Q7fmZj8yWb4igV6HgA/Qmg/WmgLJdjykiP4ig9QpDOow1RldCYWmYt1N3fQhYnnu
XUxtVRuzh2RtFwrKj+f2FFrdfF/qIgN+1/FJo4bdRlxH6OzCLylJ+Je9Mvhi72OX
JdLs0VISAT3e0Yj1lmrblpW6gPWTqdpWn6440XcCFUDZ6WIBEWHKQWcf1a/ucoE6
6Hc5tjou/PZvoCtSrYe/EQYkaJfqL7svAHuip8aSn490NxVAJXGx4Cgp7WgJSUDr
nr1K3OPp8kWH9cWq0zKv7OxmQs+BFNb8ntr3KCa+ii3y1AbHOFJNGu5NxaGTO/+S
5RW4cn8vGhfZ5BND7r1ae0ir/29Qx/IUklF7b5rW9rLhpleCOEj3o+RiF3so3K7o
bmUGjyFBamGI2jADvE7vp+LXyim4/OejblHqosmi2xlGSHu+pTiqMONjTj7u7Edr
HFQIfFNRAWH9SA5Jm+L/pesSqVpPs6aBrwRkw+VXH/333pD4I85r9qeJcYvUUHYh
qaDBlLN5bc8HMlmQupJ1LRy/2vRquC6ya30IehZUGJmBioA81ctcWeUFj1pdlNKx
59mhuyekNRFwjiUa89Xhsik20vBXssnd7yUEwnGXL0DhPGfmRCeQyN0MQ1BWg2dh
rKha68YjCpvjyVVU/BAvJlnGNKXjFelukFxFWbO8vY4wuAObkdFw9rUMTsyOH5BU
MAtKmYd8ZEefS0PyGRigjOqyABOlVA3yrfwvQFF4w4L+5IIBGjG/BdWooXS030WG
0Pqpayd/XtRwDRWZ+qgP/MeXkoSGFiFiiTib9LshijGjXdLOSgmuBcFMwDeJEcSV
fEIReMdt5O0Im/vGJs6ceRappdueCs22+UAnwUj7eadyhgbVEJGefJCgFpEn3Hkt
ZMhcvFcC5e6Yz5Q7Y5c3hN7O65157mMBkPhStgpQmYBJPH//vpViXdAH5JWe7DYs
EDrOxJe+FQV2L/pp3zzfl+NglPERHqV1I4UeloqLdK6YEqORDu5PX0dN4FkIocHE
J5TEufB4y67dAOvJyS2tHQcb+JaiZcYChZRM+3Tf0lEF01NV4M0UdncU8HdaRKVg
T3e/vn2gXnykFK2uHAGJCrsHKMR13YA2pAoRu/UMsVxMZfeO/tRlXlx1/8sFre26
DLtb14e1RLePCjkjrfwLrFB8g6B03xf63SFeCZCpvfnS3lwf7+71vUalvcw7z0m+
6t9ULMV1zxZe9APLEba7yPPaPFBurrQIM+dsmxIa/8IfV5l25g6zvHA3MvwV+foH
+jQNFH+w+y9ahy9OoMOuf2G/vM6YLaLA502fruweT8lb0NTkhdaetdP5FMkyFg+2
kT7XT7tLxWdbABceLRmvktOwlNurjHF/HP65b9FiyuPOwR3wEsrnweM9Jywrk5g6
IiX+PwkRxH1cHEkKajW3fwOC3m1AZ9LgQEPDU5tHlV355botb57fX/rp+S4HuOeX
za0gBvyrWXspvfJHdyxGzHjbZZXYqbCQvnJfyJr8RgGRuUh33TEVICj6GIB0Ritw
9CjGsACVxijBLPGmlPVpJH+PTb9+77oyPmFiUa9Xg0U58r17AloQSybtN8CfwgEM
U4pWD+vOjtmr+Pa2kjGJGNu4VS3N5MYvCdudXy2cBxiialejAzWetwroO5V4l5kL
8mxFPPLZF8mJ2Sxnf9NRiDYM58Pd9l4u/ep5DKg1QyPAwqGPMqzqipC09XJurU2+
6/d5dareqytUD6a6LwC5RGiLIpyva+HtiUl1/9yv5FkkGSKPXN9LVIU98pEsSyXW
h5YxPlQ+GmzVtEAkUg0PABOxOM7MOi9ErbTwzgTteLxQGU7vzmeCgVqWssKg8FH9
EEcS9IyJbs4jmq7uARwHx3nUBtY21qBN5kF186MvxzBrkbWagF/1LvE1c4Kx4J9v
csuKdlHuXKsCQrIjMakYYv3al6ln0cew+cX2jIdyMakizKULe9w5tnD9ttco3JcD
RmQxwY1MyJanZUr/029SMqLOwMiHg6FkhQdxRJEKAJXiELArCqZDtAOzkMUpjs0m
jpBESgNF0xA3M2Hn+ZesTiIIj5/4OCG0uL9RCFsvmPzzayJ6EK9laCQZc8X96zBA
+iB0CZ5qwF0f4U74jhs+mzMghkbK3XChebpim3V5q6BtcV8oxvjbK2TqGT7mxzT3
I7Y/hY2BNIO1QwMZxAevsi7ssvxqdmQ46xy8XgZi01oaf/QnNi6K2X6bs+7dAP4p
bYmDoytHI/p9qQyr1Sp2qGg2mg9Vw24aNmqokxFdzc6KDW68LG83P2EUP4Ycd3Fd
Ciy+eTHfdHSOrnNGKYzxUx0sbmL0cQibGKH7PpwBL59Ojskiz76/4TPkTPlZU39a
18tsaJLtYKCgug1YBZBtJFCdsiCUIdf+cxX7dHoFay+vluynkX1KVkMxlMLo+wqW
HQ0DKZ7ddbzZNyMFKUIqE2vYxiwi/1DLHykt7jW/UZOfyJgi5wRtHLH2+NhVlIIK
4WjOS03ThxQu378eLJhIDhhHcF9HKkodw1wxDtSMy/jjZ6VthkAbTF8FB+MgZlNH
2ie1GHVz2TdmRqNpWGgk7GjX506ytSuROSKxSXAeYOO7F+lIAjMDaiFI0/EQG1Fh
Q1/9O0H02Eqz08qZ51jXr1hlnp1hR+7VSOQizlHtuzbf63TjuJV/yewihAcVvsc9
wZaUVvpeGCW2z7yzBLwDhvbJcEFEknbYONLUnZH7FZR3+0UWJ5Iqyr2WS0zsn+eK
+qtGzPqxS98Uce6Ak9e9qGAglk7Fhe7DUlt8LkETw0SJSdnjT4BAbgJ1Py76uy3a
7503rIHR8FRvnRpIVo0TR8UOMUyydezGHLEZh/1pAXfblQZ4zun4tbETXBatrDh9
FsjOxhCg+xxPdhf+qw43d5f0MmHpW8LeVyAKuduCpZvkZsUG4TpVE0IqKOxVLC9V
rUWtt5WhMhlrCckAe6gEDGwdFX3ZLcQPBoW63ijXptyACDFC1UUOsuqPttCxEC+C
dG9DwKgajsVrCikunnnUhOcX2iW6126NiFrQqR9csr3Ecv4LHlArCGgqnq5itpHH
yjPC8qfShxoEmygelEJpEJMJPc0Vd4eIGAiTS3uhh3NJdPZHMN+lkSs7zUq9ElTs
Rf6PLcr3G+BBJLz4CMBtx8u0tgh635YfCrVChhhe4VWeDAWxgQ7GmdwPcpjwiJEI
E1DfaXu95mHF86QVL+CdKDmnMiR0rg18IOxDbHrke6a67dJji9IGLD8PCMjoiaVK
qHavQCez85IiHKZTceRRUENJ8uWxdlF65TTzEV6x0FuqfIq48lUfWvY1yQ973UyA
e3ItSEztG7fczFsYXJCk53BSvCUIeQROL/dc/PiwDm+jBz+fk3h0Wdu0pxN+QUpF
r1aU3VHDflouUMr+1blzeKlBT7lD5qERnJRUq1u2q1yarBy3pJvClwf6vozdHGKC
ND45lhaZNL3cQDIqQvx4+qu6wpDrcMuGF+h6Tl8tKKZFlcv7U2PFfl01BaxfY/cM
i78RvWqrJRI5AvZeY8mAJRFWExwqxYBLDShYB7h9usvBFm09Rh2AdQrtmiJCI7to
SZBv1OxTXsZELmXEgzkl/TXWk7yl2q8eS3Rt41A1TaO50TE59XjoFYqXJViPCiiZ
MnO2FN3MPixAq72IdaWUegieyZQQQt8dSf05u3ERYsFEHjLriyamJPllyWAhVIbQ
5lJR0XxFBtxgTmIoK/5G8+h5oZYxJNL9c8K5XiZHpnINneVBTDsZcwE5R0ddF0s0
YPx8YCbHDriHa2un9zC0Jz1M28F00ABUksNseN2p5guSCgehe26AYIU7vi9Z9zWd
yG+GUapKxDZiLfASRoztB0+KGM6ai908We/g4hogcLGcEXyn2sD1mLXYBBGaK4Er
ADaVSkWzTAe6HPeEPYTg1RqvF4MX2LO86xbfceppRjZoUjqPv4ziODYOaqRgK5+y
+Y2vB9UcDFnS4Jhi8Hc33B+7CtM7VO/dN5WFtJagFD+KiZ92IrWw4g2Q9Wd5DktJ
pdJ4gqvGVEkRHlgPtJ+gYZjlfvUG3kAla1NnivlQVE3AIHrTmm/Cs6gXVAuBZ/q+
L5mewDcq3j68eioL2eMrZx3CsKIv4fEQ6C9XU7LSmrVcrVGiCfTDFQgvBTm6UdM3
/pCcGwc6C5sW64gHBlGnVhPcRBGmOZSlJSoc47FYSPIvlZPht43tVm/aKkEqKXER
MRw3UGLYjacpAMnDUHd647IuBrFHu3S60Fj4lR3xChJ6H49IVknnbMK5DYnm6yP/
4KEEICSFUD4PU+XGBPwLwdx22ActTcD9TmJe1ogXdk7oGcmF1Gsr8Vf/TRDUiqU1
AwL5ACtokL3tj+zdsVW2OFppANwXztUkOthHrGfr62njOFWeK7JJa1yYjPYqwj1z
5LPkGlEHGu5ASmSxU5W5uwk+MqkaCwzd3oWYyIa6bvPFZVzdoKv5wsOl43fVaENy
u0fSBI4n/fEnwazZwYVEBgGf4xYK9wfaHzqvGpscqnza8XGEDJ5nNll+OD5AjnT3
YZtXLMiwZchm55bokIFVFSj6sv4vCDACwcHYylGXZK41Zus2BZ1ajR/QqsxSWqg5
4sDrZD4ne375jhhVMB1NPH5bz5Dq0qA0oRZi+s0asnvnOo233HuE2O3oOkZuxpSa
5IyB1OCFNgVmv5L6A7vuVUPGTCoxYe3OKs7uue7vPMKGBU/VsN1UaTu0lBlzc98Z
B7iXlSn4tqcp5ZFz/YtC1e9nBR9ynQ/IemRXhkq12iRm47dyLXQJuPtHuDVI/GJE
YEGo89lpkN0LbIa2Gg4/Z15aJG4kS2mu2D9aFYcj4F9Mi8ht/Th10446N0tYrIIs
dZHylB18Dwtsm0sDML3uGW0zgqX/c2mykfpEjmJ7B4k7b+g/CX5mcNeLKpJvV0C+
KkzfztTH1xHPyAUMy8BM+JS4UEonIK+re3x7wQ4EaxEZKYDTPYXhV/gBZ7WRyJAn
009/DA0GthZC27Ar8qImAj8SbAXoNe3PVGfUNW5u8gYlM9wGKY3cnriZX5MIo0Wq
i/SDAIk4dwibI0RPfvq9tA8O1ZV9NcktM3QjARcoXQGXh8QXvjOXWZ1Ea7hB01RB
Jib0UiLE7yds4An3U1CKhtVjbQOnAlf04fGQuBWNBklYr2TqbJjFmsfMKUfFZg86
vh/tcjPjnW5rwN7PPj4z7eAH2RTeJu24pNtQCC33WhWiB6eZ/hypOfiGlLhgDT9m
XAuxQ43lGaYwWkBTRMOof2BLEfQAN3DmAlCjAfbqDaymUra5OGvdiWlF0E4gfw0h
/GmHQACb1KcQXgtF6HS34smtcoK3oUzrRm7Eghq4YNf4ADDzY6Z5F+16Bfk3S1x8
4g6ug1UJ2CZ+X31vSb6+rKQPyuXYHNfXAtyNNYV0J3tBmNDwlDMF+4Zzsr8SLsi8
jKgWhIOLCcmVLI+TvvdWqV9rvPkIDWusdn2d2xs6ztjoGautiYuOPhQtv1zkxwyn
ief+2m+X8rNF7eRtPB0+3CCyFy7MBiqTocwdTon3AwgboN4vZfJ20f2kL4wvfWEp
MGMJ8hfDCtJv0mF/OZonqlaaWLxmcbELInHBJ3I6YPB5rJy8hJK/SHMAdRyzuq2N
2fj6FzBpud6nNdupKeF5v+eU29lvRctW2QnQSjZwu+2VsWGSQMJfXYk/H0UxdUMX
95oMXmsAEmHWX5OHmlI4AjBicFyOlPwjZGucPL7iXNBFGiSABbkW7fs+YXDBPzD3
kVa+dYUD9FSc1fyfjxY8A/J6dJpv+aolT9/JhOGs9UBDh3pwwv3MJ9Bcg3aKm51X
XymREpdJUGwTsJFRc5jS+zukDWvMxEHMBFbZACeeuaxUB9NnOWbLH0uqugzv2+s9
EcTBfHUxYsUrYZoNy3EEiMugRkkCAMXmDjgluxXyPpoEaxexElafvfyBM7ViQ35I
gaqBJvhNA/LU6TklXV9LOI2LTl/IZciarKD3RHpawFJ7H/peQZkpo7wDC1jrtnWd
/rUMiZlyxuBV27PhLFRWLgJ2ugT4PwspjLdRaf34TieQUWC9fyK9n4C05UWsqwec
HAKg8iGwP+k3zfrNPoBmUgp+QXkk2tu+2BEPsQrqaF12HGQC3selppd6jCLCo1gr
BSo7jqQQYXBFum0b7oU08/wkemrRGzTXsQsgeG8SasvbH56GPwEAm4mPyhuR6SDt
b0hFUjetSeTfLXwVB8urv4FibezXqEEpVlYSJZBPDiKNBY5QCe0CbwiEAQehCln9
YsoPnXtTLFnFDdaZty2AgS3GQknfbkOTUNoqffhISth9Iq1ciJ8NuT0GUXB7Lary
zGagBj26A6bG4HUhA+HlCLGWHy5x9zM2VlpEDoedqZvqCm0GJs7dMh/RfzR+Csbz
Q0IAdIQyFrOvRPzx9ERXtfWSTpJW6Owr20bqpHnn+tUwdY5zXgWj61VkXbVxVmZW
ugfmak6/hQsvt50yL4UEZi4sitSWbGVmDjXvv1omKt120hP3E+1b8U5SM+OhL1d1
Fda1+qKgRAXMXxRPMMsk9q08YcqBAYi5ghvPnJvkHerNvZPknduJ15di53zAmCPm
GLGYomk8OdXZ6htHPVuaL3fLVyHYUS4wtF4ODNyLdCrKI7pmNMWekdpCTQKgvcDB
O9hOWXT13yw7OYPrUu7rxkj957CYADmO17vxwVhM2OeMSUXAF+h+lC95e+PtdmAG
9+q3du24NKWlqRE3FUP4jFRM/Z5ZFcpF6RWmwMN3X1bJstfp5bpT0vUhu2uEffL5
ebEDaGZOloYliY+/Ih74Im7Oayy89os5dzeax35PZSwLgKvzNbbjuMQ0C3A9LcBO
YKfVmA3wQcdlJIUki2Rceb8dhy84DSwuqxQS/DWg3nV1pnEWv3bcVIzggUzxXhnG
SHM0nFoSqrjA9IgB1921HJVhjDBBrvbaKMP2TRgGpHTfC3O97o11AlyKL8UPYjD7
rzQqGkIpmR852swX9j1quilDujMSSZgWYe1BOhdAR28pKEpk5Hzt5XE421EYPc8A
vLRLnRONIbHw1eq0VokpYEahDPX2bSlM6XNuvi1i2pHSSkSgU4l/Cit0cMKB8edO
c0sB2K2xNZO9KMtn12r9cgXpOg5QERQcSAso3xoObbeYTUipKRcj9d9QXL7MRzDj
0kQwWnPeClLqfHlAHCjyzT0QcZII2mTFfWlkXu+TDJr/bMOU/7rZq1olZQ56McQg
x4IJeEILihnXhbgKRk1vRYYq/sbiJM6FMWeoErN5iVW4yYNqmF/GKsAr1CMueD56
yiQHyBQqXlYAWONVzHMzjb3yVmrT+hZFiuwjZTplwI8ve8AHpFu58D/9B0MsvFl1
hIVyvNXJEFgEVuDet83ITcDDbcJ/vyM87Lw9vhi4TmbBEW5c/lyYW9Dvoi3xcosh
TZgEYINZ1ABj1apG0JL6UqbCn7AAjDPIUO4oOk1HxqeO7lco1vlEaTLELfML9Mrw
rEDRJJES6ou2eKG/7S3n26W0IjBK934xMLRRhKiy9uKUf/G41FX6UJDmEqGE9bax
BGoQiu7s0aSNXJ2FMtF1Ru3uNzl5G5Ac6H4ykc+MSXsGJBorpzCKEPqY9c8K+mgG
RX7/cff68qh44pZjyPBPdjKldzRolxjdZ8lfEnXcFErBu23270cfd/aoXJwQaVjp
Ht6iCs1kN9Bw96+e3xocmiGH245+O5FBm3EvPZXyaoIwHP9MCw2yk04eXDEX4iCw
13xJq4C4M+GNnzlzDBjPp7EXjPSCvzzR0xZJcPxFGbhsPIkrS1XGQE1Mo9igtzl1
lEA6WYVb4FaJNMTs3QuSMNRF24cvxa6FbMvc+RccND3Z686ai6G8gIRrLTLCV/sp
MAqKJaYIz13eAsPxoPGUbyZTdE4nZ9ghTVs3ygdNh5L3nGuOzcjPk3RwuHHvO5Ps
ZmbYLvPrWPpheFz9OmnbbifSRVICvbiyu9vrJAtFJ/osToW/YMiXzbzIsBGq0w1o
opnuAA/QfMwfw1ptk+N8wjsp0az2wLeNm1Pf03YUrDUhlwuf/DRnpfvA9zu6CN7M
m27S4/RMbpWxI+8ZUjNTMOFz70OUPwYHtVHiCL3q7KqEzafO3KfUyUIiZaNqDGHJ
N8Fjn+HxuAq0Hovfcyg18NHPWWRY86p2PjmUKtZDOe36Q5vO8+w7pBU2gCdmLrM5
7NvhBhyrW560ccEHokFTLyVNtjhyJOX+Gjd76vajgbreo+Ho9So3zbL7Xte59nZT
eUbSZIqad7jSI1e33ZMSrqKyEQ0WN6G3SRAefNdlJSmwEyW4NM34yw9au/QMzWig
SsGcd/peSkA2v4Ds5yYdE12MxUYs585+FW2D00YLBZHftQ4S3yNpitH1I7mKmKqJ
50trSz1QzOC1PvfK574ovuuulpLaBO3m4LTrpz3gnOEPkeu8z0z7iixkNNFV4AKz
c4AuUQURWaf/AWk8C0lZ/jXDJVl2oUqwusDaC1kq+Xo9PlcCZiDnso5YJgMUFWL3
Tla7LHX9ztn2u1dWC2qPAovghiiuKAIUsMMHwN6DEvkNAzjSmVGoZ+H57qkG5Pwt
zZZOVhI624nOogLQ1FKruH8T9YgJPDpZ4w/ecQysyP/8GQtlb4TCRpRzZO2ZBKBc
mlNLlKg80bhMbn3A864pKV+evoL3LvbohJAx0npQ+E92fjC4R7jIti3hNmqQtuv+
lxhZUA1JMETe7iIJxj7m+/Fv0r8za1TxrpJdaQ7eCHcWvmRVKBcQpeIQW/FLia9S
m6TWugPDjXJ/TAROjduy/xyvjrM6QxF/ZIH097PsJpgQeoxnk3e62Tc6PJ5gDwrw
RvPtfwSS7kutCStsF9GjcbnwlcVc0jc2W1frFFefXmJQVt+w22yt6Uc32HfFcz8S
hs6fiChsT2ERsxFbq4UArfSnN9JKVLWm3mTH0uDyexIIHqHWeDvUG0k9t3Ml6VKm
uegIhjEdfALlhNCmm2Xqm4Gdm8un6qy4uf0eE6+9wFAlDWhCuFcMkBGm+uATnVAR
sYstlGH4Yreb93ROL/z+kHT4WjSXttmq5HKFHimFGxW8EZOK/1/sgF6cWpk8PmR5
GqwmVlT+8AU2ElhWKy4x9h661apSmu/ojoblYVGb4R7G5FNXeL8dKHaSKYFFVMTF
IizTkyGyFNMdc9mHAA6UYJA2iFuv55pGnorzGiKMn8tZ3ZXbR5C9d2K/CX/el2W4
UIQ0Vy0xFBevS025Ya1nVIo1Jlgy4opJgk3p16v/ph/uzFt10X5eg9sThaj5hT83
dQ3Mqc+6HOYB6R2WkqKekhgI3ItPFO1N/7DywR0OwOaSOzg9ayK2pdLr4hBI5Ryh
P+asj6g8zOtAfE/8vV0Sn/hw5cLDTISrpB8QCgI3pME1/8DAOVwfkJz/Asjb9Bmf
l13LedLm7B/017qY00O9WnI/578SkBh7G3E6XD+oy9rXlYGYjJspOXMb+iKWLPrs
aakCuMwA8HSHIFdQgq9nHClWHviTTC4ufwPGV7yI0S2fsYzJa4VqJBEG1SOmEqLu
cOsVylYsH9GOd7CbcdEhgzErMLHHoHsBV/dJ9JtyR0mVGGTam3WhSmQPtC/bfnuq
3QNpzcTiReuriZW5ybvp1UvlcZALBx8dPpXz3zuV9efaKYPIKghIAx0BtArgJECG
ID+1ZD1CI4MuglrR/Ya5xjf5LPZocgWxW1h7WGh3hm9OX3JkoiwbdlyLA0+Py5IA
/JJZ7If/58WM6m8j+9LwWufKTBhmXzvXvNQXwTfDKjbESxCbbokGI7dPEUF5da6O
GcrhK6grjbavIRHiOYrzjrpycNSCbkBnKrkUx2NN0t7DYce0Ighuu366HpRAIQ7l
mZqCODryjXcHPO8DJvOTUvQGYtg3BmowjfzxK9nSl7S4Mw4sWaBIZJub4sSvkSmA
RPmXKn5G1G0n3psPJeoB55edJcxJm159FRf1tj61BJAw0bk0t8V5/yjKVSQ/zfuk
zux2N6kPQRh1TL7Ip2uICL85qaeXQ3tomv+xedpfYgyNifnpQyHh2teDrIFwIURA
AQCK5pbjg9536VmkdVaCPkfqWTGUG5DBcgYNxEDgem8SoKBo7qgam0PP0ZRSu+aF
/P/KCZ9eCyGWVbeBel2KhYk/JfUBWeiPwXhXtRt5vDbyQC0/oyO1weEzLrCW5QC7
tBf5gEaXXM2w1HFeYG+CLiDf1Y3ek9FxNU1bzpZAElUvM0DEnDxCr2I9/54ZEbSF
RV5Ppq0Rzppk+KxDnXUu3xfQ1uNatFpfAIAyBX/+1SsYM3BtMlbihWfhhvFKkua3
EzMMUyNPL0FjVBsfxEy47vDABXFk3R4IcnEpHF6/vZO84zfyELxdu7Uoe05HgPHK
Wl3LYx5FymPocE/Z2Ar5ycoqZgu2h4WPkQNCN9aEK5uhWuVPdHa+aWV+QXsKuIDU
OiHxAEDzqreoEKekmX1NYz01AcnbEbOB/D8E5pKbo7ARO+LgfdnuZaghOCdnjcco
lc36jhR2/gP3hJzlsrnPBmikWOjjI5vDUBWY7oVoRoN5ydNKAYdhQeTSfV4bEZ91
sMyYgukLMGn6A2O2ppR+alV+gRQUKhgsXR6WNNy/Duv1KZZHXyG3pHQyMz6P9LbA
iZwMf+/2JU3uRmmxU5qI1OHtac+eeklUtuVxsLdqkLIbc7eBHkYRsPDFcqVzkxOA
uFSJ3twMu+RE/5ZOWX01zsNMIJMFXEdvswXJlSVlY6Au05RL9yAGFpiYpjAI/Vbf
MzujitGN9OhsPXVUbDeR1BJtRyMgxcmAPnqVTNovm3A+u/RlCOaRZMrxDiOomAhN
iylyk/eCimHpOkTMuKPkVCfN+jg9wmW9hwmx1Gv2QzoR6PaSuqeGqvic0ieJkNBs
TMWKTRzOcsZHMkueNyKHlecpmwr/I9s1PxLOGsuP1xnU4xKzlVaFPOZ7BN6zky9L
9zFghKtEQd/2PzfA4TH6KscCGbIc8eoYOpMPILZf3TJP0q7EykrtpKd0P7uFxW4D
qXaJU74bDqeXWxFQrb1VJOPkWAfV3W4r87xv/OdU2z++szPRK32HsFtl5Yt2AH2I
ZEc8cVdpnFTcTfGOhZsr2uTHao2s50P+LkCaCYCOAIbacmhsMs9TgjUDMPBLxPJp
7NXHVIqFz0gkF1ADsHum9aXiXDhqolF4qIgVDAtdyjmUoRW7m9JjKz0/Zt4isuNj
WAehD1x9oBGlS9+bi9IWeJ2l8EsMQphK7J45D3bTKVvF+IAZJn2jBLlmNVOhDQJd
8ptdu7WlXK9Xp7m52SPcAPyXnGG0rMFMkcn+KyUs6Le/7/TQqPly6ifeUmZPglJ8
r+oqM0jf4xO9Se9vjaYcDewmseppWe5k2L1EYuw82JUrkBbON6FozXrHC/w/RmIz
PhONn6wYIjrdAKPNmI+PyQwwR0hu+npi6LXoQ62PZCXRS9oaXe7Sj5Xl4UCweK++
MpwfWcC40RxO2JCx1tVrGHwnPa74f9/Jxgbe4P6lqm5P+PnuptYQe0ziF02xIVL0
xcFDXySJ5ogMci/xhKsszM6xZPvWElbMpc1nw2RAXhjG/P7Kb9LJ+GMp93P2R+nJ
b0eDiLC2otsIH2yWp2gbH5//9uAvVJnZR4T2k22UE+uEnUUx2NXJzTi4Z+v4tcx4
WT08b0e7Ogk9OOTjsJ6pKEdb/8L5HOvxbEm+PoNgng6CBlhWo0Xqqi5+LKK7Lg8O
EpH6Bt/OlBpoDmqFutoCyEvjID+FZOrA2Cg7xYyh6AFiqpdPRqMxRcLQGp2kPIfs
Jk/Zah9jhkMGOLdbcGSj6UFHXo6zKNY7zlUp5ae2cD2w5VcUZ0I5LhZ3Ah4SjAzI
xOQq4axKwDY+Mtzf0G32AaGc60xrgaKXSxxgAyQm4KICJcw6VaqrG3E/8yw5M6Ze
gUWLUwiRgQT+1ng3858iFE2dMAvoYOwrO2U5feX5c52Ai3S+8PLc+LdEa5JYmoHr
e9mUzx1ab6UEzpJbvTMx1Zii+J6I17KS+u3g4l/WqMbsphYw7aNwo0Uj1fPO46Ij
GMwFVBqV0lhwby8Vp9dOsmDHC2VxHLTqhsnGJ6DJqMurK3WTCAq5+2hxG1aBwv4H
pWBosRBCO/ij95PFUJ2sJyr7us7sfRflqAyjIYK9E41CtUPga4w7trgWYWlnlXMT
Kjqb6dG+cXfgygINQfYtdbVzqnfVCIeSO84UnRxgUkHlIfLOfblQuTt/noFb7RYC
q1DOBN0TpUbCs1F2cJAGkCHdffCD5e+Ofyh215aUOr7qeusP6Nk1lhWVjbcVBObt
BOtwjakR4bBaUhSeyjh8Q1uL7Af2+hre2uxC8Qw/Q+xe1tQUiCxV9vX7wVxaXvXj
z+UO6tW3t7im75p/iQ0T5xRcckYs/n3vco6+nvqruP+LNMVqyK9HZWmcnaYKPKOE
8LD7M/CzDju3kgwb107a6fL8znV3f5qyWgAtD4ZpRLHtuuHKmLKudgVri3gYVSGj
7gmi3cDrme1APaPP9T1M7Cl8ATNMXi4V/BNGMCx34US6tj7sRJfoS2C8ujFZ9XCD
YMsaMB1RFJrCX35vKUuwPUZ50uBJUBzf9x4rHxfTVvTHDeXPPS9+RxXAbo8KWliG
5j5kB5gPYTnS5UdwDVviOOfzCFmWKDa07rkhtDRfsFS4ZvpcH1IS+/H3WYyXAk8w
J/4JPBAXw20xmHbD5AaCEVyCkDsY16Xg2vZdN4I04x4wGZoVgflat2wKApdhW5xh
hjn4aWSEafzPknWtQ7j7SZdJFiI5qubtIF50pClHKlOWPIWeSDdFTqyLTfZHgZqk
UlfrVQ+APdVEbh3AV9OAla5a8aNR/mpNMIDyLWp4LxmvlTqgL27uurwbcR6I9Sw2
SbFEe1aHa4HgZd5NTghVjHyKQC0sNLVIzLRUOu1ZFHH8SVw3ojA/Rbn98aG6fnoU
Chd/xq+OPG4Opu9ww9/YKjyg8V7rg2omN6mD9sOuz1R7SsPz37yhcD0CfduneFsq
6nmz9xNFXistsCnWYLAuTvu7pD2+kFFcRAWPrw0ar2WxirwRLjNq2LnTz1webB2Z
a+Dpgqk/5qJNh/+0j6xa2T2tK8KHdzmlRK0uwVrXw++iRSOiHFbqFUhYNqNpfs0U
HZwemBxtrVQUYmQZYjEu6LaT9rT1s+oF3rlARmwBPHgmOfKYF83FSucqk9LobZFX
r3OtoXOuuv7B7ztp+v+78PIspV8HLoh7R0bZqOX34HhK3MZbuK9GHLJVnUsKBoeP
+LBhVdWAYI7mecMxbnFw77JkR7+o9c5J1J1VDjKv7hu1RFmeXTq9YIAFSwJvdz8z
PT1PuqlKBzirjYHDUZEy2GfGlAV/LrYbYBKloAn/1fM55JMujuBrbPWgB0ZV8UqB
fRXS8dSPBO29dEgqG+lVpCYyBmj8T+zEwAwN386GaLD63m0/2ddM/PfmbCRu2Nlq
TX6bKmqqBJ1kZ0F26SxV81+I7x/4AcGItpBXu3NXZhoEI9CdfHv1xH7P5iIHn87p
EBh8wyB4EphM6PyRisyHtaY7kRHcQDYqSTRIUwZIeFhnGW14Axm1GKonhKxpX2bA
gOpe3M6z4phoq9HFwfN1/N2WKKe8Dgr+KTsmOjXNmn+QgdRqSnUpNjUaTyQKkkRe
L9JDzZTP/3Z5nPSPsgL0oSlgAM9nbAbJe5bUNrcxNzsz4zhW6C4HL68EgIvSOnaw
LGaE0qhW/mM5g5CFYD+UkCYCRDK/uH0b8zOCJd96vA8o85d9QgRDyNPf4MS/WAzQ
GfF7yvRkqWYNJOfEQBEyVqBvyCj/v4wUjp/XROcBSAomA9PPEjwcP69II9DH6atm
LzOuwc2bZC3e0AemaVIIz2ulicYP7efkrd1hyEnVFpxxz/Y60dbGCsTcEf9lgft/
uSovuqV8FDNzJubJ7KkI3vCyhuRocjTeMNOH7NAsGlYWBgp3wNWpMkogR9zUAs83
tauEArD0rwB7aiZlKIhwYs/v10VwixRoMPo+Tp+aiveSNKCnkaa00yR3DB17GaGf
tSEO/D7zLotN9UeQrpHzk/jg/93G0L41C8KJWf2p4BDWRZNWLojSfalBuX7Phr2k
M3nEvLCFyie023vNaIck7mNrebayn4+lnCeGjl9zZdqR5mdDrad3t7esMgwFcVGB
Z4yMbVfGspy5/fTAuzDPbvU6D8AzdkVtfQNAKnGlp0mKvXUxb7TgWHt7WQg1ivQG
88pwF77kD2tmUVmvoW9XK+vkHmk/zsxAdTOU1eKl8mAoBw4yUhGt0GVQvvUGjdaQ
43o8j62urrBDTm26D9xdiLyRj7nqF324ran/xr/tvw4Oa8ZONh9gj+CDGxw6zgez
xb3DZi97yWyDBOlmAWOQOlEUOtyM04S1R9Z0aVKbQjU+uG6XhJw+j5/+5rXt9ZCa
bSS/DkfXN6iN0hEvJn85U+g7bFSGuMORwYiOnLDC1UyXeDFicMUM0wzwM060tkJi
zBkqr969eD2UsnVgnbliTQU1v+EFtKXjy/b8h531dhtVDe1GVRVlrwuaR8sGo4og
8xEXDIPwbDGEP0KQNg1s/6pxIlJ9Q2P3fuW7FybTTnBMNk/g3PVt7vSi+tM4E3Q9
bdqOeGRXq6/UYWpsrtcVmNO5Vd4smZB9hrvQI2mtjU76PkT1MIea1ywq7LmTuQF9
L6iYpd7n3wykkTD9fV0mNrwKI8XVBPfXgOw+5Odt5Fbfy2VO/CWd6I7r4HCyyQXz
slKROua2hzQZGm/9jvV/hegU47LZeuu/ckk6TX6QSZHNYAI6N2wKK/b/mkpxDf7T
oT3LPl4X3uw8a4o25fT13KeThgAW1OJ36HXDMQ4TQ9sbBXCL5AF7AF/CYgmbOGDY
Q4ExYAh6YxfOL8RX4GyOp1+F05RzbGGVVozeu28EVZYnXiq3R6Hr0C6xp3zUCJWg
RIoUuYhCTku1oeH2V7e1BCA074c/Gvpc5quygZ85xYWC6ovVtx8u3SmLT2jdSu5H
50/oCoRC5oTFcn6WeAXIH1lzmemGvKU5wPYUpJ/m+Vxa/ctLbhxEO+5RXmcxJRn1
XKRMvHIDZvuqPSYfhEv7hOTVXbNH6OmkR2OKC7D+Yj3RY7Ji2D1qBXJHpzABkzQS
+ubSGPlEb4wq81cu7RvJP3MJ9gZ/Gm/F+HYGkYRsERaLcRXu0IBUhBM99SQoAtBe
APCSZEVZXJ7vLY9EYRrd63qp87dwLmW1Ds9y5fRS8YnzgMB+qqFbWCvipZaaAkuB
xDijyuWYwPq7P4Nt84G3jt/cTQdItllygI8KM0tyF8DhYga6d7daUTqQ77GJH9Ui
rEmxACEhtwfmDO9r9bxwN0RRgQd+DlH3l5vKieLBtjXUuZNbguvOiWsDn38IIkrY
YYFUbLYu64+8/3mhudIv9606fAyf3on0iZIqFp87T7YTjX1/cmisAn+5KcpVROhN
ST2Z83J+kRWTTbwvN0+9V8hBvISLdW+4syyX/0QgIbtjgQZFEOhnH20Kr7Y3Dvq6
t3apgjgxFk1PYJnwA6NTxSrVS/JNyv7i+YzbQLpkxgVH6zQRdc87/2bh0E4evWI9
m5FTXYQhECTRBchRmX4WWWlb8Oc+l2kXppx1ADhJez4UZ4alRMsjY9stQ62C3bAY
js5PlwL5yiobskH54jssQAcJH/x7AiX7IlvTB1ngZuWCiN5dBxQ3TfW5l0OIoLi8
y7w8A/XAuX/J98tiAE/lKF5QbpUY70x4rTiH1/x5pxIL9A3kI19hPQDrdqEDuHOx
hecoLaRfzNr0ikc/Vq9jWNlsN9HtOFdahX9Zv7JpZpnFunqe60mXdA6rJxVOMQ1k
iCMwSZA50Q+XGVJYMytSudVssEIhcgUIS6sgBL1wRFXynfnLlQxFQX0q8Kve9oB9
R0VrcPb4rFuzMJADi3k4YrT52+ldhWi3dLXxUQAa9+43wy/0pF7k5lg7gwby7Z+1
99YA94RcxmI7B5xp6/2Jlqk37nzme5VFtiWv3oi9fQjdK4bdLZtq/Ku2WOyWRYK9
PCpyPezBBw3YGs3cxAlu4PvriDdQR3ozhF5xnI6J4shCgqgWdI53MoykHRi5e5lv
jkbh5t+FkBNDaoFI66IhXu1SNOiH1g25q+X0/WUH3VXoOhE1P818AhmTZHV6X5uS
T3CEvBJoMHHcjjK5mUvBoPNlfX3dC/8w89Ps/rNdXVePUKJ943YYNzt7hIW9qWWL
AyGwLZj0OhST33cnjgauuo1s0rXkL1zXOBY5SVxdeJhWV+by6x4uQ0nLQ9nXUUyR
/ooWoLOFjDgTg5F01pd9rhUGNY7zHW2s366UWt1Rd4WJWmvCXwwVkorgvlLzZO5c
mbt59ekEovymXQjrYqw16G712u+ufQU2FXi6KCoYTlQqsCwnb1ANhiomboFikq6x
+xX+/pKH8qhnZ/UAaecyGk7XhJhEXDNnWTb7GZK48ZMD3BjsqQ7hFj6rc8xYNaa8
RL+y8eKCnbYgTsiUMB8yrAETac4syel4P/p7C07SL23IXFG7bzxpDkrCLRWRErwl
r85foSviMoVffUvXWHePJBPlA6zmgE4WFOfvp8jUvE7JStBGBWxZi+h3wJDKnWgu
l6uPB80mN07l5AmpWsgVaDoTXWSeDcIsn1fZIkTUVfZ4Vymugq5BjLyuadJocFYm
tKRGQMoMwDs5DsfOu+9lCvY8os4GL5/yv6oFjW7uBTSWgRlwkuVBnObHlDc6XSqs
TznR2MWJjFhSHH/PTLUYRDAMIPVLdbqS6PR/hr0e3HcxnGNKFZzynxnuXzzluoHu
3IUc2ocUOMKULIMoxyfpeF7dNzAorCZm+W9WGoNGi579rrxxN7x4r2I6/R0QR5vB
enWKphYNBpUCM0xfPIqF57rY4A01gcgZRGTMh4YlQkcw7mX6mZ3TUhvOWpr9WWfb
2to9u9BODiZ0LlRiOHc+BAZ2zMcPs+alynb4g1PI1NvwSmt7UluRA0CreZMrdQTn
hA4/lYXRpK6uSQct45UaeT2ANFfnaeJWVImptgaR75DlG3fnRIXBOU4O8XQLgOQH
oRn7mCG7C3BYLIheJZDyIGY3Npyl3byEZkLzKN965Jr3TgBaHrduQeJDpmGlb613
op0Va2vjOrmhtSoSqs+WkjZvJtVM2OjgUfeyDw1x/ERG2oh1Y1meMocvE1gx329j
YNUcnh1xKCFB5ap3qbZEHfAJ0osMHquQT1/8QroHiJBJPqZZ629Vc2WVNdUr7tFq
leAs2d5DtDGw3CGM9gdlS+1vg+kp5qb+sdW0+7tUVeknuXOoRU7+TF6TYw/SJt3Q
3oydoOsjiTA1nnCUOj8vpg4asrLXomQ8Dwvl2mKczdB7BbHq3KvfpsdnwNJotoJv
9RfOyvwzMaTYsRRbexfmoJmBFNn2sXfPg/5KMsTlXhVfzDyHwq2R3Yl6DbTSUWLF
hHgA5m0GDLJcoMYQFbESvt2JHS1GEDrwojIjuxSsL8SteiKzWVV95ArbFeKhRrFO
MUXBMXLSsMaMEvacl6LW47zc/hms+IOsW8rZJI9ZEPcCRYn3NjC9VBhBaW97w3mS
NaSqjvVc7u3F0s4I0HsIW6tyjdMDagplmPoUkSolbXbm1/cCAqrZAhlz5DiAtLvO
reOzKn82F7SSl7fPCv2C85mfdVbZKX25AETbGRs0MkWvKgBp1HdUx+Pe/lB4kGlv
/PAbmBMK3YttNxSIOuA7L1aJo2l0ZBU5E57v7Qsx/eeKfO8QHzO5I/t4qOXh1O9M
MGy9IyB4u+GZUUgDuQyz7Lot6pKeRudLg4BPV7pzn3FZ5rjRDo3BuN+Dz6r56C1p
Yx4gdQq5La4pxHulfnXiRdG3pebvDput5kPkS9AcGi4Vq156ptfTPvO2vi1cdM6P
8d5oJoVbfW4IreJ0GfnZqJNgwOGr+tfP18CBkB3cF3y6CpA6+LvLCI1UY5PadzC8
DYYNSqc0H+CJIdIzzgUL9QP20n+It+vvAfft7mEe+Qq+9AHVfURzDfkTrEgLdd1H
c0PDc1i2ch8uW5GNdPflKGYt6UfgOsGfPgbuYaBZonS/onZo8U/KbLMlXjcZTvKN
XMB6yJWEds0ZJfR+IOSQ7WqimniYBoU56fa7jsaGFM8EC3KJHQepg+6EvDRnztuu
f+cu+2yJGe4pjbxGYya+zYZfaSnMfYcHDxLriYhhd755VMUDqCvMVql729nLmWqk
Z6tE4sYUQt+8TTjR9kTbdmoKvSBz75fitZldqqHv2dULMRrFUIdaSk4WPobe6aL9
xJKzVCqXtTZ3WWtNurufdn76YLdiPh4CiO1zna4FQ+uT46fxGLkxruv03T5Bujbd
JqeZBDn0VsY0JcBGCKOQxjS+koRr1PUuOCyuf3R6xZgTd3YqVR39W6z70BK++W/4
blPU9Yjg+H/qIn0fJBVuxkrB/qc2KLqiEDL3EvtdfgtuVOg17vfRHKKMp3ocNGVC
Wvx/u2I8otq6we5SV+BuABv0bIQfY41Ld4gToszvmuUrut7pbFdmikuRe+/d5/Rg
w8MXypoWGu7wvpHURaE9AzYCCVgrK9ust1Do2UutUClJ/83vZQ2uBr/cxZy1E5Tw
Q9SKKSBz0z3gMtlv3pggfIvAZLjVb+Xr4iiE2Q8Ci6shKGC9/JcD4uZn2eGa8Fbu
Z5oJ1Hx0voBGXjJrlMDstk4LGfsyBLxjuomA1O24u2iLc5ERGOY3JzxpXPJlQsJV
CbINvQu4mhRJPQ3cRIIB4ji01I62yxUTqvm+Gzp92Rs2QktFIwP+c8aVvq5PmMSv
oVFGjY8y3GCCe4AYzh1eZ0QEdPeA0C361VDRgRcjL9jexIgFgtX/JcgVnKdpmckn
91Qrp24oFJgj273CKTQkNT2iAPrmeFZM6clRiF3wS9icyF6YM3GlTxlU4o1qTXD6
zG4NCnckxkNg4usxEcua30hpdJdBLxiYDkszGRqSfeUDyv6n/btFueiTvXOuv+/f
V0XL96Ch2t8aiaO6YS7W5gGy0BYiwQwhAaBP3EHu1pePcZl2ik5mtV/lOEe/SIHS
9TNw6QkLwRbcw9lOGfPOTgyzR+jKmKHxh/o3XmPtJP+A3+I/CvbdM9DlT3jCl9t4
rbJp4gKZp4M+QAicS2OSmMjThkz3Ctt4erq2+I2KodJnedjWMt/GFIcUR0hXGfty
D8DGjTfh677IqEaUrgTEjzSXLgSwGFEyyWyz0fECYGpaoeB++X5cJUAd5AEmYvgm
M2UWNx4zveL86HA8CzXmOrgaHERHKO8ecwH6VX0O2o3RhLFCZk8jqWy2HyxUSbml
/GmRU6dTcYbqlNWJqpN1eAo7LFn7BQ+yaxwF0ck7JiT8we8ZKHE8OvsKGXvptWcu
vhtKtl7Gct1RNkCgN+fe1ftvDY1VzpjUwlzrFG5zOj3iqoehq2BcLxRp/NVGq5Df
Clz67Fuwm0KmIOh3FKsU3Y2MNTPR4k9bO538p65DJ7UNW6SQ6F35AR92HAa5VGNL
dr5fiO0SH54To4sq33+aiqM71Lr5kaVg8OlTMSxCvcXsKbvSyGClzJEZDOsN3tnQ
JedGbWR96RrN+A0hIMp44270f+kR+P5itrA7ymYkYZDtlWKAWYerg5Q0MKqKyivC
kSppsNivGH6tp9ahEBgW+3aOBKjei5QGas4scEilwQzGerCyhLkFVxXMd8B6gNRF
fhGjP9V2ayZJxM9ZDZRPzzSvlMTLvnw5nx9TfZxWwNJjgN5NDkWrHsMDiXJqfed9
lX3fvQx9Zi1kVst2UZfz6aTzzIgQfneeEe4hwNpmtCGlNqgsIc2xm6oNWY7tJWSU
UgIm1H6BFgwtyb6uFuNhVghd+LSLa0M/Dfviz4qtKM6w9JwBshwWJRXEwTFaXEiA
RW0vMjFTV6Ho9BR/xi3DgRtHgdKJqiIsAM/3VqHMotPiKrlzHYjlrB6rJnKmeuB3
cM9I0LBjlu38XWOe5lamG+gQEJJxs4BVmefzMD6Okx9sdpA9fdEBdnTpmGf9vd0K
dUvFQqa0lCcLPEOx4D/L3aF/nFXSi9BW6AUe6fvoHWPBU018NYe9oLXdpJZCDbnq
+o2MM1dwS9ZbmEOnOEPDb25FNPJXzxkFqCwQUoOt8k9Hygh/rgVVb9SJMadRx/pE
XrhNvEn6jbgz92EQI48Z2lnFW/yn1/Oe6VwTVGgigNMDvDTee4j3olnO+9Gxn15p
8ZiT+9QAZAhyEfO9a41UcKYdhiFxkvLRGVlBuYDi57xkDxgJNt8pl2pZMqLobSzJ
Pe1E4oE0yXSYCOse1Xx494B5XKTGyiZXeTbkzHsiCBXyHpTKaNinNtAKCt1dJhjb
bhMUzVabBCgH8n32+e5nHnm2ugqVlMNX778N93GTSWR7Y8FTU+FqDDcJxdqX2odZ
YUkJ8hFxcEoTp4HoTJDqCTI8wAueUhJX14QL2w49QAjysDRDyyYhXqbjU1KEwrCA
Wv2cFASD+XElB8nMOrhwICpfq6RIouktUonjK9hi7B1jDw91+Tp6Ks2sEOfr6M6G
rZHvyKlH0vlR5HelUlk8xs4feXZlIHJtRZtXV8Lira3O0+bfWzj+hQ9OLieLVkDs
LHTwzfxWPk9zy5i63xKiRHKcQHZ0RbVr98DkOh9j0qgG/CKSLXnh+mLyym4ET1iT
urQkkvI5vvdqwiLY4IwvB/6NG0mIatVGV2GMHLOnemJaSt/r7RDoygOP1aG/xTIo
i9lfYgyXGcCvz30RgEAb91x5HHWERWB5S0FIG2ofUHasuGsAZYBAJBNInbAQd4y6
p9rR8k03DaRxptgtevpUZJphq/d05EIXA4IFvmxN72wK+5VHtNmsFxHlEqPFHzPr
meSukFXtkpsjZrXfDgBXcnbtfFCr1hHZH3lbeWBQhrBHefbxsdxru836ws0UmzxH
FXZwJZdfkLNgCzFTPxFZKUxvj1vj9AUThvKExvynwzgdnwbN2M7iIqvPDgolr+ZV
wYlDLkzanxC47SYp37E/Ig5BsHRk9dhrCJ7SR4nAXwnrQd73iZ5XdhiwIceJEUh8
ay0GMYDpODIkjCa/paVg6T1GQk3Vt2PvbXcEbqkDtDydYKr7Q3N1fHEEwNnYRkEq
YUVam2l6RgQ3nkLv/iHi/Uw8673SfqDr/GPBK1YUJcviTgD+OrohYOuhF4n0+4V6
e/j486S5VsV+eCohGGQHgv/0WYkmbrDNbw2YkDfz5XVf86xajqug1BVsaKFjaRxb
O8pnEL9C7pSew/xBNsTftA1EShn/i/vCDUN1qR5FDo5dUIsY8rQN+y3DkaPl/q7P
77hIX2Uc04L+BswxEeibGF9Aoj1yrSywEa4goE+DdVNIcI9d3PvYE2E4DfogTKcI
ls1m32f8TrQWwVY9pDjfWNeWylV30VXOE6ngPmmeoWwXOGE3bv1yhzm2mgTBmZlg
MWSVzh4vAJ6VULFXEtpqXhk+22Mx38MInXu+ySlwSO+nWrZdYKGt8n00e4AwgtKp
8F5FCf8YD2ByhM5YQJNhcoHk6iZXmd2j7O8Sfi7N4c2ss3HFdTMDFeZJ8mwI9qP8
fRpgM5zPpZVEyWrxAso6h7VD5xbUkxiQjHOeshnBbQncjHvr1O5ssnZvDFRowp2F
ldBQMECfN94KFJBD/HtXoc6isaDbOycFTFU9jKvk+u15zUDZNNwCZHq0hlrtT6DM
BRKfoTkIKKqB237RkB1lU/iQ+yuiHNRyP2jDn2cDjy9a9mHC3UUAu2QntehmivAt
OHR4WmlP14NjOA/unw/piL+5XPH5TqPLJ4YAzsNGDjwc2JbO/QlrEraf6OrIl6Tn
aoWE3e5Tc4wXGDo3OEhfgKa9A2BTJ8RsPYJmFe8d1u/ZOinKy8VMsprN6iYwRaeT
ITLe82GrnZf+5kxxbzeGvERNjqCudwINi4hVfi52yVzVt0/n3vsROoywgeiodJ9E
aFi0zKiUVO7Fl1NheFxCe3crjmruYb7eMG38g9OeEQOWDw0ISSDvw8TuLE4c+2zL
c4BK/M8j5PA9Qmv1ltHyD40/SOUlOoobL2v4Hzo8pQXIKTpf4NBlTzfDRlzBQXDS
gMGaTlItBl7z+/qE2ZCLXfq/HdGmyoGLfx6skeafCXpNTYmskQU0M75Pa8UNr3Fc
uZvXEQOdfTzywNbHtuxSgnIAsPmvM+AUMJNvVuM6wzm0uxZCgXDElkbENTMI1BFY
/HxCknglqm2Pe48FImxCrYfj7BCUhv9DaOC2NzDF4grydzfs7HVCK1Pi4OQHL6BD
JiKnI7OUZoJqvmxSfhw5TvODitx5APfpTv1c5sP6CwN9JMlujCUMefweu6jmW0uK
HZYuWAdxbH78SzHT7l86zXgBl+tQI4ev7yLypoeWnFXiCENBPv26oru/cJUV29WW
mtWx0J6WmvoGA7iayF/6k3VcgHytjf738KZeAgp35i5OOXnggCYvcF2jR8uOW4/i
pcT6IYTN/M/dvIL1sisOHIly+qAC+00VYpClZJUwuBiQT0zynvdmgbor4ZTKiiMY
HwUhX9vOI/DEQTwSOrkDhVqU6F0RbQxsarGfCT5nA2ubhmp/rTxHYZxA/U6oKP9v
fDBgS8Xwt3FSzALomDDRzUYToyOqecMBvBVtUqvq5Wf1w4We2t5koUrEdRjZlxl9
0aVqPflYcLFrqsvYGaV102us8HiRHC716Dv8rERRTyyx7TKaZ7LoO0leRrDouWB4
gBiQIn0Zh6oGLL9qIwObZBdSBA6xplyzxAxVVuFNYUTNHXqCEdT2krsNnrmqINGx
x4nPQ/l0RQTkosL+L7xLjEpV8hdi3169iJIWaOib6/WwAxOr9wcDP3LwIAOIfTST
AwC2GqQl5qYBn/wQhjk+YjUO2Ev+YcE/pQ6BgcLQ9+wG0wcfRlm6Qndg/Si6F2fC
GICYUMZtvH9/4B+pkOQDndBM+mwQ1vdrQcs5H6yaJPlo3tMpby7RCIfaTDkS3k1V
KuqpIx6Mnuj87XHvPLjMoW5VKsjjthSo/o0Y9KeYkO2Uv+eXFoi6joL1VHSmDj6j
TmO1ZbUR+mLE2fhxw2ILiUwwJ8Fmi5Qa8RgYOEPDH/o3FnR69vj2JMk1fTjjnQkQ
UYf2M83QyyN4qDQMsdObySc4pD4bwVOnGrtqEPJq/OA0fExaUA9Xiv801P93QaXH
HJrnOXgHrc6mytqKdKNUh0SICSdq+POOzWSsZZhmqTSN3x7ZOx84EV2AHjiSdUlW
KwqCoVhRJZQJOmaVYD30NNP8VqgTMrfoLQvVKCCmeOekdKggvxIPNfjYdbdTGfUt
gtytVpER8eBX0YyYMG/B0hy0iYN6JmQNlL0n09JtUrRT7rreCJainIVpOqzzqHrO
Dl8fGU54zmwC9L4zXW2JRlLI1dj1xXRLrFK8Nqi2u6swl7NmOlkZpaQeMTYlXjiV
ygdSMaVaFA1ixDlUwkhzAXMmpV1wx7EQLGztcaggi6PRNwPE/j33+s91EpUzGDoE
+kcglMd8mdg6RzqoMK2ibUkuuzET9CBprLlEWDIJKB3FYsAgpQGt9lqnmwdY1+q8
ku1elLskcf15V8IJno5udy2Fk7sTJ05CmGzHBriPDucVoXLS1NmOWycr3l1b2Uyi
Y4hQmlGPyqQWIvfAV/+zgd2wyJG15hFuaEpmj3U5YSJ5X2CZRTyl6/YLqCDQdxk6
5sssw8GyBLPV2r93M2iFqqn4wLpDIbnauo16lzseIwrRCpzFaMp8xau3cjuPOjJD
aqhZAagMl5UhqkJ8QnIysIrmXtdqW4FWR93qGuBETFDeGuGp5y8Go0L9/awpqmoQ
M25/uFIVVcv4oL0PAxm23YmB7fY4Y79VZWBnjBRnchjiyCpFHYBpKNWsQN/QR83j
n4mi0KFMsdBEesu+PR7pvBJ0T92XFHpm9zSVDXHuExDG9jXgzsVduh9Yn84G/LMh
tPWvBNNGKdnDVygwgpYoQ2na0mY8Daxg+ooqaa85hgGXpgzOJfjGtL0pvk8I3BIP
US7S/mRKMB1o8NdiFMx1Z2/wu/NAqDFxBwpOJpTgtS6Pu0XjDgt8dO1wXmIwEyyk
/tXgPFz1Gu+//fOGaW+HM7W4Ts5cKR/oVdEwxE4i3N/Tabyu+TGr6SHW7WiNfg4v
V0oTMnKBngSqep+oEFVDp6X9F14RzsWvwy/8K14Hgmv0kMf5FBmygz9JZuA8N5eu
VifBJ0ihO96+NX5goyMvC2cn2gdlribbOIesFVDDqOSnt43UUm8YQsGK0WkkQX6E
l6MfpbcR0zMXxw7CF8+eep4UyrryMrB4Le8ugChbM7zlDF3lFaNOoVKw0XaIjW+t
8svHgJMSqzvtzZgN3CeoBAB+6jEB1CAQuWDFTRCDdf6Ei9haEnE1X6f8QnNTdZmK
f/i47Un+81NzBEGf8CJqm2sTTwJh+87K5ZgMfqOvn+zYW0jVMIIoyIHRN+DI6ao7
4q0qM6/G4pt+/j6o5ZV/L5SrC46Yp0OBVzUmZ3DhDZialnPphBY8W42LqWcYRqaM
yvrfQ3p1nVjmatt53hWJBzbZ2X9NbL6rGg53WlTNm2zLNRTsUZ8qLmwuVUAxiugs
srvM+RwJ9Cik5mm7AdVgnFJLXu3qg7aScnyGK/gDsZXq6X6in6jHmMJJNMufGnUt
FsPM1iQgxEK9EMY+97qAC9R63rOMy5ClkdUbG+n53KmrrRWycfxgtiBD1OnmOky4
EhDbJgs+tY2OiuPxiaVKxfbPsKIXdaDqucI80fOKHOSj1vsNKV1nVTMnh7wGJLxJ
P+sLY6LwAHvBJgjs74o+orQGyXuiKXWHdolfDxYfbwgkHYxYglCUzgPgg3w0Tf4H
Pf9P0KvUXRDzi/D6rCk2s+7qNKse6cRfBNmIlb0B3LHvMsbXMPInClCY2bl9bXfb
T6l8b3Xy3BCl9kxTeuAkMHFHppYE5W68ZzK4m8SLj/XGgAnoWPS4VTG+QezTYjMG
qRxjjHHRXUF2iSeEdFtQw38IqPX3Uo/dmZYpaNV8NdGKexoqj/js0vfgLAWfXK7X
VzeuZfw5Zfx95SWAOkxPk+FfjC/VWXQnKHzJ/1EXtcflBAC82rhZrSN/AfSMPtww
Em5I+FLEHgSJUO2VUP6B2j8fTOmH9fWHRegsvv6+u8Z8nB7EhXc7/BWJXaXIG1eV
lgjaglDeCn6AFD6fCQwcTI0FfC9bEqRBvEDRtgMj1xwW+Cbv7wL6axWAeKscxo9H
V6u+q9Ik/c+q2EooeapKVHaw1UAnkoYLw3GBOHsByJ1Zn7QrgMfMpU7W61kdTWdK
D81JxTbcm8utC88/akQVJDfzDPRJfFk/3iZiiUafCZxXAn9SSl1RzdzHHk73Qb1P
QCvwriA5Hx1zgvRkgFWHrsZIgw+4es76g2jE/yKwly+r0OaeNdLlKQgap81er/g4
lmmMXaPccpmZ0opBoQk0CxOWhY9LfMLXw/V7Bnk3CIEHb1Gb0IueNWSEjr04KOc9
qr/TXgKKeeNuqjyiMVWFO0w9sWGR9ZtA7RBPJXOotX8r2hIlouA0NUKVJ3SaML7O
YEAw/ze4Wdj440z6SK6sG9Gh4mLIhlCO62vvbA6SzxCi/bERM1npb4nBC9FQSV3v
b9BXXL9x4TCGVuejfeHhn2np3vJirAHl9vYPNCcudC+TIIvQNb5Z6vYInxTnVKGk
3sgiDAmXazIQfS3d5CZmbICSyQ5CdhzDwVVVyQQoXLCIEXx9mnU6gs6xMFigV7D3
Hz1xjcVaBniipUXF0xWL0hGBM/UlMEnulGZ5B2qn2ZdQfddDffeMS46E+u2yFzEx
VTIMmY5CR1n54O050Z0AL4YJ9QQ7V38VmWJ51gxIn0jKFXafDDwE81G+77Kbr0Bk
xJkdntMlxMniC5lcxrp+LLYo59mo54vXU8Lv1/jNTSSy1RMF2D2TAY+ARtBy2n7l
OF+5GohRM71dDkqXpROugxm3Do5nwNi4jMeFZfXW2jQ7vy6FwTLNcNXqh3R3gDk5
2++qskN9yVDFPmoQ16EQnrI3CYCDnU77GOdZBVWdT0K6r3J/ookF3Qy9a6ZjSOlN
gTMhcYfU8C7DBbhTGopvgSIK6OFaUW/DRCIY9fM8pqJeUNvuwR+QPEenFlBuPj0K
CCKheAncCyusCSQoC0ukulkeFfE2M/P06t5IaKpZaXFHv/D3ajZbXkQsTrvARQJy
8eHInB4g96rE1vvAfnCYgZ8CNwuPcZKOAepp69Wci/MESqrfmXCe1U6yN8+Jt3tZ
0rYOxySiP/q8NnUuPxxlC73KT416fn+NvDuCEy+eywvqYq1M5QusWrEpBrG+wY5/
ebSv3MVRFBFmUtoPtBLzT6RKA9OjNMwCe4zXvGFrd7UUhSsC0SavSCOeZYUDV4Rp
m2BdgcZkXXTGbisVzLyPf07VVfk8ithz3RBfJ4ropMIk6rMKp97PpSntj3kApVLy
Fy68vZusYGobg0Wd7yo7XkWfivE4hH2HP3qlwlznrBWYjodud6sba5fcLFBPaGHY
c2zSCdB8fMyOTlnn/1MvAelonwvCIVimjsp1f6eiBm/FeD0e/Rhxb1NUedhAxtOM
55uWWuWkCzIWkdMVIzaCoTxzApIIhmbYMxMqdtYKTWAeJOssR0a0wvISsuz51Lfh
EKMyOm0V2KRlyALLAzbqAFUg2DS+2K6HYidqIP+uWRl6f7yEqL1T9OL99DbOnc0u
jm0ZtHSB55OF3arRtaT6q+dVStzhD4sNwQnPE3nGf1FDwUEk/adtgzthWdjdHuNa
4D/L9HvkCfz8o6X/TL0NKh90GgExC2Qclgl5bo1zegeJxtmHW52nW/1hpriUhOV3
39pxlwwP5TN5Uqn/6pOCRfmH836zO2MVl66oPnCE5N9uNuvwDkxwfyirNREhPukM
Vm0i9QeQ4+UGZDaF8HxfqDzDrbvwEkIsrIgWZkT7rPOAmaZG9mie//ICSV13ciyE
35n6v8bN53BfRONzw41+hzBeJ1MPRccBJKxWHziWYGpNRsKM6pvptwtn0OabjGO3
7xqIUddq7DC0ri5tAn6nVVdu/IoQ7BpHk1MEnDoa2ihdn08G+GrAKFuRR+yoWQnL
F4B3f8rijEiOdS3LiEKZPNjzmygmaARFJdkHLup3myjyEHW/Zbr4OauXILHuvg39
OyFIFTxWsJRbW/YOR7kJGfvtSCQei6jmyBDzzZmxvJhA49Ztq4ogDY3WuDUEeeL0
EigV4J+t7LRd14qQds6w7960wojqHaEEf6rR9g2m6Pvf91mBqY9eNTi5+VlTSs/S
eB3S3PnWRB/odxa2zd8Ln3bBuYp+55tklmZLFljge+PGMNaquoREK2UqVFESg76e
RoqFOoSZo9Wb6HoHFkUqxSfZvUkCzVIJWoQyQZznYfLX8ceS3bXXPshgeqUbllR7
c4fSrUyc+UoKCQDWOj4D8EYKX0+xbVW5HdJhIA25B3cJAkm8AnmUMCtOBJFai1p4
FLZWorbv6ZU0d4EFqMek4+lZa8u7Vc6cIuUHdRM7F/M22zfMQcANgJ+3xYje4MbP
kPpjiy3HVnZyWvM0SG4t+MXyd0A4P4l7NCb+8tS9jrxbNxgUF/OSJ3IyrIvza1Cj
WTTuxnjN5qzwZrgSrixAFcsyTIprzaO0sISlgoswbtHhl/cw+40369ObMwrMIeYt
JOWOXOh9Wa0OkUEMSClK/v3pvkx6jrbdc236r94oPTTSot5Ogr+FOb7WKP3Pp5ds
2hezv7dhz0ZMPswQ+CWbpApDWqwHcOdt81YKtcEv3kNKWY9R4AGy2cgO91e6r06J
gKw9pzo0z5T7TjI8fkuqsx7w/jCHfYXQ4ttTjawY15he68f/E9gOijawir10eHwu
FWOwUt52m2nCvGGTVa+UwGFvbTVrA5Wwtszown49IRkAU80NY1oVcCNYBmyFGEam
XJTJSxHPF9y+1z9pVgoy2RDj2vx3sVNrzaSHbt/dNccY3lXkSRbjFv1cUzTYHYB2
KV5dyC1SoMMHB0XGS7NABPa9dwjTI+5siqim/bjgTeR075HtIfxL+pSD/bj25qfb
Z7av7aiGfxij7tzwNdiMq5brasqmlPT/H9cNXpgOQDYchqndzCDElHHUF8Zm975D
o/uxVNzSbGiqqSoUeLiW42aYbjwoVSLvYnli020VrR4E6kcSD2IqtJf27bbO9+Pg
3sdVHgHb+Y7s2xzIMG5KALTnU3B0haYX+Lj5BFZi2chtHYJAMcvQNXVfqKYkM1Zs
lpYx3KIY26bPnqYGVnDiNAs63VS2zDkeNKbQdkeQBhQOGIya/hamwIfTJ306TLA5
68W1L0jS97Y8vg7PynJuiNzdouLKGgs5BXHJHvkkERcKiIJ+7NxvdTn3QJh4oBtN
3OgUoPlfv1xNI70VuPADl2QR93jiGvWf3H4rPOEY1tisxouIb4iSRJhJ+ZhTkZ6u
SQgOSbbxJYGxZ45TA4JK7mkqseNEMn29ECSaPCdFF9lCZbPo/2dVSBH4OmJ3E0eh
IOs+HGP1i88IIbrRDMCgNoMe0ChOZ7gsvStphUhotQKImC2CpZ+eqt4KaPaYJpU5
Ny2aig1Sxprr1x+kOBPML1OZJ2KX3NKuEfsN+R7IOqtRqgO/h+blAvTofZHvlkRU
d/4bYehm2EPx6+QYpWQvky+N4oereGPNPYsNKdO2xPAuMI1qeQ764xgrx7/KZ1OB
2At3zPm1uIpgyN1TU5UZB6MQQo1EbwftOjX7t4fZAW4CI0c9AX4ISXaXSowvQ5fy
sU6SuMPPJPNDSMK1SC3vnc3utYtE2VFwAhstCTEKrPryCiKlxmoQQcG+x9one7kx
5AXi/jayDSNNJ8EKpQ1bIOWlbBN6grFS61vqLuOAksNUipeD3YzN7Yw/2aL/Rsz7
PkpBZsNW4JGOBaRtscciGfMqwthr1657WDqO0xY/VJOLu6UKB5BH9CgofskcocNW
MpBLipsUv8a7n+g3qkYms7yYwMObL+qFxTZ5PtYjEy6OKFDws2u+M5ePqu3a1JMI
sicbNWoxIRa4nfhaKhmtCn0TApdJ5iecb9PNougkmf+SFNmMHfHtMegSLDoEyhh5
mppW5fnxQe5t3e9nQJWSC40P8lg7ULYqPUUsDa/uZeViJIC61Dv6P1Wy/baKDHZ3
0GgZ+8sFt6MvIZss6RqiqYaq5orfb3e/6RdxL4Zmux5Ro8O230rQ85B27bCLp0Qo
J9P7VP1B9io3Qcn9lAAi1Y9ZAEwg/ZBqM2i4FWIUyPZvhPq0aOux0iF+YkvtmYAU
BzX14l15SZ6UVqlP9ue+CS+w5WqmZkVlO/VlyqEamfqfVT4lN/3ESKq5eUVQ5iLZ
SsjwGm6mlsoFswFP3Cen6AoE4O8RWNClYz8O2fsu0CrNTTUuAJVUB2r0AxD0PKKb
XzGekRFtcPFcFNvLhrOmqiBC5H1ohV69V4SSJIu+2Hl0ht6HYRM7ZOzqAkiHFKZW
qskIMVr2viqIl6Egt3ZioYXbhSi34HfgewmDERyn4ZMgJ9F+VGMGChkcKlMBhh/J
+CnC2WGUqyRh9l0sr9gMoE69AEW8QCO0gd3IVgGk2QENJ8f2HsrqHQQgYuwr8TgJ
Y+qpsvi6R7FnINL1zOqbLchR/A3aevU/077DSyohzzdz5BSoi1KFx/9pOpBMJHhK
Gn//dSRPksF8ATCY/RoCVVuc7Vt1HkfKmbQSYau67r7911Vywvvxntc5Y6C2KyWf
d92tAFzDKCMnrtyzZ/AqndxdLz4ciGtJlCfJeYfqrf+vOf9tZY5E9G9+SpjqkA77
3kv6dnZSJN3PYPH4eD4Yve8dmw9dcJAXjlHLDVaEyxBA0NWVNwYHdCt2ATfkobSF
PqFOpZJG3b32+CVVprl6ugFiYt7GN0kwlYULv8WNaQe3gMsZGsdwVRnVLzuLOm5i
AXp3oroTF65129QAR6Yw/WaDYukZuMMUq0iZnsr4YlE4+Ll3pe0ZiK4AHzWvxlx1
tyQRwMcwMoJ9t8eeqPMq6bfirrh3Vafvfje0cYeL1jCnTNt1J1SUVIE+A4MD5D6M
D9tlYAHZUCYvYOf1r5SCxfuyFEF7OZdhbMPAMk5ncW4fCJ6snRzJ1H4BYBK5YDnk
UzYkjPGBes6LjbPiY+D/o1R1biyJwM9jAKhaNM36wHju3FKv6HEYkrfMqPDCy6Bl
C4RFfhPalGIATql/RnzNJT13aTbr2dbJ54XBLF7pkD4GLkRxyyfKocc0oWCPUqld
BeR7K+vIVfG51OGmCYmkIf6sBKtzHV6Ej7NKlGUwFH22rCFDARP2GEi3GpjBWqej
b6/0WKIJnt2wzWTDYKbwUj7XcFEuMkH1FhdCXgoXIAYIqXpfe61qcDRopGJSJCK0
U8yMxzRNw3UDqLvbuA5/HIL1X3m5ufjCMyG870OZ94xDNaqH7615uTh5F+RrSM1B
pb1zJZHah8ihbfQy5V6jcpyAcnAWNo5wq48eJgx8PADr2YhKHytfGO9JVkKk81sx
qM3Lvfoocpf9GpK2ogc7eG/DSWqvqYPofuSPIFLVCltPqeBaNID1h6dg453gPanz
dbyq6vvOeh+egHU2FGQJD2JHzftQNGLhPBoimG8sf1EFAlkv20IE4KH2mFbCmxav
jXuBxyhi56Q3ZimH8OIGxl/PaPx3vKnc8L8a1g2mWdbdj7mTpfqET+UXwt4GQ22F
5oATjcPOUKy2cJwuu9nWihsqWjjtP3nY9EjxAptJIMJl1p4kMKz7hof/ptutUR1m
si6/5nItg17LTC6aE1qvPbq765CUiDu7fzp+xSHG9PxQe7nRvXhBAiffxbit4rx6
0IfUmyIWYj7baI5Ugs7oPFKmitD9Iy24yhJJv8f8yYhWyuq9hSeYnwZLRje+CatG
ttXvhf9WpWHSupOwbMTmsd7BLEZMwJYtiYpkNNYdijVR+49ZZBRr5CA2B1iuSLAB
EQ/h0CT/KLyyWaEjrklnVfZLkLXgpd0REyyktjRpU9O2LrurHPm5OuJGRDERiBCW
aGlc/kXtHm1+SmG4k6hkZLQGJsx+COQPIiyLVZRpimiFpGUw/AZD5oJAxWO0+u/S
H11YRnDRqfSVhBAvs2ujNx74ygwzKiEX8Rb3jFmnPrrRqvXjrQ7+pa1AntCZxi7R
FkBi1YDmtBKQAqAZ77jDEh4L3DoCbFx759d2fadQGMSbOLTRoBfUy0EodYG+a8l+
4+bEABh0R98iPCbVI+rP49OFAbqppdM4aNjjVopqVc7cIb/Tz0E3/ntETfXcJ7a7
RRrgwz12TGDuROWv9Q/t6kvxA5OZrPk5wPI7uaUCTQbJZXfkcLg4MZu6QQ3bW+Y3
LjvMcGsHcynBP89Q3YWjLytxYu7zDPQcnSAi9wto7ZMYjQUgNUGprLGrw4sVOhpT
i6k8SeGA9oNOlg4eAz8cdDQtbT8bdIu3UKQZeqqjYa3nC7uZh0x2jG/L0qGC1Bl7
tAskjlv6qEFnQTSrZJTXKh9iBNZYeU3z739VNhQAfj/DqBTSA5ZpZLJxJ0eOeWfk
JER4I5Ow/URrbI+7yKLWN+wWXVQEzuOmzhg9lCJlQM/8cxUGYwvolhMXiZG+S6L+
Iw2riP4BxGTY8CSQVfn/w75HtI6uyDNphkpnFRQeiKOMD8n19M2qlZORFshGNZFp
2DHTe9OIV9W7Hxd0P/P4KxmW5+GKI6cgvf/TDTqGTVT3mtrqF/47j19vSzSgBNd5
F/p8EHc9IGSHJk0WLikFkh79yNyv0EM3F/zb2HeG3cEC9BZ4dSNGMamEJ7q2Vi8L
03ZFNAk42VCgB+kV8ZEKrIHpQx1xJE6CwFDASmu811FtV0wI/b1PM+MOCeHHnaMu
2gamTceb59TVU/vLge3qtMpZ00x6iRagdbTHv9nK0qkiFQqMyHdisDcHxLWnwEqf
44wBVl15VkEOzG7i7RKHQWgf68/twApiVyTnJrOs7qpxbyBO9nJZNOgESLtLKHlf
ahbVw6bDDiA570kToiF7uIXzsr7hM8YgzwYWJzS/vfmbqOhYlCsHmCFgdUY0GPd0
/DdV4bL9x2na56B5aQuYMxi3aduw+Ycs0XV0zosNkQCfRQqmIoPhPTijcRAMzTyf
KFRt4NyCxyvgNOSUKhdfxJTFGn9Z6sv+oahvClu0kie4Trzl3e6YwrXbqROB3kV8
mfJLfbquAvxnHR7wYW0e/HG1RpjdF7uoUhURvlvh7XGcETYbmEWXVtC0CXS+7Hh7
zTOTCPq4drozoplpX5jNRheZtqwzAnH/qOpazS1TEF6+rNL4V2G+SI5/CCS5VRaL
QUf/nZViETp9/F+w5T1cR0ahQYNtT06gFe40XqARqJvKhMWxxOCMmbNb3vVZZ1GH
1qbFXmHfvVNqBFMGwS0zgL4b26velxZIyRkSIcDpKcK56oNhEsB66n5Num42Qvss
JdUJaDTO7nB8yLwb3+QDjR+szjCR4jG6l//bLfbB4p/MStMrwwNIr9pUTAQqVWC4
m/HkOcVc8xcD60j+7dqGN8OK7kvJklRveUK8kNSuLy/ro8hf4T+H2wIxK457s78n
ooCTkWfS2wygHT3hCg7scGaLM+r8wl+HfRmIgMUUsbqc8biCuY3t+F3Gh+WIm+H0
yuq5Lw/1rMSf2d5eaCpxcuzJotQI4vWS0GpXmJ6XYLm86FyoXwgCT1NFGI3h93AD
FZ3odkozyHq3tCdLf6L1/Mu7H+bHKHChs5/KhMLeRNGmPdt6AgNsdsrQgqSF9DTo
RaHoETfGS0y7y77SpqrIxhmiHD6GOlNH1WX5oTogf5YKWZ/xwJPC56WBNgdT+SJn
8wvCSSMl0NGDvRSzMLXUXbL53ayWUyPIe1jZW5PLI1dCtSqKEMuT743RrtdO62SU
Ky/YYKdTdEMAkz8DqWIFyjSBkD853NDanAAG6apQeOlIYUdsaI1az9urfpf5U5tw
Xgy7qyrExB/R1KrX/HvVnDx8GVpBrV+o4HR3OWS7Fkh/q7gObhBR+8GYFmOSGYMS
5NXizcc1bFmS6pZTYMA55h6hheZFP6A4zfZFrRmJHlKBinfRNIQHi/MItw2fsqM5
rlPxBQUOj9fBkfj25jAE8Wqhgojjkwf0bMaesNTGWtkVoz6VanGJ6Gq4/NT/lODx
fhEyGQN80B65wK+ggmD736wieP78uBG519+pTcPKnj+YQuQzyhyjCtOwpUYMdsG1
TdmGVZxxJTIcDHf7RU6pZ+5n/6hGX2wPkfcEpv0C7C7Ep3B3qDYyMo27Qb4sduWI
U5Q/2vGhfn4Gipb9iaFU9hDY/hHcYw1TQA2kRhLhTYvutMlbMrwOYA8tdKUg3Lqv
lo8MHhW8TFLwzk7K9TgK2KTVv8kT0eq+8RiPr+beeUiz+OMcC4j8rWhzGwr6OEPY
7OPP/OVVLwhZsaz9rrZZjpHb2RvJ+KrpfCOk2P5hb8+Si8JxCvI0MtsS6Oenoh1d
ddGIyusnX4zIxUXAYHrUOi+5eelJZ59PkUuJW6AGwesfp8aEQbNTevDbNUwZgY5l
AlgqbxkeykvgI3KPZ70fGuu3NXR3RyZfFELE5dAkFLRxBWpTs1gOkUL5WLSRuU/P
vjnR/U4bKz7HZ5jKXRT7V2B2av4gLVJ9bI2BBkNuX8PCxsX/GF0XuXaVpUorSrCg
UBMWxeNbspYs3hdHhi1Iqq6V0Tms8TmCj/iV/907WmHbZHHxc0Gd2ADoPONXX7fk
dnlfZDRtlJ2tFgGRaD72nZ4trpxkH8bc7rWwij0FZ2A9CxAgb/VpEAv4zG4PgDDB
SCnKu33gbKTzjyf6LxqC9NW2knIECX6GhKRbpbYMnzsCa90LTwlQN4yT4ffFgN6q
1t20kp6rDSIoRvdVTLQsigdkLhgYnwl81TmONtx29dDMzDxFDhUrRV+Lfw0WXt7H
Lohm9A6yX9/RK35o9inbkvrWaaY9YnKqK3atclzWrpohrIwBDz4XIHmc0PmHGrtv
JWnd8hdSKyc3unV+948XeubSKDZUnulzMaDtXoFdkPtp1NtYDV2IM67wvctQMV1u
oBV7LmM1vQmO4ZARtnHwRKl2kPnQM4sx1jGxzAQJgnYtKIS6vtl7cXI17d0R9b9r
d/M0LyyaYD6tbVPhda8JJrZ8zVUaJYqPcyxq8h8zD5qTVXZ7fdGSuQgHST8loNJ0
XeufKO/ZfpZMwD5clkWCdhJZ9c7PIHBhTBzDr4pO8gKn75AvmEE5WsbAze0ATKlt
QOEZq/2vBDZp00mGCCmlcdRIOfZ54doPirOKKuz1eZOQwP71rLBF0t77wqcZhsJ3
mprsEPnVNkRaf14tmDI/1XJrWFco+GzXy5jaAozteNZeemk/ZOiw+i4Yd2P0mGap
ng+mrhaBhjRsB1R6mOVKUUb0k37Wnci0Q16q5Jh5MLW+LiLeabcyiLngaJwy0cbZ
uQRIgw9klFo4MkWZ1/HYHV4xWASH10kJxy4j3g/QwwCYO197JF/H9uKnWb7h4TAw
hufwBcuXss3ct2JsYkefulzeP+HhKDDt6z9whwN26JWOgeD0zMH1PcydjiAhJnoz
QBgTozrRnF8/vqCQabOPnyli7iE+hrg5QCXYkCB5wy5+qAkh771xhJQmufSroOxs
Ak+cQHje6JguVjX5iCcgZMYDxefkefiEgnmBBskkI4pTHivHKugknUrSCPYJIsbP
wH+Zx5SCwlVIXf1sKk1QtdNxh4lejCj+Eihju0NGbpfQgkF00ga/DDfFLmgDXlua
SN5hi34Et/YmvYWS9nf+SYkgrH92PHo1v6S57Qa8RS7ncRGgVwKlto/nAQ7JGzXV
rV9JI3OT/dxwiQ5pq2t53rqjB2SIiiQlxfxg6zQJBsahK5LIBdlggb8Zt05Vk20I
nx18MKjWKykhdO0srm4G/YACueAF88jgbWHUMPAt/KCO/X0FlV9Chn2M1QRWbbBq
0k/cgRnMqiwmlhcnTE8KGNfSm0PXI0n4MtI3yYSd16DNBWAErAptv8laaePAF1wG
ICus1uj7HxY7fJ+wgLLKZfDTFVnzODv6skVU0nUxjOnw1XaZ4umQKYtvDssbDwtC
zS6c7ua8M4XODKzPleZZ+VElNwGxJt8hmH+g44MvpXFVNfjzMg3n6Bgvt2Y4p/EE
0eotshKOKHfxyxMDva/jzRKY4R9hQSLKqaMBePMUZ0Mjbhp+9c3++8NJjcv2pqQJ
QCwUD0nUdiFtjlAIUXcomzztrwveOlNBBeR8sO5Nmom+vAUMGzmQzavxD21/EFcB
0ocym/MSMebAkQTTS8MMeG8ky2MglGpkKA4vuUCMti/Pxdr0hxRNySDnpSIaOmch
2BfKSS6mrG0tpIh8QJl1XVuPdEssd0QLipdxlaC+ACWxyLEH4AzGJNrOuQq+qlVK
HWRloua6N5w4ua/U0LpsNMIyU/edDkuS5TnlUMRcPVu1KXEUDUzNOmC2Yf40rKQE
4v8A3NHiN2YGsDx4j7vLzPrfifgQ/SNHePSVnog+lBQRjiRG1z7Wk+3+dfTOPTm9
DJQ7j0zbT48nflLqpe/IWA9F4RBF9r3XGYLM8Aly/H9ApUeybDWBgVs2qRPDblOV
ws/iIVn2DgIjKNyIKS3OccmW8flVxoKzUE1mWwcUIahsebqQRTBnGcixVxLscuvh
yizLMRYZ/a5CTWVZwSYNRjQT4TjVwM9F7wd1mVWE1ZHXBv5k4AQ+lXna/gCKLr7M
ZpnL7JNo1HGJotEoK12jfA8Cs7urvgqILHCXT7zkRERA4rgx9rjRG5zLYxBZyCnX
JvpGYIR/cBTPuULV+LE6bksXH4KxK8mbvmfBMFMUZ6VFobRZQMO+e9BBO3i76OKv
nSVUzSpMtf11AwJVbs0+XpGoP4Uk5y4WXrfsNkkvUet48txTAMOo5gLoW2yZ6ro8
krfln14loZkJBnv+lsFAxqo+os6rvayg1IY77SIlAgF/pNzs+dZBJp7gi0wER5W6
3o80NwJbL5/iKePXqNNUMl+NytMli8ATCUfWpSKAlwhAIqWCXwF0IGOnGjN7PYN5
Fz8432+VX0oxPFsFEEF3bXJFIQe26QWAS8ZOi6JVUPoIMvo7JiqurumioTkMaGvT
m3rRui8jYeA74TgE5OOpIOz7onL6t966q22CuBK7KOyLp2HEfALI/IEGXt6jYhOh
7PjpPNeOZvyLWKGa8QsZBZlUyVvW9QWCTT/AFbdFwijUIhFTitBCisKuy/N5cgjG
LJooI1O9UduTx4J9uh+6sjF6W9DegJjC5lWk0y5EGfbAjVyCkW+ZWNpv3Av4yKjx
AgROGPd41R7fv+dPbCdBdwPfhXFf1eRJ1lhOGHKcqFxYvmFo1So9gEFANBpOu5dc
6t/BYGpq0i1Ya2f/UrJNznheHull+aeyD1jSHS35xeJh0uycB/nCurXuDfad9Gy6
5sW2MJvZiTfgki5F39y9QAz6fg7KPL+G8oz6bFfUB0CHCZsQM6607i4Ds7aiTKzW
S0/+hlRT4nYGzY618bj13GJ+MMw4C5A0JF21zN3GfZhsRUz1HUwOolPRVZcWQgV1
dWH7QEgKfymtMvGZNDJPRJ7Ugx0vwaVNseXn8Di92cjRZdY1ukSgDfzqgd4/yTNh
1abtQ8JR8Uil6SzUFQYpmP+QbZ4IaCebyiJveuXLUs4U6qpoPKXjyqFCZfZGnAgA
y9Kg/aSeZonAtdCT6GDkigY+etxLzHVtC+TICSRkfFth3C9f2C/Ie0cN4hWMKFJj
nw86EmC/0WyKDL4P1Ts2GDJS/IgVAmObqckPpApl+2rkgH1BfnPF+qAsVBUJw6kE
9dnjz4e8jbF+Q2jGQZ241m8VgVvMW2/4akALnexiJyVOuG/f/z+h5ndwZXtsSFFo
/8F++4tA89CjxVa7rGn0UoQfAA6uGKp7SWYcDaiZMTQ/8ucOTT1JAZ761mgOzgLR
lOPYDDFrRTi2Ncs30NsRY7Hc7C9utZBJXzsYza4466juK/s07pHMpo9l6Ml7gNUY
Uxk96z1jYvgSkU0vEwDsKXSOFqWkBrAJoTsNL91oIVs3Ay324ezdphgdQU11RYzT
kjduj/X22B1ez6dIKLulAgRb6xh3C+w3RA/XU8EJph2XIU0hpfdz8mzZ8ZQ7mJSA
5DqvdFtzhL8nTBOX1YGriDWA7io9B0m7yIqWz4GFcZtJF/dmoSWk/qstk328qzCc
8XEOJVrCpL1LyxnVv0WKSYGdBP/rWdaxhQhvsIkpKmZ9z1J2Y5FLg9atAh8XTrHl
VJIw/xCljg/h4DEKZ8RZr3X4K+WpXQeiIQT4ctMI1ClVtiEQsrzfQ7OuSpqeMzst
k+nlPHkB4KRbpr1mKo767qhPWpupuRcNilRo2eYiPeBDvmq/pQWbyUml9eUDS1SE
OkmX8AHeXL9nYGMPeN5TMiEQVicaA9S05fIomrTzwbzQVD87jDLnHN3n2d3hJdVP
1+mCKprKZ3QjS+tIOOLNa0ordzuMjnFmDJHxc5NvJDkyURE+XIwGdk2ACqUFDeFd
SogfNiTPZrBrrYtRt6/LA1nugt2tuGtdlZbdbmLiPJzP/QL9MwK4qV0g8vmXRaul
R+RxaEM6UckJsw1r83Fw6UTUd3/ynohKYuTPCAh+w6ArO87W8aT7YRw41VeKsiFr
PUgQofJrNG4QSl8u/QOdrrWrFL/39yvz6SXCpiytabCyvjLU8Vx7YFUkoOGF6+Nj
7jiD3HshC0OQm5q7GEDyOAI5br9o7OYkI6oTHL2sGkT4WSSmuQBoH5s/BhNI5sRx
kuucjWxpw0xzDLPV734/blQwYX7WbIc7pjlTrBOqbJp0La4ZCxgLv2ma76a4Uy9x
SClFq1W7rwy8aCn7tpMi7tP4NrWIlhQ1JwgCV5ALB0quFfp2ydVTEiHl3hYc3VNF
epaBt14BgH3mwiUWvFjReuzWJyX9vDQB0Ks2NTpAmSPelqnkWWntfuzAfC9HD80F
kAOWYR/kBEzNQcNSbd9Y3knOF0a0DYVdeks9dDCPXMneqKIwPrKNLkz3VdkBhlVT
N59+Mw5flgwpC/hnNiyuC12l+aElSXSa1/BafVqEBV29dmBfHg9SAbve5/lx2iRa
9HA7/BdW9ZOMGAFjXRCbwAyiri/QUBHuETIgke17O+ZPnrg/iIVrYRRoEAlOENX9
2TFyh1o+WnlnjnfkP+A4FEDDzzE4MeGpDCSloZocfPCXy0nEE8JE9bgtpfrDHA2Q
9QUYWySn/RWmJIJqe/YPRW/bNBzPrAIOnjKpXyxR2tOB6CKy1Egg1trP52T2ODW1
GkERiHQ3unyjinAUDmmQC0VV5vKPGoyBECh1O3hVWaf7Q138QmTCzxsoAuie9+9/
nrwZMiEhhsPsA9raOagS+JiMwOpEVmimmkN2tKll8MK040wYmb8Mm3IiyWYy0D2R
/4gt1FTKNs4ApJOwNLmaJCnBeZum4tFkh7emqdju0IpwiUZN6FxzP7jJxDKpan9I
VdD99TsjZzNfOQgV3pudRBfCU72hShV6JXP/hZUh32WewSSTynPj93OenitBQr7U
3V6Ltw8G/Fg2uqDpas/oRs0yTKe6kaO3V3OgM9EEe6z1LaS3ltYk6L5ekPuqIfUz
DAK+l6L3XwhcW4x8574UTRDC7igoiGgegN33DWjDe3OZvc/TiorAf7AK9EStSUhp
OoFrhHSDz+g3AvAfR2DW1QVhyT+jA0LNfqsq9djSUiZf9rfRXD65Nw3ks+u4WJTj
EKDUasYkhcOY/otr8YZlE4NGd+aVGQjFBoNjTajthJAW69sglutLKLiX+0jrVx9B
KonF2H55FeG72eGTO5ivlp8ijP+kkeiqGJvY9d1U227Vj5Hpk4TiY3e3k6nbenKT
2uvadZ8DZBWHRR8CItVeDPXdzdH8zg0IepCQ0mTIY809kgOJUs2TwUuN7m+q6GhE
xxSb05Jxb3IBLCsAUajmn5j2TgixGpFFOaPMq/1mbZI90PEF5zfUDy3Zlaiko2et
vX1G1kDemNxFWRq/WHr/72HZPX/ffQTkp9ybcS6mnJ5BuHftx6/FELr9EGSj5Uy7
gKQqWpY7hSuk4BEYBWNNbyA1aO2oa1NDmEHF6Z7Cp6MWQv5yAlJBMHRzYzDH/xhO
9Ooz0v1048lqgIFETYMKL7iOct1E1c2ppAlWSdEeh74kftkMV/vdgFqxaWKcIfse
WEEDWeBjh7U6XZFzXR11On0kMBDI1HEflsA0QlCFt7kTavnK7E9JuxpAaBB+Y2zU
SUmvE8zuP68iUx6vVV16G4L2f64Ofo4C2SiynpfgzOFzNrPYRdUABfrFbn9WU3x5
pKXAlhe+bz0qdkav72ssALv9s6BPt/kObMlMYIK4E3HZI0hwOSulpHJKCKnB6RDT
UJG1hl4jMcySeetngZ45uNOKQQlt/y46GpjDJKj4R3CsZ1S54M5ZGj7yoAd3gaB+
0aIBMHJf/hqvMn5jD1UX/uJwr9NhozK4/AinIUbI+WVQU9rUIoXmbcVBo+uD8FCK
Nar9o+bO0DgHhj/Z2M+5ZOWZYg/6CJML851LfVpmQN+UGkxDCJucDD15DkdZ/mEd
Y6zI8OnGxfBe6EqQtoVSvgtF/EIqDXqg9SuvuowdDRqcGpgMLYMkb73AVBnplPic
VtUr3g56P4mwoP0V/XQiq44HszRCDd5GsEKrNjnLLJzD3/PHNIaPVMMPU2v05ND2
nGGwj62Z/pA/2sKwc8DBFWS8E5IcIZBJqTrOHrvTXYzPFK0RfYUmtp0n0/lSAXm1
I7JPOGETRBKypkpjkxeg+KnhFO7E8iqbqFcXJZdW0nEIpSYEJ0CZB4gD0AsE9FkV
QrtVatt36RyofCSWlLAumx6gxphpxMJlwzXDfn1K2RJSi8vs3qMMs6e4RA4aaJaC
Fjj+ro3HIN/4ezVqXNsGFugfGnUm75t6cLQwkP6ffWFgR97km/PoGrnNNGGn/v3f
SockCIvWqrrFeCy3t4U8PCyCliK2MAFA1qScAIHWcdpY4FSYyP6NIR/h/daKNLjs
40ojMoMAOR1fOQybJB9weKc756KivRBqnJyv7b9bN4odthkxlpv+cSSdOn2u8PB9
hfXU4tILcOBM+ocwjV17/Lq6X5e9KxxZld3+tqoBlY9ICxWW2StivPqoEwNkGa4K
M6QogIGjRFEGySMicKstjqbY7rg8AqtSUqyeIDW5tA6ZO3scnFlRIIgAa9q+R93i
ihdWg5sMChyHcY2JasTNNdF0YLNyiiVx59kxN3Q/6H5vECmsgWPSZm3IVWXQgk3r
E7HAj1MBnldmgUcE+wA0WjHySDISxdDWQiirU41ftxSainhYnBOqFFyQVaLnlzd+
PueTuX0Hcefs8wErOf/ezWvubqT2S+4roRKqBXmaY4oinb0rhP3SPYlPJHaJPqum
kp8jO3YZDKFu+x2nw8ccUoCTEuZcuyL3Oy2v+WNGej2pGFX469AbXYs7ucPwAMPI
XGYgs9Jz9PggjXb72rLaU2fQwHhJsrmCID9GpWEWYcjsCSp3aPeHQvGFY4wLORQj
rchym278q0dtMpxAe7RBdK3umtBHt/oaGJ5TNsrsd9mGJ2EPk09RZ2PT8Kg1InQQ
TvMRNr1kBZ7NfMxJqAr2NeKUAvIt3LIjgYv8aie3/Hp8VYxnRWZ5St7Qe7apUCnZ
U66wWRHXCLwMWsCMeZiWhfWWev1usXZNSqhD5KL1O0ntAHAduULzsrY2izhYsf6r
F1vw8aFvZlscYaW2f0+jMBnU+6sUVipRuwDlfnEcVU41g7U/k69BpLYYFlef9rqZ
nk649wEjmrPapu3lauz+EVbzU/Vf6nkTk4ym3VlQA79JJelE5iSJ4cT0hsytXRZJ
2zVFIP8yZG18154pAtwrxZ8LRt3fLBrrsVNbusBAUijsaubwgnaY+V2hKVgvQ3PU
/bPMKgxnFd2O1AkPtyoIMU+/6rKmBBJH5fkcZ6TfKiXgUAUn0kQwTugRVT6OA4SP
eHAQ7kS35fl66K6OoLtrI+cn1fNERLpHEm0LNmsJZI6Sk3Of4vAazIfhNkBnn6BX
yzMuXzTjf8UUd1Lk3e7osZ9zQUPG/pd+ygefomWCfeUI3Ez9XGINI6C8g87hBylf
Yt2YZ2zOe6WPYLZOObkxB+qgjr2z15JyGdxoKlh/tdoX7fK+8QTj7eBxoLd7eu1E
scIoUM9Q2D/lrmKCILuIxgbUBTEK56pWCLiQmBIQcJN577U0oYbUTptj1o0bLCHl
xc2bfIa07+nQZCMe6eTjmTcwxbvunozfKzxgeN50GVsK+sN9NbugtZOV0SHUVyOR
wIsQq4mvg6DEcHmTCt0esermg+4PJxbbheCIMBrbaq7K3zRmey+vr9TmOxQmE5nj
CRJGMSThuSQ03kefOXcaUVVp2TDVSJxrrNn4HBHJ2yZ37q6z6SLRmrhJVzPqQLuM
YaUMabMki46wlol15WEwSqBBh8bCfxv5mN1wGJa+nK1bkjXuTIeC51g+r6sN4p/n
QrYMvdHQD2gdzo5gHFzmsMTlCK/5+kdjtBPArBsuiGgq78za5d3vvK9iZS1w/vts
c2ZnXfwB0yj+yYbPntUxOunL5nlpGZunkl1M/j399sZF9YWikKokTYsZONaoLDWi
P4p8Mz2176lOGmCE9dT+bc3pT2C+ancKOKPhxBMBN8c4rcb5xYhc3HNM6BQHbeXq
wwQHMAYNFDv70UwDrSDFwrllrrpXK3j4R2TwCqM/XYPp2tmuaVjx+vxn0DAcQKHm
wmsMUurG0yBC2ovCZugfB84nr/h4V5SUevqPM0PG1N68YLmsEzrOHpcj/tcKzC7V
LNd1Po3Dgx1iF7lE5n+bPC6C7vwiQf+HwsIdmTqygY8FyNW8n8E7Vr46/rJ67HSA
Xv1Od71B/3uN9Z32SdtFNW0BSYlzc862OKvLxGK0KZDD9ImwfM0vLuD9S2lRsJRf
Gx8PF9l+5r8F6hQjMsiG61IC5c588dUuitUAGM9mRDa+mnMiXywITA07mTGphvT5
khJfGDGnXOHEYqqO5iVCAYZgTB28jUkQ1Jk/dUaI5ixlpzF3CZMWYWz4TsDQj41M
ZfXph6jANKiI4HWp9BZmnrojXQa0YInNshuXO2Cqp3Vh9vueijjLvot+qE0xNRVm
RO+tJicYWSwVvCxICjTz2EoaWGLPyHLmui0+nG2K6Dm2x9KHCCA0rtRnvFUWUQ5t
9m8PqWISsrZPtghu3HOKSrlP3zn4/lgcmWjHDBhRvAkHkBEJMwsKMW35NUWFyiG6
yjDB7WFNjP56/0Y/XsWkI8bAxwmNE3mC3Qx2mOKk5oj4P9lxknRa+ThVg5kMGj1j
NsucTQDeqPpH7DVAZ1rAyhORwas+jbOI62eVacxcfOiSVgCqGu+3FKBxT5cX+DP0
w39FtpdhSDMVaT6/OrA+deWWj1fDTRCLXNrctizbm7x2tL4o50T9iHWG1MHsij/+
6d5I3w9mA+cGSCFBvIxO8f6srQjXMNz5W1poHE8S+Xoyrr1rflASsoWgAKS+Kr+Q
AtipPyvXEfRVmopIkH4QNfEjPnD5eFM1Gw8HN2NTgwVxuDD+O5oHhJxGUP/5CGXN
RbMzCE5EIDmNWeykiwuvHTqIqBAiJ3XO4UN4ZgqbjBwpPKSmLQ7zZOBUPisIQ91J
QNQt6sI6q993AxN5bVx6hWzsP/SbTwlZPcY0zwEiUTiNHpD20hqF8OGwmnsOyvZV
piXye/nUUi2m8YY02uru4WxwYPo7ib1jwOMORbz2SJP+V/WkLtWu/5Xc1jSi4ajU
gy3TjRmUggUOMZF+cHhQgsBvHyWv6n3JGc3dBoV3ce4P2ICLvUxiF3OBe0CJEaMo
pvgzqsnYl8NGO0SDdLlqnSaANyPjl7mzeyB3hMr0B3zC8hJCHyGkQ0OS2MyYTQiP
HTJu2c0igRK61bxZEMpTZ0firUPbuUcpdJZwERPrVODHjij0WBpQgJwakEfTHrhS
RCVa26q/WrcOk+vekqkEi2nIdL4SiPB1kMD8jPP8R5FoDSYl9IOZUgakVTE0HE6Z
fWobNB0n6z9K5J8qfw1Izivh8tpK9oYYFIHnK+WfAV0cvYxIG5kPPuRjJ2UZL8aC
V02LjB3Rt4iu947HHKer3PbYq07YlYBZGJByVUDyfzJx2upVnSgqueh2yUaDUXnq
0QQA2ypJLXM1/hkvMsrdu6Dt9zkc2Me2m81joTFa7T2oRacGAXYUc+TKcawrGKYs
k138sD/3fexyBpSwyAh5RvBs5zRBZWoRrqg+PN0nuDD8UtnFt2ZX8ioHVaDhxDDk
tVLpTpkmSvjHs9gXHzZ0AKwIrpdL9g3kQTmRSRsIgRWrvDaUacvmQFikBir4nkku
jje93E5Rvo4J19o9YK0EKWoMTutY3Ww5R3NUDozkwLp/KbzQSqUbZiYD6Pxt2M7B
0a3sOvGNG6UUY9k4HNzmuSfP4805TYygT3oPOjtDf3kF442Yj+jf/Kw13uA/xmwk
WQ08UKtSzwb4UFxTPKVpyZp1PxRYeoaeEsFXHhkepF8FKMjjbEu4zeOCGNYUCoxk
k6QJpq/WQCy4A6HRJYkeRDNk2h24xZYPnzzlMgEGT2kVYQ48grwqzHb2hZKKrQNY
RtzcvIv9j7nQPoLrdgDijMNBTlLVBfDjdc9qMVdO2Iv6j5HWNP0YYQfMnhMbxAEN
T2JSe7oJKhVzv8sRhaJ3DM6L9LOFa1fZ7sebEF6pZose2Sjvvq8AJWy3vcDcmnaL
0UkkaxfxHe7nPZFQjbRQHpfAUUPxr9YT6Yjq01jrRCXH2KbZ7jjidvnvfrkUwZB2
68Jv/9EC62ERFyO4bB2xhOwxLg6CTIOWyjAX9bvn1/FSXUOZrNUrwwHRHiIAGkX6
+LziTF2lw0faG/4BEt9zqXCgqbom+8HulaYqLtm+5nAQPOVTRKbym81R5I2xyMWV
s5qMXGtVRrxB56nRY0Uh3k2hyzRynVi+Xp7z+vYD9qW2py/7zHP0NEl1wsSz2QQG
UBPJN98r+fUaet+NJBYyBPHtLuPCqwQ4S33eahPvUHZS/vo9DZMYoH2wk7aBISeX
VKCdRLfq0GZ98K8JaJDtiKSr57A2vMjGrZbcN2E6C2GzEn3UTaDIKupAl2kezrZ1
6XMQgpq/cE50erJkZKZN00KAIbVlXtuMqyMT+D1RESDYVR3b+yUflVaIenlT0TIA
EkRNCkKqCp3LXVJcuEVSihXYB6PQwfXAbEBNiF5QyHiTGt2B2Qp+7FCJoW2kjYlO
0VAUdvf/p2x0JxoU/nDSlX0ucCc1xuY3un6NX2YtqqZPCLQvcpdMVgCVq2iIWR5L
kxnN8RzW1ArxmQI4b3gDsQvky9kW4VvBnzBngOeza6z9DoHy5wW13HRAuJt85CF5
wCgT8Vpo67jv9v4HeclRfFrBBoEKCUe7HqqCWV1cuOm91peZRzFJl+IJVC+/ygcV
MA1C1+i9PAnKMcZO1tz06wAjEXKQaqrSZXTUUv5wYoiK9RG3weHI/PkJ5hJNLKhQ
L/aJOo5RYLTZFk1KpgO1Ba34nVqLp6tQK26T8PnD3fIdIsegnM1xlGribWXeOtWa
JxzjBcp5kvHXrDeXsJMSreOLYTqVuD1in8B3sCxWbY6AUX2B5CiwNBwwXntCl4uV
A+PfwG0DyFN47AnhGoiqg2k5Z4j7c/HkRZLzqPKF75sBQLAlsbnfxoy7Hm0dIlVz
rHN8xToVUe8olBZiHIFWBmQVujC8/XEyrGE/QGz7+kNMkrFbEOXLFLbDAw3gEyjh
HzhzMqvRp9PX8ekQpR/K88kypjEH8nhG3dGoo4MAoOoyzG/VSaTyzwMdjkjdcN3/
GbEZOqS177wsGQ4zBOMIdNlSJ5Bh948A0dX22gg4fa8MfH9hXqi9tyVSTtsR0DAP
xNF94hTO0J84I6T0tSCTzE4Uu734M9RolFvUhkX+jdo5JqFIY/FoGkOeYqn4lHPO
wlV5uEIOFtOxDnRzpkJN3QuquERlKc+dLjx6QWpi+EclXW2LNMg1yZ9Ls/VK2mpg
Ojs4FNjRGfVqwlLkoub34Bn5MfC+AKqma4rE2sbhW8Jckjja5kHcRlhV29cd6fbo
g/erItNOCVMeDDPBSjM86edtp+5lYgOx5AKWzVssxSyG+Ni57uz5YY95qdZL1Bvj
kiYx52SLvimd5e/90l1xhJ0atPpgTEMFAz2Jx70A00JBh2J6EpyKHVZa9QX4Q9y7
3t1oxfhN9mtvB+N6/cX7lJ8QV8sxXH2CKWOYw0pzloXavnX/IqgeaGMtx+DsrIZC
8o70edu2ahiGNLCj4PqvDue0/VVDE3gVgrucYb7zYS6KOgyZIHuZOGKidPAvBYmq
36iv+RZVaEA1cz4iz43fBvBhXDe5CCNUmJ6JDPjJ7LY59dSD1rc8wlH2tIPiX/tl
mMKqQNPfZ5orGpGScQzmCB1jE/LEgVCXdbVxAWD5ikGdqcDw5OfNmr9hfeZNjy8k
t3uFHXlnOIWO+z1rGPaTz26oy8Sp2k+1kZZ79u/RJp0GAsgB18eTkfrU6KJEOo/m
zp/1FwQNKSuY26zdJJg/j3DRqId/xPAl4W/MhOnJKfqaxlp2qlocpBZgO5GPGGan
ebCui9wfZGgWsvSUocUPOG2oR96xQAefffDXQE3UL6j2KKSOWes+lxNaUal6NH6Q
Y0291sVltgzTkuphp+QpecnYaokMiKCK7gZWrIW94/EdnMrZV8oBR7wZS5gkHPSm
B4sLSsFi6qf12CcJfOMZq//LiiUUSXpad8+ObI6gm+fDzp0eez79XotzpWr35PP3
xlJ2sTcE2OdVlYzH88lVMg/YuHRO+SIHO35rAKdRJlHjp0zweQlbGax7NWSLLhDS
0EirjuDjEn17+TNEaQkaXaD4+eTCqaNa11dDroUm7uqqyxFEe9YOWUHnevlMRGGV
kxLk1QYmdM23AoxSatIvYWFsdaQ0+V9krsxPigQdhitpKxky8rfbpguZHFbs6is4
69l98GSTaRfxxQx1xyNQcUYZsj++IeuY1YduYhAjiLFpqWKVGo59kwnUhP1V9jJP
25rNef2AmQro9gRyy3Br9Y2p2uT6oPQkW3i049usMkzADZy3eScuaONm/qPJFtWj
6xsVZcLjfmNFl0p/3EcGPE4rZS8St+OemOSzXUz9B1tKyZnu3HbWp25GaZab8gJv
e+kqGHhA7KrUcn13uOgcTrCvtlcreF8AZmLzoQvRh/ZJ73pQ2TFo85BaT98x4uxJ
Y2xlaDqIqQfuHPzHdned0oNBD8eHMi0irfkG5jjJ5nRVM5/IF4yIZ32XM4y8vwIK
Cs7qZR0mgMW8E0jYH1O5RVnzhLoGOhAyApOEJbgwY4PFIpkckhhjtk8N/e4W7uTa
ZrqSUokw5Tmgdie+oJR5LHvCUaR8PPrNDfK7HgaW8SX96KC8ZQ92F/aU5DWDvobL
wFq2uCKdnF9OnbTrF3fFiBqo34l7aFBVnSEf2G8n2Y1YFzViio8yCzUUf/mNNM/y
TUxRavap/BfLGBSdd3ZF9pV0LPQOMxld//jEbUDbTW6n4t36JEmmT0S14tpNm4qh
A8i5wjGH5XrGnYi2z8FfImJmLaFdlKciV8iWepIpVzCC2W+lN7/oAzSW5gErEXwI
uHEinooDRDiV196Or6D1BienbkZlSCnQ1kM6lP/pDfEWhLNtFnTLOB7cei6VsJ8I
obRBucbbriAQPm/ntmZAVw7b711J6kabmGPM8oJbekhbVseh83YGFgeUV+3ABVZ2
pJhcp4camtABvTtf9hn9GtbDcGyfQQrqsVA4TsutxntoKG2PXxGKzO+ezP4F6wHE
CQEUvg+d915GdIxbCKikx/0bN9mPClPrMhOQyRT0dOLh0nWsc2OhvMVPce/365w9
aOevzaPwF3T31givuocvq8wO1JIiD496cjp+18u+lqLwqNIlb19VBhRHApJZDNs6
3BKwNS1qWyroYL4zjNM6+9kVd/1fxQoh3fX4MtCAL/BRrhnzMCC/xrXVt6R2Z/i1
y0TwRjFENyzzDotZ4tJcbNQYFn8hXjndyua705OkmlDRvXajUttsVq0aukRL50yd
4ZHdIrAf0L9RNDAEXPfNYIbz8jAX8N9y76HEwWOhAVK5Z2+zrGX9gwZBJP+EDLR1
8dKiApm9iEZiiYTNAeWKpEW+FaN1QZRYVt3UfJBtytXXF+YMT2TZCV53ByIP1E2r
ktBBc9S7OarTQW8xAzMslHytCbNyEnJlSgpZ4IR9qQAkqFfi0duB7qvXitX/Y2wA
dJGIsNhBm4WEwJ3UQmtFoQyWRJAVg/8xI/Jz36JfOYBQf1HYJF+AIRiFbFIzHR6o
uB7vrBYgdp1R4hXr8p4IWkcTbIPybu2atGDeukqm4jBzRP+BBJSXkNjFOcjZVaWw
Vre168P4V895fjcjo+rIJzTerO3m7Bs3IG2SrBRzt8IupMMs1u5tRkkfhwp97M8e
H+c0MF+aib0ylOp98NYB5bk8TsnjzkQ+I0bS7bP0FZc/UwFjEyjyqI+gdjXvjM1x
kIQQeuJVTHhIOaGn3Xuox9TYpAfW8Yv/UupJxVDPmqwSgk56sAGyHxEkCGXNLaAS
uX4cYqvyhC5fZZWC3wvrm8+W/6B5Lal2s7IkiDgHgwM5XO/WWGPrT60zb2WVOopk
jNA8F8JMfS1J+Wch7mAc0lS43H/GjRzVwsMWkIvP9BEeTR+2+d3iryQs4dyFlEBW
8BRfvD5yHyGQwYYdOTAHyqLMzZ6BxnmiB/HE6bku5phviYsBd43UVTqyJCxuY9UI
zvrTo60wwbKyaEBWV51SpRZr6BPrtCbD1czbhAl/b07Zrhdbx91WYtdfpUpy8yvh
AeMe3M3KjHbm6Yhrtv415VgMh0qN/pqdVSGRYk1/TDY9sLN85VSbdusXDbqZw2PN
9WYh87r5cniY/8qdxP9uriLS0jud7uU5Fa/WhuQvFAW3Hfed5/+4xyMpMR7wo5Tw
W79cGmX0pxebzVjJbiGFTg619qG0+4ESSUzp1C4xR3D/B3NEdqW1rWt4LdyzosOh
MnGMcKJANTjLzxx4Trgs1VfUwC7gWRAXh2O7OvFQYI1xun3IdkWSpjyT25jtPtnD
DrCu9YIrIiHHt/BrYhpgqATIwMpiMvLvf8lRuxObLm88IvNxOPbHUczlT+1YRBCs
niOX6mrYb0JwH9fcubNwyF29ZPA90d8Ij/Lkg/5szwd+aP40Se1KyfXes7phkIya
15XkgFuUIcC8Jp9XVznS9lzh5qKcP6QdiiDn+8ruNvTZyrFW0mEmxafINj9M02Ow
r1Cz+ku8xHbvYeVKruRy7J+N5YCHY1Nsal9RslFTQZl3Q+gTnthbSSIEh4VYU7JN
JjpybUzzIcwFjQz2oVaVTDaJMQVMc+CRPrTRQADqdL61tNsVVS2GCE1iijL5l99e
5+0cHs+YBHT4WQeuVnvGyCBfjkHIFlqkQeCziI/sv8byJ7ajLQ8wnjJBJYJ4bydK
fsiPKVFCU254xaeMFeSDbp3iJhgiAMJ59aC1YuM9RdJ/a5WzV4NZ0tGLgmv27nZU
FNFWG8fbWMosoJAY2+1BW1mXpnI6p9wQ+s3rvgP2ZT54aVd2mhQxExfldVVL8Gmf
kuHAvKc5prxmnUKu44b5W8KlJgWyzXWI+/OlFtM+4IhWgpkA9ZvAehq5oXKCIdQe
hNBYa5rjXizbwWDrWO3yBrnJGhi/ZZTcDmiO4gqYJ5mYTfmlnYf/RPSonKeVNVtU
ebz3QUYLiRHjUNfE+kRAroX9oEBWAZLBXRJemyQBeHTCgs0BDHi6x1SMvqebUlxW
xRi4sX/3wg7sANwFgB/88a07hnHYZrMF1ZffJIMY8/LCcxnJnQAPoPa5fZwiJG6q
WHmzDP0L4nfg5CW3Mrkss2xXKoOW0yxFc4HALGrxMZ6dW+w2NVMvbPtynQkocmZh
JybgH7WfusXevlKk7KWhGMNCeCiV+gdJ0TWjrIVLY6Xhm+IjAroW0ObwyXaZlMhb
Efhf47t//Sb7bbkytBOtF+wJXXNwlrSIDVzMX73jD/s0OtSBdSGpCI96JgYEOJzg
x03OwM8aILmhyY66XbSQTrQGKc+kINddbNWAyn2fj8LIz4H5+jprj6hJ4iLHKpR2
/PQaH3bWaZLpYfjQPEOoL7J4cCrE2gEzfUjzmfvdzK35iMPv7odVTn36AwPoIISQ
CxZKFLhEL0BM89GmhDF+3arZxQeYUCCxqPWwPf7EGKxYHRN0yXO0DR6oyVzpSbhZ
a4Vr07KN74ZSqaqD3NBRsTq7YubOimoPqjyGp6Fm7oL89P+IYpmL4ecvSFKHgadu
S54zOYHzFQQEQAfg2RjOyL+aqxw5Lwp7gCt2IER5fv3imv3EZrhVO7hmMHPv8TTZ
TUrznNdtZSL8ZVrXHi70ZUWit3u+DZw4PAN1A0Dp/hJsDcGRY6JRauPdsDURSgf0
CY90tAJnov5npzemvIDPV0WRinwRDJo6+OZ1Uqseym/aS0R9QVzWRhZ+tMnSmN0t
PHu48NH1zXqAGmG+E3AbC/naz592n3ExJX7paiTMWTefdq6MVDsR85OQI/OYevLO
k0rfmnIlmiFffCuSaONejwTVkzfeGZBm7ZSUq7+91hJmTzdJm+NqZt1vU73cu0F8
RWNH0iiXPTf+TB97zlLciko5U4XZuoF7ruN4EkQMaltfTw7H7qG8NRZbebecPgYe
WiTtcQ0+UqVoYb0+DJvsAER78R5vLmtG9r9KbUJaB+0hv2J9fIxz2ALjLOijM8gq
o5Nl4vCY3TtvUaI+XPwIFeXC1GfpPWoHNOmI6WoEmc8SKA8Sp8v7YqovnUKAdS1K
uhTIGWlnVpeNle82LUtkvffq1QMM6ZlGNsqZIutVBoqv8M0AihIQMew4qvpJ42sG
vfs+VK/yKRDk4ksP5TFn5kRI1N6HZtrF7TCTqhkloqnbvxmAHhlIt2MO1TNsGBlg
PeFaMfndnmpDrmdD+LGIb5zFxUPXyELrkW8W1MTn6ZnBc3V/lE+QBPb+SgM1oUdc
LY9xu7QLP6v5blD7qZkHV89MzWHEa6CEqE8KdXIJPyA9g4Ku4NBklG26ia7ZSHDf
AC82yWIA51mIM3G0157DXWaukaXvp8Xjt+3DyOMgQdrDLT2eTNzZiWtAKDb/KQk9
rwmWYzNHEep7KtqyqKWDV2jYUFCUQpvV3XpjncdcXvQkDlQVyBIxCyUgK6vPVSKC
k/0zMVK/XjC0nX/tjpOGD8ZzOB5dXK572PEnCq+Y8hL8OyTCMSIXrgAdT4euDhdo
78VvPOmx/yM7ou37vgyRvBUjHQewElDElO2l8fUwwaKT7PyBWCZp97y/26TqfQdR
/FdpSgqdQ0w04vVyF6TkA7+ie5TNrnybHpsgGXX49g3IyKk0nAY5BrVf6LL/M4Lp
+eZywdEoMuD+TleMzx3JAxCLEklYpNWAeYmqfw6agys9dMsNcki4UEHXzZQZfWss
Jv83xaAf3YAPnJ6+o3LuuiQrx9i7FB6CFjmR0BnG30GNX2tyQCFAcCb6TjR+m7O2
Bul4lF8WRvgjTvxcooT3wWIInzQFEQjnPmWvqbyTIZAjdinqMYPmPr9qmOhfvpbl
vIA6xp33ERb4x8MOEdRDJCZZRuF6HYpoX91ERpvBMpwkN/F21QUXj6DQrlIZGjBC
0NB77oGlSTpSz2sPwOdpjlzS5VMqumCjqByaS21cakOwokGvD85F7bq26BP4R6Ww
p/QGr30tscX3O7G1JbbmUzTBR1SMLOE4VR6aNrNwe3KOX7zLEAClqduxYz7ke+z9
lRK6zu9XjNyYEorR8XIMfbgl7MKronBRI/nVsdSqpX2F6Af4E744ZFVrFWL6bJbB
oi+lK96uFncrZU9tbfMbJRbHE8GHiL24Y2v58kdL5+O0fIRaPR3f6jU+Lau5Uj3+
/2g8Ox+hDUMZbMXfgOnW+6gYu9tx1Mc+5yIdwYYbNDkz9P6x2ZkzbJSG7tTsJQ5g
Z4ig54VDtqh5pNyAWTMtA1RbuEteUvby1dZt0E5JR2i59tllhMNVUTGhGSVino6N
zfYVscx8fmVPiVyCOuHCCzWkZ35uET5T6gOAuZ9ohGcpNvPaiPFcYz0VeT4GTkiB
kmQuJ127ZIGvmFDhw2KYQlGu4CDJphG4xJYfHnlFdSdeoP2J9M1Nr8c2YJDIB9RK
dpF9nOFcabsUwVGYfmqQXA3z67tkLC0IYwtiASFrYw+gI2ZC0SHdtb//vodgK1il
6qtoP3vKPTR+bWE6j86nwtTCXkv71EQdf9P1f2GSz1NHlRIvucBPuQmekztxeRrt
GdEoS9wL7yFc1siMk+o53DoJrLwbb0Br/dW8jlH4vrw3drMH4VBktPao8wjgR6LJ
42uXIz+pLIQ65StGEwC5GtKrPk8njsVegetjrl9pPq1/RyCxSt6j4dHh3UbKs3x6
QErdTpVKAV9+RfKMWSKP0B8fwimmfu6gv7GGhoPiDb0g+r5xG0kfiszyfB2zJDfi
Sls+3nIJaO3HwHk1YhTl+sBNZCKA6X88/AUIwwzqRxgnBeq/P7gqplWXmzIMzgOH
5ZjmtjKmlf3B22sW65fIJRppOVWkOZSMJJ3Pfq570OBZZm8TK9poGSFdR4rUOc5J
ua5dIAHYVe1K5IYbZ0Fq5mOZnyqt7DLSyK/xpwwmpMJxSG0241DRK28hW3omJyN/
PkS5358jZjWoKxsx+HsWPoYiYMef43z/JALNPZrNUzIanCvHgUX8hpU6Z0xchZ0p
Khe5EVutnzVfcC2CCmbPZ/l3k84KhqQmSM87Kzhj47s+2FhE3gZypuITl9GKB5bv
Ko/mhrVFUIvq4Y8qthfCL+pPRRGRg8wX3Rns/zs4LzTjYAnBUyt2vtjFL+Z8WhUW
r1enmEAWSILYx8VwCF+bTfXGgdnebLznnSXurB+6WuFPkdKa9XYHfe9iBX1xyMGn
j7yV8Ymq9mhHiCmGVVITEMNc+2JwUFFaf/AOG6pj4N7V54YPHk6HiAdyzniHE0jR
DxaBQtGKlUA9yUCNu55POAEj1Vk01y/J2qkXmY5IlNfQFClyF/aCpRdiPCvUC4Pr
/jApo893+Y7jASDKhpwfcOf6LFp0c/NvVM40EzVOdCaOPHnDqB3gj0tzdWp4uy0e
g7YH9iadrqCBYb1+F50wIaXy5eBRJZBwN1NgrHOY8NywCDV7C6QwzJp1DQw3KAwp
qxTB7OAwaiCd8Fv4bri3czqoJNZOJbKHWBUa8qne0ALHDHjozqRBllytBOGpjZcr
F4W4iECXq8W57Ru7Ti9G2ERm1OQrgvJhFeRkLSwHu8YtHKplqlEIW8CDMULTQy95
N4REwG12+h8u7AUjDfKqjZK8ky5gS7vab9ZQ4T3hDvF291p6XSnExZT+zxFtjitt
4srbrjPxR7LoLr5iWdGJMuUiPR49zgYaXxzElG4/fzQB1keEGstevVj1jURgHnMp
RfD5Uiq6O/+dRwUUbRm62rundsVwOEsv7SuX2OERtulT7sKZUVw41iu8ZEEufSd9
Y55VczBGL/tJq0EzdJGEYAaYwXAKvtMhDjoF77cabUVcwje/MY552YNw7sF7rkWN
HxuEsfO/ulIsqfCbmj+LWcR2KPbMEcoSo9UCGA/54lNYFjOunxXrEu1MRvRCaKBO
GaLriJGIlV9b4NLBm1VRhAt2LIDlCRvUsxebkWX5Nka3wenZQZ3TsoD7KBORjVbB
fUfGkHf+4CGFxe6o8+W+L/I1v8abLEi91RqI6NmKysQVfrt1Y29wrwbCw/dmjAgW
Jao2BF0otY3wd/9Z0W/qjBABH2pk/8cCPDOWzE/xZzKwCNJYRSrhZ5+NmqxUquOH
kZrXJmspMA594FWXKru22NKXScAmxgSciWlP/BzHpUH7Nxg9tY43E43lm6UZQlwk
w/v0U1SRxuePyDLgBK3xpWNEYvfHcKCEb2lzWzSFeRIGbP2QMvTZp/rGyExC6BQw
jR3fS2ltMQdeZ90BR7NrG+KTkzP+5yKEhzZ4wqsgIlxeHZpY3CIpa/K2S6qYWA6Q
r/9pBShLq0DCIH0oITe3Bx3+SLJepvf/rZVu3sH85Dx4VvCFjfKH1aQdca5sDUDd
P2JGjO/1luukdvqoKblnQr1Sz5cqFO7DF3sadrjzfcrqBWU+KX6fYtgiyFmjGvNb
5ApO+uYX5IPpHEYz7A9x9ghz9BXcgeWjyQzdz9OI7rPo7+U046MGdW6udt7wApvo
u7Oau1o88j+/O1t3TtFOPPmgiOQB9qS/1uGOMEP3kdMm8AEJFt0Cl+Llp6+7EjQw
vnw/UAFlPV1i0hes4+q92YIe3/C+q1vRWBppoyaEWArVTzn2KgeuI9JdACn17x67
wKerMUDpfFmQv70UYRsVqLIosGTz8HrX8YYuEmAnwHxnXxNpPTaQbSwpRcmQsJUs
1mo9t01Nwc1RzTEAM8woUeuQjVG0K0SbJw3BmTY6wkFrXuytSbmQ2wT2FpIaX4MU
CFafFacob7YSVrRPKlv/3TGAV2+mxPFxk6HonvAGlWRriCiY6fx0Ie3n/X6HzgrP
/NRXAc3+XlmB0wuoYTjpeWwvsK1nXXe6FBDoSkhf1rgzCwx/V0/YWCBWz9M8NQnh
3EMYMSP3ZIMz+rNPkjVFi7NH4h7ATHF3p7ZCiC6LDfAgcrzktP2llaVsH17kyDPi
D2EkQAdaqFw8YFw9aWw8swBwu8TC/S07yWh36mMdmA89O+tstf7s+H7NYoN/JPm/
7ecAfsLIXNxrv4GjAdVPIC5ssPDaNnNUvFecbf8t/wSIO1pKfzMCv0L1edVAWbsL
VLHwFx8s3+ipGQMjcm8n4W6c15YX58AmuhSOhySmOgrh5vtbY5QZvR/Hn9TnLrFA
Du0bjQeasCEr2h7WfcnuzEtKi8Jjb0DkXrTyvJ0E0ihqJUcsjbrlRgdhBEVJargo
4Rlvi/LuSa1CsNWqZtVZdQ+iJjmVG7YqvwX1a4j/paoj+pFhFlGK0IUDmebevS3T
vo5i9G2TJVf5rACVYwcdkSUZabSR5J3bG5EE/fcmup3CBBcWX4C3LgcUBeBJHw3O
nU9vMXF5em/0Dj53xfR0pbrkWSJf70UHkiqW/kU6C+WxoqMaRoF5vmmoWDnSfjWY
bceU9TOWlNVSITVlxDjO4JUS+AtQk0UTLFbJ7jQOICZjHZLtRSt5o3FJhZo23cYM
dk2oOmWkqH9BNrq1WyJ1DSIE16tW+BXBEwGzF/LbdFPfqMUKhj12JgGCKf1C4vxN
tR1+/qBIV/WpZDl1qL3jASgYp018ZGM2thWTD8kY99HagkkwossRVY8eYmE7kI4b
zn1dp3mxCfHjt621JQpd6Yqn6FYYizWlLKQ0igcKAwBD2X3ReLBl32daA7wJXQB0
bMUhCOtyKoCZ6YWsV3vQt/0LkGvP9HfP8QGCFMJlw8zuLBcVUt7Qa/o20mGvzKsV
anfDD3n61T6dqL9tOJLqNViqeB1S8Ldlt2md4tthGLHaeQIXYq19EIV01OJzZv0u
2+g11wRoH9ARAorTd3eGld2dCuw9QmR47WgGACpKmPOD1JeBjW+btgGXABhaXH8S
lpGlDRCHfRlZIJqZ2ZtB65UZJFNyb1gWCCuxv6NsIlNb+7/AuHKI6xvux+6cu6Yo
2IXQYypWzdJzsVQ0ArP1zcLM+DX32yza7POJ/4upGr+pSTki5zHn/qg7zFHI+1RU
Z2kXrqklIgXFRM0noSx3ucz/N0X6VA+B5PPov8mnkzmnA3fBgleNME9LITfOFKbU
KWQv+DMRs3Qh8wYc9lQSZs8ZabBBHSkKmQr/QWV/HyugRs3ZPm1U5z72BRskcar5
b5pxcC6k349mgSjGWLsTlKFFD1xDVtlaBjEiARgIz8jPxnIPNeJGdE98KJcSzeyk
jZn49QEf9fE+oKbneFObRuzMRg0YyZX9S3/VrXtjSu2W2l7hNq32G/jgcta/Oqsd
EPLw7lUbEoTKSoida/0EgwlMJMJPve+k8mhs+xARSPplesaGCcUDmL5RQmhE9dvg
MsPmX8hr19HaoGSSYkiDG6f4l6Fg8g0Yy4342XmpuUXblPZnbAqr2rqSVYG/E5fK
K4f1waQWWWSX68fnTPR8E1Snx/77Ii2A8tDQHrWN+/uF3Q6FsO28ueB0m2GA8b8f
EJua41PmUA/9EO7ScD7eBMVOiKXJhnXPDFAJPf2tMgXoVWaLFJl2CJQB23vuT02P
7qao+vae0cv+je26NtHyQdMYsA6+pQqOxKjcqDRDeg9dMgdNF+BqUOdfe96T1hHS
8qKwnhILZQm77Du7yIdy+vwaQ1OnM4A7+PWRjZV8B23o1U6Rz1/inZ7zR1oSccFO
R6b9OC/NlFEx4wEWRsO6umI9uOprDu33hhilv97gQoCKGDCkpHWV5OG9CwU0Flma
f8TXAk4x5KirMNb0rx/PczDfpvR7Kaeq3gBE+uYRYoVUDgLtPSzGX2UEDtAzeWDX
DqhrnURd9uREn9z6GL8LMhjYUPRJuJawlGHfvnp/s8/ZSzuQxMBWYPidKnYQPV/g
OGeUjRHPV+knwjsou/zP5ouDgTB3x3N5Ueys9nqW2dvm1Fay3FM72Ww/Tjd4WfEg
mVeeNeuj6l30t+mVXgppyDxqPYIH/HYQ5GlPy/BDb77e5uF7hPg+PyKmuyGjoBWS
Bn4/gyDv2Qo1gkD4WIJFj0uWDfswfcrVbehKHZW0LlUTB3c7N8kr8BgVC9MiZe3N
Kdj0cWTATB2LJjn0/0IFnSrpuY2GWN3TIQmgGYS1YbnWVKW9ApJa9/XGXrKqiiR2
zanEXVZXNUxm49iHjn5oKBOW+mev3nMRIE9dJQ+vyIJhuyOv6L0MIs/EvxCl4U5D
HluU36ponVc3Ukldfe2WWcqndzT2LwdGFbjGdPsCy1B30QSQl6zat8MmpTQyHMJf
8MS75Cze/iLeIZINJc/tm5pcAw+xSUVtVSkhSDSsnPMykP9bGDFcjx/09DxwxERD
7Vx08GlvEK54oJFX270HC7GEnOOBOgfm7YAgdQUmrSgGEnLoZ9jaaSCKUJLoK4xy
E4/hGoSPNKHsOHcqG4RJeeRQ5BK1KreDJMaMOfdsrtuRvp9piNqvGBIKy3eYOA/1
iMnX1j0UPmt64ZfshOgHd/1r9OvlFhH+rfT4sAzQwL+9oE41604a4m0WSz4CB46S
eSjjAKXK5Vv22IEBOyNYhdl0PaxTjj2l1yFAu80M/Q7MRGZ70cuofsju4Eu7fGVE
4Z3/URyysJ1O+tWRFozfzSjP+2lI+xxvjJqShFHeLkmF6451m63dDX4ePF30SwNc
+nXyK1lwIMBX0pKGamj0CGBWkOn9WdTHy7Xj7H355JqYnmRcKyjaNQpC59SYw6+C
DYx5AK90kezMQnZEFwTB4EHuIddlU9YqyVondtnqeiQrBF/9EhXX37ow6gQidFAu
ftZtBkgWbNLrrWF/G2xuwvfY8x3vFBiVXL/jU6eibWKuy2E8hrlNftcirKoz294x
lvmVM6C0t3NNvl3oHMZcmuTuIeGlJeiSV3Usvi7cWfS+RkcFYqW6XDPM2T7Yibzh
YeiIcuZTHADyzcmTq7BLU/CGYCLqxnCJphtEClcBnGTrFQ4QVHw/FyEv/+A3YsHi
Cam25kRZ59uctwSeYIybxgcOsmQBgPd3Uep8eSA8gYQSGd4djlyuT/lMJubL5Ewc
fuXm6sHtBYFsRxXIbmqQTM7Ak2NrDkPUaY84OlrKSAurkPE1/1AGRiFdw1kiz3nD
wsncUQVDkgXAN43EYUO5nwtvD4+WZ3/bGFBNgg6YXb600f9WACQbm3jIW3dRdq5D
KI+uRxZ3ujX3pLv4sCHBIqp/UGB2YaCyQI3mRcceJIabCALc9mLsWaNkKsqVUa7y
MG4OKjRSXpjI2GDgjiCiaRi4onSWuVN6aLFkcymBWImZ3g/+s4P0isGhUr0Rf1VH
hWSy88aTCC2rK7pwyAAjx3ZAtYDrFQguMr3cRSvtEjeAFRET7PC8cJwWNizMTC+N
h/14NtXBoDFgq/Wxa0BQgo5Gci4bPqmRFLMMWNbYpvDDLHJSRoROFtChshgRdQdp
rEARdfa/eLYVfBlmrmSV/MVHzMnJEiDvShFKD+9T838xntOlTS0IlZnB21sS57eu
k7oT+kdMUXckQDzGjjmzTuliXUn3ArOhC4IPgSq6n2uoWlZ2EgsvXFKEhztEmzAj
wQDZf6m/yMsOp82p2AMFhSxMxrSLujQjkcLI6sR66CD33w7nkxn8Pp7rxYYJAG2y
vEzDBOfGS5H2WIrPYhaLRxvshNogSGQ2EyMBCv2SnuswNRaD2QiNxyraiSicXuLW
WO4p0LOEzQC3aQBSDFxP5usbkzX3/76ehhBdGpVfYxlxt+QTpSwEEQ2xM2fGcKVW
kZZ+KcEzcHTVBNkgsa6RWDMj4vo23rSlSyNgz46QKXphTTz0a4vHZ0x8xM/N2A+3
Jvttn+j52C1T4JHVa7Rw+gl7TJOMOr62ZY71pGZVaGZeagUKvU5jgxODCYH4rCYf
tXvpyLYPWswyqpLR09HOOJMlECyMlOKIBdrGQK6KwiUkSkjFogQ2WzDLzA3UevhP
7EKnqVp4pnOXFLKSn7gVwOpLH+FVcJQEno5m++ow+OXzghukKxmDQFSQcZHFzfzy
WqNWnWEQgoquQQVBE3F2ht9Aeg0f4ip+Zbl49IztndpZQ96fu2EFaKmIpzXQ0Zwp
AwWCVXgrooS05oevRjqB9gSxK31AW4ngDwNmtdNaNYOykYioBlzruPVXb7mK+rBH
kHeOmdlh2jgtMYKTfAEulKDG0gdFS+Gln60TlY9dzZtxjtbYlOlGbpnY71MmKagI
pzfzWYiwDC9DC3t6cZlol8dKJ+5/NY85S+vxbHTf/E5+QFONLaKZ/k68sUq+nm0B
C3s554hoVAW5/nNHb0Kg6ROphr6csZtLriJ/8O771hb3vFsUb8b1qBTffjWMj40I
akC4cNByT0NpG1ePWTx9+ADqwMeUo5lnffXIekn/0KVayj241bdTGKUoC9uC5ltc
Xi5aS8YtM9GAaPHXaG3txxYjaJ8BZpxVu647HOwwaMNw71L5BHMNpH3J4oVyZNcS
u/FjYN8ctn4WCNJxfil8xIKfGde/txouvvStUNRk18OR+inaENB+LsUq6SnH9m8C
tTktZugnROBJOFcXOeCSDvs3tZ7eViEzngisdwcoiokCpFZCi0KOs8vKkW2RS6NU
pmDDq6hJF1XQsj8+/JFZJ2yCzsO12gmfbEEhkVAb8WOuwB1L9pqp+9DWJfYFfoLe
VwZrKnlvw8aDa8gDA8QP4ldrE7N6RLeaiAVGRNb5n5NsG6OXEarTihasaBuRT8RQ
ZWwV54Jmf0SGevhvRX4x6UhbOsRUaDvDPD/TwkQzJlHR5tVUlx9PyXTHI/n/mW4h
AiBL2xhmAcn7OtmrtE84Y5L90+VA0ZO7WAIdrBSCl+ojA/fn+nRJbOJrMBPLXGJf
v1EXjfflApcVjngjj0fcWOpElUfKFlDQ06a3cg9Q9861+Yu7VD1TQ6Z3xn8Vq2Gs
SOa6X8BkoEHffXFBlbdc+yy5aIWlT2b8/5BIbe2FW6ZXgpDUpJ8/N+0k7F9sJCw+
1piEPJ4aQaUbT8VuU+pEGmmRFvZ6w1SsEQoeOT8tfrL5Tf4HoD7EY0rBH/VyIy5l
517fh9ORiO1+deYJbNyBJlIS0Zj1FrnVhiId9C14fJCC1qrA30oO9thv05Sg4TrX
FwimrKuW6SZZQrzob591C28CM8Cue1BTmyKLd9XgOTlsROH4fqvPoEUYMwLeomFV
fQ8FYD/sFb+D0kbwUoqXnFhkpmYn6OnpoBewWLEuwFMk0J7ARaG16ecR2C/br1ny
J/4VeWjTjYjWkZMVTFnrjQf6EN3zUcm44kvwql9rRm4Q7+ba3oN/3cldV525pA9L
3cRTWI9HrN7ezIecZ8hD0i9ZIcTES44F8BmY1Mqia8i9wgElNOHIuZ1a5W1Lx6/2
QRX+VqrH+Hznm6kUb5RPzvBEOX8PfDCH/rJYXGK+bPg7T+ZfSbBUl4vrg/YikwWs
6PO64DPCoxrk9/bNJ/28QABVPmjQX4Jcj+rH9uSOvqk/N6JdJBYsP72MfXBgZdWF
JIFscWHKQPVQXtkjoIrqQnHFscar4Q1RR6m+nVoL8dDFV5uIUmkpBKP3KGtjKGoC
cBelp6QYIAraF98Ds8YB38gPElB7HJL6lwLF9vTAphPt/OdKf5yWH5WMCkC2iDmL
YSTCAQ3EOUUs39IRixp/h+YbtU5iZ+oNhoVWjX+AaN6FVQAnIHCbTEC36/BkZTFt
e1VF4HnAySHtK8anbUx/7/9D0rYDAI5E6CShTQ7TOOXMEpar+CSO24o4T6UHs9VB
XoMtqCwDb5RumE4tFUP/wt88QokQeaptJnn/72G2vz0+9DO72Ztmb12U2FCspquM
Ap4LXomrJHoc3JgoP65cJu+q0dmTMdgg4ENYlThZgSbA4vxIOKJog8rplYbWB7Ub
4jMJWVcKhRmg2FozRWVfKc6lZhleWJMBkn/ZAvBL9zjAVRYx+IrinQ2ev/duxeii
UTvSwxt5vLYFkMI46Ix360f0XmvsVM97esbHX4vzxZtxZ0YBZOjpSTwSgvq2oWwx
B1uVHbkhMQ3vJ7sjcYPpWDJDxEbRrlrlj2uSj5ILc//5JL4j9bcEc4bP442Zq0uK
flQ7N0/zchSWRZYjr8strit3CxblYRmq/0go2Qz+Wy8+lWcayO6FjGaD1jcvaq9h
nLLSpJivp8WnSzJWavVoys4Q3ePEIzpDwsFdbU3l4XHzfMMLAigai1GuHp3vQNh7
3wJImLfppy9ZBKEw+F7+qExdZIv+Q1eQdD2FSydCsr2BTqYlpTEkWei3qj4/Fedj
rh3ZdX2GDfZYF/kp73W9pypm34yd6yaZmxCx0Q9whFArU30iJsi0Yp6+V0viDGnK
3cLPClhF+swKHwAvlw8yueljLh3ZMBvlUb3+KvasdxPSwWanAi9L9sypQhHI/Kml
ybwFm5dYbK34dRMNrNMdpjaCAWQKDKzOvDxX5/0sI+DXeIBmFsr6nl5ZdwyMBwbl
ea4ritQXCCRPvMG7YFh0OuVRTW8dZKPczWYKCvwmyo7y6m0ZPIkm5zasRdZX5oS8
E2/OE1SaPtBfNoiq7JQrsUU4nuPyqJDNGnjho9ox8NajdBfuzWGlZ/g6JjFrTDzD
KT8ytz9x/nLMVjj7clUQOq24oiNFVmgAplY+TR6qsemfzuwC4q/GWxEbqpmxJRtQ
PFjvCLpwQSMxAKPnO1uhPKdeuUUzSrYnA9OeOZwx65qGJ7wjKTeZg7OUm2FI4CSn
3M5S7937+zrtkO1LqlNiWSP4IhK5zgWKVcXeFoRjMRZq4ohoAAnmwLX9O5IzI2By
0r0z9vJNRcLkW7EDX5LGoCgrKfGG+HhKykIm5SAktnONdpwCphSqtJt3f+GvAsY7
S34qRfKCc+Kh+IR92qCdPyjS01kAVpUlzrI4+XyKsnUr1eCajjnneqJDl0Z6bgLP
iKWjKg/dhKj+0etjAaunqz/blYjunhZOs56tdEEQh3u6ubkFv4CTDjK0IULA7fpF
tbr1q7BiisR6i8etUtMrcIuvGT8m72b6JBigxjATTOVM4WCstjVz3CxaMHnOpB0X
3qdODB+nYm9c76KQjITIhU213gqIkHP2U3F1F5OU62Ze8YZ3Uw9B6ItgKWeQhb99
8GH4FzjWK/3fcgjvhQUWO28VOzBmKNNFZ9n7YUwj5T4rg3s55b3HQ15wgi1oIMxl
qFjg3DSjm/VJJ0uZ07CYlmEcKpFhzP3RuEEXLyudJwqoPvoJssSWcN1qHJqdZNen
8bmb3W3yApJsXDmR9jWbd/Jjwo6Yh53+BY9tJWqBmxX4yXQsYh45jNtiganXaM8d
G23EODJ+6ifc74JuBWZ8lILxUVk54B5fRhwt/YA16nVAFgGo1loqDl0GaGxKQhB1
zwopPn46jV+ic4bWbuMjQlCkqL6H6w9uHCC6KgHKLgbAt06XoV+43GjYDVRAgaAA
Rs8mPCvm+AIFL2bnWSiGZ3lW7FVoKISGtzax25px0Kwvlgin2HMSd/Snh6nB5sP3
O4NgwFEJxAc9sawH7K8T5tEiC7HYIaxn5hoki8huI+BmSnCQh9Ilei7xS7Ns+HQh
ZO/KpxpEUqznnAF/tNZmbVik3c+PwN/f7vplLWcOMKAfaDT9DtdRIcukJUoSyRAC
fw/uQflCawC6yD4pOlXQcUBjhKsTEaTGZgASz/N4jCRHWjhMDGh/qcrrc/6k4ucr
PhTbhgDeUTj0zyRzC3zB3VG8bpumPLB3s1lTVJA40feAQ6ryPgvWevs/IYRExBJ0
Qyg1HeCRvBtMEEpoKjLWlCfxrmcKlvK4dd2Hs99zbS4LlSLMO6+qE33RREJLVyfM
QMVV0gu8BG2AMy33kjrYg6TrPAl32pfTtHYslxG3vIFshl79UuHUGdIKzdccMiyZ
qCisgxcoq8JJYYvqM+/xKhqoIDIlrY0Qkc4ALEd6+cAr+ViMK/v6DuuEuk0Y2zXX
uijF8b1ywakh3u+GCTJ/rqbCCCeY9G0fBIFnUu8Kay8pIXzqtOAKV7v+ym5qGre6
i4x+p+0Kj9okV0eQR6soFv9jSHXBoWAXYELwNVCCMUk6ACYshFmYwAavcp+xgiZI
bQa+iZkkLrB28Zg1CG+17hEI1s1ScwrEZJ1/pkWyPd9ZNc61b8t+dorXZAKkucs5
VtvE6LxCg1DgAA+d9URH+1BOPPWiwF2ndxXRItLBFUQ1XMp1Zx5D/X6/LwhvT61T
4L7Tim3H0+9F+jw6U2MLwiErUFALc9I5C8dvJ7irBvNkwJ8QLV+Nw0uGw1DuYxem
bd8086Cvkzcb7LiETmmfzE/HQ9nzxAU7glkw4VSPRw21Q8r3XWSxyIURd2ArnCho
LyZPhXGBamI/vAtuzvIdVNqVVd96EaJY96Tlzlc5wRn+cEttaol8u4mkLV9wooxs
+zQkM8aEd3kYO6f3Wj+4a3LMZQxYlJCxgaG5QpX0hEkRVjB2B3pnLLov3Fy1Esga
ySzKK4ZdDcJ7RjUEDkrNRyU8/76rOO9tP8HdPyLXsdUh+4r0uC/SybNinF1nD8xC
Jlj7BQL44zTsgNGdACEn+6ASCeYk6T6z/suLxgcl+xox+unPMMX4ENVg7bqktITK
6Ul2sDMwhbnGBTcfd2r2rTplpBHdo1vvNJHSQ6K7YG7ePb3gsrNOhUEjBp6osbJ7
0gFBc5loBietZwmLr1QrIV/cOdZlvOHV3u3Tw2Vc0tehnXhMQtArKk9pJTb1SnFL
c2E/hRUFfh+ykqe4kddcrY6uWbMbHqcIKldhkbDlRjcu1MtAkrgfY9nFXsaPVp74
V/UmYLwOgB8aULhIWU7eNPqVPpU+5PwC4OSY2bW9kkdBUykeEIZYa2jO3PzbL2DW
lqMB0Ls5Z4d53H6MsmW/3Cm34o8y5azGlXcclZoLXMbBikNyZ82iKeM7off2PZyj
1WxpEKIb0+WYHGTVi+bNZE9q28d/TRZZhPGi6bOcXxa0/j5xJj0Qx0B5OmPgm+3G
/w6/tam/eOqBWG5a5g47OjqUuTJKL5JYVCpPaevlgiukGdHNXzewVE/uZWe5n7aN
qPOoCnRMEU28Bvq2SpKiraD9Rg3FgsCDnSjwUecRwlogcJcnBTZ+q/VFv49Vrqet
nq4/XvFmmCMwhCvYtrwUUz1pTkDEXTJZThh1vcD50EZICj45Z7dAPMMt961gne2I
lFrKlcGCyiIy/DI1FOXJDY+seZjzWIAQeEvve5e8CZOMZvoidFoDuAifva3GiEvC
erVz8z0mCfy9jgRfIku/Dyc2S+YsiejjjrV8RsW9/wmFoYwaUZ2JZKNFUwz2xKo9
YOYqDAfxmQug1Zi/ahnzojv5Il3/OdJ7Xw+Uf5bhNGr1Xr7fjQZfOR9Q7AbIXgeu
aO+3e+fdkDIwX5acYcY1QUPYdXABeYJ1jJ55mDaE8mZKjAn48ltlZzb4mNgrUkcR
QFCKUcg1KGqKT3afqT1tzEqVxir0YTuCHu3zfvgaGZUlGFnEOOmQc8s9pnkH7N0k
Ip4BHHRSi+7zNmI+YJBGPOevA4dR7UzGqCmTRPPCFQcWC2B7Sz6TjZFK4EZ4YUKb
5cLZuww/kJ1qgdJls5L2pWNLNygQr7OrY6ucf7ah9ugYkP1n9aPhGLeLM2XwdZxv
FGAEdDeXiJm6g11f+FaLt4dRKbn/zniFTm4lGxXaFv4rdwuSLy6ljBnG2d1iFKiS
OLa7j1y6+eNJaw1d0PAHGDsODAQyhRpYJkKKNid6+cne3zFn//9Vfcjm7xgtH0q3
Yf4hZW3Z5XaEbqgMursQOElHpVyZrWUSbyP0s09rgJXEJycUp6CKOQnRw91VXdCd
TVHIbrU2CZRG5ITsTpwYhOKbmFLkJnu4ct3QbQOfCyYfOOc1ARqNgj4shV4Fcm0b
2/2MhGYPfX/fHXTq+5x8gq7dfU+VMY90dQkMj1JW/HoE9LtkCTIq86l+Dpn/KOMP
8U98Xd1JMBtdEzItW5Y/EofWQ7/dd8Z4vyssouWJ0n4YKnhv+SXXXBpPeh7w0IrP
SWUuIT4vo5vdj5W+1Rqr+9S1M5QtJ9sCPgMz3jwh7Ttxl0kEkb2cVowFL6EIGS8i
WWkeieu8TvJ+vWsNFhgIwBkuiO97UTsAEUu3SVAwIvIpiLVJOsJ4+ryBjpKvyOQY
j+2E4wSyfYB7/HJh+2smu+cGNIFnHRQIgG/8KCmqVHkdDC1SRENxst/ngeB0HiU1
SD8Oz0baURgVByE383EvcKEA01q9UQwGbD6vLlU2QMX/n5lWzajukQ+F1oxPE6Vb
T1CtMGgoqPr7oPt/OYy6jd44pAsMM4G7QzY2xAL2VAAlnx8rRR7rTDpz8mMGEsVL
WiTe7Duxt2+4P5RkM3JTg8EyuC6GDOARstGge4TlRqMWUbMmPjOWHzCosbbppvY/
o2pUv6rd9A/XMf15l4hbc9G8t6e4g124dtDuOg/BJlddwJl/jCW7Ahn1l+OSGWBv
yB+pDuOiHYjbcbKpk0abGxzpdML7GdBsHukfrttODctef8q8m1pj5Ezy+OmTh/bV
lRWvb1Iifxw389no94VyiikdZ+OOcTXN1Dg46IuVglEGGkrF+qWgrNuSrVUrtKHP
tGoru+VOkYCoqz5Lf2m+QlE5JYZ4HKPntJB0/lsGvkSK1vWGUOmvg236i4y4i0k0
JM9Jg4XXEz58whQ7MVOoU8fIBWLsDmSECRvQ3yYDwlzkF25rMgPh9zoFU0qMzQWW
4qIIdvyeNqTzuj7EVEXUlEOL8LlfWjOoopD+DtiqAliGgqv0Oiu3z782Q9VV+ooO
c+br0uTvT9yDlBEdKtxxGh9lYVisbZcyDHtzcxPWQkPOeXzKTclOudFx6N3xrNOd
X+2oAG2EdaRTuGd5QLM+hi55QaTn/dbO7FIYCAGZMMHBD1T7lsKeGuVnLO161Kmt
M91wW2ZyH/sZG+EAHmxbfk/aSDq6D3RishsnZcf+dL3us2/T+WbbTHilwK14EmWv
h6EbXUHIIs1GMRLm5gFqcmb7vHrXzZMj9mvuzWIIBXQxYvPS4lElhlvqUNzFe4OH
QLxst329KtaHgC4PbhylpE1Yacu4H7CDJx8PjoJ1GKuRZ4FIu1ihn5oGpPBtoA+V
PLHkzAsd5m+SR/zlQZuoQTy5ggA21NWa6VAr+a/OHXzxK1op8cESX49AYN4sLt5M
so8ijZq0+0FOPY1TQvf01OSG45NTUOfmu7yYbXO8c2P9sbViKUdzSIPYFCPv2LJ3
i5DizTUAmwWbs621/2fv9l9kPvj42qpHHahqv0K3VaqucIdWBYFxsMHVWv7WLBv7
FoAhM1jGwrFi6DdjdZ4TSNeAhShmkkZQWiVEN1wCbKIQvZM5WkiKOGRrY1XR8xqn
iv+91wytYl29jL8PFnM1IjJb5ZRvoOD1txVcNlZvrnF/fasxxuR+ZZagvAInOw+F
K0igYBAL0q8x3r2XJz8MnNoah9t/6u19/w3HiJv0rOt0vg2w2b1c3g+g1H5y6Ab2
AvlKdXtZicjcCNPgPHybs2yZ+qpu7aj952LxB+HUJ+3GhoP88F6cT2KLV7OCGipY
jDDvWVK2LxZZW4/YsoiPoVpx73aPpzFA/aOC/ca43qpFEVmr+PXEk+5uSxis8rvt
ZDJzeKPvC0gCw7HY6z4o6aFXqGNwtjmEhlv8U5xLgbZjTG9PaBBh5Vn8+6DmmRAL
9eLiYMx3+DO/XdRVN7n9sJ1AdK3P/53+hlfXfgxVO9WG1nCA1eiEi9WSS9tOiMpT
7ct/ywgpmT/wA2hEw5oZ7KaDe0THlAMysuxil+LfgkXyqSzOYLod0xjmdCYXWH0Q
d8G26Kph58PLbjeP6mOahYHZtlFv0DiCMKFQXgCz7kwSsB1pCBajxBoRGd09drEa
lCPN9uG4flYY2xW8sS1YvmyVKVxb98JzYbwm0hzIB7KL7SU6N/caZJUyD+zihZDy
U+3j2IEk1VerctOVhG6meryXWoScWOLxC0w6t/GyDNX+ioO/lwXDmUdlkaxBHOo6
xKFLJ/LNinrQpKysInCZUZvUQ9MzntQlLTghNHx7wQ29cF+wxqKKRcWPjq0ybNUG
av5qBC2nM0GWa6F19QqFG0necwonhBFwTQVvkyMtYLIsDnDjrAaZ87NzD0x/pGNR
I0HZANlFJeH6BisYZcSYVDNv741YQq3peV6AZuMxA1+5dEybIptFY7rgno47x6jn
SQ8bDsZUt7njslileeHOXYdlI0ytYHstyyg/P0zQhRv+2IYCxql06FeKfpxvjj0f
wDnk+LWoV//7Hao7qPzlZs6ZVOCaIHz+Al/WHSvPfk3eqcnZzhx5SnSlauLGES6G
e4Uow3L7Oc8caf74E5wyUtKd3x/HF13+0+jeZI3xkxVukqG9OouMsx6WAgqZJVM1
YiJEf/iDqiceorLwBb7qilJ6kDKJyZLVS1U3PK3a4BpFPAINB1B+oFV08dzSnfHT
T57+01ZJQlSaPsaiYQixMwZgMYXiOCOgE6v8BYyeU2KGeEhnF5/igQMkZlTy/cCi
5EFjcH9DHDy1vKaJH6+6ahe69ixT1E8FMxVcKcfPM0hGR0pTPx8fw02vaN+dks/M
5K3gT3aOzNXmtvyZPW7zyKrgABpRNu8V3x9f+rYJQtXjlYcqAxdxeJUusFMSuuPs
vvRaARJgOQSao0n3qvm7N1erLWxuJgXUx1jP2d0Mcy3KtQF3d0wLP6DdC94CJ4Zz
y9MhLLjNt4MUPS6upsYzlxyCBTa/EajOwdlxe+oDtVOtp5wOCqCbEsTei/cNr9Ba
VQ+SyA2BEtmoCJ/hs8aKwrFEqYwiryyc198kmaV0sV+lt8HiKlY8DvBVQc+A6kYz
qy1HYdwdojANikSqcbgwlbiea+ET21wEDaTgIwkXg6nF55iND8PFd9lQNSMWki2U
B6qeNGL6Ox045CapCiMxiuSmCsbucjAUt/e4xdlRiRwf+d79yUDb36essSpnSfgC
HVYFrugh4f2NjE3zDKGfxh4zMBMhSqMw5pL8u1ns5oPyFa9zCX8BqXJVYuVDeZZV
fNljHc3AZABUSaTJC6WzJKskj5Xno27AkDY4Zt+YXubSUNiSl3/rSumi1IuW/XwT
+SqEqHnUftNnu9Q2sR3meI6YRSgqghAoBjrpz22m5UsbJo5UYNwDElDUY0abIgwd
jOsJmETOE7y7FUtSzrX+h3dZi/e8diQAs5I2u3KR+K270LVudKZ7iSGtxLaLzx5U
A5hwlvmTPW58EksRdMA7nzbCp2wQRRrNgWbtzXYZ0aIHPOBxTEtwd3X1hGgF2L7m
czhbxo3AMpVHVJoQpFW6OjnKImHH59kvOFIWcYx/0Dmu2Wj9dDAuBOnGZWPmI0Ty
ZJ/HLs4ywjGK9xpglhb9X6cKi0yMHEVGC8INcWZJkv1GGZ2TA0FsIPwWwD70D5Gy
8j/8iuo+/H3BXFJyfssCnFbMNIrwqOKzjIZqRdhpeUd9P1t1mv7qHCDS+A4dq/KC
3JHpnVHC7yTYbUqKhNTHfsViUuR9At9FRmBouB136+JgsfhEUEqXpOz5hAbknKYt
dGMYwr0L4j1bqB/+PtugGS0JZy21iogMtQZzDVCQwbXijM7L4sksGD2xOtvdOpho
AiI18TSh1N4R8Hw48dtRi+X8aCSgni2LnGG1zH74tWSW8sQf890/Bpr2FhnAsgyt
j+iDovxCOiAp3NUZ+y1UV5aCLso5bB7Miz0USpMKJMvnRAgKzI3/ka+T1cn+Uon5
xShY8Gg/cG+xGlFvy32zHv8ZlP7PWV5l2+cki8C1LQDxiBqB5nTrtuwvTwrSM6ki
5g/ciwc+CLt+xY526vCBGBjGGY0VR1l/Jph1YAjOHt50sMGd2vwpADmI10B3TRH2
gifk+UfNkXd2vvwZGmyrAjQiO05k53miUgTL5qZwKO9kVrtIpyTLtkoIEIgWuMWx
HcnhGHXj7/rU386BsYeeHg58XValRMQ5O2I2Z0DR3nIUC6u8mwbdEWLuHVZpRxy7
AK2+1RdJozOqZp1CrGtY0MQpqoX/BA/uI+EP3Mo6UAY2vssgsM4bPXSPQe5DffRP
PDktPHGC8piD3PNYefbu8VI7cUeT5n5gB0BQS1SRX5VyrJpZZn4fxoUVBGkE+Emp
Qz06Hxu0q/WSqXT+r17hr3rgwORahzrR32ZXD0uCyLXSVWsN70yeW5Q9X/MDaODy
Zkkn17zNv2Op35Sj6VTBaenCDGy+ZSczWp+97ffL8sGkT8Vn9d5Psg/KHi2KbEbL
DHFj8pSmlVXeW9RpdcVE5NWhLK81i6Vl/1jSYFLksyovnR7mKo3ySAyEqt61D11Y
CMIE8xCjWVDGgmUkVwDQv4F//nF2I70MbltZtrc+t4+sl0DJeCTaJvMz7HK56OS5
JQwoKo5zT/B1k+0dLatZelOgqKUDAqERP7eo5qyoUxAO+Gmg7am2JpZdElfs+jkc
g7okOL453nmtRqE64/sOdS1StpstygKpNR3gFp6BFsv7LzkrreZgnOo0zYUFgUvS
8KxFDtLCi93uDXtTaGrQngpdrbs/18Bw4XFzlhhR51yts4GvVH1dvKJV21GgR6dS
9QvNFV/Nc5bw/Wtb73NmQlISrjoZGA8ThM8VEAUI5FXqf5D06Ao7GIWpCj8v/ZgH
yJSpt4xg8AsQrZrQ3ecOJGEJ+ijdCjBC9E1t+um70TATQUa/uvJdVqyg6ZYXpfBt
9b/+n54z+s9VD/+4+IIYpT9FA0C28LsMmfjogWYUqjg2DYtehZ3UPQivB1QR+IEy
zx6cUt2kVPhT80OeJSxT94K8cn02u+5utKJ2m1WW33b0q+Zhu0mUohRmSPYwdH6S
ms0clh3lO8seC9+NoAs+WV+7WRfrTj2WXMiM8D7X20CZzp+u6UL+j9wEF+pWkyUA
BFvknwYylzYXvSM41JBfQ4bractGt5iNRnccgCIBJ2cJDTpOGjikv9iZaySxZc82
xP94rcyemeyDxKCPiGl09Yg+cPLJJ9CMZNxszVgDi5APFB4pDudMkFxi2N/xiR2B
XT+7UvSWCPWa3ouWM06AXCJaG9x2evbEgXMSMRYks78M1DgwK6E5Y9BbN9Fa5C2H
83uDK6A1TOFqdaZ1zwJ7uRuuog1oEykysl0imI5nEuQOT4wxMmGBk0up41EJp8xN
gBpXJCvtAphBR+MfDwfOiW7SDCJxVIWC41jeXsemnFlVSg6mRx96fi+poU7tsL3w
L5lwE10mfve/wAaTcpIuQqdl5nMJvJ5ZzVW7QtlCuMvX1M7nXHt8Li/qhplL9s9l
Ic6b+pp0rj10lwOZXRoMsTT6ddkaEikaEmgtiWLTs2e3FCuB2GHYqmSvWwMZKCh6
wFxRuIuCM5Zyzop3KZmNoacBOMYk96YaWapimmNz70W1a2RnooDKkV4AxVezqbcL
FbsvzGUBri9J/d2HrPxnp6qoVjG/rCcvhTxMETHyK0qf3BO3USLdXIJ2+VdVjQDc
rIiICjS5Avtp+zv78A4tH9+0ThbP0jTo+LnYuQ20CohrnshzUULcVatogRTWo7D5
sxxRFhZZFdVO1snN8z82TGvBA2p1qae1wUmMjOeBxw0j6tEk2PeBkFixgBi8ap3o
p2e6V3xvsCIzoy7S878w0NAUOZ8whz/rvaIQSyXlnA2rc6ivvfx0uEsg7CzfN/c0
TTl4gjF+G9+/fwxqzkM8hD2rzWo9bh6qblWuYTNZeKqWuICq2JBZqgKPuK99bTa4
0Nl4Mis1LRQ2kY02ZpWE/StHSzh7m9aTXQwOV4Z7zn8Ix/QlZvWLHpUTPxvl8RPu
6pQGCePz/a/Q9stllaSMx2HgAbeM69ANTVKhRJcBY9HTf6ePoLwNW+YhMQDzMtd8
Nv8EAYGmUczj4psT9P5CxHd/kdVIE8UfKDohcIEn0L17gEpF0pW8X1+RVwFeAuLr
YUt9V94+K+tvpVfBqiy1Mxyp2faBPSu7+juLzaAna+4p4YJawyZiBOHrD4g89EWl
AcF0rV4Ll0scrasoy6qdm/iRrBfK3TFi/5kNricwlgckepFnoZFauqhv6S5QkvTi
y0VbcyAql2fWq3Msl7pJzZsy8BkmogLwX/wHtiqtqYkxQKP3YQHY5YFTGhocoNck
2FvAHbm3s5HbTYB4KzzkNkk7P33q1zy4PsQ+PZcmB+9kAqSWR7TAwifV/43cQlpW
JHyd6MaV5zBwWbVOKz33q5s49rgdnNX1Z2k7Lzn8o8pXm7lWl5Wz9V+m5AlS/mnK
ntdElIamwnRRQIffer1gI46qnpIJWwxzERpBnO/9WZTHaEzqU+JXa/lBquHQEgxH
ha3l58GavLOwYhN2Xc27sTTaM6ctZTx7kr7Vmkyt6MdheAPnBm8QcxjBcWNcuNWa
ySOPY0rXcmzghYgSyc4rlll971sEJQxI46ZXD47NRVg3NYpDRYUCW+sQ/KltVJOe
zTdwHEItHjtL36GZAvXPLmCtAQeUbJRB8QuaDYotxAp3Ve9RamcDv7MEdOqVIzhL
4Sk1Lqx9Y6YBlMDiPcTZdqhJ/KN9q2a8f6doTZfN62I6wPFWymWYp/8M68mrWj5m
yQKAJEkiJpBA2jtTcmJFF1CLoUk7aAFSCYpWon0csRhM24XCaHSxJavgMNNzINLl
8HFeRZPJKaZ9ubHVCUlZVX2Ym6aCHYTxj2OkeqrgWamcAALat9VfsCxiAbCISgBg
HBz4i2p+VpanWYyt55chw9x52D4G8+Gy+nXzrAV9B/NY0DFsWhcUoIyCRX79Xr/4
E+bsSkRS/hlKF4pnKBHwBqNCtnX+kCqb6bT0yocnCJj9dwHp0xHjZncvPg3vMoWH
+3i+VWugBZp0vr3O7dch6zGKjTJomrtFMyPVVKlyPScZIrKUOeKGNDvm/SqIokwT
KkBdOskc0NyDMCBg7ilyk/EQFC3rTlXgjAadFOEQBHPK/C0Zw6xeYBXwX+F4AO8I
67bnncy+pdZbDHr53/+/eAaXZC9DIn7cpAZT5RXm8wkVETXqk75Kg2LYImEZ/8cL
/6Ymx9Y7gq8kXhlbpsz1Src+1QLn4WV81eejkSxb1Fy2Txdh/vUGr+dbcpZUkvSo
zlgmTI7KZhOie6RoWFB94bHq6ZQCV+SqS+5HnIbt3bYUTnwsIrrSPxBzOTebALWz
CwH5gnyn++PtOSOnxGC0Ix2Rp2WuBv0GCoIgjIxvA+zjdeoseNY+uA/tSXV8Xe0F
pmnRU73hNU0i4zm9niAOKkKR9hxDvCkIAGjNoeGUeiKeSXXHkrALAT26R5BcJX9x
sd/pLFA0QYxPbq5vpDNl7zXaNX2VqJnPAFIclOrL45DocQJrOL20lf6iqFG3onpe
JcDH1HMHr2BQLc4OYN8hqm58hotxLyYL2aN8wzmVBAn7PzG15p/yQvT5K/xDHiNA
4WfnL3StpAZYlrCk6Va0uvzWmbzNsUw0L7b3DldeKy2opMw2lzIuDAF5wjpvWsk0
dElUDSFfPbKutu1lmmUo4Sv6deohrIN6IBAsJOWsaAHSpj/7PGecX20DiQAzk8M2
WlDEIT/L10U4LdVXcnMFl6k2yzWpryqcMUwRnaPVZyxpqiUAzqHtlFnl/qs3zOJ9
iVpiRkCKvgg63WoXJyHMAgi3UKJ/iWaY01uUyOsvm94yYw/SQ+krMpD+SnSoHkCJ
0edtKlWrorUb4omeuLXi1jrQDEKQFMrVmG3hRPMpbSk5EN3gIB779hl5xa3zeGbN
OxXCTh9uk1sHDSsvlgpKhR/1yfjd6EkfufxeK+PVU6/A+oMuTEcrf9dBZvOcMSPe
Wz+z/Joa1Wp7LpihTf5HsfZ+DXLrBoXupcL7rfXGZxr+PhQE8qK3Y7VdJ+Jx3L3+
UM9w8glrUesYU/6kAbZ2pAPLSpQRtqWkvP1OUYeOd4UZDucc7yy80s4y7G4q0ID8
xU20QrLah8oKZCf4CQL8aiDZZJNPJiU07S5KRjvcs98KTONEU52Ic+WNdHxwoOMN
+1WYn+rOCxUdrVSAFZH6pR2+n6uW/ywd4W7Y83jjNaO4mjSmJkacU2OsV7whv6zt
A1P7I4mLSHHYtcuKwuBR+OESsfX0o+t39CFWhlq6vnRU2MlM/jlCFFlyDv/lcOD+
1HITibIUA/XZwP1rVjOto1dObK6aicCN6Gz9wtY6h4zkh9O7F9DPrB3QnKbPSyX8
tz3Ye47GGGzfbSD2e5C8EBeZwsTQczAiw4fwEywMTabcRSArvGqlGLG1SovOh9YR
/oKI4QLRqmuVj6Ysy6PjMMzH2deeC7eGn7Uq+1Tslb6DABx8EA0A0Ee9XG+YgyLf
z9pdZJpaGSYV6s2qRpo1t1HabPPHcywqFMg10CBljje59S231pO6ZEFZ1kLbMjEs
RNIP31smmYSXdcRjX3KRRqHhqfHZvqygUgAZzqe+P5Y6Y+UhoQtK/G2xNi2q2Vsa
N+F5mDYVQ3taB9c8ZoMjocfWa7fshTcIMPx1JLtU2VaHpweH9I90NMIXmmc/CiHj
R1D/Bt3S/CtfMaEjy6FoHfJq1jnOvUMYB5ng9ZXRC+KUskuoWgKq6wVkJoqZBpDC
4H5X1l0dOdIjr47o0hg/gx7czk41kQCqf4W5qNAE5ZKj42XITHbxa7jRc9w4fOfD
+tJvJUvfgUFxLyPKmyh/H9y//GJALDxU6sZe1gD0Bb7YHk8QDNXFdRIbmISSNjBC
njuj8UxY1XOCKkLMTiJRrK7slILrZcD7fIEBIunLJCryxJ88QBb3IkHRfcickKBr
FIQcayCklxtiCkUTUJ1JGJKoQXtvz41IGmnefHoFkO7umKY8MO1v94E6ogimeUeG
E2uBcop11RBmkMY0Ju2d/aN7Zd/j3LBf0eJKvV3mLWNpAJ7ojMUXS1BdwReB5hXN
3ly4x+czMc7g9vbYiSJqV9VlmIWLQsSHM7tI1uFcHJAXFMYrh1I4La3dSjpv8WW+
SuG7eGooZugLV5o7KlpQW5qtGZVCrntPO/RRiI2eYti+mC9E2mM+HyM6V4zNo5rn
JEf3SUt2SC4Re8Djq0fbg6FysdHk4gb9XnfxgY+lkudtbnvbEUdh658Gx+RT6GYf
HyuMaWrYmh6S/z9mb9b0epc+i8DC0uQy5FTZUZMyiP/AKEMBGQL1GBkLCSXi01Af
ZnDGZq1310j/Lbs4j30TBpiGyrCXgFBHOPwUAANbGe9vkXuB7oq0zxxwxjPx7ryP
r5VPDbg0IK/NeClC05avzhywaGr2tCP1zz5WDV4LrOkR7UtZYYkMNmX/p/FMAIDL
71RMCKAGiaAPphaagqHGo8NMFEojmE5HSXNtCOlLFOQGuaXLcEKHxN73o/Z1AFAj
Fn8OuK9zCIi/aN+tZqn/pZZiMfLJKs7OuJ6wGAG0n+FaumIO8TthjdjMVHwxISpn
r5qleHLTMyPYLu3dAFDbwNVizKI/ccTXO1FfA+7Fjx60s04m9wThIG3nsriYXCSx
an+PiBORCTMX/SWNMqR/uajIgA9xBusncCkGa34PvfZX/25Z16rsXYF3fKnapmyx
gWwmcDm9lmdJh8zVHZy/bukdowBmfGEyjBaih07neOJlZMU0DQOMAgwA59quW6EL
E8s8TK0sKQUgGDHYYahGbaPZMkxQKgt+cXRoKmt07Cmj1Q/tmPvS0yFdTMPc0KNh
RSXAk+y9KadyB5QGZhkYCZR+44dk1oQs7/j1i7Y/OCa/7V4SWu02//+6s0P3NQtL
ppFjlOz+VnPPdzNbAvMszW6mp0ut1kK2iYFxmAAhW7ikJr7e+Zr/g3lPhDLpVLie
h1oGwpg+RE0jovL3xNv89wYibkToRQ9NhFIP+pqhITl9TOhHiC3XiOd8qWkWfaXk
2dWQDgAA87iYyqDqo2k+rCaCR486/I69yul2wr/ij7cOcmeRT6Z+V5T5ELbEzrEw
TDTlHznuSudsB+a8fSl0L4bHoKce5hkhSzf8zCqv5FMvGYBb2gm0e2jpnAIwMtNG
6l/8keBeyXnCY0bYmBCWmHuWflVY74iWY3TvE+8rJy9/dgwNMZ9B/8qN+414xDuG
jkZB9UNMs80f0S7xWbfCys3Im0W+DyXrgByTN4D61wAeWAH8PmlxFvuPEKjB+R6i
j1ZcYC59J8Zwn3XzNhMl4m8XSJcEhtLu+y50VzjvwwGxgYnIVc1rdQMF1mx7MeHJ
+oORK1Swhk1ACYszWkl9YDNEkgrIpYofBW6fTAnyBnOsuUgvSYUTikepQ99LX2Bu
KRpZZ5Vt0WsBMKopK7FgdmGEyceSWLcN0ZONmTL7lsJVw/lUn3d+5ohTJZ573PvK
y2+0nWGoY3eSArZjlum/GHMiWS+CNiRM7RZuiGGEVa5PQWqwdv7WPpZWwCuFAOnc
rqnoqBmwAGFnfEaA9nzM1F7fjBh/n4O/bQ/9Ba2qQSH3LPvYeqaOlxRv27EhvSNA
a/c09lfEULIn0ARO1yl/mAekHvj91rsEADbHAEYId5SWVVQECJQvN+IDzVoPZTcN
A9L2dMcp8i80fFXcZLqfOFbjYqQctl3Vu76hrcOW5UszIfZmw34MMima/a6bbCl3
YWhF/yFTBqn13sdEreSPVo7YTiI3hjAlmSf1PwjmwlAIav2XaRK+L5tt7E910she
R3dw1/xfiNlTwK1ewV5oYfjwUkcA7og5AKqXF3eLA569pN1x9UlqGxjy3YZhnaa1
UE0ih40VO59A3KvR+cr6MuONM7u0OyKa/gIIJzU3kAbadb5OV+hiy2RZosaYiwOp
UgZE+Du+E2RnpQ40y0K0UuVQjCdTnXNb+Bqw/6Km5iF7lek5JCO6dXEysvfExOBv
TlTi2eFbue1QYEjRvU2P7d/UcvHb0l/iIprfQ0r1uBwNWprK7Lmn/pEHRTtc59e6
UFfjFHhZnrqCr1+aZNDGngF6jVPaXj6Bhwy+9O+XxNevucGRLsCIowh0CddcnM2G
g9xihZARyfUZdgMp2psRHSGDiPhJLirQ4aPIumXMHFc9oo94KMuuJS6Yf53vTp9j
AafsquEw5gXkqjaFbOlUeuU/s3AD+YTEogPcNUHWNLPrAmdGx+pATX7ntbUx/rX8
9VAQSRAYkKAvf2PcbBuMHKj7RK3nW1Di4FBvpQMkCWtbmsWkCRaV7Z76BBbHMn1t
xtQO2YzaEq3KA83yxepUMRCWlay+FjVwm6NI1URh0ecdNedQoysJiYV4QHUrwmga
omLdvyIRzaujBNzZ+uFGkcVKaCM+xOUwn6M+OamCLuvSqKki5/24kART/3cfepPj
Zl7wZXvrwR/wmnvKqmjcCgptQEo4jJ6I5jkoIfRqnQRaduFLy+xal9NetQbretYz
awX0YtOQo9cGW0oqTxBA458efttzJWnf1k7fztLCytEh85l57SMqyvPe2KRiS7hS
tcj3yAYduZOnxOTRMsdD4/ZGwcrs6kuvt/OkEzSNy01JqIvpgv9e1PsrsCto2P72
JAjY8vBI/bI+KV0kNdTczG4R5oSuzcTqwU4acibA158FfB9tLLwXfdHZvav/iqtF
cOymCHDbPNLgcY5gjiNKMC0Nbu234bwwYfFXXSxhBxVPE3nFhMbywEzmcOFu0IB8
96nJ/u3TvxLPVlnAfPD0NLCRd+1XVWZyAADrqFpm+KcYRuyYJCKTjP0HTq4ElOMM
x+PIAvs0Zx8lvr8vz2TEhdhwQZw/QIzCX+zPsK/FYotHVU8Pjv0KHw7zNN4D6Vgj
n8W9pwft2Sb+Dr0zkocGcCg+YArYiSFeNAeZ6bDP8W/KpHfxKPC2Wnsl35LSuefH
Tqh2Dc5RJowsGPq7pUdZ3TOveK1aNJbp2aT3hwR0Sp2SmMpe52RdbRj/s/deqVjg
DV1VR315TjlIzFPVMjc5v9fk6t76ygL1weMkk3GUyykjFpiD3Da8iEGy+WWc8Qs7
YsDRGvH46YJPAT24DyBkNr6ZRtJ8UOw9LZlU13pO7xaaBXDCYXSIHJCF7bOWfeko
6KTHSGVQ75+CytnJfSw8Xdqe9cg4ijhl/P0Aae2OCM/k1H0YR8ARtuas9Ii45a8k
8yKIQJp6qlYyZyYS1Hr6zitO0FLZFo50Se8osC/zTCw0Kl7L47uxpuxMvOJClLwg
iZw79o/NDqBedgzTFz7l4QEfxwlNTg+43VNMIoUXk3ZZHqLPYMXfC84pcdAVgZtd
l25wm8yqQxfIrFoH9nOabGWSQ/lfhElIWImQkRKUadAczgsFH35ZdeeEAVe/JDSw
p7W0LKupe7j0LePh8HkK3PgDaHsQYelegfP/ZXml3Ci3iUoY9vVC8EMQCpwdNaE6
GheEq7JUUyOe27Qv6yRt+IBj7PtE8twh9dav9Ew2TmkuHk/mDGCZ2EXL6D3GyBnF
gAZrywITXzns+x/UZVcuujHaz/1MK1SXUUNkloDm5y4ylnVsY4qtGqkUxG2vOxRY
faSt9s3JC5szKPovjaLYAgEssGEtbAQZa8msef6ofc+3A06WDIyWp66WIGJwdFT9
Kx/vAagj6/G1AI1+iUI8sa7Ug6/1vk+2He+6kbrPwAbjrvIcjyYwx91ug5LUsebK
HFpjgfFCXVtuztGee5QJBWed8m+pdFGvQdmRmJSGbv7QgqviRYQI5xZPRfhKWtXB
Y0QnLSWcD9oZYcQg83L+vnx6JWNE/6HkZdFfL5zmYQQpmFC9OiXQ1SzPuoxoh+7N
2FclJa63SXErUZP0O+5CB06XfaBIQav33zoZbB3dtV9r+jVqjKmV3f4XI/IGFoV3
tWYHRLMkl/3gEuS3alFOACi3wJYQb3sZMchQBP81jdMd79/8aMODF8s4Hc2sC65x
FDS1h+naY21pKEQdNuAtFZTuyJuHCVdrdgw4KYgzHCfK766x/rHM7hl4yBAnTew0
v1GExSH0rk1RQbJANTI4mgK5N6q/3OmBo4cCjyLZUsfvNlIVcxGOGKK51sXO/POp
hYCILLWZtkJHHCJIHobVIH9qp2bphwQNYx0wHvJj6yjSCj5iVt/wOALfT9m6gl/i
8JyVO1b/JOLQB4M8h5n/5H+EUI+8uajECDOjRCCRwVll2eGy1CcntYRjwLLrFwmP
dQkIjYYzjosX+J+ojyQnw+Vy555EaLFLwNu9LWVPdlMqV4lYAXNKmjN/32vzUzIs
pGasl/oLZ6EAw2ODNu/iXc+06Ck42W8T+c1qzUXvMXHESSz3bSOyDDLykTvWDTFE
bLn9mllO0l9C3HchFiQ/2kBO/K5VCF6ik6fxo2bo/bWy6xOTK2jt925hdL6WuV5s
HsAWQB6Eh0Gw+YzQWL19oO+ip8rDeX1B4wX2e8B1h6VAoEBxn/aeMxszWtaBxIot
W1DtB9QVQ1+nm7IGcHu5+N+R6F/vArXjckhSjWubY5k768edV2ZRcZ5doGMwhuIj
DKnOWvKE3wOjpoXxYoALqy0FWHN1HJgNT03SRKWRtqVj2v1vY4ScEa9JasqrqkQ1
yNhwqd1N2z3O6HVp2WeNHprJtt261xmNz9sYS0kycy63FigD8Cj2PTtjJTmE+qxK
MJ5m48u4sFieEUS8JZeEJ0ZCyVClk+C9AnFfhR3QSfWjLWKC1xE0OBEAnxPeUsR4
AvQk8MtfL5VbHH4PiocIfW+3iyF5rnn7R6/9NLyEp0aKv5MXYZlCKa6cXNXLNDIb
qCit/1QZAvtxTTeybkROXiAzV1jGqL+nqB3zHnDess+HUAhE6VReZXtEpwVdVEHO
FG0X9/Q9WeO6LjQgzVjgbIqFvRKRWfzgJYQKI2Qsx6SaWdJ9rtZCoAqMbKiGRxsU
rBhYetsOChhb1hPpnkcn20fIvCbynM6dHa08NpXp6LAanJEfQgDvJE48/PvyOA+a
9RZUD2LVmsiLGowLXS7FuxSl8ALc4bjfd9eiuKlRmUsDNaIIftBcVHfer2YOCwg4
t5lzDJxy9vRrL64rNjRddYAibNWksi1tobwr5Y9tXoP29c5CrVXYiQIVx2OXZjUV
18ovSIZ9t74tCrLFcrWZhTNLrjo5Yp8jdAbp0r/GT9BnMmsp0nvNj9IkiGoVHYRv
q+pXkxf/RkZbu2E+eZqk+H/ax47Xw/ANGfJNP9t6H95IKTkhV6VGnxkjDnKoykVt
RM7Uuda1oaUZ6KMkoeI/zD0eoEUGhHX1ky6Lmw7rPRcXc0DuBoyCcviIrPdAqvIe
xnPIteXoOpxNGUvr4AmQJIrpc4lbsjsNCBZ7OqYDBamXHeZjhyX4h1WBtEpJRpQl
+Mt0xx9G7ARkLRreKV40YI5KtbrExJb441e1XNQ1QqEFFyO8r2eWTM0Et0QI7zQm
QdpmsuXiY7eFPxJdTmNLLECNofstvPvRruw8oBNa06CoMa18iJsnxF/0gdFMLEON
NksyrK5G+Cx9YGNlLVW4VXeTtCjYKTUiw1dUFoPjJpSTLb9cC1DxeI9W1V0XDfTJ
Qgg9aCdHvh9D9Mi9jupW+G/eC4PEd+2gE+CJSzDSMlT4eRLdh4zlk1G4Q+SwoBi0
TQg/UjZ1pQsccS4cfhzCN19mBodRw8e/NST/xpzVrg8mPCXucJmYP/w24lV9+3/J
hImENkWAvkp5RxWYqv4NHRf8TiYgZiTKUlumMxGvUBsLD561lHO/ve/3QNZcvaLu
CfDcMVZOnBOZEoiKuP7spFpOMO/3Dq1PNWcf8lw14lUZFHW+78FnX/C1b/KcOY8r
bhnfW2bK4+9XvIoUHFCJe2zYk/CavZTSioVMh0mz5vq9YYNCGMnH5l3HQ2Ghe4xr
GfZJf9Tvs8MGcAZ5bShjbg5BQLx6fpxiYNh49hIaiOHwI85rjpi4QuHKnEdrhTSK
+Ml7kaTAcVvA+boY+g6XPqJEuWVPlKZA4TyxqXNzV9EukRG5rhGwQWBB+5CFLseR
Le106H/sGXa1gOplSo3EmkrnazlweGGmcSkK91KVQkbePROvYelcgJZeEZJ2MA3B
cBDTrpD6NLHI1X8it9pyXdhORrcZys2IIHTBMJlBPA5y+SHcWvbUhZ0tveeFh4CK
W1i4/xJBdbOq+j195jyMeHrjpaGB93cV+vn+HCe8RKRRyRQSj3Tr5tZd4QQEWDyk
HBXJnuMLMkPK4Nl3C++uNBS9BX1m56Fm0jdevRpUDwBpWShSD7z+jhtsTyGTmqNI
rR8QNO9HEr8zNnsJ64x5NfYTTx+iKLOeGwqYvCMRY9SVBPINEwIBX7f+AdHRL8+s
dNoHxGO3V3+s+aPuW+DImk7bIaT/8MLSpOm85PuKZLlqEeneMmv7Wis80FZAF/A+
XCXRgZFByfrx9yKNMqhjpivjLcNZivNSt+/Z9pMumDb1daZjP/lna3YfyGxQNJ/o
59QVNzigFrk01r479eGYpca7LebJwD1ZhCyOXqfC5XAMAshMEivFe7xL4kBdu3Z8
5wQ0c3+k1qOFL/2TREIefNSNcIHrGqkkAueafx2dxE9dgZFRBDDrj4laRhJlbBRY
IEfQpshX/1RVDGTDRCMvDyKu6/n8AyiUNoL7pYAybxOm/jo6tKQcBZuOb7XdqAAh
FAIhsnL5xp14TXtm6nHwD+l53SHRJLN1rmCZ3hNT3usQmMORZbA1EFkyMaDi3c8o
7/g4D77crpwepbb4OBN5IrjmybDEt/nzbfApox0otUz4Kw5YB3oRrHu2hqtZksk7
sAm3qVTVA4BjJku8Wf9oFEu7k87rM+8bTbGJ9SFU0oD+ODWwMAC6g96i4PpLYoKg
l3t27Lkiiq6UBTcf7nZn9moo8cfRJUf34oz5ZLj+IK4akk4EwnosEH/9XlEG1YHQ
Z8Efs9DSwdc468kqR9lbNzZYlBZYFwxODyZaMwHkw8kba3FBaQotENVR3YzJg+7y
Bk3su0xfsTeaJ01SrphO2iPKPJRqfYXdNLOKHPnoWiGazASFakG9o6CQFV/9K+lG
H+huv9KaVYSTa+MFMxkYTG6tqd3mIvuTN9Mu5oCBeRG4sOwF2+nOHYGEhvSmkyj9
yKYYc2aoktMi1ll1MuF9kpvKzPKe9oA+NG/CmoHD+CHoRp32mX0cbcF36a1NMU4S
5rcw2eaLr/w88OXtHCFBVz15RevhQxuHZUKBC2xnoN/jqXUTVSZ80VBlchHeRYeD
lNYyiiyzF5vo7tq0yV/hncKRmTiVpOHbNcJUMbsEfyt4Go1iOX29w+DKAe9VwMfG
eZUreSQXzD/eW9/ryM4FIqzvQxoHbiM2cF5vK7eQtfiIWd/WKa4LjB1FewaJud/u
fs71N6nfxWx6ziooel3SFw49lYySDPm0oyg1X4UOPrbvPrhFgwm5hRhze/hE7r9o
7NsIiP9QxxXWQuMKYYj2tPg7m80wSpDhWEMDGSX4JX7+4evfdXGzYYh33Cw8c45K
8RgG74MPGmfDrQ4qAjDfdlLOyLO8FqpwyFhk4QzsECTLbm4HmjnspDrPR7g4lQnm
9/2n+x+J0UtjFuzdsdgl2NaYeMzr27Gp0zbVDt17MiLSIb/FrDmq3qQjwRERJjK9
kc3wqY4Y9eA6ewYe3dKk4jjzukx3Sw3yDazBDo3r8khY6UpP0q4V14fki9UHImV2
qtW/rucElUbCEN3YFcNRhmZJ7bkr4eG+o2SEH6vWt34X9lHISK+6lVzhrE6h2VFQ
9FEPGDqGjbJKf7Ah+kvxPaMnZ0hUzPxZWFAeTRHY2lFd2b+97NMgCwdVWuegWgHt
jDBXCy672EwMWpRUjvhtvRMSMJ6Swo4kxfJfSvXyIw1FhOXzYrxO0axLZ07fN4SG
qUiSPr5S99BZDztDC8D5xw4P+l1wkuJ0vZX84j6qpw11guCRFZO6XrX+2AmywX2K
uW7eamvSCDccWjxlxz8Xwh92GbnwMH6bovwM2A9DmGjpg2N0gJKpcJJKTgEtvmZl
+727r7uumeB0MjloOMiAY36o/3qUhbpO5SolE1AjgJnTSugy6zVqCnO3PrJlDEag
p6R21GW3Wrjkw1zKSFANFcxI6V6Jy3yogT5KiTGxthjtmUpDoKgUuZdoExF78PND
lOebcpnJulHKKThhhQTMvc/v2R0iSzDRebtKfg2qCDA+WBIOScAcxyy10p+yh2Wd
R0sOJT9McyDRLWBlDa+f4OsDj6B3gArVBlbRpgHz5ddq6CezuyuxSK4KURnFXi5g
2MX0gcgwTxKZ5DtGK8Ra+lmaDa5Cgxju+KU6wwQg7VPHj/EdcT/x3LlnilAodbr2
06Ckq59RsPlEkKELvYEPZCGgK9qpq+EGOdwmgE7YmbRQ9huH3NYGjwxLqQi5MGGu
N2x8bQZ3/CO/oTeUljioLKG4i0BDJ/9tz4a5KCial97CRmqNB4hJEkfKcvCVvY5F
luHzzXP4cDwL8ilBfV+ekdNB9KcHj9xFwC02XBmNub+Cv+XZY7HYTk6W1rgEs9ry
ty6y+ib28Rv8nDWOADcX5rhXND5OJI7ijZCli8b0+qLxOhFxNHU8Gjj0egcK/H3w
KKP6xcGljNW8j4fDSKxGmdDRx2J83jy+LrCSPzJvfR1dSJ3BUJJitvnJdkrGPKHP
dHmSWg17CMC2bsYbq+dRukm9J6f1eSGXI/KOsaeORp40j+UDBCo/P4MnZQtfWk8w
Wez1e8taNCi1KDq73kmWo0qywHj6e0c7pEkAv2XI40vH9+xe/OeKs1JKcnp3S+B/
yjGIK87sObV5BctlWf7cNJrc3vE9GJ+FFp6mbUmIJBHBmEnhhh+4SIHwWQrBPY/E
b66pqdWdFrymeFZ0UM6Z6ZDbFqaSzOtPGNWMC509GszVptPeQIf4+FL8VDYLftPD
jq4eOHkqEdujLjY7MCz50QzK31cYe1Oh3B2jnRQCiKhAXEOe3Ms0n4NnU0GqanyB
Fx8KfhoI0psvlPlJdcxh1SEMpMApNF9LOg7llpuec/cEHpc70bhqJ7Y9KacGfzoO
o0vaYGGxJ0bo99v6n0TlxdKlp/sRv4OTEhQ+zolXpBMPeeUJMTuTkk1jq+Slre38
1xV3+iQtpJuaE8XAZSTapDSukMqhkyaVGs1xkm2QxOC/6PYHSM+l/j0S9N2mQBH7
Zc3yVV3Pa9z6G8GwX5xkBTp5P7YI8ttbr4lc0l9e35roLq3F/chbr7ktLIGiguRY
+weGn3F7x2DvZSSLWHRGvJ4Fb/MhZ1uWWBdCWNilKSK6pdbldtL318s8nNH5bJoo
TA5zfzc25YhvzMr0rbdYoX5zVq/O1WROC39sudMSmL7eVjmRpA4XIDG9dBJNTN6z
DomBKhsaxa7WLwvvolYDV1cuNn+q3sI4gTnbvRExSdq/Hwe9EWorS/w9TSBDTefI
nZXne1T9exA4n8tmtnl/CMw0wywi2LCBhD2R2xuoAlwkn6ZXe79PPRZihMzb2dpM
IGntFbUV7R6VESV9+kF6IkNndSCObfM/O7APXsvd+yj7+kzK0Qc3iswYAjTLQ41H
rcb9o2krIEQcoEi2rK3dix5889qhNEULyDl8wSlVgGIs3nDTTEASSrBSM4W8MCJ1
HLj8AsNIN6gW7Auko74Wl5hF02sKyvJiCvLe9GYkF44mpG/NBmwD2np+GJUDW+xn
CE1lqCM0NUL0LK7sbKOBnrVGteQzRmxxgh4nHky4gV0W9raCyFkdY04NvHig2bG2
yOLUzE6cRKHXOO09umWxKoRwPKbxfSaEEWEry2c+fE1gCJGwwP0gXx/Zqb29s8iT
i5ESotHsC4uhnVrmtgoyVPvYqH0/RcGeBHk+sAVGiFs2CMB49NSzh7uUKwYQJ6Xb
GnFRXDTQkuPkXL0YpR8sI3KqRlSp4feYfzRv0DT/4TKo9pKIqTokAypO9W9YRgIu
QRF6oMdEGQVhqcYv4tinGyVk/jg1KHn8P4uAzjmw7Gol79iFYQ2/DeFihL73odtO
L5FkLciP3fR73UmxjqMlMTMV1lpO/FQdpup8ruojt6h+DxrbTksq57jco8VmmTUc
AByC7vwnsFCp5rgmAZ57+pk+QZVS5ZUHSHFHwzC4LvsV7TgiPyiGhj0UHs0atPxI
Ntpo5u9jEjAyK4a+riwUQTLU/3sB1o8qxwG3LPZtkdnfBD2RijIip6hexJgZ/rzT
lawJ78iczxOcrCId2NN1lXifJLeMKZsUuHCMkfIkX7/6qEyXUnShkhoW0NOHRnnI
dKB9bEnm5dxkJWTls43+hS11w7zkU7yReckRWPlPxVVU+sfR4iftHPJ2IUgFffWC
8R2FIRSpbZ1Sn7nBxFVMn+k4Qwy0CpQZBMZCevjFg4PjIuyPD9Jh5QDx9ice+Mas
3xNQcOzYM1ZePvPOvJQiF7OgNYJaQ4uao35xibZOWdm2cdwZOfEbi8HoK+XXob3s
+zitn6Ygv6d6no3tPQQaZaUm1Sp96uSVs6xxStt7tyF6Eb5yor8EpF2VzArlgyuv
5SRaLi9QV5qF5+Dfs/g70LO7sQz/me0iBczPHp5NWHb8yFv7R4k3RUG0DdeI17hy
fHCa//b3+/AI1tTCEP6DQj/YY8n7zJDF2eULylMN6tbaOi/WXvtGVwXAzBZ6Awg1
yGKHFD7HXZz8se/5k0IZbeasGgaO9L/Mpd0FDQ/gn2ikA1a/Jxj0dKm9ggA9macc
gHywV7U1yGxdgcIAXh5dYZ3OEBaMDKQoRvQ+5zEIORtcxmhFvlhTUA/S63W048Os
lXC+4dblA03QOTIuGXg1HUxiLUUosucCBF7SWVqZCEj/2Sfpk70cKxtmyKgwVAvf
LpwRpxINAjFwGxSdLto18iLFUjiu5FTXYMYV3FHcNBL/R4Qz4IxWldo1U3dofK6n
xEBw8aZ8NGa03RrF7vCvT9x5/zlh1FYNadLtyEpdGtvJQ0rTNosL0/ly+xFaQ4dx
6Yg26tzFGlbw0lrIfvwesKPJTCJUP4HEEQGkC58d82m57zdEMrThepiGyAyOXjFs
vMIKoPSLvWqB4Gn7jLH5Zl+LZOy3mVwaHBKl/xBhhZufMpj1guTuvtJwtCVyhRpL
QLSEG6BvGCx1nrpJBsvcwFHwnFzNnejobJByOwOt9erteMgI9Nl+jT4nRiwGxFsx
HK3LreCb4r3XwjlzrPSpjeDF97mGEM6AsA31W7nThUIcwnmkSBIcrOvfAMmRPKU3
yLnKvq3UL7Tg0LJ4bDXm9U2fGdjWu58MQGLO8pR6GfmuzFXZuKVY0CG4TXi4fJRZ
1g0+QdF9N1vaK/8Z20DnEqHl9mubQvolItfGa2lpD7bdbsEt3DYtjhO1S/t86EWn
LymqT1+DAOfKwOGFvyw+Ezh8CZL0FSPc6HFEFZhZa348QmXVa+fZVvKcohwBs7ai
5jhG2CqPjgm9i7m9QHpU9Imiu9+6LyH10O3zyCNdANoN+CTX3VBj4qz0xmGE+5BO
aPOhNHndv1ZcGgImsvrlva9/hVmBX3psZ0sM70LAdhABlWp2b8H1zCzb79lSeld9
CsroECEBuLrht+cJCpRsHrsoQZAE3LByuHWpqZNyz1dc75TEjhCZsq67SKZex3li
jDBSEaMJSv9hrPfJeLs1XfNXKbciKRcXG+Ihfu/LiYi3M4NJ7jFHzm4ErAvQ2zxs
VEDTLVhza2BERQu+rUsCmrj/srAulhfYot6ZS1kBjEaMWhO7QoaIWo+g6g/9tsvO
z5UXBq6Q23uMIAC5mTw+0xW9OKwAa4Mjfnwt8wx9ja0T6NDk9NUo0RyppKqthshy
0OF0tYRcwIf55A3EljpFiN/Auc19aVqxtv7XggU+jG6THWLjz2eNGX+HT67auHj5
ozl2/eTkVg0wqJergXKgwW4aXBqQTwn/i/QlYXpj7u8A2wNqmAdXEH6BN6sQ4zey
XRt2wRwDnlF3KnC0Sal61K9ruypgDRdVsp/9mdUSyI7Ofni/3G+9HguKonzDVhmQ
Xeqo8AccVdZggvegqVUeBbIDwdEjL1vvxkowISzBQcL8dJkMJda3piUKwYhSF/Dv
frO3Ui3id/K6iz2ZW8uAuWBs/jVgGUEwybX2DefSr5VMWCriCSYw2fHGInKgqzBa
fc3I5r7VtUl7u03vuG5cXiZH9wLG5UTQDsNALpIjh9c5P8TuRQEis/Uriab7yRFz
GZR1zBzcnzQ7ViUR+J76lOvfhYh32Seq6Ds9AI/k4z7WVaGnX2c9Fm2cqAlxv81X
sCaQXvAZNhTuL2pVpwPzwT6wnOMazB3LQgvt0aazs/tZJzi9l6O4OtYL5KW4r0Bw
0ER1jt4U7XxkquKXYabyAc+KVoKOUh6Fsqwyq2+2+/lk65JW75r0WfesGc+frPP3
PtIsXSvAu6zJaH2+uztq+/0QOKM+8DzWM/08JlCkFzyHblwXfnBDC+5+34dniHeM
PQ/sU2soOMcHQwpE8BgJmgZBajhJuIDEFneXoEwR5CrXgz/bRE5GPZGeoJYDrei0
uevwdeROcxEz7KICoOaTdS1rU76KDc8fqmnpbzFLsE5M+fUNHUS1FWjLLIrSlehO
SqlIcighTbvzzanepj/WOX2N0RtGEix5/hlTji+sI5x8puN8DXhGGltO+Ch9T4Mw
C1IFOc3n883qsetDZJ9IB8e9Z4Zhwge8Ld4f38KXo2S1PufgQyB5pStZ75utkrTc
Ll6YfH2uCE175FjUkiFELh5sqwjM82prqLv9LIPV5sspnJTtuc57N+lAd4c6NyOB
8/9+DHv2N5HM6vVnrLZ9LjEpTLwUEIOUTi1ht0hbAOIrrqcdN5zPQAtQR0lQc65j
+frT7rmf7I5GdwlRa4MZFsYPCTdVnRF9qP4RM8o2Lm2OL448lQYE+J4xs/PYe4Mv
hYGkTl62VI32nt+fK9U8VoOsSAeySs4ZDK+RFXpBeuz/nS7TXEWhYFundkWsivE8
txIcNtj19LhG8b2wFhsr2ZhjrqqyxD3trxGIWFq2+k1gWNa5Cok+eWWXyvOBjfSW
/mQlRTus5V9Tb+8uG4eycvDOoAbz7+gUbrfvYUzmjNUwQAlf87qqrmOSk+8vI6Ez
XC1LEATEEOrrzAj5nVwlvufSjH9ktgnrX/aZawODXkuVsztKfUhY0op/8sif7heZ
KE4s02B+oeGXCLed1GQyRCaEi7nledhe15Lzsp0SlvfdvKlkZ139XhgodJaU9mUy
jYRUX0En+TDFXMWEfWIteMDhRhQzvNGpcgF5n/8rIlJM7RYRrHpnGaVMCXSsURnd
C6KljJs4+BHhse3VESAXjkJ4oIQSVyLE2e0kRklBo8dm+YcnueNPM/ahwqy4yF8V
VaSqhZtNlUn488lYsG4k7nMMgN7fUrxaW+/FTWAOwDyaR0szZpD8BSPDduASDx1W
SXLnBarCG8Hx/FZml5jGULzG/9mZa+db17dvdADVWdWTvgKXENKQg247WlQHI0lZ
YitIgGGa9Eu1Gs754LmyINvwKZCqXdqDaF2rSWaqeVmKOucwOst/9XCpfqx8c5FI
VQrFF8HjU2QkxjovbIWxxDYu/XxVpDOfWABPW8n2E4qJM53CJwjb/urTWEQsM8te
3kABJhmwtZ8fcwcXfxA9yAyzfDp1Nwpya10cWwL2FnRxgOWRYBaUpEr3qQJ7FCAB
PCYQUIhARNkzE06z7czA3sCPNi8HL0VfsjHz9WUFz5rq/NhR9AP5Q9DHXq8BbXWI
8JwtB2Sep4JPiLkzCNolpSxpLQhWZN0yNde6fiUYbd2orZnxlOo3Y3riX4kLAZga
7eAQBEcMn7hifYcO6A/YjhuNyxH2jy9G6B1YQCYQm5yySSe7CvIGdR7WgSdmtN/O
OKerAoYHy7jfYRQlLR/AUbJEJc5mjnBTw+cGarqJvWsXhoMmhfMsLP0UrOmDG/ae
ZMhLQpZMBG6/sZHSbJwNbbj0cW6gyBjpQs4Z8QlsrxRCz27YjZAp052x7tDp+VU9
Uw4CDS6ylq24hiGyCiahhOEzg0cFb3fimvOFdQt184S74BcAj1OltpBFgDqy1IeD
6u3Eu+WrFH/S5N/anPNgRAl3xEAjNiXKaU/BtUir1zWnMbbnL7o66dtatSpPGo+E
benOj1/cTPEV+jFf67BZRxTR0vslMGWJ7YeHHTU8tAo8Y1H5c/dkkIxb9sWhRx8K
kkvupWAACLB3eSUZXHBgcuh5bD6rUiSMgn1aepOFGcmmKQevfl88PL7Ie/QPs2dy
778861PqueRqf+q+qfDpWQKEQFH5sjYfLy1+0utZpdM2ZmRdKI++hvUJXRgq4DT8
TDFi1CEJ6wpG+HZdYkiPD6dJOmVyZ7dJqigwrW5aOKPBUG1CE5bvYtgo4+ptyv2W
NW/I409ijysNU+58pwsUAVw5w06eEclqF94pAjJcQInBeur4CP2KOZbzajCn0sk8
UWFxqoJNKjGPsEsmIPHpo+7dyH8MNHgMzU5QQiTv20gW+pn9ovbxpwUJfv1Ip4su
HWd7tzeRmweagpBriE/0oKItmytwg9xhhQxFwPzhn6FCjzxhbLfHcyAvx8/3n2Ca
EJ0t08ADibSHOIe2bxMrEnbMB9/stvoP2+cA5gDDg7pZcEBFzFX59QblnaxRGm1R
PsIyDfcCBffd5L/kYDwfHA+UgrN65WXbR2MLQKbHuMD90TWpB/o0XWuDmYEMKQB8
pr8sFy9BkjXpfXZnXL6TgoHUPlwzuwcCsrW7EAPBJCBsPkTOei5jctDJRUR8BwdY
sCmwwbRW9daXulRGyU0W4KbOZRY/6RYUnoFT55SxKIUh6LomL148ZvNqdeK1zlKv
73OTbRYkLRwftSB49t7w/Oj/GXbF7bh4AP/gjKEST+S7IDM8JmCDi9NXFd/QS4wS
1MDEz2TsTxJdZQWfKTYkqubFB4sQ0fzbSw5bZFw5Olr3NiYVKkL7zSnZankkSSsZ
Y8MotveytH0yOYS/4AceG6btdkmrbbw8/vDcOLbm9ILFEu0lCgg5VfNdrLGFpb5m
YEv69lBRZbVt3Cyl1WzXuJL+IaXWL9SESIum6OvyyXHEsTYRZs0Hj0xAGnOwiD3a
lCYBeI1Cp+apb1aHdmZeGfVMnz6/h6NocE0Pz/tpzdvt7Xy62xyV3Y8uhq2ZFGKI
ybDeYflOeq4nvjBIMqe5YtoZ69OSGR122dSYrERiorOjrjTpGeuOX4/eBlkXOHQJ
HNff8VEUT1b8LaYc3G+Y8jCeWsfJG/B1MmH7ODkT7PuimWRt1YXnFI0ciWKEqE0Z
vepqIVq/z9MVxnUzw0AXM3f26W6sxyUo+2BeVOrJ8AmuA0gsmmGwEAjEvy5SemfX
tZxkOxzfE954ZrRPqDK5FrabQlBCK/2JrRGsW/R0+4GwAIyiI3xODsOCdRsWfL3J
97Do0AftY7bVF+mKY6e94mv8GuNJUgZHyzwxNFC2pIyZmP3XBe/GlxRFr608a1UQ
+6SxPqIcwPxHpwWnX6a+xRPYRGQwJWTRycmL/8DX9du2RULUbs6SARwvWbJb2fWU
neJSvWZDxiYtY9pNXajs2IBtLAsxStjXalkHwZopSdvhOHY3mjxEbbjv5MpvgEdA
zyNQjyiG1HQlzgW+FnCYgePGsMIgP3gProNS0GS4jxTs6TpF/xZ47exAwqkpsukE
/nRtYjeLovFNbubq7iSAj7mkCm4+D7zqK5ZaZBldKF+ZOQOtKr33Ge0UVXcxN3KG
XriA4eZkfiIhChUYSydPLcZk+KUWBbqWy8sY8QFtspdlPLhhl9SroCdDqLkIbK1k
Ic9gm+TDI83snkLYEncPZDUuMTpG9i8kU3VhqqoGUv3w6ygTjGvSLoS7P5+pBAqj
nZbdQmtE5gRqUvK+V+a1R4IRDpNp1n63sNXXR5FGcWEdcoiywbXyVxcQSpxZbiWz
WQ5iiyfs+9gSGjJlEPgAnCe884ao19NaC/shwhMMxA1SCgyWCFLsvRuMjdGtqLZP
acA3grvwy10DNXqdwqGdCBzVGVYsPdg3onRqWvXuOz4CzwWz6/VsCxSlElWWpvOw
iVxBleSmEVU+E5fByQE89YRLjuJJRfbzif6NX2QnsucOkZLrlX70YeIhB65tJvXD
FFlFdsP1l2d+Zua+pIX5sh8hJMQjl5GOSJhsYklTKOisZA1I9+wdvqpk1XHrIAT3
4IJTeaHICuyrPbkhu2BPIOJqTDD+aOLAr+P+5028zftuXCpCW2arrE0VyIWw9Kki
kz2oLXdrp55MBqnd5jtmpFvprmlIyJhVgiXT2yK059VlAjCPFFTxaKy/kNQhOQvp
oPFxqYGO36+QmmAz6QwnylVcPqDxJaUKlWcv5hVKKqTy3WGLpo9rEFeREGCRkAW2
GvnWCNqyZ7m3164IKf8z7yvEhRbmMtbNmImEmWb1rMKaw9C9kZ+lESdFfGlnX9hr
pSdKh71A0Zu7CNIzIMeyA2swc1ry9jSMN/M9K3zDlFV6dnvCz/BZdhoV7Z7KsH2f
CDsgT7UTwKzPnmPrLsBGScFMp0QxCvPxv8iPnKZauMaLW7kQKHnGwa5KGSx9B67/
dRStRhnm5ujsCRCxv81Bbp7TejdchwXrLSOxCF0bHxNIjUhhYJVSA1BB8Tq5NMJv
NKVMNtMqGzu5XdWLV4ZQDpb/GJRHRH5joFSAQcKAoEtMx6xI2Pd8yNLPwugFyUK+
e8o7qP61BxXB2y+tRQILWA8xH9WapJVIZFSQ7gyQj/hokBLI4HPIIQW5LjcgpWqE
F/+JEQsDINkgjrSrxiWA3FHRBwoDnPRhoBfu4hLt1LMJNg5zytp0YxoqnDxoIkaj
m1erDuidINtdNUcoVPGFQjsrxOgU2MUkPNzL4DS8U5VaGNNTN6BkNs4Ct+yZ/IA9
Gh01BGilWPyGO7+cnUuVMRPb4AYncW+2fL9oykoYQIRQpNKH0qTk0DTl3d9PgsPo
1e8h5Ds0FwU+mkZj3DOfYWRj9w8nqPLh2RZsBMV/kCjRA9F2mq6NKUYKssBrM6Z2
YaV+Dpbm/S7M9u0TSVa9zakJTLz9dYfDY2YPDgx/UuL58Vs3N6QiX+TMDa82YgwC
kNMYh4fjZ+JMoS90ge153MbDB+qeotebLqLy65awteOqMurD6otaJF3ts3pOD76N
qYApJNPe7div24Cyx4hze6oZhX3Xtj3ibEEB5cC3DL5GMX0IcERi7TJBlfrqyTqT
/NcjI2W3RnXMO/b+k7Xtmg0DLVnkpkskscH/C3sr2Xo3RIcq0uuOi1pe5n9r96A4
xHBn5rbJ9vXdXHHnLVdYaDjFxW360EG6YYUubACxCiR/XM+KGM4Jm5IGTWhO4Nn6
zJBx7WHIOeRZcSezOv+YzU02mMU2saZhIWRh5zNBiOgV9ijklmQ03/DnR4qP2zaB
Gb1eF+CMfXcxNiyZ+SM3sknceFVEaBUULFWw/EoU5XY6JLzz9dYc1L9Li67C5PGg
c92s7mQENXXfj4Mpx7oHSyqENTB92An/wkN2bhzAksIfOL5iFHTaUcdNjR6bRq7l
m0vh1A40GVSInq04U5W9iVFpQtNO7YO2bYFbzF5kk7K9qqzcZXGKklyhWrwCqk7i
byDd2wqIVdnlsD6Jz3bv2W8pESzMJo0V8nEcsNPIpr8XhksHIHUPHlN0KsWzp6OB
pQiEWM4EXyitcGejPq6KvzP0IJPZKquNEJobDYJuXWJg3kWCq1Nr3t00hAl8YenO
J/WcmL5lU3koTrcfsqtWaI/R3BI8YZsKmHwD3xepoL6/yNzCi1pk2Z9SP0uawGLA
Zej/zZTSSxB3c/1gE1SdP0fMOTxl/5xA31CFrAhFgPUP/m5H3inNJEiPwXr+JLrJ
UET3wTe8ebRrzgIgpl3Rqb1HiDCskZhmAv0yXBQcri69OphchLIfGbPRiT05r+mk
PYEwlNdb8uh8tseY9XZVJrg7MhRGkNXAk7cArUpc7NdvK6LpDgEZHkyqgtBNRfvn
2BcI92oiPFsFlad7UMtipTuKmMV9nfBdAm9QsxMcD/inajdIYpEQLExj6GL8hYov
exKuczxp4p1Ra69qvYacKAXnmvxGNJTFCIV4nzfwerxXAeF4CaFjVdY0votHriXw
hr1k/BJgJoAIo9j5CMFQyklliJqY5brmBYJUU+OcT4onx5usMY8/lM3aZvOUhbry
3WEIOkK9GMhepzxhZacELmWkTTpwk6T3qIgIiryQUFA56MrOiJkKuYE86VycI0nj
0izNaA4ArPIwQpwu/srUGDm508fnk3nX3HrMYBL0EJ8I3hehOLr3OUfQA945g6tx
PXwnDNeG3ofPEjEnTMoUmk598GjeEezJmv8ia2MJ7kR5uyn/5r8hwH9xxAG8z09H
XRnHEllXKWs0rTwp8tVn02tScIRlQjp471Dxqm/w0mbPzuLRbvxEHFzt3w48TNva
gDGjNWYp5fNJ9dDE+Yhv2rt+FOYyB7r+rrjnwMXHIWajR8sK+LrkZ5nHzRHPpDOp
/+5GMCCb0RTbFbi6PUTu1BZwhMB4zuLk7NBCc4LC0eyrWgP9DbtQbT7Yd83A+JA5
suZ6yzIsDO3rU6FOfmdH9KnnzViQJj4xL8U/2H2RE7fPWG3Cf/djQuzLI4iTXczw
M5ox7Q/uu4cCNTxaVhbANrFaDnlR20xU4pmTuwcvwWWCgNJYunhfPmzI9iTFWgv0
y6a5REsNEJOZb9E38PB3fQSEr1dhUL+fsi61cvGtcOC1rf+KdQFNDM4kvhzvUd6U
MK6I71sBMY06WsdwQSq3DxsdAk/cCOC/oA0zGcp2/MPbP68j0gDgUWiK+Gjnm2Pj
B0jWQLSynKsgHZOj8aq96faeWNWlXPoZlPLdp4HST1opwM9iMrbf95T8i18La+cJ
tC1YmI9aFpefWXzb9BUa34rRLw0KxetLEhh89oNH+Nt3VboLpf0rUTs43rqWutin
qD7/JyRPjf8LC0zLl982AzsfBKVWbyiyp37l5U4ELtkUVyKSowU1dq1k4F144+b5
IL8IWJ/PSfwSG+JjSolXPMz73yfn530i07WtKjlSiC5ywyLf2J8urlrXT+JCGSz4
Pez4C0Ff0mgpWzVdOUlBMsgChlpGJU6Yp3UwrWHIYxtgOCC/O6PdvsryO0HpOk7q
cFwKyz3gS7BJoGStw3ExIU8Tqy8ZIKJCOYEBNcA+hHzP3oEqjSHPmrAJJCH9kUZv
1zLwG5VRqdytmQIgTmKQNRSPJYiL45KOLYP5nBgaggPDzJbnQsFIlijazBIOLNTv
vx8Sosuy1NF65N2XHeSjqF/EJfeCYux5zw4FsZdXRK34RldPX+7PHUHPPrSqklIL
6IqPJC3KBXxvaE5a+qq4zRfSaEeaqXUEsBUDeJIpAvOVvf23kXEF9E9iyQRRFG5V
viwlHn8hk3UWzi9bB4+6ilD+PmiFGSgTKG/tZ7JNmqTFjGu+DoZbWYL6rl8/GhHQ
Mpnh4jUlkcK8BGjHfVQ8le2un9k2ylJeyeWx4nBvCT68fLI6Ka6mesPcU/CTEqdk
rvtlxKGthzl778R7UoBr/fQgRXAyPWh9hy/CP7n1qI+DZbdaA3fEn/oFlwg3gBX+
c8PHim0T1xf0Qt0sOzqP2EpKmScFKmKXqlT56pNUkQyERPTcBrmSxbxpYhjEj6gO
MhRmzwW9iiIcTHX6G2QFJn94iA7xdYCbd5Zdb8ORKNCOuFf6Wg37D6UMcrp8yd/7
6S9LLq5dzfdzQ4MA+3t8eCdrA8IriwOLRj0NnFjOCwd+kSnjqHAd3XbcBP/lFrZ4
iGcknGncrfm3LuJDpY+FagP2TlTLG6f7T5wLY5LC0MZtnvlMbm8vb7oA+wtQF3Dk
dZrRwoIOxn26WxkQHx5g5qTPB92MMedLVbPNVBpntVfzXjEB/VRQwxkx3UMQWDHf
MUlonMDyVGPjnzh8scvJBjEmkgVRGxRyG84IhM3joF2wgYZytWfrjlxP94QH89iZ
UWfOQ5bJTCW5ljR+/Al3p58isnbAFfC77i2/WepjQD8nJWnrEFxrngz1pk/z1OA1
zsavvkS8j3AFLKv5q1hbOOuroNCcNYVyx1CPk3yxEM5X5wJ8nD2Y4aVZhF2/122R
VHtcV32HYu8fmbXBCg4wMNYHGb+2SFjzEvU5q/BV7uT3x9Texk98DtgGqZ+ybSdV
gT0diIyRGDtWSnkU4hrjMI4gf3dGtZ6xI76k+gNEyUnIwLn3dGY9UeM4KEzH5Gp+
hr31KrGCPS8IkScijgRYBp8rr8tikDpdbrSR1RucFraLZPgE5PVEtRJtFvoGXk5i
YJ1xy+v2TfJE+OLgiDgOK2dfxm+2fzwbCkP5lxv7vPHU7ibmP7wzyhIYvDt1E88j
zdetkdLuEuLe3v+Ft4YnIRRwkPif56PnbD483cO/RmNdpLlT50l/CVFzMq0kmc7z
dau55UzWmffgHVglBWibJdKbVjB0/5SVkM/3JJgUZVBM+X/RcSmQGZyfdFTR+pv+
7K9K5k06eXfYwGk8JCHWAUBS9Z1MDfHZT475zQ9S1I8qyHY9EDEP4mJ5m+XApwdj
/ahJ8U1GZ43ORTxOvOKqvYMfPQXgI4dQ/vhDGOLmTVVeU0xO7qa65I/KleUuMO4L
7xD5/pGAIIKNcVfm5RwnvF2DG2lBaVrx4V6D7fhgmk+wVvWy0aNoqXqBGaEu20je
irDUtIc13r4EGMz1gvR7rNri19KRScRnry51QGoMuui4tVeE8Im0j+V3GJ3mxZ8P
x/MRIqtwhxtXu6CIn1XFj2Aj3eKaOwJkHJIQUBmdDo7LtI1IIxTYGSZdT+oPjBUV
Mvdb5WQNwg8nuj0dHVevEPHoIZZFxzCL7VgnXRhM2m6b0R8Th960qgjZhs19beSl
hCPs3Of7/w8naG8FLfVhJHTXBY3h3FqVc7wsqG1mhm+sSakb3qsV9woh4E9uSus2
UC4l0RR58949oHCZ12QbRgdLL2KAMd7P1EEFaq8O2z0ngRbYk3ZIVuCu2RmzIQi1
6xS6VDfjmt5fM8Kz4o0SkPXdYlbYoS9TR8fi460NUH1++6uDIgZEWhQF+sa59v9t
abRzSwdE7RBBrD8xP0fjf5Ekgr+el5feSHGmNIapVWHnP/c+W30x7Q95kl3O4/ov
nSIp2ns9w6jo7DTyTbF93tVIRQB6L3QNgb77EgQk4nrD2NItcGrY7n6nUxl1eFC2
98yP89PVLBWSZ8o5+6uzDN0sTiMSlR7KTCObqL6bHFt5RWEzFtyKheHmPnOCOEP6
VOX9DZnhs4ayJUjIS4gybPQgmuSHoA7uDGT1G7MsyE2LFsyCtbLvnPaRZvwQU/Pn
UWmkp0Lf5RWD77Eg0rTIg5W2XlnoX+tbKavR8oUiHMKLCY0yHqdI2Css0CLsIZR1
JnosjFavLpFFWdM4w5WlTojorH5G1PGrFaCcft04ASYjcK/OR2vS+mQUp/exxaPz
4PUbLgVLUAlaYMVn6bBQuhMyKTH45ckdfScMAqvrPHlkqKnEC27G7lGn5uNOh4Cj
UM3le3l1nOb5CpKT/mn/CHGG5W3nmxuyYYZ/r+C/oiAvRGzJZYQZKr8ZeRJhx+0E
52EIzH8iUy3yZ7DwWH0BjCQloyFw7TQHWj4Y0pw/owypESg7Y8bOujbwoL93dXlS
qWG0t56dNAk+qDaUI9OHj2wKzci/mnCDbb9Ng3/Hq3hTmSnFAI0qM6ibq2HMCCs3
8j1LLKL/iTBDsjaTRom+IqA3mSRxJEGlS6OTOeNQyNzV/ndl9gq1853v8btSJPVZ
FfKQM9x1deyK/5zLkx6rWRihyyqogE2vLHKHKgvv8uUK/GOHykF+Rhzg6w5aJXHh
LFbmhzdImqJhnNQ6PRkH5RRTLQj5wYpspgKyVSLtjWpUotF3c8GoBaJ+L0MzSLcV
UrqBMByMYWYE+KSd3rDK1DV6gS0YM4S6auc7LuhUD7d1a0Xt25bbITenkdqpoE2c
0U7W4Q77P7Z19ii+P0EPbp1sol/ewuocRmLZwrZb59nmPMtB8PpCjP5hroQpK34e
9to8Efr9q+WhUQqvW4BS8Z1wZLtryruKRBJACwGZYTl7h7/TRs8481QCyguU5Frw
vhPyu38J+eWZ/ljG481JmzpnzL48l1S2VB318l3wgCNaIvht/Bld45pByXdKZ+Sv
E9lClyjQicWbxtQVX40J8ytsKqTSX6AcV3QJEEnv05BAtWpN34h0eys9xF5yCiBn
7PZN4YmoK2M4nGhFKcmllfb7xpwrBrwjVpERzi4m9LRcujvZtlDjGpVc6BhCi+IY
pze/Q9gDsc5YLTNBLMXX4STgrvd+XQBut2kdi/aR7anwM926HDyKqQEUXtD5LdW8
MoWo7Cvr4YwLSHpSFGfqOYtXS1VhWQGthL6KDCEqm8SAsi671ZihHW9/vmgbN/GL
XRqnpH1BhXUdxcWmsgdyU/NZ4qpKtS0WkrKEyguzf+K2jaMPYorVGJIzJoLZ3krr
+qVKlRYYRDm7zKe+ws/4Degd9frExpxFLKnk6vdSdDW01+ixUA+gx2g8LepQ5JTu
StJw+gHBShKG3NZrRURHZDn2Y8cE/hUajQON9o+wQCjJsIzTxGeSWyc0HIIJ+LSK
W2L0CuXzKHlaqOODjIfWfs9/qByKp7ku16MsjDS6fLXw8FboBANfyi00VeJL48f1
SsNDBC4a5IzJqp54P+WcYbHAOr8Wv9BDr9SdrgjW445u+ynJxwjbFdfW3F/CAQIS
BktD5jkq+65FXzwfyoyapsIW7bj1uKqO6urklkOWNgY0tZ3qOzyKwcoooI1Cr8tV
oO73frqY0+9D9BBd3q3aaTqPWjDBSygZBK/PAawomLTqRMjGhqt67PEhnMnwfN9f
DRdB9vDmDd8H19XeJ4ykIC3MHMdaXaNpILyR0Xy0Ejm6oTu90IqFex8hSsk+H5KQ
JaqNkTZVWM0V95T4zAnzdwBnBnIvhRV6cE0AhkUCAPNR9nMJsNMFILtYzAUmt51z
u6j8j+V2dTF5//hW2ticfBNWfLo0l7WqI4S56mRFd7L/CmOO6bEQWH71Ke5kHivm
YxYCCa2sZ13LNr5ze6Z3tS94vmv1i1S47PXXz7lH48I5nrqUnLEUMwJ7Loe8Cibz
RuzRr4jVrHzEMaL7KGCJN8G+A51MpqQTaEVdOSW3hvxF5aOhiUR3/zI/cJOKbA6x
eyTng0eg1Z227pfTH6JyhAplM/+e+DVMRsLNCtpurEPbZ0BWBIhaIOSn7l2Zr2pq
4vi3uWgtEAYtIAUvkosMYVBqlYA0WoHsypzm3waZDbT2j7uJ9W6iD+bo0i8bEddV
EqcGibuTTxVHSJh5DrSbDykmJsBcaOCeiiFIIDXc1Veg0TImig5h/ev3Ycw1ljwd
UlRru1UqD6oRBe9bBN3agC079AGS07/QXxpoGRNNY7GPX3xKwkg2qr0H2mzjTxse
UKgw3zugQIcZJUNzkV6uQeDVSx45nYY0usP/HTFFZsfpBywMFMyggq5Gh2w9oTS6
vDPpkqiWw3kgtOUE20EGijapIOu4SVDJa1+LlNr8eDfHpMOGEmqmM4FbQ6tTyHxX
4FB9X50Qw5pGlkhZBUunVZ1uCnV3KUa3WCXzipL4ilOdXhmpsBByH18J6NIVM9wi
KKnJAtxzv2RDHuieyMzGwa5dsvR7kTF4m2EvTAGnzn0xvIrETrUkLbrxTvTyrUe8
By4OqvsiXYJ+4EKN5PxTQ1+fp+n8EtU5lmyJ0UN73tgddC5DTnIU5CVo1Dp+sph0
EIlL6R22ltJh/nHVyJhu9X/EnhG7XigBoAbQ/SnFiYBUUbHHzjeebCNsMy+ecn1O
Qn6PKUD4uG6GIwQ5UMlwhUFkUByGLuOUeeYzsmd1TDdoaINEORx9aywQMbMR0p7w
xGauxsOF5kB4TZtJeyAOV62qg/wkuvWbG2atIQXXd/c4J1vhDLiCDtd/hElxP9NA
XpVRaKvYuh0NQET0h2Bap+DL2xOTtf7NT9ju1iUCxP2uxDRTjLks+O+mGgCpsn02
ZA+0WXiOnmWUFRWVmn+G/zMrwZ9/f1WQnfuwYn6gzi2+4a2zGMVXs1r40KOJUl49
zRqP9iDIt2eC/0gz79OIOOdRSLKWfvd3hR77C+3FFuX/E+vbjaI8GB4grMIrHJBX
98FfoFuhqZumIARk8Ggp0RpOd2Tl3g8Oe/qQmWZRgO3bspWOz3FyCyrOUk4Uq0Fw
KdGcmIRj5Q/Wk3cNb40PRCsgKJAkCruxRjib7Ni6j852UGUkRapze2CbeIC9LpUv
a8sogQIUYm17i+dqJsCilC0Wx+DmupENt/CcllPunyfXYMVt5SGg3wxw2cz6fXuT
hm+EYle+pLB56ip8LgWkM2K38QPS+FR0AFx1rIvmbmBwmsMqQ3FS8AxTKxAmw5iZ
vLUD7Hn3h6tuJUASuMYGgWyJpMtoOBu7oyE4knWELK3D+fUmFDEAC3vxS9eixe5H
uYywtxY4+Lzc3FGiBhaQf1ZuiEKSP8cknDTQnUda2fWklUYs2yJ6aqWkpl5jwP0R
HpHus8q4TXuTHvfUdksthoNTPEmF4Gr9wQPN2GM15MmWHrSY7oBBIzUeeluJEryL
Rc9CN5StWlYuCv9mAUJFytbm7+lPdvXVLtwOda+9VDWzzMqzhmtasq3QYmU5JriZ
Y4YKNGpfdz7NjcT4MNtED6/cb01UQfTihpPgkmO8JswnS80Q2Cs5ERiW63Yz4GrB
JvUp0NUrgP2bcMoUsPKNoRlsqD84MCHFkmXWOm/BBvJBzk9eZ6S8Z8bTuLvfGtbX
BHSesWPVKVpjOpP9WElnKFMKiJHxT+Bn+JklUyWP00/qiBecm/r4e5GbFWhM+MBF
tVwtUzH8BrQjFLM+TPecQvme2Zugjxb6FCK1yPCTDDtx1kU6pNZZXTENnRxkkp7X
X0MTape0rTV+U5IFIkBJGq9oKJjNy35QH0P4FMlzs12hZJHfoviYOjNoewy7wILf
j+LzYiL7Ze2Sb8SNYm6cc6se57hbSoxA1/GasAM6P8PthX9rwepKpO9E4evzl/Pf
7FR0yM0eEA30869y81P8FZRgBYvKK7nwGFncswG+waHGxjB8mHffWgqtvpxQiZU4
LCzzotw/S/cVq+wGlHax1zPvgUfD+JoxSrDtcsjnUezlaYbvaGPSrHn7PeL2ZS1j
6uxy742uVc/3d5WeezN3f56UbsgDEeASg3/T7RBvTEHSwAMAKae+y4ozku5ZCmOV
Zy8drz6hcYIyK3QOw0eWjWUMM8MZCusfcEZVtIZh0GREmn9KVas1WMsbQrsnIleZ
aq08a3Vzvmin7koS5Gzx6+EvXf+/DQ8rXENB3uHJYu2Lkk4C8b0QGIYJt0+vz74o
enE75atdFr4HT5dnT+b7T3SKlaVmMQN6oX3JT7/t7+E2pk6gmxb5b9h5BdGoh+Ih
QpVHmecqvL1+9mLCs8LsV1wscQDdLscNfX5ai9Mmv18n9yojUCezEChtnJJvyg7x
o4Zg8sh8bfA+W8ih2CjG2II/vZ/zX1KMfx4DqH0fgAA/3RZRLE4CIzrHZNPjxhbc
RkK2Y71gVgaEoBEa/wbpsjwQ2nNgjlyz20XbHNT/M+Tw2itPP5NE3DFrzmBmuqVb
GH5MUitWed5LXa1awddaU/kqk2BTDEr54DFakD8PL/esUsNsAZq7QX3BkjWQZSav
ncPYHNM0PeFktgL7gWJxw0Psf1dRXi2m8NovzgUKulJjOSJGDM7QxjBdel2nqV6g
WfH36UFqKcGB6Ahti5YxUEKs8QwTHTL7sEM575HSPf6YerU7xuLWWcW4Fja1s2Wo
xh2fo17Nf7CpznERyDc81nicTCAWKARLQDwN/xYC+FYaV3TC4D9697ni1r1Rtlr5
ZFfMH852aGFyGWDHg8WKS49yDKj1fkbrK+5Og2kw5xCCkNb4I2KjvAsijA4zdqtN
n3Lk3FHf/GvrulweAGcfb4YMMxZ7w0wbA1ElBtGBw0WbEIPUEMa29Govg+NzItXZ
qIDmIxubAIc5qJ6lkna3b5YFI2g9GtOrCwwEhbh/hn5fw87e39WTGVAgIlJIyr1+
MFgPrQEDA6kq96pZsl6mPJ56q+tnI7cTMbmqOcFMNQfjJ28B0frVMHUGVd4iaUU2
W6pKrcZo3Con/RIpQ1Y+TmBf6L6yyaLKUGdQuDjZQXsansOIPXEVP8tbvxswf9ls
ZHofui3Al7QQwGmtZ6EMzE/2LAvyJALGM8T//E0qvVeFFVtWN/IJJug+ZvM6WlBz
UJLk0eXw0kqK1zENFdu274/sVIS5wrV5gtHCidt7cnVzHrCh3ZXTq7M0e08lAuQc
MKemkC7XWkwTzjJBkaToUESIt6ZKsRy/4yF1GFl9rOORZh64ZFIg6ysh4uptD6es
7KRZWo9PBGfb02uzDXQjVKw1U2avRo+55GRYitY0JH5vObpPIM/KFx+1jwyTbiv8
cQb5/xghKJapItCcwgKMl4zxMoqfpuCYaS2EulCdtyKY1bA3NBpvS+avg1o+Xl5P
yl7xLymOBxdTVX3wtFxLbcreP0Cj5lY74l+ZNP9GLa3JVFsdAEzkR/UEZGCVscG0
KmuUK4LNz+F77YsqPITGEqowQz+3FgxYLR4SMJflKkh9apM7819fZw6cnwJAOk0Q
m7oZT41nPG2fFjt+I/L1cNDkg/N1a1klrGiuuEKZJcNt7PA4T4m0JCWLndjMC9a4
CtDZ6Ck6GtVmTCoKzra8gsGJwU4iWuAuG9623LWkZp3puuOWiHKI+BCpCEAb6wu4
yy/B+EhSLZ1SKX0oC7lRcRiJU7+C7R7KuSRDM9SQuPhas7G3HwE7hR67uoFuR6xh
C91bG1mwSdn9U88rbDLWOvuj19gAH5xYW0dAOZN5OQeWv03msKEwoSARupDMVIDY
v5ahvutqA4H0Bisq+9tci4mQV8c4csFGejyMN8qrLddMRJGOq5ohu7jMZZTkawq0
hSONeprSQ65T50jh2RK6nDsk+jylcyAuUGfk2XfV997troz74/AdhZA5p1ratfp7
QkpLzuNzrsEtAggijH8YkGmAOSo0LJgkNsuX5JkUfYBAucEu21QOoMDPwsr05idM
7Mhc7d6OOmI8I+zIGib81Z8eKwwubQ/VvwhfSXj1F8GkH1Q2iB9Irkx1mu4/1Z1/
Ex6TgciPXgohyamJdi7fr0D3XXEAxTe9+joMoxrTkUHdtlJUhZ3HjVBaRMIFwvox
KNjrvAaSp5nhLV3Ic50rVtxY0S/I2HDBRLzHZ/4FRrKTPXl7wMD+hzZcjQ5slixQ
bbEd/PPGrDC+iDNnP7TzAqNORXkJ4XePBx8MsZsiDYDbWZ4ZeGw4IvjqqkiSLeTn
t/UHwfAhORHGvbIaMRWB40fBxnkFtgUINGP+5nLkFyC3VbTt4aynbtJvLKemGjdT
scitrnH0upv2OxYaHiFhwH94Wtm3u1KycdS3vmWXQLSdL3ceKlQaPtTuYeeRbaKg
DtP0HF8mtJNranetzJQzF+WJvvn33QOkwkDwchNUV+MwbX+8qoPDlOHmVt8bKriy
ggxiOBoIXN52YvyPNuE6CSQBYqXERflflyGoEX8gVXvGPqWLR805kJ3T7XCkpmDv
3XyrraFyplm1pX65/jqk46aOXZsZerGHq/F50Gs6UjppgPAA9rRIkev/pkNW8uuo
JDh83ZFCr907CQDzH1qhdIO/1KHBJefIQWD5WBs6CiERTsuv/t5VzHGc7pyMwyk7
8BHKmOmW4wvNtd/hULcrY76v6nY1zdY0aq52bzYMcDXRI/is720aLdDC8OXTIA8I
1xalq4+v9F07EP6xdqmzA1g9Jh3WjJ8cXEQ01KyjKo+brxrKx0xZZ2HkDCl73nsr
3x4M29WPj8Y7ktX4Lls/vFWLId8yCpRYg15pL9uOFCgltpamo/pUcBmHpzoihN+T
BWNFlw3Ntconv2Wa1o7h7V/R2eEEEH+qUOB4yMNpJsArQSZl3NCEMXmOJAV9+U3h
Y2J2NkH0tZOgCx85SVJThdpRbQkMLrOI48JOxRWKKwK4yG5zMZf04MsTgdS1prHC
jQPTdswuV/oNw9l87TMt0+MQWfxLpRRPzz2DeGuRuzTagl17dv9J6J5aAMLNAqGG
LPc1sedjL2cDJ/Ns4p6JEmvPsvPyOuZ0CjBEtLyZE2wnEl+UDbUPG8aRusntXG9Z
dGj5l9HorXnS32UBXKGETeA3CRhCVXrtTXTO3TE1ldVLvMs8QqqD56qFZa/RPq2V
8eMMlPh/kX9nYZUydMwu6j1dqNRfUKbGrjCx0HQy8iNqssBwuqGTpA9TmL13J1IF
7qsOqzXmmzTHHhcZEUnghaOdwlsFK3nNaSaB9AozCnZIpwLMrh+YaulOJ1EYn581
z1H1bAk8q4tSIFXlUGGKgKzqS3O+hTKK4uxJXkKbBthMP7s0tfVW+224TDi96pdG
6iKcqp9RKa3ta8/Cwl9oT54B6MCY+gq+QKKqOqZmlA4JgSeGV5Jzv0QXLU+RhLsu
Ntx5T3v9S0uV7xfBrUi7mB2dPZXqgI5h2mHngx2ZYYcLpbWzuSYR2DLenx04BJ8u
IDDljaZNNZHHN1Fybu8JbJYI6eQqSc/NfLsMvSOF8UQT7I3zrjkV9ArOkDupJXsY
g+ZOCooJtQnQwJtpSXAK63WbzvkyI9zYl6A+tlOLSsbVM8q9CbVFHWcGbLzFyfas
vN2GA2jXdLwHMEVLmNA4Q2+kEjYeQaE9zWui2DmiFzPpth0RJVRvDsHI4vsLLl9r
+iZzUfRCJ7RfXzV4SdXgu3rF7JLXkgEkA/++lsBDHyzKzqvQ/5+Qbt1MxemmfV9s
rWQHgMT6mrwz3obJ1pUy6Tx5VZmgJWVPRxGttTjkzz0a+sTX633ARbeqaANKglSf
Ck5KwYwek8L9K75SzW+v3yqk7L3Ibnig+kFDz21sNxWmU2QEhPE0NES/u0H+2g1b
z6+mdjJ4x1B3u3HPnAgFNcEallVxBhdUSiAiiOTePFdZRMMJPE2hm/G41JvxBVi3
GTXWd4fRh6UuFILOrBx9sxvrAerF6G6MxVup3+yg5b+lRdO7i1jWzanku6te9o+v
eMB6raiI+SfykFsvXC3mvxW7ey2qFcfIZ2S4YelrcJN7GQjaBqsPb6iklOBt5zQo
MTIVcd/M9FX3TIHXPGTL+jCxidbAf5lZkcazmtVC109zgOo1R0nyx1POG2cqJ18s
RkrR5T74L6Sfa8NhsRxbEgqlT2CzjPEG6kmYY9MHGQMgGA1A4vhDE1Rniisg/H62
+7Bw7lxgJ+sC6tsncve6jzfjqLEO0GUkHo1fgrzfyRXgqiRoHtKzT8MRLBAXUxkb
Byvo8qcKxOanO5P3sZtgrHAI5Yh93csZFokLFk81bXmPUIIePj87E8c0pIEt43eu
ggJRIgzk3mFRjMZxRo8zplCzcZ37Cf8nR/PohSdlHW7KaJJpcPswKg/Grl8+Z+He
+N9B9ZK0p+JNrQ9zNL02ObxE3Tqt19PpInCERnKEtOB0HQc5NTqHbWl5fHZxQmL1
SXQu8bRtwjmbi0v9cQEdj+5fUlDO3STr7I1cXOAB5RJZbOwYa4eeoL/vmkrIrlSF
Q99eq1AO6Hxb456jwNY2HDeAiBAZUybV4DpaKwXwKGBF86GhP9m/Z00UqVCmDi2z
xN/YRhusHjxTL97NkK1U0iaKnp4UXpvgQ1rSHlCOcvikh6eoLtzyEaUbb6NHYWn7
QZBfIh+hk+RT6D7Oxx3Gy6Qo48v1In+SgJNWFsUOHaomsOCzmhayT/CnjPJ7LFQH
TBfI0SG/cDVjOjlfMmFsWIK9iSaNFwphlf5oJiUtauVaS6912abIveHdQ575d3tf
ZHE6jb0ZDuTqDi3T6hdmTetZZ0x2rPpDwBxwRyziM/pR5U98jJkKTUFE9ucY4hCb
v/CnOqHMis2Q9RrwEYGNDzJb4YZtcQiIAMBlxcUXxpQRfl5xKaSxG3lZRPBg5HvW
x8jqEN7C2LTWNSNsVk+T94tUQyUI8EvHzXt4vgg0LzRT0GEYudKEwhURmi7MKxPN
CK8blY1fFgdMBQI6TASjxpG8LaUCkyXaWUsraoZlSSu6LA9BQRpPSos2MlLsrnrG
RskmvaSK+q9py5b6W3acF8urgFuj2PZiXFPmTyrYSNm0n9Y37R1lz3bvsS/9EhPl
gp3vMRn+oWM1tDERnHpqX7S/StvkFcXjT9Gev/exzvKtsOLq1xSezdOpuhbg+DrJ
G5M4mlk1brOfY4CF8FUrQEM3CYF21S6Q5ea3zvALpyVxivoma33A5UOzK38w0imq
Hcv0OnIjWbiIZ1TkWAtvyow8vsbLYHjKLix/vJqYjhcgklbeOnGC3GyO3Jusbs9o
9awAdA7Szx7o/RqcZ3nnewS10EUp3TNwHLrHH5SVDuI+MK3zi9zyaOJLvED1oPwg
ZIgdPtk6Z+61Ibr3yY+jitH0prX2nkyC77GGI0jd0OTi/QS9O8hcnZZ82sLFu0r6
gsb04A8ZYs3fTkkbNEA6XL19bBudAZpPXIhUc5djkoTSHWMr/v7vGrVtWwNh6AXO
0P7jxW1thtTi8ozHLR56NHe8pqsMsm9IOIPnn416tD1zJ8GA8nlfW1JN4AraETLo
urfQ55n6jfPSoPYyDchSt3vQSRVu95LKszZOm/RwXrR2vwvzh2U1eCy1PKHpEJxL
0mog0uGeNdJo5GJEZwNkcxptWWkZARA3kjeLrHUjVP6wfWVmasvq3d/7U+21kRnw
eSLa8Jdxl3kljE6IOxqBvcIMP+lFbvr2mtRlw8K+h5jZeGsAUI/UQH7wJB9o7GLl
Ow1WnOTQyRNog32/g2IPMR+7n9/t0r+S5v6kc/mIDoBdFa9iQagLqialVAovdMOX
ab8nqgZY3u+yGec7Va9pd8T2oB2FoR5seQUm3bHtL8QIq0QnsBVPThh05NMmUb8c
s7r5qABxZAz+eUAqAu3jZ6O5Uq5EGw9MBGk/aMYz9fFuykAUyhm47WDZ0hTcgl1K
/OVepW2/2hP+m7KeHfWw+YzVx3zUtCdH+cJMqNZe1odYrAHmD+2P/qbqOxcNrqad
wO8ohWqR4W86Va/oEDyZynK5cuO9WunFMBW8hjeGhZLTGaVQD+1tXt+ulgXee+JB
s4u0dknP916I02T1QEEucBI9lCux04OLK+42Q24LB4qBuH6CjavM5PDxLai4f4R/
QElyVqINF/clkR0/rQxzhWcWY0mvn1pkiNIaN+zpI29dgIcjz8kXLQAaB2bLsFeF
6Eo+/MBSmCtd3mnLZBAsqTx1TyvAqNOREtwoLn4cAE2hTLP89/1jb7+TThxSHbRT
7L/eLHIMB8kTOmnAXLdkubn6DJUPIZzPIm/yceeEw/qNqALMwKVODCecjQTheHn3
sV765gu6pEI1rBJvwOoAJMKDCNT///G2wKIcc46tgOdGfKziD58oMH+H5LWdb9Gl
DigsgqIJBPWEezndFA7hLcjde4wUjty4B/r2aZenrfZ9H4ciZhaxcmhhvta1dy+l
UvmEG1cQR4LOoqZbJM6C3a3yi+/RXEoEbxgH5YFkl49HxaBdRKYDA5tBgXEGHCq8
u7RZbTS9EjOY1C2gEfeHCiFBXMG3bkHlmPojAQnZm5cV4OF5G0nQC5+nlq5ozZpT
bYv/E928xJ6M3JrZayzGOh+bjcCTh5D6p0aHANTkr5YIRWxwl6JeRfntImfQ1wrT
cC+3T2lKPsXBbMcUWGbo4sp9eSfGyCyV6PCbTflXI7d2lNv0HCbYda2tsJsK0yxQ
nkoFr5Jid4GXQMKmSRNZFClyq1YdHKtn56nOOx7xtWH11MkIOKaYB4PTqIablY/i
GSZd6ec6oaCWJOSHcZr3xgtx5AuKnagDXtcnWGLexj6CsXe6S3YBgSNw4NGLPhyt
9jCxsjOUjSZHNgRyrdMQJS7eMghoyuCYE9yxPdp5tm2doc8SQX63bFp2h2pG7Jqx
NS0TiPp0xxi97PbxRfOvr9lz+hwiwdm7VRD3LYQbSYJNQhKrauw8ZlubWhz655+i
XnJT8zFRMmUPD48M8Gcg9hQSqQcPvboe6qo/f5XwguhNVUxZtZsyhZFlwDV/6gef
hrLxJSZpgEW5MsY3RuAxM3wS1E+Aa/3++/Ptl6tvSyhJjk1NnvUTBpPgL9/5UIbG
DP8bzucYV911YZ29v6Qpti+kj/NvA/q2em6KabaN09v9dyR2Z/h10jUWYAkm7lWR
UrO7C2ZnqRZQUV5nC7JnJoD6qPqyeohulZICl/QFl/S1wxNdcvwceVaO1BEdxEBw
42CBABFYNqqsfI8w7mlSOAxd9WqmeYQ3d4+Z0MG0rQ7bJr+yk4ccNQB0gynYCH5D
y+/kTRdEd11FNS5i1x9MTNr1ERYyxV7Ncjjwfs/DLAPawIV1XGaC0zJROG/ODcR9
gbTVFYO2RiXQxkeL1vbEyWTkLZvQsyteGHjDYGVspOLkS3ndShtxP8yc8dL934GZ
U7MSLjI0F9exx/iM6+8UPilgRjmuG9VAsfOh/uIHVJuAjJ52H3BeV/PnsSosucnF
ugoeQ+KMP9Akl670qY+4zyiDRCo8y9m6YqSvjHiw//jg6Me6TP6SJxPjwTpa2dJv
ApUEebDN+E4XzYYE4uxPdNYX1RVRppSNvM+DpVESIguQOnQir8lJIJe71O/9AEU6
2AnSzpiDCcP6PfTe3NF0Ag7xVwaCsbF47U946tOfUaVmFUkVb4Ylj+T+6E9CZI17
TPfPlaJI9tRg8VOWHZBHEWe8HPGGtI1KOmSOSaj3UFIi08g9Wdgru05v3guqdDmk
kU3ExSOy3EgIj9zLU676mVUHp4mv02K8qNiJpOC8GshZK9UOx4YcDJhrInXkoGFp
c2YdDkV1rS0W/GZsonqxL9pFH8prp7frM/TvQTSsD1bSLI+AT40jWc33vb1qoNLH
5VlBayObu1zGsebBxguCCNdxD37cplEbL0hF8WbkbfJMyXw6MfkdRoyC0Qp79IdF
+ArkUF4bP/0n5eQkg3I6KZ6EAMh/ZMhs5dC8bK2r0y9WRbmn+eEP2ialG9PJLirT
Mof+x1RIs5dfEYJRiCc1vMbijBK/1nXqaisICE4UDNL2cvaroP6bHHR8AG4oiGEC
rF9A02aek6VK7+HJck1zLkm0vcg//XBT2xRI85HdsQ6ZouVBaINn4iJi7HclWpFW
IYOrvviDGaqISdc4ZJmZ7SYrRVIkwowCBGai+AI3ylc77hMDt9c9WUORntAiGYPY
6WZMRZkSyvbkFDi7INfehGgWUbnINSCpL462LyJBhzUOmobZCo+Qog1/ts9D1A+S
rondIrUXFfuDxhQIO+/8+E4Qpb57VqczCC6tPc/Imtneg/46Mf1yx5uQgyuhj0X4
VgdfibdeDoTCykCDhwSxlH0nZ9XNkOCBMXUXcZvfodQ/WstOAaOBfrLCbKRFkStf
0f4dIazG5GPZ5MU+VkmgNTpKV8c4KA+RqX9Ax6W4hTCJ6ZdD2tbuRhJqVI4Ir97R
cT66fVX/TkEsx6TNmbK1PamIkJdCZOgtwzzJniMJtMHuBtA4K3PGkQmmQpK1+I59
MgTmsMb8c7aEql4+ZhDxunvECQ6jB/4JWfydGGFsOhISaP+laVei+AN+7XyTV9LT
2az+4fKaHMk7P2GEjfJyLO8lDGZnrAHgYDvmuNeQ5/cW7/vcqhRJnJvFdhq76kM6
0AJBCL1vuKVl6W+V/+51UyXfvVFCuzGW2Pi5ctGkaZxSP2RvDWK0XGQl85bDI/f3
n0T7xNxjU0JBU0zzw6CmBm+593xFtaG7wouWYhp4mwo8Sqpk1uW3pUlyvltBGobE
lFVXQVyiu4FJcsptCAhqNuB2VxWYiKcRGB8Sn8t75ni8y1L63iZWI7zGQ9dSshrE
gyvT50plrKBZPHro84AFx+LSXfOTkf8ZhZBQax/g1Aqrz2DEfBgiizhsJNfsYTUQ
MHMlPUGuAh5iIQ5mXHN3TDtS5tC2N883ybyKR3M8LPujLltAKtVjMhj2JNv8Xgvs
Awfnqsubk98niJ3NHqww64PAGq0BvjglX1CLdNUC+BV64zbaNz1lq4Fd8Csbw065
ESF2PoC+i1yj2p31Pf5HWsIuaRV9lMg0osACRRqBh87iPNffImea2J6ycrjaOdw6
f2zzoMxDrI5jZlkh634KNlPKBFBXx2Ssf3U5vXTiWb7FhfgwFAE5xiMqZthwjTvv
ydaXG3dBNvcaP00EZKHVrk4tKTb8Wdj2B1KEVG9lYSNP4kXTtql0Ziw7YlRCtGIi
Y+u1P/MO3/UEXBKIzRIPxxM+ng6guoxQcSJF/V+KRdQyCrP4+s0kYTy2niE37Yj2
Jqt2AObgOIGFdT14Eq9qP5ax2xbhT/5kleQM+Kxau0vI+xG1sr4FzUy52Ot6MiD/
TozzFXem+dT1MSAQyWYCX7uXb3zPjkMN3Km3ExII28tUtsZ11ylYq5eh6bQUg/v9
B9g37ZIAYGN1YuVC1PEE12bUaOP1UJXpKJZL/KN6+TqW7jnpBzN4RIghQSnkksvL
Db8VVq+oEoW+1llQxcYAoRh2IzOFiwK4rfbqFPRSLW5aDblK0wtGv7xP8nz4g6TP
joJJm5fVmpQXMwgkCYQJnJgmmRWQCFKOngUGAezxyi/afPwIrUyt23i0Woqwy10S
6vSaWlAaPcpNnmTNRBiOGYIy7fbRApF1L+d+6Fq8VcTvyBsuIVJeB9uZaTYf16cM
NrSPX0RTUS8mmq2wQFwZlfMOCrBAu8cRRI/eyqb/XOIMrxd05P0Z2h3GXmAI9A7y
eqvr0Fh84d64eBg3obl9MzU8hhU6QasV/qmNIOtxDfwQ5QKny8MG9UIaHUCkYB/T
ya0vRstB5rjbF/HvKm3s+plxTAQcvq0pSTuaILGmsdL2uS1+rGeMbD8gqyR0fz/k
A7MxIS9XyDvYDrszoxphuNgcvGCeb6yvGCMYm5+76jsPvSqvdUPu7QZmTzUH79Vz
tKwXN9VtAWbLGuYOHq29kEoE888LZoLMzb5kDWLdPPplEGhJFojJG5P58SdWXU7t
xzYlFtj5zbUJgL/sE7zGhmi58kAtfLFNii8f9euziNnwiaYtPeJQr1krmjiClgmw
kSrafxGEr2dzyIp6NwNMmvTqcyitgrrWPQbYQRuxm++uFSaJJC5AmOR/uDxrD5S4
9T4u5iruiCJdsaWc0MjJqgyqVTn0JdnEniTZnSszQI4/AOr6ELd2joP7tMNyM0E9
uV4z+XD8gdHsPxxKKjri7Q5gbic9AUPUnNlFNOYi7W3eYI1qyhd/JeEqQRMWNo7w
olGaJl+b60fIhWX8g5FGyJa9ftbpWbbTC8vmnyCoasVVsH+2hlxadeJLx2OdNjE9
SU4YBeSRes8dnIhfw7QLMeodvpkftJVtzE6T5gs5W8GmUTXSpSlCBppl9zCBAa8u
s0CdM2pB2GYwefWoxJ1lNSWB1XLxYNV2AdnTucVw2mE/BjywXQhj47fnGNEJsZOC
ByP9yWFVUk2IVCk5vmHFzIzG5Qty/dKLgUH44DKgI0yEDnnOE+wiMwTjh5fRUqRp
FDxWlxJD1+T0+fMiEQkC2oUniKEyu+mMuR96I7OuMceCwkSRui7sUknKnwBjNe4r
38mTXvx/lWZD6IPgs3bdX5yxVNdVbAEI3a0Q2obXmXZ08x+PiHA9Niv3JOlW9IJx
ZeO7z9iCIVX20NB0V0OBgfhmrFm/UrGjcYFzt43iR5tlAZ23+bKELbGzjbTpqK+O
kLUS+z642t8ezh8VUbOz7YeoBHPTjShw6/Y0DlO/j0QVNy6VOWUZT97wYZuMOZZn
Aks2ps8hMgzUeIQeUz913D7JhRRW4tfBkGGWOlC5a8uVv5QyonNInMISXgHvVXKK
75DdX7D/qV1Jo6QVnbTqcUwltVrk9dWpuPwHx1AjZQljIXYUqEYEbbXZzSddJH84
rettg/C5fwn8+H49RrZAqGrTUl9EY0S1u8hQOpZFzPLJejGLhxJ7JTbOzgsIgFgX
BsGkW5VtdMiAkRryYcOp1MHrBgCX7rcmN6fWfiJpbYI/kWns31DPGEQ3lE0G3TNa
4y1IGoONdUaf7Oip4hobYnXd3nruLnMlzjsFK10HjD4q41CF2tcm18b3jklvwbh1
8dLMg5+BQ/gVDx9j+sBe+moyhr1AE2WE6fFzQQl5V1huUthxIS0WQPIuAWjwMyKz
0j72+b3t8/egxxcOhkmrC+Y0dMc/TZSCxocvvYkFRK9yXUzhx4P+1nGUZQISWGuk
go/PrEeXGiU9Il242ln3Ob7gAvuOuTro1DsG2KqeQIQMnoncZwDm9/7/iC75r3iL
u7gKKmO5gaSFkjxLGCFGKgsYHdB6uiHuaHTxS4S32g4yad4Jysty5CndHy13DDK7
tbyhs6U57HVbwflj1JubutgDhGHKrVWX6JPBQLJVAVFoMZ86QZPvxok1Gi3QvnOD
sM/3H/rKvGr6YmTPJzkfTQItSJDA2R+DxAGGc6HR0ULSODVlMd6ldbEAkM14FcZV
/cdpWm8Jv8phVB/Hk0FuObomLbhwUTd2uqbeliknV00uehI2T9sBEboGMJqscB3n
j2yvDTTN+t0nooBIvjSM8dXWSLmABcy22JkCwB3YKp+FlaNZkhw6g6jHHI9dqVFD
hGLMFLjmtU8VnsOSEmB7gpjXNVJf4u/DOHMBVntIewWwFfzPPTxuB78rqd6tHKzP
SM6AHaSqQHI2JkGcgeRoBDoBMS4fNuUBtlZGpLBC+sGRodXCgfhTtlwaZLMYhRu+
pIsMesR0LdqFYCqfvTGpXZzR8c1QmJW384aagBGkdBoHamSLx9C0+zd30vK48ChI
OjuhipWjono3WAALUD66gVeHjf+dXx5gpaR3w4Y6FtrW89wWNuytbzk0I9IwNVKp
h6s3UFn/pU3oSEen4YQISGvxWcDWbsrr+xp6v7/slc4YTIxMBLC1FsZonjVhjdq/
cfPYnx9IDfQg/6gysON+S/LSwtuTuedotyW8mYlPuZj/TfTqImjLVZDq1yELfF6z
5K1uskDXpNsTT9ZGJ0g/3vJW7xthz1ac3Q8jbQ3UWGo5CdAt3jTQ9zGTbTXs9/gP
sq507Jx3Va2vicSZWuu66MB5lFVq96VIrabL0H8gA8jYxWQC94vs/wpI132hEgCN
xnv6rY92oPvH7s2i0pAy38AyLy9qDXDh7wlPZ95YhDXruYQcE4rQ+XI6tV8ieais
+HqiwRuIuADlH+O9A/u3fPvr9JlHWsGTxNAtW6aPeLyz4bh77I0iRcls18fOkLCy
qdLa3gVGssG01TVCB2efzn0+Hm8MztQa309fmzCQHZ8+7oIbnzpfMFj3YfeGhptn
eAbcxEkranRKeGEx0bXfrtYe79Bn4QFEJpG1niYKrJpqTjC1bFBGPEewxnImiZZ0
So9hUt+VTqgCOakD6OaEbK+GRafxgXJxGKeYLTvPzF/tkUZQswM5JVXYsVgdT3V9
6NK6+ZSW3OYmqjmRAJE4nTj69VF0MTGjtDf2knDY1PXI5xjFsctWfouGoGNYWTyV
QTQkiZBdDMngKv1DjpWQn5uhBURQZOJCBk4LxkaD5bhdd41LjYXnEuECxC8oaj8t
9UPF4NPYLsblIUZf1JAnkROiMTJri0sLIUAlztW3clL5vYq1lHL8hw4l/QyypFEg
bjqnM+ZFSSTRixTDuMAyLEyjvvLnEsWlledTGNwYFTmtGWDJ2QK7gFi2pr1e7/fh
K3D7D/HSWXOeY72z8nUeTNImOsoJAg/RUFT7bLvTvIV5NlNqz/r9Na8JXJAjIO26
FNrYDfnO85+NHTp2l9dQam0M4A0XIVqqB58D4Gy5+CyRDRc9Fpw36fIr6STshLtP
FTUfevQZ1y6LQuTS/R+tAUMW48i/gxvU9Q5BMUIUvY9ugFd+JHshSh4vxk5WHM/0
QeEXvhdMTDQQCEPuTyOv7GtRozy9WeUY05ihkq7wUAe3AH++tkIZcU6waSU7yPqr
02cR406072MfLCcKNaZY4/ooM9hRQybNmx2ym3FJIdu1/u/tKyF8we3RWG/r67ld
wvQROXDa3FRa8hUTSGjiEY3yXPv2A9JjwkfwQSjMzg5BntELnfv6v65hctlpIV3f
1p+Z5Ggg9TB2sR/z3F/PgLRyU97t4ZnogKuJHbZ5RQRGwD9q9vyMCES8N1w+Suj+
bO5BBzfyGu3omFyrAZjL/xxD7WFLqrKh/5wsLfmzh36FZ5qhpn8zr/kPoVot70X/
u11+ZnSfIlpQMFTtI2b3BLz/g4hJz30Vnb7JZ74EU5KbXup5lUKmWa3uQ1WaFboW
E6xD75V/nBbxFLJxGyCxc99+eCxvU/HyKsOlxjXEA7pByNTCH2pfAxrisnL1eCJw
Ssg+AuQyPY8zaWmMP+pk/GqDfYXG1nLHlAVwtdAKTKh8zclSJOMtEXc9MHsGUwht
QG0yUdQV6F7nSgnMO3+zeHz8WaH+Xi2GpleJzF4G/gqRMM5BPTUpAl5wmWUtjoHE
He0iIfZ8u/ZKSlEL9OZXMzPWa+ssa2gc7aO7fVRDKIyhlsGf8VR+Q4ugENg3Fg47
TfJw18GEETqJhIICuhPTH/wkJf2SNCrnmTDQnusRDXD2TbCosCcI7yN/c9DG3S7i
TW9Qae3vSFjrFUGjY0fGXhZhwqrgda7AqeEv+NNv5mbNCG//FnB/S1eG0z1TV6I4
1wxl4HatIFiySFSXA90CD/lRaJjRF3+FJQYXQEoabecCb3bioCtoJF8tzXzrIcWe
Vwii6tOxmkawRuCr/OHE4frU/O/n/aR1x9ctln9J25PDdqsXR/y+ymyr9zNH3gDK
q9wwHpQLwjUtG4D8YNxcaVNxdcAXMvfnoIOw/0gymd3jfm/fTqhX8GTWTPxDgxoV
N0Q8cgRgBCeZkoCiIWcZYhn+QHRT5EX3LbXWJQCMD6Fjy0+ZqGtiDsNZ/WIRbOuN
+Q+iWisvlBp6x2vYnxlO+6/s/lhxlIYbLK46lB+OBQC2I8fucXnUv9BL48taeuiQ
vygFY2jXnCceVq+3sqpHdls98mqi8Yxrb6SJ5f8aeZaBKMMmyYPatLOFHXgrJFBI
XrfZ3GCoe46cNJh/t7MsgMf7nzVhbMXvuA7hfkSzpSsNuVzYR5dxtjm0o1ywVDc4
GWotLQ5zSjwRC1It+fqrvDlZK6PO4cHADlY6yMG9LG3W/kvy0MXoq1EU++haCZDK
YKxcvSXPt5vkhmT8CGkoYMKZvTQwkM6zvotJ20zPtU2FQgMydoHH2gAzYqG3D5rR
Le11c6xYXGAkMP5z0H76W+zDlMkS0jGy6ukeepF4TsTF4qybR6+zNbQgm5yRI9vb
5wkYD/m/VeNkA1qSuMUV340gRMAVL+BHOjKtdlbUrjVd9NZLSdAIZoOTFCXD0u/2
S5fvh7q+2+wcZsvo6NAbxX+b57yDAOO8QpoQZlFcWABmb/ti4xcjRA8fT0+rNMod
t4ah0KwPJR27Ck2s/+6u0JFGLzJYFEPSlZkc6F4Jy8EhDu/ZLoeABHbi1CyaZk3f
siht2F1Ij9aQn/AbPJbjRJPQe+UCRryYzeU/btUA4Qzgv9hUo5fR3lsVUDIa0/rZ
DngQbpJ4+vH7ax8RJBMe0svSF8VTkDCryuCg1s9Jm2x29S5CVK8sKhEiivjE/06T
hiSB3/xEXcMKvqhg0JUD1evWk+UweKpAiwKkyGBVnPfh+lGtH9vJ3rEogRSSJdOa
BoOiA5xZIDsJ0bOwwukBBPGxR0tt4iRR2BQnDseyIemyzkrvuEs3rHEeuUP/KGOm
EVwtIP/ATUOWAwlC9nylHCAlZ4ukEgrH3kY5dY8vFc5VPu6g+9krncDACGjvBcuI
J7AHP/9Z808Y7iS0pBfN0RShGx6Orvz57qnuT0Y9i/Y/tJ1hlugYwNJY0BzqyUuk
JzoI66Ip0QLwEOzKHsSIFa+R169iDL9BKiRFlun5e4AuCJuyKfJ+gagjpvnvzj1l
XthXQ12sgk9se1upWLSvASIEQbgc8GiIXOGVhHsWQlm4Kf/HuwXnFxxAxkgR1gMK
dy8RkMM1X3wp+Eyy3QWsGN5YoSSOYJkJQwIPJZpg8RnYSg4XtfWBvFB7yVk6W7UV
d+qAS63BYfmbmALQvjtyRbjvltmNpKEO3RvVUzi9KetaiDDMjFETIKnxhvIKR2Tt
Gsl3lEkO+NqM9v5bkleywhvxvnuSij767DxpyIDTxbtz8YMINJ7hCacPIqeDPydd
4CLW7kCXTZ95owD9J1x220JMVaWhENLoblXSkAoXbhvCZWICih7f1z9qv8nuGsOO
O+EiWE/yXKm0xANBtesjkhXiv3kjXbgPGbnn+cK+OjWFyti45mOL4/5ARucy2uFh
56Vi0CdBcc+kP5adX7vrVoFY2GZDAcuket1AvWI+OP+fmnwo6/mz2sH9WrP4VSld
naRitn5l4gBT6MJ4D+KrwzEEW22J0qvoMjuo+O9AOAHRzPytitsEVQemqUdkU6Rj
XqyLLXnJFdj2Uy31k5HHjpesOeFO4VCWD/gdFRnHboTZKX29N2z1Lr/hOPoxsiwF
ICwnFcl2gc6WuHOCH1tUxHrOlmoyyWX02CWhURXBjZJOUAEB7VZ3mBat0NjTBZ/w
I3zX0YVdLfH48bBrPknDm98WskDRYG9T8ujPAjrtkrAifg5FcvNdXqv3fPC48n+K
ShOwJw8NnsC87RLFJs4ApaJGP+VbO8NsEwOu/FCT+k5mrjCCEuEejZP3xaQr9z1l
dKGzDUW+c510q116rabmlHWiwvvT+nXe3QWk9m5auiZSdWKTaZd/SEPChKRAIhqZ
hZMKbGgvBsP0hcEOil3lznTJtlzcOE34NEoCz84wgH7jVemfnPk9nZ1Cj6j0vUPo
0jyojwbMF2aC/oVn+rfvPh3UbQ8HjXaBsNyEgeSmlsCXtdvG6x3Ur7FHljwLrSZt
2N9i35GB/3kw8KGjDQ1WR1InHxggRRAI7gkLgZgMXX8dOliSXrskVLQoQSA5l4RU
OqvmJZX3Di+kRLjnzD+bO5aTNd5YjuFmkJxL5Uti+SuuSuFHHbQY8ESCvxM7Bz7z
JBTkzJ36yYyCxejQWn45HpTI5pnNSJXEiTp8AdZNohpLmcylzcZotFijyXyRpesF
Lax8+zZZEPv/SAs8il83xvALpAnyo/rSKqp63VgBQ+qkSC2TVSEgiTzGDcHncXdp
NBBQcdKy9Bvibpk3tesITGBVHa78exNmswT8nWBxRvzpNXwBPT5s7pH1axtSc/Ix
z5P9tGQgO1O0kOKzKiwDqqVKWTPLPMzZqWGA8f7kIgMR9aU7G/D5yPUOPh+xesic
KarbeATgkzeWgye77fuWxWQQZKEoSmmCcmdd4YP4DXMuWldsvvVioZe1yAW8kiba
QB9/gK7kU20dCnYMwI0Tk+aIgKScbIiRO3DqzETwHONedbNmzzyMBm93CTuTIU2X
CXdWAnC4hNjcdWx2eOcLgxFWtLyZXABd6Q4ZMJGvb3tqSz20XpAepaXrfl2/+xxK
sqrsmWkq+JeQRlAuKPzYv7Ev9Zp+phc/bS8e1J22J6qB4uujbkIIugHMOmBP4jE0
EPOQfTklD/fyE5PW8l3i+bMwdBpg6rGYxLA6w8Rckyw9lIWuSleCDBUnVHer/lsf
VR5uBNTsnXMN/3BQhiFOj7qoxKlbjyIBHkOqZmyTv857Y0pBI9nh71LGNO13Iz92
ot6fhgX/rCuMR9FemkJL1uEwRrI2y6hOfiV668wcD+5/P63m9YAyee5QxLq96rNh
DNS1PPxJv0l7i0DKeCCHeaKb2eYIne8nzhyoTdzhY/+gvVnY0rELhLM/uKBY4XJf
iSAXrg9dQ5iYRmouleQVcGwUVa/PxvTF5tgVc1SubCxm8iDrLYQ1xOI+3tiRyAu1
zjPA2khbA4gmEhbOZ4j2BOU0EdLwFXA8LLwvgjMw0/1AL+PeFV7TFqwK1D6JAQfR
YXzwudp6ByTUEfhdBUzTwhEabo71lZ1IDju2kiEJhLmANUUpv6JvTmhZLBQVJmBJ
LM0Ug5wu9iMHD1iEzFFf/m0UvjUUZhbdJNGWXALnS4eQUXC1Aw/BM8T4QghFb+FS
W/wMzfu1+Ynpw6MjQU9+r+3BpifXd8uiQXEiTDaf9M2AXMuJioiDYbDj+G2EVlXv
2J4qRLtv1tP++Is5rm3pUA81k1DhwQHbIyyy6f2tx+DejK9+Vp4BQSdWnLprfqQN
vf1r4epBW/v8Nm6ulotR6765SXKyL8JDuSzcAeDYM+Tfbasl+J6U69gur9ytBwlw
qTvFUs3oPQc9uqARyrXpnDRnw1wK4YO6kzjJix+mRlBN9uZBmIW2V24W1Hy3lQ/V
l1R+Z7YLiLUHH/MzYB1GeuDFpLxqMYrldnbhkNwOxEb60I/YmlDXRVip3+/rXv3d
SlMYuieLekBFUNXkzU4NFNOfalURXy4i+QeUBrM5WNhfM4KDAKhRw41B84+C4Nxw
XrAh2vOkRWJBu+zShbAVtitGHOeleAONXegBUtytoNobBbK9I5En/k5/fjTIQ3eN
8dJq/ehHwEvV7PMvtORy43uXsM56rpPH2dI6QivGJPnAt+Uxx/bosvu5z92yGkQ3
Tw5gp85l4usCfOv98XsDhtK5G5y7H4hEy/SLesj3gh4N9wYb3TIK4KrE7MjYItdS
HgBtlDkT6+Il1PMy6X259u1XU1+T04/D6JxLog+1ucvnu3fu9jfOAE8eYEGHkNZ5
6/qU3FotEQdwoAeWhYxSqmJVHijrpEna1CJXC6oDOvCRKl0hRfuU4jWowgdrJJVl
R8ZYW5p8hpFw+kW1dKpmAf1Km6Y8AmVe12XZtPjtwqNTUBnduRPpnWGmpKHjGVrl
STkgqfcfBGlfYmfvzee0CW7o44mTKHhvnlsDR+zL1emj1zzvPSf3PGvKbXiLv9N0
JXKFXFsWT/d0skTFr8phIuN3RcoqyEhrLUafYc7HezQ9TnAC4YLxH7vhGzvumpbR
R9yKCdgXqigrDEtaubGaqkVBQ7J5kUUgG94iGNoDWUQEyVZPJtRrFwShSuu4ePah
/HRLQQn0hdueTQArzF0Pi0xw/OAAuigFS3Whz8/sfRNrobm1xDrFfkCt3kmik6Kn
Pv8dgkVhBxeniNup5bjJctDLbimw6n4gksFFTB9/AG4wOQxjN+ELjWpc6AwTotT2
OFoNq/yhQrhzJfbck9xj/C6dWitrm73ngR6v98HbGxXcJcuIQUv0nVIdmbhpyHjc
nnkst9sH4h/5H68MgmDwJqob8+nJMdajG2qqbn1LbuD9RflMPTnEHYWYgZQ2z4Fi
0XQHM6aAxU+WuszAsojssu1XrAy1yciqbheG8Je3zCpCPIHJO4qUlCFwngwMPQXg
KaFLgryRDa9LERyX0IEjjGpuqaNcgqBr0W0w7a2No4mZI9/Op3GRTask0pjupLJB
eH+v01BGC8aZT19LAI8Ol827Lzi+ExScwrj2zZRALlHvFSC/Tu0sUEdX8UilPvCB
BFxivE6fG4GHl7z24vOnMrYafllmr+WJlM6mGxYmaAcxXc22IPNcZ3KDEIrCjlLu
cTJ4gRqbbXcfWR0xLmtwZDHWZ8y0M2Mo8YPTajhZaK+ApvyrPaWDH/HHXQRceir0
v0d/wxVqSuADdlZXoewwyJke9Qhbr+LmnaO8KLjTonkoiS9ejFl4gTBNCRyMgtPe
hKo8cTyi20jYY5ugVS5cwIFDSOqdEDm8RgyFltvE8XAIyLrypnR0+O42KI7uO45Q
RLGhYgXjeMLc/LWMz9SajrwwUBG+7ZX0TlDgkSFDAz4DxXuzbI8ewKLks37q0UVe
oQZsuaoAxgN21IS5hlgYGc1EODOceyBf7xF2MkVDyMK/3MGdNe99B40hDUBjvGGT
h3a3PylKs3pL2ohAVXMplphM0/ASo9r3OB9A+qK9ChwDjkRXuTI+tiIgnuQfNwPn
JLz58QeSl20rGMd5EvUsaKjl1Dlwf5NBCCXsKq70sRtb2epvAisbplhy/YaUH1Ga
qt+A1ve3sSn4sk/6Qb+WAbymabQAZSZZLEWMarguimv0pL+fKR12tQJZLkt1oBM9
JeI2x2/OetU2o+MUb6SlqeAVKJmRgwsk8n9SwpItKnFYkttKDRM4JEYdCGArTVKF
QmQIEzpgXyeWXio434ntFlUvOQhrj7Joaen3eymHATkefKKQMuTbq2vqXf1p6WfY
H87mk2QJ19G3Bv7nzwveojt99U0n2L6W89P18KAVrmGBv61YZamW7sbmLUHqpuK4
sYtwrROGqwhSdX2XXve4SHQaHH5TU1FPO+q8Lnv+BpKBqGG2D3akjRdlZfMyo/JV
vp7YLB2BbWif+NqM74ZG3J551yLjnzgjKRdPkGvI4Z8aYBNtWkC3qpYJAu23Hu4/
BHr5mJFFZQTdXY+dTwDXPsOHTRT0ljspbHJXW2LU/kVJ1TuJEgTcWL6oAW6LVUXN
pI5HtcvLIXkCmVON5zAmvlkkQ768lx1ji/LaXXkCuczG1Y/Ryrog6yEgV+DaXsWY
53ZXu8bYhRGar2KS0gpdcqQZFpZ5TLFvcUfZEjN/kEq9TgZGRLD5MqYEi88V2MuD
wTdnDBJu0mO/2dn/EwLxUdwXzsXIrTcVEzBRhLFLVQVoZeErdiIElNcpHArtXpGW
46bTudrB+I6FADsZa3oo8loZ3euMn5YG1jvvS7Lo2jxtFFkBULUFCdclKnbWpy7J
EehP6gS6+zuJHcNlpRTwUA6BsK/pYLHNXWJRfk89q4Gn4G42SIw7uvpdLIg5y3LG
3cETnlUAP6gpcsusN6mvNP1aHz6tAgDlHIzceNUqTGqk+fIX1LDXz+RXQBDW1mSu
etV6RdLPe5yLg7w2HrY/BXKre8s9dmsV0vJtBmmpUDXdilcKA63jm4eZg/yB/wHP
zyPUMTg6hexVHzim15ftYqnSK4I5x+TY3FOU3769y3ssGFlAFvlWQES3Nt7c+gIK
jwBE7D4K8zLCtS3Mlrj3ZR1uNBEDZ5dpVzHpkXJs4B2X2KwYb32U2cZfhU7y9byT
op7FJkzIEETNNKV7WvKZ2MVbue4yV5BYYebixajmPt4q48HZGPSgiquesl6KZqlf
wGUkSw5/xvquFCPk6c5rat0QBoIn+28JSdp98y9jXYp1Q6gIV8HYn5utDA2ENWgv
CFa+x8epXQ9F6VxdByFR4suoCCBMnCbzGS0UlSk6K8SuP86oLoRcoLE+NkpkPGnH
M/q68MEX34OM3dS+jsM+YRSYSGYNIJYTAR2MwPU2vD8GDqYeH/tjxiBmBFu08qh/
iO8raBXOGcC2gnxnLSb+r9JRic6l4vv9HALmJludq8fbDzbKj4tlgSsXpqUF9J11
4IUZ3fx4t1uHtcZGbSQ+2Pc9K3GTfHUUODl+QUhrnIfc9m/zCfzXPvAWlE0pMTu7
h5yRRyBdltCVm4H4t/c63NYRf7Qp6YXb50X46xPLjvDbQMvPUEgiXOaHyS3fN1Wb
1z/O7urzGrEPIdm2hq5VmQAzXF2uGoQ8X0RF2kAmq5QC7E0XUH7glHbPZiZt+lMd
YiveTRPFNyXD1+tFXkyMMwIJVBPSP3wV+cCsHcecCGl2JR1TVqaSd9rZmaHwxwQ2
gmCn7qgDLLM0oJMeTKLcVcdOCTGRyWvnOCbWaymoN8IS6rJT31Q3/msQcXi09nOL
C36FELFvtDuvcOKNl09W9zrjo9nehEtCRaO+vJs9hSt/p5QSvDuttatW5ucCaDuw
k6qrbATcqYbtdhtTiV9ClEgNNLKpFEamk4YBXBGj6r3rkbhObBHjjPoiKw8Mqrm/
e2MBKQkMNo4zMxQXKbmvtczrMlyailXaa/8zScLNizVeBgFbnW1YfQdR/SkdsF1Y
qlRjj5ypiBmb+K5zINTCEJQ6oI2naUFElj1lUg5v1l6m5jMZ2HLSh1aeK858qctu
wGzQOlsHwQEzaxigIRkb+YDEuiHjf4SVA2G9lD/xTCfuKRb/jyMbDuH0Xeiovble
X4r0PKswKGQfrkhJGgAs/4Klibk6J7su7DEZf97M3EPFOvXFaS1C0TKt8k6g0519
7WGX/j6wcu3Eg4M6F9woNN2EgXWs2k5WutdSoZAra2heePZc3NdyltzF7ROL1Vln
cf3ktZCH3IejA0euB0vEkKte6mAjaGqoklkdKyQ2od67pKQZ76wi3UT8Z8eIShBy
Zm1xj4iiq+euG60So8WBYL5wA2GvZBwhF4IiwVL2Pi+wPsX2CY8cAGgPDBFaOHeq
XNYna25JbYg14L9lgPCxla3XJu5yVJWXi/PIoPX+qPUAzt/vDF+gWSCCSoE4xIvn
ouv/LC5tqNTjf4KlCiDRGliU8PDQZx0Sc4lLv2DkPZGY6UIegkfZkRxnWpdpqYvL
/ke4S5kIiIj9CYIH71YdUX9VEuu7zTcgzVtPbN4tmz+bAGK2r+m65ln/Dxy2BFN+
wdA3HT7XmrfpMjHhTmlKbFAlarv6fM9jn9i59MugzFBF6wZdBJyCUqtLVwMQNKez
Iy2otZFgigvnnV4TZhIaH8tDejce9Wt3qQeIW6KKKuX6+f1B4Nop6Kg+r9KRShiB
sCRUOkVZTJdTygSam8PI+u5ZGHZ8PnX4kM+iHmeE9zXUifvKFBCMsrvio6mGXZ7o
r8LC8+HTp843fuuZMn3nK2RJICB0sEiYyUB7MjvTbg1/HMC5RkGIEYUOiIF5Y70Z
JzTmvZD8i4pI9eQJrvAk3/afFxdFjN55jNIp1mw47SRTD9FfYt+flFSVEUdrtCYa
cmnJmTy0Q2CgRrF+tLq88L5vIxBCtpyxZ59FNXxRfrdWXYZ+7dPe4PCicmCSPHx+
KVPnXzV2pJ7Jk4vyL8I86Nxr/maiJoV8k5qKpInbZgpAF3J8naqtCj3HPIs7r9gt
mjPxuEicmFeEPIatPWFxuFonb3AfzeJjQf0vzBTDW4//aiFz2PwlrhQAiuNmPLTI
MCQNVBqMOIbPBwrdFcZubBsCTptw9kGgVSBtZ1F5UT0V5qxW7TV+ZlqejUUfBisX
wGGH8qa9dI5dZr/ikbemoW98ue3gh4ZfXnoEpM4JfqxpiuXumaDs5TFw4wbcr+fH
xdOv8U9P71DIYNXkyF49ZmvQJKuhb7xaGa8LGMdFFJV6OPenXu5KiyT6bwO+m4Ja
66k6E0NT4tlHb8GE7NKy72FknTHQGXFuiJKeK3IBZSqSp28NawYWMV05n6GJFF9t
2pt5Rp0U7JgByZ1ZG/LxR3Ck7IwobU1pVMT+rEys8MY6LtVEe6F+mS/ujJvK5Pz0
XTH95z7p+7aVJmnDc0NcFEyQhJnhhxGHGtEi/oFwixv9d5PLO9V6wJKPipek7FEl
6SYrCB8sDVUSj85MHl2M3LI0wE72qTJjNyya9iG9/Apbp7k6+yXgfRlgOhHoOupZ
aENwrDJQ9gC+Wi1CxVUsFxXF1GG28XrVRitybyOq8j7G2LJav1zetTdIlAMOWDUN
gjYvqAz99mGchLJvisktb7ib71VbiLm9K0uKDyTjdIGsrFY63az4pDBTGuXKJGCX
P37HLuSxVCHkuoqoYKMHN/lY+T2yl5J2/N+Rxf5NxTvwrlPXd/D0TUxEvCEjIspi
ip+WxLwpBpYDyGzzgZKk+BM0kpvLprLikrl7GHws9VRoFBNzp6lLlR/wqfmk/L1Y
iAR1B4926IIqAQ+Sk2Q/hYF06kBSJu6MoIOga7zqn6EAanbVBYVEu/27Ux7uyMCI
8K6AniEWBuKje1ol+LzSynr3y/9N7D5GAzHtRRNk2vkVHPeFK/GZmglW99cN/lg0
oGYJdB8l5MOEQOyXnfl58TPj2zGlo4VTnPAAn1VM1vNZGWEwjqtWM3gdwug8j9e3
3XmazSKrTApwUpSCQeRDtxGLBWNCsvPZVLF/8f9Rj5zFdWnMuAo83+Xu8TMeG+jW
oB6a7iDWBkB8INb2gBOMXZrRn1OIECLBaccsspjmGXBTm7IlhmtRVsjTumlTmGFJ
gR1XCe4FLGq0gfZRS3JQcF9SRw8m88yg7upyr5ket9RQImio0mR+rlF+qR0uBMSx
kchtNjYZ1l4LtvPRV4IpSzZdSLNGIRDcZZjcM20O6IKTSuP/SsrDdBDweUJsqMwi
HiYJOCiny1evTQu5fd/FnnYu/MJxqrKuQzKkk2tXlM/7iNVIZa49LBkyBnEWCxq9
lEl7cuH+FsA9ikaYjoQ+pXQGwBjen1skFhY9inHKGgO/wCm8NgrnNf5BHh0nv20Q
16sUrmRAssvmHfzsGeWYC0eiKupE3b1SiIrLZEujNoOeNm1P3rKivhTNOjAJnEgP
hXsR18dJZbCYAUa1a1VNv1UwjrvrxBjqa8xwPFGRNw+KYyW1kllWr/RAhw2yMkbd
bTYENfQT78Sdgy6yPg0UokgFgcj/a34U5y7aKDZti28GWMy6BpROX2SEf8eKNUhD
BTzIuLqfI4n2vbCALE3cbwxnKuAnff5iNwLz2KdKOZFXtF20VRbKwQiuk6jvJL4o
iZ+UU35xeAo/TCW840N/vyvwC5i+Ab7P5Ez5NLYPHzOY1AMyOoCrmcQQKlTT0YrG
OQtGJOD6f6ff5hDV6bMzMbhXfKgBuQ3MPvoFjUwPcIXqO3/7kU5Ekq1Zzncs4vg2
ZvvjP/5dk3iAL70LYYvNqjUKDuI0HmqbYdze7aj2AqKTD3SiYSdDxbVeKBDTPlDo
yRGHs6RMr7Bkkh7T92YFfL42pM4LXoLPqL1dpIHeiIKg/FaftT+zmDdirfhmbYkL
KKofSqL8wlix/Qn8cosgAhnExmlOf9Y6ooiZ4u863kbfNY+wx/pTzxn+VAbnqbOJ
nG4Sv91xoVg2xj1cmzzFh//uYlWXBz89OoTJEkixptAPrHBRMmOjSrtpJ3bRR4MY
bnEmi98D4LR2rRwhxDkvcQHMJuirVsswxaYif5U87Q6/ktpdCJshWyQyUkhYSNz3
c942GuBMy4McFTmRO3Osx3MPdYO8mBlK61D8oJ53Gmy+JYgr2GmpxTcSdJOE3cmI
kLBPaxNrRvy8F1ZFdV2ap/yRYENBVQVafFYNdf+jJkAR5B4uKwQ8AxTwGiamLhsc
9H2f2pot7wEauugUTrJBtroq9kPino9rsh1o4QyiEtagKBOFhdkLugy82S9KrcsO
KhqvBUZJ83zEj1/Yy3rgBLuxveJhvkXmZiN9Cc9iDVhn7e3YbRlF+nOxeDwZslvq
//y3N2nRFRoKpQzZyCu18TSagTbciq+HtAohddJdpQyUNG/tZ8JsYjxVPUUprZFA
xhYWNsUAWs3+uQqYzq7n9dq2PbOJpyRQlkN1u9pkT6z/syfTr+yFUd85DoK0LfG3
ScxNu+DV0pPvVdytmlKkHzKpPKs4g24JsZ8yC/aZV1pS5yJRUVte0F0Z5Ac8lK97
fcyPDJVCPoxA4hyBsZWeQ51iLymb4dwGpmoHI8ZKnpZQ+u7k65fsNFdBMrMxOjFs
aEcM9GBNV/vzMLMadg6c8OSgMDqpw1kkVzDynLecU8NwC6c6vNI3WNTwkPDyG7C0
kbMt5LQJcX2Rg9nhw3RJEMClOayQsVbDwi0cQCyLZwG1MVnWX20AXLWMGdEjCR2p
Cp1yO+AeAXmcaHbtmhFiDudHBq1wy3c4KHloo3jNcU1jrQvSwLuW9f8XiPwE0fqe
U/GzdiqGNfM1uFuUVBBqODG3W9P5eJ68hfhHcIqxLbnTVGF5rELKLomePoLPZkdq
UEPPBRbUiQEYqT9jLJ2XApSjMVDodEaid76+Y7Z2C0r1BL3SJVx0IGM7mU9ceYQM
j/JNUZvBCTUnbMlM6mjn1ERuQ991vZMzeNDM05ufp7NJWA0ges3Ye+j6LNmIV3Ud
Bg1YgIHPQUw/FQFY0zw+SgmAjKBUawSp+5gpHL8Jl0R98i+yX+T7FJX59DA9ZyHU
LFYhs8gnXdoQUssw1r13K3iniAVlivFbHWL61Ac7ruQhs7JTQkgpGsIsvO4ZmSuD
PaYH/67KhpSawTzaUaDmLV7QJFKiewc0sz6r51vHA8MwuodwwX3BVcZaLk6xfpBk
AIqSu6wMJRbNQU1on8zU1tOQANBiZAzvIjfE6wGYIf4FUwxl5HOch5voHOLY7aSf
imNf+vqIu45F5uyoWpg5NaCTk+jmUjG13nM/nlGGfHIATHF62sOe2sH8ePSFl2ky
1Wl0JvA3qWye1sjTuAQWfQYQCkhzWzfKMeRP5Ev2WVXvvCcQsBdJkP6p/s1zuRgP
TZCPXwKNE3TQs6DKPpvl/wT7F5fCgilnFX6VFPQK+wnwFmskOMTZw03ebHUH+WFh
9uxq/Mzk9dRiW66mDNBqHTzFfY472WnINXyI0XzU3tZ/hKno79nhNEEM6Bmmxf5T
Tu3MJqED2bUWuiRzMSnYy6iJsnnMPb6slmcbD89nUqENn54ip0WzWrJcXphaFEnm
PtCWB6xd3rG7sHxy23ZDsACYPcCKx9S+abznvhiMU+OBh+OHnQCLEmbKBnq985FM
2pZT1YBrYuEBB8jdrNp7yflfN/fIZBfdSHaDNZLz6Ox4etaW/6BXWqMrSxXLE2es
N2UcT3X71B29SD8+Wdlfrn8aKe7C9itcWfcSw7iXNSPimQgZPcd3iAGpqCrL8w+L
acriB9j6oPry7s7rG7GgYe6LHT6WXL4TnsI8sqrpFl9swp3y4ZWg4D71fUzx0Mca
gdOhk6KT7Xr8ADRnFp+BK60KZLR3oP4V0RSszI8P2fUDZj9i9q9BvmQaFvZ6V3KZ
DYC8EiQ5b/TzW1ZupUTuyrsYb8T9II8xWOVwM6gEqBgxSJu7E/FC+bazfIoiWmtP
xZBMGhCeOwkyHwdJqSoLHHZODykuYJmnA+QtoQ+ukymtIQWYtXW38iw6+PyDgfFU
JG435OqTvJt/NDXSCN1ypWaOoTdCyeAQnFvvTDQbTK/Xe3swFCCveJ/k5mjSZY61
5vE5oLAs3yCXBURMdDISZ3+4hmn6MPUAnbjnMqcs5QlxHSrz7llCES/9N+mqrr8k
XPePAxCwCqka35XDaBiGK+nZb8TwMHuS9w67UmJlMGyXsGQ+6GxxzAKmlLEtug1R
7E5sWjGM+Unvf+LkgvhI/htFVU1ZZ96InzAcsHVMEtDGWL3ShO/a9+PeQOF1VHyf
09jzqyx3QZpF9FUTNk3GOZNdRoHElmf93+H05Bqo7g+bE15CsSijjxzVz7A7dWzr
ewMQkpMFmes7MtGQplULPrMTmRgqPHkcz1N/8txFYYeiqiwZqBcICHOO06cZekST
eHpiKLjux5Qf+WMHddgoPojHGUTs6ka30gbt1KmiRgzLz1LNZZ1PiEo67mr63K0F
WmMrmPQZHbEmaxf8g8AMZW+WUEHVhWd4+okwlgFTN7yUQz4Dg6y/Ni5RNUYHMZFk
Gwnjac7/26/5EaamxWmAtjPwF3pkm5nmkXD27uvRDtFD9AP/mtAdgaQ4kayiVGxJ
DqGwUjOD+/u7/5j6CiBH6KoUmRO5gicpoGJlfoimBYUZEUL02HQ2xCcxyPgcW6RE
+Lfi6zuhBKkztCVpReAGkRMTnyl6ks3Xsi2H96pi7a/FZyHvn7eVpOvE9VwOa6hx
1GeKEqol3daudLiyYKfYCm/D4wkRK73zTiJxGo8ZdYjqE4j4cO9ZwdIhimfDGPdI
jEQIeYOBaiE7E0+Ts7me8HA4QUL9B5xpQlpVSDrg9iAVGwJLcdZMKVz4jZmX2l+W
n1MJVvrbqgwSSdH8YpKlVRxL8ur2SBs6WHLQKa/8ssbbz+40mwY32WnmFmyvtdUp
RyD2CAIr8wK4EoHCgHApWYexLQXGYGAkr+k4NukEfOkdwKdlj21Kg2l9xk5he9xD
Eoj0BSBrhOYRGFT+RbZ70JVJk8DoBY97o85/+80C++bRVwiBX17NY1ng0TG5pfrD
kuhdvBW+waHjATeJzXKSLG3amCb3uiI0veWK75x/474R0/2yx++oR6gUhxPYSXSZ
3oeNIehOll1skvxZdY2FzxwJjH/eFZbiN70HS3wUcEGyzDZb3938wcxHAFEU9oEk
ZG2W0Tt3jj7IexjB1INGL8/ZCYDUNiaedYk/Dz9I6mMn3BNiXjknwRL+skKVoCXv
v+laBEsGPLvYS/c0Bp7MJtdlhvAiAJKQj+ekTYGImi2bCrRUJFUJvNVioCegnY42
TdZsmthsVxQfGmytlJcS+kCFyUnCoAMly9f7WqB2tFc9hu02eC3HQbeYQXvj4LM9
wX11nnujexJ65YH1D3B3TXwEErhHPuiXwj+LfU3+DPYmR+Dot8BxWyfOeaLbWfgf
rTneUD90T2pNhqkaOHWybi0fFWdR2tD/Nvtfv3l2JkeZyrQygRUaMIzOq3iU+75B
Hua8Ctx8lpRa0qxPGgaYa/fr3PzGsePqOEmUi/myTd4T+E9lPekxJEu0Ud3ToSeF
IueSZ1qFcmRxENEy+ySAQQhCPp9APnB+UMp2/ixjVomXpZbVDXGwCqtI0S8Id6OE
Brck7e0r7mq1A7F5H1qtHTJq3Li+Tdv++Mz+xzxlB+/s1My7wM1KRiVfnRzRl8Dk
NmHlgYRNKnWhQGU8Du2wy6iphwqaa1okodcgCPuucvXB6NDS3RxfJWDP4a0PxlBH
/NOcGwV9qtQW800FhB8CIjEQceFLoo4UOO8fwiALz+x9Dxjtp8eqRywr3t0/PMJg
onynmVYkjjdPwPnArGz3N5JjijL7HHVS8M59q3FXJF4MxwNZtki+AOxtMTA0GQYX
UywKNnIwA7DT1n+VV2ywg5HVVkTV5H5YayYnhK++hGcfpR1Id0t1TxH+XjT75Ehu
DAMZLFN70QaWHqreRZbix6+K1/icStrLlyz2kT/XgSSNLOXIqXDWR4s4eapP2g3c
CPUM8ijp40wyhZmBRszMGhEiKuJWFftngUErd2NpVxVrODQDT9I/JL2tfESE+6ho
+JdSWH5zOKhrLm7W8Y9tgTV4XnMKPl5i20QOelBoidKm5DbFiBstiFEtL9DRNiVH
49qFnSTpXkl6IjNmRM79QnCVYsTopIKFmUjSfAxy9iYTsrjLcz3oZj+R6GLecFUr
/14tfqrd/Q6CZf8mylXKf2GKaJfr0v0S9RV39fb++1KIwcLDw6cj4hzkpi1qTxXm
3kECKLYiEwFp8AXAVrsIknm0lDuu2x8drbeyvFVNnI0PjHeeAH/sscZyS3gfSgjW
kYTMeUfTC3x3Agf0Edn9t7GwgG/gqzp4YvTXfUkOjZTZiQ+mFuvQxW8TUUt5ZBTB
oYWu8mOlARfwnjhZWbBWquF+rYGxQXlwFKeQJH77v9sEkgJKxCq+L4dctiw009Me
IPyfPN3IW1LLqZ9ldZvR8PgjjENhqIWalU7QwZaDRriQcSyj5H2k+/ApWDJjEB5E
xQo3/CPdtbY6LSzm27N0hC6PhfdV+NPwRXbPOxBHeXCO2e9abwcZsP0fsVyzyhhe
CVur5MFpMI+kpd309quauFctLszXe0tbzJklAUGp5JUYXwcJV77BnKKsyJAbAzvp
Q05dFFC5aJ0Vh2Vpl1AZbn3s9HCEawx+q/ADGXJ8+NbWU1Xwx1THIkz/ToL0JnNz
WtKge9EcikCHfNZE4tKHhaE6O353iVnbcPwafExXyjj+YRvyyRrKuVlimHyR7lIV
hUzGNg48pbcQRCEEpfYTOe3E4N/WzdhdYjNiLKbDLOGMloydsNtldtAxsKREawCV
L7aIvdpf9rerTXnVPg1h2oXXrlqpTcg8LrQOmItD+VdH4M/HhwI5sp2KAgBT3Hht
zl3frLCLMbwZirUl2Vx9Hg5myatmnVa9e7tkq4f+u5h9ab9ZmvCK4FAgGzZp070Q
P67TeO/LGo3O5W16fzC3ckvGADfJL1XVKdsHQYSheHwfG8aT1QFqwSbVDUc84fL/
J9DnfDbz4DhzFZhVaPYG/WGtmYTo/DLktfSg/44z8NLdwnrDMl1WpZy6gOLngysX
ObV2frs0R9iLMeENJeIozhygnA1u34jbRpQHsDkfQvW2NSACJ4HTo/XusgcGmxPj
iwRbvbgWYOdAXcQaoSsLhSHiQeiSpUJhNb5wjQ3XRcghgrFKZSx75ESvig2yB0xv
QjSR7N2uMeVjyr6AiSRm7wFL6w/toKaAc2ncFwKE4gEYjMLJkg9XuAN+I8XlteF4
7HbCNOB/qI9Qj828uec9lDMUP41iA3t+3lY6GpigQfh1xl5G5RiFZgJ9CUicm1Xy
6JwY4W/YI7rtmPOLXi2ZkWU12ZxaLQ3SMwJXWeKEuHXfEp8PyeT8xNbFkDPGYeI0
v8FARxWOnEpdBc/jcw+UG+QFAaPLSLvPXOPc0elCvs2inqTyzGVtOx21AdpgUQv/
QrpR3xXsqHfX5OPspzYiXnnpQfteJe3dMovLmkPj2OWic4Go69f19IXPsCVM36fM
flu48ZVghy5Bj4UVc4myUaStNWogGGjObwEHgX/FWEAwCtZnEApr2rz1sm++1TcV
2DE93KB8AE8zC0SoRm1BCRqEPEYI/n+BgHY5YdFmmD2jyy7lcPm6hd2ga3KlRDs5
AYhl9CPHS1w40ewabvarFaSaiaPoncnJG5XHRWi6v4hfWSHY1yBrmJJ/zK/smODW
FprfJh27Lkn+/+1Ol3FHiN9LmsAZnQE9M++4ZNopoBxpHUzhzE863NF9SEdZW9Jk
qdFsg8Y/S76psEArfgHbxCP+j1nn8ZgyUnTPD2MA1/O91BXpZ3rxt2bEfgjux2/c
3JcyVQs6w4WAYaVc+g/p6OM317Mq0vfIkVngsZkRkr6AQOqpKvsZZ9tP+m0xTgtI
Hp9klcp68UEV4ZUkLOxKY5w9ojQCG8BLk/H9zk+SE59QXMBPXNTXC6bLKIpkA4wO
R7mmTYbAuLIMTML4VvV6LuXjpbBa0B9zHCl7IkU1H+UnhUUHOLvPASE6SORcat/Y
cWlXQ+aVYGjZjcPzjBXjanAUMYxJUZfcnZAHcLSd/dhN0vSUOio4Wmr76eilNRMp
Ds9WXHG/YxYuZfjyCylPN4PYpd3pY/ZpV5Ri/W5gbyYgCycAXpqvEwg4mv+bT/gu
oPzhoJYUNkWQu99P5ZDwtUu+FXssD9VNgepFvu7xtcidWX1PW0hH/7TEgO7wWSQL
ximWrqaEvFtbXZLIwjBa7QcWjfcKIIMiJDOZScpWNj7ekpKUkPXAeC02qonILG+f
FXE1zSd4Q4LQP6XHgUd1rk1dlsMOgo6nLN0bDW2EA3nPsni/Yom1X/VA/UdH/9Td
uc7v3yGEe4LR6b9dWo8p5DrCtvbBIBpf7Pv/ROvKHDjkNG91zSLcqlwzaXKhzz31
KHegPNsCa+KqxEm5tnUq4WNCtArCQxfeuKkcnKERgOoUgl4LwH4s9Ju5EWlHYjc6
gHx1Wa9SXUwYkvBbDX/GiA5FDQpzoIQzkwR/ORZTuZ+MMZ4Ji04Cs4rBaHILiZZY
nz0bPWCSulQvnefdZ0TLi8nm9mpqK7iiMPuZ9BizXZThZVnN4S5/JsnDJHJ70HWM
KSzfac9D0Jgz4Q9LuLdeM7yTwYZe26LDkdLUYCepKobFlgVsIU+fR8/paU/FDPU1
a8j5QtU5HXG2MK3VpucRrRo+OJ2ePmsgNYdAtOLHLIPk8GU1+GYgLp1F6f0Be1Io
evoSB1UzGpTzRD6IAlShGd5kyTg7ee3+GksaQ/cF18Ca1cR4PoYktNCYE9P31FNb
MjdnrvMBZ0+X2Y5G0nBSjuC+GJdwNcExQ+SRsMhehjn9yi2bhoqQe/aygWsphdeG
sJLeILV1ypqoGht9lHgWenvgSc1gshy8D8qZC3Al0MGqhmn7bchLK9Pjk2r/IxEh
bxymSG46wSNN3/XXY5FvmL+/OAyqYliUv8Jqy7C6/BJYAXBUOBIQLmcjOPI9QLNA
l23sTQacDg935Zn6GqxbLW5gEcCIblTXlCemjmh6BgA5806TsQopfYllu0u/ALJT
0bjgeFBTTImwa2a1RuXTWdgyyQ6AiCSFp97JUyA3EVhhhdio/WOEbr/fwoW7FrmI
2X165QVoOJxHkyy43DyPkFnxx8dOzs1FkKA8CfS/GE8iXazDcF5kN3y/IHN9iEtV
mpFWnJMYMr07ey6e6wqPX+TU5DSyZ09WLIBXxdorXi+lXh0O/jldwgBITE9pz9ho
gN78qtzthUO6R+AsvnjvwXlxIimdxucBRtCY7v+IMFojBLvUb8kcdaxKmyWDnhgt
CFkNag03Tkpw629EYevjptiu5NYlQokkk8YrSwRTK3BOzj3rzf4GbMBnDX6nSSUv
351PdgcPMhQMaVkQ7QR3zaYDJESY5FbMhSFT0cJiOXtoH0GyfesEwtQULh6CFvtJ
Ycn+KLpBgjWs+9UsJmeq4Qv2DwOnexCF1x4jMRAajpiqtZd5tflhoHuGr/o8QrAD
za8XMplJmuGaG2H2ba6qz964Rnf5g94y9ZxtJHibmVh8GLSUjuf8lHCMOP1Bnoc+
UgfEA4euES/n7ql7qidsl5+fiO19lR0SOy6cVTbORwJzuIeIYL97aznPjYZmCE24
iKWolZvIj3uzSkNBA2fZ1g2GPed+FxXEyWjNZrf4hc07m+0mcUJTLpijyF87JycQ
Erg+bipE6ysSypfyOTT/3f7yxL9Mke1EcYd4W+kSDobgT36KoTX1eEYLqR1Umu4F
laVPnDRWESmuPfrgaVwhK+YJTE7RjdPigbt9uC42qre2a4n4mnBQsm+4CTH3vCEN
g9SuPsfbMBUOm9ZhlxgCOhJBZkgPTJKu8WcO00P8JgQI9NLhQ+Y/sQ0bGvCasqEN
lsi9ENeRdDOkcVCyOri9Io83QNrqi+W1h/onmVELBo6BvvK1/7ytv9pRxMbGELnd
wLZJG1bUdq7xBfrOrMKrEk0Ig60ely5Lv315QVLYoEjuqhUux0QOs/xALCicD3Qx
19iHB8Od8qhOBFEeo4Bkdw3OSieUstkVtCxpNaw/c78UWFG4XL6p9qIScjoXdq1O
DsM4N/5T9UYDVjO6TMU/Pxh0YbsrxX2hMIaIqvOO3MTcb/X7iocagFu9XpCC76LM
qBVMeEIZ/u/ro/gewOyLl1wUaoyAfYqROY3jV/Woi6KNVjXM4BRmCltYpjJd0r/g
0D0Uclt4uEpLHDzVFMl3TvoT59BXuiiM5gIAZUyQNprYSB+6V0YKHcTjljNrwkUN
Q0lLJnBtrLGmrc5kLwBpu36NbGyphEkplxXX2cS+w02yqXk/xClSsl4FUq4L27oU
daDDSCBTpnB/tRIP5vRRlu2VAK2+hk1nec3OCK5RKBO15rNiCcliFzGCXDMOK4Mh
D+nwPPH/OKFHu/c0Emo66A+LaQ4jZ/tM3oipzLDnQMxvsMfVbmB9nixCRiAqwV8u
4GNl6zW89DLnZQAYxOa3Wz0axXe6PU2TXDdblFl5Sx9RkXwBys8Xdel18WSPMfcN
2gvAiPl1a3GW/DQ32xrVKJH1YMod1HaOVHb6+F5kV102rKcI15mwZ9f+LFKitlO2
BIqG4BQ7MbFmDYRps1ZkgsTJ+OXNnBD++7xYQ+/XhA1cosGqPbHuLb15Dau5Ibur
S/GgCeURCnrFnYU9qWh1ZrTuM3h8oOBVQ1OuvELRyK7p+E1NRaWaUnlJgrsNrOjj
mkdanI4FAopbfkDLFY6qtkPDAddUeW/3Ecqowd+G03eNOVvP3Jc/sfrOMu/+CHQv
88EjQt6SA+HMe9UHofNl9Zov/YQ2o5jP9E3NESWJNIWfqeQ2DmYLHZJ4WPIjgPNj
FWBMENhxUsXWWOTlXaeKSpFGJkZDy+6uwkHqDg8lvpEx/HwVghChHgXvGOelkt5o
HHcIxfcJOqIH53jNKYxiKnN5C0sH2XQPQDIPvcsYz0Lozst/5/EokrvDZA+0KNOf
iJsswp9ulhDgja4QpeIzFoAj0ReambYl3O1XDPV2nLlLQ5Cp/6ywwx+5iJAVn9OL
sgflwI/NaSpZPzjPHvyY155ukz30lkWgY3H2Y7y3sAsekIMbMx7qe3+C0H4ZqcEs
tzgw2ivpKxOFEGpGUWvUKROL7MK/psEgv9i/FwUWPG2icj7FKizaO+wSrthvGfD9
sk+4qff9C46DdgLkQcwN7dliBqVL/rD0ALWe+EUkW7T4dny6GRiarGiUvkPIwBx8
OgjN16fZz9GNcP/sPObJyVyZRCZbVYpOFwZ0JJE5Jc1sqQYvf/KSvRckR0+hrGhQ
AyYeTuXQhSmJwHW/P3WHR5MgXULsrj57cZi7+WnBY0OofvTg/YQp1V9sCom6Mi7O
C6qQrLA2n2VzfBNwleF9AvgvE3684dfUekClBndYpSEO9Hd6CSU0Wd7SU9XRli7i
SsVhP3PqPpLPJqJ7SPJk5I3aIfPLkX4DTzEUQD7/ORH929WD7gXi4oHAs96/+iEw
oi0aFJXybgvcqPew06onrr09T5ctiKjxLVhUkzsPXGLawIQ90en7W0p9balCuRmu
9uT1iRBcWVQU5pmWziXmz3NT+844PJGdiARLrr4vbObLVxVBSJ+J8W6DzqiaYAcr
TODAE6AeuJfnrbyFGTBOzR0Cnxnjuxcs/opAOQOohQpvMS4RF9Bpqe5DFCNjlk0D
a9nRvmrNPmWKqDxhadV+yP7HKWHrV6y2lMJtqMmtVi2AVE3wFKmF1FwItgHxVjw9
Fy3xsZbKKzVtctEn/VTzYjm0/mN99aIQLfI4TQrPTmQrngqe6yrzQFsqoWC7ae2q
sTNjR5NL6Ba4XsmKGtbApDw7JVfWvCTrKaCLlb9AghteAUlG9ZkxB1WmxaRtcLmU
9+I5pcul/FgFtk8pJXjQQKgA9lr3++CTBG8Htbq51+/BRGA809nTtBPjN7u5NEjY
7rpIYigfif15CD/aF3Qovud4cp16H5REXiZhqLjUby9iuoktdSOWy/0Mr0ophpqo
uetL/rwoXtLMF8MaK+cnyEz8sT9Nkn7AM24JXL4ntZXHzfDoOkhTT4s+tfArx5c7
YBqACuctIMmnHz6WiT0GEgPk/KDWXe9Vx78+ZXFLPoXuX3Wkjt+ZAwGUE9m8eBUh
pAh3SuQbKOkRyu2k+k5/DTqD8TB2Hfmog0i5A2YsiBc/aiKCR1TMcULCHjdDcqhQ
2PkqAoVtCvJrkwoOWgjOP+Y4xBrTQyG2Kr5baeldEvJ1QOX/cj32R+lwS9M3tuOE
d858Q3jkudnutGy0xIGdTHsZMDMe0l+OAw2j+QkxTmW1ri0+J1EVgnIUl1G0zCYm
tduimWNH7cCLwyFNz9AnJ0FheUUIerpBecdIT2d1OtGffcPGd3xAD8fI/52Re0Go
HPZOqW+fy4QHv1jUmTP7KM6C7eKSYM4rskc6euW9f2AwG9Ojs558zmD7Z2NiBVUD
neXG+Y+BySDVsCHBW8yt3gvoBWhFErISAWvLnOal3P/ESF56O6yjAkF6umPNVfDg
0YazEbm44MtatpciicNjltvAeS5fZ7hphNPJUKA3YU9xB/bb0cExmhl5nCS6SMs7
1jX9VcrWARm5CJVz7qgKCljP0OBh9iTjKinGq4mBlQORn1yhSVQkqQD2wf0zRtXM
uNdtClj4gF3D3+BGdwfDyzx6K/rdmlaKR8dtQoRGp3nGA4JnbOnCPZt466fieECY
1BPgS69YooGumdpq2pg/13bhsYjhAq3OFdb06rdIBHUgyopvqjxo4puCOrjyq0nN
85da0ajSSPaBDBKQmHV7lPq5aF69kX9WMYlI3JZUo2poyXlbOEXbeolAtHbX9Nzf
0juko3Bfgy8FxBhCCHsPh3U87gtlZOCGyeM2lIWN9/x/nj3Dt5zvIXafzgtoLXnJ
awWdZW4iKX7wBbrCBr5atTPiWBUGpuHo9ncry9rEHmH4c5PkfOA7MIH3iNnvw9eB
x4uFmoQomVeUyirmpbOLa6ziUt3vsDsPV9b/Y1yL6AQ2KSOlSAnZM7cSmG35BZ0/
mSAftfO1DWSyIg/uWoEs3fpRPlfluEqYyouQDRABPOAxY7uSTx1lSrmyejd3KiuG
7gXLAy/ovCCcJnUOShOO3dQB2+RKjXqi0buN7atMAbznQv5RdYDhsZP4aFOEuOuZ
mf2FNJGWL+HK3Qo2Y+XDUIP9Sd30qAiHwzbh1AIdtTThd+MacRSVu0le19wJBGYU
Dw8Bu4M9tDnRb43h30TIEYRMTE0jiXpqF0B/0GJNr+mnUsPvhrss7+ujWrL6BIG3
5eGGQZvpsYY3ayx9vwMCuE+7mR5khZpU9ELqh90w4mFuh5tGAFtluvaH8ZSHC59h
iRFXfaNL1MvbC0NtAJfG+K37g8AEWREvibn05+fKCagBUtcl+QtGawFH8ioVExrY
uPXJpNNjv/H4mn05zVTOmugzQltIIXECJGsb8gzkXJLI4CiyJI8b/rDVq0v9XPfn
YXyI4uLBHq5+0FmBIzyBrOsRDXj2nFskLFbM0qN9JG//5UTsGuO3WLXi+FiTU9qT
d/dm8Y96GIh9qptw3tvYl5Z/0Ny7/brUnnq691cvpqzBDNE+P2l8dOBJeK9NcXDb
iBlbB1gwknQlbgbu4q57VWu9iO9HbVCO394fw+Xebf9V7K/ZHjXbuj8a7ZbzWHUe
jKei3QFEDTgSkQXN/5Gpah66slTxQ6Sx/ROXkUQS+yVmzfE7Os7jJ2Mv7xkp7e4z
rgMPRBebQ3Sfz+3vsVoyF9K0+8QXk0hk7lf+jAF1ZgEVZRLYW6xLerET/AH2d5XU
b/lI6Phta476gcnHN7rRM0EOLCJSAaMY0rMalObkXvRk0INByScSYJbJe4iXXOej
YjR7m9GeSxSjGxRSMXpL6JBt9Uy+I7NflThcgBCCjSLkz1wDpKBssmud93kCB9Fx
/GSN9wmGMRVhInCR710/x1NPW2IWTUhq3c/ee5xR0d9ZNkOLruK5DB9SqXh1J2P+
d5T8m1Qe6HA6gZE525B94NG2v7ObhUhg3s6Zp5FeAmrlbO8SxV8HYeuLZvqTOuqn
BksLbpQ8IPhpQHCVRPnWFVYe62rgPxXEpEEGhjrx5MBrcVSyA7IwVU+zBL7ZG6YO
3b9DgB3+UyfnAOL9JW7hvjbLA+Y/wUnE1qGC+DoEe4yMB3LTmpHyI4mTar+LM3Tk
u9i/OCzmQsVlhZ6rKCLzruc9+xDPVzeTD/P0PNe709O2idCyF2DxuLid+AAo8gnY
pBFgMtyWypbxy0yqRhHiH9BdoW9Xpcmkq18SkDgmrgAt39yb2qvsnlmX+Isxnj40
FjxjLeXhCh1Scz3Tce3Kt4bvymkeUVypiiiFBsii/w/JKeY2bokiSEWYVpxG/2R4
SeEFi83CJk7xPoq760cSjtIsuAlKQ6NJJLOapWkpWrNdqVTrLR3/HvECe/CVb0uD
AYVmweKqpxmax+j05ITfmwz56hXQBDVZSWi3VNVDmPaDbdKYjIC3qLUfH+KNs6TG
AMaQwgWYa5WZ2OLKH/2JNCcFQq+OM3dLRSWUsoczHqUnm2MdFNJ+7rBDOum47iy6
3yYkVh2l70gxkZnpvAONBhmS7lpUQVmple94WZfSH0KEFM6T4FxbzBt3qgUywJTu
8qKOc8mFqaU17mPtK5owMb57Ou1u6UsqGVLrGZRhHY/SXnGvn5uoE0Xe7GDnK+F3
3kezQJy6oXHtft594cOqISDhKbMDPgD/zkKdNxku54l0kvH3bhp0LxN7b3W9AeBm
ZC5+kl42EcLSk9kcoD9k3QFefQouWjsY8ibDfAWdwDB/lLqnrn5c4knEFsumEvqj
AtlO+idwv0H4ZW9l+n7hUAdEgwTEEcnXQUQHcYqS28AAZoRUwhx3mk2wOJJILxtx
G2uXVK92u8+o+zeSFApmg4mwmjR6Q3OqFWYuzdgCvgZzUdOcGYHHUS4zKI/3wYrX
aDqsXLn8AQX9k39R3bAG8vwV0uBdTRCmFMczZQ0/E0SMtYMA3J0RywoP4Li6BW9m
Wo6JqmYGV7UOMhbJ9uiT3a5IKiyxM6/89vfg6lwJ9z2zvHfSxc4g4AfFWQYPzGR8
V/yuSMNvNkV/ECZwWGNPjFZnn/h38M9AC4e+v1FMrS8+d5wkTRCGejCqk8UQsV4N
G5za9eJeyhUPDr/RfUDOZsfRJTx5Uc8F0H4X7ztmbCMWV7b3M+OuY+2aex2cMTg+
H0ewN22gc3HMCPDOqgMN8hSaCVdHOVo2qbfpRLrecNIYKXl4XqqylRti2wo0wc9b
4y4rz9iqm16wH7/KRMFWQpWu/aPvlrdLw34dvTwKrPRmXFShhGewm9AGED7Sa74R
ZdoyegoATZHq4lCBQQjcBhXRl7pgQocGGdlfFRie4K9fPwtVelH/LroiJ5884K9U
PQTWETWlhowlGx2oX3eQ4vZcZ5BG2EcKNbuSac3DHChDNuqyzcoVC90GaWVal1AV
sqQP2+FEUc8py4ACjP5+KvrMSekrfIvmq7RHMkIMpZuoKxqgA0YHxSUep1K8VEhK
lD89lOHYbG9CnbzksXHWnjL/CADUcGtqaGSgVaoGTOWo3QtPrnnA2xO71aQ8kRcp
3Hra3QlnYzTuLG6D0OZKD6vk0vX33FP/ae9vCAAaouyQGNOloLI9RwDzhNysYHhk
OZCR4/Ws+QV1IRjjfENSph6p+T4Abfv/tMvj7tVSYAd8PvL8ux5ws4lG0fLf+bKP
ec9rs0ngVcd5PSr+Uy6O33G+bSikDD7lk3dmiD5WCKciVyMX1cMmyy7W/tFoy+/7
RCaVeptujX4K9WiudOVSXTW0oe9/CXOLX+QGtnzQujG56XIIjvOI+3RR6WNRlY6s
QBJPYN+FZWkBoFHmhGoNA1/7IMxCrmSBZgwfmNvZSH9aF7cTA0+ftZ7Q+blD/Uj9
VcnvyTdf0mXyrDjmn6VZQLbpPCEo7PNCSDOB6arfojxze5O+rAvPG9OOselAbNOb
vkmX3ItF07q3D2fRsSQQV/cCaRAbN6AYsVviKg9mLk/Kd0SONqwAA593eK6K8dK5
hCOYBo+iZpzXJOhbA+qXv6SQ3CpTgwTF7V9qSJNM5mBgLVI85/+6yrsEFfi5czro
nZ6AGQRVgVEuoHswYM3dwp6nb2OgQ2zVvummqlG38F7lDwV2hBJHbHcpdLGDaXdl
MkVNS0MVfPbANuIEAv1UVVX2ZIxunm/BNe1grKqRkhbZUfWynVsD+yrs1EE+OVia
Yb/95YS1XnRgEl959x5wFf5BtMg6sk2U1a/jjRhrgoSuc4Cz3/DNOdkFhvJ85gYb
1rUKyUvFRTdHEUj5ScxP3VGqa1auCk+aC+3jVUc91ZPPBr8ahl/AU6qEYxdO8huz
XyUJrS7PGNCqL8bPShzKoHsyXIE2IA7+v/wsyCBQ9AfW35E0mq7Obv+mzDKNjv1T
nNu4L7oOKYrGhcbi2PNi5cFOf85yxg9KWJ7I4AHfAGvuS2pgRawOZ5l/2b+QXjiy
y6662bLxLnjF6ztE/9gTGGlnqZSgvg/cBThO5UBvSbQn/U1kVEOe3e6XFCgQ1ufa
9cKV3xI/gU5ap8kZfAafR6pl89+BjX4o0RBhob5l+6VgUTintTSux6zo+qOLZfnM
kyiqXQxT3MqQVJZ5OR5wZ/VaULn1AVWqmJ1oqXKCM9kUAIWopjXl3lD44jH61xhz
3mJzSuKIR0++xQ973grYPa++XgGVCsy27iV8Tg7gKkvx9TlVAGXe/toJR37MpJYU
KIuvI7lq0KOgeDQ6SUR/a8fEJeFI5YLVEeNeve3Pxcf0MuGMWjxdRP3b+NAK9wJo
1/vt64tsqzQjryHHQBBb5FM3GjzSipvl++GA7+x2PGbOY5necImUdXjttbYOea62
KtUSytd/+ioIEwcnleIoGRcHgb0N2xPLJgDb2omHg6AMYJDVIyePcxOGETsGyEvF
Uk5nVup3D8wDNKoq3wCeJXDra3mUtgqOsal+GPG5HBeEHdIx4OCENI2YmaJx3+Pn
PB9dHDiKNlvhn57Ppm9804ED/Kbp7COFL9V8zAiWpKQbrI8NbhcEBNCaq4Ua+xqH
VIZq2m+ux+qymMr9T/sWVVSmedP2x0Nu7l3lv9fm6XEKYI3srbhhjNNoG9UAVAeJ
IFB2eAUZdD18D9ZofaBs9lZ6z9NRW+PWyY9LIQt4M5h2KVGJDZQoXFC17719CeCP
fJpDka3GUQFdULkWCF36191q1b4ffhO33ncVAXn27bgtlvZ7SPOZIBDTLKg1fD+Q
Ug7pfKtpO9Yi5pnBAWDxlhvLdScoIg8zHpNmO4OMhk4ShVQh5BDI7g5ukC/IoRP2
JffcVPMCO6sSRdm0ZdNEpDJxfbc0+hJlgir4F9ZT00HuFQFV+7M7+NCGXqGQWmsj
2BBAOZavFbRFWdl7VG3NMLeC+KEfP9JPpso7ep9wMRja+rmMyfgZcK93I0MyX/0b
vRcyB6MWZYBHdSr7c+F7eqnG42q5OP7emhQGfwTiQ7t1HsnsyvEEtCB6sKeW9CPD
nWyhZ8xAU39Fu+1cYCyp545w5iXhxbYhG9pae+IeJCqhQVtPJPQxyufcfVzgmmEH
tUUfWdEl5VVlb39jciYGSjnF4PbyjUpHuAIOtEQmNquiYhf0nleP8hMgiYSwsrdI
LqXzv/0MJ1jkrgAvx/9n32NN6sKait5tZLwqX9+BEs8WzkRFKWJcoiGLT8XWWWxS
j5rrezh5A8F+g/YA/x3xdZK7d+YQJG0svi7tjklvcxb6K+y2FoIWne77/P6tIAZE
f3TBRf8kdrwPQXF73yqttdm0hePvkMgeD7qfFtXwQ6jDNGlWHelabFmqi4QMbeuo
QmrD1SFNse1NEW3oSFphevI60tULHT+Xwypwk3aYk/bNNWQlGIlCG5z2jeBWrtVL
KGJNUK8dF2YC+V1QyfgChpvf39+0oXPwYDquWOUwBiMj7e8GeegMq7kBHNwTkZim
8G4P3zDraIioS4WV/UanP2Mia36kJ1a6udqiqRs8O0ZAcKI9oMA9O++1WtXqixOe
/SF0ZYFXClqs5ZmbOl/j7bqfGS03Fo99s321UXyyIyOPzLhSxuvdTWThduJhMaO9
agbQvY3mISV78dEEU/8UaAUxHn5PmaOAjYZlvFwy23DwbzKCm1nK0N4T6e2LDS+F
fxHdOtuyEqdCBAC6lVHHjP/KlgFaC4LDM5FdUMnV1nbP6QqOO1e/oPXv0GAG7QqD
499pQ3vpEB2ZGtOZGMhHmeIgu8cWzWIKETrwI24uEoMCYHLAHNMYoJIrHkkfPYC4
nf/JaG5Bbv++P5ZhBAcnHninWazj4Vv/Fqp933Cocg07u7Ldnr3/IpFuhYQizROn
f/Oli8abam+VbWCStlRo8BJ2Z75DvYJGNebund7y+M2BjCiFyXiTA1Rwy8CK6hV0
LsteGkI7vcbUsUMg+PAmTnyerxpUEfWTZjPTbmdpNMwdXblz68+pTHTF0Fo5ud/4
MGv6S8AzkzcZA5MpZad1QrHWWAi3cDCBvBYh/OHgnSCJeD0TboITMpqGKp1Z64fE
Gpsgz7S8gTyiMqMUQJwdcDgRt1CFLjmhRgct6hRKxvw0SW/0vZySgWT3vl5ZjCHw
GAl3H0g31pvjGDxTW9RrT8qxxHZXYcEQfJAC9cjv3Dn32oq3//okkmVIMkp1Kp69
RurRGe/dlxQleFLj8HK2M8vAqCJBSo7LNzrTMjPNLrnkHsqAnPSCHpFLOc0x22dT
HilpXKSKGRN2B+82trsjku7SBEZZbKLEr06wsQ/R/yMY63jVTcGrBF3ZMsoPl5AW
x4kgx/CJaSuq2zPMBM4uiHNPX1yPigtTyvWPV1Ir8e0HRWUfVrtT3OiG3rkq9xVk
WGxROcigT7q2kcnzV9QDMuJSRztRIBfmJqXJF90enE48yh56Nw45pv+wudWNk2yd
fefpUwyHeRtEmp8DedcMtK18LAK62FbSBXclj1/9eWwgIjgdVcVJ5SVIEOg+ML+V
pS2JJBF+ay3fuhxlecjO5S9Tg+SBnTlR5zmTbq+3KUW0Orc5F+CVUrEQ7GiwRrRE
sXjx7e7fJQu9CbLBS34bZOmaDl459ePB5cGoMBzuOl9fkZtZaGbZNo6XnYdOmsMf
ClLxR+r5WnyK89IxbbNYUsr+mBljVE1Vb1Bk/pXdaUTIU4UstVkmtpUBqIfZgvv6
c6zIIKgUVTW6Rhl33NXBf+j+rUeHRTxDa/uHb4xtQRlv9BK1nyp1GPVxrwN1mbOi
yx6xZiNF8c9Ore0tu+aXREDRGN85vpdxNzGi6lDD967YOgvAe1UsyHFeYef+mWqI
MLiN2pxouZrDlcbFlGLNwQtMZY3It7pzAcsZe4HcDHIWEjFPjFu/6EtavwzQQgag
TlVrwSvsegJMt/qbJKxdAfi5kDvZQ1bHy7AZBkTnaRdrPdePDxiXJMCo6SbAea3X
cbLQgUM3AvQ+I5EJgvXWX/SmzFQ+o2JxAF+zO7Njfa7uVpu06bhTygiOm/iGaHxQ
m5oUPxP+AcIulgyhL1Dy0zUxQL3WAvbD259k9maFsgFT66ce9nEym8k43W/KpT1Q
lssHxIm6GhvU2tDwCOtDFDeEY9jRFbSYmtZDWqA4Xuhw6uzZAab7iq0W+r6dgFTD
g0qSMyIb/0PwYBag7yv3An/ZH9CDUH+Snp8Siyy5qyWNFA3srnKr6CQRlBRU/QEz
9PHPScLy9MnM2gDzMRnKwFQxo8ANxt8BRcbCZw6rpA+NyVJYGO9k05RG+PDXOzTH
3s2vDFS5FCqVSA3yYSUbXlaYz/Zrs367X36SDFPA7MU3xye9oQqxKhr/LxRHOgQa
Gq2dAWOp/q3mSge5E4/hpqJvM7qP9cJyt3XRmyYVdE+frshU+nbPE3rXGnyMYR5X
6Zz12mjliJ5KHYJfTuRYgg5GJEwZfvgyPWWZqZTZBMIOrC0+1ACJ3HGynZiY2iL4
yEEeALMHeiTdD9/LtZMznRvmrQSwQseaAL2gI9CWe87YeziiGvZYpl2iBsoMWlIP
9edyNj9raBmEG4LPAGCdzqvXyqKsb8LGYj6bST21CjHZtnQ4CQPGjAKNgZr2Vk6v
Nj+7XiNAbioYBRjeL5tLIeXnxkeAxFGaBQfUYn6DsmjvxuaMvh66fs0uIH05nD8C
8273mKaRiEIPc0EZHTd4/PHOHF46gmamfNlNV+TRaqznj04k+azAB8QURlnHO1KX
EarbCTfemn5dZOlW00PyT7+ZCtJu3l/0040BY4cE1mL6wAoD5eK3QxnFjGkKditi
PDKgMH9LNNrcECnjWN9nKiqJNht1NMu430x0GWSk1Fn6hqQ5O6k2mWltOkkxtqr9
yvkg4GDtwLzYoXqqU4YClVizi18DyVvKApcX/Q6BCvHmQ4e2J7IhM0D5u1Xiw063
OtOLK8j/oZtn5V1iwqVTnhsJjYi1Av/fQZVuC4r/cf7viLoZb2io+ejA1eok2iKV
gFqzSznmIMADlTljzpbP7rDPPHbyLbRBGJxwv3/IHwweIBtvVqJxyrnvNNKutg4n
dp7KUJ0lFgJ/cA9qXw3fvPZmzfTfglpiaq60JsVXD2g5iwENZJgEWR6cmcN1xxkY
91ScRr0CNeVaoW++Ik4rETccf288Z0bhwz4WwLIJFfpwOXsy5OSI5vsHVO5HkoLt
56YM9E3B09ecKN0fOcB8LGS11GTawDeeejqloWnKYGlzyViYfQjDK3+rAPW6wNp/
QRlxv5a6P1wgZiXztDLv8XFkYa4ulRvKgFtWPO1azyNXjF6c/N9gV2J2miU2qIYD
VZ5UXTEej75w1urf5DI2gQzbPJFlJxL7OcjYpmpS2NEbs0KP61Evs6tsyW31OgD3
5IoI9I1jTe0/c6hG/SZurpCVZKoTQ8FdhKxAL2Yok6WcekoYO0QxlS8NMK6VuKCe
xnLn+0DiTAThGmMc7479YU76oWPAO3OeEoFU9txY18/oxUIsgc4d0qBL5x087idG
J4Tu2H7t8RHdOtsHZQ56a83tIVQuHv0GdT8U/KByIHahWc/AaEqsNlx8kNi5fYAn
K6WQCXM8ZdBsHG2qV9urXPfUKRJVkUYZWreBED6ZX7rUq87netlZOZ2kWODKsSZ/
Eg8UYe/P3QcjCH7zkxt5C0UVIaQzzlqpc/X6FmsHsf1KwUKU66koDZex2Jvc064N
KfJd3sF9mjc1GfeWcky9lKIWihNoCnpyjef+KRU3z/l1H0zbWtTPkhqmvvK3VfLu
+Q/HZpBbqbDhu8FYKtLKTDcXygAMXvXn1Yiz0C7r8pUSBCEd3XboeuNxIScESTd+
8UiU+Blq8uJ6MtqBWXvbSUNcbiBDm8EgBXGagTNRn+PFnrflUD29lv1pqDTw+9mO
5JwFazbNfouBeR/ZD5s3KFBHASYhMRfXI8o7XZJx6rwmKAJgBWvTi/e6SZpwHTHC
H1ZQIuhO6A10Dsx1MpyBE3D/1Om/MBkLI6SQ86nmAOy+Dfd7esG0Wg4/3gsNCqtu
mY4T5NKPPx43c/o7MO+bmqTKbfTT/jvJLLhlKDvpsJsm5K4ZKWgUe5+jAJUOekbm
Ftc0rEmxSEpBqU00XW40J5qcgAvG5aIkQam5bCe5qaE2/ScUJn/GQhfP53IuWDB9
sIID3Zasf/fQjcR2jMCiuBAoSbJQRQoIZym1rF+QeZo7cUNtyvlW9/9HEMYKg4eY
9VEKb60Urv1kUD6+azo6y5KGB4TusN40k3nQrzYmOtD7HwqTnqVCD0xGHWzn6BEn
TDzyaSqwpurn2GXUIz/InArsqETIK7fbSsJXxVi6g9jf8sYnr4/0jb4bIZyqFJTv
BneT8L6myGpwgFcWJeqE4OYeqTDH0/ZXt7/cI/zvlhp8XIJKSiFPtKWjNwX3/1Hp
bALILAp8QEUPmalOj5/xsg4yl7btrGhbWn9z74iehH6ULF2cjfyqS1qJNWtB2wpX
eWJJHVcJnA5Tf1CUz52Uk0EXRvQqEy56K6QmVEcTZhz6/VXw5wNlN6vv4z+PbGur
xlRUtJ93Vp51LGNr/OVoxKqS2guIdMZbyktqVWj0zz6/8Bh/x0JP4xmxgzYwPEqx
0EvES8ylWbOFTTfTYJcqK8ENngzm6+PNuJbVtnKLZcWK5wyVrHHJ2mV2sE9sOWsC
lCYNUjgdBGUpfpJ484sOE6dKLy5WbCdji1lfzfpK1lWiFiMnwlboYxLovNzaCJ3H
8Lgc114kbWsf3yJjPWTR4b2VKYqof5njtiLkZkvKBGH1irdBFuav0xCDzxwk0FK/
+8JvcgTpQ1QNHd2RFfsbBOKDb3ro7WceZnm3OzUal2xp1OTYCLQJT9UM568da5Ok
HvOCbElOaMJJljxkaVNuUnV5OA44WcHZ7T4+IlXZzKETApUbePxI1ukZA2Dyjw/6
PFGGe/fAADPCh+9LwqiTIEhCfUymcOEl3/7RHu0q9TuQb6Y9Lombjd5m7k7DQ20E
F/5q7y/v2+eHmLiuy50KRBHkA+0GlWKZdqK987NjfFkhMiK4zaDjDUnNAos80di8
5L5zv40XFWfqKerGL4RZ9iReYyoGeujWyHl13iwkm74h0XLDrzGhrRFQ+GyMIExW
usbwyeddkB0pkrMt7DRgnb4NIcZtGBRyjfBPtRH/oQVeCRVTk700q+OxKbhdoq0t
A34gCtmJdU4emaki7cgJ29fMMgoS0Md8j5eJaUifYf0YACiTjzBTqcSe7Km63uTq
TvimWeRa215UXnKGYqWsc15F+XgIhOLXTZKPeOh9p3gNyvD+9Kk9WArTWF90eDxh
3wM6o//lLRd1pnn1YtudLoNCK38tmiWpOzE5kaQRgxN2sBnQWC1B6SiZAk9lBeal
q3bnNU3HxbU5ZyIjj75FTgDBRxfCa44Exwjs5sRHhRc/ccXEb6f3ZAXppj9FGhgS
/uYAR/3tXUIcB9ueW6rKIs5vyouLzRJvfuEiWuViDAZoLxpTtyIcBZMLg8dW0esQ
5RB2b/K55znxiAYNUASSfAHPIQALqw8nhCQy0ZBQiB39rQQz2lhOkXTkm1RIjCAL
Dyr9ysaFOTpQ1IiJcMfdRQrx2F8lhvj/a3CvkpaoEU4oL7KaqqOQ2Yki/laO4ImF
cLAuVn2xnAaytJrNePavXFeLPpAIwZMneoehb19j1Tr4T/P3Exlety4cJFYobjwf
y1V1FQT/2DJO/Ud3GeMv5jPMaMhaC3XLoLIhx9Y2CmZNADW27zwxPsgEsRt9/aYz
ESjVbX2ueJy41vZKSa1Gl/E6IIAZfjzdaLPy/dTG+D/lrvVLJ/I4OliBm5nxvKiq
tj+gjhVYzeSRPLjjy7vxBic0HRfGEIyyS5qSO9TU5C+A3sSDf0oOfiU4bxW1Rpnb
V1FgOMqD73HAdNC7X8B+9gFDVWT6VI7t40EcfGI1rysXg2xuJWfX+tMlVgyUfabM
5svIVBI92tOlkg2SZMn9gF0PNOyO1i+Gr8HIGHpHmgaAcNhowSyyPSfiRb17VRKk
I0TwWicUo9KKEZPUs3kK7JzqaeChXO3EubttvxidHV/p377mbzLKxy5unrOcBpf4
3T+OsNYoXl1J43wCgCJEuEcpAxxRgrv53vG3Ni4Lsxn/tf72YnGQPxIvvidQ9iF9
o3WQGK09H2uSC/LLOTbT/czY6wDYw4VE7H5Cs/vj/rf8TM9dImPy8wrV/qeeDZ/2
KfVGgM+//TURTqxyfLjJW/uXPZFi2UrH050J2Rq0HhPV2GlmeDoagpsiTa5nLziy
m3U5Or4xxOjCBi3z27259ajVOL7V3P7j1/MmQzaMOcvhjl7H12jNPYuaY3LU91UG
2lirZ1cWOEsmxEyqvmDBUxgY055gZGePRlkEb/pfY+gZwmAddnksLpQLuJyYbNlg
XAs+pNAuSVo7adlgP6fyO2qpMhJzFcClx4eUIn6C/ukCBHbJ3n/kySc+9AmYEhfi
PLO39Ap7IxV7801irZ2zIrggHU+Iab1rz07mr8H5LDWofyeI9ANzdTeyHKYq+ymZ
KoJpGMkX2OAhPDUeJE2T10f4E0UJ1okou4P5xx95xHUPC3b6fbLJMdJt9iLUbqt2
BiNKgImQtdiuJRifsnlbnKsTTnh/V8DBjKSc0cEDWxbElK8/TwXDN4is2mi2Fpdv
51T+bvAh54z5YSSwfumCRyytXIrUkj94hNCKQgXcK2cHtPPCg2QwfNltTFzoKzhu
4L9oraLDSwc2D2fptQHgfNCIlwdW9+uwXuxloSuSwaWqQ7dwuQ7Ab+IRtDWKGwKC
CXcLUko8Urw03nM6LoYe1iTpI+fcsetqdzFl/+POoB/3E/npRmDbGlJJJeKKRx6f
mcSWpXX0ER3GeFgW1u/H287WJEOR0KYd9ntmkcN0BG165jO3QxW3CUchKal1PKkV
cJDPwlISZCVyASB66dxNsLUqkHZkMZvPFVdhBEm5nymrp1XQrc2gy1LdjwWuypsV
W1nNcC+/WnZ/IPK8v2zlvbfdDcKKdF88oDSqjHRxk+UBhnx5bi2oDZf/8kitx0J1
JfZHEqgXc6leoVCmQGVy8Ho/2SZzdMp0gw3A9TlOsxpBPTrBgjRQk2d2dD3mVPE6
VkKCOL1T5CqlzyS3jChgP90e3pm6sqwW+SK2+pxkWGssrAxbcZB7SDsy+bSu5THQ
MWpbKavtG03GtBidDsSUeQsTEPU9twdYNhqa/gpC/mKtdRf9e2T6s13prUBHhq79
WKfhfthjxI+jZFFlVf28+gD1QoHqQBvS08YMNyzV/SKItLLoEdfzXP0i9Jsb3jfn
5DvkMxU0by0DUia4I4bmbuuUyR5V2uVP3kabOwEqR+vrr4zoZbt+4BmTb4RZEJkE
IdNPk5GJzDEzpgKJ5N9TCq9vOrqBWOloDhPTxEiSKSAyAqXLa7n/D5AhcLtsQL4d
xstM/IXuAa0XXYnXJE1JxV1LfmHSl3JnwPLpSGFq8Rzk+nO5oPq04usoeCTcJfxB
UBRD9bCIaHRXNy7aiRsRDqMtH4Mytrrg8MFlqIhu2aNP5arGOMeUBJC21j7VXH6U
QRid8uULn8wpe4ljiu2hr17ZokcHKFhtZ8Kl6inuIzKJd9lquLIflSQ6D4g8CxZ3
ZiascQKeSVgYfZ9knaedk+IE4fYtYCpevcjImBLD+cGb6m7VFt0b1dLvBLLEBEMk
TrbW32hoj2sSIbtc3rBTqQFyl0bhoUc2dms3tBAafrgHl+6xFQzvtrT/uStmiX/R
pi1vGzr5edYpyPcHL7dLVfhJyk960hEUgJa3WnE4WaLMIGm759RvKCP0KXJBreFU
OK7DNr1iT6xGw9QAByGvgz8r5VxaU52D6NOM5sgdn9A5IoZGBEJGD0Z+FOBL2Z+B
JcMBF3MWYVkJo5cGtD/s02f9WzVJPM1uOHlJ+d/9FTnDmOPcjxdQcfGkkMPExLfO
KvfGqp6M0pWEOhBbR5mumeUS3kpA4nFmHrN2W82YMjjJ9YuRj55f76dbh8wQz+Yt
gwP8WJf8jd+rhw95+v1NjLoEfipRmthsUPzCtThofXo6u2yNv+mwHvWKWA78BUug
Vz2o7fX3rU7axt0k4ws5HiWL8xHwN2acZg8fC7PTvOgCWfY1zq9G3ZN8LPiRUWbc
1t3lJwGDMUndpK5L8jOyRZdW4CiYDZZblWEbhss5zkWEJeVFJDImRCYqdIZai0zO
IZhvESSkfU+YKRkeNN1gq6fdr71GlM0vVndmAPnW3vxvp1V2rCBXtDSz5RtoKcjh
PuMSwPM0PC+gcIKlzRqLJS/p/OYE3xLjRP48TFlwKE5G+u6UAAe8Q6ZSWztqWcCj
u6z8GOjb26JNpQsaXy/62T+G6vD1c0S09Ni8IkxQtWh8E0SDu8HCcSVXRQIHW6LJ
bAMu8XoHFnG9fPONwr/oUdwkRcgkGDEkX68wfnT2dHzJe11KymHDC57PsmuMGvjA
I0YGmzxeedpAMk3y5KiZgscobAjoYfibGqkvIKhUDHqbMPJW2/lx592NFHgvGM38
R/gGmueb+kV6E66pRjrsr8EvOt3aTeaE8OiL+h4l9U3ZWuTT8rUkUe6pIrwF+dWZ
8OgSnpWdh5blNaei74AkJhSrmiuoB0CIdhkEB8mBSXSGIzjsvRQX/necnRSuJhgN
/rSkqXFyKQWzkVnSIo5G/WY/erhgwMkDE+KFAjBpzGQB0fOzxdKic5KRNxTFye9b
ipqBDP6Sjz6fhkkGZxZUU+telR/6GgWcVDLDbadwbs8ROw3hb52LwzJNHq2pj9X/
HYVslcFSRQYgdqkPyKH3cHUi2e8QlJidlE2Sg0j7JO4eVe1VPXjo3W8GGKEowpNG
lCJQ6PGOPY0d6/POZSpYit5AxG0oC2KEYID81ZfYrDI0RD7WnYWmvabxkze+onNf
apF9Obab+d/p/3kCY3bX8u5Q1njZsvK2JrSQC6rLHqiBpeYZYRtN3OkfnATi3y9w
mjWFqFoGrQTTLrVy1M+Sf17WAecEKxttl4FLx8tCcXknwYuZ7+Ri/4/2jHMJtVsw
kH26QU/zZpIC/wOBULK0pyTRpLdgnnYsBNRTCQEPoioIus0JYdLgtBXZaDl+Dgdi
v3eYOkxpIizziwcj5GwYlYMZETLgcLmWr8we1Rqlmft/oD0KarA2+YWTtQtFu5on
cl9vLBcvQNtexzU3GXrifUAotxex+2bXekqk5il0bMmPvlhM3dSc8u3A7rvCe0fx
sBdmAmkDelavnlbh9fYS1EHEwEu9BYagNJAOjl8mLQkAEULkMX+JdNpRLxbJMMy1
tE6zkPr5TSVCE9LY1D86ypP8DqigR7Vq+WDU0Pk7SOP4ynxXbgOZWIA7X+2F14Yo
ZD67F/JfGh6j8soF//MgTaTHlLszeb8yTcE6TAEJm7pCQfJ2cEmf3Bb9SEZ1BTsp
ImC4Ha9MDpRAm16WchLaXJNquTXFL7Qux2f2LYoFew7s6wXytE6Wq0eHSrlH90kg
1IGqHAOghyHBhRuzVZwhmssMUvK//bYJCgJUCzVLBaR1Kd6qaQigv4F9hcVtppzW
0UAi2WT569ifBYMpmm44affBT/M4P0s2a5LkM0GOxOpm6UATD/l1e9MQZCo/J4F4
dsJAfMcoebJ6zJCIMmnhr/743iPsqVGGd6EZJVR9Km4Qnl7V/wTuO4VL7Jocr0yY
JE9z40GmBTLm2jqDrNhzDN7rO12fsuYCfMaoOy0F4vp+0zSO4+smttJcng+62AJy
ggTmQ1yRrtLWEvF30lePUKK2kiMYrbQr9qwarB1D64EaGEWXd7p0glHkIWTL2k6u
12EumGVDZ3KxFQkMrDwdl43RNkF8mif/5NuePs6J5AbkxEFXrfFubS5IrMz1wcXi
wFvRGsA44JkqTNs5Ul8LYB10Q43M9vDDqERQ9pXmq2O8XkZrmoZRckXWT0GJ+Ifr
eH5e5X94KEirtbFnXUtoYWhl195zv+j23NgzaPpSQiYTDqcBJCPL9ncty/Twg3i7
pZGix1MCNk8fUiqQ6j1lzjBgMnkvitpx6bVDCf6vbdbzMp5yjLC2nRcfZZwsiyIT
vLWtbHHDEaptaQBMv10ZX5AL33bayFnAs02SBxYAq8ANb8vUSEG51O5uJQKWOSQa
zJ8ROgqT9VsNMX4/cdisIFQ53adWxgmedE+qQcfiUGAnS+rCp+f41qs1/PldJMUZ
CNLgYcelQi/bZst7HLE1O/rezZgl3IW//ji22Rjgf1BxD/aaamSm4gzD7pc21vC9
zf1vwDhtHUTMIRaCQOPxg2lv6t06+LN/p067O11djnQjucKnFUsvkQqZId96LPYv
UsDbLp+oyZWIgs7WeSeUsk5MrnDpPemPo7WVb4GlV4xuBt8QFL1YSraaxVpU73rz
nosx8B5Sb/rg/32eXyzcNFqRXnQOR9Z+yrh85je3Cy6hGsdNhgPkKE+N/uNpKvIs
5LcHgxi9bw92NY6bf70SlG2BxTJu+HCf8qSkloo37X277YzKzsm05eaI+rqnTA6v
g4PyKJhid0VcKEbhF21PcIxrGCnJ0ko8JPdAKdMYo0b+AoYqwUglvrK6q2IR1oPa
GyI+grH4n33yZg8luqgGhlhtwJW0AKoUrSlwJo0CMHdVJWpLpV7yrsiHv5T/6e98
0l9cR6Oqe0eP44qvFtBQLo4LbTm/x7ojw+24sgL1oE2bCr1FKh/hG5ljUbyDd387
LrTgH1YsbwrYjUFDclyA4ds4uT1jE+NvYEcoWifqoKDx5YqNkZ9zhK2W8xFLrxzh
MkfeE/VF+jBLmKpJY+o63K3uxFrEFsvIGjq9nH4CPy6aipRYkPvVdyymPZRAD0m0
1BQLTr+HYeoOqTXFFxT8e675rHl3L81lUtIt4bk9g276GykEc6aMGH75FeCDAODO
T8sNF3zB9epG6iroKmdiDWR0Jnz2ORJeSBAmWzcICeXkvyH/aMM5z7A0IW8zXGu2
LIuD6FdPqFnpcJo5DZMsO0tvqJDLKbgDQFI2FadO2EiDuyDBLw31WsXBXU1WmB1W
2hWIylLUJ9YOGx4ton2cHBzGbzMIhu6TUcXxG0Kv1AmSe4SEZ90k8clp0KZiW9s6
BBt1PZn9RVDaO8Ivm7ijTra+bbNIOSz/SzIV9K3KV9DuhUEJ+v6kOllo7p+lXQ7n
YVlykzHj/l+0KtPDlz4o4bNeUruK28y7CNaKs2/znEVnYYCk+tPB34412pk9/Tcd
HbFRynFJzqoNH7lKQVA4CGok6aR1rxXAHtCrEko5BO5jc/KZpwRGMAWIReQocUIt
y5Gbes0Sa24vuWPWrXk+yaoQW8ACc7poLml6OS52v2e3GI1z4lL4SSTdtwDH+jNU
/f5/XuQWhIaaieI9uswVTk3iGQcqWjgAxRKXlqHbE9Ddt/tpHLSYw49Zmt28/0Po
6J44e85vVvAnSAOID3NBkTm5/0ACz3XF4Zt6OOSiumMM8zxMO/GqaSe7PVCM+uap
q4syVEiJHDQL0LQVYvU9NT/J7ZSS1SBm3RS1TTnaLzNOxcvbAPHJbM/cyF3etHtp
ogVtqCTLqmxhQeVuRT0rG/lL8xNCqEtAOK0D+qSn8uYr8cFOjwiH+0B7wV1fe8AX
8oEoGFfaKICnE1qEsGUD5NrwXYvrhsJS9an2jP4g2OsScpBOn6DGRmHt6Lgv/NA/
3kv3+2hBSDI2hw7rsRf/A0FaAoicriFRNPHiMkktD548YVda0tdnyykVt0Bt2GmP
vj4aHdh6hGz1M93uq2gXCQCmInq5R685UcVA/folgx9xdPLKK4rjyAN19R0W9JVo
0R/gy35iZqUzhGsc5LHWHttHu5IyhK983w9+FvSyY003Mntyq1sZZbctDQPccOso
fe8//En9R9zmKNYwFbsRSjF2xq6tMZHhpxARmh+tPbOSx1lDdvcYc2k4wEHObOol
7yLhSI6DkQG9bjCWc2wSv2jy+rp90hglsMdMVwYbP41WblZgl28tbwgGUJmb+T8h
Tquj25ray0R8gsDOhPPq6DjtfAlo4xMROtW2AHoy2GdbgYWv8/ptllTl6xeKaVZh
czLapSaWY3rvzPcr2V0I3ZXSZguWmkhACdXTB7xMoUY=
`pragma protect end_protected
