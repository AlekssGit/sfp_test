// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
23zYYfWHagjSGFIiprSnT97CcMZV+6NwUYIFRgeb++6meDaHzWkE3UfpoMvwfAHp
KSWog0W28AxP14BqzSkGBf0yfw8vrNX0cCrwcxkm+jyZXfwOFYLT7qT0X49HHLa4
lpEBhNIBQG/eOap7S5xmxYk3Nzczd1i/0AvlOm0Le3q7aaG1n1xAug==
//pragma protect end_key_block
//pragma protect digest_block
KGSW+0TQ7KoaiGc233X8XoeIQ8A=
//pragma protect end_digest_block
//pragma protect data_block
nR6G/NjlrykKEiseiiQq7TKreVVcU2NT4dber0tqMW1omY6Sn86qKmZT7XccDMnn
F1RvGdo0HxVg+yWbGbvXh3enYQRAlVXP2f5tJehN6Aos2anzPC5bnpWl7z5ZJPgd
/aP95LTb8MdLYptfGUdZibrYmf8taAeeSzOMBKOxA39TnHcmDdm4xGoQIfb8eAG6
eTPs5TbeYJLkRJ9cDA1BKdG8jBi0EZWMuNE/z/Q6Ztjhi4cXw0eoJZvU0e6PoXo3
37SVf5KnWKecMpBmNpZHYvGnvuhN5QXbGUXg6n0XK6IDZguDHcUVySOquW1XSTDU
kLary/9CfxZqtNKSewxLbnUFXElNCt5BCnE4YuCrzLoHntEa7AfBEfIu6wKBNd0h
Nm5UpA28MF82KMUXKnr+U+s1f8v8DZUr4sI/2Ab5VrrVB/TERow8z/i1CX/duMvy
BWFTaG9dCN8UpSXq0QzMZ9pWObVQ1wVmYLNALl1YwIKV/1yZzt+oNW4/AIzCYb+2
sdv/BLluhFrUbR2zQZIpIhPKmeS3iwQ9b/vzoMuc6fIzlIkjjUVNvcaHB8oQgsD7
i+gsouAILaH1NV7MWdOaDeGO3AOr5W+lyXNikTNuYetadttiiBpGyjvpmWPqSYgo
RoxiJTjElFnRh4n78zaRwKvX9tKm19RhYJ7s/lfzPVJtTIQ+wAsHrsMPqQJ/cbzs
F/3mRz2UQBkIwRXp0MGafN28dWFRcfDk9LKUIwR8epfT7cTTuMPdjJ7YCl4Im6TD
c9/UEaz2XI6GmKjw0pYN2ZAqXSYMi1zFIXiI5gajp/8Em1+Va6TDW3UVKITA2AiT
aCjZfOuwzOWfXRenmVo6fgj36KDIDP0f2scKek3vvKHtVQ+UnklOwulcDT9jB5R6
5k3lN5jbBvzXQqAMJ4oklfiTOXIvK6PHgsZUUEEbk3x74k+uj23I0pgdEsv4SiJc
7IXkhLoloTMlP/GpoYqtvquRz9ALu0xyJk6acH/34APSiyd4a8fblb3Y1hL0/wP5
TD856MClF4HcMTt1CK3uve+bbv/gLl46jjFPxvVRgb1dLSYHCZ3RrrGoi9u56fL0
Uq1w4uz7z45M/L/LBU2q7/1xqV334nDGDudz4qmOHAGlLBs4XapUcNp+TB/xXV5A
O97xKhz6K/BzgJT9ROSR4MbO9L5lT5+8Wm1GWi/D+GLX6IVUesda0aZB1Y2gGH/r
ReX7xBFIskOPXY12GYfCXt00LDfgNQEhe0TMF+UT9sS3an3TzzfmZr04NBEtYQHe
MHou6n9rgN+l7XdEJMFCldMVVox1DJ2sXYvdwfXpxU2nekvaJyTN6U66pshSuleb
IuJ/paYZBF828Xu25nuBlw1OuOZilg4N+4uVbzXRQjqTaC6GS/zTMMkoporHZqGH
+qQrNL+EJ9YQsASvc0cneM6Lnd0UDktqqqKKeTO/zPcpTcZOxi7hFXHo+hvHbher
wYhCHZbnvz2VigJKsWEc0aIQaUsVvDzAU+rEYNvC8c/z/CXrdNiOr/Kr+KpoGpAf
FTqGFhYogLsW8A4cVz9KaAgo/odtGHb+Sk8PhmV7s62c9SZCPu7cO+KKSLRIfbD1
X88kOeigg5p8Bxn1eo9cqJRRVdoIJdaqywUYNJsJkgys6DFP/OFtMk1I6FEVrPZm
BAW/T8QMXXV0KJ2gktL7lZYw9VGQ/WNBVExD9VKyCh4HgKxZreIqn+BCHfAOW3ni
qiPWapJahWB4k5afO0th2U6K+OXno212YvUA0J8VMCQZ9tQKKHhjdKwuiJTHtHP0
AGEhnL9p5CzFd/Y+J0PrprN+uHjhJHciv4p3g/4icF49Z2j744Oc2l3bCAfs+brT
aiRak4oqWFKGBptnfMDp0JUaNAxllfBNgD8xxyWUPeavkTTID2cwmt/XrvCkSo2S
Rhg/lNw4W/bkxNpjsDnYv+IHnLpqgObM/aalwXtMShzHqauQWQkXj5JGeNXw3AFu
MaH+mFcnsq+rTeRHWpGVLod+Ix5hbSrCVtkM3BY+iqWKhcp5SnneLng0WevChwqI
LjeJbeCEjMXGiMmNYbAexk9JkmMXpS00fZ1l5W3J4TEO8eg0Kug6VQhmRdFfT+ge
HAU0D7NjXtwmayjADAimgQRhMJqSdwsKeBNgFr4fhUiB0ZR8m+w5cAaA/Nq+5JiJ
mBupBwfHfTEE1T8WZlRSdiF9mP00NbaANUp550yxU3/HF49fWa59nykithsvaO68
1mybrt5Wbl6TGEpzVp7aziSgydhaFap/GvjIXUDFzh9jJTqqI9wQn1nhvrfNSXSF
UweqB5E07p8SmF2NfJaNicFHHGaqQceYIJrvr5Ad0NYU+vo0y7EQnfwazZEkZe7G
vDgzqi7p0LTyRaYKUhfJg7mtybaU6ZY6K+awNrixDD2qpMMDaqNhtjzeWAD1KB+k
Vv3PzfDDXJ0vvWgbAgYqZdoI9ihT+R8UND47Mq3YZWaR5f2QIyFnmLz8ecY4oQ+z
dQVM+hVt6R0zQCKIMkm0ksSPHTCwPTxT/OVJHd/CZgZW2UGT+xwMjkc6MGnjvsqg
8e/l3PJWSCdjgc1eduX8s4dJTX6y18VCPYccYCO4mANR4Ekuzs4haAiIkkNUdsvD
mYYYGkezPZ6F0BjxCVkZ+6qBbhtK3AU0s9nnL11z5L5sBvfVKHDPLuDHq/pTeQTK
X3jTm0U6oYdB3mE2ZehNM3UmIf9yLJwKTxZTslhjlsqQjPVXi3kFcp1YmdYX1jsp
s1RdnNZNEweAdCcqTdG3er5iNw8Ee6iMMLPITUB8WTo+q2njT7Vff17m2roUVidg
wQmftvU1ue+XV3cxit67ZXlZ1TnJ/0nq4J5yPLgUZUVXpOOzPleG6cLuKopIKn6G
FaCCy0t30XQdUkGLGPHTpT+YsRKxQ5id55b1RPaK+0fCBmVxnNTn4eZVEWNkmQI0
P7s5FgSFzgxDc2UdYIEtMRaw2fKvd4DXlyDJ5saY3cR+yxFIGWknURpVcWl0JBvt
iov/L21gKH776J5SFbHtf4+rZunERb5cqH9acx5wQ5X79ifYvP5u8lrNqjS45Qk4
dwY/8HpZiG3oCGpiOHL02FPN3P+v1Y0x2QC5qx8jDiNbM+K/SdPRxLWDnj6rditc
73evmnLpoKfISskqFIkmhSRY6KRcx5f0Xwv5UZogjsVCzb5/QYvXoXtlK0TdmH2F
8W+btfDpKuC1OtIq9bKtCODFkt7TBxO9yBILllPNLx4GyW2A6L5wKKGlDuO6TOGb
oVMrQZteaIWWjDJvuBBHiDiD8b9IMnK6LjJXMs4QT2HDmX9ecd4AWtxP5AtpfeXn
ef+ZyZwQeZSxHTIRu7BqByrz7zaXDqfhDHu24sAbSCv516V0JfrR2jFbYmxc6KaB
3qGpWd1f7WeKyLsXIvuI00b8vm0Fwm48bavEsyrhQie7ErojF9Uu5PPq7jGHbDdB
Wsgd1eRWAGOZ/l0VFXokTlmwZn2bpOZVUihEZ6ojeTG3Dd1UpPuXw7G5qzKAXGLQ
XKOdqq3um6DSgnVfwzhCD7O1UAIAoEtmlzJHnOTsnYYP14JpznMBDG2QIafIUKhd
PWDkz5E8PWuQaQfvaYfGTSe1TCaIVMHEbPVzbg+kF2/XvtAEbkYQ/IRdhiIoIU1w
pKEVGjqTX7pTdfi43cgol53qrPOmLduGPL2EXh5S8psGaauB8O0Mw4wtifiYcW5U
f+KknKnMuA9P0d9t0bEpCs3WY7YCQK+p+XD1Hvetqv5KBYQx9fm4aVWxqOD0DpyD
2wpEJIQDfwexguGM34ukyFwEA5WoGGHhUY8xUGFTGO4Wm2snMZCOnwCAPut3fumr
GBrjCf/UZ98ytXaeIu4K/+MHsOjGHuqKQgxVxyl0zjIbvtsd9SC1VQeShrcW+C0u
YH9SYkcvF/v2aSOyveVWj8brG/0S38Nt5Lhpy+bVnO7rhfy5Qt83shqo7rOdZJ/L
7S2onGejQdQVhQnB0iHCcShY/L9bRqFoMRIj7owZFPhUiFhi0TG90wkznPIY/zlA
1NdQrtwT78oZO4/OHW6AKFZAKQzoReRtJo7tncvFRH//isEhdBJhKeoQcqu/R4Ik
FBZ9PThp8OQijEFBIda0I2/AM+JDNN8yflWXCrqm+mSlTx/gbQgNN3tjcpiZljMS
zID9uc2h5sP1JVmsciBo0/X9MjPfM/ICpizrTMpiUe+h4pJrkVCT1u9t5B3L2Hog
EoBhxfdSe9mIBaf94O9+yknNvBvFCxlJuXcvE9dpEJQ52b8dpPNohecD0SpFs1BC
mS+rUIbKxIoKBCr6RNkKL0GQIAow5j22jEJPBRWZR+JP4qLaNfRAj1chIct+Khbc
DXNxV51AAtzW9N1PYrBTWPd0bibtyNrJdjGl9PZ8ZbP0c/8jYSz8cfiMlA+ZlwOg
aaLbO8GDt729LnW+WIXjd6kpPRV+XLG6uhzCEDdu27zxw5EPwybFYeez4+7ywvJh
t37CRj0Jh3zl/tLZnjULBPlASKreZY27r2iG0l1PwGtzNw+e8ZBWAr5tzW3KFZXl
3wKStSzg3Oj4lVhiA9nrNeCcXS4lqUHV8N3aWr0ONQ3/TfE10R9HCik0B4RCpq7K
RlUUj5mMX64+ZE288U7WFWdapJEZ6NRGlfWZ+MA/HaQJy670eClTfAjuqarCkoep
zYEeJcsDvkvYcoUBU3buaRWnoYlG6JdaAxOvZBqRZdBMB6MzU8SSa/nMcdP3ZIml
CyGTR+Yc4LlIme/jCAgJr67MXhGjmVZLLdkRm7Rt2RroYSGRkSk4bwq7E//iuo8V
ltGaIN7IzpLE+eodiLW6X0zK6TP1oIMafkf8l7KHMUTo7MBgqPAeDU+mRdqi6vje
SqRKH3GogJV1ZeTT+uDSDu1Fioh6CeVnC5YLpJBoilCkPSV6riKRDdwIAf9qdxyu
gbPdBUrCWF6p1CVBIGKV1qpBgf8xDwhohtUKSUBPGVsPqSW1qtw+t2zS7ZPCaVga
NcgsqtVrbG/t981NqJscYpdBFNDUtCmduXh9wqC3WRlXSAnbhIQbgRthfqfL3L0n
UwUoIIfwjsuIFRq8eEEZ5U8b5DyyfB1K/faqBYE4Tg12iJJkeUwqJGFmt3ySF55H
hKx8OWuIH2YnCo5QxS69jMpEdwqMrhEQfqxJMfL3WJFblshOEzlO6OZZ1aZXYVzQ
WqE4Wo0lKj3T6CNEx1I5e9NjJoBixTQfEZIqnUogTMj6QWMteeerghh8hTSMJb0t
OgiXe2C3IkUtHuYo0sRtpKi28c5UgMGwhnQ+Gerk/JPd5uvXZJGcp6KhryxvO61o
nZuu4ujz7V5qL7GvQaTZCxxxiGkYxrfxWOeg6mMtbUujwpwAab9IL98Af818+p4G
ReLLmiIH5nHYg0QKz29mCmAc4gMiItiZLBwcBnlU+7X8H6lIpt1dU4bZvXFVw/or
RarKar7xGCxx5lGEFHdL0KNBQ29r4mUtX5q2BPI3pwH0pu3f4wsaQIlRYn4m4Gev
ImSmGW+yxeJUGTF2EYjnRGxSyPPiFQlznrrskmOWk8OfZ0vLFeTrRhGf0SYExb+8
XJDrBKaaGzvfSyLxT4+vCw+/kKZ1W7yLmKcEmu1wa8v6nf5FxSGq4qe6bBH/AIKE
xjxGxH3eoCDzhS8Bof2I/k4xicLcNyFNc5olv402ozPsSljJc74/PtuUZrsN1ZWB
wQ3mo/hja+usvplMqLj6b7Qi1XZQsnFxCy4mgsxBuJ45UcIp0QSFtC6igkDTj3a3
bGkIdeBsyDj0X/5md6NK+M5MgoLxLbXkwKvlu8CT9HYb/khU7hBMJYKKLW905f66
XuQmWANfuiYrHQMRrVsMubJkKXNkAV5g6qRwn7G1R7cVM//Ms8dpI6iSHvfoCXoA
5bWu88Z6JDKjgiv+Zmoa9C4+MTlY5v8EkIOIQSAYXDvb1aXNjv0MO24Xehl5yiRj
Co0/J8S7T4EHXIvjO6lOx2t/D8aBcZv/x1zQzVfbYB9q0esaDLysUtNI1vYpoFd5
F2JdtjtSb8OHnZVzSBuXseynJWNPMDyd6pEV/rlLHBH/n44JObeIJxTOCPR7OE92
Wj/EBzBNXiWSZQhgiQJVpGG6ZA6zqLXb6l8RA6uditO6T1/ZFHEe9eFjx3m4VpjH
KQhYFM8iRBf4HR06EdjhKBHv19fWVMSPvZxtKxcsFuK9nam0ovx0FGVW7QL88y7J
bqitvSZqa548PBflPfvCeT7xU8vu4oIEPqUiT9mfXtFCJCN4Jc3pHrdxwZ1uPZpF
v5MiM4WJQBtLyFNBLyAEwFEwgA9wDmdTA0woETRbmsRINde1f9EepR5ROJiMDh7Y
II/d2nG/jyk+dmoFZOs5b/nTz9CqfFAJ1yzK82dpI8bXJnE0jaqXdyI+4BnxXcrS
yNQKTn1FmYZNsT99zIdPhcfYAn9A4m0SZC8DgPp9AwZs5O88QxZl5B5yuJ5VuhtW
/nll0psgQ30nlof3asZz+P1sn7qt7vdksCqiBSZbH1VWP7N08kgFVovWCEoodpYQ
fYkU59rK95JZHOCeUzzz3wQHm6YplA79t29uTy2zl1RL+LmpJD/Y+GtjXePYoMQ9
JTpcFfHjMKNArfKaj/w18YqIRIKH2zdDT8QTBqC5HBxeSt0vENVH18RzsBDWlmmZ
cywzuohOKtGi+kRYL1YU2bR5fm4qLFJaJEEdgNe9H3bT6waYZV0UhuFJiziQDZ8d
tYVAlE25OVGlCiX4ZiZl1xb/tzeQwCUEPwdb28w+Vsq68zrSVbiwtwsp6TcUqjAE
wKcE9JsKY9MCmE911VSNmmh2ciliXs2HEKLnI1DG0wNDZhI/ETvJXSE0163nUkDp
Nz4v5vRqN4SHcT1HSBp+uLspaqjhDTq4heOqjrW0NA3YZ++gOdRLT4goFfrT/Kcy
E1ObUIC6FUfZwATOhVTJIG2LYidrSr+RT6iQLmuvMDBwTdDgjIWzNSoJaDH0Gga9
6X/p68bPBEsvrhhG+JhdeDrb2Re3vw8DB6fmDZ5IvcORaQJ3T8VDaUlUZ7/wddeo
3zItwXIMOmoChukITbV6TwW/Dn2QHk51mJQCh0Kv2jGMQS0EpQ31PxZuur5EYr1U
6ey0vA5NBW9mXeJzZes+ABM+OwZVDsptThirN5Z1QzaWXfW0t1Cp7tkUQUeKCwba
k75txtIRLoacjM2uKl5jXgurcfxpHFNd/LMuFj6uuSag+4SoEcs6eqGW71ExSmf0
ZhNt6Ir11qpVgf7OlFU8Q2ti1JVHyLB8UIhhTShPy21MajWlj853GXj1BJ4Qxwkq
rdbj1YSod0bT/ZsqBXotBQAKvdeGsgmKJJuFvIpL6WBDVZtfEj8EBY8bRteavaOq
GIbrlj8/9K29TV7YMmRJBQHl17xSAsACGOewSB0ByEpCwZTnWTit7V45GFee9geD
E/uOIGSRxMrU0QPQ4ENxZRWeAg+HqYxS3pUeS/BVnud9CtICgzh1czahp5wdKG6P
uWCsCOeVw3+h0bVGYiP9NSn/ecvBIOzoEZHSNbRK9onqaHvriwp192UOeyNogRhM
e3eaIwON+R+ZgSLFT19UrheAfhKVkYHNcrVc/gEmuUBP0g+k1Ep4f2rwscDiAdLL
Zolh7veJStGIAZJBHuWLEAbq8OfVg1E6AQe3iqHG1vKtPgvLzucZwDAmRO2HQyEU
qXrrKm5ACebXMySaZXAPZ76QLtZ1VfiCj6eY2pvTP3er6GPkIN3J6qCFUsUjR8zz
PnmenMSjLr8n8Vo/8jB3OPO2P1OtCnQuzXeA5rxqvJ/vwPHBcuwkEryi7AD6wYTj
PXEfbBn6qZwoN1fPPVzL+wmfycS2LpIRRjQ8q08UjmnUsUjjZzG0C9SWCnnFhA6D
X3S6XJ3PIFaRx6TX9LcR49guGyMop0Bk9n6YMtvTgy7V1HHk6hicGpPjxzhIWSs2
Yeqr0Arzav6gQr7rOxwaiX+tn2pfJvOLkmwQdBMlL228Ya1KmUFR5QZnUlTlND7Z
4Nk2rwAPvHy1ZclIdsKi8V4Ni/YrALAduZNYfRVHgn+6h/1JlZK/8cuknZ1ZqGGh
BlKTCZmWzrOyqacO5BAg3Xm4R5jkZVnCO8cu3BhVLcxe9nJJ8imYnUy9CXPyo23V
Z8rdpMyBVza3fDOoPsAVqaOW4H2i6uHkEgTasJtoXNClaoSkKc5qpgybCVkSnXsg
D5irs1f8gepnUJsG1zqlLmMUsJU7xnXA4flHKTKM8etg64lgdgiKjD6YMY8F4sKk
wXtT2A1iyU9tChbe96lom6OOR7mIvJP5P229KAvd1n1YR/e7CPUGqI6X9zt+VD5o
YU4p9wDNLjGJ7hw8OoOsciXSPqFwm93E1TlwGzp8xdHi0biQji3SVQCFKf6wgGUo
PyGdlWBZtN9xF3ApAOxyqtJVFndQZ1jcNwZaXf0Ov/qzM4g/Y2zZvFTMuaxNINYl
jYBk5+lxRpnyd+WHXwK9IiR3zaO7Y1wVSiH+LjYoSUCyS9tSVKt/R53c7FqbZcae
F/6YIkaISf9E36nx3i6+Lot/ROjvgWiB/YbBUmUqZubxp0/+wyw0LFraMYxh9dEl
B5I/Zr2dNgXWNXBq0BvgmBNTSB3WHRqT3wi+7ggB9QeB791G56A+tPNclY3bvnCb
kHgmDdY/U4ckfPugybdxC5EzGS1kd4g9Mv1KaVdQV3IaNEzrIYhOQez4GmfONoGY
YqRcNQTMPd71imLPICWgwrBFRoDopcOBFTaRPOI6P4Z0jgpVNx44Qy5SGqP+zP41
FdQHL9HLyUEkCr9JLGrRr+ZGytnoO1oQJVP4Jf3hu2e/TwFZEqDeTRB1oDdOnCpd
TiQXzv6Aaa3b4VjOk1rlCuau3NUFEpChNFIDqEHqlO8v/Nzzt09N9x6Y7v49WNAk
3GDCFUdHd9Lx/gafSGTrTvWLUrT/9e+N+aiokISHBpDCBInijJbWTUpqOs/B538s
fagiPM3pAwvGnxKmdypj+PKmkS96RAGyKmarvWnnbX9IWMZasLfueKukw7KQh3iv
zR7Xqwt6HuGyUxF+BgTYbH5XMH7lUMfZlgnbXgsHg/Vb1ZyX3BEjFeNpdmTkAqR7
AlwDtwI3IxFGCcnAVpvUFrNwFLQQbyaIeC68YjcFddvK5EysgV3jfH+CZV5WkMyd
fkZ71L+8sH5bcJswZ9o8r+SiScEm0Coz17Ffv69N3UXnoqkLFgqVg9V6FRVW0U7h
aputzYE42cavvyGlX4tj9wYJnLADkWFkX4ynohyMFQkN1WCsUb5DP2ZKGIUU3X8T
0FJv36n+C4zNZfijVISN2DfuNjasYFKFXTpk+RH9Y0Ol3NagUttnu8zM+bYBAXpr
v20iHj+Qk3SHpLVM8V3X7Mnjws6ZrHynu0Ik3vlzIGmaMOS3/TTTO+nPEJ1qO11/
uqKm0zwHdc6epYUsFPK0Kar6HHhTzidZJe4ahV+Xnr0GAyRMPW6DSmdOHFY8SsdF
CWvMktCYvgRylIm08t8svAafx4xNLRNMx7FbE+7a8eOT80a91wPcq3XD49rk0/FY
wLGg6c2I7+caCDHa7eJ8cyZLWwVoe2Ge32C/1fRfJLIlagw76pLii48//svbOqiN
bCloqbO39iRniscwO/81w97fQa41PTTOP5ZvaLjfCU3Lf3ylndauLIBNOCFUbmzu
lPhKtVtSjQU0CkIzs6SOHqZQ7142B26roaHHWzTknYtHNF5y0sioJn4ZaE+3DCNi
/wQO+xRusCUI47sSE7pY6PeUSH7bJjygdKmBPvgyH8sXBnz+LROkbDV3/PpbwVc2
jzf2CfGJR7r2hNtEVESl/VXTS6frC6Yw/kHrN04IcGzKE4omHQ5C+k5/86KSM/0h
nLXyI91EigZGf3Am2b7jMBo+D7wIs/DngDfDh+hxDDoibDs1bnTG1uXH8eqQcg1h
nA4O5y4iCdG7pyCfNR5GwNSdnCBt2fh3tAEqtZZkyfjtG1c3ZlLScI4ledoEjn0Z
Dh17Z5sMKdkU1kJS6LsHmxG6Asb6pNnvG7cBHMm48nMGkFMHZMAVhx7i3MU1CWkd
oNq6gpkgt2fMrSzS1pRmhrevFL2hQUC+VexW/Rlvwg6I4ubOW+13+XoHNKTb1IMA
tlb9OEVHcixl1xhWMfz0CA+0xJehJHyprzDvtz3aJy11yhkSXBcq/dTQuU2oSH/G
yktkfn6oU0jXN0aHKZdBijMRAvBUjxVeoxURuJBoUNQ+EUrI7RjlPudtsI+ZCXyC
C6LucCkf/cXDHlpmfSaRQJ3Csst0YT6nk87oCmBNEWOm/wO0xPoSP7Eb3+h0Mt3l
hqOC52qhG5qQO2FVkNQVv8d5ALLezl4OwHSUr3zrheqc+p3omDcqFIT8sx/Czypu
vMKHzKSGjggCNWhu1itYBc03XpjIpQbNZsDb/O9MhgSNJqOERq1K+xK8sXnogs5K
6yq25mLbnQXgu4dFGtJvuevpiLEsCXudK4ZoBV1UMgZeFX6eEswwha/Iz/Rq+V0W
YWVWD7eA3/xShd99cUdJBEfXzStMOxrnHODMYQFc5wHJ5hrch6Oz0gbP+4dI5/+9
VMzr5JMDZ67mp9mhnrv+GaLa11ZqDom4HgKswk6IwP7XHafWGZh+5ipnGtDqqSDN
DyqWizHzuhi+dqvT0PQW3ASHnC27I8JV0Uhii5lxEYm+QEJ1hw2Dt/+cY/sdDYrb
EAjct1ZT2VFS/fAe0bpnJhNKgIW6ZJEZsEvQ8ubH+2eqmr9E/AT9AJbHl3SKNy3S
5NS/FCZCSXzSqhw1f0XloXmZBsrsUFBNsshcykJouVB4GCkk/4AumtIeDBlSKKPz
+QRRWGRPgCl6GIuuEc+YbH0zvIJkSnxurhSlB4GUgS6ZWZrF5aNhI90Q5yrtgW3S
beAYHykddvbkiDdJlJ0647H0Xqz1oi3/3AA56ggmWNeGyw8u1KxGYp59snFy93C4
BOp19pqOzpv1srk+wppQTxPcomlKxrvoMBhrOHj6Wtop80drQ31P5Ubu1b7du6Ma
pNi1HriZfY+5GMo6cUiVLkD0v1kf5hNZCgOOGlgNitTRnbt25hfyg2t07w6bH0jx
emwpqEC+xqAXuRcYnI6vSGCC16t7Vpr+6Hh7QXUesTTQdmnEjnbx/E9jwHy5wR4A
QU2a2HlxSKZsY18Qt3iFyNIdfDU3Y2ViFZowNepGA+yB3yF/MGVuMJmwEo7MH61p
bDyIaePVDbJqWbtVHlaplu2xYqdPmOVmkzU7hHnXPdEsX08hFozyYqHvN1U4vkE9
Jl34DZU9XFnmaqHCreRj5fIIQ+EyFoyW3LnKTPHfgxNCPxGrzrykSiSm57K9fYc5
Oy+0Lki5hAwN0tYSV9D7BprKYVFNrC/BFJn+NSAu5Wjilzel2VP1qHyuZW46RHEJ
SQN7+5w5Bfd305v4NT/L12hek694rzvE0dk19b40iGJeaJQrmRysYAgRbhjQELXh
cO2yal+i1ghd9PLfetsym5qLW3dU59TnLJ3U0T2HvLmVqFPjs3sfKnNzoEv+Ycuj
1TvLOIBikENlBC1qCUMiLCq2StX3eQ2MeWUqZLqQm6lpGJXvjQN8lmWWjry+AWuW
zz7FNOR40cMRoK9/A01FNuGaK9GZeU0dG6SIUEjq+1UUmXfKck85ll4rm7DJLD7V
6xmloaS/eKUGqGEA0rE7vmUmtMqjjpfwzs5E4VN5FwkLxQDsfcIUT3BsNjFWRocf
WWvr8QOd9G8qMLxZW9Cg/bXGRAkzEaWh3yYczvf1KgssB4Q/bZNZ/6UYBXfO22/f
ZTUcByc3wNjxLD1Si9aJLdSOLu4O6pUd8NRRDgyBozTUOrARzUctN6azYMoBveql
lJ98D9WaV8RjYOSeUoqgagmIoV/IpJ4usba6j/k4E2W4Bw7mJp/jy5sQNOWNsjEV
24UXk5s4NNTC6iCyGyw7eyfnJP9Rlhf3stmFHgi9ZQPckKO9wdjfczFlWLKdDupB
kViW6q68RrG9qn4JrTiYtB2tWOIRxxJSfdYeDPnvH9tlTJgvFY5zTevwpbGunhJF
FWt3IImz/WBP341JR53xhYke2FuWNJ4eE/6p1M9kFqc3LwUMQ8DueBklmOQ7r3ch
Ermq4PjLqvB4TjWjj5sthjt1rkVRcT/59dOPL9QE7XdrUporbSVi5Vnol+wD0VNR
8DLJLghcYWHiHYGYtiDTJjQi/3qu62bqoidZz/ZersHyZ1sAAZ7WO7EUm3ycEnzz
FlBPj30i17oZ9235sSz4M7brZRXiC60kvosZ8PN8h04Xao2X0uxER6uD7y/I4Rxk
zQRwJMAdM1g9BlLCy7FQGVt84hbuxQbd4FXXwfX35U+hkitVv1kaeZL6tqAF5jXZ
MiCGO7atHOixNWcYj8uewkUGcNYXTwcaj1+XjP+AyPjr7GAvMVZUV34Tox/eSU8A
nnu9DuFZLZe1QM4ECS26R0eOmwtIIlIfCbie5IlRU9YMbrOtvckuCD++9teFDyDc
X7LrL4DVVrS0QY1gOg7WePWtKt4vE3gTZVd3lv9WSn6qZtzHetJMvp+ei2DTNdc5
IjFr/wRnQv10+hA4Gxij8HnwTNBypNhqUmcXKvw/PcRIjMhG0/ROFTLghwz4fBXM
bv7MieoxyA6EJxrtIcOcX+qYZ+ivTAN8yJ45dUVwDoaLEvwE7FxXm1qqM3EE49vJ
23AEq5vFAZi1bw6F8qUEujXOmO8FVe/MbWNJNdCUA7erjOIe8Wwv+X91z+adeZXh
xoxXW1mtHuNUKUvgfNU/BaZlYTo27mkutXH9ctbVYlvdDAav7Pda/jArwqmJqCa7
y40m+hky+Bx/fJd1yiPfhi4+AUusYmnVCZnCF5rbCpRBWNKw+PyI7uSZ9x+i3XPL
dZOeeDrjJc1VCnoEvob/FDTBTqZkWwFZ0X/hrijv/x6qii3Hg54h5hlenYniLnCy
XsWAVa2QT4cf+qNgER5KweOzYQoPqI7LeKbrjCWK02HdY6DvLlP8i7lyWyatWaGS
ytNEjyanpiR8VFf+r5qgsol0GI0C2rUa8epvw+DKEiu1sir/hTedx21Uf/hKoF5t
R6fffvxjOUpnhhTZVoupj6bLCTZFy0vYMHGy11TFZpCBoAa8YAL89gKJmoRXvkIk
2NpTg1/KEdGLyTDGTImDbC39kdnwtp+f/9TpWrGIgfE/k7rjCNa+TinngTTLsfQD
u+oJODN2GuxmcLabKcPQlQB0OgSEv+aBHDJBb5TJtwhpptTeWxHVAi/vbKVaVNfk
qolsGY3Ab8iKhtOv+EVAQs/YgiRtkzE7+3Jm6naDGtgtyror3NyJXwRR/H9qI35J
fMFjusJNoHEl08cqU9uoAM8SyMhLVLU4bK/zUvJ03l/ghWqiTgJP7aCjJ5WiSgey
38jnYccxeSePIHWOhRQe7iD0V11RzfaAlChjwZMKyKdgJDSsOkE5R8rR4mvmckF5
e6TqonjUbkjgICNv3Vx21OZapN6Qw8enDIC2BcztSQ4+QJu7VEj3fDrjfO7Pt/ge
Gn/iiLXtabD+P2cnFqpBxs4iJ9PeJb47Zan8gEdsy5wZ3K1G2C9wiCaP1qtp9G4Z
2c6En99+eXr8pvywoKOLKEVXq55L1bmK1LwKpBVXCydVodt1j9FDy9k+wVhREibp
mbB3iqdAt0zpKgePVgOGvnh57C9SCcdKoUOikmxQm8cgJ3ZXW/z/c11RYAKyd5HX
P5L1UaqXMx1juJgMjZGnB86YgiXkNAOXQZET182ctCF5qi57NDPSOZ7uc30HH3Ix
H5ILCHe3oRIPGWsK9o2VBSh3OAPuNC4DIv6qS9UCSK9Sq/qLZoQt3mb8aFv6ZM6+
KsYYWqOjvlNC5rLwkRR1wpQv/vsdBnn0GdfGG9janYg+AqwrsZuzALCM15Fc6Kxq
cJTjA/KW+kCbozCZkGEjmPKLWpEVoV+fJRgy67TnIh7mCBjivZeSATxF+NNZygtQ
vd1IwBsHJtvKDi3eZQYe760sHDCJVCHA2KOLyW8sKBB6ZSvT5tM1wuD/XlK/brl1
PlAJGjdr7MoR7gplxuxQ4+E+hi7w8p20XyE7My5vWbnKOmlLuubw9mYOsqzChCEO
b7cPWS/0bv1aDEV2+3qI/Wl0CbENmC4xxqihvLFNqAKYcPiUOBlUcljUAoKo/Uk8
tVhIFBRIBAnYKexI8rPQtYGL8ShiF1NKJM7POezH00mx92T8pxIh9V2dTvlM9VEG
uno2ja7IY8mp0h8mmPDKYDB36SQCEVS60dtoIjeToF36r5yE6ZuSbFEcoKUti02/
NzkFoaheumPQ2snx1JBXZ/o0rriZIRI1ThiJhvDZ6VNAbQHGgw4ac//l0JDraD9F
YErp+lbHD/QqTOV4zNDkDXzp8dJCTdbnuv5W84o+yjNzdtAT89aqnq32818WA72Z
rhZOAoWAYSh0pRqVzRjIP0CeLlLi1rd+LeR2tC9xk53WqNAnRqt5Fv5crpJj+ZSK
XQ7C7yno+0oCBPrAqGss28jXOU54ppFpeOkJPhuikma5fa7XL3/uyzrnHQImXsZp
EJnjlBjsI9UFw/fGJaywAw==
//pragma protect end_data_block
//pragma protect digest_block
Rv1S0Z8VNZs+FaV1tfSxixwHJTg=
//pragma protect end_digest_block
//pragma protect end_protected
