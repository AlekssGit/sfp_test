`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
dIXSmYw9c0orX/UNqSZ0VE2M7n8f9ufmTpOGkxuUrFaFuU2YnU2s43beVni/Eug4
C6J+Wwcq+YZCFcyNpvvjklx7UpdeO9j5PTijpvq4bnWL5S7gp52diYx/Y33Ppo9N
QK3nTEBzsz1eN/SpFu8dFw8FVmLWCqYVQJd2kFjKAMw=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4080), data_block
ztDtvGukLz1xWawiNIKgl+Bq8wUxLEh1waVZEr2pU+rMZGbnENr8neY7LUzWgFvP
4atkCF3fZzVSW1WowwlvU1un6WrJhr085Jjt/c0ayunpuVxH88MVpOKso812GYRT
/cTsHF35Abw95fS+kmilqrCSYKdm2/ghjmnZqh/8+fYmLvzwtXp/2v0S4ENELCrG
Sj8tIxNDTUp/p5lBHrBnsvKLSxtUTNqvA21Uz1NAA7hAy6u2QzDoY7S9aZMv2SsO
P+HdHwHzxot7SH0yD1YbWJeFNSMs//Gnrfsjcp4cGg1cDgx9fE+iEHkuUL86CF75
KdeBeSbELlmA8DN8UvCfURJ3YCa8Q3S61sCBj/+oxuO3MGVSmAQmMJHMMeo62r1O
kmaeUnZn6ojo7gDPs5cRFRoXe43eg8Q0rrlJH2QbHkIaeO4f46L061KDAiLkOLGn
x2a5oJhhUIpU5FdG2ldcPTZQRt4CBNC8KWLtwj6TEjuVw5UMo25AyUX2zEZeT3FG
A+ySdZvgTgVhLRlKZdDQUrauyj5XL1IQRoGmkqKgFDji7Fj5vWPZLnuxL5EnOSYY
xiX2YFUw5QlK6BQI2zin2yXsI4Z9ts8xFirBAmwc4hMdCezwc3i/kdzr8k6XIr0K
dhoDo1SURBp7Y95rQoZe4735rCO2HjyIOyKNhwv5l/DNEIkB/sJB9YHGKQ2jNvDr
nAHWZwRUy9/NvlLgPUGSiNJ5t7CgvL4+Ty8KGn21RQGVenraoNRXqit7vsMhP1vv
p6C0nzWHyxpPlD+wLxCp6esN2bQhs+06YX28bJDd9I0Emd+I03a5Po8BpV2m7oED
F7PyF2X+riM//f2HDTzoV1jRPjRBvLfOnS4K9npQMNAfcJZZf/3uKyHZC1Hf+e0L
DVUqM0zihnU64COLs5ISPu7SdpEXF6NODqNsIS7H6bDbnM7nnof4/zsBF024XDsg
b1S8pfhUzc9vuuq4GrYHsJYoCd5gbKp7j4T1i5mPCRVfHwR9FguyG+wo0uWdYLPM
pNVU25OIgukWiHhlkVOF51JRaPX7p7ol6FYcHW9xv0QqMqEBKIgLN7KLHaFCGJVO
8ZcCqOtLCjO5xoOODqe4tPbnul3NzAfW4xw+kmgtXTS5v4kTa7gRJfB9nvixSPvA
WljgftFLMMGkjgo+1vleOoiW4vYtZR6so9OtItRLuZMcMtsVAVv+n+LgYYNCVM+G
6tff5UBdGsvbeiqTQI8NC4fWoYYQ1ymTvr+B9aw2kvIuaQarzzLv4g4pamSx6iX7
uuFBJF1r7wwb34gjqFk9Yh8OUPt7HLnjbhKL1xkPQlJwLyBOx/OyJ6JhL3K4E1Gq
lnLOr6KY26N4+/CyDWEiHicMLe3DUm6W05qX6HMV6OSV+N9iIGVr592GVMu1H94z
54eCdsKeskqXOT49Szjs8I+6LjLLDlRZ0pu1j6xWrVLjH8rL2v2UrKBKVevsSkgW
FLjD+tOXppkOF+Y/fm1DMsJ663+IL3foKsHwE5eWOrheubXOwVozPgF8EaINaLKE
WYHEpS7lOhQRvLRjGXzFWl4W/vlFoHzWtT4hevmTeMDc8WLai+52IOEG1PELCjwG
poyTM4wD7XuQ3k9wYinOohDeHG1TR1KzEY3qfAvvDCZDA+FK0nr1neWUjzyZyLe5
QaDuqc3lkatGQrSASjvgIMMEDfEouLzrycEALBn2DZ7cuviKbYtubPkms7q/ocSZ
EbA99NsA9Gkkl3VIUgAuLwft/13M0Q5/kW4gzSN/lnupoZZ5ClwM29v8aFAgsvwf
9/GeFS1Co9dMU3kO1Lsh1toPiXskZdKg2kTZOQy+StzskGAQc5gZ1G2D4hX3hKoQ
JAvbzqs3ufCvGAJOftYJKTRhXVRXuXfFlehPkNc4kEuUDbUwmK1h5Cu426MATNOa
Yi6k1aaN4UjvqCRY2m8FcYM+VB8lcvr/R+jn8zprZ5/2Y3fDqJmCdG5oATizpcfG
sQjbB8aQc4y8SbuBfOejPH5fEteWeJlgz65iO0dSSRKsrS9o2hbjCk4QTEmjWYpH
xdF4tKcNdslxaLxqp2JOTZxF1nugfqQr+fRsZm3fyVBlFBJH72/lQ5p/9FYzvCaA
jpLp8HpgiHAzSCk3Z+pzSyiDT2gaGaBeeUlccSVLnfiysBw+Bjqr70UlsdHduKS2
U6RsO9JX15tCJ1Ma/HPFtWhChxjK36DFutbhFHZ9GcTVXVjI5uMpGcSRUBEojvvH
865n6j/SEejCAqe+BbzgrMk5Wu/H4dcZmpdrhRhTar0eZlG/Z4ivR7fmhEz1E+oY
t/TlaizVkRqBX3A+/TyCcuxzrYCGX80GSzzK8ET8PgSg9BsbCP69xeAzi8lBethy
a/gTlVzaFVWiigMPn/hZYypzfpEIRFEkISstMZcP79XkaGQMLRfQmEhdots0mhw0
VHzqBEeOMCQRb4CfCLwyIsyEuFj5FAhNM6YY8FNHj743ps19kkGcATQtmT4uTW1P
G6t3WYMjj6BFGpKa+IAWCx74OZtAxd7czNuDzSuurGtClgUoqYU3uME5lU0GiEZb
DTrxXiAuSoZ8+Aky88r+z35xAUpDpz1UwB9nsEzcmtPNE9y/0kLSahI8uBaPXnB3
og2DyshSwZ0kgrthcxbmsXfL+LrbIIk+ecqcYMZJVI2GhQO+5i7U+GA5Z6Q/ULCi
q7at0BFjPIbMiEmgnuxwMVuC3fwnXA9OUuvsaDONzikISDb75dGjl3Rpsgej1ap0
d3JjKHmGggzOOpHBd7hodIV8IMSFllA9DDfcmOe0VWO4bbObm455qlT/UWLavfXj
p3NO5V0vpkq+BijqXFpEYb1bYGSQImSMuP1gg+5sJqbzM5k4yepn+1++Fzqp2Nh8
5GoXvGLaKmRwqCXbXUXLSN9rytVV0OsPO4BLzIjkRGSY6WT+iwPBoGbHAVACXTLm
sdLiCJIoWH7Nux2M62LR9udhel8eVA8prEtj19D0vUiV8AAixXo4fEzonHcFHi9S
QVwUI3xYfLsEmVTZXxXSWW9VQJ95+MvM+CwtNJb7O/S+hXoYIfvqtHD66kxjOgrX
Ewbbk12YgIx2ju50yfEhFRDB3nErUXgbaB30RS5JdXuHEuB0ihKbouxxUWTn4+TR
kF/C5THZL29iA4Ro0tdHRXEa6dZV7cQdJhG23b+74k7k/wrwZyM/+Z14MQmVOO2N
gCKJQXxNZN3JchTOLK1HYTWho/zuEXR1ue+aZB1k74SaSQ7HDe8cJQCtMsNdQvv9
5fbEkdtiNCtPJ8+WFM3fKVKkWS06IidIHLJ54WlCWcFqQg5CjZv8LfV2ZWde9KHG
w9mnHUQpF0wy1XnB69Of76Lex/tSYqwcg08SpAgclocWWIKx1Acq08Kc9LPizkTj
v0bGNM31lHJX5CQzbVwxcX/oBzNEp7FxENhddf6n6W1iuljS8d7uNSFSqOk/LNqB
py6AR3gLcqIihHJAXNvr8dht/b8kgamxt+f/WrfLMMirvbifF/q8n8RvSu4orP9i
Vi52s2Czbtu5lGkzFAvFTIL2Z0qpa83A4YpAOVY3rZgnZwjCpXlKSDDUDr4uTbH4
VMot5FzShrmef9uLC2xX7eWCfVBTs8Yf9+R8PI0ZHv8HVuX1f5shuHs2CsyUa1jT
bHm+n+EO9YA2fzhjZSSF7g9aQBjhx6AeX4Y0/qOFr4nxFgSZMB69u7HE+OF1BXKw
ajjvyLGFitanaBaB2nTaZ0AaeuweYuBeCZWEZ7Q25wmUfZclMGSQNsMH9BQMDRt/
l0OYx5ckO84Z8WCuFbBa0uSBiY9LWSFDvFsn1KlnukjqefVvur9bUiK18Kv72Aey
wnlZUI4PBcGvXhSgKV1vdeJodl4GaAzFztZNYBwuTeI6ojedIKLPf7XjwM9l2KVg
2O+CiQ+znEmvSdVodr5MKdMCRTbaSHi7fgoV7xL+SPdnt7hr0SlgHOmxopPKyz0s
TwpGgLb1gJ0/6vJz8oeicQmyanPPjuJAG7N2tJjPSN44P4qxGw4tjoFRaGSb1sPe
JgkMyPxx9ZqyYoLUZaOJsSqT2jzOND/CxzVD7UbPCbo8zvqrAmWidVNIjt+74s1n
RScicv9hNqvTbBTKXmITw2c9oMLXb4OMMHmrN2AX4FKew3f/QaPGehTAueJvi5A3
UqXIAuVEwZC8PYVdMtel9QH/43oFtCRuHOXS0+3zZHeOE+UdANRznvTNvM4l8TVW
/F5wqJxfG361jVSJfBezWveZdrCqDOB9vIi1ysATPLPPNI9LtlbagxJvfy24QZKw
psDgMVZcxf2BILOAbT2XjWEyNkRc9imllYUa6Hd00VEUxnCL9xqlrbvb2nZKaymr
qtHTnJ26XWXmA9uZ2QMni7PxbSQfXFuyGpEftvfkuMSqYMF1Ig5FRhIuIEqsUa/a
ubiGUlg6t0gqt/APRRVw1IwkIJSGoPnwCi725FLWfr5nxkD8XSY/VSUhOtgu1ONU
8E8J3VAUe14a15qVa+BENan/mXmEKCjnrWPFEjJmkBc/VP1lplt8qqKzVos4F5SA
+/KYItxw6T3iOlCmYVN1Bhn8Z1sIJ8TGMd1u0RjZlvofzXZs3YvOdoQKhFOcl5e5
zXrUoo/RGO2/Bfaz+1J223ekFTuOxgZRuhcqcGF1+6XnKKsbcgxvdlJvpMNrfSeA
Ge2Zh6es6WkjywQUw+WeDi9nT8t2oQmKIm4EZOsEbkzM5dNXysSo5ezwknLK/73n
P8zGhuo4LIP6QfjS6k4Aem4oZq8eBliMBIzN0gR/J5yohQLDIGtQYpEryFtvSIih
ORu+fwBt11kX+M4EauEBt6BbQNMWtVyOWZFv4Kx5HOP+vFEN+GyWQ+l/1dWZ9Bz6
s0HCAnf+tkiVsmzHa1SemMc4sDkQiLHbfP5v3duy8jzFGx9MCJCJ9KMwgtKF/cCc
FNDY8rsNbV+eSq5vuI/W9iHpQq52b7Ua74JHWfvccWTZlrtdSlHXyT3dJYqBoMfF
oZwdZO0ZAVyS5Lz1HyRzO++czwWc+Ov57L8nKHXQrVf/ul0bUvEIiIRiOXnf4v2J
oB8YIYdXQHrpDv9I2JLjqx+0FGlkK2yyutIYuT2a0AlLyvaRI5SoODOCdbVNqejq
7l6o/20xJenXEYAtZUOPyAeeQY+nuqY1lx03mGC6k03/dE9LIp+rvzB8Q5lkG8yF
ZtzqI1ML1blLVOrDMTeTCuN5SMNYZaQyK7NfbGsgGqr7rBZsTp44aIDj1pXT5+Bg
8e2PmFsChIOPyy1Mv1Vee/8SQPhRORAVXDVtzknJniGi9BAFOIa7/hftDQnO5JEF
rIW26TuWnGqalRCvRjcHFIJW7YFTOSsA40TAsO6UuBYrtjkrGxZKUsKcLxhYnAdx
QiNDKPHqlDLZp7qpUU5yXUy/RTgRtqpTOt8eRcoOlv3upC+zvqAlweEZf2FbTWvS
`pragma protect end_protected
