// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
pNDN3JiFzIU9nLhYQZWHUTBsCQvQ00xL5W//wVpFilwYAf3rkKXARnXeKc9xKMg3
QZcyjp1eqLfCGfu4VgCvxYznUZG8CGNLXn8WuWKfJefa33oivl1Khv5k4LKWj6DR
sKNyGD5fZK4ICcQSKS/AYZkVqLcRdz8OH+LjLu44MAAEYDZfEDnn0g==
//pragma protect end_key_block
//pragma protect digest_block
Ysj6+4pkFLFckL31RY+CqxvPcl0=
//pragma protect end_digest_block
//pragma protect data_block
ifVhOtQWTpE6DpSjr6XNtzq0NiYRrldtZqpAA6mLI9iPAAiJpyzY5zzB37+Ovk1B
qJQtA+myvVPmyhcfVWP/Wggm36QRKcxplIvYH2RKD1ld06EameZYEvBSgUQJtLYx
Y6jIcF6RJtaOgI/Ms6B6Dh+N6xrFjJMzxyT5seWdO/hU9HYvKz1ZmRThJmnAzH/9
lOfZLnvezzk9L8thT3OG1aPlcrK9mfBYdg/su353jyTHkVs3zLOCpMuFxCwgqQvn
2TUPP926hMwWTq4VWh6j+162Lcv11PRYAzNug6DrH6hF6vG45fk5efJqQqQ/Pqua
OEVIidwmKUJGTqYdt39ClL3tdiDFI81izTiogZV4Brs1xkLEcQo+1S3gyPg4NQsB
Eb9smTwEHvXMzRnYiVAjBNtZBRRGGhwkvk8u3rYFlPFGW4SUozp4a/GVBUNdBBy2
xStHmNMwwCMu3AdC+I3tFqUcIifzE8Jmt8gnwLV8Bo0s/DLq2J59wnaRiXccbyCp
LZkHGFTmTYF5Qhdkt2ZCEjslgxgoDpEhra4+mIixQ/Oe/RkkidW0aXGBZ1TaHi9z
lQeR0xXgdVHrIN6kxmoB4Ryie/qRMBZBabXIZ1nJh0rXk2FkM3RWLyHB1Bt+caTL
61aE3bSlFzfGnZd/q3t1oYAxgQAlpKIFL6AwT+Y2tj9+8G37Fc5NjNE8T3w0Cbxh
t1s4uIDOZXfA1RPp7YpQCDk52FDny2IrMRAi2sIPGzhlfXrTIY2yxq3wuxm0OUOJ
hSUrtviqTWX9sk+qn+Hwffvteo5QcTcT8VexvgBdmVy7no7k7aainsToc4QszCcJ
fKzPuUCcFOMUFJwmjrbYFclknw0rLt5Tja5QWsA+7xgzmnN3C5dze7v+/BrSYEBF
LAo8UXBwEuQ4OMK+BnXGfoOis+PLLbrPZtTy+QUz+8OjWLTKg8LCUGOiWNJfhYqU
COxsbMuOiyOtLxG1oCrQaaUu3xItAMcFakUb54o1Y31BMvYdMWshAJ9Zv37Ajxht
aUEkzbG2UAWG9xxMPckRtwQDr5C2/ped8HAxX2Fg9Jri/UC+HGi3ahazCA2LNDbJ
+xe/LHfV44QWXnKcXE3uoMPqgjdJ+wksqtMBxJqpcAgj/c2auY5DizJuRt1idDrn
8FVhywzprISstZf5I0nodpN8A/ks+Mqx604AHPbSbt4Ul5dtYA4883gUk6VgWgn5
oRAB3sH7p6Qfl2ij7/vbBz5TTi3tNQ3xe9ZR6i06JTL69hD4yXj85xT+LyACXkVp
2l0Gc66uobk0LFk6UxSS85OPrY50r88jNC/SmNwBZiaQ7pexZMzi13+z531LBy3y
3gRiNlDu+7gaqflPalhdIcCfYOqDuUqkJU3fq6Jk8sxxU6TCJ7gD1lVjjFmSKami
ZgoXluHdvHbXm60bIcwnRKzmMeFACrX/AlDhd1jNmAQuVdro6ovkp0NHvvCb7i0e
AxCKW5BlsWaxiHtLm6o14NEUChyn3NzBvOybktf30QHNZtETVCHjJet3iEssWcIY
NvPYv0QOJcJKGD8OndKuabbx4Tm9WUPe0gubO1EcTZXupj4EDBqo6rQclZ5Lsq2W
ncwm8Hi04fUK5EY9/S4w0/jKEJSCzebEiYYKMtGhva917sMBinLxXoRoSEIR3GKs
ix+iG5VtH/jDAiJ6d4ySXUSo3fin4+HL8pTEFHplwrXokq1mIIsZx2jG7O7B2efp
Owh36QdTPobuUp4bDwMsMV6lrRvsBBMQq/s7LOP+t0wwrzCXKx9mfTPjwWZSSZu1
suRBzbp38cDbHPsbm+BGdBHivrwuMz45q1M9a451L4b0ky3y3BSIuCc1SzrqGcea
pg6QYt7c+8xs2krJv+8KbZA8VDjxzSHEQeaOxBLi2zTcCCE6sXE/csvfWM/1WRH0
DIYUdUgcJlz7mcbF1eBzQqW7jkJAtabsKv1UUXgGDnTR4YHuWJAQQYylXFx0vcm7
01c8XIWHmekqkyr5AgC0qDMs5XWzESgJJ8K7itzwnTLpN2y+YZIikJmSIZ3igJk2
Z8kkxNtR7fpmnD2SwA3ejmUMjMsx70JlTgxshP4AHPXfmjEZHvH5uV5S+LWHovPY
2fa/EczFMP9ngnUIsYxPnTuajMYwPxnbMQJLfivxkQAmlc9o1fBP2L6goglnjsVP
WCZc09Cj51M8weoeS49XUT4yxQO53Yw/UYpSO6hnk6wkfZKPpakNvXkxi6Dmq24e
kh24q8mHUKlg5Fxka5PZ2ZqShphrh5/oJNUN2kNyfS/fXrwogFplBm9l8j3aNG2v
8hNCUnTj2KRUjSIfcy+EPT0P0i/lydMMu2tUcku67/JlfuppzLhBApYn2CsN8usC
IccpSNDy/5FtR7P9Mb+CXrYKtgifdtP3iT8+RjRNWvrZMju8S8eWeAeO2s9FHS1D
5Low+uVqobk+KbpbBSfo60VQ0NUu03LM2F3XTuwNw+quC6NoMyAKtNR340qXWUY8
gxyxiHT3d5NA7KOEO3v07Kdm/nbZ+Oz8tfn5FQU05gvHDu2Y+T5XzOw3lJU/7c3Z
Z7uBxjI/UBw5LfKaDyce0kz2WWPfcoRNVVHs3q2zswCPfNDngktSEu6oxM5nixJG
966GDJrLiK9JjMYZp8QHR+xayKB29TXSpnomHPE2L9tRMb3+r0QB56Gt0y7V814N
n4YQvgb+dNaQ3UJAhZvhuZ3Qbr9O3gWjCpuU4EtaYOnlkVtw83OXLH7jjahMSzmB
yQiZ1UKTLTxfmskw+C6123AEJBg461i5Uo0WUfaag+nAqhAXoyiNnr5tLkdK6jf0
IiMZ4xMS7Gg3jnUkkJVRoVg9+e+FYS8rGy2yhBtEr7ReRmxfo7L+H/Z50NW5hCrY
oLKwH7BXwHTSOaiRxp5FsXJY+WPGh0Q+4pIZxkgtuDtFP6CbRsGPVIl4rB3xQvPL
XzJuZjdUYaWtt9E+Zqx8XfrLA8Tpx1vlV1X9vtrikMPmWZ/DSceOqjTKOPGXCGnZ
Ka4jI+Yb9RctJrKLJQNxTKS8AU3k30Sc8CkCkbCAtBZyscDKIjjsBAZCc6Sqg8+S
iCl+lAeXYodxbi9DISFg74n7zSP61KMLBTC8qLE2ZGYXb/DXtl7fM5aJugLDmuLM
99j0BuFJczKSpjjUGQruatM5VY21hGl186h0GDX+QyaT7uJpoAZRRmXV9bDWYYr6
BEPITag70eSnU2BD3BfjhCLw8icF5lZZbbcTyGh1DjFArJpJKKrHEqijOMaFeY9K
sqqIQyCIEOGUfc6UhU23Rru1s1gEN1/pltVe6Y+IluWwQz8KkQtB18adbL4w5uiM
ErCdWCyrKuva/SuYx4boD+WjlvLGCytnQ+G0ROn6SO/czx+tOWwNklwYUOu/NFIw
xMNZl+MoPGdhzp7bwr3twRYS1hMN5WIqjS7KwAdu/KNPXJ/Gymi8sSNNR62GhINL
P2i9GyOed2L3WpR9WfaygIU0VfqfCpoRfbovePi5A8aON9MCPRm2tN7fyPzty01J
QC2/7p3kel7hHcfTrnv5rc5DTleXxlZinD6CHFcMv0RhvBtyQ6FVllY4PCXCk/iD
b+d/xcdQBGB86RJ6wATldIYVm9oAAhSgcmJ/C8ydWgyFYozFlWc5/YpJFOoEvSfm
4K7+jxl8hsuj9IR6afNchHClQPuFwohU8OP4PpYG7aphQeRLkuOUr+hWuFMuNGCQ
Sizemuo+pnkeCzFMPC4Uea+O3ZDN3d2vDfp80NcugBBTQKewLc3cYuXbARaWC6MR
0JxLNAJKxOw+V+F+FMV8w3dF7AQfs19THWAoDZ2elqo7urFe2oxy1fd8ho4rjSgQ
fdYOHujqzk699q97+y7mpRMtY4Dvs7A7jy56LLi1wzajEOVxhN0vGfuT5GsYQnRG
o6BdCLw1FcJEW73aDIT9C3Eqkms0k1YTtZK9045bU9Iz7uDd7J7o+17BtFqTVLMc
azcOTAllBkIE8z/xJVfVXmpRY4Dd46eT2pvs+MJw0dAaGwZ4L81+iTw1bCAPwv4v
lSgc0M0u9bRPw8MAvSujsbjTr/HdpCvAYtNm+VUCByNlnuvGE80S8DSfR1ifdgcb
fTnmHTkPJGmovmm7aMmBBqoA9l5H1j21hllNxCTl24J/na9yGZ3YlVS0Fg2PZikq
7n0oX8wc3QD0AHDX7jraUnBNBJzT+RQVCtTPlEd4i8WooH7mpZaoRpeQsS1Ns7gI
fOiKWJzQbZ2wxW0Q/Wn9OhcW/ev4oCmCtITfHzkaVspBLrL85jYFvfg38pS6Krtc
c5BkggXIUhosXNl68X4LW74W7tQjZJ5Hg/bQak5JwRKJ5OTbmObUeatzK3g+YjpY
VKw5qK4H0uY0YFz3KV1D0VX4gTF0gMkf/9Mog0UjEpMz6odTUKkKOc0O7whhSyvu
kYWxIlA2bBd5ODQNdLWbbO4F7Zm2iZEVNGFzd8VZDQJs1JbshksDCcz45XBjz2ru
z7VfZEtlbJH+ThlREDEolCPn73bANG8Gt9NiVMQPEEH8FpwjF4UFine0Cgmyt6vA
gaYkGGX0WRDdSoLq6BhjV03eUMreUOMON0FaGL89hmVQyhOoV/dJwfarm7SvGXob
vn3i00gFVz0fqObpHlLZkgPWP/zOYd6yzLoK71M1WKqhyP8/Abss5VFsNfIiIbQ5
eUEYgZC4yjNhRirs07iiiAT5bv6tNovR4PR3heJ156/bu0qjSflmTrvnJc6iSMKl
DwhUSAIeYRGvqkkN90dLvd+KN7pnHiMlpJ8FjirqNDNcjCtbkApfSv9l/7RCVLR8
W/AGwNlp5OWkd6DWE7uyuwTStHgaJ7TiPZX/mop47QMS1qhW+5Lhmldr0Tpcbepy
xNfVMFsvX33aSNYJncJpnUQzwPW6KwL4uVb3kBtKyxBXSsaAYxyWd5DhFM9lKGzn
5yOaasYVvRPderPgApj8D/lZa2Tf7euZUfsyfHmqH4Qbj+GK3461mdFz6pSt6UyW
DhnGIaUNepYAihynMSKQ4T2uU8TkeHF3mILcOQESDNo+NPs2t3sQQzEAfyG7QCcn
zb4UX6do6dPAoWn9jj5CecNiac+f1e3KczOVCz0JPOv5Xor2YgtC5WktR98uzASP
gP8R1SNRq9+JlKDUZ/dwM7Y38aoV/Le5PEP66GWfOxfcm0q9/WDj94mDjxOe9DV7
Uqjj7Kc6JUYRflwRMcC+G1nMhGxI81ke8jBuwsFmVvYbU/FWMDAcjew+99citETE
q2Xtt/Aw9lm0lDB7XloAokSBJ/BUMGZH28SDXAT968upzcVAbXJvUOlcgeucMxvl
j9dqQm1+pfvyd9GytqzJpuIK+KmXueOttFs0RBR8rut/W9NDFq0x8ivJH2DhwSMb
K3ZSBBIBaxZ5mwDJlO57cLvHYOc5HvttQcZSqXrjPyZ207QOi+gKjhxkBT2o2sJG
zg5oGc18QyqB1rpqonvJyUHgd3lMsNpdq4goPltPtgucn6s1nBWWn6+Mi6VijwdA
XFd81o3pDHVifioctYXMM+foGCnOrHdOvFSwZzQhU7mSB/IOGFVBJfXDc7/EZXPs
xB31uBAxUwLGAKvIR9GYYBya1owXDTPhoFK0bTZXH+NHlU6JKUpSgn9BK1wzp00T
v5REFLl2fWoIYf9BL50+7tggE2BC50OOX9LvwoQBkptATG/AYK8OQ5/Vfu85mmGp
yeamD54EzgzEP+MPgKaFKB75cYY5qDAfhS2NZW9wQOVRUm3VfoPkmc4SFMXBKUDG
hqVOCeU6cCmRF5FPfzSOW6Q0d0DVn3iIWKcKyY/vVZ/crwCvv9iARHyff+Ya8QRX
hsOkM6SRkOh8dzo7QvSnxMivTC6u45T+wXk9YM3VvfinPgTMWj+5RuyVdoRxdJpR
BdeXxm/RsL3Zf6hEvygS6f8Cexxqb14yukOS5gT2YlU9Ej4eYBg3ncY+SQ5J7gfC
K6nbclJPSq3OFiJ8fqWW7jkDOxhp+hp9TtklMdoyHfKzxQVGKUR83S/OOBfBt5mX
UubACQ6Y8MbjcufThG7aVJ2diCcjMQacaiEJmzTWZbdNVEGR975P5TW2n9MGIVCw
CQ21IKUyL4fTQ2waeCxsjY+lmmvnPOL3/cSjtw2xvVyFHEiK8K+kRWhPiv1+cNya
Nk3Rxuzqd+4u99OhL2gjKPBRY3ODLGgm0PWfe69T4FauCaE4WessJvrf0YpaNed4
fUwhbw54XNgiukI6ltG4mSJ9CiPbkSg3CZ6wxyysLxFSTFuHo53iVSYCgJ3tk2nq
nfpTOUFSYOpR9soAyfd5KNMLsUqCAREiDWun+ehkRLB7vz6sx9/hrhihvhklmtzg
7pGY1walzQK7UNFc6/GKPEo3ojIkVXh36CgCpp8Z1yWSo1iJQOM4yw18mstmM0/s
nKk/QgFuYbX5SJAyQlMwgiO4PFvNxhlNb35dtuD8F+u8jI7hShPaF15yE9eZbQaF
3rGgKcSY1waFgBC/qY/uaNDeu3N3/HVap9m+p2ewFIFwSAjySun8PJdHvYFl0Z4M
Btlr/fSQxJDUfyaK95bnKhULYCiqy6vrjYeg8D9yw0zONQLzK6R+JmWC7KowQ9iN
C6BSoj699HtU/yrwXsgUaBQ8ffwtGZzkc2Z6922pvbyooCmCFx86vy9sUHuGHPOt
2n/Jx0U5feWZXZ5ODCArcGpXwOOX0c/2qD38FbbfUrUzA3iHVXfo6fi7fVRZdrKv
C4UdyFXDDX3kSOsHdh8/jrnVzbsyFKR2c2zefjz0L3BFeB9XteYzwBSI83rKeSWB
Ke8UtbYpeEdJ5Nlrpt6g/TWexnB+uKXp7tnvIO4RE0KXTCFXchI85lsFJkuA/rlV
FH0bWjSYDS4OzZWOf92FybxTxUN10UudJ97cXwlnOPYVtGPLnMAwIa+71wgcdx4x
vrKRGgnT/IJVKG6QIJOaPnfmCEmUOO8KsUD+BuaYhkIYvkOZv/UQiRh2v+CEG0WU
+v8M9+GtpruB3z/WNKe+TC7s7AIUDqgdc7r2t20o80kMUT1SOIAhZg3+F1kV/c7+
dG8zLkCCpUKIT0h4IlN649J48zvyjKzBjIFArMEzn87N22l12Klaesg5ezsniWB0

//pragma protect end_data_block
//pragma protect digest_block
J222tTuKAQ7xle+xMbEyBcrpJmw=
//pragma protect end_digest_block
//pragma protect end_protected
