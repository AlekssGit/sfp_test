`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
dklCFk5RkbXppeUy+h5XH0rP0dtmmTuBOsdGRd4pnjJ8+Mvb+xVn64FZr1Gj/wNk
JkPS/4xKXgPf7j6ZebrGIOen5Q65RmzToF3Pf/J9Mhfe+T8XRl8rG64RX6d1zaZ+
PZ8xvR2BaFEikRZG1r3FdNhzQxjSkyNnXJGEpgCjyZ4=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 5168), data_block
MSokSYg5yKHHq1nyIQcmF/E/gxxBuImUdAzPrsoOjx+b60eEqajFCSQ6KOIQoBt7
tH3V3rbnlrunP3ydBnzjHUqbmXCJkO80P92Re4/LuyZ/el7axZ1bzXaaN3J+58Jc
x2EasRw+aSeNYC7zxzgDbbUHULYOkk7cC0ug1XaVh2TBR+ykm9HYrBGM+7uf1nAj
hkzGlnTUWVZcz8cN4Tb0KtwpWTOeBTvBnjZfHzPp3tUEnSh9qR4bLScUqkBNJbVd
mvK4srLEwSdNsjJfCsJhnV70Cg5kiLkEt88mcfrxNMS6Eb0zgDkssIC5cGw+mHIE
5CMuqI6yrvRIbvSyPUMmRGTYcUhDymyiwbl24BpjwUin+cgH1MHCAbBkubjyQOom
miLIgMC7xz/oFQD6k6PrpZJtvR/TJRQofXKHg5zLJoOVLozefiQbfXhWmQ/d+m1a
lG79KlBCRP6BBwXCVMeXw/zAeukpOiVyUTRNveDQ30Nq/d/dL4UYu6G69enat4b+
bJv4t0EatSSm+2guPAq5S1wNko2hpsiN6TiXFBtn1wwfWDgwFEy3rKCYbg2CYBdS
z9Y1tlVC/C22jmWQNKr9zXk1XPOv0bJTt++NJ4Soi6CxkPCJJ968qaYLWFhR8OCm
dY9iZylzvlFShLgq03biRSUHUGuQRNCJdZbBKnVXpEhyv1QNo2fyRN5D2D4M5/MR
PaUfZRPC7oB4196XBO5ZvxguRvIlI0khUcWbg7Y3pDp5vUxO+esavJ4WYRocu8JL
l+BlFGhcObYg+9r650MnTq2JK4Ymw+zFYdAJhLhMTaA7mfYpgLPUTqyAYhGStA0y
mvxVuUS22tjeyFPNJIlzMyPSTQvcdxL3evmhcydif5u6Sp16ktwzxToIpKstycMm
PPZFF43jr3AloS35XfDaKNZM7nQ1UtFQZhnXb/MqfMy02CGgmuHHFBffbVFZJGhM
MvHVDDapCA5d3hPrB7GHMwJurgQYtpnDQS9/WeEXjk9gEkLETKiW9DLBxcXXDYoA
jGJSpiA7/9w2B8z5cHp+joYJvp33ilNXqquAtaUKR+DTT1CAiq60wV9IrO5X3uPG
V3DpUrURqsGu2Ve1qvlbTi7cVx8DRUneNQlV8G86f8+KnKArEg3hwFDGmtMSXj7e
k8LZRPo7E/qvG5frMbJCDoj20qudQDdWL5I/uCFKLP6VYcl4oP6xw7w59X4/NAgy
BTtmgbvbYrkuVuG3tDBKaMoFcaB4I8vxAE5MeiHw1hgw1ww9iYpacTXsg5e3UX9C
1QG7Za6lCaDarsGt43LFZhmXM3NGMM8VtFACHUI5jrPhYZuXcT1deFAqjP5NUCXN
owy2Z+mgHdoosKj0kVHqn5/MokSg5R8v1uoEuKqGqJYiJ1SmQyAxjLNRYDl6Ji2o
5IVA+8Rx/qfNgjpybaiJsaGw9PqX23qF9rgDUU7agjKgBQZYKbtmfHiot/vuAe+/
j/mbE/MzyNif/xW/Py0gdrB/8B528JqIaT3mtxoG15SCD+Hwtr9yyW+b6AMURauN
OhvQaqgN2wl3GtwbiKGkdfQhz/XXLK4ttmyWto55jdnAp+ckv4cBC/3HzRQh1d4N
b/2UEOhJNNRnkXu8W3jBoQfFSUfhRoKxz/QLI0MU5gTQk3mYuGFTkVESXvgWYfoE
IC7LE9oR+NjqwRfTOf5GbKXf/zh35T8fpNTEnseW14eoYy8kNV9xAPN2KkzgoJwc
eE40NZhQSc+/7/Usjr5BoSDvqZXm2TJ5qQyGzLODUPMYAYjEWLBCxl5M1IU0S7Tf
tRWvLrjxiiv0QUg9V1wl6jVOyGIf1HTwqRHER+RSGva6mnpQ5d7Y0XmeLS84RChp
sp6hboMJbaRLzcYX/UxxAgCJIKlXJazaRn2x6HLc9fT9WETrTu/OCmFPitjJ4q6B
0NOEGDqYGC4rCB6cAvdio3twnRc2MaVYt+d1GdI2xWjZJw5WIUbSP42HrO2owqnl
AwpjV81P22WKAx0DncqeQpy80MfdlszXh26wJ9pQ24V5JCHIGVVGBFBwa1bZNWHB
M0zrOP1RgSwFgI5un2xUWwDze9o1+QT9UvfP/WJXj0eBGghGd9dBYWaB8lHmH1JC
WOK1sB6uJj1TeLKB/m2aQxcgZ5ZkthYOGnKIw04U+79c3QYZro/VTic10rx4MAo8
U4dqn3vVdKI1r1VP13zBsKCPoczbE5TX2oNZ18MiELSndTkVB5rG9nST3HNQ9b44
oaCD5zW+vvjRKhD93Jr6XJuvrSzqqYLEQho//F5GCWNY8iaz/BjC+YrnTfvRxYn8
+hQpPN8zWHcd7HN54idlOlkTR44dnu2Q4BJ1kMBI0gTWhFfqienUSi51TueyRVkm
QPN8anrtM7PjGgSKRMcQIiml1IZdx0LyomClH87XsNYWPQXLP3oe4XvXXl4x7rmW
2mX6qLf0fiZybk1ZiFIHSg1O+flg67ttvDawc98MlJUfLfD6na09c1dkVNJePfWM
B0IRM2B3GtHJWDEOt3MuC0SAkvXEhnOxJ2dbY1P9F+czanlsSuPjfOg19QHOAI3G
8m/QX7n4ieCwjPtn92Ndkk/00b4RAZ4W7Hm5/BwX9PbTk9hmfsiJ0WkfYM7xH3Le
egrb5w+C+9UwUIO2Z9ErhbLfpCmpSARBNXuHkr3yDriA7Wxpu5QRD1tXxoemFiQO
QMbhnMZvAoDWZmlbEOqyKQPk+mnH4eosMg06GC1efj2dHoW0sf5A6TmHNruSzyeM
KgkVNS6MsDyjgVtKqwDLicWEqc/cIsi5kvIrn7Pjn7zelQMSGwCdYGyrGb9jFojk
R6PkatOO6dJsPaSp5E7WllSAHLBHgVILsml3zgEqD5tYXLZAPABLEigaboDsDuSN
+HDPJ5xhBPgyZfXgmuGPCutJ+pxNzgxM+/526HOVujh7930isvVVYcXGRRCPuUTr
F0IsC6PPHe6652SbZONiVCACUDHn3qS5HJ0vpsfgd+3/v+oqqTX0e0jXWyybj0B/
mlzD8BnJR1+tGzNUJ5siyWXEGu4XGmVznS4a3H3IZ2sIUOIJFRbvC6ODFsXuQ3A8
DN0FQ4S8DCxetkkBX1AKiwrwNuD3dIEg0TR0gp3bNFDZyWJP3+2HrX49MGlC4cy3
8X3HCiwgybFc5R1oe3KlesxR4vDR3t88qUGfK8brmnx862WX6ojU1T4sji1QyvZP
7dueC94SFbzqmcKYIn4N59xYAcM0vntMylZQT6bKwtMfFoK64laXzbQqiYxqANYl
Il4jnEQxy3FW8iWIVGx30TB6aFdTXM7+PBuw0OJMXfF0sNQvmdmneXFgyQi6S5fy
en4ZRu9yk6a/+apTYOrlsSiB+enZDiwcDkTY2iQ9TCJu8tp/qWoooj9QRdUpUJPJ
069HEgDVfzVcDP8/CEwGAtNwuqD6yUF98BrNCaIG0Fr+ocPCFP2fHKEYPYhcOc3v
2gs9SUehbpMouYSqIoHTre2pbLoJgDTZW/YYJxznOwKGIpGxR6IPhvOU4R4uKBgb
j35uuBPG4sok38pzuHDVg8+RI29HRaw29sRxDBBKswQK7NxOysWaYG/N2SI9U+Uh
wMrHr/4XfeLI1izYJnAVKypXT+XFc3C5fhpycavzY2iZ0s23DCONb0/5xRh5KLyY
L0bKc/7ptOk6KJsLN3Vr4NNJ5BfsbF5BPNEAFdQjy7Yz0Rs3NJtuKRDTVkbBZrb+
p+yZLsMsBN5/fwV/qVfvapZAAzmjxLbtDLydClVbHIs3ZuoY2fepUROsM4MEPny7
ISwYE6GFlHX69rD0apql0JOy/6T2Y4kMkrzAPdQcuzpWGuUPsCen6zWIoydEpeyh
GCM9eNesf1ChUm0uTVPPIqHPHaItOGVuVWLbN7VE+4HugN48JtJQEHZ4aOQiViO1
N/hbZyy2v9PhBqzZFpBR2RNRriuoUS3gCEU/uF1f4YVJYJ9ZljYZGXwntFjmY3Ym
szVzZSY9OCWtgTFW7cZWNQqgzxFu4VcI8XvZCW+gCRtJ2hH9UrtMO/yd9DLrrQFN
rKGY/QuBK1RPY0uxyukEwvoUdQde/c0i8PETOkFvbzaKdMeZblSq0S/7Sxn7j7Ta
s1+3fHm/q13MiavQLYgXnwOiJZrQ18pqRQGoxPBlaTSAFYsTt8Xl/YAn6SdkLhvN
Ntavmzqz+YAgUUmuNQpuYHOpbZRXRdRtiKDk2WN9/q/cQswJmC9RoUTVVukxLMS2
gAvHLUIaepf1SaP5waaMF+7JTJTtxHsA9UCbsEf/V6gwpSdvGUwIhx+ERTkfp65o
nH13GaNE2Mr5BRBv4AQp1N6ujP875bqCLghkr2LdP5Hsd4XNOq886AV8ME1QwVmc
w2UoS79gbZcdIx9V1M4+rf1i//RZyRgIJEeBLe7RVghzRKii8pPYnnQoYTXTSyty
uyp689YSH5yIvY6479U8uhfsXA1Jm6cNmCzrE2QczHdeXHMVGypXINXxBhjA1NwW
UYq0dUl2W03Bjxd/bKstdT0Iz3UFEz+Og3jzev1US4VmqMDqGZeL2n5/mI5iRPpa
tvvfESuj8LoymYis5iBku/nCqMrCnpk4h170g9EVjZ31zjGagmbEb7SAkPLD5IpZ
P7Oyuh1hvHGXOfbfkkYN5kLAXnzopm7wpXXoNN9WuUvWNiGqKm1ei5HqIK29a5RK
4Y0W+8gj6CJ00qZpiLXYGzAbVOvM16LCGlr+PeE03jg1ne0jqDn596tc5kvf7ZoY
nGI2cSmox/+uXsyQnUsxaPW0vOwyID01qTsd3eSkYmdyCTHAEo1Jn3hfh3YHLEdo
mCvIuzOW+T/RDE/JucBG4x3bS+1ysbJk0mOtYZxH5v+HhsjIghcHi9Bi+6MdNjcj
cT32mafub+SNbuhHgT+gr9FufYm/vuJtMjzdgzidOVKcTiQrRQsJUwqTYCcNI4/0
aJZ8gYc05q3oSWL+mOH0M0atKPbc4O5O2yTfEnJw8tX3iSs1bLqHXySR1F9K8Tm9
JmpmQ6fHUgPXqn4J/qL/po8KI03AxC0xkCfuj2zsybUdzS5wOt2oD/1zENFsaelV
gh+3D/pvN6sEzPoDvYVoH8CiqXe09TrRFQVO55cVDPSW/jvTv0demaIjOOBntVJS
xC79SHDB4Xvr2Z+GQ7LoADy2xmH2zBxicBPzdvaUByFF6oR375HpDIewzPcKdCCg
jWYSxguPdZiCNwwMDe6M0i/XSPYcUKrCHhbHP2Zj5NzfTecWuWF4XYM0crCGmAni
XS2y+vf6e63Qn1ce0HUYTW1IHdUFr5MBXXUphiz1cVRstpuhhn/rDU2PZ0wg+Twa
mxpyhMBXGhTBLMgfA988q9PACzKCRsCBVDmHN3kKMZn5VUVkT4eEGaJ6bElgEzXW
x4967VkdgxS/pfnW9RfHZnZRicUXXqPEEi1mqPLUwEupBU9kwLlOPnt0GBa4ckMw
PDQTWIcfEIzB1rQIkzIvzhOIlBFklAYRdk3hgR8aorfXwQUIvPIqx58e+effbK/y
SH5G7g3Bf0Ge+wwbE80Wm1qTdM/Y56hd6er6k5e8y07zNm3qAZs+t0M0XrpnOK4+
pehS4gF0cmXrGXSNu9PEAqA1ErfNQH2s3lmTrTIGZt3LDapGoXcPoTXNwfKbPiHQ
zjHrz9XTicx5yzEr2pTqaPaHl+6DP/LauxGfdXN2La4HAMlLFznWa7QLk1ucYrC5
ubbWOL5hjNxJOM07/XjDbQ4KXSsnNxD3VUzEOOgEPX7IFXVKQb8DwK0lz+NWBXff
WClJqxA7WhSgp18m/+JJ6he6K/WRZ1sfqOKhoW58TIWgd3bGsXUzvqw8urqsIjLG
Pcq2uvk4UXupvYRSMyiP5TFI5ctGrarGG0/LcCPQZPr4HmZqA754169qK8td4Yyj
W8dX6RVhQJDFGWONzbxUM6m6nQuYSf7f+YLwFUQ5O08+2c7dn/GVgC+j8fq8WjkK
AXfRv+w88v6FTtuuPoS0W7bYmT445qQ6LRnNSLzr//KBpJbGg38YTsDqjEcJA8aH
PRAcKGSRmLcAfMbUPhuTQnKgE7zA511EPvBqb9b1U5oYyiWBWqHNzP9rusBan0QE
Eh6/Zx+lp0P0kmAlzWgTfdZiEYkEHmL0IYFM+VRsJun/AFIOJe+HwZE3dXtzoil7
d3xjl47vKiLkYeIjpZbUC8JEMmBiP3zKiswZ8U98cW2IJIO1YmYhB4LYm76g0H5O
UsbJ/3pUYw7fowC2Vloh/99rbmJA4i6NCseVzJiQ32YDZ1k/zqAX91A5i/XGdiMX
/igjfIbz291XhYA7Z42xysVgupmi3MZZWjXOkRAHIVEVZFt0jXoslO3mpBZEPg1H
lFJ6Qa4qXN2gBTKJQfILe5aHARn58DeoTQQiz17c/pClA24BmisQYsyjWDH0ZVDg
ewftnXJkxk562VzTA2UbYd+RPPRL8xsgkbN+F+xpCwmlVnsRfkEFqWGtXSDv24Q1
HLZKMDMhvVIU2HTAVBySTQxvOnYV0kGfCkiE5ShjlcyRNtqf0ldbpPNRIXRCVegG
pzNyOppih6aG6ws6lSDaeVleqXvPN8te8PESIrhB+tJrNkFgsS2Bshsy+PAQ39hy
6y0HQFRF8PIFdTeJr8BNFFiZzybHBETvt0kusCroBJYzMh/YL5vKsn8G1cYyYBLA
LrVYolh0gW3wzW7wN67RpAP0cDLiI/7Z8VsLXxS7sxLf4YelMTw8OLkgIvX7it3g
FHRaIls7X6cPNR54wG50G67M8vYZdYBeEOVH1JRLkPSKBj/9djpiDS7vf70z3IrL
JV48Eh5wHiyNoY9TG7BIaaJJe1MoTbbO96J+YABeXET8ht22MKbkWidTXNpW9/0E
ryPhRIjsqfC7I0jIJN6n0pgIv9ocY2PviC9Cm7xXOBw=
`pragma protect end_protected
