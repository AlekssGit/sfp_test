// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
KjUYSHtQlbGckgDYXwWiPq2v2OgZrXRc4N4/ZZSnMhnEzqBv46aVtLnS1I/bAcrO
b5HaXrw2zud/c1RjlgKhcdaNzYLwu5yCnNJCItF+zQx523HeAEfyj5XZM+JRRQZA
tJfNdn2GNPTclLjMuGJ4n0Wd3JVNGBGHUHx61Gtli5yrmn0s91wlaA==
//pragma protect end_key_block
//pragma protect digest_block
LNuyozFlI5jbLPlOOeqo8egKVDE=
//pragma protect end_digest_block
//pragma protect data_block
0EIwdwsBFEkjWGhvAeEpuGJ/su7+Iwx5njpNW0+TuAElyx9st6VR91giCXQUqZqQ
dOYxbzM3Frb5crak53Wvpu+kGI81qLnYZi3tCX0XUAoazyE66Gf0cv3v2p+vSsqb
NFA87HG4YpuDNKrgp6r6HbzBTUBmV+kfT5oyvc7AlfV1t8x8uVrNrxJU+Et++laH
L30OY+94xzBEROO89Sbpzt9NtkEaMTABw7H9x1T4VTQE16cCB/lktFd95fEsMQgX
/WrPXl1/ogs1y/VFcZVPaa2qaOC840mzyqn5JVmtabdrARt8UuefkjhIQJGie0l/
RSWb8TBdCE0zzybIi114TmESQ5HnSyKaUZlFL50QZ+wOZLzqUT+TXaEnbi3zEYEk
Q1J/zFkrAjr6pxMipYM2+wE6xb8OaYhETPlQThhqPyL4/SIkgCdCUtnteu3E3K/q
dEPCXncq49xT225LvwBp3ukaqGbeA6tw5tR4z29BNt3ZxPhzmsd97EMVwYli5a9x
TdG8HZ6ACteJpZyFLilbmHJDTAs9HnOfg4sRF369yeNJsrkppd4LH5RnyWtTD7hV
SoZHH9Rtet4sE/WJkwFnmK8yUhd34S0agYOH7cLSXzQCsrHMJvU+E9QEtwq0RzbF
iDdZ2xX6hZg08hwjHez/pSlY0KokHPr1MLkBouF+dRbC9O6fEZG/kai0Sa4wiMb6
cNEpDuKKm4soNjQS4Xb6dF3JTJMwsiqqg8EWFxBNkBsVusts4rEfTFYE2jFqqRMa
gTfNECiq5DLN82bTerWYqZSu2D81HENMOnsZ8qgxnzLQvN0hoSKx8p9E0yVoTXAU
py2dXoZL7UC8ZoImXr7j3NUdcrxoL6aVmx5bQktzT4RouA0vUP0evYlqSZ53C7Pt
chIt9Whkt0c8/pnIPOCgwOG0D3R8F2kHqWNIZn0v10gArlZaKuE89/i5VSwlUoQH
S1lyd4RPcs/uJRZ9XEX93Jcwfgx0y/bS+uGJdYcNZTp04JYFDu04UkhY2mQOgDEf
wWnrvZcOY2+cE1GlkklIbdHyTedPSL+G7HcofqGG5guiBa+DDvHlZePmplSc1aAp
WorE6XFBJeNGSPhH6BpZrFDpQzcUnRBHetA1LCr01feyCO6nJj6Wdk+oAayvNhxj
NFrpEQ7ObrdBCAW0HKezGb9ePFF2+md0ctGe4V5UxTvLmyjR1o4Udj1TnIrPKRjL
SS1LQjRuRXiMo3DpDSEybWJ2svFzRunzr52AsoHju6Jgsg8n9xQSuisSOMiP7vhx
OKsIF3Td2hdba9OFKvO2Bbdtrzgq3fkKUekAMQz+sw8kiTScDmWE58sDR9h9nmWE
a2LFiPeXgEhzJPEAcUayLmVv3rmrQQty8xRl/NzfysJDDlSSXIs6Dk1tc5QwHk9x
Xaxacu12XL9J6dEep6AZuS/1qYCLRlCYX4JMAky8NwpBY2fOlXJPoHM9BTdv+z4F
Y+zQM6REqTXVJTE/lmLGH4K4CnKPSlAeOSLIh9qmTra8GdWMA8R0ACN+0qus4HHf
vwtlhRLlOfBZOPOIXJ3AzOfDTh6a8hikbD7Zu9h5wOQOyfAZV5gqQq95XQSuIegn
0Yzca0GJ3AmpCV+oM+l//H8W0dSs/MWr1om3BRN66fGHMjHOaCZHe5zxOk5vdQQr
KPctsLnfhtsH3nbQlzsE8YQ1nru8XmqSCZt1DwSkZ5AWLeHxsGvvAoUZSCFXTyMY
3ICMRv3CbhV/+CnwN7nOdWXT5/l305K3lOoYlfZkU6FLpwM4/bbIEEgmSuJ2fn+O
MsAzdG/ef9TQ+hnaIEU5XuQegjFtqHZsigH11JWKHVqlL1/YFb2JA2QNLBwmP2CD
AXdRiuo/vGy6+5+O/xPh6a0i1cDkGP7a3rIjWXrsU179Tf+KIEOjGaQPVFo9nvJp
in3aSPdTmK0d3vkG6T4+ZtFPrPdImswkFrRSRoqo76pIZ2rVyU2PzyNBNJYUJkBt
mJso9r+1ddRLCHxoDCWHvK36Q36Vz9Hzq3pLMpBw4aWtlLNO7o7U2iSjroLYpJia
hMZVm5cGsmBO8KrF4JxyxABip/H+Xq+8CQ+VuWzL3TXkQggGPkz/QFINyWbN0Jcs
m0iKDFehC5+MOaVlCgy+VbcW07B2YpRVoIn9yzlad7WseAETF46PFOFZ71BsBoUH
PVhpFTyN0KUDSdOdO6lPttlA6iLSWxjbaySF3l/mRg2lrHRHZGDwHJ4dvBFZANUb
/2uvacl8ttLchJZifjtI+MvDddbcWIaF+TQes8p7ixNsU6iBQ01TiUxgEZuRcciG
n81EAMIBG/x1WVa9ufin2W7wC5j+L49i1cdgwYW2HowoZNZLL8ww3nOynjWyyndY
7abhGqk2ldKAzlgxl2kCEy6+kK4cDt8m856FHxXjvJfvU0iVo8/vtcOjSkRcMPuW
2ReOXsnfcdMqcnUx0HJrOm3xAJH98X0k7TUMo3HpdslYw01CpeqB83ZLh5qJ5Y8i
B2Cexho5KmpgC9frl3XCtZDRXeAB6qUDOiirZx2w7ikGJkXNS/61Ud7m2DNhDDC+
ii5PLMr6cXx4/z9SuM/oTRNBGzPBY+L+BTvsp0MEFgfBMKSMxc7TY3OjFKrifxrt
qH+hGYVEobxK8mMcClp7xG0/ZNSbG9WXQhhQ8jTU1+40LEDr8JrdKNYLEiImYCBz
dTzWrBbwKXhmmHTlbBZMTcicZ+8CDpLHLLuTdKYONxq1BkXEow0EDAHg1JU14Ss5
s9yJtRcrwbTZs0Su5oV6uf9ZYrbS6GfIEjxhR9/ZELWxSmFAkjsp+GEU/JEIR9hS
l6B++E/EEV29sQYE5T+YGcQvkHp+d9znX3FuYAG1GQH0Ou0qkFRKxYZ3IBJaGmdR
4YmBRnJECF4nVwjO4I6+UFi9NhD2LnnMKIIWavW1l3zRg7IlPq1d13xyFW5QK7+c
NVptc+/RVp+VgtNI//TAPz7apry0V9lgkvl27dRmmeZ6Kj2CGMEiw+nNftLgXKQe
dOosBBbmjPD+l7vnaRO36fBucIw7urlhzr99Us8xoPLkagfKkVS9WF/Qlx9fce5Y
EeLPEyMOhlbe4KkP4Vnfd6dP7lIJIUHbvBJX+qxEa3BatHt+iRKK31SjS2ecatxX
PTx5oFD3M2kJtJRLwBV0Z5lYcndvcxHEflGw77rRubqDljGoy8jtadznfGEF65WH
tl8rGuqt33woNYxLLzFAeuuCMtPEdX/XMLHnY/avB90KSlGGg5eLdKzRtwWKcy2j
4akGI5DLN4PCWeZgfp8RgfeApT/mD+6G3ulBFl5ZKOvwSb9PFacnDQ3cWZvwt0Ty
Dw+QVyCSENMH3WUyczOzx/Q8juUifAr16nRfWyeSgvOFVGVCrdekByrcXyD6KtgQ
3UtmKWy7ClhO8s2IvhPZnFRZyAMUKv6ptS2rkBncNbaY5JeMGyvJFzmhUNADB5KN
+RBStd9Nr6PfMhpZbVNS+E01icoPNg4joo4thOcpAKKuxa6WbHAx3xSl3OAyMc9i
BDhgy4eU8x8dr7wHRcIyy93SjXk//V/Rv+vjsjUKSIQt60F8/AfNAwRq0nQnrA/0
3NF1HieusSwGklt/gPp20zGFjf/xaBz760pfe1LOOmbbwtJEkPQb4Ql5/fp4kLX9
TrKymRsgEfYKLw+Qg5crjHkALqTWpVaWz0BY7zeU/vH4Z8xTBIrPatkw8IeRu5JF
a9rQssx43kLAuCEIXS5iO5xsw7oBodWbH9ad0oQzan3m/kJoYfDeZJNzn/zNQEwF
LFmGyMgM7P6045clUMEDsCBzd4i/AGvE39VCdCfTLy1r9oClVGfEYQXYU3MsuY9D
IKvY8UrDfMFylcXU5B//o5TkpnBcou4l4HbaGTZf6P+LG1kbPE5bWg5haGhI/LdJ
T0pdolV7CNRrCmQgpZc9Pdi1DNGzXUd3Px91oY4Jc2LJTGs5HXgGkdxoEiHKW1XE
q1c5BeAmgTri0x2xsxXwV1EcD//ZACoyYeS8TP97vVYl5APkvlAFAvZDyCeewY0B
kbiN2gEl5/ECjOBEFCmvJrARd4CGtbdIFtWYcN/nDhof8PFJfgM2GVWCaudFPB4C
AocJpfC1Gc02Qewx6sF4jrtB6tCLvbanqkSlieLjUnzdojexkvr1+Wij4R+V68w/
nfEGvpMvV83wt0tTPqGDW2pSQ4IUukPzhmdpQh570pFYoNJM4EUglNJlgO4vISsV
33N6b/zvd2J+6RenRNPA/UDV84rVjCAE/zuke3IgQXY4/7YkM13a/EoKKuLpYJ7A
f+y/FgOlXeLsTHZnCx0ngczAKz9ngQUIyEPmq7t/jDBqQgEUM/h1zzFNL1BEY8Gy
+X47MGU5LqZ1wD5UNQDf91QLayFWeBQUDFoLMCwn18D6zRksCicDfMQeQ+YqxxZa
eaFfN2hnjfJncvm72Ry77jndt7iwvhbS0I+9ZFhM9ccfCg3S5WY9QMsanXOEh+MW
gGon4V7E/HU816SHmjPHun4U7sty6xOx56Af2BouYSearlsTHjLG6bsi8kDvwktR
F0vZ1bRSCVrBBzZZx2i9pH9Bk5QhEDCPzI2etm3QhzAAmZV4CQEDmPA8jwj6YdiC
EOwnXZto2XL4Nr5DfLwx3+G/h4M9xhCnx5nn6fmv6sgQfCEx3A/OmcNFziR/NylF
F0JZLMmMJ8YgEVKNzYUAGr6MyINf+SdOOYOwdXxaAMvuaZZdOaCud4BLSgMB7LBd
tVkz7sZnBbIi3iscNaIhUd9AYwEiAjWz1k0Mr7QyuHn4a+nhK5ZgYl36D8LGTsMs
WkiSGO6Nk4Kin7d2FLByAH/iAlMRrEHglH8J+PWxaE9qKiIWjUQlE6UKbn9+mpCF
e+0h7YtJYh3FDhEg/WropmgeTfdDdaijLoaslGObuEls0RcLNv9sVo1IzQBG66II
E/+fWO0/RQNLzINxBBdaCja2KjDIO2aUk7Gm1f7/lxkrl36tfBEnL6L84VUCAw6Z
ybjy/s6PYGKbF/wKy6ZslI3rG4AwRRKCDU4kqS7tXBaUdWvwZmqg7M+fAy1Co6N3
3fGxqcvtXPE1amsbX2/Y1ebCYxD/NvtQ3iFutaB32u/5sZoa0oiSv/IBAR+Q2CzL
nxJF9uYr02SivpCyXaLT3/SFKDbzzyd7J4DPFETBexV9oa+XvNWFlJuM+vnPNw3T
26V7Mzdi0avrP4EOob4wLQHyJluAmEp8IpbAiLqkGgqTg78GNHMLioGDX1EFs9Oo
WRCHEDe/wlVH3SY8NPpgzXBKSoFbdIQRNnyu1T/PBBNYP1kiovoATmlxE1y30l0E
SKtTU5lNZewhTMvqtdw1ii/suF1bX52QM6kOS7nCHJmbTMDVyqJIO9ZlxELPJVK2
BpA2+QT+KYcMGAlsJ2M/No6ofu1uUC0GlTWsyg6FozzE0yqJuPT32wt9L9O9Nug3
efvR7XxzBXwagbhCTBU6f2M5A9vv0+DSuDTHzxu8xBPDqkcfOOtbkfkPE0CJXzeM
X7CDDuWnbZUIwOVBkwTh6TkDzDoWUjY57x/LECWwAygn5DUDIJbeBURxu9Od3RGz
PqoCkHBeoiJdYSaHxzVuLad6PPRxgqV+0OAET4KEVrVHFpfxLVw6TD8VpyPU9Yrr
xlHmQDDJ/c9ZOLJjGkRTPMpnh/9ZiUl0gMM/RCD35ujbbbWu9t1IKeHA/5gGfJho
brNsgMOXVPPE2q/bGJDaEO/7cQjm7Y69zuyq4tyG6GOrINb/ysEuADtDHJIw7JRN
B5qy5xFGioUOwwZVE2yKmCmLVcjk5P9o+oef5DdskRfbLIpdXSImDETje230u627
PwNKhwt6Ktk91eFPYXHc3FwkSs5RO1E9PoyQ/qMk8cMZ7hIppvgl3f0UeejP6dSt
hp3t1vGTqi6biGM3WSLbiQcWq+VqN/mXTytBe0MPBUj2v1qBoa43IMHNMs1WfpSM
p3OVjPQ1t+HSMZL6cXU8BAyZ5o5Om1rMbS9cFqrZ4yk1Cv0yWr7WG3UNSSwPsJlC
psHzkIBSknJsd6TsszB+DGNnJ/N89GzmF9L+BaX6m3D+WCR1bDJoQzlKPsgrOtO1
rsatLglMlps6POFyUyK9zZ9nMqAC9t4f0MZyxEqs+CiIbQbuEU+hInEVufW56Oiv
b7iZSYV9MtLQQQXOsSIZ8FTrtSRxv8puZV6tRcR7uGbflGYBVP783YuKPCf2LxPI
fGFjkT/54BJkeYeBmRCANtNgCTduH4CC7+IEjAGQLxuYawVhePMc/ojJVxO2jHMA
xKDz4vOhwcTLbj4V9WV2018we2bMZ0bibYymrvtxq+PopLQjD+DT81CZtfEdw7GG
NhXVAu+ARBo7qlE3YBbOqbAKz0yFR76TDMXUQ3aIxl/YtBt4YyNwf9EVoh66KlZ8
PczK62Nn5LzK3dSmyL8kZL/bXWO/qkZl/SZ6EKxGg/b1SOftvVus9zIcPpWSDcN5
Bpw9dmLrUh750vz1aLeQCltQ0/PUzkefV3kkSC48v5aGuhHttQ/UTXNWN0cGlC10
TbPKlcQfCquQ2Cg3cd7NKpnahBovLWvZtD/Ndoli7KSPHhsIUl4VTWPoA06fK5ct
vqVRgfGyqMTa5Vna4VHWYGDnmyJvWt0TCsqgz56RIPpEy51Wg4ARzFFJ8AdDlDG5
a4zUOvYP492XV3bvLkETQPY9TUYCkWp98u+H7N6qNG/2LNpIiOn/o/OCqxWHxWLx
73kpEYnFqvgwCQH+4ODkrPFmx5rEkSYNwbKwUS6jl5+Npu6VKXESA2Nl/SvSEmBG
Z/+YOMuSmTHiGiTad2ER6sap0EJbPCO387p54KQ9dxHbOQOOk9d72GxH6eAfczd1
1qzeyoe5jpxP8+lC07s08LZcZunJ99lODNCF6AKC7GsXstsR6dIXpNij4/fw6qZk
vSIMPoFGeoTxdBN2U84tMQZQYc1i1XpEnfvjMYElTJ2HJHbJyUBmuqw72tEfP+qu
YYMAxC7ep+AtC59dFUkRCxueReP0LEq+4giQtxCU43D2+KZp9gYaScD+Eg9YfB/s
rOXKT0HuGgAveXrNHUy3RfFrWe8lq61mopGaIwNXR/PFnBGQTtwMf0lQH+dFrVHs
KLqz31Il0BlvdWosBrz+g/iVX4dkbRvr7n4VgRr8qopAi/fFZpfGALGmSNohBJBW
ACQ9qXQxPGQJSOp2QPOS0hVccx5zH8KDnZ9iA7za9daM6c6q3SKPXfjrXzcFHPOv
9IHKN8X8l+IQWf8Auw65Rkj+S9G4G+9R/owfup4tcDZEAJsWxOtsKSe/qsIL0twD
DeJxiYbyItktylWbS3AP7Q4/oJamUxFD5QHuCINq5BZI7kNdadi6eMokTdExZHGG
VRbqHiCXOJRhDadlmI1PB8Odmn3u9S2y3A3dwJC03T+We6gUv2pxU4unKteQZIHP
Lndgwcpi9Ob1Z9HO7ZKcvxvxLrlE4NGhHKc9NPQiSurqAcPS3b06GAzUTE63m6a7
L0yd9i6DFfrhszz7cHUbsBzJAnPvRrP2oL/8Z7iBaeOWqhtYjYJ3Ae+Oks7R0oV2
MM2FQHSqq5g/qVu2UR6hjWUiD10oexRsCka/w09rI3DaEzOZsVr8+e8OYYJnJGGL
ygvAOIRhDTvx7higaTkplv3nAL4VpQ7WoaXwsri6lvVaGRyQtXYLgGBe0AOFO6/V
81O9SI16fjmkCnfAOZfXid8f3sXrXV7fQvr5TSoS/KZOhFwQVPoY1+aha5Hfx7rk
HAXT7X668JdvUk/k2O97JOeDnrOHhe7XKgLYP5yWWqVFZda6EcwqhEEer0RyB65m
m5KOPCUUjG/o1gWlP5Sc21pObgvji7P6qXSYRE79p7dCKdYgm37mofVbgkB8Ohjf
HyHrXo8EHzOSphkyhh1gZrlp8EXOP6iWBzzyFnCdmO4x/SiZI7ZTUtGFvCGxMOdb
dylPVjO9S7XoLZAZPGaQye5uCvOjx947hEpIa1ZUmtQr2g5O7r5X+EHK+YRK4Col
ld1TENEfkYIPL0C3MHFDcj0wsMSV5WpcNnYOytuTCgBrbbONA9sWEUfjf2gv5Cmv
+d8zu/nOlKlpZAFJhzJMScBgzXIMGLPtELBdYSUF99cz6DvB+L+t5uXTUkqkttZN
4UVeZkoPzhkDegzMDGa7/KJ1p6jAnAhgeMA/yzb1ZAbKAlnd2qmfHkzU0vSlR/4o
t/hXS0ontfFx8stLcprKcA+pGtC3Ty9AZcIoQQvPNf7csv9wqK6gOKrDo6OP0KrY
4xCy8U3FQ72Adc1llMcN+LshG2NeGYeam/gXYavE08x4f9mLMo0CNgIgYqnpDomD
JbTDAMj/AOGeT72ud1/kwos8dBl75eflnd8O5cSU7tIOFEJDr6PopoRsTQv+4eMw
1/kHwV1G8t5VV4esLcl54knMSqdCltepKObe4uMHSqxHkd7DFbiIl+gIdaTk5dV3
ZL6/nUNCt/6ndItxGByU6LlxbDLCWRGz4osiBX39K8yL4I1SDyVHPRh+sbr9a3l6
VYeAS7porxQ0UGIP+264Cc4trrLfLnIC26CG6mieCttgace8fScemNVbKABmacrz
mRorNVqvhUnzHPLrYYZJmlHDhgGI+XCQeHKdsQ29QTE0haFMReK8loQbXmsPuOmQ
KHvzK6vtry8XHeV+TpteYTnxUQdVGZ3eFaT3RfpbkfKYMEHUYynRWwP041xYzgNW
sOR4L7gxAyn/YIlLvVJG7x9xnokyEoYgPOy+GTzILeSQlVQ6cZbSwDR1kVv1sg42
BOlf1aaIfCLUVx2oUiDREGMvjGGYt/3eYWeUXDWW+HLrzw4nz66tgnwscCAZ3yaG
tuWA4tZYDfuPheK++1zD/CW4oMRmykzWx8UsOMQZ7dxqyCy/6MIhOpkIS5ejBIsk
ICer1lPVnd1UgeRvhjelLazFaYngL0OlI9hkHKR3FQYWCYhC4A2yyRIfaIwpelBD
lS6LEuF7IGjjx/0G2e439wKqzvIx/eFBzxfACJ+8/ZuWJBEgqUBMK+4rVfTpu8U7
AB7ZaLVf+zrImZa8bOde33oSIrZYH4SWBRnKh7SLY9ZlLRKeTCpUut7nvNRPwGcB
JKZJdg1ILAazohxIVeI0ZDFFW1wq4FWJ6czGNNYUUO/MJyBh5Q1nJBwEI+6HbU/D
GLzkTz01be76qRWITYVAup+XDcwyMs25jK++CdfweGzbj6VKwJ8i8nJLtPxe3db4
4ij71DTGpQSHC9yNuNjUYanzTG3y6flICRhgJX/POUplhl6mt3KavdE1w/nsvUa3
f0nWfdFTdBbtEzJiWWFr5VIjY0fOVd+DvHyJFU53JBRKna7j2r1hNfub1Wcp/dAy
sWwhtUUiwcfYE/IcUO/j1OGSO/z6THuftwfAsu+YbGjLsalmWGltHtikTYhkodmg
YE0Gqybtux8fnK2ljxu7A6Ooz8GJDORxAsjQFgV2VYFBR3bPzfsObJLpR/dv936W
+CHj3Yq2cc5EsdfwDrimYLIqicYqr3NOIj9E+PzIgeVzPfEYOc6JL5su+hFCOC0j
OEtQog0nNF2NISF2/IPbXtjMQ8LlggJGoDSqLx3ygw7f0HosIUSx5tosBlbua+zq
zsCL4//AzHyacnin6J7w7OxDHmLFeprxjOc2k7jGxtrQPohjAtFfRZ+vdDgJq9KN
M5HpTjhxynSeWeXeCN3rsCS2OcXgX3O3iF/xHRWJ8eXW/odseTnH4dKLbshumuxA
0a5VfiE7z2BDrQnWVbxyMLPFKvqCD0vyMdsv4zDQEQEvKznwNuuWDpLeQyMmcmof
eCoYtqNA7BYjiWD3bxfwOk6n/lfYCvOvGOw/E1qgXJvc82wPOSb9+NbzuLN4RLfQ
ArVEWcPzYKPHg+sD0O2Sy0uAA/uNHFVXYgswTXRDmWvx0fW7QZRtrA3Ub1JtPCU5
6vbwfz7PltzCwuE78uZ9fBzjWJKHf+RZh55V2Ox7LMcAY7YnfRpsSAlG1UoCQ++U
1Ss7uD1BBsrX06Tt8r7fIfXrXYJs1PeHdMJNJ4BZ2yV3hxR+s+ZCMJb8XflZNWdG
pnMdi58/4XzfKZL7KUXD4qFO1N4MYEo+nIPJIPtbsI8Pw1LKyIV5SqJF7LJsztXx
AWE/wuEmSO7/6bhvCSjTFF5w7FVvc0GlPGavCeyTGyQhVDAdigxxZ+KWLc87DCGN
/6tWdLJ1Zx6Z30SORg4ybPD6JcHBmkmi+E5vqxpwk70kTDmB39wzmEJf24OBSHGX
r6+F2oZTEvhOqENOzpd7bK0YsZtkxlyqeJ6ojr7rDvV2VKjivwcaGoo9sZbEkkmK
P4GJNftfWITtOnCvE1A5UNFA1ZkPoqFwPcEfYjuNWl+xL/D9mCP5H/f1L5uTtMGY
pf5XlNfLxJTg9Mmj1qM4cNR5Z/ZBIkYDK7OpGvHZRnZGg1uDdkUbES/VGbO50kKj
S6o2C0Rvy5Kw3M8IonW2yoGFKH5GPreiuNJ8euHDL8hLvLfhh4wuMfj0GCo5oLOm
t2XdA7KdADqnpmKBvB98EswAMn8TLD4t4Y8UVXqF4p0fnFc+SQK5OWO1TeU3qQ4n
gk582ly+61O+Z64f4piKcD5b9eqTDuHD/8Yam7uNTrJ0d4cJL+jxKfoedjFp50LQ
ANAlqD8lLXBhBVKjzfyks0s2wkKd5IVnCJmgvswFdQCba14kU0O0SkE0Vj08/FC/
06OVhjqKc603xIJ50YcgDx9mz7Q/EkmvEIbTCw3qflXXJLd+5PXZxayYpFWCng3c
J4OuJ5xBFT8xFFs7PCiHBoawQJOzhFEEbfXDx52mDjCeYgDJKImrPPg1ImKkplu+
0ZAJfLk6quRM1z6ENuMhiS2hfSm+q1+D6/s04IOC6g3JNSvGIt2dsAG1SqdSk7u4
fuvIUCjlH4ebriad6JJTgqKdhiJnOK1/gYQshdamojIv8E993iW1WZK9Ew74qzLh
NNRVAkz5+OhmhK9COiv3f/jJcNCbQgysaQPK08/2hCsV7ZkDV6U/Ll5VALoo2qAw
j0e5UXqseYCyCRxyBSAQx7a9/r35ZyW7H/B65WmqWb+kHD3urFc8H0ynL5LvLwC7
6VHs97+fu9pHQo9PJX0YeJoykk0u1Wi9R5SZ1VcutgiauA4H7xE024zoZUKdyR3C
zAgmTgzsnYzXCmjCCUQlSoKTfkW8o7SaumLMC4+NqYTR4x7n06HlRcr1zrbuTA3F
4mFaXXBZZEx7RJ1pCBCOB7UoRRCxZ6NOxDNIcowdSC6q8BJL62GJPvhOBqxX0NZ7
5tEkRrZtKdP5C0soa3WaNk9C5++nuDpJTF9huhizjSYxKWa573bzXeowB5i/ATp8
TP/ipaHNMOojBevWU0Pc+vhPo2iyAfWqx+cHEzHp4Njn+TK7gX4Eh3uMqBEYUZ/B
S2Fi2aRilmWb5luZvIZGhXMC8/+i0k+pQnA//C+a7mCNKpZI2ls6/x4MXkJ4163Y
Apaya1OgxanfRS4krMlqtLenYZ0BhFq5kKuYsRtXdV0DFxTk4cNxSi88OixdvbWQ
JUovjdI4+tednL8mhX2b2oJzW11SA8EnHvcHfi/d/it27sXF0qlICxXg5jd7HZLo
KzkjHdjoYmw1Yb8FhpCCQQYg76GbU33ELmPCzqTQ9+CKNNE8YrtlIy2lNoo0n79e
vKdDSBgYWGq0LDzacVljX5qgK9jiMtnzRRWJm71tajEgQKwZ2OmaY1o08IHufLv5
UP45n3zPlqF5Dnf7nEys/G8Y1PU6oWCKZ/A/hPbi/NDKHiQk2Z0nkgjqqeFteP36
095/OPByROXLw9l4brUheZC+ka0YJLCduMUM2Led8BIIBVUAXu/DkC3UJgyWS1KA
aA9mNyYqVk3auR1mlj91dokp1kh5+q6rFqwqF3LxvkzLldkTR8nr55WiqcDMYIjB
rrwUvVMuqLb+OElw6J/WYKVg/e3o5yA7gp4AbUhXeqjeGfLTcQNomw3HRrKmZYWy
y1WSN3TfvTs1GcBoWiwVhDPQLexPjGb9HFKaKTK9FKu24CwO2RwDYp93yavFtIR+
I26YrJHoEL57G/aLMJks7oK036QhG9hSyntbmgI9nm112B5rCISyN0k4RqBRBAdr
NZWuk0uMv6O+B3k43ko+iiNit5hJQ49uu9rHjcoQg9p/FtZJ81cnD+QhA6sYsOwm
R50c/ELl0bdqNvN0yCuE5z8nNNvdhc6YYMiVdFtsoHTya8n7VsyNnxvKxhBtgNMQ
OX/YO5jvCAmJVKCHbbKk4/Ux2RDr4ODYv5b0LvOzqJZUzjVTiVcOYjcnLcP/YgU8
cyU0X0IfcBIUg+53KoVbaNy0olUX7Gj9WiUxc1PC6wXwKZZ5PoI23Ezt3eVI5FL/
ze613GUFza69GoxLGKikNFeZ55ypK4OQXk4hmNiksA5yAeIqHTun45Hghv6JYToE
MzGT2q0UmM9URdgk6iY3+jTTAtk0rew9ZBbWZmNRiGybXjoV/cxmGTNJLSBl6uat
xGUJCSA0j/ex7A02wT2AtK1nnzFleY8FGH5qk5NoN6trRLzryuDS/JOIx6XOkoab
r7MUPf6Pb/h47OV9bSCu3Tw3ofcV9vM7euqbWOKqFNrYjeKiXTAjaCPjC7DX4Lkd
6rojPbbp1EdpY2XNF6dh8wPua8timlyP9B3mNeOkTe3hL9twS08Yl4Wgs5riEKiG
o9jMwjOMsMb7PC0CKcrjMTipbW+1N4AXbtJMuSWt/2FziXg4YYGiPGKvDys887Pb
ed3tX/wvJFQ8Hrak9WpnLEy26dL12JuvCLgVE0fYlPQ7UGuUQQBbYFSzzYcXvcRg
xbE6ceeCo5i6oD0JLLHJm2top1JFiFWfa9BPa9EAVruFd+KJujRLUE0WDtHF8WsT
dYzzHuzvLTtL+RdNswLQDy026blTWE4ZlIU8YPDq21wn98JHQyGpiiiSCepZcWi1
3CL/GkwDsNWYTLfFJWv8F75cvgNd1YewhFs52qb/gOmWcPjE3QyxxPiCeKxgv++v
5BIUvQFO++l9HkU6jI2klmeEDjYvmmBaf/ign4inToZB8fctovU821vOWcx9UifQ
pi4YGqJ1cyiae2IyxnruZWTiFXgoP+/vL733a4tOm8UsANHlGCmKEnDfU4EX9TgB
hA3IQL3O5nn0FaSth6JSGs42ZNM/3Cr5jAEeIoH0ZQCiNNnLspoFn8HPjLf+5i4L
jB1rSKMzItM0xTC8fm9cP6CzYjDOQxUZs70baoOJ3AgjKqIQY9k/RWloQfzx9JJv
T5g6cFOwrlXLlzBl4/IbxkuhuHF3E0sqmqwdZ1YfywW8lxrAKWeBMd44jAT2D8om
uYZryvQAF0JiAHjXatukTBqUV/D7MKChK4K1soONg8w7oQk53LGKoWvbLI3tVS5j
Z+fKOtosckgpjZjnnpROplAfATUokePgYAfM9CpH5k0SCe4yHqyju72nr8opZ6KP
CV5TOvOrANr60hsGyDZ3h59IRgAOR3P3vjMkj/UZAfqGNbs/DiIjuUSApcOzBGKI
NBHlCDm/4OkxqhN01Ca2e5LiY4N4723oQueym128z4pGm+P/h3oINKx9rWwlIJp7
XGHCWofuSkyf4Rin9JIlU7XTbJifJQIC6N24wVNAhFFbuXGyjR0wsO+H9gZYA7/3
cvgoPB8hkAPWwtNFeVMNHANBvWiwT/lfZC/RvzrylEpZSMQ3KkcjLzQ/6TSN4jsw
DjnWdZINIAYcD+SQQ6s0nZFDbtDhutHoOZKSY9vsFkaAJMlxMTDfZKPeU/9mHBVh
TD0xBkBmDZLFhxcJCB2JrICWyc3gXTaP/kFVQeSIFBkrCWVsluOvz9wtAuCNMFX8
cSWin6VONMdWNij1od4UoRBO00zYA/1CO8L7T81jAb8IR+r90sZvfwA7Ndgl4nO1
gScvGvY/qy/YUb8NmWxnSG+uTIICwm18/WPLY1QfSSlz9qaHOUjGF+Q6UW+ORk09
Ixi8K1PCc77+ic3D4am9+EGh85OkbqcdXX/+suIPu+Bxy4VjfyJ5zcLA2lAVVw4h
g4jWlTQ+2BMowCDqe8YggQ+9PIX7sV4x45AH84plkSq3/6SKIy9MhBZtcW3hfQX0
5ilxp18I9tr7RH2rSgPdMqyYO7gI7G0GsHmP3s8GzXfZNaP0G06NT6RqhIgE/8gx
5XlHiA95uZfoFlRGOdaW4M4oAlEySo/XgR1SN1ZBy6r+rVqGVZgKB/Ir68yww/ks
0yKGU2zrSbns7ADq6JiSyUC+eojCJ3pIpreFFY/Y6tEJPnqGmuq96uewhnvkeArn
5MIQraT6I3U58Jkv3ZqGZQEJ6Vb3VvCUmqm4kpg9PPpBTtfe4XYYb4+hh6Vj1K0F
pXQ3w1+NCl10qYimIW0tDcDbxr44exW7Nm96Ew0cBlebZxTVgXXRTT+1gmZ7AvSt
G+bYML7gY3qEikaGjxcqA6GiLZwQQMI0S3J8asnBtX5QLpwyKbcK6BnTGH/3rtxz
91TETlh2lWydlBggTRHPeRnOKOrVF0226gwOWN3FN3MPUAx4etzD+MGMPTXWSe3f
YAISdGPUE9NfI95yNcbNqA==
//pragma protect end_data_block
//pragma protect digest_block
ns3E475MBj/Gbj9Ow/VHkixsXEw=
//pragma protect end_digest_block
//pragma protect end_protected
