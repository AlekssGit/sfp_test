// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
yRid4LRfx+L/dYuUYW4TYlGJhtW+JGHmXsTHS8l4+MtYyJwzhqDGex41+nOIAEeb
iat/5BGGQc515wuKF85N7tuobQa8rHQSZxvEw3jap9WMREVFZ8d9bk4C4fvtjVnP
9sBGkuh/OwB3n3j6ELrayqyE7lSbuo/jG7Hp5xAObkg=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 3744 )
`pragma protect data_block
GO8XLSB0YlOzbG8iF4Hdu0TyYDig9aS9u2j2GHkrfj5MjmBG+CK890ibaYMNazOz
PhHtaX2n+vJLoM8cvu20gw5xmudpA6ZEb7bYORKVDd+eTIt7XacHfJ41iNM5gJvi
AWaep3xS3++WhucRpqlAiGX14c1VKbULlpEhzZv0tLHt3DrKW/AQZRFhbzHnblrq
EOJ5SAgV+/sgDR2cqCvz5eACaeL307+reg+Vlgm22B7+LHIgJHh3OPPRlYx7CIS8
gJMzdNXgpsIJviuXeJzqXEGDSXqerUZJJF77YGRY0WHXXNuTRYFNEffULnbAmTH8
yq9WslKowCMI//o8AwT8ykrLLe6TmuxbdLEAOm8X5O1TrDvsxC2kKT5lqXQV7DHy
IPV8iOVRgC1gFBCX3qsdBhIcevyp7eSmmf6A+fIxW8IPuLVuhFAtn5VE3C9HPKIO
XigjFXAPxaOVoGq/6yAJHfiJxw2of5rEdnsTTlEN9Ad9hk+gfcty8c1/6biehceQ
2W6WfVGEv7566GxWsYRM+dno0xfLo3HMhsIKbeSBpJ1kGggpiJ1uVdhMW4wmQ4VH
tE1yi56Az2hvASNEBl98zbSD0hHLBvw1YFLfBw2RVHeLtMF3UybKIZ4rNHGOp2Ht
Smx9MVjsm/wOgCO0F3ZzLIbucDv9t4U9fMooNBCLtCoF9c3xsKEwdHRv33nxwE0i
jLksCLTGARJvUePNXXPA5RGEerhGtQr1M8htujGM/0u7tKCWiidDbngbca0kYrSX
VPWE6UPLpNsWWc9kUsCj0WIT5Tamxb2k9bw1HwTdfAygVlOJ+U3xfhwYINJirYpJ
35DnD2LTS6p3i69XCwy3c8lPYvBgulCKkMKuFJoBK3/y3rylOr9pqw/ClusdEWwh
Hg4Hf7zcBrbrz0apO7fFJjSIexIQ5e7JlUMWjLQToEWOv1gPEgS77ha3NYxDHuDU
EqIx7adeOn1ZxaJxQ9eKkHz5xeYT+3FXqHVAwTNyzmDEsuaO20jfVyq1UWnq6vgG
G9OuFKydTAoxQJ+BtKbj0ku38damLyGFghEeNYbJwHqvOZYcT35+vjM4zeJ8d7SU
HYUmBtDPOkpdleuuo2bxsbOPZ9SU4CEd3WvaM39WhuQBCSs/zBwb7IoQLdgBHzec
LIxo0zW32nHqHeiFbc3snFmc2+aXMaNlguftDP3+FJoeNUUe4YTEGSJyfDMU5xPr
9RxpR9FaZzM5DhvdwTyNxvQoRolTy8ua82j3Ml10qOt7yvIjpU3NCw95NzxTar+W
0VP0QoifyNZYpZBpjxYxJnIAC5R2l1aBl+AZJptj17Fo1uLqiuF/8q8AyNxJsicE
UB9rGFrF4FNJL4zjbcxjPM/lHBS4OFvdTh55XrM4CAUe69slHPpA9T4p5ahbW0ns
C+GCo0VsgBelITtN2JXs1I0oFvqTanfHQ8+3PDCn/CuJbYfQS70O2ev/a3ecidRV
TenUsyDPFX+PSyWUCIkwQ+UtI3TAjzz1gFOMXc+iK0Gaa1nZJN9o5sbP96RZ7sjf
oKPVNmVhxeAzlYqah3fT3fGcHdlXI911zvlmUkS+S/6Xy7D+mr7LIVX8/etWOFlt
pYaBo2OnLzY+o2yigsWxbLrTE7Cz+WammPmjBWpSdZ8mINV2L14CISvDFDGKYRSM
NRUm6CYihphrd1OAenfQy+OSu7fjO64NjFq8FeZ6advrbyZVIZ4nchoGKSmucnpM
sF0Gyt9OmrXB93LLUIqxAz9N7aVBRlVvIgrtHk5wU+nfSZH/fN9lgRFrslG6floq
INwzaVN+vCSIUj71ipckmutBiLcX3yp4haTIaeJEsbAbqVWV6r6qRqwmP3XHKd3m
d9vY3kEy2Sw0gENzCGIvpADcIiHx+r6Y3lLj1aXMM1POBmq1nHONRmpDFoRa50NL
CbYe+gf7bvp9KWkr+Hys7ChmFhSN4/vvFgsILymThIJtXklhciovCWiwES4hov/v
ZlVsmhYM032KHCM3Wwpveyp6FbMifws9eh5HDdqSy60fgLsRYUORISSGg4kHvwbr
NEji+rBBnErEG8RKawjFjk97pby/+mtV7w8qYalb+3Z/UkzS4Rtg6AosKNWrsflk
R7Y5G6wtXbm3brwyIejr1lpMgWXlocUx/ookhiE0xSiT+bOBfjjnvVtPyvmR6YTJ
Bd4M6U0m728ekAHTCwuKsKHsuM+K3NZV5TYlPsIDMh95XIqG7dmRxTNsUssBob6v
a3Ucbwtwc5QJSpxtlgyHbdJvqWWxZk/pzE7Q4GpHftaQME8sBSGnzNfK3qoGXZ2c
RV17B0x92uFpEMdefE5bm43FfYZbue6lZqwpUjCydhlZxlmO5NbXVaFlQC6WT3F1
CVur308lpQtT5nqFPFCYNejuNDsOcX61FzB6k7kkJ88OcOhsgFExJAkTyJIiXOdC
9v0KBMOcTeJw1A9D95Y+2CP7f21hp3kf8uRhfb3NwG0Hwr4aj506M8xefJn99C8/
ITKjaWKfbRAOtZVlDHEpKGOSswGPVwRhuuk3F1FsQ76WlGxNkRShPnpVG56PBUy3
av610ASTDLQZwQoT/7sws+72B5wrE/ox/MQF0tgt8IqmnacGS0aWAh4GjhWtAawe
J6rTtwwY4FNWhJZ9Jqs4s2grWzPGJf0G4de84c4Yt+SIfTrMF5o2QCmIrPDu/s4D
9yOcM/VHq8Cx3+NkWJ/CeZpX0E4c+SXoftbHHmnh6Ergnzw/AHMAYk78lQxTKX7l
QcayX4LO1xkR0Szxs/NHoEI5xabxCfnlKC2WS79xdPEU6xPSxCqk4Lhb1aBk5qYh
MSSaqFj276HTpP3wz79V5rX4ekbJ0V8NJOx4qnlK0bGjGtPrCCDhYF6YzFTokIy/
OFjfIPEku+EwU4AF09RFsHSOtgW+Zlm1zu4GKjxjDS2hVYhlRMuWmkul+8PqyKyW
71gnnpF49pKA3fagTSGEXV4B1vxkU6hHDQr9ipvBoSVCSUSoIkqi/kqx7ED22n72
PaOz9Hk+S1ybQ3SRGMv3cGXvk7EZPTneDga3aNXNYHZiKGtaYw5m+ABuqx4+irBZ
FrsyE4BDf5DQe7ipm8O1NMZKWIXDMSAjkhhjxRICDJdKU4w0JGcbprGIIimde8Ya
nVfablucBgFKla60DIjICS8kBOIMWE0ggnyUOtYsnPy45BMVsIaQWPFDEwmd+LAq
D2RmM3/0Rv00DKs6dqFywsQ5+jLTB55qcTR43nYIBZF4XSmhfgwhCyFS5bRFLcAv
lcnoWwzQwhP9V5Nb5HnWAte1C3wJ0wu2Akrazb8K6U77AL3zg2TLcj6fyGCOzf11
h/ufK+UjXzOz/1yK/OBV9WI0Q5k9lGGAxcyr5vzRSslAh5zL/EJkzS00X4CHgXAh
Sw7tWXWiy7e/yIEE8t9Ehdi8ymCWfCXLQCJEJYOAN/wWMMSmoIVJ/K69lnq71Xoz
5NJJg+oKXxfyWujKCOvk7UXBQjqQ/cIQ91DJO1Urducoj+oD3U/CzgK5YMrHYAAV
p5Tqfa47FxlVJWp2GEnYAM7PmPRnwD4/tPNqo3ucO9hOKjP8R14b8+RfIYzGoYh/
c46+nHpjlZI3R+XulqYra7oZVR/SXauG91sYJHCZcko7AWp/YZTNscpMkLk9Phhr
n1o4eo5cEHXYtmxd2g+tqiEC3QSnvLnkGoGvtwebUxGScPEWhh9q4HX837B6jkyQ
nqY12tZNyyOCzC4pfCqTJYaykCs1VK637kaoI8MY3LOaHdlCTe107utxJwrPf5my
dS2iUfpKfsUkJvExsAwOJxwW8lPZH2lUP+5nU2JMt2JELwVfRLssqRRD2az+Yw5E
VAgFSkCuN2I51bO77Aj7dw+33z+iwgzbI9NpVkSwswPopD+zjI+5eC8wfXhraOE8
o6VboeIc6+s3gnPIWaUcBORa6tfxcabLqTvUf+AaAMuxdLCr2iuCkUFv+6AsV/2K
jJTY5J/80grzPYcLnc3bVaa8Kl4CQcAJkx1PpQkLKdsyemIE73tRPRRdDrYd2QkV
N1mO8wlGoaiwMIzaEAiJGTxT4GtH6bxPyl3S/59uULFj8WNoUEWZ1DF0LYQkcS03
49mqjLXLdBleBJfbuJUomgy704HTt+RUKy2EtbvBKSb2LuVLQr1edGJBtgEJuQHd
VUBr97o64sk1R2hP1f0wscWDkPD54tlnqgalxKMdNLwmheOYayj+UBWAhNJebMUl
d0n4gGnkJuR4TFGzcPvE29F/EL+hISZdEv2QqkwHyvIMovmuLkKhYRGo396jhXiJ
0TQD4ErD6p+HhyT1WEbePaQr70IJkv9Ktm1PIJtRNuKv50opUOGrWIF6j86dFBAR
/PQGy5mlCiTsheZ4eXGuoZXgQ8rNzNikUgNn9ZI2LTXeXMPH2j1O2KZTHiGm7/G8
sh8GegiMCGt4oBXyZEnfBF+edliDnjwl7Y4dIoUOE60lRo2zCqY6gw9/iohUWTDG
95DICVYVvRa85A+1Q14qqEA9WxgH1uscKyhQS8RWosp94cmrRjuSWSXX2ZOMWso+
uW1/t8AO6sF/r378TVtHEq+6+pftu8q2DmMpk2WlMbfR+YqHOBqg5BXOhaHogQBU
2bqwwo42HcExn7miyjwy2QdYM8GIAqtphPA+qCKdNm46UcQ2kqtGcQfHM2i6FoDI
5toJirn48K+Ife5cH2N9e0F+w7Qiaa4U3GkdRC0SS9gR6Nwk8M1W6aS/1FABSz9m
fv6U0HpiZ+XzpVzQTNne771QCVBq4jPOwFTX+EQ9KDFxZE7wpn5rXVOjyvVoqrr2
QWvI7oomw/VkLkQFlIl3ti5P8bREkqwq7oDTnhhaiWzpRBq+6ZllQPGhbPtWX81S
u3aMT9ARwgqL58wDo34yrd+Be+bpXi7VFsXZVal5aUDH9H1yd0CjgQlMpl4xbWUs
lizsr0Q0eNH5NkWmyZfEIFDROCPgRgGpkdSJOdUu8W4X2fKIcimDNBv57VBB9Rra

`pragma protect end_protected
