`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
RmUSF9WApELicABORwSJE54xP4GXI0QbS8qQp9vh4SPu1k3JtwXv+QVRPLs98E7F
UMtx5PWTMvlPPDzAxV40kjNc95g8KiDJMbXQVDp/fRt4TJBh/8dIpWFBG8dPSF1l
gaoDb9OFz75KyalJKw/Yxmjp+VLEyB4NvuuEH/G8FUI=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2992), data_block
cmPT5FzGR1B2gcJu/RR59UH42G3n2AInpV7Q4jja4pDtcTAwlLxkZesZhQrNxAr0
kBQbQk/5KJGEHBKg3a37ozY/dKj8mqLNQEHJ2UTDKevyyUsL5B9LXorbA/DVjInO
QXMalujPKN2RGNjE3/h3WNm2PDbwTZWAVryyv66p5AZ0/QLuu7Z8RtX4vBs17si4
J+YcGU7l4mqfHlh4k9T9SrMfOzZVP3MXWlkolmJuEePhvoRbT9BTj+rcpVLyjWVs
NLIPEDIVhce7tUD2Bzz7NnC4Gn/a0FNCm52h4Tau5Y43aOQFiM6BRVcSflsWPEqe
ksnzpB9Qh/biHbwN+kUIlKNj8UesFyhfOgLEPwKz69Uc84Kk+yof6hNNPIfH2zue
f5+dQilBndRAsrymJt1t9S2Q0xT4ChkymqInu3EELGQizdj0bQzLNgALx/2vODoR
YlqmghRyPj47swBQXkKfW4N4WES+tU2fAxfaduLm+k95BPw13HkfXhz7bJBAP4bS
KF+5i31NtzqG9jJiscwxyDGfL9AYIo6BZcWhHnVHsqqu3Ao7Cza1VqGoU13k63Rs
E9NyG6+qxWl2SAMsv3OMENxel4HIzJikvdFhuoXO7LJVCW8jTXAlagEvrAjtCOLh
5WHSsezOUIwG1CtQdGnpGewg3iUC9M7djEpVy9lcZKVxXOAeSNsrd9RI+JcACEws
F9ykzCtashA33dwShtv3b1Y0OXlnfo1MgqGaXsipAJW5siopkjXADv/YrW1ZzyPV
ol/WufJ3SsHzFAcKVhauW5wXI8dz412RjVl95Esjb85778cwbLdVDuN316Nheov2
7tdUsLEoalBcVtkyxcX5KHbWbmCCDGFZi3ybNXF+gZe76CN/vcY5Zpzh7BuPzdOe
nvEyTTygyccV8Bue/EgoWDvtaUjd7jBiXm5jRiHoBekJIKsRkV3u+N0hEi+COwZ5
lS56XdZhZeHw7z0MnlTNKaakXXAQtZwSbP8bAoD8OdiTSjPuCLAxQJBMvlXcHQm3
1RwmRCn5sr/cVI9QIYiueXg/8G1+qt4L8NiZAGrDga+mpnXaf+d0crpl2I5K5W5o
FqOzlTvlEizwtvOr6PnXi6vE61cn3S2PPkiPyR48HyG29QEZKhXcnLQPu0GeZoLp
TCeNbuPWoR9pv7kZbY4U4qZuy6sTunSKLdVpBMP9x3Isly5lx8lC7SAIeudSBBFg
LsYYTtiSHudr6VYcATAVA4+Yptyad5dTeDYIOvz8ebAYYD4gZ4Nk4iSqctlHzb1r
nS/KNKzNC4tT2Yic4GPd1kD26wt7M4u8foAVP4JCmsl5sDjDEKJOvaccqFbaF6aE
mR++36FSit1slMIn9dnCOat8YQTXqpU2cMY6Q/n4pPbYyhwB6/rml60kMabT/tUx
oEBEfilLiOy+i+e7xhX56OFkTdHg24ywc1x0e9wWRCDVVZf9vrslO3oDrZ7G8Awm
SoBssfNgtybwbNIaUDpMGkVIPf8M3/LtQiHZ+miAn6BGuuS7K++ORkD3EiK8SiYt
3KB6MsTmZAPA3+i9krVEmXzObVlomRRGIZeUMAZb02YZDxaXwLIl2lPzPuAIe8ck
jlRJ2VG9+CqfXTmSeNSRBRHgHGUPYnmkiQaz3/kwZT/vVqKJJyJxDx4kv5Vgsc16
gOOoYjX+CIYVGBwuyRMXr20oOgOoXMC/buFX15gBfWZ0A7tV+VFBvKVaJk2crYjS
BqoO74nX3GhQc7PxhkihuixSaroosHOuc1Xue1oq0wginPzXZyTQxXTgTW+WZwcD
89J3/ui+eJlnTsKThwxgqDTaUCpPSc1E2K+Stq6VdWISH0powtbTaqZVVjQz0oJ4
iOlw0D07sDIGImzBeP0jw+9ieHLwJwHJaS8A70xvHhfHy+Rbu+PVeuyW3rKCK4QX
rSnlMKJ5snHOkibB+ha6nC7jPSwi7NEI8v2xd4tfUR9oHD1pMUxmXqYejv9JPfd9
BE2/71TmYUkrMrV83C9B1QkIATRFbCls0EJ0jze8MVvXAjGhcPw5hHWeI/ADOFdE
O4+jknJHQTjRK4/HlYo8LBW+fHwZHrT+Muk7hFdYRZ8Ne9P3fC5GxVggZv870HvP
C1nCs/ppQcEkzs0RWhECYu/f1FTpGXr9QEOQOwO0vL3MPGcD2i5s37lY8k5Dgv5G
bXMn7H6HV9NEVR8CRY0b+VCdjTvHe5S5/G4udTLtVEaFyTdz3yFKsl3NUClpBOvu
g7PriOIdd21pzDip9aypIgTYsN1E7l7onVaLAHZNS6TW/Lft+3HXlXt+o26RQrvi
ic4ZdZKfhql1BIKLPZqykIsang5tM2tWpmY+tjkK7sKgCzl/Jv7Z+piygVicx66g
g0eX1Wc4LUhLNl5AxE/nZzWIUXRX1bhZFG8n67jTz9Y7Y3NI3lgK0RO0g02S4BYw
VL2WOzCIjJaoNTRNHu5hdqgfgKyJ2jqp2IHEZOINO33vQGp1sdIdHaKchXx5YdFO
arLYpj1NOH5MAfqemSLss2meTgrLx1d6QuTM/w34K5bwFPj6oC/7ypkKBokGEyEr
/xjgPWgS9Pxnnehg9nPwzcVbucIedCfGf7Zw2eAZKM8gdumXfKqKOIjPSO28XUup
sTOpg1vdJNvzFgTGF+rEzTv7ObFQgxFQMcEOVuiZPe2EKNoFA8PvTNOJrcQIOTxq
40EJ1wc4matI2IrIP2ox09HuWLqhLP7br+f/JKgp+7J4fyLt10b7chHxy5QLAkC5
FacDY/kGYR1lvE5TQFU/BvYRst66ZybqTGrnd7h76KDP1CfOPf49CZ8AfdCx1EgI
G0uF7NB2yLaXmHKpf+BcEO4INv/WdKY8ov0uUbOV9l1NsjqFIg7GcGBFMCYmDkCC
zctTY8gx4BVSXVzBuJiK+hW2PEvVbMMoLIwHll1InA62AI+15Ez9yszEyZOWr+Oh
4QZyZgwibEj9puM5jMPjDmGhpgpAzXjUNgk+NnUxhKahos35Ut7HO5jCO2zkraiN
50VLAUNucTNtRbYuAirnD8649NJ9yhAu2GWkkAoxvueCTns/D3bZ/B1Np0P8vnMM
LUk/UwLEYAUU4plvs62l+W2zG3ce3J4r1vVALqvfNPXMbRkoDjG1asoUw6LvdLCB
3t9hVDCIsNq1KdQCS2GXQR5cN3MfP9nSehjZ6vDj3016uRmbKZOH4XtM42Qp2qEY
efzPwkFdWY/21hUAyMMYGXnGsq+Ix3zth4L32Jvbzo0suPzO2kOi5qssTG2U08oD
pcLUhhQJM1JyePv2/MzY25U73WC1DZ31U09K8qYoCvbQi0J5DbHwh+Ew3LA9DuZf
rbt8K9gdBmeq7cl4RG3IyGyOwcREZsObEwgbnEcMTd+kjjpSFoPYngsuEWO8ypkQ
wJVh4I2WnIEh3ZozQzX9M3g5xix2GPdWlpt3+25nAWRQJ0/kjCvPCwyOKjEGfAcE
ddbgddlKrdUNe38CyQ9pvLJOqiu3904QvGncdLchLfMBStwAD4S8h8EMEO2RRmWa
ruufBziU4+kWEitVBpBL0iIuHPqPWRbWnKXGIaJARzNqqHsMrZ48LEUM0IZMzEWB
+Qchg2PH4fjd5uws5/lVqkkqutH6iR3sGpKJflZK7IwtGkVVflZZGeliNUoeCT3f
pNKsqgVsJlFeH1wZau9UgqEVTBONm3UGuS2CjjktDgzFqEwJpD9QNh/JejJpux74
ccdast9V8MRUqLQf4ysCFbv8493BxAICr9PweCMtJO+BLCySxvMj8ePk8KO+bf/c
SIGmqJwhCua8mxUVhfUwSofpJc9AdgEXCIpr3VvPp7L/jbnG74FBkV0IPB+9ae+a
Z7Oma5CP8uMD75pCf3q7LjCb66EC/36utzWQp2Osrj/zYv4POFFRfJbNTiKQuzdI
pDTldMkNpa4b+6cBVZSPpFLE2Lv8SB51MaBY8lCMNcLDy8wCojPlgUXn2ljF2Xzq
0AHX0YYTZDTG8Btm9qXoVg==
`pragma protect end_protected
