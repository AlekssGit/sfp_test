`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
njR2mD4+DfjyI/e2PeDV+ciHvMvi3XPTQlNkRuL7mKdCc6mfn6ZfcXijpLnO/M5H
wU1IOG437jlhGK9MilciCJmVnE/U98fdEBGKajVS+IL7QJbTvFSjRotZiCccDFix
0PDh2Eej9lYHBQ0l/9aGWwXtBYAx70SBvUVmUWbhcZ8=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10752), data_block
Kg0p5LoRITB5eSd320sRTkh21DBxp/A5rMkrh5n/fi05LWjEPUo7D9QFbFTBMDjZ
SKItSGpgb6UTGKyNiheTXUJAVQPzwS9m23LdQzQeNQxPMmc6m5AwN8ZSRzz6MatO
qa5dcn+4xjgfd8Nm+QkX+YX9w3vrJdb2UYmGKiyg1qPxV5FFRkha9G11ETweryJX
bew+E14RffN1mIGgKDpQR5JbLAZZLTgLOQjKn9yVXnkWw3xxddOpZvCXc1WSSKhl
CrEF75nBSwL7mfg4TnY4zNPFzWEtacYBq3brbfL0TEYsZ9oe6rxF53dDo3jiP4eP
5jTTVyUaxeWGqjJsNXbPE4izVaOTnZxRDZ9HuSoENDJ5NB53igiwSYH6QR1KTBYP
KTr6mXEdDasU1ZVcwR8LLydAV2ltxqCynvADBbfqfsDL8D3cJkyUms7d5divEY8z
CvFKpgvssS17dNyMWGZkxSIbiriGma7wyqpTBxMGJ6FRrw+gA73jhC6XqFbsA2zA
nw7vfZtsj4uHxfniL2UI9naoLTm32WrNBpRAk+zU4b3p7OG8bjQB24aN0ixHScVO
XIsej54XNQHRHkcZ68yP/lrYLlqaahXRH6hayidaAEf7BuU0ogdCT+pxYYkV994e
5nPfTnPUEp4cUGLNMeGJA7C5gCJgHBm2CazNSa5pq7oWbFZA5G3M0H0V6jh/ryAi
XgVsRnvmA6vGtqBv4LPXFRKbvur0uyqIW11Fm87Y3gvvakkgqWYKw8Bz7IR7HZpo
SrkzUK1Syg3RVCxAlsebB0g40uY2aUNo14peOXyRO8gh3qqa9dwthH0criTfRnd4
HvB9fPMBFNCyD4Luy0LFv6Fn61wcMptig2AhLcMGdCoc0qpumrBMpnSAw/apVaMz
Z11LjdcURihPJLhOPo1pfyrX1jw00n1MjgBGImlpkM7lbQwQWJZDosegaOFYNmgP
1PGz+xbBqsk0BhfIUwNHOp0NHFhaCkP2f5rDGNOceuBoDq4djLWu5cB00yvLKsCz
c8cSZjoOm8RFLhd2eoxHEIIBIt3KuwX/2Rs179HYU8bGG29HuIxr6wSTDoWfn5OX
AsNEA1m0DapyEc4OuVDbp3b4+Rga+f9tTCoLqNPrPp8pXHKr6zQjmXLLVc0pMCj4
vI33mmGf/r+kc0OzXx40EN2AwuBbq2skCPkdOyudu9E1zPI+SsTEPooXzfXIXREw
PkPHRzfPMeT0v0o+EZdi8NmAIHm0O6eSsLUZB223qqLq9PsmBA075UYMkGVrZKMo
SC3TgJBT6zokE2jxSpCFge0gzVDQCVjKDUbL4+HYzAYlLmNhfIK8m2eOe/T+7HCm
q5pTE8IJSWKc7hR0O3GhusFHthlnMho9Een0eLpcTdTZlIU3XkJ7pdmT7ijQbk9x
u68xOOm5kFCPUH2dLhil9X1Rjf6UBpihzdGxwv9JmYBDLpE8KXctk3aVSfpDgVwt
lWKmEew+mw/KbPV4/56aj7tJOdWQJBm0a/NSC5GNsc6XiZYIW0PxN1K7QNOmWK+x
dafEmSPEYscLpUO+D9AS4M26housV2pGUfyHZz4IYi25n/PBX4Q13FG6oPsCgV57
qRQja4vc9dj700Ore/P5/TYAVFFH8We3qri38IQsQ3yIX+uu4+Ks8H3U/zRear6h
bucB9jAH044yjXM2QAA2vIMUbhoO7ZZ7sUO5FFxPXlyQwra5O+MjfnxhJiT3Lisn
uMXKLFjSmsYpyscLT60iDh+mRawL7J8gsBNY8JhamhYC0bKJrxQX59ceYgJ9yZIC
9PSRWud1FomNY83nn/yKYNgcNyJjXCSEHZTBgi2BzpGkxkS+n6YiMKj/f6MWxpQ2
BViqpf3GyZp57F44kX2YjySxGg3tfCLBPEVYdJTgR3OQTFc4XnUxOTnqYzIu2hul
FK0QocQ056wyUlsbu0V8VzCPLgfpRr4dcwu8AbC+PSokJs2C8Sueb4N7/12Wy5GK
n18cP05zpV35+LVCBO/NdXyzmbnTWXThAGWbxsTvLj0TBnpUZDUlkepXfyjjCp7O
jvSH25F4Quw6idJoWz7l3oLGblmU0E934Mvkq6V6EPUXlQyulln/6uPHaYrcLjWz
ZrC82Htw1DnfUWededYRS3OgJMKMylwA+khzcdlMns4u5ItLyJA0FQi2SVlaNM1b
TMjKSIKeW8YI/J6JttX8RdASMKgI3pHt6cZ1n69sNyo/6XCw/QR8869EL0BQfCmb
bH/7YXVQyqfnQQyJj9COBNlWZX2u0nRb0wzKps+Wp+1+J6Bf+hU1gARy0lHL5dnY
x3woCgpovg5WP33gTNIwvPj66IyE/4W6tL0aexMjzk24xuPmv35qO+WQNrOKhYjj
ITVXBHeHlAWtU1yZxNcsUE3gCFHko9jIEj9veOoLcRPFx7i680GD0VSts2iy3ugL
a/VJg3IpBctgMx9fR2kOL//Y/d9Qv1b8dswPDs8wyb9xX5s+YpJlg9SuPnB56ekc
3VYGWxyG3XeIrRzAU7ihYJ2ZLXNpmT/0BKod2V0dJkEY7n3im5yXkpumI4IPtUja
3DnQia4G8MZe7hSCV7i8iJp58o7ZKh9GWkegVMnj30Zm7NkIXihMP0B4PJ85QX6D
ww7yz7UNBqNXcgbHbiwRLqr9dSGckcE8EADOIFy7w+seU3obBZZEDU+rfLlYZila
+B6Md/ozvAZGTNOsTkXsMNYZxX8F+oYskuy6qBxZWAx2MAmTd1y7eM38ByCRjABe
SfvzVjA8voSCH5UXGQ6zjCON3OaXaTFPP9874riF5qyRcamtlorLvD3zLS/EPvVz
fF4yVBshqKXBdJEzUBk/Ml9Ajel3Y32qUQ7n/H4crKoZvhT3jlR9Y4DF6cM7RjTm
iE76eSmeaUNas/KbjpV6DIJKLPOmFtHUMDD1NN6LfSLzDP+IIbulmrNC2klCrLlE
3uAOqTjRTaH/2As3Zsb+/XJH4rjb1sKYzjVThbVlCm+Aot5ySnoyMMFjepGdlmOx
8Ol4Ti/nI+OoPnB/mpx3rc3sami5Jvx1yi8TgJ2lOyJIqLXhmm9jo08whimG26ng
5z7coa7hsnOxW2bF7wmJZbOSP7HPOAe5p/PcKadFzpXDnQ9arBz8pJ8p/XSU4X9H
uY+FfkreSIol3yW3fDNSrctyIXBMmMfQX2Lfd+llJfj0hbYTd/oe6R9g9/9dDAa1
91RHviAdEsZ3dhwt75737IkeHvljncn9KfJ2XqvhcDlyfR9Rby4DQtMMk7dcZYyV
auWm3BOba+HiWoHLOB2c1Ll8Unl8XpkGtV4jvm0uwZQNPQy4qrSRBVKnpCAyCzaN
QB+r7X271IcUzzp5EJgA5Lvt0gh/T+5a8E3DpWKaweFqG7BYwFBQN2lEJ9yK00l4
ZwdSBRsnv/GYH28Tn5yqa3L2OMFoKgNIb4Z3ZPxyrvR2fQDkOPnuzLgKzvWXz5tQ
8WVKPoIZ0dKlREVgGAX2BIygOfgCCvUKL42TXhxv7Q6S8vj4wrQvp8N3FXhq5F8L
ZnFmepHtnpmwPWsOGHlKuOWbCACprB+60VIwdTIxRnB2m2XSDd4W7+HHCGR/UaP3
FDinyGk+YeIp9DZ9yh1kbJcNBr+TTVC4DfvGizEoclzkOazfWOBNeLUEZE92mHWx
mksbz9quIL6MCyw+zSJhuTg7+YEGh7ol/ez7yN9cInnrxAFYvzq/uUWRAOM+mFIm
OrqT5v9dwlaBbv+Tn9rytcClk4KlJCtaeACKlNenJJZH1QHht53N9QzA3l3kzL8a
Lrg4sw6Vu81cVtYiKMBe72HPk1ubT+Hkhl3S11W0adVfB61eFmJAs5Fv4u4aBeP3
nE6i0X0URru2tCd4Adf30TS3BxRi+YQJkCoSM6L+sX40W/1EbTL4w+UMlIpYnb8u
XKopZlgMFpqUyjsUJtT072IUdf4KlrjbjzlknSD4xQM2LhnmUyqwxgLigh+UroF3
Lyl+ylRLUX5VN90kgiWc8JaM72fD/bnKlCikxNij7S0SKvuFhthBoo5jKBQ/JlPm
nFSi9IYY2Dyj3SikQvH5pSy5w1RMDA8D4z8qAWX7jT88cIVluMJeyCn+7KQGykge
BlJpkOsiEt3iCiOj8j0T+yB0xrR2tqHgQvFfQOT4BxemYJLiIV3H9ebP7wO2nVUc
whm8V4buuCc+u9p3QsmFJO+S9igLmRqnouWezkPU6ApWZ4JPsgv4wijxBAFE/H+V
xcSAtIJ9snBvW0NqyvFOSvygySDPQoebdQy3qLPsNS7lNn+pjuRqos+CzurR6kIq
G/lCOmCJyNBng6nRiIjbKWzi1tT3ZA6OZo5/gdl5GEN6xpy9Y2bnIc4R0VpqpWLV
ww0X6cQNQmohcrQixZCTemkfut8L/IY1jxnR3BYokslC+0t5ATvLSkFityxeT8KY
3T7L+2rrp8TOLpzso+Jrn3lvgoTpZSTbiSAzxZIwFa3n8Mzsk5uvH8ko5cXnjT9h
zSxwAQ0vGdRYcl73CLXFpU9XDbZpfhK3O4MQQZfIZO2q042BUw+FV8B1fLRkCfPL
vpSi8IaGBS5SAPwY03xJ2U9obo75SaPsNkhDUz0PfPNlhCXCbzfFOnNzhUuMX2Do
Bn2vTVStLZtEtl2+I+fKZyuh4cjTGMDxvVepgap/g3ePBh0/QSiwz9kHdzDfdpld
QkK9RoDpq5O5ra4HQ9n/XY2L2AfbQNMD1zhecHI5gNwfNbk9Mq4A9ftZqB9bF/Ew
V51CWokd7zeb2hUv/YTsD7knJtpmvdcgUIxUb4AeU6kt8pvhPN8ftvGK44d8Cwsb
N4IO1tUKCE3v412sOMRYeFZw83CZI9NdBolWxyJ4d9i8Uet/xikIJOP5vZTZDfqm
zFi5F3Mq2B31E4XWU8a3ytqTx8Vpr+8LGgYT9/J9+m5fMpQaqULgIlWt87Fh4KgX
EtHjw9AI3nPjX/2UrqydYHjiQP1RO1RUr7oZ2TDiIJmuJnDR/QC7ml+mcMQNJ5Tm
RggwyQ9uZUe4mtl0CGZrYz2Qun+jYqja02ojgdiBr55pw2oUXGJC6EvGF7SuecGL
wuZmYDY1DrkOqUIZq9hwd2+cvux9utcHhBk3vVsVAxOoFllOL9WH5ckmS9HVEy/A
/viBdfE70ZItyYhhBny6RmffIBxc2TcaEE9MfHnGf70nQNciod6hrxYR7DBYdzM/
4NtVw1ffqVuprZxNl1q/i/uccS9HS1cfpodftulJG5XyKTdsnb/SaHuk9//9gTC4
ccSybQRpoTxQVrNhXzyWHv9+ka58T95A702ZQrpCjv0Z7dQY+HkFmAHHJ32FOnqS
KPokGjd9TuqEhQvZgIzlFOo3TGsI+TGbIb/2ssWxtIUblvZMlCv8NTAtNGNj+DaW
NsktboMa6x0ugHXqemqX2J8KTdbH87fM7OsjRYe3M25arAoc9v2X6f6o6OoDO6IM
VzknNtg0xxDAKImvmj+tyXWDaBLdyIzKhCFrwg0gfd2605OUYMqPb7n2oKhZ9cPM
EH/v0OmTBo93PFtnNKX7EC3BE8cvsTbb82SjXMKRR4IjxukfSioAt9m4lcNF+EB2
pVSdlsTxAorV0kcaRmnldomWfi6Eu3rVK1AJqjIlzGu4EONoONo/QEpmnFwq1NgO
TdKX8r+T/Yhtc47p4ej7ASndCOfvjQtyUcZwhxIGIfbM4i4BL3b/fm+p29zuwkmw
EA2T84Y3PP9ZZtLOeC7quVfXYOAiH/nDOWO5nRN1PrfDJVfXShg97MFfFbJ19mji
pJ8Z+RqmQG0tu0x21yh4AeMgcGiuxfHsxYEgb3FsalfTmO0h53ypy5I4pzDwqcAb
vg37vTID6Axe0E1NhWAzjv4hdyKtEox1jis2YcTPO4e/qvey9qLN0BC1q8bhp5Xy
fDf4KPWl7i6QqxJ1/gaQ6LVm7zfMrgE7jqwBBJ8PjfENdT0EM70tR/N+BAN0t478
7zDpCPNTc0rV0/OzHjoU5HmDDWf9ftjQ5hj1g0t1RSrGyHPYhSz4kOXAzAVA2272
+AdDd0TyPpuJ1PujtdzQIYIh1ui/q5pz3NW8xwhjtalDVQ68EtjP4n2jXADh1Jud
bxMGWp0a/s3CWO431Eqy949PhO4/l55wDo/iWT1fL2qLQPp8KebGLkOTheWzdIy+
ZXrZnpSAqmZjnYe4WDoLsqFIMszj6kMSvNARDAVF4xwgwq1WGNhseibyLl+JzaG6
V5qzmhsawYjdVYdxd+tiP7c93DimzQclzn5+9ow6jIC38MNclqagKALpbUibxzUG
TujVlDudXuE+B4Lm0oYhwPxqEXta+X4u0pIivi0HSLqyC47xQX22SUcwDHhLNjLu
8iTxu8mf3aTTtBPCW1mXeld4tSYBlMBSUYSLZJYpni52e3xggdNa4fWhHZsHbFzy
maW09QLekRWDkYFKViHFRANxpnLgua7OenjGW9pffkovnjAIY4SnMARyNV6HjUbt
uHQKqZX3Uf6ZZ7NJvKjf9CBgfhRl0MUZS6cEHdd5XWtfxbTzwk5BjI1/VB/T1B+A
rI+NJtTx8utDcfrODcjRa0CwNMfeUNZpupS/TlSX3H9bRKZ8ZQfsR3HfuqH9qyUD
HrrTwpkyuWin6jZKo1Q9NIGCM3FcF8fJOWP0tGZAEkdBX9/IJgfYsACGdevkEk+a
Ys2PtqgIuBa1X8wdqCTbmwj0SC96hSvGRvOYsRdzLXx2NkeF9+IQFYrW4rj1ZjD7
WT662nKi5YDdCFXUO+STKRXvqjmnLhESycSbTU/6FU42l6Z8GJYVlMISTKkSstAI
n4/U4cYfwBu6JwcgXgKyA69MNthG8ZCYETXYmsTJi+3SAQV4KD9Fm82DdqdEj+gX
11OW1Jq2ZJZPdGRE5xHFlX6Xce8az8X+zkTbRpKBAxIs2WS9hCW5Ep/XdR40SgHx
9J5EeF3a5eNC+Hru90aGJoA5FBmpwL2YherBQ3drrhmG9jvNcjxeLzrP01QdldMT
dvQugfBsV48a1hXWWiuJ+9A8QFFCzTrHuA6Ypls9qnJIyrcG6ZoTLad2kkUAew0d
RG78fjWWaVUwDuWJfomlQ3vTmBF8TV8C65/XEW4KKLt8YOjOZdEQSRD67X42rNmy
d3bOtF6eTvxhtTfIzkFa97CK2MaWQvQxN2gHuniv5JKP3C3eUo7MN6wIT8I1oGec
/a7Ktc/08WauP6JX6XmT28tY7Jkinf4Y4mpg+eFinDmG3IGaMAmSdu64047Nen7E
XEHM0wotIvqKQkIGx8Ij5ejDptuCvVIXHLg8Zh88QWSrLECkYUnvn0+dCfOaVYLM
jKDnnEXobK8dc6n/G3L2wqM305y6DOG4ImiH78q03ZP+8bnwUAN4aYNb+YLPHKKC
a5jzBu2mxJp4Y/dFhkfVnvUk7IlB4ibxW+fA/9j+Mtfhfhqft+gcsyWS1J7me7ep
NU713KvgIWpj+3FJdgYH5FOMN7kF4k/j90FlBLy3OucIW2HuovVwmKS8T1V8l3BQ
JrqnDnrv9E9MZWkeljSRKq49zBRqr3oSb+XBb5vOmnzHN+/+MrtLWbIs5CQR7mLI
48q0ZWTlnjrWWrACajsLgpVeMDiyQPa5fqR4cPLrs8QdKrXNbB0FHUfi37GhZqwZ
TftNrIrxPdYGJVBsYnVkUAQZCkCcYcvnpNz/OVT8ED9PJdGrISwZsHHt2paXLHUk
fZhM4F10sy+AmPQIfBVveClP0ABBzBPlU9yeDG63nb4k4zS+rMUQ1gmuy5YYZAe9
WNCSRo32K5yYiRl3JfGVdaUap2lJt72m2GRLyFctORVg00B/jsSOn3lcs7iTiNxn
uYB94qvDcO7W7+ick2exgeTncko8ZLLVIW91MhKXqEJlwtP1+5wnpFVYiOamA6Ln
yC7qXosvOVn+KIQd3QLgY6/LWUxMZNtPyQhkNz261srYCzX3Orr8KNORvKJwKg4i
/CF6e7aAr9BjKk5C6bifj1Gy7DAOhrGd005DDpUB9kjQnE15thAxeWbAt3LeBYPu
zYf97dkslzkMGBqXDde61U3RQ/5Sx3X5v26Kbb+y1k4RqDfxO/pLmc7IT7JQf5da
Fb47ygLluj7nPMiQHuNZsNvrWGXRhIzsicz7dI6eoQSrRJ41F6XDaTrSzg1EhtGA
zyAB95vCVjSwNs9SDJKOwPKbHfihohrjWk3EnNYE/duk6haoS1LLO+r1Ra7PuoQ1
2SNsDasbWR1jxPc5JFrW6mRpMRRjHMEI4Xr4vVVL/YvNCpy5lsEyWBIBG8IjNMfV
98gbRTxvBpoT5AlhO9lus/mZxyjgg2X9mqsKQZDTx9oL6RiMKtKbA4bCAeh3GgxO
HO1rnT7xHBavwYEEnO2MtWgfESxgsq4BYaQ4WFSt348qzAPGjhEuE7J9XYss8j9l
V2JrynkZePY1aEQvxkKwojQUfWs4buFXM1s284nP/Qq3hl8+QUqZtylx0ThJTJYV
EN+YspDZTjVVf3OlDD/n7ZHOesKp13wBt4aoOJrOkj/FPGfdoW0UaveaF3fmNdva
kU9u7xq0DI0jXLn3beqQ1ae+hMVM9s1SaRWEhh3XVz6jHzAaCKnwhbvA+G34N2iK
O4MbbeJ6kYaXolDjGmNZlTPNZWkUA8ePb0kgaG4jLsLZ4KkJ+6inkNJDAxOKbcRH
DVx9TfoJwd4/yri4nqRDgz1zDl/vZEfl7KDZ3ZIzD6TRbVzJ4+NIQXuuTFXV6X+g
F44o92kXAgdkhTpVkyUOLHZ7xOYCwcC4Czh4ARnHGC3LJBlr976GZKx7IQU/M7d7
71mcbkkfZnImkUpOjjBSXyDfyikgXGsk9ZPLo6hwoZPsObMQFTWPDNqVLItr1qRC
kwltISfZCSyJ81i/M7mHx+6LpWrqQH0rjOqNOz29A3VqdRixQ1U/CtQFpimk0H7N
hmuN0HtAl9ocQKIXeBT3pAjQYJr+/e0rlA6tuiqaIzZBl1olcV58YTNG4PXxyKao
LVV93huYkwOVwBuSCM4+DvB7s6yRqv3tyk8o2/DLJmGN8jAM/YlYfztR2VyPkmvP
+cLYLL8T7UnU4eWv5P9qkX90PkKkc5pBPR9Zy6SjDdIOvmg5eGea/vx4DoLmUurj
8Lwocr/uB+H7bcHavb/7BlL8X+PXN1ruuCYYtI2iNj4qMEsbFV+ezeMNzAKf/N/T
cQdGgsz/scqI+eglahe1oTpcrv1EddiKotJ8VeKjG05VN2oEuczbQvCin+vzr5uf
3m/VsjHy8E9Ydu6FPc3OfoOM6yxsgie7nlMEVj3hrl8v0pL09ttc3cVN3NWPeNIE
/bqZtQfLxYlBqdgXzglEpT49EL05IW8MKSheZK+byrsHu4jGyCZdEivryJe6H7RJ
Uc59HjCfv2OggCQZEagOe/qYQ816P2USdhAAX176y/cRcJJq6gFbFoAyhGHtlv3v
dEJMl0YZ1ybblvCNk6UoOsR2IpFRqqA2GpFoNmY1u3Q6qI4zPot81hWWi5IFJjHK
Nn7oTQuw8NwUKX2nAFUmZOq/c6LKz7MRi6BoHndSkkgZ4ma79TyFXi4qHwaO5YKd
I5UsytOfaKYA39eRAuScLi+BTnuFqtDhIMV1VCKiSsWPiAulnwWVtAGnff2GBddb
MRcuMa61lsS85LqehimyQ3/5m/2dffx5xyBE96kd+f0nXpu1eS+2UPNzoveUWDc5
6tb0QZHdbj1bR99kLzvQf8tTuBQbLy6NPzQQ2LBia7qznub4/WqkF/yQ0wDciSIQ
sWnmf2kQsgAsL1GG3lFc7ZuQCvgL4wKunpHw6UIsFxsXahqOjCfbEJgwYNcJowYO
4W3aN90J8ZKiYRR8Qq7TH0Uv+B/MRtSGeOjOeVqaLrPqqpzBk4eJla2Y/XJ9cm9N
XbLSHACfnv36HSGtk5fY+MnZcBbhKCGJBP6kM+oaq1pot9emVcnv1jMdRwFE7yDu
38IrK+3weXNpVKLP3mjk6QO31jSLgrOA69kPqPiH8TSZOhXEV/FPMuGnh4F1bZE8
LTuN1dbYX6zf8c1FDPiIBMYIzc9HBeKc6ZwKjwkfiSsOMLswQ74GjZWF0nPWirQE
T0sLXCxk6e3Sng+1FeO3iulLLu1mXv3cmtYw0RmDmorGtDubdHiuXdYsSVx3qhyg
JpDrS0U+8TsqcMs9AZyK7deNGIS0LAvgxpHLyEynak2Qq0vF4dDsU1JjBn0DFhy7
3eHxsG+iwrwYSqpCiG9wAbKRXnNvtPa5iSuvnJRyYTkMAcqeO32xlUQ6J00+4kTW
+ru0YK5SSgazDp1bSwTZuwhvVIIt0ThqY/CZEsUTr7sihMCygOxCAasc3ydGEKqL
hPJdx/QK9FslPnR+EsvjNhKq/obM37EvktHZpknqt8ZgLlPH3/IuMLvw0wSlGhol
iL/WqTDMaEW1TtgWp5v4LxBuQ20KvQnS1tmXewv4L0+c98jQB24JoUbZg+5fa4TV
MBjqS4Z7td/+K0vVoQAsBYfvppVDsyzbjtll7g4THku5WbAXwBUjcxImsdMjNxbc
H30Nm73G3F4TLPj+UJPB25Urkoaj7cE4+KXW5C6HAjiHEZRIYzPzEaJ0RiGE4aVV
N0cK0N7Kvd/TzjF0YDaxcTRE6sd6YxI02KIhoE5IxoGqnpT1ATlMQQ9DQFbEsKIo
f9eW46grEfiSsE2owgNJnMwlW59+SdK/WWpG7FRYBqiDYeaemTQ59AjJDWYTTdp/
yUxFVhE3ph24uwr48gWOWi23/rBIoHqs2194XX4XaGD2KZhWKiTrybMNFp+pEX/N
5moYlGiulai98AK3WK2RvkisRMZ2CQRR9jJNtxVMx9qaRxS0MR+VVcZ2T9oBu/kd
LpZkUJqd4TseqI+1QNCGnwuancpIiJIK4u6SFcD5tCsRgMRagf+h7+aOzAm8jPVF
cS/NXfyq8mn9dP7a8QrW3T/KEQFQOF0J7CZ7OuSbDHET0kkOAtEsTefaB6jdaZj9
8btodEEmmJS3UxUl8QBwprrxkEQG3qqmB0CpwLxFPGGQM2zMh4v0lGxfUcu5tKl3
gUi2/msMod0K8mJ06FyNklNS4Mh6K4IaEcGdqT7UgAjgl+McIccqY/+tIjLAq/Ie
/geUWFsEubERsX8/y9R7F1WvoLy/b8Voj9AJDIckrCehinP6BHRvAY5nKjoYbfcI
t9OPYqp091VJl/WsvP6Vqk/FHk6fprzvo9NGwwD7RXpeTnYI+NDPCop8Dlzs702F
s+6zXj4rLBAEYsyyqMEFDaKyrDSynJ3lwRug+tcdm12A5zfsP74jELuDuX29sD3S
+dx7uBdggnOdYZL+a6LkHDFD1+pvGcVhlP11roqxiU2QOGRESMqGNMBOyudPl4KU
hFAw5fq67sXeaUBNFbgf73HmxwoIAW2lQMa79khaqCWONQK1bJ17Yy3109DsLuN0
PEaRmkyQqhQf4vgH+nnUhBlUpyzsuNmgwfXEniIqvL1Z9aYQoR6Rm1lTrup+2Gdp
L+J/Xj04Ecmu0pX8EEMk/BnmWA11NJipwwDNuqplpRhF6LvoeE1y2o00txo8W9Y9
iSLEnAJJsdY7sJ2ZbRqONhCzIQ8mAmDs4TjNwRRwsDrE3NERsPbfY3BXyhf80I97
Upbg+hVaStUOAH7sfgbnZoWdxCa5uguJyr/VPOgcGkiqx4vfmyOSfTST36dIQGi3
jLZSDxSw4LzPfLGt255Ycd9QQbENJUEtMm+BvN3CqG6q0NdCyYC/23fqDlPSt2ya
VeyGgBv5+f6kWvdUW1BXio1FMIYT1YI3URkoVYbfvbNTjLP6YJsHiQwjEqKsp2b4
VMim75mR+qnyMKEkmoNTgJapunExI7MHGC9XnJR9hCCMv6yXL/DdUaT/Ly6dUwaL
Mj97Gb7S/ubud6EZWoQYfPVfKmqO4RVEP4MtR4rApTVOWtatPXv7Uoi0+I9Scp6Q
tDH/3Krcjgp96PPz+iepmMYzX9vPIuNbvc01cUU7NFW2cho+EGce/9LQbvD63436
18JzGnaBWvkH9kFCDt2XkYQY2oY593BJ/RlfgEuB5vAtylulfY2YbLCTYVz1h5O9
Sh9+IRJ+7dMoG00cw+0LL1R10MmfNtNtWU8p08xxsMkHXggc32BmQPK54lr8/guj
U9LZGZotb//2zbjreA3ESNTdXzqXDFzZ+VhuPeaZGzvDDXvQdaeX1bW2uwGaPjgS
IPlkhLRbI05nx9SIa12tj7pEbA6ocCs2B45zu9Ol2HMAgHoNa9CfoNZzeVAcjqBo
8LyiItMlMsmoZ0b0g3MX/22vvp1il2q+bjK934PHH1LlRESxLQJ9jEkuGjhmFeQw
Z7kSR/dtKwks8qUb55PQAA++Gxym0l4B1sbpM8fls5pOdNfznPRCgJks288JoaSA
sNfvhc+2OC4OiDFy/v3Dr2wQLSRJumE29aB9Y9TtKqD/sMMbg6RmaVCRBwK2F5Jr
Bb0f+u7lX+iDUGYeNMymg7le+fasEs1tXzLKImbHQ+Z50FvFg18EuJjSspQwuIbQ
R2jB3dvYE7uyG/1y8KcijSueHt3+5F3zRPctWlTBX7wuQvV1EuFuTJYUTNhyp/Hs
XLePZ34AcUK1bnSvMKYJzoWhujSyTY+B19z/KJDcWrSsayAR/sCoT65LV9PNLSUQ
Zs2UEbtXqPpXxoxNUGzD+4G/A21Sp4Xkc7CE0cldkyQu7acq0XZq7ccpRMyGpwyE
muXXhAGiGUbsTgyVzt6ex5nWrpsThT+qTdu5U86TuJIcUnnlsCrhfyucAICljRZ7
A0HeV/umKIOpZ/9qwYrabSKga7swkD1PhxcBcXbv93Hmlk/erSNzxrHyeCKIbY+R
VSXJD+d6cg2yyUILMNNKFMHWOohQEGTkEGcfPoiE/oyVMWT3099/l6Up0rgBEXk0
yuD+mOlLd97DRjx5RaixbV+QxIEuoqLA+15OImmf1gse4/i05I3YbyWYDK34arrl
tfSmJfaIBjayupf5O2VZNNEdqBtgg1qWvQInv1Xlb2NOXHczVYWQ0oneE0fOCnXn
0dbFVaF561QKR6vY/vAxVdFUyMNSBSZw8b63gAsdP1E0bE7joW/uaGNUSdZRLrkO
BQS7aPkaPfC1UOpFzoIpcrL/KqDwliLV9FhaO3PolDqJSX5nGfVT09tM5q7mf8IM
O1zB+1lI/h2u1hfokDLyPpta3Tw0lgKY6PSyla8ztdXouWcc2nHmQzhtiXHhkfu5
4MctUE6rZUC/HdJaokSNZUDKS/s55g8xI7LgoWAcXW2KoJ2sS5TNwbdIewi+6AA+
tsUBmYrAj+ON5dWfdEJaaOYUuvxp9/l8OyySN6ep/2Uk5GJFyP+/lIT5GWzQInxq
Ue9qRW0ogSTriWo/VmDTgTc6hlZTf5ZB5Ehc1bUU31vqZRI9omzZz2CJOQf/G0df
EeD1dHHymfVghogx0PtGWPf8HCJgSbzGNOw78KMyq2U72nGr1KnLlEIle0fObk8m
osvUNaGm29xOkM8MTJr9xx0Vy7ukt87RKAHldXmtYrlN2mo69xSvkXWChPatYTpc
Vn6I0QIq8YcjaDYTtw6VFI27Mj3FnZk+A0XBUPs51YXH3SoowIvMq4KpAjla/DZ1
pDElt6GEYkez/WnEvSuL+xP7HjnziitUuB4onG3M83BOUDXihfMK1AHIj2kELwi/
Mw6/mkA6MNYg8wra/drICkw801qixYmtfS9VDiiuLxInRRjpS71YW8PVI75JbA/8
04feFcZhM6t8kdvx+keDSIzneQoN8XofWFd7Ll0UNjGIuNyvQW3oe1d4Xq/svHso
mZZxj1j7Zd31iSI1CFzgo0SY+CSu/eFj0PiehQffSqJsbWEwfpcaeoILfcaPk3SS
oja1b88gt4Woen+SOIinTqfyHGgYA9N/2TRH4pCSoKWPt3KhQk2BVwr3rBy4k5pp
2K+x2C7M86fF+saKyD63pj5aORDAjJnMOqX8nV3CbKUbbXMvihtM+BXTlxkUyhGp
HDvpZe8aiz05GSkX+rcSXoMjQd0aByi79DA5W4TfVU0gWb6nzkM9KqUdWbd6N56Q
GG9MK5um7v0Dk1YY5DzVpwR6gfttyVNQOlLOoRYxi5XpV/2KZfqzKpN628EspQMf
p9UAald/HfGvP/6LDrnnnjZld5nno+wy9Yt2+77K306H9rCcthBMf/NLHGWOPuAG
B5ChDKK2Jtl3lCgReUpLoUW0HuDN4eNcVWVYG2b4f1y3EciD5H7Vsl8UT/MblX5t
DODjHzbNLNU25WXguDdDZeQmmyD5B+jOfXJ1GMiGQi92ACWL1bogVyHSuHnZszqa
KsvlFuxxKuT9PlqpoVjIlaKmJd4lsYJ9KtfFj9auRlc4FmD4d/yHhfeGjZWzLe7R
`pragma protect end_protected
