`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
Ur0FS7MPmHzFtAfZCi/mW0MHf8lm4xY4LmQwJcWvS+wzqwMgIE0Nopv/0AzKpeo9
y/FigAtVFKP77SJdzPivt4CGYhi4s0jYVLAV7SqjWTLiSqJpDB+QMngL92eIcWdB
BXH2r4+9oqMCbMFcP+97u7MXw0CCaLoCFD52TzKRa6k=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 2992), data_block
P+DB2MrCjnek70xItGVMS/N3AXwcpLeThYI6kExaYQk3usMlfU0n62v8nPmm02GV
XqFLSYEfnxqU4uwHHZPepFvgr3x6QeiCqhcUY9VzZzE9NwRboZlGlgx31yvLF3r6
YuF+iCXeuhqN+SERUDdo0bnVWtR/AyjdI5QgVYua33pfvMzPA8YBkmoijE02yVbn
efUfncA9wH2AGzeKz6zvYrowVxo7rJY25pOBm0kux1G8tcn3E8uKhHWzXug9DlUR
N6kS6FQD6eXpZdZg3wmPx+6zI56xKkPzRaXNOrc6jxBenS168Q3SBgAArXMnaTKj
UZNQEfKnH22C2Ppsnom/wAPIgBDYUCAn/MiN4/e84Es9r9r3zmjxxZFT5jtDJAT3
rkBGwt3va8aikqUncltstvq7tpEO8Rq/+EOLLMPqtwhQ5z8P7l4WqaHQrCTlfuPY
L/lf48hIHFUN6g2dWq2yC4/jghU6Yi7K2qo9x+GahV/d9LhXGz/WwPboLO4ctlBU
VId67v4xTPwPLXiNWzdy85TD7Nk0QJKtuQX0iZwQaihC0tIOEtxPM0B61t14aaQX
ZlnMpC2Fh5uxjGXnLhtC0nmYjQgVpL/jLex+k8GK0JpRPW5p+KgajXIYlXEAWORd
FURO1KhGfNPzB+7MQiHpy+vGhBy+9Hi92FFSgOBW89i+FOvazvjY6DZf0NdQyT3n
zacvsmt0GNazhna50bL2dP/YqctQCMy1UfJ7zWOP5lMb0r2n8Uge/qosvHrkUsKZ
me4detwk+fLWv5eEq9ZdGGXIBaof+Dz5fWzQ1mo1/DY6471VOeAFl2NJ/LCff8WM
Dsfg6tBFdLIxBGp/7LCrhxn+lhFVKWMpiQ8NRl8hDZ4FuRw4SX0FIqgGbS1/mAgf
+7Fi5lmL6Vfnh0WytEBI8mc2Cj+OgVqIm6UmCBMueNrU1+gI9VXT58gMPH87cBAy
dnKZu36wjsTHcaPgw8wDGhBUHWO72ttz2sWMfaiV+0Ix+AKYZRiuMdIr3Gdex8ff
fmwxAckUYR/z0QZklADLrsyiHiVzwtWMYLFjfj5ZY1YR/IYQDUGMbOyubYhbEMdH
L884g+PUTnxjHMwXYsUU+pgVkgssoVz7C8d1hZjLRm87avgV35TMeiJHcC5N/9Bb
/GNPnx4uxJOsUQ51HEfygtfne0ajv//MrJ3jtywQ09/qfvNrXILNI5J+wfomhgmJ
YI1Ysm+IPcfYg+1Du9YtyFpHq7cmkrLIXlz9g2oSjw8W8T3wTT3rO0R0znFgmPqN
5D57ac2KCLWNHS3/+tQXLJAMbEhIiq2ATnZYa9NG7omiufNjpxD8VEDuBKu1KQ2X
hAOusrsW0kTJbFsvvvXh0HVMH3DK4a3Q2SN9rDeDgwb2KOCdWucG7kYS/SfdyPoZ
UGCaEyVxjjVK+bvzXnp9MGJeAtWa3F+pSx3fRA1BBmO2S7W4sbzgtpaFUezbul7Z
OE7d7vYGKofDOtRuYlWya1n8ASO2VSmOy0AQ6+N9W0k619J44YGgOthrMdjLH87S
cDuztCDl0tzz2D5fpFuj18rQ+6nD/OCJ9nuKnmKhC+YcFP23dtYA4VU/76wg2Ogk
wjlAJZd67q4aAtwu4vQffvwbtz52Dm3J71ZobaB3u1mPILOIFxpcnly4gqrFx88d
bqTA/DwEv0t74efWdObCzq53Vh91QmMh77ZOx0a6tLpPmK/eTrxL+p0hjK+W2GZ+
4wvNSzWdC1Jo2A0xQmX8Q66QNGbc/U0KPgz3alrW93JeuXHLoFkx5FvuaHLY0+5o
MXG2QpFJZ9lTSqDQUKk0lvt78lesmw3j0X6UDCLRO/igZ9DeLK/YAq9CL8+s9KRW
VCziHs1ZYpTJj7ylo2cSRO90nU4H8M9AoMEtDRTXlKmh4RDhhe0ainVfp1pR/v3q
wxg/eb0bi2vNDO+aH+F1nqc3pT0VJV5VrcFPZznTzKf+3wZVDf0nBKDYmXwB6w7x
tHei4Ysr/52He/ziFVvUqm54J+KCtn7JyACrelAMovdl7ZC/3i9oZTu6Gx4mn90h
IlPqFxNxf8Je/y064QT7PhfHVyAkl2Gq5CJBhhjfQOW+6K5GtEDj1gVjiXPwKE1f
O4voMgTqrKlkYBUwpm4it2PkKXM8JM39Ie9GiWTVGX1+9TXFytgxI4MoxU4iaoRV
J+pLXIrC7ZMjUCWmn+5ZSKin7bxg/1etVKBlN29X+e0RMbRezd/vsxVLuuETAP4M
g/FH5eBN4XxJhu6UPlmyUYEjqRuByR3UHEW4KohePjkdwSp1AWfPviJuRQUm3tVX
9GCYu/fCSnZEgBAzHD/Ti4/4JDB7RhUGf/rQ31gyyBnHfcSknbKeO8/mIRSDP+ft
ZycnKHVth6W0eR8AK4Z6+qZCcCrQM0TXIhNYLE290g8LprGpAesNqiPr0QNOKToY
t39rvcnpHW25fI27ACJXIGETnZTDr/GQihPHYAFAdKF/swx2mSUAjmhHFGJWC06q
GZsvuKGgk2jEql5kb2jJ0yApHd3n7VUIpv/e8KSvqOlwrgaQUty4Ms2BRLJzKchM
Xpb5rNd2NU8vFuq0yUI+rt4CAdnjThh57qlDxEtBFoEbihLla3ZDdjueR2FZKiao
4OYcO8vIRSMcMbTKifQZzWDfysLOSi2rDqW4XHglEqgAow682c6X0cadbrh8ykUR
I/Ht6tNpUXL6/c7NpHhIG3Pk1GmU4PNQy5FTzHyDOIoMyY9uFEffJM1CYLRviiPC
EthM91N8Ez4TH12ZPLohM4qTIdcCi4805Fod5r4GnsRKMw/HVVvJAlYx7LRt8FIF
UAhqGcaAxr8zCalPJoTnljQetYTNLrb3QKcMREQltHuUkiuV8MHPl3tZPicKPIcz
U6rcAf7Yi+fenvh6cS8vjECbtKEim8iKMNfVg3Xy/u/mMrkYMzkE3JEpUteHTpQw
IuJl5PiKEdaMSVGbgzessD+elfRVqFaffU2rJC9p1prXeNFkDiGMupWThbj4J4nY
KIR275cYTO8PITEGCSGFS5+yLFiBusGDbPGDLbaK+j+bcur0YJnIpvqTslKRiWZd
gCAMRP+7Us/4HbNDDNaYkjz5Zi56EAcSX1Sr6RQs2KEvZCJpT2npkFy2hTRTNIsZ
ow3EbOVhK8dvcvktKwog2I8c0+XuGY+qyZ1W+bwr1eC3NFM9kMHks3fjfTN7WmGo
CmDxutHaxk+0SSs8+aVUbnBHJLqbuNS4gaPeKvhd3bk+TDlHQhuOlJfd3uNofyXV
D5m0efNWPcPabwappVfu6FXlkXEAu0TqWsjLTVFZ7CmJrodeOU0lwFAchB8PtWvf
bIUkx1fAa+k+pglHMyFAkO0GYSz5SS0dwJYwZpWRvc4WRcSRClZtgn+ronV5H9Hz
na8Kr0q59+mDSVSHZL2ZJxQC26tNv7mG5zB5fwHA0i3JD8Q0mASfM7q+Duwn+SKU
IoIUAPjBUw+BN5A6XXHaLxosZeoubdMYqETYyLmBvEo7nwUXYlMiOllWo/cetW2J
lZUV5N+rNHihG7Jl9g4XxWGSP0xw0bBz3/LtAN0CC9YOsg7xbDuUuadxwa46OF3A
LmMXzKWXFYsfe2Lgz6TTRLTLA+93WG4GdHDc3YGgLl5Y9rsBYOv1dFueWlMmDJTf
syIyHs6qtWKI2MBynXKt95ot5AtPJ/V2bauZknPUOZdJPoU+5LhST5jvjRTwtAWw
mGng+hQhPEo/ZTV04wqAYIi3MpMu2vTCTqu+SlfCicoDxSsH/daZqvnW7fEeERmu
qS7XJouI5MKfuSdKGlVWLmHqr3KpAk3GySP1EYDJBsfWWt8v8P+2teeXWiP8BQpq
F06VA/ykt9kR1K1aiB5w9WqdG75YvOImwdNp0LPNUF39IF3N+WO0AxN23oHnbM/O
6ULjH4tYgdq/w7ExnbdGmtA9f7frL4SJhXxURYy2O36+dFg8FK0IkEoM33b2gPUh
1mEYO/F3gcgPWEwPN/DqGg==
`pragma protect end_protected
