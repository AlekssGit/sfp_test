`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
VEcl4dBNjHvy8aZYXlo/dO5iT8ZIDfeKbs5iuKsFyy318TKHIo2UE2l/u7MbhN3s
z7rmJuUvLchhNvMBkrRCYH+Y9SYyye7eKKITX+/6ls5N5P1lL5rwQ5gcYel5+8t4
1R2l/IiaR4pcPRQFG7rV9giJCgM8NFs3REEbpBWuRgg=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 70496), data_block
XCjuWo/+exKh9H6RkNoZCVxycEq1uBrAwFyJ1yMZD3Po06DoZhQsr3n24109xb1H
gjj/wtvNtWkjVDRZPbzhEQmm92BUzeB41hZ8llNI7WsGrNX49MpZ++E5upOKimT7
1CGYftYph3RugnPRPzsbjrvxA7a56+NrxQRn6Qhlrq8NCmmaqcnUXNf0XtLQnjVZ
N0t/eWGapFTUzVsRSPMw7IkSyi3rtzHlo1v1stipi83XbPtUQVMB586jwTj6Ss3Z
dOoCnFIB3XwdVjRxNp51Bm+OR7wuPmm34JFdgk/VsK+pjW4YhDloNN61nTIyADI+
q/BCSm1W9U/iMyqkPP/7WsrukfeOjTcR/BeHvDWQDVD9JNelBV8pMVsAMR5gPihK
Zlw+VxT+DtNQjInPZdPatUD4Qd5T4TYanodkX9r3H34vjM1J8HYFF2Nufb0S86vF
XjAtSo3yLiBqq/Hgvtf3bJEXOER8DQlgW3xuQbEKTaR3TJCjx/TdfOXtaja1f7oz
vEu0LmxmdCgAGCHyhRbFAJhZDhq4vDX1LAgYhkmyIfD1MC9WJH53+ktUqVkwNcVB
cbYY0N2cpfQdazb8ptMX2Rwz8M2Pvb2MiqWhUmCnFQMGW7xMC9Fc90Q9uud+W7iF
DvCBOkVn2lQqIj4bOiuYvBVsVt14RIDdK4knv+Jm+au1fK6wzzPP/16Uc/xZd2L2
Vwgk4ZCM25euHlzcl7Tgy6Iqr2KjABlfserKEwej87FuO5L2i6m2yAg5ZteTMARO
FRu7LBqM7TDFrPWs8pomB2AhhCMG1o7mR9cWMY4DIzfpmBqOZdc6RSIu5DiOB9op
4V/vQuJFxjfAhVigctXvKpPm6t4QWNq60ivB7+U2BKHK00EAbKLqkk1EF5oiQROB
SSx0sU+kUw0Vg7gyT1dEpw31awEiMQ50KldQ/a8A2hWPTHYpqLO8ISElOpsnSnfm
D6yLR9UUt7MDnXpZ4LdjFUpuefIjQVuANuBe8a5z9iAnd0GxwfP9zYuHy+MPzux0
Xd/JMzsP8OFI2O2AB4Yv6B/LTVogRK/QRAaCEOjz0oE7CvPYzAyJluBBUfhzOHTO
gOeXLq6dzwEU3no4X/ThzaWo9Qybog31YEmk/SS5dVNLYP/8acTn7GWLp8pyZP1M
YrULJWb29h50nd/mQzcq+OCEdi8kaBM8X0Pz7RLZyhXG4tgmI1lCPpqw0O1DPKfy
uQ78jkw4qSlSNaS+6Mcie4oHxJ+R/urIXXk+O3mHM7+JoQhgwHTUR/hbKODrV9VO
fKf0JFFAGVtjHtGph2bLDa18VQFJs+8yPs6bQhfCJ3QIdc9Y7FJy8T7B9uwds9Ph
sdtESYBwpw2h61JIHmGI2ulR4d1JcWGLdYm7dLeZPWA6VcxMIaUffN5dD8U19y9F
nbJ9RTcos5N4+ScByKj9JLCENAK9weQm/sZc44HUOL0QNgpbr5PVANwDLYiKV6A0
qiXLqSYOJ2Q2GmeWPYD7E006uewb7vjqfhryovXxX868x9BEnL0klV+TcwKava7B
EURb8LP6KI6ub4hHne1ZDvNAGxec1QKr/IBTyWBk655uPJeSb2Ah4jNyQefyw2ef
8CRA+DcNvtBz9VE+kzwFUJ1xb9GCk6kap571UyvbeQuDp1WnDNUpPidsVOzxGQ6z
xSzKYf8YsjbsLrXmDWUiPenRvw+sAR6if+it8ZNwTk6ITQgb382UqfwGIi37G8ty
9feoI/JyhXZCgaLlxpX3pD3K1r1C97o8lImMRDTHZtNS5+CZ6/V9m/K08EIGRipQ
ee0p1+KUkrhPypISRD0bdOcnls+WCPfXAbzvDu8zBusmSFe8+5qjTjgznTvia6kn
Yav/b6tnaUbItLzrnz4yBLUizcPzNwYpNDFwCwPwyH3z80YM5SaO680++tjAIk0K
uR72gHe7uonUafyvu+9M7KlHtp5gWXm5P2OxJyAFA2pkM6uVWOT+vCPfTmgzcEAg
G7IG5eJaiGy4HBZwKrPLvFkH9adq8mqnnPOyTqMqkIzo7MxMl5M4VhTo5h2Uv6j0
Cn5Rrt0qx2Ct8Qr7RvthVC2h1wDUBtIqfP5MA+lm/mFBBAOLv7kE2xPgVJzPR7hb
G2Z8m2IPvtnsKl2wzfewrGKaNHu966lmf1P5y76Y8mIT2Qw3iSDdoFMUHQbPVspE
YJkHOcduNsqiqpvVEGuGavp2tSInTJzRbM/F4hJ/P8LceAmIZRVnH8RGWGw0HG6V
u9LAn2sYWfCyufhMhU1mLxnqwyu93YxQyA/UP3ymNxAvyd87kxy4ByaH7eW7D2sK
Lr9f0IQ8agGToSFHElfwMpHT5dYuGcLbymciodPeYzXsG6MPazLxc5zcyBz18jtC
rTzOie2YZ30/3CwdNxr2FOp1CFwqISp4WnWpeT4xIf/kawk3t6+MZEZBnvxzXUR2
QoithcGtoZ2cQFTUmXPkgh5wHBNkXN2kfiw0LnLQzirFHn0DoAYXcegPyYIlmbu2
+p/+nJX/WzYE4osfAS8MP8sjLPqOkOmbB6/9qAA2u6ocXwugnWbnk166hynoq0A8
gBkdi6lqyjLEnPzd0z0McETtMHMSIEPqn3ConK64Y+mA/jJSy/d5ordb9PxeuXyP
GR9RGRayJ8czr2jLu9PpPX+RLZ4m58bazQ7xme+kQH6NtmZaXzmyBqtU2YWpA11T
wNLhqveh2oGXQDZK4QOCAnA4JSMVyumq1jkqP2sWn8A60ESA8+hU/xT1IPNOwqpj
LaJltuF59nmCTBbqbBireQ593lTwnzdT7uIQVVi9H7ThGNlW+vbHnrbuCYe/bamI
/3QxFuox+jSDs9Gejhzzzud/+6OwEac7i8tXN03fvDbG81C71bSpoIku0mM/6PCX
Xv0D/AM3FdYm+vUPeY4pDcFK6vpPfEInkaOMLon2VEA9j2aTeCAO7eb5Z3bBVeOV
UrggX2F1Uahzf6Wz7dAJZU3rIMwLexQUJ7go6iJPO098hqCoR5WhPm/2MbR8lSfM
m5ynWpT0nAmZuxPqvF59uZ8/+rpALskc51GAdcxd/rW56CKhwtzzPcd6pSIRbwGl
zPntKsXt+qsB0UHpHUVNEcT0BrQ+FUU+w2ij2nyaKAIaD1KdIxl51XHA09cV7jcW
YBYOtLxZwO9j4Zt9eXSXvqSbKLXFljyT/Z7D9z38kLoHLx/yx8aSfenwbtTghugW
ur6V2KoLI0t/hw+umB2/RHmGibLkQhw0/1wUqzRoTfR5ErwjgJtZBb+wPhTx9/PB
rbSkMsjga4Vs5pqr7q1WSz4KBVhPs8zbb/9b6b6mqsDZUAo/32Bk3znKBUEj6y8E
yj8kerjm2JtDnrL3359BPzUtKeH8iMaMmT0i0Izf944/mV8OSl3YbIPxMMzjVRz+
tUnJsj9OkxGMbM9bxG7xYUqSXMYXqcdNod+FZZD+vYJOacFM1QldvRl3FBZEwk9+
M5fwZu4w2mpOmpKNbsA2uuOJjyTKNIImoYiP7oz2rMQdXgKaP2MwKWD9YmPxjKEx
iq20q1i853nZtZ7xXt5PYsK7GBvcfJQ50hDyaX38Z+u4L+5/AmoXKXKAQcLefqJ9
qaXlTNpHciEydi8JkduVjyp4iOGLMvIPwi12Huc+jgKfpSXckO7rZoqIo7r9XhKv
y1/Eu3sxHp+l5AYUAFiPAzPzJqpSweL9kiwBmKcunm52JaKPEBwZgFLPqu3yHZl7
fGKp86pl458K/Ty2XMa+V/0s/wAfDISEFAfaEzsa79HVtAmfubN3z++WzHSTIq9j
8n3rJMafHHGidbJI073GO7JWeIouzYdAc+PjWQWPb1kdIP7/SIiGkUcN4zpHIPUg
tNi/j2rY4nonyrG+U35vDExJ121tLLzIESrQG8NvLj/kE03J+hWqt3kVn5FJVz0F
NnjlpgQUisU8i7iJ68rcXJ4AC+3N61rqaAkWHMIeH6ljS3cVFqe73QbRwZRxtGk3
1KYbdbdAg1dc2qNEjV6zdzRCHoPIwJ1gflPAP82DLhLpwj2Y/GNujpKh4BrTTZkD
LBPaDO7jmSvrPBnMHNKTnZC24tEYwxQ470qAC3V73HXmzzPL2dRkC4fR6lidcR76
bUlli/GO4pIZ96gJ5CWVGbstTzS/3KXCz/YJZrOvKuikzN7t4KMLoY+xNc8E00Mb
HrBQOIAlLr9JWzapdd+uSRirCD90d+sRXKxJQys1YGc3vQsXXUl+e1ljGnGHAkF3
UuIi64Jk6LVSUXAzOGRRCF/7WqeapKihMzNG1MMWZ+Ieig0e24+RShz9VG6x0qOn
HbKLhaTZJYvEf+ZHaupOCuWuzbGlAWWzDFRAWW8bj2EkExfB+hxWBxAeQ4pIRhJL
sip0rzlef91WxVtSjt9YmHKkiXI9HiiDkjaHL7bhBH5nSUkaOp2DsaY02ywoaIJ0
s2dMdcOncpGZ0W/Y8z5aHg2gq+vTcQ13Ef5f+C+0pwnU30B+M19S6PEAmACwlBg9
60qawpmNF8K1+S0AintfgPlw/tuvVuryiIyRJBh2LJJZnuTn8twpr3xVemuPTHL4
vu8Q1Xm3FuL0XM+IZeHF5xnE4mxzsLviE4KB1mhyN5FJHKfd2xYa9ngG0xlHKzzG
6w3ka3zEjpAiGQy03dOh46020vAu9FEk4d/d1+78tucnVnCtj4fa0hI8fxe9Ygq3
yFVv/vWlbDHDpeQtdU6VUNWkU/lL+VU/kethVKuYK3YruEOoexKHJU3X+z+m7/QJ
DUbsyNuOngKb1Uumbcj4w1W4WsnAgn0wxO7OZEYP93ZqJif27RKLctUVwlB/1m2J
ZWahP4XBSaIWZqrXJrqYffFh9Mzo1bbp1QYxjnerXzXqph4TYlyGBJaoQjD0gJ/o
2KY8uFo2qs9Wl3xxs7FGQbYgpGj95s6LEd/a9opUPpUTMTOraKjDSC8ZBfZqPigD
bMl5xN2lmUETLwEQSq5G3hfbYEuOwpJjlEYGIsLBCdR3mAoFbixnoJDoiiIdu6jB
VxM3gZ8VaPFNVRkFVhurQt2IQ+0IxY6ZceWC2wJZhOpJbONIQTQCzdaBAJ/5iTWH
JVoQV5TVMvJgoHWfpg++NYCuWSfJEg+Ls+kw9ynZsfyV2MzeV3FI0azQtYyV0/dH
8eWotVrfxVZRXemHAGf9gcl6DzDdlZw4U9rtDB1N40YLXbobrZ9cEA0dli4BAsA+
JUG2WdTnWdzPyU32iKylTHwWDdf/cHWL+3XtmI76xJbCm/GGEVJ4bbX8HF1nogGC
U54Cdup+RD19eGg8MobvOvM8Eh+I/QoIUt1yPL/BJ5aaVCoQ4zljfEV2sHehR+5u
uSSE1bd83k47RwIbZSbfc49CNmGw/lrUcCoaMf5/MkMyosONoWsCETcJJsoVJlOC
MDItlSrNOGB3EwmPdyQj9pqPRAGthL8zWhOX/CfI4UO3dCKmWzh/Ikty53SEHuQX
1ghWWcSG+F653uvYZdYhEPpb0tazDLxLpnqYpO9xG67VaFGGngC7JDMCLM7gLEcM
PuPDSbSujUedhYi3StGsuHnZ0BqhIDBNb3j0HCRITp7FjjpC9UPFo4Ii8GxbdJeR
zhkowFb/GOdyCqZS/+jMXi6x/bardNsXabiC1L30+ob+OcEIMziXwCO670kE0vfZ
zsX513NGBT9XEDt7QBNkaSgEuMO9j1o0Rtg2CwmgHDpFw+NlD6Wm8JIfA2p387WH
te4pOar3txgvZMa30409FC6QjIMPYNdR5uAyokelhYamB219tqEDCq7qVvQIP471
CoDHmYvLSViW9xfjFzyC7ibHTXtYRH7SBjeoIrJQ5rEfL0UDTao/6t/SnoE6q1Qd
4BybSF3rCPXalD6G9a4jIATkfJFIdkNXE0ji/E1lJfab9bTw4tdzbdyyKvk8GYTp
AJ0wEb6gI7qTIX93r4ZfxIVdrW0NtJPXQ5YFKuOVkqeP/gb12ArZ8iQZRCFC3EEH
ILbQg+9F4uATULUq793XTO0ZYVAYbhRmjsD+ruEauhOMDNg8rG86BBwaY73jOoWC
sTGnqJMUEGphPF9TpRA94LRfYNRCP0GUoJlembcdPpYgK+hJZRbLQReh+W/vwhxB
Cmdi6gkMY1C0TqF3BCrTgBElcRUOB/T7nCIxOqlYLKxj8r3wFiH2zoWHG6pl7l9B
WasAgvm0ugvdSlBpIoxE0SNZQacfZwARlJ0qu912egoO1nA9hDn3tHqpKmEgeQrj
CQ3Z/S2P0dE6aUePVtWhub3akgjXcS08tMrXMO5yJIik+m1coJs5ojOas8d8ylpn
G7YQd2/DOr2D3lC/SCLrl2PC0bzJfbea3HRnfM8+yx6qxvmHEfggrrWdieSnWUfE
XRuWOSO1LyWNN1I+FUX5Z+k98gBBfYkrrhFB5maSrSO0XaQokENXSizwiSBesmHm
yIC66MRaWAbvJsUUHZD5xnT5bivxMBaShSsAH4FGru5+tAcPonB14N6R8HGhjcRE
rtP9DhK3PDznNddhKLwW34nlcfuHvkm9b0N3VE2Y1OaVcgaEgU38uYQxCFUmR11x
rRW4BoYYzaS37NZvB64sYPrYavPcxG/vLrOqV6r9lNGqPSlO3+Ac/+zQER0JaFP5
vWz8fct131NhCN4YaM1dPeF1BLhpOAdbe4t1anUcyAC0HQKEAyPCwoDxw3gb6y3D
3iXY4grMYCBY/wjLq7WyTe6vQl1VBOGuaebPAWbCU916OEqHmoFUDu1X4kPuv8O5
1s8mgs92LN0OzHkfx1v1xqmVAvCDdYnhpasvzt9ypP50KUhQTVnzMgyZL8JOztZl
hvijo9GmBtY3T8l2LfKRltiRgus3ZC3qLKjtnjOFG7KG63WOeDqM40cxN0kGNQH1
fnswz16cIy4iKsQ/B2I+qCFNwV7DMpTDxdsyWDwkx1Su0CavLsvBg0QvU5JtZndn
XipjATAVbh7ah5ckcaXA6EAsujg403JCyiSfFa5OxtrfN9RtAU3pipyQ6GX0mx3W
lEOGsTtH+I6joXYgu/uuvutDudts0Pca+kWYu7MqWT29Sj/hf54yA4b/QIh5R94H
v713uhKqIs/sBRHYjNbd32pkDdes97PObmEGWlY9rIlvkS6bGNq+0b+CnGu1kgjl
fkPmS0Rrskx0Q/GaBOcuGioq6sSgkB/Fa4nVvxxGg+TKIAz/Z2mp09Bzrsw5Jlvf
pMZ4hSt9JjyqMO7JmDVCbSePlW9u8UfMOrp1ug4s9sZi4AUb3/iaHPf3t1+IPaFP
xwZQSs6eF69Mvc4+4q5VAFsfiYHNJO3ipDU7yMeYsyp9mUarEFjT69ZbDdqs6OgJ
aUBdwqGeQqh/YhCLOuaoD7mbZ6mXYTcd/P0z8znZqboOfGzdha1LI4UPZ32JDiBn
vCDthqMfY0vLHjAY+huPIXqoYTTG5u9ViunM6kI8hyqMHOpFzZhC7jGpt/jYRqvC
GoFzjPKginXO43TT34Y4Lcc4FTpUaOEQgbZGSnwJgo3o54CaDA8zTNaeS2MNGTOw
x1ii2ebbmwW/0oPQUvi9+tBlcgbi2K5dcC84LgGbUAv/avrVHO93I4PypdiI/Sw2
JDreOfonOjyYontn6L7tPUabAnAli190l32GRdvRUOMSPcISLdfnhUwA5VUX+pvZ
jfA+wMvzNrwY1v8Ij2MzN8nCeIx79asAks/LccDy45QdbqYLNZMqwICzh9rohrkB
u2ADxMIWmler0T/iVTrH6w6gcmIN1ssUn9AvxlMDXfDjdGXg0E/yZJjl5e2Eic4H
70he0qHcaLTEJh6K7u2G3l4VDGPeaE5w9l7uVwOkV+YfIW6Hx7jtI7gJZccoScm4
DTqiQCr5f8NoO7BoPRUKrd9N+9tlw2vhNrkJ2B4zvbrUswZvg34d8oSNHtZUb6Vv
kHmKW9ojotRQ8Ap8++zShRwWAoygYZQ29hHOzOmmE9KWOYdmk2twzY9Uuujooqj3
hGUEyvpF9zN/vfV5KOU0lR7sUMUh7QyPpaBw8HBwJX6mCJ+BpBHN5VjZQnogwlpg
YJtjSCRaomQQuYTDDKvq+2Nnwz0EoZ9Up4e7ulx/RJCQKayazj9RxaObAEKzuIss
drBH41gf069PRslK1tVV8Hpkdi0LYk0FAEdyy+6czxnoySMjAd1lvBtvXNbZTtzm
GoODkcaIpgFOUVrg0CEKBLO2zukVKYTIv5+QTwJIGfXvkSfQE+N7Cp2yUVneHE7H
Q5rHVUPA2OCl3SDCTshkmjs6Z/6XLyDTgr6KrQD5tt+6RcKWHBEEikQw18UGSThj
imdsq2XrPyImEI4XG//hkqLHZUR6khkBz7CaMoySXDi1WQMjtrl0YRdUX1mcwSUq
fdae2vIY6Jai6sbofEJduXg50kae4V+F8nx2HFolWjJ3d3k0MK4AEbpEGJwmowsf
EHSyASwX1lEopyMEtxbtC98qoMXhj08OpOU3KozASaQOcbUBtqI86mz5ZaVa/25+
MNTaAQtwFfvzv795UzCfCK4ky6NoukpU0aO6hWtK6ylYwEy64rvlaWeO4q4wBCzI
rIlLCefdOa5E+2P3LeKE7awf/JVOsMhvKpIEnYVnd5hALnAr14Nf9+r+jO2NRN34
Em0kvlbZIZ9IZF8EUw9FnFi4ZNs6JL3M9YhBZ2HtaqaseBt57D5pNWsCY9s/oEQf
9aVxGWVuGgiQk8FmbRZbJtSVrRjeyaXvfD804WOJE/ElbQ5ete6EOCppR7l/UJLU
k8/ljuYKy7ldzp3gjcP5d9uBJEXADv+sM9UoKMF7R4QL8R5f3De4Hz8b91aOth2W
f7UKEixlGI5g6NOcaB3EK8xgr2jsIyPpHooaFNF5kzGiWeDWumwsYMQ3id5czIDd
y2NNl0DKxGiRCNrPv6Gan2ve4DvQrZ5qXZI6cbcmmXS49caqelE3vc6Fro4JnIwB
3jp57prLqj8jvzRm3MoKjhQ9Xnyhw9GrA8xXXlTpiJY3kjx/Z6hHZB9gY1JDRxf2
G+cg0SKdRY11akX8l138QhmMUjpVUNu7uvcaMR19BeuH+xPHnW76hNpwY+nBzARB
5F1+jhQ/u7hmUQk7eL1yH+vpqAIRd3OBJ7OXb2BA5fbIerhgiTAuKL2hUUm+l0Bb
Dn+vvu2oq4Lsz1QUdc8EBfyu7hxivCff4mb0MouB+UEUl207+yorxonRYUlXBRdN
yn1oKvsl5/GZMiOQAYwaie+0SjdwHPm4yzDc4jiFLE2ddMMw5tpRVUFd9mceiMIM
wunpgsi95DOOkcuzZpofzIBrfQEp2ihejdQ+J3fsC/EPgu0jIZaRXjx9++PuuSm3
C9pYUIdmUIQjUPBhlNmglH+JHv26BThA0RDPgtNRjG9cETQqDtgq+GOqtRcdwec0
jeDu8C/t4W5R0f8aff0zsL7rmdFHcGXHNSD/gEgtlFR9AnSQzNmXbKGXvRFazbE2
zPA4cldeOKYhDsWQ0fijFRcJmYtaZ1hUWk3RdtJsnDUdiuog5JXao8TefFIAQxhi
gRrRnErb/5HLmOEZzq+zT/UgcPvClGujHEKsgATNKu7GNRRNFmH3k0YHQkpqB4bP
moANIDuk7mobT//N7U0y6ToC3evLihDW69L59CGfx+J2LubmUAMfhGTxhG2uWegm
Xha06Qf4SODTKdp+Z46UqIgS+z5DO2vqPBrE7U+yWsvPL4zHZkr1BFctpEdD+yz0
hN2fKDuKcGVR4ix9R0F5eB0Loc77Z+gbOoRHqUY7RENKGPDTtAxTazkCpB2fhBKt
Q6d5DwYCdrdF0GI/jKhmTR//oTCB10Z7cIsQLri05Ufn+Bdus/HSV2SbPIMdBuN+
n23hmIwTSzxWUKRuzCMpFb+/5mJYGRE/JLva1Z5kjFiWZfYcpSRz1GsFIB/OTARG
fpqZLhWPQy58qFPIQnI+ie/V8MTuqItvLPrVCSCMvdRxdQV1IWA2aFbEeSvmS+1r
DAKrH3WgvebmU+YXJCpSUkJrw2Qnrc+u4ysknHS8Tap0RhqqE4kB+OSCBNPxRwOQ
ziAzUGcHSAkSVzFsbR0BfXM/VjwAuQ0JqCsjshuz9uxphtrtzrrGGUyIGHqzs2Zy
VthwfnOnA/guBoO18zvzojALdhpso3V4fw1d02KF1v07cucMYNIoprMEt0LfpAwy
gbZaXiG479SX6t3U+rxjW53G/lYurMYc3Jxa3fZhtUNuRqdxDKuksa4l+tOy2EjG
GeN6T/Po79cPSeWpEyNJID1beqAviZxJLKUQmCmBn1XoOR3Wz2G+UF4G7cyUbOYQ
SGYZP4PPtVIK84bWG+e28F+tabY/xMvhktymSdrMZzwWR4eqQ9Z+Ea0o1gEHM26E
8Hpunmw8mk6aDUtrN1co8pDfeAggHbxzoNakmHLmmqS0fLGq0rycUDOtzsnBTdus
ierJQXvyVeEbRL9F88FqczYSoKzx18LqwM+cIt8U3fm44SXsg2PCQjsqcHPSwdb+
7Uz0Dm2hvkBADIFA7hXPWqtTSpDMdppN1qzMXDoYDcJEbmf5iTQ2RdkRmXh05S9i
AAaExHjef7YLCgnwGt0PFNvoH0BBhYSYitVR2xEjEIbbCW/WhZpQUARXNKI4T3U4
PvJDLGIDX2GV1zxxRfkMxZ2hFnj+E60HRbHA/9jknAUIkvYvZNaR9+M8VhLsefHt
YSWye2DWdi34CQ8eF//UbiF2wj+XI5aRzAYM1nP81gdJvEOmIvlaov/grLqDngdV
72BKVQoMKXloDwi/T6Wuq2nA59h4d+RFOkIWVBWJJhOypGkUgy70Ml4nsVSl+LVI
Mo7R8CIbFv4pmXbck+Rd/5aNATU48u7qmPCSYj6r8UfVEiAnVqNYRvIDParM9D6r
1IcefFz4r7mTkOwpILUNly0piCP+Nf73L6fR0vSDO2nFerIyoDaqF7/QzR8VxiwX
//+Cd+QTr5xpM8DuPTGm0TajwG2ZObOeb40uCcp6d0NsnWU8QaMqfpLi3q8+QuKq
OLmopsOJsBz4/V+sspX70hflfzz7Vj64nSk8+0r6BYeREDa3u9deUdIqZxHgqyQG
zUGVCXqXH9qJiZSo1noU6FRVhiMKbus02Lbi0bcn63qKU9mvlueoUf1dTJsz+TMo
Njk/ZPJJpAt9varkwqHiL+wssAhP69Pd+6wvXX2+RtvTSDinhL/Nt9vQL6Y6zJZR
EJQsa3nb7Sjar3wqMYzRtjAEHrxN+8wnW5FdngRJUd7/mADnvJk8mn8rIZSxTTgZ
F+KtEdfo3f6nISxnfb1a+WclDqH5neM3bT1rDmcgldoQKLknhjPblHiODE3tbQYq
1dJyoID8O8UmjbBq7Y+ranytiTCKOflZVac+Q3zIaTz9B7J8qLhjlwVGh7lYRvox
Dg1JT5wq4z+5GHJ3C6iVTSmjHJN9A0I+pSFZrNI797o1P7CLjKqhmT37tInjxGWb
sY0txCiKNYTAr4WqsSNL3C2LKgGeritudxmOPhQJWq7yhx2VXzy6xXj9mn2PY/3f
KCPmQXKOyi2l7m+3uiRY74GRd7svtdxRVXjoezcGw0ntIJGOHSSIQBECJw7trKjq
I9o1me+gMxJ/RaRCgC85xqkpPqrUNRkUkUPR9T5JORLWwvfDXKk8btYmtyGZgRDC
IxK6y3W5rpQ36xsluGRkhXSgIqMcbU5zQ8sz1H3V3skTQbPIsiBYUTPaX/HMq5fx
a55gWyQ09PK0kcc3KbP5KVzFwRMd5cBrY7HUQnBfvLJRH93IeGBbKbEu5dkXG9tS
NaTMO1P/lqu1uBtT+4I7ZsqyCYuNz5tX5GVF+ZKh4I+KQ8qdoRBeOzpzgg0Zt23e
7WRNkIkX9AyV/fWMCRkqotlefPD3YbVKJRhC1l6DsT5/+pzRp0gK/FDywGubLUgK
nayYqVXrJVttqPoe6+yp7VqccmoTEyKLNSiHWZIk5pXXebBuj3hV7sgpYk+93jje
zQJ64FR5BToiGgTiULcQCA0JoKuKbcJp0cPhkyQkB7iFh4j8MNI2V0HvzKTABWTh
RemTbXxPa5NyN2f5opSsaO/SUsaW4Zv+jl0QkQ1dbFSNoZ5dGuI+xh/GxHYryD/s
5k5JUTQxs5XChnw72avhCo6eFAnt0hST8yWVAx2ZOMc8LeOJQWImei2/IIKzL+Wv
RKKvVUkk86ZI+C4TM1Y3TZlvORANeJsLALZIfl+OIUaqnfkFgmb9/Aay645OZvBF
8ihvweCE7U9KWlMDAefvKMi+mCipw3VAHsAZutVQJs8Q39ql5CUsZba3tF1I3YFV
Y5uXatzAMKSjyK/oUODsOmoFNy/KfNssnlc19oFLfUYy4Kmq3k93iCGQXXN4U2to
ctiyePhB/szyqkbg6Q5fbRkRBu1Tw+zKOONenMKzIenxaJbYdJizHFNGRBLJTz/O
eFH5wZ7OYBh+eV34tGVR1SfxLcKPA+vz3hhfZkL35ABAstSFN98VvoSisenhAVvM
hijeWhe3uO+D2D6N/4K2Lu2kLGphQzpoeIG0qH3Ifwy7SUwp7OvQPrJz6TylTSlW
rjH1KEEcIJqX86Cze93l1MNP6wJ9r16uEA5PdJmxcYv0n2IN3ji03mGPanWkF+x6
2/v2EkZjoeo3VqTazYxMD7Kb6nH8yTIfcGbN3bXofeAVTieuonx9IJKl1sqEVoon
xLX7IGo4sjFCMTEyN3rpQJdXiwk4SFDKU116a6xGPjZa6JX53/JjtBAL9fP1x3Rh
6og3NSLZ3yHOu8N2ujAE7HVnpbHxjQ7n5nTRbc2RfyiH3JxE2AXNOV9UbvX4FvCm
roiOrw7X9Ls2okXuSO1ZlpZQUbRNUAhFdmvHDC+ups69ZTQiHx9NAs5pmW2vN9BT
OJmMwDgoGVVHuCnZWV+NyR5pbkLB+KT8/t6SLtY2qSEJVIgDWJKtMy6C3VMwS5v6
i6Kcbew0oreR+vB7BvT6Y4SCPoU4IGPEkhZzrj3Hte4+qxPd7rC1qMvZOivEJpXP
02/w57E6X4nq51czt1CI82vVOPGnD+GGG7ypyHm9m4pDooSZNaVW7Uw7c1H2qFSx
i390kY8fISxPI1QOFZr5PH0bPeaqXurucDTLKDKICPLBO33FnWUTLIOw0rCSStHn
K0wqIbDDJAZZ98J8kGbfpoVIf2rqXQiplQRo7YOChNnh0rUex0w1p3IcTsOot7UU
94CClCb/UCQTsVFeRD6NcfiWRo/PebJAIcu4PP1TSny1OunWmam4NqdY6S1y5EPN
RxHjWImOSM3XJH3ZZ2DUktFY4m30FB4SJ71HR9q3iMBn4QK3bKrm17ZV01pw24Dr
08oOrTZIxHyyck3BIQpF0FAOdxJzcS0ugLLznUxoxnlWyJigHHc2zVTU2uTwhyGA
F27z8E4ddnrHDEtusd1XyS8XKfSQRIOPivZrLEj0WVvdYa7FSCWeNYQhAmjrvDwY
AKVASmxuIWJP3/HufgPxTQ+/AdmbWizsdCYnTSdbJLYKMzSfvNgZVzDBR0AQrvPz
0GoMLVWnD7sLOGmo9W/Cu5QTZGTiz6lg0ulCz0C4UXGaD7eeNx8Jwk97Fp8pwBNO
LXAGAwzuHU0/PhpnR6/R5gbJq9dTr7782GZpHDniTFuytO+PdhbQPrlz2u/jr1PC
0h5trbM3DRVovMZQ93IUDHvCbcqfA8lHIoF1Y2zvt5FZ+KQFmm0cY9SQDaQKOjwF
OUgw1C5oZKsbH/wUMSZedk1cGM6/cf7Ihk0PutGSxxivJbMZC3dAlRIngkcoypfK
u0LiszHEz6bGBHAOBxuNPN+4trlvfGOSc/mkI3drWTwIWjAYvv7ST4QKUbyKykNs
Mcw7ke4Jvv2gdL02UvhNgyGvgaUp1I3+EfNmAXKEpEurorMZTGHhSVVLX2lRR55S
DwKEsmPBhmVwkfRW01t6QQDIotner6r+4icdKngRfA8oMM5RgguYR+dL3tteshCk
pE/WMZ0IwYlUwBdPc2LaTGb01ifdNUT+k7w67ctRAAf5gnPN9aI7dcwrRMziIIQQ
tuZrLz6VtU4uTxOpVe5kf1kAe2lb8Evf0wU1ouc0MGOSsOX2Iz4UnVhNmPxFnIWQ
u6SLtkcLsfU8gsdsw1k3wf8MIrDfFG8IBJhUpCzkJ8Of/opJakyyHq2kLSeoQFvE
n+dTzlyPAGMdZ5ksTgCCkOGLYtMx9lkHkO21SzUp0ODZadaUXyOwbDwJYMnnNDqo
cd6S3toiocwhWWhwKNynvsPvXX498Gy2sqOSTIB6AQ0Ld4kd082N03oTBOqCynXZ
+QlwAsiwLSgeh8mpFf7ikzOjnvwUyIy7LnybD8Rda85YtQe6dTalxVCw07F2UTTj
/7Nh/kvT9AdXCiFG7gg5l31dysH9/gLEgfzi4o85rvM2deCm0ZoDglYyh1RcD7nK
cA1UJU8r9rffJgCK+G910ceFLz6cPq4XDnTEJDxfP56vGuvIeuRE2x2BUVWVepeU
K/ZsyNHbaNg/fnJuz3Ip2ozT7hmBUSQp6qQRTKwcTef2+SgM0T/C0McfJRuwUa37
XL6tIqm4Y/bjV6TnN1kc11yRrMt4IOd7i8O79DtKWZ0m6lFstuivwlKGox4JkOnn
RHa4Rp1fojzGDcqoMRlWTK93kYSDgBXnFe73O8ERwGCMyuOofWDgJY+gUzoP0+AJ
pIPfKUkS/LZOaHlGqWtJvCRMP8a+/u7qEZfisaE5WG4NJpLFA86/zxmRwTqqlft+
FuiM2brwB3MN/XEcnKRO7Rii0yK14AmX0mw9IGPG9T5r/P+Fh254jABp4otimhlX
BmaKEbKPvHnvUMdkmmYw7bI60aQpnToKfAsa3nWi63xX0iMvSWTwlQYK/tzRui9s
eVsg2VHhVJY+Yu09NdV9hT8+luGY0mc5opXj8+DL5e0U7uS5Yf6UDSb1zuR06wkG
8ALNvw80/4dcqikfJibfJGqbn5/gI5AdEMWEwiWgI6HAyOTdKaVt1m8TmkC4xmPY
H+V6qD2p9EEba60yIfXFNF+o8LOuUdNW7mpoxSomieyDKvrj4gLuBaZhVztr+MBM
+890VldhEnj+B5r/KEaE+kcLVOv5VIEzwMAgSwSGOhp4NclLW0f7BWko86jClZlP
UwYylRE8W4o1OJAJro/GxvTZEzHNnnk8OjNM4aeQaTzsv4JRFpoPy6AUtRYEBjLX
NH/CeKEF0Mv2uK/CfprMWp/5Q6jyIRSpmwhNRXX5P+pVoEcF9zQW3Iwe4dWi9nOa
Vmp4lKUe4u+1CTj9fJLui6cfcX+ih6OBrofUSjW0SxXtfuJjrcPUXmR0Wexp/yKf
oVRN59IsvUiTVE5sVcreaJmKz+tjdCGdOLzFE6zdeT1SxZyIPvj16P1Dcdwn5rZq
ZPlGIUIhFltQcNarhDk0TNjUBVomEJ/nq3yUtsdgrYdrjRm2RnXkRd1Plr4db9fI
GRPIAJwASL2lA3gv55ajSLjv5RMfUNCXl331llV82q8BVyP/1xWX7NR9bKb7LmLY
gljSm2JV9RFh3oN/WEeVawZA3pDzdl6GVPZY8PeAGHMa7pKKMGxuI1Y1PMQh71XK
PjDxKa4HZwnFvff7caUspqc9r0/bEFjMJ8edsjL+rY4sywhnrDssfA5iasMjgumg
cHMCtLiGcTmSmWFw1rsO1HTIGD3JBlwFFm8DPdk3FazXavvLt2gZN63icSnAYuQG
+CcWybJv4yAM0ybmNaISWJseAd2XucVMhd/KINUdX/RMkx7bsunSufX9j8/aM85T
fZdE3eal0BAuKXVhRWowL3oK4X6DrsvKTtjr5RGf+Zw2Tjf0IWg9h0MM+v1kWBby
rcC5507KBgEDX/3EPMlOwcFMiY89au2BSCMmxdRkLGeBgwZaxVnJS8Vk+mahaNDP
QLUsbkS0dlavBZRYhVzrA9gRany6t6pOUBHXq8HghAYQwktrr7jDUfi0nlE1DU2A
jGOaTgi00Bhmm9GXmiYPn9Ikaj5yMSxv3exjiYFVd+UR0LMKtZbAyUj31YC7rMk+
Js5N3Ph5GKqFVwmI2oHEiBnqdyduj0v0XpKW7ZZeVCq6MCLWgvlDjs8rlkP9wGt1
O1cUeYKwO3jIRSiaStdKzwMJb7GUMFNsHaPCjaI7b6eiHeKKGLwoUkAU1HwpOwmP
UdndlRyv2e9Up5VmovGxEfKQl7rIs3q+SiaJ/30EVCanA6u3Fy6pRjPpjknunKAX
2pu+vWJi4Kp8bQlGAHCu+Pw+U+xv8phZd9SOCQY88tirkVcOXDSxAhCqNzvzl1D9
NyRPBJLJFGx87QuR3cwfuvtQefp85otFVyFrGTD+UK7TkFzmHBAfgEhJuWdOO0QL
bYYrazmATrBBkR/oQTO96BP6YGC85jC3V4alTfg4YJrJAJG+HbyiYqSL3TQ/VtJ+
MoBiaMm44CtdTqXMguca6pSckBmvCc5GwBJc+y6we0yn7GsnE86ll5abINTAPAsc
BkCu++OplhXvWVCO/3SdscVKzqCpmlIrcPWv3xdns4meZaLPs9R6Kv8TINCwzdvO
cLsCKLkEHxUsvjpNCCxC+WecYzRELHgDyeN0IJUDJ9H/hJmPF9pwiseu+O2nSMvP
spoqYxOUbnk9LqEM+azjKoa7ccrDItoLFMn500YCRbuQxrlWHFxNu3ASu759qkma
HpqF+XfNPZvNzd41b/ygOY78bfias22JZQnZA6cJUecc5ijDMzFQDEPk08bP2h6J
2wgQ4QPSaSfbX2BUQaUJhGjQ8VHzReq/UsqGb8dztkDCrJ10mc3H5v8tMO7VCc66
BijaO+NAgit0FZ52WJL55NDXgt/9t2/x5cSl1or0zenjg1SP2AoIFKhH+iPuyy8g
MHAYPoF7GaX4hA0C/QdpnwcXqE0T4G+nq5oX9e/DwSiOpC3TmqGLQ2NDYpUw1rcj
4JkUysbsTPkbVbrWoihoIO4scE0a0swkO+oB4viBQc4Y70NfjLfwkgCs8/AsAHXY
mRuHPwkFaxP7N8XD6SyU6otTUy1ffXfSuoyMGFCeJ1uYixJcTPgcLQldazDDfbQL
QGCsCbw7f2rfD8U770Z4D7vr3qzx2XeCrSDpYpO8UxfUqNQwTvD4qxzeg2np9/C9
QgdEE0VZAJKu6ebadiWjyE4dRWQr9E/C85YMRRNPxRmYesmEd61zjgWFk8qD6jTt
zkGC0TyV/Ar3i0UV8BgYtCxtTbwtGH6KgZ7mpxrHUaP3WHaF21+Kh1zaUnoBxC1U
cztx9D4abkFVCe5QAUUFdExhQTTBq/QaSJOUksi1FR1KX0IQPOXIrdyaMmTnqMtp
ucSQrLBIjHgVFthFNc9ix7FAwoP9zO9j5XBO6IQ3huGQ1U2HL1t2sie19NeEtVXN
kh6wGT9Bg6A4Myc79cCyaoUrQm0xx7mAsk+k/SkykmoFPrcfFkzvJUDL6BWz+38V
BmJ37IxcsMtcVkMSC2SMx+pxtBZ18hU0JHio75uiG4fmPZlmvERkiAug0OBUQ+gp
qKWWpIObCzhpy46KBZBY4kLmBXod1S4rtkjiqp5I5igN+YbBPaXFiO1Y93M2YIpP
R/tXhF3dtRG+cUCDcuXr6gjhdBkR2Ruly86SsWpxhq3UagNjToQSQnef1Vm4cRyp
zmkOpySRs9y236SiNQg8PPQvWCpBksVmRfKjr1eLwKDfu1uMR7cu8u1KxbELmW6I
mngyyJpo1BX2LkxAJQ3q8xQYZjFlExiHfCJTcbMqUPIbsHHjddk9v/qLUOp76N4M
SqXyptg1qVXojbBlYexwKYiz9+NuEbxav8iQy8jp/RUsA/JKD/MWkNd722fS29Pz
Gd6+OHhKseclTReUwkD+KiELvIGMQQr6rDEDexXkxu5gmbO7GQF3yd9r/zYhBgSb
3oDCSmtDD+xWCnpsGOdcGPqt6Hsoi160tVY9+gYaXMRKjV0l3OIekclY5hmRGPQi
H7NZnpnYtCqU9yDrcRs8dVDmlIDyNxuPsVk2fchKredMAKp7bAliohjT8X98RMiw
tZ7xeEETIdYsfxakew4AsbE7bs5t2WpgEFe0kVO2BlY9H9ESsrpQayMe8EVv1Ppi
dcVszYvpVaq1uW1NMdbb7H2UIZ6iRkqlzkcFpt/pPyX/jTS96mHC0e1Peq0N3kYd
hpAEV4YQvPR8bLzDFc1RfeuVgETwlOeOFqMXgKmA/iCKR6PNtQvVIWdzZfcxrbvY
PVhq1Bd4MDmIblAuoXFJHhqcy9qGpw5kjHC3u2J2bJrR+wmPhwzoWn2pGQblQrYy
Vc20x+03UJ38WJtuE24zkPGKusnik3sNLpyOmUgNGoIDbn+K78xb4t48HOYd0ZyE
QH3c1J8RCbpd6D20Rm5REQjRnfnhSFWHaHiiWQmgFsaRUWCzIz2mW5WV+iasowIv
nF11NKTlMgpcHhz86otJGyySU7yfGAKG0cAMhaVtNp6ACsp+dzhcex32Ah2gjqrx
iFHJjMQ6BFR36L9vA1Ui8tTJUsju6LRUcdaxpPzmoGJEWNTF8wL45tJxWcztdQdP
jRELReV8Rij67ac50a9lvQ23WmaRR2lhFkFHeWAG8CA8sk8OWLVcRWyXMG68MKE3
nJs7ESjS2ys5X5MNh97TARUILZjeJEKQZsqPnaJWjumEYMu2LUgpJ8nc/Sl54i9D
FAY57XkTkBUOaInFg2K0XNVf2FbhCX/jN0Y0zT9Dx/ENZaksL2IqepYuB2m/Mua2
omaIy6RMGrC5ivO9Vkhy80jmna6GkAje+WUfp1x0RFotISTNoosZOgrJb+MTIr3w
b45H0Aqul65pOrzU4tRsF6nz2W5M0oAN/xlMbh4uYyNnfKkI/xxV/iVUUwE5Ts6g
oCV81+EsY36uQCcArVW67FHhaRcEjzggW0cAg0xyF3qY/qVgvmCLNwsujjcul/Sj
/moMyHNNgRi9jCFhFE4mOLEEsLNwUIceNLqMfuNeWyg4+EmlqU8CjTH5GP1/9nof
u4tAjLpKw7VyG8ArUR6i5MovaSyduPxIPhH5S4xEnfkIgN72z236+8N7kNpkgo2m
YfL1zduJLqUj6qpfTUqI8e8LFYgMWkdkh5wrGz5HfmC2j5Xl9XRB5N+lNiF8jVD5
8a1yZ1WHQ79otK1XzVJRf4zb1f2oBzTM7KB8lqHx9IY7BNZ7DrxEYp1ybyDW6SyA
p0r996y+0WmvDb5h4gD8F2bhy9u7kwxJSHdn8ThH42G1evHmBQNkJizwZPzvrlxU
0xPhzOT63XuDSmK5oqJ0g+pw2VwhHTM3q056bNjp9W0myAjczbpHbijAzKiUPyCb
fEntpRY2qALYC9/UROTnS0wFDTlRgeiOTScRqc6J6eR6J3k5k5mEExSizJ06uuGb
XHwcwfsv/cGIaPZUH6FsKcSbtivta27bqr2QGxIsnlI2C//V3ysjCHiy/vvvffiV
ngguh4bbOi26HTqpoOUMfqG8I1UEmUmeXxS3vdXpFa7HwvASJilrLJmIDKVMIiEu
RMJ3bMp094TFNrYJ5w78w6pCHB0FjVX6wJ6aS+d5JVMASiOhKDvbz7PezkYTZ4bT
3SGQCOjM1+T3xCDb3CA3fXb+22dCvBHC6EhV3Dl8hGW5xD2AakaEgr3JdNgmGSGS
Rh9PTKSK5RAr5QzHQDZbmG/R1Ykc6kuNJhhA7IbxrmufQCh9WBtwh14uPOHamHtP
aXXgQcyzu9dSjT3QuxQGRYOvg54hdIuh8QqkUgnMBrald5ivaA4mss/xfPEBKhiv
hQ+EPxMj/9UpClG0twGV7n+8gXPREmOrwR0UpXQmtoJJqlbcojbRJ3dyWEikqxIN
Yhi2bcj/sDnRduZpiZfrwZ6ELdglPVZ/9x4CkGDSWlUCf4J2ILN+QX90HL7SF6J4
aaMkGougtoe6DjNmEI5IjLZxMcTMSze7BWpJzfHNOQuwnyJ1NfRPWVLiDPRtCgYo
8HJcU8GJd5tEgJwXRM6Cr6wkH+WpttYb2AZycC5ExavXR8DA56YB0pIyvrdbcgqq
nHH5QI5KZn05/vyKfgdmR63kRzlwCqILkAxHm5tBFrAcLYbtDjLzOltEmmgvy5Yv
8mI55JWH/Dr5GqaYXlj/SfleA2ti9yRAOTcYI10K9ng5f21cDLwyr2tKqOvefThI
mcM3fH8HxEf4k0xMaSzc8H9sQs4uEGsWnfjaSctcJ7aonShltzluanq0e3QOcxmL
VkisqCM5PDHX4Es6eJ1FI9Tm/KQjO3fysiM8ZyQilvShEC+xANN0FkouWhY27x+V
8VLhHBJICpM77GAGy4B+ZMy4DIGGI8wLhDPhBDmFe70DBcPU2C9G+h4+7r2OndzR
3AKoBQJQiOlwPah+lFBFoPKzg1jLXh5wUJaCkFG2cvha3vjkmMXmZqJKheYi6NEJ
rDEFfPsOuOsqzVktber+iSRpaSvS3IHlSzmus4EcY8QO6rav5zGc+K7zAu4HQ4mm
TNO9ATyEljiPGbTMh4oFhz4VnFpwkMQQ3uN76wl/irQk7Rq83GHejpmYzVzt+9p6
SEcMvhjiCrdx7us/QPXttDwKnxeP1zF0W6w9JZy+fYXXMqdOH6ldhW7fp/zX8/lx
Tu597zUojcjTsbUDvzZCP+IemuC6CAYkgL5mpVVzFtMUDbAsJpZP9brRZ7Tjpz0N
ZN7Sq3gTMDG2XjdfjAkIIbUGJWivfU4KY5Y89oKxd8QjDPFMegFjotY+kiSuRbWj
3b0XGy097phPOE2k29NKOF39yaPf5Jp5P0YJQpnM/HuwBHiWB3jAk0B8tE4Tdsn8
60LKIMl01VOC9EUqHshcwSN5Z1v0k8bkEhYZdPXc/Prr8o9XvUStA4k/DENBKR38
l82sw/NG4fcAFHr8G9JM01XLzt50yhL2w0jvqiyq5YepBgb1TIKoLp5+KKy5Rrgf
JcKEJvt9ZTK4QWo0xK+yLCngi2qQLidu3VfGyxxblLugwWuAmvlClncmUUIQcqM6
NRoTCzszcJ6aClZSafw67HtAy8Y/Gnp2OCJL1gKfTy3AdCK3Gxd9ntSRtiEV+FYH
SDHsGJAnUiUorFWXMwFz7LRAdq+3GWE5qTPY5Jg31NTxBuy7VJVqePC5LmH54Jt8
MQ5FpZxhwyNp8e6U6X5D+z3ewMaN/FryOfxLxTRu89pN1E0MDFrFVS+34eKbjinJ
gKni8UfHEmuOW94LmX/AB/RgAD+x/IS/gT7ZlZE1waM1yC3ikWSNCkcnJFoFAZAj
bdJ3+BXUSeehpFdNNrplOgTzyHZCTF/FFDj8orQSQb/DH9ViaTogV0mDhPOfFIbM
tvFfOQauITZ0l4depEyj/LteRvbZsxJZRX+1H0R/Kze96WwwuJzU2gFIngeERqBQ
D+gs8nYi7uQ+73ZvNLd2o3Zai4ixeC8uVoOpo55nGQNxu5Mr7zgtzzvGF2itAR5Y
MLmej3Pu/wsdZD2pnWo8UWc9Lg9tA4/ttHYZoLg+6XFDeHttdStUX5my/yHOPBhf
CEseMzJ3VCNKlz4I2NFKzl4ML6kDh8EzrGfzRa2mYySz40u/xgrmfhTh52bEfOfv
k/7FnsfZi//jo/+f/kjzAuvhUky5cge3/hPmCMl1CVWZPqM62Omt72B3r7caNnaa
bPExdBNcjRNEGhwTCEnW7qjoybPC2hd+nGA7MaPRTAaDw/NkHztiiiDKnLuv65fn
lHg4gvb7hOB5I4/fxhdc97oJrWolKr0cOlD0MIQFuaFrhQQvxFhWzIaSVxaWUkkO
jazHnBpuMuGzOx/xqo1jFANKUMeQYs67lNMB5ZaX+kf3s7Xe7HIcnwcl2kWlN4Jn
BKLGrmaXekROQY6s42K1ZA80IYDPDfEkwh0Dqa1gLMUhdMTAuJQamSg/xAWyjLqB
LIXwXLyw2ftOQXHkgq9iMVepsg53y0VeMrTcYAhNFbZx3EoeZ6ssPr3chQS3cqPs
7eMfRwPTasgmLrv9J78Xnj8w+TkfMI+7400dG5hQq90A1HBRe+7EgihK1O+Kvy/p
Cw8AIQUQ0qmONKW9nAnEbnRYTKHfmIFD+DgdR11Mbq2cJ2qvHTqZI3m0X3TjG367
WtWzlLgRYPIOJ8b1Pv8l3hR3077BUYwFpCMAhWD+QgMnBMX0J2DGcu/ajelza8jz
Qimm062XlheNQrsKTjARYYHYsWJUX4sqcEQ7L9ImZMVff0oAD3fJIYsXItX2KJII
Hq125pNtBt+T7gVFtHCCVW3GyA1SfiGX+N/SJVmpQFLoAlt5c9A7dsUaGM7mmqta
tOylQX3NUuaBJ9ZF8tZCGedPJcgLweV2q/N7QRooFlg90uABFDQ5q4edPD7bwy1H
ozPMKOUg53vge1xSRDWUEFkxGTaojcl7iGi6ykT2kENK1wxk/LtFcOtJ3o/67gs2
2eC5HJMk1Ns0HPhkC6Q2DViHkumUqyOSmY7n2CywS66ispTklzdm1lAtYnwZYzXI
r3pIzZwP+vBgZu+6XQXE4aIf+8wztnnoVrcalZPcQciJofBe7Ejd2HeVyH/TUGd7
2X6PsXuulPM7P6b5Z0INzGERp+ecTKk6qlTovEoKUMqVNinp8BVAaeM+pjBm6wvc
9MbeBLRZ9dZH6JP8aISJ7Q1Us0Yc0VFnWtvIDVrvOS2Yszzat0DdegcjSl8jPJvz
0fuewbg9cgvZYGIhnVKF4zGaTsAU8/znxFzqFO8uTafkLcQHtTb1brIwxa9RmKAY
quKVxZcJtA6RN0jncr9AB9WZRg3hjpCiIEgVf+HGFNGh597/wVQ2LF2X9/XSiKw+
7x+01c6fqaObSP4vQySVkhv3byBrrKObHaOlaMkeL4GtFzB4vlUwvOWeVcYhyBrD
iUK2w0ELL91zW60BG6bFyNO0xIT3VQgqgizrfSvRJCBszS5QAhONzqa1cAjoTzLe
UwKGJyjtxAKZu17eDf2tE1GsfCNJh47ZuLwjYv4OB3LXVis8Qca3ngNFqKfPecBS
AtRjFvYFkGDeKf3xkKCSbSiN32gbl6q/ULS2QikJRN/nlE36o+kvOnaRUdjym06n
jmAROb7OGYFEMBN8pYbWc8rd4Nzh7OsvDhLdiwAPV3sYmvPskxCblt8oxnpY0c7d
VqtApsrp2n5n9jsZcDNWYOohroDOxlbzcntgTYBYeUD42nUNbx2WEXNrrLsPs/Xo
jvB1Q8qnnTdVBGWHMgGOwJt+MEsyu1IDKy4tav9R9ZvE+Ir2ijnnm62LBzT9pPQT
qsc0H07WUyLCeXOvNHn/HnBX95rzcG+wXyk5Ofx0z6EvjEaoSuXbRuODr2cnO2Yp
krkqgfXtJYAVv1bEPhZsVHItys/mSRozsrZbGe85r7gSB7uXc/Yf8USiT5gJy0jx
zUmhzW8x/wtZg8v4gjlbP+5isz81S+W40I/J3xbky6ugeMDPAX6IqN/Juj7ctG9D
BKti3Y0QoyfqfaOKJZ79CmgNofMxtEBum8vgPF7PU9xca8rrWpoA8jBsWiDXlWVZ
yAz37O3F0Qgz4ClpISQ5UhnKS1ofI5Jl16CxOVKvZ7YEAGQuCmlPWNpyUzyQkH9M
ZlA1Kz8PS7MJJSUfA91S7bevZZCBFd5xbCCQcMZTHJZR7DSn4xB6qkrGMGRkjdSV
lAtnoObDKas5IxVnVnaeexFjn/e/s7p51+ynP+owF49Ft468oY2d/sKjY/cwuvZP
FBwhANF5JTOdkgOqUem6oBZ85e1FUIB/TTsuDcidC5SI3I6wsRZNWIWVtvR/7KIv
PGT7Ng2HLdmP/VrEPLttnMOUmliMlBHrSkTO1Y2yW2waz0Dl1ytlHK2tUI/auDWJ
BHUEUQpL0D1D0mpY5gEKhU/JUWCZ0sfSmVUBWySZGZ1plDUf8zoa/ZgbZdSrEHni
NJ/tEJEMMfI+aoy1GLq0Ad0BWc7sjyGn3ByGhDkOKzDyyUmIY3hNLXJAU0sUFxLX
clPW3iCuGt0Sh7CZSGQ69eVg0uALrtdmeQ+ClD9Oqt0+QPSzL/Uw3Cr76NapU6zg
8vptH34AwhGwXl3M/gH9+u7pzTHbRdi3Z2Cg7a4oPvqOPGfb1Mumtw49t/RaLt/T
2k7dPVms0E5wxauHAcWrzauWtz5t0cTik3RW3UpyTd9OZp8oSSjKLD0tSdDo159l
eConDoaw/n9jsmlRV2Lg3jsllvM7RSUEHbJxA3fCQUIYOo2iQTd63EyNCjSEUMLG
dt4femIt0bAdwDe2XvSj8jKIVRAWNmkBE6NSv64qINqctBe/o66MKgySxS6+L6og
91LKTt28H2zFg/Zh4Rn94dlU58DMtI8ZYNCitGCQ0xRBw7EWhh4q2llfYirm4vXd
j5nb4HFE+/caXUqaX55dOHF/eRv/nN+/ae11kPgD9RoJrbSm93Qir8YU+b5ZyiZ+
4FWCNlNy2jjO7V8pccCh9irof1MctW8zR6Wzx4grSn9gyo4/rFcb/l6Ab7ANSkUF
WEnRHi8l7Z/RAbD+ouCQRlafdQ8LctqD0ocofI9njMx1mU8eyLZrJvEq2X1UYGNU
+qNQlefi3aOid9rJ1+NFI/jtOe1AK0jx8tcaFPuWYkru0ahEGaT69VHuAVdYGuoQ
F8ePoy+HdlFBGM8UipO6gh/c6sReY1nThi0JTQLDhS/Wlym2S/ivjO/rRcZ9xoDP
zZoBuHYUG0F3U96fTJPvpEZrcXEwUcNNFxgyTjF1tTKt6HLNizt76VWNODOSFrqv
wqps+LpiHu2k1oY8gep3mWyzuCZ1a2p2xw03L8KWxHKrJg6h1Z0CBOIrfxqYf6z5
7OeJepsyu6lJbE9kTrEI56nHf+g7O7FSu7znIBORD98cctfpE51TRepfUssIXetI
TZ7sbQk6iSsZHasnwElKCZehoA9Yt6u3j6sJfcRKyWcW0PBAK0ZvHZlrpth1i0CF
sY94nXDiepGh+iLOdz2r5ZEpXtxmF3TNJkqykUNSBgLt17tE4PRQJ69hBa/254hf
nq0fvRc7TEJEojzVH8gb/VzQF5mY70Y2K950V8oqgrMr0/lmiXJ+TAiEEV/QzLoO
dNUlh7pOQsodZxAsSukY5kj8VFyhE9+a1seV7zL2I0jfAd19C1jiMp58nBRJb6tD
IVU9zycT5U1ey58Ies3kXxnQfktre/8eR44vK3Mg7CPx4agtzlMhx/0gTf4NzznV
yhatC7ajMd+3hZg1AqF7/mRlgOmzN9I8wyqN1W5/ytXTwCEeKsvq096BigUWQw+n
nuLt9gFmRclge9GkMqxCo1GJAM//hNOyHY7Je2hopPt4BIvcQKzJyq0n/VjOyFAw
DG4TS4Z97561B0GlfUKzZJaMDZwfalcCnbaAfzb4U12wffFMSLGRo6eql/BihiWZ
svMPKWdcK8MWSjt0yXI4QH1Jibmt2gbKADOC1Iw0+MX966JES/cnMgY7DkopW9lC
cY/iwgrS9wppRo9NbYtaepxgCekdnXrqLtc1wJ5Wd/uElO111fy2EbOVbkBONK9n
zfvPB7akP3U5yttIHcO6tLwvI3OOIi0V9WIUV4nS1d4gI1MrDZZe2svoKae5o/rk
/pHGlvo8fUXiY0rRBpHO+nrvjHIDB6v4TX4OHMs3CB3sJZB56Oao5ifQv0mV1QxT
iHnVYo9+eCsjqYqSPK75EyjwSSK1spLppdWxLkRsUEgq3HXtveDHjp0/eVFq3tV2
RulDqsywo+Eez388HBcdCLVjiGj7PyDMCUBWJJBBD9Em9VYnpBh59j1iASMqj4BC
Zc2K+6gsc6uACA2EKMYI/r7z6jAfk7xVPPNeSMisodrkLsF0j4xsg3+b2JTb2WnI
loGBL2OUHmtrnj1sKSVMDyOYXP632HKBXTNQGLHcyFcImq7hNeJtro+EqiAAqxpm
U3usNWB5fXHIPyySWljkDKp8DfrlODH06SFnaUw+o3AgpuhuqMgM2PSaj4UVhop0
XcB8zyz9Iw1ILnwTMn4toHNRsOZSm/t1/piLO7esvw3x8gaFXhgUPBYRHWGSBt47
lVrH6MgH9rgiNlNkMtoJ6XoUaVIVEfdW/RbsgZl9mVeRwjFEu/KVcGYcAAp4xTsl
iK/4J+KeE1A6gHOwJF6ZCUXowZ4oMfLQlc7ccE2ru4TEB3lyxnvBSbGsyiy19/nI
zo/rR9IwxDv3IVQsKIr30Aq7QZyHKBXPROWp7291scE4Oan+eGxCR0t2tg+UZj8J
svybyPtkxU1cCovwRLnfvHGLUdXGbshof4lHn9DIPLxsU86v6OZ0f5+6J402R/yL
/94Nc4IdKXkRoOZlS9zpgwZN2FAHD/gj58QzaMzqQH9etwKEOYmBGQvGQjl/QL+3
ONS7iAaLQVJHGt1EbK9xRG0n2Sia3AndeCo8XN8MApjwmfQnIIHJkExKDNcIuOmK
S5zI7myiOCC5vDkt9hEkC4Ab0pNsvrxY4Zc9XgSn3qTh5iLrIBfInhEtoiafRaJQ
3fApD2+i3rYb5P3Q+v2mRXt9uulZNUDgzZMQ+jKeg3+t4vlnD08AH9JPPif/au2x
zjPtDyRlV80b43f/D7Iq758+OV1KSMx+G7ThdJxiD5QzYVMa7oF16fIpaJtyDXJv
SvsdJF8lEuV233F1oXmDJd/DbxlKB243JmjtbbkSzjiEJ8Umo86n46BS/yQNMQiv
YUq772QCFZHvh2N6LQFNUL0vESg285nsbMOPGaAcWgFoBlgJ3K/p85DZuGwTL58V
FMItAmSw624bxv8M4DoRG8DjkxQoycrNwIf5VjmmTRfVyq/lLhLlmEiyykBXcvjN
F0VuGNtOFYl5FfijSeruFfh8jWK8uTKT7xa/ifRnvQKhnR0dkPJpU6qW3zdvpquf
pIRT7BiBZOe1u5oqrTREbP91xiRgbJOR6U/xn5BDjHGoqtpmxyWMuMxfgqW3Rwtd
g8/qws7P8TDgQPC757pX4EFx0sOenAT1anzekMQtBvvOthMwpwdGuOjWCiuuPJ+P
By9Gzn07Sv/f4GRsGFmVw9YSOBicGsHans/Z3/tQC3qiaDtFj7Rypuuxi8iPXap2
ZEHsjbZ82E1eg9LRLH+qNmK9csTwI06srnXbUNeCmFNLcT0DL7j1HzGAJOuKvx9t
bRUONy2hd7gLJV4du3LrfcRJ4ZSFbTxfLdPEo2Ecls0wR2kNpOXUnsLkGefuVB8z
cmuj0ZmNjZeb6m/ZCvjKiKMQMExNavMNNp3x8jsw1UDTdSY5DOje/1O3yM90PLMV
IUEN4mTdlw/9AtlzeYcUtn7/SUCrNUl8yzr5v/6LzLhXqfU9GqrynQaA2OsokjQB
ps5jbjpEJeX2jUvGJhRE2hGzNbL3/1BUejOMbrwnxLHMCjODdooxlyF+oNrSSAnF
nsEjxvKDm7Lg0sGyUWMkCC4Kw6o8zTdNnsCpNhR/Kh+3ASnBkyKJeDe8RTnLO7JZ
T+YSIcGvSP8rIztxIevHkrFW7ZamJV02O9ygytWyAYaXQN6N70+pcGTntmpSCZq1
1M5TY1BrQwGe4uGS62g3OaGKXLnsGzltxRpikxpH6pbAND4nSWz+3u0x0mcets88
4iAvreM/8GRj24L5nSf5A1pdaHYHTgzZzfOwzaWuelLm77gednr67ItAoxiM0BwF
N46ybMNnslYBGXT6gB/tjxbXBhpqfBEVvIccenwmDldyiBpSX6oKb5Rox9gP5W4+
fwXAAtciwAmz9cjzSGnTJV6WSRn6z17MWm4estYz1JyMJvtabcEwf/7wFdE1pkRZ
Pw5M7L7RcVOIs7yrX7w2HiTzhhTBzql9IhYRtUj9+7fazgo4emxGpQ1m4YTu9EhV
KUeMQJ1De6FTptp32FadEWg3xJWwcAGBm+z7ggD3AelaU5c3Asi64VQiadHoKhfl
8wG+RxL7Kc+9EkvzzjP6PiSrDN5/bvbksResnzaNsfZlzPbv8t8ObqtJrygBkxyy
tWwQf+mVZDIScos777pIQgoOAbs1sKsPKT/Pcgg9fU3DwE9PObVqUSgzAv52gMeX
FDnf9oBV1EGU1YK6JMsiSvEpYskI+k55DGm8dkSdXvOk4wfwtgcD+w1tls5sRT//
/QCGEICsAJaXTjm/4kfgbKf6xoNkgkaetCkkwrKmaKVB41Om4Vpmj6eMoHsgxEko
xNig2y/h73K0jQlXhFS9grepxHQ/Prkrg/Kj9779LNhK/iIVYPPj1bw3breNqN0Q
ODs1HXOzPMsqcUBm1PLifbRZt/E9MUTLniVr+bjpQrQKZ9BhhSvUl+ngFc2QAmMc
PcAnqHYOKji9MuKaLnA5KYBjNp2gvi1FG5w7/EkTqiaTS4RKt/woF+nX7AmHcoAB
yosmCNPlm0DDq7I81ogrdF4t1f5OVFHlNm32h/AGZyK00/DkYuhHFbl97x98Fi1f
6JCLifHjpRI0UCIZkzAJ3ytCgdjhUHrVUbaXWgRgq6KtIpgIksvD2LC5QLeIG8Qh
A5OHjfasNHZ89N6IhikvkOQgPw3+lt2C9hH6jehPbs+05vtez5WGqQ+PQdYIt+Z1
rf82Jl2PfNUFQqhfjpVJxvJ2V7NaDkVOvLamoJjTa9nenEcFQDUBhSyQjPB79ncS
+w41GKplOhb77zi9eo7SuuxtX4q+pHM/Ch7wDfXdq1nGwmd9T6MpRXDGRt6yhXV8
2PUTbjq41YR2ZgF71rFXcUwlRFZO9aH0V2YSFp5DNNPwc7U/vkpOix3DpihJx5sJ
igzf65l86Tlhjg1hFt6qGS9wHyd2cbuEe1G1KtkWMg71qQBqDrHF56LmiMF11RlH
rmMLg3NAQsPxhtLG5LMSeO6uk4jPZ212OWpuZRKg0+S1ZSiKz9RTxuksUiXQkdjv
+HM69B4kWshsMD1snJxfDuxzizU1LfZJ97cUFnPSOf1rZA0hE6EXeHbyv7gd/M+8
no2htGRXwQvoftMg8gxRvvC/dYgzGBzUMvTRSGUT4stpSIvPes6vdOXdTz0V9ve8
E403KHqlYEsIunLftrI9iqhCnaq78zjTaqbQV2hGMo1S9srtTY96TSvIj/p99hbe
fnsVZYKbMor2bOJeTA0X2d4AjTEJwoEkRhbQ0W6yEXmPvJW+S6q3DQPagZxU/HxA
0E4JHLHWof2TROrCDM/onPNgQeb4/3Qo+zVf8uWKWvuE+pBusleBMD7ZtDphSYFz
BdwvnY6vYQWSLpGFmpiAz9T4HUFdrj8+Dsf06TQKoiC3j9hBgYVQYtcnQ5Eg94Lc
/NeVUZSThCx3pCCUlFFZGx3zjZbzEGlQg0EQyOx1ZBZyvpMiYhwbOIrL39Ktr7nX
doWujoy/C1s4ZJrADkvfAQ49WmlggafvTUgekUl3iOySqyJvtxknMzsMsEflsgN4
5DWvqFSKNuh/kwZmQq6MuZYzmEl3r/aubZwNfT1b4QD5qf3YA2JLK/Lbbtqymu5A
CLOdKzgbwtjNCo7PTtraLKWc4ZYsCbW4cTSedf/W+Org7GY3AvLcEtZ5oXY/ZDl8
aGEb5azcnJamhRZeItSC0asO5/5ZNL2hmz8yHz34obnKYhZ/ceu417QkzwRQycId
RNnRNKIZQHFoGDWau1S8E/0+Y0hN/C3nAEbJK0y53W32TWB/U2G5omv9vSieHf4Q
6aZnRCuJOw474fGQWj3mhfV3UggCTJZqrI+kuZ++ZDJjTeS6j3zFUM2IpRmC95BX
oPaeQEiuq0f7TQ5+QpJLzBZv9lMCtqZqCFd53zJKEzYVLr+v+fzZzCR6NF4Ko3Dv
gpzyaU9gJK0N5N7OGI05BjvZtzfox+GIjepdDO3Ja0p5m2WUXsRkm36lAD1rcgq2
P3jhueXTiAUtm47RE8+Iv1/VTXaMv7b2lgWmHHq0LPGKop05usVI2OihqhQ/cAwt
K6v+UGzSUR5+0njSge607hFDRiRAY+EJEPiYe/gwOJKs5lu0omW9wt2iw/eKHnEB
HAvutiMzA44ey2YxcL7eZlykdheSoFP/oqYCHW7mDuZ4GBWdoctohN2WeG2HFFRv
GPYzq03TFEXrIfyXGgk8vrlyjrrxK6AjPvyh6sNEi6iTmYgk/O52j8kqTlOCjVWP
U+8IfsrVKno+wn6ObEfZpI2vcz07pnJNAw9qof6ndIqeB7uRcUPRrOGLmrGkRQy5
sXBOH3v7pG7UgnBanf4MRjOWxZvNkYlwaeGBA3hj71lkS2TRewIuNRVfZr/343MI
xOf6IQ1ZuLwIsci3dfq+Bs+7JA6Qq0M3Qkf79F0+PrABKyzPAtICsQOGQo21bd6s
tW1u17hoe3dGUX9hBuOMs+1gPUhPfT87HBxxcSWpDUjoeNQeXWxgH89u8vpv18di
tbjFKE8BPGBL38eOoyGYM/jxaz2q5zWTieaZrzvOBq1ZeR+Y1tc8yRQQey1ULubt
cTfVL4iZvnGYr0U3LmUSVklqU8LshgnZa0PzPmYE09Vy4f4I9qDip/31FRkWE3JH
KTCUz22GJMQtSmQCybIUxSGrWsaUgmC5lO3KXRINycmGqg30f67xFvfnBMUu5cKt
fJVW5tQw4VDbSrTvTkkrx8FV9rsvqAtMIaaD5bUh/BlghB7GskytLkXpmFz5Hshb
BG8lDQpzK0KVxtU2jwvk4ihCzZnNyWPWzzkfXNRKzm2pBzyMzzgq7CBkb79O6tvm
z1TgTYyL7UKFB7meWx0rnSO2nkcB2DmpNmTla3csCC28+Zsbg7u37Luh6iPO4HxR
w2DlrU4zA91sHWl/PK1W/7Nv8w6a8VRq50eOe4p4hDSGAvTUQfUB0rRgBSGS15hU
3FDbDG2PyppiEsNbqz9xN4QE2vfLBBn1spx5WuVrAymfRp80McaeLxjUbQbaRE4u
EIccVeL0AjQChv7KyRrRpLcGiwq9fhUnLqQFO2bWfh/2NYODzoN6lM1NMkoeaRmm
SzAWQai3WqYcWec9fgIyhJSjCCOHHsSvQYA8uwhroghnUl5iioWPQvUlUBMUxyCc
Azgzn49Eg1u1cA+0+Zyg80y2IDIE3MfG1CyR5Pu2DiE04ejTRCt8Lroh3jD2SKdG
q+ZSUCwQPfhSOVSk4UC0mrXfQP19zn68o8vaY/zpPdgYb24gvtopNC3l/rC8IRTu
pr/Oee9a/fJKS1U3WlRco3jSEapmyTm7Y1gjdEQ81l9jKgzFuyw0LcHDRhGIo/jL
E7NGc4JUWLcI3Wh8scaqfy/m/XlKgf38UpFHpIMmvFNqubGileHluHRgenE7HZUR
WNeCeCdBwuXq4rJ+p8pq0vWocz38E4ckGx7J4X053ec9wh2jUeg9eU3yW7NOdPt+
4d7M9tfVc5vmLLYHwekYDtpzlm1b2t+vBOcGhVgajBkR1cW4d+8bxRP0N7K+do0i
3Hk+wzOebFxX6EkhHINkuWmaAZlkAxvXOfG3t8q2cqs26F2B35KIHg2sOu1senS6
YqCbYlvYvHbfyA/spNkKRDF30R7C7CoyxCxj1pc0HKLXx1ZxKKSdfEQllLKmXp65
aQCOL8aOjL/tRZLcm6SpR9j4jEGmKHsxyNveIq96IE7GKWrmbIlz44nXIN5mkGLu
0r96BFqMpDjGodiGaidcoday8B/rWE3+WtWlLucqmsuuGkRKxRSy8m6mzilGFxeZ
DvfnRa0NI3F0EWURr9/pFc0Xl4H4p2POlkJGrRg+8tFbQiQLlOPg3WaZufJ1/sYz
ubFTQYg8E1gbBLt2XaIWMCNptIJqqL3R60t5AlyY4FL3vA0qOt4jdeuFGZl6oixK
4TQyXA/xgFv5GX4losLp9qMJqPunYrLHHNKiCdOHE06XeRQOtXXzjIkrUqrgpAwL
Sdw8r+Q6t1tjGomdm+se28ScQjj5mPYe0RYn9YdCWjy+6jnQXqSH7kLD0+dZCkOk
NiAdrzo47xzUjPHcPcx0tJ5iOYP6d4SO4cRPxKjBaAVlY1v6lpYL6puws7s43ICT
rPAgdffdONH3eeuAgZmJT0ZbiEMehxoVwX2bcnSXElw0J18Mpo8+Ay03EABFzJNZ
f7TYWOvSZk+VKn0QL2jfncAfcJm8BFB1E9LVpK8AypdD7AUPjdTOxJdz9iGZsnnT
5go56/kNwlB076Aa0T85Arru8bxUMAX5AxYzNtFF9nGO0eQ08IuBYSmTIWFcURoP
kj8UA5KxDtEkdF9n4Rui7fUEm08LCXw0ClY66zabt9WjOSzbLB47gDMsmtKG2G2X
kaqr9HlyxXhWfa5JPASXazdUilmaJdaoJ1LDG/PFrpPpgXPlmYvv0+0jtTDoyMVG
LtrSutxwjfdX7jegsNlW2QJZpkdavT/tWYBTIYUhW1CKtYUwh/DTgkORFxqx29me
frscPCbeu+5oib+aIcq0StsdMI4ffy4yLdIo660/O3c166KUQFE8NyWRDpuxAZsZ
dNqzFlU+4ewA0e7nb0wZ/RaXn43Ws0Dj+O7/P5Osly14fJ0Z25ykiyj4AvVEaUVS
ZsQ0yy2RG7jF2OyHKZk+xubeINNxfM2rZno27+/aoQl3gk7nVW+WKIkYo8/zj4uF
P+weH1pILlFgMhsqfuNA5Fe5m33mMk/a0900atTPykKOJlYwp1U42BxLJMGJ+A1I
cUUm24WwnCCqb4OjoICEYP++Nq9QpOdcnvgpiGJLzwMvkSOhZ+dYFyK+vCF0YA27
/GjcZG7oVU1up5dAw+V/NTX2RkQ/8r2QW0fV6EEnb7p1Dnm6WbTSiNsH8qqKjjAW
dz3Ojh4tL7nc8syNK8Ddp2PIJ1WiCBIQSWCpb3PSPd58HBNA45qgKWrRoC2RpgnX
qCmMaPEZU203DE0euYq0K9yMyHBMEdO4Vbswwb17gfyypcUfTTGGu094UMqRYxPV
qXcLUGldP4nCA/f9SseV8R0KEcEaDF++hj1bfXZYQH32Zi1BJ6122OAH+HujnpFv
G1qaWLgyFda7JLo8X/CoD0ef+siFxapiNime1pWHsdvDlYavbt2iLJgiBTSW6T0/
rfhFLnGEVICJCzWjKQVWPhUq2BjnMyz31YEIrAVlqaLK/D1b4QL04cmfdPV4O+3s
xjC/9Rf2wYCNjE9xE4Mjl50CCJXK9QAxSTye690i0rwvT5WW8AnyNQI68hJZQOfw
me7Ha4ImqJvria9ABcATV7NKmw8SXheBcXxplsQwJ9AF9RNAtgUmbOrRnki+dC5W
GpvSZN8b4L/g0yeyY/H0ZaVgdoaYNDtwNnChxPaw0IMoWQWBPGEqNawDQxSnzdCH
Gipe3E5HZgfXNbwnnwL/FkGQ0Hf70NjVduedWFgJzTb3YFSjg2tLn/ib+uqrrclg
aQQxjzOKkNZpwXTjS4DPzi1OdhixEFWiEvkyERAVaS/Lxa+zWcmZ/LwdlEucTFZb
WkwMQujrSa1+lsSQH3wuA0WBscFIKVk/JZVQpTa0rddKI2+LKM8inz7pSJn4rUqD
tTjayjJUzNqO6WKmDw8jIBnAOjcrfZx6K6GzHN6ZLMFDtxoPnug/wf8dz6De4CwQ
dNcEsooxOBM0RQN+ZbyQ/y+5vyLNHME8Frc/A2V5SLOzBBjxlt84dm4hOgIVfyfV
9dUlvV8dzE9GF4ErP7Jee0Sk4WCJqVONdA1oTjebFPDxAr/Nd3AnfdnZ3ASvx4sU
HK51HNwDRexVWD/XGDak+PvY8jszNPshtAg+KuhdbGLFL2o9TfX1fcG9tm+of3wo
mazX0vyRK8LJ0TU2Azq7Q7pX/cmrslkaYFvxybfMtN9+KnPN2//mhP+BVoOyF44y
NUCuqIU7UNLeVvUPXn5dtEJYckpKtuxTfP6ZEBu8+Zf71QgDJ6KjaaFiydoGYr2P
Z3kFgZXbEqafycqT28ywRWiQH2T8qBR828SCL+7jyvrPAi03LcoF8EKyeQHLytJW
Xy7WQF79vJ2BGf3gngrVllf84+uXFc0oWQW5b+cQskKUtgA27CNkxcl4Qk5+e8jO
MoASJKmzeGuMN6qwaOwZoyMuvakb9ODe+Rgev51hSYRkXxxsmFHYNqOPEHCqK9ZL
e5IYgC1sOvuNlrfC15tdSSnRRg2PI9ruarHi/9lIvSwh6SApN5xkppf08hRiViZW
kSWi9ZiM6OZsDSCoxlNWWw5hf2e79K0CQXV3rr8xivnetbHbYYXfz8Y19sK0HQOn
qCFhyY5nnjP5mNi5odV+T3YrKMBDCiq4ETb6xcwRqZitxd25ZqH3n2BYqhM+W4K5
x0YqUhd4dWnfg60iW0Y3w3yiaPXdL+1Q3T9v/Fzjqr0S1+NoaEthkAx527FwpHeM
e6UTNlTwnbJ14662W8McT0422087DPDj4t1SOTVxtgT6XCukFamoHaIMGsMdL4qw
AbdWGHkIhTi5PX+Dp4mWWxkjysqchj855Xy54PoawgU4eSY7QkcTDKapvjKYACpY
ebm87YhmeJT8OIJpK35jzndpd0FUjoks22kebQSxHhhPsr7QfvHtYjMvjPiceKsT
RPkNz0xyS51hvUL967c33u8g74FaWVXu8UKKzMiou2f+biRAzcha9Zdd/a3wRB1/
saps4ILGwWt4UC+D9Cn5hnMsOguub55D7fwIvC7eFdeATUZnlKARgrA7+ue7fJ5f
RBiJGl/7+tw83BnoxAbvyIJ8pehChtvRGcd3zwRSmw9qyFpiCxf9JJPs9rGIkz4o
HZJFZeHL1/ky4/Up+I9YtWX9e0j+rSj2qeluRFHyK7AojCJ3mNW+kqiQodfDhvsV
9q2uA07NmixcmG1rJDj6a0UtqDNuschnUiXrxGk1X9Ma09V93UTN19o8xn0OcyEh
xYSx2JIWIXZpDifZD17ck/8/0ZvPylhPJMc29YXl1+ugZQOQmUYjNx0IspmShvhB
KMC9vE64bM9UVFmJizfGMUawEv5Py3bA60+4DTGl/EYKqS6oE8bWiYpxjCoxLZXa
J6liIDPv33p2bHDXx992tGjXR6QtX8aCZrAg2yRCnudXZP1466uJrSH9IPpznbrH
YzQCROnbQ7BjRF3qeGlpNEwhBYRLfQ5SIYPi1XHuwQ06MChUyOnUFYWhXZzPSSSQ
9CCoM63hkBTHh1cKtv6ETwGNJxKlQ4i8FqT5CEnErSlhMSC3tYafSFzNsbgnKWsK
pujMms8Kpii+zjMHok3wde/p0aVmi1vQjEspBS0hG6SprzMIVnQvLULeqm7nHn3A
+K+epj1XY27do1s4fKf0f7SoAoXh+ej5R4Zyuw6y3Pi2hu1jcWo+/uIuLI2VZcoD
f/SwCArPk4lTd+rEJTB9qyVhuKt1TQ0DKGriZNtxUpUFn8+MsI8kfdXO9bgbZW4Q
+xUmOjcvK6s0T9b+E/meuxgs1oK5TGNQ4BbmaFLQfEJw7xxKfTASV93wKskyECrd
6bXR0zOn+vqnBtYNWQYjZ5KU8C9JQRwS0WoUsmX/DdO2XrPbKdPMaa2npZeKkbVT
x8dhBMr2bafxCkFXqHVwjPmQpQ+j5nLGTaRKAiACv63YyYzgHR6G5aqqhS3w2jea
npWUEC/nQeNu3rmAeZ3JP1uJP8QRPlzaU0jjp/og3l0ASp3Vm/EFQ88DSTAsKeGW
YdUcppJF/8jn+jZsKTovo7FfXhh4Nq5+SmpNh+OumRJth6JrngCgECnh0WBRofw5
TpvloDCfD4Fib8O/BjJOyFf7MkpE6KXIdvd9IczHQXyYFnDc+sNnGIlrgAT/e0LU
yZXs3WPoP6TMHLzkSH8m4xRvjkOybS/6uWXrTZF3Mb52UfJkLc9AjopIhsQ1SMVa
do56OrAwXf1Mx4c0u8oV/yDDvrmu+uW4THkIR6Jl0BlPb4YM7PAmt0cZrHs7GEro
b3BT7FZdBrNvHW5VfzwfLAXo/r885rC50EDwJIs6TYCrTsCsuWocue4P6d0majo3
JbrhW66w9QklWKCWRfdfcNXCgZRt1/jnOZJdx95fWN+bo26fxUuyI/M30QeYIMwK
PDuvDqZI4THTrBG3+2pasSYkF9VH2tfst2UjXWqgHRNTl3bxgzKJHyLa9NWeTqjW
YkkOmwCO8qqsBurr+THZHL/zWPewrlwuKytUe1EtqLKDZzpD2w/jL8H00CbC/j7O
TLvHx9hFwy4riOMZuOjWyYs7ZJ+ORXFJtfDo7gB6+vhy2mSm0DAdhCx4Gss7zym6
OeUMcfDbTGwRmJBgo6vwoqqABnypcMjuqeSXdrQ4vDU9NlZFi2ESue5uV/XYmhw9
GHG0acMqMSeEX4Aq0RwnuIRHsVLHSmwAPOukwTO2JGobFRkwGUv/UGxCjMC33X7y
Y3cTUuWORdZ+tdOFO+zsZDgbh7SqtfD1mp4nT27Ztdb6UXzIjfx1TmCGue9oT04b
WicACMqDyy2jFFf3XIO4okVT782pIXpq2HjrvHVCLepl0MoNPZUdCSot1T5ibIgx
YnecUc6BgHEQXWPGmK1AM0nfEtKG24vJ4NGH3oB2iU08EU8pAIa3l91Ch6wYLpJ/
lNcT9zNl8cyYreIeN+yF/bAbGZ3sYuRT0su6PY6RysBaB7IaaJ7Pd6fNPVMaL3FS
qpSEZO5F0SPOw0BxDQol53nkxqVb7UZGjlBcfs9wGysqOS036080EGSW/Fr1Z0tK
Rz0mnyhW2XsLOWfELGDgueXaAl0Pv4+mgOUIxStkrd5B0qaglisL/s6D/5/SA1v6
Ks2sYOCaq5Hb4V3eOs/b16Dzs2tyQqp+ERgSVyqnHPkfvGw1pAXiiOnrYPz/vE4a
Lxv4bi+kokSAR211Rn+8d22MMGcGIlR+Qyk2CR+qDgI0MyOcC+KVn6FwvBq/YhK7
Tniy8UW8foWnJVyPJ/KQUFNqHqg3kNcWrtWs2AcLsQuEb3ucwux0GbS9nQtFcD+i
M1awydYmRPMaaT+uutthPIx9Vtp/xgvD+YNUqjntYWu8+DuS7tVxQYVNjJLXTdoN
99YKE7qPnmse/ol/v3mJ72ZIHUsL9y8ZnwPK2pRx7eyFhQ5FMaPS3+9NSr2knscT
K1loUsjt7Lv3gYx1L9Lt9vjgRH6803t6KQaClQKtPYSESeK/+FFJP7BW2HEUQDMg
9cD4QXuIjZYfK0KIVCMz3eP/GvwDAFHJjShvwSp/ATUSBt0XQivmach1J3OBPjJF
NOvRVMQqEM8XB9UBouEsX004n0j2QXMYqF22vVCK7scY/nlCMBW3i/hs22P5ceGh
XRmlbghumrZSAo02aFyqew0RypkSbr6H9p4tatX+OvzYHq/jaGS0CGguYscoN8/v
hFLsRsr2lIiuNzYNxwOE4raRUQjws7IRFwWq54M55cwZh4LM0Th3QwLTTAS6szVv
WCNMAp2bCgKmvs4sCBKmtQ0T0dAMUA/aBu1eZPt9XfI0snmP4AtEyGj80U1FWfl/
F/5PHgB6ahOtgvmpnST1pfAS1LS4z5dOUcE62E0wEDsKACbuZ1O39nfpbxwtbLen
WagSgatJWnYgR48Iganr/xMbzJ3s+MDWrpk+MkR9ovzYKahq6vQ6qzSLWhf3ouT1
ef/I1pCzaC100T8IbDw1TbTg1ShZ8jlpSBPkr5UZj8O0BBlptcxmod739Xws80IP
9jus3RvXFRXTQvXEW4ghMRNd5bfjRY9KlJkiW2vGLqGFXEqKmd2EW7lrCCtZY/Wo
YF9IYhsmqkChZpHelqpiVSfqAG3IJIBb07agZapGwAf0X6bz6p5VyGbOpUvcDWM6
63VttKN4MP+7sJ0qfnDZyfiTEqjiGCjaDn9D8CcR7x/WK6BaJ0he3Sq16k28iDie
5zeh9vVa4cDWV52p7Txj8TiaQ33N9h+Cn3q7YLUeNBa1ShVjg6vDNUOF35ihCWX5
UP6s4A0OWVsbcmrgJOlL1R2MKhgJz4hdRUjqQIT+5J3xqUreTkKUykIfwiBkOquF
bj/TvA7KQpeX+JbeEetk6Kl6jquEm7KSdDVZynKVCwEKyBBENIdvxsByuhkYdgci
2NKmzP4KEPcVVFkhdhq3UKFjRdOljl23Zp9eWb2my+Kmd1IY04D7q2fGSkqBZmat
HYSyb8not2hc1GtoZ/QZQnzZV5S1vFqhxvt/lrDf41XU/Jxpg5DCO4C/wpNUlCfu
WYy5ApU/C3LikTlEguc6FNU9ImA5zyTOqtT9N111YGC82rgTCnPZ92m9ZGVmLaZx
xlKGqTkxhwhowVcR72lY34nwhireTQVaY05p98gqo8E+QmJrFLpBJmqOzr1Q2WuZ
AsNfcfAb5C5xKZmkVLGU0Obl7RWH5XJNASMqp0U2X0FQaaQNo6ivaylOdNnAIB7X
+uA21Z3hFPqCW+ltxGgWeMVGmVrDKvh+vVFKlWSvroQJo6mbTuSh0lbF4zoN4sVG
7vUZqIoQG1kcAF1wEIKizrUJ+x00vSCqGOPzZHYP5i6hZFAjzNYXrLH+iFDgELJH
zzRo/nlDFU/vVR7UsE7QMMPtFbsfmsjVHjQqGZMGp33Xe64l5v9PmyKb0yXVsalA
XQLpMJCxeFFipVCBuJNVudCxc2IoDEp8r7AbbTNhf6N1Ofn25fj7fxm5dOUhedRe
64K85t2iZzTrtNauJxImoPN6nN8qZ9SCZ6qkR3WzVP2ceK2QkIaMb39vui0J+5pt
ePWNSZDtxC7G6WMPT8NxjwFvps18874mWngU0WUn73wK/2wMDhn5r8yyQDWosAPP
kJvmWdW9mCKnOzDtCpuHhakAaqSXZhAC5zITA1f5ay7ORjQNVKqDXkurtiPI11rV
tVMRTYmzx1AkAhkwP4fSRCc9cCSvML1blkK93C/N0jP1Oirirg0fYaAAjlxw4vmZ
1L7d+gcew0lb9X1p/SWldUeMGBw0mOriQvil1xF0Y7y+Yuro3StqWWGmH8jLGSeq
6f2nrkb5Ey6yhQuWB60HjpPqnb6rEtwOk4bthUOmyxvU/SRC6BsKg9V4fXmnjLHJ
qQ7UVcwXc+B6MpbDvTlqjIohtS8s/Q4RVbfXG7zrXKH5DI1Zri8J7SmfLs1lgmXc
d3JWXKfDAU/I9RNZ5/TDxrdKClD11UZmoJK59hVOEboDtBOAhq2I6Tvb/jJKoTR3
C/SBBrJFgefZD6uWz5tYft30OshskXbqVnxcaZEGDMkW1lVuapG4Wxeg2grHUdko
i43qghcYqc6Ij5nI+mv3kuLubQ/KppNExKgrfECCXX06ULRc6z28ywwQJI8LFX/g
h69D//+XoDIq/nM2ShB+T4Xgq69GkguciN3tyBwdfhnYGj4J4RyVtX32z82ocz0V
z0C3N9ZzsJ5udGdedgqRKcaTBxaPbr7DLZVPmjV0KPReqatsN3FLrVIUg2DFJDfZ
cCj4zA499C3VA5I0vCUn+GJE7LAiyVhKuuSNe8F9/Y43EeXLrvdLby9gHTjPXhs1
eIUYnUtsKWw44+ey7sYcIXuLELIjwE+nrtZHnXltYPNj+zPBvQYc0AqiZ6AwdNFz
9xKCEuq34VZ5ajIZ5q7RK4wTfMAc3gFMU0Ak8CZd4JcKla3qc15uUOw07P2tDdfM
ABy532RwCPal7L4s8ZnKPK3QA7J24vs/yWvtA3zXFuomZJ7qKxfKrQX40dTkZv93
rvTvFSIY1yMq+Uqo6I78R2Pp8tOkWNl++NPDh44SnmNE/0wzYj+kmUzG0EPPr3r6
Pr07OtxDs8Cc8Vd24bE6bjE3vGpJVIeKqkfUXWPFHC18od74N6PicbPOve/lTR2k
1GAzeq2NIVfO4JxhDrT+sjQ6k4WEZr8s34A44bhJwjoTK7Pg69A+mvauxqqTAS6h
3WiGIebMQgExigGCIJdey1/Xkyn4tcETrYQPFVoJDdukMiGKZLNDLGxvz8DxYk+e
PEPicRiZeMRRon6AJIGQKavWsN0Am1IEVtYuklOrclWLvhtPFIuuiwG9b3DsCq02
739z2VXnMjA5Akbn7LjLphix7Z3hQ2XP1ZPlZOAHSA2Sl18rxUUwrDh7KGL9lqyp
5EzdsqRV+8TJz39eS6zmRyrRxTmBXzKPASp73WLS+82u66KFAdnLuF2F51BOOmiJ
TJdIWAswaoETNBPpN19bFzxSKdaD9sNAm23G7HomNdMOBoBhdmSJeui0gwSO3GHq
mjhBJ0JoKuqi40K1enO2/xwLVCm1zFUvBb7bInN3VweRpzD1o80luPrq+C3nfljj
sBGtP+W1fbKQauUTaV0BKesn4Mu8whUyBRjkbMrHkWQwVLOj957i/VMZAHEdVgoI
bM0F//Bn+uEVab25mMVvacDy827nFasXKhOPJMDVD76Xbq3ipKByV3r8PiFSWmJw
5Kc80X/37nc1hHvSPoLykoorWOtYT9uBHX5pcy5Gxez3OkpbALEZunzH7C3iB8eb
qazYE93nXOr85feqH3ECEIfiCw4DQw65uoNNdN8leVfR0riLQ+Q+jF/faaZYdznY
uBdjdP6NwuIdBl/R9CiCIqp0mRoPH9X0r0EBRT7gRVIXnohmoHMnXTMGOhZy0Jw5
mv1HXnBMS0W2ESpk6tJ5X620OAtLQd0rsb583r0A+760VyalAsaM+ii/CHChNCM7
MHC/lkdVHrv9b4emFVp6SBA1WDUVRV4b1X0d2VATGVtOOx2b9bpAFysBDQmtyfPM
4qnSGuZW+w18poaLdgIS0iLTda6LXiZNOo0hC+QeiuHsLPagU58YjHKAJ2liH+a+
aTWtQrmHoaExMFM3zxgn0iwD4YP0MgW+z+p+bw73tihJ8kMApeZSwr1KkAjksJcG
/wXsAj/q+ml/0feIm7pdklUgFE8VjDqd+g0FNvTIr2jIU6/BbH/VvxTUQRIf8Xk9
XqseGiE26KuGjuyW6iGB/t37XxJx3U6waEsd19vWN21DiUr34WQzTwaf4Lcmv1Le
rsHfxGS0J0bIDoSY0pfQov0Y/Cl7z4TL05TC50fkWVHTagLoKGgQib+xzPJdeuPP
sNX0xAgdW6qHwsjxhxg5Bre5Atq4I/wmklemlhrbQsVLMT/txASR3r12U9AOElw0
uaiOjRoBoxytWGiCBacj7J4+Vf8EVBhXjUpStoqpgV3ldTCJYDQP5z8/RKEMVBs7
uOZK5RRF5Zb4WIGEUrrBev3VNt14fP20C9RCNUC4wFBMZFjvUpqfiJieSLT07tVm
dJct7QE1rGp02PwTHC8/nn8lCuJau8Zn5L6J2p3PphFtBwoCiDxtvCmD96PxvrkC
RGkUz1CUxXhAyHBBAATrHGvCEfdVIOUMBTjVgG7Kcy4zMFF3NYUPvr5gVpBW/Z4H
UDI715oMP87TcVX+pqHkYfyOJFGHF4BGPXIFmHfOP1fzL1utFkCPF7jCP/yGETKR
D6EOX62Qt3Ds2F+qqrtI0ImkCDIb4xKRSuy2Ms1B3Re4N875gSO/MEzY1qzftYuP
gE8nkoApueL/JHe9uTSOE4y7MPTFKrOiy55owgb+7eusFg9BCR+zVahr+SZw1A7E
gy9Sxu2hCOo8+Pj2Wg/XOFxyaYJfF59qDK4ITiCqDnofwZ3K1xPLjhLriKPqmB+I
+DXZrIw/eS4+0VZ10iCidUNgiym/p27RgkdoaEXyAX3YKoUe3PCpUS9rdjGE70me
sREGoOzLox+C20d0Gj/VsctgZxLkI2y098++9NhzeV06fiNSeg6uHeXPwUHxqaB9
ykKFpU+Ml7IxG50dBKZSjq6+rJT9MPQ5oYv79acQ5BUB2HKh27k/a8mFzywd97mC
8vRKO3IQCjUBL83JPFmSwVyeyXcmUPe0k4obcAF57+TrSqX8TfdvIUvHRCyzAOIl
o02ImkUIUer8eFkC1IQWoomqYlNptIDzlTjYiFx/2vr4KFvvfXkQYqxqUWa+woBW
ndV4B6luWD2Ws6jsuyGF7DhLTjadF6VEN/qaY/L/nkN51lPGBeaUKHQNUonXcdwK
nDq78LXTttlYA7dptbJnvFgKNCFa3FML+dnzflXstffuMJX3yQ5n7gjqSEzfO2yP
tMVz705utwY9oN2EG0jqUobV8rp2R/uDZxnneVprO0+S5gSJ/gGAFiBJsZA0x/Nf
Bb+2mi5oT3dAyOYO32wEL8Fh8zBIoe8yMc+QQyV+z+y2yTvIu8GMfDddlNw3ePCq
SsKX5ssZUZi9GNcM7LwYmOw8PvOhmUT5wgEf+xc6miY9HlN+dBIPSb1a7TyeVTK0
U9ttjIUZU5YoG7G2sPDFlEDdYGK9+85+qDO2QhKicMoAOYLola6CMYiS2BK1FMVI
VH8pPcFNEZTbYo6yooBBfu0+ZCJy39mu3TDlSNw1kMJTGhZqNJgNspRLQM5oByfL
JNQMjNuka7Qx1MBzlZWpsGiRFHdBcqWJm00ym6a40X1eXWYYVYB4V3VBjTZ9gv5D
3cnFdl6yU90RrNudRpLJMdakzW0zhWgi0QRj9HLwKHPdGXv1k+3HO25dtfc38o+g
/87m6jeZz+5z1tuOK27mOUgMafWIVFvK/04KnfGBx0A6PorOXyS9m4/PQ8MA/cYp
wXUDNwFRf8Q2ZrEXcPQNeh6XKFrsW8bZ/i2Ht/fA9WepOlOshRWjqAkFxvPlBeY5
lnL1v2Fj7ym/cQ5vorRNOEOKvnkuihQUDvyBva7KKLp5QkrGJ5YyVVbRL595DuPq
2okFkjC1P6GC/3W5K8QXiq7oQqo993JZRl9znvXwE8r/XhV3551y3omHu8kgEVvR
UAtMz+ee/VPnTkrx+qbUJyGATyIfMW5aqUAEuKsW/wr5/CZx/nEfYlskjJXMWt7I
6J13dwxusKcz3zuxFvISaUIGNpuhrDdOktaYY/p4Wc9bbkmhzjMf93BhwdaUkq6P
DDpRWDyYaSXq9ZgC3WkfDglRm2VUfM2FkAMjIKU7v4BjtWmaWPc4JAGt7C4jazfM
h/wQFZaecMlWWtYVlsThn6McaBLoh47STaGJOEwaDsljsRmiLooCatZP4z+Grav9
7Xdm/DCpVT016xD2ZjGrto1+WCX+pMZjiYF2A5UB28v1Ju3HZQHYMwMEswVrJVLg
eot1idfaXUyI/E35FbLU76qgjK3ybSgiQIIKaJOI5uo8DyvX6u4ci6sTjkpUkmqo
E9XNYbuqbAzOEofbyx5bYjiEsR7uChhRc4fLg2lnInMKR26OyHBAEhp8PFU051iX
9kNNXF5akpSbwD/8NV19JU/s8pZy6tZ+0r5JojK9fGfhYfY2wRBtv4BgxlOqKrDk
RxwbT94UOH1zccM+27yfW5/9b2f9ZAhZD21dUBdo3Mj8JSkXtnIUt4S0/fMIi8zx
s5j4/Cp0id1wiq7K1o7WT00wSKIeDzougLvgSKaF07RmJHQH75XG4LZbnRAbFFLN
198GOTEu/rR5TZBLej6am92YbqSL5iTDZZ3QhfjRXqyYVfb4iPun1TNS4mtwTBjc
+HjJ7IO0dzWntYGAsAFCT0RCc/x4tM3Ry9Yx7joSB17eLgeEX1Zw3IQAMTvpV9Zf
y8EAveBK3OwMpXuQMl40J+rncc/5peRQT05tvBOGotmAeHotPZeh9PIucrca5kXr
v0di/FMpGGGfLm8INSQSxg9TlodFpmtoatCOSkHIZjeuboxse0q+rrcq6/3vIHLw
Mfe9JPPejiNTsjEsM0OKoh+6CMFMd0ejxq19BzahaAeecQng/tE7P5Xk/3ZMkHnZ
iihq5GgAcGtqnXjufN++/sX4VLhwDgdqGDChcyT68C38QbRjBnS/ZkdCD2Xc7fTe
rnRs1bOEQ0QIjqaqr4ZS08/VDlujyVOugu8lmi2B6ALfmtAgfMk5LIm6MW2EHL78
T0YyD1Aag3pqmLpjY8sSL0MZWFDJD6PFrTcPJ2/8JJ3wiGp5UnLWXPgHg4EOkX36
lxvSuyAq8vMWMa7sMG76egrIgqnpaeKX9kZpdTf5INpydAch1M3jZHwkhJPYqM0X
71MQOuQ3q5eTDqoPTFnF2mliAO0zZeGj4+AmznSR/OtBIjfd9R5ZuWGY68MSCBVL
amSk018kpRBzD2WZ6DG8cLetjHeUS/qfgTWqtl8GzFBaEaAqqsQpuTC8DkVh8yVT
9hCUfr89NWkqi7UMH59nDrllrEHuLKz71te/cLAMml5AJRfcSMpm2iUDzgSEFs96
+elLbmRRbu/CZOJmJINyBnW06CByWdnzybQKK4scEHTDezWpip1UQoyi66c58d5b
iRxseoCuhO51vGp+Zj3wWzq7UOR8i4gldHfn6A3mNmRbM4aJ8ETpRz3eYP5TK5xJ
CG2igoj3jngJh8Vz3EeE9PRPL1iorTbz6z7K2e3f569tpVutgF0YiImOpRM1CyAn
sOLfwsHGbYjDsSXUx2Luj7qAhjtSv9vgh8seYQhwvGJwJjvti3fuf7kbvRdOs6BK
18vs8IXcLxRaeXRi7WEuI75ai5wt3FKoa2wzdGZSbYDjWF8Lu3wcNpOd4EWCbTsc
Sgymo37uW0QtR7gXXk0T3MTASKiSCulEZal39TKp3W1Kb7GUg66KKcQDxMZLK6W6
CAl1GqAoFL1030kWFwo4HonpA8Q/KqG+X5dCO2+Bvn3cZ+/Ag30vUprJA7m6TRCo
9RdHfslDgxq8gawcjfbj6b+quC5ohS/Cu94GNPu2rbppD/dvditWYyUGYdy+7Fau
WRsm1uhYhqFD/2Db+7PHjQmd+w5dCShI/y51ZFdGx36Aok1U6oPQSEghSqhJ2Vqi
5Utt3xsFI0chAqhVWYaaq5l96CXl8ju8sFv7hJbjPd0YhisJ/iCC+D1xmtK94dlX
Bsi2MW3/xVXO6xsW51+HeXJWe6WlGy5/fqI+XyX3KTCBnjj5j3/TrvizhVT2GRN4
PDDtgxpqHLMndzrbGwMXX7Ol8RDDnqOE1I/9CG9H2i/2rQ8EzSIKAzZntm3+Z0E8
vYB0B8lD9E7fRXVpPx6zQQh+WPDndhml+qrHu7YBqMMrAan+ZpXMtayiG2mhtQDb
0zPBach36VN14F+YNPWYFnLQJXAbMhwaiAqiEtEvtUT4Tm05cr/un5CsqCcw7MBN
7QbhPGszWgmzMWLgY6XMsedHFEnM0xuDPIdEsV9k6F+HtQg39QRXSZlaGTwTwyu6
qmkaQtAV7qzpEgSQj5vjnV4XacV4TUHDaMz1+wW1dIl29Tn8EVEwmdq6RcY93NXk
7UdMcdUP8+06Q6S9VIF8GS9s6xYiIZqH1/1Eo4oyqdwEBEKASr8Fz00MEqHEqpUe
nZ1EG+YwUlCN4lSGjLlWUBM8z+YLC96Kg9PZbOedLubx/DJX/FZ5wBwd5pDXh9Jx
PfkPQ2865c/tnNnxVBCZ+/QH37eNA+NTza2d/+gIBd0TI8BcLFaXbpOUGpSmZwX0
JlmdtW7FJReS7EoHxlbn1CcTJp6QrfspcSgSd6PrghIi4S8n0b20eQLWIFFPrR3s
ik07zbirVKL1yLmA4AuCz50OLcFT6V/ZbBk5rhYLhiGMJxRZMo3VFbtPcQd/GkHz
6l/fgvmGWqcIyh+CCyiKxTvnNnSFkSICzeCatPJwW+L8yC1yko9PtGynKoa7NZ0Z
8eBuLEbsPzzYNWi8f0ey/6rxtHnrCd34KK0DoqAjXH7nuTx6LZgDFeFiGu6IBkxG
kvua7vP8UQoqwwtSmt/c56xDLYU2qmSii0K/7V5a213yow3/1rAmbWHt2bHmpH6r
h/XJooUwbDexeBRZE5UPItg1DV495JQNTSfuMR1hCxQmgLmjqn3GrL/BMuLJV5Ea
L85UcdpPH9zbUiztbsQE38E9uWsDTWaFNBtr7P4ufrqBng8vJ70U26+ZRtw0PJK+
U9ErsaR/GuCAsxsAU2ZD7UaA8S6mrn3PbCvM3D4XLdE7lWIOpIojy3xMTfd7Gy+N
5gBIgcAw8+f6UX/c0rLxvFkNU3uwABOuLDb0NqI5FR9nv9o5UHMaPIdGy1A5QdsS
9Zq/x+pTkn7TQLa1Fs+xPrsdZmQQb+LbXotwJJWAy5UIQnaZzFm+y/Br19SSyE5m
wQ55Byu/IQis+uhhFFR0wbjA8gOI7LA6JTLz5zGp+p1m/Hnl2iz2FQCVc8GwoYT5
84CxrBomSpVJGf2BU8YABehPGkHQzv+W9h+OMYn5Naqd+RQOKx6Uu/1x5Z35K/i3
0Y1rGA70g3YfkNv26nOx+zGbucnvGSfydol28Kud0dEzkgq9rJX9x42uzaUQCnxd
yVNn0oS1DsvnMH52EaXpFDqoWtX35nj61pGoG/tBLOWHvwRkbYFKVTUd9Kcj220H
HEPvQ3D4ceSxl4pTVKTKE7rcfuVzr6IiNsPg2amPO6lQjAGvFql8jCTBpA5TU1zl
flDoRGbS8GMJk+7TxG2QToPgAPWFaY4Eo3Yt8+wyH+8xx4agOKzZZEtfKHssFHJO
e6mFxlXeEHcBYBTLuA0eHqsFP4idJQjNi+0muk3a3G/iQbRrmU+b7k75ze+5+oc3
uXZ6dv/tiN+HHT/MdTwwbZCy+fHgTycdeHqwifK15rA0oFO+Stp6G+VX8PoKotaL
uijLQebxcO96UJDXnvm5ISkceMw21DPf7PkSBEjlzfOYAlNlxJgh/NiEIHAXGdSY
suBJvhEd4PgFlrkklvqmh8Y6j0nRPT+jnQVnjJt43TYvFCUuCLLhk5KGXlsfZD7r
7p19B+Edvr1g8+1FqXVLf/wqU+Dl/hJcQBIl3rIciwTbLz5dM5MZcAftUv09H58j
17kDSWStRJTonlPpvR3cBhE3xEJ+rN2Z7/rTEIwjazTawtA0bVVCkKv8IXOjTSI6
fuuPUgZ1+Ovpv8iwcD/Ulitz4YbGat7KJopAOdOptCCMzhcYFO02kIa2ywfBHHCY
YveCJeZ5xawY64L+jMLyhzNPMJKzDaScNxv37TkLQVLI6X1/V4u4sixjse67RfpV
CNekRUtV8zEeOkDITvQlAy9vDhyPk3P8JNzy2g6IwQK3k0fdACzUJdgUVmqVtl44
hhkiWTc7wHrfbgw5IXQy8K2aBevcMWlgWGsohQ9JsluS1IpdW3ZQUabWBqNGX+S+
YspxeV1iHAn9J3+R7vLV8vrimBw4GhMFJhZp5FaSp1vhHSv2oDgoOERZUvE9FMZ2
S9LdIZnuj2wYPq0X8TXGh9f2fyFwjfZTdoRC1phAs8bgd156xHXZ3Z1HoZywmA54
jD6KSy+mqEO+fY2rxX4ntdQaLmW043r26p1ZgB/yn15g9nuC8+IKRlBgwyNJqQNb
nneSy9caF9HVWKQBIK3VD7fnsRs/r2w5mQIrt2bTgQ6xiS6amt7vs/qhpbJCFhuH
J5xlrruUzpsKPp6q98XWmWoDJC6dPdeR7n50JXW6DnuYyWgs3dFwWzc46jMJGXQv
18le+uAb3ha/uBA0HUjowC6YEx33+zPINLXYYs6B5B6AmyLZ8r4khZPRHA3hg9sD
Ar4CAJJZjXJBB6feHhmbZDhhFbIYyTzENhOtrz7iBFZzbtqHEtfZtTJgtVukTZXq
AYI2j8jKDeIsnP4ALUJcDsJWaYe34ON+4ZlWGTzT9rPHwWj618KVuQD83/wQ3RyM
sdcFOSD2KoOs/E96gGFFhYOfq/6OWJ/evBrbXfdTcktYM0kPVPYD0ZEbAtJ8asLl
MtCqRfCmwZN4LUcLQk3YEt+H8NYif4gMvoDlWdSlwm1m+fCKcw95xOS9OXUorUg+
6BXsq0uIAngSRC6dTeOgYyp8D251XrT3RSkNomoLBcDN8JX+oaw+XlarqTEam/1+
R+QLMiIHfxTwX60Lmqw+e1jusr6aNDTT2TdIFMAict4K6FTYTMY5vE8M/qx8cRGs
7vaM5xp4FCtJxn4v9eMfmfcavSe1/zFM0aWxvBzavJO5O/WLuoIoguEgRCvFERFo
RXeB1mEMjk53J/ore/vcqmkYoNCTq0tsPWGysAotqj5zLWmGFzHExlTbxqi0JyPR
Bc2ryZmZZ0taaZ178enRboec3dpaH/e/N2bxHo4KYoBQv9HyMm33v1wLYewX7C6b
ak0CrG0sv9ubDwTFIx3hNIhL1u1Cujh8STb/S1C3o/RoV7ScEplSi0KFmzeFK9vZ
KWW/b2BPD1b3RLj1Mk85cpp9ecTBLBFUtIoVUTXGMAnMDHllHL1YpgKlRld/M41W
HySq5RnpKanvJJBhyrZHbj0xBEKwZgKxWKOkymGzAjkSaK/pYF0Jt3BOFf9p7DtI
T12xrm0IAoaBn06W2mwGtnb+op635MzxkcTdFudm4zW74/xCSZzNcsYkBrk6mAl8
58MB+24AL+TRshN7qDTkKR6c9/JhDb67WolNjAbiA6BYMw/K9HdGuSZZBhv4rhbL
GN9Kk/uS06H9N3OLNxNpm+RpvMlyrmQrcofpaGDylDT/DzjRf5s2MaULjjYh82Qe
qzjGjbupEz+r3FHb2+zClZ7DPUFQosz9KTgQ2J3ZM/k+nL1O9hxKqG7sFvegtpHn
3uorTZLY1U3GvICGkw/TjfG/J96jzdlfql7LUAUjBjvQ+pQHcKqsleAvvQK0s7JW
HZWTChxmvm8ZyaPc9bljDEJQygPp9zuqpTvPTpdG7gLUIKifixX4BgFoRIFu4z6d
b/sbIzIOsJPrZ3k9w/ZoOhgt4nU2C79JXaJzIZ+Am10EwtfZ9HXUW59VF9SX7Ajp
ue0ytfsnNaUyhl4pglfEAYCfxyGUF4ZlwmgUC7zdYP62jvqzYyQ1hgHyKcCwJmI3
HewXkB47t8hUSxmzyrDPvGDgnuueAVIK1Dt3xJiozH6j1AJ0W7s+Pr5WMKIh4pBn
gkuB4Pz6fAQd1jjd+R+S6ZcrX9K0Qoc3p7IZIG29ry33FSmGXFlycdqGWyjMlPdw
huHcxTvz2kX3Z+j/QdxEZOapjg427PiXrR/XC4Ukd41+e72kIJB+mdRW5ymzuDPk
Vx6TxhoVAe57R4l2hpY8aPDbW9YRVeaoDFUBEX+BGKhZs3ibgiIgQritb0f8aWhE
kzzlxcLdNtWZWhDbcRIpKgxSjP9vWX5mXXEo2awPjRNQRMwlXMh/cXDh6ToKV5VH
dHz7wNXTbiYkE+sDPr0WdAJkKiV9wiQXwPRlMGfReJ/Kh67KyK7VqVyIrwlkkuLl
Jj8v2FSoHGQdFKSt9+uZ5SE2VTeubClnYsKH01W4uTY0ixg3UIXG+mJY47pa4tPi
pn/C1HJQqLkeN4J34CPEO5OlAmvkHXU7eptOzBzgf1Ejrq/NEYkxEu2E3b8uUlpV
18vLGlug4OhNGAa9J0DK57Pl88DHq68MfxHFUPjcFGgR94aqy7JHvcbKf6ymWIQS
AibEJochVZ5d/KVLiEF1C734YgvIqlxeg5YmJEpQme2npKyeZyQnolabRrRizaNF
4sr/06GBEDA4zQ1gHKEimeLbjXqTsrQP01MB4EZjOu8lk2rermUgDT0IvZQjO64F
vNk8+8xKNfFWuWnaXBwRd0brTVbDvM444zu4uVgWT32lDWsaSmgz29wkbCCmAiZO
5H1q4LPPnJPeBPnWIEo3M+JedKEj4H44FKxRUWh3DlrFEX68ZgFi4M+bAc7d/2PU
9+4jjBYmKMQKjkGp/wqWl4buQn0Op4qOdOXVRqDuicfSPB/pbl9dxvp76h56MRg4
YYhi9A7MaIXL4ZPLI6Z4X9H7LN3cCKEB9/wsBdc0q7Gp8M5L/qKEoxRP0ZhVgv6I
ZkT8d5lhmaTDjXl+E/qiYmCYFKZNLxqkLoQL4yJQEWxGnwlA8HMP05wTOl0MIBaC
ByjvdfaDyVIz4KB0rSCuhkgxgka+O7O87bxIZ8I0x4XEIVjk94lmDUjrpOcP4g/q
0/JHVT1lc07pXOgwyLfOBEUpSG6yzKyBmsknCPMPNihUsR/L5j6efnVilUojUECK
v1bS9yTvKoaddkMbiu571uZzSmSBxZ7beq4xoVjNANz8Y1XvE0RrijTHW2SJN8o2
JfGWyRXA6U0rj+etcLWB4DhYaT68qjfQPhcTJtk/h6IO87uHdUcIk4A9FOw02Dma
dvV96u7hvx9hPh9M2A1SLZuQn32MLA67YfzELpFgesOzzPWQJwLIELh4o+EO+sa7
uQqKCWMtXy8Dmbk0qsiZJb/oqeBsxaBwTI4y8YHBbRAV2w0LKGStEBbXFHzRGZQN
wNnOFdSQGUQ0Ou8ODGs0TbWtJIlJMwcpY7EEPOCfFVj14i0bK41NwGzOFS/4fWP3
ADewCaW+Y2zhpHkf3CjyS9YwEjquGBEzkj0r0GXHG+nic5y5C4Hig9+uO/w9YXoZ
RVjVdtRMP3jioHvjtBMPuYurZ10Vy7wEts9E2Zu7QR8akSe5CjhIS5Wv/3qGnDfx
SvGtWAlgCCNAvG7BPt9S1FrMYZhjzvRkAhPqEt6MNfwEwIVNn/kQBoXPWEGpIL5Q
dsIuqOOG4CxW0UQUQoZdIeI9ZgK4miKY5MZvFXq9tzS1DZT4kt2HEf2aATQFYnnh
FrXnk0bjXJ00wIsRqGPj26w2huVKxGJqk39iCi+VjR8nzk3rgD5IYKic43vTCQ50
QyrlnKN3ssBYmxPEdh/p6RBzVUKoslg4QqiYXb6fKBf/dA5PACBj4PBi1HZKx7Pr
2IOdwmZFcH2lFWmH4XwFwQwbAHRG+dPKNeOZ8Y6II1lrNVxFxN7y2MchxrELurku
hgDa3+rf3LAqvtOPiBs/T8fPQgt0FroUNwE+C4J3KFEzeO4Hj0xWywhnfpIJ4tIJ
NUssXHqhXoUtXUvpBUm1ie971LSqBKBFHjSV56J0F4OjhDJ3vgi2Y46y8z1lKgDg
ANEXDVcT0YzPuxVtYO9j1MOUp8sH4SaLArXNL4Oemp52rE+YgCU9jp3+rDILwbhh
oY5hkpBb2ZeNrUh57Bk/Boq166l/HABJdWsyKnuDbioOog4BG0yYzyGUu5TqoeUx
8OfcnH0XvoxAPPu86IHCHSt7P222sf5rYa6f1sFFEZ69v0FVXPEyjK+c8TYoiNJI
xK0oRHP29owOSBUYljraeKruFnwzvnarVpIPPbcdUYRnqxUOz+njc+/Wb8V9VSVe
qmBOYyTetyMP6gKtKv5YLu0PlFAnTlvbbMIg58DhGIwGEE8ZHlvVzjX8mteT81k5
b1tSK9JWbfT9WdXCEd4hlTa2/U7nZpTh1Wl8XH/y81fuGscRzFkZBAMXh5PSPf0l
zD6Vz8dm44cvFBvZynEy45/15os7AvvtkYQ+PLt7iGVolT3Yp4AaBxbRLjZWYMHc
DMlMEluut5z2kevmD8AFlX3FGD483Cc5/N/LeDDVncZGyhKnza48WwnWfE/gLS/J
WGgmjpqLkgP32aCXfmgZp6gVY3l9ZW0UmL0TADNB9q6mN8fN/X6W+TX6OfwpmVSK
tnFE6go7RJckcKS/Tcr//iBf2hbOLRekDLnkymlubV3Lz/WXTXMeMIhf+zJdTQTE
BgKQ/XWg/aRo5VTS9wno2olUqSGfIQxd+vI9oy8lJ6FRTMLrQ/u7K+K3T+9TgF5y
LKEo4Ssx8RZsf/wlmzI27tFtZ8xl2A3+/fu8OtPaGBdR6eNXsxXQa+W5GI40ECA8
S2Wj5Dp8fORNHP9m26bSkOUC/4FNroeCcKiPVEHat0WdgP1idaR5bzNSz+5hrUF6
qVGJuhJx4QYwYz7VgiazQjJhepg/sWR4v9Yu9C1RS0p2xk50XEXWz0dYUReCL0st
WvqQAkYud/0cQt+EKFeja3votS0qrIWCB6grKWZrFPP86EF+QFW9Rgi4VsWND4df
i8PR9Ov8mNmJJskReF/3EzHRVSGQIpY6EuJ2+IJUXf/stg3M5qBpEEHJmc6S+2A/
AJG+B1LyR0FPLjbCZfo2JVKVeOGHxmwXDwfBpVT4V8VmaKRU4s81Vi7EAjOykN7y
dpY/bGr1c95dbEJI67uZqwi5WQrug9iQV9frmNmsDGXS1/bWohlmTa0J3gwdwHJu
YYwmnCgVYxdJgeZ+6iBfHbIDpVh0fGQfGHbdjLuPP1xkgIbpIuib9aLXZH+BGVNM
zSdv9R0V5VpUrlRrNK7rM7a99TwwPB8XM0OXjilPcJtQdejEJxDdQMQ4tyV8g/uY
Z4NzM6cJ5SCOOGrvz2Pwun/y7CnYavFDRSWFGEywQHvsizHWoEaUCgYCwjhoJvNy
UL5cLZxUgkzFsJ1nFbRwooUAUGbAv7R7dmez9bKuBcilFGm+iPHvcC9HTIYIvJjI
ES5gtvVuMISGHPzXqhJTvV0zPvDvg4VlrMOO1hNV5YmyXXk8W0hZn8KGd7u4gbmj
n2yjKS4KQ+FP77j9214ealFJVcuzwERq2Gan0OcRjwoXq+Q/YN1uAAcqUCK876mu
nSUPbbOmrCXUovCPXQ+cIUz3pyvolzJ9GCcpbf5YxW2daPH/FmUvhvgNM4q79UZI
3inMVBUtdD93SZiG5+t8olg0KnPm9EO4PlCqz1PQKSdp08RBsAK8iVIG8ytRi83j
71UZZMrwFkdB6USc4rBMn969VJRga87j9cfDt0jGMlOXLGrVnbsR7UGDh1095d90
YmBT4uAZRbQq7uRBAjwZxFW7vFedqHPh3hkrjbAxosdjhxDsTFnpnd87JwQN9T9I
dwjaKK2Bvduazf5F13qBqX0bU1661CqxUrFlrMfRqQdMMyaKjw5SDMKoSgtvucs4
9Fjoa0bgDD+ViBvRWPEe6OTFc2yXvL6mKYxoxn7xxgio10GC/Buit55qE8lw4Lg7
0s4MjLilcHQ6vwbZjmQG92CBoY5jsM2CbrybGUufGiyz82dDVMiDhdtGOSRyc1ju
+bc0dBWCTA0x75PdkBbmjalwHC5dckjU+ufy9H10HoCEGgkymg6l0K9G/SxEbQon
rlLaVBBKhQlrm6bylOX9rVWcP0Q6t3+MNk3QPXlnfaE1N+TJIH4yLepoEIE4D4yD
BUlfpbvqeJFEt/seDqygY/C1w9wSmIXC7gqZshvAZvcB0pxcSkC1mUT5kWh3Tbq5
jl4KOL9YsC+EaYG310iigtwuRcubVTejVpHDQY8nAxDYsR9n4ez4TfepIflCSdvM
u7Iz+A5ohN7C1LYl3rxquOwkjRX07pEHXdWTP9jGnr3CJHRKgWXeC6VmrYIEuIri
N3infjZt8WE5CaVwipn9RRK1xy3xGUgtvdfxvZSiWvuuJULBtU+6zG+yA1GOFnmf
9ZjxWDvN7vhAWyPQln1M6FFUTVIf4Ii0xVDywPJ3+6/JwgKCNFCcJttEA0Wo+vER
gQnEz0bAgxfP3dq1/xYe7TVboGToXR/LODdUnL4ybH+j5kh7rAo7x6B7CzhOubjk
drq3LypJfQ3NiBdUM4q0fdr4mVH3lu+kNa8eBm7o0ZepEe1+4Ogvf0+yZ6NUlSlA
92SwEj7KAMSU5whFFdMDV8vHC20wd9d6cqblzNf6x+a/5ctDvdHAbhQYoXL3fD/D
JVWjtLI/J08NamNy6Oj5sBxQtr/M9MHCj7IQILaUqeYD3QkbiPD7M97psbhC/ZSU
kOo2OeNxsgVTbrrE/X6fqY76+zj9cXFra4tAbZ+IoLYbJV2mYAKz+w/N2Gikertf
WBh4zVd87EMzRuzmLkXGM7tLXtHtg2qk6sE2v2BAl9lHDzVC3MAOxLu0fC0CiZks
FRt1aRzTQpPr9RwBpINH0iBUCjz7pSs7aZN8FOSyfk/igdD+b827+ESKN97oXr57
ii8XvWTcq77+Xe3PNPeYDtMvohNilE2XcuTuM24hVIbf4XsxhXO4TssLNzoM/lF0
ZjIcyuwWfIsuwhez8DuvJEoH/eIjKWoAOs22HG20Q3gfGgqB2qHK1fzFfThucAzO
o11UGY57hJgXng8fEMugxhtpy4IEEpXdQSqRmPvj8HBMTXAUIpqu8ZTvtkzxiJu6
NzFZShQQufuKvXhDSLW2haCN9sRgPX5RniKOcm+HOyhvSOVvtoCYP2rP8CXVNJFz
NiwiyNQOmTxZ/IBRN3j1/DhSRUPznn7HdqinujpHshcF+UtpdTnTyvzj7JEgm/ea
jXcxRq8Y2HXmN+gt95EdEOndoxZ+rLQ83xQeq0xUGMDfC9l86zX1u1/B4lbBEyaz
drIzOFSUnnkSSTLxml29qbjhrqt5eBLVLU6sac+66DjYUnw5PALboLpV+DXcrOU9
Fbxda7uCzyVJ0llwuEdoLtck4r1hV7lc54I/HqaVAYa5iMOCvseCPdgHNq2e/RHv
Rz79kiMt2wpD6Fs7Fhgz711uWjKkijQtXfM7eo1/m3ilKYxeKdrU23ECPNWwFL3R
b1tGf1mmUBtmaSoH52ITZyLEArEjTlk21Fxkugi1uD7jc0isTninzQ645hOubZAi
CFibLBAJjV5tGz66rwv+yzbSPC/im1YB3XlY3vFY0LKLCVSjfNTqw2hzNzJAY4Zq
5JrXpnrwHCHWMl+7iDcd5KB1oXlnam6qJ6a+XqThS5Kx4oNpCnhsYbzAqHUrKbBJ
M72WzWPYjNGhrKqRuD0L+XN9aAo/8RnEoYFlZj9IeXTNkwtLoiP85MCX73H+iu5Y
LeA3P602dyGo+Lix+YeGa2R31hyrpy8JbDypY9bB7N6Qn1a1SUQte31t8NbI4gS7
BUXcIZnY0Y5tU6lUhVSiHzYpmzSGkou0Bg1ugR6OslodE4FkupUEpxEzbxohLkrC
bub9+e4wofib4m5aqpRTgXPSY7Zou/Z56ZEMzdySPGr+kSoY8bxF/+uEo5B3Wasr
+M8XqsnolvhGA59YNKA9YuoaIYWEyTk0mnEi+iZ4hlETsgo2Jg4q5U/rsfScJ9Rb
m7bJsJLKMP8LOfOrNRQRy9pAzoTHLUehe8RBezMWCu64XD0hDJeQ9yLOf1LmF0ke
tn7eoGoSZoemxTS241CfQR9QoPxUg86Yi7hG2Bk/7HnLS5TdkZMhil9A32qA538l
CABSYGgb9jD3niwx0unBxq3NksPT7CiubOFzoKaFi44F0jYfAWeXjJsIg71WLg8H
cfAFZmxqlbDKnO/ZAEjW0BNPZAigIAWvjwBlBpl5sPRb62IXyAKXEs74Gsqxfh8O
300DV9OGDIAQnkWI4JC0GRhxQ5vgcERzbbxzWzWYu2OUGLf0tGFD9/+VhELGEaaC
2VubQWapggGB+jhnfeFGM5Dvwp0h7UijVc3bFeUAeskGxp/NhUpxoRMa2cLf6zQE
1ozIjzqa2cOS+YNThiBalk9+SKXOQQ6rEI30wbuinmqxLgrnpknWhhP7uhJW4A1N
DnqiZVW368xz+fhuPxxQ+ObsORHhfgMGE+5K+2rtEkmP7h1YahOxMgWUEhDYGrvX
YvbyMKkTcF6MrShaa50s9Rw/8LeHrOvJ5jXAKplZuyWP8C1RaHEVGBPLfkLG2kga
4pAhnnIur36g24K0Hgz3w9fvD5W5wHi997at9yEbsNolKWoIBArym5yfyxHqM5dC
N9WmCnfZyTR3UWVTXnx9xcASyZMetpHxHtoExJRGqzo9OZI7A6qtOx12AR7zC5tS
OPUxzBy/zzxy5rH9DnAzN+J5LSZufTyfPEYqtfhZDNW2ANbadm1XyzwyGKbM8ZfN
UoopzLfG1CwEnLsP/S2HWfgu0oLAYI9ZytciVyYapAhh1n3A6u9d1vzvdBADDsMU
cCH1ZRuycygbEFkBIHsrzEjzK2VxtMMybXcToetnf7cdJhfqDuZOJdSGqkbBn1mn
pdhGXjQN74T5px1THhuftUspSYF0gKQ3O/i79srs71RX7q+Yx9oQzZojoOGRQZuD
yDEqv4DITWWXrmuyfC5urOboQMO11wfX71xSs+0GkQcizbKciiaIgi4sIfSlNjns
DsHQy3cEBj3RO82utvXriGRFH+MW0o4xRv8Yxz+pwl8a2/zAc7TBscqyU6s/ORqk
s1rTE8yudSZhXVV7bfuoRzMTA/prgV+T3xw2aBQhWRzplBOQ7jl82Vcm5dzsVeqC
nRM1aybQ//4t6al3EetDRzk6RTBSFyDTpiJNX2jN+70R0/msa+kaups3aExdtgOX
7/HY6qLmlGKrnYNBTGsYK0KxOLtC3Tg67f3nQ2fGTAKKjSAuF/mxELpAocsEVgkr
tlVb0BG1zC8UerOpb55MgtlsZhf93tzyOQKtzzozPLINupEDYQBhK+stpOkR4hIv
gdwpRoWD1ZbO50EN7ClyTIaCiJxIk+xxsh9dAHvLjs7AJGXloqmi1sLqg7WWSZOx
xRkjG9DEUnXZXuPjbcmnghXjHOtDIryd9mv3I1c7w0wa5uf73JiAIQpwinc17WEM
jFWprWPJupy42E2Q+rmgZab1BnIRWpXupwMaso0XGgnG4J6oOzndEoOBRAawFId1
edyA4ZYTC5Cf7uJ86xgvGFmP/vRiMXMblchhugQMUwZIZclW8ESXonma/yBQQngW
/Uj+0kOozD196EwDy+583H3T+Y06qlSrdn6Poukdj69wx2wad1pzMWd7YCgga45e
XdeBCEAVBc9AngGEkjfdIZ0Zzj0x+ZmytzfOhZe6pP81DiomeQqtPCa7vRtcorXi
jvqhxVeMFS2YDvh1VK8c6yDSDNmUyQh12pwLibZGxwrGHrMFYBZxpjnf5EWMuYBS
ayNaQoJpikw5hX+wRh40gCU+krzw651ukwlE20wqAd/1C+/+4sfi884877dms10Q
e5m28tg1lIu8bREwtoJPZThiZalfbn3TKXRC8hK4ImBMgsArKjtN/pmsv2qwGOC4
0p/83CRxwxdxFQ/7GwPL/A+7ViyU3VbsC6ehJgNuYKPB5cBpEYjL458UKXElXJ7N
gbt2zHhyHr47/WigrgB2WE6KRXGM6A4v51cvvVyqdQx1FlHetLc+aSbRvOqxixVb
LD/oqGPv9BTH8WYJhFWJPfXkVR5Dv39fdtSQGZFtN+0tMRZ836veOa4PcEd7EVgY
ATtCMWhL+nmlQXtVyoZdRB5uXDCYfDREBP/2fBrbZYXL/VtveAziLVCOyJUkjJG0
jM6/AuA/w9W7k+mJuJ+NPtjGY3YKqgrwvkRV3PLAi8N+wy5vMAh7LqKNra7KE5Bc
BCI4Fitnbu1LR9kcMRm070+lkwlRMl3bPJcRpc0q2mQre48ZDukE2jMWl/NscX5b
IDmEw0OSYR3txWYiaCaJYd0Bo5qgbsJcxp5clcM6XcVbpcETNbrXfXDQLN/XmTd4
SkyU8EwCWzNNaOXXVZaZuwUAN5Qx9ntbAtpsJXQec5smVfZb1tPREQAbS8Cc0PVd
vTU61H6mqbTFzKOFunpEJrieTk0tHdDXbtm1LSju+poAIQY+qcOFl/Quv41NmChm
CquYaTvzKvaHQiCZWNhg8m1bmOo4ruf+j9E0PLpLHVawq/IRR7m653grEvDJYpV4
TOOiQygdcYTF0nD/Ck2WJkiF5J/qTA7LkF1K7o+5erqOMvOFgOjEbR2dj6h05tDI
WNeuIKpv2tol+5qepLiRH8cviJiSJxm7rM6L6sv7pd9QT+KbmpitGzyEDWf8+nCN
CH4q5BA9HA8yJ6zqUXuRR/A8+Vja1Rf/A7bqaLwFvROGU2+NfrHZJpgMKhl+AGgI
m6dt/vFacP/XB7VA/UbjiSGHmhMxJH61/jYq9+1jTz1swUjPFqvDg5A8FM6V05Xk
KH3tpEmNO1mlLwNfR4aiZZJ3qlqqEhWQ7Il1S3W7ci7veQ1qgpoaslntwJ/5ANFK
LVbSAwqZMknekY44XT69IcTFiIyFqPdrDNoJH9JLfeExmc99M2Wv0QHj4VKF16hz
27t3Nn7Zdh4CsgFI7J5wxGrX3UFqLt0iP+yYLmHlmNXwPCIg4jeCn3qv9SrerkqF
W5rTZ99CtZFZJoA0O+1p7MoDb+een0AOpzRjiOqT6azl5HpJlOrPb0fznnTOIOfo
2NXH2NEwa0c8O2IxUsA87HmgSXCnxRQdptl8zedfk+8X46IwZPoZO8bgEsqvIqkm
0L972uTOIoD5IZYicpljbbyaBug7PI1vrOAQbB8U+X4cI5jxvcn590ORZRSE0lHI
h2qFyq8KqDJhSrogp50n2jtfIf/MdJUEdIYlqNtL/YIepcTlNURRcCaQISyubv80
VzxGefdwoj7LPkW0AtwGL88m/7YEtHtEGsnHxm3AuC+cvxUd5dW6rQyJG57EoTsj
z52U8UUtGjF9QG2xfZhskqEs4TterAEWbOqpmIJ/GSC605UusiRJEf5iTaDz+cd6
t9pT0U4nP8D6dt6YY/8RSV9oy/2Ajkxl3hT7uhI6HQJGzp3P0QCwfuRSU1SCPeow
DXTePLfv/WNLNrUCtzRjXDdBFtCo783kEryhztbRptiF37jxjnTcnlCoNkvUpw5w
L8wPoZfAQx5OqxqLa5smA0ffxzm/055dL7WwqjKhn+Yz88g21yzBz6wcc6D7lm2e
Udyx9Mncbz32TADmSZwleikrT/ck06vbjzzuzcMzbyeevWowLk2zLoCilMVWq3jv
jpoXuuobWRGOWTWcDnrrGymyd3fUwUmjjbPYSlaJ999SAoASmw+di7jv+ZBUruMl
msbFH187Bo02cLDHde4rl+PK86DEAn7x3dRRnxemMxvI0q+zORMW51aJBP0hi/T+
J7AAqhNOjrT52xOE5mlqnJ5zHT6MqoaiRhouENu2p1OUJGrV5eYJdpybeDid4TlD
MsK/gOpRhfit7ju7eO06FG/fI22iV1RCE9q9Md+iVg8vjjX6YOp1t8Bt3cxGdZGm
5ekJNMVDo6T2gFNc9mB/hS9kRxNFk/g7GDKaQhTV+a6vRhUvTxs4q+O4ilvBzKft
IdhB2YP9v5qNtA5baDKn3mdwG5xNh95hTCZdsW2eS1tLIE/EbU61AEKX2r9rFAvv
46/7p6OzIKTJKPy4VftEl+dQqYsWF9DOwySdoLxhObu9xzUiV+HxwMT4yKUH+74s
WMGxZRg1Z6xm4kXA02MpdYVWc5RxYXsCOvDlexIAol9uzhCnU+jK77jLwMo3AvXi
lA8A2lHnt31QhVezJLnUIZ6FjqMK3Mm2/glWp52s/gA78+iSQ+sN6+GS/1NLMHf4
QAKMZuiNS+4k1otosGf5wlmA4+YYlgC2eEZuZviIxTf2oB+ojfSPFEE63zC6O32k
h26tSgVn6FkbhoP1CTtt5vgNvm5pkHZFwE3amIkupoN9R1+/rLhv8t6mJf/+r/A/
jZCqgf0YhggdunRxmBZyu2u/tYpU5Mf10gZHePEWIcb6xMLx0SqPBZM+saSKfBkM
XnuKBcZr4kGQkhpXd4kGdM82VuqPdxMEkvGBrSzRM/tiZIqhq5sCvFa0uHK8l/Z8
DX6k09ovc8bqF2SHnWmvOa1pKtkG6aKUdCH5m4ZKaJFkZYoFdsVIXOzx8ls/dC+o
jbmLsW7T4/HxqaeqYjwzGk4kTTKGYIUO28a7gytpRjCLZ7HHrjS1hrNTN3cTVsxR
Dec7zcDd2eNs/avvRKti1jro+WlQiKZrxpMr1YZIXvDDZmTAdYu2Vn/by4WWhz2B
hun1KZ+TOjW/J6yqu+qrV5f7nkmMEB0Obg6PAsXYRdY9Hqe9+eiYJ2P4y03WMZEl
2Be8aYl7utdq4z/wP+Ju7LLJGaVhXY06pqpVj3KVg8ZhIGGG7YhiCAT8QwkVCbMR
vfF5fR+KUzGczaSeRZq2klaa7qydPYJFjVCN4375+P6Cq3t5CCKpBvHLdEP8ifND
u0w3uXsC7eQLlw+J3KAOQoejT5nQfYuXsWLyaHUfgHrD+XShmjC/XFduP7AxejlM
w5M+E88coxabKHFqI+GMB2fbCWlCeT8AVbUiO2UvXwHuoCpXwK9qQUmurqh6PA2h
+WkgKkXAP0FAf1c6wDh5+penZ28MtsSbEObvY1HRa8sdbS4xbtgZ2fwq2OQAQiI5
sYL54wPBTSdbGOhejd3vNk8UWZVqJPnxFi2LrBVvdBV98NMssFcTwB+VxOkIexwU
cj11FQacFkFNHr3W4QbaThihplxtSz3VUlqInvFOUe3+DMjcLJ5ZpV9TQs+/YVmL
lAZ9gxD0VbYLvS2z/zrFO/WsS8hV3UGvsBYRYpNFt1fWu8NNEXtcBEXNmIAtSpIH
IaSRxDkjwWOAjt4ozOihsSKqA/RF0ulhtZfOg6lXAOKJhe031UkJbTd2LoKJRc8f
fFzQ18z6sQ52oKbW6hRSBG2UCuQ7jP3P7m0nNPEsM3jk1OeI0CSfPik9d58SlysE
qOhRtX1YRlihFI1sWsea8TC6IYt7TdysBOJJpZlXeNoZzRVnvo+KMGUcmMkSb1XH
n6SDqKsSuhcR4ar/sEUkAhhPgugEvXR/hrG6sB3nkaAMThnedGnZtl487npr0uPp
Q6r3W+QKbVf7W30eAkTlW7C+uCzK8G9j4FIRwcbgGFdB6ly1wHYPU89FI1h7N9WJ
fQAvjHKYOXwjoFsfoIgFrJPRtCQlm/abJ5438CNOBPVQssqq5EePq2WpIxWPsB2K
bqpLijCLAFj5I5KDEuYsi4IK99Lh2+ZUdD+HMbWJb/8IlFxYAfygf34R6C84jnZg
jMdJzRFYOb+HsK+Bg0mz5ahamzYyppkmdEQYlgy9XI/NKhaBEeBh1A3VkoDpdt0R
zFLdCZpVUo5naDT/P+sCmb9hFhCUGmevNLTm/3gvmDX7CDFpop30RLXLRjTAmlxS
USzuw0v+No0QeuQ9eHDbWxmhbARwLUXiG0HyYeFRYOIiizqvxDDuXsM9SYch17gV
Mi2uizPejXokkgI85QqooQZmk5xoiu24/43bxlcK/VkGtMmBIM5YJvKAM5hdxHzB
3ge/DVoGhV6zHm3WPrUJmUUEXKkqfZD2xDy0PhiEKLdl52KCtrFRsI8bgaHLPeJd
0tdIli+/UIEmM5Vka1O9XiEV17A1JFVB1eRGUTFX9be3L8I8+LIpMY0z+XypOdfA
bYbWtUGRFirOqPCHNd45eJ96KcDhpNiVRp4LQnyy9F3s58vfMw+123DYMUaUW+Ku
jGZ5f2t52AVkaVTcuFgk+sgSY+fam4nXsKFAUrbFOiAOKytTckw8ekCAOvRm9744
T3zVjIRqHdPHYPJ/lbompMYHnLUC+gYkO1+c77mgd2eOvoEuBaWpIZwaHj+XLddJ
Dz/IeImGdCkkex50X3hwSHfYAatiK7kw04Q0gL3nRWguknJc8d0HKV3W+I7OFPKT
CC+Z9VGAaBdtXQW7GyKhY/fbUmKmsK2n1E2xOvWUOgPpODZ2UH8xec1RCrRhlqm+
cSfRjlO+B7q/koahMfIxevxpwJq7BoomiyLof4NU4o96BShmYK/sYqqrkaIOIy1n
+aWfATxwZiSNEuOhq6Ep8ZZ0/5iVXZg+AGXinR9zp4vRBHGE9GAI1c5WhAwyOt5N
jSrydx58BowLftnj20kmDg2azYIBJDKVl3nuDPPGy+ZkVBUZVnbYmUggmFYf2adn
xjHfJuE2H8skmLQyAnUPSHZz2/fJp04EivKZHz9i9ZTtnV9akrRJ4Thn2AVU38KE
jO8cqtmLWhkRoJphmJb8riI7u1d+1TUiePoN/qPVfsgiGVP7r1oWipUc5hV1bc4L
nJ5xozr+kT5K9RJkMm7ql2Z0dlW+B/BKh0HvK+BgjdFdOkJ3t9Serk4C0flLQ1u7
G12gEyDiVQMu8GPGCxTF5XTTTWs+UJpiWFzXZInjpqeH/H5I/ZCV7sUHIxG8vpXQ
dOTHeUoHvXJzfxF/pIp6CUIEKYOQIISWdEboM9rvLeaURQPPkjcf5GFtT/PEl2Lt
b6KVrxFXP481UdWrcn2uioZkrAhv0dcn/kpUQ4mA+nXh+//WeYLGth4Wsvhcyt9e
aCI2u/jWAZPyZ9QEmnybhYj2pjV2Ff9kWY5DQ5FiCFyhGjVgZM8l/D1b9yjrSiWe
+ylOuNfRdodZG9lJixcxaxP78PI+680ubg2pdykH9xTtrRSYqAeRUPiXl327xcNa
a/SOjHe41/qhUSbXsyqzcmEwlXgQENdme6kciTRn/5FlKZKalLzboz2OTvX1TdO5
muwd7WdHScehyV/SzMbk9jOb0ShpT+3Yt6H05ys81YI7N+75aPQylnjWolciKZ6D
7Ue9ipY9ckKciTyWNo2GcadmasTmbLvqKqs6XYuoMMgvGsdg68GzBbVREbL4HoXM
cTQuU9kfwuULdYAkL/mQoWPjD+/xJBMHSsAEiPhX7vbdMj1yk9RXxsdED7WHaT5F
HFPHv+L5HyWV52nGKQpW44J0bqSnjxUensbI/hIEC7xTyn//QBDNuf3PA2yWl77D
sguIYSx7ISspRF+Hz8p40uRAN022uotu1Tq9lmqaS/lP/GPiUnlUowOugfsV0S3V
/jhjT6ITncETEKEvkE7Oi7zrNihedf7BPj0DHC56Ud9an/R8AiQ/OqmEWp2FolRt
MlUoK/uDpPQF99o++5sHZe2N3HmhH24QOA6x6QTVZviNM4tMAlT7JwOAQ26COQon
pQdnMEapWxfO0XqEdRXh8CKy/fpJolIgpVJ11SNQKJe9ID6NtqmV41U6tSMLn5Fy
4B5AYxkBP4d4FdVq/Xvm/Vubc6xDIeSoU/bBK493LbG692Aiqc+ze39vve2Z4wR/
A25ZRIluljmUg+iofQoHbmBfr687sUCOvHiXQdr1R3eHKmE29D6vCG3jpsRumXDu
wsWzh10fsW/+iQmlZlxvaBcb38tH9f6YooLTEPUtMAi7phx3JD1HI8l/hseBJspI
yWY96sjixgWK9lBHhj2ftBtUuU7YaelLxO3+pKT5rzhvvx3SZmbtkpVAjxIg9l7v
pRO7NlikBul95Efq4xJTRTgri1l+D4c3V5KEW26MGZfUoiTwZ2sShzSY4wX7+3W5
L2VXPstwc/wGTQL0xhgMeu8kP1ffIi6S3mAIWlrwFv4S/Uexy7s5C9BVEuYfAK7H
p9IZq3YnruHb+KwzdLfJ+heA2KmlWrDeHuNZIv7OJH0UUNQbURXEUIDr6UgUBbun
NuQvYOSD7e87/6hKujcRI94UenWmaTbHbcWGPcfz7SVthkyGXPrn5DXh0HW69xRe
igjXIpPGr7AiBNxbs/U8cT4d8SD7UvJg0L99lR07qY9M6KfJcPPxQ47tNAMAdsQo
nrixtXDloXQ3IRZSZk+0zM7ZHRHdjGptyhWuyu9gnaxUVxvw2n8+dYDe6qF+wa6L
AwdIJ3vs9kXH/KFw1bO/cjQifpuiwReB6/1+hPC5rdYEe+Yk9IGmAlSsMHMd56UT
ekjfsKdMweaT/3fdE25UanVylR9DE15e0bmyLOV8cZf5+nrGCElicca2tWCgn1vg
xwi+YbrV08L7DbRO672LhyAkqSuZbamg+ibddZ1htkJLMasRSxk29OeEi5AHWY9b
wKU8jphTZV7Ensftsgz6WZb/G9RnPfDfTpfwc/QrVikKUrKQ/uiztKBfNFmWoKF7
pPk8Zxyjm+HOwy9ZsmWPAxrQY3QwiAsZH27C2Wt2HC5ADGuLlrUjfYSvTxRFtBWE
ZmyO2IlwBcKJoNmxXPfKj1erPAFG5ljgip0HD96GdWsy+rrGRn0Ga8yllDDhPMGQ
UfpTfxWt+nKs8O1LgSE9H9BwtofP/NAh/HqpsS7LeLWDzmYnvCmQH3vLlntw1MPR
fkaGvEKlQSfFdr/rKDxdjWmwyqMxzSNSnXMbVk0GywdR5hVj2ts7lXl66sJNWdFf
2Fh/A+5w5RO9EgrWWN2uEqw2ews97g8n08gjHXviMf5ooB6/+8xGgKPUvFHjyjHT
Uhb3LBtBLQ15B7eq9/xF68ltXzq6cfTiwQGrz/WRoZj/8oUFHzUq+AD2jnLCamue
JnlUNUIwmfUVy6XRp86lce0HQBuM+e81i5un/6pajIOh/ptX7AWO2lCGTwXz8SpF
ydeQIzQ2WZxnHRgxZk6ETlRp/ntIhDKG7HnQXfw7+xbzobFg+JrUqVa4oy1/tLki
LkquEp5ZFalzZAI7cb/enofqvbUBCGh+Lz/wqeF4qJGu/5SL2HPh4NDK2LJkSUjW
0ra5VgaVxdCZXT7n+OBMm1iZmwfNBOUMp/+T/YmuSIj6prte+xhjr6a9he2G7NHN
YMTvJzjMyQJjCClkwPeyxji542RUrjqv0HNNvohkcCezhlUGn3UcRxZYeHF4iADo
VIrKmRgF4wzwH7E70Ux3UQVeepLvKw1tMSWn6EVfFPYNPTFOCMJ8aYfRGKTQ3T2w
eRg+jWTAE9B2IY5PEyyh2TQZdABYasvejTAENaHT/A+F/WO20P1dYl/Tnx2iVTaV
VgoR2fYEil4f2OPBLZ2NDLTaNYNALnTog2f0Fz2op1H/ZKqg2Vpd4HanGOgEnvbL
fxOj9g1Nci2BfR+lU7JcP5/518HmRIz1ccxGwB7ea6ffsIt8aKnDd5LpK0ipSSQi
k0SO9zTQaKcC9OMqxxdPN4WjsM30onVzNGy76SzJAd2HacYBV5MT2AkiFNUKWNnZ
BL+wTVT7SgEaWRwyEFuG2JCMwMAghcxnqOspTid9wHyLdyRyiE+6GPms2TShDt62
IFSjb5X9rn2Tj2o/+Tjn7hAz4t8mC2v4wDRPqIDDgKDggPc5a0mSeZa8cz9S8O4H
qIwadjbpl5wfRlgeUZ2ylF/AUPQ43zLDsKkTawM7gQ5smq5D+nR665VTqRxv7T6t
TzNmd9O/Fi+1rq0h5P4n9D/o5Dq+P5gwdDNQysQ0KE1EtLkCJp24R0XV2T8SMocY
7plJIRXWXV5FmrrznJk9Mbw1EaXtKxIQzLo7JLSaQmFnmCFXpJ20LmHXfSUafXWb
KIS8ZQKP+bAmQi4oIUOw5WSsPjCTCn78F0DMpyh71MbRDGCCDkLEQc6LPzVfxY4X
/lw+4MGFVCbHMrLGj5bdOz8U8c9tfXLZYjLR5/TtomG1qMBuicckpdsZIi3C0MUB
zdR/CwFNnvTcV9+V+ggj6hdMU/so0wu76GJrSF1lF01El2Uspmn5GCvA7BevwUEQ
4GvRbQK/oANOTf6jT7wjqtBdwu6MILpA/JlADfd24MAokO/IIOJQcjJzPDzBib+q
pc6ATXC19X0Mpcatv3B5/Exr9BsW29v1MmobYDiDj5jmzhbqBQXxKdrfzmJKek2Q
tAZpHS9kTLKsJOjyZM5VD76925s15zMRuAHGzg8IMaubi/HMk1uc405vlpmyVPb6
qZyeC/4NjKJYLBNfw3+E7E2L0rH78BSvUfJv9foeb/GDlKblIdDpX6ecwV9ZRp8p
PL+O8xFhj6xByjYl0ukXTnz2y+uiNpaeetcRc3m6+l0Mz5zbbjerrRXLgVVpPBNs
0CoS6/tObv3cNhbTwLnOeY3uUOPz7f4rUnZR/FLbiJbE6SOGlcjh4v+1uIPuvPNt
on/ifHfvR5WM+J/DaiVAEbx0uPSxGAjjPQOlRi2J1UQZ/VWR9n7xF3l/7DyUwVH8
Vi0rPaAVcG7YK/Efpkoz9omIW7sPAtaOgvFJH3IbYOp/XSfeujnIwaTc5QSkYIu/
a2OsgGSqjEA8JauLfmyR8M9ea705nsJaAL5zvgLTJY0/lRfSjziBlVuhbAL5AXZP
rBSxTjOVf5wZjjOF4HdFkG7atLQBQUYtbKb1Udh5PEnztSrYN+noy5eGTILb3ZwA
Dg8ghh5wmNr7ngwV15Lki/Wv6eKxuR38wrKVFfGUJPijta7fvYMiE3I1wBNNAISd
br/HuEOP5v3HSrlKLeJHUUG6tHrkLHu7j8Xh2y4LA9pqZm9C8YVvjcheNVs52Lz1
/zeoh9KQF9bGauF6aWIRbGMJ4TrRkquLpnBPsNV6qjlE/UPR/ZribjDNls3Vvuyk
O97ge/85VQ6CZwZqvdPAHpGEZ8ZAJ83z7gvsFCGpbXdf0fjxqqUNSic7nxwOGLNh
HZhvhn8Y9Ayt18QdgH1kT+tdY4Akhl26Ulso52FyLGs4Ebwh1101nIJpvNXROj0S
TT4jS0+xg5fXB6PEdPNflA545C84fR5mLL89ep5Fzu67IigvYIjv+Xe1b4DL4Htz
pKwBtRlALK/iCdDO5Ketk8Ly7GiNS9AGhyGKHm0PMC9Em1eZFVPRxqR2oZilcJMe
HTVO5GNI8ii9KxwTXbd9bktNb1yjXwj9fnLY+HX6h8fI1wUA6xgqNeM9xOhH/PRe
OQN7dzAlYO+m7q4Dipts7oVgIxVBZvVuO5U5ZdkrRclJG5Sz73bf4Dfk+EYC+c5j
vU0eyR17DDKzNXFacz0M1fwOvA3XIbsFl9AnTVXjIKuAfKsCBfGfNITvSL85kmtQ
5ew2d4iplOUnXXaXH5Q0qssyc89bbsr0O2g2DX24zaHkYFmt8D0mkfyn2LyckYr2
/eoO5R6mdgqdLHMvqhFsoL7EblG3NRNpgNzMEgCeDOlAhWT0+5xKW9cRtP8H3UsN
r5LSSIeKAjVey+HEMRUXJh6Wwdx5zZ8datbSrhBK8TM1nZWabTjZ72JkEg0157Af
UvxXhzAT8b+nU3fG/xhtv7g6IbBm0m/wjh3nsoeU2F+3qcPYBAkKHBoyyRxv9q87
05Xv69Mceg5QbWzHP3xqlnwV9JNBgoTywJAhU/gL/Qh0MULt2/Uw0mb7UxxHjIYN
jvahLJYG3+BcMC8Xde9MpBlqvxP7o+UlBa8DMz1jw0tPX+ZKVeYmfDUXkPGxX3fD
NZK8U/ApjpwA70l8YhrSxi9tFNvQKBlin5tK9Sk7m8wHQZeSBRnF6hJr+HfwcLxR
WNiUkF9MndsHCqnLDiKWEooLYAWxKI2orYSxqUibke7m63Z5iUiQPT4BqYNvboY9
UI7Kkonxo50wwAqa2mFjZnXzYQXrUFZ9NyWgqqQu2btB0tWKly0eZDt9BzMlZo4F
40+jk5BgKjtGHUWv0v5WcOzn4z0aFQ3txUGrd6xm4pQDh92IbBl+fmeHU2DXO7nH
EkgHcyDKxmZrO9Eyf3+UUNIdNrTF/CpLPh7SZvG0ATj1MYmPJa7amcuIL1Rp/73C
0n9uG12fUZdhnbuWkxf7ZawVeOf/FRHZ4/imViy1859PcU9UVnTXt/Q15bN8uwZ4
6bVFsLDHMsBgv/oZePR1RhQwhRWJwkFOzsPhEnRWE6XbCc5fTvO1zC7OtNvyr04+
GTlV7lHUsRpARoQaK+84W/16zlLu7lFDELuofZMwq8W8iVT2MMDn+NBPEu9kFS3L
6ng/vSlKqhcxKoHt8jF9mPmcrGTtLaL71bNEY6wlMIzM1inlNL/J56xidyW5fJTr
QNcw+RBE87Tn2SUahqsYfk6byifxKX27rLAKjeVd+yULUKdtCZ/is7qVt4Y3bUfc
rt7R6lGC5K77o5XPXGX/XsHnBWZ9NhPghf6LB8W73cFlaeowa1WXnmeTV634KtWC
itTuzZUQLEG92Eiwe5hSZnUF+ZzByqfzxkVZFg2kYsVh2lOS1nd1PYxRmEFxjY7P
xUXGwe46CThtmB6LyA/oMyeYsx93ZwVMDI9LjgZff1QUIVphM69lVQe6OeGTFi7D
J7szyIC7qsAg0yERZYNGzL8wQyOIKpdEIYecUcS1B/PNon9G/QDDICkszyuEmJLY
8rxMSPDJJHJK7dJq3MDDnPPm3vUyKlcBXJZBYK9MNfE4EnCjsiUmSuXIYQtX04gN
/NTRjpukr6FmuBXXqhdvCs3LqL5cT8T6idvK+bcCv8SpWR5Q6bwbl8aw+0EFsv3+
nSnrCQ5aSi3IEBOePnUldpTzJtnJfxagHqQDv5vFEV9JpHHCIAZgQ0nPdN+WbPtJ
fQkA5Zd6sZI0bGluDNbz25GOj0J0IquxxuUaMx2Swyib1bBCNBrSegDsUJTBzUMm
knKjFD+4cz1uAAQkoTc2Mvb1Hwbx5Uu4VcrbCsTPZS1kt0Jjz1EJukrMWA0el6bp
JwiSGUmycUin4iLtiQSkP5no9xQN/ret/dcAVmaTpiYD/4QgSz+5YubjLkD/n1MC
p6YQv0BDRgGL6OVOPEQ3eaBpMDa0RkFO7x5x7JRTrr1YGxeg58LM6P2VfJXKXsWZ
v+s6dQtQqGWOeHE2LHWUtpMFTwoFleH0cnFzBHBmTSVoj9i0sosKVCKYjMhWCV/V
63QWkttl0LuPjEI8RABeT+qJ4YdV3j1hizh7L5/qUAlZsy3VA/QAUIS7mCz25KA4
HjkRTo9cNPAKqaEvKLwSyjPQxAtGrRziHd3Ge107pYOkVQGLxCKeaqB3z5Dn8lGe
u4KEA6gNdboBWjJVqAmNhYNM0pHVaYxh0P43iSDUNnLoEj7kUArN4F3rnzWQuQPO
iVbvx6Vb8sw4/cetZHqRJwDxf1Odlloj67Pcgo34nwUfH3ObOIirk+iIWQMdEldP
aVjx3salukKoVZ1qsbOUYdnuqWXjqx/hK7q8i/hawRISBfszMKCk2XEGn4wuAqMR
kJAIUCbF1IGMq18c9uAd9XeApY6a5WY4697NC0GnYxWG+U3OFEcGgnbjx06BFtoW
HTYI4DESvFRfyxc/PJO32S/tUJxYoSmBxOxRSsuf4cUeKNZmJmrlpQd6vCqC5M/h
NQoDNMHfCu6wRW6Bv62pJur8c92eEJPqRZLX2NlLfZx3PZDkz9NftVx4n/Vf7ZRg
fG77WbCyMFIVveWuir6tfvHbsetb1kwg9Ohdbb5qZeu/70jS6FozS6bVekAb/tMN
07JecJQiOt3vlR+5T/WiWMRmyP6QViIRUfEzlng5dyEqE7g3gDvupcyYGR6C6u6k
FogGOUhQ7g93qZvbkf1G1M7ThW32wK3XLxjigVuwa76TWdWR7szr9efixLKVr+fm
v4S34nzg4HFV5lvavwuqOjLXNcKG+sXcVdQiKm4QAhydE3KaeB2oZUsBlC0p2zcv
hOhrbj/Ap/AUS8cOkuBVCTvPwEB4lkOcr/HcNJgdISdDN7CTeS+F+Nygj8WR+FsF
hxfCtvkJ/bsC7x0yWkxhAx2TOc2OkLLzcDqWGMyidaLIrrncrvyx+Grl6kdosc8S
Tt/qO7VCUl4q+mTP3+YY6Rf9ymqxiGBka2vywH/6eTGdI8sNofbszI+p/wtHydOp
21onHOWnuWLuACdG5QLcrNXiQ+d6vQO0w6DzTcuMI2wYRonCBktjgmy5gqqcYXDr
koi1cRQPx6eHS7POYd3VLzl8oxP5ZkdZGsXIvqerZywCaSKzrEI/o9W/oDMp6eQf
oj+Az5CO0ThBtuG0ofdqkUoCE+5ofIOH0aqjFoYFlsK39ZOHUq7HshiiiRuy+icb
gUSihGNVbr9Y96hC940G349teE77X3IY5HplBHmiOaUXjlA1ycV/1Oa45R0pw4ni
QuLftYXrZwFmrbKmpH+C0cAf3imKI+u+HwMdcdNCKFtTNkTcYm5VMc5ZNULvCrKS
B5dKimuhFHBG8+KoJKk5aOxhUmxXaCtm4WMEWLRmM1X37jdgR1IgN31aPtMcbz15
WGeaShWdoQIdUgDpRyJ8Yrm/4ujOsXUMeatPGtKR1WdbEheuaPB8vBIjo5xal02d
JE1JSR+aAMKdutDQP6Jt4xUpocnojqDnrEUF1tY091JBelOEZ+fvBG/TKb/vmBHv
GJgfTukwrJO+e+dsLr2lGLmWVQ0M8NRJlTUY2sO82/JVjQTSWK4wQGTQD6l2PxZH
9hHEWujr+af92TIfPbn/hNTqMWxw7QaNrfzLkGvDHDXboS3Kfjla75tNgN7Amxf4
pqtskFY4a4qdCRyMu81e9feCdLpvuDM8GhhZDLpG3zS3koXYY8UvMQs9xGbObaGr
Zfyk5HwsaWuOGgZlCyzlRxCu8k20L6HdihvXNcvmHh2C/dM+BET3iwktuq1Hz9Wu
AjsgI77tparGfcTQ2DWoj3B1vvokwQ2b8feDYcQLKerEZ9GHc61P+dIQa4LBXkHB
ISP/2OcUjS8t9sCnbrn8UwbWNf5ZjOKqMYZRn6DW7xe9DfYDtS2ejawdCrTPhaM4
P1zOR9txUfBadFoDAd8Unr/jPbsHdHL7VoPMDpfua3CYTPrlMYygkZoriWPVfXaN
CiCb7ThVhY0pA/F/hMv9ZKyv7C0XMwdzyfzhA0pVUDE8QZh2QQC0w/wjyCZ7V4l3
oWPjcUyPb9jV4hbTV5qqjoD6m5tWin++kPIBTD3/2byTrvZEOnONzffZuyr+wXdd
uIbcv3L+Xy+mm82qQ4Neapk+VrGSLOnHGacWRcV5vW4wOrc1EM2hZNwehLT+Lszv
l3/RdyzB5Y5U957ntRleXK1CnvXM21RZTw/kgZEx4LOr0p8mJVpiZ6sHGsGLLywf
+NnWH707FqQa8iXyiFcJ5p5P8CjZogiWQxAUq9hN7leCDNbVgrpboKdE8u+vdTdl
w5c4nE6mKXaslV//cVNr/3GZNFSTJ9kasuHl+0dDPnAJljk0KoykCzhny65B4Nq+
qKyejiL7Ti8AIW2IfcMeurfUPw38GGAdPmafgxi0w9iEuHKHgzL9F9HMJ3iLhm1c
vUDQnx3bj4mTb72zjxnTLaCgo1YUAPBl3AZZqIQ6QOUgLJfMm2k/VB9Nx6/7MKXy
OGPq9PzUa8pcs6r09MsB3BMlLYcedqZXiv0JxC/lgGZKuQitNmRjPi0BBWUiVZiw
oIRY5twxFVhkQ+BtdPqaErFN2Clbgm7DaYlBKwpAspa7VsjMc+LfBhdO9EMCDRIg
P6bnNEiRvII+P0q+fFNDHrjl/AUPlgUksNYBwWquXQCsYoXRqBr6a+yOZsU4sYW7
XFoZaq+HIUhHPGfc6qS3BVCDLLuGj5r7IttzFNCqoewFK7oHNCoLr8jcZS4fJtTj
Wre+MEUJHNrzkXKMTlIB+CSxWZFvICdecYQpG/BukjCpVAVgO1L96IvhMLN+8rfX
KCKF3AaMCtxqJYG9DZOD7l4iUakeBWKHpByaomsuMUZXrNqQ2nDdQFTucYGrXwt0
YnM03MjDFhqzYkgkXUF5A+iGZ1Grwsrvk30yftZhpgiDXksCBQ/DcOeNW3ONwZOV
20Bm9Yym2PP4Hvm8muaL19g5JOL0tHM28QKy0ftPH8VC1Kyim1ywqdYW8HyPMBDM
zJXHilwG+P5JISZ1KxkPY9QsNzRXyaQ45uqDTs/N9RYVRWPWuWEvc3yPlSGoxyMX
UBDeHs0WhPg8jlx1El1FNQxncUdnjNVfIAtUrIFSMUGLzijH6qmKyj7phHiOUbBX
NGafMb4qOCmT9UNnFCPXbvoiQzMSi3QzudI4v34RjnbTs7Kh/5ScWtXpvLii0ILQ
BqxhiCFKBFGH8w304sMOJR47z5YCO+JmhMvyS5jzFG7fwlIBVI8SAeGxVlDZk/BO
Zt1uS31uMkwxsx7pA9G3xsV7v5RiTlKpsjZ3pGPnG1p26Qkh+pFfWi73NReRNyTg
m/YTj1EFpBNC7z6WFt9Pq3Na9gTYtqf6T4wEQATUnR8h2FEVarzE/qv4TMDseRAm
ttuoKXOngI4EQBC2zZx+wNH/t6qXW/eJ0Q1FG74jlpf0+Y9RYpoi+uQpNTDl1bYX
Kkx0B5v2UVjPmLCK9G82vzQwYxPstye8v2W6CUv9HRXUkhAZfd+uq5t0rW7OKFbg
AejdmFPfeepIdMmRVkrtGK29Bk3PGlHlRxwpuR2fn5IHLkc8Aw0anr+dcGh3j31h
YulaabEvbqePeKcBkLUB5rfhsKJl0xZr5yxzyXgoDy+KQPPZe/42+ZZ8LBNzu5mw
9PzKGaO2oT6wHavBaPNqOdOzr3dMhmV2P2rBJpqfuWxHETxooMRjEbz89FsEm2rD
wUMzuHk9hdye7Dan3BuRDRWGztcW/aw1qDRNnnIk1XUNYnytTUCBn2LBva78T9kC
VuFdsGSMYRSn9BKizve3Fro5XxkPGw5sy+0iLOHH3JusmyxMOV75tVjDTLVleUF+
LUOH4rurBWMHkSX8YOV82VIr1IFFtzVkP3KcuT5Ga7iVPZUKc3gFhlpMRrF+cMv0
SnD3BeH1HejbZcGc9JwLmP5NQ8wVP7ROk+HvbkJKbu9L31xSACs96ZxZuqlicvQc
awHT2OOqKmx5wSD3Yg7ymxk6xBZDweJJSDdnOxwHHN5k4x3xu9Tcq6+8A1HXtmMt
z8LtLjzHBC0dtWIbDJfyaLyzbDXdSouXK5iprC7AckacsmmMI+gApDXjc5otP3FN
sqm8N0GsHRwd6u4PsZg45WegU9141MvYCPViEQ5IrNWmT22jk+dR+6l4y/D7CYV1
cO/6IuZkfmTakEwMeJuT4OBaednMvUkskalVxdBWXRMZAo+cDJsQ9pPg1DXMOwL6
JmT71ywV6JRFflgMf3QXXqQx9KidzQqGeGWRyjDQrP5eXHgCEf6fHs7M6V5kyHko
BdpQLWDpCakP9UzfQiFOkhgK1LvlbcZf4GEoTyUFkjzEcf+xutwxxjEC8Ljn/Ti6
PnqiRQ7Y3a3ygxVgCmpcHOlmagtCuR5RMrpXjJvywfkepFLKU6B4vxCE1fnZy5Fd
20udNTptGxVTcD0xxd4j6NDqrDFqdLZN+hhpgvfRLAyj6MnHSpfYUjM49lltxIAT
ToFMnFzKb955aPXktEgfMLmIxQegWLXTY5Q0FMblFF/w3AIJ+lh6IypVUtLGFRcN
uAdYFNDZpAtav9ViLmOGl4dSf7Sd1BNJ4i8bOJV57cF7vZ8DtrYb4FrVVs99nzR8
WoMRWZg2J1JFvm62EevWDJmNDjjBWaS6QVg8Mgcv8YQloHmY83QCJJTmw163XBFq
82hAjyG7SbV6v7OnpX880UCMc+OzfgquOo/lbrwpiiM1TyrTFooVtqgL9imhfAfl
efK/8jXdQ9XUbTyLliFwu01QNzBoHdaAdePSejvxbjUxTR0Yd3l/35HQtcf0zXEw
jAKRG+WEpzEGlCH89paQes2evVaV30eaHWZXhDsFAZZ5cwVaZLRvOvgYNnnH8X97
grooVuHP58LJfLDqcOERL33bEVrsq20oQiv0TEY2JSMKHVS++uGD7fbxlWQ8Ml70
c7joaZnAznliDvSLzMeXF8Q0Xz+J7gzSsJ9+IsRSqT62f7CE3HsgTuNPiSpE/G/w
izvM9QzgeDGq7Ni/tRWoaVmKBT0HyVeVLtjC/+HTbNe098uf8RlJ/Fx6AGL9+DHG
CAA0f0B17tTzJQCz/Aigi3cWk4MCsXZ1jmhUJUOECIAitH0Xs1YLbGpYaPr4OoO7
deQ2+xePgp9LOnFC6d9yqMZAQmsyNe9Kktt10nfT7tMNHsdOcsdmkARUv23qPEjU
hXsp0hCTkMfgZVAhvlnBL6yLLCjpyK4riqF1BYphVciqpECaqeW8ZrLeQkOQVNBd
/JDL2txUztdh3YV9Zn5F28Xeu6XAbI4OiPa1IX6U6jqe3d5aPfbzmHwqqIZHVTrP
dmSfYUub3tP4kfbQ8/oF0eK9+W3jC8wMJxPiu6bInz2WbUgcBjod0wjJyFTDVlCo
fwcddNNfETg/pLdZ4KOYgpTEKSoDxUa2AkQCzDymG+Q80XdReanRm/4ahCdabaC7
lKzmex2L0sUYwQlMLUjHw+1uZOYQJany+O35g2LQVMaa8RGY+g8o36soUdWeQInw
mfHTQpo9opBvEYbwZPMkAMdDkcoxyNO9Kc1PL5C2NQTqTioH/QShlI24un1fIVBf
s2JTEuIK4RAlwB8JMyuaRV+Y/cs/f0GhljTm4yTUkyawY05b1wfE+3+QkdMRxdaS
J1PKvAelLpO1MuAkWGkIL9Ffd2BlMAxqoCTfzFD8su6iFb7rlIOL4x9mv+5FVWEd
i/sBaoOjYd4pHDFteG02yWxBd33M9CTycqXG9X4Cgv+UfNHkpKjnZlopYTz4HQbZ
hsS6RSNHtU5devujW4v1UIHKyQSuW0SzGcVPSFA+m2nI/sbhTa4u1M7qu+4Y7RX7
LAUFtxgGJ32RwwScRMV0Iv8kvvWSRE6IL2+pNdvYLH/kfnyjiGc/NurlMnYvN8FR
SYYCGHZFUjhxo1CwZnQUwy5khX5z/HZ7ViXTSfg7pm0+lTliHz1VaVz3Gr2N+Pgt
HpFFU5GJvtvnNxtps/yReq8UFkCqJEYj3KKAZSQbEGbBBN5Rlfdd4yHXAG2RjYx8
d75lHDWrUl38XPAL9/+vFJSfNZWqhUqv1xKE0DvKNG+vWGugoX0gAHFcVPxXxAxQ
7reSq6A6u70X0nDzvF3tYvM2TC0tJA66Xvlmmam/PX1r01CYB7gC+gbzl8f9Pcu9
n+uwqooL2D5HHvPcVHT6G5tvSSFrbPY/VKXYZNCuiCczQl3V4c+RHmUtqXSjdkwQ
1AQNBL9QjAQeQ1U1NIofmvSOBK6ijN2oDz7z2P6TowgKjdffzQ/b3K+a8dvZ7zAm
XSBV3/thjXPz0tjbAlVCMRiKq02zl6tcIeEAxxAxN9EMYEkdbv/oUUhGkNYg7X/Q
ht+cpizco7VadM5HsEonziX28taMpQwA/2wBRSX3o0gh2hdjMe7r/NUmREa89iuK
nZQD2e7WeRMulOSBBaWZGQZS58OpqqRwBmuLNooAQwTeOVAJlV6B0Rfvq30j3LlJ
j4GjQcy+l3uidl8mHla9uLdv0PlV/E0UF2BS2qbNCv7VqY8TTILuaNsmC7xGGT5x
8BmyxiN4UlIbz9qhHYPqCT+6Kel9/+6SxK16qyj+GI7eqVWzxKvQuZCTw8U7IIm5
jidcrGuboeUvkIhEelXeVlrBt/R+DYWCn3uAO8shxNa2ZXN9WnSQv/zwKFIp3d/C
mVxJJZhXG08f979YfF+0l3Vhw48QbG/51BBRrSCHkbvKTJDoSzBB+RrzaQIrvDLc
hzZIaexu685gVM8d3YqxLKa8bV24SRzp6DBmxOYagaohRsKvHA4uxewmDtfDGlVJ
iM8M8dPlas+DfwtrJWfVTKOkSjqGgnMi/G5xdmZMEgonqdp44crQLLUwgeCEqYWs
r/wLPerknzEW/Qn2etdlbYitokheml4CxpDptNEcAjKYTeDm8/WR+S7BaV6Pco3Y
hEDoJJtI9UxrNO8Y5ZiNr/2hahe7mELSxB1nn1jW5Amd1/UlGGP7mCluWoRoPkgv
LhI68j8S64nSlNyzQxJcVMXEO5nLuIugCvqdJrfp8fGZeirxrW25VlqH6hwurUbe
iOxch1MTh0f0KiglAHwhJ0MCZnMFW1ED15iAuc4/PEqyUOhnteqkUwX9KML9JQch
5ztzsmDdhcdS66lTkZmNyM0MiT7PnWogTNDrbkX4znnbO2xt0oOhYeyNy+Gu01Bl
G4G4uMp4lc8wyYEsAlVFq4kspiLd4XPEg+wffYBdlxd1B/YMY1mx+xvpKEw2Z+/3
09+WCpmDznm8L8ustaQdQRoCZuuI+0d3Bq9U6qYORonlaGZx5Gza8BWg3DRA4oKV
SOCtWySYnNM3C79mewZ3DfqH7WLtOHRl00hFlQvqUhDtj3ctZbky9A28ZK0JEpRG
8TOJEXvr2Hysm7JKBcYMWmn6h4YTxMi9N+LKwmmo6orthIBGJLB1Q+aiehzMvP5Q
IX1sn1Yd+reJzEc28dQgLZ186h3aIpFOV8hia/xq3OPDFYRGQayUGRX3vaOFt5eJ
44GNuM7YNSj3/3Id2CjaO2Q68QSdX/UNYyOPhhzS8GG5G2W/YYm8HM42vdI6Xm2f
ZQx9py0oDo/XmE1hVD7gQxblVoSz7/soQQZhJdvRj5Xj6WkOKn8PE6VkCLvzlNeV
V3zK9kmdr8g+YE1ln6GGKz+xIUCepaB2DSLUJwuNTf10ZoSyZiKP2nZo+W2AqDps
DWgI+177RMQyO6ZMhZRyPLiaXUCypF3GlYYwj6ZsDrKYLb8UbGQGPx24yqeZFIUk
FxZq1Nk55JhKHxzCQ+QbYO9wHt4JloAvETHyDacDy6/uGm++oD6pxPJ3T60+NnAf
yVi11IaGFJ2dH9MRiASQlv33UeBohEcPgOi6Q9CAgZJFJEIFZgOueRoBMYjjK4Sy
AW6m2zBWJPwFIMvCy8GepiGU55hYGpPfy4B0a077QLoye38AMQ6sDnpTIsp8G5Dx
z9y8Ud9cOlsig69s9GUaE/4OGOf/2mN/5qprP82BXsGDX/yMi+kVCXqs5JiJhb8p
uanYv6B6ZhWKn7GW8Yje9Q3josefNQGHPkNg60aRWv53kaGY8WWi9Es2R96L+hhX
fJb0owHHP/dzxt0xj4a+THAxneQY/iU2z5W2azK/CeDJWlMDEQRyo1RUPB76dAze
p0yVNBnzs2D73szhPeEir/FiUPiBDFoJYMcHSVAgTCHE1dHp2MLZ3139Hsf3XmEa
pqAzPvxVAbQXL78lhLqO+h4V6qo8BwTOWxwIkBB5ZlXZD0Juq18Bfp2Fzf0xHNXA
LBLDSPJZtCiEe2yXgHupRhDIbjRV8FUa9rWueEWhEas26C7EA8w2dPehQY+2aU+m
XGOJyjvoGKgQUjUMfINSsomz5XicmfQ+d/HLHmSWErkl+PCEcGXFRp+8jNef2zwd
/ZEFbKyeWDY21QHTSo2JUu30rqpIZymE1is8DTuQpdnbISKp0BxOPXipj3Xq2vwQ
cJtRs22w7hcUqD5nKkfh9ooSLqRzTlPuoFQjQLqif8QUT/bMDlIAVD1wrpyuQ66t
X/hCcUs0d0TLRidaRVOZ7MqOzWRTTJ0aedWfNknDOCIt2y/HBkFiAGgI39Br1ach
q3HKbpgeM3Utiyj6fuYj9uH6bZMdSUZWoCtZX3wpFeeMKo29u9a9Djl/mmTWYb5G
7HdaTJQybGJouvMQjb6yLLxDEXhWCG21fGUm3b7D8H2iziGbzNYvkUXZHH1lOrbe
XPwVlbw4vLc/k7ZLo06orxBzvq2hseW88WBXN24OvGWi3DRpIcK7GvlcA+EnKK7F
Zjb1WyQYJIzABIYGg/3ufG93Lp6woVi4fyBuIIdzXYay+BCju0rQlmZilB2W9Z93
eURxV9J3FEtnd/zQj+ma61BrYHJirZeSZCJQ6GQ64/IZsnN7p9STsC/qq/wYe7mi
rM9z3kjOS9VzyQpjWEpgVKoXcwSPBviBFQMiM1crnajxUMNqbOa9pcOlBEvhZ56Z
Sw03216Q+gsZqnQUBguy2qe8vUqdYEBE5jY7EWm5bgtnR5p3/+r8qEix4aa2VJiE
S0GHYNpvH9rrPOzH0I85lDiPtUeWw8EKDSDzKJcfH+KjDosXwV/am132qz9dxXVQ
n1U1vwV++2lTF+abKGW6yKTaDePOuU/ada5M5mT1oJa1pgzt2ZjvWslQrr+dUSbW
hoSjK+JzEKVba91PFPbU1ISK59E6sRBbke4RLGzfR4B+RTDZByrFzZe3/ysE9epS
xg+yzXfo7en2I8VPY7PlaGscpPWgpM+B6UrdhEYQR4J8ay6gM1fJRdFfzbQSW8bM
VIAMCDuCypFjOKU9YHU2hAIz6Lao4HoMf1nYOAY1zBm7KdsTEafMqWgeDG7ida8t
rRR1zVAbiwwcOIoPGigGzlqrGBYorbLbHbY0eh/SbU6bxobKv3V5b+1/SXKuFkbJ
T/r3yrSt3Hny63CodJGHQWX15FPdiqX4IZoMDGyPuZKO3+N46EqvoSYpxRwTHAsS
69oyDspBb+0ORYcSzEDtjgmHDfUeRHN4U5TGzuvRn6hDyEsSpZ5Z0XFEP60yoQES
Z3GBMK0nfMs7Z56BKBDEtUj++gQq7i1gChWaEPtQTBsfXNGtoxdB5htMLTDKORW0
p1Qb0WuhalHevHb5Ppl46ysLPvJCYlQCMuQNC6KjfXjwqxUWPsN4rqhZXcICNZTT
h7Q1jZrem1+WTAzALzREuGwlCJJOqQrCUmZU/T+RcJVCdPLRvCzLOaPfMHeOYjzm
NXzkZjSMGx1MjidTE5m/1SH9SR53ppVLrsto2cQRuIYB45CrmY3JRmQMEUacKcnm
sC02p4tPEbNNL/sZemrGDwkH8WOI9EBN++LK8V0rhDZAGY5t8BjaSwrrqpsARz9t
Li6VG8ORDz5c2ql+TLve+Sma7qZpvay2vPxWtYpVIewv4HIfbvYA6iolPfDoVbTC
FUfBqyc3UtmcN/O5AGE1pQM5gvNOfnVGb83F92iZV4ZC2FEeCw2youIHMhDXRr9D
M0KcH4HVu5B4wHm/yGscfjuBak0bJXNP6hKi8VI1g7NBfsYPPFP3+N/ErENWbmel
Jc7Q9Ur7L5OaIzb49a6eBmrxN7PRvr7qelJTB813CLTA2JIoJgAy+7klNBixyhzt
g7qjk9+73G2h+ayk+jLiDA++fC9qyLLgRYMmHXW2Id/YBxP0aggh9vvRzssJe+54
GC8pPLv1dBkToeAJR9bGgosFYfb8hcHq8Bb+BESDZR1RdVotbPPUpq+kiw/SDQnT
Pu6W/BhjA+C1eD23AS8p82bI7r7sukBgPjnUdTqmv1n99h6qQYMGQyHDN2wTb2gY
BT1LMhXc0fUI+P59QhNlOoNdaByL+tNGFg3+SeeoiYao27BZ29uvf1tRLwOHTubS
jKa9bdL5gwLi1mZxAwv6Z+E0mR9ggjAUkYxOs34SjMNF7egImg9bJii5DVf7l20e
++oovtIalALkQEu8tWzpuZ/CnVWxVFCgPS7e3cXoU+9PbP9HMubvBeWhZNkxsJzN
OyijYF35yc6hA6yWtM6K1iV2FzrJj3HPZ5vPcXY18/+YNJv6RnU4y9xUE1yulcT6
Ei462MAkirUERTPFr2KmlVp4ZdVKYFTPGMBHdcE0trLk4l4DPjhxXq8WbikMHHus
tGYAAo76nHeiOugZ6fB0UxS3ks2S2N79iHf6teFkMipl6E9gJv9XTj7XRMtYd7oU
2h9hErxg48El16Bn1M0nr3o0wrBX7g9dvK0viahfKwCPoNQw/+p+5xeQe+2MCdq+
4x3LBKlPkao68JNJon5/JixTlaAb/iThYN8nLjsTcL5DCn0YxVK20iLD71KV+Fxx
X03DU0rYsbFaTil+7qItc17V/RDV804hclxzb4Ubrn4rGtA3MhXjtWJUgiiXemra
kjXxnGXTrK0D9eA8f/+It6j/rQ9HVqP7/e632WaYs0+NICSNG0i6fDSFzwbuYS9m
wpIcduhbzAUOQzMgIBfaz9z+PtGyhTwolU+MRdHpev/UZ0sFtZklFKmOjWSi4u/F
QP7t4kmoaulWZnIOCmeu9DCBVJztjtd1Bn8XeGoJj+YOKA+zio6C3T0d9A0jzBNC
VZV9SY2N1mG25ayzv985zyYcknVkxWVrAi3Fu3HZOsMbX588III6dvbx7IEAz+Oa
iTNjzUAliUgfxpL8Sz4sgqWkggRauHgecS9ZPwBWGxkESSFCv2gAeXz87EBxAVLm
uXemWjvVoe5M1zhqrFxltEcLPKUxscS3dC8US4qZDxh6lzZATFDHsKMqFaTzDECf
KvWI9DM+vO9/C93OUVuj8L2jI5lxBPoC7/fQM4LuiSPVLjh8UXppWszbkfJhCKch
/OVCSFvuyNulDzxvV3x935ooxFtFccMVzcQZ2dv2kPz+2/R5VpAbePm2IYUfr5SC
0YRMQIYkaJCrcXWhbqKlqywoGTumr+0duaOxLr1x9m3evXsvrWQ+GtltsZmwCzpI
NquCFgSgYxSrgK3/kfTQM6QeEpvMx0ql3XeT3tNOKiDZ+Eu/RlE0WFA4cZqnYJug
2R2U0SFEXsl7PAnQryz+BeQn8uLX2cDiscOxlR4cnXkF4A1y10jX9e8ul0Lf27+q
XsIImW+N3pO50reR3TFHXBcVzlmH+FyRC/AEYfSvxQrazgJnQ9FClLWTo32VOslh
SHXcooX29mc6XIVeOcLeZ1OsDjQOZw/fZYso63VhZfYx90VEc0j7qH0BSoqaungt
gqP129U0rP9z1Qy3KdzQcZrjIG+KGdUPGE/arIRpF+Wcg2WX/8kzX50vHXPghpzf
7dVrcCpxxQfoIh00ht+4dICpjZF0umqisqMfYiebTz0CNe96JvypTdQPamIk4Mha
LRpUkKmevsWS0AordxJHAG9WB13RnlthkvIzDKSEpGsyH2icM6prW+Dozn4TAUBH
qytbW0LJnovkkVGKJ+dZA1snWixD86WD24Hhshu3t5CUXy4efd0BkWXxNgM26aQh
t8vtBLjXN5+rOg/bnSOkBp/V8BJ6kfOF/FkEu87sGGPegZ+HLUynatQHAHEMuR98
YaG0lff3qw+5u2dCMrt6mNK/WgTJidnTyPAK4gqaGPCg/Eu1zpDLPCF2Td5ADFV4
5RzaEA4mmbYClM65yASGH5Oqff1CHFJ4BOH5q0+DaDWowtrcWpriI70Rziy0VTTx
nWA/OlD8pxZsWQRl8xNjhU1+tns7MbmUxviD4o0haaeG0oszNwz28HhRetY2zXv0
XhnQxoZl3EK0KMlB5lSBRpt/TzFtpXYCn1Ao8GPL5qLuOHDPtP6a+viivxclys//
2eU7RR3fgUHm67/0UsAMwr760HtrcpzO+196uHS7Okhd0m6yE0da2z93GjGB5gAz
QPr9cCxl3G036uVCquImjizZwdg5A4GniQPSdMRrpdacPdGd+XJ+3NRQ1iLZMbkG
GH5BZo92y6yVEGKT5nlFoeV65mumnsKDQMXOaiy0NqyGYynCHuq90LgQu8VNiPyo
t7vNb9h1NBUNxamlQ0RxNEzu+LrrLgbcfji2rFKVdU/wUo+cMmmO0KeScy07UaRC
ztCacsMhLwJp5liFoqGrWWYh/ERBvjHJGx054LylNqvaP7wNCaAvPny1uACBn58Y
dFSgAc8AMnaXs16EAZk4PyAEkoRRGfR6+jpAIu/c/SOeFMmG/3RZFpGVcCW/mxjd
ASJ/hAbvXwLHx6qOeDbSPu8IhNc8s6Fqqk0NKfR69HAnpau6V4JC9/0CbqsqkEjA
L5xA8kjdnmcXl1c6prTWnt8VbsEm/57U5JOJz8fcJ4lXU2EY6ahPdVvhTm3Fygb7
fHfw6emup45lILxwhnFOBZKvPa3MXqj9KisCKVeX7GG1HmmH4u1frxLw8fUT2Ags
cAPuLphUODzel+StliZ6dqISF/SGaCX7+npZMQVonXDChkO+vHwwhvFl5PZIXPFj
BLJNxrebwE0GCn5FPglpBHkIfkfXeZCOvE9BJ04hIUuryQblP/qyKXWqUpcNDZfL
HkMg1qRPC1RPtyfyN/swxv+lcaPs4HORLMB0P0/hKBXEpVUIAYfeM0lxDEh+AdBv
oWhtdiAc6XZ3YVTMpULJZzG0vESSrRF58uxPrbyfNsqvYbAL/K5Z3AX5aWV+4X3Q
3tbp9JG4NlOSpzibNAAwvj9bGG+ABRH8x0sI11qCgd7BB5ScxQys+uq5HnPSSXr/
9/SQB5Ia1KvraL1tQ2dTXWl/Vavu3NVDHCdipjQS/HaNCpW4X/v3G81O+oRjb7kJ
h4dUIyBjHz1bKgfPWhcjzwNYp2EsjbHGSPyfzhaJtoy4i5JassVJaXMojJ2te2vC
CSmExJ7OLoW8wfT5PrVLiIpPS2eF0B+rSeHfvSWX7hkHXHQxhXBKj9fVKgqcBNxI
LFECTGChr1uSBNYaNe3ydHT+zhpotkLNh8yadzrSCeyJBEgC9uUJ1OmcUUrGF18n
YcCqHomfptVgDsh/zZnz+4tP1JJI0wZZvg3TG8j/pNw8Y4oZsBEqMl8bCHpeKTwG
RjSgKQS6XM3YYeNDUevi+f/PDEuK9DX/QzHOMbgKVeufytrS3hHhUFdWCAl7QVG6
HCAVXSFTbTM0du7N3wiq+L1eA1xnwW4wX4SZtIK+pP+918sMne7xPqZ/lyKeVxuK
+Um8Gz0Cj3DTIO97KxuFLqCfxyyzmxu1SFGdIUEcgS7H32ifgm3H9EQTCP2D6O6Z
TALfmQ7TjO5xU/kwCnJIp3tgkA2Jm0bUUylkelWcbX9HdAVmlrDcBBHSRKTJ2c8/
zhirRoHTSr2iznq+So3iW0GF/DycChKAYUm4eSs3tinkaON4vIUoYCLG9VU/jei8
QFjahl5dKQ47IayVm7ZY12Dr//zaJgRA+uWxvTktooqIWxJ42/gFUbJeuQJyoPo1
QVLCMgSbo0x4ZxWl89XluibXKN5w4ahxQLOoXBrS0r3ks53eAB+d5oFa8skr7mHe
f4IOY4cwC0mEqko/IT2hNCFCbfrAPtjzNJqT22DXQbYswskRQBLT10fyYYkVGDNb
ygYPNe3gOIf/BrqQX0mNoYB/qjFX642Qgv6H0QzPDJBXPKQctAjblMjcmG4IgB2P
SK2lmUTp5CVHrn8VwEvbjzbRNIhwhNIKQnKTedkWuXC1VFwpf4RQ5UH7kO6mH7If
2qY6UWusebsGC7yxRSHqrEZ941YkVjhlO795YUHOvFlK8KwvrxZPW2qzSs4h6eNQ
YHI567liuqJ+qGyL0zzj8/L/nXrELH2sSD/QHQKNHJLZPhVByBj/GBZDe8Ktedhb
GC1Mv8uRfRistpZ0ghAPU87IAnbRQZBz22cNBjgAKhK63leBn/bBmSZzNeukp9fw
qwR+V/tKRNiNM3yig/cdbwUH6Dbn06ukh1tdbbkbtWN2V2TAf3TZevsw9FbU7e9n
GVTIhmAdNLR3uYcJYSwoqyGMKvYDjFDLPDOXc0cSyY6Cso4MlyXskKb3wLgkxvNF
NOXZWAhn0UU2290jtlkqCBGihQB4jZy3Ddk2Ov2Z+03Apl+G6uPmjlq89+C7aopf
s8epmF09IbkbK3zWSqobgKjAcZLiTxziE9WenS0zhV4SkFaAqZm4/vGve2FlXJOM
nw6Jex9DZDf5w2HyRtuhfbQcBcP6enCe0LZz3M0NFvZo7BQ47SDZwTuAGyC9P7Jl
54ODMPjFfpv4LqU/Uq9l49By3hVo83vCPo0ArgP5/euVaSpgkWViULFQRkYOixZ1
sKyqifrrd+OAOp2G1WY14YjVwWttUFdQlyZ1q8NVXcWoOhKg2MVak0HmxAogI6kK
DBxpj9RZ/m5ln/Xf0BMoyCFfDlEUpRPhmkANEXcC0DIc+wUDAIaLojEH1fsFaATx
APsUxGE8PF+I6gFWOGjQXg8+YtCHXdTT91U512V/WbFY+I2WmzkiZAbtIyuKqLgV
ciSCyV7c+NZD/6mh5NtOFuji+UX+009A8MTZbxvHYeLX9cQfl9dRJhPLHm7YYo4a
A6267UQd6mjvny4Q5LvXslv8YV+atARv0osFsXRA51WrVcP98QLfIWY1FUqWnP/0
qVdAL6lmQbpZbu33EJ6P+l9mPM3hKPFxm9EACFK1Ozrz8PZNK9OpLIs/UwBKX6mO
Mt9GKbOMRvAA1bFnuQhFFC8VQBrFsPgRhIdUuDOnyMO/aUx6xG1Wo+O3dBap7M3r
GWPioKgyX3To6CC7fr9s3abTucXQQeZK9u1En5MnYeV+iKBNq/8GheO81AgFSbKN
g0wERg9m/4ryQSyX9QKzkjOuXuQUT55m5lUh0ztKmvFjbrm/TfS0ZC3fOyTb2rwC
RaANPUn07PkwQ6Bbfu6FA6Wap+f5MqUh84XRYBKM7eiN0dlRkPNxEBB8YytYemg/
7dqpofqEe6++zjYdrqWFcBmTgiuGkpaA50nOAsb8mdu5OYcbfwIip7SJZRxeIBNX
hUdGdB1AGeOZod4qHLIpQPCkpRpp/yIUElM3KI0X4eFc9cUPi8zyPDFQmu4HYDG6
EUy0ce3fm9X+yn1QgsarIOF+ZaqFQc2f10sCtv1J2gn817obHNvNTztVNldnMe39
gQFXBIJP1NzL7qOH0t5Jar+YDnsMaNPImuzJY+QcZ0V35ZCp9PgNxmWEsjAMHRH6
xHk9YotCbyaHQCzkLP7C/9AhYJ6NmfoYuYyBEVRJcgLZKSqoUPEC57RQPh1qjH49
mL3yRZ5NLXofsENwt1L6SkXS+1xZ3TnJkCpLxvOGY9msJ4NsartgDyyRh4jf0ZT6
+yFQf1etph3U2MZIoO4/DPhkfD4U6msErrcK0C1OcA18NLp8lRTBaDbBKDQahl2A
8TP43esdHzpVeN3LVqLQa/GKUibutkVGMUvoDmdvjK4G5V8XXWBticC757OsWcqe
WGLZ333gGT41GMLhUHYDxct+UKA6Exwtt41NWqj7jP/4QCgapPvtGAeZ/TknmnnJ
Yjr2RVkbaLcE4vfLNCX+EA0Jgepn5Up2QwOopgR5p8xND+hpqh/xWgBtSQXbVNV6
1z8cjYWHEkgg7nWuvlOCATyf5jcItQD0i6I4RAe4eDP4FU1PB/2QgTWeDub0oE+R
pqtJIBpr57ouHvxepgL3yEPSnkPpHhk/Qol/6wtK49UjSZGXktokh2PduVe0R/Yn
mjVCrVG4t1WaEWxr7ckpoOwyjh0N0Xp9SPCs7Xie898R+QUXNEzL5tZMGGkpNUB2
OwvLtHxNbaAS6vO+UPg+iPqm4uVKl9rFYpT7JpkTiswVqOO1Reypsz+daXTDO9vh
B2TjmcXSmHc1wQpq2eoJnlTa4/P4ggXQjLf/Zbmw39w1BsTLWViTCEH2C024CwP9
ZaFeJRx+/X43h9Ib2FXmKZru6ZRkUTWLAWFj7wmDheX7VRhcCmTiOxThoblZyZwB
Q1pBtGwV52UVMfTeBC5Cx/k5hWkwo3NVpAi/QFIfqsdDEUXnsfG2Q4FT1bdkuvYR
iax9mR+MKP2a7ZbhyjjsgqjWXmKYMzf/2+LNDt38xS00TH1OolgxyZfxOrWcLhtq
GrNcZRQsPelfSBsX4vzBZYbetEdMfmlp5/+9ujeiEfYAcR9rmx7JaPYCYn3vaaoG
2ycC9acFYaY2oIZrWGccLdCZtoY7pEDkVMdA03MbSjsCZzxDtJJpGnF6/LKhvIfW
1NZ0xtx9/p9PBxuEpSfs4Olqg4wvuE4YUeI/y+b7TEJkiVNycuVnDwBTLzKTxMln
LwqZ565B+Ki0Taz6+hel/cA7M+Jrl0C+CTrKhI8IkJYcHhx9SjHhzdYWa/K4Umut
PF1Itq+4ilQ9MwNGKJwncFhPRYDGxh3tVpW3muXuIMPGSwkDN/eZusGV/btMB50Y
Lz0A4sFhLuvtKv/QHCQcUPFHA/bAN1dq52dUb0Urb2JVVvjFOxW3D3An4E9AywHz
sw3T81LONu8ZgedPsGjD6CxiadOLdhaIfIedquOLyZpKCW7+799DHtFiCTJBq8Fy
Eh6j6zN8FQZh81jWF1URdqUaxTCN7WVbgcnwdlebnfYQ0YOxocjIWkt0rYWZ7m2l
lSjEIbTZhqouIzo4yL4Uh82Lq/LjqxY/ZWMQSYBOnBdrAL/GolxOsa1IzrPE5tso
6ADHYzCzaLACThjfXEOZxwTmSpQVMLWdvJMzQnh02h06jg76AWTKwW7X2jkn2fHw
tvX0Bbww5aZdv1qmSpuDGi3M8nhNylCnqZ4i4s2rLf88uqGNNAJ8jA2EFz/hmj+M
c1JBEisOoYkMhj4XpSMvVLdBf07iFTNkXprkjvk+2UQz1xws/xFx0jjNHmzQC+Fn
w4hKSQDya7rJ+tG4izR+Ve+IifAuKCiUTsDVncbPNxqtVnF1emEpV6GoT/HV+X3y
roX2kmnF6nO0q1D5oIwKNmNvd2Su19UogvTOE9nHpj1WWj8GX2rZ8y+dwrtUPvgQ
qyxNk5XxT9EU2nhh/KeondoBJx/MD73UiySEnfaetShHwnpcKUfISPvaKu5edmQP
rIElBKObelSVxIu+3wD1Hq9ujwV1093kUOuF7+1fyEhsYe3+Ox+jKdaVNb0Od4tk
olbM3473YurNZWDb3c2Jvzeiec+soF/lv0QnfvvDlHov17DajC4k5HypAwWw3tBN
RtyknfTvnMB/69CzumjNg/7hvILi3xuFlU4fuQNzkY6WorzUyIEUkNBRMJueTyGo
s6f53IfOcI56zBCbq5oFLm2ETcar+qTPE5QGwCAptNmr7iG6ZT9yjM1usJ+Z+gXj
iP9CAmqjWt0fMots3LOmXuWlFyPHXDNyR1ySUVugyvZASChAIss+jOWdIGaoI2cR
gEHShMTQkobUfujfmOSYcRb+iypByxV5cVakJ5H4Zguoy0aVVrV4LEh1AkGQbELv
+inmVxlS2Kkukz4X+JrzqVc6EGXaMBnqegI3zM60V1Eooy2FONd8caRXWqZqeOET
xBN+lD4eOiNfb1hhZyEeJt6soacCSDp9P1pcwAn2fjPmVz0ZhddULVmNIcrqh2G2
r8kq6lQPpCmXw3/TNLF84fu8lQ9SPFU3pXAJZbG5cS/7Kf12/bsinZ8v0OvU8iGY
T2/b3HJ44BXQJIY9gGC1komc+CYsQqNMbEzvLtR+AqQcGNduNnkbNwPvhQSOsWTi
VjoPFqaJm8/Lm+H5yg6OMujx+/Puhx1R+sARQ4YAlxUx4cJwr2UwVLFlh41tzSRW
0Ws+okf04+TIF84/gMmo2mQ8J+jwpgr97zBdq4WGEPv7s+VAoD+MlyObjF4WaEmi
PBfizNziCsepJ5uE5q+gBvMze3jZmPr7IB+O2sHUUvvnjl3o96NgkNcO3zPQ9m6y
sw+6LqHYdQDtYaas/eJsiUbqw/gDSP8ZMrsruR1C3bayT0cq7Q4nw1a53eXK+jb3
nhO0lJtUyUzOiTfE8VyenBMp+eCD8SiiVjez9Pk4RfYVzht4x9DsUPd2gyNhEuun
s1TD2hxMGyM9wTVLo8lpO4UBdXBQU+12c+bCrKBVxdVRoBcbz2iTyuVqWv/gHadg
hU0Iy2P2zPXHCGeIXRTVPBQOX03yi9Fgrl9/pQfV/DFJBf4b01mrnlbrHiY4yN1/
S9TuiUye+ymVWH7W9DaYDmFA0iB3c4NkylH2NxJQa1IxfMiEspMARWP3xM62Vya4
0QqGJLIG9DrBbXUgqG7SlVSrwbifzv94yScOTqi2xKAwFMB/GwEZ6GTiJCtAZVsv
z1C4X+sFT1/cO5ea45Qw4R9JyYNxjhcnGL3TGVKO+MeoZbzKSxF9jF369zzpAqoH
3a8HSbozz79Q+n54fHaa6R0ptNISCUl1X4mUoss3s73IfSadXgOuGMbxaEIn6Atj
3v0O4SpMy5xS9zqMEUTvrWW++yH/5ASpeS/STvz3phBZ0fKtq4Nhr52M7EquUf+O
Q6yxYqR1tTl1WCWcxOW4N6zsv4hCKPJ4qKBwSYt1DggeSiDoYDSQd1+q2vwXMsF4
eZWxIyvVEx2gL5wxsWc27Pbr83HRAsi/w9vMcc/JFqgLEhMuBdRt6DwZdakffdVU
Hfu2iqYzvCvvkZE62bbaXd/MD3u28Uea0K8GKw5deiNSTDi8KWwem+mhCPSS455f
Pq06ST91raulc5GMEEQY2d9ZM0OMS09qxZeVXwoWa8/VNNO+5WiR+8FyhCaIckUK
PP4S6+t+bYLdTofRwvK6vMtRpeCFUMRhN2rrh0mBOEbMgU+V/smcDVSnxlLaKoM3
6FIxIKHt5KEu3n/6HHgNKRqeicqeRZsy3Gkvritooup6u6Kan8D8dcJIo7VII8Hh
iZwauAoYnvGkhgTNLrQkvxScRj7ufMukoQNVTq34E6/yUkEgy8T+qz6kOUMl0wlH
8e2iA3c5E/ZF4vu64eja/uxUwMgjYw2+qZ8ETabF96H/vTBDhejslgVnaM2lf89m
gYejbMip8/3IgVomd5h9ank21oOc9fIhOGFm9G9n3w9RnWF8ZY8yYe6ZMXEKst08
/94Wmw7Bszr0qMOuArbUkxM8gcV/5+2t3KbtfzUiRVN0sQOtM/aW7FRDSrVc58zD
gYGhCnJYEWWjKP2bCY47ChfOO8tnqOKZ34zIFbl/eSy71Ggw3Fcv2POBMiDJRcSu
T5izDk+1EOMYhZU9lVmXAQ/nQyaRTIgmN6T5u5f/huERGgtSgxQ2Yev/J3iHp3hG
cYr6hhVh8/8xHucHv6hBmt/PNh64bDtMTKpz+236RuAy1SBrtk9ze/qjXAUq4rNS
hEf9GemxIMYHdX4k/a3OBxcJDq0Isa5/uXbyO4TogvCiTHza8tOd2RA4KapLMeR4
mIMMXdzngjFbKZjlvHanhQb97m/sc2RmunnHG9FQvuACJh1K/pJOXDkvlPt7uV2B
upYNlF0EyqIshxKFADvOZ/m6uvkdQOHPoxDmkSArJWV6P8aAdpaqLNh4lhwQTGxW
nRIXTWb1Oxgo/MipcH8Q9H5ob5Q9TyPYKfgG99E9Oh9BTnVxs8yj+BmfMGHM4FnI
Dpm9HWe1wpiWkbVuajA2nquHMnzzDu51EJcKoQqFNc1nsr5rJBgHxPMX0gYbbAqB
MUXMQSrw8yRqjrRPaiAu6SRp2TuZ2gb99Ptnf0/masvFdsO2AkvYSNZp3nlCdOLi
TNV5pPoMh4GFdj7ooKJSkOa0mNnT8tRsSbC9Zi6Zd+Twka4Kiqv0y/osfT9lhEHn
GtjqA/ZoPwsEMwf8L5s1TRKvqnGHGvbenYpNmTivkySpomenxvtRJ8+r+nQwLjFw
ADzfAO705BEOOUPSgw7X3lVA9trCjL4YTi8wuerQUsg96K8NTc0cxmYSdsjoowuD
7sFW+OtCZp8XrjFFBH1xBQO3eB6gLnGNlIsxDlztTuDPezSKwdmG+pvhdoPWhsWP
GZFWVlVDG6W+w1ED1AzKJn+dM/X54XwIARkfQK9BMaIrmvaLmDf9rfe81+YkzOLq
Qk467UH/cpPugs6CeU/+5Ipikm1IypbqJQ7khenAYM+GN6Z0Rv/9mCWb8u0iC8rh
Xk/kRBR32XWqa4VjMnsv/0d3WzIJhC17fW4v/OBWWsfE+duef88D8TyQcy9mbPXk
TAdkP6jsm2TxYMyUv/JJ3Zow8XF3lPtwbYp4OpNuWcVyq3zeZlV95AmpJB7HCeYg
fh0zzWrzJnRMlTRWeSK7IsRBAKBvPWLoHqRRQyCTXGhm9YzgXBaCo6O1G5tf3AF7
yXlZpO94O1MnT/pThQN0ns7qMVTjEvauCeMXiQKvZ8D8Fx27pTqoVBZFTbHzsMLE
Q/VFvpV6c3QIaMxeOcmgj4AEJtnOuOv0u7+7r93wR8l5YwlInbBxMIn+kWREzrUz
LDsl86JX+JbeONYuKH1mdsxxLxHJpFSU3zOeBuDdB7QKK2oVH038jYH4mjFwA1eC
GGfk2ln6FueRu4suvoG69PW208mg9LMgKEDcoSIMwx8GGpsbYvQl+9V9MhP08PY6
hW7jXo/23coJ+Hb+ZCs0JRAfxG0+nHRTVx3gWdb0RHc1UPZDQm0NKqpyhBfm+9gH
8hn3ZbmMaI1/+x/MlvMwej0+S/21tFWI3NFIQHf0evl3c5OqqtyhorpPHeFw1CWy
bDgnCdNPVQFitcVx9sijVq8U1A4tT3k1G7NHW3KaC4nydU2i015zz9lBfyfm7wbT
ZyPLa/iqp2dLg530IUgfWeqeCHsmugKhiJizTA95/sL2QXx5kUY3dDmOhwpkS856
U3h0c/iPk57OrZTKJBvDvcVyJTKb52YgzbOEGxnmPnOBYvT5F0qQ47OWxTNQyD51
wKLDrSVNT0zLSCzcY64xY0Em5ZnSQi0N7wBFAKbUppYirYbOToYrMRxREdqBhl3c
q5jdZJQGYh5y87ydN1ysQLetoq+uhACkO5lToDtw5Z+nXjTt2uj6bi9R7qgVG/Ro
GlhUgntlCS9LP3pLSbaa8rjA2bPcUuhYLmgirzMsst0WhenzP34SdAVmU3URgyy2
7lz4nw48T65bGMgbYt9TFLj9G6EPB1f8kKHmXAwQ2CBu4h1PE/4C1EPo01DazIaS
SiCMYujNVVr2t+w+D1LJFs/moO564excUv9r9KRvdY5u+KDFe8gQLqe1EEbDLe/h
qqOQY9ndMtjMPGP1194C64XGBGnk7GKpuaMPyZDXU/uPkUJqGNOpZAg3dWpvX7Xw
widkzhTF7qgG2AhXQmmRXCQ/5Eal9ojEYGUidqY1e3f7pnbpPcpNMdMU44BuH5Fl
nCQWkKTjrtvE7z+nRoExFpd2TaTCqmPdDHrJdT7VCmllisM10ZPzrnxNOtTQhoT1
3Ug277sM6X4iVP66NsN5i1q7bVnBxCwlVfc4gD7sNbgIIzerxWMVz3FR1OcogQrB
+hbGx5ygtzUl1t5EeqVF3M5O94EGOmuTeK04bFKynBFM0Mdrv+Oc6TK7f4LQ2YjV
hHkJaUA7eSJmMk+gAdH9s/6kzuNUXkEeotvbhxcC5RIEt+JWlSiCywiLiEaYC1Rm
lqpgQ9hb+x/XkIpbdzu2QWl9ZoJGB2dV1TJ9b0+xRHPJYNsnWo+hq8T5tppD2+iG
K9nRfJ3lheMEbEXX2h1BhODNHEH7DXUdRx4a2KTbz8be7ayTJIAb2P2ObGykymoF
9G+LdEutY2d70qcjqP3MNl4YOT/9akKq35AJZmRLWrj+l6gINe5nI6zgjXm4YfZc
jrcD5fh3t0bP25mj52k0ZiW67PNe60zsOcdNJSYS3gHe+BgLSj4XJnW3KO4BZV9m
vg+ns6vFWoyESiOfKbHTiu/57B9qJIY7LucR2xBzlyQsT/FBGg/+JTDqztDwqMl3
3T3yPg6M4LRaYU6M6jvRSegoQx9V02V5e49E5m6cKAmjxlenH+1sk05WQXCgqt28
U6eDLjyM90tzTgdfxv81juTJS4TUATt2zgqAArakuuUshO3lzJDbFqdKww0khXPO
vIV53oKymp0zcaeLJMv0eC4KPeHoUfZuM71Sx0kGFNrwZYXml1cOIKbHJRT96kvV
Z1LF8Hk5DUVc6s/ugu+6a9GBeLHcToN2JHDoX/s+TRtG/MjEJ+W7u+Wo1H6a9zII
sn4f53C+HcQwqwSAp+EwdkzSQVcqAwlGFcAI7RKsc+E4zQUtKbCNEY1eUuYLrSGe
gc2I4f4/mdkToX3OzmVHmpbWBxKyXejTaOHOW87V55kVRvi0eRoiRbFunEtsp33R
LdwrFUWgwgEULgzma20kuGbcg2werLEsp2hkpykd/ucEuoX5q4yesjRs2EArii6v
LjYMgzpAzOhabC9HE7mpRT7GW9quaKwnmOLkZCpSV+g003Bo2bpWTCBZGX6eVTTB
9OEXXGgLjh/fhTc2/iQc1klbPOXX50o0SReRXu9Gqkto3T6DlROk+Zw0JHHZxdYL
TPX3HF8NiNWAakL4T17woI0iv9J7+S88UGky11ke5UxlPDdVejA6NFpTYBaZv4gv
4K/SX8OHckUtaFkbZIA+wy667fTzfK9NAVvhCcPA3qasB71PWQ0h3rB7lDe2lRxH
9bpqYiGZuooWP9TebkkHGIU75u835iomofF5QclgfqC2/aMp3Snyh/TNTFnVOTcA
R0kugZvLFYe8MrNozgBPKDPrytLNQTC5N4uZawjbsAguTCLrAsUoGZhDERP8hKJF
k5echSyZkktiN0IMx9L6LYtSFhrpwPKzbGSfPCeXLDQ0EAQZqtLkK1L/jEO6i1e+
Mhf/5/Inke6lcM/Yp0T2Wx1xGhTbTBLrAzOKNPXYAiBd9JgWM22kBNb/1hx5jvn4
lihFQepVHOH9luiwxwRKZENpEmr7Mtq4BfRqrSkBuLSSbT588L5Ae8JLCAP1RGYm
wD8bKNB4eTIvuTIG1NoBkxV2cYKNPnFhQ/LpKH55jDEEA5nRMr+mBEXlaMPEgLNE
8T9M8wiAaQbgxENKdJHE/ArSwPwgdEBzSddapLjLqwZnPNEUTZ/QGjsZ/TDhUpgE
Q9EShqoAh3XX8ImPKq8mSpz1WTAgarf5YxQmfsJENwprRCXuRJhPqVi/u0LbpxKV
KJ3Z03j3Oyi56sF9FVhMQEjZUIoNZf8qXXI72hvcblhruWaouPtD2RQ6gW9Dcl8i
G4bgqX1s2BPbyRMDBOF5ASeHJn/Bhawoz2HYbT2NJljh4iNKbIWECUzOnhS+n5h8
Nfd94Ge4idT/81Pz0+qWvWvIBhsoHdBJaf60nibknBqSHdrwMZXHN7djKhaf1mRO
VNPrnUy3rtzR7tkkbGahY1JqAR2ovYS3H10KGyctWwn4tBQMZzeQklV7gf1Lox9m
7A/NXgFfrHWlDwh4AEfobQNjzaGx+QwmiUfq0wTOUD5eFP9YsYAJBZtpyGLbB7bk
6Efb/qzxTkaMtFZ5ERIetpuHlsR1ZZunLqvUoRN+TCy1fohPdGNhhgxYqir7jjHS
0Xd/7+3fEuX64GsDvTMVe0EqPPkP5JDcEtkKMOYBWCsbHH1oEny6QgBdTFTsKV6T
gSPmFMfzEuluO0TzJ0rOuHFSh4UYtojj/P031Yu/dVz9yU7xJv2Pc7xlIB1WA0LU
2RIlJl3FHES0gLbB1klvSI4spF3vQkdVF6jhktR+F7h0fUVCN30DHGSiS9RwDkF1
X//9/PORlIJ0y1jm9gcpkvvwThwHIGXJpEX4q/ElC2G3wYbufGgamqQLkN3QrvWS
cgAQPsgvti7O4kgY4XPVChBCobXyHAc/xPcTN0hC6KoYUBZnyLiDzSmK6J6dvQL0
WFOjWgKFiEg4Sej3zCzbqUSeM2Fn5o3bSUX/aOEM+ORdafvFNcWD/FjDFpHxcW0q
reZ1MxEAVhXfbKstzkokni3Q9wY+HDhHcogzKfCl3vubgSX4tvdco4G+iwY8UWoR
XBvZhkFneMdIm5T40cWtO1/WKoNmwnXuU42rjoVXfzHTa7f0lxQD/leRqPrcf5t2
ylpC/6sTlkKBTj+Stkp3Uk/OGYAxqK+bl2GBdolhIGu8gaqXq4zfmAmisfUBk/jI
b3NnhQ7ZjlL/wpbbNiyn1H57IPn4zt57lFLHoE1OsBult3/jK1OsR2GrNyiv1NSb
dAOI7NqKLsZH+Ei78RrxXE/kXJP9kN9nUYuL2bfgmfQHPwAuEOTMxIB7z79avrpV
sQz3KnZvHRQvxf1B5GDASrmFCNITbYr2GxTjtzm8a1FjPEkwOGx5aMxkiJ1/gfnl
OtFll/7xTjbBixSo+qyGqwVE+tyVMaetaGzDan0hK/M8o3T3YvoiP9FUnFd4cnMQ
d7ph4U/4Z/kygl1YiLcaoHoHKSdcjduc5nekuuQY83sRQxqXZD0exnmBt+Zx1/WV
bMKlBcTegwddwtIgUXemg6UCZ18qvkwsBFL50BWcwJt5qnbiwRTA6ISLbBdf7MJR
dQFCbH2Yt6QEziagZ4Hx4DgSOjysK/r5rmrQ5wKfbGWYoD0uuGV2wIvXFTfsk/C+
jh9qb8LJNMqJndkwKxiyeQHdL88jxiFhezefM4U3EP/9dVrP/6s0verYVfQrJFOI
vrCfsPfGZiqTGrTueAgXYcjQz9Q3xox667uKV3KQ+wVp1CWln5iNkPgbtvKUrqTk
U32kRelu4dWQNHM/15ZHci9pVbBF2mYd4tCZ61WoA6DK1Vt9734AfXrg+jvKrT6F
fEspPQ7riyfd/iSAnAkhuZrDJBJiaWUPLEN9CMNc9HwknB7gicd5s7uy73TQZBPL
mqeijTYWa4CnUXrGWbUfNLtNzvTIEx1mCGniA9Y8FtkRcXe6obZUmlP35LxNCgN0
wfFDatsVQ57r84Fj7PqXSDSMOcUdFGPVS92ofAC5yT3FCTjPh3LyhAA5WPNbevcb
Lzt8na+D8uujsWY881xN5BgsO4soKbA4I/5fFYMeIUcoXxxOTa+ocjPUUcnM/dpl
y+gIvbFLYU/IgPxV/EcbPASLM0hSqyw8J3GMBJBtI0DW4cTcVLqyvlWbr/1aTpJi
jbQBX21F93bfkenzpx+kM8KFVApTbV5UN0e2G1vPpk12wXa6RQc+hbhJnWNrVdAK
W/fEWv0ixp+Y61S+NsZB73eHvtUpcWdnzwjwZzojdBy6mFHZ4RyVGVxFFqY1CELR
LyMAh0rsYRU6z9kyPjx1IiIaOrjH0CpzlT3qGf/7vFjqb8EPmmQ6e2sFkE4B48DV
PDcAR3ycm8vB5+UcU/t50Zdz8q0W5GJSRe2Zai9rdUYuphhretb1f1eYbGJyzkUM
K73M+7lGbxBNTptbhLWaSOXPasUWPaZno/EWPBvP/Mi0N1GwIYgKy524A2Ajxekb
NQp9ba3ixreSiT5BnSjbvgHmzzl/Aq8skRJTKvwUwDkhEN4zNzRZdqvmtpCNg/JS
Pbqm1evpoCmyEuekqfDrThsskFPxTFmTn/A/izVNjviP8qx3/16pvVvmQ8c7mPwG
+/LEial7T19NSZSzDtUmQMQhqc/dTTf3ss97pWTIrVBQrUQyJuwChpJg0rXK27+7
0bLm1hsAbE9khFRLgHzVMKqW3VwVpTL1knNUJKQuDzrXK+LFlzoMZoknNYavD48m
v0udiRWdoJh6kxUMUVje+2ykkMLzEB1KJG4foi70B7THOiAzXwtvQhDKuRJvY9C7
WC8ilgq/k/EnOcVUQ46ubf6WGlLf3XeqPZvHU0ENBCXsy/Wd+n//UyC5AbW7NOy4
sPJ/UQF48+n6rbb/dVgjITmdgGCiBxSFysdsstjKX6/RU/IO6SlzSqXNo3t1gLe2
aM3W9Sxm6B0qsXU4c3uNk4Jf69YeFZ/XE7T1WGsjanm85N0xscj86igUFXuGrKbr
fnI5ogdW/e5gGdo7xJFXoIC4wCTk/7TvFDbtpfaYE0L5288diLAWwFRFF7MctEjZ
JOGXzMwElePSJxUwF6Dd87sXPWUQ3rsMS444OKN8+pIbfxOlVuCHzRHtjcvNUyTW
AGOvL5mGTl2Cll7qn+cfSaRP/fQw6OCguajxtBp9wnZoG+qA8tCjgPGGm6Ama8O2
PCYtMrQaJyVk4TyS9f4qg5YqwGPEhW0E7K0zYuR2Xpy6JUJzOH05+s3wApqJVtbl
tMfBIzxwn6t1rjIXQseYA+DbUZdEIEL74LW1NQmxOx8=
`pragma protect end_protected
