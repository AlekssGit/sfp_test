// clock_50_out.v

// Generated using ACDS version 21.3 170

`timescale 1 ps / 1 ps
module clock_50_out (
		input  wire  in_clk,  //  in_clk.clk
		output wire  out_clk  // out_clk.clk
	);

	assign out_clk = in_clk;

endmodule
