`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
tLGsHHYQjWUjvaJR+WLOaM5yuRlC+2J50VohUM+sfd8KxjNPGGN2CN1vug3EI0Er
LGY+EpTbNsDjK3h36OTUh8vRBLEWkRNcL2f4kSjZzuqMdfMSCF8WQLrqL5blyiWQ
3XXbe261AqL1nMrdHE9jCYH8Du4iqKVNeyeodEqbxxc=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 4080), data_block
AfklsbZytq40WeOMVNBjhgIdk8K4IeJWVyywQDA5c73z/b3oLsQDwb3vjBuIfrDQ
MDLjnbI/sdJUCYltorUTIEKH0/dvWk378aHGEu5XBpPksMbHBLSAZZsTFZLzjd7O
9qDef6pU0Coyoct243yZ0WO/xUvYXhQL9el+5kzjVeUl9bIuXM9nj5r3bLoe9/2m
iQv/giE4wUcSn77I48YTjNXSKMxUMxsa61VqhoLQQ/wYwXz2AXe59I1E6mveVqAu
HAn5+XjWo7gyocSCe1vxhrP+gewZRChpev+AHShOSCYB2wcR9MpDg0a7vzvu+sbV
ula3LEhfv+clUL9jGKCQkLFIwr4kjcZ7FchJVWhYtZVqiALadC/v4XOPBOsoQPve
t+EZ9jpcRmiF2M4/WiqRUjkmrDuW+jGGfDArGUzvps0//ZM1aZfef5FlXhcQTNrI
dUXpq3R+r5nMF27wugRkyOYChmeVn62/rZ8Po1uylmTQZcup8LJTYtaFJS6N7mVD
dyZEDZ/zABaGb35T2tUqaMD+trecWHxAJrc2JbGgIKfui7BuSPfkZCVplmp1fqED
nXX5a6MV9aZ+9quyfl+XwKPiP7gE7o8aDNavBvNzzkevfosXk3JgMANYMISLi8jG
PNMQjn+eZN5m50JvabvHcdq2XmhmLQQ3oXEZ3Hk5xL0RIpY7v2ERWPmDnK1cdPQP
d5rHPaGsxRU7wD8tcfb7YiM8PXPf+aQrmxdzvlufP2ABKQ+AXELtlPuOzxjkFKEy
k6om5uK1JS/fn6gwXefdLfyzt3gEgtEuUdj9/sbHfu9kTJdKho5G5gJaQJ/9zjuS
lw83S76VO6XEqDurP8nSMrXeXjSTNnZLKEiarWdWVlU/NB00M1ChKP/94skNjEY7
pJYty3bk1m0Vhvt0MjblE4GbNOAkE1t0RDg/260uD3Je0rd/U2KDLuj4JOTgp2cV
QZ6WvXzSnVAUdXm+hUbQC4UKnsBzXd0ODjdrz+sr+F8cx8h+OLAy+m02YmgC1thQ
ZN6hcYW0BBhQPUxz35W5AgtZw+eW0A6yCRTEFR5bMc4/YiVAVpQEAehKoRj12ByI
5aCUlkzaDqMdBtQjhv87Xmi5gSdHBzzkTHIjKBMfxPvQ5hzi5ztNZz+oxOgeIYM+
/b4eM7+X8RzpibTC3Ke4z4FfyVf+Upoyrbs+j5wAOw0/dRkw7KgPcjVKEvXXfeTQ
XREERSCFwOPBk/ZeDGGthkdPEpFLmkesdGbz2HYU8rrKB0gLcmto3zWFFarVLIXZ
+adFzU3a78opD7YYaWAbWj6JCkuvjlUU80W/kDqXEvvhB463vgVCcGBqBcH3FpZ3
InH9YJfdUnvQFG0ul3LBmtxdBJmPIJksgXMqZb0c36GxKCJtCA0y3frF1ZF4wj7y
ytkUyZDKlPjadk/N2fFDaCxbZ4XELsnPAphL0EAefMwkyR+rKerhVBXvzJi1Tv1J
eS0AjeoPcvWQ9WoyEjM5JAY5lkWcX8yhM5JoJA/WCvUlHJF3xT63L0CCzPUgEH/3
KjThpxPDeIEu2bLOz4VxTGAcNr+mSSKWI31GrCm/Gy2PRrF2bLiFQL9X+8PqnrJm
ryeaf9A8r6E41sr5aROHRdmmARxpy2sp4ORx0BS0B0udH/5tFfHMJZwSVLtwiJgF
2/vL5SIJZmhr1DrLysk/mMFLq+U0qt3VXoq3BF3AecoB3BK3FyUfmPNcC0dpRUxN
cSd2lLTTQqOuD9odYzN0YYAeF5IutPO9owUzd3AdTnjf57b307bFByd4jLOpkK8/
65BsH8TkfWpl3mrTuis4ikiFCjcVYz138QXCWU4kGjwhvIK+Q4vPAsc5OEC3gH63
GOYfRbWqAf7f1WqWne6aJjMgLhV2FGX4nlMXFU4tZ1qYOM8dXAeha7/31u19g2Jb
l44BO6yH2h6Eh3Ri2gxZBhRYfKtbI76YGpHfXbkNNN6WrSnD5G2pUT4112+1G8Sk
ssEf/hDaO6hszDkcDXnvAk+Q2LbNvEitMlnRKoy9O2URmPBxUJezcOEKhu63Np1p
IQtF22N3qWPoGu2zKuyeY9QzQ047BCHPMZtencz6/QldFP7mdlH0n/YCN25Dvmvf
QWrkq8tHIiYY9oc3wRouddX5EFL4JiuC/h68SiyG6IeibWA2VSKLLSLh8VGyGXn+
FsC/Ad7dWhEKYVYG+aMIEBe2NyvQO+nb/dG2uq0VxfEEmOp969Y0ckvg+2/2V13t
K6IpY5z3/D21F9Nd/PTMMkw755nq46uEEkhH5sH0NT47sS1VwCBxnaPCS7ctNJzJ
2hXTIKmRT7qVtm5UgpBTovnLZeFhpnKoBT883EBRXNT2xUdQowlBodHiH7oBYSzN
RZvaT9ubKYH3KwC0vvZfnidW37XtHFoGC0SbtAylkUjK5IkMthVe3yDyOs58cGfL
mW2Dd5/twWU/ck4IB8MZaK12wd93IC1nplf4VnA7BB0HOg4nqjPNUGLYHnwvcWy7
fFoacfTGpCWWIKlSQ6lMlO6q6aLplOL8Ks6xAbcIUliTcgagylPut2NbwRPu/Ss6
o9U5/CGMZgHpPM8ETuq9KCT2RAv/bae1oI4R1FX45xzoI3FW4Y+3FDjrV2EIlpax
Xzrn39vW0IlMQd+vn7Oc8X01IGnsWaks8FhFdcwDI+8r1LMiier+vJfLAjNsXJi8
ii4CFku9JiLtArRpSk4wUyCi/l2Z0UQ6fGtSBY7OGZxbOZrSULCmwOqhacsoGe/U
rLAfSqXajJZXlvnGzurxNI7NfVoiFajzj3J5adDOMww0Aq5b+NOqAB567Jrf+Fle
wxEFX9EaYkPn51bOGd8nqq/hfw+7K4dOioMYaBB7SYMoTeG4eYsXFu3Wo/55DvbE
HnpyorbFQKWKQh4POk5OHMF9FZfakefXsNWraa0yVvhdnKEqsg4UZ8OhvBGTfcrY
i08PLWB/51gNh3kRhFBSzTbOnbWlhAhYCvF+a5WaKzayGseo3tIOaaaMU26AkdRH
+ANlkyB/S26btWAa7Trk8j+xx3vGUiogvfXHX19FTjUmcP+kzREETmDKvJj/n4n9
Pb6Rilmyhm+eRjWwdD1e1py6Msh0NRaIpoQkaOND4o8yQTsyLvD+2+qW1eMZf1tQ
i/fJALyLqDT50Xd1kZqgJ8U+GbSvmmHRNz22ukhWfOxelqERiYm2VmHkwn1/qgW2
jJhlJ7pCD+h+CnvCu1xBEwPzj7ZQ7PFTmLC3NRGhevqufEDLIzCrXjOiyO+rAT0J
AoWzapoQ5t/U5chPDlI7vvXlf2WM2TK3RIzV0Pk5UuwR9K7bWTGAN3x7/mXgaqlT
gTs4cOTyR0/oWpXBXnL3K7+JLjqcm5PDFmBHz/VLaRmMXmQEeJOhIHhJAX42uxvP
q+EM50sN3fJuSbVGgiUUF+z17zVdLAR0f/bqPmaCtVTZUB9BKcWvn+m0dfOnYMOS
FXXq2wgXgahB6zqwvXJsIMRJAstOa6eoq94Q/478a32ibd8FEJN7wsYPZEmG7rsM
rHEtuZVcgmTztPY8fT+aRRxb9rv3mW0eeZ1wEavRnce4bK/ZOkFNsPUCEf4MUNhZ
DNFvR4n43jmd59j90qgClKEQ8YqI4D+VeZP0/qlyIp+aDroC85U2WDxMVj/hi/9I
44xkBH9abyEq+C0Chfm6fvTVxKQIRvFJP8UOzPpXUtk5C/0+dvb1EDiPROJ9VHva
0Lp8HxK7baj/+Ze4K/YmafgFnWNw1UREqr2M3H7HRD1Ry1YxEzLtqwTwFlfpz4ue
DQx2VLJ9KaaaFjk1HOTW4xBeE1lymla3s43AtDD486ot1EilxMPrtSpjuCRstgTY
h1R/5b6OpuaQxQPgg/Uu/7RoLDxjSePrUWqB3bF5FhuVcfwj/C9IKjOMbw4eeOA/
E8kInOBMrIojPt6/eD1bm8ASuh81FzxNmpUOWk9VSyna0EK4P4xcDs5Rm3N9rUTj
onFrpvlGno4YBaW3xm6NnEbN48o6lcFkmnd14vHBSPWu6n5rdRFBEi8RWKIg0hwS
nSV+08wM04L64uOuhBhOr3miGa/SWuSAcssx3pp9qGhPWJVwUZA89pgSIXPTm1Ra
6vZ/u9WV+pWupwgl4axRnXzeipIccsv2vhybpZUKdHZ7dnSYJj4alJ8wYrw+7rZF
/EwplwSA0IHK0Y3LJbQuLMMp0Jaam9Dricoc8/l0TDNbtR5rcCkCA2X9TkHBSxNA
Pqzkp1i5+2WKwuFkER/kF+ndpXJv9MdTGGsfBNAAu0Uc1GhEud7rq8UgY8F8TBAJ
fPncU2JRa58VU800SUJIrtZQ1tBHEsxXSUN2ZwVnwwIh8sCn9ygQ3Ikp4rXQdu+V
h7hk9DtlIuWm4Ae53MdT53eljDYxW3u9DtMk4qd3GrO1Rz8FQ3/LYcQuVeWRMbAi
C+WZ+rftYVgXj7M7xZh3OzfjSgiIetOaD9LEDiGRg9xV223I4kLyAlwCzrHWzUX5
WuaYhScvqDwqUWXuDi/KMt9tIB+1E3UpH6+4pWnPbgIM4DJg6JKAE/QoUvPeUBzL
5DkSxVxaEJBxLaM+ve/qO+HADtA2MXctfq56MBbrWVzdvklka0BAW9BFvMbP4bzO
OgP8bZLssw7zYFID5Zdzp7pxVCf5NHwoVbS6LN60ukOgx+YcUa8D1wdREREmTmFm
imcReLTAnE9gbJtsHO3PDvixRHyefyWtCp7cttqmH3wUBDNGWHbPuDc//KeyxYPV
EMUpajPNG8XFlsjunwtrfAzmY2ypqZNvSKi1Ho21SuxYE5nWDX4PfoOydqlq740K
424BNvdoKoKbWfMEDMoAC85wnFksMnQYZgd4h6Q1qEkROUjhgpyjIE1PAxbNqELW
G6SyLPxZK3KxUB4Ksbdf0xRPYy/uoqweXGJ1k2mi61MxkZ5AjQNoy1TGcH6O4r9Y
VkSHcW84inBUg6kLw70KR6xsY/mo//EsHWP+ipuxSewy8nYIkc0qHR7WvG0OMFtW
0Cp4LBqJbKOTb1OFZlKdp4mwRu48Kw3OG3C+q+noVKPa4Yreh/8nfu6S7OBK+AYV
K+4Q0Xdy7u9KGKbU+tJn03A1q4Y64qHY0Zs7gV1/o63SrgP47sFODI+UmtDoVnPM
ZWbNvExvEfuVLTwmsHtfQNAI8D3bgCu3ibk1SPmqSf4SCudqDnvmi5Ym5gU2ekfS
eOahMjozctTRNn9xDc0XOViI2v5T3M3IUDCdWFzw7Oat48jaOWQysrZTvDecHKC7
7V+3EwaOSpZ+j+p3dmRbm65WHlUkSJbfjm6+f6Zb4vSFMLiwLaExJDFYWzvEBNhi
PAHx5M3goL2mxJympYD+NPRzGeG+28qxO9FJ754Bu8GmwSRg63hIbZljtA6pc84u
XniXufqO/ckPMbkra68glaa80dQezm0hOngcP97D4fqP0cqjyO1GSGfddRCF9bvT
`pragma protect end_protected
