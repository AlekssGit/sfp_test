// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
wYUUIBRfNScyk69aqORoaEakRA6TJLnCEcA7d0wMKdSA+1tspy4B2SiHLwww1nGC
jj5FAXgLGRBNjMXBampRPPPSXoojqPHPSLDGgo4nNM/88kdbk72MRuGe3rez3GFR
vSkaZUdBpFC9YaJvzgogXpHtReao+8n+TF0xvEnO8o3ptY68HucVXA==
//pragma protect end_key_block
//pragma protect digest_block
el5WBWXUX0MVC4+U2TukZ0TLix4=
//pragma protect end_digest_block
//pragma protect data_block
HXX4A4A69To08ML9DjbaI8uJdbZgod9EJyGxlgEk2Cqbjr7DAwY7XulzBOhExnoh
I1vc9Dbl4YBf+GafPR/EIivWB8vBq34awNB0yZQ9BU5byATenMQl8PW3MgzIusU7
r/uBuNcfdiEK8zv7fynacmA5tEGmk7exEn/WrZjdqXuYEGcSf21qD98TWjFN2NTQ
gsLPFKNtr/NQD/InJ0bARhUVRyZ8TptUFt2Hm2uBOg1D0CT2K8tS5Q4i4/2rKtMR
IKejacqjkMnp6EDHdVRUIqBfHbjeFJjMiN0iLpXu7Ek57MYuatcdOwDZIudiX7VK
GbLUPST/zx8mKNBf4Cc3eGICnX20siBxBIv6Wiw6f1cjpyme0vn6nLqmwxQNbLjx
zaIxkTLnyPwklCMuCYFjwNa15o8KT5+2Ly2sWpiD8rJiejSOf52ABEy88ZLcBYfE
yp4RcGw+tczlBQHu2cqNAHzIhjJBuX/KhnrwQ+djbaPuDin/9qPm0fj7cdm69Zr1
Y9Ws8jQUbMhspQ5+y6BEo0ypwWSPT6FsfEaT5jUdpMQmWplR1qp0NMIkBOPJkg7Z
nrtiy4af8rey+Jq7XEmQUlz0tk6utmRnd2dTPvQ8ZKoRkoj/9W/Fjh7PCgCdzzUY
WmyYiO4hpXAZMjPq0EzHgZEjy1lHUy8vm4In3tio3esBOSIBURkLL7kkunytXNsO
C0VSMD+rDAju6+SXt7u8aFYijbJDYy7f9RbnfWHYfv0jSMMp3ojyZSIT49dQv5C8
0yNa6BzrS/d4rHae7EbsjZTVzt44lGxWIlbR75NPhufLtNGhmHsIi9h5eaozgPGu
l0rCAxB4lZjiaMZPqPygywp1v72MpcUqph6Wak/OniX0zk4N9kzyDK5UG9S60mDR
2+9K7muwvmVzZ/5EPalzBwpRMTGuy+GnLtcBzQU2kOM9ORylXZ0GmYF0zOvfnPy2
ffLUU+91jHXXOkLlb675+L0RkEjJ8ffD57sOOPX0mCF0E3FmZ19azXEYQnz/4Sp5
gN6J3jGdyvK/1PzTDMGs/J3z7LG3+3IhAYAGkNamwxobTOTJ+BUlSyk3okbopRKk
/T9kjyyRgNr+7zjzOhtQIea8zrkChIaAaYgeloTxaXsLtwrH9LSdDHxPMh5jbs0y
GqSjkNj1MWfYG/MpPtLWuAVRUKqqHUNaG+hvSLc85+hyh6I3sUeaonggAEz0/W7d
j9EkjBQaD5aaOwnk7Lsfm4SPV+zsh2LylqLSeqqUBi2p/BsiEtzX3aDXJkhQ9js6
avVpyp3Ae6AYW1t/gK9pTSgq4zAfeZJ+trUmbGTd0zPxNxUGmSsF58+YNbejGyGD
FQ2hp8mql0uf0gLYOtTODn30lAO0DwcfWmaC6l0YuKRhsTFQuAf8M0ygkNFqQuQa
qLDEG3A48YOYmgxL228pwQEwpr/4qo/p5YMPAoeFIWQhFxd1+uWfIEhkrRnl8mnw
p4MG4snWfRrJS2Pgclu1sBYMqBW6MlOGiIBmBnBFkMZ34jVZXvfurF5wuDgTqLmT
ONZEf13Xy0irFpVEMMcWTMh2/fxnDm/kG+QnYCbGwm3ebFnB+RBHzQoY1ISLs/s4
QReWshg8L+tC+rNCcTbZSgwRs663f+XP/PymqfdUI5XeXpwLxoYfv6DO0sMBz1nf
VYnnqz6NA96+ae8V9Cj4F8Asz1/JOWwi5YCkPknmtoo7lpgoTQwt+k9eiL6R1jsP
UTzoCiASsAIkWCAxmnYhl+qNrKurSOznR562r5jthXHFzflWkHy1kt2Xb+ZeuzTW
9pCl5TQSeiJPHRIJ7wKDpDEwE9EmFmit7nz2QYnHTQJNGkqLo+fJ4A5fUsYf7Leh
ZsIgC93mvkt9CP+CsY8q1X1wlcM7iEplhTLBz40bjAFJ5xQcDljF2B0Scm4XKMDh
9/YIbw4og9RI3epEnVXxL4Xi5E4AAKP9Q8V+8dl4cPxa09vfHCWwVdLjm6kQXIvJ
4lf6OU1e7ALYZLdCUW98lf/0OFCpCgvTApQqQvnrZAmOamHNZM9HKaG+w1ObnIZB
oyuqxf2IgDvZd3lEverJsR7h8+v3ytAQBCXeWsI2/188ZISyT3bOyDRt9yzaaLg3
r0Km4zHF4mNX+hrLNOaJrOrNMfTD88TsK5FotUfTUhURd00ltRHXUaC3xJaxy9C5
jjcV3A++466yONd1qVYPopmbr7NGjufRszC6qfMFfipm4YrS8qM9RM8RPanenU+X
e64pE6k44YEYQpEzBuG+LIlzh9SrPBTTPSr+9EGy5k30/VrbMi3vc8FYfAVfw4r6
zPx2coF9iuGkXuqPr0E4rQJl6RwCSgfCgYHkwgB9LNJ1QIDPCnR28q/W3/ZJlill
MahIJ+xwusYR8vHUK1t9K2S4blRaxWQWD+hXwyC9vmQWpvwiWbgO1f94xPGPn6Ao
mb35gScnxHKsjagyj/tzW7zjw88eBxvsGUTK0XJHMJZw4arcbkU5rNrinG1UisnI
dNA0WxFf5IMcMDUBh6lxKirTfcdHdBfW2Rb1nXzTGK5scMmSd+zvM+lOeXE5eM4F
G0by1hSBh22aWbTmK2lnFBEi+MUT7FP0H91O0WQydKlb8dopRBo2qe5EoZjWaof7
yGrWZL5B7QcoYCHStc8/yAJaHH/NKsNcbiCxZ6decz/swjLRD6/ttGyFqVVNMENs
uCwexSIDfS4NMoHGJIgVb4UGZaXm4zrvIR9XjcmLcci6MY4QDQJ9LgD4r84Q4xXR
gNqH4mG7M9omsJrsO8+Rps+gF/z30bGvgf+O7G4xnqm5zhhZKD1QhljxklU2ejY5
nYzluwjJGflt292M1Lmx9EkfTJwgJr5luzzFhQsIK7jUaRveAwbBGQ8VCNLSgJZv
bPkrRXiwREok9uPRyT6cOPpGNyupEQHgurpCeR4DqxW8pND2FAAZV7XvndJhREwn
ZX781mBJwyv3MxkhXJCFhTFdG11zsKUn5MNg0ia+g2Fz/ITxhEylQ4T/PO5vrUOj
LpwEx18LM1eRsy0eHdtLNTEr937ptDQ/TNesSyS6T+cwj5c8eV31l9QJN7Xb8hfb
v5Otsjq0ZedYzK3w7iLPSmwmL7RjIoex4QTpUvzVmyICH0AFN2Pk0HJ1BOUKzLlf
KPdMP3u5KnbQe1qyKThrrRyLgdM5I83Lvp03PsSTrF7iiF77U0g8/pAFOVu6MrwH
KqY0RSKHpNLjvHk84QN+D2pW5ebSLkMpl5wt5IlsSriD0UEHQdbAQt/K5FPAEQbO
WiExEDnwOuJwP2sisxutof6gOfuh25ho2X6cAFuKIe3jd/7iEU373vGwH80Lt3jo
y7xhBlURIeyWYZ9O4L+Inz8nBNhuv0ZnMJ8df0Y9SYGRl7UF6i+oeNZQALnYOrau
vBrWSGjGLpVZnpsokbtE5JrIOS9Td+RgiuuZce0BPkH3ARnzJ14YADKtlgQYc2XN
fcju/Sn+iBWDE5+uoZ0gwr3/YgybD5PrCL0Y3newZ2dRjpCPuxdXpd6wBRcNdMyX
gQ3r52s5MS+DVV7QGIshr6ZTCVYqkOUXS9Xd45kzlRsXSxGHc7vd1Ep58gAvAOtR
LJHHvuVgPX9nnq32tENW2UIU7g065Pc2njABqRrtu8hVpXxWVCdqyxa2EaKaw5go
BwXRKN3JmsfmE0Mbj2d975/9yvMolIE5z1CYBeOSxDmKqmtCYza5lxu3GPnbpVzs
Ztz38LJFTO+3aMVXMC7sou+HJLMTAzq91tvCyh9Z4ty8QpKt8b3q/XopkQY5EESF
v28kmhXD1GJdSVMf5P+XpcedMlZILWoMjeCscz54u5HVfSVegAJ7cYv/y+YrCrQU
d9lv/aDJvsKX203YVn5d4EalqszzSfOP+yFwbkuKtVB8OMc/oHYjJq0oZl99P6bN
K8EQxRnbUB9kSgub5+VPOJKFiFwO6mZXmDUidiZByYjQYH/aMQtvDbtPMRrHqzTV
YEKxU48A70vRdUzcaxnNvFuKfgrbISC6zkEfCTqlgBC5v+P9rEU85YLbG+puDQbE
N1c4l3P8fheHs1t4lbBbU9sipmCl2W4YogEtTnzmyzKp2x2X9DRuti/Q8cP004rf
p66N+mcOMbhDBRIVN5DQl0CVkWpMJq14LdY+Fh8hPP//iQRPf10dQSLCAv3/Z5kj
0VtKPQTI+Qkos/ARy9fqpkam94/vyf+fZlBWQ32WDB7Ex8/n/dQLXZH9fMP+6zTq
gbP6EQkFUUyd1O0s3y6J0v6WCKrraB6O3cwYQEGqAColfOfcBMQO9xx6PpxWE54Y
VKtSTgAjMdvBuwHWWYKPa5+NWVYRimNybdBxjv2fXQHUwxGLuq7jeZNmIppIyulT
Xi81w1KZU6pQi1gbGrFOJ1HEVKW/5XU+YS4pVi0PAhywbox5SZz70D80pjMfIEdP
b/FmP56od7BtGqQSx4x6Srcfa+iw0M/brPYGGZbXrpZPnTdNAMG5VOqzDE++lANi
gx2RE68BX7O9PTDIWZG5I4peBjJSfVQ7RseqDDAi5QZaxX52UdxuADDzrNNI1Hv+
nUxSfAf5NYtFlyatKq+iOZwTO746B5gj1Og/b4Mfkb0fzUa4DXUtq8C0SlwHpph3
4ZCbY/d+SLH0xghA2N/yVcnmrTaIlODhc9KTnTMyfCLjZ+vbiaFWgs60ZBOiQ/DN
fQeoEHVs9jiRgaFLX5WHoDsfbLrv+v+sGiLb3Q6R8FKUlzsPudIPhUOcAm82NB77
sjFEr0MpcfC0CexqZsRr2GExy2b9pjnoIvkm4YHissT9ITuyUDRc9Y2cJO3omaoe
gukGf6hK4fPU3gS82LN/LkJWv32+oe+RIC6NObvjQFT7uDvZtPs4uI3gnEkGFj4G
UwcqKlNIeqccNE/CVIe8vmSpqoQL7gjyOwZlnoWfxuqCoKCOK93ha1fITPditEet
ko/3ZOb62EODH8VnvwJXNeEw6IOn0MwisL884+u9z3eG9OPdUWOj28Bj1/2lnv2k
TPxwtO/H4powRB1zWfid6NJrBgkYyXVYKG3hvnK8wlIMlwHqHUsiaqkVlwISr9VC
BJ8occ/s/VxxhFmp7i2G+bWtfg7hJHJ4X8eSYFetflPCcra+XYRSSolK+rE+2dA7
GR95IANYxsEeDdZ05um/GUwleS6sRaulj/nE1gGcmwlVwchyFbPdcz4OQfULsgug
O7+qH/4CROfFk9jsMiYpA14qNi+y949tADZC4yG5WvFtUs7RhwjpcVlVY9f7xfGO
ZoPqOxqyvuaY9l/U1lm5+TtF/W0iTsfJFJz1iLEJ1/ywLBOX9sX+mkvLXfk8obLl
ladvTeFDLksExmqeeoQ2x+um4lAWt9e0TFndlup2m9sBNeeNOETvXQ0efoCHNFMf
X4ZTE4VN6gHmjtc05awvenO281HfvrZUdCKMgVK4BsgS+AgUCMjFiDoW7Aob06Cq
kX5gfOl2FgWXzKkK5Ak2zqmcikx1ncncUP2JNRLhxHdTFv7VkcDQPVkfXdNK6trq
p6G7OojV4Km4y6fYotfJZYjIKHV2UMiKZbV6D51TBB4hdL0VPOHV/Y3QbvBh1goP
qFbk7m4kEBVbfP39yAQ1UlPyRCtEiEc+64k0UHYBavyGgOTVHqeZj/hs+5IIWwSl
fAP1JrOMXbsMsorPZxOWXUpKCnWlsuWfrKF0Jz41Ih0yX/dsCLjF/m2TIQxjrmje
61nSGIKTdWBSqCHiUofvOEqxVyWmHKdhcnCgTcdifmSZkJy+MXPAyj6Uy+yBZmrf
JWdtpBlxtorOIhhtn1jbEleadSJas9XwPTcrwWjym/IGWsDsKD1NMWMpkkOiBwKh
2CctX+Hcza5rtHzesntJsFWtJXE3ZAmewKTDBuhfZOB+sLmvMkwACVf2ldZJYDmY
BWkPSjhBUJabthIIxPFt2oGHuHSGqI0LOSwMB7gjkqVr0stlSqz6CH0sq82gpi7E
84YbbaJi/6QJBK0DMNiqHrknYocIbxHaTfLAGf33Z74ou+ympnnyHGjhTYku5FWs
Nz99SGrnkz5zbz7GgYAZ5EHPx1btRt2jKd2R9HWYpSpDzcsb2tYPOSc8UwRykV6m
+kFvTehVJR6Fn3l9vVzhMT2m1ra73HIMt9r1RM6j6qc19PZb0N8D3KN1Aw2TJ+Su
PLcmTqKkOqBfMGqpuTZe6hpSeBrMRmOPos0Zwhox96S39T+glZeyI/ZTJ+pI2SfT
AC7Xy/0xJ6RajQXPy3Gmv391DHw3jUoV1fIy2YYuIBJgWvJatxj44blzqp5gClDJ
pxKmdY6AvWL1eoVJHut08HEv7xaggXXXQFO4C+kAjEdAxkDRLFtoFLsLGE2kbMf7
Ty7YCHWLJ4ZvTdVGiwFsD4pA9tyVyn8I+yeqBEuh33Gg+CGBIFm+SQoSj2rurNfq
2bHwDJAxm0t2pP0p0YNhVCk6xZRhNGUu0bUNZ1EmGspL2ryJSeuxTfDaoJ+w0Rr9
dIyD7T4M05Q5Qs8LKvjrdMi2ApdWGRfiZFUIsWaDC5BV4hrkqusnLFd2j4htukss
jfyPUHL9Kv5siGeDXyljb7+yCIFAQzSjp0tw51ub1FSg6c0GklxHQcIvrAxG8RZN
94g+DYQh0VRVBudvijCWGYn/fYQNBwQOL/EdUPpeuUYWnM/h4bEvCGToTUf5mw/a
Fn/knSFO4z/gsw2ORDUIRE+7R6/jET1z/4GF2koFx+G1hMhw3wsH5gkf2CTO5ii+
ZJTDBpQ8B8/gPEGdhYtVECMQYy2XeTN4SSd6IV0bM4Q3BNde//YNXorkJLCJr5+k
etTt37aQoV/gBfkkVOyA+I/2/1VtddK/++xedWUP1/vQUTTayE0/J0+coRaHaclV
3RKgoXfBejBb5NNAlGa3NRb2Sb3I7xObXpxXj/SrdvZqAIY9HA/HcNdXBsOu4t2p
vTev2Onn6TEXWYOqBQqIIwaAILZA3ZqBLrk0vA1AdY1wiQO6knfnNKBzLNm6agAY
NzxJR6P0lHRw0o8PRwfyHcoXAsXGQD4DiTQzRa2c7kMqjVzYV/Mgk5xmnazbnrO/
6fS1ceHBI/GwpgYwt6ymhekV2Q/DDaYLlISOyq5IrGN3xPyOXOs6EIQr1O3vT8LI
+MK4ODyeRLOs5cgA3UztgWRRhVofwAsuxRVgiYppmW8vImvyWu3QoCZneChc7dZr
8htNYbGwAbbd1Qq3GbSijbsVOUxOjZ/bJLHz/YrRbuGN1NCxPRZCQ4zmy/5lIkZQ
lJqMaw2g8UX+t3pJjqWL/koEwnDZVp/oLzSL0tJvPUuyB36udx/qRdrJ0jd7q0qM
igtZgwAgUMFFNGfqV69areHtylpHHoIwsQ4ugQpxgFSDIPA9Mx29j243w8y9xcrH
cJnqeRrkBTB64J8fO91eoFy0BpJRb3yxc1t4UMW9w4O4tnJwvxyu3EN/xFphnUUo
5qwBjfaLJfBTpobbsUKS+D7jJSq7jSWdEuloqK8cvwimjtH16RuVk73uNA/iZTvH
y287t4NUk9y7VYwjoAn52ksIsk8zPNn2M3UsgiVxqmd9JoFQBMh7USzr4myCrpwB
MCYoAGsTS6jrqinmIUXvhcvYcWXu3JRZqlLeDfnBiUohKo/SrbqaxsfEU+5htg3t
o9NB4daWlag8R1uMuJyZBgp44X+20zrDfJucWhfeoYBuvEDtiuEIVBEL/u6x5jGm
9R6Hefs4of4n5xhbJ+KRiMf7Ycgw15XEgfERs64Xc6MgsnWE0yrLD/Jo3VcDpFSk
8axPKsKGw9loVMP8D0Wd0Q==
//pragma protect end_data_block
//pragma protect digest_block
XygJQj1shyh0XkivlYFCfUC6JjE=
//pragma protect end_digest_block
//pragma protect end_protected
