// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
1eYIzymq/BShXVFQQ8meP6ClJAah7kn03g8A+sxlKKoQw2wS6pvXeynPzQv/svhl
BElQJt3NyKxzgDOfEzn/nyu/FTcboCebOjwgTcegnvEd2eCKpu6CUYAmEki9tkb4
MmLRT9SAjJymg7KrJJRE4eRuquVG2Zgn0tOLjiCSboQ=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 5232 )
`pragma protect data_block
PSgTTx7zKMJC0TCFHl7R0SVf1E+VDudS3E/ATk3K/YVxL18dMixG1TeRKFiDC8eP
fzqiTpNzFdLZDdghxSJhPazLxs+ZBURp3+9hMmFf8MyqpfeGom4o+jsNcu1EsBlT
wnfH+80R/WLWg/7eUP/MS0XTbIc3lg8e0px0AKMunCteqJwfbnC9Fe+KBkXN21dp
nNg0ZM4QtLqsLya5Pyr/PVMJX8P2cJKxUYt4YFZmWce6kSQH8mP3ai8JnQHTKXVo
nuRFkzDZw3NLcA4gtywkEScWjNNIHFnaBk+STrH2JyqiHnf8wlqrNm4olLxKfxGC
u0NjFAos8NuHJmXhFHq+l7oFybdGVP/4ziucWwbFAgxBWTxLtgse9FrKnFg8UWKs
x+KwhqV5MCavexClX3RGC2fQeaa0zeFVBi0TmgLVFZxVHCP3yKnljtQb+U+HIjSU
CUGdKhf/JIVceC+Yx9I04YkyScP9XF7loKqPfuzwAiEaWZk/NuiGIYIB7JlUaHEJ
xB0v9qR/sqMcOtYJKL3Y/nWAiwD20WrJI/mKhEsLTmSNx9iIT+AyxQFIwax3xVft
mmd8Xld90rz3OMQmyhuV3nv5zqyjeIM6+3y2bk3XIAxveDJbHMWmZAQ9mNxvHabf
hiT2rQZFXM7dtRLIs8F3C84V70WmQwmfD7iOiwdt7xgySIc3YsemWucqdvEG8LVK
ugxS5RkFZzK39SK71qv3aQgCSuYzBQ+uYXFQRw83pGW9tgJxpPyEwgP4BCmc/gLm
aJ7qoGCaUgQCkQ981pyiy6mf+E9F+vhwqNvNl9cuQ9Sl/ddS3xw/iWD5CDqTm2dd
qdFBg4Vtg29qgwugJgXyvqlvezr68gNrsPYmfz40kDYynT4jWBcqGmM4TkAPSnyy
r9JbL4YEmR+blCIRyInbCjV1g67ktNRGe3eOTyucDUvILxEJ5CHB16cmfkCH01yl
/TPTvLFDCLkjv4HLtUexNdxKufDnsEAO8lyjU8QvowaXQE3ei0Appn4a3kEgYVho
JO0dDBn5OU0f/Vl/gogAiApBY92uGWWo1lmVbA03oXopxeHpwZ5xy5N3NISOnIqR
Jk3sVrtzHQ4EyjWe7gNbIeMdUJQjwl1BSAAccL21iCCbiLHS08x/isP6YnufcCLe
98C8AOUmTBjKhRrpL9ME/B1jxsD8VElSu9XtLd1OPMKLJFrpdrRwQ1IkWcEL0XgH
8u496pmgZ+ZDl3/053jt018nOAWrX2p3K4Loc7d67uJ2TSWOgYtIcdaVB1ho/O0S
zS2CCdHK5xh4p6uI4e7S148C7sYRzDQyJCML3HU9Os4VsWx/6SrQB1q0JkbCMbdD
9ZvDjk2PcOYxp+AmEtQOpk8SUJXbR5ipwUIoodTeSy6SfJERfPhpvEZ1AdsxBGaF
Cig4ye8Molr79RYHrD1Ff8ogqSaF976kW8nl5Q1K2R7Iwm8hh8DFxEnHZNqcvqqE
z2c3ebEPbHJfFYuYOGMc9bB33KsZRlLZwX3qcvhN79lrFraZDBMX5HTLq3ewsk1n
ZnLXPKnJVGRUSgg7EqxcTBN8YbOyGUgeBNQcE5SRPdyQx99vk9O3x8ztQT4hehHu
34vA043n+/G6niTO3A8qZPXF7qMME+nUp2Kbt1rZ7P7mLUFRufyFtRi/5m/V7hzk
LhTOgwK6pSWG57RNbllWDWAZQQqFdNIDVhylzqFsF0oH49yfFX/7h62R/BzGfbGN
O2MXZMWRcHIuJtM3el8t0VZvwb+GqEkz9L9XPx5NDj7rG4TA3WtHaAXiUrb/Jfsz
3Pj9pwfV3b5Se17m9Te4ekr03H/d8c5UP3Ar5r4OugOUnGaKLa2O52pS9mK2YQrw
yNgYIV7jc+q9TGjDnrCoZ8JJhEBDlYXSGZ5UFzPxcYBfusyxNVTTQCRkN3HFi2jT
emHbY//p8UuUcwlF1GkNu19acFIcwkf3PYgW9zjLUmJgek+QZagFIFRjuSojiSAh
5SKKpJ0kJO+blv3E0FtsAuc5dl1ALIf17Hqy/37n+8xCmItIOprSWiHokO3IzaEp
9IDAzwjBozxciCOqUSAm/gMeJQ8kI6F2uLP4FAPYcbWR2TQK6nKjErENHRFHJ4uN
ojEbeznF5Uwpx2RzhIpwCEJxVKonQrJntsN/1ro3892DIecouQ075wnJDhSZMnHk
jszZOz8rfUGlK0qlHpfd0O2yXxtdGCZoiyhxEXPAUBfHO21/YXnZ8JYh1yRgnnE1
o3GVIgWTqpegTzjbIbTia26UaxnIMpo8p83DAmygYmdhgJ6VEpUUT9HOeoHKqZTj
Yb20glGvlTw70wmc65rkar5PTmPBi/1sN8BySSKx1G31Y0K49ZH4sxal9uya3OEJ
o1lyuX6Y8H7p29ECQNQPZeTLhxI9Bqlxk6+CeYojebM/qhKIYjvo/GJBc9cAPlB3
1d9aGh/yQxZbSeCJSI4l8DoZsChgcvfx/bvFO8XjqJdQs53pE9FPW0byrJrY5fNF
vHFgnsVdoKKl+YI/UnF7Bji+qM7/aqmsUwkhMFHXwADvgqnvzqWIK4Gpa37QoyIT
aw00NdZHY/ZucER+ky9j4RBbmQoRUk5Y12EobBOysf9+YLlbr2awufbCCd63t0eJ
KcTY5bU1ULYMhukPUsrV+JlhKyS7jcmTF9O4cXkiquIMNIOG7HbrE9MMFqcW/Mpg
6Mo10Y/XpJSqlFEeg/5SFuwjTdv+XhPYK6McDFn60aYpVeyZeCSXC2lq8cFBxlKH
HsRm52MD21SgJq117k+LPaTPlVN8gLHW5udAt2Nc2OnSHCcdV3IHn9n+fVpW1j/i
RHM5IpZLZCJI9qOdoITpS8TjwHg+2ZisgOfSeoEcwkAa0i+7G0sudZKZs2lrZIop
Zdu64nPrE/EST3qt54TMgBl9A9+I4as/NpmsfPW56/VzgRiIqC68es/yY887A2zG
tgSIM7VvbwvQ95I+AZz5S00zRoq24MS7kwf3mRuIaQ+S+MUQ0/OKoZjBWgizniQo
Rv2zsRxK8AZuCxZGPggI6mbkbKge2qK84wmjmFOorBAU4YA9GaPVA0L/jxbGJTom
m9OhJrFIMMahE/QSrlHP0D752uSRMsiHPzZKjfa8xj43fle7XhMIAh03maFvL4O/
3/7IngpRUDSdCBmLAPW6tuAWKT96+oZRSOJE50VKlmZi82GsE5yuUXxUSvlYOoi4
tn7gyz9b4L/G+gpExo0O24ErAGBkSx4n4oI2K+0BpaQSpHzi7zc/ycMIs4cqOUqv
QQCELEop3AccuGcd2/IbPbSrgpcm1UcOWShccuxP5F1GmBlakwZuR4y8fM/W170Z
KX2gu1Ze1dgQD5Slk6ABJZyals5ISO5W1jgZHPeJ5a/Xv6rZFTLsfFbFP63HybPg
Go572CQMM7Q8c6deJZ4E0oNyMW63x4rb4mXxKdPl4460GxYUIa47qkc56zQ59PKQ
38erMLlbpfXPNGlU7yB4+Xv4PoceuRUWZmpWtIu2V+sOxH8fOGk+mVvWMTBcC40x
79yMAexQbFgLElrqQlPrLVcHuhN+hJyPUhcZyLLiSZS+7M+MGXTSkSNLi3cOUX/o
dVy5AZuDydIamCyZbLmW/n9foub9Clyefu8LtiPOoIgtqFglvIZ057lW+ppaaU8p
Gkrx0rMOB9+3fa+4ukL72r8G8wnxaOdKdYBV2uJLjeDZFjhdnaqFuOFYttXc5iDt
pDprm6KAwiBOq593gY9fs/Stt/uYPd9W3D1JY0cKqmcYPIB03iG7cQ9xVAb5fKIs
VKkQLux7/F/nSC9JlnAgx8MSPfKP5Y6A0EjAPTBFc1eaW+gv1HxpxZSHR7YE9pNH
t8wyoIwAiv8yRautKUCosEA9/LNUYJDfYw6wRVQ5pmZTeSCH5Zu75COqQr3XSZ2/
Dmho9UROvPYI2epCr8v0cnXYmmYbHwIlSnma3F5VMIXn2Dk3bV8C5nask7h3KddP
Vh1an3BUJlFxcOzBkwlZb5hmAO60CYsEex5O8hPAeAHzXSEwSS8byRxGw4sjfqN+
6fz7UL0vSiHyPM0Y0uybhTRrDSYqOYBUs9U4PzZJHv0FCHCjjEcuku2r6uwB8djp
B+MXym8Csc4wBEu4/pFCr412+c7r6ZBcTEQuuB1GAs55+EU8/J4quPp13n1wvpHD
n9sOVGifJfcw1Da5X+nKjnPAOneiH1nvhsfWzFgSqVfYziac3FYfBIfSgR7hQ3dd
6CaTJy6Vf3ji16NLgy/rT+d9XF6HSV5sjyOvNrngDYN3F/yqIlaDiF9miTbsvrhc
utNPLEjJfJLzKN7Rqdpm4JbpSl9hqe0+TVF6tScydNxEKU9qHxg4w2hx4jhUMn/i
L481rDkbdaReBf4zExMa1UUfejlz21Id7SdAhILdkmkKxWcy8OHxdnoQOUvDLjLm
os6wEagqIB5I6ccVyj3GwRuv28pGbV3F77uBuJbDITGu2Khog3nGyNbNGH4gUAJ0
47FMkBiXfcEwKyjGX1ROb1fQsamRS7QgeQGq0eXJe2lXcckv10LGuh+j4zoIhTHn
Wzb0p1eiK6l0qQr4uEpbe07bWcb5HR4dKEEF7qqv/+uc4k1RECdx4gbSHeqFSJFe
/R4QhU49sSrGHrVk2gaLKRCT7yJq8rq7BrLu06nYQGX+WAbnBe7V3BCLZvOzuYbk
sinTYEMJS/IHfdH8n4RDXspJo8mT/W4kuvyO6lvxV9TrLJhsE0MGU65cracHaHk+
pO3yk2zMKq0Mwy9sjaw5WEZY5QjAmeIhB6pZQfZgFb+k+5OWbvflb5Iq6T3zahce
zxUIJSBvb3o6icsh9H3bYAyD94lrsNGiLcHxGyWfhEMKY8ECQPkI4cdus8R3gw5h
iPwAbAvABjosQfna9JUFbNLkgYD3Fem+jXwasRXdeIfp392uqsK4AO6zdnhT2SAG
+QkzxWnKDs/dxzQGU8JVl4R8vQkCzyydVYMEgPsDylIIj591TnL5xmiEq8rGtWG8
KFgjiv5ooh9r5VFtXIExsmS1Gfn5MBS7dIzII4Up0CP3ax9u9GFLg9TH1ic7N3B3
AVnUcd+EBNLPW7tUJ4YxIxrIvVNsPICGVLLYPxSaOSD4J3PsbIll74O6KrPAWUvD
3bq/cXsNPTOi3TgqHO7RDpsj1LP2Y4adh9o+0cn1SD+cqfPcZdcL/Bsly9XS1XUw
17ZUyKOW7f3pWsR6b24+dfEQRl4RjeSYfUuUVT1HgDRCHTu8S8xURu1DR0yc+3aU
Ehtv/aOXHqbyMaYBgO/A7P72WaeRUO3ZzJN+JtQO2Av1pvqO7LNOalu/jqGiJ6t/
xhYitxcWaHl6m4SsHbzlwVckpNTawyupqXrTb4zUcJQNokL/xO0GpxFTvMuIr6cW
zhLnRlf1opzmPvULVu8wJWuPtH0wmWRLCkIaWuafgCWrPZ4Z0r3oQSxbmVXVU7Ja
GM9J9C0Te+xNYFWuS4XITQquDW9YCyxXdvZCXQzHVNVLQrRYDuzPsv+UZj0LnFlG
FDVDagfG/DXD61A2wQz30bkpp2Jzx/CT7r7u16vYx4N6VuLwFZXthzDwYY/dD3J9
k3ExUdWppOMC4m5cKgekbt/5Vl31VlS5jA8LaTgfNJovYZ7T3HJUwbT1aZEf4UJa
YkcfoU99HgBomlLXveZy/aF5+JS/dAZDsUxXSgNfcWooAaji+PO4u143lM70uadq
BB/L41aop5OAHWxvkbqPm7dJwtGZ6uKFCdBFAQvvtoFZx5ZC4Mclg9jaCKdiKO4m
h34iI+n4PH3chft8N7IuJjhSC+9JEwA9bq4eTBVeVYhIkyymeLkbNNYPhzrA2iVH
pGgA6KHx9ln2Ie2aEOqLktDqN2v6RZ6S7QGbkYAIij8pJGVfm8bB230b+y7LnBGT
7oPeWHbi2ynp8DlmQTi1w4oofFTLKzMVEc5BfFMjmy1ZCYi3U9fVWAgnfPAwXGa+
VTjQsT3rTKgKokNKITkM5da4zeS9NuL5JXA1/PdL2txFJpkYgHKkVjw4n1JEpCTU
8OJcy5On87Yl4ApvNkltRw+0I/RIrbg2OFaQoEms/QznX7lk+atwvRuMLmPjHAN2
lvbMQL+afA5y8/Lhwov8ZDVsx0SIwLx6rMHAl7ALpdnXNnYj2D7V/YdWTlYkCEfs
vx6msGDoIeomM4ZJABF6xV+kMfytctRSp4D2J1v/FIdTQdAUD8WyLdij3CovesQa
70tjaF0d3k7X+u/S1+O/xZOpWqGO5Xlpd8eMzUh5+BT1StfAEQWeCeVUd0Hd+f+O
zi2PLXpeNRULzI0aclN6zemXi/21iDbwran4RDlA0S8ZIaW1dzTONWnea8q4XqLs
anOwgfaJ5TWvRf/65pUwhUQFlEVp8OMSbrmgaVUFKchVlzST+HCxqCS50nU0Yg8s
fL5oUDturoNaosru92YnXcnWFx/kfXDdMhuFL+FELhXyijP5I9xUkFqJVXGKt7U6
Zi8Z3k3W99KKjp74KFXz+ihywA0A+Heccb+70eMIMVxztDoiHyoa2coQGR9yDxwy
EmQwvAiPhVthuY/h6QrjBUlWLh/dmjdToU+SlVKDC4nAjDb2IYrivO1DUZijcR3z
TZtFMQc9X8BcIfaWoXvHif8ZERFuhygMV7W0S1XSAGCzM7fxxegerSudDX0JvSoy
eWcP39YutJdfhvIehnQ0O3yVyTtIMG3KU7S5PlTba/UG7+FH5T7pSZbI6bPsUcqc
MtEfxqK5x0BJrS6AZvxEebdxxr/BYLmPyzFl8lfv0acNvUB79871cMsjgF12m4rH
0ZrdmISEBuSuWzfkJ49YGI/BZ5iDu686crWYRRtyptsllvumuuqeNrm3z+3UQSEn
DAUue7J8XiqflW0kyPMPE0oeERXV9z30uSUO39VqMYhgR69xsFkyidQrBJVrMJa5
E7Rj4B/SuytPto/jviEhBjEwLNzK4ica4SnE3VIw0BgYw8dya8L+ksRYdUlQFgVA

`pragma protect end_protected
