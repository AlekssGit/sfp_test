// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
KVmWWvdN8klb/spi5zjVuO45ihZx12OTCIAXljXcK7i00e/AOhc1Hsv+lFZa1dMXP5P76rtPgv50
UuTJCNk4l8HuQK7tK3W2EVIgwijaOETb7uSgQxUs0jVWy0j9oXeR3LatmkS1wRIVFcUSoraFRJZJ
OGO+ro/5XZs5VR7bDLHSmQ83Ya4x+lzLBFfW+xpUhLRi/+hOn+mN7fVnXnT/Am3D4ZlDzt2i++1+
HB0tERXOn0DpdpvR0CoX1DpBWXU+3jSXh+uRpEVAqr+WUcw0nf/dG5r89Ksu/0iiAQoeFSoLu7uE
Arlr6dRzMPklnUs7lb7zfu4+oiWL5rPY951r5A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5088)
TRwbUSGdsl8XGxAKm0+4YtmP9UFPGfM26iZBZGMoiSwt1F1LXH8I/K2ddBVWtfk7HTtKajHt2Sf9
UlCvq/t+RuEzL54NuIyycmEcAwfpcy5MRyNEmMA/DsP2ewOfag381meiQV5YZRXQLcHWS8RFv43N
Gp3hn6UmQUdDgh3D6kU2rIDGgS7VVKrLppMK4BDBe7yhpIUqWGCCrPldxA8Plr5Lm3CygxkNrlkA
sL84WgWhxPtJ23Vt+Nt77wRyC51vdLF60gqHDOlcDrlA2e5yoMX3wPir3gnHlsSL6UPZF6CgkVjP
H8Jhm88bHy2+nucerTqELWcFJNQJSSWlzkxj8HKw5xM+Evw7g7NPheoeR9EzRscK5ZtCIpYpLC4v
TPOC8Kf/gV66W0O9X9bHUOSnew5k5wpaiUS7BrKWN9W1VmSHuqBLafVrxU93u5JS7dR6NQKQKV5U
6vL3s63zPaGBf3SfyIPEoOyD8Hb0n/Hh/KkiNOuT30JiE9a7L+oSFO/Z1nW5klqUbhXeMiQI7yDf
hIrzVHT0bNiYxZ6EacuwIA74S/yFHzgG+qSZxcAxdrUo14sMcpKCM4FcP1fRBIrpHrEOuWPm+lTZ
7De+LdwGhGq5MpnSBfLVffSLsaQ0Kq1cw5Tk0gdatTR/7v9jYUfL/nrCi9KiGR9M/efie3FyMOAQ
RTmG7deZ10Ll+wmc70Fyqv+DGiYq368a8yNnCrBufmFRpwJ6DUj5E+krU9cK4n8p+uuBlzJkYYs8
4nkEtdulxbqSuo3jYAL0SRmZV2AjlEqNWvRtdHN+AGersmy559DMDfaYCYoUz7JjTQ5WbvoosxQv
xP9HA6ZaVK0wRFcGkcoaB5rDheeGY9LhqD/OK8P6K7L5kxfSu5kDPwjPNMyJCpHPx4EqpUOnfApb
MK/eXFApsZ2VWGOnYf3o3DwgFsY4ZFNQgUZKbglXuxGNEJesis3t5UCXyK4Izedmj7P8Gmb4AStv
eal6PhuQzHN9GRYTC0M6KLuUT72naY/XfYHBIe/5ByC2Io4ZcbZloLJf1esxN61v0SvmujYMOXG5
Cbip55AX2lUh2/AJs4d3/mbgz40UlntY1CVOJGebPwgaScA4wDhKctL8bYQVhjFgebieQe2hSXJU
oxdvVdw+gB5O5lxLD5QpArz793C6SWxbENDHwA7W8DbXJAVbsD6HgiCGUqJdn8rI31dgKTmlaaCY
d34bOwk/+Ls161FVEIhw1cZRbY+bahn3smMV+m2gNZghWxbFwt0N9tJ6DBsOy1QbwVkSYMG9c6DQ
YYVExJUyFBSiNKSdYdDgzNK52x4C+tAqopfRgVD8/G8i451TTxqc+6I/38OKUInqJtLNrs9CEsIz
/Ij+TypNcNpiFLiMeylyZnr+hQ0UifVtClhFR4QTqttOBU99ucCFj6scTF87cdsl5frcpi4VuHS+
0rAFoqF2n1AuIYNQ7nCJ3XsnL4/2mt1kAm7SpUc/MR1dveyaEXVz994VeGpshyxYx3PiSW/0VwrP
E1beJOf9Rmk4gaLxIPb0BopkSkPwhTlHY1zCi4TuFv53r3/xn5g49+zIIc01pQ8AKrGVSk7fPc0i
xbLmtFJpLsajkld1/DPPFzyJYk7ht88ehHzNjoMgjMw4OGtXxXTYRNNj0YkRdb+mnc+jkQoGor5S
Rn5lr+N75+QJGR8vxTGnLXrYNitKYwawdqAFWc5XLHVs06/Ir9zvU4HxXiY98R5JTR8d2wl4FjN1
i9Yhz80YK/DqwmlmHc75LxB49WsvkKx0LEI0/zF5UVTS3Bgmp8BzYizSZZJG4OngINPtC8l1mBUw
480U+8qiUeD4FK/0ol/Asak+Bm+KH/YanIBU7M06SR3r4+0SRiijDoZH6AWLcQqhLz+Ic8CB9aYo
etHHE0SHd2yXxUPPBjGB64TfVrJB4QLP6csugt9gG138szRc00TofvutVL5EOqAHzUQM3z5x0grb
6OTlnx81/mjEKkcVG5i4V8VmgxVkAKpuj7f6F62uAXXouK0Esfe7Ig0uFwjpjbmP3U3tmpVoBYxe
f8W6ZMlFugE+AsftwfLLwl7r+zFcugQqYs8bWV1D0GwhVbczPln9c6IQCmXWIzZ/ksgH/eiwe+Gf
D+Nd/pDqHejCEzR4BHrrUQFBhcXQsXOaPwHNJZ98lokT0MHaREjaM3w/kb2MBKS7K7lXwUpoH2Zn
eh69RR7tRcrTn87ariSgkxd7H4mu5lz6PpTxuXAbwXHcL+FamUlni21Iv+Qn8hLL61Jdjt3diiR6
dErlITMQkrYmKBBqz8fn25eVGVUG6plTbc7SlhnEeOW3iuHQ9qQ6Vlosjz1Hf2/k+qa5fWHkGKFM
MdNmtMrmrb/z7yTUS+4nawnlY8n6KmJuXKuz8tSjHN/Oia+cb8Crfmy9AVW5Nj2EDFq+8I1tGI4g
92bnfE3+pc5XaUfpgsRstGqu/qIoSxcVlaBxplx/LVlUmS7yqRgLBXeFCn/AwjThT3C8f2/yTBqV
hs+mb5BCB9Ge99UkZPSMG2sSD/ozakWZs2Jp/aJjtjao9VsshC6qS0vZwZ8dh25rkH96EWEEFCTm
pLfoug2sGxXUJ8b32KLOXtcBaulj3RV9cc9nmPUAKxPEDCFrcrE6D+ATbLSSjorHkZNtpd8lLqkJ
C5psKG/OR/8x7pYD8pKlUfyDDb1k/zwTwAW46oApFAMwnmzkE8ETd2hkwvvnfI8u+OIATQWP2afh
siiFIeQK2sFI8sReFHkJtKcHWMr4CwvJmM7xTdY3s3L50xO2lxA6Cq/Mnm37//nr0swiE9AlAarQ
p7SRhlh3uH8rZV66/Oq5zrB5Rm0c6Y6Aay/fi8x2CndQPoxnoRFu3tfhTHeSFFKmm3UydIzHu2ZL
m1aLttNbFRyXBRLiuNgXSBUfQ/bq7OMLc8s7T1rfUaQkALgw3cU7B2TDj0haCLwcPdcna+08U3OZ
pvJjXJ13GZE5GShs2FJr7hLSEBKSMCMstBpSN71sDb8KNm0fqFoxVI/uDntHL3EB7hxarzLx6/nA
16/C7s59RuGQhtOqztU/A4v2f125sjNq7bpFOeXnGDVwOPWqCP5NhlH1Nq0J1pjCamIXtNDT+rZ/
3k4quXOAfiiEpm/Hqr5dmwHQr+XkceYp1xgiZjBoQcS1ZZgEAlWUrWNFy624fwfK+yVrDF94Z8a+
73W2DC0eTx0fogaFIg4Eu09QcxG8PrLrwCNNng6jS6O1jYV849cm0myY/cGvGEOumvL5D0dFJiCQ
YZZIzw/X/v3WIe249pjXCt20rYi9mpPMFsO7qkcC670IVS/ECqoS2tKJ0fHR73CxsHeoqjmJTKcV
T3VM/8IsEbVwEHr/7+zsFGlDhLprnR9AnfzgvjlZKGyAA/DLqer9eHg8BpRMYkgXf8Jen5Q8Oy+7
9PMOKnVydZlFhO9G2FNOoaPHzT8YCrY/uZOprdFxRken+09z+uDOw25baAkmMkKicu/DQKzNM5SQ
PbTnIgCMoikUA+g17Tw38siseqh8YMYLmS022/4Kp9gjjw7gvGJtQAYh7ViFG4iLEWMIdQx7hzKP
y+LagZgVBGItCsCoV/7HqX+vEpzF9cuIsO1hNFajqOO4PXzNob/izDYhsvcBjpOEhIVtJx6JtZXa
Ev8qv+GGUa0sREYwVVEOLrIXAYSJwCOSV/J6OEHCxrm7KcW5CbnQTuO/SqwBeXO/9AwEnXAUlTjq
7uoDtVmA9JVlIkciZQY1GKVdkf8MRxOMrPb1j87qr7DxhurATUnOiKUyClzhTBF+A52pgxeTMc35
f9irsa4IdS5w2FAvB7Jncqe2IccO6+WVvCfODTLXkRrV/54BJ9a/rNyseLSKCp2yB/KeIVdIuGnG
qWMFYs0TgQJfgJe9bm0FAnulOc8CCXIJoLFM7gFchFw5PqmrQd127ocxrusFHx8FRyaX92Bn3rqg
c9ZOdr/CDonZpykYQfk2UWm23sNQhjmYGfuIYkXyHy1W3KKj9EIQSei1tLz5qxQM/iOEXd1eul09
KFgexiOrkdjzN1ynKTTzWlqS3jvZPKvUxUTGiViFzdotF3vRASrjP4kaeOuzB8mlTWw3FxrbUNzw
0Pt9V7OHo+w+BDmQuWxeyYog2w4tBLx0ig6+F5DFu9MjqTBw/ihjjHOmUi2HxAq0B5NOBRrzC1nh
XV7qLQCCO35eSPBwuB1r4KiRRa0XaBFCr1JfkVjGYaoswU35GkldzGkh0CQn8TscnzQPBMdlCOA6
w1OrOYG/uS0v0m/nNoQTfeUbVoBpjJoF2KZMxcP3K2qRJLGupPmq3pAIKL42VOigjjP5e7Pp/KlP
OJlUce0+ef/Ob5RtUmnGmk8fV9pvFvz/C+Cr7xM9bC6NVVvT+6kO7NdYVjoYaiBhkZcgcSvaxZVh
7jTJyUeQkoxIroo/hmhByHv/mSc6UcUI8GMmMVa2oKyZpGj5HRFojgfOxDpdXVxZIFITR8m5lGGp
Ngi+6TGAJk60r3nE6y8v3+QxT8GwzHk+ruw6hPVIoF9q9vJS4bKGYl/5UOQfKouS7yhmD7KJBaBm
W9pZZr2D6LGVQAxzJt+kfvAdw15ghWGPPzug7fJ0qHHq4bYWY3nTETbzltv1ki4cFkA1GEgczPDf
OOGpz07zII68wglE55OIR77bdyB8nzDeJKeMK6v+DvfQz2nnhbjXaN/9yRalbMEV6kUPVx4fgUDk
X383Frvbn/Yi+uveJJeH6JQEKSLvjYm8s6jnmZbMVfeOmxdDEUTviSxgDmyKKHw5Z1Ub6X/DDmIn
k/Yf+n75h0HINX/RMhoDavGfHnqN1qQyyfrwlTrqQsQ3nC0q7wl0yzu2nM2zEEtwiPklVbualliY
8b5mtIXk3PM1tG2uAY3HXsUep1eEig1VzhKJXqRPoPFiaEx5kIf96Nf18hxA2aIlogsVAS8kPhQG
TOW7IgbwtBqTZy/H1sGmh8qn72U8YeWSbix1F1+pAJ0xPT1h3TyHJxHx5pWBar2C998/t3WQe372
xS8qQ6VaDZK4EnS0kEknhxkjUpMvir8Eul8uq9LUYn2zPA94+ZLNKuvLpeqjKo11luh8OuMReQ3P
kYfkMpEo/qW+08TqfB6yruyJB2CgwFsVscB3wwS+JzO+lkbg3DnQMCRItM0J/F6mBQ8+WvfefxNk
9QLIwLihKic3LZ7jwp5X9xrAshg40wC49c47JX8zyTHpLy5mYvhYGFLL3aL/bbla0M3niZXCwet5
BJJFK8udqiL8O8YJ+0wj3eMCKqvcccP4dhIGA9rQd3BbEOlQB2CeqPkXv0hbQpuxlJco3zTM6AuB
MduRPH23+gwwPZ815mRoWK4ZEEopEAv3l+FFEwfpaRBDyqiSsGeBHkTFBYusE34ZHaVQEU17Kjwg
6elJC9E123HkjtTDf/SETb6KmrdXStP1FGdGS8D8bQKpO4l42N+nip1mUcdHpNNEjgLYxam8Wh7K
qGkzUiYDpcV/J4NLMesSiA43okR6ihBYxtvynyeVHS+/CNXkIy4P1DdNJ/nJbYQKqj2n/1q6qRF9
YntsKjYP8fCKBUTLfDm6iPo6sz0tg2wjPJ9OBcXnXFDIHlpYg32fcsTtGJTZP/5iupIY6EepUPJk
x451+ZFHzcqCa7awzGGjFm0qitepPEvVF0hAv7dbvFNrK0cDPwXV4cCMB87+i/T8Dn1tASVKTN1f
lJ5jeRTLYcbAVR0vbZOrU1G7cpuZLneWCodNj0HLIEt3/oEnPOXcSvsIX2eg+1XhGwzuBluS9ymP
2JeAnLUl7HNs0Cx5l02DRGsX73XbqvBP2h7+W7z7tZ0U1upU4bn4o/8oZXLwm/4+TV/xKoCTiH3w
uYJNH4rgtGAqmImf4Kv8IFR5izdTJBK/9o3x+0ecryN4Ggi1OVDpAs5Kc3q3Sjxgp1bBa4XA4tuI
LHjCrkhS97gN3yUzMcyrGUBhqqXrDxgXFUx02ODSpYbUke+XmWb+8VJZqT3E8illVx48m7dkxvsF
OFfVK4c5maFmBPU1PVpcFQXmsgSfROFX6/MI93vZE50TCQRIO9hlJDPOAe3rQWMR8Khf9WtEEtBg
4IsRN66zgvrAX1eYbsuu/u7qJP31qjTlN+cGMf0THKYJHtegiRnydeikbMij6Us2vPRPiavmLlxJ
VZTTn5955BmviwfoPFf45yBw+siqJVvzZvx5slxuFYNpgcq+K4y5OhGcvc33BL1Wzv4nWYeyM0C6
4qJh0BFxghKIL5kUcLtK6bZlGgh2rm/SG2M+RQJb3wSnxBae2TvI8gl8QWqwCPVZ88e+yCA1is5v
aepFb+JILswXcr4iwH6YrOGW8VOS9UJ2dY46Y2Sfl7C8LFTd22O6B+69RZX/dVazNBh79xxaEjVf
ta5yGEv4agpvHOV90+fqa8d/i0bOIe4LoFaSsBeJvywy7DpoChzvLCsuflWjxHBG95ZWXvCCBO/a
SwCIqBscSJpt9Cygc0QuA1W02KLS89ZdgZqJzbbh6EoaJORp3xyOI2gIfzBfjffZ+qZ5t09DIlHl
kcmlnhy7YSz3E3ukcAKD6Zq1FlEtgKsBOmxzwRiWLU8OSsCpLx8AsBtAYUUGITj2hs3GiZ/EYzwa
DRWY1aP6V1AY5fW1bXcBqa/aPl49dcwnmKd15Pli3mtT8P7p0P1b57QAd6o3lbPGCRyCNPBWXfGG
mK5fficaRPkB3HFq+t17LienM+Acemby4IdOwY73hR3WwfPD7fPzGUPh+leRULk4ROQgBy+86AOE
ca1VBvtcFIJAiklbssKh
`pragma protect end_protected
