`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
cR6QxkesWKcB/joqatTg+ohE00vRVVhiaNj25mZrgpc9TkZkjcUWv3bnM/jDjCZu
WySIJRIjmkG/6ifJmEWqOXw5j+rn1c7yL5jASvcnpHNRk3GDZoc6cqPG6lo69GCP
uTAqm4IzhTWuU9Y+ZUlz3qt/69hksoKyQxj23Bu7Rw8=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 36496), data_block
65jjrVed3kiO1Ys3xBFAsUQpIwL8+LhxOn7U1tjgOA6Q06zqJjqM3nDmtzK5jMxr
dNPXIoT+cxe0pNv2UfJdSQxwUb0+s7KfG/fdLI8Z5HnKW29eQyEua4hBoNr3V4CB
I/IBm+ztg86XhO5/TMaevq0NGeuBqzZToP2LcFN/f0xNblwf2HXG8YbVKLwqN403
w9m80+ZF75j1NDe9Qmj0PUeYW23+Qglud4/Axb3+Da5wJo2cKYi/EIs880H1xH6m
YAuc+i7kQi1FgTIzLHclBRtWC2fQcPkxUB/jEr8jSXcMauDaBIh+VHEDvLy0Pjc8
pFasQ6IsgGzeGPHDolqAaTuh60h0tLNjLtDJYPk/Q4jq1PezvosKwh43D3PkCBuo
uey9XzpY7fUTJd2L9RyGKaGQLRa3THZl/oxyRDiBhe/R8o3hjN0ezZgFAfaUCEjd
s9h/QStVaQ93pXfFGgR3JLC+NhzT3FI8Q7lH9yVjMh5VDT4bDnfR4PNob5AdUT9g
t9p8F94DfB1Om4CgeYbWmKkh/E/LDJ7e639EEfl3oVMOsAwg4r9ItKadASgoD0iE
CVxgZGqyipLyD4pwbf18b9b2K30SqUVTg2m21gHUKrWcZsqhM5lts+v+GSs2jIf6
k3JQs5lmtl4NZAFxnxwqLlw+qG5jJx1AQk3pGZgK0uhKtkP9yzqmkD3khp/qMKnX
TLk353IfK3bgQNUSNi+pUdmST1L9LCgQkgTl9ozG76fPSbnZA75ngFEzf4ucQj+r
TlZeK7nDqG9TwRutQ88uFytSRnf+PHqz4QuQTDMobat5nio32ZOvMJDJzV/AvGMM
Lk51MrU+687iMNvMUJlysHHF0CzOy6OfG2F4E5kl2CLM4WC8SsjESMogbt+BD08E
i9WmGZuIbE4L/x27Tt/vhWy0I6xdboJMglHwcc1l3ZRjGH2n535oeMv5big0WWyG
kURE5qt4mnC95KE9EqQQiG1UTmd3voFsz0J42v9BQUV3kCJMO3d91pLAHwfoFcqx
QvmwsQNwA2+tLRL/jhXKrV+50Un2ag32jbFez8Rp06rShLFA3eYx86lQXf3RdQLu
uDy3WeCH33n3NDM+QW4Ih8l9QbN7pQ8vRPrSzR7i6snfcf8fh5jqoXH1/Wpfjwav
dr/LpLTcGgrUINUpP5ecKuU3mb2sAkTjPrGZln6L8Qfzml2cduNtUyTmPz7ym4sM
nX/gW65JKO52r7TAIKbMW3rT/d+qfTyjmx8Tm+7bHk9V7y0c7LrtrfdXmLWWH7nn
hh4kRMy8NFNqeeNMzpm4Zuh1sMQZXUV4OBKEUNKoi+COM7E0iC/94LMPqidezJA8
96W6OnhXLOhktdBJAn4B37oMeCLImBxm8jknheebYOfMr7nF9MxQ/7t5yMfA8Mhq
z2LtVCtrbUSv+Hhv7UI/GusgTAd9QEF9KYt1CEabT+t3cEkl69v8GxXkKelNYXux
rTKkEOae4+qERxgRLoog7PfEn0DMXseD615HOQO6Wn4b4GOxt4JJEcdaUIFtH41k
L7m0CSPMXVYKVIEC67O42pf5Poefq6oC3en8Y34qcvD7aTcAdfUV4J+Eh5pU+cgW
iEABvdDcOuCDTkCgM3lO5kNCaBqoK8MWSLO/kYQa1O1ZUBK38rL7cA9nNzVPdP7m
v53EywAkxEelNwM0OFQ/VKye8T9b6SeB/m3lpw0msWisqm2ds/utH9O4hRWQA6B1
69/jHuiA6ZX2rf0Q5K7/wdvqx28ata2qAaT++VMhzXQQ/DXiYG3Xa0YkTyJeqVXQ
9DcG4Tkw14kNlO16XugwY9Ci4fmkt7HcDDlmmpaEvdQt+1bQXhG1KJr4H9kG869O
GoeYCDqFN7x63qDXgHZc0QsffJK4DhMEPyPgJiHl+wcO6qqgngncmPzpFZorMkFJ
bDj3vZLUFmFBIcHMvBXmLILr6gVrKHnP0U6vhnbvAkkWbRHQ2ygPuPUXteUXoExe
WufOobqClTLMy2Dtk6ABcgJKvvwusvlUva5dH4srvQ1OTmCL/yI8zSkjv9yEY7V5
kfsPxOwg0K7h8q9+o9LaKfKcKEEviKSl/EczJCCNla3LqTh6kkcJuUbIcWCmF0++
pVCL6AUP9SzyFLsJh/hSFf3ywGlYHIBu3je2BkgNJXD2+4ut3G5HbN5qpx0/7DRt
WOZPnRrqGjSn5hmDkeOTJwuEt9zy7q7AbWEObZKLxdLpPBAZ3lJPO7QXH6M7NQWc
jDTg8fXGLT7L6l8vzShC9xJERRbQhI176sGoA9d7Ng+M2FIhfdcLF6cZZPcPslBB
gszZp3t3xBoMOfXie4BNpnf3MCnCEubn5ygdFLkExrrzL0NLKK1SjzIWT2ZMBC5v
zUlPoF5TizaWhJAH2DRuNiC6xrsaoA88L8JbZZWYc1LAu5367X1+k7sKTJznNvTw
9QdcZM7ladov5UjzmR7y40F7ImVSvZ+l2sghgSExhgqDIXbZqCcw2vvvKsCCm6LY
uni9sMJcN1wCVEZQwtBc7iuMxdqeH6YTij6V5/VvcRvBjiJIrfZmOoSpdVqYbMyk
7U/TWCRSkZoMuf+dAQaf34MNz30zFUtCVguH7xBzctiz1Hkx015wJJ677imxt5Qa
Um1XCtvSakzjgczBP9PykMY5yv8SkUDc/HcqCZewfOKlpbXWWedN15kZ4bxE9aMs
CozidD2WPPykQKqPf8UV1cIkBvfmXsgpsF+Fdf/0TVw9HG7Yq+/jm19tG5rmZbUX
5Hol2EbpGmw4K5nJ7lu1YO+pWbsIPlaoiegeTrZkYzlL3rQPOKzrnnjnKr1A7Av/
ew0F8NIDoP2n7FpW1PYW3+ibv0McNQoLM+YX7JAhuZErd9OjS8NuTOnCvajJbMED
F85Pto8iJtsrgiyqiii5R2AzmjCQ0f54H8LWvg33aU0x5NntHNg339OMfLThcCFe
416ZZYOyyTX/6jng+eCjU2KBo7dcClu0h5+2JRCuZzjKCKggL/P1VKZBLb7YgthM
rQFuLH9wuBQ/0u31VsxcoleWz/A+sHBxk/BTEHU2SC2pnYLtWiWC3aF/1tyc1TXH
gONnl+lMM3Pzz1fYrX0ZgIOK9N/p03ZllTOV7B3/L5W2rSI33r1jTbCpgnle8fih
HCdTbjR3V3h76580mmwhctdL3iyWXtH7kpiGi70X5Ko2OuKhlFe7g3pFo0A3eqR9
TPyv4PHV/WIHgV1FwRdQHXXBCUZzyj1JP7k4xvqbag8lk061hNnJ2EfeMxQeJhH0
Btit97IzHnpE0jxSyWRwpe+FiSPqNzYTeDeVroxVL603BHjyIdS+caSsk6h+9nB8
Ad8L2+3WPbGNpyHDQp9J+agOsNU4WHbNtbre0ivTJqEuXqhFrwyYq5G8RVAk9Q5S
djsMYAqaFoxIyfwKIkVfygIzif/fUa4sJWETzPBwY4rC+Cpc5rLzVxIfO0hR4GH5
eNn5OEd0lWX6F50QiWG+bsuqhjxZHzgOpG+eFO+uTWLqljkdOl4wNoflc0/0MCXH
M/balS+Xu6gmDnoPYqFwY2jXjMT53zJqh4dldecTqvNB/anjsr2JPV/78GLq/l9f
0OAkllj6FWBmM11HKi/XaWWhO4AdSD8MKl1o1mzwdp8+SDspgAmS9q3TMfCYEU0q
yUHiTEX4bbxrrd0lUhOWdxnXT0yrEUWSS9P2QHEo9yM1bYX8pvh14riRgemJgPfT
4cTFlddvGoNYBTB+tXL7aV1GDZC9UXi5ruNlewMLbFgInBodE4olF82kXKKsxTfw
ftkOegfE9LijHl4nii/xeau7YWHa6TqtE5FItQTlsArGTzUU7beon15rDyT1nWMb
9ES5jJL2WSjY3S7gydx0GlYPyGuRbF4lXFRXfoPImRo4xzk0TmBou1ahzQ0IKjYy
CNs8155L8fyFy1/rFe9zaAlcBcIkI09tu6wY4eQlEzS6CwOjdrgJ1/ez4s92orE6
K08ueaurXg0G4uHOvNsLKSBqOn6ePVENb2RnXGOExXJkVUo0kiwbUUibhnc+ZlxW
I7GO6bHEEbDp/SSLeUox+9V+D05NRnHsCxLMGIQBflamuZ9kTsw3SWX9JkJBVUZO
iFI+cc/vRzupVGt8QnbJg+EDl3Rz8EpXbBKbEPoMG4i0acTZ0tUgDxlOk9ryr341
fMDSVQFwhfS4CTDetxHHb4K1jcIUG+2UCkexeRORY+L9iroh0Hpb0c1Mhsoy6IId
4HdbIxa72EzL87RRREo/01No66YPtXWKEAHxIKlmTXKFT5hDsQJpU9uA5nNzIRHK
VvA4VdGTE4sPET/PiLLKzBujIkvAhsW/B32JUWSD5ulz0j53Y8ArbZshYMMzkqag
Zx0M8wGA5xUZLb6ZQCebQb+7EOs6MYuhPJE5FWxLFriBy/iJMSGwrLgloPWPTQyg
o5/TuLbb7mq6BjckNZADcHOlpYxmqBQlvXeMa5VCHV2vD80VECQNFtEKOyWzlZ4D
+GZmatLvsHEFmke8uCp/cEQo1GBa2qUawM99eIVOpgQbVLmTkTTnkH+/RUcfoRuX
U6EoWXU4MlF1qk1chNo/CvR9pmuhNwloO4td5w1u1oM8Q8Lm0anQEoFEUIMZfuVA
dALLFSVwMqbabQRVzvUBUZhw1VtB5swcGOV5KeLQ2cKzQ2RYisqGLyVn2B3Puylm
zAKAAEov5WXBDuAwUFzCAdJu1gpA+rwIiynweQMCOWofKi5tRmz5J7F7BiOrSnCt
MzvlgbRUnHr7z8LhsORfkN7jmIphvrLHXwOazEi8WXIJpK3+d9fvIdKK3ZZPKXIG
XvFpE8MrhyBlaY4ZTCir9A8s9avDpgidYIXeFlUlM8x7ZrFio0FlF0ioRDm7NAvE
pZXCMRYLflqN83OvQqq8ogiEfbt22GJ/N9iLOBsZNqo9H7mJDdfuJS4Hpygqdw0f
qvuZTammeWtbmqp8ImcKqwynNqJcrSokbRuIMuG7dyu9ERvlWdGNBIVqan34ANel
vJ87xQqQi5NDWipDfkZ0N+uvRNGP/+hXgWfgUADTBxjnmAiqh532c11NbaZKHzzZ
1U1HIeiBLrik3Jd9Xz6cVn2ZRO6qW3ooLu68oSxJvd/PBV1eC0JqiXvVCmGCFJOM
JOAZoVHlukVBFNoGabpxQn04KCuIfYuLrab1Y3/dGI81cAd1f+AbQBdpFw063P7T
LR8OlDercGiUCkmonqmD4uj/KtUddQO/v+G9GHoe2C7PrH6vQUAaCWjvNI3Qdg9N
oFDnLhBvjTRvXOaoqe2hHCbDXw5J3Mzb1jyq2rqGIkjvdTMKy7WUmsAVkNmEbtAg
v2iztE3tuTtVdmQWbaVXfpB3Lv/wHSWPxBkjP2bcfGfEcgXVqBccNibENCPFjabG
pyQGi597IM87VgGpIBEazIwLQghQs+vnbnPHJ2urRcZ1+NdQTRCwfTKT72Yno4An
JLAUonv1KayfnSUXtA3T6uBFfkmb2sxQ+kME53LjEihbBwt08YtHOXFBtbEZyYc1
ZLz7UrwatlKgdufkCS6icb+tmdl23L7Le6k7TYo8eenIVuZOXiPTz7JFxK09dhQO
LCgtddqAR2vHbQcuhk4QuMqFrSM81oQ6Ip0vx5Cr8c5il72aCdH6CExwQtnrE5MH
SXo6XAWp9vXxk2CvSjObGwGT0q/324PY4r00avABOV3MJpWApB5SThAn2oVoyI+9
LwGVz9Fa9EiFCz7Le0IWHPaiC8gmU1eYtSfIt6XDvfGTZX64f1SEUV7eRsKdb7n6
+w1mNFH8gT6YpcgVDM9KqW7EoI81PeJwtkU3Gzs2kfTGC7I/qBQkUt+SLwXGgog6
k8pTlwBmOy+yQmV1U7OblzBEkz3XxCKC3SHg/nWnZrna3QIGa0KY8NPyQQpgbD/A
FfGMs0v7yG8tli0C36xJ8wSTGzW6wOfmx5Rmk8V7DwDRIqikKC3gGe+NJ55TG40g
wa8yFSUhimVBsZa3PoBufN22p3c7P7ODIwAgCq5bVMs2HPgyTExg3BobVdvdsgvE
qSiLGqPVqMptECbGsmrD+UlIv0UWCWRBWirC+uHSG0ntE0L4o4T2wxU/O7GrVloz
6UwQ1LoVZM6YJ9ZyEJ73H4fjx4Almtqz8FvCnN+eXRMERLbAjfjJUpaKVD2EzTDh
aBZTJ84a9HSAB/uQBP+idqJkFJNgC8FxRHNFaMUm5/NZKKktFEOYq3WaXcv6Uuu6
laR+1cDuGX/CJwWmfD/TmhgVRINrapSoph8zZbeHGNCNEQE+24viV63iUiwxdMav
Z807hKkahv06XFxCrIGsFDknK7EKJSDgJ8h3DX4dhWXf+2iVtH6h5tOCJAHh6uD/
Wc7NwGeTuxdlyrRlVKLJgA8O+/A8Cj7uPJXlWa5ld73gjG/3y9qTYNLM6FRyAiBq
vr5c2xvwi9ZlC5rvLpvSd1Wms1oIskC1vBUS9g8UtBKu0D1ENpqS9zNE/haTUlOB
Xk+xrsCu/AwICkdsu+mlCmvdrm2FwVZo2Ul8nUuL9wNfaXT0VaI0AvBpdeDeg28a
5/Lpzq5QqsDjhDBxuWwG0BWNdemCcTDa1KsQC+PvIHaVBCkqz1/xH2ZtVrB/uSDL
q5vNYpr3YKLN+cM2wpDmpSvDgfasWs8otY+TpxajBXCDMtb0NLcGd2TJDXdjsy1P
XGGUZRAlxMshXSqa/XxbBV7jHd0gw8RSO74ES5lpSVpJ+lnh0qz802KFk6CqqnIp
JS/GhbI+snKOF4KMOAn8ojksbvqTvwJf2+kplG845LKyOol/TMfnOiT1jqBkYhnv
UeUBEy1cXhr3Ah2E3PGWcqshr/vg7V7lqpXaZW29kdYeYrSmvy3hUuKJ9Y65vRo/
HFEB15O0jD8PpCBCH8OCWZEAoDhrb4gzDW8ehHNL7mPjtmux+PooHOJ41LEAJYby
dr9g5QiNc1TsgOQuAPtFuB7YUbkYTSGlPrJTvd7Fn+5PXjD4+lKNiDErkJVQWuJF
Eo6zbczdlUnHVU+Hgi8DRkao1GT1CrAbBBCEddDKrJs2INHh08/9FruBr+it86H+
S35JIZtUs1ge+ztGXP0mQvMSJfbf+7KsIqKbYGnkswERvgo9ISIH6mVdpGZodKmd
FB5aY3ePvRWOsVtwqYK5fVAhM/DuC9ZsLFmpPeSm5Bhc32TDxwwzzsHlfTEi17IO
CV+rtZlP2wAdhFxup41C2GtTVkNwD7uAgJhr9Vt+cHE0ZQor3xA1hm2PcZ4EBOQk
HKGXLkXBHbdma8v5liCO9G0fIhALD5m9nIl3gq1hjMB3BhTKXw/BouuA/aTLcq98
WrxO8RbmHwmpVsKC9hgVswlQFK0AOTgILHASZ55wzNNNDPaO9RSSkVtA3X2wqVtY
c+tC+uHSY+B695qKxah5cMyVq0vkvJIL/7tEuALv6brB0um+cH9d0W+p4UhbTSps
7COLODZiYM3meTOFCAGg/1YixAMCD73oi2RDGFSZ2xc0LuicN7MQ5yDOdUrJzhGJ
4Q44uXpIDanhh36zFEOtSSYq0a9X9ANfXhZtYEtG4jAO7CK06gH+zWFdlKN4qSfU
nmqWEy/PHGh/502QDLxG+tVdegGG9AzSXFdvxkC+9g0QV68ArZTNnDOvLbRlBEak
2bKjdhuAzqIDfAO5/HxNcpIv/IX1uh/c1vsnbg9H8Yq6G6Ij0A2GwLMpIZpVwske
NLVY2tp+eMHDklncnulsoMf5VF4esKcA6G1biBGDLTzDD4DPwlwf0IFsjAnTru/m
lrCsjE6HrwJdQ/nkfKb65HG/LZFfAXWEm2gY+km78NJFAk5ulghSXCxU4j5YQyxt
Xj522K9TWEIFoMzHm191IMvYY9tJgesgn5DtKrvaSyRguOdtusQTOW0tWAd5YS0Z
as5R8Fk172y766xGY/C8jirSThX+Zg5XyTy3nXtHeDIJn2p2KIRk5cf1WWh41oXe
cT9l6RWw5wUTyBjDkJbAPfgxHZ79+Lw5gFZmu6vkdOngiH+PcQc0huc9ofwqs1mC
qSbXQwjOrB9xhVc7G/nGzReN4jR428AwUIbos9Gw4z069J3cGR+/WmM+RBiGDMA/
3cyn9fNdcOcqyMLxD6RSy+7NM32QYc2oOOX5OnDID/Kswa6rbMPzol5wOxEMSKkF
TKS6hm7k2Jk7Mg+bJw5+qKjAZi+3KzwE9gawkjmVai0hSGiuCX3njEgXkBLl3ruZ
SGdgwsf4OYZ0VeRu3qSyhc7YwaU7iLtzJuUU/EmwOXOnwya6CSxQi0YhE0uYFb22
xmf5p+piDsPIa3Z7BBMg5x6Ote/r8pSkbatg1Q9ES3xN9PEfns4UUWl2pRbkPmh7
58cuIn0fTiZefbZq1dOIf420owUKhq0HK3q+rc46XEBuYPvreaV7Y2GBpUQE7yup
2+1Tl5uD6QrQh9LMVeBTAZ6lXDM6BLkaQwU7QkptY6t7xv/C0ngwtiFEh7SeMp5k
f4Nq7buAWP8ITqfxKOAzYSEPKqzcR6n9G2A6QqbLr5h5LF4nzMc9aGc/RG/rnmmP
BdUag2d/NU70L9MgE7yjYnEXRDtmoKfjttIYfgmjNZpzI15S3juoXaKJKY+2iQWJ
qzeh4LoPwWl18mm+mPcKMUnYhyTTdNJ03WgiM51Kh5ZK3Yx1ka4hiKlrJ7Vn7FpT
sj2NuvE1CUnPik4KzvNlmPptapXgd35qFJ9S6i0tUg/Yjl6iHw3mSd171GLFql6t
ltGVNfyZWpUvsn5zzOUHffmo5ZZpN3QJM53xa47/Y80lvyvM34q/q4KkyK6nPVv9
Auoq95liywWhc/8Kpt864QHO4kSN/eLblf+XQkPYheZ/59vTY7lCVaPcmut8K8pD
k2w8UEtkz6WD5tMhBHgvn3ARUV8RWM4Z6scF4jXzP1Zv+QUf5hrfmwVy5Q19FE6B
1bd/49Lfq1SluxbEyb4Ng2S9/2eUooeFyai/Pml6HrRMj5tcOuwNadY5ybMv1AKZ
LrI/Xsf60AaJ3ms9MsT5+nFSnpqgFlwmCGAFMaH5/L3LepntSmdnteYeudTm+J4e
g10c4ofMBd4qor2puuXVmbnHp2y9GxMljJ3SVEzrr1/JzKMeZDUrE/gH/tPAP7dM
XMKsaGW5WHXumQfRK1ZoyH4bTBINErRA01VFgN/lsFt94B3znKPMLStxLUIaGWBH
HoPQNGDPG+aQz67XEFJ4g4O/aUOBk3Csi83WbAUYn4RIl75bMX8CjnBDyFjWumEF
g3H1bZdpW7PhE4yaeEGK6HTjlmCGHwpJBXbN/kSxPt3qOJlmlaysVFqtBLNfpImA
BGcqP4j26XjjSqQG6/0DsAS0brkHeAuuNiSiMZOCUpZKzP9irH2OZraPcGJlhj7m
FVMqwFFTHuvDbbeK5db21wThq+OmqI38DvJDvV0SeBJYzzNIcMif7STq6jSMHWWF
Bh1t3m4Xdyn5xOmwy8eyR6Qr8gTN5q8Yo10hhgFFuzMSuDWU83Nv7xNL2UUOZhG6
vZvVonHMrkf1TnqPuOHbCeYMGs5xUR7h9p2SQToHdyGe63iEG1h0wJgoKanKOlF2
80knEjCVQwWys5NGxq/i0bxuwjXu5lWZpBdJIbqNpwuE1mZHq5a2mmNeE2hBeqFf
NhlmyV+KOZrW76fxJz5ob66I8pvtcskMydAxffqdXg9aT0yoH9BtoeUNqGDcdTo/
rIgogtutvwjUEJYjUVQ3vLWGuydi47nU0mucMIDs2U8quzRyIrCravuSf+38Sn8O
x+4nMZConEz94m6GqdddssvzuRwO5wW/b/OfppEaKmaSai3v/vMDYnuJnUpGy4cr
YQPiTb4Sqe4nzdVSjMq9fueE20rAYp0S20slAqBqz6J0Oj8/eu1K1KZvPP+t8xgc
HmnMpa7WW9JQzB7cIQL6q7S64+Z3eD4A8bL7dIYJtMgIjUiEmg1qZTLL8O7p7EQc
g6QiHN5IgSuuzq84rcGao3vKcV1asiH+bzfNvepfNrc7Dq6HDfUOR1ZL48Qu0VEI
hFreXMDHob2LK27brnWufUAJZl4OpNIfeU+Cbdj42CPX5fylnywlLsGcw8cyBpu/
epU+t+RnRqdnf/s7pDQO54b3LmfBoSH8s12sTwXHnJ7XGzFNmZ/KFneomIUQFMb4
rAmjzHvDkaLcpXFwQRLZaDX+6ZAoNO+356y+Qvty/IBl8cRCGrE96BDkjolVum5p
hwdKjt26Rku+DGBLELP/NvONLd2qNAoHGgBFFTDID/CNSzyd/JtK0bfu5fgY3gTu
c0NtS00wUQ6SJpZNLsd2nUCnpCwlCi2EmGbMoV2Gv0Bl8EaTA0X9KsMKBfrhA+Ht
2tLeJkTvSQdX5RRhMXw8KUpia2hIOZ/gNmvHZWlW/yq6ktg3QRzy2NLwpG/Ce81n
lOeP1XEE+GUPsNTIgneTbD5a5cobqjRAlJg9RewMU/07SjkyvHbqmr22Db/U/9A3
klkUlv3AM+/4V50GZPyuPly7pfNhEWndlqyVRh/oZ+UK9Xoj53SkG0tAJT9XNC5G
bE7pHwqvawwTeuJsmrDJqntnehrl4secNbspZ6U9G3lh0wmFR+R0K9Aag0LAiplX
Qqn2gIStg5uJBkqz/wWlOSHosI/RJ2ntQ8NdHPWtzDIRgF9N3XhfElPw02ScbRxh
8YE0xkVsnvo0qxzmUnCp4TN6T/oQAc9QXNXCaHfUKyqAy6Wp1Zg5I0Wgm08kQAj3
EoDjxxEqFYsObIXsSlNEIYfV6mMqlwiFRxWwShT9yRTDWJr9U4s0UldZtm8XBHX3
KolM0DwIlbg9NurCzb5sKScAjG4ZZcbSD1/pgpLyB5gzF0IICHoPkzT+/TY4CU8P
1/r4FOImPcUiwUBdZEhFc4tp1c1I0rckT5AYSCF3oV+IvKRUAqx3lhOVpgjT+VAH
bwRtJ5cHdyg0UHdxSeL46EKufu7b3INpAy6Ppv+M4mszhed6wUG8c46hmxO8glZ2
8+qPGqjEnFr5ysMseGfCxrSVRN0+bi608Oo/OJOXl7uWaELe0o68THAi/EliZsfA
xK5Uqi+jEdqsEQvsnZBS59EP4U8s5lMMmnEv9SX89dz2QVfFO6rG1gqN79iTNES6
WpQVFn3a8Y5kxnuX288kYlzK362PO26GkiPQdJpDtAgJXVj88FJqhWwdqfEUX2C7
wIhiXt3iEbe80ZWoSJOF0MamzTEql20DfseM2ny1KytDT65FThA0fgkAgZm9LqUe
1m5G/avl8pb4uICQCdh0OqLXOeq/gJ2WNgXClero1T22B8milkWDqOd1qsG2Rj73
cofLQDaWPFTWtroLLvGl4NPhl2VCk35hnrgSo7v3leoVvnoF1+i7eaQ5HJHXgECp
OXgawYI38uDiqjwHceY6QSWQysBG6b1tBtKFJ7mPFg4bp6hkElKjw0LZD5BBmFXA
vtBHHPDVkUh5jrg20AlHGVymc3KiWLL8jlFhcvdfovDiPTjNhwcGbRxOfOvBaYBt
liTjt3BFL1D86cvLZ7wq/1O5i028Xe5NKR/71L2Ywvbsu3npolzHx8IQhi7svgWa
cUJGJ7kOHrV/sOJQYGssp87tbOtdqVjxcX5PNhGcjS+7CnvNzXWM5J24ufUvE09u
RlZPB53xjMZVu4s16vA5p9UWZzH12hJyoThnPWe+/EZHZ0MtB8Ok3Alm/1N6cMbU
jzCyyuxu2hG7/cJjRsvbIHSizGPsNsv+7Vj5T8GyAmA3OSxc78Jm9R1hkv2hXG92
tS6rZYTFgg4/WCSrxi9H6yMiBfElbu295JLWOBX9gmZGcAQqONz2jSIBTVZUss0t
NxwBPuEpB+7xKzYRKx8+Ts3Kz7cBKhhOhiABHx9ctX7yq6JIAsyyTGgDwvs3mtK4
pi4mJ5ifkTe9cwlTNju9un0AJSo+f+OEWNiHIHsshBRiP2cOzYZNYWe3x2n5MZZ2
ZHGDvxScVdq14sbrpfNXKcqieNcn3NWsZNnXOpNKyMCud+ExiaLq1PaZ2igG5EwD
xm5eudi95a5T2HmlRyEyJkx4T/KhwSy6ly7PAxSTdzHk9bvNJ2xRjYxGhkKuaRpD
0uwaxQOSqKKgCW2FM93kW0rCYsKM+h42bJhgH8IpmysUoYhS2F3q8o4xzgEYp9gd
ehKpqJeGPTxVt/c+e7I2EZa1R2omJqqK4bK73lmMhq2oJQsr4gS84tI1Dld1Jxuj
wF/FEq4adk7IYIvrt43PkvG+KsLADeTDuTcFlS5Pr1SU8qXe81U5jSySY4MN+ekA
YgtIR9NygbIPITTnxiw72RnIgKFDYUpWLoEeVO8ihWo2e44p5q4g9pDx3Y01mzR+
KglJkcmrZ11LYadPFFxqOFLgws7ZhY1FHlDIBf0sL6RlJcqwiW3BpzmF6CYKVXiY
hgr5dUTDhn5Zp7Fj+4c7/GwvRetNKiZbcJ2VggRhb53ov1phtBzT1361835QTCRe
65Jr7y36LcEL/GcqMqZZVho3uIEOu+yBxaQQQjAvzMdsrY5QjqtP++++lxQd+Iel
hnQdi0YA+4ukOUL5S0zlzjUfFSJ9aw74F42Mi/oIlJhDaAOODer9CAnzLHI2T7mb
/KbqCGWt6DBAJV9RzpPvFR3yZ8beGL/42Cn3WGcwpvIUJM5mpYDMWBkUGIK2NG+A
jnQB/KKWPE3VqobdGfaCXpl8TL8ktdT8GD8ePXALA6OL/3TKkChg1nfIM0iaQtf7
4TWR0FPO22iZLZy0pN+yu1Oqccj//lz1iqmzQOZ7l3GhymcXgTrTo9Fi7fvhJxnz
m3mUb9hSe3RkcXRNbU5fQHr8ylXGqx3YcrguXrI9kUNz5fwChJvL+NRMPPVp+IDC
EKp3iws3ckZIg5LBoSiqcZkmW15f+XOdiZJy6xRrMbogHCjCYDPo3KSEQ+sbJL0T
z87qsgkrQN/jWbusSrVLws1op72j1GFrpMxhcmZkAKG67Nbl5+15bukoQ6plMbFf
gg7B8XXEXE3kcErG4qcnJ2+Q1wkJWl51s5a4eutSii9FD5Huk/vLqaywM44TrAlC
q1ULq2U8lYmf8XTR6O+Qa+wEvPw29hs3mJhME9YNnRmWLM1za7WQREBngUXNtuIO
W0gvFSn175aYlWaM2GQ47+wof4cbAMX9Lt/+lNfqFNjezG3Iftw4SZ3IzWAwO/do
An39kI4GM0W8OqUEkzPd1NPerYxuzGUx8kydgyoS4TERhLl0DoO5+0fCrxSNoIlw
PPB4sWlmJVUTWlwaNamcS0I7yPHExyOY6j13Hmco+XB/fk8dO7LFgLZF8Wk4Raqk
uOEJ9cr41dyrw3vJ4MWCXJRJm+YN0wIhDfhUljFcZVaZ7/lelMrW92qAvoX/R9zn
F5Gl9az6pbAG/ElvJ9FzD/l6uSoWnekoUBKfy8HIpG9KBhvyeRUys3isXH6XNKMQ
i9OCpITbLz5UkasStNw6Qu9BBQ8ZqG/ILr+5bpOIT7rOTzVOPAvNOyYj4ss7xUCY
lhiIJ1H411PZgY4Pj0OZgNxNI9i8SY7HlKth0uwvNc9Pn1QTsHRdjJiKS6guwm+E
atPvreS70CqpMImsSB4kbBlIknIfE6NOmZdrALe2/lCakxfgwMJg1DCiaK/FastB
Vhsn3FuEGAXw2z6wRQJLaOo2dzMz2ifMTVHiLmu/D7ZW8Q5eOxphmfRjsFu0+cf5
oWSNYfnYyT4wdN6PLkQssEIE3mSUYKqKYb7rHoSRTU0WHSUPa2qFcq7PpRU1pFCT
7fjE2xE7h9JzjaBSFqIGCMhH+sMJJObaducC9m0+fS/0GO7eP1lkAVPk3JO9rjue
ZtqFpGPHm/G/2RLyib0RME8w1EKfS5j2e5c1bX5N4tzzQLobeWgCEnYV+5GBoviV
B8IOHeEtGwpF7iN6YVapQeuv8l+Xh36Ga9SyBQXhIJrp2JzwIS6a4J3XcHatvcba
htjno6pCixk9Lpws98x1Neht3XdRGSoqcz91xWzUGvYkpMpji8INVnZmZaAQIzGV
AKV9pAtaL95tQY4qDpHrSX2sV4kLK+EIuXj72jdlgmgMdvbOzBg/UUfTwFMet95i
Bg6+2adJVoJFEDIC0hc2qtqhf5TswPHN3Kjq4T5cySgBhl7Is2DiQve8MfFZl0IO
uwL3QNX+c0MmhpOI5zrR4hKahFJtEwpEShvmSVUvbDOiDjD9XCx+4HieRxeoWMEX
QFMF47V+vhXV/QfyRhh8OovoPTY9l1NXJgTmQP2oCrlUEdMvsFbpuBte97XDSzqM
zMFomXnl0MFBFscLzTbeFOtUt1nqBu+wPpdgMLX4NBf2ooT/HjsaYFnvZIbSjBQj
rbXO5cItYf7oodvtY+UGFBKqt/LPFRrNze4rLiq31sxp9iFSl/urOU37S4ZkvJ6b
EdyoLqR2m0658IhsWl9nz6B/Pfda2y8YToh4eleTMG/+JQO1G05DIzCr5I8jlgIr
9em5U/O9TKhqspBz8x5Q+vU6I9lr0jNWANqcNzJ/mKCVAmWVB9xRS92Ug+OLCChU
0WmBrDrJavVaQdvH+796xPywB3ak0yBTrVvhaiQ+/M+SSRDHSYFWElzSDhcpT7m7
Fxhajhp5r1F8VdAxd9R+3Ln7BtwWQCGpkYMQ0c6jHZgVKZ5x2mTo3kKTBZf0bbo8
FGOCBbO+jhXEmXU+CzEbScFJE1hOZi1WdwNIVRqQMybN+j3+4BbBey0kazmz9hbm
p1ir0Uik7LQoESEBx/CsX9oIn3LyjMKaMMBRAcLxGSmdQge24GRrgnY3hCsI+fag
fFOLH0I/hPMX281+zSm7VXjLElze/Jsh9k7CQOG306u7x81rn+F4w8Wl1AlRqEll
yKXvz76R8fJtZGmryEIUG0gjNSlvkVQGKodDTDgRDjfyL4yTc27G/+2Y2e2ghCSt
UM71NjHf8Bc3s87rhdu0Pop80C1ILvkIpuZUQIq+7x1j/H8o2secxppcccjqrF9D
ARl1zOzlVh+JdHd59HpY6OdEuA6J5HM689uixs4YxUtHC7fhtssYmIb35kUonZhH
87GuBzqWJBlqB2tMyXODmEQvEwV2t/6GD1W8izWP3l+gMQuNuFC4prTplzIFJH1j
uIspN3kSD8B1kFhmuaCgnZcIDQc+/ThxhkCt67AdvnvnS52Nk/ErTApMShL7yqZu
NahUyUVoQS2TvLa1qTA2SxFqD8U13/WXE1bgvmCxydFW2Ra/Q9QHLEjRcxthuA/1
6a9okJ/zVjmA5xPsLc01MtSyyeJCrBBeI/pudO4fZtGjrYMEApnLpTp5VSSdj43I
aSW8jzA/AMmpR0rXSveH2zGzy3hzDb+F1UEhXfV8u23eLmEkFTCAe8nTFilAf/64
BODxPzKfgvA1XgE6AEY/H3Yfn0gZOWAUZMmF+q6POYdEJ1DVUNqvC6kLwyjHGDIo
lZpijH6f6fYOavP/a7DoIsMqRfelxViz9dB4Fk7Pcz/8jvSl5p6UiWapLw5Fyuy5
1lflhj7K69zR0/u3jZL01wUTFg3YZ9ADiQn2B59vKyYdVOweyGRGLyfOxrqv3KZc
W3agkTU8bHaamSyXMi4ZbI3vVPwE8jDqRn2CaBTahK2839mImB7S9oN6HQPP93xO
juDdW7uOQtui/GQaGltZqI9pPvUvxMa/ywv6RnUZg0/1sO25nUl56RwBzJRfmfka
szeXlgE06CKhhaqEMtLWeCApVVnIfN1QewsFeBuuALnFHnveaP6p6Z1bCqeTdSpf
agenwo3v2UTwGxGUiHNsyYUw3yoUbR8HHxG9tbQAi9WkddJUDrqvIm5eEBN3NMtx
vHOQBnH3mn31ns34Hjf34g3wj0dUYweVI1uWOBg0PwjXlgn4+UWYqyVWMaMbf0xT
mlzylFEDwue+CewBh9GIH1vC6Ig7Kad7rC2ek2P/bpEm537GtbqW2IUziJ0VF5hW
U/vAP+/gGEE7JCDMcBLJKZHd+IXBYJFmijSM/F4QolgNaSLKR1/1OI7tMfTiidx4
Uecn0kXf8EbmZZTnoVNnVKSHJYo9ADZf8nslerug6qVluih4MlIxWNRoROI1Z5Qc
Czeoj8rnrz1rwQTRzPT7ESmEJkNBOcXS9cbyCLsxkZ97n5kk4w/YmfAPPXMTtOad
hp3D0qCk9aujWesdrAhR3s5v4VASPl1Kjz8fGuQj7bSpCUg3uvvui3OAwcJQg8cV
hSdFQFHGAyaWwAmSjLmngSVvGRdV07t5qOila+UA97QW/faDJ498ANS1oy3MHXxU
JeZ9ZOe20ATwPDBaoMgml/3IRFAoXMC2Ysyku9CrXrQMoO/Xt1iW9bgKw9HpkYAo
yLYA/ycgv9jcb+BRZkJjDyQLvDIpm3NigdZKFoHMDMC1q0eCOeOg441d2VHDFACt
+35k93AUGxK4khv+0GzZfTAAyBBwdeEQU/2mMcT6lmdaI+WT77EQqPhhBSmeFdz0
D+sTBCOAWy4YuFF9KHdcgesLaY88aKUz5PWIzKYyCA8G9Sfy4Kbg2hP2FYFQPzVX
Dz+nOyIgc0yZfZD8SoCYqMrGpm0eSBICqITvo1ouRG7n31PYDh82Vj6T+aJrMYd/
x4YvS6qO3obOcxJ0WDxnN98vHIugE01DV9twQmCbeqwM6n65GRIWZQSzw5WAZ5/K
d86mnW4Kb7hAwG6BJ71EeZ5so6HC5NK5bmkStmvMMGhMkhM4ar25qXzbDsXZXZCp
tisteglEpgdbX6rRs9S3EuoD8YM3z+NtupHxD/TTVynnG4xc60cw4Ernq/k3kvrD
xVb9cFtvWxhYgxc/LjqxvigKrs0RhekdO8ydKBrqTknIOR5nrDnvJqxf1tB3/u2/
uj5O0SH9a3z/h4ueqpNQ+mpQuCUgTSYm5qw8vigPKDwJOb1LDC7P/8itO3U1zMP1
fiXlPwqBg4EFYzReQBvxuMdlQMUxir6/4fLZO1IHrNdwL6nl60QGadK44UhVC1hl
vzb1aISVO7l8qpvtfkZ66RSviwzNgW/7WAFpqiyp37XwJBazkawp0Ry9UDWbZQ1i
zfWuj8+croXSObIVb/JJkINBVe8I55IUBPGqwuqBUGpqXJFrE/TtSNV0unnwk+oD
HjfyNwmcpcx2qrNSQ4THKq+Ygc94qdOCqw3zxsUPWIP7VgnwA90uDJXideZlrNTu
10Q3it0Lbd71uqP53WvEFUQqFbdZwrme32GiTkzJn7L3ZqUUwpJkt53tSKQ6mLZU
CTurin39j5JgY8ewNmqr4bU7m42Lp3I9GARfcMcXPRmYolgkJZTo+oeQjhNggtD6
dXZrsEcR5Cwt01YhLj6IZ17fiMf6UkaLoj8RnOBXdcX35POZDtBs8hKSQzNrKug3
bRYWpmrrITZFpnAXVvK9+ezGn+UIIrFcZGBMF8j6GNHSCsHMAKDGT5iRAjDr9FEw
KZVPrCivhQEj1SfWrGkQeMovBKIHQgFwnxoJ58GnmMBK2hKIS+Gt3JUyd+hisog1
M03hl55M/Vzwvxn7FdYa557TRKC1g5tV2DH1wJT7KWW1CZ5QMz7eCfpwIVz+WpEn
K2xVvlnvan5mmrCnCuJtmKIGW5H+zZsO6ADGLokahg/s/Ac/bQYOJ1u2CZJU31uH
yV1fvfUu94o9JF0WEdaLpwmf4mXXgVWHxO6+yZaFNd0lQzH3LouvL9G+b2NZ0sjn
U+eIUpCD+oH0eO5097slyNrGlEu0BgTX9fx+gNi39CwPrMUmBjN5YDCgmX0lIG9d
kmWsAJTNdpyKYVLG+EgGr2bLIASHoMUbVUPtMWpTIppvjtX4lc2RxmHNcKyaOCHe
IVPp+eOCHj78h6C13iqq/habwWQMzva1C0JItDekrZ9n8/jh/jt0I5l4aZc6eCXP
BW51DUgeRnGy+A/1jAW5DMLNUYq5TSIu96cRLChQKkaCf9q9SscxcLQSs4ZcQG8O
T79YBG+kNEfNUlLO8aowDq0FN2eu4/dXn97VAQl4AtLvdB9DZC6zV+rx4mXRXL9a
2SRn+7vJ0zKiYoGbrX/A3BGwxX7E6yFHhdIsskOfOM4BARKt/Yov5kuQOjBFxESc
b7kAlHITIlyK1ryOfapHb8dS4aAXixIiYqmztbzzuWiEy7PufBiXBCY/SQALka1n
1hL8RRdHFEtNGk0JbhEohhSHPRrbDKdWgv89/qCflv/Wa8oiyWA6XwKt6Z7JP8YS
CdI+ws9FT5vySP0u/01tRpn9LMakBqwq66DrDeCet/pbljiBCTISEOFfLsyCo7a4
26Kz5QfYb1ataAXscKwiGp9ERNhrD83O1p6jlBzrE3nJaR25rd6TkdQcaS5tv2ii
cVc/0vDvIlmGhnmXBU5bPT4D1TTE49V7Hgg8ZjQJUTPb8phRNoVRXui2UbNmJaBb
RkEfpbIgl0W6D1/lj4IPvZQm115zP+ichXDqhGYp9/QaR5mSQFkHd/lcGjtna4g7
99YZKIAdacZiL455mpmbCsY32CPys3dFIcIsDnBdO89SIU23CCw3Pcwg1U+I3Ld/
XeTvr1YOugS6hAHxMrvFU+IGJgr3iFt7dHGX4SIPnjzR4K0E+C8KbuJ5Lb0/LedT
hOyMzc2Qqsdb14ZJWqT8t8ZJhYpkTX1n7TH4wuvZimanLh+bsxaRJzV/WobNrbZt
KW+wTAQlGkHqSFnb1D8vvBOZ/z9qoyyorCwtSyLbTcc3MmZXVzwWubF/gFyNTbIE
ggDZHCHKt1/4xgspwFuYrzzeUqcswZCJ9g4gzcvOfh31iz7fXkTIITIp1s5GpleY
z2M6tMT8mqApTSeezQpEw9yyI25FZYo5M0o9W2Ctvt87b2QT78iJbYoKq6o8a6Pd
Xx7O61Z6UrOzcoqNlkJg6jsiV/Dbr4W9YkxCsURwq2PjkCyDBnyNCrNpLfzeHZQ4
QnCFOXES4BJ3CWw2s08e+aJLm5ODcI8xBZF21kuIG+ytcvuL09AlnCKFXsWIoAD4
GEfGNfyCbeWQCseHHmpSqwoqzIzPH4ig1Jxn+SzgW41RhC/oh5FTRzXg6h274ERA
wAse7iBpIq6guF0186h4aMzMkoWGJC5fp7Ij2n9Wg34iI1wRdJqZ36mxIclm12/P
/4CpvjpQAMyefE7vsMouMAWFWjrOKvCU3TdZTcVK56BKa0QX0sv02oI6qVh9Blsj
Sy+HVBG/RlYY5/oTvMB443L3U/0Ik0Kii3oFlTu3quXRLtx6+mqOxbewyLFT2F9a
ZfVE2sOcVZ8A+Vzkldl/gbR7FqWikKTwu0eukAEoluu0SmvTcyUsMaKQlI+bsHyf
uZRGTJJgyJOtvd2GlZkjZzueL3JCvcHE8bBh5uOBfyDSAAB5vTCWCOddSz/AyOZM
7yGwJDITvaQM72hiIzHMTnqqXmJ9zNyuw0cXHUs3sc6JeHTD1Nl3jY6u44YHdo7d
i0hGsFDvtuxLmddD6dxqogRcA/z4HkUGIfd2dF7qgubC62yiwIDxKmLGiXcPRrzT
CuYAaTOv+29Ojx+ouEgIzDg7qjFQibeoKrnl32z1/jaGdGMWUIyOsxdZQ+IhOS6i
S/Ll9ehZTb3r+08Wq3iX0PFSGMPsaB3MeO2KG7Up6bOiZP2P7QSnUDmI0Oiy2IP7
tNB3tLfg3tPzynpYGrICwTpwGQuYS2qc439RkFgW051mj1LNQhc7pU3VhbFA5jCy
tcjK8N4X+j5B4M60If2qfavgrl/eR+OvzFEKICrCMA950Qq6H76opaS1Y+YrtlSL
P4gJo+GMvRM3Nt0q6HUvOCnMm91QCL9HDf27e6n7dpttmJM/cbE3yBZJicjQjrJz
sFUcNbb80VzDsY3lEYY9VHmdyIPP2V2KQb+PGO4sfXNpoEus9XJJVDS/xwgsx4Lj
HDOY3YUb5vPh60gjhCJsULzk8+MV/tWl3Yk646cS57NHz7lAiEStUL7gwTrmq7Iu
2QvADnfAjdVNayOcp9ddvS/mDRZZLKWuG1xKSrn8vw2Fq56+SXd4MWvaq/qNgU0e
bMHBndoSj0/WccD8gplHhQ4yBk66HWUx3YvIKvPH72WS1Iy+OVMi9IYNpLJ5Kf0j
BmvuL2EGpgAsS9CwX0YXX5NABECfkm+KaJ3kiYtlv9IsF1c5uK8eSHRba0JLe7YL
sAyR6/TQRZMVVtAWfczQKcoFR6YV8OD2DUp2fn1nkqQLFliuzse9Mcq3rd1hHU+Q
r1K3tD8ih1Ld3sJxl06+CVB26HJKnAemuH1HQjzUKpQVWpyHtX0qtAqjV5CxJPMj
2b4RU7S6NKt1vtD5kBsaJVpfIy/H7BezvNgGNjPAcrEhaW6+og2I8T5iB2K3n081
ab7ZInP3k4K3USFE7bGGA2R2B1t7uDbhyi5R5nKS9wALrXVqJ2LRSVVUXD70xwgT
7nn0YdcbVUdQFCbH5r0hNRISvtnTzBtOwvGUfQ+WKvr7YTPKBCQpj+chcgHybDaQ
UlMnTZZ08XjtN3Qb9eLEe8HjsoClww/+Rwp2J4Q/OWlJAfhCKRnKdVupgsigdY8s
Oy9hwTFDnXV4tL1BDrau6FvmWl5OCfLVVPT/5UgB8SBqwgzisCOuCUt8Yyee6jdD
sgpzmiD0Y3ICZU3mKp+Sz/h09tZqrE/Qv1+zaJ7H01ShGmHMoixRmf3DX1wb1mSR
PGqEyxTdWcq4NwZAYwlZ0em6Kz713l7MiRQNYfx1pPQuj20qlz7sjBI1+1kO9n7h
Ji6A52s2+0IQ7vdS9de9Xdeb6AdqhCwF9NcP4oGLnmCifQaQL7bRgOKLxMFW2ibb
bR5gxvUVIbTU1ZQFZSsx3v2+67HSmg9glRciMAxerXeHf2CN9tPgp8YUorQxtrti
CdDiS27uGD4sDk4HQQgEmTiS6/Ke99/dXthAtQkri/Np7YMqGG5pKyUTEBVcYx40
fmGuuGTZNe10uxDLQHfcXKbRlUW42Qtfzjl1fCDLPM9k2xVxxOlpaChPae+/kFfc
7b9dSone5xgAx2TCLRD5mvqjkd+TmoEBqOJVUT5iwfo+QFMVccxvcNVrJmFJi+bE
sSKNTnBmhMLv4rRKzQO6ObqbRHBJNhxHSC5RMRbiGlGNONRBVb4P9jmiLNVJL+mT
3rsCOEHvzEYob+nTOVo8/RGeFq0N56qWsAOAk+7OjzzII69FHKC2SI4YVcyf1+TH
upy1rguRTnRMy3S7taFaOcEGrPjY9Za4ogcWn1f+gPHcZjyd/EFUlSezzAnF/sqL
hTXusyFTQOJfGTWW70mLLMd5Qsn8X6wuZiVpWz8LBJ8OooZWg+FnXBRmVAOk5TMy
osNpkIW6BLDyKGiPHUrg9KkDZJITZ8TTwBAzYmUU4tE4BbAcijBxDqoJP8WXXgl9
coeNmhuKAHQjq6v6hpxeMC7pBJrzM9zi8mBjUXvi7ExC8g8sdIECRt3Rs6oAY9yV
vpViELugh/zUvZnBTogLcpZsgnkgB9CvCIpBsu6xd8F7hT0rF3B+/6f2lmmkCZRM
YLG/ww0RbaDasTygqeHAG03w6fL51BeNELEtF5q+lpB3TqGMBC34vrIZgNshrXL5
zUsZDzAJX9GrkqLhg61V283f3Yr/cK/1kAmc0eWAyoiTvvxHa0FDRiwAwWjZLCmZ
Dp93Mylkt0CIASmYQFGVAtuRnN7M25EJyWkrYf5X0VoVnIWEy/YQIouvV0xokugz
iHILac9urA61wtWTG8XaW2nJUmgbNTdNl8HNSDWE2CN216OZMsJHjRLrgwRZVibM
6i+PLH2U1KoVxgP3hCRsKGLF6zEyEazkdU1YJ8A2JvN5g/dQ9MxATqNldhgRV0Cl
fHZJXDTLWpKS/7L8Jswye0aHefAOvbhw1nVng0TwrGNuk9DZW2/oXK6fr2Gh67h8
hy8B9dIZ3vd9HEhfhTA2t4Nf0fR9H27LXyhj7kBK0BaDavanZW/msPoiPqVqKpSo
+wa2whlg1hTVli+f3jV67AnF6IHmz9VyO/D3rM0huJO+ldDh5sDGbBbge8X2hK6/
GDdfHmFeNkuykNBCCGJyW49AzjQmU0UYhpsizSRpu9JlLPkkaXV/GKwfAX9mwZpg
Bji3IhW7k45zHCutUhClH3YD/vJmn1+A57L3kKvrbaEW1v+oAarc7qoB2kPLhUxh
q7eipfImKWlf9wwcI5C7Vt0CsOBYzepuZGlgFde0Hf9oa06+6BvEnRbjLJuSgljM
n4lUfF+7OxRgvOnJLorJHd4rwI8knu3wlKgli9834frJNhclx4m47ugGaPSoflyM
12R5LtCh7AVlBGkvm2kRXm9ygRG3/g5rel6G5UjAtPOK0zvPCYNQRee9fcvbhPWM
USHxvdA13Ov0bfaPuO7cR6xuA1MnD5axjdw5d9rXbeMOZhd+gxJSrOyfgo1OfvtZ
ocH10VEMoz8ziMGmXkmWnXj81yqEz4l6w30U2jyFxqrOZgHW94Ayok1tL1AV6PJT
iEk7ubYob5bR+RPJXzA7V4aRb/IGzV6vKxz96CFWWyo26Qs3i8BmzbNIfMryrAZP
/Uaw761k7XuewAAs3vwmwb6sGZMKg//nZW2xPfeLxHLttlF39dMfZOzrVJMhd4bt
cEgr4L8J3bkdZFCasVtTCtKxMY0KTqgQC/Q/hJotsx9luGOtuwmedsTy/dLGbPhb
C6K0kdiuzNsNp6XXgFq6k7cjWEzP3i7xpJ1dpqzCTqQjOlxBY4gmIKTttP+Bytw6
plJm19hLOPR4o0DOR12KSaQpvi+ZgShnNl7ahHRUJjfhyhnk0ZDuaNI3IrJII58w
yRgprW/bssUetfeIp1nqB6c5dzNg5dSPAmTYJqwLsFQ+quKJPVNYXUtEg4yTzRg/
IO4Rq4ervIHjy4jn+qCHo/6bfSX9pDpp90edGhJazM6MUKzGTJOXZf7kLPdlTgz4
k8UcoM2ePvWGPjrSnr+xbVwZuYA6lmBXUbkj3mkWAmbzAU2PCAQzNtcQBOBYNCr8
ynO8txQWMbTyMp/rqEqrNLG05S+IsPpm11PfKx76HktBiUMUjljyjDaZZnIESEhP
YnT4hRAZ9h+AFn3sWAzDcUH0lbdIcQwEJFJNcr7ecG9PEo1sd2clqOCaGuvY6IDp
TF5Bny8dVhhq5b232AkXEC67R5TKEMarpQCieGUSz8xJRgyFD2HLqvBwEpevaUbh
ToDjxJSrtG4f7N345YUSRfpySi1xKzOadPXLxj0yqi7e01x4mNS+5vHhSWi/QvvO
l2aayQbX4SPYb/5ANX8fNkFt+uBPVExYLIYxUQi87EV+zRtWK9KMpeVkHslPd5Pg
dAZqLEclueava9JE0nyboJP0P1qYLVMyBOJrpUB30T1Eh3GDpDCGf12a44aLvF7S
d71vu4wQglohEWFcDk72w2uvogHsPeVcqQ1cMMcERFtHU5tKcV+SyksrzGIJgWUK
urGRUEve3G8zw4ThUvV5x6kewFxdLEbW15UleMWO3QY4ddApTCo58l2YHR9VBh4K
mfPONB37liFbfIt5Qkzvuk5QUTUe3cFia8cboNu0AvrBFec96jbwra1XtnZ/7/Yd
0WTxZjQiK27OCrAGtNRbMgvPxlow6/9jfUfVpN+5L31OY/uJTxno8+MT18KPaOmw
TDCT9CDLKNln0kNZMfS4u4b4o9N8Gd5HM3hepAwDh/DUnfK2Y3S+MH8Jen+Nj06n
AIG0gizmdrmJVDMtG1EN+jGPog+FJtO1RGG6JTaS4Heruk+TMCfjrFu1xzUhNdBW
/7m4xfEHLumsISu5W1ypTy8RFMXfC3WLrLq3E3zI1LmO4RI77yczXMZrLrnmnZhE
4/C976rakb5ElYzigMR9b2c6Q5yFlGoZnZ7CMcUmQJ9Z7keue//VTHm3VhP+YcIU
URHu7kaW0eoZfAZ8izS8/3q9hYmtdHwFfZ2l+ia0YlJGjSjgOZ7E0DH078kLe3Pm
+8r/dOVBKS6f3EqvbhhbOG2zzA1rQdcQfpX8V/V2ALBPwyZv4Seob3RoLxulrXOx
nbDcvFWVZSL/OysG07yKRMNCG3YQRlmseHGiFLG0lQzQQ7yYxaT/rH0IDqg1Vtvj
ga5+cPDnjLdwPp1er5f/IFxo6GKbTSB7g9vDmERBZGOet4M4wGwdY+PZS+tSLY3t
pEkaxp69b/KNklnIMNOOMX7JqW4dHl0Ip/FuzShhkNg/9m61WUUB41Pl+HFL7kAa
zfu0ZFDcdD/gSiVZPcGEOfvdtf1AHMQoCthgltBKChrMmBFUwC8jcd9c9K2OMvDi
JUeIL3mmiV8viIn+x+iGhPYwgWJgEVTNbBcJAFDuHO/+tvMg3CLAzfY/8ie7xAEg
euJWUr89EXKiTn8iZI8jIp0qO7t0jadEr7qPlXacV9w6aRh4hGdwwpMXtd4FqxtW
Ekb3xkSGFB+weiPPTUGYPNXCu46a2Nu2T3SpPEwkWAtpabe6+dhFRYqxc5zQZwRB
tc23KLmBvq4ldZqxa+9DbGVJKORGwH52evTSTdHbl4Cutaz2/PXamsxKL51272bT
mZ2dcLRB1rmY03Mgm4QZaPZv5CpzeBM9ZTFRd42shKYj74sonBmvg1956Y6gRCIh
zIDvxQY0PNbt4Jpf1/HlrxnmDOzqxFdsZmW36bMIF09XAY24FcADkiP4dKIVQhY9
T3vO+9rv7IXdYIqta8LiIIFdwPeIsURLKREim0NIWLtXq43ggzGLPBPM8UI27qYb
qiO5vUJse5rjQpfIrNiRhlA7HL32NBhVT3ewk4N0z01wZaZjO0avusFzQ1I+H42a
vMWN6bvdgDBqn1MeaJih+KB3joZoXUsy0d2Sgq6h/5RyvUjgQv8uHtHk5aeiEuc6
DNzFK9AeOQVHkQ8n06alBG5/tgFKVEzGAdv2ZFd7wv2bvN31yhvUytZoFnixZm9h
eT1a7dInxgwaKDWttOkV6YHTUCrVW9+4hNRjprnamkjEZpjpUcz28RKgFe/LIUjd
13unEwooumweYDcBBZD38fyAwkR2bfFsMvDY27v7lHir7l8c/jC8knY+wl9h/69W
Iy5Gk18ShumRhYIqC/vMg58SmsUKTJJrSh4sfAOtRuySNmthARaTeVrrcT+yMDdC
w3INtRIpkRlfTzmXWMsqvc8eJkfzI+mBc0q8k9O7jdwWUln/kbgrLrUIVa26DS8v
talOW/gQq5vIVs4yagx+7J/AhwFIk6xXlAHizd9eeWOWrhM43M/WgkDaEeEoF/2I
1U5egKWJu5F6N57+C8kvjCXj7tHqQbbQnsOvlg6DJcZ01yALIn0EjSpfOeoRWNTT
aY2dDA5a2dLUAaKXLZ64AJVa7ZDYzul0NUmVysO1GFW+w0njgbui0Y51T/jpK3g6
V12Q6jzsNiAOnPetTOL9vxuWiOPgL4B+MSydf2GQqxpbYwSEh5XDsqenwEGNSCi2
leAGSZQhyTyd4WW8yEoncSQn7+GrP3mNJbcAXoxalpEi/fB+H0fy9rSYskvjtXbP
yp5r65aS17gHPZRIz+rjXcmvQLSvNms3Ab8zZTB2V8/hCtcifwH4n6LFxZPRFR8H
Y91i6KA+06b8pMulqMV9cwJfcPunin89P+tqrDUWhv4o7gEPY2jZSi+/P+pW5ytM
aV90vbqNH+6ldvbZb2whzKbX9m/BfbwMInORY+ivsnmQ8WlFe68Kso91PDEB7O3N
lYfFOSnuS326KpS5oqL8AwTWExiYmut0XpbH2MQUFZw35oCIuStrbdYFeUADpX9P
D+1DLuN0nJ6evrvnQ5MgKsfo2WPMY5Hn0yTiQwGUK6RD7tY+pK2VeKABh+c/2tgZ
GKxyrCA3BjGTzN8P//7trD+wAtwY4//n5sbtuMKjyntuURH8/cZFa3a8AUMIiECq
EXQT0a7D17VqYqcog5IH+/yxb3a2MVCYct6vUZYBX0eO3G2UbtjU82x0itn2BQ6h
bDCrIlthE1ryh27uNnt7US4y5JwY/5xL1YFSP8M+aDwQWWCxEqoQ1gbLjngLlomd
6NhNKzLcSuCsMBDLyy7itOTsYCsgijAE7C5wl2RjXuVrhxbVxSss1i9U38xYzsft
tqgeTZsTq9psvINWVFtA4tLCdJELmOy8IchocL71krCzBOWZwmUIVTfoshuhbXDU
3vXhIwR38EQyqBeKtxvYDP/zYf6eQZBfuEsj0CHrjqncSv0xHZ2RpaJU3ZF1s4dY
cfgzm48B8DsN+/imxoVfQIYoBGu9cGXA8ETedASDxBukjqrMuIrVGJrNgQF4Kc8V
t59ykJrSq7Vw8P5KnB/+/fD0mum6s4+Rjimgaqml16UnGM7DrpxTSKhEkIgvSmbb
EtQYVSmmAWZ43d9xVxIfl/f0v7RR1vQwyNRlgQOSEYG7pAI+c6i55l5DnUlRq/ZK
v4DHqB4RkpQuXpQsH0xJVrlGhixOzS+3XYAah5VJbpEdzqIzi6uyGwFgSUtnG4Gt
DF/AH47v7fqLNEZxNPh2DCXVnTWCsoSI31GGNswAiL0HEyJcnwq7Rge/uhqRwHln
Uei0MlIDq55CHAw8KLt+ZMO0rS0mJ9CDgeDLvST1GwgwTmvcCVu+O/wV1t6/ibWV
xqUnNZIMX9sYLrLKBel1gSg04jviQwViEcKIKJdo+8230L0n6K4E5fGX0f1uYyYy
Yr4shZcQ5/qEcjIRMpKVPIiBxVn3Z7uCId+08PYbCONlgpuxQ2K6Wqox87ZWj41u
R+LuACrOZLhskA7bAdrRljWnBHOE/CKwAj9X1WILGXQU3pBsVLOxvAFZXF3g52CU
YmGLwVrJtE8s5lXv42b7i7TkYkrYtmXCHrXsx3Px0v+TzQO7Ztqiq5ahusYR+id0
DpmlqROsfipOIoICe6nbnpQ33zwz2IRxG+cCXdWumf8ZfUItP+vGYItRQjYSpPQn
x7rIPvtdTO/W2CzytIy67cCB7sET9AexETmjbOIegdIFkhFJNln6I6ljSl0E2c/E
MW4g0OS/54ZNyxdJWUAjR0Ciq/1QIxEYRnQoDPC3XZvwkqgDQ8BvbLpXD5nMEmpH
MxjAOaOuamSyMAn4poCdJ29RzGz1IrHC+2kwliMN3X2z+1XpOBspDBZ4dY74V4hF
t6IQVUljSsNBrbX/PRwSqmcnMJ9s6Qmebn/5mieu2gWdY4T7dKgTIUUkmYmcAJkX
eZpZwBTkkLNafqiGXK8Xd1H5Eq1cnb8xIf1tfzgJwfSuYOFR1jYaTOtOUecRBY8M
JSYje3UXuoDAsfiFW81jj8Yy4csARvQYMEM8N8PmJv2S4QqzDZt+L/dS+Nuo3Rrt
StdNpDGpOKQhelE121AcpzPAGKAJ1n5ZfprnxU9O6EHqro9hVrcqD353CojvjuhE
ROVkYGK9AerGD1uNubKjMeAwFnb0K+rJVLzWZ2dK9ACd4WxiGC07y5xOXD9T2uYm
WH1W5PBdV0wzEQ1gxXquYq902QKkOFHzOFTEmqI5cfBNldZCdDNsL2Fj/UmWZ2F/
S+H+byDmnGNhPklquypBQQVXgrK6VE9jyMDvUb4+dmsK98F2ABXG/brbTV26IT1F
BrmnwQ/VQDMeKG8yABhVNVt6mVF2nWeS/YnMMjKCFhTYs8iqZH5B2yIMrfQebp3e
sdV1CgJo3uXoGzZ8HsHW8OFL22ntVb1h3f+jwid/SpO6gt2QfsA4JhUE1zdn1wg0
nJt7a3BQ+phzsH8PasVitRZW9XjPpbdZ7N5x8j4vYmILCysI3WYM3YuX+9gjvmbJ
QaEQ/+syugLFQph38rpYb0CFqtMfCUs2nTzT+kGlMyZw9/1VDlSa7kSdSLAHE3wv
H8dirMDk8c2yZksAUZ4H2hlgX4gviowgkQZg2Xy9zFRif5xfMvGqF9EqU4y4iaVR
Ug8NgHyeAsnQZs0LNjPfhLjjNuCH5TMW3EtQSCryja5RJRhf0D41DlBGMEaxrXSE
VfOKz3VchrkMQLK7a6V0H02Gz7Ii2sg3fvhzyycWeWsWrmd7VfK7gtQJlylT5lev
HrIuBPixzRR1XVniPDk313OBHcqvlio7b0zR9P7XFJ+h9op963yaiRzNMOjSygCW
1lJmiGFnYCpq2rQf1LsQcl/953UmWOftxgxNkc5CxxmxHjrKsdn8acjeIlmOX1Kx
zoIWchaY/5XondHJek3IqAvyxt4wUp3N6ecnCBRq/6WLIkishdGqr1T1Muvrdig2
GIiggt6mcLr1UizwaDbxs8vxGXGD2ImctI4CJuquq9L/vC3eKH4cn48mxfzHprdh
QK6NLJ1VV3o5GG93FVZsZofc8xC8Obqss4ocHkfZyNd/wCUe0mg8hg07wRh6kT0+
a5MpIoTLK43RC+B5cGoPAJ8Cd5nsjKoT8dMnPqV/uflgiXZj4o+DLystuFJAckO+
t+IKcKSF6kZq+0YBtEFBYk1sYPp9Hk7cuCs+iRjPAcqiM8+a9bMQotsgK0oWmTUy
Me1zd2vsaGGjuQFuEiuoM0dJbUEGyfKWZz7CfYwKdlBMyVS0zGfVpREKuOtQpB8w
ziMd3pEYBzTtXDKVlAiWnyLCmnQujHigPail3yXu2pw2vNMrJ8rBWL8m/dyqg6UK
lIwiiIOFzDEmG8+SHACIvv3/NEtUkE9H/WI6v8ILdXSlkMm7fjjEqbMf/HvkIDdS
liTQ6HItKuPaMF6+vzISVZ32n0nJJ44nEio1Ew24XtdcTVKItbzBYOS+5gNaUS4l
EPfEZdN5SagCu06iPjvDv8afFFL+2XR7jdYC46XtzfJYKK/VVS6Q9OPFvPHt2NGI
Jwcyo+aks9rXfl8Op1IBWVS/2+ARVTrkrUjoA+CIeba44nEdoz2XjOqqXSmf9vkh
U7NgAV4un0+vL7KDvk/nfL4dzel3OI053PxUODCLJUHckQh2AuKKXg9ghcmPJ1d+
sp4OoLU9BLh9kiBn4/2ha2NBkKz44/5mOLBoEXqkEjG31ugD8phdrsaJruaigMxz
FjrCxz16z1nQKxAenJf07P6FE6n47eDCqNDNtkpHudMYSJEdz+itirkcCfLdiDe+
G+cWpAnAMjVkKwMPer/84U/4a9ThpsJZWGqOSEdIapdKeJ/jKEXiMTEaZMtfffGm
FAAcr1yVd01LB2ZV43WIOE7yYMwV7kqKHL6ktSL7QD3/T4Y/5BNphTjxZ9nujD2d
mTDCgyVvwlZ4Hek6IO0f8fzWMhB1eHVfJXFvN2WjMe3EpTSMfr47UQoNuPko4gc7
X6EiGRZkL84vBFE4qsfldDLBdwsdXGRcAFUds55j6bfPSPHLqQnzTe4zLU+yjqgd
7eX441uPnY4Xu1D6KXpvw/STUhR0vFDneDq2hqbUrURWqy2KUGbS6ws6IjyXw9lE
49f6NuzYs6Pqjn+1GUIIgob9SQixuycLs+8lEMqjziPIW8R3gQ+shV8Nm7avn1Bg
b/osH85C7ZuqJLEdNNpjYY9b5/uvkqdQ1lXbNPWmiw0cD492Js7lDvavCmJib8Ga
e3NSvZQpw4emFHU+1YxyBYdLtVFmBPxHban8mcFQ+aK1rn/yRSfpEAOBERcEbwbs
vPh8YKrHHiRFkdGIWcnbKXqW5JG7oVRtnRYgez7VBudqlGS/YmiheBbxoBjGfR9v
0BxdmFRQkpTotCJu/pyW7CP0qtlryNUO5jLC1KkOf/CFr8/Ur6PkWhsu6bnhfoeO
hJwAdYBWDfcOIlfVZzLuVp06QRONxESOxMCAfI6W0W4iXxHwDKl1a1fq4LY7OhgX
YBqRl87cNKLUKDhhGtLSmRiWYDZBtoXNR8Z2Es3mwxHo6IH1zSx4fQhoW9AHlvDC
7U59ql7IgYIJMbjYoRbxeHEF1i8uMZmgusnV3jIyBPmJqH7GzTTQSd+gV9mOHm0t
G46iglNHkUmy+RvLTqiUHnCoG5VTrz38InKVsU38Ep6j9pPBJnTCx3LZQq5OSFyG
YFJcn177OYDnQ9il5K5rvPjXy+hMoenPqo9agCWuKNnRtQ1FB8m8wa9XKaJgFjsC
+dJsPVgKmSwVQ/9adlVWlYbZKz2uw98sIpC5QFnv0C5f2C/YKjjcLxcxLnKpmvA1
y7p4s+MBFh3SwWEsi2X2XLYldkrDxqtjZxKfAqCKDwUVbeb/c10cCM+is8tmonc0
xdWW9r3wE911XX/dcGEaMcqjMQ0fAxrsM4pa10VmNcaiwafxr8NPHl0UkAlf50xz
6S0dVNh7J88oQ67C9q/O12ITXzTvZhQNutx2ziePsklgA5RWc+6XUbT8VTuZImPs
QhUp/T9NnfhKt7eMnBedp2Auw6VRUJLK0AUIh2B6MyQ4RmrNA1ExkqTkODsEkeq4
5nx+HL7HZJAoasvLwhbEeYDN+63/m4+2oTTxwRadjkaeHa5LKCiSldlONoAEtUyj
2fot0JK27OUM8YVePePbHvV+vHY3Yw3qc6wecSdqMj2xWIZsj+mvVGBj5qGJw9uX
Ag52IS1S3gXb8LJWj3m75p+c+6CAVqBAEGaluplAXIfHBvFlPMi+rOCPocf1vhZJ
oSMaIi3kICdf/v1ObqcuIc11h4CZRmyPzElreVOEO9OE37v9gEPdv6G5SwjtbDu+
k4ipxSPUvET1iUzfaisC/LwFgM5NO60CWxFVkaYYo7D+gjMWS76SD0Pw7XJGAIFO
Ds1M01UG61omQWyLnNGVRFZujaRnHpqeVa6zIyZTU4Bat9OKh7qbAFlmprjk0FFt
zE0uPMDr6Gqbu5/XV5n21bKE0onhe2FdQpIUCsnY9E+5tLqphP2H9EKStAE2JEze
dsgmAWX4bhh74Fl71cuhH/2yT4Dp5KUMlXAzN7mV7PnTFV1K/SGmY6f+lVd6Gfw/
A71pFscodMBR+38QGVPywNmTJZ3YBcK82Iw9uuzi5VCwd0Q2Fk6HwqnY5TWrqI7N
iXMRfV7LvV95p8958Kb98Y0xBN9UHOm7e0G7Y7pHRpTipUaopeETcQQ6NuSQxONC
TGYPMeleGZ+37HmuaHQrG+vCCFphDqT6Sn/vxg/q4ploDyjF5QtEv9NfzGbNbB/e
ZJjFqBqN6n+rAuzRSY6V4pB5EsZOS1vOwtn8y2mAyfwJFkmEnHmJfYjTjTSXzufv
uMrR78oB0Yr5Fjo/Vf14/wE9A+viFW46/6StT1s2IdsceW4wXbzJ04Ws/221w3Lp
OW1ILpCtk75njj75pz9IMr0HTJWAKKy8nrbwyubCoa66q1WeCcpzOj2SYIJ0jgwI
QcpFr0oMsU+D46cij8TiylfMte3GbR6IYdzZ30Bj7Y9oBxUpINKb10FwVesil7DP
f8/s6joXdiW4pEy7ikaVjl+JoHIF8u0OtXSzfYf5i1slR5kQWPTpV8xBPkZDM9wV
9ptJUUlUAREgQIR9UF+bHsNfOh+WiiZMoDP97TygTZwpzj6f9KY6zRLQL5w5Y3QQ
yobFMDT+mtVzf9tdqtcf1d73Jlr9Y0p00I2F4Alo34AqxWHe+/OD1w0ys/W+zapb
lXso/SX1JpmgmvouCsoBiFUxKi1Xh+8Re0yoI2w6t7qFWu4DRAazVLLKT1ExKl5q
o2LC8DwOqds2hdJt0PZ4EI9R5CTU/xWoMMXprnHE9tbA+kU3QwPie3msyYfyG7WM
FtKbdIsdjt++VhZdDzjWznURqEhsy+X5PK1CSMWWPCkJzJJtJGO9EtVh/xRJ2WBm
2Fuzsx+9JxWbQ6ARWH/PzwhtGcRKRni2G/Ogc9kRQgJ6jSpVIiWhm69auLXt1FIe
Gf/TNy+L1I7rTiNkWtS2Os1ZGgayqtd1DAqhwqCWHDmsgpkFuVz9GXldgk8dKjYp
o5r8yed5AaI2nlxq6/9VGYrCEMSvIMVM6au+gK8KsBMh8EPSMeVhRS5Eq+kb6aEv
RajQfdH0iinXEzppKxqEKlH7kjVPrgX3d+3oR79LmEa5774m5WhZWsZrbeoJPrg7
5GzZLlxQKcEjz9s2dz6O5pqHU0wDtvzzHibQSk/1gXJX0VWEXbU+5ZTq0JKQqcHf
hqk2+ZxXNoSWilEhE0Ofme+2DDt9pxVbpE0Dxd/CKEO7f762AYUpaFYoIohPVxvi
tM0i/IGef5bLlHwk4/P5u0xIr9UKSbp5y9K/tOcySykEQQWXU0Xqxw8rbUm0eUy7
Yr2BkPIz8cu7EUv7+jcQW0Tkfb172+KWl/rYscfS91uZ6spOcR8QPpSUtaCH3t9d
OJ/s9ThezP7ah0EDC9+zvZGv877+Cg4MhzZ9iVtA3zsOQYtmnHeJMorPSUj8+BRc
wR75/IDSe51g0fYPMXOcEpDJLzP2c7bBea0y4KZzZuRO4tga/iP0DCzXq4Jg5RIH
Z46xWNvFTE1mJeIe0TROlXvbY/KMSI1KkeF6k0HuTKDJgcU9R0490XhEgP8DoU1+
tkCingnb2xe4286iMPw2mYR9IvUyB3fy388lD9d7YtGfpLi4NjPGg9o4Sl8w85gZ
yLpyCQ3lOYjbtwTqIatdqwawlUNgrizWkxsRJDi9j7B1iplie/4+s3CdVCiY64+i
yKJZch2vT47yrVgLDnJDBbH347gQKi6vbOz5X6gbu6/W1ya7cAe5xGMlOiCiuIYp
ojn/D6a1wR8EmDluLrVvV4UM7t1ebT7NRO6rotPLcIrbh1GfJmTphOY/rPKdXkZ2
cGdlDkyvoze24nvtUlVdc4vAkD6rKosUDARuBLXrg2iQr3HVWcyPOyXmz4FcUVfi
Ha3o/KyX89rh2FJMJN/3d9HQPJtzFL6GdA0RHV0CvrHtTclSwSuEw0hlqTp/V16R
gfVjbcCzR4YQ+wiGtY3Qd4Bk2o/qOKV5TOpNv2m3z591o2glJzqX/UC5KF2M5FAj
0xvDe+WcB3soRjx4xYa5OE7R4J8OiQd7eniI0Uvc3c/Lgg8CVuSfBi1nMr4a6hM/
tQ5cEVW36VeUKA8dfnH2BVmDd9R0/QIw1EthLQsn39ppY6wfpxCFVE7vWte0eflt
7ylxa6dXcJpiuJkyoHQiVBb6DPVLwyO6s00JL2RLLFux3QyigQ6IM6Ww9TVCPODT
tQ2Y0Lh1D9rrbqW6swjABAWwSvboU11O6tRafSepuAfEnYxgfcT660CeVTlN0Z9p
2FbgFCNGDD0Q6rdGKZHirfpZ18ePnWVF6jPe4+5a51cZfhPepK7A/yu5DV/4u7uV
3C4exGkevqzHDBIvCMEEV8U6pMTmYXhwGhz7bTE5ysK9KZvKsUWisvdekNsSrtMJ
dgxqQoNfmAutJJB40DCMdFOYBCp4GMqr3oJO7GwVSX8yI3yNK3ady2Fdm/K/hr7D
fa1TdbmhGcvmTIVPeSUAw9+mBdsZuBlOn6if46JBcmCdB+SCjzVeL8JnOwHNSSll
9QmMSPBUGpo2czzzSX1JGFHetue+keoKRMRbjoF7aXdJJUsK1JS/Jxx41CLmsUkR
dk7N4XYvQ+jlAwkHLfkAZMnB1StQ733FkAOWVnzQagm95ufoKwmivzTNcaNQaNRw
SgEvXspnjQNu/CJ93jlDhVyJVSKAY4TZXzI8ZOXYwviC/2dK+LMQ8nG/E8BB52eJ
ua76SJgb1HgvIf5RctArTm/u/Jp+bEh/CywUdsBi/3j1SppowRd//HHq/XVXqUEM
AwdPciEdz2Ywn2sYN5TffIlT2A9ojW23/4LRiFv7qHl2GudkvUhMtgsu9f4Jl1gw
xiz3JlLowfvfjoIfZioHEnmq13FeFwTHs/QE7EE15dAVd0/pJ8qIMriFKbAzK4xH
CVliAWMjSihpTyI1NNjYqmx7w0p4cC2v2GSxv/vdDop9eSCdDkLENyKxsVY1dS0p
oVNQfrBBR7IirGx9ogE4BYXhxHh7tEFxSLlzvF2wEu9plkyj2dX8EDakCOige6Rv
X4+AL3nFP4wwe1pwqW+aoyQmi3tEiPsxcGFQA/h+tNpDtHMAeFjcoqaPPiWRXYJk
pPij14KF/nj1EeKBkN7XGSNvbK4g7kfZjzbb+eITtz58GGeHTNzZ8TneKDtHVTs4
42Bvd0X50fWv1RJlCman9lDSRT+AtBV0WpiaI5K18VlCwOn/hNxVTbuoQXPsol6u
E1KN48uRvferdsame+uQZMS2Ud8GONqtkV8UEowbvhJlyDwJ17X90s7yoFB+j7kS
8HQ9m44E95TEakKfRjyUaQKnZufqTIL3Mwl2SrFyXkPbetd/RQpUfvAXMu2hLfqr
Z38PaUGpYhCpET0qfFObnwK//6j8ygS8HooTGUDkqJ4IBLDTiXdCSrfLcfCx2s3g
/CzfIT96ZqT1ZFCzAhY3Ja8TLmPDAqeVZCuaoZvpSIHkb59SZU1wmTyTlThn89bk
ci73qQYe/UAMp73C8LnVrzk8/qNtRkYiseonluQ7YB7bMFE2zCgks1O1YXvkiq67
baZLuqjVTyU7HDdq6P2bDljN8LkPz7ecMjH02cgam7vF0f8KclJCY+7pSigkhfuC
y4qK+eDSAgLA258gXCHs8/mLuOXXE4h6j3NWPFbrtoxeSSd64fi4rr3/zxfsk+RY
UjrAJ24CBSvuoeSZ03mWabHQRICQH2kvtxB+4wmnuZdX8MvIwZcUzAHFUhnwqAMg
+Q6T9ziIXsPOGPPbn7KiM+8tQSGFwI/YKKz4AtZ4ccP3pf0hnvf2FK7ZDkZWWsJU
V+WwLoqGSgapVraIHq9G6AnBNhrIflfZdpbwochu7WjyjPKydl0ub00UkPHB5DL2
vfsJYEHP+OZnxnFfFJXzcCLaQBi2Ys24UCZ0w6iM+g5FRU/LrbNPizqsXNwXsYiZ
BDpguKhkAT36abfWwkVFJWKRrCwzbP3aOXNB8ek3R40knhuyXvVQ/fAZavBFJn6j
r2/AztQDmC1v3cEIdausQh6t2spaPv1X2xCaWhtg+H4kdXjgHn42GDmtLE0yXTyM
2jt7Ag1e44XjfMbz6ZKiMlf6kCOStFRrhupVQSpS6cRdTeZAPUMc3GkdQGCGx38r
cuS/rabkcN6stGN4jEr+sdjvl8yaOu/2oIORwhp+uyrKF/bvONu5IQbw4fInDe4F
ZDC2WXjO0fKHCd6z97UOX0IrhSU+Qd6nIjama32Sdb7hLkVk6/IRdR3pI6NppLTL
siLjjzMvINX55/C4voQ3X4d98BxYkch4LkLfXdORwt61US7O6qpu2EvwUaGsi/xQ
CkR/d74l5RMeRBsaQIsyGeMguWIT1Qv2x0KKm8t6qDEXeuu5+2diprn4b1zISWL3
Zx5gCtESkq0OSTbn2lQCLmimNnm7wbCGF5wN2Ud5wxdkQpQDMRCUV83EpftTKfBc
XsK3VS2Z50xqo1WZW9JJYQQ2Elhs986icn15uIq8TfsAzC6CjmIo2dtaxyPfcrxB
Pt74aVHjTURvf+KWNHh5jUHEwPplrBBItDIFTcUXp5I/E5V3oPq7yHRNS8u2Qd4l
pEE9qPokC1B8HtlR8qpvwiiPzSWSBDH6+r2y1BcEBvSPFUGBanyzqS78P3sgn9pV
XIPdwXAoj42J4regKPk5TXIp462J+kB9PEllEFH3cJjy+K4wQCyagVfYLP+iYnAV
ba7LFpX1JEqMpXgB3FCJB6H53TGTOlXZKrk6zTjedZyZ0UltupCzqqJf38q5DCwO
KBa9LMlaUw5dH1jFDaauwE1ihnIgTSjFPl246DqvgYkfJRxFRYPODyTOe+ruXHND
xgkpObTuJKhIhWrTg0c9J4C6WmRihQVVjPzw7gBjbfC/ibpuYKHOH+8HoR2ablY7
cVZuBHzqqJK+ywfzyAqbC4FVETUAN0Ad7E+P6pWh8SpX8YFd6ciOzAcwTXd6Ts2R
RMv6M32o6QrT8KhM/fV0ZI9rk22MzlInLipR6kg9B0wbaF+j8Lyoovoc9q0ZN77q
ws9Q5eml6IL8+1YbMk0CAFlvm/nw790dBMSpTR4ELQmL1QODfnMjbLWwPL0LYbb8
Nlpd8vq2SuBAOemVYBX642ZivpfxD2NgW6yuE0wZtoR7oEQwFQ7DQny4riQXO5di
3g+2Il/bUiJJm1+YtBZMc6yrP43+wccuK/NbtfPnP7qdSzU4SB3wR2jV5wynQaoT
An0mDBOdBMm4Fcl+yL0KMikpbJuF+/1ENUnfhFm0PBtXtLH+PgLzHroGqSV1ChNr
Wxqx89PW72j/kob65rg0TNvbIFvdsT43uEliniVR/C/2oC82GKrwKp/4nZPqczD3
3+pZsB7rNlYfnCipoTflb6hXa/HHRo10DUhBS5hB5+BQPKT4wzecMZ7P5EyfMDhv
CkQzIpxNh9k20a3l0HsbgizRzlITlSPBnJEs29E9KssHd2MadFaI7l/P7v9dYV7E
ZxV5pN2lJ2k1tF8W1752KzaL5EFQ7AB/hfa7jwEA9CRka+AFS4G3QCxWnxYKIG6A
FbyrlM32jnv1W6dDubsmsfTw5KzYqCJDlk29yheweAadKMQfhz7KqT7gDoQeS3fZ
3A7zi3VaT0OCNzz34h547yZrj7u75jRHe4zsnLdiwiLf9pKTspBgdYuDb1wnp3uu
FKiKr5j2ryNi1WhSItBiayvDwNUhwhJJOs9ZpqQY1x9885Kuun6om015wKPm1S4O
5SvJNkeKj1J1dVr2yKCOXCiFQ24QRB2bo1A6WWsBLonTTR72CIslHRxgHeJx0Q1G
I+SbyYLJbOb70cezbwtmmr++w7TxMNlpNnWzHms5R8fDU7RoHyiRC6QfisiChJ3T
EZKCKSA/7FfOEfwKQ+NmobHAxUhxFIgxfHq2WmYYTn1BiL11uosaNlB0c4zGaNFW
U7PSwlW6rQr3ogja9W0hm9emi/ez24aPiqFxLmAuthlFsz17MBBpq7uPMoKHtrw+
TTGTvFZs4pHYU2tCOMye8CjVi/Y7ULNqNy4xcxqFJwXfmrNuLhnMsJfDGsHJ0hOo
LtYtFqXCkXfiPXwqg3kJsL3bOIVRDodh3D6jFUNNzGTqr+SRA0EFbpvEve586Ud7
Dr/76v71dhQjB/MOCVh9+OHsNuPsv57jAPd9e844E2DOBLLVfyZTZ42TxIUjfg6E
NpHadMn3lE/oDuwfPQQ2cup7cqI5q88QFslFBb9nREwYY7JLTLcn+ZodBabGo7iX
oRK7qOWPzhDuDK41QiofRUzl8cnuk0ehlIVaPVHYvGKJlbFe+FyvHXyc/7ZFuYrx
oQcKdxTuKYp0xs+nzfce/+74eVi9RpfBY2O3pdWhQa+uDgF5HRflLCtcg8qrhJKU
FYtVNFGW/na1pL0Vje1ZF05hJH+s5U71W991U1ntISrNgwzmtSTjwU4RFP/qwPBQ
EQUdc0fzHBLOIjbikmkDIwxwCl0wtUvj2KOiwmII0muLI5k8faGclT0n0nqwT+Af
lLk+JccVOpCdHrEHJtby3UQ2/C6/WOduaH8sJVB7YmshCh1T6JEty9G927DM6Rmq
9rurK3HCUz/qkPZJPiNPwFXjNnmW7fEa8ivhi6rqZA3X9R6oTrThMT2rXtF6RS1F
xWcdDLFvTgDuiMFoSfc5eJFqnky37BSKdYZ71sKclTHbRyL44BXtQ2BAF+fzpdq9
zckRa08HsctaMCH6Z6oC5TBhYuYI5QJv/WYjuY4S6DueWoV7+XanTWikiwQgSw21
0qyRu0QD8mxahTG7hE0KAqeAaP8e9/RFK2o2WX4O+oVY3VjXnpwriPrkTsFtlBpn
Xm7OwwXOZNwpqRHHzI6CRkYuUyv40tNvY5G8viMezjBe0Zem7K+msko3Cwi4GdzQ
qcfYfjAxiD3vlcW1sah14xtj3zWxeT4les4gq8BySlcIbgV8mPxGmcvkn5y/tWeB
DeUjNWbGkRiQAhC/69VxrkM4s68lFJE/Dgy4Byq6GteMfLIU0atVEAFKt254+l2P
vA67UZGVaHkwmD3rrSwAPLtNcrG0IWfkV0h7K9XdIng0lfF7Kw4Uy+xzo0zlTh5r
NJ0cQYCiOmMAr555nbvwKwcyGWjwPJMjTeB/PlFRy/PBeb09htgFovAXI5pZrsY8
R+TnCNKottKdS6GrOdRXxik8oSh0MAKDRGY0nC1iLYB8TOWy+xX842SzQjwHpFAf
DbD8qmeEWEQMBpnARSQ5mRH+rrn4Rm7q11L7h1dhptIC9HZtzGjedvF/mNfVucWu
ddsjeNx1vuAUWQdpvmC0u2yw/i4X+hWtk3XeVYtkVSlNDFBnwGM+Ega7RhNzsWxm
wc2hHc4QcTJ1ppu+H4lO4OOcKIY6gL3JNLGJmkdViSTmf71emN0c+LXL97zWIAdt
p1SuLGo6UMzhtnG1+oL92dfYRIUmQaCnvHzwIuW5mK8XkopxXP2irXg2gGNVotZs
dN8F/F6mSH+6OBJgiak69zSFldZrLydnN+kxwiIq8iptePmWfzIrYXc1ruHNOC1z
CbBEsT6DBFbSQSMevJH7FNzVoBwpDjTE8+aSpFLM/6bCEGC1vfy5LajcbkNZbuRP
Hb4VgeaL/nnPCp5jB0RcENnSvchfC83rNq8N9jGrhpO8QWlbibyS71yTrjJDU/b3
5vI2pFXcpTxVcaHHI7rpYLLdby6vU//wyOexw1l9O0ZZ5N/2+sZWafrYtDcD049P
ubXS1RQh6tMmmEXuVWnj7jgG8ROfE3ghtfXxPPf30jpkfHtL1eWKPcXu3YMR9IkF
Sdw766bxwm6fg+GUMYFqG1HZnlV92SF/wJh2iMt1411X6kerTGWJxABE/4vaYuhj
do60RDPgy9AHzWFr9U5HCk5Mou5yD6pA+wcysAYuI1NH/gTN6mKOmWDRi7OtYcgf
iU+O0TrC6BMPChMl3qhgyeDUxYQycTkyNGFHis5q5Z87GvsDZRUIj5Ezu1Tt4w4Z
+G66avU72SptAmCv/3OF8Kb2c5inbKZbH2YfDjszItmbDgUBkpM+nVvBB1na8Mj9
qDJY+qoBat1NXk1O6L7iZdkI9YRdbg2vNuU87HUwkAAAzvk550qN8wmh7TAXuu8l
xJiMUPH49etlHv5lpg5F3pLVdO6QKoyMJA0a3V8uuIgQXXFuwVJQBsLiklJx0jP+
aqZojX7HQXHp0AaZ8IssfXtgY2x6r0R4wWnaIF7JKx1SKcK7DDAIe2ESid+Ub+yi
w/8TJDuuk95XJ/9ANa6nTf4pHcPfvCI3X9ersY3ODfHObA8ol5oS+NMBqFllV1Cp
5uHDsPTF25v+kgDlzFgO74qJj8J1ukqXtlpI2kXdThEv2Vo9DzppQcdKMyC+Q8JJ
dcvw9imvZMdcpwGWnfXF76jpCvTGVkjekhIgcxp761M9mzy2f76sYk48Xn1GcC/E
LXO3BNm89PfwKuUGSvxv2HsuNbzNgoAqwXwu4s9XEDVNnJM/dxVaIOhBvUKi/e6p
0YaYNGRnQCovTto3EJr+KMBKecsB4r/ScFuEn7DksWQ+XY9HQrlLZoniQZwh1cpR
FZ74hhh2TRIs2edgwrb93ShnoFaU5D7T2owtFQOyAYJwRn004GcxcuB40D8N1sSq
yAj13bo3YTBUahcEDKeaZjXNh5t6yJswOmUQZLV5F6TGi+JZVS2Vw96+dv4Eohux
H84/XDhvTGzyV/ane1s3gHodDPs5b6avRa09YlXCylKEi1rZLiWBPWzeBhdnBvng
E8xZPktQ5gZeRjvvq/BXF3ywhVr5YYu8PVjLjBkcKrseo5TJgvShdNvECXfyGpaj
u5o5yTPVNm9npXXEvGU2Qya3Iyxfq4pQzMdBa+T4GFqAz+hNo8Ov+9fmvtVO7Av4
UTLbZPjaJi/H6hfOaqsRJaHHzD7i8tJd3bVEORFkUuBb+lfGUlbofp6wk7ok/a7l
7VUvSpLQPvNde8c5mHKJ3K0ui2JT/ESuige6P5AyI3R+jH5G3Hud21/x/PEbO0hj
wTaKEzKP814+B9EMtusFMwVCyXdJ/aBXvqsFQ+npKznL+/TBYgQ9r2V5ZaE+M/Ws
b87nzMwvZMY3PeQjd0623vW22LCvGagtCU3ZQyFJhSeGf87KmG77Gp1iUUkM/V7W
FJXC2ylSDYfhJLHEhxDvyFv9U3zdd5iwUOYszG86cpasEdE5vUxhu7VYBVRZR5VC
rtF7LYdpeB7yTH+OteOAw3xe9u5yIr6HIYavbqhTbrhLWD0UhdUGTA83HPcP2igy
vd7hpFWcBdaZqneYDYI9zkXDwTeUzpnWKdWjMEg/8Kqgg0f8Qk7/CUGGRFt+1GTG
aLiT4Kb2gseZ0pKGiKQvUlirVX7HA62wDvs+/MuHNm6NoDElKOXo6wP8nTysaiDt
KtGPo5mT/eb80KSL9PVMD1z0q0QhKIi/mnopod3sWWJKB1Ue3Tt9UX5iOM+LCB4Z
qcp+qwsd6g+cVp1Wa5cN13HcLNN3mJJf9OnJKRTLlIpG7J1i/lLrIbMJjSWRpen3
irtkf8SpXOi5qmRQ4iQ615sHARg4zhBMrmjDqF83+xojGTdf3jPmixn84MNOrpOK
LupUELjVWnEz93hdcOW8SCci4wsxDYAv/G5pVLJywK6VE89NH19Q6kTtifjCsjq8
2GXcW/tLgY6fU5UDDIugIvqowFysWyEcy9sMtzsDBQEz1dwdkIHirIAvfrzbR1TA
UcYk/8kBZoYB/WxX3nMfrtFzMbylratwrXumtREutTSLcG0CGUyboWNcUikWbi9W
DC7H1m7V2gB/OVE4F78Q5/xQuP/mPNYFsAMQE9FCd4XvLMVbYClI6iY+jKKpbJQf
hKNyavl29/pbPtoHsIVdK1RgDGQ6HT4T1WVj1ZO5VFMkAAom34kK36c234VAuOzl
jhF8aRzSRqz3J0hDzhkiJ2I13MAyGuFTCWPCUCUk3OV6TvXF5wlZq9Rw3FMdgAMd
59haD15RAmgHLFQn42TlZmmOrR0ERPJ92c62osxAj0/S9c45V3XgbfOy/hrGH2tj
ZhZpFLZCYjp3WiDZSx0cEZMtkX2t55A9fhmlq5SdKh50iWBzuLAEeZ3Lq7JtAe2+
G50JClWygQ0oeZbZ0kRMp6LnANYDvmc80wwj56XNaldVA7n27Yp/7pXOGX1CaqsR
ORP7xZaGWKKUvp69c8XRYnjI9W9TRkyi6WViW5Zbp9TIeUuEirj0Y7Tpzj0+t8xU
/aoBkTznd+vXfLnDGPBmxgs4v146wOOqRSAcUjl5RH/ObAUmc2sRNYpKMhzC4BM1
moqIt7u1P36cHCSy/zv/BSczVrFY9wD4lEoudjeoPG0+sOD6pzLA2kE0x9Erfj8G
Lb8kjq4Ooj0CfcX2DofPJLBIGhQKQKCK4CXyPFGlMkYY+5dZ5UGWveep78nA7FUd
McQYrImXd89GNGDIEO0Spr/jqlu/Fn0m+NCMLlu2xNLwsjV0yF+6nh8QArgRr2O6
Nlx1zyE+TVQb8x+fyjW84r+HsBx3w6JYBO4UDEeEjX1/0L0MBOGVrJg+jxwG3jxh
C6CufiFZOtGi15TgQjPFNVABd5e3uEDcBhtXYc6DHHjNbpkvuUXC++y8SZx8opAV
uN9fjdTQLtnuFvdOQTNIHDQE+e2PRSujdlAz9/phb1E7Qy4xiB2fdhqq43b4rwF1
h2RKlU4M0wjy4ObTAWr4DM151LQgzoeKP+WDjUq/FyIC4urscp2bClnNxF6dEZ+l
cVSwnACY/FcFLgNQ+yk/AllX8q1C0dtnxGxoK5SabGPSq1D2MVuiF/BlpbQQZCDM
DhggzB8zvcd2s0eXZTnW5pYzsLqegE08Tqg+49Mpt01TTZTY4ymyBNDuJrCT4c53
m/RPpy2o/+9+uN3L7wDSiFZHKGF3oQWGD5VNVs+M5YCjQok2LveUqkDtHWSH2FVJ
VhZZnl3Nbde5NNVt7JA37ggXfEWOiQz3gsankcHvAqDaf9L7FDcFj2SGzs4KHRFF
MtdSx5gYXCDhlApzPeqy3iwVrahq5U4eWto4AX6ZA7Jaoo5emaqE7G4lDtCmKv6L
sZB+w57HGbmjPn3IzsxpQOab2swJtiu9FDRuemhN/Q1Ao5ueXHISSLXDHjf+WzcT
YnvYf4hhqSrILrlIX2OyxGdR2bGXY/QrAuYiX/ie4JDN7CW6UBykRT4GKFpGthNy
7ds6o6lx5VR/076dUgtwO3CzQeaAq509wo4e8NW98BuinGbNEpVrFdD5/0xaArgl
B3xtpWNwPigRL68quORm14O/ag5I8H8hlGsnP4A7F02PvTjJXkzwoVtIReiC1hww
RO8+0l4UFsO+5KeKKFwaMIMzakzLeRlXe+Yu63Q539wbho3/kACb0YhLd0Z0tYKJ
r2fopoEtip7073eqxXJld5n+6F41jiuhMiK2jaAPcFNFLcbsRLeJKxgg2jeqzZUB
iEWGfzTnKVRRolfCvEWlx+YJZtv/8FqeBxdAj2Cd89KnpWPR2nVhneCqWK9aB8W8
MK75dJP9jKYc7Wki4BuBPIp72OyMW2lmaq67K3v3h5gue9HNR7zZA9lKV3yA+eGc
EQck7mqsBJWpwUklyZG+wtqwxQFdy5DsLPmTmbGag0DQXnDXg5AVfvz4r93kAXvG
g3D8lMWkxgKZ6cdDBlOl4iQHLANtbUJ3WYXlXVs2pN6zGRXIlPH/T7Hxhm2MJmLE
g4I8lGriUL0k+1a6kH2/pjycG+2l8liXHxUDugOZOg1d3+PFoHE879Bneaiht0De
RUeSOKBgvmJ0BudRZ36Wke3LUcGIrS7xYhs2f7CEcg4R/akJBKXQm6f858UQBnEq
W018Yxzhxh28Dw5+hEwxGHcrli4bGezG3EyVE4l1qPVdp79GKcUfWy1gvwePYQXe
lWKqPGE6Eh6RBFxBuuf3Fn6xBW3IW7nP0Mnbe/chtBrtJ6ga5t7fvoICTNRhLJzv
GKBR0WOaRNk35CFqJJFvdAyCcy8OqC7Ebxv/H/pu82DIKtL4lLvWK6bWtEB0iQS5
DSUEgAsnsRUPQRCz/fbQyV4+okueC9pyCeJWesPVqhkmOQXnA4crHHlrK8JtyCC6
nVtZ17SzeB3E5Dfl51ZVJWiMfnMUn4aCbeOPeIfdkPOZNrZ6hWfjBwH1XGZICcBB
YOrmquqh57lFEGqBDtlw+jP8BGXJagpeQyVOHXWaAgl7RaJEb6VIbtMs8xiPGkKx
/A+C3ylsv2HXGy6Q8w4iIYobO1S/Jik0HLovALdtasjTcvy7W/iGwfCGKMIuyzYf
iOnTuepsIknA4gqFhnSi0g6GizQye8SFtmSxTRYe6HQtSLV3FEEm6iFvt24Z3cw5
nkBqyu7gqQLpO+bTxFtUuYTZ+kOB8akcbFShTsyTcmvbASMcUFhAAF3eBBTbKdBq
Y92PnKO+9Bb/QCwJQvw38eQyw9Gjf2dXPtWO394wRvSduFgE8H+FLN6MtbkVOCdG
zKt16RIGDYPc86hRORFyGJSYYSnrzeWCtxiQwXsR+60a4stxTkVPhQpcgQ8z4CZN
cj09LxUJjkxujox463tslUMztKaalFhrWpqVV6hAKzcoQ7CvXBQyWEr1cjYjm5tm
KFRTWXDptpj9kQjonVDoVAeN1F1Bp39GiECQ+wBiK6ouZdDZRczNYxdIjd5EvNde
AYi5+2fIj946da9bdx6u+MNp3YNbZjXJmFB2W5axzbp6ThhoAFpgd3Zv+XJjLPDb
5UbWLScuCHXbLwq64QokwhsBTD5QMnorPkhxNKVOl/iirseNEmLonnL5/9T9MZ8+
2Kv0YuAvmSGtIhBURl2HqzI60uTB+5NQ/n0wvTJmSuevOtJLXV/R/FPeaMvk7ft4
WrhdY1z4gszfboLWz8B4h1lO6tZd2HXGJqXQ48t4jK1s9MqXz/fQtiM7V295Udwp
33SRyyxOoyI6MA30CBAtcM2b2Vra0XHspCELrpEwTGfhzK9sb8/v6+8qRFzVqiYx
/RPFb3jp/39PtT1nL11oTwKWYWhcRzMDI1IC0FuvFd7RzFQr590j7mXUCeNBXb1n
mvlWoBEn6Mb3kXJIZ93BZIknELa6CYWEy2RVetHyZLWqrAnbbI0WcqOoFwj56RjS
GdXS1Tw2WhxQ2f1kFN3n2hDqPCfIFdX82CSYoDz5Z2s8e1o7YZJ8FhKfIMZM+oiQ
FFtCnOd6px4iLxDs/bxGPNLUl9yI/JrzGtkKr3xF2qqQ2P1GdOkbtJTCeJtve+TM
LlPVf4/zMBlqm6rYNAzoMpZnPF/7lAZA3fJmZ6TDqewvo5WYecwP/HsnQUClDNu3
9qSQLGstbXDkeYmcwyOeWgBqFcBafouygDYrkzynPnnlQjU71H2Flc6UtUF6IjsC
Emlv3241djCgM7PBLlf1t735nWhMZp+ztC6R8VJzlNCkkcMFheC8bn6fEWTEiefY
V22s3uxNNaGz4aARQejT/H6jzTzkAnkrxT5/zTpCEXl2FdaSXFie2FmI4u2lEQAZ
eNhk/R84oYzczZgNeEFBQ2ZiwzyeRjLFrAPmxEO9h9tvjcDqLt7E8oVkPkiUJv5N
JAhMwjqqV/whjfUhdoQ0DW3+v7/D6WZCH2m3LmUnChIvudIRV9aqu5ByED5jIpQc
Y8mtvoxl3L+5m3yQKPJymKmW5tNhAJNkvqgtg0J2O7qVdwzrqonMgBb1ZUu0Q1RF
GNHI1VIKEcfpaotxaNJiA5tsARIRRPDhF8vaKPEnhQqgOjw6RDITdgtAgnVCCsbb
n0js68vhCAlJgOQZcS867PFdPKlvNcS8tKKDFTxVrOWcM/qDCm9lWFMjx0Ifwvvq
FDrBIw1Q2sRipBoNV9acAmGNle3CV/wv5IP5fAmFTEpTDp6AxjsiMJB36cpquaOW
g+4J+7tMEeR6hAFWBIQQIrmhp7WM/JpYfVUlkC4xV8fkNZ4PioLI9FWJM6Ic/i0f
GspT5HtFxRJwDr1Uq/oVa1rJrwM7HGhKWi4/KilZO4+zMcgJZm4c1wSrPmT+UqeY
od2iEE5YbMK9/dSXXJrtpb+WmwmEWgo3XLMVgPbTwvodsKpfYi1zFGk+iEjaroh9
2g8ISm9ytkFzUNbcmALoDr6qKNR9Bum6uotwdaVwjt2lz5syOL2VwwA/QrTkWR5e
jw4OUY9dnqpIAW9jjmX1h/Dxw8IyPXlsMBvpnZ+7GLdX4YUOA/vnz95XZ9EdvFlZ
hCWUpn/gHVW5fow18mS+5UG5BkB4baE32UGANUWdpCpvOMvkYCJQ2pZx3B6ER7hj
mkS35CcpQ2yseyDqB1LZe3GmSIBBPIUvE9nSHM+ZOgEa8xlpGojcjrdZu2XJ3tM2
PT1C8PlT+ab/XFxO8SXCIv3eCQDkvCq+7cVPiixtTaqHIkJJGsgdPCY4NzxhcCvi
yXxjFUFw5TbNsYJWasGRr8VCc2PmAZCJ3zMMk7+MtTBHo6LSLX9LqjN2ikPrQCMn
jdELwenknALJrNg+aXeZR7ZKrELGwRbtBJQWPNhZXfVh17OrD0fmGWR7DDO2/7h3
Ar66B4UrxBWAxWpo8aWlGyTocEEVryHwdTVQInptLQIgu4PWAsc7zqUYoj8annok
P5CtvywCWPjnYd7KemzVbCJVCHSF6ORD3EY5bWPx8ziS8MFM+dBCuZXDsB6+KOBN
DxC3rZXqngOlVN1IbJI4ryggtZz7EI70nfFWWpyESv0Aj0gS4XyavmhQ5WTsoLOA
VO/0JZtdk8dBaw0kAk/tx7q9HmVZW7ZHPQJu+qZBHNyebYAerWzPuBHN2Gkyn/7B
ebLXGLVX7R9j2NJAM7UjZIBIl0JbBMDACw/ho7hC9Le8Q7NdgejWDFpbEHkc7PBq
tgIP6KAx6g0YnZ2UuOBXNIGI089inb3XQD9dY8FO49uLDD/3i1iLuyjdNZNG75J8
HcrsmBAmB7Tkqk2z0BvQVXpBHAAujeYOM7SUQG9s4th4iaWquw5Cencvmu4v2Stj
s6Ig8x05rnNJk0Ko3sR1M7NUb1J3ipoUwhNOtk8YUeFrXrIgbd2JofoarmLZLMu+
GtYWU4gkd722bNM0zY4lzNIu90gpTOlfPQIYptzITA9LaGA1IDPbE8VIyTcbGGT/
sSLBQK2dRyYW2VLQvCOEPZKv1xvR3ctI48dd3Br5aeE+laCxMM7ObDNb2DxyhSWf
U41T9NbdDWxWS/H0syIvQuPOTkuuTgPwNqmZJubQLv8EWSKt82QNLrtW7cNjF4zZ
q8UUOAXC1s78NjPZAvpEt0iQQ7LcKDPHFlZnkAuHtRc3iH/HMWaw1zj+HNg48KkF
prdFS0QIxwSCg9jP6wmuhPCHighCYwa2guNkkkxj9Y+WRbKjqYHM0mEBgiJmHDVO
1n42D2XzujVPojtbxmUBmrZnOMbZSXthPtHxrzEJi85YEKnZ64w05ggPgKMxeRMO
TZGysKUAXf5ofu6Jrm/hGhryXT+4edICP5xM7sOfnlJzspyfI2kbUdvvOC1KGCPL
4ZCgEYOfKjEeuucJAiJpouuH2vR7jBbQRwuOZD33qkEhk97b0aswhKg7dcR08h2L
0TZqsbHRIyBOhDJgmfdgmTqvVrYrLz55/Jap6npxUB46L4G6hdx/7PhfVC2TQOEa
AuOdZoUO85ksYIeoB3rqLNkeN2jOpjLpiCm8WtEoW3XQQzEPfvdOJzyUhiFljrhc
7io4eMTOH0xKNU0Eue+1Y1fvuHTTdG9dd+7tspxEooo+uKov+7U/t7rODDTmnqW1
6KN6n++wf75AbMYZdGGwFaZgbcEeYD4xtsybyvBRROvVou/bO7CRpyp36nhNgFPn
a4iPEMvSGdIqYMvhkfyVey4Mgm+J+9PPh4uKwT6LosasOzDiJkCFj5ldYuwJ9RsQ
CU5rvkP2+xppyxr/4H7xDUetAjjY3L8KmSUKfyiHaqEY+6xi4P1+wvY0fGkw0daM
bm5zZ4gtnZbAqbyGmQBFRmKU2N51gtVx3NWVUpVpcOGkOjmK67Mnr13IPcgMXBMB
wu+S905aBC7gt68RuQIpDnLoS2BLHvEwjocy7DozVREi2NV732FSeSlIz+VcGOfV
StoSvWHtscO0pn7aj4U0GyRJkNWGBuQ6lHv+FIAKnckAzmt66zyyR5u/Sxejq6s0
7B5M4yWi1OvHDHSk8GAFFAPa2N9yj4v1JMruwg7GlDnwvWdYIvNQZ3rZkBqdg49D
VCTCXdE3vEHxd9w7P9Dxr0eS7FJGV8U+rjuyxJhBkVQAtqAN5YgGdeLjDYysQiDl
OV4pMlRV4Dih5a80+DfA5trYZSOqd5iOEENG4wve/EZbJQtOy30zd5PWQie8Jdgy
1bP2ifD06JttjHBoSDQLZ0DecSewqZclFvl1rfaczRF1a1HrKokS++ebU2X9k1Qt
Fe7KNG2SsB+TUaf7bp9D0Fji9mVe4pEi2YlAtn0TmFj7evoZzq87NN9TTVa79tqY
/5nCV0EIIqFlZlLaP8iAII7AeWnez99l8vSKu3ZVr/dT4drh/+yy+vWtvbmQy7BG
3l9PdjwUXEc9754Szxqzsu64n2QGMMxlOo3UxWLBj+TxYcPXiu0TL5qOOdyYcbcb
SqvUgnxPvy7NZOe0tcWJhVqq43Yg5S88kAHgiVWSNUT2dpvM19fKR+Q1woFIubNM
l2DoOEpxfN6ZbqFO2g2dCSkKfmZHpQ4J3cMsauFWGKuC38/rS8cXnawgoDIrFfbd
TMVj4HfMjljMS914haP6w7XH5PAPWXlbcOeDygsB99IYUWUqu4snETw522atNyxQ
rg7RewWjTlgxu1gMlZkBphxMoRdSohkfMhYi1Ra7NIBXrvZrZpNjxvfSlXiTVOXy
Ba+6STqHaEibDT1R3G7VPP/A9n6LvVURA/YDbT9bJNuqBjXqQRZftlLSFUi+DyHR
j5KDnjSR4bMutHshklT9m9YDoUq5CPD/yUXkgGuld63n15JeWkrVPsMd5UZxc8s/
U4zSqA0nJoJT6DFwEICKit6m678cT+rb95PYzBX8IYP7JxGkHK90qiDpxUQIYd1h
YmdsXHFRD0/cR0Tjuu8FGPEjDqoWyAAZzqLlF3hqyCtl7i5JHjrbiqqW3y5lP7rI
+hRSTSxGJ765xj46cjNN7iqqWwH2r8ZSq5ZXHkVEimkk2sppeIc0ZfVnK03fg6K+
ARxiNaVvPpdmvh5yd9lFEJo72Ed7xHW4YrDVmmwVMw85hzL/oNOZTa4MBFIXxme2
HBVTseYHnvALVBkEY44EC0/uuIm728AWHLq2OtWQoUckYCLIJacWYjeKc/rexhEB
9uPNldUdpY4Td1HFd/4/2k2Q3srWGlNQxHibhT/sLIEyAtW+9PI6Qpu0mnE5Qwzn
x48adiABTlttSoVGzt8Ni27EjV7zXnhoe1g66yBPtNE9SsH4LGrsp+AAh8Rffmvz
J4wjxS6Iek/9XCWm/RubM0L98R+iBm/0QgyPFw3a8Lio4zUD+lOjl/ei6LFogW40
La3PaUTVLhDmUYKQKyIB8vfzRNVR53tDmzwtCfYbd8aUBOSZRtVcRE1CDNcwDBX2
j1lIEXOSLUmeOF+294BkK8JFCCVe3X0ZiMEFQNXJu8eECC1MiBF/GeW/spDwWfy2
o7hIS5tZpdeRZkwIgaAG8hx6L1+MMq11uMiRUxgtzv1aeDNB57fcMtcWjJmltNaf
e7GhLKWYhNmVOzfLjBFyPMBkyG77vcs/jjABkOvoJtbgnjLIS1AAgnLLS7oYXXjc
ALD5rNXNgP9la7uQ8QkhnYk9SE4vFFTUiZdE6v86ttRkalx/nC7bsQCfl8uIhDsd
RoP2docPaNY3OJRwQGKUWGLGA3qLYKmmBOWKuGuwo/McZjAV6mzsyIpQEYBDoC0S
qwMQPA3wC6XMUW4oJ0W3pZ6MkboIGUKxSOOmvCHT9WHyjJNlnULpi8lXqZI9mhmW
QAViGmc4kR6g+qzwBj2Fd6zBiNVvF2YVactk6mGKZNdN7aNzCahib6NwBHDIuRS1
3Y62vzBMinQ7BJjcwuO5M1zmm8Er1TWww8MaBPM+aRhMvcStGQBltA+Q/GblH+Po
1J2lLgH2eV4jTy5trpJHsQ==
`pragma protect end_protected
