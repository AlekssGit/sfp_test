// setup_ddr.v

// Generated using ACDS version 21.4 67

`timescale 1 ps / 1 ps
module setup_ddr (
		output wire [24:0]  amm_addr,                 //   avalon_master.address
		input  wire [255:0] amm_readdata,             //                .readdata
		output wire [255:0] amm_writedata,            //                .writedata
		output wire         amm_read,                 //                .read
		output wire         amm_write,                //                .write
		output wire [31:0]  amm_byteenable,           //                .byteenable
		output wire [6:0]   amm_burstcount,           //                .burstcount
		input  wire         amm_readdatavalid,        //                .readdatavalid
		input  wire         amm_ready,                //                .waitrequest
		output wire         setup_done,               //           setup.setup_done
		input  wire         local_cal_success_avalon, //      ddr_status.local_cal_success
		input  wire         local_cal_fail_avalon,    //                .local_cal_fail
		input  wire         ram_ready,                //       ddr_ready.ram_ready
		input  wire         clk,                      // clock_125_tx_rx.clk
		input  wire         avalon_clk,               //    clock_avalon.clk
		input  wire         clk_50,                   //        clock_50.clk
		input  wire         rst_n,                    //     reset_board.reset
		input  wire         avalon_reset,             //    reset_avalon.reset
		input  wire         reset,                    //    reset_module.reset
		output wire         local_cal_success         //     cal_success.writeresponsevalid_n
	);

	setup_ddr_data_256 setup_ddr (
		.amm_addr                 (amm_addr),                 //  output,   width = 25,   avalon_master.address
		.amm_readdata             (amm_readdata),             //   input,  width = 256,                .readdata
		.amm_writedata            (amm_writedata),            //  output,  width = 256,                .writedata
		.amm_read                 (amm_read),                 //  output,    width = 1,                .read
		.amm_write                (amm_write),                //  output,    width = 1,                .write
		.amm_byteenable           (amm_byteenable),           //  output,   width = 32,                .byteenable
		.amm_burstcount           (amm_burstcount),           //  output,    width = 7,                .burstcount
		.amm_readdatavalid        (amm_readdatavalid),        //   input,    width = 1,                .readdatavalid
		.amm_ready                (amm_ready),                //   input,    width = 1,                .waitrequest
		.setup_done               (setup_done),               //  output,    width = 1,           setup.setup_done
		.local_cal_success_avalon (local_cal_success_avalon), //   input,    width = 1,      ddr_status.local_cal_success
		.local_cal_fail_avalon    (local_cal_fail_avalon),    //   input,    width = 1,                .local_cal_fail
		.ram_ready                (ram_ready),                //   input,    width = 1,       ddr_ready.ram_ready
		.clk                      (clk),                      //   input,    width = 1, clock_125_tx_rx.clk
		.avalon_clk               (avalon_clk),               //   input,    width = 1,    clock_avalon.clk
		.clk_50                   (clk_50),                   //   input,    width = 1,        clock_50.clk
		.rst_n                    (rst_n),                    //   input,    width = 1,     reset_board.reset
		.avalon_reset             (avalon_reset),             //   input,    width = 1,    reset_avalon.reset
		.reset                    (reset),                    //   input,    width = 1,    reset_module.reset
		.local_cal_success        (local_cal_success)         //  output,    width = 1,     cal_success.writeresponsevalid_n
	);

endmodule
