// system_design.v

// Generated using ACDS version 21.3 170

`timescale 1 ps / 1 ps
module system_design (
		output wire        clock_50_clk,                            //                    clock_50.clk
		output wire        ddr_avalon_clk,                          //                  ddr_avalon.clk
		input  wire        ddr3_global_reset_n_reset_n,             //         ddr3_global_reset_n.reset_n
		input  wire        ddr3_clock_clk,                          //                  ddr3_clock.clk
		input  wire        ddr3_oct_oct_rzqin,                      //                    ddr3_oct.oct_rzqin
		output wire [0:0]  ddr3_mem_mem_ck,                         //                    ddr3_mem.mem_ck
		output wire [0:0]  ddr3_mem_mem_ck_n,                       //                            .mem_ck_n
		output wire [14:0] ddr3_mem_mem_a,                          //                            .mem_a
		output wire [2:0]  ddr3_mem_mem_ba,                         //                            .mem_ba
		output wire [0:0]  ddr3_mem_mem_cke,                        //                            .mem_cke
		output wire [0:0]  ddr3_mem_mem_cs_n,                       //                            .mem_cs_n
		output wire [0:0]  ddr3_mem_mem_odt,                        //                            .mem_odt
		output wire [0:0]  ddr3_mem_mem_reset_n,                    //                            .mem_reset_n
		output wire [0:0]  ddr3_mem_mem_we_n,                       //                            .mem_we_n
		output wire [0:0]  ddr3_mem_mem_ras_n,                      //                            .mem_ras_n
		output wire [0:0]  ddr3_mem_mem_cas_n,                      //                            .mem_cas_n
		inout  wire [4:0]  ddr3_mem_mem_dqs,                        //                            .mem_dqs
		inout  wire [4:0]  ddr3_mem_mem_dqs_n,                      //                            .mem_dqs_n
		inout  wire [39:0] ddr3_mem_mem_dq,                         //                            .mem_dq
		output wire [4:0]  ddr3_mem_mem_dm,                         //                            .mem_dm
		output wire        ddr_avalon_reset_reset,                  //            ddr_avalon_reset.reset
		output wire        mac_inited_mac_inited,                   //                  mac_inited.mac_inited
		input  wire        pcie_refclk_clk,                         //                 pcie_refclk.clk
		input  wire        pcie_npor_npor,                          //                   pcie_npor.npor
		input  wire        pcie_npor_pin_perst,                     //                            .pin_perst
		input  wire        pcie_hip_serial_rx_in0,                  //             pcie_hip_serial.rx_in0
		input  wire        pcie_hip_serial_rx_in1,                  //                            .rx_in1
		input  wire        pcie_hip_serial_rx_in2,                  //                            .rx_in2
		input  wire        pcie_hip_serial_rx_in3,                  //                            .rx_in3
		output wire        pcie_hip_serial_tx_out0,                 //                            .tx_out0
		output wire        pcie_hip_serial_tx_out1,                 //                            .tx_out1
		output wire        pcie_hip_serial_tx_out2,                 //                            .tx_out2
		output wire        pcie_hip_serial_tx_out3,                 //                            .tx_out3
		input  wire        pll_refclk_clk,                          //                  pll_refclk.clk
		output wire        receive_packet_1_data_saved_data_saved,  // receive_packet_1_data_saved.data_saved
		output wire        receive_packet_2_data_saved_data_saved,  // receive_packet_2_data_saved.data_saved
		output wire        reset_main_out_reset,                    //              reset_main_out.reset
		input  wire        reset_mod_clock_clk,                     //             reset_mod_clock.clk
		input  wire        reset_mod_reset_reset_n,                 //             reset_mod_reset.reset_n
		output wire        reset_mod_reset_phy_reset,               //         reset_mod_reset_phy.reset
		output wire [5:0]  pcie_send_control_start_ram_addr,        //           pcie_send_control.start_ram_addr
		output wire        pcie_send_control_signal,                //                            .signal
		input  wire [24:0] send_packet_1_control_start_ram_addr,    //       send_packet_1_control.start_ram_addr
		input  wire        send_packet_1_control_cmd_send,          //                            .cmd_send
		input  wire [24:0] send_packet_2_control_start_ram_addr,    //       send_packet_2_control.start_ram_addr
		input  wire        send_packet_2_control_cmd_send,          //                            .cmd_send
		input  wire        ddr_ready_ram_ready,                     //                   ddr_ready.ram_ready
		input  wire        reset_board_reset,                       //                 reset_board.reset
		output wire        mem_cal_success_cal_success,             //             mem_cal_success.cal_success
		output wire        mac_misc_1_magic_wakeup,                 //                  mac_misc_1.magic_wakeup
		input  wire        mac_misc_1_magic_sleep_n,                //                            .magic_sleep_n
		input  wire        mac_misc_1_tx_crc_fwd,                   //                            .tx_crc_fwd
		output wire        mac_mdio_mdc,                            //                    mac_mdio.mdc
		input  wire        mac_mdio_mdio_in,                        //                            .mdio_in
		output wire        mac_mdio_mdio_out,                       //                            .mdio_out
		output wire        mac_mdio_mdio_oen,                       //                            .mdio_oen
		output wire        mac_misc_2_magic_wakeup,                 //                  mac_misc_2.magic_wakeup
		input  wire        mac_misc_2_magic_sleep_n,                //                            .magic_sleep_n
		input  wire        mac_misc_2_tx_crc_fwd,                   //                            .tx_crc_fwd
		input  wire        tse_ref_clk,                             //                     tse_ref.clk
		output wire        status_led_connection_0_crs,             //     status_led_connection_0.crs
		output wire        status_led_connection_0_link,            //                            .link
		output wire        status_led_connection_0_panel_link,      //                            .panel_link
		output wire        status_led_connection_0_col,             //                            .col
		output wire        status_led_connection_0_an,              //                            .an
		output wire        status_led_connection_0_char_err,        //                            .char_err
		output wire        status_led_connection_0_disp_err,        //                            .disp_err
		input  wire [0:0]  tx_analogreset_0_tx_analogreset,         //            tx_analogreset_0.tx_analogreset
		input  wire [0:0]  tx_digitalreset_0_tx_digitalreset,       //           tx_digitalreset_0.tx_digitalreset
		input  wire [0:0]  rx_analogreset_0_rx_analogreset,         //            rx_analogreset_0.rx_analogreset
		input  wire [0:0]  rx_digitalreset_0_rx_digitalreset,       //           rx_digitalreset_0.rx_digitalreset
		output wire [0:0]  tx_cal_busy_0_tx_cal_busy,               //               tx_cal_busy_0.tx_cal_busy
		output wire [0:0]  rx_cal_busy_0_rx_cal_busy,               //               rx_cal_busy_0.rx_cal_busy
		input  wire        tse_rx_cdr_refclk_0_clk,                 //         tse_rx_cdr_refclk_0.clk
		input  wire [0:0]  rx_set_locktodata_0_rx_set_locktodata,   //         rx_set_locktodata_0.rx_set_locktodata
		input  wire [0:0]  rx_set_locktoref_0_rx_set_locktoref,     //          rx_set_locktoref_0.rx_set_locktoref
		output wire [0:0]  rx_is_lockedtoref_0_rx_is_lockedtoref,   //         rx_is_lockedtoref_0.rx_is_lockedtoref
		output wire [0:0]  rx_is_lockedtodata_0_rx_is_lockedtodata, //        rx_is_lockedtodata_0.rx_is_lockedtodata
		input  wire        sgmii_1_rxp,                             //                     sgmii_1.rxp
		output wire        sgmii_1_txp,                             //                            .txp
		output wire        serdes_control_connection_0_export,      // serdes_control_connection_0.export
		output wire        status_led_connection_1_crs,             //     status_led_connection_1.crs
		output wire        status_led_connection_1_link,            //                            .link
		output wire        status_led_connection_1_panel_link,      //                            .panel_link
		output wire        status_led_connection_1_col,             //                            .col
		output wire        status_led_connection_1_an,              //                            .an
		output wire        status_led_connection_1_char_err,        //                            .char_err
		output wire        status_led_connection_1_disp_err,        //                            .disp_err
		input  wire [0:0]  tx_analogreset_1_tx_analogreset,         //            tx_analogreset_1.tx_analogreset
		input  wire [0:0]  tx_digitalreset_1_tx_digitalreset,       //           tx_digitalreset_1.tx_digitalreset
		input  wire [0:0]  rx_analogreset_1_rx_analogreset,         //            rx_analogreset_1.rx_analogreset
		input  wire [0:0]  rx_digitalreset_1_rx_digitalreset,       //           rx_digitalreset_1.rx_digitalreset
		output wire [0:0]  tx_cal_busy_1_tx_cal_busy,               //               tx_cal_busy_1.tx_cal_busy
		output wire [0:0]  rx_cal_busy_1_rx_cal_busy,               //               rx_cal_busy_1.rx_cal_busy
		input  wire        tse_rx_cdr_refclk_1_clk,                 //         tse_rx_cdr_refclk_1.clk
		input  wire [0:0]  rx_set_locktodata_1_rx_set_locktodata,   //         rx_set_locktodata_1.rx_set_locktodata
		input  wire [0:0]  rx_set_locktoref_1_rx_set_locktoref,     //          rx_set_locktoref_1.rx_set_locktoref
		output wire [0:0]  rx_is_lockedtoref_1_rx_is_lockedtoref,   //         rx_is_lockedtoref_1.rx_is_lockedtoref
		output wire [0:0]  rx_is_lockedtodata_1_rx_is_lockedtodata, //        rx_is_lockedtodata_1.rx_is_lockedtodata
		input  wire        sgmii_2_rxp,                             //                     sgmii_2.rxp
		output wire        sgmii_2_txp,                             //                            .txp
		output wire        serdes_control_connection_1_export,      // serdes_control_connection_1.export
		input  wire [0:0]  tse_tx_serial_clk_2_clk,                 //         tse_tx_serial_clk_2.clk
		input  wire        tse_rx_cdr_refclk_2_clk,                 //         tse_rx_cdr_refclk_2.clk
		input  wire        sgmii_3_rxp,                             //                     sgmii_3.rxp
		output wire        sgmii_3_txp,                             //                            .txp
		input  wire [0:0]  tse_tx_serial_clk_3_clk,                 //         tse_tx_serial_clk_3.clk
		input  wire        tse_rx_cdr_refclk_3_clk,                 //         tse_rx_cdr_refclk_3.clk
		input  wire        sgmii_4_rxp,                             //                     sgmii_4.rxp
		output wire        sgmii_4_txp,                             //                            .txp
		input  wire        xcvr_pll_powerdown_pll_powerdown,        //          xcvr_pll_powerdown.pll_powerdown
		input  wire        xcvr_pll_refclk_clk                      //             xcvr_pll_refclk.clk
	);

	wire   [31:0] init_mac_avalon_master_readdata;                            // tse:reg_data_out -> init_mac:DAT_I
	wire          init_mac_avalon_master_waitrequest;                         // tse:reg_busy -> init_mac:BUSY
	wire    [9:0] init_mac_avalon_master_address;                             // init_mac:ADR_O -> tse:reg_addr
	wire          init_mac_avalon_master_read;                                // init_mac:RD -> tse:reg_rd
	wire   [31:0] init_mac_avalon_master_writedata;                           // init_mac:DAT_O -> tse:reg_data_in
	wire          init_mac_avalon_master_write;                               // init_mac:WR -> tse:reg_wr
	wire          send_packet_1_avalon_streaming_source_valid;                // send_packet_1:ff_tx_wren -> tse:data_tx_valid_0
	wire    [7:0] send_packet_1_avalon_streaming_source_data;                 // send_packet_1:ff_tx_data -> tse:data_tx_data_0
	wire          send_packet_1_avalon_streaming_source_ready;                // tse:data_tx_ready_0 -> send_packet_1:ff_tx_rdy
	wire          send_packet_1_avalon_streaming_source_startofpacket;        // send_packet_1:ff_tx_sop -> tse:data_tx_sop_0
	wire          send_packet_1_avalon_streaming_source_endofpacket;          // send_packet_1:ff_tx_eop -> tse:data_tx_eop_0
	wire          send_packet_1_avalon_streaming_source_error;                // send_packet_1:ff_tx_err -> tse:data_tx_error_0
	wire          send_packet_2_avalon_streaming_source_valid;                // send_packet_2:ff_tx_wren -> tse:data_tx_valid_1
	wire    [7:0] send_packet_2_avalon_streaming_source_data;                 // send_packet_2:ff_tx_data -> tse:data_tx_data_1
	wire          send_packet_2_avalon_streaming_source_ready;                // tse:data_tx_ready_1 -> send_packet_2:ff_tx_rdy
	wire          send_packet_2_avalon_streaming_source_startofpacket;        // send_packet_2:ff_tx_sop -> tse:data_tx_sop_1
	wire          send_packet_2_avalon_streaming_source_endofpacket;          // send_packet_2:ff_tx_eop -> tse:data_tx_eop_1
	wire          send_packet_2_avalon_streaming_source_error;                // send_packet_2:ff_tx_err -> tse:data_tx_error_1
	wire          receive_packet_1_fifo_status_valid;                         // receive_packet_1:rx_afull_valid -> tse:rx_afull_valid
	wire    [1:0] receive_packet_1_fifo_status_data;                          // receive_packet_1:rx_afull_data -> tse:rx_afull_data
	wire    [1:0] receive_packet_1_fifo_status_channel;                       // receive_packet_1:rx_afull_channel -> tse:rx_afull_channel
	wire          tse_receive_0_valid;                                        // tse:data_rx_valid_0 -> receive_packet_1:ff_rx_dval
	wire    [7:0] tse_receive_0_data;                                         // tse:data_rx_data_0 -> receive_packet_1:ff_rx_data
	wire          tse_receive_0_ready;                                        // receive_packet_1:ff_rx_rdy -> tse:data_rx_ready_0
	wire          tse_receive_0_startofpacket;                                // tse:data_rx_sop_0 -> receive_packet_1:ff_rx_sop
	wire          tse_receive_0_endofpacket;                                  // tse:data_rx_eop_0 -> receive_packet_1:ff_rx_eop
	wire    [4:0] tse_receive_0_error;                                        // tse:data_rx_error_0 -> receive_packet_1:rx_err
	wire          tse_receive_1_valid;                                        // tse:data_rx_valid_1 -> receive_packet_2:ff_rx_dval
	wire    [7:0] tse_receive_1_data;                                         // tse:data_rx_data_1 -> receive_packet_2:ff_rx_data
	wire          tse_receive_1_ready;                                        // receive_packet_2:ff_rx_rdy -> tse:data_rx_ready_1
	wire          tse_receive_1_startofpacket;                                // tse:data_rx_sop_1 -> receive_packet_2:ff_rx_sop
	wire          tse_receive_1_endofpacket;                                  // tse:data_rx_eop_1 -> receive_packet_2:ff_rx_eop
	wire    [4:0] tse_receive_1_error;                                        // tse:data_rx_error_1 -> receive_packet_2:rx_err
	wire          pcie_coreclkout_hip_clk;                                    // pcie:coreclkout_hip -> [irq_mapper:clk, mm_interconnect_1:pcie_coreclkout_hip_clk, mm_interconnect_6:pcie_coreclkout_hip_clk, send_cmd_pcie:clk]
	wire          ddr3_emif_usr_clk_clk;                                      // ddr3:emif_usr_clk -> [clock_ddr_avalon:in_clk, mm_interconnect_1:ddr3_emif_usr_clk_clk, rst_controller_005:clk, setup_ddr:avalon_clk]
	wire          tse_mac_rx_clock_connection_0_clk;                          // tse:mac_rx_clk_0 -> [mem_rcv_1:clk, mm_interconnect_2:tse_mac_rx_clock_connection_0_clk, receive_packet_1:clk_original, rst_controller_004:clk]
	wire          tse_mac_rx_clock_connection_1_clk;                          // tse:mac_rx_clk_1 -> [mem_4:clk2, mem_rcv_2:clk, mm_interconnect_5:tse_mac_rx_clock_connection_1_clk, receive_packet_2:clk_original, rst_controller_002:clk]
	wire          tse_mac_tx_clock_connection_0_clk;                          // tse:mac_tx_clk_0 -> [mem_5:clk, mm_interconnect_4:tse_mac_tx_clock_connection_0_clk, rst_controller_003:clk, send_packet_1:clk_original]
	wire          tse_mac_tx_clock_connection_1_clk;                          // tse:mac_tx_clk_1 -> [mem_4:clk, mm_interconnect_3:tse_mac_tx_clock_connection_1_clk, rst_controller_001:clk, send_packet_2:clk_original]
	wire          pll_outclk0_clk;                                            // pll:outclk_0 -> [receive_packet_1:fifo_status_clk, setup_ddr:clk, tse:rx_afull_clk]
	wire          pll_outclk1_clk;                                            // pll:outclk_1 -> [clock_50_out:in_clk, init_mac:clk, rst_controller:clk, setup_ddr:clk_50, tse:clk]
	wire          pll_outclk2_clk;                                            // pll:outclk_2 -> receive_packet_2:fifo_status_clk
	wire          send_cmd_pcie_ddr_setup_cmd_ddr_setup_cmd;                  // send_cmd_pcie:ddr_setup_cmd -> setup_ddr:ddr_setup_cmd_pci
	wire          setup_ddr_ddr_status_out_local_cal_fail;                    // setup_ddr:ddr_local_cal_fail -> send_cmd_pcie:ddr_local_cal_fail
	wire          setup_ddr_ddr_status_out_local_cal_success;                 // setup_ddr:ddr_local_cal_success -> send_cmd_pcie:ddr_local_cal_success
	wire          setup_ddr_resets_information_main_reset;                    // setup_ddr:system_main_reset -> send_cmd_pcie:system_main_reset
	wire          setup_ddr_resets_information_board_reset;                   // setup_ddr:board_reset -> send_cmd_pcie:board_reset
	wire          setup_ddr_resets_information_ddr_avalon_reset;              // setup_ddr:ddr_avalon_rst -> send_cmd_pcie:ddr_avalon_rst
	wire          setup_ddr_setup_setup_done;                                 // setup_ddr:setup_done -> send_cmd_pcie:ddr_setup_done
	wire          ddr3_status_local_cal_fail;                                 // ddr3:local_cal_fail -> setup_ddr:local_cal_fail_avalon
	wire          ddr3_status_local_cal_success;                              // ddr3:local_cal_success -> setup_ddr:local_cal_success_avalon
	wire          xcvr_pll_tx_serial_clk_clk;                                 // xcvr_pll:tx_serial_clk -> [tse:tx_serial_clk_0, tse:tx_serial_clk_1]
	wire          pcie_app_nreset_status_reset;                               // pcie:app_nreset_status -> [irq_mapper:reset, mm_interconnect_1:pcie_rxm_bar2_translator_reset_reset_bridge_in_reset_reset, mm_interconnect_6:pcie_rxm_bar0_translator_reset_reset_bridge_in_reset_reset, send_cmd_pcie:rst_n]
	wire          ddr3_emif_usr_reset_n_reset;                                // ddr3:emif_usr_reset_n -> [ddr_avalon_reset:in_reset, rst_controller_005:reset_in0]
	wire          reset_mod_reset_main_reset;                                 // reset_mod:reset -> [pll:rst, reset_main:in_reset, rst_controller:reset_in0, rst_controller_001:reset_in0, rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_004:reset_in0, setup_ddr:reset]
	wire  [255:0] setup_ddr_avalon_master_readdata;                           // mm_interconnect_1:setup_ddr_avalon_master_readdata -> setup_ddr:amm_readdata
	wire          setup_ddr_avalon_master_waitrequest;                        // mm_interconnect_1:setup_ddr_avalon_master_waitrequest -> setup_ddr:amm_ready
	wire   [24:0] setup_ddr_avalon_master_address;                            // setup_ddr:amm_addr -> mm_interconnect_1:setup_ddr_avalon_master_address
	wire          setup_ddr_avalon_master_read;                               // setup_ddr:amm_read -> mm_interconnect_1:setup_ddr_avalon_master_read
	wire   [31:0] setup_ddr_avalon_master_byteenable;                         // setup_ddr:amm_byteenable -> mm_interconnect_1:setup_ddr_avalon_master_byteenable
	wire          setup_ddr_avalon_master_readdatavalid;                      // mm_interconnect_1:setup_ddr_avalon_master_readdatavalid -> setup_ddr:amm_readdatavalid
	wire  [255:0] setup_ddr_avalon_master_writedata;                          // setup_ddr:amm_writedata -> mm_interconnect_1:setup_ddr_avalon_master_writedata
	wire          setup_ddr_avalon_master_write;                              // setup_ddr:amm_write -> mm_interconnect_1:setup_ddr_avalon_master_write
	wire    [6:0] setup_ddr_avalon_master_burstcount;                         // setup_ddr:amm_burstcount -> mm_interconnect_1:setup_ddr_avalon_master_burstcount
	wire  [127:0] pcie_rxm_bar2_readdata;                                     // mm_interconnect_1:pcie_rxm_bar2_readdata -> pcie:rxm_bar2_readdata_i
	wire          pcie_rxm_bar2_waitrequest;                                  // mm_interconnect_1:pcie_rxm_bar2_waitrequest -> pcie:rxm_bar2_waitrequest_i
	wire   [63:0] pcie_rxm_bar2_address;                                      // pcie:rxm_bar2_address_o -> mm_interconnect_1:pcie_rxm_bar2_address
	wire   [15:0] pcie_rxm_bar2_byteenable;                                   // pcie:rxm_bar2_byteenable_o -> mm_interconnect_1:pcie_rxm_bar2_byteenable
	wire          pcie_rxm_bar2_read;                                         // pcie:rxm_bar2_read_o -> mm_interconnect_1:pcie_rxm_bar2_read
	wire          pcie_rxm_bar2_readdatavalid;                                // mm_interconnect_1:pcie_rxm_bar2_readdatavalid -> pcie:rxm_bar2_readdatavalid_i
	wire  [127:0] pcie_rxm_bar2_writedata;                                    // pcie:rxm_bar2_writedata_o -> mm_interconnect_1:pcie_rxm_bar2_writedata
	wire          pcie_rxm_bar2_write;                                        // pcie:rxm_bar2_write_o -> mm_interconnect_1:pcie_rxm_bar2_write
	wire    [5:0] pcie_rxm_bar2_burstcount;                                   // pcie:rxm_bar2_burstcount_o -> mm_interconnect_1:pcie_rxm_bar2_burstcount
	wire  [255:0] mm_interconnect_1_ddr3_ctrl_amm_0_readdata;                 // ddr3:amm_readdata_0 -> mm_interconnect_1:ddr3_ctrl_amm_0_readdata
	wire          mm_interconnect_1_ddr3_ctrl_amm_0_waitrequest;              // ddr3:amm_ready_0 -> mm_interconnect_1:ddr3_ctrl_amm_0_waitrequest
	wire   [24:0] mm_interconnect_1_ddr3_ctrl_amm_0_address;                  // mm_interconnect_1:ddr3_ctrl_amm_0_address -> ddr3:amm_address_0
	wire          mm_interconnect_1_ddr3_ctrl_amm_0_read;                     // mm_interconnect_1:ddr3_ctrl_amm_0_read -> ddr3:amm_read_0
	wire   [31:0] mm_interconnect_1_ddr3_ctrl_amm_0_byteenable;               // mm_interconnect_1:ddr3_ctrl_amm_0_byteenable -> ddr3:amm_byteenable_0
	wire          mm_interconnect_1_ddr3_ctrl_amm_0_readdatavalid;            // ddr3:amm_readdatavalid_0 -> mm_interconnect_1:ddr3_ctrl_amm_0_readdatavalid
	wire          mm_interconnect_1_ddr3_ctrl_amm_0_write;                    // mm_interconnect_1:ddr3_ctrl_amm_0_write -> ddr3:amm_write_0
	wire  [255:0] mm_interconnect_1_ddr3_ctrl_amm_0_writedata;                // mm_interconnect_1:ddr3_ctrl_amm_0_writedata -> ddr3:amm_writedata_0
	wire    [6:0] mm_interconnect_1_ddr3_ctrl_amm_0_burstcount;               // mm_interconnect_1:ddr3_ctrl_amm_0_burstcount -> ddr3:amm_burstcount_0
	wire          receive_packet_1_avalon_master_chipselect;                  // receive_packet_1:ram_chipselect -> mm_interconnect_2:receive_packet_1_avalon_master_chipselect
	wire   [31:0] receive_packet_1_avalon_master_readdata;                    // mm_interconnect_2:receive_packet_1_avalon_master_readdata -> receive_packet_1:ram_readdata
	wire          receive_packet_1_avalon_master_waitrequest;                 // mm_interconnect_2:receive_packet_1_avalon_master_waitrequest -> receive_packet_1:ram_waitrequest
	wire    [9:0] receive_packet_1_avalon_master_address;                     // receive_packet_1:ram_addr -> mm_interconnect_2:receive_packet_1_avalon_master_address
	wire    [3:0] receive_packet_1_avalon_master_byteenable;                  // receive_packet_1:ram_byteenable -> mm_interconnect_2:receive_packet_1_avalon_master_byteenable
	wire          receive_packet_1_avalon_master_write;                       // receive_packet_1:ram_write -> mm_interconnect_2:receive_packet_1_avalon_master_write
	wire   [31:0] receive_packet_1_avalon_master_writedata;                   // receive_packet_1:ram_writedata -> mm_interconnect_2:receive_packet_1_avalon_master_writedata
	wire          mm_interconnect_2_mem_rcv_1_s1_chipselect;                  // mm_interconnect_2:mem_rcv_1_s1_chipselect -> mem_rcv_1:chipselect
	wire   [31:0] mm_interconnect_2_mem_rcv_1_s1_readdata;                    // mem_rcv_1:readdata -> mm_interconnect_2:mem_rcv_1_s1_readdata
	wire    [9:0] mm_interconnect_2_mem_rcv_1_s1_address;                     // mm_interconnect_2:mem_rcv_1_s1_address -> mem_rcv_1:address
	wire    [3:0] mm_interconnect_2_mem_rcv_1_s1_byteenable;                  // mm_interconnect_2:mem_rcv_1_s1_byteenable -> mem_rcv_1:byteenable
	wire          mm_interconnect_2_mem_rcv_1_s1_write;                       // mm_interconnect_2:mem_rcv_1_s1_write -> mem_rcv_1:write
	wire   [31:0] mm_interconnect_2_mem_rcv_1_s1_writedata;                   // mm_interconnect_2:mem_rcv_1_s1_writedata -> mem_rcv_1:writedata
	wire          mm_interconnect_2_mem_rcv_1_s1_clken;                       // mm_interconnect_2:mem_rcv_1_s1_clken -> mem_rcv_1:clken
	wire          send_packet_2_avalon_master_chipselect;                     // send_packet_2:ram_chipselect -> mm_interconnect_3:send_packet_2_avalon_master_chipselect
	wire   [31:0] send_packet_2_avalon_master_readdata;                       // mm_interconnect_3:send_packet_2_avalon_master_readdata -> send_packet_2:ram_readdata
	wire          send_packet_2_avalon_master_waitrequest;                    // mm_interconnect_3:send_packet_2_avalon_master_waitrequest -> send_packet_2:ram_waitrequest
	wire    [9:0] send_packet_2_avalon_master_address;                        // send_packet_2:ram_addr -> mm_interconnect_3:send_packet_2_avalon_master_address
	wire    [3:0] send_packet_2_avalon_master_byteenable;                     // send_packet_2:ram_byteenable -> mm_interconnect_3:send_packet_2_avalon_master_byteenable
	wire          send_packet_2_avalon_master_write;                          // send_packet_2:ram_write -> mm_interconnect_3:send_packet_2_avalon_master_write
	wire   [31:0] send_packet_2_avalon_master_writedata;                      // send_packet_2:ram_writedata -> mm_interconnect_3:send_packet_2_avalon_master_writedata
	wire          mm_interconnect_3_mem_4_s1_chipselect;                      // mm_interconnect_3:mem_4_s1_chipselect -> mem_4:chipselect
	wire   [31:0] mm_interconnect_3_mem_4_s1_readdata;                        // mem_4:readdata -> mm_interconnect_3:mem_4_s1_readdata
	wire    [9:0] mm_interconnect_3_mem_4_s1_address;                         // mm_interconnect_3:mem_4_s1_address -> mem_4:address
	wire    [3:0] mm_interconnect_3_mem_4_s1_byteenable;                      // mm_interconnect_3:mem_4_s1_byteenable -> mem_4:byteenable
	wire          mm_interconnect_3_mem_4_s1_write;                           // mm_interconnect_3:mem_4_s1_write -> mem_4:write
	wire   [31:0] mm_interconnect_3_mem_4_s1_writedata;                       // mm_interconnect_3:mem_4_s1_writedata -> mem_4:writedata
	wire          mm_interconnect_3_mem_4_s1_clken;                           // mm_interconnect_3:mem_4_s1_clken -> mem_4:clken
	wire          send_packet_1_avalon_master_chipselect;                     // send_packet_1:ram_chipselect -> mm_interconnect_4:send_packet_1_avalon_master_chipselect
	wire   [31:0] send_packet_1_avalon_master_readdata;                       // mm_interconnect_4:send_packet_1_avalon_master_readdata -> send_packet_1:ram_readdata
	wire          send_packet_1_avalon_master_waitrequest;                    // mm_interconnect_4:send_packet_1_avalon_master_waitrequest -> send_packet_1:ram_waitrequest
	wire    [9:0] send_packet_1_avalon_master_address;                        // send_packet_1:ram_addr -> mm_interconnect_4:send_packet_1_avalon_master_address
	wire    [3:0] send_packet_1_avalon_master_byteenable;                     // send_packet_1:ram_byteenable -> mm_interconnect_4:send_packet_1_avalon_master_byteenable
	wire          send_packet_1_avalon_master_write;                          // send_packet_1:ram_write -> mm_interconnect_4:send_packet_1_avalon_master_write
	wire   [31:0] send_packet_1_avalon_master_writedata;                      // send_packet_1:ram_writedata -> mm_interconnect_4:send_packet_1_avalon_master_writedata
	wire          mm_interconnect_4_mem_5_s1_chipselect;                      // mm_interconnect_4:mem_5_s1_chipselect -> mem_5:chipselect
	wire   [31:0] mm_interconnect_4_mem_5_s1_readdata;                        // mem_5:readdata -> mm_interconnect_4:mem_5_s1_readdata
	wire    [9:0] mm_interconnect_4_mem_5_s1_address;                         // mm_interconnect_4:mem_5_s1_address -> mem_5:address
	wire    [3:0] mm_interconnect_4_mem_5_s1_byteenable;                      // mm_interconnect_4:mem_5_s1_byteenable -> mem_5:byteenable
	wire          mm_interconnect_4_mem_5_s1_write;                           // mm_interconnect_4:mem_5_s1_write -> mem_5:write
	wire   [31:0] mm_interconnect_4_mem_5_s1_writedata;                       // mm_interconnect_4:mem_5_s1_writedata -> mem_5:writedata
	wire          mm_interconnect_4_mem_5_s1_clken;                           // mm_interconnect_4:mem_5_s1_clken -> mem_5:clken
	wire          receive_packet_2_avalon_master_chipselect;                  // receive_packet_2:ram_chipselect -> mm_interconnect_5:receive_packet_2_avalon_master_chipselect
	wire   [31:0] receive_packet_2_avalon_master_readdata;                    // mm_interconnect_5:receive_packet_2_avalon_master_readdata -> receive_packet_2:ram_readdata
	wire          receive_packet_2_avalon_master_waitrequest;                 // mm_interconnect_5:receive_packet_2_avalon_master_waitrequest -> receive_packet_2:ram_waitrequest
	wire    [9:0] receive_packet_2_avalon_master_address;                     // receive_packet_2:ram_addr -> mm_interconnect_5:receive_packet_2_avalon_master_address
	wire    [3:0] receive_packet_2_avalon_master_byteenable;                  // receive_packet_2:ram_byteenable -> mm_interconnect_5:receive_packet_2_avalon_master_byteenable
	wire          receive_packet_2_avalon_master_write;                       // receive_packet_2:ram_write -> mm_interconnect_5:receive_packet_2_avalon_master_write
	wire   [31:0] receive_packet_2_avalon_master_writedata;                   // receive_packet_2:ram_writedata -> mm_interconnect_5:receive_packet_2_avalon_master_writedata
	wire          mm_interconnect_5_mem_4_s2_chipselect;                      // mm_interconnect_5:mem_4_s2_chipselect -> mem_4:chipselect2
	wire   [31:0] mm_interconnect_5_mem_4_s2_readdata;                        // mem_4:readdata2 -> mm_interconnect_5:mem_4_s2_readdata
	wire    [9:0] mm_interconnect_5_mem_4_s2_address;                         // mm_interconnect_5:mem_4_s2_address -> mem_4:address2
	wire    [3:0] mm_interconnect_5_mem_4_s2_byteenable;                      // mm_interconnect_5:mem_4_s2_byteenable -> mem_4:byteenable2
	wire          mm_interconnect_5_mem_4_s2_write;                           // mm_interconnect_5:mem_4_s2_write -> mem_4:write2
	wire   [31:0] mm_interconnect_5_mem_4_s2_writedata;                       // mm_interconnect_5:mem_4_s2_writedata -> mem_4:writedata2
	wire          mm_interconnect_5_mem_4_s2_clken;                           // mm_interconnect_5:mem_4_s2_clken -> mem_4:clken2
	wire  [127:0] pcie_rxm_bar0_readdata;                                     // mm_interconnect_6:pcie_rxm_bar0_readdata -> pcie:rxm_bar0_readdata_i
	wire          pcie_rxm_bar0_waitrequest;                                  // mm_interconnect_6:pcie_rxm_bar0_waitrequest -> pcie:rxm_bar0_waitrequest_i
	wire   [63:0] pcie_rxm_bar0_address;                                      // pcie:rxm_bar0_address_o -> mm_interconnect_6:pcie_rxm_bar0_address
	wire   [15:0] pcie_rxm_bar0_byteenable;                                   // pcie:rxm_bar0_byteenable_o -> mm_interconnect_6:pcie_rxm_bar0_byteenable
	wire          pcie_rxm_bar0_read;                                         // pcie:rxm_bar0_read_o -> mm_interconnect_6:pcie_rxm_bar0_read
	wire          pcie_rxm_bar0_readdatavalid;                                // mm_interconnect_6:pcie_rxm_bar0_readdatavalid -> pcie:rxm_bar0_readdatavalid_i
	wire  [127:0] pcie_rxm_bar0_writedata;                                    // pcie:rxm_bar0_writedata_o -> mm_interconnect_6:pcie_rxm_bar0_writedata
	wire          pcie_rxm_bar0_write;                                        // pcie:rxm_bar0_write_o -> mm_interconnect_6:pcie_rxm_bar0_write
	wire    [5:0] pcie_rxm_bar0_burstcount;                                   // pcie:rxm_bar0_burstcount_o -> mm_interconnect_6:pcie_rxm_bar0_burstcount
	wire   [31:0] mm_interconnect_6_send_cmd_pcie_avalon_slave_readdata;      // send_cmd_pcie:avalon_mm_read_data -> mm_interconnect_6:send_cmd_pcie_avalon_slave_readdata
	wire   [15:0] mm_interconnect_6_send_cmd_pcie_avalon_slave_address;       // mm_interconnect_6:send_cmd_pcie_avalon_slave_address -> send_cmd_pcie:avalon_mm_addr
	wire          mm_interconnect_6_send_cmd_pcie_avalon_slave_read;          // mm_interconnect_6:send_cmd_pcie_avalon_slave_read -> send_cmd_pcie:avalon_mm_read
	wire          mm_interconnect_6_send_cmd_pcie_avalon_slave_readdatavalid; // send_cmd_pcie:avalon_mm_rd_valid -> mm_interconnect_6:send_cmd_pcie_avalon_slave_readdatavalid
	wire          mm_interconnect_6_send_cmd_pcie_avalon_slave_write;         // mm_interconnect_6:send_cmd_pcie_avalon_slave_write -> send_cmd_pcie:avalon_mm_write
	wire   [31:0] mm_interconnect_6_send_cmd_pcie_avalon_slave_writedata;     // mm_interconnect_6:send_cmd_pcie_avalon_slave_writedata -> send_cmd_pcie:avalon_mm_write_data
	wire   [15:0] pcie_rxm_irq_irq;                                           // irq_mapper:sender_irq -> pcie:rxm_irq_i
	wire          rst_controller_reset_out_reset;                             // rst_controller:reset_out -> [init_mac:reset, tse:reset]
	wire          rst_controller_001_reset_out_reset;                         // rst_controller_001:reset_out -> [mem_4:reset, mm_interconnect_3:send_packet_2_reset_reset_bridge_in_reset_reset, send_packet_2:rst]
	wire          rst_controller_001_reset_out_reset_req;                     // rst_controller_001:reset_req -> [mem_4:reset_req, rst_translator:reset_req_in]
	wire          rst_controller_002_reset_out_reset;                         // rst_controller_002:reset_out -> [mem_4:reset2, mem_rcv_2:reset, mm_interconnect_5:receive_packet_2_reset_reset_bridge_in_reset_reset, receive_packet_2:rst]
	wire          rst_controller_002_reset_out_reset_req;                     // rst_controller_002:reset_req -> [mem_4:reset_req2, mem_rcv_2:reset_req, rst_translator_001:reset_req_in]
	wire          rst_controller_003_reset_out_reset;                         // rst_controller_003:reset_out -> [mem_5:reset, mm_interconnect_4:send_packet_1_reset_reset_bridge_in_reset_reset, send_packet_1:rst]
	wire          rst_controller_003_reset_out_reset_req;                     // rst_controller_003:reset_req -> [mem_5:reset_req, rst_translator_002:reset_req_in]
	wire          rst_controller_004_reset_out_reset;                         // rst_controller_004:reset_out -> [mem_rcv_1:reset, mm_interconnect_2:receive_packet_1_reset_reset_bridge_in_reset_reset, receive_packet_1:rst]
	wire          rst_controller_004_reset_out_reset_req;                     // rst_controller_004:reset_req -> [mem_rcv_1:reset_req, rst_translator_003:reset_req_in]
	wire          rst_controller_005_reset_out_reset;                         // rst_controller_005:reset_out -> [mm_interconnect_1:setup_ddr_reset_avalon_reset_bridge_in_reset_reset, setup_ddr:avalon_reset]

	clock_50_out clock_50_out (
		.in_clk  (pll_outclk1_clk), //   input,  width = 1,  in_clk.clk
		.out_clk (clock_50_clk)     //  output,  width = 1, out_clk.clk
	);

	clock_ddr_avalon clock_ddr_avalon (
		.in_clk  (ddr3_emif_usr_clk_clk), //   input,  width = 1,  in_clk.clk
		.out_clk (ddr_avalon_clk)         //  output,  width = 1, out_clk.clk
	);

	ddr3 ddr3 (
		.global_reset_n            (ddr3_global_reset_n_reset_n),                     //   input,    width = 1,            global_reset_n.reset_n
		.pll_ref_clk               (ddr3_clock_clk),                                  //   input,    width = 1,               pll_ref_clk.clk
		.oct_rzqin                 (ddr3_oct_oct_rzqin),                              //   input,    width = 1,                       oct.oct_rzqin
		.mem_ck                    (ddr3_mem_mem_ck),                                 //  output,    width = 1,                       mem.mem_ck
		.mem_ck_n                  (ddr3_mem_mem_ck_n),                               //  output,    width = 1,                          .mem_ck_n
		.mem_a                     (ddr3_mem_mem_a),                                  //  output,   width = 15,                          .mem_a
		.mem_ba                    (ddr3_mem_mem_ba),                                 //  output,    width = 3,                          .mem_ba
		.mem_cke                   (ddr3_mem_mem_cke),                                //  output,    width = 1,                          .mem_cke
		.mem_cs_n                  (ddr3_mem_mem_cs_n),                               //  output,    width = 1,                          .mem_cs_n
		.mem_odt                   (ddr3_mem_mem_odt),                                //  output,    width = 1,                          .mem_odt
		.mem_reset_n               (ddr3_mem_mem_reset_n),                            //  output,    width = 1,                          .mem_reset_n
		.mem_we_n                  (ddr3_mem_mem_we_n),                               //  output,    width = 1,                          .mem_we_n
		.mem_ras_n                 (ddr3_mem_mem_ras_n),                              //  output,    width = 1,                          .mem_ras_n
		.mem_cas_n                 (ddr3_mem_mem_cas_n),                              //  output,    width = 1,                          .mem_cas_n
		.mem_dqs                   (ddr3_mem_mem_dqs),                                //   inout,    width = 5,                          .mem_dqs
		.mem_dqs_n                 (ddr3_mem_mem_dqs_n),                              //   inout,    width = 5,                          .mem_dqs_n
		.mem_dq                    (ddr3_mem_mem_dq),                                 //   inout,   width = 40,                          .mem_dq
		.mem_dm                    (ddr3_mem_mem_dm),                                 //  output,    width = 5,                          .mem_dm
		.local_cal_success         (ddr3_status_local_cal_success),                   //  output,    width = 1,                    status.local_cal_success
		.local_cal_fail            (ddr3_status_local_cal_fail),                      //  output,    width = 1,                          .local_cal_fail
		.emif_usr_reset_n          (ddr3_emif_usr_reset_n_reset),                     //  output,    width = 1,          emif_usr_reset_n.reset_n
		.emif_usr_clk              (ddr3_emif_usr_clk_clk),                           //  output,    width = 1,              emif_usr_clk.clk
		.ctrl_ecc_user_interrupt_0 (),                                                //  output,    width = 1, ctrl_ecc_user_interrupt_0.ctrl_ecc_user_interrupt
		.amm_ready_0               (mm_interconnect_1_ddr3_ctrl_amm_0_waitrequest),   //  output,    width = 1,                ctrl_amm_0.waitrequest_n
		.amm_read_0                (mm_interconnect_1_ddr3_ctrl_amm_0_read),          //   input,    width = 1,                          .read
		.amm_write_0               (mm_interconnect_1_ddr3_ctrl_amm_0_write),         //   input,    width = 1,                          .write
		.amm_address_0             (mm_interconnect_1_ddr3_ctrl_amm_0_address),       //   input,   width = 25,                          .address
		.amm_readdata_0            (mm_interconnect_1_ddr3_ctrl_amm_0_readdata),      //  output,  width = 256,                          .readdata
		.amm_writedata_0           (mm_interconnect_1_ddr3_ctrl_amm_0_writedata),     //   input,  width = 256,                          .writedata
		.amm_burstcount_0          (mm_interconnect_1_ddr3_ctrl_amm_0_burstcount),    //   input,    width = 7,                          .burstcount
		.amm_byteenable_0          (mm_interconnect_1_ddr3_ctrl_amm_0_byteenable),    //   input,   width = 32,                          .byteenable
		.amm_readdatavalid_0       (mm_interconnect_1_ddr3_ctrl_amm_0_readdatavalid)  //  output,    width = 1,                          .readdatavalid
	);

	ddr_avalon_reset ddr_avalon_reset (
		.in_reset  (~ddr3_emif_usr_reset_n_reset), //   input,  width = 1,  in_reset.reset
		.out_reset (ddr_avalon_reset_reset)        //  output,  width = 1, out_reset.reset
	);

	init_mac init_mac (
		.clk        (pll_outclk1_clk),                    //   input,   width = 1,         clock.clk
		.reset      (rst_controller_reset_out_reset),     //   input,   width = 1,         reset.reset
		.ADR_O      (init_mac_avalon_master_address),     //  output,  width = 10, avalon_master.address
		.DAT_I      (init_mac_avalon_master_readdata),    //   input,  width = 32,              .readdata
		.DAT_O      (init_mac_avalon_master_writedata),   //  output,  width = 32,              .writedata
		.RD         (init_mac_avalon_master_read),        //  output,   width = 1,              .read
		.WR         (init_mac_avalon_master_write),       //  output,   width = 1,              .write
		.BUSY       (init_mac_avalon_master_waitrequest), //   input,   width = 1,              .waitrequest
		.mac_inited (mac_inited_mac_inited)               //  output,   width = 1,    mac_inited.mac_inited
	);

	mem_4 mem_4 (
		.clk         (tse_mac_tx_clock_connection_1_clk),      //   input,   width = 1,   clk1.clk
		.address     (mm_interconnect_3_mem_4_s1_address),     //   input,  width = 10,     s1.address
		.clken       (mm_interconnect_3_mem_4_s1_clken),       //   input,   width = 1,       .clken
		.chipselect  (mm_interconnect_3_mem_4_s1_chipselect),  //   input,   width = 1,       .chipselect
		.write       (mm_interconnect_3_mem_4_s1_write),       //   input,   width = 1,       .write
		.readdata    (mm_interconnect_3_mem_4_s1_readdata),    //  output,  width = 32,       .readdata
		.writedata   (mm_interconnect_3_mem_4_s1_writedata),   //   input,  width = 32,       .writedata
		.byteenable  (mm_interconnect_3_mem_4_s1_byteenable),  //   input,   width = 4,       .byteenable
		.reset       (rst_controller_001_reset_out_reset),     //   input,   width = 1, reset1.reset
		.reset_req   (rst_controller_001_reset_out_reset_req), //   input,   width = 1,       .reset_req
		.address2    (mm_interconnect_5_mem_4_s2_address),     //   input,  width = 10,     s2.address
		.chipselect2 (mm_interconnect_5_mem_4_s2_chipselect),  //   input,   width = 1,       .chipselect
		.clken2      (mm_interconnect_5_mem_4_s2_clken),       //   input,   width = 1,       .clken
		.write2      (mm_interconnect_5_mem_4_s2_write),       //   input,   width = 1,       .write
		.readdata2   (mm_interconnect_5_mem_4_s2_readdata),    //  output,  width = 32,       .readdata
		.writedata2  (mm_interconnect_5_mem_4_s2_writedata),   //   input,  width = 32,       .writedata
		.byteenable2 (mm_interconnect_5_mem_4_s2_byteenable),  //   input,   width = 4,       .byteenable
		.clk2        (tse_mac_rx_clock_connection_1_clk),      //   input,   width = 1,   clk2.clk
		.reset2      (rst_controller_002_reset_out_reset),     //   input,   width = 1, reset2.reset
		.reset_req2  (rst_controller_002_reset_out_reset_req)  //   input,   width = 1,       .reset_req
	);

	mem_5 mem_5 (
		.clk        (tse_mac_tx_clock_connection_0_clk),      //   input,   width = 1,   clk1.clk
		.address    (mm_interconnect_4_mem_5_s1_address),     //   input,  width = 10,     s1.address
		.clken      (mm_interconnect_4_mem_5_s1_clken),       //   input,   width = 1,       .clken
		.chipselect (mm_interconnect_4_mem_5_s1_chipselect),  //   input,   width = 1,       .chipselect
		.write      (mm_interconnect_4_mem_5_s1_write),       //   input,   width = 1,       .write
		.readdata   (mm_interconnect_4_mem_5_s1_readdata),    //  output,  width = 32,       .readdata
		.writedata  (mm_interconnect_4_mem_5_s1_writedata),   //   input,  width = 32,       .writedata
		.byteenable (mm_interconnect_4_mem_5_s1_byteenable),  //   input,   width = 4,       .byteenable
		.reset      (rst_controller_003_reset_out_reset),     //   input,   width = 1, reset1.reset
		.reset_req  (rst_controller_003_reset_out_reset_req)  //   input,   width = 1,       .reset_req
	);

	mem_3 mem_rcv_1 (
		.clk        (tse_mac_rx_clock_connection_0_clk),         //   input,   width = 1,   clk1.clk
		.address    (mm_interconnect_2_mem_rcv_1_s1_address),    //   input,  width = 10,     s1.address
		.clken      (mm_interconnect_2_mem_rcv_1_s1_clken),      //   input,   width = 1,       .clken
		.chipselect (mm_interconnect_2_mem_rcv_1_s1_chipselect), //   input,   width = 1,       .chipselect
		.write      (mm_interconnect_2_mem_rcv_1_s1_write),      //   input,   width = 1,       .write
		.readdata   (mm_interconnect_2_mem_rcv_1_s1_readdata),   //  output,  width = 32,       .readdata
		.writedata  (mm_interconnect_2_mem_rcv_1_s1_writedata),  //   input,  width = 32,       .writedata
		.byteenable (mm_interconnect_2_mem_rcv_1_s1_byteenable), //   input,   width = 4,       .byteenable
		.reset      (rst_controller_004_reset_out_reset),        //   input,   width = 1, reset1.reset
		.reset_req  (rst_controller_004_reset_out_reset_req)     //   input,   width = 1,       .reset_req
	);

	mem_rcv_0 mem_rcv_2 (
		.clk        (tse_mac_rx_clock_connection_1_clk),      //   input,   width = 1,   clk1.clk
		.address    (),                                       //   input,  width = 10,     s1.address
		.clken      (),                                       //   input,   width = 1,       .clken
		.chipselect (),                                       //   input,   width = 1,       .chipselect
		.write      (),                                       //   input,   width = 1,       .write
		.readdata   (),                                       //  output,  width = 32,       .readdata
		.writedata  (),                                       //   input,  width = 32,       .writedata
		.byteenable (),                                       //   input,   width = 4,       .byteenable
		.reset      (rst_controller_002_reset_out_reset),     //   input,   width = 1, reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req)  //   input,   width = 1,       .reset_req
	);

	pcie pcie (
		.coreclkout_hip           (pcie_coreclkout_hip_clk),      //  output,    width = 1,    coreclkout_hip.clk
		.refclk                   (pcie_refclk_clk),              //   input,    width = 1,            refclk.clk
		.npor                     (pcie_npor_npor),               //   input,    width = 1,              npor.npor
		.pin_perst                (pcie_npor_pin_perst),          //   input,    width = 1,                  .pin_perst
		.app_nreset_status        (pcie_app_nreset_status_reset), //  output,    width = 1, app_nreset_status.reset_n
		.test_in                  (),                             //   input,   width = 32,          hip_ctrl.test_in
		.simu_mode_pipe           (),                             //   input,    width = 1,                  .simu_mode_pipe
		.sim_pipe_pclk_in         (),                             //   input,    width = 1,          hip_pipe.sim_pipe_pclk_in
		.sim_pipe_rate            (),                             //  output,    width = 2,                  .sim_pipe_rate
		.sim_ltssmstate           (),                             //  output,    width = 5,                  .sim_ltssmstate
		.eidleinfersel0           (),                             //  output,    width = 3,                  .eidleinfersel0
		.eidleinfersel1           (),                             //  output,    width = 3,                  .eidleinfersel1
		.eidleinfersel2           (),                             //  output,    width = 3,                  .eidleinfersel2
		.eidleinfersel3           (),                             //  output,    width = 3,                  .eidleinfersel3
		.powerdown0               (),                             //  output,    width = 2,                  .powerdown0
		.powerdown1               (),                             //  output,    width = 2,                  .powerdown1
		.powerdown2               (),                             //  output,    width = 2,                  .powerdown2
		.powerdown3               (),                             //  output,    width = 2,                  .powerdown3
		.rxpolarity0              (),                             //  output,    width = 1,                  .rxpolarity0
		.rxpolarity1              (),                             //  output,    width = 1,                  .rxpolarity1
		.rxpolarity2              (),                             //  output,    width = 1,                  .rxpolarity2
		.rxpolarity3              (),                             //  output,    width = 1,                  .rxpolarity3
		.txcompl0                 (),                             //  output,    width = 1,                  .txcompl0
		.txcompl1                 (),                             //  output,    width = 1,                  .txcompl1
		.txcompl2                 (),                             //  output,    width = 1,                  .txcompl2
		.txcompl3                 (),                             //  output,    width = 1,                  .txcompl3
		.txdata0                  (),                             //  output,   width = 32,                  .txdata0
		.txdata1                  (),                             //  output,   width = 32,                  .txdata1
		.txdata2                  (),                             //  output,   width = 32,                  .txdata2
		.txdata3                  (),                             //  output,   width = 32,                  .txdata3
		.txdatak0                 (),                             //  output,    width = 4,                  .txdatak0
		.txdatak1                 (),                             //  output,    width = 4,                  .txdatak1
		.txdatak2                 (),                             //  output,    width = 4,                  .txdatak2
		.txdatak3                 (),                             //  output,    width = 4,                  .txdatak3
		.txdetectrx0              (),                             //  output,    width = 1,                  .txdetectrx0
		.txdetectrx1              (),                             //  output,    width = 1,                  .txdetectrx1
		.txdetectrx2              (),                             //  output,    width = 1,                  .txdetectrx2
		.txdetectrx3              (),                             //  output,    width = 1,                  .txdetectrx3
		.txelecidle0              (),                             //  output,    width = 1,                  .txelecidle0
		.txelecidle1              (),                             //  output,    width = 1,                  .txelecidle1
		.txelecidle2              (),                             //  output,    width = 1,                  .txelecidle2
		.txelecidle3              (),                             //  output,    width = 1,                  .txelecidle3
		.txdeemph0                (),                             //  output,    width = 1,                  .txdeemph0
		.txdeemph1                (),                             //  output,    width = 1,                  .txdeemph1
		.txdeemph2                (),                             //  output,    width = 1,                  .txdeemph2
		.txdeemph3                (),                             //  output,    width = 1,                  .txdeemph3
		.txmargin0                (),                             //  output,    width = 3,                  .txmargin0
		.txmargin1                (),                             //  output,    width = 3,                  .txmargin1
		.txmargin2                (),                             //  output,    width = 3,                  .txmargin2
		.txmargin3                (),                             //  output,    width = 3,                  .txmargin3
		.txswing0                 (),                             //  output,    width = 1,                  .txswing0
		.txswing1                 (),                             //  output,    width = 1,                  .txswing1
		.txswing2                 (),                             //  output,    width = 1,                  .txswing2
		.txswing3                 (),                             //  output,    width = 1,                  .txswing3
		.phystatus0               (),                             //   input,    width = 1,                  .phystatus0
		.phystatus1               (),                             //   input,    width = 1,                  .phystatus1
		.phystatus2               (),                             //   input,    width = 1,                  .phystatus2
		.phystatus3               (),                             //   input,    width = 1,                  .phystatus3
		.rxdata0                  (),                             //   input,   width = 32,                  .rxdata0
		.rxdata1                  (),                             //   input,   width = 32,                  .rxdata1
		.rxdata2                  (),                             //   input,   width = 32,                  .rxdata2
		.rxdata3                  (),                             //   input,   width = 32,                  .rxdata3
		.rxdatak0                 (),                             //   input,    width = 4,                  .rxdatak0
		.rxdatak1                 (),                             //   input,    width = 4,                  .rxdatak1
		.rxdatak2                 (),                             //   input,    width = 4,                  .rxdatak2
		.rxdatak3                 (),                             //   input,    width = 4,                  .rxdatak3
		.rxelecidle0              (),                             //   input,    width = 1,                  .rxelecidle0
		.rxelecidle1              (),                             //   input,    width = 1,                  .rxelecidle1
		.rxelecidle2              (),                             //   input,    width = 1,                  .rxelecidle2
		.rxelecidle3              (),                             //   input,    width = 1,                  .rxelecidle3
		.rxstatus0                (),                             //   input,    width = 3,                  .rxstatus0
		.rxstatus1                (),                             //   input,    width = 3,                  .rxstatus1
		.rxstatus2                (),                             //   input,    width = 3,                  .rxstatus2
		.rxstatus3                (),                             //   input,    width = 3,                  .rxstatus3
		.rxvalid0                 (),                             //   input,    width = 1,                  .rxvalid0
		.rxvalid1                 (),                             //   input,    width = 1,                  .rxvalid1
		.rxvalid2                 (),                             //   input,    width = 1,                  .rxvalid2
		.rxvalid3                 (),                             //   input,    width = 1,                  .rxvalid3
		.rxdataskip0              (),                             //   input,    width = 1,                  .rxdataskip0
		.rxdataskip1              (),                             //   input,    width = 1,                  .rxdataskip1
		.rxdataskip2              (),                             //   input,    width = 1,                  .rxdataskip2
		.rxdataskip3              (),                             //   input,    width = 1,                  .rxdataskip3
		.rxblkst0                 (),                             //   input,    width = 1,                  .rxblkst0
		.rxblkst1                 (),                             //   input,    width = 1,                  .rxblkst1
		.rxblkst2                 (),                             //   input,    width = 1,                  .rxblkst2
		.rxblkst3                 (),                             //   input,    width = 1,                  .rxblkst3
		.rxsynchd0                (),                             //   input,    width = 2,                  .rxsynchd0
		.rxsynchd1                (),                             //   input,    width = 2,                  .rxsynchd1
		.rxsynchd2                (),                             //   input,    width = 2,                  .rxsynchd2
		.rxsynchd3                (),                             //   input,    width = 2,                  .rxsynchd3
		.currentcoeff0            (),                             //  output,   width = 18,                  .currentcoeff0
		.currentcoeff1            (),                             //  output,   width = 18,                  .currentcoeff1
		.currentcoeff2            (),                             //  output,   width = 18,                  .currentcoeff2
		.currentcoeff3            (),                             //  output,   width = 18,                  .currentcoeff3
		.currentrxpreset0         (),                             //  output,    width = 3,                  .currentrxpreset0
		.currentrxpreset1         (),                             //  output,    width = 3,                  .currentrxpreset1
		.currentrxpreset2         (),                             //  output,    width = 3,                  .currentrxpreset2
		.currentrxpreset3         (),                             //  output,    width = 3,                  .currentrxpreset3
		.txsynchd0                (),                             //  output,    width = 2,                  .txsynchd0
		.txsynchd1                (),                             //  output,    width = 2,                  .txsynchd1
		.txsynchd2                (),                             //  output,    width = 2,                  .txsynchd2
		.txsynchd3                (),                             //  output,    width = 2,                  .txsynchd3
		.txblkst0                 (),                             //  output,    width = 1,                  .txblkst0
		.txblkst1                 (),                             //  output,    width = 1,                  .txblkst1
		.txblkst2                 (),                             //  output,    width = 1,                  .txblkst2
		.txblkst3                 (),                             //  output,    width = 1,                  .txblkst3
		.txdataskip0              (),                             //  output,    width = 1,                  .txdataskip0
		.txdataskip1              (),                             //  output,    width = 1,                  .txdataskip1
		.txdataskip2              (),                             //  output,    width = 1,                  .txdataskip2
		.txdataskip3              (),                             //  output,    width = 1,                  .txdataskip3
		.rate0                    (),                             //  output,    width = 2,                  .rate0
		.rate1                    (),                             //  output,    width = 2,                  .rate1
		.rate2                    (),                             //  output,    width = 2,                  .rate2
		.rate3                    (),                             //  output,    width = 2,                  .rate3
		.rx_in0                   (pcie_hip_serial_rx_in0),       //   input,    width = 1,        hip_serial.rx_in0
		.rx_in1                   (pcie_hip_serial_rx_in1),       //   input,    width = 1,                  .rx_in1
		.rx_in2                   (pcie_hip_serial_rx_in2),       //   input,    width = 1,                  .rx_in2
		.rx_in3                   (pcie_hip_serial_rx_in3),       //   input,    width = 1,                  .rx_in3
		.tx_out0                  (pcie_hip_serial_tx_out0),      //  output,    width = 1,                  .tx_out0
		.tx_out1                  (pcie_hip_serial_tx_out1),      //  output,    width = 1,                  .tx_out1
		.tx_out2                  (pcie_hip_serial_tx_out2),      //  output,    width = 1,                  .tx_out2
		.tx_out3                  (pcie_hip_serial_tx_out3),      //  output,    width = 1,                  .tx_out3
		.msi_intfc_o              (),                             //  output,   width = 82,         msi_intfc.msi_intfc
		.msi_control_o            (),                             //  output,   width = 16,       msi_control.msi_control
		.msix_intfc_o             (),                             //  output,   width = 16,        msix_intfc.msix_intfc
		.intx_req_i               (),                             //   input,    width = 1,        intx_intfc.intx_req
		.intx_ack_o               (),                             //  output,    width = 1,                  .intx_ack
		.txs_address_i            (),                             //   input,   width = 64,               txs.address
		.txs_chipselect_i         (),                             //   input,    width = 1,                  .chipselect
		.txs_byteenable_i         (),                             //   input,   width = 16,                  .byteenable
		.txs_readdata_o           (),                             //  output,  width = 128,                  .readdata
		.txs_writedata_i          (),                             //   input,  width = 128,                  .writedata
		.txs_read_i               (),                             //   input,    width = 1,                  .read
		.txs_write_i              (),                             //   input,    width = 1,                  .write
		.txs_burstcount_i         (),                             //   input,    width = 6,                  .burstcount
		.txs_readdatavalid_o      (),                             //  output,    width = 1,                  .readdatavalid
		.txs_waitrequest_o        (),                             //  output,    width = 1,                  .waitrequest
		.cra_chipselect_i         (),                             //   input,    width = 1,               cra.chipselect
		.cra_address_i            (),                             //   input,   width = 14,                  .address
		.cra_byteenable_i         (),                             //   input,    width = 4,                  .byteenable
		.cra_read_i               (),                             //   input,    width = 1,                  .read
		.cra_readdata_o           (),                             //  output,   width = 32,                  .readdata
		.cra_write_i              (),                             //   input,    width = 1,                  .write
		.cra_writedata_i          (),                             //   input,   width = 32,                  .writedata
		.cra_waitrequest_o        (),                             //  output,    width = 1,                  .waitrequest
		.cra_irq_o                (),                             //  output,    width = 1,           cra_irq.irq
		.rxm_bar0_address_o       (pcie_rxm_bar0_address),        //  output,   width = 64,          rxm_bar0.address
		.rxm_bar0_byteenable_o    (pcie_rxm_bar0_byteenable),     //  output,   width = 16,                  .byteenable
		.rxm_bar0_readdata_i      (pcie_rxm_bar0_readdata),       //   input,  width = 128,                  .readdata
		.rxm_bar0_writedata_o     (pcie_rxm_bar0_writedata),      //  output,  width = 128,                  .writedata
		.rxm_bar0_read_o          (pcie_rxm_bar0_read),           //  output,    width = 1,                  .read
		.rxm_bar0_write_o         (pcie_rxm_bar0_write),          //  output,    width = 1,                  .write
		.rxm_bar0_burstcount_o    (pcie_rxm_bar0_burstcount),     //  output,    width = 6,                  .burstcount
		.rxm_bar0_readdatavalid_i (pcie_rxm_bar0_readdatavalid),  //   input,    width = 1,                  .readdatavalid
		.rxm_bar0_waitrequest_i   (pcie_rxm_bar0_waitrequest),    //   input,    width = 1,                  .waitrequest
		.rxm_bar2_address_o       (pcie_rxm_bar2_address),        //  output,   width = 64,          rxm_bar2.address
		.rxm_bar2_byteenable_o    (pcie_rxm_bar2_byteenable),     //  output,   width = 16,                  .byteenable
		.rxm_bar2_readdata_i      (pcie_rxm_bar2_readdata),       //   input,  width = 128,                  .readdata
		.rxm_bar2_writedata_o     (pcie_rxm_bar2_writedata),      //  output,  width = 128,                  .writedata
		.rxm_bar2_read_o          (pcie_rxm_bar2_read),           //  output,    width = 1,                  .read
		.rxm_bar2_write_o         (pcie_rxm_bar2_write),          //  output,    width = 1,                  .write
		.rxm_bar2_burstcount_o    (pcie_rxm_bar2_burstcount),     //  output,    width = 6,                  .burstcount
		.rxm_bar2_readdatavalid_i (pcie_rxm_bar2_readdatavalid),  //   input,    width = 1,                  .readdatavalid
		.rxm_bar2_waitrequest_i   (pcie_rxm_bar2_waitrequest),    //   input,    width = 1,                  .waitrequest
		.rxm_irq_i                (pcie_rxm_irq_irq)              //   input,   width = 16,           rxm_irq.irq
	);

	pll pll (
		.rst      (reset_mod_reset_main_reset), //   input,  width = 1,   reset.reset
		.refclk   (pll_refclk_clk),             //   input,  width = 1,  refclk.clk
		.outclk_0 (pll_outclk0_clk),            //  output,  width = 1, outclk0.clk
		.outclk_1 (pll_outclk1_clk),            //  output,  width = 1, outclk1.clk
		.outclk_2 (pll_outclk2_clk),            //  output,  width = 1, outclk2.clk
		.outclk_3 ()                            //  output,  width = 1, outclk3.clk
	);

	receive_packet_1 receive_packet_1 (
		.ff_rx_data       (tse_receive_0_data),                         //   input,   width = 8, avalon_streaming_sink.data
		.ff_rx_eop        (tse_receive_0_endofpacket),                  //   input,   width = 1,                      .endofpacket
		.ff_rx_rdy        (tse_receive_0_ready),                        //  output,   width = 1,                      .ready
		.ff_rx_sop        (tse_receive_0_startofpacket),                //   input,   width = 1,                      .startofpacket
		.ff_rx_dval       (tse_receive_0_valid),                        //   input,   width = 1,                      .valid
		.rx_err           (tse_receive_0_error),                        //   input,   width = 5,                      .error
		.ram_addr         (receive_packet_1_avalon_master_address),     //  output,  width = 10,         avalon_master.address
		.ram_chipselect   (receive_packet_1_avalon_master_chipselect),  //  output,   width = 1,                      .chipselect
		.ram_write        (receive_packet_1_avalon_master_write),       //  output,   width = 1,                      .write
		.ram_readdata     (receive_packet_1_avalon_master_readdata),    //   input,  width = 32,                      .readdata
		.ram_writedata    (receive_packet_1_avalon_master_writedata),   //  output,  width = 32,                      .writedata
		.ram_byteenable   (receive_packet_1_avalon_master_byteenable),  //  output,   width = 4,                      .byteenable
		.ram_waitrequest  (receive_packet_1_avalon_master_waitrequest), //   input,   width = 1,                      .waitrequest
		.clk_original     (tse_mac_rx_clock_connection_0_clk),          //   input,   width = 1,                 clock.clk
		.rst              (rst_controller_004_reset_out_reset),         //   input,   width = 1,                 reset.reset
		.rx_afull_data    (receive_packet_1_fifo_status_data),          //  output,   width = 2,           fifo_status.data
		.rx_afull_valid   (receive_packet_1_fifo_status_valid),         //  output,   width = 1,                      .valid
		.rx_afull_channel (receive_packet_1_fifo_status_channel),       //  output,   width = 2,                      .channel
		.fifo_status_clk  (pll_outclk0_clk),                            //   input,   width = 1,       fifo_status_clk.clk
		.data_saved       (receive_packet_1_data_saved_data_saved)      //  output,   width = 1,            data_saved.data_saved
	);

	receive_packet_0 receive_packet_2 (
		.ff_rx_data       (tse_receive_1_data),                         //   input,   width = 8, avalon_streaming_sink.data
		.ff_rx_eop        (tse_receive_1_endofpacket),                  //   input,   width = 1,                      .endofpacket
		.ff_rx_rdy        (tse_receive_1_ready),                        //  output,   width = 1,                      .ready
		.ff_rx_sop        (tse_receive_1_startofpacket),                //   input,   width = 1,                      .startofpacket
		.ff_rx_dval       (tse_receive_1_valid),                        //   input,   width = 1,                      .valid
		.rx_err           (tse_receive_1_error),                        //   input,   width = 5,                      .error
		.ram_addr         (receive_packet_2_avalon_master_address),     //  output,  width = 10,         avalon_master.address
		.ram_chipselect   (receive_packet_2_avalon_master_chipselect),  //  output,   width = 1,                      .chipselect
		.ram_write        (receive_packet_2_avalon_master_write),       //  output,   width = 1,                      .write
		.ram_readdata     (receive_packet_2_avalon_master_readdata),    //   input,  width = 32,                      .readdata
		.ram_writedata    (receive_packet_2_avalon_master_writedata),   //  output,  width = 32,                      .writedata
		.ram_byteenable   (receive_packet_2_avalon_master_byteenable),  //  output,   width = 4,                      .byteenable
		.ram_waitrequest  (receive_packet_2_avalon_master_waitrequest), //   input,   width = 1,                      .waitrequest
		.clk_original     (tse_mac_rx_clock_connection_1_clk),          //   input,   width = 1,                 clock.clk
		.rst              (rst_controller_002_reset_out_reset),         //   input,   width = 1,                 reset.reset
		.rx_afull_data    (),                                           //  output,   width = 2,           fifo_status.data
		.rx_afull_valid   (),                                           //  output,   width = 1,                      .valid
		.rx_afull_channel (),                                           //  output,   width = 2,                      .channel
		.fifo_status_clk  (pll_outclk2_clk),                            //   input,   width = 1,       fifo_status_clk.clk
		.data_saved       (receive_packet_2_data_saved_data_saved)      //  output,   width = 1,            data_saved.data_saved
	);

	reset_main reset_main (
		.in_reset  (reset_mod_reset_main_reset), //   input,  width = 1,  in_reset.reset
		.out_reset (reset_main_out_reset)        //  output,  width = 1, out_reset.reset
	);

	reset_mod reset_mod (
		.clk       (reset_mod_clock_clk),        //   input,  width = 1,      clock.clk
		.rst_n     (reset_mod_reset_reset_n),    //   input,  width = 1,      reset.reset_n
		.reset     (reset_mod_reset_main_reset), //  output,  width = 1, reset_main.reset
		.reset_phy (reset_mod_reset_phy_reset)   //  output,  width = 1,  reset_phy.reset
	);

	send_cmd_pcie send_cmd_pcie (
		.clk                   (pcie_coreclkout_hip_clk),                                    //   input,   width = 1,              clock.clk
		.rst_n                 (pcie_app_nreset_status_reset),                               //   input,   width = 1,              reset.reset_n
		.avalon_mm_read        (mm_interconnect_6_send_cmd_pcie_avalon_slave_read),          //   input,   width = 1,       avalon_slave.read
		.avalon_mm_write       (mm_interconnect_6_send_cmd_pcie_avalon_slave_write),         //   input,   width = 1,                   .write
		.avalon_mm_addr        (mm_interconnect_6_send_cmd_pcie_avalon_slave_address),       //   input,  width = 16,                   .address
		.avalon_mm_write_data  (mm_interconnect_6_send_cmd_pcie_avalon_slave_writedata),     //   input,  width = 32,                   .writedata
		.avalon_mm_read_data   (mm_interconnect_6_send_cmd_pcie_avalon_slave_readdata),      //  output,  width = 32,                   .readdata
		.avalon_mm_rd_valid    (mm_interconnect_6_send_cmd_pcie_avalon_slave_readdatavalid), //  output,   width = 1,                   .readdatavalid
		.start_ram_addr        (pcie_send_control_start_ram_addr),                           //  output,   width = 6,       send_control.start_ram_addr
		.send_cmd              (pcie_send_control_signal),                                   //  output,   width = 1,                   .signal
		.ddr_local_cal_success (setup_ddr_ddr_status_out_local_cal_success),                 //   input,   width = 1,         ddr_status.local_cal_success
		.ddr_local_cal_fail    (setup_ddr_ddr_status_out_local_cal_fail),                    //   input,   width = 1,                   .local_cal_fail
		.ddr_setup_done        (setup_ddr_setup_setup_done),                                 //   input,   width = 1,     ddr_setup_done.setup_done
		.system_main_reset     (setup_ddr_resets_information_main_reset),                    //   input,   width = 1, resets_information.main_reset
		.ddr_avalon_rst        (setup_ddr_resets_information_ddr_avalon_reset),              //   input,   width = 1,                   .ddr_avalon_reset
		.board_reset           (setup_ddr_resets_information_board_reset),                   //   input,   width = 1,                   .board_reset
		.ddr_setup_cmd         (send_cmd_pcie_ddr_setup_cmd_ddr_setup_cmd)                   //  output,   width = 1,      ddr_setup_cmd.ddr_setup_cmd
	);

	send_packet_1 send_packet_1 (
		.clk_original    (tse_mac_tx_clock_connection_0_clk),                   //   input,   width = 1,                   clock.clk
		.rst             (rst_controller_003_reset_out_reset),                  //   input,   width = 1,                   reset.reset
		.ram_addr        (send_packet_1_avalon_master_address),                 //  output,  width = 10,           avalon_master.address
		.ram_chipselect  (send_packet_1_avalon_master_chipselect),              //  output,   width = 1,                        .chipselect
		.ram_write       (send_packet_1_avalon_master_write),                   //  output,   width = 1,                        .write
		.ram_readdata    (send_packet_1_avalon_master_readdata),                //   input,  width = 32,                        .readdata
		.ram_writedata   (send_packet_1_avalon_master_writedata),               //  output,  width = 32,                        .writedata
		.ram_byteenable  (send_packet_1_avalon_master_byteenable),              //  output,   width = 4,                        .byteenable
		.ram_waitrequest (send_packet_1_avalon_master_waitrequest),             //   input,   width = 1,                        .waitrequest
		.ff_tx_data      (send_packet_1_avalon_streaming_source_data),          //  output,   width = 8, avalon_streaming_source.data
		.ff_tx_eop       (send_packet_1_avalon_streaming_source_endofpacket),   //  output,   width = 1,                        .endofpacket
		.ff_tx_err       (send_packet_1_avalon_streaming_source_error),         //  output,   width = 1,                        .error
		.ff_tx_rdy       (send_packet_1_avalon_streaming_source_ready),         //   input,   width = 1,                        .ready
		.ff_tx_sop       (send_packet_1_avalon_streaming_source_startofpacket), //  output,   width = 1,                        .startofpacket
		.ff_tx_wren      (send_packet_1_avalon_streaming_source_valid),         //  output,   width = 1,                        .valid
		.start_ram_addr  (send_packet_1_control_start_ram_addr),                //   input,  width = 25,                 control.start_ram_addr
		.cmd_send        (send_packet_1_control_cmd_send)                       //   input,   width = 1,                        .cmd_send
	);

	send_packet_1 send_packet_2 (
		.clk_original    (tse_mac_tx_clock_connection_1_clk),                   //   input,   width = 1,                   clock.clk
		.rst             (rst_controller_001_reset_out_reset),                  //   input,   width = 1,                   reset.reset
		.ram_addr        (send_packet_2_avalon_master_address),                 //  output,  width = 10,           avalon_master.address
		.ram_chipselect  (send_packet_2_avalon_master_chipselect),              //  output,   width = 1,                        .chipselect
		.ram_write       (send_packet_2_avalon_master_write),                   //  output,   width = 1,                        .write
		.ram_readdata    (send_packet_2_avalon_master_readdata),                //   input,  width = 32,                        .readdata
		.ram_writedata   (send_packet_2_avalon_master_writedata),               //  output,  width = 32,                        .writedata
		.ram_byteenable  (send_packet_2_avalon_master_byteenable),              //  output,   width = 4,                        .byteenable
		.ram_waitrequest (send_packet_2_avalon_master_waitrequest),             //   input,   width = 1,                        .waitrequest
		.ff_tx_data      (send_packet_2_avalon_streaming_source_data),          //  output,   width = 8, avalon_streaming_source.data
		.ff_tx_eop       (send_packet_2_avalon_streaming_source_endofpacket),   //  output,   width = 1,                        .endofpacket
		.ff_tx_err       (send_packet_2_avalon_streaming_source_error),         //  output,   width = 1,                        .error
		.ff_tx_rdy       (send_packet_2_avalon_streaming_source_ready),         //   input,   width = 1,                        .ready
		.ff_tx_sop       (send_packet_2_avalon_streaming_source_startofpacket), //  output,   width = 1,                        .startofpacket
		.ff_tx_wren      (send_packet_2_avalon_streaming_source_valid),         //  output,   width = 1,                        .valid
		.start_ram_addr  (send_packet_2_control_start_ram_addr),                //   input,  width = 25,                 control.start_ram_addr
		.cmd_send        (send_packet_2_control_cmd_send)                       //   input,   width = 1,                        .cmd_send
	);

	setup_ddr setup_ddr (
		.amm_addr                 (setup_ddr_avalon_master_address),               //  output,   width = 25,      avalon_master.address
		.amm_readdata             (setup_ddr_avalon_master_readdata),              //   input,  width = 256,                   .readdata
		.amm_writedata            (setup_ddr_avalon_master_writedata),             //  output,  width = 256,                   .writedata
		.amm_read                 (setup_ddr_avalon_master_read),                  //  output,    width = 1,                   .read
		.amm_write                (setup_ddr_avalon_master_write),                 //  output,    width = 1,                   .write
		.amm_byteenable           (setup_ddr_avalon_master_byteenable),            //  output,   width = 32,                   .byteenable
		.amm_burstcount           (setup_ddr_avalon_master_burstcount),            //  output,    width = 7,                   .burstcount
		.amm_readdatavalid        (setup_ddr_avalon_master_readdatavalid),         //   input,    width = 1,                   .readdatavalid
		.amm_ready                (setup_ddr_avalon_master_waitrequest),           //   input,    width = 1,                   .waitrequest
		.setup_done               (setup_ddr_setup_setup_done),                    //  output,    width = 1,              setup.setup_done
		.local_cal_success_avalon (ddr3_status_local_cal_success),                 //   input,    width = 1,         ddr_status.local_cal_success
		.local_cal_fail_avalon    (ddr3_status_local_cal_fail),                    //   input,    width = 1,                   .local_cal_fail
		.ram_ready                (ddr_ready_ram_ready),                           //   input,    width = 1,          ddr_ready.ram_ready
		.clk                      (pll_outclk0_clk),                               //   input,    width = 1,    clock_125_tx_rx.clk
		.avalon_clk               (ddr3_emif_usr_clk_clk),                         //   input,    width = 1,       clock_avalon.clk
		.clk_50                   (pll_outclk1_clk),                               //   input,    width = 1,           clock_50.clk
		.rst_n                    (reset_board_reset),                             //   input,    width = 1,        reset_board.reset
		.avalon_reset             (rst_controller_005_reset_out_reset),            //   input,    width = 1,       reset_avalon.reset
		.reset                    (reset_mod_reset_main_reset),                    //   input,    width = 1,       reset_module.reset
		.reset_local_cal_success  (mem_cal_success_cal_success),                   //  output,    width = 1,        cal_success.cal_success
		.ddr_local_cal_success    (setup_ddr_ddr_status_out_local_cal_success),    //  output,    width = 1,     ddr_status_out.local_cal_success
		.ddr_local_cal_fail       (setup_ddr_ddr_status_out_local_cal_fail),       //  output,    width = 1,                   .local_cal_fail
		.system_main_reset        (setup_ddr_resets_information_main_reset),       //  output,    width = 1, resets_information.main_reset
		.ddr_avalon_rst           (setup_ddr_resets_information_ddr_avalon_reset), //  output,    width = 1,                   .ddr_avalon_reset
		.board_reset              (setup_ddr_resets_information_board_reset),      //  output,    width = 1,                   .board_reset
		.ddr_setup_cmd_pci        (send_cmd_pcie_ddr_setup_cmd_ddr_setup_cmd)      //   input,    width = 1,      ddr_setup_cmd.ddr_setup_cmd
	);

	tse tse (
		.clk                  (pll_outclk1_clk),                                     //   input,   width = 1,        control_port_clock_connection.clk
		.reset                (rst_controller_reset_out_reset),                      //   input,   width = 1,                     reset_connection.reset
		.reg_data_out         (init_mac_avalon_master_readdata),                     //  output,  width = 32,                         control_port.readdata
		.reg_rd               (init_mac_avalon_master_read),                         //   input,   width = 1,                                     .read
		.reg_data_in          (init_mac_avalon_master_writedata),                    //   input,  width = 32,                                     .writedata
		.reg_wr               (init_mac_avalon_master_write),                        //   input,   width = 1,                                     .write
		.reg_busy             (init_mac_avalon_master_waitrequest),                  //  output,   width = 1,                                     .waitrequest
		.reg_addr             (init_mac_avalon_master_address),                      //   input,  width = 10,                                     .address
		.rx_afull_clk         (pll_outclk0_clk),                                     //   input,   width = 1, receive_fifo_status_clock_connection.clk
		.rx_afull_data        (receive_packet_1_fifo_status_data),                   //   input,   width = 2,                  receive_fifo_status.data
		.rx_afull_valid       (receive_packet_1_fifo_status_valid),                  //   input,   width = 1,                                     .valid
		.rx_afull_channel     (receive_packet_1_fifo_status_channel),                //   input,   width = 2,                                     .channel
		.mac_rx_clk_0         (tse_mac_rx_clock_connection_0_clk),                   //  output,   width = 1,            mac_rx_clock_connection_0.clk
		.mac_tx_clk_0         (tse_mac_tx_clock_connection_0_clk),                   //  output,   width = 1,            mac_tx_clock_connection_0.clk
		.data_rx_data_0       (tse_receive_0_data),                                  //  output,   width = 8,                            receive_0.data
		.data_rx_eop_0        (tse_receive_0_endofpacket),                           //  output,   width = 1,                                     .endofpacket
		.data_rx_error_0      (tse_receive_0_error),                                 //  output,   width = 5,                                     .error
		.data_rx_ready_0      (tse_receive_0_ready),                                 //   input,   width = 1,                                     .ready
		.data_rx_sop_0        (tse_receive_0_startofpacket),                         //  output,   width = 1,                                     .startofpacket
		.data_rx_valid_0      (tse_receive_0_valid),                                 //  output,   width = 1,                                     .valid
		.data_tx_data_0       (send_packet_1_avalon_streaming_source_data),          //   input,   width = 8,                           transmit_0.data
		.data_tx_eop_0        (send_packet_1_avalon_streaming_source_endofpacket),   //   input,   width = 1,                                     .endofpacket
		.data_tx_error_0      (send_packet_1_avalon_streaming_source_error),         //   input,   width = 1,                                     .error
		.data_tx_ready_0      (send_packet_1_avalon_streaming_source_ready),         //  output,   width = 1,                                     .ready
		.data_tx_sop_0        (send_packet_1_avalon_streaming_source_startofpacket), //   input,   width = 1,                                     .startofpacket
		.data_tx_valid_0      (send_packet_1_avalon_streaming_source_valid),         //   input,   width = 1,                                     .valid
		.pkt_class_data_0     (),                                                    //  output,   width = 5,                receive_packet_type_0.data
		.pkt_class_valid_0    (),                                                    //  output,   width = 1,                                     .valid
		.magic_wakeup_0       (mac_misc_1_magic_wakeup),                             //  output,   width = 1,                mac_misc_connection_0.magic_wakeup
		.magic_sleep_n_0      (mac_misc_1_magic_sleep_n),                            //   input,   width = 1,                                     .magic_sleep_n
		.tx_crc_fwd_0         (mac_misc_1_tx_crc_fwd),                               //   input,   width = 1,                                     .tx_crc_fwd
		.mdc                  (mac_mdio_mdc),                                        //  output,   width = 1,                  mac_mdio_connection.mdc
		.mdio_in              (mac_mdio_mdio_in),                                    //   input,   width = 1,                                     .mdio_in
		.mdio_out             (mac_mdio_mdio_out),                                   //  output,   width = 1,                                     .mdio_out
		.mdio_oen             (mac_mdio_mdio_oen),                                   //  output,   width = 1,                                     .mdio_oen
		.mac_rx_clk_1         (tse_mac_rx_clock_connection_1_clk),                   //  output,   width = 1,            mac_rx_clock_connection_1.clk
		.mac_tx_clk_1         (tse_mac_tx_clock_connection_1_clk),                   //  output,   width = 1,            mac_tx_clock_connection_1.clk
		.data_rx_data_1       (tse_receive_1_data),                                  //  output,   width = 8,                            receive_1.data
		.data_rx_eop_1        (tse_receive_1_endofpacket),                           //  output,   width = 1,                                     .endofpacket
		.data_rx_error_1      (tse_receive_1_error),                                 //  output,   width = 5,                                     .error
		.data_rx_ready_1      (tse_receive_1_ready),                                 //   input,   width = 1,                                     .ready
		.data_rx_sop_1        (tse_receive_1_startofpacket),                         //  output,   width = 1,                                     .startofpacket
		.data_rx_valid_1      (tse_receive_1_valid),                                 //  output,   width = 1,                                     .valid
		.data_tx_data_1       (send_packet_2_avalon_streaming_source_data),          //   input,   width = 8,                           transmit_1.data
		.data_tx_eop_1        (send_packet_2_avalon_streaming_source_endofpacket),   //   input,   width = 1,                                     .endofpacket
		.data_tx_error_1      (send_packet_2_avalon_streaming_source_error),         //   input,   width = 1,                                     .error
		.data_tx_ready_1      (send_packet_2_avalon_streaming_source_ready),         //  output,   width = 1,                                     .ready
		.data_tx_sop_1        (send_packet_2_avalon_streaming_source_startofpacket), //   input,   width = 1,                                     .startofpacket
		.data_tx_valid_1      (send_packet_2_avalon_streaming_source_valid),         //   input,   width = 1,                                     .valid
		.pkt_class_data_1     (),                                                    //  output,   width = 5,                receive_packet_type_1.data
		.pkt_class_valid_1    (),                                                    //  output,   width = 1,                                     .valid
		.magic_wakeup_1       (mac_misc_2_magic_wakeup),                             //  output,   width = 1,                mac_misc_connection_1.magic_wakeup
		.magic_sleep_n_1      (mac_misc_2_magic_sleep_n),                            //   input,   width = 1,                                     .magic_sleep_n
		.tx_crc_fwd_1         (mac_misc_2_tx_crc_fwd),                               //   input,   width = 1,                                     .tx_crc_fwd
		.mac_rx_clk_2         (),                                                    //  output,   width = 1,            mac_rx_clock_connection_2.clk
		.mac_tx_clk_2         (),                                                    //  output,   width = 1,            mac_tx_clock_connection_2.clk
		.data_rx_data_2       (),                                                    //  output,   width = 8,                            receive_2.data
		.data_rx_eop_2        (),                                                    //  output,   width = 1,                                     .endofpacket
		.data_rx_error_2      (),                                                    //  output,   width = 5,                                     .error
		.data_rx_ready_2      (),                                                    //   input,   width = 1,                                     .ready
		.data_rx_sop_2        (),                                                    //  output,   width = 1,                                     .startofpacket
		.data_rx_valid_2      (),                                                    //  output,   width = 1,                                     .valid
		.data_tx_data_2       (),                                                    //   input,   width = 8,                           transmit_2.data
		.data_tx_eop_2        (),                                                    //   input,   width = 1,                                     .endofpacket
		.data_tx_error_2      (),                                                    //   input,   width = 1,                                     .error
		.data_tx_ready_2      (),                                                    //  output,   width = 1,                                     .ready
		.data_tx_sop_2        (),                                                    //   input,   width = 1,                                     .startofpacket
		.data_tx_valid_2      (),                                                    //   input,   width = 1,                                     .valid
		.pkt_class_data_2     (),                                                    //  output,   width = 5,                receive_packet_type_2.data
		.pkt_class_valid_2    (),                                                    //  output,   width = 1,                                     .valid
		.magic_wakeup_2       (),                                                    //  output,   width = 1,                mac_misc_connection_2.magic_wakeup
		.magic_sleep_n_2      (),                                                    //   input,   width = 1,                                     .magic_sleep_n
		.tx_crc_fwd_2         (),                                                    //   input,   width = 1,                                     .tx_crc_fwd
		.mac_rx_clk_3         (),                                                    //  output,   width = 1,            mac_rx_clock_connection_3.clk
		.mac_tx_clk_3         (),                                                    //  output,   width = 1,            mac_tx_clock_connection_3.clk
		.data_rx_data_3       (),                                                    //  output,   width = 8,                            receive_3.data
		.data_rx_eop_3        (),                                                    //  output,   width = 1,                                     .endofpacket
		.data_rx_error_3      (),                                                    //  output,   width = 5,                                     .error
		.data_rx_ready_3      (),                                                    //   input,   width = 1,                                     .ready
		.data_rx_sop_3        (),                                                    //  output,   width = 1,                                     .startofpacket
		.data_rx_valid_3      (),                                                    //  output,   width = 1,                                     .valid
		.data_tx_data_3       (),                                                    //   input,   width = 8,                           transmit_3.data
		.data_tx_eop_3        (),                                                    //   input,   width = 1,                                     .endofpacket
		.data_tx_error_3      (),                                                    //   input,   width = 1,                                     .error
		.data_tx_ready_3      (),                                                    //  output,   width = 1,                                     .ready
		.data_tx_sop_3        (),                                                    //   input,   width = 1,                                     .startofpacket
		.data_tx_valid_3      (),                                                    //   input,   width = 1,                                     .valid
		.pkt_class_data_3     (),                                                    //  output,   width = 5,                receive_packet_type_3.data
		.pkt_class_valid_3    (),                                                    //  output,   width = 1,                                     .valid
		.magic_wakeup_3       (),                                                    //  output,   width = 1,                mac_misc_connection_3.magic_wakeup
		.magic_sleep_n_3      (),                                                    //   input,   width = 1,                                     .magic_sleep_n
		.tx_crc_fwd_3         (),                                                    //   input,   width = 1,                                     .tx_crc_fwd
		.ref_clk              (tse_ref_clk),                                         //   input,   width = 1,         pcs_ref_clk_clock_connection.clk
		.led_crs_0            (status_led_connection_0_crs),                         //  output,   width = 1,              status_led_connection_0.crs
		.led_link_0           (status_led_connection_0_link),                        //  output,   width = 1,                                     .link
		.led_panel_link_0     (status_led_connection_0_panel_link),                  //  output,   width = 1,                                     .panel_link
		.led_col_0            (status_led_connection_0_col),                         //  output,   width = 1,                                     .col
		.led_an_0             (status_led_connection_0_an),                          //  output,   width = 1,                                     .an
		.led_char_err_0       (status_led_connection_0_char_err),                    //  output,   width = 1,                                     .char_err
		.led_disp_err_0       (status_led_connection_0_disp_err),                    //  output,   width = 1,                                     .disp_err
		.tx_analogreset_0     (tx_analogreset_0_tx_analogreset),                     //   input,   width = 1,                     tx_analogreset_0.tx_analogreset
		.tx_digitalreset_0    (tx_digitalreset_0_tx_digitalreset),                   //   input,   width = 1,                    tx_digitalreset_0.tx_digitalreset
		.rx_analogreset_0     (rx_analogreset_0_rx_analogreset),                     //   input,   width = 1,                     rx_analogreset_0.rx_analogreset
		.rx_digitalreset_0    (rx_digitalreset_0_rx_digitalreset),                   //   input,   width = 1,                    rx_digitalreset_0.rx_digitalreset
		.tx_cal_busy_0        (tx_cal_busy_0_tx_cal_busy),                           //  output,   width = 1,                        tx_cal_busy_0.tx_cal_busy
		.rx_cal_busy_0        (rx_cal_busy_0_rx_cal_busy),                           //  output,   width = 1,                        rx_cal_busy_0.rx_cal_busy
		.tx_serial_clk_0      (xcvr_pll_tx_serial_clk_clk),                          //   input,   width = 1,                      tx_serial_clk_0.clk
		.rx_cdr_refclk_0      (tse_rx_cdr_refclk_0_clk),                             //   input,   width = 1,                      rx_cdr_refclk_0.clk
		.rx_set_locktodata_0  (rx_set_locktodata_0_rx_set_locktodata),               //   input,   width = 1,                  rx_set_locktodata_0.rx_set_locktodata
		.rx_set_locktoref_0   (rx_set_locktoref_0_rx_set_locktoref),                 //   input,   width = 1,                   rx_set_locktoref_0.rx_set_locktoref
		.rx_is_lockedtoref_0  (rx_is_lockedtoref_0_rx_is_lockedtoref),               //  output,   width = 1,                  rx_is_lockedtoref_0.rx_is_lockedtoref
		.rx_is_lockedtodata_0 (rx_is_lockedtodata_0_rx_is_lockedtodata),             //  output,   width = 1,                 rx_is_lockedtodata_0.rx_is_lockedtodata
		.rxp_0                (sgmii_1_rxp),                                         //   input,   width = 1,                  serial_connection_0.rxp
		.txp_0                (sgmii_1_txp),                                         //  output,   width = 1,                                     .txp
		.rx_recovclkout_0     (serdes_control_connection_0_export),                  //  output,   width = 1,          serdes_control_connection_0.export
		.led_crs_1            (status_led_connection_1_crs),                         //  output,   width = 1,              status_led_connection_1.crs
		.led_link_1           (status_led_connection_1_link),                        //  output,   width = 1,                                     .link
		.led_panel_link_1     (status_led_connection_1_panel_link),                  //  output,   width = 1,                                     .panel_link
		.led_col_1            (status_led_connection_1_col),                         //  output,   width = 1,                                     .col
		.led_an_1             (status_led_connection_1_an),                          //  output,   width = 1,                                     .an
		.led_char_err_1       (status_led_connection_1_char_err),                    //  output,   width = 1,                                     .char_err
		.led_disp_err_1       (status_led_connection_1_disp_err),                    //  output,   width = 1,                                     .disp_err
		.tx_analogreset_1     (tx_analogreset_1_tx_analogreset),                     //   input,   width = 1,                     tx_analogreset_1.tx_analogreset
		.tx_digitalreset_1    (tx_digitalreset_1_tx_digitalreset),                   //   input,   width = 1,                    tx_digitalreset_1.tx_digitalreset
		.rx_analogreset_1     (rx_analogreset_1_rx_analogreset),                     //   input,   width = 1,                     rx_analogreset_1.rx_analogreset
		.rx_digitalreset_1    (rx_digitalreset_1_rx_digitalreset),                   //   input,   width = 1,                    rx_digitalreset_1.rx_digitalreset
		.tx_cal_busy_1        (tx_cal_busy_1_tx_cal_busy),                           //  output,   width = 1,                        tx_cal_busy_1.tx_cal_busy
		.rx_cal_busy_1        (rx_cal_busy_1_rx_cal_busy),                           //  output,   width = 1,                        rx_cal_busy_1.rx_cal_busy
		.tx_serial_clk_1      (xcvr_pll_tx_serial_clk_clk),                          //   input,   width = 1,                      tx_serial_clk_1.clk
		.rx_cdr_refclk_1      (tse_rx_cdr_refclk_1_clk),                             //   input,   width = 1,                      rx_cdr_refclk_1.clk
		.rx_set_locktodata_1  (rx_set_locktodata_1_rx_set_locktodata),               //   input,   width = 1,                  rx_set_locktodata_1.rx_set_locktodata
		.rx_set_locktoref_1   (rx_set_locktoref_1_rx_set_locktoref),                 //   input,   width = 1,                   rx_set_locktoref_1.rx_set_locktoref
		.rx_is_lockedtoref_1  (rx_is_lockedtoref_1_rx_is_lockedtoref),               //  output,   width = 1,                  rx_is_lockedtoref_1.rx_is_lockedtoref
		.rx_is_lockedtodata_1 (rx_is_lockedtodata_1_rx_is_lockedtodata),             //  output,   width = 1,                 rx_is_lockedtodata_1.rx_is_lockedtodata
		.rxp_1                (sgmii_2_rxp),                                         //   input,   width = 1,                  serial_connection_1.rxp
		.txp_1                (sgmii_2_txp),                                         //  output,   width = 1,                                     .txp
		.rx_recovclkout_1     (serdes_control_connection_1_export),                  //  output,   width = 1,          serdes_control_connection_1.export
		.led_crs_2            (),                                                    //  output,   width = 1,              status_led_connection_2.crs
		.led_link_2           (),                                                    //  output,   width = 1,                                     .link
		.led_panel_link_2     (),                                                    //  output,   width = 1,                                     .panel_link
		.led_col_2            (),                                                    //  output,   width = 1,                                     .col
		.led_an_2             (),                                                    //  output,   width = 1,                                     .an
		.led_char_err_2       (),                                                    //  output,   width = 1,                                     .char_err
		.led_disp_err_2       (),                                                    //  output,   width = 1,                                     .disp_err
		.tx_analogreset_2     (),                                                    //   input,   width = 1,                     tx_analogreset_2.tx_analogreset
		.tx_digitalreset_2    (),                                                    //   input,   width = 1,                    tx_digitalreset_2.tx_digitalreset
		.rx_analogreset_2     (),                                                    //   input,   width = 1,                     rx_analogreset_2.rx_analogreset
		.rx_digitalreset_2    (),                                                    //   input,   width = 1,                    rx_digitalreset_2.rx_digitalreset
		.tx_cal_busy_2        (),                                                    //  output,   width = 1,                        tx_cal_busy_2.tx_cal_busy
		.rx_cal_busy_2        (),                                                    //  output,   width = 1,                        rx_cal_busy_2.rx_cal_busy
		.tx_serial_clk_2      (tse_tx_serial_clk_2_clk),                             //   input,   width = 1,                      tx_serial_clk_2.clk
		.rx_cdr_refclk_2      (tse_rx_cdr_refclk_2_clk),                             //   input,   width = 1,                      rx_cdr_refclk_2.clk
		.rx_set_locktodata_2  (),                                                    //   input,   width = 1,                  rx_set_locktodata_2.rx_set_locktodata
		.rx_set_locktoref_2   (),                                                    //   input,   width = 1,                   rx_set_locktoref_2.rx_set_locktoref
		.rx_is_lockedtoref_2  (),                                                    //  output,   width = 1,                  rx_is_lockedtoref_2.rx_is_lockedtoref
		.rx_is_lockedtodata_2 (),                                                    //  output,   width = 1,                 rx_is_lockedtodata_2.rx_is_lockedtodata
		.rxp_2                (sgmii_3_rxp),                                         //   input,   width = 1,                  serial_connection_2.rxp
		.txp_2                (sgmii_3_txp),                                         //  output,   width = 1,                                     .txp
		.rx_recovclkout_2     (),                                                    //  output,   width = 1,          serdes_control_connection_2.export
		.led_crs_3            (),                                                    //  output,   width = 1,              status_led_connection_3.crs
		.led_link_3           (),                                                    //  output,   width = 1,                                     .link
		.led_panel_link_3     (),                                                    //  output,   width = 1,                                     .panel_link
		.led_col_3            (),                                                    //  output,   width = 1,                                     .col
		.led_an_3             (),                                                    //  output,   width = 1,                                     .an
		.led_char_err_3       (),                                                    //  output,   width = 1,                                     .char_err
		.led_disp_err_3       (),                                                    //  output,   width = 1,                                     .disp_err
		.tx_analogreset_3     (),                                                    //   input,   width = 1,                     tx_analogreset_3.tx_analogreset
		.tx_digitalreset_3    (),                                                    //   input,   width = 1,                    tx_digitalreset_3.tx_digitalreset
		.rx_analogreset_3     (),                                                    //   input,   width = 1,                     rx_analogreset_3.rx_analogreset
		.rx_digitalreset_3    (),                                                    //   input,   width = 1,                    rx_digitalreset_3.rx_digitalreset
		.tx_cal_busy_3        (),                                                    //  output,   width = 1,                        tx_cal_busy_3.tx_cal_busy
		.rx_cal_busy_3        (),                                                    //  output,   width = 1,                        rx_cal_busy_3.rx_cal_busy
		.tx_serial_clk_3      (tse_tx_serial_clk_3_clk),                             //   input,   width = 1,                      tx_serial_clk_3.clk
		.rx_cdr_refclk_3      (tse_rx_cdr_refclk_3_clk),                             //   input,   width = 1,                      rx_cdr_refclk_3.clk
		.rx_set_locktodata_3  (),                                                    //   input,   width = 1,                  rx_set_locktodata_3.rx_set_locktodata
		.rx_set_locktoref_3   (),                                                    //   input,   width = 1,                   rx_set_locktoref_3.rx_set_locktoref
		.rx_is_lockedtoref_3  (),                                                    //  output,   width = 1,                  rx_is_lockedtoref_3.rx_is_lockedtoref
		.rx_is_lockedtodata_3 (),                                                    //  output,   width = 1,                 rx_is_lockedtodata_3.rx_is_lockedtodata
		.rxp_3                (sgmii_4_rxp),                                         //   input,   width = 1,                  serial_connection_3.rxp
		.txp_3                (sgmii_4_txp),                                         //  output,   width = 1,                                     .txp
		.rx_recovclkout_3     ()                                                     //  output,   width = 1,          serdes_control_connection_3.export
	);

	xcvr_pll xcvr_pll (
		.pll_powerdown (xcvr_pll_powerdown_pll_powerdown), //   input,  width = 1, pll_powerdown.pll_powerdown
		.pll_refclk0   (xcvr_pll_refclk_clk),              //   input,  width = 1,   pll_refclk0.clk
		.tx_serial_clk (xcvr_pll_tx_serial_clk_clk),       //  output,  width = 1, tx_serial_clk.clk
		.pll_locked    (),                                 //  output,  width = 1,    pll_locked.pll_locked
		.pll_cal_busy  ()                                  //  output,  width = 1,  pll_cal_busy.pll_cal_busy
	);

	system_design_altera_mm_interconnect_1920_656hvpi mm_interconnect_1 (
		.setup_ddr_avalon_master_address                            (setup_ddr_avalon_master_address),                 //   input,   width = 25,                              setup_ddr_avalon_master.address
		.setup_ddr_avalon_master_waitrequest                        (setup_ddr_avalon_master_waitrequest),             //  output,    width = 1,                                                     .waitrequest
		.setup_ddr_avalon_master_burstcount                         (setup_ddr_avalon_master_burstcount),              //   input,    width = 7,                                                     .burstcount
		.setup_ddr_avalon_master_byteenable                         (setup_ddr_avalon_master_byteenable),              //   input,   width = 32,                                                     .byteenable
		.setup_ddr_avalon_master_read                               (setup_ddr_avalon_master_read),                    //   input,    width = 1,                                                     .read
		.setup_ddr_avalon_master_readdata                           (setup_ddr_avalon_master_readdata),                //  output,  width = 256,                                                     .readdata
		.setup_ddr_avalon_master_readdatavalid                      (setup_ddr_avalon_master_readdatavalid),           //  output,    width = 1,                                                     .readdatavalid
		.setup_ddr_avalon_master_write                              (setup_ddr_avalon_master_write),                   //   input,    width = 1,                                                     .write
		.setup_ddr_avalon_master_writedata                          (setup_ddr_avalon_master_writedata),               //   input,  width = 256,                                                     .writedata
		.pcie_rxm_bar2_address                                      (pcie_rxm_bar2_address),                           //   input,   width = 64,                                        pcie_rxm_bar2.address
		.pcie_rxm_bar2_waitrequest                                  (pcie_rxm_bar2_waitrequest),                       //  output,    width = 1,                                                     .waitrequest
		.pcie_rxm_bar2_burstcount                                   (pcie_rxm_bar2_burstcount),                        //   input,    width = 6,                                                     .burstcount
		.pcie_rxm_bar2_byteenable                                   (pcie_rxm_bar2_byteenable),                        //   input,   width = 16,                                                     .byteenable
		.pcie_rxm_bar2_read                                         (pcie_rxm_bar2_read),                              //   input,    width = 1,                                                     .read
		.pcie_rxm_bar2_readdata                                     (pcie_rxm_bar2_readdata),                          //  output,  width = 128,                                                     .readdata
		.pcie_rxm_bar2_readdatavalid                                (pcie_rxm_bar2_readdatavalid),                     //  output,    width = 1,                                                     .readdatavalid
		.pcie_rxm_bar2_write                                        (pcie_rxm_bar2_write),                             //   input,    width = 1,                                                     .write
		.pcie_rxm_bar2_writedata                                    (pcie_rxm_bar2_writedata),                         //   input,  width = 128,                                                     .writedata
		.ddr3_ctrl_amm_0_address                                    (mm_interconnect_1_ddr3_ctrl_amm_0_address),       //  output,   width = 25,                                      ddr3_ctrl_amm_0.address
		.ddr3_ctrl_amm_0_write                                      (mm_interconnect_1_ddr3_ctrl_amm_0_write),         //  output,    width = 1,                                                     .write
		.ddr3_ctrl_amm_0_read                                       (mm_interconnect_1_ddr3_ctrl_amm_0_read),          //  output,    width = 1,                                                     .read
		.ddr3_ctrl_amm_0_readdata                                   (mm_interconnect_1_ddr3_ctrl_amm_0_readdata),      //   input,  width = 256,                                                     .readdata
		.ddr3_ctrl_amm_0_writedata                                  (mm_interconnect_1_ddr3_ctrl_amm_0_writedata),     //  output,  width = 256,                                                     .writedata
		.ddr3_ctrl_amm_0_burstcount                                 (mm_interconnect_1_ddr3_ctrl_amm_0_burstcount),    //  output,    width = 7,                                                     .burstcount
		.ddr3_ctrl_amm_0_byteenable                                 (mm_interconnect_1_ddr3_ctrl_amm_0_byteenable),    //  output,   width = 32,                                                     .byteenable
		.ddr3_ctrl_amm_0_readdatavalid                              (mm_interconnect_1_ddr3_ctrl_amm_0_readdatavalid), //   input,    width = 1,                                                     .readdatavalid
		.ddr3_ctrl_amm_0_waitrequest                                (~mm_interconnect_1_ddr3_ctrl_amm_0_waitrequest),  //   input,    width = 1,                                                     .waitrequest
		.setup_ddr_reset_avalon_reset_bridge_in_reset_reset         (rst_controller_005_reset_out_reset),              //   input,    width = 1,         setup_ddr_reset_avalon_reset_bridge_in_reset.reset
		.pcie_rxm_bar2_translator_reset_reset_bridge_in_reset_reset (~pcie_app_nreset_status_reset),                   //   input,    width = 1, pcie_rxm_bar2_translator_reset_reset_bridge_in_reset.reset
		.ddr3_emif_usr_clk_clk                                      (ddr3_emif_usr_clk_clk),                           //   input,    width = 1,                                    ddr3_emif_usr_clk.clk
		.pcie_coreclkout_hip_clk                                    (pcie_coreclkout_hip_clk)                          //   input,    width = 1,                                  pcie_coreclkout_hip.clk
	);

	system_design_altera_mm_interconnect_1920_qky3gdi mm_interconnect_2 (
		.receive_packet_1_avalon_master_address             (receive_packet_1_avalon_master_address),     //   input,  width = 10,               receive_packet_1_avalon_master.address
		.receive_packet_1_avalon_master_waitrequest         (receive_packet_1_avalon_master_waitrequest), //  output,   width = 1,                                             .waitrequest
		.receive_packet_1_avalon_master_byteenable          (receive_packet_1_avalon_master_byteenable),  //   input,   width = 4,                                             .byteenable
		.receive_packet_1_avalon_master_chipselect          (receive_packet_1_avalon_master_chipselect),  //   input,   width = 1,                                             .chipselect
		.receive_packet_1_avalon_master_readdata            (receive_packet_1_avalon_master_readdata),    //  output,  width = 32,                                             .readdata
		.receive_packet_1_avalon_master_write               (receive_packet_1_avalon_master_write),       //   input,   width = 1,                                             .write
		.receive_packet_1_avalon_master_writedata           (receive_packet_1_avalon_master_writedata),   //   input,  width = 32,                                             .writedata
		.mem_rcv_1_s1_address                               (mm_interconnect_2_mem_rcv_1_s1_address),     //  output,  width = 10,                                 mem_rcv_1_s1.address
		.mem_rcv_1_s1_write                                 (mm_interconnect_2_mem_rcv_1_s1_write),       //  output,   width = 1,                                             .write
		.mem_rcv_1_s1_readdata                              (mm_interconnect_2_mem_rcv_1_s1_readdata),    //   input,  width = 32,                                             .readdata
		.mem_rcv_1_s1_writedata                             (mm_interconnect_2_mem_rcv_1_s1_writedata),   //  output,  width = 32,                                             .writedata
		.mem_rcv_1_s1_byteenable                            (mm_interconnect_2_mem_rcv_1_s1_byteenable),  //  output,   width = 4,                                             .byteenable
		.mem_rcv_1_s1_chipselect                            (mm_interconnect_2_mem_rcv_1_s1_chipselect),  //  output,   width = 1,                                             .chipselect
		.mem_rcv_1_s1_clken                                 (mm_interconnect_2_mem_rcv_1_s1_clken),       //  output,   width = 1,                                             .clken
		.receive_packet_1_reset_reset_bridge_in_reset_reset (rst_controller_004_reset_out_reset),         //   input,   width = 1, receive_packet_1_reset_reset_bridge_in_reset.reset
		.tse_mac_rx_clock_connection_0_clk                  (tse_mac_rx_clock_connection_0_clk)           //   input,   width = 1,                tse_mac_rx_clock_connection_0.clk
	);

	system_design_altera_mm_interconnect_1920_tqdmh6a mm_interconnect_3 (
		.send_packet_2_avalon_master_address             (send_packet_2_avalon_master_address),     //   input,  width = 10,               send_packet_2_avalon_master.address
		.send_packet_2_avalon_master_waitrequest         (send_packet_2_avalon_master_waitrequest), //  output,   width = 1,                                          .waitrequest
		.send_packet_2_avalon_master_byteenable          (send_packet_2_avalon_master_byteenable),  //   input,   width = 4,                                          .byteenable
		.send_packet_2_avalon_master_chipselect          (send_packet_2_avalon_master_chipselect),  //   input,   width = 1,                                          .chipselect
		.send_packet_2_avalon_master_readdata            (send_packet_2_avalon_master_readdata),    //  output,  width = 32,                                          .readdata
		.send_packet_2_avalon_master_write               (send_packet_2_avalon_master_write),       //   input,   width = 1,                                          .write
		.send_packet_2_avalon_master_writedata           (send_packet_2_avalon_master_writedata),   //   input,  width = 32,                                          .writedata
		.mem_4_s1_address                                (mm_interconnect_3_mem_4_s1_address),      //  output,  width = 10,                                  mem_4_s1.address
		.mem_4_s1_write                                  (mm_interconnect_3_mem_4_s1_write),        //  output,   width = 1,                                          .write
		.mem_4_s1_readdata                               (mm_interconnect_3_mem_4_s1_readdata),     //   input,  width = 32,                                          .readdata
		.mem_4_s1_writedata                              (mm_interconnect_3_mem_4_s1_writedata),    //  output,  width = 32,                                          .writedata
		.mem_4_s1_byteenable                             (mm_interconnect_3_mem_4_s1_byteenable),   //  output,   width = 4,                                          .byteenable
		.mem_4_s1_chipselect                             (mm_interconnect_3_mem_4_s1_chipselect),   //  output,   width = 1,                                          .chipselect
		.mem_4_s1_clken                                  (mm_interconnect_3_mem_4_s1_clken),        //  output,   width = 1,                                          .clken
		.send_packet_2_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),      //   input,   width = 1, send_packet_2_reset_reset_bridge_in_reset.reset
		.tse_mac_tx_clock_connection_1_clk               (tse_mac_tx_clock_connection_1_clk)        //   input,   width = 1,             tse_mac_tx_clock_connection_1.clk
	);

	system_design_altera_mm_interconnect_1920_nnzxfdi mm_interconnect_4 (
		.send_packet_1_avalon_master_address             (send_packet_1_avalon_master_address),     //   input,  width = 10,               send_packet_1_avalon_master.address
		.send_packet_1_avalon_master_waitrequest         (send_packet_1_avalon_master_waitrequest), //  output,   width = 1,                                          .waitrequest
		.send_packet_1_avalon_master_byteenable          (send_packet_1_avalon_master_byteenable),  //   input,   width = 4,                                          .byteenable
		.send_packet_1_avalon_master_chipselect          (send_packet_1_avalon_master_chipselect),  //   input,   width = 1,                                          .chipselect
		.send_packet_1_avalon_master_readdata            (send_packet_1_avalon_master_readdata),    //  output,  width = 32,                                          .readdata
		.send_packet_1_avalon_master_write               (send_packet_1_avalon_master_write),       //   input,   width = 1,                                          .write
		.send_packet_1_avalon_master_writedata           (send_packet_1_avalon_master_writedata),   //   input,  width = 32,                                          .writedata
		.mem_5_s1_address                                (mm_interconnect_4_mem_5_s1_address),      //  output,  width = 10,                                  mem_5_s1.address
		.mem_5_s1_write                                  (mm_interconnect_4_mem_5_s1_write),        //  output,   width = 1,                                          .write
		.mem_5_s1_readdata                               (mm_interconnect_4_mem_5_s1_readdata),     //   input,  width = 32,                                          .readdata
		.mem_5_s1_writedata                              (mm_interconnect_4_mem_5_s1_writedata),    //  output,  width = 32,                                          .writedata
		.mem_5_s1_byteenable                             (mm_interconnect_4_mem_5_s1_byteenable),   //  output,   width = 4,                                          .byteenable
		.mem_5_s1_chipselect                             (mm_interconnect_4_mem_5_s1_chipselect),   //  output,   width = 1,                                          .chipselect
		.mem_5_s1_clken                                  (mm_interconnect_4_mem_5_s1_clken),        //  output,   width = 1,                                          .clken
		.send_packet_1_reset_reset_bridge_in_reset_reset (rst_controller_003_reset_out_reset),      //   input,   width = 1, send_packet_1_reset_reset_bridge_in_reset.reset
		.tse_mac_tx_clock_connection_0_clk               (tse_mac_tx_clock_connection_0_clk)        //   input,   width = 1,             tse_mac_tx_clock_connection_0.clk
	);

	system_design_altera_mm_interconnect_1920_rvh6iyy mm_interconnect_5 (
		.receive_packet_2_avalon_master_address             (receive_packet_2_avalon_master_address),     //   input,  width = 10,               receive_packet_2_avalon_master.address
		.receive_packet_2_avalon_master_waitrequest         (receive_packet_2_avalon_master_waitrequest), //  output,   width = 1,                                             .waitrequest
		.receive_packet_2_avalon_master_byteenable          (receive_packet_2_avalon_master_byteenable),  //   input,   width = 4,                                             .byteenable
		.receive_packet_2_avalon_master_chipselect          (receive_packet_2_avalon_master_chipselect),  //   input,   width = 1,                                             .chipselect
		.receive_packet_2_avalon_master_readdata            (receive_packet_2_avalon_master_readdata),    //  output,  width = 32,                                             .readdata
		.receive_packet_2_avalon_master_write               (receive_packet_2_avalon_master_write),       //   input,   width = 1,                                             .write
		.receive_packet_2_avalon_master_writedata           (receive_packet_2_avalon_master_writedata),   //   input,  width = 32,                                             .writedata
		.mem_4_s2_address                                   (mm_interconnect_5_mem_4_s2_address),         //  output,  width = 10,                                     mem_4_s2.address
		.mem_4_s2_write                                     (mm_interconnect_5_mem_4_s2_write),           //  output,   width = 1,                                             .write
		.mem_4_s2_readdata                                  (mm_interconnect_5_mem_4_s2_readdata),        //   input,  width = 32,                                             .readdata
		.mem_4_s2_writedata                                 (mm_interconnect_5_mem_4_s2_writedata),       //  output,  width = 32,                                             .writedata
		.mem_4_s2_byteenable                                (mm_interconnect_5_mem_4_s2_byteenable),      //  output,   width = 4,                                             .byteenable
		.mem_4_s2_chipselect                                (mm_interconnect_5_mem_4_s2_chipselect),      //  output,   width = 1,                                             .chipselect
		.mem_4_s2_clken                                     (mm_interconnect_5_mem_4_s2_clken),           //  output,   width = 1,                                             .clken
		.receive_packet_2_reset_reset_bridge_in_reset_reset (rst_controller_002_reset_out_reset),         //   input,   width = 1, receive_packet_2_reset_reset_bridge_in_reset.reset
		.tse_mac_rx_clock_connection_1_clk                  (tse_mac_rx_clock_connection_1_clk)           //   input,   width = 1,                tse_mac_rx_clock_connection_1.clk
	);

	system_design_altera_mm_interconnect_1920_nmewghq mm_interconnect_6 (
		.pcie_rxm_bar0_address                                      (pcie_rxm_bar0_address),                                      //   input,   width = 64,                                        pcie_rxm_bar0.address
		.pcie_rxm_bar0_waitrequest                                  (pcie_rxm_bar0_waitrequest),                                  //  output,    width = 1,                                                     .waitrequest
		.pcie_rxm_bar0_burstcount                                   (pcie_rxm_bar0_burstcount),                                   //   input,    width = 6,                                                     .burstcount
		.pcie_rxm_bar0_byteenable                                   (pcie_rxm_bar0_byteenable),                                   //   input,   width = 16,                                                     .byteenable
		.pcie_rxm_bar0_read                                         (pcie_rxm_bar0_read),                                         //   input,    width = 1,                                                     .read
		.pcie_rxm_bar0_readdata                                     (pcie_rxm_bar0_readdata),                                     //  output,  width = 128,                                                     .readdata
		.pcie_rxm_bar0_readdatavalid                                (pcie_rxm_bar0_readdatavalid),                                //  output,    width = 1,                                                     .readdatavalid
		.pcie_rxm_bar0_write                                        (pcie_rxm_bar0_write),                                        //   input,    width = 1,                                                     .write
		.pcie_rxm_bar0_writedata                                    (pcie_rxm_bar0_writedata),                                    //   input,  width = 128,                                                     .writedata
		.send_cmd_pcie_avalon_slave_address                         (mm_interconnect_6_send_cmd_pcie_avalon_slave_address),       //  output,   width = 16,                           send_cmd_pcie_avalon_slave.address
		.send_cmd_pcie_avalon_slave_write                           (mm_interconnect_6_send_cmd_pcie_avalon_slave_write),         //  output,    width = 1,                                                     .write
		.send_cmd_pcie_avalon_slave_read                            (mm_interconnect_6_send_cmd_pcie_avalon_slave_read),          //  output,    width = 1,                                                     .read
		.send_cmd_pcie_avalon_slave_readdata                        (mm_interconnect_6_send_cmd_pcie_avalon_slave_readdata),      //   input,   width = 32,                                                     .readdata
		.send_cmd_pcie_avalon_slave_writedata                       (mm_interconnect_6_send_cmd_pcie_avalon_slave_writedata),     //  output,   width = 32,                                                     .writedata
		.send_cmd_pcie_avalon_slave_readdatavalid                   (mm_interconnect_6_send_cmd_pcie_avalon_slave_readdatavalid), //   input,    width = 1,                                                     .readdatavalid
		.pcie_rxm_bar0_translator_reset_reset_bridge_in_reset_reset (~pcie_app_nreset_status_reset),                              //   input,    width = 1, pcie_rxm_bar0_translator_reset_reset_bridge_in_reset.reset
		.pcie_coreclkout_hip_clk                                    (pcie_coreclkout_hip_clk)                                     //   input,    width = 1,                                  pcie_coreclkout_hip.clk
	);

	system_design_altera_irq_mapper_1920_66fzifq irq_mapper (
		.clk        (pcie_coreclkout_hip_clk),       //   input,   width = 1,       clk.clk
		.reset      (~pcie_app_nreset_status_reset), //   input,   width = 1, clk_reset.reset
		.sender_irq (pcie_rxm_irq_irq)               //  output,  width = 16,    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (reset_mod_reset_main_reset),     //   input,  width = 1, reset_in0.reset
		.clk            (pll_outclk1_clk),                //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                               // (terminated),                       
		.reset_req_in0  (1'b0),                           // (terminated),                       
		.reset_in1      (1'b0),                           // (terminated),                       
		.reset_req_in1  (1'b0),                           // (terminated),                       
		.reset_in2      (1'b0),                           // (terminated),                       
		.reset_req_in2  (1'b0),                           // (terminated),                       
		.reset_in3      (1'b0),                           // (terminated),                       
		.reset_req_in3  (1'b0),                           // (terminated),                       
		.reset_in4      (1'b0),                           // (terminated),                       
		.reset_req_in4  (1'b0),                           // (terminated),                       
		.reset_in5      (1'b0),                           // (terminated),                       
		.reset_req_in5  (1'b0),                           // (terminated),                       
		.reset_in6      (1'b0),                           // (terminated),                       
		.reset_req_in6  (1'b0),                           // (terminated),                       
		.reset_in7      (1'b0),                           // (terminated),                       
		.reset_req_in7  (1'b0),                           // (terminated),                       
		.reset_in8      (1'b0),                           // (terminated),                       
		.reset_req_in8  (1'b0),                           // (terminated),                       
		.reset_in9      (1'b0),                           // (terminated),                       
		.reset_req_in9  (1'b0),                           // (terminated),                       
		.reset_in10     (1'b0),                           // (terminated),                       
		.reset_req_in10 (1'b0),                           // (terminated),                       
		.reset_in11     (1'b0),                           // (terminated),                       
		.reset_req_in11 (1'b0),                           // (terminated),                       
		.reset_in12     (1'b0),                           // (terminated),                       
		.reset_req_in12 (1'b0),                           // (terminated),                       
		.reset_in13     (1'b0),                           // (terminated),                       
		.reset_req_in13 (1'b0),                           // (terminated),                       
		.reset_in14     (1'b0),                           // (terminated),                       
		.reset_req_in14 (1'b0),                           // (terminated),                       
		.reset_in15     (1'b0),                           // (terminated),                       
		.reset_req_in15 (1'b0)                            // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (reset_mod_reset_main_reset),             //   input,  width = 1, reset_in0.reset
		.clk            (tse_mac_tx_clock_connection_1_clk),      //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     //  output,  width = 1, reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //  output,  width = 1,          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated),                       
		.reset_in1      (1'b0),                                   // (terminated),                       
		.reset_req_in1  (1'b0),                                   // (terminated),                       
		.reset_in2      (1'b0),                                   // (terminated),                       
		.reset_req_in2  (1'b0),                                   // (terminated),                       
		.reset_in3      (1'b0),                                   // (terminated),                       
		.reset_req_in3  (1'b0),                                   // (terminated),                       
		.reset_in4      (1'b0),                                   // (terminated),                       
		.reset_req_in4  (1'b0),                                   // (terminated),                       
		.reset_in5      (1'b0),                                   // (terminated),                       
		.reset_req_in5  (1'b0),                                   // (terminated),                       
		.reset_in6      (1'b0),                                   // (terminated),                       
		.reset_req_in6  (1'b0),                                   // (terminated),                       
		.reset_in7      (1'b0),                                   // (terminated),                       
		.reset_req_in7  (1'b0),                                   // (terminated),                       
		.reset_in8      (1'b0),                                   // (terminated),                       
		.reset_req_in8  (1'b0),                                   // (terminated),                       
		.reset_in9      (1'b0),                                   // (terminated),                       
		.reset_req_in9  (1'b0),                                   // (terminated),                       
		.reset_in10     (1'b0),                                   // (terminated),                       
		.reset_req_in10 (1'b0),                                   // (terminated),                       
		.reset_in11     (1'b0),                                   // (terminated),                       
		.reset_req_in11 (1'b0),                                   // (terminated),                       
		.reset_in12     (1'b0),                                   // (terminated),                       
		.reset_req_in12 (1'b0),                                   // (terminated),                       
		.reset_in13     (1'b0),                                   // (terminated),                       
		.reset_req_in13 (1'b0),                                   // (terminated),                       
		.reset_in14     (1'b0),                                   // (terminated),                       
		.reset_req_in14 (1'b0),                                   // (terminated),                       
		.reset_in15     (1'b0),                                   // (terminated),                       
		.reset_req_in15 (1'b0)                                    // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (reset_mod_reset_main_reset),             //   input,  width = 1, reset_in0.reset
		.clk            (tse_mac_rx_clock_connection_1_clk),      //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     //  output,  width = 1, reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //  output,  width = 1,          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated),                       
		.reset_in1      (1'b0),                                   // (terminated),                       
		.reset_req_in1  (1'b0),                                   // (terminated),                       
		.reset_in2      (1'b0),                                   // (terminated),                       
		.reset_req_in2  (1'b0),                                   // (terminated),                       
		.reset_in3      (1'b0),                                   // (terminated),                       
		.reset_req_in3  (1'b0),                                   // (terminated),                       
		.reset_in4      (1'b0),                                   // (terminated),                       
		.reset_req_in4  (1'b0),                                   // (terminated),                       
		.reset_in5      (1'b0),                                   // (terminated),                       
		.reset_req_in5  (1'b0),                                   // (terminated),                       
		.reset_in6      (1'b0),                                   // (terminated),                       
		.reset_req_in6  (1'b0),                                   // (terminated),                       
		.reset_in7      (1'b0),                                   // (terminated),                       
		.reset_req_in7  (1'b0),                                   // (terminated),                       
		.reset_in8      (1'b0),                                   // (terminated),                       
		.reset_req_in8  (1'b0),                                   // (terminated),                       
		.reset_in9      (1'b0),                                   // (terminated),                       
		.reset_req_in9  (1'b0),                                   // (terminated),                       
		.reset_in10     (1'b0),                                   // (terminated),                       
		.reset_req_in10 (1'b0),                                   // (terminated),                       
		.reset_in11     (1'b0),                                   // (terminated),                       
		.reset_req_in11 (1'b0),                                   // (terminated),                       
		.reset_in12     (1'b0),                                   // (terminated),                       
		.reset_req_in12 (1'b0),                                   // (terminated),                       
		.reset_in13     (1'b0),                                   // (terminated),                       
		.reset_req_in13 (1'b0),                                   // (terminated),                       
		.reset_in14     (1'b0),                                   // (terminated),                       
		.reset_req_in14 (1'b0),                                   // (terminated),                       
		.reset_in15     (1'b0),                                   // (terminated),                       
		.reset_req_in15 (1'b0)                                    // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (reset_mod_reset_main_reset),             //   input,  width = 1, reset_in0.reset
		.clk            (tse_mac_tx_clock_connection_0_clk),      //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset),     //  output,  width = 1, reset_out.reset
		.reset_req      (rst_controller_003_reset_out_reset_req), //  output,  width = 1,          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated),                       
		.reset_in1      (1'b0),                                   // (terminated),                       
		.reset_req_in1  (1'b0),                                   // (terminated),                       
		.reset_in2      (1'b0),                                   // (terminated),                       
		.reset_req_in2  (1'b0),                                   // (terminated),                       
		.reset_in3      (1'b0),                                   // (terminated),                       
		.reset_req_in3  (1'b0),                                   // (terminated),                       
		.reset_in4      (1'b0),                                   // (terminated),                       
		.reset_req_in4  (1'b0),                                   // (terminated),                       
		.reset_in5      (1'b0),                                   // (terminated),                       
		.reset_req_in5  (1'b0),                                   // (terminated),                       
		.reset_in6      (1'b0),                                   // (terminated),                       
		.reset_req_in6  (1'b0),                                   // (terminated),                       
		.reset_in7      (1'b0),                                   // (terminated),                       
		.reset_req_in7  (1'b0),                                   // (terminated),                       
		.reset_in8      (1'b0),                                   // (terminated),                       
		.reset_req_in8  (1'b0),                                   // (terminated),                       
		.reset_in9      (1'b0),                                   // (terminated),                       
		.reset_req_in9  (1'b0),                                   // (terminated),                       
		.reset_in10     (1'b0),                                   // (terminated),                       
		.reset_req_in10 (1'b0),                                   // (terminated),                       
		.reset_in11     (1'b0),                                   // (terminated),                       
		.reset_req_in11 (1'b0),                                   // (terminated),                       
		.reset_in12     (1'b0),                                   // (terminated),                       
		.reset_req_in12 (1'b0),                                   // (terminated),                       
		.reset_in13     (1'b0),                                   // (terminated),                       
		.reset_req_in13 (1'b0),                                   // (terminated),                       
		.reset_in14     (1'b0),                                   // (terminated),                       
		.reset_req_in14 (1'b0),                                   // (terminated),                       
		.reset_in15     (1'b0),                                   // (terminated),                       
		.reset_req_in15 (1'b0)                                    // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (reset_mod_reset_main_reset),             //   input,  width = 1, reset_in0.reset
		.clk            (tse_mac_rx_clock_connection_0_clk),      //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset),     //  output,  width = 1, reset_out.reset
		.reset_req      (rst_controller_004_reset_out_reset_req), //  output,  width = 1,          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated),                       
		.reset_in1      (1'b0),                                   // (terminated),                       
		.reset_req_in1  (1'b0),                                   // (terminated),                       
		.reset_in2      (1'b0),                                   // (terminated),                       
		.reset_req_in2  (1'b0),                                   // (terminated),                       
		.reset_in3      (1'b0),                                   // (terminated),                       
		.reset_req_in3  (1'b0),                                   // (terminated),                       
		.reset_in4      (1'b0),                                   // (terminated),                       
		.reset_req_in4  (1'b0),                                   // (terminated),                       
		.reset_in5      (1'b0),                                   // (terminated),                       
		.reset_req_in5  (1'b0),                                   // (terminated),                       
		.reset_in6      (1'b0),                                   // (terminated),                       
		.reset_req_in6  (1'b0),                                   // (terminated),                       
		.reset_in7      (1'b0),                                   // (terminated),                       
		.reset_req_in7  (1'b0),                                   // (terminated),                       
		.reset_in8      (1'b0),                                   // (terminated),                       
		.reset_req_in8  (1'b0),                                   // (terminated),                       
		.reset_in9      (1'b0),                                   // (terminated),                       
		.reset_req_in9  (1'b0),                                   // (terminated),                       
		.reset_in10     (1'b0),                                   // (terminated),                       
		.reset_req_in10 (1'b0),                                   // (terminated),                       
		.reset_in11     (1'b0),                                   // (terminated),                       
		.reset_req_in11 (1'b0),                                   // (terminated),                       
		.reset_in12     (1'b0),                                   // (terminated),                       
		.reset_req_in12 (1'b0),                                   // (terminated),                       
		.reset_in13     (1'b0),                                   // (terminated),                       
		.reset_req_in13 (1'b0),                                   // (terminated),                       
		.reset_in14     (1'b0),                                   // (terminated),                       
		.reset_req_in14 (1'b0),                                   // (terminated),                       
		.reset_in15     (1'b0),                                   // (terminated),                       
		.reset_req_in15 (1'b0)                                    // (terminated),                       
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~ddr3_emif_usr_reset_n_reset),       //   input,  width = 1, reset_in0.reset
		.clk            (ddr3_emif_usr_clk_clk),              //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                                   // (terminated),                       
		.reset_req_in0  (1'b0),                               // (terminated),                       
		.reset_in1      (1'b0),                               // (terminated),                       
		.reset_req_in1  (1'b0),                               // (terminated),                       
		.reset_in2      (1'b0),                               // (terminated),                       
		.reset_req_in2  (1'b0),                               // (terminated),                       
		.reset_in3      (1'b0),                               // (terminated),                       
		.reset_req_in3  (1'b0),                               // (terminated),                       
		.reset_in4      (1'b0),                               // (terminated),                       
		.reset_req_in4  (1'b0),                               // (terminated),                       
		.reset_in5      (1'b0),                               // (terminated),                       
		.reset_req_in5  (1'b0),                               // (terminated),                       
		.reset_in6      (1'b0),                               // (terminated),                       
		.reset_req_in6  (1'b0),                               // (terminated),                       
		.reset_in7      (1'b0),                               // (terminated),                       
		.reset_req_in7  (1'b0),                               // (terminated),                       
		.reset_in8      (1'b0),                               // (terminated),                       
		.reset_req_in8  (1'b0),                               // (terminated),                       
		.reset_in9      (1'b0),                               // (terminated),                       
		.reset_req_in9  (1'b0),                               // (terminated),                       
		.reset_in10     (1'b0),                               // (terminated),                       
		.reset_req_in10 (1'b0),                               // (terminated),                       
		.reset_in11     (1'b0),                               // (terminated),                       
		.reset_req_in11 (1'b0),                               // (terminated),                       
		.reset_in12     (1'b0),                               // (terminated),                       
		.reset_req_in12 (1'b0),                               // (terminated),                       
		.reset_in13     (1'b0),                               // (terminated),                       
		.reset_req_in13 (1'b0),                               // (terminated),                       
		.reset_in14     (1'b0),                               // (terminated),                       
		.reset_req_in14 (1'b0),                               // (terminated),                       
		.reset_in15     (1'b0),                               // (terminated),                       
		.reset_req_in15 (1'b0)                                // (terminated),                       
	);

endmodule
