`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
DN/BfmzWEdhtzhBEn06RkZwL8EFNc2oOEF18SeM7/bjo7YZktpqGnkpA7GR3a/J0
17ySSfOKak2ehEQNOH07yQnLwv6wqotaKqUca++EjKuyAkeVhYh7PHc8xQOp6nnr
Jb1QtgXAldDlGg3iNR2x2aXRmOS445f1bjU1mkKjFmQ=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 70496), data_block
L3Sf15N2MB6XMCLK5/Ltywy1boC5ES52P2cHp7gM5UCQF/DxPiNf/Li+0qqnwRJ1
yr5E3FqVkns+77nBQ7LEBK1rMbzXjak8H8txErIPs8Rz60vSumqSV+PPingmhl3g
iZzkxq9FZLX+JMIiPirVo/7DMVAWutYQo76kGjNDpgvYJzL3jjqdmys/yxAkmkUZ
n9L6h47lsb43YqaKWHoEnyaMq3k4WIBNBKMQn39opNB81uf2EOAfTyYBaEjA08l3
3dDa7XRe9u/l/OgHfejlrfi5R+tbyzSCrI/klDDim4Lfyd4jLudfkjWhXLOqU84d
AYK5eU4UEd8NYgKvFMTy6rWzXjNrQjeWoeA/w+remwS1eJucVFDtil9l6+ZAJ43g
B8jThvTwX/x8HJe9In4eMxR96NvU53PdkkdzBxcKJdmVSPjQovh5pWyQpnmDq5RH
SJP89OvGX4AMppvPhvxOXnmtWSlVUn6XH3qtdC7mq2NkSx0lL9r1JDLo1rOMJR3/
tSZVOs/CSHuDFS1qKYHgZzyV//D7LaLqNqxv1n/o7iZxZU3sfcucu4F56SuqT0WM
ft4cdujUmO5rlUDqvkhf3oHpOTJXH1sknBDkOkeuR/XAXc9AtPRq3BIyIPtteNgG
AQ4elp32oT4rHvddhavkIKv8DkhKYHoRwdr3DTYOqtwRpBt//EnPhIsGwCNTwaWG
E7SxE7Ym/kpGLBgIDaXQGG917pO91UL1NgQ+fzK6DeOa4pZX/+/PrAhLC7NAqIDO
nO2S9J3nIyU0FK7ToQXfp+TTQgsTb5R5jIl1CkBfE1f9jjSdrgof/Lku9zldfw1b
u08ZtLsKU9FkbPvmICDujA6wGca3HEpsklj5jvzBrBJ6+kJ6s5TKicozWC9w80Jt
eJrL2e9nhgt47xmWcVMSZdJEauioCZSY0BY1ITdyT0yjp4ZNgfvFJkezxGgPpe+f
zt9O+RcFZPnzZJOFMl70ZBoN71ZrlE3D35iatcw2ERzaKNVlkZudcZ3wpZk9dFvp
/imKhJLr9b4ityfOCsbBwaSMzDaK+AndPzTDgC+enZuYmdVBn5nda2Hk7Z56m9ZV
SzhRySV5wWlqXwcyqbVuRRPqssogIVrMCpHNHc0M5uP+34iLdP/Q1UExd8nRXJuX
RlwX51ooxZdgDqBR8KUAMRSNFakh8sK5lt+vMZhPZdCqN7C9HdomLHJeEe4fQQoj
ncrWA2TwHGDKY5ctCDAj1XzIyV1g0hpggxxaAjzzzd/Tkjgoq+zUikzCFv84IVUB
u0EXs4h3nxodCv/rsc2VxJjdpwPEV5Ws9y7WlHfdDZL+gvqM7x/XCXPw5eW3XDND
3/I1c4TKvHDEV7a8/bVpD1QUL5QIHo3ALyoq2LfxY56Oo9bx1TlngZKM4hMNPSsq
TLKnvmgNjvCcD2c5L7vZZW5P1BgH99TlRYhSkHh+e9g0Bi9lUFIgbGQXCRWjE5NH
ajhqdWDdE8zNzfNA3PoPV/6mE8sxD6AGqgOJKYq1VmZUvUh3WbuZFNh7nxrk7TU+
kocznPybDZAe3sOz7nn/3M5mUp679/xwozxJBQ74Ou6KTy4KkvrwTbR61YQ2MX1d
sidcdRU8ASiJW0w9ISwzQ2HdX0e3/G4SZjL6XMpVvmIFUZLa7eP1LjsCtBL0e+vg
OC5k5NWBEKsgSXcW3WZSUjG+0x7oMYMxxEcKr+VdzuS0eaZLwLgawn5fw73ZuLeJ
luaCpE+j2FxqOG3H7qYxsAMslOqgXVx2/lo6XYIM84R1kQ1XPVxglmUIX9Et9kOp
P6AbdTKLpaRSlrVNJztHdSdqsns1gOSzsLYdV2e8er/dppf/8CtL9BvogYkJsovc
l91y4Z56R3mCv5KPFFCI5RXt6WdjE8a0PuNB5CHS+iAWkLlA4FFQpfk9j1UoghBa
EurFXyntDeraahM4ae2gnxAQycjM98xv8ITqyOQifyCsHBaHVgPrhAht2VESsHbW
a3PX6DxxMXfpjL+rNxss0e6STToU+qWerwkCIZ9w2VWu3tx/VJtRXUs9MGEw5V4Z
JOcMVVtzrljI6Egf7HuD2nHJ/6Q0jPj8aPqb03cn3i+fQb60grxY+azF8avpGF9t
iVHAbnYMDnr5i8aBSHnS0i5FQp11LPCifP+oWHw6rSxtCI5Vj8HDKlo3Uo7DPMVK
MReUDeKVO8tNHf3G8huGi595qZveGNCw57PiAjQAEZVtfrmhprg1aS6yJmLPptoJ
LLN3XEPTIfMvXw44XLouiWyT2URlVuVo+aXaYb8xrE2tJ/WCxNiiwD9pDUVE29tQ
M1+h+faq06TeQzrR9RcIZQ4Z0JdsCTBD6B9bg0vLA5bbRGpKCfAKw1g/aVo/acsL
DdriRfoh+iU/n8lhFBMVS/B+tdND5pniWFOa954Ie+dbdRcXM3Gp7XHZZSUYo1CB
ncDtLGm6BNcHRa/0KGKnNYqeAASuOdqQ6Umds0P1AH22oufzXxo17t+tdiOQk86w
IQElTLxiKno8MN7FZVtC2/Lfh5RCykWztqAXxYQPf4HBshLIbK1wbf7E0tColth8
FPUkAFjHkPLEN0SdIrMGNwbITvHAL0N190f/T3C7bLWhx2jd1uqnJDVQMQIhGHqO
s1eojHLjMcXjXKFiYWadGsqW/cm/BDzetIa94DfuFDh//ay+ikb03pTrEdtXgFd+
HLdIqb16Kvx1RsOepZcLPCGp7cPCwzfhA/UnuQn6gwQs4Ftv1MoTGUNLE0gmda11
EPEeF3+ncj6bGenRKaZ9QVjg9nn2FfNvr3KrpbO+WZ3EUsxYzulICRgMMePHrCzg
mgOSFrJ4ebqyRczj5v55oQHhFcpLO5ynlnfVdmV56KK1jJq/5bnOJ1dVtXJPwVpf
6ahSDLGG+xCyFJwn8vevCfZrWO0x2bKK9bX3AS7I2eWW0ZioHL6kl87Oj+yftLQr
kfx8X0NrX4t9zGtIIsodAArxakrggkfjHZoTezzdu5XeymGUvAndCmzFcJWWwmqs
9UgTTHLSTllotGeNH05TSp1YCIZhacZ/soa5LgxLpVsQwmQKGCWMJK1VTa/Mtjsv
UtMcmMX8+Rf09B8HzcMnKEzUsNH0A5cR1po+uN5bVsYWqTJjW5MD+3ea6mqq3p4a
qh/NcNYvwBkYOvDDWxwHyoB81CGNGENFTvRuiaRexMquLTMMyn3cmD2k4pC1Nyqi
tv4HNNLS/J/JG1+mU4JuNc2sxsSW7nUqBDLtwFnXOn33q6GycKVH9tyxIayecxJ8
5Kjg88JILsB1b20bQO8V4liSDn/LeujmzkjUQfX72CXOiUGuXixcTMi+qUbc3jIf
uu+mIpEXiMdSVfOncUy6ejwV1KXhWWzO5X+XMV3TEqSVMYH/lpelRs0/G6bqqz1L
ALMSL7FjJD15Am8M8losR/FYOiudrTDXVSf9lLQjJNk6OSHIlpNGCJQL2SQK/NUi
mvhQHsXpyPD3N1OxRRSZIvKW5FUzjgv38Opnyij5anXVNMZni2i/YZ+wO0FmxXfO
rlOu2XDCFB0DnsLMisQHiUptIDySgUCF0YZ+srd6W+m5jeVEcwT6sC4Ff4Ltu828
JGOwfCh6l7IQwWwdw7aX12ZAjMb6OTWUM7uAS0iTk1jySPGsPwD6LEDOHjDtGtaW
4rHwF4AOLmMizszK/GRYBB/aHE34Jf5sJQ0rIzFqEMRF862TwrNUY2PcEoat4DWr
R61yU0tmgZjX01jICX3ciMUMtwA7f1N+8d3pXjbqqOTOC6UV4d7R+T0BhQOL6zOI
Zp+ZPLbkDbHCgfLZcLZHBcjDmxzObNhwwOFF9N01yCbI4QFhz1k/jsDO9VcUzdfq
azlm4F1MiZ4AWEH15xk1sdOrhos6ylG8cCEHYcRS8J3vN80Len18BPd/IQsTxMAe
QxD3HSh2u8yiNSxnB0aP9MFC002VG6bPoD+iYJAlzwMw/XiKkU/CONvqMMSv6QdU
Wu/O4qUB3H+vI0zwd1MuWhJV0SPMPkgVchMudf5KnINvyyBd6XH316N56knp6r4B
pyDs6wUWWRaWaNrixZRvMptK/2Vhoz5aosgsVN25o9qum2A1WDW9L3PY1kelZu5z
HkwsxD3hJMtuGV4dW8Hkdp+gBxYhcbnoxQQyTZuT+l+4oqPbsFZsPsT/If2KG7ZX
aA6umA9cd7LGQl7DOP9eZqj16fG1l3DDzae6nW3sf97TzGNQS6NMdH0RHmJHkWia
8berIZMndooGIJJLXcN2P0oIgk0GR0esOVqWQ3vVPe7pqSIzQZgDQe/ehmxxQ5Ei
bIpbxJZfE1vS9TIdWg5YtV7XU7bnU8uLh5N+TcZmDVeUgNWs/72lnBAvexSqFNTx
4UwLhokc5t/niGUXwByfCZJI81YgJDgwQY0Q2+c3/b1TlHkIP8i8Vb9YMr13O/QK
oaeINJNPRjBBo03KXkdm+tmk1AcLwRTGnVXLaDlMcWZsVEiNkgoKjQeXuaMceorM
nEW3RWhXd/SSPGGK9JfSK5ZgAvKFb6cgYUyHDE2xGXCsaRgxqRcqsKf6tRSYMZcJ
3QCWUXumjuaOWa5WDrgM25B8P5B6JvekAJXRrRNVWTp9nTv4SPususDV7745AyVN
qz/vNlLDAouOl4roiheXJ+E72IlgOXjEt+zYwROF07bZhk+weu0I0s1/ChaaL5Px
fYHpVRsGpDAi77Xife02ydPfEbk6U1MVBC4mr+TOFLY6mzsaPo5I8yAhUndOJ4FB
e7hEu0UM/BqSfDZVw0cEih+sgs1lU9XdG/iGm8zoIe1c8d6XqiXCo5n8Ea3LvDot
EA2+eWvOEVZXAAakftpyU0qKo3EkqcobpqJqwLXtFEVboxhq2p/aNd7AIaqF0o33
iwDSwILNyB9d0Wsco9TmiACfKQsM9FrRO9OiYHuvmhEK89MOjn1WdI3wsiTQV/1K
N2ETEW89jhL2MrWsRl+ZPVa1N1N0EOUj4r5wsX2GKUYX5Om+LMTREombBjbKHqpD
Ee3Q/CLZ8cFAwvblxVsFt5YqnKTDTEW/Lmj1m5Zld7QLgQAlhQgGw3T3rFzxI2zq
18R4Gh+I0K5xA3XEewQDOCFdHR3JJIkSymJa25eydPvMHQe+PEkNnXLIAk7TpP4K
xgCAlfFrbe4JzeBoWvPz3NUce4HWN+mzDkTZ61znBt9WapGBoiMCv8EP3TmZNjng
Fx032ztMtYkfLGk5G1ezz8aPi7To55KaVYFfoM3a66TyOu3ml+YaTBkF3UJGstN4
ilNPxJLHqvdzgNosWXSf3Q9itgQy7c3YV4+7lMpx4lxF4tNZLfEOvhleTbh4HYFm
RBFfZBXvtN88qsRmbeOWmHEFp0TKFUdZyOzDCpIzjOdoNxJ7v3viqXW0c53GIVjh
VHBV+1jeq4pO0woLQoMprRpgo51QA1PyjH93cpjUeI8mLcTBOdR0+FIwFcEwnHk+
LUojzRDsujjhsptgxvYM0gc3qSE0XquXiY2I5zm0iSHlVIpqOgXsNnWrnnDMFL2s
zdmkFN8LJQ6j8dcDkDv4B34m25Q25SV5u76c8H98POz/Q/ET/RE4AOyHhr9N5sAm
IfxtZnHhs63gOHNmhSBXWBjsJfJIoeQhNwjUS6BADM5bqiXvr8nip/nQ3nTp1UqJ
C1lFPQ2xQeTFwQMR+LOTcQn4if+S2tpjjZGq9aLVDxFxFw/rrX6oDGu6JrZbXFG8
m2F+fPYs1G2P1Yc6Zlst8z8zjDfweVFlnmQDozDDrTkCpI2LYIj3nmKQY4En6Rs2
4kcxPFo3a1S7vthsLlXevGciNXvX7FRA3efj4BX+AXTyZid1/kVUdd2Tz3422JHR
4y21aq4+QmVUHw9MMsTIY0locDXXOI108VsdPmPRsHHiuW3m6joIz0OiNzep5qNM
zK34TVQ/Am5t+bTWOhZwO4A9UzboQ7Lke1fSOie55QIDECB7dSSjhZfxUZ+kk61k
KgJf20WDtn8dvWmOiZ2fmH2V4xByqspbQEd9/J0a7e6T74zWHDO8rjNe0Ub1xVan
HsTUFfivwKpjM/C8TvpZoK5kA466x6UwiHeJq15zZNGTLdA6ub+1zejK3sLRI984
kBddK9bQbxndipm59ofiF2CZn/P/+pLhu2fd33Z3D3CO5bJXdgNOju5OUuChSACP
ygENBjdHDzElGzlk6aBXEm6R355KlsWePaWjQQGOe9oiBU0ntzfyT7zICH4FRWQY
t49v9Hf2FH0gak55nYDUaNGyXjakveyRtENdvAA/+kU2GpZixWmCii3fGOSpzr+y
QSXTonMJMJOYuXRJ8Angqxd7X4qag0lIzDXi1nBZd5RqYYQq42iQcjfgV8DyrWx/
lTEX637p9ev9lzB+zs938a6+dib2nFzzQ1EHT4tVWGXIYauBd9p/hRvM4vuoX5S5
CIi/twthcZ5gh5LqHDTQeJmlWHpVP7On0X1i2WXQF47mGeowLB4J5W5USeo8b3Zs
PQ+/yLs7XUx0ygQSgHJfkNjKVfgtU71qRrjyTVy3AmkSUyXXvWsT1t4Wtm7J4PzE
r/FlQudTHhc3f4qzjGI4a9g1wZGt4ARECzg6xlgULRjWZx+UxHDDI1UgllrC3HqM
D0qXTB6feJWQg5HGjo7uefmJ3SajVgsbOO+u21BA1a16jphD3NPVfbz/3+4ycbxa
GH4frK3OyT9y+kqUhAPGW7sYYEdnV1oNk2O6ITY31C7Wu327CcX1ePAcrxjrpRg3
OceeBg4wOAiG7w8A/ELrOb0DqXWbxmpeZZ1L3LVkvAyNcs4xQMoOprLFO4CK8eA6
alctmm8WNCthRSlZrWcReZktNEmSs9tNy08xddBzL6VDiNYnPZPZyg6EY/mdZZXj
W1DsOsFtUk5nB+fzLuz/3FMjk0vlgS2gt/mlChWCsQ5kYS9eCvx4FwBJExiXARAp
P/iisg34qFZVFjRgSKygHMvbzpTKWOTKW8LgepD+dbCmlnFIbZ6rBEZehSl+G9Q3
3bdjE3DwjyqXKwYykNmyciFhfu9StbDeDLdFuucUk5f7h3VyqEdqvK2+sx6HiTK3
OBCDwg3AIgqkBNOZScP3dG/5uaifRgaDlXF405zFjDAQzyrxSGt77ymlFlE0wVN3
vMXnbnzFsFFtYto6NcftjNT/BmcXXEKIDRJLnr47RP6+JPL2gQh8Z7D8EaK3w++1
4FqPTGkdoLIpm8iEG26+1C3nmm/gdfbI+tl+QthPoJELwILIfkCMdwlaJzq6eJrV
PbuMeDlepjV0OcN8yblSKJoPXpZgWIVoKCNpxLToZmycc3OSgVYXdBQlr5/Qajf7
VBaqRWnURwrwe4fPb9idn26JoX2ccAx5puWWgaGWvdtY8lJpx/ls1yRYO6i84oPK
sh7j2KUdd/jh635VFqXpfcTyzCgbNfaDVhfQzixtu64Kx7MUQyX3NgYu/yW37Ta7
BTmfmYI1KpdESxquWv03cg0XXXApKeL7OkRFMaim60KwQnDNuV2bU0BXgK3JMqmZ
OA4prGB90rduBf6lG4M8Gzt246VO1dSuEOjRppa+iA9ftK5GzPQPyrW1Lkmzg8Xq
h7oaLVQKKCshxiBGsamwBkuTv4OkQlyS9uVhW+1M4l4Uf1M0yfWJD8QlwGk2q6Q1
+PWA9hhNKum4AZDbqBmI3RDuutnoRz9XTPobpYt151poI9VXQwguxJAreutVr1w9
VmHfYVpmckPQARPqSAY+cDTBqKB12266XMqvREjvqWMqKj/83mz87lDITWixstRk
IoGQc7hm+ErRPUfPCgn0i91OVA/ade+VhhXhTQw2z7KAHRorKmB1l/2D+rjTKN+l
L5MzRIaYcX3hDZ5izG2FJ8g7gfDBNhlm6DnaRr7xdpv8IBFpiWfYtVkSSSE8FKHQ
8A/xmnunkHSkPsxXG5O2d3xcGfvSWub+e6h+8E7rFsYuJguAUgW79l3oAqHsS0dI
Vu9KNlsFHmQ3tEpsXEmhz3GN6OaAdJoeOWSCt4Cq/ogKtzgNXLLdQMld08W7K6Kh
Ou7cFfc9p/D2fCsBTJY/PiYTGEjEqHFY8EkSHKExzUOv6SCm1qfJ0B1ul0gvWlbk
lBIqxN/lENdad/Z5J/RVwvC0xecsW6ETCVoHzUm57yu63MRvceP6zHWocfQEPcIH
8KCr5P5EZl2FMeerf6m5GecTB0yk70AooJihpH4jOzmepOTJy/zCjDJ0t3zJPXNq
nQWuncJMnQWFm71S3J7T/10ov/TAHXkO66qjBBK6U3tcbyY1pHC41WSjJGoQa7Yw
Kqz0iWwTY8ywq22BIZnOCJdKb/cwFhmw7OwjbvCon3Kf2UUEqG/qVs7iwfi2OxtY
spmjOFIk5CCYhUAGruJZ4r3i9j99ylIA68ZkHFNoVvJyGnFkt9a9ZGMdj5/agQpZ
qv+RFHPM1AET7KmwVxRZY3YL2rqGFu6Wx18DLTYQN3LzmIGzl9TUsXO5iQHecWkE
HwZ3JQzwD5Q8tqvV0ZSNk+saawTZzrrUQjTN6q0pVeW/VEPCvwuBvwBE5yOSR5S7
7yr5WOfzp55K2aap96DKvuvTNkxS7vbbejXgQaQnY9rRNveXn5ytZIJEmG7fFvFk
mDiEt9HFBNDHnuODY1NQmuWu/Pc9eITHcfFoWAZHYhNXyNbbFfHXTQN0VK8niUXJ
cQuukoP9x/q28QLleJCIJjrpE+JzF2e0ETQFlYzOcHUmQ00QL1YCNOizGudlp45P
+L1orw3EX7rs0eGXTLV3ekFOawwVXrQ9b+ucJyRbFe4BHL0wqjhfiZWRIoC18zii
malKWoPOJQJCJWQX+0Uc72nli1e94CZi2BCQh/np5CYpwk6Lo8p2wjpQQ/0+gQKx
ZQeMKKMOFg7zIa4dm0tA3s21ZHo8OxtfzTB19DRyWbSA7zRX2Af9ZfeLnL3yGQCr
ThlaM+/GKVLdm5jnwgyuZQlZYXVaJatPWK2ws98xZAs/Gy9Zg8d8QPMSrVy3HoeE
9Q2pzv/xMGwmO2u/upl9pdAJ274U0j9Nx2RGvJU3sIFlX9RNnVEETWu8qkDIIL2a
TXsB8sb5nvKMNCcvW+uy4SayEBt+0NEWYpy6x+ZJC1c5QgPOq+Uilqtb+JaFzMl8
TqAkSKe5UfSPtrSvH/9q/5yb27Mi3cimKLmgSsv0N1QrkigTQP6FBpGbpwmyc1n6
TqhMq7UYldi1OAxD+JTg4+wdROk/mdRA2R6bQ24cjjxi5fINx2s3IkSAUHyteYfQ
e9W6Bgbvo+DRTHuNLYyL41b78WntnwfR01eqbFiFPbXvYdzhB6JrgbqUGTTjUbhj
t2sMBRfTKAdJo5PuYe6r2F04/I+cLKdAmVYTptocs5+96yCZmBr1BMT/7SwV/Vh0
pZ2r0atyzMce5jRl9uCfyacp2xpTXAkfl3TizElXrdLIfUjW2dEXfUbrceAZjf6C
o7BApbcZBcEWMCeEXELq5+gz82Q/2j2GgL7VlEL5Dfp8T0SqL1Bx5kbS6EJDT2W9
s+mAu3Mrl/wceWU5lD/jwYKY0w/EUJ5hZVZjwceGKOX9/oVGoAM54OUPLuU7oKpo
tSqKBxSmlvyWpp6LS0OdIrsSRiKqqDXn6lQNfN8kbaxXl6R7URGqBgyR50rpYMzy
YZ3COpXqVAVg3ZUA3YgNdfadBtnlL91HNifvKXBczQsReZ5YtzoaYFEWPp/kHWqe
YYHmumJs1LZE3Y4EMOtgVxqQq2Qz+1ro57oxHTXyeUgBbbU+/Wgi++b+pf6qE2q1
KKnTM2QDEgbzJHPBr4utN1XxDn8gwDQdQC4uC0XQKpY6BIKWVUoPYIFko86Py+ha
CRNK+HQWEdHqywEVPDUwk/KRmuqCIsqnOkZIs6SeQ5qTYLQpxqJdydpIEiUV2d87
DXCnQM4kvH/syQDgwKLD5VG2rBoBFGOceNVj/7KiHvo7WfC+KU64ivGt40h+aUAi
otUM8D9Sdc4u3tUbnvXiVbRc3Bb2WOJT30D9rUzcnFQ3faHmD1xnXo0Rrg4rOtVx
OmbqDG2X+Ustm2PAgC0A9/srG4jZE6LhTqbN5B5T/D2LN+uok3856MEI58BQYkCC
qSxlHaeAr2AttwkeEk0iC1XRhsb2lnPxGFRizb8Ja+c4iMB7kYdTS00Vh/caMHvA
fE1hRMHqHUv0rq4M3Uuvsfk/vHVg+N9Coni9mCaPj1nD1Ud4iug5Tg4BCnCekhsL
ziicS0aQg9FCbNqet0UDkBvr8mQtz99rGcfoRquDWcP7xaEuHJTDgLUGcwcy+XSS
hhz9LF1x4L4IqBl+F62gYsKSqB6B8MmnpBQwsahGBHeTAZJ1NjqwQPJMolwNEyxe
QT4Ecr/LlFXvaMtvKyDEfuqaScQyycvPCWtKSgmw4CmWgJsxl3VfAnoHFVYAKqRo
HGQ7AvqpYYerTWGKcB7taiSs1OvOlAlhOYmSQppOd0xOtl1EZRvecp7+8R+aBcyJ
mb70tOe9I+9Ram2bh5XE9uXQH7evzr4ItuKoduLv+ZBl6rkRJn48ppLoKVOMolFT
dTMdsZfEitJGSyA5CXXSHcuKg4W9mYvHB6UKJJ88qXzzScL5c+y21fQAVl3osA1A
3V+7E4si00TIxSvZhQHBFODdjS4YUBi+OcCbtMBF9a4/FGorBJq+UhE/FYPgQHWi
sP1ifYYtPBhHcs2+eDyuFcm3Z6p5g0wuv7e2RXpWWC1a6h/oVPGnuP2MFFVTK8CW
ktZ6b9y+l76xrXRl6jUu2phEfqXcj+d8izMGWajoxOmQ3KJI494sh2r0yH6nLHGr
VueaOkrygcYYgKlYDMpKk9eVHbg7zphbaf8J0XLwUtrdyJg6L/nQV1YQy3Sv0vbW
zLcmjjoAe+ZoLMI1um0a14Kfm0rtrTZwlXT8WCotPxAxxHM2/ReFSVo2J/92/JsN
pSwuZWdjnHjc5JF3WiaVt+9q7/zI2qwpAuCiSpJG0+AlTMpXFB/bfhCj6WDmqU1A
/oMD5/JqSot2IIMZBK4SWuwMncPgi198ksu7rrbNnYZdSv0XvpmFWRyYvD5TdZUk
0GnrWPW4oD7Jg57UPqlYNUXbN1HZ4ViezmjOfX0LYB3L/V9zApclpirTLK7BLvML
wT/6u7F8zcUhHRQBjL0ObDiJSXcZLB8RfhIdih/I3jtNIURQbiFbzyGQ9kdQhBbX
Zch4kJ/D8G5pz272As0GDoiH+8PbspodJmARTp5tl/yhjxeouLtti1U7gj0WEmPs
Pc9yO0hwD93Pp9NGmbFzfQ11uX8+d9pC52GG47/ZuK4BjL9+dUArA/HQEJtuWld0
0MxIlzoNQr8AZ9tGtsiFFRx89EgRUApveSEA7fKzRvf0MAG3In7ZF+fcR2Gn5K7a
vC0ZFAjeFVoWOcDJQTJPk+oUqaLWotz6G+G9Ks052PWLzxC0ue4gv20RB99TOiZ8
EYB1OSEqgKL++rlVxf4sF1C9TQ7Bi6nCllwKHTI9KY+qj6lJUpADyI1Ai5sweoSn
T791WwpMXu64K6KOK9XAD7UCu/W4KQ6T8JDgkDQBPmWVouYFfURUUpcDCJ+k06Xh
uwIkc72X6ybWsJXS5bW2DvCebriOmB7Od6jaxxikthAm7HEf9Vv4y+hnvGmN8Elc
5tU4H8pzX2ngw6eF+lV1vqsgZCXdWU0vYUmPIV1CKeXETUYh44yaXiqaFOBSM+Vk
UcW5Ye3zoOmgpAecVC4meyz/kQM4jQXM474DhL3gUqtlUdORgMmS9SUtRNO3zhxa
SyqfHSUuYQertKx0GSzFiXx6htabwAi/Ki5ygQMdGYhrLZOodhDE2ksdheQemFKW
0ggzCdzQkAGwt2pKVCtlG7dtZoa16uYf0dV4wohQ7uJSyuCc2HwSRipGts9sKJj3
9KRoJH3U2jkStL04K/JbBf+/+SFgZ5zAvxMlWypC3nIeDBL9u0N95K/QJgmFdqcs
XHss1XIbzsWej/y+wpkTQdFA6wHVdCHQK/wzA3XIr+76BCmm5oDqI+FN0XriVWpI
/uplZ1yRfBKlbyFA8gsy7ojAcamCYPJX+2j7lHufUJvKMBVMiIET3/U+szRQuATL
VdW/NtQ1N9YHW/3/WWcKrkWwrbFe+Qz+/nQe1JFf/i7ul2J4Iavw6+8CTKeg7v7E
b1omcbI/89AsqTyG7Ihl2gatiYkQabvMRIB8EmYDzmffw28I7w5ALa9bLrPFGvy2
OFLkZOA56UaWTa2pFoZmRmUlTpubgtTeoSkqYwELikaU28OKTHh0SYnnLGH4Z8d0
7d1krU5GWREI0lPaYWlkGpBNbYfjFTt4SVR/vQNCxYPY2jxJyeLPiRxxtgoi0Xdo
5Bmn3CWfee7fMJtnVikzBON6xixH5gDs2t539qxPZPw+BuEpUBzimZqdOdkzcGyx
M6x2Cl3XHAHxZUXoIOh4m2wiqadYCw5v1RQRcc825f7yH5JkD9h9FP4phiwXjTOV
cHy8gsDZvYvNY4q/5TLY/WTqdF4V4tSF1ZWH+R2LbvBasj7ZxJo6LT+em5pWQqxr
Ir6JHcuDQdR4QCYnzkDAjP5mHZbJ7x3WP4xhiQNtf+xvMpcAv71SEz0e+MC6hv7V
MBp6McC1dGKC8wZSOHMsKQTbJU1r21qNHH5OJe+CnazZbi3BnrrswtxrkQ8Q9A5A
MvpAh0FBgPqB1KQPULNn6blNvzdH8OF5ZKPCfJ5yIHiXaoN4ODiyJ+vehuX+yNql
6ItQWg2+7+h3qApy/usCwy38C/BAZkWF3hm7XqgcXI8eraT/W3zxbNNKPXbzr0F0
ylYWmjJya4E/QfVOJgZVGYC2GtnD2KxsJ8T8Y9iHu1DqPq5uvz1HySmAeFfCOMBz
wBjOPD2yAwg7L6t6gwtGh7oUtj3K+aR+0lJSP4wbJeo0eKsoPjOm+y5sGeelr4UW
0Btf8dvLT/7alOiWDLsZ4MD0X9wa5XArHNJf22ge4lzJWTkPJjGd54MCOuH6lVO0
C9oybUO9dWJIL5SzvssgRuop7XFP/HBCRJ3aR3Rb6zkM4eEQ96XOLEt0GRhibg/V
Dw4cOGBUbMNPweh5BvCc2kBvkCLY1KtR/3EgTHe/wb0/g+uxbLKieE9QCNkBKWEg
sYHxN5GLKDxcwbWvvdaTBYJIWpvFOwPJOUEjlcqav1SAtIysT9oTZtFSpkiN93f1
4vjxhrZFI1c00OnCPl5Kj8PwqC8UJgwkElMgyj3mpNPti53cMUlVg+t+0+afqN5r
FvmEWr8cQ7DTWPahbh3g8z+P4Jqc7Rz++KzluxSy28z3o1n4f58WED+fL36A2b1v
NxQMUWmtoWU0BQvt4jvYQTz4UGBcMpbKSh94Wro2kqiEcjhANcAikG/deYr7FOQd
c/Y9OuR/Hut52Jq9E9n4jT0NzuiGX4c6uy862aocwuhV4nuD2Oh0ZpCdRKF9D3oT
ZcKopZ0I0HzfafCy9HFN5SKQMGlI97WigrUhWW79I4SkEDzElZhiBzsFKt8K3lLk
c6tEqbFhugA6qA4/St4VJzBfHOYWpN8Ve3zzm00amKNoRdW3I/LXnHik8kkJtnRF
Ec7rAPn9GgApMc4+HYsPLjtLpSgS6qH/39ZZvDFkyzpfF1VuT/nXnlFH3NgCe0Zx
xa+HeiqAjLol01tgcDQWHS5YTMhKT3V6rDz+lrTNujc+pL6hbynO4APa4aR62bD5
PBLFiPY02PS+R4+3J7BWWOemezAkgq2c1eY051Khmyn8enV0Ci5NRjiFf/3sPwZl
AzlSRm9ZHY6VYdqAbl+fxXHfK8984dC3n9C6D7d35QYRCsw0kwcOD6E6k7Ohgwuu
VbJTEvhLojSZuZmheCRiJSqWbAAD47rpsmFqKTGpY6Nza8KyToZ6qxHXO3ymYvhM
eYNYnW0rVzBCN40uvWaACYSsaUu2VBYUEtoit8xnw7rQJJmrbMLdEsYjAWd4a11g
m5BDcWHwGyo54Cbv+zxjb+4SdZXTtYX5Jo+g3lEmTh2jeJFGhSxwJeGYMCQrwMSe
1LsUBC3DAN2wqYPcBi3yJ0hAV2wz94hb2mdxcWRsj2pz8Tj1//ya9XnWlD0X4hgB
c5ZOF5VbxyVaHz3Xn/AmWO3SO+00wrW1mVken20JI2XeDXM+oS0fH/x86lUIiKeL
qRFufv6oaYHcazvNAWbA55bEROTlw7LqheYIvRMiLogJydBdYaxLpsAbqBGXRYDY
WiBRLYVTpklefxhNdPJsjo/gN3g6WQ8CnUFtWT935VFne/vnShoJ4SBm472bVqd4
fSA0sz9zmoh3ETcthNiy3Ob71XIMwNYjtB1IRWGyYkocrVUOQlNfahRDhKIowEz+
xdc8wLpl6Ga0gM6GxaaquDuMsNiOwuicarlBNX4mziP0hrpIm5gnzLm6CQc+r3o3
eRKogkxwaaixKmZjolJkdw6p9xlj6m2pMlsdGqrT6QEVn3rUlqRq75tErwMWsjoJ
o5t8xWTIf++B8YXU4ekC2CWH0ASAry0CwLzWUmhlvVlM5aIh7E6zusQWjW1ElofH
IATduKsIzeJS1L/+Igo8SZNPw1es4yQEzKWclz5Surs8YvnOO9tVvRfWlN1juPyj
NKzbAKEkJJEtj/ji4DeGY/vJD09Mbx+G0Vg77NzVWve55xueSJBJGFLj2aGEDOYq
MDax/zKsoqbxvIMu2qu1mkrwAjcb6s2K839Y6D3Fr3PXYzFZoNBlU347W63Ogu/L
CI40u71ECZeq7ZpnnFBo/4RRMMHhTAwSQxT8HAoJUuJrmQQOO544XN9zwG5nRaEM
+fnLtiCcIakomsP55sZloEH8VNi9qQY/TjSobtRRZ8i0C9rhOH0T7Sdf2AJ/ozoT
jTXb+nfT4FJIWPzx6rMc6xI9RevYR/nrnePmihSBb39ffcvZDAmO/CEJLbzscm3Y
wBW0gci5Z7EUxgUgz683PiwfbWu+Nd1J4Mm1OIuBG6vBQxJDd/eYE2exiR5C1IWC
HEfC16BAIiv+XykrqVVs6P7h9RVYG3AM0DR6WQLJ9F4ZFJ12FJcIwG+H3FIdpvcG
FZHrCjSwHzTXsM/IXvQUv7009iq955O7akjol69JbjuctXrv6DINkhu1f1YXvo0F
pc84ksFPmYeVQRFgznOFFixwjI8PCcZ+y3dCYjd3qWxQ4AiLi9hUenwoBXxjBHKE
HHR43ZyeW57utNbi4NYkzlHJacRi8zQ9/CWY++vn2fnGStyEyIhBXHDmUISGlBfe
imALVOm39iOB1ngUlAeaVP2MDsZWjvRxq/CF0KYrHBdDGywLpkULKqHMKw3SyKPO
21kRaNFqDxaRHld9FQXBOc4TSbx0FT/12pgpn9f78lExJob5wKDhRuT7UUvpOV2Z
X+w/Vf2ACbli9AIaCQCudshynwkJOO+cWqK+kYab1CcCguQgtdvA8b59V1G6tij1
PUhoDA3C0krI9wjBorL/PX4dyB0JCx1tZHZp12DAXMmU62diiaZmBdxvXcxRVfeN
hSw3PFDJfMhraxgKTnPm2U4+waupX/emRFUduKn4tfhLrw4xoJtKB0gqQBNwsRob
O7WsSn75a6wNfoIrtovE/vfwoApU1VAgv+AsgApr64z85Mr9nlGx4+sK5LX6lySo
PWRI8X6uaiAfSXpLAH4eANv+DbxycCQT+9lWD+Erq6p68dIXBqEa7qOVO1gYNJ3P
jeUg9K5qy9ZUDxEZiFnWxW3nyOHkgjiYuzhdMW874rQB1vgzoMZ/cw9YhZLkDBPF
iYTmn8ZDFAJIRL5QdySdA8Ouh6yI7QgjFaoO46fKwGpjTbiLq8nsokNTnmTtm2Ww
7jhCzXtdyhYrRptdwYge+JenFr37ZW+jCRU2LOf1FQrRjv3g15FTu4AF5IMZ75Ul
QT4PuY47ieOlmPUGasCUl+Ptu13S/d7zFRdCq1nM+4XDICdKkI9+so+VeFK7qwfz
w5hBI/prWObwk79eY9cJ9HTpMFqcZ4Owe4F7waK9WO+y5UeWdTPtcRrQfHipmjXa
HxLmVJEf45meIdoV82SbGwGwjD7DI4hcQTMGII9udK4PFwVYuKW4ZlbSPssail8u
0sh0f0maloU1Q49T9oK31KaDstASXvYnmcp4vWVNwSKwb53Ry2DT8BO7gIG3Scz4
kgO+o/lUWruMG3CtZt9nMJiEwpasY/gmfvnfxbkLb2fMH+FIXdYlWvM29HcnS3tm
JY/rzHMf4krq/diyblow5uK2ZxJk9F7i1CudtXX1gX+/Tn2V5gyJtWlS/lG/a5yC
8m4Oe8O+2IUU9HRuHaNpFgO1jT4zKWfubNS+1sIVntIfv2bX837FyUmzz5emoOMp
Wx+LFU2JSMQrHk7KB8/F/QShlsbStOhUBS3MF2crOkRgg517jCqBfPd5a2s6GbSN
7DGuA5ndOL/viKVjv6RJpkmgnGmCeifNj17NPsoIu81/TtyLD/8cP6BERBNyBYHD
z5L7lRCH0UOuoisRLECAkAGyMsnhJW4+FDCTxxRnIJZVOo4Ful/P1syRYxGIJ+5E
I/SwT30Nibie8V6pKBClYBnxqpSK5+vojX/QBJtCENVGP0iX3rRWw2zwreBRTcWi
JtXo/UnB16kinWOSNxlrFQYUhNRVh2OpZuULQlk1S39FlGxnwi55dywZbtmY7WsH
JE2E2x45U2j9vVa3w/qUzOLO/iVvGZZvVkq6f9lPFRZQ+7wA0shwfcI2/ZOVe7bT
aqbilv5er5wdvEiO1RqT/V+vnEWYFficv55c8hpNusTrWGYz+e1KkXXMozR12259
ymk6AacKJ0Txyj5MdVjoBBmpScRuynMdICSFrPvT/Bo8PpOWqMcbRXK2/7REHE8g
zyetAFUE6v/p3hhlHteWjQmziUo5JKda1YR+vOD1SKMGmTAu2q8VMEc1nFDiyekQ
U7DxAvhaZ7Apxs4rLlWtZJSd8TTfhTiYOVGJTn8ZR0KoLt8lVmJaWQnldIK13kQP
w/h2bmLMQfqFnjbHgA36k2pRqdtXtnzGWw7f8Rr8ROgY/fEpP2rDf8LSALjogPAy
Mxyjvnz6fxW+l0/cKxgS0B+8iogxo5JbqcnT36YJGF/SIfl+XrpyYCvD+KEfv147
hE4BJ7L6EkHW2fE0pdqKRlXIvhCxAReNI/eZaQYHSBCaVuT2cYXcFtrmMq5Q/Lef
6NAPhBHP1L8l51Pn73FddR0MBb4ZC6XIzk3hPKjiKvM+4++O3hEcki9Qn7nray/x
byY02aRxE+4OKhE+lr0sRxS76H/iUNHcvqq/4Cft49Jf0Kq4UISbbMRXF8PHIOPB
od4zeR034Iz0NOUSLTAfKysygxChYWJeWI6tFPi7t3gg7FCc2h21+SH3xmKwOlgp
1dujEAZsW7RYX1vCzlrfDE+/Np9vXy/w68GOUrvlnia1cSKnxpaBY3He1W3bjSbK
feNixbWlnR0hsJl48UtsMtd/2e/UiMID6AO/4wzvp2kVlDW+n3VGzNgSIdJB9kf5
uMi2s9ZPy2u0E9MwF5QWSTAOO41R9S5S93S7n5vXMW4h6NisA0J7zVDV15y2NWHs
GG8eVDiWVsRz3MfODapVGCG9L+wcP7NY4K/z+PKe+2FMPw9m9ISJmjuCX2FL2s2W
+UIuhR2eplgRrKY24A0EtWNhblCX1HYbUxPGqtLY1DoW7HatJF1Q2/wZL87af+cz
wisC2sJn6DgerJIw9DE48Lka1QsFPbtGpiJ/G0iglfY4/RK5T/DMHB+svR3+IROv
qW83I7vpa2tl9MPSxuTr2sKKbQTnzNWRg/iN0/jCWZvKMmzwXxf/oenihxguPPQv
I5EXI9VbaGRsRi1fYUyUVh7tUJBgLFoaO91klVhzpwNob1dyE6QsoVrVvfxFKCe/
zm62zPoS0P1WZj4suZ+qTvN6X8KNdb47rgni8/OEGahpWRZLmOWVjov3vCtLTWFl
L8x/M+GxNxUprJAPoqIRi8ZqHb2erbBq5V0gjQn/PQa5RQOXA87P5FDFzKPXBAAg
RuwkDnU3yIJeZ1hUyny6HMcpiKG26UeYxhbiJr3g1put38fdGyjY2oaZWRyDr9UM
hRfs54z22SXmTlJB5ahiQ6jL6BxkZO8uQUCTdOvk2ZQKcDg05DO/7g0wzWiQzT5q
W1uzjsV2sPzTIly5ZadxpW7fxkAAFfOdUULKsaa34Aw/AUMr2hDaQhMiZIk1IPxF
RTOnFa88oOu+lR4c8LlRCulrmyxUSXdvOHyJHYzAAQi8y60w6NGfuxani/f4BE7U
ejH/vWR5wrQrXpKiYEzwlATz0dnFXK8/VAwATmqek+vygpSSWZ+ofsx3BQMcmNEf
nYBPRbTKwJFKvlB9Df0EcHlwbjQRvlsXtRuFV+ZiAyWXZSFy5n+ynf4Qpe1w5LRU
fRWxOdvqpE0AcgvaCJ6TuWkTVLonsyOmHyA8BKMK+43zxg6jxP1hf5+rpFa/gVVR
1vLn4/CgYkVJi3Vgq1onZllxmCeHH3mohj6ufrdPeWGgSNCz/c7YTp4U4M9ugDqS
LGA7v745tKVrk+GnDU9Z73EqTVcgp3laW+Lv5k4xNmwlRIQJTG+T1XUwoHLNVeA3
xYX8RRVsB3/D4j8e2TKi6qnxVlI3ZWWmAPRamM1pDGvmm53mKgY/wFM/UgvBbj42
OvR8hB3hEoI5Uu1GlgO7ApJxMyuy1GJ6SRVTL2NY3x1NteviHjWoQttsDD/+e7/N
9GvDFiLtGcM0wl5QB4cm6SXSkEBh+GP6GRZXEyXF7l2H3IqhkCzHH29Q3oefqIMS
Gns2WpWIw1/gBLNbfDBqQufupAxpRmCKDWK9aGqRVu1BQdF/O84VJ4o3u0nhzt6C
y+yIGEKd4dBIIgIiVN/D6AUL0PAFJWFJSqL24hpUeFaPd79zYE5BhkRJcZBfDFWR
jAqlMQAA/rJn0aEl2c4gQc/G+624oelYc+MG5C7TGt5zTfFd0Pn/PIBNCkcwUwoH
XhcLe/26+KUpxzXNgwT7cActJjkygcF2B+C6l9VzziSyhWtxTANP3UtNXtEXYUUv
N0TG3viliJGhzKifT2MQr7hSZEHL372w7dvSYzXGxts0w2Dr4O/mZyCjW3nJ3cl6
h69eh8clLti2neVRoUkpbmkVvg/RCXWM8zmt5cPF43e3dU0FhPtlbnEBUPba0m49
PNohxF5Fn7Iw+Q7ulIn4tuwM/1jfVucnzNevSTiVIrreAkmSFvABHEuzpCDVkLQ3
0uW76C9+JE7IXV+7iFAQAMSmNnNHICmkVHmsNK5TvJjM+oS6WofLQrBR0Me5jdwd
JA+EFFwukDKpJoKVBpxSnM6TPidVkJcBxWxt3QXJk6DUxQyz7/KDdmZbbo0YUzOQ
7cURAfR8G1quoVtESzrwcmjCyREwVOXOsue788AGSQot9W+zbDCpuJrEtX7/vNVE
IZekdeq1EZNzwpjsglrEHDbj9WEhQntv2lo1uqvFZ5UWfDDHj9oyNDh68ffrtyo7
rKsxiKWc7RUxdr/FKC6WGetx3Kw01uAUYAd7ucgpCwBD0CGuBVc/gMMNdTfQnN+3
qtCALap3vr13qKVtKIyIVp5o8MoL1QwWxw+w3tSYgEmwl0bHo1515AFCjBZ+4q+n
+AqGKGcaepoAS1PTXcL7QdR0PByRCQ/Z2rw+GHH7cneKzdw4wqdwmVZADeLI8o4V
OqKCdbaRgSOVxc5pHHDjWurQw6t4kr3BQg/e8ZzwRtSRXa4uhi6HBuXqjjNHzZy8
azLezmYlkse4bco3u6+nXWIkwo+9SL/2lfyMiogudMbqAdTyTVNLNANQoviyWOs3
/H/lzLWA4q3mCXPPLULRPTqXOvsE032N60PfnJpx+w6Djl1h0U4mprWnLXCQRFVQ
jYhu837VKsmrOcB+61Y77nReYuIYz76AqZxKpm36JqVpAn4myxyB7BIWsBOG3hCu
NCQHH5a15AquwXWBcXhHbxCb7TSPP//prjxsmqXnIc/Av4rznVi5XjS6Xw1SONpU
y0wLios9uS3S8ej4jPiTnjSgvH23M3VoPiIT6+4UQJBhfewM3vJLd4hvTkcpkHDL
MjysVXRqWeFnWZ/ekNi5VNZxuYOcRSvjLK1oz5ZQwW+a6KH8fjKgVmyOLQXD/97x
9Lkz8YvdRkjVa8MvUKByoByu52GR9qUTivMpqhpOqjnwSiWiW3sGGzaLlYJwxH9d
2DU5c7pGweZNbZNkM3wXie5G4sXc/YG4ZHczYlOjGuC4rfl9CbkC7AD91QrMblfQ
Nw0EU4DruP8QU6dGScIGL5lvqzzPjK/1/WilG9ZjbJD0PQGjE5QLa7BWTbTAwcc1
KBjsUz68HmBLj1Wu5coJVbj4YfVB/8EQGIiYX4ZD3lvw02XaKybCLTVWnBzViyvM
CFLBlmIg+mUj11A6I8leobGGsT0Jjfg5mEQdTBSluQVUOOAMXdqY4x3uDj5+SsVD
8A3sL0s4Gi7AtYX2+WO61FeYfdAOyq/WEhsadz+2fuqOQ0ISZCjCthnP0+vGaXCM
OO4OV3KFpX/OxXjxWs7HNlMYnQZg7259dictLlk32fvVctk844bh3W8YkHo9NwZ+
m9x9OWR0YBSE/67QX5NtPhr1D+nWHsMkSirUEUaTUT+lG3N4WdklbsU8LGGZIa0n
1Emhci6vLdx6u3FyXMQC8TrhOI42gPxG3ORwWULpouHHqXSKaCezUQPR5bfy3jS6
Etaqs63GuIZhwi3d8wLgpPagxt/pGKm4Qv8BaZuOV6Dvl76V8mrvtDYmjCosKKpd
acBX8XEi3iFtWV0XuT4XQ9PU7ShVcEQsABLNHxlgaDIZDF8Z8pfg8sZWAmJu47Gi
qHUWU5lOcgsxf2l6q5t16GELpj9POJKQBK7FGIeR80xE7ZgZdcYlkQSQyrcJLfr/
wrZEd/cyWHN+eeMCdvP4aYm9LXELibOl77GJ3Cvdjl5SbznjwG/KGm8G8ELtiEYC
gH2FeijaPmAmnXQo/BXaPBZhjRPcp5gRDycMQuRhouBzCOH78UcKiI66G0jwb5iH
Jxwp4scyX5uBGLceqo7emVDrc3iMUa42rpMOAh1Gx5i5wOH9pMp282mgnhlOb2I3
zoAAk/U7iKaAwbmRjc7UyNpM1ioBneLArnuLFdUcrpiFEszwGBpuaGbhGG23ARGV
tLz/orVydOEucAAeHVM/cA7snNgBJZYOOi362tYfiHKE3GNxlub3hZq53AOkxXwu
7tgxVJyhoK6bZmYyI0eMozSWmAFeqvpAhwj7Kw4cryIvqd1zw3/Viw66kY4vOxS5
Fb2ZtKDswckwWxSORseMKYY0VF8oCIuTzcrZxRC1DnE3Ej2PDAxRk5J0mMmSnnUw
AJ7XG3fpWGnQnAwbZxTMV+38Qxd1N0SUlKLfBsu8orLT2XhtzAXXry3pf/7lRAkY
EfywoZtvq9ZwoGwfiNqaDK7je+zXZ1BcMDd3enMzUOSjDGAYaxI/3HSLZo/tKzlf
BkfKEGiYZUOxEnYpDMGKL8OhUh25OGLjjMsOg+nOkWn9WGs+QKqbzefkOQjgi50l
k+5FNxxU4Kblp+qD6xQs5Tw1oSqFKVAvdP9uREcHvLWpDwOzywl7LC6wnlvakDQ7
c16fuBpgqtY3statZU4qtS3iYFxcYLR8rm3zIZjn6KA10T5PICjERViqdA7TF/18
8rWO9sLHlpys4UUO1Ub7vl8D7KKuteYmlHlE/A7yb7VZriv3ubbC4h+X6pRP4KNR
M02+6z1mjsibW0N0kMymjf0y+b8QjIwMqO1RMsVE4kHoPV7dCtKMqR8N3ctSen96
yv6Uu0kIyq7k6YG84wML78HuZQp7V8uEIb9OPZiH15pBcf2YwN0tYsv2OrYxJXmg
vrlY7HxXdI2DcvnY1Y+n0me9PdQb4oAJ8sK8SO6NsJgvBkJWqhDZycOaf+OQqWpK
t3bNksovaaf1mIWHncWvafdxIaDpWD4xx4pi/78jWch6pQq0kzA7qBGye7x5uHNK
p90AjtZdrchoHySz149Auhh5XYaNIi0N1IxmfQ9V6rDUwcU/+JWhFtrCumgbM6kI
rUsWbrNTKRydr0Og3CC8pUtdg2wcXo0mcysrf68diWUIx2bKldKQZ+TCtrSTU8OK
/pf4b5aMWHy71p49FEs72SOv/CoZ0QJeexc8APAFGJr16l6/BYxZ54Y5Y23Kj45A
VfH79+7bDMnrTWooqJrBkVEeHd8A66R+hhGESbziVQjUSDADZIrO5mFTuukUn2Fq
/mCZexgEPtShJU7Kf8IykeQ8AZS/Oqih+vC+6bMp+7/nV6xouz/5OjEwlst7VoUH
+UdUm4J8y/VHq3G4x/0VoXYwqvHzkpMrJmdZ5+yivIwJvoUKrBjIeUomkcROA99G
m7pZ8PoDbciEMUmDktSHjGX5a7gmeBaMk4tUWGRFSz/hHoH30ryqi25ym7fNscIT
5brBZoG0OAT7IPfzUqiJwDYTY7rFs3U0+/ODfPILuSoF4KiDKXKr8SDKZOLywJzs
MtNE7WCTcGy+VrlhRf5OjLze5eqKx8E+Ljmu8TRyTjv8ZOez4/RtxnfQZ6OBcVvD
Y2j91cB2n4LzN86cuVg/t3wa67TCTwpkXaHTK6Es/KGZ8UFCmFH74dw9aDH0A5ST
iQPq1w4xw3VnukBduW+W+CKyJb6YlDuXoCKNCPibLl+f+/lC//KqwAN0S+gZIFuP
b3nnwCbuJpYsTVFNF5rkUrOHQ/iyj2MkGtbDRPH4rtwirWDBFYUl9fH38pqAeqo2
tNGpStJOyE66qDRPcnGTXwK5C9qrYmpdTMso3jQdLuFx4RNgmTJSCmd7BEpX3DJX
ajFEFAm43HuCMXq2c7Z7tAftmZGOEpCbr0EWtcc5+G8RRXl2Pq5omEYeCjY/684Q
qJjOHfG27zazm1D0zsLqpfQCl9AvK/kkdWdo7g9SFFOvcsznopMxkSkQufC6WT71
HnlP5vkz24bmxHMrkNK6HiIJugnSmU89D97btzP5diZ3g7kIxmukcyJXyl2FSJ7N
pTpb5Bolji9eRNcSHINwLxRik+cJLNA3sXGbhVzXgT4yhBqOd1fNfY1V0smjJXzR
OKV5OVFT0eaBDaWUE8unFru34sL9pORFfOsgK2yzTACZRe0k2LTAP0vEi/AdJSAy
fJCCJqpevLTWiDoT0Ac5IHjeTkZZSpCr8U/RDlQM2n/tjLSQg728plwFbbAkJoyy
v4/lwZ5vjKEqLt7Uc7W8spF5GPbyHh1ooSXpv1zSQEl3k2zUSuPmdGdOZLduRf5+
2FtnvB9LEe8xfpl8PBu/2cdkCxFa317ryEZm5NTD6O2dU6RGx9msDjipve63uyml
McC+h5f0/0iIwvIfteCAzH4OBt5mqBjfvfR+TzR81vuF/d+p6KbK+cq5RmJ6gIRs
M4PsYbNGvpR41QeTHo8GdLqr2RSLOWvibwg3Q5dB0qN278LfawgjGvptPTswD5Nh
Bihy0moo9qywtokk35qQ9fWNwcpzqnhSpC0vIJvtMiBkPFNOM1LgUQWLTnK0Y6w6
EnkeXHrudt+KzLHs5mPaWvSa1Z9VMSULwTZTh8FePmIBDSlwSof91CfEbplGjTNI
0V2Qjm/jZtE5yzq6DdBMO8PNmbr6aXI1JU10xSmNJJRZ5a9GJJlPNlnarkrOtkzl
l5CmYl9C2Iyq9lvOlj0ZVsaA1CjYzAvdqPo/8p+HdLNJl5r0bqBSGzrPb5wjWmH2
skQ5dbb/8DV8sdPOY7nu4bUPg0tmuQWhubloQkVHmKZdKbPuU31XPLJ8jkNU21zS
YuqLGgPvyperuH0Y4GCWvbUePFYgIOJ018tjIyQU9+iWX63Ybxu+0IW584v7XmFP
Ti3sM2O6O/cgfMy5tWmpYkY/vpLZcBEywdjB/XVYPp0webatfd3EbfGGyHWB8rKj
SwUcBUmYe0pO9aXeLieCtnD6ROxViherduKdCcfEmzIg+YZW6rz1poLoS3dotZGc
V6uWbRcOHdciLs4jhJUS3TQssom6u76NxjLa92TI1+YV1enRolrmJVxafT0c6rlY
lo5QuCXLuymolKQxQ/Y37UPdRBXnCHJDMagLbFV3oL3VUYwAg4Z/tT1XLeUOl0yb
wddxmjv6zVwdd+QLqp6RNxVK6TU41Li+BgebeU6CCWrInP/T0DGSqbYHunvBYT0O
6okgbTkR5wypYhA9RZilcq931/M+OFX2Zf6CgSEXevWcLoBg4nNjQtdf9fPN57Xe
6jld/4SSG6gu1Y36Z7Lyu/MNb9v7KkfchsC418MB6sHaKreAdnHVdRrcuJjn5GGW
Jna79dePeDcU3LK7aYwV3k8tN/dX39Jfw6NW8rJ/jTZFyUIX/BVaqIPiVMO1IP94
7OL5W7UDszMHcK+hJP/Bn5QhfK6Yih7Ia2VKeiIleemhZoMYS6jl8sig4OjH9HkN
xBJcrNNnoRilfSlSPSp3W8eTa9Z6i4Uwg0/4PLSZTW2a/yFcgIFWCw+2HrQuaWHP
lvoRYzg9/i9ghyE3RyYm24SnF3qMGhiVcXHPei5p8eHT3a5ktasimCl+JJG9HbZ5
WyX5zAq5zlG1eHwSxZtphJtfETWL83pOUv2+fTClVaRPlq4O+Nz0rXXDsBgHcVma
pcyS8nF94gP85mIetbf148uzAIKfM8q/IKae/YD/O12ih165kxAy5J6kYojDaM56
y/hI7xThALezla4qLXik79ZIB+zmwdsygSHOXFasIGxv4OjR1hGh70kZTSiP2RV3
QaTNuFu9AokvtzrQ6JxSxtosCSDLyjRBxzQAa58RlnPxr0VZ0baqPy55wsi2cglb
FO5rmrO2sY3buC91pBkKH8NsQmnskbj2UwLA2gL/jRo6M7bN91dAct7U/asUuWRP
/1xqn/kWUcwbo2bR/NCCMvPpCBaxYyLuIwyqFuuxGTCq4AHVsLbGZLOis10VuhKM
WytBvqKBITGHIhkfuGoj61IERc5MgS5gorN9XbfkauSe3kszA09RQiCrQU4vOpGM
GLT546xV11AA0jMbylPM53A4gwrn4GzviMMhy1V/3vAuz4kF9eFbruKpfj/fMZ8x
N6XlHdQKsC+QJlMT/wnxJgBTXUKZrCLchTyqQzc+Jpe15Z3s8SK1CSlsRib/zgeA
TUcsmytOfPpfdSncWC/PIL9fRJGSewSLOkx5oOTqR8j1GbDqNsv698yT8iqeBIAM
fCeL2RCXAOWPPR38oj12QSDR6wUPVqCTI2p0BgIE2U9SJax/WheZOT13EhfV3rbl
Eb7qY9dz9vzeSycUu+VMIltN3oOd9ViHzLKgCk/+Z9AYPuttD9f1mChZv/4oBo/5
rts5IgXOSnjEj4eKASeeebp51EPfj14y9g9fEd8r2qCP6MYfgo0RUi4c4nR4uoY6
zbZKXmIAeG9IP5swWCi7137M8IfYd/Fc6pU0MFBCqV5PU/zGs5VbJbc4Zl18aa9T
ow+OZkqltD5fvvi/bDHCJy0knPdnjmRalC94iyz2356uevXJW1iPzjO5ufp+0WSZ
s0FO9SyoaZ6neTmEDBuMa/ZJsbyGsYkMdW98qae6OC1Ck4640d0G97hM3jpAG6Ay
EGnOEVs7pLP/Voec6o+P8KrIYdw15T9b+uhjpmbyTbB5UY7EHKiVr+hMW38Z1RaY
bn0PISiA2yTNSL87ZnHe8js5pGfp+uIWB3oUQvviJfSML3sEJz4aX5KUxMjDaMpY
GYY8E4uzY8NS1TfmnGg4V7v4fgeQpcuWiEtNkoek9oQqyRqPBc8kaoOu6ucwNLMh
q/jQXFqShZDouxtmmvGvS/UpQ991qpX4vIHXZUhETPHyZ3S5tisBu8SJSPwGTyvi
AsZkBK3+oigC3VdUzk/Bl3zCv1IBOj8ivZcYoUd3awL3kqLZHJhpFFh5GEk9CMsM
DflU0zuVH+LvIdd2RvdyHeWp/YTfDy0U88P0mVP8KfgDjGY8DiOzXLcT1w6zCLbJ
TGnuWf8AMt87l+CQCOevExRgo+o7noM4XPOhzlxclLUP0AIo70hMOhMDusM7IbEU
rr5dnu07Dx2z3XL3TYlTMtaCZuYtp/SnvF+KDN33qQJw3eB/76qIL+AdMKNdrdrE
rNE6NnVYQ0OFy0mfh6/e/asUeCWf/nFEgIiUJRHVGBp1vEXjyIOQsSBNc8YL7yLJ
ejoBCnxqOOo91t7CvgrxPgx2dn0HY//Ue4mdc28wQXJROcFPhOZR4H+VqC4f3Qqi
zoBjRcdfI5KyjXMyV+1alRNJ6E7Bfs1IttAAJ7ml660ON2rSPUHvR6ONEdWijyf8
DsFOjrbAvMEg7OhzwfM8paZF23xt1GKrHmmWFzZ8nhNP/+Ns8qB5m9f4pJUZbWjE
TlNMvIuN13OOlxTAVcCF0LW2luWHt91Z8RbVvJfdjcODPmbWVMkhInxyO2faXiEN
dYv1XgHavoKx2o9hToVJXZGlYgOjm7sl/HnJu8CPf2MGselHsxSp3oJyyytbHWDR
d2YoNlHtuyPH5ii83+xPmQui1xqgSjviA87k+i2o1GMJwo/ML3BOGGf3epXFghzG
KWbxJs901bG9LeGIwU6sLAfR4Gw/hoTwA75w5GSiYLbbAFZQSiMydeKDWxgYeuPi
hcueOfJ+wDFDGSLbCki340e/T8TY2rUGDTiJIkvyD0aGYTuxit6emc0jSIldcjrG
Ni4m+xjbGS6njtH4n0WgLM24R3H3syTs8bDTvJwb2bcLVQsmSNLdw9gO3puQxLc8
LOUHLwni0N1uuMtK1pkS3mxNFgeOBoKr4agoJUQh7FLOlQI9RacIofWnbOE3b9gZ
LJhlEtW+3A9Uk5V6fUsH5SKYcb5vJFH51kZSlF6C5abf0FshSSfH3u1G/2Yv/3RH
DdbCDDgsEI+w28y8/Wynu5/gbXPyngSrw6cBvOyji4k/tXXHs8BBNAFAoW9d9VPd
5IoMlpnQgVFZVlAaLTPm2bE0UwgbmamoOvOiwXa+wO/l0PgnKM9FrPKMGft9zyZI
pZS7jtlT9Nu5NskDfxdbF2OY3/JB9VJ0m3nGasI+y38mnZ5utILQ8M1BR0FEN9pV
VQaWLYcLCuw75EVYTSQLUcSKOMhGCuzrNq5iUAmhHBCzfPTWiKh+VGorpJbrxBw3
uHzRDPzTY3x+LBTfSDShP9mQCRxm1KjTBJoMh3afrAecv7VGoKj9e4sCHOcum023
UeM2rTWuHy3rlwcT7XXwwcfMi9xIYWI9ilyZ0e82agLpAP0vdcRmHKCQB2WtAVij
Htm5MJT47oUn1iHyMjtoKW/24ikAtX5Jnn7/tzUlDCjeSe5toLhbnuPSA0aNI6i9
KzPx/J4Al1MDKBqMuMWwzuWuHcG84FXJRN+SJYVg9ZXzBqin99fu4F1mZQzyCHt6
p8dnToKLgMiR17TRmK/UwVCpQRTbNntPfGy9Hb6Cu9bWj6T3/KeL5V3Leq+lNSXG
EScnzc9KzRaXdpmjHNpJBtsqiUQoUvxXEcZZ689BW7L944Krv6DLxQcptKYYhoNt
yWmrz7sVwqZ1MYjpsyM4KG560sjWgVAK4rybKUQvjYnI8rKyUYTaNZm2h7zzcJxy
e/DktzGcucCCZVON6OJXFDbd8HdMVpqH21YFqeHNrf9D3MLG8WpwtA7Dv3ihrNam
4npJxn904NozPnjtXmGInM3MjaNIP8WglJBJLAX7OU0iOWwyZsPfYGGpUnKjhNU6
ORV1JK+Na3q7PATuEwhLnX2SVjuBvIPymNZwK1GXJBfU6rKXk4DzGHEUK7QqtdNu
dSt3dY0FjmYjqvP9sIC3hn+O14UuS6g0xrQFV5ZmjmmrjY4nw0JfYrVTwIDcocWF
OD95gTrTjUCRbN9mImJto24IPBWQB8ZNSgCGRb355CIdAUjqta9SadDARJkNga0K
wULIZxIGcyQzeIwFRwJsOWSLF72HtvvW2yjJRHnkwVEZCJmzczW2DSFSrXgUbA/W
o2zUod+3NYvyGSuqgcCsqYoOZ0cJX45l1OfJ+OZPSN+sRtJp5d+WK/MTEB3LE/mw
MtNwhF0N/rdjN8HE+xxEZSZ8wMwQsMROzXO0ysE5yBXe68+Ig3llYPZhSi2liTRK
KxaCGxdDVFGyxdTjOhuTl09gR6nv++ZtRmqhY/Z4maBKvAJt7m7GA64WGUv5gy0T
6qrVn806xs5BKXq0wMRWkd117ugS1sYNLamcLouj30S7+G9BEQz28kYfujYVZzMe
fqPmqCJbbCtMbv0Iq6wKX9bgGKZCGaZ2P4U92AfkPypumyx6xyuLXP+S1ZiVQ6Aq
nPMmZXxquv2Iau4ukSsFdmVONcpcXth+rFflr0lvg9ylyb63zhErGq5PiaoKLm4M
5hBW/eEB6Dev4R2/zCorC/OLeUmDLvJuwkO4xTBgQ0Hmr/Yksi+HqrCYpierEl7Q
rHXQxIHaK4dLz0xyDFUOaeK0zquxKzp+B4EvJBSskTYnrM7MkJ//J8CP1R9G4HKe
jnObCTdE5aYQXC28zf2J90HQlAFkk8OUAh7CH2/tnksU1XEgO2UHBuprT0+0iKVc
5hNazXpUpBW+AWRsZqtTuP6ZsoYFD5CI9hyjphfgdhnD+E06Aqc/4cJTa0W2Nz1C
nS2HSGZG09PTr7v02ErY3LVtJFGyNmrtSPBu4FRVSoe7MP/POBy999oV4vlHIRGZ
N2LMKV99a7QVHO6UMIHiA7wEBxtz0mL3tjWh5XtK5nRpDeFy1WZTcOPD2TIoC31e
1bLRnNlIvwn4xp9SdfcgMa7l5GpUhliag/RkrKpaGZM8eeWXgfsmDbxyfR7v9iTO
544HLlBjc1ntU2p68XyUCQbZlFVVaLjxxM8kbzQbSnKXGCZkGMPH3GkmloixUjEB
fc89tBRZn2bnyHky1jHbf5G6IuOZW5QFnTRUL5IWKIWeH6Zdlw45wy28Vbga2UXY
4M5/B6FeHzuE0QzG/UHSusuBBzLc4Ku1foXWFJxnJKUE48Tip4cd8tXMSpX0maqM
qeIIgEAMoq+IKBPQ+qswGzKKqJuwM0IBjnPCRSHQOrom5CC92VzK8eIwCsntvQe3
fqciutUYWfsoTIhZdQjILRUkLnd0AANTgZVlvEhH5/9IlXATatuUMSbf0nsJeWa2
JQzJScrZW5F/oeiPYEwDXpiBwyZbGAeoQCJvfoCVcTkI8ye7k1so0Q8eQqkMmIvt
qfRjcKyAgMYRZOBZtlU1/88P9HT6OJzUrUtxE5darwMGaJN3ue9PkhF3buL8W1WY
mszsv+mxZrgG+tjLa3G7Pi9b1DY4aAqAeEsIbao7GsKp+cP9Vfp1isVjaW8eVDA0
uaEFaxMBDoQILXy5BfDoPOjAOMi7BaecdMpRxM7VpT9ALytsJ2VVD/mCU8C8Q6Jq
AMgt6RqJXzhD/mLAnzgw88O0fsT29zS54GVChcFG0wUkvnmqyScaky2WRHkxR1ar
JJ4cxiMWbaKbWY4cHKymRQ0ThRRq/mzKSaZGOQQqKWGegKhBglQdVp61n0E3bED1
BVnnUkykGx7GGr2LsyxJhN+uSjFacLz5L0ZAdxWqtk6sTYvVDVdctCL3OVzki1ui
/4kwJoGYh5rtT49fS7H6qURjB25b+KeDPOAFd77CyXDHtC79xo90IK7q2flzCdyo
eKW/pZW442+PaoEpbROrTskMgJ72FhOQz38XlSl+QcFFN1iApQLLrEocC+qhBDeH
ekiITN7Oh9jq1oAKRc8KhjTGhjEu28pU4KSmtHEU99ovj3fX9cQJtLUxcKAYVZQC
ZO1pGNlZrdcmh9s7Q+zGel08FUhQcP1/06gMHYihU1O4syRKZ5P7hrTc/mdrLorV
B8gJcn4IXeK55UDPFhvcdarPK35u2T7O6vf7bu91wymIU4Z+P6hfmSYQNJ+jyfSu
EkNVQL3CX0FYw3AAjAYJRtgQLJ2AJ8NHkETTjTy03AttEluXI3l82UD7qrgGzyKM
g11OQYJZ8sQuLbb+XJJoqCE3ytXDMGU09uEZhVZeqDJNiKnJZURGm74mghKzJljY
Q/QbX+35//V7HsBhKZ44eP5nR0tuqzt+/pEyhmGdVid1PYDNDsWuH+ngGok8/pm6
ulBz7O5ekQ4PyOjIq8kdPnbsWs+nksU32bMapiJgt+f/w/p2g2iQcDRHohwJk/LK
ToLVuvnxlx/JQzlzxhqLK2I1f0FwyE1BdlooLzy8OX5RB6QvkLPeqm+hxi6wyWxG
RW1LbOADZZSxIyi/P4sDPg8GTvYV+06du3tYf9fpEMEcyc/wFQH38FvwKTNxukny
B8xdIeiinwJ2n+L+Lp5+riMbKXM/Z6CCw5plLOzffdbBNPSr68H18K5C/vTpt/0B
ueecA0g65AyQLBwjC3qtl3UZnlOCyD/bqwAqJXSbLYuI+OUpYVgdULyW4eTuu+uQ
tL3rBNuae+s2CeOa0nxDcXTShHT9CCZLrIyNgGMmDdvumKLj/dRZ9D9IMipEDGF0
SKV2ZFBMAreeke/rwHrCxEPwoRy9nyMMAF2M3Hun1Wc2vfdMjEKbETEQicrCJLQi
sAh/ylSQn8zTOivO5v0igU/ib1VLtn30FXzKYQVc/fGWQQgAKWmyynAfPVolOz83
sLHULM8j+2NG47T9FZUBApx7ETdRf4LTv/2g7nkh0fv0PdvLfnQMuUfOQ83ji7zJ
SS+523/TyxpbPAfM9f/0HUZdrM/N2n73FsCwiadTnB/Dca+64ZSIm2dTxEAwVXz0
CrO3asRA2lrd18g3ZQ2zJYgjcEPp4SfK1SnPODKJeB5N0MiIzO9HHeO/bb1hYr3V
mlM0re+tGzA4pS3dlArpwfa/cilufGDttKdYs65TMb20eO/JT9S06+xau5ZQmzLX
tadhUGChII3ELVkj7/6RI+3RGu6fhdmmYVse8dpgYX93zA1NGCHmDk9lFUEHnMGQ
vi6kJ/Xj7M1RVwR4B8aWdHmrgyvAD5WLEkxw3MEq/WuaxigCLu4T62kqnu7jxcUc
6LVX65nIzqV7yRrVq0oXZj78egU1MWhEHQ2nNdEafpZ1RWPe81XVYHDUzChNidSE
Xuq1grJT3hx1Y1eV6+wBxSDbOPSO/8mzUGlQZPdv9uVq+pG+Mcj66bvTavORZRFE
sd0MDON+B1rnPq52Kl8hQe1kjCA/dXyjJUywLGEEBFKSUMHSfNt2Y+UQKHtN1sjT
+IAmSAg/aHMgS+1JofZEb60w/c3oKICO/+LkYOyCQLC9dznHuvRgXDpc35v+xmtU
4Ak8qtqORH/ogn6MPqZot7tRk8XXcUW5tNowWJef/gwtcplM1gN61sD8/i8wE/ii
JnEroyVU5CSfaGaXi08VBF93LLT3BN3NdAUW+Insws+6eT3iz9K7lWZGLqz5jhPP
8EN18TROLMnk1VQlPyaiFH2Nhqvl7YhPvBrh4h5wo5Y8I+nAPmaBD8EyW6Lkw9IK
O8N4g48PMENcbCwrj/9Yq3j2mIIFoTks8vMHdVSb91eRidTs5kceODC4OD81alwr
IXWkF8ooT+gLRTw7RT1dkpTOFjekp3qUS9Z5Vpu20yMre29J1HC/USw9zmSrr+Ce
NWs0x2c+k5rhgi/k5BPuljxf/7gNJ0komHI0kCCNhL6epGYb7krI9KO9NG4vKGZH
Jl2Ks5IONVLP8XLGirKUsHWu9lmoQRTLNz3wGmR/zb9pG8eE8NpLHpUJfd8KPh1r
59ylU0QgD4lcwb6EAEKwDM5J1rs+LGJsgn45fp++xgUt+TvcfVBJbTx9qI7TjGDG
c9jUWrVCr25yzNxPbf+BWROZgGtivwtyo43kfhXZkVz1XfUbSpw28H8b5zOeZCOR
0jnQ9cgUyh8QOdrpTcHdct+gcSZpt3p/FaVaz8lBLMFqiO6o+52QkMNFO3XE/w2C
5+4k+Mp+FsBFN2WkK2REXnmC2r2/jVZL6SUXN21iuI2Sgwj3wcJV8umcqqjJq/Gj
euTn7qBoTITBS7a2NKCXFxyWr8Sb7cmYTV5kLHRQh5ajGh8dq7GR3vgG7oIPczQg
EkiZrWF2xWFmj3H7MR4eeWNPdbHBi+RfIr4QpmDWySRBqEpHnKwJ0HHkjogru5Vl
Sqfk7kAoAGNQ+5A707y4huta9oWTmvz7uSiRO144BymAw+4IgguhYoQCh3puPjmC
fHXLwjKTNC19+5SySiq7p1uSK4Q9uylroOTfpFUhjSiHQpZbA1ikyv9H5ij1v7jr
rynqY0DnQi2LOFUwewntw1AVT8tWGukLvL5cw7AC9X4Xmm84XuZEKXB6CuBIk61U
drClSQD3oPH4+1xbd7GakiEAHhAV+7J+z77aU4Ij4rT8C6Y0n0kz5xEadY1g0/nx
NcUqnGO8/Xqj8ya8IFVv+ywsQJ9vk1f8klJlkHXlGIcwikiV67npUU72YbWcALzi
W4vLqawYLpo3uPJwNYuMi1brKfPYWrqQQd4n3ihnPxn0jH4WY2JvIynoseZyMBsH
04bICdoUyuVfn+XqWynSqw9ZZIvCwPQUmpb2sN3M0K7l4xPgEr8lT8p/SXKsqi+i
PWK/r1qaxaDI+22v6DWVppcdr1gb7jpEEIuMSRorAr7Dh4nW4kHx18rvuoNoIQN6
XCMeXQmMxfFANZbgPSYObcpnH0wW2wKJ/qAFRFBd4V38YgsadZn80WLmnmzqChDS
V8xf6vKYbF4aLHtupq/Umzz/Ypi/KdkUSk9SlNcwgZP6xDIY3k2vvqDRBLePKzoP
++3r7Lxg1TY2NCe6okRJXa5N+UINOjFcYHA+u2YNyNnQny5ca55DY/8pbEjBF19n
0zBeVQ8OLXnRdKpKgMDVZrMFuWAu+3BAHl3bIiYuEal2+GdLhuAv6sjvcDvGwY/q
mSpOVehk2+RelrMmmWJvn0EEqCY3lbhuoQTXe5Q2WJT+EdiTF6cvvNvr7JnADG/l
P0z0ohQRsxMgpGeYMexW7RGE8I2ryBiBZvsetQgRc74TPp5bsPzOzGuXfjg8pXPz
pUlxnJgWEl/zOukH7RXLJrBmQFmNK/D/VlGFWUCVCYLswPcgNEjxyAPAVjiHTei1
WqQEvDAEHBmwJZ64xafvDX088NHSM++pRWkHxlnUSTID+JQaf2zixX82RhmAVzDF
qAWaJh4OLcW+gmERLfJ98eYpR/G9jHGxLYQtzR1XpSeR8KvisH3YdENMGzBw7soo
Cr8itqiles/WQfI1Y6ms5zuWHGOJoF12cYtFmWSSO1IFMcHd3+n6MAgdPaV/4prS
mDWTPN9Gw+4MWylx/yv7KGReb7IEdb7tyosi8Wsl4gTi2rgEfCO7w7EFHaG1kXyB
SZ0HLUccaC1xLtsI9FDNYyIB324z/71SeBnNxaWcTwuF+5qSKgk7jHdwAhWdykUD
TkYJTPsIP0Havq5EgL1W0jNvuOO5ElefDRaoz8xeTylymPiWhAIE4Kgu7HFvPByg
C6Tr0L3O37A4rUNXjEZwRWaZYy0r2mLNFvWMZOxXUsR5O2xW4nJD5FtXCS5OUROP
jMCHIEbOiDivo8QaOH7hqGLYWcZ1+8NGhKxrH4uF9sE+rOStRXQFZ3c8q45orOe7
7Dz9cJvhsuFV2pWRRGX2Q6tY2UygTdJPuk1dXbw0cvKESqiRNIaXQYiTqyPb8ulk
zyGNOw9VuK7Pzv2SnSBiBsjwXzQ2ZijhRTNhmhKSRPrCRXvF92YV8P4u6f7sOZP5
i27I65vY1/lmvIYWO5HbSlHCJnKFSD3YugNWguhv4pBI40df7bWEL2I6xIcTAkVf
9BrV4lgFXHhigcXSRDBU0slGpZD/JTJ6LPXYB5woyUy5zByz7sxEs5ZH4uFxezkP
0W7HrlUaoCadwApUvADYBdfhGF1kLtPFK0yZIan8ftfxWm9ymplUYyTJ8NpRiLi0
2NaV1Zr0RFoBHJOFqGDfudRfaGBChWkAWwQQUWZxvy1w0NmQjAc6PekflBH322du
QdsqnWuvmpeRu8gacRNRxgtmiBbSywGXPwcF/gRaNf5dqN7AVr+WPV69C/uLLCfL
cAMw4YSa6/W2fm0iKJbJ5k1oognvIFNJWFPgIRywK+gqzwbIf1Tu4bLR+UasWJMl
vXKvx/jXJr3ivzjqb+h2Ue7CIKmO0Azd3jnhyWmXdHGh1vAvoPtSIW9zOV5irE2Z
El6HwAKG2fU1ZNCtyj4jmoT4qbnS8ztV8fHNhffH76a5lAMP3Gox6xHkkCvVQAhG
JhMzqpXXOIdvzuvMIjIjTDFlrU8Ge3YcpvN5CaiBreci8jh7BML18u9Fmr1D6VO5
BJlawHmyS+sPEsBesUO72e+xxJ7m+rC5nVdmundAT8QNqwihXb4GF0GB0lL/8Um6
F9SjEOLlwtlvucZqo1mu/wFRZY5VWWzPSQteZpnBvzycegVM52I/l1U1dVeFKqvv
eXOZGQ3lpYM1Bb+JWj3EZZRhrURjA2VMgFtuoagDoBkKum6IhClB6X5K88HuEdQH
bXNNuaQLzSikWJVJKg+VhWcvpXGIThkRP/tJXDTAhpc6VROgd9YOXwz4ggafZHPN
LQr3/XrBzSpKqvqtf8EU8nUN+UOShC+kQfnqZONj9gsRNtVj7AXJL6kihYLI5f3W
YcJjoCnvsNlRSkR5+1TJ96gBYnJ5yT/1klXlLw6wQe6IvtYno3mSBuBSp+FLtA0f
CVnI2xXmO/H6XsgmWM52TGqS0mhQyHLqOigglWsLO1Cg80t2rvvYDGHca7BMKY2K
Hp+z+jKdY38/08W7tfTaGiEaKZJXxRci7WV2QA6i5Q5daukB+zT6iIykrtiKJq10
eUHYIy9BsYxfU4AAsORgojf5lyEllUAAby2zmtgp5fUnaerdVvbhs7BHNYH0KcgG
ncAfir882UX+pYf7JMOvK0V3ax61ErlS3GEIq05GVadV5xmhumaZc9ezoU9lXsdG
AY7tO0SerW54MXwTumaoMzJaRo7aXhS9WsSNtf6rv7R1tNRw/shjD0psrek7W+Y5
YdXV6GQ2oalnWuHbrMTE8WzRwsezo+GGj8E807y5YkLtwx4Do22z6uEoK/arhNbO
AznF13ORr0dxvLbW7+Ya/xfaW8uYZGRz909WnMX+ADzdNKOndd652rw2ctSspbe0
j4eWmm0Zzte1sBXS1/Yz+y+V6sCPy9PNwRuhACcrAqOUXidIZOdg5BdV2MlZOceL
SjTmkttVfdvncagXBYGMfzqiiaoKd8X+SQYF3iNUkLlDY6OKMNafYzaLFWk7W0zy
aGdB6Hm0i74dcUAUGkauoU5DL2J44PtGJslojBjLWVg74eiNibUUo0Gbr57StqGe
+1gMxARwymFt/JIVVdoDoE2RUTvJAVw/7pH9saOJrqJ9EXwKajiJpeVqiyExJnPM
G+yRwA1Z+zpjEYXuMuhrlVqR7/0n1tap464Kzv2QLsvuj/dvpakyyMn7ShNDalNm
l8IUjdukGnz42cnyv/9lStStko0DMuDaAeJGaorrNPWzhZk2uK448X2WbgskjOci
Mm41/42TH3Gk2fBWumAtv57ssQM1N7v/z5M7QBqKYNyQ4GJuWlOhBj/RWGEYB8uY
L2pyFHFBJlHHoaQ4rgcp4MhOMo2CpAMnPxtEDLHOGvlximZ5jJp5ep3qIpA/4V1G
imjGZufxdpCrhGM9RW2qQv7+GXKA3F3oihllZQlm9B6k1LjByfvNW9g9BweYc+w4
dBBND+NMpIkuNxNlaePC+5UDjur4PNA4SAZwP1V98bzp9YH4004dVcsIhQMfpg7j
O1YQQZGHPHLq+W/NDQBRBDykQVPeX/Ue32bmhQJE51qe4z9Kx7fFK2kQ2MWKy61Z
tqVIvqtystlLggKvAb1c6MTyWSizdalrFIBbve72XAHBfA1TXZbySn89SCydb+K4
QK1GASH8EHycNZW3OA3ABHV/Wc9fS5p70fQxpJiRvdI2OyNcfT7aiD32g3+T2KHH
UQ3TbYRPYbgUxuyd2AvK9iT4FdW0BUd7miazOyINnwujPEgk0XXAjMgEdLAmzlW+
g42kHIaMLpiNHtQQNYSimsgxoqR7Lw/VLZFyTtXUIHaAhQgOr9haYXAxQ/UN/dPS
GDJopQnurSd+gTvX2N57tHJGnn94K8AyYX/5bXR+q2VgOKur8IaRk5cV/pfDTtH4
IsttlwNUoZfp2uDcYMACFnJoftJDjgkEl01YkvxQnckxetbaourFfRRStM7/B1qU
JXqZ2wjmQ9epGoR35kICS9bVGP4kms4CurPtyrV/M22ye0d92pOSsKa4MYYHOQYk
bDPaHvWjBdvcOfBj16W1XnrritpR7pGgTY+p5MMGPe/5aqtWTGu3uQvOKeR2Gboj
RNpLenSQ4/DccTNYGGA8Ck7FsmeARqCJYkjzA/wz99vK81lpWQVJzxvSnkTPRHKs
yrZX1fVGP0w4sRmijyg1+0QUdoz6BLTOLB90cX72jD/pIsNjmZZBH9Y/tt5GUhIq
q0fbG1DbfzGi+L6qGDJaKw1Qezr6gAMxc7Drzn04C6fPvCyLym/bQ3jXmGOcEy2R
OY0d7oQPfxDGYYC0J8S5KQ3bTtbzMkcSfaV7lXtFrJEGg/GsPr19Gk3ooT+4/qC4
R7NGrourmlvR3/4qS8PTqTycY9jTatMIR2Ru+opd3DdEg+mOFnxuz0ukHkuDDOOj
QN19IRWn/0OarbWiqcerIjofMvYOcJctUw2Cny+ow1CAZn32PjjEkNziZeHrZS+S
aCIAY553y7JXjA9pOjxNmta45TkXyJP452gM7J/TJHa14Jz1W/84hNw/2IpdUaoW
R2m6TYlQMhGfHjmsXBJdh7bGCbTF/PK1K4JRIMAV10AoGuoJSMK7az7bn2Z4C2kz
cuerwNlKO7RqlhHCPasBxyQ0KBRb5fzcufLAwTiLsKKUnqbD7z1dy0XY5NH4lUyc
7nVH6wypeNo910WNEeldK3WaUSoel1PNtnGPyIpQEdGmaddyX1bslk/Y0h+sMUOJ
wAqfu3gKixes6uO4EILcgseu3TyaeK+N1LDAiXOkhxpGyti/XV2M1C9eRQpDzwYb
ROIrs6DFBhmHwnHvq0eCX6CkC8cErRG2PqxTdI/Bf404P9fn49Raf0xt52vl8waI
dEYHeh3FtGGIUuIf9XSbmVTBcaXMZEMFjLGrPf3NfvpnZMFvTqnt5QqsXxD8Uaow
LZFKIOmXzQTCpUxvgj+B8uAqr4eITnrijrcskNGhEbhCw5WHbGulh+c1LsQhOmHn
eZ2U2+2DKOOUh5XlLH3phfQuGBQzFbLXXsKjn87pjpeAvQy1hDhZcz0d2uUkys4w
1/qP31CugQlKl91ztLYruY/odAQn0+Z8SnlqZrFyQ0zonHVKHXBetgMqGvRiyuJa
Y0t3CDemOwct5eLlYhddWhJ3TGO1nnFebSkRl8AUKzlvRME0PaLF6MSaFbeN0HNI
ZcwCKCKwGMh7ZC8ZxYxaFW2vV2Wf320cBuyo/p94b0x3OXo+2/L7aPm/tsJt7KAn
Z3S7QPkXKSvMeT7FV7b9ukYnFPfzreBLQgR7PXiRloAOS7ZCs64OLbhmJVrOS3gW
ovUBr1cvMzKaAudE2fOUHJ5QglOXPhGc6iqCMcyObUoHrkZDwwikSVMjXdPW2zjd
tXCRRXY6bAoKmH6EtHQTpSOHgccgPa/Wx7Wk1vafiJ4JT7g1BerpiKE05fGx3ItA
iQmum4MpPsZOvLaCAwkVR97vIWFxGVlmMftsqh8yzIfS5ODeUsWLoh8m79lo9wUp
SClE7tQ+RfWEOJzrOgXzUkM6LmIO7h3XvX4qiORM0K2Yz3f4sHz4C4wC/rK89o3f
wWCRmSEicTUildwmvySSR+Kr2RkiNkItcCbHs6Nk8NtLbgNx9plxju/KkiJ1cyX2
N05qWttTceRmVw73w3l8wGif9QghSPFarxLA+EMFXLkOFu9yDu8WenJkyQ9wqAC7
c+ziPWPJEVA79WSCuDY7IucxnIryQE3g2aHJG9dq6/c269GelG50y03cUGGFR4EM
OcSjJHiglZmCl8r0QLTSXoF5OYvkWz1AJlAM6BTbZmHG5e7sac14c1yFCCjIjZZj
WJ/s7Yfl6V5yK2WQmlOWcVk/0HzfG7uYcL9NfKoF58tWXfrdFjM7KiMZPEDCR7Q7
4AuaS6XKLlg6+D0jltWAFoTlIvbpUG5acbVAL60t0cdDpsbBtt+2mB93iRT3ZyNQ
qJ2UvBK6a+HjV9ec4DxNnFcVih+MYjrbK6i6HTlk2OVL0SJywWcfqPF4jfLMjL52
I53QVJHnypV9sGvfaY2pnV+H/bq/6zYGNiuibiqB9wGb6zEBZUsJBzDaaitGdHMY
trT/+mMjUGX2J9qxcH/eTVLNXMawSceQFpov7w0zvHLIyFcSlTghzaxjc4vwoIcB
gOqeTLORxc+XVqhgevBPgyUCg9dHUWROrKcIopVuQLF/vuhoBIFE6aFxUdVVB83W
Z64n/Pe9UnUIp8WCTjKQQd/S6jhC1ybBNN1uar/AsTEh1spQDYS+fmVrEP0T3jop
+k6KytAf2Ki+mfKpERwdQGeUox3JeCvlK1rv2N7jRIkwqDUdDa7R7k4tLdXzFKnz
NK1lXg9tTRDTUvVSbyxPqKoCCLs+djtBhYMdzLh3LWLF6s1tWfnS7GWk4XLMXhR1
3ex8m04Ex6xcwR3B+hLve6kKuH4nts/xIoj8zu7k3WD4D0qzzmTXQbR+R1/gSb8s
2G1rCcUHQZy4svuDKHjlfbuN7QMJSUEvfBZ0Xo9cu2EP3mEFQ5ZgolsiRbVKCm6E
k7OAXjh2l/Q9CbH5QNwcLeT5Tfb1NeEDjckPKnci5+jVyOn8u8IPoq9M3nDLN6tA
pdZSbkap1Jf2j1KAUy1r7nbsc1H8/QQO/S0q5xZL66nG2sqcly7qICYFq311Dgzh
0k2MNFo461yQMSkw4vJupm+cOtEV8FgLPYkcemb3qSA4dt14iDR67skcrTNQVi/Q
g8w3bgwrH4SEOgxRzs1KWWPUQXR/YG4ZTfbIDgG9nGYC1exwJW4GFb7f4ELrzSWA
gyI5hrSS6xVy0qzKGfE4K78Gl4n3zcKmYfRB6rk5GhiCXPUjbOj3PfTJCtmwgu7y
Kf2UH1KfrvsPfNmYPZAihNMRBAu2ytR63n5eBn+y37C0jptpESFjvRkTAEgrzLgA
fJ2+jzoxdAyH+Ly06DXa49cJyoV28P+FN0anRBF9+MMNR50CaD6NAYYYj4hPcA+m
krJddqy7+G8B1SoDOmxwKO+BpyMJKObT8C0I6m0dbgq4HclxSMI92jPHzcQExJ4M
+9jo6HnHaOKFJsTGrFhjqU+mTTW5SWhHUKb+h7kdBq6gDVfZsxtuWrSOuGlv+N21
gSDMQ2pk4aGjbbuCEfO2IbWXWsl7jSzmVar2MIo0D05P4jxfI1zg1jKn/cLlcebL
fXisux9LrWkQMwlMUKghEnwFjl5mF7GV+KVQ66wayp7Fo0/9R24xkHAEmk+O9He6
PVxaarkKXN3qmKlyqqFvzWuIBvaZpWgims1wr7B1/KgE6AKWEQojizLkPGwSHcP+
QoQyA30vn7t6xkx9Loih9FGAxHffuqWjpKLbnwhIAp8hvRekwpuG/6/UEZ7GGYkV
q1OOiX8HHufJX2ibCj0YQPb0GewmdDuzy5w/sJLw6/zmq12ZklGUuf8ccbjm6Wco
0p4YyfURAeLftxFgonkB8u8zdPfiOsCeDvsc+s5zShbECMCtNrKVjNaibgIt7Oru
hdQvQUIdlwQFoJDm7USK+3mleeoGfJ+Wjh1vsTddg3JTH8HDGU6/OBLSprLG2q0k
vjeo1Gkr1rs5b+BRWTDKHcaoYKvE8pFpp4XdiFakpXarxLjB25dK4m+uVeLMrYJu
36mRD0c/HRR1C3QBMkhL4HoOtURnfG1p2CnU8cbITn4PiJh1uhSi0nGPYg7QANSW
YTA4Qv3XGitPoF06FfP72ZnQDq2P0pDQYIxqO2brUtx7NQIVs9hV+aod8y6AYZsJ
rb5YBtDdL1hnU7BOn582gfY9mf5AbBjX7yRw16gcAgzJFXG72A5bDVXpgBU/2t/z
PPfOzNHd2WFAh8SwyzX8TKdp04anUBtXKnU6Ad1ZePDYhmwNZQKMFwM3AqMiGhE9
a9ikkrhOmWc3YpIYoioJjEsLRNrYgGweKKkGsUXa+gjZKcowhtHzYG7MgLSiv+nk
xMJ3kgrdRk242N9quzoClLrMcApQqP4eKNjj9pFrpyQnbRAsL9daiyCKosZlxryA
E7eXNJy7HUhPEXTDiOGrpdAWqHD1ZSn2IfpI/k5o/CkXv85NR0oVtXk0ui4d8p9Z
U0W3U+6zaCUrNYQK6MPi5vTQsHxdUh8fTzTWRy1ACkwb2lbbMT+h7ZgBiVBTXLSe
l/5be9jrMxECeDrzR3dhw2y37MewhxRmciY5j4kD5q22/hdCDgA9khTKg1yG374B
tee4oo7ywqrFBbueqBmIj6p02CCdssJ4ha1Ta/RztjMJlmR0KqZnnlmQ/e5ygPsa
lkdwyMo1v0EpZbeEiZvVwpUBcMR4aWjcjo4iA272XvPflIv4KkgH1FiikBM++ZVl
f3nM92nAm62FPS6I35/u741MUYLASXeVDRARjF0lDij60iBVylDEwdlea2/n2qcq
r74vhhCX0gJD/1TnsaaAosxCEXh2A+QUSGrA6acclXb9X2yiXw3YWCPHmLAlBXEa
Z6ha8GGSCceYK9XBBCvVAjm3P2s3lzTYPNzgc3G74L0iPsQHtSQNeka2f/l9tbEd
6UQWaOpkiTxN1RJ6PEqFyZB++EgoKBN0vLDQP23s4fv+IsndVHCsbyhiqn3SYPq4
5XTAOT9ANDTnW6A1qkqrUQfxx4qZyhb3kRTM+KJ7zvdAvKxa6XIX2BUAkMyBo8Nc
UDkWEjgOM9Qofi/ce9cCjTfmmh8Y9QpQufj4DjxzcLph4FGpy8h258Vk4mNa+1Qh
rflS1bv+2YbgayEWm9+TMrHazYrbLEaX4PN+kZ3imnIUgKJOnFrjaMZF/OC8nmZp
F94LOJb0ioWkb8WbOXEDmlKxfk/PVr6KXUfACc1pjsW0I4POki56mCwb7KkUAPq+
IaaGivj74+0wt7gdRRK4WwpxxSn1hpLINoE4GHbVsIZxCMwjxJpqoL5LPq9444t8
5gb46L+ZsP1A5fyH91hH9Jh9tEMRlx3pkujuacJX38PQljyGF674kUW9XTrnlXFR
w43ZRg8FudeKctb+xVs/LVIgcjHq1K8LMbP8axvkqlBpISqzKfbHEyuPRtaiuOQz
qpCtZ3V3+E7JAs0zgEndBzVO3S+AMfHn5cDYjt0JRgy1IdbkDVepH5wh/xrkh2iX
wuDRQ/otyoukaIaDTas72q6I/gy/goj99e9eKJCZ2ny7xVASh8Rde3TYdc/QHMCI
5QsXoS6z49erfA45fx2eyKmx3dLM5H8Ft2kSteRy4z5C4/KWZQX4RxQnMDsrsw/P
Gwl/Dfu73emPRZmF7Yy2WDXwOoVrUT7/CXblQ+ONer0IQSDkReiAcJaNqicfM79r
U1eHLoWJMXp7yUL4Z+/Yr1nmERmjrKcjUU0ahmO4G4FWL6xunRH+LQo4oEk0Oa0K
1ikCY0odwr0mt4hjjxQ8SvalgnHMxvrloPkhB7scdXsD3QrieDfj5w0iOIuxbjfC
ON4vE1N9KMTPX0Q96yQ7ln99Rz9dyP9wHXPb4h2REjv/oeKXGJrWSszZB2qR49nP
W3rqx/8ooSmiJzvKX+0K7JBZ4dcjjMBQfvoe76MHSOVCpl7YkhWI6pVSMVeYJuWG
TQgtbGzbQT0KMBGB0HDfiSHHCqxp/N1I97ESbkFNrYQyiWN8NG/Rnlk84QY6sLHV
PkVDkKGcS8w7SyF8Vt4ecyidYMfHxzQCUNnCqIg5TdEx1dDqYWYm1GfT8GxMmjy+
M3jtYbwZcGZsl62SDyJKc1S2rDtwTr5wkIUoSSm1Y7uTBtBRO0ssokZ8zyd3NKh7
khlkxTFVOz+hKgdhLvF5pvLngDVj05tFio0FxIMuPmU/7aPU8ZcaUUUMccT5pHv/
+kGlD/kHWZfOO5oU3R33nn6OIhMVUiMEbds0ofCzjubT6h9k2PY+s1e1VW0vo8uh
bduJ4+rUiryRTlSqSSl18PCTsdDHaA7zaojPFH2NxMxeM1oeuP6i18xBV0toJcaa
gkfEUrkYb0TZ6sYI3DXyuQPkutALHNrVP3skibC4DwOnrfhBzP6AYj8LCntceITL
YSljxKeOqGH4wjk4n0F4lratw5OgnEEft+uzJEX3X1MGBgXMTbtd8h7UC9g/0jAP
AlKtd17RiVQK/6u5r9hrpCa0vtH8QSxa2UtE8EcMaFGlmmF9CcI21sQy8moMIYH6
Uoui7vv56SqNFaV2lYyMIuv5To0/GxdLaU/FrHayAfu1cBzKg14pI5J7U1cHgmLg
XqAFkg6P2UCUFj8il3xoZTCYIeuJL/4oKaqDM6QN4Z/HjGtROZWzOCW0rhpA60sI
N+XPtsBMsM+kAgKFaJaG18X8acZGCrOi/UOJkdXIGUAsRWAJsMBaV+5oghuQsSZR
DK2/Kcj+lDlod5zNElYxUEbw+7Z95mfINLTn7a/SDROkxVptk6LhsvzByW1z+e0K
ITidiNk6Mvk4c24RxwDu7MbCTr+9t0/wH/tUmrjrWFLypj/dOZL6oFwzTXOVFR5+
9H7J+Xo7WQI5RZUJbKyX7+5QcDBcH8fZLfHP2S6K6v2NDSEUb17J5I4HENb6bA+3
Y60PipxPN37qF+Vns8hDPu2LZ0sCMmUpiHa3fwRhkYbXR8hYZhZCZEvPB+eAtGWa
Wm3ZPrawfp8PpP56ObV/qSTYPM0MM1/twf2JQY5Q7X1uX80IrjCQXzKEiDC4SylE
ZEXTnhsvi+1l+xTCeAH52EsyfiLF7LgFiB5Tj0x8GBr5IyIPJHnBNqh94RqAYoLm
Ezb+hdgG6mIFzFQNlrIRc2ulyZOnB3DRqBbncDOXAW3GpdUFLqA48Ym/l68u4eAh
redHIdpE+COOM+nwgd10f+G/7988WAyjVqaCmfnqBBsNMVDM8mFXkQWXo2iY1YTf
onA5YaOn9W38SQ7iOhT8IwjNU/hZ7ngaF+Gig1fiRaWP0/l+j1saMErjK5xmDL//
a2FWkihyv9TfFXFML1/nJ4to1+o4Pe+2hmeSmtSP8qW4G1ShjwAeD2QzWcAFJhZz
c79Jcx1K5sHa0q4kRUW1JpZEUPWgsDP5mwuR0cu2GfeOA6T6jH/ot4rOU/gYA35L
OUYfR91dBmEJE101f81w1pmhm1C55CyhYW8XYB5BlYdECGZWwkdpmbGn8ZyFSmL+
1e1g+1pIsL9b3G0nZnBEf81BNq/Myqus5RTUyYtielzp3utL9m68XIj3GmqQqH9r
fhUeQEa60IurSlF8fXR63qDevfHVF5uA1n2+NZ4ej3xSpG7ApGpPXHhmS+iJQTVn
ePL6TNa2zZSHKVAsXm1mggGYSfVVstcHwS3mf4noyVSsqI7XumN058Z/amaGOx4K
M1AJVtH7X4YnwAxVSHz2fXA/qqW3M337xL1tRhpkFBV/XcpRzaJH18FRfGh9dTqO
zIPBtPK8U+iSXvNkcXjPUVhyGm2x4hIZusqIe1bPRNI6VoJwv7DNuYvU8QK4PYyv
QaN+DycqLHxbAE9n+7kXoYMpCUVH8sHN6uHno8i6RoDTKmcXzaenadMsO53imYIh
DW3ee3dOF5JAtt9QtAtQTcbuB2gI1ZxqUr6AWwxUG6hIaamVvRRS9oHGTYYYmPgZ
lUZ+9LdWHpTnSuJLnQHKAYZtvASJa6SBU3xuvq1za0zRLFUXkSks9GlEx1Zaj3BP
ZwUP4XPJMyhhHnX3AaY8x1b5avc4Hh7wrkg8JTMWaCMlflREepLWXrlY7hKJaW/Y
+9L9ETzrjQTFAQSgbli5IGJdBiao8IWu3q2K51/AB0/jVhxF/2SOGeFJ0A80EZDB
padHySo7CuWgmFqOfR8jrIJD2Ri0vIuLTiBzMk7VbxIuNtnlcdt55dt2cRpd6alt
XnArH1trZdSS7nV2wYl7oU0R/XXhXaP0GMwJh1qk5PJtfXm7y9b8yrA7jLYSCQW4
OBrnPy7qB78fM9c3Cvb8QSDP38B3/jl8/t2LDWM5JjEEIlgJH79pAqvgxrodMYmE
MHRa9WID3XPXVBiffoV+AscLFgKiiV0J9m5BcplfZSEwb48ujQfnhGQL0mPg1ftR
UDv7Y+S/lfwHYQu7Zwf1wq2zle+xwVYkgar7424ZeFCSBs8QebFKb2/4N54JNYgj
8tXRTWo1jWEU9qXAdRoHG9qPx0Pw42VFxLiJpp816Mi0UnNNauRY2jFeCsCJ6gTO
QbtN28KqbX/YUJy14kIIKAdnyXPH2+JM48+YMHd6eWtGa4uc2rKPM1+NjS0BzB3+
IoBFoKGgjGadhFCzCKeNn3c+5iPrwbuB89E4bgiDe//+FbJv0t8Ato0K2/6KFQ6e
9C4MwLgnQmfcgSV7uJL8qVB6BDKsIUXhAODdnVufGNBLw1mXZdCiFKXVxEM1sA6z
kJJvmgZKUBp0058OV0f+Ver4JuLgc8TDiKmnmEEk4T+gVPI8HJtrddtudOjP5Bpe
/zeob7Y0+UBF3CsYZekH7YIGTrmWW4+jrHWL2FqWFZRlUN0AtQat2wEV2plu3XGP
SHXxm0CHgMITPLN8p6D/NXkH64BoCG8DWeSFQmx9HN3QWUEdq/ZluYZEL63G+8M5
rbAr2z09LlZjyzHnUAZKdYYVD2yqTTcn2UiIVkAtefn84/bjdZsMH25gAlM0U0JB
GwrfHKkQ9YFgqCvpKUiQvwzZ7Di7jTfzyXVqXTwpj5n1GeRfMfqR/QihGjlfkQQz
VrOkONgRs7ISehwzoqxc7WiZp4i4T/qDxISKSwlsv0S6ra1RBzNsooj4LGVfljPL
T+69I+xobyWMAmveZ3Pe+DgHtCLzkj/2Tm3RnNyy5JYDl3MxYhXMKTgzkhABILs0
QrgfV5z2GaQgNd/5iZczb5gsVJgxtzSfANx6BG9wLOxVa6Zw8miHhdw0VTCBnHGm
xx5V+BlrXRMN1X2n9smZbHsHuY8Ls+BRH2IBrd5cVlnHiMj1H2cSmGzR4IhsKkkA
Menai9Yq0l9rpZUwqjwwjCsMh8XGyef20G/5BIEbCkcUA7K//vz+sGTBMv4bEOWN
eX+zg31Gl3KQZJxGEeUEQQciuRMRELgSLbcGRw9AW4Tl6D5hdaeiJM8+svhPRNx1
9+VCtqs8tk0/qgVBeluWjJefRmvjZL/WdYR4nYarsNRgCorJs2Zb0tF10fmO84VK
o1AaMx2KRM4VplninBqgR6KxWh91DjTDyiU3FADpiU8vB6vflUblQL7rnfCu2put
Y83gv1RUlL6dnyYGtYO1STLWIPGlcdc/KumsnB2Mxhe8jfewMS+BzhLuomnighNz
Aje0lTIA91iMd1HDHXUShHa6l7W8eaVwzGVRcDiRncOjqPlYKXft+SI0fu86ntmd
6eWNBrJ5puNxF7rMZc5j1QPMUnVJy4DyAJ+PsiqsWwUJxchomfPreB4WyYZaSDJl
uT/MW7vCcaFkXlITWkkfp+mqVgvvTilYtd3Ob+KiD2HqDCstdfcRlFwVVoTHWZRA
1TkMj6xoIsJFfOH7BTnEPCBWnwJW4YTzRwIScdsZFUxcUrBthWkvU2UB8WrGMkKQ
W062qubAu6Xb6R/hIsQ9hfThsppF3P93hmGS3PWaZLgidssSobkVHFRXdqDORe2V
1lk3YdwSnPHHTemIBCUbsymj3Z4haYpqJFNt6nRFCNxyhHYQ5ai/0GGT0i8uJYpV
VuT+f9h5B3sRH7CoXdsmqN7WyE0S5c56uX7Pd8Xj1YgyjMhkmTR+82rxJbZw900s
xWwYA2j4RVSGP9wzFXzH9w/tsyI5sFNm6IW/o2MWIF/t9P44D8y9kkHJw8RXRm+F
YXUl6t/eLgSVcFPXUa2XQXQ9ROF/LrWgyy0qsX2ttGepz+RlW9T2IoZtLAU9Aob4
zfo2JcZv1VUzTYCUpIZQbBQu7+mscs5iu/ex28UkW3PpZazHsmjp/n6ojS5ID3TT
izieJq08ERev42SEVJeL4jnevC+g3e0Ci1KvmCOEUFmxA5VAtommnbUlNq5j2fD/
lzhERN/AiU/EqEgX4uOEemuOwihJ05xq+9kJbquF1OCRJKeHT1wv6wWGT44G5LN5
CZUUCNlZyT5pH+53j1jixU0F0UoUJN9oHpNk/P8GdObJqGR8naB6C3Xpzt7IojPa
bWlEVHb7q3n8tKY0AHpt7XNqxIFI37ATfrGhzKt/63385sWRx/nUlY/aYloiWJ8m
RBT1YxsYR1e6cHAhghEwNBID01PKHFIUqCRW0BUp3Vubw18fw0XaAKW0uofT/zcl
E/yveqqyQdvk0WakhefmvMwNhBMt/OmuZq4ML1FeO2fweFqOToyi3y55Ovpxtw/u
fSCrC+1V/+j4h0iqj/73Tu8PEtFp0hiRzmaR6pfo5FgTB3/IeR79n/rzyXpOScvy
tpD03ZcrScZczLs649gs7jP/vxFTXY33MTjQ0cW1SPydOCspXrzyrkqn0kv6MjhN
PdmHXElEdMikwCSTr5wC/pUnpsO3GBk13earhtQwomMv8kfywR8UKz//O/afAzLR
OsOCWtEiTt4jWs4CndK8Q+2JdXklJCW+HaG4vQ43XZvSWKuKjly1fSn/K7CRXXIf
q/MnCi9nrH80oHKWdQVA8e2ClrdfarYSUL06sVMJZOb3M8xzG/SNUXI+8Nonvzzy
mKYF3+8rznQGXRFOOyjF9UjawANVh24dMVhAUayuxTVzTKfUXXjErQhBsnEIja51
prnEIeTSHyXvGjJu5NTysuR6bxVvyBGSjYEOedA8Pxj1U35MQRt3/Ec7uCQggmhs
JOs0NVfwP6sA6S+/YwX7XhE6anDi1upk1DmMSSrbJ7mvUcXMWpvkhQwIbY3tY8pw
WTzn7JE0SQJv3Re8f2+5iTmA8bnEjACGOuRyNe1hNJAA76RyVBRANXID9KOpjfCJ
7D6eWGXyx3boaFECFlWlW5MuoR9ikV7hfVaOOQEKxV1FBUGv0fNbmjl7TtYkw0mb
g0H3dhCSM/dRYg/p7gaM6cXipdWa9xcxwge5X5WaoHvt9PulPb0IJ8Ak5Hoo0cvx
iaj3kqs0dgqRQzWkhgVEbvX7a1Lku0dWQ4jYlshj1HmEDl5i0aTZerOlfbfZf3Kk
w0HhAduiuDKPhgQnIrnW3s1j5zdm1tuLFiT+2P5DSKc+PAMqJ3E9zJchOzBmLBSD
xkA2SgH1sYh26HsyaNwVimmn4wlNgLzLlw4Alb3dgvDU+xH/ce/N1fzphiPZgPvG
k0uUbS/rxGuT6HN5tHp9TGMufQEi5BMrggE8CeU7vYOFNQEyleG1QG+dBhGdKJbk
SgEXJr3+LwG/LWgyJEi7k1AIZn0D2Hs8uNrcgXt3ukEHCPtbxwirAJUFLZV2qaZp
jchLfaNl237s/W5wUbVktX2sWM3/ZnR5UgjEcgfyoACiEkVAx46oV395GtA+k+M9
OyBx9LZHXeccv9DhLN4GZqO03E4CBeJBuhTfJjtAQ2LZ5oKPSyovOkAyzhCoaGJv
F/vw2b/iEDNRAnR6NUXOpMyebx134XqSAP4D81AS2YbOBXm3RTCy044y+BrB7vAE
8CCUst3WPqFVEcIPrWh2cVBQsdwLijneXQP5160a50pb07/juMXTh9lsanyzUXIG
4gNorgPYBIEhly8FyRyecQiCj8D9D0SH7+2lx0GKzuGETAGMyhtXbOeNqq7KI/gI
oPQ2ZDUyNXWmcZZ7kW3GcWVmMAJsqW/qq9iZVKslPTu68kHIjEOQl+dd8RENEMYk
9C03MMAZOjJEigbjOzWRNww86IiCcF2OTNstMJTv1n+geCS4mqgMagiz2iboN/ho
WD/jusYtXmQCVkr3Wxvf31TVPWAN77mZMI9sMsQ1hwDQydlvvXINB5Fr1Eg/58s9
LTymOcaJ1yHDNy37KQp/Gf9TlRUO6fOYTs4GqQEKqp95a4rMUD2ebkI1LHDC4qnD
6q2YwyTjnPZ4pH2xxvLjv1mtdPGhl0EqFO34VF5RsQCZ8sRLTXEY+B7QiukS4zKK
yVr612s54tkphAHqOnSJJ9ITappeexngGCrBnkEATl/jfGFpA1Nz1yqc79hivM2q
YwCgVVqhFCuzAkwa2lHH+C1My2yBp1byufAbe7WadHSdcLJiqtWdGRN2+lU1dYOX
pqMme0I05eNQe1fVbEGmVevo/1rruNzULJNqmnnXrl/aJSSH/Rm67niu91Zox7Ds
qgosoyNwqK1BahMj4IPCkiXsxLtC8/N1BhXhTlqMzl7p8XkwoPOGTtMNjrIv9ff+
so8iylJHKcqBsY8KyWYeNp2KrHmZR98Mi0Q70zFumP2fq8UR2ExUM7hg3oojANOd
Mq9pqmQ8JgAIX8fTmmTGiKBbdHagRtd0yarMV6jl9quIWiActH/ijW6vmjFyv/DV
rVdXzoig0QTsBlODQHhsZTFsgfBPEtcCojRupLkVDY+G+uOjaqRtJT0sPTMMx9oR
m1mJxXk/OSCTqRBPt+ieev+JZBsvPXhWt7yUEQuGzcce3ZQhBhuHZDoZtA31k5oF
VX5gf4MbHc0X8EDCG5StEmj9vVPbB/3d6PXwAmaEjNKcpKNHj4+Aqw+7bSlDTga4
viqR0VbvGoyFYTqNg2tE/4S2WtM4MtbvuoLjdK9WfDeGCv1VIKe77PqUqbZIFdgI
Qh3u09a6GQdUSn7h1yv1UVudn7r3WSN5mD5xpUR6rkl+Jj9K3Ie9haFkCdH23u4y
C2ToEjQD86nrYRQbTQ6xUpZrqxxxa/80jtTNaXILLC4JmG4yJxdsIB0WiJPEMdrY
RC38hgdXB2C4Ft/1v61gELbjD10+izZMt6HzqUYgwtDDuNxdWvbq7m5hNmfBBloJ
9vOBxQIrVuo115E5tZsGAJ2PVmnF20RBcwP6Wd6JrFZsBZCskqI361L9yTZMZHmb
IqxivEYp781VEbbdZYDUGvONYfvrUxRVrqulS1jtN8UtGLp/xk1CKjDwNONBPe0h
h7/m6p5JTvrTN+jJcqofs1Dimk5+v5SwM+3e1vM9BDEf5l2B6pDcu41/xm7p6nVp
4cRk/dr5julv+7K4p+y8rCxYObK0eDXVgWjvaMlLEx8BH+pxTChXprOKUoAm+PAj
z6w2Vmiw475IUfQPWvEAgGVu5F3X7QDJXUd5LWQsM19hKEKeXYUNG6HKTifqFKJQ
0nwnOltZ/0lhgrwrERg6mJwI+KGe1ugWqqH6WaCSH15U9u5NvsZ6CTkecrrrMZnG
0z5B4iuQOcm/TuQn6dMY3yvNw1Gh82boB2lN6bYGyusOHYa0wiKon3wdltxy4UiP
iKn0OBSKrP+nLMVgQVyE1n9NPyUCd+dv/gvWICUt1yXdFYiszSnSd3kngVUN6o0S
YvQ8xTNX0GIkWK8DROPqi4tVqfHHdxm/Vnmc4cxJ7mNQz7nIprg3ieLfp+U53u+J
0Y06MUX2PTdZ2cp9NCwlZOispSBJauWqXGf5zOC+pxDS2IRwwWxfECfaAEt+9QU6
8RudhtPF46O9DR61ZJgny5sAJtbctGq9bzuSNiqXqN7ye8Bm5lQ1PLmqb0ZkmFV1
1DMzZ78slXOTGiuBU6hDR+d9x43g2Hip6XaKEFcD/0i8e/NqweFzR0cl/v85+5gC
HscZJO/VUJyWntBYCWcLS1KByQJaZW5NF5qwbHcUQnaD82D1O9QPXlN4uolzHYhm
WYdzBDqqPVp/RY0W1kdN9BBtSaJbR2iCMevl4IXCAQlgY7U67E4xZarnbIkT7Sh8
kDiDb1lnilL6ApzwTaEuU2hkjaJQAeyIL0/13mzrI5S9OO3fowkOQA4enHKJ9v50
LGEXSj2nAF5uofWscc9kZBHGjuxuvgGexk/Uoadg8C8BdQaixUBfzJZU4cpbuFPy
DdhuLYXPkxLkELf2d7jcolGXVo7Xg1RmXxQdId8d4zROJL4ylHpafBgLx+msSd94
82thY8mATmw00l5/b3XjI8w0/IgFsLDQKJoIkaS4CPGkc8zh8ZiVr5ePPlEeR8oX
MGxGbvAsr7nrWF16HfBeIp+xDl8GXRATEusR+M7VR8jBE5lN90JQjvE4DEWnsWQ2
qlnn8LIdJuzb5vdZjgvMTPEKBIpei2sG+Z/8cjTDKpf7M3W+CgRblwKXjg+wBWrD
nRNQ4XtVomYFmrvHaaYohTf5aIW1ZVma3qLMytMHszyAmzalp6OA/HaF1UdTXbym
gTmRTHailsxkYL9UOXzUH8Oa90XB3h9VJ+AiPojxfuwY5XBMfdGMPfEK15Qsb1SD
bnb55yLjGk5J5CAAQvZ9Hd3fchkKU206hmrTF+1WhlHPw/HOA8mLdE8cTXAXgLOj
LSLU5OhwwqDeVb988oB6RZDk79DtQ/mnqK8OKezegnEIhRfqUtZuUwD6FUbzMJqK
isDXHznqWs/IFWCvE1qVc5CAjdDXfh7+JdK40Trn4pkSb+heTQgkRHC4xBF3UaMy
Q8xK1emY3j0CzMau/M9WaZuO0DL8PzXQFeM0R0/BZBRqxXr/CE2YzJgvUHAr1lmL
m6qVRgkI02VmYDqs0iVcGo9UfbI+SZ5+0fpgPxMu7nSgEUlsE8nNLfp0dn3JG0AO
CMIegwrS5C7tVs7I9CRVJ31MYk0Dgp+r6LcP2ktFSqPi55wnjv6iK6BUHGaCvdi+
ijOF+iznJgyGSlSMWQRcDBKtNKkx2bgmi15q+0zFdNd89JDtc9lAT3Q10LydJEeB
wRrL9t/Lo7KAikVhiDbCoLsiGQKwWvLMPKoUhB1mcHz2U4V4vMlVjTuKMpJR6s5W
badp2m8hPU3PFoZqUynfTMNo+pcttx3LQkDo7DJWI/NtE34y2xQ8Mu1DitKihogw
cwVjD32j55045DrDvHefFf/7PL5zc47GDV3C1+pYkigTufKayUCr35jBcZhZhYa2
JIlpwOT80SOg6TPnVvS1Q6xbyQEQ09AGRb/7vZMiHUQ6W1CG+yjWGEUdLriYS2wR
J4o61AkfKmEeSVjR4C41dtEnFg7hM4oelPlx74swIZto61SBzMWv8IAUBQjSS8eJ
uyTYOhzKPO8XOiRgdisr+AVEHmUlwmjf+FYuiPZNgjZaDXtRPJ4kr37JLGw5oItq
Hj0KZh/CEgrsexFfZE2qDHmSQaS4+UWwwPeJHubMVX0tTDq5WRie4GM+uUxTO4SB
ODjnYHjvvZLZsbgz79vIyY+V7idRd2RffmbG570riwbT0l4ygTqnvUaqQVG5G8Pf
eb/zIAl0CAXX7zVEDhQN6v4jruVZ7MhTfBRHAy2qD/U7mkXoZsSXNBs0g4HsTXfH
MdjfKaqBdl4wFOdZ9cwveJvxW5Eqsez182WJLRzLp/dNq9dGlI6zq7mrl4dRc0bG
tF9pZlpOSUpoNOBGoRl0qwVdaM5y//XMSfL51CgGQ2o923VAb/RqKRzrgn14QE8v
wILcRLbKhF3zgNUCHMBnI1f85VBF8GRt4nOtMmksY1B/QWX5LyZwhm9quylbC9MT
3ckl+CftSiLVJn/weICNiXZvag4yvrfmrZFQOt9CyUPlK08VB/mf8NcGZ0UAHuTS
+Y0UzCNBk0CH8k/AMeYFyJVwApMFlfjRMqEkSmA4SqtkwzefZ0XbRPNIQ2fXqTK3
W0TkyKODsCHTzSUb78c1Pyf0A0xDxUxQoYKCIU+nVXkFwCutw/BbbnrunReMNuAe
eVjZkibisY7NnA7bmGwKgA1BVrSM1uQjFRdpVsw/bFIM8/f2mE5xcDJNDpv7IwVW
6LywUTsU3xzcilv2kuTVlRwn916KAMV6XYNlb0QHMZt3blqbkhVwYucX+v39ICyi
rWKrwz2XoNB/OynT3VOivS15kpRlY+p+KNKlWu/KG3B/PtD+5U1/C8jzBCDj3m3q
K1puqtTiSC1TNOeCJFh5JIzzj4uRWSF/Je2xdTqtycUHWJBv7RN9+o+BbWH5bWqQ
yuu3SoApi1RKQKOvSONY6P/nWop2CNfPfJEz41OzENOPajJbAT6JTO5CttBgCo4b
BTq+JC2yjsqK2G0LTCIuzN64nlsbKEYUFvPBN6tIat5wZpZXDJ2L2NA2w1AWVVCH
AkLINbdPiNopYtjbEns9T/+eQXB1WCsPMfc2dPB7u6GQ94vvqyEronIH9yUxIdIh
cUcmIOfO/kYRNmXDq5Uub92LIqTI0HKF8RMEVYRLfWxNeegOhbBxp2FgEUAYuTPZ
dHYbgZp1/giL+VIBnAUHQ/QCpDpFK9OETm7C65+MWpVkJ/IKuTIyf/EW7lab+JAe
qNegzIfwg2yslqFXzC0WFb/a5ATjg8lJdS+gcGyamUKo5ZJ+bbNZECRKzLUjd0sj
yPYhlcNhojjFC9C1e9MW5mF28Ym8uoc6YFHL/qraUo+soHOxIX4pZ2rgpUHfEWO8
xOVDyKy3CwbA/g+IczwvgRpWXdNPJzCICoRfWGriLMjCLl+ASBUiw+TCQxEZMbNa
4zxNiC6WP0jA4+pRgw9G6Z1hoP1xgG5GdfmONRmjrocT+plWn46KNbV6wAw5okhS
7k+LUjYqhKjgEK5z2TN9UcarUq/0EicOTDhT9nq6mrZJW4CUx5RKM0ZMxRBV7UKV
fbI+LLGZVySfe4tMCV8GPCRkVoeOqdMguggiLOaxRSmZOJMNoGLtycI7Quf35trT
MFKLk6VeHT783JhL1BZMcFoizk1h9S4GbHjDWN0cGMCuZfWv9MyjSI65wp9bIl1t
HJFLBWpuvUl3q5tpOzQjRwn875h5niJr3u21SDJHAEbAWgPj9k+ryCNK9ifF2qJs
A7XxjtQEQednabpwpTfsCG/+neGrA8CLf293VpNxdNAqKbKiYzkqTTb0oXFgAqpW
D9ahHyph6hMqgEETzq3YYQIRZpXiqqky5p42OSqhqTvi3+VR2aCnUy4Q+Pt6gOGJ
9L5n6Ig5u5Rgv7iY0ZQYUKKfovpkidffN45Va8Jc7dICX9eyqT8K3n1ZhM5cpZGH
2t6PSlznJFdPzLcyYHTDtczjYwg1kOMYGBkbqg+T9il8YuGrhaw157oLjxjJcLq6
5HPrt/J2n2vnRq3dwGCwKGsJeQkGJ8XP1BG5SAMkokA1N+4FVpTIRlOt0uH5yndl
NH5Oo5XKjcz9NeKro1Sc8chU30vDEbPlzIoYrWqLo23sqPB/Ey2MjRX8FauuXsIr
BGXLe6y4cIDBGLjoxQ/A+DEjQljYyJsqZJC0WuLy1ABuuvkLewt/MsObpcFidQqA
mGS2w3S4evxExRlvOAOixZomMWsvHto1dD50hZcdy8bHzIzDOMdG9sMl50beOMlT
pSZXQO/1I/ElzikAh4hRTsNo6nlc7OPl/Powqj8HWHSdTRBOg65YU71TACa/y0rB
Kdrrw61CF3ektJm9CTI/E1aOQN1za59i6lIzjWBEEtXbRfgRBYuiJGFgCzWOOyJq
cqL4tJf7PY1KUZ9SWqko7SRAb0jX3iFSFrQI+hUuM2AyDYu+VkLCa5h6S0Q1iWqg
jyP+RwPNYdGB5NW66yIt5P5aWGAN5dfMYA82llpkfsNpUg+J5RxDnWQjnGm3/6SB
rnOMoaYMbKOAAkf+9ZQu4fa+Z66IZcFc5lK96ovfwKtwoyaAu91JlMgTLP5ptj9O
mg4LxIEDaR05V7dTSIkWiWVEJJp2dKDVWwWltvHPGwn2fRWM3Vl8OsVftgo/2/ap
QHcNd78/P4iJmXhGxd0FlNSY6cxpy2Kc2mSzMxaRX4EmJ0ko0uL6RHHaf9IyqRv4
AEV8ATfZEy/c0cZ5RfLq6tkRwULe7++1+4zl1NjmdC5G7nVUHbuG5akTiHGzd42P
WF0Bkbo5m5ly6fKMDmBLHD/ftUqYr4KC+R/tSMWVw93INlCzmdMqoWgRYHgqZ4u8
UCUYyF0cwIiof2xC/fqE6ElTYsfjgTNHp6wYsi6nFMxUyH1Bk51nq/MC0p9ctV4G
3oMqeAwtXFjUQRC6da3TSHXQ4MmxrfLuT5iZNuTIUqsQfyIlXYofUpvmRh3jhnPi
jVwbSESp98uIUKcbTMnLHeKp5ikvSq//B34qpwudlIrVP/gNVZFjs0iq4o1BL6sQ
66Sgai0q/aIq0AHBnP/f/NE4ao1JM/lk240fdD9wpgmk12kbHFRJVNFo/91iOtcF
AMnrYHbvKfKakw8GRjfYnQrq/dArx11MAWUGTAzRaL4r3F+MIqBQ2CzKQvn0roi1
Q6YBYVi/4KmSzi9eH2sOewF8snPGBzSkDOGlwgSQ9a94xs2B66GyLFIxkCA/nfYJ
am74je+LZpviQ7Xdf5vsGy0J1VoEwdou13bb2E1AvLkIGUWGKajl97d5aQhs++9+
Yg9z45zuLb1nfI18N+SGjD5z1vcUq4UGJ1E4bwXX6csxvZ3Pfm4XLCqtYu028oB3
pZTgPpMGDSj5c6AauuP4GMeJ3+ZBVrNug0ExeU+QSCYeleGrAfO0cbrdW16czrAd
mYNQLovOcJyIY2MVm0sOLutu1sNQxPMgLxyA9yj0vsKjIJBIEMnZ9XZ6B1/QVYld
kqjroXFWGMWJvZq1VnMKcnSpaut19Uc90o8Jv86G3dAhjod/jjB+AMir33lkkdU6
mi4RMOC+YltHZfca06fRjYZterLuHety61k41dWqQJAE9eDq+sYQYigRo5a9xZ4c
Dr2FkV3b5xQJoun3NE/QuQ0SSUk3KNUTLyiGTt5UhtupFROgxL+5sJR6S9O4NnpR
mGXKcv1oLrRcH2qKWG9arGQynxPEVXUcnRO4Kmgn4gpk0OLuvJ6LqcERPyd8L7P2
DFjX4FVZvYM6HIU3zabsgroIeTB5dGNkQN2Dx7elFQUZ+AvLixia8eYI0LSk5zrk
coIFqoGJbdIVjO3Db9SMQOiLEW3VHtWWY33DyPd2JfPUcmVkoYWG5hsLeC1QDBBG
8/0u1TCnQIOJUjNlq6G/DLFjLSOB/50xF0AeN/+Fsty4Cx0Wbedv/BGh6BBq9v+n
WIT+Ohv0+l3mgJ99MruJ6GYatZb7jOaxnHVJmfwoLgblOQi+B7Zh1ZQs25IQSm0U
yex5Fsh91/ZvY7WeSNEBfLUmNu1b6P6P1pk0wQa7PyXhgTllGhIaHGKbTjDS4Kar
FkAGIKt/GXV8ZsxFGaUShBdlZDG2Gnr0FHgJIZdAEBN9k2T0r9bxZ8PM1FY6cPWX
6PQJZDDxajYdWTM2Prst20jQYEZ5ya5/UerN8NZsPsns0TGe6b8XNzEDUr5B4N9Y
swBOXp3MCav3/bxNVIrerxs2P4FehzPOrl66cCCSuORzb4uI9HvEIXii2Bzb39h9
pT43YCuO2fpSOoiuwzPDYepcbRBnLqkLU4dEM0KiofADQZecFaLgTaG0YTylUkKz
UsUu8fKvI0/reFK6fiPOKS++LvUy1jLZUEgGx4MEOtNsZt/YUSJIlAwzLQgcQUjV
/GxGcjfaq0bI8J6yXGp/+Sd4Ke1Q0se/uKSvq8JuhDKx7sXOlzXgK21cTSCIp8af
7NzBo5lkDTnLb+rN/RT/5c59/8wiseoyXSQW/VVIXtV6Wpl0L3G8GUdZXlAv1r4n
wNzjci8FyN9tHFCrfGmyAtwUhNcDanJAOVqFP58CKD8WXFLccMBbQTJSicZtKR0x
C0j5gB4ygHE0EdHvM5vn8vKsRwZrYpaegkew6J4dHxpYxeh+VJ52PV2HszlK03Tw
k2hWcctFYcFOZvT1EVi7bW9NRZtfXrcZJiWYgKDVh24u4JQREpxC22VSp3Z7wN4t
Wb2I13u4QiTxRTlK3eshXNU62lPU1YYvWpKWla3zaZOAbaIEAQ68gwqxqZFhUKzH
CzRLt7OSZc7ebPigzajr8pjNXE4ZL647tiHMVXuW0qmKAvovjlQ3vrYbGXpPoC1t
6Qgjr5ZzWAT5+9V7jV/Ih1ZIIf06rHq4lAOBMLZEA/f1CfvDfSPSxJ74JtDeGjkv
yKFPR4hU5QyBJ+FjqkjpkkU6qhw5Uzs1eGDuq+SUSsdhhlF9z8eBEsVV0+b52VJ9
gX0c9BP2rBbtg1NUwgJWjNngGDYcZGIacK4wGmVdfvtAxtkZo51gi2LYtSor/3eD
abyA2HN1Q4TmM9uGMplqF624GsUU+vxgw2etn5Ko0BZxCxkARBw3bpV7pTogNhxE
PrS9Vg3lJPJlXTr9jfBK9kpZ4e61GF8aTYrfqNzpWLgyT00P62IzMsbh+RJtY0vA
E0gxmO1RAgA2UMn5IO7d8UlKQJje+krrKrjGQ4aW3NdvvWqDkuSFz3tvQSxt7PZl
sbZb6wwPaNroLCL6+R7WBCdgz8eHAbJ6388jS7bA8Tr1ngxCTVhZqVoBjPcGSW3I
yvjWP0pfTco1Lope/AfHPfu+Zt6MQyL+j1umQGnrj0hUPVxk2MioOIBTNKGADVWI
NCIEqJBQonb8PQ7JFWI0egqdXdWbBgnVC0+57lEbZra+WhDTNL/54OS6hMrb+qQl
G6f+h5fkmAV46ilKzVZ+XNDldfCymLp/F/PIrlrumgOTU46ldWjIf16crK6kccJR
ZEfSBiJZ5FrGZGOuBurBizYUvwGLjWlYeAqsgm+X/hpg0g40f1wW/XYhYwQnrZak
gd4CdL1GgfzbnGJUC3l9gQCRHnDe74zcZN3HElh/RMDQ2ajPNlf8Qo/e/+rXi5OU
Zor9Nik67AfseHQkSoF4KQl7DTr/okEz9MO8YcebClLM7QMeLkZAOVlUwtymB7Vc
HA8BtRGuhvgPRPIgpe91YnI9gAf36Gy/81n+H6MKK9bCAe3iqHURsmcuj9s8wGxL
dhrVF6CM05Czx8hRoNg3lAb6erbebxtNuZ38f3VK3VDNk8IeKhPnSHb+lymaK22E
YWC2MEI213AS7/Tx6qWtjf04l+onZxf+EvK7++oTscSYP6gcqQyWjrL3V125SZsJ
LRkQIZMdWrib6zMrJzqKWTOgMBPGjK5WBPdHUaUB2fNlhq2gyu9o/jgc7kHu7WWR
I+szoMaXA5xODLlSma9cwBkQyxp1iTvchvs+/VRRUQ/DFZqJ+oONHGLMMCjZQnyF
mb1rM5B1bwp6mjgbcAEDLiKVlN/DAitQvBImP5/46aQILKQYgDX+zMytyQ/DrK39
PohtORed24efe+MW2Z9puc9WdLyAi7yD1QbrgkwkKuWauPXBEwW2I3ha8ZonvdPW
GGWus0o7KlfheH9TBWRKXZDZmH63poMcFYyxR2SMqH2dGKHW1estSSkWKA7a58X0
aie4NSNFBaXl8Yjg91c1NFlSWeLHSApv12iDcmZFhMmUWvZwLRbyT59UucneM4Sy
EEENMQScJQxM7l737UjRqPbHliWOdB9ffz4AjwUaCUCJ+7F+3RvjQOvev0ZU9Boo
lvkVhxa5UX+HB3QA5uAD2GauP7LBcbG2myQiffH2hKvseJ5Sxd3sYPBfgs1aIpXL
7JfN0rR8ME6alZaem+lVY39ExE7MPTq9SKXCzp50R3zX2wg6kJM0CzveWo5tYNjE
oFOKAoociU/XZBRgSTfcrorLH++Uv99DqRP4dlRmZ/vmNU2wvKXkxnu6+vDZdBxB
bp82JSFhjt44MrQbPRmY2WlFyEHHRaDs3AtBrJd6KMu93NbPu2iRgt8WcBXw2FcC
/DGBnPTOvMsNS/HAggocmhKwUPQqtbrqwMghwI/d1uR4mfMMFH3ZizXBPwqefujf
lfwtEkDNK6dQJkdlHnhuuEE+a2l1qHdNq2dJDBqlMmzv3PRF9oJm3pmdjGA7oFxZ
AAXmDiHr0kPSCVdB9Otn29Q91i2719salDENswy9PNpWeLElseMPwirxukEuaQ3z
UCQZradzZV/BQ8aySEI7bRMPhCJmUC+U91sYJ9jRtnH1cXKd+lDDuoMrYH0LoclA
iY4J6rTumoXyQl8eDta5IX1EM8KNMoezWcWx7k+X2KX6v73QfHYL2+Vi/RQmMUrI
tvqul/uHe2iVVzYHnb+OFOj8Cz6NoqqaKDDiBAr5GR1Hc8h0Y6ZXngqbegJVAaJP
7otFWIBXcQ6gwVetdzK8QyVhwdcFfNiy1U0YC0nwErrkp6pOvNWfRiMrpLWg2FjE
CKluIbVvlmEJc/BqgGsw2IqDXrDuCHVKijLKCUo3ULobsZElYZ4IzXPmQGzjNfbE
na4FZzMYt5RumI9tfKxJBZaUi5nX6YQV7ze+L7r75KFygfe4Fxt8LSyeD4v7q+ZZ
P77LfhAYqYSDAY7PWjQrMBtjfIHyXVSvAu7iDK67dTkf3ELSKLEKy9CaiMifqvYg
U84SqlMwnYLLYgesepxVe8DnKSWybBjMgveC1zEjhqKb9TQ9rpfPaP+TtnkarM08
LPaTpS2uyaeO8aKOGGIKsJkhg8+4i0jN9eo18X+PbrTSXUIKhWuAFq9L2t1AI1vA
QYzXypEmMQKfS07Y0NHC79qX9ZboeWPZEqc6E16TtvqoHYCzT7X4AiahzVsE0NN9
5uCpQwSGK05/lak+9uqs0k3+bH6xXL5FLjm0BnsbD7pYgUL+QXf2d7Y9a744Qud9
QOV0U8fGFACpHBzpND6pMANaflPWoBbDFI2s4NEPHc4LuPmsdX+AquHvrU8SGnsO
MQrnD83eLlXf9etLskiL9gidGXyxAcbbGMWAcEgWj9+91nWySIWNJIpUIo3QGWOk
83ySUE8M2uQP06ge0FpSUsSMpwzRY4BthGB5IpSnDGNrDDYyvtwsp7MXJDFQRK2D
nD6BqX2Bht2NCXBmBfgieHYW//t4b87W5JNAmRcq7qfmwBkjKhkrsIzu207KEBNk
ac16Ypr0nTFtI3vpFbqU/U4Ae9NDqYBt6q0Gxg/7SOXMAp9lZp1eHm+Cwfxaybuu
fSqrzH7z2vMNsBcm7xx0PUqxoYXVmzzjVALKzBsvhhJjMid6RRpdVtC8jCsdelS1
/IxzCVgQ/bXdvNpvFerrd8nLe9MyWi3mfuElJB92Ft6IcKe0PTYygt5HqvxIGPTJ
sqKSbvlt416utIgDhGtGsShKBu+C+qnygpsdreHrkhiiiTCZURj7bNxAJXLXKhgu
ZRm4O4nDZbbHXoBak4AkojXk0CbIS/a8ua1ppbG2Ae6SBhldM8kEei/oODua8KQm
rcLrzwGLJLL2fJp0UN5uGPzW58xKzBgctY5YAK25Sx/jkgedckTrGKDr5p7ICeR0
BO56r65Eq68deI6f1ShfsmLN1WGEK9o9zlDdScoRABIAXws++JoPNEFta03ji2Ob
BpGkMdl+jVYMKo5dGAOe7lGALRLkgICg1jEAMJOaUJjbQ0a117qBHHOOOf35NaDW
IWUL/xZyroTUO7E4WknaTr76EOJ8TNkZhfy82LymypAXA9Q9itQKN1aBCY4Es/8s
s0ZZucKVYk2q5XLOEVCnUKumFNy/bIDCM0x1IEMen3ughvJ6AhNYePIb3SkmhGTs
jtjuJ4bsZ+uLspA0+PsjCmTlt2dXL6Mak0z97LDKufKd0rNY3CmqU9kDbxXDyXyh
zmZZB5be74PrxU5SCfu0CYv+Il5EjO80pybigkSz4ZwzTKWAw4oOAfljrpWYCmet
A3is5U7q/7KUyT9r2YWcaN1uFsObMirudr0BSq5xDaiK0kFGMko6l48hTqrZaO3M
xtAmFJdBs0U60yXPVRUx7eWQo77VA4yLuo2TnnQ12aXGMSCnKWWEOwfKOna6/cEw
yWrJcj3Gx6+F1efSYhACiUjbkMZTwvFe8+IHOdtokTwxxsz9MDeLrbajGo7wzMnv
qiM/DPJUfNOw8uuYGnFCNLxPiHjOU9hVSTUOfjXTYEPkL4J3sF9qTr0vEr3RKlbQ
keazouc7/iJw81sCQxQXqOUCmiWk5ioC3i8VHjapgdSaCk3q92c2Ft8EkPjAShXZ
zBk1i/D3Iy5fpXaaFFjJI6I1yKVYWVZRws4fS1tfHtylLZjBOeyxegW+V13uNrVQ
cxaXi+kN2Kz7R855dyeZJImxl9J5ZnUwdk/gv1EiVC0JSXFQF5b/11H3bmkcr6Y1
JOUOx5MZhbjFKfOP3N+kYGgDryMnj89G/mPD0yaXo1zeeKsnMYQY/D1EXdxzTTn6
q9esjTiput4czQaJ8gQQYJyvreYDt1dHTOCQhzh8YhPDhWThsDv3cYf1o2LJxn61
6XyEEfVEuGuHuQpqtr4HDvtR5wzMWPO0/D3auV47fKsuYfdi+52O2JIY/B4qbgn8
NzKPRnvXPUtXQAaxiwCp5Q3InWvtHd3mGxhii8+hZ7v20d6UPsO1vfwvjOK/kbzp
itn/ZHYPhVeW1/aXiUgpfz3VkNxKeQxJ1Ug4ObnoMx5xSK2DwhszCHiXj1xTjEx8
HJfBbjjAJWKbJVCrkguOcV3izR18VOES3BloL2b8Ark7eEgzUcHto4vhZgZo5jdd
OqbXSr5ZlnFmm0WrnUKWrrXK8A1GUTKOpQXZRlwl+1A5Zwvyo+aPVcwT1u42epGs
H7MQN0CP0vZNC+9MF4S0qCZ+0+p94Y0+go0syD01GYPOHtqQSX7m/sW/oMwguQXb
DMelQrJDxw2LrkXJHKkCW8LF2pEjcrMw8/NlECeRxk4IXwKAX3KghIj6dRCURDcM
lZGF3VDjfYTV7WrcoFIohRQv0aapB8xVV+jT4OXkkJGkN2SaVeDiIMDgqSfnIaPe
EJ2D7Yk3lyHs45sPr9d+7uio8wdjpXmHyOEFBTSPEWA2+q/e5ZfOnUTyw762BZsa
q1+po1+BmE8pYab1BxZpvsfmY6wkDNB7/03MRTaPC323IO+6HoSa2YNQaFQD6q1c
G6h/pADLkOlSorYhyOrLr3TtWe6JYlWtzafZb4lVLL5YymwC0+qyf0Yk7Msjvc9V
u0NwjFqsmUPRYK2xRP0ggnv+6d00rW+OlhqipmIMEqDwex0+tK95UcUGophf3fjJ
diL6vc5aubnjqx5Ki6FhdCRrR4jsz9eXZDj0IXKovj29nFrrX57vF+f8V3TLxZAF
+OzV1Tlh5ixDMlh/l4PjH49qhlGmuOpnc25LgJbbOg6e/b5aNdBSiINN/khKVsP5
7xzKqXL+jTGs7GdVKOarQoGTZDAlIHna7zW7jSS8wX2DskVk7ahHqRI5Mi+fzQYz
s27yNdWLSHyzs2tf2IjV+N1lAT2tkaBBGuVVzj/I6Uy4MTglbIzYFls4lOWEDcWb
/XFGV+wPhLe03a3CN9tJnHv77sxbl5N7zycYRuaBigYsAw4S+lPh9NmnXAE3oiKD
d92u2aVf+HUgMB4NM0hU4NRfwhpJWf3nDEqS0HxQpSrQuWPBv8HtHCAQnQrwur4p
2WnlW6AyK1Bi47GjW+Wp/szp4mY6l8XjIT9Z3amaBkpajoz5eI+dfg54AdUZIV5v
Kg5ZvIqMBOD1vIf0rXQ8kmLBeLGbJ043KBvvLsELrqPSKDZxEL6f+ntXlodYyb0y
vyBHzjMm3lrQt4H9yqFTVF8Z57mKGxFek4mwwfkXrHwI6x7EVG4qNJYPcvHQUgmr
GGN17GPfQjV4OAZ5oBEsYTmMEARhN/QRglmjhcOCLMVmp+TfQnJA+PbJIbFhlvjM
s+JauChK5aWCjUhMnATtmYroDEs31iKwraSiAjW0zCX4StA7FOvUVRF2Vv3p4y0I
hxWiliSep9FHYHM7RiMVF0wYVPHS6ThQMQ8AqqAA0v+n1G+T9qou1SBQN7v8ilWY
I46oHc9tKUZLrJP0DTDHySEFrkI9PzI61nn9S4z2Cp3t3sd5IwADOgh9+wjUDiV5
kv81iQznZN69DXk2UPxQeQBuKzTa5q2BtCX+m5Q308FV3LyzEI6gESHtKtBYjgx+
TqwTq4jt6PBwxdPvkFEnGk7IiWatY6vrUCIdHBQlXSfbbTgBwMhOZmyV9fdnd1pF
ewsDC49rhzSpdFGZFy/2Q3AqM/1x4gFoxdnt5724NndUx59d6RPPOn0/98Bx9G/t
LUQi0CfzLKPpFdIf0ena0YWEBPCUN9tHVtkpxqkGUMDA9QNRYf8GhHZwJJOYeC8K
As8iUmsr/8IKPrAy+lwWjPBs0P82FdnOlEeC+OiBjYhpNYAwvSJobLpCSD6kFIh1
vmgXVAk//NLh1ntoBRJ0HqKYu4FECtdYKURoEgrXSIDXG2DglxpGiAahS71iubcX
hBQ/j9iWoZ8/cnxkqsExQKLTAg9o4NmaZ4YnwawTcezmqKUkag0lufvNyFq6zhN9
MNW1cTZYhDNOx8aUnOcdSI0wpqhAX9eXwsf8QmzIc1OPNuR9+2yFB4VYLcMPk7Vj
oK7Zr1H4+TYQmoA4fNdcM5NH2Efg40PlDO25dCjXdPcyaZyBtxGM6GSc+4rP/Nef
BPf2FC5X1RWTRTDYXXV4a/mbtoNjoVrdi9nvmIlJdSboPsRBmnZOGkmxndW1jp6t
YarGKtdPYkPqmhPGNxNmDRRstBY7Q4s+Tmxd9KQgGAZ/iNWY3QnNS0VQIzMUBq59
eTAvhzyzYsCz51gkzVaGUnDnMfldp+ANIZDPMPqx5K6iAttcDUY0/f/XquuuFOxQ
XJQkNIQWUs84eEX4V9tJB2X8w3gpaOE1LvuL4imbDUGgct8v/vL5rMNymJBjoKhQ
x3X09ExKjHgfrBN3isCMBXO0i7/0CIZLTZAa0bGrPKoaRG02Yt5bHZ7BWSHe76cd
YS45mfK8srFwW5m0/2cQ57UUneOnZcPVOnfS5zJDXVVFeLyaowq8Ko/XIPYvoVo3
6UqjHgvc1NoDR7WkwllHQczfoCocRgX64Nnjd32xDBmE+2bdYmARJ1q1PwOPOgPQ
xDaCON+xEjdC7nZtTd1gzmjSwa6yhbV1JcWLHZ7+M6ubVQqI8fSVrwHdzPBuoN4j
iUToiUWHb6q5KF8mB0oKx4Xghy1fJgZ0xO1KvfZlINpWoo+YS5+1D/r6XzF2w9VL
NpdYzcdxlq6xRcGM3/bAoO6GP68IWe2+oQV9CtW7IeCiihusNRXVeecakFOU0976
0TQcxJ1EYG5GMmUvMIPXjRLa7FgLgyTkuZYop821YkhGdiIAFBmfh1vuP/V3aD5l
ta7BzWZpU0G7K7TwuqBiGI7amTSwjzxBfptcmkNaWoJUX1uwA/lQjUW8dsa7ocvt
v/fTe+/jYz44gV+h/QY6IpYDqzO1qJDz58pvI6Hj+Up9gIpVrJP28odTD98Y8+Ok
ZNbdkl+5B7LT91fO+YCf92RFc1Hjg7zaY6snOZBqh65VJRECtzH17VJxLYhArFZh
hEoZmseBxd2DIUXjAPSfFgdLnR3AZJwgc37faXf1jQAWOo5Kdrm64utM+e5MyAtF
+Lz0Jox434iWDuGcW1FMtgL7P3x41qINzs3CQUx+pCACzDwTs/YFHjwGsDBu/S7X
uljHDqSBMCLxXtLXal8oWPTGO6sMmtXtDXXypdlxDyygDWF3g1cJ4bCda24TM1TQ
9zeZlzl5CY3DodwDE3NGDXQb0cvXkGFdU9JIy5Cg7r9YVkxIYji6Bl141hjytUv2
1yilaBZDVUEDmLOkNEalObPjg2Uje76dpJmx5kXrtmS/rTpM3uFiqfAQi7Gav6Ls
jZOAPv98dq232Ol3flq/3j2MlGSDDQv8pLqZwNTYXmevS+RyPfZTWVp40NJwbRfF
nIIFTvgcqwGRP6diW+mv8G3g3xG7UDEHrw5E3q9hegd4wVFzW4nHR1/t0Ee0h5XS
R75mfqUFLCAumYnz2uxd/lj1Kcu1iQyiPKPRvW1RumgPjFAGpolEoES4EvWkYkj1
ghnsZxspxk6SUuzMUpoeM1cl2oSgq5dnZ8wNEYd0cgV4KCtdgDO5KKHJB2NqYmqa
MacufmPnzzzIpoG4F4jl+IAE55UaUbe9JqXQFm/No1kSq25FR8OLKA7/3xrmcs1D
QiEdQEs1DDJpAI7kA91C09Ltbfv2SBI4oNzVlggRVUFIvvJzrK2ZlgqD4vLN39Ni
w/oZplUxeg+FGkf07VNy6Vx+doLSRx72824Pjxahv05GaZTZORvF0qrnBTg/vYMk
+R1ZscFU98upoaXW3gkPf0IvP2BRP3iuxkthP0DWkyR7Z51ntC7WB/zwZhh7gxUs
L7MRALmIlEPSE7pcqpauxOvtxymQm9lijEP2Du2V56PQR7+JnJLQ3YhSBxfAmyg8
1VFmUaq2f5ncSnwsTwyyfvDOkY0V/qcdy+2wOtRUd430Z2SjNF5Jt8e4ikV1tWRA
vsZLBvHIkROi3mAQjbK+6S0K1z4eDIpZUEGbJQmHAaNR7oe5fVHBWzNKvKJeV+q8
emP40mrYcKDeHd4svIG4swCAI86sfje+3XCrC1Wig37Xcc75F7QX6eXU0sxWpJou
EI7Bb4vWuhiNtfvhxOmT57CFeb0QrbZvlAwANh/KojmrJ3gk+NqJ8t7D7Nho5vBP
A/ekqcBEJup3ftoiQNb6bnZnNRM/5hEeOzfJqUQJs7mGO6cIAgZKZALNzqwI/gxu
MCE8JLpNIP/ruhWgalB//A8qgQO1BK7I9lhFYYpHAQmNao3FZtwtr+aXveq7rF4X
w2cG8lwIrlJ5DBSfy+lqbcKwqwTdVPORowPjEYuC99zsEXj8utRvJLe9Cp/RNZm/
cDp1l61xZjorIwUkfCR7Z61jF6HxTXQar/w3/ph+DQJq4f6O6BXgxdSx88XQxhbX
0kEAt3dKxotW/MF2FDl3pSCzNvI5f409ueGAvJO6M6V220MIW8MRIcMhFeSzeQ4M
chYM7gWNp8dm88ej+fL0gldJw136QnI3ZU/ynm7Ihr8/HL25fdxECFwGVOVKu6SK
8Mo98nZTKh5rAS6Lcyn71c2Wbiq0KF1qCP9/KVrl5M58Zn5Wn2JWVgFhm0ZPM6Bq
nPQN8wTpf3gbdhjmnm3TmWt5enppVBl+cXMCvnniBVv1MZm+mO66gNfdVlgh91zk
iw3otKyUVZE2I4RRzskIFDOAOhibk5n6dXfx6QM55mKiFdDmoOj6x1mX4/NX3xhs
IHmLh0GnE8eyKVZSp2oWuU5WCXQYh6dUeKsUKtPzwGncEwMWDjq0H49G+7x+2Rov
H/JAX/hNqs1NubumZjUoPaZ3KDj+g9pyBrOmLMrYwWr/QTqmL0I13BdDRQLAVFz7
VWsNwHWMZ1G8LAVtwPofPJ03Pzr1b8WBPFYDM20ty4OpuVzy3XDCd9bdUdQKOcwk
rScYde3DHSTo64+71+UjlSEqW+yf79IlpwY2TxoONVCQNfX3+3jtxRbBQvPerSbs
MqhG6aV71+iqoMhPBJ777gwwSheFm9F1rf9ebUTtzoIiv4Fv+Gv0dErxCZF2vaRQ
KOy9DHpEpody2wRjt09DlqUjwC4kBECD07Ab2p9VYT4OmJj1ON0xv6r6lDFWhgkl
siOTg9Ltgahsw0xuajKvlmCUlaxYIliZpp96ErM8lof9pGMiTdpaU32QwztVNzMU
Be+FqPfaMKiQNwsQAqKVs0DkE8K+zfQ1jINmkKNRLVTUczYaEN2l5TKyDVIFHqSe
Q0OgLvAgLgOjd/0kXWV0dy5i/UgRWms/QvOowUIOGtJyyQqYbiG/IcGJq4z5g5OO
89ZXBHHq7vSVQQ27+iKlYH95ytDpqV9AaCN3wPNMCo+bjjryfWhz4yPIZoOm90iK
y3lhCTEjZKUKQSgImBJ09adGWla5eBltsJOOL0vzaHHz+h65C3fdGeeW0w1vICNs
ruZudEYl2oxWDEy8tvB9OzMydRHaCbuTvUNjB5Vmy/n5rnBrSCaxJlgUBTBkngH8
oWCLI5nA3NDgAcKthxhMyZkz0V2qSq3t/nPwTcbHLxMee/vXAfDJ+keLBM/voLie
LvKQeyt51CJeJS33+jg4MQhLQ/n8Y+c/VjZuvp6wO2SxGUejZBC3HQh1kuOpKsWo
5p67brWGTXOmvk3DVwRnbyjy26SHO2wQnRgZ4jB8aq9wpJYIvXkP3dRComOXKbkt
18JV7ZBP3PbnU9WiCTesuEZpiQsP+87vqqpB7LNF2wbxJrq2/BHnLB5z7f03RXCc
mZ9Fcv/Wvpz2c37dgPH0lo/8Ir1WdzFDQBeEdI2XW4fdM+g/6UYyVf+VUw/fgsS5
Zd6LEmFTjhVF8kYEie8N0SdjFnthvrgI8RmlAP20gXYf+4Wvb+ZDJZHvJWPJx1Me
zE8r0JKcSTxfi4AMbdZNyy+UfgAnIqtuYpe+89JTwlexKVZvElrzINSKS7lSApzo
TvzVEJzU1pVDqQqJlFjVTDP0T88cG0rN6toa+mILfqaeDANzG9yXNwQQtbyUrcsM
Q9xarqVAERUcischPBlt1MoYLB0bv0jPBm7XmLKVTpz/DrGfeY8T+8g6Zzen0108
L8VJv0phWF7D9i/FbqqrGZ5n+Pt2WiUQ2uz5fb0D/y4i7IoJulmPtO5tKgykoVR7
Df4iaA0uWkysYli9pVXEdlobxjU+latmwFGZ4EtAKD7mSsZRUGjtGvcGgIV61jGG
LicgqQdOYSHN76gJH3CiIS5pje1+YoMCcrXtj92xt1iu6Xm4kMvdSJ+UrZa+31VI
+2UESL5p3088cxfjn6MZgxF9DELUEWe30sTDmkTAlm2TXl5TazQqStGZJh17B1IQ
aPn9Jw/KbXntEHz4HM059n+uKB75f5avQXEeRwPzm9IjE97B4oI5jl3ex8qdyKjK
TI11Z/06QZHql+WFpNRipTXYf0QV8ZVZofhQKzFdkvII7yI8FGOTF8nWkDY9wO7T
O9RiIgfwKvsV6U3Af0FH6RGS02y2FgsxmV6UzQeMFzZayDBQ7RX5L0EsUtV3QBvY
J3n0tRvy18Yc0gE3Fv0xLJU90Ng+ssiubk4EAXfZYT/H4tSPyDf9p0UgyR9ZdF67
hB6Pt6sNBD7g3eBVxPTda3PTRS9wNrix36spxLOgECPWch0MNRrHFSWZQ+GyGXqc
OS8B0hEJFdjXRtD/hb+CPz0AcQnxENPQTTTYodhHAd9Qgx2TL9rSJ2EUTqxlT6Va
p3RObIhfA4R+ZQUk279vFYpBDG14xO7lnUEdC2qgyV0iUOoGpZP/4TEdYPYNTKUV
qaS2Hbzj9U/Su3mimfox/PqAyICDISzsNFrgTEzhtxv74SiR3yitKCrrXbDeAlWf
AtvN4xRvYpuuPPEHxoI7ac+3dyNWYyo+oWRkL5CFDWCQ9Y+GjuO6FKn2MJAmk95l
+EqjnTOomT6QdjCt6RkR546OK6c0HCLrHry1b4a30U6JdNY6lEciqBUfjLnGBQjn
9AVQsoXUWAy90p72QeGrVoaxJXWoLyVfUBnf5+y8thHvocMGb2GAf2yE+QlWIz6o
N1ndkVDbphjatr4VYfpp5ZfG9SGb6uJp3Vl8C/8buGzLXTDqaA2gezp3THe4/yt+
4MrmSe8ou+P+EbXDDWi4ELNWDM7L+PbAoXTa+JVIcP8Cp6bnfbftFdonB4i6OH9x
OTpO/5dhgnW+5sWGEmR+bXGwESQYsrAI0uP9Ff2sddfGbyjAXDMPDwhyEuRw11rZ
+Frv9n9k5uJc9n4yhh9R/d44zjOqKW0zWgD923yl/9lyguX/JH+mJUqzoUv+9fPK
bA1GBEoirKBZlwwNEWCH3Aajk5l6jKowqplyhvDiUlPC85331ZPlrao9tOC5oUHC
jjiWsdmTr7Sp4hpkySE59cOZapCoeWjPFckl3S6HkbyFpvVLFC5SdDhpeMm5jeii
+Wm6lpS+PYzLm1zvD9liOOyHMi0SZyGP+fB/u3TZZ64o6ebvjLkAh2EOmaXI+lG9
quKSJMVUV47VSl3sMCvkoR+F07VIlPyBi1Pem9JMTmAZPKaTsMcrhHE1uKxBWNER
PDpIpjvnGwQ7v7c5ZHWMCdC5oqapBt1msuQN8RiDc+RYE2/PYyddP+f7aOJS9Pc7
7eLb+bTTXRtS8A+ejw2IEO+t7Ttgkcu6/Kt89MyWwQhAaM1TgyCTO/kpxGWbwkdY
oTtA6l0l3nXWy/cpUl+KvGdr1z81IObB+o8Z8QrkgjKJ9Jt0nUS0NIIyQxGIDkqK
OrXTTy39q25s1tMHgRx5oPTWRUem6ylKMnH41NLUCz/zrjGOmGXssEwKJRuFXkbg
Qj8JZvefKgPpf+httDthRXsedQkyD86gvui6AzwCXzY4I6zF/mqDZudH/5aAXQUZ
0fo6VNc3Ntdz93VrbGRYbsjGrOR7idwHJg8QB2xGa352UjJJVp5glEaOm8XR7tpv
w2PyCsBTpfQpobSgS1Tnr9F9MT9jUSK+792obTtKXhfx12PeB3WsdpKyzShmn5BV
XosQkheTWzJbHSL8G01BtWc9BCQHgta4DXABPweguneJDLQTPBzB8zjp8ctRdIhq
ZU0/VvyP/25NLkf1UL7IP6NUVWfx52Srd/DdqPnCTAMLhvyROdt1jrfIqa7CFl5E
ZsLiArNDxp2rAnAJ6PjoLi0YFrIhpPfLqKvKfW8P3Li5d/vuwxraS1/CmLI3ZLlP
e/p+abx9jXO0PmzYwmGePmsGnI9jwPw60v0JxvQ65x40/rJ26nJwSczS0A/N7y4o
DdTE0eAqXdF72eWaRX03CWNWalDTLvH7kxZHiWk+ErxjaWzDJOXnbaaPjnnt5kiJ
IZbCPEPV/wjx/fY4plGNOsYwjsthfk+YERBxCyvuY3JMUhFPCkrUN/Fx/1dJYbOb
N34AH39qSbirKm823clot4dtYatiKgNpiJe7RB3wuHCfW+jwsCEStR+qi7NwE2CY
6wYgxk2otx4iG5NJkzy1YuE4O+nt0BD3cLdN3SrWmGrmi02S8mM2DpwBSjky0QUx
hdPmfXKegJ2j5IzBITOfFspLUMmDXL0MUPH66xbT01Onf45W+B31j+PVMx33d34l
6JuF+EunmBX2UEMSIs08HKJAy08gggtZZzs3pUEG/mf/2KSxv/rHE+N4po+ufPgY
tSVGIqZTPwhBu3gtSJVw6m4AvEFzStNDkLtuMiiDv+7nbpWaRTkDEdJTFgd1oqWB
qCsCyV45mAonYeh8q4J7ci7V5hTqQTnR3cVfp1ZY2+P79IK0JwOBRvONHthkxGw4
Oz8pkI6hyznlk/mBLet1prts9mdUbzm4m8oIKPPorFtjXZbODtO3mTRG1071tvau
Rb0lz617/rq1zZ9IHDDGvFpUNLqPT6KySEb5C4+Sur8p9Lvb6+adjs8/JoBXYON5
EcDz8F/FFJy0OM1bf8LIYiotAw5GyJ6cDU91zGMmPoh5HGLRs17HoTDPrODQqxwD
NXzcjiqV4WqCivzjuvLHnvY3iGGs/z3wMykwnxZNRI7aknd6E1dQe2lZ0csBncr5
jLXeBXFuqB0Zcs6+Mwn0hIk9N34SO8io+ECWg6i19ZCQyo6feljKU1Ah3YmSqwrO
OSM3loo1yNNZwlW/QUBQh0foa4y4KaapvXxB11U4jT3sPm3se1vmEFGIQJsJeoem
NESNkXqit6Jm4Gik5zjXybtMpQgzrq4Dp4h5nFXfDI+uoDEDAsUbvpGV9FHQYB6E
ds5QYvUl7bVyNDYyXZQ+S1mZUt07f9lCOIDCKyxTAfPcs35IgABhrP+A4rSto0iM
4TX0deVEXaBvTUIAW8mDEqOZGcx7gTZsivcr1erIsk/gC6xUhusvUrTCNobk4rQQ
u/8hIHU7rFGNtsh/8m4G3iQcpJZtHXsmKKaEHrdg4hvykEPHk0/WTg2HoGrC32MN
A+9RE3aqXyC9NuqeJHbklAV1wCek0BoupsyYI/pCMYzyvx3O+SaX+zK5Q17JVpVD
tpBsPfyuhEXjIQVivQ99ziemyjshJyjN6lJ7a51gcXdmpdzssJG6slS0B3PBC7Hh
mSckstkDGG0f3carf8AIFpWXYDXD5vggNFVXSE8/kEvqpWG3qjbGC49EIBZUcq3P
pLr0GPFbNHYHn64PfnbAaHG1619D8eZ6fFCbcDKh5jxiB5M0oQfXLFai3KJMj91L
kMmelJ4vxpSe14spREPhFZMx6IzqPTm+AitJ0REM/j544fIVNa8c2t2YA3M/+4zw
tKTvP7+Hyo4Jedt+pg9aM16CmB/hWuWxcbHVWxwDALwzK/pu5JaygkeKBOTsaxj9
sxJi/iifz4mekPOLeuVrtDnOs5fmlzEzj9XOoz2L1thZcKqcjGTUeLpabWSYeeIs
41wP085do463lPMuG5zArIJ9aAa62rzOt/AqsEpRK7a+3URvN/LgyEwJgk9IC6ve
Gc9Z6iJCe+JTtl4mYxTEqW93Fjj1N4Gn4JLL5ktru8+/B0rtkwFgyl77mCweaPBs
8peXiQPuCRPqasi9xDY8NiEVLgrmprbGOTYc8EUE4zvR3kZaCUfFCL05n0MiuSOw
RjeXv16Zssc0vRgiTV19v+w+qToREKtXjr5wUIqhcWe/+InE7RpGPWQmttiBWThL
UjVUBMW0rejtkpbvZos8tRV6GiHaN224VQR+LO0BRQHihxmNjMks1FFWuu+TYgNp
Q0U/vUG2CFUycfNttWELw2S0FkuJe+eoPfzRWfKuTcCNsE1bYWPTkA51lpRkxgfm
IPeAvbD6GPEL3stUf3eGqG5BbdSzs4GXQ4i211nKiTm2YqR1RL2lYUNeJ/mfFAYu
vTakXcJ4OxggvwjQFfm2tG23dhPaFZl0onbqaVb1YzCS4PtKPcowfgzOYAGJeGsG
+0nSwPQbqjeZviyQVcFipHs7WPU6gEZhF0x9ewebkUTyF1FKTbboK2N0cviSZg1E
MVvOwP7hlMW/d/kkPi+EHi/fP1CV/r4UX41GzhA3x0/xqZef7KxCa8GvWfYjeURO
nkUoovACsXX+z8uCz5OgxUgY2kornzwJ39bJI3d512m93KledzXLiJIDyjwWq+3v
Y7vjK/8fAlXXXxrEvYdqkTFiVVSQLFnLbeKUEa4qzHhDwRj4PIUNyIpobbUSwSl3
aeXw8KRw7L5qyuL5WJZ+iRrn58HtFRxRYh0YWMF4MPSLg5CxuqGRConOQwScI89O
mA7xqqi1eqyz6aScBW+nQ8qk0IGIb72lK43kb8uC6zQC4RYThkNsftLQ9rFSfAu4
tobGbitn/dvmKdstyL300dcDSSj8zSrrGcRZd1Avlgx9iglDWKcz4vJDjyoeOP6E
0M32okbmPW6h9BnB5od6cKNcN8DFJzRzfmW0astfMoJVk64hOK6Z2AhRCnGJH3kw
cPTsprXCSEYqufOyipFAylS2MWXc2Emx9e7YFmwFaHGwPpCok2y3bID+cVQqFeCG
repeKY5yIqWArfegD5EcfAEwyRMlDxbwGJd9sCCQpejHVOB+FmDYR3vFXumwFlMp
IiPchyBXWHt2RAYYP0L7lY/mINp7bZfo/uHdU84J83pVgQ50C1l2YErSvY9CceDj
vPGCB0jCzjkGQLtlisBmtJwIdwXGFwQTJ/5rE0OFVy/NKN4YJ0tQRXFokUD/vslu
M2IjwhEb4Z0eoccsN66yRHI3FA+7siFE5r/vUXkFG4/rHk+eGYxwbqQt6QliG9Z5
kKBMIVDDrz41Ds8hrQecC8XUQeVogOWKs9NzuhJmLhT1RcMLOVIpezwlpLPaThW8
QYG3LhH2Ganj/DVJLEC4zxRnvwa6nJPza7aDWeqlWNQ+JWIWpM7XxYVmPklDTvcp
ULBlfqP+QlwKQ+Aa3qgoynFTW3jQ2TvIjYauj8g5nNN4e/tGcu21FbaKQuLRmmc6
CzxCQahGCfRNI9XjJjwMZMCAwRoTmApG15+6Ji38nYtOgSprh/+wj9Asb/GmzmAr
42z+65fWzNOpyJz6S5+zqlE8VulEI+OFSHiOv2RkfsS0UJeBBy4fXcLApqtUhxLw
e8GuhXWpaI+k1mkxzGMJJMHrZhysD1FLPcrhjMJJIgah+WDZnWPDN7FisM+WTmbO
vWa565IwflA++4LNnU4/HiadnCoaph2CA9fo+2J2LHZllIJanzxhOB7ZBvTgbPS5
aOL9gmeNSX3GyXb7dLYCrXhzudbBfZ3kmi8/Ysts7CiOp7rBXjF6urDzMvFebDmW
/1uwD4xu8+KVG7bW1ZB2GEcD7r3SCZ7TTL18BuN4BQ4zfcheV6NRm23wQq2MeBFh
EhBFlMrmPGSbHNYki288g4wJMGP9t4ZTvumGKRg108duVduys5zqdZSv4LojRDfW
voIM9TWXPgtE70u4VNUcRP5/FE6l3UFmufzMA9S+sJw1P6RIg/K/9phsHDT/g4tg
P7Io56wR/WJ5g9XzyGZO0QhboTocPhiEFwamC7EP1tBws7rf1fh/pqCRoK48yg8I
0Saa2w4g3t2XY4vEHRxLki7wunn1mu//JJ02OrrFRDILCfykgIjhMBXXXWrnG9uq
uNU5FQ+4YaWrzOLulVcuB05vkgjAhi6HCrl9Tyu6IYfCG7OTc731y7UNNQGxS0Jz
ioRz1RcXWrB4PoJVwHYkUp2lpEZ0SNzft0ev+wLD50RANulnZ6t1phoC96W4h2Ch
izUF6VLp+2QklFRNEw/KEnY/m6eVfGy3WqlGPjMhwjFYJJLpVqAFB6CD0Vbfo6Pt
DbqQfcSjStg3ndu0H8Ve/0do8htYtK7gmHmMfFIdxTDqHlmGh3IfThd9CL8EQ+F/
6sERP4jczEILwKs4yvfmUJ+zkp3oatuUVmae9C29KJAuJ9P0Q+yX/gHTSHS64PxK
W7FG2VZbqdF3XtV4GFEyc9QbpTE6Pq+mrmRZjErvbGaJWxVlGoiuZ9NTuaHAcinl
XcbUkcRhu5BkchjWsZk+LINMMFrT7Qola2sXxRACRfSoIKhgG5dLsTPBRBOTvhE1
9Q7qtbhrkaKtzCdCl8nqE3s364BGbL0cq6Nj+iptTuHqEHjqMuv6zXvqG+VdsrDJ
TX24q//h0UbnVAQvbQvtiGmASov+ksmAwMQxzACep1K/FSydxA8baq0DgmTDo+rD
smOaHA7Dd86JteGNmHNDi/eBpO35Hczjn8Y8a9+F1KlJC4mejQTAKBz3cUgSJpCL
Qzb/dXgUzhoGc8NEWQWxZl4zqcWUeg+j+0MGxTFCN7DByn78QSV09lSBskD0vQor
QhlR0Fb2p/l95N8Uc0oSwRbn+b/lipElFsnjKZtEahMBKNuSD8LIaZwHbcR0WvTv
ukYPeeXt2qEUtj7H36eEnWJ9f903V/264PmK6qCq1gl+h3GFGy+2HrxIFOgQoC6d
4qxfqaCdaprWPOy7WWMtQfZ352U3QXEhfAvAAaAb74oioUpbSdJkA2j/yzmzZYHW
XIlAkM1daqTxYbD9IH/s7cKIGV5TSusSrbQ+MbcK9n6Odg90t85fEhCt/ne/Jj78
H0LUAjyrhh/AP2JNix7y/LNX/QFd1x/F+4Xp/yMYRIWbh8TnmBuTcw/92MebWDIm
k8QIE/zTpbEu+QHHy+njK4F80Uz12feh7PPvKfcUkwAt+ZvW8frdhJU3W9xtb/TK
e6RD3VNbjYcuf9U6ietj5UnB5bSfUYRPVJCsno0W7SeQITgddyu+8oZhr/trAwIm
sy6q9jcrXMbUMdyHRzUeW3cAvoZRPJ135dQlWDQocFRFAOAy4dCd2Opr7hc3GeK2
8dRIawXBVxuRICQcs9FtRs/K+q6tB3fG7h040pC0Zcj81uGjUC4aAM35LYnr2UNW
ZladBlty650eB5NPW8bmp+RQvEvX3tnBWdiLfOHxlzjvNJBftGCdZTpoUAPJr0Nm
YlZhbrBhA6y9H9oEfCMVK+bjboYfv+zbizfCPzWfjN+uMYcO3fnAvpvJvzG4lUPj
cZM8BbQP/xqHiaap1zijVUh9dbbPHcNfSiFMBmGu7twskTPCOXE8LuCVBWTE9VWR
Pa+Bs9iARTeSUjbIWR7iCo+1ZHwLFg80ht30t5ysFrY+13YLB3YYpgMbN6V24InW
cl3PaQnrw29CV5BofXTYTOkwuxiaW6pgf6zjHmUuXcxNZpp49CgPx+to0/mDa0SH
Sq5byogNJkYfA0Js0UfFf2xmSAg3/Y1BfT599C/cwVKY6aW4n+8E+iL+7bJw7vLM
TcnEjKPgeu3hztF6R0amTmPotsZkGurObZe6xgQiqYzMiEMg6SsVze8skrAYzLod
OZMThHNrzyotEgZnT0hAROh9QTjH5t9zrC39BjF6OWotcqpSKkVR4y8ZqGXt3SQw
i1RftVpUirVvLFx0eQaD72s+XgEBqc5uP3oCk7thRiRKks3c9EA2yaxSwLn9qVUy
KAlAKeW5XUXdYIHEdmSkzlSQwRGl7YCkCIfNgCsnINE67e1waZ6kYCGZ/qinrcwh
o9D62r4BvzWJ1w/KtuKWgPqB+/39ELIV/4LSgiyqh7FLf5mbvHpXt4cTsiF3/I5R
wU/U3D4xQQYOILjqQ07o1/vD7JtupQYGZjj/Dre5SlB5kPs2uJ10g31ltnY4vQQI
KK8ub0asBFZ+EiwKC95UjLaMRY/KfdpUbPq6MJlzkXhcGDo67V0Cw5jp+qdJR94q
3O1rOCHoYle8Taz91cyOSmAzcyIYpG8El6b4Ay3RKcJ7lGyLFNyJkBmqzEFp0jeL
C+uW7TkZFW0JkbsOanI+XytdYF56kV1pVecn2i29QsJUWIkKeuvQTOstYmwrrTuB
OTvHY31es8yr79Bo/lDcNwjhFNRw1gvEHdVEML1Iq2OeKMIKRMayoKUM5ZMCanf4
N98763XGGXCmajiaCnrA5ilTq5g5ONzILeL+UyVYsKl76WPDpu+sYJroicbt7POG
eTXqqj8SWMMRNJUtEa7D99PsfxZEca31n5VPo+zMxPRyJlnAlNcQ2kZCHlsW4nXJ
jW+VM0BZYcTYMmXqHLrvR3opzwODwjZBkENadhOWl1LcntOR1nbM34U1QvSXi+tZ
R0lfFHVurXJS91l2yBGY97iXhFzy02Jn1Ydl6OzpEHtLnxaKKswmZ3SfYYixcUX5
XBuuuEXMzFXXNLnngmKKwq46X5A85LhewyK36fNflwpwFsFvVjIKISasDFfxZ7Wv
Wy/DwVpcYngriUijFJtifs01BbcH2nBaqs4unTjijpwIEogQmLKrvqk0vVbQ24kT
RwkO2u65zk44kuB1lMIeRIvRGJf+IFzTgY968xXCI1F8e5my1Cd4mkaqpBT5zfiC
+4yNFcAEiPvAL7g9GjQBGu97TpSQIEEDQIKzgtMFVCI5qP8NXtnFhmB+v5hyMJJV
xajbhg2X/d2LtBpRCWDsUrgXfn2ElfwJU6W0QbC0emgCK5eHpPKPfh34eW9CkMdq
eCjXS+bvXWJ5wpIGoxv65j1cO7czqE5FdKUeCDeNeAwoD/8Swa7U76Sm9GzdJnFJ
Vx5GLEkG02CH3uwF5wyrR7sFqqzzLaSFjFyFSouQ8zkWcqIZk1J451kmeSG0OGLf
MkicI44Z+fNKqUbPO1JdofE4iViTF2MkoAvwimRGagjSVFruQ7WeJLvV71a3Y/h4
br+pAw0W6ET0FEkzaO/KTLodFHHVZMZB2+YZqlQB6Te8m7jHXJ5b2+36EQyhmb0Q
5r2+434j7ssVryuWDuGWRIRHtOUddhPDvk6fCRV7Mj/D2JOohg7Talnog5A+JCZl
jYZRaBbCS4br1EMZfWBGhhh93GqmP7kQpzBB5CGNKbec5N2XXZFxOKCoei0L5gTK
d4DbosgPHzNvbjj2mtdqlmDnRu7njzoQe99zU4SkfrU8HGXBazOfU4AovYEH1cEN
e4tMl80i4nzP6wUiLzKVelSNqn0uqaX+oKhTcPaFit8vl5wfUPEpLKjmaAiGiTJt
peWiqMg4gERgq5M/HxjTvIOfBDF32Gjr7wrkC73kZwHZGUPJ8qRtRvJmzgWHsz2Y
//8H3pongUEahBc4L0RD4boKQroKkZCaUEmrIj1IQ/rucxd7kBv2WYx8yfBT9Zke
Wx3Gzc6XtlOiRZb2gLa/da1CxlrmbfBfgRHJHmvZde83hWLaKUVlsojl7Dg9ekll
NirTGjxO6xilUhzGTO17WNw9DILbNO9YjpCA2oc2aQvIG5Q7R/SY40z9kIF5EBGP
Ocubnyy/nxkh/YPDWodYgxe1BKAwmDOkk3ppTZpgHyxAUsz7LZoywxDCuChZIrcr
AkxcI/wIWioDF4SBiVpDBxGt8Rkw9olFmNkj47Kx/S8yH0ZSvYZ2Qnf7D+a9etKr
13OygDaPIlqQIkohk8h+5klmhmPom5W6ZDaZvrpLjohlKQlYELhSocCZ1xlJ4AOn
ciscrHOc7EMOIPl/0PhWEO05SpUxT33KDE95UEqVSFFM62QGsSnZIGB37yZG/a3z
x+m5zwf0a7MF0qrlYdNR0hqEMgptdwOcGnRkkL8lhlQTKnR/RczIrIHAM//LDtWZ
lWji0tVno3uXX7LgQe8p6t4WKybvLAdyakLCiU/CmWi18lMRxRPCWGo4ZzzeQCJA
mpRu8SNQAFl9/9MRtSFCWsuIreaNBWzK78NwNZAnpn/mVinNp4tO444eSxGOHUeP
LhQgouhjTnIp4u2k8Vrx7h2LHBKX5tROpDB7/Rt/3JRXIxjS0yZw3MOqedJIeYEb
Wi2morwgA/QJW23Zv1yCbErEiqhN2nbKDMSWXjliiId+7bzXUcn7oeFkRK3tAFU2
nCFKYeap5HVKD7zbUqBPZSxlRatzIkUWgl7M5gWcB6aVFOYrHNFoWQT2qVY18QA+
2j7Z+UFk76E5J/DWTR1EHkCTipo6ULYhw/FdIORFyCX17WpfMRmdcNLC9sMKnj23
B38RttnQNaf38OuSqs2IME135wRR/7m1Izh3i0TZD68OPB59/9O5G9nrJ2awS8QN
NI9/dUTElDnskx28TQwQsETyhVTOrI9B3USWvsf/Mu8LCjLsmgirg0mxr7rKWfHZ
0EaBVLo8d9VY8jJZZTlTnJGrduv4fiNnZ/1lWZULrWQNIzSU49iWrkOPmK1wCoJG
cdhHGKs5PjAdgpan0HnDUvVLF3HNnYtVfaRSnjNwniwJJuzHIWgLHWWOCquJ9DZP
2VXpIoH8UgMa2Q86CALOWGa/mHqN/ffdV8O5hlOubEqhgeA8eoq2oKqgdeqCO1uw
70dW37A5FNaWtzyodXlMlcnSrFJuXyBPpfWWueEHLk5PIqhxRY2nb6EUbctNzlZB
B3uft5CaVIjRl3f1NRfRL7oVqlO4itPoVzysnmcBlS2yErJCVdIzh5CbxuV0fFWL
q0J9B0h2YpM0coZK4VLan4UscPcY3u08x9tWHMYWfulp9R4pzz1Q88N1cTiR2SPb
G/KG9Di+WC/spaX8RkbtMuY11gT5iTMA2R7RrrBQgWKRSnyQMpGJAuNx7/43q31/
OOdQ6Cn6ORJvJ0s2CZIWmQhSYrNLwUtc4DyfGNmJ2C7Fs3ASw0AXuQVbueIvE/HY
HkBVQNZePyz7/G2CojVVP0NN18bsnTg/RBdTd+n1qtNRbRm8IaVFGUmotWkPXkaP
ygWIKVPq7lHpTFkAB9UXXgkdRPm10WFn2e0ykk68iAFGg+hXOKqAnvhUeAg841/k
4JxSTgykYvxcXygVt0Pe+1v3BfZ+nW+ojFFASgbxH1WmGEULrSjy/tYMuX4iI1ve
d0l0biwmwpbbsUbFfnk5aYcTloNIJIgKbvWY8geZzmP8cqNgzp5vzkPiXv+dVGR0
fB8vDDuvv0r4+tRsT80d5AGLRIX9FVbRX9SkqqJMv/RO4tqYKBQMhA/eBz3tMrqc
DGIDHQlcpk5amKjbyjbceXnQAWlEMSOgn5NtzXMpvUHrPXZqTNX9iQbrQJSu24mm
DR/3jUbi7k2/hyTcb+dIJNT/Ct0zgdHl1QtTiwzYHEo/JMwvqpTF3ieuH/RLnfkc
NS9Ax4qRIZKTNRye7KKAe4ny0oHBFx4AxoTqQ77m8jJxlmSdcaXFVApMeX6ZeENJ
Mik0ZNxD7vqLiXMz8kj+qOLwFOUJyOvotR3bNegXR0++oir/+0sflcorxHye8xao
0ZZDgaSI8m+rhkCUVRN+OT2zzjqXcihN3S2nxSa3ySsyB1CmG4s6TkUP3e9SCG74
F4cbfclY5SUKFOuk0LdLyvdvJayJggbMn2tCCqf+ayHQppO+bmUBE0dQ6GWOu4+p
cY8SJJLIX8t8/zseesTphTwXBKjmcCBzTBi8HFwbaRXelLJM8bKOcZ4MvWp8J4Mq
DKCriiHsc2EGQB6TGZ1HzbqsObUIPMT0zGbejUZS3OCM1dAgM69H/OkFBZP/b1AF
VxX4OKd2iYR/HEJz51fXTG7B1FajvWNOoLtwFaEiDdl5RTN8f1tG5+kaNW98qpbY
6anElwm3qIcluxspUfNuGcbZGxTufzGUGDlW+RjMHqLtuqjGv6DSHiQfjOFtK4jr
6PJddUV5ED1OjLVOviP08EJ28LSc0aZmTnFt+SurhhXQNyW3AL3MybbnobqUW6I9
NAlsiip/X0ZlayjcHLOwNrpg+W2JMs4Fxq/SULDnUkPL5U/w8cb9SeBBNjPCKp6C
BGDvn/SRHC07rApwCkjmPZJuSEmZLvAQzdr2m7r/rkrSJVS8pmYpgJWXGb0bJOtS
JaMD1Jnex7qAN/J4hEZWtFkhN3jyZ+rGEfk3qM3tZsNLaYlIKAPx/9FbDFrd1Her
APY0Zfd9bEEMsLNrFs/j5xByR9OVzAia4wVksYoW8vcY97+QGamPcqoKk/gYv983
9LO/fN6Td00P7wXaVbsnz7LMx7xMf1oDr2k1Ye0cwVoR1yU3RSPWaoPMA/uWQRKF
JXVPh0CWtgKTAZ632CjHdAcDqW2Etmk5eto5o86J9TqBvrnjM/kRyXr68dB3uwhQ
r8Jq/wdclPwTnxglCkulYrvu83/yTge9t63eARS1zlCbkq9YluYPhLGF80hQNEWF
P45GW/kMxRgjZl4Xx/+IHqjbzLJcMttpps9rd7hPHs/L0kYj2UeUXN38duYAjCVU
YtNBGW73wyjd9PPjfJykfRUOjmz+V7M9UBJts0uj6vdQXwmIjEUZAoI8uXgeMasj
gTuQv1L1IQl/WdRdkvZnsh6CnMP4anDYpJWv/wP81dzMLFbV+tcyzpWOGkSxOwhj
xNKSiVBrsXzaZY2Hm+jBphWfhVHZBVDq3HIx5MEzrbQ/zeA+x+rqQayAi5A5/X9e
vnOg8s5QD/QSRDkkXm6oy839QXLrOAsxmR25IKRVj6226VDYJO7O8IjXiwCauz5y
Q+Az/j+d0IqrdM0na5ufZvn+vp/mqNQxjSUsCjT9DsHEezBdHz0jvP/pg2JcMdpL
skgrblm5fk/8q/PoqiMNI/IpjXvNHEtDViooSN/fpv5wVyhkB/U+gFP4lnoxKX57
U/iMCmmt15Nd8Z3eKTn48Z+/lRMWhwmKdKWGpB2r7TmL2QRq+JXSN3aPOf6tf3yy
m2LWx5RJiRqkONXx2m8mDtBmiBLvKPEgiJOlAK2h892Pj1CAj3mABx/hOnQPME6R
tm48n+N0S3Y1jUcHwChALZJVaqpylBbJLZvRM80TF/4ewSxE0G22rhKtsWY7884x
aGhoDTRhW8XcBsbWQUAiTFV+E6cGIahD06BzdLZh5BVjlwC8Lz2/C59KNbSTbfW6
1r2Q9OTw9aXRFWwln0j/Vf4S0HuLkfVJ6FMrwItJoJCs+Dg3RBNtrBlCPIC/qqlM
z9PqzFbecSxkt70KMOkVXQp76nug3pYUXlVipphW4Isj57J+r03IdZaQso771rLG
1XPYj508Ffpl+MCB49jSq8AR5/QPh163TsVDqGzLePl5n8A3hA5w4u4t/lfLEA3w
Byw1/+g3QeGYilN1feno5yi3qR+KurqsQFsmFjRoPXBiEWjfGm2D3j4Pn21E57AG
8hFXTZFQxNHlrPCfWF8rs/UBGy4es+/aUCcgU6Dal5DJVO+Cl/Tl6mDV7IJ5c2WS
I1hER4xOiMVKk3sUX+IPQIggu7nG8H82LJ8fOQMBho+AMASvFVXLKFBz/h7uvkcV
rGK5BXBoJn7PoR9NRp0uyGa+Oekw9p3Vist4OYH2OxTLMSZ83Kc4/8x/tTkyQ6SF
Ho4NOEiulBGDYMyQXl81q3rKTYFxcPjWsXqOl2mdjTKZcLujFU8Se/rSi1xkejIs
qT+VLzHhSdZTMWDFPEn8xInJR7O3bCCTZzYINj5FnKVxrJKvNTKkg04W0dp1/kbV
v1Ix0FcieKO0ugi/WeEkYA3dmcQb4NmKcs424tMIVK3rK9fJpBuN+weVCN6Xu+tD
zEpL3k/rNuC5AI9N7WGxZ39OxpSw7fUKnbG00ouRPp2Dlb5oJE2jj0rKqoAIVN2Y
3uTbFiN0hqYJfRJ73helM4tyEM7ReN7Hctz/AToqNGzVy4TkaLSohBrEdaFwSUSp
ThSDqGAkP5scTcRsAN+VmflZcegDFTU0H98rV512NUKsjpnpm1hyfvgzKmSaxJ/e
5zQQ0uNo2BABtaeEIDfdyb48zeVjo0yKKDWvrjIL+FihapoH6VIshZaTHEdkVPVD
mOo+dTdjvbowS3Cqf5O2wiqJvmxirEgtW6jhhOtv5htmLjvQnTAV73KbGluDC6Zd
fnxJdzoW1y5KEDkLqlOEYE6i/dxnv7D1/WX5xl6d7KsV0P15l1sqz09Umf6S1btN
LG6ao3wflK+RvOWmzkWLKHmHwhNcah0vGYXBDyYsRSv81EseDHj9GqOt4oF1ByDe
64kgjJ48tOKSkY3Jz1tg3Y+8oOTxsFJ6H/5IDlMKuusFB7iBJnHngDuRk3HsTavf
FDv0GlVXzFX8iLve+vgG4i5M6t3gF36+WpbqXhWJ8yZzJSy3MZorh4QVFE9fvsdD
jVpGxIelC/tPkgjLafJsxVHNKvv/B/5okfYySxCGylXxfqjQImsRAxgiDJI8S+Es
i5jD4/VlzEPFzZ83vsJW+OkXXuP46G0N3ZoxuvjcyhhzmCVPmHoc99abBbQ6RmbJ
MuBNBJ9bodquhFCu9CRtBt1IHdC5Xz+Ny+zgK3fx91H8oR14+RXiWAlXAng+TZMx
rZWQBk+55TtAE62zIUeRvKG2NUVjqroiHnBVcX/rDopxwfO75JSV/UwmRGS5ERxm
pHWGNBERSMtqXO2JDA2IK8yxD5aBYSDD3EUusFmOsK3R06AMkikQF2mehMSOT3eG
c7/PezbHwQzPtNTedhPcMHk5aJnFqP6IIyc5gCBUUePJ3N8dqH+NZZVKs0O9JECl
wEq8vctuSGaKUI1aClWwoyGjJk/gcfd51ibXKRA5jQDRTq/AeEd0KncGY47EgDRJ
/G1y2otu/a0hOMgVdmWZuR/HUnLlZJmPExQBIoajTH2dOVHagzJYmic9T9suCDrA
hvjlDhj9CBcTrceiGuvIrLUB05FyfmtF53jY41BdntUfSRLKT2C3V/T0SK1Sc1CT
zBFNRqmPHNfbQ4SaU0oHCU3SKD5FCq+Hp7gOq3M2DwrkJ34xPHm6OL1TBk6dNz9O
cyM18s/UwZKhUf2ovwK4Qf2z+TMHJySgULlblv686IAJFOtSCTC8U3upiOofjr0J
RVjuHOGZVxSsMmXQC32RDfe05f3YLr+TrpQecr8gUKerttUjuyno5kUrmjGtjadY
Gi8lSbDbDrRgrGilqzkcdbUci85Sl1HgaCQyY/EWED9OyYrDgOabcu5NZs3gCAHX
3zjUMeyjet3vorxrp26N6KGlMZk862p0ERVz/4ILGkgJ7APLL+t16InsWCxw9DB6
2BB1V0UaUaWcCplOrxtE/xGWUx8sjzGlKCdyrA17Xktq21U149BxrOET7IKBj+FW
XnYPpEMJ4k3xxBh3ahzX00wbO+6AvmhN3oEWOqNw/vApCOHTq/XTXC4v108wb1SS
C6VY5nkDZ5vwyL828YZ6jZg2eR3TvgQt7CAL8FxxlD2pnTNnU4EOHXuWRd/8Jxqz
8q6ln4CNJfMw4/otxnY9Ydi4s6LraTjGPVxi320WfqNGdvl7uoWjo7yeMNXCBMjv
zxexsxp9Eo2J+fuqVAdZHNpr0im1aHCkvHryLw63YRLCpcSmrSWu2s/cM3oa+cp9
Y/cuzL+W+Iw/tp7CE2drHJRVDbNNsP49xDawq4gDoea/aqZusSyDyModUNz4jxo6
W+rTpWsfh7ZTmkADq7Yeq70gqszUqzqHUn04vLhj7fRFesMW3d/fBkeD9gVwVTio
eNiLJFd5ZjVh8ijgzPYGWZO3+nWvwmkHGR1sBVHWGCQXqd4rTaY0ZKT7h0C7N9CY
rv+/wrcI2xfKCwuQzyXY6wbzhLh8DJEVHrZR8RNrypLW1BCZFlW0sRjijNzSvajh
XrEUdTGxHpfOOo3b0XtWmDJNJj8Rpl2DcRvzEDNcY6lXzrehBTt5SICTV2d3ffx+
oMdFK98cTR5u3Oy+rq6VH+Ied6sOJgwQMGX0uLymEY+PVML7isxmwKEXV1TZs8sD
sbwMSS/iYteAP932CX1907azSFK102DKAnqLr5QX8iMiL96BlmQ6gM0oJNItVjx5
vruZwohO71JdRX7ybF6HHof4eyDLd6mYwmBGxE77WouBJb0bXi5YcKmtoxtikDqy
hUhUthSCMZ9xQrcG9sUuP4NjQQwUrRONXbPSoxuShvAbScLAVa8jLU9QNlg5Y3kV
OApeU012HMH9qp7H1IE9UKgacjn+pXRTM2i+mM3Jz80G4JSvgZnEaAELOWimouoz
VOGVtFSbvQuAchg0PgOpohpIOh09mlkm0/yItwHiOiJKeXDZq1Sn87MgXXQo3txr
Ikn2LEPu0rgHX45mQaWrdPU9f3ydkt2V3nm9yVrVBdUgyNGDuUHu9BiOjW5tCPxP
/kgWVgdT0eQGitIactD/nhKmdj2S2CWfDOAfMaJYDFtAa9idLExang5fs1/3AI7U
UP5qexUxy6TGeUQD4Eb6LiR2YaEo/1VatKTqXFQ2U7O3Q6gMIsyJPRro/qzSBXwZ
KIoThjaRptadlI+pCgyvJ1YRjEyr4qEHzEmwqlIXhQKpzaZPRBr+cNU2qTxp7hQg
681a0BJknPRhHcFjabq5SMIBVQBJGkbh7y7c+pNuYwOXh2hvK9M0RGHA5ypydhCP
/bo6IOqSI3OU/ElSNpmdCYhKlZTsiNSYZx/VomambUtrHJbV7ef265UB1iQIUSmV
a4/fuFqD9OxoghQgBIcIFli+EyyX6GCC00rPqaJS882UILBGYPM6A6kp4LTLXU3I
R4YBwIw56apkHmFmjaJrTRK/v7grLoOTF6pfd5xDPWY3KHk1z7ycQ/VwS7e3Pg3s
lVV8BlbiMiFn9bbjnIi/7gf6GrBiiyTKy4z9HN/t7v82ZyKYqnZPRIUR7NTVgHK3
8A3Wjfjv6Toy5XK6t+MG53QPpl+IcxRQpLGdckRVyToZLabRPGNs1VW1fqHsyLjV
Of6ttTScwEbZoQwFBRhOw2Y4B3/ZPyySqE6JucJvkakhkH0GbsVVZxEE3R49h9qh
mzp/lOvZxXfIe6kl4nVspJehHvkuewc4mYRttCifldpiv6xsam0jsNhO2APIR3Jg
AJSJUwa7XuVAN0EZ4KyRJMmxhGdD/wXhI5cbU03cLp1QrBMkK2Ko64ciAdWgRzCc
3D1JoSgVPGQF9pJfLFSverjultzILKvOqKMMbaxBMoA4NSwJ3nxUHO5X0NBJ6tuL
w1qWC9b+cOjm0SdlIOjzGezZwhbx188p+nbkAR40I8u6X7W0Q5ij7+xqPoIlw0iR
/jG2o00NXrrO9vdnZmrPyVvm0fa0r5hgMDfh1DqqMqRcc9skFxoOr8aKytqJH0jq
2WDWkheJ0GK0JpWGrBEJcYneNbwz4yNcvfv5KcWHpa0s9lFtUCoWeqYwFWkjYecX
1LM1mm10vzHAljkmY2HetZxZYEpAmVbN6Jx1njQlVOMnCtyvPDQY6XQtmQvLDSzM
5Wrx3AKUJqIa/yZVoCJoiavaHr0wBL0WWpn2vnLwtHJDbKyYd45uo6Ov5kvr/lID
9CQ9BulyjsIBZAoc8wSK7Us8sBE6yd+F9UJBylH5JF1XJQ2PHu8i+QgeOu99uz9L
k0Yi8mfes4782NUlLvv+8LWcaQD1B5LJEd0Gxr+52mqS0gA5//0cLgdQ2hKLRwX6
XndNyp4O82QVfHP257LjNb4YhlnXJGEaTpyd6nL0sOh/nYf2bwwapD5gK5VyNCFs
cEXnEwvfyoYIEjZOLT4bY9jkd1ga2qclBgrBC8xUE+VxrAoOdpi1X1goqgrRFvhn
2ogyCPEPJxupKKWbffWSERZ/DCpYdb8CVqyckASufecIlbWAH1zqqWXScMZSTR3l
inHVz6PS4zS7imww5Ou9OpRtE7SpKFZohFTlr6jn5EY3WjN7/RD6Vo3Zl4Bdmx/G
yMgjS7k3yjOHolBbvjn2axg0F3uGg/9i/rh3vW8VoPkKS7wn/FiHQID2Lrbk4PZs
iXokEmmGi4KesNBmENTI6gtV8WJH9y5QiuB6OlHgH7uw11Mna0mE9ZBCfEZURmRs
eQy/x3M7YqgSzGAKmtmZaUulgMyUxP4IsRlvZjHTPb2/5golXFSy1eq76iVltYJX
SEq7463WdWGVF7DM3vkD+k+vNQgO9UFPR/SAH+WHde9Z1/oIk2mXtn9KRpL0E6no
+Wjs4VDFjpeBNydBgOJDzsYfN65cle8fukH5p4DpAh5S9gAOsLt1R5to5Eckptem
OixJ/P0ij/Qw8yYSQnQRKbamOTLz6pfSMmzPgStOTM96+AF1skh/BkN9AuwbtEus
PFGMCdn7aRuvGK3OJ/VjkroEwOfcYx70xAnpDFZPGI2BZBrD98PssFkCaVIPTess
S6Bd6I31aLVDjRHm+PZoYmhKEjHI/vf3h0OtpH+4ZvQTNDX2zKkfc618SkEOFy7H
4eU9Jckv4DIgApxDFkaBSv+Ol4qT2wK77n+IcXH8QuTA0Kr7BnIx/mK2GZy7ZuxB
AB7lZ7zHEA6pJdfsIX4jjiFAUgMGvs417MfHr1xGUOA5NOPZvfrPNru+OcNs38U4
D/7wcFrgkVS9Ik6+lQGZpaqrYgSK2VYaCAoIoBMwKRAhGl3WsOUdwLcCyBOVsH5F
VH4OM7BEqAdZE8dD/6GfV5hU0SCqQq2A1SG1q4jFE1uURtHMwCrpz/VSwuE82rIl
QdI1kfXAS/3UzGmWNFITdhvpvAlgv2pGx+kLkY3/Wr2+HmP17VCPdV510RUXsjju
w4cwev3GcrxdrIbB9XdNgRQlcuxU+y3HSjJMSrtrCOXl3ZXjmymiPMif3MPnkRPh
Lgmp6vnSIc8hIw2VTlD7Vt1L5MN1PkTaPBQ+78Tec2w+Tik60ZxJ1MTnIqOBJ0Oz
ViIeIdlh7sYhMK1lzSB7FQIznlMklqv+Kn//JW2y9oBUGsDO+yFddifrlDSe1RCs
e0oCRprxypDv3azMMnmBpWBR3iXMDJqdo93rILM12OQ9pP6ZN5BJjwdWF9Hm6ik8
txuXxr5sqnP9qp0lly5YeDpZhXlWDwOvMrnj86aAe+lrNiA5OfM/FfJsA3nhnYXW
kc2Rc4WtC4js3QOPlCXr+nz9PLDdPPkp/HiQCLGANdrOl/1hSqo5HRu+VxyG4slr
wl/abEnFlXh1ch1vxyxYOKrRKePq8WWeq5h7FtxKs5o8KDWWeCeQS+4qB0Qkjn2D
M92Q8pCgUiYf/9IFJmA6F1ZHRDCjsxH/5DFFMiXugPETKY9qRUZySbRyGH+G6cOU
6uhvZ0aluzCIfgelkntZ5hDZ44B3ZUnQJlvDjW4662Mk90j5VQTVeg/88bF7pbr6
Xuy9RS7q5U/tssGyM/nI7vO6NQUiNOqCwfCfGaSjuD6S4Pry4NZwKyZ4dRcUg0RP
yAm6LRLwwum0yeX1rnRsiyqxVde9Wi7DKNEAD5qJwdNyhzCSWtd0ZvHJhKfW1ocm
POTPwqkEdyZL17r1zP0ynEnTFVHxR5Ap4aHjcmkPd/AOreeMd9lYhEs5WuRutjck
oXHyqUV5gzIjGOBHPZfcVJz9T/E5Ffwbh8Wjp9uMJ8lODhTYBnoxnoOiCsRyI+6g
JJamtOP7Nfoo61UkL6iSE6dUPXYPplRaEFRYQVqZ7+CnscceZJXxtBFAmDHR2uG1
qQR+mjHqc3ZShwvgQd54/2Q/aNTi8DLgSFFr75QjqWn3FPUruT0s4gTmmCS8k4iU
sDtLJrzg8lt6W6bnK9sgy14IkYZc5I1c5DudjXoX8TM1yKh2OlDblwBMDgRS8nKt
38MLtUoOqpxJuCyko/mOQW/jquG8eRtoDDp7TzKobGWDxK3jf/tseEqc6/0Hx6c0
tnjRVpPii95mO7cuxLB/3J91I3YykAMAegS8hR7MUUwXf69KOsax7x9Hohc/fYET
ACVKf6bB/K0runDOZIgyK0dJ2sZN46HbGjU8XSf+AyTe/G8AdNlcUQpprRGmjlSl
3rB1n/dbv+QZSxyrct5QP7RC6WsWTsjcRTlKhFb6DV1Xu0OA5mwZoczylV9g6PkH
ncuUGxtDoRoryPnqHcviV9OSeIg2MJTylH2Dd2Z9vLxpxYkuzba38OG/QY/AYG69
vE7tkN3y4KHrYXaUpoEVKkMAXbNYB67u9eByjqwp9qKEPzX135IibWySMYHvwn05
d8JhlIQHaHded8jxZhtnmO6hDypEyNPVryjGiVPNAgWJpG9uIGZgfoTvltvV8sY4
u5qVHNdwriN3OiX/aza6jxF7dfGkSWqJNa/LyyKgR+PD3RtTcIrWp55mdf9ix0V0
GlLHeSNOc0ztQv20/b6rl+/g3nZoi36QhC0OyodCEjuIVLB+i+W3ZaRPxcqz07We
G43dHu/nJToGadDnY5Tgj/DXGexGJqCXWWUGHPI+z89RvDUZGZEXkUkuBqq4uWTo
nTNY7B1veUDphjKxHD9z3qJN3pjZ1ni44d7zUrZfq8jLP1zV3Lg7x52OBtZ9MHfu
cyAi2xTwqYY34Rd3iaU3EX61ymaqs11ctwfhjxwUQDZn69ihHstLsmqYuxGfBTfh
0P6wgXWJBboR9siOZwUjI04sz4XU/fUYxAZXOMw65huvENuqgGFXGEtDZ7FMtfiN
hXP8Yyka2RLMzLI5Ckg8Ova6ssRAQe1pIFSMMD3zKl5oCgiiW+2rtW4LRc6inKIR
FWLH14s/JzYrQl1lr2GkNdYyWQZb4kNQPLOi/jIsOdnwRBHnS3glz78I4MKc+tGM
3OCagPR5vAy7ZuMV2DHLH/scVcG3plqQmCZNTtKvWAOSSYertE+8VVUp1Hl+IBTq
i0YbpiAr8XfS2hMXZPMHV7s5PJmaJEzpQsldQ79hB7NeFVtDSGSKi7hfhpOJijCV
M1o4SF7UsUMMvg5U1WGs8Yj9y5WdOjTydIoC38ScwpmeSouC0wsGXdd2khai9V0j
vOtjT9/jsMO+hgzd7WMbXs001NUS0qTg67DCfgMd0fQdA395vatRCEiJin4jkeQZ
YqSA/ipt9kYTEGQQu71YRS9zCWbKM8HTZcl5ogX7D14QwnzDGX5W3AA90XalpsDO
vaz2+cOj0kI6avuFS8Dy2l4qFePWlz1vbyDFWI5mibzTFeoWW0HY8S03uS/0bXU8
FnzpWcfjZIqnTKSQ07snc08X2UIyRWn07XtfwhisjLClT0pWy6FOeLre79ohJA/1
HhGjm2TJTMHUZdYdb/mI7C4ya4RuMlEu05XmJW06/DbNk8FJaVIJr7aASQ01e1Ss
oLN3Ix3lddYf9KjOR2CLGSz2CzWixSBG5P3/tDegHJLBxEpXBqOF6DBl+6XLl/vT
jZSqGDyNIkITq4MzV9VJxsF4N/fMCtJHANq/jHr3GClk3JzfngWsf1pGR+CQcpHd
GDMiTVQBe8EXROsOlOroL6Jfvja5d5HEpAAp17nKGPkDAv3lHNzeOncEFwrmaR+h
2hzG5BEN8LeQUk7REx2vE8FxBaLCHJ8k9cuh/fhZ5DPAjt92LG3sUvRW7QQCj9Xj
gS69BYXSOX1nLPQs4thhFPosmuE7tc6w21Sn5ce1ZUVELaSectlyoQuKc5uu0Khf
oD3+5v2ytx75uO83dO4HTZFHUNfEQKxoAkQyNhsOpktli6NDHpklmvHrnHxn646e
vrN8J+v2Q8sIWd8DiJIUb1XwSLgUJDNISBmOrejbkrEJVNksshPNTyKEMySFeoYj
ZCYKGJ9zRBtuYg27hvAkaaWZWahteSy4UxVNr9+gdRYX7NS3a3uIwZ2Z8p7a8wa2
NVAIg1cCoD14c++RodNmNUyZmlvcpO0cWoWnLwk47eyqsIgxbc8ymY29oPS+WYX8
PfnR11BOCMr5+c+Ar/IiIt/ne1N3+37/ZHfiwDWeF1yRJjeAyhnC17HMl0d/XIQS
lfkQ37ygJ/dxuTEx4D5yrZNrPg/mAHEXOSggeOSbVnmU1tVsPIukdq3QEGJZokp4
f8OFy0PveeZmY2YPUuGVZ+lL68lc7O79T4/bERor6CLnsWqW43U+PBDAzmffsZjc
aGijkUVSF6lt52t5FyQaz0PKbInbZGEopjbMpOOofyUXwJq8XN2QR6UfR1QZYbO3
cvcHhxI+lwyjvbiVOAlDxhnPv5FcjtTs6l4dacXAR54sDxOhjk7nF/VZ/a+d2Zng
kZDaXzaPgZ+OpanIIiAJyI1s6XSxAI2xLjrM3SCLIYBN1UNQjznqbn8OchdS8H0m
ypZEEynzYdm2/ZUI4JyE08vJhX5XfLaJWNbP6XKgWGRraewFDNjiaNXPiCste1I5
YpfvTxrJtzMvi6HJst2/QMngVT+uxdQT0EhjaI8NmHBFNOrBA6aMU0d5lDeN+tyg
/d/QJc2bld1n41yGsxtVIw/IMFA8Se3yr9E8QIjtddkHgeR3RLaDtzWru3/C4Wne
CyPxsoo4uFebdePrVzXWR87s/ZD0XQVRbOfGasv2evaC1NVQX4QI7TmXydrDQsy4
ADJPuNGi8/ll9Gr6Ep8cGMFoko6JRc5lWiIYFz1LFK3Rtue9kVYK2bQ56PK1XHFB
dG31BMzegJ18cUPodszd2zuS1Rlh0S8AZlzEy7Ig/3Ull6zz8VYPN8l4mjXKsNvf
XwSnYYydvF8gjHRXSCVAaZ22kCeWdadvLdKNMHGslb2feKAV0LxEob1LJ7RYUTP2
VIHcqPtbaH4ye5+5XZ2pmfVNwJXve4Fhn/HwTPkWEnHnhkS2MsFPHwlgr8NIDorw
PDq3fTGdY/wSCwJSSV2+s68SEXTbegJxkT751AeK6rq/eyE9GHfhRvA3dl+K+mWX
1dg8Qm1lKIiymH51VEwe84aICH1uRrWXrNZ8peiK432eCRzKmx+MkDbYO28o3oQB
L1Ma+fHuvMFpxxJj2hWkJjFuih/qtMHFJtF5sHvnV8pgzChY1cvqU50/c6eTsVKt
VfnrXZObHKUNnlFHiwwtl7tGwyT9NlvSqodfRPgmlR5GJwhmwlqh7U5hUOBhpUjk
+ehwC7YKyQzeMfC9UEpagb66jwPPAIyZo/BB3y1XUpx0batlxoPSi3s8fbMagGAj
vm3x2Jpmt476qq9ttWyxVpNK/yJenolLiZ+2Igiwk59BrQ0cYohxuKITrIsry+jF
9a/iFIH9GquqfKJ1kkcj7gvJkk2GBPP233fmNTXN4SOic37Hnni14gCBsyDvkVB4
pogIUGntLZ43H3el9Y092IJn56rC2+0e+OPAO5SH7mKL2FKwYNpEjUHbVGmOjH8D
IKS1QGrJAVeHvEY/SAWK+Y7/IQbFggKRgIraYAomgdiO6ddBxwFzW0JEoqDEHHtj
G5EmxaORtsRx22YgbDBd7k3/PO/tCkDpVGhV0vY24P1wuOAATqpP3o0rLK0xknxu
l+Xl4pCNLKtAKFEIwGO21YMu68HSoNtu/qYNWykTusLmZzL4o3dw+wKFEpc6lIvJ
jc0YUPxgN/5cLIKt6iU4amjGQ3FArXd4eo5ztDWpKr3OMXHdR+G/vsM0k6J28YTJ
TxBz/v7SUXRsXsfKiAyTR1HWfd+/B4ar2O7sHGgpbgI9sNkINweEjj7vkdb4Yw5K
p8mJJ30imskxnhxaps1GjIQ74RCOEQZ0TsOtnWY9mU8aZeaHvkUeAen9e8yN1Hq5
F2m6D4gJRQsW2YQRsh4JHhjAgdi4nyA4OCPt4en4w8x6nBFEEhKEzyj5jyTP2jLy
6F8k3QsOVHOmnnobTHa3v++aA8xhi4jra0OBBBfC9W6p0vThwSs94s+oERlJkqy9
liNQkB8tz7I8GBGoFb+ueHB38BBITkbM9At9NKTk24jI0t6RykVYutr5VrKfsxQW
EWPx0TLPBkyy8Hg0a8wpcC57Um/Bz2LFSdLH/JEO2lGvdxNCcoDV0kyy2RX/LfU9
IMlJh3oDcRVEe8icpHXR0yRvpmfgOIMe7CMuyB4Mn3aPi11ukIRFr8Akd9K43LRn
3J+zOFqqA45mvHAfPBYWX/J9YlL7Mqut2uxZYQPsErGO22dkajcfzRC4uhrEUHTM
gOQKwC3SSVD6iihU7iaoBArXBaP2IHrrxGER+bAT5OKRUjQ/qOWyKE+qgPdpAzUs
qmTAhJ5qcPB10BfyoaP853aqiEe2JDwvQQQ3RL/+X9fuSulJFYVGFWadq0OhIcR8
ob3GarYpqDEZVwY6/Qf0G20Ky55HA0jerIaV/pdi0eqeJqvwTXPmGOUVLl091Avi
UlAKhRdnmr8Uc2f77FYoBP/x0M7K8tpeBR9Cp3ZDkAerk7JDZFzUCfMWFFP70FQu
GF/DxpC9xQuJYHpPH6xkp8avFqHyb7HcOGdPmoFxylifJqxyOLqLhUQ+UxRqnSWJ
qpMBJA2yyeOI3WrmtxVBfWG7jMp8NVYP9kGeJnulIagrZoLyzVStoQAtvf/ysUyi
bYiixvaOwW+/7yp0pNVQiRd35qXC0sM7RR4goULAg5Oh04c2EFibC+V9HbzKuD6W
Mk2WmwPZcbv+iYZ8D6lRO3lDCo39qh+/1gphLCoJgZSi/yoSPYJpV9kNFKLlbTVf
6Au3UiB4ReAkxwe6Ojxl34RGAfzclkeX6UIxbz+pGLL23XV+pweLJnP/cyxC5eZS
b2OO0Bhc+8hMN27yh9TLsrN/MAaZhf6IeIv89NPgPa05ZfQ7jYarW3SUcMlWBxeR
GXd/6DqhT62gB+1SAobBZ3VUibuowxgTIbQJQBNPFRXdSQGbHF8DvR5vMYDNz7ON
5XTbAl0W4QFQ8/r15QaArtZThjtzbfYnlSUZPxwwJuk9WLpgzP9P2UQPsRZVzVrA
XSy7hHjWOZTiQTcyj1LNjBq/JI1HZqWLKKmuj2QCEMo5r2eYY5MQ45jsoSbzQ+uB
UEWCnftrdbDD3RD8O4Aer3bupq5Au+vJ1FT+OEZ4DsQheMODUPpNLIZwkHsJYdU2
GoMO9QsArJzA9IbedOYTrfFNYWBs6NkZIwq5HlICUOS70o3gbUELaITcNagEN5Sa
hwqcU1VGSHbJoAq2NG8hfPTdFvx9FlNaZzl7YIGaSDEoJ6tLbwGd7rJQUwjoAI4d
LO9cRl8AkPmvG4v+V1BYWN+uAJKUWTvFl5NhHF7dejXHd+fLEKQtGwLY8Zt1aitk
LI7IChxjqqq0wZawQjOr3PRC7MQ8kwVABGntkacJmTVn6B9LKRr9DtMKd1EFTutf
XJxdm+EBJMj+9gi+qv9oQMgPMHWTOxP6bSVio174MN341R953OlHeBsscJMgf9k+
afkTQLgN3iJjibMgh+Dpya21TwsMUwu9dwNsrAccXOkh5DlKTZmlwdZbzZgNZKqB
af2t2ucA40tu5YEzy1+1+BHu88O7Ns6vXMwRstNwUZo44gT9uu+Yjhna59/pWysn
iLDTpwj6fxp70LTGiEru4YadLVXUHU8av4X9tYCh1afTzEcXe8nF824pg6x4QfgG
jPIADHAt/i8jy5yj/mzqSiH646lYjLSSb1SIcJPZNgnxXbCRvnc5UKoeyrY4MZY6
adwDvvvMQSWG5mxdQW7CD7u3YVf1K/eKXV5Nc9VheiCCiGwRV0WJ9yZ18LiQzCmH
cGdYSbq3nzrs6n4NmnVR3wXR5naeLoQeMXwdH8Ynl1ZGaGs7723dFPIQOFotYQas
5HTjJDsaSNyIhgDF7ZfCFzJtAhaQLwIWrLckDn0N7CuAk8iS5tBXKcxFXcbDVLdA
iyxTFnAkwfV+QTYe6gcfvbPiQKMxvDB+SfrkRmVJwYfZei0GR/SzImItriMPKvkV
CU0CEQqGT68uPHahwCDjM5Xh7xPOYTwpSMK0JnvltBjQz8v5+dhn+BQNIa+9aHss
xMNxraCNjYi8smNWb68SmfOZJkp1o6RAXNeh7OH0zVCelAsUgaM9LvfHSGiFj4i6
k+EQ+tUwDycKKGsPlIWk3wrEY9jgaU2S+4hbBuhUrrLvoSVemt/RKk+/3nJNAjUo
J354+H3md8/1DDfnT7EPyfmqvLTuMgv2fNra1umdB+IiYj424WFQt+N6nYnFqYYJ
rME3qI9YdfNiqrUtXB/p6j8HI6YC6bMC9MVyTOfatb4v8fsDyf4SGc2F/xS3MIW0
sWd5QiNpvvzKtksSa8R7YuaE6v8Riz9PkImtrOsAVQOyICisinCnmxS6VzMkXhwH
nhFnpYH52k2/zDo5aPpyLKQwjo7tAx4UeEcx6KyzYTewgnI07DUc4iD3lnwkSn0X
h+BvqCOVF8l6yuEeOlfqmiruuOTrz+1X+90EK8cQRIkdfKG1uIaWI5mJCK7Kdhis
SYkY1rwZ9FS7Q47NSbys3J2UfOX9qfxCPoI2cznDs9XYJyX1f+THtk8+OJStcf6a
Ho2bNLGl72c07hmWt6MJSUYHJOhgxZ3JK3CSR8ap/IFiZhMuR2Z6nRfdM/Bmj1jc
wFren3lM970St1kPXpKtTwuQmUDBLVvkDoP5M1tW1c5RG80mElQldVnpMfTcL9Vj
FZd8VuBLJDigr9d8CJN0NKHT3z3V0tmXk7GvRRqwIlFG+Qz32mV5WkAQNAljowuS
TsLB/Gnt41PPLTvOMPKXxHSjc/ORSxQpoiUucoReBBgiP/ImRVSJN0on8WS3bzKQ
y0fhpp3tQyYd4HpdN7UfZdU21GjTe6GY5i6QJ44+CRPNrn9aOINe5X/e1/JYwz0Y
RoocJuzNsrTvF4XloOqtUlQYzsRB1H/QzGi/5wyGVJPqfhU1j4wOrFATAzHcIiz/
VM5rygKagZ777sH23Zfw+5/ZohUeGvLZsJyKYvhQDcx8U0D5LK1mcur2rVsdt1YX
YMjq5MhDLHWKkpqokkSGfsUbKDn1q7N3BQtv2WFhG3S3UG39qT69NK0jPtoZNRnL
ZEsQLzVBK+K+4LuqSfXsPBQwayFMqecHgZHLz1PY+BS81alnUGPOUrhyCJzmB2DL
W0d7/jF/sice6YXb1UuTqPyMgqGIHXcUUca/3QnopKs3lF8WsezQyiG2fR8gjq9p
Xv8IG9Q+rPEqHwJKTlLAYtRLSCJBjVZdcQ3JtltsEAfQMpDJiOyO+SS2wQagqTzE
4OSfizU4jtnrkHUNvWyMIV3V4NBy88XT9yV6xASKEOy0sd1v0BLse/pu4i6XCEFC
GNAjZjHcuJe2MuOqooBz34kIa/C3PMJ31uIp/S35T0jBB8bJAtkS17PgbkDELHDw
14PnGElzgz9bFmB10jRA6ivvn2INRyMM+9AUE8aV0IOzIb4/zNsItVWJNrLCTE73
BLLbu4ETFUDEzYjmJFNrsETI0PTfN5uF2I9dEaaJkvz5HWygi1J1y7o0v1rDmmid
441yZeK4csL3Fi3/eaXI3u19upkv7+lSzLNMN9PgltQiDtCx34bHa3GnbRxIV4dw
E5V3Cr7yod3N3S7TriY0lQLOQr43NuYYeI1wIMq4rksoEjFm5oeBFe6MRKY/W6a+
cJdfx5PmbJWFrnpOw/vS+iFjgRnlc9jLn18+BOqxzc7x+EhLLqEFKGxW/aAdkRTs
aywldE3I0P62vDOZuI29wKMYDxapdIJgXP1hlqtggj76kybhuW9SGG1FsSEfmNwO
ntJ1gYsKzIZzTw7fAUWzLUr3hPCT2HMaEFQL3NXg0eSUurg4ecSqnzCMCJ9jVA+0
71kRnfvff3BIE45UhsPKHVp4O9OVNWyDwNBLwcwIxgI352EwiV1RM9th/lClEsUQ
vkFPXwdLd1dDXWo5zDUFROnu1GZEdEe6YOdrsbyM0Y3liYTwEFLYVxboQtGfD0f7
zxkyw6ngj06x78r37GemFwBi18kz/+5WBAxh/Vc22vVyFSx9aFaDqJyl+dYpFLRp
Qj3ievWz7h7OyPjnft8s5yF1WJ2npsi5QZj8zH6dQD0P3KkNJVRbp0VMQEf0Hel4
zbbHE5Ch/GeDttMBrpGl/zdQzyYIXmwy+wR8rOC5wulTLXCJure+UhB02ZGyPU6B
ykMyXHZt0d/FLbLuwfYWQzVkHJXL9E83/11d+Ktiehk=
`pragma protect end_protected
