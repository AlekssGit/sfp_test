// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
nnCqc7ivfSpDA7ZaPbqG0EnRcs3Ol6KAVE+IRylQlI0aAxxRuGtXlIuuVGDOofVP+a/v2qyoof5l
IQco8ACuTDewbsGr1wyZj1B9toDG2rPU6xDgtMaRyn3VNt+CPMdIPAFiNg/tsGhC/gt40JxOZaSa
JYV6+/sV82ICHmMNJABKnbQkhwdtShhaeWV7/SqtgTueYz0q1uh9zFww4h/gu++WTc0oLC6uaeJm
cYxXUmXghPOx6uUQroaS/X8TN7cTJigTzrDDaLOSgPi+LGXt8sQaz5QQ59XHI4MkRSkRfeDE/b8y
jHjrCfVAjyhxVW8PJblMQ7cKmYTmaOvJ3kJqpw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 5088)
6zI6tif0ZX1NL5LgNZWSEq1JawrKyO9FcILiJ6+Oe8ZRBQmZz5E6/PZXi6XNQ1qreuL3xyo4td7+
PvqrydTsp9TMUPFqHD2T6SJ2guAzN+q0qclyMRi8dQMwnggimYC2rHfcHNar0BYKpG0zIQlIkN2u
8nIn1BpGAMLeQOXVNdf6Ce1SXfArHEBrgmlDopnhlnQyPCrNVVgsGq7uP73QFXyOtFntyx43Rk4K
tjvH/DCUNFlZ4bOpoTlSL/JvzI8AN5UCZ85e1l5ItPGvfzw2VmAp7OG1uto98RznSq8LNpAl+JFs
9qCG7jrcloWELr+0daLRVMN+pa57rf9OqQHmCA1xIMpAtl/wlOJBvYodysEJzwcX744uC9fvs8Un
XfoIOxPjfosEK6R7OqQfxRvVgF1/cerOq1BZkjksQxjB+1jnwkZ3Xoj3cSH+LYHcvGQc/Ll8VuK/
5HewZQXeADMLK4SjcE5Qt99eEcg61vY7/8H+L3S6REo8l7B3YLVp82D3zQ/NBZ+xNH0yTo3ptNVy
5Eg9KYFy3MSkJ3rdhKOzpd9DzIChiN7VE0BDhJPdRGd4tY3uqUZKKc1OPvT5TrQVcQsxeVhcXL/T
rDUhICIoisogc04hpFOzOFZmy9NB6LicX+cm0CszWrnOBw+ds9LcAeW2sqVlaG7oN+hCJ5TaAuQE
F8aEbms/bh92Mf60Um+cC8E42ftJrRWRTHbo3tkZmhXkQcqKE5RiuAPflSbkkpVOPyqIekNro5Hx
j80yoeU7YvwTfNzB82/TjRRQHJpdGFq0kCo/zou3Lv9L1c+xFMaHqcUf1m3w+HpI9J2yVCBr6t3i
LyD6jlAK4QqBCSey2wPuAcfuCidcfmEsrNlv+nc+vQWXgUO5CNtLE9XyN0cy4Ky0fU2NjL18MTYk
TYOlXVNLTao5J5wPvdukr37wz+ZtHMX2xuwqMi9KBSE6rmgkDl0/qWh0ZqL7GnAu6e+ZSFa6OW5x
Kvntn+wznLXFyCnC3cmvnNSJwkp6D3Lplv4YfRKW2Bz5KhTWCxDG0gPiMANzSA6zvjUAzDsF63AT
Jc/UdRC+ZFZBAt8vv57kE3echyRCn08RgLT5U8HmhQ+gcUyNVQECYxUo+ror0Mtz5qGnK8wcU1I5
jf7Gbua++y2TgNEY0kkwldduY3SN2ryC3cRFcIoUSu7B4jFrCFE/JL0Nl/qrrNwPzMe1ED+G8zcM
QAjXX30alyJebhWmLz6Le7f8thZZvC1AO9S8pNyQqmd5087237N78fUg9fPjhx3avuWmEJPJVNVy
AfCmiHwdVC5wsWZ4fB4+RxDf1ro92hzNIlxupbgirIz+uveiWMBtFUT0IbqrFohrw6Cu+svDghhS
JsvF6QAsY9jw7NDqP/0Iaq/YnbFNdE06q+AIv0qUyPOaoxc8bKfVA0ShtrrGJDXeiPAkCJ+K3Dor
X/q2kJJsuJOgMGi+r9jCWQ/eGGMdal5JTndyPOGYIjNrX/P+TnDZItpdSnCgmjdzMLlNAQqvSZCM
8xg6QZdv9y8TdZ833WEx2cS5aKhz3qp78mRoAO08dtgv0xOYXBkLDPfWgqJaWcuZVZxXUGBdXKIu
DdUKlOFfxSySjhrxja2keIFVXbwnXVEJ6ycbMfSLGLX7B6rdc+xjLabplXzGm8n1W9jxEqrVQ+0F
82/pJfTd/A/dVQj9KsAytkGMSWcoURcZMANVcVdNjAQDR/RLjzZkZEwVdfZpwzVrGhLAYYehLQI+
SUik4ntfsgBWQuKB8ShiQtLvVat4AhLRY516bNYVm1n7l+6pFL5RFkrwyuXHU+FTXa9jizd5FTKO
Z4If+kkhb252yORXYX8crsyU8Iu8ra22zsp6PvmsnHD+hGoorc1U2HpuvyTv8FkQjgROaEx1bNZW
1cqVkc4w/RNGlo2TPkJWFXyr4Q/UPrqi4jgaAdzLEt65xxfUxLOvsnU4yJBJKL+tmijXwNBx89AS
FWh/lMXZ8lGvGcz++V7vK1ybBAI5cMPF0+Ec8oJRQWhqXaQQ+DdZz7BIlgJOXT+u2YXcHUb0BH/8
KOo/zAFjNV2GL1nBaXWheuOA1lxdBqjqIGmyxVckqdi/TXHeif0VeYLPxtBFJW0npYUpFEvtw6LH
XCiY5XAtLASY8av6L0KX2EFpdydE1qDtg+0rDDC7gIf3W2dk9AGU05/U+MKcMkGYV8IYmaKErRdB
LXhVUZFasW+JXorkluYAaD8fDLTY4nooYzLyaB65s0bEdFaYMlAGnFzogjQWi8Bh7gLGkCDZhIn1
Q3FWCBhJi0PeaFjAWKIC/Vd8zB9bQzfa08zI+ozdas1s2h/3+q3+YkUof55+fwGPRedp0ANOqvhT
odHEmFnbSyivdtaM2IelhTd4TY53rtY0iw3TJmDF/DFrteBSyS2dD17rOM3pePRJ+sZ8OdNFe/be
uqlOMtRYbHosVHdxI7O5iKNW4nGB5qzbYtWBEQ2wBGUcUIpqIFaQdetnwnm/xSSjSwu1zvH66/Vz
6CI1ypHVIauINl9u/lWC363Zo+j2tVusovF6EnO/eOUO3kSiVrJXy+NYtd3OPswuytc3YoNFoiVV
xK3FuFTLgicRiuNL98KnuFPgjCzOB1PTfs+yLqMuJ5g4FkGTZ9vBAuhkjOTfj4z4cpyvnVXisOi/
n4MMkKqMWRl0aVkyQJOCA6hi2BZNaOQ49Yj1Mf5KX/V4nX9IYK4MYi/I+65cnj7vuO6or/qX5OgD
sV1nXJdz0ZrGmeEW/esT4Hoksd9Zc46zcKdKl2vgc1HcIIXHh5uvEmE7JDvdIsWaXpqrVDvqtLTA
wtsyWgz0VV5Www2Y8JfZs6rf0v8a5zMEoKwNkrGpTn847ylj1S50EDjwByAJmjlXWPMm4DizNLhs
j5lJn5mCGRw+v0yEnp8gqsCEWLHMdink8FgTcqbWkRQFBPX5OjuhiHxfr5WMuny6EA1mqba6cs1c
vY9eYCkHjMhACgCTOpFMtfYnRBD2GeOseLbi23F8Lmi2Cz4yZHq4GjJ3123a6Mhezr8JisI/maQX
5g1uFjQD9ahx6fKYjAxN2xScFqQWvxkFcqVImYyYHN97l3jWoYRs8BK93w1mjqzJh0/EeELiFibE
Ka9d8D5Pgk1OopY2gQyW5einu8bVlo/nkqtnuhdjwk0INq/mxNHkH/zr2Y4vusZLcDOKgLiUhBAp
G8r4vg/bBZFLtGYP8upGXixCF0A6/UCyFjSMKeefyw4kH5OzDIzQY6MYSCOpSeYL/cJK6LNPcxgq
Qdc3bkQPoWSbCdZTwBmSV/D12rWKdu20ZPUFMtVZKalMRza1wG0Bc8waX7cELeVCmJHWquVK9Z59
nuaoJc5LlHVHmO/NAI1Ux8ChiJ3G1PnrT7PG6h4RrwHjiNGUpm6mT/5TyNaApwiwFxXQi5dQd+zQ
nSnFJyPv8Mu+CTDYkbFYoONnn94ya/JMHgPyxoppRquGpWHNMNRQBoIYgQjm/INasLu0T9L/l9ST
szpt5Hf1Mnrqn1v8IQ3IRG35vBck1DLIa0aRjENejkQOmB0aiJlKwO6og26qA/d7trNih1EmiVSN
c2Q7futd2E8jv1I0s1XpJDrLluAbDZyF6xISfHRUfbwGj/jDggf0w9TfzXl5MBU46mpZCcow9HBV
L98FMvR0EUYIv7oJo+V0cjcb1BzZEWzQU3e5sLUHpjcRmXVDLNv0/3HgE9sgXc1mH/bi5fUIuo0k
uUC0iT+Ypmbjg6G7trcTATC9PFLOPyg/fJd6YtSREfCLqasO2v/h32Nmy023s6RjjFHQolAn5xDB
cSiDypDJpT+nxFOPBaxqE2h47BBFYhkm7HJWoT26/tHg0KXzUbG+MaATeSHcHlKXy3Tdua0ohMXC
ZRRMi3cvVFXnXTnSFAU9jygLHPNxs+LKJipEkMU1CFK1q5FkXI+hUUPWo87Vc74H1o2s7jxAHkIw
5JOs7uRirf2/TsAhFyVh9E+VUfl78hIHAhl1uoKy2FcyUDQpqvkxpULxrYKaRZdLldmw1H0EGvH3
i7WcjWkmbFUYX7econvvEzYriLgcmTk0Jlk4CbN9NWtyEa4LQ1JN3H0GJUatyoyIEjIiHujNEeac
qtogga3dEOo4GrAFf8KulAvS+CJB14DjYiQ0r7pivKu9BnwDNyzDwiZVN+MXQmeXspB7n6F42HRm
jh/Z2LzGTh+iorf/cAk120RNEu+OzmCxKS2q7AUweS9whVDL5qceeupSzUuiWXu0DOppnkK0MeGD
1k6PmcH8JDfCKcXHq0kK60KNSqH+q1g1HnwtQLjpKtOFwIuhKmmWWzxRch/LaHRQv/PX4Wqclo7z
J6lpSh13EKXAKdMUIdK+EwxQtq1mGFDUcJlbGKXnRIi2mkywOktfGH65uP79eWiNfX58cUZFBNqX
Pe5aE3skmJHWgAFPoRTj6iwYlzR1Mby4/Rr6uqyJDu4uQo7EPoJiE57TFRsVE4hFcsPqYBM2R6QT
0utFdoQgos7vuJVb5uPU4DLnZMLFuqlmxNDrYUyArobwUhkEpULvJi9UrDe7SvjQHMvWxLLCpe1f
iTII51p6DPnyW15fjOd8LNtyh4gWEPntNf6ckiZu53k7mvj5IEjZPfAGq2vxiFRvPybevs9Tahz3
tY3Hr9eGCjJQwbg3Gz8IEHFBkQRNq7+bM4HfKxVa8jq72EX4tYBVeRPLsLx7xoIgmb57rFhUi1W9
Z0rkKeS3aIXbFtO68WlE5D/DBotvea09f5jXD4t+0SbeO5BB+vhrTG+EVz73lovj/od4UPMi6Jqm
svG7A2rwC+Kxp0kr+TB6xpP7DIqecwyFa8zQYV4cSI+CZ61xsq5nUznpNEwiy1jq7PK8uPOlvELl
TaKACsmueg1yk4yTqt1Eu2vIWqaM3G3Yz5VHFzqsRUJ9QQM4Zy4afiEKvrcfQEG0zidvTE0PBU+V
bQhDk3ni6/acm+2auVXLGFgpgpCZ1/pwLABX+EhIIBJh5/y5sEVZ/A6pjID+PiEl8qRzDmSBZqHu
jCW8B/GQB7pJnA6Tm+AN8HcS2XBVl0mPfGD6QYCS9bN4pY40HlfEvRVwLzOy54rNVGN36vj/PYBR
U7z7vyKoxLRL9W8c9J9SF0/OYAOBjbt2CJjs2c/sT4VT20UoQOqbvj8xe7Udka99Of5Nm8y+qOEh
mJrEkHcegrNWel+LTUjDqub4Qk+RYk0DvjoM1hwfZFmJEVEQETBkYpOJ5dEVy0wnozmwX4JSe7Uf
WNl232Ts0hlpsFUvpi9/K61QlhLeGqT/fjErsYWjh9Utqetqf6SzAoDXiiRUPZHzZ/sz9UZYhGGO
/qyQLnBRwS0Irf7gLzzy6twpzrhWqRpxpGUkBcfW2leFao8W+FA0nAq3U6K+rCn3smoMaNIM2JdN
1eLU5HDI8gTCmiM7EifVvRvJXcwl9GCs4b3KiPKGscu+9B5u9LEKI9QwgApl9ypTZv+5yVCIw2QY
TITAbtLNNlmxWK5+DF8iFYRyKManuDpQ2Zi/lymaQ4ZlmKOcZxy7+AU2/8bxmtR6i3HanqtSm/LT
TeE8/wqDRz1Ypfh3Jhrd+K993I9qMSndBkOotdHphtFWW9nxJgO5nMEr19vTwEhOaQxskMelzg07
3cXMtUrRAW49SyZ5/QFCFHSPh8ZiqVWAsOm9sNxKQHmGv9cm3lmvk/O0iBmlKXzolqFFXeQ8FVmv
3PIq7W/GzVSW+erDfQbRzBF7QcmYH6oqRyz1+Cfe/YFyn26k5YWGUNluF8hQjFAettgj6bJ4Xn3A
mrXIUZq9n6nT+t4i5aJsWm9yovdAMuLB8t+i/DAYXZvq5effaAwMGmWo6Rk5dK/Cgf1Y5bi8tfcT
arKcZI++P3VLKwj4Y2K7nY1Q29t6ViuUA972gAJXqqqU+QqDvgZCwgkvmhW4UHCVFgxj861hPxNQ
LJuFdR0+X+3WhBbED1AAtnT2hRqnG/VgEEMPWMytscNMhxP8EqXuIR7CBEYoUOowV3QMcL73c17Z
sepTEAFVcxnbNFnC3Z4XqPTPcJdmgB/HwF3HAfA7OYp0hAvUmRnBALClBHRWn7wdBQkZ0vmFzmEY
Hmz7AqEXT2DBSotbnxqVVBrAl4EsYu/wgfn7AeBRcbi2oEPPML7awbd6lgPt1K0U8BXms5gz2Z1/
LhyhKNE17LzPdHODjGl4CAOQwa5DQD9rJNXXO+6AugQoaj8EdZ8aD1dJc8+j6ck317rhRI/gthmw
Tiw7ACWoHBCkFlhnJs0HKxS+qxTvQorcwI+W/qehO1QojdrJbXbH61wSgq6koqdXdMnKozLrFQNo
M4olg8hQYdOmZDKxD2Lwt5e3SGzyIt1zdG24AnjkCcq+EIi6ITm2nb9CriYWp3VN0BT8h1oAfxlk
y2W+2s8IxC0mEc5sCMaSEkskVDM9CO0hJLkDF8f2L9eStp1TYh5xvOiFjKrD7rWfLgbKFs4B/6pR
R/Cg9hzZkdYruP/zNF5swEk2aEnxSUqfA74b3UMAVPWMV6iwPuomTAsbIk/pr0XKgn0guiBLzdyN
O8g0jNLpSRBiV7dgLT/527sW4mma3ipb5S2TkWwLBmnVRmWVY26J/k/pyz14lRp3kxj1y0Esu/x6
QOY2gq6AEysmJ1hBS2R76X+HqhTQkebTSW4tosc6ttQVmHct58MoVxB5sLOnOCGB2NL+WwPrFCIx
Ce6T8nLJYqeI2F5nOsAOt0UFH9ntWg0TF6Ts5j5gehpzumZQqHqkL0LKXP1HugrHEcNG7OTOmYvC
VPnCsttFk4gNFH2ky5In
`pragma protect end_protected
