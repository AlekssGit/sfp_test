`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
Ga5IT02wHzk6fn2Daxihr4vUVO536Oc232Vv4kUsp1NzGXqoiuwyvM0le8V4UTg9
lg3UjdgE37N4lmcfx+8cXGOEK5FsSjCH0+hgo08N8DwpXDYotNFcgJyI9AbmW/MQ
hLZ7xtPeUBT+mJDtJPB+69X7LIZF/NgvTsZYKvIJaFU=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 36496), data_block
CNlfvxL1WNVUdDuMLdSSctZANEskiKxVKizwfjShcDsNCtheEeBOp+dlJx3tgraE
prtScZiuxC+P3n2gI+ICR65gGI9/OlEl+CWSKREnoQGjD7MiqsPtGw867ZjNvmCU
csztYG4JfFAz6ceFMfzEmJLjiAWm/9SJ3qD8iQPX40pLpmvVBHYf964T4GV1POT0
NX5KdJj6A97WS/u+VUKm18emZHoyh0Obt0Gc5VbisONYvuYGUYetAsc99KRopnNb
AIkKGwlRHmMOQzELkiK1FgBLUTg2OrotK5sQhyeSJhDgDUvg7dZKGkAVELEGpMIn
CXyjUTgCezCRs59gzLH11iSAPBw8PHiJkg4Dqpz4yGABctvecK0QUuRkTtA8qLrW
cZv2GJlx2hIANhlUYz5NZ4hh5ruXaggfa6ENBeYP5SUmLgn2Kp+Gac85DKI1tCbq
PKqUBa5VnfwKCKr9TGL0cGhbMmH1lyBtZilVtj8MGoti29c5tiU+cVIyly/Y/wTx
aIyIX+9NGScqVDyWi39AhzGi4MDRo3QSNbuwgD7J2ovf4Mp57rgTtvadtV44HLcM
2gb2AzUoQ4nLX2qyZwA4KIN0iDS8ndvhBUpLYQppKm7znneSjrhRQhx1afy7188t
6EE8zOudQvA2//u2oX3x09NAA1zXR+Jpjq6PMtl/yc7CHkalXiwv60sbyY67EBIs
kMFUrMeEjm/qR31DItJj3QZenoPaqkpZKkGwEEDajXXK4hT610exKf/8I0IOsavv
pnO+y8PwHyEivKJ3Roo+RSYHXPkzeCmXRmtAVFEMOSXQaJ59iWpqy1GRg2SBsybM
sLrwke5K2xnnbOhvr4/s+x/C7eBoItI8AzTxbuGoq4NMiqT4WC3jXx/1ziC4JZwF
oZ+V4WSlb/+I9JYxksAExI6QQiRX6r0052CIlEP3Zd37ulh2fyATlAA2r7lod2PU
/K81A79VhxHZJQ11pbAdSbyo/PF0KqpNhnRvEbdUiZaFQcsmOc7bgl8f0evEOqT3
wCimqRfDkSKkE+ZQ36QXqwLFY3RZtk0az+v4gXmRCTD/NMXWTVulReA/7i0sRojQ
YjOUuO7TXxA+RNhjTruwEza5a2XnPSIBeobWWTAUxCro9L5DAm/u7/vYtQYMLiKJ
A/0e7QWWqaLcI3x3wAy+scOnUplJsZdBQ/eQglyASCwDx61mKN2utmHb19/4g8U+
nuSO5UDdTwUNjGIVzX1t3JB51Fc8UDHXxincRRBbMNyF77yrIErOgfjq88SrTjqZ
zAA71hm52yTOaWZ7vktHZGVddOGm9A7ax8OT8WevBD0IYzu4AI9JIQITpv6McmcW
Z3ZeDuvhRYp9jKjGau4jSO+k6uh8M3HHL2v9wQDm5tdFsfOMzIcxpBd6zbwmi2AP
nJ8T69952IwMrx+RbXSal3JJfwPqIb5I/9Y1AVUdr5p8L4GpTQ+1XPqYYIY39+Jy
CwFboKkj7+UnboumUzxOhBaGDyJGZb8pvvq/LIhEbLqc64wzjpwBoDudvkrGCyE1
qhqfjGqnEB7ZlAPLYyFvKa86nsjSvCdDgxDhR5zYheh6qqqe0EC3TaDZX1LUzfup
sV38hrootO3+pvm6ul/0FVg2Wbx2R6JzrU50zLXaUHODkqloLn0pqhHKanRyMEeR
Hoga9etLVLxB+C/9V4Jye0ISsB61v2Qky5kb3PyQtwf2fGzJuobyk2hZWpVRhyqJ
S+ZDixGGK8z9UZOHEQOmkcJnUmYIGKBVasYve9UMqzIK3wWoKzUdEKNFKN9DvXhC
Y+0H5pJFi+k0E4s3lyqqitQPXbXeBnNbkV5n76RkdPzxr/AwQvBrdAvvOiFEoPix
KG+Uuzx7K7MPBYp8KQDDcbKwOg1HTyfSm06t7L3Z25LzvVe8MisXe5x98wXlCwSG
oZ1mJTflVhq5kwx1byzX+LiSref4194pxiDiyzaF6Gbxtkf5raX0i+cnWAPhYBpT
MbZS2libTC3YOY9JSx722JR1W3DR7kHf2va1ydctRyQGDvNMJGf5oJbTNBbiRvXX
/CSNKrNhJxlo5w8pIcZc5oJDF6WAoFhzbR3hIYPa87iwGmx1SUbFFBPARFJUJKC4
sTJnyj7ygR1PPbD87rU0WeVo+zOFxdmO3d7Tqwr0clO/8zenfV0TuOOCYNAW1iG3
mYc2MdBvKje9eDRSRuFWOp+K70O3OZnUbLxlKW7fFlcEcQ9X7Yvskj4e6cFjX/oB
4cidg3WwG5e3ALspK9nKYtkiZzmXtv8RwiVr+yplgrqN0t7cSyJ9vIL/Y4ZfGno3
jyeqBm2nUpSXS+UdWaeVhTuod1CB+0H58/NX+5UKfZm6O7xqtL4OBiQhC/S25kmb
yqZ20m9oqt3TdEjNTcxcxT/kMaGHvs7kxb16ImLHOGzFq8f3lctEjioffMRQIUPr
YBVniAWQqW3YCK4T2uQbmvFyuOa7FWpi9ypwxZfXNkkez5ZjU9ZY5Lhup8IyBsCf
SICsJF5FaCkhuIKTx3ofPX02Rj5PFJpy37E/qNShns2bI7i5yScKia5ZMmBZIxti
exI/EXT60ZX2Ty0rKm8mJE8Xrdzq1rqKC71UNloWwojSkPLICvoFlhmgETALOCQ+
sC67/kOmelyOgMQ31VO37DDb8LsDIe/Sh4Bf8T+QQoo9OEj6iN7FmM9NENyZVABD
v7OxX2HGJBQcrww6X2pjEboHhnOZfvgGXgNh82Q7IAiRygu5ZCOtD3tzFjvOc2fL
9pDqYbb4LqKKAbbk2wVGQWdgoW0bCOKkWE5jtT8XmpMc/mgrVCp6Gn74i99xu0SE
ftziDTfU03jQpwERTR/Uo9uN8kdYO/iiYz72oKi22OuvRKEyECFjMu59cs0dsDCw
3fUzfXInA9e1cLTeX+5HoYLrKiDAt6H97oboi6SRkNexcUQjV4TG+A72cUIarVwo
yjkxDJO7dgRbOo5dzMDJ6wBZCeKGuu5lUKDP1ukDj/OnGubFNpDW4ZNIeaoRRdja
C2ugcJxrXeZIHlPUhEQllfENHl3+SC4ZUjltbylUX45vHbb5V7uVH4Ly9enYYbPd
asuU3Grop4Dsk5c637OLmj7UlASnYmpDq5jgJ07PuQ6cf7HW9lPhTuLLBX+emePZ
eWQiR8+tX/1byqRafO4B23BXHkcuO6Jyb0n8HxVlyC47dHzh85frWNkWCODkbNwn
VzRvLNR8ha71VMP8/axTv3Ku2GtWDoUnDox7Yb8boN0ZAHdqEc5F+rnkx+kKYvat
6UDuabywHMBRZ2AmvH0Qv1z37Uh5lzQWGCGxZScf6ClBPhOB1S72g5XXGVzfFIC+
RawrDZqSF07QiXjMZ5Z5n/HoFEqzIfMMtipnNlBSC4k8ksHrvqZbfsmLys7KessZ
S6xCFlb3wQ6oUUqFGR9yjOktHUJRgqwAeSM81JaSlDL8v3udUX9YF91O/BJifYfY
kR0T75vWLvVFO7S5iv5T/NzlIBEyO/gOyy6rdihKJheHK3NM9p2uUvCdSE/TyV1z
e+tkIgK6liRwGBSVqGKdBkNQToEduHXyIiXihB9QCoLx3gZZZVVwCRpCd0rqIMUw
bkXwMLvLKoOFR1J31WmhHE7z4mGVuVAfbD/nNW3VFrGY+HdUUJMvE8dk4A49GsDW
vLZ+6RDHoGuaNzIom9st6Gxc/sJ9mC9eoFeQBQPX/6mFIydOxH/B7TmTKHrr1PVn
WmOq2O1pzP4oiPPqsdgHx5pUA9nrGH+PsN7+mCU66938MnHOLEwjLOwEHM69wbi8
yvy9SjBduaFnBoj0mtpqajMFYipc0BNXyuW8fCRI20g/0mXrMAaDwnIsGIRcJmHl
6nLuxn/jNiHoUibKNTPJwx0KrTUcl6jNOY1doZjtZ9NLoFss4drERhv3ze7WUACH
BvsZGX4oBoDEAhhhS9Iq73HUqIXP2lrONG41+HpsOD1qTb2SlzwCaYb9p3smsVdg
FHocK6QSZZXBjmTb4bHrD2SSTr0NXump9YM4ZBqynShDHT63ob1R0EC0kjwniljV
KD36ZKqpOcNWF4CrlmhtvgPH0uV6TEm4lzNxEOMt2fTlB3Pbe7TBRBgbcE+8kQ59
Kx8riGJ5gO+cPRaD495Cny7ZakwPDxJs2kO6eEaSWvx8MUwTWXd7jx8y9iAL6A2v
pMRHvEnPlvWjgKJ1MW4GKp3b0COdFMYHGcsBq9671IqScPDYNzLSgCckqUe4Vkc3
Zw7XeW0yO4kFKde7enHvAcRKKMvMkD/Xrx7oajAsWAB/CUolIxO+5CB/y5HAfZcn
VFTPS+rmZReLkYP1O4p4sRqT2mxtOhZG8dK9LFBFoRjvyq/CG9VUaIfzgFZomRze
zVTG2KcWMpsX/PsGmzCvXAjzZD3w+0JBligsK7nasvgHVpuqxKTHXpYhp3w4qoBy
0whvc65mcCYORKt18Gy95chfcFi3fX7kJabrQVhjD2rkD6YcWXNEKkLiUweEfXLN
gTHIFIqtSoAbZVkA+PPkgMr1zfhZ5JIYdaqDF3wRzvSqkAGEOIxv6A8AdpokBkE0
xdABebsY0W0wfyERdrD0Wy8/vBu6ZxRoAh9S/TRug7Dyu2bxQeBVntyqZDldCy3j
DKXLcnl6nDeEKqNiQG95bAiWGovNz1Y/uJtAEcksvwFVor43ukuIeoUwUmQYAVmQ
5EgWGMdjqkq/6orcawJAEHTWIlUBHmPdigNIKRDbD7X3et22QTaZJEqVZBwp9rUt
+6Bql+1yIGkYgyif2Ir/vJjXuWgpwDRR6gXKIaOt4EOFYue3ZhuEuPteIhFOhx7d
OkLaZlnxv7+QWrt8PYIcIwhdV9O6NgjK6DKXKggBSjM1hgqm7WJ0k3/VGSOmf3yb
YXG8F2VWXic6vodMGghJ8+66nXJFczgfDqdaaxhnQ8pOusBHT0kBIWQRqwxm9reB
nG1aze4RfEK9khaHNgH9WTGLoowrYOy4z7MQZv2VU2McMmIDt+/Xw8L958FItcOM
135ZZRce6vDRoVjV5Jd0B0r4Sm29CbrF1nRx1zRyjEqyM9ZQvepH30EmWa2B4AFZ
5Wz+1OQ51NFWh4AU6WFXnKqHyvRJR4CYFWsgMi4652E+LuGdrLKoAtFbZkdR2/Qx
Kd7H2LthzX9efb6qENp3XrkLmgD+WEWdC7Ze0KW05jY8WWfk4PMZsaa650ZFcbmq
2+tZw3vxco5/SRHueXQhEArK5NMKb5IGKklFXGJJXqAyjnv/Qs+GrMiqdlLcUC/g
L9OD7G2h04Ghh5DK3Xqij8rHZOolTM2aDtLTz6kMYkuYR1wQmKr4FNIrzmUhmDF5
82t3gWKhOshi5MH1KVHn7mw2QvFqy5A9m0v3n57TMMktLvcHuYqLmcfLPh1J30pm
sywRTV/40OcnA6FlbculpDEen+1QNou0RTYtPeQMlyWtSvwooIHqrmH+z1nbPF/V
IPK9PEEuhCx/RD8Q8PdqIV4BEmb4V3iUh7Wvd1VQP+6F7RF8TDMxgBwhDSUxQ8AK
ITFFbq/YFSeahYDvY39LeXm0HneO7WOUag+8j8t9776qtmk127RD8tT7qHrtqfmo
l8vevdfm90PptQdwu6jXrFC+BVNVrSqAC18fJ29lPLGw0DthzvDdEaxcAjqmp31c
uwyVu52kvDS0YDKLEniT5BUBNp9YT1wgGdj8ZFgmz7lwR7SUXQDEwHV0SIeq+Zey
xczVYO0R0Nr9FnBE74EBa5LoUZAFmr39ebCJkuWV+RSMBu8xGq9OvA04gFZhbpK8
8Gmnk93FPNF/l9eOXR2R539xKCYjradtQfnhXeu3Wq6O1fAPFnEijyg96RmZ33Bo
wrmnkUeO0P6tuEXZYdhW2jMuGX5Z2bubQDFZmdQ5xEdZq/cOiYlF513ueHCf6nH8
c7zB0Ewt5S1J0lfaXSQc5kfKoNORcv4eTPDtdYPd/yK6tFUFkrfBOIGDARZ7ZahC
rowMZ54xQBiRYNmFeGa+RarjY5VByD7ocGUyuCezXIiH6j79KLxPHA6Hh3+pehsU
u93AGsTiapxAQZ9fDLduFZbLxWf/4kC4438uaXHTlujImHnG6gkAQbJlwhmHBhqR
jIgHBPmL3tkzm+t7z4VNogct56prbRbk5zM80Fty2yZQOKCxfE2F4OH9oBWZuVvc
+yGBWSDORIMmvrVQwc7UYML0PBsimyoKX+LexrBpct87CkcRRpX1LU13vAPtiLlX
iNwKcl67uFMhnRXXFS6UfNcLbfjD4npW6O/nyG20TRokcxZOIdLPzSKG3x/imWNs
tDTUJE6yqlp4+0Jpl9GFZ980n3fEPvOrNUaqIvIc4dAvjFiKm6W4c/C+HxF+u0wo
LGr776WeRSFN+WmhjdL/ypKeK1Optn0GqtN5zDloqBPUtT1efATWKFzRiIfEs4zH
FhivjC9tabQuwbFcWKq8D27J7zUJTmMP8q/bXsTNSYlTtDmco1wdsF1IDbC2WN1K
KRqq7R9tHxnn/c69V4/9mfTmnxpVT7L6iKJWZccyq7kvuc/0mAhjeuRuoeqWUOKz
OShLUpzRaqStFiIO44+/qF9JwfrnRv+zYoyQ2XTWFLSJk0Y8moBvcF6E6Cu9xxVs
1PrzapHXLly3oa8Oon36gYDuoB/GkohCXgIneEo+5fIWMOdDwgfk2vTqdyt+APlX
PtOpnzg11+3kJC795+1EUGI9v8lUPF/4/TzVSgQMEq1XeIr/AIyaTFCbp8IJm1/2
CxeSr5bLcMsJ6fRDh6j6MCTygHQe0JwxjayjNQB8+Ep5IvdHS/Y8TDEtzqBrLYiu
j5LBRcE/GbGiqBM9oRJ13+uSkoN/uQD6mDEV/gKaW/a/6J0LeREowdmC+aUoL0Tk
rQJs95x5mCM8mrqcs4RpKpRbQYUNRH/pQ+cfEcyRhxJ8eP4J5OmKmB9jtloSjxGf
Ppm234rBBS27QzxNkesEb+C7/k//WL82oH6gJKJKfTK0kgFz41PUvwo6OpmzV5Fe
NWJ1oCqnpGPcwQNGnckd+c9UUrTxN8u0gcKrqVLFmOVMDTNFGnoOAuDtwhOlfW8p
Pgw3DbpVKlD4WJBqbAdlwUM8lU6v/ox2pIzWN8nQTFZfbBZHoKW42ZNP/LodYhwg
HDLcLDuq6D/Iivs33M4/QgymJCElbnAVNqMVBjal0HiAyALK5f3rBEjz5y1HCWjB
jHO1hg/XRlBuUtypxRoW33ehUp/hVwy8yecSRkOncP/1cFjFbaJy49JWIwFq+crG
YG/JRionCoOr+TXXwffEI+Ndp5qrNcvqxAoRSl+Vx7C01DTGhVTq9c264MwdYsga
ZX29o2b4TYIvYn2vwSt9YBaiRx6dr/nmoxbD2P6+Y1hQ7vbzPWyhFFObe25Yl0oY
Cas7T2ktr6ZQnOawWiS2EgVa6W/UmcQAEMI8yv73gAT73od9sG638MTzNIt4TWBD
URjYfg0WPTCHHenwXegxOf3IlVVsZiSJLxZyN7vJwwi54OsysNf5ME1YCUa6MMga
EaVf+ovxXR1ngICzwSrE58ZJpDZjFbNRCSNs1MJWQlCo6ohoRz0MV5XcwefV48ta
7VTFK6hWoiq131F4D/jarCJLHvdL6mT8Yak5I8gPzKplfGb04bucVSaf0RF//Jsg
4IHJ1s2Dt712jjBL3jl4hr4mXJG8jNr67836YjIR9fzgQoR/dNy2ioBOZirz0yYq
+heJXLcNYtzFqwzYbR7u/wZmyvBDdq9yvTErKKcFcQMAGmrBWqLJGkIA765DsZ0y
nE1Y/Tgo5mefkXlt2ji+DgC6JbXM8U/ZizMdwxpAMNuOQ77xxmPlxnvozpuTPg0+
4KX7HpKZCFoQay8yZBpn5Vov75wNoKKVNWkFl2rVXS1Dq6QoTymALt8a0Qi2i4G/
d5R5E34FJrEXOv/a8IO8/cW2AOI1tHKPtPS2kamOQz818k0SwnW+P/gQjxHm2uCv
CnxpwjOqzUyK+pgYqj0vrlw07VC/rDr+IKMqECnkEzrryFLuBHgTrVjpNOvD5txw
Nv/ew6AMiO3ZKQJXsVBsd6dGsxBi9Qi7BehVQ8t+UTOfzHz2AjSk4BO24UiI53X7
ljSyaHJT+dXO0Yx+arajNwmZ2ASC9929R5U8cGAK7vCf7hAeh+i1gXFK2uwDvZrz
JX9ACV3V+2anio6g4rMMui96xzDJ32AHnOnY5O2ORnP0HwyB7AT8K+bkJc9HW8k1
AgS737PsGHLBam6kpjLbPuwEy8meFtO/9hTxwTWHBScloEBBEnIVAW0yqlIZQtgo
/FiUYk044r6IQxI1ymaGJaevzSup7OC2ynHG5tMapNhTupYdPPPuOaUgGcqq9Pp8
jdLmssuYr/EuR0yYo6IB/aAzCanudzHFYrrwv/MBZIv8PLLrUkQ6563gwK4AuLXa
aSnaMbXzXo1/31n6cKohBYfFJpNlOcZ4ux4tM58z9UfSV+kNW+xDf+8bJv0H94Uv
hrmXV5rklB2UIiMtP+O/UxnOxA0OGslsgmJHeqmos+MpngVDPIHvfsCLAQOgzl+k
b307UPeGulE83JQH01Hf7+0ZJFotkWb7vmfKhuXJq4G2jkqaxOY5O0YwykvEGjpo
hGVWTtxYEI1aQV8vssVlHgccYvF0ZjCFMf7KuKbxw4fy3lUSVAdq5j+8q5CjhFxm
dPN0BhlyghGEk078FJTTM9l+7gCKksCE8Ulh7QqBKPST4tJ8RVvlwTqj4jDxmmL9
UaGHJUZ+GcYaXvNqGpWUf3OS5gGrI+5h/xzpIwTNiawF0Po/VP0wUfI5KbAyXEBi
bV810GvspKnHUS0tXDa41I+kQh/HBy0o/nAc0/TFGj+Atf4uxYKbc+tFhBTSk9yU
xczJh7rxpnU46e+t2NPlgmlyPY5RRuB86qUkdtdJqsuYTS0MNwHKRBpBUioN/ZYK
GCXRNcP+4V1hKYDw1zBRhJf1oi3LnKvfHfQS/eFW20IRsmpRr0mvJx3Zjly1mFZ6
cTmazL8r+awAMwhePnn7761YneYNys1kXMsJNT9m+YW0pkU9fQ42xJyAMlfxxSl7
3qyjuIVtbnj46qgXhkaGUXwiU/ykC1R3NoZLyNJD6UowRWYwXmegS2U1pOXZsOir
lwxqnpk0F7AhWBJPUr0lHG6nm/AA9WQBDTm3htZ3/LwBDIcWLqEheNz/GU5U6nww
aSLh+MYX0aNWt5nrgRmftmoHg630C6o1pBIG8ZuIJ9SHNoJPtC6VR3g8lrausp0P
FUV/9qaWksY9se8m2cltCFWcMb68LY7H/Eejk4i5vSzJVYAz6AfjzxU/B87jz/Kr
7qFcIlrl9fn/ntEnFYUf4rU359o1eCrV8aSX5tjjngkapbzMQHpeT+rehHCYzWqR
DNsctvITKFTkcgAFKc78aVDWU4I6jRZQ0VTWSD5/s5YY1uLzYL3CPRDozlBjxQWa
NVIcaki25qQj0q3RWtVi0VmZfTeB+youv/y+5Ot0bQieWxbl+V3Ry+M2aKG585+T
8WQdCRBDZ5ErjB6nL3Q/PTTo6J3inBj1FgKh1OGrx363MS7PUtv0DYaRKvuMZUN9
FbN535jn9tr1v0mGYIQX63sD/OQ0rJqhVw9CKMEXkPiAg42YG7UQ556YL5MBF87V
RUppz5Tj4XH01gPKcq2s69okziy8ijmAyB4cQoab9PLtzaJiC6wd4xqfCcNvYD4+
a7YYdk9I/7bAvYDoagk9auDulgONNvbZhhTPE/TcTk0EOsTwLBvuk7tRB2ZBLrug
Zkpbiad4+CAYD/dHy75jzKwg0JdGjeGqAiiTRzwNBdKG2WYGMiMcH+pWKLDxYDvA
1bRK828EHU/xG+r7WmjdJCgqN+W2z4Zjk4yJ7UbT6I356zchxlpbxD1xoekIW82d
Z+sjlFe53iavvjGfs+qwegxGRfm0oHOgdsvKRDtOq+M7Frg67PZRF+kizVy0n9rp
QS0bkQFIkf8a0F/feaOpEHxLD52KxxFEMI0rUQ+70rZiIy7F86OKPn/vjCpnsVph
gWWJcRnheWyeZsIsiYDeeMVT67PQt8iWO3J/Gr9RjYGUPsU01RG8f32tXY7bt8PQ
JOUUWvg18p9T3bR+XewkcByYtuY7oUhwFX1VHMkXJIYrTdDTbeGWnTazS5d7k9HI
w2H1Hpmin0NxNgMDopzxipK8117bGqIV7P78s8arQTI/j3OuykTwUw9W2yX8ybWL
7CnyA8Fduo+JrmqfpZG/+E44FNWRbjjfCePmx+pl0or4LC/O9Vd/lnQqY3V+mB4B
GfRIz5t1OATO7pjspQrYAdO2QVOmcfy6rn721zsFuX33M7dZL5RFOvU6RFudHwQW
KtknYErP5Z/O/4vV06nJMCjbXx+DjrKkDNAAEq38Z9rsveV1m4Ejg8JSkermifIA
nEyyy9mnpre//cbC/FTZb5Rc1HDWn0CpYVBJvf411XyYwc2wKFfJlRw093iGt9Wq
Wau3HQPQuA5/cIzA5tWp7mW5l5bnsEdGpNz1bnRH0Rc0Jyc32BTfiNR3eKgGo395
vbKbGWbWYPqm615Hfohh0HEo8reg7fbgmaJcvK/erqDveGK7Ty3Jt8xCayOYSuX2
nz/8IFcmt5ZptPTx8HkP1rOsUAYZdEDw7A6ei5lDFrXZOx8czq0B4vwvQhAbZ+y4
0xbkbpqEwZm/YeZN/oq4/j1XG8xtRm3qaIWfkE8llX9p+XyxC08OznNTYbVNKcSN
zgm9eug362W1OHpIZRQ16xivQt5tB7hf7RVddG7Pz5UYyeDzphwz55xkD9ME/kpW
tPdfnGKiu9bzNYFXsJOlII+k0EGVgRY7cvZdi7WH7qKm/kLEmBvx/21ugu0a7P6D
4VJOUrVZGcG8iVLsrhHQEPnc7UDzKRjV+8Nx8D4/DOCuFxqCNc4qzzqXpS6G4/gm
MvFLhPwI0J4/inYmgWRcsFC8/XnUSbcuS8c+e+OsBp073Ngm7k+QQCdNx8SBSMQi
H5GXJBCvxHDkgQX7ras1Eamx+LROou3etj68L5JPTXq4OCiRR+szu/K9aeiJUTdX
Uh2sJnB8FA6LUd0tJdhAa0nF3rRytC19vS+CLv6tM+Mm+AXWPYEEuawRFwl4T1MW
sivwZAnHjMDJg6XI2FCaFWRKexOW4/X2b4YWRstCMkxaMY1v9K8YLud/IPHW7pJg
p1Ub7N8agxTQJqpwEPgIdUtdGqxjUBZ/fLoikPnWVOB+wZUUgVm7p9nZlIB7hUyA
UOAv5POxsRymA/JapcZOR3mc2fJ4ncgYKvU7wJwzmM10Azztx34PauxriNXO3OPO
wtKQqegbnm5HRxjVBrefgAdK5XY379YtSbGO/bFuK81WtH7wFWnLWUrWQmkbJI/Z
AFXiPhmPDYTIGx+APVQ/SBzcGtRWLYA/OmA3m5oydrnGqB1pLvMdaIWav8QqDdn/
pT3QBk70SOqnuttFvjYUJmM/BUarFYhqkLNUh1prH6qJYr47vCAOtefSAx1F9Y++
P9IEnMguJrZp9AjOYyAZa35SQwfv7FHrX7cAkXEtx37zIvaVYg2X3VTPBPYZn5Ou
dusU136sJMTlbqkhmBdC7cbFcWDnRCCb8/mMs6cecMF2ogaBHvC9uG0ImlbgZMLo
pVAeuxk+ncr+Y5QvdufLlf5J6PXXzY1xsifZsd2qw584FfaB63mf1RCaosBVMFco
ERlGu8Co38oE44TkCEDZ4frDYFmixDpqmPy47YnbFhtXBG17dcRkgpqpOCQF+oU3
yco0xU8xSOBw32QwBpav2o5eGnQuhCYAaWkEkiVrCkLgyX8isj42yDQ7lmWDtsf/
ccLl6Hzqz+HpGpxg6ioyWUtHsJm4jQYD+IVcDyrolijuGC3fwGSpEvonSTAipsaK
n2nBn71Tu7s6+4TkY4Jkl7Oi8nXOmnQIAmn40LmmTa6BiZnRO+fX/mMv+vYgn7hH
MgzzlEbRHjGz9UFT0l+rnONS+wn94eZm6X7NPubfensIJhONiro8d0KdqVWMQpG8
ARnSlpzDK660buxqioCMtfBOToYz+DSyOQ2lZAFUXys9lWFwqXW0k1nu8q/tZTbf
KfILsCixpLHaZ+zI7HUf0VoTBiWKAbLtdi2gu+wP5P0EzLuSjzAw6I9UqEx42zdW
TOOZJki7Usbko1DcxfoN1b67g1j4mrCF9XmkYKPcasT8xgZG1LY9+Xd4iSabOS6K
PVKPlGIL5sLzElF1F5sBQ2szB8zpbVxVflIZI2pTq4QrJf/MuhMZUTMa5Jg3Myqv
YSmpzGz+oNY8mdWw5W26f1+2Kz2L+ZjfHB4esos8tENo+Tn5HArKRIsdwM3QqCVU
1QeL0cWye3yQCTwcPuaxicm+z+VDA230IM6gnfTOHmc3pREnzb+E6+Uh09gagyNB
GLEczrW26JEvWDjQg+QUYMlSJVXvt1YyZuJg5KeZqEH7VbQ8Pgm1ObBM60EhGXBb
+fmKapK8wxm0eGNZBMmMnZNiBLVrAu+ru/3qMGAYUmfdra8XyOvLbWBGM7KSOWYV
dG4kY6spOV18K/I2Ze+4qpgBKavSqarSvke0vVtTkfkkOM0+W5axBlTWjr1uMInD
8Nb9ERC2u9FI/2zZDM+/ZVw3Q0xiPToJgeG7yYSdgo9YmOj9c7VpdJP6jV5XA1tv
52PaWN75IR5dSMgL0ih3VDK7ZNgFIo7pjGRQNGScKyZbnOyVmezfrlk3vhBn+Nb6
GuGonxyJAEypgvOxo25OMROoSvZMV8TxExuaYtlqVn7RqzNQzV3y7qtHiRp8jWgl
M0zalzZ556nBRcqX0YegsXJNmLrTwLwaw44bk7GMXAB4v5Kxt6v0kWWdrDUqEaue
GGceINqOisWggRBuEtgZWYWqU4wXZ4i569lDSXstWdnTtyQNlrZE5tuCulVHzzZ9
Zm08kF1ZQDyakzpVc1CYpdZbWsqHRjJDjHRvSANwm/dsk+KFNCP4LtMOzjalCgTJ
RGHHBnhxC5Zufe0yUCqCVIFuQRXlUcR8s5WWn7kxodKjm0DiC1i2r/R7d4Yn1q/f
MwrRGiE7ZfbNvxL9h3VAAdor2VM3vRTbgC6He2yaQK7OQWh/ni2TWQYUq71rv4kI
ksxu6o1uonhVmTkpxytw7Yl7lYU5gplv+tMuZQBlFI1zGObZvutpEf+3pnkXY3TU
G3jSNftv69tj4vvaQ1QWf4huAkckcpbAzwQ7roEzMwSktInsqPKiz2mcXns033fM
cYufz71PbpqQWt9ZfjvGPlteTdB4iGkP3l83UKaN50iwaPlf7+fxC5iOfj1j2nDD
QVVRw+fhVWvFZDvYDHffJsWk5EjXYR2qIXA/4yWWa0br14Ci8PdH96judiqG7MVD
COben1O/IpQ1CVaWOhKYGWzG3/OtUfRRejnrwHcRR+yRo3KOU57ZteXsp2JPvTfe
EEydt/XDF+/439y30YekvWDd7eYFQq0e2NmphTX+O2LONrfJ/XqRQZKw42QyTwj/
Ly487uynONYZ3mT1VAj9aVrDaBdWUb2hh49Lb5dEn7UiR7nQgkclQ3F5AjlU7/Jw
N9aNSShqPX/V6iHerZHdxXK5snUHVW14QEHqDAoPAC9ZJQmu9tQO7xIlb9iCcPtw
f1gPcyZEI5HWw5A+Mbgq6cbVYBO4i2ea9GFoKL1djc47anYAqm5Kq8Vd9Vzv4wZA
LNjipxUATK2+sp1bacnHKbdYRBe9BQ/k639LZ6iJ0bqrs3n+gZwNx5fdfpwCMuNy
BFzU61sDN9GY/iHsM0x/PD90uApmI2ch5e3whLcaDC5nFf0JY7g5xS8gCN+8ezDu
u+9UHd6D1hNb6Q7EOy1lRivL3Q2ppXaT+VAXulkW1Wl9fqGK5rSRIHELB803j/Vj
JGnOpst+GYRmoWBRGgyk/mAOwgzaCea4+8YGFUGBYarGrr5xH90ZkVtdSZuDdf8D
9EVaoPuMtkXop05FjOXwGhwcmrN8UMCYPE56p11XbPlv/gz8UE7IfY3Ph1bpYvZc
VEVIdQuIGACer5YruvOwIJb+g3ZFXJyg9hvW8KOidDOsDeljHXxH0Hvv2gNFmVx4
3ZnUvV1MXRpTs8oFAbJWUlKpo573/3KLC48ly3ddpGtsCPQMmXWxUY78JdJVygg3
jtaKXzQey0YYU1RRNeeU9o5eGaAHCBPUt3UKmto1qQ9ZzS84JTeoMteUZjuOUs2j
D2mdYgOqnMrME5zC951jwlIxeqgU1M8ysGu5DcuzPMy/Evi3nnCcmxOlain2SsWZ
65hWhw4GOYet04yhnpsYAZnasl5W16UHTkFrmbmzDr/yC7BG0n96Jh+tO7QO/zO2
5NrtMOTYDNbNWUT7/fzL+1GNXFugfZHvSRczw5eiagxLiRN/ibfKXKTzlx+lyT6p
uZBaP/DO/liL3hDQ4fTknckIUgu3SMSj4jfBfZrFezGxzDfi8hwcgZTyvwvbdoS5
CKuiPlKJHmurL6VO/87pO+cNobs8s9G8dr4ffTzcqsTzbb2nVGupcTc0/hBbX+7C
o6ImeWVF1tqme17wX3zIAlc1V/smOWpEyEbAC33RbhJAtZZJIrQR/Evkmyme/DW6
5rNN8YKRyWPj5RjagmziEpOgtBmgcgKsDOnzvmEBCJ9qIswZn/p5ZZ2G3Muv+kDq
hRdmDobx1Kdouv/sy71jnTZvnuMVbJ/Q4E5vfOg0DWlF26wsHQYolxsw3JyObc9k
TRJInIvXW8wYpRl1VfxGJXXxBea/RmWsjhGOgKD7wKGOQvHiQcVOVw39IYGdNKOF
ZDGqq6+9TXEiN3tHEHb5WdShL+px9ZeMX+8GpyArSGY6R7rFidvwDtgIHtIZ1aVJ
9I+SrkDay9+yTinux4imy/BbVNTPlVyU+UWSKUjmQmYme14MdWIrILMkOsbFfPsj
QlsPGtV7eBWa/nX8WHJ7Vb/iQyXmgTZlfaU4ZHumLdA5DN8jo3zfvf3jPlYDZkGp
4SfZRedfOM09LxfM4GMw28/foap5VKdIOSzDg1JaJDk/xrZmgqcgXDjVFl1msdk6
HT/MLdPuuabmR9uPlYLk4lhCmLfJIClJfDPSKqxvUI8GaIcuFAcWAWJAZgbjyC52
ru19nXTUXzFGM9Ki7rovKYROMwm7+RuXBSfVxdHZGfp/NXyuIumrQbzRrLDnhe8e
g0lHsqz4iX9pEco7jRyobH4Z+RfvqzQrcu4eu78FeBONtOW2PAWiVZZ4AdKTzNQf
Wg3lIgT1svY7+ldbQg0f9CTyv/erDCV34oQPFUG3tYUJc+AuMzTdWh+ySdUks6p9
8Z6nMwa4SB95zXHJ1Wve4Iaia728Y0AyTtfD4rmfrfIayrRV1pK3GOynthI4TeFM
tcWyVovmftfea4vZxzPEgLgE+DEpxIKPViUnEP6ouIbipdESFoKCSzPRXPikh8v2
+1vnaGCrLskvkUnN0lGWvmv7qb5YLqvQM88bdsqJbUyf0utTbxPCcyVr8spFYs05
31FIVNVl2Pd9Ee1NGp0K11N7K/eU+DiL3joVP2G99Qg6Ed5xKQfOKzndhbZCjpAh
mKR42ZaBpsdk1HflitUjtIUqJoncr4RAkaXbxES5FsRJbOA2XW3zxHhz60atkKGx
5F9Ts3jpdFwY8tPJ7m4ijGPdf+fGo+OeMFK+8+c1tAMOdW1n0edLV2eIniPsP3gp
rgemd+WgtD/nQlwrydpMgrOtQalcQZ6apTeWOsROP3dc4SXC5qGRcHAG2/VPH7nD
ygBm8diLsh4zyiDxc1jqs2qlyr5lbM3BmeFREZ+BTMPjjUqvgr80a9OLw6j18BoY
y8JTTGSfnP/1MrtiN8n7CWGzjUN5+kHDgtPEJwta1hEuZ67JcNro1XZVX+NpSsb1
XulgSdSIef/1mcmN4jCgQWJ8QSufX6ZZhxiDMZsFLyCCjss/upSG8QWiLb0CpIO5
7JSu6YXA2QSKVTkWlt20x5XkFn+WKOb7M1lYGH8NMfWraGT2+obhRo8T/JeLiSE7
OzrG5ym7B13KCcm/ceD+QpoKwGEOhhhCUoes+VsXd3fe191wjur8blUAKED0apSl
fm7aE8bHuH7q6wIXxtMIY0bK/igtSrkCauGbjP/rhHHmm6lu9BgMHsd+bfXJFyND
x4jpkyLR9BReMy27T/3gxTpLhxHjadLRMDDGEYp/raA1OHqBiqJ+lmw7yg4O9PZe
KHB7aTrY7MPUgjFaAC0wxsYmgFZKjS0OYZng9K20ffVBW7Aldi2lA7GR3qN/2vtd
2wrPBQE9F1BDa57Obn1Z/zYeLqBoGLPu2ZLwbigsUcwoRxF4+/oNJBVitu+VxgPN
eQZxc23K3bRHujvkkp4FbxXb9hb6Wbzimm0tfln45O7Jb6x5v/1jYBwnZLJjAYhL
DaJc40tq88mCXEAZ0qpxBvwU65FGP5JA5opd5Rdtd12FVoECco66HWgSR4h7N/7v
jw/yfwSrMfQUI4w00/lC+V7o5K5zudLjdIQqUXfiUHCceJpEzV2aPKZeoEoDk/3+
hO/6T0ibeQhCRmlX4Dc+4TqseyKn6d3DUJcL+99CqFdq09i13H6WRWo/RJML5D1f
uHZN0kGxTf1BejyvVlgMMkRJAj82jdBqJzZXw0Ym9L2TwSJr6Upn6dNG2wzMCTN2
rJWeh21aE8smMt35WIkIpx9Iml72C+AkaCkiULgUlpBgZWoMmp601z6/7Xqi5T6/
nC6VQ8ty2V7Eax+GWEzM99UWM4IuwgIrD1ED76+LL1knBYDBd90k0en+dOZEWP5Z
CoXstYAgZjd+WBu6q/tvvQcB9tH76VwX4oTRheUqeGOgzGDjhGImMBShk0WzHW1c
FXYoPZFmS8au0wN8Rxuwlq696bEH12tyHgW+q7oEHB9bLDcP5njc+oDgsGtLv+cl
qB5pzvUGUmnqhSJEzqffWnTNh/HPF/K4hItuAsdIv/EKTu5OZ2N7YwH2QrnYSq45
TjYACsO1rRhXV82j9fS8ljuaEAG/XhnQ1xPiEPjZ2YLt7LO1MPpM9OZMT37s/3Pa
VXpO/1l55hsmDXJLaPI2IXCg2++freIHbHD8rYWNy/e1x0iAfh699Yfx+FpPCgeR
HCUvELVdghJyCwvpVZKj5ZYaoNk5Dd3+kr0/B8u4rJ930DfWNJ+fsHaw0TvImtPa
SBLxCs0F0C7dn8x6ILc+hTl5iqhVzvfM3TWnn5R370v+kHXg9cbuVutob7fFpQ24
+PSgdumnY3DK/zKH5QSCo/TVW/cFor3+C9rE9AgJNFINfO97I0kOKcIWoCTrGYao
dgN4/7XzFfc/Y0082pnsl1V5bdUFpitwKvhTsY4x1k951Zt1ePCxh2FFB/CXAYo5
SbQeXsrJs/p/zd1xt9MWi8DOA0KZFCL4Pi6+BRva6m3fF6vl2ZA0xxSjCD6bwpsu
nILGb/ss0s9XatOLDndXxawf7JON3GSVCxlwFvZjIwXPvOS3eG1mxuAfn32dfZyy
db8vJZzLnfPFzDCqeho66XFVxOKXk33KbkUfEs8xb5Om+vlObcWcp2Ac1oE3LyaR
5afpqH2NdO9EXZ0OH1Pc0zZsagOqxFSq74PNzCdLCom9T3IVCN/xf/GyJKiSdUMO
5V0KPpqdsX6HgGYYYWiHZQyXROMc7cVBVARxIwp9Sqxihq90uK20UqkBzzDE4Rmh
1vMUVH6Vl+i2wzGjP1wXZgs1p3iEdiaJh6u9DV3T94ayzVirVG0mJ00faVlrMLz6
UOzZSHZMN6lA/L98rHxDUllehUBCLjreh83qxs+hBJ3JyrvzWxXAIEFQg7gPISrg
J0MGmZCk4D9q17CoMDu4nY8rqKlYLOGGw62vZ44n0nr6+XTWJHD7Ku68WxBsZq/c
QL7ObRMqbOffK7V8j4eqKxTsDTj5c+Ch9u3DrqdBXdCV/vdxX7hrtNsUchAFjt9V
aQNUWtK97bsG5ZmMpu+RIITbNdx2Huaa0loWRAmN44sDYdxLsLq1pF3e0iEZTfxu
C2nhOTxqlGIZkNiXFFHUUtEvbSrPijmU3AZAVUgtrd31BShnR7U8s7RUIYHo0nrB
Hrrkx6V+V2y4Sz3nImPV38S9Pdv/ucgiTA2XNAtVI+dYNz2CClBZGy+aRy5xvniN
UeKnMeDKLyIe4B/IxRkYhj5oPv6wFZ88I1w74SJLL+RFgNkxWGOeFwygExzWgVg6
Sq4oJ9xOWPe5TOa5zY9i4L+SfHP6PfPesS4FxmfBk6NIrx8L9FDANNzU34DjbJOZ
pKBw6IKi/I6n9OyYqOohTj3JeXPL+YDP2eSA17Rmo5ArG9J9GjObgpQDpRswC7jr
ff5a84/NoRf9yw9m7+qHrnIve7ScpXo4qXZwis4kqWguk1K0zvyiYIVx8LSarZtZ
4PxRNulRWHzAU5DcMT01Nl1bOazI/rCaUgK00SexBvVEINWIB3aWUtWQjLguW6R2
ygqdFmI6+2pML/5n13h+QTo9cBrOvOX84dT2Gg+Ve4a3h7a8V3aUj+V7vmqbTMfh
1CoI88PfMpI+iF3Zz8IBOSmMnhH4Xndl4qMErtVwkCzm74nHpZHaIw3rcY+K7eCa
lNJIO/ZzQrFmN0VtFvr0KARxK0xEcndC4hE9wn0qD5jBUbzYd7mawieKFMufYzct
BswW9obqoFl2SPNdbeIjgHtO31S+6HS8lZwVyd9B9XIU1lYG3z8VXAUkrxyrcms8
8OTW7gvGZNyfC6nTbDb17ZPcCiuqYKMzSENoK8OJ3MMEWHQ8529rtDmBUSGvo1Qx
ZV/nUZQweLloafqVZEvJkubI6sbKatiBjeHIxb7r9CdVV2qYv1pTQqqOHLL7SgLM
IRLKPv82vWJaI0ly0Ysqh/fR5xvgWrpaSC38T3o2cR1hFOc3MFA2WQ+9aemhAxdF
1wShbNpjeSwcQz+cKYyRie8tfkU8HR6xj/UOdupPLMp0lZUroRcvVVxpY2fEoj7Q
ZOqNuALNopQR4GSmgPF35gPj2U1wa7FgP6Wzcoc5UOV/gvjCLB6tQS/97H2Y+8pM
FeI8jnDitnBXZNR7OKOQBseh4W7JJoEr0U2JMcb8kDe9U9nRUK3SFzuCQrXVw44C
JeyFfCSLbhS6RUXLxFYtAyjWfSXt63iCSvnYO6JUMYJvPSd8rsb/lCXj4AkCD8Tl
4Z1/KjOv1Vtuldq6Ujjg6SUNO7Qy4Aih05UIZ5rVg9JUQDoTrk8WcrqOmyea/wJU
9NKGX32u9AahlU0FeqWYrjkDl8fb/Y4OLHkn0qZzYlB2yvtZSHZz5Y32TYAbRiNk
s5WMgrpvqmt1UoRsSuO5PzGq755Pp5kIVvpqU86o6NnCChn+p7t5kzIdXqZHFt5O
m6qGlH5wNV6d9gdgPoLAybRaAL5y8wq5m3y7HBg0GOSAuWS5J0dMBMePw1c6Avfg
s1idyBzU7ZqWiDWcbE9ulg/L1i8Ua8OtRz9g7WTKLNRD0g3Z28LMJibyg/zAPG7r
8E1OJEF/ZGPj/d5LhTTEKW4Eq1vxPI/DzkdgUioGOuhI7yPwX9ZjsQvN6xUYKnA3
y4eTVKGhFuQyfDJeGR5vaD5Mdj1ng2kS9RkVKDibNZeOThaTTcdGNo0ivribkW+s
mnlb2ihFC26dqCm+ig7c6Q8l3qIw2gx4ndxAffjTuoiobSbmLhp24Kvxp1UXA9gM
NLsJCwcvnBs/wGfZpR1JlKOsL8P+wKYjf70qpfn3FpX7bOrkXGzMSdIxnqbnPYuM
8BsJOZlcimoPeS6yU3LcAMhWDrQTVWMMpJtLhvHrVvloJZ/MgqQPChfJn1kLjEcJ
Kg6gACtHbfGhP5/E78gsnZ/TqweEt34pLQTu/FZLCqZbbrpdVoomHegOJFRL5xb0
reu6LR1P+lCGhBPymUBpfqx7aaZ2OAC5bDTON01JHVmnt0iA0heKX2dCgZxWIfmZ
jZtQogF9+Qof2owZd3cPLUSxctiKhlAgdUd2mVqb6SaM4k0w6ajmC0bYLY1hQi8Y
wJErwkhKyubAmPLof/ay2VsSXoxlV2egW2EpQsyNkNVDxsZEnw5THZ4KpvCTn4J1
p6cpvQyd2qTO9vaKE72ujjQ/9dUWjPVFnGnL0pcn2Nw5DKjit10RZfdYIVWsCphE
pJWtzPat8EyQpMVaQ+Gm11F0K1mhPMVDDEnP40VSNYrZOnYQp9FIpna8d4QjVKD2
kCZHdjG47H1qMw08yHuVmLGy18UuI5gc8M6Qt/I59L7je5ZcuqTCAf0+pe45v+nt
ZFqGKSaB5LnN8Ah5szg/5+PYV/S3727QoMOAfYT3LERkPEIpaKlO7Xg+iYk5FHn+
NN1lXk6bhwz37LC88Asylx5NnP8S1tWpZi66UhU/hL19kU2mm6ZdzQI745838jGr
XWxsP44EB2uCiM8z94iV42SqEem9/8RU/fBdoSsO8mm3Ys7LNtMZ+L8wPiZcGe/v
F+1cwQTPv+Zr7InV1AS2acbGWZ4Wv2yVrkum+xmvypHGufIkjibQvub9QEsghN0e
tnDpY86t8MXH2JE0zNAlApuMsCQSA9LJoHKpX+H/HK8mu3oLCKMJY/MOeRbHh5/0
xXlvKtoqY/EUucwhtP62rxK6sBeYXufZ14Z5HABf630gb1h19eu9mjE53hXTNlNV
M36hazyAjyy1BO6NQjINug1z3wEjhGHnGmcydsaSXQ+edAJnAfolLKnF9wkioMFe
mT71Drp/aBcUmi645dExbEb8IXWCUa3EJb4sWUFhcb6c1CzOaifra+wW7nJHWquA
XRM056cZywHg7sswxq1Ar0CpnajtQoy9244Oyh2n2xLjMwKQFHaYRZc6GVRm3xVW
aYcZxg3gwVydWxIcQY31Q4WfFWJvL1sMYjn1ZDs5DepLwRvVg4AWzjgAOsZ0lwM3
JdIGlOd47ddahFi9MYdVFWpHcjagCQFWEVo+PZI4ASTypU1CH5mTtt3/qw4lSPD9
OCqUs9mzlYDxNtq66nWHufO3rnppP4kV1yxC4N8MR0ewZNWvA5nyIK2Y4hagqOPz
2AEZEvKgB87n+T/gZ34evMDIbZIowogVgxXNlSxgqbOX3cWw6fNOjGdGgNDAVrQG
nJfGpoBlzVzMdAksG2PihdXftMzmOfOcI0Y07YfEm+4gh2FS6p8uMkVdzdVqhmHC
ndDeiyFh+XMehOIXByUITtMUZOZAuH7BeWNYB84AsVYWCZfhEFNvWgOWE9YJaoAu
5Ume5npqQQ9nAIx1sXD2e1Clw76wSkKT1KDDiGfswgFdzy3VJg/jrqSTXfhkUDSg
PHc4CGzAIx0xFtIBQ8iZNekw4ImN8xZ4Jmy+OBb/9hvb6MEuTk5uX9hZ2vohK562
UPYtielAFpoQjkB5zmKn9z7hM0G+QRxZQT82o/l1rqQKSUF0viDAhld3TmkaKndf
NIvtEWGalVL4daf0cfz7HN2TF3mRmhoeQwNQ4ZTO2qVluEjGDHnutsFy18/p6zcR
wcrpD0EfxNNpl3Ds5VX+KQ8iIiw0DKM2JnWOkup71NOSFGpgI66WgrMGFh2KJf6s
Dqs1caPlTCEHoabM8pa2E9ndL/eN2RmFbKwfFWsgJka4+4t8/MKthFb7USHhnqti
0VFYcSf4fEiLow1kkkRlIBItuMKDUk8A/msxwgZ89uNGJqAPn4awlbCsUh3RLsOU
bLaMXH2N5P3hMpHvrSZ+oxS4oSbPYzt5pZ8oL/OL/mRrzbuhOobOoe6iThobsXqy
34+G5QGWKI4RzZTt8uSff338piDXtLNlE6Wa9KIDA7Xux6s1nGA0RennL5aB9EUe
v31pMF7IlcPiUOMldotTfObgCtUNx/NsL+R/+axNxqlTsfscp8X8OQZXmBG7QBgA
Duo8wApatJBgnmZrHGiJlw87a4vBJzEAb1qdfQafUYlKJTVwctMPB1FgW1Y8jNG0
PDoTdi5Yjjs2aMQzS6oYXj/mOor67eULw9ruuvjKY+vtKywBkL8QWPlu4xJLuDuL
RyJpeSgS2lNK02cjpDeIFbceVFR09ONzqRMZVD8LMIQ1YvuHsf06OeS53/7s08g5
PDXFLwptrCCAbIWvloDvIX+rTXwREGbBIcOF/pvog30tdF+Hj4/EH39s8mAXbptI
F0BOLrjdUuEVbydeRioUVH9SD7zDISltPS+vBzEyuuRDXNUblOPEGMmjiHf/jTJd
ej6rev23NOixgaSXckGICZPCsc0caMuaPx5REaouawPxKzzvUv4/27WKAAiLyHsh
QFa2zTQ6am6dTrFdysXAK3dpgAE9O52BKE6XMc2uQEh0Gp33qDRQ4KD/5dAVjR1I
MmY803EgNdL7LZ6rQbMqVQJ5r66ufTIOsxHsnePPKKdqC1N2fA2m63h2Utbvb0Bg
P/xGi+fH96aWbUeu9zrHLD1rrBpuBkI2QKJaIpDwnElxIUpGyuWdqx6nrWQg24bU
urV0euEaJWzMwG18fDAL3fv3qzWctdlj7d+TfQPErgMh6IlNMUvUFuidMdNW3fOD
1Kug2RJCWNfhafWxBPZ2BIy0Zl3dJvrCIq8aKA+J45gKcsqFW42J2SnQs3+I3/ua
TCmyGkr0JO+HMT/vs84IW6Wn4tRQNHPbHBJgO6dPyuTOD9eWg+52LFim6eyKO16O
aG7yid4m9acTnmyKzhnPj3qF1i1zfBiPGICYsTsWVkOhar/0+Bb0HJv7OZSyKy8g
Gk19WOO4pmr1WHZ3nrItlWHxi5EaC+1fOEET3jVpbyzuQEO0JSZQNeB63iajG/sB
5vvag6efGKR6yKX1/AL5sea2cg/FrRlJZLyj5XJPqSO6tC+dvTwQv0ppQu4tSPvm
YacWUT88ZJEuMNbgayvbfrD7MflZ7i4uNu1XGHjrNgB/zLw1/XRWVh1OBzUSYE+i
ZhhPBRxLx+JmnjFOW37Iyxm6qyXj0uhMu01nJLNLD52zwsqMoBOJG0ScB8WhbxAO
oy6VG9EChw3MRwzykWHjPJ71o5rmUZHtp7o7CCfSrVbVZrLX3BUB5nigHdC2WXNz
dKL1RxQk+Lx3zapeEBUlby4V6p2TLqHUvwG24PesAC2arZTqaPxABuqleG2RwY9S
cwfeZXJ12/FSFz/8wCdJu3W3/i4SySV5RijPxgXc8hOpc7u792knJCEmdI9Ht0W1
xBoLPCuDx1JDFDRF8WI9PY0dpvewU/BOpp4fD3MYUGeDGq/KuTzPyWrWdNyeA4cp
RYqGLVpiKPRTSaY/Rvs4EbRUAd58yPB+WPSjM0gAyuP6WTqZap3nG8yQKou8miy9
PoLHsrJpWHnGwDh/U2pMEC+iYZTLKnMTVpRmcASpXAUbGnS/d7CJozsq0rcsA3GL
k39BOvJ7aZYDrc4Ni/cUHpO21gY8kVny9By8q34ToX4ugNkZlBX6XDKs/UhsUSQU
ebM+JKXj8cVBmloNUq9Hhh/LvoqVHdPvrUeYukxWC+v07yhB4XNcpi+B9kRflihr
P3JoqNzmDE7+zYI2Guxvz75hfSQXE9nLanW02bpWwe4eVNl0A/Ot6ZTHAmLuexG8
3dzC0nDwj3+iVJ/N7+mAJW7UMA/vNiVdnfG7MB5tQvGyf0WmRJCOutNc0hKnibZC
o5TVajt/sHgDJMMmbcHisgIX0gyZyhZ5H1Op8KvAPzRCej2W3nOAJlA1X0J63JDe
k+GBZTPGhOiiVnzavhEC8DantqYVynNpsYcA0jC6Nl0bWp8G0yv5X8fHf+Gvg6Jb
zgjp06coEZaQBGWzJgRFXaswe8SsLUcBuuVeSDgNOlSNvhfbAbWYtUCwHIHzaaug
zLtDBpidmn+ul5+3p0EPQDimQC0S0Y/bFOBK2kR4MWcuPUF7LG/rGDrJZfonMPm8
o5rIE0g4lDWGZ/QpCwHml4QdAiHJ3Kc5wNLbcHSrM2lwm/BqBYgvCISmowAR3GeU
NtyMl6hc7r9xwyZsL+QEFtG6aX0VSG0QsSZ36y5AOESL2hUE8g9qofhLJN9uVCJK
yD9/I8M7J0xsp6+qncI2hXuDTeZmyS8cfHGIuEbwHZ4TWfkKkeF7ukvd7HigMEkS
bu/Amwz9xcQoKYDi84Qu80r7DSf6XyXLw894TeXet78WCwaHK9ULTPZvr5TKmZty
VdeS5x8XjigrhZlkekHKeR0lKGikJ+PwTQNXY97+ELy5vrxyDEf1MiJjX+ZXIpJ4
qYftMXoh+RHzIlzQDR+21QJ/onlpjB8N1rvvv7kzWOU09ClGQVKuBtTY9I84vQc0
S03QA3Osqb4KNTreXzJN2TCvvmDUVEY0HWbkKqkL6rRHvpybWS/Dt7VduuOdFpqE
q5jFSiCddnNYCt7YbYjDW9niiH+WPd1tt1yJmaNeqkvC5lPuUe6ljfNTAEqEx72K
VpDHwM8FEFAJR6z0bySUYeKpLoMf8qvmuiYCZSpewWUUKgPVLoJyGwxdI17YLexw
+fNH9Uu5iJuE5llKUtlc1RI6SB2igdmd6KSZaoqTav8np+4aBE9gePkNN7obAECJ
v22U5CnGRn/Zgeer5ET3ll2Z4aDtbCqXyPb9b62khQWgfe8iZwDhNDOBvDjMld+L
/DcgGfsltZjF+wUkQrIYku6XMdyQkHC9PnLCk5vDEYoP6/Ijrx+SSgQ1vUp/whV/
iAe4hABzlDkc49kAP6leWOglLUl3xTaQJM8hJsBc9DYwI10rrspKS8Tc8CXGTrN+
T/qUUnizu9UPf6tG8/pJUqLc94/libCTEu8qxn1XsMx62Q15QJe/qppw71FceEFd
c7sJCvL3d57pskk+moqQGfVwk1h7BMvivlr4pahTCRJy8XbtCoDXl3yZ2yPZAynr
vTD6hmM3Qp4uazKL5Dx60PQV3NmizPA+sJUvrSLPt41Ru+YoLZwvsIISwYiHb7w9
9ROr1m5gPtiF7WMOQEiYLjX7w7JmjE2pxHPujUQe1qb6sPY2j8xrod+fFQJtiWbz
wzSxZBtjwxwfpPw2gMML9KWhBXTrR8ZRjvryK0cYPe0BMQijwrjdHxG+48ag2Nmw
A1WVzNEnrLe/Vu4ypk9KJxVCz/QBlXCCp6euFlS1+ktJ8Y03beME9rOk4QLcFdru
bwgoTijK3+B9UuPr0gMOx/DG/0yazWziUmUcwRd8ebqPitW2luDDZ7soAvWgWSYP
qHYbiVDiuceu703+oxfMkREiMsvmAtEg4bA35C8imBMXZXEO73vJZhcAbRE8wx30
X7CsElQoyURnqlYW2NAC2JtWdYZFxka5nqva+1wU/CqE9BdShgAWurr72QGAtJZ/
b+vAARf8OMEuX0KR7OJNwa/EndntjxE3tZb5PHJ1U4J8Y9PGsgA7I03q4GQLXvy0
91RMdJBKx98rBd0FPRzN0hTLhvKP829ZL/h9TgoUsDcUjlWH3irZtpEvPKp5JukL
c0BLdhrSflEpFiX5e0bF+H0Q9CuGfprqFq5V6DpKDb+4NYq1GtTKO9yMTqIM3v+c
1pWyxFcGLKHXUaor6ExYl3SNaWCOOKkAD9gYidYFII8yunqvQBKRcAM/R8FN+nix
cEwMgdrHUBptDPbLqI7XpG+v07T+8xOlS0wF9K4OOf/gi3yuQHA8ABMMfBMt4R67
D6vmKJsdEiEafm5Sxv3tHKTqLrodgmSpuYsZ6x1TWcn603wi23iJKO/qh/567UNj
mDZMTqgA3otyxWoKo5N+LHk9pG/UkyporReszTqOeeBeV6e5rhYuBPbMvcMtI87F
XynVETZtFrv/fFlWd6WqNtmL+qedByLXfguCyB4tr0T3Eq8AoVigQSbiYjz8i79h
/ugWHMG86ZeJFTZvZlVvsET6mbaNcf4MyNelvu9ixNtyIZKoeegO5IxTkJQN+1Nt
697im6Rc2j2VKSJ288jkYqOxNlzCmDIDWvYNyJWm56zxqUT3IDjwAZFAUSwan8Wc
q8BIqXltonGf4oQFCSg+MvR8FX1Zr9nnjtDXSkcIoE8pJZQCidX2K4RiqJwkpznx
fFhVq6Lpk+5DN4F/nxGrn/7eSPiBdjdxKKG1nYnXO7W3RiFhMJmg9Ye/zNMJbPSA
iWIhiaD5hs8sLqbvvwdP/JwXh5SQ78oN5xvB0rHxPcw1+MiUU0Bd+YWVl9g8kPPT
HOURU9yYM9XzGOXmtjPZ+U5nV/VDYhaPLpmOolGYmlMwBNnIekw4L+IIj4i7+HJw
lBxlkXGez02qBy7eiv5sz4HASpz7p83zBOyXpuSzrBfExhPpFmXlgGFuCO6qUkHu
HkgTr1dJhO/evC3gUc5FdxYeZzjeQtHrvAQCDNdHA2KDSaK2ygbuSyAd16ZIB+R3
kgY0EG0SiRiJMCqJtEXe30pU4KZpoM7cJ+jCTQsgNFWT5VAIiFvcx5kifJkh89n1
2uIOAThwDZ6NIcAciAshoBd8luemwfF9WdQQ9FQyzlzilzXWFV8WvnyqWXjZLjNo
pyzQiiMCHpWzbhOEflNhsVcYgBqa9oHqBanbfYNFtOs21kvYVlsSHBYR/1lbmS76
cd59PGd62pnjU7+3rVJx608+O8JRfNCMplh8PV13tgYR9uzOC/U/h00Mt41Njrul
tPMb16SAwYYr4QiOeiQdDk20P6txYJs7Z9D8S0YSBq5pEudJEyFtTzxjBHvQcJV7
2c9Vgugbyn50yh9TlS+KPoVarD607h783FdVE53jg8Z7mwYbHNu8vOTpL0AF+yXA
9D1D+DBTFItc1/tLfI/QMZ0a7r+mVqApN26TrZdm+Vq7O/17V896saA2+oO1lCPP
mq2Rm27/DGD9IGajxalRniBF2mv7YOSV6zMwQl9PC8y0dAXHrneZe0D/3MBRl5+k
bvUD4CXc+J5Tav6a7JgzMiSHU37vZIXk+I/74ZFUY50cmI/kfX771wQkZFoErZI7
IGZJhPXRHXdaxu9F9YW3Bon6pjNJZxZ3TocfzTWCaBZTnhyAezKJY1BPRjwgJkDF
IzS3QwFvA176X5voxH8HQIWzMRr0rI7FRbwEI4y8cmmaZ0NCmlltFLcEwglEh9JN
WFINB8J+Q5eH+ZGd4pdQKwY+sX3bfMOp+GF9XlZe9pgsKajMUA2QvWku4SkUYUlQ
acWosRwPnhB1rXmeSBlg7lq5SznqK0W8+zhGN9onGDUHg4LTrX+8QZTWNJ0wxSaC
icycdhwNsHbZLArgdEjHAGqJe1oWJ3sLcRVGozLX7fDpSKhz/ncYoNSkox56G6f2
1D7gQStsSXP/pcIoCOxewFTZri5PQucPAhkU/AK//Lq7fxUXNJL/Cosg6xzeusp2
RuvpAZAkHDdBABqnCC4HrRfNBl0SLOCrwFD8I4c8tLvFrJxYicvi+OBziUqhY5qD
RMDAzmoBzGfneE8/PDkL7EL+NhUOdxo3zf1xfDNM+xTEtXnzfTwgGPTX5HIEiSko
VDsGJCF22BHeoVHBbsa/lNxftVH0JenJGH9eY0Ye7M/TtXi1keOcs49Ibo3GZqPd
5dnTx29sKeHV+9eFLZMlKNQqpQLuDlaYp2XCJ4Mt1XmQFoHeHhS+ZCWNO5Cdmzp7
OiYMu4vqPfAtXkx+YdhzUyct1pAapn/h4hGOJzybnZWk2byyMlw14JQWb9FPPZe0
FuIwE6ycnBDM/QWin/spb0lNmpL6FlB+A6wfXTxwrXhSIxkUpNXMpIFTRNrwQ9/w
I41xOOGp5opO7PLisV1SVyc0PaFM5KVrcNRyx8rOfEUsN+sYfHxHoPB1EEZE8XMP
zxIFtXFgBDy6NNW49aWlT4nEmhTYdiKKNSALDNh8cU4ZT9InPhSdSCus6QgNTNQL
qhAw413cQBzyG6OSGHDcKUSY9/E/r2xSkO85r1lXoeP0ranOHi6C4x2n4+yVujmP
NwKzQhv1bJs1wM2rS9HjGE4Fcscf3A/ttl4Z8RntuYau0ZpkqnnXMwgNbcsICxt1
IqrnGgbYmaQ/vm/6SHyNDTLlx5WhWr4fvw4u6RX8DKxtBCKsQdiwznGTkLdX1ZW8
wUEeqAcg3Z2VsUGyaCklCwq0cMohC9KBtbzIZwbnOYw00qqsM3r0wpNlfU06hsqc
o1IgiLsvtzv+QlMa/GLKbURWf8wr9yhHee/qgX+qhxIUMnH4kszLgGNTpH43Uhps
UyJm82gaVTSHMtIp+25tyjVRMffieyGRFxnGpSRnU0ySyCDsXJ+8cIHBYKtiLmXo
bDwXzlTr0ny9lg1K+b+CzInL6TvVuLHYl+Q4m+lTUmY+87RM2cQPyrpTfoxrELqP
/Lf9K88Cc1F3OzswCZl9OhuA29jE8E/ViKfHSKtl4G3p3X+xp+jBkBO7G0LVwG3P
x0QQYZm8MjSId2kbnNQjtpT6OXftiNyBs6RybX6y2jbNDypOHjW4RugN4emdu1uK
nfZ0on2Nx+zjUZEQN6sx5I4K+aqPc0tuH9y26GqiVpoTbCDGxpiRlBRYWkfva/Lo
zwPWuUd3CpzSVhmWgFrl1bpqGUstLvQfnUNE1ryvhI40vEbrHz9gWrszkVM6ui2O
ncRx+KBYo6v2IEYe5BfkaarOmFG0YKsmEIx8Usvji4tSmDaBTeyBNbXGFTuZI0x4
71HXCUld9Slglk9R9njMlqOpmbmBcMrMVVR153zrstURhD9rwFSFLapoEUhwiOj3
wUnvegerym9TRdjnDx+sR+3rSDjLcmefk0KiGnst359OebmaW4f9qA4scsoGPZ4V
YLj3g3j8qG1J7UpQWc1/uxn8IqBoixlEziJc6hrc3sZWLjck0eNZvUYTmJqHPxjg
fV4QDj4P+o4yKOW8VgKnAX0xy72pPVhTMwQEcxJ+HrJ5h/5PxKUZVbk1IRretzQD
UvEuZ15hfhpQTTFlwA5Hxmp+/ixtTcqmZdks4pUCxxPFGdzFWNN0TI0+2NRXjwiF
LleqrzXNmX3zibRlq4zVpqtfcBeZOjBYi2YGd9/3TXjXEahwVu8PhcxQSB6oGnAt
Vy7R14MiH3fcdn3pgTICexjIad4FhBFoquKxqVfsHk1BZJOs5FCtn7YRM/A5QRTP
71VLBSnIruQv2JCAD/F6wZOaM2ZjKQChfggaHPf9Pm2NpJslNCmTYRvjC9sQRyeD
RAajpOJzd3nPt+topeLG5UCp96WPK8qiNzsjcVVShkSN3Qp+UXw18Fcx/mYFk+c2
OnINg+KBw9PY7dF+mXOu/Z/NarkG4SwK2lFSjt4k/wjOe4XWf0DXsG5aojOip0AN
T55vThq5NbDHID1kyfkCW+t+yyVLAx9HrBScTX5KMBycVdfBqZvMAw8rzIRwI4yY
fguxidRtVb+6dRXEf0VkUcVVsusbNDysCIFSMpMeSqPvpxHh3cXXoW9+xWE8zIkZ
EK1vqbCpWO+e9mskWjFjjqv4vyQGll7YdJyBhro9RM7Wz9pXH+v4MckCBzsWTxwD
YaHkKK2v1rRmVutKqE7I0wz0OM27u8LXD0J/duSDxQW7785j8rvcRmdJm4lHjoT0
vOhrsf+vGqQE6uPgmIK8XsbI6Hz5C9voL+qj3h8R6yaPB9/Vv9M6phbwSSrctqYP
jmqcOpcpeaTU8HxRotUOBtant6IGGgg/w4LCdOtzy5zdl54LX64nfhrPKIDdayO6
i84H12vmw7kDHGSaSHMXbH6MZNyEe7mhOZ4gdIummOHdg4hnfm1VvHJvbnf4pSJe
Icp9VwqGXBwXKg0691XS18oOUI6fTs20Q311loH8cnUaFQY2Uyb/Rsj+0qD9NP5s
QPhGi721WvnPnDKRH6x8Oiwoqqt7nJrYHnTf2OTY+Sttlo8NEYhF67CG1FTJAW5c
8tCa8cJ0d6F31bWHiB6CJUPun2InRSs6rkSXsH88PabA2RspUzfBf6DY3PD2f9bE
dJ8a1EQ9jC9QVWZEOuFsqVqre4IFBXdFip36O7j9Tei6qMuJlPFvfaXbW6426Iqv
rIoo9ziEwPjr/HLp12fNc77/PsKsAsUH+GAYKkX66U6ndMDP0Fo1vkkP9jdCdXIL
vUBN5a+nrJNN3FhNvsI4M1xIEYWd26F8FUfuX0Vf2xbzTtbNR+jHumiItxjxQYVg
SRdjpPNHuLNKCI5V6WdiUJwjnqTAW/2ktiNhjahGu+DR2vrsBGC2sEqBORfsdWfl
3n+FJjYrZq/5nhiYnX/yqlBa8vx/eE2kKTp3M46he7xSVHDmqB7Rq1nF0KbpgIEe
nScngis4MhQkM1LlONT9zqOLPNyOG8PyvlkF4mLZ4X/feT6g3tOY9OuxMMRmGUwg
ATTOJM294aSgMD4MZxIo20daUeqLkgfA9tSVVJQDP2fCeOcX/tiwPWHgdy2Gh2R2
d01pYH+bfCFwveftrzuwW0GRJ6UGoAclzUPtF9IBlo5f5C2swo+P0t9rng8FhE7B
cbKKc6yAxVzjNTcVZel7SYrzrrAenAx0ezYLT9iCrK5UAKLk5R+aqWQ5SjbKjpdB
rop+2VKq+oh9y66V1yuQpxyBDYG7KEJHWFYwkf+KtGiFnrOpquWlnzeMQ1GTMZb8
oWbIBioNpx0xyP8mitkqaH9xpBDRilYV8x1SunOoXq/1bCJKA/5RfyCfi9AipWBP
oLogW2fcw6VRKsdnGUcG2oxN2D9jsaGOYWIG5zIKu20i3oJ4X9pfzUZWXQv2+4fc
LzcbBqDqfZiMJZhWE3yU2MjXUWWfp/OLTYZSawLKe7pXNZR18+9RQCCMWnn2n1cW
szWMTqBS+o/1IWZrcVhWZbC4f4qU9QxvKXebYmPBMXjJb3WMz1jqJ5jaroAFA6s0
0cDLgX/6mVFGrZ9tfw+gNHazfgv4/eAH5BUWnpth7IPcUfwBpg0KPL8OfRT5HQnc
fopLQPl8ClfyDMgerule32E2H+4vqrDese3YqZm6hr7HZuINRT2nR/seT5STWdsi
Y0BbcUSEJQjTj7ZqEX4NNmHzH81jv2VIZuG6boUWvrRY7Vapq7LUCXrHr6kDGCpS
r0BAGX0DCAr020hOPcnivVOn3h+B6mKHLInZcHwqi/Xg7Q1Js6ZHq2wu+2c9YXZo
kVzawFehCWOfm8cDkgEeiaAg3d9TVY9CzC7JnbFwN4jZs84Bg3Y1uhkmM5ekYIbf
stISC7XWes5tRU3RZRRH9V+ymjzCnl4QXjX5NxTvb6SojG/RugxJonD9HHqWNeCS
81gG/eUuig7VkUrgSD4Y9I6YiWUvExlNnaMjcqgZ9ixjw02q1EJ6AW85FWFOvEkC
BN3l82Fy0bDrTA79pgrbhgB/sxb/m30qRafPf5Umj2lAZm65vSID/LGMQufz9p3w
qIufVcnzX7Ccg2RbjdMxO5fBnosXyYu1kfHi/mJfLmC3Dpf2wWzznCUh9S2Sklj7
jf7nLmI+bb3XjqtKqVs60bJXP0l5l5mNNJ5oaeufcGlK0ERgcnXVrO5hGH1ob1TU
64lPq7kWKqWIg6mk/pH1sLTw9dYSfZAnIZiOYajoGiGXobGJiZFzU2Go4zANQFjA
yiqlk7ZESaypVO5gywHxccaJZiMAzg7zz77LU7hptgMlSNX/M0ZndrHyQkSMi/fH
riVujyNwjF/EumUkGMWa/LriQWWXVjg45R10cXBUkmm32Q366ytRFtE099ufAr8s
2ZAZdbDyBpMu+Hm2zp9aI6zcN0dMSakvlKC9iK6J8pjbdAxhICe4gM5H0Syeyfjb
wElsGPrgpVM69TYrMdERmEMK3AeWohYkeokf2Ceor/kh0jV4hzINyau+f95z1Rq4
E32xztgY3TAKAKwF0wQiYRSwsq9eDaI0dykY+Sz42wL/EInMPXcuHvBoN9T+j+p8
59iDix69dIOOux708+Cpz0wQUfI46C4avXoTSSdCLsI3D6BQ/7C9U3Tquy01vj56
5jvcoiaQFXhbFbzDieBvMf+1bpFwRSlEIIFbNPoj0PAuT8gk3xhCtwFk3oFAuywh
HSmAoGG992IZq8c3xTuhqx0xosmS7nNp9ldnqAQHv+QlWY/1sQ3dPHmYoSn26xJX
OpRbfAEYQDW8c/RFaqn+WhttAwJjuObmM/hqA5iFgCNGFJTY8TQ43dALYN960LBD
jBqLxu+OKaXSh1FHoAqbDcAlamFIiqBZOCayWt5PByJe3I5Dz+ijoDUKJ6B1U0na
lT6PYRYkll7A6uhD8zf9ElScA/tyf0aJiK/Xo2q10NxhTwCpZFITIAlaoYNReikn
C5Ur0GcZSPQXTb5Fudk3UtJ1/FjXBqL7Mc5F8mV+WaE9EcVgQgYYqSWO7DOZKmlM
UcyghrIajhmM7vry0ceq5tYaObVrNTCwUndvS81l1XAbRzuIX+S/Yk4uuzfzG+MU
1ycTeO+sHogzJCu0B/T1uNkxl0bGIEDi6E6IhNs//DG9HEQjPY4EqpUa8IfQaePM
fEi6krWkclpAKDzuvaXbun8ITiFJAOXYHuCLveiW7IGuzChaScjsWfMz6rtBqyTK
Y5c6cmsxpmGiI/1cbg0R+Y0RU+MM1A7CO9JbLOqJJyHdrSBzkkXRMlkkqhbJtijl
119Kj+eYxN3EkZjvSy3jspcsIgdwncQzfsB3NXliJa+pzQe5/nQpVc4gM6KiOcgD
mp9QCDpmd0wc8UDpxu7G5XL7kCjUVg/rjYpjyon2x0wnkcCDtCfzUjAQdX5AXekr
AbNQnU1BbVIxCB1Qur0rl2WzwSVzvYStFLpMkE+KqEp8kDdgU2LFT2YUELcyuBQe
kh57NVfA26eyKovMZx8eUkxHjuC7pO4AWyMeFjaCH66RYWv7d9X/Y36HX3W6oUjZ
vyNaXpoznj4RqX07FxFbhNF9srNmyErFq3JMlQ24n7sNnnhjysqHIr9UxLhz1mZg
PfreEHKFsyUmbRXs/1yv5qlPmcdgxk2iPSfNWNFnILW0wTDIRGwZzJ6cvEmyyVVh
Xv1U6O7mHRl1zSpuIupfWVlqOV7vNdrGqa9R71DgQzAvmwWV6pNy6ig/CH53z8m7
AXYVpDDq4FSExxu4LY4JiNt5c7PVCsTw3Dqx2VVhpxJEWAjDJPaOhIWIdzDKnV6y
IL/qWp7WfG12MwxQAGzgn+Gyr1Bb3IHkhhP8k0hegK9ED0I0hXc5n29rmRg0l8RT
FK4PO4wdd1VFxCKAkirtXP1X2rCjrEUldXPC+Xkm8pXpYIqswplJkTazOzJ79kzy
PnCrC1xpTYtPD41pcngChIvup1FppGABa/KdzgaXd8rwwfeEGPACeI4APCODgeCt
JZvjRS65SkiXnd+OkfQ6LjiOdCID4CZ2vaV7Ai0pbGbohSWPqxWpQVZ/wYwL2lYX
2PSuTj6faTw8nt/wxCbieN1IsuiEgicNuPQjTgL4ol0whs7X5iJrSL1PZWG6Zyfv
lPZ8dJiJkmXEvxENNL6P9QlILEo5nVP6Y8r1XgyT47qVzMLubwSrZTP4fD9PDuqY
aCjQ2IimBtumhN7poK+g4Jfp/+lUCLts5XUMAeu/h25YsOe5otC1wh3tQkxT4ubW
vMtb+v3Fr7qtT/+ahDXOmTmBR5S6uijgjOQeGUZGTerxdzRQePj+3DE4GvrtT///
+J9ZXG98vbcOWbEUaYL5toLxt0y1p+umEM2Y8xTMNWamAZpHrmOBBrRcwrXw5l4b
0qAS2H1i3wzEg0caGo8cs2QyQlcQZtzahsvLlxA/ML0Blvu/EF8pD88iEeMPcekB
CcfEfv0tHsiEy0rXWsPjexx/4GdXHvOXF1ZByHcsQWFwohauqW3AOxvkfPi1MDwl
xRtPwZjvmQTv6sdeBziIW4+f7YuyD5Qy7jzC9312oTUiXhhI5rugRgWKifIUS4uA
T2+UlnmHTIFnBSpanpJhrT7j/ySRFXq2Kk/IKHHFtBZaC0CvO0WV8ptfMPWF7scV
J6RlQc1CrZrIbVP+EumqM/CJqISlvpn6Uh8y5avILgmcrSu/x3fHb81xPy8cNPOG
LbSeUsPShwuJ92vWdhEI2CJe9csv5tHuGAA64R6+wsDzZ+zeRs1TpG1WMj4OrLuC
Uar5rdzzw7LBASyBnY+WV6mutChQVmIq6GRXos9pXpVIu/gWEqvlq1fUHuUSPBp2
j+DiYtgfzsqltq+yRE/c+3C/zpTMt4pTyLLjtC29/ForKXRmgQixGvqcSfmG5Pg8
0jxGXDOfGqI+pJUTY0tVCaN7m+Urn8j4Y0zSSrlOplg/WqE36R+KZClhK7RfKKLH
7ifXjNLoIV9gwB28Myoq/pVrPmFJnX7hQoj918lN0KDex/EZx3PETo9i1ZPiEBQ6
g2vPWO7UisD+myCaM1cFRg8qNjnGL8ey3+08lRSk1P+Ad0VvehWjGjC7RwZczK8K
3ZROodL0UGmKua0cLvtMO9m/ztNuqvNyZ62BjDJRHvzDA3Eayz9M1TF3fxYY30z2
H14sWr9ZQe2YPPcDfwXZ83/FZ7lI9qlGVoKk4Eed7pgVl/gss8jt476HXhifK2BF
CvsovJxpznWr0cPJYmepRisqgoa+YheB71ealDd9H0wZIS3VP0oqZfoC3rhLQxD/
yAY03esFVT7VHjOxQvjvJSGqH46fd88kkkXWZpFuBTFARJeUfo39t39S3F89lKJL
JZO9hvFWVjVLZAyoqoJ/zKtra3T4s2OUbsoO0lDhHESv6EzMD4qDz+wmM8zsW6nG
LDYdHWi9XB6MTOQxLXO8fFxkBfhVjcP13kWMA2J9tOAA6Xr4XSfgUz5NZR3WRRYU
45j9IsxXJ3P6K6R7rrpELeA/UBPHK2mFKo55pfTjZthWbaqwO743FaAeMXy4KG8u
tb0RDt0cq+Rf8CgNaWTdTRZZFvitAOIFn8t2lgTH5JGHTYVrnEfMyRIUNGaji5x8
PTfQrjFIBkQUi/47rnqlL7KiNcAvAj/krQZpF01eKxwjv4+s7+Ww+G1PoLpOfzb3
dLVtGsIQJex3P9xloF6DFv0iS8k7LMHsItW8HdVWe/f0ztE5izKckNRa36V5lhug
d4uhc5xwqQnxeP9EPmEhWgkCmhYZCQ/k6BCOtNoonnLKIyV3+Ue1iLlcVeJiZSeE
PlJTM4+FODYOe9HSep5pKD7bhY+lKCkviAYQz/uJ3eUFlff5geTJ+CASzGiswpMs
Xx73pYVxaqmOCul3v+MdOzvalzKvcrIjzFPGDLfe4BsWJbWd3fJP+7XCZl54GN1J
0R/zyScmcwlrVhjZajUMs+xSumgyugXyu00hSzIlbvzB/DA6q5IQMKfa6nORrKIc
1moTE1CEiO5n2pwGwPRO9HNO3BTKZOoAbdV1C9NivaEBZcCadjTMIm5szex3guT4
/nQTcgIiAuI10KzTvOXs1dd95Nq2VJFfjs1SkBPbUf2PzkrzhCpLIGXPo/kuCLzJ
qiXcK+khnjRIzYKI2Fvvzkl6kAbLodp0VRW3AdzH4rWhdue0eRpeqFoq80MdUEW6
e0DaTHYmsogZDlUYPK9csp6T9nxrMOZizMxd4QNcTHjIINOB94pwliZwoCp3iVz7
FWXqaLyM0bBK84ZA7BbChgM6w2UNYZGMAUIatZDaLuhM2jCeOFxGAe8X64iEjnPH
2+TPG0loBtCzEZWYBz/3nf4EZkLCeEO9ZO0ImQOusUvfnSfNF9+ETzIKti0v5EzT
NevvdMGYcFab9WEgOVRVd9Jz4HeOlZK6qZSksut+L4mbyyF4lHN1CUxHXWWOhwlQ
um/y8NaIj1dZVawCAk5wMPh1hTOWdcXr6hLzrBRC5Pteqz0n05gXrmcR3Wyfzceq
ZNWh0BLaZ7tkZQ+CWhrcKybUymAgwpAIZvCgmh0SerYHO+Ks2AmqhHMN1JeMSMaG
DqLi01bPf620TlbH3Ev8qhx+JJt6k3lQxqWUrZXXLy9LaFBlNufIOmAeCA3gts5p
pEk64NNc+UmFhOtX/qRBPupM4AyAg0RugG5YK5kJFADGZS+T4VF7eaKDlHhZMtW8
wIKZoYM46xDs6i2p9z5y+QGk92q/wZp7K8J9Y8XGxbtzd8z78G1/Lo7ZcvRjBOkF
wH4V8035z9jMiOH6cO695H303s7lcqi9uEX90wzYZ5n9RD1GGJLMwwUtVNL4EePQ
cUURaD+7ktggQPnM839XizodbvWLsjyZ2u89bP88TOO8AN7Vt07HB/fffAbtX0H9
aZdPW/zI09STVqKWUU4ZW/g9Fy7P3hXUDmeJD0YJVS8FTDzgo3xZcZVntc+1nhFY
lItNSblSRXemxekB+Pera79w8faH2JpmOSKtMfPQyDS2NjGSmNYdvhYrBgDS4pK2
1wYn3uCDV9V7qsOxcrwu4nUd1rIo67ixlrpVR78wKpdaVC+throQQAmzko+zQ3+Z
DLNIRNtN6HWDWe6l4hmK5ctr0TM15VSHI+NqJ+pILFzogwaaD1VhDthlh1XvzTJd
Bzq23IZXdjN3g+rMKDG/r/8Orlv1UYZU2lMUJaaTKqxsBocZvQPxZQ0VgSRQKbdr
XH+2QKl5H+4KgLXFHvn4tWas8dbRa0MdskKMbz31GcK6Is1ba2N2pW6MnrhXA/wg
d0E33bXdRDLOLvEVS5MHQj+Cb9/An9kKbWHfa1J4DIRIXi2jHLG1MORG2+9uE5sQ
Nx4MQ4AGFEklZFeuTGO+ZkKQn+faRXKEFKfi+XRGHPm3EPgIvMdC9l/dgX7S00eA
LGTIz/it5RRupz2r68wcD5TWzkXdhnceBSRgLrdOnAPDEMyFCxi6lb1bwgfR8nYE
1fG8AGZeXQrDMLzdwJVa+nFwPPZFAHgY0Jl6NUQKX46IfZ6+wY0Q/iqDwBwhqDWI
ddZjhZuedGGpI5UMZIMxsSt0RwY/PoYHqpb1ZawNcdJuIiDq0MSNoe9PDYW/cndE
rL3s0Fkl2OypwMKpiWLcrTzzBKbCZIe/87b74vhHOh0zSzxNMOZoPtuZ8XLk6gn5
oy/mVXvw/8B8xsLDI7tge3PmGYGGRb6q3ZnQDcWawcLS6v5pfTVqLq0aiXFS3Fcr
oFmuGBcPVnkVE9v6AINVhPTjbgeBRXZ+mcTBlsw9u3cuhkhKPh+0fYlwaEKS8bas
LacuEVubV4kzBqy0nlmU1/NY9oO807P6h8sHdqaiQLUFKGCNox/CALzNLOMR4efa
rhnxV2UPywdR/c73ESgEtqFXTS66Qu1e+nSCF7pnD3+BnXj95/tTiA/mLhz1Sgzt
K93oBY37apW+RHtWh7oqc9ai3wXbdTOZHdMxTwrkFVZX3aP1UGhMf7IwK7S/xros
/Fi6wPrusNKfzTFUW0Y5p/7M5gT5kOPF4nDh5WhYDbBnRbIZ2ZIWuAQqaabnjPuZ
Aki9Eim4nqaJb34D3r7P+fZjmow8bVOmTLM8/0qS/i71UP4rj6Kk4FSW34zlY7vt
siYqQGgoGvqlABgZKgXF3u6qajXpbiZ2yC6gKf11W/WAkLeJjxfGxA/3dlkELXim
pbP9OQvD+h6dGwUeC8ORljIAZIN2CKKBvhIiGvbDlva0VvHbPVANHLgwe9yHXv19
YxFHaPWzV4zubAOju4F8WWgLmN7m0H7xVI0Gj5Z82ug9hwHuTJ9C4S4/O7jlKqqa
/acMlubNprvBnOrE4CqPsshdFFuygEiB4RE3fmJDs/lsbMTK9+eKH6/KW6IPcqPa
R2zR8s/0pC3m7viI5dFn9Qbb6zGFsKY4g+PAJbHw6W55z7xeLQyuo1lE+x6llDg+
lgoAHPygr/qG2cMoN8c0969n3Fj5avfNqSawO6XiqtBcFmYPmzFJVfCJknLCoXnd
C5LDvNDb6ffAxKlBIjzAmHVo1hT9dYPp1E1hFBigcXDjM48lBId1+d/iJLIMJWwN
bDZI1gUv9M136FTJArWbimmUfBlipCAWqzfs8Ku+dc2d93KDc63FESP9ef9CWnqK
XflfQeawQudsaDtrrtqduwFHVHT6utvvCswuBGC0uoNf+huaLDOYeipLRBpViSFX
u9gf9dK1dBmj7idh5+MrWOqiBvU7iCrg98XQcutcOaLCFuJ6sGfvwzhQBmp7cSMI
Xvj4gmJHcsBVjoGabgEyb/+TiRFCZTti0mvBDKJuQaNm0PzL1olugblu3N4DkTqG
039tTDlUm2VTmQ0eH0MekgjFJNon7B3feeGSMgkLjMzsSn1MJaIOM1mBR7yzp3Gh
nfMVJMrX/9kmV95Pk++U5cVluoI4MPUsLFiDu5zKCOa70CtoDHxfhziDaLR4BXgh
wAUzncknjGA3W7a7DzmuXru3TbjMwN94JsQ2tu/FXoHZhgCMFsgrzUrVnOUhayhi
F+9/g1fy5aePFUXaE/Yeb8hQtQ8lTH0iRx/h2tz9CP9dZwcUbwOWsEsz99wgrzvY
TNSCMykl7QGVyMdfYq8WXirDg3RSAFz2Zmhh4jber4oTBEhIOYEy/7QpdiYiEAFL
Ch1/UYMhySwb3GhB2H5Bf/ND0MxFO0y7zYjfa40y/tNJG/okrPa895DvttMcP7Ki
t6xOPDhZ5VpriAq4HhIjDHD20WO1lNO15zZ0V0IfF6OPXjYy0igZy8u+vXFoE1Jn
fVJahh/VzvvMxqNeGpWg+31MBGPX6T044BNVXJylsOlciGVXRPLEdHrdvIxda1JJ
yYhGX1k2vdDGj0jQTVBgSK0RKqNAbDSLSIj1vh57oigVI93zWZfqp8P7p8YhuIdu
WAoarUWkJWZUBsNYX8oE9kgTGlJ1GYXkNptFfsqzTfBhUURsAAA3u71caf2TxXEz
0IU00z4/NM6mCkJw1sPxrZzkawCbFQ+we49MdfQxhn4KZMixyGuBzqL0Fk3FSzW1
Mz1qjISyEdPpsTz1m7WZ9JTaL7BcsOKhK6WsbVAlbjmoBFk4EENalvcYlOJwcgJG
NMqu/GUgCuBf3eNkoDSAvydCsc2oYHROw78gcdxmUbQQuLryZMxByyQGS1DQHWy3
DOhRYh6LvOZrVwMlM0PsBq7suL48RKosiECKUIMOeYKKNFuzXtkxwX6at+M59ttx
NQYkVp92IGxWZx3ZCaONigdz9Kwks2tSEU3mwMargFP1dfd8z+pDI1q0Iy6sGnma
FhKmKJpwA9l1elm14AalfryUGKZVJke1kbba21Ct5Y8g3D8SGkoeRM7Q31YhaN6j
5XMLX2sNif7ONJzkDk/8ggz7/WuoQqZ71SkwMRrfh0yT3uL0RCYq3/UnmBrqUTQi
PdxarDyQot6W6/Pq8aWhntbL1bpnOcCfwomM4kCB+6CFW00oF/e/wcBIFgWeQ+j8
0l2FO5hDx6nvIBUFhJDgksbqNTaQBPc0/VNyIpmE4jbhTiH7mqejYTW4SGn/+BN7
nINykcVuTUq+dK+3eNu2OVbG4Yy8FicwyyJa+8FvnOHVN4JmpTzBlPp27kuR8e4C
Y6nW5OhX7tCtP4XnQ+DE5EfZhvhyOJxJT13Xk20VH4egKPRQVF2yw4C0JXGHQUtq
EqXVK9kLo807DggXTylz9peB9BP3a2PlzsZjkGUsdIPm5QCa3xEQGyHIh2ea6fC2
NX8UOEiI20jMRBSSIfDksE7B8b3N3/KVSPNGAgzy3QceCXGn35zcGWjkL0qGOe/z
Ybx0npZezSw/4tYRPeepy2wJydeLp6NAghxQq3ELWJbJrfIbX3hW98x2V3A2Rd40
fsvpGGlhr5Cw0HaSMmUgG3pmjx5NGqgkOXV62p09/oU8wOc6Pgg3gWxDdm1zJO0a
awHMyHptY7cZBSgvF1D+lnvL6jS1fGX+Xv2hWoRGE/06Ey2Z6xXXqJCSfrZAj19g
E/qQgv5FeJan4OnSMPxjsLyCJOn5iYoivtEkKfCF2wlweJh5CM+8ouGMOUgysS4/
5UD/um0pgFovHx74Q8l+1r/LGpc8eesrvYbHlcQX6AgD+H3C3BHoeXjGaaiDL66o
ZPnwXwrTm2HfpFzManvT0I0XcfQUrqLjrRetoLfBOv3jz3FiS8VdYGGEm8OyFR9S
Q9gkQywX+k0MKHxnTXYGo53iP+29gKpGCMB+lFXcHRDuu/ruyf1WOMr06wLpQCum
lJKYYXXtamj0KZuxn6Jq7pGqniz5gL5PvtlT11zdn0bii749UPb3Ee3gNcW2ASJv
YlC6xVum41085eXt/aKM3uudvbH11sNOe3vZ28v4hC2vRUk0qecS6GnOJ6y7WPu3
a86tmgIl9dwza8/+TnOOvWT2zY7JgAaLMoXpJ65diuTF3B1GcpGvcApwqL/2exCo
kLU+H2FF7mcVvk2C/NRLXiqIv51z6StLz7RO1df8AVWzeRmPHayy2CXbpY1Hm1Qh
/NkyMNHZdytZ+fQbsHq+vFa4bxUVk2Hq6XdH/2iXMt/iC0mbRiWhPe3zwY1BeZ6l
uzH09ZwDeioiWaXLt1WYOAyACz/49RhkT9KauAmnjgN4RDKpORngNE2Nh9muMelY
ypOYm1BmbJdGzegt5V1VUwft+AmmRFAT1vdGH5MkseJQN3ndd3VL/ENp+GoaWFRs
LojrUeEDwLBCeLHUu5MQGiSt+OT3oeMb96nnYCcoWEWQrjVQhi7HrZq2ujCnMPnB
02TNI4TlS7e8gPlVHxH96NRE6P0tAOdgn9YQyloGHP/ErWm9WVkTDP8yMI3RO9j+
hScnOoZzMcsqBGPsXQ3xwf2ICKi5rB/05v80EmBvHo+w1YonL/cKyGuexpXR2b4/
jmeMS3HtsvRE6d920N7DxcAydx/JQjQQydpCpiMc5LfJXi75ZeDebmO8BaTF00L8
esNXFVGGzyZYaayTjlsx/XMBoeCjHY9KmrwvdmYORyf3AxXm68Ry2rWh23FVvDDF
UZkihRiAGhm6rHfIP2k15IUiqwgi7J9JMhGhSHlu2KGURYbD+tWZGI6CJKlqn8t9
RssYSng4aQA4hJezuhuPNl/vQpL+tiS7dq1SlMnnpeKqtn+1JMrKzXwFJgpi5pe6
D96GabAoeif2H9T18ovyz5cn5Obzs+hlQiljguqWLzs0kaXimzI3q+WidxV6bJHB
hd4Zo9ttRgrmafoayMgPEjSv5HX4/X12Sl3P5YPIzowGgoJZd2DqDTAYvJoUuNdV
2I94CLGgvd6bI9Wp7mNtRz2qV/BhbouebfsznhHNGs7q/aQbjwktFakaTiQRAgNK
HP34eLp/86KHSpiBZ0t2ZpKQ2vHACn1qHVAUIcwiQQ2cPMiM/sSL+Dq+e8S72YuZ
4WpLoBouTsR1ys08MhWWgNJgXXmVDQbZcB8tObeDRjMAt3J5lrmbs2zTq2B+Ociu
HX21jVEnL0vP4UaEPio7SqVUQmW09arW1gFUCUWLc2BcCqJkjxqMskoGkCQ8GBbF
P3jfOrsOPkmdEsGdmnYAbGTPO7qrYg5PwmGlEVowggE+krPARuGIa9kROf2rsUci
PfAeA046fAAtRMfSr899JYku4MU79g1dm5/fjJpSEgCo1cwU1glwo7N9+Ji4Ud7m
80/SA3Ff5HNMIiy/2y4fDZK/XyaBbvGRIzORaK87vMl8rfURmfvTUNerWaZrYvHp
5y1lE7IBov1UatgIISB0zRDEFpl1qHq9yG/xb/A/pzp95dB5qIbtFDECCxSBXq2B
uRYm04k7W1vg1Am+dOmbHfGEc6By/xUENRkW1FjjZp0lwml6CsoKj3ysbjLdTEoD
gclID4tvxaIcZcEoxTbfKxODjRKKNl5+02SHAE8zbQzs0Y4Lx8GS08JdTICqhL+b
4Wrl1kcTKnPOsChyAEeqa+U0Iqh1BQp6mzj1VJv4Ltaaf59b+1ik2RB7jwszmZ40
/5pHJjHP7GNSzLlCQcHJr9QTPIEFMlk0paTvACFAd5ZulWouNuvRutLruV1AkBUg
NIOtwBBa0jNcIXmecY+YcV0KQA/Ci2dYYxuzmpa0UZcw1wyOEIvIJWx0GFpPG0of
IiP2HHnJ66bXR13CE9LcTlDJydD3oUxHtK4q/aIFdS/fMh7KTqkg+l4P4KG4buNE
PYirMx+J3vcxWPgE0WeS5L6b4tR8za7dWtqFAsl7Sw7mMTyQ22VTYvoCUbX/5YhB
qz5b5l55XClWucSTX9fKCQWeZJYyyAKv5pQV/0lv4Cm275CRvwoz8wWfvTbhpAWH
WqHF0zWJK0HXFkKupj7cQtkfui0LRAshl3BM7IMd09P4omhEEz3Ixi8WAXzoLCiO
zEwF2HYnAQXutzIFnspJy/twxuL2ifuBJUUdJho/HOhfobqgNzTOY4kP6kWorSb4
2qOXg7tkimRIDDSskDGIAAwG9R/zZXqvs74E5OlKiS02X8Ri8viAsdOiCcScR/cd
phHO0fPQfUJWEiWC+Hpw0d/Shz8mzsQa6VldxFCCWIG6zMMFTkjjvjW4MDPTkRu/
Lr45P6GY6b8cPDccqRmmYqx3BzOsPemL2ci21N6pZFnOyDZpjBQvXWqMGRNHQVZ8
p8f0Md4W8UqUhRgkL9BIwSs6aXHpGN1Rk9m3UNUO1JxQtE0OeZ+6UwLuGAWIyS7c
ufa+WMzYjxy6tkyutBQTDTYHzLsqQYwo+fO6Yy9Amf7AptYpWCeE63nwNsRY1+AF
waKFLiZTG8u+QDlcu+/uvkS76zSEJ2pcXQITptoi0LyKX2o//DDvkVVquF7cxsCm
R9gKQTV2i5yMBZzhAfhFz+c6xdk7OzB3fFp8adi2L/OIMW9mWaq3gfIWdmpQAXiP
eb2jWgJZMycv9KvSvPNyiExaU4Dhxt78FLDqJ/14nsYk0f+7YwBLJLIijDO+0yTV
un0nVR08q0Vv17oUUDQLR8XDBr5CI+Wc6Y+V45ATLEA9rJzFbnA+iD8kEwnXqBH6
+fjXQH5SAalTm59/tPqmZDbu3hwgS8c3763lAihrBKLrBzPXc5f6KLLBlxM6C9a3
cmDcom8EWE+tmTwHaelXaxXDuFCyu4FtgnDol5XNYCwvk8xevzkPWMnGHETcgIwA
qjWtc1d5xOAhbae5glsZznuUYsfYWsyFuaysn1U5bmPImjcne0q9XpLMdXzKJiUS
C1Dh8XcIZZQ2ovkZi9SvXOxXetyngLkiVj4P1R49dlqoE6dc7bWbAY1kxu+y6NYM
btzSb6kUSAPfxcDL8d8WDlKRYaQt98LHAOdaHnPoEEF3CWjpWpGyLBNPTHSe0isS
27H4hITd7mrvRqqC0c1fO4z1PpXsTJtwztD7q1XmWQe3YMM+WlApAl/R/+wrvT+e
79AivLJ8SReUxk40a3/VSUnjBSxvTjZrUqShwIbgCWXxtN2Ngm74QMdGApRFtRWZ
NYMWIAU+b0ZaDpBk1wQ+Hu5vyPfo0q7/6orQcsUvLhCA+i4GbTsJJyLBbfTXA8oH
wlElZVWrg85AGTQcqU8JHcbSJzZ6sq0V9nSIz3iSrqkQ/wVk9tSoV9po25VsDql4
EYyQiLIXanidnydT7htw/QXd2nTRa5EFR5IWa1hGGpoCwE9vYDUoCDO/M+5tO4oH
veo2a8mTFv/zw88rz+XdmW+bpurTbNCDZI6IOuTXeIThx63Yi9GshE0UGho/PsO6
hLoZh56ZqpC28wMHAF3gTWAcxdjq0wx45tGIR5Ztq/cBuGJBw8LGKwE7Q7In9ey5
dXIB4CcDlQCpgXJYd/eyKqHo0RY/HcFQkW+ZhDdvcBY6vji5x1FEIUNTkL1DMCDt
MqvnUqiqYG0jnYlKEHa9OhdXzqsVyNBqZY8VSj8TTdDGSVXnZz7smHXzpOaT0+lL
AxvZdmaMk3jrJ0sMai6YxEaiu7Uy+UsnqYL9qzqZ0LMmk6wdv+jhsBrZAVyoZPoN
5lKdrUIe+jwZGU8GYjO4iZaAzh0DhEBp2B4No79wGpPzEYA8ExhDcIo1oByzN+2T
FNdPGWueAiKOV5TBCGc48v9DQHWrsVyDrpyy5+hEnFtv3E6GvUWGgbkOZ6XGaqdm
7DZ4VIz5pgg2c3+4Qfk9JlTh3Z0oM2TXuLbC/kjfACF+1KGx6f/Aane7sfgGxao7
VyV3lT5NFTny4Cx6B9lJjqMNI639Xsez69jWJwL03ZmkSZpzxnAoFEsoN7/nhVvd
ShCYoMcMi33o4VfTdvz0v3v9T8RUEKWhCgm968lbiw7tI9d7NL5W34BvZZQEtG2A
7FUPVMTaezGHOCe0qzCzuHgXYt/Sa854L2ueskpiosBLjzq6WaeruZKjfbf7/40V
USMryteFDJi1glGtORV9SwPTrCtylTUOGGp/RPylbcUJtCLa+1uCCnz36GqYAqcR
vwDVHLlWRmL5az7KpG5cyMk4LlIBu2Gdhxxd3qnETbiu+wYTzqfqgY0rTULw4dcv
eV0/Mg1LYVbQztYlH63mGPoUncxetnDaIgXQ9X5N8sGbbO4xv6RK7doknfCKOV3W
JQ6Dwqnwm3fbgMdHxNyTcEStTvdu2yfqalQy3BLazVk2Hc6doqOFJxASzcDSlHXt
vm4VD7L+23shQLz2YVTyfl2oDnYmhFYuLMLeYE3IKWMeowACfGTz1WyE+/GLaObM
i9JzRxgTyeSwkAVBUpsE1FaUFtGESrTAuj5EwwrjpQFksPArMqpRvC/DqKTTB2MF
3mpXDgtzKIZVLcA7QJGUcbjfoChPfhvNMVbB1bGPInDKfWAQ/MNjV9yBkFhUxBMg
KuS64MlTdB19QMskHxJT+V4GdGr6Q3FSk4EJQjO27rZJQ4/zWQeSl5za/69am8Sj
/fu6kQE24TSosseKzZEBPKKZB4vRKppyuH9qjoYwiRmrcfm85fNDS8dFE2BajqEW
IhyVoz5k1McgteTD4Tw37ntUVYFXvSR/uTCoggnniI4UIPNP8iw90R49617oqGs+
PqsbtrSet6XL5hWmPqUHh8nnk9cqhR3T33EstTtMrpD/xIl7H4f4y6P2P1yFNPDs
1nkks2asiOBoQRBOwRCVZGIZHJLO3UHSGYGd2fcowb0K+72T2FI8AZo8X6bAaGqZ
NJhJ/Z3U5/Fahh1oKMj0KbV+mZUYQBnhJl7rhVqNbrjahojFFAg/RNCu1TrTqHIw
aT5vcWwktMAUkL17lVS74VbH0bOM9naKb5Pp7lYV3J3pY3TxIk08u+EICxJAcvME
Re59SZRK8gGdnqBlw6rqN8RwUGMDwbUUOsA9aWw/b1kUCXJJAOALdRvRB1XPJn5f
0+Bv1Haeo0vPTC0AFAmIkfprHtOn0E1p5fdEjOMbQ16bH5GGe4URqXCg0y001bG0
y0k1Cgm6f8SsA72UCWINLbLnMAAxec0wCz1aApfhZ4eV8hF50S0AptpKBE5i4g1F
0ctaapxkYDckuULGrgkZwXEEvVfkVG+S0fMmbpFWQi/IkD9j6zLUN4tl3/5J8hN5
5m+AcnUmhPs7W/aaASi7VbCyHkfp+ghYeFWRdQRCcoxbUl04BlapkOwPix8vzU/T
sg5Qx0ZZadVWyAR9WEpMRQ2E/2e9/Z+DgNXSlfFvUfUAyISXFBQrJMDT4HJ8nHZK
hVbOr157kIs4P2O5iZN2F7V6YZ/YL5wsyJ9LGHSplcLeBddtGP35hXpY7tHHViSx
rfVkkky3SXfjjvK4iJdOBN4vkTZD56lCccufhKZSuTndXobj2XPLaKUIn/rscKHF
G6wB74wH5fkZEtiwAJ1RFpWoZKyck0+dJsOnb1O+bcLhVdMwWE0UI+LXKH5Pet5I
AFhhcxr9KWvJppHb1kHK4uZeAKJuAeYlSu0Ocrer1r7Qo067sIR9YjMDh92JM+zn
rwwv6HWeQpagHKT3+o3tST/KFh9JA7MN2D5LQJsUcRMc5dvr0MsJHMl1TgP/mDpd
wcJ2sggimUksBLwhXxspAkRjYcSGqmKvwXzfFA5Gr5voijS49v3eE+MYkBBcRZuA
fhv3PNykmTnVfeC6dZ2dznoRDcRcbEGv/NmHmoT6l7APrWpK+DgMPMpLsgti8L6n
qWV5ZLJ/iWJO8Hr69A3fSVWPwsAjGt9zS1zQtB+rdPqTAXPHRYIOecLU86Sqsy9G
0MmKPjFrBzMyleOqhcAOwyh+IhDdH/htp7dUvedvllsvrrC3E80I0JTl2D4s65DS
wOim2InjQYTqsmqJBJPsgQVqxdTqJrgsNl2E7y7ukesOqlqgAls9BSQKkd8Vg665
iPj2Ss6u4tPou6pV/kiwP+WBS2LQSqyXrgfV9HME63OkeYX5vfbVDqXPsyR5YTQT
qSc+WQ7x5J874aFBp4mNBGa+tDV1V1oEuR7RSkHlxFMpBeTksqq7QdqmyCXtzLYG
JddHFo8h8JPomC6c7BZD3nlewGwRRHZfMbOBIR40UaS5RSE+FL1xRv9+NQ122Pn8
NKtIXy3NgnsE/akzDvtijhJCI73vTmZiuD6fPBLp8QPDnaIac41KCVfGKYFUv5kQ
wxQjUdd9LqpZAdov15mxETath4uY8uoNM85oCibZaPSAy1L0zw/ZliL93IZHbRqd
yyQ6DoYoU0j7WUPe+wEJQz+aqLZ7EmCRm6nfne/GY6BDOCCoUTq4roNEkn4glBqW
sJcD9bxEmoc5jHk1fZEdwpFTukrn2LcEB/TbhSsvjrVUSGSBzxvTH7cgnwkTSrTs
YRU0CA1wesxzjXk3z2BiWSbTsmMWqAY3Od1kpockaL4xe6FuMfLSj1jSXiYjuqgs
I2MdLj/8IfA67AHK64NxtWA9L/YYhmmgeOQsVScc3B++Qj6GO4RoU1wbia/+T/l5
/xaQCixw9MgLvOMFqJ6uXmIK4mUH2AcVzSBThhE0TP1HsGrNudeg/LLUL8OVhH0f
DR9OQVcnUlolnvKi+tnd2pZULXOI5YOmpCEt8RF1MtF7V3kUVNWjZ8KrvhQDBofN
5OC924ofIwkwv/1NTkKXkTtOkkmqDjLBgEYOCbCtOfZIpo+Qc4yAkSa9Lo4UU1JX
jNLxl9vNF53aeMVVzGBiEXH0Z2w99E2XzXdUMU4qMlNS3yBmao4S8Z2vvX6n6roh
0oxvZvI8xTOGEYVX63GDN2iYgRj24gVNRQqEJmjYUwj+h2Jeo9sVCVWW+6Qq+Jyd
6Yd/VnXIj1PPvudMRf0bUvHvMs8ngF1+7WGYQ4cpRo1dHoatWYJqX1ZmbUoHOgyM
y1V/fmXtO+DR1CVccTkRHLn9WekwUIWSNPEOgaYly3CCJvUPIUhy74JYXIR6qRK6
xr3ilyvk2TqeJd2/Yze8Fx/p8OqoP4j+bDG+UnA/DHf+Y7ilqf8YeFLJweyCImLN
Cs+5PvS5u3a39ZfZRjCotTraswPy0Y+8rcPiYnfKK8Iku+TnPlHcXpAyeYdravM4
FiVebceE4aQ8uH7QPTi3Kj1vjUGvyGBgjVwsv2bDFczLPEFA5Z41eRjm3mPhd+0V
AeH0FLNFawTpTIWlovqqk/e37Og2aBdhFO5+ofU5DX58IEUVjYTuqb2aeWaL/so3
OvJFMHMR+jTNUuMmX1pNo6K7HPvfDZbslE3+Gu7gF1WHmMBb+wUNgp551pBS6hDE
aFLVkKS8ecr55GGx4pe4d6qytl+cWWb3/w8vPM8jRZmVcfjGUh6k9Mf/3Mp9uLTw
ULsRLkVYFwxkfZ+kanvhA6Lawj6AEZuUERC3n4eBKxpBkB0Af6R+Mjs5GZyJ05u7
iVfAMBZfv1utVqv3yA7TdAtemmpiCpIZdntbVxnbfitKGrsJUlSYO95bUjifRjHW
DZtHflcC/L9pjVzaGZxoGDNqIsnced79QNKXDTuVzglP1Y1Nlyc1Yn9Ji/Sbs9Rh
WGoOdtSx3duoz1l43AEnnnMTH1phlPxkbuggest9hTi83vox8R0mPl+IiBtBb91C
R/cI3Iuo4NY6MT2Fk8qaQ0atjFFcduDj/bBbF/0dRXBvEtc0eLpsQsk70ngQ/Srt
VPiDjyEjxhEHMgftjtVM9D5uENa2WWd0TT+ux3FwGKU0hwqbqKGAhllnbFJNfcGJ
wPLgyKXKmLRFvbco2NVBaLjlCFzXVrUCaHB4TAYNhC1MupwdH0TWwNp5Tu+lUPcz
eYIPHgqIy1oyA9TRwIui1EpbrKcbzqsi0z/o9UdPMwUGQkuU0SiOVANubO0VHq3/
VY56sPY2nuwMz44bRVXygJFvjUUNGCYn6S6DRg+ocp6/DeBK/+TryfdDTagjDneq
DF/L2Ao8xyGJ6stmys4+OZRN7i9zSeTbipfp3jDbr7bNUExO9rEAQOjAqi1VM5qW
msFx3Rih1NIOIGF+0t6bXg7JEAvK0hQW4LdKb+PA4mAlhCbtkUl+RMMsKeryKe/G
G0M+UAFyUne+wVJVmgY2L6zmCXUIAHl3AZhKU3zMODXgFcUT87+Q9taj9pQta8ji
EA8a8GSFpd3tLaGriEC3/s0V096ecDZIXwbtyTfFeS01rL04yzxMw3mB3EBp/Dpv
v/F1rgBshcaQeDldO7h2p3pk24I8Yr7yZNLGoUIjKY5C3xY87gv1FMC/942JDkF6
a7rZnArl9p4QbnBqT2AxC+4BSWjflIINrXPEmZK6g9ulk2sybfduRkzrfkqdQeA0
UIyFScrXJ9JaktYkd2Z9hH1mQrXBo6DZ2NWQybYUsr1jHpPsiDZpmMmy3yoA/Zc2
Pv2pcL68MsawwxNmMYBwvvPmn3UisBaoKCnfJsilSVIlSuYsirCPBkSWpmkusBM8
+o/UzP8CjizcQt5P1rai/SGcq+O9AyJvlxbt+68DGW5wOYEPoh7U5B7wT7hPx5Mu
6j2OUxjsYiNW60QOdX02aQybnaH4r5DF2sEHlIevt/Up5Xe0e5NS/cgsJL1blnb8
VRtFHjARgvzmZJixYG9phuIMdUsgPliLqCtWibZwiEig2Sqvu0CzWt7GPdZDj4aD
3fvn60zc25AOS08cPCzhL5GnqhqUDaRNlClMXL02HYhKTTSSk7D4lKx9NLN/SGGw
XZCf/sR8TBeU2BQ3sGPd45VfxNn0ulYeZadNSy+Q22zH2h2YhJhIrjQd7j8/c1gE
Tsmvx9l+/Gh66tQcf5dYn/bA96XF3NBC3SwNZhQlevlS6IuB034Ek+XHvBJ7xt40
7PSL2ak4UcOHaUrQNcdgBQ==
`pragma protect end_protected
