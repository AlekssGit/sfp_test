// ed_sim.v

// Generated using ACDS version 21.4 67

`timescale 1 ps / 1 ps
module ed_sim (
		output wire  sim_checker_traffic_gen_pass,         //        sim_checker.traffic_gen_pass
		output wire  sim_checker_traffic_gen_fail,         //                   .traffic_gen_fail
		output wire  sim_checker_traffic_gen_timeout,      //                   .traffic_gen_timeout
		output wire  cal_status_checker_local_cal_success, // cal_status_checker.local_cal_success
		output wire  cal_status_checker_local_cal_fail     //                   .local_cal_fail
	);

	wire          pll_ref_clk_source_clk_clk;                             // pll_ref_clk_source:clk -> [ddr3:pll_ref_clk, global_reset_n_source:clk]
	wire          ddr3_emif_usr_clk_clk;                                  // ddr3:emif_usr_clk -> [mm_interconnect_0:ddr3_emif_usr_clk_clk, rst_controller:clk, tg:emif_usr_clk]
	wire          ddr3_ctrl_ecc_user_interrupt_0_ctrl_ecc_user_interrupt; // ddr3:ctrl_ecc_user_interrupt_0 -> tg:ctrl_ecc_user_interrupt_0
	wire    [0:0] ddr3_mem_mem_reset_n;                                   // ddr3:mem_reset_n -> mem:mem_reset_n
	wire    [0:0] ddr3_mem_mem_cas_n;                                     // ddr3:mem_cas_n -> mem:mem_cas_n
	wire    [2:0] ddr3_mem_mem_ba;                                        // ddr3:mem_ba -> mem:mem_ba
	wire    [0:0] ddr3_mem_mem_we_n;                                      // ddr3:mem_we_n -> mem:mem_we_n
	wire    [0:0] ddr3_mem_mem_ck;                                        // ddr3:mem_ck -> mem:mem_ck
	wire    [4:0] ddr3_mem_mem_dqs;                                       // [] -> [ddr3:mem_dqs, mem:mem_dqs]
	wire    [4:0] ddr3_mem_mem_dm;                                        // ddr3:mem_dm -> mem:mem_dm
	wire   [39:0] ddr3_mem_mem_dq;                                        // [] -> [ddr3:mem_dq, mem:mem_dq]
	wire    [0:0] ddr3_mem_mem_cs_n;                                      // ddr3:mem_cs_n -> mem:mem_cs_n
	wire   [14:0] ddr3_mem_mem_a;                                         // ddr3:mem_a -> mem:mem_a
	wire    [0:0] ddr3_mem_mem_odt;                                       // ddr3:mem_odt -> mem:mem_odt
	wire    [0:0] ddr3_mem_mem_ras_n;                                     // ddr3:mem_ras_n -> mem:mem_ras_n
	wire    [4:0] ddr3_mem_mem_dqs_n;                                     // [] -> [ddr3:mem_dqs_n, mem:mem_dqs_n]
	wire    [0:0] ddr3_mem_mem_ck_n;                                      // ddr3:mem_ck_n -> mem:mem_ck_n
	wire    [0:0] ddr3_mem_mem_cke;                                       // ddr3:mem_cke -> mem:mem_cke
	wire          ddr3_status_local_cal_fail;                             // ddr3:local_cal_fail -> sim_checker:local_cal_fail_0
	wire          ddr3_status_local_cal_success;                          // ddr3:local_cal_success -> sim_checker:local_cal_success_0
	wire          tg_tg_status_0_traffic_gen_fail;                        // tg:traffic_gen_fail_0 -> sim_checker:traffic_gen_fail_0
	wire          tg_tg_status_0_traffic_gen_timeout;                     // tg:traffic_gen_timeout_0 -> sim_checker:traffic_gen_timeout_0
	wire          tg_tg_status_0_traffic_gen_pass;                        // tg:traffic_gen_pass_0 -> sim_checker:traffic_gen_pass_0
	wire          ddr3_emif_usr_reset_n_reset;                            // ddr3:emif_usr_reset_n -> [rst_controller:reset_in0, tg:emif_usr_reset_n]
	wire          global_reset_n_source_reset_reset;                      // global_reset_n_source:reset -> global_reset_n_splitter:sig_input
	wire          global_reset_n_splitter_sig_output_if_0_reset;          // global_reset_n_splitter:sig_output_0 -> ddr3:global_reset_n
	wire          tg_ctrl_amm_0_waitrequest;                              // mm_interconnect_0:tg_ctrl_amm_0_waitrequest -> tg:amm_ready_0
	wire  [255:0] tg_ctrl_amm_0_readdata;                                 // mm_interconnect_0:tg_ctrl_amm_0_readdata -> tg:amm_readdata_0
	wire          tg_ctrl_amm_0_read;                                     // tg:amm_read_0 -> mm_interconnect_0:tg_ctrl_amm_0_read
	wire   [29:0] tg_ctrl_amm_0_address;                                  // tg:amm_address_0 -> mm_interconnect_0:tg_ctrl_amm_0_address
	wire   [31:0] tg_ctrl_amm_0_byteenable;                               // tg:amm_byteenable_0 -> mm_interconnect_0:tg_ctrl_amm_0_byteenable
	wire          tg_ctrl_amm_0_readdatavalid;                            // mm_interconnect_0:tg_ctrl_amm_0_readdatavalid -> tg:amm_readdatavalid_0
	wire          tg_ctrl_amm_0_write;                                    // tg:amm_write_0 -> mm_interconnect_0:tg_ctrl_amm_0_write
	wire  [255:0] tg_ctrl_amm_0_writedata;                                // tg:amm_writedata_0 -> mm_interconnect_0:tg_ctrl_amm_0_writedata
	wire    [6:0] tg_ctrl_amm_0_burstcount;                               // tg:amm_burstcount_0 -> mm_interconnect_0:tg_ctrl_amm_0_burstcount
	wire  [255:0] mm_interconnect_0_ddr3_ctrl_amm_0_readdata;             // ddr3:amm_readdata_0 -> mm_interconnect_0:ddr3_ctrl_amm_0_readdata
	wire          mm_interconnect_0_ddr3_ctrl_amm_0_waitrequest;          // ddr3:amm_ready_0 -> mm_interconnect_0:ddr3_ctrl_amm_0_waitrequest
	wire   [24:0] mm_interconnect_0_ddr3_ctrl_amm_0_address;              // mm_interconnect_0:ddr3_ctrl_amm_0_address -> ddr3:amm_address_0
	wire          mm_interconnect_0_ddr3_ctrl_amm_0_read;                 // mm_interconnect_0:ddr3_ctrl_amm_0_read -> ddr3:amm_read_0
	wire   [31:0] mm_interconnect_0_ddr3_ctrl_amm_0_byteenable;           // mm_interconnect_0:ddr3_ctrl_amm_0_byteenable -> ddr3:amm_byteenable_0
	wire          mm_interconnect_0_ddr3_ctrl_amm_0_readdatavalid;        // ddr3:amm_readdatavalid_0 -> mm_interconnect_0:ddr3_ctrl_amm_0_readdatavalid
	wire          mm_interconnect_0_ddr3_ctrl_amm_0_write;                // mm_interconnect_0:ddr3_ctrl_amm_0_write -> ddr3:amm_write_0
	wire  [255:0] mm_interconnect_0_ddr3_ctrl_amm_0_writedata;            // mm_interconnect_0:ddr3_ctrl_amm_0_writedata -> ddr3:amm_writedata_0
	wire    [6:0] mm_interconnect_0_ddr3_ctrl_amm_0_burstcount;           // mm_interconnect_0:ddr3_ctrl_amm_0_burstcount -> ddr3:amm_burstcount_0
	wire          rst_controller_reset_out_reset;                         // rst_controller:reset_out -> mm_interconnect_0:tg_ctrl_amm_0_translator_reset_reset_bridge_in_reset_reset

	ed_sim_ddr3 ddr3 (
		.global_reset_n            (global_reset_n_splitter_sig_output_if_0_reset),          //   input,    width = 1,            global_reset_n.reset_n
		.pll_ref_clk               (pll_ref_clk_source_clk_clk),                             //   input,    width = 1,               pll_ref_clk.clk
		.oct_rzqin                 (),                                                       //   input,    width = 1,                       oct.oct_rzqin
		.mem_ck                    (ddr3_mem_mem_ck),                                        //  output,    width = 1,                       mem.mem_ck
		.mem_ck_n                  (ddr3_mem_mem_ck_n),                                      //  output,    width = 1,                          .mem_ck_n
		.mem_a                     (ddr3_mem_mem_a),                                         //  output,   width = 15,                          .mem_a
		.mem_ba                    (ddr3_mem_mem_ba),                                        //  output,    width = 3,                          .mem_ba
		.mem_cke                   (ddr3_mem_mem_cke),                                       //  output,    width = 1,                          .mem_cke
		.mem_cs_n                  (ddr3_mem_mem_cs_n),                                      //  output,    width = 1,                          .mem_cs_n
		.mem_odt                   (ddr3_mem_mem_odt),                                       //  output,    width = 1,                          .mem_odt
		.mem_reset_n               (ddr3_mem_mem_reset_n),                                   //  output,    width = 1,                          .mem_reset_n
		.mem_we_n                  (ddr3_mem_mem_we_n),                                      //  output,    width = 1,                          .mem_we_n
		.mem_ras_n                 (ddr3_mem_mem_ras_n),                                     //  output,    width = 1,                          .mem_ras_n
		.mem_cas_n                 (ddr3_mem_mem_cas_n),                                     //  output,    width = 1,                          .mem_cas_n
		.mem_dqs                   (ddr3_mem_mem_dqs),                                       //   inout,    width = 5,                          .mem_dqs
		.mem_dqs_n                 (ddr3_mem_mem_dqs_n),                                     //   inout,    width = 5,                          .mem_dqs_n
		.mem_dq                    (ddr3_mem_mem_dq),                                        //   inout,   width = 40,                          .mem_dq
		.mem_dm                    (ddr3_mem_mem_dm),                                        //  output,    width = 5,                          .mem_dm
		.local_cal_success         (ddr3_status_local_cal_success),                          //  output,    width = 1,                    status.local_cal_success
		.local_cal_fail            (ddr3_status_local_cal_fail),                             //  output,    width = 1,                          .local_cal_fail
		.emif_usr_reset_n          (ddr3_emif_usr_reset_n_reset),                            //  output,    width = 1,          emif_usr_reset_n.reset_n
		.emif_usr_clk              (ddr3_emif_usr_clk_clk),                                  //  output,    width = 1,              emif_usr_clk.clk
		.ctrl_ecc_user_interrupt_0 (ddr3_ctrl_ecc_user_interrupt_0_ctrl_ecc_user_interrupt), //  output,    width = 1, ctrl_ecc_user_interrupt_0.ctrl_ecc_user_interrupt
		.amm_ready_0               (mm_interconnect_0_ddr3_ctrl_amm_0_waitrequest),          //  output,    width = 1,                ctrl_amm_0.waitrequest_n
		.amm_read_0                (mm_interconnect_0_ddr3_ctrl_amm_0_read),                 //   input,    width = 1,                          .read
		.amm_write_0               (mm_interconnect_0_ddr3_ctrl_amm_0_write),                //   input,    width = 1,                          .write
		.amm_address_0             (mm_interconnect_0_ddr3_ctrl_amm_0_address),              //   input,   width = 25,                          .address
		.amm_readdata_0            (mm_interconnect_0_ddr3_ctrl_amm_0_readdata),             //  output,  width = 256,                          .readdata
		.amm_writedata_0           (mm_interconnect_0_ddr3_ctrl_amm_0_writedata),            //   input,  width = 256,                          .writedata
		.amm_burstcount_0          (mm_interconnect_0_ddr3_ctrl_amm_0_burstcount),           //   input,    width = 7,                          .burstcount
		.amm_byteenable_0          (mm_interconnect_0_ddr3_ctrl_amm_0_byteenable),           //   input,   width = 32,                          .byteenable
		.amm_readdatavalid_0       (mm_interconnect_0_ddr3_ctrl_amm_0_readdatavalid)         //  output,    width = 1,                          .readdatavalid
	);

	ed_sim_global_reset_n_source global_reset_n_source (
		.reset (global_reset_n_source_reset_reset), //  output,  width = 1, reset.reset_n
		.clk   (pll_ref_clk_source_clk_clk)         //   input,  width = 1,   clk.clk
	);

	ed_sim_global_reset_n_splitter global_reset_n_splitter (
		.sig_input    (global_reset_n_source_reset_reset),             //   input,  width = 1,    sig_input_if.reset_n
		.sig_output_0 (global_reset_n_splitter_sig_output_if_0_reset)  //  output,  width = 1, sig_output_if_0.reset_n
	);

	ed_sim_mem mem (
		.mem_ck      (ddr3_mem_mem_ck),      //   input,   width = 1, mem.mem_ck
		.mem_ck_n    (ddr3_mem_mem_ck_n),    //   input,   width = 1,    .mem_ck_n
		.mem_a       (ddr3_mem_mem_a),       //   input,  width = 15,    .mem_a
		.mem_ba      (ddr3_mem_mem_ba),      //   input,   width = 3,    .mem_ba
		.mem_cke     (ddr3_mem_mem_cke),     //   input,   width = 1,    .mem_cke
		.mem_cs_n    (ddr3_mem_mem_cs_n),    //   input,   width = 1,    .mem_cs_n
		.mem_odt     (ddr3_mem_mem_odt),     //   input,   width = 1,    .mem_odt
		.mem_reset_n (ddr3_mem_mem_reset_n), //   input,   width = 1,    .mem_reset_n
		.mem_we_n    (ddr3_mem_mem_we_n),    //   input,   width = 1,    .mem_we_n
		.mem_ras_n   (ddr3_mem_mem_ras_n),   //   input,   width = 1,    .mem_ras_n
		.mem_cas_n   (ddr3_mem_mem_cas_n),   //   input,   width = 1,    .mem_cas_n
		.mem_dqs     (ddr3_mem_mem_dqs),     //   inout,   width = 5,    .mem_dqs
		.mem_dqs_n   (ddr3_mem_mem_dqs_n),   //   inout,   width = 5,    .mem_dqs_n
		.mem_dq      (ddr3_mem_mem_dq),      //   inout,  width = 40,    .mem_dq
		.mem_dm      (ddr3_mem_mem_dm)       //   input,   width = 5,    .mem_dm
	);

	ed_sim_pll_ref_clk_source pll_ref_clk_source (
		.clk (pll_ref_clk_source_clk_clk)  //  output,  width = 1, clk.clk
	);

	ed_sim_sim_checker sim_checker (
		.traffic_gen_pass_0    (tg_tg_status_0_traffic_gen_pass),      //   input,  width = 1, tg_status_0.traffic_gen_pass
		.traffic_gen_fail_0    (tg_tg_status_0_traffic_gen_fail),      //   input,  width = 1,            .traffic_gen_fail
		.traffic_gen_timeout_0 (tg_tg_status_0_traffic_gen_timeout),   //   input,  width = 1,            .traffic_gen_timeout
		.traffic_gen_pass      (sim_checker_traffic_gen_pass),         //  output,  width = 1,   tg_status.traffic_gen_pass
		.traffic_gen_fail      (sim_checker_traffic_gen_fail),         //  output,  width = 1,            .traffic_gen_fail
		.traffic_gen_timeout   (sim_checker_traffic_gen_timeout),      //  output,  width = 1,            .traffic_gen_timeout
		.local_cal_success_0   (ddr3_status_local_cal_success),        //   input,  width = 1,    status_0.local_cal_success
		.local_cal_fail_0      (ddr3_status_local_cal_fail),           //   input,  width = 1,            .local_cal_fail
		.local_cal_success     (cal_status_checker_local_cal_success), //  output,  width = 1,      status.local_cal_success
		.local_cal_fail        (cal_status_checker_local_cal_fail)     //  output,  width = 1,            .local_cal_fail
	);

	ed_sim_tg tg (
		.emif_usr_reset_n          (ddr3_emif_usr_reset_n_reset),                            //   input,    width = 1,          emif_usr_reset_n.reset_n
		.ninit_done                (),                                                       //   input,    width = 1,                ninit_done.ninit_done
		.emif_usr_clk              (ddr3_emif_usr_clk_clk),                                  //   input,    width = 1,              emif_usr_clk.clk
		.amm_ready_0               (~tg_ctrl_amm_0_waitrequest),                             //   input,    width = 1,                ctrl_amm_0.waitrequest_n
		.amm_read_0                (tg_ctrl_amm_0_read),                                     //  output,    width = 1,                          .read
		.amm_write_0               (tg_ctrl_amm_0_write),                                    //  output,    width = 1,                          .write
		.amm_address_0             (tg_ctrl_amm_0_address),                                  //  output,   width = 30,                          .address
		.amm_readdata_0            (tg_ctrl_amm_0_readdata),                                 //   input,  width = 256,                          .readdata
		.amm_writedata_0           (tg_ctrl_amm_0_writedata),                                //  output,  width = 256,                          .writedata
		.amm_burstcount_0          (tg_ctrl_amm_0_burstcount),                               //  output,    width = 7,                          .burstcount
		.amm_byteenable_0          (tg_ctrl_amm_0_byteenable),                               //  output,   width = 32,                          .byteenable
		.amm_readdatavalid_0       (tg_ctrl_amm_0_readdatavalid),                            //   input,    width = 1,                          .readdatavalid
		.traffic_gen_pass_0        (tg_tg_status_0_traffic_gen_pass),                        //  output,    width = 1,               tg_status_0.traffic_gen_pass
		.traffic_gen_fail_0        (tg_tg_status_0_traffic_gen_fail),                        //  output,    width = 1,                          .traffic_gen_fail
		.traffic_gen_timeout_0     (tg_tg_status_0_traffic_gen_timeout),                     //  output,    width = 1,                          .traffic_gen_timeout
		.ctrl_ecc_user_interrupt_0 (ddr3_ctrl_ecc_user_interrupt_0_ctrl_ecc_user_interrupt)  //   input,    width = 1, ctrl_ecc_user_interrupt_0.ctrl_ecc_user_interrupt
	);

	ed_sim_altera_mm_interconnect_1920_3ogrq5i mm_interconnect_0 (
		.tg_ctrl_amm_0_address                                      (tg_ctrl_amm_0_address),                           //   input,   width = 30,                                        tg_ctrl_amm_0.address
		.tg_ctrl_amm_0_waitrequest                                  (tg_ctrl_amm_0_waitrequest),                       //  output,    width = 1,                                                     .waitrequest
		.tg_ctrl_amm_0_burstcount                                   (tg_ctrl_amm_0_burstcount),                        //   input,    width = 7,                                                     .burstcount
		.tg_ctrl_amm_0_byteenable                                   (tg_ctrl_amm_0_byteenable),                        //   input,   width = 32,                                                     .byteenable
		.tg_ctrl_amm_0_read                                         (tg_ctrl_amm_0_read),                              //   input,    width = 1,                                                     .read
		.tg_ctrl_amm_0_readdata                                     (tg_ctrl_amm_0_readdata),                          //  output,  width = 256,                                                     .readdata
		.tg_ctrl_amm_0_readdatavalid                                (tg_ctrl_amm_0_readdatavalid),                     //  output,    width = 1,                                                     .readdatavalid
		.tg_ctrl_amm_0_write                                        (tg_ctrl_amm_0_write),                             //   input,    width = 1,                                                     .write
		.tg_ctrl_amm_0_writedata                                    (tg_ctrl_amm_0_writedata),                         //   input,  width = 256,                                                     .writedata
		.ddr3_ctrl_amm_0_address                                    (mm_interconnect_0_ddr3_ctrl_amm_0_address),       //  output,   width = 25,                                      ddr3_ctrl_amm_0.address
		.ddr3_ctrl_amm_0_write                                      (mm_interconnect_0_ddr3_ctrl_amm_0_write),         //  output,    width = 1,                                                     .write
		.ddr3_ctrl_amm_0_read                                       (mm_interconnect_0_ddr3_ctrl_amm_0_read),          //  output,    width = 1,                                                     .read
		.ddr3_ctrl_amm_0_readdata                                   (mm_interconnect_0_ddr3_ctrl_amm_0_readdata),      //   input,  width = 256,                                                     .readdata
		.ddr3_ctrl_amm_0_writedata                                  (mm_interconnect_0_ddr3_ctrl_amm_0_writedata),     //  output,  width = 256,                                                     .writedata
		.ddr3_ctrl_amm_0_burstcount                                 (mm_interconnect_0_ddr3_ctrl_amm_0_burstcount),    //  output,    width = 7,                                                     .burstcount
		.ddr3_ctrl_amm_0_byteenable                                 (mm_interconnect_0_ddr3_ctrl_amm_0_byteenable),    //  output,   width = 32,                                                     .byteenable
		.ddr3_ctrl_amm_0_readdatavalid                              (mm_interconnect_0_ddr3_ctrl_amm_0_readdatavalid), //   input,    width = 1,                                                     .readdatavalid
		.ddr3_ctrl_amm_0_waitrequest                                (~mm_interconnect_0_ddr3_ctrl_amm_0_waitrequest),  //   input,    width = 1,                                                     .waitrequest
		.tg_ctrl_amm_0_translator_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                  //   input,    width = 1, tg_ctrl_amm_0_translator_reset_reset_bridge_in_reset.reset
		.ddr3_emif_usr_clk_clk                                      (ddr3_emif_usr_clk_clk)                            //   input,    width = 1,                                    ddr3_emif_usr_clk.clk
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~ddr3_emif_usr_reset_n_reset),   //   input,  width = 1, reset_in0.reset
		.clk            (ddr3_emif_usr_clk_clk),          //   input,  width = 1,       clk.clk
		.reset_out      (rst_controller_reset_out_reset), //  output,  width = 1, reset_out.reset
		.reset_req      (),                               // (terminated),                       
		.reset_req_in0  (1'b0),                           // (terminated),                       
		.reset_in1      (1'b0),                           // (terminated),                       
		.reset_req_in1  (1'b0),                           // (terminated),                       
		.reset_in2      (1'b0),                           // (terminated),                       
		.reset_req_in2  (1'b0),                           // (terminated),                       
		.reset_in3      (1'b0),                           // (terminated),                       
		.reset_req_in3  (1'b0),                           // (terminated),                       
		.reset_in4      (1'b0),                           // (terminated),                       
		.reset_req_in4  (1'b0),                           // (terminated),                       
		.reset_in5      (1'b0),                           // (terminated),                       
		.reset_req_in5  (1'b0),                           // (terminated),                       
		.reset_in6      (1'b0),                           // (terminated),                       
		.reset_req_in6  (1'b0),                           // (terminated),                       
		.reset_in7      (1'b0),                           // (terminated),                       
		.reset_req_in7  (1'b0),                           // (terminated),                       
		.reset_in8      (1'b0),                           // (terminated),                       
		.reset_req_in8  (1'b0),                           // (terminated),                       
		.reset_in9      (1'b0),                           // (terminated),                       
		.reset_req_in9  (1'b0),                           // (terminated),                       
		.reset_in10     (1'b0),                           // (terminated),                       
		.reset_req_in10 (1'b0),                           // (terminated),                       
		.reset_in11     (1'b0),                           // (terminated),                       
		.reset_req_in11 (1'b0),                           // (terminated),                       
		.reset_in12     (1'b0),                           // (terminated),                       
		.reset_req_in12 (1'b0),                           // (terminated),                       
		.reset_in13     (1'b0),                           // (terminated),                       
		.reset_req_in13 (1'b0),                           // (terminated),                       
		.reset_in14     (1'b0),                           // (terminated),                       
		.reset_req_in14 (1'b0),                           // (terminated),                       
		.reset_in15     (1'b0),                           // (terminated),                       
		.reset_req_in15 (1'b0)                            // (terminated),                       
	);

endmodule
