`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
HGbDbPTH5xl8JxohLHftYIPGzACSAkCdcXnSDcZySu0fj7m88PXJBzUsjPBXLM5m
W8YoEQGknKKvxTWicpaD8sq8r1SzdCTrlAseKR7v/EKgpnj+2wysnxbxsJRz6AuD
rOGJkwJFk8jTYoYjJYnXiVLZfysL3Oywx9jroveFbuk=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 5168), data_block
OsXZl4U1gRDTYpSHX03hWh8vPIZZrwD3bBdNIGzppOiCJfLwRbGIdftMwxuboE3f
EPFtMT6vJ4SWUTDIADck2ZKZWFgX+meFMDdvxhDoOoOEjdM/8e8MSR0xaLi/bUf9
PqloJiTiR8YhCKuQv3oUdRVAz8rQtR4OVxKx5AyPlHTzT5rIYNZ+cl3XG+j6llXG
ObDy5epf/Sgo3HinYGYZmJyY24o3TSUunszcUAmHHcQN70bSOO92Y1GCgbTylFjb
ckvLfAU+Z002uFlcuefvPvm+wVS9flQp0RRq0UiEykM+Mu8MG89FBVkoJqcikk0r
3+5F5pWADpEoXHUhYaRDrNG4ztc/1TfE5w/WWH5EOGJa60JymeAzeroM+jhotLCg
h46oQwzHXEHI3wwfmoeLvdLDdPzoiqrVMz0T+1jlsqUrdlAFmUciEO1TgWSx/Xsu
SAoPH7VVwgT/VKSuIej6kQoV+e/K4dG1eylcDidMV7eba0pbI3OJ/PPgGrXolaj4
UxelAasF/QoljynwDf+YUP+bTewUBU3Jqkg+onub56/zez/4YR9A1mYlnTOGjurl
zA9AnNaXia/QMqvTx/RF0hbARcaw2YvlqsHtrodTyLSzlfyHp/IAhSKmDyBEZfse
Ye9zJrHaEWaVDMIbGWWupyjEOR3vaU1iDRBkpX1h+n+kU3b/LjVtQl/C0t5ylLtE
FSkXiSZT+jqmTc42oeTt7nlNcDMccMMIPGGKXNGwbjgaTFlFuGVlZHvx6Jds31xu
Yuf9WlzmAa7hwN64lLJsLa4jFJVHg+ixztbXv+DijRoMU9DofjzkDl6cKYrId5Vt
/a/R47Z23d+UKB97o0GZwBH402TeIOlxZ8mNlNAaJMe366v+HQchj9cveL40gnxg
oNXzhyRaDdFm2pSckEauddr9Bh4bL5gArrQ0b8UWM/Ig+rV9UQ2C5w5F/KzJ1r3X
f70smnlzTXmIpObrehOBHmpmfIUFQZLqTP/7i1fZLNkNoVvYrSOFCmLiMgpYypFn
YiaB1zPcDPoT5QD3epSGXoIICNss8mQ6whhxeoXCvi1rBUcE3dPoJujrbRnqvNTS
yHC8eX0Q1YzRO5E1goxOTAvb4v8T7tOmr7f484x0NT0rXtIoTM7z5yv5FYrUJKNd
27JgX4tXcgnGseSx1nk2rRmCCUpcyh6QTbUhfPYO8bjC6slysdf9KBh/UnT76Xer
eNo4wK2QIYYJ5P70cqNJooNSsQijli02NCXipNdvjqHMrXzOw4WfQ0IrADwTn4GI
aupUnM67iWB0IJqaplK8g6q5TlWlGeABH+aLjfAcw0UBQ9XKWzxfA/iHvnYzvTii
r+VdPvg8AdsKko9DsWyDTqEBvDDYcH3AaHzuNwdhzC2GxrOlouvCv+becupIT1Y0
f60DYUWV4iceO2nb9OdZiOz5L+1e2Gtu8kaYJNF1XqlVUcYVJuc6K3KIXM/tncoP
0ui3S8T965vxNNInvbns//IOXjafOBBhcHuBiaC2rQ3MDgpYGl7pZW3kAx7EDMH3
gxs5E+oPCUqPrFPYKv8ZpO3mjeHsQq8F7QpYRxJjUVpFeaf7xi5gXwNKKpHIL0KP
cXJZK+gyF5DVz7FtNQKHY/t6t02JokRWkEd8b06nx4lOQzitdfn8uQfFR/0LiPz4
Lnbpbq4UWLrIMjvMky30FmvLf0qa/xbSxbWr06LKTQOd7z8O6Hln5FfvZiJcRsaQ
t8tm45HwW9FNPLHZednj6mLGqdkBRI+Pv6+VwG4U0Ae5VOnS5O1H2Z9JTxs3IdeE
AEjSRHHXokk3E0a1w7eO+Y6Pew0q5A7nwCzSCzf87yPigwVfhQvPMt2JgK6NCLdo
Wx1asCKhvovPFRYlZpadHwSQyEJl05R6hMRkmZJArTLWH8qza/NnJ/r8KXRKgMja
wZxDqLfZdUtSUVXBfuOsNGt4/LIXbKCWCPeMryxgqqmyJPgeXNYV9aVfSZRKjSDG
fKp6PWfBGhjwGY+ge2kmahdRPap6XHcS8BHuOwCpSkaVUaxqA+lPIOYdTaWDtTG+
iXYmtmCq3HcJY6r00CKQVrGxV27oSaXk+B/9L+pnG7wEoDBzEHAD0sY/2EiMNVh/
4CSwS6dLi6UTUsg9bUd2nnbMBF4431OCfW82PHKDZRgw3PT8JhGCQtthFWIrOu/n
zjBj26z+ehCi0kPuMs4+B/ETJFXj4moIH50oJF6JCD+XBBer1bnnnGxLaMNn1FLS
mcg8Nua0lIsFXNo5QQn0Ilbg6DYuVGRCTuQu6dI9KCiCm8jsrBcAFAXdCxP2rpxW
qWV46gsMOmmzcwVKArk1dxXPSD69VdoZxI9Zj5kCAVcAh9up66V5PCK71AZbVpej
oiA36YkD127YqEZKXXD0wJVPrg6CG8xkMdXINFOnPVEKPuX+k2bb/ZWjcjkLvYg0
qSCbJqzCxaLxVWzMzsSSEp/+rra8TWlWyc7jl1VvIBH8eBATT55Byk0/1yTkGzti
NBfp3s00wDiIRpsdUR/HCVu3pmKtVRtT84NuBGYC5p3pHE5a3zNgogpJ9fQIUFKb
KPBoki4+pQSLGBeWwHqBXdcXjAzsWJLl4RQ72EHWwHl9E+TyQ7xix6j7juFYd+Uw
Keba/RM7b/hePQ3pBld5BQnguVBFXgnKRrY1tbmCSDpjDoEUArp5/9HfXBaY+xT7
f+EOnWfrDDCaw1Xfe3j4OfPMRWlq/RvBKGjnLPtwSEhp29OZvG5QaGOy/BW32lae
KzgveYkPTEknws9uCr+lV7Ziq0/NiYg1PwUCnxh4Wtx3kDG/g8vf4ZHvX8SuRTXw
JrnYVJzy/qiog1RaMdji4KOY81bifWodWJ94dLTjOCZhUEDqY5Z6fkTnLpMAD8Gm
Np8+h7+/C2ilkE9XliniIQsH4VTJiCNK2O+1T7HQDUe9Yhl84YFq+dv8eEzPQRuS
qPKHA0AJQYmk3gw0r3Fb50zNGPRhGqihmFRxDhKYD/SxL0ZJjOUqgv31A8AXOczr
fwU7ApF6HRzhuGON69VemMmkWe/zTNvW/mNkdtGLM0YAO1+L3k7oVbqDW6egDLFo
WAjyGkQR8QktyVmAvYp1t/Awb02F6AunvCvZuJ2V+5qxZjxOGafvWMY2jnzu7nmM
jmloXNW8QROT4vjww56PE6FZsKrRhRrD6d4nMVkoN3EqbO2F5aH5MuP4v1AULk53
9sakHFqEpiwq7uO1WKv4kS2v6C9LNgCuBx4F6Qp72PUhgdbR/sEdwoecNFpWkRzo
i+H2+9QJAfaxjmQMBtW86jyRWCSSzMPzKoAhgYhcPCyQkYS/S1Vi/DZYIkra38ba
7nuNaEIjxWbS1zdQKCWicArlW7/bKFWRTAnvf3hxcjihkHRxMhVn3Q41utzM+yHH
/UujPxYguabYz2t1AUYEzUyGRkLwGYW44gMbsMOvorXfFeSPl99/1n40sXKmOq3/
pxoiSTEuYx1CH0rKtKxCD+/lJUgwr1DYstzh7Mnyw0RRZ8IMPMQtuf7CRHWQeQLx
ztWnhmUtdfrzdY7znBqiNjJMjncio6lL7jtHgecNbdGO4Jr+heyg4pYH1qSb9AYq
02rp3et6upMTEa4y6VhgxaMOJ7ckJzCXnVX2kJxWbKoONxDZC7sKE9h0SA/1q9P4
nI3CufUZRAvPAsX8MjL1v5V1ClpAlacinbSniqKxGMseJjQcPbjpCCAH/KWvtVFQ
uJtcdxgn97qDc1nJ77NH96InJxh/Nyeb3+CVBAsfzVaZgwOCYCo7LbRZ4988PCI1
UojlWYBs6B4pp49EbRc1oO0q+zbIcc1rGSwsKUoH/qhiI/ZnWfZLuUbCeHHx91AO
IWW8myr3qj46tnwy2wkAnE0thhQvS7leLPcHMCUR/8kkEYy+jUB5wSXGFczh0dke
KJySWf1/F2tXFF3+fInsLTYMFmChCTyp7nbfJP/sp2/s6uT9O3XCy0aRmlKNeI/m
KrTMITuowqRmiixC9STQfeWtv6SBfZy0RLX+pmHNOVwXyrMTogAmBVJeXDPo1oXv
GVrUlLl58zG0yZYwOkHN6fFvo4DxP4SstD3SI8YPr3rtyBXqNfghZ41JtMJfBWnI
taeyotf9c2WKDmEpNheRqf6uiM8wX6RG6IwA+zG8Zlc0SnWDyyBA7E/TSEBG5Omh
zcCqWF18QnCLhEjlK6yi4BQ9TFwYUJLM8CPQIW84XgtzMKbw1iok6M+vGgqc+pd6
aapZZJgUu1Zk1Mz2sB4FgtavKTNxqE+nF9beekdM1LPFsNd5V3AXafdoPWDSPdht
mrVjoOQfsi0fjro/XHlVo34MpGoFPIJz+dgtGIVtw+hwKuSNb51ftZFUSNAxaWIZ
znfcTFndoCdvowMjODVkbcptCz8k8N1wcP5gLLYweEPd0fC/0Z/62KbBzC1uS6pQ
9ZNq9BhFlxLJUNLK1WXMbhnQKGgeR9dWdZBTCoeAw8RgFb7yJgyktqUhmovB7/pZ
61Kbz9OZ1LsOJTehGvypM6FHdGVkO0dWfQeu1uZN5McMoytUR3yGP0sW383T8nt/
4HlUlSFCEZESae/s4VdE+mxCo1OmIs7C9YRTZXV6gsbg2SFEngky4VgtrTWsL5cL
4aoNJyq/718xzvdZXoPCZDd/FpeAIkDaFmYbSBeANPcIH6FCWiGZaq7lsPL/FhR6
gBZwpTht/Y9rgTXYCRe7BE9G+Z/J63IbPw+B2P+BcEA5oTlkawsed52GT3CPE498
wb0BW6NbGHtYIyg51Vwgltr4wp4gtSkL+HfIhUESvPgoaRJg5ZuQ/38Ns/XbF8+q
cjVhPu/QrHVRaUXxFhWkWepy+JMho3dU0pNtUGy3c/glBq0pL18miXv+YK1STdHM
EsmJ6Av2//llgtId7YFDkOOCsB2T3Zk28DClSBa8KCdPrzI+2uYRcVPxRkKrGk8B
fxwsyGcPxAZAaZ1RxuUbMw21Nn8S8YKoXk94sKwIcE4O/WYok0mRyIPmHQlCmwOp
WAE++BxtNMnpdYwmJnVxB/G2LRt3YV0MkRlaHfGOd5oBLTmiFAlD/zJ/Nbp4kTIU
H2lCrEQGnCF7Sqq08sZkAEvQBCVYREIqbJR/Va5nreFDMEJNvAdBgSJdPGTgjT8v
1rROQSmGUTHzjecj30HtQud0+chuJaROLxl8gcwlARawG0tQjm8z59EDTl62Acfb
o/QNN0jtIsUTPAeGo6Tv5vO4LMm+88RLzk9uB568jJVttJJkgIpVOzfCr3OfJV1H
f0PF4g9jZmfskF7xLsyG/uRrj1HNkIRwODvtC8zf3XQZC5F7rrqsQnKmX1/s9ham
bv9cXcHsZKrMgR0WyHDod0GCcz2Q844sKGyzJ6CvBXMo7JooMqFgrVMBD03GtIBN
TBOTHqDvxYAIoHrkd4xjJQhJlpYybA/iUDaD9UYKQiUhdLjdwa+/1jHcjrx1+kG/
bHWTOGmK4SllUsPZp5jBCYd0xODA/0Cmff9In3WI0/ikzGWbyeRO+AOMw293QKh2
1vxm4x9o890dR0E/REidIlcKRTrMiCj5INEevfCo/IQTzbyR9qsRhpESik9QTmb9
1C/eqvHoqX7g5RJ3WlL7ytIdzgxrVxaJZcj1dIDOMWFIyzQsi80pwVJL3Pnxqpso
0152Y62HFJ1OMZqDtlQKSnPhoaIUexh2/iCHdplWK/OGgpuNsCk6P1PvdbqRaL0Y
K9jKSRxaJFoS68aAYMQTYjl3ObW9+f+wQTuSIBSqAPaPLJG3+l/JM13Sj+wWpk8n
eqEK6zKpE/ZZuvojOzG3Ip7vxay8+lIshTK+mAWPo0LMZbN/0L12C6OUa1iwbShb
aWWjTDdHso25ZF1aatC+p6F5tAFNPq/5EmkQq4GrXRFkrWIbp5vajcKKl+JBCexp
GgXOAhvBtXX+Ys3H6Oaw8GfswYZ4lVHWxkbNfscL5a/rXcp9tGjX7SDxPxA2Qa9F
fqsyZrbBTzWJs2KHCKXb3ghPh78vlcR9DFIINnl+eCqRNr9rQPkIs4TMqBJL2Svk
Qsl4nVGZGHzXsU7O7uYQoCNWJdA6kl+WIY7WejnZs2TLhTPi+Vd6+Yk1Z5Z6wqe+
NSjgR/HQKKENGJOCKxJ77hi6wwGF+ImCSALWjNimI16uzbc1gkwXna2PejBBnqmb
uKcLkmKtuCrCFiE8jhEoI5swoBvLsoYDfrg17txD5+lqvs2Wm7w3yE2dDQbFM8qq
UUm8MKfu6bPXKlYhRBhyUBRcYuUNyrinYufR35rtUYRhRreO3rS/qAn4OzCnUhtD
DUq4z9+O2JLJMlMVdIeAFY+xrtCsv4aBt9mBECLVVkVFRiI+ljKC1K5bQC4HRrt+
cb+z3RP7E7ULXxRjdPocRbbWVQ6rRlujo9hN8TYG9DUhK/4dNrEYRlxxEPyux7o+
oz5OMnw40OcIMfwKH7JBixOhgO30/m1Zavv1fkzxOmJ9lWNVKITCIg91tbBn2akK
r+Xq6alBXSWZxT1+T37GbDahTxglXvYruHrHIzHIKcNfrFBKcIIZzNrEDNu0VIqR
djCu7HeCv1wYUSzE4luKUyMpQdP6ksyAMuBuo3PTjfQB6xX0vs/Cu9Z/AyYNqI3d
3fuhWN8S4BzwVwhKKXurNIAzQK1uxWeiHmUbo21Wq5A+xFe2olcme6LHKx6ytdWi
PUXeX7S38blHZbHiFjT+AH2/yv2PLbidAHRE6XGB148RHAK6CV5luEYj+1nhrttJ
TOBwPcz/Pzrwx36aWREJTemSPCN8eXZyCb3Y6K1MGlwwWX79Pmth5boYR+UbIadF
d/N6sI2aYbQzW5aa//OOHlnjL9f2UZd+Tlt80Nw6yw4wR+GjimYDZmRoMriqcrOF
iJisgHHG7kraN11oCtZPV2k1SRQ/WMkEeC/Hv7b1Ltc=
`pragma protect end_protected
