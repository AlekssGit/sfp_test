// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
WCnO4edaMxELqhiY4fH1xBODnBSQD++xbCXgNwOtepi+ZfG4RtVy4S/+g7oIqh92
MrUtbGBKM1fhlIqshUs0d77TexLly8XtLB7WLfF/+t0HxHXRzc7kh1XFIyY+PwoU
2CAQYdD/EwH83nZW/RRZeYlgYjaUZh/b2ls81e/oVvc=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 5280 )
`pragma protect data_block
lySsWLJ/AEP/h1N34Xo+FVO6eZ1tLVJkNABK4o6a/f/rdO+MLgBJDGhmg6QLHnNu
lPbQ1wQPA+bNxbUH2sJEyreuj7vicy6VKY+FS/MNcQfrgfw2ZDViskY9i08qVxZ1
vDLo7ejyqWUn4jc4pCGmDeN3NqJA9cuin1axC+bSMJ5ZOoW/vkHFrZPjvY21sSNq
dSfAJwdPJl7Jy2sIAXMpLe6QQoWTeNRC1QNEwwJdjARYd5y7uy7sJ0PRe2aQy7as
kiSlN1M0/y1gSmgF64V+yeU4lo+XRCFHUPqaAC3Yxxt7orBniDJqQVHK4MHoPJwj
GwQEU9B75pnnzLdiDMBSTLuBjqzez0qgkHwwUmJT8yzZHAdAkUIcbvlcWR9T75Fa
nx/lyEVFvRFKZ0aNTlT/gZ8l3EykLIwWytrCHkiDexH9353xTQrjJ5G8LkapUaFM
bnT88J1SYGTxH1UmxD8WxyRfPAWKR/o0Kv6Ctc5XTCUwXfhizqskPUaeveOoyzOr
6XRjYo6f3YDTtER1a+s2TFHb0+Kibkn8faxdsbtzgMlw2MieXSat1k+r4nH8JS+2
opwPut+Nv6NTtBGOBooegTpxDElKgU1smhK8/+5Ty7PT/Gb96hMzSeCkkgjnwWGD
tLiBCpyyKz0Srf3n3AvE6Upt2ActMMrJ0x29BuHZI3LkfP6/MlqdpaR/gCQxpedK
cK7n5fot8QKCnDH+nKDjBVfQIh9Ohg6NmacyvbsC3STguAvjKuB5xKeanIV02VnG
AJL6XQXvuPBmgUGd1qQQ16goCngZLhuK/QekCoHozG9kfHjcrZUcQ64hkEdn6mNu
5G/5eNo2UiY08kRleKPbM/PGfRNnbHaU82EBTVmQnvO7X/lK4zooxah8lYDjOaV7
Ne6svq96S3/SeKnhU3IL+qaVZ+JC0AmjHYcpSkmoWIpvNEet6CdwD+g5n29t7uEz
qfCWlSiYOKgzQqFsDuUmfDdEO+KctvV/hBezK8X3pMbArDNpBKPECUt6Sb4FqYxH
8b4DURRwKhDbwfIxR7VK0IqBlcfF+SKSzYKiOfNpR7zXh23xpTxC0Z89tmzW+3Pl
cHIwQji7LGxETqyocJ3dP74NIEqpBSFc9oRi3FICwIej5dqTv52FggnwA797SHac
VXapPtFu+rWWBQi0MHiG9N6UgSLx4DD26QQqPAKB+u6LXLsro8nz5KW7Q3we6Osr
yLywXEv1wjaPFk6e1KklmShBdbwXUNczcipUHDW8dtgCUvd20eMoT+xW0ueTqBlk
cGt1x0w7YlvxOqg+palgiJ03UzvH/iW/j5v0OVEXZFYoXHHL8rCagS0CbSh8lsRG
iZNabO/ixntv+bQYBey6/AE4rxWOj2yTTKE2OnO+BBwGxVC5g/ArTH6dpt7EyUcp
codmsy+ynStD/jcYhWdlGJPROaFg6+PLXTmv4W67qJbVC47be+9MJGtjToYG7Epe
c4e6Jc1Fl+DiISYXH/O1P/OndMuuaAq841VgaHxAB6ab1NM2liYjQoUyukzYClXc
kzzWZy5qhNiyoXd/grK/WG/Aq3hPUKugiOrgX+stirYBkXEBD81OXgd1rvD+i2/k
m3BlrsNqjO2MbUtp86Ie3EArw/vKiYRiOneUCxBaqS1lyMi+kTZEFkzMlMez2ued
Nx1W8u1ZurzJFyv0O+dW7to/gzD4UIHPiNQaWIayOB8j8jSf9C1fzOSIxST5ajtC
Nm0HayhtPXWr1AWCGfre9yraRpJ0sa0xeeIT+MOp+/+LDTAz28raL6sZGEd4qJvB
TPN8uETqYSWdTgrQf1GU26SO++sAoJmyL8wv+I8g7PeDBXKj+OzUHbik7z4JWnvL
gzqaPfpOzwfIbUze2/ch1U6zsdgIK+LUrZXJH8yO/wbEKM6PHcQORZx40LhU+p9V
x+0YbaLso9+/VuIq3X3xWTeZ6fC3/+l4nC7r/DJBHNnzm+llbC449sU8FQgYsXEp
j+RKbr7lS4E6RhqufxvwgtmVjQiFJld7Zg+rzPh2NVAgPfmLW1oQzGjHuwfG7M1X
hlEsTi4FyxLr+GFDLgsyndlecVQKnir8Pc+zf5YIOjFBKVF/YlPGDvX/248jPA/K
QqsMaNER82gkikI/FLUuNnG22ji4OC0cjNzv9spAk7TCxlGkCYQhiYWD8tiNkaBD
Q5n8YThd0VDHDzJ8qSqjS0RvDJDvqKrADuIkncHQmwfKYGkn3Q5QAvtW7ogAUHGx
Xbnywano3kj5Me85l6r1wNLJqRvxEs6pYy8P2deQEsw/UsXEpOUZflC8BfsLr2QO
zileKL2hWFq7EK6KjtlyfjjU7s23THRM9tL/+5La2NZIIm4f1dBaTV33BUNbqBwV
sLiMuMB6EOdQ/wOv6BR0xkGLyR66y+uHj+eLwDjR9/dD6eftV1zo0npQay1G7fUk
NKlxKtKOhHJiAbp8mAqRHTL9O7o+RrkGRep03BbUnfNF2TxmbEAB70dtXVzcHh1N
Xg/Ga94CDwnnNv7Wtab3SwxRKmDW1b0Jth9t57FOJvRMWFFa45LBl/iL+DZzTPIM
WNGhgF/Z8DdrXlujVDXcO5B4kRWYiyoGx0tuqiD/6FuMpDeY+RL0GPXNG06O2aev
0rLP/p1gyxz0omSUx82JH7xdt4nsj8cjJNCAR5n3S5+YJ+onEBcSgKuI5V27hiNB
/5vW8NUPhXVPU08u3kSIdnMO1NnprzDjYgful2E5qsLqfOfglJ21owsowNizHn/N
GCgx+ZyQeIogyXurW/Bv81aNvgNKQzBSbFkeD3ScLAqAS5E+/dJKNMB3EZBiJWp8
k6DYHxBw0Tn/kmBot9LJIO2GqTrv+uUOnpaM+70kYV6NYtwQcEHB2Bj/SHqYN0c1
kVjj5U4iiaxVugpiZJaKrBDAmQYRDYKyh2+46qcNATraZipoQiskD8Y4NIjU/ysM
/zLIQVPqjtUGS1iDaGmF8zpAZBhzwGjErtdSoW0eMFr4BrG6KbdFrsHuOV9W/LIV
sfnPmjYME/rHSkKo4LJuTIfvSL3qKI9imrjxJqnXBfpwkyb0N8noHg4juhIWDkVR
gYZfJDWFIsqkTTTAnxFHN+Xl0HzeOxAUtI8gwUk1CwqvN+XNp2XKYXPdvcoD0HWJ
cTRMzVVbHRhX3Y9+X3Ggjw0zLaLwkb/5x4UUbyvchlJSNNkSg25X1ebrNhQC3zC3
rbA/7KT2BL1LRrXn8FWyHw9iCQCZiV1gh8or0FYpjs+0vLQ6ZmK4cHL9fqU7Z+q2
u3kwUhmKqQqC6tJvRFljRrnvtpwJoIktt6DKa4wwIYC2x0iS/YwWMXHy1Dy5gbZd
eZN9cNoC3an6VQeeQpP4zkK8F3yQwkQs0J6wVVWA0H88uq8oFIcGSP/xoTf2aCTd
ep4ApXaY2Aug0WnXfhP0cgD3RbFjVrStFNR6rpZSsS0GdN+R2/VNE6z+rs14QrZi
u18+kdPppFNRGJAU0m9qFjWk3XYbvEz6cxxF+8cvfWExJ8MY+Uvf2/cIAMof7Q1j
fwb4dgntGsk8ei7QGy0/wD6N8M0QotCCOoWcV0bkm0uGxRo9vcoe4Voe0QA53PG9
smuMjBnEK5iYKB9Z0zEi1ycvAC0p9juYIF3yvyzh6gZz8NU7aPGLHdnnEk3l8qAP
dWthp4rzH4B7WyRaJ98IoAiqY0ZKmSqJZbj4ERDfTwOQfMa2fSJTD9YAdJ4IJWAp
zLHxjSxFq4OAyg3UR/kjXUoV+T7PM6QMDi49tGl7lGcQ6B2vZf3YTnVO97lgYhRD
KTLNDzCiNrzpGzQUNE6sHWBMQ0zGEIxx7+v/nKQEkZnpkJTESjXy/UWZoXFEBEuW
dX5wgebnsJp/8VwbUimERN1ur4wzU0E4+fGD543664u3l4hY/52nZCX6hIehT+u/
ElpQvGflGTrGb0cpDPloBUr5uC3ABOLGwkTNb8unNM6ZAgXRM5oXnUHhHnCIHmNc
yJANLefFuZBqW+cIjrsnf0X++oT5zxa3lTvcUwPOYzw1y9hgIAn//w+8xRw9Jgvw
/3BlErkvJxH//zBYREvuZbvjARNwocJutj+wakb4uBN4hkY6Aem1L11PDxTgjsA1
L/T+YsAycP0raWcy7mr447VgzlKMh5xxaYJVU5boLeXNrPSLbKCs+yILmTNn3gqe
Yu7gNX3qDFYyGupRA+Na2k86jHSLDMPgUNipwK+LoM9Nh5CKXLxp9ksUEpe7JntV
d8oulj2kZRLPtKkoaYoclHnt+L0xUUCwCuoEOyYbsx+k2REsmZ5eUhgbCt3/am7F
bFduxglo8Ilo4RcF8u2gt4Jc/d9AokhIuN+9rl+StN/olRrVpOZgor85eX+djnXx
Ed4yWdB2FNSV0k9BTxetAAamsZV3OUPd1I1gIC/hnht+b/PIRtX5JMpav14smHgk
Wy2csCHrTHyPF2lCGJfNyN+bq53sGrBw35Ctwyu7TqQqyws0YsQdDYRrdXN5vI1c
40kpfq8KahHMPIGTDIq8JP041TiPN6JEB6an2WqJmw9IM5Vy9Hcrut9aq2m5lzwE
04MGMDpqoZvJqT8d3jOVh8YyFT5lZoo/q72+Jcfjh0eYUYDNFbWqNmMJ+SqarZuZ
64LSiZ6t/0i5HQVJ6E0/dms3nAH7TVzZKOvImTI2eWjwAXIJsWPFolcNNQ18LifH
jzBg7UhI+lwCLvqEJdyeQnG8Xjxt9rEcqk4LTFpUXNLl3IgaSeEopWhyb0XFHZwT
1wT2OrKdy2RDuTc8cCGEpzqnma4TraTTVEb7U1uPmBUu3c2oTe2Iqg7+GAvtnk5L
+/28/lIIQ9yLxkDtxeD9eXIBJd8HKeWpsQkv6IG45CW9SHrhljGT5BI/ROxHuNpI
oBCvEcRcdK6R9AAhvkjPENZV5n2XbpvsW5cE3W6eK2JCaBhG2jaQIxmINFhN3ie3
5bPahrvlv+3KFDoVVzRxqvliuHkbCG9hKyo1hTB2o9YWiIeFgJvx/m4+GPslRjaF
Zq0D1IrmbatPx7eKo+5W2mZwPsTWpOjd4SfCBiO9W5pJCzAhzQUs9q+3I2KUMFLS
Cy+KsrWMAmK+zN0zPyKpvMhx3/cKskRBFmEfqz6BtIRR/Mky9IB4wGTQyTeHTPLr
UwieaKJihhlLFF14gIqpMybcyXTcyGcY+HqOXY4BlUC8+lxcBcX1HOCS+g7iKBTj
V2QNRboR1zsFrgC2nOjSk8LN+vw6NPwxJunjMjLFj1199E46io2usScem8Hhfqmk
+yTQsBwPeVpIPPpFQNSNw3Dpa9gffTkBbD/7rJ/VaPs5FcPO+3iKxHPVLIl1S9gl
wNNZTlx8am+QRbHaOoIdp0DjTA30Na1/t3IJyYlH27AGk5jKj/4j15YniPrlvKTo
Yof+4hGjDNqeEq3cKmqyaiDTHye8iGj1PfKXESL6RImIcw0tuTpEHZShArJyrotF
/fDe65l3zB1ItLEqJtsJZBuPR/rX83Hga/q0GIgPIddbobO7uzz2bh+cnwkGFKQU
VnQcfns9DIl9rijFKFkt93mCDke/mLkKofG2sQ2QiuwvHSvRZvSa+T6vLgPaRDOB
DarfY/fMOZGayw7fLjeq+2Kr0TRY3SqO+bxKiqHHIijK1juLLHxoTXNVN9eyNchj
DOmSIII9ALiO2YUL+qZ6+PEAakRplwniLdBCzrR+QCImmLqXiFXL6g2kDM59+9L0
KnrjZcTxuCXEmNPIRT/Llz//uWDbT1dr/Xtl5Zz/7tCx1vJdc0UrrigWFv2Kw88R
O1pb1bNMdNuffF02jOltQ8CPkAAg6M7HkmBXumPkTNNHxU3hhWOyBRbWxT4M8XYf
kAopcKzJm4mQB/WtMoEET2VuCzw9nuNXPcjCWvfxcjYo0A7KUrNWUOehfwiotV+t
5xPv/515jcWk+1Fqn+CRowtuze8QMdJmZJXVQ8zFZOVF1r3jz+eBOkfxGcgx4gAM
Tp3qJCQ5tUrXdoiBL4jtwNSo2/Vh69G54GahA1A3mCaK3RuzCm8d35ZVAcWi//QR
+Da/7xjME7rcN/vEHLnf/ohOKnNEcSBXi+3C1fHiKXt6bzDRmcJJtEiHEwUnDwDe
Uno6IVX0bwQE/VQm6Syd1bFKRt/OkwkdiP44bpxIpGxLoQJo0Eas+AKqUAdvYiJm
QKdeMbIJob1NjMvtMa5dDYQoO1Bc+OYcLZeLAdm6p+tI/8+TIboJ4QUGZmz3CNkq
4ViIGBSo+0/yomRAHtr3IliCw/6PW34JYSHDM9RIbNrTAv55PYnebRwYaJVXymFf
pqJ6hQtv+scGaN1K9IxwHOtiwq4lYQ5p1pZ7YPz82GPTpUxuQSthBnQkJkOq6Gec
G82aaQ1GPNsULRi06cBo2UId3FZYyUvBUZpzhYVp2IqZWk97Q5Y5vf6sJuAFO2Aj
Mas4+C5KOBWrAXYXaGFXq3U2ijUjWcg6t9pZRZBqMOMj80G4lWBJsl71bK3U44bh
+jQ+Un07xvJxoI1aszQ7dw2MKrWW9LJpUtI2UEe32VZ+izgd6ekWlubeKcXpmkNq
vn5Jd1BlrK92ky1oVxW2Cx7vIDCuC0xbduHZxP2vuxi/L8dFGooOThmFDOOxtO6j
UJb5jW8RVrUJRF3lolyBK8mA2idSE4wapK1GETP8DGenpEZj+6eAMucCtRj+5dCr
sxvy+QgEmR6Lh7msYpXYewhXIzJ5rQM/BG7OisQZSdMXwaCzS4JnmKJzYspxOACx
rFUvO3hKatHzfK2VF482CVirXyNJudsi6XZYfo/w2rPB/FITg26C0paDbgclm2li
mjY2AZUwLmcvO3er06lwo78D8xg6WhdSMobqoWGYwEAJl81pjq+S0HNhx4NhasA2
E0XIIRpH3Wh+V7yET/P3zl4o4ex8dU3i/oNbuE8mFg1OTnMI8ueqMECmxx6dUoOI
8k26VmJiBnqtz1GFRC/eZOZRBAWPPT2+MdR/Bag9uOMJ1I+kEScJFwMrMpfb2+sg
YToO2/KHDaoQVrjiCWjGNyuX/NzoHqQjk9YZFVUKEQiIPY8Q68HGewOPUzmkCb9i

`pragma protect end_protected
