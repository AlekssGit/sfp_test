// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
kJOppMNhY3TbMPQ8/v9dXsabmNRlqQlKKfqG/HIXU8MGW3Cnrg7iLoof+QoZFZuq+mQlDSWplpBI
bww56FeTqrnMagDFLfRShass80e/RGsg0GDsslMZnFVplcNYnOayzWSK1PGsBd2WJo3kaR4VPMNv
QtVu1eNOnzjKghWJA6lsBFP12eRr7AN4UJsJTlu3zuG84lxxUCyiJGtWESqjuo3P3/mXJm1SNbfR
0ylItwe+YblR97giNxtI3EUEDxhDMfTVkK0ZjgRzQSj0dLqjzguaQsY6ISZ1Iz485mekkQExY2dj
0AFdBnghGJj4N8dpZOP89YOgona2W8GBifQ0bg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10672)
cUvlmsytcWU1CI6T1LgrArprvk7FZisNih/Zl5EpUhUTaMYiGqQSrKaPrCm9dT+aj0387lSEYPhD
QWdKLwaiuKllzHtu94RW7oIZEjXhyc0bAU3GoNrvq0MS5XEql4cPAYhNZSSHV0kuU4BG5tgZ01lm
Ff3VpgyJ1cuCpEiRuqHeX/jUpyqwENKGDO8PVO6BmQU7zLDfZ1gfLTzZoIDO4u9Cfy14JOdtKJrr
dVtEGDNNcmynw9VXgAZRkx1Kj6IeGAzG86fHyKtJ+xn8QFW20XSNqyZr0n9jnpdPYdsmqNENQPsU
PBnD/hQRSircHmuy5MHKfPF/SIhg2G6BmXN5YsQzsRjzHNJ8jUu/NSf5KvZvYAMdQGQeFyEnAkTe
Sj3hvVx8DEXJXaqwsEM+SS4D1QR9rVkLurE52YgB2goGhMVrAXfgWYU+OuMIphKZsKu6URRRvhju
uSVtZXJVvRy2+8E3BnOxCzoj5OjNmH45Ex5CxfiWoYTNCa1KUTyYdL7zYAD4EiWuwX9MmRxm2klH
F46OUXvEcCJ7579M7JsYMecwYeG5dDRIsdib745hT7J37WeKigz6CZB21GWc42DAWWBvBAU/g/om
7Tz6J0QpT1Dala/I4O2Js1z/J09m5C9DYA8HBE3JFjwDk72j17vZOVcQOqzC+VxHSRk+iY6IXtgV
eUawUoy6UfcF6DUyZ78NPZHpVohY+mIfpR7WuR0NcHt5gQEMlIYKgtCERGOA2ZzNMCoidvNeDZ8W
5ZGQ/hKtDSV4SQeGGQef36hY+u2RSxwYoVmAh1cHt5LjQ6O20SSSf0H9uyLeBgbpuziY4VWvreIU
wuhdJYaNQhfsV1U7B6JU2cE2Z9bboKK/pFdM8eVfblfwUSJmPEt+3Z9hjPJ8cfA07dbfPDbBBSsr
4PhJBjNzbcC/0cvzT5I9NgZUv86mKD5V51pGDFfqwVNDZQ/zSm+H0trZIyjCdz5oOH8H3L0iyqpJ
gT6ICUejhkLLz5jvTwjyJldHVPYz1Bkm/fvipTual381olquP5Dr7TWmWbgBylxjvdV0bLv57dRD
d3LZPfjw6gTHMG34N/w9/SJqIEoqDM9RtnEhTBOvn1pGieqZoKO5DJ4HjuAWX9i6VT9Vh5qodrCA
P30VUgsYxHTXmTMBqErz/eSNlI2VWUBerZirGFFfZ1VbZGC7Pl+f/ahZMkAWcxTUm1xJ44u5vsf4
6Z9vCmcn0NBwzVqcjx0NS44sAZBAj0AIBeKzoovYg4HEfjz3NyIlpbAhgGaELI01Dh2IHMuCyjlZ
tl7XB8TFw/6BINtLHFWUHj0iNbO2FFk7LV2AK4SgUwBHpNdaHWotr49MiP1jzka6e90dd0+h9s8U
Lmu9qQyTp0WQU7TRW2bv4OIRprCyfIKH+eMDvTPNhUzzrjhFGwAxqD7AvJQYvp0ZlQFXZkzfYLZH
4uIRbq0E2rpNCBUWbKmlnyAducQV6vG3nq3f7qgTT1n3qMYJFod3OvLxDnAix7N1EAIP/ImcaEtV
ubgn0O5v7z0pfTkSeVdsXdSps76X5Xo/utqRwloNYss29QzcA8KQfyYG41sgMU8uvS8DLIhrlcXq
B1doy/EkHl/NmxaDZKZvvOSSNgE+xd1gPyEAqwhce9EERZTZv3RNjkd256VAjg/Wlf2y9OqT3zqW
c9QECrl5IzILtaXsGvdBsrCoJpr2DyBNz11apBBt6eiuUKZCYAqxJpoX5ZdfJnU1EdeIL6iQ+PQf
wbIeuMk7hjdTb08LhcRK/MUVzxN5OnmpH0tCbpNLE/Ca734nnvCC8tlY6WAf56guMyFVNCQvyOUF
JOZJwXynHV+MFesBNelWWoAvUw3ujjSn89uZZ1N0bDtq3+1NhVs2wBbcebzikY7CTuMh5O9rSG68
rpk/1jsFm0R8GMP/qX0oa+TkVq4Swh1BxQ2VBgVfMWAI56lTd3CxmTHdekuF7b8Tv2DQ1lUFRB+c
Vh+cE4+O50o1Vyx7M/2palhA+yORxyv2FSEhO5137nu63mzsq2vFk/LWQO4G9p9t+Zrw5XDDePeB
zl8iamOaV7rWi+tuihK+xfyLftZyDGzz2IEeq6NElB/Ai+iQDxPubpH3kGdISvkjRpEsGGk5OddJ
zcsjUitzYZVVc9HH8OR1L0XKklvThGZCXyuxFjnzSW+czLKyy0+5SjpBFKKXeesoDatikSUxIhCS
U4fKtzDctJcKJrwtdhpeubyxfYfLApby0CHsGaawlicq0bC58ZGf+EoyBBPtYlobd+r0dAR47JP/
iZvZazGVwfmrsuVzjSwpzXG1Xc+j9QbZ0kqckzi8AT5TPq9NLGDcQRbJGsXJ1GfshXkjb1EPlp2H
Ff4gupkbQzoEeZNwQ9siVbnGyrmbmYrZDZdQJdrC8Pr1ESoWu5c3FEr1nDfsdHBhPyzcu0unQJn+
59A7Q3TlbkB+3XL3OoJqFfiT0uY9NwXwi43Q4yGAJg7O+BeE6lJ9TRGu8fU91Y545MgLEWaJZjDT
/iXLlXtnTIIwTZYuuZHcb/FpbG43/ScoDetekpyXa7aSzS63GnOz0bdunssFsZJCaBeGyq8HY81L
PC2MhEbo6EuoF2PrJgWdWTjHoclCiipyHvQVf4cslQe3OXDd73RONYbEh2FmdXirvJRvLtnCyxCj
m3po99g35MQvSoNmkMRwAQ4tPU5TLDRCQG2PizZ5rMyZ7Vw6kS7RCLJX6RAmx5XU821Df7mwWHT1
lMphjfl7OMPcR4AoLbT7Jl+alnRYyl+XyNbnE1y9i/0mU7qi0V1amakGlkFebZDxE8zgNZF58HD2
MpvKhgBicW6VFnZ/yr8k56crYPKLVng+S0GmieH5Ru9E40YLZAyoa1jUQsI6fSmJk5H1HNylI0ly
0RsJ+KW4QgMc+fYhuKd5iBs/uQa2XqajVxw//nwaTnVcvvcKqLbM8PKEJ+RZG6m0CPjb0RINDwbM
yK1ndVjPHE2niPbZ24JwpBu0WSLKRbZw2u1IQfwKVDavwIV3GTURm4wYltm7zJGVJhyzEK/UnRx9
0NExmGKN80kJT1A0t/U8flOUPuWVGqz5rPSC9MUg0PXQvdzbEIAxV96FUaWdsnJANztfHCdlH5SS
NG9xoBRsDHZWCQ79x5MPSyJLr3zUKQouZ3C8Ajlztsro9LyqONzrOsY44YAQ0CpH35Bkwos2X8rL
zTPBzsVIyH6W6ekOxKvnqROGm7EqCeIS10b6Rl/4LhZvpmfiepgv7LsDtFiw8wyk72+Ro/T2lYFr
rQf1qZmG5D4IqFUHIIxX5aWiVnnU1v2rjbvDNl0oe6jPyfP1VYvx8+/Bm8W0EiTb/jwKkweeerBa
fqxa5VTIxYqTZlWewL3ByXIXaHeJZvpEqgo5xEcRSZGTnq7iy0PUlJjB20Pi7pNIThuWPaPmm8uX
rUn87jUmiPz/7xpvYASWF2473A3E1Os/5UzUjCYh0GkIVB7ck3lZLpKXmPSj/iTyUwCm+HjyDCVi
tNDFk2X3Odbfv4Is5ds5+RTOjTUN9zJn4VR6sU0mMm3xw+Pz3h5nS+yF1iaDGSA9whKbfU54g4pa
CsMIcEXZsCxU3rX8L5xwbYL3cOHmym9ysBiRd5rj6/Jqenl8C4ryo+dN7FoXa1FP8s9Muf75alQa
CTshCmO7k80wvW61z4dW17AfkpFJmTE7c2t+HzANSWLUQN8PqELd1W7NZbQlDtYIodx7tIzxefu5
edHK0ESsv5Of7pAWs0ZWkRhMOxB0nGzoeBhPqZvvl6X7+WxMx7Ct09kRldMilSk6hjrt4V3VuGOt
L0zmibPeg/zXJt+kH4RQnVF4dwkjSTOQb2ZHI6vdV6uzoulBcS/u5K2GglQoEOa8MpNIME5Irf7O
2irwBzQ8iEOLXJ9Mi3mwiwBm/0Q/gv6iie8H1yPE0qxpig3KEfbpDSU2C8zRTd0YXVjxeoApUVP8
MSy8euVAmIa2vu3RoUvf3vLvIqBLBsbuz8257X6xCma0wfM9+dGE8wAexAi9X9V3R3yne9efoohz
QiSmqT548h5hkbj3FpIWoX1Dl13XJerT6ItAqP8mv1Hei+ebNkDnyCphCypwIv8Jv4ba0Y9Hsjb3
XcbcxXPUolyNNEnxNHRaKrjFX0VEdTzThsCQX08r7I0kcZ3nLG6DdMpFyInZ2ZX+p8KTTBWTrpAc
U/n2FiQLjar9FBfl99jph+BjD6r5rnBGt+no2yPZfbqhGth/qQpTN0QWpy0MG4AcdF51tXAw7iyM
b/7x0EH2Q0CVhv5NwQGYaAVcOoTr2ikntc5YdC6zabJMICmjqK59JkzcmjpnVOZy0bT3WSbNkSed
RmlcPB4giQBTZZXQK7XfltY3KrTK593LlXLo3DNzqVg/tvnR0XsJMXpFf2yCMSYwwjRmthXyH9Up
XV9yq3ipuEDTICr5IaYe1778OF5AA+owfb1xZogXdCpMsMT64ZrwkXXqjn2AtqLBj1PQdibXKSN5
UL0zFRbP6AbGeFZzOZNvGxgBF6Bc7vNC9JEu5MTRmAauoRUpCxMyFuZmH2cPvjwujKwGorZoNKbt
fuNtwA12myv/67DDqyuzYQFYHOT9Zv5Ob+NBWSimjaO1oatsKoos3YKj272rolcj2oBMQEUGlaUo
B2SmUgbrSkkLsT58YLlxIv1jQ5DaPW5lvU09IKOKHgz7sddgbkt6ILLX3atCRgLBpJUeY4T9JGnP
BAH1cqg/PC7qJ9MaSB6t13m7iuS7cn+M5hAd9qZ1poPG7xBArRuoxoYTPC9kMr/pAy0cbOipJIKO
N/l679QNLjhrL9VnqP8LSDpP7sjzVewWq7jrKhRH6PofTFD4N6o6t7PKUPrOTa9vaDATSYI5W/8k
3WsWBtV9t/aBQxehrW/tGKYvbrnyGZIx/c8PhiujJ+qIa7CKAg3K0/fGfiOL80unOL43yU+8BpQU
Y7oxUHQTmzQDTIxxSOuroYQkxF0LwZe9tdr9CAMYNak9sjwLAnzepFHxMlDkUpCG6d4ekRNkWkYk
Y6Q6HpeeoYlTS0LN/C2u1DggXmpmNmOlRWFYnyVTn86Jv+EzwZFdyI+glKgUYsmDUTqKtjmxPpfL
lqHBaOwwtyvQlujGDj9/usXDs8wAU2gVGzK0ONcK1t4AfYl2wBMZSPKDqWIxfQo0/8oKJnon1btd
X4eN3ZqeuLgW81tFAvfX1U2aYZC0M62vsq3iu2vAi3SBwtE8FINlV3wJm3+lYM+Tw5GQPQ+5fPoz
QRGb5+DnG9zChQJzFL881yUSa8qzGTiAS2yf5NNB/MVpxKmqyNPwaXPK2LK/r3TZMA5vR4wo/Z9M
2QO5cAmHXX6/NuYi3U4q2d6dFs7ikNFc+R8bVGpYrFM+262XjHeVZnqp4+p37XQaPzI9aMi9OOu6
Tn5E3KDZOgS3k4eaYt5CsBpnfbEhub/p5BP5hWvlkqrt4Utl/umi/z7Cm+w/OKEDHQO51Glrrz2t
1aGjvVJ1d5dcPCIsZpEvWQVwnwRZyIlD2O8YHVXJVqbP2fdz0/p78LQnOfF+Ls3ujyCuMJeucVML
l2aOVIbRbmAl9Q8fLlP/ybocZLY5wRdPl4cxaloETtOebnbXCnGoHbY9KFHXxvF8sG3PlQFKrXV2
vTY8Oi3jSk31WtSTvW1ALYg0BFubRA6ItJTtrJcznvX+4ZXoMXMAhl10WUkO6XUCT2f65wMvjbk3
W8awM20SyffeQghellFTLTgdMWDBE67ikRR3AmmTc1wRJnULIwxA5n9qeAN/yh2fUeWCwIO9BK6R
TYfFkENiDqo9rdRnzBlyQKcgXttplGLVAN7Xuu0SUCWc2JLO5TwEnA/L9F4cIe23vGHml/UiMvc8
vMrBkgIJ3OQ+s8iutV+0Ge4zM53S3LrH3xSqnv9dYJM3V2FJD5vYTggfGjR+yp66pxnd+G8zXtxL
08/l3BlpeNG3ddJbpW2iZoJOP24pqwe92egUatMpArOftYLzmhBfsy+EdrvfhQeR4XqlHZnNjuti
ph6qParOyK59iY+/itBiDB7BvPbcPTfjRkpvkZmYE0dgzWbIuP3QE2a2lw7OXzO4BzImypRG3BBq
E8IuKAkQX9yB2VTML4JzYtr9MFBJiQmWF5anMYDBl70wn6+ez5hWWxm3OKby6JyHMyqNluG7rV8j
E7a/vYGMz3K5ShGlqrCLDUQfzeu4HtPIgcrMAiI2cRdNq1pm//XfSTDFxANVmZXknMO+it9I8HCA
ugm7/PEPhwFORQ2EVWO71o2NJQs45x0XxOiM1hxIZwlOmmKELuk+S4zSU0ah17ZSmnjiFJtErlyX
TVrJgb40p0Sxp5TY02ogzIZwSSZ0toOU+/clSTTjr4ImRnJCq4Ev5gD8HrFDuxW57Yqsmejd8NNz
GxpZxZYAVtzan26hzBuWcC36dXGPPpy5fovEVYiCNu1EzHhPSCJhi77RcJEPDHz///e4RgYYKB6e
eNmzHE90AvPPt1Lkv7RPXgs7v+4xaBV6EL5sWUTNICq71bF6SQVCaBTrGpNyBTuS9i2SsQoyYBTb
pEkmv4Z5meJ3Dz85i2dwYaqlZ/62Ofq1SSiNdWLA3v5FBNXEr+G6Tx8uzRP7R1UrYAo60NpwE7IV
nvinaMCFI328D4yq3K/+a2gQO4BdcGZ6JH4QReN3GaksX5s7wEwqoKwCc29OSciYw1OVHOxHL3Bu
WHXF2yMmMf9SBSkB3b7/0qiJGlL6DZnNhnh3t40h+trTW+uqPmo52wutjJaDCvWshVw+FWWHrGlD
HxySdlEie2VAR6/2H+ZrB3CgHCJ2H+vbdD7LHxLZiS5+bGcTy+R4T2wXZDTgkhGlm1dWJ21FwFnc
Kg7QygcPlOmWgt9Qsuwd9M6wpU/m3oMdj0m+KaPnqK9uDMAlTpfbgNF1o1aVT1mvQ3Pj9ubKPGHy
wM+XA0JrN/0TR8LmvyQi7QJrLdha51XFz0wd2gti7Vp7IyaryYSsDjvvYM2I37Hf3d84RpLOElMI
Dc1v2f3FwvqeEBSsJUzwPDubaa3PTn6QTl1JPYkj4rNuRu76z+xPbHeeyx7B0pCDdE9VPBZbR7vY
sfWC8UBJyzjlkZYUUpA/FNDOvsTcmjU5hiLZ+bZkwRPdy/JYlPJLN7A5YWPXWcKC9eGXhSFI3qgf
LIpMQnlWUmdQCQbc78fBnJ0h7j4cmdCip/KV+QeZA3njv8PH6V7jtppQ9igv5Md6lu3EGUEQflvb
r7bG79FiiQjas7vtsVLGpNjl9D1apBqdxUL2j6Kb/XudE+yAhA/W71+sFUTnfwnvLWNjqvCLXZum
SqOcaSPG2g2/HmsTkzZ8Ls54GNQFe1VokY0tu8juEw2NN0YHheD7dscwnMm/cK2BF60dAO6pmfKC
KH5CSPHL1qCQ3NB2JNvGE9X7z+dpAKsTzGxDTlZ5JmmZ9cjzgzxFFV2VCbgSXyfbvWzD3rhtSJlA
yFbQXhCp8bL6HW/B6SODCXD3wuQBueuV8113VqpeoVPF+GRI6d/MjrDbFy6ujri2EzgOjDFpUzJd
oBoRn1YVemjVqq2gWjtFT/s9idhmRQpOXmNNEqqcCUfHVfHIYUzN//Wx3V40ZG4Q9g+IUl2UpinH
uFLDtNqIhW5Us8zBOTUgKzqHV4tfnlFl0Mv2FNmVnDiNU0Wuqhhsl0V5D2DbXTx9ZaTFMF9I+drl
nXoN0STU71a+rCak0+IsED5VTVb5rhjnoqVqmmSpLt5/tEMs1dValj6R/ZJoJSjQmWlV4M/5oZNz
M1nOjNwHO6btiq92gB9nVwI+b4T0m/5YvHjhzKldJkr8isGhmehO0BQOfqS0KECFnjHXn6wGKf4F
RtLDyO5vP5idlnn7Cs4MciFGz4JPEHDuM/JDAhOrJ75GlEm7GuCq3bZrWY26M3DwBp3V34f4paYd
7/qhcooxxifHjrmeXFTqDSZRMrSYKzde5E0Gdl4EGaYvki4v3Rw++JRI51F5rw7F3kAXHjaS2xv3
MbpukEOCJ+bhip2HIcqbcEvocz1OCqjbVUOTPUPTFUxiPhorZq3VycobGV7bMTLFZCtVxs8m/umb
J3Alh9fWbIgijHwpVMbDuYHPCL5P+V//+i+oaE1pcz4Ib8V3rC71Y9GtXFmkiQKOyKj7/iRGoO0x
tDgIfUD68j3ePbO/1yEMn70szC+qLvKNeGh3dzXAAfN+OFV2IvbKLQz4LzSDpRdpzCO+NNFyrUdl
bbiLCVKl9TytYDMAIsSF29iQFd8+k3zmE4qlFWTz/frE2s7Ft5EqEY91OfntBHr0EUfo1DfYiCAz
k6dB+t+3kouZhd4oZmt7ZigtXsOJvo3MxCWbqb91NIFWo+BLB8CvXFvTlT/IdL5u/rI10LIgFbH6
3LsPcc2v5vxb9u8Y0M6lRalfrR5QVPwIqB3FP2LOzn7bZ3FgSTUiqTTaAd1z7FZz4JPuBU2yYrtr
52zcrhBkGPHCSBRQovkhRXnTJ15WHrQ2COomeoAk2w2sbzhLoVfgz4F/RhAuJmVVbD84HbcoMmFA
/KTwQ1RQZGd7ZvEX9Rmj6qEydo75cnYacD8RmsnSHZKgSlz3GDiVigjMThozLid7Q6GhC7INYrPR
mKOmvCnghu8+2yrhH5T0BFuRfm3Y7srcVFs+ZcCNhYq3Xf8aQ4tSTPyI1cFZApgYcK3mGKKfSw7I
HXnI9q36huDBBwFjs5IMdrjfmL/GQMdBDXoJxntvkYJsJKRI4UoavmxI/OMGefpTAy1QWwO0VqMc
rHgoyC+/0BGmsNJq8e9cnNbYMf8z6uhfN9Ta2qjZhQRqeBJqNoIBSAV6QvPtLJ/BvapzqyY7SCHA
QxyddZs2lfnXCHGSVCeuWCYx5Msn8emZ7Cz3a155ZBk8FMPkSKA0DFI2Tee6cs8k5albofuFwGKH
TfhMxSlq2nI/bntIeS9AW0HB04WFYFuuff1qwj0CXBVpxpws2uvpcoBIQajmsZtoiXoTamyd64Fk
fSMLSlFUuKkqcY+qJGqOyvCc9Smi/cRHFLt9ZpZ1edxtbMKTFLtU93IWQBK3ij3Pnf9ImbCZquMA
oq2AQkIw5qthaQmc9/pVoh8v6UFV+xwJ6S5PDY3HX/SAVj81c2y63Hjy5ebzdieiOd+Vzc0EKA1Z
UxJdZldCZNGarm8Zpg0BA5j90LSRLtMhMZv1PDbq6znpGvoXaGr312pPQzXjorPy9cSF3fcz88A5
NRRacYD/NR42A2aLJ6fIhS+l9w/zMDaxHMmGtdwPf5J1GrVwnzn6DfOQiO1sz4EAYPjeUEmgvvSD
LhuoAFg1SiJHqB1M6ygtuZ57ColMe3rMRVPCJ1u5aa7b2n7lohJVzGEEht9imSPXIcyCHmAFe2yM
WLrgPen+0qnHDPOFmi36bZ+IyeONaIvGSPdr3dVGx2AKT0HZNHtig1MBI+DZQpb3eVtn8th37SHy
CRTyZhhm5WcIEvgpp4EAEiD30Ia2EqPkLSG6dET5Miuyi6FRGfj1L4ul5PZwZxCK9LNqjAt9vfRR
MoNW5J461ScEBkKqvHNiRAIMgv4D6m/Y34u8RtGI1TZKlnKWWC2VHpIEi42MPBP5WabHi8TIc10D
8yTaW5iX6jEJ8ojsUYDrRmqxU0QHXN/fZ1BynkTvbamOVxk6U9Q2qViI2Vtsv9qA6KWz9zxUtobq
lRgFrO34Xd3RwTAfrNLimSsrT32SOVfrcBl5vGkWXhUz3lxrj2bVX+saIjYZImBp0pETxPi/ibFX
UETErbIkUlujKkHe/DUF30SJPdMoiKnoibcGR5TGGqDwGvD6eIaYRX1c6ek1Dx4+ypFq81CbE3aN
XDLsySZORdvzEBLKCJSJkZ5kPzpEBYlZB8sbLXu+ZYMVn0AqOZ+AA+vgqM8GtEv29O29Q1ltoiKf
FIgE7Uaz0LhftnKOFBLvvN3b/ZGcjiSKCQSlNGlGMZ9xLji13xq960E80pCKwxyU7MIvkQzw79HV
cNalCwkz641yRJ+FGaBrXvBjXpL/4FcITAcm0FBhIDC83LM2wPg1LmsJObmwDNooSqWP9Y8tTlcs
EXOLU8ojs/bK3xTdmWnQKXMgXoFsHiThCROIwvwcL6Hju4N8HbPm+h7PL2HSekbG+DdryLF77da2
Pk8/enmUp44XS1MtFPgGkrBAYt2gN36VDI/tfeinllbfPbSWubu+zcEdBG45QX9OLn2pi/pVvPmb
NabPFyyzos5TZ6PV9u/JkD4NcNtA/2Q5f5nMySXKeFfwf994AkN+oIyFBvbxdw3ThrlQyF9zTkjn
nzDSXQMkTQ4XPWqLxN3ck/VxWQuo7fnSAx10gEIZGiY4L4rg+HtTAfiuBfUJjrx/Hq0mwgT/yQ4D
9m5eG3cp6oIY9IYxN5+ENLp1T8ZHJMQscFdJdNpOlP/DWu6WwBUm8h02y2A8X0KVsy51m0LLdR4F
QJmWNzqhiN1LXoN3mpVpGwy+4UPHL8+lADUMS9FPBqpL2yYjWFHbiarUDcbLJGcKH5xikXWc90+G
WkKolxFxA1MSYmFWSSB0q3m8EKLg3T2rEnK06LzzgO5E7EbX5wOmQmPUT1YQiOhBFsmrMisjhiGS
z49z2TLwBanrymxYw+6yRihUI71inp6PjNvOWPDKcGlU3WTaGwm8qz3buVABccOGaFc9L3L8eiv1
9I5yTuIUdv1h9cRwQZegAagVuFciRKPxWSQYSy4mpPxQ3jaSmsBtShcNSft4sVeSe5nqjBZDRDfu
mGRE+wqC5ZJdDQmo4wLHFWKxtyOdafslv8L1gylHDDTTmzl1EwzqtAtKjxzWyXdUvRYhiE99dpWV
8IUNZ1w1kwvbTNHc2o/ko/aVen6ehpTaEVpS2wAZH3aLyEe+LaUxC/8JhMo1p64o7IJCtsOrZQx4
LC02sDV9ZONxdu5kJETgGttWYAhO8s5MjDv1o2xPvF8JQJIOObDs7NHAdTmPMNFYc0HDnA/LLdFw
0h9IYqwxVGACdqyDFe3pFAJzexoMLNVfDUkPe89a2RGPlBCDJjsh79Y2DGWrD5Gpr8lF6wLJOn1D
twGSyR6+2F4aPDXbnCuXhuJagDvrThf5+oZv7NpTVJmG5ibuw5qe+AkOZRbtC6e9CQMiy4Jnu29+
PXqUzTVsegWtLZ7AMpJpShwqqueRdzd2EoMj+BTfEGULnxJg1ACVWdkvMonqsOYxj6b+A/Gi9Nk8
DHWXiMsJUrnSrOY3LZ/rwCHNKXPiL09YNasbNn4emaF58eZurJWbae7wyJZs6Ib42xOn4fTqAUqs
ikV+7KcDBaykxZUxaJTzBNJKL0/vf4GGiAXIdQxppg7bohChxprhUuoSkg7GsyuLXmUMK6TjdWKH
TR2dXoA4T6XH7PPsbdQRxrOQReHWOuOFsJiSP7yZ/BKbCFAJxRrG10mJ8sUwWZpuPU1r2x33Yd5C
EkyE/TFnED6pDcz7POz+U6txbM6y1GWQwmbmVdGZ0njspQtOwyd1IqeCpNjJ5jGD6Jj+miYqumPg
bODe54yKIsn0MegfQKfLzQ57i90Ge5bl/cplwhRWVVVdFCECcX79vWeWi8fNWAvfgqi/CEWetyZv
BgTxv8o+RWdcU2gNQLFTEA/8Lc8r7DZUDgohmk+KDZcLffEvo4kgMN5CH8OFwNy/lLPSgJkQHuy0
FEcjuTVt3T8a7N45bFOTGqtRCh81FSa3O2UExkvF3o1o/Iv8qlM1J0SzJULkLATAeT44H3jmIUAz
ziwk6ewYw9VwefsmB5Q1XkiEolO4+HcIeL/vplzRz8o96mU2e5ZfMm3ZYx10PLc02YR/ajHkC7it
/uZhLsB0uK7dyBu3GY6rhqP9etyiO3DKtECKCT5K7ZwN4UzGer1paxpTVd6W6wLEGBX/gOpxamvz
br4Dt7S3+MxqEsWTlFgKReUTnzUGxRgasJOD6Q7QH9CZD9scVpVO4OQGxBR1NbmWt4ybJS4XcnbT
nynbGsQt4GTmd+VtNoJuCjW+f7SoiE6YUtgyzXq69MxbbAdHwBhEAthszzW8hWYm5O9TPfePjGNc
K8p0uQUW4ab/yVOCT4a8jkC6zLW/8c3LXmkZVCGLFLu0svq3KQLc8sZaeuRVv92cZ/U72yqDkfKB
sLb+a3sJMXrIw+q8Rp2wSvmbjg0s5RRHoKvL/N8M/vkzLnoYAkGKZnVJ5Jye/gXA2J/gjpfxy996
KQjQkB/B6mqC4PdSUpsgXGtLDZUieb5YdRQursVDpTyM0xTsvRJcik224TNAHDBib+lmXtZxNcI4
BV+Sw+VSqI1kBnJe1KZ7D76RyQjwGPmRZsMfhsL3+i5ydTJesPtA71ZVbiqysLlD4GG8Xa84CU4Q
vP/Um2lne+lWHfRG340vGswlp9V5OkBxzsDRMsVovN3/CFZmD+q6CJ97q22iZpuwMDjNddQXHO1m
miYUSwJAiJaGZZx34f3+MLef9YT1VC7BgRT/JI5YfigESbEDqv5BCHURuxviBPjjBQxX28grnR+s
A0KgU5xscc63n/S+6GbsEiHlMIEuheDQPpbCGFv1GjaFq6DpBw8Y3G0Q5YPo8gBjtNEAz0bMRH+K
1YZv1Wj1yGuhoxMoyh/lBgji73a+SV5ymQ1W4XyL8FJhkOiKWd8n0O4A387N3D4zlKu8x4NSfNss
p9CrlNO7F1KiGDLDpxxDx/oZGpx6VPeBJkqet+/HhtgSQl09ToCCWIZ+0Sfscm1zDZGjOYmlzarV
GUWVd7xYM6BxqIld4somZHBJCi/2VswZ+dWocclmA1lZtMOxyM7ggc5wsW5l2zdi0q4FDbLyOMVP
sqWTYdsRnhhME/GI+U2Lw0CLFhLJBdNBz/Rb67uWLq5bYkCYE7j+neoWoAPpAR9CLuzRl1bqgyEQ
Mpl4YJ+PIM6+tRqDOitHeRbQXTquk5YxJfivPUSWcwj1SgB41qvYp5FryrzOT4nQfCdbb0wapXBW
wx4T/IWLJ/BK6nbfmjZJKgOPdPAP2/3POOkUL0CBqeMOHmVCCHfHL1xM8n4L9YAykLtjXk80l4FK
yuxwxTX/SUPcfOhNElflOhPkYXE9Z+BraeLQGDHf/Q36ARoCJ91eXU/UVYhW9PoFuPPtJssOX0L5
ZFKzkGEcaIA6BT51uOQ2EvNUApn/tuJdkdFmmmsjLnzO9an2xpZ/m5U9RBnr5fo9jeLO+Xcgr3NC
CBhkgoGN4wml1qSWA8ssc8OuwCx6tqckb/GVy7T53+2xcJe2BjEA79Pohw2yIOoZGbUkd4+ZDNeY
+DnwwkrWT3F2A4pIFOF9touyWbS/ZTsVjcmnvU5UQEoYzwi7nRCsZdtmNZ85PdxINjR2z4snKqiN
PASu4jO6F5mp9+YpxVR9hZAUnF2NGlhbkDrfs37RpB4otNo4tEwep49nycspgIh5w8epzDUkrDUi
rfhfHYp5u7N6S+DXffAYXjqtQI/craIilXo8Jntf7qz7Ta7l3MW6hxsDKDlir9MhFOIN7M8G53l1
d75+2yIKs8p+4GQsXPAKeJ62CY423L+E3LmUEBRGwraa6sp2hl1RUeRvRcXwEMdKzorbu5hU+dQV
qrygnNkPjQkOi4Jam6MtWxR9ad5F61xDvdmpGF104J+xOIxaJO9zR693Q8Oj+3lE4+db+HNsWGkf
BSka9OJ2DGlxVMuS3ilGLydLUudneYuktjppmDVMmPQw5F40rOfK8LYeQiCEhfPgsmTTlefqCNHh
HnrgIIYfP8FPGd/LEbXgpC+yZL1xXUm17NNEd1ZPybcaek/R4K0sfe2DA5udRh3iP3FshHX3Ytnr
iDNto48TJibrVNiLmGbZukGpH9QEDpYs0A5WKXg5ANYIE0DOSb3RREBWXD9tOA+GAWldKFGvSk1E
QpL4veqopqlca2/NhQ86AXRuVym6svTGnF6nVZnD5hn/zPngczxSsW58bVLavpRrrYa/ua70p2Wu
K7N8Dx6lYJHk2+bUoou50Yr7BkJra8NVSHGZhnydSw+/nybBjFSfPOozmcgcCEfQ39nnVz6KfV1q
MZFkrSHDVwUNmC64QLAui8R4o/1aeOyckdK6rEEGhbmmj5/+4XhSZq5Rtx5OMkwg+r9tHgwOtSg/
eTTqtUo9HiTR5w5Kbjc2Cgh0AGmWrjWuN0N5/3koneoowthkcCjPyidgiU37+9yF6+t8yYnq3NM0
ttuwF7nF/IGY87oI2ZI9DKqaUdf7A44DniE3zySQgn9rQQOU/HNLklY233nAWXVIGKTtybuiyzxE
9gJbhpMWtGUxL1pBkQ==
`pragma protect end_protected
