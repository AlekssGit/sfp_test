// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
/weaLbWV3fYQK8RACGCMl9V0tLVt4+nZobXwL/OXU9O1IGb13QyfgfbGiFrW2GSZ
tpB/N2WOP3al0l4zqSzx4pnAQnVBxvsEKsxLvWqy2IRWBH7AMAdR9PAAOgvy3tBE
2t4LYw6cDY/yIQ/hERmn3PwS3fnwJjwrT4SimRx7Csys96sxh7bKCQ==
//pragma protect end_key_block
//pragma protect digest_block
Pd99PJjqPjFeqZpEV8h9oZawnCs=
//pragma protect end_digest_block
//pragma protect data_block
MyoeoSWBIV1iQXX5qsLfsvb+NyZCQnKhOEf0MnPJLXyOZWqP3chkFsyPFH+egES/
/+EKowWZIyULLU3Vx6qESEsW51KpSLfvv6DecrOeTuRxQMxdAbS3fXwUdCe7KJTz
mWIBk5f1OeQjo40X+/fL70KbX5X9vs4s4TlcqO2tecTxUjgVHMq3jxOrrRxllBxR
qc3v2AuJjUwXN7VaV7G45pKH1hebsTLFIaT5curIZl/L6i1s8FdBz3Yxfvr0Qy5p
KoIbxBsFMkSvyrMOqEvGUNSq9DJ+CjkyQTf2q3nRQU9aDjRXX60CoGcvOsiNQKHA
Z+w9YF3xxMKj1H0nvgdnC9SZnG0rKjvVyeE8Zg7vhFhj7u0PHW7oialrO569MhfY
bPh+nNSQyv9hCTDqognGRX+J8P87e5fPY3oKV5wkNrqNogZtRDYrEARIkxqkuWRn
tOEY5DNMvdoXDpDXmQUIRqoUFlyawN4g8n1MkX8YBH+THhpXEPhDl/6Hk/N7ahLq
vMW7DGwVIut9rteMz4oVeqiobCG3H8nKM1OPkZse4ao9+FR2mztyM1n0fXxbKrsW
4YEH/EBl44QOCQZx53j6Iyzp771u/1Tb1uNvpZo88xFQ4rYVqVBvGGVsNs8z8Zdk
53MujUI17T78jIh/iDyVF3Q0ZgSht2+tfmOxfRxnWt+HAoWJtB5Fr8G171s8ahRZ
SWhmxoN/PkdIi3Ump9uKThP/cHUrcsTnu/kPsaMuS8zzL50sx5/vMOzBRS2yqqRx
ImjUv+1YBIsEuFQEVhcAwzSvKEHaRiR55/yms57h/SkvdhMzrLwGdGD3ZcnJee1l
mAVe0lIAgZhxDymlxH05E/SwWbYt8GTfHFosO6JZ+7ZAyxKZK0PicWfWsXL452+G
L4yxn5uySE8BRbSBstJum9B1FEo6B5SyEM4I14hTscEX///V92oEpqQ78Sy2G76E
iPXKVFM83+RinqlX7NhtYf/rUNC/eN4jaXWJrg+2dDVHtP1lA9Ts5VtYOwuq8bRZ
LaZ0DeAFjaldaE2ih+fP8EmXLqRVtC81QowO6JLzawKUStMbrtEA5P0EVlss/IyJ
mgJiPPBzpdcCqYuXX1mRuJ8WaSMjBBRjZLT930k0AlDbL0I6LHXJW1CNZo7iDioy
RuFUr6uj55P1LgzbzQ0JGzZMw/xLLf4Yb1mYeGoq+E7EtXlhwItz0z0gjNsbgnq6
5ksWx9D7+1wDocReZUQnCdJlw1sCuL6I3zey44Tj5LzFNku6xVyPRZrRtcMye7Bl
AVs2/aI8tKedImLs0n7vM0iD+ANIhtzslBD+bMuFa7JElqFGNWj1S7Oeom3PrqUG
AtymWPDvhB50WxHPD2+R6IQI4lX901LQ1NGNidyzg1bKOxa43bf68l/B+RMWg8yD
mEDQn/xbp2RyHTOm/3yPtF5eA7A77y9GhxICLPNEgYXkdsU28VbWGPqQxxnnhYXF
UCRoiYG1PbvhTBeG059oycWzHD3rjs5xAvAEfoiO1dmyeecfEptox0o2OROlc7xQ
WsT1AG6n4cG3QjxEGeVknQ6mJ7NSGhTNU7dn1A9lWxRO/5JFjD9TsQ//aiYZq6NA
873UqCQVHSMq13C7KdR+gLSnz6gsHPdjFAavExzoxTM8/wu79UlnsvBpa7TYiVV3
4+tJZK7dG5/pGNKWcNZ8w8N30hcXYAFX0QdnLN26DkiIbHRcLn1roIWul+8AOxEW
+GNWv+1eKuelCnC92J7Wh913296YWzdFiqtKsVAwOunu81ZNLRnYMoPIcD8ZuuGU
SFnBPK/6wro2nZh5pkh5g4n4nD4nKQSz+2V1epbqBpoGpWPL9ZKLTeMle05w8ikW
axMp9sjQNjjkDX9Anr/tYyQMoLGFJrASrbMvo+wNzeIYUSoekTlrcTwJ8dvwODjF
JtdpcMvT6+T7r9ASpqLTazZMabEmaUhcKWURaYu2Xq2B7kCY+z0fDpdIX3SR06/X
HFpJJm2rIcC7+mloiNCkzDVj4WS4/Yzr5gLFqHubWWRiHja25QQkS/jHSQpZ1Haq
UF8nCEY8Eqf6uA1Fdk0qJYN4fXs2wmV3gWcPqMw+Q3kEQAGxWth3B5xYEIG4Vt73
eZ+/Wq6d2F1HITeDYlrm/nf4rNmrOgaPDiLa8mWUip0gFTY9Lst+Rg322cKmsoih
YreJ/LF7ff1EXYDzxaeiTur+II6Gt4CJEYvfgCYlkaIaSDnrxQL3Fo9waIXTa4V/
1rbxjx1rDsqtatMamO5ELplvgGxAHTq/8IbUlo4EFJ0Ewb3a2sBnIhHK04e+pmKQ
qoJZASR93l7jX0LDczYVFpEpbXwvy3RujignLllDsNRxcZ8bRnF03Z320XaHVdfA
pc3GP1i1hThkw0bqolJ2RSrKoR5vQ/fV6LLVAY1GNwfREj+Vxar0UU8gs3Ru7g5b
chtB8nBcrcrmxSF/8H90Xd8b8b3Phf8xm4++Bfr2DW7bQsmkaqrRrZL2RdB9aXCK
mQnHWFSmjd7ZlJ5HKSuusacyNlJTiw+xmuaNvSRXrAGENBCSlx3ULfNeHXDLWLDu
dvTqIFeo1O7X24uq+aqs9Zqh79vS4gM5Y4fq2N2tTgJRjHpNdpb8pZVqIzuPFGf6
c2h8k5E0HiN3kSUplNN3Sd+w9bx+ySqbKeR63w5yCSTUuNHOmD8vw9AMTTAh6p7Q
nanMV84fcAy4W6yCcTnH4cgiRen/9yZmI/j6PGNDogAghu/AZ0s/+u9ubVufZ0w6
YfqDO7K5quzw9+FPY5dYpDQi+CcfCiYj/Dz3R+knz5hGTrlk8p3PTqwkHPJac9at
huSfAy4l1BxPWA/+iAfxKe60KjFWeZ+e1uU+k7SmFCly+h3DoQEHesUksJ0eQO35
71IOTd66Shi+20Gh9+0VnO2yO1RqzSDd9AtXtksP3rFMCXmDqxMIV/+JTJ5Qjgok
TjZEzfqy3Z2QWKWIkJL3XPeNgO7382T9etKzQpKk66PGRLTBBtUds3/dywjsg8i6
O5iXBpTeiLo2F8nWDmw3SItYpQeeMazkTfqz1hWImJciSLqPQNF+ycs6pxRqRMtj
1FaTtMUaYvGw+uOD14UH7VLIxNqrK4QwMJtUpPzIjP+N0MMhTGuncF/2eOjBisOE
FJ2CK3En6nltYoA0hhpEYqi45KwyO6QmRqV27JrJYf07YpLOxRPPmlcnOaC86CjI
KjQo9cUKThxtP1UivB/eKaj0AL8qLiSR0YH9lR9nNPWw8+mVFLGu2MZaVLglHrfK
E1UQPOhJPOqWHj9fZgBtODIV34yeZXoJab+KqS+Qo3ZfIyelOe7jMsgbYuIVLA4t
jrp0YrM7DNYB7pkN3c9NABNUS8ZxAYC+IEDETLKQtNBLzayiziW8tf67V61Jdy5j
0XTg4uGN1+w9DY0hhr3sDmHrBh+7aGnsyCyG9f94NQJnpZ8ESlc8gSGBbz5pxOlC
fotkaw/hpiP5bwb0+t1mB8xGfAjYf42wm3oob2GXJXlT9xGX6w1wP3bN7yqGctgE
w+nvMhPxnYJVh2HnyLNWDJaxtYDaa7NvPsAsUKLlhN5bWXZHBenBE0kJ8SWKoRyh
S8R4IDMzHF2nmWZJoL8qNmgdAfxHToX8fZnfOqdloyo+UF90l8Vp4jEDgqoT3Epz
U1o1fYWPUecGpQ8oK7GrglQvDh2Dd7b+hnjkp7Uh4EHTcU0uiG0frzDkWcCwxYMa
NNJO4EQ8e0NUTJqoDI7Y9wgKM3151J48pI693CfIH6VaIJeecqwKeiMUv1z3F0qE
wMYWabneG/wKAMP6qKc7D9SjTRYd7fmDdSk3N/I8xVrdE4lavAS8E2aI7UR2EuIt
VK7PK+XeEqr3EHLBt8OY95uMdpG3PGRVNSc9/rsfBA0/fd7kaGe08b0moKsQFx6v
UvErdu51X9esGx8afIw+9OkeYphcDCDDwwuGSCWoLsKek2hlF/Hz5BP7JgVwvXBA
nXLyBzlekc76wlKI4d1VUDsQy9zYzy/LiCpCYyNwOPnrDxq//YhRmkEWIx/o4qTP
BGppKheVAQZ8aid2iT2qUFPVTV6qjxt4LzIRBmXHeqhgNoT2p56kk5RLsjcvfLAx
XXWIHMcA3Vvcjaj2VCH8uqlMtVWS6o7yFCVT8VMcSIYGNJ1amwPy5W6UXLqu9z9v
B1+NS2arjtvnA8t3LutY2opCt2oCtqcCfRm90D6Cu4vlnG437AWT1+NOsRUusjvr
xeAQ17E+MM+4EWhyD5krI187bV/bRXFN4b0Qjuw7vSrH/8HH7HuJ5xfnX08JNYEI
nShyQhGmMUuW8sMvXpUM9w6Rbioxx3yFUHfLoj9Z15nsiXVyTrgVk25bLb1V14mE
27trxwXEjImUH41Gw0a7oVZNbrJ4ayCs0Eu0BsHyxIwRmprXTRWb6ZZ+7T/qSxP9
qa42JH7UThyt/HbPTNAfy200Ot4hS2msAuU6yHXZMRH8D9SOvY4ks+77bqAW/5TV
55gOeECa2NrvsSPmuV77Br2H1shZL+uZVAo6vSQ+Q119HbH+wt/vZxV+Eh/bAAWd
609ezb2ArP6IdUR2yZ32QN0xH/OU7W8rwKOcDxQOpeZcCcbfTSbhVKIGavbl/TuF
uWvwpJmZnqdwYhz5MGnLk4NG08Jas7hSVRWAtwYjrOU4yCreaavxw4DXb2lxT2Km
a6qOgJJPSYSceyoaym9EX2loNYhEkIDX/2ZsZEMC4pKzerBqqm+XSvyzrapmEs7u
dwzf9rfBUzqNX1/zmo6TkSSG0CeyTzpIcpDsVKhU3EvmDv6ojWfG10OsbIQGrpFV
1zUTk9xJntNTKA5koscUSJLHPpHUdUvOcHpd++nn076FqCrW/1kTv5qHo4Qlnz9m
iDbmdzo5KJtbMEQEDkQrZ75fAt40k03w4ZSNPxNh/c25aZo7FWLyD6+tm/WXq8Av
F5BJZmE2QvisTKmrrubyIv1sti1LfUPa21JcivlEqPBMkhOjxN9WWe30zsj8JWPe
FxhDm83wzISHd0oWAr5cf/hADXO2jvJpYlH74aJrOQGqa0TcmUy2BYSrFzNJQ6E8
Gh8xJjI6pmr102TZLUTqzFSja8wlp7icZrE8qaAhCP1O4Oye6GKMfccs11fFkvlV
qhbQrvbSvh8BsPn8PkYrNUvdWcF1QjxEC8EK0GC7JFShfwqUqFhRocqjB6I10Ecs
ajXdxHLfKR3LzTOvideRLZ1kpBOmajfLedN/ymxSNe7LTK/Fn+G1hlrHCv3yidyV
XfblRzGkPz2FjuDpKTaPaifjeLpFDsMu4j86JTvdg1UIKvpkiiiU28+tHRGcliQG
ECmRsPHI+JMiKAy/70YmfcIVwo/J98oIxqA6C8cOuqUiYWMvsVRZWQzRtsvnAJsH
vbXH3x2WF1sBcNvCX4pOuwicRi/bJw5GUZAT9gjdqKnZvNC6DORCNRi69dk1Pb/U
JMUALafyd5w7dhjmE+ND5RwT5KK/41zFw0Qr2k+6rlsYJ64/8rHPOv4rY4A25umo
25SD/QV4yPlS2UIlYGF5S42vt/KS5Cfwb2YJGQdikFQsR+CyZhtrTw5EbNpun68w
wzxnpKmqbWZtndA2C7UZ5UWQYg7DpYmqMx6b1G3v8JdJTqMbCEo9/jcURhlif7b2
LZeqVW23bFsSSyJ2zHAlfcM2AfrlCwS+kM8JPdP43J218gNZmD1IHxPDsO92uXGO
I2GpPJXno3hHQhav3t4qTQk3wBLvWM0y9o+Q5vTwL/+Uubktlps1VTRlgeNYTxtb
kootByNEyJQAt6LIFwPLZChpDkGiYVzvc+DPf6Gpp9tCu9Hw0rCKLPRwwgywRmGA
C777Zd/5Z1Asu9FSy104L7wKkoYwmwdpFsL17kkRHSfZG9VGGplCM21D0dC0+ZTF
v+/lMEh5UwSg9HhHKJNI+tYX/cL/XlyMyPB+4UfpSmwf/6FRoiqEugbmyf/4HC5n
jGl1RP5PCJKnN33R/G1CcKoY9gtl0wsyn1SJtfggmVzr2O06FmOTjaLz9CRW2u/p
oFnW+xegBs2d5uLxFEkdvaA59XyZJuCHtFKYdh490HkRc/whQfj8RFKSYVdhE2JL
07VqAgC3CR2OQAvxufgCtl9Jjiy6LYYv3V9lAvbDMQO1asGGo8qzTa84KPcXYh9b
NM3vqDGTgGNNit8sEWyxLArPS121Z20HXxBVEAwmmU9Z+m0gKAAjzZ4nMfEZ6aci
Q2j8mikQCsDH5n9LGM5yY6ZucnMQ2Xub8UcQpGrhoILjx2G9q91RSeLAKp3HjqXL
yGShTqE9OHzd5U/qSfbZlmpbwOQODy9lh+n2y2nMLVcgjbqx0tOncEHiKJtuhpN/
2hdA9AX36wnp2HjtNir7wmjb86w/EtoMDPQRCYQ/5FnWraHl0G97UeI+VsXKBjGS
li3tyGloUIMpvo4RfpoewvtvrItueFdFLccu/DOVPkY7P8SliwDL6D7UCncNWvPL
iLM7X/D0ol3jMe9vSeQssmMO6mRY54KwqRhxk1TwLNBJvDv8mT6nH+tfKL1V4bkA
AF9ATCmoj8iViB/OyDf8oBWTwMj11YE1p2Ke4Tylegu4NpgrqJjFliPg3dZM1hhy
n4qyc7EQxj6SRmx0ibgWf7Bv7g+G68gjyQWT/+S/bat0gsbJ3TQ7eupqjvChjplv
yxHZ5VMB4ZNMcWxfmC/B+mI5moDhvvHjsuwfAh4JbVKkgvE808OQLtfFrFcPpMLF
8rRrwLOn3x2X9bvtXV+z3LVxlIc+FBp/3/JwWLoRrCozX4au/Vs/6lvCjsoDCz5B
X2a5UQr+MBkUKBolfYOtTWaDTYoRaUuVmthuzVZfDlhB/kfMEQmLd3U2AHkLf2tE
66c6vc9y1Ik/RmrKpBLZknGzSKaRUQd39H+3aHpkhluA18h8YPUjtlagRI7vGcAb
8t5IhDBnDCAFbbD1Yu5KiWC53z4D4ezaeUCAqlZgLuKVsBiQWHJv3BTWH0pQJqU9
2bt1xZ1yWexrJCuOff6H0Ly1DZjGPDcekiYPGOxBgQ73i4YxS/kVtYT//o9XfkzV
YPeqgbuNWHDHQqkroQfQ/fe9+idpaRpReUp24bAxao6LhHdWfScpJdIvCX5f+wD3
Hsz+5AqAFPT/NGDFwKje2fSiE/oYfYmid1LGw0N8hUH9qdehFJLNes4X5iDIIGB9
lUgcjJyVfGdSoeQjb8n18W4nJyA10U6Cm2LYlMPbhwDLRC5MX/uSxwfnRo1lnD8t
Q6KIHTgTcsjh5U+hasMqs1yxJYauMyNVp48vy8eFxQYx2D1JzVMmLZofO08spYwK
0OUGqNdPMs9Dg8Fm/uRO4+YL0vYsa0Q/UT08xObg8dhxfMjzeDadPQqIWnYWr/Ne
Em8EBhM9q6GJIsjMKaL6vQ+Q7wyw1qvKdDSrTdSt9vCobeqVQSBH++ooTgYxqz14
IidsrfJkITRFXAvQgg/pVjldQTlP+ow9e/ZGfz3rd/FbQ4FxpR61/GIQqMq/MbnE
ywdPBAlzMc/h7PqT0bE7hcdtHJD9t3xNccBrPS2nqVxmCg0CMbbag1TYJTnf+xkV
0XwFGEhSC+EotitqP0yWFWYkgV9WY1wDr0rsZ2lgOx4+YDWrwF/p7cPiPzkfnTEV
C72Wfd8fONpFa3zZNyNCgHEutFcmtH6QcpSrpwJAmXNG/VcXn7KDvUu2eOpJKLBA
XeDk8OqHNc3r8ZbSdnRR+gPx2UhzuPb0O+JGf2smhvusbSvaHCgn/ugghYWTcN/1
NFN34+vBAKjmyfxFQbU8/W1aurgf1CZQbQTQHPKndDhwDg7Tc2mfTJ5rwK4F7zBx
66bRDU/Me4D1zNQk79ipbrIfpdesQ5OjJ+N4wesm2jqmqkuXI8YMM1z2haI9trG+
9J071xuOBgdg4gYtAiKjHiLYNN5e9j7eLmZ/gYrIsezjYkokhaxkNOXbTUgaotH3
+R2hxLROR5fk4fBPIMrvYhUeuva9FlJg5E+9B38o/7lDScL9tj7bXl6Z5xHuBz+q
sycvXGPgpseuLr4L3vZTC3FNXg91/OhKCBaWnQpSHZCHaLH8zNpTCVWvLel9jMp8
+7au0F+N+6kRQN/BPb9dLuZyQScWBmkZ9h9C6fAhKCz7kyBuxr+7tS27Hmd9ZYyX
K3bonsR2M2RA1XPTfW3+S/4268/V2NB/FRE3SYHE5xe5NFejo2G1i+uQPJJ5vhVi
1UjDjz6E5eOEdv4hwctpI57EcJVFrpaceOTXgpxQqtS8uHUHx2WTfce3TUCPcAo4
Ucswtesf1DWRFLidBl5hJtEWT/Az7vnww80GaG2+ofmK8nxqCHd2H0mmcTUfJHx1
wt4b5MyFr7NQ583cchS+6MXB8WN2jbYheGC74ZSz14PZUd05zgoF0RjA7Z9voQ2N
h2tLoYJw8+VZZ78hBPOKNQb/9FJBqq7sNRpyqOpxpC+JlNdhQm6R9TuZsnH0mrZi
Sucn2rZrc/vg10jrblRDTpW654blFB7WWDVysUQAe5e/nk8EWh6jWu+RiOiUU4zg
Hc1J84YoUNLDbZzK4bBcyWViJMKVkkv+QwA2cm4AEqjUUBt3kJZ0fEP72dXhuRIT
LXzA3Sz20csz1YHSczhRh7j5xrq5XoPGFmJjqM4nwyLJrvgVIW8hF4sE6VYvEdoB
LuOrAXC4dJBTBJ+rE/oHfSRpDJX1GDRRmzPEduHjz2SwsA9Nb6UIDtkgGah0faQy
Wb+SHslMir3Y/iH6IQLZW5NZkrcnGcmijjeMZLGME7SR5hW0g197ugm8iCzUChie
VRNPdtibb/Ey9inv1wlLEonlvi5FRea0ak9n2wwsFNEh4+HiKaw8Gyi0JsKxHNko
L0yX0k4Hoeme/pf3bjg//d8RPDgwMv+XbAi00QYead44DEj7VM6O1fUBNa1SpuxX
3VX3CtfHuNfp064SjUu5oOIzdDDr0FI7y0uEpjGxvWISNYadm6rMaxdZRDMjVYMp
iaHJCK0kIHpJwU3BZ8nerVxxHUnFSnpFLtPSDSEr65adbCF0FP1GOOZ1ODYj2/A0
znPpryn1FZNeg1DHLu4Bho5y9NqIN6sFjkA34zy2jVaeTNU2itPSa20yphzBIAH9
QBWOr1JpJ8BQqhG9zV91Hl8AfwnAPHuw1mqzbUnC/OxSxXCJyM5OYF7JfKYvb/GZ
iGaoabHuE+hIlf+gXLlbzzcVxFWt3O8Rq/zvZ4IkYAyzxBgJgMaqc3gYEvjg1YOb
V+bRN+PiTrsxGPGCWY9gtPUTcLPz0sohxnFrVJ/yZLPrA3ls8H0S6tefqvaEo5Ft
XCPOguqu75uB+uFhd95PlxGk7KXTbg39OJmC8xKbiX4xi47mcbntkcIH0MYQfZS5
9EgHPTtCwjS2Fz+BKNdgNeyrvWRHwYzfhUAEQYLAPF5GhbBagoPha6Aj0G4Oma6+
lIxqgVf+uVxmK5j3v+G75U8vwQ6EntaE8+Rpax/pyLCix0YTUsZebZP+6mVFUu+0
ofZfCzsp9kX1i8Y15isM8kVfo6v1cNj2vAJnoUkwsP1WxOJyb9z6kS5uJXqMqBk1
wp3Q7R/P8GzkcZ9w12xHz1tgSMfMVCLLRxPT8IlZMANEutnxg+qsHbvOdi8Rv0WE
vzyW98kLKXxXIczH9CpPM8XIPQqwFN+s45a6NzODgdBGu+IDdU+8kOOW5cZAb8HP
UVt/OHnkA7a6ikoTRjqHFnWi/ObLU3YKfmmNGB1lVIRVJeb3D23G3aV4+MzEi+1L
7GTWqRHQk7Y9+Go4WiCYCnplQhUhjOk1X01MVIkP702F/zLhqC+zyWJjIb46NdSa
zEOWIjpaR6+N8Y56PStpaM5hLgdrbk89Y8pF6AlhthFGuQBwF+q8OdKmtLmBqK+2
RQX8qvvLAQF+R9TW1vZNiit10xueA1+XPTmg6t/rRNd7op6G8uXF3/Yw2No7q3vl
Duh/LGbO4yeNQuHzVOzrsixoyyMeKsN68l5I7DtP25tZJf2PbB1sddpNi6F12YI1
a/XZentXHvws9gVfvt8fBeRAw5tmtzJ5jBMO11lw/0zRwOQ7eDiRweuPJJs9W1sZ
JZqBTP50S9uZgJ1ydGT2AD7HYGCnzdfsRoBs30NckYV9iM7ebizlrcOIM5xMhi+T
KY3Tb6IbgYFum1LCdNP91UJIHWJK79cQQqFE/ZiTOSnoI/Y6I/vbmsK/eIWLK3sW
2JUNhlXK2OF3LFwfJxPcPGeU0twwrLOOlP0PrtVIB5r/76fVWvR3Lp3wcsxGMI2p
RFj/Nuj86UjP51uO8CsZkHDXTaruxPGUqXlFhCQkp58YQZ6jO8nbzAVB8V8qWcvR
cTXk3hY5pY3AQFfxPgyDbx76Rps5VZ9z40vwJ6Dc1+1Hn20xbfs08M/wYDuQ6lyt
3IzZoy/3C7OWXR7cuPUPvRm3rTOQGOa7nHfgTGOmrji+KaLXAsBA+40uP5rp1kv+
mswb+zib9dnlkktYDw1B3VKm8WqBm0vm5HqLZh9enKrGYPMcjFbcDMEr7Y3cxJq1
2evY4EZ7moL502EkPBgxaOTX1S6+s/5k2KxgrAIYBtXfOE5WAhn5LeMbFJ5MKLtD
VqU1a5+ihSjOhymELgOFgJxJrvFy63Cg5m4dEgQn0Cncu82h8VkDqtg9Cb+H2KVu
Na5URzV4NAlXAsR+4NKMGy0oHlAawq/xI5g/HNuOSYbd26F1zAvdCQv0YdxsVzFe
LQZv01PPQkyj33UpZW6XfM19GXqvkGzGed1ffNPlNgcoBRrqcOBcZg9104TuDrOm
umvEH2QkY2ZirazerfCHvZLGZ/OsSJe6ayHRXzzTwmFcw+Rrct6dmMpkMVwMyBk4
+seVFqmAUCDLmDhy1Ok5kugUr06GV2K6GJyGW/Bpu4aNzWSN71v1bksEdn0MqYEF
6vrmwzu1rZapIrUMGuerOsm1Ud2CgbzJ9J0lgl6/p9qBCgQLa+xx1YSL7SHshKKR
FVXLw+0qwWfgBeFMDVCxOEhJFKBpHwt41a5PFMVGvi600ktOVjxrxq3H/6ZPuK33
iHNo3weAMQJW9xUgoXZVuG3VtfuYDd8GhictRDvYB/4OQ43vFVNDRG6DKW6NtWn3
J4mI3bIoQQstd+AGmolA99KCrb4oXihliLBg9ujCAMidPrcp7ON2NauhnQDCeO68
Jf2voGajrkCxQD75fgxdrm23va2nusjO8SVUzIW12QhJhEd8ldWIKWcNiL8IcqBu
by2sMMGR+sBhG/c7T962VwjCrEG5ClLc1paLSrWk1xrVdcSSUMvqKcX/QsmPAzHm
2XMzDi4bP/4Dwt1GOCcwAqQI7mYtnwGJig/OPDpgQuf1pM5S7KVSg5w2aqzlOnQZ
fKs/Dr6+fP+kssARcmMxBrbz6PJACYb7qsfIzJ5rJoxQfNuq+j4q11wK9ay+kr1/
QRp+rQ4NMcQ0QjOfq7GRF3c5dGgyF3Wz9iaadio2jrV5+5PrYS8doxza5LLlJwZ2
L5YgBegB9RCJyh7DOOcyJvyh7A+xW2cFesyHZzyfLlPRONLzrDcCE0JIjHUx+m19
HHrqkahUEOXyLOE4NdpGqV6Lr3yo9vIQIln8Qvhzejw2VcZgb8vD6t9WV1icoYEf
ql76r7zDbR+llPs3QrvqBpRBqDFyOnctpPJcieqGH0J5jDMvN/Ij3DfUgc6VFgZ+
72GQ2l4O3ZGCig9NjBMedR5ROpamZWIFiycTzYD6npRvrKbg23doZUySmrB5/gaF
b+fon9DAwJTxgFx76Ql+aa63My8Qc2B2KNHdFtlBC9GEsVXu/VwN75HiC6garY9U
9eRxSm9IAx2FGkHAgp/SUcTBaM/hXN3Sha/fai3k254ZS7h/k6MV0b0AiG8qWPXY
VHggHdzfllXOWJgwxiaiRH6vz5K6m5WYqsB51n4ZS98Z+hp62R0Kz8a6y9Hes1QI
7k7U2Eb3Gx/f8/1jIX1S9+hPjjQY1AnjQrJuvSqG/PjmOIkawXkiLgm0rjlUSMQG
b3gndCiyhLrFADp8YrexvqHcgOlmwisaCuoB9eop8AqvkVS5wuPKfm55Ax1R9hFF
rcHfpLrsROqsTX7F35A3O4zivrS+07j1vM5t08UgSr02l7bQrmY0kIL1CFxCU0mC
hnU015rrjYdDQ0lhIG1DY0lV/wDXlDiNPL2CSJo3Im0h90rgzYRZT7HXMVAqUUpC
QogBh1FQFt4e+n7iQTku3fhZui/OXM6QvENOiFwgEJotfXF+NkC47xhtLojtvNUI
GDnzw7eedB5YAUeo5pKdbPYkkdMtwxdBzd3XAB2SQ5+6dU7qhPL1tH7h7qpE39/M
20dYbgIshih5R105glNo1DE3ZIMWIgkaaHi3HEVXmswxFn0ggc3KkbJWFFsEhIO1
eMHTK/RvVBKL/GjSPgZmnLyuNbuibLXL+NPp2EqZO9KaTkK8GivtlmCHGCTzzm+B

//pragma protect end_data_block
//pragma protect digest_block
/je2T8VfaX6r5LZHmt8KCQjEA3Y=
//pragma protect end_digest_block
//pragma protect end_protected
