`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
LH0UX1j3lZK1DBNNGlnTYvxMeWeYSJwOGuOo17WIT/wcJDOqrJHrbtIXKNM8mUWo
wVaDJfolic/8lo1Jm42/kAYcLdMx0HD20LwsrriLUo6GlbS9lMNJtU/jY/6XLeDg
syWanh1UZ3Yge0krR/EcavBhDiYXDnMXzr+l8uDipCU=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 468768), data_block
j7EfOKVYoFbKAA4SomKSrcMZTHM2ul+GuYQjyTdI8DmbWJmAZCUscurehM3yLkGE
PrhYl8s+fgkWJYpPmp10zMpfhPaFHH3CkEieWvOxa5bdsbogVpExgEENho25nU10
Rjtk9WA9PhuS+sSZ8iPSFHyuOB/vWJCf6RzDbtY+H/b3LFoHAh3HwXw/H/HgWPoT
FKBRHlT7buEaK2jd9x7rTiSjpvJwWhTLdgm+o9+riUTztudaJLFf/GDGYZ20Ucar
kwuJ1ibnfSFS3calV91AqTrkF+Xvb6knJ9BSVZvFpxuxO82MGInZ8z2LPGvZVGRh
NfS2lNCW63zKueM5CD732UGcizCJHMtcXV7BTJqEa6txZjWJUS7EphM5KvAR4jMh
UDGlsY3QXdnR3uQOhmqDaYbze2q8anrakviyFGLVg67yT63Vs73c7pYPcQDaCMV6
y4pb7KWYQof4SMk/K9KqEiKUpmTcaN13q4/To2dNrVIQrzCfx7FoASPZxrj7IIna
McwnduSG7y9tzxS1lz/KaLK813jRUC0utzw3Gk4wiG1IOzpctFspZkYg+S9CBppR
tF1+6htwB9NxCr7IkuTr/1Fk+LDC/ZJWXViVD9dK+lt3j90FiNnTUcHygzCwV2SO
fhLfPsN6YMXhMcELt5zRDNLi276x7W8WEagtsfDdP8RgDZ241v/zWuMwYilng3t7
l9jQEsOihoOUdrvbxdc1I3jbdniOVUB/kT+ZTTfiBfgEm0otJWSa2actP0CsuAvM
lvQ493bK6OgHvXpVCdBLh12x/vSHs+OantjD6Z70ekQwMIggf0OpcQeJZSPAB2sS
EJutDlBJlQ39Sl33SwJ+PgoKjaUlP+noXTKf+7wnIcg0p7DEd34dj6xJatxubIUp
h/M6E6XiXcffMXa2TyMBud3bK9+gHsjDL1zOA901uOgD1StaPjd0skUwjkHy4G4M
1u9Lrn1j+IpMpky8+MobIX9ZEKoA0JMzkEQB5a1yhugo/3jZT9D6XkDTFFosOq96
55YHbdZs01GBKh6a/HG1lIAy7bKRCk+uxwCDS2zTGmo7Hz/VEC2P94h4/1ldlorj
Iy4wGF1EFoPO5ySXWInQFQrhMWePPxGbqJ35vLaSjb2MO6RKrtHByxS7Z89xmvaL
FxitLK6fPuHwPTHk+iAmX28Tjysdfvw23kMsHEeOqlwsH+bNUWAGzXaJ8+/Sbr8L
bkLWwWhQ3Rms/vsvU0rhtpRrLnMsHrFymryuge+b1vCSr5RsmUZd0LSMxapCS9t7
lNs4Of21pcJgPWtkV11COMT5YQQGmU7NN3sesshcja0CUV31Pdcbo0gbd39RxwWX
tDNSHeT5JJmBywQ2HfZmrZPvvB/cCKoRBpUjTHjqXGXVQWubpLO7+m2k1uI1lY+m
B8WISUvebOKBKJx1kbq09xT9iz4eT6jW3aD2SC1YYAZK58A/Kl+BUSZoDPlPIQm2
s62rrUj++wvzdjaFDsxg4+X57XmKLQq5hyd2D9FGkYX02ntCbAbycB1hdhFMUkGl
t9o7qEVRBakwJkDarQcpopAFNc2PBYXRXjTr4JO5eNpM9vM62xcdxxnm9a6fziLw
EBe9804AUyBli3BMywE+eD4HiGGjb4xVsGJ+58l1qijZbAP55erRuNiD3dN03cU2
lOAdowaaITuKfKpeZXxzWMutneY0VQZp/8N7xz/PA7uJmO8ji9IPPk4PvjlKb5Nf
iXAsHtBM1sgOSRxsZNOD3XjWpP9ct218ahmHicqtuLfoyZocTXz6q+yFzTmK+uCF
ORScXgnfDh0aaK+5kIocdu9LjMOzPzZg3emaDFTwshmrVB/qEIfLR85Qxl1d2Qeb
la8Qt2FHHgIbXNaEx85VmSGN917vsVJmfHRlMCg45bEFiSblW6vAV94wA8S6+U65
T7zRh2Hs+QTsWf75Mcxvr/p7ftRkpsWMnFKI6BGAqHlgodSoURD6RMhNLnD9THyv
+vnUKjSde3+gOxQK9uoxEIkszTVOPxD2inr4wXGQ2zmzzNGgaDmqcvzbMO/XF+BF
1zgsF3eCUQdwecQJQkLjFxuDuCqZvFyywxL6s8sM4LNxoovIG+A4WW2TRZ6driNq
9nd/Yn939cWnvZUFh9x+Fm2uLCxIngpTtcA29mCdOLIFKRiUmr10/8215mWDf51S
UXrcwF/MKan2FpBefgyAIiK6UNFdm2j4PmXjoAWAKTNAYi60EQl6WmsIyfVATWLa
UZInB1tGU6XDeSPFnGHjblT+7W/bLbhMI+HQ9E7RirTTHWrr8Jp3wkXKWPYXeKcF
rkJIDrfYEYEfdrBj7zPd+c6RzJkKy+uWi1D/ELsDu7u4COBmPrT73WI9A//wqkFV
D6uu14vZTZm65aVJV1lHvA8XJR+Pqta7LzH8putGiB7N1WKAEHEk6yh4uwJ93KBj
N/VXZF+i51CmhJaYcP48idPjl4awro5rv9NC844CZTBLghYktBTjT82SD9cp8V+7
ZUvf5HZZrPmxUYdRjVDvCc/qbwY9UDl443mhROGjYFmfBa0gOpCnpOa2hCYSchmx
1HhT+7GLtkfvLEcaux6Z04Nghkeq8YiU8fo+NLSJzSLEFDnqo+qkgoNFL/Ps/w61
u4hF8UNgdgkf/72c88zCcQxnzVeb7xQ+gshcMelIMsJNuIOd7J415Ti5Jg81OZdq
bzzVRhO7DrPJ+JSzakJNX8W+rXfPogBxQ5xzEq2i4Z4NPIeMm7wbaK5Dqoom60sM
FqiPSYERJ5Aii9BFwdSDX6N858K7jDrTYZW7vLIEsNOd544tAw++SC61onUUf0az
SdL3oQvjQZef3FT69KXcDRX5UALNPW2lUv+CWlUNOpSE16XvV/w7i5Nm9dVrfsvE
BrAXWOGZlx4hoxZM8f1b1RPLB+K1VzpeaRFJ+Xj7sLnjSmDIy8cBmhIUtnf4qQzL
h/tDLjMjfgqL4sFv4lnaL65n2Uro+A984KvXUkQq0ILxleCjwy4YkZuGbpEWKGli
Z4ZYRWzgd2WVqq3Ke8RcTmIibpG3n5GwVfOw1DmSjYWUWm40O9uNbyPpgaIOOQ6e
UmXXMVSdLX7tMufOFirHPkp92tgeNSvJ9PxQeXgCqIq67Q6dHmMknVBd0Y87M7Bv
t0pllxzc7ycwNyJ6lVDQbC3CJSLVD4nuKgnHnNIQXFh1lu/xdaMU9Ey4xi9U5pe/
6CVqDKaqNAc1XXQhyyFNlbBoJYQpm3T0EQtj1zOT8A/ZKTGui4F2ZwfDk7FnxlhP
AyDLOZyTPPnXCfGPwqxgA43/qEvdcMoJLdrtMttNJmicDKC9qItUps3lKHEq/dVQ
tGHq6fM0TnBcJq6Gz+GkhtMB2LO2mgBWBFAbl8626lXvbUIZjyUubhDYIQe+SGI6
l4uBBeA1CMd+ZxnbvdmGwawcv4ewn/KGWGkcrW2N66m1mjFr38IK4Nh9PQJgCWBK
DU1Sp9PlxyBhcNov1IHr0aBEEZ9P6WN3GsMBpHJXABVWn/ijvJRG+9Ojk/heX+3d
MZDZQRAFsNpnPHpIrgKWIIat4qAXBCxDH9luTmCCmTNmbrKF1pQwDdm0uL/bJkvi
wx0BjZQRXzFRlkwtopEyiX0/gvDoW1WmG/bti5xnUbk/LX1ac38pIvq0EBZx5Zjd
cqIlqnVBrpgRIqupIONpKfwLVBXQ+Y29fTw45DndyWfoYFQeku7MKHfgDqGbV2Zt
uj5EUY7GI5cyT9P31uPKuAYjRv+cWz50sBrAiwsp1ysxVvQ5ARSmfc9vU2nBVFG1
XvATZV4FdoRjDHEEvmhGbGZJflJKfWb632LDM+hIhl9GBihIfF1mDe6cYcQ+7mAy
DGnW+WacHjRtaM17Z1iXcV5wtB+kxH1W5Mqb4Hi0zngPyZsoacFM5pgbSpYcuZiR
vEbSb4RW2V/vmxa9tWredAUuK2FyIv6E9wllV9lPsCy5R+YIQscR3vVMgWA4QJKa
LDyBMrpZIOeQePOa91NzJHGEd53KvJeCm3cxrfXHOmNcjxN9L+AUiXPSpZ5IBMYu
HZKljItcrKlW2z2VW6rw61x3sl0Cx2kV7qEq+kb+6J++oJDzJLUWSQ/G2D2jVyIr
IL9FdVw7n4C2lSDHITUEy74E32Z0u6bb5IzHzuGy48CxXcLyMBB3SlLHvs6m6lBn
W/lgNABYe+4dLlYHuKVsGvFudMkcEMGAXp97zfqD9f4A9Xa5EVN6D5TTWgKju9HH
jCaoSbkjlF5RvZOPDsw0vkYclTKYFTFikkFl7+qKbRr0qfNih3EpSVlS8mzsztiD
oO5OIG8OeFCbAJe5b7U2d2K1k+J1DaZ8NCJVBzcbKqOk1dDC6hBsZ4AT8SWrwgcj
FEklAp7JnZndPVYxoRvic4Y/uRXtYUCm3NArG5GeB4RERFD49NW8T5JMNqSS5PZJ
sPS+5QKcnoNUnU+yFWwiIqf6ECNUQBw7IiB6BVuyZSMQL6nYdms2uTuI/b2/gTU9
V8rbpMYDF7wataj7fMOBUPDz3cVhZ3am4AysiMmQNbtYLM1y5/dZcTcKt8hpCvgw
PcGnM2I2mHbaTsRParp1/BkSSuXru7X8tnH18xZRF9fqDZ4SlqhkW+T5doVtjTA+
oZsrhCFDO4zxVtBEBF2wpzgBSl5PUMtPrtQ9f8JQ9q58BbKTKjG0IkAYwT5/jbwH
MvXEYtV8Z774Nz9HYR9Ckf58nJagzRgw6YltSOxO6CYpenbukxoNsbtYf8374faG
ARyO1i6mUhlbputnmsGZe0NgCSteHtqfv9MvNtwym6usCM1PXL1aB64mGjt/eD6m
KJh28vbgfJQGvNr4So8pihLDMC9Dn7vE4mVVnQQXNbumZw5mtWISTOBgnbRCDJHe
C/9gjy2kVg+pz1S1EVUya7R5HQrRlCyq5A8uAx7SDqD/nzUL1Sc8DW9GStI+Lq/A
DcEMVHU+aETpwA4O/Y3rZrkdJMyj4KHbKDHzfmqxOT7Z5EpUecylPSbdzBEyurk1
tUqBWKr1emsiOOjFnphLBDIt5tM9N+96bp6wpB1w2Qifv3Ro3r6TMYGgMq0gQrQP
uVgcG7tiy9qdstto2Ju1tJGtL0jOSNvsYQB7sF7bzaHc/3bsObggkPftOAvaDUr6
cQSnaobHFnEMfT6JLkadlXCGghJ7ryUNvGWTZAn8kK7NntOTgtBN3jxuT1rzniGB
fCRsAi0oOWAr5jQLSqibZvAhxZj6oOoN9qgd1DvbpEFl5HyNYUJ3H5LxDAsi2Inr
VlbRbB1Fv/cnnEDqJBiWXw2hIt00tWRDrYUaNd/Wz9Xh0bhCM6O/bBuofkK83Aw4
56fch9mUg9LaICX+sMNmfWolpNRw5VS3bvYSPFNjicKa3hduj8HkUzT6pgBn2Bld
YB4+rX+FG+Sj8EehMcI+h8KornyYmoG4/u7jBV0aoGnNh+UqO/my7IEQAPbzk++5
rFKSfTP8e6J4YiEZZ6HEvWEunZ5lHDPQ/uDhcpDQcCHCVUEVn3rybc1ZPuhVgjC2
RmQcmQQQu9DY4ECMtAnb7QKFYk9ElQ2Hyu50Tjj44wgFXlX/QFIihI6fMRMXxldO
OS6EG3hIUIcztC+vF1Xolgt48hXEJbLyCco6poB0WAhT+cpoInRwLz/sBsT9PNd6
S0an6Cw5RWuEicdqqFtIgKAuF5/csv+E6XXl7uSlPID5eCLEpAmPz5GMOJ7/Nh7M
ZVVmNYhc6UaICDOhE9hbbB0ofsle19Wr1szNvUf/CQxOSO0d2RZYvAdSk/0lQJLk
MxmGZfughTPsbnlikIKrgFAZbOP2ITc5ZUylPooyOrzlP6BhSyOWitqiF7rYlQK0
yqlIgDmzYhUYhEL6GApvp2pcO2tCNm0pYy/fzl0J85Jp5XbzVx8N5pMfee6iH8lL
MlB+rzrpKjMsUf/m4Yv/XrWnHxaFzB8UOSygqIrS8Sk/v8It+9oYsOMkEFfZC0bO
6X6hbIraJJ5EWZOD/7ogIcF6mVEgID7+EMD/Ra6RKhAGzBVen1AEYhDoBWOl2kJA
b+P+H4w1N7XSoqRWqWYge/8Shd0jyBIclvtWqmUXrUl1FlJbfjaHHrVk54Di93vB
pDfjWm9eb0rZikqLO1uQWV+L0IY25sa87mnBLRUn6e11O1ZxldMjYHbLMI2q7rhd
LtXLrRhrBtnEKM8pl7tkUh6BfoX/EF48GfFxJYGZEK04HnbYgN0VmM+WVzaQSykq
HwzIRrbuZp29fEhizrRg4wXiyqA1zltRh/jIicilC67PQQjsshputtfwdllE1QNf
4sAPnlouCmE+Su566qUDHOdKNN9XJLCsMtYpTL2lry/MgSOqcpc3DMAJhI5DvpvW
Lsp+62DR8Pe/XtwZhj+FxyeNJ632xBdT/trf7sGbnxdN4yh8fc5xaYFj4yK3eOhV
Cuhnv10eefEdLnoajYMkp3zGi6d9zMTr2xwFJ64BjICu5rtHeEIpZ7l/drOlJD4i
w4+yLT3FDG7IvYPnarxy7Bdeipu1ymXH+nqG2PqilkuJV4olnMitty6l++A6iC8c
Hds8WICI4V23FomKTskz2fa/4zsPakUWfgRsOTARcDoYYnEQUzmpl7DOybkxH5Oy
bRRs10bkp2ivXtC/nrXtsIssVXdXtuvXvPFEX7HmjEdhtog98AGJq5ewFsMaMzPV
EbCCSqZONMnlLtb/gTQWTQrwu3eUdvNya7pClqa6Z17wyoAWP3GXAQncawaOdvEo
vqWIYG3uLc7FSNOXl5eZpy5fxCyWk+aMpxTqhHHTQVraUvQ+jiB6Jjz5HO209T1V
WJMFQRiObDWDSEje+JR1pHoh3fr9ygW/ZyKG6ALouwNBx0pDCksZOAHlC66l1rEl
UDtIZYdPotiWhnUmOP0dzBi0Q7wS0yJaB+gAADFaBqDWJovU3QdDyOCR8dfiu+Ye
vyUyTf0gcOJQ97Xeethfvf3bzjfuc/sjYwUKq81pHPx6vhIDBKLEEdwVBQBkG4wb
pP5I43YFUawgc2b8J4cabdZ2ZYSVVEL5gUxLbgBCeHmTgFHYSbUsHyUMS7wYlSnz
c9PsFepVZsOwuzIgU3+fcREQvvVaWzkkwO3AlrqyXnyYk4Cd0wBFH7H15tCeyOd7
bwz/uEODIbyHbwJOVISpjdWAW307M4JVV4DTiGvFUBYXsj5u9tYQud2dyr8ggkH8
Rb6Z7LrF9nuKy7OnxsY2C9/j6UiBKGRPNsWNwxnoBBNMfAf9s70aOmVMNs59qISv
XkkqNK4gNR9lV2qiFAuL8McZ9SDy4RNVDePF/4huRsF+Gl+SdJkI7TM1tweKTtcK
A7FWWE/XK90wKMHio9HxFV4tyy1yDdUBsMp2cbJcFqReqciO3tnOwYZoI6fwvzoi
NGCAhpbRVDS/+0iH3w6h1IaWtQzogs87K5cYcnrfSawX2Kn4DHKRcx9W260XLV2C
ChaKQVcxxtR3XyZ0Kb5SIkIiRdfviob5VOkMNS4iYu/btAYYzI/FNOjr/W0CE9nx
sJjy08J9aiMwTZrFtAIile1+nQcrQrRsSiELsfLwcIHbMln2KBcWzL0JbyR+ewpd
SC/zFHWp6kJs4wmfnK1Oo+V6CSDGA6Ynu6aVAp26lzQvWexNx4K9SzVR2W2JIl6N
rOiA01kXU5NHPqM/hx7pSm4PCiN9YXfnRrz7EHnYATPXhKV19p4qn2FIzDVI2YVS
v7XJcXQmKkNHpKwW8LyDDqz8COoVm/SBPqVNcfwwntkU4tQPBhc1n/8R4eHjWEDk
VBN5zjoZ1jE49Hlmrp5mMrYKiKgKnSedbRiAgMEZub2ti7IRYyLw8wW5flT1GvPA
wDnoIatPOWLnzRrlwwBGLoN+Fwkxfi2S2U264MT19iuUWTG1HfAq4+RqZrApVeLw
y9LDU97dDXAQUvJy3IPxZSBKv/fd2vqOYlBzXPnbVqaKT6e2zWWvjrpDVfvvTDF6
dYCuASzOIOKjWJGKqhXc468HwklatS8Bo5J5+huF4eVopa5TELeygSnms72yTeap
jRvO+C+8rTrnrP+ZMn/9lhsZHy62r+/23a6gap1g5KfGYgyHmxS+nlZih1Rzfbd0
znIRaOG/i+8gNFzqDqgc0wUjRuNE9WsxkYfueSbcf1WPNX0gMrUT1r/9mA5sDtEZ
GlTIeEyCfLotnjj5Q2QBxNcwyw00xRT5+BchxX07On8ouGRD9tfWDSsjDSCj8TSt
j6asjcKbWRNlEzlCbJ8GqYhOoCGqwh7kIk+yAZlVtkhRnLQTGWNOVGDeMcGykjI5
K7cUgB7ypPwKj7FFJ9PWABGSBUXTs4UIl6Vth5//wKV+H2ZZsBvLUMAXC9ez/+Rb
JkxiShSAH24/3dvlE/FMyzVIqABHgk35iL7YC6zJ8yvcMFUzTjzLrjXUHKd1Rz7P
oJhpsXYrhKqUkOMYtHf/3osDAOaEFj3NcJCbvcD36ZYs67up03BnfCEkuslbhQlm
C+M8djFSbNePplG4NtEtD13i0AGOF8RrQJjNHA03nCamULr9/j06ZWZslZmKn1Z6
V01KygR8Ecgmp2nN7jL8Vjc98GcCNJU3KszWmSBilj+pUgf2KUNIY9oS5DmQaFay
hl2VfiXJbND3wB/2pOojFV/stJsaDx0LL7oKx2XhMQEceRQOzHycySBlPgxSQZ72
jTGm9QpXOw7M0D48Za38bCvdh+U7sYXDueF8Z7iY6QwEdpbaEOZfjrQzorb/bj15
uGcL3gnMfvW5tdIoi2Ib7V8tuaG4AMjRzh4ymJ/NnY3+AKp4jb3RTuTCC9vjpWKW
K+aAXx0tdKd3p4LeN/edrSM+g73kDxxL+Y9z+4G1iEoa5C/3ztrjSab75f+dJ7Ta
jO6H74eIQ9zDrn0iNdgKZUWIjcTJ7WiebFQCR89rTTr49wPn9/lpYPzWjsifOE1t
8Rs+tFTBg7nzRRXWMlABgioCjGYeNdiAwBjPKH+sFjvRfE2cC4S0JJinpxiWjox0
k1JCLK5jY/mNYQXulp+yJfDoYKH/NtPYv7psSoBw6aegdbfVuyd/OGDXah6rKK9D
7T62ct7a3j3RzUYVAy5mXwPEc0OcVncTDvWWqH6LDy8ZuFRF3P9JIt48TKS/bHS9
GpbU5CoeXFINMpGqAUogcnLX7p5/SLTILUpNX9Vt9NgxTqLrNvs2xAJgLyCGx3bf
wF0nyFSFu+8F6uvXpZ/H1Vqc7gj3oHmGu9TpdC4Nl94G7Z2if10VEpdKGDbG9PSE
RxMmQYgHshOunJ3TbhHfuvH6P9PZ/mMHTBCRZSZwK31oy/i7KLb1+6oxr+POZZnT
5oSiVqUxwSZX/4I0qpkKGd+5bBlIHbtdr1c0vv/P5X7+0bosuvka0jAtXVHRH93h
BsH2ftKxEEt9bENpudB1fi3UrETyPLcvjzTWi09UuS6J0uVdgeDiz2upFkV7uYIM
CSRgo+EJ3QIvsdKCX0IBQ/+KwAMYZ+L+1UF1dZ+ybAjLuMIIb1uvL8VXnXFQnmBt
8CRp1euApyIzvB29FKggyJqY0TfRodPdw8Kwa5CT8VqWlf2+rGDZI4T6TFZbgUCc
8BKrgVhBZuOfTtawuHqwclceaaTgkScfv8F6QyNTtxwsNhFf0nnUvRP79KJRAml3
NNrpnhAHrc8TJ6hwKfWfzIrnVSwIgdEbP8fPydELdSMoUqo4UBq9cRtBgwFM/R/4
fXHbxIF0RgOGWq9iH2s+x7JeWD3gOWL6N/JQ0VVdP56oUL6Hdr8a3LmiOpBRtW5O
l8a8MBOZHk9KR12P8olCd9IgGPRaaRBh2Zi99yubMQusH0Cu7Y73F8T40Vs022sJ
SaG4V7DTctvEWfrFKbxLQqv/1pAv1vsZbV59AL6QPDPSQXPZ7Tc0m1oqg4/FQH6j
mVXOb+olHMSLS3mH55MVTs0j3WY661v+SoWUlQLJ9OWAA37t6/XboybAtvQTWHfL
A7ioTFVB5Fo0pMpMx0rBvlxKctv4IQj7mroA3iitZvYH5LNjtcu2pc1oOdosGU+k
SCd4PErwR1uIhgDUlvJLEPoDj34vezqoPwgoiCPomVunPseF+isyfun7eDNMTy2O
GU/JAlHYMo9lTbltmDA8e+j9k02JhNd6qUo/Vd4lbrVOh8ezRLCqX7FPT0Kpx5Fk
RaTY8SJ2djIlSOqNCl3wgO+9wBMp30gl7x0WsPPWp79LTBKeDGdQg1pyk8qNRcT5
sARN2m8O3qTq6utlqBmlC34c2Us9PTOdZtyw9X+sTno9ucQ8q/mck9VIpU3faqmN
NZj2YYj9zAY2LAdRUpeAdHVtcXdckJJrT2NIwYqCffFvMRLdoWFYcDdVjrxBJ7Zw
8WZZU3wHPmbbF0DJONCmEKNpztvF4rZd0HmmMCy0tHZCgFYH/1EcMVd7XBXLggbN
WUz4N8/+65y7hy5PNUHBVG9veGakMsY+QHpHWlDZmCEmzjv9Z+i7S/gRPGkSoVem
bT9qfu+5js3/k/Lcoa2VrU+bCniMSe0Zw/HyQ9DJRDZB5O39A/C0Zf59SrQLdgXk
l18pUsLOdaXUU2x+0s4kF9eIyj+2FC22u8YAKzpqXY3r/BIVMwM7wKo2KKGtm16I
8OkAedO9NK+mE/j2S5+nEepnSSeFuXXrZifIWjDJBk+YjV3VFn6kWAZ7sQN7E7Kq
iUdeS/g/lGSfmzthzUXQ/lo8olKRai1oQKQPGk7b2+IxwsXbqsqW9U7Gr3oqutCj
j+Z0SKUwPIPeblBsMCabLZppqhi9OSa+wrjDtos+MZ5pq03BgdHjU1eBa1nNPc0R
R/QCmjMg9TRD4cOhj9BJBzhCpX26pleA+sczh0alRfi53q3KpyozBcVytydpDEts
Lp2vu7+VtOJctAQ7bzymYpqFJtm6PIbVwGe6PuV18moIM+jbujsql/8/xKJ0TAQ3
XGp1s8MAiEe0t9qUpoFsXiFjnAfYox1kUwxrpD7jT0MddiIryw91h/Bp08YTLEKB
Y1fzx6hLQM7UFeymn0lVwHcMyyk2WtwL8Z/pzEKYtdndvND1cL1Fv04mGodiTVoA
TRWCbT30LYIsxzaLZiR9nmC2GPBKo+zGePotZhFrWmijwecmApnRtKMJ6fIFlhTs
VfAxvr/OHWrRtEgTvz+ppmGHyJozd8nr6teX+7+izh9/EZ4OaDuC20HJeGRQWPGF
p5SiT/5n/x9Yw9FPBgrwgQgfhps3qD/qE9YpcM7/R93rScy16FuCBmQS+3H1hIIL
7Cq9aHi0ayxtTEYtHuyIbMKSg/DMr2kMfKCjsEXFGV3v/xq/i6VEJWpxcjCP1tyd
jNZsC/uYr4TEL/NKNuvKSPcpgJ1Cj7RrzmBqVwV9RUeSLE16fENP1FyduV2VzPRi
MAigGYaIodGP/0LkA3KaUGA7H01MYuzyVvII0QM3tJKFp1bi3fp1BpgP5gTzV096
1pAQWGeJ12pGLCQYKZhdbNUPCUEdDgWnpLPQKTtxrHcqv24cE2hEBMfL6/Say7LE
Le71uCjldbiDsQhA6/ffRUBHPLz7gyX57SHsbKpstyz9FB2+zTL/fAcuAJfBd+Zq
7WeSTPd9YiG4sixJDJFn/LDzVpwG5Wy3B62SsiCoZ8+Sr/suITAq/q3f0EsyaNp/
0e4tHZRZeXx+/zI3RtRqmfEIVFFmoURXFk2F+u6UMICSA6ZVaYBmQkx3ymTBbGCI
KojL07Okl9hwtkYP8roSVlq+x9QmXe3b0JKrGqVUzsvRlclQxekitvdvmMuK1nPl
Gdl4R6WmhkQZiay4ast1bc6PMTy0sBFO8b8fYNSbBqtrsHvOJfwHnN9SbmZIuirn
7fv6ujCiUS395W4VgkKBs/WCQPRw6nOya0wW0Sq6L3vJGnoyHv3EwiuuNmMmmyXq
bc8QCtMD/q+26GFg6YK4jiLNtmOZrPafVbPxgslspHbmsgSFz2vQ5EJQ6InnXJBk
yd52R3gBhGvHvbnXOZ6UewxW553OciIYbRt2KtNtPLvswoH0cYpDPUL37fQ5yElJ
VBCPGhYU/bssIRWaO245d/NKbYcujZgMg7Db9mNFupoOCkl1eVKbDdSMZnMP3CZ1
KQoSZi5qh4XbLL8SLqyPy1JLQDEv6UhqKIxyzrnbCsg16s5w88i0R7uIn1huhlEO
MDPIbv2osChPH0Xf/eJFB+eqf1ryhhk18F9ro73bcTTd9GCN8BMEUwMNUg5JKBeO
1zpTGYZxPv9oiiGYrenXgCmurXwIAxsdQY/xeaphdgxfKXq6HnLiALik9o81Qy/W
T4l1mrExAM0jux+J8qgRIqHnt6qGmAmU3pEUkSAv3Xz3XEV9krsEmCgJnxAA0ecn
muHkBoKmaBBvi0hhSLnbvpgPWzGjo8Q8aeEz3Yb6xM1gWb2mOw97EROAor3B+AJI
lxo9+0oweLcxA799It5UEwyAPiU+e5eOkd8ntTpSlbNC94w/O3Hwr8Hrpi3Zt6q+
InhycUzZikyhZlAq3MsgPINYdoyIgiBLS1Xu2FoFLqvd8xglP+JJCC0mjpOTPkB1
4sBdllz7s38LPXcxEuIxHtsvaxPVnmkJ9qV4zhBCNSvLS3JcyuUeaTScRKir2oEL
rODwm4Q1GRxKyCSOzLell3QWQWeeFeOooBjmwSijlNc0zo04w2kmCrKfZI/lo9Jp
obZ9aAn7oCUitc6K1NxSvGqLqzMjfhStoWAbrSywipzg0hGSkIYjzXe8bJJUnq5O
RbDXbGmzJH/SmIe9o8Z8JTXamyx86Uzwy0W2WkeX+6mzhPSjB21X7MqaBCJihUTs
1B7ykI4+Hvnlwasc5ogCtkoqHfiduHA5Ef9vVI6rKtRtYvem7vfUXMfmCX/Apkd7
JSEb8SrZdnirZk3iDZ+2q+GmNerr/ytifjpxEl7Ch8QafAN+tzN+bGyFHQfFMXYE
3S1jNGS3nJ/76XCgmtOgK0GLrwSuGqzAdZLN/LgXKYLM66XEI+9RDyuQAxUWs5JT
9iJZ9NA0d3vpm1IAXAfqyhGjiWSuoQ9Mj+MYin9jiolVO5idNdlmLRmxSSgHHMsB
iG5qFwBvDHa2wFSkWGcjYzStjjY1hOlucmtoNjm5czw8JSPgDzi7hfjPOK5n3WLo
boYxUYHNrvpjnEARIvdqfW8M0NDfy/Huw+Op0zYjPiyopPuUspjvaKeRsYnGZXvc
SgilmTp1k5YGSqn5VY/2tZP4k69RDqXTbH/iREr3Tdj7eR/Db3iWh5STvnbiSwm5
dKsYlgl56BAdYJk3JedRTb1dvg+VcTZw2fTpwlr5Dp4e3QruHCRsK0ZYX7IAcKHT
+2hYDOxLWkSg+5QvyDsHw0QRhnHGQnSkKld1bWMjKHpvofg3c0oG1l15f0naa6Wk
0FdL73tA2+1SEAxdU0Yj49aEd6BsHxmKJdndnXEAUZy6dBTtql5Ml5Z/qdmx+YfS
Ps7X3lesvL/tyxcgS31zsiA2s922P2jUWERGnBaKpCbZG2dmU+aegqAZs0knx1N0
ri/Xd1RYO/ZnLc8Y5egXnJyFzKY3zNBY0mVzaV2DtFYTo+dPAcINAYPzdKe5aH62
wEYxs7F3QOc6Ht4uVTL6vipqeSt+jIf2pvQGGf7jt6mT1P55Ql8kvpzm2FLVa+ey
EbkuBQsMDT0Jhkd7K6+QJtFcfb/Pub7KAt9e3tNtoduzIr4mDvigbBAZ/8hwbjcu
EFpA3s+IOsJdRbvFWPDBeeRMM3Oj+FSaUeRN1g5Sg8s9ON0buWwUgufuulJfRo4a
LF07qm02GL+slfi3RI/VEk9TuhcGd1xgcUiuPsc5Exr2rjKnq2V9wdk1Wb4Z1+OY
BEeSwg311kvUI0fOBTMMRfEOWattF5p8HIb52QvI8ofQC8SiZdP89HW0WuwbcMXj
vZy4IienQMlbgFeYZHKNpwAKknSk/HnwwuVpSUJXUkaMG2A91HK9atNH9pvpxv6U
sAuMc5yYtQwqryNuFO/EpLFxoeLIcgh8Yp/qhxgUzR1jiS2PM7eDgz1eLGUeTQFN
rbUG8mHVX3otXm8oZKxwHeiE7JNxRXnGJcNNivFBoEyj4utkZ9KpSgOxzHY5S8ih
b2rfkv+fhvSZ/SXI7900cBzaOjgMQZFtKhAap2T6SQFWNXY/kefo6LABL+xwAoDp
tmVLdGOdLSkMHfnH9lOKFotB9Z6yAqP34vHa4Yn4kXYeOnNMXLLrSluV2IpdF1vL
htLzLI4tnhmDOo3zGvYBSUD7JwXQ8kRHjxEV844sZH6t8fic0EckWp/6pX7F0dMZ
08OAexPdgblMdR5nz0SpuihBxzf6uB2+XDcMLabTi7MzvjLoPepkn+Io23QHPFfh
LSxJvRedSRBalesrUkRdLrzXCM7vB6Qs5whHZws8q0A4EdaDF4TW3hqLOAGG7TZU
rJLbmWuvVfan2hYFKgDkbMI/giNsP6Tqf5fvy7f53sdRip3FyOctFI9x+Z/RmMW9
usCfYTPNnzHQ8cgpmlQFheZaETV5xP8Nkd/Gs39y7x5zFL70hRJHwQK7n22D+J2e
uJuczE7k0LL8xC4ikmOOVU3Pt757UCbmyUMiCvvE5dha2lXELCZXSAuJ/p+7A9bV
VmZrRtacMQrJk3XvCT/ZVdkXRAX4T7YcWWGPIPv0qHoK76dJtIQ7/dijaYgUysA+
g0GCKGULhtY1qwSD+TDReFdE3Q/fHFDLVPEACCoG/FWxwfUjgAq5U/1l3xzPUt+D
NSo9pdwqP73JshfSYYdrbndmgBamlbTJuuN2j6tNc9owz6Hpd5hWpOvo6c1agWRa
kzf79N5yP+e7BaqHbNf2es31rG/1SHlG3ahgQsQ5Bz9Dy44ghT+N4nGqE56JVG+6
o5hOT8SspuYsUZa9m48/Lx6J9nIt8Ya/yVL66vTaGFElJJ/JoPv4VcWE2H+1hIVs
DuCXM1Pf2/BBy1G9Nx+CaDpjFMdY1IalMOiUTXeVhqyr8jG8uxzkppAuSiPJPPBJ
/iX6TKLA7OEW5LKs6R48uXVaLwUfw9OUZXFQk5aXh5Q4eGx1NSClvzn05Bpgui6C
jCPX1MU7M+zvQcg2o35B9nVqfowyL1Z8IgoZqEelPEw8SdOHC0o+tYilyO/gieAg
3Bj9dHOO64XAklozffp6t5qqIXApJyf9BdgZ2PK2dqeL94sxhEcbcTtUv4kNL6VR
QWWHmsw6qxD0LLAG6i5EleMZKgYa63ykFHZuLkXcUQxUzzkhVvFeLsYjrlHpcgl5
ll6Eg0UPXD6oAs1nbcu3K+CWggAncUfeo3HXP/IAa7l0FTaLg2icTauKI7lseP8b
JZ/kIYLict1nW29cnh9yXy8KqUDIO/dTNZRax1n5oMDhkkBRyRYF/4VslH+UyAWU
DmHSWoSAC0fkW46EyvAzziYDzdCgS2zUgvWD27xnsu+vdAaiLcp5ATHZdHeuK+bc
CCAeamRxBIrkpB9L8/ydiMrQqktRzGwBso8Dk09krmSpAMCkBwNbKzEINRwWbNYc
L9iPkORi/WfhI2k5+a/JCzRcTe/koOouHFiRFPHCEKKnKttQkX9DFW7jTPrrfkRl
2G+HqnM246EFYBpVSI8T6DP7ZLgdBsChr1NzDFflxBHJgOsAFaIlw94sJHIKgTs9
Czz+mgWsINHVouE2ZlvqpjmDIQEXyMwg9lkA195HcYFrYqDD5bmp5EY1ZRorFOKH
SSOb0xBNJfQmRTFpKEz0lONqDT2v2lgIsRNOOPzzLp+RyHlr3Bakc8bkf+3N5L6t
InCLxYbAKDo2YwUQxA6Qqapw3VREMnKdq32JyY1psJ8TYdSlF49IgfAEfgHoyqNB
ByhHhGZmFPprJxL8wxAlFZoV4uFOcCNn5OKufudGQPteB9dsWmm2KM/+ZC9VQ/To
1U6Zbl2VCyQsH7jOkUqz6CzqLrLcffh4AmHNCtJTCDag209+sod4JjslG4aqJ79H
nK0MxooW6bBmAVfeLP8ecr/FQYz3Xj9boZhdnpQyxXOeZ6bEYaJh6rBaWgGAqSmD
QQQCxtNH89A04iGiYQ3SL/6H7HRVBGAVdK08Gj5fJU09JYTMAHx7HlunxZMdM/hd
uQgDeflWvf7WpKqmqZeI3UHoNrDUmZ5D3/6LBKo5b73N+3DTIoWKvfPVZ2QeDoLm
xbN0h6H8SnAWb5HIQnqp4k5ZhQeeFlTujN3ihy1YwD5LYSwcJoLQBlfHrBOhefSR
TJA71GyG5acF8tz6j0dHwVv82txQEHhJdjO7yM25eOFMHIerqgEZhEq5Ghd+Xf7K
w8zcGEcLzZIq0vVmOhJWwTkIgPPeELBYW5qh/WFi+p5dbj7v8mK9OhzCiOP6iXqO
RECYRNdvZeO1NSYLROjTzDyRLki6rzSmkRWIpwRpc0s6CyaGTNxE/ZJUOoakHgQL
MUMKUEEYab7gJy0ZjbmgcEqoVNxUqxV1RpcrWqiqvbDMhzESLunHCok2FDbaE1OA
GJS9tkCfegeoiyKCQGYVyjOyH2aIxarzGUPYGa+2T+TBZTJ6zvv+5COUS03I0iOh
AmXsp77nPnmrW4RSeSoZ6oUQlROP/WWjIe/LGG0QASPfn0nic/UsYc/v67YXfXie
Tc0UTIsL8491CoOdSKTl+6mhwz7ppsYr9sdJ4yU11LBvUCXY7JjZHE4//rGWVTSx
OCl4uBEnXXFlKf9XjNOWRC+0kmU70oo4cmkxwtKKgIlmYeSZiWFA5fgdrt3G5puA
SqHXSHufCRSbFnnPmNuovFYpeBljPoD9AH1GzYN75F8bSPEWICDKK8w+SR9VVh9u
Yb4EBKEgmVTCtV8C9WYVlVWSwBErXgCZwi3RlZHl/8y+jlZyoLIf5X4FLyoeybSP
eOPc8+OAWLY2Qy7lRhUHuub9EUOoValiX9mgyyX+5KesElhnNlvLFYxvH+t+Z4Xr
zGA4QcgA16qtN9Mp5g7cund1D4RW3etgKBqE3dq8ojyu9kBodB/iKtWQVvkBVkf0
L5LfourBHw2TOJPj293CNncE3QKq6/NjDXAa7TL79fdWfb0VpQip6OyKqRHT6uxY
CmxQMMdLl4JsYcOVGmcBpHBfAJi1MhYXP3zzFmitxn/FMqKkiYEk6bTT3E2IW7dp
+L1j8GcBv3RKxteak1LULgyvlDpSLdzm7glE5d7OvJ1dhplFOtDhc9AYVGkLkLyn
jt3VPyT69bSrWStyo0EVgUnw1oWl3lNC9eFBGlFTXvF27iT8xLI+vc4HttI5gZht
/RQA+j8AG8sfvJGBvVecnmThhAoAH6fI5qnJAS3szZzFfV1fX3/f5Qm0980tSsJX
ebX+lHruyxWsnuu2SvlYg3RIKpLWqy7VKZc/uwsH0fQHyug4q9SbzEIRrRa7CFKX
eA5YI4I9nR0aZmuUQbvwv/J5X0lVKShBmmYvKcMqr6t5K7pxyk1XpoREmBbC7gvu
SSwwuzEi5P7N5d8xfVYtVOIS/p2gNkIN+5jSJlE/+ui/SymJx09osx6iMYGB7wyz
B60iQ6F97aHudiLT/zkJeHoaBeuUm5xFCW1tGaTiqIciEwI2XV2p/Je1CeUR063z
UqAFjB39l0q6Jnx3koALeMsYwB0YdTSK1ku7EeyEisITbtuF/uo0yPiwbsY3PK3K
zpyQkM1fyPVCVdyQnTsflXtEjURHsCr5t6JeB/Dct4G0WMr+hoyUo5jd6RZsy/+D
N6+ZW0uXooRxNSi1hpz2nPXlYHZogp/2KnmVsfXgrFje4mLHn925FOo3TQZsLosH
tvDyqkEnBs335t0ZJYNDC3TvHWSdnCLoPC8E3UkxwjwWXrOKWVznCpNlYe/rP+mm
/ZYm6LGikhuK59nWzYCtZDO090Wb0t86qe8QZIfCYEQaPL3C888sS/Z/TNJsta3v
WMeHsqLMG638ntqSilhjnYNVEpPU9qZUqO32Oh2x6xsm2zVXn53LB4ID5vFBJ9+X
Gi31ea8i2pUBBpyvxYt3JJ3zTNFWsjJIVibUayxPaR2EjrECFx49qSXnUA61049a
69diHoDCxJDQD9ZViapsTNazQcawFOejklndF0EYf0nQGE/NhCRdQ6w59lCHDDT8
WvNP6XpAdTewh6ua8ESjupyumMJyIZW2RZHDwELzLtj76ExEs3CRRV645cFjjRI/
ZRfJP6X2w7M12IEHGAN1v/y44AA/+SU8BfRTtTV0NCkrwBFms4D2m/uSXMY5wnHX
BqJI2L8D08JhCAxfivnmB13jqsTRHOKhvvaNEEvQHcOZ3KXwgEbI4e5UZ7dhkg4R
Zp7As9UVPiyv1D3pxDJLDkBBGEmb5KTl5X9C/VQKbEmcImfnpidTrbKG1/1G8D/T
7tK3JNbdbE1rMR88PvSZhieIzSupvcpyP2QrKn9RNVISvlZbW0uUZ2DKXSQTrqR7
5BNDJ2jTmnHQ69IAXHm4Kw6rOhFMFjzhAawbE97PKUbGDE6H9cR5F1UnBN2wmvA/
RzDBx/MIga1vgPwH7frbJgWcUobP1W5DrBUK3B0Y/X9xUsAPL622wIfuTmrb+aSy
4QuQ9txsL0+CKvmBmIKUyprd7Ob8O5zlZH/HCx2DqIkeTYTPVh/udAIhli3wA7JP
KLKm4TGU9/yNIM3VnQyg+Pg4wWlltb8YUyGgepO9Vvb3hLlYzbaeqfx++Bdu8VYR
OLjSPhs/5wbHpJDMzKdPMqpPpGDjC3kz+psC6YI4OmMyahctDEA+5J3w4rg4Sp9f
Syc/3c0DrbzWltJR021RPaCEvRahk7Inwcu/R5kqs3CPUuaKekPg8+kAVNQ/IaD2
uGcjpDWi04v3ZgZtF9SY8+ksgt/odrMC6Pd3ZxVb2qmLyDzRzpwXmcHnZ3ikwO2P
VRvMiWjhUtWgioUFtI58TzLoEDChvBFRdihRY+bMWtU2OVBpc62rMaZqsjAo4MWx
v18fLTLSgrfMUN9/2UxWKB681OIJo5h/PCLcu3B7s1GR8zHta8GqhRXOuaRanEau
z8riqw2OLfDaNBzb9Yi3Yd/8Zxbko6aWLHM6SDFkUhnlVty+vkdhCIdkbgdl29/8
PaKrDReVEhPRstX2Wtfbk62y0qjFbPAel3s8z+7p/S1+iDVZ2a4gNuYXJtGOJp9O
fWMHiMYxFq97kr6opFh2XqaTj9mJHSEWj16IPwLCv2mSFtILSYkJTsTdlYerYzD5
HC+SFDwXqMnEgjta1uECYf1cGGpx4BEVSalbRpaUwWit2sCU//d/I1Ae2OvQS1qy
S1qVPYaIRXEKNRX01egfT0Y5U8ysL4b6G+SYTgdoIadx6gRTxtVCiR18h5qLYB/Q
a7ylVJMlRwe03l8ZIvmDI/SNkqbKxSrgXr4CBsM8ScVps4SK+bSVz81olyPAMVxu
IUV0Oxn+mv4R2i2lkW3GnU1iv1PYx5SddqzqrRCx1ZzoxR1tgo4GP57XFG6/l63u
T5pTyOmmBNneKiEyYnQUfj3bMlYcvR2YbPyYy2jtsQ/TgmNlnoPlxgcTJ8MbjxK3
TNAGs8tjoHEHAdulz0GeKQ51oUlwrm4r+q3fxSDyCbRr/6EyMiXGYetgbNvOZKAW
9kGJLTLi9Ic2nr5hkQI1wcz6Q9Me4Mc7ekHPHIgwpG+ykVFco0AXrGXyODxTjkLZ
hHEO6WGp0rL/i84EK/hEKc2uIjwvJpzF/bkwyCqte9KvhXod+FMfGjYRvegpWilz
Rfjuk9wOwagqqnw5+VRlkkijHr9/wfGubTAsprPytK0GABH90NZX2hciByhMH6fL
RoPcbLSdwVRDl4JIdueytwuw0NlXhlfjRLlSrn6kvV/SBUTauusWcXOVMNvsLDzb
TFO3fndLDlh2eWkFJFZrW2AMfxVqd4gcEhZIwjomWjMF73fv938wOGoaO0VyZyIG
s9W6QSNT7bTv11DNNgngo55w2uwydEF/vzOG9lmx7oAJCN/d9U6EV1q5uV0YrIAA
RYnRs+D5W8tYAh1kqi/T6uFbFgj9l9cLzQBiJApEcGg7ABOD3HITiSOiOKgJxypF
VATTwxKGuHWwoJgJPlNx1WBjrMtyQHhavs6GEMNxU7aX0vQMxUsgaQsCcc8RMWlD
psOSopIIykE3hhSakeY7FFzjKPkRaiaHkQcpe20CrRr02XVeakFZFR1oQqEHB5Zp
qs6LHoHRFxwmTElvukNNywYo+nOraFleUKSSjqs/AGWU5Dc/UXoSD68UqmhnXnZc
K96rqy5sPdOKA039cGdykGeQPWacxfXzoJO3vfwEN/02Es5Qjzd8LtXBClpL+L0P
8Lvm7crf2QN3kz60NMmAYniaZ6Y1siERJ3S4sqYM/u69t2/CgTy+FXyUKnwIp7E0
qogUUiszPXY4GeAwCReQYCaqMFKBj05xQWkxjJIVnSG7x8Td2JDm8eIE6pi2yxBd
n/QjR8dPDJ0KO2UfJR8MYYKBuEABeQCA6vL8BlpYR6AysPc73gXtbfmwJCxDtj3n
q1rPrwA3bNmtPvGLDe7gAbuBq5/zmj9IE8pXMdyPV/XU7lRFV++FC6vaAi7tkqF/
TADnPgnUR++07EM9JKz/neAS+riykeg5QbXFs+cHHOuOzaE4p7LOBS3F+idaq2Nq
qYoXrcr50Bc+r6lCP+8q3tCudewQ+qVE1qZDmNGHv1JIUpqHtYHtHak8EyBOi1eK
J7VP4TsQWpQekMEkwx8w1IkLQF2RQL/VefkZYSyOa/1WzKkJn3HJQz2+Pe7IxAsQ
C18I9sjwqf3SKGIrJmz+Syy66ip3jkP0XssntS0KEY00zRuK4UhILUvnJ/avJMcr
rT2vIoWeFFMBp3JU5eudfwmPcACmQsyy2CGcNS+fCd9pMK9huFrN99O+5ZendyK5
DAB+52JhGH5p78lp6ayKrgcxYNSidTpYkyQBsuPEH4Xe4bcp0JbBdIgiUeNM090b
/eL3XuLJh00tBH5Xprtnq+SSCV4JBiJ8x93gQKpStkQ15rC9oAXhkKrjFcum8ztf
6MPhuxRb/AQ8B3iAUVANS3u71HtTXcedCa35hJiATyzO3ldE/58tcr+wEFkP2ncb
QkIZF3NKkUI/QWSbVziX2DCB+/7TldC1Xosv17lyfICO9PbFOfea5Fsr75Z8kyev
zbG3dwGCXgu1UdII2PIb9qr4l719shUrFT3hBaJxiKpI2C9bDyhtq/Tqg6yf+4xg
v1EXo5LCfrpCCk12Yczda0g5wb7pvYTO1RjyHpkx/UDGdAfAui3NdwCIyEo2hXtW
CDDtguXxDDjQV6L/HQMAxEvWLmhzrtNUHoCdejXUKVwT8CjSm4jy071eWXAp9++y
8EBX0l+I8hLwGBI1TPcP8GSI5OiG/bWJ8+6dVjyBnB4Jbvdz2qtZm5NmfaYSyV3u
hU1SRXxYRNcCIV6wtAgY8+KB5BBWBmiTdy6bfUo+fEyeYLLEXkRs19+YuVO52zD2
yONOMRpswjH0FLzdFuQdgsxUHxkzB4bcQlcxboKq6j2dTNQJEYGy2z2kuN2cFUsP
/f+St4PQ4BXFNd5YtjYAlMpqNOFGENgQCIZln2kKHY9kmv/0lO3GtFYMozf+VwOR
MiqoQQajc6sHeCq0nPNIr1kFmNVZ8ubFU5QZRataJB9LEpZzfVZ9+vk8UynG8kj2
b/M4RQa/JYBiV37jxpNkwRRbeTDtzp0rlUFgLzU9GVYj7nvr3dPkj2/j/KTA8rAA
dOrt0IghcmRvQGEThL7iF7J9Y/GKDtbCAmD6PcnReE0sDDkxy5IooJoLkjQ1STfQ
ErHiZYU3rXpbfEn7/YslNK5pyGEG2QtnjJ5XdL1UR0whI+3xICJcj8dufqhW6Vtc
CkkC6KU82FGlbM+ftbO+xiu7mdSUMVTP8mry0k8OdmBPXjWIzFsa7oGP54uz1J5d
aq585yD1Jn15k4GLkaKq5K73+Q132dhyGaqNnTWQOxJbPueikP+OWmCc4vy5ZIht
hcaSODCx/oZsPXW7gFgh5TYSwKl7wnQW6dL1WSq+GiCC/eqZ1IREI1gGGZrtxxx7
2Qd07enktTXBtkkhWbMP7ji7va2KrUjMFbNYo3P381PKLysPeuUSTXskR5NYw+wA
Xu/EKpWTWysF5XrvyR+baVbpUezd5/D02itT9jzt9ab0qylH1pIDr3Nlrm3qg/Cw
1981Tbh4DD7gFR6PckxHJDGHyUa06Ka4gWnXWmDwIkFEyG/AgyTnNw0GjIGu99cD
yKeU6iKjBaD7RZdImA13V/maAQB+Bod+iemUXYXgJbm0Vq01HQ18gZPCoHwLLSI1
+pJCV3CTiT2JemUh0eHlTYibKuay7pnmxD6fEZb2kcd/C8SIXF0OycDX2T3iWx3A
yEksEGHtCJt2i8zmyLhJAVLh0GGeiPKoyowPUqQmUB984ApSjYT9qDl4CUdalgh0
0UX3BahZE9DKE2dTAJWs9Utzt1H8e5cg62fbbRiuTdzErIW2lasL3S3bj9ZQNDnK
u7DjGFC3lfMZCd7eyXkVO7Gbr4AMtClXOjG+WACtFcKhgybV9y2TfgkUNAouwPE1
6ubCTgGCQlqVkjchIJ29+S9CM6kXkZpXa/BqFsZD6RoTusmii0zj2qfyCEGWuJ/V
YS/e1Um00djTmPQxDw/oAHTM0USlDllPz03FMrYqIV+eFwFz16gtNZgnd+IE3okF
gm0NRzGIsA/GqQg7ZNzn2VwAMoP7Pm8FZdexPT/5TxUMHzNp66E03FbBFEuWF/AT
MM+70kOI1S9J7wedQtXr2XHGDAPf+pVNZedO0Zh7LBQFALDOnwWGpcu/Fb2TZFl0
FMaMD3vOy5WHAWqIFw60A0lZnzt+yTvG+6HOVdrO/o4MIhogy5IsmgBlt6G5pZlR
E9E2PjiOEq6PEMOxQYa8XxkIq9T3YPW4QejHtUzwKUg/a8Ok8PqSnxptLSOh9+hk
xpjqrl3jeDy/D3fdP5qEtIzfzRyG0MWPqLwN9W493b9beEDEIlp/ysNhdXgHPjRR
+wQ+zavHJPv4w6c6ZI5BDvg3CKj1dHtuUrSRCF5g/Ba+RbOgpXUpbYZG7exH5ySG
lNBNmhbFuhSZa4jRk1t6KaBk8jtjVvkwY/uiQMLz6avn9wQ+MW7Er+K+/s3M/J6j
0iDWDYpjIiZAz8f19efWuk+gHiNy7AQMtGJB3If9ZVNXAUHdwN4ol8iEyLGMd/4H
CYRVZZ/pDPkNZKHOqrjLAXBW6o6GKUlm1azrb4B+rRuW8x0RFmCwd/pImKylKS3S
b6MgsZ8Co1BhxluD5gFMgVZmHJ+1MKDT71bxv3lV1ZashFmLO3berUZ3KT9MF2Ug
UqClnVgv7vAWHeo8uQsJs1DZucMZMUaZTXHHoejy1zhJ3JvUyLJd8TnlJeNitg0C
TLKOWHFyh4Gyuru3f9dr0wsEjx3ltGrpgNzWUBlYiUEnWPRIJh91CqBJQtlbrmqV
TDIEV3j9v/zs+N6DLH+6I60lxgyn4l/Sj+lRjV5v+mqVw9vwSqIzVNT6PP1DmmuH
y2vDR6mE5/JToQQ6lWrwFbcm9Jr/T1mLQFFcx5MCz3Tvlsr03tAG8O5acpvwEPI2
mfzhze9URU/hQJ+Cq1HhXxMTbDkMlzueSppnBA7ias3bTRg7Tqfmw4CDwckjCzZR
zZtIRl88uPpvjFULJbIfCgtMS28OnXTTTRXPo435sViBcwIqOvDZQqzB2xPY5AQj
WlZ+2U7jXBrmLQqX2Ec/8AZiLk+tYkZCzagPFySoCXlUM4+YTOR7dLzt8C5ogpgF
8hVy22DwZz5dWJLTNDFAqnRnOQUVfm6J8tCWUeyAQ8fpknClI9blgQe/DitQU9JI
x3EC+5YHbOBNA7JFqEketcjGBYmFSPm2wN1O5lSFDzb/K847s0gZboOFISCdcIiX
qbanfHYwrB372Ihyou05Olgri9OlWJ/znQjozA0Q0awMClLid5UYn6A5vvW0LGQ7
oUAy8pVM4uI9lkYrfN/hK9bcmsUHOGL8dnhjNm1ji35L1GCbQGFq/ZOlB1N68Hok
6k8C/7EY0EZ12x1HOLRijCA3PM2HUOOxCYA2dwsy5z4zN4NAvpuHmp3x0oRZSqBU
0+VJd20AlVzKQHiP0LAFEvvPi8MQch8cGu3Y3AkD3mXWd1Sd/EY1+XDrQcwy8Vb/
ng6B00l8CFY8z9IcxHlvSQZwHAv+RD685VCzqGfTIe8ePWluJ9cfBv3mi38SZvM+
P1lUuC7Vxh4yJ4sEwkB6Eipn56GpIilUhIt0XrTleTKB0qYhmsHrR+MKGH6CM5IR
cLi85kbXZuIrF3mJ75S8ujgKKSpcF8ZWj/X6eNO9dvnMIjRgTiMeKrKUyw5Bjk1I
obDoQ7uac5HysILVREriKT31a23gp00Q9QkkLW9fhr7HJX77ixhXqO9TplwpV97R
UKDQMMYuTtopKfm/YHyx3y0PRu4Tu45N4jR4OQdA8fIP1aNTxMDVev0mhcgYLfuP
k0Sf/EdJyjAdxiKr8LAEeokEVQsuGRiBNu/MnpXex73he2o0lTBbyLxOkrqhCanN
gI9XcuLr0zbpQ+vJEnN9Rhv75Bcv+JWO/93U/z7wubg5UrmyzuSKAl9gaMmRyGlv
2oOKvMLX9sy+IzMfdg6YKlcZOXrN2nsb+NOjq9UQ8+j5R8DelMe0lYf5q+Hvb4Xg
ionJVC+UMeuX9k4sHlfJY+VUCB5XJyntgewOjJhPV//BvRwbO/j4YfDUb2gEy9AF
IaZLOsC+3UQf5REmjCsRPZNwltwtti+yJh8Mg7BXMQ+edRS2JUsSYhuSaMpMiqD+
zhbQ8zrAZMstMnyXRot3H1yFm+qSLlh6BLKcc0hvlE8FlG6620UsIG9Af791jxHC
VaOMhMrb5PdMjcvPp6Ct0jMKDDTkfKtWQtHvBAA+epsPqoy/I6gjZthhmzx2J2vS
TY/+SfnxJ3f0oCZqEhF8KqnVaJN0QYSBzs4hRdeKZ01SJQxMH4OOFbFbEDv0pRPO
Dwry91a5NZILxzz4d6PHxYJDZm7w1HG78dtZIEHTXJHSA4pQdz1ajOdpw3jnUjsP
RNXoGjez7pMLSQIxnGRUfWYGczh7u1awb7IQjTM4BL73RtN3GtWHdGJ82PC4obod
T6P7H8VjLRpG0sADlo8vQ/Ijh133QbwM59v56cND818HSh4H9Wk1tdirIRhbYeTj
bHHyJmCsjJVhM/xV7Z/+ZS1AaHljPa9SFl81gHDqMK5qHvvF8erBACwnt7tay6go
8LOVuWObtHsg81tFzJSIIe7rt08bb+oAzHrVLOZ+8R7nZXKvlx/ZxaTcsOt1yDnv
WjF8Flfh9eSVLumJs589LwDPCUtE0+g0jiJWFhzgTykvj4uQq04mXwRY7DTVKsg4
kUkZ0lBgBtzFpvGiQ8+dTNdX/ypaQKogo/i4Xb4zPAaLEQHpmHTbfcu976SALtPN
WbEGzggWLM2fDwVXrg1y/vmlfccL8E8dwsFCT5auEiuksFHut1QUUL67A9+RbhPK
pY1wSgI9KmDl9VMqoqiDyXj0YKv1OXeV1TKbZE9WV4nC6qgxhSadgRAWBhWbWuNx
WBVHzsHEJcU4AVa35LD1JXKiLgPyYnY4P0fddoJ9FslttaLfw/BJ3FKJC6NHspoL
OsATbLvvP/iaz7LgX7gmTGJ28fzmM3v6w7EBVQVoWXxvC8jZioycRwkrQc/E9ZD5
t/NyRAc/tFU+EmcWnkN1Ar4x96RZMFmgKXG8x0DNJzrvX/NUcQJ4l0GEslJnu2Uv
VXAu1DUyRTea15A9gj2vz2WPOy6kAY3VHlrAqs2GpiCPJ2/GYj1YiZUzHrMEJ5by
i9OtQy4yt5BMY5m+lE+aQpWMPrmkFkAIdF9uRRow1Ss/qS8E2BJtcjFd9u5nKo0v
gXh6AOB/ZfEVGPxrDNwqG5LKQ+8D2VqgJTytfd2oKLYFLmYrSQV3rhMis+IdwHsp
ik+zaovGlH39xSSlYGvFoXvYDGC4ogAkz9mycdqWT6YgsZ/UBB3PFUFxO1uRLx37
aPOH9+qV1146/8fqaiu/F+BEPEQDirWM24dnCZA6zYG9vwObB9qasCJZkRXyDrXM
bp0r7sK3URByz0WpxBGOH/h8kk+ZTwTnwZH8uY3lHYx2NlRK9l2MFbWoK1EVt9s5
oel+8vR2P6vEByZKEv9hMU0n3Vg24boHmoq5iGAkC8T4m+j7u5ZUIk0qxFxGQmkz
QVuIlrFLWu7dkzOPH4D9nvmYo617XGRLa3vebSLuGHHzLZdpDc36dH7Axbcl5MUZ
4VRdxOmJ6Rh6rFCQA/7SLbA9V4LIRtCJhphRoA1/VQCd7ITe4jhINHXM3dsCRJ1O
cjm8Es2g3jsbEkWrYsOVKqdjIu60YUnGk108FdIgnZQvfQscorqAf2Vn0AbN88dM
VZAnxVcFejM5Z6wUwY+quZU+p3Ol2BDjfjU/DvDXrDa+1SNNvUKy48oyjhHhXJO9
k6sGiTAnwRL6/zzpiglJ78fnsiQi8HFl3M3b0T2uFaMbG4MhP2aMGJJQL4iD7ID3
7XF8SH/iV8VGVTkUiMFWdjceHzLjvkZdtSaIXm0lJowIuQ2j4/sPZxbkbis2dLR7
buto8Z3t0kBbtg9hBeyI6wG5dSYdDtCyEKuha+GbBjqMJB7Lw19g9TJPQ+4SnYVF
tdTpnMGrPx8DTTP2Q8DmZ8Gzx7tuEf47/uo6UPRKOxgUT0ebcNqroVBWn3IvCgnb
5d8Myfjtm+1FtHdqmnr+Yt4nyDzYFZdimjrt6jvqbrrgHKKfcHcmsxRgpjnn9k9u
1Z87f3BP1XXpuiTbvleaQlREs2RpjWmomcsWNRxhnbUqV0BAh+JY8TSVro5Jd+xs
+aH/IVepFgwp3rN2JuJmsSCqq7w4SaXari/26GLZmwn/HTR0DB3BseKk12sOnvOB
09X3REhsOL2P2KASbcwCB3EncEJztKA85B0TCE3w76323dRDBhZYbTbgtJn17U9Y
EwoONQAo5Gki2xjP6h5eEqDnf+1e4RrDeEGU5B2gg9u3taE7TuJyf4w0LVRrExAE
ZX9ICt15GMXHDSPfp1Ib+qrmNFr9Wb9ImxZ/K1eNiANDz34uPtetoS+bijgG1HUS
vaR/xKjWx4BIAkebg+dak7k9RlrHPY8JT5gPTMvWvdztXOfsJMDcvAARd7BkSgVZ
FiRSI+WEZJ2d617lzgtB4mSe2nW11wo6meWlDtUE6QuUDa7EBvsEq/SfASbSlVMV
VxB1atNgaahEh1Mz04DQ6fieeTFvQHwVqaYFQ9FaXf+K9Wf7k2RNBqXmt3d+pYtD
SjtwJronY3ymSILLXEQVBpB+z4hEMD7HYxrhE5FpROWKFF9HDnmNAacY3mhIOS90
g0KJ3crRNNWJRXxhlil/EE+1S/C0q0phEBOyejK/1m97hhp8YJOXWLCGgULeGYFY
WWMjCROXgxsR5B5DnOob0KuMO7oEiS+oTsVK32SZ57OMhJNp/GNpnBMFlLyP2opb
M0k8p/PsI3ueX51PREhuzM2IgpampFQhtKnnEkKvDiIa6cCuYrXz7nN8rOdsC2Gh
nnNKeIO/EPDt4qtmEZSvoM+2D16bD70Xcki9hKGlNvm4fNpxKFvTOdnTxovhadKo
Hr1SPqzFZ7fXr8Dndt85Ofsja0mdvf4Eat1Kz9hQ0tf0HzbECOgLsaeVya5caTTY
vR8LyLq12f/Fg0lmcp+56mjKMT5PlKt0kz454lT2H7hHzmPU1mhhR5AyVuinWK7y
WwDaG/LUdaGys8VdfLcO3eoam9LIE+3mIwgfmKJUG4f/vTqJCSGf3sq1rHkAiTPq
rpiTg+0mmrvFec2d/XoQQof1yhDyBfTn8j4wpHAyNfvnqEExLOQUJDZxA5AMyiMK
yYMlt3meSGfQnWv9U/zR21yZOF5vUzN0xD5G/tTRCiyCBVvnPDtyRjzZU85lJGvR
vCCNnLhJ75GCNnhk5UZWROb1IEUX3/S3CDOX2aJfSpWu6ygNxAPk7jt25D4bN+3/
SYns/XvzuYsAsO9MsuFePapza5GF+dEfmrtkmfXW/OyLmV5A/THNLj17ycFGSeCV
3Flpzkmomk2kCdl22QsbSMKj1ubzsvJ/2v1Uafh2vXPLG2/N1rNUgWqvQ63SpDWT
l9yYXNZcKflFpVWQR19uNbP9iAsR1tyljpw9vj4s8Ys84PZeDLiXkqtnwTZj/NdH
JudTdgeyE2LcHeoDx2r7m+0Ckd5oZwOfWSkgtI+dezqHT0hFOKFCZhmzQRdeftBV
ADo/HuOEMaSQxOXRMunfWZjpLXVejt37ITWr4sk9FkOVUUjQ4tqAbBleDOvOcql6
Zl/Jxr7X0BWk7RYHtb/nAWmvqY812R/9zxAsDvejF5q4uzRIgvAMGUAKlXNFJpa8
bg0Z7j+UASJ7Hof8xxUHlNw0693/sxGoNfxV4y8RL31ENvGt14q5iEx0ERgx0GNo
bj/DEnIm/4XNegdXAoiJ4xLsV6G5gEkGXF1898AOxhXfMytUtNt4MFoYjt9hzdRY
R3znE9a6ZETu36jP2eGzo98ysMocMjtdEWLKX2SkPwHB9MF1LRLpIspPTdE+tRnQ
aByVibPlNfwz/1M7Er9PtZKxzLWm3h3dKVr1G5faQEWOJNVIp0LuRapWw1FH7ct6
MHetlOfVoDEaRQfmM1KTuiGq71DZSkmzUYfMBllBt8QEro49HOPFxjUHwm17MguD
sxU1PtlfaI9VNBUPrxS5ALKHAMSd2kWVaQszZ7Rxmmhn0Mu+Hd5da46dWH3xijMk
Seqe4RRRfCR94/KPlU1s0rLKAjMUsXSqz+/4iXH7FaaipTDqBUM4M7I46qopBj8Y
uWZwcEa8K5mj95quIhkD7g8SYpmKMqq1h+SrRIuDl64tbC3yVCyzkLU2Rjj3iG4V
ND7wwlSt9vchqVaIaA72hJ5/Bxed34kYyQdMHgC3EYAHIjVoCeHm2rNd40PuvO/v
MP9GM7whN0eo3X7ZmmgdzxKY+daAtPGAVyvcEBh8bYyqIA0yhlp3ekqr0dlhR/4K
XrpvlAclXAF+tMqKRrl9GWg8ecKK8gErcAPm5f/6zb8At4tm7iQlu9IITYxyFK9/
4Dw2Ia6r95/EX0dTK9SOAwOApH9z4Hk0ak1qSCPdn3JvuDkGmUGhWCM6cA6RBXM/
c49F3L/K4UlZ9yiJld09yyhQM8jGlLkcEz/tZ4Rz56fc73t5gEuLF06pncZRWiFh
N8MCWwLvXHB14WuwDCY5CbmsJpKIqoD7gQaZQIW2e+NMvQwBYY+vO/ws5bBcdfnT
MJ42mXDXu4KKGD+S/1ezUuxu6Yjl27asdlF35Pe02MAxAsbL7PVd0+kW50IvzOUG
GGnMlwji0csQu0PpMn7EqXdx9PN4X6BmDv0SESFSY+WH+hkE/Fip8GxnVPYDE7n4
VHckWGfoIDf87FGmpl3M8IAJ3Fa7mQfkwESQWaB9ddOb1pLD9M+ytmlFkoZN+C+f
v+n2phy6EPwz5Pqb8mqQ+uI86ge0qmES1cIP2UxXje2CSLs2iRe4NOMmuwbN7DhJ
2FNydHmra10Vs6EGsvqfm1aAC4+8gLc8fLtsautJc64Yhr/FmgD0qgOuEd2ZP13r
F6YKgPhTjAU+dCdGtI+Gg4NP3sodquTjH1RjaSq6lot/2IiM6cU09AK47wL33T8a
4terFXUFUWoxgWnnEdr9L1JyQMAO0uEUezo+i8zjZzcmufuAUX6hsGjY9ubAABhO
2kO6dqeK3IdHd3ZlYgvVR+dwDlaJSinS+M4YSA7S+KDiPazuo1Nx17lz2POqd816
ofNmnnivn3QG6/cfd10erjUouE4K6Y2rN1ZCCMH65N/9AqqEML0ZdETxOGrsH3oT
d6YM7ghoQWFZV0DFR5e3gRzb7/eEvb5HXxt/8b+9XleqR5T78EJvfPS9SF6ZcZ0i
tbKX4WVy6Ust/yPwbh5afGbZ9gBFVEcjJF+geP1AYATCChF2VdSYsjajq+0SfpIE
y0sC9VWhKFAsQNNTXkCPnzHpWLTicWKnTN4T7HOvfjxb3SwC007PRGTScPz8FSDe
WnDnCdSS58tgjmj2+fEM381qAamEaROi6I/76U/f+DpkpWdihbX1KxLGStchnZK5
lSXxNOk2G6obfMDl78QbegXmDDy32wmXkUqNDuSZR0JXADIv3ZV5bMBM4gtBPS0E
T6m4BWASc2URxPi87CqQhpx6zOoZQdyW3X6Z0NKAaBc81XNfX7NogPU9uV4bae5j
JrQKi0qItTVygx3X/RgKhBJU3ElWE1EtG2Fh8aAZV5tVpu6n6zqL0YwX7wYQ9F31
0p9V+M3zE5IuKsLtsJWTFSasDUON1QGvVh5osRvDIAL/XOvlUt1A2rwDYp8XZ8RP
Q07TIXF3WBkXSOVJuYjuXlIFR7h/BiRGkUJ1VkEKIZO9b1TS5ruyrlORebWuJVTQ
Z4XtU4Ef4IStJ6CKo0RH2cUstWpN/AvvKcTj8QmKtxoDJ+W9F4tpcw1iCJP52W8D
Q1MbbDBukAvNgeNACUlfTaZIQ2I800Y5rk0upZm6zdTmx7p8dC+pk7/3oGreBTpt
p27cmjcC7UO+C8hqdW014JnsIh+sFc+sKQqH8MGKJDM4joIBPyKwSvT4LdaDfLP4
j2avFfpDdptv7Ez3eq68hf8MV5HgQl/9zAL9tAe7ddGFK8wjbl2F4Bg3lJrTaTkK
ScBnH13mZv6jgOSTPV4R2JyD4Km4dREtZzLVxr12hx99Ou2/UbzTudax1l7ZhNS3
a2laSqlAG6B06/ri+0x+dGOx9bbNkfhLixPqaOhWngbWtZ4qyiuOyGu1P/FylHvJ
MihIywy87nq0CdqsWoh4VJ6gFIJWEjG2f9RzcodbM6bjXEfEhlb/G5hKrEdAJAfY
3Ji2EvbYI35B935bv3CQ/DWyGCjuFs3tpAggmF0adOf4f5AjzfQ+KNVwV2PE1hgd
bIeTk+eph28RVqaUzDTI9xTBE76Pt6ZMbLtOfgBPujHQCOTDndabLBC4LSoBzNbS
R8aCva07d6K4XdncRg0HeapOe1y9SD94Fh6z3m+o4JuGUd8F2UwRrosX2FQtxeNw
jXDYOiIldfZ4kOZ6Fbs+QpHAx5KV9f4Vx+U3bIGRwbm8hPtB7qz0JtaI5Be3KGoS
yQkRgagwbrNLbuOG8vz+JnbruzjABffh4LDXsufUmBKvqyXjiYEqWbBr2OE5PqaE
9z/NiK3k7RETOfy7A1qG6XxdxQU3SN40SClggWkS+3DfHP0NYzeKtQxwvKzY5IF0
3dyRJKa+tCtSAUS4xve2dtre7A61A382QV09oRMUzEULeitRTdSmCbGlc6C85wp+
kIfoT4xuBLjpc7EAZDnZOh6CJZnfyg9wvKHxsS7D0YPQsSkrtGTGZOn6roqaLn3K
ZLuSUkMloKhBdMcg+fEmDwITRPrkOW+d+zwdvQR3ZXBfNQBmzacFyZaBUbPXH3Uc
W14f4Je6ECDYR9kq25wrj275/FrA02TtV4yTEU5uOgLPIAqLnamlC94Hafwf8ulm
GK+T2P6XtMpQTs3RtXoxSGBh6fRrrNIpG4KzN8zMebGRcd2IJ7c6brnnWbifgVq9
tyHTV1XSyrn9Y7baznRpPvEKx7tREXAV/YEFBAhgVGOiDsHLOcTg3smXw7WuP+Lj
zBpqQKvnV8yyljI+P8pDTfzh/JHZGQqE8DiQEoCH5/OuIdEojqqVqfIe+d+u1Iwb
E4G95suSUxAghbnQIKgxNHe1rtDaPuJzW/EVYGQI1X9g9MPdrYLpSIF3kTqbMcub
16G/zLRboKIeaG8htU+dRkZkWKqBRqWWN//nYwTR9VVgsFtzm+SDUaC9I7ILpNV0
lf1R9R2uRJJyePEOsfrGZ18QScFD6b9dIo1rjSkIiQ/779YLM3M3WcGqFr314oy/
pH++mlCZDAGY33UcsC5TGZravXDSma0exm88TlBUI5r65Hg46/8mc96LHbY1nbuy
9nxiLgKtOZqd9t9WEGu7x3HI+e7+WrATbDcSSUDJrKO4jJjyLrAWVektFiMIV9WX
iSdWuC8vrAD++RmYVoQMTtE3mmPXjYFkhR9vJ/iHHCa9o+pATypePfGOmZW+kl57
dUcY8lTYZpAPvRR+3yFHvf78sX9cspjV4mf16ZvYjeeMmHZgMu5QSStqVGR+9mWY
58UFkPTjcJpgu+EUQTtvhvz9mex/g9sa7XxXuvsmq4ZDBbx4bypIkJHzrvYPq4LP
KRTXU1M7VLOQxLwEbCnbj5cOSg96WBt1Xrl8x/9IxovXPSyKa/3Km0i89fB4W8eb
oPCeti8/kRSvOggRmO60WMSfDAs2y1QwJJqV9Hr3aScbMIbcCnp8hPwOc9Jj9wc5
yr9LC9FwQ91v1EVhCDQjEVYXZiCUuTIBR2RU2+1eVBQWa14sbs+HzrlyW2/sdl7U
AtnwUYNQmj6nWQgIVfBQ1hjYL272kJSORsdREe9x7tWEMRl3V2AQJ99KIJUd1upR
K2ZivZx0lQv722eMN5+CMveKAtyrTm4IV0BkeH0JkHqm44NYuCyGjMVGXSEhUesk
sn8GIp3lV31T9dqB5gg1qgxv1TO8BVDQLDWgGZF9kjPDOBJvtIfgfVmGiirjmows
GKn3oq9I5BnsGps4Jfap8ZtAdV0LlBqLTq8xqCzpWAB2dapfjxXcD0smS504kemj
+NfW95/A9YVQ0vwBIbPgHp1xcsAmVpQeji7kVXAdLFQq4tLxjrEnYayHeNkm3+HG
k5nQFi6/t+YvjxZ3mJQGLAvSFumSjDR1Dc5AEISOhYY7f2xP+BVSrQ02CTedgXro
0BN+5/k9M8jTXCtPFqtFKw5twsCwxQzFI6QfhDNenu+CWlhf8qraoI2muP88P1Xl
d1rr8h8MrcD/xKz5XL+CIV8HgE2VYZa60WkYojm2nkgzmsVXq8zxDVrsluDGknld
2LCMUrVzxzOEEDZ0HTIjM3W5H/0lv9UruOXzkNF5SVWJt9fIIedPh+G1SOFeigTT
aWrJOZZKbJ3JsNMoWaWojLdSJupsmmAYV11SMxtkjHgJQybx9vDMPDpVeuy9eNEi
sXcw21njeisHRkE+5AIAFoiX6y8AcPRF77h6bJ9XsNycHffk+b++KOHQD095ur+n
ufwaEi2MZBXI1NqNStmMrX6F8Mv922QXbYq6AXESmBCwWiPjrEA8ALUFW9DK/j19
F+N6v1lI4XYld31sg5uI48Aba4S/kCm7zYqywE6qCMwS2NiFwaJi7X0n0rr9lkhj
bD4DW0gZ3glsg08KeQO+xqriSK+Zw6qSAO9oy0mVFRyZklVBSgdNOzubb1WkXgkP
4lALXIbuXGDeohMRKvuRF2/Usf1Fas91Rqv8Vw4swz/1QhoFcgwbDiVd1OQEYAhO
lA+xdmoGG2jaBWDNqWYrWSRbTEeYQxzMIxtBds3CZviwQqr1N9UJTn+Ta8PlrImW
pEx+kTWnw1bg+YKEXwZeQR3tILtt+WgagxNouZ9sVFOEDlpltLBrfpqa4bDxpYol
S7pdaXL9l0KOwGpLT3Ere6HhHCMGPD7l/m2QqqQRXV8fhd/mtgJWsKq30Xv56/mk
tvnTvoyt1VuwrxKAgzu1pQFIF+LR8jOwn3oHEZZbjNTb7N1wyLtS0qz4Qruy3whv
HxfBkA0u1ajQVAVtS6xTBUPT72/4jM5l0AFbk6rieXK7cbJ2gFYM/tC+Y6iXeXA8
SdgHjcUl/TfYDb92UVYg8DHgRPUEuky4htRgwE/ZzFIbFKoeFIyeK8LW3ljWxboj
+HahXzXPh3w6n/yRAUkxn987PYmJtL3r3o4W/xzEf/yGVa2NI9kXpqU11V9kOW5q
/h9bSAAsmSXaOW6pKirW6boCJ9R6hN/73oit07opewmxQU/Z7uWjdNdOX+CkxNlJ
rOCAON9rTqK4jISXVkKL2GRHMf2cWlQs7k+zl+9SMgIdxy88YJZkzMc4NNmJj0i2
sj/KGY92mXV83NiIAxn9c/3sZP+Bsxdcdy25M/YW2Rc2L1M85fZXG/eJf2Sf8tOW
4MFCTpyEMffXIMmlksqAIkryWfc8DqnjivzDy7uRPSduTk1ABeODpOqG4Dy76PAz
lggt6BYsaewNaBP5ZW+Zj+o8Yxkgcu7sGan7s8bxDCGIpywhEt+tMqhHngTvje5p
+cMEwgsNGLKwMKW6BZTAgpRbG6ihk4Ulep5ty0nYUie2kmG1gabzWvwAjO0/GPX8
fZLo26JXNetf2GLzgHVX3RPd6OHw6GZUSy2Fg1l1+vVPqtxJpo2KTPcH+2CaNck8
9EV1BWSdRKRSkXtntwR6PDw/V8gHyDRv5rtlsqrXlstqAuxBYcgp45qgZTVvs2Oi
nS/8KW0QesRCHls3xOefYQa581crcxGrGDS+/iglFY0Akq9Hlfc+vTqX8mtfdPds
IHgF6TZdXGVBjSVzZgMsmP89SiTuFCYLdge2CXRQQHDYLfQPS7n+kvh9xquuSCPU
NXTAiW4JoxR1zj8Q/ZdmwKd6G9M+K96EVRkxx1Dp1aD3yCvh5QA4gAy1H2TBndyC
oiMEHuoCJ+yE8pGqnCIpXPIedkmVQCC+pCMzQIAu6YPQqJrUUIBT0bzGXlFAL+2y
E0bf1EBp/q7VBhzcm3Xki/UI4JIYRGX1onIVFxq1FJ+cEvqkQm2pfJV72dP4pxNo
kDAPOmZ6Q3jHLBmQOoSnRWdX3LsAQXn+SxLYeqSsLgTGepJ7IZfTAfvePNdN6grQ
MYBoqbsvS64DAYF+yMnfCvyK+bviM08215ej1ih8y1smYmCW9iRQSA9MOFasx2jT
N6e7SgXYwA65JF6vQEmSFKwqF8tsqdhQcfEUPNoB3ImT+mPNqrdX4Id2D66g3ulZ
7qTEJ0cp/3Epji9uVuYpzfTDeeJQjCwCBBQPMCOgUj+FBjfq9og+ca7g/KsZgSN0
FFb/AI6AALko4N58M5GS9ccXsuUNiE/JigxVYnSFBAY0a6Wb7B5rq6j9ONOzqbSJ
RwtFJ7D5RYdi2mKmy+IaSCiyBS5aCU/KaVUvbZrVYm0gmt5EG78nnfneB2IMZy9y
4sKF9zDI6ivnq/6GB2g4mlHcGdoEJBHqm875cVItFtjNgSZEJSsPQrwUVXuC+G4C
rmQeFfQhka5l9uVPzxGfrvXhB1RvuDgnQciTndgiQjBi8NDhnQkPgqtzSfOCLuQV
CdGKjjtkBz80nT5jWYRnOjZN5LUurV9LgLSyze2R8oZ2N0RUL05cHszOD7mbIGqR
qpfnRN1/mncXtpe8GkqH78JLtr3EpYSe8GIds7q+sobcr2TKj2Xlqr6EqA8HwOZ0
1bBNHjBpLEeHGikCOvkZMg3kamwF18mXz//vLE4V90ATAKvJTxTDt0W+FlBJbZS8
KsQhzZGGWgU+Jh6XN1VlDhOMMi5IPUDT9tnogEk377c2LhpIGrvGk0/SUEAYlkaq
ks7C47AFVckTauXoUFDer98EyfiWPPyos0CjPuW4G2X7UYfT9GDmD6vCdObM6pYS
hS+RO3vqvIthGpz3zVCzpOgNDNur2qFXbiglkXEehfLI1eFQjQNohAwfKuWyde3n
1kjwDxG5jJ3lP0JiZD/wMvNclm05bnpIIyNqTNcXw39mOvPl2zI0A0gh/RHaOGu+
cZpTRfKHX58O6GD90rRvS/3Kml9FQ1HU8LBgYBJwvbPt66r7yjFnC9kLDT7rufs5
Oh03EyaVUzH79XJw2ZVlrwUHbScZexy4NoOZ4OCnBlAWJFqzMJXqK7wSskU+g23+
N+xaNc1jnGue/BrHKVCHZRK8+gYAwqYeJsP8LnR1q4xEY8t4XO+M+gXK9nM9V8tU
BHewojOe/6sSLsai8eMvcFkMf9a2/E9afDsR82CXBEjY2Va4E67agwxRyePkxQUa
ij3AiPDFUnELPTdnnJ0wC4ZeI1wc0lM0W83z5qtoaZ+h1TP8kyRs/cep3mRgO1R3
dewHXgZ/Nne+jgQkFOynjUt1K05nmYhFG1FsNeZ8GmcB3asfuHCDWTz/g/tiKXBj
w+2tUJB02OpPJr4YkvGgvyvkF4AEiXPxoET7bQzKEuyEfCXW3TX5eHoQVKwFTZ+d
YtG7fNzhgh5ER5lOq69sgnkEGQLiLVNqS8bv2UsumaalFVBCViWnMVVVOuX7XHn1
npA8JS45p9NhRXLZ6KdlYPBN6+kmk/4+vXLKx9ULgRuQDtR9oV+0zUfeIaWmcM91
HF66tPWsnhWGIw4Xg/XRwuNhBja9TcYluhu3PA+UR97kyUwG4Xl+SSahkRbYgG79
4dW0joe2AISfVPOeYdNEhAP3HFtcijFWaeuU4oGTB9CJeHUHPCxoumIIjDrW8nBl
UfUzSQ+VEiH1Nt3B6ACrwGa7TYxzew4Yky9AMm9sgQko6MFXIdd3cVKKFIoJHnu/
Q+mPBJJVkLcFIZkuJi0GVuQXSCpdcbr6h3CCVbNwlwJ7K92DcqzaC9o/pc+YMnHY
eCc4/bgIOcG+QrLcVNTHTZvvnB+vx5Ygso6EKt9QLFQkWTsMtPSMYtDituiixyCT
4qa9PZpxANAWhS2yG2u53Kd/QopL1ymiq/iwSMMstqPFUsRaxa/Mxtiq6wcpYzsV
toIGc0vc0oc7ghLNcwRjhjAcmDMlqmgdvoJ+eD5UhTCOhp4WD42Tp71YpWXPMiUV
Am2gYpA5w/BDhmH7yRAdW6GP3X8tyBKyuYfA83gyU0meglTbODEps4Jc3dSaDhpq
kRsHgVpw7/P7JrRKmqAfOrTlaYchCxz1H09zjtkfKEpEY1TeA/qpkDQMjJ+/pwkC
uS2Z/R8HZa7pzj9LZpbWTkiK8Wg5tngjLqBefyFUb2qkn8tHt7Dx2Z6J1sRyOecE
unKXLBrApSmLfeP6H/E9WSJRvTsUwEn5FKxGlo7Lgd3AfjncfeDGnDRDxNOBHmlJ
1XkZ8Iy8mU902ZjU3WRQbCTGIIR//Z++ZC4SeEbG2KUp+nnV8/1dB2jxkJNV3a63
24V4VahYQCKymA7l/Gll8jhJOIHquTptfgAXuebgVJqaU4fn4246m3XCb3Lgw5KY
YugT/pLI6aaVF3bfHYFBg0HbBO/bGL/e9xGLmsUk8qCK1MafS4HGW0vaZZGpaOhi
XAUiEHeFS3IxDiIJpg5GH1Pd28F3zU86bUi5Q2RS4QsbPjwJvHWGYjIZJLq4uZ3i
Wj9k78IvRNbQSA+5tBAeGtZwCb6AvCRGI4WRoVRaJfSdGUuJ4/exHu5uJIdCJeY4
0xX5ru1K4iQYdQt0uT9HwARK9fAWReZhNqt5WgM/vRZokfOK/WdixLb1NoIs8aua
lH1jUC97rTRk+Rhpejpr5CC9jf4shnBlCfCGo7trXoYa9TNErEKg87/8YX3HhF7w
5WO5ZeQQ4Wd+oTmJJhe4OcVkE6QWEeN6cpCkAXB13MKu/teDLBvDkw8iHf3wqLiz
QRox7MJlFQmUdAChoWsPqSaeFejUSKBLKl0yXs9Q8j8qNofx7pydWc5jdtXzaP+n
Tvx2shwTkcTmPEZKaHK1BpOZ9TcckbmCv7fEQFKQOA+zmODR+Lf/bfVamKGEG89V
3B5LCar+FPjuzpO3H/946ropA+dSyPEAfFpVAgA8e07Zi7xBQ0PCpvQ4embWE3gY
iCB+zDos13i8f8VtH9m+KmtKb/2wUVKuWiySCIR99aez/vDW/FZ66epVibjGCKFg
xdFQcNxoXcJKVH2mID6PyZTschI7MxCzlqRs4LCHMmEIzsD8J9tDOVDWadXXgGJN
n9TQD3ddfqLjMdUNPUaLpIUF76jTcYgnZ4ShKEzWPWYQniJpSMOs8Hw7wAkO8ZAZ
jDh4D22V8oL2JiY3Bt0d47afPDZ0dx2NpcY8b78HOkm7lAmpWFrmX/itGOw5Y1AP
B+qCqVW34SaHK/wUZQV2XTTJem20miqLXVOAy87Cw0DcoJOaKFTVpqVA2CJrJ+SA
cJZkxnS+59i8nK1dd0OGhRxKG/ZW6PUglxrG5COfs4pNN1zPWQma1fQz/gGuBhaG
0IODWIAEBKPVyVmG7Cu+UvRvKPHWEHf2IKmoRJSTXbAIXLVe7kI+VG/O8xULYvEB
Udc/BqbtvS4gV5+7CeI6/0dQ4GhWuys0i+kCSXc8wvMdKAJhzAqlwTXfhVKc74cO
71rcjjpM8SGs9WBBWjGrpNbPmlOXjA4cbsaZyHIEeKY8Ew9GZPwENXinsYqSsR0h
uMW4SqDZyppMInev3lcF++uJIVeeEYYx4g3SoHg0QJt3iBtPJANIVvHhqFdUDFwu
Vpq7JCdYOnNJPCnJ31XVDau0EcmyWTglgN20FJMVRUkbaza/lAqC37fU6aiTB89R
kDzay/YOhtshLvGJ/UwWkiCQAmOo+uOLrG7Hq8DH4IyrTb8WfPAsaV1j8vNZL6VR
+2n9FWi1+9t2ytZUj6bHE8l9kZZpCqP/aVD4l87bROHNcsVbywjraamdtlQZqOSP
jwdk02GzBLhXxbHx/SBMmJgc2XsYaMjgxayvhhRGpw6A9u+8K3G/+kdQfjCXXsQQ
X3dC33OlL0em6hk+kq57zLjO5rl10tMo6Ge3UI2IumxEn7N2qf83ebBDrL6fnTrN
0emOEHszw6j02aUwoQ2qnEdjah4xVePDTT3qkvGARz3ep0YoufLGfZIhStttqIWS
j+S8+pkn/CN3OBL1y1eaqGAIaLupMUSh1clbgpQ8E+yzHTPhU/QVJ4vUdxleV96j
JQkBaH+ykcz1L9C6Jht9HoGCbRengw5tE0TDmJFDbd/UqW4GxcZRfhpUASpKtPjJ
H2Vht1vMP4aWGId+hGKV/ley4zTLWgcMYeJRmAJjsyPMxKmkDwkZKTXGvB+2IEkA
dmqQil4Q+MSa2tA3UYGUGrFMcndulHGEp2TaC6cjZNgwUa6thGQdTJrawMwynLiD
/JNsAnvNj16xgDIdp4GcSeS7618+35WYrBY0DVhOd8c8HZNUztn+CYmg+srvF7KL
tdSY0czVEytco7qayTDawP7t9eGjJb4n9SLNzj3XmLvidCnMimihwaCa7d1rCcjF
l8QxJkzFDIqrKWkZHsmKpAhnSPi8rsMgL663K6JpLgLsePU1hwhONISgBCGPZOsU
M8FMDX/b/G47eRHgoAiqxpL/ei9AvkVfUVCTiYO1n426eHOD3/jlm1nnlWwutgKz
I4rWxXVzz7kd77DhQNzO7vACro9k2k86nLDWtuoPlimtLn63qqaR+30ts4DwWrcM
cQhm1s5wKQJQ7dlKhVYvTPdWbx33S8EgAMnd7FCGHNfrM4OJHTjjN9/1CnRpFzNc
sirvEOVmFYbsKVPX42jGh2L4xUIN5ghg9CoPhvwbCwiow3X0NL2i0IgtSOrbYe7C
06XkIPMQTap5in+ch2HVHm1jMHVKNVV1d7mWH0FsMN3b4tcjY5VWLUM5VKeOBcez
SKrC9nfmfdCqcKp5JdV9n2CpYtBFVdT8OvKPqSLL4i4EheDUZik4Px4NlO7X5TSx
8FiN6Mc1Lcp0yrECj/ubgWLbyQGFaIJEWixWPfFhV11OCztasZaeFK48dpWHQuNR
jo1tI0VXShdPUi8EpXJKI733BJKuQu+6C/cItnWmoAhRg0pXC940mdCxwHHLYHMt
Ntxxqj5fJ8VxUuB0JKDvWBs6FJlBI/ndkNuUHi9tKuqhiqhqJSPkBdNDgU3yCO2+
aejwEKrT6DFb5DtBardqsh75VqLKvsUO6Wh3GeYHbrV/HKTfP7PxK12uHcyvip6s
ga7X6/6li61uWqc5XaaSxuL6qpzZ4NTrkfv8KHKXC6h/iP5fgmbZdBpoLSJN74XM
Qj4wBIEXRKHGpdDzEqt0bvmj2D6D7luhhchLk0Td2Awjq/QjTdbdY5R4S/je5NII
0Cevo4GQ4G53gnJwhaT7v5/MJwGh23Oy8VL2Jo55tM0lg0rTd7YTvLjwPF29z5jd
mV838i6mqp3itcmFbk/j8VcWYfPG2+F1kLtwue/h+WCNpOqq1x/OXyrOHHc1y/7O
NKXxnj5Q+IwUuR3+8bWFML+BeuG27jsfr7I0IC0GolmATDV1RqqGyFoADpxX30gu
cqjWl9cmh0hLn+IT/EZ5oEdX4WpU8Q1GDhyDwbKv752cZpi0YeVd05gsrzf6sAak
jxRb0IpJwPcEAxVTCF1S0220jTl8injLK/x+cT9TRJU7NLzfZZSGe+yXT5r2720m
eOObKUx1OlIt+YAQdWUJvsVYEioSNrMZdijgY845ROGAoggAl3Imb9HF3VJAN949
MwE+QHsX8eCH8SPhwv61EhNcya/Q1IelyvkUdZLcsbCD9HzA/dhIJn0ng2kIoirI
w/5AaVoJceQz0xNdn9gVjc2lHfd9vjuG0bgQjPLXehKd+XA0IssDO1+R/8tdzhEJ
/aCd1eWKK7Hy21ltYG34ctbkUGlXQaZMEOL4CM3ivGzG3sjnxohiGy3d12fnnTXd
HoSscNOYAJ3rvOK7lmqeurDxmtWw/KxDyKS2tdKS7Ovm2AsLkrqPrSjJBAszIt+h
S0BCC6NgdNuHoFeYewWv/cGvb+f/pBg+CUQXVgpdE07Wr51hwPkrHf8sN1PNOFJW
S7hyBrplyOBQplnNeZY5iC2m+W+g+5l60oME4xfpXjkV7IUFgOkhS6+srDy+2jOa
E8ClgN4M2gU1sBJdQYai+zF2Ra15WvPnBvHsn9YaAfQpU0pmNsaccvnA+pTAyP5L
IKQCDsxWB6iebRKbO+FHRrxGFdpwfZQyM6h+xKC8QOBzj7ZTjlOqp08rHmK00ZkR
9lvXWqoQQ2yuGNtxaY9JkKUtxwpe0Gh6XPPhe8nHdK3QXz58CIhoskI8OF10wFis
R9DJzJ8S9ngNSTRw5aeBJjGBjPDJkzkdtfTwjdGITiDECnN05WfaZniXqyn0whmh
8NzO+IKKkUXJAaDa8uve0hse7mOPgTQFgUtR0Jd/3H8fPwioHP/w3quxtlqbBtAh
R5j+dL1seSc08iS6OkTsPFkNmCSZSkvlvTwPdpWH/dc6C9E85zx9D7fLS9M+QhPv
05GeQyb3F6Ms4AmjKGM7qqJRJk37tscs+oIX6glxs1uf1iqLc+MNCQq8YVAKB1MY
4QaEzt2fg5eW1NwKryLWDLMiZ3IswnEzve/vkh2/CdZNHYpPD4cDiI9uFOCbVCGq
oKFxdxyc8/ljo7N14A/IrV5I8fT0xJ3ysXPY07QIH65C8a50WF4/GVTh4EY0HI2R
LoK8NWzIPoqje8auKWU48Zua8SIKr1FoY3RlrXAkDAf8IbdHujqHTW4PsncsO5Aw
znuotWGW6sQ2O+IIdNP+nc69g7dvY1zUJqHw1xEr8xV97FqYMa2+h2Lri9Psh5qL
l1GpWqBiABdKCWXff8XP37WEc1bukLqNjX43pswjU2oevD0L7Q7dhrgsRlccrfWI
u4K89fyWDwVnYFa6Rs3MCvEJyMYwqWyyedciDifX/DFTIvIcmGhEnhwbZlLtGDCg
5lzBgo0zVWWCB94s0P0wFWT0r9sJEaikUdKA5uLrbA820O+61nOvOjtncCddRYWJ
VZt3Hn8n82Swxyv3KstmSmU7l8Ei9rQ/bdqFbS1+ccFf3hl4xWANF9odnXHEeBOx
+LTzmthuaMCt7mfS1n/RdifTAQ1bdoT+kHwnpJk4RNZLHMYU8o8BRy9kugb8Y0eF
U5vWIdH1MAC56jzX6ZyQD+SjHRBBjs/9UO/nRomBREJpAiTono4ScRBCoxNJofRE
3SwNrW6cnQG8nr5wUGLsMT+xLzJGoM23tBt1gmIikXv3nat9U+MV4J5hLeeWWcg3
Pl360zpID5Fn1fXZwU6O8/sYLEU89oftkXKohDIh9NACy4u/cSSM/tdffUCymLaG
SERjHEutziUk2qqNqGODuXDS2jxBzWNh9+eR53pE0+HGBzFHji/w2+Oo1aNknujk
HbUQOGRb8+2Inb1ZHLmil1W/ho+/VQ0gXhpMLzXHcNyQuka++OlEZbb1Av2iXUog
XiJyRQCpM5u/YcABQqt89gPos0K60zTZkg/X3SMfq/IzS+1q/Ex/WZGslMTJSKAy
X5TW3CQCJLL1um4OSX/IKprUyzd+rfUPE0tDqYYGWQlkRhgrCj6bdsN5wbACNSjF
IvQxjYMoxvRcnnJCdFhnGc73LOSEvXi4u/HR25H2ynQxl0IpPJud5oygdRyjdWEE
reDFj8sEbOkthC06o5w8uInRocDQgdnh9+eu5p7udlZlhg60+HW0K5BArin9dapd
XtqlpU8D/cAcO6zF26UGWcqIkwYeZOXCl4XyF14u24NGX1hffShtiNsSNhhoLLDE
W0bao0IjEaUw14sYIifG/UU7UTd+D7ivKNuWGhGy+S9TykDaybmCd5KnEX3+SVGj
uuPMoJbYz0e2rjxxuaVrvw6mq2Q/ysTxZ/Y7jZonvQMmPaSzqvotysEOWKc4UbbB
vektK13Ql00TlbtRrwHM3mayguFhZKr5OM0mcNCV2wHyWzzE50gS9vgeyHHVZ0kw
MXEF9ygcSqaew+DxwaT+gwU2aAmfoVDNeAnQEe8KMtV33RZvleSmIXW0KLM8wgLA
kd9/FnyYcPQ54nKzkB5DZk7JS6IOi8Ze+5Ts15Z3BYbpI8Ly3Pm/DLDaCwshxymq
K+zIxdZ1ZhTuxJhUKQFCBI9iMEcakX2k3yduqz/xGOK4DVzFlWNUFZaZHCBE/Q8P
dHIE8x80ddqWJ65eG2hqjik2ghhwb+KJWrWSsf8Fn0+t0J1qwIAG2deYl1FIkPTX
3JoA2eThdXX/6tphKjcJ5qLsFwwkMTKHRuQ7RQz7halHAh8K3QhorqRbyu6nekI2
uJWpBPYy/xD8zT/U2hsOoAxD04Z1Tb9MbuG2YF5W2xpDFAsXADOMfrKkf21yKKZI
syL1wrwhLx/MyJOy/nJ4a/uMTnG5qow4aymohutoSfzTnIoC3qgyFBsjtDQnMqvl
CiZmNn0fy9phoQ7jg8rSK2Za7dnJAd+4ysWf2Or74A+xePAZ+2HHCqqAZcW3EXxn
l/+/5FN72uI6OYPOPycuD/jEULtKu5a05A7KA3Ci165r13C37vDEXfYPNg2LILlp
k08F416Vg60uF/SJdsULBK58Hwfd96av1eU5tYtU2oYh7GQv1+jbmHEC/V+NJWlT
ZYdd1VL8asoFtPJ7KVn22ZF3sFMjJC8JySoVo4coFIJt0SW6OqX3bFx3i2nyK7T1
e4icU74fs21rniYtdZEHle+QCv2DTQqRF2YL3UgZlDQEshMATU9WULf/oB05HCH4
2NJAroO6op3CTyty1uyc0E3Vjeuc0K+y1a0xWo51FbXlfasT76+lELtSeY4o3N9u
ydGbvgLMfI+Vxji7RSSMzt+29eVZLgJ/Z/e0UljkGWDismMSyxuWgmFzAhBoceVJ
o90/lDba8Ybe1wD/lg+fq6x5vWXjP37mCwnaJ1xIxGwDOqVIM4ejFALxFB9bt81O
J3fD290Itxm2pYZbiba1DExV8BFxTHj8wOCPviScKJi115lQDPYnVeZ2J1fSMI6c
t931qgu40RDwWR60cvK8H3a/6pGJTtFHce9BIYDipSptNcb8/+oHqKE30r056AW8
w1PwqSMa/CrHv8PQ8uYZ9aiV0HEyNvbdHtZlXNWWC1x7VtBrLmimZmU6k2XN8rmr
QMiKAw0ToxAWt7Og2HUx/n27etHQjnAM8D4weJU5K4UORxCuzmef+lGcrJdUWBNY
Iw4vlsB4b2J8tQZajkqQ7jtxNxWbpi0z79byUe8as7qbfQZ8d/vFypvqosnLSXJx
J9/0LOP0/VeMmaWNJp0JFGd2Nbc6b4h7lGgDIGMkC5nQ4OitnRBoE58LembW/+Lu
Yld2CYIYQlszWBBQbv4b07NVIItmEt+Vjtfhy2BRYXHjTGHEh9rea9zxIO9apMh/
SYrPbaCe9N8SzQBp0WERweM/jmm9HJFSTJ4lgNgTssD1LhVopFSDM2MzGjnajUiI
hz58oNEjNB24Qoktr99H1AZcWmBLhJBoUyuMTeybHzuQYd527kQZlv42auUNluwl
JFIzfQf8Tnk0IAEZmEXdCF4LeyH8wksz+MYXuYifw1OLTf6bFU/AXLvKXiLy9xnZ
JkdZCacKstgKsgQY/MWkYAyrGTOTh7/KYJQ1xJjE51W8wdprLKeQtzrufqwemKUu
ub7tCmIPF4IdUuQtzeIDms+pvet1ecBRMNZtccN8a1IMIwsJsN35XiCe7uTlZDuN
A8DCC7sYGmGvgiOBg/gDAE83MbgRInARoJBxFQaNGyMYjrhAxviKoOXF31TdJLgA
hJFtzcw0/tgpkPtUerRBQ2AXgWeKQfLghU3fyy4bQ207oSBAYe4yEK0uwKetq6rw
fJoc9wCMNEPCZntJSvrI/XjDPyIBd+Lsj4U+ElIKDKURDG4sCmXBcJeZ3WQGUZId
k7vf5cubWzGNrVf1JkjnlSmJbbSQbHqDoIQme5fZ2vD2OjpdtKDRrbt1a8jvZEZO
pJXN6cwQjmS6iVM7Xb/AB9fVwNj2wmsUKxqVmwuBdMNTgq8PrYq7mttqRk7BK6f3
qQ9f6Cc+l0zkCSiSP2A/bx5ZEIohc2I2Do3NqsTRV/uusz2U53ccCvr8uaBYCwkH
oKpUmcsbm4vheBfqnCt/aQ5bBD81qi6+a0pnKYIjRzEEU9Pt4W95iyTXNT9Sj5ua
MospOa+T6VhrMkAg2kMheL/mjQpMSxvxZMqmQRyJINDn/tCPHUV/LLrZgpoLoCDY
f7I1JeZ+DVu4LW2LZaeZ0+OM4NHqq4EjNXgKGJbDYoFX8Jof0EPTSHyxLY3GdIvw
EMpi4mVQCBXp1nhMXF+4ZopmYj4igkF5CXW3QIN6Gv9Sr+sSSTrfJ5zRx6yKfE7V
gB96EA9f3AUOPrE/S24bQ8gXeomMLODU6Fs5UftnLa1xHQAeCXvT4vmdeIVOV9O/
+thTbp2g2ZJALNWRCUdYFGpMhuRci7Y4Z5iTVNFAEy3RFtC3RFlhS/zVXdiggERs
+1N/sWIyCAUnJOCXrbGtLziYag1r+efP7MljLJ8k7ZM2xfEoGL0Vg3KH9anP2obf
N0kSXe783qbmTI7xmAiqrCRZ+UDxDF22/4UBEq7ZktR+uiDGL8q/ywCVDJ+skJZv
d7JDyu7CQYTar23mNofbCfuFcKLeOThWDURHOt43kDxFDDOSpeAsdBE/DeoEAvYR
kDFV6Ju+11NbV7/IKgOx/hMCr6w8X6MIzKVTVUKBqQaNtMq+OfsBC6K3tceeJpSE
SEEho7f0jB0f0wt4BdPsFYAiAdfrq9dFe24QtfiMpQAgK3kQJfb7wtvoUJ2l/FWM
UX6FGuDdXUhT88Yg6zUAM9L3KXmxkaRR/mmr8/5Es3HlK8ngOn3QYuwy83THmeQg
RreU0n7lc5Xv8W2zKuIHGUyYWuWIIt941/iPtmcOlYxhFlDdVcenmqRqUPK4MGzu
5GOwDvFVdNws4lbo346QVY8XytewhVlLScQpopNUk9MnJqvnPsizUPK7pV7jKkMC
SFKHeuNkvBmm5y7pkr2r75PQ1txxUce/S6srXvTTRwqzMaHAnc6Zk8SQATc007IR
Zopq+d7amG41Dl/+rsjwGHWYPhznMLuIuXlnnBL64OZBQ5PnDdOKkNMgy4AnK7Xo
4wlKBLBMMHWPyxjuaYurq7i1gDtF+cTpcSKz0neMd7lXDdSEzx45z4UqaKDf2P7D
KUYUfigfRoZP8uRPFeM0ddpWwps9HaWk9DWTSSiap7qjSWU6hF1BtAlwKFiMgIF+
3K2ARmdTfPcoNsT/DvIpjFiTuC40CHo5jDJj+uOnKhQwnGm6C/NxX/lAcRqochpu
cSWoKIVLBDJVHBmfvNSt8fS/nifhKEzPnesY3D2+k0s+7nk/bZw5MQnVYr84oyRw
TRUOVCNoJBBLgu7gxnmyZ9cLe4gHRKhvB/Po+RWHVRI2tOpw0FeFxJGoUNqS19fu
d2y1XZVIMB+25pI/9p+q0Cq+b9SnD2sZD9ukp9ljOUqxAdA0j4FdCyY4+IK/usC6
SJUV0M7BPhH3JW0hUxUinwUF5tGGGPBYVy/AvJAGbDuaezjwd8sempWzuii7RhST
Uox8CYFbuliug++00/LiXRleANy58aOZzyRy7SO1y+w/u0qRaDryJ7lFNUjbdnmP
JdBf/Gi2c7FrbP5qWEqXEuoLI5VPRzIdKeU+KxaW9bMEXeA8D3zB2N4SvN/y2NA1
ykOperZ3yA+GP83QAiag4Mz39I+4w+MtRz+3gatxJyTH2YCu2ae42oRgN+ia3Qht
SbesCyqB/aZ+CLTsxZKG3iuBbIIn9m7oLfbXZuVWXr0R3iwLq/maxGwn9h2j7SpM
CUDVbmLcUvEdxyUt7yo4noDRScffyzewNqLfVfVohiXXSei7uNT/rLpbx5xnw+By
bjrKDdbzFhwvPR6E7FD7pj3Vjja7liimSGY7p1Bm4qsup8QvB3rLHkWdyAftdLgL
tGkvwL2rxb5D+JMikF66CKbmPZNd3PIZWyray5YPxXGKxSssA1eG1SlWjfzDFRjj
0jK14nGJivcHkEyY0Yn3yNCiEvwtp4TJdtI/0s4mqP/LVilpDQ2XnoS36demwOol
Nlgy3R3F65D1CzsHpJAQX34bW5e54SVC7qD3zMKbupNDyIdnh6e+awTOKQX/8kE7
Y1h67KkZerE8iKRBIUYJkKeUiQRhBeuEbmk+LaHEho8kePNVIo9QYgKKd3iNz4vT
qRzTvSZrnw5EZ4eP/XIyM0d51Y8utuSkiRumTV2eaJ7bTil/0X3COASqo+g4ZO7J
MjAfA7EVOlQD2fz9IrU1eevITFDa/6v7a9q7XIA0QXNeQ0MWdwU1mrO8lOIonQG8
m6AiBGJxSLUS1DOh/YHkkbWu5fIttuqfwddlLiL6vj2fC7ltpCOtwfYq8ZSlj5ut
Aqnd6yzs8HKxxVpHreHf1yJSOiFPUVx1WSR6EkazNJeP45aJYUS4rxVeSoTZxhmj
Ezoq5ZPXNiaqFbHjGJ0f0rZ5jk3mPtw+8KU/1MiC6+mQyA6+KTIZb3SjvZn/3IMO
IUpOop3b4LFlOODEmSNutefOT05bVo0Rnq7IffbRp4T4mHL8mSGOYSdB9Oa58thu
iw7Z5U2FGm2YbGbHu8KxEMEdwgZj3tf2r9wVWBGbdVw6OfOOeQ3xmYyF84AOZCRB
hXK1SAWWRxejXdjAntjsNZBiI4jG5SB9BnJvGOfmgojvvB3VAynYdHveEXia+ZVO
Mg5GBL+sDnYFkmW5aIGIbuvqfTWJ5PdAgtotJfa0kf+iOKiD6k1AwqqoDqQ1rzVn
Pi0huy1vIe4KWYz41jAf/AgttZiCDdnM+zpxJ++hE94Z8PS5RwRJLzQzOyZ5KEsK
cQrb19+5+nvvNHuXGSweIXnTNuz7I45P5BkPleu0ObwmPuiMpdk8KLLrHdDp2WFF
L5hpkS3VPzd9OSXF1hIWdhe+r1wqVgzBHwldu64e/RcA53DBhz52/ZeIgUC3B+H6
1uo9mHCLxfJE4IdfBby8VWKldRQREwz+nOdlskAtqKoMZY+PG5FFD1TmXeAd7d1N
351Ro/a3yvAt9ii7efWNUNkayWaYu+aP1Q+Kz+bBu9LKUUeZzY8Ti4ZHeGKkRvUE
R4c28aay6rkvboUXRPVy/jkgmnyFEaCDGXbXLY4mSu7sWa6iGltt8zSe+CZhROXO
E1kUrO2QNs3uoF+1cqkn8xfbEEhAJqFp18WdlhekBVVWSkzYiUuRZW8h8ULIPuma
ZLYpqtxf47+Qlyj1dsdkbAJPp+q+j6emn3loWNIKj5AFqUXwbKbv3zad5StPJxrN
lTdNAMMF9lYEt77CzZB1w/etKV/0CFJFH+OpMXoCwMd7HoKxek/ITUnkJE0J+2pP
pATAo9GwCfUTJhbCsxftLlhkwWHYv2zoSozeL2qSyxtBrARQT7hAx6ed/8Xp565e
Tq++ODtikDMMOZuerVuc21fe8gJHIDMcgQmc4eeOMLGfrMIpkZViwOSHKT1ya77W
VcMoknDa0lxaqyRK8Ho3I0nkpVmlQtR3yNTU2KJBS7QDJKmYl4VRlJNiwkCoT6e8
xBn7oJVg0wRu6gN1M6LiLtus3Hjr03EeZbnNeupU53eOp3TdDi7gP33FjBVcTevv
LTU/RoPF0G4GNcOAMjkTEXN0rkYU/IgTlh6p8+9fKn+2uXJe094xOa4odPJJ1eKH
A4wCRZjML/2JuUhr5YpRtB7FC+b70MOIds2XVVIj9c/hugeuA7nuQ3tunCmsOHG/
PfmMvQ8hdWFzk+/UtTWz3xZOtL3go2tc9+s/zm8UBuQPjYghqHnyy45Yh9Ac4f5z
zE1xo58xeiN90JkISvTD1KTxRVzw+mExroUWytcgHeF+GQ8keteuhBV52Kb/Oz0I
LrkZnPAjHxpachVqLyToXlbix3hwXNgL1BVEo6mxiIDiCdeZ41Zh6LO/5QU5bfvR
oxRUJZO9qHIzQqv3aCoqcKlixHOBo9usUhKsMzhqtz4N3FsjDpUrfC00SaaxIFO3
XvaNsUKfHcW9zlTd5d/q4j9yZR62mj29Zbqb4wrFgqqN++auGRf/9FyMvQtT2VMw
5gRmTh5YPz/AD259YaNRE8QBRAR7iVhf/mVs8wQOxDgaBKqldqujXBfWT1IFNzGZ
tX/Cq0aAEGALXKKNAwfZ6nlaUArN19Fm2GJSYgcVDq6VFGhoqq9haWaL+7fiv9Oh
LHzdhCH2cEDdbDUj2XickqXL/0fV12fmwr0uzCcxL6wdZIwNU7n3wA/6nQFH0Hau
h4P47AKvXX4bNC+CFYkD5ydIwGTzQvueNihSi3YRSlX2g/il2vw6eWinO4es8/SR
SgG0iF+rkZT+84XTRKrwRyopBznP8Airfp+KWOVERL3z0n9bvbuNktUaTOdAIYnJ
Nyxc0L1PllYeGSWWHlBqeNSgLim1bBZ8XkrbPKsJKH3nebzWjUC5pQrih6E16aM2
aV+hW+bC3J2gv8/Nd+ppTsg8HAlk8E8GfRq3XZWEkwvFdEUDcxSardycJgGqkUDh
zmwrjTGxzaGkhQYX5s4GdG8ZNvk9O4DQU0C9cFVL1CX8RYaFGHMd8U/aWuGxuFxl
LYS88Gy8l3Cv9m8TA84LGCDHfyGKGwjzxyRjy4ZSh5BHw9kwA5BiQj4lIqSjQzNi
7Hiwe0aMW2BpuhCZq+ONtD/wXBJz6UNA/EwnSBc3vW6sSl6ljjyOwZs+iSw9aw7i
FqYgTIK+/d5m2N8vTBf61kzedBStsyjyXh2RL2fswvJG03m9v9m3G3sEuoNeiTRh
/UoQhZbFeUZYIZBfOcoU4zO2pc5TLu7knHOjHBQDK+rhuLr3+URGC1A0/n8oQm55
8dVFFfMt3i9sy41O64Sex3ULFs7qzspIUDMUUTO0NcnAQ3eDGs/jvgGzcU1g53YM
94VUxSGhq3bxFFr5cKCudX3VQJDr67lrMGU03tnS2MK/GT5rYCxQnWMb+qs0RhhW
Ai0Qe5oLpej76bC//AxTe2CjHQIHD+aWZpVGb42O/BjLacOTJguXHBuUThiGWEmB
1NlaQalw1rXvLgeZWqFE24Y/5hu4jDTN44WNryzox2PLacwqUZoHGaUu1zoa9RgK
Oc8snV60ZJf+ddAEAcUuf4WJFezxm3OcguxBGHuUruGUdMq8O9kuDfsuGgFNYCyx
j2+pNii/n0uWXOBoluZKvmRn8PAHEEmgIOvWcAN+Wm0io2eYLx33OwYKTbWa2eGb
JdJwFz3TJBvrqrvj+ijiRTbOff2kPa0js0w1xsj9UHrhHWF8+/JiwcewVwj22xO0
oFnJ5guNYmeOFO0B6tpF3476GjhpWvp9Z01DSpNYOu+w3w9NAvEiPDR25ft+d7pO
Op/klrYbgXTYSeVR8MXIZGmphENd2AuBQ9zLfLBbJP6FsgfNRKjc7VV5uLX1E6cD
pCpqObK8NaJJgTHnTjDRLpXn7WJkMTetTpl1xW4rqTo+d0lLM7LmddYEdrXnPvjJ
ftzD7PbD4fG4vP/EFN3QGG83wmFcAM70qF6HN0dK89MxdzxRkDZZOeTmRoYjPXFR
MHCOEuunkbABwlcudNfGwsFeAftZk/VBsppvs+4oaIWj1xQWKWwKPkvK5Vfrzq3I
HJ//SRDhVFt91wZmAe6jV47vWmBsJnNOlRp1HIPah6s9YVCSC2Pudy7x9FtvDRhB
eDK4W2N7kM+dE3X82XZOgTFchjS0L6pKaopY5CTAEGG8Kn+nsoSuktp+tDgkrDuw
wcBYBhIleh8uhcakI00wD6UcUpMhTpi0F7yrthC/xzhW2Dxhgd36oU7A2CbNChhn
2S3DC7zIcV8JDU8JX0zYK98gM9d2OlHDyaOo9FfPisw7UTWqmchA0dP1QdveVRyb
zD7TE0jCLjY7cKaIls/NSE+N1wCr78WjXwJ/+pSAVwgCbJ2vdzWe0oNJ0PuP+2Ra
kIGO+0cAJICLbOsB+eCA2P+me7ss9KYP753RFOd4aKxLIaRsCpdool+I1WQXBxEw
R4vQyA+hxB6xCBTvF+Ag1lJrzTS2cfUsD6beulIxHaX+jD2DPhsT7SccSeRFQ3qn
ptHWXflbOJvFr6eD3sJB9pCYlvEDdImQ/IlMHErovyAlcjtGFjDJCtbh7zEAlw/0
J6Ujnbfl8jvKRsHKU2/lSAkMxJTXZ1itcfwt6Ez3vKAMhyAdKfd4bvsZG9DVGhDE
DST1cEjlahzw9EAPObTAB9BABN9iAPq7IbqhKhLt0fW9ItiZix5EmpBOLPfto4Sg
mGNPyPqHHNOhgZIQ3VMocde4fvCxKkjpl9WY2ayCouLlFemnQtb2TxOBhQWLrfI8
o/VE2PTGy7SSFhCIU4D0OpHSNYJOBH2BLbxlHN2VZcRzVKX3iQeB8Fekq/UjcGgD
OOLxxFeeq1oF9mCc0y+fdOLZGvpEkCKvRAOxTiNAVA7/PrzFYDvYybjIE2MTk5Ag
W2CBXNryZ0CezdPXMaUjJRajwkUDUM0E2rIywwBx15At5RB+6UQZYj3MCh4QCEuW
GLlIJelFTloqPoxdPKrMM+Ld/yZEbzlW217eaqdiMZmI4GkIIOR1n/9kssKbKN3X
0p68lNpTPkiTVTmV9jTCEAwfjBHpq8J84RtBx7FrIQo+GeM12SAhlRnJNcZVKRJ4
MA4Xj0P8Xb7n+fJAYEqRDD4pc9/ecmWIqWqwZp99DP9rLG372wVJMU8SdPW3pfPU
ij5cyfUWLtVHyoIh+9xTfRovtlTihLF3Wu5vjY0qMQ4Kb3HOCOWQEFhG6zBLR1Uv
LKdtbLwSp0S6p/tOouItWgayZO36PYkzzj4Sg/wmRwO8Mf3BcGk1QeNrVIvPNbd2
z1QpJNX0gFgb6oFhbZGytEJdL7Ws9oDLfyDLikigGc2NDKb34Dei+dNZQOEZdHJ+
Uta5GjmbQ+VZShT/aclDdtv+lZAAckJqcJMLQDWUQSZpTQHF56/Bi3dUH3zEqgO1
3dmRyWBBgy8KdewF44YqViaJA8A3Z3h6VWNF/oJqCPTrP2LR8UpzMlwVYBZlyOvc
I5dvI8f8EIYySYnGzrDt+92MTGVJH8umq9m75MsVauVAFi+suWJcjkPqQjWEZK+Q
sIyakgySBnplZwqjH26V+9yC790LqtTDUXE4ChL9a0BGo9s64BEZtywbVK7b9O5x
5I/wP6vW0fCE61uKnagiIznl0dJ3BzCVr+v6bLiJqm16LqVXqo5E9yyM4Kp3k5WR
p3f9EsiX8dEpdS/u1zb2e+AZ914cQxAF/zgkcR3jbZfxVT0es9LJ2VdFx4SrvdY8
8lLMnwc6pdra9ml4WSgbDTI1X5mvCKd+jcn3IItuiRH3GzAVX6yl9qjxtVCqNji1
QUr1elLgYkHFLDJjg/OlukwWYnN3t5heHgVLWUWByFMr7NGk15YzviFS+GTCY1Uj
K/BfPjJ/SLuRHgD8sZr00wAs57mabYHIq5mf7FEz897KEdU6Nh3zDj4nEogWUjl3
P0J8SjAx9xlVJr7jXKuYCFuyDRHw3HiBNTG0T+cPS+gPYTwqn2e6xO12u8SubMo5
AVxydLPr3wRAvf5V08L93LBMYk0Pg6mkiq65HBHStK3Te/53/zfjY1oqCf+VcpM8
JQRbv+aRzRSTXeOD7EnZa9ZNoArmmdz4Ry1KsLOmCU6QoRti+w7Bl+Xriy/6fE7x
fS25tAGLNUgVJaI6BnWT4LnzKtKColXBY2eoGhJni1BhZONd62IvDUYxpYe+5pWW
60AnDhyweuoXwNx4h3H5i/s3xJ8iwky3//rFK2IXyL1QuchuQCM1TzubaSeIUK5H
uFVjn6z4t+tX/1UmLUxylvBvNYrgZbwFPMdJ02guKmz8zexh4ZK7kRA/jS2/1fIA
PF3UXsxxcAnA4uK2VC7+jxALysPflQ1XKkRk4nfbge63kbWdBm93vhuMRar8pLo6
k/VLtT1QhfXGmiEA2ABOH+iz37vDHsjvY/lS33QOmXBgR6qjkXyEmN7XtC0l36od
o1vAp9K2WLBVPDYsLsIFn6vScJcOk3dUFYqkP98C9uLNIEbD1L9FPFrw8+ELzuHG
ZmnGwUkVTSN95S4FXN8b6W15FWudjlkyBFG0DVXR8ObLqc7dkOBDUWVZH8AmnAq7
zwD/IxWmGwjRsRD8+k11Spa4wwNIN0tg7lzm0sMDEZkBy0VgKrzqsCx/icHRJK+v
OEhxf28X5yH2iUwLWRahhmSmL+MBSmj3J+2O3HbMW0PFX3SIiGmAjV4OweCklG+s
b4ru7FjezOQ06HuQ5Vs1qgTYNzKWBpshGZHANmTB8EWHvJc1eLUbjUDqmfYRm5Mx
GV2ELNG7b+C0GyZAawiV8sB9W8Fc6fNKGdd68WHijiauMdqpF2CjTpKHeMxQ9yay
V6SEUsNdr0hLnlBZfyJM9BH6Vov/v6Dq2aGHK6bNXvaIXQ6ucbaQj3AWD6n93z9/
t5oGe3Skg1rRYDqRm8Z/Qiwu/C5EtSAwwJT4oWw3xFmuo6mWwVzfI8yPua/rwZmD
MVWAcedjzi/bdQ4lDaoz5JEYu0XO262m3R52YMb+D076HK5BzlqCzMQIPODbsFAI
YYjc+A8GAhp/F4kS/yN2lYX/CssDXcYIzU1dfQzPZ+P9RntciDnFEUHzwK/hFDTH
m86+Jjuj4XIgf7lvnwIZlw8NmptnpQLf9XwiO2nGJOusvELsBIEME1VqiKVm5XON
YTIqa1WjVD1cVWZNgaAll2f+SYJ0JDEvTkPDaLpIrlLyKuazepUgNofaB5EUhWuj
atvTrQAZpF56wX7aYxuciXfPmOEzV88uUPkXSpnWtmxoaCHEfIo+f3D2ymME0uSm
nIzTl0LWvv9mBzsSAPRcJtNFS0ODVzYjLtp5v6o5Jb1D2A2cyg1/WWWu88rLzxjr
SksGSV9yvgWgJlMqmnqhwPjycg/UjTo7X5wzT++oF3e0M4XD9yEt8L6f5X1VUY4Y
GA1zKPPY/usxhc3lfzLOQECeGkRhjdWIJsuJSs94dJlfC7NmSWLLCgrSbilwIXNb
pHGPWK7OQHS6quN04xhrlPJVhMjlXyWbAp/vpwKLwnYETKD40zUOl3OBOFJOZp+E
7TnUF8ezY/m/jALSZT3YWYYBQc8TZKK2OzRTjpwtrqLcMZzEEG1tUh2pfC7D505z
friCYdKhpQkGmc53Dxzqq5l4gnRmJqKGG2S6MncsjB/vYaVAmV6dVR63QWp0FM7m
uxwQsVq7szvS73+HbQpAhf7qqDZmFfnTAJqkkuUbR8AVi4bv/eqwz0ovl8/eZfpd
89xeXTOweCDlgJpu0rGq9ETr8fOPkQhYhm6FARoD2VF9SM8Sc6uWgig3DKIjEroS
rsjr54nGSQt6ooRJwgh1o81U7vy/lhk5HXHlMLRAso2OLlFo4p+B7QnkGu8k4EeT
6yhdPdEXNFGFqDD6+IJg5EaVy0OQ4q/WUTQ0Lh48mxoI7MnE6+Z48eQVPWjLhqBO
8E8TxYJYGL+ayyC1bgxpDMLKRVhl5Tl+MclaWKRHoFrIO4CJOHJRGn/BDnSEuY0j
Euc19AUEUeB4yStdFCUV9aHbOK26RO8DhHfl9JJv6TbvdrLqC0cWwesGpcWK0pif
zUrIldLfZ3Qqw8Fp6X3Mptf49csTXnW64aT7hgM+D6vvldB9aQKhBdUn+OW8kMoZ
9m+MX10S82i7ulICFkEHtwDAGTn5E61LmmfA9A+TXigxsUlsmBWFp4NF9dVAk8G8
Wcuno6sbAy8FXpPjjwH5KBorxVoom9hdDI9cA1gGI3EMx+pYAuiDb5rxxfJ4rN77
PjOjAvdUATRmYQHlifrfKTDwnzL+hWOs/yi26G+nU0GEtDKp/6HwMQvzR/s0LFms
4/EIpJzNbzGYO35XfsLuv/2R4Dq/LxIPMjZUoxlRuKShOWa4wsuUXk9ODWOmqSf0
w4MDhslXGmsNELIA6k8lOsoGq3tBx4P0Q+sXPEUG882btVfZmcWYk01ut+4al3bM
KUFNychpR4yUYjGvBeSEUkNnulTeHQ0No2ugAWryE/W88Iliamnh3elpBhfGprxj
56zgWXohtLG0KzPI008Nkzw2JWYe2Fo5eal6cerNtV1DYe7g83FChUVe2/GYvgYz
JEvs6FsB6K9t91frFGCM+8yxt5ZbvkkF28aPX+wLe6HGotJTU9JZBUTK5HCnR7wp
TLpQK2rvklE7xd5gP6wss5EWY4iDyr4u7DDnCmDwwUsuQR+VJsipXiSGJP2dOhHz
BucmxSXRPRI0J2Ey8iNiukFc2SNDqKt98t5KYzS1zj+cMZS4uTNH4OwCm7KiBYue
ch9mT7lzYVN0Uvz3iemC93Zxcsk43nU46qZUkdKpXhlJ/9POj9EtWo30UDDL2+cA
Z4ZKyQyl8+EvekA8qr7o32E1aFbynlNi/r1uDFTu16xuubUTZuaF7WzcUc3j/GBE
OfimIYINtN9xtfhzeCDVzJF/trYjXCR7N2bW3xC7+JDlD4598p8sxsfU14mseDEt
TyecNtk69J/9b+pYcWJaG1kJEaQpjWX5RWKozw1CUoyNEJT3yrQMOr3WZyYCZ31R
7C1JK9wM3Ku2mo6hVddUAZ6arXmDPWz3pHyLnlc6ayPi+y8aadPVHjjC1q85MI7q
xFliJCcxU5kQtYk7q/TzLLcxIRRif2Is69NZoftDqT+o2dVhWeAbhbl3nAw505mD
SJflqwrIRFyPfsaVxwiHvyMp2kxYeG4LfsMoU/G4ae7Z6iQtrQY7p5o0bS5MWO6D
rnleGMUfcb1CES64CAnGKOvWZ3w9TvIaWF2tAlAyrzAqjzqG77dUXIhOVlEkrpuH
wQ5CbEufQ2syTXgKD/PqEzRZop0CROfBZaTl2lFktKYi8raEtf5mHrypufPOzEmV
Ug64arBTSbZZ0nDOqSXABMUPjdQob46Ip3Id2MIWvKJFr/Q4I6cgwrZ7dSKG/kn8
hTXne97VfPESd00MPzYtphdD9Zc+/pWqVc2HKXFlA/FrAHi9Hui66mLIq0PjV0Mj
n2dqSy7xWgrOb9UfWTAP3rdcDGA8dD0+iphpLor+8FdstfDkiPP3XyBeMWNdPqld
vspll1xBqZSVVEG7c2QhrCSxLJ5W1J0RXoUvDDQXtDxnUzpjGykZXhTXoa1g8cpY
l+2/2MzCL+s6xxfQvGxkJ1vxtLe7uKjk8Dlx6QSC2L92WJf6r79mE6/vyuLbnTrO
rItTZWSqtySo8DhBt+NGAeYY5vtrlgCknUgKtvpd8Cg/yH7rKrrY4mPKsecUJUZF
BhXpmaVZOJHwGQCW5XtqZELYXLh+hPQV6UhNxidpS9DQpkoCwd5aLzuxnYzELCAm
uRh8FmRlw3uCKFq1+H9TwMZX8nTc8v4l2p4rhwUB+PeZbFbKt/FRGQX4WSL3m9fB
/d/rt7Pf/Cwzde4Mn3hHKnokwtrGKWxzC1FdbW8xy/JluSBt/oW9LYyhYM3DBqgC
2nu5VqEAcDlWaIKNX4W6KtHIcDe9Mha7KZCvue+wmkEujg2w71QsfYX4O9ckM999
79+bsz6cblNvz+qnMNxr0ymq6nCuXbakHsxflHec2SuE6KEtGNL1LRJK6rvnEaKh
+WiXV1Q4i3JHudOCwbX693gDE6E3+bICQV4td2ayU8ipO99h0m/x3jcgcTTmaEaa
0Gs4miopP55ygXJ3kd5l3GaG/tnxweoBrZJi0MV3VJSIP33StUBoWGHVLDfJZIJ9
2pRcJ5vH9LbvbxpdUYyDN7yKo/UfkVmrGawls1v3nftEbL3ynaLHJ3tS0muTAt/L
wFDyR/jU0LrJoqRyMMi72gO57nbZP7UqfPuETT3hbchCuVUe3K9fVKU2aIBwqVoK
4Nqc5C28sy0ztDsru/7gxLjEI4kxEffUD6n3eYwJzXryCmwglcdu5YPrH53CLy0z
PxkFwWD0Qgifs2KZs1qNDX3nBYD3l0XdKy5cHi9wcT1h3dH/xBjzM8IzYYu/ndk7
lQUDV/WmlsCgVZKFY8al5euodnyQaoKOLtm4l0R6VsZVHGxWmPfBNVkYc9qCdTmx
PWwurHG94Ci2DH/AqvlPiuaF5YBB47RTXH/lhj0litsZeGtMgMT1qocw4mivVyJl
3OU//Srmiz+KpG89afH2MIJhdeEoX6Z2kkQFlOLicFvuJ+epRqvoa5KRPhEGXL/u
bVY30LHEjVhys2H61i9o48d0TtclxbD6BM3D/E00nBa8RTYOKRp7tPRV5XzEK+4t
Sa5oRBB32wIyYtKX1+u5vyKXNjAr0ecxVeMFF56AEEeyRPQZ4otNtSe5cD6+ftSu
t9QF/ttvyvOjEgWa3OBmZw1MRKiUCLS3Q6jh0lApqRsQRTJ7lcYzoJHI2Hb016Xt
5Dpl4c4EO57Os11ABqSi7dTCohtb9mz6xz2/4wKcdwyO1BiOpvExR5J7EFK/VWwL
gexXr0VVRt5LjA7+ThEX62oKeFYXX5fq6H7cqi2y4xGV2CWuTEiS89laN4PHDQUn
GcUfAtmzo+Fr/jfU6py4qgTRwCa5pm4f+fEBMXtL2w3YI+Kzl/OUyZtFNfNo7h1+
VGLXgZlut6n+Zcgt4Av8ghh609m2LxCo4MV9+uJfdZ5fQ+5z3isRQvzYvTKOyGeT
Tp7k82R6OdrBSwHSxolXy2QyLii0jXZ8t9eycL+LEjxPPx+ssGSkrNY0U282SyDq
uwRrJGmCDTAPUqyhkoyIXvRCpuKsKR2uyehMBGMSCBgAETVouXsgQQ7L+3rh3Km8
jwoXEXj61ROqb96AqYImhytvq5HchnUd7+0NVz3kjeuep/KAPe+0ySpvSGmxomfZ
oa3yE6TSa+TyMs2Y+IWvObp15KaVG45K4mNmu3wwOZ8DNh9DMX+AvhehWTDHt32J
3/5kOM6Had59gD3qSRXhI2vg1abg3rGxlMQqQ/74hayZOl9bM+pQOahxBLvqFwrV
G+GGvqs0abkzz3BMoREzyihadlXCTVM2jKL0h9Gu4Dmos2YOfHgs9BuktPjcvCDG
UKiHF1owWZH79Chyfy1geTE9bSGMLnOYF3MdPwWgT4fzF+WJoQKNYhyL7+T0mFye
NsgPPqHwoawu7dclEpxRYCB7D8wfTq2OFPcfcEmOU49HRQCNvmJuBgSfh1FNpOb8
0ZdO8pUUed69sx/n3vRpTXX3m//8fMJ3kpf62e5TFpMtToQBYLXH7o5LoDl+32Y4
x9hIvVKpOznRu+3HBQYP+MsCRdRGvcQ3s1BRidOgg7oukMdb53nUes9Bu8SNAOwl
U9Gnsc3szJp7lYop6eH2AVkvffE9YWfH++R3cnl/dcJW60GVjp7Xtnd/+erUB/19
kUyJiQLqOa5lGdHdQMLp8d1rR+tw3GRT1Cok4ma8SNE6dornWVTlKh2kgMkUFOnk
bCq//aF+Mm8hjD7SIUWSg61i87LTGs4ZymAOAveLFeV6tFruIhGFljEbc07I5cQU
y59R/q2hs2yr8R9XkKfCJlnMfmbqDrAs/EJkciaPvYa3lrOJNcU31kud/ctHCacP
n52ljF/pHsqMQjOzPKMHXIMQxxw1R7yq3qNNt1qrQg/kMT7E9vjtVxgz7+pdpCvC
o5JR8wCFguQBalTQzDspfy5Lraqc5xGDCcgoVAyPqCUXt9UPVDKKj8diyUeh9BnE
5r4XA4+kwwo2MIUkcLZQ11vl40nGa/WOMIr9bry1k9YW8NHod7p5g95IadxtVa83
0He8JKO6dZ2Obu9taEe+UiOEWAJ+nIcIyRgO35DgpYmZcl2Nf/2WATwDyIilPQ+d
rSVRVCAPwd0vS3fsnojjyqKBNxJKt3eGJhJ7kUhEPHlpMumxhE7xEtSCc0EJmCK5
4UJBx6+CiK20fpl4C8aFgZlwzERU8SD762lN86v3/0fdfHh3bbPaK7gfnmLFkBEb
+2J+hao5mjHGB9yu0XO/z4rgGx4bkM5iuncPrHtW6vqd75lAHj1+Ph7+bdLlzqCE
8Lc/yxr6rZVaGKKBq4WrgoMERJJ+7HS4fNuf47hdtAb820te8O1BDLojTGzxOjXX
97dhCLElpLgmtvP3IOztBMfsfcs4Cf8RgjvBuPk0BRTreSDmBTPKNs53RtBrrL5+
1OCycG9U/hnCR8afUXVxjammVWiCDqmJK5uKrepNjKUq372hWq4yTaUBaOQlZGpQ
spbFc1VTLqzEqrAeEjvX2C/aCqsoPOkwRdQkEezePcMdnmwo8kRVOP/q0jcyp98Q
SzM+/YJDCh16dgYfDUaV+auSrIlArbBeVWOrZHe+i/SM3Sl/xBAGpOlNpUOws5m4
z0RWPT03n3CY4hFMtqGAJ8CE8UraAFMjc4eRHcu0BHgIDwhjRyV0VbqxrcPD1MqI
PS1r4Wngc4JcQQNTN7MGMqUtsddL576DBEFskgOiS3PkSYrePPkpT7nqPWc+KpuP
/QtKDRyotnbvFqWG3rAI0zKAAFZss3VBijILsiWOMKlIA4NPx6L37iAK+KM2fYDE
iy+YhJqU7VY/76+rmkZXbPFxhIpTCuQDNnvUbXB7eusez5KbYBvnofE0hfCQK1JO
dglMD05FJlPZAyTu2MNnJ+Osev6DX3Pg9/tZhrs4LIVOOygAF6DMq18INs2w13ZX
xHtyvbNvlRB3pB3B9jL7WOO19yf3CfK5gp38CeR+bNLD4kE36V66eFXPFakjosZt
t7NiebFD2Oq0ujYm9BrySrtq4Hw4D+WTunctMNl7e+sqp+YiUZSOU6ix8exbKA1Q
MEgv1mcHAPD0uD6JfBRIpIiwwGTr1Sy1A009Uv99vDbrPrhlZTtIRtxcjcQIAQn1
DPqtdOUoqDUF1oid3h17WlaBEHgSK5nM5lZsloVe9fM1XqPT1t+dill2pROEHVRN
IaZ8kIsBHoA0PQ/vboFFP5wR1Fu52lTxccXt7ol9fpNPTiDIVsD0wpa6CE0kp580
q+nHP/dU5pdrc70Fo5a9FKbhcrJMf5xpP4EmS2Ei6l1Sz2wnoLmrikDNxVSC6ZuS
LWGifH8y0rkKeqUIgLID7G5606KgY5DJyJfeWFNfy02UXfwb5ARS9JMwzovnR847
JbFUokIRLV9qDuDbKO46x7Ka0oCLzfBe58e86SpTop2HSjqcbxEE7ZAKELeWHBNm
YwhWWa0K0rlVma1J4xxAUh8FUFpj9DQSpvwx8JC0UiVGcasghLy5YDADOHpcwgym
WTF5/E40WvEKsP3MS1gZcSXUHVxQpjFRX8srj1oXC61IvvyBjKa5tnxHK7bLL2fw
64TX6WugDPQF+7vxCtj4dktKTb/D8c/s3BD8ThXcox6Z0ENSS1UG/aadQK9mPsLc
Ty+AH6FCWnl2UNmy86z7heC5Wer09wpdma09v0sXSsLkBC/ANKJ3iMYdHF5bSl1b
q5x/PViJybyAisHzQYVBcpeI+3ux7dfM/HoOamGOl9llJFewvpy9hmz1LoE40d6N
15rhoaMcjdRurMK9EIgyucsc+0Jc/mFidRPe9x3Q/gBjIgmh4Xk6tHEDlBng1MQD
BNTND2+EAUO5OcnTVFlSo1/f3a3ldNMYuQNVdkeQ9F4jF0N3V/semkdK1ZJxWpEA
fQPsFJIyDcekt/kif+hbftROSxzG15jUWj0tfuts68zFCVGGPL8zNX9DMMLuTzBU
UlTDK5lhuBb6Wj5CGgx1q5ivioKmIvqnHgsQjVffw0maLbBZSHTFkcstXd2sECiG
e1Gq62MeIIRr6bm+CEhHSlV8hWWUyfcLc7KmpsR6bbOD1CVnNxNv7GCSJItAQOoy
SjQEXX2F1WYYm90bkY2tt6y3rQP57lNNXkyDTmU3Tf01fZuF/agGJx4jRsLtgD3L
X+drHHWf1LysQMuEtyvJ9pjaXqDwpTnbDJ4A2XQ2qLf5vFRUwrLUnr1Z8vq/IV5G
WMS8ilx9tPt94vosNrQNn+ne3ta9mk0GURBdRlt99BT9Z9oGVTjNVubL8g5xgQyH
BGdB/Tz0CDlkkoXFAhNqShA/M3sIoYIcvxUZNBSZ6G4AAug+jbO6kdEK01O//5Js
B3y38TZ9DymPnBsKOZ2ehvc0lpAvxyP8d+S/1otf+QpQiiTJrGlgJXlMlT/t00w0
PzBMOZBzEuSh4SyVBzYjqsPEXOKFJDIhZb3x/2c85oNBnYKLCK1dVsEWE7qZm/gP
oglk9dUqFw4gYOWgn8JKVwX0HGjaVa/QbTJgEGuVw3Pg1WpBkg3eauTiLECZgJ7y
BUh71AoRZ8HgT/UWaSgFN/7VG0VEQ6grORh4wBeGGKc8SFSEgX9Fp9chxyrxMHWO
DZxm2CUMeL3mT3O0QmY296ZEvrqfUqQs0EyUy1HonGkKILe1r9uNbX1f7JLzRQEh
JCHE2c4xFqxPJHwwOgSupw4OkTHNlHrJ7WHBZlo5m0vkJZfeHwsi61ecHuRO8YYd
TngGDen2H23UMfz6aKWt9IlcKl7oN5MYg+HvDaE9dkvJ0198h9Kx/b4eAS5bd72R
3+SNK1kSIjnJSXdZFULlipPwJLnXmuETVNN1jJlnDTLHMNWZpXtlRDM9zmh62rxE
S4IW5hox0WpaQzvRRf0viT5gmBH4RG8n4f9N1X6rcCmjnphhSuE+NdOWPGlhFFQ5
A8cT7MW7ifDk1wczvBk/doM2/9fDepOZ8qjzXfMAv88Ql5GbBTGGdrB7IZbEzSFk
Lc2GRadm9YXIuCa4lZ5NGhAr/08R0n8woRl5IxIUJJ+x+zXl7nwdIB4vPxwiqgND
xuxPSIBY/jdFzd59Q9fcSxqXm8f26tQIEirecYaszQ6+CVT3Ok9Zls9GAsQqLvCA
6XrfyT4jM7keqecee1mULTaNNP5Tkp3RKHNopODlVEpbnwfmvxlA7IjOEdhRP/P/
y4+9S5w2jCRLvUPcuTO2MI8FyIXhXGmmBYi4wvQAKG1LvEijvJeSWlmquXvDUBiP
jDhsMQfLuF4ehT2HiG0o3q6bln+8liHQtumbkGlgEuzfPPx+ts4Rza3V6025mL81
9C4J21uN/8mJ8ec8UZ/pMzMrpBUiuoicAEj710GFeR9NSm0kputkp3pFmwzivo6y
sqiW/w476j4lAM+FHU0hvJpk8ArlpZGYvYKdTTVMumNUezjh6OZ3z+mMN9+cA5sy
/QWab1v6tPdOrgGSAs/QGLlze+sQSiZUB8MZ7bRo8Cd8EwxWmUcrJyD8hmJM5xmc
ULeXc1zO4roVdwokzYgaNJ5n0KeoXgO14ytJo3jMMJYOaxdHw8pCZNjZILmq3Nis
W3gafA9/tcOR3JUHZHhG3OBOolK2Ns92hD4lka1eiIv0/+CrZXdSx49/pjmcT9/g
H/Oy2Y/0WhjPBJPZU7fkjHL1nR49y0F7bbltwouc3a0A7fR4apL3FKcvRrt5dJGs
iJNEIRkFNkUcW9HvV3e9IFF8QgDGAspOXp1tIAOlCBOPJSPXHEKVmIyf+ur87lUD
uO0BsfuqUz9f5QwvwV8iceCrmsnXE2QtWHDJywxmwLaNXDbfUErLAMvFi6pK5YXT
WJJwPCMpxa8TFJMDTwhADot+Iss2OhpKacbdtg5tHRtXEW9LXw1YwDd0fuFRG+Ck
qk/yvGZJ96oFP+Km4X8ZAwG6WzXvrCZraXMeEOMYxs0gCGwz+AtxcWQqlstpoQO0
Zc8g73V76ekXbmyLumqfqXcMjTY6N7hUfKavxrEcg5b2a5OxF2yHnW/sYZNDnX1t
XdJc8YGbxn8ygxo1kAUKTe8b1PpLa+/Sn28hRc1514wVchiieQXKwYvF+BHcdN5A
G4zICT0o2xko6jKlHmRzvhRrfdWv2lj/w8VWuCuWs66QPxJdV9q47PIq4lVrfYdF
hyMZ3G1zyIxonIvrE5ZFNd4zELBGxfCqjcSvEr3mS5dNslYakIpxiiLOy03Pu9nm
i8+QZyFusosIkBNT+nMYlEyauKXcnoPtvakau10I5cq7HDiIfBbRp8YYirro8NUW
P611AbznGLplsdk+3i7LTrGvT4OI6OH5D9upKHjqeNtzo3DCjiMj0hR1b8ZAIgwp
mabhIhjeJ7Iypl3Z06r8NtuVfrmpHZZ6QRMvEhbxLE2aCbJ4sxs8mUJaatFA7Vqt
UH0VSXXERfwqY3lxcFAaZlK43NIuXsD6Ar32e8W+52T6EkCb4yaAwOfD47U/tJ8J
pv0uG/ZKWBdHrOMm15eej3WJnjopIR0pYOv8gWWsFN28NzBYW+va4PeZ0VnO2Ffp
ZkFJrGCgls9Q370PE2GXToSIr2djc3icDTSgHtx2NPWRbB9GQWQW2wQnxsBicQsA
OR2PLc3Gg3WlTrQCP7l0r963p17JPusQ3CBJ2d38Tx6KCuBXwV15keQnPn4fc+x7
snQv/9ZFLRPjJ6fREZ+7bqPeYN8vullf8KVImkWmAJD2zwE6cZF/iRnxeXYa0TGL
uwmaLSknL05ZdjVAbpODXIDz4Ah20t9s8dte+pEtW0pN1otxfzE3dL+qf8Mk7FF4
ciKSVHhbbllrSCYWLJmF0PuDGJVdnjQaQlu8VvU2tobRm0hWEQ1rLXlZYf61W28f
TITxKU/nFu5bhf7UbMTMF/jjUgAJfe3qNcig4tB6UqGMPJht+FJOIXsJKoYZkGxO
Ep0tAJK4vhtem1rEVdwzHupTVzWpphv2EttWOC54rRsBtHbIvBH0OE+N8mHXLlNH
IsgaXoE2FCRIsagFryC90x2mT79A1eLY0UhuCFU4l0iILjXwnqkMUNTgnbKQ9F4l
0sWgsNcqvWTpCbC406rxJYvqG6y/ENSFvmzqNqHNtMdGgcVYhIQjC5UqZFbOJM79
5R9jpRO8ZxbG3kVXCtoBK7pjWXUi0YQBzLJEY3pK77gga8KxtwLSBowrswWZoHuG
N4lo5x8K+qmu6tkutL2ZeMzStOpHNwjcycHkvW6NgYTiAsKGOcY06tQZQ0/4ki6V
8eOHy82B9WhN71GhG0BXBiqq/NnRc6lcjIK+A4qTn+oVf6ZexrPluJMhxAvwnIPr
VNnq8f6WPcfHZQjcEAC6YDnDs6vyEZHeHn7SNDvL9BYzFPahOlXaOBv4srOx+Vtb
aRDUsHLERsLQmT2DIUpItDDVIztU/aM7eBMAgBS7wLC9wKT9A2AWL9dEunJk97nC
tZtXMJ7hzaAg9MZPNc11JW5aN0yfD83TCzSMdS/9S6slKZBIANbx7aTm7OxIkGmL
Qkmg+TpwcoC/wx6/cjHobypmy6+BCRJHszhaeoxOGaGVy3pyGYUTrGOBhRK1DCOO
0x9seWyxl6QVBkXcow4yR4jwB9jZ4Q13/6rgfH8tBs/ETpBlFq6rnalTk2Sk2kiV
Hqm3aS0aKdntmxrUJI6sHdSxC/EFlC1c0W22UOcWnrDe6K3qr2kVNFdY1x8FWzHL
e759NmO/jG2Rfdjrp7zSAoNapgdDVdVQE4fC8C9zQL5bljqfA84j817SRuaVUtAe
+LKR+hfTrHLiTqM7vbVljRS/e95GHTJM+Zqivm6S9vfaU9T+hiMGsna1nfFj8a1l
Z7xC3FsjVwQHnx6oN/YHpILLUEgTK36aQALpvRJzl6+YGuC/DpGLTOY+gBFsMcoj
M3woABulzg0ln7trLE2UobVa7BSTWOvAOZBN3C3iUC9hadT0+eBHwt0ClsFnATHy
H8mn6Z3B3XTK8SdNH+nbKRTw/e1ri/hB7RVDhONxdLD6inkQcN41jhgY6cSW2/ZA
rO07t1xq+lGwVaI6t+uC9OP8bYPHpDHl4tHEgqd4dCB+fqF/SvMv2SYGg+ommpPi
lX8E0b+PigIqwGdSO7u6RMDDMxprvDhYTYvNk1rA0/Fp3KEdpRKUYA8Tw2rjLohT
BBcBmkj5nwj9HWqxTZS91cDk+eaO2gZnEv3fn/hWuprFvvA8/JuRFGER3AFBL3p4
hznZCri8ARHiEmYGiYxiiGVoMHqI0B85ROi5Dk75Yn4t86GQu0tlSQFAwt9fh18B
MwGGcjpdapr7XHxFfAAEz6lhVdpIx4kTPq9b2piKAwrMstKz1C1NXOuvX04PpxRT
rrxbDuer4SrO+bsPQXguTfht7ptRsHrUe3T0ntusktnDMp51DBng18IVKJ55rX8j
yjWuqkKqoxLjzy+eHTjJspmj6wVXK20gYyZToJIMCDGxUmVkKpea5NzGtv1Oku1W
dZJgRMTBEeslf3USMQ6L5TKi5gfmLglkuBqSJEmfUzu2m/ezdaMW2/+yLktrOnqT
dBpLG0t1ZcLvB2YU5UVsmUC4WZ8dwlVUkMZ6nS07gg302UzKOvCl/6dk37IkWiM9
eJS2OjqTFDaOly7FydStpIzXVE3wrhIUAgSMXYR2Qk0mtv73bXeEmddWkrwYfyKv
F7bIC/rdAsztQ2QfgMwg3/3rnhWRJp0CDrbnBxhhq/fopcOGO/YoPAPvjQ9KtV1V
URxvyWl0K01Ezn4dKwo8Vc36P4J5v/hWZGbeOATPVnS057bEAlicryK8HOCP9MC9
xyiZOFIECwSSS3RpladcpNwl7rTQbK+9b+A9MV69K1WJ3gaQllKLqPnLUPkm/f7N
Ea7daAlrGP5h6rQGuJl2uD4rnIhSz88oJhD86fRuQTWpxLo0c3cPTI4Ao906mwi+
PJ0dJGx4GLI/Z9XhqRkyZ6Drqd9iSBYEr1ROU7agLuj5nILod0kIenoc1ynxYYce
38QEPV3DSld6Et6rBywde2bbe/pqV8H+uucxDeS+v6eFtr1rhwrJZJwgA5VNWNhP
zmRexX2vZLb6SHJze5APEOWMAmKo2F6+LfwZNoQAmHzAgz4aHBg+fkdvCMe0CApL
pwtu65kEY5vdKCev9h1L6xnipfbjUyAQAb+ZIKBVmFxJHnoxm8uKtGyhx4p1FUIF
bmnTu353svmtB0KvlvYGb3DqC6P3PIR3A+xWFbzzkfUcp8m1w5qi74LAZBrVPo7v
ZUsrTRMvoZud9KhHfN9KMPVjvdgstoru9tAnTvJiU97IU/XzFU5XWZGEaArAAI4n
sT0NmFPgW8wVFkhgijPWRG0+yTMfKrNQY3rbtYp8GYl9QffTe69Z4LDVc1pNs1SH
rE4gLjwMphAAA46fSE/AayaKsg/aUOyB/PjuAh2VFrYroJ34KV5SXs7qhmX2CIEp
ejpsavYd7sUoWg7jV/ZSHyXmY/pnWxCptHROtCC7ZmGtj4Jn7nX/V1lkly4qIsd5
rxklJ1BYMBaFO4kcR0DFVMpl1OG3G2Sk3tHIIOEm17hfbuFYQJ3oZSZTUSTw8k0a
/cH0ulGZhRnpy8LTwYzJEVxtAt17sPhbazGcF5Q3tfn95JapfSgZBirDjGv1hr97
XPCUtV0yPyafu//Uj7zKj6zqCLPEk5yRCv3td2/RECB8uPWcs14YjOBGUdf/fQdx
rjAFCSURbKxJcq4AEJ780j1U2895hqBEMgnlFKV5NMTyoFQnVZbVDjWYfI5U8cdb
lGNTyt4bXQ0cHx7uObF5ZZVBi1G3QfKfcPjowepIL4nq3iT+NuW9LWjwWV/aYO6N
7p6DH2qy5a+MZnRczUABozwC/3q93YptYVdgUgEuxHnjjBykj1FZ9lavrWOjCO4V
09lFrIN/yxkwa1JQ7uHG+ZbYJ6qmAOcmMRuGb+SvJUcJghNSXtcUESKiIJ+sMSVJ
Ia4N5TLcHpfopCKyhTz2W7tcQhJsMkj+SUu1DZp5vZV1U1gnlGZQkCxsj98NZL2l
oVYMAtHg2kCXvcf6JRattmljHTTF0eiUwIxPzhJzPoEb2N6ODuqj/oqIRkLvzaN2
2WLdqR5jRxnStwqgvadUsK5EBSKhDX0JWFOd3h3dwRVGMsHDpM+0TaJgOPnaV10p
ajnLui7fS0IBIInxb7RG5CQHiHgzVjWt5e69tX/q3Ij4V5TUVn9VeupXi8bWuMbj
HOw/xUbxaUNGJWM8eBJvkLxPbPsd1NBPAWhy/V3jf3Hn+3ehYKcd1y8zfHIOolO9
kqomvtb9kqXG8vYrd8nCS5T3NAICeCCMK2/Gxwt5dFHfseHcpemHVf9Oj1/8b2Bf
iLv7/SPaVR3yGWynSkMljhFruCopGiWbAlHHp9lVKJtHROJsddUZ6KXEQKVvMcEh
hlQ2+BsW5NzHXM2Y/yuSmz5I0r4tTKdpFFdyEARunMCwlpgjmyeVOJN+KJlGYkxk
TbpvTVea5Esi3NzJm9mYpB04iZsqie8CB/7vs+7vumkBu/jqg+Ei+c2KavQgiZqe
97z1TDZjAsoW644uxgN5NsxWAfa/TnBTTMMxHHxCEfKy5oXbRIFWqbeGQykhyeoH
zK1dp0Q8AyGSCkuz4H1NdrOFGGSUUIkBINbUZMIREn8QTJxMwc3cczopWE2J34uM
U8A9fl2GT9JLFDxPzLtP6FuEbbHtlA72JSmwr7pk+0PDb7hBqJ4xEzdNk2BHueKJ
oMTPMeICv4auajzuHd83sddPydQ9FRLj8rpg8e4a4EKjnMCIZS9GE1sNOfXvbNLZ
/C9MwECwX7uLv7ypeVBBTj76Lft/7fPk1+1BTYbRV+Qj2i8U8RhInSr/1p/bQv3m
AzupoNuEupxE9b7k1F1z+uhkSjMJs3PH4HLPfdPIWqYLKL+lR4KBh3LAhD+f99q+
HclH6u4q5xPlF3rAtJztSn0dCcqSDJi3gOmITppxtgMAcHb/osRDUume68hTeifM
7FqhvzdtUAqbQ0v3JF4Ehhomvf6HsaW6HRE1cVwHSd5ivQQwaYsFM9RJpylOopLK
Avy09g4n5cU8Ejz2imBnsEBPE1sEGVw4/4BPfRW+RfwFHYnTHVvPP3Sk2PqenyCi
ZQocR5eeb687epr3LZGVlGjBhvjLcNCd2jeMDhKmQ5mJ8Qd6y9fTniE1uNbL9Mt/
62vsfRK8KcBJDlT10NJGbyBsUiKWc7tueTFhXU9afshrmTABK9wlbzgXMnZJMJUo
6Qmel57qsJWsqp94t5vpbo9KKFzJosuOa8fyvxwZS375z5t896xopuU6QBXUsajx
MQpMJ2r74A7cBJHAexF7V5AZr37SMHR8/HOxqiy+L9f1NoDLAkex33VeaJjyRZWX
u8o7z9bkZD7hLgGlc03EIqPQiMEkujl+hwtb+j2uHQcy0xJS/W/K/3Lja1Yk/xTk
5ID2UpECphNiFvD6/xztAvdZGaz9HoFTqOfcBk2pGupmf1H864W18+d0iXDr1yHc
4kLXk4+5hpLCcEJUcGXzEfoiY6wq12BFAWglgwVClqWIEhv+waFurIwa3AvKJCzE
drS4noap+EcFAl+YYiuWgOw1anROyHjVJD0njEFouNQHB0HCzyswBB6vtUM6VUh7
yhpbqM0rt/nx1JmISabekyjB3USIokWb306FJhLLr7AKUMttNSc4yxI9alOgQJJD
NIUTChg2c7tNW38vT6N7RC3f/Qr3xMmOPcMb5aGEkuiBy9GoE8kDV1uFN+vdDo4q
ZVqBLwRNQwOf0MYI2sj1rkpZ2e4oi/PYtvRHrO+bzShJHhDfZivFbgs8QfHfJg0I
BbWgbqgCuThLfvBK7SxQjLoK+j2cbLXvvLLvNPt2iVjUnhbvlz9P86lnjVffKtB6
Ke0ERQtRzcH1X9fqg7nX0KkwUaTpkQ6IEDHlMG170kwpZ/chmM5HKqhOLVMUYuX5
+cHtD8r2Up49aaLYQnOMmw9ciyP5nVyOXHdicbGLIfwMgpwd1b+RGeNka73r0F4z
/LvETY1Fwx/FQcve+Q+wpVDz/hS9xdqfEoBIvgF/ErqNCUhC/GvKosERM6YI2AhV
meoBHxcJA1nt3LVU1iYLe2PhVzxo0BZHv/Ca5+5SZNSZCh5edj3t3V5quqYbNn/5
4qmza/5FEqd0YGaRN6qCYLuiged/bVNz1sb/BQIAGkjzdg2I+xLJVmmJRnSuyNmC
8tKFNdMNNVJ3vy/qGrz/A0ATkD1lFm1Nad6jbDyky++tm7iCYkQJj7F9eGeDHikl
lgDueOJWqIGj3b9iDO4ooJYeh0wUKLyFUfNX1xeeoAX/lYd1w6OQ9b8EJ2qKcrVA
mBhvTwfecrMm4l7MbBbRmEHhBcG2oxFwfEbVaDhhHUH1uo9GRkEob+aLpbIzWAMP
DuTsjrACOsbDoi7h0BAA6OFAyO5hW+Zzf65YgzKsPBqPkv22sdP3XeLIoi/QMNh2
/sy5Mmw0/yRy/EqqKWmGfqX3cJ0m53TtedfYAVK99R54gamYQ+6kc87/ziipzxqI
TSRBguk8QPe5HiW2jVPqgfBkEZ9fpBC9sJI4sJnoJBlWI3k+Ta/yPo1nIeHIEcHY
BFc5TvqOuSTaKrDglm3iKra671ejZZqYyzoCEqbsf81n3vn4NzM1I8eLzg22Q4e6
pkf6MTyaxXRSB/4JeY/wILXGsYjqv1xVqqSwFbJAJXRt7u6L6nXWvb24NmNlEMpT
6YlKC+ErRsbeGWcSLR6ngHrhpJt1krotDEsV/09yUo0r+Iw7OKSqqWnfh7USsfnR
45rlLbigKdGVm1gE3/h/OgLrQb2G3/Tfgt/XGhTuUOnAOMll40DAmjvmlMiJrQ5s
WhxGUph0eJ/T9x9or+8KAVwFD5iSoD94H8QgYrZSkczLGKkfIuUrRMCKF36Q01R/
avoVJAvMpnztF9dAcSGMURaxTSrcA3ApeffbIGL77qKHE8pN688DBl6cDu/QOWZl
2xI/l01xb4D2nzBIHtsClrVMtv0z3IhGFQNnL06IkCsvNI1Z5YaRV85v6rreH99k
dGr9BzYmJb1iWBLrfwz1NpR+B9+xKRrhJIKryUBvFY6AxeAdFoilcsPmGEJFY8Wk
xpBPok7EH/a64qUjXDu3fJ/0vOMYTdfB3x8nzLRPg3YsF0QvWJ5d2qUNcpgP7btd
NdcUqhUzQM118lXAzo0mqGjjG0n7yqSy+uUc8aiDaNFplni3igS3dK1JzZ6pc6cg
I88wTSA+Tk9i0QE5l6m3f13CXfwYYl0cpSWp6Phb/tGZM8SC6pfjnr9ckaHwOjsI
k78wCwEATG4S6X+F5FrCA0B7uTada0PT+ah1YReKT38n5MRIvJ+5dYS3ud31HS8R
QdW0xWBOC8tDDp+TOXwKXa7A24jAk/X+Y6gNq/sj1JL0hqAcjBqvrG9aJriZ8r1g
A7pd5iYcBnGGikGx1k9vN+ykFRooqUTnMKYWzGBssW6CEuzb8LC/6Fg3Q8xU2+uE
uDbg15t8GbmkvbA4+BXMGCSLCdYFz/Gv+jkXHxNngzbc8UWVAfGGrkqYBCHlFMU8
q8UlLsS/FFsxMtKG+TUPuE5M+pLa+RlYj3dHuX9eFLcxVs4ABtOO4zOtmkQbCTA0
OuxOIsUNm2taWPCYJi3w0ApBZFXS6cm5W3MDl+ydJwgvRc/liC22WYp3246+tMX9
lmDKs9u+hDgVHAjCF1m200rzoGBzV7NG+unOARwbs3jTRUZlE7sNodwMtFGepUJC
QMWCfV95XFykz/JZfT3RUekesADU2+UatVQO1OEK5ihmg/9UaM7w/ZFuGfs3DqkI
Z2eRPzf778y2sxJubsUaBiik2/S0oSvVd22u9V4bF0Sdbq8+WbhRus9X4xigEQwC
RzwQJpfCoZZh5lxXVOZ4hmTVnJkfmwNdUgMU2cLE2+hy1BhN6gN+WRLjunP4e/d5
eNa/MQaYAjBZRZy+WvoJ4DXF2JLw1hQJ4F4jBP+bHm7DxVH1P7AVRMsYTdwwymQS
9WoeBNHGkK76hT2GCPcnRb8f6WzC5uc+9cqDZFiODcAwGPbBudpvEDFLeO4nagZ8
a0dXHyKq+uO1rrwgpbd3jupoYNweMlPmQF/NUaXo1GAKwu8CLILXQEEbqF+2PRP+
zaseNgb8Nco7AaPrhYitMlq0yEkdFJJdmDW8+y12HjRmY192D5G3oXZ9OI/i9V0V
RfcBKlh8nhujPjGgLgF9Rtz3S7DrbZk2GcFTrcqLXGIuyulPjTWXiEuBtsTUIuWe
XliUVsYf06q5LykZNle8OGAE6T/MHB/UqGpPAuG2RpdTeOEzgGL+xfDeFF53845/
IHAjyGMoypNjby+ihzntSDxX0BscBdhm40sBqkrRxLF3t/aJwBVSDCI/aPb7o4sj
2A5jHHB4az2tG2jq+TCLZYP0Q8DzzJ7wwW/nfIiip0fLE56nUtcm2v3tP20HNr1H
y440HDy1LfnAAaHlruVOXXz8s2ykMdHL3F2Gb5avuG8Fa5dUFeftL6Gpw61HWQT+
Ya//dZQzPr1sJfrHIhIWrEEu8ANbOBS6iJfI/UO4yhZl7Q/mwsmxXyO2SJXkUpS/
QesJJtMBVh+Je4sj+EnJTOIGSqYSTlHQNhnqh2PaZ+77AeB32rRbsxQnJo/P9V4e
nUSAaowy1eH/DKNmaRGhktSEMEnGZX2s8JoJtumRit2ZqUt586POyJhBYAbGzyDY
StpH2Jv1u8FFg1Y2s3EErBCg7dzYLQcG17Xee+ydDwQWILk9OdWhHPul6vUCug7A
JgtWJ9tXzYaLgWRWe/VWYJYfU52kihnYSkltEfOSSKkP49WWbarGfcUGzjyC8IAw
tUOHweeHbg4YAO3mwpnHzvqlhV/Cd9/IUWFArZHwg93vEDH6lJZF+GjANxAFM2Zs
Qzc36F8/17Zh3c0MREThLUtWNOBPygvXlmFWR8VpJbU7J2rqmt7c/UjkV9Ma1ydY
V+MiA7TYqjOnkEG0wIHqzowTFYDl31cYbBBkrwZVIPnptyqP6mbDwGfQRbtlE1Cs
oXX4rLUNrDF+mdcpJDHJShcfr2rGTk5J5CvJmAqNHlqX/URJyy6wZKhRycT94Vk6
M1W46wpbE9JD1JiR56kmgYIYGNyFZa4xS8qU2CKN0UfWjl13S8Kas+Ff/KbJnumQ
jt95U/XyCYMIAScC86JCus84swDRdjhsOF3ReEahg1rruR0X9s2/1qdTQZnuyRMG
4qrEawR2bO2pLHyZhcuTnn9AIb71tfs7T7AyHqa8XUN/oKSAzlXR7Qq88flHnp1f
RZ2iTaHoeeVWvmJx3+sLTLd5I/caX24fkhP5XgTFeVccwiT5eQFzb7bWwg7OqU1r
V/4+87hXsfhP7q5HkW0LUR22rry5nGyMwVCGpL0recR/nmTfi++JO9n1kX9l9j5u
jk0Xdq9XliU7+1H17XixQs5DR/evfcEjbuhDkMpaw+lmj9+P12IjRypvBuBUWAPl
eJuAL3AEEZvULG0qo7foqdiTon42onKgHtZa1QWekdpc+F3qaIPvX2SjwhI2xREW
LS/FnnNFq6IXiD9SXzg0AlXnXrKR1joLBC7Z5d0g0QYqfMawHgQNUHTe2EEQZiMT
6pXbt7GeT7b/0G8ggDTaz63jhV/4B6a6HR8y3WYd7kSuhZLiHacwOFgEQ/riZJqO
sTg2UQsmKPIfc8Aq4DeoAEvJDhem1i0qsN+yKhHA253i7+6sOoktd7ElekmYrcjy
U5bGrsRRptHVocv2iJEInBNiDAtmfPnGVPJuyn3z3LHGYoP6amqfkLAQqovpSOoq
tcPEiD9lmML81DKyl8k2GRRza3joUPwpSrtDIuWhifzd1KcvCaZntQHWOmyMpesK
6dJg18Ch6Z66L7XlfXojZlUIbsGvc6nKmLbPcrNmSt1MA6x4OtCd7AWNGIlzH6Pw
5QkpK4o5DnyDyR4ury9XSzySa/OMV7RRvHmWPRCB4KHke19JhiSqko1tKFfZbK0V
JUnShDE5CScDzzzgYDzTBwx5dldzPZ0gQ0vhVOCy/RY/A9hALMyvC3+DM1lvA/vJ
+Wd2I+Jj/1kZV8XQrwd+Md3T8XXh8AMoUadx3oHtpXVr1cD1uQCoxrQLNu9isUwz
dTss4IGIO9t3+0hMT4D/lJuw1Y9i9F9ErIx3m11dgv8+krr6CPTI8fnSopBg4Lpf
GCNolCA6sJ0fzq7ZTkvxfYmtzfJXBrBA1dOeI4Zrpnkx3wjy+w86X6z/185bp1Ok
5iwtkogAJeAdq0POoBhMpVCqZFEsNhyiGw7PKm3H4AnZ6ru3UUK8pELl7LQrGyvx
cXSnr8O+AigVleo51kziV/MQzCD/7SbkebV9TW95DlzXPBctSz61STU73DlxNQFz
eM+eLZow0eRY3bNHaDBkfAhVQ5iR2sM0N7G7OzFp/ZleXZc6qffssbMCCwNa0MJO
Oekg0vDpiMfnc0nH74aasskpJaMfcYu1ZGMYhxvj29mp0/bIOzyFBBO9ePnKBjIE
XLOux6nHl5qyqTZzwbM3TIQQc4p73Rf5Gq4UNlq+R1I8Tpe7UfkChvZam+HJP+2X
jwMo7qkUCOwH++WkpZRcLCDqNsGeVxzVoiQWIo1fZv5zQq+hSfULLd1XMj/ED5FN
ybnIi7Is4/aT2RGLaeQhdU4kPVBoAWQms0cAKVKLgyVl6y46AMH5NkalP0zSE+V0
YK5IQK1epqvRN9DI2myjZBUELAZNDvctN2fAXhtYz2IhJ4Sru1RafQUfa++uWNef
q8tE48qlsm86qUJ9gqXB8q65eTsbgrTN+Sb92YTZF/Wo6zcmLw+Uwxey4TBoEJvJ
tQidcZ+dFTfAK6OY0FLp4JsqnKc5rlmseBTekUH1UFWSKIh/T6OvgS71KBsXtXYO
GJHPWT6FX7C1h2byNCDMwX9CX311hLzXHzc7lXlt9gcMHRMnPD+Loc47fX52emMG
fT/F7aP286FVSMvS8HWXdi4S7RJmmuu/POM1/thn0uni2Wq55QxHFzkzTaKKfh6y
W/j0Ii6RXVUn+MCdu0JyxOQxqdStg2ZCr3lChc/GDdMxWF4eNGIcqWf2cUk/aX7v
fftPfi7X0eLobeu+3Jt/DjhjO1GO/ON/6k2I/8xVv+ZdkdbM7uiD7DtaESmYuZxx
As6U623GGLAgciQx5mTPOQFAiA+1jlW0PwpqcwdE0qXDUVDHv3BKhwQhrTtOM+l6
RO9n3iI7jgceXbLKfBlOZvnXDoM6siZpZwdgI0+73taGfrEh6QqeUOYWYH/DyVIv
LFz5c/NMaZ/moJ6rljW1sF91zviv22Gl+8eMKiHxrMf/M0aOrGZMbI31+qJfZcPX
bbZDeyuNbv1SoZKktNTyDqWefp39j0qSLr8NPWgby8PrGQjhS+8EoeI8t/Iu5Ces
LWSCPmf6g0ie50E5YJDuVcLVRARAXR1YFCnSOyqqT6XIMgQnPSL16aAOPHeapec8
CdC6a3+h7fJENZI+mtoXSJwHdsyz1ZgPOXx0xVGSVOviEK65UgU0UrXAPYOepUto
YEpp1EzjKsedY2PZtyu2IWVhIPCH3oPt6yDdEQHAGIbqTlfNNdHdod7zbHe3s59i
32RRZC/Gb3xXCMabqdjMep6jewnXWW75pSFtUraGBZlt6TxTbxkJnARF7fVxvMDy
VQi+53R4dfRJNMIfIqgDL5LSB0SKF+5IyJsnqPQBcrblIleb2X8DROHaB7JfghK0
spxL10JzhysbJnQ54JjOH5uWTv2eteDyWhISOUFm/nL0hbyYVxQQm+ev3kNLbXGR
7sy/MvxWSb2tCUXKUXBejrsI1gS/LmfkF8yK9uyInJqO/tFvYiAmqFH5+zx+dz23
o8+IU7mB8AsAfsJdE9+3AwogxZMuePqjtxPdKeF0s8wb3Y2Thh5TUXrwqBFbpOtD
AozUHMaNUJqgCtBxmlGATm9YwFL+gihpVeg601osvhOGqgvkl8/C8cjnccWHEdoN
JFRQavIo306BQ9O4oxOA79NRA5poG/nvVjRPH67ejXsSDJz6yAAd+pJ/zgaTegUo
hg9divVxhF5tCHK7hnjIFxPX28RyfnmRDfBkN6WEsK3l7XpjP5Nwh0qjwLU2jemp
6iCjHSGbqNtXn7mPuPje+VIRwZxc4Wpcu0BsinOBFjRQ0UPLSoJgx9p9cDRaRBgH
qiB8fTmAeeLf7DhNSAbwomsDfZQDBlvV5jBkp8dHF7Iqt0tJh/kJKAhcUy/xzWwR
pS1LPe/M+G0dS3mGvU0k5FTXgMlhX5TnjHHgflsDHmszopH0cocBGw7QQsJ6kxMl
ywRFIJHXyl6ETUkMtyHBQ4SMQcgTF1s0WjcjfwqbnO16HPCWOi3f19dIQTGIX3vN
v0gxchT8lAbEuAT239mfxAXZcT8bvszuQf0UB1qkhqbQATbvSKvv6J1a2WEao769
jyS8M5tilHgtqyT3GdfVUIOUkElgxhUnI4ZmPXUSz5aNMt4K0RN8HAdUYCPJ7V1r
SpIbJe/IEo/aUw3o7rGkA376Z78HZrCgrb/8QjVRfxiLCpd+WH9mmGVjDh+mpZ4G
qyvPld081zRMS+guy+oSYKj1KmqXSx8kA4BfnBjcIHjZU5BB5oqm96iR7kbVE5bq
/fKb8X1TGUIPwwEVR6y9vLMaeooeoIFedfoJ3kcJA1UIBv390kpbvHgi2pUfoxaH
gbcwJPyOrJblcl61pmkfztiZpezrZKOr7hKLHCea0mNDOAU8uVLSsrkJAhIM4aZ5
jaTJWiIJM1ktthFWnBJhowT6TBCRlnIh1NFVa+0+Mx2filz47i1iuB60g94fHOBK
eOGikMazpzJj8D9noSmVUtzNDaohzk3UdpJXdEKWF/s42k4MQKTV7uVfkJnoRPlY
Kn07VmRmsLWPqxiakzZUtu+DOSkjTmFYPd+F9kbz4x1dra/IwrIp+f3QKq+FLQtp
wILkJYe6Hnzom006MN3SBqjG6CbdwAcE/Dkln+9aSLjK5z2BA+1IO57jtRUeKkYl
1toCsQcAkKQmxr+uy9M+d3zupX2W4/gdzMJNaFMq7/KvyscFQEmczWK4GFWDo+xy
K46M0giD9UheBTIP99W41rVrdoRYIXOGm1DvBREH2LKWsrlKH9gfbCxQZ8T5t2Q+
A0yIRZOFgg/XMx8H3+JeDTt3mox4J0gqdGgrF2E44V7VUE9qnBvi13vOH4mzp8vB
lhPjl+tW1RkDDAoR4V+9/qiwqT0tub6vE1DwPUMh9jVj9D8w3Gqy6MObhJihJYNB
sxWeo8Z/affRGgRq71NV4UGvTFhFFfKzrfkzON0TjoHaiWbhp52ZkEPxff4oxjU5
pzzOt4aVNTPNuQxWeYaF0rH+3Wl38nAQkdLwJ3XiPGFetiExN4QASj/RveXZkgfF
v/RxQlTiblrFLAYsO3veLSbI/DWjjVHBpmFfK/XOvzfiEi/4kE1wjHZXk6jihJWk
j+HsNdRaSjSf11qIGL15SB77KuwXPxTDYpcmivqQxO02UZdrE9NWh5j5sNtIkXQn
pT2YzAWLfhIHrYoahmICCZFAKDJAegpLqrUv3yjmufZooT0FNJwkn31Y4D0Om901
u0RpiPovadWADNIer0hv80DohBBF2owrTgxnfzmdC4qF8/ffvnud3L7xtXbIDPcy
O/YX+S9pDpjtz4YZVyJ/cM21Fa2uYDrs4u5AxgvxI9CqT2S/pTRd4Ivn17xDjShY
wbhprYXXBKLaiYKsr/gQ2SCrsVcaw371jpmEnwJelTVM364OsBqWeA6jEroe7c15
zdLjiNOXDq/RHhJgWuNMIYjmJ+vpJBedII0PxDPWPR8onsUKtABBidpCVfO3vT/j
ZpmNuGKGw8og/60RJJYary7WAFIIWOVyGuXjrNkp0ZI8PY4n8KARLh/HRnckeNz9
KHl7O03ahGgOxnVkXG5UHw/A7KmZuXgCyK2timq3F83wUMbC983iWEUDU5mGHlrb
7bcpdP8QChucP06nCeTQjSeTc4kmW83KDK1uig4XGLAU23lnt2rxjwnJ0BLul8Xi
iQMFTRaLeF9qTKjkbuexCjN8lNe22iKBvF6tvQBkpF3HlhVVhnkh+rkyV/2iLPOl
PF7dBJ16ylXG8SN3LB0F6bNS7I/ugZ11M4rD+qdj/9dBogb47+jG58SWHFhzZZCh
k71Y6ywPQNdPDvhW/eqYd2iRukIPOzLegirBI1QYu5jQvNruIthVjBqQP73yLDPv
XMXP+g+njm7pgziL7uDyaciGAqW5kLefVLE/VwazFmPSqheJwekqWBSWfi9J/HZr
qOAOhYpG8qdpwP8AxPG52ymKblqK3UJzlXTzC8Hpv2lQ2LeFCYGBRd6wZsz5y7WZ
dXDTWr2eAph3ddtSyk+sSO8cWHSsmZmZp1gNzFfo0jD0zxFBWT3C3vyFDGmJda9/
/vvZKf60ULq1RXoNU5sXbq8c8gj9MHV0sH7x399VCACVh8WqPnzNVn3xsluU5/xe
qslxDY3ambcDD3uwP8K9MNKBdWSTam2iugNWr0UCfJc2l0Foh5j/Ggs1KMLy9GAk
k9TtxMmgcxj53KkcgpqvfQAuyQin5/aSBcd7aH3aiRZjPE2mQ0nEW1VPgwMQMOo3
4Q+nPYIMV82upse9QppugtCeaG9kmNhJCTXC7GS+mmGViCrI0T1sKV+9LJJGXn+5
t3fKrqwGI3NSiTwjImZRUXwVhFOgJScwWKPMgXtJab7gtb8n7XaU5UpMBxZ70kIX
p6x9f+PRK6TQ7IS+qm00agiicfD3Xdo/BXFklTseGPtgLGH6yFs9OcGFmxlifKrp
ig7qd8Mj5XzL1sFlladgOptG8qthqtrfrCtTVt6cUAZp4FhbQdBw3q/BoXpzgv9C
uV/XvhJT6DoRcocrkp31EhxSfQ2USuyJYFGZktYYENxWDJl08/BIkBX5VXFJwHSk
PI5vAzTm5xEzY493ks2UvAlEQfUoCw3y3E6+TlTZhDyMmfWrPkwZ94fVc3vC5jP7
DEFn/C1+s+45/8enbqXTFv0JWjkmOByVY0pXILUSQ+P20cxxYpOJFKngPcPOGDWz
NnzBnYDHl2d+HYHwS9RnmHQeKjeWh6pd+1FSdtbGihKMg26q+NRdqoel6/92YDhq
Vwx//JSuuRcgc9yJLc526PtjWpQqzgN78pdRpTpjYk1XmjLg/SY3oEBAQRkV05sO
3wYnU2QvF0iS7wTblDJIGFYJRufpX1t4ORhdcKpdcvqZJhQWIXVn7flB7yaF60xV
UcGSvN0KP+QTNG/OsiMkO/p3sPRziGh1GT+7cu59fBAMzCqU3toO0U0St6aL1DYn
W+1QMw/U/b+9lxqhlsh1PegsL1GCe0rlQ76HiUdGD+u/e9PU9o3shaYiSzIecFbF
htF/KNDmQtky0RG3n8ZJ8U5jfq1O6L1X2or+Gqld5UOfJDzeLkS/xw3LM0QaTqGE
A9cuJsJZ3oii0Zs5i/J5akxktQh5nomXDxU9QerhX+T7ArJ8/3Taqno8HolCkWyp
f4ZkzXsgdwfBN4VEF4k3f8do/o6mGNZxow5kGBnvWn/5pI2Bqq1BwrXksmSEUvVP
fpBQvHu3EBU52hYwTvvjskzvHbtgMnlkbHDPxmE8IRPEqsCnZAQqAMjcsuD7JOJn
03l6R3kkNnbUhBnL2I2ENjsfV7OImeGf5F0H2a7F5SYMqAd/qlSGo5Y0t/LKzpUE
7DYRYGumuG9qZbaBCQCo+/9TnsB2vDYdl7tTjc7cbxhh1BMh2MSqiwRNtAMFA1AP
YoOdq/ScUlvzoj4ZFOxJy2SRASsnpPt7sI0ZJ9HLod+OqduP95Beu6FpkDBQ9YEe
mlxiCYMerAaLU4TZKF4BjDgtlCa+b8fdk/CeXws4sQmxuyReyvqXkY37S3I66ZkQ
N7z8egHuP980TalCX3ZDaMvzg9T8I96FHVtCqeTUQGSEMubG1EzDaY18qJKINl/W
8BlF/vA3HyRQFjaI7ZVwWxop01PZM1SQukyfHWTTHK98pi/JJZz+ZaRgpq10/Ok7
Pc5a7S8RBAJcH5B+RfhxtF1l+bFirjW5c7AG4pa4092Ixa1Wnn1wWvES31KNk2Uv
hC2lQ+ghtGFrmIxokiXjfupqueHurs5VQRuFLrRcbsFqNDlPNbVLZCiStWESxplX
NFpAX+acXTv4+CPoCT0MVfsAsgoyvRaQlv30pRRk8Vv2+sUXcsFq+LqLjDUULUDa
CJnRjt3TWPmfiWlMi9IWhkJaY1ROdm+JXAWORKxgtRFEDESm4Mgyvv67i4mmtsmp
QBVuMLAPcYdVmNRatZkPDInpkWTcc7K5mxcaczZxFeGIrkLJMI6Ego32lVpbB78e
thbwlI3sfW/b1F8CISBJmWKnVlYCjsW57kWkP29HFQgTt55NNm850CTjDYBiTVjf
mF/az85TU9Ssdk5hbNWBeEvws7Yab72sBcQGUqQqFWJ62C0MLgkysujBlNzfynlp
ETnyn2Auhh87Uu+O23uw15zUFpv3JygGu1FpvBrsaf67mI5F1Fdl1F/CRk2aQa1G
60lsjOCeU0Xdr0SOVEnvgUrK0PiwLePxfUyNPsJFuZT02fxQeFG0nT5NMekiAE74
dMoUzXIc3KMD9ocTckyLhoTDqMXVC/2b960quTWcNER7CUKrZpDvA6gpjMEzpI3S
bjScHi1P8UlQB0rvEZb2p1+l/6PNQVq0PtMLNXjEBMu+itv/y2hec7pWt14Cs6pU
6e6r4zl+LGRWrr11u3obbR89Jdoo79hSu0m1i6o8gt1UQokMU+Q0gH9zOFJg14wo
2BoosvTfAOorgTBqI+PyERtCDG9Uy9rz2pZz6HQkiKUdPqSDOVcaSNXiEcWHAtr0
jlnKJlbefVy7ixqlU5zNvmRt18WmqNSTqGewYJF0p9YP/JoeqXrXGUYGLlJfKCXo
UNzcVqpfD5P0IIQcCIfOrPm75XRbXM10rd2wvRebYM4w2m46bbG3gUkPAW7rlVqk
dvBOACo1tUooa0jN1jZ8VWHoXmQSEnJsyV3LoAajoxkNHTLtsi3MXHMcGpDVPOlG
nvkeaNOBIwcJwltnZS/u1aGSV24w3SJwA08snszp+52/xrp7IrSq80Bu2BzZ3ueb
pVYLfUhqM1Rt3Yl2KM3VOaUfpdrtXHgMdo7dL9NMit+w7RbDJrBtWT/AxV9PNcrp
oOWF1xQG2jzqHK9fvFQZFWQYM5QiZQfUNoXWTOGFbSMcTJ2L3cCMhPmG5rJa1HZw
/6x/Rk0fK/tglCaM/cgIJaGZ37IRk+zYvibfdXV/l0I9L1rlpEQ3nQeicTponAzP
gAt5Tofiau9my7e13C7V49hJHz7mv8CmcHiZaU+p8ER6aLuqBz6td0Lq0ptmTwT6
F37YNdDx5Gy1GR+rDYiZB8mzFoG/6Nh0FQPnnYMuY6ukrzx4MLpQ7fe3YfHR2FnV
RT4QDrGrp1eo56Q2G7Knz+8V3GnccbFpv49jSOVKn7ov5zxthOu7wJg7Rlx1ijN7
b2Kv/fiHc5MpBp3n83DMUYwOwKCUInoj81gQI8p6tIOeeZID7O8yde9N7F1f4cYN
+A1qcJSg7yot4zNgZhsp1BmcbWBtBIdjD+Whib+pYARZKmqBjGwmQr6O9s25UgQJ
Y2smiEU9yBAQIWOEz01C9hahjEibUeHzTKkPFpUhXH37eqNZyRx11jXYkowKjKT5
zDqr+Xtbyri+hsueTvUtRVj1x/lu8V3iWghs5LaTivuJLJt1SdnjNUdQ8pMjFhcd
w81CfjbRw4EMuM4+odBmb75z7LxWZNID3BBNLlh8Vd4kbQbq/iGyRip9kr5TXgj8
9IR7nUBUGjEN23V47sEYjIrSVNmwG6WXeL08ipi/ehcZICU//ZfAsJZAAgRW9PQ2
K7XAMesOPHYKsIxLQTlW1zU1cOAtcip77Xh/q6EDUS3EKnwYj5xJHNrf//HzLJEy
ts9mVe+2v80EtMP8L34jfWlKhsFhLb7tdqhtquNmXV0hu+6gKLVUEpY8Juh8NDKo
I7udEGgktaIAvV7unxo1nt+bHuGartcIMFcFPVUPpqFkpfW9+PEZfsuSXahIi6Yx
aRWOQO64OzE0yYdUivkpMUytprQjGWIy4WwY7K9IZ6WZa/Pu7/QFT5T6tclAv4OP
oYswV1IrWWLT2ySsPEf4UwDcwyhYu1B77QXgKNpiZBZAnhp5OLe5TMIUlrZcGaFs
Y6fXIlb3IGimJYA+ZYQaVw3quAC127cR01u3+dTQyxf9X2XjXDn+jsMXGfEg2IjC
vRD2ZsbIdmIrU7xWU7VRhZJS0++Yz8c1eKnv++CCPkH2kXoIodppzil2rbDm5PTP
w+uZK/s5pXY0k9mfbLAR54jyIkr5KB6zgcrnu6OWhH6kMfgk55yqxttdoWdmMtHK
3e+BpnnKGjuxt602AiS/JF2BrdCpvg1nYI2gJUfofkkAfu5W7Vw3axZt4QUz54Ec
RoUX/faSOnD0a4bAWxrNEV8EI5KxqI2F0f/m/9CiadyeLexhH0owWSWqBXSj+EvX
uDpRTx7nOv0M97jWn+LiAIMDBSgz5cYvAVljzBufoQn59bCaayl3PBa847X568ru
9my6rnnT2vC/pHFd/d6D3Od0l0XPUA/ASUnqJ6ZTxMPd9U2SvOgVDAf7c87OT+er
4R0DylprPCeOMTIT68EDrBBUWnSpNftzbId+5tcNvrkrxXMRbqFRcADSemcbZxJD
sow7RPwHCU9e4AmnneYLY5KczsRNOz91BG9br1mZUTk0Sv6b0pWvIXlxibpMNgw7
nTX4zfGmLRBnTPQjE7Ho23s5tjCjihzuNLF528MD1Mka+p6arYU8etTbSMhPvzfY
Mpve24Nl59ZurULUk98nT6JttjSCv3DZ9I2VUy5phpJ7SVCz9tjcbH50F+B07m1Z
zq7X4UGb+3bk6f8zGMf2jixbcywn1z6OS6BY1nZrYRVG2tWvViyE3Nh7EiYzAe5B
/zosIh49VHem3ET3d861lViqAFFaHL3+s821GdoE3X3IEwDqbXiH2UmkyoBz7QSD
VZyCBXAYwnwQvClxKZpmOdcGmqbeU5TVFJ9/a3bqPadiI/YV0UKftjghclLpJ9hA
mXIU4b585ChK61FwD7eiupBMk1rpMV7fXR2uWNCGKIyu6paP6qlEwYpGpf3XKVJl
V/9A7xYo5ZjC5Ea6cGvfULvZLitcjkTxb94UsPhA5jVKxVghEmwsxLlWzwLZ4RTG
Toz4GY6zYZm/qa9mCzCSfgoCEIOpFVeOxmUQsiOLXufVuQG0w5ELiM0gtYGc7U8v
ouFoV2GKK5EDQMiBaq7mMLH2Kr5zLNTiBBK2vfxuAYxYuuiy1zLHEqrrb92q2yyS
TNbZJSodQsL1QpVGa+pYepyz4byUeDwVhwnUWnw77vXNgQglCwu4ukEwr4B9XLe8
oFwyB+py6cqBmPMkPq4Uqi9Uh4b7HUy7xeOzm1P3aqdwzN+i0OCSSu1h8Hp9dhM+
FVOHG3xj4ZrCF1R0EjwkSazv0aaqnSyde25E3IOvs1ZiaT/D2uKzjxMnypVgs3lm
ffw5gUyxZsYjUxEdVyVO6PcrLguN13na3eZtZ/Pjy7e4FjP0kBkWcAYyl1eFLMXb
+TDHoqOgv9YXKBGkb7IUkDblxAQCHfFOmphZCIxkDNE734ZTjBol9i2uDqMEFwUU
kiX5J5JCUEi5F4qNeHyjR5Y0vOUh9JC6mrb/Eahc+DVc5ft15qRL3zpT/zYsenv4
rtwgGkcntptgZsh6RFPULk6r4NNFqnECi9TCWJxiGaP85UWK/ei9vSdNtVZjOXKn
qlg2e1EXkCB6Unvs7Hxt7mxOlfNpiyRh+nkRTXFO+W6Qp5z+aKLud66lmLrNEuVx
7cP+pJ7Un6DG8Ldp1tjzb55XEhaM7CHn/vV36eiIEIgrowgheJpPwU05tnlkoe38
gFpaI0yGx0QJpd1Abv00oX6BqOnrdaPl0jibynTcjZn715brO4BuZNba5UXvMWpA
l06ir+jan0yYSLLHMBbJPLfGFQhWCubSVSrbf+btbJLalBu1QZrZ3e7dtS42zDT3
ht7VCDQJxFoiRQ0YDMW2qwTV0ZCNojn5WjBob/SJ2cr5NUpQTh5H3ixcwLgOI7dK
SX9grYof9BDxyhvUX5CQgy/aCg8R/Ba2Cx1FMwVusJdtVq4IyLdXbt43Ry+btAsb
dCCqnbjx621NwpVUT8aRuzmeCiTVojjktxBUFD2/Kk7B7iNPdtRMss+Mmgw7NYRK
PSRFdX0N4BNv52iUrGJUt3Yw8w9SzfyTlcZaCd3VoZu+uNGJBLdJDIiXu2d17PeH
EVPzOLdwwHdbpWENM2I/yFvuQGm/X2QO39aXp9Fx+VeUNxFp6qAEvf0TWQOchgyn
THwgj+vLsYeeRJRYwWuDrTvhGGMYW0+ingCiU+tz22vsJcF++rPNuGm5g/N6NVY/
MEAqh0S8h+HBbJOqwJcN8mXy6C/A/QBPfmwUYeGCO6bdFYz+QPyPE69Yxx3Xp5DB
/hM/V4kB607Hb+WddQlfMRzDzNT4B3WJDVQHFRJTPjSyQnm59m0uqEwFAveD0I1X
vmTJlWatGpLEQiClc+zpZxEOxwZYTLp1LbatxrH/svjMaLGQtZ/Z7ucvHws90IwQ
v9gs53CTDL7fBI9ldzZ7PN/Wc1YZ9yAeKS6PeGCPhgir2XQescfRfI8ofkpCckUB
zWMZYY34ssAfOQCrRCB1VD2HxG8EMaJBAgsILNp6rWcqBu86CbV9GBU1zDkUPjPK
HBkr5RZ2ZtPbb6B9zMA52k5w2VYLv2OtV3IKhDQ7Ms0tnMsgM8dD1lp8IWMv5mr0
1SxgH1Uulu3OzPTtBLvSnHWFVaz2w8a2U2KOiYY4IhNsh9gnOyinpOZ1Rp7dq2/0
R7Sjk+UNdVQojZTT7/jhf4DGD+Fy/cPpqcXCEBfnGJPAMR/lWnjBon8t7A1OwW6n
cBghRyhqpTX+e+yymhAE/8PfUVtKQhPjiprl6y5FHehUYwnki8Q/4gLvPtcGu8C+
AebI/05w7rvt6uuwJicv5fFO5avjZg9XMcN3BoZ6YjjhV5RlMWdl64lhEnZE3gtp
BYocfzSjecoonwuZQiNx6jZe/V28DwjbSgUOKdkX2VLauQZoqd/v9h1Qo7IrY3uR
OPnLtZ1k7hsjBrNPCA/kbMTfi94FnMx0pUGhHGhNOWUVQpXDf3BcwLuZlshzpp5D
zBihupwkbSJNaeszDC3pOdnf4Q5Y6pBnZco++rkVXPdsGftj/PfIJQ1tUYhnb6Cb
EWapVUzbvQRH2SMK6XQmmhcIweHQ5Wk+rjiPHCa4XpAVX1faPLzWLXz7ozqQdMGt
/1xozCnCG0V0InsDzp7NT2VP3liG54rZ8IoS2gymRYOkLuR3NISQ8PjWsPgypaPY
nzVSum1OSSnyCeiGkwqrVyAON0C9VGfGjoZ0+78LNFFIRMoNvJUPTGCSuHAuIAKa
J3nNgAviNl7P6fKm2GTAfWJ8VW01NCybsxpFRZW+Wb34PG2A/gdJm5S7SMa5yUnN
7IB7O33i0y4LUdlNWcXKr4VfeZU8FP6UqRJqHbUKap8hEiyBhLVqOpxScIJ9hfKt
KcBh0e6PUgCeLfvUnWt8Swzz1+ZsgysstlLJdoobm8rvFO70fSIVKSmONcj8+JMi
E+f54nE8IkRQvo9yahnV0OHF/QznmvLUx8nWhde2Ss4HRug+4sa5d9xnGWBVp71A
cRRsYEKsUOqwp/UvRFKjrlu3DWumQxkIrPbKM2YFZt/ETcOryljiBFkg2EZeAFXb
wliEgeBfP62xOrmui1oZoLEInN1OXlmjuB5vcC5yi02T99obPrzMyMXJUcgO2K2L
PjlNQMujpQ5e3FDhAmysTZ2pkB782qddKdPwcQaXkHY08as7ziUNTql7jFH43VAN
2lNMhVaI5KYQLcnmGb7pVE7T+qrBNic9Fps48piRVMY/2g1lEObcaq4QMqHB67eY
nB6p3dR0fIU8Pac1pc+yZSp+dFdbuinetggnOqYHbj7ygIEYHLxf+I5J9MPDqqo6
NhVKNNVUmHbEqMN5whP9r6kWROIV4+Uiiim2GlZ3/v7WhyTAwmCMv0LoDSJo7ZGf
piqJ/422U8PO/TpdquRr7ljYeoc21MR2btSPtIwHJAuUe9LfzkNp4xLY/RxiEsLw
TBVEbLHcUgY5PdTLi4QmHgOQBdGHbs2oHnw8phCyuarC/n/3rvZbeiqugdRDiub6
vHlHVBp35m8wIklQ2v4T9Pw3+6HHHZaaLGsCUuDowDVonHhex9HZLoUhtOXagqgu
H+sg+qEgy9un4gopq3OcFhoeuCIgXzfv82TK/lROQhbJvOjQp0WnegHaBhKMNGrL
6Y/YHmXTD1V4wtvhclnBVmckJADfTzaA1fS77FrvG6W3XrN1IjEbJTXPECktQdpG
Ln0m1YU2kMfQz17S2+Dh/xfArs467vGWIt1ls26wlAIT3RSs0sWrLAsZiQipmOpF
UcatupYHq8zRLYLzVrcpVUuyUgAlrCU/tiIXY6bisArPkbiyDT3dV+nr8Z63VXIn
AKrZpqJy+vAvs7YRETUBkLLBIUyoV9u851Bo5QB7Q900E+S4ZgFmriRV+s48eyWS
k4tlUX/TT0x1RVdNSHuWN8Wvas6omVvOUgAOpDtQqfXfL22P1sqStVxSZ8WTeNIk
ddIKJE8e3z6tcVB4JAMqoDlbYweS9GwVJpVKvsYXpA7iQhNTUOLdGqoIA4mCEgdy
nxPz13kGohUZHdlFr4TBPu1W0KiMmRAXgM1a93SLdKupiXMGspoD014dtK9dRZAP
7p1Gy4pLYbeCTBWMOoKe5n0tScIgxRvybGsbPG1SvByRKMWL2WxX37WAZfXGfoNq
rb8PJqFQ6wfDjHCnrnSmVDfcCP8VHg2L7xAGAeOgVuh60Hz3zKmsdop2jCuF+g4z
zU6AXxiK5qwR1TSFzuR217G7Rb0lvEq/CSgAoCTiwH6tNKPr1YeLd/USGal96Qvz
xVaH7KyGhhCeT9JirFqSI65hbuaJbziwc4QiJrOGpJGetjeuhXO42T5Okgce5+9W
EgHA9WR08xBgJHNgWbs/0xLITIneOqMRvxlCKIdlGSGW7Q+T9LsQCefCKMYXWj4W
XKVae7q4NOUN0kRIO1WrKz5uDroQVAs7mqqWGn4X2tkfb2qdPQwRoZC+1RTZQsza
SiCiuX9hQw2dZowStQzLfmM2SOenFGFkgX0ioGwkMfSvxthG7kQ5bxAt8o/w8Ihs
N3lJZR0GC5Pn6mpKreAf8ZTQqdmIarKfvX63oZKtHyRyxgrL1kbXsgWviDXe7qc2
sMFoCpbb0ZdbqaW0LfZ9ZXgB7I6/CLZVwl5PlBsMPbmWGgXIZFTbdQD+gnLXNGpP
USxtAaN/9gJU9YjOZSatm22LRL6MrC1rZ6OXys/WrpZInbdNf5JClERWX7kXA+ti
RqepuH3aXYJWlvMEkldn1FmSu5eQA7Gms2ckiNqZyrhG87M9APgqtezUXKGs/kCo
m+aTe9LjJOdQkHpnmOnpfUe19nZE1XZknSjLcb85lvGpsOf4K/4T0yj2Jh90i4+y
hDUHUk+AJvV+9RvARuIIIPAK/Aq9yAfJs/IQno/DZlz/WxNQVc/jBuRIULuLpiru
W+AvCOdCMNtM4LyX9ZTocEeqrVRryNAiTF1v77T5r4yUs7LRvFnBFL0BmpHeBllk
AUcv0084TO25Xo3wfU6GnKJLZFDugeMHZCH3pB8Uqjr/rODUHbVLh1Bpq3iQkVf8
TMsiSXxk5bxyvU3BCsA8YXK5gQzCJECrT8HQMec5zSmx86WTwlqJ2k/MfdRWPsbw
QZ+PesuYD6MZcj91UHZwTF8PCf7IDWyluc2ihz/9kEH90wL2s7aFgGKP96mW1BqC
gc5YXIjjVXakNJWvDduX8ms0DIwgEQe1DhjINHKgLQmsQFvwT5UKhsV7JMkjL354
pfrkLK5rerXAiVu4ukVUirRbVrK8p/C6LwNIcx7z9iuCqWuUQUImcm660XmI1Jpr
6fu44OfUZI9ZUt1rjmMPgteEvGGCMg4Sg9i3Agebrzn8J6jWI4Y3adeJvVGvOA0b
yhT1boAI1UUAqhPJPs+gA4TIKvZNAehnO2WtymMTn0HoUucEZVS/LZo90YWpkrNs
WADsZNf2dYuQqsmWT0x5rZyK8Yls/+yRMFC1g4+50xaPBZwiy/UnIvMH6QWdqM8G
COi3YPWzgi3hbmdJ+5zdcvw0oTRVKnh5y72NZ9smvctSP1/RrS7Cd2aa/cBHOV8l
E5W99JWSoO2xsxxgt7PZm7dZFDtWSQrUxP0/4+KTa0JqzS0QJ7SoWytusSJG06id
3orS5EcXPORm4YbpyDPiPR/3zSRgV1eaAzUsxigqr6t9/rjn/EJdn7O7DfKnEtUa
M3lejT6qKgMcbZF5eBbEBNVn8EketaAvFJOVhux0ji2DvVMC3WnsSXbjYYhKOlR3
RN7ZHEliLLipnAbgB6km60liZd8+e8Q0KuqQpYtw9L0WrsK1jT8+pw+rmv3nXZLX
6DH1+utI8Oy+4+Mvz1ilRCY11keDUNYY9sZju3ig9lk+wZre7iS/fEwYzSVqa7uV
0zHmz3GxZjGgJK9mr79XtteHVXI6+Llef3/vh9KkA2Glglq6FHnM3pC6sb58P2ZZ
lRmYpFwsDjMfhjwWp1n/18sAH0+u1CGnhuhRWsM1N7RWTuBqao88CwTmF3CLsxX6
pBRvRq4Hj6Oi4pKvTJuVksy5efxpid2AQMz/AbT2d9p6bPY9CZ2olURa3K715cRi
joMf7LVho35Lq21Xhxv+BNe7FgaX/WkxN71iFicMpANgKg/dv5daRPo7KLHXWbMR
lyw96tnLkIR7IiuOvY4WEYTq4JRG5/7KEIZGh8QpYj253d47RprU/jiMdF2PZ96B
GtHDu9mWWExfH4cZOEJYjssIHuguKTXUyf0FCYgyZTSR4v2LXbkizyqy06lxBtlK
5BZrztaXpZ+CzVFUcj/GMvOxt/Oo/utbnnbJeqv+0ziP0zQZows/r6rEj1+/AnPb
INqJpJcSIjHCOFvqOfxP/llMyrSLRi3ngCYFknF4/q69lWxI1Yr9x6sj6HVBaajM
dRNM0BcFc1BDqO3j8870wegyzKmqrg4e7fS0AJ+CZt2g5RtDdteCZkfZjChAomip
+UVoLL7GboBSzDJ0mu+XKr28i/+NowE/s3FhIyoZNNwfUOJV7X3H1JTj/Di1qY3d
DZehRWzLQSV8iwceodl1zzlDnvGkNBQy7nwpfZPipW7fZQe+LkZ5FVc4S+Xv3WMl
CzM9wNr4tv06MelwnrJQLAC7VtnwDtNV+cEYl1pKpFcV2rGxp4LkawVa08GNIXoP
1NaGwZ1awe3rMeZs5BNAd2/sPk0UR+ZW4nlPRC0xyeEMk9U3uPPzJkaPTk2p6Eig
koSjpPKfUzGIdCyMfsgX8ObofuOBFBPj3r4lnfgabKdXL6IGiB3FI+RerisxvZ3+
1F7Ar++GtSDtNBoqxov21iIgaBNRpV/ZP98BoVfVveUgUMjefIQP1Ps6PkFJ0z4Y
O3t94gWn4PPgZGkXCB2tISndkPdJlI+jWcGfg56TaRosBaxP4moP1L59fF8BIj/K
fOCcPUWQPMAfq1hL3Pz0GUAI12IwkzcoeFEz2tPsjkWqhukSVsMz8Mv02zD37v+C
NhJUx1ZmPlw1t/Sf+ARG/DeUy7761rvZvfCRYI3A4HG5eAQNGK3lYdFYySrOw0iO
BMQGE8Lz5GJuP4a7NtSkMLDfxDXU046JTn56Zf1qaY7Do9quE87Ab0YiCSECpPe4
7nsH9vx7wJkK/DgoBTN3n7BJ9koomYC5pFUoehaQDSlUcAH96NUJSfN8ZfpxA8cI
rFGxM6iry0NpyKbrwCKtIHqohT+dAk4rgKKMAFrC4MaTBpoLlRgbLsyAWK/ZYwmU
F1ZRzM1LnBfYvE+u/qk3h1xcKviLXCw8xMIn1jeZF7lF7jQS77GOytP8SX0M7k7m
PkRAKOchxrQf6l3PiZeGKPx/yCwKN920v9r9Aw9PEoH6NqDPU+veuB2Oggm6zW74
/LeJYFAHCoe37P30KRr0dfbJV2ne0agNjrRYT/X55C4BmELc/AHFmDNWB2bUNMdx
7NpCivwEdwd9IfO+A5qdZgC+xN2oqm5dvdZLa3sl5E/5Z6TW41M0WJNlCxmSl4VX
VFRpdqjRObqDo2JCzWxbEX25IyXrJcz2+++a/o8tuqgTeeiLt2XYjiW9soLULvLA
wYg7gs8EMIwqXSyeFjIU7sCMFjmYQJy0hL5GC+55SFPuuME1Qpg4QBbRYJW54z+m
Kx9QEy+3kPnC4JIQI6gaSKhQHzreAJRfVO838KHlagkLfPxnPl5d/JElOoadfsYK
mx55V9Bul0fOc0JJfVuzLLCSB8GXRcBGNQvYisvAZFbQ6dYQp/erXNe6rfRTjj07
7cln/Z1E1/bSKalY5OvpJ4Md0DZPov52F706vN9e46/+jCxwTTibHuFI7oeGzabl
3ERlTYZiQUkzTUNhjDZd1PKCCfwWrOaI4bCMOPAN70Cu32OnYK/6xsSeSB5PVzly
kDb2+CFft9E4W/fRcUWG+/488r9cWCMrRHUq/BSDx1dVW5sN7MsTLx1wi5O4jS2i
mDkOMsIdNtWXOjlMUktDa8+Pk57dIaNkBFocUyZYamw15VMw0HZ143hxjOb+ZBs6
sLQ+bedmgpiw+vRbjfte/e76f08yzvuQHUoU/E267nv+wHFTuJfVvKp3VxQr1McL
ZNaIFq9WDtBDD/z7PjxjkilOxU7X7mTsZwdqbCX2rhDnATpGItkjyA10OQplITOO
PZV3drh424LA98WaAXIj+YbJ1QTwBKeySKCEFHavs2Q1REFBeDaIgimdF2q1kPnb
USp/MDX8FWUjif9ZxOpPUhFFraAlKthNQCEX7oeyDiGDXhOpjneznug3SpII2fK5
cG8CK0fLvjb8HkdLOf4Auz8Ms3VA1dAkLDjqoKDcaVzgo8UAO84XLKgjqCAf68Yd
shlLXyAwbbD/fr5/4H9786FEs4+mklWboVbFJPjVvWRxohkFDzr1d1Zyt3wqciXl
/+kHt69p/4As0WS+w0Ve2pYVDgC5vnYg/lMXH0GrLcabiM1vHpm9HymAttcP/y1g
oNndXTM0vJykuD6eae7YmxCN2uf85wuYtCHUr+xttAOSIbREWtBscanVNVzKhxjO
qS791pIKh+kiImuOibWfUYAP39jhAa6KXHgdYf8NuGJLeaS0k9y0J5YSzMUJc5oK
MIlpLXFwh0Mg8mlu9HKwdxeZMej13d8SzNR18e/4pE6KXPHQwOjUI7T6w5TCvHHy
m5UK5ODCZ+IytX/UW0Lj6E8TBlC4hloDrEiN9hMFkDrfjvwSqPFKEhUAFjHk1Ma4
L00S+kexYnJ8z4XkGOVKOszklZgrSo/ewEJfswOzPev00hFGcy7KqGoeBJv2YiaV
+q++YKgsj7YTsd/QmKf0lF4QDqw85Yt/1yeU68kt1H9rsJ+veuE09SCwGudeZ5+T
EFn6IxHAnZTQvVNxv5fUnfZWqF5P/2oJC4EVV9J5/JJhGw/xYovSmkXWj9kmSalb
Du4YlIscH6Sp1XgSPw2+bZzxvehftHFUhH68EvmoQ2WidHehmb0uEIk2gXM64TIF
43PNKwylOsWiEP/tjqqx9KukoIkgBTLUzqGOlV4Q/la6HwdRr2NrWhshqMbsvSvp
PzPWXU9IpUI/Z9799NYwjaiO7/yRXqSW8LkvUV1fvfyuxN7WlnJFQck0txUdpfXz
D/owpx56E9eXWmRThjhCiQChm0NVbXkzmPMAp9tgI3STTguAktU1K1XmvmP7F8St
fOFTGTofIS5wwp/r5prBzx3B+MOX5dPkWSbsYvbuh3w0f3odsFoTDFCucxI0XnnP
cuqiuyKZYLnhyHbUuF2ClIerLsjaY0rzpwSGQTd8s+qNDKyAatQpBVijtVrCLbK3
ji2FEh5pnzj+anrYpDBkDdZJ3NuBN47X+gYhpZe5BnQjY33QuQ/1f4BHP/oO5FlF
DelvrhL2bf44Q14vUyFTuqNwV43KCSnFdpAnj/Rm3xaXbN4bD7+Jm+xXwwCiNX8z
iHiht1oVDPuQTSWg4PvLEfMv4812xkiw3k8o3atDpYrd7zd0IuDg/hedZx8tIT6t
7gpw0CfVbmsSN4abZrrrxjumyfO9mOisa0Tn071nS6AubBAg5xHoYZocrlU/4q+s
/zCfMNBV9wdik2AtcxZ+Ysd4heZmY5GmpYdxL1cNHUI42xocpMnywQamr63WJgt9
tf62zBfm8g5oVqDDC+ANgofo4W+z9Nikzsf+kwYwpMMt6hOAVZQ09b3DSKQwb/Pg
6hv5gfs4tDMxzTCtzEwn2p6KUpFJzneeYs60GK7+rVePc0T4wn9tio6/kabd26nR
7SEBfzWh+Atja+H+UXilYr3e4UAHeO7e1weCvrcpnQC5Bh2Ll77TcvyMvZDswH8f
iAPQHh/1uVQyo/hPAzgSeiCeul+9xNxjgGFNdBr0QT8evrMSE1fe6wNmM+hMgZJG
gLMLTklm4UlC7pcmsuuUhidJlzagOaXsDITaO2KrjPIY2UTaiZeDFRwU7crVLHvR
pfZfOAVcMlFs+V9UTqx7VyrHPnQQNWbNZOQBV8UjhQhpqWOQEYZOpgunXg04h3NU
hAEXhIeJdSdOdSN+3mDJNFucy7rtsp2cReGj2Xx0cyU5Gz0QNEBUeDVHlHH0J6+e
pkGA2r/fTrgq9F7M764DKhHTJ82U9wO8ie9FGk7thzJiixXygmUScLdT+sPHkhtt
9aDRwnjlQVU/5yF6mZbaRcgp2zI126fCYnwST0VrbhVmMGPeoEpS4OyNFAP73HR4
I5hnagSZTmh5WsqeYN3+Nr9K8CAVg9NgkZkw9dEJtyTOJdczdec2dWKfSSalmD+k
L9umRINCees0sQEt6sfmseN/6PZdXvezK0MGNgkVr4YeGkfjR8D+0Olf++DlDIt6
mV0X+frjWUrFQb7rPS88UtYy2pe4/TAUeY6s6MGFpaXDeH5cidp7YGdZ4b1Rw8EG
Js82dfQ+ZphBKOGkCx8whm3+JEjNiC9zIPzRi2nz+9P5JqTYnOn7x9UeZqm+auJB
hg49TBsLroxlrPW1Q1R/XKv9fTJpS1NiaHxQe1OMI7CKGhKgLVUJ1JXVjq0pZYs7
Yk/s5kp3rXhwrhfb8nmTOlTSybqPXdkDNdLo1JoyrQJa4WqBEWwSnHoglQ/LnHv7
cukDzWDLdjg3L0fqAqArnLmoOWFVycyzJ1paU07v3R7ibh2HCm4giZvDRVudN7z5
EsmrlWYKnjrxs7AGTd9XJbFDUCj9sPVeD3dTEroMbklE+6EoczB2npBqN9mI1RzX
wgVD55ZNGfMEJZx8UIFZUs9pUpVuWBNM+5ITRq+SLPr56aF/UDxQzpuuTtgGl+UP
EhJtJoXeTLhNvcStpxD0H1MA1JOtlQePoCqDD0WzHyd0Hlt/VCWfYUVInN5EyQ3R
TRNaKykMk3TAxvg7YyrsBUJQUlk8OT4CcElq3JC97dMxQghW71pTSSenzG6By9hT
8v4wehWZNyal/Ap2R3UYvyF8SSz/g3jo7X1frz162t06aHpQm6K2n5J0DCm6O7Oa
UZjS9I2GF4cSrfiljW2Ull1VOFq2upD10p0KXey/5/V4vt2XP45cBtdoXuyM43pb
v8F7+0lP9XsXpZDxoVLYQMHRlPF/gK/OHEaju+GX2LX1EAn6aTPvxz2GM5OLiCQF
Tu2z+aBU0yxSsWba/pR5xL52Nraq1EkzAWB0QGe69Kwl44hm8XKEWHaTWn9Eh/QD
IPylpAW1UJu5KFyDToG2rXt8mvyHBKEtFyfzwfk2TgbFBlhblYBr/ccANFqFX+jQ
uk20AJFmxNJcIgV099/aM902gtIIEGhcLCNGwngBjRk1afKcbIRpa4nVdzw4oqC8
9xkuxh7XJJQteKxLZO+Z6S71e2vjNg99pcD3PmwH2x6n4URMNuyINrt42hdfaL6j
kpifdJldt+TSKQISVqgpmI9lOkkux14ZTMOSEx3aoztLLXE1wrwgK8GHXadHBWKi
2ptml8WOaDg1t7CeDkCQZgmxzgurTgQgIrcBY+fObqxR3YUd57TkvQh2wSqxPXOi
Synd+lSGY/S8EfkEf9XFvmvoNdqI/PXNL2aOz75vWhkM3EzcLLmv1aVvqhj0Sxqc
/PzIdtq9xiPScgjzyNR90bFovz/jShkPCFz3LoOAa+sot+2e0jbcOgJi8250L3O7
mQOrtkgw8ICZlw6TiwrOhag/KlHSvis8HBj5LdmJnsESQxAfLOxSQ0WEmLG6PM1d
jCzpUzlRA5o4Ib2JWheiI55+tDSIdjdQj5erDgckIba/aXW1oryMHrAiOekfE17b
WaLYQmsKPcu+6CFF1xdY+kDdg/zbglHhQwWX/H0fg8YDsCc43/MFjBtmcRRunX1x
SnU1ByUQ29QaEC0gzu1fVm5OqZqgdHyZJY/eJk4qr/njnDw5qNZWmhe2W9Zwojpc
A2vUaDgEBsFVgENgxuBL0FS953Q4zgKAaOwRpqtZCMFX1Jyr9at6aR6T2kltjQNo
WjYoGFo+weXguktHYwUg3ROce1MfG4ldBrQ+6bdSFuEuCIZ01jvpgHWO6DFt7Gaa
hd9WPo98eEd3JP8LSWmorK3jADjAyQn844z6FIVzMQjCURUQBh+Ndu/U83MzKDqj
atQafifuKWFwE5omEFUu/FhZvrTd6SVnY1/WkUNLtKHbGXu7fRzCxI5YB/hl9HbP
suRWOGX+eJHFYL6vF9ksnJPTtgvGbZdV9/n/cw5of99rSmyNlnQoQX1foxPBCyMK
2w0PMzoHtBAA6Km1wr5aVzmZYhtarekXlo6DEkCYaUIf+4DQlM3/98ERh4GEccy0
OdqJFPszr+FgifqkkLhChf3fvFN8e07dVR5ADZaP35mM+l7po6Q7PQpShto7tcEM
LWW4emEv48rJc8YyezCJVG5ZVMyihCg8j11KbVrTxKkTT1X0fOcOS+M8Mw7vZ3Pi
BgMZJL84Uc5JgJLU7UFkQoSDdQaE+6pvYvdl00ILLbSl35OAxS5K+Be/A8MRqWne
qJMffiZV2gA5CZ6IB6dOjapTPqh6hxRN2AsMK+cvTqIjI4DxflUDp9nd5Pea9Oxu
tcSwaEk/TBmG0yqCMfLOrmKLF4CJZLjBcUgCLZfBwNNt/azqazGzDgpcmPLKTrP8
BGVa6Qjxpg1drNp5D5IMe9F9KR47P6SLhajQ9D1zFZHZXnf48lkDKK1NLk3Iz6P+
NZYRCFB4rQV9PxgyJaeX4zK1z6Imye8yYb8Ih4otmkAArMF2KY7W0YnwUBeLQ/1P
COXHwKfAyIBKpIaohLIGgmdGNHygOBJ2mKLRQmnjyYLILjneKGd5ky8l+uhuJC+E
y2yKDZ2H0D/oSIuNEbaJ48thNh1+QppmU09HBgh+hScXP5UhynnIeZxDnSHPpFNp
PQu/U5Qm0xlZyRUgyvez6mmC9I/7FBIFzC0OChxFLKUUbBopsBVAZM6IEe0zbv26
tjsvA5aNQIfp5JufSma6bXBkRjDj+CtzlXZfGqwA5ZmXaKh6RLigGIprxAUvfKgD
dad8v4qIHA8uJufMX8AGYPc4pl8MG2y8Ax2tW+H6nfZCtabitxm8YFHtvHB5bxtw
VW5pkey1IlSsXDMfEOldomvzjwH8yUBbB+9uXdvpJUyCiFbHyxCkLlyGoEXjhpek
IHtxGpQ+KCiz9sPggwlD9YU3x0nFrBadLPH7siNQUCB9HgRI6Z7Ata8mlX+YPH61
Mk8p8RzHrMBImujgloiV6PRnjS0yTwZzJFu8UxrW3ZDdm/UDlTfdAkpRXPsEpDQ/
deo4tB8C0f4t8DpLKJU21K4TMV4zFP6Py++I8jSc3UU0o0/NGefchCvOBk/SpX4h
ZcV+6XDx0ACr1r6YJuo3j5dZBV5bEm2rwBIeCaJhl7blMNij6VR0KSmimfO63yNg
89jOKtDlFoIofvLSjmZnyhThgYdcCOhYTzMuxb18A1sXwVeNFfHc3FJq3UCl3zvO
aNOi0DH6GH9C4FC8pK/PtB3U3yBjNn4EqMYvNClWgTLo+1Qud/Atvf4+rRBdvBV0
5VzprkLlhjNSdOrl5X7KayjmHgbvb45FWaGFj77QRTfcfFVnzcOXdosQSb1xbdMR
7PGkWzjT4uxYOH8sA+fX4cO+y2PtcJfqzFb62dnmwZ62o5MwRcKVlOCbH+iBc61f
0sdznl80qm5zZktDKYM48YbWzwBIz0exwf5XAaej+kIZyfsYMPDm0qzKisam44ef
pvZeQw+70xQIGbpVbCWu5+BV40E544OIGP8ykLuOsOjSf7yUi6v6nck6t7XSo20C
4lE5lN/pufp09YybjqRgF4SHWQrsXnGqAw7f5/BHnXCfT9XRduaGPE5CiD5KNBDw
fMsekjFGCaplTY0KYR6Q+Bt3RAGENhOyFAZd6TH8SmtGbnYOCYctKo47Rw4iMUcP
4qdfQkPB4i31fDu2m4XHJ3RiI4viYFeJxjZzqV16PLM6onvZOOL8YBa+kGbFPY0P
ncCTZToqYK01XxS/P/DMZZ0OXoAPz7ggf85762+Zuzo2l/JjTAcb9esvbo7fetnv
7ioM6nTSvRtrmvE7/YIMjzPDTIlLNff5o1bJPZ5LG65G5Opsz6aru4uGXu0QkjjW
CunejyVWb4vFzV6rYTDs+eUtnCqQlevs64JL4pp2JCkWSnmemNOAv+9Yk1wRqOTV
1HqcxScs88yEUmfJYfao6JqrFnjpceNd1A1VKM6+3IEjoIPfuC85X7h401pHB3NS
RLwRt8ncirbuefZzp8PBrgqaaarKD7eUEHs8ClJDSeCfeeUM6yDWJgd60KpSsj0+
K1wUaF5GStFz4YaNUONtF7JJ3e6uT3csFK7ib5nQcPhnc2ZuT/xTCqWAUEa2zfc5
BQDqZkpeV8Pmd+yiedO13WDLwdlf8GF0cyXbnUPhFDbGquAZhL+CYtlIn8DLHNqF
JZ8Q6EXQ9e3ViVeXzNzcgFlYqjY7sWilnTH4klcPdeZB45jre8b3ovUPj9zlKiax
IHCcYGMb86ZtvS4Yinjb01dRZiUH/REh8yPp2hZpXdcAX5wITCv+m/w/T8xUrSdK
hYg4hxKxDzhLPfERnqjTC9E86TNTn4oXGdxG3/7VSSwZQuNmZ4D932fYhASlr3ZE
q+gb+Vazc2Rg4vrz2Ro8vzjEhP07lkY2HUTQTwmec96u566YV7If9R+U5YOf4BC+
/2kzUwkGSg39LE1EPe5TtLioXDglE8uEw/1MTvmLYb3rzZ8CAEE5aHd4MJU2kdRZ
8MaigOGZYIHNbzxggGI/tIvaXe6wjadWOamy0DwbDfHbvmD6B52Znv+DBOv7EQYg
GqeVPohmgokcEJ8b6c8RIcT0rhQcgm80kv/ga2kDRF3vlU0ye4EcLUvqS6U7AXYB
PhSeVzMaSL66c7p7DaQ81xKu3q/Wlnt4TFqvSDeHo386tlRRH4E20VkfBx40cwWO
cFc/Uasl/bc4ZJK+Nq+3ATjpgE4HFq5pIO+Rxpd7mI4HVt34Xus8p+aGyGzjWK75
SJnJEJ48fxzo80pKD2GiAFBRjg8fPqNtr5AQynVHEnwoXxsGhz+p7gCPHrhCHf9W
rvmhvsRTila+/bZN/oFHeMElrOKIGemgyZLcY8Z92NeEHtTfLXMw2WGpLSmrnuAA
ahp7m61a2LnlJ+2sv9O7GeEwWt7DyYxJyc5pnaXF/++btNA4O7JRvBhdQxFh//Rf
98jcP3jumorm/drTOY+O+ZPfiYTa8ObBNzRRgTWbLWXNY6tUnrlP4VrxPcusVhtL
9bXj2N6oCmRXmJjjWR6VNaBdGHsKISyHNA4m/gu9fclSeCLNa87xQggppZuPC/Ke
C/9+y994eKO1iEo9UWRnX6HX+k4mhqnfXPXDn881oKiJAtTtjk0CMnhuUgdY9VW+
3klU+J71zJBIK8x6tcbHJOooC0eRiW17YqN35uO4O5RxhFCkqx+LKNqxMB8ifMrK
etYffD+Fikk8RWypa7UlV3dt7f+vCmJo8OnBVpaWKYkv2YcjAa/VW01ydzMTbKUt
IK3PhNl9ZW/wUOWjSXv353ilE859SnHJU2p/6J+5G+MdluQqR8IF7wlxK6hC5VYU
9UtLj/CVC7hXEbnvLuwLDHtjLs1pNdao4+KfO6qHDKe6PyEJG56LnTpYU17IULGJ
JtAtyhZp0Su9bjPOjnRej1LB4Id5yI0996CszEqB6ID1rzBjpuOn+VgcyOpnyCB5
6lhtGG1bWTgGNZjF44Hy9DJrFPX0ieth1cgxCl/bqV7SucdANZ3eOgTAA2ZmVPU0
jBATIliOBpugKUsLBWNhFYonDzR5WugbhH/1HuEpPf9HPwEF7YtSvuSDHs5CAMo+
JZuEWbIVILnY60mhwZPh8JH5XC8nCwfPsbnPeysck8yYsfVAJy+a2KYm6Pycvgp9
SyFNfPmVsqeek5Jf+jS7Jm7eBuOHOgEmq4LO3pc7JcUgkhmB6puaqtExEWqXeMe3
ZfMhhKFhqt4o4x/YQXWfKw56jkWaA1H4JhgeDEIKFT7+9qCwrWgJjB3j3HXli0NL
/O2H2zueubfFdjepwB9tlDvIqN/V0QDgCf/w0aL/z5mdfa9Rby3OVMACwmaWSMd2
xYurZgbl6EueaV2xj9YiK2SEmOiwGLAbgMxZTCcOYNEwDmrAFGGjmfWbjdQhTSwL
Sr8IKf3LE1+ELE08X276hfly/I9RMEUwNq0wYeNPRtimMk5cFXzlo94MNliCIRVP
JctpnxsHo9JLV1c1wohGe5uON3h6VJ9WSt5VlEQHa1UEv+pn+y11PKEUPF2MLjsa
6NStoHf09XMAm5FeJMCmZH0w49p81RCBz/SGTW2tVV8gdFh4c+/LQWdCcQf5QYVB
iLqLfKc7yKbVeL0ms/Wr1/l0XdGX2QAlgHfQ0R/ibAG0NQReXpfVkw/OcvA20xn4
LGLUFYZUP4rxcFCky2JtIT0PVD40LGQHLZZH5F+RWmMNSE5NyLVsvE/YnZVdbDph
1EEMioOnC+p3Tkv1cQo9JyG2UEIyyzHWjra2xwjyVvwx7fS0EJt/CqQ4cjfq9iiG
a2jLRRCI29Y7I1QbUbVe0xuIUcMdv7XO9x8apEtdB605yT6SjU9bgTjKpDYUrdrV
ud+eGeS2Fr8sDeucrYGmMEChr3d4HlhF8F1MdMzB/OjcoEfyDZLChIjpQ9gK6aCL
j9WtVcy6llFgirsxxKZrJzdY7hryL9cHmif5HyuL9so6T3BCfIYyKG/IS6KdVW1Z
NSRnM8buqKs6R6SDtBXB3lMHgFlDT4mxxaxSx2KG0oEDhtT1VKkXPtv6Xpd51yyY
7LfvdXZSJbC2/PsvizN4QdIdKOacn7JoVLIcYFcvc/4Y9A/JHAwvWIkNJcobXAAz
iV+crCM8kl1x5uCw8rmNFfwuXaX3E6HLDW2dHWRK3Nghd1F9GcyGXilufl08eh/0
AotK+5UKLZoQiiDc0oew+vzJOY6LFTeLK5umKal40r039xg0xEfrU8rxYh8aWfts
+b672XDBT1NLyTuBOUEX/GKXIXhFuvZw6hT62DHXE5BnfwXMaSFOqa41KOmgm+sQ
BsjkPd04ukZnPiQzI7xfoC2vbBNWSHQvmSsuqLncvkVCfwOFd02l2ZbtY/8cryNm
ssFScKgVS8Rk8dN3pNgLYBDoRq8tvJLFxqhIO+kytxpvkIQAbLqG/gW4SYNrV2BF
GFmUs1B3xdXlPZXd7jTngCM/ZBAExdLDleRK1Yls3Nx4U2MfJRs/ePkaohWj72gw
CEdvwoaosDEQfu58SZ4gXcritr3JDE/tlDfz8Qr4JBVRMDHlIZyo3bhKpcFGIlgM
mCAEF85x0eUG6Gs1V+UPQ3eGnIt+jVNc5MHUJPbNSHrHYKLKCSoXm9mw8iULLvJv
8aq/58I9GCwk4Nkbosnez61rQbzvE7hAnjjfW7cmpnytnxrU0FbE64LvIDd2N2N3
8gUA7h/UXUydzcrSkq/n5Xy8T0mg54cBI90yxkpfZWqJHnk5bnToGRgWBTdJLYkm
FMy7toxYp8AaaOJWDmhnfSpLkdfw/kE9XtrcX2JlaZXSXt+Z7JWNUbn0N0oiIz0g
uqJ/mogLp4P5VsGkVppVKQ44b/BkjP48JynToxQ9i9cW+EWuftE+LqTp9kIR8Ja5
9I9/QUDYsw4lXD2BUaOLnN4REFqV4MivbMJWUjZqRIcAoooL3423a4gp2cRgR1Ri
+rh+eVuEeQ2JXEBPplziR2/wIVBKt+joVunEjWdFJjQmguwFST9R73ibnWRCiQkS
9J2xjAnCQtiSyWlNpDpPWCWwdQnAkpCIPGQ7W9X01ta4sGHBLQVi2J0pjvu9xx1a
I1TtUecH3DtthRoXnGxjlMLDkphGngenJsewEvxDOVsYrKFKJTVx6X5Lr8kRd9ax
sT528ER8JK33XGCBpXyocBRmFeYfMKT4T8RBcvfRGmCaobjw/le0Audo7nwiIvP4
sjFuGRdnPgxsFqm7xEO8CifkaOGK3ZY42zQ+l7UnP4KdUUtVYVk4eH5tny4y41iV
lTKMD703gKia4DOGs3dKIx6AOGBi/qEhyS0B/kfjxlRTlPY4WTez98NJPWRsEBAT
ICD1LororfTWlDL0sVq75eICTFwO9n7q7omBRY5h+uzmfUo46eItueHHBfHbRCFt
cGd6hPUmcO9CdGZ0DrynUDLA9rGctOZKo0NleiVd/DYCv+cDvKTJvj/MJCX2L+1H
E+ZYi4ovH7kK7vuytR6/HtV1dX1NWGbHJH2lmhIImeasumf7LEjPCAtf4nMO86Il
NIRxHtko2sw9M3YTWx37uVrYoeYoZFJqvr7tyT7BGwbMVPxdn5Y5dvgpnMlBxoFL
jVQPlgtrwYcbeau63s+8QUYQ8Y2LW7010nDGELQlRYBN51xmktbFCfz0l1GBxIAE
iE1rjn3hZXM0f1v9Q4KwFy/0oOfBLCAwp2XZsv4mHpsSZR8JXh9naChljJSOhuCU
oWL+6A4mg/rMTt8YOlLUwoqsuAXrKri/i5nEp3TA9Rq/ou2dSBOtwBPfx0CjFenV
v/Cgz7pzK4VPwcFmGCvBYsrxIGKIpkTzHREQL32HTh4NtTiUiMWebLVm4zfw51BR
ac+s2SV7erMWJJMKudrWIaI4z5tTSFNeYJjwyH60yFB/Yujuu1pYsW7Hu4AG772f
Xbys7VlqmGLW+ls/ez2sJl8HsuaMOFUQLk980+tbhN2WAlJt5vLwF78gFGp78uIZ
PWDF98TAcz8jyVTfv9rOnG4QqDI7UMocEY4/bl1ejy1Xoq8AoU0HDvUw46mAn5+d
GegYQ7bT+W+Bx7dpaPNIGLVXKIhnTAKnST48jNjdKPoRim93xracBNnALg9iXHd2
yYHs8WqbqbXJYatslLdXGeYt7tuH9CubEslfBE8NCGKTLssw/6eyi6TEGx8V/+QN
M9bVcZzAZd0Gvo35bazCpIfXqGFmur65hjXw0BsA5i6/nfAJ4GOZvGtKE/oQtV29
FTQionD7GxCCnKUcOulbdHVCD53kM/G3X6X6/RiiP8m06DCRDzGQAhtHNDVMSJrL
esb9sgjgdFfEwUU/WDoQ4yXwXjEkaSQ37wqbbUelF6y0zlFqJmuM3PrWzsJl1SD7
jfYFhpeSpiu077y3YIhRBYKrY0L143WAr42+5lYLpVKdfiFVQMu3LX+O0nEc4+u8
X/IXYGCGGFPuaJZmNhNhrmwMqBNBTl3aKyEq1ilojocEw8qENdDZMiw7NEl8IG0f
nQZvjhqLLgbPgSRyb19SiAgV34Z4KunMVwbrg7/LYfwmI/DamYESjL1EzSZJd9fX
9MsLoBX9P+wiwX9wGeO9VB2Osd3J5xqC6K6hbV6ERM5Aq57RZhChKVyxtk/3z7VA
gNsLg9vQGUG8LjFGll97ASkMAOe7obzbYuNq99tUKl1Zm7vmLynPZEP7d7J20qUy
g87e1ejLB1EY2cKLOjO9Fsuvocj21n4bwPB3gDiWGaCPTV8N6qY+Kgt5S8zp2rLN
mtLH2602IBxDrFj0S7Jho3scZAryi8Hcd31+n3ejanOHY47ZDwoG2UyepMzIu6Ck
LmvGxgNka9WX8+T1SISUVdtxPDjxtsu9lMVJzTxVqAwy+gRjxCUoLChkvTfPRvO1
C2LIKKE/YWyrNuKASol68HJJzlwRZWTW6UqUZq6ht+2ak/MaQxDuXtHRWp4EQ8NT
XtA3pRUx3vNUPKj4Kvd2rirBmDZnYDn6bhFBy5k0YFOnrdyk+OQhGNKjnhQEJv3p
c1fQ57bEsNQdM06hKvAgdpyi33UkQmFp1Cf39veXBghjaAom7IglTqQCvppq5kv6
XvLfiFsyv2+3cqo62ADdmpd/kV9F1VMdbRcT2/E92PHcsAbBpYweJd5rx0SnnALm
eaPJ/Gl0hMekn4uA8G4eENKQynoETX1Fmd2cNN5uONnwIOKFsELlm00Spep1NPLR
/EK8CNV6ZUI1tTkqw/PeHUMYabzkV5dkSE8Oks5bmNapA5fwIO7FTX5ykSXpyibI
XCLvdLXS8/nbW3Qme7XZSCtLDlrKWMSG6gev7LFqEifCKoo/CLrR5qObwYW/EY8I
y2atQeYkOFhLVkylV1qUdM0V+YcHKKrcUlvm7xLRXmwWh9ZuF+mzdPnSriDeH2/g
etF7ZoLvobkvdDNfXFZW37l7z4b9rQgJx6uS/lLv77jzbxdEQW0EEgoSTli9a/Ve
5VvxcTILvEXqYbrqNPFPTfiMWmqKjbxbF3S3CnVgqacIOFx4Fa1JmmlGU2/I/l5s
umpKX9BmNqCFPz6VOCgqv1H1+5mKechZNlSnZA/CzoFyGXhnE7AHJp43fEYSxfTu
DwCrNlpDXfwaZmcjt+9/WOKh5P3lYuKEmqXdYRx74/fy1l9l3BHvUc9ZH7NWo41j
PFd8Y25I6zKYhfXciCzbtEPUr1V6+UmHd/hADHe11BSFTu4xghZjLzXiXaCCEI9m
U2wKr+uH49ghbJvVyJt3wsK8kX3zBn6lsO5jonfyKhlRinCsqeOZkRxjK9TTWwiv
slYw5QzEcO3PMf4ETab9Xa9hDeX1EVNFwnQl9XNaX67AP/PAiRLYayMSORyMtect
uNWz0aHXOsOgucms7zRdbLBb2NuVqDA2nngN9/z9dPIUSQ/8fBALRnKr1Wj/XVKv
qjDmQ3fjkp53rFpgu3XAfGJDYZl97z9O/8sHvaR+R3HSD7jjG3h1zF0/TQIHAtiF
gQE6UI0cGOn82gQiRd1E0Xi8lqDW+GV2Scv7heZZ68BhCPtpLkIKPTwcKs3tv1VB
1K8YSHvysOO2syBiWcJDr/o/Neo3ZijIUShW0yzn+Fisuu3Dk/IxBPBuxk+irigG
r9v+9R9Ixg0mbpo9Wri9Dou2si1agWxej++dEqpr2JXMa3RgM0n5mxJEvMPHdmgi
fj2FQYRui5NK/qsOPK8y/lCofDroLcLGP9C2yQReEsJz6B96ylDZwT0/6NAKJrWA
xrUie0DlJ4/WWAHWsYziy7i2BDTBTg0HqrqUubb55vKHIvLuSjs7DZukH5oesUj7
KABmNBYo1Js1ZEHiKFEpZTvvCg1gYHGAZA4Ek8TznIvDr51QoOwgOmem0mv6FuBL
WVgJAiNdYWad6VuClAnteT3yUUtzFfUR4LROLUaQjHul7DcxayJuD6Ik1DGQXzTb
CAydnFdgfWHaX10WxW4o3qe8S6/3MrtPy+6LiF+jkIbO8O61HIRyApe6WLu+O60X
PKPZHYSKwcASK0+DfpAnI3Fdm6aLk1QVAGGX2+//Ewv2l9MHioOBD6VOJDpehcDX
0BRdDlKU11ql5CmjlddWPwf6XZbnScCp+Nf0K6xaAArYpgjJkXZodvGCBmu5qWPi
RrJ1rJ0nfY0LtEmflPqf+0L0eWfouye+etj1FB5cu+iWcP1C0x13Sv3yn3QMVqWo
GwDxoyoe4Yb40kZdnqQLrezBsRvhqfWc6bWfVdMwyOOoHxEv61D2YzbfrBcxgDmL
FXn5hUQp/MFC9A+8uKkCjvTbEb7TCFkoonmqo4Oy7dN7S/KUndnw3dzYoNPZSx0R
qk0/iVDsl+RWcLaY1se4HRgxLc3obtkwvrZatB/2MkdM9Ah3Yf/60a7TqyCU9WKA
jFqNDcg0drYVj4Gwzu86ZIl4t21llsikia8K+KY4dhJL7bpyLKjkHavIRwqBzmdr
b6yMYQa7JQRldFdyUjMU3bpgk0Q4OEqKGiCmzn/E1+udJzv/wbtCjSZyTBiKQd0D
TIdkUAwdbsvIe2QpQpjpzFsw3vpBEFmctak68zBKMCgx19AkqGIXaUMJ93bPSYQg
eSjmqOqZ2uJAAN/Xa9ZjpiyCz4Cr5XfywYFyCHrBi1uhX9Fq1WMVypH55FX0JnqE
AdyeCDASzd/XqNq2lu5Z+p1huiW953RUpWiGJwAwsfIqFZxc2zfVZWZB/3Wp2MO8
LGIJml7M9DtmgwxIQGtjV8q7gpdjzuLjuGTSAQyAhiphQm88GbrcJRYYF7eZIsC2
t4DY+LOeWUX+o7KUvPMwO9JossSZjUnL/b58HEBfAz5swfqum7nSkaZPjZ+10ES6
ehEjbDbB1VngahHHofkDvzh/HvgYEYoYHEsGancXxEyOCsKFVQMW7GlVqmss35rt
wChjCbykajiiG9+7MksigxJ+SapXRr7V934QINdYzF8kWrNoZzAUie/25kH6Z2Ne
ppHvEuwznAFDqnes7pI9qCVTuVEGciX7GyaTHkaySFP5FhS34XYxc9K45Qw1iNQ9
BElKVHXqTJhw5evCzsxzKeD5fuiC5SNH1QdfQSY8knLX7XrkZPqt5s1V2M4e1tki
x3gGcyMF9URjWK1tR3eLGcO+6QjD5Q+xheonCZwnZnzK8x1NlYCYi6lbNRlqWExL
bqxmXHeo2K5i8VRqdRZg6DmpTyoWEvY2/4Y0nPy1+ma67Qbo6Hexkq7iD8wEgqEP
byjnD84TIrXqStwUX//2LaCzkN0NbWqkjgcVoIDwePo9PyNpCiR1dEHZDB66CTsz
pnNnEJHXTmzMPOMktnwTd7qUBIkjb3FtWJ7rAPlgE1ZU2rT0xX6lCz2YLESUHdtr
Gv5Y4Mb/GikkjE7O9UX7usT8p8sTix1mtI9groeIFAnPtW9hB+RTOFu3ARFu/jpw
/pK6ARwn9okljNJssT29DyfE2XIMqDD4aViHf+23qK+i+Ph64pfoK41e480Dg7Mh
mlEKwBwL2G7BXRwsvYU/RrhThRYNgY9u+RgYOzpWdgq2Ek7ORSOBCfL8c+Hbi2LH
BLMQFw1cq36uBLY5hzo/bxBB8F1jiNQXI9K9KaCMh234b1AQ8qpQw0++nu+i2dgT
vvfW3+c3oLPJ5gkoz8pB60R/yPnc7d8HJ0g42G7PGZ/OXXGq/BUnt9yxBCwGeWQP
VO0RgVF4UJYg7uxs4jQG8SbP09pxmdrZW1kwTnTrwNxWNrBd7+xVC4V91uypdm76
pSY3r4xggmH+Wf3QkEkhYaxxQlFeqWTKtjmeoYVecQtHvgzTU1vRQcg90AGHxGIV
McV+JtBw9OhGXvzuXGd6IX60KZoIxzwSVuRUoSlSUsUg/6lpdvMPEDgBErW5TqgB
/8cTvr9flKvgBnaU1ZycOpnaDkSDCZthOtnHQkswosjGB1Yx8dMxxkwv5xNBH3Uv
vPas0llY1Z4WnNHavdOQrdSggvkiNLDdEzkeeHmmaCN/TA9GoF3141bItdJ89CVG
5BpY/C5c7QhxOBMUOswSH8WIzK//J7ahkAHXvOKZD9kAAuE+46Ot7Hz+fqUrMdod
xBEQgPU4puFIXQqxpPsHXMEUZonsqZ0jCfeUqgEp+DtzyBTLBr0NyNeX2rPUgwFD
HM/NjZIEYqu4MpE2ZAO+DSIAYDgULWC6Ys5OIkXcb2zi3YCndadjKdOSmgo3p5hh
/DA2YpVG3gadvS/jiTqsqIA5NgSOjA3ldrjk8b3xuwhH+ADd1X7ggZ+BcpayXCdm
A9db0Y7+QO2nWpYD8mEyyyybf0nVraF0/AGoszyB+4EkIRThBSqf5Mu95CzqYaJP
WLhyyVjFGDqVoKe5yKHezwxKsYd/I7bL89BVXuW6KLsI0SDyM1cRvLxHsWDrc0ya
OrEIRPdJ136uvEV6/a5Lq9FRRTUDz9owA8ktz3UYbxtYRmhOcKmUx9lfr6mwKNXz
s/WQT950TKKY3y0Cs7gTsWkMfq3kMaMcEoFFKb0mEsf8CeDHt/sdik0JlUM7R+6o
VeOBBm9jUngElfeMjUGd8PBAOiZoQtzLDAOU3HPOuX8u1Jfw2Oi/x/4dz/l06e1Z
OM/p1E120gcLl4fNhCNg/ANkJO3fihMm8nN9KWVjXE6DdNdeCbkjI4YSSwolY5cJ
ooJ9TJtBo0UlJXWoaqsnaqEZ0bP+mnbbof75jbRzttceAsmtn9PlMy6ZaT5SBwfO
27yJRjkUOPYrRmXY1nXi2ATOs4Pby2qSlYzyOBpeD2tNNenmAF9bKPqVLjuOqq7s
EEWN5D+pUPTWiVA8JZ9piI9F7qZBLQwo8MsPG8YJkTys3b+k0iTMxaS1HJ2us+HZ
AHlOW9qqcKvu87enGSwfjYoNoGgdbveEDoYmxoMflWEMBT4fPA/ShBFFkAbxEBsc
iHaEv/m262oWlyhAlGm95lx0tI99lbOLBOpsDuHf19dIJhHG0uDXDVAPJ9LbKQbc
g/85AhL5a0+JX1Wu7RAZtbRR7U2kiHGNWY5PkCLNxylo9g7fDKYvCgjHDyKwN3Qc
xeNuD7+AfcwVYO+zY+n4S1eETHrVsn7kQPVDETOQJZ1CGIYaj2vyOj69uaPd5eSi
KO1pcxqKFcOQq6ieYJeG7Sd0Lm8tH+5mrcNoaUU5pNd/rkB2OcJ9a/3PXAva2pRC
oodCJ3tZeQUe6td/3eg54rBaKJz1M4KXH+h8F0VkUki9MrrvdXXJyMuWrv6ydnUH
GhTm6rR257AhLi28mKkmfhb2jSelVtZDVOHfhLxupmgiW8+5hVVbtstilwfWNTOY
HGzDEQYjleop/sVNZuUcgCBJOO/MSLmYYuwEbsQW7y5CUGYs0oUYlIEZBKVPxGpz
uCHcBE72ueCfGnetpiY42MrXZOCsEPD4QwyBtZ/OHzk19fSxVRTYLrB2y7qq/EJT
VK99CNL887ZRzNqAVtoG/fLTlfjSHe4wrNGnEnQDVbNU6NeIwpwf8Yowp4hZGvw+
kiyaD9SefiSoyecUeZMUKilD8Mv5MEZeUKOpXm55xQorTnFnp3sMFvXOtWbDWCs3
33bJC40nYXAHKPLoQUKV5evubOI96COQ8Yz5zgCDVPHWQtdQ6kjW/9ZTppHN+Adk
aPRhVzQ3bab5BHVvUfcmnMX90lbY8B6xzTxZenqn0iH4G19g7bWwqLSD5ZljVWF+
UImjTx33/fb97dFE0jpkiXBZTqTo3grgCnCrKLf9Kvc4PAMlwxn7Cd9gzoeDmFbQ
F8qzUoeGSr/oYsWLDIxR+AMKJ0tFoS15Yv5zKmbtTrbUXqeLcQMP83nMFeIjkD/L
ikGnM+K/GT/IfO+RL8QebKoNby7daUhqwnSjFNLDjCW2yJ29zeiEAj8whzLvNYZ0
GrgKgpDkdf4VwwK9N5dSg1HKlzK2Y0ws0juYen03Bjp2+pPK0H7gkA6cbzgtnKLr
sIgIKXdZXSkcFvW7Opz2sJ+qqXFWAky/gIUr8YaRSjHQ2Hs9JGSFgFeSTGlUNJk0
JF40pDeJdcuVf7rerYrhgBTTx/R5HkUYzlMDX1ydaVZ/NOt+5aruo8kPruTacYEk
w1OL1lZMLj2C2oxo+vhyhkk9GKyvrqSRHA120lEp91KuGNxT+zCfnyKlEBlUIek7
Qti3evDo4r3AcmqF91TRhd417oWHEN+CGHTrXCgw1LQDC734+fSF1QipYBEuCbd5
7DtXZfR//b5OYhKaSk69qSF5YDV2vGj1xYhj0ow3+ImkUbw2dmMajL/TfuOx0WdO
V1FTHS3Re6FGRVN/KZkVDNWp3tLmV9sfzU+2frk9uOYLkiFNulkSivx+zLqMJeUd
4PN20G9ylCTQtdKjDu8OjcRDL6JANqGnMEkh1trgDVFHEFY1NS7nuzzeyIWuqqrp
qjECpltp2+TudVlt1AWwCssAMbqdfkL3nzvQyRUtOdpzvf4qMh987pcJ5zu43qfs
Ft6GCNe/Cd1nMiKXxVTR3TRLPDhOp8Qnszx8h10k03DFVgyl8XmSTzzuV/zM9m6Q
ndkoVYqPSd+JXB7xSfE3MrvuJh5wL5MjdkHMAHDd/On41adsr3YDVfNzFeql1eaO
ZQ3aaTZsWyJTZxDWwJ9UHe5uT+9X2PnB19Y8uQ0A52Z1c6peJsre0iaqBQRLfXH1
54WlhHZjEsr5x+J+rKTjzOZu0ERoCJRwUUwTynWVStXAQOT3zBY8cmepuqg6rrCv
1cb5Peg+hdZgF5Hyar3SOxplX0No5DnxSzzRFD9yXJascOGRky7xm3cTEaYcdJg0
TylmZLVJP2AVvEPOCY2IMq7LhogpBiqMfLHdLOa+MwxvckDtPGcMamZI/cijp3eW
D6vax4btwi1uYvB4SLm+vHduc5tT8ogL7sh8rh8F6RWO/jKpniS4qiZE/vRPklT5
hF6jyYQsHluiAb6n00TIRRNNP4qRwT48qJcHTE7a4pkdT7RDAo7Baq5/KDU7tAuM
wQGI8DJrpq4GG1JLGFB0+eVkiP7ddu/SPmgFoM5/DK1WSc1PuvT4N3g84D/aOZFf
nC5zU7iwvcolkMTVzcs5Cp1Yl4ib4hw+XQVunZVdT3obuJBxyc1MMdXvx9ph7buK
Dxh9JWQj36dKans7FebTz9a5ZlNos3/SXhSpPCUmjd323yzkQTVTNePsYy7IHHYA
Lo5DZ3VtgyO3aGnSs0pslnBYUXr0W2b9JRoZ6j2oMRZJGF5aPO+UAMFrGYw6hjyF
55iqDHLzeMSvUpE1ce15qZveiDO6mFq/rbd5/tZQvtxlU8uf1uco5iHrFZjgpFkY
0Ztcuu/Y1B352g8Y7RxpMn4qLwapIa6TInoBb0iIJbdXnTiAB8p2U1BKGs7Q+9QC
NwdMTxocNKdgtSVqhQDaa7+i0eQ6m/ngh7TZG9239ebI4d3THaWXNgQ1TqQPJdBx
IQT+C/cadSD0AsJT4W9yubky2+MEqla95PWTH5BSJ48eE61ICj2aLj5CnnNIm9LA
qNreVkjGGKeRzz+N3nHeRWFGf45WWvqu7iHqgkj+ny9WKjrSUEzzgseasJ9H3Zi7
TA6wc2NhVS5Fqn4UDW3B5zoQuh9hFUT0CQYkJR2T63xYUEkiFIHCskBbGD63UgBf
paA4P7f/7HffYvudIWNqC0mBggPN0atAuJSoBZPFmU04TiKoEbPFDrjZFre1ZbIw
PL8IKF/VUxEBxVZcp/QW9bL7d44Yneo+pLdBBHnTLTECQTO/LvcCg1E0E/4VTCg9
1S8ZX3+/F9XR+ixK/BudjNtG4mHx7N7qi26gxfvKa7SFL0TuXTrX/CtlffZVRwid
qdYBtZ/BsFIyP9ukxGVatDimk8TUd8SiNrbx1k/WXBoQaYH6ivsmvgrEmbV2SdYw
KpDcqUh3HJcoiG4X9GTDQ0s5zE02mYN4CJfc1eaEZ2GtvUCOoNlaDLLzkO+5TINx
ghiTZn8LzP+lfgLQDwhmh1AMpAmgSvhdEWmpseKnyEUKKUWRwUZbpX64mNVG9hTS
V/ndaE6CiIE0lMKvN/jNiNKgTg3374w5Js5+pd5i48Wf/vLOTXpRSeWANJB4P1gT
osCZqvnahx6Ue5dfDWrqyOhSyHvxAntt82Rq9lATymngD/pF4YCPvgP8zgW/VRpf
8vKYogWVtJvV44cZKokvjYauYnwrPgsR9FjYkTcrz/oMLPPyXsOwUX2tpH+DmHvz
yT7gCBH12/RqA13OUOkwzHxChLGgDg3zhKE4JK8ArLbFcqfNdzBw4v2ETR6SEfte
DqoIXco/8e4i6MIDJ2iuaIZO82ndixPdcqkvpB5JQZ/Vmd0UFZ2RL5Cd/wFO83JT
spg8zgGfrp/R+2KsNsZcQKZm2oiWZ2MzOe9JZ+bErNyeE2Zaa2M2g6f/FmkDXCsF
SupWa8g1oP8ScnrrtKM/r/V7dd6bZZDlLQaiJ91ujim8RXLadcpTszdKILspukvZ
p/LI0X9Kyy1aHpsyPfR19OM6bXhktYnO+qbg3L+LWY1tOgQ13KI5m6H0DKJulFIm
F37sPJWYkW7tXidboBPObVF0s2XM7i4svRgLT8b24yZJfq80iX/LtkIhsLh1Ovpc
NGiliYNKTdUSompvE1541DBcNhLZS39OeynG0TyawCi1cuGiEzqsw2XEUTo5+Nir
JvHaSAzdA24b+ZGlXRseMG9poej1Dsxb0/C9lF7pNFrJp7hbi8OVXm5RtE5tlfc6
rqVDBQKMRf8/KhsnOjAitiOAFpsBdGl+w/RNoFfWHQ/tWnLqssDx7STvvLmGiNbD
sHoD4lMU589xK7WtNgDq8BWyG/zWl3yHIiNw34CcaxBRGrtZw9XRZICq7+Igo6tw
ZL4Zd8B1kHNSPUWsmpQIVBafB9Ga2xHOZnk94FAZ39nMIDRwY1kSBwGb9l9dmCmA
9UzYBZVOOL/Vtw6yHvufeKDCOM1VrV/Aq2qHF7Z6WuhQWr2CQi8VpS00y94ubgX9
DbhAdsZNXPLEMZCcEi8mfmt0dn6TWoa9ub8hC99Rqf1GU4N/xjWWehFuNhav9t44
5aVs9mtvObqeZLJvE6mZH7TJR66Vf+niJsMcQDB4wAtL7TZWaWIBSgjsVsdG67U9
3Uq0aOdcPFMf1dRPQ6aCgpEJdvdExruVGvzaoj1lpPHsS9j1R+lFEiTxlRTUwnKB
liBUX+H+5l5dBvOl2vA2vvTm/3t3Zjv+ITzTU3/peyPxvl62gaJpHzhJnxI4ZXlH
qmi2EYjrs6R+6C782JcXyOlGJw2fWpDRmRuLziiUFyJUHuZcTlDXWoH+UfMIl14a
zAKbZX30Md6PDffNXFdOfUZoTOYA4YDOLOiZbGcy3hXCIKBrjuHq1jStQMY+Zqc1
CpiCdB8n+G5CYRdNgGi16ss1SJmIoJmB03ni6eYuApSr8yCZT5fKu6FV9HowYJ49
BbT3MybJX4fqp5NWmKG5fglXKigBLNRWVoQhkLJ/mYozNW5I19EVAnfzGhg2bqLr
uCU+y82E8DE8HDVqcJz8fmlP/I0aiJA5favaLUZa2soKYllK1m01XQNZDBAOWg6g
HS8eGQEm9mOttSxHYwMMTAx+u25m6GvC+4SZpkKatHymb4rwD8/FvWYNVq0Z55bE
9c6Js4M7UrdbkNyo2dQDsJKzpHg/WGXwNrmlsjf7FxotCbwnA4QKtjRBj4Tjzkra
P3Abj1dmWQy8MaARzEjcdf/SzKYrIEj8qVOq+pJi4/H4CGg3PJvn9wt/ZjbNB5fn
sMw3uGIxlT+WyseHH0KNZLyzxqxiYxV92ioqvyVdyFOm+DAt20OHVn/BGErrNUUn
EknU4l8EJE7L7611NJTi7ryKeKZAOjbyomU+6TE55bl+g2GioivHMS15R6FEU8x6
PnQv830PVCF01COUzRupTSHwUYv0CpiAgvFr27cD37jqYvIDMpGIfrUgrXbwWwJb
tNwN0z7KTwwCQxtZfYkYViOfoBE+3cMp0+6gBifF6XEUMrER65SiZE8pn+l+Dche
YuWshyNGmetHU6YBD8NG7k1pz5KnOcX/2J1M4kFf3mINCtbu7st99fH12klHNwCq
/7wC31oT5fgIdEQuA2D9xnbB9RY7GJBW7HAM19lW58zKy85fkbgwoz+wQpkgpbwH
71AguF2q8T3ct5q1XFOnKP9gHJL00StYWWhHpx53fP2Tu+Hm+0AIs8sJyzH5SLuF
+JnMsMkGbnhFDuCC0KDg+0gfe9ieE0CwL4hQK4jbkRcDpnIcKK0a42pAa+hUl7K7
659UZ2yYNRejA6bE3QAHKSUXlDsJZdJlw3NcJbBJMtFDa+OLuvrk+GD6F1Gd2t72
/RecKse1ci7rS+lLm1eXdW9QU1XDX8YQHlVwP4MvrmimHgdn8SEz5SC0PZRccQT/
XNdG8Hlr2vMG7ZEXFgHbJij8Ge/Yq2IHTdesQE+ldxfOm8Sj2anAB6EmCdCeHJQg
p+yXkWTc1dtN8/oLVTp3gRT6hVp8+su6WAb1cr8LmQbRmMHrYR+zSwzwq0roGV3H
iNdQETrO4z5GMOTxytTMC+VP0OztJIwOg85af1UjeuzWYl0+zqLbeLJXJCnwPf8k
C6rbgxhn4y12aOqyD6kvl/ETAa0cAJORHuddnulKrEHGAoWynPq8YaXw7t+ozHq1
JjBLxlfZ6GqeKyqMzOt6klzr0WDw2aMqb0zX3ZuYHcR4s5XHpRVZSAFR4Z+VfRP2
LYsSm6K/omXpf6kYlPFbkY+f+IQAUf4tXoYOpna3VzzzU1t9aXxJqH9jx3Sh7L7M
zynuSwlEJgJANM1QlV2TjyxD8ligQAg4GRJR37nWnz+uyQNKAqJ4RXuHbDA4o96G
E5VTuKTxFtGAi0U7gsIf85+UcKhYOfQRdDaN/UYuF/8TOiuOexD0ncaCXHuCb7Q+
Y47VUVU3B5iVpXJf/r4uTgHVBqbR2516ygmV7TfCIxWYmQs/SgslhfzFDHy6b2Me
csGaOBxylYoXcYvsXQDa6hsQZabNyZh6M9ZWDzWnX6KuvPVMKANSVLoyfoX1ZPVx
SbrkldFgkH5xWuuemY0L70utW01A0m7X7LMsRxizRfK0Pn9QWP+W9mr1TMM+WdUt
qyuhYIeeh+QW7MtoGs6eHFTd7XmcGb7L9dCUk4DCGSnA5FJWlkCu+abf/tCM/lGw
2fHlh/FEl4e/Snt/E9idlQ8i9a06/LPHsk6duq1ppE/N/mZvbzSo13ILj3rGWGR+
7+jIDUDQ5NgWJ9xhcopR6ipQtpV/yGMfHRHyh+6Y4xazjA8Rw3tZuDR/3iNBYccD
YJXVWYRLSELSYakFNMNqQQa4ZisnMqSaiwibhERmO65v99cw3NoQM7D2Pg10ukA3
sfaPXJ1ciXWJ+s52VdQk3DMwq1IQ8py21zNRp/rcvMGZzcfzm//mOCpkZCqDFlDx
8A0Fsgx6ue4f+61eyYhkoVxDR756QuwUb4gqcAIme+IcQ9p4amPBuGKXpV3+Bt+w
YjNVnKkXgXNdlkF408ddETS7JmmT7wDPR8JEkmpY7JCi1pm3g6ThVNvmbjsl//ES
puNchhsVshnqE+VY6s0oo9JxDn46f2lILZqvB5KktrRQRZYm9XWgT01xmroLfQ3T
zcq5Rq/FPTJyksDSKXtiCOzzh6zwdMuCAZz1A40B/TDI+GXkwRQQJbsDWrmqSr8G
eo3298GB1NoSxTX0CBdSf/5Oh3zVPKApWRv1VZvWkJNmM3fzm3w2KHkawZ6oxUEy
HAKtmHvE5Nmel3B9SiMNIAEZII8NVjT4rHkWOiGO+JK3UD/h6KzZ10GZr/WWnwAk
VhHr+6Qd4qeavsmR3MjcQu5CBjW1drOkEgmfAMAymxQmB4RqOxl5q209ngEwturf
UAjImOSO3jkOgMARMKTwZwvlYrdVgQOw+gICgDWZQWu7bu7y+/10W4M+2VAhpXCG
k4TYDVovwcjtII2Q5YHHcDt+jvnvDVZX7qMPrqwKpHi+toEaa3lEEBPC65ReX5ae
hIxFuILA9iMPHHMRfazxzsSL8zJnY5W7eKkPLzlZC9KWdnY8bIbzg5B5oLXuK0iy
JhU6gZl+W+U5vCH08oAs+30TH4KaGVHEjB5ZOvjBf6TdFUYyoZMdF7DOyiwZElmV
6FzmWVHKOUCmWxCJJOL94Tv6xo6sZO+IvNxBYFVvfM7LkXZNtAVb1A2Qg+VxYvT+
yKNAEYTlvp7eD6UKRaj5i0eb6Gf7ImrQNzTg4iFe6xTFd7AtGCmneCHWunjcac9d
jd0iC60YFkYqBwkMz1FIsjGobXylOd8FpE5GSnFJ0aeHZLu+xblsk8Fy7mQuG6B6
jTz384W9K5n2hKbGx5ymoLZzNQ09ZF2c/x+Ua5NOZHCMbejOTOEkZzMOe1w66Auj
73Figpc4Vekiquy+2IH2vkIgn8njPcMSVJAiTq/SwmFTA9+eA9VWE+4Sb3XGeoyH
LYrHGL4KCNlaZ74x0bTH7Z+nykhSVPRABE624Z7IdcspKxcH/qG102UyczXTqYvI
AlTP1fqGmX/0u2kmnJ/HAYXO8NQdus4RFcqgjL+KgDhmmK1Kuuk23XdvB1GWntxl
Qzvn5cDpRwBvOBAIjJD2bDwUw0k9UeBft6tThHtSargYvyX0VAMJEUJ1E9Ay6oZv
JXTtEOC3cVEhbQ91bOtG+I2XpQRRFWCxLL9bRoFnfySSRgkO9B4ydjrAFjg1hQDy
Uc07r82ndG48GJTaBkgeMTMJqf0qpsSFrr4ICV3AoKgp6KA3U4KLF1uIZEDd+DpY
V60Fw1D+GVxPuZDlxfKySq2M+J0c0iYGnPGJPYTqSEKCtw3us+th9nUPxEqz/5+o
ngy1DyDgkYEs41bwB+TfRogTHAGD5jWl5NuCuo5LPeYijU0boLMnE2tPIU2Q3oqo
kstBgiQ2sphr3O4K9jNPZ+q+zMuUwzLKdHBopj+IeUGSc2AWrDnCb9Azc2YB2xSs
4POjybGOwaZIpYZtQb/216mLHD4EeDnuEy28MSagjhjIOF5r3pZfiAbJ0er/7sd2
wNYUk8hCZoNQX/21EUp+1d6aN5CFLu8x8gniO/kq1QwyvXG/d+2wHpQH746bjKJm
7pJI3DKzSa5Hk+HLIZhKO6iCG9vZpxdsqTfHoCGY9tEIxSbeoUqmHd35uXOCtXzJ
OFqkcCOXJFi/9pf4Luh3Xn+dPJ1DdoD0LqHjHVgOvcrNK0vUZp1St+Kl63pKVSw1
aQzajwQMM9LMMKUZws31NlmNqyiIlYpdaySf9xHcatteBTv6CazqtHhvitHWVNdr
bONC7oSmkWwJz/REwbRvBeys3cb6xJ94fwULRskL9xc6l8g8BvMt9nztjyEnVUr0
I+VYX2v0hsQAr7IKbjqgaPeIdnmmUCvrYK1XfSeoTDBEz3HAomlliRVXwUFbOUZC
qoMIWD5aof5/ZaByXQ4FFxXbtGw0iViz0NP0rua30DhmTCjdp0TNx7pxBLzVjUT2
WxU3rbDPxieWiHns2jTcwdkM5n0ZTQbMIb2masu/+39/cFPc3ACOdDmeO7YSySEi
uKocVwOxJJe81ZALTMx+lf4VioZiKvtMAmkmeWeFqslRpHxwpUw+p3HuHoPIrTDD
YlQsIF9uvvx3Lrak5j+RWJiRBKYAw2Fcoy+0zSOoI2asuiUzBZwYhTLa/S5fjpMQ
9Wqvr0Jmr507Vww5BlDkeSWkainE/DMOZSF7PNZgS9joF/SOxDfnjlkZRrAzVOJS
afngQ1PnkQx5R8MZ9LcaT4OJCAbHuDa7N5/PKgzXy1QtoflqUL1w11pQPfHvmlL+
1F/ba4Mzs1+JVqsReFhXbaQIAGfG9ukq68BJMZfhQb5zconP4VFLiszz2hndmNsL
xttFrRla7Vv7XVQHghzLVxZ2Q9n0L3tDIbkXgehlkjyfkMW4oKGAFa6xiQ/j9XQ2
Ih6W5mnbplArLWRuKBDmMrrMtibF0A4RSJfgipbyk71moiM816EpZdXeJ2eaaiqF
IcUr58Uv1F30idOKZElWgZsb2qj3xcAzv5fP3HSX2l5AjHIoqxT/HxH3dEZHI8kW
B0tvgJEaLSMfca44L+rHN6TCmacDDnk5G/lcLDtB0i7uynLNvV0NQsL9WDzh0CvQ
mpeTuY48kBFFPILB4e7pmtVakXZSw4/458DfdFM0WIzbsazKf68Kz/Cbu3Z4iTF4
JkGwVywEz8iBH2K0fVewMgmiq9PLLKUqe0S8VJCqyOUzTEIZR+c76i5p4T4o5E50
0m5YOhf/TuTvqjcSwXl6H2za8ryKMKhaUKb+uq2VDVa3lk78Nkwb7X4rysa3KPX/
8hfno2ifE9yXUUkDKYBIaT+bV4eqgfEZ/YFLhQsLjorCAJuqj3Q5ixFrk6k1OsAk
/L6Wrn2K0QUZ1jpbR/rqCbObHgxwwzepkuJsuFEl3mLfLFZzP695zOLDFW/2leUT
J+mWKEaRxQf9AgBAeD3qTUGJMDH4f2z9KNGlpDnSt6VK30kK1aZs5l81xe6oJtGX
T5mB9wDj1YhFKQsn1m1aJSRdn2uKdEvEXUE4nAaVzU/8wbKF2R7r3MNrsEqFYFSK
kOopKJKkkKJRZKGpHa+nBeOG124Lm8K3yVtWfPHBVBzUV3bbTijnb2qQVixa+RvV
jgagC5queRWtrhBbF55IXGqZuj4pNlFBPZb2jmFgbXgypiB7cgBw5t8Q9EHfQl/k
xn3arqMaYestDH1iq0KcOYNQaQPYY9p8HB+oTIhRvP15cjsvtcQQa22ZGBGFLDGL
bCoYc6wp0rrUlxLSftPlquOPlvkgc9cuzBXFJXfr67paS3KxB/d/+Ic/q5FWDs+4
m+O9z7UWO5prS0bsSqyDns3mbGUpC4dSNf39M5Jl/AV04HDsN4Ptw8s+9P37dOx4
6bixI/IfYOTF/3Jh7fv8L7sIQ/oQNNkk2y7ytKg88/G3KtuuUnkk04xjJap3K8fk
qhAa1NxpkisXqB6XsKYGBVSTvrFDYEAtcJjZO7aK3smEHga6aRDP5Ehcukhhk4D/
sCPy5/qmpeSxK6SZsE9Usiwrnjr+Qy8uAqGu1M4DrV97gcPVl1nkZFIVCW9CScqi
sGVBOX7OQpJuOQRxjdNMQGIIA88N6D17PbzbfkcJ6+BX69Ty0KOIODwYhHrmMnGk
f6SgAOxhSCKWRDVbX7Eq1WqkoVLBd5keXt//Z0HjHsJaZbE9wa19xpIYZBL7yBFy
Gul2VkQS22rX1DMt0fYI+T+fwfIlfuKVnJ7IVb9oMfb2z4hJlC5Y99anSODN6NZ6
XmIK1l8mAyIJ/m87NquXD4Fbu10NLnDQppBnh6IIrlZm/M2e3AWsiXG6Jgm/VJwe
g06ET/lu1LUAK1snHiRO/Wy91E1oCxUg2ELKjQ7PLBHmDa7bOZBjFsRe0kDLMCN8
dOWeBansIi1ChEJYq2sf5KMTDgvBak0BZSrUbCEJawcjMNraD1iArtkONIZJXJJe
lvkZm8TRNwfLUhoa835tV9vvGe96P63cYIyrTXp1ZkXlCSONfBCq1DRREMRXbMzE
PpXQnmEYZcJO5TOFhzqTEkgN8mzV1ljYJbv6Diy6UtJ24jok0i23lWxS+20DD8EL
SiLtl7YN0lBgvi9Lt5oXF2mPzvdJBwGYGkI/SKopuieAiWFDalrG5tcDLU+mIUIA
OBOouW9hDfz2TnMKp7++SEWk58zeoYpVxHvJXbIzAJh7z352x1CiIYViD3Cia/HH
1rDSS8UY5WKc6YVBqLqwEukGoaOtHlWipzjp2/Za8Un7zepXTFkMcu7h3b7dpBV9
QV4zZbCNfDVcjVLe2jP/n1BvgUfpPEqe6wCcxGAOZhY040JZucaNtOANMCkXIHE3
P6sURJWU81nFsesg5P1cYCuMxK2DhTEgGePrBqHHnyNPpIrdYGi82KMGiE8s4EOS
dTu46stkm4fxWOMQGNYuFJxpgLm6IFMC4yM48rd2tZesJP33jEcGXbfmJ1d3Yqav
WpH/OHIWEFIuomwyhqTTcSNsLZFpZqhPdQIpkTHA9cUihjAy5Xu8AFg6K0D6ebzP
A9PkJGoOuwTZUujY9/3R+vNS3E1HRLVV93m2dY1bHZSjeLurDn3CDXflJ4K52D4U
cvIRGnV+fTPyYjeWdP3TFgKrMbCQJ724IvK2Xm9KmDUgD71gnRMUBAcwSq6hsAw5
ngJylx9EvMywIYx0ugv/sgiPhy/3UUFmi9QY3r1TeQzZUusrNyWkpraWuGqM2RK0
rdPsM094ks9LKNXfCIWpUOKwnHW682IRVejq/TdaMvVgqzpXII33aadRqKG8Lltk
dH/igQsLPr83CUInZmVmd4Hz2aP1TCHiITVoeoAhVa1EVzHcYw3fVZth5DvhMH2Z
kM6p4TVB+fYXKc6zirOkV5xuASFKu6pwcUiLxb8LDqDch7qpSWWYeSFQTTp8e51k
AoIWChnfAG5xYyEg4dPNsD8ZwLaRfa+G9GV2GabP42wXa5eZeBNr4K/qoFLib464
OBj14raglVMGZFsymS/vgWDoEFi+Q5W465ER+fQ6NcQQUNj/nxPxXWOFDodFyxeQ
ra+Jzaq4hGBcg672YOkPibyKuK057IB0H/7VqeDX1kcc6wRotNTimxiEOXDSKQA8
t/lD9CwNUs+oxAqBTqm95XiQTEWyfmj0AtgQ+1Wqc6oOQOvW5YAPhTy/9RD1ZuaG
et/r0ljXvsK6qg8seHQGODYMRAfj78ZgDBCWyu/wcq1UdT67RIb6wshrww3Sj4aH
VXUlr67IvQbk1OYv0h1gsAec8QiWCC7XPsflILXNWFdWfANth97Fc7H3XORtt5Ti
ywCuqwWan3qUUJpwdHB+waAgAsDLWvmRO2d6/821wc9ucPupDbnkn4EjQgm+jiaw
Ex0NyuDsDqLVJPDFsGW+Vmy9QOOvIbzd/yE/cOdZiqWYiEmbwdA+mXihwUCiW/Qw
84mQ4qxTy3/nMxNPGTiJxgs4/Qjcv0OONprjbYxcyfXmzCN2sJYdoep7GMzZ4UOY
MD1VArSGhfkr5C8nMhjD9/AFVzfVv5XZnR+8UAnS67x1RonbACr0NcQ0zuLmXMWC
f0LYaQcX3cD9FjevMwp7wRQcY065hE+HAlE8VNSSgJIuf1BO0bXtP68g+ZgqwvHc
VoXqxg23FGdfOVeW22C5aOdvpf8vhoQtMyGNgykag2AwJYlQ7wRqXckbvzqmSjIG
DYf66qjMIfT4haolmOAk5DlXThKVvVWMH+aQnpsTRLE1CmdlBcvD+FhQYk/H5Xbi
RhxP/fsTaFzHkiNiIjI8J4K9izjHMCZx+sJ5HGzLmAFhdf8YJWJzaG+Eb1GMcWwO
pDidvWgW8XVPo38/Tiwx/chFOj/I81C/i8NJ2ELmguHICDhFTVfHU0q1wfz1QbsE
ZYOlEGTQpOR4L63bdjkHOSRYsPKt0ytVBXO4pd4pt3mCA2JxPKY+AgLDhocJIxvb
DjrPLNbopMOGyAL4EXWjPq7d1UYHTHW3SqCjyJogcIstSipzR8l7TXDi2N416daJ
vbhCAYUhXtpWQcw3ourjo9J/5wDW43PEGvoDmjDGfZ+7vxZ4g0AwBgIDVNaKYf3t
eAXk0DWCVLCeltHAbKFpjH84HTNHdu7HlHR4vScK6lCFbMqADcR01rqCzEH8Xbi8
6xikAYJCElV3SUkW9KLlSJ7gQw5JoT8QDODcQNeFJmTO8AqPIBX0IsrnlljUGzz7
dNo7hFHVlecGoTsGM+vefOR6xQ57pw8uf61Ga0HTaM00R2TboN5Mjd+TCILa44El
eO0gy6x2zZl5hR1Ta5EON30+tEGD+0t+hNUTEutRpRb0FEb7VD1Pcf4Li1At0Zi6
7zEevZFMMEzuSLfaiyk1USzK7L+8ycn3FmNv069hq/ioALuXn6UcLSzb+uflZ8io
rucCBBDGVshjN+NvJ5hs4kpJ93s3Df8Yb4yRHneOT8Hgt9BV3RY6IZFg/KlE/rof
cz7n6BlMWyb7ZW7C7yT6UUhElAG1WzUZ26rVpaX4X2+chNFAUSbNkpaYQbzEdzOJ
mDB0ZbUhThTwrGu2EIgCelB16fMEh+9PgIu5j3BvXUAeA8kyIKTYhaIEHA6/vwJV
jc/7k+2RDogd2kuWV29oyemwKYul2SacTb5P22WMQbTLorYYlsfSWqBA3D5OCGvA
TeeH+AJG1z17+K9w4wFYnPlieE8+oo1AV21gKFzjKFWRhwsMObKEu/GsTtTj5ke6
J8IXzVjkJLtfngP95z5pvDm+B96vz80GVSZ1ZdPPFdkCT7bu010xFxnSI5qVpH2R
i8oV+LnzlOYN5yWnoUxUsMYEQXcK1wZNPG9HfYpXGB4Fsifj6lQuXnrKhuMiefVN
gZ01DifkBQWX6v752SK+YsDwjS9IC5ROw4Fjty6Vd8jSA1AHIey9iO9f9koodwrr
DRHVpfUxP534G8NuQLkCcQabRnvC0I1y+9P/2OA+wDsW442EjSo9of3SLAAsxDbI
RKbbGsVhRb0twoGECRpC6Vo3zbEmlRKBLaWq6+bRpnIy7G4190rUd974+QsAYAo0
5kZ9axpxSRyc4JNQ8T4EY6HlAyC1Flrx++9hsw1xNqIRc1BmmHwPqEiJlFhDBikf
iPZjKwyvdiY0DdffTTZR6g4R459Xk+rCT7mTeL+BUsLe8674wEwL1oht+N4vcCU3
9JYULNAy5MfqxDDec9PeoX+/tmSJnWgcmjUGD7aZdJBS4sFiQL5ESZ/KwLyezuPJ
9HYKL9jwnF5nS6TWMwMV0rGytloSjsw1gt+kc52hQ5aVCehyQdyv29fjC3im79Rs
Ajz0yvRkgvwgfifcGTcxQJkt0yMiJOPv6dTywxDHPS1KKxW2qWgWDv118f6By8wK
TU1cr0pqPmN7aN+FOpl3dJh8zUuhbd/hgS2ndYay95+EjZVwrSGI9qopXDq6s0pA
6swxVopzVwX7UM9F4le9LAH0mWsg3uZB0GgsOup57+xvBXB3af3PY0SByaku46Aw
39yU12PVswVdUMu9fh+2RAdFURVXzKAKku1PnINk9d84oWgvfoe0Qi/GTUNOUTA4
rRc5Gd5vhe6o3ClVRxUzcWJe3W5rWlM0bxV1daBp7YYY6pN0GiLryynALY36HRdn
HH0dybKtC9b95OHSWQdfKrN1wvDYHhAk6UhDySWotRHnZrVYpl6GwExhSldnwO8a
yMsN3IvrY/eW6b/XuVuMRbamfjdGORgt9zVJoIYBuKcBPn1hKp1rFYE3yNSGJmvw
/09WwblwLpMERki4RFC/lKcR7kqpu1EDUKFqjIlCyOdFKedliPSTRrWqBeymv6Nl
QSI6f2ppsfA4RQYP7HcjhgX3bdxJFAirSujzfF0sMq+KDMi1IsKr+3EDaG38DaWc
DkrmAtXfSOQQLH43MchFjqmiU41qI0VwBvqrJHt5cpMQ1lg6llaKfHhC9SkgNVxu
I9HK6WlvFFYVIH1YG3jJJ8PVjdKRGvWuli0IaVvGKxEEy4nhpDScigPLgavYhysH
+E9mtteofvgPloLbI7MDkp6HFY48ushyitlNzCI8mXrkdSTBTaiLqUcn63UXNjks
ulYLIMK7DXBGIddAxStG5nOuJ7nehau2Vyef8hnOcdznY6xFLmJtMZ7/LAqGSb+b
YuUOweW0GkT6TCIEFTJrCCsQibxJK+muemKNjW7h0KGCM513aVm4mIpZFuA2huR4
5H2RqJ59xKzDZVkC2DW29yo3YiLgzIwePUV4y4ZCoZH6NG8eFXgj302c1RtzD6Q1
DPYpdLVwpIHMIYjIrwLM/ESqjJ2c6CSaBonIMhqjpXZVrVWkFVu0wNimOBkWPEnt
Ewqh9XP94RgDywEiayDuEDzxEJq7+c7acKbECLXCMe1y7AZhTjQYUc1Mlw/FF10B
Zra4Zfz5KWEbgOz8TC+fgb7XgrUbPdMb2KY12EprymFgnS4buzhGTppffGxS7AX+
kO4D8bPcDaTtUMYtx0Rd9Fog3nvX825ZKjtzAJ91Qz1cuzQtp31gEB+hlhT9a/An
kvLiDayGKCECr+dKclCLyIzH57iR8Sv8xqttFrRoeOdcIUpjlS7UJtEwWDOac60K
7D1iK+GgF7sm+lsMcIOvbUGUF6VCzKbZ1TWRVl2iSSn4FXMZ4rYV0VWEhGOAmPhX
i6dJKzMD84rviAGNOe2re6yTiEtr+8woTeBx86o4kycE3lUptOkhcTg8tVgUL+JB
KVeCwmkSjXJM2uuoqc4ERAgs1Yiovkza90mV820ghhukI7xJxlmavpPWtMypAcmF
jjvmAbIUs9qmaiAfr+yJsXZIId5QWtvupMi4CSuCI1ApOEglmk8et4YWzuu4fiyH
Js5eMIvSHKut9F8ejabVBtXLADBNuc8f/x8hUJ9yYXhQ+G/x5/EjBli3ZQICSTFj
JI5chlxzxtcU8VX9DnenS/6AQEJ2nUuFMXC4Vk1zErTVLjVC8u+Ud5mjhcfkKCOS
ckkYpbdYuVYzMTL5I1Vd0KXZjkXaDoonbfBfDTpDpwj3bkDAQtGV2fboMtGCQrWZ
1pkJp37YVMLDw2VzG2TJvU2ZGxI3SCimzXZMkxC8OXH+50Txq39m3GQNmMxsiPPn
+9LjXKH22sdyhMVGmXTx8zWdRDmFbqTZtvMz5fj8WFMwfmCquXZsktBlEa9mNLcK
2Kn8QwEvbOXXTYf1S2sMYhpX1iHMTwvNYeJ9P/wJsXKxgPwqBhGgayKZQ0jTwo9B
ON3xABOc7EeazN+9UlzWdBFLX/LYnFWmsYwYcoPps/kkoC9gU9hm6Gjqf3Nwkhr6
HVg4pQn0fs3rZGenBKZcJ6SJnMXBEpUjWCHwQKIrMv5D9KA6H7mLw5rFtGq/18jX
epRl+GOkN7AQeMtUmS4YOSHA7upDww8b6Vuxci9U+soBac4nYFyGUzeecj67HR3b
/L5CmOoZWHSQVNJug7oyhdCHDxsa17myorfOQtElykl37cyL/KM1ZI1jpP9U1cRc
N0iaePBwl9R+XQ638yluKl8olF98GLnDgzjiMN1KQTTG5upx6R+0Hl77ZizUxwUh
zRV1KTgRaRjtz3qeNANZ8MDLrxb3F67TLUSGhOpx05X7hOGSYliXUid39jiw2zLF
mE3l/Je71nPZ5/W0MbNOwjebOUZ/UbeJvgg6k9uJrjRG14RVI/bA/lcDj7+/vN3y
VihX/1cz2gQ7yFyuRF4P5aM+Ge+qZbVq4XPxJJIhmrVNEKSWGCIhIv7Omn0eVdb6
qpHPR9fozxvbVq6E47wZh6JP+PLMVVAsirgMtimJwcjY7L8t90J9Wv1QVbBPTR1T
ZE6p8urF7wHngpM3joPoq2L3Hl1QbwrB0A/qv8zSGGqAF7RoVtVT0cxr+NuT6SG1
Tj9S7gc4VZ+Fzaxmtg+KQMBwUceeS60TUEQ6NYM1yskZPA45zCvPIQRCpssrZ306
Ln2ZzJtwQDgIh0M4fqPISCbSdeF8duj+E5jsua4HyjO0gaYhhJO/1yL+pIZkhazk
IQooEt8PIXKb3+bZjZSCcm8/P7O0h56qjb7LoU8WlLo8aeB3GGfUcpyeUoM7/jj0
opt4zMjaao8TECtn+UCExTEDWF9wg1ZOachPfr/SGZ2YGEHB36F/vOgTs41RhrYq
eskQFQgS6vvEMPfZzRZjMemjpY+fvoWt95bZqm3lc0TyOKPVjmv6T7j09AbhJlaP
kAY4f3HAK9HNIXsDlp1nKJWz5n5kc3s10JqRqF2nx40jJyo/NaTa2Bxx64ddSC0z
OvT/TIsIwvNq9EHq5YJqwAlpTyeWb7mG3Pj+XW0Wcg4QbOtXZUCgsI6nuT1Sxbyh
pTolJaUDJ/IImtPHQuRITTtT291jktw0e0AcI+bbOOutH4b6KlLHzCG6VhkoD/2S
Hu9JXUsVuWS1NgC4ig71akiH7VjznLrxcJ0L10ZZkLl+dc6n6IBI1hBfZuDQm5IS
q2CNojeSXYSIcG2VXOxQgJDYewZ4LvL5uHrzhL/RwAmEnzgQWkG95LGSjYyA59lt
RYuP3VYxMTcBJ4Wuw32tiKAMpXAZRqJeWKhlwc8K8aX4l++fx4Sz9LyFrrBnxwaI
e1B6GGjC13HBRPXJBnTWBk266Fg+HzzBBFbG6NrRot0FOvydOV85ixBNLePHGRTW
h5Orc4BEBtTaqgLl/l57vqp7aoqI/+rILFhe+y+frKlTpbZY7mWWtT0lGlSSjNzo
St/Q7eeBNEJ658I7z1befhmSy2/b4Gy6wPEJtkl68oV8H0LiV7izEJRVUWJ203pO
FDNmjJeq1PcjNOJRWUwcm3FlrP4ehNZGuaj5PTyHpwnQ9gQhXog21SauseFJBll5
C4UikChplVMAPBC5CmrwlX9hyAOwDUS1kYm96iTqwtc8bGIp1sRNRTu+qC3QQQap
LIkWYQVCv3ZicHscS7kzUfrh9Ev8oQDYTmd/ikKxbpT2vEAytD6KBptxGpN3L0qc
QiEnYIv/rub5Jb5Nk/gfSTt2zDUORalFJkehX+8pyKwn2DD+rEm+fIvGoeRDvcSg
lc4OmNNl+qSD/jAfqGZnXCdmVhBnxKD5qopbYAzfGjllUXwEnpAN+N0hA9sH2/sx
UjcCDjpqGsfQgmr4peo5k0KewC7fgEd5C5H5lkBDOddH+/O0YBIgo2cCtZO+zSss
4ZzMrNl2sKEAsrBoUEpGBUpCkSjPfUv3r0eOjx24hohi53/TifGtLZYt/U2KIJS2
shsh+nwKNS61A8O6SxJXdzl/tE9eu4cF9zRIjb2PBjrKkcBFIkxHvzUtGcffnXVB
mwn6jgava1Bfzbqm5yQJ5wh+R6BWD91nbLp9UF6ABU8L7A+9i5aVgRDBW7dMuBrh
KJeWC79F3jCivZLLtSspP+TrqyjqaPCa1xMwmImAqy0HRAdl8UsNUIiYFcsmvD5j
sPANDHz1NsyflJCMRwXEzU+PE7Oyxe9QDa0o7ZVINdffCHxAYTcWNH10XWCCisE6
WfOpTy7OV7ThsBblWOSf/rMLIYIyCEq7evn1KdYmYG59N38qUc0MZF6fNOpGxGmX
LmlFGLKElCu/yIw/NZhSpUgCbPi0a+NvATKTuhOVQOGun2xiwzWOx5dkAAd5b7pF
15tNgb/Ut38ml8YexVXCfqfk5U3ehWiMtY69RPK65dtVuxKeWp1q13jlaXKloOzE
Ngzg1VHGQGfiaR+Q25sOLpg77Yz32xklQwxOXNI3sKoQl7ZZjwZu87kXEcrnIPMr
xH3gv/PkoBQzd/6A/vYpS2A7udnx4mTsXxXkWJS/Pdd8C7svKMNOtGbqmnYzE2Ot
3+fju8OC6EgPhJYnkSng/CM+JY7zT7qwEc9Az6NkHWb6200u0a+VPRvqpbGuocGC
QFLzxMlmARUafxu/VBOXWHJ+s0kqWC/wOJzrYeHmh6heBp28PppOR7SiThvLLoFk
/t5pxNa6jKCQPx8h2ZMBDhVRtSpFuraUcyNj3iXut8FbKb8yVlqZzIpBo+vLVrkG
fzi/GdnB0jhnylrBQPWscXi1b/KkBNho3f5mddwK5LvTExkiq87kV1Jo507R1vUW
O8qQzlG8pZI87IPyI3pgbUgOyydUF163M3WxIH22VqJ8MRPKDdNgFuuxQk9oCu1z
oeEHbPjwAK+xpkPH8XHzZ/ppMXf2689QTFg+ckmrxWv30gnlbRFzvdLVvU/CZ3Sw
aLrMoJE34jQqcJUt1F3LNky73w4Y3TUOT2KdJKpMsygBkT3d8DW+8qTVVNSjjE3F
dI5OHbGqe+d2uqJIF1nz76UGC8qqY0RcYDHALTbhCLVLbM4rig/cUM6+J1M13av7
hWpdnbPzWaPJsBfrBcsa32oSqnKwjfnBz+2QBtcSMCgfwkZK0R5DUiPgIqHEo7sf
Es62KdbTrlGV/DruZJPv6y2YHtjNBuaznGGlx4bLthOLncm2HhUF+W5I7JpitguS
3QrywDmIP/pcFQCn2C6izkN359QELwj3jhPxRH6RXvawPSHhStjwNAJFBUrsVq4y
95VPnRZ/OD/CBi2mKA6lK0BUNJbzxIHc1EgMqZWa3bCcC/ZYulYs4sXHmUEYnJ9i
a+Z6wnaqFYPgkFsErwtesfp7Wt84aFYX02pgEVQTxHF1dWGEuhJ9j1CU7U+EKjVk
Q4hKyUadr0yJSaKpsO60BDT6wI3thHl3O1iWvSPdGefakY7eG/xUP2nHDYomeeED
sCdbCK5fWy3gdfxq9vjiSGKmXSw1KQfSQ28P0VoNFLp9AK/5RnWBagzu6Zs9Wxyr
hhPFACcPqh/90hUv16yCz9/hhx3220x4qc3LvkAAIYJACc3k9bOihjA7K3sUnD0Y
YDRwcDSRNl394Wl7kuaPmSx1HTUi9zwSISCZOXbwrPzKdBVlbS7/x9N1B+WOG7Hf
xhZEu4mI8YAwydBjuoax564vAWHrJ2ZdGXGwR9luiVIYDPTGw2oeociw8XnxFSWQ
5Oe3+7Zjc7mv2AAG8hPkucxNy8EO/0UYTyfKx0/YLvafcZMaK2Pc3xSLf6s6DvQU
3jzbPj/LCpBV20uzRHrEpcbhNvozRSPH8l9Kwdxhen1YXTLMIF82eihwYo5EihOj
aAFPZyFRcy5yUAprg6Gn51ldJ34XMlu/rrxtWEAYbF7zGwiuYQQrFz3S0lD5ctYA
m2lO1etOJwlUhYi88bv9lOjud4jOoGTQSqbx2zRya12WSwzclogxC/VsbHCeXbHJ
OLkLesKOGk9I653Ckaf/chWNrElaXwpAzz0tvsMUiB36Fc7gzguRlA8m1nSQ3gFf
ekpXhDIVsdu7gqH2xq89YCmqKzd4aJ3j9vMlYto9RD42M1FNX1wZV5kH51SFhteT
R0g4reef9UHpoABSqXrANgWLL4MvnjmKF7sKgpB0bMnmTbrn38savfSdfrBxKmUc
cDwEnmmMNTmC7uhXrHpAfQoUsvYkPV0l0pqA55FtvWSuoCYTO4vFIsJR8zqWpfVX
moxKvDwqwh0yQ1XQVlnglyhw4EUZvkiJomAKP1jwxBtIXlynbQWpNL5qMysNNHgC
LEasrCRp7OrRDiiMPtPEj26gFfz1U1UJQ3EJic2rJuaSEG4MIiwBF34KZxYGJFik
k6Vl3BcTbW2bD4cWNtAnQSA9FRiGqEdYd6bAnauReC0BmUhkRUoPfi7CDLUvoQqI
CzMHpn0Tdn2QmedBr1lPW39S+POLdBMRtB7ZIYwSW1n5h7NnA2Ekfq/iH0S8enWc
+CHFIgs1g4scoEieBOo03QIG764aWReRO2YIQ4MDNjtNaTAHETUC0SMGaZu3PXaZ
FzTFdX7778H9ez6iGVRD3y3tS+kzJ6wgEvERuQhRumT9rGwmoPo/eIUSCP7OnHtX
V1WxHGYZR+7cZgohNcKZMVNxV9Jnnxf8EbivDPV2IY/eNEXGLCaWiNOlCtci2bcJ
Ujrz3qYNMk/MfOnpjoTM/Uq8WyjagbVLNrNhJ3GXCzOvtmV9GMgYbTZmEqJ75Xz0
tgwFoCj4RTe5au5LarOklxyco48zitVcj7fk2hTm1x3Bvf1Om6q+QmQGSrWtpbj3
ZjFjYVl2rURVdBS4pBBabBcbJI5takMFY5uUzmJNBUWznkHfhKqvQLn0R6TekTty
nfLkWlK4jeRpocPSdSlm1vemvTqW9LRAL5QB1g8cMDdDcMNz9Ou5Hse4SxCSk1uH
Tc2++s/x0Ye8K0NYaQptOQnMYmahFPN3JgkV9W/Sz8Rkj502MrLFtnLf9NO+0zo4
aboOlC0U89IsgtgV1O+L/HzFRIqmXpjs1tPTPniF2S3eDgEyUAyqE3Y9LoEd5nki
ECx9CWYyaufg6BL5Kggig687lm2vPftkWkkjD1rEfofxrX12S0ln8OuMlspzgRrr
Q39D9t7/zhC0zcJgBEOcKeiGIc1UxoHuRSr7CyoT8vfnLSD3t6Rpj2sNkXRQs/4m
kAAragLGdUMT2VyHhL8d87pz+1WP7nNJCb2ZrWCs6z1ehr4WRZZxapRpND6kiD3Y
FIu17WaDwkkwFX51BY9/6q029ri4JFDhsemdmVHwaioZEJBv+sKOUai6NMxj8kbL
4C2MubUDpRI5PFMPc/uDOZbAgZEqak6qU76EddzmeVxNeLBkbUCN6CPAaz3PZe2X
cmBkngxJz/IUzCv+0O518x+HLmceYANbuLbE8BCPWK6FLlioDMN5XeFtMhVtL43m
+3hk4MMxX2Jw/EvbdP5ROUelD19TafrsFNM0E7fDaENlFjxe058AT22YEEEt6unl
CEcmMAZqhf1htr5PbqGges/Aaf/NcPJh08551CKlmNIpEwcKiHe7imepdhzrdZ+D
SZ9b9m3vKaUavYLoUpFNYP9dqms+Y+l/bMxuwB2MHsm9fOlY6Ne98yRO6jDjK4CW
x6r2VrkXtyfBnYkrtXvN6plB2wlkEOZ0TACGkPKPFXMD/dnlGheY9elpp3Mwu6zJ
PyJ1jBRrZ280Bc9adnq5NchTDN8+J9AaJf+HIg+azGyIY14gCE1rdkY0VpPBIKd8
JtxdJTzx/GbZyB0FRXehvXVrK19ecjVxJ6BfNIo2MsTr8qSKOiBp4dKgMzEpvG1v
glGXEZmyc1wewVhFclz0iZ0bLW1gUEgKEpHWXiWNLh4q0DuNrfK/08pxLyfa50F5
rEvPwbNu5i9J9EseGAcC+rGH//1KQVLnbUkLcn47M9yf+19AtpnFfLO8SaFIEAfr
qGlXgyh/yyScKsc2o17K8Xzdnwz3jkJTP63jO3WHLrBeVCFV4+SIi3GAgAd5CBVl
ffVyV8qdulkU6lnbnDS4Uhqib2MJZ6bMgw7E6rMgl3Ohelaw07XvKl0mzSCKiKko
TLiEGcc+9c4+dIhb94xBr0kUzHMGUL59eUljpUpkt9iqwCXEI7T88P8NRBQ8y0z2
YFuMbdWuVRJGxgLLeFRpjGdOSnkz4hpJsJwS9+shusse15yG1bz7uBlKdGeeNoP1
KfuwxPbZO95e8qFwHbDKn2C3mBJdAWDgmfz/7Db/rq9ENoyAYvXvoLXgkg/f2UFZ
AyhaOpFkfTXR91ZYavoXpvFimP7OLR+Nxs3nfc16ZM78I+BBMWooqBOykrbg7YyR
UlE3vWC1ohsHmm4YaaubCzRJyLOySv6s+F7WOSJRaAtvzgmcWSRlUKWr0WJec0+K
BYI1bJbs9XIhjPbAqaks3xoEbJJnQajUgVWp0N6l5cyU0bKOmxKwLKUJ+CeKno7e
/2yJ2EErgti5t1tfFP3uV9/u1+wXFgThUlkxszwRfGtNcH054BhIiE1hK7ALqDYW
m9uN3lRBhDBBkFmiutpnJPWB3xcP5MW7IN2zEBI7QkwFDfHfLy0HW1m4gBsVrClW
NcBJoiTs9CqdxJV0mW5aYdIPScsSz5KaV+LVyc3JAt1Vrd5k3Dh+dtSgQsK37FeT
Mzg1Ydaa2vwiM8CGvx3PKxN7FA76s8ZiMt/JwnzbnkTOWg7YL9y2Pg5GT4F6UbMI
g1Q/KPu4stpVUJZv2F3lgDz/eHe8RAUTtt2BxZWpZAhRbnkvrIzYWlT5fWLId3Tq
vB/PG+zTIYD0jkoyste2jQBsaWNS44+YnItFI1x9Je8n1eNF10wJ0RHmhJpA656r
iSWsDgiX+D0hKGaWHeFg/vJ4M8Un6M1I4qDHmFS1N29gjnbUdtOQxBAnq1VwR1Ga
ET5cMNgwxgYePuNM+GMfjIlO4vOUMNh44DdG8gdlsXKm6sMLOwJtB9fdDEbKuF9H
xaj7x3fxP0Ubai3tl3/sspTDdosgoH5IX9izrLeg9uOhRvqDiNax7sK8vLsE/2Md
6DEgPeT+p9h6REhIKvB5vdOhTnMUK8Y7i/6czjlgPLqaV8vH7XoiBZq+V/JKiaGx
1vTFmC7dBDCA767VO0TAMRKYHtG8LIaC3+gd2GyXFy7ZvaUd1yx0JLfBcd6CBPz1
EU693ce38WXd76UMjS2fXMhenf1VhrRlZiiuizmFHcaFBTmMehHi0RLqS1qGbYEs
LPtYb+vxrGnlRcAfElojQ6D38ENEkqb0TmAzmFCPYwGnpkgfm3J9OyLZfahPJ8da
9l3IJfWhH3n2VSEOfp+Nxn56n0ROtIJ0YJjLOar97TCPMJ/OaYRcHv7JfOxzlzE+
nVYB5rvYPZdVpmS9G3kncOtct5lTSTmsJ+Z9m8bWciDZxaRBriQBbfCVaWwh1T9/
MN7uc4DT4OwBameafyoA2+naBjSiX97hac3LuMvGcexPaR2pnB7mDLmleErrPjJD
hcj2RfA5Na0MHVlNJ/DgQ0pcXzTY+mnnZE9gVy0KWeM3GyhbTZdce3EuChFtBdzW
FAixhnJfPLnZtJBXBXjDaab8g/r+PWCY3/yD3Jf7nuWj9MtWH3mS5IfLwRJ35rEF
JmHd8suxRQ3kZDq00IuC06x24cnojMAdTB6m+KT9XxoxKSmktAp0YSp8BTiptZ0Z
1Gk/2VufKhFli1vN5Vj1ICgM7pODd1Z7gHNQntktRYhnFcbUPlHfIdZ+3Dl80mmQ
HDzfNYelnZixbKSVEuSWmDQBnazmczjnnVV0lTL28zp1E6PQBt7fAP40ZMvLP5Qb
eHSu9YU+pNMWjbDnrrBHdmlZkq3oM7V7Wp9v/cDkfJsSvWyqs+Kt+fmAuSc7/63d
xwrdNafukbRKSuc9+x7RfymzGdwHb1+2NccTeyktj4E/jQRIiVpCh5VUgVWH6WKz
FzuWOEmbHSbk3/PV2RmjN5vo20gTp9wUL7Y/4B2yin7kAjS6PU+BELY/9Akv0rpM
y5r4Del58qxOjXJVYlxK13iNOkqONwoal7rfkVh8uZ2IeomhWvvjNglB4ak1aBQ2
2GuJBK8Ftc91eKQelwtpL5TSP5lTy1SP33KAmRPoZY45ayWCWQGSlLNqaY3nALQ4
KgiWUY0s5W5Rl7JOPlQVeXaCakAMwht1gwgZ7PBtksORA9W3V9/IS5Iz3ntfLNKC
8q9Hf/d0VFF9zsoiYzxiDLT/yZlTfTp9dgZsk30sQhYpYdkgDajfT96crA96qLGG
bDxY3teu+/zuuzCbY+jHd4UEvZOcQ9Jt+r2YCDyvM5jjwNbzxAWz1gmwON4pc4Ja
nn8T9KYHbrJ2XfGv4bqT7aIYFLnwKZbHs5Bvdx7rmMDgqtOOVcGbwjcle50e2x1Z
1LBnPkQRRS5O+P5GmBQb3grj0Qmst+l0yhq57erHqp8uLZMZxs21k7phim/2ccK7
lO2JZkGLL2y3ton0H0E1ASNZ4NUEjQZxlvxFQDZeLz5BeJMvmIsbgry6dp+HFdDl
G3lPIgtIUHGDtJzqHgQXh1i/p+KvE8h+NINBALwX13nX7PAmrLnUgkC166r/qzqo
Lf3Yjqo+khhr2LHDa1pOpX4ZAXm15ZyOXUJCjZ5hwiZBq5rctXIw14YRyXuwLfv/
4EQiMxiMN+nNkkCTB7sSCGVv3sCfnjliIRGXQKD2j6JX0sj7EF7kOaxeUf3uOFZa
0yGv6+lEmD3KqVRHtXduWEwO+s6CVUeUejKu05FJiIoGe+O85Oy51BhArcSE46P0
mJpuUa4xmSYBhwdlzhqnz6+7lQxiZ/q/0h+SYGRjbAt6pjARjXQcmHivsDZT5A4y
I31Q4W6xbvZORT+jaVzej5T4SacBYq0WbT1P1JRQ8CzsgC1E1SA+IfVZrbDNH8rO
I5ivgBKOQqbn0w9Fs3nNLhdY7LZsoPY47H1UgWvj5kBMmVDfkgDfrAUG7Pv6b0Kf
QRJvBliB+pKBdk5vgoT8QeAw0E+j6jhd1NVYcHTdTpc/XHPlHyCOUBCzTnpzCoXQ
EuXrU/vfmcDsQjHv+toZBoILu4N8Lwcn7OrxWHQOo8RohrgMpTZHGo9HnPkQGRou
mYj1u4jEolCeQcn+isHepjnD8XV8n5kN99EOy6K/zRcYdZ5ViQt6Dr+8IDQOJEfE
I9ZeKOa6OkeUcXUvLTnsUWQcSehpz6LOFKLb+bGO6x5liL0bUJvvXP0ySJC1Qglg
kjFYawal0nm5QvITh2ZWzJMyZbUEtOtK/jxMSNPX/Zujw2IZ2Cdgo1YWNyrLLxTf
1U03O6Ks7EfZpupJ+Hmcm4QOp4ywhV3qwlLv8VxfbWoZuwivWLRp2f7AsEVgNsTo
+uJXeF7/T9seZ3Rj44IoJkwssDNd5HWOheRIYHKbuRjITRNaJjii1oej3nHaeX68
23RHa8BRKnDXQCmXL8WV2SPf3JCF1OoR408OvEpb1VZ3DgzzGwHGGWKdw3kAazrq
4+jUP98coQCZ0+5yavUcVUhEcY0cMVeZ4DpTtB81y4tyFOlJhK7D+N7LSUKB85uS
0kGACNDGprpdW3PD9OtKXCRyVi+nKkNIl6+JAKB13kOUI/7qtNEvV2ziyhMjz67V
qTCaRUfdAtTELtaf8zJdL1zh6acNUGL3kOZ1sqddCdiIp9aLjkmPi+1xnFP3q3+b
G29c2uRBiD7kJj7XK0nowDBtgYsi5SS/blHvD8PkNxRUdSEk2YHpozD557PnZ5rt
1vkTls9BrAFrw1EuMVtPpLJAAvU5O1Mrbr9R9rmVGj0kVyr38LUj81Y8TMX03nbv
zzorN5nvSqkT3uZF4SIfGL1JfD708WnAVoj/wQxAwkKu6+k4nrg1ViqRi7ipNd24
zMkJgsXW2MBfJhzmVX/lJUIZ87sUFTEU/GITqyvWzc2o4U4KKp14e1wiTBV88jyH
8/dS4XlRS/eBKCGb8KmTGFsCzX/vHc492P7rn5ndXG/d7EBbKmYcubaolpC4LzhN
VjYM6cfOU4553KwWRiGQ4uZozYioF+LDN6ig84oEwFDxmJ36+4HTBYxHcZLpsSqY
brJXtF81d7A11ye9Rg2hBPFA8ahBQerASHP3HhUp2f33Brymi+1LebQSJBZAv8IW
1Wy0KYUmSqWjfs5Yu0IsILyloTxro7avcHX8cam6ZClG0JbhAa4UpKlpHbPHuWXp
tgp/KubUXQaWApsEIye+z+kJNPXeeA84VElQpbjIqqrlBxrcUppgzcnzbywTFozX
6b1Oc6fXs9rveMFFEvTm/0bE9iCkKZjmk8EkPouHEAya6tCvvRRUStTjM5fh3Q7l
Kc4QQKHvhzI49/+dq1Xrjs0oh7YnV9dsbTIo/dQdj65E/n6auTE72QLsqPS0UI3b
da7YuaNJiIsV1bYhTyCBqzNNwtJqgEubase8loA85rhW2NM/eZh2kcfwNXd+6XsN
oYuvFpU3UrmBqv7FYsVLhJC3WeVE7/7bzyIkTAz2aXwmQL/ZMFphjv4QF7AdMoC+
iobPXulYGr9ZaL8D4WvvdZLOmM9U7AegFoox6iYL4zRWs6alu5oaRb/nb92FcF2A
Vx//QV70YYdsedkPaDIjeCfjOmiKNzKKisofMgNtwM+7ICtoDCt3wDB7NpLyzsuv
HV906ZsnffEYFjzedYrvFsS5i7MwG/CudfIzpbChUGcWtT+Alreb0J1gNE23kGKS
duhwY5/ZrwXGZ8JmeFNHJ73boX9k+vBvT2rtXX/JZlBjMgNe5PJd5zVxP2DnMOsE
ll90pqzaUUoerWvvWnRPH4sXKF3BFEQ8oKZhV56/vadMzuA9Hx3yidSkLXDK8Hf3
6knZ99PcUcASFW48sAdNs8ZsmMUQdn/0NrveDWm7H4xO2ehWTNR6XC+M5flKxsfa
GvUvjNRL7eu5H9mprGMYT/LhYqQ8fYBwtTrwrwybINgkpjxy8mMBnvuweuJI059v
2qwDoIv1Mbd3DHwBjuAaE6WqVFxyMQCU7oc0LVYnJzZVpEuLQ8tmsU5kq7V1gHU9
TrP6lFcLS2FdldJj7g7wh4yXuz7XoIBsjYf1NzhdqNx32+emyaZ7Mz5qB2hf8lMP
dmhQbHcmRxatq9zJQv0fkuaKpfK+oqg9m1ExNRUZGCc3ewrW2fUF4nXMuBptd7Lw
TRS6/4MS63lLUHRMUfPPzLDngkjsZZUu2vHbI5STuY2vmupYuju6QZeXr/YgPKfw
qE8zImOizWNv+8uTXaEx4XtZPJyuIYIqrEhXHqIH0EE5iEmjF37jt5pFq4AigsEQ
d4GSdaCOLAn81T/B35JPQMSrBr23UrO67j+dnu4IbppgIc85U0h0xa0xz7riIKnn
Z4qtd6FGeBjDffAWLdmsr4izljX/z+szRLoWWI7s9FMOrlTEUkRDBTUSZXzmIwuD
dT/FhuwjCQjvw+Tzxq3mkb2Br1JXFtXi43mF0JstDIZQjv1vqfUSgFdtcE2yZsP7
5ooGzkIC6/YZ6RmszmxfFHhtvrdhqOYlZAVcan3xSV/IV7YfElpvBukzv3Rf2OSM
9jnUsRClvcTcrYfezXSViP9NI1nZ6IBht7P1ZMNHxUZOIae/su9i01zzn3u11M71
m/kOI/xNAKMKvZyat1lCUngj0Y9IMfp5uFJWUmmD3HSTSPu7dn2nB3BAZ/dA6Iqi
aj8oNMmWx3W+MPN0+9kMMrYiqKgxKOi30TVoPssYx9FGjhAOjDD4fqy89cnc04oX
vZIgJ1n8NsJ5VAgPZddltXpsl5WHMZCGnpuD+QXD2+v7yRR3fHSGsd2ST+jfOdVN
3+Tqueuud6Fgfv3DoGLbDADiQTL54f4ic3X1Uw07eiBGO06YJQDyQOPDoTbIw1Uj
ABYGy4Vm031ASsebF9/RfFtOk0y84PkyDah3ejxw19zE2zOFvSi9tzGrrzIjPqQX
vmCyavUglmc91U+nMCnHwil7DPOABuSHLDkUfXRKDQ20jMg6X5WXFLcPJusdHDEJ
Y/ww/iz/Vfb4nZC1vH/r1xyN73b8nZLI7VH1/H+qXWEoBS2+HG7bRyOO/knTpiux
Gr+zR+BEhKw88JsiAP02L6bWsW/K8NYq75GzYFAhyXTuJRA+6uJqAdD1cxEqyfCh
ciA94Z7+MOv/gxfFnTdl5OHwgfn7v0tMx8/M01hTscVD8gwvMo9dQcldcPeoz+aM
xzzWkesrzMroZtSluM2wEZDebqplrXT2hD718KaplwMRO+2dV6Pl3Mf2C+idKDpe
CEHUJO+BeG6UfZzJwCkPCRv8C+A7a7TcQJfV/KmBODIMxHnDC5hHgUGlJbh7MhkY
nXbnytF5BPTUugqBYEFyr7eQ77iK205LAiXCLAwSbVtXAZPqoRnCfAF9JytNughp
/hdNKugKAdpMQpoqZFK+oQ5Mv+8dy0tUUU6Xx8Hzhg2ttQf0oxTlDY1nKaKOP7TP
aPUbSRXPtJonaAGW8zOgQz3vW6GwEaDxCjWbpbFC8SH9I94xQLsq9LIIg+awsdkG
GbmT0weAbaJ1pT7LZdYc/282HAYqh9dyB0rw7RYm9H6NkfVm1G6u5WkldMk+ZTTR
er32B6Tkb3hfMOdcG/9cMncUKVDsYCWHBvuaEsD5xDCdlXFd9Opht1jJLs3iPHIJ
0d2pe+n0S51jcUfVc3eufRlZjbS0S0Y4+H//51axkwd8q7ZLWaE3RRGIDD9q51xK
F1FXVQQzOMRWZQ+rZ0q6CwAeyyhMDlYvzqru8JF72MSDKD1IfU5L35IoSiAnPTsN
MWYfgrQUH0QniqQet9w5WucR9EUNozT+XX3Ue5niPnvRX6ndDE5y1PUQpKgXQOX0
CCaSiNgjB5QvhTJU7rxCsZ6kFrrHy8hL2FSynETEdaTI1E60eFzXL/DqiQbQ82Sl
vNIwQIxjXaX7qRqb9TEJS69zcNC77nU/TdBYNCpBJAmSHczcD2gw6f+oniiJKfAx
3sIOYdy+117UWIXuHVf2jHSAYQvyerqslR7hmES8NC5ldzDnyBWzHHhYKwAf30mm
9Pq7Q89i1aJhUmjZ0LY6JKkr550jqL4i3tZUY+StjQUMrf41b8zobrFsCEjthi/K
CV+ZMTZFEpHF1yz/1i4pdv0mLUczxBuRkvLHil1DOdGWz6AwgJ4kuXVpnkha4c3d
2Wner0GcUiu3FtRxT/YplXUdshBExoWrd6RByY7Z0AThipafDzRiV8nEpirT8OMQ
K2pxv8SFZaahX3nTjyMCK0DtdBvR1+Qo/NNCFwYHdWFLPZAuCGOyYCX8PfhbksG3
qHACIiCpYlnQ9jo1GhdOJwgqCh5AR8j5Laws5PU7W3xBEvPwEfxDeBGZR/Rt/7Ej
uivO3wx9a3SAyX4mvTjkynZ3AZKXqbi66lf4/ira0pnwPfNga4ZYpG0M/f0gXXkW
1BX7AjUsNvUrMz+uW18j6sKPPxv7T+1XUs+wmOKe07H0aKmRiZGE/Vu6oQpL6o5o
GmzEzBLKq8ShbZMh/wIESn+Si0N/5F5qL6wCV9E69chwI1AMrRr+eXw2yNO8pdo/
4iY9NVsfWmX4IiJoBvxBtRPctKR49Ekx6pIpRyh7zB/VD/fruDETLqmR/LiNFJwz
BQgRnCJRjO5Da5NAyCgj+D0ZpYP0Dc3UDIPGCnKBkAEDyKesGN+YrzVPRuZfUMcQ
FM9m6q/A86GGCUWdbetuO4aBSxYWBzo1+fcKHkuhJF5J06DhCrP89qNJ5Z5YzIXz
ieIDCHzuPoYgAaz5xXpnGoJ3zrRCoH3hxasIE8K+JGl+e5yTBcxCkv6gT+F4NPIX
urQRPcVAQtH0aVJR0tUBDcK5e2bDJPl1+9bvyTzQwV7QmJno6lAPo4jvPfij4OJA
OagKkLlheyX6wiohIVufIJpAc6iFyXYmaDLla32R6v6CJkMKN4/bVB8OTwi02MXd
PXdC+AvfaQKukCmFJ2NMixLDfNWC0VQjdKIwBss9YxJiN4g9dZTRnSzvoWVWENaZ
aW9ZlKjbsxYY2xjkWmmwLPGMNYhH+x4FGbUEoYzAjYeHLxHOyFw4pMtyy7/BC77S
8KIMvUgVpe7qVEe+o1Du6RMc0p3UlKbY+fD2OI6wSH0J+mnoLh4XLmSoYAuGe/1n
Qm8tbOnc3oV1eSG7GryDfC1qH/3uVCzgm3AzWxuuZJMo6UaCOlnKB1uIN4A2nAu+
aWSwH6VIIzKcyIan8w6lwbeXi/6KFqGcMQvcm+DuVJcs0h3YFa6gnQTdzgv2uyHb
WxNtpkHsHLOWZwewd/yyL83NIxEKpO+hO7VA2wuAewLQAIS9YbKaqWZdiC8eTQTt
rXu6CW8qtEjdB8FyZhzztsO4ITYH9R9ojyhk1o9jcQ48M25ossFiKhGXKKqn2fz6
zRMtk4lirz0mPmimVp6KOQIDp1tDKI2fV7V7KXD1582HUta4ctaOkNNOl5VpvDiO
9XQXftBgH0ybNCuENQHbKoTPu2zzB8dkYmQeF5s7X7J8JAz1r3y6Z1CVe+5mHf8g
HUULO9fnqIpd1BOAxOZO4A5bWeZluhnmKFAzEjpXyj3R8F6QLzDITyDUXZvPj+2w
YAylEiXA94TJDm08va2jqXr/Kh6pfW3BkhG9IN50ZRdIkvc4viyOJIUrCLQQBYDc
1F6IaQi07Ucna5BLy+MC1mcIBsFRKMVQjS0ne+8U07I5NshKFLEmTY7riqSGvxEA
zRFvei1/SG2SrfKEYh8ZS+P5foWpzSlOLJqsrgHaNjRxYDhlRgiZvB3UXXdbx05J
t4CAnwDzp3laEwiINdUo+tFq5rDEao16Bx8kU+h/o94eLPBBJe1AS21uhUk/fXzm
uMukiFRTFoqArRwT1ib5WDuo1+VsjSDE6aN4QfCUwCKvM987ASLWlHkH3iBQcgzt
/s/sIAgontEOh6esKSq4vSvqmYil9DAOANRnhitZ6S8BvVnEzocJ/w9ymlgiU/Q0
Uuj/HIdFo9Qm67dTrJREzEqMdlUEaL9SumFFsh2HC72W8D9R7UQSpljBO67GLzOy
J+WCgzBv3mZ9EoVDuJn3dELSpmd/vbPVaFMdfG8SpA/gK8vRmNsThhgX2wPUUicd
itQUJbMgpD+1W5zlIswjqfXHTgmIc8sqk0QmmYY42qVSHCnRjkB9lQb4SzVp6a8/
37oB3naSPnK8aZRDtILAzG1StSiXjTKTsASo/JGdiuPmTkHbfSAofeoYXvowyQdR
NL2Pv1n5xUAYmUKUHPbAfmbxyUhrXShsryXLIV8EOcCOe3l2ik1E+wyAmFQNLYd5
YUnQED1QI3Pt+8/WE10pLdMs1wplT0JBgBsM7ip8ngGzIN6otI84uTiMgbtukdVa
FvW0dzCV+P5TgJMwSJpOm8dRqoAQUdhZfT7x0xr7SPjprGrSVpXkqWWRwHnGiMtH
Qf2/6kgKe1y1HsCKhWZK9Lv1DvyUFverxGRTvGH1L4VSP3eQToteIUI1MwODwBHb
L5wX6URymjWrnnFmOpPHLZUrL4vtC43iqPN6I9Mo1sQNwAmSEt07j7agn/QIkgVY
fd7zKD4sJaVJ0fKJ8L1Mmv9wfTy5BgG/vTl6F85ZsriyWF1FQJfbVQw0FeNxBOMf
lIbGAD6vsIUNKrLTSTrN01VtgdH+jo/8QJK2qEq/E2GXPgUhXot98/X8DExmbtuQ
F8vdZRNWYe3TPW5VKmg69vTzFpmBQJlI8kLZB/No5Bl500ggucVTQFbMt/hNczmK
nwiflGYny6hej8Hc5Fo9ZKpbbpb4eXAh3esccgWAjh4wynQ9QRQMAd2CiNEz4imG
fJVWELsMmBVhX4pJE4VNawMFMyh37f1WVE2AqIhJoV3vv+hFp6O2FxWoYZcPPsTi
WOBYTp/9pll1ekT2X0kop9eiGg6V8FdU7voms2nw+9HA9C5t2RbYqCFdxhjOS0IA
oA4O6+1yjnWW6jG9+f4aqr7Bi1qQFFRoGLtIivzblq0OtJsIA0XjuE3aNuLhjF58
WUQa2Pkj4s8z+xFKb9jfSDT4s/Qd8ab5XWDT/w0bbfIJPJp8mTIhqe9aqW+5jwCa
ohMlJgQNo5f+rm+gUUHDdJ5MIfeJnUUHYD8swAiV9ZcBLrMyLxMV6w+Z1FkDTJMX
o7X3PhCubuRX58SeqbIIT4W727Y4sfyIgz99ALDMZkvtWYMo2TwBJ/7MOkl/wbpu
hIotJe8pYlXeIQ25xZX6Y83iSzmlRLKQVVyT1Vv04b7p4rryXxin2PbjE51u7/2D
2wpc1o61suSnctF1smcp+XCy523G7Kjv+guBAx/yiLPsDci1xSBx0Bj2edKMWa3G
iPzvP9ALj+cersfLsF45LB2RliiCYSn1S3GurvzFkE4l0ULVKKkrwRxLb4l4zFby
B66O7nDhF772VK8sN02ksJOwDwbf8ZfaaOSsk7chQpI+JPudPTULOddMLjksAk1K
vp6nWRiUwbpaR5CDhaT+bEwG585PQMMkZowXvnigO5QKppw5hAF8paNS412l2O40
z+ryOzRVs9rBi/9fbQTP6eHcv/RaQObVZgqIpxPl6YJFwF8Rcnkx1YcVaF7gRVhB
OzCDNxlr6btxSepG+DBvuHGDOX1i2XCUiguMrGuV8rEF+zqgYxymkCcXNmX8TtnX
5ihsUezhwVN5HIxlrmIU8rrA8wQTIwPROUYa8TmwF2nnc3uVDvBpYmj8tY0vPM7h
XK05AmAQEKyHTaWM0TnDkllnl8KcWJbw9XR8gLnh4d+sXjh2JacxIWu1yEgJiXSG
MMhZZmBUJrQjzmOtIQsn63s0ARZTwXHq+Ru4t5IulhRrXBLEM8sifI+Jnn3oK7Q7
zHdfvKfCWB5UdCIyhL2TSuvk2fpcbZjtpqdozFprADvrDrXh4YNjO77EJcpST/vg
1Q4LgiIOrBdu63cxGs6evOL5LS/DwSjI+tdPOVltP8ZGUX17gNIa72tNpzbh8vye
7kOyBn1XFTzazBjln+PqIy5sQOaEiWQ1yBNj60ZgoMbWnVK89aWE21dr0EBLxWwF
Tltr23oHgzK2iPpmpCTrIKjLxVdHaL1la4g2qjXiBgEgDNdPOnTgg6Q7rvM2j4iD
VjrnJCbEkn2LdRT/aqYD+KEjtHMcIjnL7cM3AT39gJyZvw0Ikup5+b8EMtbJk2U7
YwuFp4feanCa+07AU1ufLlLkp0hVhqQsIuwPuar4cuK1OWfzM9TOEDF3marRO98s
EQX/aKtSyUrgY7qW3CFHYuWNIrA8qH+fFyDdE3jH2C1Qqu+uWUdpIS5FYS/zl2Iy
+tiAYVX4iFBQ4EMuHN2iSOHzNCEJ853sU5SR/zEKikts5Dik5fR/IanArAt5uEQv
yjh2Ih5+H+mXoWb4Vq2jBfZaofipOANkzEa8o9rAOvOl+LCYkXMrZY8aJDWoSvSo
8NuSrbGKxHEMKTkc5UmlrspHF/b6c7cCQY6fA8P1EJEiFViYL6qDrEGobSqOtmvh
vbQNqqe+VGSw7xXdSMf0+la/AVtPxl7CFpp7W9+fwjnGyOz9avo7bSi92Ajp22Ww
5GIJeFz56JaLVfJuONFB4Z/0N9BofK5Itvxh0B34B17WXOhZj3dRLozU/bXzHgo1
czxm2kxlng24/JnvyO8eZrlb3VQC4XoANiAule616L4UdMkIFTp8azyglpSaSxvn
Nmq3rfbJFHUtN/h4kdtA3TCI20mLyPOg4hIuvM5Is9kfDZ+tlTv6jkaVSbWqAgqF
7ukahSJ+AMOZ+U8dAupzKevqxCahOOYdal6U9y3Vq4bmxyUpNEiMN4BsmmOc++GD
F/S20DyA2qEaTd4W/hnbpZfpDhMOx8VwC1BmGNJcurK8uPFYZk6ZydsDbicH2i1T
KHfPzA+pzRWwEvU2u0REMvSu5vcDtzS7qt+i8ViLAzRPj1Wt8e/Ii8pQ3XbeOIhx
D1EbcK4RDYwetFxOGiHTjNiKlRD05VnAUQR3JYJlbq3PNWDr7e/91o1JyA5Bke6B
3MHIcwyKUucSRp/bdmzqVPTdYDB+kbpfKMSaWi3HsV+qK4FSW/z9XdVRguFvRpfg
CyP6CI/rwKQQf+VexP4HzCoSl8I+i8WOBBtPw1NJxTJizJ8MjXHtZjdYeTDKCDs1
z3T/Tu9BsZnTglcYr9DdeT5/Rq1PgfHJEzD9WZAdnjpDGU5d0oOexlA3ofKUuxWU
GwYiFiJntiPlm+uBzc2D2dDfTvRIJ5b/VcEKfTrzmdlQnIM2z2J6eqNvsH6HJhjb
8Q4qmk/ZHnAGrI2ffkdI/bVptc1hiUXznn61DwFrUw1m3uqmdP0WsALATlXpDCnX
dTLoKF/1/DHCHjtEr5NMFTL71oj6Z+ewUqjTETlflFUr8eRsE4NZjDBiODH6A6DJ
dmu75iLXUR6X7aP9W24xbetTwjN8F6LIkpwhYdytH6AdVzrKLpPXfa5TyFSqm3Lp
oxJAFHxCrZcyKbsVefxWWGP1iHMNBQIDRXMkFsJXWRDRR2esiTPw1Do2iOWEmJAB
RylPpm3DcEdcnhCZ9W0OhJBJsS+eimy9nQWj8dEzjDHRq/hRlS4QSViZUf/SL74b
CQUnFvY7vYKNUvB4nPYke7c44qjT2s8KXmfoxdDTfVAaLSFGmNv8Nr0CR8N6aqZG
1ZwkSC3T0/+t/jth0f7AwGyvG2LiNxQYlUMWCD1XNxV6u9DQWI87993+ve1GfNWw
NKwQXYHv3DmrqfLRTkbWeLjHfwGmhgew14MDtIFt+9h0y6cKBfG1gdGmEy33qUP4
CG9hUp1qNyCc/n3xH8vRdRbj59W4LG4nuVtxqDxZyT1Hc6kvLWWRV9O7h/rK1NCX
eAANPzlg5jFWrdD8mCJieA1LnJHEt1yS11cx4uZFCEHTjoP9KvaTnfu3vtwysI8F
N3OvzyjlL8moZ52PtYQDrE2vSC4+v6Rc1p2W3W98MK7XO7bkGm6L+JN5uYTB4pnY
WXOZmEomYittF48t9qiE2HTSWmDtXKvYDnYJ5B5Nw4s7lJnDBq2RzPW6Rtp6iGKm
8zr4TwwFBtOLjZ3bT0IzZ6S5Ptm7k6aSareBLGLHY/c+GaEmCKmN9so8ESnU9hev
OLsuVGwEFW+A28TsVpoRcjDxkkfn5V0ub0IqJ0V1nSfoVc4mSu65BEJ3ZFgLqvXC
LJRw6+1gTFvvKnhrx8LmmIOHQXolWXuNEDSZexdyKpP2qMrpK9Rzrsc8rPGLH3Rw
bLWHkyWQRzjys+iU2Vgf1zmhL2f22J8tB8JSjU4F4KiqvG0woVJNPVWgENfpFak1
W+D0b/zAwmU4Rytgb1JS1TweN+aNQSxZdx4+pA4kXo12L6GJk8Cb6kIRO5Cm1im8
pJj6MThh6g2sNnhHx2qn1sUdXBIDp5BHnGqNEaEKJCnhYh7Y3Pl1na15v2OYoksR
rCdTWDjw52PEfmAQ92VCMaubmWshwPOOXWkfVUhHZPAFf6JCViBOx1DZPRyFkq+8
gygoC3p00+nC+bLmmub0QSCzfuOduF8MVWAAJU6ykYMmEGVZzH2vIhr/+mb7nvT0
hlvgfZSajBfhYhz0WDgDQUNT2AkY+tdUpOPOoiUVV4L9/Dn5CidqRAd43sOd4LvS
otUlExAspDzko4PRJVxHXQp5EG73l+sHXVd+ZwjxKv3q5kQV5N1wXXWcxazyzTkr
N7/g42UgpXEpfh0BbbNFX6RupdsQ9u/8d7ayjyo/mfH3BgPKBLwMuZOSvEFI1ZG7
x9zfeB8RSwfP0dDNaEMG2H5C07OAR7LRt/n4pHltTuTpcgUFmEuVCcCSl47Q5zPu
kB1I+vjdwbuZqTzzl/oPu9H14OiA9VWxUrVpjf8oLZpkzB1JA4VoKKZ8pJnWtHD+
2pHujfyjMHq8hwmq9fIbutX0xN5OkN0MDhvNBgLKLGqZOHqdhrNrFf75WN+5usEk
6cqzNt1bgNcrBl1rkq8DQG3OQlINjOltNnxQKFmq5zX1DVApoB65GRblxgRaw9lp
ygVsDqPTaLgd0rIPqHe1u2Ok8H9SLloVJAtdP8RZUyYB9Ra+6bfw8xJLFcBNPMYg
TGZUu5XtcB8ia5HGpUuOVtH9eSQRderMFN1voVHgS2N9bDgG9y3FLaX1bpmIEtKz
/tDTTq4GXO/Yl4cFE/VvjN4dvSezttUW7KdYTFCMHAYZV1BGBl7ViZh6qFwvoiZs
Gv3JiT0rgDB6jJFGVzbnq6/EQqALcHQaZqsCuu9yiSmolqsA71ZLVlinJllDZ5TG
2MYk/ZvX/354Jfw+xVnCiXa3Mt2tfsn2lj79ECWct/jtCClX2SvrGQdLcEAZ1FC9
YTtCyeuJUmgMVqBGviyY4CLN1avSDEm90u+Lm2pFIiVoZQDetIj2hNJCxuEhlaTp
ARS/I3Jh6QdurwuNYjEAoPikTyUrz4WYLBjLtOB8Oh8k4k3RrEAW0BYZOnChPKGO
L48IfqqrQAcyE9wUCgstjp18/KB94x6DpOs5AWkuF6R72uQUdnN4cCgJU2VNv1zY
rL1unRcqMQ4x2n5AUb2/71hVsMLrBZiFc/E5nAUadfQit2OGpraYD/Jz8/C9ZBdb
03gl7P/QshWVLegpVVolFaFSB7kU121aFbc54nBTxGqpPzZAFmTbCsmNuIY4j9j1
9Df0bZfxE/Z9tE8jjhJeboAbwkeAAR3YRqLdpb3R36nxVObxa53N42DHAb2E5aMz
a63a6bu6w6R24o7u/qynZ28bkMRGFJAFb3sDmVGQQJn+s85HMuBAcE6rGIYQhGDW
eDsukisFQuv/uQf6v6n8VpB3ZBi/tydHIdIXkFnjBKgZyACBU0P0V1m/LWkWPAkN
vR8ruxFIm2Uc3+HkfhuC5URyGuWygartDELSS3JMmimDjLjjZexZi5evlkiTOpmx
+D9SdYbOf+/uIMqTqWFoxorJ2o0d4XCtG9HKOqqXFHg0Av8pVrs+yZaraPHmPY7E
jU7rGXvsSqN8MKbCgLOB2XECJoX5RDMkQs1WnLKjUTsszZOyv/7J3MLVn0FFA0Yk
gFcX7843LD3FtuPtaU2/UgzGDNAqEsmmgAWEE6iPB2Yi6HaEsAGMdP4P6RrwIQCQ
DT0PakdpyS8v2Vxa+dtRHyL1OYe/KUttCThFtE06O2CF4z1sDRoNUiRU2sHMEBpv
VUX4DHBZtct/K9g1KZCdl7obJFNwHlFiuhwBc/54nIJNuKhldROp0TWuQkYZaMcD
nqytXvF1qQjq8G5MpopcRFGh4Q6Zlr3oFIdZmLs7WDNtM+tx28+hwPjCh7Y0PN5i
jhnFPh2gR/s2Nt98FQUl5ZhpJbTnmxHRMTVQIj6d10leR+iJGUKNi+H9emDypKNp
mDsF9jyoySvQRKV0zT3ntCQBoElzyKueyW+F21Zs7hbQEF/TLse6Y4AcaNCowK5f
neRnwGtmAs9QZ04WztciYdoPndoxbkySZiMKR20xK2n4ofybZWKuAd5zUZH3bDw9
o+n1lwC6iAjbGG+5CSCg1Lo6u7At+fGwuR1MGMHgeEbo/f+F0zs3F6uYsHeRfytE
BSgf+jzHH+eZLBsV/ekbxpZ2CE//t/mFDF3qCvrp/Ydq/7mJer574DailAb8GDe9
JIjqHgsHG8PKeluCtbdwRrdBil3vvFFzw1hPkFKgNfHWD62rxuS8nPZjSaY+2xlp
Htu6JVlmBhqGIIIP/GO0tzGppH5RDnK/fI5jKWut03BO9lQNQ4frF6FmdoVwJMCf
GthIQCBeKIviye6GdXUkjFwGxydos3ubHAXio4wXW7r4rez2LGII9e92KMJlD/ao
W7ulWmGw3BTupIiDiNEyvTI8N41tGt5q6mYUJwkz9fPCM/qU5afnFdJ26lUIBRg6
GNDUKXMV5ELf+aprnfeJyllgjAI+/t9I77htpy6TFNayGtjVguwfhRplbNduc4S7
o395N1olQ+ICU+tAR+LsVt0Q3t1nCd4F6ZnJPFBt7hbNjMd3/zJKPKADcrzQv4tH
YcRTCx+/w+1xEfGIN4PNuCc3609zjKfkSc0MBIRBntGfeCL1aBzMVyadK69MORRL
GvjisTCBpr9sSWDOSc8VvTPi+9VpmV2V2xFT3Bh+6tUiQaJPoMRhmNagyo3vMFtb
3iikJpwqPGvVoiYmC4EjRsHk7/ziY+K9GnPbplX0vs9P8MPcPb1ALtt8Zpfr8po/
Ir7xCp3gSjMrfZ1SyfyzKtQEeQB0EAqkO0t6WMdJgNaLyU+vJrjo1Bzlsvf43j2/
6+UcMPcP4xnLgVsR6gP2h0VHikuCY8gNZi+2XS729tCIBqJqnk0l0D+HbogWDWTr
A5Wjy4Ri71+pPdCdcwMIaeBFQHeCYH7eBLRXzAwevgz9siizIFcDEuIIAf7RmcVW
KnR29fnj9akd8AAXLHM48Nj+bIF4UVVyJ3zwPSTLb/HfxQsfDR82iR1pgcBc1dBe
nAof0MUfIxvn88vpnPrMU/+hbBa197U0S7ka0/PETAfnMZCWJni7AV9BYzEpnCo6
lycTXMeERHl5IwuX81vIlLPTfRO9Pk5WIu4GIfEYHKY4pM7A21n4G9ixOp+CJI9s
701COaXD39mzD3REdcO/fHvxLtaOIwyqfaWrwD/RDWIIjZa5GLpHuiM5Emr7rX1f
88GKhxq9MOSunW/jg15p9eIUd1OQDL1YK5MbLBPsQTpsQiBawXMh5FF8Hr8TPD5s
+nhXrA8zLWsdCyYr1u5xryW+TYNZGxWFfxs1/XllGbUZYrTt+l6iUtvdtNJ9ansj
JlE1s3Lmc43ylB8IJjvQ8W/w6KhqWQw5OImK5450h8bnlXbprfa5sxshR7Zp3CTd
N7u2AUWi79FHknmtHHIJfGjy+SsN1kkA7M+JvoTeOmrraI38sd06d4oSaFNxrHw1
cls8oNYQDyTcnqdNZHapbGWIq2I2RpYChfwamo8cz+fsp5M8II6YaNCvBDuC4Pxs
gjEgfgs2SWxSXAZFv11x6/QGBL7eD2dl8CsAXpy0GpTzewE7iHTLBYnqwz/O4dXF
9zOoZ8T5R8kPeXJiQjBubEnWSdSv4L3900gf+JHDujOAzD3RP/Yrye0yK4TV61rO
qWJDFA1Wj3ftsD+GROliFyJn//WTaQJnLZJmiLr/6k9eoC5sMUW7Gg/AbqixAv+l
vWbb0zDOeZA7ZUBN63rwRtn4DNcG7Gof2TkktggYXuNaSu024ikItxiiRcYa11uH
Yeqsvp2cMEXCWITf1HX/6z6xUjVtS6xcD3s2gxjY7oSg9SCNxjweLXte2z+hzrDR
nYEzMtx0mwLaqwETlS4Sj2NZNLHVvRMcBf3eumJ0W2VJVrfcHlQcZwOhppByR9Je
cy8esrAC9kZhszO8nG9TZvCej9oylLsUFB92VOMG+xsWh92l5tcsjSHlyjML1dbN
ga4biVIxerUz6PXbSs+9DgjVZUbOtzUt6eB5P8bKG/ZmDcEScYDGRlXl4kidrgFo
447qRf3hpf5xKUJp00Og3JvGmrg9yKGtzYGgL3XNIygSWcQQ5rE2ERQC9a0sJZzm
mffO56tdOK3HYsFPT8x0wll/bGPBvpSReHENQQja7Qw0wzYljv/rvKFvaqezdrl2
4Q4QFN+BLVh939mIRcr8Q27UTEhZP5/uOmcE98zjndF4C72d4g1RWuCloToXD6NQ
YxMwdmsG8RwpAAEVc/0I2s+hS54NSVhIAj3yagv/J+rAPWE9KatjcdUQeKxA4CK6
rMVzVc6gEIM+Jka8600ifpvzRqJ81Hp9Wvp78AZ9Nk5JeKSnL97K3RgQGhdStSl8
b3libCXLwngTq20GJJKHdPrUyqKpa2gUOyMjM4t6JMTSdyUccB5ZVA9vlOL1RvEi
WxADUnGVseyFmtOu+s0mBU8HNNqiJuFfe6e2oqYNnpUuNyD/O4Pzz9Wr5S8soog5
CGANxOb8GPjJh25rdd+7Dl8vUGpQ8SN/KcAXEKd0qkOV/Tr6zAoNvS8v2zHPiGfG
P/A7+cxX9a/+AnsqBAUwledpqchVRQqHeV3GoG+uFcoXzdmr4moEzjScxBVt1W4h
GF3A+vDXE6kDBF2x+PzOmqCMgr4N/ZYc0CUMIRvYgrXbuyqmRCjp5id6UvvQq3vl
eSCLZyfWbTgFZ5DPIJMIe8YkXiD+61fsibscU72psawP2RPtyrMVFBanaC5DUoOm
pkvlg70cJfipFQ0Xru26lgeXgBb72kTY6GRqPUigi8pNP0YQFDypVMO8wQg+bRq+
2JM9l8x6QxHpSPtgRis5vyYUVGXI8hQF+rLMNF9W0MMKwZjRwsagbitQIpgK/iZC
xrJLxhtp326U0RLxUIuKt4NrJla+f0prtA7DvMh7N4tjiRsFQpIPgjNTQyhMyTiV
6+PYGieY4im59Kundiqxpwf16/+HqDjpKBTjj7yxrykt+6m8bGgPdsFTpylBPPme
AajQKAll+pkDCVib+0OQq5L4kOgYX4kaHTGOSItJbZlC9mwYSReqKBwqvQNVChb+
xd/x5CtgB1rbroK0jMgxY3jHwxSNrr/Xab8tuZjlyMJwbqqRmCMhOsuepyYmd7AN
92AFWdoVorOSkm7KjiwBpf/RpaSh/QUWnEOKq5jrrdRtVaQHcApQ/4cX+S8TZ5A4
s6PaD+3Qse/66UJc5e+RLMU5bANiimMioLNa3N7qTqp3ALvVY1H1BFACUixavEyp
yCe86aVVOdW4KyhaP3zMCwHIzsrvvDkStNNYhEJMxOlmMEroUkBGXQWha8y5uk/L
AVoqYHRSb/KU4ZXOJl1N2W+vW4elc/zyy1r167fbzBGpx/JrjFEOcp+LuK2zMmqK
rjfjCE9cJ7fsiGTSNzDcS454yFFjcfYBWcCNhtl+HEBETFf+9knzvaJtWTg1K5WX
dnhNlWydILyqfeyVMVNqhNDJKHTlNCtw2lOyK+eDjOXyyu9F/0gIwTYtavgRNGuI
ovt6kChbm32X9XjJyNr5PVDm7bdE4b9GRBtFSem7tdUeWCtmX3Ci9QdvwPTysWCj
YOTfJxuatKbP3mlMkc7+1AMvOHYDH7zzrhEqtEQhaFG88opm50zpMFdmMC+g4PkO
skGAxSpu92gs+K8oAc0/YrHacLu3PgOx5tTxx/w/0Uzw3D7TKnhGNZIjeE25ecm9
zU1cO883NpGRJV3j0dWjQtqIoZ/lwk44YXHru7NcZyMR122zoqG0KXGn65JpRZez
187VQmrhKBsE6FSO/WPww9juyS2F7jUyZxe1uzfXgTN99pyebv4Zb6ys50c7EccC
8mWkK5s+9thVaPcsb2dK9198KoVSqLEFS46pHtvjcYdnOFKDTRVpccTJqbuU525o
5HHTq+7zqL8mlPLGcx+u5X/OLbw+QC6QGqhjeTt7++o5RTiO+FhoQzP0W8TzKV6+
n7JcAtH/NlIv2DRtwEzqQ4VILJaBp/YicKZV2nqX7gek7n1rFecuAtQ81akzUF1U
tujDB0f3b41qLVnx2TDNixbZySu85SG0EunfwSAL8bZbzoYnKRAJMq1ZEe9M9nl/
hr3pquwajznZErfXF5GM2HcjgFwMzTmSthMq7dm1xT4qAeFmfyNMLmczNDSj4+XS
BJS1nxt8stpBxkp4WrmP4j40TVhnPwwbRrKC/NPGsdaUqyOBRYamEbQyr1PalJ7g
u2YKIlW594wOj9bJqrscK9cAVk6fckloRsGs0OpkK18vfXiIBHYv2gtrZMe8zuik
ipurDaiEPGadJi5QfIMRsOGLVquraWfukWsS6sS6d/zI4LIAGdElnkKNd5HB5XSE
nL7SsMCnSTv8TczpnmL4oQMiklIsOSou2f/+TaTMKmPg4ubpbwOzbBKvCcjJ04E9
IzSj2jrgh6b72/Dt1tKPxTCt+7c/aADVbott2lCVLZnJq1TOPOBo9dGj/QmrJ285
OACMus8PJjj/POIna7TTTos9DpBcZU2sQvERsr2bFx1jZhPmoojLU3pwiVfHVDdu
4kVn2q6IVd3T25gH8NYDSjt6Ji0zXUHUVQ5IT47+P/0byoGfMXcDUHLMlS6n4Pyx
0j07V6ICTc9ECjErANpef32D4uk0c7+pbX5wx+TBG+7SATOrUAj6KbXPeAuka370
BJng5ImWQ6EcmzqgBfOprhcXGSMlbNZo6G6PjRBFadHBQ6Mao0NMOODJvtQ8zlhB
wfUUSfot6D3RKYp2P0A3X1aBQKIsCH8hQXI2SP9lt9DAEq5rormb8gVCON/66V2F
5HQ+zw8DdE0uUYkfsz8js/b979dZg07blO6+Jof5EChJfLPFB3iuKS1/rl1G/uiM
W6Z5HwBCtIOYQAtkpMqdcsHYCV4/X4RT/Gbd4uQHk/79Bz/UGrYZXLoljYz9cH0G
MJIqUZjmkaCcL0OaNyiMAqMo8CNgMQk6SDVzxg7NZY1mA4wOfx/sOAbjPD0mZ2Nh
TpBXXDo4IQ6rKWVRsirLYncPlfCFVsZGtCIdnK6NQHJOD6gVcNvbGsdjKOItvruy
fLLPPEpwSJS90YujKuuLaoWCtn0U2j7JHqTV0tcyoVMDkQajT6jBptvtr/cbi6I4
B+BYEs3pP8o9R4zeh5YEXvl4x1qLIPSf+rmIbVR2XQBHwjPO9jJZT9a9tPzSQJC+
YIUre6426Ovc0hPJwQVv8YflLhT/292rq9hRGvGc7GgogORKChujwSB6aJFnTpqF
ResLSspIyaF7glcaQm18y92uDFP0FOzrKc0qKuKTiVo2nxtDSSZ0eRh/cZd0c09u
0uPgDuSzDHIUv0Pzt1NMSXss/11MuvbnQRuLDPkig0c8Gw1vqhcglopwTYRw3NVh
AeKDD1PLUblKeyjn5UxfzXRglb7lp9qd6OXGSGzn3fZ89DWBkdlHYviW0LG02bOr
/RhLdr7FEZwZ4Xor+bB8gWKrooLNLlNXQytgNiDfIXw4aQjJVCIlSfYAV2duxn4J
364nkDkPCdK9prSdVuGnYz/71tw2Sf65Bh2TpLo9/tfMSiydmpZgBAsVCVAqU2cS
UFmFMPOxuBwmhlMqaOtS5GQSzGy7wmPa6Ra3iSFjYflqtoGPK+vGTnPsepfP/xZK
G/Yg9LYN2CqiTcJfb6ZgTenQFfYc+6ZyMVa1Z95aB9Yj/Ija+VFSdfgbIVi/qoEL
AI0UrjkkSmDM4Bfwl5rWv23wQQJENSAZqT3xA+dT4GnhXx8+4deInaRdpB2Cbomf
Xr5/FTG1pXb37DenZBqwGm49qieT8TuaGj4zPM4OjuGi6bxJQwBww6mCaMoeuDYW
+cM9Au3/g+N/a9j3lu0FWa7F0t+IDDp6lVitT+UGZY3dsw2z2kbt0UJpLglUETNM
d6qkYLYMCJb3gfWJ6Z1cyvr2X85K/kTa4X4qCYQA/a1PVDWond9YXc4/5y6riwZ0
urb2hr8vn6XtdUN4uKE2jR7rAGb1aaK7cdwmMgrcfI4Lb9aR1yLKUzZquDc5A+Un
g5rZUSFE/avRdnLslC64jBhzKDYqH5O0T7n6LHWCvcrXgQfue4C1Rw0uupLRHRwF
kAYa09IbSU6KbBdFCSigsFNg0OUJWJXHfezQ1oKDL9dcAQ7UzIRo+Ao3qDcYjiUe
7yzIpGKRz4bvzqShpqW5OCUIXV3B+Xa7kfu36+uqXLpIj+MeWMe156+8iQzyyXTu
fjGi+aGkmzUz4vjkz9hX72WUi9LvJRf2kY1dUy9d4P6UytlRAHtvc/yxtSNowkMZ
GexqevbE0YuowY4bV9HvD26DunCrYgC+s36lKVFIx858o9a5TU3TB0o3oZ22iUNN
sMmBwqeVSLXyLz1ex59WIN8iYE7Pp7B4FxKa/Ko1tIZDJbXUr7mtG0ICXhSuCvKZ
0iEu2rp1V1ck2oLUcOxYzZxFjoCGOJA7lfLjRpIjeL1hX2yr2S3nXbyoLvmY9b21
2buykaeSOXDMaA9IUVHIrQgTeTl3UyxR/8zWQH+bl4qLDN3AU3fsM/VAFOOSX07L
NpltH4Piw5LyZuTNyygn0Wl3tB6GDDK9XkKGIxziHMbVCUrYTfrfpHBMYty58xEa
SvcxLRP3oxXxLtI8PiIVZ6HOp8M3cru/bR1RXC0U2r/uXYLQtspsBEfFrTq94Xwm
zsLoaiEXEgEcS7zEXvU/5nujrnARWBc5qWkWSrQcSAePGHpOUpCjqsHANeK4jsZq
UednPB3T8+l3b2BRtFQjUM8BIzhavxHwlRjKQN6ifge5Z5oTBzGkiwxD1+v5WOIE
FKuNB+W6weFlTZWFZMS9lt9zb3eF0rhdzXcmvr+rtUnjYW/HKpkWfBhh1+2qs9AO
FtNI6ndl2mVQqmnOd+oUK3G2H2xBdaAI1HExvNlQSSXezSCXFrd0uFFbhqLCLcOI
b+htDECzdjNlrldxFFyUxd5gkGOblX6W4K5wkfMmSyQMGDT5EpMKn6nDP/xoN4Ja
7fpbUWBTjnXje1Kpif9wkmHLWtN/f/IuhuQgre1aIlIonqwoKd1kZnqZmfyBw7wu
GNld7lf8Zr66oYOl8c0ykrNBW1T7Im+90IpLFXE5z+tquAWoU654r6oCN/ACttrI
8HEpCwf0nKyw7tYXp+j8+HhUYDLbRLoLjjPBsa9WFyPUKttQnKqSUM05qwQjVQFT
OvRL/+4+rR0x+nywLvqE5KIkyuH7ufPHQL2gGwCxQyXgulWtA2MjyNzr5wexJ8Xm
oDYr7/jzOcNQAS7n7akOpCTAikTqsELBmOT7Ja6jr5VUpTdnABQ+IVCnqxg9EJM+
Ck8Gg5izgSIoIG3q16jLPfE70vCihupRU3ZEeyniNMgazwaikqatNWuM7kC2rj5I
W8MABCKseHSl49GDPaeh3lBbL3psBZ5uuFd5jlMTjBW62XSNGx/f6gfHRFpMfNRs
yDfK9/kZETf2JN0XoX/kQgGMWqQzvHxDTALBY7StXKh/ldxjW0ZDwJpb7Ppjvxzb
Fxn0lpNPwsWmIx6NwM3gewqTZfEpBCmfo/+rDoBvxoBJv63DlHUCsNOLzDVfqWOV
PXFoARx8Zoj4AlwGK9lzH2JOEwm4oQM23KvHeAUcHtsuLWT13natj+Gd4Dahr8wo
5ZtKrCsR6jeAx5EMsOnlIXtjAt1paKrjeKlNoEqtjqp/rdybq3NpbpECNt7DRhu2
EAw3sMtBJ8qZ6EOBLHEueS+r65mdp4zGXxUO/L4wPAhJMsJlJC7RN2krPK5gOGJ5
/0GSJwuMnXRY/B00Fiy6tNE5PpI+slb2QQvG7O+Cqe6/Z+ApGpF2E9dM/bgfBPhS
xxTwHqF2U+9toECPBydLEXPPPlLIufK/JcYiJNVDB8QG5kNC894t/p+4TYmEcmHM
f96POvRCpF0ILmjASgAaB2eV1qfsmbWSZPMTiD9h6jXSGDlytt6itvhkUVKxKon7
9Dpc776f1mHxzRL/yNGC0n5STeqvueMn/WWatkJzvN8P9dbYtt4oCNk5fJFIdejE
+6taIfmorG4UQ7hVMAw9P8mPZ30TqlbesF8OOBNwftCxVbEpg2jMCYnSrHKiK4+4
i9bvolwD9B6/r4AiqZmL///PCz1NwZwnONusPeAxDzNlVPYzLslO2SiI4D0Kbsvv
vUO208lbZbMOIQyirC02JSeMhr+lCiUQn8pxUz6rL9kb7Co7PIclsfKWjYJKdQ0L
6U8ElSvtFudm+MxH0UWcICSfMLqJNyo52CTwJDu/XL9XMX6dVlMe6ECmh23CoxKW
+NZmY5rjchLUV6byeMQh+6eNcKPyP44u6Z3HRZi8OO6Lmc2MOeX77VUYX8ZvCqIN
ozR44eUc5kiIIL5ir2k45G414/1TuY7R69PheDUFLuUdpoCl4tBcOVDNzM8ksiS/
j2BMsoM+u2KReQGPwTVthIfLfmUcZAg2HE1bbkDbRL8ExLbrVOcEhglDXlhOBoo/
myU0Gmdhwc78WaQWRtbtNWCdENkRryd/Awpt+g3BOwXJvKQbxvsxFTwC6D+4uMVw
F7hAyUx9ST2ar3nmV1HslmZ6+nlUD2vc44mwxCvlLc87Pkm0z2LOClUWXwqJmqDz
Wl92H18oMtwnBT404pinMC102WEXywrKHNICnVuOM7W9Xf4YRB0YK7ItxgI9m0mt
C7e8bir9ajL+oS+oF3n5gGkT6d+GDpjgPe679lOiyif1P0UjmeJ5DXJHUVCxnJfi
yrZFQguE9PlQFpP7bOMn+I/BC3+4ppeHWYshzvnvP94XMN04ZWXFOiBoKL8BpK6I
VrH0llVZbl09iv2jNeRJBAwA03fu5HFP5nQ6xSI6pfLyZXyqZR31TsymbF5LEyaJ
KZOYIycI7HGAYNoy4wkLAyk/KHKvI0JEroxgn6h//1rW43ne9Izqh+mqe7Vd541G
DXwbI0sOWk8NsqFBe4S2IqD9DGfzYyNy/qhq7IXObQmwBgoCuRWQztmZQJOCgyX6
BSMmWM/sTWcGGKTfMRoY8pRB/0jayrDh3GBSWKWb+Zqsr1lNuqH55LnHlDXvHDeP
yYN4AdPkyoc4XJfQ6umry6VMR6KsiNB52xkD7q5CmMZLzjrv5VBwBNyvS5xD5MeC
u2EQaGbuPFNNmYYaJJmhL1LmhESGsXd0VTh0xKBpnyBEh9A91WfUrJoDxTkQNkge
DcTpccLxpY9YibARzsB8adHvkNvLnD8YufVw5JCe95MIsNt7e6wjd7D9kpsxXotF
kzCfFplLhxfofWr2fR1aqtCMd+qpRiKg5+rDxWC8tEBIzXCkiSlFI3aOCsW8f5M3
Z33ouSFEZdduhfg+HZ2dnRz5f5Jqm5/lAy2jhVtFOJrc0p5YHjUvCXw3HqZrXYKn
fPcijYK5PcaPpLvpPAzA1gJrp8YqYpUKFqp4YOlFxnwe4mO2XOp1DOvHS9187i6R
kldxaPBUjOkFO1l2Homkp9qCxU8Iot3me9YViw/L+Wsz9ROGCdMHpYwu4e+olnUX
YXiLGXzA4VfscBk1755cmr+HkLFzxl7Si6OdZGJIs+c96ua2ecwqdHNsPhU+4nqX
AjKd7Gi6XxaHY6RrT1knwIqbPM6PCGK39MBsYA4k5dKrOQ2tFD3oJV9yrM8LzYge
tlqC0OV9S0E6a2AI9r963erowBx7+ZYec+iHnfyAQvscnDQaNaPsZoO8YEXuvPc1
XrJhenJmN6z56lWaxzqBU9UVNCy7KlXgwe31rSKD/OSzUgWDsFO6IRqcd0advVDg
TVKscFgoMBHsfvvjM/zODdJou+lXA2V0pkXEluvWsyhWhxPkQPbR8MYa/5egaQAs
Kjxx5QGcB/0TrmuVm+1GKx0LsYKEwxmiba8Xb8XIFRfqsaaENND5kPdZEqpiMfKC
oP2JHP0IzAKubURYpZNQS6XLPHI22trGDxPu1X08ipK6DRQ8FBokzXsDAS0RrIXJ
6qtwonMNBG9yswVmhe65pb//I7aWlayNFE5KXyHYznKxxQtYip6YcxIzaC2nWtef
iFaCrmAUOPg8eo3+0uKX2xE7zSE2+/FUUkgXX6RU8OVzxcBwKn5ulJQF7Qe7MLYL
langLwFgLq1gQ4I6m9mFki9DgIzzcnRkospDmJyLxltC5hK00IqbtkcMo0RUjN4C
kYwk5/Jo98njv2JuzKTJMVLD+7obMYOQosokCb7o0flsSUKnWQTJ/bxHwdUFZQc3
ha/KZJwClvPHgGZ5q4/nD7IwJhNP4mmlnGNIgpc9aVuSW4aSt0Qcowfdz3ehYyQ3
HitPfc3fsYxKlNrckMZXVQtm/9wDmjiHGZbUmJP2Sb665CNucYo5YDmkpfD/Zrbp
wGWo3yiFMZ4wNsaoLAqbEshWhqsCbUoFmteYG6Pxro2wcqq7GptbPiR9w6V184gJ
V97Vkfne9zgf6TsmrVhThNX60P6bxn63/ah3P4+1uyZ+qfu/eGKIom8FltYLHS1+
PxkJJv1VccAXTfez/8MJgjNQMJVx3aNKmOwo4wsoO8hjeuSjheJzq8vwLAkuzbug
Ji550LvtDMddkFRdv2jWi/r8U/GiiVGNK4ObP1SeVhDlZARuimO/ZnHYbr+u8NYy
CBpoEto6wRjM99mCC3WSODfGCMj8wC1/GFBJCHQ0XtPnZWkLwkRI39/H/Z4lTmZu
S3+srI47KOFuCVz3HVPst90lEykIPm9BVrI7p1WCbuT4N/0unAXMS3KX/4k9EurY
re+C8ttzA4C8tkzKYRlS25+hs0VbunO423HehfnONgfPReZi502ilQn5mZ3oBseO
9AJhCBaEHoCe8dRo1M5uxbBxHu8lSxPQowVYf5XBTCDeagsgSSt7YjX6veo4OmqP
0nIuuJ59WBwrokVtyzCEPnU5217kGSDj72uCZYgDdBuPK4zbuPdmM947iTAWozV6
9M8SfC9LvgIe5Z9HSYxPHY+lZO6QGhmst55NkFnFIZx3qpJCMwAlfU/nStLDx37e
crakrb9sdNRl7ncFZoEtNIZaPDQH8XRFvSThszsmf8Nu7NYLrqlCO9TCrs6Dxjej
yU8We4vFYRzVhk7YoUv2OqaNLIcDjMHuTsNUv6AulMKAGiqc3fKE7DOU2/TV82jF
3PxRGNFYotZ153/GMo48AuBa14aV4i/YW5boQo8aJngleu6jDBVO9/LG6I8FR4LM
mqdd8UFTjIFMKDNhMNFl5KCtK9mq+UAA3sN2+nrLY/Q1A+iuXmElHvjJBkqHr07c
leuJjCH1GYLNAhIUFxrIuxH8Dlgh/Ab0dgK+FnlQreP/ctneH3dYAl2RV5QS3gM/
nqiJEkbhuGRZ5dfX+i3Eaf89YNlUU7uPrkxBQYEExgAXxh1vYSoYsle5CKVMWfND
PboohDuzu8QVRN7bVo2Zif7LG3qvo1kY1LRQzqxllOWlieoQI3t7Il7Y8JH02tSH
5Hh/x+jjbrGxr4C+udJEax82QeyCuURKPHV6l+Tb1+Zza94phAAMZ6pzUC4pMnUO
6P7Rcsbv7tL66BpClc1wg5d/eAXWSmF6TqM/iNtKgEYilp/Njn38VOl/Fw6Zsh74
yIu8faTunUOQj8A2alFB0ZShvjIivEyNv3qvoVZXS7+V/ILJQmN4QOKQnOdeeafG
2oqV+WiOF1QsHBOryH2cXsW3tRk1zlG02zpqb1ODwFiDeu2iCZKdKOmYav3xEMza
gG8hUBNGgvtw5QGCbMDVvAGE1Meg3FWyqgxEphBCY12jFiXwvv/ZM4TLgbgXRkvY
YJVse4cuteaHDzqduKepPJ4GwXuq9rKhkNOdOr0MsMYVt900xSheog0cYpod28lf
dQU23xCbf4dcWp5sqRRb4YMEn7FeEfWk4yqIZOze/nnMA1XrvrTnBJfLgTj8WVCE
5bhoEEoPsrf8Hc+SwHrnDjCeUJ+7gfZ1XyzBvR8xbtSO+lhJEYJCBL2icbxM61im
M/ArXSbK90gIoSfAwYuCp9IjHLKYCoIoAeECQCLUsZ7N9iJOt9PUWTSR+BYH7I5x
xwIBqKNDnB3vQZoi399a+CX9k3E3qOLBb+CTjs2JTVeZKQooPsqYB+XyUphxaGr3
MatHT6B5YKaxLMAZ8YZd8Y2thXmyP732d5cxmsjvwH8EQj78JKgeoXHUl0kTFiqO
J16VrumyV6Glt+MqXeOTDEGcyWxyWKi3afpALCQJtn14VsXfC9K+lFvnX3wJdgbY
n3omCEf9boX/IObluRzK1AWVL8cWFA7Cky9EZmvKtIkCFxcebvGadUQK/K5hyugq
1iA33zt78a9J6ZsRLYc5qdgKzJuhI8lrZU6fbDsum2xptRTi3pLBPAH+f/z6BoaT
ohSHs1NwsGlCPur02K3AwjSD8bnFMurI4ZtzVypU0z/fxxbDAVrCLUqDDrCxKS9d
QBLwEkSYh8lnd9yfMOSud6y6ypuERBSb9nLYZltTrAtrCb/LokPw5vSJo8GOaiRj
m40oBWoquZiofC64/Ht253Xt0xpOdGVQuBxFhgVbHqG67fYzsrXbrejCOCPqIYOO
Ef7WhUYOUu0nil6VYV3O9ymFlslQuFyVg9VqDHBPGsCoHyT7/p1PzyxtOEgmtifZ
Qi2GpkWJ0IaJLiZfIZ3kD/Je57BTiv14MrvPak+WeOgnVeN3B+IXcOVl0MPaOPme
wp8XBvlW2SNK/XAKx9GSznS7f20I6P0eKWBcNFv1FOn5x5G54Hy96sVYo7uwdiC3
rxSwttXT/USyqBpjOuhzvaUhzEDOTrKuJlWs3a5itky3N6EOeNNN2YZdCPq2r69p
cp7LTiGvf31oEqRi1YXfndjFAtCYibDR7r3g2IAD1RH0XRcRvRZbb1+FLpIUuoOc
Np8XZghKWoDcCGUOxz/ioUTfqq5kZ3sHtxTYhS6tWxGbr0XFiy75+X7bp0cvKqjv
nMwQruhbMi0x/LqCUbVIA+CsBrAAzqBaOziA/h2yJH3lwbP0C5+WTB+b1CElxo1S
ieGeirKWUc5AoeZ/yeCnWv89KzWtVz8PxCyxZ7eWFb6OslXcPxnjM45Qkt41radx
gtFT0JZw+DwNg+ILXLeyUZxf3NLiZ+aDJB0sOReSmt6q3jWLN6lXDG3nJDoqiAEw
WEpPYHTcOxsQ+IkCmVpXArCKRq5ayKaV960vEnSb50aLVjVe5fWLZUDVVNUl27SZ
G8Vf2mY5lp+oDtre501lJxwel/fxq6EJiMjy0mj6nvSnUQ5X4pxQbD+5pXz3ESc3
ipOZY7BmHeY7p+QEiQbAtf0lkxNMDVOtzI67nZ5yj65Dra1IjKmxPcdc7sfdwJw5
phi479373RJf8GOt9fQse+A65d68oMK+H3o2EXfj1eajFJDu1drwog28Ro6YtYV6
qbnQS7kPLiM/m2tK9G4cjfez/PB0mo3uiLtV2h/5KGSoKJyxJtD5fVU99gk78cUh
ZJnRdxWFwgjHQV8lT4JjZVNbn49DmZQiEiycTlCYvUjvgvWTXKa2z1/6j40fGIw7
l/RIoVpC9p0Eq/bLIjrXRiF+oKHaG74K/lSYfv8/mP6+uAVth/SIYfs/BntGjT3U
4zhQG6YDG+8n000Iv5xUig4FVVakMaMKw4LoKJEcPQL2/J39JyhJqXbFV/vRuKLL
F1aKC19cimVfSo3ffA2Zxu9bC3r/TXna7fsb6Q09L+WU/Q0Ww482HqwURhdAJjo4
6MueScLTjrBnc2V9u97A6mpwpKj/mQbEoYFX6xJPSamE55VJzS61svBz40YVM9xR
jMcsr4lS6bazjmXwpvdXL1D6I3BaFw+jzXbLPRjK45v7+ztqU4ktff0YFxe7k4sS
ZZoLx4AALRTLDHwA7x7yMmfYJV3wiYp0/NlR7FCvyz7/5NAA1vuM2ug6QmEjLeTM
qvMeRqYvDXaf/jzJGq1ca+UuIS7JOyVY/Emz1CEgbikYNjyGfis5Zk5wATt6s69K
q//KCAuOq1V/8fWo5Wp2fCBOvUuSHk3WyW7eVCviS7MwJnkx1Kq1bAuCuV4qntRa
/B2m6FVQQpgeSzXE+PWB3yLs7d2kl0oHpL/5xpu9C1tkBsrKq3H7cFKS8bbHPLgG
LAv5DHH1FHy/XNF1AFnZWURX4zd5LhmWLFESv9eiuBgcooFKA8Ogt7Pr27SSKQqH
8MJ/Q27IOIH0aDYlQPH1Q90a9f178lAg2uIGAAVX0+N1rmK21s9E+wQYTB2851I/
EAp8MHFP/pef8Uv0Xb1XCcJEloMP1eMNC9diMN2Hlq1IaabMz4aTN0Qwzlbu6wOe
9Q5WfB/dBYf5qKN0RDY6AqL3sum25GcACYNxggg/kVOfJgdyC+Dw1VlxCYpReMuW
nsMyBi20aoeIFu4hVGundewHxhNdm0psXZkxqKUJs82rHunhZ7VdMJZsElagv69k
oUWFN/gYF9Y6pMlL04rj6J9Z4UAaT4pNdmlg/y7kWdEbu5CE7O3cakZ9g07/Xhfg
sfdbv8ZqIupWUn8uxqL5tbkNfkvp7/sqhnmpnrB+BRUihJhD5N8AsAdeYFOsSz0l
ikfeDqHbK6IQAzJHNsJrARhOPdT/soczv09E8CidBuaMfKmvhkmQt3/ldbHsczD7
Dnjmr4sZFKY9AGjXlck6rgNFFs46ja2b+8Ab0NrTP3QKLldUvs18/hZD4IFyLTTB
l5yi2v/Qb4ayW2sH3EE1V4/vbAk2mks89mUtVBTAGUpaZFYx/jJnLFAthFCR7EcI
UaPVthwvqN6ZLlimGstyQmMaUTndjchCbzH4M+kmPpHnGQh7FjN3ZcZ8OkYuvN5B
8gaEkg93Ivc76UWxpXqAb6Yuhev492FB7LUOa5qzR0ekpUOl4lACgGb6qodEjQCg
Aw9l70oNiJ4jdf+MSR9baCYneLHlhDwPUKU/TVgncRcHQsxdArUtTiEcOeRZOoji
Es6T67PCLOI+d3v3zZvu4hSx4NNCv6qN6FQFr7hU1IgQMdl9emwPexAzf+01tRpB
eD1AB95Xj68Db3j6OxiRP7LAoIxyVyzoQ3C1GbY1PVxedwFpHOOAKNrSbbmAZOxu
h/GHSL+UgLzmxYpXltDGRWC556e1eZR5egLvw/Di82YgODFmKUfyTUvA2Sv64NTd
9lPWXKe7/4WfqzYISVOC2CoKpDIYLeQHZT763Ll899ZndBm35pyDhYv2Bja4KSSO
qvSzRj3E/w8YsZT/lk1RmRpnlDmVKFGu64Qwx3LalH7hjc4mTs5TM+gXmZiorvYU
JfTBwA/6hmABlJZeagQJHyAspCtrrt/GEqoqcpY+8J04a+x1LsydlnRrDvK/nrbB
HHaowWnNdBrUXN/dOd3+BG3SVQv3mWDAhsVL8K/EKjQJjMM4Adz0/TXcGncZPutv
RlI9F69ceJzknTUJTqSsnydt5suh6lFH9FltpqryXQ9Lu73pBrvXyaY/iVLyC+SA
mXw0Xwn3AF+rh1gOkExmxpsrRIo+sDSqrZKXq8PyygBS2ulJTA7u2Ag8EMpGa8D9
wYyRUyqbdtDBK5h6ZodVhKAs7B+wcLmq8sbq0LRAmIFWsBaJWFMM9KvqtlDOED4k
czFEvzXPOZWSb49HHFTwiWXlpA7SwO7JeT8gIwtA0JvFMEMsVqnf1n50Ays3rg4j
6tkIDaZGzvt5B7zsNjf2Eiuq2R8/jsD0sUGB0aQFJQTeR7Va+sQAzi8QU3rwm3L+
5StuvJbE4MFkiCpURv/JBw0Ms8eWvSv6sUranrK+DR0i/rohbB7M/TwN0Icin99y
tz02GLlsAcVlnFhqnIY6M0xEWfcNylcvR3fpIuMkLiNWov1Yr5jHrpSD0O/a12aQ
PeIARBXUnd3VRPaQVvrY0/nDVxGtbTHH7ktRI7kE+/0OnMDPIY+FgO9reU1uHhZi
HLyAOfUH9QNmOrQnDHWdbOOhq1i3q2SlN4rcYvcyfV8OagJvO1EWgK/6KVJGlGZi
svp+Z5UgEtTY7eFb7kU94qBiN45TAzhySYVYPBON2DlIV0sdbm3/Se5+GrctXnHh
XglSJkZGJoi4mRgSChHqAZzJfc0LNFUl+FPBUoyza4mDlALoc/A4npt2ckaeXeQo
O6USmNODTkaKLvNk9dIQIp7QLt9F2c6h2eN2+gfhM9XqU2DkZVdpW2j8BqNnAEI8
MvjPDDNjum3dQywxGKMWq5PLI+GVeYmAmoWAAJt3iFVJN/9XYpe24Ve+xBV7FG3U
P2D747w+BQFY9URQc9mlOI4SyyEUtBE/8lOjf1WRmiLeR4u0mu/pMeYmNI300kmj
YTztIe0IOU55KkRrdq+0BHb31BRKYpLHE6AeGH5LKeiuRG9/65ctwzEFn542ltLw
GYLBxEi+XETxCrGp3so0G2cIa+KURSXoxZAVUIScEbok1bEz8IzPKpF9e1ZK+UgJ
qHW7JaHoAhhpYtGEYraxcjTEAeBhdDeTxeMvVfAnJ5GbdzijtBCo98c9TjDM7vbw
dgdBMiTvmAQZ4/K87UjnLd5YtXWVaJdVKVKkEwjSuuLt87oLoCUIfzT03zomea46
gVv9rEMKSqgfAV5/fmXBtlHXMwreBThNgK7OPCK2ueAhjeIGvG2ta5anhy8HwaJX
clZNArYAZivWB6HFsoJoxZ13pHcMRrxQqeYSyHWhCQvT0gH4j4GPCM4ScdMnwIoO
1Y5haMmf5x0Bc2LD0fCgEB/PeRSJ51c9Gz2itRanIQL850HohbKFjgfclEgN+FHy
A5/MN5XkVTsLCJPKdlx9lHfeLR7dxAYuS3c19LgCwKpjNPMjhyzc58GHo4V20KcX
jtkg6Kt31xkelByduMbiCHggqy2pVMPh29VYh4eCjFYAJBpWcKG6LpbqqQyVEgrq
rGIjXpl5onBAm4SUlImtuEzwAfWYFfaJ0fqHw4kZwLnrA4oWrB42lzHbBXzoSYXE
0rvreBhXiiVU3TXvQuZMWKeky/6SAFIDo/xSE+k+yiftfEHKciNQVYGq09sO2f+I
vLbHNCvRvHIfris72gGr4xDx/an01dOC+KnNpypTjQBklotB/HgeJ3wZiwvtAAXO
/Qsq1Pq5ZTtqGebMS3wpilgUw9K5tvj9iYa6UxTz+ShncZYCWs2A+KAr19GzAIbt
jR7AHF85otK9EtScRjQLwfzQig1/8Vddk6f7VpBmEKbzGcpsd6/xEDj7zRBuHGAx
DYGAUFmuvEmzxiR1bYR4mkF51tEC3OMWfSDFl2mZ5GjgP33rRNcS9VHfl8MbP3JK
fOR8fSQbdtRi+zP8aZ+c4BRercPYn7kTEeNWFChQ7k9mKlNG4pMHFxOwvhosE9fU
0/i/zLTrQ/0In8/dH27QiExsjwnjm489LIA3T531RxAj7AJ8P0l4H1YjQC242Gvl
Q935jTgQPMjUJuron+oQ1qoLjap0SJJmtT89JbhttnyNs6+GzPcKgFW06YSfXXYF
LLmQ8UW35dX+X9XdK1BptkS//2BLQWx1i2Bnh+g+K11lS8ZCMnKILXMqB3xmMu93
yV9zNEaHn/E6osCkJN2ihtDZwTNo0hLfd014Qun5BCYDksYCNm0+W0IX6bzSZE6l
BTK8KwEKkJo/DsAlsInXblezk2IQuSQaDNbeUO5bzzqcOOdREN6ncKIui+9sLxRe
eHp8yq9VoqWaZH/V69RtskuaAM7Ow2gcvnHsbKZgF1pf4qwKK7L9SFYdxgsjlLUZ
uplUncC890akICxzhXq4F+XPYcqjoca1Iqn/2ZhqeLuCleoJTCsrxaxK/D7kYq8m
dher2GwVr3T3VqN2NRqaJ2tngxDBT+vbnfUE0KC42dYnj3cV6DTDEGKE6VG9KFsa
kjpO5Vk/Ej8je19oMYc22gshKJfGf83I7Oh4874BrfN8hHuTQOxMCCkITcD9tt2W
bJG4PEF0bc6dVU9HHqpF4b11jS1bpNpwTwk7R1U+p26mLKoc3nkCWzQYhayYmX26
NY2W10o2zF8AwhRnFGUh+buVdYojrOCWn3nGaodOgSeSPTszvNXwzrNzA5Q4HYPJ
wf+L9BR9C90OiAWlzkQVjfvD12wDTk14HlxxKX/NbVoD/A1qesIqWols2vqsQ3P5
Fg2mc/znKUsxt7uoaTplJvw/yJDASTDrCZ7lixVwB4nWLuQz2pd870ExIttTlDgE
IE4Uj6yz34lJM3iGfYvuZL/SS75h++xf/PaOsSfnG9ow49tJIRu1U43uYWX5pMaB
mBzrTD0qRTfHXliMXlRP9CGfzeHOsxtIvd440UhqasOWEu4bXHVLQXULkRcVKGdE
/s296V79HslPsmacNoulMMOzL04BQSZqiBbmth8Pyf7TPMWJ5J+G/wgMjp/q0jdV
MqNunsBEN7Rp8PVZdteUnDktKoZaCWL7DE0BuCpzjQ/0653TtnRoXZ83FoRUnSVv
XLAVbhKk3aEsnRMjQA5SbuxtAQ2HtKahLcgEVvv4XX2CvzmQtZNhqO7QesDtHGzE
YDPSt4lkT96Zc6FVE9imumYMvfhwj/Z7VHEN72Kzc1LXWulEDBdNLTPd5f8g2VD2
bzYGkH+HjA/RNL8vdyhoKKLe5lNludN187gnofX8aMzKsFrbXcPrS5VeQfOEIGuS
7oHQpWGOHQTaZfFKeVzYgk34ojTSe2jI8gkBG5eMB4I4Rv99Vf6zDaP2Q5Pp5BJ8
uOL4Bk/Kesd+2dnGUC1jcYG48Ul1CcZbaVN5JwCnQdFV4K3F2JNgPvlerFhBHUrN
pBOrSiiPrLV6SDgr76WSyEYZh3biWAdZ7hDJlMeyvgRyr5pz7iSyv2vrinG1Xg9O
oTpzQnvsto6cpiFLdKSAE1sGBNj3BqmGz6dshYqjAlUyy4iAN02UyOQICqRiL/XJ
QxYTkW+ujEuTpjwrKolkKnSYLo49D/wm+SLcg7EQ0ZzTdEmb1CVhrVnGs3PRNgUZ
6bOWf0m8OL9jirUtyPjIbtD9oTrlwQyger8OogK09Y2TkkOt2FPTpXSPxdcDOgHD
lDlchnAdOAJV4g47WvsjupaOW/Akk3ijafQk/WyLM1cEzlWiFIQPfxFl9ecEWfmU
KIP+V4f5CYdkMS30jJmEI/FZzOe9kWE4ApF2+JVkcIsQjgXzjlY+h6+DitctsCky
dvfhgS7cxwGLYXD3YwiGyPsDhj79lQOwl+3NR35UD7YGUYAVM1GXm0017EkX0blY
HXbs/h6oMIQ7TQ8sJ7ctwxFlmwXCG1FHhlNM3Z/zFhB2ZglDy0xGzvV2Kv17YmDK
kDsIZBKjFZwL3b49Xyhdr1VxHv7btYSkyGpl94nWZj40R8bUHk/YYiv7rEd536W0
c1ZQLnQClkSliGr2yWS6vtrCTiMaYYfSd2TrQAump1m9mKU8qzo7qMqGCMww1Eir
SzhQCmvLRJd+CTlMJ8SdAV3rF7uK+thuqSRBBnSvTcs6oCFNe1VXkRumovLEeRbO
dGCCUIJ27My+25OKF5tQjOOJnN4sVmPLQjKXHvr9+EtGMgreBu/5KravZCPinzsc
uhK5Y4Wq0131Y1HaN+4kGDk/8WRFiUfd1odQkPTIRyZqlo/kR0ZnXDkQkgVZSsZV
xY8sY6VDx8NEkEjL9nOhrHb0NLKaBtu/7Yw//Xlc6qm3cvBebTevQQXgPH+VLwAm
mj3jquds89GWY7bnxcRBzA6HxY6QsJ1Iv4SSWO/+hwkeEyDchMbXTdlre2YtLZea
GUxNJfe0CwHi+BxgIMGY36USjUYEN7xq12pH5aeaUsPUar967URUZ4pwg/rB0uwp
OcXovTZeRcl53Zg0ZFNrk3ui0P3VHcAoHT0SVerDSe8J2lGqS8pzNMrbaX5AhkEn
k0DKIGOvGXsQwtx8NB10iSM9Kw0vUhzrVXmlUFfRqqZ970pWPjgJzY/jLRpJVhOc
hZQHNaorCCl3OIzNIVAeMGCP3NT4ydBnxYfTGCMX6aWO48HCqkfK+2VoW7Rt6wif
HoMtkJF0HNMvGma5xkPIHLpZUUG41cvhOwrAjgImgDIYoQ89EuYoRqYbCk6HG51M
JomN66fq0lJCpyrg98vvdYjvNZmsWSoX/uXdQdmA1vTApdGgknBlO61lmfMC9tvR
96homkfU7vTVM5Pggl2h8n2FPaH2Kf5G6ztFmd9e3f9x34UAAK8oqA34/erqDVaN
5Xl71OaldPZHoeBMw+9Rg/XWrlE5xG82TWrlayId5T70l+eEd6mWcghoMJmUsKvK
OjHnFTxDLkzrh35d7alhFsn8LNgK3MeEV7Bhd/XwUvNScNdoVUpfgjAQdqeEvVe9
vW3TYuhyEfawDR0H3au9TPWqwkDyhTcV4Gfz3vLJeq/SuX+g/nlFrGQHGm0Ig6TW
008THt4aND7CXpQiLNE+lDzqWVFaD3YOWVmYTpXYdDHHQ34kF9gQp6cYnfDR+u8G
SIypxIDjJ+9MipRqUw/QsKhxs0gUOLdYT1Lj81k267FYYwbi/O8pfE+JWl9nDzrM
c+0FSin/PwGeFGEeE3oz7kCakix2tW5ZMAo1ajLZlRGVHHDVPz+bTGbT+YUWhB6t
1JfK3/ysScFJmf90pR90el0RFkNEEMKLQV5Ln6sP0pmR2wtStr2RgiZ0DFnOM89c
cBqkXJ1d0Bz7RFvOd9LXLcWiF6X1mYd5V9g2/6/JH/xaH6iiNJP5PJ0OZSMK8SO+
kQJYf5j+bShoscfPy0H1q4ELMZ/Wo7G8Igb5YbSAoOtgK575aQSHG9wrJhA/1Dng
ch5nHcby/CASZeaktdMh0W37BEkIIziuxhyHTe5eVtcEfg/FljZCFkvs/TncYJju
uzWamJxD/ebWslRUXdWToRnMUfNCJUqlfzfSbJCanzs9NnExQb12vF9WPg8mc3hb
ZISv/bBh5Iv3GXRwn4RS3ebKYj5xzE6EVGCxbjoM0/gm8eXLHT9UZgJUy8PJD8+W
lSsxXwD51IwRS+X9tU4jVgr2dPx3fGUD+tIk0xmApf5cBVu92YaUBysCONFhng2a
bkVZp5EoGzzRCg+giupITlkSbWi63zg3WKI32+DNwe+i9XvowBUhBdr4ZrAKPRL1
NonZVPj2aTyIQmZkOfSrDpUbnNo1McIXrDIITBQDlhQXeOrZyyeYyVYTdxssePc4
We7ufesr0Or3k6jzg8DNwWiubF3coA9B0UkES2yY7guJmhSAKOhuwDCa/qHvPspr
qjK9BdIxGSlNvshexoxNvzxNhc0Sm9fr5/aTODBa9Lqdi1JCnuMq+KD0FK+JhXrW
MKoLUm5CVcxK6R2lny2oJ7TBFGFx8icGUqfvXOjqinLOT07++jmd9QXyW6fdBB8l
C3Ur/RDNFh0wof8oya17Co5/+jSoK4bIwVBpDlmMm5o5Rra08O2kbdJWomLdRzGW
Vuyyg0gkFwSweNKDWlY/BDoj27VFBlZ5fo0YacKXInzvsvqo4H9tlIFsVX76owqm
Z7sZAv7Evv2mCbzqbuZb5DbNGKV/VPTxhhESMrmekT31aqCAcJ1k86z17z6aWvo9
OxnLWgMSrIVQZ8qSe80+OveZPL88dmwAYBo0QdP+Ls9Ujba8cl3s6RLOitS18Z9j
93IhOHI48gYq8J5LoHwMCoHm1fcyovXf/GisO90xerW8Tddorccz1yboPbURgc56
6jZF3PyohiX7aw2dPTURR9ATmXPO+DE0CTseiLlKT+3WEfOA7+tOzNC4nKOsSG54
hJe6K0xNVi9HVAF9U4rJChhENE5lKDXDrNvFrc44tOP26sSRj4n68W2TfC9NhJ/0
2MIkui7XZVQMcBtiuBAvYtCLWb79e5sdqzfDG9LSOzx/ZHtbdpngvVCMgNQiWnNp
ATQg1qoLWYj0LwjGBlVjRaHqYfUjIyZg5dPZdyc+vylOitBpYfQiEiynpHce9e4i
wcxYilOekeMKABZwUlWLk5xXQIeKe7XRgzLmQqJCORdkJ5xEWjbx9G8mlFqfuYi2
tT3lblqasB7MoVvi1DIL0YcjKfXsrr+JukSZwUSMSI7620hznjqnz4oiICAWX48/
4szS04pRLxr21omyMi3GUxduG++/ybMmK8qFImVSQudPqdqETNgcrC6oFI2G5mi3
kiB+CmV6Kju1o0/jvEzXnCXqjDSzZ0TqyxYZ2s/RIGTfVB1LktqLB062sexHL9pG
VdKq2bFMWbcVaydaS9GJJEhH3h7q6eQxmAa+EDWXpql8INKWnHzx5TN87245l81a
if66riVvwphmn37bg9ez04dM27MtwRzK254oaq0TRjitoQpH/WJLdZ9TXWrW40fG
DbU/7hBB01bBSO4NaeluHo+gYPmH+s5cWPmkXM9VwTN1YGBsM2Xc4OHcKu12Sdx9
t31rFcA/LXsDQYjB1Y1AHGL7wUlxfNO2ATdG5MuXkbKouYZNQycpLFi6MQudbxFD
KvPhgghoN09cViBd/FBQs8vGeZNQ90kbIlVvGNZDjM13/dgFM8aq8PZ+DIbcwbYj
tn+A2jShyoQLqT1wc0hRYnnvxZqU80hhAdH8kABZ0K/nKgjHqTqVxdODRU/2oyjh
trm7knaPzan0k5kboOO+0bFnXfp9TFtxMLYPbM5RK3Tgv964dOqhoZM1YYcw3YMu
aULfcCRFy6oYavr3PMfGtCfb40BYPcG5BmwIhlM7OwOQgxjYkIjrD5YhQaA7I7ME
XC31DsdWQNwB/RWIhC49B22PAbNGpSQ5Kqy6zUyC/3U+uJB2exq9IcIfVzzlwWye
xjoaCLJ5260e18FhgFO1Y+0pZEKn8bgXxwe79XSL81HuPPFqLF4G3bHTPzZ/37u8
eyAwqW2TeQE6hV62VLgFEX4Yg56mAE7pMU01Xhh05c0tupaMCY+hWdoKuXyGcVV1
RpeWwcBS70cSENd/T+XlJpHXjEjrpZpWGxSUUpIoQSAjdzM1OAl3hY/citl7Dyq7
1jLp0vxqDhhDuB7YXJ58PIXBmphr+AR4ICpPn82FuATZGQdJ8JPITlcIO35+vbqy
seuqT45YnK9VKx1RNADK4dD6swFnXjllFrFcBJHx8FwEpG1JXOnbVktVtPBTNUr2
CC5W/HJAJdgTt3Ai7tUmlkWNA3zk699Ym4zzup+qrcLuC0rmbe6OoRGCY07ErJSG
SbYIp9YpscAolLPsgycKyhqrhfDykZhfGW+o4GyhufG0xdkprw2kAVT0ieU7Y4e8
juIROqh0F8O1dXfyqqDKei2S2T1qjQIo2qBfYp8OsWrIw1DsQYCVicSbA0Bx1Dix
Y7mFmUevV4kNe00cfg3WQ1fa3I7x8si5cRFuh5uumdRA2B08qqTyKOYorX4M4aS/
2Db3d6HjL/XxDFuGWLcZGyz1LqPrujJU+DKB+os7sDJDSmZ5subtYk6+Dq6Qommk
JvWJlVBLVYSwUlVxerxzs0ug6qXf8q2JlrWxh7rj8Wx5l9+fnMbtPCxjEQBlElR+
8WlzW4lvuFjzDTznos2nNog2ib/AEo34Z+qeDLq/fCWhTD0jqYFLHgRgzGEpTlhi
8K9G/UPemjO1H6WK+a62aqSOeGjwHuWv9aBaUKKPmduXRLtcY98V2xlnFNKCnjPV
7nA5OZ4m2eY7UvTeXfepDD5uY+XMDaBlHNqfRBYfOzy9ZeoNUCWh0TrDm3No9sx3
n8P+YNgBnKG26hJuTF3IZKKd5w4vTUWCDLE6pc8IB7apFfyPwgP1R1y5DB/88UP1
nV2ouBGuU8i/0Ft2L2kKfKT/mI+AE8VHMbfjncb4zSR2LoEKuNVu9mvYR5gPyGF0
dMNmWrwhnPmVZudENMuNpCtYbNzQJbDqacmBGTeCuIZDy6L7rk016g+zUsW0FzjH
grM/kXwsMmgHGmtf7PoNTj3qUmayns2OGgSyjbOWMdTtt3CUDFzuF2c14+Cgqeo/
Sos9IrQQDpeC2CKXpm3Sx9329qM0f/iijv6nQ3TBuGnSnrZDP9S3IkVWeK5U9RHM
wzg3CXFt9kOSN2DQySN/JtgHojBXhszAdwRwk/cGIJFEwgYAkdvKtyW1UTkKTv/Q
Adi+/Zdji7k2wkYa/xKRI4Gsev0EaiRZMmWCPuNTuO7pfx++2cj2E1h5DBBHjpqf
aq1BpYZsecuz2PwQ0S715U/trBPqjaTy144pZo5/yndqXFYEt9x4BAecOjhQV+G0
i0Lmh/laLfu+UxcuxDX6C2/QsRCGkAezbqrPIW+34qJXXf4NYoqGkkrcaiP8VaQO
b7fkO8lWGXWHqQ00eP1qWN4gNMrQkSvcJIm9DzgxSHKJhUDFsL5+Fg/JVETzcIHi
VyL96qx3bVWdc7925TaeGWcD452XQ5nl8btozLI878xQY+/lEN9RTpM1jEdFpkWH
bLeGanTO4WgDvS//FWZQmwQR6wlRoA4heGyXAdQ4fwCPx60tvSBZRrMS01Kec2JF
/b/RqM4YgXqQUYh40+fEo07hgSYYx1shS3xz3oOHq/i02wPSmY8L+/h0GD+XMpzO
xTfWcresw0/nA9ijZ2934Q17tkAXWw4Au5sqXR15koHgI53vVNi2sdInfoTjprLa
vP9J8UNMfbA11Uc3NUKKw9/Ly/wvijTpENetZ7eJXeEFHmmt8pZsZ71Y/tFB4Y8y
Wh3XdiNCktDNeypFo7K69vKcZUSEJOAq+foF1axg38qBAeoagpwXlkiljPsd/aPd
oq+EnFPlrJpPfBkR0Dm/9fA1YAjOnBL+SZueg9TFm/jOhSzt7TCTQWz1fL+wSvW0
JaXxMpv5Ip+AiXfk3z0cm4AQhnIY1Ae9goMpCXWQ/HveEDhkZMwJaXlY9d9zludz
RUr9+d9JEDU3yEwrQtvflYqeW3bAydGhNjttiqtd7tyqMUl9kQ3mpLyB5OReo60h
aq9um6uR2mni9j8/Pj4R7la6Idb1rLpPwyVnD60v56mysilhXRX6zCZJ7fDPRDK0
5RV2RFTYRQTE0OzuIkvRYmJHdLU29lTaO2eosDo2kMgiEoholHEDutLFWiHdBZfd
R1U7u29CyF/LrY3zEnIFgVvLCHKimeYX2UdBIUjjXisXxqA/lc5Rgud4iqgc6Tek
RME2IEan1p8bCt6pvvK8cwin9CEuZtDGRs3OSoJy1tD3t0e2mkvDbg4L/xE/Elzd
2PINahhHwaM8D1DVK+b1ZRltgy5h8y4TQXk20XrxhQ+DdRsHhx6dR8hNH81IDdbe
6pEbhAetPIQOF1lEp+UKkVhuGwIOM8uG2Hoi1CoxW0tfPFlODG1OVEg0clR8j1iu
SS2da2Ih+FISvkUZeRQc423LXzcuPshNAu8k+Iub2j1Qf78HRo+718AXhG+BXH9F
crdetcTHcn93TdS3/ZMLKjD0Try6/nwsOArlo15ZVOpsu2FNk+u2ScPXJojqsqtA
1Z6n4MpQ/GSvCluzZueqj8HYCymyzUHTY52uz4X8gqWR54xCyRyDta6iTvKpKnEV
pFQsu/3Or1Fu+AeyP4yp3LizUG8bGly1k3TCpBzfOvH9jKv+sEeAZvmxC5SZ/NKL
4xgqHNvp5nhKxscZyQPh41hogvnPev526TFob0txvNXeQS975MkaC0DZlNweB0Rx
yQex2LSf7T+cS90ECImSWoxRDFR21PhEaUJyG+MEhhLdVauRtmzuGedxuyVPBmXJ
tS7s6HHFzDasiwJsVhcC6DTWqtyzg6JbYmJatqwt1ArhPs7/KPVI1kX8YDK/77uT
IDNcWDPGPPhLeAu05xmgDaarztKwmPuBLcWYX4IAfumW3eIzDge+vdSyoOZOk5WQ
NrEJuosh647dEiCSBCCZkYCDEJBVgwMYD7iyyejdRx+MbCuupyKgM+nVreYWYrMS
sKY6M3xcCGTbza17PzT547IAS8oY/WJoEeuecgfpRE60IwA1PFLYnvaZsC1mGDs9
crMQ77ijVgfBlaju6JNCeusNbaqRnq4zfnMYlfJdi8+poWkr5ziRWi1wrR4AjhVH
IujVZ6dzevMuBFrMjWQz6a9fzAGeTvf4Z5MrqbO7ZJ/L/A98p3+/n7hY6nWqNpRh
GzliEF+Eijpg+VQWfPP1VlA3dEwLilziur531eUh4YTza5w1YSaxIdmiYaDWoF/z
asHl7I1iMejfjVsz24+YN8feMaGdBDrbY4agtASmXQJnxOkkHS8QhDxzeyeWuqhB
2dnqS3euaShpaXBTciOyJVrRaA6GR45oebFM0n87QAYRkQcA6qL33Z5ReoMQ/jEt
TH9OyxHr6sdIQmfFLqqa5iA0ZABEFeMVBY62/48WQxjmKfQuch7fIgzA4rBp8BbV
RdUAqGszm6kk4YvCy3kC4r9EfO8AnCsDn7e6SUxdGi2DsU93xyrTBlIGBRA1nulT
H0FnqFHfxcwckisjYOuRI4myxOQBrFd6z8qg2nVNyattp9qRTFQ8Nr7kjP89ADu1
IRI9SgNGcRTWu+BSZN3pbbmbvwsPWrtYQFXs25P7+8ULRnIl8W+Vyr9PBsH7E/Hv
D6iV2h9HSmkKF8dAZ+29NuBSdjZGlILDBYa0/EySICTJRgcNkxFeZ4I0byJZRN/9
OJgdXyfNPpyC0O7Yw+CK1OK4O0P1WfHVKzwPWFJFs8FZPE5XO6tFmRDUb5VHZS2u
jTNNIOUyKab0p2GHV4D3xnqekysFXHMchtbFR4CjdqaBqIiWaoK/3ULvAQenHtGa
oCjz1LlU9oOjqP0x4BTSCz7K1obYHBsrIbmQ2yi++nNd2yJvhucg30xMJte+UVVv
22RcDM+uvjl8NzbmQ3dh4+9z3TR/2bXDuFf+V6FQ4E/g5JN/z2zcQHp+HWkHh/Pv
lBcFdJWaOewdPtpJc70ET2qMyWOrbzlhi6oZ0w6dWvZVn8g8IPBxVxEVrsK/EUDk
bKNpWLgj0T5e0DtaEC4chVXtYYyotl4I7/8OjTd41qW1om3mnwx5RLB9iJRv3twv
DuI7KahbnnTwVrkptQcrTHyylRHQzQXa8xSRLQaCUfQ83Bs2ZFHXEO5nV9+fs96K
mTZRQXpMhWMAD1zA9dXE/HznI2Td+cBgnXknZZi3aCWZdaQeFQMSzZ3iX0RWjLLY
rJLpEvPYHm9xP7PFl4IPRO/C9U2LPuWsGpdBKbndcY9BIAMA0zxAJ5Ni+7A1ltbm
1c6SViXnYR+/so7D8U2cbdG+3NpdudctGejbM2GOHM1jonJ8fsD4HFtGOQ8zqDnd
wo2kAKDmkFbEOM+eQetNptmVnUZilhvctVPdxmwKJaPRqoDrCwI6xEL30r4ZlWfO
ta2q8cFMwfw65TOTvjjgXTskohgEnaHvNepSILh4dJ9G/47kQC6N21xgQ0yztr0u
Gs3FIMZXAo3EzGgsI2kh1jwKaXKH1EPfCmXkGIObjmrbt9e1BYOI4XI1U3nX/I0S
2GPLvuiP/2f0kz0F76pbulAL+t/qwBrQLUqVywldZDdtCc5OLoUl2IFLd43wKR+k
2cSOZdcxs4tHkXNEz0U1J9yVNHG4rJOX8vgcoGV/AgOr0dIktisp9/T1UkuHddOZ
ZNUN3a6YjbnfaW/Llo9yWAgok+wBYtKsoypxwjt8xCc6uRbty8wVVJeEDFaH3x93
mMZFPnAaqjD24CS3/hCaOXFr0f8XhlR4woW3npGZwLHJEON9iOCZ5Dh6KA1DhyAc
WIh07I17GOX5A5cfi7Pu0K6CONaf5KZxKsZqB5gYK74eU+FgA0ybnMH3QWBZY7Qh
bg8lP/Ndaqc6ke3824Kwj9b5a90CBxmhTQREUnwynpO6sGgz/RbUhRSW+cH7+iza
9RycC3FVVBKkw+L4A4ihW2QbsnGR+LBcpyyJTwIqwf24trScEMRKRUIDEfXKtQXP
aLH+UnTM4/tIk7bX0mYzIosurexBXu5VJLB9tO+ZmBd0xvbapLhaT5L/zR5LO5we
1FY4vTiHobeTSom12kVJ72h0XkmymlnCUV4VyeIewRDI4VgeeGxXmhKOtJbcECl9
MM/GcOazemu97Vmrpd3EQLw4MN84wBhcrjxxrJBFNFGXSAKFEqmCrbd0AopO/klF
W9HMjvV0gja3d4QnxRHiyA270e83tnPVDEQMsIK0mHqHlaQFHw3O/GHNA6a6Odjn
gUfdxISoHvvbyoBuWKW/pqVC4VK/tnNnqxgjDRb97uhK7mfJDLebExPPpR3ikSzr
ND6XeEMkcOeNFgBdbQLPsp9ZEfkUsjjBiNybh/9b63ukRMpUHUMeAjiQTn4UDXtW
887LtVh6KnxgdD+adO/9ALvzz96VduVXO4glugIAQGfu+ZzTGkd5EzeDBrxIlo/n
k2HKMsjX4I2l8cwPI0DP/P7kCs+WY4B0ZH35c7CN+xw6pWYAJjzsfnc7WAZeIOLE
rjh6Rh+1gbwhNgENQtUi6gKV8+JbdZrkZ+VSYKCik5gAhT5vu6u4khzN9J6GTFCk
/EhemedjY6XbNXzEI16vCXXCcuJB8Bs3gxcvfR0f4eZZ/1I3S4F6bbZ77rd1yRAQ
zg6uxFCa7AIGyhHVsnaUFjzOj0OROzUUTWvIf3Fnt9IzNB2aVpJfM24eICxnpK9v
9G0c5YntTQNdTSufkAGtarppZ/qLoGKk8EqtchiIDqYYK2nowiIyB2sA7s9Xps+7
N/dym6MM4W8Wfrr7aqSLODwkILSeDuFfR7yZ18KVA9GNHw3EBV96hLvSq1d9uSgP
6Vmd97nJE+xhBSimvdhhWh6RA/qthyUPlme530Un9cqNR6mDflRnJ5jP559y2Hir
oCo0B4smpNBGdZ6JLeXCXXGnHwr8iQ0qs/I8lxIBZSy2aVDIjpZSC/uoz4h0IUcH
uF4WI+E2XctB+bqQmbsPl5U2eOOaGqbHOWp5vTTMs/D+kkrgS/kmz74OFziVcpnp
E4fhj0MQZouPQNRGCTNLaEiPBitBjTs1u+kxFCY/CMM8PqRuJYFbmqKp2jpU/7RT
06ehMELmGYU3Ne/2H+Ernnb8hgHQr2N9SFc4bVP4kVedkTKPmv8GTBZrGmZS4jGa
UtxG3gxTaESEChABWRTMI1ltq+ksRA4gmRtfnI/wOdgRmCzP1YfQSl9YvzINI4FN
GIluLKByYG1y6E7Jz74cBxKZfBAKCE7tyT9ZbsAlDVAcHwpdYPtFTluXSRe3I9AH
MuY7Yyjwgw0cj9MDiDOVSgxk4XELWRwi3UB8nk6uzhOzH1dTg+DdoJ6fqsuXi4E1
M8bXi6BlD+TBYeHSoJYich1nCZWSkt+W8aVfdINSdr+WA/fOylgK/SPfWwi3UF4r
q/PXJI/cw45SzqqR/873eNRHNYXcXeh7tdXzZ8xkxoU4nyAATPQbeF14gEbaK87c
nPVhuFhgyrvgEtkMuV9NPuDiDUcV4VCnF7IlTVjA2cug/jZSdXK/gNgbLLdqIoQz
nyu8LDPDmvGm3041xm3Ui67jHnGFAJdYbO9tyLKJCcXGhVcwB9vmk6iO8wp1tmkM
DeUlMXfFPvpxEQQYBplCkr3dADaMLJW9nLKXwr4fjElNHtb+8k9o7N6x123xXK4N
UjaX6GC+YmDffoWu2gCsjeq9DhsUQgS+mBUy/y/FlqAXb3Fg0EgOodNtiU/LKJjF
ijcq+2/gwioccpbudlhiJeyaEpyRfCKsM7wK91BswgCMfmQ/N+GBuv5Dh5xq+3xw
eDJtlCXfzUIlP7dDYvNisZi3mPuXLOI1OKnoc6v4tdC9LocoLQHek0HRpTp07c44
T6BxaUl3CX8wzgSmZZjLGtvwDfOHBQ+Vlh1BhjBpCTAI2H+OeP1mZ/IxuQg9vwzv
fOzm6jrfvNJkmgM7/O3MeNvjNAn9jx/SRLu9GsZFui3JvyxwjzQw46u1iasunZl/
d3B3JKc7iDiEuOtML7tYUdmvL4WC1FWhPgvCqjmlmX+XMBmTlJX6D1pX5F8AHDxH
XkbNQTbjNUr3jBwGw/RayWaz/axlK/OUidndktKSjNDNy7KQlm9NBfnjAE8oWNr6
ukciaBsxACaDOcUHNBNdm2gBQMo4BR9cy2Rxx6FgbB4z31GTAp176DWxUEHRmJrF
u0bbel2Qa1zuypZka/HUbZhQ8bF+IuP8mH/GQexeYeJeum3J4ESaSeMuWGi7W6V6
HnR/cqV1VLNW5VOe1d5fPPM3ZoH20uN2qSTInxYAHcJZQXKwjiqo5Exrd5sDvwer
CUoJ8fWbDOpIaSmeccHrX1qOalWfwCJmFO/2449USe0fcMO7MzJU1i46VpbXGnFR
lP6ToC4m1hLC+9iiTbpIgOeg9R1Gvx6N1WT8FUS+PBUTzurmTZUP8V8ip40yFvmN
ar/R7YG2QRtK77NJUPW4shYDP1rsaCGAKzDFd5J6hZomVxASIAvanvAunCZM/520
yEoQldXePXIRKmjzNatlezsYzTFqEoZKupIz0tjOWRtSxBnQuIvEKc8FFM6l02aw
Yd1B7Et04ynkPh9pjG+dSRn6vgbVqguHdw6nrkwdbvkWlDelQdFi/OaMDUWx2Hxt
hhwYFnE34gx9vmUmtaEYdxVe5LrwrDTanWzbgtVOvGf3UL70Pq+PBpE6B0/H9N+y
TQnAvkODT/pYVQWt6JvgIFHZ7XE67eTvki2qRczjWVl+2l6lTJFK7qLGkkZbsY9v
nZzEIXurv5b14UG2La4WJtSnApO6g4832kjmrS74tQ6brEdqc/rWgY8Ii6HqGmF/
SAfsJGES/UNncJ0g7T6LzU8KqxbnQTiKIQoVt6vV4ErUPl5veIlup9pnoObrvuqA
5P7MDcyd0/tHpkS4eTNRDlsXVgn2QESUJxBJQ75mjf72QI29do7dLs1HTPQhkcCt
EFy2l/vXAXKsn2OwSJg4AAza00uxMZe5dHVEwjbcW6Pp8GxZ3xfhvng7LKMss41C
vp8T8mzJ4s94BeM7jQWhDwmTY4EFPsCzfz1A2xZAkXota9TusupVtEa0C3QV0CVz
S7vhD1AM7Qz45Ts75cD2MWjFUYFWfwzSWLZwxaYzqZFF+8QZ38TCKExGnLhlQdz/
Rz6oNWp8BN5zdGOukSZFDNEzkTMjpOwc3EZCJC5PBNicM90Vmfed5Es5+FcibyhL
TqWAsegcPP9te5loaO+knMzYE01404JmVugj2FyuiCoL2ezbSqChryzex58hDMZ8
mTOJSrfQ+qyPDrkJZRDV3nQ6tXmPrqh7Ik3XST6gs7zwSuBLt05u27TA9zUeyxpY
hv3yDzNFLOjXmNXrsBE8xyMdiUsbNDD+CI+qg/W/uoLBo3qvS+erSTNtZ+a+patA
i0h+lHlaXLd3CQhY5yEguG0ARWEr++z61NV4asNCctjl42omZGUp+EMVLpSkQaET
Nl5ZCyXSAOuKRQGZSV8GEODNm1rA1gBFp3NXNH9T9J8n1jw/Ru+PWQYQXnq4c1Wm
8CFVLa+6Qi2c0X58NeGPxRtitjkdSZ0htpzSO/dpq1pjYqYBq+5+JY6oIUiBHsEO
dMVY/CZCQli2aX9qi5nJAvWCnqcgpevH/DnNA4ZqPzlxaJU6RjAKyLc3t61eDqx6
nBq5twAmZ2el9SCU7y1EUJhH9bJv08ekiUWm/FzfEmi1egeJfUa4Nr1b+qgWPcfd
LQFXrZ1Eukozr1dCIpnVR0VqPySR0gpWK9kXyvy0GOebWT0LFPnOn+jut81XBXTN
1h99zDPlMMShGd1xFSThSTEdGWTuEmgIMlBi1kH5rS+Q8kGsXtQHOCZL0Pc8k7tg
U1nIcSpyHiac2BnoOXPlpSg7ApuPKhxSfUnDsO5fgwsFdLzlrwy9+1iVXwREI/j/
9uzh9odhU6OHdkmltS+64v1KBN7F3Lq9NGyIg0+2hSZ6/GsOuGDST8VTpCi7jgLT
S13qZx34Rjozd169msXLDEWxK1r/cxBGfUhTgHiMLYtAEIzTPe9opEQt+h8a2GEG
fT9VO/he3tAWK+fwmspzkyf8OrX1GRIFth87Aq/wqIpOpEl6X5ApJXzhBKQBrXHW
uLv94Am2fa4JlDAvr17ARu3PEM/kjK51a6WEHzbRShg/DnzRB5IpzMpWs57bf5Q+
2VfVmbKTOC84kU0WuMzeCJVH2qe/rYaMkGvNO9isDWZayBVGcND9Og3nu/bLU6a6
ZyZbbRcae5OHxsqnUzYEcs9jXNv0qwvijS0TdCgQULfns93yhksWM9HLVBv3Ogbf
vjTwlPYmR5brTkdCv+YuIGJao3s4buv05DJL/uogy5hV2oziNNYbtE1cJr8G5aQ2
+Khw4C5EIH6dKk+ho/ylnqMqpLaREfSspM9GltFbV+WOuVgpX9uDUgZFD7wnfQlY
cPEjp98SdpD30Tf26IgP/rctvCZIqxsThBygpicfkuh2z9JeeAqQF4ZV5A9Qf0n1
Uarfl4nBrTmC4euId4SIpA1obAb2bzrPHrrUBwJ/kPxvNlJtiu+5CCbvcG+Q+PIw
K2laSa599GSwiNh9lcY20ZkfkYgWwDZCvtX7/nVlUHUoBrnTPTggX5PtENyuu1zi
d/0RKtJkaCokv0B59gEaS5qU80CDbrZIIk06UBrBZnwkd9j33pEqREvdshGTJGll
W5n8nOPOu8D72V4yv6EMuvNaBdYqjZfZt6YNOvIM1Q/O/Ue2cNxSCOqzQ0L+xHqw
hmYHKQ7fZYWKNgvEEHYzP36+i9oYRsRY6aNpKbyfDhNZLFLHUfH7kUhgkXmNN46S
IzHnxrGbh6hxpTwzLP1k91KkJ+6LIu+y4uN6FFbESKz+vMBxk02RMFZ7kZGM7sru
xZkw/YnrFPkZ488tCgQ+v9sQsnzCP4OKwe5/K53/YJ9BCKNhoZj1J1WLL6Lox1rs
rPY88/Wv2NXPgLgd0TL/xyesJTZiwS5FfOJbro7yi1U2GhHM+2o2T08GfjvHPOTs
Y+ieFuYFAWoLHH5V8RDU7Fitveub1CV/zbOdpglmlRxNRvDhiMCcWc7MdfeqM93J
AlhMd1B1VqENAjUBYu3+/4GfyruOnR0yMXHNN71yttQ9x3sXu3SJb5YvvEnm9hut
S2n4tE6cyrSBmZxX5YzYmUCLKGLfJZP8zzOeOv3Xe9wykY/RbGft7rR7hnwlnQcs
GfuOOqxvS930aUW5yPXoboVWzk6UIaZLp6uJQs6SCHO2rl+w79LNNYoiD8ROPENv
d+tJzZNaOU8YB5K5pwihiQ2hKWevZMv+AlaLJOY99ESanUKM5bq3WFI5Jp6+Lhix
48e/M49O9GmcYmqpOxVrtX6r5XGJfHyS6qqko3JgbrlG5OypQfOeKGK1fI0Sl0uk
RuETfjMekaCGc/gWnbNP26KA22Sx/5APb4AojIt1YftLPPpr/WKYngxknE+LFliA
DspfJZue4cFNhi3emSUnKwX8mAelyjiD1fZddmnk6mXQfTwGNXSNS59tfaJLA7SG
ZEK5TIrYvgswe/H75kG7kXe3XIouWDMxKz7hypqLG73Y/gDvedF6JsJ3Dhwf3+LC
KJ/CGhqYstIMriEgSEMIr7Dt8cfkTpLv0rTI+8pJ2IdNyziFOQh0GZvdvbWMOVry
g5d7IfZ8TUGfuRUzfQJ3FPU13W1mhu/mzx4de0WUUXc+0esolD0fKdSMEOFm5nJ+
7YSrz7CnFDtKYBO0FCtnN/lHMD/oHCh/nGxII4EM57fpi/oeJOR2As9VkRYZdTdf
8AhudGs3qrx3R0vP8AW+biQRGtZ3mL8weECw2R0PxQ1qN7FMVSW9vIr1aRMxJxCq
hCw0b8B7CBW/Nv5KzpFsGw9GUFS9qJYdJI1FuYJTNTSPNu7rS/lpaeAIj5bIJwNl
J+y1exV4NArrHN0wUUOkSRTsmdLrmjw2pQ2/K8bLeLs9pLHvjNyZpAntl/4t1/i7
xhYTwTYESzwkA3RTZYEdRBAsSAFgDV+Y8+qCw3ctF2PKxbKXlJ3V1lnq4qvh1iSY
25bhh0I9jAduSEYUi/vlByOVTjdqJY0EcItqQdOS/sXBkoIn5I4x7N2VLnKJmjnk
FHhyNiI8QKLkglOIB6JjGrBXJ1iZx+uPFNRZCGJK5qOIaaSy6ULyKcpDKf9WzLxG
gr9vAWGAQDRjXKJTtcyaxm/sbBfwGaVdMZZwtEp1M79peI4TgHaS/90fObjQu8Ws
IrmjipI3+LK7Eq6JMKMbGmgX0abn2ZF5puAViBJl89c+4TkE08zQll2Zp2PDC0AD
cPQoqsJ1Sedo+lQrU5rGABeWYhCv2p20zMbYyl1zJ9GkQQ4vjQxL4srQcL5sePmJ
sgR25Ewb4wfdplsSmbdsrosJ+QXafjLRkkAgvQkEwC3gCCkRmZxpvAgaAg4pmd1l
WaL9M4iNkAVM58fBeH7VAUvN4HoFqz+6HZafGfQGKCaWQnFmiwhuulBA4OWi1dnI
Z6x2ruJdLdJR6CllvcUJ9k9rTnhoWwJTzFlYFQcjvdTz3bTGfsbWWGUUGvn8+Llv
YVhr4FGXlcdDCbFMNJxKLTtCLL9PplK00InIqNPKePL+deE4nN9Dl1xwSXjMYD/9
OY0nCSad9Le0wHQtqFMZSUv2kedI9IGpXPMc7yufxXHizUM76SS4UtgsV46ift/d
fghqjb0iTMj56OvzRoL1k//I1T43Jm4oR71+CynvkumFqUMpusO4xk9LHvFVxc0l
ZliGEY5piSHoR4KXF9jY9yilr860ynxJ8SlBm1K910K/H5AY+hcUGU+5h5Pta3Qc
uYllebT8DYTx5gA8ntdZrJ6pulIuEax0YbW1+s0QDDbjPbh2SmsEnx7OQP6l6VN8
28EEeLNi9P+Pi4/3XiLlDbGa7I7EgqiBaXTf13Mosbd3lDR5v1ccmLVfSxJZW5G/
SUjHCZXNb9Q7dDm+SoCHPDnHipqXVubl3GcK8RQP4sKKFFewSQ/N74+bH5o3bUU/
OS9iUkMKEWS4MbhSPn5Mge3b1Tp+kOq+6GFBJs7wq8/S6suhEPYi7qFA9Seb9ii7
NaHgRdPSJ5vfz2/BNAT5NfyUI2pftkSur1MgoVz1Gwa1mA/syWKNds4hyzGnVzqJ
hIQwkVwNmWR0maguAuvx4IrSL21V2xsdem/bzi6mOL52a0XB0Wh4gQ+cWdjso9sk
ofL3zOWDu96RUeyzgzIXRoC3U6WYEM5U7u/VXp8mkRX6Vu7dMRjU7pu61vOAVHJq
1VgSpp9/LtgPxC8TjnYdzCBKdZCeFk6NOTSidMBeJ6xrpf83ISoR8/8a8aXQbdbt
5LNDQ44/VUXRQK7lmwxKxVwfKItKjefb76ko30zBujr7k1Qu9cAzkK+cktVPImGr
DpKgXNFkq3/x97yz1+F9W2gBzpvJieVstiwbJPk7ZNOXXmjd6cEZvW29qYvYxW8x
pL2gXaJDxC0imIKI6huFOW4d7TAKo9tXVXREUoe1Jr0kHs2YrRKS2srLpA2Blgfv
VDdbaTfdVX4iMaAactQW+hY4kg52WIzYVC1n9vp9ORqtgZ9UGRA405lW8WsOq2mt
WLwi0j1XjeSwEvY4IYbcAhSgWDnogbBU4tGAe9U2nR2zt4qNoeU294DamLZG7tA0
WJddCjoqJtLeCLH6//57EvvrfedTwPOG/YTo8f8xKWBWKzjaWoAW7F2IK4Dka71G
knyAtXoZi6Co/chuFr65KYT6Yvdm5Ih0Dg1knw5BE/O/YTc/zdf8VMI4RysNFvfz
1ns5l6VP/21ncPg2KRI9DAPGoWUalnKpojzaZ5IhAeod6a7dZXJBmR6rVIUzR/8I
vdc99tUucrKKKF9XU7fE5Ah8h+deVXxWUy+q7b0CZmV7J/VjyC7XyTaMcVlvGaYo
RTk1kjnbZmiGvwkrYuOlQNNnFGSYpDaaAxvsTRsOPSE3iHjfk3jekjZTx9R7eIQj
ycyTnQxXfU00FQHlyIlj6vPv9lgg7fBDOjzSdYkSJKuhY+ykrxY+rAM9hOaNcp0h
NZcy+lh4rNvnCSsCBAQ9qKaFXE2VaNphGy1X40urtbKT7XDVOOHQjl1iKdiQysG2
kfGoNl8RYSJs0ePVoDXSGRL2ghtRubUFowbtAjRtOdX9AEEQfoY6ysFzbVg9raOh
oyACcpKRwNDqVVDbgpxn/LemFH2SZCN085th6oPr/ZItzg3mwPksAreAGABjtxnr
m1xOKxs2VtBVhJS+aY6cUSVmlbulkAHsAluqnQwIUMU2wSr3Rfo1O9AFppqJk4Go
Qg+/57ujUXqeMsIZFTN0tIyBDlaATEKXmuNLfCFNqFy2laGuej9CvcEDf/1izFAk
K2i7qk6Csk9jwrRuPEhoTtZv6lx/10Es+8fRSA2suzuD1Rrp0eFTjbgMWoxGYR77
LyEBwvZi5Sqj5JqdSFJq2CxyR1+Sfm6AwdS+qweK5Hh3y7yZX2+1lxv+AShPPpFJ
JKYtgyGH0m1rBcFn9R+AOZqPqB/tjI3p2z2BzpuYDShevH+Dl2yKl3ucA+RAVjaX
XUCh6VXUo1BfEL/DXVZtle0Mh5CE5Qn0Qi4haiNaOZMHAoC8l1pTDcZisZYJCmB5
gV/YIinaQWdfLqWIHDTvIAh9VOJ+g1UAVh39YoSngIt7In43ilfLEU2W+hDbjxTj
7WJJ7XFicsuMIdVRfIeAElD5JTIrDsvy+ATZ1vRJeN76sgdhbk0odVCy09V9TKAV
UhnF5MqVX61HRi2Q0AeWjadc97OcVyUwRZxzQspMhJQlkcM7NOzCtiTv1Bwf+4+N
otchiFGgQL7JrnDiFOiS6BlRKOY7NhhtxXMVKmn2dk7pkDmy5sFuCdQbu/cdKnlv
WeOhkc2nRnfxVEcyhppxcpWtT5clzS2PP2ulJi1Lv2fo52gdd/n3gv1pz9tDGV20
88bY8RHr7TILpdnPZJHVv9+jU+IDG8KVQ3e23VYCzTuCWGLSToYXNluH55BLvEek
909YNwNi8jVpTbhAtBo5TXAsKoRHZsyKALTSOvxm7Yifta5rlXOQYOPrtLgUj/sq
ifAWtRVqfUfaY1jkWIJHq4I6T86R42xZfbIWoNtr1Qy1uAoByAxjeQDKA+HjA/bO
IdTqYk3yN4SP1snRUUfPuHkjC58YXwZupZBG676wLaqPvQa/43M6IvwrBu2hM0lB
38fjhu2+Hg2ARVzbqIihJbTVzMqYYUMpQocAZNktPLsRvEFDVKjeJKfnDT/dCAiK
npM0CwHU5gT+0811wG6cpZ2rGBuyaMxF3WTRD+phBI8he8kV3hQwsCBPbNkpU5ye
5G3MHE7odys3RQY82nuDehXR8cTAEGDpKsFwyKQxVvAyG+uapbbHfrz7jeXfexDw
WZAJudp/589eBTKtmzo9gWgUmaZPe540ya597qLGu4JZwdwNWCSnEf9RqKhiBoWn
0fKksLXKxrHq9HGRzIgXpIY/CWqWsVtw+IORfkSDEbLjP/QhaBvYlONsjlNW3V1U
FI2rurUkwfphffsuHLlHhPoDN0WmcVOCmvHIkJubp095G+8qdD0AE6SdfiIfzzzq
C0SToak5lmiPAlrHy1VWBj3fxy8jlqXCz+4yp5R4AXrIetsYj0yYnkg+aTxp5Nj5
KeUv/5K/8CA5dQY6gA4NBgno2mAW4lBqOp+WjXVPxnB1F21bB+GFUEUXIDgh4yV/
M+grquvUub+zxmDFNaFcc/QykuOpBIJlR2y1xjhVHT+XKDNJVFi83NfrCLcINn9d
8b6hdx2Of/O+oE+Yn9qFJrcmw6zfgxveQqyYUBIGidwdkVbFHiNTI0vaBQfWJs3g
/vgj986q13+kjBXDQYaxEekwrU+pi4Nb5E3OO5754eblRuY2kDkTKJ80sNpUDOqr
ykrzCMeqvPaIL9am6ki2e5LDMC1bOyomlTuh3ZoZsNYKWmW8Xtz3JZyaO/hREqRR
82806YO+xTYFZekZHTxf1vIj1kpB8v8ga+GxvqNb6yiuUNDaLonrdH23mSbHHuem
PS3EyUq/f4V6PX5RsWzg+NtZIrKT3J1X3+VmtuHOMQXmdyFtiBmu/QKWVVrr8toG
ca8EZiavu10UfIMN4hTbvQBy0KW7oix8BElX2xzcFgN0YR7Zs5CovrKR8XS61+Il
kQCoXtcZ9ekTesZtUmgzilkD/OVfsJ9IlgiObbdiMfjiKorliEaqWqcHgVBiuY0q
SMXEGWMFETUuNkskRUFC964Bi/G6EZ0iasvCnWuwpa6F8VjzTS95CGfvO9Pfykd1
OuvoBtLJWnuOnTWIv5a2AuykanEQUYCmnaNMQDg+a9eyOm4/2jqaul0OU6INga47
nq+quEd3C70Ejp04CdkRU8cfQN+kl8DP2Y1jaj6Punk82pBRqEqNltvUyzJOagcH
xShxaBowDzj2R+KdnQIDpKnxfccg9Ldkkb1rj5OacCubg9R+WEPGVwvXWVqab8Tc
XXujCMw0U8B2tfLKWyvvK8aww3/nhn4awL4s5FozP6BdYD1yiPQinRRXEksxbGZZ
Nve0zEiqMqHFlsHTZMa8Wx1dL1EtK4/Zq5NpQ7TkzKpn9MgoikrDOWiQpu5J7rnq
CfFhZgeg1BEE4GYjbNXOlCjqNqqIj8Mx1NzEzzu6qe9thvZFHhG19BJe8c3Ihq0s
PL2z6Dkzic9x0/k2aJoRY4mRAeLrISTSJPV23nvjJF1T3dKbKrvKjb161we1nOE9
fbTH4MOT3QydmZIZWLzvx//kc/SNYy1oMp9sruasEzNdSeZcuI26Zi6kQugme37O
v0sqQdCtt/vwW7YEQalZmu1/wyPk5v0R8x6qPESkgtNJndrK+8es0vhEqF/5zM1P
EjCpIWHdQ9v3FFvf25Ct0cCddOzTAx5Xn/bIDD/6HwJpbPuvpUChZNCRiAqsjPx8
iRFVV/sjfcz+1pCVAYFrUiEhQb7LRNrG2e/uxPopSM8Mw6XF8Bv+xvgF9jjIrN5c
4cmvEQD7tX3inLT9WPNzm0K3TgJsTQDPEk7i91z9+0qSj5iClHm0+JXur2ptPYu3
WAK0ow81iH+yVaZdWNfgcejaqyMziWMa1W9OGSQyLJdcqqOOLFQecF5n2A0wCevl
IwUcQt/NQlFNH4wBKbLJxzEHEY2uoR6wJnu1SNg5r9gOJlWHybLU/E5fOrLnSY6X
WFvbeDQRg/3L3dVd/k9kb+OME38LRtIoX1D9voJbE1Q+qKufkboHrh623od1dqW7
gpvntXNQ3I4M00blNRF8AvzClX18hEuMjyquzcFM4rbF8/fyWnQUZ077rjQKKW+H
7wHmbSgUUk9xShK2ohWRHYSHvyaqCigfezwwGjR4A78OaX36gJE3QTOhe3Ldl3yt
y4Bah2Xwak4/uaDOd2+7LUqI00zEuR13M63B0UVZHD2TCNPEqcg2PariuE4tQL4h
PuYhhwuVylz92GXyytovzPMmHAkhKCEjmPekwUcxAIz9za7HTi9LT1K3QiZwsDvN
WEp8+cQlfrORJmcuhFY6YmZon5SUxX5jvuDAAn/FJsRAu/3e0EHr/rPxB4a6+6uL
GRagbPUoUzskEHwF9T7FbqZZSvFtfdClMqfCHtjBrstCPcgsbz8j03Umwc2mWRRD
AVGcDvV5LVvLaCahJnwBbbgz/EtAyKij1m5itR00zdJRR0nvZtyBoFNhnk1d9/Ko
7AUTbHeSyFNllcF9MxFddtoH2EhuQ3ryjY3putgFNG0kWPBVHH9x5F2ihV+XcMi4
roncJc0KNSfwKUpBLfGoSPlshWCL25cTUbJAWroaQcmZwlMnJ373PBEg9B1T6qSI
zNAw8Uu2cyM7SBT0hTcpaigZpNhVBWaeHV+zybtDM4WWle8XDQAtdNfKTt7Ay5L6
Ty66NRvVE1dAttnQRIkY4KME+hyj+5pcEOW5s4/lcOJyHQ+/PIw81bAnKw1+fdPl
PCvPMgZx5E4sOuqncZAV4P6QBUXzz0iLpLKvAGmAvmJG75NjsMSycnto2/+S2h4O
msmhyJI3u8gqCMEu8lr02dx3atVT35LQCuyBcDCCMJcAlSC9/eW+ulgcfh8ojL+J
U4KZkt1/9NOwRfwQyp0HZnFF/1Za8Y3/rBrdwM+prCHl/z+wr8JA70ZGms3PWE+8
19XU91/HRPQOKfIJk0LdtzEBLdpFnDF4X3Ym8+f92Tkq7RmCll03TmehUYdJukD/
zjcuMUniPgpsK963rHmRp11y21iL7jq3U5uDK/BLTXJX8Ix105sLXuoUAwlV8JU3
/qUzytUZrRWH67ahJt3Hz7A0meLCcjpvEm0Sve5YgCPMsu7ZJOfKGKw/499d9Iz9
qWHrwMirS6rkSaJEygi00kCJ4EOZyFcZwQdQZyeTmyltFTnr0WH4j0uCM2dOS8n3
zI+DDDzkyehc8H3W3/EMLAXSKyGjahnp4Im4iNl0s7nTILp5DStyxalWPBewWrvH
Gc1tKy7KA2K9y4qfeAB47WOpVRW4KwBjnGBR1/iylfnNgx2zEjJk0Rkz2A355dtg
0/yjOaJKdUG3dDq8ynSjM9z786EOYWBPNP63fmfCkChR72Kakil2k9heKYYA1z/U
/25PpGVdqpK4KDwaDrcthTAQMiZar1j7oQKi/54vQrsrZ2xIjUTQKrAT5fim8GSP
mCS3apzzERB4diQdgRplIHY7kDhELShE35QmKkjXbFqU7QA/TKn9Vm12JejxTplS
zLBfrUv3M+3qoZZDBzCOXojp855s6EHizWtsq91P3qDCMK5oDXfPS4mlHB8V6Akc
ZUvAt4QOH+Ffqag/+/POY0i5M4xtnnLJZiEbr3+8i5UM9cuTv7qd1u8uKEHb0BXl
/e1IiknyWV4xSuLXsvi0pz4k/Q/dM5AwxXe+ljxJ5bjBeLIdT8SJ4mqbbeEqOtZf
9vHNvhBLXfkjjpJli4+imu6zzzhloEShf8t2J8DZ0b5aNVJoQHIxvEMa77iTfKAE
DjOQ7l6LdCCvpBhnjQxILDdR4s1xgw5MAEKAUOsaZWhXsNXHoVE2UN/Bfa+DioiN
wuXlbz49OkjA/qO/JAwfaLlc2Xk6yyFAKiMmty/HDlhklt3dewOJrT3VoNZtLJui
G/vb9Elk6MHhaS5+Mgciux6P+Nt3fKQ3TN+J445J7vMqA+/InlePGKgFfp6jay6i
ZvgfuHt2exygmdnh1Ex2VMLsMKKWJbivl6pBHXEx90Olcyawj+sDW7CV8oO3g+pQ
pUxFM2oBi/3I1QUNssjOyBI9yLeFIV4iTgC5CpDmLrSb55WZV9T9AzASFRLXiOvy
AUDqb9xbwN8NyH5iOGzn3rHcXw/q0bmnUQxdq8iu1OchDE/QevMAtmo1MwCZHfdz
6ynxSnxwSf3s3lOOFykOzHCwYURaia7INF8qQ8NbTeRlMmSJs9gcjV5z0OKN+EZF
FA56NKYm02TY9RTVYmZnEQ2JVbCoY7/4BD1IBLvXymn1d8JAEYWVyugY/JR3UMjo
X2WHzVWlJyd6Q9pNYCof3Dsxum/WnejooI8+MPkkgCDfPfTWZhzwB4jtP/0JHtkH
+KK+kz04G5vDECFr+8BL5qZoTozt2GFSn++tNZz9oeRib0qdoe93SDbdeiqIwI/P
lVuqh0p6EM2vXsb21hNImVRBqLYAHE/ZU05RgVm8cva5//qYbVZA57boQt7VadDT
9Okj7o9YHUxFtK23h3et6XMDx2707NzqbVDgXbuCimvG/wFhNrFB/g6IujPVhxyB
r70f/zdOrz81xAERNbA7Ze+O11kGnfl4d8bnUHArqRi7NvtznonO+8ry5xbqKpb9
LWulQx0qlESEowtd9LlySFKe0EHFOtPu7svugPm5+l0G4RY4k01wFtxVihSBU8LZ
kKJTPEAGPV0KOT5Miq/wvEJBFggYBaWCTxm16ZLyfItIISTtCyESZqpjLtxGDVD3
l1iuMX/8WS8wZLa+AYXll7PM4X29g09G2TqGveBuaJnPrbPCEfRxyRp8cXEXjJBA
CqMm8k3EH0tvnsJ9oAxvXzKnDMLDSiBM2P55WFAom/XnQui6h/elBymgABgmAMbZ
GBvXIaOG27iWVAVPZB9e6ZeLvSBCXO7YydPlohL/SgXI5CkHDkwXEot81hIjAZZO
/zscAVij+201GMSLHHg3Z74/3VkpTfIirk1bnwN4d9R1kkaNjUL6RFXdGb/rizTM
43HVLOMq7PeNTSjoit5O2dXIzyKK562riGFSBNacpDszMoXczdDVDQmxobSllIOF
DDrB+Q6CgxhHuKdj/fhBlp9JrUVm8PYvzcnoUmG3tnXF8ANYXppFUxEnwPLKTzCG
Kkz6Bc/aruwDi/W3X4Xu8OM4E9ZBB5CNuN4chzkJRX+BzcgiwiWwCCVMAyTC5xTi
GjFK+FQiT+qlGOJMZbEX0s7xvOddkSvev0xkyO/klDdfrcBf5G4G4KFZOqPLRseu
4+TRSU7Gyyqx26ZNRd52OY9WRj8FV9F7WVF5qsB+M1F/Redrw88B6zqZRLIqlTCc
2OsO9oBiKYHk7uyFLpwA0rtbvDk+Qro8ncywjnBmCNaiWrhlNTxiSE8p/iCryxFw
pSPg7gbbnldpApjGdatOUxKhkkJ8YrKvdXMv2KCR9CVE91LL+TsZ6uyoK2A0IEBp
zPbWfmucunj+ZGzqeK5PEKaieS8VJPP3cq/8I2WC9NBmtuvTgJHlbJXagvnLPLgU
rsWw3FvarmGqS172le79qOnQ9pL48EhDX6tHUyo3nGkhpjPRolWGSrzRmZ+VVkG/
OT2ZY9UrgNIgTHj46orM38nBJHC8WHV2Fl0zB+m1fo7RxMWmvTEcURNRK1xCp+mQ
uSZztM51n8d7/VN+z7zVE1rThwY1mXJbDmMzuBNMUXwWXhaif0KnLgcVgFo1etlm
8Sk/Ne5ItL0gKvKu+vSO9PpPdrtys4Au+W1ta1lF5chLs4KtIS4NzdSiGVqQaLS3
r9DUUlQdUzhAPR/NqZ+e2ttnZda8CSMEN8H4L9NY7rNRkr7uZWh2BjolgmMifE3y
xkb8Dzg4/0ZTXB6gfYZDtG3MQ79iNuxKu6cqqSQEGQuXHwGSlnTPP7lmqjdCEFS2
K/lGQIpdceyRliBfAuRlMoCIZxF0dSLJUgdij49hSc/ANw9j1K/SjXi6LNQsOgBS
5Pljhq9dyhqKoSmg1Py6tOYAGHJjvy+Y0DUBH7W3lSIjh5xb4OvNApuistTozEHv
9fcMN6YVU9MkDfNVJY2b+FWbXSeG/EoxF9r9sSUS6U6PhA47HhyrEBMl1NMZx8RV
l2bJ1a+f/7mqBbSCmKwTHatxje/6kRQkTu5OIJOaOcxjDK5R7Itf87y433nLZ4JW
3bjjncJz8Al2TAuLm35mja/5G2Pk8EuUgocW9nta1OJgDtZv/iY2AMudfeLFfJqn
tfTmg6nZ+BKV0uGod0HfjUMCHyta9jVQfI133qfEQNoDo6AMBJcPSEtyV6xp8pcV
ZZZbN/Wkrjgo8ft75/TEi58vP/grGz9Q3WprGDvoqp67UaqFlCv4hyyVkRGB/R7q
rfPeVVHHwp6OGK0nEv1Um5x6S2Px2JabUyfqq99bZwGwM1yoTdiWcoCTKT0n6q04
3f1rxh9vzD7+Ima5lvZWEKKf9y3vRFQtNgbR3CR7Wgp0BgJVMM7JDMicVK4NAhdM
pQgG9/iw+Nw93yhInFMNStTmaSmOSpCABe0tkwCeQ9BwPMJHM7fluStwKVAC0L9Z
RTHpt4icxZiEIgpIGFzmJpPg2VmebJu3nRN1l/1yFHo/foXe8rJtkV3+P/fAsAYS
lQEmcEaO5ahUkYeuGGPqIucKgLW/ZLjaVvAGmuUszbRh2o4y+hR22Vj6PSmlSLzW
PNShNBVKDmPkHOjCUZ4mkKMlQTBvxnbvx8EM5kMoWsORrHnQ+SMaPSy+TQ9tzVgw
pojkgMImpoYL3+x8tsFZFYvZYxNbx5+jRetYXWwFFr/mKbz15c6420PvY5LOCsrL
pEyvEGS4kCwMY0rFDDLb4OFzC5xaClhrd4CxEl0SpGC40Jo51Bh7HH/HZKx2mg1E
91WDQnn73SysXdiWnyRaudVbp3Hvl4VHTvKqTeWvcWDkIyj1Ruy/Df1r48whrGgB
xDVlTJAo4LDBc2LrEgyPvhmB/ApmeiYu4ChhntSDj89COYMMIdtxZWPxi51cyats
3HVfbfA/jVPZgzb/KPS+cDmkwRBCvkFIFTTM45XOunKsLRgxh8X2lPkH8glCHtvy
3LzEJG6grr7Z5FfRZ1yQnlg94YXY4ojVNPFOM/cEQ5uVN6i65LnK6qfaFGwoua2C
4Fs+LhuCigaT3088nzQdsh8UQ7RkERFhGK8tuNRL2kqzNPIqCT+DItt37a+Qqmco
aadBohMcVYrdIgz9SR5+JnovhuQ5LPn3qDmOrkN/0JscrDmrbQmqgrT2aoAejLj4
l4d9hmfeQLjMKEiBJUvVfMwK5khyvUYpLIxRe7nruZ1PKGgdySPF0Masq6grbPMY
BsYdOFw4hoSMW2Jq1SUFJXUA6Ya5WtOJ6HvRibBAReOCHfvEQ/Xn0QWN8bUPV8qE
xg9FA2iLz3pLGSkyx91wqZrSWIFyomfFtnPKAwwdHp8y17k49nQerfDKNLDpJA4o
dzfId781mzL2IHc/2GM5WOii7StbnawZds8W2Rk8BQsnRI/s/ErkhhXIt9sIIQJn
+fntk0CteAEsUYa2FohLsqNY06u2isTZAzdDSgmGKnwFtrx9gKBjyBsnA4MWjZQc
k/n0OEiO+sTqSGHka44I9P0gsCNfyZ5gfg3QdpW6opxUh0mTAYVRuUdDy/XrLE3H
MBfbXqWMoi3mPcjZeX3zWvLwnUZMGL++APxpKvIcL3uiGN3hu94dDsC/blayirVw
GFIuno6WTv8opjBaNAFpDHzaaRhtxMLny5L/aOXgG3AV77Lz9eZ/qwnGvU9NNt/0
Sn7QxZ673G5FH+ejBwpE1TtqwKKtQF3F27eKZ9kdNTdVl5/hsf1phwDDCspBHHSM
a14To48PKCYuy6wbJ9bHzpJuPp8qFCtlSHYxPybLBQwjnWuXvRyDMXNgkV39F4/s
35yicVaGsUO9eAm/LKVSCZURxlpFo71J2yUGbT6i3fW0TIaed1WM43I7jPl5YqNa
+8bWKcMUMLVw6x0TYFkyR94igkbsdgn5rljPkbcCbGlqxkEZoymd9qauZEwF9UIL
/ltxBt62kmPkS1kbKYRq4InMZCyTEpShtbHfSVFU5xNMn/Sy5FMJlA2GnXjOA2lW
V4x4Zt3VCv8PeUhbLe96VdnJpMXKpu7gAbUDz6wiwa0Le7dsmSx7FwY/9loxhMUA
LLMiDvkNhktTiQP3y8Tf9jzQup0gyOt906u8PNNjFaP4T7W17+VJuOtl1OG0HzkY
uVpVzKt3dPsoU/XM3LmRc5S/ktkPqywLWJ7ihcLmmF2//5OCL5DcGfHillCZuKnN
S8kBbB4NKYVxDkDT572CHCe4EzRnl6mbotDGID3RaiM+0uw3iRIvaK4aS7892PAc
OiiFtYD9btU5tiPjzZ/hbBQf/OlX9LCNF+igJk2j+8sVUjDJNmuhVPtkntAwYsP5
0OssYoNn42fKXFGLECdXyWfWhsk0SZBBY58viccvl2BppnK4Vc3NVJAcuulTlYw0
ATfsDSckr/v9bnOIPfKftfGy9D6AQfGL4OT4uy5w80djNpk/1chXr17m5exK0kum
RDpXk2rFSdc2t73fOXh267Qz1N507NO53yHs76KyTRpZZpuS/Eq1lT/oJJota+dl
QqHNTY5iP9mSvXWa1nhmmhLPnxagYGadeOGupB9+uu2rMroQbFxJZh3l/FQ6yh2D
DbbvIONksyGCY5GoQ5BPiLS0l1kxMPTC9XkkEH8Qg1yQe2Kzu+uQwqT1zB7zzGBF
c3nn2joI1UZlGFtMUjW9hV30uaFQGcKxf1mOwvZwhFHFzzBv6DPzh8i/Sh1RJg78
p6bBf+oLomQzFWazS5XQU7d6aT//tLUSNKClbZH2Eo6hkPi1JA1qEcO40Rvl5JW1
Xu4MCLmzadUT6Hj/KJMEKJYQJTDploF268BWUz/fLbE7W5H1D6awr/rRTl5e8FpZ
0yNjKuV4ZhIFhUgI8CMMsk0c2GpdNA8QdFwUzLwL0jE9kcJAk9TqSxiVZPCi0qNl
WTw9sHcPUTBwMym7ZH1TWqCmg7ITBM/dFTcxVrDKQ9rmJhGwfv5cjpiRX9VuVhL1
Jh/Ocx4skbJcXNlHMMQ/vIIFwlMkhxxGVhLGaeUPRNB8I6J6zKGQN90k0KcTcvhh
rgqvRCJb573GF1od0l1jQZ2ueIqEZvI+LgsPmlh9Hw3HsHZjRyXeC2GCVQIsPsHT
z7f81/Nj+MaL9xPUj4drvruJiHbyq5CwYwxTD/pOKnvhUJfFlFc/d5nyeNWNd9RS
O4LI+c1ySNWwgIzGcOjzAtbbQ/T3LK1+/pG9GEzaLTGHiTvGvtdwFSx6HpUrPd+w
ouCLosrf6yMl4uA8ZRYUZxVaIboZWYyb+ghPBsvNZZQA3o3hJsz4wX/L5RZ3HrTC
S92bx37QiPIK5ADxQHaXqondmD/JHeMo5SVLjGdq12m3S60sU3cdA1yjTOaxf6DK
f0QnSDVLLb3ZPkq8dnwqnfocUhGuc+QvScJOX9h3lJHPJVDRy9tEX6cXdC+VYM+B
iU5Qrj9LXvv5Lcha+yOPumX0w9Mh4BiTQ6YnrF3IXmQyS2nJPQ76zT5a8tMQNmj8
CiPrgPuFt+5ci/yUAf4e3fqegyHhnFqE2gr9mV3/PamcARis985wUykNafArhQYj
EqCY4y1YxcG3uheUGd3QCPH5cbTHsLDegY4Aj4D2moJ2BtJZ+YrmFT/2dWPBBGkR
/rsN7T4SJZ75bCOQSYp7vd6kiOwSOtw7rPgzd4K3sEOGSjyGYCPkE1GCUDZV9Btm
Gpd1RNmipvY+2fL9UWzDnU4d6gxOn7MIYKc2MZpL3YJN01gt04bxQtXTRoFMHjlu
GyP6VuJrgvTEXUMtumfuHnWh1q82DsKmn6fp69Ip4RPoeVy86bZz9jK3ohQEKmqL
6BAmc+0CIMBOwHjM6XWKgxHd21+t97HfwiRFoIOmNiHhj1iO31BUJvnVBwJxBUDH
s5m6u0NWFCHgWnXXlxPIRsZx8idWDnPS0bWy0QDHYQ2swmPfIOnJoMqha0c8rGxB
zaOQxIGKGVvy0QD1dIx6Bbaowi8EtSDj9EyOIkw4Ky1v7vo/NLmdx1H+YXy5m7aC
Anosy1UPL5ou7qm54C+u2kJlx71A7ChVKiAzRlgNTb1pK46ak9+TL2e3+XfhqB1W
lt6JsApfwkBNCOLTV55RYUo6VgOpZbImXRN8eEDmmMlVOP9zBU60GKbxiAY6x9iD
anILEt927OLapO1qj6v48RboL/um+FCYwkPscw0RW8Zh6iv4xf1CY1ciY5Y+Gye3
bud23CqfKEjCN9BRYBP/n06nI0VNRNVnMdIeZHWo1cITm1WF1QyZI8SQEx1y1587
Q3VP1vL3eODzWRLxLDjwFl1jcgL1zFA7zHdwomR4R8Tucm07nktodVcNuLPeMk6t
NofkaxNeLb+Lo/0O4b50djZiinWtCCbaL3fe//kSsXSaNWK05Twhmy1mfi3fEsOH
9ySOvXQN3zFGR15V5sjhRcICLI13ZQQt5FOwg2YkJ2z2Ln6j1OKLktnVh+bblcL7
AjAChyUM5PSWVUzbvm3YICo49EqlVRGjAI2F0OUDMjMp5dAMrdcZtFYy1PLms+hq
P+hWD+Y6fQz+1Of58srzNN3tVKYta9+iyJVnRQx9ayTGWVxnjjnTWVRVtctdWsmV
ETGqRR/lvVMm6U8BeIirLFgHOYdezd86oDDHMVG2ukwVLx2mvOl854/GUkNhZ1U3
bmuTHdAqqlYlLIX0mey4IIN1kHh5t7vB1laTOh+yC3uta35csPhAA16tgjo6se2d
amkJ602Yrg07TA9o0b2jZORFmX15wvpm/+otLeKXzJDdoGT8WgMqsVOhsbPvf5RF
GgQ+mTiSbbfuzYbmsTIQDf3SLNudrZElXiRccL+RblYasZvrRtLJugyurDH5+x3V
r3B1aYU/53R7XPorCZ9E1wq1LNDY/hpLQVnRy3nV6rsal6hDRj9H8gs6ThNibC0Q
e1EO3NGx9wKN4otR28uZ9e3Qp55KqCWHaXoxpchHEizEPFikcJ1krEn2hRt3VYkh
o7cGMPA5NIrBzPIw3iEv/rvY+on2YEVmUWyTsOg7dWnpV526wLJa4ZyUoVTgiA1e
N4Ce+AxW2mxmPeHcIIrijEVbuB/wa03P7B6jS764W4/U4eeZZUZUmJ1TTmYhfSvY
T9TslH9KfhsnOnBtSDLsnp1E0oQOsKr393cO/cDYigFVMabQ5YjyHA1h+4zpAuph
0QuNKstBejeZ5aUZwwzyvW5NaCBfGLfqVLVbezR9+1wJd/zlhvyGiXSSXyJcw3P1
/d1iKg1DT0CECP7zjw4Sc30hmzpQL8Tdd84XjJ0tleMXJl40sKOu31d/hrUuiqIh
Xr6kZN79zIzDKOZcDuHZpgT3OVnRWlCaJ3egK+bDh6fUaaxo9DgU79Q+lNskRpKV
0a82GF2+cXnMv5qlmm1G15Mp6jpeTxxivQsYUPN+iEQZIa0sCnIi5dMkoQKSi/34
doMj5NkWj5wvn5CGX9drjNZxim8YDAkznnpqbIVS7QYprMcJfnrmCk460c8biAlX
anUlrGIC975Qowne+GmfgBO0EfcEPiPJvEIbDiG5PMz/MDEX1LHF00GNKLIrwEdp
zUy05qOPn6HgHKX54THf0XZXFORii0+yZhe9yzkgb/JCDz4N2jAa+UdCS5qSwjsQ
Fp7Fuabg1kNjUDz5JmOoXLz0vrnDmWbcuYRQFQTBnGim51H1uxWKFnUYmZNrGgyR
MgF4EOw+fqwAQnqa1663BRKTrjNfs5rzEzTXGSseoG9vKDhVLKaQKVa/zikLuBPB
V6V6dOuNemsCdDPy8aFC1QWK45hV4nKdKndOtG8MC/3tQ2bo3b6ipCUHTiB/BSrq
BBe2hfZa4gkiG2+9sVyQ4mquwZeAEDedHIMn3idPuuUGLYZHAXlwOqdqw6olEZtt
1JD9FcYS5REiXIgqVNlxNdYoY/KH71Y2DH+Qf5Kzq6NLQzR6rZmZqX7fqWzyCIaB
JtVHqE0lBFnb+eXU4/En8ubKAaDIgoGrw9wEwwKvXRSV31k+Db9zfQPsTVl9jkeH
Iy5kfOKm466LPAB4sWLy8CpZcQH5k0zNWGZe1el6yalstEFAIp3pSDWuWM371ZGW
kU09RKDNAGYQvXDFdMSr8x5LCANkw1yaJhbuRYholG1+6mph8Wa4eq8qf5Jo5kuQ
jFdwfSLwUZF7I+ShbBDrdaeDh2TQCEV/ySBY4ARelprHTLnzvsvnZg28xyHBrnH2
BN9oMSbjNgWU86hb5EPBKoppeAkbwbNfUWhPrrbvGntbZM5gb4U1Dil69oLWhiD1
xSLFnRx48znuHllmRTdUO1icuMMzeN60FJLtZwSALONkMNtytVCEND0+OH4qabHS
xmKzKf+r2xKbqfzxbb1i9DWjhWY8x5O+jdsRJJjn3XL7c5ByLo+gooiHmF2Ctkyi
MvAaDiTZZx0q1EOSQM1s6rMa3lVKqegqQwKM3airKUReQmkoPmekI8KDh7uFHNBU
enRHUrhjiJtE4QVc7MHG+RyCwfdtB+5KHJTradcwXO3xsx0aj8pS5WjTMPEz4pl/
t6+aIDSMhJcKsS367y+4102Rjnc4vPB7+8B8te4qPoP5RMzpuIbR51QHxJ4JwPzP
vC6O2Us8+uXcB6vR2slYBiSIyeqc6Jfsp6vFTjE44FTSicrStbT7Wd4bi1o93zog
807171OEoNnEOaxtDomvMbwhG/VNYkEwjawvGuCwejDK2NuilE2nPrFfpbp1MyLL
AY4RLZ+xDiDa7oSavN9VzzGv8HYjzC+L8+BdJXz0RnNv0xqAGRNp56viwtyrvOHo
OfBQjLiQ6HEofzxDhv7qCHUe/I/NCLvqa96Ygz/YYGIxUep8yjo3Z7MOUFy75tt7
PQoDffyD8oabZjX1ECp/L200S/T+Cref3laKiuY4sO2h9ltAp5Dtl9alUhUGtkcy
i+ZIKETZpH+xcrYUfWpbzcGxEq7Eqxfi+d5cUbeA4aiApNjJlDmpbAdDwo8ZwwHO
EToaiVmvhqgj9qaEPZvI6z6gdmMWTd9aiXpUokyO3XgGm3hcN/fL0P4VAnKRw4lf
1ikqx152XX0LIs8MRhikyFdR85ratNzXCiYfZ2fGiWd1VQxfwQwnrvTFTXyzRGaz
SGmcsH69ubi8pLJV4y6MUkvLP6MLTEkFnTcCTR+v/yj+E/yk9zgZ0ktzOI+el1gL
r/v4I2yhrQExFaJQBVSV8lXIMAcj0xB0zjvUmEkm69hcNZsGwDY13vYmE18rR2uD
AwDo+b0oihElR5OXQGSoz8F+mx9zieWMIjcAdN7L5EeEqgDilfcFR9RVzW16/g5l
fI/B/OD6H32ErybSDggolmb7wzxOq8MaVxLm+G7mK0TWrI/kONLI2oB6EjRGHysf
4Tv7z4xPImd0wlTOkUFemdK9LwdwohjcXK+h7GEMELY9yRyuwheeabNAMXNOmNec
Z/q4AAfXHdVC63MgPE6VeunRkoa2+xmRAHiNwHTtsUzq4kNouhYvam1LZbHfD1eR
4pMic55qgqTLb04blt7eSlDpWISK6ILYyvN/7ZuZFQJkeZWvX6PwJbQF8A1o2s8o
orcIALNPKgorhinpmXN0LVxoMyd86jOprWhT698imyWDMVfs6/MKUU/wv13H9H36
hK2qysZDj6CAiY5vlWLrRiBZ0OPA+9nAYb+02TZP+ceelV8UF+OONv1uTJB2+NZz
jPxDlRQn60UuTGvMsiSZRSUO2r0hQC++sINGIeaujxsYWsL8t+QMwsd40EjmmNZh
jO/RJps+/lvfROg3jm4EQejagcZClGTOr4Hi5lQ5rYE6mKDr1zVQdJ02BA4wk2JD
59NdyNMy77p/nzqJTb2Me15rTvnN2jd9PFvFY2GeonX0sIm7pm6vh/myruXv/0v5
RUfnq3MFO0RdLO1aW4yepygfulOVZX89H3vlTCVHW4F319tw7OPRNem/7LMtfeqH
VJNuVpEOIDlxtauGEHGIWPFW6k/ZpfiHb5TwnAL5PVFFsl1tkoV9I6t0VK2HKdmO
bNeJNvx+9ofYn+B7cCKv5bJboqBkHZxXPaGSsPJiuN8qce/eKjP+R1cURPPtXCrk
CVoXGcVDv/hiklw7EArYmwazFxvPNJh639jY3S6ChRczFdEBTBjl6P7OmArU/i5t
Fz3lvCVsr7sSkkVFRR5aKh7TQxDxvsaDJM2JyT7k1B5ooQgejV2Qhml647Zy9J4R
YUomPGplW5UeQZmXKHAWAAL5IP78LtBTxScpuEhLq+m/z6AbibWXyQt4XpOe4xLn
MqN0UQZQetQgyTQJNOz3SRMYWgTTNsSUqtMgbw6yQe9H0hM7Mgl4P/ADqpzbmq+X
y8D9qnqtkE5YS1ts1q1nDKNebj2XrS6DaRhQnGWhdceze6bwctO3C/1THHMAGsYf
bWyHvnGnNAS1e1rHGOnzRp8I+FgrA7ZM3oR2D6W0bP5mxp3qw2/ANZ028vJw1QXb
dIL69s5cPcORqJNDoCekW4C5PEmxr3uv+wNztONxtqLfFqN0pzqSy0xSd0fLj9Gm
P1FzZ5hUbuGd/Y1ZwK4o+lscpS91YHE2M4049UzpkuJi9/n+NlUMLWx5iT3sAhZx
+hUPbvx0x87poQxOOqRf/i9bitI5v+GfBXAMDxVlwCq9yAjccRllkz2+0DvvloSl
wNe5PIjo4OI+1GPGM/16kOAaqgIyH6/wu3vwXG/sryh6mT6Mr+HRkJ9LXrXgU4Cx
ygZjrpQP/u7C+E42jXHnNVOhhBkaY/gqr6BBENjQo/8fLmhfO1Oo95yKVnp3huJh
scxLOq+7xXypnby6hhI+QyLsKSCkx9nU8Z09+0Zi5s9KWlu+OhknazEtZTXCLAtG
L1Xn9StOEc1BW5i/GdJ0HoA+ECnK148QzZ6QhMoR9haVEsrtJs+qYVBRAtPSFxjk
HUrNHO1atqbtoXiLHiqtzy93k6RfA2q4djlr7oeo2/bAgM8PNDih1BvMfCJwsAnZ
GG+vyD6kEThw8cy9OYmy2R8FzAub+IIYd1w5dnjlqKuC+9uZU5wBdggDP/V/vfcz
PwtspzPt5FeXlBQH9/hS51Wc+8ttqb0zlavWhRWUgoNwA6l0zr/4pCRuaOgiJORy
jihSWpk/0oPBuljplkVOl4KATZ05dodvB73UhY5yi0fjgXeun9GY+iDodJwbyXZM
tg8eMpU8fbYfoj/Te6Hr944VKiWBJCazE3jxbrei/PAgndN5B46chG0VVmwRf6/9
0Ch2zMzouADOYSftdWWcaOC2BWhITpVPrDzoatabX1VT/dTN7/YMC9iohMiGysNo
BQuHaqFLvYdBgi0UiML7rWrjizGgjQsiHdT4Ppy3Y19hE9AppW/bmrFNGnjIwud5
r6+cr/7j5G2lMy0tTwEE1n5t/CIDUNZOHHTcKgJ8SkL2fFlRJ7MX1QAesMLBzoHD
DLbPCOTJCxmjCKL4VJ+UJB28ZoA847QCYygGkz3uYirwOmoqgPPr/yEjcdNHHE66
zAMgW8MrrC8Ug30MWuQjqbKYv+AttHluaCFHHpBsGxa6bxad/c8GMh4IJw438Cyq
coP5Zua+ruBmuvrzmdR/TCf7HJKrXY1REAroUqBhyBxj+9Jdph41Wr8IcbX8ng9L
AfTFS3wWMN07ZKxptP6Z/EPMJHxDROBqGz9M3q2uaUGBLw0pRyFJ81SAPaQfvCpD
hJ+O2YxNVEvnVssiRp3MiBgexCLwBQUq54OJu7CfHfMZQVOJ9lqD3Is0Rkix3p5I
Zy9Cy4A4tb8d1onx/iGFAo4LO2b4gFl3jhdWSZ+cmOhv7uZmm9S7xT0eIPP/rhLB
vUk8DdgVcrsg8Ff/76/R6Gb2V8k9gkVb/5lv8Oqt6CQapOl18EHN7oZnVCDvh8zh
WoFQV0xmDc1JknyF/aY5YER4YatwJJLpJdc7vCt7W1xlJRO5yY0Lyd8j4XnHnvnK
s1xgcWDUYs0hb+y2LHVW2PyI7VwCBu9TUlbd0pA2jXvsryo7wA5xmwrqbRCxdVhV
uoslOL2huEsqddGwCV7YNZ0ohT4DcKNKS5ZMwaEMh0P/yrkYPjuaVvPDx5iSZ6QP
/YgpYtPTQ4FuGglRaay/3xhWW3zY5U1bieQN5zi3TpshDvvYmDy/TSIeCR5qJyaN
/Q/M486s1liJfuETVtuyZnswqtlT4276rB4dAOG4dMpkW9JLJQB3EupTBfi8oSTd
LKti93Z3twZjMTmwGC5Wsemy4K027uuQibfntoE8cae0Oh6v4DKP4sK7EYmkIDrL
NT8g+cDm8iXdOVRmJjHkhG0DbPZJcFxzzsMXFMl3KlLNtycvshfwtlDHUtbrCicL
uRk8P69V2Anw1KhkdHLWlh7WuKaUALFZvfLFzLxglw6U3PZdl5jKP2cQPpPvAK3e
nrvyuLtT2XU9sA+UqQUuzEiBVhWUS7aFfnyMovXU1BFesctcwbWve430GQurpucQ
ag77TEPtCVVtgA/cvnEkyQJVNNBXzhN0c70Z1PPnI5vsdUcv9TzYCtjN/BO5TXWA
waRKwplpfsLJFfdt9tGNp3sKZ7Lv10PDd/6xo58H18Bs+Cr+/eZV/to18mWIz9H4
zPpuk/sVgKRI1qUMHxAf7w3BWJg8WlwsxfEwJfI4uA9HNxWkvLd0R5wFzIfWiuWS
XdJNsSD9MeZhnGrGSCzJEmDcx7oHbb7/ltmvUgPvjhWqhw9+55vWzf2rbLOgXQjA
bZkq+aGpRENcJmmkKURb2ga3bQjarB/33y30coVEavMVHrKu/3ZWWXtGHUHZrq5I
UgUoL2M1JK25g8AhxzaR6skohoiu9CbBfrpVj6Ojwt72fW1nFsSKMy3iJrwoEag0
0SDQaC73TO9I0vQnUFj5VcMAAs73VER/flYet/VShQ64tLMEo0aBjAiKKpaQjwm0
qqZdCNCIal/gQpD1KBql44Ju3eQcIr+kEg3SrxQj4spzOM9jwPfykqshLYMInbDy
kYfNEQVidFsqEH1BrH5L7JlFwAZJy3mHgUnURZwdmztQSRZbGzsUnEJV1vE9g8Ae
Cxz/SNJELqUErxGqdKA0Wm4FTORe9/G7TL6IJTSZ8Z3Uyp7tcRND7AsUJr66upv8
G5smnTFkfVu+SqAl7nxO1fP5+IY7XHYWyhfCV7aWBff1ow/q948aeC+dk/X1VaFE
34YkidXAf5i6PWR9TeElTwMfsvCJjzk76NyeaObv13KKKLf4gQ6QCrh2bxokTi0A
aAUeAY/utimNdSx/XQ+1UblcJi9Gu1X2v6KE8Ry3XpZdvFqlW1pGdHWnjTrUUuzz
eC4qtATWG2ZZ0tRTh5VfQohQoyBDaobz9iFmxEHCFOJwY8F2aJ3gMsRVIltR+yN1
5eUppKcJrBKXJLKGy3FndGyo1lcLdawH32smHxtpCnBqh+NnKHFvKWGRuhZ/kGCn
9TWpzzza3Z1O58Od71wgjcuLImeUF+8rFpbbb05Xu3v12/YGX5JeMU9Y5D37HX0o
WA0GafKQ02McVJN8EBn4yRKessX59+34GtlWhNfj8RTwlplxnHCpHVz2aZTddb4k
hoDDcg3wbGf3yVSdNuDYtiMMgjfnWEGiE2prGEDwbLlFc4U4oXz3/FmcmP6aGpOH
+KAHhG4qpK39rIheW60Q+2cdaMv3uzvlraxDCh3lsLCeoxDvod4KuDIRziCFNLZs
3YbnstNBd/s68hTJew3lXfqAi/ypRf063wc2x/1LDuEluraWDVaqLnPA03NrNrcF
KaIjwvXCNbSENB2f5TETKzlpQ/eUrlyV6ZQ/e+6p71I5w5nIpYnBDnwDowmdDuMJ
VZ0JZYWzWIR41I1ryQI8jcNrAdWstnL+KVfI1AtHzjz8GCq5BLRqD9MDBD/nN4kZ
JVfLX28CAGe90tEpanXDdsHkdpJ7O7a7BeBCQc7WF9HKsp9Km9lQYlDD8AkrjnQa
6jSAldqVulxPXo8/hAJEHEOTQBZBMKmfKlEZ31CXO+kktgxl2j/ipzVmgfz2iAo/
iOq9U+9lA6wRZJkMbwjbzddXlklqEFD7M3O4XYCtInB8/ht0eZszraYSCXsm2Lg6
Jn8J3lkfY6xsKsk6AdxxL1MrRBDdsKw4qMaW1sYSHcQRKPnsAWMGUwVu3dQT5+ne
BkBo+REjqa6Sw4r7WcL699yYpivKJt00COmQ20UrvyO65Qtimkv6oNZ9HOQlQxMP
/wNjtA5vZIEU1pR0VhpE+FgM9OMOtUvGeT83laGRycNg1ZGwfm6/O7WgT1foVDMh
VoDtfTUHeFONYbrh1uf1Hj9kSHqvVDn4RW3XAQOAUtqy3iG4KmcIsCpsLoq71L2C
uAn9wRZQvN4pynVr0qDDuSFkZNj6WUOc/u0eu54WSqwwKD/eFSLhGo2ZdbZ9N6vB
JJrX0rjBGrfKC4WK6MyBX1q9iw5hxQclGwFT4PuFzwwscTKqtaB7Wqx6FHrNPbi5
9mLCkRveU7w4yo2zhPyInT1jhC0/qwt6A38T6Op8wrYkOFOSBgy36BP2lNACq96V
5011NYJnW3Z9V6s5Wnb883DDXih1mAeSpHGcVZnPrxybKAPT57Nar3wrOAUGuhUO
J4A8xFmkzyu21/Qz1c+OWKVskrBknYKuNE++5URNYz+EjdtQ1cgxMjk6D3Fv9T7H
tbFo3b/j1tYqdfZuTcWMEJkpNGRwQfq/2hlNjJ++GD6bDaWjnYHxkDJaCgKcDTOo
wsXAyiy2g9UiWhDaSRWuTpFbwo0tTUjz5Pcencdm3FABMebbBFxpvXkVMyndjMqO
f4tQ0XnCTwtwyglvWqQV8oi0MtricNMnouB7tKr4iaHo2di6TNZ+YDSPaHOS24i7
WKPYPUWnv/2SQUMog/vw80bfFoItLUYt7HUMkXiBIbQvEjlrr2jR1IwBspOhFVJQ
Yq0lXK9nWhnZLKO/8ZzJY1Sgftp2ySka1SvU+Hg3ssfR9/xKPG0jK/BfHIzc32xj
kXjdP1xaXtOiPArp7ZejdF2T3HEohr93yIMUgTnlBtUz8VeIAdjpJcmxDBmakCzH
QN73PcQ+HgfUu6pSkmAIY/we7TFgmbPl+V41NQcIwjaQAQL+xGcia9bot4IBi/em
u3FTiE32SguN/tY6AtjkI+QsiNdkJJOoG5+f++B6FJ8Lt6JqvYsDJjkWp9A8VhFY
gtJvxf4J4TIALWa9HSSoMZFueTGFCFU9tHMq+xN0ectlRLTwwCgLLTZInkxjmUek
mvzHHkIMvTSHbZ0sn0mrJ7gyqASj07NFGHB5CjBbtbOiDMPfm4lwtKiSM0tTevkz
j7BpssTea8emthD4D4ztB2PX/c5zaUHkwqW5fVpMvb6XfQcwjUHvbh9XEO1xHkIB
sxd5MnueCj5rxTL61ce+3M/AZr2+aEWZ7ZepmL4XKnw7VhzGsoT7mLfrLirF3mGL
nyuonMEGc9oLKH550gJyIffJSKR019zbTr8Lt0ofGhaARkhxPR/hoUNyTnf9GhQ3
/hWtqk0zmzwWcm+HaWF0535PnQdrr55zfvN+OENzcxLo+6dWiTjoW4jg3Sda7EAd
u4fp+QN0wodm4YVC6Y+aXS/cE9b2YzbuIJlk4nhDau74mjq9tJJh1W9WxKgdEKLu
uGZsgoIYIsTF34jIAM5UAf7qy7lX3SM+/s7rOAqfnxmWS9HZD+SbEZNGJuCnHG/1
URZdYwRG0bISfuIMFysEoSFxV9uu5dk9YVX4Iw93g/lQf1OUET4a7UdfVp+cBVid
q1Eb0zXr/8M6Awl9pdMWh5CfS8UIyVR0pACh06U4q4/D5DJ+D1+56wQfdK7rxLWa
oIhyh1ajnOwqEHnoU5axDQQ2W34725u2fVTqvnH3PC5BpgBDlqu/KsfJbglDrA30
fcLewPy6lwVgf7KtcdLYnx+GIoKrZmR3yD9+/RGX5GYuzOSs5aoFXZx56eTss4AS
zQIptP+sYiMDS016OoE8RfBHWqtLooIJq7WyZAoc/68CtBwBI2Ncwj9L1YQ8VHEX
tiB+ExM8wZy1yBBPkn+83k+nAnUhLKC7fXdrhfOBsqSG6u1PDClGiSvxGCt5lPmU
7zv2UR1zuQXoCkGs2NQUbwwgFdwKefXujewcT9t+rzMvbSPPw9DPhn+N8TZB/jT6
6+tQoquvciYhkiutpA0r1Y32TQeewAEB10/TAurLx0obgjT4zPZWuZ2Fp73xILDq
O6nm/gFjGbhL7lQ8Uq5xhFVGvzncGDko6nBMfPVzlGR3Agq7OFG8W+rd2qaoQntA
Sx2LY74hbu8sJ+Wqvj8S4I5m9kgdxuEFRdytPVSO0p99FZm9L79QNats3rzfNC4G
jk3eN6UU/mpDZL+Oa3NO5Q+MYE1nRzbafFVRKnu3FH5PNceNr+wcZHGm7bYEosc/
NP3nvNScJucOl1et7tYxdSnKU3PmDkcxqU12YagteeIKMQCce2eoZ+uNbZFl2hBH
zcUb6fL5Xypu8QDZ4JP+2lcnCSR81oQm9l2wgfUJ9iCFIpQapaVvCmLPnVQPAwlQ
2idDm/CXanwpisWYiLCfD/xgZL1GIPYsNptjyA9LCV/srea0QhofCbRSTP0/hzxe
K6qWIDWjDVT92d0+QiAkhbRSMfz8LZsgQESHWwbvLxg3Y6tTGjWSsWLbx2/8LPMT
1o3QVLZr6FYJBam/lT5/6UqdNkdqLdvHuCKdhn4ro4gUIUFMS7SVtrqXxFCbLxTT
gY1xPp+vmh2LMf1Uy8GNXIsyBFZUF7Ij7XkiheC3rq+t6QFsBRvSyCR3o6rZB6vv
pTopJtjyoVo3efySTR6t0j69jrc6JIiCO1WZsZaILQmMyLrwIHJOkvAeh/SCRTU0
EBBatwDLuxGl4Hw3NXo/YitCzxudKi8tGMd9/ZPCq7ds036MHjodK6rd3D7dUjIv
gkx/vOcwW19A0nUhw0rORmxxfbd6odGVXqa3J6cD6AtDuq7SbC/XnOSgOnTLCQsh
P5mgvOjLHgVdCwAJtQQ0JYEqr+cwvO1UeuyLKIFWfDtiW3UwrtJQ77IEJn68r8XU
ygZfhut5VufcasePd8Eifx92WLYVp8vHJSwp26TIWq3VuiRMbm/yQe8wffiBsXo5
/AOFytEbdgfOdx9fIVh80Vz9KGGRwaAQeCWRCXMTGgEaZTT1+xAJ60/3fBCdE5Ps
R3naDOXjmCYSt3ZMG5z9qzAYEcwEsK/VkqJ4u+l1iYQgHr/MYBJ7+yH5EvW7ZLa7
Wk63CybAw5ysJMrwsH184UctonT1IhtkRG6I8HFFumF5C2eaYoCKHN8Z5uUDMKa5
F+deGp52XDCvPur85QwR5u/GKlihRp9n+Zg/DORksAROZ683/bpEThPo7F5be7yN
7H6po6UosecZnksYcWRHZyTuYmqroZwGSe+513GLfdkGXjacowLKNeHrfBCjHHLa
caCQW5r6xCSvOOTAxwcwkmB3ZfxzKOW/28UOkPfhohJmQgEQ6rgzzefSE/ObEwmz
J7nWLUSYIZRLirsZMYa0guOkdEIRVJUeYgJNioMabH27B/baDQYwUvWzEMRQYQzf
kAgUpy/7Um6P6CZj9yNQoIiO4bY+oe3nC1CYDtYOCdCDH4mmUX0GdRyP+pQbdTl1
lDyc4MTDc3CC4ya67YBMK4oUYAmHmNc6FieHrv9SKujKh+ydzCJAkZl0GxjOl4QX
FfR4KMbUZ8PzYKDusM2X0X0NmYvV9oCNj0QMeyRO/N0ravs4ppHIKZMGhRY1GnX4
YQIAwA5C81VORuexLjnBKFIvGgjKkHMPyDM/5/xFdJ2NkBwDnM+KNLSaMpGULIX/
lSismfjmp1ng59E5A3cPA3VaTTYf+P4gsRw+YG+msVAkZGyWOknr9xD+y8xGDwXk
sytVnjS4i3og9pvC/mz0lsJEl5Z2OA2mpxzXPxMiyDJ3M1J+RhyJ5P2rLa3JiNNw
YuWpORipe7ZPSfzEW/N+PYFgXQFb7Cv3Ej/CUURXb0IFwIx8I62oNZ/xPExP2XVq
vrheplqhAQqqrNUguMmXShg8I9CKx28t7khNcfnjW8OH4t0vItm1HzPZLE+3wxaW
8PhGWZcP+vS4DSjcgaserWPOyKMtMU9iGb/kavWwWHdQyutVy9Jei9Z1CCY0FVH6
/IVP1qLjxmGPpGvH6AcIuvVa/sngd3r8devbhpifhCol69hx/7SCRwDjG+gM4FqW
+tYXZ5Rq04SsOrmFyvS/uUuCbqt7WsLTzu5QGFftm+iqZhyuHAKqOmdJFMimVrB7
AA3kwSHczbJqJDPKd8iZi30FjKICqz3ERpivdkYiV/Y376bcpjaSWXKNauubZFvm
1LEN0w7pvmT2wbUkpLoa64IJsMyDtbsHxqaCg7KfFfa3LhJIR/VLEoZv9bqwXRw4
G9g6xHIBYtB7bdz7r2XzMgnRxg5+1auI9EXh3bM0Oq007IW54Ty3W8zGq4LfL732
xSAgh+s1nbl+QXIGMWyO1sG0j/f/ZU4jAatplIDNIu5csPLNFiENR31RaqrN8RGO
N/nKqJyFxcGNRvH4kJzhqM6zufTMCHE0UWWaVm1JrYegqOCjFCaQTOWqj7s14xts
4kBG92+26IU+LOLpFbuo62oMIJN/F5648X8Dx8rvAhQTHS9iXogH2yDCjp3miEOm
nRUr1+qzeETNXjnyNjPcN3N7aSd70TOTKd+6RG2LbOtuKKCC1JrRVbKNOCRDOfUp
yMJGNCahhXt/VT5i6xVj8e5PBi6Y4Fdz6rGwbxtyEoF2OBaGooy+qkIJbaIWm1hd
8mWPu+poxTRmzm4e1qZfP8z+asi/wkaNl6gFfxKdieJgnd+4rRh+HnFbimrixX2r
8E1TXI8bXLT2mudVyItHQvhltc6GGWzUgbgtXTNaewb4C/s2qe+On06HNJg9BHkc
b2dZ8H6VxRbI9pwlTkmtrH4418DWUxvpQxUq0NVScsKnACAJH96FKIt4Gw5iN4rv
0Z5jswJuKOjWVGznplmmdivh3pohcwZ8R2NsfbXJPFyXiDvsmJXC9nwfME5WJDwq
XgSa+JpcmW5rGQkEiTOGtuZcBN6EGgVMquoL/U4akP9mC4C4A1jAcmCZHZvm725C
YcYDKQcWIBSPrWjo0xHDaDCjlcZ+P4FAUHnh8I+S4LZvtIuveVN9f5kHtbdBtHvF
Rup/fRYdtko/5zzyrxn3A1IusM9CWRexENHYVN63ffJXlt+sNny3qDxkphZYzHjO
Cg07TPKz9mrZPr20W9nO7EzEw7UnT4IduvzW09kMaVdjfoS0lfeherBe82qhYpC4
qJR7GgkNPFt2IZfdl+Lf9l5N8VRCokPVL0yQDz4e8ANGKUMxNHTD43a2p4J8kZHQ
c9WFwE0lrOkOCtqJ7UNmSEhSlG/cSZ9R6I4ZvPdtI+wgqlTAww3tZ2hMpXagDZEk
oy1OONRd4rGT3/uPyA0oVMv3Cu83EtGnop0R8md5L7wCHBjxdWj62q0Z8z7bbh5O
KbaiROPY3gJ7qveaV23zTEgdYUivv8R0BjYJboftKjzCA1S2YZQr8O9bbW/crUBh
16gqUQm4IUQRXltWa1yBHCBznc+ywm1Xe8O2etYPf/QixTeY25oAAJ2yBDuzZ0kw
qDnOtq/K5ll4lnhZErSOPpoo7ntT10pzta+hm3NPaveCKmpYOUZz9pgfO6mKLsVp
CSdJK9vNcnMnBLHjOupkQi8x4xEg3BSGZQAhrDfdxK1FmwRbSJuwe4EfIXRsWO1f
eiB/OV0HJOjWv/whv4RipCzhM15VN50R0CHOJfcWSuG5GojuGPYDeNvj7qlhrwK/
FWcKfDhVDgioKIuBxXbFzzgcdwLzsx/ERvb4zDQNSSJkeDYbPl7YBREH4geST+9r
eKCYBtSVrtajZ4NOAnV5cIMJ044D8YvP2UTk08c6k5xxMh+SYfiJVFZ9r/EfHDFu
6PMD092ReY7PvQcvZNEXRVsj9LXEMfjACXMvFQ+8DzUmZaP3DycYGpNiaMKsJVOG
Wlcl8amrHhBdMENEZQAXWmyB4sPKrEjVev2wvB04MvLKvVKB9eiW+6sxcpdYVvJw
jzOqdBc8Fi49quLwDBNfYbmO0vkFQd/qwMyy4Vocodnj1MU3F79zL4WFMb4gmPdP
MHWtsB9n8AusaJp9xWW4xwaCVLttzQwk5K/gzJsxhT1rbCQA+QDBHQk7UiR1fZbB
aW6M6sHeA7Y6R4CMFuMZQl37E/AVF7koP8Rw2RX0k8oK0m9jI5J+zuSn5K2dLG3y
/HDoW8yXghcU5kY5mXMk1RINEhUKq1cKRV8X34CdvnfmWAb+PV/R/3MBVnlMPotL
cPqE9TDcn7vQw4XPGmYHrIp3N6KzasdLzv05ITV7CSdRA2UItdkN5Cva7mEEuIFF
iOMKtP+2gfQ8XRAETo/ysflpI4uOEmwflFSq3hItqrOSxCK3dazcclki4r5m4ah8
03vCp72rUMKB48Q9S2WJaB7wqjmoTgsxdGuvBdbW5Q32Lgbk6aon3CJFyiSj8bWW
YpjXVoG82gx5GFJpCncFcmjQhDiKEFzyZBMnaY+qMYM/4aj00bGRAbsJ9Ki2+VO9
OR/GPUyOw8S0XxeMlKQJDqZBGAjVMKZ4Ze2gk5aA/QffUb9Hl59xdYX7DZ/6Rz2K
evHC96c7nGgmscC1gIIdUhHYfAi9g5UD78rVb3swsMGcUs6PiLPg8K7KlsdxOS5Y
HxDYCZH2aLo930X4+SR610n8ESaaI1pY2VEWja8vglrkwIPqec3xyjiFdFpgygGg
5wyu4Ffe6xHMD5LD0CgY4TiUbtRVHHkcWziY5xhaonTt6IPSLCDWa+4Kta1GYSIa
u+VMmUfB+2MSPH+6QVi2InJurCMixVkwxtaHGh3BapkXKxhG/Z0SGKqK96bSDHoX
DvIhRLIxdNwzn83s1f7DKVqVWIKbxzNTpzOGCYNUnmiYpvh+PEmnxXML6/bohPET
FhGWO+qyOTOKs4vzhCgPLt+BiCOU7ciRAOXUeEK7T9x5azZZp9rlUSTOLXIRkO/n
g+e5u5p/T7AQ7SfiFQlVetgjqveGnRBHvcxHIOTwkyIjnb/hlMXWsAauuVXXnOwB
XK/Fxsrj3HGPI0XXXd6MEZRqremMipo/jpT1Tq/m7XsduiDqJoLt2PnKnRSn4Soq
+J8X/e05eUR7tO0AF6/KK1H2HEneGNzcqJ4otxgikqHEaIi/QZAUfBGJlOWy7PjE
uUK7ztH5xg1sgiZPdiliQwLSMp/YqJSaWGllsoNWn6RrpVdLeGAX8LNJFBIR3KWp
w/Um67HFH5oe3k4+upgQswAgsnv+OBhGpJkOageNjfFVLEjJIXKBk5nEmxsZqOYW
8pGp8D6A5wffyTe842EPKTkmFgw+m2dSY1v6JgFXb0Lcp420OB7U1maSH4ixhFFD
GiUgOJdmeW2wX7KjNIiLvR5/LT+Lh+Zn6FBAi/qCnf1OrP1FnLb0Ob/X5XGpznI6
OC8HzoLdCvaZvYCz59ykuETEKzZlSbrOFP5ahkuqq6OhQ8MVQxzns/nfGMIXLQXf
4mabrGg47JoYX4DRlQi02sgGZQeXtxtr1S4dLyejUnKn0cSTsknL+SQBr9WoRhqI
y7+Qe8Thi5MALH2N6jjEjI4MLSVePEF4BgMkFA4C+55xUYIIhw0QHfhlIenW3Yhr
yBoQSwrdHzdvxJydTCVhp8Fv7TA/6MrJoKirR0SKM1Lbq+Cy0FZkD1JSI3vYtx8Y
Hl9F94e0Ol8fkN6wajEFmn5CFn3Z32kwkd1yOk0H5E7hJSdG7djDen6Kh4eHUbvX
lzPNUdqgV+fDvqyoGsEwMXs3asGXz6vs6VWwds7/8A9OsXRmd416zDoR0e3U/6Po
CI/0L3FrvOmuXZJraRBHl5BlTgwUzI6AV8DkBBoRcQypO+IfdzGNB0ps4v+oi57+
D4o/Nk7biNQ2903WPsj67Bb7BPB+IJ7iOsCAkEckjh321d34rWqcAT4N6bvqD8UN
JA5fVFHBkgRwPRTD/fGrDLFYPR2d1aGZmPruhquoMLr8XX6EZ3j3cr/8R2Ey3jpo
Ct+olnWLstni2RT0/VSfXVi/Rs0Tdwm2e0zIYBu0NwdjLZmDE25e/dbU4i8DnYZP
m9Ny07fNuMq64xLxA/xCmfMa5fQ2+WpJrOGe3QBWHq1H2OHJ8HA1HYLNU1EWIFRg
LBMaiuy4KVLeggZYf+3XPNXyPJEVJBwG1LldZim4m4eNPC5CeHvKrZ/pBNIdjRUp
yq5DYii+J+j45nNhelu8ontAgRVhAmFCbSex4vqojqP5gAuEUu8C/EpOh0t/Ey5V
I1C9NOZVJm2ISf5dwdqrC10OISi50YhOKJatFkmBrTkTeH+S/io0YDhuoruAGaT4
chD+cIkQXe23ieabRwQnww3XTOrR8EphyeWrKRrBFVC7QILhFRWUgAkTIHQbDUyw
ORbbfw9v5jKpWtFY38BNRQg0xvM8c6nAqTUT8kz+VhYaeDTXCp7bqV4DNJJB1xxm
wrhVOypBL9Jp2vnoMtMxdbOjg4vdVahgHb/a6kn1yQnRpGIbljHVO1x1Z+Cj4uGz
f5hdP//SxUqNsRkYR5GKu3QGvNXQ3xY/qzndoSiUiURJiT/eyOlSK1V1d+Twrcy8
bGXYH3xGLzXsPpGFbMbYhh3t0XoNphjLS/rWkc500LJ6z+uz3AOlW0ijnVi2lgi8
LeIDzs1mD9IR8NX+BcKijO/nwOH31bdVZcKex7GjsiYZU2uA9bc6ZWwz0AtkXClV
K6tJK+Rr+cYrXYTMWqcvH9/SyCSlzsOTsiBjYrRYHrx1D4+dqBsmQTmckcpQ9P+K
/a4KCNGoC5JUDRqYlAZaKKYDQoslYKzpWgkt0J4I/zPDglqrSFsZ/5Lv+hohrJBM
GF5VFu6kTmLqSUIzQbbjcwK5RfHaRwYvTTrcYZ7B1p3A16hVcLNDZX+BbyL5XxYT
DXgGyzKVZp7YyypX95CgJfG6MIF8zB+CjQTk5nrM0Zfa2VWcYmF7c15dfjfS5Eno
mnpaaKq+cKs5NIezxV4dgV75YhZSzde3fRfe3uS16tT/RNvau7AetpUZ7QFLrOb5
cnL4VHyhSmH5o5ExrIHVFykZ1OxpvLZC5Uid6twdDCFEjgKI0cXtKBYME8Qnw777
Gri3bdHUVLIzcQHaQ/WB+RzJiT5x36dNIXnAezkatfqgZbxG4e9CAMS3YapQkfxI
/hz8vdgOOf1vkjeZ98raZzNz9c3PuOrkCc73TrWz6hv10IKXoCKyLpbWk2fm7CRC
ObOXElP4hioSsL4Frckv/k1Ih0aorlXZKIGd/1MnvVXB3Ps88BCfD96E0Ltlb4EJ
+3WV6VCrft+u8CfilIT9IbKAQQTZBXQe6nll51v/vFuQNNFMhYF80YrEHfu3koLl
Comn12C+x+FWOMGSiXP/vAUJTULyDpKqXjB15VPF4QunMIyIXXnh8z8rzGNPgmzy
moqQxjIQIzY1tq0jl19QqrAJFHbmKlbp9TJzJnIPcxm19hcMPFgGwcQ9oTI+oVTe
Yuoo2mNym81+m8hPi3W0zB9RU7jULrEl/nYvmZ/KZw20xw2BAgFHmGKaKHmIzD9M
gD2rOup1jtf2SBjXAJNtr53zCe9m2QsLYl7+EvcB4zNpV6XBa0tAAJ7Dt4Gzv3B3
DKzBX/qcyjgyZfBeV195BRYw8H8fUe/SAw2eNEijk6B8s/isYPDY6eCfcJopuRkR
rkQKpd6vZZE6ntJEGIVK/Lr6JlDC6qkafyoYEFJZ3uQo+e4j9CNJ6e50js3tAHlj
TevkG6wYWTAeu3rVORr96RthmVTxQlMmg79efEoT33pk8J/CZVSgCRwUEx9mqtZ+
yRv+gzqxlgqPcq+IGz/KfBtQwd9h2GsZ7RVZpKNttCCjbeRE5MVADknSH8KPpwhf
QDqZe+ph9OIq0kBbITm0xgAfeLl9qTo4w9nCSCF23mmOTcuS2Wj+Mvvhgs0MBOzS
QMJ5ba7/z4KB2DopZqVzjf+lJclewayLMO/n26pEUCA1OoyIDQQTkEAe54nteFsm
4pEtaZlwQis+Dkr7vjJr8CUHvPJ5RLAHP3R9lEusX93Ez/yKcMd/htJ89wWXGyqA
Hr9o4TDJnUTGersj2zeFrI2Zixb2gv9AIRKgDTpp2k+0O59fVaJh2E49YS0CK359
OgWdgY+UzZp+5GyRBjHrRnW1bawmVvX0eFzbxzDCuSNi1BJp4nO+4+4PZ5geWtaC
dbYK68PBaG+W/pNwp4GkW8T7PYP4OzGXgcgaWlwxD0Nh6lB5FGFxekMwwkuTjgz9
kUvk5eG0oOH6l+hzD9/LBlKNcNosEhY0ZD7r0yFJskYWfoO4FBOpO8cblEDaFSnv
LBn+unQB53IeHBRDKvLMjw6gQoAIotKKQqfgJeshEIF2flQjPebYl/Erzewpo+l0
cmcqi1VF5qs7yM4AH7fyV+TDy8wVcKGnl2aN6N7aVQqgXlg2yrTHbGfc+LQ5RrA6
+bk83il+z7bIP5D1/P9PL1LO5bDpGKong4ZjakKS8NBc9ImZH1Qbo4JrGBqlpQKL
UILObTwCf4WwneWX/otqe3CO3PNQaarjKK71bXIsZaK89sKh9Pz/M53oxeDDx6c5
qwzajZ7OEiggkuRTHjTRb9JyWhlLmBtOuX3IfjF0BJzBVbjBNlUG4BxRrxAt6y2D
vPy3D+KlGVXahkHUDawecB2e850pU+uLH7hWN2PFm0+qGY23NovDRNsfIvYn4mg1
lhbhiqAha9y4sWoWSDrZy4Q7APVKGDxh6ocul65Zv4kixwLkdHQ5h3Z1emG8tLpL
df+h5aD9QvGFLh1N7r2NwBWplK1ZtHgAqojLv5tvsBawYvGkpvHrWRvs9gF+Dstu
T7L4KwBARM8kv+TLJeWgBG2q1D771ovOBQbwkmugo6b8yoR43AKa4xx/2Tu4jiN/
zpGAN3Cr8I4688gX8xyaiySZgaG4W2t0bS8BUGSB0Gllroq2TQfSUbujge/K/uAR
0LyI2VuBvG7/fjHmq0tTxoTrFogjumAxAtMicdLi+7FTfHO7LLXgZeI7AvwyaLJH
Z+znQBAmYVBbYQw3fbIb+xCnYSFZlFP9eHBT6rgp/DU+c2DPI3S/CNXWPWbzd41T
7tf7NMfxDCIrq2JJgp7vqoo5RWIiIby/wdge0Xu5wkLnsxahd+cI/U3QoVvfbQLQ
jwh5+SfgknLDf6HIM4ituQI0cUlvBN/BwhxkHCq3uovFlN08Pp+eDG4AzhenY9VC
XjlljY9q6X1xrHr/RXVJSl1spE49wMdwImsRMHpoLhbbX9ix4cVvYUeXvWcUd2yD
cnMn2j9kDx1jcdK97Uqfw0fVb9g6KntzniEc/89syjzACxZeQTNhVzpU8vqijAA3
bIjljAO9uuhhlFsenmafBCTLOXdcjMWMO2ES1Kqbe/CU+h/CpkfXJF49Vdt9NoSK
1kB5VM66I2yAqz2zbd+DoNtxqYR4frxeN76aVsNcv5J9XcPYzY7/SnK1hEQSFzeZ
dz3xQjbeU6n+jqRafJ86naS121bOkLmlwYRHh0krpnrOSHbUVKsw+62X+7r1YnCf
0sXDX+726X7iLBnlXeBNSw7BqF2L7XBMfOUc6I7A/cN2wsytJ3ufbwgxI+Gjy9Tz
ysXohtbY3QDNbfI8zzLTyNrFI/vrHgAAN5ClnCW0ZskX4HuRqqUI4WOxyrxNqHDc
Y3IA5QAgRR6ugB88kb8jFfPn5R6lr3RQXCKzKYkGtNL/SZx+2ZDDbGPi3ihn+GIC
KQ4+mo8XksjBxD3Gb6hXhRlTgYjS7kKqwS4uzt5aD2F0fkY1Ez7nwIiSPgeRQRo8
gHFFFQzPeFMRtvLEKEKdrTEeBqqO0oeukLPDmlILQANftj3uN8qvKCzPRCRH4TiR
beY9MnLmIiHQvG4GspZ3htdXoYvtu8j2p0/icCgPH9gza7voefWbGYD88MR+J+dc
DxftLpXAK+7TzE/hHVd6QALakibXKzSL2XVp8zwyzDrFgeSF5HGTr0HGgDt5zmew
UA6sw+nrUDUpnNFRIwNTShAQG4Ht0o6OMCTsKawq6vjybWK3iCVGXAgdYfaIcP1J
/t73RdtzPQw4CD7T6QLRyZQdJVcK9ekX7t5yonbCvEA7A+0SrXEOHdBZLVMZ3CW7
UFbQZlrYcABD9XC/jIzGyziAbTLQ+7d3Qs57mxGVyr5W2sFtqf3lERvcOT1D293T
KOuclIhOzSY+NqzPMRNA89ZShRqqXdvca00hU8Z6THODUJRwGpQek9rqCnhY7cm/
hpxEdlATH/CeKJf/j2Txgp2dygU9yF8WOGlUohPEV03PkfBmN7HpnF8Prz6QsuxR
+YzdPBYTVBR5WW8zOJPWugEidrwO1IifsMQmcEZW7WcL7Nn5ZXudHnVonQ1HZI1g
9U1a84G7hBMnb1R9SYWEQUTOHYfVIqnoGnWQdmXFpp4Zt5Z/zL/mSc5PVFGHDtac
Yo6mfDaZJ/euKtP9A85h/epjuYVtIxZMRUuIXCWLTM+CtNRC+7O4D3AzwiaMxZt6
Zf0qhm7SroWLPo6AFH/vkNkSD0qelsJdAhPqFxyDA66/BDMwBjBjd9NASUU6QN+g
wYhJoaxJvYTHBuGWLqkPsULXwvJJr2N7Cab7Yrtx1/z0bxaNS60OzlvBXXEz+rlC
qYfS18d2rG5AnOPmKcqdFMD1i9/Ph00Py6oH49wVu9HVtA0zN8TI5Y8ad71Z9RoU
PTUQnkeG7B/iaGKJspAx3A9h73eEyH5foA/HTo6KEnsKEyCgHvCXhQSC4TeLulvI
wMkUJ+KiSmazXN4Dd0m6ae2bJTZq1e1YkXJPcTjsVu8l5NjS/SSR52kPSms/lom+
uZXnpvK763NKTeWhG/mz4BeRvbXOAJ1byyDfoxw0z7ETZkrGXisE9QEMQHECwB9z
xrHnbI+8Z8Xvm3riTnbw+Z6OKNnKfrca+25GdGIavkUvAhi8IfzLhjqi/h/TtM7x
8bJlvVX2SydHxmoeSzJUYLCi9hSCOEMv/hJ0FA18eHyOMPQx6EZEeBmlBcJ7z2/q
74DJ3z4yO3MH6BRnRevbcOM7iB2Bcwz+LY06FaBZ8tLE9vp8pz7A6zPoBIUUJriX
DmUNduG68ZnESViIJj00FHzphy4QYtuiNPmlqEymzxBrMsn0L/szDFsr/hFsQ9bk
JlvmW5AxqMoOkRW9ReSFoCHoR9KHX2ddZ8mJ3U/QMFufOk9C+n2jKNAGF9Hx50pO
UcZU8xSuKCXkz+Vq83UNfDs2mMce35/bUUj9sNxKM/hu9KoXNjneQFQHkrknp6c5
SLiDf7T/gUvF7RffQVvM0iOg/b1YMYFqcOP18x5TCsGLbmvYR+CzyryryjQQfAIW
HSElZQVVAgv9gi5LEm+ziYIe7hULooVBSGyzyw6VnbU2qFDacHdVsimIWrcpxO5/
iU8/bRAGu5+6/I6XuDl1qVxOl+CGCZqkusEfX34Evr6pxpYs+MdRh2UpvncSqJQZ
/LgpuGPT5TGg5qHPdhlbVMQ67/yHG9NnMXpHLCobP0WGC2IDD5WErfe3OwAo12BV
UgOGcxzloSillHAdPO2IHxSuXjtVLZRIMYPZ6S8j+1Oe+ahzz9fH2p0iT/O9iCc2
kwwqpimMl6r03/42Ll73K845NDBtwVz7NPmEyjMQMBabdz+tAzMnsNYE5TSzPPLA
A8jWr17Do510MmNPiR52fepD+DXk9HpBDW+1IP6ikkZT+BKUD3bVHay9+CedGa+i
xkw5w88rQiBrZ0tkzlkkjbo2hhfH7gqu6q13F/5BOaHG/DohWovA3OzAymP9LjPL
NciQNfVSdf3c41hc24mLi9+AVRmqqA7cjvs5lIBjNgGt1+A1lU7Ye3RItBAoLTj9
KF9c63DLxp6U6ha1pyXO5dyUJ4Ld2mwgrJivntPG40RczHAcBFyAikFwOvMhVCCx
hYFxOWXxudQ880C0S5Anr/5VWHwSHgtFqBtjs9422eKWnficVxe6U4NiQwQTkgie
w0StXX9JyVUYx6riGWylviFvNqw4zuwBz+QoQeJgmVsEvAgmNAyKdfuo3O5MIoPV
hBFTll89nREIc3qMTQKDpfqFMWlaD/IjCKntp9LKfuCh9XK6dv1/4E/JeITHyhYD
1fPSS35Rgb6qTNuqVyKsixARH7bMA1jMhkLGtEFzKdQFNzGFhGrDB/nk7fuiu5k4
703hjysvLEzl7eLwYBB3UqJedOWgkQGCNzQltXKkJoJTs0LBvl5issu/SxsWMW9v
RsDC5UyikHpy0An4bDgnjzdtNmmEaqxuZYfDV+PvcrHfsGeSoh+znik4hnx1Gmmy
ugX2lHL8vqW8hXx6qHHI27JV/ietrV9lM7UGzbZaJJkU2jEfqBSjSnABGt/Pfowi
1JetvKeCm7RqFkn/0xwj3jkwT7THpvnh2sTdnwrEot4b6DKOpQaLpA/UWGOmw/YW
PWu+ifrDZxNZY/5pSC3JJZfvHqOVSLixDEqsg2ptKf0wEa98ph/Rx/gDNg6V689i
PtD4vH2Se6Cnx1/3df1vol60Apr07F6qjMGM9DpaOk9Y9gHkUL0hdKpR21vF6csT
8Tq8P82Jet3XUnww+D+4ZFFBkhNEXEhdQWfuZ7Uo0cznMBdv92oc6S13UJzu3+wb
UygeX5ure9M4S/LrQQasLszHH6bVpnytw/dBmXnEraR+x43jzEtvBmIM31dtWthZ
05GPnh3QBAWJkYXOpKuFV551htgzt3BlCxufXwNwOWIjDAfK73eK/xd65J3R9WZx
wKn4f4ZuQs+RE0gRu5HJQCmCRF4zuzY8DogVagWR12G95sIV54xJ1bYK4QcYePMj
vWlfXtJ/dv2RkvwsFksdnunFyE5bvqKOnqrl29Rv0k+naESJY6WyUIPBiKtZBXV0
uHM50RmLJarMx+RIfM0cPDjfniCV/UKrFcmaBqUUSD1iHc9UDSWU0z7XVgf+3MdE
oETFyP1jyxN/8C1ElsPjii4Zk0LTQLMJ9gDeeMFPoIm38uCerHc+t08/YOHvnsLq
gZCzph/0b4rpJVesK9ATb0ANIu6sTneB200clTSN+Vd2OuJRUJ+CPUVeVT2MRhWo
2fxtvbbFEcAScF04a+Z9238gz6kbTupNH43NgeIKVRFxjdHSE5kr7oeTp5sQRJ6R
vw3hKGKOguEYr5l+vahk/CXlOzKOA/SotqI6e7hZxzw5baV0qNNST7JkjJmYf9jI
dkQJlHtm50GsuZhbSKVBslHSIcnudIT+5eBLWvcngvhL6J/msHutq1Vfz0WxUGaQ
VyD9Nmq/04R7J7W4ex18VgIUG+vgEai20Y829KmzCoupQTxeb3WWYFRwkRIUh0Uc
R7QB2zZ6HHQXQapucYmoxdl0ZPvIypaISRDL2GOUOWwapUyj2ZjFulYvCyW3l+4U
meixQS4GiTgzhilU6Nyl/jwbt5fm38V3rzui1sv92oUIbB7DycRyarnybpTXEt7Z
iEeCLS89EhgbPZblXs1HGNLb+R8R5sCccvoiXQncvaemdZj4+rh+jnIOzhUjKYZj
zO0QIBU/IJPbjmy/ii9XPVxouSD64s8nFRGez46gfPd/sG4fzKsBbn9a4vs8xaOv
UvYn/8BukrDVWwb89tQ3aoaAm38izq83dQzwGF8KFkv5gzKSVf/Gi0UOhr3y7zb4
EWPpGhCeTwJ+LTKyiIh9wymZNYwyCXD9gpefq9Ak/k4d4WSeFxdaa4dz1UhCudUl
hdq54mjjf90IfrQLyxp8qlIFsdQ2rD1wWueNlJWE9T4kJuIABBHKCoDDq1ZlF/Uk
6bwcURkcJivoPxjlZ5mhk7cf7it4NhKfEneAI2y2C4/GkCjYwzeBV2vLhQ+biqE0
NqcXL44GmbMoi8gnyPHSPCNFEGHUi1BAzeuA3gzODQFg/Gtd+a66DjgL9hCLlwke
JlGbK5CoLKfbZyuVqsGvwH/TM1Ai/nvEl4jqhJF9MJC6nL9XffhFpQJR1wbhQFRU
rmTREbeirU41xSfp/5GBvfO8L6pbRCmmRf7Z/pJ88yKYr1bnImhk3Kh5MSSoxMgp
9cHDRdIWaKLGXfsErGMnrI64R877GxhqN8X8bjD4SsJZT7MmrtIPvBGwlcqDunbj
/Znl85ie3mkHuvFWQACwUHSuqo6WeJ+6b/xiI6GFLOHPwpDn0SuELwJTBkApcDbT
fEtdC6tsLt1DMA8YGMq5jig0tuB9hd/rkHWtMUXD79OQAPKb5zeToN1N54TVLu5Z
f9gq+cgvWn3ymDv34k8J2HvNqQ62obUTO/yePb8Gb8JhlZ5hRM58Ghfv/OrqxjAL
3vp1EsTCnc7oEUQrE+5LLnKUUDFu061Z3Nq1mmqCGR1F4afABhtjetrZRixanLOy
QZ4R4IDx/13NnoK0q+zhHYq8ejkZVlBnwIUOvvl44pgtdziHzGv/58TnoUQ0GODZ
RJQNd36zjhK/wFWto2QqfvlECh1MffmPsKAxG8rjrNhAFR+ZDHZXE0s/cjWL3MBO
iGidYDe9wVzn3hai70EgqkiMy/NQ9T+zrW6Amyo9mvWyGdy2PLoactHNEunlLfJp
GjIxdRbOD4ZePUD/wRUROUtiC7zXpHYYoc+KDh4YmJ5qEkJhxtcjh4HJRrk5NrHn
q82KHIyhLzmWpp+qcvo0fIJA7WpE/zUKwUiVpmrhKH7KptOcSv8+qwk4yyDQ16Yd
h8qCLQndcDzi21lM3fl4IENdTAvARpMx9nhudJRiihbHXMcbnos/Ce+bSw8iNDFt
lfpzfm64yX1HRpjqw17MKNc1XvgUNQxQKYqbztOTVVGeXxOKE3ZtWtKUH2uLaZ4V
mDUvfydxvHObfGgEFvJp784HGbHHI/s57D6NpvsS++S+fw/JM6xvaTWaRJEiWWZR
iyNamQxo5p6RgAQFpoHXI+zTc0XNas9Lx/pQFQctwXDCuUaQ8/25ahxiZiERxOdm
SudmOKEEW8N4W/hOaDH2+LXDYL3XrrzKBhrbzb+7mbgHES7/n4qe0fjezzOPVlTq
bN/HasAOuUrw2KWuPYd1zcM6dKKuJghRu1aOrY0LHlM8kUTfUGqiWB9QWnPuXiD+
788VkMyMa60sgst/Rs1TF4U3AXNNXPugac9KJgA4DuhjVYa/9BqirvmiR02jpX0q
3MeSvazZndcovcriWoj9nI/hJMVKau2SyWN7l+4eeNcJHXFnzDr5p/PRoeCQw44F
30YqO4KFu4+QWst/uqSHrOG2oDez5oYYWICDy8/2t++kizZXALYeD2QL75SXMS1U
98pS9/7uiJykL7DVr2NdRVd/mBZW5OFRi30EmeRWJa8cTf61EqYg+ZhUHoyTF9GC
8BVC1SOfK+hXliL91s8wvV674IdTgLaRT6pP/Rv2YiKEkzGRiw5vWZSHM/m+iRQM
hCWO6bQ6gbg3g7YujPxE5zQLHOg1zy4nWuJwtuP4MB2+Xkmhea2RoAecj3LTKHe1
/mGIJjM9SfEgSZXHwAEtcKGUSGPaMVeD7VhJJabmSRj2RD6hZQt9nvlq2UMRpmao
eBWI9HuY+dcUJQopGkxd8V5EhyJpzM88AIL/a+87yISXzv4LX2Cm4GANuAC/uahu
zJmYibwONK6dTU0sRGlE3Ecm3BivQSRm2rKwZQlMwWPTXVOMWrN4deiMYVdFBkpo
WICPCqliiLSKafsgQ8eqliqqutRnnnjpjQvo7tB5J8gfJiCshsjn1F4w7mj6JJwu
quybhUX7PKqRpV+CMC6IMDOSRH0EYNP524D2O1+Rq1mpTR4lRt948TRq7GwafAGu
cXrejfXIKoMyeb2sw8MroSRq8yPPzjOW+uwDMBa/2hw+cV0916bN4ThtLyu96JDM
/Lv0TeJZ0CB685Ndts2wF1E18318bzBziKQ5dct4UygaUaI4n2zVtpdu6Hw0cnGI
tVJO85Bwm3W3bEyOVF2YohfXPKSE9e2PrKeBzQrvgI2ychKLNfH1pFfjC2/8v/PN
w34zzLC+Rx/9P8Uh8RqHAzx0XGNqL1VCGADol86YrOtEijvB8XsQMg0nUS+fiivg
f613lLe/Jp/1AjMVK2oKWQy9jsbmuJGF1ENeTX/R0/MhLMixqJA8jSDcqw0QZk3i
PywPg/++cuftYxXaxTSx2mgTTgcKTIvk/5CaMmG50dw36eE9PG/1PlINHHMo8hSn
9ZUORMClunAkRfK63+nny+5E0br0w4WcdUYoKHpe7PxVdMKCNR8gLr3/kmcSEpKv
fSyeIWfp1bCjnv3aCCy5Z/ItHPUmfXH+lI46QYfErNmp99VxeC2jo8W5Nmpkw3O3
dGaIjeDM+DNYz3pry5slOTQdg9tEFLa0OaxvUV5j9TjocvhMFuAicxRiBd/vUUOJ
WllzHlnA5FXhawdGt7Gl5PX4AfcLADKuwZqzzKDrdHkqY3WqVJod9q2AD6MLBtm0
qJhvcbmq0Jbxeqw1u6US6RDFiKQSo6Q5uRJvNJRBjW7/4pLNr36RGUlNcD62Tf5c
P5fLlfz8qcKKk/YAorHre/CLohoy1sqApp5nmykiD1+Fnmvn2cSQjsF9oo4D2eUd
wm1NrfiR8ntqO9g63OGs9dzq41BU/un34+lqWrJwHHErze5cvE4QUqbyF6HLWzIe
nRoSA6V/KUgblaiGL7JKuDKUyZF2BiI2uKpJm4d7/1PFhVz/cVo7t8SXxXr8EvXV
q4KMe97o4Xa4iFXD3IHeWdubaFiyuDOKoqo4w5U0y2Z28Ib1IrasgGWHkRRHkOHo
nDcOd7v07dNFfhthpdyuxdZPz39fUPx8DH7F1peC4iHYVzlqCtff9LvnR5GhiCke
S/dK6xfS05N8VCnu3UcR029N9EOmx5VNNs5Ee4daTOHAIyStQziNOfGwjyNYi9h5
AG3sz0L28NQnjcCbmh/N2A+2fA7cGU8zdzRcfMuj9z5JSFu8fbmG3UGGoLFvz5J7
4FrA/ACmCrt3BnQr507KRn1RA1UkHdXMSckNgdVb/w/XaA82TgecCpqK808FtDFh
8X2siYGrn0n3cgnHvma9NEspj/9bBj/GFiKbew4/SkfYqBWO7KzJoynQjL1hCnN/
wMrSBQ6IaHDbWRyT7BcO2cGXesn+YV4ponkMPSHRzzz/uaqcc5acAKFReGMngh17
nmOLOsXVh1iqpmiO4mBfjHyzZb5aAaRy9qo6b2UnB+OtNIBq0OPKophB+r08lHb2
asRW2zmbTIQgwfUCO9jjBBWS+mlJ25oKTWDKZAWgNapd4KkCTdYRWtyZoSP4ek3s
pS545b7GMbxLkdPIiWzl1WqaHe0/kwO3YKJhyXad4MVwOf5FcpyZP6+ssVEAXLhE
ohAfqLhjmcdNGJVTynBT40zisMo3xttb+fVzPuoia9xNVgVdp4vJ4TdUGtLpc24a
+Ze3LpN/kr0qjlIiBT/luaeunHzzFJ4yOMOzY/nTB1mwGyri9a/hLkP4vf86aTZF
OZ2gvRTzYTNDf89CxiqxbZFLD1jXQmsRejo71ARqbqlGNjg6enUy0eV1txJdrBAc
qrHUqz31pQlRhaAtbNk8PkugC2lkdxoohVxT6Snes6vF+GwzbVe9y1XFYHgc9S9k
6cX3s4Ry2baULRQLbw0+F+NP30WTzn1EN/z9kkVJQbaK7xYoFSUEe6TTPvmE8MAc
eWV2a6r7fF2BQSKiQuPh8ZBM4kxHw2ZlZ/s/CeEhwsDIPkAYtfiTRERHglnoTFbD
+seO/e2vdDjl5Od8IRY955exg+UATsGu6AvZHsRJ+N+r11t6ODny4+LtTu347NdB
TMyAxLbZb2euym6up9jxWYG5I7IcmqYjKR9E/ID+fu54sVtYfzcwDKsS4M3OyGcO
h1vH9JPmY9FeZ862TCEpuVhn/BZUIoro1tPUUuIfG57seRy/D4kDz368SKUNmnP1
Hrv1yMvno8xNWTzTHVpRBV13Q7A+yexal4mvXVQ8xz6gWmIw4LnJ8pZdxNbgr6Oe
myN86oFjtxVZnRjb8v62ed0fnCc45cGdGAKgisDBYtIaZ5pL9P4oef7G5wg9UwpX
E1CYr0OinRwFFx1BXb47VA9idX1+HyZlmbr1BX1qfj4N0mqh2kbu7X14E5jZ3cSH
zm8qXWDaKij3BV7EKTsGLPkvLYHNF9RaKha9EUX1WYWb+r1Lbvha7/28jXxPKi8A
2OfIaTBssbxvLtf+V3uIPQ39u+8iBuKhp0HU11N9oDbbffgfVGAGPmpZL5SjlhN5
JatLr57X5iKvASRXpmIBIUEPC4uYE6OUC1F/X4X1UbTNojYtlYNruTr2V0acGNN9
0cC7X1YVVZIUL+TF1i4Wv8oER9EIV2L+G+0heC62qCPGB+5Q8DtRJ6Kp8nJFGrof
DIUkpgwtrc5rqHPGhXgWK38DHc67QHr8sIFCZ+2ecVTsrJ4TgpbCqEaQyKlvEp4p
Wz5nLVcYXXclQTOD8JB0Dt54/WrzPT3QzF2rAd2CzkwYx274ZWdkajdEMt8xMFWa
5XYY3idDoDO5AS++DjuGQ3/rXjSte5AJulsq6kRJWbSM/caYH+/VUGSR6PJWCp+9
mbt2QVowOPjpkXUUc2NuCwY40vYfJXhCUilh8c0vRvDeC73r8GT+BRxkMisdWpPj
ggdG5Ery1OE0KiwXrv8HtQGlrStwjCl29bJiZ8hqTncbAFJxw1x8+DycTtfyvFFS
0mPV6ynmDGnRGYu6TcUx2j6j7dVA1+v3wQc0KRre1lfERqzV0ALWv3fG1SG8Ir5B
ral/bDt0tJMuor5sfGtnVOsCxT6/dL6UYHOdzktS4jSjs1x8YlykzZxaeY0Q24pq
YI6kjVK1BsHelU+G59rWcS8C6OI2ifMYrjUZYnP2gCm76CffqRAGPkFFhBAsYFXV
4uS1tRuK9gy2r6S3xI/ZmHXhGjgfA3cLXLqekKVoeLCM4kMWq9J7koD6Le7+qFSs
BKHyHwdAAIOab5PJYubfeupAWwD6xcfuwi5GblXTKnmM84DBNyS93wGL7vcOjB47
3TLDrrS0o8GtLTlqxgnqJqGdYEuFHeGZPwHQ73b4o8NUZe8xttB0lH4Fk23uRV64
BOhauvKppWCVSuzAhHGFIQSYJaQsQFAl2JtdOCa975X6nFD9UsC29G7sL3Vwh7Jt
a/mqY8acnvjlox7Skc3Sb5nDlMupOt3Yg41sDGR1sdorz+l/cf/+W2QnFvMHUpVZ
I3JqILUUGnrtvCQs6wCX3Msy6kp3xlXxnqDHmzQ914J0Crh1+cOdQy+oUkDajKYi
h1xLbM/9iOZCWAzqE80Rq3cwcRquPd5u/WVyQu9U8YAxnZjjmcK6vE0XelflbGwo
MLcvX2/2kV2L2iPIKlBeePdc8vBt0hGlJ0wb/sKzHvVDrtqEX1UJcK+NccO80nXo
IZ/yZUssZkpcGpQaf1MO1RfQnACNiE4d/gN9Uu2qE8cAiZNmzCb218Av+zY0nCrL
jyqrIGp6bEzMfQMrqe5o+To4aGPoDQWHjIzHiwVwrXt+mYSfCVL59CIcyeJPwR+k
Oln9vq4t0FBqbZ+YjuqlHeorT2fzrJ/WaHr55MfEKcvlW7uxsysGqI8AtEVmDR8R
rvlKGnl8IzkIEZ3W8WyMjYpFTCEcQLo6bk7Pd4izqxwqpRkMtvTifyYACtQdI/DO
kCg2KN5ic3kEMyqMKMU7J3VszDm8cVeeokmAMy+QrqdqHSIgPKSGaU/NPfN47Tmn
80h/4Pd99uIaB9voBHm8t6bCS1oPXhrsjqFPUe+GmPTWzFU8cPo0ajICNgwOzZRx
ilHQzH35uZoC0MyZGKdgJ8CgCVULDfibAWBIhfYWUhZDLsc9sC56AFvRl6niAmQI
iTgvspvXUg7JEOQdHEiesMFJ6OK+gwB971V9WUHHMdu/Ij7uj5bDRCGwN/ZHcp0q
Owrof6s9GBDPBJNo9E2RUxOakZeB934qcNbRYpttSvBk32hIp5HbGDJraVzfeyJS
WHYvvZ7eNUN61P3MC/mpMo51qKaLwyemGsk0yT8ZgzNJb/F09fwZfAzZalcCr6RI
qGrR6qycVU+u6pcfps/uLuBVPJ4DRvGoQsGr/zVOMXREs3Fl3dleOwCH65w7O3br
NCkZS45UxD9ciYqDda+XdiHc64OEST12dncLlGfdvJ3xvnXIuVC2x9P16giR8Ivj
ot8O2HE31Vj+mGFJi+/rjOR3XdCpX/zq9c8pKYakrXH6oZS337aEyGVfHjUAbDUv
45I9fq4Dh+J0uSccxIfzJP/a2xjnKUucXYP4AtAaAVpEZmnbyTY9YwzH7e/vy46x
+djgvTxb52Nloupui58CVq/1RWfCFsb+qbCscf8MtE76cVIcNgLt/a2fFFcwgCIE
PRyIp0jluJ9j7MDIoRnz4k9BVXD4tzYow4MpIiwzP+YrZfJimImON115RVDdYWbr
AGzynfNVv8U7eSSaNDZ2FH5PLchQ/ILc9sgMu46jZtGVNdtFZmfLW1Efp/Vz03Ew
Jk/iOD84HyGO9YmONd14N2PPdNLAPLqTLyom2QdT9+Msahkr9zv+FJHBT6iZu1wV
07WF8ZX629WL9IE7U6yuL80F35QF4sbdiEjRHHlWDff83/tZ5Rdt78qnn6/3r218
5hXtdmOXBSATmcVgVd4Hs310lxrf5cPeCvn3Q+D1TFPlYckpIk/GtrFtoA4QgUXO
10Ankb7Kkjxg/znUa1HT050DnYgt5BtoC5O8EM4gqPeqPU82gQV/0D82SwQ6UeDM
ufNwcafnMqiyJgaSZdLPrNcqodi1aL5NlMiPpeziCPEN26vtl3FuWOSfIGAfoAgV
eRUcQW6EODd912j0SkCxZgr27mEP/XYHcUzcgHXhKqDeFjt3U/cjycYmgYyxPdSW
n7/ttD1rzpbJaaVtmekccPM8PXIGdiNqDPAQOG5WyEe1oxkKNqzGxmXUlJONgJNX
5UXXPmHPUUgHJ0hN5RaDeGiZPiq1ReevxCdKPSle2SeCYo232/jeG7jlrSTJrDgQ
BgvP15cJCeyJ6413zlbv1EB4GLpYLOzse/TM6Edc1lyTrPnRoeYDKxChjL7kRhhM
YZH1XSP1cJTAI6nRjg5T+Egm6HJbo0mEd0nUWdLIrW+xedBL0CkY5wFDpBNdn9JY
LqOLT/FfifBVBw+7QB3fYi1GYhBQCxk9CiMOHeK5B5uMxmmBmYSbqPNtQqF3FUbX
/0HjJ2cTJwHM/N4h6YaUYtmcRptNV3Dx0F6LDDgsELazqYfGn+7BDKL8Ussd7Ea6
Yxop2EJIqByYjsxhO5ao6GB9OpBGdnJzw59N8ru5JTRVwlSmNgtOgbX3oiqXlApX
w5KzWpiNBFZWTwcJd5Wzotg8s4spcfHz0w+/6twN2o+x7U0b17rn7PsHIdFHUq+V
+R+cRfHlY4TUQU/MQ7TbmzM320P3XzGBvZx2ODFWdQrsr/0ZaB7DrWirzpz4lfTh
AQd78bp1b2R8rA5uaX6WvRD9qjJ1JMI/tZI5VitB0NGfona6/q8/iL4pKseD1Fa4
JjWXmnT6fZSDJRIa8/Mj67/uE7c2eA84CMhTKvDjgP99nFIdK4MvVHXkQT1A8+Ll
ZALk9PyYW0pCN1ueIClR0W+Djb/TffFgc0fMt/ljmprSObJEzxMLpqgM1/DpkSUF
6Nt5iX68n3eiJ074Mg6L07Yi06cPtoq+MGuUb3EITtpqPsMyxwrUb47y8yDBHS06
6dM5GkUPOsnXMQkGsckKZQoNpMOUxVTX/N4Bdgsh/azhFJ4ziCbXjQJfFZ6nSk+k
iDJkbazaH1kyNy2kwJBD57uCBhRD7bIY89yr61hrfi7RgGACbVxy/kCznSTxrAFK
xPzBhY+J8UsVq2stjBNvE4dAegJDPk2No0VTGn/paW86zUy66VeatbgHoOo7acqb
GQEQdg3jSVzc4xHeUy83dvSZjWWsrwqUJnueSkpeoW7VjavCqor+GG/FnVpPPP3G
aEN2T7BD6Cllie8p9Hivp2sShepLpSX2yBT6GrDrLHKRNgzaaeY2EkEcK4CSX0Gy
lUPymKGn1XS4O7hGeUtlllgvoJC3G80f1upyysVGEuRE+1MP6QlsshE5PczGAC+B
Pc0Xi+xNgDtHQUfvmA8Jkj/M2x6n8xg1wRGyq8uestbsrgCrIVxCGl49T8+i/lKm
wcsJtC9voXp+Hf/V9Rt3EbCzA/iZCSEpDquybf+aKJ0N+xdSBG1a9tr0q9joQV2e
1mmlupECvn1n9Ncu3Qyyl0fBz8x+xryjm2ZBW4cC0h0B1+rrP1nVlV9TAf76qnI0
971pAGjg1mP67CU0NDbgXCcovEXfWPP1oCwxUz5lMFbaj46RpFHv2ye9V3PmIRhs
Qcvpslj1gEjWfhpgYrDwqWtPMKGZ0EiOE9vDamKl8o3OxkjelMCii/NFlzyRBb4h
oovrajcJrb5UOzplJYMaBXyWX5QxjYncWCWFkY4j4MrDGxncKHWfTMwZAYjDkCLr
q1zUzYBe3U+jKjEXzgPBXXRU5gN7A1y7UBUByHUelqxdBe87auj2LOjoNvLkzpu2
FnbuM2JNBlu4eEnzagK6HfK13ePsEuMyjQ6sW2PR1tAHQVMLQJ7fi3l0nTmGh+8f
ZbgCX3MUPlO7+qnMQjD5Dk6ws9/7jdzDVPB/CW7BO7W3FrR/dMBzUsN13fYjvuMo
bKS3Fn8JoEUjb9kB1hUxeQZ++EBGHkoLdq5w0cW04StVQyNIpDMxK/v5Hu+AwUvV
+fm9tUPAwnGvqgL3V0Si2Nc6ebgU4JujQ034rJK545FMkKU9xRwntFLdNBy+M1kf
S5AhVflltN7YjS19qhbJave1n/0BAJdloh/EXhyPq1rdu17GRHsu0KGDL5/WSJqZ
K+xO2UfPLqHqu8nHkTkAAtjVBJxUrAWJeL/TqIainPqh6PiJVpaSkCQ6rRwdxIob
1N/jupmDYTvxBbTLC8z63ozCsslg3CnHAaCrylHB9VttfPSGN0rAuVwDysSRDJJe
Lm2mMWTww+rHesU2INwA7XlOdRSHTw9GEGAdWQu4+zLCdO6GCjI9AinABL9ESN8c
Dxe8dRwcxI4DlORsImbJzqm8vGO2BMlBUVWTAciYlYNk+FPi1YJrwOD4oqWLSqBZ
Tlh4aQdXd2jhJdHPdpjtXmVQxW1I0SDFFsMLw0lXT2CUbSp+ik7UEoKzwVK5HmPf
N6NtdUI2YcJeTs0Udtb9d3m3K4OVQx8S/pv9bvgpncM3Q73oGvC+PUKQZ3VWd8OK
ZIwUaFaQpwiEVApT3cXzYoYwV+xO+b2Qay+n3rcLB5sTF7IbeTmdf68zJaRuFg6d
ZwWFMtL6kfNG0ZlE+AhxHT5rFK8mPHY1H18zUCBPXsoBS7tu8nA/yVCU9iFEqWum
yheLEDTA4ShKvmtvaelxzHQN2k4d8V/Gf8uyruh1lOrwDsz0vhOOpIWYF1wfEwaF
bP6Eg7bVO7j124VqAVTz1l3n1oKQW2Hr3Lj8IcrWa8/et8MOyc0YZs7L/XXk6xKi
fyvknTD2r5F4TgrvokrUhpY62Ditez5zYB13uNnoOd35kDiJ+WrEPrxlIgck/03u
dg4t0Y3sRrklzQBOsoUMJ2cjUnp2A5wP+gmvEh/ejPpB8XiDk9Tin6sC46qe2/Ep
YknoVfSuwadZsLel5qJd16pEslog8AHcpGEgTlIqJIKUsu+MaRfIbvX356I/E7KE
jYBiBCmRd8pa4vxR/Pq7/yMbCkPUrnrF1vzQXwXQpAJzGhPM+0j2j3q+/GP9+e5Q
T6jvvCTsy0GO3fMs3ZPSvk2RPOxsoyzfDOqMoIle+dN8AQAhwyZA9fZhxF6Fu2V3
ZGcdV8ph3S4EAASjyxP3+j/z1dReeH70eLDlcj5+YRJQm72fb9a9UCni4Kt6GM1i
oyzGijdoevmAv6p+ki/43mEbCekKKZWfTi3irDHTBlcuAlfIxNmMuQsWNhOLgh+d
0uSHCQ/hpJlM1Cx+DebyITA8sZ24xQ1bV2dsOMgq4IH4Sk25oKfVZokc0vn0Qta0
GvcVXACexWC28Z8285HYM/LruN8D5kInHlcTV6xs0IrAbziKd/cTabIsSO3uZJmQ
qtTazZHLyfQxf87/BjKXFMC9RGAspvwdZ/o5/gemTnQv2SqyiiX27QYwTQFna6Bl
KWqGzxFVpJWSmTg83pipYtl4vGRxBfl+MPthTezg93iEnk1Af7/UbrqJDxYrEAVJ
m9l7J5s19G7gEBFUSvpZuAWzV8WX4FdqwUXdRO66PbZOqDGxGX891sHX3ql5r3+1
TQi46vf6QDURVtliazTw1ReUtbBofW1JjKjTUHGpwwfeudvxFN34LqRTnjCZzQ8T
0CDUo7bzcfW//JVLQMe8MC9uSpvpoSqQmzGB6Lo9/m5CsvM6/DKfbc7WJpZN+ioE
J6eyvN2NYwZc0S10LvUqvWImgA0t0OlCp9FRAZqow+t1BCgc2HK533L+5w1Ldi/j
8YZTScFm7K7Wo8dTZ5I5MAiOZiMZjUtAcaNo/N3oiHkp1eKw8xGvamAHacStjEkY
cGZx8Vc39hndt0fdtF6Bn5+s4MjJl0DU5Q5nXXEC8AZM7lPfbxuHJ1kO5gF+y+3J
Ru7CMS+nSvBl4G+1sBz3NPcguhE91IHbPn83spDlmlAYGxFc1vU1lhc+lQ+NPvq3
woJwxB0AaiAo0rTB2i2g+z/MLoSsZ8muOQecXut5tCoZ6UVmPiTnlTzwQRnMElP0
+gGjs0L6bq4Tw1GPh1vSjMoKW2wVa4g1FF4P23JXA83CmXhW4MFwf3pWdOVTKcJ/
reLaxTgjYwThZSSZfy9M+uxfzMX+K7Aqar050rxtrCx6+4NyaytILS6ToSRryBrM
IZiRsVb+EF5c6/WolsMLdJ1bxlCMc9586JecVxE3AYZKsQhkV+aesyVa0R5gNywE
rcXfLoU0RcDUBuGCP+fCHSo0jqleBgyJ5XV0D0MfzGiDfr6Z2cRsPZU/JUo8emaa
Kna2qBW6fflgwFltcHIx7DDcO8Jj8Vonsg8kqy2hBxzrSdc9deJIRtfDa66fSRLk
pJv4Poi4wSGx37gA/JhztgXjvXGDilOozk5E7sHt5wr3yJqlo46OuhprZonb6VGt
P084VldevIXZ03PNh3bRo54ilNx07WDXy0ieKhPnNhZ2BQL3vMDa0duBVhsn7jsJ
CEU9PPNs/k29bdtmc+mY+zV84pWaOMs2KwJ9ptW5qunrYBgKFpwrmDE0dkDbmstx
/KD3XEhO2yDC+sxBpNCCf5iwUA5rdMIbhj3V+yMTVh98YG8yVDyA9urW4HUigjZm
CfpdRTIgkS11rGGcZY8XIiP+ipqINquVlDL4vcaZw5zoqrecQbDc0kx8S6UWOD4r
Jeiytp+c25YZlawftN3+AiP4Tr5HV1cX4kDpbolhYCKm+jrVK/nC8gnquKyaJFGi
6SLELwfGoSZOIOK/DAwInNeeZSHkJ/z/2NEyw1ot1jT3S9PZLkdC4VlU74Yrej9v
ftymbawixU6k1ZYtS2MKncC+GRhsmsyJ1VOsO0jnC0RjdhwU1AvVnBP8oIfqHTq7
rTae7ssjpI31ytMCgsoL3hru8xTwm+NVHvuaLmqL2Rt2weIeHLmYGgRPTPOtQw8n
G9FWajswC6+pgt+Itt/S0gyOBwfQba38zkv5g/gg8EgN1qCOofFwG2GpWZCIZj8W
TGjYzd3N/0BhLjlxx7g8KG5iJZ6s7/Jb0fHM4+5jtKhz6vmKdUKC2J2pzcAvVloJ
15OEe5eCFqd4VS4C7HPJRmUZqEdGAjLgI6MT/6hmWUnn2d9dN9z2ihPjDeiZxo68
BisG08hRRabQ8GuuN4btT5AZzk9ltdSOtEG6/y2v1BzVUuAjq1bf5mYvwvHINxW3
GQEBT/nQttUA93uetIs4VX4DsmYmsh5e4ZPLXwfvMfLSsKLiPXnvlD8cAwkN0kgg
68jfThYl1zQVASRgMbnnZW4UbpO2AmMzyWdOTLxHbJYrSoeIM+XYaHWDKo1qyvaW
51LmUc9HE/mRk44j/VCzPjuxSrvFgP2mhJXQgiqRU28e0tNtwnYeAIe9t0bdR3y+
g+Vpfy3QViUgb06T3QvR+QERRZQSkQqcH5TxZk/wfVuCseQHlEIYVpC9DxHG6CFc
NXZ5tS8S5sHKukhlCBWWX49UVal39l11Fo4FltDpkKbm+hsCUvDS+Q7dQV6Ise3O
2tVVS7/aT8+XHv978rpbkqCwFszJ8oDgECeHHigbKQoOMD2hSn0xP79w7aza8SPG
9ojmEtc8iKBCwLCcyqYdZPryd1DePiTi4RHLaiTskq7x3PaS1g5ACWRApL232qL2
KsxLtf4dzxZVAmpU3GlnyUgbgvG9ZkkRAJZr+4pQSI8NaAZH2Q+iUWbUHEF4cRCF
dxLlPve+DSLGK0wElmRkW+pmmjVfm8mImLSJoJ4ABQK3LPBl0C1Ui4mrJgokcZpf
u5sMynxOfWrepKPDusfk68O9iu/rMWA36pW5Rdmeg8+JUk+zL7j5+bj8xXr2zF9u
/3W4gt75B+JH85h4G8ligbDHhv9BLq1fpOuFUWae2oDNUj/2qmhiXVtumMUFh1l2
4IWOBkrbMjk9ETSt+8e3pRWpEREGbTKqv5sWacoqdPmwPVx9/V+emhGLC7/3gqbQ
e6HfxbUDbb7mWij5uVorC5GMLcuuMUbOUhxJ2VBaqsPnZOvf9p9mB0X3ahL43t6t
D2uxWYSO4+vXrhUTVFUBm6C+cZTqFw5tahXVFFtCFY7GmYQkUwAA93veNX0WtoAW
tBCOSPOuuLPVQdRLjimWrJlWl6rLeGc/Ci+UOC+Y+29LlIdUi140kdhonVNHcbvY
jKEXGfb5tpZroc75HMO+BA/RjLYUHi9pdYFwGaMsPaDpIcJ9I1yZuMKG2LNH6UOZ
XcSWL7TTZkWnl6g980IU+pfwgCWD7PpHXqbw4KjJhwnJ8muS4QTcgmOL/rQAOdmR
XI8pGy3CJ+mT/XC6zQbzkz0rvlj8o++YVUgMBMRBBcrJW7i+NHYEGRa8W43Hakrw
KvWoeWgRwozkBLq4P+2luHYvWGR/SHI0M9RWfFqilYed5JFMNN/BSZHaO31k94PT
hquCyyNr0nMzO4dQaVZVHG+gytR3LD4F4KJ8H0NczOIl50cwOBEKful1Y0DqxNsx
HXQBgEmoVckS5Tntb3qGkY3x4shP95GRYkdLS63SoJtp72rcTzLqcX9KosI4XGvU
IsE/xQQYvTohVdAY/ygN+cWKS0SvhrHe5YSVuwXQShZTUdWo2PmcCfnYSjPlzmXn
QJPQgUZT+bcRJ01TAXpUOyJ2oIQv7W7OULyvMa0HmGWHTdL8Wl2pm3Avai0fB2T4
JsMe6mrV7ISw2NkCaVr7cvzMIHxpRSNnrnFDB/xd1ruc96HxjlcAcro6wR535ieJ
ik+8QRaJbXB8hRth3KyokBdjIGdbT7eMqKUfACC6yZn3DLCC9F1kqVI7jNRTrr+s
zBgC8keUVnarFAcr2fNjQKRSNVoUTnRyEXM76amSRamcmqbHCq+Y0hIKeeEKZ8vW
sAkbCK2oqCsQpeRDcXUf34XD1yjGuvr1eL+TG8uin+9CniOCS6XaL/7SYJtvm1Js
u/HvGHC52DjrR5bfR2zbN+LMVEFTa68gXokdnIre7au2+UR26aMM8iD7YSDSxZ3P
f0Na4EGm7XeTHab0K+fao3kyGOhNh+sG3V2IruIQZ1DZKaxyaZ9XAehlDu8YE/kY
FPy1VINiKpw4tzBjB1xO9UsrI3sCGabFt7Sy2D4kwB2P8XutFOEmA1jBRaWclw7I
mGvWW/VBWeAa3f3aZkAlQr1xzrFzMFhOiSwIgABeUxU3NugFRPd8UV0haxocqntD
VIUvrkvRo6xAwyaPKTyB/QNgk9iJ0cwbTtn5BSzuEO7tMMGD+JwWlnIHDZybE+LB
F+jjyb0uIqfP8wp/fSkelK3GlodratY8GOdR6pyUmNRDoSihdq9fPaTaUEkHA1uw
EyC8eIMxiJzQGK1Xjzy/fzFsKutxjkcnfIIlV8TGKqNdlFUW8K0UTMFWpjhx6Gda
E2RLOTS6j1t30zKxcR1/h4u5e4WR7fZaR2iqYyY2hFJ9eCvZ0n3/ClwiMqoWejGR
IMqoDU7QDlndoQ3jcntXxSZtAhRVlY2KK5ZvKLXcPiTCJScSKXe8/OJLGFQ4Bm2s
iey+0l/mPMfE5Vrip1BgO5L1nTuGIBKIcTGnDYj9CzNThqG6ovw7O2jYyuyUNxmC
yPNwZDHe6OjRNRI1SJ/Xe7U+XBzuoAfHIn2blJEsBpb2wIpfP/Vc1Hm6Sj6NOyeA
M69FaVgFntRFShUeAhvkqFAnUtVcGISs8L2upLC083MHERobhRxHqLXF6kmwHYID
3KMWFwO85ClGAZibtDQ1GXLy4S/MYbhxo4xqFg4zuJBuhAUAyKLgLYidZyVcckJb
c3WD8AuExPb2i0J2d310kWWNEES8zlhFPyf/u8CiJh/fpGNuviV6G1aZhdBv+B83
nspU0nDxPBBfk4G/qf19OFnlY8DeGK09z3/FNJGsGTwg4WqlsB44i8VUrZ1rbFTR
KivqBiwGLvIBIyjVXuCBT4FfE8TJN4emCIFyocjBbV80GQsaTXR3l7BvjCoVKHXF
LhVQbMn7bfCP76BnMuj+pOo3LWJSo2VS97C/cQWiMM4FaU0+laEfcZpUSikuu/GC
W8/HXAtciK657oodOKh5fSQ9TcvD1jl6zimMewDnZ1LZEltEoQwOEspxGPPk00xw
RbJwcp1gW7x86qf6niyVM0mgz1ogdLLnbbAPNjABjgW9wYjArzuUGNvtCjkHuSrv
cESQKCzNjF+X9nHBeFzBqiS0QZOPzrzscXildJP5sCXem+B/ZnK9E+84ahbBim9v
TUfuxKat4oQEEby1JWiktSPMcHQdcDHZl0GqzZn8Z3r6i5jT9r/IY7rtz+wmOhrD
4bGemytOIZFi0f7ehwlHZAiFduwKtBq46DEcGgoQMA9j/lL8u38gK6r0JoaDzo3F
AJrBre92XExNFN7VFYk9KFtK3KQvJkl/O8Ev+LxeCT8R8kuDL5DmqtcB5BsDe3PU
2rB4P3soKwqUhYjptOA9z4VB4/2jiBcwHt59DEt1Z/VZBWBfKgmjAyXr9odCDhQF
ckHPOtUHBEWfnq/ryzXC4JljpZ9QfJIq3yPepu4fAWOnkMV8HBXBVw4hX1+a4nM8
ADOE9MDedFC4fNbUasIEBwRDELZujCmgyukhrbXNeWoZ1yrlEIODpeJfNthsifd5
okID4TsSHc81JjzxQUhNJqffhLwk4qJB/yl/J8d72rLoPXbP5yL9s9B8Pfu2nwrp
uD1/AmlBwWAK1y5Jq898c9zyMzDn+B0o4vsH9Nv2HUjZQL2TX12Fd4u8erYB4Ttm
FR5o6/YSAksS0fP0qc5mHdEmnYV5L9Tq/YmSn6VpB3ce49jnYi8y5LIE73PpQXgK
2jo6cWaynOaAIP8U6KJ2rP/x7dgfFVKtYfUHLvzHXrsSCDgnnUoSyrkLNbPtaAIX
vim2ATBzvVavxX99pJAb9OXiFrUBRAPLlJrgssoRCEkXfDV9vj8nd2cOAQYJSMTx
/yMACXdmITClbE7fj5cCmhNVEjZGD82UjSFhT4uNfKUPIhQc3SZoiRse8P9oWF6G
b2p5E5IL2Iarbnlvktb9FVAylmcT6JVbyzPIyHtNM6TWwH4u/jPEoX9L3iOwYErD
wNsoPPV3P/3gieGjEfTs3SO1iDq+zY/QyPu3sbG68yrlgaNsAaVIsN3WwIQX9Thz
lpjDPicXDRNSAlw0dA4jFFd0Zxlyt+9aKWrRrfi69RHAWygIEwRUfZgp8is7zxvE
XprBjlZGSh++HACJDFBMqKRUafeF18+IvnJk2N3HUr1kiv7VZmpA69N9ZbQ+9FhR
im/v82JVapKqEazwEE0pNUi3ge+1SDFc+KwizrqfaV4OrFUl5OZzWsDlzCQU8hMy
Ff/9oe0CXTNtUGk0TP0w8P2rsVOgA/ayxH4259xvzqZcVJ7r0CoXrzxuVsOYHzQL
c/xIt1X6K+FbqezHnjDj/ekZZvY3Cc73IgG++SgTb7ptzeiWE0+C9Qi/h0UKdFgf
R2cT0x+X9tWGZULFg9GyP4lAo0EgHBW8L3qRjTDs4vLjs9TT8lAR6aeVGSMy/s62
3VqBdd747ayWZPD2flSZfzr/CT2OEdd+UiN0qrTX2RsOtheYTiRqhsO/H9lOrPtD
y3ZgEPaovnRz5/DamDpL4LH71oKbdN50Lsa49ts1G6wOVMWMhhbKqF594cQe/oms
C39z+NKQuXuotOU4k8H54ptz3fi+YDup3Nnl9c01Fvk3DA2dVQ+HWIQg+QDaSc4z
1IG0YIbqnkD1tWdFaZJTAetEsgC9e4QMJKeGFhTtToZNArMrp4NXzxckxY7IYW1T
fg+i6qT6aIiTVg9Cql2K35itFzZOiBr7f1KzERYM5WspGAH23RC5UD0Ybch7eFUa
1rxBssyovk1PfTuU1vEeRpt/XsrsUhJZM+hs7O+GgXBpssKXKBGkrsPswlwrsaDG
QBNu5dF0tsP8L/DhcandSEZ3cCCxsaM/K3ZH7uh0AVqzIS6VgxCzWsb77Pu6kcXv
/YeGmvleWFhK6XpTBJxFkntB+OV2W+1QEVDXOje5wU9SyQNGNt0M/l6coKw6gJUE
qPIW5yLLm9XBk97KhQYUbsYaly3ChcO+aeDKCw/5BECUfVqpVl8knuUc6RNP5VYc
ZJwYJ+MGXPCQTUaoosCv2m3pf95eEmPB8UKRRCBIoC/lGNAQSRDmqwhIBIZ1f5T8
TC7kzr8wIOjKKIx6szPpR2bpvx6BXrC3qUhYVnz2rSceZoHQnBru2vuW9fp+pYid
Km3uqNHO+NYMuNuWLdWf7LxYaLaV8N/2O4XL4Ft3CRqX/IHX02z37E0lSMOxM/bb
PySXeX1dY6+qOEd0rvPBfCoMdGnDbtlIgs14E8RmsbOaz3b/Te9M41TmM4u8u7sO
E+Y8qvO61dr1PjHPsdgABJQfyMqdrro6TEBHKxjHiZy8+Kr5DyE5s5XksW8LX/AI
mCv5vwJ1AEdAgRf775UEu9yMh0i9wUFjzUVfrEaxAcI5aoEGNIxBMqZ+yEjkBpQJ
Qk5smx62b4FSCg+BkCpVy5ND2Nv0tR/PNrFizVOfI78sgEsdcf/Iq2mjTTkrgHgm
ZbTFi1vqHpT3KG2rminsFoDOZWW1HNYV/ofehbL2cFcQ5bwcP8DPAwJ1ErCzfDlF
oQwlmc/mM93BWfrau/LxPsCC47JFK7W0H47zPDySLD6fai2XieHlK+dLJ5/p8dqF
9aBlbcujjkHJmN70Nz4Zv1L/D3Edr035mbhevcvPYx9irJP2Tze7CXMek/Neat4I
bcCyVLl16wc+7kQRo9hblkWoBaMkmu45jg6B6oBIek0hBLrLF/wqvHOnt987uVcW
1R64oPDbIxU5goESfKOTC920EAj9lDxOkeTLLm0UzQf2FsjfdQ/7POmpYfq8PdWQ
Xjn82kTCa4gg8SqtDqDuqqVbjz+1D/J+Ceq0dvZqRVGsykV8PDdaD4Uhc4pTXT85
pKhMks5b6VVcT23OMLEVgUUmoilYhPkt4TJ60OnT7nOwJoTGrNyY6N6wjpAQPcgl
/IsBAPpqbSG587aqOyfR8+WmwMvyNa+sNE+ZdJ8+wmlA48/LlE/4wV4FH6BTNcEw
crutoxkTbT4dguLtzFxcXMpxUo/ontyzMSM/ZdUmXr5BkhcDtTrNs2VVmMwi3x/s
rjrFt6CnBoXUz9UqCGY5tFwOOIn1xwI7lyFJRFHRRmXm6WQXdEtVCe+hHfs4qpPJ
6B0eGraheYEwv7XooOmCm9fVrD9T81KARrRP5mgiySi6Cy1xfSRmrFrj8dQG9GJG
6QjxU25/bYnIK3p0chRWNyzoCp7heAzT6fW/LYlZ6faNPTYqFpdDRY49nrdjBTuq
baATV1eb3RDnzsUAWbuldESeqrhJpAB7y9RjB7xfeZnmDAzX3E//k2tw4VI4B9G0
MoIGm+FPMpG/H8hotYad5WZfIu55JCMjIbrynCpufpGA3weY7Yusc42XCZNwn6nw
83LDtQzKlRimVMuLWbUITI2YTCk/JQyM9NGh78RNvHo6i2SxJSE+oAVlOCim56E3
8pfifrXRFLlw2ZMT1kWqoD0wEwwjW7qyDMIYssfZnTpBYBQtLHSsYxVCFRJzu531
t9ek1FH5BoOhE7nf1QYFhcZNTmVh7E3w+rP4cIHui0vMnSf3sBaVFnHgTqPI6KsF
M+w7DZDxk2ll1fTKn7L4pDTO38NLjMzYRcLhy5yr+qL7/KjkWBywI8DYtkKz30Kz
Y1Z+QUBKyFdjuRZE20WcOI/NkA9apja6GMqamPa3+IXkRpi/u21SVsT3y8HlKM9B
xA753HlHjH5STQG4/hD4XTmiZl0FuZ1trEYuxxFBZOOodA2Tz32orMcVuMUjYXNG
vsnDhHfW0TZjkPrwPD5fjcMRCnqXnwm18AmkDkct73Gf21uqPS2G5+1baS0+l4Y+
LNBztLHNNBjvsJ7OJsjpwpPBkQGv0BqLZ/403ZW5qViv2Ua7FiyMxxf0aZ7mypof
1r4r4247XSxEoECiwFbr9P8LDn8N77XCe47RfAq7UjHqVkO+7zPC/eDV2ZYDyxiX
Q9Wy1YKd/r653siZpwqQwtaa7w/eSzjkFlNaETg+MUuZ9yyTk2jp+kIFj/gGndBb
x6IuV5DiJQBE6XAZ7Faar0Syjhvs7DgXabOm2onS7x0l1TyI1wFLjjzo1Eu5gNX2
94BYIgCzM+Lxflvap/MGqJYhr5vFfW+S4ynyIkWQaR/dYCV9FtZRcaPLRP/P6l60
PsTjbzRbKt1tdyPz9ZJ7vZdCUCt/DmqL7mkKwmPiMrlI7JoljgkpYj3BpdtW04Iz
s0YdJCAddA8DMXPbv1Yfp1m8h6XW0U8MO3gKNWn3NPxfcyjuuRB6NIbDWg7QpOPH
jsUFHcwFlktRikAfLUOueP0ALoJzJYaTHbOY3ZnBSrw5xfxOGWWfiGwZ+qDz4eGe
9bhFPnL6ykGgUhLUn85iUYH9cjZZ4wjvEokGMzkhpzwDqAH5I56Hn++Yu/Eja/YF
rdi//zg5wM+a0stGHudGZQUfB08n/Eg6GUQ2l8VWftx+vVCHzXH3QqZrIjrM3UUN
k61VHHl6+arqLvzs4EnEaSkL/0JqBQKjj7QZAF94q5rHkv4KI3wxY3LD+ySyMQlj
sDOrP4wby0SSgHos7Z/JGLjGwBc8jnrP2ZJIJ3C9rMiW21vLm1qEcPsTo2m13MY0
5hEyZMoCgTJvc8OyTlEIqC2aAfuH4qbAXoRQce/dVMY9KWeO0y/GeU4wrX9zzEWy
gSE2ZbIhIzIvUQ7dA7KON32coJ7lN1olkRttapVP7J/afat9j55BnykGVYxbwAD6
g6R17OVDz0WoGqSWSoZIq1zCoswhTE01hNrZkdCJN0fbxyxjtqvO09IEz675Eser
zAxyThYX5IiFp/fHOQJWesFNYYFBvtZZBpCdf9wOI8o1E5+K3p9/YWORjASMxn0H
XOM03pbobR066vKrYvgQNt7TWJ5U276U1xkFtf2L+oxRcQB3qp+lIYVXFwS3jKNw
yEkCPqkiSCMHRkO+XWmDDpHOd2OyeKS7MJASFkM187R4YiHZlZtxio1Y5XcSGpXL
UHM+6n7eIIswSqfnPLzgmhixyllFjvZ7YcAhvXi02MMXv6NrOSu4rlg8ilyWK0kF
s4zCQtqQSQGb+Rel/0CHi9RgB5cF1MUiw78RSms2/xoMwvXomtvY1yS+E4gBKBU2
Vbkqi3WdR3Or6URzmOhflUgxHbEANFMEU4+dN6oBXfpyGym2HzY/Ruz1oaF7Lz4f
85AbParjdG6TVXGxh8FRKfDIEOQo09zuHeKTVH2wZ+L9rvq1CTvB7/0+vpDtydzL
oiUXa5bHkORvOHnsIwWi5xdEm7q8FrpvPpgxGuFyvzk3xES8yaStlHb2om3lH0xA
zXFZOWCL+xc0J9dClRD7jiqk08ADrXiO/+e4F1aKHi6jltXRtgcGYOR/tpdNtCdB
SVKSv0ruguXC2TZJqB48ORQYypqZwF7U2PEylYCgsEq2nbOM0qIBkQsB8ze23vX+
EATlWa6se28y62ScfLIdGMp3NPucyale261o8UpLIJUWFjxtv/6Q7wHlZZDf/zz/
wO/2wZ3NMzc6v8wtS9t1mzSD1aU3kw5gUoVENY7L7djJDcD3vjZLBpzjzlZs6CuB
lL9kk4cGoXb+SNNVedM3rwyrJ9+Re+4OmelvCQdyEZBtHk+co/gqFDeS7jbUUzNu
MUHwtvctETZCstQ26trekkEO5LCxMnkVUjKhMuE8NvP8xbJBOC2Ad59WSi97VEtg
7KycA/fRqRo8zpy403Kv2DW7GMvlyy4aqUUY3ggIo/J2RNMST/aFfBRpLPA3WoXd
S0vGVpNjh/yRwisnt9LrcOG/JUKB80/whgSb7I8ck5D+jPVUxiD7opaSRbxSjkTU
K0dQb6DIEbkEZQdqdulIP/tusAJVHyuzEWLtIX7sjinZ9C0kEx9AssqkEJUXg5//
R89TN51vMe5TLKhRo533nyo3lwhODgYmT0K9JcorglfjDcuKFsHmeFLYlH72qMQ1
TWJRMu67/04kWuL9YPly0dz7TkTgq9Bzl2kw0mw1zGp5ujSd4x4t3ZcnM1PDMMX5
Vy1WC5G/D3DSBEpK56kLTZ/e2+32mbLFfRbMOAtQxDACvhucaUOgeVPgdHGcinkA
hjRtSzUVRwFQIS+MwIX7sW8f25psOHr5FPPuaxgsZ8TYbdJCEe1nyYzhv9UfjIr0
A2kbAjHeV1eBXcIj4vj8wSYkI3EjKnOKGeTZTvFk4Zz4SH3+rDr75vUShKep3pUn
Sx0KZ+elMJAfkSDX+TGwqnRIzxUIQeAXBhdZGlrGkCGi6dRbEzbRK6Fwfi9HLxGj
6COkQCx/3+3cw8gRzngiKtjEax7kP/yS5OKETSvBY/iwpXnodMQrXAkHY0+6psXR
9D+DQJB8jYdfD//BthuKv4xqNxQQT0RiGzPYiDgjhxw2zHR21Q4l14iyvSRWeSF6
7RAoECeL6xgZhVjiG0ndL7wUxm2QouQy8P4hXEtcUWnApbplYj5vMK27GYHc6X3e
iZYt/Q1Vb2q6RzGOrZZLnnMkn20Nvfr9UpsNytRqJXIxc0p5CQqv9eBFQquFqy3u
Ex0+pJ+6URwZX4y1pu4op2P4j00tR1T42cdbeC+MMHgUXVRjF7wPtqIUV6NrRXXs
iIEIIIEmhSofpVCEJBR5rrbqAE+zwHSaEOGIAUOfIcfEhyMu00/MJMYr/RVQ1IIn
h24GfraFPehkTWISmpdlSv9UCNvLL8cw43bUDs4KJ7Hp+kqp8IoiHPPXv+HQrigs
jYpMh1yE25JqIP/31WLcX0Rcf3e/dqCnvJ0X8ZSX0/gaVUNsbZFrNbHQt6MNpA0z
TreUIl/WUte5ZqgUzrNDEAjBR21sFAzIHlSekPitbfUuFdAEHvbBxKQlXZyKch57
KZKjdMSnqPfMZsAVBQVXZiNmYA+uqFb5qo/0o8isuFeWj35BQr7gJw+qYlGlwaRU
kMLFlEcC+DTEs4iOydFqXW7aVvvz2WhzLnuZZyzKf3UAS67Ws+HuQIQToxDEadUQ
zvX9ITFCpf3hHLBphQCQlYVpwy3mBiwdVbLU3YmLYHlbxyB5WINIMiVqEJc3nTWm
6vXThtKALr+182yZpZFMsfVtKvgnjhqs/s4eihhNSdSeD9pWyqvgklrREo25xRjD
Ko4X5QYl/8Kub3zxxL87KJXsdXfhk4aI8H6y85Zy0hjNeRTRxJPv99ro9vSQcrxs
zRX1tANitmW9QuolYbj3k3uAjbZv26SJv9Fj39xBDO4mi78Kj7PzHAN++O1y+mPx
NWhIAeE3JM1PDsQEvx8lx2diJCjYnkEyU2ghZEXH9pmNmz1uYB87eytQwXMqhaEc
TaMLmxxu5fCLOuHlqMDG29IseIgJL4nXyTRqAd39uNtxcow9dwA+F0gS2OdB+YIn
lAAViZiWgiEGA/NR9MgYZJosAsHWgvo2qUXkwaTvyg+7zV/WUrTKVnB5OxX6K/1V
UFqgv5mkfhnk23tyJFFlHWnX+LEsSGE18DgA10tDw4L26cEMQnhr4t5ur2P9uqDi
OHrWE9A6qs8WsJFsYA+JZ+YN3ZzM90/0/OXLxiJrzjF/ETq+X0ULF/tpXitdcodt
IjxkaOHnhaOekIxBI7TIfXOCXoc0KZZwxMXjjnxU+OA+JPIqw8KgW1Htfw8anGcn
Pt2n6t0xiwxsR1jxl/aX4Wa7L4+/gbcUAktmlrxta1u0BApOvZuDvEtFmneDvl4O
5SbrZR/TTreXf0XklC/ceWgiEzj4qx4ztLr8o6raG9hzWVPFhWbcOVsCDHZpSb03
1dUkvsluLDKOMHkdSB6HCuHcmJGJaZ25o6Twrnl4OSqRt3TL+bdKDoKo4SGi+rjZ
b6iUb9jq/4iS16WXTvGTZ8KfDW892uZfQ9EU417Wlirg8/yMjk8KuSiTS0a48Vw9
3/1SNzL/y6pO8PYo9jpiR7Vpf/S4HEBWl9wTJLzD33Pkty7vG77yK+Ed4yzOQER8
lEIL6DV+ETozrLOMr0GVk/dCb1QojjLfgV4o5L4JMtMqMH9kiniv5qaH98yWCeLx
AmNS9dA+vaDTCONaxWYLogUz3axaeMxv7c5TnVgZ/y2nMEyoP78lU1epMe2gG9tW
lsi8vDKV9gFV5jfqC/+0/xA6pofq03mWIeVq9E2SJlLMnGL+J8iWY/rPv1WroKXs
CT4tfQWVIUZ3evGQ9We+8rdadS7aL+vJabxqeafaX14/0IVNwoQWBUdIfM5CwfIl
Z0MLfWtNESQ0m0fmml7QMfY/G/dOGe8FyhavEuvUZNQ5SlhqXplDdzb/kk7GpZzu
uGPZNQJxo33LpbYp5oHXmBj7KFqzdKNdFJc/vm4fN1p0HbxGxeYrgbyulJqrn8nk
mZjS5Yjj8Glx7C3RQTqG3KgrxDt3OWmTfWu3rt1CNq/aYq/6QrQu13CySARXaiWe
nn4dHMUFBc9F6lj2kn6eaVV5wfaCVY/s7Vw/FkO3czXEv6Z0CPX+NYuC1xC4R4bM
B9ixoTzOw3ubTG6CCUx3fYKSRtPc9IUBE3ZfIX8npmWCiCWP5tar3KAa5ekgcr3E
HRPLxey1BzhZiouk/zTqKfEetnxGN4RjPjmSUFPVlYul07a2zLtEsGH5PULRh0Bs
xZ2QdBlnS2DlMy4pGllNvv+xx5fGYwdFGnGoa/zMTDXJt9ZK5F5bytPfSzMDsGt4
NTI5alf371pDW66vY68W1XEAdK7gYj0dwqOMJqdf6Hix6Wfc13d6rno5vdrbDepZ
39kPfrckX4EBFlWu/UGRGtE8oNlTOsYhI85riufiY/eTtaRuizvJ99vhhDabhEJb
fYbrEkkLhbZ7ao5LZcbzvNlUYFouzQXbDsUGZ2w6vL9LWeDNoFRkd12Lnr7zpsm1
kb0oxiUmgRGRgxKpYWZDpCzioblXcGILMALyq55+uB3Wv7grSj7MqUWT/p5adTwo
5XZacCfUhHF45uJ1puUUbluY7g+Md9EZp/h9MImbkoD4UcvsFShesHJVi+i13kc2
Bn7GlbQ+ww3dhKLSIg0GupGUzHq9RmMcDCa4GXuA3cBzfbvPRrAm4vnc383IQ3wN
ZW3TTsQz8klylqqJHNI19VVBT38XRV6d48hfz83y6D2eXqUx5SPHk80fPrmxyxcj
W4PRGiBNQWDcYb0gLdp5axdxVjsl+YNUxBCippHDR9MgfLjZTnaY3buAO79U+sPQ
XgunFhOaanIH4aR/tBf3FMrpVCguAAWwvVRHpzi+yo/PaWNoCa5l9DUkjkMUafh7
GaCoAoeF46TSjh7vGjsrPBC/iJba9o0BC4jMxUkx5J8dW5Clmh3K2X70EAxo3gLU
FXFWs4UkLQvEsRu4/mxjCgmRHUceNit27ZcKHPpEk3EYp/kHjdqEEMZnX88KzwyH
Twfz0hbhO2s9TUrit2Jza42XFwym1XLTYU+047+ZkjwXNI0YtM6obvw0qy+moydx
gfWEyDNXh6DBo/MWDpnyZTi8cNsQM2J6UdaqpCylDjyUPQjzG1U3Bv3i1IVHd/uu
XNdlt1VlnVgIprayvKaI/CH6Cgg7gE5JNpmr6Esf9YEPvir/E4lSZvYNlU+AKyZO
lDrAWoZWO2YjMgzdtPeXrO5axu2G0+XUat33QEqVuUBFBxmu7gOeIO63w+ijwP72
YJ8lKhWxAmir395fmHxmWkIG8aQgVyjuMOAoOBDJdD8A7GU+dqMrf8HDSNIGhG4i
mSMPqH1A+y95WtVHygNnqAWAtA6D6xsUn68em+e1qxG+7Y6l0U4x4D4Ymc6FY4tH
xMMx0Cf4RInOzTxQOHoaumDwnmItXiidCXnm6L79iqyYMYYeI072qLM4Tm8Vs5T6
XF1YvucAKxdmIJJbQFe4M0LhV2tMDwx+iB/eXJmtrT6ZLJJKjrWRZiZp90YrZYvH
4pofuVaekSQlg1DV7IZME0iuPD5cv+fQS4l05zf0uSqTfuaE2CNZV6nQAlklPCSO
d+LHeY9r0zzI2acoJWrMKj3zab56uSbtW71SeIKL7twEECU4VR3Z/SyAXbDVMV4b
K49OsHXiRXtyMnx9p9/WdUYhf6lwA3GEoY56+UatcWIjwraRuNku4Mg9nsoO/QmA
uDvatUkpZx1uHpaz3NHmdgLzNpjDHtPAQKgASNo+ajebiJEn6dzq1Z12Oo+036PK
cCmfJHUF2Wqj5GGENF+dxhr46sWHoCo1UjM13WoC1yEA0PAydWxLmkDBwxd9xenn
QzjJfwF2KzZshKE2Q0lXL7jqSW/eTOPg50CG8qa/wCT9k9P84A4kjTHT7o3FN0ch
kLHTcLWv0/oCIQocggnRxQtZ9/JIQna+Q25cObEtMKGeCv2gJ/SUuqbDSMdzmeIa
ZxoYsdQUm1UWH7WCO8bevc2W8itRDo6m8HLcHKaxp41K5FVeP5PCrxEbxADhaLq4
8Zw1SuDnEl62TUV2EaE8usd02EDY1tP09qLB6dm/7olq4FVAMtGrNYZCn4OHJBb1
7FLe+pLHdVx+m2dAgqAPj0KCvGCtIBbe87v3oprha4ivQS2IybzLAcvQz8pYIOTB
rgb/hci4cPMPYnMtwH8tWMQ6KoBkE9Z0EzGBk2TfddfmlrYF8vXW6OPCXYicWPoF
4jJS+aZ6VOW4CMsnnRNTbnSWjqh5J6O6ESeVKi16djWezwf/n2xPM+qDYqsfdHe4
EfNR333RsoxTwk+5Jm18uG36ZvvhGvqL/V8HcJr3MHNQYKl05KFUDB5k0lOK1R7s
AwajysENCDH54prcxFa6cLQzvn+bUBrCSihv36q3yq1gAxOoDRaY/+BnyyhQHrsY
8vt2fomIojR2soGVeKzRR1usro7EBrL48TMb38kHWbPZMvfT0T3R3itv2qhVNRS+
f7+uqLTdLWZy5/mBgIjAczpvB5LhCuBYivjT6lCioToQZiOiB2fv+3xk2UPqpz9S
TtGYEIJfw/1j8xDWb7SUcTp+wVKf30DDEW7DHPwIy4OVN+kytkHumAN6mWKcRa0R
/yMYePOKeBwnYqLFHrXJYBNMDAzfFqsxb5yVHg39yw+2epG0HCNPf01efltserGr
YyUOFEBhtcbjgzcOKg74gqHWwkjecPG1Y19e+I8dtqqqIKsr9tZ0X5m/I/vDwZSc
ggODDHO1TwpVQ1fmRgl4KJuVcMLeyi+O8+1Sioe176Wm+RKslsw5kUi2Lbwogho9
a0aOA6glrOUQNsU0iobihL9TZ7UlgTH1Rv4KXl6u2Jd485rhYdDxMcnfgG+chu+w
gxCpziTx3TOEJmnoxTbKmlXTfZWUyW3q5Boi81ejbgW7MGoE6Kd3/sAXuPSsypRB
HrkOadjBWWlB3Yub7vvtUzHZzMwGlNVcbpzn3oaE1YCClobSEsnE0h4Zva533Bmk
+WJtZqdrXHDLM68rP7hOC7qoYcYswv3GgTAVOl2BtWN8TR9S/PHw7hV4h0iky8DT
MZ9oJ4yU7mwXurRWPFz6VGfdoF2oeqPx/pbq1iDZz1xF9wdsfXuJoXOCr9VzPa9U
X/WvgXc0owClif/J6o07Cy10OJTszYCuqcq29IUVf0VHTSKAWrWRsvbG7qDPAvfQ
N11hXHbLTeO0WJkrSjMPHPttOrO8DpSBDyKOGlD2qeE5qTi1Bq5l4CwyHi7ZNQOO
OXwrqwP19CaskdEaLK5W4mDK+hGFykZcV7/L0M3KrRp7bzMbMOm8T0PA1UxAgCJd
7oLG8MjhE9S09qPeJOi0LGrQ5YOO1c/v/3yXsP1YvORg6sW5Vp++AsN+H5xjY8kk
JlScqAD9dd+ASHTP6HQGKTjnjZD/axYavrJRmlDM0E6+I2uYidGWSKu4u+R/EIIm
xBpzq+YqlZbLBjMLceQHgMU0wygQ/VskXabQzVg7I3mU7YJeMsEkbQilys2BR4gr
arfXXPCeP16i/byhcU4Oa4Wup8WbAfusXZ5bcnOLPS8ioCvlECaEV6Jxb7I6nChI
Ns1Uxja1MPRLYWd3GB99JDjJg3C1OXPQ4k138CYCwbtvYeK+MgrA/150jNSxscOF
97kw5oERgAy8Gkjv8jkKw46NvRMgVteHkb2IaMpVGiQzn5fUYtEf7xMcoiwFvtmX
Csf6ZsTXca5bv2RpqFT8m9boIEdWHm4NyJoDCDYxUJ5O1u7JD86HRtyeyum1znN2
7HGGThPW/vhn/K8WEWPKgOwvQIRVeL+AAQg1COMteENoiXY0sG42t4YFiecZQy7k
JVckXgB0yvNwXO1WiGPWn0I7QBf/tI6gqB95uUVz1wjcYVskZSuEuO7ddaYH8ndy
9h8WSobxIaOyxyG+zmFOHVIvpKGhM3ZczjOeotxmK5ohhoWTSK4zK7cZjuxhDQxp
dRSsxegRlwIu1A2YdLOq6w0gG0ueElpj/+nPbAskO+fNRF+yf7WDxgFvmqehno8c
Q6GoXgeHX6HuqbLDBqL+oT4AsA3QHKgQn3uHGC5gaojvin2ywZMqEbmNBcgRvHM7
nnh42jmforDpGhYbcdTI90Wn2+kPx8Ck5pFqe1NyP6YSAgEYMKOaO68+CeSuMzBM
emCUVjvubwvnDkvb355pkVUB2wp/WZWz0MMlFg/oTmONlXS3bGMzF4liTeNsttgf
5vW7Cczx+GuqRSkHkOTgvoc9gzVozalYhH9p9n1bT50TRPDvsv+R5jw6OqDymIyp
JbHfae1cV2YVSsbRrryGu4V7ZCnfSfk/pUs2zMLwj4AFT5ovhTGiX5u6+3lujipo
cgFwbh+yaeMOjcKrPUFE6QiqWEuTUoGwZbBmrzHBOBB08Hu/OTAq7oTE90jAFF02
9Nb54yT55cEVi4tUbytFLJULiAMy+PE+ba9o7oImy+Sb5uKdrVDrdvGecQDvWU0D
gejgMpu7/Qd88jJU6TBq3iM6+1QCYObYXnvWjJqXdsF6b+f+9vinSJPwGHqDV/NR
txKEvpURc+0L+eQj7qxXjTF8DaDxMT1Km8DYp4T9ZcS9fAUm3o9CBmg8BpR0KJbJ
7LGF3H4iUmsba12oTQicWXtEaJUl+qMybqCod9C5uotLlj1oJOojNDJ99BEWJape
IOp2zVxlVtkQRtiCtADbJrvd7eNbHKpgy0dYPp2h9fUGwcU/JVMnQj0nSSa2YkLx
nn86iUc/MNmQLxqSxzHmKyZmkRsVhzYaSOHTrXaWbPyI1PATZSM7mg5eDAgarPo6
voMjsvfZuD3NHYZ4iwqh2q5SGnwmBacGBXGxnxTwW2wvn/paL1Ve0UJE3plZdL0I
2j+plK7BmODNgcinTIqHtQoNObkpvm0u/3ZtZRq51XHHXTJ58ftQFA9PHhC2/nIS
i/7943u7tVKSaTd9T5Wz+2f6NZbUOusy23enVni7vVwh6Fu8HBhRjjQPMMZY9c6k
ThVW5toWfsFzwKBWlBHL+KunzG81je+glYjuwTcMs247ddUETLLZ4+i8pMWnfpcf
oFFywWr9iGm36+jrT59S7dkQhtUplC9Bg81QaFePnzvxgn07nGvB4UvkUjqS+PQC
h+6yBPlNB9svWu5eMTtj9UUtxnemHwR1hKyAk0Hrq5TV2Si/uT2FTLmGrWhAtIrQ
5vjk62Ya4XtlFnETqfD5s4l5YleDAxVf41DhRdt3uJ8lMrzO8rFs1ab3jrx7x/le
XxemLtWsjIgDcwCA8FeZ6zAEW9RXY6fzSHz3xGRJM3i/oQg3XLffFnwQYXbeJEbV
W2uaWkPbJM622lkP1cTqf/BnU5wgFynzRbFoTLaqQ8ll8b5rNg3bXpUW9rHxKqZD
fO4BFxvNi663ty0Iqg/bMuNXzvZOrlwyK/Z3z4ORJZa52yq2dLxsteSt7Om7nSHH
TgabCAX9EOzXIB/CWNs2TNT9RnZc9tMGzX+foAqDPG6JEGQW34anuC/iRw1dhloX
/ZjIy9fc0pm3yY0MYMskQks1YezytpcvKgkePQzc2EA8HCPHnTzk32aY77nYxT75
+iZQUfasusmHlbpXnsgq4OcIkS22RA2ugbryGfvHiIlqkmcYUkRujRLsNQ7ZGqSh
wmLusZ6YgOHw0e7qWFUkWuZKPYwRRMKhSpLi63PaOVlnJPfpGZg4QuSMg36tnUxb
RoIFtUTh/gzK27h/p98b0D3q80Xk04crXeb5fZKRlF7miAwPPPONLw2Z1r6/xTeo
KcGi+Y+s0bzpTkcRmreBIdUe38byODtQkItmO9creJAAA8X9ZRAQBqRxZcDkhNm+
ZsJBy2+Kk9VsnVCH/0vdAF+ZmmS16Sp8BhJmQvNL7aPp05TRVr9GdWbAfd1TX8kg
H2e+/Ca20S4LYqnIONlibymUj3hzDnFfPW8mKGj88yI8ovywsAjd1PJl1f/sI/KO
SedFPTlm43+Pl+JB/F+caaAXkyQVSiCLsLobRcS2qukxNzsm5RRUM18XWWSvO0SQ
A5yGay4KXBbmwQnLqBbuz858bSmgx17S3aJ1PeYiqWM5ZVvVcblT/KFDJeEpoZhB
LzWqiHd2JVcB3dzJMMhZhUuiXrCQ0nwEvxaLzYCrTGWKFZzJwqYJSVUfUfB/jSyi
sUAhgHP2Knq9v/Bp3Ge8bV45Egj4NQX8HRi7Qiv6baWizGYTgjrhGvJjVYCgvRIS
2M2y1IDoDxtCARgEMjub0/FCjYvc1B/n6cK9RJXZXlZLlp54yz0EyCUKXhrdFutq
K0pLCibM1mfM6jj+MV1Iq9WioecZzefKWjXaPGpOQ8+kZ48eIrGW2uYXrIM8oFyA
oxiP4ZcM+j55/EWz9xyiMV7upU6j/SpGeJjsXIQ4rdXxrmYDRmujXBsb8kqBV52v
TXIw/BHv5rOxdXl4Fo7nndPhslIuywqp5yVewfwE3DzyBbQL37ci8h3rWbbYiSRN
mRLDBuDDW00+1m8DaRFlUFTd3j5qiqKTBSw2tnSgMH4mbNyb2pAoEwF9coVxcyTF
Vmhd2dm2WhwmCNZUwj8GZhC/MzgcMK/vgYKQJpKX5cYIsMpkk7ciKAUis7KaHaiP
e6iEXqugma/nUmSX4qZrfevwXF4Pjha47THUPHyD4VF9kQS5b+AlzK7p2m1BtaZo
vONnhMY1T9XOdYJsGitUyLD8ZrhYsbDkKfeUfVRPErE5l/Mht8BeY4+KbXjmqfNH
Dc8V84jyxUFzCAy0txbBiGT/K0Tx+wh/IvnZIvNOIi6Loth4yTa4bkAnfVnaqSY6
ZDmXgee85FWZX4tVEG5pKO56cFAgDrMeRe8/bkqe0eBSim83eMQvcBeJP7Yuv1m9
sMuHnZNyg4+i2i5XVsp9uIWwKUkqo5PvRpNNjTn84OWpu+5PD0yMPlFGJ96mQVqE
wEKvxqCuB2upi9sN0z1y+QA7tIHSEhsBC4kqGieGzFt5S8zvNbMjUsDW9xm0nBH+
Yq9mWnXAta/kX6hzr/gzt/4aRLP0HfEvNWRpfv8CdXsOVkDw2lOjEVDcL4M4mPVU
IWJAjRDUuewSifxb0lsSgycYkXk1GzRev8sPQfNvAdEw/FOpX/MQ1cads8lPf9wE
gzPf69o6nX42zpbL7MewN5QTMPslgMFnm2tzhIQ4b9bMbuwzVc2xymBPuuKbz7th
Yz2dwAmks8LJRuYMDyRAHw45S9BTWS94mjiXBl5PAAZ1A4/1NVugdTFFx6fH2fqC
KTTuLiBna7y3k2f8xmEMc3QKSSgw/W6YyzFRTsMR5GobinppLPrz8iHyAGWJccyd
bKBWpcrnxyuWAjOvSWCybxSppaRVsxTUn7p35riq/CRJtBZ7VDs5p52RvSOYjfI3
rciFKm89EVBlBTYtWb3LrkKUOa0fiGzHML/1hHxEGYEjnV1Qb9YCthwzYkBMasob
KCde+S3pTMw3+D5Vxn18BahlOz80sH/3SkmpA+rIXnnh6kUPsaOB7VjUBynXGVSS
B/tm8SaUNpTv3PwyMFLhdNhKkkmbt5HvyY1t00iyHxSxm5A4V+16F2KFMezs2e2J
74VqnSR4fPvzthAgzXAgQikcVNPEVJ9axQ0O8IZkVqZLnDCuDaFVXof0jwjuDfPa
0oDKebL6zieK6P04jK7puGbFZ/mTJrbQjXTKOgQvqGeiuvAEG4khqBMMyNTYCGRk
uyJIlvUkjIeB103BXKw9EjxMePyt/7jo09fPM2pVteyvrWZFC1LMjNnqGjTniyWE
ZRNX1aag2mbWAL+1TROwz6vdMOFBjHWPFcowRRo6JND818dlUnK5EtkNvYZA7YLr
D1S9inf8ehHYT88eR7MV1p8I8Q9v1F1B4dVA6owCutxXCHOLunpO8Pv14qTF6GAu
CPJ6FFSKhVHmRUSOH0AvLLiwyTw+vBEp5V7Y1vNQ4SEAyu4sldzapVKLz9ZkKrqy
OtKtG3EpvAB5WwbpIqz0AfY3aCWLd5V9CZ1yPMjdxgCXcqoY1glDcZvaZiK49O8p
kPnMyM8m3cwHp+EZ2GwmUYagLFVTiSIKVCH5i7qpVKiFauW47B6iNM3Xo0tUrFyI
bDpxCMkn6JlrdlQr1YBHCW4hj5J+d0T0MQX9sNOxwSz1XkOZw37Q1dghyAsLDYvA
z/XlGKSpcOwyZ3F/N1OURWOLzFkpOdRreDh9vkhFbPIT2CVXMZshxKSJlbNczQoz
yIhkeNdDihVUaNP+ks/uY4NP89LwGC0kvCRZshKcg9+yshcbhpVThIA1VbeQwo9M
27EhULRoupXAoXTesZvoY+vJE8+99eyHkP4ouCUcARVkutduTfJBEdTRNE/gQIst
NpGq+5WkHuGXs5TL4AJydtm2glKtMyUKJKIXVjZnIbUuhbEyqB/Y91Q30dpjf9U/
7TZmzL8WpcHE2T5sgIcsGMS2ifOEuC0MgPQF2+BIfFRdphxc3+/BHGtu31G9Ih1R
R8B/uc6Hdsbgmb85qoj8PuBPuujYvlIc4SN+JoJboh/vFUhxNMAmeZbDmGhetHF7
KpA7XDeG2IQ30Ql8dNHMMX9Dy2UVLTfQCRhOkJhqTTlz7x/Y8n9Fd1XZJn8L4J/V
iSLLWaVq+4j6EJ7J4xdzdRFHBHD6xf/YjYVrlmA644N8soeuSvy9IVtvrLR3Jlpz
yZcQjDYFoFoH9lSInl9+324TGsVw+1DMqmn1WnDHi3RdZGa2Em/5nA0AXcSiNnlv
Yug9vTQYT6ngM+VRd5ri+SkIQyBtP9qJA0nAFrBc71GhwJ2h6cV5RpMDncZ9MUW7
8wJBEdDDqp+iWee6aZaS4YmGkLfoD0LcpetYK/nCXa5kF6kEYGst+1dkI73UQOmP
4ItkhqbolfqE0S0scagZP2hR1MbKhGaNopwXjmF75o+udvI9MCc2t/+whAeL/tKo
c9S/kSA1xkF4dTLbX9QVwwPn57F7TXvqlYHpOMtlie+5orsRBAuL7grQv0TEcFZG
nM1iW+TjtF064yAWfxD2sFZD6jp41tCaC91jTGe15l3HU8GCAJaHdWGyoXzEvkdf
fxwBQBShve61z4XbFHsdD6mZynU4xpUXAAJT4Jw7p5DbihUnVAVe1+GMPhuQ8HbV
WGsn2JuUvmSikw+juIR255xcLS8GkG3d3J+hGxb535xnVH0tmcU/IuYcSYg4TR3/
X51iIED/UWymjZyG0BYCdEqLGrpw9laVd1dUApHa1CpeVmcpY4DApaomX1mUVfca
+jigQfqud5mgVbtaXhndyvYOSBEAe/buYZ2TTwwgCwIh5kFUsTWWu1V4mZF+wHdd
rAGEcMkMaUHuwgkAaAUhtkN7PPMDdvCdfnzQEoLwbpJwJ+sVsNmCUP4t9ZcJnaUi
RQRGOhP9TypCFq855Ccw5x+f33SCwxdEet5haBLtKmdSSTpiL+3ybAI3wqVKdXjX
i8ItqAJSqRq/lUQK+SU234+g3qxBoTyw4QaK6tIipTuZieaHx+dmfyCYwd+u2yge
ZiX8FOGJztoSKyAiNsOp1IpO523w9WC8FjLpkLkFtLz8hrd99iViaHJKGMc5oNsi
9zv86w8IQ7uQVVaOvdML8H/6ODJ5L3Z+akZk+ujNRF/xMqEGEcjHYvT3+Xw4jwVF
BqScNH0RT5X6uxnONuBY9ZZyuAy03BDJ6KaMrLSCgXikNZAZb/F8jAKdEDtDB6Y/
F06LO+0JMFsEsyxkb+9aSRrd4ALUhCZ2svyaeYkaWGf3+K2Uq+nnCBHpvXpuzAdm
3lCpXNr0iURXjdKA/5YViXwOlBdpJTm6GeGj+m6jJiRYSxE1UsoTRCuMIqJDKVNB
ZYjkYa1r1OBbEv9RWjHl/FtTf1jeBN6xCrl74MOxoZ+fT2vhua/OV4fpNKhZNBfn
V2R5Sw2a/lfJywjtHd9eAwsQ5hlE/g4l8oyFgYp3HFqhAGXdI+bXa8H/lOwtpFEf
pYp4bEEZ5VtsiCmor1Y5y9xEsYGLKV3LX2xUG5yqmHGNfGf98bBBhUndu9z/iJxY
LvOFK5UNHHwgfhMJUhCiL9Lv9bJNUksjgJeME8gCSas7OXZI1vmb/48Td7jYRabw
nx3trTDI2WJQK2CFCtOgzeoG3UrtDZQUpiM/XV/Fwg5MBehK8iX3BlczjcppP6M3
31rFIxd1f6WSh74Oi+QXI+u6OzmsJWShkK5Ben9Fp3RRMLwIJB1vtHFMoHYeue6V
LD3N4s4KFyo003YBUvQnbtvVWOKLlfpDiGMXjrmBkqTAj0ZBXFTh9adhV0bfG3cV
qc73FuPdtoyvKAli+y9XPFjFgUpQ9FNljfrTB3vKXnUpwqMRcVotmpub6I9iKoPZ
1BKcwhLBVDxj/vW69M6gESHKwluQ2qtUlpVi1h0XqVtbzeLA3mYGJkIiKEB+3tSP
4jBxFJocbfx9N2RtuC40+erzNiyo8Eub9NcGjkTHxwnt/+8U+GcI8RWGQUjo36GK
7mxUACawYzkRMfSBHFE0EJwE2Yucde8QC4ojiLSfiDftUtO+oCkH3smoSUm0ouO8
o66qVoRoWHiLl+nntCJ8I1kl7C/LFvC2n1SmGTc4VqCDepnHVEPNJixJSMdmcEU6
wmR51zbwGGeaOWd9xB5348QQs7j2reJn1X2Qkm/GF4/g2nsOMWGcc6/xf4tGsNNb
GimAKJU9bpH/Uy8KeL1/E7RJJgnT0SNl158+fwduZoEBmpEQUzjhPr0LBjAQYozM
QEsxH41bBdGBQ7ZnGlo8G7T63oRYxHQITemJM2bOrNeGWrqWuEJg5OxR5qgZXN4K
M5epwjzxSWOebRn8P7o1eqXM1TFZe3TrwU39nhRZlNu2935yYWeTmhKQN0JHzAil
WnznIdzNCuGrAxL2YixPABrI4nYXHBD/164ohtrXB95C84w47KpKsSoNwH2+1U5O
NkOocqhA4GvnYW3zEjEY7Vcrg9KBMUR0pA/wUzhNi+hYquJ4uz1exfrW6Apg6BWZ
isPGFSXK3f27HDg37jBB9ScDGsZnHAUW+MyY6J/8waTUxjxAYydvnJwXtD/vVXfP
gkhKEOL5D1Gg/xYLEQ0s6GOfKicd1GBqOBQrlieR25OfKQWX6fa+Cwlibf2GbV0c
qn5f6I9O1Di0I54Ag6pSDZbTBGTgKeBD5DcZrz7wZDITcA9yuDVTFtS+UPwdyXir
bolOs4gHUv9aewMvNRr5s/QrsE5EM6V7w0i96JduYYY+msXgYlyiecmTfFFPs26C
BFGhTKBQ6Hbf9S4RIUBad1g7PkGPspH6RAubNByVXEWr9xyyd/kmNFB0sOOVbDPl
CmPZWVXYFjgJTJSBRniaBfhdbq3hHPAEEo+wLHsfveIds7GN0RGiRW0LVrbbDEcN
YzA+cUlB4l9d8uz4xaB5Q1YOLbfROZIADh5LupxPL1HO4JI/WvnOmBsH2z8LqhGk
C/6Np83esF31pE9mmspF3EUi9RU9MOX6d/tolnonfL9TGJlDGgTi8CelyIj/SWrv
i7fdLhKC3oGJLHXHkN4gewlB95l3oYttfsARdG2sg/jbWChJDV9esGq7k3Q+Y3YC
5ULFfd6Tyxn4qQdf0diAgAdahUFsEBPzcOlLwiS0iQcfEnSS8UXEMY4Y/omC0BV3
8EAyh8fMOuZMXEEEZON6pDD4QU9EbiTJp2aHOp49OxoDHrNAOL0drE8N7KXCaKCu
vFi7qZXJlJV6JxA05D7PyGetZaP0u6aPpF2PuXBOJStCoYDkSr8Wi20ukmyszADU
Sszs2Q0NDrFmwBBd+RHHkvFY8sw3Pkf1isiIUY06N3OpKvIyvAafVdWXCPhs+ywK
iPFIDXkqJeuf1UEgEETa+v4XOz7Cyx6xyrM45rHkCCNKt/AJSTkJIVPsf2niW15v
1dk9HJB1Z2m1kf6wFxVjm/vNJrlMJ4DPv2UDsoiANUxCpbEwjEH9Plg3LaBOUHzi
2xTbPkcCGK/LyWh2A1O1FqmhD/UVxtDBmc/EPsfHKPDLwNmh7+PzfcgTLkm/mzKp
+DI/H4zn2MSa5oGGh1mqqjVERHTDXmXD70/f4nQtkHnPKMq6A/6g+jHkT+MnG9VA
ikZoeOc0q18GJ09BHhbh84kAZdUDUGDp+mCUjLSBDh3JHScOuOFb2Y1X3ywVSD6R
mUoeBloRMuXKBaIvt2OG/0kGVlJkFHNurEzorhp26lAeWYxx0Z5zaVxVjfBhM9w8
zEHZGR/2uqTvyAYUBBv/99mSodx1MyRxy12CRFiZaVnNTYqTwo4V+A2ntsjM43DK
4MnhkUDxJjYbGygeuyOhwXDGdQT++L/urgRJodCE1xvBcyg2EoDzDjvRdPSy8/+2
UgG301nWsWYy5A5t2bN7pjsEyiRRYqU9fRlhxYGr2zwljvaJR5K0v2OGOZXuBJd9
xZV+gp7Z+uocwHZlBgv0dJhJN4YFVGXHthtbkwye60eyiUz/Oo8cUYKt4nZrr1DT
21vF+xePD8mHy1SI0PZoF5Ruq0WTxduwsBf6Kr5jzjkLavDNovLHX2Co4JZsE+Ry
KSLEVevbfzzgdHc80DKEZfZ/wjHLKO/Mp6LbhjcpQpgO18y4mMRDSKDQ85zZmW0x
Kq/8a0jRGQ1W+BdVKg3fdQp4IeqQmzl5eDLuMOBv0Gs7clQLlmFe87RIZXNq7nme
ggb7o0YoHS1nRoIDuDfv8lN5vjlqYM2I3PJNN9qBtoVtR1lh9nvMQ5qfgFVmcvpW
7wqYBzJfRXyjVgsNgk2iaWGhuAko7yxXxB4B8l/oWa8QYerzLpF24cB0jiNwIefl
qrBKz6idl0R5j8m3avBZyhO2mFtAMBvGj42TKnNK+iWk3LyXMbbTonO591sJ7ru1
qqDkOhcBd4zy65l1cD6Z2Xl6ZPr6VmiG4zYFsDWwedQ/7UOrfMddkL4p9ETeCh/m
foqjSu2CdgtNkmYanWiadls6FlP/aroIosV2yVNyFafdFiWHkkirIpfIgLZKTKQJ
FPuLySJ8B+UnbGdWhpbNeV6S7fw+E4i3qV1Tcm0H9ZOW+DuYB/JErnPVEbPswHht
iMzNJzMriI0umIp0VaVRMFrBjfTv7XXyxbIyIXZdPuZX9xfc+IAMf1QEa7IvaT2l
QnRdSQD0Z/F6khzbPgxTH1D+PKQBMOWI18B/6hdZXIl4yr0rbhJIEbd/sMoj+QCP
/sI0gbb8CbYBLfg8GvNFKiJmKobIYiFzsbBQlnB100C1BbD6Bgzb1u2QVVz5HhCE
FQSKiDHlSFG7kdIX/L+7hhRN1PkP2/QvImxDbw9SOj/W8Bha1h9OEqkHq2UAPaJf
sCN2l+T62kpoWrsL6IEwhQz9mn0F3Ti/KzI4GL3zJ2jO7yt9QIl8q1VxzJJMA0N/
pO+fvQQprWQPlJnnFO0tQKYItoGsTA+Kl0AIlwv1vWXCzdJVlesLEQUyh5caxLoc
w9GMF9sWG8Vcr5d/bsfjGYEalsandh60+W957CeLr9253RCJd8nF6fsB2Jk66+2C
CMqH/X3t2c9LDlJDGXHotUuh7t6AkFNyLTxelEpOrVcvBSIlCrKKAPLPFdKHJ2xh
hDXJdwycNb37sesQZCXz78QwhQVlQv4bgXL0/sKgZtwB6YJhDilGm72kpYnyvZy2
LRcQD58R3c+MUy1AcOqugjjWALWwtbgOGCfhxuc2dsiw/8U705oThv6PKMoTz+IR
l1buOs5/5ieu2KclrhsPSFhitKDarv6aw9U2HF9109TTWc922VNeIM+b7aJWRGb2
rxZRDWcH4NLueZzBpHzKsYg5nkFTXJun/OtoWYmJbpvyONo2bdOa6G9QQLXYTw1A
g9CZFXgj6MY+iBQzCsn1g4h+aq2Hb+7gJKZPAd4fH82w0erK7Ty0D3b8jM/RWALs
Y+Aaxg5EMl6hXKfgaVLCRRl+SqLAEYOPksFwAdYoDSf3F/NlM1W3ZQWEMsChHJBJ
knokgE/doc0kQleHfYolzilW6UE7tm98KgIgjvftgWvF9ynApVHzR2FTwmgsu4je
Lp/8gja29rs782MSYoJTLJ9uTHVmVff0k6k4PY+gk94L2sn22t/CNp4SRdPGIS3B
i17XGgYm1JsbkL1gbweQMizHbz3PQXkI8n5p8RSdJ04PxtHxQkHTu4W9GSA9hfP1
ufOZBticok8vTz0fHVOqFm+9IKBev4FAx84eqe12XmWLms/6Q2waU8MRld1eKoBy
YRgkRafqphdT+5x+ShBRis+hTDk4spVJkx74X9cLuJURVw4PITFapusp/ovDOXQL
CiDJB+u3J0Y8AbqYkCzq5jNlV32Q3S4yMwnfKkzDDMOnq2nJrrWkscWfshJhwBoU
fjW4GtglBLDBS8ONHPhTNlPBbz4oOQakhi6KX8aK/EljOEq9Vl9B+mCgN3Qr1hSa
4L6roXY1481e5zwhR3b17eIxnEcbCCmMtgK0A0CpkzTSQoyOxRqMr9IQ8r+5kaoF
O1tlHoWDcwUOecxZFCDbqwAViCIbTeSFI0cKiT8E81oHiX59b0WhZRI775Dj2CXT
GJdI4P5S0C32yE4sPk8zFiZDxlayOzUzQoqOrJN2zRCe2zL2/BIOBTMY/HwrwokA
kICEk8sIF3ABgRupnheFQI+8mnfWmI1ZCaNX+bi60JSpIvMoSlRc1J+lIdbLuI8K
80pwUzFbY4gj8besKToRvucUYyLPJu9isK1zy2HbzhdBVv0D7+9TTxya46Pnl/hA
n57vNa3gcrk0AGfNDjx6GvxIQdWE6FfgUoSnVblQxh2wCEa7HpKyt80tCoupmNjm
gUUw8NrXwT3gvcXnA9L61QYFKL+TdQJZLuiMetJys0EMRxLxASpwGtI2QW7Pyr5q
v5olUzDgXRwKlan8DLOyretK33Jve1i6hzo8JfnJRrwWCT7HXHHzoFLePsTChLu+
bUtaM9EgpcBKZ1zibLQYwhPvzdySOzTceTyfkrdK58bB6Sxpou3+OeLZhNWnTdaL
1BZqsVmwxwdSxMQm6/a+Sx5ivuU/Bt3gz8CwoKcMZdcIQTz/Ej8CvP/+2VwGMnmv
RZMe61e5HdIfWILy5AcMjpmALfGR9KIR1+BNFr1kvJtfXEdzH5FQv+tUvS0Y967n
Pu9DkB2bmfDHiD6WStfBCGzf7g5TyTOkNR5XarVZHV416AyslunaOF3YKL8Fkbfn
H9scrPbQPZxfWNMHliNQalPsYMd7sEVtGIDSaLI4K1Hf/3K3lGkhYfDFNO/YZgLu
Xy68t9HUZtFtiuoPxyjk4AkapHHVYp3ZIw3xhn/C6/dwKG4d6mFlIxTIUKZOdUqi
TZ8Z6eDUUOYwCrYNRtxXcC+tUFHe5EoL1KdEBszOuuxMrK1em5AnFyupfLyjhHL2
PhLYprU0QR63JwtY1gSOiUmBndX0cC1ORsxssdPHfklZ0dDJrTppmyDxGBskODbm
OO/huCnWZIlEKEEgUoNqWEQLoEOjIv/3bXxgB03fD6T709AA8st5D8Oz1HPWhFC/
IFIVWtjAd68Q0MKIFqSjvNFcMuMnCujn+XfHiUOX9//CmolEI0AsKDJi/5fp9/BL
PVInEQDsbB0N2H6AK9uRgq6uhjITsYJwga/o/9z+Goolk5wLct704/Q1UBeEMjOd
4dEUqZpjgFCsY8pyHvyGMTRtF7KyFIS691tlrZP2Hnge1V7XCAyfSabv7fBmwBnC
5JVfK8XQefazSYKDWm+KvYshtylpwRMpFl6Djh7P09kW845KrEKmr+Y+uO3+J4SA
Dc8IMByW7UjVI6p0FkuckEYh5gfs+RfPW9EiURSuspq8rp4HNBl29XUBRzKU6PP7
k2qh8UH1qEHznueNOSXLKsB30NijgURMZJ3uft9Kc6Aq2GKOtn7ve4S3zzmKbz9g
LqF1BzpRID+IN2ayoYNwa/IstbE2+sgtw37CnJ6y4VxF3/WwJ5yg1eTRP9Cm2sZL
QU6/Bq5gwyRZRW0wJKit61tUWDjo+bq2bxB3LdkcPP2DcACLWTpuIKr44+Fu3Z7d
2WSHD0vGMoplqcUiBivC4UDiMDFQZ7mpLRy+oS+TjtllQ9CGOF84M6Hw/5XTy1Qv
TKiLXPZchEeQfdmCqcNTkMsXBOFPffIqMmEGtGDtgdk0t3LExaUS/IBJ97m7XxpK
+vj4zG4cUHiJwELe3LMfzXEtE6y2wfxFpWMIynpjFjtj2oG9yDY47BxprJokwUxC
f0zfRjmeyJQUlrGqBO89h40HqVMcL3x91iiF+DMcpZeLTV81EJjdTRA5wM4u3psY
vXh4DWWa0FmfjqkpJKKarvxs7SEbI2eqpyy3nTvP1xrzOXIOje9HfGk0bHulIOtb
0uI2cj9irj7dBlUPJpNaFPuREq5qJedfq5PYCZbhkeM4xROIp5RpcKc5zehuTYdv
JE5JHepskTwLKFlzUfssoveLyGwMNCNgYgRCXBq1SXFCR2LJLRCwbxF02qtvr1Zu
DU3NObwqykVsneCfef8qvRGmvKYoFBCbjOawGiEn6ziynXa9+9WfRV4LSAA5GA4C
MmXuXcaylWlq1nlheMo3zG1L3Fh96gtHKb9LmOOYXEHPCdeQ5VgwKk7EYorE0fXW
GvbbENna5LQTAfJQink/x24ZAfhtwXjG7HS/+9Xt4uDhH53zC5ol0wJ4MtxM3ler
u3RbNxXbwJSo4gT0RsmgFniIqhZkdVtULODb4fGiL66sfDnXtfRVuWSQQqUK5tv1
8Gu4pagLg96zXKpkZdK+Q9icJxPlItcU00YcJZbXoo3HWtT101CeL4GamslbJesr
d42RrCW7cJjlW/+hUi+denoeOLP9Z0h4/8U418fC0VZU8mi3V4Ge89nDg3zK4v9F
xYlJC7I7oUV5aI85IN7QC9DhlJIcSFfGy4v4qqX4OcfYQ3abD+0UN36v5/NxZrB8
L5o5D9M75H+SYrod0JYGWuNlKSHTRGOyb2/Z5FJk+PO2QG/Lmm7/5xEsJXOAbKQg
jrr6JK7vmCvWWseAUzufiSuk+CWCxhSTun6FaNQHdm680tMjto269EmIW7YJEhWy
WMmu9cRhFGpq25CCkeg4kWzeKUzErXZB61WpVdGtW2VuIx64lJvDqDshalRBO8XM
zJo7/ALrXxrWh3hH4nB3rXncDZYLhMJTTnurQJXyuE1q/WukOkNtBXo1OVeSMIFA
tc0iTAR1JomfwHIhgEvgnm2U6UUXo0AgBgA3qkh9MoZJ/JI2W1yGmVdueCccXsSP
XGJJhY5NnAJRGTlmt+2xBGQH0oRDB46sxIlRo4NOT/U32HvsQIDbP2Y+6xeU24bE
hG5VtltnS6Xzn3C9Pcb6l+L9gYhklhd9WUodtU8K8gdVKo9VBdEBFBBiCjLP/7gZ
9aQsL/Slxxq5uvPjJnYCBtqrtFKZ72U7dW+ya/FA2h9D6joTdtyOSQ8c/tJ+zMQ7
5T27bwtxTmDwa3vdHI27eNwszPflErySwYPhHYO+chOTiQ+h/Z8jngC9ThKlmvyZ
NLXDaJFeeK2L9cCe/BXalHDO3RTiyAJL+OiCWFZ8ywv3NDhbsQ4DlXxlXHrLdc1I
KgCRCYQTQL77zyd6zFyOFjGFlIB8A4lx7xNE1FyAUIYKN3UeOjcJKPfmu3CWbDXo
xAvDM0/Sm4us2BavyCcLzGHw7SaB9hoyWuo2iLTHwiMHhqyu7Vugp5daa457OQaG
aSQTIzm2QN5fToCXqUX19aAA13p8Wwdas37u+33XgCBS6gf1l1hIrhTiRACdmZT7
xgrDKB6qDI/x8OwdnVP8ZmNGruTd+LKOLfsaVMLvM+vLRGz0xoRo5o3hlOwnbFn4
90YsPT2yJLJCjN3M6T22wSN4aRrqXidqTvuCn+kny+YOVCeU7W7MCZCTw7/MUe6L
u4/jlYN2vBbwhQK+yUwL0l9mcbI1Oao6jmjpz0755Uc5c7MAl3zIqvnfZDM2nYJE
xqqM+ku3YnI897JjLX7nZPHJwmj4+LWSQK3T8OqG34YtTDt41WaFoLZsOQBFzXI5
QgRJRWuKwJbE2VZqFDs9FxfnLnQ4x+Jgksi+9M8QnujogxRif1RXd9iaMLR4xUtq
DGYvhBVf+JzWOS/1OpuxUa1j2jJuXIKxuQ/GlDc5KVleuT8rWqBcXiEzfK9EpGG5
l/VMu1nYfrNDoxZiU1GkCKiNGpX7Tk5XwQ5zbrOTsh0Irk2c7530iOPKLGV2T/Xc
3rVcFHFC2kcY0PH+b+YPcm6QCQne3FfOU6Dn7zSnAC4DMW9Rhyj09TWp8agHBzGt
rVsqBQc7TZhPmVXJenVb2/FXcMr5JNDumihEub8jJcjl4H53/oyCgdplpCyZYcwp
vM+YUfh61Pr4j4DI8iFi/M8brWSsy8Otnm2lwlNXiBlCUgEHo9C4N381pEkWgNZh
OjnTntYhqxHS/RK9iU2P9zpLQriFCstMIGX4PS7RjMvMmKUMWJHYVJCqT0Jmz9nJ
EJdXdGvJct+TtrjrxUtdjG7O0qNpZFLomcCUc0RnX7K0w7KVRpfVEPC1fylRwTkG
oqZ6+yF6x0R0xWiyyB3XAqAeuXkvemxn84au6HlGiaTc9JdMvC2U1EMEQ6iuJMRx
ESYYzT//E1yHNgc1+02PAzBmQSRz8ptLWc45dRB7pRSOym+qucM8Pj0Uh0vU/BpV
c1RHwylYmYLCV5v9W3bzhzUqQNtcmIHkmbuT1JFyEOtUei9ARZl7DltAW8gImtHB
ZSB8ehvY8kjVYchay2eEgy06KTOl1jOkNBFK+Iv4AkI0DDGPEAitpP+kzFhim6bo
FM4JPSTZXXL6KPfie2HzCHKtVPzQZ3YCva84DtxZwJBXhB5qBs4WDPGF/C9Qyzr2
LcOgoZbMisE60ixsT7TgxogzvEecxH3AnG1ZBmahmz6lZlNKOoEWew9lDN86zcAT
JW44fWY88nVF0F6ZornSr2rstq6hU/i9hoEN2lXNTE+5VYmiz2qlnAK86vkh6p16
3Sx8CT/yKQXnTaFNIjza0lz4JjC8rp620kQNCmR9C3CZRyHqUi/eBSTJmHmKbujD
pmgsdUs5gVSvFch5iUBODCUeeEs6/zECKh9qVCXpcKcp6gJSiXDhje/Btqzrdmk2
Yix7N2om3c6ITi+MatD5VOeNaQmSBZh5+zXNJPniN2QLPf19ru5WN5HF2gmJzPbY
tYpBhEBRw7qfTUUHfYJebIVSU6IQOSCn9x0IUmyozMCfV1tP2uEQlm5q91JbFjMT
5AWW0eCVdwkh24tjdsK2h83yGxIRDtCSz+n86klfFcMSZx8HrnnxKc63E7hoWlRb
LRDdMCzejDlRfLh6u95pROPN/qxqfDdgPRqtHidpM96ufFCP3/gAmD5ErEVX/e1r
dCOWBZFklKFOhHqFL5n1+CxzT/zBKtIqgdIbUomTHfuqYX/D7GthYQ5LONCFZgH4
rzrio4H2b00D0s34eOzhrRkXJSRhB/iruRDX9ivmro+y5No1hIoDbNiOXCiqPXxs
Zsb6CeDMb/1Dnkxnzumoo0dyFwzbgNQKLHyYjnHpLx76GHUYByFLAYfsRF+5UTP8
+vwaY2bzaVGv1gAj1DCTpvgjx+USrmN4QVtwkk5glQgpQdqFp59f+q+hZ87VeRqJ
YULMGQzMXZgIUs3ya9IpBpUc9wLMFrlXXrxTPECTi0kYgCX6gi7k+B7idH7o40J8
JkXcFjQZpoGb7JTBAU/2jplsDpI6paqgtYiTnKqgRhmMq6sRTWBYYtOwPCyanEzs
SvW04ZPy+92IJg3qpH5Kt6WAg2642LhbUFl9QZJXA1Fkt7tvh92sMvgO+hEWcFlV
J+MW8C/0U5VqsT/mJNI0J/c5xSMBVKRzu3XzLs6U2+XR0474r5IQquyzC3sZVRKu
BJp8kN+1tVCiq4H5p/fIGXW59ImAC/Zj1Q7+r9XwjBWKlBTnwRMtYHXFUDjurnWf
OA+por6ZqaOXZIIo8gWpXpkEWkW99vEWMDGHZY9NeYI0NPEUCMdfyvM3RPsjtbLU
1EucTqsSNULz1YIC3VPQ7Gs+3ATF/p0sNrOySeu9TJ69LTzP6DBdSaqU8XnHgYRJ
1uExUypBOF+1jEPqs7zAuureUdOozJ4FDgMOBQhxET/K1vCgn9Pr3SarKHv7NhzQ
6hNDax6QgxjbEd/gz92OItZEt8cFhcJ6tx4sA6R5/1kb3PQfUtHPS9pk7iz/gqil
z06DtKY0FQm5Vg80wXrrzP+2MoEuGcFPGxUqEuI7OCSsMXX/1ZB6eHrdHed7fkMJ
B4mt3tpuAzlmP55wCMjQ6QbhoAcT2gy5dw3POX8IuLtysC7yQkn+fHI8ZjEWjwEh
LRmmEW2hJY6wHC0ott77QBYaiHfcOlYV+JSrNC0g0nBDDmGdvHs23HlgR8S5L3Yp
IFOUbREZYhulrNjsGE+YYouNZMkUmMr+Y5eX5fO2AB32C/g8qZi20tjKD82XIA9E
oyu/8XHTZ4s6QbqfuBAQNcfvxqePI8daIxKVrEVnqfz4LsHEXgFRTZD0A1pUK8ru
3Pat/4WV0UKyt4NvEe0PFFPqnChy8yjONja8bAjmv1GxPW5q2ud2XIqkcBTPVgTG
WY8aW54rK2tZCc9F8+d1ZOA/FSf9muOWZyHll6D8m/Advf+S8cRiQBhqHvZJsV4U
60v0b8Thr8hdIZBgFTABgVRpZ2qGvZg1WoOs9CUSzmUvzifwWmVE+u5mB8zJ4cNC
SIcbSoCA9vRJA1mW9zOArVP91HtY3yl0odHLn79HFY8x+fqHHRaJpJnFzH7UQw2D
9UGJNhrJG8rXgkEk45cpTsuYHHWFX3eXFsOA34t/E5Ltw5JqIyhcZMvSUASx0rN/
QOd7BqqmT8/KHdb1NSomsw0hajm6GGuk3n6fKjSClTPf4HLG4A6UxkdoYYnNp9kP
UQxm7iLUBDwaeqjOnBH8RmmnD0rcW00JdnmRGeaZ5HxsDHvQ4LR/8XC4kTuoeChV
NQdfHnSrFDeuLjUmjjD1Jzt0UDqXrcphZAtld0vJCqhfxl34nxsOKbfXjntJ4prr
yeFBNpMVaqBvJDnIQgbOBcZrdpfkwsjUjsyBSjhTZX2kHNovtkVlPmGx/E34HL9r
J4jzQk6YK6VV9VJLZyjQSrV7esHhL9lb31o4G89XrTJADAeEMU6Z6fmjTPUotn38
nCnbRrW8GItIvdGEJS3Z8eGh3H0CsUrCUXN+sq95umTQQQDUiWRuUZsM0T1HMWtT
c2xYnhmLkkkq8C5gjwRlIY9qlYJLI5/r/+fSDxS2lTpbEvXp0Ey2fr7MlPeLlXV1
lozv/LJN1Sxd/wPaPlyiumaFIeKbQrBlinvUxHkvNGGMQ5IxR/hiILtIGnAxJGrJ
LO+I9nYsvm8kYmu4gHup4bn+dHehSFy1IAXQJWjsBFkrHVJQIklLYAzWlsfFGWE2
hGFhDXFPyJSyZTfLnUOfsJiR2rif4VcgPxF2FW88jR/62MCClKse6Wo8Lkfz7yYA
WAzOqAjkdcctq97Jm1dmDB1p6BoiD2ZXGydYx7Z13UaiOn7LLYceJ7F/FBRjt+wQ
ZbIIBO+A//FsihqubxMUiXNKY/MXhqwoxAroujPhU4OSSn/CivY7TcX8D/OCAIZQ
UZOcJ6rE1MGc7FTEjnRC+qrU5f5bHxbbDtequ9wyioBecviS8YnleS8c5mPmj/hj
1uDV02d+8XkzC2HBJpYMWhEFpl2s2gUZMod4DjZ0umI3S8DKjLvGxCZr6UcvJNkb
OKgRqXCFIgVz03VNGe8BSdNLTrnHjDANNishlH7DBAOm+OTBbK3rrkSGN8iBUqpD
zwBnasbEgMD/zNh2p+qI3nFFbN+poRk0/cjo70CQhragCm/EQ+zCs7jvidrp6A3n
xxWMFjnFxY5uW3vQ8aeqJG6qpmBXyaOCh61hDXCQwFw6Bld9tLVoZT2nmz+mxT95
IDIwD32Ydl+cJZRwKVCnTZsWVWmeyNGniwTCtr5QGzWYZJClRXoNI4eoVhDsK2g7
N5SiR+MqCEIl8LgApPPdCp0zyPgZXh8ZbXfrDE/0CS3DZXowqwH8cpdo7NIsCESD
qZaKZU/e3ekdyhr+qrMu1X5UIjPBsQlsopVUBzY+CT9oD47XWnxGm+nNMrXPLs5d
oKWFVIu+PS8AJg8EctIo/i6GPzjY7zI3t+aHopqbrZtHkWM6vm7UkE9FBCARkqJp
42qhfyrA30EmVMzOQU/AlVgrAEpFSA40fCH+VbyHhe8+nTSuXwirS/VkD/shXcwz
udOLpLSB7reRVZDiNKiSVNkcnGU2lqlfGJtdFj/M3wPvstm/RAmtNCsl6nTm94fh
+Padnj4iaYp+KwhRQSpdAuElsMkHX+Y57rSK0MjDRWr9QxmznpapamNpG6wrg7PV
Me6mD6ugQ/OAZgY/i+SqP7p4enGyjNd7fQ1gORTKUOcKg4haF0vLeCfDrbI1eZag
6qK1F+4+98i6gOUg+GiBPzh1XNdMNfqP6ZenUjCcJgGlJsanWXT2oa2FPJSuaAx1
Tpix3hqcAyfdnH1nJs8uhEaXRTJZcntgN+xqHWVlwZMtrYnHM1CijmGIa5j6I8Se
7iIRgtRDdvzzdEy4rwsvyEXj678Ao1lAkpC1qOBdygu56oa+mQimLiaVva6Zmf0y
d/LipF4/RvypqQNuphDtyQj1Rxxqnx23RAwQ163Pkk2wlZYRFCL/FqDXRQC7rXFg
jvzwmSCqj9HHh1oRwLO+fpkc46j0f+1JmqVt36URb33gZEkvh1efKqcm5LaI3zfE
rnnHEEWamOzDXTRQ4re9TegYfp10Rq6wJOVSOGXXmPzHe+vnMlHihdWKsrZNRVS2
rViRZ6H3JoZuJlcNB638FyYIlBPeY4c0txF8JVy1oBvdEazBiWolgZP3MLsW+a5d
8mvcQPfgeZVucmRVW734JbP8O9tAwtSCPeL8uvGoql4SFYvXdMSjmZM2sqWU24yn
4mbbrj3ntXPe2Sci6n1KFLJY1Ct4GauOL0JGfrnxmw7JCV4YNfgXJffq4lEFfJ6Y
CTcEB1e9hh6OXXs8OADTuzFQcUfFkT9/MDzq8Uz/MWcKYq25rVrYJx4k/gTiNkJt
24+NJjoW7vxD73P6g0WCVMwHtAydQy2MyWX8GDH9ITaCsfwqSEptpgcJ5AuNpwsU
fb0CunPhxQF1mvbGJdrdiuC0C/e91/EKqqIrKXbAXJryb/VOsw3wnBwhje2Ou2TN
Pfk+96IrMdza0YNhm3KIHR4GyQNnw7jV1q0ufpHxgVPmIhbS2cM30Cz2rgP4x1Xr
DBpALVhDhmSIkKT3tlyivGfojZQ8qFqzotvFCY5FojvVua9UXQj0UENmeARSL1SU
CDmJWfNehglcXYDB5oIR0rJBFeir3+fQqDBvcx4PwMBd643q1Ivww9qiENgiIqrx
dje6tN0BeCd1QCxJyY9Atp0Mp4LDCzxNH5upPNby4xpufS24MkSSPymF5x6l1ZAr
TrEPk2XSPlBfVtW5hkumzQjiHcl/XwKl0meG2r3JS12P/6DVbyFY3OiYHDhg/ulH
sthEDelvX37fe8UJPM0ZrPDGZHbK8NdvShNaXzZE0BSsg+I1giKVTThRDxwG8nqt
X+7zQxC4PrlwnmVBB5CUYHi0WIoizUFlLCIUV565M8b2vlPNRrL/UFMypX9SOVoX
VWv9iYeWdJ+3T3VbaSCC1O4HNH84L5fcDnYMTnWrCxsECLn+zQZu72SQQOE7GQAs
0D7iTEMsKeOABb2/DTL6dac9XtPb5b1qyu3EQ4n+7WnRT5tNbgDjqBw5WaUNrQHk
E/+LwE9rfAoLIaOQsEmIbOr8psKbyF1CKcG++9pLJWGr8IerGL/WA+JkQX1EpoT2
PaZolPGP6+kIpD5FzkRU6AcOCu2JNeAXetpUvqoWqXW88LzDR2W6W/af7QQG4pXj
5H7dYF7I0UK38+p9OfYSJ3EsipIqeU7v0GVqEoWKKdM6OmlHEqRfO8SV+TwY0qU2
ZikWe4tEQRVNDpelUGPxghJ0zH0u2jZ8veuiJpiRbIXaI4afLZmOBX3HdPOS550w
XEO8wLDhgMN8hPCwiUlLY23Ip/6gSvx4Q9R4871zDlgejQ9HvmyCkqPe0WuxfpIF
51ik25F59VENNnJbCX0bKk1W+gKUmlSf5MeWJL5DvIl7hzzJVYRK93Ne7GBmIJ/b
Wqw04ouWnLORAMe5Ozcyaos0k7bDMIhOto46968S+0I1I7i6qPEL7riZ4t2MKYUS
8WNTiHinEXjfJFZufNKgbQXWQ8AkbSeudNJfNwmOcPfGsScb1qRaoz17auQw8pk8
LtueidjKPDiUCTl2iUokeYvqJQKPhoZ1DqY9sgeka1Jsie9ti9A0BiYQbrSU/75T
1+D/P949i4HHQxdf45bXWeo65b3BfVfqldd54Y2yKX50oBeV/CEn4GiIk4kmSDh0
8rpulQBQAgz8Vffk0GcJtN0yDTS42Tfvv3wRYojGnRG3fMDRh7cszDr1yr5Hbm9n
/prZqye0AoK6ogrv6+NJ3guiFVDhXJIDdGyaKVallljY+GynbgFZYqG4FoYDRLBR
S/XMVqhh/Xa0ZPAx161azXpha3pfg22D5/msBX3YOpL1FVSsw07gQogR2q5vqKVE
njdkraR/XjxnD7hpRKzmRJIGzaRxzarFjcPqgqBhNXXjZk6WJTJ6JdCQBLvpVuEG
BOe5NaZhtMqDtIhume0fjeA+HrLk8H4M3Eco6pUVcvmKb3LaYKFOatcJ1R57VWF/
yuDdXtrOD0gPdjzQvlunLA7G0NopRaxyyFQMaWCLFzvIEtsB08VWZlcGQWmCUc39
8MODpFGJZAPz8MoHMH/SqaQbi1ALeJTK1YLaEe22jk3qeoJUSVk9hEYNwlZ+WnqR
5J+tDRFc+BK6m3gVOS3VDD5glgJVK0z3iYB+H+iH7chVU51AcVBZ/WB4DTH07IkT
qAT2YYt+mNZkupuUpaM+7eNdZJul60yY8O0Ab7qcgYV/YSBrv7ZaTEjv1UwTDU5s
E6xd9gQvio3GXvGGIOK/O24XychKrcRQTeBB4nWlmHC7e4jwVSDIcGIftvg0+hjk
LY1j5BjjZdGPDuYxGMRDaJEDs/NzwGNzQjKJRsJdSkNdOS9fUoCN6zAojMLFDpU0
Ec2fTVjvHeHh3QLSolb0/HaHgG7/9bLOiz/juB9RvF1KpVYENiO4GEG++nqngRiw
1ikypRAR1MgZ7DVkRJMucvgbh7KH6mruErel3bQwg9jGEM9arDj4YG2cwMzuFqCc
/yybeBumyxhNsP1y8/qhCtzdgDqzO4S7kggMfWGDJ/rVm5A2OpU78LqqGqRlLah8
daTUtBnQovv1ga9hNtYNwr6r1FRGa9/arErlWDipqMtHihWrPP9OKbeIG0HM4iFv
pJgIjZ12kS1HUYCDzGqoWDppaPuM4MLlnfo990/Hq6qpolCNyoYwiwgYKpNcQiIr
9pIsJ7op/bLUSxSwl2wjYU2L5S/pR7td4EpFawX5H3kbcr41mLWbxs3RZYTx7/wq
OuhCIgLznTx5iRGFfeceaoxjHrK/hw+DC43t+wacpmiu+F19ctn4RytjoipXnPIy
m4FIYgsbpSZc37qsk5Pj2FDOfcVtFD+XlVFROnc+fIHvb8k53Ck7DwIhiZkdebG7
zoCsqyWzeQyUeuLaUuVZ0oPTQvr0CpDBRYA7K5Xecwn/g1advHbFJi4ukjV2r+aG
E8PWOHpDLGm+dfUzVGLoYAsl7mZBNPiS2WgVE9QGFhZs+WulN95khTL3i/jz4uis
sychKR4UFDrzTMXXnhf6Lg15HsV7mFg9pPaLHuj4mGln4OLZMz1I3xzbP7NdZvpP
MpjEMaFaiBW5QB+Jev9allUKhsr2NkLLtnEg/kxpDiNl/ILXzYeR5Nnx0p8ibMd7
9tsXqbx4uTE8InCdEC2Wk+XgZlcllE/7RKVe865af1/gJdn0gdNFN95IoBMOC2Sy
hwyGm8bhlJqdMUN5qgmGyTO+vSRjlo9o/RfqO2XeDOkQmzuiGLVMGa7VSVNmUV4G
1GepeKhnk8kYxKlP3VCMgJ0UOIPniPxXnnSeuwD593pecaZl3RBzvYIHwI3PU0Cf
wKgXAaPaARXl+/htsKSADg7277y6Fp2pP8yr4iUKChwX1P/ZVbuWqHYP7tLjbmNS
ZT5wy8uTc0WtQGeyyDCEbwtZ2KGJCJs3V5tgKn6LqXIt+EnYw7ejupl6P/nB9pOv
WQlRZ7RsJeiHL77szhm2wYCiNet1VJn0SUCoVOdEWYthSDLszkTibxzmZ34Mj9Cp
OH8oVB4fP8VAOdg1dDIBk+EDLd7J1nD4Ay+9rE/LuPsKJ8/wdv3rv+C6ubx+SjQc
0FiVpC2lo4gN8pvkAt86CdzHJX5QIu+wlz9KDAPhVIokDfkENOQlB0nlvzGNAE16
lQFm8jPFkJ/E/L/19BhSYD+YL7M5/mfOmNOgwCqPW7Ay0uKholyZWrRIfv99Lz3F
fvQP45HliY/E5M7POa5nJojAxL0Krx7S8pU7fml25iOBWtHlJobv2WY31as37dSm
cd8gmsa/gBxvG29SIX50+LnJP6j2eCKRYTs3abXPBJllP5VyejPR2+FMl5EMXOBY
au1CzjUOX839B0o0OWSj9ZNvPCUXJSh78uNPmzHpqziwR/GcBLoXOysSOqE8gxgn
TARJthcy9Ja8cfC9S1TN4vfQrkJZimwyQyCHtC7E9YkEg2QtESYtMR7teXi6K6rj
itx5VV0yDp2OFLF0XHuhGPTGQqHVvX0GyPh+mC2+ns9FyFRBrDp+Uy4GmHm7WemC
E3bAs7+RKmP856pKtCJjLQ1JqxsFJ7uPMH3tZM8X0KYyDpN2CjcizZJM8b6Mnkj8
xGXUzNJD+OvwyupGvNtwCVl5jlEE7mDqv61Eplya8dc4u8t85LNKP1YHFsaWRwzR
DBxkZlnZ46otkf1dWGoxUPCQF+SHJ4ZKXfDpcfLQYVkv2x3DiXxLOaKTopCrpCWR
CR8rG/ZKw4TOwFEcqeSZuAj42spxoXb6oszJU4EswxRYalCGXanIPrWIa2z91T3S
5SSsCvxWG3e96CUNEhupDKW2K402g2YfJJJy1A199EUKE/pWO+wCmpvIsuzxhBGY
pdM8FUSIdYU+Ax8O62S6VSov1Scozo7DD4yJnYpcVNVdTTVJmz6PFseowZ2npKZO
FP7HWU2hAMTDca4Mk08Nylu94aycsc5txmcqhPiuAe7foPlIXPyWkJK8Hfxh4HQC
4OywTjaLub6olQS8IKQRBolCnfTsrAnlEI8HZj5njh9Es/X15WtfO2kobvwICE+p
3c6tvDxQu4HwOUsxyHjgqC8jThYrFSAX3nHZL0gtVwd7yobg7jvb1OccTAZaIx7T
qswK8PRKMjElDcOsGLbPtmsKXPsGAnl7nPRARGpWrorrGoRDeMcRm0trf35PNF/i
/gKhIt7xaRy/o3uLCqyORIv+E5vMS1Kj32nUMFGHvap7qQuyy3poC/zNp9E0bkIa
jZoy4gwGEu+RApoC8oalN36CuNGYcg3zoNpjYJFwcvTg4I5zPPOOdfi26mn9/emS
mRc3WdsbVRNWZwKbc81dK1O7zZT60ejYlzXviFhBwNnvUJmKgVqpoYfaYwN8tVyQ
GnqD9D9JHc+hR/IckEwSF4tnbJht3qYU0KsfccObPiUR5RVf4nIPVAEFvWgxKjBT
zyh2nZOubQjb5Z1/8imlV0WPkqUJ7Sc3APpEUpowcoiZ1TriO8vP/nQHrhWCMCLU
Qupg9Z7PcmPHG7/XCwRlEiYpyAIYjoW4vFA/qv0QZ2FBpw0TT4v3msDiaaUmfL2c
yF5wpeGNhsWvRXtGwDV2iNkSQsabaU44oQAwVVSh7ZfgU3SESyhqiF4dCIPm9h4G
AnLK8ZncMl0ZZGbZe5A0aS0CV47lspyHzUKAxPyG+mSAJM8e80ojMfUgN4TvnhaQ
izvv7LCxCgriyVQKSN1Oze3viaLoMqsuLghXIHw4cvNVY6W+8tpc7QQg/F9ef/kK
6Ka39Zr8/eEQMLBYwU3/NlJi7NVFGoMN2T7rNZcyMzsZfr8apvIobl3BN+93cWY4
Bzkfrs0wOO7aqH37UYkmGl4L8fxhhhtWWPH98UkFa5Oo1RGXMuDltcxIqJwCbYPi
iD44jMn3Lwdu4ut3SAHeRph5YswN+ka6ZItSSS6aKQQ4wvRYBuuPCbLdDfqmwwYy
k1zLsBR8ZQDpEs8BAynEfj+5YRAwml+qyNJ5JTyCUqhWhSSNarQKgUAUVAUKAdbG
SmGn03DFGau+j6ufMiwtM3qzmapM/7ZNN0qmMQOgZQJaUje6YeXok7PIRqM/hDxI
xbjLSxaOu+PVBWcUTwlBOWd4+jho2zX2CBCZi+dJKuN2T1NM3ELwacW5qyWtgQDi
WSs5rHK1wSrnVwc0F95f1Ca22zW4D2lN3kvLjV2/lGPV+8DY72rV02dv7jyEYJ/0
K1fTim7AsFilD47hBy3/r3mizk2dENWe7iEX+zvw3xJDnvKdvy5WuN74o/EYULF+
61uPjBCkLStaoblIul/HuFfd6gHEzaVkNCpHUSufGYihgEaCoRB1DRMcJ3Fl68sI
lr2exF9gs57Y9p6kDN3EWKF/GPIbl8aYmttiCjL2swH07i/9CLeuONUX+u/AmfTE
l8rGz7XZrHhBK597iger/FE8adm822CI/EakoTBKDVsbOyBuYVZ5rLnHDg280ooP
hMCf3ZZL3g6BnDp66hjd2WL+GynjTaMdw9iBAmWU9Zh0zSD60lUdebI58/zY7DtZ
Ml6CdHSix03XUGsYEw4NbyviNri7K5r/kds5yDeptVXkEOvsG8SbT7BD04Cu4h0R
vX3Yhjc8/yb86VpeC0UrXbehHgkWYe8bfT/+cnp3XyiNZ+vGwiA3jnNP4vi3aihD
KXkXJ7F0B0/D/xpOp1/apFhyWXkM5p1rNPeYd371Te90p56WmvAcL6Q1tbuUSRc2
WSsy737DOx1WELjdoM9kZIeV6UdIyw8PPRDP1a4q8d+WTflIDBuVZcuImemtnTQK
Zd4deotm/blEXCPuk+Ob7KDrkbA20+fLZlwW+W5ObTInOvdj65Zvt51sdnRqKkDu
nbFB2qnZQL3a9s/KswciKCUlJP2PYmartJeMNSkeC7pqFXaVasXNGOcGczDxP8HL
h4HT9O5MVw8pNiD87+MMTXK8rAHXZGeMFlhM7DOpPzEiC8zo6sl34QzJ0sTJE8CF
195iPyl+bmAIJewtLsmmrqD7DMaFBhL2KtkS8lEGC1N0pezbR7HAh2n/6SUoQEw+
bRT1xA7v7hP8JFM+Erg8BeO7/6qGWDg3JDU5FyJYcJ/gwvLqXdH24+wVCLsJLdjV
9GuhSzWG0hvTM2m/WuGscUvg0Nx/Eg/URb7ADneSXu8OJD72CzVshb227KYCR9Af
wDuELdZuBkrSd4c02cxpKrhTm6kujzbZAQNVOjc12oWtntRp+aFRO7clEwxWNwJW
mgF1Ow2+wu65QZoqKez3v89myPL+LvZXdZp/eVAnvI7hA59vnFOPGHxsT0GyavNm
+kggcAD1D/JILO+IsNw3iP+UVNwhc3KvS760bZDn8GyFWc7YKKVtE7mA+2A+Xy9h
wrVHGv1z5SRGMMSd/6ClbZ+r5tFw5TkEvgQ24C8ckG0xUNcEV2iweGUkQduIuHBe
HVtQhUr8kuZfw/S33JCT5LmcKGaqZYEp0asKXaTosaHl9wFuf0tVn5HMfa46p1hB
IYFubdn36H8WiTL4UoTL6gCQ8d3gFHhoXv2u4criP9i1BQZgsdRsCad9wpJhUDTW
9hWv7HdfIhD4bxGvJ+KjWsWZG40gc/VTgmzd40Z5iunMAMIVXZ5cbNI7885k0UTo
m4J1O0N4JLA41eDXEc/SA7jMUvYOqOjuwv5cEefEFpBwHSlR4USZCpjK/bCncBaV
bjrrTUdDcbY6C/utA/l6TjaTWcCrRxIsYoTM/97Gw6cXvGCEDcwBaEjxyP4NdHhG
w4/SKpGWNYkocvvJeBKAVXLc1RJOu7RAHALSDD7Ie7cTcjaWSWX+GoXjN0dtNAiN
3wkmFnval4/buEKaV10ztoWgcUl7J3Prs/tROD+hyYBHOEpGRH409KFtcUGLe7I5
50kDz/3Mcuj1wQ0BEIRz94xHbOHEQN27FXoGahWSeGbKkVpZY2EmCsivnm7olUSr
bG4vzbzGMSJ6cKwwgTPaO70gGOuddt0R4s/y8K86W55Wu7Xktz+AeYbUcGZpz2hC
pfaALhiCBufSL/d5NfBBS9Fc9vIkiUusk8J3r+DH36E9OFUPXW8TuZeF7vj6o/Qa
Hc0fg4EXykfNC5xm3Qe7WUh8RenTgz4a9vhFmfUik3GomQEubG/ldbvXq0tprUoB
6gseju8mgvxku3fNzotDKwSHPxzqClMigplWVQgf3DJ0+1cIVha8ote6FlJ0aFN3
Cc6KxCX9hgGMuCVX2RcWutokqosA1WT9gWOdxThI/m2VcPFY1wnvF2GzJdOpcMDp
IEOGsCI9InlClbaiKMQM124FrK5QqlqR0Y/mnrs0Zb2LahQFTal7fcvBKNHBwzh7
FvmRmICVa8qT12PNDLURI8zXkssSUFTuT4PHQmAayurk1xDLNfEdLX+pvB/+xuj1
jIs9xKuhBI1OrvNXNI+zMLlbmpAeLowYIG/RAdx9ZL3b+Y4g86plfSoNwozufnbW
y+T+MbGv+qF0ApzyHXKVqDahRNvxwvm5Ou4/McOZaC3ZPQT94G9NMCHvJhUJy850
nUNho/9grx6KFOOZKLJNLaoRE73f1NygqxHQp8rX2gmBX6joCwlgezp/vkhM3mmn
P0XZj35FgLhJcJfmd6Ub4XCw1fSs4oU9XxTRU764sqAaFZidE6ZAXu5by41r6Xi2
3frCUTfSVKxS0TUf5OUOrJzaYpVeEcWUa3jzcODZJ5tFR4A+R+HM+C6XjWnW00RQ
juLZX0wPzZi6NQbzzEQJHpeAvEz39DCDnPCFjehGDSSBATqs6qi/FE0UbYFlCGWq
2uJiZ3WcpA03aVamaUJvgBm6fNaToJa+UrVtd6G+WQYu6YLoG+TYiFWib7Sahyd4
JxTY3etZrMsqMCkcx393N8NLMWmRetNxD89tQ7ZJgSYKzvhgvKiWPP9N0r++hapO
MXak/IZiTeYfQSmH50fhEZ8EU9nOOumcagaEkt28mBiODDyK+WuwOlGx8ROomkb4
7F+XlSPe6zFWXPekV+HCqd5vcCTP4PGjqpN360b5j637dcfY8sUYttuEm2WF2f3j
9jGfYwkJdeckJ6Zhhm5iWZBDClETaLH4RtK1PCEB2FFZWgTY/wlyRmCMbux2nrYF
VoFcHzB3kpvoUYuWyT8+CjdPKBHbeuOHIDtOT25i3ywlpPaohdlL8OE+dV0RuzFn
qaxvloXsYkDOdsCg01gazUQMDEWf8O90+GKdObcUFbx0F1ZLgASWWnf9LPJ0fQtI
HZmbDvIwL6bL6rc5bPDiAtG6UVa7AY9SJkxOPsPai7YE70tCteZN9lm57Ql96vEx
QhkHTAMJgNEs9cH2So1mB9cD/qFaAV1DZ0SU774afYr8a11VL73iEgV74e2qmKXc
XN2rqLlO0qs/LH7Iq6jINmEEuUN5EKi42/qyzEZpFjEfqDSJ6Vksv1B8snKOuqoo
HNDexP70x3FZefLxtJYeSpeuBqcoymPA5cUgpcBfpKgudSUA8NeRDXtkpLNrN1Uc
j0ZL1Jv8j7RRbjslLVjWc0xK7w4BNy1g/wyx3++yz1UUe/XSOhVfzh3RGR27PVhm
i684saTDmptkIjF/GyZKbH1b9mIVAsnAYyHvO2iCBN3JrD9RcVXp6miYvIAU5WYO
rvNo5XB7bgDCRZdlcLSzyz60wKxze/BzXEKAbfGrOf1LTy8chKPdInMUclPrCdMj
2GgMrFK9cx4NyX8sENVi1UXrwhLJvWwv3dk/Edo5QZflCMO03DNxS7EVFgdK9GuE
EN56/+FM1/JkHHV9Acgbcv8c1D5hK0vLVJCpExI6UObMP0nZwQ/Mxt3xN30dfeed
IavLLl4jlmExAx5BAVut/4w0UVbNYTV+UeUHNg638bppkMBBC5jrvfeit041jO/+
EW3a8iCTfSmYmpcQ95CD2L3sCghJRoVOzKd1xStz7Eb6aVxOKM2ErKuPFJmmYzVu
8Pi7Xb+zEh1kekyYZo2hYvXUnn8cGxnNZ1cxU8s2i1MeeL96SVaHKRiQZtiVU1KU
rf8ZHpwp/mI8ALXXcHbWcjW+YYDGwFokx2wsCrZlDLdZj7cRgN/VzfANaWubcfG/
lqsrTWHZJGcA8zFNIDdlRsiqgZILuzA/fQp0lYKWCBbdjBIPgYe2vl8nZji29snJ
1/68luGuRrnqBC9GIeFk68lbCSQKTrS1SC/XLl5BxjajTzBnNYkAXoeqsv+R+lSn
U6jyy+YFkSWtqsTXguDKEMOQzcf+kn2+VVrYgdW3ZSfxExpWFsrgNoOcbMHs5hJc
rq4/BH2AgIWI31gN0IqzJVMsHZs7Cgac7aSBH0pOZnRVxpWgftdbDtUq7sdbYoWG
7LmiLFv/CuetOs4WKuscveghYsG3NxgffQ0daznEeWI2NWP7Jp2I+rtZg6GjDBsB
apt47WSop6I2F0BzIhs78KOwuq+HoRmvbELJLpDr/RYttc0+7xEB2xTgwmeGiOr0
0fA6ofTNQ5bGuInESSAlfQ6lN/L9inPKtMYsfvMt1vkpjB42zGm3qGGsvSX7/xYf
NFD5SgeJfUvn6j8n3aNdrYnoJkiVHhWEGk8k7arkii0N4pe4BnxXmj0U2WmT0r70
l4mN83q9GgPo9lsdXQkvyvris7ZjKuO1t2/GpFQ9QBBAQPCQKsgAwCVoE+y+wRdT
hUsTAhI5ODvB9PyhPFuSOQseNykX6dw1PqryFLgmuGXRB8+G/IEnGhL/Urt6rRwO
KiyTJu3ZI714JLHKI/565gHapCMpqzq5SRAbBStS7nCnfHUMEHeeZZRro25Bhigt
c9TUn53nTCzdV9sNXPQbjYXlgXh97AQQZYjx1Pou9gAFIum40IbiKvcMPWIcFFLi
mXOeM1O9Y8/zXVBPQaF2Up5l6xIPLj5M/TiYqx0fNG9C+MUZ1wI5DZztqt1RSSjr
NsuAhBIIXC7MiJ3vtIX85nC/fq2dksfKTLbDpSjJDrWMQKjcf6MljCmZ6M5yCdI8
83mhLgsxcwWAQ3Xn+1Oc+NMLb7/Oh7ClQz6YtWrmU0svaMYMGy6uIre3E0qJOIe9
Wy41g/SoqRgCGjQ/Ex7IzkA/9MzfXPjclJtMtXwlWvoz8l93bR+2aI08LFgm/WHO
z95a8CKEVBpn10No0XM5H3dfD6cI7QvLpEDd5sqYgTXsPB2QnICvMAtDnpzRzjVR
M1w6ISxTW0IOxy41/tMX4dasi5BuWeztFXyIPkst0Dz5Ig/Se1ZzsbxPbdCcDd14
Bo8TBX+XVms4xW6eVBRLZBLJsILoYXunahzIDuwGYONqtnDvzmAsku9LDH4LJoSE
tUsRQyov2uG+vOvBSVLZT87Bw+9OaXmhNGuu3mGuIsyxkDWvou6YdSGpGWA1f9Mu
pmDzGvKxtEqUDrRiSnLUciKU7yD8wG4t0VUhoA+9GQz246ByRKFPrAiZF0E3CjH1
vq39FMVOyQomCzhsnd/DnZMJkM9LD23pBlOvkfV/j86Flq+yXjufoR2uYlAwbXzZ
Hz5z5WPKla3jYMQVUvYfFnA7ntIMOy3WvrL/+baFX5yyb5DcHPns/NHroTAua+MZ
IddZheXUwQe3dAFHpqlRxYRaYxbd5wUa/t05v9Pvs5dgcG8dRdpafXOLqjUT92sX
44bwVrH/DZ0Fs09HNwumdFyrstSkTP2y1RPtc0wgpaZSbvo6JOEla4ex4ocffKLj
Lb4dOL/3Dc3J8i9uUzAk9S3Bcaqz5zEz1c/B37V1BMQzQ4A2YqeSi2fNUzeLppaO
/p53vJJQJjeTdi0PkstO0G5rIKtNyP4OMYo+bFfQ2qgsIPYTIms0AbmmqTv1RYyf
SB7fgR2r4h28ysdtBuziWozbB0G2gdwTCrVdPL+WqVC8B6i9EuFFNnZYncY8gyYl
11xJAueyOiDXSqXZcbNByHnNzhYdtBW6BRv4hO6rpgQxsu8BlOTyStu+zUQM0CMv
eCAIyU2XpYIslytl1fGjJcJcV1a/r5eclcSe8iojA0K9TIx0AdwDBfTfuDw5gGAL
Oyfee9QzWaNFsmNUOrLtt/a/3BLMc75B/tQJEJAElTMin5+EsPHKhBw5ltj1GYRk
y1xdOnLCsZNccrmbGsNNTL/4XxWNpa3Ae9Ur2l7JLinBCZHw0AOMlcVtw74wiLad
3ajguKMHg1o4tcdAd76dSGYe+30z7Y7G/EFrnXsc6MQJU0Md/GFslCg2vP7seXWl
7u9gsY5r9lGzcWScklx6l6O7bIhFn9DwAKCjUHMsjAwmTum2iwYQcK+tdwpYqNf8
zt9zU1r2UdAl4x00S0hizvlLDb9Y0BesSObLfL/+FMuY4NtMt0g5c8YN9OMDHb9b
3Tiwp3xWCzyprxtB8zfpGyZ2tOIypx+YMXa2h5sVOHPs7+O/yH7C2vJfVjF2A7IJ
zm4DPtefFnswQy6b6VUyqUm4B5AMrudzZ7PiodVfC3a0QV5/QVBuvNhSJGlTDdQZ
GcZpSwuQAeUzdQ/awB6hNyJ/2SkAuZBRLqsJAAHtDd26h0tzotIwkEf+o1Rv2fFh
RTsh3NaPsZ5jyXF8Kky1t8tgQWmeB4hhi3UVd4l8rVECnHqfgKWCWnwKYEyG6T5X
q9sCsKQM2EKEYLlqthARcbZy9wBSYrwFywsnFWmHmRr4pqGSeJS3X65GSghx8BBK
Ip16c6F/hls8PdcZGt2bzrjQr2Dj29QDS9dHdL7p1BcmKy8MkwlIKLU1GlAHIGaf
ym7LL8wNudOOxDAeoueTtsV5KKEq9ZLwb5RD0ixMNHnACLX+DqM2kMYzw0I/+ju1
tWklGNUud0tHK8I33IajkIJZvWPHDpPvf1u7e4ghs6IzgS/F4RPaBxVYgLvq6xmJ
Gf5K7ky1TnjY1+hnS9wapwcogr1i9Do2HNY0oLOHhvKuRF9+zfR9H5KzzTdUI2J8
2+H6cDjJ6+/03fidF91Hcpsy/wJR7lpigLcE3xiPWaqPVgu6DpyMDbAZOU3BpLQH
rI77O1pD7xbOvUmjRa0tCSuD//1+DrtGG6HmuvQFFkNHXKym9bkkL0lCCmAVlECf
kNRo5aRX1ax2OT+ICBjr3wI/X8akaqwOQCwwXM9FGaeABEM1kpaplgz6Gi0z11Wr
0Z2edo9Zz2PetQInJ9o+32UQOpMfxMPpU8bnFKyvkH/x2t71W8UIMWwzH2/jq+cX
mV+JgIRLGM7lby8v/omp7wEKvEVUvoishNGve/ftdYqx/NnYR01FyjiXRnSRUrFM
4MeNy9YiTAcs85h/bmnOOpIa7EZjUopHZViHOHdm1ML7TqpM3A65DOgCd4L//Ezg
TXjbBnS5KBfohn0wubStLS/YHlc8mEaQTwSnl6zklN1hcVrWD43Ci8omFI979LJ8
VyrqUdLxHQkkI1XG69Hfti3K7W1PDU9AfAHOdCc+ULQVUBVzKCpfEisFxLEJ/wa9
ANGE6e8iyn1G4ZkN85wrckovt1WKg1eDZXrXweFsjJsr9CiHYr4ITQCYoZML1Hlj
3oGKKRIhgoC9Uwl9qyzgjDjio1MlddH7ikLC3ewFjKsIGiUzzDxcIHWhMA67H0qs
fkCxac/IdjEwIAvaIwgQyWKYTy9w04mhQC3+8X1agZdbX9j3gRmszgnsMPdI99vI
R7PQ4ta8G+TYeK8aVo09g+rjjEUzwWH0QyAHYrQTCDtHsOgchAZmqylO/Wb05H/u
of5wz5DWN5EkkbvsHGSrOQbnMsi670R4kkPPKxn3Eg3EUAlgByHfswBOEBvVNwSS
u41Z1nsW6TnBZHWq4HYNSV640YVC5iz+HxgSEv5cMHVNYhM3Twr58aCWh5ZIBVB0
wlmC1KpVAavUqn4b4k8ShwGytIg5ys/nXj9eolgbMiWzZiX1ThdmA2UUwO1DKaLN
DkFvaOnm79gIybYcrgUEYIcT224aoOF6AbC4m83ZlOaIAELTJUnxP27zOrpT4BHC
YwyKsg/asrCQQuw350JE1nrsjUt9dvzVz4cZZ6z8bVVvXBrWLLiZCDxzmW/Rl5LK
zvHSY2Rf4dP8I4HkJLk4UIm5/MQuOoi6Llh2hN0RMMzZpGxxPS8r7s115Rb9b6iJ
8cR/Ste861dOqe1jF3MTmjD88W6KhU+t9dfDj6Uqke/OIVtkHQ13VdlcjH0Cjb43
sUMrwROEQBqrcobbzgtNcdyJ1mojNQyM31KGmOgUtbMOd/STPdSNdvwZIV11Wsrj
ql72fMAjflsSHLIf8eHvCQTPHU1Pdrj+HCYlEiJnT0KUF1mwjEu4c+p1fwfQyszX
LH8Q/A1CQo6UQRZvcA81ALDr07pnr4ZcI5djsIBRc/dFvhcH5Sp08/r4VUcK1Cps
WyzwhEPILyIoEgDSsxFAM/JZwbwBkamhbCEm2eZYT3eLXui32LrX8UzI1otzp6hC
71AUMfKlUOTK21t1RNExHTF1vwNHy8MRB33MO/zSe+zZBtPa9DO3E40picpPP6Oq
QqMy1PVfoVTZVPCwuhp25Ye5tGA9tBZ9dz986ZwR7XeknQ6Tpm5Znu1LAveD7vL3
9XFzRUd45onZQeOzM40DXgxyN5aCpUv5oou66jZdF8Wdb56Hbg0WQIgh56mIOsR1
oPf6F6fB7OII3vKr7VEpRw/B4+connVWXkac8Ntd8MNIuIqHypUCdw33k96gZrNw
SiwLXqLiUHlVaYt+g3Kg0JvPHvt+UccMp8ujiHLx8ceIeW5loxljAKnOBwxjKwzG
KzFg4BuSiv1XUCVBIhk2Ioybutu+07iI/bSw+W7FljuNSkKs6GtyEnys5byxbJzh
gse7CDF9ier7kAhmXIZkbplUTBrDqFU5qknT6akfEpY6dlleEubm/IaW0gZIYpGg
pItnNmDXnIDNj6U/tCJkYDGhSOydMNQH4hyHQhWbM+AY+tmqGr4MmNXvaPziFMHx
a/dboGUFAhKcbe/WWLw+5FVXNCJeFLBvpqJFuGFwzZJVfsTUnznJdl4+dBJmHKX3
A9jt5MANYzfpbwTSQD4kWA7+NzSoGd1NrUCYdXd+7tMLcZVAdfOeyl2FqZdWWALY
Bl3YFB7ZQvVLcLper9VXw7RUFUr7OowVNwqNKXxWFo9fHKF9MFPAk4/R9tV1fyQ0
D9icE23kJ6Ye1u++Fy34hGhCI1a0cTNV3XszR4nS685oTeGQVIr06QL0kOdspNdN
Zg0UA8jjMMXB5/np4V3VxgNREIXRTYc9uY0iGP3mS675hhcCpyU6eNwxK1ZG982V
BpBnucvA0+R9vYJMMNWSjx/Q3RQ+F9uQkwtl/alLr5dppsusZ1HpfRaw9y4MQD5k
mdjVo0bZFYYG1td5spIeVjCMjxhleUatYTbrVselYFRxh1zbrEkKeqt1MwikGr/y
/j1TBzRbU2x5leECldNmvxJgtgyhin3PfZJXnGPcWrm1HJ/3dgq0ISXAkhC15983
VOFGF9gwhqc1ODY2JBRZr+vdRFPKO+5ybLfPnSUkEDqKzDORo3kfsabTMHF7jitL
ZTN9FJpzEPjFRTYg4IZEOK9Z1kuWx0pH7oGivC8RhRU1b6wmCBQSV3PoeF3C9EDB
mmJjiapZyG16rNKbghncmQ7zMhWenOSexW/nQ1OzkJ1F5YGigWWWCkgt38W9x8MZ
cQ/TRP//xfK/AcfGKv4NFpVYwYgDBA3GH7YcOWdb6h9+WG2LUHjVG2reF8nDWeNe
CNd3mDN/LhgKtt73xpInHuq7M/DhNIaXWpGcM139ylcKRmafDw6v3j0YOCUNrCrW
C7x4zvmvEXn9mFB44r/uFLyF+131ejn3MqiUu7iVVC729Uq2VzKszrnirTkmz9pB
v30m+wu8Kvms47tXXC8jVwUIYwmqM5oFSA2bg2GDdHYGNax7vKMr1Q0dznT2zCpN
5DSldVEBJG13ucT+ejVhBI9AZs7IOcUTF2nhW0BzWJVMyvjGsHc7vuqZAi4NVDPS
sl+BdhyYXD3wk1v6RXWiGgwYLWcPM9JgF31a78+5t5qbjH0EajBBtYXd64NtLJnH
EbPN9aoqM67+U4zHU0RmQ5nDzgqZGdBKvSFZgBjL24u6aW0XjtlcSFW/nB6/lRwo
TV1Z8AZYTSkYFg/XZ0ZMee0nOzTiPWgbvRrhLpDfKDDWFa63ZhgYq9k0S73yQDI4
0Cz31IrIE4La+mbc48A0xvw7A3g/CBH1wggSNJeRv762JNKMqkymubhnH3wfDTn/
rJHkTEGBHsbUAeg/F2VWiVQjvNzPPY47rmq5zJCXUKyWhHQSU6h+ZVqk9J2xRMSw
lKSJLnI8wKlXxbtLUxItnk2gqRDNEKUWWdYzS6AGU4LklfQvth2mGBIudCbl18oi
+nI4MQpVjE9JzxaO5NHX7C41cbcuk+/RNyYxMqdWpDVCv+lMJbOhTkT0dDQ3S14V
LGlTBqduXe8YJcYfdc6/yZSxoEIzPJhaFsASkfFJq5HpZH+9xuUqfRscHk2AFNQD
ba6cJnt8htIQFF9zZ/zBcHjYcSl/EdciNXG3luRsMC7UOVR6IFVKsBOZHGoZfINp
cWqEUKwZDY6CisoSEdBjuK0eGRoUwY93Px6PioFvICtVo6fZ3thbyjCGVK++aIvY
bdWj77+zecfBcThmgAcEh0MMGzecikWovELx5CasfIdt/GPB+6TpXRlRUXlLOyak
uj/rhkz4Pz/CHD10czQcwjIvT94MEg6EchPDsPGujuSqyLj5F71aAvRS71tHEaB6
KYcuXqcekAD1G8KMUap6pcYwLXB/zwWgS00A0HutYizYvfq/Nz5JK5JnsmmInfJa
Zvxm0QTUoaAxWwtdzuXkCEiAjWP/Arb2OW1LsSzPu2c+IEx7XfHb9Bf5vDvp/ZDh
udN6PVfLkObaA/tcK+qnQVzZ8/rgwNdEUM1wiVjjBHjJKa64M4OpRX5En391ASgE
vDu9SSWCDacsTWWHnUUr4qSnnfHzptf9nfVFmMhTs11bxwkY/ErxUafnWVQWLz6Q
Aktq6F23aSQ8OtCjIg2CAx2dZ6kDwHmcjWaftIk7OmVlocOIx2rCPZC17Wu1wzQU
JxUL1t50h8Riv15vvueUpmEUwL0/3nOQn7Xc+ea6JmKyP1yl8DHlVeA5iEQ7qO9f
u07f1nYjvJsaXbG9Yhbz09C1z0ONHeFLmRPojkevV5F+/aWg7zloFR0P1cI7fw1g
N4Rc9oahqzWEl6zRQOVORIcLRtnK6tqI6FFB6cgPFudqDAqi7DgGtNkqEomek7Vi
8QM3MHfknQiC/tN4iclAYM863XCtUm9jmOWKhokT6/8Ww2O8o7Ur0uopL8fYq24O
diSM50JTAlm9V6ZZmq6Fy/YLbJAD+QQYFySE5Sn2OLSJ9LkwDPMR08c7Dn68EpzK
5bTgHNsIW1IXec7aAb7I+Mb+x4Qi8pieAY4jlnH/F3vjd61OkMzelrUoNmc/Nazv
G/m7p1Y6vSYNUd1lI7bYz0vVsht/xx11gmTWxLSWs2igIYM3RPVji0GE7hP7c+uD
nSKMxYYauEJGvHWdyv0MqbyiTQ+K06mZRQ3TyEw1maYzvMLxT4KDmT8GKdWN+Vjt
2SIBXILvO3kx5bvN36O26+GBK6GkR+/xD1XAI1YTEd0rmlYWLjN58TsBKuHNjOVR
WQEeVfRk1ScjSNTLUbsTVIAxDWSc4evXLfTeMyqmLJvHWFu074LXNb2G1OGpa5Dh
Mtpm3mVoCdAdSxNCJUrt+Wl/7CijKWQTOX/n4/j68q+dKgGhHIbqzQr6QEgfLddv
7yVEpXeJuYxeLzJh4O9fxGEBYQdWeRF55Gdy8afRkGYnRpGzCo5AAc+pTSfra2EB
IlB3FWtUnJxnghsAAJuXwFYT2iGRK0EafJyjKv0oaIreLJnU3gU848N3uvIgRMUx
oG1kEHcCGXBXpkK1CIDjlrLT4K5iZh94VZJ238pH5IN9y9oypuWFHU7ZVHOMwfWM
yMO82Ec8WgOIFKV/O0bKIllKAwf0AEYcr9bsDixh5jqm9KLr/MphNJlwH+5Tbexd
M4uZDXYjBvxPYidmpC2N4KPj/g5KywHGM5kh5g8NPU7/sYln2Wru+yewLPdzY2mv
T6WU9ClZ4JhFxoal1PcZz7X9Vy3DvddUZhWf4lkk6ieOWDtHLntA+VnbMi+1KJDy
kvm+2OJJOClX8azcZIIUPQ2c3tb/Rpm8Ykl6SHXGuMSDmbFIM3vXXG/GT/s064MK
Rs9YnBHJsPAPnIeCiv12rBJ43hyJP6Y+Fl2Z3PNCvcAamIWvVjlGludPNSeku2bi
jshxGByZtSzCr08A4MyFKf0kmk2zdVN04J12XM7/fmrSqJmw+fdiKWFcVf9tigoL
qw/xB0UKgrun3I86LwB+Qg/yKcnBspkkNiRsHhOup3TfL6202NBFcSMZ7C7uqWtG
RegNXP5dyDpLpIMOCeRJkT3vIjx8Yn1NmPoxnD1aqBZa59GAbJzyl3tVjaoCGf1y
wsW0IF6BtBFwV62iRebIWrrTWpADmpmmiHVrxLLvBnsxPOwHofQFBhwKISE0XXBe
xIS0+vjFzVqpasxwgGjRNYvv1yiTDVvmJzVnOFmKY1BWsPCXLP+8EIFp5h/I0rCF
gQX0N88wTvzSV7xJI9OJxop9L9DNnwDx5KuxgWEViuD1yI61GcFnTNw1wWcftLWT
VcX2XTURlVv8sRJC+eSAPKd+HF1kJO4BsRBx9Zc4VLowAixLv2Ec+yTfNpTnl0/z
HWZizD94Uuwra8Pzmqp8AcEBvtfGNlKMwk7TwrbNf6EsgeJ6eMHX93Mj7q8Zlwy0
BVjVmwDNClDKKKemkV71v02WS3cB2vW2kI7VsFdmNt+GbpGtZ96LE4Bi6utM6nLG
QMnWDbAeEFhrEe5lZrM/Gko8b2F+3e8d4D6IIqdAGnSDuPONKW80cPX8x1bnFzk4
3jUYxXxqy9e9ejrpJj2dorLS8W6QoqUC9guzgGXWoW5UMgfp4xltYEay09WcW+8i
/675dV4l/NzqX3taxAc50tbcgVuGo4KdIdtebdhxUgbAsRg1ttSdxQa476ugyIjQ
AZ61VAqVSBDJjkh1JfUr2rb6a3Xe99/MnqKoa1Xt+pSLuF6RrnQy3LGXKl5W9bS+
JhB1xhNJK/NPo4XjuAp1Kh7eaAz5BhcU3grlbC7PzAnAcXxL2qZ1SSMDxIl8HHkY
i+AzoQ408GNxAAFv3ihXrgDiX7ug8B29E4vrH05SLV/WRLY85WUBUDlQaeHHY+dZ
QDf/G33m4JfXsqld/Vi9MRMTRcHwwgMzJjoeKy0Dv6qJ4kJGS12UYsUvUTjDrOg+
I8MWZsx9K6toEIKTaxXm9fMkAUZgaDGXtvla3NiOY37cx91gd6Oyn3PqBFvyPUn2
GAirRxp/2d208icrXY106d0Kc4Ak6lOLpntGfSLqzWiy3/cXrH7juS0/Mg9txnRy
jtU4CAH196k7KPYc9riQMOJ0Nss3zUkU5DslVIsnauuT9Q3yYS/ogDHNVdylnvni
U7ajzMy1ap3hsejPpJta+ktw8q573clPQ9kZd8aS0ohgtdaYYWryVeCxjDXGnfW/
XWw4BzjxvXSeqbajCf2bAjfbYkuB5w+qCilpE4H0NjkluIMOUdu4CKrkxHeRn/hp
BB0eBkHatyLhAnDJYIDcpPzh4obcTkolhHKtWT1F5hPg0fHE3zcp/lsB0LZmluVT
my5aZM7XjgMd8eCKikCD9wPYw/zK8uAKLqKgho84bUtkYxZGo4vwn4OVw/X8qi72
plFHpZH5LkC9gbStJ51YymASxhL6kuwBlUrk+H8LbKTVt762F4U1ri5nzuiPHuK5
XjgyAss1UL3NPwUD51xtB4hnXt9M+fDQcsLrp4VkpLSsHMHxBwVZHoKH5wisRzdW
SrF20Jn0i4XD4oYH40YSFkW15q31DxzqN2Z5CD95Lt1/4avnIossgYfiFnVBRv0b
9oridszybd2Pv+fmW/INei8MivLM2/+03MZBlY7ip+wTNYo2nYezBjsVypBC6tzO
tMM+3xqemh6BLXSzzv2Q23TsQddyQOEx0vMfqRpGkZ4m1/1JVCOkpP1g5fqUMygX
eiwxp5C3l/mQs2nEatjzo9PRSSCznPkBqyJ84+xOKIA3WEft6I+Vu/n0DIc6np0X
ul0vEXsh5uOSqIFdZGZrH7Heh/ld3bFWw8xqh5ar9bejsYKu/BNrh9hRjl5pciwx
bb3SXmSStG8cNgK4UZrx9hfx3NQ6UGReAxXXhEJgDGnbbfLigA2vA0TlJoL3pSMH
YBF3/LaI1lDMuhjCiTWEV3T+fhycjWVfpHMinAaFQE7tGSAjam52ZoGRHN2NkTqU
MTk37SjPUmKYB35MScrup7LecclKhBMviFTpptSkUWNmSHc+2QbfAs9051Q3Nv9s
OpSfIIPsduqlNzrmBHlfDMPLVqNJa2vktzPfB4CIMIsewMmSUun1lOmHda+i2Jlt
pqJ2v+nB082FBZXE9K86nqGOGa+zh0rz/wU/uzmOEvpSGOEFLrYo1i+Gyx/nxSR/
zJhcVoNEKMwkhfkHpVCmj/p+EWG/2BKzLw6fLsHqXkStrRwJS66uqUAjqkKWOPZk
Fgihw2S08wUEpEcGVVBBOrYLCOiyolqnmz2v4FJOQJO77lvArnKPBkHrJLWx1WC3
Y97g5s7nmkrdqzDVLw/o5lvrrtNnR/kMdoGqtFYO/xWN2E030/L0cZEjQnGwZzvZ
axL6onRA3HRIsJDnSrIwP4cmqtWvFmERhIH2Db34tnbtVzxQGOYL+b7n6lhqy8HV
a4AzyT7mfRgElbiBGzvr5YIKn4Cj3mEFy+PZ/y+B/IBkheWYuLS81mVTc1SNxlxZ
JyP35EB38D+VzGCs8u/GyAulyCtkjVPbPcdOFSE7KUMx7LU+QiPyFuymc6EXekED
W/Nu0bW0f2KJSZaLFkOPtSYwLWyle09pqmYHlIipJIMQ90IbZwVigIPfUus2dkVR
kaOp9Wh5MymrYisFxXSl8bHkhJ28KDYo/xLOW8iYpGbBduA2R8A8YNqFEqOpMGB1
Qarwmi22fBGoJgmV/YJygrBnmZLKG2MXbMNwfulW9jHmkUW+XTKzG7hvYKhAm88m
V0LslA4J5bzT5oX2+rmIIdycczqIV4GEcqw0ejzqoRzx4FYxNTM1DT1Fd5IL8Dxj
9xC0GKF1HWx8hIOUFgIS2/1ADpx71DZyJ8JL14odlcbkpKYHD/E0wAIspB3SVi23
BZmlaQ2ZPDamAn9VBHV88HiA0X4qayrk6KJQeTVpEgMhDZErCEeSXDZY7cNQ9dhf
agLQseqDTL15SARU1cWgGRIDk3Z24658PZd7RNDwaUat276xgQfnUfTxFWCJ/vSP
UuVUo0WEDxb1KN/MYwdcPaEzrw515AfW/gsEuLNth7McIyuGPYKF7dkydRZNxOx4
MQbxi/9pCt1Git1y1l90C9QfeQHmqmzE9Gfw1nz80okdsBbvvjD61K8V+WnzLC3J
LxI/ecnAsWucOEOtZ89nHWijfq3370DyQvXOkWeRp23SkAVn8Rzk03FymEIsl1v0
mvia1og8qXaYV+XPFIdUc72mwagCUEIjC12Ru6gbPdWT/GOvLIS2AwOC9Su+vFAd
2ozs1DoVn/LOOAufIGAWyj4TprbEHiet9Ba7e4W5UTSlrYSp70ECYysTqXb9ts1B
xBa6eOEVq3qrtbNJPQzphoC4ndo8xTUNVCH4ZIvWGGdd7TGh2aQa/tscnq/x+F7e
QTzZkagEk3w3YoYkAVHFLTuVRnu6cBQQsLoU5FLOcqeL0QV5+IUUStPt6ukoeCts
yR+6M59VL/mq7FSpmFavQuBwCcZ4qKRXvrxYjA3Hnd6QlVkeaN5puwxTXhZRsR9T
RtjfuV8bbI8iWAadUBTX6CttE1no9noLXAhArsw3gzn3K98I0tqBCJUXhRcc4Bgn
epImKU1ggFZFj4fh8iL8bhBuuNcJqmSJ1NmXp3J+VVhwldzWID/ClsU84BPAL/Ui
kDpiypmyvX9jzZx2eh//3MxIZ7QOG0xilyDzJY9W5q2HtqTI9NQ7+wYfG7CTYGlD
gWlurMQB907OhevZzGR8/n14tSupwy1UW8m2SQz6ZmUYfNLJmRowCLTsgs0SBYE4
XKEVPOxiaeL6O8DFpdunFNNAqcJ7Tif3FUx67nA547AUPK3WlzkPnZcO61IOGDBs
Hoz4Qy2kxqOj2EMbIVXGum5NzqfgkUASD9BoFDZ3FPufAruOr83t4PwSpFfG4erG
7uzbPJdaMzxOBgaFYvOsQZAM/fNhbHLdd/+ovWm2ziqLHaNyrRU98vfilCodMhGj
nVLNRgUv8GZKOnpRbFDjW9RhBMt4S6nB+Ye+5DqiR/pdHGAgNv12JzzOFmpeiTNk
J4/inarFSeZXHLYf5LwjD75boIgcF0EiiZZrw7KzRDCgA+rT3hCgtb3R2Fv2yBV3
webxX50Ga2faHROxKSAw9pLtxwwHQMtTGhqmI2CsUyvim1MuwiiF2FhPte3u+8f3
RddQsZb8NMoMpEa1D+gmCMAyAjVR+d4yr/6B8EfGr2Gru6PvBl5pDqquuimZHe7B
FWMP8/6HL/dLaecu4I0ik0sJLpDWRtFnz6RNFxBqFOZkgbBbLWgb+5XDdDjCADhq
8mlGhQ328JLgjkz6e8oAq0ZvmzBeKqOG7sPxjqqj7oRtYzpmqLeEcJ/GeYP6WNW4
v84bFKmdaARYUHCNeVU4y2QCRCrA65byq/tFhMAIVt7/9q9nz1acImxtw0meagun
AN5ccA5Pj8Gn1u4CeJN/d0/wejjLGidayCp2+E4ebVhZhw1C+XbqWiTnJBHgSmqF
v5t49rIuMO+G79cB7fpmiz/z9fJGTMYnm+rVlub6hhVjSkOWrbz6fz97FM+ejnjj
7ZqI6imBIxnPq0A0eE4SzwFgneTBrKJjCYwvPSbEzLtc413aIBSlZOi6hmITo8Ai
H0vz82f6w8UeKpBR7GEtpoQr0CRkdqGsHbFKiYI3MI2MQobtZ4rpw8gXT9eMS1R+
yolH21x9QAfzBc6hCkLa2QO7e7Hg+JyKtS1rypOpFW2KBlGA8uTxmOvQkENLkmle
jeoktWODLHTNpU1KGNIqm2QtKBjtswvS1JdPmFVDtLloZq1dDGlwqaeAXJWvCorB
v+fGK3f2fI25uZd8A5IUWaz35pXbqV8klD+bvDKuI8H6g9x6voDvo50xrRKnoFiQ
APj3MJrQwVdlOdX2jJSy1XjroxFVyRAqL0YalRuzpLPQnWZT3MLk2Gdf3ETkiT9r
igqkHIyZMYhCqgvXj7Exi2AZsFV1zHTch5wxwlSdXs0ccqufRxFhEUUl87EhIhGt
KBtDgW/7wBYfLhKWd/tml87IJfpWm4uRDKtZ3vj+U0MJUP8GSZpYQjPqAcKrVVEZ
yk58tAeimj+Ga6+LpisCTRRwbP1GZqhRgnhOJebYk4W6b7EjFu3AME2zHhTB4ZWo
U/4n7+Q7mKREetU+ds5hUsA6Wd6r6f602PtjvjQvnCOoN2wVjBnMQ0UdbqHr+ai2
JegVgvkHHx0KCULpV1w86byJ2YKmac9vWrstTRJIoEgCdPkr9U/+EXwEZqTL+60B
0CxIgWssAuPPC9ryuxG1tKGTz2dkGveqmxLHd3wpef7AT5KcM81Cdr0T2PGOZUB2
ylYYsOv13peWKzIKwgcLkHlyTka60oke4iOBE3095eqBgWX3mpoc1S30wDIiGShL
kv3ZbvMeTBKa8Tar/+2xksIpaVVBTpcDt4P3yKFFX3btTRrqwNP9pkWcXUt4gczc
kKSwA0+Jigob9HbKfz9kLK01hWaFmTJx3z9WpWD8CNAWkcns4KsufME+2wYuHbRO
J0MW8q3be9OUBggA+CS7M8lQZxYi0lfPuhNJEnnxqGnu3Igdhgj5R9qnAhqUHZ9f
c5uG3WaZ0dJal0d7BOtq+5XwArrIbxp4TolcyZvfXtoocZbvGBDck9StwY/jRuMD
beQkiS6xEorKX5Zb+PKutcg6cW1ysxmK9GrRvrYh129vVH5NcYSnJkHChGKUnIjm
XvQFOzbmosWGHbFqx21wd1ifwQ/3hFWjjmS2+e2Nfldg/4Y2CGMD6QtOdUO4mC5v
u4FzIpy5wHP0m3aCbgkSU8lvkMDT2QR21+08vjTexATIh33VQkRhV0+iLe5ZBXwC
yGDcbQUSW6O6pAXiaFoXyVo86LCHI62+3k9fIkqpqfVYvaUnQdoHr50hgJziJ2UG
OpK7WxAegWDNbPHiSjVR3q1WSomBOWoqVFk7+UIM550xNDDnpJ+xJaUyDO0aog0h
g5D6puqifIrJ+1Ala27HCmf2KngHTAH8iLyi/MkR/xaNkg6RHYa6KuRZJqfekUpJ
o/XvTzgB6g1dgBxQQn3EJlVjYPEXizqzcPwRAAt/5ZiM4WfJRDvMSKsJ17UUlenb
vbFeeIbfK1vVOCp9ZH7mNziI/VzU4kl2NHtYuN9OZ6wBsKLDkFEHBSdH9SBt1arP
KAcLHrZS/P3mfv540xzQP1hgEYg5ZaiMYmhengoyMc7lAWKee42AJShTEcw9a3xA
llFZka2jswzz6FB+ThF615U5W9wASmcPWzQ63xMdcDQRj3vRSUgRblSvgbUjvVVh
GoIC44ZolK0h5mlBFksDN8RgplpnmGDH+Dt9F3Nzlvqk0/cyxPd0gN1WXarMGpra
uMHvJs/k7w55xVFF965LU19P5yg6shUuw2m9kSQ8/YDgaI4ngYTIklbVZCstHtkB
yup4wkmWsb6PVWb4lh1LQWnATmKqUDAvrl1elC7gYix302WZtDO/h52UN/lREbsP
6IgMOFIeRX3a111Qdts8gRmsm6Pxx7fnoEGDmSDGsc4FjjIQlwnYKDLXkB3IfOfs
gLH/2TamCrN5ad9jnJmJfQflZNHNL8T3v8jyh2mCxoxfyVSDFsj+q+D9YrbWo3KZ
z7XK9JAlrqrlUvlf614VAzqDq/FNXRX605Zd5jFZbZDe6EWAtBMvnqA/OHZVFEBB
d2pNDgsXECnGoNqGoMJk4niKSJPdrZnr9LULd/8XnSue0Pqe2KNM5Zd9BS7b81Cv
9Zk5Nnr8tUGb0pgByCy8JpoVNQzBaXiYFeTuurdN1e6Va/Xr47A+ptrHJNLn/Muv
fgg1nVqV7iIccOE0/DBHrPjrlq1KnveLb5IepDlP2Ns7TVue95v4e+ufS15dIryV
BmK12yi62oSafJBAzFU2HoA33YvtsYjuhPf6ZYu1v6rp12+u8vSKqkK+Ql2pT7QY
YyWpr5LQBQogy8Iheryjuxfrqpuoxql90Sqa2W+gcYHhnO4qMP/6IXiI7FgsmPlH
fJsjoG86JshLU3iEaNnrB3YB7dWksVIVC7q4Xq1L6pokE4h5XanMz4VS/LMKSc2c
uEXFGQJZefKuUeoZPjBArDiaFrXmbLNBdjTEN063ZY6+aoZjd1wpkON7DgDY+YR1
TKgf/JpjNAzEjzxIwx/WNKhAPT/da1QMgo7ups0uVuSYktL85mHxVHlrFToEnbdg
caasL4tzuTLQ6dzds/HnXgKSq+Jm9uhQeE+B65NFCz4t5empx448WOaltODWco3G
ryij8sIC4s4vyeGDPDQlWA+0dmgya4wqcor+N+OLfiLMnfMzDZasPtGV/wKeDlOx
UJoz2D6PN0OwdOKqswRQxY5YXYGJlJ2lnE2ptIxkqOFJwdAu4qJLJdejz17bn6yO
KCqZR6cbIQe83Zn9JV89KT7U1l9zRuCjWgeF44Y3TH0UTCoepu/0Cw4P3iWzo7B6
4btDFCL+B1vVuoSscEo5Bi29KbxRmasKR49Y+Hk9ttxP3h3RyDDOwxV25nJSn30d
OGE0Y92zeCsUT6M98K0ayZiuJytq/YnFPiQD7Iu2bM/t+l/sWb/9PjL2P0vvpCOJ
p8j63/MmGcTuLtPNupNX/UhbsOMqhKlZDL1j6snQ+Te6cO1itTCoI9xZ5o9B1UsQ
p8flj7OnbbEP4K71RVepp0YFaC4+8Ii4xiE7ZNF3SlsZgNqqux2JclEt3H7k8AF7
oPVjmDjzb5wLGB0j3Q/ktHdr73Mxyag3tIwpbh6OBq4U5fZSzAakdDMMag1UDQOl
vW908QGLqFiG4zSwzCeUXYaazosfvyrQkQdALsxQMIjeF91Ups3JB5Tpkf0yd8Vp
evDV1YBLDBDCI3gC5mV2G/xgUpffs7KjQySkPY6M6GM5ZDsN8LWdRBQO4eRn10q6
kKpZkTB93oTfDFiYtV81OewASOxcmuv8C3nI4d/TLXd+XlSNlLGFtVsuiwQi0Q9Z
ox7lEA3RouKsE5zEH9phBTGM40fcJzx41RuFLjf8RQjs8CFWdwdnK8k/AeKrdh8r
u60KlryhBs+f7X759tRc3pOBzmmHkwQLPshl7odUIsT0akK79unDh/Se7mFLRog0
1npSZQJr0veTVJS4YPU73OQW8bBfFZRCHyQYQaL7/+Hq8Evz6Dc6SnY6dtNwhBsI
zIkwUJSygRZ0ntx17TKSQik+Gdjm0G0jL9FOZdM0fmTmF8N9ga9M8XSuR9sKjaW+
OuqPG18T5FdsTxPVrCg75JBHEG0Mopo0dEf50b3f1FaEuFz6gKJdzLud3jOXlFOv
IYMJGHsPH3gjP1eR9iXmkuZP1R4eoNE5gxKie3x2sM3bUQ7SEXm2QXVfE0niX+Pk
PKQPLP09tPR2WOEaplXYPgffrFEe/ZP1S/mkOJ/bU8IL9fF5j2wasXcejJ8dvgvR
Z+Zzq7DT1IYvfGNDDLRabURCAzbXBqyGRMwi2XbWec/5+mSnsKKAQzm0so8Yo6lT
nSRP2Pnnk11b+Tp75419g9EsAQWVYcOPHEqUAJAxuZZsFTc56AFk4pq7m/s9AZpN
/MyuksQb28yGqmXJfD8oZmF2VNqhYzuGJGH/GZEzIwUoQSB1EXQ3J07cF96ccVTU
gL4ybHaCD7QJqPhfMYidRPIDdZqpnGCG5Hryw5vMPKssUTGO7eTEMOcs/e7gTHwH
6BkheX6p5SRrBkoY4o/memG1j86AobLkNk0xJODTmm4vfufaDm4rOgKS07N4boh7
5su1XkDuy3zXPUv7Pk/eJst4+nDlq/zbzuZFEtDfXkNhJBDW20H4w5jojaGxeXn1
vQYVOmwT3xvA0+MJGRKH67HtFOgCUnr8Jt3q8oOJUHH/S1r/fgjanFhGOWo2PPj4
3goP1A9kYH6QE3bdzVjY3FIN/dIh2hTA5w6m90Ubcw/BGe8fIGZhUvPMaFs5pZgs
Yugdwry60jIH3HTs0Oa5ZxUXw8bo7MObrdqjZsoFvd7iIbT4gcP9H66zhIEKbEQP
msEPdKHRex+k2SDR71+ipojyYQtiGLdsN1L15M8BP6lN2g3DEoAUP9WRgnq5RJ3U
2Vdv4YBHsRVQ2OfciJ5jD0Bp9f+h/DsdAWaWoAGnWGHXB5REkncFzL1Z9ONCyR4H
0k+kkmcsZ0rYFYxC7mGMV8Mky5E1mnOLBYcfRbqlT5dJpjAKAWaRhaF09AeGoovz
lCACBeiZfENxLxsarEEuuXr+8rMz61ZgcYQ+/vhmB+lM2UXQsTcnPUFVd8vQ1FbG
dTC+G0LH2eyi91EEmtzHCPkgOQENSzltVlaUGFEYUneh1rTxsaO0dtC6cMEzXsTA
X8C42qF9mql0wMueUHkocLO/T/e/x5UIuzUbUY/mKY5fJt2VpxuFcpp355c8Tl0w
UcsNc5Y2tY+pfj4r4qZeT3hjOQ9YE91htK1UiTkuRGK7w96GhAhVDvV2JYP1WtLj
NWnXJoUnWJukLZSeB2V6FxnMlreyy5zcNAAVXyJaTZGQfaKVvByOzn1ltyjXcVZ/
WYl+69kFJaw1wlOx2301a3bkUux96+q+xG8uh/7MH5WprUWahd5AiGTaXUs/mDZR
x7f1VPEXjWa6I5xamrxEx49TkqUMV6prdh00h+JRyNJvaP1OR+KgiffBHfztOUoo
DdoxBufU3vl/um7GL6ROKvDYSiS/oBsxughPOPOvnzgumOGdIiXdmWtUPuGx75mC
tamgL5CgyFCeTBOWIwkO0O4+7BKigQ74RemjgGekivAyelc+0nUCFCpA0A3pcz5d
tKrPvBz0FhuC4+DUXSIG80P/vd7y2rsUZ3dQ4rzVHdAPfCtfY5lJbutX4O0iM2Us
ivitfmqPNEzRPCDqEsKSIOQ/S4HQaymhLklx9c6ljQu6r2dFlaoPVDj8DCK8XtAP
saoYYiqvsB35cfaMlPIrT21giD4cz1x/JDVPva4D2fUwE9MpLdt/GC7ATJtE5jd1
1+aFNqP98pZVQNelXRRHaD5z6BO5J7OeZattYVTTBvd2mpYbiCjrcHu0pvv30nIH
kim+g+DSvqEXHzzqRuc0Hy0u43OsU+G9U49kdGnEnbWPQjXh7IQoXjfKgzc0/ul3
hsNUsuH1aI+dW9+Mhdsq1NwhozqlCbynAy54GxCRaI9yXZ0ITSdzruD6EjzNJoRO
4hrhoBMbf5w9SbilQAy0PTaaU24VEJBKqBZujNmCmIIA+Ax/l42umIa1JZ/I9QYY
RKycgPyD++5t4cHXGzb4sUUGJhnVNS+xRnb5ufiM1mQm6GogdT3Wtq7O2S97Bo/z
ld6zAgwk0dnGG8eByNQQ33uM/qCZV5eMzURMTsTqgQQvnUWkID1e0uq+LblutY3G
CeOsE/QNgU3OXWupJBV3S9nVRCc/xs+p0PurMJeaYb6abJAw6BPaLtDlsgy24QQ9
gnqniItFQI2NGq+CTPowRCFwF6Dy/4GfR7O4VHYqB+W8kHWY8tVo7NSP4+kl4cCM
UcP0OAg7oVpa1uXE+H8kI4c3TI657XZtoZNpmPpOxg9IaW+CaDVyZhxaVemYHrbf
XsImqVJP4tBWBDaiZ/E7LGm9g/dYmz3OSexIm8nUnc12sGx9S/cGXb5HV9vfUqBH
PZ2VbCDEAEWVcpGv+AHxRh4GDkt12kHMy2+P8dRc8av6aqx40Do1av7GBDsvRR47
o46Hp3eLpySQYJ3G5FPotAQIVP2ufNedSE0wvMl9vKlcyo0jaO/+ToysXzw2+zFX
z2Bb9ApcaevlEk1plwLh7G0HZfHepaqhDlyiuWEQpJBvx3axR4onm1hOjH/b1K7J
FExDMapsak80SxfZwpMTIor8wekvNvqvdNMm+a6Lzb1/1RiSgvjFPhobOwrR+8Rj
uBN0PES5su3ybBz022MBBiYSJweWVp4shvLZnJRkrj4IJhUARFuYxmGj8kkMd9q9
7FbBaCZV3KhALorEXT8EK+oo5HYVgAtFjc98a/LIrlwaGfrrz8JUBu0cH/iPzGie
kP/vSvQeI7iC+LVJnqCiESH94vQloig4AUEYmDG4RbOQ3xMzXNWVmS7jDdv1s0q5
N7PfVpSy4dwYr6RiyPlfCeTIvkiImGj4gHXA5VkTDX9AEoB4w5jjPKQLfsuR/wbk
8l4gKkFboKG4fK4Fopzs78K5HtYR9Bz4qfzX0Lr8bihh4beNBSokmoQF361d2eWB
MhSPzJgvCxaTiV+HrGgq/2RKZldx41A8jBEuY8pmxRfuP/adNJnv2O5NT94yrteY
2/Qm1D42B9LbhT5AmGq3JJGPTrWMZCTJT5RmXNj5CTvMM/GfDhwmXISe+3AJrgcn
93XYKiNs1IiB3H0cCk4AuNbT0KS6LOUGmlxSQz76/StMpa4TpaXz3NzwzOZ+3fUU
7MQju97DFeqTyOHuGPGpojqamUww6jTNCPOuqDM2yDUapTsHOoX61gsUuNDLe7sd
4qOeexYcxK8rtnjIlNcoPCunPBN3TwrIDxmzngZjTAGJJCwVqirVEBc/qPFsRwxJ
PRmphum5s4UL1dSUtcnd8GOJG3JcOSC8K3ubXkoPMryeCGZ4JcNv6s9evHd1TqTV
zTshXoKredpzv/A3mvmvAsBMHDu4ynCkYmPS1v7aBpT40N7dqnJlwFOJ+ULjp02H
WlUzNOmXvx9XilC2cDU9roVt2kO6SMIrwJwObHzakJ7yN8Gluqy2HQt0E3XT6RRf
Rxx+4Z+05Y23n++enKZwLuSDhHG4t9acRaaUmuXWzxGRscNLP8wS7a+R6q/49ayE
mjr8ild86zQ/WXRtFYD1GJhzbnEbJQzGypzNhx2JxL2Dd/ael4GLM2SpZIcs2ui9
TvMMdloCnZnXKaKYB9B98pktr0qI1D94EXW9zDIrP978wK+rerRs2mFXMmkLZheF
+hvSM4C01ShxD9B6xviF0cbt8wUs/AGnPOtn9Low49y9Ix/0LLOfVzLvuTHXorjv
Mym5XBgxbA/kPrYw/RrdfW8islWy8oSxiU7PLL4Dn5myDq8VzEvomeMeRCJ7RcS1
wKgQaeEs7DjmHNaLG6Pxj/7E6CnR0xOv8DI2Mo2H6pHrjDgAih3OLrJPNWsk3ekM
H8q2IfDPR+bA9grmDTKPcPkefXx0h9EnT9C5TSTtY3Kr+Ct0trx/QjwFAijMyKzh
rpEB+2ShJnv/smAeySQyaQZGRo1h/YlDQuZjfTdl87zLZaQThRhlLhqIOtbPA5FE
XO+5HPQ0Lhn3pXtIFjepPqmaUeQlm+3LuXR904/CPe6IN5CrSvxMsXGUEy1907rL
oTlYkjn+z7mu21hPopeh9XasxJkRW/Sz2/sqW8aSoZ2GwhxYEgKCRkIzGH5KO56l
iYe9py94AHHI8o/82kiHiltGD8C+R2JtMyPFxQRba12atYaK4MQ5ityY4bDZf+Gd
L5s4bmSEXz0LNFj84HLupRlDxvi9vm1y/DZZax8UUxSW05ABkefh0crkDZOmv5eu
IHGwNG63mt9jHLf93EjMSfdRPMayBOF1y2BTWVls3VrLK6tbiATK/v0+aShPRUyx
n8Nvo3BpY4ZbDSRRX5JE8s406tRZ4x2p51tfTfGtWb7jV5l7c/1/HOrXDaenapSn
0WE5dIBRWp4A9Vg6pCc934KkjlDXXSAYc4IqITe61HMc0zDCR1uvp6+CW7d5ZxF+
bdhnUI8nGL2dVlZIVHb2ZKWQyO5rTST67KM/Zl9dxWvfrJLR97E4Ekyd9/FpKDEv
65xBo/H9lS/RYFm/yCNTPVLNDoyA2WKmjPTkJmZrXh5uqelp3xQnJKhe+1n9rdEM
9tECyoeL43uhxhQ3VCTbMvWZrrcXsScMqDz7yDzUBtGRHNnWHpp+SpBTQPC+Cef6
Oudi2QQSDqdFb5e8hojMvHDPszVm4nh4oEv9ovmO7sPbqkPDBOlqA6BC0WJ/VNgK
K/M+pJziPRArQaRkwsr5ws7Bohr1F2ES3rYSFmYMIj83e0ACBw9LmJtHOy2AYqft
y/KkJqzzVWgtiTSBVCFBU2SPy4uTSuaRpHEQSKlutOTmM6H8CP+mGie0gvLATQ4s
UL4M+fSlFJNBrPMguWYbsY7PKN7cXaBDQMBgwqkS1AAV6riO7buD64fjhEAnSlA3
nIXvKQrwaatFHn6ogF7utxKGCANIKBtWr9zqvIKHroEWDSf4/zEADVp96tjUYeZp
RwZNt0lcc+EYOlyAiAyHc/iWCY3uYA5Q1UeGcwscNkWvl4V9ZjHboScgG/m+30lU
EVA6Tbyb5V4TBKLHeTDo7JfkD8IpHCntjKbhruDQry1sE09uPwK/t2qSzDExa6Xe
qbrwQK/6ZsvwytUxJcuHGmuB+WVSBz8BThClPLKg4BB1itiq4VfURsq1gnPBqT38
902OPF9QzZ4ooVfE8fRwDeTYCz1MWx1IrfbD84agDBhXjBo9HxIepNI9RkxwYbHo
7Bss620ZmBLy9aPjb94/INSmKHe6UQfo2yCPMAvt/jfJtsr1AlGDgrDHBof+Aei7
v845K3m0nMdWqsLiTdKtva7wRDwZbGGeWEGUBhyU59Q/I59+7k6Q06D/N9fI+wqB
v/5xmt7yDdduZhTmWugYBrZtA0CFMuS7gLOb1gmxyI4EAgN+RgXOAtjt/eRz7Shr
kmqEUFk4yL1wN6lnhThk/KS2/UM/VY3cTHK/Bx0Sz0w2/k1RrTN+fmKFWQjpc4+q
+iPhz8+xS+npABhHJH4BpeFvc8CCx9/GZqJvrCj9T+6Is/AvFHiqSsQIBFkIEMkt
4Gby/VfQ70n18wbZdBUUVW+MioRxNrXlPlFBSst8GCLmuqzC7zzHI3u1GiwjQDTj
Pg3z1LO774TV72rwVs7llFoM/ZgiD/fjYOzchYVWCVoB/TFtaDZ7dJ0dHoliINXk
PjaNeIYH5X4SQqU0QL4wiO5RdTbkC9zTukWi5v6c7QLv/ZwJTwK2K1h34Dl5qx6C
7vCfvOSDNHP5nnGKUAwLTgfOdjGyiZ6e/e+XouYVt4Zy3igyVTubdamCQ7zDM82d
FVXr/mT3ua1fdKk28FlwHsC1xEYx+JjDAdTXDnP/1rSg1MHd24dENYzSLkT7VI9W
9tI45c0fU7tXxwyWFjdfNx8NUt7XWpbPu112H7qL9mZae0jcopLnF9YoM8sx7Z/H
fxDRFyPt+np5oXI9dERtq5w2aEuocfXNn4Eb5nbtvfexADxVNfu0sZC+2eDQfJyh
xqFTT43FYC9uh1txAtE7pU+63c5gDBLom2UOgj9QAghh2Le38sVE7H6DpnQVLC7P
2BDQ+l7gtzyn7/cQBz9aonSRqzAQLsiRIxPFKSW8SRl601gP4He2jmz0s1QJ+MRo
zkKbYaTdAHYzghpe6/1iUkxBGTSal5Cnw1RdTP296B9orE7o0zOg70iIYMQMmku8
XKHXNX5EU591W0686ZiHqBO0828ZTiTNoGF/5OZAIxgljOTOn4uqaBXt3WtQ0zdH
9DnMfgWJarEcPmcFONQmWjtcRoagIkmVHLFudtnmAjs2CcJFVPmUlHcMVv2EJjy9
MTM6lycwK3ayCXbm74tbv74MqkZkUljwVElBl3rwmRnT9CK8xl7BAH7aG3epdlcZ
KTPk5bamWgZRofZnDSdKTm3W+lsvjySkyI30c4D0tSwIMP019vHWAQ2fEjzsZzbp
EOqo6tOJRESl8FZnIAO7SVOj9zZWN645XzGltXiwbMM10qRL1HZ+hJtlmK+X0yby
TGKS6yZjo45FwtuBB6frb4B5bGmzH664ffak1TLiDk1qFLagmhUS3Bg8RCw/Sq12
RPV6mkiRxBvGNsqaYVzqRs6Br83Bo/qCpzifZf4oretx9qXBMixsDyea5mjzEEv2
sBV+oTfgq6m4LBPJrefUIIJyexgNvfcnFYIXmaxdaXmPcfz0R/Rxc6Q7UwZBYMOr
DIGor17GVJyPwSR4FoHm3oN0RYsal3VBGXg3v4isTJK7Gi51WM4MS74l6xvLg8or
xvusRtw3tfIezujorvcaw1q0ADmk2SzavZEtU12O4hzh652FUi1YEEXBbXjplwYY
fewSQBXjPi/+rIm0CZ1Gj1pIWMslA3WPtKnlzIKIBmCnCz8vHtkPtE2nxYZ3nME5
s5RqrAfqynewUfc5dvs6dmLLOD1KrdhAJmOgJaY3LIHeY3Plr7tb0WfGdDAV56xq
JnWjOO8mnXutmmyGk7N0AK7yEFpkjj61bs59EvqDtyoMI/m5NSBemB7oD7Z6Bflm
rC7vhgt1myUxTGjpVUVzhcM40qTjD1pIgzRB41HpSLs8jg/nYWaji9pEGUtds/NB
OB6ZLIaoNh35qnHa7FOe5ru1KAdCH6QJmV7EC4CuH3bvoLR74/fwkyKnfb/4+lDm
vYGfmZqSTiIEbcHR0HfDSDuEN2Sg/P3GuzOt65HGW1eZqQZ9UsbzBngewd2OIX8q
yqAGiXI5ciS3KKdWNzbzjjl/M+SfYJadGWnwlEWXTP+iwzrYXnJlp0aNk/h4E3cP
zpEW8cJ/qZDWFulfNcuu/xLJpCspMtGb0q7t1IMldiHgBFfFiON8kwhCyZpHpQ1s
tUpAy7abQJFmMI3cvCWy2SKJq4nNouJ27mYt5rTtWNKpxa2DPLM0bbPdoC96Jgez
9kTEboMUxSDZAfWXsQkuFgSP9LhPIREyl/3Je9RafzrdFz7FZXwSBHvf5AAul7PC
L4q1o1URRIQ4E5iVFuTpvDTCyHKUtaiAiwsUMF1EHZ73A/HLfAcsbT65HqV/qpS/
HkdMnD3ZIdS8x6UcR8PLMDBVFtRmMMXyHhkAIG+zR/GTHS6cMVZpuPVHKTHAYOyJ
vyyxLo4BuIPMcDzoqz8yVELOSuuAZrP65uGW8T8pvEF6eVG6OkG6y4eCKfgkNQXS
gGsja8e+SwxBs3GIU39kRuK4dViz/t7lU5H9BlcjHcRkfGiODOf2B8OHRaeYrX1n
/qhGEjpw4tKfVdR/NhH9z7nOoUM3rFfkNcyAvmyx1XkB53YHnJvM5KM2NQYrMhs8
fFLp6mLxjhNB6i5rZAJ6XeZLaQxjWgUoVc7oVHRyir6P1YJKBegKuRa0+4j267IP
0wQ/EjWdC9J7zvCbgQBVhh6kTPSugMysPcvz3M7Dzhji+bi30G3rzcm+fs8Too+A
/7FgtoyB/VQIF8l1h/chVtfsRno6UO6AHMTLho5DlVIY/3QcIhhlq/c4CN6UHFWE
hFvnxIUox3fdH9mLT9JewYdrl6qVRqnUpW4cgmUYr8jtWmUjRcebFmFReWUTUHhg
QQU/IekcMrrA4k4xPErXz4NqmSKxj+iKGT0B79E+7gYmdqdwkBSKF3VicfXoorda
XewCRC4v24dKG2WC7GgdqLIVhyhZtIUvdynqy7RQlDW7skWnW411287SJNT5WvWu
nXtNygu5o1CaLOHEZaSOEzKJCigQqbGEOkLU8BVoVE4HX13GrPFnXAo4nnAzWe7Q
nIunNVLpgDWKRGXGHi9Fa/V7M53gh9gaWW2Cy71qNU6O/tEMvGn9/0kqN3wtwqtG
TngFi3U0eJilvN9qv1z3WOWNZwTvtikmDffXnFGtz7Ed+5x2KhhHkUtXd06+Xnb7
l+twH+EGb32/OrZTZUVNTaniTORKARjptkvm71vdyVPJF3EeKu6MqyMoMuv6EHhe
erxpgXWh0rXCsbRwbii33KmNTVEYY3yWkghfmGFJI4/wyxHND+bssKAvXTHVjpgV
lAEFY0thgwlbI8Y3pfsMfQEkiDHyswguig5gH8S5S4FVbZm3PGhbiegGuwFzgvNX
YNt0x7fnD72v4LLLBGV3BVoo6G7soUha9K0IWr48x95TmtGDN2lJqIT+I3zzijY8
pPqQVxwcnAnCvmeGW3JixlOSvaDSHXiaTBLLDCfHOuzMfcxK5mP6Nd5S6Cc4FTFm
FO7K8i5BODt/FwdNV5rZkz/gMD9Tzw83VKPR1ccG2p701lQnPfkJOGN2YMBhm8rH
2RmIwRYzv8iFL8+OZyQKaYWxg7CN/iU+5LzHcaTKQ8bFkEvZ84TC5u0pd66xW23o
X6BnGM2kx0HSm5+tVZ8VGZxMk3yZ784S6JUFJzQd/06/bchMzBQEp9K7Pb7k6BaY
FIwHtBPecylUIurTYZaf8tuPnR0CqgscJGzeX3p0hjUr++ZrHJO3UBoR5asyLaH6
yzGxXsH6Q3Ljs/UP8BddeTe1jxB8gIoZwMfuT8r9Yqfd+V+9KDK6tx1Vif/Afo6P
wGeeTQAuSTbroE/kIh5ztUruej+bD3oqvKWm73GPdJzF9K5FqeitxHnA3twx2wq1
XF0RwGCA9d2qEOA0EtUkxJFtja4MMZS5+sMWvo5GHFpfFV9oe7BMEab9/7iywLHj
XJzgasqgdnqJLLbzNtnVrjhPDbO88mpy5L0vtbt1AI+eL961HTBNkBHUPl4yEqRz
f9T+zMWreIFTWoCMlrKHgGEoWDrVOeYBkobapADHAM1q0JnG61XQ+zKp8ZP1N7E/
LTjp3a3TYjWW4e4q7Fh4nnKgPLxduhvvAoS9C82GBhx2rrw6VYKz3Zn3Bk63OeRd
VRk01YorksVnbQJ6I1/ISEtvjSZv0L4ia/GvlJfh1mbRIh+7iAFL1+CTRxHSGnOs
demhtEGRcDy6WvXZYvP1gCUW4tHIWIsi3VcQYIYxLRrzjBnetqD10w9WxbbWxTDx
C/G2+2hkQAuOxohYTfBIRs4NDbd2NRqd8+NrdvsCvVxMy2iaq5vfW1EeWql0sjm/
x9sXNzBEll/U26e+6MSDdIZDBb6vkT5f+YHdxzTdVoXc0zAkKoK1xBItG563eMQG
Lbi4EJjYZlV/gedYuPTWDPxlv1U2ifPc86Q7kL7xIqrvWIUuw7TVjXgwROh4X7No
XMrgcZVuEABsQbKdf41NMwbm/lem/NBCf6PodGEBbJ195P6meaTPp/aBT1mwH9Hf
4GqlJ8P7gnHZNyiKaGpA7YdhpZWKYVhBUNy2ZjKfXcVG6dRjNvAfSff+O08tGQ39
Ym2yiG1zPklfrXwX5dYKiLxlQrgiutu/YUUDDXoFtDUgVJEMEYyOkJg0Lw/t0Bc9
SObjFi0WTMUDotGGak6X4YLKkVaXuHwNo7r3xDCPZPqh4Z156G72xlhwoSPi3z0X
ns8mwFJsiNsfNY1CBo57kR32exyFPFRbyXmxyhOhDSWWesrDuohzEHi9xBMXdam3
29biYhoABx7/B/LQHdtTQz+lw5f7jkCwJMoihJqUJt9lLkg3zRAaQeYrh06acUWP
Kj8muKRtSDIDBubRCW2OzFsQ5MNyfCWa2l0MgdWfRpljKN0x4LpZnLgsH+aVCS1E
PgksZ96Wcd7yx96bigX8+rCxWI25/hXpVBfd16lwyRe6yxEvrqrngt/dU4gjqh4g
u/hWtWZUkyye1UrVBnRE4WzUq6tgp8FRxdajZtlnlZh2qJbSB9nFIGDfHPWNDJW7
4v7Gl8fbULAef8dl2Kx6ZxVNB6Fq8M9JLxlFYkqls7pVSzkZWHT3fgGnrBAXDTOL
33CGgdzPN5+wBnj2iTDcAQVB950kuzB6z3oHretY5MapfAc57rRkmTUZpBhiOu1v
Fm1E3r+lbzAXzamEbE3y7S/XU3xY1NBL1sFpfn3QOHZfmuhNQshHnrktin91pxkO
Te16blMMlRkj7rmjIoT0RGG3+/lNm/Dm3qNCOhjPbakkx2JhahE+BQcrq+QUYIXM
dC07biyQN3yHqrf7urRAjPGAkk9Jy3jrA97HnSXioBcea6RLA1Y0r9Ccluh5w1vn
2JuqO5sQmLGJfSemN039TplYbDOv3P+r6S539kbN/Zv5YMUlLpWjkvzDVHcbXVCk
3dlQygTFZaYlztjQ9qP3PW21idjPWfU0ZTd9cuff3BNPvbe3jR7ntV8nKhXkGGD8
QKwiNo8IxkL7cJtLZjXz3BsRhQxnJNbvETz+2zxGgE7QFDyJyyJP0JbmfVZux8oS
v5Ag4Rc3FZaN4INEHrpewAjJO5c5yR1j9R0Euc/D2vexDcD//0QDyRyB0fJqVaia
ICknLL3/K8zYgPJvtheiVxvcnZvkZDaEXqJC/WHpXL1REXdNe8Q6pqvYxH8VFujW
oNjH9t8bVe1SN5U89/uuxjul7h+6lpIlJs8ETFMvEAB2mxoe1WommlaHvOYS+Tx0
D6YNuoKfja2GzFO12+wNmcXDRpQxX4Bppg6SQM/O4DJ6+hQSjiKJ+ZBKOxlvN6sW
L0WNUi5ZoK76ohrjwYmhdRPuOh9xtD5C96+bz3pW4KkP3xIoeGX7pN1qSRnLyaMM
i+CBfcjKB0l19ma7QOnnBLjeClUqZrmQNZBUu1bCGbBGeM6fgzvSA+Gzi7wVal9g
sznM7FBAuW22VeBiuyZCWX4Fazw7sy4XveGdXW5F+/lUPb4S/wr0fuo7v3Hb2Ls6
zlbpGCFB0Nho2J2FmzO3H0I2cOHuxAECfzA+1Kwva4cxp3x9DVJcNHkRRhuf4ZmU
ibvsaEjwvmsyD31xEk3nGtocuMbiBz2hLi6h/kYMazuvWGd/ry8pn/1+0+9dlt8b
Xmd+DIyhmx2kxKS8Uc0WRur6zsgFqltAC8uaDBX6QoPVfy9fvj7R96PSoiPrTqud
9gTq3FW22P/IKBkkvprkuMJvbXQzKTA3DiU1ygjvlJ3URyMhxLqhkCBYUQ923BDJ
iSXakD+ZLIMqjXh0HpBl3Q+aPF3a1QOTkitJlMy/SnaV2BPUermObdJaZFyhkeE+
H+ZwQ6XJjjVyBw0bWSlrksvUhXEHN6qexjGF+eaVbSqQTyIJEuwgqbFi88Lkd4s5
JAvC99yxfC33VxUJU2tJnWnMtV65jf290LOfddmajOgPJYzlbHthQByWJDAjaxBU
B2qFfupCRtcoMFxshwzqPthWDg5Wk1vUi9QrqvzSRcO6zCV5pQzrD9Z0/S/iIUAz
8WmwvdZVgrAGUuBmFeuI4VyxLYPw9DM2gM5FOGGp0APiJUlU3mWh4RhlrD1Lq/KY
l0kwbxf4iJqPxDMNE+7oaALJe9/+YJJTF14QBleH+E57rS6SO7aa8WujOQIonPdJ
4Xb7tFwBJh/zJ95j9Yv+WY9Rl1fIyaeUxGFZRwA4xzlOwmVPUNVOP27sq5FwBVK+
2zlF6z51VO1vlsD9UmQ8Hku9wTe4uXUXrJLoYpnyE9tDaoOtR/tB26PIOJRJTn9D
sv9f2f2loYYPFhE8MPGAlY/JTNmYX/KUBE2PqQMosCWs1x72Ea676VmBarOMJrWE
P4wLDwAeqAkD5dwVLjJCF9klqSAucU7pBWM3zMWfeq+O2Obc1OQf97UNQgZHgQTb
5mSXf2TKnLLdztoMJCnV6s9CoD3ti2yV4BBB3WdYrkzJCjf6y70hsAIdeVTZ8dpV
pYIOoDEy4dFBUHNOGXJZxloqhDHYmKnOhrl7BfdP3qPjsfiMXhy/pib689J8OU0Y
BLqgKfDYP2Xc5gX47vI0+1P9S/p7S/ZSWr2KMZtEubXaiMXRYQBOrJkSFupEDyyP
LQbNs8u1R9u3SCvp+x7IZURWAgVJW0M13I7XSjd9J/SZZTeqQ+sKG3Uf+QMCbGRn
ZAaeKjreMtI7x/Nm0bOLpfDVpBitAAz/gXP0nR+JabYrTnpsAuWnxdcxDrm4WdUY
fp99vl2lmUhqnzDQ9jaoy+JZB1V0MBL0jP21iV8Cx+yX1MtfBwGhDVsAOdYo+vQQ
dn9GCg6/aUYYvxUj6NT9eXOICKonpwRPl1ZkXAarlrrBoQiPLlPo/kSl6hc0Cnef
HJkP7uv6FxQpMSGaW5pzT3vZs/K0Wcsb5Hecm7oTPR+cVbj2gb3QFLlNc6fhraH5
Vr1fI6V0Q2jvXbLUPpdASG1fkGBx36fQXEF0ZdHElKJOeYe6Ar32TSyoh2EtVFRE
FvOsEGouGD90g3GE84SNhp9Ur5nsG1WkcrTssFC1yseN8RlZNvGM2KuSJ/b7GOd1
BQm1yDWSVrManxZRXX0AfAq7dRuE27ONwymEdN9HbiUBwQT+hvvC7ce2MttTVoNR
cPsqnMK6s/C+oiVg25QwcVFc8nHWbYbUC9nOeVjHUwgrwyl+uzbzjiHwVEtqq7nT
tcmBl2AmW9GyRHdHd8ELIlyyCqV8xeOh+fq+ouDwBBRPf2n00cCCoz9krmNzqN8C
rVuuwkpfvAppoFKjHB+fo6z1KPOdqZWddHPzUiNIgvyFoBHpJvobHfm8oxZoQbyx
1kAdjVLztC9Cp8afrPmnmFOwQadR552XjBz7R9LUoJo2/YO23iJdrYBaChv5nwa1
EgJ+hf6OEUM4BM5dSAa/Rz996ofDpS6NajBUvm7C73tBF7KoIC+t3mg5j97akeRF
mbVyo/Q5TXGLee0GdsQILyL38rpGIx0PYIZlGiceffE9wbB/1XMNePwzcrIHak24
4mfxJO9NrJFFYOGJV+WU1sN9dfsTGO/NgVNIEIl3HO89mUpdKPvmwes42PYoILPA
JXHsYK4LsZGowG4h/8m2KZuudfQ1s4ca745tjrj5aFUpD+Vcwbu7TxpCY8F8oIGP
k72uQr/HAvYhPqpyEhrrubPN+7wFEpurD/uLmkOeKYF4vhBNcRsdsD4fYwmEmCEd
DrDjN/x/mnIgnbJanm2BSMU19GYsqWQbX/wHiIC13ciW0rZcN5DyOnaNxnHYASaN
6v0Gp86WPfgSa7GljMpCPSTM7DIgCywJ2xssWJLad2hdcJMeFqXe5+ffIGcMFxqU
tEH+WOI7b+8GLhlDM5PXhIEZSSWU2u9VK8Unrn1DTl0Da+ODAbhSrUBcNsLDrEd8
o6O/+ENPq7f1Wv1euOvZ4yXQEF5ocJ11qiWAdaHM6+SZpSnqsBLnXSxMcU0cIzUv
M8B/ZptgjJK4T0UVTe2jnLMYpo7f5jgQEptPgES4KAMt80TF2nN1vGrQleo4SJUu
dEZrAHLHGWg6wd66w9ahhu2CguNCz2hmmtSI3re3+aDM8o3n7LKhYxlptLBlEbrC
GsxW7L4CVyHhri+yquqkRq1fSlSS4+cLb28xaSidVzIhYxoHvHLKH7qbEcTO07JG
fOMH/3wfM+W6bvMxtP4/h1DYeKgbn+wmeb2Or1K8NqDH8HoX3gDeTDVETV+sdzMy
x8SxWDThv5Sd1NB6hoytIXN9pwwD8NnTC5vmW3Rq8n0ozcdc6AkKo1yuebEG7ugR
VfPOTrljyCmBX5N8jS3wRDtVUT/gz7+kd1bH2g3Fj5tycm7hIxijFcOd9yvVqaw4
QY/iR6u0ZD/Wby6/fqwOVpKDWG3+2d6tIIs7x7Jix7n9yA02tCMGSjXWhi/L3oJH
uiyTAf7K9V51phITLTG9YUKe0SgL5Lvn/ryS1O07JPiJIo4QBLZf0m/eF1hLPLjy
G9xZKYaVAZNt+R5CPny6zVap81zMRTvxGKMwk2UkLYUbklQEX0EQlXB4dEgJEy/H
8Wo27aAarpBj/R/wZDoJFJvfL1/AjCsDP3FOnC3XjNf+cE16TTZaJS0F9qhHxajA
hI8EgoAr/WmGaRYLHYTB4wfYLuP9p/mn95xKP8coHdWo0l8sjfJWVXviR2l9sTb+
yZOEf51v0/RJSLCpMj5GEGQIZfmKaQOQRhjb0k1164mI1TeBrHYYLlLeLbDcEbjr
3cARwTBe9sNkRZRHGJp9KMPYQ0+ITba1UbkEwMnTRx+S5DNH1V1aNYoYpdk2rX76
1H2HwbI/mBZO4eVipme5Ab+7keGIUpNqYFw9SDeQ2W12c6vUFUFXOERJEEJ+BTj+
HXDx9x0kEWEZq3/Ntz5B4Jw6qSM2vA08OwgIQRgqI0CTBtU2iENr+pBhwqoNUf7S
VqTjUQfYSpdH3iVb3u5xb4A/MKEdFxXwPaTMcV3kmAYtQ4r3pQYb4rYg56BDqgEE
g04z4veAT21LhdTErb6cdEG7bNAVkd+mxT/wBaW7tolhFgB6eUzgQjpjEv+A8/ab
2SLA1izgCUYt3SteQyXAF9t4j4BOPXVBqKpZmMhoR6NklLPVuVC4YfYBoQG6G2e3
q2DEdVnQx8UcbaudaoJKkPxozJ/et6qjA1+eMnf+ZY4WxHfqjEOQTApUL9QLaWr+
9IwnPtwNy3QCSJhmigJdKk5+f/CApLczsv1NI8s5gkd+30ZImofYHYLE8q9qy2ij
6CWNjtm2WqP6ZEOgE8Mm+aOydvp/dOrREGRiWUO/U9Sw5+6m1TqO5rwSNqZIq93u
QixVXMRMC7Q+E5J7Dv0n7MrgY9SdmSFyUBgdQDLiocLjGap1GwIo7jgT0CwWDSkt
mK149X4LlXY4fPZ8fIuvOL/CihwyHvs+dC4039+17iNXu2ZyvrGS83R54+tBMChx
W5++GereVN8xC7FbTqVw5xQjRIuxkm8tMn7bbgANi3ZQQ3KdRskXjqrKoparS6MN
cM6YGi1ZUq3TcKp4YkeSUB3Ws94qAsV495PnZSA2N1zbpZEs9c/NvyrCX87jogtu
DvjVmfCU8Hl5YKoH6XgvRZrbroWs8lK/vbQceLs/Jl+OGUKKndFZJQvDVZ7jHC4C
FZGGtZQU2JGYgcFoAVaAffcv2ruQr8u5LDZqBjqVmGbXj4iDvtiemWsGqFNY7cEc
5rdW/Bgv6cyqo912pdGQlRu22jZA4hXvYZFO6Y2iLWuq1EubuUV4Q5anBbF0DW3q
0QksmC7tIRlvGzRskleViBcJrsuMZ7REBCIhs1xuxwe5oF1FrTBlE0VFIN02T4RN
VAhJmFmYPc4k6g7fWaG+poA3X2/KhkKZPjzbfR1ksALckxMbcNibOhLgpfbgrmqK
+kBAqaw7Dbpz9LnxfGlRyW9ctsB4Mcxgof9OMgYSGhndd/ryXEmC9PmqsuhLKDg7
ADbhwhebLf2DV/aBr6paJX1poXCFL6dolGGLuzVHW9Fd331V22GWj06SIX+39jZ7
hISK/uw3IKEUJ2lUYBq7/oPfYA0HaSOeU98BnFTawfETqNbvi0I1KJE39bdW6x3O
bllA0AARWrSyRrteFXnTGQ213vof0juGbpqLJXtT09dXUm5KSUAz4HOfVPom/wOt
6s7+nlxWwpA0NbzUdd7z6ReWehI1w516J2/t9dZHFUr1OM/n6oo+Nj3XQf/s0G6x
TImCntLgcvK2nwc/6Ff3XwFKM8uaXsat0X5rChJTnn/wCK7vYXOOnE098CqSp9GW
tzfPo0dMwte4bS3PBTe0+kZ7tJswk4QczB98ci6n9QNm3dL2x8rEAZo4ohJ/b57O
uZdttPKQrrlp9CoeubuZMEhdUn/HFaiXp0W31t4x+a8LJsZBYCANmCXthFkM2LhJ
CVdcevVOU7RSnLSF21fJtxV+uMk8zjoatDaAJFiBorsWf0109OTJeLxvRH+CPOLR
GuoTdSlYwFDIxoFnh60rndONOsZY8Z/DJuKChdZl22nJDgNqkspzPTRF2d/umQBE
NIAfSdISeJCrCzTsf3imUaU0LjAtj4KZStiHSxVNrYBwM20df3WFMUnXpbXLqBXW
+uNrQWu8gFV3t7p4/HrksM7n6pfgp4KoAjY0CpgDGzip+UUUj/hDQbS+Ksob3S80
G1iMA7x/dK3pNTm9ts7l+gZL17yNau3Wcdvk5LrOj4jfiFTRTECZxSuOHp9ahYPO
INJlkm8uEfjeWNNa9COxgV/jguOdRhmRb6lzCSbwzvbWVNCxlxOw3hI6drQ4hgyF
AgGglJ3kFRcD508NEXC4Ur82zZnVSWVjPKZtJlnPhbyMz5DzBN+sKR6M08WoJGyE
rwarB87hRCXn+OInIK+Cn2D83XVTXxAKvx3a+FZyn9Df34A2g/bvbS9jlHaNMJ2C
Hrrj5HfbGrFM2cjVp6ZdPcX4XbGcJYXX28HLY69e6SGxUfwMi0LCCsBqdAzNjJUD
7DFmzGQUIwJlseUYPNcd80iPOHkZAVleomDf2+U/+0NSNqnqLxs0OBVqMWoIn/Dg
eFTj7QPPIaJ4B4qtlXcxxj7mgjZHuo+Jzo+pCHEVF/LbM0ZtCfSbjWKAsdTXzB7W
8mFb+aQJGx3jkV42D/oV9CAehFeWmRkrBK07y/6EYbsDsEkZsSYOuXHUUJCHQpBV
HaaTGrU3bZzo/GzhLgvEkGc0qm34a+GNDboK7ICPg3IWqihDmHKbt31MD14lvwa9
JPVv4krTtmvoIDoYDt9/W3ezmKcVeHuM+pLMPscjawKLwgV9zO36yLSzhR6qbJg0
0XGz9XEZWJ+jk+G/2NXxV1xdioMGgX9SYFdXZ7aHEqCFX/08roomRXXSjG7Jh8bh
o7f0z/xytJw0tTfVIQYBySx4Tk+DTvL4+KfCRXqx0n26RfrpPVDhOoAUQGs2a2Bc
FNc4dE/Dky17ptPyhYZ6Iqv1D2J+iuTTYvAimKxgXyZpJ+gNQHZ8/XmJ6tCyrhaU
zd4v7NVPckPXen/rAAF8SKGybOtmx0CJJaT+XzlQ0PYaYKG04ztK9t1eZQPpL/SU
UgP1mE6dyFM/d1A7DIkJXgqF7mUw1arhJiS7h0CZCQG93I3+va2glSAHmyYDQlBY
nFtj40hn3Ybs2QLXbF4rDBTGFe6qSx9sd2C4E/uTgI1AYuUmaF36AspkTTaQTeni
A5Zmu68YpzbyZil6eS8Gqxz1A8br1B3DqxqnscV9sx4puEcJhIbmjecm2PPpuUj4
aofb2YHibhdhdl/CflyHt1wlR7JS8H8me+bOKXTqJjj7X7UUFtXbWHnPYgf+sqZm
94irXmjn0YbY5o+4DelOk6a209cODX8ZdNkBGq8+ZKgcIS+ngGY6BjSftU/Q2Fay
JdeqOdmd5wSTlsuJtDeU4RH+DymSfpxciCdtXBQrjsFEfGdgOa5JVPw6upF7LWRJ
2+BBATNk39xyE7BJ2mNnq6fq8qXR72oVh9WQ5a0BpVgI8bUYBXv9hgBgGNE8XUfD
ZgorrAhJCwPPDoTEZvF49BvCeHA4z4ZgQElYv7x1egY9+JXd+2xW0PzdHxCQecj8
Dc8BggWYC4KLcl/OO1dCPpTYIeTcGzCJLMtE8NPsE4KQsS6zYlzdRE6w5U1Ze5R7
58SV81mYx8j7me10M9uv1xIWr1vwSpHBzuEFXosw5CLJBLuswDgchFNFxEtUluWD
2BNq3j5NKSl955M/1f68uS2FxE02pdBcuz2zWov+u9/NTEmu8HtScsfEGfeGfKIc
BwAMxaHLUKx4J+hyOAUdp7fOZ5EYr7EbfXho9Y5J+oMnO/w5iTEUpuxhrWd4Nl30
NjFWGxlW+M9hWW9C/nEAmhc2tEvx7YvTyilVJbSnt7H+8qNGv1uV3SBTQGGHHkp+
7fxUTO1IpLS73Y1J18aJ4SSRWles+JvsgBv6JD1qaJHpyzYYJxf1yLJuBPvgMoa8
Y4edVTTOgomtH3RudL4LFSPg8KDSZdLfhUbxN7snrhHQtJQBGwe1rLe8M1lv7Y+8
2QuY+0xC8svstUq7mSUWVkIcxpDXyWTpjo0Zt4uM6QnnxPPKsV2/8Tr5TqIaf5np
RPoieqsRCo8O7q4MFTJ3AX/WGAX3Cjc7n1ypztIp/H9VJpOX/BYbDjxGsxVypwOr
SpLmtcBZFVL5APwdOSkyMMIheoDFAxP/4Zuw5t5is897JqT+OOLt3XQ+3rVFNakF
sOkAl3v21i1yX7QuytCZBcaRZjanMX0I4fedvqXr+C1hVwNfBbr2X4LkrQflK7BW
z1S+JdBStLa+Xm16H9C9I1TQ3JEsl3HVyZsV4nx2b6uMIYfC4pQuXRSsdZqvZmf6
0XEVZKlxWuM0020Dxp9A8ibupi6a9GcEr78OFJ9Hu9yawC5fLjLByDUhrxUqAs5m
73s9msT2yBD+D2hQYpc++UtB4WmEuM46hfXqViOVPvUgdKiRlFQuz7/bUvZ1JKxv
Z1KIX+CdVa9V3SoK+0mW0YHdvyNiFrHCyqO/h8Hb297wG1EAHt9uRYJQ8vhNUnrl
d/o++eqe2TzJ/Q5CtvLXvwhtwqeaQJVYpcwtZSUkyag4rfQOuZbv9EDBBEKCQe+d
ENgKCghCbul2jFeA+VdkI2Z+VzC4/DliMZQPbHW4GjFRCQjX1MftMO7k/g4+Nfp3
M82E1delvbMukOm6yTYLfH23VfTVXkdNiVWd6+VKBzOQjXuNZBO1B71oQssdRj/O
2fAVbiyae/UPmtrHI0U+P/5+kRC9hOVLiV3R18YLevnZ8ERkrDGsl7AQm7mRYRem
Nt8fi6fcm4c5PNFH/S5d8ESlW/7Et5MFpcJq8TJxHH+ZIgsH2GpU61CB6h/Z55ht
920enKVmXKl9ym9U6X+eZ3dcG1l1cZi+g97FfEmotCheSwnZG0SmUEed8xmPGlyf
xXEVHzCJrsXthf8SL6Ge4/aGh0X4s5XDJ3RKXeReJLFGdM2OiU8kb8afNomMMovy
gKz1XF2X8InANK3M4HVWkHJSDL3olIAZlYW4S05+wLlTgkf4NDyOYoXBXCbOkfVP
DVdcq9290mRpnnyVlv5JS+vtt6URwnb1PS+NoM6suPtCi7wCQ/mpHVOCL2EzN4hE
QBkjlz0LAT2zEwmB5BDZHJWqAeK5HEgUQb47F9bx/5NDNjeLEYHphkqPw9EuMYzB
eIohgbG8GoGOKttPmZs9nR832V7WPyHxmEEVBXt52zcnGVRmk0mS22TCkkb6+X8X
Gye7mP5WelbTre5O74x+AQBi4jPJnh1Zr7ZMDBShVhbpWYgRnXXdinWOPLfzVfL3
c9VBw+S7rkP39iE8GZhNiqzBberH6sRDxwhqn44AQbqdZj94FqJVQmDPDV6MnYSj
WInZXYLB6lR1qXZa/jydQV+K0WOodpW4kNa8HvXwUgkHhEKDplG2q6mINhsYjg2v
LGZ4kjsItv6NPZ6k1YfN9YV4UkNfAPRmpOlnOn0mIiRmt0P3fUDGdwNwGA0vSMOu
KPLQvG7I5sr6l9ef0lbhMb+ayszeaPJJujww3o2TsnzDvwAnCyHwZAW/szcuqB5E
fLfxr7pR1GV1FatAooYk20gdVEHXZjrszf2XkIwog3mvnPTSEwmwLbmVTz8gejCd
Qpvm+IyEvjaMpFH3Jal/DiQiySgWDOf94VU5jUdwN+afeZj6BTty5wNlT8W7IplJ
BQBgz2Nb9D303w6Go+HPH6m1YBCqoZEFEDuSLSRxlLVQkl3o7EBU+v+u9dwfxvId
yLAz71BXBP0Zy2vPQcVmOxR2u/1KPM43K/vOzilfEl5gwLfhL4XB6BM2ju5SOMA1
hdUIpySlQX1+GH4c3SM1o5m8ret5FYkvDh2/MkkQNu7vRPTFRVmxoQZr3iE4hdTz
5C7zsnU0IMo8De3ltXoWNbVSh61rONKc87Bx1JK9usKBVXB3xW1sIuYjalr9uYho
pyBmN2q9Ro4xiN6lxymbo/iI0JkbFYwwEiv9UWuKTx+AwbRhkXQU97HSmHI2U9NZ
N98Nqku/MVnKrcjssjVHfzbnt1LIHz2txvzS3u5AQuZT+MOgYoPz3qGfHiu+1IeN
23/Ri0xRk9ZUVooZLYO+dCEhOOHOVbRGOyRY+qNTAkFpac0jcfMhBTj6QpM4Z0y8
AKnk+jfdq6KYPLLfgwXyHLa5HHjEZ8t6QWF5YY8Tbxlq2KMj/mUiFVROetMxRG3R
mH5rbrqJXTpnBPVMGLZ6hxqi28vzOsz6lLAviCLV2EhkVWjIDmLVAXk3b/x0G/Nh
1IK5hoaw5owlSgL244K+mbepacm2MI5k4+hsQwE7Gsk/KmXqCCFjQdVHLK8P1V6Z
gp8rfWyDgWKPJrYj8CFHM4U4Sn/kAphzNoeFJko4g9ka4HoIwjFrlcrEXdMaIUa7
LIghsdNoIsOR0ySiMBdj4assT57MkMJqteHWAbuP8UVod3o7SMQ3OJnlnqAHWFpF
C5a4ZF+addeqoOrnG6TpDNaKtQs94tI72lYV4JhyHm4Uq1GFVIz2A5jM688FfTiL
u1Xsd39mxiYqd/2iycy2wjBNgz9pI7S1sSERLdDLPKxcAKQAUB6VOtuYXB6N6COX
2XU95cMViSvEayqIHCRfXc5jir6vWDYcaDIWn68lIJDHdeDYtFNAH123JOR4wFnT
VEj2/29Uv3g3P+YSjh+WH697VWxDHGtEzWQDn7KvmsOPSHM2Db2ko8ch0R3I2vPo
uR+4Uz1QSLEDLWCLMJ5pAwDcyvYkAzdj20fWB8v4jr3jb+fuhZe7Z+g85zkD0IwS
RiOF0ZgvYEqRvTupFvva4VcxjLcAaDktVIfbo7YgiKPRxp5dD9FETV3/+vcZsOVI
cXJOxFyqDHCqylamNbEKAUPyqKSy3LJDWSkX6WUlW+rFRKKFBbnnGAhjfOqcIrLh
cM1cIbp+W1HHtOMRo/lnXrGDZxXZl1erVA4KyS/pJFdx+VPRFWkwLTCMgNy2dcx+
NmNl+z99Usj7cUeOIjFEV/wa7RX6iooze+SKcO0HpSI3XCi4RMRkGNDA+XwRzThu
vzoGrKok+Jk8HKeOGfOHfFH5d7ySuhLJx+KO0YVY0r9Oov5yBm5sYcAP3mjewrID
nl3F5djNZ/WUJu6zmjD281o/XrXpyePXKiR4zC6OAG0ufA06KUVfmy8UtdOHX9R2
Tdp16vwWw73pYlRSbTGc3+BVY3om1T2ED6Rp1cCVOti+UNrpfi6vVdWDKbixiqb5
8reqM6jhoUAqlYAtbz9VgsXg4StLRKUpY9mD32OvUevZFeoXeV9ECyZU+9T+rpNh
DQL502t9N/3MIkvtdfyJvL++bc+umJp1FKqchMNzHeadThQBxFpa60qPib8WruAZ
tbMgU/OWLZAaZhCow8dxLrVqZe2OW1BZ0g4yMj6okU1wSXipP2/bXYgHmpF06zKo
gnzz1vUZhH1SKhwwiB2cWWz5zatJQw3OLyPPUfWXyBD3gWyeFg655kCWwY800dmg
e8LswGwbTGcMhkvUGrgxhYEMiULYaHDcwHzy7SOVphL40lDSlcc1wKy9hq1v8uZD
fJldUG79ENstH5BRLbYiValNETjQ2NoA4Ct5LbuNH7iM9kQnZEwN7mLOtfMUCUE+
gyGkxSNArDXAzT5v7iV0y9edWql6IFyq0JwlsvpNdCqOL5JRzIeuYXqpBMzdVywr
UcWwr0DpibK2I21EKExrcUT9LhoXplHOGfSdfmZTZBq6p+TvLPwJAKUKP3W7fkVY
ZS1rAjwW/cKH/GyxPuj8q2EmJc5ckuldCjtYbWQwk0JAfg5phxooWnq4DItkNnPh
Wv4w/6OpLqjXnV4Ow6m+HfB67PPQsWgSvKDtwySptNKG8KJ7/v537veE5trsFqKE
U06Qf7JSflJditVEwvCujhgk9pxhXFsoxAZO4AYwY7UxRfbY3tEXODdIqAxwgH/e
VtnpxdjXLxtnzqCyBpyBuzsqDCuaqnxSEDLy24vhn5BYT3CslFuyFOkCcz5I+PAV
P5B6nkMeJtBBcwhhR6Dtq4DWzwN+UUPp8WTgcRSg2XESn2B/MHUelpD6wLEbp3M8
5uceOQ71MntajQZcXvgEgAvxruf3g+Jjrr2Q35Y8yWy3ELJYcl/MqnjYHRTejIyj
WGmY1czyuo74lXpDpqBNDmKBICbzzMJ+AKEWIwuxBSsexkGmTTJIsWjez2ADFB7m
mBuBEdplStvqvyoLHh8Z54dFt+Be8n+gK+En9uEvK/0kqTpvpK6y+fodd6BEoLcG
H10+m/MwulVC5PStWXjgoIoKz2deZWF9V5FNfO7+jN/nXyHlmFJdGVcVgn59OpiO
0jlsmPe1TeIJspQI1UMYwpIJ8FfQtyIwFYAry0HlHa6edcl5S8Hl7p1RoIpyhMQJ
91l+tqHmNuTX//E9ebMn2HhQXDfAp6vGQGq91zA1HhpKOzA97tQSIqVW9yDJ5Pr5
3/yMGRc6EbUjStcq2T2zAbO1lBLU5EipKyH2enEmj++kAth+L4vRzYu2fGfKj1+H
VYLMG7EI4s12jRx6izqdDJFR9ir1XLfeLzgJ+0DlzDoRnopNbDY7UWQtdHyAFzuN
SLuoYiymt7qcRtYD1gZXCmEoPDdu4LnB82Cj9q+XVUuIikjNqLRG22s+Nris5NRK
jPuD5Efcl69qXiYlNH0eM5oHay5OLdMCUvofH+dyByDyyzPDFRGYZwobuwKSPNCN
tpmkRQC1FF6k2IgGBU1szdpFxuyARb5GZnHhi56Oo0oIiDLXBupPzCRA/A4YSpE6
5ynEgKiaAzzgOAUdBcVW96EeteHr7MekoSzsUo11mqDZRl9/iGG4zv2fIE4hyGoB
pDUj0uMN4bL1dTqH0S7xBfZTh5iSIuIEzfh33xVI12nN/hMM9HbcF7jrqc+TtGRt
pwMnqKiCp5FsWF3hKg7Rt5plfFHslPdQ7oqyCKtDh7C58OjTarJlmsMWZB+prsJG
Vhu9KeUk7fgkLwHop4GLBflkId0Mbt1PTvvncKPBir99xvBx8zf4G6a0nHbqSd72
y8NsCRMJrCaVtS/okNSv0x6kB/Zvaxwlp66ZcJy5rNEA2XUQRkjvO52YT7bxylOY
uOqjtqpljtiAbNEjX1e0K3jEM4YmSvmR/1pkm3Bq6CDdeHsOP3/nT3zmuwENayVV
x2Lwwb42s6M9anUPFY61bROBqbfnKs42d9dCnkXNWPfEPUausg6x9+SiecryeZsY
T7UKWogWN9nPT1VXg1SDkscTjWjMe2/6iPG8Wp/JTElhX5reYpHQINpXcfH0QlDN
ffetJBTPPhX4qOSdp8KrgdUDCTTpSbl7lCCJPCxjzEmgBKqNYvHhl0s0QPrfhpsS
QQTFQ+aGRcwK+6rKGjftlyzhjjYVyTEq4pjjhdpqAHwvm3TsDFC3Zdy7z54dA/ob
OD/i6MoMy+6s9mHZrH8DAodX9Rdv0BEb5b+y0dLRtf1FyuumpCeY3cPojSDGKO/d
mtpDO/k41VJw2mHatLNRO5Y/FjFA1aOMDvQoDm/jrmLUjWhPsZzQLVokOO76sdWF
Rc+M+1467mhtw7BWqHkbMlK8n6w/wVln4ehrYvX588pvW4vbyBdoxoTcOvIVrHgX
cxtCKMbxkQ5H+rG1+3wCmoqQl2xdxjHEoK9IRea3UOeyWYrIrXDBiW6Ya5K2K6vK
iWRDtDuynEz/SNl3rqPfch2q+CXxciKGbswpMVvNLfnMJI2endnW0PtMUEt5SVO4
biSWWi7tgXIWU30DOTQwSr/WQZ8vRgNadoXxCc6I2wviKa7DBL9eJk9fvZnbTiZU
inyZqAi7SzzRER6ukOHDauVXM4xwSiIdXxPpp1k72qST2rsq5N4AdK+JbiHaxgXr
CEqNY+hCiFNdfn7K1p/iJ4ycOfeMwt+12q0a3D9DotiClMloHTQs95dGX9NdJ2eo
QqEtH5AOJzXe7VycubYtjL4VNPXAfBqtamV7PfIQfTx5hUBdCG+D8t82yiEByGA1
a0B0b0Jza/TX6dfOcuXue8gdOcEHWg4lyeNYBDtZqUlz6R5ASTAIsNPPHLGTeGti
5JGcProqIwhj4qYCGRSOL0YXCd7lmHX9BU+3NCev2x04z75Os8WlRBjkB4okK/Ya
Scsg2Db20NTCK/a8OY9diDaylDhBs5HXQYnpNhcQmVcUqWQXfAlXGCs04tKmIvsz
+eR5n3KDXkdYDHK1APlG5fEkAaFL3nJsoVAPqScN6A8rf4LFWecBhHoGXtosv+Gh
yOr/8Jc/MiSqlLnI4yZxlclHRSEvK7CiaL2HFEK1hT9SO04IavAcg4/kwJgCgu1N
PmPpIfZqyHrJjsuhsSvpnoTWyI7KTuWyoKAmFIfY4ZSRb9zuxDM52HM8AFuXCoeo
OOchM0mtOS+VhuIe2ey1HvloqgL2NkH5NB+xLmia4DAl84W1jwASg8ybRfC4j8zb
dZiYsI3qgORjORR6Ipun0263sIW6r7UAL13Eij9F/jSKWh/67IXdcqvQPUyMJUxq
EHkne7oItww6z8PEMYOM6BPcB/yniqsErDW8c0vgQpt378mGj+y8KHIyTvhjBz1j
4eojKjIFh5lXYpdXHylZ4ScfQlyeqrKbkPSe7azMGoN5B/AfhafcU3hPdHdhKyEY
LDjQQZ1UHZTTrQ/pPY49gA2M9sl/4X6JMrEVrY7k1f5WnilJmxkhaGkQU86iUkr2
qWR5z7MPxIQuxugkBrL7hVAe7vmuywB6teg/WOy+GkdN8bKl+uQYVl/xnIpgivYt
iq4L22G081BJkQrMPllD9xH9p4kpTqmuNsjLbf7RNZWggwLX1/JPlM8KBVjmX6Qq
Ck/Oqxpp3SuWZmsEqT2eweB87kLJwnRO71veUvs4fpmhp4JSEb0RfKrmbJi39xRJ
xSGQ831jo12w4ui0hjA48yhWbGd5rO9TcBii2bZEiQffSmhaFyDHisKE5fwpKGYv
UwCSRXzrXUOvbhVwV+sRHb2alIziw/PQp8PV90w1X+7Wt4rJtgYSPyck+BfQhd+q
VEcR2reLixKCDd7M3YcTDj8GupftTML7XfA9sQBDsvbXU22BWPs0/VF4506BFVSk
sQbFFUze+uMNaemQPmTejDDJRv0rLONLCTf4fQw5J7pxqU6BdnFbT6BJttxy89SB
hDAB5HKZcZUJ/alY5f21/MJfX6/S3AYWgVNva+a6p0cYHBulztJIW4nRuQlSTGP2
YdS21wWH/5N4u8mTEnxjIo7RraBjRFQ7ScY7vebNet2HvyGF54AiVEhtTkqYlMFf
wig55UEUTGentbR4a/I1j6OYHanPgXjpd0Bz2TTHFvjFAlOBs+ErjK0U5PFLr+7f
IUOPb7n7q9G56pHx0HORiTkYpmQRzngmuSGmdGr3hGIfYUbHDtuCqyfCTpmyVq8G
NH24GtO34qR5IDjA8TDD/BN3ZMz2KKX8Q8acy2fi1AZi2c3Iwp7F8F/cT7NJzxyc
nvu/3vTENFhc44N6YiwrFr9C3/HIQpnropxVpWIQ7YYa3Y0t60AY630KX8kZ6jEC
Hmn2BUJXuVol6xh9QPl7BJ2E3D1XPTTOGh2UlEAenQr9icJRo0AWKrIPI0RZKb5D
oxfsFtbJlJEUrlPMrFQmshNR/N56FlBVKC7rqmBFbNktZvdOb/9kZOTbIc8gp9D0
U8CD8jsbR0gzS0RQTlX2xpg3djPhov0PnUqjzLHwXLhaEcewxTvSJcn2MlMTUvGK
zqAbuUmOHpmGxusam27yYruh86v1UCCRKH1mHC56elK55VVStY9FWK5AILiN0Jal
dMpGmUfSKL1VohpgdOvvzfNUB3wBNCBrNpheCzmSPjp94FhF94PldSqzGL9ZGNR7
uPrFnJ07WFZ4f2jQ0P16sRod+Ishd46LMra3vZOBm7D5Q30saY27IBHLIK2gefZE
WIDIsxZPW1//2yjt82TKnDgf+4Qj+6NFBcMGHPAlQIYrpgvVJT3x8Iz6xv59HZjm
eS1vN5H2IE611lxFXucuAkBa6kkkv2dgLrAMg6mRrfWTylYdC6ZbBnOTKJjg5wV/
eK4HdPp5zCnw3JbYytm/Iv19stLx0sdwBSAjgy4hWN27nbbhso13GeN6w/o1Xiv3
LgEHJM4aHK8KcmsbNF8MzhHTMBphuYDVnUf+n6lAlD1QFAs9/ISFmkdEyvHflsk7
f1pmmJ3SjG9EeVK1ii+v6Ts7+xma61BuaMUCpGyYx1ISNRVsnenKB6BnJPEG5DvO
Mbygk5utTaqEzKLdF7RtldcEO/c953D40gCr3Y4pFmnSvGoKT4zQ+iCvzVsE6F0k
1vlSjOmPyt4J55rE/iZFihp8p/FUz+r5qLitp7y0fwvt5SZhr8TU0K98d6+/+EQl
6DSmCYBI4BefNo/o6pRMjVDrA12KX4drUo5/xY56neRBN/AS+j09+vBefHsIOCMb
4FuMIooqnh3TBzHAOhJv/3O9wDc6DBYMvkhQ0KaBbWOd7iV/GaD6pyyZ8iiaWjSt
oaxtLOp6Cn/1uSPijSlrj57UrlPXCTP6ct5S7ppV6GJbzdE8O8tmNs1jW5eNFPuJ
HbwXv+3TuQ2GHf+y52qygPBi+QA/ttq+HqeU/reY5z1lqgT6FEwGk/62Vpmemzqa
H11Jz4yy+ms7dJKIIfXA49aqKA4ScvZ8XPV/dq/uooYsYj4JTvhx9fsEFs6lvEqT
OBEB8Gh5QQ6MbOKhu91rhaLHK0p5RbtOYuMDA/gwj1+7RXpR5z8wS68UPbauRHCz
da4dgN3I5WhUVf32S72u4bpkzNS9oLwqPlPkcCniDrWgZ3j+r1bYo8gg6RNqXq+T
AMZgnw/AboJxZGrwbavsjrBx3fx7bZGhZON9+Xi6Qi3NBqW1l1SeRdlvJwgVLrKW
n9Pq9ZQDaFv6pIHmg8VZpoyvNqc5e6LQNd9/3T4OBgWpdZ2J8/eoSm0zG1WHsXU/
UGQ3ZA2cbWTG/au/HyJQKyZrfAhJeeSORyxT718qOIFqFK9WWkGH2CW6hIsiWpuo
G8XnMQXy4bCAfJ4bhtyWlqwaOyv3a8na/TfqSY3FI3ddnhBp0kmlnid6R329SYnQ
bjZhCYXLFnKQ23DWKTo68nzCjy1NVD5Z0pyr48AJxxuP8Xd4sndNn2COy4R1GA+t
7JE3RZ6wGj5DgAEvsz8ZqP3scKXoQq6fgL4RpvWwns+rPC60YnFpK99RnSFjJPsX
tlf8fp8XG4ODyj6/RAkscraju/vbj+st+jqpxou0GiXMRPBIsdzhuZ68L0VTjfJ8
xiSTGYJb2RqWlFk7PZDWVZhxjqsuanr+S86UYe7zrX99gw0/472QnRyacRbG9aTF
u528YvobsE3fuL3sLcqjJoMGd4YVgsh91+RLRJiZPMJ2oytxIYcoOE7WPQvSOrs+
51dwNEVtbZHXpUSwCkqMebqx7fFdvfma+5yrmURACkBNY4zSgPL1VoltfFyWMf7b
GgAE1p1szWDtznfnjR5PmJMZPQna74DBHej4R9JogUWRoICyG66FU6MBn6vUyVwf
fTdokzhgiTfYP0xYxOm4ymx70+M/WZ2W6tv5l836OGZ/cqRH/vJ58QqLS1D8hycE
W8hyntm5lFgfJYaL2fT1+I2i9xAwlHwGNXMgJ0Fm3H4Z3T8cYWTATvhQ6hdZmh1p
ZEhUaR9gK5XsuMXNjTgAfqRP+RCW0DlNvm/QbQ51IeNYqRBqQxqKrRHF8hOySRNf
Pd6KJnDTRgNqxsrmXnEkLnBaMaBuOd6xOvNr/9ItZ0Ggr0Hy8p7ZouXv3Q+MWl+K
paxvZ4meQ5Ffz/sjZndJqKtr9BP/XcVKLb0dYci580yco/mjtP5gT4KFLSx/FS52
2EXxlVjcYqDyUixpOTSble29A3vPT/6K+GGJBxSRIW/Jp06HgZ7jAiakWS1vfkzp
bQrFxu6unn0GgjDioChibCTUpEJwf2F9waXnxdEoJuuq6klRXkEfseHWW1SMuDUu
M398wTmVVj3RwLr6ZzHwpDFc5dGJyHfOi/Va76RPPGGaN2xiI1n19UAL3OuUJmAG
S8jKT5DwrBD6IdZHn2lIbD1Uctq1kmk7SvP8VKrPDEch4HanYhoy8yT41g6cVwzN
iFQTah1wSoQIbKwnhmDS4LGcNZ1fca7H/O9fuGKs/HGhJ50JAkYy1gV8m9M242vZ
Vr/bFUlyWiXMJAUao8pWO6uNS60gWNAf01TtgzpZFEPiPht+HW3+oeVzK4Uq/YTt
9MSNTPXD/RPAywJIyuthU68H4yBu/TVEkPbUdfC28T/vBI6gU/qQsQAM5+L1wdNN
Mpm8kyV0TxwohUxpCu4q98tyYe2wLdyIJ4eW4U347IoWNosHvNUegb1lEpI7XsJL
UPY4KVv/o934g33y9i8VayvkeVcxq7QjqxoPpJkrlIY8L3L3MqUnMqyHYWein+ZL
3eJ7C1KtoLoIypbhhcNnNCpFSY150If2Zgk5JuRz0E385rfUoSDz2SjSx1qb1E/i
NfqVXXaLL1fuWrrf9m4KZKZCZq5f4IwBn3pDbuCZDKbNdGjTDzKg5rmR120mpR+o
L64yOExTrb2cCEz1XnM3kSfzyH1bRdTT2Ccr+gP2SmIJx9NbDcUlyLOFDDZ8eDWm
G6VvJujy7BSjVvW1bNAuH13h6wg4/EwDMbFsjP7fATlNIzHAAj1QOrT+DrXUQhr4
nMeK3ipGODPk/X4gBmsO43MivHT/mMTcF05zbcDJr1bvQKoImQ6Ux85sXmNQyw4k
61bI0rCshnmmIc1YzjytLl5y4nlJPttjFvFNR95qbGqkFE4cOd4vxBcaWSrG1A9t
3J9ASlyJiFvWiVY8NrjEGcITD+sLXprIZYmvwRWgvXdE60PWiEKD4n4t/6zbtiyi
FUZMLoLSno9/lGX4spPYb/rwPFyK4W4cY9qjxcEHDPY88Ni3EJW7+XzIqRF/FsYy
GaL4jyFAdtMkHWdtdY88Zww3Bc+K0ynfREh/clkMnhDyy6MIc2AffyVFBAI8cQJk
Kl1R/yvQauxuvllvebGyfcegW4j/6zs6L2uvptwM+gUeqomh2vNuXdjML7BO9dj7
fPiXwqY4HttlrYgkt9iIjCT0sI8H4HgxmAY0BF72Ai1FzAg+BJdHTqeGs/g9JR2C
+Hu0N5gzmuHcDPFXZHsS8b6bSI3Avz1LrSTYQVpOXEKO+cz7vWCA9ji/YqpPmBtA
2rVBH7pgaO419hlDPQyF/m9SNS6pA0uHMh7foOjxRVskhQzbckkDgO579jtOgxAY
bEJlnSYnFIiZRWtMeOmmkMh0ZltmBgbK9mud4T4XpOzHgG2pR06NPDS8lW9Vu1j3
cNDdvTyAMIx1plRFCpPSOHzZBgeK2WIWtt/Z0Bh4qY+g63vVSRQm8Kj2UtnEcXKl
Bf/cIzwoFwGT6N9v6qOBN7DIiLx8idHDQts3KIuk4sh/1JzrNDJXrjjVY2usZ2rq
Ts33+wUrCZCV7J9VaJOB4F6pvuk0o+G2waXcXLk4CSR/9GOxtpvmiQt0cfJrgPeS
l2BQ04kOyKd1M/l8Xps83Q/vYxWsX4pYIy+fwuPCkwYPDeYRYZk7qQEazGmT+qz5
F5RwWpts/WJG5WahP0GzwFgwSNTmgB04cJ15kDH7sMEn+j7nCWMDDrduiK0I7oR5
AqWzODSUPYIxgKnikWsoV21PT9JdimpmZYmYLCSdyGpZCxqHsX62BoU8b0rs98D0
efMOOI29v4ggP+DsgCTJK6HHc3IueXnXtKb6hCDdjQPizpQ/mdN52P0a5vvEaU5E
8moCNUEnXR3o4ap+xyXFcbmVOyAMxCvwXXW65VfdkSV9QouIViIuehOK8Mp4Opj8
ko5SlreXLjPG+TZ5X7hSfbqe9wclZGuS4O9UzSIZlAS9JS1JaStF623+YPLITlJN
C033n1P8l2Ni2QMzkvQt0Hb/C45F72cDmMTZGHI0CTVOeGANF78FQQoHiIrEHzgr
QSU5IFUFyU0QGgVrif/ISCn6tQbyppns73Oce8zjPFV4gR3v/oLKDhr7LlA4UfpS
uP0qUKmFNZLHm/OU32QYOVBJ3Ee7kCKIbjFK5jAXp6HnK+pfTYNujW6k8SeeE6Wo
09vI6509DHUckRCjzZ/iOc0qqeP4WJPzELHNcLfZj6IFBnDdJBmRIPnARdDI5yjU
+Sqpun4iY7MsodMNCIN+u88vqRrpsovK7iiMmKkC+XtrY9RIuwG1HvVw5PNea20/
KMdJivROoJNnWwZywb7eT0W5pW0oXRrQMqXwTou//fe82i8qhnG2fn3hBmjAlBPS
vRDN/GgMBS//UDCR0UPv5SRyYVXpiNbcgolj9OYyM/2eUG8sPxcNpYEP0JbHOkkL
SlhX90bfUJgYmEZemnoPfAfFYe5FuNXj1uqYkfX0hwxBLHpYsAc/27YOh2LeLyls
2e0lNnbueA4Y+frtvGrWL4VniJ0SA6K2AA4FpAOkLbd2E2U8E+ssO4V7WB/ZPF2y
TiHtakP6Q7MBWLG1oP7z3QBi4qL5O5zHTbk0vsYv91zxHOMydY2cvekleweW1Dvd
oXjZv7wTgZc2qExmZnHac9CEy25lTs2G2xRo4MGf7/mFUubgDS57JambFtzOn88V
8yG3vAuMyl0z0gx/hj4oSQ1MPEXAuujKuKSU9a26sVtKfgTbqPBZ74ptk4GSVMV/
Kbjy7BcdngRIkjcZcde4aHL/xK55e0oVPZNbg92IP0COmd0yPdVBNdZTp6kU8NT7
QHa9Bhfu2N6+zQ1BcYSnYli1DuxJR3yB0PPnwzJOQ2l9a7rE/xpbtV4JeB+B9sVH
FwKkyr01p0kLcn1SZZKn39jITxqlEnWUUu2NUAa4SXiwJEFHkRQKw8CD1ZhUQDw2
Vu7fkTvH3t62aXPXWS/hdz2jfGxut94LiairBACk2fkrNEC6fHT8nRSMfBFM5Svx
Qr2EQcLs+XOejPAYZRket/4ixbteNcFfzZo9XuWZ1wPFm5YEnD+i9rDKj4IvJk5U
aA4myAlzTyAEMcoQhwFXZY0REyWyQBtjBZ88cxzIBI6O7uMEYsGPq6Me8ip1NeDS
uJNY6eD/c6u1p+PcLq6SZm39k7yD53CBVWHDhkYfcrpYHp5hXgnTgq8kL4yQqwbJ
UeB5RVQCTgIkXtKj4qhSykI8g8UwQ6jrca/qMVTrmSMFjHh+wbs3b5Zzu6Ve7hW7
sJm3wrmItaicwzoGeSEkfX8vRQacnPYMqau45UrhsGR4BqlC/gmqYN1Kj3lLR5nt
R/ZunnZeDHYpSHFhUi4+Yf5rOsizsYJisCoo02M+15EgZIqSAZjRpqhQD3cQjraF
J7ai+ctiiaLfMsLbT9An3kEZW9neo3ZMeeF2Xf9pTjntPy2via01hQWeic+pgCYL
wBzrUxMratv2fND8t278CkSYSnCAGdhkBzwpSA4ISVmgYlgXSBNFEo78GJBPThvt
MLaL2Podo4cFiY1ltJ78Tv4OERqviiB4AcHCqiaoZ4incmY8uebR2Sz1UqQKwsJ2
Nxmg6Q5ip/ubgGTDCPnTs8kTSc7Q9a8bYsJtzeDsmMxOWQYWcLmILwp51OGwAwEk
jfMPK0h/ZjZeYIFvOeRAfzZByP+33WQpa6fwKF8mt5Zhyv8qrNiFp7TzKWbBfriV
qe1B3Ha0rLyVdyDHu5fVLDo30FEMvo4XzXVolqGHSYD0j/BMDhJUW2TK2g6v4q8i
ODqwp0E3wBaDM6T9VKbsodM0scJuZXE7FioWvWoomEHIP001Tr+wyA8NEvCiZAyc
tCXXeUNn9+bEA/TPQpGtNVEPUz0OkMxNs7NnfChWLAaML3Sb8uT08iXMSViHgNqK
5SZUvVUkaW9ZlZQaU+pZmZvyqFvqhnUIuXoKJlcungymbXlQiN/caX/RR30ELGWt
RNqBSwyf6b9oDcsQIvhZE1Ce3iOGCaNhE5QGz2sPN3V8NzcPkp2xOYuF6PSe97dc
k9eJy5bMD89I9FpAjXldC5Dc4bpBcrcL0QsLo1DZFXZEUjCoMQaaC3zshDiBAdq/
4W+Pbma9ghcvf03IXrnWPxMEG2eRZIYp4aesvjxNrpBXPG7BKYhvapm0JXiSjkVb
Fzc1TGCgeju+gXToo+V3fAJT1eBXC9xopvP1cSdiXOyPusltKETQ+q9rDlZBbAzj
c3C9/7d4ZQyPv+zfg1VP62g2MZm/N+eoOZUEQlAF6aigGBJoxQssdazBaipwsKnQ
Hix+S4PA2zVByYpGKwpKKKdPhEPo0TkDBqWAa+2ZfUoT4ECK+NuO29MDj/gUeLlU
S0FKxd2HtaLp637swtYi8kZVGq70fpRIUFl46sjFPZljW8RhNxfhMJmgjc9Ro0Jg
82KRFocpKRbGhSnwJ6XqHP6it/MkBapv/9ZZy1/XKXjKM4bYjqCioWcGadulkAaJ
IMnFwriqwV9m89VRfMse88/PYEUsiUmocu0toppJUg5qGtUSyt3FlSPezzUT/zab
aOLQvkpDOpRzggOU4vSMSGty0EHWPPxzbvz6NzRpUoNzg5TmGsRScl+83IVYVRou
1ErPZ22P9HKHSHPVR+0NPvwgSQwaX38FJKSqmMDJu1fcud8oDfg3D1Twjw3h3evm
Ggr8U16xEbyqkRJrgiM5TzPXkcnyc3SRoRI0DEjuz1pbT3wexboamaRJlEOgc1Bk
Dr+KicNyXGsUCS5aCaKNcrf6pH+1k6l6yScrTeMDRzOeodBwiT1tukeHryGZqkpo
yzn+4r1WU8jXnEuWfqBxeNgxwaG2XShL8uuCRnlPjmqr1agMZlEXV/A+hcxq9qHk
T9OWE1Sl+BR55/B0vP1te58xBMis8xumbuVNoybNet48w0DJzOcSsyQFrCSOMHqf
3t6PZdCnRst2VFcWLKFlWS3fJ5rQ3p/A/H/on/5yWbqwFhPB7bayseRoywMs0bsD
+VcqvAyC2S3KUDVrYJVqC2BvUR3vM11pVEAck0cTRtnqH/mGE3AU6AgrMA4ExTsX
ONDYv7d/bXbvX8zuOTV8OlLf/Kj4BJ+GDflDzE5sFseyjJ7exLc3ZH13O+GB+fgl
M8tHsejv4s6K2vL/vc4en2IQpLpzYs3wYpxxYMNFq6hcRV+wUFhboB9AehmFP0L5
WBd7UJHWuGIzpo1tF7PCtqTrAWdTch27jWdgFYv49vcKKUUsDmgvZxVW6wxsktmQ
eVzhKDJOT4f+6P0rwhlW0S5esZCmNL8jpM6UpfzH4F74weim4Xqz+79y5IT5yObN
eglV/MAj66H2m8BOEgXvmE2y8KBs1gjr6xcGqoo95WyuvcjUnEgsoiCWnAJLNdqM
NVY/DOk5jaZO+9ioL4V/NQADFka5wMvIsXTnFUv6n88kYdRsaMdjfC3U4EqMTRFt
/F9NkFnPABvMy2ctBlBIVvauPf9gtLpJkVJw9qCZWBvP7ciEAoUi775mpua5pMqs
7014yiGBt7S92rFEekrB2QgZtNbhYMezcbzrree8ru0oLvui6cZLxyGDnMszYsnI
eflvS14uWFLvX+dCMtgf2eyBRETXka0K9iruU8nEWcQPqTLTHiwXSqXca2xJ+IUv
sOfsDiN7o+xiPIRULlhJApvQ+GElc8pRtvstPmFZxXdbVxOn841k9yE7aWic34Hu
rpJl6dqZ8z/MTwuvfaj2UGF7FvIPeWMSs7eLedb5sxe9upzQtxqJd744v/Us+ZQV
GbJppLM4ttweknWq/4S4szixGuxBaeKw81ia52ttb6YM0gTHj6dFOA2BI0aThTxn
NicG7uBOjVsiZZLnem/q5HEQXYMfn3ZCGS6L1zLOlkvP5hmguWycffs1jHYaQ0FQ
0qWk/Btr5tlvK81QvF75NbZNCOd62FLCEO3xGKLS5CXscwgH5UZS5WqX3M44dy9E
CWcUqaxDTqtgzeuDqPAffre6WSclJOr+AwXnlJ262OV1bUzXmM1sfpJ0o1H+g7ZI
iSBaeNoXvsQJy3WJrwgDgjw0EpEAh9zxBlNZTd1BWAaMNk+QKmTf7v5LdwDGt2jv
kdzlx1i+3ypUHkPN8CQWDngUN7e0dvROkKBCIm4u2ta1kxvh7gkdvzGOPMtynaq4
gUZCZkCeNQwEW49BiqQ+Z3xnONGbUCcntRI035h+Mn9d5Mkt71V1wSCkpRk+ITLW
mOdoqIV/H67B1d6Z93nmGdzpgnrC+LNID07GO8PnynhqVQKpKAJnEsHh6RvooBV6
PsaXX0biNk8A0HJwKCHh4ltRNhX1Z2rkYMdwVOTfTzKFmQjgoCgOaltGJ0CMQWM1
hw0lC/iTf+FGyOjrXVmoRufJ+e010Jy8BWNMyfkrblyP2lHNaRjln9B3PfluA4uc
tOhxXcnibJItPRbtxSdR8pgloCnx+7KZsLJdNvzybPkcLM6vXIcjbGmJajx7lwEq
gJLzJipAuNQ4Gk+l3VTabKz31p2kMaPw2SSaNQK1BfCHB/HvyzrIELmODs/D3YkF
9Rm9mvE0HFiuD2Rl03UY/WYdYpHL0Hc2TwsT43tK01IzboOjfYlgTXT78Wz22eG3
64VWnWynhn4HPMWQzmkqXxSElGHIClHQjxpbV7wDzAWR82sdpt7JPQ0TvVXAz+Qo
YVvM0Rc4EPnwfN4UFt9gCfYMdbrEqcsxXsaOPYkv8rrVyiDbUZUyKm4PYqGpfOTY
0ZKAxI14GyIvd4zlpZFNU7XCMLo7oHnCTiPlOCZ+F0AnEYMzqejdUIXKaZUmD235
GboXBARdBFCT5pacH91STPvIU39nksPYzD4jbyHhj5KVTTy0UtfXDDRb5OuG300T
yBMoZKBB/BAcYCr9O/lyhRtmdSwA8YAmsU9SRJXIKqlDXge8MXmst5K0w58FtEg8
jFCgdKww/Jmpzg+nFVAfrHlx6YsIGXKDOw15XKizFgDAv4bxC7a+Q17fPwyW8szC
KEjAa4P27/G4LLyuCT4YPg6mqSVITfRvEz6okpFNKpvZWU3trKsmnlDo+9yXdYht
wSUcchSpvrezTvp1BnaDaNIXUbxjK2BzdJkH7KwUpQBQbfAmtDFy7s7gKA4oGfAo
tkCxPcP4S/tZcaqAT9CZ1comhGIRQr2aivXWW60tDi2yW6LcTYR0CpvFagtuuT37
tNOkUXh9X1B8PezGhou38KYCKcgyxECxkFDtdSWtiRffj2ocqpNUl0WfpS7T39TI
gSVW+rpUNSz+XkiyDr6Zv7WNIR3VUkOjrqIxpQbqxQ7To0rf7EqqiUxRll6Jv36/
raPmemFFa5eMlTmcUqp0FMeIQn4pSJIuQJVwEXup4YL06NsaRQJklMaA/uVB9X0I
Jnz51zRtehYOKHpxWaHI+H47m8r9eaV6+O4yyVLZY9ZIXmiVb2yYX7N+XfDUZ28S
8VK2vfKloDqOjFQf2oqk7R4xecjl7/FdmV4EdH0h1Q4NQlzwi3MJUOiEEURVBx+K
EaXLEl3RkTHtqRMxybxQMV5+SLba1ljwdQMZRc/sPGPAxNFFrE4Z8LAj1GrZVY9I
ma8MmQCUirn/k0ebhgbijEkrBTt1XfM/yATCARtIjtNL89Kqmx7UGDq6JrsAP0P0
SK7167KMsDXWGkwG6XVHeIGbJSjMW3LTFUb6FsPTtI5RMsn1wpHEK0n0oRbWWnQy
9uOzkN90Fm3pxp16gm/ELL0yon6LQBUDSGZTaaeaZqD/3FWU9oIJaDn6efgDjvlf
3jBX+GCa7TjvLrledBu4H3zJxTed83QSPFYNnH49ytIJmrdIoB1Y8UjiRByrlscF
jaY0oFTFEbRF2U8MW+tL6PrDBOeJf13KEXKZpuAUDVOX4YwNh5qfYhE1gn+Q255h
Ac7bZZx9pCbXjym71CEEgIyTnVd8rgVeMC0mOdt/qNHwtc3qWyAygylu10xmryhy
qb3j7GSDFRtg5vkhAbTYd5yAmzunVVI0A+J+UaVDDFxYP/zx+VYkv6CpswDJKYfa
B9+MC99t3Fz7I7Zx/wvhmMGrjHNp99qyI1k3wze8dZc7uYPwQpjyAK/6Jx4/t6H6
2Qix78gDM+a/uA0yUcoAXMibX++edJHYQNXxekvHQ031FcFtP1j0u2w0eHudbN9G
2lpLHCJv6elsL3lHsuq++uSuAVsMziByvP10wegiBi8eBx1y34n8F7jG1btWqwQb
x8ZdFZuCte2Qx68uos0Cbie+Imb+/mH9JB/RnxhVzQCTnTyIwypNOcLbZUT+Doh1
pVF+GV8wR0HhfZfjCE+VpT2mv5GRubqJe+usHRvo+ivpS8FbxQxew+UeghP/budN
JA7tXHLNZvpzEsnnvaXtdSlYnkDz2AAFrpZdCGWN96SM2IJCchpONNQnRNcjqXOx
IAJ+/ffBD9hvOF8PeJpaYv+1XKJn7Gcowz/k/ngySD6+4NnYt6Yt/m9G58F8rbP5
4/Wpm4m6O+WQu/DgPflIO85EqHmA7a2ZHjJVy1dPF0+jlzvvANtZXz7agQESzb6Z
ibY6VaRHTrmN69YvhMNis2jkzDRb2xyF3ruhG/qrGdkCEu6+Wme6WJ9NYPnyEXqh
TPXitV7mglZRojn383hrfHs8NCz4vHdd/4JkuO2OCLbCbT9I9GXqe90tlynHyyyw
/uYdrARpSefV+Pv7RC8c4cHM5yTIRLWya3Q0D6TJxv/nqu/sJ0JIsHnTe3d5rTQw
1xf2aoPWtEHnQldsVsp/1m20dfnWpujvGGZxar7+PpKlPvTpP+ITDgbpvXCdaKDE
l7piCQHZzoD+Omr1FMEtgPz3ozOCL9jXBP3QMlmeMsCdf5Vujy59Qh+RbZY3VpEu
+5v38qVhZJ71vqbuxxJm1SuhYkahTaMYM1B0Z6YfeEjYZZluvu0Q+mXVftbuvDeY
yOgOx2ezb2b/qfZzhbJbQruecc+2ToledTTT9pyKDMvqs2Qi8cYBraeTc80M3Cy2
aqJoI37ketYMCzwmTaunGAcQKU6R5S3Vy3R05EDU3WC1EKYMNd97cyZhRuVvz6LF
ZE3V6JneHM9+XpSpn5hJQ40k4qyxJNMHngRJTlOpOSeXD3o9rBws6MgIvcEqlmLv
p9XPyfy2rLTpMsiOH5CbPcBRrwd+vC8b0mseDJl4XW6VUemBlXDOVI46WOlR4vd1
6Zg47H1RcbWIX/AYX0e6rRx1dSkkRx2gbxIapqrk+7ffMKopVIxGkSNmhSpN8j1G
AHkWZrkX8spJJyKu3/ZcA7TeKZBxnsH54dCrjq72TybP7YZQr/1BrDa9/rl2jZaP
hLY/aRcb2mBnSDG9qY6dypVAvYrYVD4u2e3r0tt7SLViROGPKhgkfvd9uU74c5qN
h29Ujsk6tiL88tWVMpPANQuoz+aniplERWLhKWqfCZl5y9l89py+D2VVUdjsJTeg
QTGyzCwKHqoYz6bquw3Ske403GPz7osVYeVbz0EGEjAfB8ZiLy7fkBt2LWu+mOcc
cHyjkjIf7t95+U7PYWlUQu5/sxIh8CuHpi0K+d2QWDO/YmBxXap4/xR5zoUOQFCO
WbCJyocXdtvdI72jwWVKuKOKohQx4GuxnYuaX981zU70744GW+rZK3n0A1F6wmO2
9GjDUhKjSGI+UHYa7Lm2CIM3QBvm2VRaQhpyASkiZY2yOjiGWxCND20t9MEIrIvQ
HzyEcxZtLsEB3AiZOdsq/sSUwx31DmnUADPBF2OitERWD6T8o5YYHiC3hupQckX3
nbpArE5AqHvTrC6iZrHkrXxNQ2VJJh3GM+7Gj+2OO+Qpf47yIm5aUnnBz+E0KuUr
rNl8guKVskg3ljld+2gkfS+eGu9Nh8TLYzva17mZ2OT4Khxv5F98ybonwE6bifI+
dZFVJEIQiOl3Z4h5STkxj52XGeo0xJfx8ILVyi/4Bs9z6IS4RquaCGO+Wte06iCA
cX5vCmljni+JZYrLdcS0aMPQxPGj92OHZ9V/ptkHMsNxqrrR4z7vpcuCeNc6e2py
E+3yOlI+Ua8EheOxrLX0ztRtXvFtrs/WO4MO6/IospeY2bYxrNgAyssCqDGk4xpF
P9AJpGYq8Lfnxg1in0/HICtdRjOyE9nuWbhaTOdc1+/EYXdLNkm9F+YecUTU6Gz7
+m+Bj8tDX6VqMZasN2SnJzaAEh6FrlqVeW+F43h+x1KTJNp4ctFbeZeaWRSYOequ
KTjyoddmVb3YRyNVtb8YUfCWOMx/qX6kryDKOrpA/Jxa17PCWoy1U9iRdr8n3OiO
gLfJmzsBl82ywI/kL+LsXRl9/FxS2HOB5KfLIMS3xfPWN+Ye/HjXr71OWgtFLrI3
n5phFe9Lna6b1hJWAVhj5NhvyebWF95OycFs4tlCvzHWTZXJgVxB9A8vGVmEh4d8
i9PSvpagcILhTuBJOvOvN+V+VvVqdJE0svtefaP694KSyjStL6yF2hBT2o4X50UO
3wprfmBPhOH3c3GNwmmPySteWqTPd/wB3CmtqnLyNUABczvenUUqeHenSLU2u9Pj
meCRjhZs7SLCNfmlIji36+mluc6p+v7cFBukDvRd19OpjTy4yUXLBWc+zu64NRvV
VINNEWtIjqwlWrlh+6NpSEHL+vh6GzYLPYUnYlWH7blojg4vGnlVDz+DVrsGxO8A
QT56CptT9gWvffeW2OvZfnvtRoQv727JTnpWxkQYet+yhuWCClIA49jmp8IcUQ8A
VP+yXiUZHUixekmNTsedAf8Y+QESRy980uhdO+vgH7ZzHM+gI/dOyuwl/Gkb1OBc
2aCuCQVnfzsYc9j2Tpy059x+lHtgWY6f95xgS4+r2aV2ZKYsdcfblXgXC8T++TZq
7NXDcLj6NiDapMpUh58M0f2aDVANee0Murki8f/la4HROu//qjnZZnyd+WCdJm4I
8eOEU2y5juUNFPrRGkyeSSk6Yo0T3Xp/Cq71fdTRTQVO8U3fXlKi/0a4QIkGi2H5
2cImY5eOZ9XgVHPppaG/EKeUtvRO8lYFoF0hCuYkhjJRroJxMhiAPNx2D8zVqVdl
iy7zenNr78kdLX6fFYJFqS5F6w9R1I67QLYpY6b6GWjiUsQQ+s7D0VtF/FKrvfZ5
p04kUVzQoZdXXq+i5832RgBN33Co8pf6g79iRbseEr1KAxbcl91RobQoDkqwn45i
RjuXZG2hxH/haUa7Jjx7b5BzibH/ONn8G7X+Y2YWFt/dNkYmJ+06W4Hpz3wtUCDd
JOnkHZeIicHvxnKpmsqX49p5uWniUuomLbhfBa0i8ZjSfqB/tGDW53bcAsmV3pJ6
ErILD5G/w1Df7ebpDXVDb0XYGi4Do5pRHBCtVyeZksm6j1siTC6ojfVJxA+PRkir
/Aoi+dGzoBzckkWnk7yL/rHSpJ/yZDKygcVFmh1371v72IgaavH/qzwgYMJg8TN8
7XM864jEWlB6agm6d+IIbvzzYCZPCfZt9Db4osawWffXH2jVAi5PdeqhJRbasltn
GQxQjNFUsYX6FLpqWS2tDjpz+FuSTfsvnj2Md7WdwzcjCVXgkikrzJ2QPNmyKJVt
QdCGYF54TnZIebR/Hf/tCplo+iefU8W8+mVRyGQJTXBaKSWpL5wwtkosy6uVL7EE
4zLWElZWQlyp8mb2uy5Sm+8vsZ/Z7fT+O4qqVrbojdGPD4XQL+hS0A6+e1cnVi+L
BLBpweiwdMqE4xA3yci04CNdBRb+hFu8Lj08Z8kEjkmVGy2x+uPyz7H2LvxM43c4
L+dn9cITO2ZX3kRV6u4o2sjusOPRssMWM6A/v0KQIZDNaC8IqGtd11nQq77sRymu
ir+seLu+Sz8PCg4s/QEkGGvmnoAdNF3fVG0OROptcfZ+mTeEFFP/AaDmj8FG5ihM
q+dvTMk5zN47kEs9b2wwHRp8kAYjA1LBn2PMInF4er3g7Ysoe9Ksp//cnjvxjGtI
hgVaFQuuQKuFfwn7fgJYD83Pej+yAEUVjbIC0DjiW7aliSClcDCtqHOM6t2pYnrn
19YvSJUQz0rTP2vjzQx+6i0vty6KMbKupQZdUxd+NUw5AceF8hM8D6sUKAndj61T
LNhwod33Or11TgmPbWT964gakCaLq6L108F+HT5F7DNHkO7dNof0Y+smtoWjlIzY
jPNiyhZNkRYxc+Q151g+ws1vwtD1/BiyrALXJqzkQ4CeaMwJbaClkBomB4uqxuyZ
6MXvBF4hhIxPs8HcaHGen1Zj/S3kzIf5WbdZK0a0DoNCB6Mk++kGrC8dE7IZxD+f
In6p8fVP/Ce6P8zGk1Ezj+rP1K3THk8ekAeU+SaSpoPmYIibnyBaDVoDhlZltB/q
IZHNA8qHLaDXD9chS7ofkYwUberNQUSGpIrPqtNirXWz2OPJ19AxHra7gxLHos07
zRinucgSPutCtP2TPdZBaeHk8RJTZ9C1TvUzvNr/p8m+P+CgLnExsgsSzW4RbOLs
65TJNxU2pPk/RvKI1qhJvOo01cmu82q7qOQ2SCaBxYgm/ScFkWRW9L9mt2YAYulc
Uayp+SrLpj7nOO50NeXkZsCZiwD9y7G3DtY3th+FM4UjX8p9iMv9OPu+9vOdTSS/
EnxY2N8osVaDnAQUDbmuoRbSv+3FFXt04s3EZeZyAigFMYjfwZl0RsfEhrAbuIRd
j4gE//VgRJ/hMMQvtRGsLfwlJSHV2AMZ5YR4TdaRNafXjUjZrVyWj5vm111MewFS
+ae0BBEsCoUff+ZvkhpFb6fT5j3FNa+Q+Xma5ulcsRtLMAa0bOUQUMEqnSk6iNxa
QitUvnxmLVsYm0aL+mCe4kFP6/hCq3b/QEegrajOz9bVnB+EgizNKG2vMiiFLh4j
Xn/xuecIfC7Hg1jSe7TRjl3qPKTZ60Q/dXbpj0uFNf4HXluJW8ZuhK5MfzFY2H1D
n/Ba0SVy+QmfkqiN/pv1/+D4D63SziqRnUAG633Ay7ng/qSJunHeE+zSumTmCwzu
g22dKyVH1/Yh5wVnjpWtjKc2DdmtYeEcOeXCt9hbsBjtwAAs5wbHF9vx3SoOQmMu
LtmhsVMCOtVE1KRAdeIYQLK5LPmZ6HoG118Xu/Yopis2KjZ2T7rIgw2mUssX8ZnK
joRy5GNwoMejN7yVGiDQDHr8SyV72gx+qLv65mX+5KeXgNBM5EbzZJ0iKmJaCXuy
NsebhQ/OwQS5Axpv3HTZhZPkzb6CrNJdeIab8XtLKf6jFENWgAAbL6rtioQI02PP
got5oamthR6lPWRxOZH2xvf5/Ywqk7foGUeCl7n7TY1lKRp6wzxZRkEvWosCijXu
iDuaa29IDmUT0IWP3w59e8NnTpDQrzb75epQ1+hbcMIJEpxeXag5iIyaSF2FBupD
3G7Ne9oYsDz+pyNJoV4a0ULl7htAM9VqerrgxxLZkEAI9HQp8cbCW2Qnugvhj4gC
bQZ2MXE/m4wUrnJno/++rWooQbATV9N7ZVk/ipjWRjCMHQtpwlBuIG5Yq8Fv/+YZ
UJKdmjULoNGhylR/DVyKYlkeaeacJQIBwV+B9/d6dY8OxLAmbuH+zoxXcHsLxWdo
ivjgckTiVjDNUwIHHknOgA/21ER3zEKYJXjysRTxfAkMN9rzSzuT0ZssbxVHIcZE
TlZGgVQlvhEY9hiTqvwrD2Sd7RyKh7FItBuFuPrLrfFZFBVSxULZ+IiFPu0gg3Kt
AJ43O6nDOEzY0dk/u7Et7TWCECoO+DGi6KPNd2UrM8pjbjzKUiRfxLh/TfOdYhKf
3MFuTnHWbtg9Fqw56sfMQRlMsZzkjSykNm3wrz0ymx9ET6TZv8QGHCQtSDHLOiI3
dJxRo56qmwM0fCAaRONiIBI4yMju6HR4FMgorE3Cj3Y2bBwMyyPaUSa+1sdAc6LL
s+ZR5ehjNZ4Iu7A7EAouh5cKgUyg4nYbyN5gXFTDEUBjwsqDZdsrmezJQdxjKVY1
jYBZZGIxnF7O7X/SJnsDn/W/pKE53HN56xiiVuqm4rWKqTY+YhD9n+xNYufe0z3J
1/cv75KBSIukzHYBmIEQRYC905Wqg/jD6zsbvCcdDuYJnbTES7aEbUE7JTZ6H6Od
uLom7di+6dcnQUZHZptRo/IqQFqKaFGbMRZC2uLIori9l2afzbhIO+k7wKPVwO9I
FrhXJrYPZ/v6AjMHNZp1mI8CbmUXrP8FefFr74r4wwoCQqQZCDWlYQWiloC1Wa66
8R7pmVQrVH1leNz79/DIySEx4mYLQtb9PEmWmmV5lhvQlgiTK8ZcG7sM8kjL1Yf6
lByTIyoz5ILe1sJXzxFvi97BWKLKGagoMhSpClbJDF3thYhVNh6GhE2wUTzgOwBl
JClAGhzZXN9vYBrskxUzdbIrn8YXjQjo/ybg4E1iLKCfe1HQ2RPoVugzKTZTLNld
bYMFZjp4rkrF0IFhnxMXnTqJD3JKKHvnk1vZVaKnW4GBwI20gCBJPHPZSIk6ziHE
EcdshjWTkB4EXGkckL51ikrDwC7YbNIm6ttfT7L2YaJ4DLANqkpGReCFzL2LCAHc
i8RT0v10TaTPeZfrU96MP8ktvlN0GPuuo76NqiVvkBq9FlTU5zpn0LKd2UqcWYre
k6YldJRKsU6kUfte6SJvQXLn9tXudiKGACl5eV0zAIy1uXGX7ddkZurcCPqWuFQ1
l10gIVKCLUiMNJ7KuBU2h0ha9AMSw3Gy/MeV9jN862hhvTuR3KLZQA+hGwMdBC1l
A4ocp0jMJqKl2i9VilVgH184SNuvl56x3+M6X1CU2EMpNYQLbzGzBXWsRmelypPN
X3rhgcW4a7cgRU7Q8FyW3PDUhlOeIH6TJeBrsS1tSzSc3OWECGM8mjYk8ZN6+DGc
x3s0Sz+2xRVj1qI++20FlUwvTbdJnbkP7F7YKFkKk0mlaUmHmYw8o5F+pM7DT+yS
bcxdcdaQ+F3NjKpaVwSad8ZIt/a/ZpchcQOhOyPa+6zauyUMgkKTeI5l94bHwI26
eQwiFVqGY0XHqWiVipRbgYrTiV97VEnSpB9YOSRR7Bk6FjW8WDoJ4F/5V3rTzIDD
vsuSipFcpelovN5nYgBwV06rt5eeTtAg4vzpSfxJ+zl5hudxuPxgoJmqTFqHeW0l
HepCUI5FjbGLai6DqUsYGv4bReuH0Nvdw2WnBBHsHobIz9RiPpjU6svaMEtziPDK
qISd8J2lX8WqcYBcVsVJeJ786wD+wHb3QZhgkOv1ULdwmbeV0lwyM1FT6KvBWlvy
jSDmO2Cwse7JMjIHsnqSuyQWxQcNjXigMgvFwLA2LXLvjdPNWMy28MVuIUUaYgU7
gAemG5pE3fol57xmebEF+8LB/X/N70N77UtYSJmDqhbv+8pAE/GHemskZ2i+WT/t
lKJsyj2sugxuPPUePqrwaBG8Z67lnLD/YA8ChIrD3XUXeeiwgSpvnHYebe6A5wj3
DdyPQxWC5oeOjcTspycUy43NWlXvQ1+802LOwV6UxYP/n6lRPKn2aoFPk7FZGvL3
PbVRZ7xwVY2B8OUGSLKqRns08EfZf/R4RSEqVLOAXjcf/uHRjZ+x4bDwNn2S43Yb
NwocpGhWPxotIdKnoCJlSM0hwvnFzGyuQBHfF/c/mO9bqt3Ybx+1HeqHHkXsFEjr
I1IcskUc6wA8oPff6MSm+GVOX//0bdcf5SEmJyawaEcfqVBZ5dniPpd349vqitys
/tSvcUW7XkP/fmtr6/bCluGPQEbPizTN4qbYrimv82Uk0wp2LxTRHcrw5Qjhr/xH
a8wpiFHRHvEjQOUeFkj0p6CeRlr3vxL3JjolfzJUHkCBIhRgmQHex0NsQ++b6ap8
NwP9PCzPVCytlxg5qUYgtCglcBBOurJu1tvea+2Kg3hiTv5WQ4GQb78x3iHpVJ0x
zhVkcGYZzG/whbMAG4QzWJjMX8Ayt38NkxXHysnXdyLt5iPjIU+6UyRpcKjBeX5j
wb9Eeo1YJUwg1/AlJTL4POIq3eR//3S5gCzzZJijnnQ/3sBed4wJieelT7vx7/x4
kH7rQWbR0c0Ga8OKcgSIE2bW/NaHiAw8j5DUMvNS7FhFCRAqrLajMm+9/QFAKt1w
jefNdVw5VAAI5mD3dvlLY9ib1VtfsR+0ttNLGr1fGRP0u7C6VPkP4CENijlzlMDw
cQiOnsEOO89p+xPAQFvX/TULuyDcdzvHpanzqaWtsqatp9eC/d5NVkGwYHRR18/q
0EBXx8/hAAhtLr8FcEDnChNuGj6dg2ibWR6fQcUnEGIi1U6ZknfXi1vjzkCrJfm0
Kx0YoO/9a4HtWEPANGQfcOsSZqWlZKZkbHmsn6TwZPbYmgvNmkYCXlbKOqSQFjwt
dOVJnVNbr03np49lNfkfzjKGpZ/ZTueoFJ9Wm6u9h6jSdDg91yH9AzJ1OmY/qyvZ
eZHjevyNZaCo0O6cuLQNgpI5z/ADV/QZg6MvrDvvVzpP8e9v6XgVPqtZ+0ou9wdf
guZZHficawdGvAxgzgOBg6rvUskJrbv20H2VMaSr2g9MsqyCvWayWKmsmk/wH65P
4IR7XAXW+RwojGBCvnes1DEl/SFGT0iXjYFbM5NzIijlil9R3bgPYku0XkLm/i12
LGw63ePCIOwgVWkUXfhaos17GWKkLix76B5ajKmDdMZGn/c0EVv0pSkyrFNLmHMs
ECNNIBbXbqAC7q9DNZun66ZQsgi9pMkvC8XNSmA22TeL3oJvVlo4IKgFhIcCJ2jy
WfzgiKGejP7FDALKNO1/Xska227KE8uDeMCLHq87OHDFA5JKCgRtOSNovklUH/op
6OKoKnLNBitSs32ts2RUbsRRJtKeUB40c0xjWppVP/dzcgrZASigHiXn55W3mdAV
TzII6nOJoWWG6CFLb2/DMBfgmpTHwt7ZFcLvIn26yeVAEuN2T6pRfSqS027ImTnN
htvZsJnFS8LFKEkgmzJQotTDMw9evXhNZWm73Dd/vXjB0rkpETMd1Pd+aOKgYBk/
srPpPSmcUZomrJNC8qxln2fTJoKc9vfvk5aJoEdxRcr9jRGR61u/otywLhzP9Z8S
on7ArKQIlAjWmMNsptpMU2H2727/V7DjS63tGKWim4olSHoDMpvZrrspP93sw5o0
kLFjtKRvPUhCY5RqgX0KdccMsHWnkI/PhPUTxdHNjA2sf70yATpSsu+QdJkCuo0s
liI0/k4gnBjuURHs6qK+/ouCscW7s0beYsq/N9V15ew1ZOpowu1+drbmzXMxumJ+
I3j0Cis0x2Tubdn0fBfQMXW9/aC9CHQmMAsm684YUg/e5/opzPnbalxrl50Ie+A3
lLsbD8zpH3aLJMIO1sYDfgzfaKlbSd9pLqxE+4s32eAeLSLHm4T/4159R3xDyI2N
TMJ/Hp8JOf45i3oDBAdI0r8ERquU2oecGvTnivZt57p/NHUo7ct210oIVhT62TMN
ALD2HKmNXgGZe1+Mshct275FTbbYdfmZ23kvbsH0yjyEXFvH5okvbbt/w754MCiv
oH+yNFZk93bMjVQOW/vGwY91Hbf1xIz+tg9rLArrRrNGmL4PkXTB2DqyLgNj1TBm
9Xtb2b3/46fcetjqq71nZed6QvlbYz3sgUccPBePLyydW3gqBBTaMR7nt8Aj3OXV
4gP04lKUKZq4V2xbfKXVtYJGu4R0sLHu1izV2U5PD1Yp/jGsvLBIbmnu3xEdz7K5
ypanZilOgIpSz0Tdo//74+rEKBOl6pFKJ74VskkAk0pbchZsU+CGFWxyA5e0UNhx
bkxtecu0pIU8r0htW8QHSm3y/lUt7icJTzpSt0mtPEMHMuRcSQ5C8/bjBJlXe4lP
oGlitmYwbbG8tVMJBsWfKAjhwNE6gmWd7vqmYRDLqdqDFvpT2wyaGXC9iUIb0Syo
Rm1YKgux1Q+bkCZAYyiUPeNsIOYIwG+gPWHwyqk60Tck+dOoDrNfPoAW/S3Uwtku
gBfH5Gv4cYs4ut3rNFnu1yolfotxFt11DxtTBYxBulGUE2cCfsVMXS5qyw94itgy
xCB2/LUOW9CFfarS7SoFboN1wtykeAZvxFaUkUQRQAZlIHsWbmGRGhUiXdt6OwjT
AohLB3RMQI0zn6OZwv3iUWJNJ5O95bEqor/R/T3B3ob8lfb7jr2TeQlZQCSCyUhi
IldSEFlLVhT+usTr1Fpb3g9juCOmS8P7SyllGBFXoq24aYJDKH8gTNL0y3dN0zer
nZvsB4VUbXIquCUSwHdLLl4+SsgIzS3W08PrLAQvR44pThnFTS5k9wStWNzwO+wX
qtORzUb4638Owh1He06Nch6z2fw9mmfi7w4czBMGwp2VRLA2B5EfaAYL8PCjnGIE
Crolbzpja9loUrGaWtv84/RbQAEIU8ghNTGowwxeZSoMIg8FHuar30c9io1J+Yhs
im2uG54hOSRxS1ZnLr21cq9wCY/2rnFjkL+DV1n5EzupCCPA+1rSXW1H+9p5rJyY
vt8TZE+Ma30oO/Q1vTe/X8yspX5zsoxBWiwS4yJa9FlRdOzJpTzPWi8ikdT83bfa
XtH+JgFnUtPs7cGzeZcHvs0nEDLPgGXlNNm9LYpZ3WWFCTlj8z7gOXoJmihV3HBj
VsAxcNonC/3Wk9RbJ3RW0j+vdOyAvPcj3AAj7U8/SnbjoQ4DsKzW+qvSMHcqipoh
DuBc/QGy9RgDYKWu27ylFEWS1nJNU3up0OYUjaQhGj7L+wtUQc/hXhofcS0KuW7X
7lEI1nBue0Ubp4Jif+Az8VzlIU1HW2xnvCP44DuzZ1CHRaEcqYHyjNwOSFqFZfax
y59yUP2MXPlDIUDJdEP031cV4pQ99Wg/38D5Tmj47IhpC21O5Y47JLe0f78Gdwcv
eHTUfgiU+DFqNUPXiL3+xbWXFU/aspqWgVZLTySRYIreQQEbq16eAGZPObkZQDMJ
GnwYn5c/O9ItleeRPCuM8Ji2i5E87ajFxGj3rTkd39mW5A6lJks5kgGhNZpG/SJv
NDOMkOPrn5PVsOPGmp1EyWpkeTVn4FE5YiiGnZ936ujyqS4h1vKINeZKRudLTREt
3a4K2Vbrm4WfJh09eYIThMtYO108eTiOQyuXQaNT1PDh0NWxzgjS1aNKDsU6J/4N
tOg5jFLTiz8ZyXa65AuxV/V2NuUHmx71yZmSbuVI2HO9kJvabP54ifpV7F1X+t5N
ieB8p10+uQoBUt8I051QPi1cYol43J7P0cZ5FSIHRsWZjZo7trT+7Um9TE5rV9w1
e54THKFYbzc+ECPj25HrmyDw6keDzhEdUJsIwHuW+6SAtvzt/AH+43yE0bpVDGfr
Pdu4m/vlYqpupeQdYsZjUDYARTEoUQ/RKbK7npMnI6Ebk7BM13rUxMoBevPtvdAC
0jMZWHrwj50LTZbFk3lR58HVszvDqXhnqMHYa94qpxSV7pbMFkmrU9/cOx6abXMM
w9Xm3QQxuHwRxbZug/lrRRO3Te4i9IJXwVEZhp5oA4V0VwwEoVqS1gF8ITg6zLyk
RDKyo74kPBR9uV0Tt5wDwqoxOlbabbphupi4l+5WHn02h7CYMcqmsxcS3D5PRN+k
vqZGD/rkzF2yfR+b7vDYnL/8tb6redrARl95/XYHJ7ngC2BsnXOCjaJFz7Nk0bWf
bWPzH1nnog+ekCUMhGPsuL3Hx4jAiIu+y8Pxw0pS6/ZVHXSh8r3IhgC6jHlXhL/y
7WiHpv5J0fq7XjUs08KEFyCfooik/39i6l61SqtXoYFOwb4ne4nGi3RNEYvDWs4s
bU06i8ttYNKCcIGBStTJyV6ZmAPKywyDhc42a94aU2tRhA+2gO1ZdjwZqI1PnpOA
nO6PsemA0vV4dlX84pUrzMysCuOGebIccSR5DGPKKXhit8kXehpU6hMUdvIFA6Cg
Kq5C4HcsrwNf+01Q0B6ULxAAMNG8bc+O65nE+Fu68N3jbx+sSYyWCAmrfUa9A3wS
yJsf0QDmCPpb0MLlWBPTHqpQ93sqE8l+QCmr/IyP4aSS5F8VkI8RYNohk9ZP91jt
ZHElYA3NPQf+Cb/SbVR7feoyRtEDduWUH+pjdKFWq8ZEbIEYdpYPc1MVbOyoQiWM
N+o31vg/IS9YGoAIsFf/BHCvXPF9LH3uyJt8uUFixsmjiziRIs4tAJ4cXddlQGnc
6Hnlyyd20yAv1LQK8dnhKLdE73u3EwSoY88XjD9eFIMnGARgUIrzjuFfVwgEad/b
/RvEIoPvb/hXSS2nnG8euvOA35zL1VF66aTQwQMAv/WM433SlWDOSSQxHq5FKSqr
bZNs1536YqJ1TeqsceJZsFYGNX9lRTwNG8+q5CrjZjlakMladzHdPwOEHjeUQDXP
XMuA590RABMFbW6P3KITH4/iEUsyDFVowAlU6zizH5OujE+0RdxiD5zFuQPlSTi8
8quKoQCXtxbObEb9x2o91V12PAGGzdYmATcaJE0b1GrMjMYjjD9LeKIBU9WEWpYW
3DK0cCtW5cYZRGiZbtEVIDGIRev5lnMpFxgE9fC5QQw+WN1Kz6uZZCXjqVc++Zds
jrH9oGUQpAsLT7uB0533KgaCwmm6S5jCgoh+SDv/GA2PKRMXrjz1KWJ3VT4Txo1t
jK4DrWqV6Vh1DorSfJjfB/PbJWcZT6pgo5QEWdlVoUhGIAF2cNICM57VNMam20R2
PJ2BT3LRL2qMM+SrI2nhoqo7KTP0U1jBz2ouP4k3FeYOPUwsHxdLnOfPI3nqPpS9
Zvj0FQzxKAQXtwFLiEaJ1FK2q8qORyzCyoo3enweQGrrRYFtXHN8jDsAKki91KXm
iEeXyelM+NAb5fHadREGy0C2IIA6t8Fv7FCQHZOeBT7W7S5b5P9vNsRTnoFuK1o1
T9M3LGXzyxUeHGtts7XXmAMXRh0zu9NwPbZTwfitIUR7/tR5dY9YSYqpGJBmDyL6
bPqWajzKnsMGJ1HQKa2s1K/qy/oH5+QjTg0vLbyjIPivbqEpQMNW4XsoHY1p1cAy
Xm4fJCNyzSSFs+ja0ggfuctMQVC2PYvLcG1kePOAEbWY7jDk2SwF77ZoaMqV/t4N
bry7lUj0vJ1K3+l+Sz4SwZ0037I0vFJYvQ/rnJ7VApfQyP7v8Qeged7GxuRqRe1j
mY0muDu8TSK8q2QLue4j13/EwAYqa5Vv2DGxmJuQ2pCzg7b9qwImrGSV7foGPiRG
sBcE1xtb3gu4XQ4xT3dlS6PtyIKUdLWrUYwD0yGd5fSBKctZhTDOc8w0PN+FdUSa
KufguNqYBzPdmvPqt5bbnjFbDB7wZSeovuri4UuJn+eOQsFdb2HGAzSPeHkjGGLH
MIOTRxWeZzQVnFiBB4XliUvkEphaAYktky6AM9riVU7aAngbTYShaxDza7ktAiyA
jbkov5f9xxAbT2AOzibSd0Ns1NE8tdVgaE8c5vWSOQKUwG9U9RXWGh7ogjYUFkFG
PFzhViGDngPWQWwJHlcf2mHzI1K3/MxOmxM35efHxP51mMmkiPWc821DseQafvtd
wsXjvWjlqarPuPStfHEHsRfNMm2FB13yah/sA45wWGp2rC9wcctUXW7OPoVYH7LS
xcwKdyewLlB9exFo6v3DuY2WmrjhKO8PmutMajBuavybSEj0TmQj4twogVzJexBe
SYDVmXkQFUQwxk1w/BBXA7Cz1hi1YzelMS8kldveUGvXPKOSJFzKmRwrk0e0+5jk
VClX+Q9ApGnkFJLNyBCQGPrfrUstf8Tn+d5CpejUqFRKyt61ZlbSKUGdMnZMCr/Q
ybhaeRWGLbZF1/pV3is5U0b3znedFyqfIxxsCOe9tLJXDKzHMKuKsHLbATCl+5UJ
4QUxAfiQe3AUMOxILK9mWAIRmjoCnSkYXiS6BYydY+XgpI32qdybI5PGzMnRZJou
Uf5bX8XyLoXTrYKcyweAxqwCoNrI8U/OD5WAtL3MQQ6Gs3gIgMTho3YebeJvOD3a
fAvYweJzXJT+1uwAG342w7eivBMYR/EK0JiUSLlC8zNjdR/ObveNT9Tg6Hs4xCc8
kKAolhsu69YQdwnZHhprJBJ3mbCRrEwm2YgZEZHdjXhhnPtnOq4yNRISjIff2HFm
dfktEtCrGGICIK4HHs8X6OZskeqr/AxIHoKmLKIVMrCFDXJa/OM8xGQCLKDZ6IQ+
u/ARyp0PJvSX2OIJf8ow5dRiGK6O6+TlrYrpV5YMe53vKh8MrWtcE85mpvCwHrCQ
gCTrnHtZyQB9najStuirs43Vvuok3fNoHFxh/ZIgSF4tQzNe4T3kuGH0nkuI1i8d
BcaHWZEUArqtFgV+79z7YGb37kMOOEj1oRbfKpIwX49KDXoF94Wmcu98EfHabuIC
C7ouFrXAXkej4f6vCjkzpl8jouYPhyx0ViRKNRXoJ1oNVTrfMMfWsy7PqmHcaqt7
SUyGGGZbzcEv/30z7A3HokpgEyNLBL3jikLRVPWH4OghudHt3FPnWQtoREQdEIX8
4NtRgvtuF4GHWlQeKy76bQ+3IclWHeNa2C3wu/GFyCOsDn1Og8khW9pUD7/rQ0pa
j2dMO24zju/S4z7DucfKi7JWwf+8Tu1J5xH3gaMKbMs1V+pHEtrb/IbKZmPNXqsg
cDt+ChQPudJsA2S+YbRYCiALlLuLUh+7zZ7s+EpQslhv7b8KE/PfclLWlPhokOx8
jgHSFo9JRW1kzw2uXgEwdrEN8J7DxvVgaYVRjwF1JxFgqr6xBQGZV43nB/N5KUSj
6lbuCEYyEVsYz2nCVlMDcIYl2cACzyGycLdRKiPdnPnc0pY3lQU1muBOVzB2LGF1
Sjg706xlgERuNU/3YJm7BS8dhfbTiaWA1yFuGVsZttfQBvEmB4z9+gjz4zQguNZA
dgvfTkOhN2wJTjk+Xo6q5NN9jEeNKZ0wc3V0GsUV7xHHVY9Sy0CO30lUgA7cFB0q
uKOzdCQ2ZCoAzxILCWPVXKQyeB7S78WKCx23HheF3cKjZvSN4/Pav77G/q0epud9
StYLalxGMYVjmoVVd64GtY8O+MQCzOkuiWB8hcMJpn2uzdZmn3fiHXQ8Pumso0dp
XQh2TWAlKBO/01zW6hZXz1ZR1bOosFR8pS9hP82mZli6Q7GF7eisN6hqKtI6jEqT
MMA8WtAhuCqIlVLDkOLw+zeZ4K908katflQGCkXepvJYbZHIYUrZ1OgEvFNSY2Mv
PdIrNvHngryUgtF/2WrqewvL1CXfXcslJnDaaJzppsagJ8F8/SZb4MdsY3fbGQzY
B2fBdXSAH+CcWl5tzv7Jj2SVVcbY1xM8wGLAJlKE9RRiC1YCl/P1X4QLpKpZEK7y
CdwoSXpW2F0N6DRj28atJ4x6JuSh3ilheBEn54eTSBrPBE3MA687apLFy3MQfLUx
UpjGfATF4/tQLAn4Yidyt3IT59Gpl4xFDjnCQmRdaaXlXCE3rSTTtvehdo5nqAIE
aw0pdveCWm0vKJSIyWQK0a9f6r6qy+XcZlRe3z/WED6M41PvKegXInpcEk68oRe4
18prEBl5VN88fcyKRkdsddr+ZBKlpfAYMFXvl+CF5aHjiHS/Gcyzsi6Qykho41OO
OB2U+E1ec3BJGXjLMbWV+v1BBj5U+Cl+jcXF58omlz0Wr4ZZj/BwoIk/tdoEzSga
LNc9mfYEPyiFD9otpgmWahtwnCa5RupUamiNOYyAM7tbQD/ZCBCMtg/1lC1ayfLB
tUG4e15urTnjSoEA4oCT3vIXBQl6ZnQUZ4DF9Cg7dExzh7Ul+aMCN06JDkL3GNkS
lgeJBf/KxcFFOHmTkHh+d6VA3RtpGuCeYHV0ZiKdLc9pDR1Qj8agJtY5CuoEgIOA
5pbu2QHQx0xAxFER07TJmozXnbxFBvLP814ESavX6jDgab1jwk5ipi3Dp5vvFohF
zxhaBoIT2Q2l4uF5yZTQjCO80zAEs26UGd2AjfmTe0pXH81b2zYOuJ3rt8Jz7Npb
H3JVAqtUihqmwQCeykSnvunCdEIbcTvty55cCtzGQJR2m3+g20/YFpWAi9lUjIwA
FkA5ZkcbxjRH6swtEaSWIka/yUKnCjqcZyCIGU6/P/n1/VxOCTIe3Z4wRuSAb1BP
sWEya6kNyb/z6OYBO/ZU25gg+mbIhtgTKX0EzgXTNIeq2u0Ufl0Tk8nPF9zkKHua
LnVcKQ7DGu4+VdIdu7C8zcCEWYYq/ZQTqvadbZRCJArST7ySrp0EpZCJJYg07hb7
40iYvYSE3v339yFEN3jyd66/22xMxxoedkEbL0LGYLxaOAw+HaXq2IadloNu3X3W
G1KOovyfUvPF/03wXOB/3rdSWJtAKfodzh6IU+uQXDo4Yc/CdsAmp6zVaEN0La42
uweySmP1Sm8kpCdDyaDL4m+uICx0FHmHsiqP2n5UXl9mvLJQmTTuHINdkEuZXasE
Nvb4bMBnGOXv9dCYTgXAskK73Dt9tqoKK/tEhtGdxlD48yqpcTaMGHRrHvZktTZY
QpouMUPFbpSipRYK8n93ttbam+349lnZMq5OvMl6I435dQ67a5FtO6yCcUzFi3IZ
zsXhGTGnowJdpIq8U01MLxPlQQS2gc+La2KOuhlXXp4Sf4ZJD93foHlxTy15eLoQ
8Tw7dgBKb6EGlNuKzsMAAJ9lBf/MI7UhHL141QozIhNP3jR0DKb/Aiv3DEerbfeA
Ex/srLBEFsEEApUi6elpdmMvk5r888RyO5Ji6NacxBEAjCxW2ZWQjDVz5EoZDWBo
DmmV6mSo6WTHWSP0U13zr1hor/hJUD1dyJd/sAPeDYiMtwhpCFPxAjBQQ2soBF4I
q50UaQOUTqd1iuhlqDeBhDYzefhF1pj4uNRmT4XrFhJ+/A9gIhKm7+/OpGgDe3Cs
OEGYciMQsVrPpSvzs0j6aJpxXXAPNiP2+baUxYGLXlJB6bnfFbU4GA7fGZk1E+jw
6cv9EEEpsY1qDklkbggEgmsKt4xZOjNVk/uo2f4LWxpY5n/LQQ5dipy0NjS6jUwF
wAKA+4WxIxGFtzNkFaVib5fWYb93JCp2bxwHTxTj3bUq+qnTQL5rlh5VMp1giEiJ
l9jfX6wbkh0Kj1YsIJOKJM0n7z5d002rJJ43c1b92f6HO2SMQ87oFAHqOoI4wqV3
wyEKfDUJHt9gCdPBRQuNbfb43M3BagbkhbqG1vfd6d9umVAw6WPGNvPwGE86Oa6g
h3nEizDxzm31k0EHScTUnvrQGZdxnS3cvBlRPYKOktH0E06suoyJSb8upanTBZbl
E6GdN/VYBYU2gadCHF5/dQtXRY1ExxUuHG8yy9tqN5n3lFZsXDkblwtzsWTAtZpd
h+akOBH1DRBlAkM+/ErOQ8ifwt91UyJG91bl+h8yfIz3vKkYE24JdVH/+PJvqwBT
YXy901WnFuWYy7/jDcMgGiRXB2Fd3h0fa6rAr55lwIBwLE6q5j7NqVG5uFDjMHtK
1CGmsxAKsxc0vHoGU6XP25/RkezJu/w1HualvK7Im6t+vpP5FLsGv4Dp9ulYlqet
esHdf5GfDeek+xKK0SC8XDPQx/MHUA/nV1TkmrKT19HxbsRVMpUzp6EmcAPdMEf3
hERWb+ZHDMnQBtJ0itv6/Q+QbCj2Xc9S/zTrK/lfs3412ow6E9xNlLJ9YVQzuC17
nWyoHwdhUX074Dp3ZGfc0lMni1S/3T2wMBjXFhL4HoEpSMWzMI/UFzAZUB8MK+i3
q2rMYxqJiXzu+KutnMqtnqEaqCRHjEeX3ZcTwKephuCSFNi61bQWCcveInQ/grIg
+qnzX1lvAQeJqve8Jfz9yZ9sX9Jc3MeAVxMcNynTpLCXgaSBBSiLcqmLigPXFLF6
nCQsD4K0xDy+VMmytaTE6tuoDuWERFP3QuHGYRiFrNGk6Ae+PSVeSm8HOWVEFJIY
WsjCx6V/BmUBMjRaSFw56bYCGjCIb8ekt3nFEdT5PDtHTObg01U9XybMfBiWCWPy
3i4JKdBba6m45xfPTuzKbZ6q5RUuUEKlYUGiDvBFKZzhMyR2R46LVwIs0UswZ2rr
3yUPX8YzE3iJXeW8f6jltZvNMGn0408EZ3w1ugLL1Q1K/2zQ6sPnqASu2EHRdqHW
KjwhDLddfZqVKjbteeN3uhUBxoSmaKIpT9RMzq/v8C4VVy3B3OxSnEIMNi9abxMM
/EOnP+l2CXLTo2Y90y4wypjB2RTwek+76Z54VumDsPcn4s4ip6uilXSk31zwZpez
uuZiVSfkjBKaJpwaT7cTjgJUgrOWVEMgnlwrpVIHwKakkVr0YceOSQ7ZTA0CctgV
8VvEBOQ4ueacykTyK2+u/HrnCdmwTUOdsG1Opf+QP+cifeCJKzSnlFCc4A8ZA6As
TI0/rz/xMAbugET/HR8PKafPlYzTRq1bC3LHX4Kyzz/WoQD+C+fJRlJiSiQ8Pr+4
zH6bWqWwaq1KMZ6WBfK0f1rh5QfhhmnXKmBxXg7f1uzwPH29x7RsLZ/H/1lTTfor
8gwaD6jDM7ZpnEa+fHcLu0FNqlBTRyn9vFnjMNS4zszjd2oFu3bgB10kKzSjCO3x
NizMuyYtcq5zrhfBZFBnGZ5eaUQwcSZE3yKcaBiOinfaVlJbtiIXIA0jHc0X/ZLc
WU+r7hJyOB6J0FJvLF4gPSnkdZvvzvn968A7lpbHtYaWu8YCQmKHAb0OD5SbSYJf
HSk7n7Lxj9AtPRySLrGXlqexEo83DvYsajN6uQd96HslFzdGc+LIJC3jMrlEkL5C
GDAU1TIdT74PIIzbbUGPrtXXRAB8OguigYpjMsN6Q5C4OwNLE358AbZCcwce1Lok
mdgzvnwE4NJP6sN+dicbBeNgp0Vd9RD7HSCs3s86schgAiEOnpTNFwLccB40sgUv
ZWm8L+JFLd+O8b83gsjj0N7PKgqpbNkGYO4TEq7TPZGnPO4ZeyVI+8AQtLRp0QvI
pGJnrhWtbebnvGa8BiUrxC6A9iFAHmwk/BIQKNph5bv7VaUuF95YYD4v6tvFM3LX
11NNW4kHdcgojVCDciyhOvy79Fa0fV80AyEousHoeJRTQoku9dsoj5M92K9u6LUV
9PTD25heF6vzN2GMz39xs6hKy9FCAJxphI6+HdWm+rMlTYeRFgBiAnGDg0hx79m+
cgBhX2WwJfIpoJxxpE0DfskMMfIS2v3kmHvszs9cEXEBOteZQjGfFrOzmqMpPRUj
I9V573MM3D/coMlgKqVmvlQJ+XlcsgtlDGhsza9XB3lg4gVV2KFPI9cjEPxJ2G4x
jnNGEMXPNhonhgACzKjk5j1Gt2htK9zzc5rEOg5CcE3c07X7GZYwxspHmRnAGtDu
tyyxk6vIB/+e+GM+wjMqXZXYvjFCBYxJW29teQJyocB5KUC5pwK3po0NC+IsNvE6
nOx6qX8zaBhOMnPEauFaQRhnrGCLVnaWv7TM1+ET1sS5QHOvjjrzP/mq0n2Uo1jW
gu00BrZhcTFjrNa1bTLlVMSL6RUuUy2RQq47tKdUxh3ZwwgnQvbzUFV/8MX36E9A
fmuJYWRHzGVjt8NXudZD5JkB/RVBlaKH76PpcRXcba9JNis+czwccIzr+t5i/+oq
LXmdslzFoH0YCT8asAGsex1klAvUx5MvP+mBLQacUGhQQtvlx/x5N7bx7j/e0Gw+
XxAzUYipFSqbVSpPr+nbAnzSrk91NL7foHqPF9ybJ9uEWlkNUMqjmM+3IaUr4hUn
LaQhgCh1GrT5dcuk3k9UudTFFsrXEO1RoBgRc1lN1btX/97kS9k1DQfmVXn+W0ue
za/93mHEoQ6I3rBss5kQ5yEi79LyL+S/ckD7IjCEY0wrDgqzA0pVnXqdCwJsWBmp
fLMcPC/fsTG6ccEmMBMJ4toZyLfsE+Jdj1aPl5/5mv2jH6PGbkYgtqC2mUN28F+P
gUxWJa3j+CGaIbKGblAjqPPeZlPxk5ZxcKqp/rGfd9vRNmwtx+pgZDG0lKQIGQUG
Q/eYw5HFAorH9wydzmNyB96AIYyzgUlhAofeGqzCf/gqKdybmrgMPBbZbOYD1Pw9
VshN3HMLo2J/PN8Tq7gshypi2BfyiUUUZlhUXQOiSutE3YZWt7I8QbfbKNRJNCeG
69wfHQiCKxH1z2SnKK0XRia38eal+cnGtDQxg7evNB8Vx0dfzZX5XJYoaLmEobDC
4D60nKYjoIUYRnMRahvfpQvTDTpexuQHVoyvlRyRI0EOojce7lNLoKGm9x2thgpe
kZpf++/qTMXq5uDlZ+AVAg+9X8IHBguL3ORu5tediVSkfynU1fTA0HMGKtHr7y7f
f/uzBHXc4NpllAJbwFHViGuZwuSc8ajz8eQqob8b1MZnfOaShm7Aejgln0auC6wd
ihQy2NnvMCshGypUI6SmWwRHcXX3YgjQdjd3azeY5PRvXbA+3XIVNIVI1XHx+GtA
mIh2Z03muEdXb9qDrTvpONJ3EjbITO4BqXjSeiViURQS9KonOelPDZPunkaLWxUF
2DLZ9yBzFSxFhbSKY/tk1fl1g7SC9rCYXOASErS+cpVEo7w1DGbot4PhS2wjZjl6
cV/KILBz7OSQcFH4o4EeV9LQUjRPxMk5Cml0UP2vX6FuevetX7+LeKwXorQfLWLs
mJTepy3synQo3cxtjZa4mZEE9ljUASUVzIH5subU76ADyxBNfw6/rprdKe5T2BYk
4/OuoriwjOrgNpdVoesTPmRbRRtP0LDcOnZpLXjvnS5EAJ1ezH9U9OQf1/frAFrO
PLeZ4mh+xzJ7gws8VmPXRdFRn6lA+0ma0csx5a2MsUbELS1FRxDahe/f8DRXbVBH
ZmbA+p8ecsN3PDFIPgLd2ClAOBfIGKk+J4pDymPcDrJ8LNiKoHt9gt79ibzBweR5
RCYF5NkUMQscUGsxuI//Kkq56sdKQdf7JcVoDd8eKUzqLuEQdczgBQdCQJES3WPo
a8/Mfy8cOg+zkxXNwn8CPSprdnbP7nJSh3K9AD3R8IJe19wCrZKu0yEVc8joAZqc
xNGooGPxuENIH5dkTNXqOpRm6U2zvyM0mMsB50UBcMC/Isg0pRnUaB9XPP5paaI8
gKqeIvBugQUHMhrtX+60npSbfD4Kem5Hy3Ma+Uuz2G/Bb6o3ujrZQx3a+3R7vvQs
9Kwp6uB03COssj6WZTWR5/WGfAQiz62dPtIDfQ6pNLMiUiKWSxdxynl5BJc5p5WU
NKeHfJA9tscWgwWiiwCFxaei4fy2hQKTfqq6mXoVa6Jm1rNfQAUwgCejHFtY4HOO
7EJI9AGY1dXk/UGcXrCkyS11Gc42WGSE3kpAuA5x86OJtlk1+OvugqUO8u/oplIZ
owZYcYzNFXmY8zT4nxpGlUFPJYMSzIMbP7Nt0nVZbasjtjokOanZQl0ARQ4p3g0J
ifRt5fowIRTunHmjinxJzPVx06K5Jyo6HJnJmLuKQENVfGrlya3Yvs/dPxUaaeP1
KJI3+vfNRyaz2Yjk+oVAMTIfyoUxtMvTa/1G0RFrTijkHXM9VYmnYP9vy1SuFOEA
aPG+H5aeGwn9Seh8XruU09aE4jp3LRUEdaVLi8F6w2wX0Q6gwqZUhs75n+989sO5
gyvN3d/+yuJltxR6kXJf3Rs9Mku379kW1PufG9hpBSeNTm98tQN82yBZHCN3qg7Z
jU1dCWb6vchoSFV13wAvGJPNN9hZwddsWqEWhzt4s5lqWZfI8vV8BPlK0vmet1oI
72O5gn3Sgkdb//IZB7ff0JA82pbyVOowckp9HiBpPg86IzBf9o8+Pc/x+6oJfp3a
yxmT9t0qOnCfcHTpEg5fsUp1IHmGZ2cml2vX1qIRFpqemtB9Ip4bSbwb/HMVgsXp
4+JZExkz8sX/dA3f2JeLlEGd516xf8uBQ7pHW5fT2oTferSotogWMmRZPOxNH12Y
V3shYmljZh/oXurvaSSFU/rMvIRoqWxdvtJ+C7VOHVa/4d4SUeSGzZ+WTj73z7jD
n1OeXArfaH+iXvAm//RREEk89PEmO5ZQwdybvnXaQmF0U/+48omlxF46/41swWE0
yl3VJ4mOKfSkpBHSb7O3fUigWOBec6Z4s4wVf3LxZLJ0WfdLrnjoYz2bwtFKfxSN
ukfDBfWv/uJ4FntrpSVwgaosZfuCuQQA4gh0ZIk/IQr85GdhQIMhWzdXyMZ4Yybi
YxqXcGklGFkUDZyeMbmoU+DXq21RGzWvrJRk7OMUwZ7HvNhzOKD9XveFClyg6rd5
wW+7Jx/D/4bz17IyQ86grShvIDT97+djouKpkwyoY46RL9dDX3qDGVIDk6HBmV7I
kFPdljlUOt2TbPanIUYFETOGTVy7W//r7u56xc/QQC4lHEILUyQJLYZ3uxKUVC4L
L8rMxtb6djsi6Neij3ZyvLGz/Inz5DyKA3yj6aHLsmd6sO67hr54msNf4kj4DL54
bt01bSDEwBZQOigx9VKo132sA6sz8ZEYqn+/FXDaVWMS2nAEGOdVFGRogZT7U7LG
eqv2AAaz6Awn6yj0sMu0+/ssa9H+ckOZyqKSnKPCcYCgdoWaZW2xOJiFgimhQ05T
oitqUn0ve4SGN4C8QYoM50sxZ/QeGs0mOTYf/wzZxS9fC6qNcs05W9Q+dDAaP8nb
BTmvSYuqwzQe61ldmxGoxVPnLYJitVedCM2kA9BCw+PM4/B2FUKCfp1cgCvALjAZ
V1iw02Wajov0mb7uCa+Ky5eqlm0qlGUfrkLXva0JM875DguaZKwJyiLDUWp1G6vU
P1DT2vQNyQMGnstupOMyr0KScsf5t+6SmqlO+sEk6SC2hBH2jhn83ZWjdWCYnwNv
KAb1Z6kczp1bjRM9gUk9m7O4qqtYNv6fO5bGYeRz9z7TqFfdgL45SBd4UXS8VkBf
8J7touUv+wn8lzserNbbJnaT46e6kdkGnb6vZdp3+MpP2vtcUMq33YyQOiHPELYE
p6Vfdu9RkU7k7Bw2u20CtpVPhKrGCFCYI6u6nsq2G3wLOS/i3+E3S9yylx4wMk+r
LPifzgP6Zp0FZ8S1JKJVaI2ISOMPKDF7on3qRFKpWidvIoZJ8hzSQmcH6fJrODah
wVl4YGRiap94UMpntu0YS+ePRAEmLugOzycq5vuWCeW2GoUK2KGtdfBVQQnlfEhx
dE8LAbAuunnp7t8XqL4lPjqQ7ntMe4W93ZyBbbpvBIOJu6epPDLY6dnntf4OOZyo
FUSy5sNyqdTj0HB5nACVf9hNSlOZnhRgyTFH/MLmpy4JULIaQhXHu2kvVdIZWAEi
P5hEMl9WnuOYP6Ggi7egQ4KoHgPd50gQnp7pWLtb17KQ9z1nxjpxuAsDLHg0LhFG
FzPht407UaDgqaATBRipBaajAtNm8pHlX1jVoe8VcnA7F9iQbZwFw2by8xHu9Gpb
EQi0gUoxH19GC0+NGD8EBpZigwufw32AaSxMYfV8/VQQqiTznvn2dHK4V7toOt1K
qh51AO7+RHWO5AGLFvcXEAL+dXJMw3pJibDyxDU99+7x5gDShixv0j/kUkF6ZQ++
rWK/chBCIfine63JESq6dCtsZRHRLJ4l+wsuJ4ifzFV6mfFM10y0/9V39tuRcT++
oatSGyCU1GVxcdOZuzIBgW7OCGXrGQey7loQwFrHiE0H1ClKH00a2IPvjFJaeWZ6
NkHdXMjhRtEZ4IkZ6aEm5V3sKkM53O1QIkS8Rlihd5OvdtBBvO+qTC5wRD3fQFuB
3mQLWAPmRKlNqrPQlBDbrgOOuIS9BnBC8osPy3lEcFqKMJJrRG21OC2GO+yzEUMm
YzxpDadZeXzbBczLRwvKvIjbpPHgLTkjGZiN3E3Htsjjqnx4T/ijgBXmKsZ0Ftoa
plnTbO8UyEegsdMpEEHSNPHVOHejVNuzi4xSVEOKY4ui5DdjajcL0NdI/tvq/j3S
nKWh/chwUPtL0UXyxLu52LLgNJU1lKtAKcHTrMGMmnqdrBY/9cONpgmiOeCjdmyI
eJV4+rlaZoDfGgaLy8sndqSiqQ/jvgQbIMFgdM4UL7zz4WJL9jXZY4vreJZlAFWD
F1xpSEJSiKymOgZ+dVhfxFjCTmQ4L80uRZ54Lb0/a8AgG2i8rtJQdium5cRwAD74
7OBggiQ/OI1MdzQPDhKOWGcYLJW5cMDgOG1wUM7HoyajdlFq33KGQymTVLWLPeV2
/dG0FUnxjeI80uGrZeLUbSZ4DLrfEGkPPOblhXnhFpW1Jv3NfhGgAChD+II6Srmd
iXwWzsvpi6YPKJR9KgLX9NUCOJmRaUlrI/nYJKgO6HaVCvXwnUttAD2mWna89cKJ
wbwlPxqyTFUTdb1XciB5l+98R+EjKbcsbn8KWL1gXEz4B0NdzcuNxef+K0ChUKIY
fuo1QDWi3aqWiQX+pnzTaiK/CWC92FYSFVQQBYB6AuDx2qEzzth5XW4xO33aScMw
WW1CEYpBkFOIPuDVUDv4jDg2DHra+/HIa1w7VqwaO4LnBrawqG/uQ0/Yvr1IXDB7
mXQd4X2SRpom0CLeZ7QXwoe7VUcWv07NiUICRTHJO8blPZuo4C0q0RKT9Av2P6aJ
HH67tJ5JA2FvGeBtCFoF4mpgLgoUXA5At7O0OxtrRA2uyHxxU8QZ4wsdnDKXx/O2
+4NwlXSa2uEF+yIn4YHTsERB8ZTXdStUYF8mFITHmHE3oXTk+gGNtkvaQEmLK8O5
N0yqbANvUoFQ9hnoodGvDcZphsmjaitlaTIP6jfS4J86iA1ksVu8zM5jF9pUg7lj
0hEjChTT9xK4xKENOCOfnZWbgI5tk4gv1oJd2r5eLplMgMeEV0A3tUARwUTDSGqW
rxXWr19cTUGaAbz+UqpzPycrjhqsbaocY54kcKQbEOunRJcVQnMJv1v6E7H8C1Wt
NrfCNYwVQ8iWh13MxN5VHmermNMqSkbgvGqhpJMTOinF7aM0BTxpfukW0gi6jYxZ
YUhLsQ3GjhkExlAN4QBTRzM4KNcUXsIjfZdTSKMtouWRHzkMtrLQ5vFw1Kcndqvq
WRq5Shdq5jhGE/C7DA1UFZu0GLwkSbJZSUBrRKbA0ODin/fTTVjMHHZVdzNOcGnw
KpHQ7GU7fOzWJgi0XTefFWzx99fx3z84qHYpg7HD6iFDfsZmQYwo4yZqgMpU7qyL
eBXudULvfmRxoUe3qu3N++LHpBnTRKoaPYIPEh3+RhFz/hcbLVtrSN7SN02WmMjm
Mbd4suPIDIBnZyWDq7jiQmeKCSQvmO9cxL+atw5BRwbq2J6GwZvbsSwu+VBKLocX
jBXVixw/hR0hS3qUeyxqj+XjWjyPwwbIGuDTWdlqcTfzr7tfDVNgMKgNC9Sk8JdB
00G5sZNmrsY6C3k/lk/sip+FW/slxCNL7x0jYzELJILskTL4d7EkTMmg0EnE1Beu
7niG4LPH2sYHIaje6IaFCeEjK0Wo38Y9/v6Bs0rBpQBdr27Jb1zKha42SnijDDRt
E6kISDrU1/vCdSlfAkXS5f6Fh41WTBRzJnoVVaOsTnCj4pBfuNQEyNGrLbsXOIOM
QXopvCWVKT1apustFg/x+nsWJp7zQ/KqnoD2ylvBYqzDMBv97klzwOlNqD+r19Cs
kPJ7wI9egpDBEn2wLwUVS5K6ZSTPrJET97JgLAohyecX+LAI4KDKFAyov/5luWER
DN+/aCWJ5MWxH/fYjTTytqPYNwProwpGtmf71sCGn5ZLfUnc5OkknTpm8UyI2yV6
0uhuvvm3rwFzWbSMQ+QKCSYqkavVPvBfx6dTZCUV1e9pOe8ewhrA+cusPBcTFEHV
Lb1AxRNiAefpWA73lJUlQjL8/nxMJMGd3UfXXk2+EUVKqR8/cZoNVpMUY9tImSgY
QGszWIBk21MuzQ9/8y/nu8XuZiouoJukDTBMMC8tKh8ns6HvZzQDxdGbLJU3u4YF
az2fXAcELcGBu5N3H/LJTObdTMMAWZyv01Rh5ED5LMjK8DOgsiV5tSE1Rb2+zn/r
fYWm7K0fP9/btmQRm7yfCxXCvseU0M9A0N1dz4aTlDN6g3fHzrRBPxfQx3hVKhKN
VBxxLmDP/Fpur+lrvaWI2ERoUK63rlGOBx+Buk0uZw8RhI3HFgI/5w5U2lTO2PvE
xQ2SjbNzGCxQDVk3rjT5EtNN8VZ03Sxijqdo0al1l0d9ogl0DxmnPn8PQxmSdTPb
Gz2hac93bOWUYDvHUhSVVEtpMMbS9fJavAJeGTxmiOblALGVY9kQI3DokiQASWJJ
EQlRU2DWsRPEZAvVOPZGLEM/1G7O0fsF3PwayHl2sBGFuDKCAmsa2Ib9ro2j8uV7
Eqk0axyf2U1ZXQPCLPLQRaN5oS1obceSVgqwyN5q0PLeEP2QIvZin61gtq+UsF3o
7KMLdWe4DyyMsBiY7BVvA5oAYsAiQJXoCeIgKYbLU6bbRA5srjXOshvP3okhr5cC
NWF15qafizqnbKaS+FauMEUhy91Xu9jKpulq+Wcs+imEhsy7fXYF0oM/3GzZgrCh
VZFNL8eCtnxgNtyq3PiOIotjWEQ5Y8nEm17dkjreDAnulN9T49g17kJDQAzbZYzt
6oyCizRhPok6bXFt+SCXhbCRUXZdKD3yust8k0IE5CbRDEQ3S+ufaY33C6XL8tVz
2u5I8sR/hGk5G1m7CeCaQBXmTdQ3rz9XImsQBP4OajK8SJbCFt6YF//LR5kMwMIp
I5KnBgu+xDK2vurhenYHiRuWIoznGBc5HFERkhCOTHneOLGcSV0ZqhUhDNJa5J34
ArdyqWZbSBusfMGc4xk6+CP+yRCyuZpJCwC4r1lKv1SEl+Cqb8qfD3JTFqkmIshl
5+oOkL6E7q0GUpaA0Xzvdalu+esuzWjLt5HVhMYRzf3B9mHrGhXwz5Evdarld/3n
S5I3Wht9QgLLFuFPt4xhpSbkge/mjU8K7rPS3CISVAkKUzb290Vy4WMJkH8H6gTe
FkGwBNhxWiluExZlBJ7n5xz1F0M56wNnJMtRWOIN/fyb1wV+5rZxgzIYEyB9h6qp
YCnaUHVrovFUxPbUwAmcwq50bwYXwpvwdflWO2rGZyH2FeNp49ouHJ+OWfB1Ejv+
RBqp7oKcFcASEbVMP7ogR6sSfDVeduNNZongM+K4VhVyghX8RSemELSBiLj+Uryn
B4cvWepG0rzAILOHpxKAO22FKzNkY+V3KykaB3V9mfUR8VHAcZFJ3YAqLsxSuuw4
ZUmxVEJaBTC9akkkSiMW0szt/VeRQgLVl2dZNqvWYzL32Y1aRPo+db7jb9PSgInK
y1tDEI8vYq8gI70+bFcP64jN6x5wgxkz7jHENdV489VL38b54rn3/P4w5KCvZzZm
3aOSf713bVRbM2YoSE0JX1cTsM13eFhxpiM7xsfzNlDA3eIIeHwtfGscJuZLFG9k
dShahUVYI9ullbbbYA1CWTbOTxEt6dL5fkibkIxaSnJStZhBvT43nCptDgbng11w
TGWPZPFeZsbcghU2AR0iJtCXgGFuYnnnL7JrnvOw3uYIt3A/Ezu8/P+9SiNVV8/v
LceLQexfoYEBs7yQKceBiGhkKv4vt45el42EH+uRNDQegfAkj/yTnec73Id7gOWG
C8m365yPs/okDtdv38JlAM6XWNtUb2GxscaYE09ijReyMj5+2zUGgazyanpv98rd
BxT8SnxFKG7qDaumPI6wSs976LU8pYJEqZMEVdleHZVcWz2SzOli4M1UL9QEYF18
s/vVXTXKc1wiiff9eG18T66z5Ng4NLaCdm4kdrM8oR7wsvUE2xXp40ZxTGwvdlWL
KrpLLQnoplNdabXQ9zrx4cRyKbRkqJ9nSkiBgBaoBFmopuqJHzlnOenmMgtBILF8
J9UzU/5GixEiOHm02ADmERM5jb5mHKEcoWuUvMYqoAFkPzAN43fJCQF+070LXFRz
SEoQYAM6GmVstVgKBn6X+MiYTz4ioVs8aQWgSrSZig0m6wXQsDQ4YmLDziuYf8Fi
eADdH0TUjqMr5F8jNquw/X11nt/8/yrWYjETRhZtF3ROtJyZqCb/V9yXb7w3Iws2
1Mzw0daCOeaIPuprHxkekrb3Z0CsTaBHITkwF3BOTYBcv0FVOxoZv66GhHttGiwq
lOfuMI6j6B9nr7oy1FSCSJ5z7Y2lqixWSquZPZE6gq65+qRDbCFY0E3x4h/CjKDV
dg6v2GPfJ/rtPGJ8yPMnsJrZXcqktuJJoaaieLHznVueHe22rNE1wshOH6jMioVq
j/ostBq4Js2GbcGzOJqZ3v0tCdBAPdQw7jXLODggOGi9U1aJPaSHRvwn+265D7GQ
hrofPe8XOXMLdAQr3d69ZGrX1LwkyZ+1C0bUPI1rrXUT2fXvGOWegWeRTTMOPn4W
Ccnyt0cSNSnAxhgOzvxA4OSfojN6iXTf/agGkp0LA8P1kUGCkJO8ghttaX/igw+b
CWSH3uEjU8ZXoPQIzKYmzcFyMw3V4IKteNSIeQB63XWld4+NccQDMa/IFwZDP+Nr
JdRFjjoCwly1PCNUfgkLHvgU5Vkf9tHbDy90uzK3HBxBYjWooiu7d32hLafigyU6
tZrtDdUSu8ZWOHkU625GdlTAO6y+6F/NMdSnTMIAh6yFExVPUwnyuH8Dglqj8lPM
9wwGfq1fR+DH904Wdv1M7mYCmwNU1qc6xyFmkpCamM3w13j9REDJhlVxG2D/eEk7
Z/G7roEKupvmprxA79Ndb9gLz+2DoZbYa1gqMpSbuwEHEZ9sr7wXjJloXffRaacL
xKMnSCt3IvIkWeXqYK7u8Go+cs6WKnHevLfSXH3k0sKrTd8koa5PaSyuO25c/yhJ
dsFN4e0sCEgQPTvVoWN4kSR3Vlajf/r/EsC/1PABSsLKV4X7s6joh1XQ6FHkpPSB
WEqiT7rfge3DSET65OgF1R/nxRidvJFN9sv53AUE5+pLqWhIeBljdOyZBdlOKgf3
jsPyv7qhkzeC2K9AHukMvW88DZiha1T19alFlDg8xXLl+n1kNL654JQKDaWF+ZG+
iMjgzzSCGVsHcqhJEqiIfNGltr2bwuXt5ctxTRu1X4t07RTxcEs5SEbql3frcjnj
KHTTmg5s2nmoleOdQXbRphfY3lunvHdtMIdEZUhPJg2Kr8XHyJku5Lm4jzVn+L5t
4nVeR1y3DHl8z81skGRV3xVDCRb8+4sCDRGgA1ui9n0mZeFUF5o0rqT/tNAbLY6D
UPtORGdMnOZd2+ACPahTow+mcbPyn+OHxJemYq0/0DJD6TjfxpYKFFCfqwHBEbKU
f4ITwpYsluH1e/JK/8DBLOnBr65lZCD8P4rX2UvZofafiqe8LGD6Ht/wWm5nTDhO
Sa5iuNvMkFfMXO2o9spH3vcf411dJBpK3RR4mb6/h/mXsII6juH4Y+Ist2NOo4Ps
WNPOosk1JpzYhZKks6sBIluY+91zsD9l7hRDSBvqNZzQbzY9M4tpbCbSMU8157Vx
brCqQyD0+y54ceUTQsUtgH4Ax4JHM/LdUSFzu2QSQd8R/O9jQtps6AHo7w3lWjwA
5UwlG7gPxGxq7L8GEkmLRaHsBh5Nx5xaid7RS2uRZqEkeW0H4woLB9oWCCAxks40
lxthSeMPYz3oFWhzXTNMpwVb2qnZKM7ke/+LNSnPEKTdut7dKz+nt+POSfNUHcKa
05wSyGedrW72Isu32qJYB4wG+srlBJ5EETup/HaJU7f9CFt7fhXm0vw5gbrFV9oK
4SSKO52X2ciSGTghFpOf+7dJ9/13+m1TvAFUQR94C2XoOfM/4o+E/8kfwx6PrB6I
RuW5rNwJKDz43oDcXu0FmDcjL2jSwnifFLu8PXnOAl03w8GACqo4gPTp0zh29l3k
Q04jDiqxCzpXmtBSzT4WGrV41bbfaeh8t8M8ibz7ymS97H1Sj+ubrjp3x9iTTA4D
UzOYqQc+TxPeljHSZZ81BrMAVazT902vN+kORglaXt+xaDZVayUMBbq4FKXFUWOi
z7nyJ8jmvyUDpKBW2nNSUFn5Y4si/yLFlQO+5r0kvIrpqS00fq1Di8/20XFqsU4j
b4G+slzqLn5rQjHyCRTvtw5mPHiPi9nMFzNjml6UjotZLHa7+y4yV3HCPQkEd9Is
aOrPg5S+ENmwmIPxPS1PMNrVxn+HSHs/+Ag4VKgJoKcGw+ZxQ9zYA/iVDpiWdAwK
bYujYwT0HyhxgHPd6xnEyH8evovoxY9MEw4SGAjj6Z8/jjt80sMKzW4+8cDbNW+2
96xd5fIsNNaqiJ+lPVE2vIeGEaK76UeTGoRAb7efcqCja4vqqYUoDsVPqOP69a/K
Qrl4rdKZkoIW/emeY3LiPZy3LkqudKxIt1yFwisZN7y1UOk7wEUFkdNSi12STLWt
n+VOSomcHYCB9L/lt/uQCpf5JD0IIBOyUuZfgnG6fAg0Tqy0818/QqUo9Eixn5tU
Ean7jdC1O17MlbrfC470VhZqfQroP2rv9vsUGGgeInt8I7sLoV5U4CrIMw8Hyy+6
jhoHgG3yuAMJvgQwR6kQQnW3PdtODw+JYLESVxjp8Ka06lV1l0Ay17DL96mPQs/s
NgKvLLsbGcooxV/3XLIZynk9GeI72kpJuB1LHCC/yrVeRhR3yyHmZigNWwMtinwV
UbO5K/1nMH+sJEEOtUU9ug2rxa269hZpoNMzu+fV9m4bqbUDe/FQXUJusZgp9zxp
hzzJlzNFDH4LANPoGKchCslCsknX7U7J8msXYnHIng1JCrtTgeahs/jcPKhYkTkl
RiQ3qZk6jU8UAjUrgsd534KZy0Af3jlKw3g37M05onew2CSoRAeFT3HxZVF+GreC
zjDAKXiFWNX93NN3MU2OaddYpMnjlRxyVb82zqSU7PR2xp7/BRFFLQV4ZchX+GGW
UzY4lY8tBYX2A7dnR3Vcn7VfJi4A6z3sCk/13gxRsr6zHXTbryth16afXRyS3hYr
C4br47qjWtPBHN0P4toan5ziqLup4JYvi0ql5tofwNp1aKdKqUtlOovYbDK+AFmO
mxXTxE/Dtqsd5s3LRctU+zJ75gL9ELESwLKNXrkDYHJRWuNJPRysomUwIM724JUC
szYkCHMC4NLBXwuBUfqjNJ6osWhaziWyFVoj0QeOWCW137gWc7ZnGekotqApjg64
cjGc+zwZZO0v0SVcIFSniBNjKpHoO/7azfUud492eQ6KPNfEiTDfs6xP2fvDF9zP
LTVc2U3zBPXcHWWcpFs2oEBXOpLvtLcYmcTaKvqtuNWZ+glf8kAIlMIi+HP8dqbd
c59qAzUSUEKvjOQVvxdZxnfJOa8XutU8vEkCARSr/8r90dOj2jAARXqiZ87SZEKi
UdBcdaeTK6/DZ0qQDnvaq+q/uh8taCTCmRAjCxf2Om/4kAYSXXpIJjzWRVeVwgM9
JhFm+DCYBZUI0KT/36bXFItQ24z1tVT+Xt8q2rDv8JEU44kUHRv7P/NoOEoEzDV9
bfqqLs1fwSQlp7hSCOQZJgrwuHO6x5QQ0bBN5GAy2hvWN9OoC4f1ULoQjCjt9R/P
0lvg6pwE8RV6hx3Q4c2il/FiZLmoHGY+lMwX0m8OThL4H6Euvf4eviPN99C1eNNI
D2beOi/ABCRJPRwe9PktyMvI5BVV/cznMeZXP6E2HNwA1hiM4pmqr7PJouAJ/Wod
EzeJPsKjqeC5LBnyjN+LwrLMke2+M82gHvS5R1aKqGzxJMVkKHN6p5TOF3s2SaYD
5zbRSX3Y5lKMQ6mGbFKMZdBS9S2N+ruHQvViaXBVP+RzbkR8FzOlT5ThLWlPpxMC
N7qHoyxUT7ZzjvYvNLd/dPMq1BOIDCgrbw1Br1bRZ37WhWFkIorKFO2MBQ3tK4Gt
Kau48pkBM2Cd8YK37lW0RRyc5Io9lWT30YScKCgRlnZQ1jUogDv3IKJlGAZ6yYHK
f65VmiE3vONEXABFs/4E96cB7IEV9gn3JPeVW6clC//ghS65LaBuyY5DdJpZtlrN
sftqoPcgF2lw+YlkGBMHXu8mk1Xjfv1E+zR1BrwyQ4lXbSg65oAlITQLqev6CC15
AwuW129haVTHBDJ5QLeHgWNcwjq4jcRHjR/Q8WdqSFg/xAQ9Ye5P3drqFj1EbEqA
V49fjIQv+xtGRtHmjKXUu4T6MKbloWsYFVUBvHWZo+E4T401omzAptRjPgFmIsD9
VWgbQzio4p7yqfSDRkI2fFZ5Ox8DO184CFG6TOJzhi9WZIpLsqvqZyrtBwNR8cpL
cqymF+f4VAwSDbgfThdfHRoWBg/wli8+AtxSphKy+FRbI2BY4WXs7xkcT26pxYpZ
tBKVzIUMaoyIsNCiI8ZY/bp61B48Mq90+MdspOMnqrKgXffLPFEIiP4Ok41Splw8
OOMWmsT6OnVYSId1MwJxTDQqPLXwBNDcEyPYYTGj7qVbeyf0wMvaaDI7fIGWKy4M
TOlh+qT2Q3cMYscfgHgXoshzALdBVLmxaBWaWnnQXFONVlAxKbjFxo8d7VT17/fq
zbLzan0/hHYb19WbRwhcGF8NlVeTxr20Ezgj12RKnXxou6cz0OlH0++B4ZBKl5cy
1adhD/seHQIXMZboU2vIg9bCVoGhbPppMsy34zbfq3nx/4/1HiZNETYuresbZzbv
ltmRlKhpokpJ6hmvcvWtUnnxPYUoEa4ra/8AuXPCbr1Bj+Lb5Ar/H/LOilVxyBbn
3QSP0na9D08CapT92pYBOCBQ5yG+fAaigWBvCYw7Nu/6CPjH5WGGvS6TNTgjFy3i
QdP08HHmA2X/7AXWMdxrV0MffOOZ1HdY8jPOdnPWyGCb04zdM1wruCppXY79Cb88
zyDmGOlvRfSxTMK2Mun+93t9L4VQkiinZJPXJG32pfewbyLvEhCj5rmp1XeKWkui
RugfvF4a4QFD0RuHJ0TuvKSLGW0yNXAsWPL4Xzj6unLS+JAchiqH5M6pmfTzY2XH
VWIS264KunvsFZzs8RQvFs+lTuAeUYcHnsj+v4zBhchb5pmHlELJPH/N/f3BHktr
1BHZl2q4CsB1iLz5GoCtDbOkq+ig+yrLMceq49OiTD9sK9Ui+CjFL0Wtuvk3iAY+
2pnpfQWDJRisT57rOqhA/5OO2fUJ3tBqUu0qr5jnRmtmnfsB2tr3wu50J9S9QIsB
rccYAGkO3fQdwSlMVkuTIgXB50iHkAtQIUWN2Oct35HBcPQFTDBWkpj0XXc5eAtn
GbJsHLA9Z1w77jIq69uHdTW+pDcE1Wihd0VnOHFMkRi3Mab5k6etKc1VpkhuD0Rp
J6DBxdqQqr4e6CvCWFHqduKZyGED6v29ejNdCeHkqHxLe0G+eSWkG4n1mhCal09c
w03OADZhGePjZjBxCKNil2wULfnmDVSL4ZLFiSQFKNdhHrZazJlzuJGDNOZJkJMM
y0J5D/neovZom52snQT5qUi+UYEn8H1emIHLDDh6cNfRbifVmvMYos1thM3k4Qhg
56cKmdmdupnLK7nSYdTDBZBjZHsYeZHcjyJsdPejSuqp7lDb8JHlUR7F5PXgaqCt
taKX57svx/UAF3FfnYJulEGOS7irPWbf+Bnx3wSZWqSfSHrgMLwBorCIUuRueUt8
5BykYp9w/QlCrHlG5NF2ZDxGXhGgvDwU1T/oIiafNz8DEz3jHCsS9DkAZgtwP63r
JUb2Gqq/gPbrLx/cfiIY4cwx1q/GXkVWLphWjhx4Ek7vKqFK7RnmG0ZwfDi33KW0
Zhe5g0/60HkEia4M7YbmBRDu2hBvYjvaFVO/WVWLiyII+L/yHEhG8AswypxbA5sI
5qSOwMbSComlTIz8TLo/XCUUhev6h0QLvQyQXIrvr7tc3eaBlHDb92QQpnN158FT
5RxDttVhiqx4HRzWyc4+enJ+t6wQic84j6BgWOlZg42WuQoTHDQXTEWgfCmAqjiR
9Ph8RbqHJNNGFbhYAEEOAv6rKuAG/25v8gHMHLoVhuOYZK/q17O2AiV6kBcCOR5R
UwxKZSbwoEY+blCi28BR10g6E9C8+kFNjSjG3Mds8vjwKNG6y0YE55TAg3AC3ZEZ
sI2sftmNFjSCq0L6Ss9nGRYmiBCKG5XWlk+6rR/6tmHLAQzHL1UgAarwB53uG8rt
sZT8EaRqVXa6aswopbq+2M4/svaucI3Rr22XBE6+Gth7A7VgegLKFT+CvGtWHLHU
qZiw85d4Xg9C3xhAMGEgxcML+H1tzuc6COVrSZ059V0oEhN3WtRFhGg3Xe21lOSl
kN2C+BXXR8hBcSvkJFsU5soY7Db1Mx6GQ55jQL40AvsFTyfGMg85+//pdVy54h9f
RByaZLsgPL8oyzqwlg3+8eatgEB/i74m9y8NXZfaIGQb6VL4GTwP2VkDxEr7Ubft
ppvkbZ82tpsvNaVGOJlDKouDrnPmcpun1W+EeaqYXEKJriXNNZPZHm7khFXqL+QN
eFRcnRltlQx9HWIRJDeHFB4e7vNI+0PLKvI2t4Awj5ZokWioUpHpE7BAXtDwc9Hs
I4f4nxTzHrmoRzkOdAQNIHOU1daxiT8DskgJBWGrdmgcZJtt72Wvp/v/w2J0SaPS
gQ4QsRfFUP9Vxn0s8dUceRerPyxVcagdFRHdPD2FWObU5KnQu01vXSro2B07Sg9l
n9LSOVGCk2jepJazILrPvoh/KDDNpkRUAmqOkaUsdLle9+l1qox5rD7jSVi09SBi
BZqJvv6Mt6G3HpeKarmPikQxv4kixjo21EUYLB0UPPxTCgz7wO0Ra3OQMh6xWH4/
OJbY/dywxVz3OxO/eONbl4sA+HoALCkioXAorwJ5Nz0hR7S/i7LIKMn+roHZTe57
CWYpAZJ8RoH1p8WceJRWtNLBg5XiubWd1Qn9G0Qz0yCgZKLl6ABbtfZUiVch9SHu
tzieYINXyZMgvTODVMekd+kPTY4DOr0wmTZR/IwmJNEf3t8AvalI2KX5zFS4RNIt
NiJhsDcWQkN+95d9ORa0GPcyn8thVx2dUjFemj0JoZqRWpIrQpUb3s4pP7CfOFPj
XD/ox/265s4nD1uZKXcBhI5s948A6DRf+tIDoJ89216hy3Hxy8whSHba0TrGL1D6
d11/Ak9UzVUrUwdWbfKzaCzdg6CW9HTCYPcHC5EEpWe5Mp0yeVBCxi8Ou7fxgcSh
30k8fy56eLwk316wE1+sWUYa3F6Q3aFn1VEafUpsF/tYdxVnFOTwEdvGQpfGfC9E
ruXFTOWWGy6KT6SZsF9IZe3txKmu//pyYxq09nJePrwZo0IcP50KzYaKYK8konud
P9l9ceue2vCHESpKZXvi1r4bGGLhA0CSQJBOYA1yyGFhIVMa4gVs/Jmh58LX1NyY
9rxFIpLKhFA38yxJDMb7DkeDTCg4wQjlcYUIvPC/wTRZmoSjDmYBnmSq8xkP8voK
H2BD4m8K4FtU7L2peEL27m97IeMmG0B4PCl12zi+kCvzDc7jS0sxdd0f9uLfDfI1
LBM7i6KHyDrfiYaBXIDm0WcvoBszCHwXQ6ii2Z+6dGDPETxlgJ/W0JUBd/dRpjEY
KNtZq5pWc6i7hOrAvF2w2Fk3UjeLTDRIUPZPaIHhA3GriLalgdFNz2G40S3JOwEg
otGG+0S6jPcmCF5qtRiPemehZVfy9Aoqol+Pl/o521tClP0WA/K3L9A4deZ78XPs
drFaLlnszDcno8fUH0f7XY5/l0XlThBEp97dgzpdSYZsxU0PBjWvMhscSRp6pLUK
DJq9RR9ZUrDPmTUkn2SpzvdPAi5vtV5cJivpfIA+ssYFqBRKEXxRTHzTjiLHozHg
LC5kMbFtjeJpglBN6ygCUHSJCVADipEX5vTEOtSiBLtdWN+tqnVfrV4FRxzKyFMJ
yjtTAKUKIxCjp03AlTuaJtWe7zbQ6LDqIsUMdykL/8V6P2r5N+LLcV746q0HqIef
4Z8UlBdidVUqVImSb5b8M+PiD0ptQGWVro5UibQv34tVaVWbJ6x+c7d6CrIYV91+
/5xPt33VSNOU7gbceWGfRSYXK5jS0NovaHCNEKqeYeml12W7BQ5skNAN9L1NT6vh
29Fj3qctIljGIYsUIUGzMdWsx+nhTkfKvRm0hTDqSuONLuHOQGa4wzfh5PrtlyJ7
z6w0xda38/IuTijXzKQq9h1av76XEC0ED1iix3x9iFviOOv4rGUGVG2RWWoG3giO
HYQFznyNnBJYbg0K6KpkcYZEtnu7rSO9k6CmyMS8t2kr+22KwRZDwkur8inULpTb
0ixpjHi3fhFxkyJ6uF+Ve7hswPOUSkzrkf9yuluOrkActJyRWClRsmrFQCb3XQFF
JjiQJBHm9QKnhagVVxXdzHtKkrU5maiCPi9+zVMRLa4CT3LP9VyrQarm1CzvD6kD
vanj+hc3pv1M0oxFAaBuCzc0GRdGvXMnRCoITBMxUNJ0L/Qpzpu3alo4UAF3BHU5
fneeFp/ivB+SdCjE7pkAhb8OeozULY8GtbrL0+a6w7E2b5a6sXh2PPGTT50AwpEs
+WQV3AMNY9funRf6E5dWKi7Pv24/cZq1qH0otcFJzg6b1y6f4F9vSTCnOz5eaOOA
SE2CWPLa4bR3ejoh7g7j5n72gJkcUd0xXM7xoVv01HaauJbsjjT6HiULmgJgPyRl
SlrwNkQsZ6QIFneNvm1CiI+0wE4SdojEMg8qG7cJw31xwM/psMChoX4pyd82Hv2r
oxglfkGpKiB8FaNlGZh6ZWjlQvF2ou2pLsVjrKq+RxajMOILj9DrYct4KnFLQOPr
cwLhSDeBwDrMt0zu7wUatn/8xIzBlL2J2rT+ev/AVocGpN/WZFDmIl38HHyW0k6B
2pMFe+MICYWayDnGc2zKLCOQt/NWOH2iAi3egDohe/SRbPubN32UCLjIgATfALZT
RAp18AViR4QfVt7gjAfSgbNU5pgcWmDtJUkRAvA1HQP8Ty7aJdV/LhIapdkw0+CM
rBjEo6ZgbN6Ir7U+Q3aAdj8m7pQyRAg+aNE4T2Qeb4XcE+4C5dT42tYjptGfMBsR
uZ4N5Oi9kx+gbTJogdJwETyN04jAsq3OWGZ/R8KJC4vWK8jYPVtaWSp/zcJ+c4K0
/WIUHysijRlaFHHS9uEVcQhUYDPdEFMlZrsdZzVBzRgAQA3GHsWiqrjvDerMmza/
f9jXCM96WQg+Hd+yAf0khY/SDx5bbeytAmKr6NG8ipAsdrKWZwipLWwP+3/kWdlS
3l+Jeb6//CoWNNxFzt3hdwUhYPi3XJggKN7ufCcovs3im1S+bkCt9xvdx3lO0Ygs
nmlDflxGqJk4RJqGDjo/N8PsXGtF+K07AHD+GexgDyVFa+DWgGKLCRqExsdhtCcY
D1exCeAjPCDDSPuHMwiwDm9IfQyrtPKjlNzCKUeYZISjMYPVLlUOnbCKa8ONr+qA
8Pg6TtAhCY9lYnq41FB49PDJOgDJcMgu2sbtGuNWdu9ytM35dhx3G+YqRsbNCxC9
Ufnm48uL0uVH7bG2mctd96CJClheEUNOrob1Yy1/ipHWoFUUh37YEAE7RHgeafpr
5pQNxmGHTo1yKiNEzkGfSHOF7YShf/Ji+KXZyroUwhU3E8ZZ2MAYrKOAR0HcCAMU
uYnlGZWYYB4uQ2KHVrIldIqsmq1PrUcFgnV3qZ56RqFCyc3eyRHctFDmgtBtI/UM
nK8RCRXDQjrKmbsc/RIy476elGi7K4GlffV96YHT+0JUOLXsnfJzlk99EHkSyW+u
yLlJIGcaPSSc/t165/bilQzD6QURac15LNvSl0yHOpDL6RIwcsByLUUgJBsT53Q1
RPhNLuWzCS8CKavVK5Ef8lazYkyKHE36/Oo5YCibr6pxjQo7DY28Chb5q9MjNKws
yf9mUKhZv5ffyQnwJQt+AFJ2xjHutZjGUnS28eMoUcXrbOcQWrbH/IEIy1vheMUA
1JWUEfZPsg4lh5uQw9Ckq608BPXgz5Ca1u3ZzpJe9A2S0L82i+WQE9l7zzgp6wdl
hRHMQbMx6zowYp2d9W3A6RglsQYpO/ZIwoUeukfn67gGYGMVGhPPvO6H7LcXJ+tn
8c8mUS2l6dVVZnMQAtPpEEfGmlUKJb+b8mS9YXpiGOdJOwSESwP/uerWxwdIHYrB
IHmzBbHyQ9ixaKx+dRrgTzYvPbedBWBMAMT/FtL8kIpZbQkH2WlVZSGm9y2YZXK9
mkRoyO4uy10ubKLDBNa4mZGodeW9PTuopMH3Y4q+hxzQN0R+DVt8bqlJY70jsDsG
SWR4ggvZEmrFaQo3LHFcmy1treRsepyXy0ltWd5V1K/XfTBlcMDNafIfo++JcOVi
0Uyzzuwb6tUE+ClTOZxz3/BV/aJAah7gbGyGi8GO4nn3fvZ9DkvgvVaUJrNVWQWc
3M5raePyLQjNOTKwnMInP97CWKMiovc6jxESkMO4yjlfkm4Dbn0o4XV98iZbVDHz
N/ynjZKb3OoXmwqCN9FKKt78LSvapIQeCoMgjSpOGeLe/9lPSSep3GsEBl790Xrn
Pl/O5LcSwHJSKJCMk41Vy0IMkkqZ9quiM2WdTDNq2RHwj/YXZUxlGjd9zrKA4KqI
+TPXXmrsTgYrHH55kA4dGeTkFqYRaNZqG6QnO9o4y0vkAKnNI3rEtECy18x1WZxx
tdS3hbq6i3CMr/BEywxcqczPCEPgwDYpH1YhvPrZvSks1HKANaix9IyZCM/90pGm
TZzUZi/UpvYbeuus+yUUDEbqA/JfUPbDCCx6YDTzw5fwEBIjhPMegYblk00U7zKB
Ki7cs8cPWY8wXWA/Z7WwOwgEGwHIB1E86V8rOF5qCf1s14FriXYLwEVaEhz5O07v
mOj42csyF/+49TX7YTM0ExWUvd4mOSpVbCQ79Sji9Hf5P/tNtFhVcE5QdCDofxq5
CJAVRUWRB9URNJeiCOacMuLZEjPmEu4VxVtDFf531qle7JEYOzfSQMHzIpdAYjy2
Pur+1GPXTm2U/nV2T8PMFg7nfKL5AWbJjCXyrk7ZOg4Xfb8lnsNw+SgH23VRuugQ
DmV3CmKisawDE+fGNuYJL5UMFhAIR8tcoapo0ZOwtwQ45gYZWRUcq0oNUy6wk35a
ZiX05T1tOE9XNuXoPe72UeC2Z0qv15iDxHy9R9zsNb2aakM0Vqp02ipZyZxVk+f9
zt6fSr5QYGPcW9dEd4fRDBbPvcfT03mjsCsjrTDH591TtKqg728tLsHJ+EFh7u0p
GgStK3k/PEf3o0GjZtXpV6cmqvrysLQ1Z8qwJ0Ovd3WGwpPqjCNmO+8JRgmL2M9K
jhUw3mhdeNmblcBnkYN7vAHR9bS0lFJMgdERysRVXAl3uML3ea5YS4843rCirNB2
4awdy4xCWwX0D82QmHYLTE9rq3nvsxQU+cN6VWu+43DUAlraWdEZdqz69LMKWq0R
TF6y92u9RoBuRA4rlq9hGsiiV9iTvKqCbhendj+I88kMy2MEmMct/88lv1v6/qC7
reGwGQpjo82ttymZEwvPmFuCXA5wdbofcpiGyIkPkg8mU3kDYNChaCEcoLOXDvA/
jifR6yq2XkedR2aMZUHUVgiZhqSElY9K6MVg+YAGXMp6jnX9qGQbp8+rzR3KJ8KM
JIx4iqxS4CUQKCdhX/ETXdNy7IUjPUfbO/LBpUKO/Sgm2tB4IVMbxq6UQezPNBPU
wBQk9Jcds6fGqu8EBQ6lv3mgay3/Q8AI1SpAXLQE9h0XqnTjHnahJelvkXfLJ34r
hTy1mD+QqgRa38pYPmCottVXl9fXR7XPQyHAVq0XAFoR6BZe4sEZilUSPfy1Kfk0
MVUMUPvmPPJ2qLQvmbNT1rkQY4t1ezXMHY/1m2bGDfxS7RmT2lr46wU9ML8xWuJ4
E6K9xwveaN+X1mPqdy7EtBh1bKYJSO6tTGgPiPcbu1rO4WqlOe7E8kPSzi7VRV5U
hDk+iw6JHRePldeKzD5xbFwrO6aUpr96uSmjZDAGJe6M/EWPfRvbKpOPUNN0DXb6
UyOZZuE2bziIWSZ7XZngjMQnlh26qEsVU4RlsDR06+NM8ykTKoB/IowrEuyrhLoA
lwoT6DgU1hhOeEdGRcROzK1LIm+p36xF/RM1kGR1VK70KFsRpSEJ1OZDMxnrlLg1
Mlrf0e4ebxu5PMTybjcuAvgLo9WF7sB4HCDqEH7YoKw1tGK5Wix6/JrW0KhWrLCU
XndlmBREXrRjoSnzBYGy/tnGypUeGWQpLPxvrw/L3FXfHhG3NYvbpYZkBU6QpimX
lx6oDGP5ZcVU0netNm3/ixZvzvhZfz4VcK3hNgo39hTlQYiq7cLMu5NAM4o9jVSQ
i4WlcSy8SAGoUUZElvKRpJ6xdAk++xIY7XaAwVrC8zmh9xDzsv4M7JcRwYAtEYF9
QZ4NQGaBOUd62PtnD0DJ19ucdQUGUAc3wk8XVYCyXsh68zCX3ijBc048XuJxraR8
3HqkuHHo5IjCPK8PjqXHQCb04ZloQJIkHQ091DAB/wN0lt2eQDpXVm3EItLdqeBA
vGOhRtOqySRB2E2F1OY9GaBGWnjBovQd8ITwrb4Z/Xhb777l4eCysuNKVTyJzqiF
yEkaPZOaA1EGLVCkLLS59TO5oUniF9Bn9Y8Oi90+BahxzrHKo9IgkQGigbU4RMeq
gg7oe/ve5tkxnIjegW6F46zaKQynzmL9a1EYdmtD6Yg0+kc55umiiHb6tyK+jyOl
5JDg8XmNpenlpyOt+HE7Ch5YlpjC6IiOnGaSqfQg/1K/nXOSxpAvvaGsPxgevoox
ybENRwS67TN3Wye0Q7f9nwU5Axs76T6VVIwCMm0AKjXLI14Ru5UIx4vw6UwJfmm3
c3gCRyQba/97pqm/ouCG3yDPh9w2kmc47HG/ic9jwgYzHQW7ajOn39LXZmWsbmwE
RhozlBmbdtNWWiKktZbn8ywcoipTy9OsI8YGDV41UJMZDqrqA7FJTpIwx89jfpMz
AzE/Rb8yngCdf33JfnzvhdH9+31qJ73/dLkw3R2QJ50YIMWAakSbkv3lgPGfDmxz
kYWC+YlD5D0y0M274f4akB6LUIiWSbu4HfZ6tL8ngthfYmu3CwdLoMvUbTJWK8oB
XVa1vOkhyzDL7zbkgaGK2X9RCYm6fKsv6gCGIny7tr8KtL+g2nUJo/UYMRmvpSxA
TnhSSynsYq/ZPIZndOBS4NRDdbUHtf3Q030N1FXrTuTzdEQNmvE8OmFxuo/m3M8C
ygtoD4RblP8k1oG5ayH3mlGRmtxVmws6exGK4+YoQuGPeo/0gO0NQ648qnGPfjZn
B7fGPViRS5ph31WGivHMNR4byWqQbHS92lOX6O+HMAoRSYiJtS2WYb+ZO9Hix8Dc
yyxTDIQEq88cFrTTE8SHiLEeuD31u+F/aKr70XilZw48TCzpMnSepNO54LWvhey3
zXW8KUmtpLOOShBxcQwng4bXh6NqdOLiow24EETzstnPlC4KRQleHxn86MMwLNni
9FoegLKntTwgAwgakEjFay6qNd+LrwTp9RJ3EgaNtkPWNwogVYk8wAWLnA2pVPhK
0Xm/i/0frELWW7XWbtCYao8TCWttHdlEIKuLvjn+5J2tKsHCjEh25TFFn92GhV5D
uYYkOJdEYCgS8ZXRPrbmqnnpzrxP5mmGL7/22NcydRnXOibD7N3MYaKfKWiUfCVY
3V9R3JDau5anR9fkIkhSlGI35iadnUFFhHU8VIV2f8cvriZaWKZ8GJh46MlmrhQ0
PUurFg8Q4rz0jViXBOHx+uECn+3Iolyo5+zo9217pUK1M/yK6jMqay+vyGl8PovH
5rLWvbJdo5UQWa9BatafVVm3pTSyrrU4+dhEjJrqnkbW/l14MFJ6DbfrfNWQyplG
RRtMh0Fb25b87WjQ0EnQQLAe/rVRjXL04BNTekC+itR9SxxIleJE8395a5g/jtAi
kkZHTDVrsW/YAi8Gr3Lx8s2qdxwOkSl/GXnT8+L7ZiR6lsGB4EtuZfmMpGyGd6GA
izyLJXJsrMg0rL6EYa8WS/VzwCUnVBjQ0Ppn8mPLYwJoQ35cijlmhHlyU6zGJpGb
ISLws8iTRk7d7hG4R1p96zEueoaqC/PJ9uRUIOBKIyBdhIltefxsTjcTnPke2+aE
yEwV4qGsLSesLYuJTUoWCJvOxRaULICi7G6R/as69bWMsuogNQVw6CzYj2qTVLK1
9NM3iSVxtZ4ssWDicjVnUp8+WoS+YYPWan6qMOGNeudAROAnqBoZvaxDyakRwu6d
L4YADm/L5Gjh2knyQOEM70XpytyHXIByw9Vw+eZ9pTZ4FBveIdvlkQ8SGajLbEqf
uErv8dHFtLxcIV6OB2M9IzwjAXqqUM1+dgZ9KyDmTKaDy8bYr+dW90BTfru+J+oB
cZ+Vk6+q5ntHMImslCfcN/htGY9YARdG7qTWIix6BJN9FXtesP6Ri22IcGOD4twZ
gGyxx8jUjxL/iSAhL6skAKKBWlK8oy02a0GjYgEeTxya+sK5RXhmkudY54LMW4kK
b8w4FEfoR5xciouQbEUpoKYdEsvAqBpNZLyGbnuCjNnGnjvpGoywX6hsQCncGhSw
MYLwclYEy7PJgiuApYEo+z2cPM6ectvUJbPxn9V8EZDHUo1vhp+FlWfEsOAl0/h1
wxjtKNypKDeGAOxJRZCJjXIkuomzB3ky2QoN+UWYThcbdUe57/z99I8HTRw4AcDy
W77C+BghsQZceq1N+Vy+vlqipCoF7J9IuweXWsTKLDSMWP9fSDL2bTP5t0WUjbg9
6DHx+eLh2TC5nw3NMlBTURJAZbQEZVLFha6oE6pMu3ApNfHDmf1lDZgwwL390rqa
65BEJLfQ2/SlfQAXkJy/AdJcXT2P+BVI90VURKadQHZF3E3bhYggq9CPKlnkh480
AkUqa18eh4oER5THmhLnSpv+dP8AaL9giJwtIoHxby+hilfbngmF/nVm+Fo6jgnx
41sNVsj9jeYbB1eCZ6ixBnavv0dHD3tArEBXeH9sko4Q5oSZdrbejBFx06C6z9U7
j2vw89cEeivksvsXrLlRYzbMRaZ9bjxfVNkx9ZVderKquv6+FNzmUxo6JNvpWaw7
cMX7sDuOOVCugc93Z39GFO1HOLrv5zduSxQwOypWKERqHMjuky4TxE1pyjmROb7o
xu/PwVVUZbQ9Sk1RY3qvqymKuxqlBo3vz+ZlJBfV8+kLk3VOlamzlGHFUhWghyHW
opZ43r6jXajyx+g+IzyF3XU6e7oMwGn27bHLnKmIj0L8BW8PaxHgkySIU2TkOZ6Y
s0wTOxJTy3ZESYOz0OsJVO+Kojm9Ut1RiOK/Oy6dJdpi6WfaYJ+AYUQL05Thqb2q
SQqgWBqGM3On0tsqL7t9SB51y83/ZRZxF0BkhbQ8OVkLLeSqYqLX3G1wDM7RURyX
137cG0Mhj5w2GSgqAwb2Yz6jnzJJ2ecbC/M0uWdRNY1MPt1556T8UuIIVMaXthBn
Z9POYhMDjJtCW3jNLPZPWqeeRC2A+uwJZYh+vVf/RkpzP6FYpfotsa46obyD+T3P
PFG3p+KvAYsPvma3Rw34/q/iT7a+1nIlMWIk6944JmA3nw92sTuI7HldTKXz7BIk
96UztYkufOmD8EakMip3PyI2B67cxELYl3YM+jBddkTfdXl68CxQ+u7P70Mq1S31
Yy18y9Fpnck9TJ/UFnwIA6TzW2enmRoVEeO+51zu/YdQF8R3rd84+gs0718KgD/K
tRb+GimjRMwmWXmL3coAtdEF8PBFM9KItl0ZUqGkxynT1ZxE7YO3UNE19iz2TZd9
eqYtCMyqiFR7+ikGDNg9cswunvBdi7Kz9LHjN4mbYF8C2g3zw5bnXiR//A0SxesA
brjtO9ykFxE2jZu/Mu5j4DuF3mjBVwLEY8Pa0K6MGEcSw1MBdExz62vF5shVHWBu
ZihQ3zuePduFo1uf3hGUaELhxBMsC99LImiNayT1E8461SWYSCK7n327FmU3+1cK
RlmhcIrI+eioY76zVjMWM9GaKThoqPSys1CMDab/A7dsmvswxv2i23QBa149w0HD
t2stocJmTcUv9QmPSSsqxeeDRFq4kdIYbXGxQtW97ZanZahMrrcd34nfGes4kvvd
Qavhy4BF3LIT5Yw0MNAM2y4upeZ5rh5T94WqUpH4fECCCaFfIE/gJv2orrdEFJ5m
NQ9AewErkIcQEJkxO+HEqQtp9XgL4x8bJIiJlABUG2V/Ji8pS9ZQSchlI/QMckge
CTFkSlWXVLfnaTYSxn3G9Z5wyJqCL8Cm4HenzP/ZvbbJUliAuFotdd5/mg+fdAeq
ThizGu/i3BbaKHbFJpFR58GlXzVKVLSYODQyXv+hzAhGcetWOM4w6+Ryqe+Pi3Ue
inU+qaGdBMHIQ/EH3Q/aIIVHwOVDO36XXGNpPBMIW0/OUTu1hC+2aLcYHYysfj8G
mao7/a89/MjC2Uu1+qOaUWYga0M56Wmktb2kdcMAXBEkLjWxLr3YQnvG0L5mwfnn
n3/JY1uohlfG02plwcKAMBhG9gcpjcymWCVpt2gybLh3tLL/Eb3msppxawfdez6i
QNdXZvfs4QhNwjN4w6T9HZeazyRg0z4wtkv+Ma4h9tNa4yLEUv/+uUNtwrIGawEM
fHSht3weX/+P6hkyhs9iA1eLoOV+wybTH63zyN/HrgtDNK1XmAWIDF7/eQI6v0EU
kmMatJ0UzyqdjghtQ2J75i1v62NvZ/NNEkFzrNpjEPSavH7GbsVoMiRbLKeV9dI8
HopM51GvWLxeXZC2L3BlRB2UIqmb/WqnQqZiRdkqUoUYT9DWpn3wCvRD5eCcYskD
MkZg9ELXct4QUvQdxiOphohuhyv/7LY9IFsfqOdUM52QXomWhmwXKZWnJ3Fc4i8+
K0Mc71S8FA8fDoomE5PSmpnRcexsHeyte/1WS7/2z7pbOpr/KS9drb9kaNyGbXu7
dEBDYwPDuPWtOP4i2Lvo5XOyXtHLYkKiPS4sus5oQVjoT6TgJO3Riht9yG7DppnJ
akCQo2qpfTRwh0aczflwQSC3Sx07En2OWfObLTTti6/SicRh4l0ytwpbMlC8kNiq
/iMzJZ0E8bzRzQr2xLcmMqUvFE3dr+TA2Ta/ObDs3wI1RUDeRJNDOafCvCkpLK9w
x7P0dDs82FfxyUNunMZZ0R0z4/MpjumvDtWAGdJb7vaqMfWQL3kBdlrlEd5XFtTz
qzZroTgao+IAqzVFho9fCNtjIt3qT4dO7dLk06tXOzgHBeOsY932+0kbFiDxCjPM
n1xvNwsfPoHpLMrRKpSkyR7C29xVdAQW7csOJJMyDFGOZ+De8SOvA2JohVXDtgu4
QoDA2FvU4zDQAz73Pu3Q2/qF3DIwFTV94HRlvsFXAJ1yJleHt6yYSxKZPGV9ncf2
/IrdJCb4ENnIfWkZcl61PgwbQGOFUVHX69lEfWAuwOO60a6Hip6QygDhAofGZYRi
yiZfqzi/XSYj3L3YaJb3UyEBCwYrcSyiHbnyaNUApeZw5xqziJVF+xMa9yZNuAkj
VsJYcEMyyqoHj1z22oimR1X6uDX5IBp80JEQBVC3zjPppr8u/JAVVppklNqpmviS
QU2+z/fFhoQ1ZNATQGGn+JZByKYCLFepdS2DUPI5+rck3m6sMgyNWt2WQVmLlfr1
2qhubR3EnAAR9SRciJB4kbylcBynDuN2hd3yIPo7vuUBiCKWamLSNCN46pMwl0NW
7uIgZO2LKjStFKJgniPfrpZy4Rv07aulDW8TiQF930HhhI+9t1APEucMJaIe/lgv
glmWdjce3G+5aH79GPlCNjKxa07uogov4zIoslDLELanIpRbyEKcaAP4kOVthU7d
WnEq4n/T5zHx1wGfzAD63Xp/w+5A7t1qglivjdbCr/PRvhTsEpWQvR/RALkmj/3u
NA/uSnj5rfN4Y29aXqNz1ei2yj6rfe0EjL6iwpoZBNmd8++K9B4epRBFclgsoYT/
jnLxtsHvqDbLSTEbnVumM8a0yQHa8k/ZOWPf96uks0BjmiooGVFb6lH/yQQSuXSi
NpKOXM43j/fe7LMxzc5IME5PTiozQhp9GBIvgNZgCy9JTYi1PB2kQcAde/oLyo2K
bYwHaEZZpHtSmQMpRpQ3XzRgK8SD9P5CItT5yxa6k45FH+jefpIgbBeQXqRLKmjr
E7FFXZ5CNKDl1noo8XhEV11ghry1iGZQTwTKTy17t0nm7fwYToLQT6IyOtCEl27O
pAQ4DDdxY4oZfzgEE20ORc874kUNvary+rTQeKUj0quUFXacT7M2seRHkkAsNOY6
dGsE2R4IbiGvospM0fd9okiOnpZTRKFpUtsFkY/sIPgXJLGL/PUl2ze0+cVY3Xx3
QbNqXvFrF807AfZnbLVsLiIdr7c6GNecOdyLDb7u6CwiiBy4/3cu3kSH8+NbGpUL
uqqO1w3BbBCMpVyhdEyiNuOUYx2wguhOhp/sWDrM60P72OYZKuhTMX4ePoDgluev
F2HPmbgTEdGg957MDTdYtxvJXUtjSP9Yh8KQh2HlQVCdBCNRuo72woGxNiRTaAIp
nXRQk4VDECVP5eTbfZJ2Fe9R8XbmMBN4diuWFLVCUmGHpIE6gQL+9nUNfnfbU2Q4
lrZH7uHEk4q7O1insUYXU5ASiIHBqliiUwqk//Hwi7vRaxKUXa/k/Yq36c7gqOgH
6hN1iGP/M9SGlrZt3lS5rxGfi2ocuBHiiPaf4hCFA/tXbQvo61pYDOr54q8szrpx
jQBigIuSBtsXYhT3f1rplfOWx1+ZzEv1gjU8HPD29EeTierpHGi/bkuRu8mZT/Bb
N+MBbGGERiLRFcXBhUogkTzE3ZOTvvZB43q8B5m+zDmBm6uNW0jjf1JQ8SWEG4dn
bypwQ/Sgj0GSfZ6LTpgSHi9vRUPnHHVQQoGcaZ3JChxEXc4mdy1XHSjYe55fYcW+
UY+TbMz7SBM8ZTMjK2ScA6lpuz0jFmIKWDiX4K0J/A9aYFpKJad4aKQNGBmpswqa
BLznAjM/Bi0GAwFJiz1AcWuV5FRsupBkOwF1F7IYs24Tjj579Hv6lSi2jSPIAhBN
WXz9HIo5DmvJqeACTiC6C2weO7zO0AjYkyIh9lhKitKxU13MWWEIBpBUaqqvdKCW
t8sZn+XawoNVhq9FjkSdfCHaouHDvIGNoRutRL2ba0jLE/Lo86SJMwEDisMQTm+d
Y99cVlBI6392gAUIenbelcgxy/+YuXbrkFZQyVhlvWvLErcsAP0+2VdteJa2F9CU
hAYhkuVVR4CfZNFXlcrTttk4SJqvvnEN9L4+DFExrRfQYtvmfK1g+qyGG/b+GsSw
9XSudHeHmv8NbOe30XWRSEZwmLn7lVmnIQ8yQBCgG+17uWvRUMzskWejxvOb/wUf
vdWOIdGaH4lDb4GNjenbUQSU1AMhSPzpd+VYj4LoACGzH97GZB3Q7toSghkW8C7m
1NuXDMitNlMFVqqsVXDjw716N20j/911XYKhY5XeJU0sUZ0a6c2F1XFYA//F+FYD
Tqou2ugfSsd2+9qG5sfQXtiNGQfWXGEX0XKDpReG75ENmiLsBwrMqFiJKfAhSX7K
2vn+TUIITO4NcaXqRGH7zjJYMpyf/ugOofvhSGwDwtL5dV+pReqr03mmQXfXN/Qs
/PKIIRrroptsPVLHXUV/XlO08ez7MCez+UolKxwoZzLcVN5kO74EzNGW4crIcZNT
gD7XyhQy2WsHovpPYJQ9qz44FoQeeTLHdOCl6GI8YNE6PpealdfF/K69Aea6VUlN
C6UtuaJbmw0TTBghWydcd8sj3eO7HKVnlgpklu8Ljoda2FfZTJIREkJ9yRpOfb3P
cAiiB6lStX+SSWMXZsDdrkHDyuAVyOf6QB7FQPMYr/6ccFC9xbB7xSKC5E9T8R+/
AW1leW3CWr60/8uOtun0cXoEi3JlShP5j7AKN/o4FwQPoEmqlHzZ6fTd7ro2IOuC
QVvuTehtZ9Qve6fC0+2czWVfjQTB+a22s3iZIRNRXlrLbHdJFUtHGDoDuY6QnFJB
NWbEJnj568Z1tZaPaf3wDu4AHZubJT61bpsCjdrl5TapVI2aaUfWtDgYa1P4hfI0
erAhhyJBroCTpxIB1/9p0SBge29hyXme+11Y0nsOynOn/H2jjII6D661d6p7UR1y
Es5r0FWIbXFXeQaqY1Vq3MfdfbOoww/omubP9A8QbCkw43Lrgsada6LJ07WzHN2R
SNRVCQH6v9aMMNwRejI8S0MKdVJuJVf6W2kVPdstRWUkGo2b3TPp7fIy16cwNYnY
cjn4d39KvisfTq7GKuxlETMqvuEmzSYwNMpMt5viH7JxFBRq5UUIeY5/6iVuVy0H
rb1cbvIypGsroZNYZYHc/Cd0LwkFTWK0jx/st9RzaDePtRSVOiUA88YjuVetWfM7
JlFOGZh3wRBSxFSoRN87KOCh3IcsZ0TKY6+4LTfCCHIc0Ce7HR4GDk2dzaFXUpon
69QFFJZJozVeUs9/jOxbcdVgAeRA/26umWaraOEcpDRdy3JZkWAS3+lGya7Zgw90
zIrtjvlGMnezYUTo8gYzCIxm4F5ZSiuhP5dNldyerjQZd3nQ/66LSkxEk/IfdSZe
8CwTV3H/QS7bHx9Tj0fv9JOOx3SvL8N1ttXI2Swe8S7CmDHLWFv3FVMKkIIMgTI6
FpCVnJrSQFl7nKdqyQPsawt+cIp9OrYz8KG0ozMQa9lP/6RLlfxu8MIN2VkJI3f2
RRBPeHAwFG+s4FoasRreZfmc2t6MRh63W+LS8ZaR8S2u+ZNly5J7vzNE6x5V6mRO
FG67IFQz1TMwlcEjrUyJAj+J8oya8Sm16jhCnMIDpetc/94Roccp4rUYKpHVKYsA
bwIvK6kriBSFf2Y9Qsq2CpVGbf3OEsgPT4uNRczpu+ZSfIS63vxwYDPJ/AipYUuB
Z6guVn1NWq7Xqem4ROqy+SI1ln0hf3vfDQ6EBbtxo0m6Rva717PsgNQqiQ4oALfs
/vKxRITM+cY7D/ixjhd5/zzXMNCw6aNcZOmYdXjQs6y6HME1D1IKiXiYA+67NLmr
fug13DUoS9xUUXyubAkCxDod8LSF5CUbnUBVM3giaKbweb5bDjK8nOB3NweXj/Uj
3sKU0TnnWFG//DlPsvgTbod0cg2hjtbSnYvxon8JMQeGuwyyFZ7LvTjV9Kcvmu4+
dA4OlPFUShP4wj9C+J5ESY4lAFW/bQBGd/zMX+Trx/pomxLkRAe1SJZsc+Im+JEf
pgDCluF/kPKHGU0kS7hqLw9T0IVcCWhgRJ5Ev2jziqt7wNf1TBb+L/mAoRUlb3lm
TQD20hiSNm4d430mKeceNpXdXX9mJsyq1RjjxYlNVZ4Af3xq0RAwhudnirCFH+ea
Du04zVRGUhe4LJF8v45tbU3GOEGSO5dz4+CavLPnxi1n4Vl7PSf36TgA6mV8rL70
H0t913A/iJxib/RzhSFWV0Y6lShjXPRriiJxy/RfrsBb9dQBrQWlqongGw5jMBCF
NW9Robd45yDGE5v0IvW5Enb/thsjdEEkWvVSPEx/EQqW8fNZco3WkP8eculz158g
DnXe99qH3S2Rf9gOUzr1gWSkzIixBIVHy35nZ/R8MUR8SieQwxndJn1Evh/4RMYO
cYqW/f2x0JdkCXaPdlfsuRaZtEmkt2EE4/U9hE9rqOPrOA9Zs94/mrlmL2IXPqOY
JNhlqA1p1hlap6k63a5tyqf/yFmEOOolmZBSNczsUm+H3VQLCeItzui6jDZQM76b
uCqChMYtNv36Tu5psEPsSTFVc1UWcFS5ABdJAzAqTZvp83DDbiLaB0tg+J/Vyvfo
/IBNYDkjYZ28kLW51hVTl4MFT6JHNSENoe7Ryk1ES9URcGxT0Eh/694gNLsUY5S7
rGrd+73C735TxQ4PxVlg10sDOpelfGww/r4pjGMjdFFmP+IgCQa9+PAGKt9iY+o9
AUdv7Gy8ey8UuKkqGe1qZ/tw9U61Dxv+P6A9AEQLOFPEnUvvsyILN8VKFZ5F/Etk
gRYZwO7qck/PGwup06ueWmfcrqmt1S8h769/MhNyXnyTi8q6F3kKOOJFVwBChcma
X/Spk9gqVezTumYfHmeXf0ZN/kCfvVc4XNl22bC17PUzGx2QZK1fytZWtTFZxyXz
ZMySTdhH0vb4mmF6hgr5YLhlzpZfaAhlNvrNVwzPrRkse1G+OUrRUpf/9uPFytjQ
qJc0BbnpOpFcz/oh1918V6f0V8cYGNJ6v1Vt7VfgFSOBgF2HzAf/ni/epkLGa6tO
bd0SVgJ0r0XF7y66ZibKoBJEZx5lG2wq9xmhUsa5XjB/a/OoVtzt8gZVTaJp4q5a
WGqcLQnOzbSml/qNMPhELV9GwiBNZ9mN0kGWFHbBs7jqn/5OBMX7RKomTDBNzoIs
MGLxOuD4x/CkCLlClT1Mja4tZP2fVDY2zkuCWISMp1MzNSVjZTrApkaOlZm1MdSd
M/SPAjg37kN/LTtA8m5Iv9eW/f/RNiA4zss+WJTbEf7iMpcd5IQWItV6Du8+GlX0
smX89ecgava8S49PBOdsB+TsSDkfkbikagielj9+krI2Ged0M//nf+Qq0QnwvULu
zzHlqfHWq4h8VM+5XRU+HRqt9PQQgnbihBMQllRz3+vh8dSVCwCwG1Man5kzqUJv
NSwIiXWaV1dsPLlw4fFXP0uVIAAylzG+MvIa4lRceUCC4+yUI3uj+QiTiB1g6OlC
jidHwZVgdMaehigwnscHKdHDP2KZhtwLunf6oN66VubQjN9MSQ3+IteLUDS3b92G
YkgfeNuBQTl5PFTyZn3Vhh2ofcQxX77iHTJeIopOnF0/zlUin44rz6nGslYO46g7
tFdVMP89138c9S1IZx6bbZhDVyp1u3cFvy8SIALfFz1BbpG9nfRgOJNLuLa7n9mw
IiyC+9CjswcgIju6slDT7rpwfgA8GoNID7HT/VqC/go3P1O4FfFd9B2RKNTlNHnM
iJDlF+OkiSnwXmhQsg9F4jqUBMhgXBCvlMSe+LsnLwhhuWqVJvJjVPAVmvWJEV9E
hdHimid8ieXz+GNDAnWukLZFMWQGM0FW/dqmRm1kadymxMhG9GnlhK8bl733ahP9
znD6BO8hsIhLGkAKrpDq31tNnxvhblecAKIcnQpSsoe5NBF4awm7XgExXFOzJEFD
HFASZRir7W54uIxBdLZkuBFVYU0bRGfO40Uk+61uMPAqKzXDn9FY0kyKOLe0Ff2K
wNJVAgNoFTZih3LNndATM6N6y+YRFCHGnO6WJKSs6SDwACjJCBccZFdV7lGV1Cyu
aEMsWscI25vgVUQtmuphXTc8q8EHJvSCMlJsuknJK6qjezccY7vIQR7RQnv25PD2
O0RlPuwGl/I149BEw5KZSD/WKLE034vPrMj6HGPKQQIi238S21EpxhZTj6BzjP1C
KDctQE8z3rQ112Nw+/ZgiW9PgtK2/SmmIBnKwgituSDCaz0IAYZj7ip+nXMBEh2W
MtN2ZHagScMeZgZK9X2sDNDPYr1WTPQxRj0585h4gQ9C8/E5NcOH0lxuKMycuH3M
uAFYsxoEHhUoLW+Cy2mha8M21qrvbwfiby3ktBIOON31wv4+pE2JdQE1se3EFRnQ
/P28yk89/Xw+mFMNeQ6Q1fAs/ZvDYRbBZhnPnTEsz2SpJRd4JFjaSB6j+UWYEC0d
V41rdWvst0/dDupFdvxh690uOrSLCAMiY26oPb3sfiCgDw+EYEsrSRDqUS+zCyQy
XhrUgATDfQST5Jc/luJmL1Ex95m5bNpcJJPJi3ycumPMfUrxKBNY2z+SXFOA49+3
S5W4boH8gW4iZYkApGjbQxrTmEn0RVAUdcu1xTRXS4XIWBxdWJxFRlya/hLohOtZ
xbHXeHiC6hSaphJKm1K9/SFbdEKJSsxERiyup4to4pf9VxUIKJL+p9RVyI6Ot1b/
6mV9WQlHU6JRwA5bM8DqW6kAGzHaAf0wsaEhfSAcggQeWN/osi6pYDfGaYwJdrHY
FX5r/VxmWITOndeE23miy0qQ6xlzRY4ldLjkjGGyRnWokRWhoXU3eWwfQMqkykAz
PJL+I09HSGyJURCFdUmwpR7Nwy/5n0trRtjteziBg9pnh3MKGxJmJ1mxI0ymkY3b
lahHc1woiefu1WbHGujNZYOypLs2U8a5DOWWGnMcNh69pMP11+ESrdIJJMG69oXr
bzg3pxLghApqs2mltCjQSDj5sopxi8fKx65iy0E0Xg2hG0ogHnRQ9eLSJpjTZ9ZL
Joqd8IAP7CLAthSblDA6sOnHSTNn+51U11D58RJZy7WAzpy9xw6hMuP53sQlC4a4
qFNz2Gai+pjmtsOk4QQtJEtnvI9yCCPiGfrSl7eKX9o/Zx51jiJKxk9w3eCN/sX9
ICckOy/m9hTgfN44zZEYRjalIou8ba6yqWbqjt0roWFtYkVQETrl3chpie5EBdwT
bsd+9skw3KybrISA+UkyTXPFCUQ7PMdp6vPtMJpkrusnxdWpU9ZAPPBXRvsi1PLs
bu+u+9F8dq0UB+P2jBO+clrVKMZPyTZZlzstD1AqwJdBJTMkwDkdtRQLtR9Vt5OB
zgMfa+LT9yRKF4lMM3k/12QQo0byxGrx5CRaIh3Fx8UTfNRx72YlIn6JSmC34IQ0
S5IsbglEFzqx236njmdzJE3RHm9AzfAskvl5XsSOFldvqEr2/ciGtRRF1vOC5zXX
za3a2DILLRDYbACnL/xNHVVjv/vkn/MIoFe8ERkM+7hssVbNllwwIRjHF2D0i4ff
WQ5FqLJQp/7O5RnJKfanP/eMSZNK7fPMjttDfXCm9ZMTs8087SOqSbb9hkivvBv0
bGHz2Z5OeuLFIJPnUnVBOQJfckaO9+mjSBSyFh6SnKEMzwhQTl1oxufjmiJmICmi
Qj0pgahJDxO7C0cWfPyAEu5Xrm3XPHE1pZlMImlTnJo1feD6vUdM60uEEBLaFOtw
SsqzQ88JoW/Ynlg1fHlzz1HffBOir1mV+s7Gf57tE8xUYYwCGorZwELFoIH1c4cW
rEag5sr2jTJDKCgWFW9XjPr4AE3TPgBJciY300wQV6AMwuYaCutFuOcB5MwB/FWz
Tx7f6QgEHnYHt5hWh2GrSMwOapF27MNb/g14cz1dRFmR43iTWYlx2gipuK4+ozmH
E6y64eNgPUyRr6Q3nEOpvbCWrzYVrPkYBxRTN0YoIsNubahiLF2qaLKc0pYt+X+m
wd/VgJ8dOLRkGo82FkB1j7z4fQoX1hJcgI1vY1x8D7TYwi0uF/WGjGxvjjbpEzMw
WIo71IG9rSEl7YOChQcOJczPQDwjTEnQr50+aItURJOFxUUz0LvhLHsXGtXYQK/c
MGXvqkXIIy9Qkw2zhdEidc+UVmsNh72qSoj/IqUBGFoV3crf+zW2E15PuIr7E4zy
jPZCPgC7j4qWqWS/4UhIyiprmZfTzkU52gLgxOE1bkOustsXMISl4HDdVFkoRgdU
QkbxR6fvODpsHhPF8zSgiVTbj/LA5zmIVrGz3eJhod74hLpoERV7tt7U07ekCYGB
MrUGrn65+O3hpx4EFutENylsVOZ9ZxawZj8XBFQD/nf5B8kEE5X05bY4nAO+1fOH
mEv2V/dil9UeIyJi8XzbX6p+3KiQtdpcJNc6e349krkva2p3zFaQAWvZyY8ORmu2
ah7y6db3PWoXtbeJlQbRAG8FhtIC9b21Fq7Plk6tSfSiATochQZnQ3RKbV4c1ekp
eF0fOxC5nW5quXwhPbEJuya/H8Ui+C0TXLNCKm+l/BbJu/myw9z8D3WtZwA1W/Jg
NVBpstSlN51q3++spP4NNQ5/+W4yoXpoMADj9WHp2oRpQSOmKaucBcLOlPY9ke4c
w7IiB/zBqfV9By33IPEneKsjuf6qGGWg/gYhFikQKsukaBy82vxOPaUT7x1Gp2GC
FThXjqHjpkg87srYGM/zSu/WB98GPHALUjKAnXpaPM+qFlsURunFns8/NlYUIjyO
4J2d3Jmbwh7wIsfMRSy8IfR82meP4hAuagmdTS2HAmTAgZUvkplVR3H8QdJEidq8
KOdqU5BiS2Pu17bxq7l357mZZp516AsAx0JQaLovnleaqynEScXrJ5CdWp6qiMJG
SmJbFG9Q251G1RazqY+M2Ku6ahkaGLro49OyAOi/0iyaq4xWYxEdnQuBrT+0t8Ed
URZV2PbEMHzOlkB3g+2Ubh0f2LDK7UvINMbd2JVfUsjf4p4JMCKKPS9e8D8/I2DM
BqB/spVVPxoe2UEVN+f5Ke9xl5r/hQKtUxzQgqqy+s4tkOIzfwEatALU7rwNA+0a
rNXfAUovTVqyex40DtBcl6R1h6Uppp4Er+U0u7n1cerprzVgR7VDMJ8Ie027d4d6
UdLiD7i+k7wN3oYV3rnOLzZ23VuuXnICxmVaDTdsabIkgD12p+Kobsd6eksdvF8E
GdEcnjPU2Polk77vtSwXQI84v6RRtdj6QMI4IQHATO1wPtiXAH2aVD5HY+0bS7vP
LSV03y+us2Gff4q4zwwrN7+1ZqQTPs3dDdxqL9U1UYc7u/hzVMmLTufmLvJfjKtW
SASgbA7XaQOFP/Pt90++SLHJv2rO9Gyuul7ajpjLlajB6puPrxWzpXEkKIImJgB+
C2SuFKXGZZwfpHCetGxQ9RuuD+AQvhgoY0MHs+djfWCd6+y1SfLirhk+XQToK8rM
dzkh3YdEpX6aoUzqejHcaZ2LeidGH8dB1DRq9j/QPvIq3NTnbblya85InzIQthte
KFjQ4YOagP9rrRDZk68q8tbWY+UbKiJPI8MjJ0GUZWnMLNxMXEbFixOYzKdSlvLp
ny2R1ftdvEYQ4XALHxs22SZxVHaRI/Y2slVHVBpftxE19stMx2EY5a5641lfXqaX
c0Dn6cAwGZy+rW+0mLeH5R6SP/esRAetL0AMhR6WUFKT+FGqzDZ1JvERV+GUpC7G
NT9Xn4KYB2tk09qLxQ+SEmLIQgvqDHxUH8ylDL2OlHNZ6OQGdxRd4j32rJh8JKTo
qYl9VGw6hk7WQgpLTeMrsx/3XNfN+ayFWRecApT4VzPK7kcHQJurM4d16xOYjNN4
I6Od3A79PAwLmVToPJluvb5K37+jUXfuN0vQSuUqJyEObUA12Y8uBpTY3NJIw970
8xLyhOWfa+luTdPO6P/G1hZUDpXNRAwdgA4ayhPyAVE+HdiSAfp2FpJ+SpPZ75O6
PUtrTVOT6I0IOnrOCYlHA/ZLBrjasTT56zV97T3AiV+z0g+rSr9hwLpQt9UnAJt7
nUkduLlx5t7ysAARrro1qfjFtU1HZgwDYxyjvv+9qy+Xk74bqcuR1dNcwl5+DeJ1
ggRGvV4XM8kThf59sOPTGbeu7CuBiYushSNk6dB4xWsIHecoU8/IKSgsKiydlMi8
57KLsEFeUwdTFVev4T5l01JmQy9MowDoGTAYfMNtrw6W5gWe5l/n4CQqyH1fARCV
YWPTCjvr6uzASjoFP76hd/aROWmMTU2m1LBTc/R033CEUGr/qwxTAEJs44Hcp6uX
Pw+DyOMszUlyFSqBe7vUVH5mMhDijoBMBVJUETGypNloGsDbm7F1CSLYQnLJJ6+9
4BxeZ8QlrG67IrTSSv5JNnTTWJqAfqFAixOVsBAAZvHeq3LnUe7daDjm7GOr7x9i
93ASx3ko5R/UA5vPQuoAXrqc5kEOyNYQ2hjV9qDIXvG2V/JhqjEvQ7aA8q23LQ97
r9i5YnjdVQ3+/gRXqRK7IKQoGVtJmnJrgp4V31IPd97moHw4QQH/K1f2ce4CNQJF
otq7iYN4Sy7Tg7vwfIXh+MjvbHnqAQd5fxTIyuLr/IvYSTsrHC3HFMM9kN3h2ZD6
lVF2NX/AE6XMIapDv5pYwYHSerAn1QjTdMo0edzOOk+7tvGFDhjw4a9Wk+i8H55d
ExspzmJvKY6QmJEk2ENsEHv5kyMKzgf59RLxxtIx9DDg5h7agJkHrOCm6BWvPO1w
N92RNKJmFkd4byE7pwlNSdEyBrYblXN0uAWXYoOWgUk8kJkgBaxloTADJtiCNY0X
budHtFl5RUZKxOcISVM0YuP3zURAQxZl4G2TNbA+jgSOU1e6T+8Nw0/SRhJ9qJBU
/FAVNyoT+Lo8GEQJIkHXEbBcexmxzy5L+lrxtix6DD8KTqE9vgwamz0nBMgoLgw0
D10pkoTnnbTaTItS76rNU0aYdrho1K8UE23HvLuMEPcu08wEZtLe2Vk54ttDw6k/
H6nUjjHyKJgQslv7dW46w6G1cy7mkWr9E7wvdUqVPCnqb3DTccZQXpo5nRPzwpj7
7SSGvp5+NzcuxZ9+rA1yfhGcuu8H+WRfzpy8mS3oSvCiFO1idrm+VwQnm+b/RWcV
n2psoUCRLOImgh8hFch7r09W6pc90boCUWQB18txEKv6o8EmG+9JvpTU/S0nbdI/
xVQPoeuOblU/iHeTMfSZ80YvPd0++UEZ11qx1eh1E60173yfeJobNmJLnWsjv6cR
RXpwAZ0HUvsEurm4ooRXEZkkc09gi0T55r9sL+LlzYZkpi30NIDOqcuBZP92SSLb
CTYe5y7bZdtnLjk4mT9674URxPRmTpgLHRgG6DPuUM+3LD2p9QlUcw5SGRkeSjGf
V+NSL/DunDM4fkkZL8ENFR0QVoIlsB8JX5Lj//Z+7Xzd9T4GS2y3o25tbKm2f5aG
nsXS85qkpTNbTGWqrcjC5/E1/iRHFzCjKvHQxHks5cyigxRAbQISOw1cYHdPj54d
11egPvc6Frqc5oAqYlsJnvYGOANf9TJ+g8DvjV6ofJvIdRX8iG5e/zhwoWahKHZl
PdQ/bw8KGIn6rTHNbe3V8stqawawDPIVpOuQEKSU2q8gomGK4SC2u208kA4ABigf
E/X0nRZs81tHUu2HxAs3+2+A9knk7P306bFjqktfBs9I2di3AyXt0XdVsgsKKU4V
wJ0DoYPHgAuntl4FWNClk9kmSwdsPn8tbyM4gtighYd+agCpQkCywrYVvp9N+tTv
eeutw0E3+q1T2IiiWrtmxzu+aOpnLvZdcB3U8S4pyoCknAXmyF/5kCp01nXDtWiK
0TbUjXqGII1nPiLPBP7zoba6AKMHtbuZcaNgLWGn0/ERYlh25/LW1ON6n1vhqRYi
vUTbIcQtazZJILqzXIuV/e4egcCosamPPT5u97XCv0P2ySwy+ytCy0lrk7ozKHpH
lHVsXPEkHtdvtLEoyi8fGSOkXAqTLkRUfBkiTpkR4TcjvgW+vdfLCD4xZkXg1ADz
kD0y/slXuoMMpC6cPpHA1H/NIRfiqAWGuGRee6Rcwzc4yOUlAIQcU8h03Hsgk13E
lxDvU6lUeVHriiPD3hFlL9eXi/3mfS9C/3LOOVfXuxvRVh8rIHb1vqJ7N0zHfagA
iKi67GHo52ce9XBsoxLcb/fMHSietUak6s410OAULOC77AYyeWcJ29eoyleU1YS1
ZYvvPqV7dxbbxw32zUsHIc4fNy9iRhwsMxwaHH0V/QAez9EpYAIyxIXwc8l5wV/6
UcVKqEaNDGLPxZFzNGk8xkoAio+s/Yf+0bz5YQ/CNOBi2wJxQnJ/8Ju8vUea2u2V
xj8n7ImbfP6MFfT2OkI8s4jMC90UhKXFYWI96kDomfDVRUaZnCM68xgq8zAluAbe
cUCWN3p+cMtGStTicyZEobvVVhj9nybkQCRrzYiAVV4E+Lt8zr+maRkpBTk2I/P7
8D24Jh7Hb7xNA625caTBfeqwilvKvCDCJPzjJNB+r1e5bnQe7Z/gSJAz+o49Dmg7
ilFqJ6aN16xY/wxpWhpfxR5xUeaMAzRUfH//90+XCrfB4BNybXycIgdHm6IKBov1
NlsGqmaH+ycMyyzZG1YlGP0icECSv5Yu+Ik7GmQ5srccBcGb6j8r/L3cDcTg+GVc
CHlC5b1ZPXneKPzIo39ULRAVkWsOVISfPhjOj6aEMplr1CHQ8YMbLEKI9YgHeeEA
h+6p1NbEnvjJv2/ZgIKx5K5ujA/8IFowI4GA1+wXisoqunIWUNrKTpgTH9msgOxS
FWKGNPy058WpcxL3CtnhMcQF+g6UDbQsUHeqhvwO09ZR8LEAdwrER+eCgMnRtfE8
ysXp2bMG3Og1DDDYV2vMOIFhexCn9ndGp6ceWxsh1/xBNEk/9F7sThPCyHPF2jqf
aNaHs7kPIC9YzHm4IQNPyWOBv3LGCLmqAHkkwidLAQOz0WXGQlEgZTzF1BTB5wH1
WZB7yro2TI7RvRLgcoSysF6d7fFUQYIsXDDVuRiN7RxPp3hQTQROV9FdI5WFfgSS
sWrEu+4YdbUV+TyfNiSE+9oIEAu43TBdUieOUMQHH+dYVume1kKJU0/7M9c+/Hpk
1O/N06kLomjKs2aO9CQgh/XOpQ4SVJrIGyTdPl1cP/Lv/7yoYdChkJjiUL5CWLBH
HYIUE8UtH08gDc3yJMRW+RwNhHdu0IcYmOU5kHWjWV3D6I6zbHiMs5MJaS0hVCMB
ic2PfKB7vA8dPZCFes9eZS9FlBMNmW/IXj/T5dHadrfPGRqRnVC0t4OZBq/4mi7Y
pFdElBFVPOGtF4g7+Qbqe99Ae8IhyCXthAIAcq7prXBwJ7n16DRnA2HMD0SjGzCu
ICb22fmulvIeq7mkHMGYghiKX0mGM9tm1Cra4JVB/WRD0wkYSz8BGx9yG4m7VfJF
qhT0H/33DaxtHbYz4xGEH1LsA9G7tm01kbF4gWfIvS35qaeR1RZ6O+r1GMM1bz0l
RrTr8vTXSZccMAzXid+nYB2wTwT/PJNX55+/L5h2GdfjISAqiLcLL2XQ4TZ7y5lU
H62qNOV/mhz1tzfoDpqs8Hwn+TzjD0c+kOLHSBhaSSNt0XZAeTQZ/pBkJSWYGfrv
caQsxUlRX+1mjGNw7cNU2pVs0uKXIC+OHzjpyvAAXPDz9ROLkLEufcpUczI7CyJx
Ix+hVTyG51wWDiz3zZcF8ZkTDyiLCBUJ5+dVuDDqwrqz05HLVJSPgc/jZMEQZiTy
I4BUBUZmOp0ZTR+dmi1sGOWh48TxL0u9y0zz0dkTyR6lPCWNGlpDQDfqMNFZs38Y
V/o0pYBUyPsjaqoesxwiDnsoymLD2iG+diFO7b7XL1WMJtk1Hj+su8SyjuGmZCEg
qtpamJunASgLIQMfY2o5GZzdRMyd2iSk2Z0LG5GcCEyKRMfAyTJUeg+r0PnWhHOe
W9L0wG5NFAkHND9YLD+vXhCf1OXsPlhsu3e52k9PYkSdVJpFtE0F3D4qtIBRwilz
DizG+Bczd3UffVDL2/fh3WwAl2ixah5WkJVPY+cCv7kaNNeARxz8aMpe9GbvL9zw
SHL8nnEacdFdkAgqc6hDuVJtInCWKlyMVgQMKjbu00JORvSWXGZ+t1nSq1HQ9uip
zHspuquNO47D2mq8BG2ONCLs3L48cZYfc/mYYIYP19f/xJod0YJejXSpWHDt7Sxl
oWVn2YLfzvUgx5Zh4JIwgE7ckiimIU091SREOMktF77YzFi2j5S4L1dpHuasr5Dh
gIapQC2waON6luD07agCyUP6X/vF6AJ6Fl0uMlsFqZyZhGtyZppnmH0QjQyrJkhm
4zBffJkmSOs4UnTO2loAm5LLincHSMoDN9FXr6sE9yVFrK0VwmdtbX4/7nC0eygd
RCOmhsXYTALdnGvvasWK+Zv8mvkNHoUEsgTO5/U91sGcSHFKv7y4wzJWxlTeNqL8
7+bDiigrEhf8v0vi4R8SLJAIZpHeGDC8uSuQkFrpErnRnrmmCDkzcaZX8TpYCkZh
PNxMkObqsnzxlBrGNA6pbual1OCjVkqzHKOxtxrh7pLA/Vr6zKhCBwRzRZaC+hKk
p5TT3aBiPTIaHPtp7gReOMBz2gbD7JZieA/PL12Z1enDHxVtERtsS0O8pxPqCvU5
Qu9l4LsSzQLhtYA/2I2cdtB2IzL5br/RjlGEy8grlzitCuIJQJrFERfL85ofsm6f
lqttfYISITjWERLu2le6OfLcF3gcQio37hhxaUBmTtINAezmQwoZ4CVdahfGLCNI
gRoc4/SWsYX10mf/CpbnZLSPoQ/Mp+CYDUqTnjg3j6J0i1fDujw5xD0aJsFtrs9H
0Nr/mT4Fjg7Fhry2bIz0f0NiemcMJ9Biv1uVrGhHlb1EDrNEyKT4CITwpR9VJ4S7
obVmlijrABjMRyLOSritvKk6fWCtyFFOWcukhn111yhXij79BEmkk8kv45n1zvKK
tBRvKLAzIuzCR14uNqs9A977zhOuceNP2tqfoZuyrc3ZbgmnbodkcMwYNqpJNvLo
aNyrhk90pCZmfabVVoYMOVoL6hsRhTBRwrjHoFw2iABibIJdlykH1SFsveDxb5Nb
M26UjjBDFMKgGiTGPBM7KClbb3TpyPT2SbhwFbYun2h9EEDFwXY57er4xogaWiEH
kBKUPvWjRfEUkIQpgGY5lPImlDkoP/EzHgKQVbwiNrwG5GxWl0rA2jD1zaQyUFe3
3LIOTjSLFOVFTAn12QS+UfEGiWTzrS0O7WEIMX/AU0Z5k6kWQRgEk8fWEF4qwhQo
icic8PoSGt9eFwatQRy5vtIKunlQNHyIM7vzHTr+KcWBf9xAMr+HHJhUmXHZ8qAv
5ibsudQPifTOwIWCIaUqOa2lkQmCMx5yo1gImet7YqSzqa2jXjNIoOsa0XHhsWnX
EvIEDz+EYQCOx+nBrD58Lk2P0IpOVCEkCfnRVTgEyh11NXzG8l2A11dEaCMKdEla
5i1SRMnJiwp/QgQiawqaekB3eKV2splQU1J4lG86guLDWlVqE6MRbYN9seyOEF0E
CDSj/EdcIVee2kEh+UxlKWGJYFOtCcduvS2dzlW8kqJSeDyT/APF2QpFntB+1PPQ
J9J1GyMSp5fgAWz09mp+uTr421+UblLo5L10bx4PHTPVlZG0Rbm1F9tfnP6oxh0O
xvqbJE7yMeCjBdWi19TXAdA0b1Rn2tvoGytNvCLw2eXuwun8nThJo2LAiJ+kK1Y6
gVDU5CECmjKBJwvx3bvhXzVTlBaxLl7hWybyX/gsbX8fUnPJC9amAQjwS8J3j+KD
el5JEjIncjkts/yV+/+XnwiUkZExgZE2hggPceOKptOeLImlFAFckcPrljv8/PWP
AKQ7l6NqKs384OdLI/YAPJ5yZkXykpdxzbkictp7OfWLi8Aq74OAf2uex2ZG2xaP
eMgh871JhGpk4HHjmLl1cqvKKy23W0jitZgpXkZrbu5gOoH4VwfBKcoU4ZqZ7OAH
0RVA1burftjvRpTYlo4pNXAsJigSUNrH3URNY0KaNK/KXqieVXUvIGOW2RU4MofN
ZhQKXU3nTms+CKAMcxS/LBxssuzHmnSNmwV/liCRb/zGgfw4XVeWljOhmfecI+pi
mq3287N62jjFGnpk8vB5/ntiRP7h4MnZ2aSfkngMT24FgUBBxs9qUaBiqGRxhW+Y
w934H/wP8IOlSYeJhfRNyx/7Hf/xDo3i5xlU2+fPOw9+qUCeZ8CP6FWno4zUAOlh
kj1VoZPNQdPhiaI+qubbeKk1lZZ7F9c56IAQMUQidTB3IiRy6FpoOE0G7Gfh9wvi
016YV3n6B2eLDFDjeCbjyAOo0xIxRgfCUVAMjDrXD/4A16HHa2PB/C18YLAEED3O
gEyqTxMOn20U0FS/bnKqOKi1QjiBQShB7KMjW9j+hjLbEw1vX6dbSn2KzGzfZ8lc
XPiGFfMjBawY9JXF4mMI0iGKWjjT/2ABtZKlLMTlXs610o+OeSRa5TSmAYIhiYok
yI2qSLTqpVohxAPPLtuohALLjWTiKZLo/zYGfgYmXt1SIBfxK7gTkk8N3qFN06Ag
j9QQ4blGy76b3WIEwgLzJA9O/js0maCYIfMIvAGC2Wp2pBXKVkOfG5r+x8akNWjw
rPhDY2uOHwYD5k2CAIpVznnNv6V0kUTUFdrcj7N347pjfKJEaL/4jj6abauAePdO
ghGNAWvCYUMYM7ItIqyPPIMaCvMbmYW/bNdm7lddt7oc3GRoUW1bJX/9XcqeFe+q
3lCWmOmM0caTmD+BBGZPBWbYLIrkSVPG64Y0tvqKMPlfZSWBD4t2HLztgh3Cs7AF
yW7O+JfZjKZhVPWV1vT7GPJKcWyV9GMmMPyDv4oeIX1/UYzu+Z6j/jc/nPWvr3KE
le5FRD4XvkOD7ydGQSXbpePiOdmoppBS8wgF3bL8goEutj/i9hm5gtWuSEu9Ljkt
X5ohZz1IWEraIXCQFZ3e1FbMm6/YstJuPA5ApSJrf1WrKLOuWpVR5NusFG9mjB/s
UVdCyamGnVOF3rXzA0wfnT/Rhb8Jyo8Lu16h+lK+XXUHelOXKRMyuK+dPhDcVYaH
VmVWIQKRxt8lvqfb1ONhy3vJW9q9bPgEnqvcYgYnNOgLbIyE6fMcgmCkXvUXa/Wh
aCRddmgwXn7cc8xCUg5u740iQaTQuzFhKPDDad4ITvaUF5I5drQ8vIW8XIVPId8V
u3+b3d4jbfYz3vJucNu/3aDEzvqzqAfwHphk/9qFZLd45c4Dzk0LIrHu4xGA3XUW
rl+hGyjmMe3aM9YVq2eRr5aT8BaVV8LVj1Lfq7LJk2BCmAPihvjINxQ3nOxH04Jd
Vr9YYeksobQhAc6dlUwIo2prYBmk1OBJwVRqmynWgY51x11eTJgNOcXY3u9CDzp+
8BlOvTrkNj6tER76NZYb38otIVQgS4FY9O79hkateAq/4WYb1dLaVsDvHMQ20RoY
sbaHxvlnue9fNUYEJz8X/XxAgdUEDUSiLPu3APwOwjeLQMbIbgCxADE0Dl4o69hq
OgpHkOKZRagoaB2n58ahATTg0c/qSEMdfrPRm91yUair6u89fTOfxDAgHzXn1OLi
axhbtDe80h+QifqjBXGkGEn8b8b5X2T49UAOoVB0NZTzcQqM6f8KOTOTh1SprX28
XwZdRr9jH+J265GJtzymhODQzXMJ/McMYa0BY1npPfhEn0lNA4IBz8hMVPtJIUw+
IfTpfKmtEEOmvYRdrs6yhADI+jIkFGgF79FXTa1Yy8EUFfgpX1t8Ka4pq8frOuI4
9N38RC+F4xESFyagM5gucqRJpe/FTSwq2UqBqYal5gQ8yFhwjO9Vw0OaSBLGF19k
tvypt/rNZ5L8HRFN+mWd3cic8vL8gKb0QIXRjs68tUTlp7jVKPyFPGlYSbDdkpP7
ITAOFxEV7mT6kxiKm9GMn29xubWZbTN3jnngRpzdjGGGDG7uEFs7Tb14VYhaarPL
/tlO2ttjH8N2JDtLEfGRSdiyFm0aeeZ/dVlAQg8JbPbYyjVjcd41FXRWmx+O/X6q
72LgxCuNbxIklDTLtNc20s1bFDLHFYcj9K3UPIHoj7ut7KaPYoGwmmR5jJLYKMl3
ijADZNVDjc7R7Ym4zU7B5RNUfEVqguz88h+hg+BZruVYp939AUZLMF48AqeH+iPu
nJwIzluF++BLxU3oksiO4LbDx1GWlbbOpeqt9Mt4dX9o0aVKWxxa6RxsgakcLdsk
fol8ec4gIulRBafpicwP3IrlruRHeDijYdzxOCfn7cVxo6mcudbhoLzSBdSfjFAL
RpnA6FsRILshjNTt3WkGC45VwiNFO66C/CyiE6WcSPVV8B2biwVTonkBrLi+JCUr
61ToP8aPbDvJSpKHpxJ6rdpHbu0zZCRDyPkqH1H0Wak6yz04uwgFRSkjruM6gx1W
j2Ml2XYwrqlmtzXEJgTf1e5gVWs5LO5tFKQSZCm2gkpO5mTnoNvTSJEa71zM2QX7
u4Se3U2bTIHhm6rzTG0eTuMl9Ct8TDKgKjRurWVkC5/DhFqqnemWO4H2/Ethh4sl
ayz2bVB7te7l0wtQl8pAMr1OJOsHX1YNT8V5r+wHO7qfb9fPWl/Gc8c2Q0SV7/YE
3ckxst76y0L8nH0VU9NljBwMqSZRNkdts+YD5VZYwJEc+lhOOSXXmePK1Ra9Ly6Y
P7BTIvDJgNDin84KLeu4VYQsGYZj7XQEP22pej5PCAmQawdc6mTIBhpyoq89fEWj
DcRUpW+P+9TN5a3me7AfkBWw7iWAR/SLIfR6l+Y23EJuxIXJsMv2ll96HyaKACMg
QW66MvHmyzClkTKRCHAQyfemY3q2+ygDUg9HrB1DzXGvA7M8WrANpNqY0Z/Ae8P+
yUbafVD8P7m+83LhMRSQU8PzHDYVyOG+S/JKHB4Gaf15lcvgXVcpeBnj7aUgfvWo
yVRs57++/D9LHn8+fhMbrg9gqYs2cbgu0qLpOxpeUVuK23eV6uhtGMopVdfCif+c
xJ21/w9c1VKiC/3uB2l9zPlFNA4HUH9KXhG4mwONQNzUooU4SXWHbeGZ5nkWml4B
HZOrwRu7Yf7O0fTGPYnIG/fnnG832EWcY83f63fldyLHEUt9ZvSwhbY4Pmkn45VT
coButpDe3NELtKnuJOEvyzKYy5s5PDO33ws7pt9NmKwUgmSe5ED0ZTVV9eltD1zR
4bdzmbVJysEFxBC9L5VkaAOHj9hnMTl9w+ICl6nWHGbMcnAyhe9HuQq4Uyy0fAAt
W0/afbvjJI2y4WOLKajsXkMCORcvxCqrq8fPBlTiMjYV0V6MlgXM+NMwz4ya87UY
i2QRzr/+Jh+Cu5MjTvAFdQKGXaUR7SYQbcD21c9riN2pdzRZ52faoR+SM4IDuvWQ
AK2BhtDqQYDlKBoptFvWn9SiX7KpmpXA25c/WtVakaMeZ5Lfiz2xsB/SrxnwkA50
9z6NkYY4RIZxiCHrKu++R8EWTlN63kv/S0KEzECykVM4n9MyVKy39nq+GrtuVvHc
Iiexda+Dx5zm7Vd0AA7SxUEysbY4WQjojYKoO7AEJDLMnBtW9XSngUitTVeth673
LrVsESVOGDWKmrAyK7Vqu1YBelDDUXFJOIaEe1JLBxQmbtw4Txd+7A51FCOVHXDL
YM/emEoJeDJi698RvQ6mlCww/Oi54q+/GLue1o+Oovn4Do0Bkr+X8vlrmAztZboR
SYQ5NULZys4O6w7q7rICIoUQ5QbjVjBuu8PUXCgGImBaXln1YNP4lhL8XVF3HCra
vhNaVrjYiH7WTrkRA3ZIOJpYkYheP13h6rmnrzmgRxSbCLsco9pyvN+yIyBIk75R
WddnBffDY85lcP9VXpiNL3YgCnoT95bT2f5/vL8SO7urrWREzof+3lbiJ8dGQGdg
XZfxVsUVhpxvwf5djiUatwABsoTBuMdRpHlM4UCGX4zfkHzFP+Y8Bd7UaMnHndBZ
QeIoCnQpU7eEj4Dc8woJpxUChohuk2+G2Q+aX0Xjpg98hEpni/YPW2YA/KUKLumP
YIC3Lqf+3BZchFMYSIIxdnR3y9LvJKm94OjrkUqFne3xhlCACwdIgiE7X5sPtClq
WvCTav0ZRKs75NgO0vJB8IDGVpuK0tbTmNICON2xASbL1NmyRce/2754PQrNVvaJ
OmmzpPyv9DtdsgarOybCfTgz7SGRBuomSYrJQvYBZTAh1whf8yrH+qcUhAA30D8D
5SbDdWCdRxHAHnMOgmP1YmwHiblVQf1DCgatW7hvDRDGaq/lX5YK9gCyaiI7qnlr
D8qkb4YvDRhWhp/v5whKc4R5biVtCgqPCqrjI5hNrd7m4WjRc60Rw7d+s8uG/kyz
leGq5hsgYjH4yW6J630Wr0ftv68gk8awMZhC+b7gOjeQH9ooJvIejVsleEtGXD2C
nZEh87HW1EMVXeIKNBZakCw1Z5eEuO43UtmivksduY9ZkAxKDuiks+skX8A7YChD
2P7pZAnagG0oPo9Ogg+oniw98Zpro7Nkr+ubP/K+Wdx4WThtDrmy2/in0CAm3nrx
c1HISlzUiRVEyXLX39eCIuGDccWJ/QU+wQQFLZdaHohcntFCF4TOkUBTKQw7jhba
dSJat+UJxsXYy6rwWABtC2L9mDspcDMFlzp2nFsVSpMKT2Zf8PbDB0EZrn1WFzOK
rVSmJCQqRASYgX3slXVKqwn1D2JOCKBUhetgJnjb4vqthcGibYWhq4QfQMKM4XEb
Wsqvp8lwD4CptzRiDZzabQ3w9IlxQEq5YKZBhh5Xuh6NMgr4nA9NZWp+XhYIwZA7
IUn+JDMd8wYnUcgNmsGt5fbWYAQmRq3PSprMwMaaRaWE2dOVVmjEZMeE5+pRHwzP
bR19Gx3IcU2a6pFkaWK1KfkNL+q8UZhE1JZLf8kP9uCcoqOGz3goqs5A84ze6Mqd
Hf/h9fkc0sxgkmohoj/M9D5Yc5rINHDyuCDc68RumZRk4t4gEZA2xkB1KMVJSRz2
dsAKiN/7FqdYvsJUIl29sytS3x6mjC+TV6NjEQl5ii21/wC0ZMakjOMoePhZ+gQl
AmzuqGpc8c97NEVEfDkoUGamwDyXFp3A2hpJTe1LGBFDlEeXgDdg9BA7oBPvHq2X
+G4OkfepWuvVmDM1ZfpAPnuGm/Hch9OyOklyEFpM3dj6acYAsI/YROj0gXbpdqUA
p0G3bSPBTpaZa57+K2ql2M2ywQ1gfViarm/ogBKHvWpXDmldIJLFAymjzxBgvrIX
6OPzSr55R2lM28WzU67gjxT8wvDVaCj9jz2Y67llA13ooLmmU9PpZlljqKZa6/yl
H4pXLpfefOqdew5N01lE0xH+hsppj/ABiErBRghkijwslSF2/r7yaat39XTs/K3/
fWZ/vyUikbycj5N9sn8FwE8f/TXAEVYBBNfSalCETVzaWQmQ8lUUD/VxRQh20W7c
U2XteLBiqiJC9SVtQBEPJ/uPdU1ditwEmG1JwXZ/nqo8v+wsvQ+mLTOS22Q5DTx1
BQJQpsaTei9O45vyQBxgo6XOOeDLxrjQgqxvhZXzBwv6BOGsa+bt4RrjVHaeQeIU
K4iBoPyHcP5RxhvQtRypHV9AnpzTbDtKPVwnTLyf6Ckia+ofrark98ruz93kBPLa
+iplvrJtFnwXNG0PETJVjUY/CJVsGIp/FILu5EH+Z1OSroo8NCFdelDFoZSqRdNa
cd+vRsWHkbfDuDtImCbTNPsILuUx0cd8d4/eaEHzh6UwEnF1kzoJQRmMPgdGqa+W
iVNocR0eLztEhLPnKL1Cu+2KUcEyi75uZOi3ERbkbK1AhS0zqkjxjzOl//woLeEF
38/vdBJpzChXt1pQLvikm/8gfXqiKlArcY07p0D7vdju/wQcQXfMbeMQw1N/OBz3
asbaQFp080dVWCGEb2ExXd6+xwe+svphkIwqsFSANyrU5TxvtCfR+Ak5D4it1GGm
oCEqqaBh9y80758lGeq5N3JqfOS9pifnwHh+WhRZJjga+mVJO3P6LuBMNZZNSjV7
7tgYR1qNNxkKrJAaMabpoUCV+gPCb/1gRCYsrgPEF3yXQdt+SH8xWi/8d6RvlD/C
0JQKRNN7/Z3ej1SNwtVAu7koIL9FdrE/pdZtNI4dcYCHnpTRAQdzUOoAMfaRFlaJ
n0WaJAWfc0R/g59D3Tz9yc4aGMaJyw0GV5Z7lL7CoUd9dvY3k/1UHNo6YcmiO9tw
LkofeKDIqw516oT3Yh+CR4kmv0xFB5WgwK3i8PJqXIvqeJuPjNZ4dWGAgHh1XgVQ
Rvz1Q7+Ue1SiCsCPNtPN/WhsJm7jAdMv2s43RVbMnQAl3gE8KIMclM2OxVcuZBYU
yrm1fV04dgzr8LDsxsRKnXzUdDUftN7OT73Ubg1wZ7MGBn0aQjaWDVFxd6/j1z5Q
OxFYMhfcoK0E66PMz6We99EXUAC6Os45I0Sct+WKZj4GHKDbrd5AINUk3X0fJc1U
Ykj+NZ0de4rt3cn+wzvj0hz1CMSdxUWUuUqzgumVqHDL3Uc093uC45lG3jBJoACp
t6D+uWtGtBTcNblfiOuvJkzAuCiknFjaa0YNtZM3AigtbkjPwTg0fTXDXq4pw8/o
46tSi9UK3t7R6NbbJNJQs4rkBPWEApWwrRzzear6QkhDwPnTOeLAEDcAhONWBlph
3b+nOeyGEH6tAKmFWbU0ypXxqiqKSeRaiDJUe9LBTHquAmO6R1Yn7dtBqNd+3VqQ
5yloYqwUoEPTCgprkfdOwJCTNUcyVzesr5NjPkdej5q4HB6MTuVxsvJh+aBmtNEa
od6ji6EFRBwSVC1IOpXY/2EbFKUXu7Y/syjgyj3Yfp7LR+Q6HMePUMgJ+w2pnlSY
7p3baMv0WsQBJHnaoU+EwqYDNM7uWREs9p1iBoW+c5xCFJu01FkPcwgtDbNb8FCr
CIURDE+CoKv+stfvxdGZJ5mEFWNhXU2zQ9qfOc7PF09HtgVFy5SBCUvZxSGoWMQN
CpRsFRnF0NR87DuM1GtOhnUkK6YBkDCdEUyVxB4wqredoptgffMA8ZZpoYIGCQpO
Lz8NLnXPKGkxHZKUi74tujmc0F7a7npIxD/TxYdpHHtr5b+UL99Zbx+1vhjVjjgp
4hv7jR+k4PVTpriCKU05Ap5I3tJtV8KpneCsyIHfRc1BnS4bK+alSZJMbI6Zh1q9
w9LCOhxaeupVB5h1uJcNrefTyf4zzDp1t3tZhGjPjuiuTOoB6WKsN6iN97t1bnC0
1DbkmI2ClyCaRM1hl3RTPgz9qkz2kPn+C2Kr12WOS9sYMgIMZ1cpVAItqzEB/6cw
tcOOzFLlaOQ939k9hcQ2fbGFxg16GMeXs4a65UZuILN60MIgnsQ2VWftKAuCl7Ms
ksfx7BMBqjS3OsMWIJXtdeXRZx/I6lcg8wR2pvdc0p239iVNcjrpcSn24iR/7z3Q
vyIXq55Pskcb6tOGfQv83np9nKq56ERJRkOtmffAlSDk4pQ4n7pRfgU95UY0F+sC
Bz7jANPpZlA3MeufXT+wdchcbFd9B1/0qnL801aYFJyG8WdUbP5MMQASnm/RjMP8
12vWxY85h8f+ubu4udZvjnrDbV6ZBKO8aNNg07VPL2vqCEhBzpS3u/REH9w8mTW9
Y/yRnAYMwBZccfxURyGQbQmTzfYA29KLrspsq5lNXoY0bmyE5Ndf73AboEnyGah7
oe/IzLm4TCzrJjnbTKD62RIMR/lqRIWybdyze6Uf5T71rY7VLa2FeyG3KAQn/Bse
wnVDOzB7n15S38HK5Zvjh+V/Jp7KdCM+xko8qLa6GqNucsylV+TysjmTIcfZDnSY
fFaE3rDibZBMw1iXjfxAtFVJ50HGX6EPHp7F+46y3iUZzZePq3fE1dy4stJ6Zbi3
Kn9dvDDeklfi3BCtmhUxyuAx12kYU9s5DfAszmDFIq/fjSFWbAp71KKZOVc+2h2e
tQZnI5G1Q3AdcQrPc/fyNt73Iy9BSHB7Q5Bkm1tIhkpqa+Labk/mqIHK6S16RKxh
/UWVqunTFtWizXgW4ue4UwiIGVIiBi0PhwE/eP5YnG/btPOQvrYGmBFBWC6h0VWL
fcjY7wbMUuOiljS/FczncsLqEixsNFpIZXtXUtyZmeTQ2qdfpM7J1m2k7g8HGoQT
c6zadm62VF3jwu4olGuBxwvDMeFOFSs0Mn/8TcNtwsdEZJheHs+aIF3dIT/hMEc1
6K/vHnVnkSkHUl9rbwlh57SIlj8wNlk/0hl5R1RzJmNq7BncwETa2GYD0ZHtv6XB
GysoV1I/QHscTcMXfXlhn5RLeE7bQsTkFpEY+rEEQWE1DLGu1/NQkeyTP+lvrhv/
gZtvkHNEB3sFPoVH5XRia0fYGsf6uEnqv/tmeVZcYvzVEcj2At6XRqniOPV0qETR
LHNIBFKfFX+u6vEIsK5Th3761wLzen7hjoXsQnr1Mt8pC6YnXamM3R3b6o52YVjg
c85jRe3AfNAuJ0RvnC2L9yvYq+PDlV8SWpnka+aw/o5lIp6rHgUCBchgRX9G2qd5
vw+3EUqoIkbQR/wRg5P/AFL1w1UlVHtSH+metDUFfpAt46zoENf22a4P2Croj4Gc
sT9bB/Qed9zYPG77pETtB3rCl1LvRjfwT5Sjm49rpZJdYvmr10p24V3MNRauvguE
RylSY9tFYE1HTIDRxpu6O6wVGIxmKHt42pPK2vBM8yTWLdZraL8k/NX+nUnjfqyj
rCOzHKa/1+go9g21J6v1ATQmHmW+S8qP0y6kaY51jfTuJ5VdsQkedNWi4qf9DhHY
d7hk2hNybKrKFoT5XhYul5if/a15l4/0NVWdv6tSq0WeIez1LPRgZht8wKE+7z2+
k693oP4k5ldS6FbdyTi3YharKigPulCDoEeq9IL5UEg7A9tINyMxgBYWQCxK9w/t
rUZXzYGQ4h2k5uHUrAc39xEiwqXWH/2Dk6KnJk96QywrKPkbYiU0e3y51JyKFPR+
RguKSncqW2XZ9iB+1QKCF5yp6Z3U3D9wlktbxKk5KROrfR4iV5F5LZXy4AI9/lnE
QYeWsLALBYY8cE9bk6FsvmlM7a6+BPwPSc24E0WDUWO9k3nmskPZ5kdhj59dXB6X
IAJ73CtDGSkxuAYnVKfLZRiqoyUPNTmD5itrC6HKiRr8wlFob2RCl8kKAKwh7aPn
cd78WN8BYxtD4Rw48N+0XGCgN4ERmtq7hQlCn4EgazWZ4i8eMGLaDkR7mTUC0WiD
wrW0ZLNQq65UtDmpduropd4pApv44ZpZ16Ie2K9sDsPv8LKRgWoKaX3llocNTILj
eohYTTw+0SCZ35khcSJu5/jjncqWV8JL2rNlZjXEgtfcFZXCIUKr8syV6O3uFaPU
Yt4zhkqH95KsXmPCJOIRGwngQ7dI3Z51c/uN+gkXSenrmFfdGouGVlcDSEGscOfC
1f5bf7wNaczVA3pR0WJYmFESAQUXum7F3pJ1oMtThgsBv8HHpyWttI+AYSLRGxU0
m9MeiBZ4mxJDP87NuDBQpkypxUEqU+rTSnnPqY8TYmuybCOYNgkE3Faqpr/p47FO
yzqN2XMaSuDk0A08iRY7sJStWBp7bM5Jy0cFB2sttUiNJOdkQN2jFOkT97vo5olf
PcrRuuscRgPwfw2L9O3WW0DFMFn0NZQ6Iw/O7BjfxuyWebZCxqqc5duaJ7zz3fwC
Vd+umPYnQVbi9FOsSvzt5G24dGFgK/ZonpblmcQwv+gXCejpZ7FOUc7ZyV4TjIr0
HzJQ2OmsyhJGD1sm0lfXE3P91nbYahlQA15vhJ/ApDRH49RhclcH8FT5HBULmQJS
6jMlep/ePzk4nqkeWeMo7xiGyuAAo3Tru/Xyb964skPrbQzJI4Tsn9Z+oQWAuWv3
a+xHu73J639HuG+8DVJ6ClrkeNOJ5ZaRdYk8fYlNdTUyOSWEdElwS7UK4psLkpG9
XvDVAp1oTWo3Ic11VuqGGKucQYRvWTJX7UF4yJuGKWT1xK+E1qk/Bac0l4+tRTZW
uGM19zjAEPfvo+qJnkBKsYK/Wj87d+AM7X7Iy+EWtCVX93A95fuXmbKcuEqaf1K+
nbCHjf8lSL5KGDi0T8qqP9lNxievrIxLeLcscNXPSHM6ld/pqIro5H121yHsuf5P
UWyB2/EGMJdCfBj4kY7TujmNcsGhPq3YUgxpMOHc+fjj9VipfdKldVGgcpuQAqQC
2bL6fsvA70WZR8nu9Rb+0X8ko7iDDjujZeP4O5fkysxpNeegebJ6DNykUhY/DC1D
mY6fk3dmgl4XpjLXTbJNcEuJRBpbUYmzycK/DQRPloPpi+GYDSnOF5PRm5KKfyph
hBTMRtIjII14zLfwuFxnDfoK82nfBFGrK09NVZ1lhsyRwNzf0oIrFdLhba2ZjmR5
WCVv7ETkkj/M9KmaXTL4ta4EC7Ootc4wAO+Y7i9x0yb9CittapjsXn4ZWNV7zFep
PTNmsAp91VzSM4ZHCr0+/4KrKf0PAJkQMta2Z/8dQvD2fDfYltgTyJmzhgU+nT5O
9dRus9I/Go++eZOlcROVVsD253TfIr/pkPcrWZICBphE5ZDys1U+rXVvUkfCg/XF
nHIdRn5Xk1L/9XnPj3zDMkcF5JUQj3dOtiRBQ3DlmUReDOwhUdwnh0gvdcmaYnGV
KE+w3/h2bSa9IsdQ+ty2qs++99jzxIs5dL6xdcAhqdtnkCmkbjO2FK7VAnzlZvkn
0wbfaw0yQMwwGcfEmoQW3eCSPzlmrI19PDORAQI70Xk8lJidG5NGHL7bMUroK/Zw
v2e76uTL3Jjcj6tiOg5Grd9JJ//mMWbLvCZfQnGTffkAyLDZGT7DVzVFl4CXrzDx
Acyy5ZoRJ6hefmZDA0JZuZ1MLZdqPq2sQMSqHEUKRPeYB9MJW7W/5uVmwPMRPL8j
zvl3HlFkGaSPLRYhwz3udZkDnfRbav+K94alNlGMuP1NO1zY+gSu/8UxffP25G+b
4JI+tRS4sC8fIqlnAK3FGztrs4NT6robL+P7z5kB7f5mrfyOzpb24v2wL8dDYqZU
51EacTTosLvMeAPLK9/kUA/2N9ErKivi8Bxe+q98XVHNl8bpf5nGwYSnWQ92hqNW
4XpE+v+4XhsMtILjM/YmTAh/XMHAA74pnJtjYNPob6Ebq++V9lwHLK2vTLv4ufhk
s7QNYSHBD7rDD42p29Vk7/gqOLPfieLWquOlYpkco7XomqmnRSh3PEp+t4F4bEZA
oKG74HNDqD+QwxdloWTRaNm82VkAPeqUhTaSbVI/56ePRryQqHVLodGVS42tIBv7
jAVJAh1CS28y97nVQ6l/b9pETn3PQGt0EptNu4aIZ5PzL2aUe1iMsTdIZ8SO/pxY
FO2QkBXFcERF0/BOJ6HMjbyMpm9+eVqEBfvxRetb4+h9tQaj3/B5gqgBsE8lrcrK
5u6tCz9iHVSc2EsxWZqp9AG6YQe3IOEDlLkbTzfWKkQrp1nj0wT/5bCYXmjkI5Up
Qb1WiBfwrHviCSFFxLVZxnFm12tJxoF07OCL88ViU3HLwHxeToVG8QgPgAbsNgkw
GtT+HkVMbv2i9NLlvp08PDpn0nEuWjguSY92wmoN3dD/WsFm4FJ4HyYbc9hd0lBw
gWjg0ks6eXiaUNujP6UOspVcUb6h+wA6SzBSb1fcRhkz1pY6ntxEuacscFeKly82
cayIGxWVAsA1y0UWmvRHXeYqyAsuybs8Co3qxFovTe/GEoeB7FbON2r7hY8N67zn
Is5qOz2N3rBiPseK3G1pu1qVObwmJrEoqC2XNRYhWs1w5Ng77rHTXpQVhFyR9dyQ
UsCE9WgteddL8awJm20EME3pBHDdwK3xQNH8lOoTXYkrgqdJUZO93teeaFSPXqbf
o4+/9AJNMZtu3QXBw0zcyYcBbsZrCtQh9rmT4Z7z1HCvlLAM9mNZwvJWykHeZszo
U45I+HLZPxuZ+blSac8k8Kr3zcb/bDIa5vlTWHaKn6lh3qbd2+YiWit5H4xev10P
rdJ7ZoN+slCHi1IklBYWwsWAycWy5aIOcG8DH8tKNBb7ePd+B27OyickKQVfKv3V
TkmrZSUm7hG1KB6HlcMsozOiw/cIWooHa4r8M49Y1RhWS3BqsuCplul92Ud3Tzrc
WAguBRWyUgUKgS6R1fRJrcLuw9cdIQ11yfSxBC2J+zK6/f126tRzG5HFfPZG9vJy
QKWBdEeKq0uDxHhXzciiDSF9+sxtCiCh2lRAlef/aECHbje3fTbQQ2tg0JK0+7e8
1ml10svj1Led6ks8MRsGut+iQOp5LLoddp8KuI/aAocNmRxMiAvCHkjkcvEoYByv
m64mvG7eqi3hcUC3pPFC4HV2WAjaLu1Fn5Gc6uKaBX9Nj0UNgfqAsfyB3Qctid2n
p8H9E5ysWATcsoqRWC3JqqnMwncUKvIRLcR0HHCmMqIE86pwuuD1DkGkVi2CT9ne
IM2Galp2q68z7xwVR8WLY/hhNWhTH+ArYX1xg8geS+ysWHY5LSlNRRk4pTVjaENp
HNaTevnsrAmDfKcoxvZyefXKTbsSi+DR3uHeuPl667m3wCDHOSYK2FPC/mcVkB/q
MgTGrJlINkHtpKHltYr/wVjK+LqdAs0X5jy5WY4Nsz1wwVJvVPGnTI2c7QCatgQi
qZzt7GsD3DYzCBAdi31dV3tSabLoU5ADFFtSurgtbownSG+Q92ObW9Dr6sCElV6n
lavTBk74xOeRgZRH+kaFZiaMtSrdFNvUSfTHi+1oYgW2qAl+K3hEIbUzLlSnx0BT
KWKK2wytSEOjYpF7/oTx/bzqFPJxrpx2sWqk/QZn1ib39Q5EwvcapglYtwFlEx0m
+0hl8NBX9fGTs6pWRgOCTxuMySmqI4uEBw0HcZux1PxN0x/n7ohu7G7cPtRw3BGn
bNScml5Nkhproxr4VZroNSHwjInNg+odIdjC0im11PQip7ixU0J6f/A6UiZbGu5r
unB+2VzA1r8Dltn4EGp4TuCZ8p0A7TSEn6AhYakYWkykAEl3eEdePgE1DOMIGUVb
DJzWQSiVHFOAml92usIVDyYF8LgNdR2LQqYmVb82XOJ+GewVAV1J3nyNtm/eaNfh
kEyohP9OFuuD+mY/Z9lkXbAkRE+VTEFsmZ5QmQKjMgguzHtSD8eTWreFsWjvu98K
tRyNcxxWAqpaxdDh4lnitwPteXH+KsAS7QIi0s7IuUG8uN0tqpK2iZ7AcwBaiqau
aXYAfV11xtCxYt36W5ekZj/ZbTlbAzxFTjKnu6IKrc1IfmkkdxiK9UC+iaPNxVmC
uPD1NYB68GwLEhjPrAZ1mSN1Vd+f1rw2+ekKS+dulid/Af3ylDLMbOMhRfk6ug3Y
9Alb5uY2Ui5/OJLwQaWKTIl2ZRaHCEA4KROB8GsLbXthn5Eiq8Xv6xUx/oGqAnEs
lgNusEieuPorNZwJVmsYGIQ5TrZnZP24zHwGWH8cUHpRMBUVpfhvg8dLF7+ZG1J+
fZWbWM6YuP24zjGCt6vKnYF4f8cdBu+uGr+GC/1gv6+KmdENdx5LbR9Cuz4tHfwY
ScmqIrFyDUw2nC4u8euiUoRCruAEhFy0sy1A5Tj63xvCOcxUXEHV+oGC+DfmXa8V
bR+iLCDrLdseoww7DDue2dI8Y6Ef4U2pRcYMhTLpDAUqNPT3BvpLdc3BjiiAFvoA
F20lgpunjZWJGyGKoiXz2ia5rH5/pSk7EBrQQBW7oBvQUNDfya8KZIurJZwbh/3y
O+eHDyMahCEtE/NuojwdDwUnZR0YnkFGWG6VohKgqITcLRrXB3YSPzN+ErU/cbvr
DHJGyN7aoXPsn5tb2lcaCuew0DQKz914cX18h7XnyQWmCvDmZ3lVJvgCxveJeFkt
CR1j/S8KFRwGrSb5+nKR+73bt6dn7kSLdQu63Z3bfCRZPnelu276Wkt7rMGM9i6y
z8YQHpXNUjQ2SqPMcVkSRryEAdLai2oYoCwvlSBFdLItNp3LfaHudHs+PPPMsQ6m
tjhHFIaURNQ+OH/CC372prac9Wonicd9QqTJ5NwzNcXlCjKiiUaCR44kojDu+EmN
4+w2yqH2zmMEYv2onwakiRhm8c786VXqq0PY2Z5CwikrpX4IFfjKXUYHgkO5ef0o
zmdfnte3hdN4lwS430Fg03FjLswffjkTddkUfp/T+UbPu1gAo+GXloTo5I4HdV/K
DQPATH1W9MePDskFeRba50cUak+WH3/nVSIETOB9nSHjDnZZXIT6yvkypH4kCC2d
u1R5z5SCimp+cMyWa1vi+xqjzvbeu9resZhDL6rTE9pVULTQaeDG5IktWjhP4x3m
PF9VFJWaPWGMl7acm37Tk1imxrU/D7svn8/sPysRTIsahFJnjhNFjZeOXd4Q3f7k
j2OVrIXxgZSnmO1hW2AVPpBxkBceOWQyrM3WDWGzeW67T5CLnKbfEH7f+pZJxb4J
7NGvcrhUWzjfIplIwCDvaqcf72mAj9z6GIvJi2oAm7cLHiMSqk6/VY8sv3edcK1I
EmdXe08TIHo4Cj5HURkDeMyk26TbPWZfXwRp0pw8LjVlYVTftzSVc5W3U3W0PaZ/
EGRRbbQh9Zbg4xexJoPV5OWs8iiT8w3l8KLXC/otqbNqKuKGJHF+8+DFmkc7PFiF
wWuLu5LQyPXLIzmbpwmnpVSV9di5qUvOTnxazCbdEGgcIlZiUDJd8i4oBE3KQH+K
Lz9lqY2goGqGsYfmVg/VylIs0SYIf6BqFIqMUKEmgpFqWBrx+5p6C/ZxdDmt6jVo
ltFiubrn/BVg1FgAdyN+8KS5oPAmzt5Ni1wCJUEy2hznGuT3mX8CWZqJ2caXuK3+
uvkT8XrHLq6LU/+iOtgXzg0271V2utr1MiQSPlInue4pCT+6Pd712+fbs9b3o/aM
O+wXnIjfwykkoMZpo9fOj3LHtIiIfw0PU0JLqcIaItzlJt9ZOMGyARkneo6lQUud
KkQP5Vm3J73obmy5N4yhNILIOw3fklk+YIgqYgkvHCFG2gNlSDxANLHgHzEbZ1V+
Z+BanWCH0Khs9Cc6hRzaC9OesT4HjRRxum2i1/T6OqgtaCOa5iZoN2xTihtMl+Eu
EOFpNi9d2q04OF6u6YnmsMvAXTOk4TPiibX7MoNxUG0v5LGhuGkXSwnK373On1Ox
TPYLEiChgqkJDVuCtE29xMQqXS4JvSlwvORIKV/34x37HhAEB9wJC5G6c/wJfwwW
yYdzHrqRAWDFQ1nFOA9VwyNxRBgzymnRLg5DY8XTK4MOHWgWdXjZBe47Ua4dB8Ax
NW63NSQpi6DxDTbVeIVpdm5OnVYtK6L89WPMnWS3r2MXv8SE2JTZH2ibOYX/00Kw
DkvbWvV/xCd+JFtQTEgaDQ1+hqFYXVaNcJdZR1UpPI9aSlZeNCThhEGZelt7x9rh
0X1fec2dvAI5uCWOtvVTYuXsEAeYx20BjpV6aEFHuQqiuJBbZwSkAZ8yv7yy6GV8
Rv5hgC/L/gnYiA2wue6vqWuqREaGkYrtoMKdCeCK/7Zx1PPQzeeZ/mrKCGp01sOg
Tlkp0+P/W2nXNSGfcpuv719qTXbsXGxLSyED/GW6KM+S6dpF+Kpys2LNaT4YgfGX
1MoRQCgxMpQcNsMJgr8+1AMJ8HprUJImxcJMRt0M6aR74t0jSzAu7HqNCFTYcJlM
4OTqvaQFRTvbHdCDgV9zCyGSwLUZ51w4WZBy+A/Z61fSdv2G0aRN5cQA0JvnP2qR
IGRUwvcFalasZUF553QUrcu2efRHID4RPdCHeBHVpoHOVKhp65h5LtqwSGGruIuN
PlFi6Ui7FwvYY+uB0gjVNo6hA62m5fFvkOOMSlfDzgObDVa1nz3Rp2UnelftmMFI
A/F8J9ZiqMbZgoqESnE/Z5zE8ahjkpxVoVd0OVQ0/USYWiHOQ6kIwzpZDIlm65Fh
AAs8TR1ScovNaDsxNhJXUXWWBvEHfvRXkTMT43fjK1EVpud5XkvJlYkLW/ituEKK
G4I8a0RC1s7uEH0sk9VeUl/1oD8/vNXvavxaksbcuJ+b5JpI6V+Wm8xHZN0SuzfZ
8qev7R1Wd/W8TNuT/6OVmyjclRTc4EbBUF8uZoTESu3K4KrcjM2J7FpaopW/a+MY
/CY+6/ehNjaHVKmFUJ3NVlNAkpXVrXEgJEPmVvNglTkAGL3Y39K9pJ2yRE7+3BdV
OcvlLqIQKocl39oSDFx0+WR9rkBhUzC3EaAUDGPYP/5fl2Qb1499D05V2QsnssQF
HJAFzaR1Vbx4bCICn6AiotMoVWqftDhR7TL1ShKCKo5/4HyCmz8PA3OemXfNs5pb
/S2Qyqowm7P1wIoQT8HCSw/rDS7Soz6+sMH4Yrdf24dIanz4ek7Wy/wUsmRD8T8S
nqyr4JbPr6vFAHGh9rn6yav4j4r3sJzmg3wzBSfdFONVUzE3JfgMsRVNwO9cIjy9
O0/KgEnEaA8nLYE1pYo5WzbrdkQNyRdcG8/BTHjU0EyFd8u1Ko9hjrOf9V3GxLhv
7l/OJ3Tvq9ynYAbwvRvvnMw6OZto6sCEpG7afULQBFOYuElXtyJOTNllCirctNqB
Taw4jrG1YaAi3uNS9tEk0aoDTUoM1U+WksPxeRMGcVQByuT/Hv3EePDMZPZ/p4AL
m1ofpLQhhfReB0tlXmQzlOXtAW1L2C6RJkcBefP/LULwiydBqBxgJMK0cFvQuIf0
cZg6pCqjpk60jcir6XSHJiYgkELGtmCDPWSmg6kCz6S++57sr5YvG8i5Nt0HlI6m
4gX20HDSyFST2K3BLpO9fRB29qeVp8G8ULwpgrN5V4G5rD8MA/tIAyQ6xvHyATQw
ADoKMo7kXCl1gLQbf4DDmHCXd7MzPK/+tX+AejIWN4xoeIZzOeFywMuuCTLRLHqr
M2j07vu0bmUAqcm81PwnboY2Iz3qP3YTQ92PeTx9820h0ghm5RvdjsdMnD/x+fVk
SfEfT7rlwHih5NJxSKrRcADVE3W2Tf22FSHrw+KPHPzJH/ziYNzHtRrY1d5VkqgH
otGsiGhP3kbLfpAOsa7HF2u8XDv8TXodOlbNT2irIA9m/twoRqsC5DH0kXRaPjs7
RSSKHgpMaWMjbby1y5I7l67PGcmzky6Pi1pElt2iVwLOx1Hw0sq2a+3AceNB+Pp/
yUExJmUKsgWmgqwp7LeLYnwauLRs0NvrnAUMT6+VOnh5R5WcRYLAEc/L0RUAchA9
oDGJXjUqxbRfdqJXHsatPo3PjsiC0wHAYYlTU7KRPkl3Q78iWrGyMyqFREmCCo33
0mcxTsr1xCPe0eyiyG9xRJaBni2zySwP6I3F+xyKmd0JfpjZNI3RyDqDULAxFzmh
X+wx7DUOlJsSHl9xMTMvIpLjonbX/Os/kcGaJ7CX5fLfGatvwpn6nqwJi8BzkbIr
vCaBoozFG87OfbS9IsKXfIRWKsgFTCZ4HBlXXSHAjQvsLMqAihAMbkn+7X6MenWW
eqMqakSLEsNQUY59kU5XiVCADK5H7LAU6jXils3iGp9hvz+FCHGJCHx37YOYmCBZ
XViemaaMQKuVl17AB00zlG3e+F38Dv/8iWImDNZqMKsn9P2PW/oKsYgh/gKgSN0E
/Uz0ruea+LZQ9HXX7uFY4/N29fBy96YhyPIv6PBfQoDT0/Kxfh4L51+YwuZJ3+Da
L83IDRWM6yNwPEXqmOuQi5n4Kj9pFi4sVzm15ONTwPmkHsQuDyuLGPVeFmFEip8K
gERQ/02hieZ2Ri+qiIVST28Eyx3HFkb2rLZinScQTRPCl8v0MK5G6DmQIePOVWhP
yXa9xO5fjjkPxKqRtl/zWZsN/951UqTkklkNXMDrCFygB4+NgyrkBhwF0VKB6Qxt
SSjeFvFrWtKsf6R6xFjLu78k3MR5nBw2qbq8ZSGC/BtgJ1HXnOjlIkn/tleZkasj
9ReXmp8T7eFJEbKZghnSFzZM3l279U4tp0git1Lmr+lfehXIEGN8XJyid2yJ0C42
sfTtoUD7SYRJrHms7mAbt19Aky7wg8+SMUwNdnALpPwC8vBxECodYcXOfxuW8Wh+
aE1T1RxuNaSh7O67+PBzQqJLWcOuHMcaxwmQ0UxLFbhMOPkCM+GFmJw9DEELFlqq
jsiB4ukdtlxWPUgbG5P75qBada9a2kMEEP5EB5E3uVZsYcAvaIib2a6c1ELVl4gd
HFNem18tVo5wEN34fIRWhydv/3PbTTdr6AvE9RYSWJfyG+9XnF8AmiyQvY9nPqlx
FEkpjDEdAzTNQGNy73SfMq+bbj+RN/uMN/lxDoVS5zmX2gYmEBSrOBQWSG9nT0Te
Smqmbe8/9d+ugDHPM1XMHB2RwH00c3sY4d50baKF0xNDWNF9rq4waZ3nc6TVNrly
ydGx7RAJ7wSdkXsqo/y3zMg04hanlSPSKwz84EVX2C+IWVLT6OJW6itrSboROVmT
4f4Zbb/JBerBGumxO4Amyr7IauOPFsaSwA/ABq09PyUdr1jsVMWNslSuFqiPZCmT
vl4GCdDdCdq0T+nKabYKKef75mEA5LagvNhlTARcf7hy96kGdgOXyZC4PttubFTB
v6e+9b49XYr0v3KYhCyDKkk2uVP8cqEPWCJAOtcBZ9T1tT0uI5Z5KrW+Yax6D+49
EKNE7gpAzm02NhFbZ9FV8JnY29kBe+CBO5t4TJSadFYsqyxGddLu2R7WZki2LnRE
iPY2MMKXzMM2qS1KEA2ccSaowP/775LLJHkyEkd0lZZmGTZQreNUZJX8UYk+o6HQ
xmpNuS6zSBnLYyWjd0vayZMaGGIPUy77ABCcRyF+bqj20ty2j+IxeX3wWVoTY3X2
SkibhsKkqxYjAJ1lw6u+i9L3nU+aeCMO0gU3bG5Pg80RGxU11lEBbPrXxzUHZqNB
vcXYYnXLHLoWEh8vwJwDvAaytZqxQpzRXj7LdEP83VBbufYMR6SbJMDyGIxu8R/a
asCS31XZtqCqXB3dp07zSeI6yvjQglGBF6ibwAmXwaSrI7okGiWBX7KckGqVqjKQ
COZNDgZzLG6XTxrpI9jkUE7Ltl7G5bJriOYx8ILhsndkRpeOG4D3foqSLtk6m1Kr
KNUeSlNhTB4RGq+BsutqgRuG1WwbFrjGdaE/yfZJti+OCXEvxjTNtZNaCE8s9Z53
Lv0gQm9V2OtfyjjMvq/Bm2l698rCQcR3fQtMntD5w+WTZayG/UnDkEELxyrcWfcz
TGLJmFzInQKP62BeGTEvZxorgilML/UebnV7JdFwL+CW1mMuSnY5Ja8+ElKLAMjY
hpi5URTzKN3gAmEMgPTKfOze5KBlMqWuBBWIk1nCsQ9AwoYZxNZb5xCYGBFKn2DC
GHS8EOyO9KRNEWKx77KKFlnSrc/TRzrx8h2aHIZyrBhj+o+dd/skjf3rqX/xParl
LLsPe6iR/IO/1MrQnK98wvxOWdVAO7mHifgF6LOOsUsij4M+e5BKBtMbzeyuFN2m
1JFuHtYIbCcnnuHZUNJ/iHFAj8OjNdPuUbuB+lEWUMDgsHd7+JgdkswWd+V8vNpZ
835l9BF8BTOMdAUU6fNAixM4+LZPJZub0jclxKyKCxKGGlAJSSw1PKqm6qA8mA4Z
hphDRpYxSitB3r6923qrW5mDOnOUjARhf9hCXVrNIjGYXuWvLyB87tITkVNOUzfV
7SAAozleg9p62zlQ7u8R9B/DS3NeESCPxkrgQsGI9Rh7tmfmTB5ckl46g6T9EHcm
s4fLv266PZaKkHJGNSIxgoMyN+e9cJBo0KrrWAUr2DbrpoQVq/SoTSLn0zHxqyU5
VyRhd6N9rKzdlzyOEpeprU7NDcZx0qoVQ9mhbEjrj9bsuT0juRVmU7N5HDJex1C4
LD0ZBl1n2yF5IKmljhfKgqex0NTG8NYNqHSzxWgUkONBen5aDgP3WmU0pzc63ZQa
B4dEQXPVc5sE+I+UiZ3H/iewLlT8DasBYdK9SCh6uOCUmUi2yVFza/m1Dr81Mclj
vPOyRnj86A9s5Kq8GueLuyb9tM4nRk7mqSgJBx3GHOc18EFlkUOLajuBAvZL+qej
ohKkYjX+xV6hJaR9wfz2pKp+z6flAUD3YOdGOhLneqY7Is7bk8dXvVuIH2Ua39U8
2VgiaSyPZO9MNEyhmRrOcb548jsoglmFrcugekJeTuNV5OEHbtoMDeu92MQfqG8o
nf3/6Kd/nXTY0zGMJyTxaLKrOXmpTfU0Mx2BvUd4fLUSzyVpJz172/6L1f9P+NbE
nmpKz/Di1UEpDT3a/xo456Dp048mKo23pTYuWkpuJIp2oPT8w7OiBLAEaqE+zOMs
5nwlnZAc6JZhVUr9iAahbot8izt1e7iqZGnRSAuF0Yui+ijvzcu6ZFluSuvLf7x5
0Ebv3QQiqU5OfIlwwkSsX2bpg2XmIoGDY9dDxHjHxL+pQvA0Mufn/3+eBZNv7AOz
/5qXWoB6/8YJfoh09/OovphJuYlxU0dNvWd5qQUhbd30ZH1v+dfPxeUg5cNU3IvN
+ovjh0NAgtVO8zazamd5460baKQTI4uuJm7Zi6JI9G4l/eZ4UJP+mOWH5mrDEyTG
Efu6o8iSOJqKWNU55O2Xfql7MVmzWJcmKt+kjJP8dFqfyxEJYr/oTIFhFk/N8jjq
1KPYMEr4xapIsJPXXzSFsZ9fTcMThGGX1fWXB6nr/ncxPo5n/gQNrb2bIeJhsHA7
ZnK9xHC/1+59nun54im779BrObFH0sSlVN/6CiqykPcsV3y6I37V0zCP3PPWuKig
L6LcZqjbZ3EhOCDOVKC1wfcFe33xLd6H9+FwUE/vuRCyLmDMGHNRYSHD9fO5hzxu
7CAndbpiK9GHpXGFNCxtgwGBLTTnKWNGbA+B8jXEjFY27xewCMxlu8somc9h7Lsj
heny819Ao4DSNFDXHZU6jLqOjRr+ti714uenfsjg9F+7IvOxP3b4YvNUmojCJF/c
nQY/UZWqRCZapNRbgI2JiDSQ2aJRh6eDqjnQvWEfgyK1k7LYPxaxywnD0agbFAhQ
Q2UmONSRvqxpM68l81jEa7uiviAVfveKldrZ4pn6RPc4DlCHZcwOPsPzk5bGSWSH
ZLc+PE0D4uL4JR/Zdptn18XZVqM4tZvig71UnUfVNPo3BfrlVbeIiSlZO1DoZJd4
aFkkBQPNXz6PMR3bJLxDtw0xk1Hsl0uJnmvzLXAGyNziDyRhZ9MdQpVkaeOWS63I
vLxqWCXUFhFK48WffXl9r9Uo8upM3zldNEQbXXFOyxknkKFg1+vp3pHR96bcvIaD
t7R1DMys/BjA7RCDR8TJGddcz42t1kQSZXIMXqbDijPVLF3LNHkjnb/w90aypuvY
uqrdSJtf+6osGKp73Q9dI+FN0DHIBimY8IY8COEgUYRtxlDGjhz0Dn/FiwHCckhA
OeusNOM8BuOXMMGjGOBdIhH89LoW511uHO/dl4Owsqs/W0/hi5QzfgyXSgRR6wpj
h6bkWio3K6bkLJw2XTJdYmj+owVHuk0LIPsj42n3YPQca84VnEOFxthS8zdNdd/u
YOHz/RZdMESnoxs77zvoFSz1tILyZ6Fb2ktQ71Q2u/jTif731tE63B7Kno29kezK
suk8vyWvKIwd5h+dbOI1/3R0S8ETHN9DXBwi36GfcEI0FzrsvnXrYPE9kyDdBBlw
RGIvpS8kBSOg3lxL/cSz25c4Ed1urnb8ZzF6hA1n2F9+APTFl4tGph0NMMIUaDgw
cF+SUfhOw3P/eAscZKmiH6VHxNFOnC0KqS0cxAzVhPwuJJ+ej3aYXMaRX8asWp0K
2NZngvUGoKvBSqqBCySJU3lRm7OOp+fAc1hdYLn1a8Jt0uITHf02OK2pnXiMIw5m
HiJVs+D7aMz//THoHDRv/u96yOWahj5zq2Lnlafa2C43DS16C4YajNqyR6Nnh8je
NK+kTHDwLUXe5xTJaesw5p9njcqee/CYCjGyXU6cwrwYdBufRZCvCxslihfg6ofN
ZbTZWuUfCo+dJNESOuYbsQIhnSUxlsGgMZPf6tyinXtIsYShBcPFql7Ip2q5r8e9
xZvyFLTEfuoSxiFuvVzrLeSVKr/ZBc2+T0UFWUz2n2m0fpjCatThar4aIAFxNfYv
sWuNYHmzeMPLqXtgjS1bzjSZpZXC8h+QlPulxoluBnbS2WkVI5xEGdcAM3QuhGDa
5b4mGM47wmkJCG2XNxV9/TUqOkmdytmOvVPo5rh1/YYWVoBvQ4hXiwT4uOBmxvRm
iCCq/ChlLzveb0obvY5pzM+Ip6GcPFFplY20pVNM6fG7/duBJNHYElAIWvI+tTCb
0z8vbVngTdeWg2tJEI5d068P2QnHb72478WrnC0qoFXUWYQRdQWIm/nRfnSvT96u
0WY4J0E3A0bkKEmWqfyIRkzeTodUsIYdEZOfXFANljlAkRDfnHj8LBqKYGPRFW0a
xjKuFeAvYM8hheBmKHrWl0BJmry+JQhysyqnKK2kETJxFh4Nhx7qbGqkjW9zfSRu
nEU113sPbKZsAtROoXU58jdfRQkN8456r7Q0VAsjH/VnzC/y+sZkRW2Bs9VDIr4R
u/C4b7uzgBdIdRAtQAatP8hmGTamynNCeCABucLR8ZEutUCO/pUAdJr4ibCgPkVg
cCf/KqTJ+sy0sriS3rOqw/9lCkoR/DIeLeeZdZK/L9taALnZeYPcVKdYkGEHG8kU
mHL74wmiRFQbRf51y6UrKNotJ+vOHgzDNLmGhudXqgeFXl8Mq2MWJOGsEoSubc8c
H2AGNbW8v5R2FBlmAeDXRDqLyWOWzC/gcKj4F37OVijCC7uZ7jUdXR51DjfXeI7u
Hzo8ymUgm5w/ZsFxD3w2gNbN73nM66UOsM6zyZHuP9znTDqSK0P9KtL8QfIlFJLQ
FEarIybhUdf9P1IlijoA3JkvC7RNqvaHnVU+aa1v3abOmzcclVCoZILDi3ZhjDBP
roD1hOfALCaJQjPs8SD7ekwIZe2iolIDZvxTRmX7rKyuEDAI4x6UROXQwiMbp72e
JFDOtXvakzVjxI0yLyLRKA/QErGKO1F5VnfC7fK+S/UExiTfSQ3xiRZuat2iidow
SilRMFkscGNxJpfTSQ41b6rHJ7ScnCbdPl4zDtvKqBd/ru020i3Eo7HEub80S5oZ
d2JuoovmMq+iMO4tZUHmR5B1XqoRRuRH3XqkJV2hFgqJuL8MDU81YWgTs240R23F
fym/GWu8/181mZ8v1Whdf6RBS5z77hXjosGsgChG4ZlgQJGd/lCQfjsK/8cUf7qB
XTsgIV2LVSlABL+FAIb3uCSv22VvYCu5zxKC1X75FjkFWc+3x2ONl9bj96dg0hPq
bBPzvfXSYZwvm1sR7f8x2wuxZBW3TnMFBL6lB9KrnJA+aTHhL6OxktuUMg6p7wal
LGoUbQMJv3vyKktvw0KUmIXHFSRGPgavaqGLq3tyIMfOgZUICu1YUYrjbQiPnTYV
fSsJYgekOW5jQQlHcg/rMwa4OrTOooVN2DTBY781VY/lc36IdygdP+Q1U5UzEDZ1
pf8Fja1+oPdx0ot7yR4sSk4HZmVRhf6qFy4f1Ebda6eaun2tur89GVLzklexh2CW
qIZSZnnoXhILTw9ndovwdZLr+Aq5Io4Rn5O1TILf4v0O1oIwzY1s8YvUPzcXwXgx
x09KNoaUnUrxqHCtuR8EerKn9xqYD4CkRGYo9FPg2Fn7nqdQoN+pX11QxWm1KZ6L
vCoSoLUG6JTHRul+uoJu8ZwmIYkVWv2w8Xagdn64o9oYTAM0xoHT1bO1r1do3R51
RVa22ei7BptWEacvDJwvwZvuveKcWkm0xza92XV8P6a6q71teMzFKERgVyNfFepb
v1AlCSSqSKInzRmN6ebzr71aksujvSfgvsID/l8sIaaDszal8KUsn70xr3klfrAu
yNxVv3cIXhMsWmPROpztH6AAIaMzM1ufxnertKSuhuRTfv477t4W7uFzbDzzc7NR
ELSBVbwVT6YHNNI7ijze+WitzElQGV8BlZ/VHJ9WRThnqOSjU8rpu+O8a96bMt5a
S7vlJf5ZWFOeDA0zvd7ydoLh/MdzmfqT+Cv63LKAiTrcnGrKpklkvKmcHEDMPL3H
tBr4vbtyl1v+VYn5ZP3ly6xdsgyiR0NTdeThYQULgsiPT43HDoPO9V6p8H1Mz2CV
5Z4Biyu+M0S6JftQzB9mV+uXjOdEvdAXzOCP5XnvWZBcD8GMER8FFnReOZV40THj
KDV/czx4lnXZ8QUDtUpQstli9a5oGtMcpWNmlm6oOoB7Auo7Y2etbLAYQ3cyTvF4
9+X0DaPcRvlQ9a0C8d6dSXKpLW5/ccX7H2ehXnvIuyFyhVs5/uSckz0YqjU6U5NC
ZzBMV2zqI4zQAbzFJYnmahrEXSI8lL1exUKaSCpUAcNiF4B4LdL58HGswzJwgtze
rpdV6e2dBJ4emcfoN04Xv4nxiZTDGV54lt6wAkDEQMRQ2ey9u+0XC1STV9XJ4w3A
cfQi2LPE8rspwzLzn5Jf8lrFGjn8/pvZq4z6ZR+91WXe+G6nBDQfWMEaXjMiCW3f
O08h6PgQ37alBzwb1/ZxR89gT6epC2jmnrLQHC/8ZmEOt07hCXhwKr6gXrIpg5X+
SAs2CZnImngxqLOe7D2sLa6925AbfqPmjwIbmZrrKnYhYYAzWdf6BpTG23vXf+ko
zunjG4Wx74KlhwsZo9qyuBJLwDOgJuQM1gnlN28m6zKf+zXWVL3dn/bIfiWgl+M/
p3o8B4RKv+4YBpsmEEWiB7/tsrq7w/VDlEqkO/lfQT6cWzBUyqc9TwnMW1jHM3T6
h2sJwq4PJ4+f4wvKkAM9A6A68Hg0+YIGrq93n7ZhNVf9FQhqz0XNqYYWDa/ulDl9
qHMSCEftIXSEka0Y1c2qvhya1mNUPBiJ6yZhpEqo05addrG16Jhazxq2HeT7vfCk
AGiiRI4a4oed7jKoDgQtVaG22GDoiEOXdJCNdSigUjN3at77Lq2s6Wazof50Jg4t
9TP6UviAhFP7WfYMyLa99X7JcUUIB+zaKUEEUU5L4Sp8qZkqCBMhCe9XyXZ7oc/U
yBBNPpVtpaq0hhG3+3d45T/T1YMhqes7DQfN31gqnDQBIsnmBIhQa8YseQZ+4CZ/
644zRMh5cXM2XCHSl1pFMY4Wqo4zKZR8GUflx5EZnI7F9QsTGE7rXO9d7h1E3RnB
dYu7Ny18iOZ9cK3o8mZhOHkoEQOQOUaJbLfs0C/BKNi9vg6S8MizuBMMqUAmVgoZ
GzXyV8JCw1PgUGc84cGpdP/7eDMkxu6PoYxCjkqupivADWgzj+FxaRlB+SZaw4ew
97SomDqTnFRbyYQ5gRQgksDPksi62HLXG5eiOeC/smlaAkW0izECkRqp1kVtfnJw
DNQDeMWJMmOMC0mJz5DtExoH/xSL9EZqFMZtTsAGNnt6gtSJmCuqTs6dUJUUejQ2
nRJYVuHyub20vqaldqPy9TP0niTj7c1A+d4gOiVhSxZ8xC4gRRE3qCnMI/x6VhQ9
IhMQfgaF7TGSwzmTMY9MS8UAGYahZO/74dK9c9lgW8d1RKqYpZ0q47weAXXSK+vA
KuguLe8eI/krKE9pVQiRoAIWmwFmwUqP03nahzqKNCGtxGXeg8kIegb7qz/5vgpc
SwB7oXiKWEYicq3YyuCLQF9so+qI8WSfaHav4pRBBH6tIYgZqnHvg8ZDktneYpcS
gyXxRxGrUYQ4hOkg68T8Sq9O2sAH5XJZmmqfYxdKbD3BW25lMhDKubtTWnp8vQV4
rU1IVS7Maa3VjpLwnc8nYu2iEUmXRjpnYNvL1wtxuh/J/FEIHGNMfCyGcwIFtjxp
t+Jg2OQ78Aq1YNlFSS3JiefkaUOiU8R9xNnPDXQsuI97cHdYqjCFuWC7C6vL8QUe
xWNdJpOPFwdIS4U4gHZXv4aOWTXX/tWoeH75acKJKYOImOXv/MFFhiFsPxfS/L/u
j3Q0Sgsx3g/L6fR6f7Qb+GVp5c+FvNbkcLhasTYemrmrgjwSSZ+dqPFFu6iZmBxt
LKT6FOlQVddccN40mzoWl2v9qFOPTHIFTwcoBJ0bPflSCLX3ELI5MP81fm7QVU+E
psugsCdnUOZDN1f5H55BzG7mWd8t0UuXhGBKD1RxFMw3mAgxVfC2w3rioseBvrC8
oGmkEhMFkHOdqzy+MHCNOQpPafCB+zPbOCN2hSouQYLqJzjq8/du98fAUPThMwLz
bCvth+WkLkXfld8m+u4W0AQe+d04JwrCX3RJ/U7+qLgch4d8lA3mFbe0wOKAkZ5b
zRJDruYKHh7aKcgr9gY5uG3HVNuWLy0mAO0DenCVTKD2+YG0uSwf7IK/aK9w0+g3
6IVkLS+1nhD7QhQPclkGxTgTFHxt4wp9dsF2Bl/j4RfCEE4x+6GzrwN3NYAmhpLT
7LZ+YURIHdo/Dd8oFQeFZJlb3rwH5od66GDgO3ZQnDUrfeAP64m4jYoAgaV3ItGS
BcMoQtuKG4gAD/6bsrJE3Fh4zoch5r1UkKpfuifG68dbs6N4rIi41g7JrQhjJJmM
rF4VTv7qWE2G9sFrkVA0+vFRNEu6jgpiSfdF54M6dZMPwpwtrg2E8pJXx4qjmz60
JYxTjpI1cMaNWzppGcHAUAUgLqgoTKf9YJB/NDiJVNv/78B80GO/dZ7x8rDZSB24
3Kp61B9JRwJntxRVsQBFjs8VuOfoNl/PlLpZk1IEYmXN9/DxMK8PzbdzhFZirVVh
JBB5kcVNVFP5mjNkSPIDNo2a9XOwRA4TuZ0KOkcF9AzsyIYySkDbgG9UkysmfAOD
c0McK3dwex1EawYLC209qoTw0ft+/ySy7Unoenz0ZEk5Jcy/XpzbT8wmrWeUQ7DR
Qwvyv18LEtCdRMP9IgmfQuXcXCUQrgICvdPp8F01fsvIDoc8o0bw/dYwvT0VB8NY
o4uJ0AVqJKCxMBPA6y2th86PtExVt2M1K3Ld3taoT9A8WfZw74R+JyphmYx3957g
qjIGWddQRr6AuKhAWybeGVoY9x6kefW031XmV2paLTZ283vS6iK9QNfv5Ok/wtec
uL2d8r3FCrVuMmTGuP7l7pWz/Ob3+7Ji5ClKfexODFCQQ/wvc8PHdgPX3yfBC7DC
HFCbiExk9abXgAz5/paeNFk3m3AH8YUJauepq+O6cMzbogHy8DUNYt6TvvlVTDad
1zRyuGU2HDVES5cm7JNe/qoG/m5imlMHrNlvpjIOBEvFyiZ/bMkgYJqihcjEhO1w
W6uZMRotZ1J2SIQ3l+fF1pJrKem5ZMb28QlAFM8tAGy/8ansbt4DaNDz9FchPM4K
wG2t0tU2CvD+7QXtVc3Gz9mNmD4qv+OcjgyoazIzcqE31+/eCESoyu9hHe902r6y
vn0RpsOVX+NAKAzmhFNu0wgfZNknxxfVU5TpF9c+yeyQ6pMQpMCnjJ8WFCK9snpd
NLxy1317DtE2Gmlt3CSziy9dxa5JxbSrLT81mr0Sw6ZCZZjzy3dS0C56+8tNXr1A
fO0J9psiv//xTAi7uK2fjBWcZ2r/iaqj1elRCtUa5NM0YILZTu8XESrAynkICgHH
wDuWAWByVSwxmw6OBVVbqtayuqtU5V0yvkuSOBR70g9rpjqFRMhsXkIIS8zDz4sl
EO/itmwdHzil5g99YUDd87m6VjtNSwSa26PTsQwJ5v5B0CaPiaAhG5EtMxpa1UC3
K/H1H7sldjLYtSDV/a+f2Kqp/T15SETQbMJCGKYPOR/zgMPC36MVsqhHtWPKKwhp
ae9Znn11O2j7pVZLfwIhnY3GX0yX6WnJXq4ioSxjCyfIXHWRbXcOo54XUxgByjx0
yh4B2/dezBke4YF4dWBCeMaw49qX/Qfa/onetYzNGQhqoR2ZXVWC15tOpUW1z228
RAiOG24Eoip8Z3kmekGXMj9tqLCBhLGejS+C0V9G546/EDW2EqDx/Q6tIZ3apwmQ
loU8ItCgL0kDu4f/RZBJQrtfZAWOFzQxJT21itIh219UJN3w6y9mZpIbOy33Vy9P
1GFSYdetMey/9jRH1e7IxSxSfXOdqEnvvq0aUyHo8cz07y5CEum+a5oiKE3TVH7B
Nwy3LWWKIsZUOTTfJV5Rv1RoUU/kHvSrBlmniSoIAoDH0yHgvBMKh55AMlOxBGoN
vF2SHBY/5HeifcxVKibK17caAnHWVFFZVdPoU4NuxEs276RZxavSf5PToUds6vEy
2tGVTQ2Fuu9Rgil7/tTEq+GuWaYe4qG5RvbfR+y7oAZwsT56b3FNawC5bvs1qmOt
+84XYxj5oJcbKpHmI+ob94t6tyQUQwOeRx4e8/myQJ/lwE09MvlARaB4tAmvs4OS
V5Ad/cYU+BsB1Pj+qMG1e82iMmN9Auk2YeNcTl01+f+jyqJ0kGcRZ8r1EuCeb1Lb
ihgYA+FIRVsQmPesHOtjCN1r+H/RxgJL4caDuG9YXfoEKLJq4mwjZaBZ10+gwUbv
mz7UH4FKYlsYkizxAKJdT5W++Dv9WxvSSRv2Wq31vCcVHtHNdBluawJgDFsvVct+
aAHCHFLwm2D3Z+f0MscXleQHq166zdUXsWRa5W6DhzuAFMoEt9aXClmAORtt+pIR
uyIb8LWzw654cFFW2k9k+IOlSAgcIEUb60gYXwrC2uDZ7+jEYwwanZF8icGgynHj
mrCP1E5DWaLAHiVroMHGbCWn9LmCGycpTRmU0u7YKs7FjC5NmeIsGCE+MUptkCvA
Zt94M+ts+p3oy+zlMsMMzOFfrKQQHjWkTdSQBSNg0AtKYPeIYzuopeeFBfpns+UP
ZJoulcD0FrFk4KJ58Beo1w1ns1i1va4KedQO8Boh/9TYCRuHsRgu6lurAZpWL8Ji
RwbvFZ9ViEFbjIQCgyE5nUytmrey2FS2CHb2bXZ+SQ5xQpQoUmDW8JE4Tyl+znv5
vhcR9dDGVcKAzjOatZ0g4cg2p2o735Y0hZB8DMuOxE8eoLnAtWwpnkrUCTQu2Phq
T82gbccTs3unxHo/IPCni+iUBOhyiOodwQWub00MXEYQ5FqUXy11MAeA8lShGYvC
uDNJIIoVTl2TU8LxAHIeYz9FUxpgb2U9/rUltcFcrZPm8/PWUqhxMUXPGcK6X0cK
fT9GCUbntlRpW1vPJydpPak9BiMVthV6SOEvfVSP5u/PR03l5iNV9WwRQhf/mOY/
Av+CFhI3lPzQhQCKrn4FsTL3f8TgTJMw7nYEyaK8nyBx40TOJXv/hJihSnNOgc8a
Dz4dwvvU1zizJvLUnj2IUBuQmd9Px0qRAjSotio7jvbVrWqRd0zFJ4gnW6lyhreC
NgDnCPT1ITYrWtydqKt1Gz85jQtbsFxSbrpKag7bRaSBOrf8k6h63Oy0KangMF5q
xRu1UsxHIVYqpD31870QZPU6y++SM2PptDNixcVGTuyEgAuCVxfEbIHvmmMT951Z
fip84ZzK1DwUGM+CRJdFGOMHCjcTQPSYUdwPkuYUofv20clWW6PI11GCDER9x+ur
CI8Cr+1cbFREepezZE7Kdn5UxCe4kmqTOWzM1WEw/db9eHAA16ZLMOdJkJSD9ML8
oPIqlP0xRoCdCmeO/2dlYhyZXPj1e4OJJ0xPBiWgT44JAOfXrjupxW3FTS+hnvSs
f4O7dVi5fTb1IQY7M9Os12oLEmJw0M4nwqCplwFrU5tZwLLEzdJCY2OhSvZNRyrm
trbK4odkfGUQtzGBLzne3+42plecHBH7pFVk9dhiltws21mTKRGWAcd0D0xyxfN2
cfPwHiXHEF/Rgrq2c+nq4sahL/P8RiDTe84IkbGLEaDNks30mQ9vW9TVhSh29tVK
HYazjsdpAqQKMCvrSX5aONf6nb29nIZucK8ws8Fnkrpe8NGn+IWU+0b7rDDdXX+U
E9xQFbIx/v2YShi4zV8rIehRdO5cM9aAILkJoeIlHuF9RPPIlyH/dEJjPCN4lOAm
/vLBcHDy9bEWlLZMifPye2vHpJCgyRgsT9xyqUGQIaonS2m77Vh00aQDmkJVANPM
LGQWrjvO2edchCLG3vpFuz8zTGvcoRm9TjR5qCrOKPOzSqKiH/9Es2/31pcfT1E2
LlpEI9xcSpKvW2yPV2+qtiaY1ujAZbAjFo0nEDacKAh1dTrhy1jMporIcw3c+L93
7jQ8xn5rsQebxiIFhZdr9OajKaPUBkQe1NB7AYgz2+VCSK76NUWEZjgkGQrSqigm
nJnkbLl+aFfYwWAJBr8f9pDwwoUKfMjVWDPeagHfi9WubdMraka4ibsIqHCBGEOd
Wam6XQsALOAcmCSpljv+aTQ4Pp14FF27utsd83jipFeB2HWEY8v+o355MYKEbHCw
sh+brtURMlrzaRuWe82mZ2rsLbS61yXbD6zS5nThHlILswTKMsMp4StG0+KNcerF
4A7KAbLIjwcxQpMyMvToipJUkQ2zr8oofY4FBy6U2CppXhj6Qyr5AI0MLp/r0QjD
EnRPrYgdIFAksGZGgRYVCp8cg3saoK/Lyq9s1bhn03jaQ29vBuAwqNm4naHLmFo3
dC2eSCECQp5snsbqlo0Q6OtB/AHSJuGdoOy/aCZ0rS8yMFa/lEt9y2qbbZN8y3tI
wdV6xKSUnKVCn+42ZqPIcanFy3DZ13uNb8TQ1oElABBuvDDvnJ63+0ClU9sy1kOs
ymulWx+wLnrt5I673MmIN4SBglDgFVg11tsupR+1Ggec+PRe7t9gJoRMQrUPc5M3
eIx1aBsvMPsZpg7GUTO7wuywvJbxT5C9mZ26mszxf8U38NUcgyhnRGgwJG0bw63q
W61e6P4IY4Mx5l8f/yQQPuIyBoidqR9sHqUbDZp8lSdlP5yCTpSZKxZtcCRnfAEB
NSKIOw2NNwTGUF0GMsKU2nbZoh3d+7EjUDeH4L2x/CcNgEVziIDONeAoo0+routH
CAwbCebRbGGqutCUDxyhivGYFpmBE2qJH7u/hDNfgjqzEmQb7+/ffyqZuQu/Fqyd
4gwSQ0FtheNqElRFc4wWmUOZkaxCdDDIVHe/J5HDpo6FzbUDy8ONm8FPuJBQGQmP
rP/ZqpTjepgPNQC+jaTAOytNoKBcd4rLPedQanVFP6JvaMLtXHY03n4Jd5T7JpGr
xc40ZN4cKS+kJzLQsb+jztbh0m/0ym/Nrm1IuQjLxo5TOFhYAcMhvB3TF0ihvJ9k
lE0UFfexk0l9IYtSEEQE53fc3tWzY774O3mjo9sG8iao4e1M/9+zzPz2VlwD8aFB
+GQWWHS+pb1xdX/hMFx0B5HU9wGK+WVslmVcGpkOUnQ2cnVnif36VafxwHN0ffAZ
DLWh/pvpFrN1J0tHejYlczzMpQ1eAS5upty0yCQofxDL/9wJqMh5pGCDTcal+IK/
Q06L2lsOHqWcvuc0eP6OXvo5lfbF4kO8DkrNuYsd6HoYq1ka0GNJm1jB5rXkj59V
9xq0UKacaaRKSFPUX0zSEvH6yYnvNNGYFMohuCC4+bP2/C0la8uDqKN0BSGEDuEe
1pEmRB7lokHKkutaeHw14rwIYnRa4JJ87zguhUZC/aD3no5jfdfGAiXWobqa+tib
Vv1uj/lfjMrK+g9wCuZpHAimMIa3zLN2ELS148dN6kTAuF5UGtff1mq32Qw5lruu
82MWfZycOcEOtWgUTFQqk/gIry/Fjo90sRXg7DUkyHJdZvteupCibAIIoGGUXDuN
XsDb61Yx4nsHm9b1ufQiIY+h7wr+7BzU4PXy3j8mWtvKwopn4r4BbsbFu80bcr1n
tCSzgyrybyX0hiNcKLV5nK90JPFwAy/cYrtYYhAuAvI59FeEZir9KTG0OB60UjQr
GGxaF5rorANKgbvm7KHIBZEAq5QD1DN0gdlEflts5JtvqjsVYMbevJt0mA1L4JoZ
d7gn7NOEcpFU+WChmJ652pZXNiKluDzJLIud+nrIuxo9l+TwnmvbpswSdczGlLAp
SUJQ3DGzdUnmiH77MIBvJf/TLukZD0fj8QvnGi2Q95UEUMN6fr+aWUG342urDvW5
pjFNknjFA3P6nKrAS+VFsgPVXWfcBX/DRW7ujJ8lOrYlb3yDGNjWtVKxDi5TC/Qc
fGOyTbPvv/Dfy5L2IqWqxvGGKSYsS6QwKVpqXd6FRrgUcTsPRAcoSbBg6ogOzlVq
YXkXDqvv/TuUv/Zoyq/vk6f3TrQ7EriH+HljjTC9Didc029oVya0lbPi9+2BX4X6
fmiHK6dwAe9PSwfAUg9DwYm1mNu7cci3fODIW+L4Ye9xFhGOMbPKn11/jAX7tgwD
ogUOCyCxSYBNg9YTzB0zapmJ/Vlkj/gEfIg96ecLuXF8VMljnlxSCL0SVlWCNisu
Z6qHM0AHP5Yi9Bv4fugi89sGDOgbC6imnqQT6LEfq7HJ5GrZFf6rXbcmqSbUPBYz
drYOesR92kxCQ+QYkEEoAtUeP1QE66mDzDLhnj1XroqKwSGhwc6d/gxpH73nSMqI
5Ms0ZTOIwJrri0xq3HMTtj0VDbAMmnxzPqIZ7CFo39Kuwf4DQOqi8QDOntuFc1np
iJSJW08INtjqd3AdSWz9vQ2caY1JhpTMYXCxsyDe41LOMdFJYrc7gwaEaxMnLq16
FacYWRES6FZaLhZr58vuD9w+0COR7gfD0s50B8BYVvR/fSKTypC7/tmaN9dw68kH
Eatb6WkprhnFvySqUHmfitPdQR4EyVAPRnwHEQbk2ymg4shTgnWcFvx5beuRTrzn
2epW3Lzl92sI4w0Hr4MmcLjGUc/uLJYZckoV0nK47+N4u6yxlQOmPEYGcGEsP2Ts
vSFkM92lcodg0gpGJAca6swdvG3ftia9z9VOxrzQRRrOcNrm4EedZ84NZlxGkAp7
xGus4w8+chtgngYjTEwjvMBXIOEGgUUMVHkyHGs8abLTb1WhnHpd4P3TK07xik23
QHsJgfehirmPPnPQVuQPll+K1iePPxmEeQN+M1MlVZsus6C1mLSH561yB4Fdqjlc
dZikuH0S2POW5x6CHiku33lbE1TzrM47Xw+PQYUVnSi+88WGYmSYuI8sxIzWtyCC
S2brbkIy4sV7AnUp61M3l0nuKItunIKNw1lAAirP6o8qfDYFLd8uGOt4Ps1+c4IP
wzbr+U9QXaaudWd7RzkNNuXHuVNsYlU3WMGzJ9JGIv/2v+mw4+xDgXGaLdDQ09WT
nBLXB616XQVaS9My0Zc5enJyOnaGxD+1+oYKGVDhnt4wKtjS86pasz2vrjFR5MWn
M4Or4wWeXxD8eWsAgQMPoaZZqNTtA38hPXK7tuou1kemEdRxZfcOqM+d9yNqHcT7
1c5sTRqhH8PbVCiy2uxTZWP5JrXJQlYIWkSDFhpCB8M77q/1kHhL1YWGLaupwd+O
4oMhqbjN9kWsXcuqnzKrhP7esMRXO6fKHs1+MbNyKUqosFPuZEC+imMJxFcV1OKm
7Cq1ax2TYhr+imIyeYrG3PCOz6FRakt4ngI9s/UwTL8zz7A+Rz9A4mhdCJ5vdB54
6pTTMkTI6JzSAsxSr8scOSV+9a/N4S0dHotDV9G3ZQEBvNRrgAK6c6OFSjj2mPoZ
3Gv9m4+LZRb18IkAI94aLOV+GDpaEYTPu4IEEHsu2tOFtghOxszNZazJWUh0A7eS
qZYj+sjfOBlyK0IPVPbLLqJ6bA1W1va7ioAAT2L48gFFT5cStCETImavCcMQ8jyJ
b4qgzCBUan7gAxZDnY8NTYRlVohIPs67/drJnh7UfS5bEuzEMF91h/nF6jT7HFeS
16fVPq/wvuX5IEaQE6k0CuU+6ZySmK7khw6ARkHWWNG3eydGt08dnJAEufLYLBRR
zk9LZt7SOHGP3aLYfXJycL3vTY4OAUEQJXYa3QvwXuZqg0a2Z+GWJXxZEdtTU7vR
LbzchnyUAGQKO9t1euA4rphUQoezC+Fzip+MmrFirfT7+SN/30nZ8CYqcwlC3NFf
kf59orZMGWrVn0/r1zEusF/AkDmuXBQOTg0BJntDsd8j+9gBOq4SwpbsY/3hEnle
/dgPAnn3BJWpcAPQ8zoMR8mVuvxRyB/j8s9fLRTlcBQliIPjdhODc9jnX0/AOQo+
zP/zN+B1Teinxva7oKpRa4rtRKgjMr6GOUnpzxPUorw5uQwxAwciFGnZG0yDyYXa
PNGhX8EFurk38AdcWSoudp3L+673y/3EvdvwAywHTY9Z1dfIFpPw0Sqaqsrx4RDB
gdMNBCBrOEhFLtQ/72fGi8+BfX7SSQdeMbQ0q77mbahUE8d8WOHjp/8syUrPzok4
aKM3XC48zZJtxXy3b9qun+gWx1YkiKwsDq39v56dQwKRBucbRwChbl3w7GVJJ9kq
ddmheHRG4qrM232OnRmBQopuMn+bHYjdT8oJQOu5X379rtja+j8RDdwaWcE1jTEQ
kCPh76jwVqJvMLC3/scP7wxpOrpQDaaGQG6eg3t0IqgU1AG8D5+x2lS+Ege4Q3KA
MNpOajlIIOcNzfiO4Fi3kQmgEFXBWqgYU3/wr2XU+Gtn7psyXgykgLghcQOjJ6CZ
RjGKHiLuurGTlAcJ9yXq4a5K95GPOaBkfi6GTbmyl4osmTSV+ewrZW9FRzPzIT2Y
EYpG/Gm/qLpHV2NfNwp86ydaYqhed1f4651M3W4/sx67WDywaLdVaXEE5Dt4DfQ8
6NduSebPeHc6oBV7op/oGZ0pgkQHBbiNjjl/yJAOzbR1Zqpj1qy9zzjltxi53tq8
iA402s6mJGP9k8+UW6bxMVgfAnY95wTL1y1z0H+y0W6QWTn6Fz4ujJRJ4jlFBBJE
N0JnQdA7lqzn46rXD3/fAp0TloRtifmvLfxSX8dWe0fSyzJCj/VwNUTdKTuQCvsr
5yF57TieeoLP2D27Q4PbkA9aptWiewMP1p77UzHMU69c+mV9kZraITSVEKyGUNI/
05Up6zoJ9RvcYaNpTYKOyOqQGxi3Y6irbSPK1oiXbTojx2qZ47Y7pzUeG7xFSotS
T2/2N+hg75LX07nscuabq1sVHc0MB3mUGYzyKwyeIwuPCDPrPnmmOdPYpEnWQwNh
20yh6lzUzT1/191mJP8PW7CEoP6AWFWFmPL4xtrGJP9ToGXwv9cqJY6LBOiBswf0
ZM8XfS+XTeXikrIcqcegvDws6fI2rJqvKQoLY3CZKt1Aiu15DUqRfnBo4/GebGZb
ESUw86ZY22nNjIMhstML/AMb554Vhn+heyti53FaXifqeGfWIyNqoA51LkQhjxSQ
KsU2ICZJxPQITBMndY8sXpO6hOlKIrx3V4FZ9IJ29ScSES4ueRI0JZ98JZxJZfK7
Z6ntxliL3HxQ3u8jPilK2DVankMMxUbKRLd8Tl0SnD4MKnBFESgznu4afUjO/NCM
9cldGIYNpd+NUNs8h6pOcR1dbW2NOE2fWraGKvgMTBCxX7OYU4+QX0xit1tzs+vb
R8izFXniVe9YmH6PeiM5F6oALx99i1B+FQt7SYSgK2DjuYp9zh3JKP7wXwwnSy9T
feMsy8LGZXUC7vKJdE1YiBHKuPrtBt+7tsZDdgbVhyDibrFeGPyAVYZoadmySNxn
wGJLibi0e8bR835VldRgC876RjvgS9/PxCBVRkezguzOw4hI9bG7h3WAKtUzXdDP
onyTZzjqLGU3o9SmYR2Agzc3L4sX8w7aIt5ZgK6G+4IRPJjNB+nTVB49WG9PzY0h
/GPZzdiJWFFIVCBwsaUKdy+CAIUlQSS5dtSXNpdOO6atNgYdr3T/wv2xU3uMH3vF
bGtgNrTClovwzGwzq8nfTyYngcwY1HJXoi/hlwlzWlFglofF12OQdmO6rYTPijsL
XzZqqTXF526LrrwOpvEXITDQGF54ZA0ciV1pOK2UUegByJDg7tQixg6wpZS3qM7R
mHOScUmS4bkdpUZ3KsTrd5hnMQZmKUd81g9sux5bWwaQ4kxd/m3pMEMU0JravrY0
q14abyb28cJt1CloVJDn53Zjr0QWmt6yhh0bvsGxbsELxfWdW3ZvXesD6cjFTbQb
CcnMY7GSeztKgjyNCwk9dRLXimFMQjQ+Nq136KlzNc2lHtcMtHzj1Gprovi7bxj0
lAlu1aKA1rOa+lUiE+7rOWSWbyTa1evHQ6ZFb5arokTMUB9gcLEOkzQmfMr2kG1C
SUZ9++gOVFeteyAOOImwwXQR2r/tbNuAC69X/+wo95662kW0KjJyvs0scst2sYNt
H94vAZLjl7eCCCoIWfybdeVG2l6RTV+LVAjlpdS2IX9HK7nS2m1edXD0xPwOVYt3
0CYbaTIOCiqemw6OkqHrjk//uqJjUY4Xe/t1QLbiJhtV/EK7SgfJJAmP5tDWE235
NHx38QiMldzf6CFCqSV7RQ6dDDJ35FvmZSVISZAhBnkE5qNfmnGh4WUlPFQMWA9k
reLa1KE44LpWXEUuZFLaRWVx8kjoPgoML3wweCWjYgrPZrKDflyy7SLXBOCGOIkh
DK7vr78JVPeHYSkISPo0Fc5ugdRavCPXzRfGgUB74+/bqca5s9GqBr+xC+mCjqhP
XYqMNG9viz0uTHXX2PxBezm8jFsGWxH2bpSxP2vMHkPB9WdsMmXJz5+JxdjC27j8
tqY0BmfXmg8nkwrxoPUUYqYjtPMMzLtdMLWLGux7LQEzdCG/ZmtEWvKsOvBybLR3
3dQElrhrsURKIN+8rjZFgxurJ+RYbLklce7yBZ1bMft2wAIPs2XK8e0qAqk/uxRD
EX8vHIQNgMoljci5865Drgwud+QhOoQ07+bGciIFQmNmQt7JfGqWg2F+eiQVmqTI
y19m48lIMS9yoM7q+Q1INVnfhU3MjENJtydpNI/ZlxfwzZ4UF9O2sf0cBfLnbl7T
Mco/7Kqsx8MCjRyHaspjQqanX9yR1aG0C2+6j1Nj8xGO0bKwmpJb98WZmkKHCqaD
mMrikZBLvHm7gwVjwYBnjjhOBonegqtUzP+qohcekFKZVnURbjP/jVtH5X61O9h3
jL/dGc+NTz2ncsTLfvVavu4BrSYAt4sD+lDpo9/MZugzc0/gn5jZ9P7itcwns55p
nF857eTlAUQS74l4uV/E9Ip5ofE52PytfP23PwwANs/1bTXOO+UGbtKgSB4+Cr72
SmyzMHHSPkfryQZZZVuePgrDo30plfRmhna1AOH6G3J36cC45Z/M2YzGfXLSW4MK
IgAL4h5eVvJMTQSe7pKkP/UGPiue+IwybPXxSrKWwKqY8obOmP5dBUFq8Zkgnbo5
B+ZztaXFIrKjCg5siI4WaA0ShhaEOhTa6lWX1JMxlpQG7FhXPZUIzeHQmVKXA3je
e57UwXnWYP3GOYU/bwgjJRVKl3bVo0tpsm54oOTO46fGsZ7ZW1/i6e/YSndjnskz
9aaU1n3n3zlOJJZkvFmwblWgw9q6wNzMTYyGC6HFL7LmIR/95VDDvE4Tx1rOkuWH
g7Jx9BjDIU2j+ucWVAlYiISSKjGrfj0H1EMBejdXuO0zJOnTQqPhmR2DNqwKZZ6R
yZtjtei64hxExbjsmNySTsAQHrSwla3o0YFwqfha4qSTZE4By/SS0ppVu6rkZuDi
KZX8TRIQ4qo4v9/DVtBvCfB6d2Q+bC4VgCFl0RSt1YL4JX28tAZjOJI/n5RQ3CkS
cmUxZaznmLynarFMrP9HLtSppy6uHWrtpkpkPVWyo3fsaindSdaglby7sTUNYtAW
rvWKZjwRVc9cyqzQPQqd5XopFoEadjOycVY5voaShJDTnIl/fovGSg4QEoEhX/Gx
XvD5aDIIa7QV3hhkMouxQMhR8miT8ghg0BM10pkeFXVCUv+fUADN3rsSJKZs/Tri
p/H3w4sJBWU4oUhfVCVoMwLqnCNEsm/CtWU77U3UdRQBC0IV74em07lEXCPC4Vqc
/FG0t/ME5kGYlllcoeoPYLPZdXOP5FcK87eV6zcH7wzwFxbRQPHdsO3RHmdGH8Se
s4d25yGXfW5fyV2u2g+gjchIibK386AiuEc2UO0Oq00Ng7e69PFyhB2EnRpXXKUK
m4xOpUcLnQ1LRGg9bcYfhRBLE6xjo879UReOuoJxfyUMtaq85ehGTkMvS+CmlpmJ
E86K9vx8fEwBjE8ha/bPDaG6cga24I3QGqSCDTEZzg7rWFvSkBKuFMJfrOSVyDA6
TsfH0xwzeVKwxoKDLznquOPJOX2T3AKHVsJgfd5YeT3Xrtr7cR0TbDS/3ugrpdbH
mGL6Bkg784xWC98XtjZgjbdurLGXRNFvSzSpYQFWbhZk7SINGXl2Q3h07DrRReps
H3NA0UX/Ji6WgeIUPaviOsDW/rTesyZsNQdlIw2ywMmkFo6bb/Nyx/mO9/AmhpQu
V8cpNIRgzTuWJXWX6Gi7eZgbHwiDS3OexRjglmK8oi5KWzkPm/7UuNbpZ3He6VQl
f9bYMsJ2mxbJn1VtLiuA0VX/3eJ7uCMnVOPmBB0HWaDUsTTcPvUoJumO/Foy82Sc
DWumQU/G37HTGd0ru4MLsDPSWFzIi0nxjFCANzdXFaSZAmIv5f6UnQt0L0ujyuW6
2QWdz63q47BKjIzSPVj2hbOiwzIPnt+Zx/hYPEA9YtVdI96wb9LmCtpv4ULfKp/y
Tpy4lXx7n4F7q+Osv5yUzzd63wakfIikS7nDXG3QQmFtWP3GOvGfHg0TwI6bZgSZ
Wp9yxYD5uGB2ktypsEtwM1Idr94zVPCVi2W3RZoc2G9zbmKjYpH5y0sBwXQzm52t
w0kICnfQ6ecg4tl4WzGfTzp/S6YVeBME3S48OFwgc1HE7qhn4W3vEXU/rTIHh9qZ
Un4ChXSHQexIkKz7tm5F9huDbvurpm0BAsgfv9TRc/abYAu5s2PjhyHgs1yAp4C9
GxdtJ1P8SPKhHpMmjSbxMZfUDug/9OfZOQkN8Wcx/HO7YSMtODNWGqQFyWyMg0A8
GonyaejulTdcrmg5ep0OgSlnSm6oJYaFx2hSfi2eOf5C2FA0dKf3KOk0NEl3m64H
e0AvssqXlNnNbVcmmpFhtS8CK2IkLI2gxrOOCAo3gDN3U3HVp85m3lDPo1GTpk9o
zUVl5Jt1HJ7ShHpEG6id2xYw801unaAZ5MHgSIKgKYlEyIQnreIh6v/3JPVS+Cgi
pY/FhJsOEBLQcdsmX7eMMI9jaLfL/TzzAs280NHUd61rnz1OUrV9ArUlHGr+oRP9
aLsV6qyfjyZJ9leMmt1j+PS+NWkGRiskFuS6NPQn9A1xm8Omrxo7nA+KTFnPg1BU
4jXTXoge5kyw9+6e3z2eUOi+mWqzH9YfMr1+5OjncLvpUYIsuSkDAZZDj+Ir6yqn
4kMBsZ5XqYPd9XXQsifuivVqaq7NA3tL6YgiVn1qsUPvLUNBHXwqjjwcKPNXGFUU
lM/f1rMiRh8AngtDC/CReD3rfTcZ9VBS0CLTTb0pgEi7Say24e9Q5WHqVW6+lGHs
AQz44ZN3XCDiYAHgtFVpzJV2EK6cSOmuIWZNA8GBIuCGUlUOxPXSbL7oyfiKffXz
JaK0CTwLZt9ALAiLiUcDXbZ9JEZUcmZ3I7qTs8CKyyFI6WYTjSZSMmqqTN8hh8Hm
w5p7ADIq1I7A/ytyJbHB/P41DFUNizPhSSJU1XoT5E1CSfFe4yjw8gZsMHIbk8f1
htlxv0LRiGCVZ25QE7Y+WX72hWEXcYO1gqF0ffIp/4nMqeLTmLMa4YCU9Wf3kmOv
bTWTPsPlpK/FB76KkMDVAb62x5FM1Eyr6ZNQ1xIegwsgo1OBlxlesdZS26Fp4sED
P5Mv/a372icTGhYKRzze0YfvK4nWDLG62vO5cT4VfBO3SL95rcmHzV5lkmJHicej
9cnq6yDMFyV3AsBQbJXLFf9CvcizUGTmjkYrYdH5T+C0DDADBIbCWj3II/EZVOI7
gTTMvOwmwgAllE96IYm10eANTkosc0dg90NZNX931qtasWTA/GBt78ZyoVXONHJ0
cLzAfJpX34ovEOjXKBPw+aQa+TCGkXs8NyrBIgnqQ0uLQhR5MQ29O8XTl4JS1p6Y
KRi/maTGEteRcrL0ac0Ywi9ljkWGY2/GRccpAcWl0KdaUelF19Crm1FSAHk00bBP
Gm0MA+hM38jXOoUpwEfYC7kCd1ZkmAMIdAWdz3XyGAgdkh4RhY1apDED64tTZwia
0+FRzgO3eYLetMMEUBwviFJBTdOYVVqu/MiEVA0oTejjWbA0PGJx8DKfhYM3dzvE
bw9M8bIRlC2Tcyx4RVzFPosq+tPoTCntyv90X0k6YQpIQWsSKYM5Xyva2CtfdUVF
iSxK5F8/zdSE/pHfrln1GRQOu+qSLtSm71Dbsj5x5ipA+lAwmnROFxLGuQmGc//s
T+1N1+yPvh2z6l3ebegxKKW19uuv0JDCPJrm9BsWPXKyUdwQCXpv7NvOgsu2yOxT
4fre3DYwJcS7U9kfock2iALAKhRYYYXjDdOqKOMUg2tN3UgWUbRNXZgd81RXcJIi
4KY2xwy107QbanoFFC4yFkpqkZewvpjaSxFjR0DsuYS2IW36YTgV8Gn5MdkEy09Z
sZNDS60StoAM1Ve9H7SInwtXamIayIkUIrdf6iO187mlrYfldZ53ovh8FRHn3qfR
lrtexHLJTMPEaIUdCUxmDlfOTy7BHW+6lCzgyhoamoeo0PNUOhuy+w4WOw6fCyax
jVEVMRDcV2p/Eb51/Sp5ykkAxohdAZbeEiQS5bD1M4oHiT2ZoQRWkJDHKsXwrdok
SRimb6CIleZCu0ZLv4hg2wYFwSeiwEVBeZ93kx3KKqbblooe4EDta27n/WvPgyOk
mfzUldGf9ADaRV7OHBdd+FIjVeU0vHwkUr82NBCNwYCN5/zn1h1Gz8A8POtNHmYS
d0yPV/DH7hDzmR6uEpXYJexrQw77K/kzjS/9czVyLjdW/uxxgIZGKk8gF18gZuOy
1ZSU7Y/MlgBi8VLt0gx/MtnDOhPr+nHsgMRdhbVjgn9xrLqEh8uI275HHr1VBP6c
mXQpzyS1+4zoaSndOedRvDzkk2c5zouDcBorfuHDkKjyMgAVfHXlwpNoixp+8E9F
9JMQ4G/kDo1/cyk7m10tg1NGxjTiFJ66mv/QiDQkfsuabXl9ioWYnroG7MxvWp8/
w7jXwCPX9lohSojUQcThYr9i32HzOqgtQAdAdkWsxfvYpHGNM8EJ7PnnG2FEbrSh
bLjJZ9DKF61gqp34/jdiG2D++J/KmLCoYb+8Y+l6pMiGwv6Rpuwai0qkOhiAIGBS
H8F3m7UG4lAqEyWCDbhnSZVE2jFiVBX73nNzD4qb0KZc3bS9SvXppq5wJcLg03dr
QMhU2QspIqOo+QVbZyS0JEpDk9gI3d1WsA9euKt8DDDTwfltA/2ViE1nWsKiW2rE
oYQr+0hZlGKvN+ICKeNXKoFXNllpb926m2ZcxNqHb1b0sek108kpTrzvK9DGMK91
lcKcwU6fa9SteeiZ+zsge+AwCknL3XS5NcxLTNMfEobNfuJsOKvDMQzmjbEWLrZb
YHPRfIhIypsa62P1S80ngsHAhnJur5GOafOL1LcgiDEfJAhadTzZiuXgidkKdckp
4LPeuKjgRxmlMTQQCNGjUORFe6CEF/VpSy8zl45npYjujyM+mRvrcv9PCYIaBaSQ
HWkZqmvdl2x94RnJgdyBRmupcJws0StB50t1LyCeRLTlu9+Y83VNEgaW5FZkM+2U
QrZdDsphntK/A8cyvfSd7pTdhzIICxVghjyr5nVUVtQr3dVijaA6INxAvxNnbCdM
4YZ1Kkfz3CyRw4rqauXWAg3EyGj6nLkmqRveNCuGaMuU3MBDosg92mstEj2kaALc
4NJcNaaqqq4l3a6YjripEubX3weXA8ugM5EUI71lKBG7RkE7EqOaMOCxtTk8i707
c0zSuIsM8v0fGkmUIyhtA2GobBqA4BS/AsXX6xnn9troDazhMynXI3XhTWJOfiSm
5IYM8x//av7168ARzrn4C5SslKS8q6Px8p1voKyQBJwxTYIR9RGqeDzyBJjMLPVH
GdoYXRl9VVtrtGgzLzEhpFkM8ckg3cQ5erJAoi3Gi1YgHzFBvGsFRFsEhrayp6BV
cwmLvY0H331u1BdAYLSzHm4LZmr/z9GYG5qDIGcW2tQRUwqrl0FSh5NYrB2dVQui
hCDP9+NwXLnjPcybB1QtqSrCJjQe/T5azKwTtdsWtWOlscyzo380VRIIGBUE94W0
e5cARkoAn06JxL877HR/k9oPh6SYVs9INo7eZfn3+uJB5xrphoUTGnO6YEQcSZTc
RwaXWkKyCo4mGV52ZcKJ9A95FvI62FgOiS6iojOY3R0kkyrqxyTaUXdKAQxBzhed
12ZWdFYn85Z6ONqSUXRggilKApXc0TsCCF6KuyYxiTQgEtrd1TIsEwofOvr0WwjE
P6VZOcz9hMlbHnK8JrtlDmcriXxHaB/+z3QjAQvWvVi0Jx/5obFgDHvSh4kjqcBy
rNcSREQNE9pgxmvREDF980dI4do5albSOMYC7j/E0OvnnfgWLee7EX/ph4sE9y36
pkP+ZDT81fI9LYmuvCraj9pJNYAfqDxwh3ZptI3s4kK4y2aNWf4Znk1XhpLSLNg1
IKVNMrAKesYzG+pNLwYF9E/IT3qp556i+5PIrkfJ3ABGkfmLJPW+3xXhH2ryAZKX
03YMP+kXusuOchaSSTsG7zUycmfvFGqlxhKcre8lgVxECAejkmccyNyXJ7UP4Yvp
j48TtIaM2vuRJ7B4pzx4/ZEN250yL3ubnex9x0KApDcCDVWK7sUNELZHva3ju/Vu
8Qh89OXGSHlmt3kp4G42QJiP6Z1FDngv76C8mndj5S4Ay/p18aLJbgYluM3n9jAf
/QBZPZbZgOYaiyFVtizY6BKD0LN6PaOMLwEtcvUMVndSWNzdwvF0Uijks8X1/7XN
3C0uCTkwAcAIP/IoeueoNSRBd7eVeHggTIrux41Tbq7gbc4PP0l2ivMnUOdF4rwW
tw42ogMwKX2x7BgOnS6m70quPS+JyXENjcO3cVCtkAmu2wmwoYTZ+uGBBU04GXEO
URu2pys1eEhZ8f78YJ+emmxFMV9xC5zZ+LZQGVE9g4LC0ak3LFmb+IevA73UOi5i
2C+oKmlR8k1JV3V0LncEp/H+a+/i6Xpkr8IzaqjdYlJafVqJprWaKdhdkRgN1jtv
DK9RLOwgFHeF+MPgdeP2FgHpWfRQ9jdvVSpd2x7yhoB7z+kTLAT5nsY9xZnlfNmL
HvEKTgTBScwBRvsxWcxVyHRwOmIb0oYu2smOZUPeWVEwatrauY9TPLETttXtlYxU
YjWYkIiKMiHZfpRQmcAdWiSoHP8qgZ4xLgVW16Ks+14LGUj7EL21O5Q6NPKw5+xQ
AKBUBGdtPV1ls4/0PsEjVFUHEq9cUj9x94a5Huk+Db/VGHd3sSpd10NQ4iHnPeuD
tHJLgF2bFslFOP0xDtKDDxkfw6VCQnBYBw8m+a9loFshsK364rw6ZwVC0VdKGoE4
TMDusjPJhdB15iR//VywXuH+/qZZPpE7F8Avrfs1u2xSU0mrRagK8LRv+NIrhILK
fzMT9ov/17z271e1MP006EEMhOIirB70y5Rtjnkm5hRnDUMHCFBnj19C6DhkwqhT
qhL5xL9DifRR2EU1jdyJ2btKLX1yHXiqnCeLKia16Zb1mtzFHRZ477imtlX1vPWK
Dwt2C3olzionOE6mVufGyBu5ixnWRbzed7iAuast2/DCPUGQd6TVSeDDfgCsiU4U
W6qBMK5g7B1qqkZPSTmASPmJlrL2jE3VHm5niSHPMe4Q9aTFEaWZ0uI3Tq+Rgogb
NX8rNEqvJuvyVhX/CXdqCe6tWMkNQwdIgQgJVjVv4CRut+0i4aNqTxayskWY738S
rCT9NGUKxOVKwn4yQLx/MYC0D8jbCM9ewUeMRR4MxQxCUTl1aRwf1+UUtZfd15dR
YE6GcXTDMGc4ObYPF/wBlWFq1XweB2v6Dr+INzwr1kh/av9+JP/CRcwjpAxQvEeI
cgZSzNXIClCwlngbv2fS1NJoS/C9IYVz8oBo9PnVAqnB+qMa/Y1e9vMnJVNLYOg0
vnSnuSw455GItadcPmuQ2tZDzgYH9xr3ag32SS/PVaupYQjA/ee+Pfd/LwEqIBWP
TSW8lt1SwQOe4abFzRqU3HfRCD+N9N3de/Z3Dx/jTPTi8hpQalISPuCVU/zjwBU1
BnQ3w8X5fGkOdKoxCeHrhBqTeTh+Ok5dXeUxF3AUdROa97vkYMLdmEcBxYrFeKRh
pF64A99Pf2tW3i3mSLba9mmVGz3NXuzS6HbtBWEiMNkzz6WBucd4EHaekbC9UTjO
ATrZ0KjBpl0XJ7HeYMmfS+WkG//sl22h9cPJGw1ZUHlGRCxVhoLbqGKadqnaO/KW
3QgFZzNpZ32/Opyv2u/w7dbDlkfg6H3tMKqppPFH6xMip/yUteL/AfB1wUMKJ1Ao
9Zevzap2nG1M+7GM+k8GdZxCUuM8E9HGY3BIw6TOQOkpvELZWCQBQwhgwhAEzOFH
81mEblYApdAqYPdLHDJM9quMAnLL9d+5czQz5mWYZnA+ST2s8CZwWHn5szOMJmzG
sGyNAdRxLFqMK20GMg8WeLIKJQ8F9OinRO+akiVl/5FzekqaVM6/qlddRPvcNqcU
6AzYnzKdaYLNQmmSORHTCHMHLsgrjqWHK9Um95HnUlUqGQo9oxLjMGWY03wIDfoi
+TwX5sYn+M+ThmTglf+4DWrAZZ0TrVFgJAGLm+8yUmuHXuPJXMendp9MIsdsDnFN
4fDjmE082ujPfLDuxzItxvAOOwC7PmXXytU78ddZIt8SFjmZ0OlLgwOMAZ3svtKl
N5qTUgbmDKygWkdWT+X+jJq1msfvjx2DYDmaJcC6hfdWAuCYztabgjWJaOA+Zkqt
PftUivML0v7zcLARV5tvhdjYAb+r0RV1EWPfWYYu99etasP9MwcIjeYxJ7r0wDuy
DC02lVMV7W5ZkXFpU6yyK1vQvX7F0kB0h4tbQwXaj0w1fUSjTVTvNHFQ/OGqZ7nk
imz8wpRbTk0wqRdTfVJCf0D3EPqMryDHJJnlD9eOUyASQRY22Zm0mDmErOqqy5zS
1pdY37Y557I7h66c/o2VrZkPOSUD6zsxYsMaJAp9ZMYIvgNbl8eG/fmu34vRUk9e
yYEcK4/NiiPvF+WaEwRFssfEMucdjO1ztnSsneXXI9h+Mp+jO9WHYfCAWwCPN0w1
y/AjP3wvNBIdT8TgvEt6CC8qXT7XsHtzNCNZtg/49Xcemkzm61iAv61WtptHolkT
39lQY9lCQTA+YOXdSS5/ttXkI/k5hitBBLX2UjeC7a/seWyHj8cBd6IKV7Jc9qOj
zNTxOQABGXbryTdEvlOLTVDdYdi32cgADGK77p8l6qxC63zbItUbR286R6FdI8Og
B6sE3sAs0I7tgaP1egpodOkWc5BnpBxschgZ2RntPJUOXBmJGwD7FzY/9/ttDu9M
Zg1znqgWMw8lymIbzPffx48jyyFfroBMe0yZ6sOEyK/4BNa4HbXVD9For06fvmQb
SHWhWixQVQuXvNVrT1q3OfikR+efyQestfGrZ7zaH1c+33Z6Tq+a/fv4OzR+3enH
jsVwh6GNMsRf8dJGRSnsd0p3+1psUx5ONn4/1PrMj83+70RmTS1JEjE/M3io4xeS
YAfX1jgzU/kT1YGCYapqpmoO8l8gQSzV3nfWBGxP/vtsHV9p94nj6WfFGlpkvvSD
z2UkY7fSxo4EGwLMZi8gSm5KFIJZiY+rc3T5htfyAvi87La3a6JoeKPEGkxDpiMV
dRNkZS8j2GMDC/1JJ0EB36INWkaRDWV6grzGbrMBPKVLFbaaj7g6SZ1lhZ6tYS45
KEKF1U4dNLmSA4N4ILD0KvIs+hG8WXkp5iJvsyYYy19GAJGSm0G7KmtJA+PQ4s7S
NehaITzre8kBr7ieLRTi2soE6cwBo1tkZ3sj5lLIkRwpcN7/2gfHSwtZQmxBuHHt
KA99Npae/i681qhR6NhKtknesN3Lxi7BtQrMhDGq/6F19NqdMZ3NlGei/vCXpfCM
jqmyXNfsGXo8eU5n7SVQ1OYrNex1dtsButcbbzMkezjW/29ZhfjvmLzFQOSZAgMK
hW61sJJReaSza8+QEvt9Wz6+2DaKuNVIMWi+ZXDuNOlkWiszS1ctGkLPpTXAA9yv
KjiuxIIzx6NYdpQxURuSTWEY6Do5qGwN3MtwMFzSDx+W24Zfw0h73pVDjxvrzmXv
LHVJv0H8LblAFa+qfyH6lURdPMc0K6y7bfmaL5LDtGMpuu0dJQZRxyGrNCu9U3mt
KIb6+HTJDAx1hrOg63tcWmY/VJW6892NcmutGk4Rc+c5pqaVXXG5CkbzcOIGX7Sx
ol55hesJyIlxLtyn9JGwJW0wv2iaks1a6itlFUE2MhyvQ4UFMYufC1KCNXfI9b1E
OD5NxhV4Tygc1oEqQmIZBqA2AGZJBR599AbYVkhkHOiUzpTbd+DI9Ap7z2+Lagpc
JIF2AnMJtOkFlMlcqgYRai4nJGQ6q1MS+eK/0mHAc4GGFkxkH2sHXpfv6syclQ38
V2GPDntPxB0pbl7S9u43V67GTbzz16obiA1ibayiU02icA6lE1frjPu6BtofhXns
qK12vX15HEP8TFg+8g/uGQLioyTDvuJ6t9idE/0HGFd20VVxgEf08rVdQYBZ0nze
KtLnfC6/LZr1YNk27VGlwSMBfMPMzm/hC7PiIHGCDJuibE+rgxrfTu6dQUXMMQ1I
HVGjD4AbdsnOUWiJTVKxfA760zXsiMlKg8sUyuriJ9ragI/ET4DoWmgCISRGl+hV
ZZnnFcqgy7JmDuyq+tABHH5cnFRdv8ykZFQGNRX1C8Cy/iFEphr7aOF/8r7hb/rq
Rg0HcWXgDGNdkwfiWOv1GeeTdGp8evVZ6wQmaSuPJ2Pxa9a5/e3Yu5JM/SOk8Lpl
9kkbjMmJ4lQbS3O2n7hIjAHzVAxI0otgxhHyPniP3zZb6R1jpv64aZNvCk+Ou8AW
LhdUhWpQ/ML4odzcnPgiPslrSeYT8Uqk4cia+7T6Az6CFfm0uKxL3oBzAfz6GhPr
9bUKTHU2BNmxYsS5xlyufSj7blL+RcubsSDKm+Ai9NyKTdXDgCpPqW1Yz7oWzz57
YPkrM8yyg+xvV1ObAffIRW1YLR3TL9WH2/ADZix/Ri5d7LPFXUR+6WMg6Pl5ICgu
Bqd7bwsBONOGWAG/DaKnFGEJlwOAiFSSUGeDMX5EWQ7xrJghYUVc1JjAar7IyZed
6hiug7k9bpTDy89nkyqGtzyy637N5puBo6MiswsFYtRl+niaapld2L/kCruF5+/A
L7sa6BxjELss6v1tjDJJf1D+T+UEyQoozScCk80yxKnvN5VHVv9XuY6g7dGtlNCb
mpmrCWVbuyfSFYAgl1+aM94MfEluUu8PiVQegZQ8I6cnFYBL7w5jeMkZOMKUdZD5
UV1fPiJrrSAcgFtHIuWQdUS2Q8n5C12wh51OpQbOTne51MKU6W64ZT8yWDtUj0xN
USDZ3hXsp0gmOEm3/jG8oExT/ld9B5oJmOF87Ul3W+nqloMvcbB98GNgRMi9Rg4h
Jzbh+1CK1jbam2L8C+L8aj+v3oRydiDBeA9yzg8UKqV/2KzdhOajNuMXPukV5Qrr
X1Wdokpd2yzTFj25BhfPAFt3MNHADxilpZAE4PcJceauXnWQGZ+y91NWeNv9kIgF
7XpBgQdy1N464CrP9C9yGHp4H739QfL6A+NmiXX1u2bdhl9K/gAF495v4aqkvj+K
et1iGI1ukmuSjq0nUuOgrsfsTVOaffxyUkjNGAXinPhBXuVMsjExz0z0xtPuS6T1
TDlHOYVzO0ngVzjBzpPo8c6YaE2SSyzUy7UYGjIbsXpmho6K2pd+RFZz3FyZC1FR
szmLM6p0tAnmZPBSIwOQZdOtB5gHBq1z0C/ZJAScdtySd1cc8pLQpsvt6eTBTqL8
Bcy3pbNnPvANZoP4OeG+c9a3xRrvVv3uoqubhxmYUDa97MwzljiqFMjnVtRMnLBX
h9+UBfj977/Y1eLPbTO8KHaez1oUjfMDzgShYHJeIGlBBA9aO/ZNjgAnj7tMck6C
i2a+OsPH8Nlbi7jBNtKFp/qcCWyODJOL5nQj3cQL5l02y3+NiIHEMdWRNe88F0vM
4As32KMyCIiHNur63UJBCtF4/02s2ANjLojnqWzQlA3iaY9imF3Kts+t/a471xmo
NfHrEunwclzI1fA/rsXX+KkmHgd641mNo6RFKnWSYREE5OqtsNudmRmZCttfzxDW
tZjjNny76TNHf6H0ZG5azxcWQF5VBWqc2/VJv5dwd2MmMzBclva2vRwxPG0ZtvZQ
0BTloKva/NDtXP4UYsJnX+TKXiPpw4sE/p9B4a0+LFE4ogXkwxYk+dIcQ3dDiKlw
KyeT7bWtdXuRi0s67WNBHi7dGfDQzd0shFdsEP6IPlAW1w2QtJ8bRWLpq3Jif5p0
gPWVgfrxJgFX66VpOB/rzmoLWu+79CjMogCygFnuIRju6zc/egOOb/uCCBiBPVtc
U2NIfs+f3wixbB+D8K1T4YfKdFF9w2qMKk5kbDFtAlv+JBQihmAwcVzbBGk8d9LB
9aQHrzp1kjiJZUZt/Dd/K3wcHp4aSb3G5RFFiV+nSj+xXvOfaCXf1S/0r2DVgHmq
Tlhk1swwFb9/bNaQ20bXooBkgimdTB8EPDqEkSHznI53mHZgYgFQ6w2rVjfFO9Ku
AZsAnuQYGQOX+ZPSedbLj8w/I9423co1Tlg6DAO1V+jegtTp1tbnPgxiDaFKymsm
Q4ZSEYFmnkG2vP2zfun5fS32DlCpO79pP9aBwDDLvhWxpLNfv04/8iPC9gt25Al7
DoyktMdk8mPGw5LHuPWVij0Ht0vIeS1rk9nRIAdHO5SdvNxGO1Ag9j97hfOxG2j0
p93Jxw+mkeJwDXdSZ7D0v9Nxo8rlLnLS5BHJlNiRTewm0tjNTgAxQgtwT9wVoR1i
ln5wobgmNs8FiJdzx1Tmklt5OcDYh7ZRSEedJzTAbJvtrJBnfghxdqYkHxpa/zuP
FubQqu2vPL145TqPsEJiLh0T9BLHT8MiYoY6nK4Jv09sDY1Vdel7px8K36gIDN+q
AiGF7Le6R4kEIk15cJIwFpYAtxAle97JK7pFmA/0mfg+ndV2ClwmteLGmQ/pL9Lw
Uy+4wBkv4H47RFYx/Lyw5jYR8r97ZBvfAYEC358M9trzviWYv7myjQNVVH2oZqnf
Ql4bG41FuJYFnW8qGGUISdOFbZPFPOo0B9X9RAMFaWcPrWZJWknTQ9iZ5tC8oZI4
b7PwZxfCFXTWwkuvSq8o8WNhiU+xNdQBYZTxmM0KwuRD7E33cbBXlsIukEVNUEfm
7NgtHVCOjYx6ZhAN0MVxeIfT1hGG0xRrxCqJBT5lMKNtXqrTN6aaVNDtyvptACHG
9Cr2X2JmsWra5EaNJ2TTlvPeVDX1voE+rHkttwNur6t12QpexitCA5Gjr70YRnh9
UxexluCsHsOX4q7is7MLKYqRiQmrF+YatLZheHuUWfAbqO9n1V0H3uxv6aVciQIH
Y3ukji4rqPBDf1jE2eci3nSa9/7qpzOtRRvQVVsl5q1H9cu8T6GUtLCDlt4Q3QNG
e9dzR4ZL8K29IHGYbZ5W+/XaPpnPwIvzAL2uVitW2UJ4rI6M7MJLsngTqQGId0Ho
Nz7mSZ3P3T2HnW5duMOsioDke35SWlV8ocTvRt6s8cWH2o+aYHjLaJhs6cChDIf5
L0vgZn+Itet87jyTSXZeXlrmL/qHzOeBHQ972ZhoYE0xFFrchNMArBo/797xbZJD
MlMsAlGh5kSkH6RTYjC59kMbJ2qGkC0+WyJnuB/Yu8389OzuSCCjzwuZLVPALTKG
Mr5cPq2u1n1BmLnPzPu631lGMbepA6PRJxiAZhC9V1csK67PvlUwEkXtKaJpOsyQ
A+ePI3Ku2mlgt2f3kt+JjJeU2lCiPjJJ8921Dxqgo87nEnkjdZ7sSZPWMGj2yZza
sbRul2Kyfw5onv/wYLMHDYqhYxvxfM6kh9nGvCmWADVzwtTSGW+ccHmOG8lFZMc3
0Nh+hLJG8Q+wvJYlhtz/AT+kNt2DKFeaEu74Oq92MX9Bv52eVMapMTtDGW+HI4WP
5PQpk6jW0dr5llrUnwNJwrOkPztO0fCch+d5uZtsdy03TxFW5XoHy6bXjOZvJogE
RMxqOp5xGb7KXSnxSpl49XrkIxEO925siiQGp1ELqG+YDjUf8AbqnDPQYbM5MSzt
hmIaARB0PnEHUaB6o8HoCSjF5I4+b7h7ALv1lUu+IWNXMv0qgousdoWvv3jQuHDb
L9mdhx0fKepjGuh96XHhk8sijWWzPW5j4v47cj8kLDzmk9YPsKwprcfU66Nvslwt
RdCaXGAGUeJZ72c9qSpzY2OjBTydp3Hab0bEKO8o7YX+KeStY5kdeDWgLzDdSzrj
CJMP54s5RmqgzITIgddHj9HHjocV0nADo26CezdHKoQFn04/ciD4Bv2menpwOIZP
izr1ZKipT4G/SXPa+tPdwBOVBkstlskdtCG1dHoX5SpXplGmraewtJ8pmlqeWlo1
k8nZjQeXhn2FsFoBb1P5Z10RQLKQVAj4xwqdmOqAOp3/uNZ+emQMA8Ei0Uc4v3FC
hkbKq8n6+dER44jBIKsfFJ9n2KXFopDWIL3CXr+nX4Dz56dAi1pcr9qWD4YV20mq
AwTkr2ZRQ9f3+cBXdGluZ0WKXgngLBNPF/V2tmNmrC724v53aD3nHnu4Y7Xvj6Sk
6AV7/z+nr6bvPFw4DE8SvzkX1+LWYd8MAN80oSNPchsmZ1nFz6OXt6CsP6CR2qKw
sPzjMqiXySHMFk+ZIzmdkBVjPOGmMoZ5Tk6X446ofP8XKxsxesOJD0CS1l8QDBBb
KYdEuHuLw4RTWtJk5k1RQEoCdTMpO4mvd+StpuGPfGAvFb7wrJ/R3oTMxUaS2ie7
U7rFsFapy7c6dfVDZR2HnuJvWElqdkhzffErpeuTh4hxrxYztDSRHgDvywX27j1z
jyyXR50s0sxLmRg5e+pg/26+T8Z0WUTZjRlYaWDCNyJHknRWPOcQrzeE6TtXj/Nw
lpGjVGjRdsXNtRZOiKEh5296ZHH4ewoR8aBjlyDtEhTxGFPFvEnJ+3bPwyAYWD4c
OTMppOHXLLC1AiHqFIAUp1WlDNqRro2Y1kNA9Q5cp7IoDX3pKmdWSTMXX2s3nYak
5C9/5UEhQY0H/AxJZUeUfRAQu4gRtRU8wW7Gomvu4D9brstVJH0LLyxC2x1eA3IN
zq4GJo78xKCyTG59zGuM+KL+4r49JWnKNw5x2Ff0VAJyqBANJNlIZRwuTYwW9o2o
c4k+oeGMtAGn1a0X9AAVkmeWQbr6gxyh//7YyOyPNlr7jbQe0Hq3yrYGW1Zpi3Vk
JZI1VgQmmXyNe1gSATj0o6oYHMnbtoNUsj4Ugjg7ES7xT2X42EbpdrvktaRgPOOs
eTB0Bt2pepNYjAD7fC1CNQovAuYUtd7vHq4JflXUQyPUtKc0NQBCHhJjcQVd/7ZY
594WoOEb3fszGFDxDUkqgnfw7zlp0/D8lUEh7DbKI4oWD+uWY5EXecAegtNqlbtd
C5l2eWSlLStdwtUUQDX8MRZ/5a+CzFDe7OFruUCizsZ3CCKOhuG7wAT2trD9w1Ew
Kdu068wh08LOWUQzhZYx/oNyswH2A5jdhjw7E+klClI4ofHmPCs6jh93RYAGpkJ0
OXOtlmGZOqSzAFav7GJdBgiuBQhz+yJgZiEohEjkuo7Y09dsLhIG0ppnuhUSeAEc
MWBu18wXcry5kjCu8PIfKPg96g4REOMFvihiNyg7FB07wkrmfhUlUTzoZzcbE47H
CDMEyuIv078qxQmXMPQXZwdLuU9BfLrIyTBQWMMJFywIonKnMNHbiQykC6kBBFn4
miUggvskes4LpoL2AsVv9/Uq32LZfV1pE2cS6aAjD8mt6OclX1dxvlnr38h9vlBs
WYZ6u21x0EGEPFKl9K14Zbed+VJCFRZ4dyYDyDTX0cF2G9/EoclfLmgbHS+jKw3B
MfE+bOftQlCxsXQ+/MckU/fowikSsYNiGPhnu2yk0OGSd/R+FG4nY6kLSGZ9D1aK
KnwHrAkB+1ebi/a3KTf7zdf5gNIng5YFfHHfrVMCRHGH2bTDvNit5F3HQpMnbQHd
Fuy0hkxOPbKH/4mpoGzEfpy9I4dRAoZEAEnVaYP3Ghnl3se/J38+jfdc+7Dc065B
OPbczA1YS34LF00Ru+D7LyxI/3tWZrIHj4Arrv/fwHRT2rVo6ldQnxpBC4TNaE/c
oi1WG4Wm3sq76EMjOGlZ29vTj1XymLjugGkXPXBRN+CTJdVzIOFtDx3pncy7Gw+v
5h7A1FuX/X8i4ctN9f2PWL1n7YVmQAB/90O+41sNQpNjG/HST5RmT16X9XQn5QDZ
co8sRYmCEmWg/UHokedXitez10KVll41+UQhQAkK4Bydm1f+xj8m6sZBLAjKSBHR
l0BG9AW43nxJbG9OklyAe8f7Wa89983Nxy3/1OgJ9gwz76BTW69WDQwaXcgkgLdx
1e7cMY7pCFbC9xrKiLMPlUums8sHuQWsTroaeCKNlkIktvtecROKILAPsDGFd+5n
A+YSFqbMGq3+ioWBU607spAKg0QHz6n4hH1HQRY5f95U2WsOZQ9PyJMqrgSTvhXX
My1YO4qDkij7KG67Rtz6t5NhkFcKYsFuEdmQhEHNzbXHkmMnF8VxYQN+gLlMjVgU
uguqGUGBY+NKH7svzi3wnyquakP22SrVBXH4sFabGiKCNlnnfq4GophzJ4w2vLoi
BdrWSbiwvLuJJ7QyqqGrrCqeBfGZv4Y2HY9jfYhLuMHQCD62byfKJzgkSgP1VsSL
ApG4yttQCGZb5cTa9XP1u+xjR8ADw9jdK16O0NQnUtqHLQ6hKUCwcBbVqGJaGIcF
O+2GqRoVjgnumnIciEq+hdE/UsR8DOoXArfiBtpjJoniLslDiapZPAhkM/N6Qkt9
A6vsjTdRcJCsOon7qN9dGNLs3AefcKWK70ECO/M7dvS4uKwGuenuZw0+4Cga4jK8
bJJzzucmVFc93wgMy0ReVQNdGApVkmsrfqcKaaRyPohCublDmiK0w0qgzdJHo25d
5VjbYUXX7PJ8ISKW6bEgdLI8I7WUfEjRO07S/D0DDP2Ct6QPMWEgV2yOD64T2pah
i1HTJVp8+h7/LzlgBEP7IE1p62gyhDrtrz9f9IdEQnGpAi90JymtL3UgvzbCmyRl
vXvaQ7sOZ/fZO842a+KLPsqXW/KF4B7/FP1pLUtVETxTTNpMBm6kvgZ7IWwj1Gw0
aXRnywc2QyzF6svTPKIN45EhkUcmn/J2RzO2UTF8mApcsTG4EZF8tfLc1Nfc8gpz
0i75z+sEanXpn1qd+orizgv2+sDcvvzAlbBFiZ3kYpHMTcr+/q7MATNGTYv9v1MZ
AEJiLQjj4mXgSekwEdkdsinVHJ83gLZiRZ05W3hCdKE4ltWncmT0r92YDcrRHaNX
y27WRlQa7QByHAxdRj7DsXJrIozQzQ/1woAubANZhbDWKJ93JyZTsR0PdvEN1fmX
Gv6AVMBllbix/rCxiL4ZREESnkNYWjd5CUySSYKxLZNiliHxpm0rfsEwV9RZ0mFX
sd7DTsbzbKMURM+WRvi+9fSCC7RZt8tOMdMKmmH4/jPxSbO/di5IaYYi7tznlntA
9wwbilEzmz2r9mhtRG+62Lgd8KZNBC9NltutCr2lMJmWLf36Lo2po+TeKms1YZzz
UgcTxCqkL6Jchgjk4/kL2oUIqexINt+tVp2lKnJP2CS/N5RGw1S1avlmBmNq86gG
z/858BnR1dnEATrLYhjVYIdgGq1h8V2ZVmFkprrp7sEh0FYUZ4qtG5OQG/33WfKk
taz8EsliWk6nOctntV8BphemzyBgDGioNJRwdo7c5Wf9/YUB0+MIAomMZeOQWzur
wyFgjvGGf132dSKhL19TKSEU2rWiE2G36DizgSpD8F9C3hPeExIvDulxdYV++oak
GsshAEzg07yELjyLsCv8Ddf7rWyfZV+3yxxxs15/P6i6zZZVJdqBc/dYgFk+88zn
Io3MD+sozdRJCcn1ZRcxrvJECjbxGKYKtVhTL1iskwoqLyfOvv6eiGzyNRhclYrs
xhKVB/BuLg+RfXYev+Z7kTBZHQ1phcU7fg0i1plT05895dgDVNOf6ZvEsn7PSZmI
yDNvP/vFvgmjP7DA/ooKDtTdvkIcrvNzyJtvz1N1QlF7b/ZPa7j/k8iGy9TpGUCd
RU0rNcd05YErtR4geadRu85LqLmiU714lRTfs83uJqe7WO0modbdZbJaDg+4vfaB
Dex7idCLNs0l/sQXegtPA95AdAUXCCwTnR66Y5uGI876R5AyDLBxdY6i0DpNZOz6
juey58wKFhZm2u/nLWwyW6J8wE9r66TETGyRCJtxF9tlgAtUGT0WQG5cxjN7WLGd
kxR+tv4/VDRU+ybkKHdb2c15mAzMUCrG6GcGxewXORRlubGQyZzfDiFiP6FTDd94
uvpcX6GwiiGa+LVg0S2/iiuf6nLqtwknwHzdL5VLzNy2et+4dvBE9IobZjXUdzGU
eRX/7InOdyTehw9AzkDmgGZr0FkfI47KMnB7jJ4vA5VgJhs77mOCEzIp8ejSJ6KD
0COIsoKqXeTJXlRPg5LTEM0KtgJSbSrZRVG7666hGY1phKq31voV2Igg9ZmjYT92
/rWgAFpVssAuKHLGVI+xhyFxqMFhe1w5RAflO8bYCB2PG0NM3JDiITWYJHXBl4l+
+IwaPES3NvQHEESunKYgxDSFPE7CgvwAiVzzA52h51LJJTLQNHJlWaKwqjQCLTh7
LKEiWcbPKB6S2UFgfI6oLq4eGTBNRmpDDkZpN0o12Xd8hO3aI1DBANkwYeeWRu7P
SWTj5WhuYY1fKOC7eVnbfVWIS1dGEpTP9Lb4V9YePTagVOILT2peiaseRLoPVxYy
Q36/1Wr+oAGBsHSvFRQCkzCVtgUUc9SLzCA85gjz2/7BfUsPpubxamvd+N/ErqYF
Rs7Pks3YwHlHncBObFdLM+Qg21FshNucatPQsAYxu+Z2G74RNH3k2jUsgsnCCNFb
WGXbL/xvFTFZAPCAEe1WAvtlZcZbdWeE2JjDz99ggoQMulpvKUpB5x+N6qrlIcBS
ff6bpLLnUVPmZ+4h/HOxiNNd1QtvCD8Cmdk4INuTsz8MnirBgyxwzNNYnjH7q6iZ
o3HUJa4/OeJubk29eOyAbS1OUIXzhwBLOJK4talh7OrSvY2zDAritzKxr96sogII
LGDvl49JmYKCAmHRa3qHXksEOGDuTVssTWk9IfOrs2W0FoBQCy/ubWBHFy875Kiy
ihuOGWvXNr1V5Oo/q18hUtkGYnaNGi7UyweQEOIxasHA0WKquI+VsMopjYKCJXmL
jbxuEv48VRTbbW94D5yqujv62hXSkGy7iabpUWZKLmNk/dE8cK9pKNkR0m3wWeLv
NkGplScXb+gO2vstwHZX5tGxmR51uaKjFjWg+Q605X86fSTx/pN29RrCBqaq3fWe
N3KiFxfB8vAliMQ/rzeQUQqgPe/PcISpoFiPQ6QhTXsfZu/cD6KJxNiHFqhtzO6p
Niybj0Zj8ao4XoPgBzkIVjvq7aWY7odN99HGGQNdx8BJDm+ExQCA6eKTOcPawxUX
PiNc6WrFki5hbO7uiPv2+LvQ5QskfboO9ot4Ygf+koCj+STwyMk6lGubu+pCD2w/
jp9NhmDxSVnyNkIjhn+Hh1dMW0bWgbm0tNXqKQsnpXhvCO3O0sVMZHqVZj3WeQyP
0Xvo/9FqPBbLh8gyaS3XTNQTV7sPjTXxOKFvwNMZJB1+2Kss0K0uFctZJqEkP3Wu
mw/N8RWBZ6t/9C0fU/OKj46B3ItOa6zpvozSn9LrbKLhbAjCVuEfvrGBm47VyxNt
1HZ5xS1Rmuy6ynZh2mpjkiBQbPuamqXAP2rS+bhP9LQUz6wsmfr8rDDO506UHFjX
0+UzmvI9rKaSTjXMaJ1IAe8SDj/+f7PuJRlhM86usW6VGo+c6CUf9P+X0ofAk+ib
TMyE7yWSLvxX6sCmg+lFaGtRD/w8hOCvA9Yxpy5YdCM2K6rz3F6LxaKVjCA2VMD1
WrzKiQMK66rmUlAPF9i3KLdH58uc+pYWwQsioqyDMhyr2kUjTSZOkZ7UCTrAQD5C
0C5b5BDM7pWmTiFQ1KZWDYL/khVupKBPt0LYXVvt8OuJr+L9hmF5tc7/dDhNW1TU
XRc2OFbCW6ACMp1wPiONP3b/RkcecBWUSizd9DAwpu0IxihI3f7uBuCmddIyF9B9
yiW0k/6782Ks7ciemz9yOo0R+xPsgmmPX2bf+/Ehxlx4lY/ICdXjWpkpS6JVTy3m
ub6xKbC7dFityClusKVcwv9+e2ioJx4ow+p0/HYkEatn5z2jjwkJz8DwaYZU/O8q
VmeLulNGSYH0xeyMLDrahVU8yTMBqRFu97mSRcQjM+HVxURPO/M2cOys+KbNgRFb
WDpxjUj7cSsW/c4CCQDNoFHzybM6aqPsFtgOn+MpgvwcBVutlVoPBfw8inDRPNKZ
kXeEppzxBbfgi1VSFAeVhfHRSIGTgAfBnwcgkfZseTShVQPxVVfVINLB/0iK/tBX
VNks+BARcEzKvPh2xAYzAXVcAY79BVym6TBHFE9clHh8k7FQO22polaNtAc2+h7w
OZDyxsYzQTntqJnw5wRopFytAK7m4mw8EJKFPyQKVnpQFIuwzCsjk5OcgjoFAWUN
HBwqyc9RbMseqIhsY8CxhYvHNm5IRsTc0PBejoJBfoLoOjl1yvpIhKhTRiUjlX7/
SU9UdpKzQVgHr+S8GWuawL7Pf9F3wjvyAm9OBUTqB/DRrc/sG+L2HUXnoPQT/elG
DkxlFrMsdDyp61uyEY8IdiQsjZ3l633/prqG5HSU1iYvJw2lUAmFQ6x197D0Ek4v
FRRSuAjRzNcfhavHjidkRic90FJXNYZ4TzKK0ddfWYY5Z4RVn0YwE2yrXXmWxgH0
2n8HChwvFZ9OvY5fe2N/vtKZcFyFiMQ0su/ns1QA2tO2MuPt6ixLQ0ztkh+EdddJ
4nL1AuYc8shzl4y/HpDqZxuHLWDfFSLd1nZOQbTpryPS/LrbgqG40LiLOqMwdVQF
IhaqftiRyZ/IpBNGMNuFKsPVu0Rnk5w0KG8s13yauXnVOKQW7P4RXVM7VEQO7kNZ
9vm8IWflSDE8gOc4SOZnu75gfOlcjbngNbmlxxtofsYXHJN08Yv3Pk5Cm9z57qt6
x/uxhUHazQ1SZAca0cFJ9jShQJM8dk0cVRu6fKiInvH0u4BVaVRN4g2ClSDD9lb1
BtrELYbPP17S5eyvesLN4NSmegdOEoBWgcIsvWLjKTmQDh6lT04z6PCe2+ihIOj4
twX2RQN7uIU8zkZP4NRRNkvrFZNW49Fdn9BHKFbH6IM0hmjarU1sSe8KXOWD9sn5
pxgX4sFBt0Tdh3GOnMKbMP1Oicrg0sAoA9g9wn5T1lbE8MCXIHCUzR3Vl3HZ/ENV
7oxXn6VmsUO7oNe+wYwzEExitDFL/d8SnizO5gN4HZe5v8P/FQZA+pNF3tmlkbh6
4mG2aapaVXItsAf3I3+H9LVl8GBcQDUdy72t5KITNtd6NHQ8EMUNBMT433v0y+tr
sy2AP9VQuWJZ1V9fK7LWzmX/N+T9BZKo/J7wdOylGxYhySWpTUXz6D/XcWYfWVxo
TJM2LXxGDCE8mueN3t1aCnI4EKYeuDQDsOz/GRNVGqlVagOcKiM2ISTj1QGVst0p
FeHtDpFIa4EtYrXzKxWWbqBC+9rRx9ojMrIrF6dyZZEDLIHwDnOHhyuQMmT51KQ+
LrKDWtFI85Swz7zmdSIeEtPib3Cj9D+Vvdz4tEAYs7pVr55lxpz4G6AU7AwrkvK5
Q74mAaYcAd7g4TRZZ8KVG5cgnZOnytPHqJv3gjIoMha+AFtvz06jMYKYYa0+asvn
flPcXAs72pcC1AE1TNvBjt0e8nJOqXxniEA6A6hIfEVpKW2XWE21nrJ9V50BuVfm
sIvnJ8RCHaGAcFUVFsE+bMcM8o/4ZC7w4WfSpNWeedkSwWudih2fdxsJYnVsnTLT
Oq5HUJHqPcs9oLb/ohsYFa/ZbWjhvXRCeK9ryGGapQJ2K1z/qnTgp6m6efEsVMkS
kbCXLnH0ziNTMoSb75c31D8KHnlvQNPD/0+ccOKFjxzNEH6VHs9vCX7l8yQeosh3
dPCDdxcnxC0OOCygm5u5bekLeY8sBt6iCd7cvtnggX2duVYnEQfP/mfMH3wJZJfs
pBK8Ik4vSdbCNFVuQMBCLKFswyOKMbeT24JDMhdVMx7BjiXkWuNHJw7t+34odL7s
6zx5Tw+KM4e9lbLS7Ul410nWWJHB9LjcdmYbRNsVvsD692AvlBDDSU2eyUlfMdGe
nRD6aoXi090tjOpuErJkbI5gtkLrwJbS/aHAVzP43HAvYxMRENp/XJCk+G7sLw36
gFYO1OB6RkPN0RRSwCFi4AYKy71/0B/azovLcUPacSbTVNr0pDCk5IC0YlgoAz0w
JgjOVyeq3qAtXltjVk9B0hnjNVqotC6XwhJFjy5g4ni1wScAPtoqrKEtXZt9IRiG
RGGBBZh/odGO32gnYmXmeU/mZub/WHbRUnqMf0RyMXLSynwYvWOgsOCVjMvc0H+Y
k2Oy2iYbcUHcER+Qsh7KZza1gnChBq+WxfCFpPdhQvntx8RjWdHSaPC0xXBMNPt9
kUgHVNH7qqU5aHcMcSkVNizmIL9H56XQ0CBYn0WVuD8+Rgosk6+OAn97iOIEEMSX
DJni9ryy8SZOiYm80L4oJZ2JaE6gipDpPjQ64rY8AfROESCNChRcFNyyoCk4HrGT
lfHzgRwuH5T/a/xqrNepyBfAGU1raws0NxEaYg1RNxaDQu4e2+gMgiv+dNLow343
iGJIbQSbm8ppEsLhjphznZIHPdEARmX1Jj0Do4jO3Pd/icEuRgF+T453iQIk62Fl
YPdVbmLw2rdPlHkIbJq404aYhmzXuXuGqPB4lNN547D5RJ8YrTZnq+CBGoP6SEf7
Qs++J1+OzvzBx16pre7mX6SRRUTvUcxjtMMoj81kEoA/L8ZPJTeyq2rIaovmSqej
29DuvaM9IDVBChTT3RyPWwEILx8WSI6Zn85VHxG1c50OSab5VvY0Pgy6Uc8LYp95
hfT3mPilhVOCUl/rQp4OdSFmZpWjPuPvCF6aXDUNmPYQIiVm3fqnvimvg0H9/oJ8
kSrfrNn2YF8oe/ssWSJrxAJX3inBPZj7NRuafi8FE0Sr4+5ZDpi/WkQeGaMa1wTW
V+9RW7lQD2Q1mHpNKaeZcqW5xkr42BWI6eriL9PwUxDCKFPbMqu2vpCFw5mI2Ylx
xoBD6YeUYm2gxLLeZNw4tEm3ECc92R5ATopJwdUhcVN5rpp5rckWYaXA35UlW16A
qSdMiq/rPNi0wAUOiudbFjV6HgAkchmFoNtqeBG98ypWYlvjmlWmZov649vRxtaf
Nb8flttLGDUUCYpf+MWCBeiqMshdaCv6W3VF/9OBJp3d3e1Y9nOGP8G4Qpkd1p/+
gzuZFtFmpc78Wq3E6uPPA8y14phuKzLkn0B2icjWg0zK0wDPJTP5PgUErPBuMpDT
BlLZzc0lfQ3SOxNkxUR3Nn3s+3m/EeVrmB95z3bmOs71AapWfgvWSrqJmjr+uzbo
5pD8zgXp8WYKfqpZoRBA2KaQJAsdEjeqoyYC3zbe3eW8xLraokuc+xQRGrIW+8qs
K4C6dpFCvYlKMqiUshRlWVOPWfMFQs5AvM+jtuoybcZJ79OPjmFEi3v+doMTcE3V
uY75LRTUtPbuACovgnXnF9UB/I7bStYBvjhb6TDwGXYrYDBWQ0kw+ADELXgo6QdO
zifoaFuNvHZw55lBtvbBlSInP52tySwVepdZW6l2bWurJgm06cOPfTdl62z3Z+nu
VEpqoU/6vcUFIlBgXBlhwqHj8CQgGlILcAIcxAYxhqcPtUIae2lQqWHkt1I+mZvO
dLimutH7X6srF16sxoms5WlpeMnxFxSxUHRAQJcehSWshkN/cOQNC/sroARrqW47
hWgJ3BaUc6KksuSWZoVtvMTy+qXxj4X2jq3aw4EN3AjqoeVxwg7s8wwyP+qbRJ83
vSvD+ieVx7pdHtGVJ2LmCF3XouZL8NqfBPejdFHqyRSS4OKgaO1G9Idf1CIWfPLw
GJ29IYS6hmVrzd03n04U1rRyCX7mdKKDDPZjjnBaFR5Kqf3V7oarHIA2A8Gzpauc
cX2n5X3Frv55AxiKYCAOTIL4hppk90VhzQWbyEp+cqxs4bX/Qv/zsC72o+zNIGa4
Bi7G+feX0WO1G9H+FkSlk6LhWw4hDHMIBqR3UK26ciW4biATz+nmFwclOyGq/kKV
QMXtDLqcIxRnxeNdmijCx5JdQ6bM6w+mMA8upFY0l75tfuXbsnXMI+MX/pElhOZl
5GsEhACAFvPbr5XkBvn3M8smXoWy5sheSqm/kpx5ZoQyNG8pFfriw1My5RKQklTq
nQjXzphMcG7mMtZ80xg7lJKCkgTfsdzGJiM4hZfaYlbsjErrLFhP9vCaf/wgeA3g
v2ERDVhM1Lue3NeuApaLkP5aEwl0UT8XJoPq9NN9RiBLHu/tUZiaYrrGKatTlm7A
pMb2M/pDbcMsWbqUbOD5r1vTsCoLDf5hcn7tj7C4mGeDjitXnfG6gOw48x2pqmb5
/AbPQ0xZf5d7bWS/+BnqeaK/pGwGX502+AziHa1P7sX5p0y3oJ13XmRIg7k+tFbm
HK7ktaQKNqZPrl7bddNC+Fzl2p4QsQDKb3Od0cvUyyg0hiZKkjPk0BgZjVG9Eg1k
nf3gLdl7JJ2ri/RrRw1APR89aNF5groE2hHk5f2mLVmXk8dOZCIuJ18+vYhXbUah
7YUuzeMi9b+m9NcrgovZIA0ULavNToSVPQK4IvacxPAD2FeGFSCpdyQTgZg+ie4u
WImIVYzD7AR7ktP29eXB829ERvGqUNC8xVAOqqB4tNkZYi4spTYMYZ51XnOzg6Bc
JvYKL6ppAaByf/9gurhb952nJyryB6tsVFnZmSG+mYw38RDEt8zXGEX/USwLxPtv
p+zehKK0aF+q7QxWPUmC9h42AEShAHErOB6i9z8ougTjnHkg5SqTjwPpFa1MT4ig
1SBx61j8qbgQpq2vgs/5kr8FF/AhQRBjENr/O5y79RHrNI1S+FohxbAtCzQr+nO0
8cZG2f/Ag7AmjjvIdCZzJ8R3UUW6DgLf0m+3d6O4bBZzgAVlh/sqXermfW9P3Faz
M+kqciQt3Opd0kELD+7t3tgyRurTJ7urvUao9sB90eu5RoZn6QqtpPK6+i9zWwn/
sOD67gACjKuaQZYVsVv5JN65BhyFaPZCQaYnjM/vb4CK7+grcFGITHd3xsW2XAvZ
yz5tr9NvaIqk0YXwPV79K5eThkouq8IcpuTqQ6d3+WR0DsS4nk/14oSPveWn9q/x
GJiPpjLzeDKpLKvNGARHPqZu/jrNrknxwttDELflNuyOZ0YZ8D4hMPxjAQ7+djs6
UGgMWg534swQku0hj/Hm8+A8nE4f8IBGd2ow5ZEZ84D8pqqVpsgUUkmUgSrPP6Jf
xp33wuXX7FFAe4vg1sH2t31vl+lQV4p/53vYLpuxKDeuWAC/GIrHYcAmlKI8SyhQ
dmrJePeuIZQzMFVOoaohDeQYhqcG3phT8rfBbz99i3TYwCpFamBwGIbmTTXpg1qv
ZYI7onspxHuDDEdYWhL32Pt9ES2uHpM+1nA1UhIKhdNCLLmFA1YGCyJjiDBjM7Pv
oTCNzACShLN1pnnB+o48lOfrdw3GTGk/jrWPQ0/dQpJxMtrQA4jV+eL/5TQN4+4i
U1ry2qUJUQira0q1Z72gOvUNUcSQW9Tu5mE2Hmz+64SI5T7tGnzoXbBeBTebYFA1
LMtae3EA3pcVKuW99j2z/Y7QSw+hUDXCbqFw7UyDxenSBNkekBY7Gon6aTpDljI7
CeIYTMHKtc10RHnRrPQ24SkvdRalql1nE+O1K/k5DBLsBAhZ68RiAMvDtUKq0tZ8
Gizy4ZCUdsdwZKWzzBfXz8NzowFhgw+AS3b5wl+1IB4WvRpWqKPcI/0vyF6uMDBr
XDZRG5QAoCB7q7bgJrk6zaY/5r+TdQTv/tEvEP61W5Y7ydm/P4wKkP4o/SuVcUCh
WONnkhdTqmPoUycRiNwy104avS1+u9X0oM3yGjkqtwWGLhhN6/qrP+7b4fydO4OZ
gRfPZUPzam63CnMZ/MdH2KITmGad1Pd4DNztgAriXTmn9KjTxSrr5QTUClvMJRZl
0AtafW0BPzo5yZoFAmlDfM5uP0r6I89Bth4RcWerZ3RMMm7rtBwP675w5cu7IJiu
XGxC0cBVtn6nlZfaEErTM1CcgPnnJgBQq6GM5Qc2FjG6kIVJXM/pPvmQPRgZFTee
0vxvC+LgqXiyIZDWzeMZU32qfxPJmkPkSyit2tY1AJzNJmVmSZs7Wqf5X2St5Fz9
YT6slO6Zjw7jkVMVNlZ0lAS47RcPxpmrJZnlvOA9C94sAKK6VK/KS0GFzOarnj9E
sCoz06I2fY2ZspX3FZlwjAbG2RY27SI1z3XlNiuuHy+UbQakLH33PrPKVmuIxONO
3R45s+YiqQSANFDlVIIV/xjXvpunq6PicJWqBoQOZsgbuANeMbUHXlzIO2jlEBFy
JpwhQh3AgA1/U9nkndBUviVOzZlWXHCtpfO43LsXdR/N5ikktGfTSU52l7Gu25dx
VbpYHjvWJ8dcM2FckhP2WPSYyraX2Sb4eVVvxQY9g0e29eZfzqTykXrFnm57qYyu
8M9ui6GwUkmYNHXpya4B5ZefG4dNDWfcO9n3eu3cpqNxZP8X2IXUAw+Jw24Ua98j
1+E+5xKFudwArYfRxsGmTOvgO5GdjOvicXN17RhKPKh3CuHtle4l1SXCMac8VddL
+ypyUSW+KLB2r9OWTKBknFtS4RB31WFpOsFCryKzdK2r6NC7zljshLERQbQS5Q4m
0Roi6mgfNX2YcN7TD7SHJom/y1bZn3284xlsFn3BPCeDv9aAcIWPvVdz9naJasSa
jtU0ZY7YlNeQIQTVWYertK1IwgFidWl0X+lM1CF/xSUFYwOHGNEv6W5/xX5mkvnq
Jk76c6EqqOm2rG9HtyR5vITvgLP0CtFT3IWq78B+YdRP7qZF2lKulOgDhCi1GVLy
Sk0r9vrHNhs9tPDTpY9YQSktc1q17jRI+7uuP+qvmZ1zXq3oSnzrnmZR4XxNE+C5
C7sw7DA35dJ90CZ/hPCUdAD5O5+zQmR0N6+pKAWsSrS6x6JSJvxJSnKi2BhWRF9z
fdESonX5JNtDtCjmBQJFqhoxmcDPjxX/nKfrPz7cqNitxxR82gAZhxzixVSWDQ9K
D/BU6KA60qkNsZGcuEE9TxgaRGd2THpQgnennfzg6egUzyMiWntICoaZQI+NTBkr
R15g6km83ybUNBVPbPB6nkfv1Q8vErVtZSn8P9eq8lCBcVuJpwppk1c2zi94aLH+
QcHSkftERZB04wQtpVa/VV95Lne5A5WOVUyoOp+18qiuGcLIRFYqz/YCwGtfMnHj
k9Ppd8/A98L8YTQgsqlKT4z+AxBB6b/+Q6Y1XbsDtuwQuw7G7EJJzUOI91qIZK3n
gNVrJluJOmWdiqM40H7gL2AAzKOSRO+JFPcMqRzFVw90Zefr1MyfwGItdZZg4uK6
p3nfy6WFZILjiJAQNCKcJmzpX0kFGG8zS0mOqeMExtEV7Kil8Nd877ZfespXMQin
oJY/hrxoNrqhCOEza1iIIq/to03sQFb3VGtQOeRUg8lKtJb6AdpZI+oxvqZA6FLZ
GKl9LQLBXEvduInLKQoqWhtxQn1DHloXEbeR3s5oIGeriw098lZE2bftjkiBrOwy
xXC+cDOXsEllsKOQH3nrXGYRJGz/V7IuLuVUbYY+Du1sql84cbphOYpWOmmrHOo3
moIlO3OlktC3DwSZ6wzSwHwK76OWSVJCkbRyh/SwKPBRT4Bai0rBK5oHcGGpsbol
B9X9S9hy5Rgytv8hNdk++cZYezKHOhwkIMmLWG6ZKSyMRlb9PNZcMN8ue4zS1Ag8
FbiKRRKVOBTOI+lnizjiD60zm0oqFG9go7dokUXTOhxMGJ/mvol26s/eksij5dvN
rroPVSTx6vasz6CCbSfhFpLJE6pVbQtt8u3/Smsykj94HH1CMdORj7gRVpmnfM2x
ukAFzqZFS737nlSEH+oIsqv9GJjozFo2Gg9meJIjJXm/pUxYiyjxVGs1EF1bamR/
dGQoHjfqHhDHm6fBqjNGTnq/5E7R2EqzFtJT0/i0QteH+HIVUF+7xsZzE0P1wGnR
ZarZ0phKjqwRuV2+NET45g2UjRrgUX64RewxR5oO9gf8HP9viDgjVEX5YXKTZfHV
HptMPO/fAASLIeH4an33wuJK8FtPIdPNjJ290qztcImN7Or3YTETyYQlVn9mYyNi
KvzL6x7M0AFzMT21Azqco3e+VNezShvOwWjPl481SsQYRlsmPeDvBRMvLNzaxp0h
kAIAGJAn9nlRssVXT0v9mn5Lmsl4QbeqsX/J297lnt9a9eZYib6A4XItcVx/H13a
mRxvi6jsCx1eoaB+rRH5QVwQbETcULg+u022v9vXGGdr94IhpHcVhFzYiHQTxCk2
3XJ98qBkmUgn7cFECUtnMIVlCKqCX9/Rx/Js1zaz7zcKWDAPYp8rYcMpVvjDqA29
K7NHIxuxI3VlVMQ7pvdDBKYTRWxPAvMYSDBDrcnvDYQowcAZYdF4s8W6gIhzBp3z
f48y73FdHEd/aN8X6JVSsdFG2Ztsj3WmxbZuHkZAEIx7yL6DCRwgpQ8mqCopjiSl
TcUcLxn/S3osNTW4h6kOXfOo2b8t9mhcUDZ794cm/8nosxl+ju1oZMT/Csgqby+w
NWNRMkZg3UW+7ngspRzIe6kajcRDDzJAErDaK9SGgmZKY4t76wAf3Yv0xF7wypo5
Ar0ehp1YfAmbBXUclI9b4QZHmRNX0HQtQc3BugtoC51jXAd1ZKeFMQcZWUNeuibx
ryQdYFua7Hix5eC6uU8yzXLlL15tgpaj2jTpjUU8o1Iw5f0/6pckiMro0LJ1OEp2
OthrzCXezgCP3UYqwGPLkbnQL4xSNaUNAfsY57ly3peCiWDdoQSaGcDMARO0uKNk
w6USDIkBtqIzAtgwWkz2YjtN8G+NLR6HnVd4wKPTRoWCqK2L0OynWQYNRc2OOXvN
ZYN7qSX2gaP2mwOeNP2PkePajgnLqoNfHvDHc/FHbLGd9NdDI62jLAwSG0nTDYkk
E/BFVbSo+A+lQfS/OX8OWmEzJyabK0oA8Wn4rbRN/pA1jPwR2uaH1liQr2BX8LuP
rcWfl90D+KCjiviaUha7Bi4zdSDIA6R9GTMM+KlIwmncJ2poi33HZeCjRA82ucc1
/SEMji14SFJjGZBwkZ1F7sBRhzCf3TpZuzPwhCMaGO/92MEYaqQFeishw0+/pOjk
73ySjhLu9wUohny9Lg/ncXk4o8BDso+JuiEEbC+H1eerXx4/IWsLNsac275TQSw8
Zk8vsIuiqDmpcqlaTkzvAXffRDfOwvlC5K/pAOP2z2O4X17B6F5KFWyJ9Pr2lwZM
9OIKxED7s/WGvqwwppUvdQ52X90YLjbfUgxm08L4dZR0sgcVHk6OTSIE44qNZAMr
x9QZit9JPxIoZhPuYTLVQy3FVyzeju4+cJjv13E6V+Vr07KiOEFbOiyQersoPjAv
1bUBwmB8D+EiomVUVt2dJU1m/12GHB6fqNvAyKGi/thXRkVW9+V46pFHvx58jqnH
Dt/TWdV9UQCCZ+faGr4WzpVqTMbLgPYR1u2PSySLriFiYxzuRX80pv94/aHnOHQm
R6v4FKtuvEwXUnYDW64SLN8/od8fDkZtHhihjCItV2qT4Rns/i/4O0dbaQACG3/g
wkM3Z3e//ndd53hA/NoHwtF8J4F+N63i2shVNBVXiY57+NizMX6yybl1I80PvDNl
WkIyDp3wmOIpWvSzC9Z8Lu4lcFho5yXBvvi4are6ZtZCq+PfyDbxsck7eO+dzHqM
5T6bpJF0JwYJ5UaDHqpcIjKP4jfS8ydq/iGSToz9AhWRZW1oV1jhMhN/UE/PknXi
Hkq8vEEX2TeSquYlwymY8O/8dKmw8gxBudWw8GxtiF18Ftjfb4oYqk6dJ5x8EfUi
f2SSW/Pz3NcjAtkHvo/d+HSRO8sI++ifM9Io1YWtmvO6e4I0mjAgWeRAJw5aQyb4
kqR2RqO1XtONvrVWLQ+8HSlPOFkKRHRHAE706KclCpMgiiO/Rp5azCstnNcSMS9O
H2JHU1HJr58PjF0dD+U2MJ5IesQk9bSgPH7O4zvsVR/fa+50TCUKez2kwpBw9pXv
z6+1wDT5f1PwZHdgmYjbaN4d8pW2BqPqVf+d7fCgxfwYj0Ozbbx42nqiIKa/uXlX
73ldcIGYeQXM4qbNeX/peM7Sli+n/MS/kclKROvfKEl9dEcOGOMPxzv8oEhvYnei
vi9eu2R4LrvJ/TZC+84SlUurpMdkadxd7N+w/DgVyIO5gyVGRALh4OyQpsvuKen4
hfphOdUseY/qBqTlB/5hj9y+G24mI3m6MIrRA41MIv4bk2I+w5M8cienqbk/VyIl
ZZqKnQ2POkdH9w0ipWlk9L2yEph0L5VQQt44St+GAH3pFupIGi+U7gAjNBv9ybCO
HnqfHZsPdUUW0NJ6U2WVQ4RL9RZmt7FvPFYQ0nMnSI+W9vxdOKicfa1voOvRPl1A
ClW3wg0x81RcAIIz1vZBKXXTcMA8vj1uaXYbMhgFV7bSuAZdhnTlhN4zNmMcG0sr
X6TiNLAJltcQ3dD/65JksWOvmaPKHtn52yciX1BY0A/y5mcVvyFASfaGHHKVSvZX
fVPS3LCgRjzKteS7P/2WG2Hc1eghSGZvXOfy5Hgl5kPvP6NDAzxtakSHiA9vVf8f
5eb0RA+8z6H65B9Wx/16K22ANyx0x1gY1TkathmWO9w9dlsplgqaQC/Qe6UJdlbJ
RwsgcFP2iP+IQ3asBPKTKabgvsa1eXaHcjSahbDl8L90XxR99iPTgCrbaJok0qV+
aLJRyxcR263eFt8wn9ROZfmyKpx4s0HA+H9jRZUpzOCz2IRDGUn8tN1sUre43i5d
XnZooDZMJc0Mf6ML3YdABvk5TEN7F6AhM2iOW+OwnLgoU3qZd7gVVkkauOWO0aLI
In379V1XZf9mRfN+cfE/YOXc2pxts9DloWPRGCZVj9QHkWB2yHLl5Bh6MKVcO0f7
B3RAP0uTP2SfSQhih/eRIGUTqT19hArBFq5X+GoIVV3re0xo+WYravzCduzUAEir
P6JXRQZeNGTBmm5As/j0tAohsp3s9dhZeraiQyqfA0oZ37dyydp6gfKy6mFk9yA1
MTlQ2o32olbqPX5vLRRLa5gGt56wgtwLucTI4DSifSCknD8TwXzSsGujBq8si+zn
Jc+uYkha72GpMzic9cma7uKX9nw3vZ/EPnC0NHqrT5f2OUlPdWcTghllGg1xwlEp
jvpxUfrcPdx9peO/ej3aHeS4rLHIOw4zjgmKm2o1MY9zWkz1hzPtU6Zj24O9bKZg
IWFE4WdLWuVu4YFijq0tC/oPNiTnLxh6oSEC3ObostxrIqCkWZWa5EbUFk3rF0AW
GkFz2KT+/32tq79Y8uPLTvrm2MIhwmIKjesO9Y4YgDwP5fDh3Km0evtEKLF12M5C
f8ziGYI5ibsxkkDRCpeoVt+mtzC0qUTsfgRIIIQ54bR9XtGr7MOBJ6DHhBk/4xJq
jnrKD39+pdRJPFrIKgxsk4RGUPKwf0Q9mZah00xhVoIix1dxiJ2EI/x1+q4bt2IC
VibTG9CyozNTbFhNybIL49OA6KSZe6maG1D/C7BZADjFMXZqCbuRTRPYLxsWtL7h
MLl0ZJ4gZQgf8VG/xsJsYCZ2JtCJO2UtBAFmYFZOE3pR49PZq/R3EOXrpQswzQmP
5nhqFSiKWAnll+/Dc7kmNoZPIUh42ZP+EwsnuaGOtVLuUPqVIOvAsUIAo6Nz0wdK
lZaKXgPIIIpabFYC1H6M3H+mkO/MPWEKAsX+ws81hFSsa19HNgH+LUwVSRpaiU6Y
lW4Z/RavpIjA3Xpl7BIRcZix1otcA/wWMkEk8sBTLcsBdZZ9g8hJUrG8mc6XQyzD
h7LZfAdn0pg6vK3CdW6I1Qcz/Vq8rGUW7rTC9RB7y3W4esVjBvVVIdOV19+WhsVq
cDSnagSQkHHDT5YgxRfacdL/SCrCBXqkYwo65+xJiG3hvO6Cb9wOLaOwJNgIicf4
qbrJbVAMAfSK8zFzP8GCX2lOdpTr42VFW6GdqR1isKJSU+2hoeG5Di7+cUB6R48r
gtj4LKmWH4sDDhjE6+tGrNpCxHW/cKods+cCikFCe3j+3ElWTkaVCJRZ59w9ZRbe
qwl6vCjjj6kj0yEjknK3HbVjcSaVY1Cj16Bz8rXGQI5s2zQ1fkGqU1ug/wdMg1VM
Bi68sdu4xJcQPALkHwwd7VBtKo/7AoZzyAnToKYtxczpB4e+3/4LtyCQm/VU7M/a
iuJw5YMr4vMM1tLZbF2Ji9+q4mKb4sNPDjW5dDqKgUuxZwlBkcQF7e9G5WBIgx2d
ao9qs07kcUylZ2vb7x/vamVER1W0qvwcHjXLcJwBSPDOCxjPwakbC8RkhECBRHIx
AVrxG2o8m0/7PJ00NEORBqbGqEopfwoB3PhFKgRX0W/i2EIAoHVD8yENqUpIrNur
k1hKSqTy+/Zxi12Z3zg86KmGiyg1ScpFWVpj4UthbYK2b6Ygl2AtQusbWcuc1Nlk
nUCZPcQhrKDaH2V82iGeaG0UyYHwy+HOmiNPY+58Q5KSYQR1ZO0442INQYGYDkNn
+uUZRpqPSbLz+O1IAhobxmW7SWEArK11omOD/UnqzTRyPjjyE2zAWx8/SzrN08NC
qsL5F2bv3U9LCVAM+N703tu2WVUMcfxFZFsP+h4tvS1wOH/iGVmeSQhf0XubaWpv
PTNSsbRChWR4VCGvMlAndTYhP+zyG4X9v7ic4xCX8Ry8ycWl4PrGtecxzy5gC3cS
cHcQrI4W6ROO8NHExNOIwrrgEEsBOmsUyzGRuMdu9Xqs5FZVVSak347sh1UisU4U
pT//cjIyBsI7BAEl8axldI/Vzt3nv/+6m/lS/RaBs4WYQnqonY591EpB9mkZFcg1
uQiP6llfUi5WUdqZkyBvFTm7VQdW0birRsoks2OrNk5uZf7ibjfX1USoTgTay8BX
dMXDRBU4oVqEw0ShnOPwbySoTxW8YT/gYspXmGcxJrT5eFg7CX9m//Pzw+nEIyJh
HiN7H0UcK4qjl6L8NkOqQ7aiJQaOaMQb9usIVfmWJ0mXBGv7Zk7iai58rRC5fPUJ
R0zlBFDKqRQMo6oqkaG6vWOFbd7vXRQPib08DpOWSvzPF1LKGweF6+z8c+n70bvk
FzodvnHoLwW9Ag+7K3DRDQLmsl3p/gV3FFXHA/gJKbz7SVR+7dZpxD8vQ5nUV7mZ
zavdaqIVRdto+wkANTJ60HvBsPKGgF0xA7MK8dHlV+RQw/oX5ZK/UFjfWTuamhQU
lqDfe0d4zQUien65nx2k8B7oVfDUpY7ysh8Vfd184eG29n+YExS+pR2z5/3e0c6J
qf6r9Mw3Pw89hYME1IuEKrkaTpgTqKLQ9rQMJp2DPs4L5DmRU0T7ibO8aR79rkrJ
a9ER56oQOj9Qr+2sBlgy96SOqGItCLTergRVKwQGkZboaX8BtJUy/6d396xpIUZ6
Ne2+cDOkVZQb/cqjj48DxfuyYynE+sgkKhZnwyVpEKY4vbSBE/Lvp8wYjtvLm1eY
42g42oi3IvaOZNVRxPM7LvuJ6/e4zfFpZonUJFwbCO/zyifBUa+i/nppkhbspxQY
oMIQ56OxYMw7WzzsyzKtPqlLzhniIc5FlT/avilHnG6DZZYfOubcyiBAHD9verup
QZn+IQqwfjPaGd+4JiRm+CKVirIXtckBJnupYPYNnNv3mFFQDhwqlptavnBrD7q0
/K8KCdb4eoue4Is6yqsGZt1LsbiaHxE1Z3Yi8g2C7aBTPH6MUCpXQZ8UCVHBW9sB
n9EpXDADoz6xHw8PeNYjTHGfOzmyM10y5Mr6Ej3yQg1dziwaGABneBxzkk/xhC/y
X2XolfY7wS+suqI5NsMx7h9uW8MKz+LRe2AirsoHffPgpvIiSRVzwqkJGDLwhW2c
KTu0g0M9PuH/Af5Paaiaa6QUSU07RewHMe5y6lhG8y/6plqwL8kfNh8nrIZFchJP
7MY79vthhV6TwyA3jXzlCvLzu1AFIiHlKUTGxuwHHbtbLQT6uD0XbICzsRT6jNdS
gUowHBKVTNTU0mrshMh+Fed2Q1gnYQIEnO3V5ZbB80/xhtE4G8DlvGJ4ObkAgOI8
Lk2UUG1oD2ZRe3sjiyj/QAEQP4EVUHUTI3v3VOnghdYqIkehwnoHZHDAadRenzty
sQww/cd4qcH8MKgOlLW3ueimiDmaa8M9G0x6wTJIzJfG7l8EKxOQqxCnyYL400fT
ai30Eyjz0rKmLaSTgOIOGGv1ez+AiWKEtErt773Fbl31wdfMvG7zDI9zx42XujIR
SUV3ZxKiq9f0mvRERC6tyQoMnUooeFcDi7o9jQ27hTHxU3Uyw9KmKcTkMGesglwD
nIs87ysMs43RgPg4l5MfqYPiqAutSUMtxa3jk1XiXsWJ/b8btXwsmt9tfpU/Z68Y
lgO/ocMdpm76LrVNzC7265cUPXfhabysUBwuaq9JqFw7tHbhLHo9ZL42+JyihYQs
wQE4Lq2Ex34c8om3sohXD4Fw5pDjqhSUOZNirX3bW3PTDwP7moIKYWq6hmulllHV
VllUJX+Jsa6Xs37DVXQtq/SU2/Fys9GDRLDoLkW/FbQveY1WlxxQ5L9ullq1Wxm4
eysn3E+WleVljPo9eC46iDjj+pq/NnVG2GiPgTlCJ8XxlTF0dskeLqMN9u1xF6M5
2PB9IVDWNaNOOwwcRglAJ7QrK606xOVnoTXeQbYVnR/0XpUie/Zitxe2pZAzK6CU
+1E7K5zLu8iibqA/9gYznHT1ENYngeVyuLDh1CDMUvueb4QMrmiTa1+HcONJnqe0
/N161+qkXnpOUP5ut0sCiUnZTsoRR7BlpAjF9zWfAAZh0zUH8dwd8KAQxZjW7Y8P
fEVbDNjjcrCmvePPj9wGd7J+YkqSPF1aLyoRbBe7U9/Qwcs1eGjUz4kxaQkMqIxo
AscxxtH+pkcxp6xsbp19a1Db7C/EB+vJxWVQuXX8kaUC0OA2yw47SFHY/cXLpe49
xlt3BlQH3kz8LUNW5I8YO8FSwD/0pqDhx3/gpzzw0wUK5pmupcT3E2Ipe9cYgGmN
ef9TTgFEVISW5+yY4Q/XEVeIXWwrw9mWdGtPt6l1iDMHUtQXlc9NUkFvi4kxYiak
NutzuMar9bPixdHbsXvQtLMB2Xam+YBWLYB4rYimtI6aH9iVaQtFanBtVFlzbg37
YQ+2Xngh/SGfWKhyIeXoH5BWF7OvQ1FW5XrLlwUwNkIVsWJqgUQI4vT7hC7qk507
h4nU5Coalh5G9GPQ+i1OSC2E0+jAsLT+NPCOI3F3LLT4vkg3REN9PhTP5v8eMsh7
9bSRKiVoiNThidQVB9PIXNnNNHrrdh0GnFEakfWk5vR0xP1LyOj3GC/cbNoQvSmR
uGWkw7kmej6vEnkMUOrkLaOKC61aA8kTNaMjRpyEwXKXSUHvZ8zTIhgXEwPqvyYH
Q35BmKQ3i5mNvUCUwAVmg1l0ueGv5IxtdZyRRVVJYQ5ui3Mi8LvyFzmSDBivkvXy
bLHsW00Z8EKqpdbASKYfqr/j5bP8Awb+IRxqyRhSGGUfb1sB1hYgZsQXV+nWLu+k
Yo7iXL9hR5pm9PiFWRM1ZzNrK/EYVUhLkqQ4qGZ9BpEDOljALGI7rXIj3Njx7LEt
ZvwKwAypCvt32CMkpjSd5YcDAOesJfsP4zWn1YepBCJ9iRxNi1aMIUQXZiUUjel2
uG3Zp7SSENLIgnNsz8Yg9vWuKGIyE0qqMsx0nF5a4FcpCi/jR4FyxI7ULIjoTkiV
8cn9uyHqQZLBz0vA/9qAgRGPiM1DBc6Ol8+uYnM1TNqJfrFZm5vjPZtO4GemYjl8
0oXbKyPo3n2OrBDfmHkmm0u/qI8K+tNyhDZwJ+fuSsrj58t1cPOmKM7Ofh0YeQdc
ubO9F5cEVFryST3qHJEufOvnQYn88U/2mk60vzclpGv3rgRdcJsBIuUgBkmqc5QD
l3K2esqLGGFBRj9zqD3lpeyn0hOO3G9HHno9bBww2+Yz0GNh6zz/lYV71WBK6GSU
slK3qQsY1riQ0j9lKHc9GzuDZyUBf7DtvFkhHIdOAYrbioiM69OHNnJI5T+qmVy3
Pa42ug9Sk4uFMpcZvfUjAngjbhaHjWfM800eAR/f9cptcM7Wv+wdF8ay5D8pbmnG
JAgmYPWAUK/HRlqz44Zfsndo+MwO7zYvgQHDg8h+vJo9inpA+O0WAKzve+nCxGGL
csTGut64YB/TtxhRX/F1wNibsxLKxnzlQVSKFEQvY3CY5/iVsiWZHEEyrWslbyyC
tSjWNnJKEJixFuJtMxgPJO+/aBNX6WHpwYuNhp3GqIzCDjKdZwImmQhP3jbSvvth
jlSNkKgBClUs9aQnQwP0eIIEE6ZcA56JRYqqDU11muv3y/CnR+hWifRByzxp1bwm
mr2PK+D9+ZJdM8hOqqeiQEH4NkiR34eu6w6VUyMvFQN0/VC4YOsMhdWAhvnjguro
xitTq/gCmtusyZqjAU1xYxLcouJLUjJVzohfiBMRdoqA7VTMXWOBAGi5Fqv2Anb+
AQWL6Srjsl/heIpvu9e482aK5EljjxKe6JDPt3tCjTSPU9zecNMly2IdfhH0lZ/c
qf3r4/CYd5kRPOFZ/Kk4vg+H8ErK6O8KEk3o4YOyt73WXdHfvEYJrUCbbL5Hk9BG
AaMw27Hb9mb9mwGtOMobQR9k+vp/OueNuZd0hNIlQdgUa0J6WHIkvoJe75fy4Pax
5hL6lh0GpGGyay6LNVbgkNOcGeQe8E2s5NjvItE8zezE5+0dt+Ld90qLSKIrj0jV
YDs+OOOSL3bN5P9GIcpr/WfQSHzgMy5YxLkslcYTkS0sUeCgKeFWjw1BaQ4wvfMv
X8FTukjK0H+d0DO/YmuOZ55wjjJ/g3JqdQIMgNgvBxTJtydA1A6xLxlxq5VXfz/L
878FbPErl4+H4RrfJqrSjWOvryuWXgG8r7GsCi8lJSzzkEt5To3ihIy5JnVNN4u0
yJZfonsVEVURPbkBxxBqHe8BgSoTpQ7OqC4uD+O7ywFDQLxldYDQVUkeJIWN6Slq
C/dv12Q+PeVoyE0t2Y0LidxpINHB3n1TA5+HAl26PkJDyPebhCMSr1bSV5IvDX12
DyioTsWImti3JYqrr7qF8gDoMebt242iLMoGZytw5T8WWnieyZ7UiMyNO5JCIdj/
Rt7Gn1SgzUxXf/ufwjrpS9n58D+eCzXaqiQh0Kqzg2odWzQX3Ak91msQW6b74lWb
6XZYWqlnL3wNhPuXVR8w5yhq3xb7vcwW0FXMMdmVQaS36ysm/3sS38Q4aCkPS0Hi
7qoeI46WLikfNnaLe8HOh7pJJkXTLfzdHnM9DmrqhzJWo4Pbb4D8N3Pawd1oYy2P
zEiZ3J7WI3uJAh4gdOwu/ZE5UKbClSPdaQFSPUD615Cb5c3VpF89vTB3BZgvf2Ko
APgMm4X+WD59TP/ZxFYub1EIj6Mr64i3qhB/1cQ8moYNskgN1MOLyP+wuIUTYGrk
DVuPhUHx1Ye3fszl+ztAElrsPcamfpIGva7WSaszSF1ASU6CNf+YbgzfCBOHEIqW
IkXf1dhE9fs+47/M331hSp6RQBo6JkahNdYW/8sQszvwcktqu50/WHw50PNDC7uq
r7iniMJwnRtOgKLMglUTj/j6wdQ4NY1+2GpV5V3RgGfMcp+BPrD8CsBcKxCELrPX
VLXqAG+VUPuuSUyduP+PicZYfs909hjqvaULrSK41B49PVIx4UdljdyB15iZHMio
AB2eXHwN9HYCWUxhBzx5gHD1VgdfPhKvInizLxrkusTAowuFEeC6hthBQl9+a94i
DbJ/smX/uFBK6oblleE/CTrFWmALuvr16IVGTPpZBUl4J0LSo3rqUXDBVXkj2Uxg
Q23Q9i91bU7WQ80aGqP2pDWVdXrsQVVrkCDzXPASjO2qYLumejmvzz+AtA6mYaKy
uitlQzSbl+WlV/jdZLS8CKz60t+wj0bULd+Le4AX4VX1jt2P9V3/cf1qAHMnG2gs
+LuV8ukHNjVwhbBHRTm4MJTATdsTVY3S/e34cdgpMgMIzKkT570OQL0l3ZHBaaAb
RL34dxweUykaekZHBeM9dt81ftSsddJrdMWxfne6Luuvb7jqT3CJtH8g+a7r6hal
Lg28MQaXNFd3sLHXLLRCfLEV+NHrwdTJM0jD16Ih61cO/zjoNnaEtzrT3k8rjRto
P3o1DvYfWMCfzlWU3ufYX1AeTbmvEiTZ8eWeaw3AJk4UaeGqkW6Nkgh2NKfvSlAv
FlYgp0mRm6HC42tyMw63s6hM4LCjOA+OjkEW8aZ1HcJ6H6/jB448Tffo+zTC26RB
16GjXYlH6q4TtjRqEiQsdTCIWX2qm15CFDEIEK3+rAJ44J5C/kdET3dJDSD8Vob/
p7iy+J2StUR2N4blYTTsHXDg9sjezC8yWHXEr1lfDRK/IPrWvS2ZsZ+XZ6dMOnVT
c6SciyJvWxlG70k4rLEv1uTJJ8mSSua2JtcJArFQs7igDrX9OTg8pEoWrTDQ5Rqb
33ryvPphhJrsexjbblsgV8bnDilydTtQI375b6CA0jZy7/x6KO7qgZjBF8Rps0mO
RH9zxri8alyiRnjG7Gz13ULOCO2JFDSj72iNQVFcf6ZB/DlHOMS93YgBbyuMj//e
c2OuETcu83NrIsZ9FcLKPz8gN0j9ELMwA28YbGmPpN08zvhuxDaxIqPqpzlQAoCn
LtcGkUWQHFNfsjA7ybSLgNPfCaq28LQLBDms2NwgghvSxZS2DstrBsb8M/oy9crS
rgnV4fjX8FrR+kVIIzcsInJOq1ml8ddCgcTyWV6sLURgx27uYq4Wr3Ibrseyl0vl
H3GaHwPx+FRdJK3KT+IYnOrevIi5ClPW7YyTpTK7kq0jwI4K+rQvqxcGhNhrguz6
cwiDBCB7Xtaz5uUg3M3GCz6bCfFz0iWMNgJ9O570r6zJ7BgPcpWujkwF6w6Aniry
NXTQUdVhFRvuD5snluXrz/i0qWZrs3pzEiNyZJsN6XPuDY631uBh7IKcU/Sd0kuv
jvz1Qw4/sRYTCcrxSK4RcsnD9Fi+jHoVCQ77hARSZjJgKMY+gVen/DZBZtEBAlsZ
sElOFSgrWr2P1DNS/2ZNxy4Yk4/QiXlrqU3vofYkp8j0+F6fLcmlll1ZdMetllgn
WYrxixPemJiw/hWkH0HHcyDQkM4ck4iiHxtBXULUTtfK9z6f21cinkw40qZ1TScD
lUXVPP9oGl95WZPGbgyX+0ZYOlR2gN49Ibh3r6kFfmYps6h+CUTq4P97Ycjf1VFm
Y9J8tQSzLO6LKi18rdx2ryTzRTic5o562aRzWGvmIRYGP0a3/Dno1MtsSmPFlZMF
qjKcpsQNgXnEXlE70KrIWtHYhby/+AXFDpUBBEzvOO931IQ9P71J2IVshTHPpiwQ
cPMXEfVk7v+NKouqEUdzKYiaIrOQRIHvfMyUQvazZRqVkv0+1bXxkP4ecvyRjUYe
NIpZMTxzpvoAYUkmQhc1z1lbexy4zAf+6V5d3RCGJEPntah+nA+0erF/S7plftXI
I9jEvZYVNgKrqzspN+Ypb9q5YGh3tK9cDQ7NAn/OUAN3UtkKErZnFmbVYCZZsMhj
QWWzhP2w6Uyv3Aam/UsjJWZaxdzzAbQePuTNJGjlSqVqq4aFU9BvfBeNcFfATae2
q7qvsyxAc+Cg3C/5p8e38oxk8Bkg6NKq5P8RjCGwEuqo8OAYkXEbTuQj4eFP1UEO
TkfMRX7oFbTXlla9LqDyjqVt1d/rPltbeq6RvNs+q+PnNUih3vvcCX+lUxJbkcsd
Y6d5ew0aXf9j2XFLzmXhwMFzf8+5lZ0MTRJdhpeV6NkfW+aXpoXX1cHMqNDH90WQ
SeyiLkMj5YkT+IlZmbPDszAvs2O92hRQ7LZQj+/mwH1t1mNQrLiAUs3lAN87ZjGr
j5/qbyBYQ+Iopkfg+3ygRf37g7ZhWcCQ7ePZfgPSjRR/Lzh+EWbu/0LPDhvjHUgZ
IWMd2bink7FYwnLC1LTzpYOTaGDU4JLtrL04LyKSRg33DtXrrH6LmbtnjunMkUxf
RdH0sTM9Id0J4X3H5Tj1ej/SJO77KyIXmZOr3etyQJCqrkZr56STmpD9jUu255Wl
/MpXUx8sBTjKBjOuWIFude53oRhm5tqV0HRWBspR9bIn/UTy7J+DIX4QMHsMoTnk
r8utKrcyScM8JylpTPnGOXlL53BzuL8BEmT+C8JV3y2eapD5A+0mVuPHt0PZzRvE
OFcDDZRBWFRVjqUxAaERegClRW9/CmY/KmR+WVGRcIZF2yVWLcoI/lFHixHsMrYL
cEcBNJA5bRc8FRQjgQYmE4J13lRV/RAsv9Fd/jGO1wv3067w3CGuJtLlhMajixso
7QwxmbD4GGRZUoN6MxvoJc5rsB4sbIBj4XSbYrupnjMOmTw6OfJjmHaRmVOlkWPV
D6cm5xqOkboK50vG3HXoTiK7i/iLSF7oDFtLu8oEBa0jS7GbKVHfPSCUGktLcFT4
Ga7aXDa8MbwP+wlMEulTzHXacWBV2lRnUAJqBh97DN2vW70ob3HDwYocOgEBMGQE
4rWQAqgE1zJifV8eVxbCwMNCAGYkZ8iUfQ5uxCoI4cT7FuL64lRf9BCtsjUuaEsM
VOucqGtANXb+c8KOMYmSJ/iH2rlDY+rrkp0NkcMwgxpIiPKNQeJRvX/cJk5/w+V+
iQ8+xZTxBTqt7r42+PeSpo9cEpTBohZIJJAyCkgv79S5q6D1n90EeUa1gv6bVBHO
eEQv63ZyZLLhBrGDXdO7qi96CDnOkkxAkjkQdoq/8eiogZzQIaL4pfHLEQUKUTnW
P21PD+vfv/wg+TKmdKdhe3cPqZk0pP9oHDlHzO1sMIhcRDnvNLv2GyLoEKoOO9wy
/rHTnWll2VFB55OfVNJdwpn9wTbwyNj+FcU2Bj3Ht5kLMEUCltZ0K1beMgTSAdwg
BcyVUmSDllTtwVh7QgQwfdIaEE7mH93EGF6NF8R70SDY1B3myHDtuqHX2onfne3A
yO0UHt8ouMyrrgYUrA5kSP6asgUN+av2jGhyfGEANL3c7a/t8ZwMzdDEDwOXzCnF
rUyuCsIbhTfBODk2T3VA1Hl1kfQOaMpdj4MywbaevmV3gVLBgXrVfdvCQFnGnkrx
7d/X0huHn44KGtFJBfu9ZZyN5YAK2e6GepRueyi1VuaQ4gb4Rf+sxedAO0xVHSCF
8KTgamrlR7w57OOAIQKkRizIZCE9un791Xwe768DdyS5/qs33WKOjujFwlsyy91q
4Lc9Knztx2zlJOZdM2o69i697BzfcKxOU3L3boAx5EviHX2g/4VTBwpPF6WFMrfQ
RHg6cOrk0swXMHuthkRliW/fGK8Wj/2Oa4WiYjkAW4IK6ByyJU4da+9wGUTZoflk
32m6kr5UQ75w8jWtBBFiT+qzCnVAxJA6CKAeza06E20texcC/nqfNHx3KtKQVcmp
vUllqCkG99N4yUtHFpoNWTpxmQdOQ5y7PjGCAfczWP0IX9+3+4VKwdokMz29Sh2+
ZTrSrwmmXNNydJHkbmWxo6Ei7gBchpIuKhLBMdc5s9fxjyzZB7r5W4JhezGh0COo
qFKE2h8K1dQ5kKoiwkAERGnmaaetz5S38nu7QPlkAvL4rMzi1iTylb1gbsNZJ1vL
wXndDTrpQJTPLKIdhsuvPnOjVgknFKdxAu6RbBFjsAgQkABR8pReZR3E61BjpGhe
kx85748/b1m6yeJrD9ebJlbbz1FyqPpWAlQJs1Ny2DRi7bERaLSAvBofD0dSsBkz
jdewDRW5j2W2a2XGUMZBR8l98F9HtBrvPGli8G4RU/6H+ZjQp+IuOGUOuTbaIrYk
G1gWUbZPvOEGScGzIXkARIkYTXags27ZS9k7AOcswpaggq+LApznk3N7my9ZNefB
UIdYwLeEFTMwLKx+brhx2FxK/0onCxg55O9wjprB2rifo502PuWhst91BO2SHDYJ
kwjz2t+mOl+Tc4hy2cGiEgSPB9nZrxFWr5VUyAWQieSI05HD3JKwsv6OIvgEC/2L
IHsH2M4XF+7xrJx+xrE6Wr2zjEGh2tN3VKX5k71UBzm10j28VBonOjs5gdBsoFje
J0V+3ea8m96tLknnj7gadkXE8W5xUv1j3Cvh1Ae7LIXfcdEwro+rY6+QWXHuVzsQ
KS3pLxn9ls2UXDhIG6V15yZEaSNt6u+b526F3uwXnjbotlBaSq+Noh6wdpgeN/8t
YA1UsHQrewmL1qOOajqlfljOKtLRZTDtbSc2JtmTxaDis64+wgHWBYc/VZFsoMmp
TJvbvffCQfYMxDm5UJvpsposSJlRycg+JXt6WByEVb0g49kQKWyjf+0jl01vdYMD
2Vyz6aN3CaRueGvMAQIMX3SRLlBJF2sIM0zYS7Q/JetHlHHv8D73q/x+YecVohYc
aes4pBmgadNCljicMgc5t5THIRylQPEvj/3fYkPA0G/xpbdyRSRHLK9JFpOl72yC
znQyn5+uf7dmlS/BWUqu4oTAcqmbmUbUsesKCv32YBIA3uYmTY7KYndWUmSiX7uc
rRhKQhG4J9yxaanYFxfFlGqWlQ1BxEL1wB2EtZwpskuc1VEI6vE07iGAES/BkslZ
eC015sWmU07cWeKSfF5P6j3XrNahjWIt23vvkv/F0JE4E3GFko5Ps45f87qG6FJG
ZzNXDYxN9uWL5iQzGN4HMo5+fHrKJftxdqhQxR9cuPt2oE77Al5LvCTB5m5yUr32
junGK6C/1iUWieLgvTbwYpYr4KWhjDyBQfn6yur0ieAaKuhkDEX8hRhcz3veGr0D
LHtBjyulnUW/jD7m+EXBOhtFIL+OeLcoIMsZFuSmDypVyN4escGs8R3eh8dbk2Eg
AvO7Erc21oUfleVJdOSW+S6n0jMCsJjFmLnQA2WDoqDcaGYsn+JDEsMLdo65Raex
jpgdU/ja8+4klTWX1z76EQ3OzBQqxognYFGLpcJKdfQmKEi+1rYo4ypcrmPtrHqY
50JIKi10DkMBRJcL1CrBzYQaak0SxQTz7H9caTXa4kqzsgBeo4eeITZiZTCCR8xF
21jNpfmxzrfJJ+Mjk/XSGl2/Pojzk55P6SoX3n1VsiT+hf4Gz7cIYjA0IGhsLP41
ou1TP75edLdO8CjsdO9om+ThA8jETZzdPUxRBkJ0m0zji5xdvTa98tlRbNLspotr
wFSE+v7Y2yG1vqzVGbas/L5uXsRjhUprlk4bG5wN3holuYAE6oszX2ypHriGMvuz
BrpVM3/S5mekalwgnJuNVap4VBaWBIOeg9FhVe7fEUlWnb6EljH9lU8a4msXcMXe
E+yAki25/eyb26iLBHXRdGhNq48BGfItGLdzWbuX8RdJUmEu65bz/xrg4E9dFaRs
vyd8488LchvT7ZWWhUixra989WK4QG2WgVNgdOdY2MIIx0j5H7ehXw69v9C63Pke
dLU5mNSf3zTlcgzBYLOUWdYvd/iUFIS33BsIKVaNcv6P/dyWWK0P5gqwnueud6Li
pNdxyy7ENo+/mx31o+8Liho/oBhcUUbgxva0uxYk42dDeZI6aiBHfH/6TidguREb
osA6hLFTbdsa8worigwsi2Ex+bHa+OFZ+kHWLWCWaB0GCcZtmeJBvtGABz3uWI6d
b4rWrGpc1pf/iAzak9oqmoEsqkUgWNf1E1CjofnY4FJHBkFazSmU31fdDLV+wwN7
IC2czhdp0fdWod/q6lws9Hm9JogqtrH+66HyqQ3URaqGZdrVSIaxI87Oeg7G63Sd
U/rt53FEHd7b7aUo3QisDG6szNvijS/UAHFrth5gNFJlKBc8RzCahwFgC3GxYYW3
DWxsWn9aEfAiFfFFzNuKqDqnyO0wz3ncBOhEp0BqH8HdI5Jy8LCeSPWt50gwH2c+
bvSiBiC60ey69bojmIcnfXULQtFj6DcKNn0pN8j2gBX2mLQeIdboIyXUdaKloMal
KBZUQQCScc8O01kV88lPSDYoWHq1Yx9sX5hm/qVQBaxzv9JDncDcKGIRcRpEDaRH
gmT49HsC1iEe0Kp2snxwGQ0+sP0K5XR4u+Q/lL/6hEF6BMTZPZUqZtB5E1/cfZsy
KrkW37NvLFgNRfW8QDCJFuBdXzdTN4oYfCtXCPnGhIcp+Pr1MjxKrfAz3blXUXZD
W1sbKETp5BeIbD2QSFRVQ4l/Jg6fdAQpsfqjlZPATz5oJHah9pxLNgVWnusbD5VC
5SJfAHGjo0vvxCXYR1tXLkxkyMifLp/3qHOAjjT+b9hynihcokaZ73iWfWRjY68i
aJuUBgczv11vFpjmFxY9B2jH2yTXn5nTJs1U/uxifbOhGKvCpCmLxKRw5nDNP4Ue
ya5fpsEUXST3NFi9rAsIBKoeL6DPY6n8dtTbYr6p9P1iESH7g6Wnr1oAnom8OqrP
/6mjfvJ0fjimrzGmvmUtLw5t1fgArib0XqOYlaYvpoqTUGPv1+FCo2NxxJR6x9za
nvTFuSWyuU0ysd6Dx3oxEFjT7SyWINgxz4XXxz4ciriYTqZmoCqxOodJcufH7tQ0
SfWbZcq0W41fhqxKEp9A3DvvJcTDQIceuZ1wGbkadvKi6zembqGKqcfNKTVemqeD
x0VvATjJzSkrnz6jOjxuaJWLibbFOcV0Ux9gONSfNqtW/+7DzCE+3o26zkYXNfoV
fwxhXuR6cMoxY/IkwiJCUbDYqwTWW+oI/01pmiTePZiJwvy47lTXNnaQ5f7vAQ+q
r+TJhZRT4vMj3Kj35Up7RX4PqOy9N8c7pltqQXdExHUKWIOYbHaTkBRh2T+56oub
65aio9hXZdxY81qYjTn68srzvvIjy8YsC57xEcH78oFEPA/BwOTKyLmIdQGmdOd2
lEBLR6TUT8vgf4K0W3BwcnTmwanL0xKAT+zgn5RXSchPc9y9YMk8/1jBHmjaIc69
EYqRltAh6K5uCTCkPLI+14/9m/iMRAAHJydzzQfolNkkSN5Pv4AFnUVOzUkhkxrt
zNgs2A2/1jvKKoZ3FSYLqCXGch27HSre5t44tMYxAIaLvD1zG3zfb7Z+0cZok0eP
kyUsD1RRiODwhzUSLH4HyueZsjogpILJRWtfNSZm8qSWSpq9i/HF8Xw74Iri91p/
5rp5kkTZZijhqiy97WMgUJZ2GBdq9XxldcAfO/hTmZTIGT4EtwdwXmuVMCV9n91c
kui00CVzquhqGhRB6UdPkWsjUZAk6kHDo5XEix7kvJufFjhCoqne2H9whCyzIPpK
S3d+W+HyEhroqTZ1oZyPGcAVrBiVZfULAm0UUMozcF3KUiH2H95Fbp+cS2Q0DjoK
d3shbFbIsrIPrSdf1VbZWshxohsucWc6Jkb9W1NGabtiJlbcmXZpRJ7D0UIm3bfc
GmRKYi0Q4DFOGoOOAOEHHlLkpqr1J2xHXQb2T9CchGHG3v+oI83PecVuOdnR+97X
y6ExdrsF1k0d1cwrsyO9bUuwCN+7DgSRJqS1pngN4jt651SFfNwv3p+nGgY6gOQM
rCSz2rXxynlWIZY98p7tF0mOvnxlXYF8UAk/9JFqPvx6o/6F6r5cDhL/dQYwZjaQ
8fJBLAjrjx7N8FEJGpMpwXy7LJ4u3xyx5hkV29JQl8ttg/m4WDQx9GVkukNZ1/Cb
+0eAtGyj+GsKujXzFKoVAoztfLEOYd7AM4tZIA5z4tmtCtr14wM0UB5Of8JLPZly
yQS6v1qvFcoV2KgtoAPKKQNsianYae0G5D1NQHakS29thQIM7zgvTeqIYdvetnWb
Se1+d9ikC6FFNPkNONv2yrPAUadrgdCAWjNDnqMeTv56sHs5de4oZnHE3+Pn50PU
CHVNjK3V+FTJHacSgoEPET2LsWXZpYVxIGwbJCT9N04NZAUmMC1cejPTJWhDZ65V
m4UbUwk6Oc2ZTT2ZZVbU476y6pxo4Gd6Sv5fakNkjNFSSi7rzIn7XR86QCifK0Am
EazqCVHmMRngb2Mt5GXL3ffZ9PhbTFVcgUnP0S2oPYrtCDwBXNSjPK/0oFM4wcU+
wzMNFy9786WpSJuuAoA2YePqII89SesMBwZF4vxU93XKMRQsNtGykCk80WE4SssO
E5pJ+LCHd7u2hlMPY0j+REkKdzp5DdCkjaO0zKAORtvfVX2Ss4QyM4Cau9rXmF9C
C3dWC+rTH8GTzZ5iJRTB4OjcPLjLorKeNimLKPYB7k30WWtRgGefALwQF6FIYZ2C
G2BvLZI/fOQFBuUDJJToy0Azq/vs4Vo0EAUPgPuLGnCOSIH2d2iMJZ8H3CuZ1sNq
jOw7FxXaTVJ2L+PLrbujohQ0qILLiP4+uxF8IFVeb9x8yok3Z3FYI6I2vK01Legz
IaE8d5h3DOZD+4wZ3UZkeoy7dowdbFYJ07Bhs7v9vQ/U8sk0Hpm0XwbWBSM97Lr2
Iyr4EbgvV4G1Q8cfvFlBtYewiH2ouWzSZPbOAbVyPg4LpaGwMPBB23JJrkMAyml7
x87IqnXVoykajx0N6Ol2eOo+deHc+K9uCBCbSFnjzDj6arOUIdTlWUND43L5eOJ7
MaSjq/6bnqovPMYLGJdDqO4QVGKPrzmolreKzA+xEjqGlvIZFXp2n884TT28nKi5
matW12oHV6fjQYaB+u8WQqZV8CSV4mVfEStrHC6WnMS1QeUQngvfXzDyN5/dXgTR
bXu9y3s8picYa0KYTPhXvKjkkXtCP+YOesJivEH3wArHZfsBMPCnEFRlNtkD6Q0Z
94Ixra+50CQfpWnkk6c33tZHV15iwSAGqC6Fm0umm5UTN2wFXkJooxjBl5Xfx82n
gonzX4r1nRT1DhKX6t9Taxe9Vp4gTDC9ULvKtJyY9YY4A7juMMHAxws7kGNU9ane
x7/mZXAWSHICngOWoedpov6UWfIztnufhwnWX7EYYO5J/+JdOTkWWChGOjT0/v8e
PVEyndk5ueOlwdCGNGg58wx+/1kErRcJnV8p0xEXnYFsZIBxyE9DFBxBPZBBo8PJ
kgXgCQ1sdNSl9KNxOAG4lrliG7TeuS05+NFSWWnwZYx3+2W1d04R7VuIBUgvNf7p
VrPtBz6PQOtCqvthM60cMwcGGE8QTxy/8EnOuOX1uXKo/I9Upkwpfhxc/5BUYkD1
m8yE5mUD83cMDfVEwFhAqJxJExsqQ/LaFge6EUEKrRuILdDLnOEDvU5DRaCkZlqP
rq8iigTY+F0Lg1dPXg9tGyKFjs4dEQnKo1vNRBZCpJPGZfFPIhzFKTTuFbr6Kg27
16/TpRXimVfLL4SJbFaYnZys6SMuMASQ4t7Rme5oyWoLTsk9kE3+ipX7w9c+XCgc
stUAWb3Y/Lvfuhtq0x7nm8hwyuP3KrBCCA1IbAH9UB5XlPxepUyZoHro2IJK9VsL
jWDI4tNpBxPTUeJWm3T5dUdYL/Ax/aDRvkmVDSe02K87GxXSbdD3QliJDJ/3KbHE
hLlmArLpjf3N264lQK0qx5dTsPyOkMx0Oe6tJa+NovPpOWrvatHdxumg/KeFQzgI
ubtn4wIrznmKg0rAFePgr6Pfrhia61Vg5nRvlwJ/l881R0i5oW4zDksS2G+DPFjE
Iia1bYncanV1lOgZwYv3x1QgXazscIezGNmlihnalLysUdryaIfLB3gZUTVuEZf7
RIJ8ZrBWU/XC5HDNElCR+p3Q5XArKoco2b2KCpAhjQRnonMM377L5BSZgJQWazDV
bydQY/ePSBz/3nHEXn0VWjYRkpENP7miiaqe3aGd0LHiSK3QHn3/aIvpkYGUfCdj
m8yNGXnoy86NtkizBkuTAMpFFZK+OnYL4fkuFVx09q8/OCjcGHj/0MDvAcgsqpyW
onaTQ45jxzBsEstLZlygeF72l9i9NwaklDFHU3YVpsqu6vv4ewbB/tN5BQN0QkAc
J6Up6J6Y43YtYW2a38ByRgg7/CW0hvr6QuLQvqE5cQbNuWBtOy+WvUTihMWeFNnu
Yq3DAh/xbECDNGmw2VwQCQsJkn/jq6Tg+KvzB7etoBzL/908ybk7NBSt1OfQGRUj
BNGmYIhkK8Qapm5qGk3Mn+l85ApdcVM6UTC6nDGBGs05J/ZY8CIrRT/CHfxKAcZr
df3vvWWBU+G/GQM8h74Bin9cvN1EtS06Dz2Pxp+RyN1Bz4oZ4IQqC4HTrLqfiCLg
uc7ncIZsHpH5DASKxUDJ2+XQyrWYtnaxGwrdenqyaQ0jMEEIncouktjl9TeYC99Q
DEIVxFveE4Fswx0RkO6qbgIf8KgdXXijFeQqMlAs+azkx6BDYHUmy59WCLgm/pTl
Bk/80uTY6NaZrKeLEVuHk9TROOTLCOB4PxXYUN4EMULXTUD1NkYlOR7biz/j2WYJ
JMJqhMqZmpZ9JA0Tjni1/8DCw7mBsao5SH7lD74FuS1k2EdYddHUQZFdyhVlckxc
4z1E1z1jerL5MCLI8isTFOjUb7bLiSJWxNjYyOF5wauCVkPV7DAaO2WVK3A5H5wN
hwMOH3Kedzb6AO1PlWaJeSe2odrriLvWPcRNUx8NmfBhXDbmDWu6D4hGGKxe9vov
whruEkMkkPlX2eIgO6he+2vL49Oa65Z9ywcCKyfa+RlY5yhY71lB87kZ5I8/NZru
04x0w+Rw3CesEcON7y8YvYvWZV4OlwgmIdo6gL/IC5L+ePbdV+rOswdg0D8sG/jw
8xREutd0tjyyFhOWfP+RJuv8R1271LRlw2JAHeDsGlyQS17t5JCn6bm8ioR/BJqc
AT3NpiQPwX1wyg05hvnvtczGseVhVGtOvWYFkQk3w4WZhCdjktsH3cCycjtBYCOd
XPAOjvNYaymr/K6N35Yc23Uk8bTDz6S3KtwLx+pPMCavhw/dxe3zZN+nYty1ghaZ
p+1ijDZOXx3VLqW5r2S1d1P+x6Mqcd5HXR+nTl9SusvEiJOoS65LUHzMQkwGN9Sq
BQHkmiRT7iYJEjUFdY79XyoN/x8aeKYAilX7l7PYW5mti7MV1M+7Rer19YGLY7D8
80pgykNt+wsZ8WtH54SHJxoCsR0mSDkLwtdjf2WDI4bbP6oq7w9MnwIo9LZzIHcS
R/iKTuMuNS+BcudiRjE1ctJxpJbOVupS5hyM9IoIeVG6F42eLNyrA85yacmxBqkm
Sxc25Fjr8BCojRfmSc2glNrsfsCknWannDT2PJSWD1trqDhouC82TLa6M4+nZN0V
a+msQB/O2dftDm3+PL1aag2IrTKLTGxJADvtkOJflXV+YCTa3WtyNRtLPmPD8y1C
KR4U1jmRLix0wfjMIcwiIQGGgepgxjXHoG+VZP3iNdBPtQxzEkbzXoDWaPk/pt65
UB3RQ5PQg+7u5UYVv6xlHxhHD0SwotrhNomXYVfV73zk7FnWjtS8d5tPioImAbPP
wFZsZ0eXHgFs2N735T2aee9GPo4n9MRin2TAa9oDLmHoEUQ3Z2Go3W1Zf2yJ7ZMk
KlwAZgOhAeknRWQ+onukyvd/2U/7GMUJV9amlp/lIXiNLfEoSKzucIze6eSKMWk+
z5le7RAj3rUBCyIQ5FKOH52xkKZor2LGKpO1oBxwnzeHM1zro0ysWuJWXhHLVXMm
bUfM96g2skgsPCp+lpyyGUc2W5qi4GYSGxzj94qmBc/j3jzwj4DZABt/q04saF8W
sAasMmJZ4UTC6a/iZXuxMZeSFwYxPE3/J8KxtxUnn5b6YZQYfa6QfKk37rgFY1on
TL109F2bCAQpX5Pil55lFw6Eh0fIIx2Te5hEEjEiQY9ht/XvJNhcUZjmtFFey+D3
wUovkGthay+HpXW4v+6SKri96c+B3zjKfv/xt9Cd9zJDEzpRs0Oxvaqn1xn5I3QX
2jxMqMXO3ZboJEXqmb8a7KqS2wVI+oR5RhsPEWXO3jZwhrgGfY8ufQY2ka5auurV
Rns/clFCbWDJGrUMh3Qubcy+NM8S8HDWJan66P1bgK6NMCxPwJIb7atyDUbUMSUK
FYKQbP+mWZaRXF+qK3v88ifp+t1J1kWkgAbumeGh6io6ToJoO/E7AQvCsxWQ5B/0
LfuxAEnXkxIlCIawAKto+sIht6rZ8VpqkTMFyVaPxTdjvIW3RM+7Fb+RCF4i8T3P
14wsF+aBhylL9aqWwg0ISuQ9lASdqXZKQlREC6eNWJS+UtIPc1eDsGHAs+JXhaYH
XoR8cCXjqgcJ6n1Fs1ZVCtqlFKy5wvDS5pv/0xl/G9uVv7iK8k0js7ycXmGsJoyZ
VLNzBV55oyVgkluuImIlIL8bUEQAQwAZcDzfMLesR59nFPeCKeq0NK85WrTQdkdc
9tNqjULHb4+naFVvmZZDQGLk5tjxeirSVZOtC5H/H4W7iJuBSjN+s2r4ZoIzztNf
QryCeFKOZGmnMmwF/gnHRk7WW525vWvcLzuqmg6a02Jy9HptLDlgZlVirChRDKfI
Vb/zxhHMywpdoZKDl2/xa+HglIXX1kvKdyjg86ZsdgJzZutVxBDg8ILz9m9XFvFB
6b3dYG8poP25L20k31kXqOymuoThGIAPAHst4Sj5dUf99RHnSu2C/YRO1Vd5RUEb
8ewGkzv/yhvSYBetQIXckczOTm4FsdV+UQXera9nk7oyPcxxV3zr56asXnQ/bzBQ
9te6FyKu9hnzS2OVhc9S+DndMLkwo8vpjD8fjdHLk3oR/Ufr+G6dmGIPEiQ56LXN
GP2gHTxJLje62pDTkFcMztaw0ldWrn6UdjghQsNV4PI7YelwTGTmID2LoYITJz7O
CuORN8maInQevXXW1GO3sVKgfbx4gmtCEMXACFHpOEfK2k8j3CGO8XtkZoGCxn4r
9V5rnT/Bnz+t2LEOe0OwwnKz4tv9ay9PY5dxkDgs1sqKHPNPyF5AaaLK+GgGbciZ
gTL/SrpaOMqSlTL5wxCiuCCnZKHa2eq+zrVCB+rePNfMGza/sMjMM35IqyuYVnGk
UjmEHBBWhg/d28uhOhTtAF1YsZWzOf5FHk9HdeJAU7fMpazhy1tiUSYjDxnkdaHc
lbbKK7WrwaRWUigCSx1MIp75P8EvcPM90GO5Ddy3cw6FOZ83BMWcFAy+NaG27BeI
ScYi9om6A7ujMhpDuY0dh2rJF7b+07HxNdO5sT2YdbZX+Vc6fHLpYoQ/UjqgJgum
LpR3UGiz1PruC0EoGFBzJkK7lNhuf0nc7h6zGJSmapECBWz5z9RhmTbjZoy3uU3J
wzPnlO6y+A4EhBE6RzyWMrmbhhW6ayjvY8D7WO1JRvNcNkgaATTs0q15w9KWGAHx
N2POgHNRFqpRU/OCFoBIeT9K+ERRRMrTDuEZuV/WakcWMiCrjA7YQhR7rnFxkLQ3
iC5+8J4wsYo22JE7eaRDPo+KLLfyeZTRRiicTt3D8bfA3qraZcjgIapBa6Z6gGf/
yp1EmjtrUqmXciUPGJ9dWNb3Mt+HtD0MNQhb8NmsslTumcFnDJslA+1gggWDMiC7
DOdbojedHpTSudpfsMfzAGESgj0G1RIqAqsb3xZMZMdAyKVMCHL+VfoERfnO4qe8
ItiPlw7BnEh82LEnDHyAxGokzzc2oXyopigMJl00PkcgQ5RF2czR+WN6zUTC2ogv
tG5NE8YZhGecB1sYV5v1/ERAMbxi/PjfyW3WsiMvr/g6L8/1N/Y4YktasPfOmQkE
Yy0QUQSlQSrzcfJvNrHXioA9zkEBAJjKzvX12dfl4Ukalzj8UIWbHkfD5PiaOMi+
mdXCpz/nyXkwz8hHmJTtd/pK795q5R2Z3S4h3Shj8TLFVt+AV+1GYQJVM9+dhOuN
6J2dhfmn85VmCFxHmXUVp21XHorSXe/1LdTAqW88r0EasDf9IxfQxYR8+V9DwoC5
coOgrjbNnBF3bv0gbYJNEXYSUJY6uG3PaGN2YROQuPPK+jPoNb32QWjf9oey1sns
zDZ8PDCXQP9zL/YeT7XTZA7DcwVabctIrZI1jjt3BYwzh3Jx5J/zuJKKWK9oSB7B
9kA0xCmSJMBO9EzoKHMtoq7E33MhgnNwCKvUlyzoPvpHN32aOmyh2VxRkc7nAD/z
oLmoCYZfnXkMd+F01Z0kvpB5ym9gh6ZuYjt2Bqk5+uTGYnlnlnZrObaM3XExA56t
M0jYTZ6QAZkijiZ3UzeAwYgj8hgUjl55ybM9AMY6Q2NnAtGz2CO+PkYsiSC98qsS
CcTI0l4zrGaMjDEIN4e4mup5S6g3Nfzh+yqMXlfqMnWy97YY9+v6fiz2O4goY9/Z
y8EOI2M57olNVmrqxyzP3W1WbpYS46sEZHNk9fJqhBgqHB4D4FA2Bynsu+xq0Km8
G6MQBa5AeRsX9W6/4A6hVAfeHXEhd4f/6fkm164F65cFjJRw2jVbcwLRRxxZ5Euz
7AMoAPUqVx0tMGY6JMePP1n5c+UoJO4XT1ApmG3G+8Abju6rsfcAK6sGyyBVGLsz
Voo+7uwpqq/7KcFFDs9NrqvvyKzoC8RMkLLz6RXf/34TJ6cVZ64xqa2YSqcImWf6
Tv69HJ15fB6pPOStAWK50CIaUeY1+XmHCT/GV4/5s1tU3tbAau6+GcWffurPO9MJ
SERhD5kLL8Z/qcARh4BOIkruotXX8+u0mTLqMaXwSP/ColRUpENAEoKOcMfc46B2
9hBxfNNLJvwzGF354WmqAhIdrw3JM+mwESK0Ao8aBt9bx9Lisle24SJsdvqDaxqG
Su2DQ63kVSE/W7yCl1/KRHL5HRuz43o6tsskBH20g+RIcCkNshPmopQeyZ+ICDUb
whS0a3+snONL9QgM+SrwJXk+ZjijNWG/8+JVr6PZ8mt6OAHvaY+g5hKR7UlOqyN1
0849wbZBTQbFmS+EoAsYkfRepLfrFIyN0GioghtunQpnBaz5o8+u0oGW4PJcMITr
b43jLXn9c8rvU3pmAhZ26weru9L80uLd8jLF93F1smKycAuAw2a/PI43DbTK2mc7
7ioyaXEhB3mJH3Xz3khi49gm6Dw5M+A6ibAUrN+3Z0vXq08lEt5OW9YRhpeQyjJT
uA1bPz8+Mku4ojBK534LBdtdbFD8uOVV1hR1cIeUHtAFdrVQJjmNCj76u1GWW/s2
uFepziZ0+GIu3XbD9easeWkFdM++sivclqAlwY84EzVl/KBCGIv/TbkXebBT7bm8
zEyRmOAxIgd7P8h+zx0R1PgP2XtKF22lEpqx5wSynEPPGqRnil7ulW09z6ki/ONT
hZuPounWIN60hNPKPkxNIocGnchHSYTIgh1KjHTfDKiQ2ypvfhfZY3J8rzrXYJNw
E3QuLe/XUe83sSxTnPGKxpS7QLzmS2tMCg36jlFNlYpda4Fv7aHSmvdMZ7AHdNgI
1hPheODLt2cfzuKqjG5TOtst9+oFrNK/kS4Jz5fGDIBAG2ftAMT/PfLJhmOwrR/F
L/xI/tPzPDxrA5b3V9wdykErudhUnJlyID3TEmBQk0NJ/24MTHKt8H6xrkbiofCb
wPIqMGJVA5NZD/PcQ5s/orGAWzXJ+jfJiYROKiAmST/LJSE/JS0eNH05KtIolu/3
v6Y9GjMhq6Qxum8sFC4nr6wOaLwd5o9OR3lPeVP1T3Av/50j6Dy/pMz879iJExjd
SvdlesYO3LWhCfkey4Lb3jCW6Rn3wVZBjLtff5c74Sm4Xwrc+TgN11Y+ovaCdc8C
UZYp1YJ0BXwwn2UmTcN2qwb0ZQ3kxWRxvqav3uCmu9SfGRZzyIZiLaMV8IbIHhkq
gpNLCwei0Brip0QY1i1DgNqw+7Noa+6PhmCChdcQ1v63Irg01OVGMmi22PhkltsY
oRHSdXyT85atxlhMA0bdnTo99qziUmLTsHkL/ivAVUXTgciUtISp3LaXbDuk1NwI
HjkR6Tr2L0cWxHzW1sXujTOpl/9HVyVGtEPhGuiG8Wnh2rxhSUFsHWWrtuHGlb4S
AXvbM2FhB5sOgjG1chIsbLC4ktmbRmjhYLSzaHTX7AAwEzAdzqQZ/KKKFWSLQP0n
osF1LfHBNOmd8McHA1df3F3Ca/kYAeU5F0j9udE6NVGhlBP3aoNZsJQKWMNLelv5
fA6zENkuzzoyY1QmSRVNsOvC8aZFJIe06WGiAuYNiJQeMnvMcYlD5M+cUUU4wgJP
voi9/Ylp5+c+WrjGdXWabckp+afhXHV39V7nPdWtJHb6/0xPu54J3f0tXaRw9WpR
q61WdGRJjA90RyJae1//3mm3UAueHhaDcR9JFHls31RcEmQ9RS4bG4Cd5+4BZQ1m
mSSGgOjXsI1jwIar9m9xuBIR0vWMq5ca8cKUoZUeh5QNk9lvYYoIA497iXZ0ed4f
ptLlCnysq5fOUBEOQhxJDmisJGg/KkbzK2j1mzQSKULN3m1tDPEzE5Ay2MV9tRh1
b+MYmi7X7BgqoSxnRDutTQtVTu/XMQyYjsmqxXgBHKS5cuRnNUlT+ujFpcFmD4Mr
s6q/q3qSVnufcizUlASrVrXSZo9zzjJuK0/L432TvsqI7cWeGa49wpKx134ONA3B
OE5sX7k8u/Vs2f0RKTfTKhZu62FFPAu70Yp78Wn+7N0kjGSzg0P7AWoSIo1CsHgQ
wyu5n636QvffVtrQ7TkDFLzUaiaJScwQyQIrpdT20STUIawwA5OSXS82mc1tIg3L
uX0u6dsYmuM4C7ifBKqPZLaE69jyBe+nhaH5uwZ6sldGfxUY184OoqcErk82m8gd
uiPo24kSmdqweMtF7NkuJcn2FBLNrbmB9HCWrwK1+pySYXl/tsnNSbyEjygTL6vv
MgwwhbxUlD6RJXLAH9kDCVxcr/PoACU/UhNamlSB1kgZbmvnC8cAE1d6jtJJZgI7
cXMc1A4B7e9PT/AiDdJ/YWMzgfvOWVbVTophmFdOZ6BNOe9isKvSUIr2z/IFzaCW
s2mzQh5C4dj8l0tcDiAI2S4WhhZUa1KgKsiWLeBqRSCPQ5dv9/Xeo4SAoJscvX9e
rnBYmwYvD2kKIS1wSEwBCJtkxcK4kEZPx4bGaxq2zOSCgcfgPqOCILzFUB/ywTqO
d4LyPWWAyqDMYHWSuQdLfFr7T0mQyfjIlGSdo9DfM66h6XeyCqszmQdut39uJ3st
ShFwopNMk7yibrWtvS3dBIVO9+4fXTH5I373KB/CaL+02sHrYIOm06g/Ibs+5Anx
G2IrpgG1lTKcVmrFbp2y7tiGhQSDCIU/Ftp3G0cb3UjJ2cL8Ks7hvlR+URlfskpZ
vScZFGWL1k3gQDCD+IRze7TFQ0PKarGuOPGVmXhAbRol1GZTxya8HLfnaLs77G7j
rK1LGM2oUBsifLiYDYhsUUXqOQWv4rGmgV8yVC6R52vr9uZGsdo2l0xuwUcGPDEm
99/Rq+rKZ4/k6ftcxAOydGaHrqaBPUy7BDzbXFcjVyMVxHx5lg6YHVok4iq31BFG
aX8jR2jcoPQlLuF2QmGiuGY6AzeEQ60PUr/hYYLuWAFdWKDAbSuOPSIRxwot7Ucf
C7ePBSsWIaE0JORu/YcOrRj9sCTJyZ3xY9sUmbd/zWB4J73gvSBRwVGXPZvgYb9y
mkUrpQZ4CbtGVbTSeRGTC7mw1jwhOKAAwWWppFcBiC8iLHmsmUaVFv4mRA6usOlV
V5/QGjKz/3RVrPhqOxQpKD2sNfpDy02oOT7xpOxLJsobnVUC31r6U3mIRjqN1t7p
iywmdWhTM0/k1bymqejRyi5nC/D0J755/sqlnj3EEDnlxkO741q9bRByMygMoyZK
kMY12Ldoq11GcMrX+DSCkx9VkDUE4lOkAE29ui8i4zm6uTGTeFGEfs0iTADlapyP
aNWWovh19USRgYRjNeQRLwBslvH6iTP/vkIWm//rp6HIaZ4Rcsy4dF8imtXyIUK4
+b5+6h7KC4b8q7YbZ/umq1HUY5aYkMQsJYL/U7r8RKZj0Q9lm86qT6BMXe0B/ASf
ocdGR+txFKpZMmnfrCXndE8Z4bVYJsHqReFG/4HYv0ytF85NWQqIYNAOx0mIurGd
ndq8blJG9PEpqPCYwt/lJRGRDCKEC/5B/l1jStQ8tHqGN8+MEzfrKrMWieXukHft
aFfDDrwxQEbcVduaR1lzdm/wYCOCBEC40s7ioGLscnbTjEwosq9qRtcXEJIudWyp
bImZYPwJGaz6TwiGPmA5EOmvn2EptgpZPvenukpsNXKsNTJYVButG/ArPlMTQX8s
gvU1mwJJreED3yZUvRA0C2mmtK1fkWNe4bmOpMYacM3eiVPiejo42zTtpbSIz3Yp
6Ld47Zi+xhFInmzSkwvnRJuaqNAN53fXwFKdOcQ3MSNTHceBgr9LkoVBHt8kMxAX
rmwvwGgv66P5Ie15Vj2mQInOVGB4p7kfFWMSl5S5KnCEOune0Ui9LnVSIG5ysYGQ
lJXRg96caqCO/jkyDB0IDi76Rpp7A0BzNNPV9aFHJIjMOjJmmBnrxh7gA3xifZNs
KkAAMGI6IbbDr2AIW1DhyjiuW+HvtC7w31HbNoFmHo5b6W2S3UzawW1sox3Af/o8
lPMizQNetyazyaeGphRgWCX7UzwzyyTQJNte79WbkZSWcOOd5dXMzOpqLM9MeIsq
w/Dij2bFLePfr0EGOdbKyB1PN5/nQM2GXNvj0SSCk9XzI45AwAgGIDpNzeZO93qF
Ag3UbblRIaHJIVYVwk4HBL2kL4R/sAxvvPt2GFefwdMcOVP+B5A3j3fmjvrQYSrn
T+9wi3zJu0Bx1iDhxVDKdhem3RD1bUyL+GUuj9XylFqmKgZ0qg2z/KjqSPb2PZxI
XVpvac2G86uddMIUuocQqTbx4qm/aLWJ3nilaRdv0FMJTldberzT3WQcff1Dp3df
YaAi7jt4jhFoeoVn9bDkqq5syLjwozqXFppBHxJd7ZzRKQhu/VcmpnoQSfBueAwf
G3u9G+UAXXS7e5PKe7HmRcXqtxWlEyOiQq1t9EpYWAhQhRLEjJsVP5AGyUW4nGRH
br+LPzp7OUka9DCuay/pYbXLAeHk88pDevqMgsQibEX/qqHTS+HaJQgmTjWHP4eo
mUmHRoGDhAaqSXz0+o/EmxAb3SjKa0hfZLuT0ELC7q3DnN5IIo8F1ZJCjCdNcgB0
Bbfz1LYiYSaP763Embl88aGIP8Ta4IAA/nZnB2R8yeM0MOY1ND6BCnPpJSAEyO1Q
C6CSJyeR+zSNOqLEl+8PlpmCnZ9uuF9QVk7tJeDkrRcYp9ojt1rHXHJRyMoFBZb0
ozV1xGoKwuYAT0z1YzOmUaRkeFGdYnjdMyfut9tJyg0JjfqAyuoZVq6RCogQF+ap
IMvwsp8P0cNECIppQjcdNQllEkbbDIxm5SYdyXxnu7MgfHhdBRawq3dx4/NuIP44
MFbsFUwfuBVfR7LwD1/SNWr1uvP3+j5Oxv6VBnho8MiwtctpIIXtQCMbLZ41zfUH
O07hMrIOsOElF51X10tNgJX+gzU84STZHQVslheZf/KoPR2HYxPuDMmRM9gXW3vu
8dKipibrdw7uSi++qAl1pNtgyaLRmSLpnsmFJTqP0dAcvQr+u0JEuNC130AgCP+O
oQjiHf50cr5y0MCowHjC/GNwaFc6Nx0kwwopvSxg1YG5J4eqFpyof5Dszi4zr52b
UaG4nfIhucDZdd1jv3zIOsR4RPAt/CnR43aS7H0DpGthqEui5UbAm0zTnCGwLiTs
Kc2qVNtOecjf1qW6Ba6/3e++aE8leB7lnT/T98JzHQsMRRMQPOupjGPnRdgMo+M5
dbDVTLxS9RPm+jGeihRFGdMnwQHm8ENP9v5Z9elB9fp117aWg9ckk32v4YsaYgFx
fAB+V5R9gYk/LFqybTkxgci2bwwRJ1n2+Z2ueWN0o7xcIlrElG9PJp8LI4GtOKeC
/jJXJHkC3mUY90BgY5hpY9+O9RDV7rTZaTnn/CMcXV9e6tAfBD+QJc3yy6ol0NXa
MteicBZBSIRXLl6gHJ06YpkKsglUT8/8byJ5gUD37hJABq851rCeOv99QtNFp6Ha
5a3SxlmFaZ4amvp9h8L1dRsijCFek1KpzV4QC1gvYzhfdgZN84kG38OhaB/FDKwn
TlLedkNb/wf3T/wT7/3f7Bc7B/aplb+wia2+8ubOI4rv/YwaZN4RQDMoX4ipOWQC
Kic1Qosabq+v8y7OOBXT+ZVh2t5qxJvj6caUOffichLvMAEzLQ3qKHuyfC4NqNq2
K7jcKwV8lufRKRZDBNHms1zJBiyJQBfDhSks173h3WP/vOkDQVwW9O+sE45kUgPy
JKjwT9H/PqwIRCeE6MpsNcI+Iw0E7KgrrH9lSrV8b+2SnXaTrJCKdwLz+8QdBSkV
wh1wgl1dbCDR9MxXP7iQwELLww5BonCqrtMqK3bwAuZjd6cfnDWUOUshu18MlUnT
amVsICN3Hrecx26g1cozL1B0C7ynssk07KnPH4AfBsc1yvt+g6NnQ1nSs0Nmf25t
wD8wFhVje9e/lJLGEv0eO7N022D3YyiFLHVJNZ3ggAGZUsnhuO3sb6zxS7D7G9iA
/y3TP8xIgNNZMSBS/KDiu7Wf85m51ZXTu4nMaJyYFnFdRVv2pZkGW9WXJfdpnI0i
zRBcf1opN8eC+aQg2o9FfSzYBK4qk6qW222iQ5DQdbou3w03ypvyQ4VGt5huVYbU
FNa3K3pqkKWxcZxw0Ev4OU2Fr66rzvMmOEcRu1d0JY9ijNw7GTQhluOjZJcg01dZ
gTPIp8Jkd+O8qyQgXcB79Psj3x9xPBjGS/BI6YSMvoGtx31glfMQqyIX20Hvle3Q
YwN2nVpO/LNsOqDA2M2YHUS0y9dEh+Rb6GKaFRr0dnsIZz4AwUyGwH8ecTT/pf6H
BbaffpU8VvI8HC6IIkIqtI0wjpFJZCErO7ojr2T8697dUgEhrnSEDCweL8p7C+BC
f/dQFojadnuuPyo2h4YaM9oslPBji8QQKSp+fYdtfoyHxxh1uB8vAE0Fp8Z6Mg58
v+2ek3Ouw2XMCGRilRyVQ26g1QRhJdhgTNtz+ufdHzbQ3ZjyQvrNHdoRuyN1XLKe
YY+ljHElK7xW9r1Sbt+juHCsIw9bjm2BTV7CM/LTpeCyfGVunqOsK9hYZupCXQh5
SwoIsiAfJtURiQfD54GRN9pX8clDwLyq1C1ZCbtpHr3BIjbRHVfKFQ2CDPh+VkFs
P0O+JB9kxaKEmweO5zNVBmW/Xpa+ScnnaGwKazUcsMTJzGfE8GtKX57h1YKiD1Ky
Kqr6bKWkXF+6XcWnKZep4SLi8Lu/YHTj7EBeGhqZ4L2U3JdUEEM9wEu6YKYMPoqP
9GdXu7/YoFj2m65vhStsrvdug+zRSxUx4pm9qAliC/Sak4WljX5c6tw7BdATBW+g
jMnQyFARAAysfj6wSN+XQozZSypQ3NEtysQRkM+Fxomu6zQ9kWMJ/TGAqUC73vFr
6pR+GrE1o/nmAtJtEsgCLaJB+f4huL11wBcB1EtzN40h/5PZa9LLJeHK+Nr4ipJJ
fK3QJA15uxVl0V4BDMrcg5bnLA+X8tSrCSxT89KyXVI3tuPRZwiF9aA4ZZtMPMJm
DhyTllTIU+W5yUyElFEqkbUUY9ND4rO5j51hnZ7GanQyou4HMDEJmdDAJi8nGvu+
qHxNZlwEpE9JmPnsg2n1bYw/CkN8F/vH/VMDpC2ClOLufUUWZ4v8sVTGjaphIUko
dMFUmBlX1u4P9wAt+9F151aDEgQOrnPyLO0o+rSECmbmWG8Ls+dTbuhuiPFPJIhk
2Nn2SmWEs+/tBKlEkaLUrnzzfZ/S/33yMCmpnjNlVYG5tk2fP/e9V/GGRkwgHIee
/2iPBgVkfNgrqthsIQzY6kHxe32g6yBDxrUatfs3g/fRkF9f4M+PxVUb+T55z1ZJ
4vEQI2R32WTPVuaL8zju12m2Etqijwmlv/JGYlYa5nQLfHolEt3zjp+kUjXowVSY
zrO6XeZCbdS2NG7qdb9fDF+bKirO+i1dgAyJwOPkFMWYI1/CGQOnm/tnj1R/EZq0
qsNJDr6dWe+QFh8EEsS30NRuzpAw6lrBqm4nqEWLcibbOdA3nfGvn6ZdvwHAUOBL
JvIIugsQahAHMXDRdMDuUzjRIhxzEA0LBdZkuwntutvXpMfLDyTeyED78C8YUAaB
Vs90DBMnIVzvRhqtSSteCQkvdiCMNP+4u4+vdZuUanSB4mpN4idyh029nkNB0R3e
ODDE7wpTvUyENJwz/Bid+Hjm1vg1Eg91A2G0pyobPoBGCgysXrzFsVPzxvXo3PGU
GealbwP8NfsW/9TjnsH0zdlA4Iz/1t4l4NGauD6sibf4GHzGc/uwxQVuPB/J/8Nn
tUAP/7b44oXxu1vUBhhNXQItjxy6RebNPjqzjuk/TOf4Tl1RMNZ7gUDjznNxyHFb
DS+uRVxrN4lIY4gsXLN0iI13xEf+EgBjBKrg3sbJmuWgmdoUez8UQ03LWpyktNE+
2n4rhL5QbrrSgl61+of0N8o2FFN8201j1BjKQfKXzPUiC/bI4DFi0C2lvihKzmgy
a1l3M3yM/4y91xRPQfz1dCxfvv1FRf6LxUhdB7k5XrE34aRKL0NZmMgFkrCNJ1dO
pxRIZGrKe+VlMj2SsI5hqYCFxC6xwMrGCVrHy7gVu0GFgDcqWCGu/oq1j93l4BLT
rpGAE6oVr1VUCp+sdRjyNr15AzWBphYnVN0+iarO1Burjznzy42gYjz28fhudQC+
I97d71XfPP7zd1cgzHKollvYGHPgXoFtq4qSWwKyxNd6U6wPQkJReSAKRXen0Zw5
JenDsuifAfiIm4DGLCDd+Sl4euvhJ5M87d9QSogfS8ZameBkoLPgLe4cYsMciPGI
L33jrDCGGFnwh7L5YF9wnrQXbPS8w+VZWUtSbw3duninqJkjE52OM7zaXBqhEusR
AwU2+cO9eVnhO1IbjZepP+qbfIApQAiKXTNCawDwVT53/e/yOhp7EqWcE1nMw7x2
+uUNAMQef2BjG5IW1w2Hl/iYzAwoo5ebNQ9uHfJ2qcqUkzrmBFhXR+muGDyuAlKR
yO2MOdl75OWNBabOSnMaqVEt4u0oH4dS6c54cIktl71dWvGFf7MDFTA8/2cGm7Jx
WAngS2/e7K+BPDqqiyFTfQQPclHuhBKed8TGxg95sthmq5MdlT7K1iPD5jyneifO
lQQqeG7SVLsknT1o/KpkHz2EbDvy6zbyBHxUFGmrwqCIDgKfllZVNVUTLCxb0C59
SosMLtrL6cvCcEKBxwT8CPy4Kj2Y9nxis4MMjAaLPx4gzDXw6kCpbmnUlixKi9y9
7fIiiDSBMyGgKbJuzvz2EKVv1Vv165qCWi+tgKKAyPv9L/3hlEWQ9a6Lw0dpOrOK
pkzJMHFpmAO5Crc6/zibkMZ6ReHCcrekTSe0pW9eKk7GmTnC5plnJEJQHMDb+Z5W
CopRoMjnqDyBuxvAHvvbljkkbmX8rWipi+XQ7idXrybu7Fzxc2sj/cp1oysx9TLm
tBjNWCRnhzpiEuYL5eNVgrkqDSaKZ/a+fnh2Ih3nBC0jHOXVhBLZ+Jczx2Kgvbci
G9SugG7xzdhMp2TMsQAP0oKl8oZ/EzH4xAvi+23jLgJoNMIJmS6ScXkQ5NR9izin
iMDVfG8H3lLnye95SzTxnQe+JlRmrW8puT35+flWzZ+vZezBvsAvn1OLDo+4nhw1
C1YqH+RMCZhH2EKg56g7oGPZwbDRtIlfP94iWLzWHgbHon37GdGeRfQEH3Igkfcn
1UubzQpRzbtJ8aBZNUmEeLQ7ydKTgz5ucbGkTJbLa1IIP7C+xtEIEWKSomWF0Uc1
CRO6nf86IJ7iE/YY18tDxTdkbZkRyj7AnIC1/43xLgZ+mrOEK+qrSyXYvcsKJ3Xi
/RZv7myhdESsU10Pa4AQARNsun6KvmtWG+MKEEc6QrFsFh/V3cFpwMEDS/uCaSmb
Bj38iiK9ECpvjLGoZ3w/10n5wQ8j2tDxraK4Bei4HypEt/D+HpReza9JLoqvVzqX
pTwSOfAVJHMIGNTFigEWmYFMd4ZI6JrNGqP9Yr+8yyGp9gjGxefShaERg5d5kY/M
YW9irmZLQpNsDtYPoKhcyveyonbFtODqS4l2UXWVcd/VlpMeK74cli1csNxs03V2
YpD2AbuEONG1I1OQKZvTmt3ZRhn6aR2pqVqFKq3DnW7bZYWkYLda7YdopHaqDAku
GKuNj07Hww5weCCiC0T4795Py9BrQx7cQ+a4v41yrFcGG2JdNWerWF6ZsAoz2n2W
4wKoNvc0eFBOX/VloR6RRbWqO7AV8hwcBpA9x7LMHfTf1eAOhryq6Y2QV/8zXhmd
H6ielfwukZLQ75Jd9gUq2TGbP7dBqXDMa+RUxMhXnuAMbTP6xJzjgD8KDFXTatqX
f/mkxLkY+J1eqqMUTRE9dRla777gMY1A2cc5dJyfImItzlWN0Gep+Q0O+va+Dcig
fjvVtALxswroHnRsgg7HLueZNXuSu2Cq2ejC3OJx7NBNsJy4uAzCq0IKUL4pjFUq
aTITcXw6utGN+F2UZ4MZT8YMLB7sf8zzy1/J+razK5yvjoYaX36FOhJA9ims0BjR
JgOb/KUqawlTm0F8RjeOnwleiXIQfa3Ldr1plUAMEA6A4hMahW0i82V7foZn+l4t
qEC7zLa/wScjPSTI1+I3X83+L5CM8JnkLB072he5USD2Z2JbU4+b+/kf4hytgeod
1XKAu0Nz+Qy4bLQevD5Y3EzKXxNNWoJNcjfYY1OOqY7kvdvqgc5Yc9zoynkIL59B
XYZfuGrkQm/ZRTH/2SAIZaMEnaxj1bQkANdgvBgFScK4kSF5pNlfaJj9MghWtP8S
pwEZw2N0LHH5KSxudlyAX26WZ6cVsjpow2iuGU/oVFSuCuO2YETS5mNqq7oDyRZT
wtlJYobnActvH4HT0rU7ixyTDOJka1mOg6Ek3ruyoxrMMEHm2/iRYoNUyP4N/3Mm
0kVp2p3Pnf14drPjM1QHK2VJgTRKz6ExXyv8EhgLILRuJ8UAD2HBtZedxZAqG0eS
6WWLPi5Cx4MTN96OOGuAOuwd2ECRrX3sB5hSz4qp3R7emQqpjLaVGA50hv8wANZl
IYtzsfDllqtHrH11WKvsdL2EQF4CvzdCFoXd51d3Whg2arZqhnFcMbHCdG2RFdkp
qhIjtGgH0PhDO9pvRLSR1x3toiHyu6Y7N3A7PooMX/Gw9B8q7T17iY71EzaJjYbV
yaRpP/wtGPw+NBCnusVZUzr6LEaL2fbpCM6pqxOwSOLT/ovD8LUO9e6bppsTbyRg
hn0+15YMAN3CS5GyERr3oksQH+4uPU0Lysb6d51H7vzTUhuOoxBrCwbzlpx0IFxk
01Gweco3S/OJ2jzEWxU8BnRGrRBCIFuIqHgDNTMDi2oPbTHYoX7XkxFnwBt/tu2c
a6fS8QUo3T7hQweMFDYGT9NxkSjE+ANMQPnHqRR9dCt/frHn8UtGtf+Lcp6QpEBh
u/rxMUtaCmYfJ8x99FGgBIWUnYtC5MHDcBvNIURNJ/jRzfcE5GlYbZAYtZ14PbhP
FDgsRz6gS1TiHPKhvhRtTkVZKKOykU8xbo+Yt96lxBlhpk44EBYje3Qt3W71CkZk
fdQzux0w9oumvw44QrPB8yOZ5RCtUyz8JVBemPOuBPnaK+l/29b+0Qe95MKfpBKR
bph/gfg4Lk6P2MoycdRHC3sdQNVo9THsugZXmQ/1mophBgeBVXgd7iqG9Io4PMrq
9OUTNwdM/ARq9PzRBmcvPCUmqycScVqfe5l5KGWE6/Fpb+IXAhvE5DEFWOneZreG
8t8Gs0fmw03NSaGp9u0CRWcu7N6PC9FnPTLoELxdnoDi7id2xJq+amfydTcltIdB
YyXkYnEHqTcZMbohNXYv81KNmtE98PylRcBjm66gVXrpeoUTBXta36tnob5z6LEO
sDLbui3/Yc9q+8HzusbLFThxvMlgZUJYZEUSxKYHJOjSBBrKDb0dyR/vpMRN0EOn
UIl6I1Pu4B4/EB9g+bVPZ6ydzzKUin4z6J4CqJbP+P3QF5ay9sR+rVFC9c+8aWtj
KRJy0dJBjvzP4Hj1Xrv6a23HSGLGsp4eMc+lmDnRUKbbarkRrKF4H8m4/pR8E1Av
au3jFH4C+7c0lETdEPyZXbNDZW0S4zLMQwYlFqB1KIBtDO9rRvEUWGFP/admoomO
/U4TbCtEn4Xf6eTHEFNdKfU8GnkzzevOy3SplX2X5Ix87mvbArmUX8Are/B+34G1
xGpyjD41/pTWFOpTK5J0rAIMDgs63kolxwf60jYfDFkdg7/R5cpVNGnQclLQ1h+C
NJCH8gtZ0F7y36dVnhT8JoWLmqFdQWqzrj92NKqmXkfG48RnJA4jZfDeOYKBgOcE
f/OKed1eY6FEuYGElNUJ1iTwfXWyF+9+xJwlDiKURjqJ2SjA9CalVTnlwIeNItKM
/8xqFkQoY62aH0NB20Sf7FE9hccXEOL92jM/DzrpIGw+MC+TuZHuYYe80dgvBhOC
G3eaqlCUbiy/i9hXgRtaDYoUMknTIgx7QuigCSbtsJKo0Hzp0HT2zlJuywDuJlXx
OdXKm/uCeIzZOtWBwtd7gmhEVbqTBvUQxlIGQj477glsV6JHjegPCMnHlUZ1YYIs
yr54+n87e5WaFZkyT1Z3w9oVqDUh6vMRDkln39V7w87H4cblu1/6mfvPpeSSLJ3j
QeY1n1jZZ1zhdCsCiWuhq25VKJVvRJ0nyfwuvz3FRY4SChHjt9YFhRPR3OYFKfzj
1QMOongiPMkA+gVtzWMyVaqRNefJIWo9GXfwdAzjhydp5px962IHA9eHzziqJRWE
otgEITJf7/XRj5FqoXyaWoLKG3Ka4tmWr+hQ4xwv53+QWTXU2iB42NzuTut6r505
r7/z7FWR5p1OfhC1Q3maul13DfK3f3OPZGqKe5sE0jEaHJaacG4z87VCYs6HMESw
oVI3Zo0LirPvPUJbcsHNl9G6aH+YmIJmqDyfpO2T1ZGKxL/c5kHM9phddja3Amfm
6vsJFE/3ImLh1mDvuGwW30csGtV35zujosL7Rfb6e4Fg2/pnddzC7MqEdZi/+k9r
udmRoIydNDA8vhuBmUtYUxelNKUdwEP6DJQ5sZVRJOqukk7wZhHw+gsocjvbsdNj
3SO1ZcLC95yztHxxOm0bOgR5E4Sset9smiMJH5FUptbebtFO4ZULZ+5DaNnCmL81
OEeHd8HNaBQS1bGWUFkw2txvYgOBeBv8u9Iap+oudoproHw0xddB/d5FiVljhe6F
3zBPJwuAfu0b3vVmU6M9V43bLBA40dFMRWWjGnBrO1FNkRvsc01f26kNHcB7ooDV
XkGYSygCn/L9GkcJd3z91812r76eUHAWf8fWwCzDIvylQl2a7vA3pzUCneU4oyPE
BNzvp4kFfkGh9ymJNahhI5uoJ17ibZwsuE/T9gpaHG4vO00gWCr23Qb5koJks0MP
4cwyx0TiUwekXAVKSZP5cH/4U08RE1BJ2Jik2ccpAdghQHuEnOCuxH3swZRSj3ba
r6i6jtHD6mAgNxAbGjA1nQWAix6r2M/WaHBpGpxhhcYvWF5bsagaJmhm0AbXF+PS
N6gYjsKApbuXqlaCZkqdIacsS6SPzk0UVLaxbzV1p/YvS65nZRzft7vvDHW8scU9
upTytt6V2DH6kdyVW6C6CNZQpOJ1aYZLEkols/D4YJcpNrUWFEXpJ+/Ere0x9Sdl
/srAjjizIwpZyM0qygUqB0sQkUGdXDsyW/LY7lVHjvYJAXnc7h5yNvkxinMniSHb
z7jKh5ATTQHtc3aa3dVQsRabE+/7HisSK/gdt0fmPBWD0kDEwbNbP+rL6kuZwarp
vU1EHa97+E6dV+2Djy/77qLpdQ5WTizhUe9rtPVYTjlMyqGnwnklo/tNXEi6zyLX
sN3g2CrCHvlhyUgd/k0p91tSl4ZP/kqCzOUavo/2PnOJTRKZzc57uPmDicR9nASb
QyWY8DuAKIp6HUxwcSKW5c+yuLolymwPxwp4mMrAHIsMu1Bl8SLxYJQqsFuhhYYq
p4h0d8VZfNO10s2PO08trodCjcteyBiut1nTEpT3tXUgcVV8IAYl6fqSg5J3RFgm
e4bh/d2wjjIkC04JCy8Jc9aeuIXJWW7s7Y0ZKjhOvRA1ZEkJEkAH45L5SBayNhpy
58Lc5btBLbuGjhrmQaB2WdX4Hma1yejx4+J2K2HDQPKrKEg07BKOsZ81BpZZf/q7
Fe7d4bAIm/ol9R/WBcR53jyGxLtKTyKEGCQZSvwfqQCXW1MtRFBTHQAkvqBuCo/m
s5PQHIXwJbWCEuFNFMIuD8F7hh0SM+VbK1IFYvBaktqM2esUWyDY7GeomoN5ICzy
UrA/CitbM8uehEnLrqnXbAAy5B4rbYXdije/XF+W3pDx5qxri6JJX/9yydkOUdyF
hZFZ2lXScmtrFZd7aItdxyFucbgdlm53PrrrfYqBzSKSPPLdWPWEVJjcBFFyvuDB
B5hgpBz6e2ABAV79scoXDX8dIDofbxItcaZTrDygq7AECkev1Bw2BKXJp2RUG9h7
oJLfK6azHHz6rdcTxEp+O1AXpIoguaU3zzImOKZzOKfVdKDhH2FdU6la/tOUxOru
GH+nv1n+d/HCqqnkw67owpTdnB3GR9abQCMXtXFaBRFGlqNGBI4ndMTeDhL0hkqb
0P8IgmGEb+ff94H9MSiZ+t+9nD+us5kCE1RukbkAUu/3GvBO7n22rqbdhgQWzsv/
Murn2s5EgjQKbhCkFeoNVCj7Dx2XSMmrUCYnzD1PdvhHz7heut/M82m4j6pO6RWs
EMUgohBKrWsBHyZoL5IkmAAJJO6NURal5HsricWnCFy6Fj+ek8ZmxlZpMhxUEMw7
8u7jMH1+s93TxtRvksuZ3yJoQp0/f0ksoRi5e5cRx0LXPlQG2Q/wAX7kk0nPago6
hrz1O1Me6/QcwAuGqqnBKfBfjb9FfmXS/KC5mclYaGdqOGw0jlY7iILOr1WX9h/Y
bvyoU9sc+03zy3Xxr/zcitWUuFj768DNgNG9Q3Db6h8Z30VglXkUSCH5uedq6Oao
UysKcCjjEfkizY0peBsq3f4YdBfKzQwZ/v/5vtfT9yTpN2ktiXrW/sV1T3iQoje+
kkyhZJqIf7INIj5m59EB756QVUSiuaQV60+QAwHzOmSf8ZE8oEvCaao5t2QbQ/pA
+gXuX4aH1z01rVQnYcHr4AUqglkNzvnrJ+X5MIC1tzCbMyyvI/T8pTQV8fEJSzS4
3V9ye3pfTLdIy3Sm1hqNZPQPQMJ+i0v8miADBH1ntDtWU1RB+USL96ZKHuqM5XBs
h0pF676Kh4tYpJgAlAOSLt/DPiTVrMffXSBLBZZGuOPGwqHpD4MctmJm430KwzoP
X59y0U7O7TaAeZrIB2mVDWgEFJ2GoHEjnqZvbnxt1qrV9K7YlI5WZ88gSCgoQhjd
NIfOi/8rBpf3uWtz5Eiq07s/lez0wUKfRPAtly3+slrcoDhRSLzGK05dK14woqiN
er2R/CcAwBH/BSdgwhsd0ZV8li82bHsY/N5s8xMTZ5Guq8lyk8iO1/enQ+RGtVhv
VaAHae+kryC/x0SECt1YryzWx/S6FRD6Iv66w7zvK/kE4fgWnad5lyetZyqnHny9
wk8Xj3d1FnO+l3ykNxADpzZNm0sWi1swH3ClrpTdZ7mlJOq8WLTVd9MNN8qDb9ve
A4hvNlJq75HRS2hyjPYpKjdrit5QD/hBtUX9fTNXd4rRgH6Ptk9AITWm+i+VDz+g
DLF3igRmmY1eMcP2BUfKvyZ8ZXOMqUupfXQ/n1H+No4+iyr83ANEMiSNyR7Ptd8P
wBVRUywek7SOI5KOZ9M4Qk68KiuE3h0WJORVSo3fxR+YzUUPiTV/h00hE6O1/kcL
Y2nSTmoNEEX+0A1Ph6NF5tROgzqNvEsZqeZuoMpzuKW22wVW2leQBzMqSVJU7mD6
LHI+mzedxKLnv5KdNeJVE1Sy2ecGO+pSdyVzwwFqte1XR6qyyfIT5cNuA9wJ0fdb
23daNiooFoyl6AwLLKgK/5Vcun/iR/ldk6cZhii+T3lpm0fm21eFByTM0+GiX33U
EUmsR+eoGtZQWckzzhgNa7xDNeCKgGzGW1+iTP2V+yZN6YdomCnqs/7Y5wAn/onq
vnqrlna/GRNB4kmcMnLhvWrckSvel09uSClj1U5ngRtSq+RFyYU587x4KfqfUYm1
WE4J99FyYl2teFee5WVhLGv6mfVIKNDWT4gO98NYajRIC1xbi4PIOBUWES7/mFmE
AkTTcs3TWP04qO+0f+lTzhC3N/E2mpHbnx24DQP/JGUc5abD5cPt4B8qyzWNG7NA
H3KjaNwXExqrGwEREPrfR5WLdPLlazbgrTakhoRMeokTygpzQgaO6Aonyuo9WeEf
V+Nz/kedttkY2C2fQ9K/nJyn/z3Ml8/om1P7FudAXSoaIgn8P62cqtHHPrlmSHyi
YEFxigajrJ1AKxhnvlP+6kQrS1BqeSlVjBkU0AB3/DKLwM4FNZA+idQtWWboimyl
1OaVCFDYmT7g0fIDbYQHCOU9YFVTtgS5XfuexYxSylbjSNKHQ7v4UlewQ9VY3Iw9
GQzMAl82AlyzvKyGveYXsR58xEPmPtNViZRPch1lnzPa+CMPObQ1/sBEHF51de27
Def70btTWefuCexH7JD2ZUDtqX8L87KJY3WEaxPWVmZqXeSFKCXM54FrOARIpZxH
W9OajoX8zLnTkFYxWXcYqnozQNJCVE8ZpfILfqadPylzMEVonxqHTnidfONVHHDo
Onuvve20FlNJV9CDCXnW5trA+/vhHh79w0/BvD1lJfmKKwm4Ewi0At53/qByHXD0
1mBXMWX/aCWzQxY0ded++huxUFFI4Qrhdh7C9lxwQNCGNgN3s2/H65PylQpsFXJQ
cntmP+o3V+u2nE+v7k/bDN4qabUctlnNQVDs+S6VTK+36SbTUyI6e9i+/ffqAsyQ
6j2qZ13AlOZ0pEiFuSku6e0njZUhazJiHM19U7duLvs80dzLXcBJBKETp213wasa
RS2axQHOGUddIGQCg4ZKO8jGIx8HfIGnj4HiGEGsWc2mO+5hXl02nNhJiqkMjzR1
B3qq5ie9HyiGxDfPCGaEmOKScVuHJCylLQRYb7L1EYnki4E9nw/MRqTvm+AcaiHL
DbJ9aPWzkSkeQ3M5cIXtVtBNzvW2vReBbor804X7Vj+8hJTD/AKv3Uxd52Exoj0o
FTTojzt7cxfDkNgVw89HHESVnfq+6LVTAIoBm6jxmegkQy2jYeU/L9mZKAcytpo+
VH8FYiQzue6FE98SraqbnYdBEueQHloYgSKmhjPAXlFAfASW314Rho1i7xU+UNUY
8RuKte1/MNVHlyq7dmW1cV+luNw6ITDjCi4QtIlEtD6R1e42wA6ppJyDArvpYKQP
rYTjkguAcxPrLlRPd5GRjzk+ot9Rlkuy455ypXy8Q2bqS70tl2mufRokDUYzKobj
QZcoXINpnR8XIWHMUijiI09VzzsHeL0cnSN6yWPkpVYAPSMoiNVyiEx0fAM8KrHj
FYCxekc5ZYnrU3Xx4QJ8epQfkgy+vDqrnyiD4WEWJ5vwaJ+/VuNbRBd5D8zk6oj/
P1Ztp1nFKnVLCOaP1vlhtBzyGF5+bT/psEvO4GogNs23g3n6MaU2CocRFRYnuUU+
ufOZNF3sWxE0ng+1wl3P6+xtfzxgNRkKfoxuXwlK+rTPHs3cir++bb5fWL5ePHV3
NkU6ZyWcO5uxpLf/pbzPSxsVKqNvioYZi+v97A4g54JZk0UMEmtjuOOX0lbk8ErT
Gy61m/JPTTIfiKq1gykJh+ZkK1LA4yxGHo11b1B/hy7CqyVzRFoAl9HT4JSXwTnT
ixcXlghR6yN9syI4Z5kizaBXTtJn1VsQKT0nC/BZEVqN4L5r3+9rm4aUigCpG6Aj
TsO89MAgBQzvtKPlyjEx3SJYgoPoT86eayMCd2SxIGds3Sn9P5WBnyO+Bm72btIN
/yeiBUWVY8fI6PcUEd5h/7eeUKII4V2dRydRPHQN50NcJyPk0GjZPRjMpE5owq49
5OysVjj+58eyJ7jLzZAHFng9Hjn5KaAjnbDCs9XBMAe9NCwtw8vwIsszh8BTltAI
bNQIohe+t6P/DDfIa6ihm1iL/ErPi8jI5cLoWfyVewezUC/wro8GjN2pWfphFtVH
T90F3gQdwAW0ebreb3388GvW31leZJxO7AheRjV23u+iyTgR7RphHEG/7qe5isIx
Ihyc7dPF6s6npj6XB1HOOnG4ZeTwNoBlZuAGEwvk2WoxBGQMFh3zNCRi33fHhD4Y
BZlciC+PsQSX58qZBqjtqaLxgFXjvAJ4lciqqX+JEjy12YbPfsT3y142eBPoD+1u
JsfloRkzN6nwcfPNr1dymoO9u9yNyXoB0Whl9VYyLlNLOtsx5PS5PMilXDRqudyj
9mCtb6DLHGWV4EvUilYtRuaDREhCx4LHKaDAzhcwQDm9qlqDtLDPW3sxlhUCIIjs
CwrBSJd0eurdrFW/nMaad2M16r7sqpXfCxNT6vJwgfujZpdmN5PJJwrNMHXyiN1x
Yn39PoKoLrPF58n2EYPArcToeT6RrRyZgT9MbspwonVz8IC+2DjJaNHzCFAQtsLn
Byzhle9dOQm2a5L4lwpCh7i/jJAHswEOA+QH3TJh3UWq/o+5poKpSb4rMmhS7XJf
CEk9sbcvLaf1x46GprKOO0SU5i5wmxE4IKE6/VuBDLeAD0thMBI63b9rpY25yqLU
YT1fze/L1X9QuDULRGpV+jypXmdoEcTXiLs0fKAOy2VPI63L3H87B0Zqw+L7ztaV
VCGemsL8nLqhx5Rx5DsaedCv1diLqRFMNIaRJP10PndcQLbFSw46udIdr9HDe/p3
Ho/9vlP/4ZYGjGNYv6E03rNTxryxRUW1sEhvg6ilATWsVMmURRV7d/wknYi4vWIo
TJSLgy29nvcN5rgwqXRTzuWRo4kxIy7BGtJgcU4pLTzMjPcaJh/YFWVXLpCvhtbQ
kFll60jJAAJE5aV3p+TTGUFIAYqDahPffZzLQhWiL+kKrdrSVOYvgIu2XqPGQ5Hm
W0CMwhUhlvCAxRSeI1/kVB1EEL7bDP5fAu8QY1E4HlNl2HvYvcVTmjssc4M/e133
+mZE/EY12h06HQ8meT/Vcj8AF0q4OkVEdbNbNe2ETOh/KFF/a51akv7NJKW6s+bD
eIWywB5YKaImePB15uG2xXGwL9hcmHYGKpiC2MbuDwlVInw+CZKnnIK+cyjv30YS
SxPAThPIWMcc04qFhXVm/cQpSusCiExfriiaykYsrbeuR03Dj1cDSUE2WcQr2dPg
Uh9yIz7wMjc0gbtB0ol3Lz40JFiZIxRfmY3F6Ikx+5rdIdiJIWkBDjFV5nI5sr9A
Hcc7SVJkLu2UB7owEWytfkEZ8bMsU8QGbCkTuUhXflCJqX4dqfRXWIWVabh/188d
PxvmpnUhQSOd9x4ocIH2kodfKI6ggeT9QbB7X/2+hddfALEpxQR8GcbDjVV9zBD0
eC4UkrByxR23uVgidHEh71vH5zNqfJyEte06gPPnPUA8pJOeidAxeE6ZnAZwaJKO
95Geo7+bHBpX6u7G2ZySuHCeElfbtHd622M83OMJPlg19lmODVlWpB56GUFs5ng8
4zOIGaS5OffMy+rsEQ75IS8vSS59/AiOJgplAXTtQAv3rjRIwEjKXqv1OQZ/VhQ3
eQXv2D3iuxxGlr97bXh8GGvWnKPwu7z2Ri5/OhzF2SxHt2P4bi9drQUJGKK+V+hU
QhDWro3bdclqMA43rCVk0nX7BWLtrOCsxPmOuOFtX9GHeDA4UrV8vVucLHw6KKAw
dZMnXPf9Klkxtk4Mz6PZxz0ZoplfjXeFrlmyf88G6xB8SDBc9gId1m2LT1EjJ4g3
LYNZOANRSfl9X9h9oLvSurdABVca2jq0FBXMe1InHvzBkcBF7aLUw4gtANW4njMj
kE+zx/WXEMMhKgMVROQfZq6SbAHg3UGJXkugjz0vWHSiDISqEnJpdSb6HywJ2382
5ZkLsTYa+K4o/3HADtSCBX8nhjd3voNj9i1zYDpCru8/Tsb8XN/2N9BdtB+/YIPc
i3CwsTD806XxMRlD4bntinTdwmRx2SGgVtLhMqOxe0qslECiQXvimSYC0X9Q+KWw
oCVgB0tG5jm494e+KkeV96eqm7CKlmsG04rFwWCgcTBrECsefIKLe9ZItNnjLapj
dAFdMAnDPgyVLap9Bp5hjNXkvQAKqwef8BxvuxmTJs1ifVB5M0oUqvBWfHJaJAe2
32x9GAJeP5xEtPzRo8QYAKUDRFrXjT2V2m+t3v2dSFjeMzHFrcUM2VRSWcHSZsKd
3RINPyQX+Zw607sWAlKUK65hH5ZGlGG3igqGyg9Xslcc7fscZE5DsDLT6D7BYlhv
y0zCFbe6MV0VAxgEYLnu7D1gbom93Tb/UFx3k366hUewockbu7SoV8k9ov94nEU9
/TktxeU3ve+WObvrpY+A8/AgjDbbdiL3QVyq1Gm73Ife/vKhzgq1IIGGvnQLgENk
kY//MmQL9KOBfOgxyDXJ26L9Dq1T+3DouJAzGvEgW45J1gkXpqQWZqaLOhAVZUfw
umaXx88YGjI/hz8jW/g7OOilFkx/SlJ98GfEDLl+YN5eIv4e3w48tvakzHPLoFMH
76yDSEjQMxGejSr3jqLHNZ2v66fMwjYFEhQVi28nJzzuRtVB+yIEiYQqMlFJ9+hu
ITXs2ODUTHCEI3tRZDQImhnzaoGXu3ZP1k0XhKuq69vV9X98RwyVP8E4VWUwOmPM
dlEsQZvvcHM+ILBgX6AVhgZ9jfghJRxz5z+UACbpb3bYELytjYMxSiXwvKq0dvI8
kjp/uUZ8cY/p3nIdxtk/EF9aP1geM1hpGuwfXnD9AU6T18P/dsjui3/v4gGbJuWF
HyY0L0VMViB2YxwjRNoSs0x4DkuV+zqhiPHfuRP+7ff/idJgSciF0wFf6sfvJc8F
Wx79yfrNoTPhmXCaU0mO5lw88KY66XqPusSSujS5T8R4+nXcyPA94gtkGsfymxXi
0hc0LnkT6t+bwLFqBiCojpKWkodzayJP/pGs1LO0PnykPr3iw8FD5DG0WOA5jZnJ
6Idm999Mi8QT8ByMiiR8Pos5VDO0ICxjxeg3ETPOiw4EdJwIkApiTUrWVQFHe+hf
axHV2kPsnrJXsYfCLQ06nb9cL83azcTM4RQcZ1S2adwSZxf5F4YkqEtMn2Yetcf3
R1H/uP1mgWJIXuOFKmz928tZmIqKiCRf4XATVWxBHibpe1jxqokLTs6UHOBxsm2D
/uQ6uFhmUotIr32puoobkIyVmgANRbvxk8cV6AzWxKJTSkqHYGNcmGOYkq8SzDAD
IQCNZSy2Wf5ZTmK4dffTHOkEkgkRTfLi8bsVgAocAVK/1OVvmX524KQp/3yzb8aI
omc6J5ZU8gwRvWL3aTV6TIh2iJr/5ZXPXw4l6VNhy1Zg6+7r5cPxW572giph76rl
JRk+bSnHyAlwJxCJpFpHcftHg8aIf3yT1X5PmQxyV2b7cssSDUcxmhuyIwHRz515
/ci9ymGmjcR3Sn5sjCe+x1qrjTzWRmvivIAv5UN6Q9RUGkw24Jm5MpDWnAJ0Sm+U
XVZQXIFJj3pK6OjAV4Ingdj+uVXQ1Be+3VtMgRIDLnNPCETvt749O2KGFI9smUus
FxNk1qUzW72nwi1V9zrGh7mCWfL8sG/UF/HapnZjqI0lkBBBLiTAbpKHTGI0Qdcj
QlDmkLILCOU/Ajih5BbeXPm/j97sQtlpg3cGbWAPuVDMCZz7EZH0Vz4TDWs9E2FI
hgOInc+DRGrMx0qNHOgvlXErPQfsWVCVVedinbvtjRZmak6ksKwkNAl9pUeiwGJh
s+aZT5PaFRzlm5VCNEgf9eSiwGLc2DJVQPYjgH0w+SSw0Y3gcn2UcKd3GY+Exvk5
yQca6QOCDycobrjVwSmq3bCYQRZb3JQsDkHf5HxoSefl/tSKBZNhHZImkNnM29uT
fHhuxLeTtErAkaxEJjK7G/feIfNG5p1Y4Oume4K+6Do+6YcqaWgNLcENMtD+NIOC
fPa9u9j03Px6mzoJ2m8SPaw79PT4un5aqrFXYjxHN+a5krfN/i2TdFgMKqz1R2en
6j4IcQ+smVKPzJqOjgCJ3ViGJrnqFybAdvCrPZVpZU1qRzURw33tHf3gR4y3IC/F
M41x1DVoT4sr177fisEbazvygVjoItikQdG9RDddlFy6GHxgWvcnN9skjMwBGPq6
pQwWpFG0+Q5VxJK6QEV6HuU4QoPX44APzkVYlS9vYJGGxc6UULrgWYF8801D5iT1
7CqzHNaJY4z++fktcms+Jio4auaN6dSxxPcLfFbDl7825HRNtGwuMqxOVfS28TDG
4ZEuBhNSugUidadjFiICFA8Vtca4zQQYMEfAYoKo4wpxvkGnbS36IGk9rB9DAfQS
IS5Redvl6R9VJYPbiU7hak4nSSZC88jCZrYsvXiMaTCA/BtQ0sV9W4XtNiWZR1NM
3XQWDudRiZWfd6TdkHDzXLzsJLeOU2yfw9qDZ5++DW00/zQBbyVxNKUThGPA+ekf
OGwPqqTqCy3oPDvXkLLUazzy1rlygqqw5AUesF8DXUhGL01y/CeJYamg0xX8cUCW
esHkzUN57TCPDx9qSsJglObLuHzLpGfwRFQGPqIdGr/zi1sm9yum3cbfwcSRzKpB
r/UqWhCAFiRo/Cd8v923iftKPfW93in8SZBapGIZCgmnzxPtfHIr1l0wnxs1fcot
Q0SVmxWD6oE7hj2F7wwwtORzHFoRxNtlhtduKIEY3zHiWcvtBdv6MU35eJLvEKHd
/Vd4CNXa2ocKm1xpKWgdc2G250Ce6uWhwDTStFnYBo1QE+uP7ViaHz7vv64lk2f6
gNb7270Lx1lehbeTbZcle7Ov9Eh8cWrUdItwH6exQ6gEPz+V8zsloluUjeytH2Yy
fFAA8JLzOi5g64Jn3ZXT1BLh5vsoWukWcpcsR2X3HvD5+kvbaaUI2jXI+fLSGfmo
csI3X1VRPSiMkOiIY0Garc6uCizn22DiVO658fFrkPTR4slmPtn69AKfsO3qRDuc
pkO6LCo2cDshPZ5BeTD/J593d2ogwXpMH81keLXthlSMu2EVz20jqPRIJu/5Ukug
SDnAENXhXcowWZjDbr1LYIfhjpFjnnVWoasznyk+S9PBTTJy/XiYhHXTTAgSIuuB
0aJj2unm4AIDcgYtJuMSpgkyJ62F2qmBSx7jjvLVRpf9v3mAiKSdSZE2U2BXbS+U
R3caiSnzGSpQxAxhY4C6eqLghJtXuKgesfCgL6SaHWW/HOLMdXhaNgyYRH1WQy98
UeKVeSv08v7hbgXbo8ooMXH7fgaNbdZfyzvAQ8Rp4PlQn3EpdKrAtCY854uylIaV
rVdBaVzn3CW8tG/hWxM7O01eEQ+lj7wuaMPJMInzQJbkipwDHzs7SB0No3g7QyvP
f+mQv8vfF2yTEc+OZYTBD74NDGj09u5YAuu6uKMBGITZywwSEX8VDhmwzsMgzLv6
9ix4HrpQfb2Ft8hMhX1vOWnaw98clR6dHnK51nZA6sMbRgTihe+oY87MLA1AZI+L
r9wdNKkG0bDy2i0B1dlIYXrQ4EBh1OyCO9rhrCMrSX1IQ3wMmaku4S4XzS+M9Tt7
gwuaYq/pB2sgq3aKc7SLEdbBAXnBbot0F5CMr5Mzk8fMy4Hy+47F87K83Ymm6Dhx
CoYm/ZrssCl5IZ0oVWsYnDlUvMHaRkuUEG9ZzV48KSp5IrZu0z4GhGLXhMqTjJCv
7EUIEQVZS6phJClSxSlY5s4GbNZITr0D51cgxs6mNZ+GTm5U+5a0bmQrlot+mvZJ
xzUom9nLu1cbY1QveULUcUhYarZZvjuNQvx9udmL0RSRJ796UXsqG57+ASO1/AMC
qHKOf09zDhIuTyFAtMgHmRyp6e2P5gVANpl2DQPDHPqwr7GAOOhnK3O8k5w99Dyl
YF+3nlw7iJIVCoM4pZbs6DHx6JWi4HjuoxKXdtromFs6ERLi1+H/b+D5jruH4Qat
4RQ/ZyZDtcB5i/uoaToWGH7KjLdp+A4aPTbeV6Nu2OEJNQmCf7VrPhv0I2pdvgqF
49ijZ2AE5oCfSN4rhrXEwKqnU+VeMczCJJZVrhAwTfxKnRbyPRFflth4NN5GFGt0
/RR7aCHj34xkO/0K8grk1PQf+CxtVvy176/+WGs/0adWtVJSK+ONWNft8ALUGSwX
izeyhWTk0HXzVtw/Fgjd7tWmhGq28PFA7IefYQCeqLDmGc4JnnHPtmIfSy5huOVY
QOjBzF9OeHjE+AOiToB9LYm3MKe2voZH942BL6Eus/utbC0C518ev853XdOw7ILr
VCxuYcTdXrqmv0LrYlMb+Q4fM9GWGJuLNgARvMdb1t2qn5RJvYZ764huRvm1vCxi
0ATG4ql/XR7U9o8jMyY566Eel8IOgtOu5/xZNN9GkmXcFXrHSsqRvrfw6mghxLV8
Sb/nNBqu6YhLBhLyRUrfgnayBliRhddBj/wz6qqPNyaIrSiVCjAEltDFxNdT9Uv5
R3mgL1yQUtlTpq+ISQtpU/D8zW4bg05vv7VZD4Vn0GQCSfqpjW/BNJFKQSsEerbU
EZwBISz0jfI2s1xJAdTSF80bRHhU0IEkK6zVKpZ3V1SUtS6b7mJWUVoPaqgPAalw
bnamS96+1oc2IjQUMIV6vSE0GVwYok3GuFDRWKA1zOgEeFtuxWO+P+IuAZAVn6Hh
a51hd6O/Iv5Rr1fXUd0PAgsTKgrTehiirBHey7+RYyn1GETX+x21g+s5DDVKXrOc
OSu4NZsQA5QvrYjv3m5TUub9B45QXLk4vPcA7XY4+2wa+xa5lk1kDpaUQJh2iIdd
T6Nx7vA3bVHuFOCVuvGXKBxDp+RWP+beJzrWlT8dxq2tJC+fk6H7BAthL3gFyFB8
29JsDRH8UXZl+q/4VxpNwcwTxnyRXMB041OfHqgLdlIx+oo5uQ0WtbP1NrGXu7sn
7IozbL+7X1ceQ01BMLtNNv2aDfoil/IB6dDZJezKuqN1YFitDYNQzkKJ9VcKwbDE
vrbLXEy3+/7hpS5Cjp2JZH9mnWa+qjApi1nUWIU4EfvFrSqBDJ5ZhspMabH1X11w
EYG4PQqpyOoigmN8SUwBnSW0kngIpqKtZcJdXn/N5goC8IYHTWoxfqDO0ucRYTPm
fYXCHtiIrfrrasa2H7McBeqv98sbb9Zm1Xn7PDFmNF6RXEaNB+xejDZcemhxFPTp
x6yIFIp2p0nejUQihx3TqTv0+4FS8/+JKxi9SSpUT1ws9qCffScD/dnT2EMUeHL7
hCLOB5V3p1elFMBKxMKLZOHgES28yShjD0+HKlECDJZ7Emx7pDJgKsosJYCrvBGC
MyDJefjBdB1Yk4MR7lRPWYtW+lWFSqAdOU7PlXySbGqU7+kj99lSQa9/rMXSNOua
W+PG20EPkOOdDrnzj86sHVek7gUN0lfnMEAFP0EFuPvwr6tV4QCwBOGVIfOxj1V5
7ok3NtMES6PnG9DgxBml6K13y3eeKZTzGd3HR/cKkyOJ7WLfbw4t/WYS4wr1d2mn
y31yDVkRClnBpwbwpSwXte5Cb+wip2Wz6bMQJe+V4BVG+ORWZKIlHFWgC7ENPsPi
suW4Z0zeQFwurhA61f9DKgR6lv9js205FrKi23uCCBJZl1yG558zWDAnktHwsvEt
vDGNas2ltLNwxB6Yb5vQKXzEqo3UUJlOZAxaPVN8UmL/vdkaYvH/DE8qTMSQvPo0
JuCAsCRg/vyGQlpe/qk7kLraSUGd5g9klqzderD6FwuRlLp98hwpYVlClLHQtmuP
V//Y7XkLwztkmgwq7QUSrx0rBjGYdvzAepgIUmTQhud/Nz8K3jRxvLJCQaZkvRvM
0qfNpc6J6IH8r1r1NbAZHiX7ZhOE57bHzDOHaaH8rE6CVrnYcypCA1HsC2K2rhdm
uLn+n7c/Fpxa5oF76A5+IedWgzZIrvFWbX+ccb6/M1M9nElGZfUGyFwZEfXj0XIw
uWPekkZY0Ys7NqZ5J9TJwASj7IqsR2uASMwxrACH8eRelfI5H/H/7xMNmpWVc1yp
dJ9MbmQDXNCdB7kyhA8ZEhZZdPRoaTjA4VsDHW9MqP7li71neZC9RF1wpInqwopd
3Ub17gEwbO6vlNuiJvLtW0ELJySVBGDfCGatcYpvA/bJRxja1FQ5cxkf5hJsM1pT
dMZQVodnboZntdqKicq/T4ToNcHMS2CTyIozRJ49jYQt7yTQWVxJAip6PfcJS54R
0evqOdqyaSUu6a5chpVLfhjJqTEsWaG3GgZXEQMMbZs0Gn7TdO/vL1XktZuv4Hg3
xaeDt9FZfi2MOV5iLtL+KYKnCb4CbHsvf0OdU01FgjqBLP9fh/e1JE2P7IjiJO/w
zuGTU0Cmzp6eG9rLuKYUg6nP1V7DeHK7evRuNWXWKwkbEDvK2jtl/sHnWc3zvQHG
TmbVFBKuLLSPzb+erAB60pMH+/Uzvlu+RhUn2mPoVXkdUhK6BHRU9f7yhAM9lBy1
7I8ENseqIwAvBpZszeAobAc1Tx8+F8UJofd/uKKEYUKdc6G91EdwUhLi32SSeCyn
A5uQUlf7y5iD8HoxhrNOf9RotrfkgFbaAgpmB46OsR1KuVq4GUCvsMiTf14Zr7MW
omF1NWkiIg37nAnZiV9eCUra8pcjCHZohj4694vRkZV27iE8FDiUfGwcAiPLe02D
xTKENo92VvB5Y5e3fTCCgbqN5CG4iDLxUMBakfAObadF7z2czDdXE7SmtBZshY7U
D7Kydpq12Jjn+HhnYyOD9SaK56kcMN43beNHC73EFfWg7K5rWz7HTaZlnaqbr89v
M5sbWe81Am9P/v15ebtC6MjoRkTBBP9Duq1qEeLEyNGgak7iBC6yiKyCxvuMj6bp
q7F1aFqd1V8NypPqV5ZTDgNRSOkkx5JZeC0z1kfd7t8k5EJb7CZQCacVZykL8We+
GNnCm9t6suxtd11/5WPcEMGETa+HaU5ZfaK2zldmzP9ckqDRNYeFZUYlZHWKNbsl
rk5taGQWl5RztyE3A9R7Ikhgkr/8ow+6bHLN9R3DtdoZxh8yxcWpw0uZsqIKD3eA
cwVQ4IePyY1CX3mLpDPdfX6AUokglEt9C0lFxyNpopsIisEIdf3Fe6K4y+s7niHD
Kiy0CCjRLnunA4hihEotsolzodDQL1mN5KeivlT2/sK0Zv3eqGnCndqDKoVRn7zA
SXo5D6+JV18wkGj35IeSuw1J74mU03zTyahH2w86bmztnWlkGMqE6GNYcFP3S0D6
giqof5chip22/fYes5QAtGAALcbr/mwPiu0vFwqC9jzfhbJp3x9Rh3dip09WcLl0
RwEFIbkCZcA+c9M+FfITKabpDoYqzPEifWAtJy1v0hIiuTFz7tGSCkpQ1Z5jAXnV
dBXFyE0wspTVXg1+f2WdtaVApH2stFnc9UONWSyk6EzRxvPH7TcewMICEkjD3Ksf
fGnlQBqeQkAhEs/dgn7rpXeGQ3PfHwjdE2DwpE7sIC5eq0g8vkOi1O9uSJzWA4UZ
p8YazN/S2HKreiY2aMqeVOAB8mu7jUy+PYv16P2h+tj7ax2v1MKzPi+mGWRB31Vd
6AcRzu/KMNDMYBtoVWMkpr2dbjNiTfqgwuEIB6bWqB4C836twMX9E9XbYLVDti+Q
fORUgBWFeh/fc1QaKtxZgkhAjQiKBHdmNHQ+5XtfMeFNFZOomCQ8cYZbDOJvQrap
UpLpRm9XKwR9HLt6kg2F7UYwytsxyaYwy73jlJ4jBFEDOYYqCmrjk8UaaSNKMK/b
3QSFqNq+G0FLZDFvoz5WyoPDL5nyXv9Ttq5g/5Gb/pSasUSAYpFMAFXDjT2Dh9Ji
nzAy1hEXergQAzLQCXxphZk06qAiyCPpvz1VnlAoQyBJAk4DXAISQVEAMdBe5Eq9
NGGPZ1EVQ3bE4k8E1aisoSVE0n25+jutQ6B8y+MbwlHyK0H3XBqvb4xbnr7z3vzg
LQq83MYP8DeTAIB/+QaTxCk5w9KFXFYXYn0F7yFzLZYJUAzbEdbeZCj2jiPefGb8
MqwwLWNoWBoY10nWa/B2FEEPaMrQbTO7DDe54YoU5wKU4vfM3+3aS6KT2pUUQr4Z
ZLZp/EXMoEQdUuchHl6gCRzWnbnyL5vw+N/VU3Pdsp4EJFqJuZJaKEvTBcWN7AtW
ICl7b44HWMGfvkh+/5KePh4p7YQP5f2cCawbywaAH9hrZDGHQ9LOjGZBMMs7uMBe
LhYY0FQ6HqdCL6+oFy0wbhpqsd1A8W2ryD4oVKqgd5HkpRTTW+tZFBTS4AsPLljy
7j3soLdvP+/tbysAgwcU6Czo3G+49JYrilFi4r4NiPurtYtsGQHdoIon1O5e/yu1
lpxmUXnPeLDvEqX2FfoHAldvBfgzesJn8XUisqsNeP29GNNOhkeiYUBft+1/L/dO
OTp2TzqSlTvRHGTBm9LxzkXPUmYzSCTtmgDoUzoT2cKGmHBb8pRzYjX91jTa+J79
YRxuCn10sw4vD7OS+4xOx8d/CzLoPDcFUQLSfYTvlmSRvxbwuMURtL9ZQcYizIaL
HNuYDB/1k/wRvx7TFCG7UnglWuSxzPX36OqSonqG01eaZ7KsW89pBBltoiJP4kMi
BjW3q8IjYhsMr8PcBkURC5/vRaXJ0jZq+csYJ7vvT8io/bnUXv19jTUSiuyVzWGX
grEdNhJ24evnB9hnD0KKALDun6UDmIxdGEKx4RNxhtlZbk6hOeaCVFxZReaEBlk5
C8zDlzPK7NePfZpRW2OzMcQOBoP9Xkqvqzct1CVdzdWxjxGYuOW5ElxcNte4dFMY
/za2jofobfgVyUjBwOTg+VasiCrt7hD+JpFUvopf2C368dzHOBIcuHqplgfd9SIP
DMSKYUjyjsbszLbzMEkiz4Y7RBmP8iuHs1HmUDky65oX/SgjAiEucAdEQDcZW5m7
YwHgI3qY6jsNxpt9r09IrszdckPlvdfWc+ESq9Y3tv8IYWF1ldwVsyNiwGGejkfN
X4yRDmXaXP4yxLSnZATxgwn9fuANH2IvJrAxqkKaQpjdQiYLW0GzUSAbuM8+8j7C
A/186VNXYpp5E3it+MH7XolpI87WMw5Rt+kMjw72ad3Kz0tlIfm6pZ5uNg4/P3kz
OFoS0Z4SB0UwNR8Jh5S6fKO2+dEBDOiLVlH1udg3MJuIsvm4JHwQSC21oDhZeYpq
1dmiSbA044J4AkY5/fbcmN9gGJ9+7RH79Zb46cbR2E7HtL9zAg3JonrgvTCCFEcC
xyu70gcmetSE10YGBA3KGFH+C1VisPCYRqy90EYVNc/uGawDZ+5N5WNy4NoQka1d
bW6AKZyxXwz1WpLTXEQ+YpFgPKmMaBTTPaU74qG2f0l6u3g5tEMklUzAHXcB3lgX
8Asng+YsDOH1oJKeMTJncRHSk/Bs8tsZD0sK9ZuaCpF/Opj65rA42J/6QnsTMA1X
noyraF9UxmFCrczB3w2q1YZVBwRs9RD3bvDppXo5O6qJMlvajWD0jXGbaT1TTldT
/dbvQS/v8H7UjCXZXVxn70bVw6T82AuU+abkfQIxBLQoYwnGn+YH7H+udonyHviw
J22Q7wmHr79hSjF2JBb04tmy46IRbm9p9dmL2ILadDGoPPkuiW1hHd4bgU6iXF5C
84ntqpPZ4Ep13GMRyNdjIjntNtzkCdWJAwVlvnGoyfzvlM7jSsr0UTKRaeVvycof
7+fY3N6YXUCrtEmGDMRe4qOI56glYyk2541OC5Da3ZVZa9TVPtW1hlHjnLpGrFeN
8PKhdHTU9kvH2PGsx8OaBlVUMp/3fc8csBhAhTPeJFjd/kDjvkAwNt8oArzrbBqV
r11jAvHen5yCKDgZtF0FLpKcSErFwId8TOOguW0vaPxPQCaoPUYmnV00dwImI+po
l6QbXAd8euTxPZfmdLFxvvOTgXH88pJQs5qQGjiUJu+V7UEgdB5I8YsFX/WFq/HS
uYIGQg0FJRnNtTKsV0RuS80Gny1poqJ14Pj3WjyseUgYuneEoyYjhEH7uXB1GCRA
psBIkSrxiZvQN7LBoqvmuRe09L3NN2KXBwKlKccgDP8ECYj2cvdG9xUceVnipMJn
nH97rcmkYANSygXuJTDkBPhMi1jFsj4BURqu2UclqDI3Xd7irA3YLpvtyslIFHEq
1tDimzEFgGBg7te93ehnAOy4Y2fELkvGYX3MGyf0pZrPXTEXp26k+wIxOf0nPU5o
WhdunOxba9xsAGuGuAh3sDTdhdFtL2YIofikVqvsgkVOcZLVKPqRITj51+XEnT6r
QYVu8sXnaat2V6YEaSCF4FKa7l0mvrfAm/hMY4mwRaZ6E0Z7rHW86LW7l3zBrrI8
w2EXwk3FsAQYmxdyaTN0mQd+GffTkbGr2OaljOI3pnoYjcNHz3iHhr4tyj0+Cmjo
NajIlttN1f6o1HrvSHIbth92VXpZ1PlwnDBoXBReIiEmTsfOI61kVGftC253dqiK
m6OX+ngj07HbavTNBokXSg0RH5sCTqHi2HFjAMuYVSPDWeX3oLwtaObJfmBOkJgZ
Y2mBNDkQTZ1vgkuFiBx9TwWQW5EOBhWZwIzIqzyurb1HN5k/mXgZeqj2Ys6OE45h
am8u0dV5knQmSLp+sJiBb2ciPuu/0T+qxzMTLrOMBVqVH+BSXr8meik5oZEA8+8u
fpzJjvlMXAScWimjvw8JgmdGTibl6zeCtKx+gU+79nv2ENmoqqkKANXBFbOt2V2Y
V0KRds0erlraY1EBTKYZX3cxksiZ6NsmI4E2Ig8L2PCIt/STb1+rFnA1btaUqOBS
ym2WaCGnsnXeFSYXvxnRnGhV7vVpuM1wpZ6nd6reX2BPO3LE74JKdFfUNTUEMNVM
aZF813Bm+YCG8rIdGJV+auaVBAmRQjlInulGQsUwpm6HO1u+wqVv87jv1dwfPc2L
hK5/Ppd279fmY3Cixo1SozgKrjhSgVYG6oh3usK/bvx4dgasFxf7oOG8x11t0ANe
+4hulzq6hAH5r5UqdwCkGSGbT6g8NqYgt0BcL4SsZyKPzsGjvObVDwe+lDTLbik6
6iBiACC3rMpL3S348q3whOxYgDqgeeyP9J04VYN11UaFNnSgMzZPGN6rwfRX3197
AtZ52D7poe2Vw4rhD59d7Xna1NaRRRdZ8zqdpRZ9sHd8XFmSjdxHeseOQa7vhUUI
/GWQ1VTVM3x0SZefR133E3q93wFmCoM8T29Wnak2k3MZeUy12QNDaAwoRTYktDmT
rpTTvbFt6OSlTdsXU8VsYYVWWFq/Gj5mdbAQFjwYQz8m8NaDQSwiIn6iVgySXihC
hJfOH4/lnH9G7oujMGo97O2+Mn3r6TF1/kDG7LL3rXMvZ30G7B6w8qtbmRr0dIkc
qeORHc7CyEEWKF+fdiuH7Cq6HLsccXxV2F1WWF6t0y7eXVmypW6Ntidseycq7VZ8
5XwJTqXrUgbZ6mqp++Ji3lB4g/8gdKmz+ZNSb9ecROLnxyaeLF/tp9J3WutQvTbA
3tS4oCCMYzTt2gfaYzqIM526PMTvQE7Gp6p1mTKe1ID0Rk1sJZMX5PsiEokwasNP
8vivtBwBBmH/e2NUCN/y9ooMuxh9DtbGvUtMyVyUHknZWrjLmbBQxNbmGPLScR6z
UCrdwpUzE8ClnjkKdobFhH+mnHQgqZNW+ZyadpG4w2tp59Z1OfGqC2xswHB8qEn8
zikZH/x+fp7Iz5Mtj3JtCI/WP2qkLeB1X506T5WAx6lHOBV0W/Xg1E6/FIb4H7os
vtMgKCwuPIuIK8VCgRIw8gLLsByOYIVkqgxa7gGoyFVZMeMBhNmaB2EEK94jBWah
4dlPbt9tTBhSsbRwW+O7wp4BcErbwnAbYTIC60kAAysNPs7WfpSDZ6rdJ+z611NC
ylGWybik8LrKUG2uMl37a/xC3KMdB5lDG6s+coVRmcoPd4zdTYbcPez9bs5iSlX2
DWxoeVePZL4ZGnP3UavOx6MYyOSyy9P79FBX/wDTUldo68Qe2mFzGp7+UXDXMEdF
08fKqpLtgOULyqwhBau0skLRqV8+t3EfQaPIb8D1eR8hutQhgJU+1B8ms5gFmKr8
XiAvx2q55BOqHUWUwHypREtDU9/AZuj6NnQ7QUjG3mlHMbsv0Q991uMe3BvGCHQm
y6u1RYhTPw1lHdQbqpkxlqbwsxVr+l5C3TgMg5p+J/xcGomHx1McraeAPk1WqkuK
Hn0jNY9iE2CBesvZ6VyUkHxcKrSImHCeAcR+bQZjSVp2lODTBwT3vNiQB2gpFMRF
7ZBSJKoarpsPLdxx5StQ70C5zdu7BNxsj4JDOKeu6XAxKe0NAuUepTkgneyJHaR2
oSZba/flVLmgaHsne1nGgaMuYFCWG0SR6min/YOQcEuJtCKm4eG/PvtDpEjAVVqF
lao4ozdbUqq3qWpgNWPVP3Y4iYVV7Qa4kPb/en7hqiRE+CzXSlntxeiMHvnTjEFX
g7l60F4FxarkNs4w9D8NtR+PlNmihI9GUW0al2cC0z0TD7qRCxJD313c6prHP4kZ
2ZltyV9MC4iZPcjc2U9gHJqnhby1czDcAubtymGEbjgXcWBIsvPTiZIb9nBPBuOZ
EA1rLVUL922KvvzQIpjlqK6mIHnSNeLXtyJGD4yA2Mx97vmh9WG9spwmlzM3yAMG
aSN9FU3EwMDvqILuT79s+hSCL8Yq+RYEIpGJbn2X/ppAnUAi8PV1oULGXLhYU+x9
7WdocDOGwnAYj23FByWWPLCXaXHO6rxXO+MmVlluZKAI1Nbg2HY/KPuCtOuCq3kS
Ru1SANv4Vew04Y9rL0EX18+b5BMigNOKwHF2JNwrjIqfiQ08G2b5OceB4FwzsyLu
rsKNc2I2FBhfz4nze8Ar5IDJwhd0dq1DslIWar3jUj9GCBtQk45BtySuGkFqhWc8
DZ7Ar5JirFhGpVf2+EP5wzScRPn0gjqb0EUUulhBcYddP1JJvMIG+Dts3Tu3zlUn
AGBTkmpdfnrjctR9waQuFvhiwwpGUrkve/FT8C4hZVnMjMnlvYgeGvwcFzdpTXHh
HtoxMMMNZsRLhO+Lsb9F5uQSguGfeYvESJtCKU1jwPKeEzgQCZ0lO7CfdJLgoyfd
76Gl8rYn7/+9z3exFIkpDtPlhUvkaaciC6vlFx2gd0vBwaPOdgax2LyIvBTeI0QG
dLhJ7SRUVZvggB4GBJrzknCv2aTFohqZgmUJqlLxV0fhEE0vZFe1f4VmKQC+Zf+e
x7hE0BurbY8rk/RZqVXDRjgqt8T9VAlpV/c9eU56i0vmM3o1XF8E0QITwVvCY4LL
PXYxn+5AmqjCQgdDP7XS6z6cjdgFtRUW1m8w83+UZZ78D7GeG/oSQu0BWsUr6PP9
FC/n4E4xTqACaU9ayQnB8KAjHMIzQafugYMoOggCUM6/ZQMwbcTlBcOYYrZZd2rG
ME2EB2AyEEAxh6JgPRGFyojNe4RqgVERsjRno6oJ0nsFU9c5a7QR9sT2ppmC/1Ik
Zn8erccKjsDhnx3qbkkohZ3sw89kIBJY+gSeWDcCrsEM+LPbmfNQCeelVpDvIys5
fGdGDMOLAXdx3WtT+l66v+h5uppAaUlaiR45N7wJp3NoJIAJtspyPDYb4gpyfxFM
obiuqnra7byh5dB39NqWBZsR1RnyH2Krh7YiVwkBNCKdvOmc174piw0NduXVcDOD
/+w0tcwSqbwg3GHBLS1IQyS276SYaYICqMHDtvhMDwUQCVX6IriYbnziUC8ZlP7j
cOSgwVyJDELrnaYvoatDUp8dSnCs9I5xP+6yllQ9k5XVwlc36YVJiCNkuccOlcIB
v5uK9H66PF0Yi1Dn694/hR5qrtQPuICrk2lsvTua/tAsOQtU6g7E8/Oui/UeZWKe
Ay0ClTk70WFVg+ot2w5HSlasWSLO7uXCL5IeIlRqTUy1JMZecUdKrsk69G53yG0e
L7IJym9XF8lUvMmKMMbXhIa8mRcDKZmHO25NplR8R5Zl8vXtrfNLvXH5orSY+YhT
QuTFMtxyafrPsWTQgXm4i4rablmVWJIcGbBlQtpssyGstAklVMgtx81eAxTzIIL3
wqTtZ17WspSWuJh98wfKjgou6brtU8wGs0kxWoMP3GZD7/rfamOsaWCkDXmulzoS
J+DDS2B1oMzzsVWlmidqK+0lyOxLy5+iRM7EMYajwI+rbQ5dTPARzTJxWbmABhEU
cqoHPJ9gnbBr44k/OZbW3LVeFDSz0fTmn0v6iKIDonnEBDwS4aM/uRnDDCfUpyqL
cyXUf9c8c39+u6gnEzcqEQj5JnQE+s5UyNHSqV9smaUBKntzt0Ba2DwDAvV0NpKX
uP8H9wrlWmKHqvJLKPdAhod8sH3F0Q+IOixmyKvLRyQuFne4/TwjPuRq5B/Wa/2w
PB/aMPbs7i40u71OzLjt+VGsW+SxIpcu+SMXlBOmXEMzLPQG9bae4hSS1qJRX6CI
tego15/Hp7q/Vqe7iZs6rSN3v7bg/DZGMyRrOhdYUOqTfAKrghyL9+DGgfvQtdKy
R9fBbM1hNlOEPg9B3xPf+EXgXUKs9I5Olh8r1it904YauD6bIoqP870n8u4dpEZ2
1koI8X/Ux8oba8o1Jz+6cj5rTUb/jzydKX24a90LekI8x3C3vq4OONhe+nJXe7vt
6gPqkqciVhEpQP+Up37HWwNFDpWm1jncFGCYU54WpyvDkdMtfIesAHY0BEespbLF
5WG4QK7er+WvGmJSlKGXle4P9Z3AJGEC74VR9fqqGYomU+dnseIOJzn+uapffPb4
fwgsuDkpSOwyV82/OkbImIqDLHPOqzDEbWIp6U4vBrOdORxoZesflMoLcgOrk7vh
V0c2QdhLqEC97EkVyXK+SX1HlHihkh6hn3dDYsbyaJG/MGlphjocaaNxWPxZIs0Y
CmUse2GzBs5d+UAsUlLqWOj3FdcUDbn8jkEkLiGGjN/4e9Laq6Fb3W1RhbG1WxMQ
jpRL3qawsCtNvqY4hlXUdgoWIHFqplFg9gEBaQ1bU7mb+9+mYMAyGFoK0uiDqSCg
Uwvtq6R4gijWNcLCZQZHefO7zdmhvCDubdIo+HVCvmtAP14ET5J3V6jjZZmzNFCj
qEyostCGOBAeu34h3OBYu/0h4/vJj1Ks9DBcJBIa1B9ur0iAG91N1gnAmWhxJEsn
k9Dqr96LRps0ACVykf6a1dQNnGRA6lY+X9zBiZw0GjzJnHlUM4jhwH3Iicgk8PUa
Pq4gFhiiViOLG1FFymViM+b45aClNHfC60/NTB44Pfvnr5TC0rabJQquUkv4FDPG
pL4i6HHgu7OpYVlThp9sfhng2P7GKubJt+xIaYS9qZR2EAFKDDjkdjriOcYRH3/6
m6VbRGx/Ym3G0XGKXCbRl6DPKRJgAviVXuMHrfD8kmzYQXD8u8s2rwRzrfynjDVA
/ThcQb9dlJQDzwJSQxBE8VN2NgzxP1ddJwz5hsQ67m0hnIeme4QaEj1vzowUXmnq
7QSFK6hP/2ei0bxPOEhwlNkrwiE/6FidusgqdSr33ppzf8h2k8SiA5nXMnzGePyC
0xdaPifUeiFLaA5H28XUqcc/pwUqQRoxYFbnrwH7nnjhVUz50iEU36tvKnWzjaLi
CLCZxMXGFvvuoN22BJzrauBorvjIYsm0ZjTL+Kucm7Dlrr6vRkMpVUdm6V/rI60E
RuX9g7AVV8yWjta84lTcSNf4LVFqwVxNUhW3f7xURyKoTPtQe+Uskm41aXaP3JaS
cxJ5AvRdY2SJJXcrvkym/xu1WAWs507qV5PNrE4x7ra4DcK7wlzBRW5h9o/BKBJb
UDCoFARc+aobvbm0hK0B7iY9/qcMMNvEKAClDNxfPavBoRULDQ6scKiLSNlpLGre
Pg7NewKyw8jBXM0zSJSD4cpOgXLeuj7D+KWo8sZUSDN1I8gg1Pu4ugwGmNuF9r2t
GQrHn7rEFlRMwIjdV8fZ911tjmGpHdmXByk+XRkD1fdh2IrUPRBGmJ8vCYfZRKWw
sjqn6UBxqurnPmOi+kecmtxSEbV6g6eriyVlTcYFbs6OmU6UM/14Wd9ilyZEMeOL
zMHdecgDEYoYzfwJjO0r6/lwHxO+fzlN+nnbFc66B5IoZfLfa6ssXOSbwfpx5Gu9
QCMQlti5WaYWU7dlqQHW7NBJ06dUm9tWkqsK9TECOx8qGwBrnnNUKnWpU9Zz8RqZ
dRXYgiztKADbv03EvN3rt8IQ3f43s+fFNlUL/yNOtSkuPb/SoDhRCyR2nyXbTPMv
4XXFpOy3uKfd8aBAUrW2xidotZxTwZgZjeXypTD3Kwt/VyeLlLJEjHOfwyThp4Lp
a9XWV95G/Jj9oS34rpAI/KaK9gNk8Ac8u+MlNYUmdRlnVLy6SNXR3uEfenJITAg+
H7ABXC849EPzBkPs38d0vsVEj/aK0EawaLQwCebO37wPmLECUr+qWPHPKp3QkCNq
+10/mosqPJXKuz+Tn9caLnfxcpRy6c9tDJ3oA0xqLu3tC5yqwn0r/kevpeGCRNqs
mM6dR6udChPYwUgu1D4xUNuyfTShbO5TjfPZrSr3DeIZb+OjRwtnPuyXDtNDWb+R
jKU7bnVbCbvvfxewuZPsplwhb4cvDd5McVJktMp5tOzDeUsYIZV93GtOQ+9cgcBq
ST7IMH9GzuopLL1UyU4tAdA6wxvt9vCTYzoOS8HUrJKKU0FPjcRqPYnQocL3orAe
ojIzHsvTVaDxwYhwZ270ua9ah52LvMMI5qCGzx+Iih6mULuIH/GLERqQYPbg+kJU
tOaC9+geZ4o3dU2+49oT1SEBMsNTcuyIfaGEgqQl7r1DruR1lKRUt9g4TTHKjpla
LJ/6sFn7Rj2RtXwXRkD+DEkdDRh3zNCkYDNkL2GHajOZuJSmwPd8k2EbnRRCirjp
/+HrHYDWAHzSONT79RiXAkf0KNpOXJRfY2G6XYRmoJQaDNK6SRl8Zp6Cdi16PK9c
SRMDHXqEPc6dZsOuCwujMbKD6VtNGYc3SOwptNl1zwpilIoK68qVeScf5Ht+lbpx
bz8bsOeCpH2SljWaWi79TkVYFllgQrQk/GQMqhrARzTWnSkBi3vWQZHRbzBydgyc
vfyzSAmk4h9AqiURBXr+5/+ZUe7Nr4xv2f3P+pRA2t+xvHvsCXl8wUk2r8IYKkOB
3B06co4GsSoSiQ8x+mFChT+GNiXo6AzuV6ZIZGYNEP2PuDpzyj6N0BJHXryjKHE3
jGkvZ/bNpr6rWBEOCrJS4Abq0SJpvwtMB5PrwgHryI3udMF1wP8vEwJBnk1ZaSu5
2KrGgrEJONV1S1l/yNiIYmZMQBBU23lIdizpabVZ6gqJxtjQQLRgX0UgbNWsVII5
ucyoUpzzmlPw/bHJc2+CwvAH0wlFY/9Bn2s7RlV5m1YfIJ9K1gOGZrpfTiOsTlyI
gFD2o1WeyFj2jcANKIGlMNLiiHCceDV6/2qNIlBsi/OpmjxhgC7KGebH3ORm+BcM
2ifm0DZJOTiHgwlSroda5wQTj2GNng68oAHPlXP/l8Sk/SC1yENIUZYPF9Gf088z
xSGBoMMlSzxGukDoYXZjjVwtbfNH0KtTpda+p68klSbUhbUul7QwEp1J9oK9HZd2
uQBe53uUWNU+rp9E4QN+Q6lhS2NlqOOVX/hjYX5rh4AknGisQaoVb5I2tTKL6Sx1
jyFjSNDAW88e+85U9V3DjJxu9qW6i5bev5MUVdBx0xTy7IrzsWC0PBxFZ4ydBW0s
0ClI3P4iafp+mURZuio7CZDF2pqPZ+NxgKweKLSPmlehYcgOKYkf7PJU7WRrLqyE
5PFW+67jSd2ELciBTsgClr1+UiUB75NcDwE1WbEKt751AIlm8iz0ukygIvGFCOfa
FJOq62xGxpGDCFkc3RAQbK4q4Xr5vydHEpcAHerTxhCjYBlj11YjErUfMtRh3Wsm
53BwlPM0A3TP7cmOjWxXqdWAZXREXUJlQvHpuSpfyHifYfxgmd2tZ5XQSnbl0iN3
W32yC2WWgIn9ll2jSLpHYTdQC8Nh7KEoog6RpKWysyiagcoo6ykoK028S/nCm7ep
s63HBBrf9My0WT8EP5223BLS6lkysEBHN33IKbIsFPwkSu8aEAc6K2Ye1eg8WGm4
AZLqv0EpgpIyEROAwyKcaToDVc73mo17dcC9LL+Xk7nzH3swLOv2G7G/RBo9lKMP
X6T5o+wjm83C9xTbAetHGQO3w1HQMp3IpyGeRPa2n5TVQqb0j2jMQiGebTpGtL41
ry0P3YgUOPE/R4of9hCHhDCM9tU7mY63MlYvbxIzUX/TDQDOdamBVYb63F1iUXf1
spyiIGTOiMNxrxrzLKeuSyuqb2nxl+2WtpngDYCojXFhej+4D+PsfibWxBTpwV8T
kLVd+Ll+o85TNt5J7AyAS/w4u3jB1gigEBkJCX59m2bC9lGexPv2vIUr1Vqq1hnb
WWbXAM5gU0WqqCZBiS3bth6u0Py26yupDOIrCxdjwRZZ9TQKLoi9izgJPFQ/05bl
YhYvD1WyaWaLTKsesCuB2BhYJIkoju8eU+EZnkczXUEh/Bub01fDlI+QSMIr2cJZ
gVFIXEEHHSSfJnhPYd3NQYj53nj4FPbtJak9cbwAqvZ0GMcISddj9N4zPTrDlIFW
p/ksegOb53blExy1i9vgyJ0LvhtL6ZTAjgHZmFjd5L/Mg7z9TbHETa4X2I3/BuOq
rWfn2gfILf9TWw2czT3zFlw+wMHncnF3GKP1Qa3irBVVqbRlvZVWAIixcwZTyZ1V
+TE6PTJ4J9RFhqYsXzm49UT+KvFowtwCvC3xmAuYHPMJ3HA29Bm1BoiZnQSSAsRS
fDjJ73B5O11+29TNtJd3SUzQfogfl05ywqvoqmm1sY/g7o5ogQ9uoxz6uzHAwdhx
l8jJXuFW+NPBY90wBO7riQt2kPtSolXclyEl0DSrQ12R8qYY2wL+Txpd7EZxBN09
2vZUscAa+41bMqQW+PHaU5aqtqdKVXTH6uJcHEzD4GUjPmAG7vAcvBrG0+IJ1T2y
ZchJNQwxfo6nmCpvLAfgMmiFcd+OOoYbDZakomhZp8vLgRpkeJw7ZaDuel9DcpKn
94ZvULVu43E7S9bqBwhYRSBE7QQSAo0QBu1ZNUnn/9yFsQp5wqtusowyUrPPn4Y9
WXRvKEKxVw8k3TQ4pcRhRfxGujOrRYoRdBCMnGQ6cXwsAfhjfXDaco8kMt6G2eNX
e2lk8sS/dHgrS1VU60X9bjkZ3RntUFDOeFDF4b7tZLfie6ABuSO2tycPOedV7kso
8K0WDG5j1KzXfot/3Gca5HLA/sCgmrjLCbNLkSSvzgJIa1mrIFuLrVgSEKL2qmKk
Jqmuzg1zv3tT5fiaiLFTu9P0rLRAINXYj1KiGngLRDh0o/ji+OfVN6VGGlY9ecl8
OtCY1B0U0nWRWGY52Mnuh1qQV0IDFm1dJ2czAwBy6xzzfuH+On6NkRqqiG8SlTVx
GoHLAl82GXEG9OdFXhqVu1b6ml1kEx5BmP18dt9t+3Kj8N7KK5yNzSxU6YiN79Py
q+o0HJU0OjtDsy1qO5JsHDE2XTrXreCLWeGQdErQBMwtR/k+F2aZc/4EVP8+EHp2
Dw5HRyfu/RWXmZM/JpRzWGb87oYOJPb2FRswd82jXkvA7LNkqXdGagMonRC7gb/d
CQZAoapPPig+x44Dhce5C1+VWreoUTVwW4TLdJQM3aCJyusNMkBpyxZPRn7y1Lda
JAR0+CMC/tqVau9rfT5g00hFHy3yZjOG08Oo3Eu8F7+Z7zaVsn8UuH7jQk1cj9MA
AkylYL/D9WAacD+Ss5gTY0ht+nZac+ythlMX/8wpbk53rhCbEoQh5+ceu59K5oWs
GuJexqPJd3j7hZBN60QIJ77SEgBYFB2NOGVvOW3Pu5/Xg9QeCMroueNtv39hC+27
Ci0QGYgyIjVca9MtDFOPXMH7JahtB+PukQ1aMBoqyvtXDnlbYizebt/y/Yh4a+6f
g7dlZrtGu4hfvp5/lUlQPd83FWJPxmr0KjycbwGtP3La+j8KLXydV02E6h7IfweY
I9BKPKUuAUvTpLw2w4KhCWtsr/BMKn00LU1ygYFZH59OWdfPf+2IvwKqZfjHts+1
AXRVxwgCNtfFIBrhMgpmEMJKmBZ5E/cjfx+NTdrg2orU6RoTBd8KAGnFrU/m6VZp
aPXlbBXSE8n2LztbRnKBJvOhsGZE5JISTaVtzRvTfIjsPEASmWV6UHnd6vhuOcxX
qKiaM3FVKb8SiAlvKrN40WnL+c60sU1zFs+IsVUzGDEFpg/tpJMkCIYT9rADhWQu
2mgbQ2igCRgLrkNTZ+H5wWWf82R4xPaDSGIexafNSFYHrze+4411oJLtlmYFc8bg
6lQLoUDTLBhshtFHV9CEXeEcPRVDdPWYTC4my/b7XF7f/w4bddKLkIofoz23GQqX
wPzJaNqlMzP/LlAGTGGrxiovBbqSJGvGiHTC5NUoX6TtZVqCWrdhRliNOfNwjrWs
cjaGI77TgM/xzA3e2sGbRMa+lEo7sIrDZM5GbjGq5lCLYQk9BndRCNKeH81ZBCU4
9vLkt8l+mL7AdFHJ2iSOXIvJGJo3iVPFO0qRNTfsvypvQNpL2HPqgIENqQwg+AYn
F3OG/tgh3wuomDLkh0KCIZSGYiNIdhiPJNfH40IO+B67q2vfU0A5alYIme+prwXQ
dIZbFId86CZ6s5mhPTKEHC8PBnG74TaLpw7FP9VLMud7PtJ47qb5EJJBelJrXcs+
J6RHsS5m+KSv2zq2bqFhC3t/rEm2gWrtFQse4hYf/UuxIycPiGcEHFO3nreNht7L
5nd9JKueWGmre/1jHM+ESjbsS3tkSjJCsVs0fX/qFfeDoNljoFgvqRRJo55di7+N
wHTcwCNmI9l5qW1EEjMGjZqI4PCWjwsOIaTxMTKG3g3Tliys2tAu5gc5iGRFk8jJ
duR3EiTvwR7AMwOWC8GfDjPR+6rrA5A8GeNAtvsrge7KaNXyjn5TAa9BYmqxsuPm
48xr5azubHGuDaGmAkT68tSw9K74BMjMVBUs6vTZspsNsLf9shJRcbjOb6xJtKLG
xX6mioUusrp/wnb+allo/OLRjm2S6LacuvJ/RYuNIF0hEjg5vzDjcDsyPmb3xUkk
2KJfk7f8k8bOGQHTvSYX1erPgunrLFN62rWz5Z6ChiGsg5OU2Tyi8kU0SeZW578f
jZDvas+UuxHsGlISSaHxKd2wMJjRB+lEEtekMJO2bS+hoTJl+qL2mE7tKIftmBSM
XgWYlCISNdoZbmgWSI7LPz5HLMVtmqA314nF9BpRApf0OHhpi2V496EHams5XDHJ
1VBs7cMTea4/c89RoGPQK7GkZuk2TBz+b83HNMvzA7asYKe8V7JZAKrNqjBfaP2m
OkmF7Dchlzhbu1/8k5A3QcXSv0TCCighcl7ote71476w2V3M7dLmZI1rJQsjXI0C
KOMReaj5d0bVa/5H/IFSHA5Qe7thMIKc8NXuKOU16+pjPYRxnoY2AP/FJxEyvyee
O6sdL+bgqEIUyjQKvOYhPclsvCV9rDgb7BeFHOBpQ4+AmrFy2yEYYiwy72XonjVG
y3BPi+8pbNNDM+YL69/P8QO8fUuqJNXbj0aKhBmB4wCuJOCK/0mK5H6sIptehF7P
8Op/Stho9VGwhADN7HP8k5nIE3vaa8YO4IRbBE8d7Wb23IJY2HL10VCycgOhtZT0
UhW/tBKNHlSuWlHVapLDh06H+M3e9Ehfyp1a6ghS386xpht9jlJtLOdn+IBQ0VQL
xTC8VEnRWCOll2Gkwe2/h4Xe1iqUTGc6Ov2g61CkzqO40MJDmjuIAN4rA7m8vmtd
lqJrR3U2SKs3OmsYMrK0Fn4x8M8kVIUGocqv4vwlSb77bV6u3ihIK6MyTdb6ykGY
cGymd675zBn7NZxyY9g9yUZjuL77MbJ67Uj6ZJ8CuGBe6ly4RNk96yBNYpWjvSh+
wecZydWfhZlzLjAo4ihoweGx/8bok2MRdIun3pABOT1UJgWlZGsViWn3rHqNtp2r
zITPL80xyJdKxkY1Gye6o3tD5c46CcvZVDWVAa/Li8TqIZi0LOBiwKseZxiL+5qa
cGQXQhJVgiMixsKGWgXZ+2J2NaL5Kl6qHFOo0R5RdHBhgF1l2i5o+RvIW9J8aRFg
eI2J2WIK2OEsbSECCraOuA496ZCLcjNrPGS77MgAV0XbNmdMSerZT8izN2eWniR4
5FIQQ7poZ0INY8SPCJfBQIAyp4XI0alWA6GHSAWGeYVmurQXZhjpZD7mttDVqlpR
RQdhH5QJyVkffmfCglWkiOpWBAvi6tIBzwHhDc2ZtpRQQU/xEYL5Vc5LxK7YBCbu
nmkfEMBjGPl6swEQAYdnEpuFH1BLajPoDN6NHjvmyfKxfr6QpE7N3Po+hjco/knI
B7gFUHDVU94quZEFG1/51QfKAnXXDNBR/ZhURMw9cZgwxwbomhg01/I+8ALZsu6B
6CcOfv4WWqmTKStewn8NimpmHbvvxJ9HHp2mHeq26kCxM0kYCGkBTtSPIiUqds4I
i/dn7HaDZW7Guz95XPnhHGZZX7jyN9ZESaze9BZ9SYKkvnkycgHA4H6eyy4uOhUg
wjwLMmnjB7fuvFtdj2ZwOpOlybb8xi+HYCtTjB+65mqRpbLn0MyfUGpLORtqUXRQ
UxZyKRmC3DigB+8L1Jwu7G3+eWwMR5kpiGSeIo4Lr3wMZon5bBj43JPcN4zrWnta
J9amKXVDGsUW9IpuUG0hjG5+iivecMcMsioTNvzOJyg/Ts3uNUoyjMsxHKr2N3pf
/chPlapP7d6OdA+d046L/8z2G0wztuTbAue57cAZfNAiuAbYuWctQ4/07xshhsEk
WAfoEtm9KhB9UfGCxIrflBHoG4DbdVNWz0km+7ShVRbGYUTZ4JCEQpaUcaE8ghwx
NltAp8QpcvmCUvDuIIk/UpaMW5FsWppA+yOc4S6yOZth+Q4zYizupvWziGyHyrQW
Gs5VUaJMt41PSbtHq1ibNZvyETrV+8rlktk4SuLgL9mn9+76OsWtuF2AH5zlOd38
RNL/AeG78x1PWl4K1a5R+RarQf0YrIezE5ebp29sz/EL5D0utPRPnq3K1lAQUNQB
/7ys+MAGCrhbnGJvz9hNIwXr6qiybncoHT3AfcqxxJHNEOrhp3eu2SHUd/fmpKtb
spAaM9WRGr0ENGl8+omR1MNmwyVrvG51uQ6PM5KMRK6LXVF3JA99QnoD3DeOncMF
lqijb9bivZP8nxMLVEHhD+CC+agHdTP/O8yYW+Cy0tL5/duy+dvRk/rkZGAuhqUA
PvLjMRolw6GyLoqIR2WsrTB103MfjgEISiU3GmsvQtFusB4kcjrajKN0o6a189Qg
wkD0mw2LHmhxOR0bejRPY/1Pj3dsvFbPkqAvsRweLn7ukJX2F2Vox0nTaNsJuPs/
FLAUhaUpKbEz6M5zs8xOEFqjbJ5CTaM5tCIT0JFWqIgBZndniDsxbGYY9IgmPrL8
5AqZ8CjLFglRQOGJEygMnjBc2yM5meDbjrdvcuxWpXMrfZOqIDtXWuqRo1axXB+j
gWtFk9Wo45G44dz4WPIMzPTcPE1MixN3SnGaxLyHDQjct9vC2bGCO0bb61Iy4E28
Tr4zvScaBywlOeqUww8zn11D6nrJ6fSJ8S6YiKykI6czw82jjrB/jJjPUjapfW52
nqZ5xXnxn1TJz5N4Jc/Vpn+JANUmBsss/Iqa/T4Cl/788zDa9REXORYVucJBZvlx
b7g3QqvEvE9OxOJCSx/Oyg0S961Fitwht3KEQzA4s1BE9jcvIoixMt0+z2HOVLvn
XD8sGTvDvzufLDmlnMsg2tXsCtYYdwQ7yUf0GaRLqtt/XcP89CZcWv7tkYnwikQb
2ghquswqQWz1Z++BqVOlmzgf9/Zn02n+D7wBRCah4V8Zt7wG9jZirZBvfpFvNXiv
Lp3hkxgY7NhdRo1ZpzPq1Aaavkh5CwhYVdEaLjgDtxTWTWefBXEzyxf4Omaa/mUr
kfcz346NSCK0IfMf9djFnZ+GDOwpISpacqoYiW/dFXg0coLPzNtwU49Zo1q/QO3a
8GUKI4jukrUwvXguCmy6rlcx00zf7PR/T12UohaGRl1PrU25o4Ma7NSYMUfpIQ7n
IYTcLUwDu59Ld54h36WQuRn6NabUEpQ1+UQXtqVrzTrriKygtFoVAHRABpZM2WHC
+zNud3EE1K0osm8v7nVVh/z+kd9D/xyKm0Yns5siMX8tOkiDST6x9arqiJ6P0txu
1vYQQ8qmOhtGe/oBWELFg0IVvtan1wDR3qgTWtqMgaGdeAxj8Qya1QvQUishN8jo
gW0kx/lJdllXHxPiNf57+Geax8BlpDqo/fBzKq/HvNLqlTb2Q25YT00zfm/1jZcr
tQw+q8IbJ1eejByeDPMvT54cgUktWEnp0s81li+tEgttzfuV9NWn4cq9lnVLUTNM
wWds1hRV/AHTce2Q1x8E87CPMW7ZNO6FNxSc1L2Fif0e+20Uhmc2akIGIa0xm8Km
DBwDQhXCqROETajDC/yTXXllT8d3rqpuJ76Y05xAyNC8ZbJCA3Xec5bI3Q+4ANKB
FbMaeGlZ0piXnYt7GAUEIxopbYBZQ8WKYwfQjPhi9At3ACMj0vNMSVQjNE7BUf8a
tgFyOLkVMtNtYZQeeu+FbnXDMA+4PbGZc4JABpvktcXiM1ieE0+nNrLqJqmRJweD
BLb8ktrD+rmgbcJB2uhI/5tpWt9Rrv9mFq3LUxWSjwdtnEbVvM9792MnHRiCDIHd
6AirPUbM4uILlg9MWU99Fm8cDegY6mLD4SK5373QHeyhmCphn9fY15a78r4awRH+
Mrw8pC973sk9SrVAliFDyTce+BmTVSFvYWStur5TJSIFmphYB6B/RidV7gnN1gqP
QqYJ6swfLEqa4mC72Jkc7HoENXgkajzgLKtDuohFEnAoyK7ml5ri1kRbNbpMoxxT
a+mQ4MyqpySQ2i0uvBsQfsX6ND7YlrwbnUF7tus5XEx1wik6FNhytZIU7uOWhul1
rqTPEAXQ8V1+wPXuwhMs+E+nOMvPTxSE9GMv3Munh1EW2bj4EYfX3+vRdM9AsQ4o
wDbdRisub7o7uzkraWBFg6ErFX71m78lq2mUk8UjwhGY8SY+ezAq6zJ17tvkJeye
4Ra/OAnWHBbH3ZaXRXiNhq5yC6fIL5VSx5ubq3B71wNuJWzoLfnEcWnS6Z8nt8BO
V/4KTIVMLs8KozuSGxgdI/DO/upR6tjexX/6CF+9OOv0i+H5hLOrqjzLRf84/CA5
dXk+Wiv/2WfsnRxEpXMgFcuuIVYUEgDzMr7jOXZ6bxRSuKaldjHKt4Bb3ppPxXJh
DVuyzvtT+sh+Xl4VJMhFcv1JR8VqJVfUA71/3W3TA0c9kIk/jnGMjnbcf2iIT/A5
iCIWN1oRr50UZP3p1YsiMCMt9arm1Yt1ETgw5/cArLjejuXTKWCajuaVJNiqnrG9
BA4bJ+uCjIhvMnkMi1k8j+4TqS+5jF9VETZ3zJ5je+4Gp27opBmwu2Vngsi3I+TI
kEZJg0bkl5s5+madfk97FWQR9wSMUJTvNPvjSeFwFk/nA/kFsF9xrzR284Mr67tS
ZJF8W3/aUDEPEKyTepxuPKQM4Pp+mDn09Pz8t/ifv2EUS7Vj+XaN0duLJsR9YcIc
6mudyAZFoQGayOsHLGxskdzYx4tRbh4rBZI+aZkRtAxce+G2WM6qYwAoC0CQHY3A
nxCEoCdsY/Z28v5P3AZFgodL5MsQ4Lqra1VIYvL7sGhvIB5GrEI+VnqBtljPi394
miiaFvg2eDbyv3q17nYg4HTGxBzWGbaoomVjqXQ8mEykZOpK1cbYKIDHt6zl6S2q
/tJo1xCmm9NC8KrphMhG6uxet8b10lo2g+aq1nM05k3MPdZydvVndozYCux5bBIG
tB3eJy427r1wa0Ucj4MBXo1pIz56PeD5fMQ0u94sLeOVgPsGFnZV92XpK1Cx1q+N
RNBWYhmrZGpXdW3jGZXZ/bnk6jikTIn5X/UpJB6tt93JZasObzTbF8NfF/2bQ5SQ
y8n4mVAEo1zjs80EGN/vvbu7oxChDXsDyIHIVfTrWv6AmelIWigz9Ca0aJ2XlELF
YCvvHMB/aAJ6VUHb5y6NJfwf21+fGSFd1LM0hPKVS8VgVOHCDFGjk/mu8v+Fv3UW
hLLlK7+GN4gCh59VqA3aPxOOh/LqjgdWmQ1ciDDcAR5/ieN8PGNbNR+0/fVrv2H6
p0LwcfzY4k/nV1Ilta42a7PviA+Fy8Ul0dt2F251dfsO6Qg/PXCwcNAlpmBkCumf
B4DwCjGMu4bFLf1cXyCf4K9UJixo1hiUpy8PvbRoYRavyqhAQEEYC3SG4gNhoV77
Eg986KbIQ2dv1xPvqLylea92sjTSMSPPEawQUCGTruHn2/QckYL1KfDKoQbP5twT
2jlvMOq+S0MrHVE4pvk2s/pK29Vn9ZPSufm6fPwf03BOGs6AbYoCMqAFtlah6Z4s
QecC526tdUZlImCjNj6YSApssmYDsXqcjEgrDoCrOk54QOA2RCKKSvsDnSPNIwSP
fGloTrFvKbKPpKG/J2br7UzgUD3ozBGOwSrZSUYs/j5k8W8hbgvy7lG4fC9o0N+D
QGgN/TIhlLpUWyVxYOi5pAn9ZzLXioOOq22RN4h0RkklZSuZuHR2hay0x6m5Qef6
xKdt055qk0wQmPkdNPoq1g+RPGNrdnmiIfDZDIekU/JSGyW65UhoxMWc5RVbLzea
/5+o9vLYseEE9eYYjWdZ0r2mc7ONLVSndV00yNXISJq0QC7QupM9bHTO0UNmraqq
I5kklE1ZG9yeTkma6E8M4pdmM3We6YlBUrNk5EgrUxz04kfNnJFz3kaKX/b+m3wZ
NpwE1896Br1PpmNKHrRKfQ4vCc3qf7aJD/OIRkfIkT5npf89Jw0Td7Z1348rnOl9
dcVSKW0tbHORqI6rFJ1LT8KqQJpEFn+cOxvJmx4ZTZkXUe3ukiadbJobqB9LW6qB
2wfHrTncW8KdPtPEjqYX6rpNmHABaHiwmbvP3n6eOXTsqh6KWU7OSJoKyRqUCE5G
SFUd6LTqEuJHyjLc4Z54ov4eAoG8BcsHwO09TqJCe467qZkf5LtZbtK6473PCTXC
z5xlzB258tqCJN9bqJ21tTOsXE/QdFp9LJ7yLjpJ/NY2A2434pd49t3Tl2nrp6u+
BXs6q3TlrS47yV+B226uAPaj5J51i0uTIg8YbWyGej0aNoS6iXoAdLN6KFa5ijcP
AUn/cIfrCPy0qMTRqANowB1hJxWu/76Ev205vEH4E9Pc4SYeIDtT4hWfU3SyuaYe
kQrGYnHO+aUoLL9TkxWFED1HzmI6fdhkYRJz0ClpvWk76Mz5n17gegW9pw8DGVDn
H7ysRcj/Nv45czxlFP+KyABnLI9cqlodIucyQ3DUwoVI50EdW84eXo8rkzSvyfL3
TZpPHN0WmeRYOiSICcqr8tgiAd2DlL6gOTXLoqgxNCh/WBTSBChR+NnMxrOQOf2a
QRR0OyrbnfYYl6Yjy+pV9zBH52PwDsSiRMNAhOWkloqX7A2CrL0UwIFZ4rH2Huf9
vVpcQiJ1jWcxF107sDT+dLcTH4JaB8Q2E3BCkSB/kYRiWEUHFsW0en6G3I96mQAu
GaNb/vmDm3JjiF/WE4x7vWVSzY+nU59j6MyghKRsS/fDeji9MRiZLeYFgPJ/SPxv
EEZgCwsljAhLuPC08bVcmNksjIwbRkBgVfkpqKp1hB9+TpbUeFY/pSEIpHxHLOEg
nPeQnG66PmXXgkf0a4CVld+oi6iD6PR+xWXNNl5fRwkT/nlR7JJvRqmPb/66CF8d
xoc9nV06JfkNHyV55u94xHABM06NDqCTD5azDeIRqFn1/XvP69iqG3KhKhtJOcNy
YCzOZKfQwKxY4NfmSLNCpTDZuSuEb6HndbKMF0W107F9qLkwD/vdGFuPAscEVqWL
1WY434LD+WozGmQJedm8P7IdVta1Li9iixoaF2VviR+1WdJgjCBDm0E6UdeaQvPv
Jhsj2FkfBOSHQ28JQ5IYi9UgL8p/Yt1O71w8yAuJTvA6UdeN03cWa3BBSJHiiEYB
aTE4GzESz2gVv4nnjds/yvyRmKx9sOOheCKiQRFUb4+5r8mPk0aZFD3G6smUPOaA
8Pb+MkECpI7cidxZKcB+J8sov0yhUUg84vG77c7b90iNYOvFM+NAHrhIh2RXOHTK
pUAxozsX7av5UDI2DyGybTHABCcOZ2iEf8upn+c/aWjiAbiJAsOIYHvnLukdTyGt
3yD5AfU4h+DgUSS68HWQ90iNCCisHctvv8Ly+8dCQej5u+Ht1cAznujzfK679UC/
UkDU8q/b6Bi4zm4sCpvB2Kj8ZYo6Zv2Two280NJhTOq+JUkCLUk49ekwDo0rTUkJ
mJUZuk52dbyXgTV0tI8ikbwoMxYDz7g3NuwkzSpijJ+TLk/9hX/YH5mUZ/ykgqPe
gydwRBf/KaHMVxeqxOaC4y3SLTCFT8mz/m9vKzleIJre7XOvIaArIl0O0MypqTsg
wyxOytAmTiYcCQZZv084gS2XjPj8tl3rIWYGWXnaCXOuRFR0jin6ozFoBWtXAz6j
CK6rV4e+xfAkkNT+QOAwkpllP0kL0Dqy5wHgyMGJucKY3QJ7zQO7VBeRArjZlcGB
/Zgi0oin5P4x73oKyQq8u+LYjRVNGpTOzz4ZgUsGyNqyXsgDN+sbhiUigwmIrx/c
TsUDcFGg4U8eMxvKM7DALezrebFxNCFfEylcgi+4lXDQ21AXVOk+slYxq8n8jYCm
WglthKvHFGNNPimvmv+I1eWevLm9D4heUudpx7Vl+h9w7D3mUjmuXzCwS0brvxS6
0tToPC8zeFm0DFKmJmAAt4IUmJUAKJIKK844irZ+vJ6uMjF7Cw5Aoiohy3O9asqJ
ygxeNo/0JNlY1rzIZYeZwfri0FsA5YnWd2eik9f6O2clzpJAdlh/pklzQmtBrbU9
dVYHARo+kFLH74DJda7HXKdqXlrTKNziCXOUJu65XxV64Dur3u5dx9uemPPqnvOP
cT/8QFaZxTgOcj2jGmlAonVD2iEFyJ2Ti49VS5+lRv2b7wDbkcuZc1iO1Cabjw3T
iKHsrSKMxSjD31Mcb8mkbAVYS8ndk0RuflyKDwhTiTDxvRHkAENjOXsd0Shtawwj
VHh9GLo3auu7bTxBr+Sjl8QO5bCaMtyw0XOjtq7NNx6NHlkZ7cNELc86R20yvYcq
hQiSQ28JKXAXgLk5iICV2C2p/3R43Xb9fRpDpC7NfNq5OGCs/5RZKxFJlDtF1rTa
28JEN4xaCHz3ahJtg2LZBvKB9pltwt9bCqJDHVNfEjbCOmeeBP1IxBv/hvkxdQvU
4/HpS5/G+HjBQzG9/kvglEbQEjV8fX05jeWC0gPb1LnW4QtcbYci2thobL6AhptD
j6lYifB49ceSVG6x2O8ol9//S6Fr3zFm0YzvsSN9TDhROEAEYF9y7wrtb/1uNvYt
+Pu6BE0jzNBTPMiWwEIk5ay0dqWX2TDdNwhacTGxZiBYKID0KFmRsyWHzZU+G1Cy
MkdWoj9eEVRx/H5JXEwMpP/WSkLD8P2qnL8xp3PDequhpQ+D9Q7Q+BlmPIPAz3g7
qko+xX45PwRLPP8glExqK7KQ860B4ljgWNu/ltJP3s7Xzkuiu8lCvlxLT/nzWjor
nDgrvJi+gtYOAcKCcz+yWfNsc4tlwW8vIpLZsa3xCcECAALICddqOTqkW/0/a4XK
UXGGQUSVeo2tNqx49oyhn7lfyRa66hme5Y35oTiw90mRdOZoDouaiDvluhVbf0Fy
miPuPyVs/IlWLY6HjVKsfN4iiSaAKQJNYJT0qBwPxsyuDA6RAFPisgRVnvJtEZSj
4h2UETQX04SOImDhKAlJEuRmA7pJu3RCJJHwQBi6dO7hf1RN2Kwl116qVUy0hTZD
KB7isgmh+W/87OATjvnIc7AHouVzIaBNjkKK0d1hVzwjoUT02uW6F9/cyTFGczac
eZNuke1cXhBcA5ZIkoXOIL/4tIDQXnVEdnP3mBrdepUwfy8VCCQeCnXCJv/29Cbf
HlszFrExFISM8cxsOVwXuF6cu5f2Ujc0MPJbjtzK5ElBRAYMNbmGsyI2kZpqkOfz
RoHVcLuTLyO2Pko55VHvvbyK+5c6jUWCCkDxc15wWJMoFmi6pI3bdKrm74aJ9Bt3
fkmFSMWRs0nheb1j5hNyc3Gh50pYVWxXr356wWGHTRlfF9DamgMsV/XuivQIrkKD
Cj1FJvlVNB/64iOera/iHPGtVKRSZufceUxRGnlB/ZJu1ch9OcdfT4mISk3niGSs
OUfvO9h393MzFiRjVQ/wr51NmmoXKVWLwxKQS9A3MBWENR0WtDeG/kqwPiEVvZxw
oD3G/RWwHYkjfAvnrxwckB/zolBvLaWDgu2loKp1f+8Ml2Hk7D6Y/LXEbjNW4K8u
tvQq8Nu/PzQxUeR9+7itnFeX2IrjRAQdcLGCLlRIo9WMncANEf2vMRFJ2l0ZLrvj
BNzRxK76+WxA7nZ0EjYZDuTLMGwITEdmyhBVseLJgdi5Lm2tKsEwjvc8auJkj/bA
fiQt4qodf4PJSPCC9dWwLowYMIXMWOLjFu6cbSEpyMNk8lMNJahQ/mvMy5DAX53n
jcjPJ+fVm+T3wrdQE6GqcqB9LSf8wPINOczBIENIZPIkI4c/bhkTTy8raidllWG5
YUT5aE+0Tywgsgq4JlmcP7l7GMmDGY3blWtgbvmAXdDKLKVy7dwjYO1BVL5yySGn
x7+7pxSpDrOl1RCzPeIquwzCBrHQ/OESAQEVQx/Cd7IFX/LgP9T29aD0dpH09lW6
nz39KA2pjhXakHD/zOyGW29Bfsly1ZioINYFxh4+wNHhgPr/CRtc5Ssx/hv+eZVh
AYgDOLC4Hd1yIl+aD9mBq/gePTfyxRZn7ntkhP4xnDxUdgx5ANG54qdjaUU3pnjQ
w864Gd/WvVXGdl/n1gjelF0ypLPaQXzP4pODcFK1IopzpieX6GXTwxsmheOojtjc
Rs87AobHXVkuEUYWbFz4YigCRnrHW8m3xmwieq05bFBqIqMw5bW5YJ/Ooq7umhga
DrtAMV1dOdz4LNu5Rc5NjVBkip56B85VteL6EEiTfy4PG56DtpGIvGhiW2j4W73Z
oP8NViCFPjpECkk7OS59ha3XyerVEAc3t+sjV09ok+PhvbCiNA9XXl1qxDkHS5YE
49brcXmjVK7x6znNs7yVPykPoPKY1k8V/B1MjRsvCVMaBoH+JF8NqOogThgdRSTA
MXUt4/m+mDAc9Hp6+wXNE/aX0d4kkatQt0pUiEDx42kQD4kdJ/FBOGbk2yvMI1Gg
ffKkgAEyA/Udim/sHiSR020ruPGiTjE9Ots1s2V/pcbBxFVZvXPB8UcxIeryWEmu
Epen59xOeVXhEIzZ8h9xIFmkPgpWn0g/h+3w62Cs/cqgfMwgcpXuujVSVRigm2TF
GIloMInGRgHu6zLN1kpJGYvx1FTiF3LrcfvALgdolZuK6NcuiY17YIzMemFrJJF1
iyJ0u2JoBGga6LViOZJLwbQ89TbeCXionhC0sFrB+3ruqmozOUudyw89ZH8dNcW1
FP0QE4MLPyvE05PdhXbL0/BrVjP300QDbpUSCF9R/Z28PpIG14rxUtYBAeml11DE
pc3BGXNsUZ5ki96hQfcRZvqj9PgcQ4AjefScTtDg848P4YvieC4eLasnNF/Oq8Wj
6oiN8P7soNps2kEDYE97zQVEI810+VpYcbc/DlSp60lsnBa3ztiXcB6z2CvW3V4j
KKnnOqYXAKJS1r7+NfRrmlvxRgUTszJi6G1Ax0fuwEmc792Hy3JDP55pW4WiNdLy
QSWqFT2OP7eOREYxUC6aPULVblCFm5t4t3ht7cZ2/gv8ra2oIHl14ycTPenTPMYo
jshHbpQ2g2o20R5tuxGpfSgskPAAK30SPdb9sj/iQ13cMLV9KE7tqNmNErRXUw2K
QXctZRKWqZJYyCoo8UtCRGZEm7fhvCw5lkY8skUgVTCPV5PmLKG2qyYrbSwJGsgE
9bMHbFMonQYEHt31vAV+aBKhvlp8v38N2lPjI3+72QuL1briOljy6ZxMKqtYsQVw
4kRbvR22vpBhkGq7gry+XC201SdMlwdfWM34FUWxmBvWLQmz+L0XqIxfBHhpYnk1
Msr50KjWLww4l/3wRcSa6YWoJF7j9k6bmT7/uJng+leey4gzFqHvPhtAEfFtO8i+
QVnuDfmLE+QGP68NmoNSsyhKZ71r4CVnOyeYu8Rtu785E/eED8txPZJ4mQS4vAs4
HFJybo9dL0aDNohiDwrp38aYciqdjJ3L7IRjq/qFWDIF/8Vl5xlgJJ1a9JYVulTr
UyGcoWmdPvzZQVXzyYpZDYWbBuVwN54PTCmds1P465HX17REUrlitBX8bwMbI5Y+
CPDWu+xN+4c/ntg9+4nHzXeDLR62S8kpPaeCwaZlqvJA4qJFfJQfSODr6uOMvw/H
dyqnHc2K73HwWdShE2sKmH+h57YTm8DHP4ZPqP6jPe0KYTNtEwWJgmPveAVYuZcY
0k8/11YVzOrJDOQrU9gssUWPw1K9nLi+FKw1ZU2hiYxeFrcBZ5Pl37zjWib5Nprb
KT5ksPbSL49lJWlba1CO2qBqCwZ9szly2iMx3qTQQbQwa4uyhYoqb1e+9gEM8UrM
E9cS8CFoVVRzmf/4iWLiZry9mxv/1z1dxN+1k86APIqhpkmXA/qByaTsDdh/pEXY
BRqaKcMbsfHEiMcSnWeoIFQ9gY4qLw/+vk7egFktlLVJgmIY5PXK3kFtIpwlwtVs
ICUEDn9ZgyBJYouy6okh0s/3mveyTK3XgtH1fSpm87dUAzoDstiSQNfYg7pR/mpP
hgd/2dWJJO7TF9VOkOeAZ5C1L8+0mFVZnfmi5uJiLD1fOYIS+wASXmFLkIxOOn9S
QEtS9lKtH9HJ27foqtpNdwieNgT1FAUMrbNRBSjFBgV6ml7BAw7PjE0fWuKJHhLi
8vM+vet39H8tH7cwJkDefp2WEXuIJYU1x/WltCx5HgtN7YNA7AVGJuAfOjK737L3
lHyzgvVeUbTrRpFt4UIUo2g+LhjBGo1S5Zbhb0MGeXOIFPkUCtCiQXS4GB8zIA9J
Cy75pk0kVdX6IW+p2COeIJM58BE5wmZfYsVECtaoUqDzkXuzVMcJGWX95x11hhRu
0Whzl2oXr5mtG8mFOaJs2E6zKETzAxBPwxBwlHEHJsi9v8i17GUe6NinsK8B7Lh/
YZ6KbgXNrMT22h6UeXl5o69cURI6DzPA9dkOrNbCSDh9kK61/pO7G+JnQokYZ4DB
D644FazrXfs92GMwHgDS5k9r7Ymjaq74tLb+xtR5Enfl4vdvCYqHxWDwZ1zsKURu
qaBGGqgyMNNrZ55ayd2DcV/NpVDAulCs73PbUww7prKLlZh/f2lmDJhyVqtUXV/E
0awOh7ed8tD5tBXOplWPlQDkNX2okYAPJUdUhNQ4nHxJA4Z1Iyfc7S1NDMW4frCQ
fzMZO49iGJgN2g3O/e9P6JIDEyhnl5MQMk+rwWAqcXvjv4L3BtXPl74wIpnmRYuZ
4r9qB1k+iBAytSOgZjITirRgIHGBk2ym+kRduD4quMszJps3RIsLTSu7OfPXUK7d
Y2FSi9SFEzPsV+UkKVIh7YW1QFPz+uB9ROSmK1WJPfiqGr/gQIxw7JkaLTHl6EPT
82t/p1t2AbzHaDHrgLiijKKJ+UhUtmcqffGNCsaDwcK2VIarSokpMiktzLGOgW7S
zqxkc0HIJ0K0lIf3E6HEb9PT8tDqnXcqjbclsIbIsr/L7Z/rnVVsJE9vl9MFx+La
zISvL6bb3BdCtng2hCkQXyCMlPzhJRIaYLrFVAeYUC21K267fDH0yvyxfX6LFsF8
cMp0pL6/Tfm7DGoDAyyJpNY2zn0LFHf86uKB92igLgiUAAtYxbZDVCxjXxodkJtN
qJcmkLg0JUF0I3scT3KGHIGN+8FFBycY92hfBT6qexA57aC37ESi/SxmQLxe64F8
yDstzZh8HS514y/+SuiVVpk07koBho8tl5R68g9HqB623gHR8QM2nrkqaLL6Ir2q
DQ1iT3P4gegwfzmxAWefwamUFeOrz7sO7zjVCR6GawjT4KOdIK+n4MhUcV80pbEb
E1DCD9P5k0SkbNd86GVTQhsuGL0MQ28eJyPgetSVpH4T0C14hy46KpzWJG6+lcWP
3MXrYF/CKdCv9hvn2UHOFknGv9Qwk5yhUrtgUXYIpQ5CQo5NeOo+vaw9BjpwBDyI
HSz1DSEaUAqYBgola+R+/elux0kfmQKBwLmveLKwG4UkxwvdmBKcSbu/2PuLTA5M
xp50v/J5GRoKdc4klWTSUJ4plA0BUvOFVUsBgU/XGRWW1LWkxZanPlLLeSO81Wdx
H/Ef6A6z6V4osjIbpU/ys9VKLf1rizHP7x90qvy+zcZiQuCKGK0dTOdqDEG/UVgl
kPFntMr89/RdKZwKJ6xCbXWvnGHsKR6Fjcvm1OwfIYZaat46rUVHZa/DB4+feRtz
Vr4u7d4vbFOmSzDaS3+x/hSqUBWcSmrBMzjB3tIWRo68J9qcvq3yg6gALYHhst2k
nNy1rJouLzAEDFEb9zNld9n/8H5Pbf+QNFSPeObXD0MkNuZEIznD0fDfXWhiNYff
I7L6DdGGm+wD2CQPS4GvneijKLEZEjfkTmheYr0IV+S63DB2LV6AUEmOYLPqvfZB
/S1PDhJi/ThQgzcKXacSlut4YdCSpHathA98CWlwH/WsFbmq5BKXaRnssxCwc+7I
oPQzGhGVqO4yqmkdqcbAXMZ9lv3zSFsrvBZPauVF1L27uz/LiM/w6YwwUJyCb8Yv
YYJJ6qqvUw5rha0rmf1GFF7vhcX7nRxd9nCwCYooSmMkEkQiwoedbnJ5ba1mnVn1
vg5rSKXzoD1oZhnkX1WfevSicfKMxhRWKh0FOSwsK+QqY/A2t3gWUbudLETn633Q
uvsdoDPmXipZSpPYQN1v7BvMapZEm/XkVMzf1n2JXdawl4wLaM45JxhAHxZ96hCV
ctA8mXxISK38v2iiUJE6ORH47lttS70MrxbHig3/Qp0Qb60QXvjnDmmoD3EiQjf2
EVnc8km/KtKOGifzitGVfQ/2jPg/n+ElYDUGPRL9ZlHBncS+MRVDy9y1DyToN4Mc
18L7LaP6sH+oC5RiP650pzpt6krLcX1t9QMzOed/VP6ZyUaLgBEUCcTDlr5OG0lN
V7981ytPpDh+1I7pntfnto4OAxUqeIo4XvM8zEyamvDoieND4vjJWjYZeTFtMH/Y
x9EUoA3pQhm5/PWFUUzGd+zi2xR+A+pjicUl0OcO9grqTgJVRhYosZkD+uD1Zbj3
UNgDf1uw4Lh/62bjs1wK5HGXZRuxzx8TrS2qMZKii7rln8I7Dw2uskq1m87Pt2RP
sLbgd3AylsWiGUL8LCQEM35mYqdEqFdULoPnrxnsqz1Ddlotal+6gG4HhQajTuSB
YZqITOP+6rj0YSoxuXMZawevNLJRdCGMwRwttbL0Yorf2oT/MyPkRK2QNrSdHKTW
jZueMKq2SnoLi1Qw0VxSbEMhbN5KQqep4ltLR42TaK7XJt/5/ANJaWPkx/g51lui
G0r1kqY2WHzw49o/h09VF7r8dzhHQCDxYwnnBljaSZ5fEv5Tw+beQSPO9tJWHsSk
beQWS3+YasVBcVBreFo8gsq3a5CoVU208YFT2V19tqDuZdazWGCmC2Um98MZQ0V4
dur7nVD1KlZMKOLX/QKajk4Tcab/C/yPuJpf1Rh5jhrvzuwmrMu+uBhA4TLvW3Lh
YNNywn7wND8D2ZMp+w7tO9GcDrCCSjcXPSLwj1ne02XCkweem6hSm1MOa9U3vZIp
MsPY0iaENtCdWRTxk9dD26QyE150Nr+tdaahj+ymLpJcnvPknLUxleC9XNUP724i
PceK/Yczw9mVWQ/e+iZv7vy2UqrvbSqGQkiG9OdwxJSiyialyWsBvhiaghhn1HYU
+6BZMenNuhuUr7nc11C+s8VvDfdLKVHH6i5Wc1zqtes+sTByZs8egpUiP0DSGILd
RYKCxQHoDDVBMZyzLMQFphq+MCBRHgaqqQfiYzy8lCFG1m8sLyPMEZxbJX9buNfH
cjitN1bAF8NXj/3vTDk/IAw2cct+WjsRnNenQzn1tpXJkxfkGaw+ce5EjAN6/Hh3
Mjdbzb5b3o/ycGZxamotlPR0rEezAmssW5bfacd93X91RHbTcp5yBOA6uNjGmJE7
0YZOOh6vcKCN35GPBvzpgi0WYL1QLUWkGK3NSZRlVHcm1VO6E3wYZSXyDMnjmhIW
xWLyp7OCnFl5ydE9wdJEFdUynVQSu9Jnc9uWX87z07TZO6NGl3JpgqxEyyhmb60I
uM4msClGTQ9iZv0QdRAKH2SZsnoH2Zudh6010mOzKIlRCpJdmolln12S8tWkJKc5
VUc0IchIlszBx3no1rgK/ZrFt16cB1ypN9USAPs5ZklRYwMmwkmBeq96YpPS9rnq
3FaSThSrjDNeAnHF5wxNWZHZofklSd6OI+HL+myoH/LzBh2I+M82DxtYkPZF4Wrt
7SImspzAgV4FgSO4GRj35VIiyFHvLMtE8OE46tPGhr6/ZrHazGmjeTikvv5BtZim
2yYl68Z+os5VDixoLwNj36vg4lXsLOZyVC2kMq1niqIwlpVJZaw5p7T566BLwKAC
uIxJfGA61H6mmMROmSljPQhAp8uEY9BPnJUCzaRGaMt2gXSQ7w4rUZ0J+f+YxKpf
i4QnGcv17bh19nJoJusEuXPTuW8XDBGAhj0aYzF+pPRYoRV68hWYPtCxkhKiGGZ+
pLBYnBqxQxc6eUV4zqjBcGrh5oybKN4W9zjXqVseS1ZcK/FlWk1zO90ZtCSDZb/w
RzWak1jgfF/rsGmWoHxh9vS8uUz21O+QHD5jYCBU0F3VTh9eZGdDqVOPnZtHYN7Q
G13EiV0KR7SInW7VBcdWdOLWrlBfu6kmXcE6GFJzOnrEePwUBcfplE4c9CrYHlZy
jsJ3Anv8R7sfykeXnQyfZHmfLrgAQSzqaEe4WYbfP6LA3qmEoutp69rQrlxnIIss
hFH4te3u0T3z54q0TowlL4q+c8VIKNmG4lMlEiim0GlU+ItK++zJJozDqXEGRxKC
fg1vSuzuJcmGb03K7fn2CAvBHIyFhsW7PWATEMWT5R0Pc/9AYU0RWqx+x/NlsKUP
dNdrxVb4+3ll85HL/qadN3+xiGV7SbnzORTDaJIo2qMiHhLMnJQKmmz7t1B/1J8l
oCmMDXmPKnVKsd5jmne75wExMm6gki8i95pJ4GpP/cbPmPyCOu6N7epc1c8UQglS
WrZT3Y1lWAjM7oiXUWRb3qO4G5bWUuivcxvmx9lI+cEGpK47tLz+5aAsbKmaIYtI
mYaCgO4Q31FTCs81kFg/DDZ2QudYGPbg4ublPkPXNnli4608PbE74LQCqjIYc9PU
ARmnO5systNgzs6+0Xy4YvR92tzTYbw9gFqQLVVh4PT18KVju+tLXwX0qS48eEWK
/ah42CNEOhuEXeFqparTVAGkIimxUgnd0ogOH2PJQ/H9pTqR5J+s938W7Y1uxCwM
TDz6AzUEzsNfyXnYp/V3AsL76xx1Zon3Y2qSIQfULkp1O9Vz6TLhboBL+cpZVIbS
u2sISmV7Nv0mduKNJfa19IOMs/vAk0vCet+Oy81YAhx78TDXyN0OhQtnEXhFACfF
fL4RO22zWNwFrsAnwpfsn9bwiZjVrXwpSk9eLDAuvfkCqm0fp2RXB69Jsj13G4m8
poNXJ7104B0fNIMA1Jq6wapJslTVWBM+NsKHIDJ67NxePTz3hp+i38mugBDKsIOV
wUKdpFiNot7fS2pvf/9zfRyf3nlLiKreoB67PGitZNq2aY+ZISCTt8Bccc89AClu
5vNMBRIy3D6q/nULrlewM2VeBsgYtzahKeeAQsX3Q4T1EY7PZJ1cBIkYVMVmptNB
PjyFdA0OIVIDHkbQWk1Mh9u5H32sUjFfsTiAOwRuLX+NZi98dpuWKe4tasEbNiwZ
SC+Tvc0i8A1s0zldsoyN7VeTL2+j9UmJ7Mif/q3xRklwSvGmJqM4vubXARQjXoc+
wgV3OqouRnUIa3iHW5xWHK9OJnrglQbxZLM2wNIxRlOZcFYfiaZ17cKqL7TK8LoY
a9VbVxzrLM3S8YWiS+bUc53KzvkPTmbVrCIic69JuDZGngGfFzx4ZuMkDCE9Ol91
bOMPEBN/eGe4tGP7ArZGLcJhJ1oxLqg3qk3xWlEj3/2nLTvZcWpA7bRcomuDY53y
2de6oJvjpDtv4QPrljPUDugPtdk9KaWEN+js0oDs+QrrgHJKkUwa7eQSTLWOk+Q9
f7U76ujUaW0ne9MaD0i70yUxf2vyp+0ZfWu2PoYbPFHIjTRW1HQ6mNVoIMSfDZW7
UJu3fCjuciGddOCaF9HrNo2U/CcZTYeE6/7m61CoeyD3+BtksBU+o+QdM1jaIUVI
A5LpUzRX2O3cTDq7AtvK4CuCUae1MXj1oi5NSqXmT8QWGpLrP2bhphBNahxfJB+w
rx4UefeWh0U1qoYR96GdeuWQTj2XxqPtw9Q5TV3tRZFWG8YeMf3hdappCRlvNO/a
DmEJe08tAd7AC9OT7JPq3aW8KJg5BXWEwSxxs4MKcrPpV0ueJMIFiOwiydUdv3Nl
OTnBy0ycuDLut8aLEtFczCHXaZXRsb53Kq2QGzgP7mbdqdwIx/xCblaPIyjIWYjB
YrG3lXKTCXQ1isAhvo8XE4JN7p+Z8GNNLfZ+mWV4CvC2p6K4RjugwHywtcaYXNRw
GFXdiucKhEBOaZ3OzRl872c5w0SUl/y/N83yFYDztI2W+M1BCmCpBcY/I0Zvi/zr
7Z/j8qnV8imHuT5OceExZRQ4JpzEKV9PoyMmOk35vYkmGLwQSWA1ESfUVsbZqYCr
F4s7dcS0q0Qtx8kDnbvjbiP4uC9jmSam2wYFtyW7QP+QrUT/nQkg9JwXoI1Bp3Tj
vpl4/CgYukvM2aOwTfAI2+uHS2rkIC4ffNNh5dmImpEyIVpw+626LfvkgPVeYjme
GUKOoBmWlYh8Rco3S0QFm6Q0IeYiUyBShH2zj7jvD3kqxgIHvDkhsMkwze4b2joc
gRrBf31SYaQ03dgws+uYq/njLcQz1iOfjpLD2hjcSryKkXOd/wIYyQz851Wv2qL7
iEaAmmBDrN2nQNkvyc9CabI2SrYB9wrl5Rz+C2MWUPectWMU9PJeIGTudqlJ1FSH
gpAiKCZoNCdW21Z5pwXNhY4t6TxOnnWhGQaIdVM3PU+9+K7K7/dh8dun4nU1wKJO
dyJLoEbTQXavSwvOHkBm3uRTEYZZ9TD+vCIeTHI6FuuhSq6+VRN0h5jmG+cVpXw+
NzVqTaL12srUKiEa/pqDM+YIM8FzgWvBJHMgNYT7SHvNKmoNEg6ILqGQhAJMtA5m
tQWa7NlTjQqRa+kkIL3XpMRWFr5eyK3fY58oAwd7ZbVsy6O/9HaUYSt1locZFcfW
dCjswyssh0eORqpSbQR4M09zv9PLpufclyRciJZU5E7IEid3YLpaNIvhmcvGOnvk
uau4izP8hI+/S4JIgse/Ga2cgAFeaejMm9+p19ttIsJoV6sJ9B+lBuXhMJTZPc5u
55/3SDMMzG7o6xEMKyGMqmxTsxOHw4tuJupaYJVfm12ym+96ehbPnHmXrUX6dLmC
oPwSCloJSetKZZgmkTxFfUr+ki/00GQ3QL5I6I1qVc3kwN+cslAiOzQkwPXv/+05
euFs4et4KNGVDV8tNPsSq67ugYit59M2BM8Cf872MMrDw7pBBMyC4UjkeBqH0RZ5
k1Z4IaJCBxljr7GKxd2NAUyI+1Tg3zgV+fpBOtm6YdRHxRgrN+4iyjBs2TngLLkg
U9kSCevcFTbZjOiRlM5Xo4D84S3JJv0XJjxZc5OAxoLLehVW87Tjcn+Bjj03PVW0
5vaQ/vH3s51e5emxpWeqkKfQabf0mS7SAvtUmTWDyvTQfQo0SmTR20gJGCErkeQR
zSiroUSgkgEsFrGvBVQTNge72DzSfKoHiwE77wHq25cjyhDVnigcIxK2qN4GlW/m
BW5GAvEUdkZ8JX2rstp6ShFGB5L+mxRoB5mrrHJN4/Vw8mF7Op/CGSlOrhaeyFsL
qQX2c0jDX8Dt0JPTzFi/ASmdn/c5sFYk/mvaEAHrwUJtTUS8rdvM9aWfK+ccs2qq
cui4TQDcLnxjss4DYGYgOfjATWwAZ5HcFEIRSYWOcTXZ0JfLTwUvOkb/QRw35eL3
h/IlG4KifQy8oNsaDbdRPmZB4al2MveSOoc12KA/W0NA6ioLQS83VuZkqjb9+9yA
z9VfapaJfzJgNW4QWA+HPzLATfzTWSN2QRmyHjF5bg8XZrYP5maAisYPLS4hIMVu
2VRoIDNgOjv0yWKpg/wslDXXq+lpUtU6GknaEbiK88lpk+KvRFJ40HI+I19NzdzA
dLlmzC6mrTMsxzIp6W7j74aubPiT570BKUUkt7akBEM0m6rzFXhVtjY2TrDv/emA
4EjLf3DFPRDknqLZKp8F7BgqkjcO0JhujtRMBRCi/Aktm1QUYeW4nk7wut4G/fAC
Q4EzTafMBWs+CuZ58zmLw7/LsyXjeYGct0yeU2lOs+Qz6H3o+U1u3iIJNk7GH0Jh
Fz5WgedxH1n5hJQ9fQYw4tZh+ijDhkmkRq+gAuqbBufvxAdpNVaam7ubUZkI3pqd
XI4NjnSnAmHatFflocGQRDziHhNZ4/XOYDX3td5murkhY7kiJ4+bmtAJir0Tj4gc
FblUXpjeYfvT4QwVyihefVd0qVFPmmj8tPJ+rPxd6dN3UjiAAr6k7d9QEdSCwv92
30xOq8Gy7wnSFeabQyRC7LwfZRu0S3t2vzZ4C/cst4t0nDEycFL1A+qbIuXLvQ2U
CzmqcZFk8dt8sjMlG9iAbFN2Tb44LhdiB08MQXKkYdGjj6F0f0rSjIR1yEfzDg6U
VwCM4m3b4XUSuxmFAhbud+1R0d77f4NHUpUuv0NU9sIpyfAnXA6LyWXih1JuQQal
vJIw0ASWTVApla+QdsR2d26remXagM7zTYLMYsRdF+R7A8IfSxtQHjGQSpYfMtfJ
AAowxJ6tY94r7IWWSHiUvUlGXUk71MQ1cpMGYwgaNI+JNIKbF1tnMQY1j+fQ8eoO
qLNk6sulhsB/xkjhpeaI2mWvS+f3IDxz9FQ4o6lAXw6TjzLojKrMaERRDlG52B4c
Lmwg4MvMEctBcCQWd7EThotkaLZTH9AH9FebB6U3CRzWRAJFoNaziPLh2ZpQGUX5
zzb+rLHsG5NybiIib9N9iup4ryBBwOm4k3y5xdjGOorwBFBVZNdnEXzq6rrJrD6m
4N11i4cGjPsiZtUbLoVF1EDWqEMbTpFYGxSd/C2vXDS1RhRnwfk9/inXlAyPe/PT
BpxhjF7AUDwjewOkCX48u4j/fUnX2Oe68fGzLNxMRgXScKBulKv3cqweQv3DWJu/
LcyQnQFq16Ye1Dnvva/q6YGDGCS4LLSBv2CsNzIogQn9m15tyZTX7md6nRqjNyjP
oyajPFFshbPvXxRw4L4UPR6EU3q6bL/mHyD0PSB26GF8USk/jbH9DAMrs8MITJIJ
pC7XxLdaBoMF9v0NkujPvc73pHx0obMYL66iZx+DcTZbimz/3efSsTPpc/i8O5IU
GVIDWjWsI0zmsD5oGpiFaAGbyX3oWXS/Grg4Wmg4+vIxCoOgnu/e13bnbuyuEd6H
witkOKnAvlZYmNG8My4RZpZ7XS/vpR3SwYd5wyJjct5wG5YXrOR2OU77Uor/5pxk
jOUPmG73gYXPevWKOtph/dbwYTAWaZt2x9kgqB441rWaLM/78vty7lNQrMMeJnJ2
T4dIXXAlt35VRIg4b4hEVSB+7lkI0ds63EadY4dD1XY/hi/0vfwp2Vb7dQjTmXDE
LUNqqmvP7wglXDRzHDqkbfAYch2QgJNlgzUakRm0Jh7uBPQj8DAdBouHT2OqFFGs
iRQYFNE3A4l/Rwr1LDPx2BUJr/OmiJIXBzzU82ZhCTQ+kGSd6NLAap8o2G/Mk4mF
tj15u67RpscSrZgSZhX/vjpo9tQwDgAXCPzbcOSwl2w4juKR6BBFKO3ghd/+dwsH
F3Yg8dAQesQIXKmg+XciqDNe9Wl3S1KevZcLi2M+9u3xTp6Ek1YTArdkjUPnWXXS
VOb53mqHn5aM1UZFtz9rFu+LHMNusaLHc4U6zxcTbaQETdUSvg54OaGEMXRXwTmd
X2M7pz9Pkjy8teOQ4/WngDct4NTnBQ3bCNWeZ9EHJB5DLSAarv+6iC4l8OK13j0Q
s9XraBb8Pgv7uu2F2P/BChkRCN0yQ4yiYgdAr9a68rBiE3wdxzp9Mg7tNnvQ9HIh
bdUS4X36MwvLTxKkmzRR9Hl0NTEPU0J4/nYhP0TMCEzJgKfC9qboFwBIyOGSljiS
soXbkXGRqAjfG+ssV7TpxknwEs89XRpbYDBCNXvKWu19N1tcKNTjDjyi+R+pReVx
UvxM4dad8ewEPWUu1q0b98SVFVlTcsdJ1e6/kvy3wJWJwghnsA8POzZcUZKdqW0E
Cj9PVQ8r3VrY8MX1BwjzrEL4LbaVgsKGc2e/QhweF57jH+rkd8xB4wrQZZbf14Xs
PWX42aI5c1MVYLDM3tY3EMmnp4In09vQm8DcvOQi3Ts3ibdVg81pbkyeL21bFKWF
U1jducopSmYhZXy4YJ+5TrPaFGq9MyqKalMoo41OygFKGMfMx11FTlcl/F0XbP/P
QgNd8TBOd4t9uEP7iFzUKAIbrFigCNyooDsMOBRofkuwunxWtxH8JMX0+aJQ3Wc1
OkgmSujRLi3tJgTI5AhrK2ZV48kv4P1F3BUXlu3r4YLmOwpC9UyyJs1qyMZ4KiII
2n0L34+EnY8W9elQkgQgL1k84+eZEi1JVRlAaJNnUHlRH3V00VlMSEPddjCiRBKB
tJA4pBMtGLX4mcJ2puXMwieBzoEC8q3H2gkGnqKyXRqG+WUYlxybXp/fhO4iEeas
7RgwG6z0BhDx+37xLze4XBUK3bDcXPmIm+IUjthv6QIYz/PwBoKFdqxc59VrvpKJ
KzzeaFJMRvfS3YBqUS7T6hNT8x5nTRKp0rxDC1JIID0EhNpqVwXOUBXnC29TLiMn
gWqBQty3cbefssb0Smih7otSNWvyEVuyeUiPgAABdi6yRFG2S89AkWCP81nhH4q1
3STNEw3eD6nM1IwKL9aSAaey01X2G0Yo6DjQHF2Q3L0WBfc+/UTUWjgNPRO95kGN
k0/cbJ3UzXXp02MTuAzfKQXr2yRXZy7pwz/1X/SPGR00kp8iBFGKEUAi+q6EmMwY
oiWYgpf4z7MrrsDjfqMsceq9K2tZKs9CNMNPBj0qAix4+leXxnyvrok6+DJST4ov
9n1n8tasKyDqPGAeuBjAhdApYuxXtDKkzt8lcdGRHP4+gieORw4/2rpa2EMcJyjW
sxtA4gULg/BxsmWaoAdEi3NtKmpDxQrh8LR5bmEqvqNbK/h3TAqbMWpjxmi4XXoW
e1qSxZre2Wxr5XUmoM75GpG2TeHifTyplPXFWnNX/jBuv1hBDeP3GYOpxQx7H8ZE
8GU+oEn4QEXD0RI8ETo+QSdZMM7verlYVjw5hQfGfyQcoBw1bAzn/g7mcBdHroVi
SfPDcO0NiYJv1vjE2ukgLk6TjqbnGUQlnRtIxnmnMbgm6Y7LV6SWQSyR42395peZ
o0E8TZRMU9Ab8ijj1KC2HpPuROnGhW95rlk8PUmUubeTkNvgO6W75nYHmfY8Bm0+
mh9QJnSpU/xk2ylcIY3JdAZB4AU38stIufA26+eWbKx2+4ICtQ4i6uVAOO2+9sJZ
D2fQoSZx5uprQ3ZUVNrV7vmIhEO2B9tshlqNXmf3iI/o962DL8dD/9ivHUWf14px
eXCmz8aJK4B6lyXo0TatasCjzBGb8F/eVHpX4Pgd7uPKUnm2exLZYamqdgZ0DNZ0
NmaFX+Lggik/TuGBmcHIbOieS7QjQnCS6PnA7Yqg+wXBl36op4mlRB2J1BREriu5
HLL6vSUf9MFeQPyYSZdTU2UpXaqqAjy0Ti8XeubcOCNeiMX4sJFparKBaw28IM+2
MoqLaa7heYsyY4x8G0xGs30EEB1pSB6C/q4+pyptjwjknHc03u8BD8ejkjqddbnX
oKgvf1j5b2+mQGfxj1OKJbHBE0gzOq2AR/qZc+FS78jW1V7rGZzkVmBbHjLnpRt5
yqf+lozSyiZyd0Bhz9B1xyxtKKdO8zDpPSltU1Z3sTTC4+6xrX4C1VKB2aPH1TLH
Zym+tB4Xmbq+Rx0ij8tV9SmnTwwNHxInF2YeheLRbZOKZz/rLBNu1o2u1aNWtS15
xP1Wvs+d7GPmVEvmsbJx0WNO/bcK8UgrXCbkZYUkvpUpVQztXUj8CifaeYuXT1Ap
IiyuGAvh8cBChrcWTQjS2IhgmDQZhnbQpuX2Z7KJqQ1eeslAM/1tG/6ghaermTHe
AX06NKoswguBtS8idZcnZ2OANOhlcp6nZk9GIs5201RwCiLzTHC2gIIKrkPzKrCD
3Licgpcsu+tUqFQoskzS2p10kD2o0M36DPcn1gzdNABUMhRWpGUBwm9jRaHCUah2
Nm2HfTBvguBL9NTMrg41aM50qsThtWVU2lXvpNncyqqZJWUDky5/+1PgVVszCWge
8ImVKA2l1wUeXX962uA0RrWf5E8wtcRxcgrOxNWKEUNnrAwzERto4ZetNS+dI+mg
u22PoJRjbpqxsyPOX5gIiBWAEzKIsOiGLBvLAD+bRsyTT2LQJ6wBltEjKiJPXoE4
MN0YsFxyJkXPC/CBRGvOBRJVFxnOC3gYT8P7nsLwTSFBHidWs2OFh4TdUeepvx1/
1dZO9HEoiCbHSCmdUOfPf6QaTmsaBhaNpKwUn9Zbyt2X+2Rfzp3pAyVBtNgUsTNA
JsQVbPuAEtu7BjDek14ZQbqzDqYlKu0P60X978aKGCBYLn8DA3xzNtPnfyoSSXUR
QKAdmYOgs0meUp63Eh0Qek64eFY9Ucrr1ovkB6qJDUXHC+TpnXxip3ZEw62OMaKv
N4JaQ9B+/Zx71x0YP4mWKOPagkMYeqzULqiLCBadYeEOY3vQ5ObR2KA5SBxBL/5H
IQFKQzugbXS0PZs6pr/VPJ3eOICwTJPWD5fV0H6ORfZWeYNbIrOJnEScdPv5PKnu
TZh7FOLcTlZonUqd65P0QZROvEa9NKZgCl3bnWODTjA1Px6D/gDadkE8hDFP6SNr
jW6rx0VSlXB1qT0v/Clp0ixtWaJc5SbVcdekcZ9LkdyntjU0VTgniVq2N1fv5S3A
9Av2N7Yb6+jsFKHSEItTZux+INWA1VThVsFHgHkCEuLACWpqQF+VdyXZgY1J/Yz6
WYPGP8vsClErLOfgNKoZm9ZPYcnUSKIswS48cT+GTQMxNbTOENK5k55V/8wyzD4Y
IzgZ9A8/ylS9awMUl8rtSfO0+a6TezKxku1caFEASQHY3rrT058Z4mJY3tAXDJay
MMOsBqY0d+v62fUXE0DEaaMYsApDMrgcw7zGdwbIe61ZLiUTypN7K4QX8zQwXigx
PwsyJuq2cnaN7YcbBHHHoyNtuLPXL6py3M7ulSWClblR+VhVGois/co34M3OLsiQ
higPHENPRyZHwUGfX2Y0YXInZmCqnE4v1pK2IeaTc7rDSa5Nya1XLxRH47Fh/912
cGnuHWUVAkL41eu7F605ykZRKUJy6l5A/weP+2Mw3REISrXqXsQEej69t917Xwu1
K1FvghKRMwlIn6BFQUmi1Nl9NcH+4aT1DIMsO05aTpYtCr+WU7XWcaOF2l6/g/Jb
Uze6O9h+5UGDb75E4HZjmhb1W+0HbNjmhSMfztdQhHI877LzWezSDE96rMgLGdEY
OWbLbsSX9qrul2N/a6SczfRnO7HOuIBXraHGcS7y1jmUPAj0kb4up+jpznsAM2yE
HplV/TPzJcIfeNKx+Se4Norr5o7GLieIIEI+WAr96WF1KZPlgBwA/4hY1wMbnjz9
iqJTcqkunSaVXXUn2CWVytgE7MzRhGcBDENAlTwsi0ExsEF0nJX42RWUDfW3ASJ8
xcWqXExxNRd3Kg0QokhTifPIko3ps8nprhu5hxBMK53zE5pa4NSpAQRxxRyjeipz
nyedUv4P/dTL1PEx7oDyrLj51lcYD3av02CDzR+ezJhtEXpXKJnjvNbBqqBAOS5w
+DpEysCKk0Ultb43TbamXVrZUpd4+bCKnd9TuO0925ohElUCj4IIkmfmcUkJDM2S
KFNgUaFwxibj+Cz4YOlBSIY7DWBZuix/nsIdW8Do4tIomDXZIf4tyg8ez2/hMH7l
TEplokxGuZQ5EPQ2aKmhh2TH0JVpnLNcY30lQHtKcx4gyxqRqJxvjdyqLBpEuWrA
XRIAVCyrFdZ2zWu52zoh5ke/8sHs+lTXFCOITzsIqTBw+RGsAN87CiTmCdCxtcQ4
k6L75DsieEQSTCKriT+Ag8JDQYPinZ2pPdAEHf3Qv39IZ+wX1M5W5y3W/5ooH4op
o/FzOit6SIJGY4dyicrhUwU5eVMmmLnUAfjrjnTG6OUuzTIDgBKnI14ogLoKF2tt
Zq8UVDMlhTw0jPfQ2xV7WZDk5S2vwA4gTJtrEBDP91b1kQWf4B+AfA/MdWCMavDH
81+k/iz/46Hu2UkqxYqkkHcdf3q7sWOxnFmhUc2nZthT8NhcGA2M70WiG/fEXqU+
sZ1kQNqEq8WxdGL4x9MG+mhsBW4/5jwtS6XMTGkROmeIPHmTmSRsRPSlEbQyz9Pn
t/qY9XhBWkqZxsIcfS6pOVpLwkZzzbt5+/78vGJ+fggLicPZ90Z0t4ebDrUSuV6i
cVo4uG7M2O4LfGvYYGEzEcodBAmUjyUunwa2Mv7oGynl98KDZmXnPVNN+J0z5DWj
yRvAdMyZ6/FGFHllVoh7GlkwUeWm5AcFJkHLxdAfS+LSAX+tcMhcWPJRncwsqhH7
631suRU5NheLkTM/gE93DCIsXCdDlxpqYFavyMD8oBEwegP7azFK0zt0QJENJPuK
q8mCtJe9cpJoL9BESH7uhRN1adPBLG87KId9wHrkyZd5/vJuqRHiLvH3M9CZbidk
Uevzxgd+E9A6oD71vzkFYUWE72XIX3wJSjlTeKhb3BCnN0/TDHhjySkwfKM3E7fI
5t6wGzsfoLnjQt09w/pOKYhGo2gd59ViOwZM3q0xQI8DI7EpBidbx0CJKjuHm+es
p/qPcn6pL/uUrAan8/nOA6Rox9H0Rbw8+x3TdrXltVcMQ5Ub7vWyg51PKpL0hOfN
mVrteV9KFsm3fdUn6Qb6kTY0rdAJvHEX35j5cCmKWNmTHIee/4RaCQOoEPKR7New
hkqbxidCxvvbTi4XvvvJ+zBKAKCCjW8E0N7A5eLzo65OW5yi86/GKmjFZBEnuB8e
yPubnP21PmRpYm6hun8l/WaDAw15lY+Qfi37lTZ9h4VD4ULW8FZSRd9IJv3h7Jha
ZNxU8zjg2gPgwQNcrBAfnMWwhU/5l6tQ1J7CZ0wDb4PbEb8oSf6CJPMGv6YfnnI+
RvTFS9lHfefsRXszH4A+PXXHTuH4/OPT1ZuKUl6yagYLT0dIwUHOL+rhpMZKjugN
vLF8QYaCe2DoOwdl6A9MWa2JVXED0UkG502uv7MBeJQg5Is/Z5H9WHSHcCSmOtSc
u7YlIFsXZGkdlCHvmdRhQYgfZhXqJk6YMcPtMeDqkyX7T+NPKZ6zuhs3yiZHEDb8
40Dtt90ZAbdgpHcKyvVLmEComMPNG28iwzWZtESrIbCw9uxsLLHqkIuM//eejz6z
cuNHZCSJaMBCT+BsNzjEhwXiex0CEpPRvbrFxq7S6fHA62esLofswxgdWWoFXYMT
88kHnUuMyef68/bzk1B2+N7fImtzuczY1DyN71VlMKfJ2fqWnthxoM9wZSBry+6K
3EeXHnI6J9UM1bCHrheKcHts/G9RPsedNldtmP0/op7bqd7Zr1G+dC0bPzfpQK+d
hUVxNLZW7L7UUPGcl0g/E2cO/so2KxEUCKTVhx3WhO3I3r1HTK7oEP4x/fMEGCv/
wXeFPDJwokvne8nyQFm3XUBClOygkEtNACqD6QEC0mKis3pDsFO5UYcI2OCC8rnD
gMwVejcVQVVLzMzcpaDeb7jbzdFiyekc7sHHZdcPfnjvclhllHvmjrf2B9VFJ+3W
EJAdoYVC+u28qm2H8zLS+ECE/VOSD8wZ1WAMo7/gdXc0ZFaue57QZQLPHXMSnrsR
plI9t2l4HA1nvch4UDL79LcukmBrH9UwR6NhMe8Hu06u5T5sxS+HesUD1F3AUwqw
JEzB+voGzz+oP89ZfDF710zvAaJTElpYuYBjnTR0Z1s+SUKzWAqJwWUE0Q/81Yss
jg5RiE98MRVv9L1njAPHl3scHoE2dPFHFNzz11Di99sFYN3eAVashZEjHxMA1VSN
PE8JNnkp2eD6D2IGgbiu+lRaqcj0Xr1LJpZW7Pk8SvoThq359x1eLA9N6frUyFDE
Vq/svAeXykX8WPJMm6ZaQXObd/2XPdZBoWWjiXeZH7TVET/Y2fjR8JVnHu/+QH26
RXVzATv/lCl8pSH+oaeTVso3lpZHfWoDXQ+3i2ZDGi6Wk2RsUwg48AJ4ULs25YmZ
KUDrtMUenbaIsQ97bnoP2YJSNMlwc5ib2R9iCxRaoWldGklr+2uEpo/kmtYJU+EY
5DoRC4iZ4+dol0H3eDtVK9an/S+mPkBvkfwJyHR0kccso+a6rVc3e1ScpwdseUqZ
hhFoKj16q6EN6wG71wXzV7VWNEiY3FarOn7jqMi1NtR6DhmOSBCMeK+5oFhIuwvU
jJukQhTk/sdKyQ6ufhfrtzg99/Zon5Rn0l5YFdJJtfsFCFrGn4FsNlY669AiOshX
OGE4/9emwKvoI7mlj12PuxkHub7e1tivw/BSsBEZID3+Z4fDRqvKCQqJlXHDGp1P
kUVDLxyNDN4g+GsumqBUK+o9yai9gDUaenEbHTl9d88R6Pn/l08pBRS1H0af5RYL
emFsNjD29DJeAb0qh7Tj2pg0FIKFLlSqD9uzOp3S4MJctTXZfLrps9e2bK0PqMTJ
NyFacxiQsRWWcnJwZ2gbHzQBD2BSUSjxLhQgaRH+wEFM1VPWCwyluB7k/RMVCalb
PyDeQylep8yEPRmcSP9rghVH484KppkGqaPjyBl+CSZ/D9rFPY1nuM4YCrC8AWXR
FIj5yQwLCW83BR76iou28H8XJbRSoeS6YHHDtQfCqUpxGse2cHJ53jlK4PxRO+rl
lBzyVjcFcqWzDKYf3CiIJotjVs7ooN1l5/EjahuRkDsO9Uyc9OUcNFwgZgue/ou5
kBmNWLb8L8SnD/5/OFT9Aay0uGr59OBllW1NjuxDWwg4MknfZKI9WdU6IBK0Qm/7
/5Zv4Oc+wd7vhVmfRRWnHK4l61/OamfjYmnPtoPKNi42VQ4n4xDXL9zpFWNuXHgx
6/MlyDIKqKZqYAqKhVgwqnAFpJOlc8Fb3rZWLBownVXqokx4YwOA9V9nsCeRmz20
2MtEx3xUaqmv6VCsNrXwBt/R3ifExy0qz//ogaQmT3BOQwgcmklmXEt7+BP1XKjd
RPoVrvQOqeLyswcDiTK+sjaFHGr61BkSRpUFHBUQaV8nPHFcZvvysbZvex+08kbZ
lOoKsDbZJgLYmqPVWAPq1TVUG1rFls1EGUw7Y93r18xXjWOVSrY1sPVaQZddDPhI
prAWxa0z8JRBqDnHWfb/iEp1ZdmZ2742LHFEgIiHYI29jq06KOHo4H9QtMmzK7VA
selQSV8f1HqlhSOL+dY9wZVhHJhPq4+J5pi4IOAFIfL8smEUyaIV9oHscbVdW6FQ
Pe7YimLKrHKyxk69BDLypqSHuEQQojnf0ZqYqw73YLdqRCwqF1ysKIcM4e4G1s8b
y0v3lH5OSajl9QBNn8wH2wPGCwZxmRzcai0c2RVSQ6XnMI9ibU/X3HOlpsAtdoJF
IHi0AohybF/aPNuYezAm8l3HDPOJZ9dw7hbiRGshRH6l2f26An94h8bW0gF5dNRu
NmzJlSX5xga0Aver+UQ+moiX75EulKaZqhmPhMiNimZ1JQGJeC6hEY0zqiXzJbtf
8nS5nCzJHDulsBAiugAigz9gfpvAIn8cuB9NE/JbKEBLQkx64rvch/1U0q6STx3U
nEMWlgCJaJPREYdbhotrQFDYLwtNIbk9jUJsC+WMfHA964ygZPRJaKBazELJ2TUQ
JRUss69tDX2L6NddJMZz+iA2vgaOX3iqACkjS99VSRmWgIrhs/r+yGf8palZiFkg
/ZQZUtCc5kF2w5bSasGcRXdTa7RHy+ZfiaKwXzIawt579kAzSM8SHvL5PmhvqCCD
SlIvYM9QV4IF3Z8SLAhbQo6Me4XqHwO5oZ+lmR6bNA05c514Jib8Ck6ok5o8NTJz
eYu8bxKmRwyA1nhAzhF1r+3J6nJeV812/FVj8TsKjl3ZQzrVBnqgaCd8ZYie1vnJ
4mfPCKBo9OfQJwGyNdHzJi+njqZ59IPvxWM/SL77I4pDvADvuYjtpW6MAEoVq8Hi
G9GLnYY5gk9qL3JzCEEq8wsuGap1Ch6OG8CHSr3QKFTtzH2XDxpxKdwqXjmswSb/
Xy1QPCR3CCvsarItr1ONBjJloAmwJe/eCJeXGAOJDd4mVVHdVSjIy/rDYqoQsGZJ
HsfIRszL23KKEISVJHdOS33Cc27DNBZr8HLIn98AL2ZA/oMtUF1Bx9B6ELPo5RBR
Net0WDx+kJbQly91Jsq4ZW2Ixg7BRJz04gDc/BG3gnZY0tVJ5gQ7sdvkd+Wt9B/j
M6KM431OkGW2CYurpshD4yPAzJscuU2fX3Zmw8hnFTO48iLQH1eGb+mh3p6d7zmI
eRyqMnCcl1JfMyB52LqCSjvJjrnO0b1L9ukS62n0qpxeC3skk4Dh7vQQp0mSwOJ4
WQ7WLpK56X9V8o8d/dzO9nDImMCFZwwwxEwXZ2mJD6fmj3O8UyCwkt4EKF7ZyZho
tL8GCZ8jIh5kaWkjJ4myWUk+LptHveOSsXKZvzFn+Rj5OJsbYAAPyUqHq+wSviNj
jZu9DQRsvmJBej0Kp7jZNhlbMemV+ntjprlR0p3SsbQnjwyYl/mQPnnzMqgLqn/h
RF2+x6uJjC1QcOCQOiQMCj1QfUxo4NHn0gbQES3jjOs07ZCl8f8lcUQ6N2Ls9HI9
3nmERbeiJ3Y8LlnEEiXayI84xyxm3x3q+ZTkZQH/CtCMHwOXv41F3INScae4qjK/
CjDuyLvj5JUwA+LSmIV///ldxIhpWBhDRQOSJu0K+0HQAaUrJzxulvDA0MHUPbn1
2naczk7yj37UrmhigfQBbG5IcYBDCi1L5fFIAi/AY/OP2F1a/EGrtVs7roMUg/wY
2a5JBH798zfnD8QbWCk+ZXATTf+ccmf3GlJKoPTh77BrGg6Im5Mn26QurBRheGVd
Ww/ZtgqgjSVgZuo2mN1hsUrUvWziD8au3/IzqB3dl5RpZGNfmyWXMtnaKWj8pLat
6/Wzz/VvZOD5TUbPFpW4FmWaJ5CyqmBtJLYkhHrlF7FJy+HjboOeEmb3gGf4Rg3x
3JYBLFCdy8xjKCtHK018vAcW8PslGl8B2HooflMef7HpjRqGSn8r7DYuW1xL1EgS
ODEYudovIqxFtSuAKesO1WJx3Yq/Fath1DDs554hKmjE/Z9H7FO9dTkolBT44pkV
rtY2FO1kFcYnA57Nf3EDC1HGfv8IC9IPoc9PohaR1YEFvRRGAu7cEF9lNOqT+zny
UwYVaFIj34xDkVjsuOil2eJ9ORQnl8mMbfhRXjkL1NJoHJM6h1hRBoJDwbZEiHaz
01zsPP7PaA0fCHNlZBtumHe4AISE/v2+b9jA9hYWTzt3gUvNAiCtri+q/A/XdIjZ
eh6JTXWDaqX+47ftWyYQRb6b8qoONK+APx6+GHCp0JhqIHuFaR3bV163rh6kryE0
9XIxi8ZAHARBq8HVJvDuu7UFABwI+gB/TZuQDC3j5N8FB65zwDMqXErNDeSbnSX0
x2JIz1Dt8yKSvfIaljrlkuot7mfbCvSSEL3EscUQXJ7K+cetYWB9v5rUra78nzzL
mXMW8qaus60GUAGzxNxTUM+PwjwY3+uN76pdGyAgQxOyTx3jUws44HnWMqIK27cT
fVg3zbOW5UmrCwl0pmoTgJwBuB4JYv2NBMA74GPGmuATGnEzsDRvzghjGECKD4sc
zdGt6EBwShyBTDe2DJYTwvW+3BQzvEB3peBA5XZ4unYis8IZYZbLV9cewEVCI9cY
QZ522yZGHwxFlgCTK8+ts54He5X+YmQqkUiUf8sPrEjedTewwPplmvFADqMqYoOn
qhYgfAFV5BJBU5R7y6CxrmZ1kEU7mqsIYax0ayw+Qye2Z8auZblM0uhLv9DRwWD/
+f16FsuqgtyIHM3Qlq1bYJybLzjxmJgdQSrJFd1kXu8zyIfzbdRgKZyUhIo7OHnZ
wHjhQEnIhmLCk8jIme29HKSkLRF25EKo2wwBQ7K43m6Dp3RxTvnwOfA53ji1oIrA
vLIv69mSdEXS1VYI/ERX0KuKoyMZuzhOwV1LS79TulYhtURWvm5lNKVcwA2N0gfs
LAd0GqPzQzm8a6sU8jPdPchuvqoGd4MOibzNy4GvjQ+olpACa48JoBD0YjX2C9GR
DEzGipAXgkKupq5lOOQhpkfq95+8vDNC/Ddx/Xfr8QN0y+cHwVijiUYHpaKSJSln
8QukoGpBD2ZwROf2pKnP9EmT0F77U0exlWaalW4ge6taoxkRoMe90ZTpx/+luKbt
dA3mFvav3/Kv6j6oHiqC7W2W/C9JD8UcLSgoxQJukuz2+r5lyURCtBInbb3M1Ggv
ybZeTsG+ma3uE2t2ElCOAx8S3ivQN3WsPu2PbWDjfA1tc7pEBnLVR/OL1W8rVziB
iqrEFdCg75D24yqmVhCda/K7wFw+YKjiZAuo3GPSc1YC0JNNVXawABCLSSliZkR/
JSb2PC7Fuzp/QI0Xd2avTDkAPDl//7LvpY6LaYShKNgQY84y9gkvCpVV4x3Mk/OF
GKU1oL2g7NR7xWqVi2pSXfI8RDxPCczL+yaE36lgvTtuIqnlor/ozpKU3/pQzeai
xMrq+xaoG8zUVRtYAuujmlhJlm5FUlNn1yZZ5O/3EC+4CHFcLRPjBu4kxKptPsYS
4dRe59BsThogsmW5WM8mxuAHyBFPZqld9QlcJiwVKpcPccXqqV571fCRejES8vCf
TXgnfCVKeyccERld63GILABV6RDGDdpsFh47V964fkbpjKfGfyd1Gf/Sud7+a+m7
lmUrJxNxyzMOjc1h2ly0txa5HBkAp4lFSR5FKQ5m+tg/3OAG6ly+WY00sgVe8Ied
a0TvvlKOIxs46SIdp2vldDlDGb+uj49EsP7OU4PWkesT3XRg1lM5rQmz5fPvG+FQ
uusY+DGEvUTModcRFvUIcM2GF2SM3SQVfir70AR1j0T59V0Z4zpRJn4xBKD8zs+J
KvEJuVRBfmEYl2wWEC8dtELCJbdiGD+dBaqn6mLU5ogTYmy1Y9Jmy1mIgxReURuz
y0fElIuNg8fiKf0GNqVMxA6pn/tHBalQYFK0M4QA8gDf3D73r6+5g57kR+u9H3XG
bWzKddQp0PmgyqAgWqvWzY409kzVkoN54b6Moha/G9NN0M+I8ugKXURqdUsKz+hB
PeAd3vM5ZMBFT0Ft4BQcSNjpQkhwlzCJpE2I0zCv0kZ5ynez786MzhhK/fusC3Qk
sTCASugq8hvXD6IANcFSwGNNtfcv1zPrYPEshkCID1j/RdXP1DN16ookp9IcvbXA
/RZPoVKcOrJwdlkkY21xCxE90xYjF6hwaPup9KuHonTUsMexgV3mA27DXs1ehYHU
+XskEj2sZU+8Jkdw+f6OWOfTGFVEyrYsc03iuEj2OrqlaGb4RKwFISqmBx36662a
BBxpF+3TfYUfWQlxyFr71/yEsASquqOsuMWLsAV+LS/X5W53yxbGwZp1zARUKrUW
7QjBCkG3Mdw0Xt02xtcbgAxsVtOtxaCBaQGJij6PGMQhVjRCdH4Xiv5J2pCchQRV
yGjoYnYr0lUzhwCTrJiMzwUM/w9T45VdFGqULl3emqVqKfPOceQlqSN7oZ8wexQD
4dQaIrFelimS/f4GsioDJT+VkM7PyX59tGb1q96MzIn2pfBDoW6e6cRMqs3Xj9K9
+J4KfN/Zq61NMYySIU0XbEJO2hRLvcOE2mt/KyJG2W49N++/RR2w6C55bfDpR4lR
KR8phtUe4BZvGNrBKJ90CSU0WzZ3IUKyhmTbRKVj65fAExVZvCDb2eEJs8VgFWMl
q/Q4xwgLNgo4mDfLcQ113XWYgDXaVrJLqawkqMX7UTx2yKBblF1MI5ko7HrzWKa0
9FXUZ3hZd15nSaLM0pLaRbl5mokNkNPmr7ZGBP0wInZj8+ca26mYGWTCCAWeKStr
HG7vwqMu3iRoVlfk1q5TZYDCaRMTQ6t2fHSpVUgU8Qj1NQaEk+uqThhQzFXmXP7J
xx37mZMO9CiVtnHZslAsVpUnOnk3iCwRDRaVi90sTB5QN7CPKkvmvOFlyPS6pRc5
2ynBDt95L7nZ0WTCIuyJFmY2kFqwgeESzMqkSWY5Ww24G0xBlflCUcrA3onzxz6Y
DcrXPyE90O8k/v8M/s+KR3eYTx/eCBt2N1Sz+WJ3XPPeaWyCG+X2dBmJH6aRfxw/
XvNtA9C22FFMoFO9WgtdYHO/9V1p2eM9r0fEdFNw9yP6+uo/+mfPQMp82OIb/VkW
lvff5iM1oc/QEyhyIe5dFhEDD/4aq2FdeP7WjMtcdjjBqUtPEDuIRkvQDB6huspz
mVQGIRIOBiWQi6rMZOTfdRbIXll+vID4VRiPgutNJyKcHj5A1EbLV3sgYm424n6S
QLkLc0WxzC/tyfwftGvHXmmaqE7KBbqZPy9z5HgrODRHc6VxkHA5CVtndB/mC32W
ETemmXacjll60FGb5svM3ei1mbyLjhZE5sj/teUiNyyx5gNPaUGG38upNMrvokLI
ZdS4HHqwwfMB/4NhhGwmaiFiw3fn51BoIZtV81ICuM0NQ6aYfxDB3ZhNFy8sdJyf
YeahvKEW5sAULnoYYOHveDJnff6jonWgxcaZcsIKPQHkHqm4x2o7dVbhI0VWtOaQ
P09VnEMcPi2q/ydcuSoD8/mL7SdQbyDtord0Odt5T0HXt7rVoywAvKDHtsba3qoM
Bch7gtMQqK3csPTEXoS1W9FvS0+cpQa084k8Ri8nhRGWmVR69CYgq2GS0m9O1EF4
BEBOQSGgmthvG48XSfrol6tnQxKYNEER0NvPSYN/CZIIzju7lj+YlDSRusnb4Ei1
PxUl/aRbrfTax/Szvsci/cGvD+znuIBRnWIVZNKSQ52mp8P8N5ZyMmlFZVmhAElM
v2GyVWIcmWNnqlaReCxoWtQs6J/7RGX1rq+CNB8tKVTKRWhHR0x8XiMGEWwurcy/
CfNQ8AVMWETL6iN/eeCE6aWfBVCfFAbF+E5rwA2/HJyaikR7Yjk2yKcgYl09ECKA
V4/GQt4XdDlfQdq3pDOkXcqX7plmaOhOj+RatQ3Y9WRXKsaxEuDIRSF0rCe4YQ4c
6xYL5RNhGrp+eakGvBqfv/3XyKmJCWjhC+acaPwWQM+GBjCc/fJpPL/HxO0esUoa
qICrDvXVnH00UQ+7L3qnvtW6vx1nIqN/0+7tmZlPrCN/o+S1kZZNwbhNoc/fGy2U
UhI8WTV7Gqkpi2FBHRruqn2fxJGkLhXgd1bZLB7jGkX/Cj+8Dy/1mcbutTengMN8
cCZjcWHYCGwega3VjwoYGDRKewYLxg8l8YI88YNmmgjfn764CIU/w63s8RjskupG
5fqtXy13lf5IKX7MMbRoLkkFdck+z7mwzYTpTZ9v59ak5jNxPKvpE39VTxVi1fEg
7k0OKv8fJ55pXpuW4MoCrdCPmxZw0EO4bvgLGo7NKWf0Woyah7ma5P7H11hwOxt1
0xaR/eabGx66Jc0a3CcJMaFJ39kKUKKYY3Fwm2xnWG2jyNAZCE4WWVSofvUrJsQR
Qcp1zz2sMvO4cC1mAhWZgJE53pvpcktrFDzUzulTtBooXGzX/H31du3wK7Xh3MTn
92Bs7B4wriU0yt9Z2B0u4GphWaqgEtI/pKCKFRRBZ/DSHTrNRcD8bZuIqK7VUYEi
pjEPILUxv4DP5LbXfB5k+T2L0tCzZLKASpeL8gC8QeLJMinCoyzMsw1llFKC2hlS
AdcqpKvUnJe6nNdRJxvD1ZxU66iepSMlMLQ9hv/k46kAPNLnNLuARj40hAc9B9/0
g+EcaQ/5D9s4ooYC1v1D43ZbTPRzUADPBtHf4mxhMm7f1ljI37OfI/eObThOMI28
Z8CLgsI8zypsKBpPJbS5cqd5Ox0XLY+uo+e9KZULt0ica0BlbJqAEqtH8VRY9eni
5KNvrxz25kW1MV/Z9c9tmzcSeWN3cOjNKuT0csoGZKy/7wrZx2dDdgdgBIGsWADV
EPG7HYHie9WIOoPEhXy6TNPQVQZx+Er1Ef7owkmSzW9XApbdN6mti3Rli00tJryQ
JmVEGoeOgFeyKFZn5PPPOb4Ey88VqthuhXS4T0q+TMCwQ67ClWocWvk2/a+dpRLf
DVb7N9Wq8n/z8UkO4M5kjup1alregFt0R8b5+XS9PosyfaZcaQvelkwsO7ePeKeO
OWl+5lFDcFjbcg9AZCsqq3wv67+DsVuB5sGfdNxlnj9wwPCWninBA8F1nQnBYVu4
m/4WFo8AqoM1HcRPCjP+KHZQOAF8lHa5SAo0vI82oKWLvjbkJXjIhQHGY4Gm3dzG
0UjgXPJCPAtOasSWeBTjddjst2Wc9fzinoVxkvfI/VMkeUW72j1lrTEOlk6TMuXb
G742WsbkRqkCU/kXaoLHyHziOTDjCxVeoCGwyetSuou/5eXKeC6+KlXtjYzAWMUB
yMp/Izo+5OBkziCW5T7dcKq6Yp5aNMai66mD8eJGC2YuFHMNPquTiGmH1FXhqTVR
/qJLqMY6b0FRxZ8ALPnGGrsIzyqXAsnExwXNu1eu0z61rLnHYupN7OS42DuL/n52
9iMWKr+qhYu/DCIiYXo5KJP5UdbExlfKiPEVS1YNBfYOdiZ70JBKQ/quy0QSiDj+
7N0GrqiYMj6T2prdaFtHVcQdrGDHQ0MWnfzGRJyg9RhxNvIhGhIpfSj1/Lz44g/b
eEuC6oVDRtLcSulDhffJAuga5oVpnDfiibGlhOZAmpbaQ+3WOOHBrDD0IuTvydXL
LS9ZN/ikeAJHIRV6HUfx4EEMZFNNwnEskAeYZ/pPMlICKc8OFNOJPLaWg/U26Mhe
5+l+bGvi8OXxhTnD22+e/RFVUYMnVuUvQYDbar907vOyn7LUC5coDQ4x99I4dySQ
6wAPyWk2xbFqnKytWy+1pvkZb6/iq2c+T6nnMxaMVzm4OTu80hF8kBg26XS7JtCY
YDSbpifdhFRAnY2TY2jVXQrRxqBLMJR/abUY5vyC67usavlIc+CNp2l/fmkjXw4N
1Y68SE3/w398iVCvi8Via/d67/LAfZ3BDd8MQ0o65/I0bBNdfT6shINBaRUbk8Cy
c5+j/Tw20EhMpAL8f7mVoBF+Lb45y6udPEeJwHvjjZ7+KYfbBZQJ+ZWTVt2KJQml
F5lnSjp6U/+EwoWRrhlZXgLBQT0GwI68UHgGKafs4ORSL8tguLV48OMGi62SspkR
kixtRJzXaPOzyDj7LOaE5JOxNmzgHXZLhXa/uQoc9Hu8SzR7nR4+5WoRax94pE+E
wyPmxCQnNyns52cHPAjMECW03titVsRPO7G7uExcpt6uIyCg1MI9YGqk2Gw0Qkdp
AMg23fnOQS0LZRCuTPcfZxeRVoGd9o+CbUEgPmMoe7uoyNe9f+4YnStuzq1/2GD7
FBOGFSfvLr8GdrIaiYUbV3K8AYWWElOOFFOjjXeEIAdTmsC3mLu8eOQ7i5XtZ+5u
glfJGyNt9w46g88Tywz6hGRJoNVSjtExYbBD5L7HbW9XvZ7kHFJoao6D6vzNOm2/
TXN6LjdUFT6ggvvZ6PMIWuvfTtl78hDZhLJV8dPngeWdt66txQwG4R22fAfKzxof
zVojepHhA3LILVFoubt3KQSr8WeZaslYr4hyulIH7GBeV0TYXt6vwkidxKkVMsyk
mcPg/K9flmajXbQYDdC55EYvWIl+E4v9JZQltOZ6tV0bax2igAmTrDESQUAFnXLr
UDGxR3NkxitYQkv+StSQmiH2QA7hGnmNXUffXjIAkvEa468KB9IEJg1bJvY/LHrZ
Ai3tNlxstr+RudKub5d+i4/vYLBNDVwBSpf4vmrhEIiCzp4QG9fD41DpCFiyvTmv
htuHnVZdgv9QpI64YfZKee6QeI9unY0Kf/FQUf8ZGo9GPsYrq6Za2l3I/KH6F0m/
zU3MgLzv/Ug1A/WV3DlVgJXNYuk/ljKlFq28sy1eQm+1lAu8RyAc58kUBybDgHso
QqeuvlCRQB1uPY6e6rO5mPDfXHv862CoqRVyZu5Qd+1njz9djQhilcgfixhbDrLw
auYH/jx0vlX7TJD2QWMCkvoS9iQe1E0tqvWUs82VMGMyZFXKzuDSvl6N50i4G+Py
7mjfIold8WwOsfirL+1dIJIK+VLJYR4eAYMT9GnKVSi3o8+OTN8b5uXtp8SCvr+k
7pSc44SFvQRiZ798+wPHhOrGbsKPP15cAhlv8/Sf4V86jmsuHMgCOQrJTPgGUnKR
DZiACxTcqGr0UJuL4r1Oznj49Whmsqjn2+2G+aHWKqmTNTzOdvP3AQLHFMlCZXTv
xUANb15HcTOXCqVtIx5yvFo/eelYYePq1e7gkwiT8noTNScYqMNsWk7rcqk+M/lL
bVMTgqgEV4/6WZiI+mlT2HfQE+QeFOhl1a4puvX7BHv9msB0nA/fWH7rThgEcUpj
XWnYSli9DiqpllvSEj949qdQcS2eW9pTDJazi6hJagWrvRQLlHLcIcLNru/QpcQ8
X+njqKonofiC+z0SnsTCbWINsUPq8LEXFLoZMN7a4i6Uxr7tduBhKUj7BkU3FeUE
nQGzC6Y0sn+TOzfnz/ZYKDaVJouJgbGiqgFWxSgm1+mctvc7PMLhL+mjSQAjwn/w
xJyvzc4qmgt0HnZM6bw92J2OOo57Uerz7upw0V1iz2ZETBiUiIO18dQRn/assCK5
DxTZ4ozjxHnv9DzOwpXSL7DhyfpAvEW8RTC5gCw2SRMCgJVv+Z0nEWqz1QGM/0E1
QecZZPobkMjV6Fc+87zYp5lPk7YCAzjJlz5NblcMyVwvK3OAn9Y+kyLb337jSEjF
WaFwaSt8UaeCYq3Y53lfTIO26KIE1bKXCZfMmNzSQ/0OBP4IbWvvCGPSxQwNIxrx
0SwiofT7TQa2j1hBRqTCquEGT6jtYryc+6KL/nVhVVnvIm6Hfxrh8YptgAevKhJc
sEpXA6o2qyn4/fa1dLVuyMjwOnP9I8+FA/n+3tHzrKRgPRrpIBKAh/bOE77k7vFj
SFLvOxXem1ZhsaEbca1jrIpDjtH4+mJHNEezWcASUkIaIAGQgb+0uUFjCiBbxncg
E9S3vyJd3cehSym3xbH4AJ4WNWjboRrWGLoGhaAB8UV+iTE4bDcYIm/xZEHJtNXp
nXsUaPNg6Xo6ZEbTRZA0kUCMgH36O5e2so6labcio0O3mOx0hi2i98YviJE42+tW
KX0NkZDyqynglAn5xfbbTDUtZimrUVLZZgVZ99HqHsWwpbzKazjs+p9iNElfsaIX
xJTxqN/ZKPmrCzmD9RQbg77U+1kcRins7rgNYzSEmgkOa7THvknBIAP1IWSkfGaP
gOgXOLZTpY8YY/I5ulmsf4HBLeFJlEImBMiiRNpPk7edy5bUHLxdTJF/ZzL4Xt+q
tGrFhVA07DNRgr5c0Tl7g+gIxooDCaAF/mVoE9BmySM5Z/4DV1B2yj4uzcsrcvzA
1OhRL/SnRd6C5PWohCak92vPCi9t1p+NNpk9NpaufKMamXLgK9N6deUW5aRcZi+B
JJ9LAPEF8k4rYe87RWesylpuTfzvKMWpS1zPM0wwJzcwUBe9DuLk6/uNQ6QouFk8
wvwqNsS3czMOtgbCEhF9wiAPI1cMAUy+Sx+BznUbNBC+KZT/CGHK2GhuhQi/dSCE
RA2sRSExctjsJhXgOY2Iqy/BJRXtg75WS7oZ/ZfqNebHdTWRtCKNLSub4Q9UGHNW
rI+tDL4+heB6RJiA5M7EE5JWnpkr7wAz55sfArexji3J/Gtc6eaHXntshBcAb/Ok
Cq5gy0cKiJlrnumOFBt8ygNYgl1JlbTheAWwPJggdJ63JiUaa7OEbyBQvl8glyH7
MoF7pcf6fIRbyIBNYuBIyu8Cs6GXnniCzIVfxmfoYHB2O2jQvMBeCA/UXsXkU0Oa
0xS2BcerL/HIGC9YTDDAogmPMTyuIggqG7LtqFU2/kTlQ6jqXJ2Z3Dv8hXUZgeou
ujf/2mjWgOn4d6FJ8+TBq2o1aTzo+ca8rchkVKfSFg0OgANyebHjS/8mQtHxLW0w
YFn//aoIEymyMs+SalJLueIFJghxQoVBTDp6TGP7RapwWeHyzFtONRu6U1bSIy/r
lZ2Xfuer2IGVeGeIE/ObGnblpwDk1mdm2t3IaCzyhNpTNJMfx+6qpawptUsLqpXN
dK5Ke9VeU/xkj3t7xygHD4mv5GP7APsNUzxA3TIYQZBXv/6Yb5g4FsjSeI6Fdsio
sIt385kxfKcQ2reQAM3L4Gte7m0onz6sD9FApNt218Dny6a6+MCaeBkxzA7YX7xR
7tWkPVoDwYVkb7Kj6tI/ooF6a49LTA+Sxr3E++xtC7qJb/1Fqpqa7/llzaUQqW/T
0wC7LpFqSfmDZ5wck6xR9HtYH6F05bX0dK/88dEvAEcivPK1zr+YnSlcDaVhqdyQ
4F6KSJvaB8r7TmG5fWjMVyR8zv86nmaFtp35+Pt5K0c7S95qabargv/67KVy0UCG
MUwYKeIQKy+y4DbYwkPbKZu+jbAB0RF5pc+rnXj2PxI+46TwkU4cmEbQaF5hyI2z
tOpa4dPMakU+eH+G6P3txDKz1GRTimBeJZCwY3UW/gpqWl20G9R/SUZXt74W0Ttm
CfHb5LiJIYCBrK972Ksjo1Ewxi7o+AePPogzuMb6ZPKrjUXwbQdCsdHhUG1CcfkS
Ev66GuCMVnLg9gyy/zINyCMTC8oV2+8MnmivvhKI04+GVV6bCl+dxpuEimIxaKvW
nu5ytGnybIGRSv2zsxYnqR+enknXFQpHyHF23h9f+BvESpnltQwNPkRqWR6Zm90n
cqihi1//fke5AdYZOEqq85pU4+yej7JIWVDsEpcxkFXM+W5Dp5biMoJAb/XwWDrl
QT+n5dMTaloxrBqCRfO93XOaaWLpntzrVhyvaq6APH32xrsdS+5mFwkFNs06N0Nv
PxD5yuus5EUifctLg6o2/DIINz2ZX+GxXQA7vr91lSWJvR1QyJK5wSZ0vhwofqFE
Gc4oUaQdPjc8zKGawqLQBRNLNkM4v+4P6OGX9wrhC6UEjzvyA6c1ZFJHaBGhitmt
+VNrvVLfMjVB86NudQPZ6LBhFAV5sKQHBGvyYy5ff6E4lAjebBnar6/X7TfXRsq8
6MoW605mtGJxCcV/Er5yOMB0nhbU0rV/OQSUWhB5I/n045mQLx7o+yrsFKMd4WhR
yIMleGnuAWqqVPbNJ6HbUBx9NskEL+bkPgfRbPg5L/zAzdq9bHe2K0zm15UNIc63
yI7twNdptCGkf6OD4nOPzKUR4rsSOoGxQGTMHuU/xNCYivNpj5G0iXcAmTeDzHky
ivWqEyxgwMexWBKX9J4x9dspMA0rwYHPVgeSz2cC3Cnd9kLi0zIvmWaWDHy16h3Z
xCiWzYR6dp77dkytHObb2WqXjfkq0Bnio58yrpYQ2GUl6uQ8TYYF56vbhDlKnT1p
nhsYoLhvUURDUxC5wT2gV2VpEKzhMkP7Rg8tvw6Q+GJMi+ZkC2MOihW5KsNbr15e
eFqqPkTAdIcLbxwTzl1GtEJgjc7AIl7qFr7UHRbx8BrorxvE4yvIBVnrHWqVXnPz
M2e0LhJ7kwUr6y45+1ej1cCuuCF0gAaaomdqElDIoWNo3vaeE6G7ZipcKDNLEspe
NhhC+chkIFeDFIC+Vu0TWmRcwYy28Nwz4x/g8qe3bKnSRVOijIoWiIe3tyirLOYD
xeNyDNoEgfUfRHYIklkdosjEtiAgEep1LF1Ilz1uFbatvGwS2NFVBq5VF8ySHZpt
C5lesoBaHGKctv/WVh6DNj5dHStWKbAZWQ2BASbg/YMlB0B+1D0dbp4ldZXNpvr7
HJ0nFsXKXo8g+noFvyyDWeSqLggcn19XQOLiyp6Yf6RBmJrHVnCyj78bjG7M12sJ
zC7B/04nVNkHtdufObkf/ge8LXRIL0kr1QO750NQZ6k6VGpyXBRWsutpVeOuxFRj
J2iqkRd+6xbSSKxy1DjCSJxU3pXjyEIyOSn3/NLKb6d+AHULL/4MKlSikJ9SNwCX
yxuvjG3LdLnyAr2qTTE9GnnCHsWuFDzuuqRkWeotbRlZzV4W8QlFqRBJjV49PY8a
UdTQ+ZvqWxzx9acEOBMZ05NMK6jHu4WeOp4qPVyGStO6406ejy4amL+hzDdJ1ty3
GWU+ZwJ6g5ApMM0E9FKIhZZ5urNc08GCRnjfayg79Wk4+6cNc3ltOa+7gc+kJ5oO
T82kAXHkQT72mZ1TxAvQrzijSu2hfLEXrrZrPfRr7VSORas0UU/ivHruA/O/WDdG
yaFSjEruuoHVN6W8C/CSys9pJswCTlCOgjdTLgL3U1EkkoXtVvsxoD4FGZGo4cdf
hgwznVLZGvNCNV56Z7zPJpwIdO56BRM8dR9Ysknz69+mra5AfJ1at8dOjqAHMMfF
2LqcUY7Zr74Gb344vuZWQXsRflD4zSxJ1hJw0g0+OJvGXB84cRmqXSQaGpsbdzlf
+YZmKyPaGHQqIOMQz8MCBvwtbEMo6GuqQhoOrzEUAJQTgxQu/aKRPgueiC9Jo1PI
72hWOb1TJBfjS6elclC5XyEFVkFqOQntAhBCcr7PHadIZ0sn0qq0ns+N2CRy6HmS
sDuyXnK7e81VJ6sce4nyzqmvvv/779ZEFsFkHLVVUBUpruifOWuN5OWjBackqfGh
31GmvGmk6tJhAe0z+fudYQbx+FhdYBrW2WuDLQo5A+lCO7iAiBhHe53T82NDb4K4
qs34b136ybWb4Pvthq7d+fOK+Xc1XtmApfQQKwIxcv7ADxxt88ru1ls5PqCb521W
sySz4mSEGMn7PdQSYBf7lG8FL/5LSZ3bksxbNjUym+RDwVB8pNfmH8h0+6prp5Qs
CLZM/KkzewBhUeLX9JU6cheLgxGD7qJzzkb3OpiJfSuOn93pokg6igrZi1711N7c
y7uSIoWookGOrnbc7H4uRRpS88DnunTIcMYq3nS64f2rXXF/evVH1LpuSxP5CyDn
s0ZVJgpKd5/jOgevHZSEVyFUbQhCWPHlD65Rs7syCZMpvvfEdcBjZrERr2jckSaS
xWAPo207hehHkte/VO//Yr5H4Bgakomi4uUlKtAkrACEvyLz80u4UaAEHQHAlq8H
bkrhHKK4mJWZ3W1T326q3UayCOQHwPCBe6s2YggiNnvbo8Hgt+nO2Oe5t/trVAF1
+wF/RVBaLLcOyKXFS2Pb8nPbVf2oTyJRBBvihYOqOB7M/q61EoHowPPvSjxkBiNj
dGJJvH0NzHnEfHRwHvnnqWlHn2CcVvJ6nsgHaIsYjvD7QPjtfRQdJnTnfphkhohV
49qTyC0Ict30y9utNjgH2OpudGdx+0bJ6Fn0C8uOz7JrQzcmIzBptAhixn1J4OCZ
brzeUf72+rw4ByofuoMGFWJRBdxzlsPoHhmWfRdVlRNPRBeljp/Q9e3DAr2rokzy
wW0q0xmZelfGf5K2ISAhWRdIV9gAfZ6U25Vct5BnCBshRDVK7uzptCfe3kflplj+
Lei/nj5g9WodCiTwJ2nV1fIzntPDDGP54CHY+SiySb1Z1cbvfmT8qD0fxuX/AqD8
88JDKGo3/VdnaDzES0G73SgZEcrQcNA/kmfYXU7ryHIKhrHauLZ6PUQLCn0xa/PL
52nQKcElMugdp0c3cUTPsb17nLtY11AbqiswALsMI12etuhYdvm/FZ3OuBlNJvu6
2vOohvjFso4Mylm9fpIw8WZNSfhEkfLh7bdlmP21PtfoaEPa7E1faTugVaE9CfTS
ddzhwAyeYPP0wha11TRS3di3b59JXYuRjerhU0jFKX3QLSImJ4eFSdTgyD0qshla
jFztl2NqUZsP2G5O4WY6rbbza/JiFKPiieRO5ANbbiBc+MtD467eU9WM+k94ZIWs
rRTVM4Mm6p3mHEbgc4TSLD30hQSMFpr6QDK8zXNEUy3tBx6RmwaL8bYLulGB9phT
8CkWGOaGQOI914xBWJK2Oqj9dLzNE2whRL6zkdsst77bjX6L1SDwTZsWgOClsLwk
/rT//y9BJeXk960DO4BNQWK+eRlMn4YwwbdTLjAOJwS7Pex5lSjdjBud+wa4nXVW
EMk46jLGFkQZhj/Av8vM4oASs+HVMPi/+9iIBQgEiuhl3vSsujUjf63xyvBjXjn5
ylaMIqgdK/IWigmVjOv4ZtDsyfb4KqSz1AKiTtDjs+F1e4apKP4w4eCnOSCIICP0
iEGR8zC63ZqjfCGc5ArtF6Jv1/uZXj472MhnTf9jPLw7gFsEbWripz6QYy2WWLzZ
azQn3rgPbzPGevo+xmIOSnCbTuYi96FMoHPlOrtqQqRMKNPqSu7CsxXCw6i2Ci35
ZughkMVsp6fwrDf/i/3AiGG1GVzAbNoIm69HJGEiCBhE7i1wqOEkO5xUpUQdwHrB
N2WUGi1Eh+/zdOfTvt3jsyb40aTOckTZW3pvUP87Z3+j+fKTkitBMrib76bmv0pG
Bngv0cin5xlEk4r0i4vkIYWsTWPITPdDlZj8XXzGSHo8dvo7LJCg3soF8g8QyZBx
OhbspxApYoMU28tPEVj2yZDEhYzUsSwBoFtBnyVnL1l54uUYlJS2Om54kcFQgBS3
XbiTbKKN61QZD1BApWYKoCRAlEV9rmgEVg4xf4cFvZQG6/CO1Elbsb1Bdkbb3rvH
pndq8KjnkGQbXaFlpIRKwb2EMCjMFzY5dHQlM721YGHOyS6QXsdllzi6FcNoPyHg
RolwJATFxv3ud7kDrz9+83TNZUJrB89fWPOmlfZ1Ny9pHczJKO+J4dy+tKKRAZXO
Sw0g5lOr0ztQu/qPQ7G/GOmJ6CvVj66fdege+agPCmd9HCYaJm10gY3cVaPXFcVl
HsQknPJ3BWFK0/XThPEnMn+QJ+V8B9XawmJoiYxy5zi2bhDVidsQkB6gp4My8Mtl
xI8K9L+NPvwP9eU1Ykr4jyVhWVm/J7ho+Rr4BJk+RYnsA+SfGWYBDBcsSkvjsZjL
Qb+Qv2rzZ2DEOwZhDUh+T16veEH7vdayN2BzG/Qe6BKTzufUJz1D1HtPiP2fNlXR
F8j95UqkERTv0VQDLfor4iYIT6XrZdnJjcZniFBUo9OX7fsRhFfXLsUcAeZgSp3+
JFP5uZpDoZB5R+EThQNi4J2blTZDJ+XDa2SiirQUvn4uJn/m1DRlu3yRnDs+H8Th
YVi8uGESc7fimoDecqMPBo7j8pWFY+lYScTJ1/1YajQiHNOcU0/OmzvrW1LhQNeK
uBbfDHlliktRDTY1pDHQP5jWqHXmO4IBpzohBeqT73bCvV0u+oQwKW3AptxVYmTb
au4s/zGg5nrcdM9Uh8/umZhcdftJKOME/hiCMMTQVD34irLzN1JJqgubs7Ac/gzV
XiJsyJO26DpYVuTcyHKFgiVH7mrvgcuhH7ydkIweSfMWMDBPd0QV9JlrRA0EYKCr
8EdZcKwCzmDCcShOC6D10OAO8g+rw/Cn463eN5gdkOb/7uU5CZ67helkgexuh/M0
r3TXt9far1DD23d/OfNKu5ZGtXhWhf6Hl/kvLEPFL71PbBvdQU1cOET9hpJBeFLU
twAMt9eHPXkgnFRNvG4fIDv0YZGj9Xq+QCWGrK/FI9K9zY1w3VHZUUgxa4lsv8La
g7LI9QV3NqU/4RDu2RgL4R/+DE42/Na5kXitkccmitgkRhQS8OHLvzWk3rB7Ge4i
/LLJYDx3PMkFm/G/Phc13tbUk9l4DuzOUG07NpNV+Xnba4TEBoMfrCQfAT41R0TW
yqqxIqSi36DIMUgL/roVQs+xzz19TmNrcmXiC/OxVqtkExrVXMzSv2XMu0toq99P
/KD484UTnNWLEdwxiPVIHMNgCHWn+WyycCgL8eXhuPbsKcEGxSdRCV6bc3R6j+Ux
70uP9xb3h2QJVtIoxAD5s7wjTTAa7jJvbTOESHvPoLNA3M4Y1n3paWplhz50Pp4d
2Hp/7tSK/B3Yg8hZoF2eaVZ0n8K8T7K81d7CJZElH6qtXy6Fp2eMvg+3ZMQqs4Vh
EDc6aCJAZtgl39/yTn4yygm9ICl4EbjZ9dgddviShZR7w5X7qPouL+x5UdevBA4H
jivsbQ/usZ2jYYd10W4mXpF6XJenytpKtQEkp83crpkRSd6o6sZcXDFBFg5c8Cmq
y+rMZ1+Rsh9prJJNHejv3CCsSX9iBMLE+Vor9QboIamz+PfaM/b9+DN0cdZ7r9Dh
k6a2QGg1MquZtdUC5lG0WRh9g+lRzR8/J0JQyu88TSMzRceNojxEPzk93vcslvOy
9B07U4FfoZnHL+y/ktrBQOX4id8trsqznWKlfR09kGtFua4j///iiVqMyXIpjGgG
F9p/yTtiGSG8houRdDXkMvyqMkm86/wxmheAADT94NSrQhlzw4SLONprcZHL1ehL
cqeiY2tayc434vb2+vv7KdKVNKWMIfXBSCDr39WPPG9K8g8zNkItUrSDfHZQR/e/
2xRpKlUPJ0tzmZFc/Kk9C2gbpSMRkvfxHpqlKB5wcRsxKrCkCFNzqtlDZdJKf8Un
85zRYulLKjG1TLRQe5oPw9JVdS+GQ0LE9kFavw2GEd/XQ/ApHFiSiHVFiK+Hy0yZ
/xDoAwxhdNrh6HIQmUfcgt3ISt9X53b9R4dqZaGUAAaRwws6qrRzODVjUOZm2cii
uRFMGr6ARmaQppoLGeTn4JW6XAyyO0XkhugJnNPOIC4qPXuXNJ5azRb8iwQGpHPG
ttwH+9//br1OinY21kusg6GIVLvtXL61HUda0qyh5IrZHPEeVKq8k6zPyv6r/rvq
idPNN/r6tjVN0Q5QsNF44XMT35VqYMtwNOz+Wf9iSGVoWfR34Ut+DXhtkc4kSbei
uKF7A5+vRhCPsl3AuA0gbEr4qGDUv4vmWtzm5ZhdgYXboMj6OVITLPzmkrPU51iY
YThT62ciqrVDXotJeFa660uZDW/7bc8lX29zbNNMdSWpZRJX+czh7wej6/6OFyli
X2/lPBphuJ1yWZoTUkUO1XvzlC6XhGoCaQs1EeFw5HqQAz1R6f4zvvFXH2L0OXRK
bNkaDAeAmk7H3bpHntYWaSHcKE8LHskSnVtxhDBO54g4Pfu2/+JQ6ugGHoQFf4j7
Z7jWGnGvpbOVUWjIrnF8NM1aXGimmGrIiJ6TbFQd921LxWSii+YuMHKoY7g48/am
x4wlG1QhZvbZQefSfeprczQY4nvc5sGP338agxg/9o+JvFmUzQwldgmhrlx4n9ol
t/UJkiP1xnk/a9FMu/JeRfUf1tLKwnKw0498DjGb6W4OYC4lGRGWLfOYTT9OsY/P
DIM7Z8ygrYQk3yh6mN9cxp7ZX6+Uv06iJ8KTXcPkSVlEKpzzrlqLT/F1NWEBcBjU
rAPpQz7+dbndsF4AjkMh4qVU72NO0ShJ7ukxWzF/n3spEFiP6eUA28vAgvx+uO9i
CV67oOeHhxTKyVbdY2x4keM8jcg156vSKOJNeuUK2PRzSMho8eC3lk/YA15WDfsj
fmBuzjW4q0rzOy1DtK0HunArYwbSHWAMDACTKkJePl/D0x5i5o9kLISVSIjJFnlQ
pnNA/bBfqjPaXqhCXWVLWI4EvSHZAMR39pbvBm/HHo3T6sTGOPJU50D6T4vWrfzD
Apix4fk0dn3DKribJ0l6c/P3A2GEesEmEwyMpcsVhto31DfPeoDobvjF+SHU0BxW
Z5V1knZOf0qWq8R1rw7PzP/HvFilfEf9j7R1rVTKM+kjSqNhqh3Rv18qnC1R5o5G
IOM9umjHnDxoL6aBu1mDSx4ZPNIUqXxcXxvY/nhQHSt2kwF4p/zxMVJRpiBO56x9
sOTGTDDXaiJXaZKfzUvXNWkYaSfzLk3US3H0OpahnnVkBVMdXlVHFh7ZLxKhRtkv
Cut2j5lAgLSWBUIv0dFPY+KYOrm9kE/E6BLo7wP3RhZNJUC9O2xnbHKkjq4r4fkS
ZL8jKcli17Ce6sTMBA0DyoYRuLHjCp40YTEz5n684qR1OEBNF0IndYOpcs0mEU8n
ebjRTUoYpsvgWI8E3xk92a77wSojqFDYZynttNfqTMy7VFsiT8LPbl0Rp/Ghm+BZ
7FsW+hsIIVVzdYOl+8usXWArr0uSX+2edp/Ppj0krVKptj21lnZ1keMGgZXzTR1w
rWvAbZAjZogqXHHnATqDihQXLvLuEneQzLdi2JWalchML6DSESWeSiaNKt6CqT1b
Hwa2vjda7ZwWjDARY96pfHUpODpBlij3HrJQvlKMKE+zHFXZBc2+TWaf/yVAcpjE
3YStsfEE4TzWkTdyIAIc6Pz1BB7yR1bfLmtYT64TryV24j6OL2TpwuWVZbiSFOqr
PhhxcBMKYLtID0rWHLWsKNvAckPFR6LNzEeFPbBcmDxZ8tdS+y90c/Gmul6RZuMM
Rtli099kUQwJuZZVxjqdQfCsde0TwfblxDzt5UTOy+lWFS0n0J1jBrCrv+YCnL+G
d9AIxdU1hiW9rkO2I89CZlfIST5sbmUIyIqGwcDFirzOHzQJZXP6xHSM0+oI2pI0
PFNqAogdwJIZj7h/u2YBJA2I/hV1JfZrcnh6hJ8uvdXfXaiO91SJVuFNxQpOST/6
KnMS9TW+yHl2e2C/GVdjK5BC9+9XY4DJKYgo93XhAHZbb8vVIuJJUn/q6rQwe0xd
L9QSQ19fAOibUVJ87rD5g14mbTqyQuDNeBfA1Y1+1bXu3G/f8ccQs7RwZ4SIKcA+
c2uaE9TufPNKigzhSPoUP6la6UyZtmXHW0IV8qLXrcM3KB+rCdGLllQlU8/ysoSF
cRwChqpdbTREdbK3ic7USDRGONjx4lck8IZPjtY5chmiUwoAAXrjcgNHtqMdP8nw
aOLvrnn56eGgy4KAZx3z98ls85upzb/kqVTMqxIKlSw4d0SGCiUjEmga3bNbYdrj
HotCOaTJUPmWupKCaGF8ag6zKqEGSS/twpv645qMCRDVhbg4xt7XcKypR9DLfrqR
nxDwPCOFO04x8tzRqRghnMkhB3nUJMfBztMN/Z+U3+xFbVyZGh+4Eq3uFtxlkLhw
tF37kk2oDtMf0OkY9e77scVsGV6a3qi3zGJhBXrlSyJRUl4ORGLgO9SR7O/mEwmy
2LkjnWak1mLbkGZw04pX7iHe8+RPd3W0iqRweo0NMN28SA6nCBHVSYHZ1hgp9gx/
g8JxvuuKz3jopVeUD8sEhFFXkxclwpWc9nDxA4KaFE2H/UDc+psYabAmLh6/NDR/
khGgxoRD149jQUaFMkKkkn5ctSurF/z2UX01JfwhnEI/6PnZhizbVytcBYSnRH55
hzjY8fydRQc8S1Ie6GUblF1sJcBa22SnXHlY9PrKTZ9Ilq0fN6qnIS0kcxIqPpRQ
3DNFi287p37TrJ12x5cgx3fXnv3F/VWImTQfRf68R2cWQru3tTkwFjihPMIvmWv5
kbgLA//NL5G6hvDID2ZbPrrthgpkV3kWjeR2/F8AHBv6QR11gm5lRThVP1CT+u0S
5x7MmVvVUDT003vUS5y3Z7Cofp6KjgEO6Ty5w27LjVRCqxJWiZb5/GDm0Dve1MXb
3erX727v5OLO5SHjmAMGgBhjWSQLcEHw9sHEUrs7dpRSAIZZ0dTkf7OD+eLDtAf6
WEHlEHhY880ZLiJZjtpK47akITQOLgb6YY+xJAvdNjqITyAl/80kV8e/F7scokh2
upEzKnwty0AtYG9nCqY79aLf+ZbHmwg0hyxR7Pec6xYhIdIK8JWpAVr+aL2/0/IM
/Wsb2KOx8UxWm2AgQFciH9KeTkYfRlOyv1C2yZNfPDv2b6hlLDOVACgLamt4tj1o
0+quWhZMlwMYcYAGc26M0uqoEVbLFSqUsAWdHYlscrY9gO77nXzZlFkC0VM5A3QA
pJSjfAOH2bJngihBet40UpS2Kq+ViMGZeENgBa88QmgC7UAaiqY41ydaisdWTFhW
NUEC9nw/ICXhRhgFm7Af4+g7aruA22xKv7WgOOQ/+TAmru9r/A3bWqLO7eRWpQLx
iWaL8SfqdeDgR7pS+iFaJ6gPr6mYc4uxFjzCjMyzZ5U9/GPUQ03FQk9V2OJ9zTNR
xUU8HHc8K2U0F4RPldvah7a3xNbbw240twslA0B4IJB0C5JZDq/k7MXIzSvJcH/h
AJzyCnb9AN6YxV2ML8OpXsq6b6g4u0CzxelQYd1gqeTtf+tnfkgB7YKcnTMYzmpY
3CPncdrR8TSZxbePrOS4tNrh/d9BmUpNvAiexlSG3LtySxa9ugwfIi45rYNRSkaD
9ZHKRHUff+a6d5AvqOJpdsprjQKCA5VMvyKHeQuMqrIK0tMCde0Iqq8IybNdkUR2
H3MqVKabPaU9S7UsfJs+A1lytUARVq8h8E/Hhq3uDhryyWCbn627u0E928lc+7x0
J0YLDq+QyXcNOOmSeOOkg9RdSgdQY23nA0riUfWeWKmQJ1AhClpStb814QfzG4gy
uaNCn4S6dd+AFP/Qxu5iO07127seJEmc7x8kPmj6BsBwSUVRpn3Mqa1fvx8b6+S7
/RiMhmLU24+jJvExa9X1JIpIzcPpdn6PE6mhnQQ3YKT77n3BAUTxEHEMSiDkPpbw
l1SUnozP3BEHtZVzMdiwVAvRelC7Zj4qx7RTvsIGuCIRC167068y8tftNT2kWnqr
A70cUBOJ5zJpY/7Ey9OdaMS8f8NQVba5peULqSaouafw3bGQE+QGHonKd/Sd4raH
cbTaVSvczf1W/OaykNzLIXy+o8SVkbyFsUcoxUEs+CIc9QnEY+G7wcjKUiejqCQF
8Artu5JxPZek3FfRIwIpfB2tGtlK9fPINnt8lYDyRbfm/8c4BsYbTAxg+ik+iBr+
L4PqBzOG0zf2hQOVuINQN1fjnbdFDf9CoSTSBH9m2XfPA8MQPIMJOM22ZX2MgmNm
D0O8astPT8VBS0EL5A5foh5Aark0SbhcHVlAIyr1aqSQ3PuBA/yxJ283wt6JV3k4
Poo0vNu16fJFm1qOcC6XYSOuiT8Q50k/7eTHXfsnreI2SNW9KTjUoGduY2id4ltE
Sp6GcpEgr9zb0SK8xAqushEyWAinJpQBDgrArDgYqGlxqqvTEUstSIQGwatXlMlR
5+5CeTUiMz6oEK1YNyqwYBrxBbIm6cA8KRblW1vg8WImzTqDWNO4EC2KoGFHQpmp
lRKJnUKS66n/COLaD1X8JRHB95GEwv8nKMfsflQuCoFtDguUeIJoZQhuyPKlXAFp
pob6NrElSYwVju92rm9jj9S5H5Zec9wJd3CSpqIK6tgm8uYcDwL1Fx7LPyBwHwFs
9ev062szuq8ck2MlD2SMWUa2eQIUGEk4yKL4VC6QF4hi7zuARtsh8yMAo4yFVP3E
+Z5YogSekGt9A5T3hKKtg3db9/kYeUgmNX+0/2bIeXfOCmEhm5amPXDU3pTN80lF
51EoRGUpArMMdd5myw3NugVDJ0gxnhvj87OtNseaWJY7nkrYG/rWH94bwCdPkL8M
+g80fA4VhGi8iRcS5SxlEWBiJofACVBcGaho5vgaxCUEGfbhXOkyA/7cuMpWWG6q
+qLpUwgclUofmhvnmLU7xTvResM1JLIoAQAWkUif+tTGwQSf0Qtm9z5g80lptdjm
5YIK+cq5UCUPWFrrLovcj7kV+JSSbw3ztOjO+bepAUxTmnoqVdU/5Ce5ouHbYw2N
qVXNqiMa0NoQ9CEEihT1WgUhvLVfPwDlaCKVgCcjvRW66SkZ07VO5pZ6SC7yaHXN
GGMhzbVevYln4pWBEf8V6oqyPA6g8PneXmfjZAY8A76kU/c8C5QpezSAHYIMRReJ
Y07YIsSR1xw2vxJ2Bon7XF9p+fu42mufnHIDcvIRKDBZsmYXafsd0r04gVwMxkd8
pktkrPR7z5k9lMArXvHfalgxuP6g5qYrKRjVhM91HLGgVFIzrILXiX+K8khtv/oL
U/eZk010V15fBc1emr9o7sbymcTjSOF/WAcJ2EEQD9AUwF42ruKFoQN8NhdrIT1x
LpSui0pD7iUHdxSwCpLK8xMg6DXf5iFoIbKZakiyZDQrqJhW1lXeyB8cqIcxpwJg
EoSl1iPy1x4+68qmzG0/UIC6muSS5y600S3nUPPYC/PTY5FN+TjKKKLRs0ccWpDi
P0p/6zzdf4q8dzvfGTqaIAb52De5k6eU0RgdGGomF89k+Kq1NRObKyJQGVMoOkKO
rkZjzkxUoDjDc4CltjPEfjdk1DntIDoSycONAjs6e7DcyY6Nrr3ASwRw43Q0CWLv
iML3ZH2t5yPEIyRCDbs7TZ3OinOQTcUhI39XU6TUMYPTFfGomcTDJzjoKfSbOC0F
t9wIlJuVUULZ0RZf113TwOmTM+u8YgE1j7Z1wmhK0CnIzpibwHevM5CnIdcMeBVs
dhxA8o+h687nwfnBDqO6oTBGnTNrCYWDxwDJbWYE4PEZdrLBZ9nrKIMQ2HBKAeBE
Fz1xEqckgBb3QV2EdfSXqeIG36r/MxnyG3CuZzMQtAz+dAY2gZR4VCCU5xU3lkEK
ssOfk0Azn8WcWSMYKEyROa2S+LM5eXdJPKq+ykRh4al7HBC8X8hElHS/T/L9ZOrV
Ryr1G3Mj6QKziIvnu6ie9k5q2xJiN6+1RLRa0/j/oX84xKo/sUWn6/IcuP1HtcgZ
AK1szF+OLKhQkop0EPYgVhu1jKaIGmPcbHCAbmJk/9gwxBad0gsRTF1bD9B59WZL
oXvfmepBq86IcAlFa67TC/Xr5W2NRleevHA5zNZQfpmV2v/RYr0VtRF7nPZybVM5
1RINcmZHMmrqpmP+mlPdElg+Bg8g4C75iZFM6nbuD9W+fvX5Pm9IK17ggLIjD+Vt
7zyCvpsyM729w07sdzFC6kZvjMmigcc2uKv22PPukHoZUh3bhEB3lto60RPA8WjB
HMUeik6oReXom5U6IwILGa9WMHz65kbqdiGhBxVzPSCPKYanjeeqfwhZvuTVIcVu
MU5RUt5607dZQ78M3jkkW0XB0sOvluqAL9XDu51oB8soPK5Ite1mIQ1Eru9jVEur
9R6X/E8IjSuHQAdsq823dioUnOEtb9qDU/pfAp+wBbAZDe5DhLYyx3wf8rqSeKNr
hZH81Jt3QeJO+KX5lMFBV/vT/zSE5kNXNzQsahK8iUA9Mo+gK4K5wrs0bxOinVrE
QOysUt72/G2w4OUplBlMLDpKAXlLwNhyUoFtoZ2XRaFPr4R+anUQDWxtkkR07aiR
5SDCcO4gkQAkHHbThU6TFzKr5CmXeRnmOtrAT0V4zX0F0ZUs1R9fDnW9jYws1Fch
5NhEjrgNz7lhMIy9sOyiwWTGNyQWItO2soWwLhxDWhG4wwShfF878w1dytWzudmY
zfCjIJkCEYa/Gj67McTCPm4mGCqchcBie0LtMXyxk5x1OySwScX6vhNgrCyXFEMC
3a1zAasPcBrClzaRJxMB3xW007iiB3/54ljZiZ4HK1gYQiZut7oZjR3BGEs1hcQM
R1jz3DkcwsIGjlm/XVG/C6LGDq0zJUQDJzrCYqJidlVHie1iAZMjtmHv7cJg4L4N
S27Cx0hW35JdARffOfiIs3KAau2IhXCjCsxrYFQHZr6MglrCNhbeHb7vV0xL/RRE
VmFMTIgwNq7kUMi6YVz4J/vdZLJT+ApBHM6DBbyjqVG/3GXGiAOT/H6mIS+UBcEI
El7MYrzlnYpMC7PP5k5S38Ztjd5mvHxPBmhEKTUsXMoxCHs2KBT6gkhQLwBjiLD6
0X8GyEpBdYjxRjyhS3Diyb4ZvOEOGah6gaIAGPvb5mpPQZhmxyiD7gQecQRpk6EY
vdfzaora9rAD2nFB2XfuHaAT0AooQR55z/2/y37t5pFY43GzMSnVzAPv2G19Hj8z
sKPU/faIHLhVPOugVj0hb+XFPLCAgZEstb7BEXPODSCDFh3zIkCfiaebRQ9MdSWc
qT9okj7/6yEMpJHqlVHx+iDmKODUfxGhTNN4j/a83lNHKoG+KbvsiUi+uys8IFGm
9wKMuPJqdieBzdeN/wEd6YdpxL4wVJP/+w6CtTgx3Vt0ssg2AO8CgHdGAAl2wUq8
0DC6nJOke8Qb02cMVsxRV7mToTm4k5CJv5SHg3cj63fHU/unPopUIYHlu336CQds
i5VDGIGGt66I+QE4xlW2WrCOvBhJNLrlX082pS/MCa7W9yW+o1MUMKIaokfag3e3
YXQNTbxbrvSMQqyGy5VBORh2qQmmU0WzA6l1BoEWj/oXy0uiHTUuuRPVYljkr+MO
BuXy+wkf19NlG9L3qv7gTHR1+JfqlOjCjGjF3uTzQDcGylnOhEjJIUOGdDX+kFAH
xAmZpfQulC6ClAk9+2e2D1hiS0bcKYvwHtbMA+9w9UgXdwKwgdya54UXOxFN0uyA
IG3OeDanz+heW4G/Q1t2FaVQrdhFVfuRbcDl5Hj2NeWOTNRm6gMfwzko8Yn+eGFM
pVKny/sIVlDHl4W7t6VQel7/NgiQ6J8fEMIMX+WFFe25QhG8L4jVYOF8rrCktsGX
QoVckcWhqlPbZJiXZKMXB6anFYnypDZDwE3C1yvqbiB/TasVJhg+xh/hXGkuhWCP
cNkyPmLNOxjYMmA1UFJ4n+t96Lmt/u/+DYlU3EnTDEAFQr/fEazHxbWQEJS1uq9D
tTxA7istRGWRwhB7x4O0X86qKI/Hbjd2VSer66OhAXEfzE2PzecBLOjyIji/JxOP
pYsGDNHiMy++TgfGlirDG9FTqugkD8ZbfPt/tzmL2LHjeNdmcOG+fY9yydJ9Wr0P
0muifVq34hitmmyfFE4Ei6UDl5V9+K769njxRth3//jTNFyL3O+2ZWplY6rIzftQ
JIjzB7XGYjv2v35utD5i6nIGFowWfi6uTI/4Prw11HRzC0ZxKHX9+kM09B7c9+Uc
VKcoJRJiraOvvp80SsNbDSPT9moncJOAdkprKvex4gha5GRFPEKOKo+LZWsYbF22
1U9y2IEmMX/z58Lr/4B0HnQuRM4QfCV42RV3B7tkaGqMOhpCr7WfE0LwUldzK93o
dmbp8rPeL0SF+21C2fAzsUETajkCeWGscLV7KoDeN4h7BT4ytcLcNk/DkqdUQgEO
l5W+mJvndacMM3zYBVnP/JwZXJbM3moGB2FnCUPpC0hq/fGwqjKlphPqnwRxAC09
mpibcq6MyTkwkTdCCMfJ6+J9ZHNBUVB4es2uSHqbcA471a6Bujsi8Cqge+A5r1+b
6tTgzGsP+3Qn76csudRZTaNicrXrNdHz3g2amctC3yRYR/r95upqAt4JrTe7LmpR
2kttxG7I4y2WedlBmhyh5RdvH8VSWkDH31DL6LvKUldBii0GZ8wqRfvhDmkMORUK
FpipqbtZEU3rZxmUvoWwK2qDjdRfR6LaftCZAzkpNHq9ABCkU/V+ETsmTGgEH2bR
P502sF+zupCDWISSJNIct+ijS4xJmi+azAaxBC2t392vcFyFZI1QxklcEX8aCNRS
iS4dmEvcRFJLv+aP6JniDCXx+vjscanBmeGcKN/7+WoTI0oJNTvw6MwA6v+INkbP
oxfZfM0JX8tsqJcjRSsJ5YubPTE6ONeSoC9osg6E5QrT9ccAQpjCjpuPDp2vOKCS
EP44YmI5Ya41dYTRmA2wvha0pzWySIZdRtS0Vxz5gcz0X2cLYcwNXUcQSJ1FxIdK
tsInRxZX0MuHYCXo/HYLmsBJ1zJBvLp7TS+rINJqbtWP75i1ARQ7hk+aWgTHIj9M
zkDF6gRZt5ARZflUTals0VORXEaWccL2krWLfU+octRohCHgDylLt7djIuwEvE9c
mpF2z2L1iW110LZ7rB2j/T21Z4TFMYqCi/aH9nW1E1j08Glz4S5nvjCOc7OnPkRI
KM25TAwkWSvktfUXJf4e+Ebch7CJdnqw1AcBX/Vkr5zGnhyJMo7/2SNeakMQWPh7
/aJAXjPrY1vLIn6oUfY/wPLECJBvgoze+g3vUcruyaFT7JJ1KtsjJ7vdBxX3wFOn
GdvqWoxSghwtzaEmTdSyDJDkrBp09Fr5QJGcsfb8hT2RTUjFiMwLywDp2eARXfC5
+n3uTnDyZ+/uzua8raGowcAIWJUONORLHJg/0peHpJ4xz9n9hJsQiOTv6l0cV/6t
YYGKCeBSyBuGvu5umNrkxdYMX2CumienYn4rssuej5SotIYLimc/UollAV9/tMUU
lHBIi4+rgMkpL59EsfkdkkzfB0EmbKqnLKW+vWGdFVDtot3jDxpw5K1lzDjmeLnR
OsH5TmfWArp7dnSfnevtgPfyCuCl6m/jm9a/R0NRDX9y6Wpwq67e0bqX6pkiC/+K
BvdcVu8JcDZrHkVtswzkuVALkAFigTEzssAcY1/UOSbd/JwZ79MH8WYRAlD4iZNI
F6mLCnW20sfRfb7MtIdyMSJhsaOczOOvrLVx9IJhYHNy/+ClUE4X2Fh57Uc5JJwn
0ViIetzpSUvDulp6xXYo9WCDJAbbnELJxAVEEZD47AMZ6aDn+fZfRXu2zNfEgkRx
MWtV6oCkG5Z6atsDP4grsA8crVhKfqYI3s//kmzgPmIujiexLXhJdgFDA2Alj5wd
bvYQuZYuQPRyTmM1zlcrrov/mAFI9mHwERgwb5F3doaFd/bgJNlmt4g8Qn2VLS7E
Qg89APwvnhMUMaPnUnDFaQH9hY2spQbJxJbNgE5VCuGrVkDaul4LXh7cbp+6GIrd
Q3e7i+fRJVP9VT31oy39AT0JqhDECgkWBZ87YO821jSibXikrdm+3w54vPUENFOc
22w9PfQLgh/8GafvmnNaxsGUtJ57Vyx2l9rZXm2Cfg8k8xMqEWp1wcMsOrmJgp5j
8Mo2vnl/o7e7sI1+2xNmswD+0HP/FQ1KkQrEUI4y2OWfPz8cKVl6yd6BFsSQb7th
dk5lC+9uVnIsVsJxJ1cnqFE3J59aE/aLkmi4ozsG+06dC9QJHJh2gY3wVV/IWonr
4A1RRHazoIORi+E0RDzAra/A4iC3oYtQr0SUIz25199HoHH6A0ci9/DjYz1BSnI/
WkyFIyARbIZU0zVxmlSQV4ScnSkf7Ts+EfBLBxa9lEwuW1VSbDmoSPsY35CuLMlL
3QqKq2d1rXfTuYN7x9rzCy9TbXdNJY67cHAPFou2gPKvxJcWdsjZYs0Ow2xwPRF7
bcZDMqddrbjVAgIeJ26ztmjp3U1MK9Lz0GiHpW9oZ8eyxFUR1sb/wszszAO3J1zH
e5dbxtCcNZvG3spS33l7OKpnlxiRGd257MxKPiYTz08MTHsErQ7O0EBhXMOs/GBI
8K9zyf8YTVltF2cJ3AzgkM3etdJ2Y8rXAF6r7r6/i1VDeLuj0wjr52FbbRF0+VD+
vagQ+b6FcE3DfPggTS3Tm7gnBZBPHMv7CpqKS/SVOuzkV8qPWhdJb6KI1RXxeZmD
CRw2evfGiunqBK+TqBXGDL2XzpYB2PZubSUox/cmSP0ECiYsGLUyW2bioXdIlRkh
OG01r1EhN0/XrJpKeXiR6dC+elKWJs2f+6kHPQTQ2TkA4JrtLS5iIbkbd+PSO30U
BMAlxoy2Owu9sBT6O87W0THG+LvyRZX0TQrj1Mfkc+P65hLajXfrEQz4oHpmNqhG
yZhOC0r2YaItSKSGD6uWD0zv5+4lWDVnMoIpSgp36kQXJPRF74J4ueGbsClcwiFZ
mW0zC8alg+YiGXVnlNiTQa3zWvVSprF73otME0hagvKrk0ii9pGnpY8dBZW0DKPa
0Ts8mvKBexRKiFSkVK6cisw+QhzeN7AqyZL2kBKRs87ZBRwWBkm8SeOKYe6DJJ2A
BWmIUvOX3lt4sFUhstENiIlM/PlOq1CduwxuLwtuBaLfPkcdWkIHW/oLpua+aWyK
vm/WO7fzoeD36URtKc64wqxOnUm0VMp54Bq94vfq9MiP6lxNHGWiBAORTvAzbZ6P
esK3D2J9OriuL+2xM+79GQiiPQ1AZ1jG0wOn9z0yMJMdahdtuE7jPYcW+0oP92pW
yyctk+1qdyISL7nknZgzu7EHvZZZxNa8/PdTjL0CkM38EXEJVIGodzJH0yjOshIW
PxntWADkbQ5uizj2TZIV3ZQIxwnPN5LQkr4ziiMY3dMCh5ZIeiWrqYDT5HOjaf/A
x+RUN37yDVK6J6zKhI6kJXp67UCUJ6krwQjhNTIksGFjciRK8vrxVlDjVLqKPdri
ZZwTneO42ByYPVXJUY3ghpZ3VANxTj6IiGLyaHnMven9syX2iY7l1/X2bMQ9eFdx
ft+iaBG/Ew3bT03CAqn+zZ9vERyWwDXCxvMzd0e3XNDDGZ4HkQO7pnRMntPegl9Q
Kdj3h4dULUtbJbwfXTbOaXpI6zsKpQitc8LPyVN2hSOsEDLNMCTgK2RPSYOBQS66
kXEV6S99Ci/+MKgX2unHnbZeknZlIvI5eZsiOaCWgfX0zb5sMtmTh2cCBBURGECZ
/BmkAwCd8TxcO9WN1dqqClug4Ag7fDoqsdfyysejaQJcuUiN+5f7fB4Yj+boxIsH
RQIdmUuv3VL132a2HSqGVV1E8DMuo5/BG8hz4kGxbezsnUy5NPsb64Bz3LlQvwGx
zUUlgRmzragOmjoG4WN/97ztN92z5+1PHjDrLfvXS27FtYIi0eaaDHGljZ6zlqMd
PNLQ9WewDGBuPb5OuKQOCutwOg/jQ02068eNdVww4mPcnJykDqrKe2gRzPdq53by
TLSAaDpn24bXz/mDzAio7KhaRg3eWlnvVocBPdbYPeSt0FQSRva9HvKkt9iIlz/Y
FAFCRMD4aRPVv3upRgty1una/wUdPkBNYttuXlUu2qZOZ/MuKAPE1d8/qa16ZyLv
tTXhSwqmnBu5mxN34yPc0r+JHnthr2tsiGci+eT4ILIu/7QymlfoJ3Ze6iiSlob7
1+ygP4L7jXzwwbFw+ZJ+QHQboeHaD/QqSFNOrV3cUy5XqyWvEr4pKKGSOGzbBC+a
J2C/PR8810S/zaOxzE6Cno0cy445WPpuoy+TIQ9I20PZ/pVGJeJDx+DnX8lwpeZP
DqLkHSRxhD0B4MEC4e7oyS8VW007Ttlu607QgPzD05X3pQsKdprD1GUXYQOHBuhe
QNPk/kKBBfsTHUtbaGCj+qY6jbHF4hDKwjMsyyPFA73KsnsxjdT1gkCTDUfe6Bya
WAUPQYzFfxqxrnzf7gQ+dni88J35OYkQ46SKeGPlJLpt6eLz1KxNFnZm2umVI+yK
NKxEYeifV4gKCMfgkveF3my95YTt64tqGG9Mxjp22H9Oo1L4LaDGgop02ueNAE9A
ILZqeft82vCLv2q7LNjS5Nx5H4Pd/eVJHEx8fBgmzyg475fIcoi64dPmQ+MXbKHq
dPfv9r1KOMY+Zt0W1BeTpRHwcOrUzWDI0sHObVbJgumFojG0Ka6YZkiWvtqzGMOR
x2X3+JdIjZ4UptxSfIqhyLo7JdlM1sGmSk60RJCS6RiJL5rBTkrYveQo+j5ZeDM9
M808vt9iPuhfHNy0e9QZdetO4KTFcEr+86zTrO7ybJG5YOLiwa28Czt2Tu8j89bQ
vSQA17VfpBpIXzcYt9X2V4UtMO4CQfST+KnSKaQLJRu6bEitERX7cYStl3tA+MNv
YxfrZVmh6jdhxG/R6An6pMFUfXOuwNrW8pkzWNsmLoN5Al/EAOvtYZQQGJwZNdB6
mpQGEU/Wwu4zHZGNR+pN4UnbVGqqYh7hzUng19yoFE5y+AUe1mhh7xgEaIL6+91Y
7EEVkr+LCMrKV46MYo5yUZ1X3UNcvdaX90cg4cgtfYWI7u/ACmFBJrQLksbpry8v
OAEb1KDF4Gs84mXp1COgoH2rb87KdVp35U15Jo1qL3v+lh/UbJ8GxBbmsuLB43b7
GAxqXTRbvdzCtICNU3cj2pYmWVHA2LLljnG+BiSDE8YWAoJI9fKNHA3YOwunC7T+
ZnjpQ225ijV+61Z+BD5MfZ6f21lkHcppyfy7inRd6ve4g0JU+hbKtCPyatLZLdSi
V6o7AqjZoI20m9xd08Kg0zYvmZ6oF814zr+QKi3/UMBesC2FqNmXQiwLp9az+Us1
VREx1peuesr/D3NkH/kq8Avv1WTC0eQJeWcTBPrOIW0IlrySDyYW+FX0Re0HZIiO
yJ43W4FkzGufpuqeRy8H4evMMfgpGY+44+YNPqnZ4NpPBvSIdK0OeATDUdIlSMUU
wWuMYgqK0ClIsMx65lAwdZqFjFNGmTU6FsC5HzCFjk/Ty2Jn5GJfx7Krolnm+Dkj
htGzrizp8jUjEyMtH9TvJLA1ZEIodY4phRNoCM5rkli4sFMmDvWO0+SQbA2sr0cd
HHokzha0gCX0A6LH1qTrGVUW9PHpoDTBER6dEZUwRrPdrOc9j539/TeejAOo6WRx
YOiaIeihqiNkfNsiG4RR+hLwjENSBAWFliiNwNp6APDOgF02K8yuSEq4qKFx+Zzo
VZZC8MZ74nV/a/ueXGmyKPrygfA9UP6Bk9KfZc9HOAnCsPUVNRis+miKIy8ni1dA
jB3O7vw87m0giEx1eFz5LicA+8M3Pm1koOK5Hj6tcefrJdaXav4Br6b+7koLOJiD
2pGMQYrsEw23+haDXl8naH8WCzALtqnPgvr2EuhfBUzmat5BBfIegbbttBSPaepN
LVEfrhgmGK4QfVo+Pcg18sWjfwLVoARmYAe8az55IUa+/Rls1denqqLKIpzvKkIp
ykVODcRK4hGqv020OvyJozD2RvMHEd0OB3EJRM9h9VtW+cgNfBOLyDzfUF9Fr3Wf
W6dYweZL95LUw32HzOUl5ttzDXZzB8zvxPCpm6GWLFDcBnlvuM6K50ws6UN7X87I
7BMzH2HLFB07TTiID8UBGPvHkht0EO2oOK51YvF1DPqqwYecID383OkZ0lQFrvs7
oX5lXwzUlHZZhW07sDCCqJRFVjKcZWicfMDbVGxfYIZfl8Zn3nkprDyq9T8MKGKU
GupGXTxTgNWe5vRkRVLTWxqo+vioAPDNlZ0Nx3CW+Y3Ru1aeEqgNDXeJjNaPBOc4
3uvHNQdRer0l7vpIXFaELhpURh2W1JDladqlO+kHC7csToCTB10yDN5fcEBowbbZ
By6/OTffH1vJSb0cNIpPIS8glu7gXscMxvluNAy1MxCp+aNon8lJKxBIATYmmS8I
TExTvf2MAXAmzrpsFk+T74dHCm7GjRJs8CithE+fMg/WrsaBWXnWIFf6HD1FcZiq
YIteESi6aoeVEZ7s+MsmMU19++Bh0FCH9ihafFGcJLO5U2P5ziV6e5rvbWIOy+pP
lMtWJe9shW8UlPGciC+zhFauiZ3rhHyrlHdFwvjyNzFctxteT7xch+VEaLV0GvPy
Q5X6jPMXAcxCzc02MteS1+6EWfuhJVsn/ZeRSS0EM794IUviTmLhjNqdNB4Rzqfu
MMURyoFSqaYL9JlNLaZ9aqKGSQpmIMLt0ztPbvtYUQEVc4r3vgP6ItBKwR8mTIyV
XJ2nyLbmbfoGgkSvYwQ8xM5CyFtutpk7w0yVbj7lh5uKiAECvq9LowFKiPaOxQYC
z2A2xVA8VwDh5X04b8l4Rr1eFRm21S9L1ZBxDDMEZN6VFl+yJzkYZ0T2leLcD2hV
eNUUgG7niKy+QS90GfGSGyCNOKEe6+klCeGrqyx0AdjLwKXEs6BCfVKTk9KLMMHH
qJ2BBgmR1Xu/0Q84L2ZnrYm/WItNyUup8TykyyXyAo47V0DKpMFW8606bq6O3CLk
MAECaNPclRF1TB6vZEPEmnrI4pDotWtYZCkNCaCe3mvU94/KfieFRF5LYa6w4c87
vaylMijXmUyW/lgr7g3CvvbMYs1X6UDY9MOhSlVhIhteRurFGi84JhcP67UlbuC7
WQWjM6WafUYLDeUuQ9bj6cBZIvGjMygxqjqG3vBwTPVhfze0rctVRfUjeG5Ld1m+
2nTfYQFqCbm7wR6aZAtbmT5hfj5hhlL6Tkztjv4PwSPFFDwDKgNGEfY1RgAKd92P
NSq9QNT9pHgHH8My13v9uFB2WfYkdwuQahQUole78g37fOWRtQEw5nx40u4c9Cnq
RB/Y4O2SCDv9g6Ub0lsbQyTyKBpB4zngRpreOEV5nciN7ggCFu1ioSkplsLKfBb3
EVW4nPSwunNV6k2jnI1njX0oGIk1pPJO7PWO8Jzl3DyWCwxL24I6lp5Cdt6rIEWV
QjJnWwVz3oYbfY/repHj9CMuS4A3qTIinS2QroOBWgE3VCybaGsgZdy+qo67fYNu
jQ3Bs5QrKEEmhFyqQPed0Jf4cH1KSe3Z4K/5RFVd/udYiU99VDhFz3H2ijGDkh9J
G+iV5VctXDhB3326dReCkk+2unMmmAy3y0ZIcY8qmcMwDDSI3pbYk2IHB1tOeUS2
Ts0j9omJsmJvb4t2I6vBEUtkqhSfBegwsJ2eSLj9BN3URDKcDF+9cCyhtc+tsJzB
LdG28LKgoiiIeyQ3OdtpRdysYDlCPwJRqdv/0v8cobWaaImHTI/wqt+rUmgQLCbV
uezRSTAU5vdp7quPkvDHDXA2GCUcYyX+fF8JZVYijIbDtj6t3y4DfUhip+CtZoxF
SVmZIjyAbW7+dsWKtW6nP9+uUJEx3YFeHRIUSsKJcaFrZQ1pkdDY3PQIxtMf6OKN
uhk2coGTbEpt6keVjQjBeDobKWlijsjdrqEW43DDukHohKP1ZT21PjpFiU3+uj2U
9RxUmhTd7dMq4ip3uHA+OVVX25VpbEom2SRK73BJt/4lqf0+i2vMSPsMg1lcpus4
FSe+oSzKLKx5B/7DSxLJ5bJSBxJj076mwUGsO3R0I91uHoJXhrkOPl9zjJPcvBcy
qsiZatR46YOU/3MOWl4NFSntJhzlqvqnVyRvkIwP3wSZFwpv3OUYvSxbHhbLhAKc
KwTYZ0B5sXaPNowXoQ32Bdgp0/e58VctBBJgHpNuh9hU2g/EAcLNotf0wks2q5kj
KRhDIcRjvJUStWEDfFUVSDZvVtMA3cqLLWl351S2njU9mJNfOEEEB+ZZEQj7OmtA
YTMqrVhrRBYIcuesBlLk3kjKZQzGZWfvFavjax1NqV/q/X36Ehl3fIYqbjxnnOB5
k9zcwO3EVx8q5WDZ9zQ6t8LbM7dS4P/OcJT5KzemYHUV28pKhZH8940GRHK9C5Jp
rO4lLPu8z8EyKJAHsvIs8phBMvIHSPgV+ar9h7469+9VVqf9atKMzI0balt5YZB1
dzuCR06rqdIuzprAGpjMb6cLzM+qkTgHPC5hdaJQEhxlUKjNbY5DihmnwC7Ua3fm
dijOxUBrrc6H+zq4GrnQkTskVVtRhd5mnbNcNZdGgmaug5A5yESvKjIid+5v4A+B
SNxgDrX1lDRxaY/oSX7hxcJgT7jUTmkBhkoRJhZjtybBCQfMTig/NuxrVu6pviHh
8gq1q8VsJf6PgNiahf4H4TCNmmhEr4+J6cjSI0xpcQHCs4k+r5/YSt7jD5yhUp1L
jx1gpk8NmO0ulB0O7rne4kXGNS5OBjpwSKChjUSX3iVuyFPI4EYvqqqyX1v3cpFO
0DzxlaV4YnjhlLIQwxkKzQMFzDT9g21xVTqa36NKmwHiUKIMVo6WHOezj4ItN0Zf
vwgxyEf4yCp2BOzOWoZQJgAFMWsBPlvTGImni4qcmGcEHcqkn6GbrHbqRox9LoMq
lLv4W8NVwQ0fk6XvnV9b7fGYC3k633EnlKt0CJ+QNsT7s/KHk87oVhd6C1q+FQIY
6aIxG73mvwxrZwndRf2TG7G1bMHA7hRl1oPAoRcMXpWiYu6cAzLKSpMSUTs+2Z3s
NtI+guijKvmIt4x52lTr541ldKCMNUBG3XjMtQwS6BmpV1M38iwWQEkzjTEO7bYe
Q6Q3GIEJp2zh7JuGTR8prfno/9+t2BgFui/JD1tzVQczTmoK3XrJ8Jo8V7DT5JDN
HV/vNT5XlFqQhONMadubPDrvvq6e/8HAgzupgydzaZ9lkbuWEf8kNIQ03hLSa8zC
Xp9r/OpP7AMnEbCu7nng1mFn7emg8PNI+eln6SvZ3Mbsx3bkQHNTZSFExMeyDdAQ
HSjGdjrk69IYd19U+pe9zXYBwFxkx8VPwc1ZKWs/lUgT/Hq8t5lDcWrGLU/sr+0U
TOnkNR5UUfsUKW+Kp0PIOglnadghCS8kyzI4RzKRreGqpYABpuqgHG8+3PJgSD0I
Sbmxry284mmifgMK0PdHgwDy4RuP06lyWewDBBBB5ATzXlWwqHEkT0fWioOviLlD
RffnhhLAKmXCbAFMpIjSBHumXzpI3n52h5WBtOatcfY5iDpRxI/vzQ7zDSmS7JfA
2yhyu2JCUE5bDfc262j08z+sS939vSddDEthqYcQ6ciOLnBHmEnbAhkncS8Nbxgg
OvEKRF5SOaa11WQY0vYhzx6SZdQSYTOe+RhwSYi+wHqjq1ll+1/FYrR6tju5NChx
Li/SbH50mKHtsTopcR9YsxGDdmlLQNJAWWmKnPT9lzCCD/wl5W4GWjGbzzZYsabV
+yQbCkG7yynDona/Zp1J9WkK7+3CDjGWGAQ5x/28in7l3urpSlIWP/7tINpHpq6l
oaF2lXRP7IAS07TsBA0E0S04fO54zx4h1Gb4IMD2xjD90WDp1XBZxVb8iT1kOBrN
AFcbucYcggzpY6msjFKCjlqoxHISJZeqXT6aKJvg9zfKHwUaTO7iJ0HdtzHdvfFN
858k7/ptttXKBgsxNJzfakgUeDd2Ss0WmkTByxZDiDPPqMMdEIohb+aE8cDttpX8
i+g5k2/BphfararuduFR5BxymeTIVetszeR6WaFM/RSmPH7bW39UNnZ2JK5f0VRb
dDoK+TElEeCAiu1nYXhavcp0MbsHjhlzMEe6YmqES3yvfDbsATks7+cyBwjyD8vN
yeT9KEz0gRh6izdcITYYpYEy1HUgFxmtScpp83u6WT741tHTQ117QwcMhijY+jYZ
9/OMjHfP4PkAIIii/yDWl8JmGqd6vwBKo+5Rhi80kaX2kgkyPitI88/KXA/NDRHS
6NGf3aQZ+Nlm41sg/5XAP64w8GODpfFkvw2ZyKshPdKVCudZdDkuLsVDo4A4PR3b
6pqSArhY6ut5B8NUhjbQVszAg4rN5gil1iRbAKURPa7y0DP31lsRu7QrarNR7v3E
N79dF+v+PIrtR8M7UOfP0/rYpaB2jj/GfaHDmadVxKiC11eV5hz1wwA2tKLmvt9J
b16C/wBs1QF8wIDutN7hv1IE7NoP46mfElwKuyOl+VDwp9C93rPdqzt2HIzrB5D0
kswQ45p2iWSkFpeGSgfvSwTkMOmykCSr0PqxjDF/WajRcoeWuIXaLb3IKEF+t/uT
S3xE7MYCnpaocfvjlZTMqbGT79mq4tvRMOGIGBlBR1u2UNcbIs2a8aaTZVIBbJNf
y8bTNLRvc3hX5VKCfcU6INT7bX7RR+gayKn8gvRLJ6ZPBM90q82Z9D9//24V0be3
LE6/PeSNi1LnQxUbuksDO6z9Q2IMub7UCt7XQXOraVwYdaUZjGGSIqAPAaVQb5dp
tQwdl6cbHpT6ysBAEmyT4Sy+tCGLaG8sv//XsHOWVTIBJvXSALY7QnG7N93Wy+Ui
bhbJ0btjNiDT2qT3MsVCCwgeVGkCCJVskPSQNkHbHNnJDdr/GPLIWCjUw5isiOOQ
xUzIVg6XSI+Uo5wQreSGZk09afxYqySvh0bbjQ/8Ojl8QmOVIFIMyoOxSHa68zaa
l6wC1pbrKNEBmWv8mTGZat6FKVb5bCNYffQ1kClfcOGOBGRAiSOUX7aQj2GLjhfG
RpY4NoEuxyrOsW+A746WgymfWcuF93iZvBK9ICOR6ATxwyQxD5PMtxndkOm+MVyR
l4fn5nQCB+k1q9ST6X0TW3cwh+BZ12l3iUgWQ5ODj9/FIOddMwl0zu7o+7MadM2O
aB+2MkUTZZ98dkSZJpjewFZxQ2Vk9rQage5MMxRgUgPbGzKXDnkAzSBFFtCdbF+U
azpNCfyoUXGCLm4/M32wokID/3eyJSlKZXSzN8DsSUAQFw6Dsr8PX9BcExtZmQNT
rhRMD/skAtwckmlnr99riqQN16SkAVd9Jc3U8ysNXK4WlwSmMy7chcJWY/jfelAb
FhymFatMRCGTFmcQgQfp1xeB7crR9bCY+jFGQTX9XLxSC/8WoVjmGeSaQc9pMxYm
gj9SuvBdTOH4cykJOph5fh9z5Fzh7xkVgfiOycv04wWuWGl4VSFprOEThsDmzT8P
4joIVmSqSchBT5kfkmqTCQJi5vSUjiNzOevjy04MkHAv2njcWrf46EeMs46TErOg
/NHfD4civK3RxLBFraNHiDS+pIUIliReDrfu6oVHnzfU4SjDLyhgypjl8L7F3VTZ
HPRJIuUY3jpOb7nhAW8wXCjWTLfeEK4G6I8uT4Vzk/uScQhkw/XAI+9/EhIt4GPY
PpHX5Gp+zjQb1xbMBY1U16KT29BLpkueExXwFBuN6fjawW88mBbr8gF6GrL+BoLD
PeYoTYzzr/7cI88VaVUCijGdhk0eaKFWkn/OWXgmIFF71XDarIlpQBnrWuf+RKg/
HvDATOOqMdHMXmOqNc8OPB88BZVlrgzGVEzwAwHB1XJg4VdTm7OzcU/ui1CSoayr
DueZesgYkPMHplTEklWAhI4S8+D8vEMlsM8+TM1LI+q/ATLvn+Kkzdt4UtxpTTVo
T6VtjB+/gN+EivGgU6RsBZkjFr10TmmiU74JtMPbYr1bfiESw5FaQ36Qr/o8tMHL
ygdnIWZvGq1itUM+jYsvkbsmfF5xvCHUFIB62y80YPtzULBmXi6Ucfyi4nbJ+gab
cbuUdF6lHZP9l1xVyGcEEycwPWM2ACtUWpdYJvQ/mV8NZiEli7f518TwrNc5V7E3
7kGinOGzt3p6pv9Vf+nbf96TVuxZjXl38dWuISupNG9gYhgnRoBXXRBqkIPEY6pH
SrRaryQ6wefhB+wS8orqjMUM8oiAh82EJFErbPqAH6JRpqu20zhpAjnRAFvBrH6f
ujgfMs4z7eXKBxscdJ/xM4XxmaiFRCi5pbRwudAMwU6GYTssTloV1yz/jGdrdpd4
yNN7wXReG7CJ7wql57KqGmjFqeMnu+jIoTms2XnhsImfDQVz2uIoVTCXfB+kgVG4
1HeVjEFN4TfZBTEFlSTe0/T48mVaYHmSPPf7cB55NWtL3VIe+QTHsl7rXFGC3zlz
5pwNR+WyG3VGXitl89NWta6Xt+MlBl2EhNGhnSuxrjMRgN65PmV+WERpF4eiW3Dq
x6UL3RNbhEZRkY1BIBdrfc8YyR80uO1NgP9QsEzF0UBoZz4JFocroJXf6T8Fnqto
yiPRPpQr+eXVZNx6SAlGzqQGZ6ffP9ULojzs1ssjIavXi4DqWfFozUQ0QnU80oxa
P9oL+kN/dpWujODzdYYn7HTEkXOVvSYDyFRNl8BfH/uclLAnIXkeqyiSxaeRsaGh
ltLubRVCNcRuU7r+FG6t3LgLbjrcTnkPAiZei+AqU7uXyiBtLFiyz1vptdYU7twL
ObCbHRRBWZsoEoUL71uDKN/zrwECF5KvCoAyLFqsW0nExOUUpxz0YWHx0VmKTPrv
jeHENRgwxMDs0O/kcKLy6nx6lEinPmN87GignY5HVZ0s4//zKmWMIKxtA08Bj+ak
XgZAJVdtv8SMK/LRG5U5ojZloWcr0FP4G+Hg7/s2jp2EadO2Wo1PLm1w4jSvJfYO
HMLlrxZrXSm+APM+yqibAZGmXz0RQMUQqfffBxthBQjbMSJ6UX/UPZTfXHRylH2P
AJ+xpUl/WAbIe5PI26yI/MmSoK8kAN5efDU1TWsgGXpAk21zazLKDid0Ki1blvRJ
1jRc72ChZZyH1ux1V4s6ysTXnHawNgqYFx9NsZNZhcp6ZliUMLzlqmjhDRBz1L1G
zuln9elU+UaxAjW2NxfuEdi7fs/8OYOb8QSQSb6tGKaxhWi3221X5geWU5IVH610
maBN7TNCRy1qqYdElW8Ar3l6EEzI2NroCeLdn+bWgh1srRyyir0GQhfcOcGuwQ4J
OaumEouc8qC9Hs7onMYmAGrUEQwBCJSftxG1AyRse6s1AcolqrzO1MCt69/0lxzl
YU/ZvGusFP6eN0KWWNDxxT8RxEqP3M0vYw98hLwrroQSPuFgLCvmSi4R0aqcXBTF
RfGbFNew+i5Fmj/QA6kajAKVNS4FDU6F56swOIjDp/5mLXkofPRei/zYrTicNOR2
gqKBVf/3zuozNYzUJksUp1CKj8oHQ/Ae5I2UBU9YdE/2d2lEL3axSwYWWVpGQr0B
ADWM0vdtItlhL9OXu5nQ6/e8Rbj+57OdkGIQiTZnUbFNqZi6NEyi28Dujb4XARsX
GykhbjCNhUqLb3UnYL8n28K0U49HX+TzkAXsYKu8ecDVYZVJag/v/QdTkfH3y67a
UHu3HUkU18+gJ7MvEB1v47Ri+QlfHF3pyHZ6SlJizIAJYJuBgRqv7Uh3nEvKvrLZ
iNMIsk0njMUlHMxI8GB6cQVsgrqADBXnafnWbI2FdtdgIoiNGyQ2QQf/nA1PD+dI
ruSbB1gipgOtEzO7UhuFSni2tcvHsEhlrrB+3gutPx7Zl1W3lPE454vhJ/lNfciN
+oXRlS0IgF7inkTG/fQlLWtWKRpbjueRYCl2fr9PhHzUzZmgUePsXMGsNbXcZvoW
2GRgGTQrn5au6z99SyMoMomGqjhrHcvAgXUZ+TZu8vwUhlB6BwlUyqpxbQzEAS98
/IYGqm5OIq1fXmHIo+DEGrGS0JOj6SfmDTV2KhGzfGTkSMu+55yyYEbiVVVntqkr
tOYlAOD5Wl5AWxxYowPx9nZT2zXoAP+AG80qKqiXmfklD0oV1+SpHy5EkYSaRc5L
L/BJXKyvxxHLlkQ8344Ac3LO5Ji6DjY8t3nq1zIMBGyBTjeFHzJV/kcSxnQnGaM5
g+lzdHJlEmdE6wPhgM54XCnwV7mcBA1pHAx10gOoD/my3I/IySQoHw2jE5I+G/er
EV7QO6sejd8+/522U6ZJu89BRQ9g0hQamI5AjkTC8xdXu5zOPFRwlxkIvbrbgt5I
RqA56Nhvwc1q2elnrELr4pAtz6QiyEwPvIKhR1Pn6c2P+7EzNsVQ8szeAzWICen0
8PaSQJX7Y23TkJIorcKGil1O4qrtRNXUx5TthWVrJ+v1xoSDyGXf9e0TYXa5Kv0n
/yii1najRq2S1Zj1LNh0Gb+yQSzgyVjJ+m/qYiAjUhSDOEqnuTlgmGFH1wIYxX3S
y4nyHJGKsj/bQO3hCj1M63w8w6ecLXCKEK2grsY37ddSnJFpRb85V6UJcHrb7NyC
8J0my95JSYQhpcqXhnHE+YlIoHjOGOY3YsEHcOun8dWsd9jSup1nulY2jJT2Ljsq
6l7YzptQZ/XSc1hskHBCNA/MYsbMIyeiwM41+6heKcuOx7I9nu2jsLQh+Gjl9FiN
2BbKK+15piu/5XDJ5uJFpwWCoaBKrO4theJNXyFfXNss1KIrKYWpPQQURT/GxOBb
0g0pzdIOvVZYZZDnZxuB0Ad4tKz3p4NlJ/aNlk2Wcm/ot93t83l8wxbEGzNi+j5n
GcItdLwtviDm0Evp4gj3fUhUW1GnkeS49MtvsZtNcHCewEZaU+7COoLfCGqr5EJB
xdrbGt98S1dYNctwQo/0Ei54BGeTE4ReWgKe4nMGsS2WJsykQ2dWpXpPkb5cRNIv
DaDSgMkX8tHs7HwlH5jY82c+OsaMVvnb4ZfSrvVUjQUmit++eg09YfR9Qhv9CRn7
uWp5qKxMY1MpshZ3I9/FTVEVi2uBdh9FU+RCRTp0gxLbLu8fSuRVSHpz/niR03uc
gLqzBQVSXkWeHsBOfhncLkbg5SNIcG8lSQrXXAsgI/Ft7IV7nae2qbui/tOuokWn
SnaeeT1TgrdKZdo4g8YladzWfgom+N1dlPagdzT/fIbzYswrDhO6jtSA2QeNwO2M
P/uJmenAJJSlVPxJ3OSWklFEUCasWKJCnoNzBGoiQNxvVRADD+DdFaxPGxBeJPdY
IaUICBndxsGuCszsUF9ML1rOftX35AMBisQ4UpvKmwLfw19HzftvSmcdZXFgAaUI
pyHLt8u2gRcVI+SSzCeMKWFzzNF2SLhd0cECNwOIX9vfkyqvoTYKrfVy3FaeIBVX
H4ojgKmTWFoH7RT7JfFbmDCdnALhpE1nhFKdRKTEs+gmgOzrSO6m8ixevO9THctW
aufpqV3gMFEJSYeWWhcqD3AdYWpenFtuCurGmYClrps3EXU1Jkc8BvJYMAa3a5nw
ONAdwMzVAi5Z00dwcGb0BTht8MR6v3r7LUssaQUYRKqwx1WG/s/tee18mXpq5zSt
O94BKDwkXBSZQN4s7B56JLHe7Ppd2jZrpAlB77i0Ar2HOLiSFwUtPmaxOdLu1azK
2r3BO23pmahkVjpwfXgti8EhGhLjIHvbDffB7Jsg4d6NfZwBbl+5yDPMnxnu1Ewu
nbg8GxCy0wKLGiAqGTKK5+nssEv7vbtIhF7IxDI7SwSI1FzACDt+0Cx1Go+rcdWI
NViitDOLOEpQ3YM4jAXWZjLzdQWoJx04bgHUPuBA6FrpRuCQHoqjSaoPDeuXg5M9
aoYbIUIv6is3Go1JdlvyxC3lDgOeizOp2M+C2G7cF/0Mp7CI10so0N85O2at+RgY
FxGqkL4cIBYGNuPL+wI+Co4PlPtCOdoe4hWQXheC2ml5A9mvDPlVWLPOi3zwbYC8
0moXlHn4nAhUJt1x8EkTr5tWpZCckfrAGSNX1bomA9Hb7GSH5XlrYFEMnnea82zH
Lkj545BOX8NaS/gqDejvGgIzjpvd0nzEu2OY9ENaSeNWdiXoyHc6XbAgixXIMH6M
e6DlBE8Tesgl5olJLkDzFFN64NYWyZ3bAOOIeKLzeu0iplF5hPPNpz3Dr8TCVU8f
kGrSxLVdRcmAMOS7u1JSV1co6UI7lSIEEikIF0yLA5dLhFMS7A66Rd5PNHkNd8DZ
/bKld6ZXx1SJwGD2K5tmLYTmJUQpW0yd/QxGZmOzIjzfogrIxscP/TujZZ4SuEnm
7wY6cWKkNLS8Z3C+3gIEJEiIiboQXUf0lwRZcAHx+DGItgCEx92pzI8kgkDpm05z
B4Wu8GMJlQav30p6tSRKg6mNOR5cdzZ+cXEXGPRX0vcELC4xkz6dxIybcCMWvG2Y
qizJvCLZdiEMjw7sj2sPghl2TNCKHVCv+FnJxdO2h/+AU/JEsc1VEniZL1yKbDzA
XtJfuzx4rzII19fUfSMHnMe+MQi9ImePQ6GoiCkLOvWuA9ew320pkO+1t7WFzQnD
jgfVCpOrzw5nAVP43E5O3nPYqfM7Io4PsyyX2RSXfXsugHEk9v/C8hduNHztaMTq
NGBGOWK07RrGmcOlT2j7507y476oNPSAuEDKlSn0LiagCUOeKxQwjZPZ5QuooQpO
JC5phirjz2wYNAQuGE+/mAAIQmKCrQi5LDKZfFpY/iCyWyldIEpLTvT65Cz1pg05
wZ+MbhrsMThqkb4PVv36I+TTC8X1ZE2/c3O3g+tDYd3PdEBTCPgppwOPFt2PxeRt
BGR5LsKtR6MBiRkAaUQ4JxxIbxcAQ4IhdQjfN/BFQO92YOUOcAVC7Z3hxpsf3KYl
wE0Z8X3anWqHb9jijGoC+x30Twnv2jWgzr8RZr1CfdIIBSrqKXqarZLMoAAdwhfD
A4dlxJwxKFFtv9k55ZXRBreiDsi9ed8FjQbye1blh6sd2Jvq3RLDK1ecN0iCxg2I
uyrPqx45fSmDZ+/rDhx24iHkrGBlrq53c26uzl7pv+A5q8Qw1QoYb6QotsZJq0Vw
j6KhdVpG6gGheAxTXD6q1huTq8wdF4Nt91bIQGRVKUFhrDFVkP2iZ9ASnCFILZPf
eicQE0voLfnJIZNi7oWUhYOEDPu5X/QMAQYafLOB6PZNyLYHLMb397Xetpmhqu+a
5noCO4wZVjsf7MEfk39FsXGZTy40/s+S6C3tlAylRA4JIq1uF/2TBYUGEBxGcxyr
VTbzJRT2m1aofFNxORDDp/c9AWCodtLBcwg+cagp3snU5FvY/HGSrOkYAY5Z5EU+
KssJLA/QTrrI1KJ6MszwE1CuBwrbgGOlFdnR43/L6JCaL8mfAdboOg1DIn3c5obG
SnK3QOrZ3q2sb0Tss1yzW7VNjHHq86j/boSsR5ANl12m3whpbwG0NZUB8UWiTj+Y
C6TqcQ947Jwz+BfKGc+ThP7Jd5/PkQkuvxvyo007jr3DBlfnkTpklZACpQIiKS61
Cd6UFP4v+fy06LxPwaZaa/qA8dYuu72blOLix5TgQJfrEz6jV1BNaf/Kv4y3rFYQ
oNQAsW1XE/fPsWOUpbHKNd1zGLpo1Q933qDhwbuQmkmUni7B9AR6sL81L7IbeAsB
lpg3kQKj4C3J+2hmFUds9pM9Um+AaYu1ziRDd3NF7/Vp4Z9jh9m9/qcvz1aTkk2B
P71cr31/2cMD1SbFVWMPN1itOCQz1XyGa1xM6aGtmOIRadZFsLBetpjGvyzfMtGs
Bc3zeCSIzCuigFFmELQIFFqmeZkV97/+Ho/DMCmgNd8z7GW9KggmKK5gPtn6sCJV
Y0IZMyIzc7ONtIcS5ub20FjdxpY/o1tNawOdUZ+pEOm9uPoZEHcd+ZV/zsf3oJDz
DDzrnx799lXaF7MlwZMqo+WDHxD1RVFp2iBf2lQ02PuilHbnzxFvViXNQp63T0MG
w1zd5qQx0NSjYa1hV9cK1HJHcJwWIueaeCX9GH3lmvp8CEBUJjsQimcuCpIp4kP6
L2suDVA2/ppkPuv3c1PI3ss9HMK79vaVA1Kljg+higzspI3zB9gsQ+VoPv/plrk9
/AZejPhty2g9qzpVjypDFMWjTnRmBQrv8lfN07sMy70G48It2N/tVChTdJX/L804
xNjvbV5FmvTuV6RSoaOutVBZZi6PbkzLeLTSDdxFR/ZEkABGRE62REUwoHlRONlY
74FBCfnJAVN7dLSd/V+ariQyugm9hsrQ1/aijzotBKj9lWYPr3PRXdNLAA0aKb9l
BQ8E2tqqgybS53E4A4MZTXU17SC8UEpujdlpoUPdw3W/3zA6q/d4C0wjmSwK3Rhm
gANZNkVn1zPbyj8yQoKCEzPtC8ZKNyF2GvGCKWkfJI0qB6oLcNXybgc1e2BGGM2G
Yr+DZWrYmvkRW1u5H/KKQ/GF8J0YGMUeSB9/+itLEumP0IbIh3NlAYsXMRpLlmmN
DR75Enbpt7tvps7gahD3NirEIOcnBGNG+mLrXWFScR30G7n6DBVIPBfcUl9Uon8X
rH1H+iBvzhCu193BVmysx29Y4+TObALQdT94umvFu3KzJwnAUwtzt9lTc59eUOZj
9heGMNSDkgXK9dGhIDKKsuC7mKTBVN0HfvsW7aVsTMX8BSIcMSdma3ltQ9/MZbrP
VWclAnrXNwCMSeJNl339KOxRbUn97jHR0lMBVUrCtIHnpAUWt9SxqnMzXRtf2pRt
zyjdhX56+6CGib/taDGEAzmpk+DIotawXjcCUzJzLeTC6SRopVrIxQhPLbfW6H76
Apy9S9Au97KGShfCWDx+fKPXfenMsZVZAa0LMKzszrmbJ9N1P9VjeeY4MHX3LVlU
CAjuSIjwdVausFaS15UjXEzFZ151zB+9Anv1230ogRzB1motYKx/wSI6vZhdBPCH
GJMlbx5CtBwAaVAv2xA4P+U+JlspdWVQ2JPD+kwYMasglQsOeNwYDA1BmFdwVDmY
+pPXRruYLYOHtIAsgRBGsg4ITUzThZN3dfAOUnRR4/O7LYUpynFa03+4hULSMPnP
MWR9a2WO/m54Gg66wjWHWYIecy/eDs77u0OtjiTkz9LZq040smUP4OI9KbcPPAk0
dsP4NrUAVwW0qhhqKobXU6MFm1IF9Fl6B2bKVI8gpTZ5Towy1rYup+ijkHy6jspK
0J4QitJTJmaCpGxgeNLyKkul0cLwYPydLhk8gsy61e3nYcjQnsjxdnLQ2c+G0KDd
/o0BwJTAFV8FbmT1ivPY5H9WdeYEpLC9n4Wo1+6rZ8TIezs5zE7YjdgxWbXR0Ttv
kuB5Fsy1u49qmdsjGjifbzuWpgyg+m0xwhP7rez7mNpwGsd0b7OgdYVkOXyMyrMG
9XOt3TTIK6yoyPFM+MW9myK+qU3pR3VwSAaqmVuNmGSfal0oGYbXN07UftFGoPT+
a+2WkYKuz7yQtalJEL3nbypDVsH/O6QR8i7W+Bk+jkfOpU/f/DNGN17sMo/QJF6A
ncCvvsKFBRQ+0ttFWN51+dYSx+ReSuCqA4F9+Y41rr3gWE+ImIa56aIV9qAdhXRf
1YaXOMIHABdNRO+VlAwLM+qJrtQq/VCyWThsIzzvPThuW4wP6X+HnVnksLtJh+RC
Q9KLnhYmaymU6DtVJkCpeazG8c5m/iQkAdbmQ+Bli4LpQY4K6xvJEqoblPVhC4CM
/WqoudK+MRCi3+LPgEpGYq2jJrIwwpI+gE5p5tAqOVLGlm8fE30nGWnQC9xwWKfm
HPjpYg/yzrzUBCfiONEjs/RS3Lk0I/u5OHZ0dmdZinmW1VBBLCoL5LagxtERvcvQ
wf730kHIjDyj20tBxTHEjY34su5fsg4AcDVpqN+xTWaAZu73hinv7CExb2C5PIdh
6VJhf/+SMnw30hC3ORL6gJrFNNiiDlgKcux/Uj6qQc6G8Y/2MUmOgTbq5Fv7NtxO
ppBTzUy1Tf+u4flCiSIf6xHQbJKd97/suZOx/fjNFl5dNHV06Brql7+eU35j47D/
0LP4oE+PNYdBsMGv55/+xJypCQPhT08xwXTOEeaKFSAtYWI/Jg58Pm1UwsZPqXFG
BUx4r0GcWwxlebduVnZ7nmnie/XNisete5QHRsE13NESD21o8BD4f3qjIjxkG04A
G2ojgcY0tC1ACxwRPCniQfjex9PCWLy0ixWJmN23xVQlGt8wdnP8sn6QxkikCSoL
wKl6GIgCMTjrNg1JA8kk+qqBBig/ntDOC9JtgA+KPhkcBB0bdTTNP1pxjm98bii9
Jqs6ginjrA6t2LEpWZZWesRx8/m7V7C4xhvr8dpHRrBa3uZCT/taWHaoU5j+aIQT
ZJnjR6eCFVvHzlWriCQmMoMk0UoEOkf3qGTApvCZjd5WTFfD/eCl8N/rrwCzfKO3
v8x5+vW18/rvZOel7WEj+CTyNDK5fAO8mSz5os83nlth6/vMgF0v2B+6zyDaReB7
S56Jc6DhARJkQc9yyjOg3N9SnMF0X52yVPNj5RJrBr9rdh+VHMCnl2jIQi8gFCo8
ii3FN41eT85Ql4qt3o7uiCLxMlgLqrLocQepMzmklCp9X7BMTRIItBX2FgMrIoUe
ynR8pBso9bYG6XnOppDHK9yvK4bh+DNM78mMFRQhelwhVkhVmWPxSf5EMO24ERQE
oMMAMobOxwZ+kz3AFQgJ8pvqFdoPyT/+EL7EFpN4fqJu/GT4T1JiMNX1/iIMJV/4
fo9qgJIuBWttWN+ahJeDOqLcL3Www5H4bcQnF80auB6LsLBA7/yJ++DWnwaA4nVR
d2mlccnQKwwCrJX47GFcIcqx5ijcBAbA5EoajQLoi9utzSfV+89m+stueNAC3i0m
3DRQC/RaIgjn016i9pSs8lofQHNRlf6AulY04v6rWhV63NCaFjex8YIJqq1Vffs+
ivwDPl8MjBZodY3Y19JJtR6VZyR5WOOEoNGqrKuE26SsIb9eI2ZHhGIhw0ElsSds
gW4u/zfYe5XrxMPYGnMRX6mUncoVcbYCLKRyXMn8vj3jngcHyhDATwxboED8ZC0G
z5+t8ZauypxOiayLHUB9qGFnBP+FmAx/tM4I51ShQUImsdK7MBVlT5QWLaPIGhMF
OT/kyeefNSP/KFbukSjTGbwfJqiN9ZwyqvOqwdGUXFCAZEHwmxQsOzSfXdutbvgI
s9jjcOdDcxb2pvnWdMmNUBcorwDJYs7nHrlFT7AZWPbn3tDFKjImm/ZERipXFKQ9
ylaIlFO3bqcGI2Gj/z65poxJ38dTJMqZnz6W0gYWmEkH22Cs//a6Z4NJjlUC3xp4
Eq2L9FN8wbEHCDZwmbBqViRRts6RhtdDlDLCZ2XdI/HEv9VVsqeKXszHK+vR5iPu
iJpo8bfZ4RpZcLdxwubDbAfyuu1Kd1ckVEEgP6w1pu3eG6emWeAjyMedycWTDOj0
So3vj0+FexON9pDQsByyY9mKgyTToq4Ta2w8Zvxt1k7H1s12gFWG+zdPNmK45Axw
SDgjdh/ArNFhm4srJAvirqoZjeT8/2qJPF7lJ8dxB0khfcVB5fn0tAp6Nu6kK09/
lAQWzt2jclJtsGsPsy3JNR6xsckGkUKNcARFDqh5qUjJgKdnOdROeSt/3/OwSSHE
GznJ3SeTouhAzODC7kCdKRaZzAIxbFppGzLjfwoQ4nZLUe9ov5dbqjp6Ms3DVWCU
ZBZ8ysbXUXw5F2LXoOZrOda34NUEGHadyhAaGH9qYj2VYtSf8S5VPUhH8s8n5Y6k
zyunrDGiSzcQtIRSb33rMx38/NFmMtbBNB06QXuZAPKKj7jqjr9myd9+yACE+/JH
G+QrQm05xbsGO+0kKxEBuZMQibrqxMm+wCxdRg0F4lIP7MBKX48grB2aBQtNmxGY
cz3FCTrInDKOrSiklWqG9rGaqtRh+MnED4NzLy4i//nzlORDPKR/0FVfTMzfgwtK
0JA6CwaRiwAfD8ZLfLZEQ1ENMhrDSqPYJlV/MXevN/i8Bz2aNAvWrnYTbYZtFCkO
ZZWd0FWFncSkhUhSc/Iu3Kr0ZUI6p2yTTMHh+s100NN6ZFBTvRGCcfEhDsMzLU+A
G9dIgJVAM1T/vnApXC3mgomEfe5fNrHxWiDbrI0VR4jmZgdfBxdtmWd0ZM57A8U9
iabdO/svoJQhL8VF+Wd/Z5nSVC2WEAmbOu6JPE+GKILiwhP1vcF+OZQaunjes+8i
3iaB/tXXm1tCNGe+/xN5cqnq8HpBdneQ8HXgsYnlwkcU4oAAnqNSeBV/G4AkDr6D
rJQ1va2rfhsKbXYeydvWR1Nc75FDo9KRkgtdCjNUwlGUiQaq/CWVhcdIZ3UV5e77
4a5+pxzoW8SwSHePlPJeWmBMTcXhWzWOXvLKuLoGbWa50PQJPHHtGwWdBuXg9gBI
7xyNiqN4Cei0WVIrcgCXSXw0trhvztQAbUTTCzAIUaKlshLxXRem8qUlSVlfxNwp
s7XUIyP0ZJMzc5+L9sdqYoWYZ9OkiPK7Kh0KGLBrXvkH9utogfmryF1cK1ebRqTQ
8k5nCOvOf0nBIGZMgwXXVqpgUqxSIImD1UHsfKIDwBKzHGoYSJZ+vIkO58brGNJV
ZlAnLEqA4W4OUYW7xYKH1e29TVMRZlNJuzypu2F144seNcJs+qq8wHwcnyi59beM
B6AVKIdnkFJve0Nqb8OTRSdxk1+B71Q/xQMmeXkMavZHpxvsp/bWVw68qs/m0UZa
4463pGaBZLsc/bCtm78NJT+d5jN6yrnf2zPE5WwPjQkBxN8kdZNcAL6nXQgTMVVB
EXHOTyhsYPE19+FdblNMGVRiIUPhmFEA9H5S411rAwB3Bs4OQue6WE64RicfpQ7C
JEDNvxGkIVU5YDf2OnEHY8MiQtJwQTRVaHSDSJ21swCIUc30J5DSpDAOP6+wIRMj
xFYk+LqoIR+5zpEfP9Kl+MtTvlSuR2VucEPSFnOnm830di2HYtC4wjhrf+soJSDT
/6Saz3ZRcjoPSmtGFfUi50U1+BbEJuZm3ZF+dOTaUWsF2bCz1v0lhIIq0fQ1yoNL
Gr41qSsLf3BXW1DFIVuSYeoPTRGm5Zrs8TTGvf02F6aA6rErrJu01i4KH8ukJHAA
cURr2r10HV1XmFlFXtWA6tONr3MaG73x6VvmV+bQFJPXyMTgftp4C7yh4FTCV+DY
wYajcoBeJqv23tZGi06tWe9vXgtZl/z4kDf1eX+nnrOQ3CcbDVfs7vDhPIq6Fby5
9wcjXANsSJ3OqkoCZd4r3idwfMzZPZu7oFvSavYsV4uoINejay13NM6spCXm4GDb
GDrHb+tHtiaLVGCe7J8KVAc1XiHW14r2/XyJwsCJ24i/Vze7vO8cQ58j8Yn/De5A
GUw+PpBgNKGrggNh9XFPgu+2SPom6egTouGGA7fCNZtF8ecIJWd0k9dJ3qo6VZSV
utBM895Y5rgOrj/67oiAOJKiJDFB4cf80M3ykvakPC34s6fK/93wSBqlg6V+XtPT
XmYFSvvn0C1BZVqKWKNW5dfK87LbfyiXS58BuTsTaq5amfTrbpID6/3cNSuE4OPB
weSh3GCKtSSyjsZDKsNX+BrVdkpGX9kwLyOB167ETlf3+vqk1yQmLk7Pgu4XNEFf
BoikAbaNaHylO/Uu4eLKzxOsXXIOipOUap24924eEMEnGtd9wp/kdNDtaTxSGf5X
xowKwk7oAR+Akeryw8eHbtVHb2Az2gVZSdYHJDhr08R0+f+MuYZ/ZH3b2H22yb9x
yIDEX8YZUuykzP6tDhuM9Ebw/NN/csnmt84j4TYWFUZF9iaSPB7GgGVI/zUg4FbI
EBPFcv7hsLzTShewOP4G75B8U/uRNAoLhzYRB95P8HWhKYvA8B12USDJsCyj2V6Y
/UHFx49XUkmYzf1clQGcXdQaLJUkU9vrvjj2xWt3SrnM39IMb0hGyU/NJ0ogyDP0
a+ywq9wchQDxqeojAu3n+M7CB2g7bWdtg8WttQmyA3FvUPOGBeQpxCuSPUL5M6a1
r0050cR0a/Ji1J3OEDO5vxYV2H71yII0hLTroYdGFZfIqeHbiIKu6hjIgVTJUzJ6
nBxBtdqspaXDjQPjrBacNomBDtLnyOgisiWSmGR54tqP5H+B8dYnI+G1VJ1dYs6T
7WS23PYFYxdslmz35PHfn75/TSazZn2eT8xJ3S7DO8LWf+uzrD56g/Z41WcXqiUr
LP97OWZV8lfvxVvqfEhCJYBVclDlVhNC058UrVQp5PryVuWA0ziBtasQ/Yu6LN+j
JITQXomirzlxJhijkAHQZFyN44snFe1cTzEBKukg6CJlzWdVj4ZwAnxteEmvZ44e
+DiMLLHDEfBEnWNANCl7wBbToHEoFNqTr86bqpTyo+zI3fVQUJAAAa1m8xmwTjy/
SFV5do8ocF7/BgJFE72ecqE54t30lqdGjfvvThw7ngwx+85Q4cr8aQFZjfrp5RRQ
I1RZYWJDlHHElC2pfXk+6neR3QT7eKdcHqB0vFEox4KzLkja9R8LTCzWf+Q7iKMv
JHUcmt/qGGyuXBccNCvhOoQv1uHtITH6ouCGst40PrQVTMnZq9zjyh4KDdNhqg1A
qYoZOHfXi75xwH2WqrpeIZKegmqOZ+UneVYqwUXeMNVatgir9+vlozgZG64aXXX8
IZyC7xRildNsOBQ+MW7o9j77YZnVA3Qd1Q1Rz6yRjoxVX133AtxTPez3r0Aob98D
whIJBZ8QUKPlkHTqkqh6NBXZkxW7auRCE0UiIBgAnn5bNwKstFteoDNOEuw7O+Rn
y67/YdRYFhSNUuy0UCj315D0nf/nqylfuiXGSSOUqZkzAktftrbhcfHiORF0Rq3I
B0iXmos5tCLYBBV25shErybmuHnx+jPedEXjgtBgt8jqJP0SBG224lAwTPezhBQ5
srXonN6gycECAte9AWf+P2nSj8kxegaG4QjUPL8YNbut9NEnbfc9MenaVmU7mAfo
BXai40TeRH3EhM5zTCeQIznWkvQBiG9LVLu3OKm0FN/j9wt/I5ZBWKEw9uGLqcmM
WHt5FqBHt8V0+GYgUK/cPoaKMPgN32pZNwB3sipD2uWCaCJwm862AfXVvlARJedW
ctZPXh/OFPfGh9QaxnfJKGhdTcQHGrv4cb2ze9MTn16tbOSaJMi6FFtQDgtUHOo2
sg9eCtfNnRFhAUhOtxYnBmz2UYgDAYDxLvbGhfhg2IEcBNv4so2hsynsAMwwd36v
aVOcHflNdW9ax8kJg7Pp3uyiEH/TzpayaDARBjmJ3sDh8mJdpDqULucHDmzCh0Sl
XzC/umZeFN6EjqNjHrBjYnsc5iSTplSxKgsCb9sAu5o/eEOOC6Oc60zkSFbv63Zp
M+uyuKlFoVMqEFUWPC0/hcDREI8xEk27hqt7dnOPYH5b19y7j6hZSMpMNTAjBzMf
LbmbbfBHCe3AwoWqcdWb2VaqaR5g5arRcb1o4JOrA5PKZ2GMcxAVENAIFVEIamvx
AVE2FrGJI3/BqysWy1YtAw5fhV2VvrGze1F29heZYW2r5gqT/PD8YWWfPtkyPwmS
QUl1x8o4zX+DbiBhje3yIF6+xlNQPUL5sh8YxhnC8JmluvEEvuM2UoJqr/1QWFB7
Q/T+L+qVzp5MtR8DWVCJ/gIQGpF470p+XZ1rNbuV6+tF1b7hXMGrZxNI0xHGkK7e
BbfjfZmY4Xf2c6pdq1/uhYAn0FcmFObHWcp38x/Nser02MxdVrDyp/V42Mz5T2vm
7BCVGN1twe++kfCSfYt0I7ZO4PApgvdSxKe3XS46G9xbK0TaPlRMLH9kI/KEqXd8
E6AYHkxGZALke4vIOZZA0i+6u0FUV9nTDUahGq3pFhkvzgPUxb78xoMbVXu+1tCV
gmU8WoCiWhoWkSAJztCQ7g7bhi4mvDsqXyK32wrbnNJK0AEvYJhR5M2He1RHzLty
LeyxUjVTS+QQw7nDwfFiG1PdIioBwtC1BlHDeT2738a//5SM0UX36GBcwLYcnpzh
0dEbQs25N3SzQUeN2KGLvdwjG764/Lb95OoGQAygJ19mVqui8FR1fxCd1qD2K7c0
9NPGNMG2AhI/8+FrpbSsveiFZwtn70NuxJs8MBjlg5wTb3a8NlqeK7nIn6cZorvc
9An9UA3tfMQiH0IDgUiuhb2j3NhU5RF+mAN33/sYBvTBfgAfWLa5bY0TuKMC/N4U
Cfsps+AyWgZvujU8yXgJU9fth1uQH4bBLg3+HsLJMsuU3YCAYu0vrMFTFADtquRl
Afs5wZi+VTFJDEQgo/az2P1ZgeJ5Dz2FeYwoBTk1ZdnKkrz1emgfywGDTwJyMEjr
QrSfhPrYLeSTseiU5g2V/1aaG/8XLbf5QWGUhlFqO1aR+uPP2AQglQ5zm8cyPOy6
JNrbplqMbOG5QEG9TppCWx4zu2PwU7vSzMQLK3EIkFeS3SSG6GNbS7lmoBZYHWqM
jwqb/7W8xkd8klCcyyUjlITRiWUMBHzR+7HnQ4J0HaICSArXwHlCpu8+rrlgd0l1
jTtwXA4XKAGDIZDjZQULMxQRku2HJOyBVtSaXlldCASPJQ57RPIvMBCu55rnv2gV
2H5XybabUXtmXw/te2JN/9WvITIZrrXR+cNKKytDU2+9hFqCGuM2ngiAKdAdMjTL
Ru121+t5boQJY9c1rXfOQ8ePm10JSyLBdhPYUb1QghL0WbDQSI3l0EUhxXgnaHyS
vO7gjnAa50y5cLwiQwjONTTpJdxK4Y3+aqNUBVIpjLxI/1ii1e/2U3EQ2+OG4WR2
7rbaJgm3HMf9/uvQrZ8z3Fzpp5OAFBI6jEqmq7X228COjJ3l7QJCdCj+M+bxgecr
dF+GaEaLALxFVFmyin6+zSrXlPzeLd6e6sYZ8yQyvXvul0+gfJQHdQfvtwzTxGux
oglS8gUGjqwSQK5IRt1gPHeJ+SaWF1JB8+AsxrUW6VomSiwJ+J5jFfjkoBABPJ52
l9UJagN8YWAtGrezpFWb9XWq8hKX/m9DQj3kkZnkKZzCN3+ob/p6gRxKeXfDSP9Q
arxj942kAGgOfeZC+5mjvs1vJv9NW/HZPHavcJL87LahbEimdLw/LafsUFA4JKwk
LIHmrUeo4SEtVbLJMOWGDOWNqy+OV1JOMzK62p6YG6F6dujbymWjzZsV0NqHi9Kd
R+sV9f43vbWslMwd2ngdNm2dNl1E3JDRZdoODu6sLPeeO+jThzXbWRX855tXOetz
wiWIKsxjhGJ9vaKleuz/RvXM0OgIqoZTU/fZTeSbCNrxCl4XaWbG8WIF2QlkZELc
iCXJct7uoOQ1KPFGkfIThZ6ci7NG/2077+LeFyXjU5XL5wKzGdwQW4uHL3hcww5u
t0hsf/WbHpHTt3Wm5JvE2ExxobrZJ18+ejRXYGbpqyTwoD9r1epH8URUHlLpyOwA
vcvGxiGEYK6x54/mY3B1cowtMaxBLkb01UcUYJHAiPKB3M2+3t6pSPfWzQiAiHod
6QY2TFQmDIfI5bgxPRtruOMl2sSixA8FIzRXhMcUx2pfkPB0Ehoxs4oRJCkLb7aj
PiNLzA5lcPW1F2p8fwB+xoVct9bAdKazaCVwsgPiV+XTXX/SXwXViu5YnVa6Qer2
LcewPPuQk6F5HwBsho63GrXkUaCBWqgRGvckvgKL1CIxWpS0Ns4FSAB2KidVquA4
7vqfneKoryifUeVZ5xxGct8EZvJ9OZDk3sWwatv0y6NBHEGjsyVMOU4usgMDpDTT
igl1F3pQ0oLEaAU2vW3MY5Z0HpwFASxCcIV/srjmRZ5mX4UGxwsX7FNsaKYUNERc
m0LBd2g846EDYqok7PptH3a1kP+nK1BF8zQ4fgiDoFLJVp6DTVzPozAL2cRAFrhh
Lnet6L5qFAyqKBm0m7SF5tYCr35TKKugqco0X8cuzyuIQzLgYfDm5VRJY44Pawe+
i1ZtCG2bwtN2Qk78yRBibNIjsmo5FdVc8JwTaaRZ/JtqBIlhafndH/uO9fxZWBoa
4eA7Xvi+MEi2FBFkgTLuvT9gjZdalUfYeCqpkzX+D29N38qNH3T+E6WF9w4VrvZ/
jk5pSNJy7ZtLk0avYX3TZPwN8ATl+Yb+7LhMw/jBoQpBAt1YkpJ/xy99GHrzXCGR
OVB86gEfO+kmZ+5du9REpAn7SkfK/KQyrYICK/dcXA1Ir/vTBztbzWfE/NzBwQcQ
at1SoYxm8tPryzswDUSAR43FU8Gqb2BE+AgDo5GWE5naK9safglzwPNEq6VV+llL
XKQsdBehYHEydTTb6/sAB0LN+dB44CiUZNAO1c2EH7JO3015R6R4oSj2A2eKd61c
MQVrHVQz7pUgBCiB4djd5QQbu7D1LQWWjZhjmV+VgAT6wj5b5moqKz28SMUBpr8b
c6ep7O9hefJeiMKHk614ElGc2qmLBrjCNQ6dSq0Qv/Wvqa5pOyj4uNd2w3Bt7krA
ZZDTTklrHrqFKIwRU4iVN+PpEQcLG0brXwF0Fv4upI32mzRPB1dyw+DRLWfM9KnS
3DyLnpKx45sOiNfKWYDBvysk0OLHKvFDy6b7cILrBCGSS+bNdw1EdI8hk8ng4jzi
m5PWhfk3+rA+6JF292CZXaUGMOEpuq7HndM4ZKze2AuQ0l4vPSoNfv9MOzJdr2CB
5J+ii+NjU2KISGf5JW1G+T5vW5ugFUjqCB8vFMFulzV0BJm7bNOdCSeoMifARkSB
PFazHBFwwtCCDeSzbMBCMzY1iYYzZbWUTVxmCC3UurX49sIqDPMJMkoFupol4j9u
8T9OpOuMtrdNhu6DWTmQ9OfjNKVtEteBSDU9dr3zl1QTMp0Ns9llyIHfeH/syQMR
4TzXU1dUXDT2nGaWzmI5iQrOIFAKTtZI0HBJSLBpFXXI/8MDIc2Z3A2yjRhY0W17
xxS+fU6XMY9O5BII5WoJhEcM9lt7Sn/MPy8Rcguw0s9hEJjvicZs8qVx4+Gua9Ac
G0onkSalQeTAbnLhFfxA5XNGTi2LihUdKNe3Aql4BqL1BOk3mj4rVP098ekKtWiB
ccPf0OmjqmzYJXJxGnC7ytEw9nnCSPZUf1D2JFK6UW9Ay7omxrLY9wpa8L0Axwp2
D4RO1wOVOdY8dhuN49kgmiQZ3LC9ydYoyUb4Y5lweJvbVo56A5eyCw4P4/fT+GPa
Cjsi3xpxhm27ysh1rFt3WrbDVO6l9CesWmS06xHZwjCO4PtptQPHxFrS3dVnqiRW
I0m2joeNPm82BY/84ezB67OS886F8593JY+W61TzFgpEjbfbUrUtwAIqoyiisfBs
uIwcPmOQvlCNDyo2HKHfzpsuqDv3rXlBwa2IdOZRXo0JbFZ83t51fvqD4wDGH/Rc
1yuBhHlaFz+CrOgU7ddctV3aJNt/zPdlkpLPt3zNhpMcIZIjUotXB1hCOrvlX4We
tWuiX3SL64Rmj63DVEP6vfBrDo1yXmQtXnQiP2TabP/SFPjdGUk7evzTBO0VzfUy
wHgrxPtCSqd3M6m6/9wiws3eucMFvgTOqgvnfpbGaa8B24dU6O+aPPPxs1GduI+O
Ryf/eWPGMTWHlV675DwqQLFSe1q9SMU06tsV4nPSSYpYM+C3YRytNyHb74dSRE+W
c+EvW9vZuhwKwiTZdwRzU1OMCXD2R6eHQHTWw4oANeVyHxoYBOOx7jSYmTU0QDvr
4klmK/I0hJ3Zgn24HE+AntKD/k4YrTubDK7d8XvxHwaWpNoeDk+ZRQKXTtk8QoQJ
LSFLEzc5iyfn/ZJWMZyWVIldTHDw0q/FsfSNJl7ivhmkpuERh2cyDwfBz+ro4F6l
ytF3qxdaqyeQ0Ev/68eQ7zt1fG5r39xHrfIvC+GECFeWNw3yJ/C0dO+hz7fumoHQ
jBZ7m0oqRJRTxZ4HyI4fFtqZ6tV6iwtI541uBy5WzFMkk9YYOaZAc88J3cgMBKlu
zltUpfJufjP1b30KQwHQN4IyKgp8Q4ZqAUhgrsdq/RP7dvOMSRa0iF+cAM8jajbp
2V/E+a7/rmbB8txzQixK7RIWlruJC3+a/Mpn8tj7cIiD9SzD8PUrfPbDf5TK4GNo
sLsTmcu8gnAH09UuxXIAASJVe1Bv82Cpert/O3vGmU3PKBzaoXcIDfU9eejv0D+W
CZHkEtbw11mfBLwgdUJpJvbdZaZTyZEXeewAfjtRX3GLRC6/bY2EdbNuaZQw+/ii
FVZswoZi6St1/iZ7uHExlH6aeScS18eiYolRK8JnRCQxvCLzVWo1c/c8e0ynTL1F
TfSdG5XDaBrwdppY8OGv8TkDYtsmLa7teAdCtq1k0KuPmI7SrBS0K9qzj1fYHEmP
nwwU+3oJONvZz2JVwwDq4yclAFUS5o3trqwzYo6LCorMn4E6FQwMJ+90kBA3ddoP
lH5V6JT+6xRrLOAQfACj9LyyIdhN+SmSDXrzpDHGQhXlbZVxQFRE8qLAsvLGQXUL
PYVGQGoCRTCOWlzNC8OrT+eFaVfSeBwjAMPpA7710gtZQiJ24RXic8Tx1H1Hy7nT
zjr7/n+bezI6TXpk4iu8w8Xr95yIwUFe4HiCPK+A8kcTZAclyK/Lc57FCkT4WbyG
I5CMQYLEIuDv67w9V19tN8W9cKEKTMk1f4x9pZpMenFccCxuujjGNCBW5qPjf5OB
6HL0iyUH0Zh1evuzm50/Ouu2lhiD+gUpjkSRmvojzj+j3qqKUNN2YTGLFZex9WND
7fm+/DzRGdz3v7meAKUgyvNkY287mx3Cwl5PQwQLVVHnYoRsy1JpF4TxbUyIMOGY
2iG9SxeAEdywPPsSUu2FdkgJxNMLf0C13lXoX5G9e8RKnnW3BEO+PU3hOYoTCa+T
o8CZVyVEy1VdfUAOGijAWOjtPKGfchzjCoY8ivWoeo0t0Tm07OvbGpFU9nqHTF8K
ycP1i1wkgkIqvqeddndWmlFvoBYIqta5uMWGjO12hidfQWCUARufsnOxHqrETIQP
6MPl7CSuSvO8VQpXuIQmbJIoWvP0AbLlHQvVxYj80HbCwk197qbLk3iUQZSe71wm
jSK6V7JGO5VLZw+0tJg82YwGkqOLjv2NfRpevrzzBGAmfvlStCL9MAScG4pNzkbM
FBZgXsp5+5qBMDe7EZipJ6z1l3sGflmqi+tdxvgewhIaGLXga9Tj9Awo+FztW6aB
/uJhPWelKifTNjM/eWkY1EST8vUAFephxN3/ASMYE5i+/9lrF1X+Yz1wjZRwOGqB
JSQUgkCZToEw/gAb2ez7V46f/VXUHzD3kswawGJJMsojlWszY/5w+405shhbxztE
iAarNm2HyFivU87kv+lblbBoKRwReu0mCVj27+QitoMW4fAJSt8bWTMj0Abe5B/t
9Gew5os1owemsGhehu8ttgHvp8sjNk/97+i92zr2D8lc9HBzjesGJbeVbIACofJd
gmaxMcGLnpZTWAJbl97ePdhg55wIK0HhBfobKySVviF7a9VIZIPMxwJno3RFfNha
di+m+Dew57YHjjWlni7tHJIQOJyerlunmMkLheNe5eFs+e2zgrElm3ojRRaIBxnT
VW4klLmuRgaxnABRaChc4LWUmlRnIq93QtkpAbOVkIClVPCaolNcLB3GT0yhgnYK
bBdWge3vEfceY/c8QqvYYefa+wDvnvRB9yIXxiwjsMdCM93NmvGcR39UVn/Y8sYg
TaYAuUZJdYx6s/OPQnRSHDExx49HnxKAp6sU1z5qOEYu/H/fdCsaefc7ZZ8yU/+8
mCv5dYaoKR/lj1hFi1EJ5sKoK1kPl/ruIb6/KEY774o/hO9Tg9zZ7X61o+Xh1aGd
eBm+I0PEiPaL7tvqqBSnbojHZYYPiZzs4vl1QFCwnMz25q1/WcguHaNvG+zoMZDU
kdtnZl1hGcwoLCdpPw0rwlhiaMSG59U862gavERBWCW2/Zb5URd5JWbiKESB/P8r
AssY95HGPcbf4vHeQ5sFOwcgPDePz9YmNgLarD3JcmaYV2lfhEWSlwX20Hzgo3jH
VmivyJCrjW3M2LDWJIaohuP+pDaXHstrWVwpFeNoo++UqLAQ2BQYh6ONZRDFIsBO
nH+H0DKx+8H8Yb27sls0Onz/m/RajKZFAiUkcMKy3PY8h4KMIB2SfYJMtSFxxHQG
df6iblg2h4/DF4/fvSYd/pTew6uPgVNvbml+VUV6C+y2GAZU5/L5q6IUmrTlhkXE
Ctm8+cVtrxqOjFV6P8WyTox6QjBl8zvjxcivYOAPoK7FYWr7joHb+XrYa5FXZAqV
9M01VVRJXjtfk9yRZB4w+cWM4E2s26IpQlip2B/snZnK682T40sPt8Nb0PxkKHfo
DkA/q8Y6/dMQVNHhwDooYdMPATtoDHYA+p5oT7rglRtr5ADBIl2iPr7Bi6JcTeP0
zy7qFJGPIbATPqAV+3a9IZJs6w3VnDdeTv5YV7GkdkBZFWRswwN9Md05sbudiMIy
dbwPbo+594YJRIqucI/7SCb7EtR/ac8cWOO3ifv9yvc7W5MZ1/oWTsFbyBMBDFA9
rI2DfjVeko61gky2q9x1pp+dvs1WDsV/5BDp+jBvq9fyHTig6vxMCiFdczd9Pi3/
hODmPSRhqY8o/ssFoauIu5HpETRvZw2uLo1RI7ZaHEm8MLNwK/hmbVY7qrZNefd/
uWrW667e9SB2WVqZn7MgNd9GVWniYN3CFpSCl7WIKk5xDpaLIasswL0eIE985/0V
nqdmk2JG2rlHJbafEfTMa8xYvlyGCLVZO3CRltvl7B5YRi8ngTS7qpHBRlztDURT
j7lS4RsC3Dmc1FnMrfd+l/VNXit24QowT7dGt8SNcdBXRdVhBrp/wdir8yzJuBmy
qZcmeGv9hS8Yi/dYqUH+kRj0JI/Hj3EmzIY/DStkhsuB6lvCS2oOE1lYF68gmrTY
naWHNlU80CPn2jTQv+kedEYrIvbMpFak4R2hTUt8ZRuRkLvs+qbeN/JYNw4tbWVC
x7IpAFxzFhZ77enC7NS2EjbnbwBrWfvIoPMDr2+ly4GBQcaZH7dQrC855dexeqMn
6TQufEROnGsYBOzq5Td6Epv/0nRJwpSF8NChGu0Cw+6pCzrv5OH7HLNcetsQm4Mz
YZCil5mPzlW/v40bGMOpKexJoXSUzPyjIVE0ZduOIYNYIeu0JLdDlrByQEd3BWJN
SCnJdNxeg3+jJmUafPuV94uTVl76E5D0xDdEbmgCXYNgvKTIE1rWDybEIvjtoVfR
CQhIpe4uRXNLDjvy9D8dTGmdhXIKGJrUaBhYwpKfBKlhvPSj473jjibxjVc5hrKY
gaHerjJTSd0K1arGN9f/L1x2cxYX5LWDJAf0j9mQSVCSBZMtCVuhzRWCE7sFd2dC
ckmb73adWBDHyT8wXzFT8y9ZpI+/OUdQlAJ2yDnvvTuifzWyF2C1Hx6uGXlDCyZL
hDyoq2RPiH5KF08VKZ0X038rmhLk6UqPAUL7JXeDgw5NP8SajrXo3fCIn/kEdUDZ
Eua8hmRCA87r6FGNMYC2cB37cRZBWAJOj4R2dhZw6pDlxYsNfmiyrunYjg3/lAzA
sX9RVnIyTzhpNBTrNyO2zx0G0KIbEwviteSQK/a25WWxJ8AT9/2h7tIuGHEJG5nI
ck6gGrVJrPXX/G2ZFLUNXqmFrIOizH5ZfJN5RFZs559jhadgbrWgVKspiO5cVmgR
YruMve8O/b0TyYUW8Lgy79HW6sCxaIjeffkQYxqSDshNxn3g9OJAoeSVH3PzQIit
yJYifGl+s6YIapUlkfnpxp1nKTBQtbnrFdA0VOuNQ02P86tUDDRfM6z+o8TfvPJ7
eM4jarycbKZoUl9gEZdgFVpjhWD0LPIYEed2DWyV9SHqYkFp4FJA1RnrfjPdrv9A
P1dPKnnfgiOrIpKpi2JK5nDOOm9B6JRznB04DXN7x9jPLUylgSN/vQch+0/0TW9R
DphgJAPToXaRYznoPAQ7rO3yM4YIiuj73TDAk4JtnlJ+uOKg4neNQv3eClUQ3odU
nV2dMy9E4n9IU+fkv9Wycoluy1zXYFGUSAjLO5UhkvgzmG1YpNlz4EleVyzui0mx
aMc+ibDWuompTZK793ZbKZKj7dxUAr0btL1X2zOIDkDl9vuSz1FjsGMWo8K+vUW/
RItA7LXihPO1dAtnep4qAgrqCmvlasj6Nv9/TPQpX6SlZXCiUqVvx9crg7wr8Gf2
bAMEqfHd/vMcpccMoxhT4f6gp0hM3CSAk3dVN7jdLUTmxzpI14NyfMJTSKatI4dD
kqtLywzUGkdanGdoTuCFS4bsBZEKBXGSU+ejjiXhP/GIo//L70TnzoNvdzLe2X63
blyPrmR8A0hj09Q+NFnUrkt4eOU5DaQG/RWJ37SZzjDH2W2FwvBynVXldIy4ZjlD
PlefuIVl0H5DLyIiXyLOvqFSNWmtJN03/G3BFXDxO4+9SBxK+TuzqO0dHb9aQBI1
uWb5F9goyYbtjKuLyiuxi8GTjsfFxIAMPqoxrW3mo3ArhqfrU/h9sPHIT6EzG511
Tz5/rHmAjlg0c/DlorC/qOSbiPjh0DlFdH1fEIqPcpua2bSTv/o46CODKpDkx27S
IAYChkSZLugNdvOWho7GI1R97X1E+Ec6eoLGCVqoypK39/INSPOCKzPtR+eRByPQ
0wnUJQ11ECihYeq+0UksZr2d2Yz9zn7wHwVsioidCpBv2x/TKsqE6xAuDlm2J2Ki
I9xr99bfZiiN2MuuZo8cT8VWdZ++9Qte5EMRNW5HsVaQIpPEbGPsrYr9Sb74Dy6Z
UzECSo7CgJfHuX8YyLB84B+xOCOxSvBlbTBhlF3uj4IIbeYxU8Ma+YY5TtlMtTfS
R2Jitj64jmNKN8u+TPfpyAwDplk+/Cathd8OtwAu1bmbrnhK6xL2UsxHxqshNw1z
+U60rDbQh5s9AE4qBvGljKVDUL/XuQ1gmce7FHJfJqesX7bcKzUOS4vxsWF8YBWN
sWHVdC9aCUp5Sm9vFWaCcgAH8eJDm/9GClziuSd/kgZX4oqQO4bCaKBgcOfq4vB9
PI2JszU5Djxu4PW66gQaIjEtrEuxb3ASDSUnyIDWlcXgj8NSLpuqqAVc0RV79tf8
MVsCiBavIIxLxFf6qRpQBHDYkli+EqTws2U/c54Gd90e2R01RixbWta0YNamz4DW
UPrMTNlnsXhgzpNoNRMX8Fnh+QW2d4be1FyXtjF94he1b3mGOQm+NzDT6qoWL2W8
7oSfKuGLaM6hapU6uLxN1nlyngzPylb2TC1LVvnJ5wSKImAtmNBq9LX22hIzj6dc
yIqVMVDdjtn/twoLUft4Ore/0QEb/yHpjx6obP/+MThqWOAqqiwLiM2C+AgIkvFe
1kvohDZ7PKpvsJLcpBp9t2xEWYbNXcxgRNeAjJz7D7B9/UDlJoOsgyNoPO+vRd1m
i6BrhChJ3LvCVCp3OYOBp3imVOYnS+lPyowqCfsJ5LIShELM/XZ9XcSeiXMQgbow
UyIRLVZT8gzOaKShHPEB9JHeNYLzjhPK/LdQAvY5RxCJBxlQyFkVSIcSmUPaQx+1
RXtk4wCCcwIFAfhvd9Ks8PSXRMlAUKKgAcvRDQ6XAD4Rxl/igF1xhCYqdloLvZGv
YU/GEwc58fwwD4HPKlMMjlLcPNU+det+0Ujwb8WV15gRsq9oNgBFi8sSNVz6wc7l
KerDUiSDPBqKmuy0zqgiAkMsNjAspSPYarZCVUW8NEll6t+6FuAw4USMUKsFkoIy
w0TK1KkU4PP0Pp0YEY+sZQIXfgnVn0IYnxkIf5/3Uv3XfF/e1UCqDQh3sHXGazE2
LOtWRTK/+VU6bKmTiAtoLdaBE4Kv09WAM8gVTXUYKgs2GyUf7TmPOkUh+dxynOF6
T2UBMbLzV2LX6LSgVNfRS5x5neIoxDtCGJu7cop1BkOlxTAhmUZCmobrSvD5xyOJ
LHBee5Go0PsQQixgXb87VZHPvh8g5uFT4siPOMMo0AaXJPCMrW5Yz+Olp22P8CeZ
cztfrf6W/Lz7TtH0LcFxx2XlMbemKH8IC7l16tzo2Ibcl0WBKT3iiqecGlmoG30I
wNqPyIuvkaVTK4j9adglXrksPfHUpUmJvFogPmhNgZkZU+WF9HweJbJii91HPYLW
OQZkI7+KV2FFlktlEF/DDOMPyrkY6bo7yjSNHy9zYu+CqrNbrUESoqL8vPpMeR3r
Rbf9HAJHtt5kCCifvNTDeGkmB2I2CLARka+U7+kiZF5Bt28+YDXrqeuMLWOS0VSo
+Qg72tlsXSErUXySWn+uG7oaPo7pZrdb62RXKDuMYdugOsPTPUd3gcZ00oL+AdWn
dTgdpVyasDEq8ctI0fI9zWgLwVrwa3sXWvlswRgxArDMk8Gho8vyZqXNcQZHqY+C
c/7krPvERAg4u8N2l4GIOTRpdKn8FIFnGXd13GvQQpl6ZNctfitBo+K83tVnDVEl
EmyJPtv/9FjF44IjczKoSHidGRoWdYRUw4Mxj4Qjv5+MqIDjl6BfHrSCsFi2jxAA
5pFli7Im/TCBc4fJsRsTg7Re7dm6dDYuUwzFgV+thncDk2er1KHtWJnIWp7kdYxx
6BvuAHu4MI4do41iZaDDDYYFAviZMIPgs5Ofo97v+PEgLL32kLYslyMRF8D76w/X
s18YtK8qHJ2vZOzyubud2cyw++0nhZAJAndNwTTdh0OV9GUser9ZTrYwF0PYqhhY
WJ7gmhmq753kiEHa5p98FOLcQA+b/OmpKrgIzIvoqsKglvNU2jbnQYloNr1ItBFu
EhntzPhSUlSsMZBx9OoMM35JGGABUL0Angb1MHc8Kzktigxx/PKLWcUke27jDKiy
5BVbcxWo7hJ6VlVWy2uzuX1il6vB7EwRH4jJG22PxCfYcVgJyVwiu0PlU0z6XCTd
jz0Eo1WJoAm//iycKGIko/6Jy+LbIX2dN/3Lp70X5AAlIJFTqYuyg/hphSzgXZMp
+tnAnMAlscOYQPNiZWN1LfapeSzRrLrTC5BC0qF3FBop1OIDV3Cxkvyn3X1Ru6S6
Dggj1DBs+612P66MJHrEjKzr+F64cPKOj1NqMVAje0waPkaOP4TFzvy9zRwnDC97
YmP4t3EFcG3KvjplRgqjLaRjYlt854b/aCctcuwUt3Fl597GYi2unrqtjyPolspr
LonqbKpPJWdPVBQp6Y9eKr0AMEt/lPxUEe9m50BVljThutmQZ9ASC3TRUkLFtb7j
BO6Bf6/wegzIc3bFlxAkTKiObtDdnuF83OhFiLLG/lLzarOQq0ezUUfXB7HVM6TV
74qFNxKy6kY4OzM5X+I2TlkiY+vP74REPxrgEKngxT+sbAghC4B4tUtQyFG+vtX8
mLk7gY04V5pF9a7X3Wh/Xj0XupezEMxCMIw3g/PCqKJZZmu0nn8bDMhXCWeinbf3
o/BcrkTCDlA7s0SFRcB5JSTBy3joh7/q9O117E0ZC/343b2CuU+MqX/Pi9YLTQzj
6H+yjK8fCWLqDN9uQjv09hAHn6elkf78O2GtZGFsGQ0RfA7ukXNDzF/dpXRqRblw
vJL+5uONI4CvxKsSg4L5BtkidPXikgRcWEzRMydAGwxBn9c3Mgv0TwtvhzAz56CO
cpyKB/5GAd4f24hNKUMUwDighxVhyPrfQ5uoj+C2lRxrh6RabCpswnuOBRZLlWVI
zZTky0uKVKvoO3cWKskFbE54HWNlAQG+WJhvY0pszc8HWCxuvYCkX8+As33x0uAS
ghM+beNcJFklgAt4Hjbds9nNvUWuXWGyhgI2+2GraU/45FzBqjHIvIEVy3TYWocO
k1wtQKg/DdeMuWfmz0lV9gpoCfOW3U/nRcRSg6EkryJldOhzZEVg9C1oCc/8kI7P
Lxpbf+E94Lh6/PQrFwiFWeLi31iTL2DQknNjT8CT3nW/iQr9hhCVHs0xJx9Z/Htd
0VenkZucxlzhF4C+3H0iyWmXpKNYqrUBP15enRFX7rY0zDgDYQZ3k9G7iJUxNdZg
IaBN1xIs2/0JbPGb4OXzzXSjJyduVgNPUfU5YX+gVcuK+8aUNxaBMtl1erFJkFZP
DouEBr0WD9UCUO7ZUbh4hPkJqCa9IJb24u6R5QQauDlRB9tUAuyckHc+puW71qO5
vAXb7gmS75hcG42sBx/xrGvD9AxXUoFVMUrwQSuzSpdvFN6/VdQPFfRXG7WG7oyK
OazRSBkDsjkXMapv9zX7bm0WFuUCv5xlNZE7NLeYqhdIF3b29cqtDDo6GVC5DjsX
A9A4RnUL7uuegs9zkF1vhtwG+CblYy8s0qvdlMBUjH7RkbV0emnLy0MNUec5qryS
yosxJgZwtCsEdLzP9JpmTemJvi7cNogC8Kuf5iNf+E/cOxuHZcHcE4mawYcEL4xv
rzvRpxK33xsPmeUxnD+WTmc6IhppItlrD9qxp01g76j+83SG7wWldt1+oiMZ3VTt
dW1BwTLOqkN9Yj51hsHN3x1f9UTFp3mq9jt72K0NG/noJTKaaf4Oe8iampceMLfw
e3psaKoEHUSJcG1o6hXxmpvK369HOnvehgFe2HdmlNji3vBkXm4fZoPJ/vDHz769
tGyJqbgs7cGczUeRlLA9fLVV2hq0hOmkYa4DDmH8y7Z0Ul5cAbUf5z9U8uYSYrxh
bPwyPttErgyuD8YRc8o6Qo7LXcQUrraBPopaDw0BNF4tuK38H5jyYxanCtV4E5aR
eP1wlnadQhqrxoxsKe1X5pE8PUJBUEfyHvspj93UcAyseLCp/l5eRA0DHQ9bX34a
37VS2vIF4CRKXBnauDQa2DJKPfiVeKS6SzlvCl3FKi2te0w6ZmbLU/aeNE7VWv87
yrZZ10Zo9CIf3Zo5I7DRXs9v0qS2g75OFcxukzkTIBlU8mj5tv44INlzQuYcBl5N
Tjp+ntudgAOoMWJohsp3u4kvzNjYfbS0GqmvEFk1BQaNT4Sl1T7BT6lUq+OHgiVR
vkiQLjGnvVCnTg3s0ZzC6R0pb5QgRoJppxY+j7fc//ax5Jm2ec8TcMX8uZMV1OFi
cFJ5uTN6nM8eWe47vUVe0rQrz0z7e5d30owV2TcWlzt9MGa0pTFlpPmccQYg24Ga
L99QFdQFZQXIuPkXnOFCiIZ2O/v1bHGHJYd4KrFmq2jlvfauQvnKId9FUPHh4NQ8
6Q8RpElenMiGx/cjr+dRscKl7dZfwP49LDmb4w67FGNvXz+PdUI84PJz5mutYTg8
FK56rQS21CnBEYaSb3/M/36ZYKz+CW+XGgsxUJomCROCnYeOQeJJFXGXutW+2Oo8
8qeAj1AxJwr1AnHQeI1W9cO/ZErrY1ZVCZmTgZxxxh7EPneyDiyrGZ/m3zPSh83h
9+M6SnKcsSjUFjVoIHdUIgkEHGmU9l36MVZmMlGenbduSH8x7xRfr/UID0b1zHx5
ENvE8VTysjgGlnQTCLRR4Wqos6H8Lfvbn9vX51/uBzsLwq1uTA4/4Ff1bsFjHG8r
xlpt8Ta3FRa82pAr7JjynaUB7AXZu+tu3zMSKo4lxJMlW3ukHuItGrjEZiWt817W
czYjOHMK5w0tsv9NhpCXEeuTPAsmTKqkfdtRgvtSgdm7AMdFrkONM8AmDrsEgYwp
F9t7qaN+WRbQO+WdgPT3d8Agt+hd0gGGcQGNrAQ5vCNjT6ITgZ+/cXXHMqU7LyiM
vnWqtV3jHvHhXSc+EigQX0+zdfMyF5d9W22vxj03Z/25kuGxksPh2JiywowHha0Q
iO8YXQKClE0338c8ZXtOCpb30xmFwDehp67BtsvWTRzmdcJJANbK5D8S4zS/31BN
yxIToRkKKJ4AeCwk+FtvHSANVQHPw4p6R+Wh8Wwkp8ewYy+OdDP/+wN2jNyEDvxZ
g3gB6WEi5Xv8dbYCk/oBoRPpjUeRVZvrwv5dkCJj55vFCCFo8qhIUC6/WvJ1XSje
RtVltgQTuDg1Mx2bjmftZe2vKMPaV9fw0jrGDY+TbgWCVxozqV5/NB2MkGJxx1jD
bjj8pS+r8ufmWAXAg2SrTNl13ZCKI324fW4TSGurO6SVUgnIPZMMQysWKydKRSee
rOj80dRSsWLMTu/w1dfk9+MVKp9y0auQXnkQuv8AAtGL/tThumpXO4KFFUkD60hL
aNBxH3PeXgKwSyq+5N9oh75ETGLEe9lOPGguZ0T2p4AGRli5jPfteSmwUuVxA2zK
apfrE1L5ZYO3vUfcOyMsPuKY8OPR0QNZOG4Avq/GVWekk0LbUywISQcZiOq6JOwO
wwwli70tj3ACalxkw+jkNAdDJAFSv6GfKFWyN4JDZWSYLK9u7CbeDvPwKfgtQ6X/
pXH9BC5VcnOC+SE2i/ALTXg+z3lAcExAuG56qy1n/aCC07r0eE5hy4v+0z/lOKbb
WcP5ec6zy/6cccwPsLNgiid0L21AZsvZhTIOoltQH7bVDex9DxfBcRaWsQt3snVN
b7ihMaDOcmVtUk0Shngq9fazC9ORARg4yHxz6+1H1k3OvjxPbY3VgRDwptdoQO9E
BMN7fylRnOnGmbM8J2WY526bKULf16dCMRK31/KQGV8TnF72hR/uM6ixo4ZpE2Sl
WKPzdQTqraG073IrnzNN1Y1jIIyiEs/kmR956wxNT3psoZxPwXfeziYsFfoDqdVw
OhH36Lu9xyaJKL5jTvrAGrqe39wsFaq3AoKaGVMEyYpLy0nHN6z8RD7frfEtvZQ8
B11o0aTKM72NyJtBkfYqyjB9dQyzGS0CbTNnoBcOPZ55w2fKrvocIZ2/uZmcIoP5
XetJIY0LZiRGhz4U3Uv9WQGePZH5JlU7lj0aXMAyESk//dZKWI2VE7wgU0GHIqBD
UqDFMKA4pemgAxOmbg0CDEtrcsPfV/3TadVQoIDaVCgLgzFTNHkc6+2r/XVRr2gS
sZrUNBbTmpEgKIsSgf5HvE1IMLM/rKUh4RYnW0spH8iLhT4Lxj5xDifbTD59dZxg
Qwk6uXLttNJA3JuM1tEW74na3Lc6jRIUpccVGFkORMgr4uLLot/abABifp5U+462
IkzesfXEz9+AK6kq09hw9Q0LB9OAPPPz4Lik6J4w5+xNLBW5hTQbshho74tWwhRs
NQdUS+MUwufJ2VxB06boOWKN7LCiCX5QnnpJ6CGlMbz/is+U0HgMXYJndggDo6wK
XRMIu6IqQ3COFFSpNovGwbuG3ErDGzjA51is9gvImzoGyAZdebnF7Yv0Eqbv8ch5
stHTNnMQCYGxcNvZ4CTF9wm2FUoYALSazsoJvdfIf7WQwx4s7HqKaNi02l5mOxsv
TrJ7Bmq8Pe1mMS6l1vpo5UPoNGdOUTlItr5t54sBHN66grp7Z/GuC2dQiTSZezOd
538DkUcWxwlOUhYP20v8fd07Gzqw+s2OmwqLpFEUul5p3peHaVcjyts4j74pt7p4
nfYMbVxbstGcIDUYLlKA7SBRjWlY+5idRya2GdslUQOihAZ5oTCgIzjKVuk4P3OJ
XRqCTd5vOsNDJmJTPs74Q7uYIS5ED6XAcH9vd4qVNzdLqEUXyoSGmpLXk3yAmEXC
0qhJ9I5Fr79+x/pcqm3EeOXafT03QqkeG24it8EVWmHHsLEJGNXO3YSS5o/1aHyr
kGDT+R4JzzpZC0WnPD0ZRReRk4ObstQFhKIbheMpHlU+G/Boxt97AjJemEwdVww3
+bMqM0yxxYc14TUq+ltW5jukXqAAiYfk9IgkYFAV9vcD8ysZiQ/dH0e9ktCCAgr+
nkHKkRye4sYibLHjqJZGrhkVCCynymquVyiWN5myO7OT71Zwi4dbwgGnYCK5Nn9b
oWW9eo0sC8IPzw6ZU7tRwipBgz6S6EpsP+us8Hu+8aVa7M3GkbnV2EIQfGNUJ2ci
b4n261EljfnH1v628pOzPH+iD3ZNJ9YX4otOTr2Ekflu8gmv9zhVpq2on++Kwg+i
ehRDODuPE79c+VrpA7K+RpIJfOXKT9MutDYSxFdFjEv78LstRZClHuheTGexwQS4
VN2blEPuYikIXuYdzkPlRl49CF1ROoNii7szesTZgtGBXCbUSvcZY+K4LGq/NqEs
eeVpnh3fpJ7+YOcMCKOUehqfTOFo2edNtBeRm0115vO6/ojkh/zJcKuxgaex9ZJk
8BJmpat4n4W9w4smHl9FjPEI4tmVEIjj+qASsOkaawE7ZkpsPmUbd0WfsVScRz+H
qhdH9Hb8TZCEOV+pwZQR/hgYaiy2ftbFEHjtkI6/Ajs8RQSqQ6BASSAi/ajQ0hJy
vUzCtG+TevKbK0gyMNU6uyfVXlBYQwW8w75Jpea/sBsM+KR4KHiXnchabHJdX2Aj
it0UFRwKbvczRQlh70+tmRePXF0+fE7IuBK37J1gI+uG9ZMNp3Km5t4xFViEF1u4
n8Rui6l0ogCfgmSC+B2e3yp3f16vPeIELKILp6yHJVMuxo75lBMtjXwpcpVsZMcR
hmPmX/+bX943/bJTjw31yOlU1ty91lGkxgDmabriTTJ61ylcFQSj/jUmoV+OeCQN
yWE9aZ8WQVARCOT+FlW0olvP0oXgTe3uHblp7xFaLpTmTNv8UEmh9V9fg3ti0DRz
b1d/OAIFaEiXWgb2sDvEn3JlE4qMLHYeulE0lpXmJRw87mRU35RxkjX/Dw+jUzbx
usGjmKVcEXnDpLdGvV3yjwpTN5msdngaRAtCKxvRaHU7+I8teQLabPUR6fuITvzt
PntTqoAxdG7h92v99UeGgJHNxQGM34snzPxbkWQ/MooJQRocYPVhostAoqaYz5IZ
bpHU1/lDzv5rjNgCPL40msDryxMPQROtmQjK6H0VSEYy1BlOwXJ2Glez9usvaBBo
f2swrC8SNXXbcmxjk4WXKpHCJfoswxliguo+2dfyAs/dN4SY61DmtLJPIoFZzFes
UzGDgtoPSX56X8jaijf1qikzatfpMqe15XZtLWrUK98BIqueHu+yI88dmf68Mv+z
YXl0oJxIbdrXBRqNYX8SM0DXddM04hCsS2UUj0ZZOZFlcSw2IN4Cnqxi+pkAo5OV
k+0SGRAfTG7ENVZjTt2fiuE0qEZkN0SGAF1dydxG67LaZ6TYqjN59OeyKHjLvs0S
5/3RcWVjHYLMtzdr8FWkpeZgnVHrR0smtZPPPZ7ttpP/I2d7mLOTpGXqbv+Cgo8f
3o58vz5s3TYrJk58d34nNZiO000/FGdrD8JrwU3TKWqUpHNbki50QtUbdwWInz9K
57IWM79mZQHeMEWZHruC3RqhWRH8eHdhEZw1k4GevA2YkX0O5gu/l9iiZWXIVbwy
JKH6Sy3tZzhADPNbrFLrTFOUD7otlulUiINU4mAfsjGk4J5kAHvB0/w+M22UCJPw
V4K1Um/NoOGiv6mXD2XEQZ1INWvS12h0Nv1Fber+Mb43s4lLTa8lb/34IBWXyZWP
zU2br7mS5xpGIlktX+QqAkFTqCmVoYUvv73g5TzNftKTPSs6DwBek0CPbcmSVNO3
KnGKhBCF5zCBPIFDUCtxaqAmgbiR2DfqpiHwIQfhvy0+RErqmsMahPHGO8UxWZ84
4CYEjOvsOqAB7TDmfQS3nz69oAo4OUiyvdkbjfhH+7tMYMMvIsVTZaeYWzeiDfBl
39gs1Fht6Xs1Xk57DGyUk60KhVOHucHYqmfdILORczYFEFcxjbv4HN7VWoPxNVFq
+6A2LKPxdVmQIAenwWZR0lAWSs7zarDd7P67EzPdXrOkBif4Rlm8V33pz2P5KFy7
SgxtDAPdXm3vISMHmFg8X3H5WuJrxW9d4H/iUMFqLHBBw/NaPih2uDW8DPsi8fbT
ZOH5H1B7fqQb02cHvh9j3DIq159K3CwMkotaiqPXi14DAydmgjazrB04CGloVDVC
Q4PdavEiIzZB1sr+nYp/z76hIpnXzv/PghLi+Qv+AnByl1xkdN+oNPJjRn2WjR44
QEXdmbA4fc/mKHpSWHRSvTBPugolx6CwZA1LdG6omr7y0Ct/IKq5Exg0pwSwjEeT
ax3Pl86DOvjUHIuWSfVFHeGgCDbKkjkpSVLwcGlW1yDaDC4hiGijU+ug8QEQ42Ks
mkVw2KFEb4pRmBu7QMgBFxNRk9YOzZg9myb/ENa5dBjm3s2Crf7TH+oUEPxn/A+p
OZDqeKX0CNWH7eTxcnxORy6FyG0XrmCanoTfaTx3IXY6Y2HyjFeNcy71vgf7cv1C
+feAQfBDUU5slnL8LZUYul+IYPY4rAhG/KMbdG2hPtUvu7PRzLPJpFcoG/JlmLp1
wdO3RZV8b1e6oF2/FG7b8eOGC/Vx0UhlBOrME7YN5EbdEaqSGJ44juU8B8ELU/ga
Tt/2xD/nl+ttQy8SjK5XIO7MEyB3TWfmMKfQ9GOBIJFdOvfHoLYFayNEjd6428yY
BHkzPIVTwFwZagoMrtTXsa7uNu5DADDfjvNRJ1Scp7bcfR0p60ppbSzKkv00nU1M
E10sgh2rCR4aXbF4A/dWjadRlrwH9tW6kQj8XKc2Mi8euMo0krSwSM3ALi7UBXzH
ZJMpPrkpjYiyghEFdxiTVblWjVuKy2cXS68BBkMZvQ8G+itBmN+DzrqD540HMKhd
BrMEmY9zseJWud3uy1EfvW0PiBKAhCx3AaHNmiJOSunlrj+WPdpvticNhKLKUFlQ
mHt0r+T0aJ27WAIgLRq7r7q4j7wdNCS2p6FVj2RAipgZJyQ9H4RlKpQ+GdhHiarp
afs/ogHhuRCEcWiOw9WXvREFe18oH4DIHiXLFiAIUnGiN/DRShOtWJxQwPHIQ/mj
t/inVJKNDL8qr4GLLYB1rV2gcu/iOr/KZY5h6NwMkkcnErsuNmD/PAIdPqW91+Tx
a++lq6+3wFNJjJeAJ+S7Tasq3/SkXqsCTWFufWgjwytT5vw/oyOxSkiFfSGXAo7F
4IQPCb8XmhPtYjfnyJi1uRFmc4Zu+rWVimgeWxiSTOgkqDCpoPBSNaM/8jrDCsbB
9vhNz6yjHQ9Xx2UIcBqLIZYayWJYE+qBmJ3UJMlCjxOAioc/xpxiP8UhHx0lIlX3
nwVPBIBAv0UW4VC4lH+XEG79xeb+RCGDzLlySmpNc77tfCdZgDdAAgPI8RS3mdgx
HsTOV6UdStMMp6oOHB5RqyTzUn85zMRWXCQEXPmbj0bmNV3qUaTBocdJ5pE5RGXl
7V1v5psJbznqZOefPNeZqk0YmFlwWQIlIDiINIvrNPbjQkYxmfrFY51pVNZyLgps
zTrevpfaXylfVW1MYkmRxOG4tK8L5TBSGz9aUFj9EDuyk0KzuDZsL2Rr2iiCs/bx
0swJO+bYNSdGfAjvwagtVhDGm+bfLSGtBwhg663pOHQYlb0q7rkzShXDdmgW+n51
274Akt7uW1W8KuPfW6SYHkN64Qs+XVEusYkSZqBwF55/bVTa308FKONgsDG/JFU5
ZIhIVW37qSkip0IP42+pjI+uoOZ3DimIAv3WcQUkHeF042Q0jqh9BuJOlnzD0OSP
7d4923SPzjqJsrW9GzG4cbnUbdAmNHBT1/glBguM6KW9qIQO54nahJznItw3PLNX
VyshpyRcLkwEv2Az2QAdzp86QBkpgmT/SlNVJgMCeKMDoWgbhB2M5Qojh31E8eIK
OxNe+f4TtXJaO5ePJJBb8kzZekRRHL5eUaiRGjPlH4TP1DT+vqtvrMiTXcoRMbh6
ihFxfRZ3PBrv+mSsnKrULKBoWtOQWJIwV1RB7Cyrs+IeAiiit7e0Mjuqw0p+qVy7
K5tonTjj4Ob8h4xWoINs0UqgXSdufw5Y8SRj6ngvXeGs4JtpLe6p1SkLnSGYtD8W
miXq6dPVJFgVaQa0l4UjJGGl4FVGlaO5QD5Vm3M/3XkzcW7kEQiSlw5y/aTsikzL
O6/t5BAooU00T5ZxcaXmJk7NPhDid4E6pazaTdFrt8cnIImNU1wPlrg/ddi3Tlek
KerQz224wEC11yhrBrJcVpiKEdLQe4Ijjp3/3mquAWVPpWDGyUkQ1zDOKi5zTOLn
1LKR+OjWfgKOcJ9Og/KVubOYtY/a2f7RH+AOx9O8m1cdAu4GYAj41CZZy1tH8lOz
08vl4JMmfn/yDBJuuH7cuefhY+FCLa9OUOp3DYarTXGRpOnunHiSk/C2rtIjHwcV
+Ja1UAB2mqtPVessh2FGDQih/4x0pEwGfgkRsiYx1GXMjHjw3wpz4Jh+UI5GPb7s
It4bPN5XKTFcpwjE2mNPt0VP6hW02lI8izYkyjzJf7cBO2YlDfkI1enVD7uR9PbJ
kqDsE5ePWG+PSmTNv0X0mGAE1nYKUIdsm7ANH7DjAGTOn3SpDDG29oAvSscIcwzo
uGpyHQaXPr6kdhG3Ipl2VpzTxBtyfFk9bVWC7x3vqgBGYysaodGO7+N1Yq3oJNqq
TJb9xv3B+6ncPjjdomlp5T2VQ3mbyTaKuf7D4+ltZJoFcWnCwFzKjdnv3Bp6+on5
njWJNnLTtqAymJjRk/qZvAzPSnTJaqmo8JhP5dKAjveQEoSM0RLaXJVcEeq6ngfa
WucKBYqg9XyHIUFo9LtY0DUH3dZ0PQdD2JkPPiIgu1BIEDm9SoJPmVup5wXLILuh
hTAaoDkFabdMrhy+WQgP5Xlt5ONsypcY9XxkvGZg8JEnE/Tmb4E5xcporoJHJpT0
gs6yuHDXayIMQP24tLJ3ovQhmBDoowcX85SVDUwzla+3BZsR13bmxIElO7lEm9XP
aN93SLQxvND3m431ZP5RZNjhuN1feU3pacVQvv30kg27dPAB5aKtkehuw8TZNi1t
2AjzeB+RyS2J3l7icz8W2ulzoIfJGYU1prRBWmK517LGc13lHhE62dvl5GhGLtEg
pZzC34dwPrAZTAacEBsQaUfHIwYJwD7v0ORqtfLqk4ikdch5SfU0DPWIsik7PAFN
Pz3Q337I79i+uX9pStG5nJrBGdVsyY3/DREMZ0ztFWUBObJ0wQU/TTFO9IUnBop4
B7ciRZ1Q3BQNrm1iiLnXaZ+Wi6QQH8wWdpJS4vxyTQRm0Kjm9UWplrVT6GIrxPaz
wT1GoVXn7H1OzPtQbgfd4VaOs2hpm1q0ERi2Pxi96R3BKa9CBTUVdTMyETqTmbdE
ew2XqSvqYcjBloGJQE575yGapRqbtk9n33+8D8RgIDMKGW4VnQ8AhZaf/AH2GaOD
KqjqskWMno80cl75VDP7FVMJ2+zMBo7yOmg4yf6IaJdJRm66jIimK5uLwcixFrKU
ZZcFw9fhHY298kdy9pN4sllF+yll4qy9wb23Yr42EVnyzcA/RIYtZTNSIy0IXun3
tzhodiCKlefY12AXg6bt1LrMnEq3JlPrYLtPfYQT5FXB93K4/x9JLiWeOXgaZhse
pxXy5bqpvnNNc/kTVG/o0Gu86pv2DdZcNr07kn/2/5iSw6GCaw9kxWeqmEtbJ/BY
hqUnCzR88Y1WUm+hGF8PR+U6gvzZ6tCw9e0EefBgusQ9oMBVgfL2SOdp8QDMbRYw
lyoaGtwykcWSUa8EYqirv+wcT8Ahy7/uWrB178xlcEPkvgXE9C6zoB/MlqdXZsFD
FnE7lx+ARuu+igMR0zG5m8rqIYvM3mtor90URNlVjBEK3mdxhJ+prBqSGfzSV68S
94btCltWjY0hahwripPfVbXQArJ5l9qwv334XHzGBvrKkQ7F4jOu2YVc8ezz3EMd
WI1BN748HCYtuzpU0axus+2XNQT4um0KqRD6cBVvfpN/p1Y0EmiF1mI7Mphmo4jA
TWSzsm33J1OSJEzYnGn91DbbMrxtrMunxIas0KHUs/ColbRNaRy8Mnc63QX3zUsr
VioK70ogi1N5nJz+qG2StK6ZAdJC/XwXnNEtQQmneOtDM/17AJtxm+ORQdRFRcAJ
mG9C04RZb06ipoC04nT/0jAIoqpCqXUiwVv6wPd1TDyQEXOcneH1z12QLsDMAaNU
5PfLjZOKK1ifnOz1O/gzVdMWVELCBBJy/McC55SzCKO2Uqv8hVXxig7M0M7X0fcb
zrAwxBlEqr/53wncrD4imilr1md20k/yGLkaddE724QhSAbWCxHXNqME1z34/zOf
hhhHH7hi7T+K6fcsOCwlzKq4i6cXgqt37UF3ue5FvmW6o0pwQqxFodJMtsa3SPc/
qprc/HyGrTPEVBRTEHmMtMaEPza/9EAdDER0yG8HxcYKjrbDn7KgdUWg8mpE5+xq
mg/jcj8mqq4dLtdzwLu+gWd7oOP+crhUeP3/DT7MX/N0YW3tMWgAuNE+Jhtj+GZN
D18wC07MULGz+E4Vjpoh/YotBzXGzmqbJCFFx5xBHrh2p1thXSXGxqB3CdzLx/fl
dp7FVc/h/m+zM86MYleJzutiIMKgg9K3/RE/8PkR+E6Ba4DAhAr7LDsL6TisAMbp
Dm3lRzbbKApeKAYb/h3oupkFNhL4MIETwCyVmLFj/BP11e28xKJ58M2tn2Nsid8U
zI/rT56Sn6R4qOhncBpcWj9JsJwgRnt+FgiJ7byAm9szBBsxrj5eaqyr4P4iEsFe
fLu9htLcdYInnxM2CpOpXrsNtPPGoi8OL5gjq0uhEb0G+WbcZ5ZCYnb+o37Vxz63
0miMTl3TMcmqD8mC0PWfEgbl+9vrQlAhDcNgxtWhGs99fSjhjzq3C5zftRrrvr1q
CgBwq28NOwcUuqOMU6Lw/XrwIpJUcyuce2zd/bqebA5StMnJxbLZ4Dn5Ce6QvdBx
HL7slIiLc5DpTYg/DnYeD7X5MDv+cwtDd72iIrW3uqS+QnO0YWf/QsF4L4z89X3x
iwTqXvBAks+5eHlQjMuNk8H2k8jdBoSRR+lxNv6q4hqp2UQaWDII69HNXLwyEoYH
9wB5SKfcvau4+jirSPXMtD/2+KLFlHpBZaIJQ+0ChO7vU/l5L63nzt7zWiz8+qXm
tWYewcaON8lX622KIcm1fnAli3qk+r7taOd9j74mWO0TVvIsuJs0u98oSPYBKg4t
zXkZai5qnF4G3O6lvkpUqRTAOowt0mljg5NFPAEvIc8vyxo2MCn0I8KuKm2vfetF
N0lkyRr83zylbC8AQxwIxC1AV57OvLNAWL4TNSIu7zEPcAirAUD3glpBS4+HEI4h
vHlRb4CPOsHaGjJuXLlZv/Rq/7SPHBr4LHRVnQN4jUSkiXbF1O2bqQcnqX5aKCA2
oR43pCYIquQXzcLx9kIonrCLd9xCAS6DmrrpZVilgXdYDvSjpVZn2mZfYXPiXgNm
j3YpIIrY6CKC/OeSTJkA+YQlB+usAFULFK2bi0sP8SBKdnwrtYTk6GPRjeamYNOF
xinvJbUGsO6oBCeb0TjMb1tey/MbjKgZhs6m5gA9nvNoKjlmMaZUubsK2F8NfU3v
WNFexDtl4/j+wFvlXLkoADcy5/09qTLohcmEzPF+KJeALNDVCDdKqMUvaSvjcHL6
ApXhtOPdsNRZKgkbR5qh/EwF5V3NtuIukHc1tCJ6S+sTIbLO8RgKiSvWCJJLM2A9
t4EfKdNiK5bUiUUhoWvEwspms9Uyl/lsbw6RBpZXD3LACHqDVu5Dj4GpYkpKnGBO
EIHESg1K4iOABs6lw7870obZd7whbC+sEDd+tJpMEtozTJDcNl1V8UDOvilR8z8E
SMA1HtQTwv3ojceMANf0p2nz5fPHeK4diS4PJMdkItgkEnKNrtzF8Ebi2Ybey4tE
IljNybSBVv8qZGVD1w1lO5iJYXUC7gVzisSJYQNsH75o/sJ6Q7AvJerWlEPZajMV
pZPlGXi4hUuRfCoqUgUxA3iXURpoyro+xUuda/2BTUVgXKtwJbFjxeCYo2cQYfhJ
/4SGwagI7I0ahR1VlxSdJQSQeaLhqNRcy+PsIZtkWS7jcaDwnmyIRv02MHQDd3LB
za0F/nj8haRJxlr6Ksl1XnTkBbIkFoXJxgm4fSPD7Y0z0bcZQfwGC+nbNw2CN+T2
XwnEXAaKFg8fyRN5TKyvsyFHW8IJx/N8zar4Rmdo9IttrFUy20c4sEgzHVlGA+tI
sY4bO06VsoWOI69xb93wDnCfTWfxb4K6Xknf9k4kgyiVnwQ9WZFGPsGfBfXPSfIy
mtj3QN7OobC2FlbxfCt/yEUhyoEuwRhTWFZDvshkgzGvxm2Ec5avX6sEOXjrk4so
3f+7sjYYE8w8WLEu1FyNo+pTGjN+FPDc9JGsSncctm3Rjcd3mg1iM6IFLiEYYu0l
cH3BWOvGiAYv8poMVqt08i3nA5ouUtQxe5KkOaVAlglGXfaE5kTcYD2xjHnjHJH5
K9ju+/Q9Lw9OH+JwKfak3GP5ygpC/tjT657I0WwMHksYTsiLm7j+TTXbzgodjQVU
y3O910Axf0Ai/u5TfJYI/h90gdSqMPStDPbIg2vmQOLCNI4oxvN1nkbks3T7Y9iI
7oTEG91uEUOnjiIAJiTH/N5DvLvPDpLwncd6vZoOCoKfABQIG2/ZHKhAoMacvoM2
3TAGgJG4VZ/7rYZxj5k79saqrYvG0+4A8FRtft1N6fI8ISeJ+lnYQY3DPdh7/gG4
epBgg4m41XUnJmwis/rJ1KR0lkvasj718osWlxi6DyQHlyfpeVGxmc0haXda1aVH
YwtYl33cb5FmHcIrZ8todqedmItY43I1JQtOEDRncfjfJS/AlH7r49eZQKJOHAC0
4FqO/alhswFNKBAkddtSiu3eTs9QskK1+Wsb2mpQs0C1K+qZJLoyW+CsBI2no3KL
AjcMHkcfVz3p4kJxR7eTM1/H0jdDNbBw8NmpFBEJwH3kSsJyBxSksYcS3v06ELA2
sg58FKtpHycWjpnudehVwvvnX7C4IUjDaoOLYacLjwoWqo1cRE4spU+0csIceKAS
1mRqNIa8SWa6DNM2eEgSJgskWta0qWGe9qD0laASs8nhEJ+JnDgWcCaLuQA6IixO
R4EmOPqZXk0e5g7e6fSeZ8gQ0QlX1bIhrftRpiOV852Xc04N9gtMMjpo9Jbnw3pU
Ir45BqOMnU1Jju6gQ9sHATYtrK4JWGDBg2bez534nVs37RhM650IXDJQb37MET0j
fsmmTOLKu1IAPgs2H/WxzAAEragAYEUc56wDQJgroneCXFnnSi0Tt9JIthZGkxBp
XlgWQPwCGOBjRpsvomx8XEoWTqAex8sN8/hgGAAvbGRlPQlXNwPvmY1atSEHsePf
RqXVIgYGUWYRyIctVXk7cgGVzjg0h1/J1lRB4vZq7LGJ3xzTJ/0igZSZ3mv7HszM
TbO6eiCO133EgHu1oXdiKFpdIGfRuz9JwyTTe8d88UcHtgKLJna2b6tORsRkASwX
TW1Mxkkw+k2XD5hvlxVbe4dcofSXMRfZdvUTr8XNuHHO8fgJaTv4e9Y6wqAAxd36
yDs4Oc/oV1xLIfqtCP+Qs53gA8JaLLgE0dt27MUkAFszeG4xk3x+6LvMB5faLQYm
ryjSYoON5b8ne06Ocj304AEHLy2hwuERtNQTs/iAI8S4PvZcEcK79IVw/bPrYaEv
QMC23Wce0vtsDJfDFq4DOfuE7YtaxQSWmkfdjT0OHlMTqGRW+mPcnNxM1UkxqaWC
Y3tHg9DORvvGxHdGu64h4eLV/14lj5db/MulkZh6uxZD6dQzmN3BZ1Rl+YKLcZBH
roUtV5pgmZeQZp7pzrldZ/SxL8ePGck3ftYLE1/J+9k3EhP9esLGz13ntbJevgIl
aCI+cgu/fZAbyKEC81sSbxxnYirdRUQV41czXQyh9sH1l/BBfWirlejeaxDU+355
a34odNiLNyGPE3Yfe89hHf/a8pxfeby4IMz4z1Hfd39BjUHAEiv/9IHTdIcqU7u8
YPf3SXdLxv2jeFVHHLe+7A5TAUoHBlt1UZu3L4RdJek6whmiF4d7VwHEZw9PyvMS
TR8FdG9gF9nS4ctDGb/KdL4vKfWxKtHvrcI7F87u8sJkFK8nFjhAHncLFTdAEbAX
xYqYiJLkhUBh++spdlse+2RlP9KzLhsbql4og7Qa1VvcjbDuWQ3AodH22WOabAk4
3uqhWpgBqY6quf3Vu+By4xGQSBc5IPPf0EM1z4HPT2dBmWun186XMcyBk8kG2KL6
crsKHNRMG5SY8FT+Nlj9x/SiqDW0c4joa8XqZyd2/O8le+uaVLmMEzkzol3NJqAi
ZTmGbKldVkmr45NSCUO+3QiP1FyXbXBe89v91fLXiW4OfIly8SqsyQ2FoASRkAL9
VarBb9IRKz4OsjxP6AkfLk4+dGcUfT5ZGFgbqe25esyXPT28yKvzEiYGQxScPIGq
Pij0yrPFuelhtruzArn6TtnTvasGM5YzGmzxs0UqGVVLWkf02+eKBockpSsACVH8
mK8d+09FpBjrwXiGqEl+T4mKvnZ764tSgSh1GdGjY/Y1mTcOFb4fwlxchJHOMzgD
7MYU39O56awNxj9TFuH3BjGNJq3fs7ITuvZofu3iExrLXlqm09q0Zie4od3RtnS6
rKtZ3jJ6+kbR9bvZVIDn88BIALPQKTjG3+0rbz+OQqojAafOzbyHF4YG9f+EeVkt
GkaHT0EESxZa90SijliqNuC611ePnCu/zSwoKku14/Kt5H+OLayzqeKtUhMxH/lP
nraPuQtJb0orhdA6uAkEyZH+bQjWRPmj6c0aUTnWCTetzWtL6H3Awq44CZXhDzJu
CLPhda91C1+/3kwGXfeSmfj47hYTGa1Pdj4Kkh4UPNiJOQ24XNOAGhtjsARUfQsG
VcEtdiSwG0NfR1zLqylas2s+df+Fq6H0eddXud7ujKm9QI/Ri1rR9nBgGCEEqwwC
ctmsq8KnSHjGGV2f3uGSMJaEdT4fPY9gpI5YxSXlWo4jGKetMF0RtsT6nInNlFZS
WHl9HKHPGyl/rNNDo6VdG4C0vMFswyrp3cthOZFcaQqJQPFhUkGpm2+v8kZtYfrm
YeoZHgFs2PBM/0AZsFhC6bC8XkJj0yHykBc3Krbjh29N1xU6/LYRv1JEVHsXoy6T
oBs96hhq26cn4C+/BZJXwrnKdPqGGyx1biVTLX71o4omKNAPjDvie07auQketk08
hnjKupS7Uck9XrWmWvOjgGG4I82kg5TGpFAKUxLy0U0rktqUFfUDRCrwG0dSVFlt
C/6osYtz1hY+TYLkqN0Z5ps4M1MUXuwlIvnwz1702hw+DgUxkgszBmj5j7HPr4jo
Q9LSOud+n1e5BhBy7exPMXc3WtF+2FblWiH/wVZ6RoSaGko6+Y3ccCl71hHau8X7
e4Kptabk3IexOeSIidBytt9LwFg0qk5qPDqtvKG8WqKiKfws4ltmvKPM0OlJWIms
TDv+1x4VBstdF82PWtzpl6ZxOIUd7iAreDn2PIukImIgCNgeTgjE69RUJt6tkzf8
dfsOwVOGI4qDOmQ4x9uukIncqZtmFpY3+qdtd7kyT7jvz6W+VGoPkW3+gCbiyYgo
zgCRRPJBULDl8x9DXrz0e0yUEfl86a67b56W6z6jQQdbVYKzf5BTLR2fSlzKy9NT
w8vVroju8p3rms7HNaDrFtVvuW2DWv0LYUIGlZhEF1yIny0aUUIAyCz1Ap/d4Q+M
uyH/5cU3mWlotIzWgu8WWnzI2Hpw8MXI8rONTATviTZw6DrRz+CUt+r3cSyITh3k
9IIL2+Dup+ZHoVOWAEB5rbi8cAkBYuEX/DXJNmimmur+bG5GW3bNLrQiyull7DpR
1+GEt/ii8u6vvzsBElENOrSQuTZpUO6l0MK42/+rhr6Q7ZBZL17gFIb/XJbC1MyB
kA83+Dl/OtqD8PTs1fzYjh5fwyqcd1iHFiG8xYXT4h6bmmcfuriim0LYtfIbLPAd
NLGwr+lOmzZq4715b/Fdr4kY4GvN/5rVBGjGTvBgHUCbvaW/XVuS3P3Fa+TG8k6t
UxIgqgxd/frmqfIXuz2L4oc3+DsXURE0OUXcbXGgKstMIu5Zm/5K6prZsKjvly4x
D//PAo1TaTDA0njQMZOGprALKvX2aNdg/VraCK/A4ZrF/Rc0D9fsI372XfiH7KUL
k87I4ugCod0c8DztzpjyIiE8+A+8tNU08GHTlDYklJAcjky2tlCZVp1E6dsuAH0D
/pkJkfnpbY9Bz7JNaoIcR+udnr+WtKTnk1iYt3rKyBD8bSab18tWxOLvls686f1E
Dr53ILmxEGCw+CekTzO8UKZygm/vzTYPL8ckxIaklqRyh9N89Dz+RQ1kea4DyLIm
NPTNsPg6cnDjSUQnsmQw7op2XC8lAdvmv+2RFLIypIsLkrpbbVpqgi+40HU248QO
VvBMCylx/AaKTeD7qt2m/U56bkDA1ZJU/E2SxFV+0L5cIwIuLvClwoumVNQf2m5X
in/y2HReoPl6/oCPQip7WmX7vemSzm35Ivpnf/WIMEYLqRDIIE6+g4zrKkSeSEBQ
43RlowXRcVi4eDbc6qvzv4alT8fhlf5VrfRTWrCVUwD2BI0aowRgVOb0BA682Idg
pC2lQFrkl8ok0ZXedRPWXmxMpb8cu8WoTReGtCWtXopzZcn/wqedJCgA9ONc213m
DBugOvM6pfKPePD2djTvif5Cui5cRtBf4gvk+CZ6YnbQ/cJvyg6k9Dij1GMDdDMd
CryqWFdb5MQ2aRTHg1RfGmwLKlKLw116o7g6mVIiZ2E3YQxGhfSlldAvA0UqDSHj
34av+tzjkW6Un+ql9w6oOBZj25k9unWea9zrU581v+l8YS2j/IBKzTSVGKgjKLIq
8KR4LojMimHTIMRJ4WXNDVPej2kQeL6llIgVRJ0MdDLzgv8TzVLtU9Bf0BCYO3qZ
y+8LiZIJiagSjwoCiaLgpH+INgjfbC17Tse5ivKD1775A32fzVlTJzI8Rb6uMEoz
Li2KQymHPZAPXXd5EGDdasM7KtegLPu1mzdWFC5A+PKR3No8wZaxXEvXKPc6aqhH
p2sIp0Z4y7t+VED2wHtOIkzMkEWiXabqQAX8bhgaQGwVWdcbTo41UDqHuqJ+GjdL
aN56ChlsnGQnGK4k5i8CyxBUnKL40Lr2MBVW2YbirVJDjG6VOv/s/VBNS13w3pYD
O3R+qG7ES1S00aUEs7cWEA/EwOj7Xu8st++KYDK74CilKgHFzxjHxDxb33kqjwhy
8tfUX4i+vqxZEy2UWNY1ZuuXM8RF/HpE2OZUiqQDgK+gQ2txJmbf1/zuWQKKDJNe
A3FgyWawxsRxScgle3j3BgG3OAy5/k0VPMuVKUHJpKENTDmR6EZ2eifeT9oWyRWZ
hXj/zOvRdYYjcuVAZVNrNl+uzza2PnSXi6K4vySSu+d8iPNLQ76+Up0QfBY3K1xB
cF8oLL3gDXNNOj8vvzuvQHCo/dKaRcSwBvR/5CWEhFJ0Y1iD39lVlnloG4CGF7MG
AfYM+gVxle2rMtuh0DQTILgxQBqNse3nLB2yLLQnpA+yzTewhSYLfDRAYpAhCMJt
X52KiYFxeQCWcoqxwNTWzXoknL2VP9NUu8dG3NDE3xjXgXiKi+ohA2Dn54/pQ+hk
GfBMIhCjqH5xX+n2hZom5H14a+gIwRPnngWaLdloHh4bUdZLEclKiKvLv2/YqfPU
bZ1nF06arRBZ5W+3NGDXni1kxhdGJPJJGk4knLh6Vq31T1t2detRbqVgr2lC7jXW
SOQeRQxzpl4nq5sRp2sj7XEsRCWivyAXcvqTZe38tPqkas9iV3q039MD9Ew6pG6s
VdL32ydnR0u+GVlCEzJju7d+VLotnhT4HfIBfHBGcrY75ugdAWbEarCyhYsZRkrt
7Y1l+CcN57E0X92KNC/fXWOvbTc4snhsCj7IOBl9FKmrtnpOkZ7WiEH9zMiJXJ8x
ZCf6yKAlY3sK5ha81F/bLI8l4YYzMSQWFVaQkSsbXWDoJSRENecTYHn79mRmNYsT
j4jFfiuc8xpQcPK8Sxnq5G2hx3wRqcvmzyv3gd5vyMblmUQGbVKSw9eWqYUURPIX
S0+/fMRT49qq8fEgYlrefcYUeSa1vwONezfTXtcnJCYI9tQ0IB9eRmn52fRM1h+/
jsqKRcsDHy4PY3Imk3aqYItYqz4fL3mf5xTFi4Kd9w3zF7mtcxIEXxK16BBhnvuZ
leeazPyStSy7WDcB7noR3y0gY9RDmbxsk2Bz6kdBQlLlbpoCl06+9mm3vVT94uBt
9tscLVB1ZWW2yyPzV+4lx7BVhyAtk2fu8sOfFkKSkS1/RNWdkQsF6/JgnH5e6QIm
CwWNP27OePsvSFGN07tKbj2cyUm6YSeJVeLiwOgFONnQI2GlcjlL+OomiAYOMZlb
O0PU3p3hDCvY2tmsx8hOjxgxPFUCHRL/QubAD6Q5eJu2EA6SOObjs/cWyjZZlQYw
gG9zzR/o3kRgUBRzus/1IEmspqoVI+4uT13WyO9jjrmeIK01uGGlnWzwzV096d5R
moayOc7d1+lykHUxL1vDB3bWOA3mOnlA+8NMWwdSwt9HYKbyj1RpswIGgPirauXR
wCUNk+rr0Cev853FO1hNk01dHBX+Y8SYa3RNVWu0/iuMZt91sxsphpSMH9g5PKx+
CDz42ROYoZoqGGC8NswyoIAEiwXvKYiCeA3haTq6V2JYyG7CVi+ldOUcgMxDv0ts
XUQvCsYxQw1bGCUBc7yhDmcEgFEalpXSzFyN0n0kmrWtHge+e9JzYCj7qZ2TfBKs
A1mrB8a1veoyQp0MDT4GlP+TWPdEgDPERPq5Myh7315LIh2DHXPHoD93uKXsxGR2
zdJTUdmoGT6SNt8MmEO/DWdvEATtj3E/HCm66XQ6GiP4V0axzZgFPel0/a7rdwrk
ExrMEoUiHrQQVleINMpzKMkFReEyEl/gqhKxIeMdjh32FAdndvYYXonpo4VwOzbO
OBssv9PRGHu/NposENxG0FY9U/2s7+bRVkqnmfhUMjWQLmSjv4bHc8uj5TBD4bLZ
qs429UGjLgkDOeDmJmdbk8UStpWcnlM45gNIjXJKDwjI7xYcA1IF3SEbW0qsm6Jo
832s5fB9Xc3PLPHqoqjwDQMamdnPBaeKNeP4GSeDYQIl3s1kgua1ZTomaiO0d6y+
LBuqCx6Cva4yEFCcdsbS6eqEpUEJrsvdGM1EvUsMd777dyGOW6Y1cnBPecSoi+FL
FktM10OmVs8tvQDREpqBZaGPb8/1KOlmlPLyloEauL49bV+dvSRx3CJ0F2tlkGCO
S5YCkud56A9BzCjcFg4m7Iqqejt6OMthhemh9WiWIhwc7bAADDnCMFYuMfttcPIT
Ag83zIwPICO5uFiI92399f8BkBNu0kiJegngkVsCT1aWFCvzfVYah86FlKULQl1O
N542f6nB8zh6QThGgahQ6IkQIvjsG37BLS2W+V3r1yek3j9Xbr+uC0aHJpNcztwy
dwRZsBuLNjQqu3z3aUmFDt4nnqP5auCTF4ea3Am/D5OD5FZfQtoi13aYhbPmYOQ7
i4sGbcYgOJIVfUtlckyTqd5H2WruoHJgFZvfMpJMOE9VhdmcJMtt5QBx7d3J3gpM
2RrehF2vETKoiCzb0LMqZZXRoTB32O+ciYLyCDR9V3ZWC8yuTfy80xYH84Pj6WWE
yKgMFRBepNItyt/oeu8mzBPPTS8L27ZeaAkvovKOnOLlxLkS9/GftuSs1WZQAXHi
d9TMeFbCHM6cgBuxWnDWv97hWyjqULuDDSyKP1XQGuPXS2zrSASU/GbtCKRWxsl1
nXYS/XSPlpfDBRupipvAklpHLWviXB8ukTppsQyDWZamGQmIygltMnwFiO5i+DZw
07hmAt+R6y7i6342gad7s4ImuZoGo5wAmJYrUcddxCDEJx8JjL7BqBLKHPav7JxL
17rhRZIRD5DCUB4OX7a3VTWkQnrsf5MUp5o3gflQGMfU3WJCBKeOnuSCJbPrxg62
t/I/ErcDSTKLnLkhX0hGD3eqzaPWgzjVCjJjMdnqyI6BFLcCHDhtSt9M8Kz0i2Ox
4HRuGK1PAVJpKnT83m3isVPgTmX9XLvb5XkV+64Z3V/8xCM/S553WnJ1g9T57tWB
7HCQe9uzUeRvD8mirFSUPSA53xKG40AvcwwjwMTQJqDAwfwudpItBDxLiD5WRFED
Xef2lZNRTFD2XaEZPBSJ/lPhd1c9hb4HF4EmEVcG67q7dDsDY4WfV/9blkfcmtqJ
+okEJH5KMFOQI3H1XWgstIq6OqB4BGMGSCqr5bAMqD1VfjISm0s01FEum0FhmWqm
IZPB2KZsW57VLBTyd5UZoq9zxwtx/S/BaEez6aJi/DweOpC923FKN9wpxbolclVK
WQPLWXnX8Y3LKo0qawpEpyoJFsJAG3oQSf0uQDHu8DO1d3dq9nQuReH8i/CMZR25
j0bEN5avqmb7xghUBTeHpK60iFWR0BBeI+/ahrDHcXlPmH0sGnIM9tb4o4ga+ntM
Ey94BCZzrFsBvsaC5x4wXQ/NX1qlTLm1wPyPiiplCyo2K7ELEryCD/k3j3L8QYBA
ksKo2WTDx/dX57b9mTA84fuNW6kuphbSsmlO9gHuqYGnLvT1X4gydou5yz5Lh0wf
tsN0BWiRp+CJ/EyeAuIiqYTrsx7Dmdu/Sv3EriTRh7h5z9YxdwKPVm/3lrDj9ELl
QmVbErWmwJF0Jjg+ujjgd4vz1yLhfP5N874tCtCdcBgr82I9jqc32StrLMlHvSLr
hZ6DuQGbHwQyqGyGjndg2Smv1wmeufpCkDaVXkfoJUVJ/PBrxmwTrdRCuBaMR90A
tK1oTx7V4lAwTnvKyC80t17U0VL+JIp/BVcnXqGtFE6Zv0ntsV2j1lxIvxZx33ZX
w5Jj4mlbS9UdFe9hPAP+n4gbQj+zu3UMbj4tfZfLpYUXff1rpIlJICyXk2DP1dQC
BGpwndusvxdkw6pdrtIn0rCkrbGrIkq1Je3u0llzH+F8O/iwjWcAF6W1x07G/Sz1
vY7rtBA/1AVysPZWKvF4LDIdSsLEEeEXsKjSIxmA13yHh1xcB8QlGH8hol/S9I1p
JAO5qne8lHePStL/arU/FxJpIOOSXeOQAQqDiyUqtH0SLCSaPLLRXE1zGDadRqVs
kUT1PUNZgnquCaAGWLZYgj3bAo8o0tOqOpaSQY5kiEulpcXxT0RzdSS+EqMo5YV9
rAAWEqyq8wJG9PnNj0qKfbLhKus/6gYm5XBKuDBs/tCFNvpnDGKVAPtOcH9VXO2f
gRKOp99+OCsGoXyK3hzl7IkLLYiGJe7yAvt6cJJo7whm0MYUCV3zY/V2P6ahNkL7
cm9cdoUPyX+ZWQeDA5VtBv1KZBLHf7+lrr3dmJeb5oGlbr3UPnu0PW6OBJqWCuAq
5otzXUx4GFdlVEomPa+RMMFQ19OnhmgYTAn/VmPV/6J6fHFBZ4U7hhGyTCI72k+s
CMxajoviOIyxy85tDtzSjX8YUKbJMuJVCuHY4jz518nji+3eI9DxLlX9cqwUq5e5
JhQR+DVIsck1GIB//YTox9VQr9CcvX3taBCz0ms2j8N7fjsQxMy7CYhdFSugOosP
SB5AFBNAr+wzQ8ZqBU857gn8rSSaeYYFM2hR4AybGvfhlQGDfgrLzR3HMmNDOwlW
22YWWde6ToAN/HPBMgvU+70qKpeY3j9KB3jLjkV+eEmUn5o6V89T+HprwTTH/RKr
wDLKAVF5u+/yWJFqCxyhGtZ5ww8+Ut1uswUYIbAqNVq94HYlHXWH3W43kSLDI5jO
ov9l/G8v00MvNLbcCyW/1y0tvRrQ20P1feGfnMX5/Riv4Eu6MdvzWxZMZztqlYsE
cOHYzL0HSSFKv+2CErV9/q2TIHUG8lQBBwYFblPcFl2mTeU4GH4BwF2wBWMxPMgY
X3YR8PdpePszXL9vSBn2ub2+9M/0DKVnXuztuPOW9SPEk447DTzJ0/4nv2tyrsz4
4PZ0OkIEJOOPqNFXLH7dSp40O4xdC338po25q6mhPfVUjwqhQwGAOSiXmozwGCwy
tLiej3NeySQ5r1KXrKYp9gN+wjQ2irAEkfa7LdUdd2Y5/Hfza0pgxTmlzD/hGGT/
P1VJRe5IGJi9U9yzSaT13o7gO/5yVliSKLwUE6L2um5BTiMiQXwkjlpZIRF2otyn
lTPx/kk1GZftMhgYiDuz85OKODBsiN2Sx86+HwS2moA0o2m60t9tXyQefxqTqSFH
2sY/wqFXuNgdgT4yjXCEBs6/TwbSNc2IH0vzB1gfEBnEOt1LMTrV+Md7DU96aAo8
zq+WDCK1nc6kYyodNQhfpRcVySfjrwzjq74b0ByhW4I6nudYt4ZFB3CJkfCKo+AJ
C7q3oOaNkB8JHm2dCwsB/xK0h1e1IjcmN378gm59bwTkk1opKhpqHc8pc3+fxVrz
lTScPHeMkXc5b4hYFX8jUYslWm/SYjv2CmfYMCTqyd9tD5DvftOVMLMQqCv+AHLP
BIfpPMQxoCb9Ci1QVJcc6XfkBaDTMIAJa1TkJgUeb6tpyD1rfv1p8AEIi9QYH5Lz
6hfO8fjicPye0S1lr5mp29mYYclZ6QyUPfsFGGPpms+9uz6mTRLa8FHSCUpFWKJ/
K5zsVVQraaBLYRNac2StX7sML9LO0ldCz2wSyZC3Yin76AkW63fkboVEqlKsNL7e
LunD3gbiwM2r7cBososumTJy4l2lqk4qGb2QMwVWlGVRo924EeImI7Wiy/dcqC/Z
+LcPgwMQj6odu7cm0IoH0WWDgQYsW2pUSmsi1x6HdItpgjki7PeGdmuizJUtfCCu
kP2DR5Lld7Ln5L9FFWm0yEjhwXAcSYQorq3AODDMWtdQXGIyt9W449kAVqA9HQFb
+BAjFJITLvVz6PaNUt3ZYq6dMiDpM4BecFheLBPVJG9CF8hpWS5F+4xzqzH1CqGH
BUX9nLgYQcb2GwGUU7+ZZ3ph628xCoj/fDaQl3OJAksP7y6d1KYc52YRV0ECSy0m
UgtMk4n8PbNoYQmquprFaS/UGDRXUUI2NnJYlVWGs+enMvgJj0SMNHkwn800DcCO
4a1L7Athv5dcZfyCtoV76CwPX9ndxY/DaiOe5888caLGl6Ho9ODFlYuh0M9Dux+P
Ko5BoqdnzrvwrLLJS5do8WTYPMaJHMOK5IGFOgmxsy/tJjbY9kpKEqFTgIX3TMXP
9cJw5rG7cHd6rsywJ/65ZSjMEA1cuKpkVv8/kgusrUqpQhgHeOGULw9mRU2zvzHw
aGNdpn7PlPWDZGNZ5YtKgqmyQLCGJjqDp1+rLDiSMOCPyfrSyarDAT/jzhCKFVZG
J2ur/LsfudfrBCQ0u2rshBil57hx9tGS77U5lfHTWoGrKpkFvKZGzWcspG5Raidu
m1thCzUSIrz8cTnKwN0ljxmjaYQSBKhmQLjqa2a4Bhy6spB+iwwXrKlIflfwJh4U
KRexwT8gYSFflKsqIYxe8HLXScvdy1AQ+c6PPHZ8j7nmCVmJ+AeH0ntJ30hesNW2
krA2J/i2EMespPKPqoacpE4aUpyDagxpIqCJaUA3DriEnpQ4a+q2sXNlGcIOtP3V
`pragma protect end_protected
