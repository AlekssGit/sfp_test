// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.

`pragma protect begin_protected
`pragma protect version=1
`pragma protect encrypt_agent="VCS"
`pragma protect encrypt_agent_info="J-2014.12-SP1 Build Date Feb 26 2015 20:50:25"
`pragma protect author="IP Provider"
`pragma protect key_keyowner="Synopsys"
`pragma protect key_keyname="SNPS-VCS-RSA-1"
`pragma protect key_method="rsa"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 128 )
`pragma protect key_block
CEDevu0B/hebfO4dKE2QC5alpPHjaR82PTROg2ltEHa37kDXeRUkmE/CLXxZACYX
RRzBd0UPaOhQyBRd7MCX0fymKNR7DC9XRonof9eB4a8wGlY8QO/tAoNEBySzIkvZ
luosf9wI1e5jDRLJMoABP8Y4Wgby4yv/Eg81tKqZaTM=

`pragma protect data_method="aes128-cbc"
`pragma protect encoding = (enctype = "base64", line_length = 76, bytes = 5280 )
`pragma protect data_block
tKQI12kPlb+1FcUcjUTaoYSTsvRbYfBNtZ+wPaSI43UuiiUHp/C0PRqvvYTCfq8v
tVBQf/30vc9I6wNN7Ujrk52Onx4eKfynWB+2Q25Y7ArdXWkmn45KxI5+h6zhtF9v
xIPqCNqSHPjSBKMHbj4r/ByfJa4605pUZnhXn+zez26O17r1f5afh1nINMYl9adV
h/K91nftaBra/FTtnA91mNW5d/PebFWAP4kfIivyyQhWfuAgLgAdvwLagbyOoAJ0
GjHYnlWG3Mt2cokRGtU6AWFgx+qGXYYlgWR/Je+f5m5oWEi0B/Adi9PqDaUeCHfN
CruI0ynH9Z2UJL+88W+Y+qjiAHXHZKb0SHMk3ORN2n/WQIYYz/NEYKfoWw6iEy2t
ON889EpgEpzs5N12XAHEGI59QSZ4k7bFNT23jnxxTTdAgVi6a+JEwZ9WzYSbI6oe
LXRDrX5PIT6YXM1Odawsw6uBBKl8wUBEaw2ELJIijPssGbB7HxPYJJtTIcwncf1l
yGz3S/+rtf8ww2d7ov+LdzetX+MZBCAgudUk3I0kNQJCwaaZrnSH9QsrXOEytfjH
ksmm22BeausxCK5oggUmiKgNZVHSdFNdpsQ1UaI4f0Vskbh+YACzVUHMyKp/3uQZ
7Qkc3Cp4SsyIZX2t/6n+u4JpIP42hwo7LE6QqJIpnBbp4ZYHHfvS6ivQVvCB9Tbk
7i/NOOE4Vxt7SBZCPZqEljmSi7vMYPA8S6fPNdkmY/oATQ3okEo6w7r35J9JXyM+
0zJFAMDJf+oX+O8ajYjApdmtFWh1pDx1csfbpIBwrovkIp+KHHxK9l67y41TNs1R
4L/+RMwEgmMs2+r3M4knqvL6007daa34nreMp97wE3QSbXTJVHM2HB5plEJ+ez+s
Q7jlRGNBIgfPAAUF71uuKG5Yx41+sIv/nH20cZ6dUgqBKS76438PupEP+D/ZGNin
XTnkTqvv0Tt1MU7EPg3A1R6Nhp7lhAfIHh5q/mtdTtOse4zDlia6z+LQ9y5ln/A7
z7fCBOnw7IJo3OX1RUPbrCzj8jCRNTloJbnfmWUjJV+d3WOYWip1dJi9zVB7QFlE
nEChYC1CSopN+G5rrn+vMa1eJNmrDKBxm3/Y3B6DU+Q0CifGCZeBvQu8ga8/DQBL
AsELvnBE2AOMD4Pg7GDz0qKj1k9mDN+n0QzuVGU7pRZ259JexPeXglbRwVJStZ6P
t6VbfXG3V+YqVWECSw2Ow6Mr0CGvXnh/vhqjfE4Lm/jrA0gL90w+rqRktt1eYPMH
Tmd5VmaVH9JZptegd12k7n6Ce2dk0Qv73Wu/zdLrFvP+hJbt54KBdUY/mfs9wx79
cx1HN441AqCSF6OXHPU4u0ypAj0J2nlkf2GeMN4xVToLwRwEwt2mDDuilUoVC4qJ
hT4zFlk7p8X+XjN3K8QW7UToGzyMGai8Mf/zay6S90UWJJCXI4mdXasi8BP1YQsP
tdqAQpz2ulCbfLkrVqPDRBagksxV55rpayNLGuWvrkw7NAQZE3j6jDt3WGqfm4Cw
47x+N34KbARa0knsFR10P97KIG2JrN80eG4s3/9iIn96BbdW/pZUQ/yISGxNh2aJ
IbsvSa/LE26xwmuJ1yReNwcjbv3cA4VSziKQhFMoFkKyT530GfaXqOWpRvZL47PA
EgkuY81Jprd1kqtKvtU/KRAVWsn69pIB8xp/B4Cv/mrYLSMF+hwdIi7cxlOyrwi5
7SVFENIEYy5yR/ZwnUBCt0u8uS/XJDresSZkKTtIbbvMx2xhG3XgzUq5wpXVdcyw
F9FeOpxDvmwNde6WdbslrGCspDB1W7xoyiKEdh1L9wS9DaSw8tuQigcTzJ4fGW5d
0kisb3uRLVZSLcsHGtIN4LVhcJfxUR4eTsSu3K+Yt8y35/anWb2XntFNA6aRwIZu
L1Pev6aoPWtxAuOEblNgmwQCXWhhskQfzyIF3/zuW49UI7T8L3kgFTzf+qu8MOCb
Mt4Xp8gl22OhULhBljpXCxQG5Iv0gcdj2NAEEa/BZI5tqgWuf/QbybhN4M3Chlmj
EWK3Oq23lKuIPioewFdi527y4F0C0oxlmQQPgFWPh5SYWEm8DgVo4KYGwfZ8a5LC
uLxX5i5QggneS1zxRZudycBsclrJdBO5MiSWgnAeoYf8dvUOfS4LaaoBGYx+7PAu
hfu2i02yuWFiCaXH5Kykk+XV8tYxqsfMtmRkQBgP8ymuJHDg6CUFzh/VFzwR8e9x
5HZU9l0iIe7MhXt/+VLYUzVz2IWGvW9zAFx+YEGwGaymX++VOEwkuo+j415Y2lZ0
Xosun3p/UrLRGk0euFejbTxx2two626Qlt9U9zYy5VdMestpQjCpwAuQwO7wbsrT
FArVCQrGlKOodEiY/nHJHUi5sedxL0vCMbE60YDArYndqqjtDKwXrdhfxIYTtcfZ
24eUnBgkajR0ZrqKTPwVhu6HJOZNnxgE794H7G5n2vcIag63z0JFXa6WwzNBAReE
n0mX/m+KQDN6nDQjgJSDQL5H38w4+d5kReDBcXWN15Xj0tCQdxXZug47jEKYOsLr
lIui/34BWyy6DY7W5EAflIEPBUx4WfmVXMVAAI8JdhAJT1IS8SsG8JT4/h3ezBLQ
tVMSGx2v+zMJS6Ki5XvLkyLKdg8/26atfCJrFrElJWK6nbeSnvR5aHxzvxpbh2sL
xWOfh7IjF2hqtFy2gzc4LLGT86dOmE1RzGSZa8XGbE3B/J/EoffR56zKv9hbjtaa
F8hDqywflqZ5nNDppTz9U8sTS81fMqgHelzcVkhL5DKzMOd5UGsfW4i7iQjnfmy7
DJLLahq6KWBKJBzc3LNeZI+RN+b+hK8U7Dejf077h6nn6AyN+rSxoHO4gWbOJcYr
yKemdPGYL9sBt9LULqJzWHOrlwtT/5M6DAwTAEnVJQiFkd1cIpUZPqupBBgLe3lD
FiIgikIfNsaC4jONYx53JclfxP6lNZujpLq3RaFbZcPVCUBzHyvSUhrSIcgRD90R
RZ5MTV5RwKtVoNpIlQ+7X6rsV3Kq7hCWNmvDzolNLb0i3/NN+7HkxgqWb3rz+1h0
hyPr1GoIAUN51rsn8vqipJAjLmTIwfwyfvY4KHYyam6vwQbYjdlyek4vRUQZScnl
7Fxq5rltqnF4jEax/5Zjg3tJsfEKgfWLrMOLAgq1kqrYdxsyHPOQgaJKrWNTRcx2
EPImK6RJm9YQCBWv9xzkrvhjxR4gpRmJ3DhX2Gq3BHIooId2Q4oP8rRcxRb/tXIk
B0+AeniMkAEkPsK5eAtTeluAzex2huTafG1Vq2WkDzn/I8tfy6Qkcz1Hz4OlenIT
L1XQ8Jl7ivkXBLDZZ9+02bBqjFfJr5Ngyal1mhc87ObyTfAD646N23kXP6tUsBQf
Hksh50Qob6fGFkMga2bfmL+2M7P+fV7aSx5QFZEKhb3u7mrQK2mwK8K0l3jFfeZ0
SWba4xn5bdC3wk+Anjal/S/YlDcO5X4sQBpg/17O+0Z6eowNUQJv0g534opWuv/8
P/YsUNTuwTa8bOWw3DJEDCGnszJwcOq5bWK+b/2u5/w72E2RV9K0iJCRiiIS7gZX
pcC/JrWy+s5ldZA8UKyl3LQBXAXTRrwbUb4FFod9BVtFCMZbmQmKlVO15EqG6Hop
QCoNJ4cJw0d2aOYQeg/SkbfSn2RmJZqa3hhGFVrNQgIgZEI3DBj47orsWOlOhBuv
sXrGoWXvMM2L1YQ20n2NXyymkRMGB5VXOaixmuTfWwS0yJIcTxq7N5Flcr5tBQ8b
I00fLpVH5srS1R+J6gRK8v1cKnlhjzda1BC8ci2tonQBSKR69/PDy67XYhXUuUk9
R6irp4elvcdeugs2J0NcxxApFaJMJH+2V+nao3Z6AKUEG7mOK5sMPYcFbNPUVpM7
53ifwLOUvOUvy2JN5XGwBSvntAu6c2JNdwOE1WTRaUOPbpn/WXXNyQAyaSI3dwR4
HcFnTCsqF2YBS+thtIQgiuLVnEuSi5Ld+/TAOeIG1h/8A9TmgrNKQOWlOpT/RwG8
nC7OxK4PF1OJ1YoRrEDsmaw+VQp2Hztzji0OFDHG2oprCF0kwEGAjGHgsM48wA0m
UYSsadcBghveIGQYBGdG+UpGDBkNWFEijpxMm/ImeOikZgK4/sRaayA+ZhHNje05
TrTAMOH1wKRdGpooPNkPdlDkWma68UK/HCirNo3ilXVCcSfsRzAtlZeUp/3qdzbm
U9WZx568qJLaI5z5TVBI2qOjyigVp0JF3MQaP9pFojFVaOlr7SzkvUfV/Zf629iH
9Zrvl+E5DQ2hro23rVVp1uiLcncHxhV7Z/jXndOTq1RB2+ivQh4hEhtYQmgMv+7s
3D41JDanVbm0YdrFBAJ5dRhOtBPiDhXitdnZfouGuE+sBQiL0Ag0c56WqiQVRGpZ
HiKQRBfj9QeOn66V7lDrrSZG30YTwan7FnDcOD9Zp35oyqhZC5Pzza2NBVZKXLMZ
yVss5V8upMIMzo0xR6FhR4x8b10hN8J+5DaZJ6bg1kjTalV742EFkzgjp6rz4KlT
W3ODfgyeFZjKUYszQwoBUjjaryK08r2Zq/BOGbPXJAEi1cv4+uo4A5Vma0E8b1xr
5el9E/y+Ky1cJW3kZrgUxUT3fmgfdXtYsOQwKar9DNmrOr/1oTnaIUapSGoQoetT
Frr/BzMvaTR+gEN5lT/kEJRWLNZNnFQg4SWsXqh2muWz3lUt3vxNMjadJ6dptEG/
Md0pIUrjRglUwsBkG5F9825vul0ju4+pGRRPRwm7wBm6cW55Tica0F6E9sBUDcl0
S4Nw89L1zxDhvlS4mWFCR+D8QdO7dBF9KYPFsc+mTzQDcPrW7N0LKaYcRoMkoYJu
352+2qXv316T/H4Xn1Z7LE3HkHsQ5+hxNQa8Ju/LD9Tdq+yqIYoG4augi/+T4Sfz
gn1S/tMH0tV4oFxuRo9Lz3j4CI2kdEzR9gsDZQfKHsrLoQ8JBA7Q8y4DDWohhs+k
7sXaIs2j/Nq4wbLq/d4h815Lrj5d372Z7ckOsHs4fsyPeplRWTaPpOfSPTJBk5sI
dDFN+pdwXUFYSsUk3JZHxe8v4Yk9AESNd5bqkh2ROWNYc444IjGD8WLLpmfs42tR
2sMVNe53JN1mRTK0hok6EAv7dkMbW7im9zwFzyOlu99WcG44Y4et63n7NmE+J5Am
psqKcc4HfJ1qrl3HFf4rvVojJjg66JoNbAFTYtjEYZhBSSDNbkLancftFYvJMlOd
Mp92vfmV8CJsixTGthprUV8c8IapBVQVIct6hO3fCUytbVAspXzFweuK93U815BD
GbG8i16u8UPA8FBe2CwIp7bVL1StsJcRzMZxizbLZQrOTyaWj/w5fLxEMHFx/w+H
PxZObRmgjeGFVOhAtBgLRDjjdW2+5U43CF+xySEDMxzZdiLdCEahrWIIxXgMuAWK
k0txm6xulUzav+Qn9B4B4HUfcCb72G76Fnu+L/odoOK2zLiexdW9E4fN0u9zoBMs
mc40pJfYF502FCzJVsaRVm3ffMhxHVtsPTtvlUKisu89BeLlPaaK3rY75NoKJW+/
P3FiK+6VqB3HEAK+RrocGe+kMaMf2GxRxrItCAJiwHzKRLrsCrUhhI9H1ndKASSw
C9Rsu4tUepeXOo+nlWl4XBQycwPMIraahJz4szEFcexDhx0nh06p+med9UdN7Fo+
6NmciYoN/aiAFE1V4vgQWnqf6T9ogy4ZYUPuci5U1EiY7Q3amBrLKMpzDEAuSCPC
gpSaGHHz1d1JlMeEVBUyp8MG7hM12OW+fgdUwqXUpXvOIJ2sC1NwFcY8zS25UOMU
tvQyFSrPbgvKGPuO0FP+VoABf/rpGZRNWYuSEGmazdSn/f0cJ7GYvm0oHODvWIpU
XDqwKFAgX2zzcq02HFrJn7FdGoY3YLqAVe19VGUN0VdtJ1jhCMsR0jgUsnUh9LKm
Qsv4yu1Ww7vjQ9F2h384dYE1uQ+q0WIdRNhXiVgR55wXU2xi+2WHsjqtWHZ3rFCm
xquNBWjL0EwfJ7d2OjoFz5gCWpX6sobiif6eGqzniMF26IDFzPrLnMP6Thes0vUd
6yD+z7ENPEwe9jV0Rpe84XfkpauTdypfYoJRjrypRvOVPVSm/9D4IyrY8MstvxuV
dOa3tktqHsE4E0JeqFws6On5nNbo4s/oH+RwQSkkzhmRhZ9MjsjBYyWydzpsqvBI
Q5zl5KPODreAJ+fRCrn4Lbhm7TT/uWn3fS6qAG6ocGPGcgjxgFWFc5mO81IFLX+0
hwKJ7v2oX85asf3Yjb7K1V/f23GyaJ4ODXVNB0eXHPwho9Q3Tfp0wFY0gl15dtV8
zz0NlwmMIWVHEGQdK+nu5r/Pe/CNcE4XKQI9AUIg+5R3WehTc+RA+dNbsfBCXx6E
0wWNjvGPzRUL/kKBF0BPwzyAzer76H5OetnjiK2ZSFGom2TnqJ90KFPzYM+hV9Ca
no9fI9WXS7OCd2i6wRIlTZd43muENAnYSecLXpHoC1iau8TtdPEeA/rSqetB87U3
WZsHfcRFksquJoPw42anauj2Pc7kH9Y5xdYrHhEhrv4CN3Gt6Oks4d1rn41dX/li
sGXmegmzAaoCkT8t1On4Micr6ofz4YnNL2tdHzI2xrCgS3trOJc+w1jhiJQOOKdZ
J4HU2Wqs58biO6l6Fy3vMsz9JojGEUDMyf1SHAYtfSm4byy15GwaHIX96Nw2BFJR
Eapo1ML9WxFHMG5zZreK4ZzJO1q9B5dgdZcmr8GjG2mAFKJAaFlE4kfTxtg1KW8/
P0qbZUvuc5yh2TXvtWoDd2Z1HCzu6OsbmahcC2Ra8sP8qfGbo06mlnecnwsEg8FL
9rNconu7sdEdQplS9gyh2wS9wVmV7sYdif+yVQT4dnzqtiQytzDfxIgu8JuJOh+S
Q+Y7dYQ/5zP67FyziyA1zCKPfZVq5quFEQEBNgzYy65rggbTAb3B0SEfRrarQPc2
EWaNwvwJm2hC0vd+/b7V+6W/kAtGu99dp1oDeerklD7pC/eT6T8kaAEJV2r4aFK9

`pragma protect end_protected
