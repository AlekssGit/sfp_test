`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
jARUisgLYsXu4v5q0VEWY0u99HVxjgRlMq8pKCkWk/PRb1/CQhGXq73gbZnu7P9m
45hcYPE2Bq2wKoYFp1rz0gMh3LFufSkJEHaCo70BVVA/Vm6N9GLv9uxgAaNT8+kd
6AddHcjtZrSXgMwFnyb/X7bcZxzd+IW/6vDQFjq/O3k=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 5680), data_block
9VfhF9dcklObHDkGaq6av/nxv/sDtJR1GKbokJ/T2HbtNHajFAnvTPTkePI3pwp5
wmghYYmWEt2fj9C9SgUf0npvFtv6SYkh11cb8ByiBe9rV5/xA2UjfCeVKTHHKJj3
pfmHBdOmRvQ9yMIPKRZcnFVKCuFYOZLj2QV3FDmHQjvSL7YGRaNa2DEpVlwaWr8P
mnJTLouv5hTUpd7iZaPj+D5NRj1q7rrkFIy3ucinEEs90D+1cg8T0C1gUJT9fjfH
h/j1Pr+SSR3D9FVb2aVkdWhtambPEUr59YuTvY0rxAFY+a8pcu6mpiF31AiPrjSP
8pRQJZJQjk6RVNF54v0ThWOY0oDr/EaO+lGFGRL/2tOp0MFwxlNl6H7lqY4G0492
iMfw/YqzmFW94Aj2rckWcGzEfN9zTTxpn+Z4TvU28fhSc+tA16twL6advlCY1btC
ue7fPQnGdn1Nqoe6c71Lq3/jmhpAhYu102tr0GRoAUDEGXFkjScvS1Ok5D8yZsaN
+eKNRnDMO6ede73fJL9GxouqgzWvcsol6VSW5zU6nMe+mt11Mzn8QH7rPEluzi25
0Msge5JHsRz1nwLTrVq+oOyDOm9JlFO5R2jWGy7/m/amnjhsZpTo+bAlALavi7zf
DhsGhQNbDCfTjrY28gxeryQP9gZPykQWyUdRhM5QioW2aYuMGY1NB2K5FMpUo0gH
zLM8S49SdTrBn+R9KDuWOh1HxgZ8D5sMNFsUTaEs/2yLohg3OQpQ3br672sCIzrO
X9FBkzeC2XbnWvXihsVtdE8Bc0jngiIg5h5VMEE8TiHPciFqho3T5lVoqdXm9d29
SBdHq8jVHNJT0dPeVPueASHrS2GXUygXmMjLdfPfSEF61L5nWrZiTEa6c+Rq60u1
7q668NutTpMcVrzReAmpYcK/Kli8YUYbabqUUsJLmpITm0T02ktINuFJuamVZ2Kk
q3fRPag9F2ap6FSRX6OOobQOb/nELpuZsy70xK/sFNQOgwSF9jXnV1ft8B66ZClz
0gjrUrv2dxg6j18c6l8oBZzGP+xm9s//dr0Ptv+Ip8DtDUAuS+4jDhiZVwXSmNZL
KUb8oSCSnZ6RLFgFoQ3upkuEBnn3YJSeWKx29AAi7YQuzr45dGpSuHGH4E/ebBRt
npGHMZrT03MFLSuVgVgjwytcjedTAVAUIp72uaMAiFAkvgEO2ZzL7/aVlcTM/wSN
JoyfHMyXewB2/y2wZg10dSMbqSQesASv8zZ26EpBIGUO5hy4WUA0wetu3cbuzr+k
0h06gNOlyjTUFqJQP6cVNEXrUjR5ykDLLGKarJhS6q/bgwh7kjXnTsxRv8OIAc+s
1iO7tTId4UQQbIZPemVHp+yANyH3bX+RMLDBUdwoCRwGUw4cD5Y6lCFbpeyjyqyx
jw6o6erOzIzUMv60sib5qs+sNPNJWguzW8dqxOdUeOen1HNEbV0tDn11MYt2ZdiX
N7O48QEC2aEyQ93awgKp8kCJhxMFutOvpDsLD4yuC+kL1hHtzBfCyc/NDGYo9yee
B8LF1EkIOc6OSn4Y5sDUbIdrgIJZlkdXvRh+a8em2ukb+A35Rxzgb67n+iecFx25
Ezm4jB6OMQL0XdZVrw68xx0nQE9j4W10vO2owjk3qKEv24P2akG4PyY/flaj5FvJ
JJ2fPkJFxzzjjFThEblodueNOBQD3941yelyvez5uvXs/09IvpqpkomvK4Q3z4jC
gcYEMB393l4yYB8+dDBvls4CvvnPgP/LDZdxVLlOs1d2NjtDg8uYcECvdfHslP7r
JsMpUdW+BB1WVQzgOZjRIcw3qKlHwek5hwO0JtaboFTpjSaKItkAKWWoekVlSL4F
OhEVaDVStA4dT7jT4CTcVD049od42n532mdlOoAWCOAFHiVSt5Q8L4zeLi92kgBt
gGNmXmNXa5i+o3jDn4zNVA9w6+pphtcDnNTSPmgPJXFE9nae6KRdpcdpYfmq7Img
eg8aviWGecxn1BdPoAfLBAMQHWLhXLQQiSNOdZGUWzl634cw80GUBICrFjyCLIP9
LdjrIdKQKyq2CKnc3GLGPCYn1QJrIIyV3ZUwA3JT5g6/3rfc2TdMvWPZS28PZtcb
vohGp/AeFqXgG7yziuNlcptGV9qKLfzHCoySBr06INMgFLE361BVh4dpkzbFdYai
LAgHo/IcLN7vATis297ITSYAEjxDO39tzh1ZyoGC3xItGjzKaOh26vDqtx+IcBTO
FvmidjKaKv3CkZl6/Vi+r/9uRjp5iEHgu94d2lWjg7aoKDkb01YFTD5DPQZyabQe
lFIIyoB5YfwrlRSnNQSyymNQImBPd+UOmzrvktG/Adw2yl3EQmeFY3/H7Y8qso8T
xuh25VDYAnl1u38VssxxAl6OCzwJAqiSqL6c5w+fQmtv+6ZLN+8W5qdlaspHtzjD
fDIN64T3g1neaAsr7BAz8Udkk6K0d/zGMrxuGokgIelvygucoK45zSG+C2YkbIeP
W9YgctjdB30myHkPdvlUudICRnGjVuH1u7uURdU5+tE+ZEVr5gPwPLZVFtWfQKGI
LBL34h2sDo/pKebhkdQfyMGqUbe9IEHwPk/MxzxVyCsCS4OIF+9R/qa9DRs51PYS
N+tDRn2nbtOccAE3L5l4LHQmY+GthV8qbbzF8j7jACeEvza2R/Vb5glMi5pICIW+
sPm9+lWPG1s3SNBQDLr9oCNu67yC5LrrQJDCR3z4O+0rDabFZ9IYJ9LJ7d9/S+q+
1fIirE3y/YuL4IAA+1u9o6/hGMw99k2KJ9eHCuMp5CMVEEa9dci9uQeyU+phsN+f
eyX7/TsUDgObESclxGqAL1jHa65C2uTuhPM9RnIgK4p0NlF794bm8OPjG2NMnSM5
qitQaOTEIewpz0TpmZWxRcOmdYziPSSMyuTGIdBwD+Wph/XJimrfRwwEjaVl+0eL
m5QIScVxLoTbvukeKwNnyNAnbCdPJDQirW0E6RxY3U1mZgTWYfoXlBNikly2I+lu
1PtCOZlSZYnuY87W/wfOQgtc/GEOCUsHY3XVAalAUvPvqzaG802ndRqeKHp3ZbN1
zuptK26vt2Y56LT/XM7hDZ7pdDYWuqwnwLbQ6VvJb9QR6Jp1dp5nMHg4M1tk7gg/
hwTjtbF1SuiSMOJk104y0IZYIl4ooSi6LoEP6nlUNv4Ndr7BsA7JalFBKamERuoQ
5fWuzexdPa75xYyjaY+VdGLR5xcy0dRRxhYLa/cyr6ZyT6PdNN+Qf9hFKUZoIaQd
aHIMor46RtBSzEWkoapf+nCQZSJzxypLEPItRgVKOXVwBknqMOb0nqTu2y9kUpKx
jfpcvNjOe1FJsok7SfBWTLPOHNRIcXeIIiPFZLhbAwlOrL/ESbIZl1uSebphXopv
N/8WHJYAfeLvm0gGUMc/WI5YIlrl2fynRMZa5lY64v+NYCq0IVkf7dkCqDyjIlFX
6NFuGHRwtzWJvb1St4XTti6YC39F6giYPjEKJal671Ve0vK//aaxoYwnkPybqvH4
IM2UKf73+32/jf/COpICJrPDU+ijbXcKJesu1MbAYb5ZdOFT12zdVoSogaWqINV5
XDRNMpwoqcl9XK/jbuwX1HNcS2k5POBKgJzcDGuJhdpRUuzKc2l8go7NfpOdkl98
RyuB6U0NS2y22YyFbToC5ZoChT/mLgxS83UMmVtD1XNGMQ1HnxUnyBYWOrtG6zuk
u+YZklR7Ij3sOyHSfzrsbvQajmjsm6RsyvG0aILCA04p9R+ZqqbXGWOsU++6JuE/
TK41Iun351Tk7bfbXq1Uo0/iEZzaLDgdxIYrkfQ+aIm0bTZVLPXjHI/7WFDsZoXJ
K89q7kDf2QzyX1bXEVpkIxaGAXqlUBzbO9dYlkAqdegH8/2+1RgnKNIKXJU4JloF
GGblDuwNpRetwTVrM4wdYwgZar/rmYsrDsWNQuL3u2TUxQRSNRbflVvE7ROiljlx
tItnIQjfJmCHptL2FlMCXBm+eTgyPcQ7+pTmt3+Aif3z/pyryAJmKHw1rCsle0PF
khQgvFPOa3mZS4hbdyhe01gsvfaArJfdvEzx9W7Xi5om41h2oHoujL8fnsU/Yn6V
IE71CujtUzPFEO/6ISfjWlJv++MaCW+iH53+p7yDFZ+Sv+cLdt/Yhr5NlgyK7+6x
vmthRi48LFPak2T5Qf/w+xxO1Amw21HjfEY5Tr+P7qUrYUa5n+sTcNK+rUv6Sv96
d3MprIM9v5NU6OikO4xBr145CFaq2x/qSIryNH0viyS5CiqFFAL3BPrV0E4Cs7cK
HhACq8CFCgKQ/HbEF+IxAwHOoJsP1/H8FdeLsKoIwwa93jfKKdNeROmSgMwg78uP
oGgthxcAsiryU5mjBlSvYrx2n5YkJWpiYOGgHsq1i2IWLOK9yTBgiiJHpFAW9xJu
8VnTiZeCc0tKeW/2R76WiMmEEpF53qXQtLAOvKjh+XnpSGXjmWZPaOgMxaSap2bl
oGWwvprrwQJ1K+hlH7SE38V4zLrva+DrP6+f5uqXQQBht3+zyQsPtsC2RPX+86k2
cCjtDLaB67teEHj+L5uKeUYEqLFLeiKrXWYw89zGD3+WTUGIFPPbWsuP1rNEE6g7
ipwchRgId7+zvCI01AUOF7D8HBsX/VHTUiMtJhaJwIXEPDT6TPazHetraf0SHnnG
kYhnDU63Yu73dDCzukekbbOM8zLGkkxBTqO+eA2XHf+6ZPU1sKfBkPg8HQXqbSBs
sG2RDW8euw4xsI7b9bVVwZVHKly/RvXdODDezPC8QdtVdwrjG6WQTDK3m21gXJjs
6uc0bNPOQ1Vg+h/XaIkQR+TWE+4T3e6oP3OFQtXnGDvrZWS3uejcC05NQE6FRk2y
DUKStUqh4EoY3dkjgklIXmuW6ldtCFFKIalC5ch+xro9ri8GVWtE7OQw3ksbFAVj
SpfGcYTTVC0PGNEWOMLsjIFZok2Es3J2QWKi/RKIdO+VRROosYI44p/TUDNOf+i0
hWa5VkdXo7trVUTtVpnqDaZNlmEjQ/LbAqMsn3Ss3GyAPEViISml9FECMT/e3nch
Wgc8gyyCO1eP9yJX6tGmrqS2NxYXX8RhwET/9xg05JLfV7diy/4QR0hrKkxA9ZDN
sWz4NG3HIopXpwh5TFea/qlMRDdOEY9My1HtF5dA730QlwlzzPx+zfwADjUfWDkR
MUQyXjjFT/ha3U+ZddkwjW2jH83GvKt+ujnfzw15kR/R7Zk4mibrgiBt6sZBwW2K
CNENQpoTlGa0Z8RusZwaVJKfhMHE4so/EIg/cmUHBbQABVNgECuMfplSN6yw+qGv
RZRQeCsSF6mnF0EKv+tedPoV8VKtD0huNyVRXshmyGRAfshwvxEgcWkMci1KJU0J
JTJpevJmGftqyheXqv5CMP2bxksSzemmExFIsZn6n1R6QAVta8Micsk81DHy9dT7
yKph6wdQ2AlLoMNTnBb+GEA02PphVnyELeqh1vWLD3m+o6bJE8HK1Y9B5P1yYis4
YfMBp/h5Sti0xYyU3vB+nPEIFvApzfRFhETHguTgWGHwy34En94vE/xantt75BrE
IogQnQ7iIev10U4Kx9NDyOt6+j5Noq3zrNKwZqZNpW7vPNp0Hshcis+vJ+9wwdSm
nj9vVpVkY0s2VtPsmfzn51d+T607w2Idi5QAKr3Bg2IraFj08lPtV4ibDyWduKZU
UpWxZzVwRnuHvaKhErPQjVj0Wg1rM8WpS3akaqwQhbIJWxG7ADKYzoWiX8vREd39
/89vGde3GB4TrJjGFbO/JrhvzZw5rA3eVCdxhRKWGwXQQEtuQpCi0ugERNU0pbKp
T8N83jpfnXHKXZwjY/ISn8C7YDARGwEtzD3kZgyI+yFaKXlTX6XHFZDY+MhXuhQT
+AbvJ8FFJhy+6MJtfipGtbIgU2Cw36UqouzXFHYy5lecWS+TsInnPW7Bs5ZFKaJp
b12xt9czjp+baVYfmACFb4q2KDwMDhfl8v1t4KJm5kXSAGADFcSIeqdBEeYRTjmy
DB8eIIL7QduXrstHmEr9Og21FqySIdNBCcqkk+gS7DLmOsNUZNABWStCDSfX5z7v
REd2j1mN6MTVfnBqzhs8UgczwoZbXZoQljBVmAA6KrwqBdqIRRVrlcSciuEFe/Me
mmyz1SI+VyUpAzIkCWwlWNaO0X1H89V3+eZLuHBdIzh781lJeIQ8vH8SFvLOiz0i
/+3pfem5Ssvpq9xQhEA0k+cy5sorLeGd9KQxjKiVlA7KC1k1uF/8fizSQyPBYrRQ
Yqn3Gd1XoZMn3lBYi0ZxOv0VqeZ5N9mEBoezQw3rCZzVTzPUFDqXhHLw3nsBSd/9
7xAe+EurRZ7EUf6kRwCYN0MASeQOmUlML8Qivzws2lnWNPhh+knN9c+zzoPAXegI
V8Sj5PWWUriw4ZqNVf/69Lnl5qW1YJMDv6vf2iyenvrbaqXVDbv9ytgmxdw6PmTi
vtlcge6tfMHk7sJfNSjlktkj+hbPNFuxZXbKgs5w607fbrHP1SJbZKAEfKhoV1tg
jnlQppf4AOdrcJxx68m+lu793hYFlEiX6OurMRZfjzkFy9fuYSCfUlfun4IJkkkX
RMj2bobuHzIRWr5p9qEcsqdOeLcsT4YrWaGXdDs7fLO129lBLyz5F1nm+z9IpCRx
t5Wx+cUp9CXvgY3joPAjDllWDYAwGGfQgjwafKagclJw4Nb21hLDfJ6Hea7TfoUO
J4bosf2+yt7K1E7P6zJdOhXi82ck8G/EuoP3EV5OeMH4JB4U5KjU5wz1VAsajCFs
uc0Zjg9Mknpb4X1k414JmhPTzHTKGniXZxyJgeQMJ0AAlsOcJY1zCRKd4vCvWoN/
EgxFEs1/lapEI7EvgAuIOdkNnnT55oCCZDTXKR0rdqpUOXm6AjjEKmD67vi8xsoN
5jxvkzYtiPRK8MhGeuf9NtbBmaUZB/QlUfz6mdl5WGMIWdgJ9Plw4EZHLZeU0/dZ
DX/Sl8Tm9JDETy4TMLTQyd1wU7aYwwJ6DLVtqqn8foacEKKVyNi/01U+hxe/0WPY
q11cfm6wfFwhC23axp8K+v8+7YbVbBHEx9Vc/qTLkTR6R/B/pGICe4FbQY9MvDR+
0EKfrYb10BSdR6KfuLnHyG/qPlN88NTquirQqgrfDcrzV2KyywxQcacWAaQQPvR6
bqKaMqWh7lKy6oho7om7fdlwb0F/k6p4mRY2usgdtaIuZ5H8BsIH1ccgGTWF0KY/
uMBFd7MLNNulYREqQ15sKCmyv+a34DxNHBa1/9R4u8+f9BaKwuL2jijrEvAsIuoU
PoAldPT7w0e94Q47fkjJU9Zzyey6OZooII2xOUdk8tW+cbrjno1cCHhqyWMH7WQL
Dh8pqLcRoFdb2VvnXAmTfBffIQtdJguRUYxThaxziSV00LcfWqy7ilw57mJtQLaz
6x8g7Ric6rgLXMzz3mT5HIPUZGAziWZreq/0hEOssR5I2TmBGTkJ5GOzm9Bho11m
ijapOc75neUD8dsEeT1m82I5Ht+EkhIHrTBA/KDfLUFAynqkv7unxAs+ld/VWBzh
IT4drJFuZftJ3KbNLwhdcQ==
`pragma protect end_protected
