`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
UiVTLE5nbuiT/X3povhUycxU0xA2kgAsjLQNA69eha8PKC0ZmVsZ351RdIPpjOUU
1sJEUQW1YKyYgKcVGFdaU3hWvXOiebdzgftGn0DUpDvvjuCI7z4HupRMdEsYWTJz
83RGqFaWtghHR0bDhmEnPaCOLqo7CfpmEMDKnTa0byM=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 6208), data_block
MWI4qpYDgQ7FXKH5c1FcfevNYexgccXf88QGkkTTTM1X+4Z++HcTez7YWwDfGUHo
rJVBVIiI0H2ww1L2s/ZxOlMzqXtVM0x4Flg24g0DvvOEdQGaUGxIrhGUlHuzLyKa
zDZaIjReVK0gv/b6S+NkKNIOiAqDCgrau3aeLOnvgsGGyFvAxGBXagNnL0unSrqg
6Q9wU7gvMDOOGwnnWZSp/k1HEijAz6gxfv4B35xl36ZoU/zjUX4ROcYOjaXjblkx
aZksU/btoeT359anDfkRPa/ZXdPWI21uTqKl4jtMufd1lfwFYIidaIsPLVDXE3M0
dC3IHZ4iigpyXztAFWczQh07lvMGmzZXcmiPj/Ov8EgpE+VhMEa8aYcd0Q8dGOLN
TSkeFk6aTjAZ6Q+d614yFZm8aNq1vaB/3CVyUvMnrT8Sd7N+OJ8yZV4gOZpUS+/c
F9tZEyPQTV//XynufiKf0o4HD4M3inYLZO+LCrx483+V5jt7ZuSsEYli6pRpxWu7
qjmsmAA0paDg0tFsXaojF6MLaeyrt0CDofsl+Ego7QdkrWq10w3k/qXroewYCVhG
9VtOaA68QH6TNHAn139FCW6pAqa8Qr+OTE9Tp+m71VfXSloyAkGh9DSFP9j5P0Bb
bVgB5SrGPjHz9y9de6IChspY47+0DknpgmJjOHsOYish7a8KyUEsX/e1S6fqTLtc
l4ZJOnKH+DYmfbRQN7IjPEo5lTQX/yV2zHyCJiNiRvLfuznJ5XIkobbaJ/Jufewe
7FTaGx5yQ5wyzRQqa/sKGjnSt3rcagZ4T5W64srFbX5Ge6eVRDZCb6t7v4Vl9tyr
KUKVnUCEZhBRTxY/k8g99h7IR/EHXIuuE1wAF4zLfo5Jzg7M0YwI9D15ei0Sy1zX
sr0k9pgsBOMfraAL7mtTk3U8o4KTqdT8XJWnuTxmEOM+wb0Lh3Ybgc9WF3He7yn6
LOyXaIk6+DZYYE/7nG9Js+vSmv5cV1iTJTG3KtNuUeuQ/8eZOO5LzTohqq+P2nb6
BhETYIKvSPpw9lDNRs44MNoNH4HQz/sgne5R9MulPtQn+nlk5NXkeZZzWLr5Bh4W
ApGQLmSLrpE82+wXlkWJkw4/zNpy3rZr2wCvBdyjn0f/cuRMeNsMpf+mwXEstC9Q
qJagmQH82p5VBUZk4QiTnqidNnvv8PdnNepAzT2ZzersBM6oxYl27eCB+Qfn47pq
LJ1Dkjg9LxeG1BxFQtvyGtyP/0EMN7xWW/WBbDhomWevCGxEKobjnhomYWYuADLm
Mts8Slmcd90QobLKgE3zD/qQsc6eYVnukvDinedkc0Zjom+Dj8AqmbTZJDIclsmY
LIPZV2ZqUFS+iPpEzNvTt6bvaaiHy+TGM4UKg4ZEwK7qhGIdRZKROnndhfwvjLkI
u4D80IU/a6w6b3W0jrCv+HP4mQDNXOOuzfMimSKuHFXN0DXgrgLCU6cReXQDYEBm
pefgS33Xc7E7j8ph/TK8wK1Y0I0OiTEZbTzSt5f6xiVUz+3y2zbqneCY6hSkPd2k
b8FjRkYrFTAhiJCxlWOQ/OxwmkQt/ttonOw4GsdP2eLOIrVunp4HwcUaWmkUlTIk
R38MfvXgjhsOhEsrfxfnxWAkH7VDhPNtDPg/JLQlOKvT1idy8ojzIIrZKUSkT2Al
KvIntJ3ZtH1RQLlgu1QKTrwgyEKQWYfqOH7X0wb+no71ed255I4ryxzoFZ7BHkdS
rv0SvDg9HHYefegQJ1DdqHlZRwXLiC5ylHmOoptwq4TQ6JH1FntzJbe6yxv9MiiK
Jtlo/uaBfCbivdXLkIiXFJIcXGPc4VB2mptyRuMmY/9uIYt1ZQmVx2aG80elgcVW
ZU0T103WJ/n8fXrMfLHpl3QZIno30fwuiyZzGUbKop4F6WBZJUzuajWEGSm35dVH
YwcGzCvtbxlgy7mXYutxDaKIqZEVsOWtDFqwsQTo5Ny1ofqBICoXbwVlcwanDEb8
CQESI3ZGATCR0+PlK7vD7AE5nA3vrOAv9zm+Czgio9fd2X/DmHyOFLnSyWu7aTIz
MKn3b/aVRZBgavra4jFIclk2CU1FI0N3BBWJKrxi1l9SSDqhI/mxEZVzOa5yu6AM
DEQar+llyFOXyv1KWby2F0IcG3R3yN9nJmGOgCb8OmyXSB/CyzI5ce0L5avOkcIv
Wv0446tb1EFziRqiJ6HXT4UuoyhUR3nr3QdhJX3OB0zQUoZAR3F608U4ous4PCuq
FlPj5H0UZZSXOAPy3rsKTen46yLtATLF2Q3MihWTmbipCNCyHmki+QdTivmrSDLH
miojCKSUgSuUwWCz8skff9p3AVsXrP8io2ubDFd0nhSSAYlNpxLobAmOqwGFu5OR
l+J86LhpXzD87gEbv7dyboZA3YZfkJ0KCAvf96JEbq+h5/+f9c9jsK49PFNNNQ/F
73l4gC9gLwKpYVBtwAsHPUAAZRxwUQKb0wmH6OgdSJmurjoWbLG0iBCmViXzuaJC
/sRzNjtj/MI5/x9MR1NuY5njuz/l9OCuAp4fyk6aqICFg6oVat7vCyDb+KgTN+Qq
XSPWDonxs3DPENhYQeOqq0+7gmTUxNepA0VeFY4NWZxHdKAAF73mvFfP9KzwU9C4
eYcsNzcn+XtS8D4pLDIXueeAWZAne0hTQCMZC6DDBMn1eoOXtZPwbwKqmV24RmlN
oDkIgagyInEYfL1Sy17dS57vUYa0vDunrEo3lkQT6PHG2z2C6MkmzSJdWXbXNClo
GjhgIOB7ppAbT9oi9YpxdxzTt874m//CHzRtRs3yPbGYkuo9kzz7uNZCZSpIHDAS
vDQpJONW0XPN8tQVnmNmf79kT9EFgr8EIsUeLGsZ4ui5dGMUDpElccNIi2lNjbQu
psoDC6B5J/UrGzrH9BfdxWFUBmCovff3kZEwXr0BMJKWTBX1GqfY/LNrl5r+dTLF
BYY9R9MpeqwXmSCe4N8A56ZW2jxd/s3LrCCan6VqUl6QhgyI6r44EmGpk15VzIDW
cz27ysCYvxB7nvPDsZpqMJVFuAyakYS6kUHf9Y2T79TCAGRYZxt6jLGnUYc1k7hN
4ZeQCPQPhnKlo0L2ATHyb2ChfrzBZ+6xvWpkxA5l8xQ/MHRPqpfBvE1dIpw5OO5m
Gy/1W9jk2FgTlqWdPjMWDxYIkKoobAr5lI87TRrxWsxH2MkjrYuSoGByY9K7fMyx
OJGrweDLyBheSTfea0jOV+NZkXWiGyegczg5gtAstNrvOQHjk16oZRQ4Cm3bxpeG
Uzs4az9lfX5J9FL8L4TCsIADdaMixjawFZR0WDcB24/CAibzspctFvZUoF7JHDmM
nKUW9C+zG7L7zIV4so7nDRu6l57dd4ceZ1+UAEusJAVaGUegTS51Ok38Srin4kWP
rij7lbwqUTev0+gbco64X7q4t+FSE8/51Mr+tT0MPfIZhKAcELwwtlAoVOr0u8AJ
TyZLulX/3e6WsN4JLqjHBVOqlrCB1BYkU6RrOB4QAIfFP6MqHc1vvK985ZXyu6BB
GTImL9Yh92r60x42eIvXvDTAhxFtxdV2R0jxG2YcrbJajd7Yt2xOE+4ZFbQPfGy2
gc4UKDc92qZEC5AkXFf/0vF13PpaL1HNMtJZdqxkHKmGKDBMtcdi8FKSxHCqNNBB
4RsyukCcxtTd0AlFEZ3NEjmQ9ZdSXZ93VUuUQj4Ks8g8Kjfblk8mghQrPqJ02XXp
DZkoiC7lxX00SqryIJ97s5+GPeXKkOTaztOSLayX3pj6YxGVSdQRCeAwNDghoRUb
F6QsWXqj66W5KBXwhrRSVq1cDGrvKOLjukneRGXjBJHO1ZaCkKvnkpzxeh73F7Sk
VYKxzgieVEg/mbjfr0NpJ2UodvNtN2Y5ZK3Tf2yP1bvCLZ3HD8N0lKLOY8IkS5Dk
34aydNsMYmFge3MgCO2BjyDKd5PPCnXbzLpmVLqXrMQdCIt3yf06ImiOdUx6Et88
zeRTv662okrDLqCpWf0wAgUuP1wRRWUXfCHS0EsxsXjCxn0rRX45tQyJPMIRDpcO
U9xbPvn5MoPQ9ZRtavFyyiev1S54BZCUXbwLToiejvYnZ7SQuNb+BLaXBqRefRDs
oyfwPkolv5V5YdcevSMPyuYHxqrxr6aOLDWhv7FsATUYBDogTXOlbGYs8TEoC2c2
EnNHclZMsomMfp5DamD3PrsOiwlavLTrX/j6I8aLlHh/CsW4Wi3t0QTTeQrivjWj
PddbuZK1lVQDTRXemAsSe6x33RvTnruU0Hw2xQi4pqRzkpvFLoss1Evz7iX5IFJ3
OuvFcUa1GC4tmknE/4Zo4tfLYORxzZN1g1ZKviDuI4s4UbduFyvmoEaZ2+XuIL5v
qkYjnyOAuld/dDgEw7vd1iR48+aDfNfRnvRjJ1rmHJPxeNMOHVZpuoUV1Wf97RFQ
2sSK9GFdTn1MqSYIbCMDhNgQ/5Ub7Qf+hnMdAzODenOaomkXLf1DMc3ZlcirgHMj
bEvjHQIxrsCdJVrZH2EhgV/3TnIMzYyXO8vMy8/YFJbnXqGp2jet9jq7vFQ1567N
W7S0hpYNqy9pgGfMfSJjoslyaIHTd72E8JU9zR63BcssOy+NZ0vo7Xe5Fly8WDJU
OFgZHLMifNNi6B1DWzJdfeXakPxyre+XlwEAD578v1lpi/TikXxOClN2mNnA1DqT
kruK+VpszC+AK2icShhilh3Yek7NQBVmgpC0EyDHdBVAbQhI29mB3aZ/Igg51Xqe
zXcskwMZhnbjNAflWQfMmDE5nxhtfa2FJnSP7d7ISmrTTglQuCrQhFLzYVmvoQ7W
oXjwNRGyDJNfvN8fBCCavhCWXPUrYlAAygx0S6j1ZqsE6HjgPIlxnJjSb+ZOjAmN
5vk0CkMYL+uI+w2mC5hqpBIt+vZxE8X2t2JRFLzOPmI5sIRfd8dKToEVI0hRqkrG
8VqhBbtFQk8xMBEAux5u4653FL10TRkrZQuWVU82G6wyf//JL7xRhVcK6ZwueMkT
/3FuE4L0TDTpWPKmXd3qMh3gwVSKj77RZ9iBGip6XMbHQn+ifjnXneGDpK2TKztN
8q0Q4YiOeBJ4pgmx0DclfEXj2lhQyW89iiBum4auX/qDh9oW3ZEQkZTa3Hdw0y3X
9sqhwcpHCU8Mbee2tfFWpYquNz3eWtxQpkkGcBdMT7qPwkoNjrJIPBMHM1rMnL00
fIFCWLprcUFgYWHNrccTgdSFpmTeOIiVGLlVL+H70/zwn9LozfdqMp0iB3afeCbH
arwOvbRT9m2rlJsfxOzEF/7LKDoyko+EdRZOmZ8z8VukjLom5DiOaBehc2MyIo3/
JPPWMruke7NMUIh26XuWPDp10Ma9dnSPkcuQHHeVajydod2BUl1kd+gqnpbQOSQ4
Z7++qk6paEgVT4wItxy3IE2577ZmiBNsjncJMGyZHL4wpe9IxYmInfwzAKgR1hhL
5XZRA1VfZCnd8PGJlVAxbtElIRWXwcU56fFj3vDaleveW9mnfPfj4bzYPTIrgLkv
qm2HLox0GHN61rXAFmUTQGhKGd6lTGqzn+eKWfHN+kKGBLORtIpZ21fAHAr7YWuP
ABf0jsqZqbBqlb6c+Gb64MEOTmdK2TXsywMjtFSqVYZ+c5YRPRcjaYM+e9SQFTWy
T5ETxPqHpSqT64+3JdqzQLdV15oolE1NMfx58xYsqAV9na912FcYUmrnakYMzTkZ
iQKQt2vh9AjCrJ82CPMFWQRg02wD/MOxf8yIT4lkeDc+e6KgFboiUAi5g6q3eXhu
SwSrsuRtESZN975al5hpdUThhrHpbgH0MOr7EtwqMMFH5/XDzFLvXtgZZOrg0RT6
OhlWAmStB6bzffGRSIj7egdGLSw3YTEU9m81r9ys7jH1UXBmkHBSnUVGYloiRzuF
ZfNEgDLMx8Wj674Oa4zc6LGTAgGDKSNGrc07r2A4vmtxt4TTZkbKoyo0wCDu0T1j
U5CBCFHIyvumD0tX7Yg1yZgSixL33pc1zefSMoDlKatuTW8IrUU2vWvOxuzCTg11
Jn4p6wh5ABD6XED/DgSlNj9fibhEQB6FNJnpGvuBFHcmJ4J31Ia6TPxRPzGdnzIk
OZXPcqnVBXSR8bGGTepod2DD5XNOJT5ciDsEdPhPv2+MulPX5aBZlgbBeSwjAUOX
CQZ5hqspN9/l+CN39VILS9a0Yg9c7pqcyTQ8fjiPOJ2ttPGGpOOskhEuo5mvUSbT
/ajgAOL/fJkN2K1q1M53b7avKxzgnGIQqyou5whTOR4v76oqVF3KlxSf6ZcdnwTg
vKwbbQea5akv2JSTHXbwXE5qGkBE3mIvq9jwDuNosYyMu+OGMYG5SwMuCleWYdLD
LJsT5PpiQg0REzsPImb1Sezkoo9bfJIvDw753G6jrAto8N3yXJh0Z2fJOyVkFrAU
5uJPaP3SMrzAptEeTHMqhRa5dLCR+lYaPttKKRQxf8FPZQmogSNYuIuVytdn859o
zeZ0rgCIdVe3GtKaCZvMsVNx+5d0P9evi4P4JDVhR3cEz+vnhyZzLSVjImpO6F7X
3JLdEKjopuMdPWuF6KGsECDBuGkeztT5ApINLILVxOGOkuwaAdkgabLvXRfkzyhs
QwtF/P4WwUY/dNiZdErivRF7wjpTZWaIyPtykglRvr3/JrSwcuKhL8gj5iQbHPmb
pubut812lrD7YbNKCMDMXq1i5gKiiGC1ZFXusyazTXWzRcEDMNveyISoh+T/IRPK
veSXLX5i0G6pK+hp4mFAW2el0yTOcUKc76UsTTPkrMKP8HQdQBOoEyX5+nJeW6Nd
S7kWrk1emS474R6L1vjCnZtRBYs4p2NWOjSgRlXthC9O7JEPbOrjCaGHr1/TyH+K
p0Ac9GOGk8ODxkKI2ujRsvNCM/8lI74k2FgkqIm/vUjACtMSXgAjJTa896RDOtzq
6HqBMM31UAIhkVbhBlR4XNK1X+NRG3KAc8tq5rENG58oUjmew0pkUzKQkjiBUnAY
PpzlbJgy74YjaHJ9999wrPflRvai7/Qw7URThRaZXEWfKk+J/zLjf4Fh/u6yfywH
V09JvaCRad5DD6gtTD/b+snVIjG1tU86amb0waB3pqZZjGM2fo2zJ6JjZkT1kfio
R8ry6iEJpO8sGtLehpZEHXYy6VS39FfLgqdSr1a2mWmiQGOZo/sk4TJ3FTaful7y
Wlvn/+CSJ3AjqCrZfV0+Di5w9lBO2ACMXz2FyMFKJstscyYs2yN1IkFDuCB2+y9H
fSeqPQBNxno6vRj5RAMokKTvxpWFPdUqIsYhRZaYMukWfhhYnly8+v7qbYBNWYbw
vbJO7zs7XVhkKc0TSy6Uu2D9cyL2DPw7DTerGWN8X20wmdPmwatQnF0ShERiox35
V+cF/7XD9BlpapfRwRi24zLovTUNwNAU5bwlFBumlBRM1HIgW2V13JZfbWmAhwan
0U0Iy9pZzpssYj+Pf6Xgsmf4sRAf8FZ3aVzx9H1S+kRnYHGBoCspwpsUuPqSjt68
5m+9xP8XcWPorlc3tVGCblQgOhMpmjXpiKelbykth30n0WWSsQPXlzH2xGYhBlcY
MBSrn7XMUZQ1eMQ3l2UlT/eJzxq0GC0yXOsfZ7FjyB3mbeQyMECp0XvY8WDz7h9w
g8tGmOS5fu6eDRxJlqvAHEalgIjUwVfrilUv6WNfYFFEXs8nGSDXI3s682QykpmT
MufB576m9a4xia6LNiW36xLhKAlkaDcqRKElFwbqRx5c312J+7qC2c/gZqkvhLfV
7CYRSessFh6NT3gwVO3E4ME+lL7RQyO1QrGPfZ0GAaJJmSApBsCXORPBwCa+A9hd
/jFuSr7AC+05p7IeprCA2zaep6L0/d+a0ysMSjy3KtJUZoJp2mJBKfSr2BHTgAPp
W2sBdUwy7R61WiWALo2+5Pa4/ykF9IFYRWWF89ZOreawJJoET9QJny/5vl9pIJ5e
FMT5WFY7zGUWvIlVEumXEZMaaL6ojQOEFqYuQcZrgXaUCfpq5A7BCBkcEjyWXR9v
UORRGedK5HdR+vfTXaVoOGESVL2iB/ycI/twlhnp741kOjibpHisnNbf5lR4cW3B
u/cpLmr7356L7JDeffr3bKQrLsUM+g5MNUkhD7X3KBzbFz+nPCIjFbd4ta5mJcoe
7V03Mp5ZUkrUh518KZXAfskiVqex1D/z0UhDdlu3jOuoz9xmkP25/mXbqdGBNAMN
Rh2wFiJM5DX/GgLm6bPB1HcV8e8HnkPN2vVblAHm03s0A/fOS+O+U862ejtHWuu3
6qF35KAWC/ZtJoxIRxd/7A==
`pragma protect end_protected
