// (C) 2001-2021 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
ba0hP4Np3FgMGg1JbiHo0CG3/sQYuY+AmokSkOB9tAYjscmxQNqVszaJDtKhjZ9sPabaSOHSFSul
6COPTs8DBCavDDI7ZI05I9MESBT0OY0c/AllqhFwC2kx1Q4lKWeWrNkSb3+Fvr8nzteXMDcfTnT/
uzIJE7NlIaqzdr3F+oLU1xcIl2oewHCUJ6RGBufxjVMV3wGCck9rrpvJp28o6K62XyfxYJVV94d1
C3gKJ2QObV9NNHXsbV4wNTZqI82biDhulv+INzbRU/AUiDo7H62qkgmHko5RvC+A1U00Q55OyFoO
O8laTmaskiryO2n8cXvR1rSDGjCp+d/Dyu3Wlw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 9248)
kiCLUV4udTV7jRYbQkZ4JA8CXt1RWLUpJy+oLVylRiMNt2iyDnvLCXoSSsk0lRwOoWhcdP9fjlLF
5boLGrU+0uMLydmFxafm2Ljen/0CDG+FhBbIyZW1KK8eOpKdpAoCSPofCkzno9nCKspdm/tKQ6dj
Z8L3hdrbSakepIhuU593kIQFGKtTpN6bULC/uQjIw9tp1thGMSO6TmjrcVJjEhRwZHzOAVtWkdtF
ZQpiphS7gg97ozXVEyp2rAtYvYJz8mfaIcub2GHsEe+xBPAmi7FsEOGobJdNRaS5Lw9fPiHrfOnk
9OIBNSlesArMqfq2smrns98fQKY36YVX8ykvuYId4pwkS4n0ONI5TgRBG/DWUTdXJAI4N6RBh17M
qV97S/a3CMPO74/Wmtcrr7Xuk367y92WlI5Rx61XBIDRA6at+sn35S6YgNdmpq2MzdKoYOjuCyZL
GtnEa7mK7E/GWzoYCqGMCfk2ZPq5nTd1mixQx2jXF352B0RzMJS1sN/glP21Xddvng/iSg1oeNWP
gZte73gcjtb3tDE+cVByvoB+VdQj6QjBS+4thLW4pm6syzL7uuohR+gIxHtUiBqKXbAiSajak2wR
HxdByhxIxzQ3IgKwCYfagGF1+YESfHn8nj1t+G/66Jl1GiiJFdXbU2PMfsEhOo3cB3O275I+gG9G
M604FMyQEELvynEZojiLKNtEVpZNnJqrN35CpwDV41a0SkemH0lT0AcRosuMhgYV3it7bp+p3Mo5
+WfSFh+PW4/hBexvzw9lGmfe7+jNlz6L5t0T/CtBfdv0r4el+NBC/UE+BPbJ75UYAvyF17y0yQdb
KYZRfNMILRYvHnhlunBv5SNt+foZIOWiJ38UndfP7JGuC9GZdPZ9zpXz7KTL3l4R52K1KZygf4Uj
q+ny5S9X2E7/IrUlmLU0DeY75KrOaOeV4aGwns7DNWWQKHCp7ghiXgR3E1IjDL1INFGihF4ZPYOi
BmdnAr/DYPJxS1n0iSL9nIC16itfHW4MVWF1vwndCGZ+GgBrx2IjmgwXUEMnM4zI4z630hU6wBcE
Ckcy4tsG31i+a8o8pp0+T7Zno5jTcaO2nGCUWLT7XDaWqp6SjKZYwVk9rWrOeIBYUeQpB6H3gYYj
9qiKIJQYNbrOFsYkTzQp0a/+buC0nytPIvq1ZIdqMzERYPZ04eyobrhILjHaeLKPYIoopxntInPJ
huq82lZnfvbBuaYzhK7inczrOcgy2JRJmgw1cbbTii+wlKkv7FS6zY2RKVn1CxBpDGCtpeZ14vkV
esGC7ojIjeQ4tBNlRNK9zfLUgC+xrwT4oMgbWPv2YSvYuSZjRLxqo/ZZojFGwuGNECZWxxSHlouH
nVTdXT0xq7qIULM9r4+nt6HYBxvo8Lhpn2dByvaxBOdNW4aSXcb4IiBOBx2uVFjs3qJSVpos9Wkr
KStsfahf4C+0PT2bhWWyDhTLujJAkhwWjcsv71TpHyaWlYJ3pW6tURQkObPbUwWKJnKwxd87EATs
Pfw/5tPRhWNehbCw71u3nUrEZQ3DrjlKlamrgzvCSIUqmk3gfSfwHozElB575YTiJYK/eoZlSwlQ
mj+6Zo+rb7a/+RzuukGOQHq33qor1HqjZklhNy0pqmxmuZ0ziWQTSz+v0XWvVXV5rNjP5jOsJqbi
89ecf7BGmeTg4zQBPmmIoYUooaiY/Ik8bjwBw4yZp1T1B7yEQMtJuMS/NkbuCWdn8W40r2jDkkVV
7I/oq8D+DSgTT1fQaGuAH6ULdOw/mTqD9ZU2sBT6gi7+lCr9xQuA5gMOwnkloZ090pTkloeCQUMF
7QaKfrDR/oY1h74k/gFQfE9sDt6mgAEta3kWE2d4Z+9PUU5h72y/dgtwheo1Z0kl3o7Rq93yJKkw
Q/4UkQjyC0oXqV73kegZQ9fhqjM1Xmxv1Gyc1qnBlQBbwoOOTNFQIN6WtGk3nqHBWCUpeiG1Da51
KVzYt8jSAjjMwHTs1hQHL/h/JVonubt6UBB+0KRDhp34XT51vWsjidaXC3GtjXuMZIy5BFFiYTzk
opfQxYtPF0PbUme5Ot4Jb7EIMMwZHeFJ55n1aCxe8C7Ia/qR2lyCNwz1HBlnuEogUNyzZxYuqTpz
S24liEkrzPoACkz/kZfjrSvyXEAAkA+gRSo2COb2tURn/DoTsVINsdiDPrpNMeaFtUNGBzStfg0E
zBWwRl8TKlPuiEm+r2Ek8wQzQaW4MK9i1JH65QNlwMkFIzAOJEEjZM/uYaBW/IoNrmVJCMKrBjgz
0VUsRGDc2Lbf7CxySRa81mX9m6Uwgkvd6i0OEtpOE3EgHr+sz2j9LYUxDGTCgmaau/7pZzG/ANZ2
yiAhCe8vt22AIFxCQuZs4WX0oTEErHT0VSD4WcHH/gPtF94qKoKLh3MBgbMj936ZKHyt0ini9g5z
anEjSp6GLDhWpsWuI0D3Y2ozy9mkw2B9bYuove8Kg92ikWZit34MrvSY8TWslO+LeZVmSPMoPOlE
oJdTwTp+jP3U/YtrTJ3JiIhSpi3kleefy3R1ylqp5DSftI08a2VSgNYjFpUJ6abKZFneiXSedD7A
Moi3z4zX7kw0p9Vbtbm0wgBU1FqvJkzG1Ar5XMYFnA88rSXNh0cXSrrlEus6bjusb7+Mt9DJkGUO
f/+9Y3/SQVnp23cwopwT8yWRFG3Ba0UyA3mfM3TbUhF/TLZIVCNZxlRU/EwHIlL8fa1ANJf1t70e
zeueA+T5EUGBayBSj68wbnEIiWVmb/DVlT7uMWn0voLYPpkvsSAFHiXdn/ME7lHzCZuEUEg2qLE8
GDSXJ0TRoe+YsP0g89NArMU9pMxWYjiaoTe3oCoY0aRoq3QH9ZWa2IXCovUGlrJd4nFHsrRRwHEK
aP4y//hUkhH8MpPIvauMBF9Y/IDs0W0cJk3+2UgFS8SnG8/xOWZouBYgNY/u7LiUMHaZfEXRpLda
MQ8dSfwGkzfR6lAYqW2twZ2364iJKFYuYNFDKSW9rM1my3zlZ4EmYkN7wnE9EDEvptnViGl5i+2e
REbJmcmh4ZwPkjGj+yEXuzuNPdVTzT/l2RbP6wPoRRvd9kMh1KxhIdQE0suS7AEIyAbkenNZike7
ekcrjtzt1fX5soxTue878bGTT5+/XoV7Z/2Xn7N6P950mtmmvixj075ZB9jmLTaBuQhgEVlG0hHm
mqq4gAsRgL1shjBLh4I+Qllno5LzJ5fSZ/LXzxWvG0kyxetlPTgvYTnjy3VzahROVkrTkzG8oWfV
CLIYddjpUOFNI1kB5lZnq5ruJMiQK98b7l8EJZEZCMy+u1YHNFzgd6c7+m6HB4oYYhcjOTTS6BqO
MVjx0W+ObCjzUgFxp1k6CUuowl/H9nwoN36KAM+9TYo4jzI14yRWo6hojlCq6DTs4YXVLvoq9XBz
IhtMTiIxI3Hzxr+/eCG/2Nm/axmGzpH6KaUPzVeFAYNWAHfF9kjbPLz6M6JKLRtm9kK5hniDeYi2
JbQibMgm1mgMi5CvFsS4jlE+93cQejlY1b1Hmo7XrvE812vDL5cmtkAoymNsS9rxVGEEsXcGOA6U
7doH/77pzE70772GB5p7dlt/+Vi51SqIA5S/LV72q6KOhJMaaEwjRLaTQx4J1HlIemi2NnySgBfS
l8PVvmjNfH70ckat9WrS+coSRqwkLbAYHwIEPlkZZjrD8Ke3iL7PvU3jmNT7opa4r7zYb1IahHmD
2RelKGMFUWdEUkgryuz8kxPk5KZRhBEqAO0u7p6tELWvWMS4rstbYo0GFwDldKwXvbP4N38sGLO5
c/oqh9ievb+LqdgPv/SdwHdLxbh+Zt3Be4zAIEOJoLl9oLmLHlbpVSFHog36Cw22LS2eeszoNOsG
d8mqc69FAyxtGEh3jiPTeMPG/yqsaoWbKhyQJP4AYNOsUHe2Wu3N5IP+VA1iIZVykpSC0JfyVXi5
PNw+pHXA8DMNzE/EZTiWaLEdcOhAjuNfC4YNCcrAaB/alnmCDC5aek7syFmi2aNQHrtqf//KqBnP
zeZsV4UkW1Uth7hBhycRBMiMLOFN6iZfQMp7QC28r8HsYMESZJQp2f68ziGozCDbBBcMHTA2h2kI
SFWVzDdB0U1S78UyKLZysaxiB4HQ5QJvOUQmGNWksXx/HoY0GIl3+11aJaSn8GkroM5HISir5xRx
Y5MwNemJmUzLquXvjVEbNHi2qtUjcHzhi3beNmzWb1kaFgDkvUFRJ8B8llO6zaIEHTXVZBw/oVjE
zh2In82tA01G9ZBWGy8Pr4ZC3ibLg9x8AMAT6YiEQG2hHDm88Ts/BMZCmGPFOq0XludQIyDmIAma
f8i//BLZyKFiRhdZYTwScGX7Vjad55eU7IwVPdEUjjaqpFEtrIGH+cFgzI6SXNs3uyqh8egqKDYA
sW0u+QhhaBD8m4kX6SdITEzH1ApR0F4rqToO4rSmqyIXkc8MZ8e+64vPa2hcUr1TZVgf7DTutXUB
wTWk+JCXkC2P8/lKHQZuCIbKplctzl8wfI68FKbkQQqdmRNKCk6Abb0ok5N8npzt3MQw7tnEe+qU
vel/M8Z+rgmqJu/RWGDZb34Q290gsMuKOSfvxkYBB4jy4bU18+BoSRwmznhZnyGfPM/g6ujh0IVn
GuQ0HIGbbxb7Txy1vsosKuvUpSvrD4mfpLP6zCGDWI6cRFSBHi0VnEUi0oORBUCIykz417z7Gsie
oejVpiqo8m5mQWy/1cLz3B4xhvq1hOnuRSY4tLE+UO/CC+v77Y++dH7CsVaHsPhnq7CXXxm0+wk5
Z39/JhrrTKyU0b4WnEq1E31jous9NH0oyvcdo7MbP8jBPnWIvoCnA+Q+xEaqZA1ZypbR5BowHLT5
LSv2HIDRqIq01X0XydET9TpksjMDGh/LIHP2MCc8rHINJ/dnvSY+Hwg4YtAV0ippZ6p/+S9uRcuI
urW975/uZPjt6+P9RWmwxT2p6aIypydsCc1sbLXJwyyclLL5Aq9uA740f+SeV1o5dLtqYxpbf+5s
SWjHQg1HGR9MclLsAZMBqNJLghiNDyOKExqF9iPkpxetMgSGIAPfO0fFPnV5KyyouzkRouvtr91f
H0vcYyEiXg635HVF0MQYzAgO49bzHi+LYqNhV7C8itAsSkMv1SNl6lxLd2fnQvE3diZXFs0zb7Gx
LtbXha/22UpvKZqpkzuhb4c4WZgIxtQUfkBwM+CWnD9yLeobOsWLchABHjjmk84SYDoXIXFDq9zX
11qXo9YnY9C+R368YsZPYpSs5V7HRvsXkKzq9mlSi1JXMZGbbG1dk1kKEjx2ekhm1QxGeGg604Pa
GDytVLQ4UpCgv0M2kkvWBTpAMRlc1twjVbzWXdpqbqNWo/ZG55jQb2MmjVUkgZepnWjdrecPH7GI
J537/rFdKXy2oIs2cuyWwEolDZgcTPn9IEBXtC6d/PTI2MRX7bsjUZeBQlwAX47dsI+PlqP6OAns
eYi9XQkNAjMwkIEXjtw8wTjt8g2n3o5MUErkj4xuMaglTMaLyJVQLg6SMO+8qoOoiNYfP0uFllDG
iYyBrrEtGufxW0aO1PqNs0S0/GaZcvjSJZX9A6gABDPM3+/hk5R3Z6mhKb/Csz511yto7KxPBvMq
glaHyyAxz5zS8ZSuqsT5S70TyYVT+Sq/MGW991+W54+AKVXxOFGjqF4+cgzBUGKVK3d02ATbimjc
OFXGWKrnN+Y6eIqXi0eDfFE4qAzz7q7yfh6ff8M2DBsr6ia0Bfhh9F0noddzWaUyTWDyBnyg6pxN
RiaKDu91YsOaF8KYyFjNZjUq92ZCx4h+ASH5g0TZurflYZl6u89bpC5LDM4I3/o+b0NxM/a9K38a
6qNrB83x5sYY+m/pIliXQpzXva/Fo4JjVh20u9XqP4wr/t4TZIC2V7wHcWGaefmYep+aveZmIU5s
XlBrihQAPm2kdwjGMq3tf69ijTgTCBrVb6GHwN/YRXR0Y208Sj85zr+Vhn5UDWBCi4Ivt8YeoUVY
cClWFupsy9lZsBz5QHHu2g9iu9KsUzU3MhgMTyYT47YvGExi87K8TAYk/U0RZjl02EsrCdPkAAn8
ylCMrCAhTlQLlzZexaXZeD2NMm0P+KWHP95sESldifB0D4OQFgZLhzgTz6tUUxvRK1B8j2z3pqi4
BFTgrFhZdYNiybKfSqCbYhw+dmxnSPLdcXfN2hSV4XaX/6I0zEKxai7jj0NYFgWVERjRBQS+1yyw
V7JJN8PuxdQTbKaYS0PBwn5cF3Duo8OCzaVfsbOZLtHtPvLdGNwlufunxK749nxkd0NbeQXJtApW
MddxmmxNWVOUFeT5faDXY2soIfMgUUbO0v0UMiFHLB3cuU1bxINNPMyEF/8fCqghMq+Lz0KaNTX8
g2gF7ZIP1GkC4bErBT6UFCRL5Zthm3O90GaGwvk0fTdlUnR+kpnIWwv5EscGK+Hw552Y1v7hDpwr
Le2h52/KIlqXuDpH42Vz6D7bP3xP/tBSSOmA/k36S936UzX3uMzY1+0I7PE9txgf3dIOqsTQlvxF
wfDrNgtqLbq833yJxhdsjv/HssWkWJOrVFhGL0ByUTjr7et95rjNqOdJmaoEwnbvtQgoz0+mK40x
Mi/N95vyqtvl9AIQfqH34pX+BxUmtmzxHxNd2xCX3HeU6v6tiAJEzl+GJg+G68/UtEOQrXdmd6gj
1oD1OaSkObUiTDQMRQF0fd09uZ8wc+F4IBG0cSc3kQQo5WtUqcl04/y+9UfhJFrvKUq1YoAcTC9N
TfSZlnZEv1vO0UruDJjnkN3XumfMVJtfSnOP7Qvhchv5VJ78LXjj/ZC9UOAkOEtQe4gup+aQpFBX
OuaCzVHHUfIi0/iJO2yTAxhbZu4J4zbt4K2T/0I/il4JeLAXgP3rcHAdPga1TL8htkS/5e97ne06
5I+2PEQG8jw/05EB/hhTXbYsJV+SXqTMTWeT+PhNn/py1QvJTDvUlpxNJlmsNbzA9vl0s1V2QlNq
oUltHGTOhiPDa6e2VI9+7yxlQpLzgpV5GiJgvYm5mfG+SApbS4DwodcsFy4gtPRMDculYDZpAJDe
ZcQE5I/EHWa82K0+azH3JQpzBX1P/5EpvD6klLOchYyISgdRqeHPKEGHBixVhYZRW5kA9OREgrvE
7/L0AsBlZGLJD9XuwgXVwyDsJ/MrS/F5hU9juhb3+iRdGlX9kemkIGLWmOPLuRGxT3zTsJKF94tL
LGB7yfvjSM/oqOorpKnwS/ZowTPWrL06eApF2PDHJE1Yc2YyrRIrA3QH3zPPN4wWRJkZhIHwHSAG
NHSYaIr5KVptPSkaej/F+h/EutnHkN6N+4ff4KxFJF5xKQYPmIrgsMTrV9tf0vdeXnHjyda/JUhQ
OGEPKTZDwgl6Ntyy/Crc2djgdgSl9NNH0E7nX8hdluT8yeuuaZbvJfEHkL7YIFZHy5CPWZrCeO2t
Fn9aIwTRiYTz9VRUgJ97OvIDpOMn4XYvxbC3FD8zpV/MW46GNRhA911sou6mEwd3GKudbXj20ZdR
RRiOCJVmkhZ5meNXsDgxFn5STpwbTvrQ2w+b0xUsZ1t3+X7sC0PIHaJGpW0GtlOreSq/fkpNH+BH
ljrHRJwSR7sSgR02Vfec3INSmhYC9Oe3RwyAiC5LPpcBgmam2QOXlEr6kTh1A1VHE2Z2YrPM960h
trta99f3Bvm415+XvTZWwK9nvsk0+HNLuszaakSOhMcxuSGrqsAofdJapLjd+S2yV91obdQ7bBuC
kkLCk/xGEgwP/twVH1PDu9pq2RMrrt1qv1Nml1l9dgMmQDSYGSclYeo5Xd5fDPlogDHhrbDbNV1R
dWpmgmkMd8aeN0GwTvF6htetFsQ4JSgsHCNcZXZl3/iKwxWfm1R0mMcVPZlwHkHnZoCMWYdTpcI8
42g9A0AkOV//rHjBVywTqejqvYkURqaQomc/xclpwIMJOTpJRhFc/yWGAiNwYFpdK7um1FEMlOud
UPN9iU5czPnYcuNKHfu9SMTp+4RsXj8JF6s2imoKCkIWTQq3P6MOVlOu5E7Z0Hr0LgramaLyQ+Qb
piFfuPZTnL2kqkhYkLrbWYmOiEKHiD2kABXkyQYjogz4Mus8XB3x6vYCLmt4bmsjuLtTii8VnJMQ
O3UT2wHsTSqLHnO990IVggg1lYxi6sKpbztrB4wurl0Ll2FXu6CHC4qmXUxhdsY283eAim5705EP
ccA+h4w+8gbk1/6hTOVbsz3vCzxQxvHscZHnUBETLAC6fJ1jioH6uNuiyLmkgFwlSL3Ff3N4LSg4
cCwpSfTVYHe65eIabGrygeHm+x9OmBYs3T2iA0vwHoBVeQ7EEGDPRlkoGtKE70xRsHBxADFcmKHp
waO5BS1Qt3QVaFW50DP1aoul9xxVA5H/7BtoqnEP6Yc2Zb74Ts/0xVg8KeLr2HidmmUXmgby3nLf
rQ+EjEeiXsdO89ii1hhhY5sY/fyo2VYTeSyIs8zkpPnMUuQiQ9flePTl9CMvQxd8mlguZQNL/oOE
uUbOSFes80gV7b3zNxvV4yRkfy+LEnHGVskmqCfqOycD/lgTCZW/6vhIsmEx3uQ6NJoi4Zv35ZAv
WkIrvrxB4lV17090V93x9dDrFmCPZobguiUfKCWXzJ9C2NKGj5aarKBqEc0Dx0+SycPTrsBs/tdv
NH3vTdK7WKayEp0+41lOvGMqjpx/7HIiO1AuLRRRLO82NXurvP5e2/A40Jatm/be4HxbMPVp6mLM
8JQpeqFlYsQ1WVnPZK3u1HEigq1WPcr9y9ZGU8wEwRgOZiUSpywd6lAYOhSIXAHO6s9YJ4zeJth0
IuzWB0QAr8raZV4VwwPYyRlcI9tfT3hqnSElVgwCTCP5jUVxgLELc0kU/Av9TYJwMd9OaoU7joiQ
KCzqOuGK6purjrz3/UXfMkzydFO4J9P7KH52O79ACird663r/aTox6l8FUeCBdNHgfV7BPIokQIQ
87CqgfP3JcHwf8Pk46+yPT7dON+Tdo2ZSYl3Tcr7he1PTJNTajrrz9teBKfiD45AOIuAMHRAmN0m
eFsho++Tfda6ocRqMpcItlrHuThuqgAuE14TY+1k5Nh2kWq7hdr/jbMkeE16cIsoSQ4VbYgn1fvc
EG4VsQBga9p/e8eYSH1WpOy87nhrlRwqyj6DfQWtyjImj16FqSfDgeOxsaQhdBEpewjEJOi+2FBd
DaBSypktFhBXmrQJJOvXq9LubKhuhJH2nRuL+v9wFY1UvQaFN8J8Sbxe3Tja+SIqIbE5wL6Q/L+V
swiLFHx+lNv8lZ6i4JHc68ev4NO6/ubo1Bh/om1WrBXr9Jvmw42FaNwcgWvKC0SwcCmv9uz//tWe
HLuZtz31pxnYbhwpD/H5JVpnbSwXipiixvvBahGyyC33znqkGudiOTWl0HIJlO9oolcS/XOE8yIL
jvbKIcTIoIaH7Hbi0M59sLTljQLVToDHxgMBOwcHkd6KhWtQaZr0a2GQNZvxaDqvSPS/2m1YjTe5
hf0TODBmhWsSOem9G9ete6sa2AvkYxPuJOykxOBypxbW9QPi95jN9vHSFiP+p13+NF22niTO7VOG
k0xmr5dgfaIck5/AaOvHoZ+ohO8CzbkAyAKB4BoLakKw7zAQqNW2fL95KgRgtGlEencMDYgw74EK
XRoWgEtR8LniD0x+ktZrGN7T4kqn+Z1rSvp8Nvz+YETWG8EgJBAKk746un3h74NiCNmu7R3gHY3D
hnGBEGPdHUn4lHhlMwXPUiBgCvF4Os7J6Xc+XpFwBTDsUcw6S2LTzJU7pRlGeG6EOHw0YdWNPiL/
ubCvofqwt+B/b3BIn11GmmB4rUYHZSygM/6sWz1urp+ZVveAuxpVPhgn9vFX/H7AmZYL0Emupdvd
235/aMBAxgXKPENTrlDxnE7CCePfxvKccXaTCXpBsx9EaqegZZgRV1yG8YZj57P+YNMeu5jWORbu
uc7pYdHA+TDGk0dTXxvcVHUaGNyB8aqXWa6ZHzlGelZulNss1f0de2TQ6wjIZ8xLLuc2FIJXiy6b
kiJkrYHFoC5UKfZV1dxHsv2C3Pf6D2FMBCzEDmaUAq87oRNUPnjAMAbjUt6tkxupSYq6c5iLO9hC
gp3O4EKFrAckLTpvx6kKf0qBGUz5WPwft8mClMR1MDDejjQ0vSaZHI3BK7yyFWIAk9NeqcbJA6yo
Uj8FAhuGsh2cFsnJdU+ejn/ljdF/nUgXqjo/22NRdNlpZLEGtXWezqC2Adfhv189P82SzV6kqLv3
nBsS22LA4rUxEAhnOR2Dj7BEsyt2Rqt63Vzaq6OBjGWbfbqrJfr6cQMd0oH2UZihy92I7j6zHfvk
8XmGDOfDP5ssXQd4OhwWwmLPDJU5VdiDrz1yDt/yBmVzz0GwwElHlqDPmMJ+N87cTAeebDAgybut
lHVHBBG1FujwJdAjN+igPXwngKbAP4Cumtmnjv9MG2GzWcMa63G4LasiLfgY9ApgF29h32jLHx5m
97jrV8sci/2lhK2YSYrG3KAvBSgfISYz8vJg3xN4t8fqTuD7pKat/8KoAwpN4/9JLZhOTKF9iXWz
D3GqNwLXF4MIowFhDuX8dBfDEGiHup5IdfWG0qsu8kl7AaCWu2xswOnG24IFeN0OSZsxKr378/DH
qnYDkoEpDXT4ewwfvBjT5FSGQ170iZyy2z4L1coC+y9+6KlFBwxUqhC44Gige32Tk2t2jQTnbk//
HQ5LLm2A3D/K/IPCjAm3BtRjiZ0ubUQSggaM8Jb78OaTdlojsJYf8Om3OW7XXfV9Ycc8lQYLu4Z6
ddj6lFSJk4QcDBoDYPqHqVSqkPiactGxqNlNd9bisCip7LHVqDOOuPtfn0XkoG8i08u4n53peXWW
Ff5dd45S40nWJMQJm/WdtmsjhlIC0Q9wxypasjKNNQjgImRTw/uMk7OLsIXV9pa4HPy/20W4NuGK
mPGoV+gIti5dm4DCYRjMrmPXPIZHZkn49+3V/ZPpVroEKbmXjtmm2bzyqipAssTMW+f/vld2QrwX
j3gTT9CrU6H4VyWmENylaGrkXppLpgL2aH3mkoJlzOrVXFWSkacnEnoNSSm2AVJCdvAsVreguZJh
GLnrGyu87oVX1SsjBE9LT3oELu/ax6tSpJbzPNUIXeTpMatSG9yJbe7jmlJFDX2Iyv6sO97VBOQi
MObgQ0WSjk/UnQOXs5hBc3KhqrmqJyFGDT44diMQvASP0s6rJB3LalIaU17GtpzOR1X0Uali385e
rjhee7QT6X0R3MwNBRh0Sers+u6vaqypr84pAb0ZNZcLMY7FtncQwHRujyBYW9Yp1pfIcOyDs7j1
ZzqWWmoMcSQG7aDR6nRy+k74rTXuBItiiz76W9YWiQWZO1QODDUq34p1ECNkb0zEnxfxZAsbiclM
Y70AvuqZ6uXuE1WWX30B0fspz1ACEgnSmZCWLpCdPr0et+HkbVvIUChJik/nIKPOgW9MZmyx0/zK
mTetmt0Jt+Y2mfLJjtTCW4wQTaz9Uj13SIYhuWNorTEZaM0saks9IagdkWgIrNe4wdrVSFDSb9wo
bgLugNfet0JMEtTKihgrVki8xolzjPZJU8llMqDVUP4Wm1Y8CCKWjpUDOBJeACtnCIZRXVFrl5Pg
9vlAXMtqxIZz+lzuNnCId2/vQLlRN6/WeOtWmKskku/q5KfixULx7+LRF6+2qEo/C+tGFHAFod2g
yRS/CMZ0nyhjmAozJJM90uRQyEm+fOAiMx90oITtSA9AZUVgxdkWkvGxOz4ObsW+1C8sNzDCPvlr
cp5gSnN/FrB2xs/cnncPZ4Dv8pgMhqhNXSs6YFcH5CDQ3j/IULPir+AaybdsygKQfREoPcN0gqT2
QnC+aLJpZblGozSIwZR69zZjqi3ULit+jH2xKsOhgpblHc/fF+Xq8U8Ka7zNZG9iRA5dw7bI6u0+
+6XievchVGv+iPH8SuK116sbRoHIfGaYIcgZvy5NBQPmpNWHYtu+S9WY4FycP0Qif4gEzl/XZvRu
q0KzYiwSV15S1Ctk7TGKBBAk+bF6ZO8Et/Mnyhb32xOuFY7NdeSxU1AaWYtmMuv17JzcUNzonULq
diLnUTYSVkBFZFIrRuaVmfps7GUtjOR24YJJ3NhuP6Q0XcuBYeUkjkPHCnXyzo/kVIUHcREwr+h2
ImDYG4szI+LAEKWSO+NVb4jtueF3ziCIgHYhpUfUdxXC9ltougCKQz33X4+z2tj/ErolYeaJQXyr
7cxJjpEcWG89pZrW3b47OCSyopc2G0tpmT+R5jIFwTJv49u8Cmk5cO26ICoVhqd/9x67jt0d18j/
ELJJ9WLnK8SI49RJ/i8=
`pragma protect end_protected
