// reset_main.v

// Generated using ACDS version 21.3 170

`timescale 1 ps / 1 ps
module reset_main (
		input  wire  in_reset,  //  in_reset.reset
		output wire  out_reset  // out_reset.reset
	);

	assign out_reset = in_reset;

endmodule
