`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
UNXM1C7NiyNTDTsiMIg9Rm2x0imsJtN5ayba4/Tuf7YJ0kU/7OX+kq2ZC8I74/Sc
duQKqq4xb4Am5Wn869eYhb1euvxl12KCt9bvjQPnzjzHhvnOEfqT0UL2sNdzjUyu
omEn6dTP3Jpkbr9FS/RVQeqNQFb9aVg2sApJI6oGMus=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 10528), data_block
hh/L4cQBhL/nHk5h0C9nZItR91ofMuhknT5lPp6LnDy9m6TYVBpap5ejI6Tol8yM
WLHLzSPx/+eS/Hiq9cOHXNPUXnp/VeJKZ9PEv6mgXoL6aQLsa/PCjXG16xUS/xqo
KqirJLlKc0CpXxNPcQ9BD5xl00H1yMg9QGSv0Fu2u6dHRziTNmcmFuG5mD9Q+VGX
lV7lG/ngHUYFLDsymrXx79vHz+/2UPdZL5lsG2v1yRVk6uCorgFmxM0TWlg+bdcI
b1hUZFGyqaxZ1HAhgI3tC6Fp51yvtO9QAkqV1a19pG5+1UcReaELFX5gHLAs2uJq
z1FatM/EgBezC6T/0jj2A3SuNe431cuUWD8JbcS91WcD9avhN64L1mnf8+SfEjwB
hVS1UtrYjUuBMAlijH+TPf1WRrwYcCmyuP4TRRAbPzSFHico9ITFFdGFl92LKtH0
0//pbfaZPD+j0z8dJoTDiFG49yq+bbBb7810cWWMCTbpRe+VB411EhwG5nxhxWtH
D2qYCpBqDKJRrs20hxBPW2wTgy9YVrshRV2nIjmE4R4V6lLbZzGtKdWkGZ6YTxnX
kPl0R09iIUlRNNyolC6Wl7eHv7hZGRSUPnJHWqW10iyUMBb4OfUrdlDS4WOW5UVJ
5O9Vu/F5DHYJhV8MOv0iYOGdsqfGhz4oc4/h63K1ECrEsEluAZeeyKLO/mtLjICr
CUNO4WlHs0QzEjrwwTpXVTVPe51a9n5E/fKAS5QMMc7/3R0kvPur0sKiTnz2a2Mz
RN1sCuKyqj7RoSOqna+UWqHZEdDgJtc8U7/ENgrc9YfS7ITmRQKW/tEpkMoGC1dB
RQE9bQO8UVTic+/pC6wTheQVb7f5pU/Qpd9Nzmg1ZogYAeo8+9ZSuDCFoK6ZOvli
dlviE2JV6a5nqEln0XYChLXaX57PPeg39N2xwhKPYQ+W/4EPv9ye42NK0hsNFOKX
JoTmQs2ex1qqOyl6gHYulCbGoUPlLBdUEhycQTpcr0dlgZXMf1BXMkDJhbjL7AKk
badVnMWEB6ziv6y0uhuvjD7XNh6tu7ze/erZLict4SA716VjKaJmmdnTWYixcHQS
/ucdgI663T3gnSuQqXB+eWSzXlQXwyO1FNSP/UuMPQqEELTVXhC5zP6vtTauC8sX
XTGQ3dtp/bs4ryCeHsusvMgJEEfixM5hp3PuZ8d8vPLDZMWK0107DNcl8UCH9uAJ
GBpy06KwJ/TNYioT7dtbYvGR9kBS+48vkyqJPxT/OJlbt/WHwJTF6QisPTzXSWMH
YAL+PhQleibCDJknVUlefVDskPPr3fzxyNDjJ4k5kDSXtjnmV56k4KujU9kiqUCT
2liEHP9yszuSuHsIESOPeH/6wqHsqLs+ptzEF+4Rusi4DSS85qPE22lUlp4Z2MBQ
It4CQZ056PeZcxBCAa+k02QkEwQr0GcwFMLKGqePHliKssrD2+2XKf9Enaon9VQo
cQz7Ime2eAKhJF6gcbZkHVcXq9J7afYeXbn1biNFEOHULUYRwwNTpgLqipTT5Cz8
rYn3ljuSdHzw/mzXZsBaSuxHEntOt9tZFnaVuT1SPEaueyncziQbEKHihvxDwigi
Zw7uC/1/9yoCEWpR7JrMhzCkzjtwZzUi9dq84MgULLDy4pgpzKpVTfNsJWVpqhfp
PjB3qIJpMR9ZRxJkgS2iAbv8s7vJHz8H/dN3kguut6CxdfPyiDSTKYEoJWd02Zf/
bqQ2cdwF5f5TJ2b7iqvk1VpUdbw9zCsu4DBWQRlsq7YWozjHB1t1gOgG23Dl7Maq
BkOZKtkpvEdnis4yxFhdfMPJj9iyXb0CIBCVyvoWevFs5xLKDv6WWd7/j68KURXU
u3diRqmb7HjWiP5hpg7Oqbyt7O3MdhN1npUXNaqyhzvBSd1ErPhvxGMZpnPzfrej
dtSq+8gsvJXKNB7KYpehtg3eBxKLixfPu2RiLNkj4VSXJ5qSLx5gZXFvLMfgZk7f
JRKXkB9yBMjGyIBnqJEtcZq/5AYtQD7PTr+o47AyhyVqUYK4+3krA+PGiGoMgpdO
EXJ0gMw9Rll+LZbsaP2EpFtzWxNkaQvSFEDR7PPPNOUfhcNsoJGpuizPrQomSaU1
N/f6TEEBkVCxLFM5p49nqbU3caCBmN9wx/QczE9JA+9/EYHXwiVe9iGHQ6gDdw0W
EplDYP7WxplYT7xyVUFlvsYtSlCt7QTIvUbWox74QlGd9Nq2pBkmB2FmoCYCRk1v
HcUrwXOm7nEKiIpdL/KgcX62TopxLzF0wie1zgVhgIuPHnKdPGmGtLbwID7sj4FQ
YPZwhEVZztGIEpedtXRDxrCspYqLqOghFoTZiorUxrphOHL1TAMl6UXtsT4vZpMW
EAdb1uiIm3T1Rtn8mljCKlUxXOcFTo7n7tgMWpArbj2qD9j9K9zymVHGdiJD63C1
uOVZ/7YxBtcmMt/w/yAOyuJSpnn3mbMoev07dHc1inlekpkLc1eaWg+tRi3cLRIn
Md0RkuJ1R3aAcCRqc/iwlMV+mu4HZoFPdI43TI+As509gJlDAZPzj0shomNK9tk1
OLq0LB+NdGFSbvFWbkRsrnTI1s6OMxb42gvjrmSvAz27S1ZfY7PI7MfURF3Eisus
IoGZx4Py5vA5FKQGpfAk//0YcLE7THDK2DWbm/HhsWiaznKD3pksNRiyZ/AhR/OB
0LGGFFFni/t+K/FnjsuUVYfvMCFLkxKcu3gJEm0mMyf/aULXOP18pDuefuHb4X3X
uiCaA+e+Q7v2bfmgDH7JEFzTD3aWAoiRvKEPKksI2OqauKzkTvuGgPUAqjy7myiW
U/ZtilAVnVB16vjamJb3YFgEgvhHOJzX6/RbihdKieSxQjCXq8f+sk1zXXJaMjhr
HthHhXO+ZQcbQ7gwllx9SVIre+UJkyCHvX1cxV4ntGBW43wuyF4nNTUoUbBePmNp
B/L2GbM0bVAZB84YuoSK/xRCGcjngK3WFZ3rx9nTE5HP+PC/AqNzwz/SSEbrRAHr
JVdFu1iFo26V2c41ZtM+japrU6lR9W3pVgEN3sQGd+aIKB5p2JdBDIj88HozXaDz
tqGg61f1Z+1bIuumOASK/QuKdTPo34OtvcLvrwVbNDis8kz4/hJxUpBfL//Qtn/m
TdTR8SG3jjOzaA2rp/k2fEA95XkBRkCqMgXkIZylamx0fFR956TkddvOYvYW/Efe
l2ifSA8fftFMZhzHIFbPB5sfBi7MHFrcv8FYC9eeNOv5bVFffGHoj+tpAVBXvDnb
8oFtcVP3X4Nwi7ofuNIMnN3ap0tkbv6p3E4f9viA5x7T/+jIbDFWMOuwRPhU4tbZ
Nuj3LhRZhgFnkVPX2Pz55nJq4fKQ8tyk7R/H8B6+BuLkZXzXPEIgIJRdBwzt/BD/
UA2ZZEi00DknT6vVq5suDRE0s/1pC5fEcBTC5HY/qQYruGFQ3VcXJtRFP5uNvUTB
XSkE+YJlQ17DfRCRm0D7APIKcScD1YEniXhGp5HGhon2lzD/8hqiyqQ1+JJGsY+P
XrSD4uwa3AAftn9Wa8i8qzzb+1UezhHjmUM67BGcMXawNb7fsHByCq3fcwsF8aBz
4HPcajUeBIN0qCZLSnkFQ8mSnhwTKRZC/+JQs+2ukqCfyi41DOkBzS0FczfKA3ej
Y3VtzLkgkQw29V4n9viRIjYl1hOwTWTilsGLhD3JPcNka6CPThDoZQe0W5R8yKhA
Qz3bDhfLeoz/Y9vxquu7fOhJwMNB8zeK8efXUT7aKC0ZJGNMcC7sZ51mS0LMGJGR
+4lLA8Mp5BqMmkxD4auQb9l6nvrQ5cERcA1AMTkRG4a1iT9upBn3RwV4CLMYNweE
svM1r7Bo/y/TxFeQ+PmqoJbF++kht5GXbMqaLLwRxa7dFn/NYlaDP7dTUUQLpi9E
t3DgaGrxbxRiAlyz/vhGF2k9QIsId85e7q/ONv+TQlpuehmrH0yEeB28m6QVFUic
v953wNYIQb1zUCDBaY4dl0CIpyuFuAHYn4Uin+PCxYKxVOWtr/BMBwL3PkADq9zI
mGR74+C3BXv5IzC+u7Zll5NhCvl5YOwHa301V3dXjM6TiMmtTp4kudHtLT17MA5o
GbUwb66fZTe9Nwk+KKDUis0JkWamsvxFszc9hr0va9Om7LxnA3JBap1GGGytHW4m
YpxMr/JdDk64KJE7ALW96dxUH/j5C658O1KJ6I5VgMq8FEMSQfw33pTD5h+91VpR
tquhZX5ny8p1RMgyFjS7eUEPShd9e1rTwH+3msZsWSeTpk15/H8/4fW+6bai8w8O
LBVraLaXNrtOS8XEA2z9pLuaCnrprD1cdUnP4Sd6xXCnHXLx8o8H801VLh9AmnZy
QP/LCwdFLzDNAebP+ABa0eFnjnZaRu77hzEDCpUObGVz09ej78e8i3Tdymw8rDhJ
F54Surszui1sK6lvy/+jDQmr8jZ+bM4n+6NNUCtIhaurK6mBMVQDxlSpi1hOuoqt
NWiYwdk5QV+6uc3GX61U2GDGpFUVBCELPdR/8MNXS1p3yRD9QQVONlt662557fyN
Mw/NkOSnkLFRS3FJzF4v7hguQEzbDiuvQLelPC4BpNvgS2yhU7TBM553a1iJZpcg
RT7kRTi2FvXM2zfFLpRBSvuF7Bgq9fg9+YzMHrbFxdFAGpRhRySTePikYl92Zatg
eg67tz6OanxrsYAEBWdjU7RGfoLdIw/6yJ/YGnS+D0RuXKAcQNG7NtdlNwM4g5ih
MjSbbRZx8SlkcEbPsiN+a3H0O2kmjPe/aClYeTcdAtFgejaql14Ap4N7blSk4ewv
Jn3eL/FsQMGSqsF5/Dh0tsnYhoCEAk4VbJT9FhTQayz2HpILXb2UefamDQ9e9fj4
EwCG6XDsr/9Fg80oAk/szbQuG+/o3sHM7dvGzTlnVm08tBp40jm0yQibvuUyCBLe
wTa0qGmohK7Q03QvOUDrSeRHIU17pfeCaCg93TC8h9e/Ct/48e64Zx/gZZwLVqMD
y+zptr8ZRgmUlz/uqJGMQAOIIfczP+/4iS7Ed57Fl3ptQb7miHNA9AbbCK0dHpFo
Z7ve3RMhN9foFciWpdVYhptshdNuDAizOXTpSlEs0I+tLfvX3X7EMR+GiZUIE9Jj
vAp8JMMM2O7ZaUHNtVx6QeFXFnP3CbytI9E+qcXwYciMbbvPw6iJ/3WHkV6UGMYd
lNEB6n90UtXvtYeuQ76S8pjkmNgcUdKhgNQLKGIqi7MwQOkYQ/6IoWzC2VZzL2i4
TYsWTErnfsTStSV+4JhpBM6w9ZN7Oo/woQErnCHsToIk9Nl2nI8x8PNaTvqeY+6X
nwdgWLMPN5ip0vYrtx5iiwGkCxkjWU4FSTuE+cpJ9TdsJe4Ec6FY8bFoBvlN0Tm5
7TpkLry8NfKxF+zsHfqm4D+lw1QOoVsQwPazyVDxCWTFVCYcxlwUxPsrPvEoCUOh
5jVTm6VM2y1swEhM5M+e2fSrVn8GsLDRZQn8z0N1yP4Gi8HPWGnnmjELysDHqrVT
4KAEyQ5HxnLzoOiDh7oCiVkKPU4aZmSS0G4k1ArVZRs70pfjuWZu8eivLuTVhEAL
J18J9KZxg59no0sP1gi4FAM4bN1REIDm9Ri2nGRKB0Ou3HMgWqFiwiRQJ1IXMxuO
xJUzh+xFMiGydhvbWYoz0LpgOzBUoUs6Rnj7QqP8fTfN8iqqtlNq9l9+yFInQKbV
J9SxLqmdITdya2yucnr7ByyZSPXVOtZqg05WQn2J8EapIzNzCGLrQuqGtmy8SLHJ
xb5LAJ3TWq5yw+qe5zO4CV1nICvkh7Du6Ij2pjghCApJM+t2n3f8F5zeuIg0opMW
i0Kys8zYOEzZ3Fia6OmswJ0zbIghAOeNVelzQEUQM3dDVxizQgTx4spsdWp/BexW
i/suRVISFzLRQe00dnSzLtO5vu6eNSDuL1WRAKlzU7OKgmKdlWzOn06lQYaibVz0
T6IBks5F30VPjENVZ4iHaV22xloAboTpXf+VSZRr0y3fsd9X+qG7QcTRhBhPBXD4
eH6lvGxJYMUFf/nFkMXYlBNizb8TEhxvMLnGANj76cl3adDs5/br3m51i2ch6mcR
9/MgxbKYWDJ6gL0DATbMElozfMK0j48OmNiUjKdsZv1eJ2hE7GGSQ3mpqbKwuAht
KEqaGnIusmd5rFJnDgStkXEthqu/WWLdMjWRusF0HapTm87P7DfhWt+OsXz+bDnp
Wan1fEx+iY17zKrNVw8Hds3PYjZLBLoX8WUsxNIH0yHlZnU/tiRWeAt6DZvWRZPw
hTMtfyck5GvIZtTt8vvrAEBa1dY458btjVojq+4mo9V5vK1fEEKwiERuhduNfusZ
yvCuSiKY7GjBhI+QWEJMTy3uaw7uWc2Dt7enRGASt5Ue/wSgHoJ6ojbdKEJs6P/d
5aZyaGj+pyK4x3vBXh0v1h5DpCXSE/lrK0/g2uU6oZCJUoBW4aESlNGCC9URtDDh
eOWPIXIBQjcsCKdpwwcDkHNbkrUAWULazohcSEQK4EllFScwnqQz2P07X3NMkjYf
4VDsTJzoOvffBQCPpfWtuGuQ5OLko6m+6Lj0S1Bq7Zih5N8i54iXHsIB41vGPx0Q
KOG5LxgEdOGkmrnsvujP4FcX2vKLKSdqgk4Y4cN45fZr/XbCg+duL4G0iDKnzA0e
iKUzSiUsaRNJQpUZoaBFx3+Q0IF8et+DoLvnPwphoSnq/O+zoty26uxbPrGoPEn7
gkQZnMsGqS866fJnHNwHB2tGepVoQsVZgp/UHHfuDnOAhlar+bKklzfjuPXiYM84
oqqKQFfRqWgdtZQaghd1PBMZWRBI2bBNShL3qTcjYyrgVAsRNLzAqrygqOYXQWjP
tY+vtsNudwC5jqO2Cry0NlNvcMEcl7+3yvFXhmsrsyuNeV7tA/oFSevfx+9EQjJH
HxTBOO2LxjqModHBjDQwOz5WIs1mOwrCJJlprCa6AxPHv+7AHe699xCS0pJLP8g5
BBLbLVySu+78Pl2gxZQxwukRbhd2XbNgT39jq+BovLGkKpGBpm3TT15TiDQqqttc
OffBkZusoYN9z4c4XMVfUQRAODGs9/8XFL6tYS+YtkA0R7leYgVbT9+NgCLBO2AD
HY56y+WV/uIHxNd6b+7m+eTzU4Aobfdq5CtC2ov4FmTTYVH+og1ePOm2Plit9dOT
xv80bauUalUnLY+odky5yIBE2zC8DRIJUHvtNoICq6ztr/4jTcXvoI6AM/LII3ow
SgmU+3R38TQ/58ZvSbGUStUpqMwlxE/Oi10eZaHdaVOWZINcZuu+ABlSSb/tlKuU
qbcXTj6errsbPWNizHMfs3Hmt2fL1ZDyH1M8GmCfFyB7mE4Puljje10S/O+VjOtD
SC5vzqzZ6XB9wuNwWqjMzpjPXJXz9o7CMirDBjnXmOGir96Xvy7WF0HD0SvLZgx0
2hvk6fDD3B1++qB18gc/3jZxKCVJtzK/8sOAfPhze0TOkhta9NfBQISxUMaPrVBU
LOVEB1WbVLEoPzWGgFW+wn+iSLQgaW5oiepJa+hDNl2ukou2V+Dzjd5WeVQlo+Oc
NMlNpRNKdNRYTgNlvzfeC/G4ET2S8OLtfqiZ0P9BhGWsknU0uUoFfkBjvPkZs74N
K8epVUmIFUN4sCR60gJuf5VeNbxGdkyZ7ISMa8h6t7zMpnD6QibyM7BFzc716cKh
1e66+pb8sW0lx4nETo6P/rsCTt8nS5UgNDAL8js7JT6UjeRvG6EuaDMj460EqZ3o
OMfI1YWv/B9aQeiszZ5KfvmAQUN7O5KFF9FOUKM6KuXKP6izpmV6qyleXJOywBx6
cJMLHyVuW5VPVtKuUKosHoxxrlShTY7JTsgzl5+el4BKhbpc5uCbJy3odN8s/KT/
r5wEPmQcEMqWcO9N/zt8bCErAzUkO1EXDZqZ72eCpwp60Jb5CDZJVr687Sz6rxpr
SAgFa4+mrIKZNWj+yBpmn7W5nimpZ73LqPJ1+1LyuZuCrRaUtQiNAiKrLhAoMm+s
x7G5JuiufZVrxcXQmDhbYFrY/0CQF5eM3yUcRSh/P9+BVyjLLqODkjsZ02/MgkZ8
zHHFf66pC2IC/dEAX7yZa8bDceS4x4WW1rAyA1rn6Q/g66MqHDMuybXeVl4OxKLX
3WGS/KNrAZFYVMS0IbnLU5IG5MHPI7mP7kCRnhFId36i9Z6+ngH0zf9w5zww3lkF
ypFrolENmOEs7RalgnmdCOpk4hi+Gh5Uh4bJq95y9yGLch3nh24YsemGcagEMrXu
xfnT4Vd5u3pP7k6jAHCuxbZgUBiQOuGe4JgHsQLGPRhvAcGnMLXWWbDv4sYnFFcg
0OWTz4c9BxklZI52JrbxwQyNm6mR6PazGYtEnsxH6F4cY2lbJmoNnWngBHmMaMli
HGz7HPlTnNxSY1ZPWsIyaoQdGZPnGEN81otG9gvMHv2Gfr01h+yqVqKMb01/sy/y
IpifoTBVBFKfqmVm8CoGN60ZCeB7KWzkWJ+9hOAvGlffFKu3xBafns2Dwsi7am7p
El8aM7YdGo6p17ypTrqrRW1TB94RnNOBOBNKAtu9m5tCL8IkFIdJDM3TkaK4kp1M
juQkyE6uF3pIaqAk1NaBPXNmGNL49DNgA3QF3sayQ9WnDw2JLDygScXUZxA/iEtP
ceDfsvhzhLx9+xDmZZiKFU4U95AuB8bGMQG7BAzEaBe9RPb/HLeCxbiy1++ixvT+
WsKzDdfP7aXEFDtaGAHpKHFny/OEBf0RNURADCr/uYNkoPDsMaTT6bqZAqc8IXJ2
luqQqrusTW7nNvFXfJi/gRv3Y7BvbVY9mzLlh0TE3r2Un0S5SMa3VWjfWgzunRhR
OVQFVPFQHwk8PT1SAd/RBJO4sAOW4niQGpcS9smag78N78bFW/EJzJ8uOnFErv/A
fGkGVxwmKhaq2kK3NCAmOOKrTWAU9ochZu2EJ+23KPqrHmi2VYLI0c4fD3laFcJb
JE18VPIyC1q9c2pOpjZL1lQaT7Skz5XQQMRWDgDpn4hJ8xQq05pE76g9Uu4gTAb3
nu2OxLU3+FevCQJOQcqNsPyOS+eS9hIU4pRMOP95DqJWMVgRyD+vXtHuNG8eE4I4
oWBb8fbfON4MjMY1EHxAAsO89vP9aqbV6WPzHXMcKym+QjWRB7e+R1cSp0InMTIa
8aurYeUGSA5aytRpnupULAovMWvoO8JKl1kLEWha2gYLYpzRPGjyJfQu+UysXHsn
rUFvsfwXq2WWUJuFt8TgSwAnHsCKDVjm/MgDG2cBJ0l5WX4PcG3hfiHCVsdziLnp
ktBRWzlLr+6N1+NF9lWlWFcq5Fg0K9lY2rB4K1LDZISWizANTZTwAkBMMpcNLg97
piOpLsm/yiaXt92y2JrCjzizYI6QF5upYZmXr3KfDHntMUP/ROrzF3oNGj+X22Uz
i9UcTRGs8OxExxu52CFkPDEND5xRm8FpURFESYg2uFkmmTOWRSuobYJ1p7LSMbAj
uRMNHJ48BDgJ/Y1xDtn66VO72yWdyyBaU4eqesyDHhxKloELnSDQeP5CQFwNoneR
2+zvHu/t/0c5+6nw44SMEUOcvs6HoXvm3CHR1AVpY4TopDXhMqTjY5BTzbmMSrBY
aMQvQX7OSjDQQ4PIB4H8Ti62YbI2cVDmBSloE3vNDEtXMFs9qos1PdR3gZIw1mpk
2pGCsGoMXk56Q9F6n9gUne+ab7N5UPJuwdx2GpQYy+VBh6oc/ed42Opvaw5lwg3s
TZNY2RfIDE19YMEVO1yqefHenfO7t2y/YUUnDXbBZJSN0iIYJOCruk0gDpsZAKDV
9af4bM3UVyhDvIlAYx1YVxY1jYE3iNauvslpvG9hnahTdn6fpZZI7CriuoZaYXGO
3QJAY0cIIpEoz2M0J8rRjyKhsKLfPzo/LESTtkUn3rKZyg/iFpct3pbJ/ayFZHoC
TCr68ubjnZ6uJt1iMIrnvWh47Zlno1/19XuGBifd+r82IeChUyzVW/YGN0C+hobZ
tYChEXmAf80ilj5S+T9sUKeRRiT5dbyz+lkFpz6q2cTwx3a7McRcBSAqhON1L8vh
O+iJTD+mW6Zsv68FUZkT7DKt/58AeZXod75HGzFUVVYlxO9aKi74/Qobc2TUrXLx
KMkybrynNZKqF/kkGdJbdBx6ay+oTOGXB9Qp7s4xy/oTlDC5tfXCcbFoV1g6Z9il
oVZMnLE6rTK1VQYeGvsC0qesO8UY96sDcb2oL8t4Rbe79I8Ly+zTe3y6mqeurAOD
3oOQ5t4ycCU1111Ytn5U9JuyyWBpznvHHUj2LF60lm5iRYfqvKAdn8HhwX/CuoIj
JuFfL+6WFQEYFV0NVZHDQhNiA+CjSmtLJ1nXzBKngFc3WBs8+jA30SHvlmPpCN1q
eaHUZdBrdQN3Sg7qdgbA/3RbcVD09lJIjDniFFnj3efmougwIqpwa+Vf/Txe6RZL
I6JxvwkNPDN83dSS8zUfze9hgbnA+1XJwkB017U1aICBl2RSgvHFE9CqWxOIpKpO
5+0VJOtjHY3ReM/bmN49IucW2fgKU5qYbRwXhzGodRwayMmPSlKgXWesAEQjqK50
bvAm8fK/2boEgHBLELzFFwfOoMxQga2PrKmMMnCjDapFhMy2nnY9P285YTjvGQpo
IWq4BgkRuIucEtibr/nEgC4A9uaUzFSzpgdKUCYj7BGRCgAInFWAERXc//tku2el
NZPTCX7QHNz4WYzlmODtK+0oQt4pbIg3LucQghp+lQrN3UrGcIS5+X/Q3xudgcLi
rk/xJu5FVOamho5HNXmiHN0vUWqWsPUGHN0eVk0XtQIZadVSgDxhhyCpIs1n0U+L
l0GUEDRNylShROQ1tWImVs36uno2hTXXwLytdPTOeaq28BbL7hGSFHuS+2SbecsV
lHL0v3z92+y5wmd6h1GqdyCKZ/y+YcZKLWqP8VopH5AiQQ+lIWWFr9k2+hWtHraW
ao6Cfo4X/eLiU+3AczTZ1t1eSwlMN/eh1IG6aK3v/Me9vAbcIKBorVX+SUbIBjPF
kWflCxfzCMJSEFwicYzAN4YPyD5jpZcOqBr1KdL9+w1ywXmVQDKb13v+f3KQQTCn
KpuvJNress5ErkZaA8MUiMSbHpCKkK1EyYhljESkpfCh/CHk3/h2VYxRdVcRAXHI
OHYINwA+7fqVwQd9f+MWuvMNrdFIAnjWUEwpIIan/ntVt/5x5k2fQkG6nSkVyqls
dhh89mt11HWf8tVtb7n87rMgI9jkXefhp8Ub9nDOc+TYyekyCkVL3mxssQqpYOBE
42njiie0ThxsIrWgcrlw5C2c7dZC1Zuh7Cvtv8Brgtoi7LE1yx0M13fP0PDGJ+yc
peFOF3O6qCVmun+bh395/DJ+IwQSwn0JgNlHS2cPXHD5Xi0DfeN9bngb6Yz+5W2r
wOMcOQf4EgPOjGj8/VnL5xCUPW8z8kzMCZhytc/Z6C9tn8uo2uk2WGC8mJs5fiHb
XB580KhnT8liZxJoFrY3RA9sXvOu/YOpW37FrnAnZ20P7uBQXkLLVMQs9dRG0r76
8jDoc7tYzWLMwlZlQjjtOui2Yg9/RKrlyDsCW66I5nQUqFlEC34INvGv5KoSsYbO
UwPyzEKJWqAFLbds7gUCHWVXmf101S5K9DfNcsZJM2huRfAcAehJQduDDhGIdbZB
m+GVrreuem8YEpfMv1D0vdhV/7/FEc0/8kkfk76PPxZaigWT1iDOvdrCLNfxDZQ/
2DuyS3RfrJXNnT5yEZV3oM41efrIW5NmM8kBPsptT7PusnjMwz7H+RbjohbuOJY4
59XFcQ7zfLbPZxsR+C8Njent8HU+g+LxujKjjE72rngT1H85U53NdKc3AX0T5sFH
5DByKYS6FAUaOua6jkOQePgnyrw54GZpNWpwagRqZW227c5PlZtZJC/aSIh2C0pY
/M+cFtQ0+62OkuMt6mcekKxWtYPLclochXiDmEFaOkX5h++UvG8Oc8CjimKGzcIo
B60QFfWwEP5bvTOjLIlnmTCu9qnhO7VVxpCg6lkgOHUR9CC1B5ebncWjG7+NT7es
uNIlfDLxYXQeRT7C4f2OPczj6/k30vdKn6Qr+Bdv3q6UVZQBptdxTdBmIFpHXeTq
xBVlmq04oFUesyX6QoP6Si2MBaxKzW35lNynwR53K4cGam3sGCh//EY8l7vrFUV8
0rbPA1O5nfOXkBvbkXZE2QjmIdEBfrE5GDdIXxaGBXPjxPCgJXveLv8EOX7FI28C
unflNF1rZ+67A58S1Y9t6u8sbFqd00snn2QumbvIGu+4593iUXPybGkqDJSwSuwn
1cb/PiOBs/JR18VmRf6KLhs4QX/tWcCtoWYxP3cpIDUL1rqQJqwnbLbdUvq6kbaP
/XMuZZXV66kEb6XC81ehcZ8fuFIxa+HobIdSq9DgoByXpsmmsDXL4nrugBfrxxut
NWBq/YIEAhpIC8HKFRqx8SOK2/tpmlTSuiTT6P9oIqzB0qs1+G8B/LPapZizsYha
MagvKvLn62MuV7AkWQcHoGugoJWca+YaeHQi0lwzP8mrKM/6CfDjVwoGfWwF7pE9
B3jy9tbKAyT4nz8e1mSapzCpW00TRPTPOzq2qC2Djj4ToAecHmnqQH0Grnk1uJ2A
OnHZKtUdRlFkYKA50pGLFQfwB/xu/HbBvlWQDPh2TT//VC8ddrWuXogqkkUi8KMq
JIAXwBIXHqEzi2iNY+jk+ketDWlLYJQLPj7GtS38z7h3yI42Tet6QuQFOZzEOV4b
NZM9IKTMs1QLAOi/rP9o1RsCObIuZDdwSJvXwVjKX4dBvCWbcAxIT+vtuXjwxg+r
yfoYNtj2LCknDyv3XG1gCWRXyj7HujvqzYT7lDpR3HYCsYjc2AECwf99/sitTS2U
GGGfD0B7DRFPc254+9D2UvpFSIexe7zJdXbBbbd8T/GzVktBKn9OfF/Ds6RcSttK
CXG0uTMi+brvcsbpaZagCZjSZcP8zi6NxIUabyVs+M62GGvIvgl9JqQ/Lc9qlgwC
JK7qaNfmIz1lOR3fYgJ1PhQGLlxSxz+5xukS6oxg5usfEL3SjVMg0W/QM2oYBQY2
NrMVJN6xREKPKtuPmlJrxMdVYOvvuxB81kJSOnavujp8w3pR3f9YRpgVuPe/3Kes
MpCrSVc5sWkJWLRG8FlnCS+ZI8YAzTBEZ6x/vSUqKMuhl+Gt0FYG75DINxYlDIAr
GbAL0fnDoQge1Z1b5jWDq5uYFjdXVnbGoZD9sy1lABBFvx+OKtSauLD40O+tEdCA
lX15MvGnPpNAVGj3lq0kj8HOATgzqnkMLFAwCiyMq6FjSloIgeb8je89WaD4QP3g
CZH4Fkg8SrCrDM7siaTljObEvxSnIv3WhdmPVugJK7VIuL5QZE/zw/fXR6l0v3Gc
P8jK+laXAImFTnoKUINQdp3l6Cod1yq4QPBr2LlGeHmVPwnJjHey+LeWX97koPlw
LgsQZfGD8fnYmKnmwsFn97HblWyGBuLsP0J0AKSFqzefnfiO68qgcD+Qnb3nz4Y6
OE/DqYYOWzmbSVyc3dMVQHpF6JrSVIIWgBkKJ0BHAsJbbiKQo2ndVjCKY2yo3vBM
tJr92dYsUoqSQ96pK5idpcO80/ekLsgYPKjJ7L0KCuoYF6pE+ThCu8T7XjKPrWi1
VPO7lLMh17uOjPwMXG2LmXSI1GI6x75tkpSD0EQxGhhkXKsOd5NNTsdZpcFUyEkG
zhZDWOVDxi4yhfaqaEiAeeMAOUZ9IAcqd2NPywr/avGJ3vw9wr53LCW1dcdQ20Cb
exjBcAjlajKiZ5GAj5/nwsnCoSnL4TiNoRAJWS+XWmesnEke8gFJkTgUJ23CFkKF
9Xiyi/S/VAMcf5Dbs+0QCPUd+cDtAMRyU2Xe6J3vNF+FmokgOKe/CBWNp2WZYEPD
IuegOD0NMB+y7Jz72K6SojbvZAtCFdwnDsta7Ske/Kr/V3M3aeqS4BFnCadS8aHV
mm5fOHf/1Cadzd1HQsSKzOvEXL0iweOU4ImP8trblCBc8JDCsRzER97UgyFhbRL5
87HSJnLe8CuAcBNlqR1Tzg==
`pragma protect end_protected
