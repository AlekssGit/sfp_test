`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "10.4d"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 128), key_block
YrulVpTRHNj1UIR+Fn+MMFojL8kcUyrhAwtD1sgxhhLceP8DqVFBXG3H6AmJ8loO
pYi/KK2wFoYvRv1D96h99lW25E4buTiMPbr4beyLzvCnMtLtMofGpW0pRV14ABwo
8ynvfR9YoZwd8V9lLtzmTWUC+AfJCf+E7ZY644JA7cU=
`pragma protect encoding = (enctype = "base64", line_length = 64, bytes = 31712), data_block
Z3nr/UdYykVL1DVWrKytFRWpEetZ1F53bSTxQTK7Qm5zvsTxRdxmNYJsJC/biIi1
nBq0IA8S/m7AfT5veO+ck+EmyFdLrx4pEZXyjs75ifWhRdd766w5ZmQKyT/dC+6P
B7KnPKdyCOy1nCZqxryDL2I7Fn5xm30O7RFf/uXbEHceb0/3dP38IE/efkgs/4nr
Dr6cmFIcy2UheDP7xVX/0hjvKkx1kA9eDYDG26FF0ncEEEA4+teHi8qSZmtqv70Y
naXxOk4cnhjRsbBaTYzg2xW9Lut+rPaC6iTvKcojwZhtC+wuaUCTeaoMMRJeIjym
GVkJEk+DyP/VUQztYasnChejTEm+kgf6luFS6pH6reFABB36e8jSNMjOQ1iwalBD
gTTzC0bRluTxWcjVrI5lPC1+zQAdau8zaXB7XG5NN+z7EUw4na0gaktWoEuw6yaS
CnFUblD7VEfqpQoQavAek9kjql/uw1AuaOnB4KdlY30LdP0AdlZD6LAk599Z+FjY
JlkgnAOdvzbAM/CmHJJ+x59xJPzRJLbORu+0QDfo5y5MzTYG/3C623UIthcMew63
d0U83FpA4THD9okrYTd+t62GiGF7nhZreuG/52Ed+KioGDuQHuD2kMdUeYA7Ez/s
qi39lvyPKCG4zg+A+QqvqV0KpS3Rr0J+gH5P1FgTGGZnJYbrKh2lnwpgw4zYGLuO
QoHQuRW7h7R4WRqWHxIO637a7LWH6qQ+UcVFJtKde57gfQF0Q0UF/uhziXynVcz6
/vmN95hiJNsTPen4vSjBZqJFdyp80274msGQBH21Ir3ObS5dHPw2eKMS2hCa89rr
0gWhKfx8fAvAh20DtM3cb7f0U6w05BZrotcVAjgt2oQVddS64djx/YvwTd6MvQe0
h+4hWS0hAPyQ4hlRzkk/8YvRElMZgCT/mnWt91ZgOpGXSzGxPUIQRzzfzSG9Z7kH
Lkca0Nqb+TxBf0tOvEWvdsM8orpoDA+sOdqAna7oBR2GIULNlN/xTDz7i9cMW8bI
iaQCpL5cy0G8Q8MB6R5fUB5icn3wKMxozAYOULJywgTmwMqBhi/mPMERA6+eIoNL
IuQo+0eNr6NwJxPyAu1F+UdTIbWII/1SXXtD9AfrX5TBEW2Rf8q1MSDVibQaK6XB
0d0Rqn2iK0Zbn1TxKHCnKx+TsZEdyYrMCt9rq8pFT0+J6ZJuC4glxxYuoD9irxpw
2rpFEku9dziSyDjm3leUhS3feced5F1BJqJU8a8ZPNAGd+Clol+kUkQ/eErtFOot
pFCzbQj0A7WNeHKrp4i98sBIVVQXJMn/dBj64UGYSqONLj97C5R1Ti1AoZSpJHZG
vx4qyTixaeoqlY2LuLEyn61VQWLNNog8YB3jJWKl+NFvCoqRD0U94TI0qsBQminj
aiBt9HA8SZZTx5Jsqwy+2D8Agfz2u8LAujqYQPR1dPk4sgzcxJbkdJHZf/4IPn8Z
j97ssdNbikcSPyHihEN93h82OPbRLS32f5jpVRlqhRvTg5AakNfz9o8R6azYtT8x
ihCHbe7IM+iFQh1Mia/yhD+E87NNvc1VO1OFA+Te7A3ck7dlg1ubMAM8sQOzmNcs
8awF/vPMK9IdaZvAqlrUJlbW+QQH4VqyfH6Jdo8I0SNP7nHGsYozxTuaNluvtDoC
41coR6i9nwu1ezWT3p8vGOV+P2T8ywIUTvHO0szKqnIiIzY2pMKVGUrmtOjB2uIm
QE0BUklpu+zY9jdkp6jauX6jyu6XBZW6Qhe/u+QRH8yfuVLNYlSLCXdceC/4qyRz
l6/yVNsOCgfYL3A25yHjZQwjXVdjTR9jPM+aVQ+0WHwr48GBuQiBIRQpR+8BH0jz
m8o9rlDV6CzySc1dls0VPyZijuL6n6KN+3pfod3AHb+a839v5CNo+HCrgqZ5MBuB
HHiefkIiNbkoBT9saFmRiLivQFGbBGqE0Ml9sHbXVjq/ZRx/VnecTbQmANE20XA1
+GRfxJxXSGe4DMZsZllbLUoD0QF5WmWoyWfvfB+8Zt08W2HTTVzSVuWrQvT1Kgye
TvCsOxzNnxMvEoXa5YDTItEztjFrD4+I974jFkbGrcJyK4ygEzHUV81H/n3sBy/e
I2tiWNDYM6wM3vtU84AQblh0Bm8K3UQnR781cZQzlcs8PCKrfSsOIZlSWlzljj0k
avcTnIYV//bfyQAcY35y3NVMd79EIt+iQiyale0zwSyIhePHVEjELZCbGhYiX2ZS
KEVDcmxWFzYGuVJryBk+Sd0n7clrl+1Cma7JF0mspoA8kv9uP26Z2ghO/236hTBK
VuZxRhppdA7hbIAvZ6I1hwEAKQJLnxeSW6/LcufqzVHzmNlIprS8s3Jr3usTusSE
So9j8y79kenavkIYKG6PUjKTiarIOmeUJ0ErBeXc7ke9GQ52+ABlstqVUj6BmgqD
RA9S/i/g4nFA00aXW3M7MFbdVi293aJoXcNM6QnytrOFCl/LzN5a53JfkktcM8hJ
iwiDhBHNnPPVLDzQ++NcdGFL17zJ9EkK30B12QI3hLjRJuxKdGameGfYOfvCK+OS
X+xyA8GXhT7BURKYXSz/AJCM06QeaUooq4Em/dNzURfdGtt8N/VmvlOd4wO9pvA/
9sYjMVU+75IQ5ZehgzO/fYrbNkNAwwA1rKvhhKF1sJcs0kg+nyh7kqTgPAmFUu6U
Q5rO+7eTKW65YUEjYIBYv6d6DQ4ASpwp0UeXkcYIIRvcpTEeMwg/Gxz8NOyd4fqA
R7nAHnxiYBEdIZXcXRXBdxuzoG3esQG8yO7f0Gfh9+s1w+EdIUBiGsiOBKg/+Mxi
6Yu8hR/ABJgmKuJYwg13SuhoRb7TEpQqYoBPpmLePeqAjWoWa45NvccVuhfTdxZE
Rrrj0NldMm9xTnt54Hy0QbhHWgEBew+s9JCA/Sj44G8drMZqZ4zBTVnS42NxUS16
P4LTsuR/PrCaw68UPNu4I4acTYb+6DM5rgSPERmuk1WNtX134d8akdBFq3Cch5H8
8uTftLz4wTn949IgEn8BvEsivWAs+66uX1P7XvpUMZyT0sxnpmuNUlCx0AZYq38C
YgO01RlhdN0DKLvVtZdkGtIrw68CMbuBpg/NtjTe5W7IJX6SX106V/MeDs5Ibjuo
WqwpWBR4zjDWroTY88Evp/ajLZYqfB2t4ApgqknZP453x+7+GH0QoNywcY2vwybb
TeQB8iDkKld9AZoxjlfpfHFHNErKQmVIYnBAKtZEmrbwgfVBfD8CngjLPS0/ldBQ
4EyAuHOHMxxZ4K7wstZ0Ugav4py6db2S1lGr7JZg8JdSYdQfQiOWwvnHF9HI9UC4
6hSQQXkb6+gvQ8TQIjxX/OO1vGfjD4T5hOs85a4sRa2enc9dcNAIoLeO9YkNggUh
8OKGmdmTQ5h0ZSwaO1DQwNo70XlWmyTKsTjFNwpCS5Dqg3Hk/pKAstx/iOkQ77jk
dm3TcdoJN7HDGkjRMUuqifqsJWrOIFnE+9xXpYJd9kiR4H4x8bv0103omBh/omnh
YM7Cui3+WlC/OQPUgyPZ23lvSWDSCBeu8Alt+gnacVEVhsoOjfqndFBAoRnC5zB2
xil7+k2h16qysd9Mp0Gw19H8DG1+VlFviiCe8M/XhwU5DQKKWTbtjTgpNEdlBLw5
q0zKT6I/Rvq4hR6XLIw0hrquS8W8rFQSvQom3gO4bKKJ0xoaaiMgwgiuicm8F+Bg
90zj3dOKF8NhTTsIv734P1rpIb5U67oqAwhbXjxRMcVbwtx7aqrVWcE5KWCZemyj
GjGn//4SlA5Gpw+WriJgde7TO8SRy+gaavVGaCIuNexXB/NI1nTG3mUVr/uMnePF
pCYGrwTN9CDAPnrgNsQ3Bbp7zVmPBYOKQjkYgSlI8pBdGKAqL2uRGW2f4hW5oZgo
Iz05tUAkQTWKlLBjwfpZVzoyxBWpIFOUnARp0Iw8JIghE8IWIw3ETBoo3/MDaUom
Mt+iEZkGAhS9GkesFpbEyabZjm7jo0EZLONhzftKIeiggdWMEVr98vl6p5eDmtoT
iHj31jGjGO9IURloONAD6y5b6FSoTykD0rzbalIiUheSdIitxG4I/vhhp7wFndSj
lyDBpm71c1Fpa4huffzlQWIfRVyh2sGGQB7xpaNEWTfPtFJ4pLznW3d1YGh18kW+
eJxSbks6vD0Vhq9kW7vqSJdAbLTF1xurYUVvrCHpqpcYvia+4bhpgh4F3Q3yWOwS
trr58CNIzP9hv725HTmgcvQOBHW4fswMVl0Pp3bZ8OZg2LtZivp/+dToNjAISUl2
xWCiGdgPJgW4OifxbhwXMoWqigbdNU3jL1QKMleQSPqzqz6ehVUwVlZvJJlq2iL/
qtOyqb+4/N7q0nwvBVLWZNG6PnM6NPXe0eZlHo/Jdu8tP6n2TOQn5OaFXAYr23ol
98DGJoMtC6gHf8rkcTGT+lOsaHJIIzQd0B7pEYRcNwtUiWS0Kg6B35D7JzMeGk5q
IaE03rSYu5wXHwSfo2Qqu3FkNjdQnsw4K2L9HC1PcJmnq8M1zbh8yT0Z/FdCTbIy
AnE0F7iLiU0rD2iHTBb01HdpvrR8WLCMRf+ic8T0UhkWu1kOJNbcKa/S1dBLN8QQ
mQAS5Rg56NTmJ4Yl+F7lpaSnGgn3cSmeaus+wNwoKA+6b/BbD3FfY/BjFG2OmQvA
eFEj3SHU5xxBvr3mjk3EJ1HANfSi7B1UBDJoiXTqRlDyieVo/Mq/KVpqkqUWcw0p
QQLxpkzegv8euRZqomaZX5b+wY03OHdMuonM6vsesglN4sLogz7rZHskuRtUEEVm
0thnssUw6VxUfVOsW/M876JZqqJkCXKi4sTlfVxijE3iu4WxPH2iJu/d884e+G7S
XizfUVSuUEa6GtDY8p0zlb8pNOpgQKq+YMIjJDcM54nNsSzUjFLCn2eTTDcR8/zO
3b4PFl3A4+pr+PaPrGef7zFZULsWV5bPr65/hlmQhbcVDTgXeS6UOleNdP2UndGJ
nFAkLWKKW38u3BxfIUKPd3d/5B+e/mK9ymsxcvH87ujnNhlDwY727wROmQr3sLOV
sn93e6ENLMvG3pIALMqG4f+2flJeW7W6cqTulrumlFdh/Lrmyx5Exgl8q+2wl3UG
NHb1baSCHL1UphJNXg0ucyRj4/KvO5q0ooB+T2SbQ5VSvgealarn4QyszwUBe5T8
Q0jTF5MdqfjKQMq/V8NG8wi215okd1xLm3e0mpyBk4zrDrlyzFhT3RTR6+bdkDow
3enaXi98N+gEtXkjs3+OMs5zqzNTAcOHnt8tmvwV+42wEZ1CmRfVIE6A8KPh25i4
LylgGTqv+KrKcIR8qX6GjnThERZ5cCpSgc/OfvsM+B8MoJooWjaLyxChfusK6orv
Kdd6caYT6O1EOEKT2JcIOTAmdhNhAaSrFugl49k6QZuwsvsDM0jjj/OOhvZ6c6HI
U0o21x/rC95QO7Ht9Zi+rFJrZpUi4rOEPAUZi8QE5kcGXyw2VF+TIQEaKur3Eh8+
eB2zUz/2X/ab0Or0OEgq8OrwC2njIJiusIzRpamZrwKc29GYAmG8dS8dty7QFJzr
2+Z/0euc6v//xBEhxg7hjDCmt8pNIUealLdIuB4FzKkVeXjJhlC0jMfjxYahsAAr
h0LMQ9CLYBx1b5lC5iyzHAoO8EoXBMu/DOBKxS9/6BWw1789mGqM82JWIQL96nK6
TPVFs8rtLPawRtmOfjx2p+QkRYuTOeLUoPN/yKN4eqcvKqUGfnbi0/hPfbU8rpfM
VW5M877X1NbXNizzws5XVbmgE4/ctnyUJdIMQyj809kmWfImdJKZrmN8wENYqLwu
kh1lmcJtquG7goPBlzHfc5v+uq7c1Lq55HjqKpWkOLeyGHC3VtZoUd+5StDfvxiP
i38nUJqZ2t1H9Iu9CGKKt5+oA+afkQcR7ICfty1MP5qcdyxd61CxL3gvAKarGGxU
lp3DpiUE3g52Le4T1TzrJvOxiabv2bGpYk4yHAknNt5xqiTmiI45zWSLu/ybcJku
yFRXw8LowmNMfJQ0+7s29KJleivBGNJaTNCTuPmCR3b3boM4kybjoNcslEdLW+t1
1k/hCCIKSax9xjXdgq8FZwE+2My7vOi85LcskaDcplTwIAAYW0eFNvIrbpBTviHY
GXESc4olQXOrlNKM8OWNtEbuCc136QHZYCYQFrfSV+UHmFvR0UPlqT053qC8Tg5F
SakUdeiVuBSqdBc6YMa8bridB20Lk9sFxDhFjbJPxApfA3yN4jX7fv8QxMhz0Cb5
PpdJYvN7wbz59Htfy0rpCLdGsv/c9zmeqG07MPkP6BJOeuiqXM634Nhq6XGDdFvI
hs9buyAKLW8IkWtKdahxhzoj1NDRC3CxnKDlCNh34BsDOrL4k+NuxngveHfNQR6V
xbasmGHgumxwapV4kjrE8RI3i1glzx5Rk6pGTr8B4NqI8vUZclPwyQOgMgNwgT7X
/lttCnqFcS5N1Pt18yf3VlcM39PUA9OsScSAf0PdqxSvkBKnqm5IY1Oc6ILOEyF/
l3VYtRxhmxSRHNn3tc8P6GlzZFlARIyoaXTXNlLHNXbBiqqgUNNn8USMCtNqZDEU
cyaTu/vTrV09/JHJwQbY1xzP35CjEKJ6Jir+7iiStS8wI3aWBjXys/Crd1isnaVo
Fim9PhMVwkLYDvzdZMxGtfL6SBdt/PRPrtSVcfViqeVxPw0AIxw4KJ50GODVXMqH
l7+KT+2EaxBxlz7VBY6nArVzTcz7ovUfGHyJ80r6XzUZ4W97xqOsCi4Bgag5IFQo
N52ZGF/fdVnZ14OBmz5Zp8M703Ej+BBCT8bUfBKaMZNgGMD3i1cCWxm1eIBgj0TW
QUWv1E3BgVvZwCwYsHz3uYb/8KhmJjlQQHTqZ4J7/5cuGylJflrJUF1Hr5HWRRBg
nHYHBVx28FhVPaAiwVl+/SLR1LKdauL8gy+REVSUSGZFQpZBzy8hAXdkb9KtCq/o
MOpSB0sS/tg/a9nEj88o1CE1bq9tlYEM9yLOkQMffVNK7jh/r0peq1FofS2ameBu
qel6/AEYXXaLoBm2zvML4eCGI0fRY8GP21NQ6298MkheqXKRe0HSH/5F1HdCsptZ
GdGnK/YV5YFSdJdVsRSvJtNRyYS8irNj/LgftkEFRQszNO9W/C/LP5LiKJV61GTW
+wljKoNC0+K2hutKj1Y3bkR9lubwmlxkcS6eHhOhhKDuA1iS67j7lKpMOYWdq0fC
0i0KHLWH5j9KvAuryIuZ70zyBkiGCRCqFknB6WCZ18O8l+3tO0sadUONmlaZZjNC
80jDtrmTHgRTx0nFendTZE81WrOeNcImWdp/j47OzkQ7zP5/CagyKxzVq8zp1fBh
D4wHS7j04B95/M+THbfP6BwNrXzq8bjsz7nXjo11+fGddJe9ztY6Hk0xh0NuKtEZ
3dw7XGmhEvCfp0qkmfld9UwR7Qits6/DBTwYLdyuFpMKhbCj7HsLyGyJVjKkpP92
vVhu0QHpJH6x6hM4SnDZK1UKugCfpKSn1ZX5ixlnTT9JU6DaM5zsPMdL6vYP4VMv
RmjdBmChNsVmwcuV1SGoRtVmRABofsucnQWBVG+8bdG2FfpZeDz+gjM06bqOwD9x
RJPqnCJDvycGlAXF/oT6j2gIzxQ2fr2aOjBSkjij1RGRi79hMKvFWP5jtTo7bbHz
O9KAvIlxHTWACiG6XS2bGEybVD8Q3a2IFwj5WuMBx5E/2jkGoLjywEOV+3HBa8Ra
dPpxUlvqTvGpvl7sxeW6lhyMu1qDdz6j0k1DQJUqrb6SdX/ywtery7tdwIPim1+v
1dtBlWZ0kXSViiQj6GYgdM62+YpBcyLhBwEAKpfZJMC5L7yRmh0cScJ4Us6cEx/q
1y2e2sgaSaR9BifQAE2YY0n+Z4PBSiqxuRdZvEP5WvUSX+/s1gRTyfp9s3sfIGfK
umP15EyREt2zzzMwznTexYAgjLjI2g36kh5LogaHeUNPegz9gGCa9Iaj12D5hR1J
NIB/XlRZidsyc7N5JEIQ5AMyOutX0XJXSI2H0uGOsRSgllPAkXuFFHJy0i+t8rB7
zNR27r3DpLm2mm5N4+b1jSWvEV11GB4DDwrjJP77tqUCnWbkAwm64tXHwcWxpq9R
c2B9gE60hSjBJEfUNyFPCwq24sZIy1D59Nyrpg4B/kVNfjcU9g+8FaE8VCqUtWPM
AE4gFtrmfUM0zIjckl5IQKDUONTfuxFlLxCIyNssYmo9MYiXptBrGaDq4wBW2/1D
2hLj+HWOuM1du4mArCaUl08EONIHCzoDX0sEkVeZPIYOot9WLHTWoIW5Pw9ecxww
MTcqhKNk6+T7kw1rJHlaY5i84BmDgZEiK11ucF03DmDWG7KY989DUfIMT4DOWKgx
oY9ycBP2aGJEgwYCAY6BlqA2zQ8Ll2CqyrWRgHpdELw4F2BoUy6tyk6fcmVpMAWQ
1a/JEWtwoAxQ8eTkS4BVu3lAaVYLqWXVil8DyN/c21568dKOUnTfF7n0nWyroCt+
DGoZB/OvyV96gmYB3Iili7CJlNKWUpr7Cftg5G1/DtYLIIyTO5FxsFptWBcQbn4W
Hx3+/NO7W2FzTvtS8z36K46AxJSjPjXM+42YE1QMxVIgPLTKi3tdurGQb6k4Wimb
3sesJeivJiytW5lUdxnI9w36oRu1vYfFt4WJp9UvHHjeCel9bZKyQudi5EIVVNRs
fP4VnU+4RLZcddmytz6n0cRsk45DL0swrFgdCPo1LsTLmOtz1quHx6HTFkKGscqP
v1tRsV+cbdj817urQqE8d9ff2KqEiKkq+gRedPdg5EAqxINhkasqpvj7P7sRPAkg
ff0ziMxSHba1yyRoyeqvJaPdW7/2Gggv30kbQ2SN4ZIjdsRm8dmylFj3hAUnF5xS
YzecnutCslTI8zhjXuaslaGtDrLsdqvbZDkJT6wgLasLE8f6baYxmYHdz2K04r5m
9555quJaVkz1uVOvmDRiMpmxCZlqPKS7QyJkIApkgX5gk5McPfqrO2knyo9Tebq0
pQqivLeQWtPDpU4vU7bBit6jTtwNHmd0mBolM+8jZYgtsok3skm4I8WDNdkzLT7g
+gzLVCQI4Avqxu/CEz3DvyIhJtGnWwPfOTwt/9wewk1/GYslKjHzLHYoE14/aysC
EKh1XU8bB58w2T8S3tqv7wMW1SDP/AXW5lphpaDb1rNTbJkxsH7U+MGyGYOdWKOz
VFoTSf4DtZZXH0DOgFh2KE/awbzyPpgWXRfzcSuEozKB9YxceKsnEbEeJroXQ+Kp
QAi87vr11qKCOpkoI/mWG5oC++ffozME6cHDE3pehHbsNgpuJK3QW1ub1VseWd+g
VmxcarDyOmwmA0m54mQYeOY9ehMHOm5mOWKm3xHtY+JYR5b1M5KwU1Zz1sYur+Ra
BsK+SEreYdkI7iJ/szNh5gWhNGVL5BqIkFF4Gxt7zLZGgXYCXyg/VGmaCsoiTaLu
0PQ5dnd4XQFhqVgbZQmd4c5hOdIJnHgFkMg2JydQW+RH/gF76Rv9ucNaehRGKo7N
74DFyBwZOjZwcAQfCHeWtbh+ZX4MGPTdJ4cQXUNSnhAzWLLyLDXPXgzPPcYSDHe5
Qzbgm/vcDuGjoHDjTK7iFip2yoRqZWIJILNdlC2v2r1NWrnv2A7v1Mc2ocKjgNTL
e/xgZ4pGNBnzKZlP6EI6+SymyjYwbKCC1dACn7RswSxarfdfgaqXuCANtN/bXpiC
qCmpv4YHDYH1u+utub/lAK4UO/93yme2UquU1JQIwD7sa96+9cPxolnoiQgGKeTM
W3n63dGkiHkRc+dqaaBb+Oqazs8eJlEuhi2ppLbHWaG3472zD5DnNSPFpiMe73dA
Ky28RvFMMt3cLcun8bfO8dmt/fzJGaZQAoDSphPPjxxxTZJKHjAd6Vg028MQjn9u
x8GUH6UBh2H+YUxcsut9MjT/g4qg431Irkk7J5cNDPrKbT1VeP4+vaGWWeachdoZ
50BBWEDyrZeN6OySZoq70KSBoxR0by9Jz7hb3s8rqfPMYwLvBJVLJB9Itmq7KGTJ
2p5mKwfOysB7GZH4i0KIU1AiwCywO/30KUZ1Iu4wPo5jgHNslhkf7j1qdjixH++7
NlEasL3/c6Cfy9cLee/KMcL9TizisUIyNDU+9fRwyMOvFmyjPpYcESahOeLVUJ4h
u/DBmAdWRQMx/xz/NoLZhI1V0kQaUx4FfZ8bnYe5G8y0wj0gI+NgSPX/Pl8UnbBY
IzVF/6YxkWZa/JJh80TEA0ClYed97xcNZPWKmF0sacUqWuwf8Ik2zM5N7ZABGhm+
L5w9l2YASZVHdcunvZVfaTdt4I1aRpV8YuP6lJl5cCMYmKb7H/1Hkeizdx08VdKd
VZSkMrspHTyo6eHmMrGx2SynypLpt8w01mPnXUOfHD0NYCNwfyc2Y6gv+yJbeoLm
gvaQzI6Rlft7o3Bml4pNzWB5iizsFuQYiPAWOFV2sZsbguduSCqxJSV+AQdO9ygS
8879jRmALt28E38LOldPVq6o8YazsDcmutjVB180ABa5pZmBHVsk71GQsFRVLEp9
iZX5Ts+7iwR/A8g4l8bpGJSvb4doXkFz5P7/Mx1iIz4XNV64omY1ptV8YRz6zK6f
qJZ/+Cfq/gJRNgH1RE9/AmuV55LgmniU5U+IRyY26cG2GacopcupyJ4/5j/7o4uv
Ja3okug2v/EWnwa0v6+3sW9hGHzJim+AasymCwjAGcec7EKpS2Qo0hKmDn5xQ/nF
9JWoRVtFUHgY6iYHG4MphnLXlEUe+JVfPPutdeW+nwUFHNAlUctXrVJ26B3+z3ba
hSd2TXJqj3oqfMCzUvmnAAMr4ASBxyoOQPu9cWdLbHR9E4CgJVMfJSPwfPVvy1DX
Rrm9atCZR6Jf2xj7djZjwq0mztBsRLLT8VIIsDUqWqdQuXqY8D+Tme7Kyi1x1DR8
QrazdcQJcaST10zHp19eCoOG6qu5C69GsA+obyPvIw0eJ/kgZ8pJqps1mOqI+6fd
Ky2NvV+BT7D3OsIMeFuNsjJST33fDwS5UweHzZkGJk/bAlv6n4wmN3YE+VXWmEMY
ZQX5A3rmKDuy2KlH+LWen656rBeA3q9i72HvfMXHdbUaQ/xyYd7TyrWrjRIVAuUO
C+nUoHf+uTgmkUO35zHpGMadj7kEhkKZkxYYwRRocTkGO/thnT3cGNbIvRC6jXgu
0wyUEzHm4SxbxlwDwXhpPe4i3Ndu6wlkq19ivC6T/FVlKZjcdy8qie3a9FC30YbJ
NFHJ3sN8wueKTpTu+gFtTzlavl6cmFNE+GmBZN9N+hBHJ+luvPwuHAisE3EyOHA0
eLy0dJWhYfXV2fj00DEjjOiL6k1Fi9d09WJznEZDriZLfLd+UZQVIXQ86mVY0f7a
Sg/p9IZSv3UEsHVo7JVeSFIcGVEY90Xl3BMaDp2+dkjAKqhn3i3oDYrCtVITYVdZ
OLjmH267R3PmCn9xQw1dtKbTYtcOQVxRnkuWDFpnbA+4dn6epDuDhsYBt1jZo8yR
16fNV8VQTw6xqWPMFAqf02qBCjhmA3bJgc7bGrOhredu5/hogarlLpNXflA2kb5n
4T9VwsNxqq4ymwoTPHyDulTBIkzknT1fXBBI694D1PJi88JHk6MRyTvtD0r82IFt
wbzDV86ghx1ckBxqlM7Pr8LZci7HdkQ5it01Gq52ppY2Qc22dGEpBL5p3I9qv/au
2RxiAjatD9UOJsmMQe2vRsUgQiBPOoP7eeNJvt6BKyxWtT/Z3OiLCm0uGHxX5bnz
G/28mvcxhsa5xbFWSfuyIdtdvTVrTA0ZSjxj/L2TWvQx3+BVXrA47D9Np03pGH7F
IHv1TEA4SY5hgumjtswMACHLgLUDf4xdOHcjjQoXQrdHaRrB8TYczCSI6RgKIJB2
s03fElv3FHfMocfnJLczM9EkyS84FT8500qs8q9Ples3XZZ+UFrOf06BktyF23gS
uQ0bVAaAjyCnDgVs/sS33+l6HVxZkbZV02douiBsagWVoW+5TN+AZM1ijutiiuKI
gdX9obN49rRua+SLhPgRgepGwLXroPzk0ZTJSKwmxFedzzQnzXdxf/bLvxmiCs42
5rbnlnrVWihCOY0wt0VEhjam7Yu6cLJGFXj3/NeNA3fyZxUwimqmkdAYUNQOxA13
CQOFceUalVPHdL4Dl443BYGnr08Cwyy+l/iEQCwa1SB/9gl1tJb7gpt0nAiFliGS
tNea1y/puUrLk1cIm5NJi4YvfPG34Q67pzHL6y5PHaiMS/nRa11a9ESeRP+YSmEw
M1BhrCsLDEZLPT2dYzNEYhXCPn8u+noopkBQuR83WHdKqOGxom54BdqyMZ8rx7ui
+5yN/9bUxUej0IayvI8PtqcR0HYqdj0fK60X+bkvYg21YcD6pyunqxLK9FMdG9S6
InkmQEbl6ah8LjVwR3RkGIwcGiVsCUTS/bWKzRx+B0xNcZsmkcqVg2In5mGENlPp
VGeledbLMv0k16ueMzLrOYddz/m3u5Y0IstXZjvkUhuXCAXtkhFr6MFHlCtgmDMA
rsSBOcZtZZIyGpSuSNiVAc6NUyyu8HP0t50/8YfPLkllnSaz81Y4MVifpxSd9UnN
kcdp3NL8O314+pi4AMSgQ25JG4eVRD4uQTEw77zi5SaNLTD0n3Dcm0cXHhGL64D/
2J25qPPqe5x3b6hmwdAPGwqWbLVSmy7InXZ5aTFGWhpYaOJ9CuRNFfoUg/GhD86l
IiY4LLiBqmM1uOl/I8KlYnrQsY19fQh9khEkbXGiboV/Q0fAl4qvMNb1MhenMo1z
d/Ub7pqXxvmFob1DkBLaNgC9377kewe1ArY+SAQ7+U3k6fRckjrLT0kbj4BqZ8kb
9pcZ/IHUc+2r7eS0AyxHXHFoE22yJTJ06VcTbt1QF+ASZkKayABMmHzrZ/RK0yGs
xIMF1QnjKtBD8TiqgZ9JoINybpHtMnf054wQL+gf9BIaa/pGVSbsN+p1Q6w9+wKB
O1sIog/vYV9QicKL03msek7KXS7jhmB55uvBy/HlC7ScDe2PtbFxBqNiRCIKy7G6
ZCpwjjGQXw5nm0frpMdCzl8oHFnnwi1OLWHtS9WAbZblN8r6QpD7KFnHuiFxc5mS
yClinxq+t906QFBEjcvmrLXoMuHWE3CrKytU0rD0bAokleoj0SIs5vrrNTZvenCr
6TZUrm1myz3dmUh+/y8kmPgjCliP49TlOActGIpd0tZSSyn99DqdljD0oilII098
PqPqhqwKCHhCBY4Zg2pvngkJTc8HlXYhOVnwT09/0NEI0Oh1gwS7DFUrnYzuoppk
v+KmpJOmj06ZL5jBYBHiyxJ95L0BKH+A0tgLNlejmemLRBMBO8aT9ZCbHeiA12jk
S0apUcBGgb06AJHcB1+DprzCOBdbk7X9+dozfqghj8TAMxiWypUJbeB4Uj+9TEzT
+P3xyQoQjKHMrwPnJsIz6Kra3fiS3XLrxZAt74lPTeC9IP+fvhaCWqDLWibmKuUp
V32aAtDOPZrhXyG052MuftwUu7RGm/ddMwJC9zATjZ08ogCtaSVgyEG52sTjUBpT
TIkXLSr8EpkMg0B275z+EYvk6Mf2zKauVz+t1A4cCBiyqZ9yWT/WIUYjxIql8ruN
ooQCnR7iiMsSg8yvKJvF4KMcZVlW3yTpCx61aXg/EJyJspygA96rOd0kMfio4pKX
OZCD41n5YfKIhCju06IDmyzt4YbcctCeKNzjO9KPT4RLakNyk81Im62HOQVmdimT
LRLsv+GHiR6bSQXMK5rVyrIJQkpv5BAmfZapyQ6PGMBZIMEQ8O9Rf8fddCYP0X4s
X5motlq2/GWnC0XbbsCrxO1+YCEIwjjxsmdYoGmgXvBdf8l1WYmNFokg0uofL2dz
5WEqXB4qUPMnOVrRNUA4ZX8l5vWeS+2aLHD1qVdcKgmcSJTYS1ernDjnanqWDGmD
vC/xulKDKz9b2889eEfJL+Ijm09QK9ylg4MZAMfb7VRHGPYy/0GoH1xXapeSO25y
2ONhGpwGYeTFMZtkvWfeBZ3IwiTc8POr7ET1xoN3LPOKhLe1ST5rkVoD77eEQ2nz
yk8aTW6wNqGny7LHoiYj5hklebgsFSPo/R786O2E2S8kbnx3/ZMNcVEZVmBm2pJf
ih3zgARXyzFwDyWfLeg17kRt55VMOBQVEe6XIy3j4L+9fMtH+PLgDMa5vEuv3MQr
oPVt+PXgRoL4XYc1CIMQbGQQGI1QrXCSjUic/Jjv3W9GAlYTxYIl8AmT/MqboSgo
nGa4vJPTXWI91Jg3RBOJdOF2/52YhuSPXtCE7HjLH/m6T0VxLBi3V0xBiUWED1AN
z8lLAMS4Wo2mVzt5rGnigYuNyz/58Nm0cECuyNP6nNNbgBVFlZ/DhFVvIjO4R2Nm
i9eq4KbkfoxFFmot3cMqq8yWljKdksFFkkF8BiQGca8q3s8ateHSaWl3fry3Chzu
EFIpoZfZNh0CUEglk989KQYNGNz798u6ONRf/NkC94fA10a5jPvFe+MJtYBwjXgJ
6Xnux1UBbJi+QdUNq4GRddQlzF+8pywbavRpAQ41IhIRJz4Bum6+FytnjZOt/4i9
QvRoICMSZ9K9JsGF5XNjdaXNMLvfEL36KN9ZwpM2cWHtKo3coNP3m/tlVQ/2a1Pb
50H0QTsQ9msihUatExMXvlaHpIoECUn2/Kw67HtwjulCuXQEO7jEubT4lvpT8m2C
7vAaMWKQlZCtzB3wiX8CWc5AWPHCenoBg+ppW7xrnUUByF3jWGLSkbWgZtKI+riw
c00onRClUooTVlqbEi1NXsjD4P4pyKx3m4hXJPwXvhMzh+2T+iQ3noygjxwIKEc6
SlgX5Rv+iDYeQ9l7YJZSfFbejmTu9BXkqBeqKCjmdzOrieVwM/H4HTCYERNeaQEB
2Ev47B9fLFEfvjewxUyKngmPdSrftK8mhymgVyqCcLbKkCTgW9C6QNau2Ps9uPXx
VjKzbHUbvkLYuLpkH4TvkV/n14jfXgk5Czz5ezM5l43GM8zdg7k/2vj4mM6BXw7p
3yyDcoakaGfCTkKv24c2syLCgcv0K0sz5myb/pkK0r2xG7r6vLE8DfE2f2mG0Uco
4Hq40gc1LcX7zkEUHUAGu0KWwl34X2L+4RHOYm0dbxgAubaLP9D+u2DCEqlwiXja
m75F8yPgcZq2uVUwmNSoYXTTJVjuSpEn0V/rQwJXJLKZ5GSQjowe3xmB8WhQmgXi
Rq6Xl5N/ZHxOsNNOCoQoVWtEfeNVL7BlnT17bFYOQKcfwN9bHslTbqMJ78Ej50ep
xiM97lP/MBOvFVhj9frBvEiPYHDFjm/EOMJ79SnwZucOHugFBM+w9IE52XXMQhvx
22p9kCUIdK5nLrh1V+zcpPthJochHu1VzNKZlO2NEyv7R9HcrkXyZVozNrxArmWi
vylwXWN3Z5K6NRJPjiXWyRvAiKq9ejN+TsUen2O8mQoVP6biM9uyWGfKOsJUBgDO
f2fqmzhaolYiNlMMvZp7aHDdVr20eY59ddQR/uGCRuVGVGKOaT71AL4vT2BVJlbD
GDGNRejiVSupn/2b0KIQD2wLLVh3Ur6ReHM0jecINJzgZ6amc+p8+D4CZnQzA/rw
PRdO++H96PzoHRbqffN7qfeQx+PARzu5xXKztkrn0l7aTJIHGaujCdNS9lBZz75L
RAstDBUsCTgPVnnvYzh9FF7rfIf0K8w/bQqui8SjF/+FBSqi4w5SZPSyw5+fl+0o
m9sU257U7uxhNdZEVMDh/oHpU1cl8bnmOUEGDSq+UbJBx85Lk8yqt63QgAK1ZgEl
NyCE2IzLaV1McXdBS3EjUWdE5fwyerlFs5PcCmK/GBvhp4niKTZ7YVgoHREhDikh
wIKltMF2z3b6XNDNhqtI7GfxZBDb0B9j38OeH+sDFcep+juwILn1xct17hKD+iAj
Ore+1kElfa3Oizthn3IvnZqrNqLEYoDCzYobVmk0NMWaMtMoBda4YNgl+ROHbqBd
GYNZdIBoYMpA8P2Dk+APejtNF/RkOfCq0dZvc6KeRuOvUYgM+3p/7Iu2n/ni87Bi
UbQTK3/KqcbD1K2pKNoPkBR0Lfigcu4Ah40fiGcyJprLXKM6Ez7BlMt5pdjleRhG
FroGTF8Z1oDI1sGtSBY9E7K91EMeXpbS0X3pP/QrVdhQr5FiSOKVEKIfDEB3CwC0
VBgv7WgDApj4bRD0qJ7865zqxyZnvaj3wuY76dAUACRZI08wNIzWrAestRUhUthj
TJyjBaFVvE2IeWKwzXfkFz1Aqgjx/HSgAOlDjjoFbRJk7h/E3379Hqh+R4JlOJie
Vp2CUmbzoNhf5G/puPUrt7d7YprclOV9qljPVqpAx3MXzgK9J4WlA6chjnAy7ZvH
RXzrBAo4fVpCIG1rGoAbcx0sg/sFIonP94CE7LulP1v2Q59gAnEhQ4Jznsin7itY
aaqPHzNVZWa5AyHA84V9BSk0jOyNT/lRWux94NJtjwRHzFUoEcl0YmrfNzifkVdB
Ku5udRiMqbARp9h9fHkORrE0tEM3+zs4KHwUdZoKDlYhpSE6wH3Ds6IzhzuT12Uq
vcBh4v5FW/raIhG4hXYXSLpOEPZMpBPKuUNBwXiAxb2yKh2Qrs3QFvJa8ka1mplT
s1zpFNRdaf8NwyHcCWAYMay2c19F7/8RVaafPlJndiyR12G155cN5TKk3tWbUa0K
o3lRDrBAcAxZ4pkG+LGUJndrOspJONEXLrLkMg1wbnpsdkf1lNSMeR/uA9nXNxzO
mDliZBSVD93rn1d0XMNGa9X6G/mJ+t5jP5S708PSa8n4UlhRwTGM08/8OEk87njC
17e/rVsHRRP1hekX7LG6/A4jwwPlUGC5QcnjKv4swArMLmFp3850uDriBPzOsYha
bZWAWGHlIvqq/gSOnemgQpzKVFVIAbmTgUqII6DbcSwUOZGERdXGBL+uJbM7RzgP
Q9AQ5FNn51zmekgL3+rD5dpfz3ddI5agCoXRXaF313CdF5SiDKQiVcqJp6WQLpHL
U1ciDc44NfFjZ4RM2kUGxCFj2EU5X/I0LotnBgfV/ET7Y6XI8mpouN28QPhuzX/D
1SSlza3KNvPYHHjv9gB5aYP0BhM1vQORYkfzQdWui1rrEvoq2IqMzf7dYxb150AV
Ns57/8CK5xO65bQQRBUKdW/uKugHDDWNlAVa2XCb3vQljtLxwZXq5BY8c5HaUiXV
dJ3LNfETZoHPypZiLYkYWSsYYTRYmRXrwqFhxDX193medOxEGbC8SnqiVD5eR6yB
f4gqQB2meKk0UNVQ3zE1bm5tn44hXPSmNnUrv7bDJ2rNQObUfcJoIrs8CYtan1WA
vQkL6CvWWfcJeLL0YdnAIFfVNz8+rTlq6IR5g1Q+kjIJKDs6d8L9Ai5Np0Fszsyo
0XR/IB5pnvenF16IeUCR0VcCNpvS6pmKU6UhOf64jVVuO7qeBULBwIy96rDPsusG
tc7ZanI7vbEmzsFs0lppnLqDlrh2VAea9mqwimO6EOypkS2dB75avAfHTO3aVeqH
M2tlgZoW1DMMpacJC6YH37OLNW8HAa3Vj2YGiSLxdV/5grn5F6bT74frEr3h9lY3
rFH5tQTzDO6y5GCKAnYnUsT2xRAfUqxORO4ByJzl0GwrgacuoxHrzI5H48rFuFvz
i6ZVxDTzQp0bUx9ZIhq/lFlv2M0SVhC8rquPMZvD9/A81y3jcC2wapL2mSWvcgZi
NiE75Kf0SSDqWsioeEEICM4u94cNhmix1JPo2D6D77utlz0y8HCMYeP4AWiASW/8
28jk+HNkyiE5rhH47bysDv8Vvp1t+wwGgxwU8eNRVA1kx3B5JRFf08nliHsCd8uw
1AYPKszMAsgOM43fbyg/PiKYmvB94X2T5Z61T/NHCEHndOIaijo56ACo8DfbgjKo
Qpr6WgA1y3gLuS67H3jkAMaVKObdtCEY7W5l/5Y3AmVU0WVbrnMMh84DdphujFqC
VRq/GdXDSL9l2ozGwlXgT+rAVlS1BqQQxFG/ywD0hKdkPL7vEjhPAUiyoEhK68DQ
Qdsg7YcLBwiXkSHB1AsIEwpxYU8A/jGV56unZ/yTjH+KKIlla/MS1go1zFjB3A4i
EXEitJS41k3GJuvEqHRFfePRthakJs1gLjGfEXU9DFFayy+7WptHkm3jWMTAZPtn
qkuwsLuQdA2bbVXlvsRZ5XqT5x5/LEbd4+hqkaNSkVF4cL9jTvxdYaKbpFzfuEGo
S39j8DT4xnFhvc6wGj7nDlmglPZGux4/0L8bFbDQyweJPzuJRlY65fXfleXGy27M
YwOlZeLBSOI6AY5WeTTfjsXk2IteOBDLXv14Nc6HPai7qaGeXzSOPQaqe7aARloq
oIJhkb5EhgjU2f72e3vtRvm5vHX+qqXqVTz1oE67lerEw6w2JNRna0X2/06m43Bo
l3KtnNX73O2QXfSYRZ7bsXhHYSfUOwdF49m5Hob/ZpV4S4BelsdXCn9RW/L9RP1h
/BRPrMdUiv1qi2ezz/uW4KQweFuPKo45N/Mqhr2jxQMiNzIrTY+ddZKVrGYlc5My
hGa+M0Nl/wlTLV1Cs4IFLDgXUi5yczHjL7Kl0OyktF4TDqhWXJ/N/cZ0dhPnKjie
aIMecQjguNWdpGZs8CFP6CkNHK6FnAP2KxRgk2TvD+rgsdnJVWXoWy0uGYl/jCN9
ctgTVn/OwczTDTd8H9Y7l2VAWabIIxckPjOG4iKNemf6hgWBgjPrRgxL2wlINkvL
olz2GjBPtXk0caxvT2G4xgVs9eViea6C5v0g8k1C00weHSqdUfhe9sveiH966g/x
n8AnKOeMS7DzYJye/ERul3QCSvhkhGY557LEb1HNaGyngFbeHD3lJu8kd4atnota
4OVpugZR6l+ak6PPbUZUCX4vkpudmLA7YBuIT9SRJef7CFm8kfjvSI7FpmuDW0ad
tIZHb9qIp1DPUgqta28WDcsc8W1sz6E8+YgFm8vCJOqS3ueero2UQ1Qb3+fn1DdM
/P2fprkAZRYKX5pjO2c7hmDpl2xPbKsg5XU3faer331SgZ1XxSUYvv3t9jOqVuUF
0EMhi+yKceCQRtgdVbZzNxlsX8nmiUeNiFouvQ8KHIrIvR/U+c6aH8qTp3unk03X
aItAFqIhwarFrpL38gj/Faev3V4LNDrsFT4xAxsBrb10NXT6W11cMf5GON7n9TTE
1OHg9WRny7XaoVL7dj71IDNJUGiDTg7bBrEavTlZeHCNRxrv1o1cJPpbikQPWyDY
QM/6JgfIoK4mvAGynZu3GDMlZheErsVu8wHiA4eAERuV2aw7OFKGGK+yT35VpF7J
ql1A7jeal983n8gpheNpdALG9lNZcWZ8WRToTI3PTxq5bRprILmAyc6iuvW7hs62
UCz5m2+cf3DMqw6rMziEq6VsfvGjLe8DbBoWx9oLWaQ34VsWVsndtPVTMFS4ewwG
wrR4wEnFrp2rKygAFoNAGSdQ7rkYTIGzEjZq9crupG9ji5mZd+/LLwnTvdmYRLoS
A+oXuXfRk6yOIU3ls5fm78Oip3xjxV2ZGpGPHWbo15tjqLJ9Kd7bQZaPQXA4OjMR
v/fA4D2LDyZKRL7WDcSeoevXsjdw1Hc7eRUmSU3jnYlAN9KG++KgXWiGsnMmSbcR
ZQFJLaFzGV4du2eltaJrxKnm0HUeoWJRhpMYC8pwcVyRr5Wr07hhhxxaIKlIDTo0
wFzlGomUbm+L7Y14wOdeLaziezuzojXS0bkZRqyNrggE+kX03kMhpr/iSWODUyt5
w9eGdAG70bX/37bjgGeqlGR/DqJQtI1VonX8vnBoHcKhfzpOapcjpmqS5f5kQigk
wRfI2wAIkEtAVutF4UgOtgS4LsfrSOak9zGw1aZGZokq1PcrHveayJE5FQH2wUpM
X+0bItgLffPyUXh6YjrFFNcZb3R6pWRJYK96g0QowIFP+1Kx0F8AwnylqZZ7vd3W
BioFXLIifVLiKyf9IGiUtEhG1rvymvFfb9gmwsDo2aBAt1l4fKBQfceWwoMtakrq
QSLCt6vowIUOyAqJXcRMo1bmWjlAl06lxM11CO4Ur9Y57FKltnhl1PD5uAvLpwIb
ZBW/i5dfkeoNNtJdlhuO5xJ4RObzqpBZehhbGlRrACVl8wcjAw3Ugt1jrj8rJQ3G
uOceeYSOVifC95d6O6qYtqzHJs7qhp0jnHO8LLFFNXqN9pfwraCksX+1fjlh/N/B
pE7BP6T6HROKVbJp1groEQ2BssnhuUMxMcHrld7bUigmGARtCk8sjFYzFiejSLRq
K6XlmyaNHXIE1UEjICdm+71IvxsjGg+AZTwwSp+XT3P8IlWiwDYW+UxKGGIv80JC
VABStXrM/dsn8Oxo3K6mSMjmQZyeGDHV1W418YtEOX72PWh7Bvg1g9dZ+2Lh1sG9
d57XDPJnjaVV1EW8pBetLcx9hDQ1PJwT0rsNSbs7f3yg+wHwoSMdPEH3p3+0BLku
2fEkKH9kV8jC64EW3J/En/Q3YLP4pn7/i02L+rTwWnHQE+0CE2+RXnJRHycZR3qW
ZP1DZXumhNpwTCoXcVUA1Xf5hiKGj2Gb7r0fTtwwk3dCAevu5Q7Eu4+O2CHCltqI
F6/6NT/kjCxgQol20heAsOMAhhv96VHAYX058O71anP/JX9L/xE3OuqkWExIg8mV
YRGZ8Ea4tAvhPJccVg7JH2JG3qgysidpS5ccRv29yPZf211SqOg4IzTqY5hujlDI
7Xs4U/hIj4bXyFxPhsXMPJOTo2G8mr1dKAOHbzn6WXMD53nDk2ANBV3h2b3rjtIz
PmGiNbxxbKfZsGPgcPJWPAM0cDv4xTRDYIE6Rw3TBQo1tE90p5xOZozJ9vu7IbYg
/wL0fSo6ACgNvmvs1sx7tmj6lT1nYWGL2PN1KZvJNe6I70Dhko4jZz69aK2HcgI3
wCs4Ue5GFTx+Wvma3k0hFwyl7kAZvt/5riR1/VLp1jFFdc9ADq1oBl94Gw/86ARP
5Q38/Np/J5xurLWfwzdO2uIwhJGClRoot9I2SYbphPeHS6wmFkF6rBzMhoUxaAqd
WTzVSpqSwm4PHkUEODRPTwvGoSR/UIt4LfLfx2EWdHoCUERBdPChAALJEXBas+/o
/7hE+Nrjn9q9RCui8kHKBy6aI49b6TgZjEeXgDU4Hte8mWeF/fK/JcPizqt9BOJ1
H0Qiv6G8OWAKBHX/aydSwB6AZCYxdaECtyxEvJpYma7UkL+lf0iQLc2ZcCYS20em
3Vnyi2N1A8JVE+WlwddfSFrZ2kJ0+MVf08OO6N9XpF+nrLLB5jcoKkBvcA+Lyu1u
TIsZz0Nq9Tst0UwYG6C0V+R+twUCZk0XmItORbP8e23q36LqQf4uK+rgmUdQI5Vw
SMfny3ZeO6S6egjc6kFSb2rrpi6sgKxRXZJcGry+p+h4nYbeDlThh/aBTTksqnnq
QozCyjbiOzVZrZbrXGoO3EChBMdVUptI0P9MAEa2Gk71ZXSNm31wFREiN6ksXmKy
S0rbwul5V3p98TCPt8Jft8vtQwqOH6nNSCHPoAOh56lL6KQqyJXSurN6WefZxHXz
88pp2jARxA2QF8jvWEST1sqs1HEDDC4nrRsMHM5lFCaK2i8AUkUcDlqoRX326EiT
Ha5FZfhuOHfUQKpCRxv/mPJ67bqoH0+T6HWULmwb28/rpV4OzOgsWwVRa23faM1T
zyo0MEHWHUGmS8Sib4mQBxkty4NfMDnoOnV46IbsUFX0eVCAUuPfjPMuzgyd4LrJ
lJ70ti9ANeortS/Iqp68gShkXFHCTsRTFyJ4yUJQSjWG9frLMyWapVmJXBYLr/7N
55Pa0mGOcvlRV/0GHu4viIrv2OyRlkcIY+fCOYm8lYHrvPKyeRqrpDc23l6yrQSk
nTZ/bmDJxMsK9kyXBP4aRh52oKfOtrhbcwg51XlsyRW9t1CXq89BHIwdbK4Vm6+S
tvVDA+yVDZJ6kVTPF9YGNS8m7/LO3owwABR2VirMPEl+WP2YAMy/PaqEvVxx7fdb
O+2vphGZiYvohkKjliQiL86kO/3OucfKff3qRLf1SFr0xfFVyDqMYfyJVcmodBu2
poLyTa3HnbCdVM77/cZ02aWEz/GaRxbAj019/LWFEsvMowOLetL+Jn7O7Hhm5tyJ
38f94anA+80RduEW9GT4/QgKdktsmszOiYkc31A9mxDicq8nnJ5UFXhyv8blqUbf
f29tVT3i7qjsrTDtpEa7E9yuDGlFYSNfFYm1VZMhsJX6eoaBlDJM+yi3J10Xx9b+
dVTUqsUjjU8vlNK2HQCMENQMnntiUVU3gJIcp8v94Wh6gwnvqCOQDmcLmJY1npaI
2IxVUTQsXImM4WoeIMRswQZwQWgj/ZRcCvp9iHsf5fdUoH66XAfmm59aY6ZoRm3Y
vw4MsHT1ZhW7hVymGdRLwByz+a53vY76qf4d3crX+3W0nwKCs+h+5Id/HKpzA36h
aqcpBHY8r9IqOmeASiuKw/StyHp8tYLAfTUcdC7AGPIGC/foWh3EdRRQA4wMO2VY
2HHc7lz2moFlxsE1AyXshpRaulkfyvb+fZNw1QFExRB8nJJORnRh/Vy9Mve7VdM9
D8AliIUgJ5ALGoq1pEi0kML6afEamBUJO9tUJLXp6M8xYII9XtFEOiiJo8i/lo+V
U0rJBqly7ih8RRJ1C7zTLRJDAAOAXhT1YrvDfjkeE2p6IG+0kNA/rJpNRiTstn+5
+sWgIS49h1oenCYFM4uylOTuBXaUlPa++LSM9QWVuiWoacCgraYbpHc/LHwuGE50
B1OnK7ufPenHhW9FBMdyz+V6JWqNs+HOQ5Q/AnnNjVEpjZzQc89RXOCJLs4OY9gY
S0Hg3ll4a5oiK9oKTrjgIWo8brdD52QU5w0XFytqoW+Y7r/j6Caixsa2KGjhz0Od
XJ6zSVsyf6gbqpuGrEIfvPZgUB09i5LQNq12++xij7zvwXdgimMuzweLLEzgPlRn
+fcBpfKAkQ8FU05flOJ1uqtPNh4bG9Bo12jYfNkJheKx1unnh1l8Y+9J0ELyHBEL
aEb3rWayppGTCkNr4YLC3refgg99lSuZNZ5nCry3MZzlz4kYhTPLu1t2kij54C+u
dhBKxtxDQ1Zr0H49wPEvTuRijYgj0giDcLgK2sROD1StdlG/x+KJIR+w2UWcaFFC
tb6OiEfIdKHEPxF4yae0iFl5gmPhJ1UB6ZCQ48rw5nJrWGAp48Fkxobp38DbG3Ph
RY63woa+m8TUdm+dTH7dHdAsLFVHLnp8ElSp2ZJcqtj3Cv4JEyqvxn3ubomh2iV/
EdON2GxubjRdKVGr5O53KbRHR/w20b0T8BS4joxmmfVlKxvv9wKTJkD2jJPwNumR
RQj2htJVuYdqNyNenvwx9RWiF4PBURduQQHFhh7cJrgtidMiAAAgqXRJX/nOakde
VEsJFatn0e4rj41WqrNuyxgfSSnOFWo6Ogqz3W10k5flvOzNTtIHfVn0g+IZoqnq
TA9TsVgzF997Su7oUkmmJo70akL9DE7n1+3SEx0pYjoZzcfOeMafrPbPMz8hos7g
GLWQPjXCcr7KQGNsQfJPY07/W4cJ0sk9bQk/4VjPK3l1IgTCWMzMDYdt9RbUtTFp
W9oJMIvTn9/SzQ0FHYcvBaUHAG6ASJrueXthbHoAcsKRByLn6vct5vjZ+Z1juTXb
7D4/1J+mCeKXVTSfkRzU+mbFZc1sSFWgGylQHjteVfte1Kmc9TfYzp+bVrOFQwpA
yMcSOllXNXTCoozomFKaHtqsyFcku0oi5vGiGoaqNCvt1MVpaAZonFsKPZNsmaid
/MqciC/ce/2jtVTqehK8TOpLN3FvXVD/T1R8DuOG7pRUtBudaWPgLuZpGit8V/u8
j8u5N3hRMB0Y7ovXN8NxUwMBK/MLwAai7o5xCIyzP1kT+LiXbDQWeR/FH7cKTa32
Ygo/CS3Lxi9t3Ec30HM8uyfXFHJynkzdSfEFqGXomkqTzXpXgJVd+mkTVlczsqP4
0EFvmEGDw1ejmtQ6BE4Amf59HCDRxS3BBNybEkE1gO7XWkQBT+HA1QTBVgK/sajB
nOoUQXFgAuONFbe3DV3eJkjX71nuodmBCtoMVk4hGRK/JN4Boy/ewuN/+PxGySVW
xTEyvpyEXfgIsVvsk/gzZex8untkUHOzZRNZ3pg70nrkupAScH7dbiUJr/HeV7x6
zQuxRmw6+jjODDEsTqchHMCfVwTWcM38NewJEW7L6idVVpPqqkO8T1RPdoWNotxu
SmMf2MvrRid7lPuqgoPa4m9345luf6JYF5OyZa362utFM2T0MBUlQ0yvawVgeDjV
pITKHajYyi7ZpGpqmsFrNSlktu6r5nQQZVDXKL0EsH5DXkMz4Zw/t5cZwUQxrhO1
Z7kNJSxIH59WTdaagzKCM4ztAcODCfUJkMJmW4XfahYnLVof3F6t6pvZo6HwI448
FVD4y6ssSEdJb5Q7/BTueRwa00h/dDlN8+r/zwn0AkLISu9OPlBJ1BbEZZUjlVxO
MFWH++4kKMkiX3Bqsr+HkTbKOGt+Zu6TRN5v8pEatl2+cHMWhvDX9KaBd/my+9f5
D+uKtfujNl33pwAcja9FFku0bUlIuNBDscfMuH1DjHsBP4EeAob8YQQIXRnAVxwt
Xdsrp0EsVXSWYICVDzzwsOiHkB25jbkLRL4ISKSestM0P3TC1D89r8W2dxrawsVc
ex5xSDEWQoeq90fRhPeU6P6CxgPzzJfolw1eQy/p55eIPJjyKpPUimFUPSrZB8VF
/1JDNjXTn/ZkRFL35MFoTjiM+d9StUtTIDzMy4c5xuKyzDBT/PStmQXvFMfiGyH5
D7pbWwqr1Q3IrzAk+jeoW87lp57ooImFzsfhqDL3Izs4F6Q00Rt1YUbYd15IodO0
RScCen0lwXfyJKkgW+i4uVl3uaenHaj0kkhsl+t/XedEX7bcir9ajbFmFBdPXCUA
lTowV29+6tTKQhgylBwRNvuB7eIrBULTPSAPKn79m5hiIuUydM9jzCBeoPot0rV1
utkSI5q4aTFfKKCFVd67ZW050yCk4EXwu5ZgnsnU1QJM5/QxmircQsB/Edbe0BST
a1xFMu0Ga3cBM2z9IWr5taEa/FaaRIIQBvGXa1WEYoRlMFZb42hw/rlQQZzO3t2k
glI3giSIM4tkfEGJhANAwXzxozCvXoTELHx2RxU3Trywa1c8JWhCssL0Dc4cZCJP
ub38irOzy7fOLXS7GPBkIS3jjQnRzsVWZMqq2WmgRL9q7WmcuHEhc6QbrsiSUZfJ
bENKyl9OzouksS+Su6ktYICr5xQij92Sn0HuHI6QboMU3zmI16X6Q8TVGPeuxajl
8gp1CkQhT1yalwDOXAVT6ULNVmPFyGR2aezvK4idotBQeRe63GPnJ42Rh35o57ki
F+wUg2jqb2Jq8HU5+OMWdMgCuk9T52bmOoCdyFMGuSzX5GPqwduac6kGYB0fFJ4+
UsOsVJsfGBELH3Opmy2YkSE9aHAu2+lGa1cjU0fEyP/ZiRNuLVQfy2UEWTaigRvn
xeQlBgvIzXRdXRqrB3N+R+z6fECZBOB21UW/zVbVBxb+R9AsAVOqWo4VmxxWx5F/
CEb++g6r3gEqDlu0izQ3aX5I2klGgReDqJL3nTMZawuPIP2Y7gPOL+Q5vz/H5aYg
wfBDGS1E7zXVr7KycTkXV9iXcL2sIXQ4NAjRo6ZuqIAwpEp304yv/xQVWNTkATNf
+PzMUOzm/396PuvEgdesoML5d3/j6u6Syf+Pa9GZEoohqlwFG632kf3jKZ2nqFcx
aO9l7BxAJ7Rmz1Rd1rbeCed8Hrc1JiyUkJdItK14eKlL7w+g3cXMKVBPx1ehmKSn
VV1mjoP/j0XyP7diYNTdrkATm9e0xYS8qV4LBxinWcSmnjLRvSwWxZM9VN+Mw9FT
iurE9HudXHvKTdNqgvnlvHfl/qGSHZ8QWJ9kMx9Pd/I1qWWMDaLBVphrFRQBljiG
OtdtM+fRrhEcbCDlrpDFj/z6XdiQQ21Ewd9t28E8RyCmjg2xLR147iLNDB0ADuJ3
Enu0WrcZkeY8NypH65SkaRLHtLidnbQrd73XFD86xmdbY9D9KMhEE5Z/hATAkCiR
poAGMT9nJhKtOPAFJoc2AE7ckUqQpYahIGEA+zyqI9olo2+pbozS/4eZPEi/wRd2
FQ5/1zGkojsgmLnfpJisgtNhwHngtDIFxjw4GnqQJut6z8akXZrZtfSzOGzhxEFA
pQxKCITvo3fmRhxqceC4RYZEeTIw43cOflKSe9GF1SzshpR+MS1hS/kZqDVS4WGA
QcBzMj+RlG4hOxHfcYnWC/NaXZIeXS44QVqbz8ZR7+WOD1LT8PaP1UPxe3rqKXZt
dT2cEfrvWAz9krEtK429KkW5hizci9QlYAejatuCN6BzSUXKes+Tocj7AQ8Mhyhv
B1sg0eXyIXn3vXQ7KMcHCeKd6GEE77W3NkoHfYAtKjZ2sTfl3ZEqJB1d0ufLiZ+Y
SO8bzkQDLdaGlBxIswXDPkrmLYcarLPR10Yf9JReBq1+TUnvsQVEPZgbUfFOkDdA
olo5Kpqqjh6EK6pI2KMfFeIFUMSguQNTq56/WAbhENgYy77CsqEyAOSsgw+Ts6NX
Xj5Y24BWhalDzURwYexYn5m/LXtDykPK/nXGzTVXPHP+9GDcOtToKURXfhoL1fan
hCondYzR4qxWuuQvbyM1OUe0OBq9Ey9vRwcT0yK+0BNjw7d2WBS8K0yQKoQc5KHJ
1+/96DufJOe0E6lkvOZTIskGcu4yIe+P20XgJopj3qZCJ6QY4dv/lDszzGd2OfO6
8AE1c5VdYHfJducC7PLquUnqle8TgjHLyhktOT7N4iPJYBzaYURNiRR0fj+V2qg/
RUew/Z74c31OYbHAOaPNIGPV3zLvcrr0hn8by6k9bklk/CaRHy6PvCpnih7EszhJ
ftSC6kGiZJomQapxRy7K/bRwH/5/1O2kFsst0WLAxMOIkLh3KlmFw0FyU/TbW+qx
LKfkafeKfuj6A+4obKW7tLpaoU7yfIxMCuynOG14hDOXQog8p6x5ysMG1E5ty5tS
fhUQSFSFft+CzOhl9Uu3FChItAeyRkYNc4arjP/sTTk5Cr3MXGU7H4mOsEdZ8LWJ
PPGTl7RAljEM2wx+MBbV8xHPIlevRTVMhVOClFoOhdYjqDA4q982KU6THb/2vCVn
SyrOugC4xAsZONarHLS85mZvFK+rBjOYwFy3FlSWLniAIX+3un09+/N9IFs8Kkv7
N5QbsnkiflngGHekh0809WMTtliCssjeGqWKa0QUO2iutOlgCgycoMevRiM1HMgF
LnLPDUdO9YGITfWg6yOJwpkAisgbd0PeD49657j5IUL8O83PZgrpwqY7H4QjULfZ
usEGfrKiaZWlpqGGG2rs2XT83jf2ct4fD7Kl0x4SWoFu/itx02y0PYHwpc0jVOPL
5QmrR7TqT8ruw9D2X8MtAVQsf/rm79IBv+wgugLRc/BQqDsvkLe/zCPiH0yLH7rL
CJPq0eV+Ft/ivYkM0M+s7/yY0C+4eokJtBqWY71manqihSlqOtdO4KGw530GTYXy
nCWigb19E9yJCTTeL82csveYGa6RN65JVp/2zOOkN8whE4KpBi0/+ypbbq2az5O7
gWI7NAX4dsINesO7ejy1iNK1k2f5B64mU6O0UDoigQAMIobDhl15JAUFJ6NVRSqz
sYg98NxLuTL0kVl2l4MBwZxEgXWA8UINO5bOvb6UCx2mKcflnyfOaZXDlsAOWbP8
g3MrslaExsKd4R47f2UuBW4YXd55kOjQcf3dvrhEV5N+GsVTuXS+Llyhh7JUz5z5
GkvVlbpE0l6LJdtCR+N7a9WnM2lsOxSBNL8jxCVpfX59UpPmvwk4q4muBAev1mj6
titMWtjLP+yizOkoNGGxd9CzYvW0inVgA+/61ZImgUxsQ8pdhCypArP7y1iCf1vn
Vq5ofs/pIGmpO7oqXl2hb2+TvoiC/UCuM11u20JZ/uOqBG9tlybTW7E7Ho+55l27
8TvtKM68R1FajILRHSPKkd5sQdvfi4yxOCQJICCdGqmKBbJMNOSxCZ2m1iDIinYm
QvaPpQ4zpL5higG2s/GIuDZqzzWiGYU2qG4/QrIZ6++TmyZCtFi5Udlu4aOmTS2v
8UQb+c5vNLSIka8mN8oBG7E8mxIAZOUd1RehsvDcajiNQYhdcywIZCXLZDlqRiCL
G92kPFtsrFBQtgavo1d+082a0qPuaYwjYzxxK+/qaIHWMt+G6R3LfjXmbFo6kQO1
111tG0sY+0cvMLkVrWdkVsaG55RRxFGJ57259Oa16rFV6bR3GTXlLQT7Lm/QXtoM
n1sXTKJw8XptQItIov9bGYDk8maMzr6B4CCjCwMA2L6hdLHa+5gMKHolsRlMa1Is
AKGdUNF+tYvZ2sLY9rQmavrg+LqOlB0lmKgerY4lHqfZY2G/i600bfLk3UP8J5We
lj3ZD75hFztTv/XUGjiW5OXWvt1Q03Y6zMKUHqLByGgkRttZ/RFKDkT3uCgk0rWU
WjP9tBYEVhD8jSJ+8MPHOHFcsqZKtC7vzz980hquzkA1CEdm0cqgIWjn/1BI4pf2
1+VhPWbxlv0m3ZM51ffkZGihjUaD4trZHEqYiPy3vdLWPisbhVMRuxJer2TCKGcb
1vQCcRDNGrUdvK8EVunJdmL0F8sjJ1b8Sfwo9GKmluww9jFJqN+cN0nX85x2Gw16
ffKzy3NPftkvn9OqcyKZ4IpcqiMr6uFKy5h1qiaVsa6CgJQ7fjYKoGewoACg+IGC
iYoqvhyS8/tIi+VxLHRTnxoPd4yTRDcweYduIuDgT9dzGGaFbhRIYE8T7kvvnW74
ECdOUwbaNXmXbtWW2t5Tnn7sg25uKOFYoT9JkcIXlp4lBlOvqispqwT+zrYstla4
PM35bYWvDeRLw7XqmnqFPSMkRcPzV4o7Yky9j6zGQ65itlTejHPWNTrPPCvHPHLS
hQkrD0RmPfqxW0T/zxEkpNRspyrKangbi0g2NSE5q8YC8mSEur3Ojqzl1RKXBsR8
VNsTl3S5IA8kJp2Wx7jj/k0OQ89WtPCch01u+NltRXeOsua0qMyWrUyQ6Lxf/80Q
YALN8cMQV6pVUpdMqzJc8aAk+/yh+3wkgEwStlmzuhJA0bnDgIgE+fP6x+SL/OJf
yezq+mYaTEzGWK+8EqN//NLCOHgn42EVADHfNcIXxstFclGxnj2fu3R99osuOYkd
V5lgnTynUwT6U7l9Pqipqic4/5cNpG2s44woUg2j+OZ0/vfHh6WUdJipm8Q+t/2c
ymqHxFsaRxcWQ4bMblaRo+WdVYABMPoR+93930hPOeolT9NNRJQJN+spwmr43NeY
SdKMYIAh9May8mlVcnxEqw9fedbCds7rCJ1ReNVN4m5zGrEcDhgKQhhMbEgS6GyG
RctYAkKpEg3tX1tTE1jxT/txYIvwM+5LisT6eAospQQ2VPUct/hzKRJtSL4QnhHW
O4eh2XVm67YDIJkqM43WOqoBjdBPrMbDlkZfcG8770AEPprGBraMO5XQhHC4BGL/
tRVOJicVEIihJnwFoiMoIuWka+RUNJR8F1XMvIX/1YEOoPcjGfRc5pLHMvZsCV2g
9O/9qil/Gk43GUdIwj1j6HZ/rWpf3dhZzvO1WoR4UelgQLI28BR1a4LctpYPDwAK
JbxktnjH9oqdD3aCgLp+ObUVokXTC443CKZ1+3CQJ1xwWoPW1aHonG5xiDQyZAUO
VAifrmfzT6zrAJeRMnZelatfzhm7aiIGtbVTIcPciakpP1w3BGjiuLaOkCnX8Ltp
Wxqf6iwvQC91KzdbjWaAa3qSRV+QBB6V4Vj5r6W0Hwby5hz6fk4uIzsy5Pf6LL+s
thFpWtooggiTpMDRsE7K5A/51iZMtsD/clUvstTUsGoQ2HryhZRSvTKUO4rQ8dVK
CfPQW4PaX6GqpM/ET4L8gkDKxdkRzbGKNiBWfTwfeXBXZzbGLaIvMD5AnGTRPhuF
qyju8bFriyZugCYqi00z7+Pc3PSMWz9MfdrILwYJwdftxvk3QldSGf14kTniwfbJ
8RG0NdSs7SLwMDyzy6L6qrnTWMU9B/cMZZ2denVgCPjK7Ln24Ri90i3fj/85EgH3
dd5pHtE7TYQ7/Zl9S33kCwUMdkh9mHPuHvkzOoSzioGpVaog8OvpJL7DdQ0kF7E0
lUyIMUY35bpyHlqs5yUh4BbdSShSsESLopS3pMkd8OpdLiXTU9GVEa0glRpsAtgQ
yCYBKn0I7WQYXL8+fTkbMdyXOVfrOirKJiOuhsTlHDSpPpjJLKRiy+JLoIslLZYw
ff7S65nNjPfweeneLZWkmlRUVfGDx2j3YmsiUxCHrETTiyOvm9LOtJaT3MgaRDmA
lDAkeWmqyJTgJIpv4yW2AYpx+lNOzwnDy+Pw8IGJ1mcWMElMDXorBebrSdYRz8EC
d5s6J09x7gxxV+d6pFBwGidLH/xFMGi773B3jl0py2ga8J4weMp10Ln/lNp7/MZw
uNzwbG802EtHVT1m0u8bD+NhOhblNtWfJxxTh2/HcDpnQuJC3+aU/NYDstDMy2/3
Q21orcxvAAgMdmOx/ubAwulxCsMJsv0kDdyx2a5xJJFDrHpozasu5QMdPsIHqQGS
kwYcOuEhSDVwxryFnwskt8N+YEdHnrrZxX1pjhRZ0WB20LbSz1gD3PPHV6fGiY5j
1eiEiiimkC0J1mPz973SP48+sXN3iqSpsZPPQ658qp62R0csYBaCAkauRZreCXaR
qSlTfPpZ7t9O0OkDCBAmAiyRuwTcyucuGZOMVFGclOuXv9F1knzd2M9dqZbI2LMt
BjL8rjMlJO93N2t+LbKnvHA58HJfnuHA+2ngBCjJ/l3rvOxq1mgImi9yv9NYIQVc
UVPwqUisc2wolPNYVRpEK84J9MV4wOA2QnwL11AzBw4K6ygPuAbtF4jlRhbYD8ms
qvxLZ03Qh45fVPiAh01Rf36Ez1Fiuy4BSYWZkXKAdGjxQo4OAuukLGeKAMptag7I
ZEIU821eonhbctOuVDuCX8IvBTiyvxix1fYc8qJfhfGfV3h08GQ5rw0srOpj8Ef8
xyWT2ursxIVdH/bvHechYfql0Au/6fCNUED05zbHhGu42djQoiasP8rTLLPHHt72
RByB1CPD5mI1z9FdRRLiEZNWpp+Sc2aqZkhr5xcGgrjSJ8h6icmxNe5QWjV0BGkY
35PwJvR8yU9OLgYBBOy7RWk3hOycxlBZveLoYJvSuTR2w92IgxBllcYlFfKU/6ti
FQnxU3f5iR/19vdllVPFgytzGduu+mW1OEgVjQh1kDhxRbMOE16RTbAMEZsYRj60
DVn6/ffgRBvEy/5ls10lHQpYRWuzHGA7xjey0xVIPD2wJPQTLyo7naJuqiusxDbi
syfNPdVGBKO/e7YZbKG1lq2K9RlJCETiVdmJH3/GXA3av486tu4iKa21MKk8U46J
AhXYuyOsmaEVPwAVLcBhiVWnDCEiZ80b2hPZYkISv7ah7/bYO0hRx8EJK30aUC03
suiJEQPm4yVzJXqtQNuKu1pmu4s8R5sNBxkxitFlaZQcxj7jdVQCj5jjYpUfVWnS
musva5i9kNiMLT7HOrZGARB1uTWg0bDU+vvO6XwIAKJ8owdHB4NorEQRIgfQfu94
iL77g4GRirfw3p0WICs20Wz5ylkzk/sHbetse294mZ6+I2p6YDt2AbgRs5AjcQPD
NmA5oc9xczxKOBOahkESi0lPGCjNsSeshl00pF8jH721ia5HmzGJ4rTvWA4M6t2x
9mAglW2k77C8c55ThG+g9EPWq0VBWF3IFzsPLRPs/U6bxlU52Bqj3kK6CgpSH24r
cAiinEfusOzEUUCpOVijs84qH4tT2COl1/o5gvHpwBXgKZCYRPufHcBjJUDwH3By
fiKlzJ9c7gCM50O82Xdx6UxTwO6GngFPpafQTowfmoyBanI0LzQDi4YhtmDKIUm5
GFImTXVdLEK4702K23YJfhzAllYtpTdw/1tAaZzR1kEHvmb2U9tzKwNWPsXkwWco
iJi112VCT/xJavJoRlfMmL8VuLHfVhv3KrV7T1POh1cyLBiu8V5ttA/A2lw0ub/S
nHy98qAH/e29SK7r6EWirH6ERifJ6RwO2kHVMZxqepG5PMAIAuJIl7n7/oSoWsOA
pE1U/+jiU/u8pUpZya1q7xA2QjtwpSOw/oH+RXE+CYKkzNVanbrGGEv/TKEO018K
ExfKMjv9oKSbLsDvz9nnbRYOtNnvte5dSEQWPhEysHsTj3lFIhCcAB4lYGjyhOLe
LshLjFkzp0KNfxSpu4It9u/Wl8oRdqrbzI1D6aLBwxbdFNZ5ZeECmDKt7Y0pthuR
PfXwfDMznQ0kaCc5ji1557eOoa1AUFcJh3dIeNgK9URlPSZ5n0n/cxGyPYy8ysB7
fe62MoRcwZB5IVzBMd1tmDoTO34e6Rop5MPf/a/EtzMWFOc+5LW2n6gmLmvbmsTt
0TME92kEoy6HM/FuT5FVhslGbmfWVo0PAYvd40B62dzpWBR6TAAqktVmsWXuO3ma
36VxyFfOHVFijy7HzJQAB1ri0SVujQfde+/YHDTrFgVOHWEJ+3rzvY79hJPlFn/t
TeF6j1DUxeLzfwS1I/CurL6i/Wzy64LluAXoGvLoKfWCKBRGvrW1k/QLGO5zPqDv
CIFPM3qTcRkLgcKNm/opt2sWIcYDTUjFuivXEdHfWCBB36bILaszGO2tFtH0Zkx9
oUNY3krQK8BqbesAA3WE7+tYUZNodJ8M6dgITEtBN95KtCjY4hw1dlElireu39MC
FyKiKU7ZBz07BUUClJ8eEY40Y23FCDz6zHoS/8pjYkSAT5CaVOxZvpTVePpSE00p
wfLegolOOQtyivr54FMoDoFBGTM3sP1fOMu7U3apSymhWjZPiiAM3qCZi+pxGPTl
cwYPh+SyqAtToHxM2PFcalt3BECOx6eDpw5VFxlZUp1+PJFwwddUpw6UyzJZQ2Et
k3Qzd0gXmlHWJ0HnZLH5NW20Dj4eDXYfmWn1XCtdvgFBn8AibalgqgR+7Eo0X+7d
vKEmJ3kZBF3KSV58dszwLUsHWG21j0HSaOt3gzIWOE/Yr5ahqLR/jKoxJH+1O5Fs
vISUVAdbCq5J3BDjsIFagnghW2NvWK1DPDLqwzPYLMHT8xEuXTRnzT8RdmNBxxO8
l8Sg4lEGqFLyShHCXkMTZqrWOCU0qjyncF4yTWmm6WOXySSvLuG+RO/DZoJqxh1B
p2GanfCtWTaHNlrF3dkjBKnDuJiH4kQ/gcRHYs4aVc0uOXRSfOMVVMEoKftCoyoJ
CvoNrqNojdZ0j7c3AL7/qjJg2DFghtuCmSNsGELtSWiwkFda23QybYF28SdoPksr
Zj6xf9LRTS30xvC5MZnoaQDrLQK2/bNq88rTc+hNH34tJJlMRIAOS3P9IImApPuB
RM3mZU+HwbJp6V02AIH54ITJWSP0lawu/sC0wOLEUNs5EQfQXm+NbnJWnMmikSnk
pjXWhg4zlXsKXUtyT9H+y3e+REITDGmAJQYCpVbd3W7A7MsZEZchEZWMi6WZTGGe
gIlPpWMNQz2rXP75GgXLdiqYLKCXMSz4MiDa9juWw0Q1Uu2p7tE1a85S8hpBmOd/
QPKg+SFAQ8fy1ar8ABR/u1HK4n2ZhIu2oUR6VAMNfPmYeWbzJ7HQDe2pV2FFOuY7
EpaTrOT9LX5DbGgJP95rBomdYj5jfo7LdbTqUdkM+OaZeRTNIEU+S8nuT9kymqHs
s3sVMRcERgPdBLWNqp+XIk3iR51svYWkq/y7InfMZJbjn2sTi1qtixrEcdoXTO2d
U4q9UZcnflnyGhRXfKwMxglNy8DWLFS4weX8u/KNNlNhJKJ8qXp5KVAWAtAB6h7G
lZHsyPDOB0N/3cgvzBxIXUHTln9MsC0NC4LnFNFewpGysId4oGvu5io86LSUW5vA
QPCXdby7NxWG7yqYeSh2wniSy4AbAjloKpbuPLSRZ/cH7Nf+t7QWQrC2f/5vZ9ak
9f3tlcO70pc5dv3WWEFpOaJuXq9+llpFzAeCV4gI7SPzGJ9wIoqxCH1H7bUFYKbg
Xc8ERWfwp2uirle3Zwe7gAYwue/Wab9Z4ezJcD3i4NbwMnvcPXXFNjy5hxcdrYPT
Bl/+rwaiQgyTb/Bnuc+8chQrtxRfibuY0yMbCf77unN2TJK8Uy+K2ehT/+L857a+
5h6GuiD/zkj9Payv8alYZu/LlTXBjil1PC9qTpqY9S7bRpzH/yaY+t3+FbakRa/R
OxJUJ6ZKiTSu554FYgSMIhhe++A7CGTjeTMlsPegHjD85YqehKl80BVLgfqrINuA
I6Am2t6+uhWULEudlhj7wiiKKoDPpICpU8SmArv/5ZmFX/RTlWmFMy3TTGc7IreW
D4dizWpJ0vU2nBgN6l4THtwmNG22LxWDXaTyQFhH4vm+mjIWoVMFRC2XjvndfFuQ
b9Q0Gm41BKjmF2RVj0Mwvk3VoWXlCwNJg6N1cz6gAgNqUTfw5Io2uDORY5uzb8r5
lWH60VqTi8dM2t2MMg7ViBnDLKThtrQE4J/FMmpUg0H9Xgetn1CPuh6xbJ0xwccy
arc5FiyP+P9QaRyIY4rOBPGLlkMa2S4aFYIhH/GU7bVaO5TGxdmgAHHCjhN2j06C
24edbt2Dh0e/HHPUVVCarAeqn7IgokHX5W8xmXfdrZqq9AjBAnQN6d7nI+m2/dlV
6L1hQEGVWh3kT2tlxh1xIqKJKsHykNpa5mVrrlOP7iksgo8tnjZt8NHpamve6tW9
FjATYozUl5eD2CLbxhl7aIP+T5XIH7XflSXLII4wIoVc0WjAze1pWetg58LoyHFV
PSoKDHoqB7i3h95CpT7EWbjxGv6NzbbRk+Bsd6/aeNtq0g9F5V8/F6ScDOhff1zj
Yd0qf1r3O9LN5aRKzKuGHvDECFK30qd8Jz7+2OMhzCCBC3mt+pccKQZxZXGUFcgX
/kacnDoKHloq6AISgL+tC5nBePmljKrYWFHN60aVnOWLHMzd+aZVI931fgLi8Do5
NoTStxL0SsKM2f6Kz2BPYROwGQEJYWKoQAO857Exmf05FhskrI0UEwazVLhkT7iW
NcTMCUtCYLxVXRUZ++nFGcu+5Vs/xKD8eKwd9mAUpD2bZWS9YiMH/7+nVqi8PBHX
+IelBOStv219G0h9ze1b0jrYaWOS5kmBkGadntzx+cJBQjFzZrG5SxczkLJxKRMz
eHQ37Tno1uzin5MP1FwOP6ZNBzqvJBh5lKAMZIoi5+7/268EGb8YTNkKtGE6QEKf
lEGfov7UPHekipoJBDB8WUmIYEif4G2PM5x+1aB2pnTnT/wyNTYgvTtZidFqD2v0
jQ/pfFfcPpr34VrvJHLaupziYHLma55laQh8QS4vwYEySkBl7Wip+TR4hdE+tM5n
eJlWRHBAcJaH1iBkbMFhiFsdIDYjNhsiZNd9qOM1a2hU0eVWU8itq1qTZBnvdGHu
zGP+frjQ5XJLzTOVlJbpcsy+yjQjqtBkbrGlF1t2ToRpqnQVO8TgEJj+o5iSaiqn
UYW7viFCoPif0+JrMEq1drY00qWFaZvNsOqBaiN+dZMIGiOx1Wt/eVV/4RNVnO8R
kbq0mdoK+hCCfsdYCL9qgzdBrYCVmOBLzoF5UT0oONhVKX9od5oTG/+mVjFYToCr
RwRniRCYufauf8smy12YIjv/vRAkRPmWDurA2X2UPN63e+Pw8hstpMquj3ARen7B
4Q12ppVbJFV2gUoDqm1AZ9AhCLTAA1M8xWyXuHtxvutVW3QRrWiDLxd33mOCtGQB
hLkjgiC9GeMrDXAxU0r9nLlvpggfnuIN3/GrENkWQolLKClWkQkH0ysFEcTQtHGU
dkNDdKbyrsfwstKSSdwvTy93O1CFYSuUoF13+JyUC5RpqGY/VPepohJhKUdp9eGc
pkUbEIwo5QUn9lOWfOsMGbwr6w63d5ZtLXQDZrqCT0YblmJbRSwtCjQU1WwRPneG
8shWXGZ9VUwMbzmamZ8kcplbRNcC0b+70oO92Whqqx21ZMHiBy73Tjg6WPIGaLJE
jWn0IZ9i/7V/X62915gtE5Dev9G2l5nGIvZS4fQl6wG5jhrM49aOmptfwZbJuzix
pTqa398D67LEtmyX0/h7bUx55lHL6wXDR9EcSIMwrjh2eIaZjAYtcJbPSgHOO0zr
2ArfAD3Ia0uWuS4qGdjh+OcHWes/bkaXD9SzBRS5OFYAeI/DYz3qdP63AafakeBE
c5ZGM54Merd9yaj3+ITk1WOlKVngcZ/YnWkgmT7nP2y5Nfi1Z/rJtEeo3Ed6yD0l
04QgCxa4Z94vjy5cdB2EiLDtUt06s5ieuiA4DlzlO92yMgfeGJ0mYDPNggtCIPVj
R+A9Jxfe0TZpEWg0VFlVWCGg0q+9tt90bPlnkxK2as4kZVnLn6aZlGhnWp/Jx1F+
vU6gEiVyR1qC/flAtbuwruGVmo5EfOmxRka03dJzahq8pNCb6+gpQhtqG29pNFG5
3zyYKfX25QCeembUNCgdy5caj7hSFlQDOLW0qIw3Rh2CDwAYDJ+3lToEYSU6dA7F
c+pSGdMvspKDNBRcdryOJqIaQFyjidHOdM4C0Vd722Ycy4nJ6zJq6szikH94teYA
ZdjhEZeBoGNOd1CvpCrVD/4DAA1+RRoWrr1/femwCjwPq/V8dE0NxhxEYQ5gEzDr
iXYWUhKviVfpImSQGV8OpTLEjgfQyipcoc5D983+jchoo51btMUXMulPfsgF2mSE
AfRa5BQgurex3XPa/V1OnF0rm5DitJBrN+bSMvfgkjpBTz7syuuRWPw1CUE1h1fV
xaP2Ty7P3Ix3AzWv4L3tb0JudZlcQdklCIGsBNcqDlLAycO+wINkKHQJcGMsiVyo
kjOcirBtWuuhckAjZC8jrwAuu6Q71rrMXp2BJOkEm8fEQZBuYZea1+mPlbGioXGb
X9Ydt6iN0eDg11N7VjjMbyLxspRAKZMqoeUu/p51rORMwrbIP/YO9WsUXzgNn31k
WYzfWLh1qJtIgGKs0SybiIMqwTm5VF8KoEsqcSRVZUanfURE2mNmMfCZFa1BjwoT
ftxR9euC71FjNMJiFL0x9DaSwEzx3uVTUMdRIXdeykwHzsFDkQYkMuNykWgNALpA
87QwlK6Ro3CYCh61mboop0frp1vK0GSjKRdX03UhLyQeKu2soXQ+w7m12+Vxn8DP
AtZdi3xE76c89iMOf8aN8PLK6lwEA9UkveUXH/oBDkgI41kNh7t1lHC8zJMXwFNS
L5XPcUvrEh2K7Msouh66rM6xL2vjsj6FT0jk+B1qC36C6S1igciNB9ILofRsEUZ/
wLPFc9uoDK+MgItkKL5GHMgwLYjzT1tHjI/kkHxZOdJnjGumcj/HaUebDcb9EyGV
uNVY7XiBSWtmZU0fYuu7Zylwbp5JiMca0qz7Pp4Qh2ZMSXhwL02y2hLp8FMScQG4
u2O6WjfJrFsdQ3Y7UU/2g50hN+153Gf+pF627RuFUTYgxAh5VpbeX8HDT89o1/1k
ObGk6E4F6gAVf5ONJ3yHTAJjiNPazPIFWNBOOG79szMW6+pRwpMWWYuXkJRWPCjh
Gp/yJ/L1SV02FBX812qh843/VIZTTzQxK+STM2kRjqmdutbzaHUEEYTemH+CIH2o
o2k2W6FGyxIPDVIpz9z8wv5ROeIMDJzJtIarIh0XT6QIjRpVjwcev7+r2cskeCd7
Hh1yZMZPjcsP49RnXXXWde0FSxOpJzpi9DzpoSl9z1Ps5eQHEDA6Ml5r7dxPtH+z
zkxVYUX/KAZXLWchn8br0HrnV4pkIHxHO3Wf4xXW/D4jrDrYO008FfgAnLYBTkVc
fW9lI4bwTz//4wvARDQgo2//SalpAOw3bLxc+uEURJsL+RZi1oY28ZOrPIBvJzjs
UGPAKlmjbEzlfcVrawltGKsfFH3lRfWKWey/4e1+ZH4LnnQz3eH7IpEOxGQV3gAf
OV6KCxNZVbCmvzMbjfJhKkBjUVsZH8OS09rPXQFdVBg0KNyrzJd3uNYSiJmIJCJQ
tIKC1dowKnWMMvIrQWl5R6sCjWkz465GL5eke+//94zgnjtOZVVc6mZ64Kxzx/xT
MoLNdRImMOJwJtakYVDc0CawQ+c0BFIvNO6Tht7Bkwa9T7x1d4JbeSVJ9zZjeV7T
hJX1ZSKPgfWj+hpXe8ktrSataVjm4mNdK5DJxP74ODM6yg3TRg5ZycBb4vhH1Mt/
hwpH9Rdu+lrdt+nZ1Lod3KMgk5/F88Xqbck9pw+2SqmvdPDhFwPWi+stPNCg+CHp
Xl8X/9ouZhddZhZoKJ77RO4blxzF66hgM5i5VW/D20+/RR3lS9DS6SuvSriMrM57
1iLaxqZYtooDQSuEszo+QSujyMz0T5q0eB83GeXbAp8GUi/PXlNRjl88bXmicXmU
zX2ej/p8TxF68NQT4XKwJIxiPLpmBXQrvHuQWz3hYyXhRhXeRiHS+2d8D+AhvVJV
+WTKz5BNeVXpK854dcw4Ji0a9zRSRNVcTjdzUVD9JfzV/ZwIx9taeEnWnZSGPDiz
GCw1hgdCSyLE+GOsZ3dNikO00bTs99ZVqIxkGOtHc7KlOUg9kBO85sCkQWuH815v
Y6Ujq/C8GPS+sX0+CPNhkJrrjzxvBY4ifeyAUKmd0Bmk6tJY5/Y7wTkLNKNYSCgy
7dxKR47eHCYjtGFVzqB1uXFmatV6FirDrUXc6S7ez7HUkMnTx5awcTDbUvoYt3Hu
lPpn+hx39qpikKidwy6FZ3QcN0wL5MVxsWW6LR1hQte2axEQtC3S5XOJRKnpfLSb
9yxHpW42XC7oXnl1Kg2O3AF0TMxJ6ptXp62airn6o44vZ9Pa3p4g6XqzGrkYBWtx
NOhom312jzvnvYisP2lRHTpBrEVhBQ03MNj2RbiURDbHCL0JBMUdLBOhD9wYM5FK
uoxK7q9ujOFeNuVy60yBx0gAJY+aB5ZfOf5r4l+aaOE8wUbPpFN///1qGx/iXG48
nhRVdNieetmo2qed9vw6lsoMnif0LUA4i9YUXjY7eVxdYX+lef5r4arRXhlrwCpb
kn1HzksTfhbVSICUEe1yk1aOhzxciaRq6Ryj8Je7ssvTmLY/nUG/+rH11zk7OufL
+++4zDz0X8jNQqTjroMiaQZdBU1CMFj6U774qXbt7OWFPgfRU64b5c4srLwnzn4B
0x8u7pn3S/VwFf96x3j9e/ZRJ8c2VUcrLDGhViRCQ/B13+PzRXdYMyTyWo9SX30a
WWqaAPm5BKt/8MoZgnYeRvywJoRzcIjJXlVgpLJnwkmeEYWWnwA43HpGKHRQhx4T
FPubNabj67KGNK4XFpLLS4bN3NUpSERvgr5DnaZ0vMHnnqz4P0Y4rrWAoVz3Y81E
hA0cknA2EKZw30oXS3eoLhtqGHLPBcHGVvrVmui2CyN+yJlWMla6/o/1AY5KYi+6
l4xSz8skJyviHz1FcszS0Bz8WU95sK6ZVLgScjnErEbRbcYp4P9PK9Kkv5+SEoy8
Ob5QppwqyUmI27DyUe7o3EZ7IAhR65uRBRj701iZpdm36eHILwyaxApB0jdHRfK4
YVRDdMZHrIrgg7MxAbh4wd7YB1AxwqmjVLq1XOPrphG5xPFYnT8879xaqSg7Z+6c
lZnFSpwRR2Rjp+ugyyfJSajsmEOPAReBeq1u7cdZKdTg5e7mvlmkg1L0wePkgs2S
cRBcvG3I4Gg9xyI1i+UT487c6XWQt8nEYznsX/rs+GlroNCl6v/JEJG9qcJiHqfY
ParS9QBYyGw/LYEAMSYrJkPh4lChzywBHJhKCKDPjSuT0JD6Ip7PUbdNsoObWLq8
nc31YgiIrjGYKUrdhxo04NnjWbXk40TRuvRcd6y2TUQRqBfu20AM44seUkQZhtPx
PX+oP3YwclHEWF4gAP0niKmkT+vSTohkU2yqYycdPv1Sz6xSD2/q2YqZUBfd0zN/
NlPdeKKUoxxTszyPO7nTukhHQJDTiJTW+ZrfyrcwTZs33eGNmukYFtsV1Tdxf5uK
FkBuegyXz8BpUh9tmgmtJ4ALAZXZ6wHPuYO7T5kWqEoRCLPHl6Ie6Nh7dmy8kJKW
11NMnmXakv0os2pDpeUc/7tpHW042Bva3wfbL/wg4F0LZ/nd4FEDGe0ik0iL1I0N
aWsZ5a/FjT6n/eMuMAi+Ydzm1VN0OqO8gnRW30gvGIAHR0vWXFNKRnOAC6IzC6OV
NVcFf7VLXhAYD0ekPtdydgjdrQkKZr/mvN/NOclvqilmIluQb0c5JS4FfSLu1dxk
4ZkafkK6j1Icdu2O+pRexfLbTOiKbvaQ9aPhl1dI+XFgMSp3qSX8Srg31H1dSl9M
LH6MJFmcdeIkOxrdKBZmhAugqLnrVOuJRDtJqudGcpJTELAX7DC6l1EqL/kQ99J4
RwKQCPpr0PyZKVhuMVEhGgaWE3e5SiglLLZafeBQPjVeLSB5TWaGtj0wNfruWAnm
05EfeS0/7wliPbny2usBZi24eQN7njJQ0Mv/Acc0PLTBqa89215n8VfUP2CDUCPm
MvxyiqqeQHwgXQO2MQMtnmKKPklShYAoyBKleK2/WTlBNO2jX49Lin27ULfNoi39
YGWJMgNcR1rODFUAuRq3MGr6iAz+Vh/xfI6lRhliUXuzGZByRp3VmlWj+bx6Kwm7
LzXf3qNnT4plZJ5DXVt5KGRyTdgQURNP3vuCnctMW3XAEThGlhu2omazWdD5h2PV
GWyBqbw3sUTHg1+V/NDoA71P1Sj0OvWgSLZpjCFmKJsdw9uqFMBcuafTYdlm8tKp
RLavD2dPXqU+mYx3OXIG1DjD9pwtzCv/l+E+OVyjUr7vHkp/assebbkp/SWaN+FK
iI0df/6lX0CisNzbkiu1atxSfa5qdv+pDqBZdH6xZCNWJ2DibqVo18hHnPqQnfJY
JG3YSm+sQ9cgXX9GkwF6OlhwQGizfAG/uylvpiP7x2p3APoRfkEUJ/yiG5u8fE5J
Oy6Ia8kW1EmFVUToeekMmB6JYeUSG4PuQ+/geH05zWd96/Mj0C8Mtv9DH/Le8tL7
wBwXbTw9+aNfW8mjbvQwA84Tqx8p1t1bcSzxq9wEyclPIfxtF+Ci3opRL6tQhiVu
ZqfH08Pwd9VrqzBs/Q+9P4wKZeo6FdpSfIZCEGWcDqJYnLYE+tVy0XVMYYoFQXDh
c+StNn7fHBigBdAbZ3weGFojRd9bY9YyETam0NIpuvgNfLUP2x3htoiMcv1kn0NS
+VZ7xUh8u4kMU1ONQDhoQXVqehjeY/zfXs20IKYE8d2IKup/EBhEIx8jtZyz+QrU
Y9PdEd8NvSL9susZVrXWUNghO6shpca8LyBoY++xEUbGrGwCDEYZ3v6uLJ/8C8xi
896K58plqx9IoRAjGkeY7uVXCZyu16ArDCQf5+NtPUupvwmRZAMHeEUPM4RdbiLa
cBWbfM9OauFhqCsP+ducFHreaCgv73yKgW1rw7+px+1O2R2eGu9e54KnhsxIUkL5
EaLg8gRVBsRXwvhjHEpXUiDrosEl2FPgQcFRCiDSZ5YH+xXNTblaV6LqBXC8E3aj
9Tw7ciNwh7xBQci4geFxXlAVrzO0OPNNww06ju3un6pMeJZ+rxecfeDygWyWuzsG
kQrUCgWoilb2qquYkJvb7n7Qn1LXw67SES+f7TBjJt0NKOKI3LJ/k6jpCdn2Kf9j
xxEoSmrr0/9V5tTbtmJ/VwEKml48L16LWoyCcr9Tk7N6B1DRStCpMj1f5Ir4A00R
pgTKQcZX0z944uYLhF3ymJxqskxJVbuT4HoOZHy7hk0r0Sw0k9THco59u0CL4VX3
vWUk2VDWLodh83DYcFD38pfzKkkqgKJxFFv/ZM74iIrLnJvrgGZce777mxM8HQsp
Yb1+uZqAE8SYtRpFVeAD1dkWrtewTxirO1Zlxad+Xvu4KiPrCV2Q6sH/BCoDERCW
3EYRCUYQQ0x4yKtpyG68Aly4zItPZOwktefaMD+c1arx/P3PRj3+VhVoUOGaKpO1
/G+hT/KwFK2qR4tUiLoJ47b/Wsgt3UcBAwVzwXsMyYVNTFtG/aNQg0hgx1ufkVHt
eJRbG5U5GMLJpxMINLtMUabFqzmdN+wqeI022QmszA9256uYQ50oN9uyn4e/V7O8
cKTvS+JSyDQtDQ1OPd8cTZVGvG8WACzSWPXx5x8rFSfhMQI42JlAUBkvw45X9YRA
I4SkOHYyTSdwKoe+5T/j9ZiMRrKdz6F9E22z0cBkE6g=
`pragma protect end_protected
